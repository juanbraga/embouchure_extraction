BZh91AY&SY:x�`�5_�`p��"� ����a��0��U*�B��im��JBن���"(ETL�I�[RD�"�j4-�֊R�"������M�JB�P�U(�D��� 	��R�UH �J!@�D*�� R�TE ��UI
��R[T*��$D�T��g
��)B��Pv̶�
ݮ�aw5V��q�:����u����5m�,��wq�%S�;���v��i�Su͹�I��  �r��*�B��ְ��ŧ,.���j4A�%6w8��
滎��X殶D�n���k��i7u�F�	�5�l��������

�n�((
�2V��mN�vZӣ+��vݍ\�9*��s��F���.H;q�풨0gq6�w;�hhc�+Mku��R��P�%�J�ts �sn�]��q�Pݚ3ur��wg\�e*ma���+wq�t�Ν�qk�*����e(hvq�u�]���hJ��EJ�RGj����9�75Ͱ0�.[�Wl͜Μ�Xk����WN�tR���MZf�rs�E.��Gm�[08R�)P%A@�Aي۫��R���:�ɵ���*�`gwkWv����$«�w����R����՘kإt`*��j

.�+�u��wlmtp�F�d,�nUk]���.ҋ[���j�(�YD��k�m�mڨ9M�m]�iI��U!V�b!RUP�p
���\PiE�r��wիnf��fv�Fֶm\�sM5�&6�-�ͷ9ժ�*�s�m&۶��@�� T(���v�up-N)���������dm��R�g\��Z��;��7d�\�5&��veStJ*�Qʐ��QHvl3Z��J�����Vmڵws0�Ī��PW0c��9�F�q�R�� d�J�     )�IJ�=@i�� @4 �@�)�1$�OA4h<�MiOj��	JT�     ��  �    i ����&�@MM&��v��OI�iKI�&P������t�Rվ'9��u����TU��"���DEDT� �*�Ud�EAX�� Dg`�PDi�|�A_Z�J3�~a8������RW]���*P	I-V��It�n`�Cs&�70��t��6��dY(jtB2]�����OpK�롆�R�X��@f�Z�**e�Z�£�ֺ7+�����YN����;��R���N=jd��&���ńAWA��j�Ӧ�M��1JT2��]Y&Qz�Yy4�;���)�H��F��P��4�X���@่ɋ,��Y�;B9�G6ڏ�D:�&h��z5@�А����j�R���ʀ�1�,УȅG���퉕c`XA��m��������ǣ/�B��Z�ޅ��K�q�0�,4AM�����Nf�H��fFƜii��
hKdŤV'�%�B�flfM���X�vkb��Kf:����[NZV�6S��#cf��6'�,�]S(h7�I,+�jJ��;�䎪��4,bgn��[�������D��1o�	�g�����z�
�t���f�!p�$��EX2���nd�2A���1��n��PFcgvJj���Ә�[%��S^�{uh��Y��6�&%�S�-1j����N�d�@��K�4k+I��d둊!�N^��k�[{Bj�X��m��vobk��nl�d�;��Z�L��'�R���@��7�uXaںP�P��+A��S06�ʥDm Y��յ���5��l�Jʤ��z���yi��Z��	j;L��ᤒ ����y�k&��lku!Ѡ�e�ꬹJBd��ڵn��Ī�\Ǭ��V�{����v�T��M�&��;^*���*V�+!Y���%���n-[Z��ѩc"�'xӳA�$ն�9)к$@��P���$n&��s���[�M�7,���iy�'���5�tm�*#Jf!#��_"���J�g;`��)��M[1�4�q�Z�]�)��̩�����YF�絺�3�����GJ�i�M�EZ���Q�Ni�grJ�Ӥm�?&wJ��Й�Vb�b�f��{1�V��)�	��,��!�"�
��e*��#ۥ���6cԀi:
aPՖ�-�h#��P�0��w�v��*�f�dp�U6U�C����5cVK"��*�V�d�I�I\�"3
uM�ƼouTL$KY�T{f�n�cŅ�=ڭb-�)���<T��h-��)�F��-岯����ٺ֞g5�yJ�DeJ #�&�B�+D��#�l�M2�FИ�L�+!�.�N٨i<@���ާN�zh\'n�&�s����rɉц�'w�֒�:]�s\�<-R�kA񠉯*;')AD���#ZP�PCH��$��_F�@��4�ev�K�M��IFh���43�s�o[ۘ��9�;�deR��W���Q"ܱJ���铤}L���Xe�ۛ8��J�
+��:�sSA���#c���f�-חy��������Q��kr*ʕi����k������ֈæh���a �5�؆�\�V9U�K7l�lT��1H�+(�ّH���Ku�(P ��K"���X�nҳ[�����Қ��Ԭf+��^Ba1І�&Dе�j�1���"�3`X�0閩cd#$���*M���9�B�Ȼ�Ō;�35�����9i$���7Va�b=�b",�h��iF����`��N�-%}y��Re�̪�R����$�E��¾�Bc�a6e��[j�ت�]9����5��q}*�B�v�Itop�0�g�1�Os%�Q�]b�3��m��z	2Ň�k�C5�%��F�7yAӈeďێR�vs[������WWR�Ŗ�<J�JP�3t��6�vȼ�n�RѪ�婱�����b��#;�e]������r�����d�ϝ B�)�&0b��g�D
�9��*,Kj۩p��tmf-�����(U+¥g�+QI�S�ݍ�yYs�ª^��L��N��#Y�6��acYh[[�Y	��ߖ��G�A�d%� $V�P�_ A5("j�Q:�Zw��T�f���߇�<��,b���Q[!	�g,T��%zN<�8����� l�7)�a�&���$�t�~ �E
Vh����F�5d̎��h!
I_D�?QA�_|6�1B��
A�4�T�&�h�;l�l�n��l��*_QF���|���n����rܨ��D=ԍ,K�oU�Lӛ��t�ԇ��[J���pM$ځ�Q��=�4�yi+��m-��V��!LJw����W$r�,C/~+//Y�wL��.o�<��ƚ�_0Dqm�`]Z�PQvU�x�[��1bVI���Jm�
���7r��Ў�B�U��r��"�AL�V��F�u���wg>���[IA�)4�*�ĝ�m��kE0�l(7{����d%�v����(V�ݛ7c+-���K[��ѭ� j���}�e�#6:0�٢ho�Q8ș+t<U��\�������F/��� �;�򭖅L���r��cR�ЬemJ6�,;w�n><��v�g%�V�a|�1��I��Z;Y��_9cP�E��>��®�`����B/�y�R%�ϑs��fF~!����G(5v��wOH&ȡV�o��3D���L�W�-M���j�Yc5�- u��f7�:N>��b�s6�4�����0"kl��t�-mZM݈%�Lm�����9j�f�ڧ���wv�ڳ���	�YEh�*�X�6�-E\hX���`V:I�q`/�em97i�@a����Ef�1�-��G9,5�W���U�� !��̖KG�֐����0�M�#ӂ���Բ�+��d�f�����f�L�߳q�M,U���RY���jO]�U˕ �Y(#�,�+IW�D`�v6�������ƍ����Am�<u,l�)�A�[E�T�b���5$JY�[yU/%���m<X��j q٣b�4�O������X[��'B.�R��-H`�R���2�+�hn�b��@1f�)���y�э޺���P:"�Ub�С:P�oZhcxu�R��xY\4�.Lz��٬��"�� lwnf��X4~��%�U�?�������I�b�R�0�U`�mm
/]T)R�@7i1�o �P4��#y������8����s���~�<��`T"j����n�o:en�[�` �3m�F�1V���l/�$a|�o�T�?j�>f�H\k��
B4F��,��i�Z
I+s�Ak~w\��a^38i�a�P���ȉ�1���P��[j��#_�@�H��A�x"�B�U���s
;�P��b��}���s"�f��˦�B���O]A�1Ex�Eb�	��tU�9��>��� �� ����&
�0ݢ*=�EPm�\�I�F�Z�n2�8v�	'�(��"�?�;b��m��B�f��P�R�tܑX(jd�.�e�x�Ǒ_*�Q�)��HA�QZ�di�:���i(A��d���Q�#Bj�f�&���A�UkC���4�@�+e��	۰B�
�B�$d	��������l��i��6��.�ؾAF�T 
c\������',�cP�[V�n�m�r�����5�wAPamR��浭��5��Jk�Kƨ���`����r�����l�	��{����(���������h�-�?U|H'�5�JW�g����dMP`�-��
%:y[(+�E�����X�!�F�j���ݪ4����g���CX3(Uƨ�]��o4SmN���ݩH	t�$�6�9�J�X��I�pm,5_I���\�a�Fi�ݥ5�N���E��%��>4p�N�_�˺E^-`\�	��UHh0A���	���i�J42Dp���U��n�6����ڒ�M��
הVnP�b��X�l����%������_Z���{+�T�iH���J]|C`�wu#���煔�I6�������ZB4%*:�T-��<n9�^c��cf=�sV��FΌ�0�?��!��TŬ@Pp�_f^2)4C[z�A��.��8E����rބU�xe̲4���N(��[$KϮ�"�"�a! ���ir�a)�%hA١Y����V�7q
nX���w�t�[�Y�޴���J]'[crl[b�`�މ�AV?�B+.0�(^'4!%*,2�����a<#\�@�5P
 BN(��f���0�� ��Lk�QL�sETA��(���[J�Y����bZ��ç5�$�hb�5���U��X����H�c�[�t(��J�4�ڸ�L�y���wsz(#�gP��Z:�IA��
��[X��b�h���P�-D�9�iI���C� e���8�k~y�����e��Ȋߥ�2��54��/M��(��dts�p[�)\�X!V�|���LG�>���tA ��ʉ׎�*Q�i��&�n�j�W/:��N�<��Z!Wh��T
������������r��@��*�c	0�ت�?��o�L���5M�f���	�`����0�8	
5W���s���c2J���)���o�7�Żךww;��i8V�75ݹtK�ܡ�T0Q�
G6�WT��M�t����w@i�E�$�u��j��$N����\�sdZ�NU5>lLʥ���˵[��N�sc�f�\����"���f���k�@�~j^<a�Р#>�̶C5�O��
&B*�'d���������$ ~�1��ڪ(����K@�b2��1u�7�CSݗ�P�6�4J��2U�ݡ�K5o2������7�0�D�֝(�Ƌ��(�yt&P����b#A��x5H����a�Z��a��@
���ۓv�Z��d��O����Ki�! ��,F�t��d0�!��f�Yj�X��A�魔��[��Eaeӂ�w7+3)T��*�p�x$��^X��ʓ������q̶v���pi�5��{�ۅ�\�19[,1l�/j�R륪7`֗T ���i*��{��I�b��{B
�}�S��E�@�ׇS��R�(:۹��T�f�SK�s6�d�`f찈m�yR|�>�9�US�t�m)��ɭU��������#S5,(f�R��R&�Zkhd����ۂ`9B��I-J�	P9������nZVޝd�s��������5���(k,���(ځ�O!����h�������d��j��
������6�b�Y��t\��eg�X"L�hdv�� (x��Zf��Qfm^��'�݋E��T0`�`]�r��Q��m-ͽLӻ6V���QkL�@ݳ.Y�b
��N�k��ݭ���ݬH)j����I�r�ح�D)T��f���Y٥��ܻ�4V�6[/0���Q@
�4Y�Ab�pz`�(5�J��Nb,���X^�B^�'$u��i��29h��m]]�kf�-*���В%�CT�ʴ�L���͂���Y����љ4�x���Ѥn���n69ai��"6����+wmkԍe��*�7[8���,��,AvA��7�ߦ-�boY��GO�f�Y�)�ڡ)۰s�ϖ�D#�͌�K��fm��Qյ�C�ݿ��;��"�
t�<�c��E��n82���ࣚ���R�azZ��ӷ�Z7�(��RX"I"8�V�w_z�i*t�0�n�RYY�d{���5��1'R�S�%�)lQd0�ۘ%5���EGA�5�;̚.7x2}fMd���Oc�Cr�`7O*3>��_e,
�%�DA�c
,�sF<z#�*����_^;�-�CiIN��ww#ݛ��
�����|ww�r��󧖝75h���UC$���[7a��)YX+u�ib�;���y&�4k<���v�y��b,X;��QtFۢbk"ɩ&m��H٬hU��B/�:H:��l[���*�1A��0�/�X���I�gj��ȋe\��V���˘U�`?3��saP��A��LY�hޡy��6��9����LrSӘ�ӻ������@�X.����J�-.�8�f��݅�J�E[oI�t��Wv�z�M��՘$Ѕ��:�Cd`�;)��*��+�\��.�Ub��IXl�rV�Hm^�]���X1뫇E^���8�A��gH�\8�h�K#3C	�Xt|(T�2��i��h+��=6 �['MT�����e��0(h s�i	��j�H�h݉%��ZB�cx��I<�e�@�L։�p�ok(��ġ���݄^�F����Y	Р�*��Ff��3e�/4�.=ܓ�꤅�{Fu\�`���ըj�F��B�͕�aRI@�� ���_dӦ����6���P���c�1j��a�"�F��ɨf ,nB����Mkv��V:f�X�-	�*Ǭ�MǬb9�����p�*Y��)���Ї�Z#ѫ�wURj����T�� o�QQб}b���e�N^�\�$\z\��K�+�YvB��K��6�;3bʻ�3U4u�w����s���pe��3�[��F�X�n���7V5�&�����ZX���֞�֎k�b(�C�A���)�?T80��52"E7*�
�j@��S�D^�����"'�L[a�����s44�=z[�{��ja��T��o\Ѹ��A�Y����s0����+�5�����y������ew������NT��ح���U���М̅��7Z�P���jvt>����R�l�!��.)D��Fn��R�G��Ys.]e��nH�&�������v����g:T��Rs�"��ѨY�e\@�Xǘg!ژw}��D�q�Q�G_̽F����.d=���].�8�����{�h������OL�4�Ò򷻱F�k��+[�G"C6�mk-�����)�Rb���
0�}���)�/m��OUu���Z]�;&`��ge)t�-Ȑ.\v�NwJ�Eջ���0�ӵG/�\��;n���xy弚�]@.��&��M���t��N�zn�«K��/�]�v.�k����UUO��'�j�N�����%��Ӻ}�1�톮1ٝ5�G����:��W�uf�3_�y���mm�'5. n����BA��F�0�����������r��u�MS���Hة����/G��)dl�9�<┴��S%*���y8�{wbe�x��vЋ;�\�{��Q�ܫ�ӏ7���@���wB���U��o/��nFy��
�A�lq�&i�2ѽvqծF�F�ۮʹyJ�%�YC���[�ul�4h�G��tD�+��^�k��Ä\��b��{{�W_f�t����aEd��ͦS�/��=%���c���t��nk{-;{A2�kW�ᵑ},f�{�I�}}5�@��ZV���R�:K���7G�?6�ZN���Un�v���z"̄EK8=�WY�#)ɺ�0^�{t�רE�N4���Xq�]	w�Wu���(�8ZI��
L��hޢ�ZC� ���Џ+��E�uJ��ʏ�WeuUѸ�Ӧdp���]�VM�[��yv�֒؀qZ�����<2:9�6���*�Tv>7��׼!�q䇺���y_��v������q�[���D��\&��S�̡ۨ:Aӗ�D�K#K}J�h�lwntm���Ayy�Y�GU��m�B���>���!�f�'[�>����ᖫ7v$���I7���(�z����悽o��ѽ�,"�+���^*������x��+H����ٻ�h�ۏ1P�rL>z"�y҃���A)*�%[}f�s{x�I�h7��v�����N�wu�rK���p{�K��wW-�d{�r�Gd˷pt�s�\^\�}X�N�HKt�q��\5�Ɩ��Z��}\�6r��P�]�Wv�ܝ-�uE�6����$�4�9#�'��ws�"�\�|c�"h���F�P�d�Y�_ɬ�*����'�wsoU5F���E���In���]�[&˼������w+s���r�j�R�����T��o�M�V�_<Js]\�e8����4�j �Yi��W�'W-��_X�ѹ'��פx�}���͞�Zݙx�hX$w"��%O�-<�zY��mIө�"�V�.��N�ά���ts˹;ZIF�K�F�ݝ�ر�rOwuι���I��/���Ϸ�K���$�Kd[���wRޭm��!ƹo%��ؔ��k6�{�]�oy����ə!�n�w���y.wL���}3��$����-��3.���Ŕ��wt�����Ի���%˹n�J6�y.|�݅wIۺ��w0]��$�K���B73�F��k2�`����K���1C"��u�#`٨���2�u 8q�`gZ�^fuH��رRs�mM=8m��6�ڜ%2���Zw�f^G�������ܮ�t���L�}��iZ)>T�^eumܓ�.���S�f�T���y�>ӈ�ƨ��
EB���eܹ��I$m������I%�Z�>ܯ�v��`W���Z�� �[u5�-���]��9�Xfѩ�K����{-󴢤�hfN8K�a���ﲀ����,��eZN����4��D+����w{75�%<�+afܴn��έ}������'^��9�����;]#�	VF�]@C@���ڝ+�R}R�#�u����+p����Ar�J��
L2퉂]��u{Ң�p�{#��Wv��}9e��&��@�r�]�	�#1�*��7���X8N	X��gtһ�j��M�K�S���$9���3z��m�+��
Y�BV��L�Kf��һ��Uٓj�u��:��l�\챦q����z�In���GH�*'�D�`��������$�[��ZZ�Z�����1�drZK]t"�j5���̜��&�vjU��٬�-PvJ;���Z�S�;%���"e��6�{G>&n����	�����|�pWh9
2�U挙�L�T�[M�B ���,�~Qc�^��/��2��h�]��r������w���[�^'�V>䛙}�C��O^�)fJ�6 "��Ĭ\�6=�y,��H����<c��a���\�S��ŗ�����[+6�ڎ׬�mc�g���텈����o]�oz��nc�́wb��:�8����7KY}I]췄����/9���e�qKW�����r���01�x�˅�z���y�d�<�i�h�]�^�5������*N5���^��wA`�fm�oZOC�엹�����;�t���렗v�%��z�{�t�_V<�x��Y�b��M6��cm#��]���w�{��W���=Ɵ]#�i`K"����OE�h�,U�R��
��C;\��Cm�]��Ew67k�Ե�Ym�iws��+����?Y�e�iӪ��ԇ+c�g��Os��k��Xn�_r޻�����6&�L����;rЖ�����z���w`�od���uG�єx Jn�p��wc���7o0ڵ�J۽IL�|4��ߝ�h湕{zTװ���!)e���h��kYea�B����+��H�u�h���_��P+/h4���籫�n�2΍Y���	��uw'	�Y$}���\3��H$n��0;3�_/�`V�?bΓfv�9���Z����p"eMӳ�����j�j�b�ӓ@[�{��N'+ F\�n�;�Z�v��j�_R,�D��h�m���=�<W���>���V��H+U����K��-���yg�t�G�]G/5�=*�q�GO��n�q��J�nNeU2u5���}M*5�Y�{3��4���ykA\hJ|;4�-��J���1	����/��;/�L�}�[[ܖ� ̓�s&�S�2��o-𺘮+Sz4Y}x׉f�*(�S�͊�:�,G�����p,�mw*���'>�y��1�uJ�u[�Ü�L������q�ۺK���Ź�z��}Ҩ��v��y���������w���.仉T,�U�n �A��e\aZ۶�����=7^��ۜT�a��Y]����1]%|�zԨ#Ǣ���b��k˺ټ�I����4�YbӕO�`�Jn�Fq�:�Ԫ7v��ja��S)t�Ļ�j��a�Ż�1��A����r�jAwv�Tvwg~�C�遒B�ph�[33�[#��a]�Z�����t���M�0����)\��A������U����x���^�޴�>.�R��``N�ʏ��wU�m����˅S�_H���w�6��dA��1kQJ�b�2TΨr��K��E\��;e���WQʹQ���cV,SY�-�:Ҿ�e�9X�}o��9�����k#�_�n��^��W@�%6��\��.�ī�L��w�0]���-ZmZ:��`�I6w��[tF�0]���؇=�kv�g[[�P�u	%e�{����ek��H�L�ĵ�u���|�gA^��j�bX���G��o��ɆҤ�6�,45�X7Pj�����bK	0�Bv��֢�:��t��w':�ڛ�}�y�gudp��I9[
�P�w��;���j]yG�G�\q����1�=EV:�l��*���Ӽ.ݕ���/m�$L�}d#yܯ�Nm��bZ�V��pp���6�ձ���`^iꏒQ�ͨ��iθ�(�Ԇ��n�,�[�;t1���ھ٦en����q��ݔa�p6��s������[4�r��*YT�X�R9j������#GW>Z�(.���/�P����$ 5�,���Yұv�8�h����:�q1�3/u%Bk�Ye�	":ZN����D��3-�]MT�r;W��%�̜�v-��[�w�7�NH)Z�(����W�'*룲�-����7z��)���WDz�nd�Qװi�l����P�گV�Ş���{��ʼ�s��[�Ϧ�Xd�w#��̹�������FS��#��[:�Gw"v��o.���+2<AZ.�v��F�{�m_P��J�Y�����X�]�����MS��5d�ڊ�9�*;o�1]L�����	�Ӑj�k��c42:j9ۯV!'K�KD�N�n��hf"�9�S)Ю��.VNw���-�vFЧ��{��Ӳk��m�Q��&�i�uVɖ���!Q��#��L���� n�FqUYs���>�Lp3��Uٳ�xI[5Χg`� !vf�Pg+Rۺpc*4e��rta�ٵRtm쬘���3�8�w_2k-�z�uB��J�M\d� :��Ȧ_<l<�i��������ѽ�Ԕ0��л�}�8��rm���:�m��z�c���Dvq��c�)� �[��<�l�9E[��c�|��T��q雠s�F//;v�M
bvgwh�vl��m��@{��ˆ��d%����X@V�\�-�fQ�-	ǭ+W]��{F
�7�ڻ�1ɗ���6A���̍vIN�>�S�v��4XZӔ�E��w\���N��\�\���k�97`���y�����bKN_L
�oP��45��̆+�ۧ��+U��di�i�ۚA��Ñ|1�w��w�d�/ԍW�̎I�N��-��їڂɓ��Ҏ�ʀ>:ʧ�b�G;�Š���&�8e�)q�!�2>��9/p+�{�~�D����&v��t�&����[9i\��#7�v!N��vydܽ�
]�ff�-x���t3��Q�E�t�F�y8v��WO�uF+��p�p�U�^f���^n�*9�v�Nw9�:S��6��SV��4ZT���3j9���(h�agW5F�Wg���P+:k��B����]O�����5Һ���,���8N�SU�V���;�}y�*,�0�a�I����Vz���K����z(���Ig#jE��E�[��3nX��1S٤eJ@��J�[�E��og�IvA,�Sogu����s���dE<C�}z�5��nM�;�g[s��U&��������,ɸ��XP� �����'9y��)t:���[�n��	�	ac���})��*]���],sz��G�e����`X6���l��Q���y�^)�ѭ��Ư3nֈ
������sI�[�=��>�N�.�ێ�48=U`�td�׮bj��J�nQ�r�G��,�[�z;dr�V�Y.����-���wp���[{�=�+,e��'b܁��P��������w��U���R/�����
 /�C.�����9� ^^�'oU�=�Ի�$y�ֹ]�M.��tV�fm;Tm� �Q�ˌ��UWN���2���\YU՛w��b��>���C���,��]��|�W\;1"Y�I�ձ�+Lͺӂ���v�Vx����闸�`$��K�LN�w,����-����"�eԲ�Z�N[�
�q�4�6��tz�m�Vry]�c��`�ok�G+Z���`鶰�u:�N���:bKz��L�d�8�t�;xv䵽�0�Z��RR�v�,�e�=b�^��+�w�8��(c�I����3C�^�\�*��,i�&�)�PZ��.�^l�(��6�=x�"�U������07)d�K)Uʴ�׀�����fs��Pg,�ih�͚�gCE
8�\5.t�1����&�%�r����!*���m��m�஻����r���ո�v�vv�M��U�����ˌn��]>b��o4i �꥙LQս���>1e�}yKAٔ�.p�d�j+Vv�9�qu|u��N�p+��[/��rvo]���@[��{�GY�\'`��'�u�%KɊ���O�=|qu����)Z���JH �����v��#m�g�t�W�p���'���*�dus��B$(��2�fE�{_^'{U�sb�z<�R�|��86�L���Q��T(]�0M��|rͬ6;���^<�sz�/�\�'@p�����>��cs/6s'+P{���W_e�k���ñk���wZ*
�J��wf��u��Ãl���2d�v��q)9�cqݝ�Ԫ=���4I��0q��V:=6�1R�o�*T��X�٧Y�X�)���^f������򵶫6�ɫ�lS��
�[ΪU6�C�;���P�6=�c�/��.���N�����"��Pзs�+ҹ���[זօ�7hV�����x/(N�;�E�.펪�^�;�ښ`��������P��;+*C.��e��<�E�|{��qԫ*:W��os%�+r�(������9#�)`��ƇYM�:��n�l��w��8��=:�]�z��١1��M�5��"���^�ȏO��*D�{�a�jЊ�;��M7r����~�ɒ�ܴ�͹a]`�y���/T��\R���0���v2��<' ��u9�1 +:T�#����CJ=U&5�|������u�i���nt=���+���w���*�/D��\zp���ڎ����8Jɂ�a�p�(���Y�b�J���PA�M!�U�b�wr�t���j�,f��j�K���x�`��;�,Vգ�K���s�m��40B�@�w��]]��cښ�2��v��Y\F�z<4Z�z����$���9�r�	ggSe)�ӦgK��Ǽ֫���,�2�[j�p��ggc�vu����\���K��c��e�Ԧ��s�6:��{��������sp�)�,B�q�Y�U"�	I���X��!�[��X74P�(��ھu�
�M��8F�����n^��ٵ%Ͷh��,r\�	�J�rU�hjj�+6\^�Q��ئ"1ɕ>�+�ox�u�އm��Z8bZ�]n����fӢ�h��ט�0�O�Vj=�9���f�\����(=N�5�WC����8XOE��S[�!"4.��V��в�\��`
 ���/���

�G$PAW<|��\��đ~�Ry�U�X���AO$͈Ź�VEXq:�՚B�[�m-���n!	�s�٭��P�x]7�1�8VXda�K��%�v�����iL����ׄ\�:ҶJr=��:)g#��A��p����Mt�a�7���e^���%	K{�](�Y�Q��M�ܗ[�Z*��+_U��H)Cx��}|h.gf
�DǇ_���P��q�!��Zft�y���M��1csu�V�&:��Q�Kv�pe:}3�M-C���p�y�c�����\:y��~z��s	=CnQZ�Gk�Oe,!���J��-�WP (��4��*���3�����)�1�%u��r�1Ǘ�6L��F�8�q���ױ��ۛm)H����9�wO�oK:YsXpPt�7�ip?q���Ư��v��T�\1��7Ա��|/w�WVC��wyo�3�4v+�}i�J妻8ޙy1Yn�%�4��]ZKi�4ѭ	w�J�C!���n�}2��ܫLdU�7�ܹ���Wpܚ��].\(�e�d"�j�	e̹xt��zؽ�]\���j����!o6���������[���o��<�_d��!�5P�yL�9�F7��F�[�!:��)X|���j�6�p2v�u�M��U�&9�5Gt,mɄR,ɖֻq�#.tU�^�Vu�ɭm�+*J͗�j�G6\y-,;�q��e�%K���e�J���M��n�ˬ����w�
��Ā@�M����X��
��+���.KG��Vfv��6/�����agGJ���-�k�hR.��7����{nNֻ�9�=��T3	�ᓫX̣�1m����dl�%�m��:�|%���y��zi@���e2��2|�����������7O)}����5����G�J����_pL�ii��c��#�Ԯ��ul��[�u���G?{���+ؑã˳�U�(�� �7WU��^�� 6w
��hE����ܤ�� ���G�~����gcZ����
i�Mz�0�wL���R��H'	E;�r�"	�={Y�|�Ed�"B����G�},ur���^��]ڜ_�:��'iV��/pRa�J^��&���8{�ūVB��\MYK!��z�#ѯ!��w�c�y���>^�
��1��!�O.�T���V��Vh�wE�{QCV��#ՙ9��whp&n��.�߷9Y��u��u�m�c]�Nq�Q��R��I��[�W՝-2EMN��]�xC����˺���=���v�7%�M�w{�p�:�H��_�$��=��{N ��9��3��[�H�pa�y!��K�
��!���:8N%1��֮�;A�g� 79m��I������9�Ռ1*M��3{����+z"��Ə�mC��B��v<�}�/ �[�'�~R ��RHDC��w�7����҄�Q�>��KT��G�>F!7�Y�AfQ^T��t��W%Gy��wS�mK�|��}���Ӹ������Vd�"�C�v���s_�m�}���ˤ��7%�1�2;pf�8d��E����H�UTEcH#PFDDPQTE�X�#�E��U���YcDH,��`��E�PDI���Ѷ2C�}�:��z�l�H�#�/aE,�����,���ry}�(U
�L����S�`�|��k[y�i�p�-�J��j��͍s�ß;+���u:��r����[֮��u��<��s���zb��1��֗�����gB����1�se����mN�*둞��r������[�TAɊ�=������%��cL��  o��%>Ƥ8;��V��=J/"MNfJW������~��%H��y��Uh6"�.��x}� G��_����g%w.4y�SGy�����V{}5�@���zü^���f�z[��-��9ϐ�UW��C�j��x\T���ኪ���3�#�ec�7 �贺���U�u૪N�������$�`���~�OQUv�)��+Nu�a��?E��Xf�Y/��-�
�7�Ky}$!>;�!U+mF��$�dQR(�*�VB�Tm�	lj��R
6�R�)X�]�� l�g����:���d���B�O'Zʜ�@��{Q6/�����Һ��m` v���\^)bE\F0�b]�./Y�%%�(��+�j����mw�9V���VSG*'�V��+��i(*�u�o��}_W�L������M,q@����L�p̭��R��R�jޛ��v�j��8��<0��ƛ_|+}��|>��Lu�Wk��E���Ӝ�W���R=��bج7Y]�/��%u�/�����U��8��*5ec���y����}ջ���CUg:e���n�)��n��4��vH�����odg��̋��#����DcX1"���0�`	(1@F �I!�
1�,Uot��3Ýﹿ��Lײ�л�<�^�m"����{�ч��ʗ�c
���nwu����Z����|>(7���v+�B�q�h���i����˱��*ج����Kslܜ�X������3��kuueJ�Zz��3ZG���ǯ��Y��k\W7*����WH��\����ݾ׫up�nx/s�@��>��'�(��̏� > �7���rD�z������{O"�k7������)�}ΰ���E��i�ʋغ��D�.�=׺� ��sY-@�.�K:�ٖ_���IN�=w���?Ut�=~�3��leK��8�ɟ@N"#��R��:�nz�,�|����7:]ԉ|:�^���&�/gEh����K%JT;;�8Q]�< |*�\�?��z�]�8�T�ht\����G�����0�m׶U������,s��uVI�Y� |8W����>������|>:�w^l��S�B�t��Hfv�""�Ϋ����1����������w�'v�;/m�!��):�q'-,U�[1�&��WxX]P	W�m�*�q^M����s��u�[��z���}RNX�gt��J�_W~����`I����yjr����t��p�M��\g8Y) �&Sx.����G�}U�*=!��]e��V	�r� |
��XH#ߠ�s���}��|�W�V���bu9���jY�f�ڽ�]���O_]����L1o��<.J��#��P���O0c錭�9iev~v�u�-�������s���S���}���ƻ����o�$桝�������b#�#$a��ȫ��F`Ŋ!I��P }��yH��{����|y$!XOt��T��4��zg��͚�N��4�볩��m��4;}-P����Cղ��F8�����ҳ�7MM(�7ծ��l�R��G��'�2l�p#�|�{�����	!k��M,�CmAAVQRI`�F(��2"�0��@�Vj�U`��F,B��X�*�"�
��ZfQF1cj0�}�h����},������bY�r��	�_i��`�p��ϭ�+�z���ʵ��Xvح��a�{'&�ٱ>t9�Q�ǐ��f�D=�8�l�������;���V���ξ���ê����������|[�����+={Tb�fR�rt ��t�nsBt�6�5�Oo"E���.�q(�HOF�z=�^�x��k�(?z|1�y͚�%0��f����u)׾��i�WY�]B2�[���dj]
�Zӱ����T����z�s;ԡ�z�Tk����f8�4(-���꣹�p�M��/��~�`��nKڋ�rWH�l{�脤���Dz�zz��s�8�8)��Q;1T�Ot\m���81GnY�pmT���v��2z=���bOe�)���3����P핖�� �"���(����ba�,bF$dEPE��AY%imEE��J�\!X�������m�>3.���W)OR��ץF�C�0v�c9aC�.-t�r��S��i�GlͲ��×׸[���5\�6,�[Є�.��&wb�0�b| ��;�9^�V�7���DD%���n�xSe���q�$�u7V��LT���c��*W�4z�2C~�ڬ��6�s��|}���9�4�S������t��W�J�����m	���F<�5�!�Ũ�����"1`��(FEA��d@Qa$X�(*���<�@�����>�><nJ����w��}���WVw�ө�ڵ6�ZWf��u&�p����I�슗�G�!��k�ʲ0����]drղ�(���Qގ�4[Cr^���u�c��o0���^Us̬U���>ȵ���(�V->��v�x��T������g}��q�W����$F,���V(�� )�Ag�C�@�Xˑ}���r¼��˧)�ԍ��/i����V*f��uͨ�1�W%��Sb���ߍr*�Q9S�0υ�\Z�&�H/n�j:����.���� >��}�n{�a�QЂeo4�e+�ص���qU���4m�jk����rw9�v5��s�U��  �8P��}�Lt���8`���d`�2�!�®Z�SC���#���:���Y#�Q�ػn5f�p���S�{"ݬeR���ħ��9��U0v̸�����#�Vvk.�|�.����O.��wV����x�d�8��g�$��]���І����Q�x+&� �+xouUCEa�k�j��sjW��\�[�[�����Am��=������=2GmMD[�Z�m	��ywG����{n_L�M{R �p�������U_z��k�0U�bU��i*�,UEb�(�"���PX�Y# "�QPE���J�FET*�DVJ�(���"E�2*#-%B�T�\�{����_<����Ѿ�t����ɽ|��}G�_M�kw@5;�	x�no$L9�К7M塷����ܔr_�n*�Wq�wM��{Ѿ�1U ya�7�']{��N�K̅���Z��4vk3`�P���*�`�
Ү�����4ڕ(��9�3Z}p�d<ã���'m�<4�X�ۙ���Dd��e�ڬ��${�����E��"T��# A��D� �@�0+� �$��ʺ��	<�{e��Fga��eӽu�]5���4=y�~��o�7��z��Q�gD�����h&6���/���r�vSDڥP���ұ����W�������ۃhc��!�G�� �}��y�#������S�4�r�%�Ù9L��թy����w�˧�<�˴��e�,=��[h��O��{Ր��#��9��5\V\K ����U��Q�j�r懹��x��Kc/XD;V��.�%�f��!�
�ה!�~��������Ġs�R��v7�4m��p�p�
�{��j�0�Xi�����*҂0Z�V{�ư��&&����w��-%��t�kN�PQuh7Xb�'��2���(�حm՘��
��FaE<�aɤ.�UM�l0bcQ�������d5��ѭ�jӸ[ӛ��2��C�&3���meue*���x�[���:.�zw�n{��x�L@[吣2�XKVS��r�љ���Y��]��#%o�r"�[�%��*VH�Ȧ�1,��Ab)�X�#N�ÉU�rRi�J�.kn�6nBh�����n��%�e����uk1�M���y�x;�3I���̸ �GvhӬC���o|�Zٍp,��o�.6��pנ���: �P ���Tr�e�	g�C#�J�0֍feP�n�dr�K�k���n�뉐����;s]�Ň_��T���d�M8,ݲ��W�U�<9�eF����$J�v�(���P#kZ�D��b�Z
� �0��Χ�Z�ә�J���p��yfL��������wPLc�:�q�:�2*��m"����Z*�|��;�\�]f��@�Vk����i��X�7�z����N���*����1g;Ժ�̡Wm�s�2��s���Q����y�ەnh��M�5N�|�U^Я�3d�vl�8=λer;d��P�e�W�zo/^ކ�����I��NڳwL�b̵�wU����{&ԗBÝ��m����Ņ���a#�ٝgz��L�0�.��%uH	��W��`��mˬɪ��ϳ0���kw�y�F��v�L�}&Z&Ico%���TVGJ5��P�]���#�[0��}lU��ز���MM�0f�ҏ���(�Cx�j�^v��6a�x�k�:,�����P�������׵z��V�ɳ�(����@��C��v�V)�u�� {�rL���Wg4۴�w=��58�|�S	�n�S�����W��z�T���Ƕ=x޾�$���]���`5;l�ƹږn<���핈�t�ї�521��9og)����1d��><��Ň�:���ɹ�^�&��K�gz��zĘ+���ܼ$�KZg�Щ藴�;�K���χU̗)��j�X�j�N,N����A��y�Ǘ��Wρ�V,��w�}��Sܦ�#"(;�vt�Y=|ڽ�"9�����4�zmjT��xC�ڗ�r=�xz`<�^�s;�a��L�V{�1�K=���v��gD��;��g.�o)�a
�B�K��/[�\���h��G�9@��ծ����ޣ�zfoew���\_�7Fإ�0��ט�g�G�'V=��9	�{9�$�+_ވ�����w���n���EI#��p&� -1�x��NP�$:z�gavL��W�������΂��W=�M泿O�$�H���!����g���?~7�,�r�����f���hU�\���j�^M��rp�s���?���b����yw�l�����	{��]l�X^��6_�{����V�d����9�wꁐߛvO�#�%���7"o��|"�(7�I��LH�(N��>�z={돕��<���;���z�z���we�7�h�  ��B��!�}Up>�M.��8ܕ�ػ��6%5?Q��g�PO���@��|�|3.w�L�wy� �t�zs%�ه�
 �z�!`��7n��|�<j�z���	�¼	v�U$������V{�L�:�\YNM�²�'&�nf�&��Or��v�ݵ�IYW���v�4uh'
�.F�GQXIIn�xT���_����������˱s�fO�ǣ;%=��&�A���fV��_���->�j�>i<�wn�����.��x����`�|G��
!"�	#$XEX ��0�đ" ��A � ��jOʱZ��v���Yݿ�Ae���u�t�6�.���/�ft�b����U&3d	w�c��»o���܇�rb�v�������Ӓy��Y��'.�_�
i�<�c����c���[�����=!��|��/�R�G�k�A��x���I�~{\��@~��?�m��� �D��F��XV(ª���!RR0-�Q�R�#X�@�մm-�h=������̏����ЊXG}P�e)��B�V�4���8�	�*Z�a1u�T[�kU�4Z�A��YD}	w�~��Ϸ�W"��(�Sr؎xz��. FvD��ݯ���Q|��Z�V�+�B2�!G��e���,�5�E!��> �^���<��w�5c ե��2)%�*QE� �$ @���Kj���GP����9	��XQanѤ�ox$!%�)T��S��:R�M�!���ua��3"5:����S�u����5%���	Dg@BQ��13\5�C@���d[(�ƶj'(���-�wm��F�@�Piw#߳�����.��OВu��[�}�um�S���twh����~{%X�P�ڑ�h������b��kr�ܻ����Y�}%��2�Ћu�`N�&r=�}�E�0Q��"����TT�(�db,V1Y#d# �(��UE`�DF*1A`��	H��Q5J
'�������w���VEry`PU�U9��l�C����Zg�t"��%�&��=�S�t"��"�p�����s�f�p��=�g��|>k��������Yn����rލ��>��n�N�T�����>�Nn���M���SX!��~�wv���z�^�ts���bc�?G�����Nc��?!_;�Cd�cB�&�suv�
�nq�]�Qp��S�{-�</�M��%���4�:+{t��Xq����w��G�_r)�sO>��M�z>�W��=�}�����.>,c[�Um�������,Ǎ:�鵹�n�L#j��E�T�[���2����o&�u?��3�� ��ܾۏ���]��TN��S�c'(����6>c�n۔x�Z��ծB�@J�w>lt�JS
<�dU�X�"��aH���"����QD�3�����ۺi����}<�-:�\9��q���j������7�T����r����&*J�0" �2�}���F}O�+s�ǧ[���]��4g.О,��qs�I��vYA��͑��<��Wz�ȝGҪ)�l^+��Gd��2:��� ���?G���G'+�e��۷�o s�='��Z����1'�I}�p'&�d�!�����h�%�כj���JУ�S���Jb'%�r�A�=��G�#g���.����.:��{Y[���D�����@Ѫ��$������U�9�m�{ny���V�sO���T�!&2�>�{��`�|_㿠b���x����`¡��/D�*g2�ݑ��k��*�.>�e�=:�gǥ�r�X���f�@�9�e�B.�����x(�n���ے��v��g���u��1��7����`$X��y?�z���.��Gs�,N�w���o:]�4}�z{�Q�}�:�uy���Y$��-��|�W�ipG|"�{�c3��ܨ�]� 4:IRcm,�`F�!NBݺ�%����ı�"2c��yk]н��{F#���3���}+�� ud�������}ċ�
s��sO<�Ϫm���2�+:@#����pfn�w��|&%W.��w�x e��t���R�����{׽�N����}����|We�FmN#�Cc�w��G���#���|�U׶	�3�]�I���q�J�m�L�h���G����g�3?#Qf�-���§3�j�]G��0č�,���&���«g���"�Gl �^�z���8��YBEW\jy�c�		�a����6~�B ��yě�*D���̑u;.oY�YA���&.�Vd[���΅�����Y$�Hy��~V2,d�ȑ�P"2E�E�
E���9�{������؊""
�������T�hTE|G���k����'uu�|��ﻸ噽�x-%_q pv��l���	u��]t�!�j�¶�.����eo.�F�7ܟU�e�P�a[�7�|���A�w�1��^�,�yxܧZ0g0�McF-iW�C���e����Y����?��}s��[^��f����ܿ5��zǞ����jtW�m��s&��8A�2�GY����gVTOv�:�!lY�U�ѻEm�����菎Ͼ������dP�r�=�s�=s9ٮ�a)�zO�Ӂe��2����h�Cn�=\�1Av�=}��â���}������+S��ޠg��s�1���
�������?!�}b�ƃ�c�3Z���1m�q��|>���w;�;-o��V1O������$H�?s�Q��ߊ�S߿J"�X����q?�WZ�-��s�UN�C���}��2�!	��)��)َ�%9��]�����jb��_����	��]űoG�~�5�J9�h{����^8� I ��(��*��"��P{J�"�Y`0V1F" � (�RAAd�$`
*X+��c"�A�X"�1U�* G�ϵ���ޜ2�OXk j�;��2h�4�}1ڛ���k��'e�ۙ��Y��"�^�����TЏ�/��;L���X��nW�rtdw��?%�d}p}{!K��3�O�5p5�zqUf<%F���Aʛ��g��ޏz	����ۛ𙟣h�D��1��r�*�TL�}:�:o��Ü��L���˻�TQ�/e�#$�z=7�	G�q�z�[�ә�اÈ�\[F,�D�\%oQah�}�|�]��u�3?I=��x��|�6!�1�����e�kn�� �;Q��?��r�3N�����Qo���m�}���,�[�x��fb���<o�V�AS�����64�����N�bE��9�jrc�����Ɗ�~�>*��{[
�ِ�)ia���}��+��
�ۡ�k_M�yZ}-^�<��&{D��`Ω	x9���y�����,T�(�H� (H� ***�f��>���O�_V�faO��z=N�)Ɍp����N��gDܞ�c�<��v��s;��>���6�,!`�dT��~��x>}ϻ���l�@�ݻ���	ԯ4�oS�Ǎ���{o�7k�E�v���rG5������\�����c�+�Fe+��ޒxG����6���pd�<�z�����קO���'���b'Ԭ�A8Y7'C���?u{�(����KnA��)��z�*�<r^N���� שn𞚶_Jv���� 9|�w߿s���?�s���U�0�WĔ&�2�Y^���̠�-6M�Om�h�����>�`#���f8S�95C�C��N.�m�6=�,i�_��u�t}	>���l���$��G��jF��l����݇W9tc��g�~Z}������2"
I�G�	QP{/��?����O���1��"����c<�"6j�`D�✌֣Fm��d��k�ʁf7oz��<�K�~՟#���m��~���? 8UJV�ߵ��oqp�ͣN h�w�#u*��1[���|{FN��5�����PJB��|KݎY�:���Gy��_cГ�#Q��DB,R$"1$PB  0 �*�F(
#PATVEQb��b��:�����'D-,�m�Y
��"H�� �AAB) � ���������J�/���_f�u� �y�^M�0K��9W"������y,rY]�&v��nr�n�]Ѳ�V�L�
ѽݛw2�t��NL�޵�$&�j�R��7-�>�;�܉b���GF���^���ܴ�v���W̡;�:��v�	�ވ��B�f�6]������GHT�u�o�#�̥���EV����1�I����81X�V����x)��Q��e�[�����?y���~�ey������,I�������=R�˩���P%Uy�hT�t7S���3B*��ΐނ=М��R�}�D�Ó�����#dj�����:����N9���Fĩ+L�OF�:�I8�a�G�$�3�k�؍v�;�l�X����	"*H�20� �� �P���ϗ
��xjva&sk�6T��&��/(�����~buګ�	As��*�O<J뭡�יV������dU�7�Ѽ>��B����H߾9=�:�g����>��|��]>7aQZ���*�Q�UmR�XZZZ!͋��T�r��5N:��&C����x(�;\sC��ٝ��c��w!�}���L�ri"�r_T�]�֯'5�\�����ʷ<ӳ��7�sW�����eҳ���8��A ������QտDz#��ə�7uH���.�l�!MY1ۂOM�*�pY�^���I	�!��ENX���FB5!l�0� �$�
���=荭��0�`��$���C��єX��^�+b,#�k��ޚZ^��ް�����noU��С��Y���n�Ϻj\�}���q��Vf�Ʒ�%�ʻhS��=t\�,���F^|^�Mt�Q/��ͪ�޵*j"rx��6��T^
���]�~� |I �3p�z����V�O���/$`�v�uq�H�EdO����iO�~0Ｘ��#���Vke����;T�����dU��T� �@R
"�$U�RȌZ���#a �'��:b!y�����_5~�Ss��?x��&��||��ֲٗ��@tǅV�<�0<==����, G�yx�Zs����%���rK���wD�m�o����T����7���m�x��T�rZ�5	,>i3BJo=}��xh�s;]z��І��.�
E�k�+�p۫[�ַ���s0ְ����C�lͅж^\���M',� ���f���£�e�WMB�+GZ;K�:�˾v�mv���k�R�
[���5Mas��{��Ni:��)7���|Q����m�J�"M$h�A��K`H��7����2�e[m�LıR�j�[uwnh��6��,E���7� �&��T���J��gv��3}/L��G�X#7ܙZ�7�a�;u��.�9��м�4)�X����hAH��H��\�/%Z[S�s�lMs!��hf:O.^[��%��Q�I���;�'C	�I�M6MA�;`ƓD�j�
�s]�m�8!��Mi��u�.ir��:neyAT��%�WuD+oP�q�i�����U���j�t[�Vk�˦@��k��(�$;����t$�A*#X���Mq){g.NԪ/�]��i<ƹ�����U7)mV��۬ˉ�zc[0��ߊ���P%p��4��`b�i>�vZRKU�Jަ�]���z�.<�6a�,�b��S�U�(�U�Iٵ��̪���������Q)����ꉽ��v�*�8^�Mޗ9��x�&$�"���f�:'`y%�?��${Vp��Wlzk�͇dG���H����%�U�����=A[����؞�hf���9��-u�=��}�Υ�i�����R��k텾�}�x��r�mh��
���O�m�odM�L�]�z��a��{q��+���a�t&�G�G�U7+�*��L3�յ/2�4�Vv��4��Te������:.!�:�_o,��T����]dkH�]�v�Gw`F�q�6��l����IB�U�9�8��V��֎�|d�֝�BU.Ei���mL�6��YZ�|{��v+�:���b>��C/K~"�r���ۗ��^L��mr�&�O�G^8�,L�+��ə�f��!5��d\�Go
��kV�u<�d�]��VV���Ъ�tnv���p�
�����ѻD���9�G(-�&��r�U�Y��Mpy:�r�W�]c�Lu�z���\�lᔐ����C\�6z�	�b[Rp�\�r(hC�-<�7G�-:�Wq�-�t$��޶*�ܭ���a5o����٫6,gA��oLq���3�Xž�ܫ[J�;u���$��7�k�̪����epɢJ��y'Z�����vM�L�u��[�[	��N#�F�d
5������cB�k��NiLl��EӺ�Y;���G��C�T���yˤӽ~	'��r�a��]�t� ��X��+��R>���g��`�����r�g���׷3�H�������p������&Uo��*�O�x�����9�hCZ����7z߅��.� "�vA$E�~>��a���5f�N�)��uL�]m��I�ũߡv��Ю��c~�4l���!�C�un�b9����~���"$A�"
Ȱ��	$D��U�`�?y�e�9�����KTk��o%R�JC��^�!D��wy�ryD�1ͺl`��B��b*�U�wy��֫� �k�����|�o�NK�Ovʺ�TL7F.�Uʉ�a,<��)�aM��|2_Qcy�\W���?c�>,U�1w�8�w�,���}��y���/�{��*��J�V0�B*���P-��e������;����T��l;���O��,��NQ����f�Q�e�H-��McW@,ob�m�9L����7�c-���ԉ>8A����{�ex���aB���3_��y��ڝg�!gA�P�G�,�~yF�_}ㄹX�oe���	m��PINk��ʀ�FJ.���a£|'�3��OZ�Ʀ^ 	�9}���=��seq�Y0�(~�+>=�yg`;��G��dC;�ˆ]v?X�`z|�Li�e�����+y����>�?W�ݝ�H���Ҽ���f���F�����	��?����XG��6|-i���o�}�짱��	Lلx�F�*�}���Y錇�@���[.+���h�}��>����:~%dr��$�s���ߩQ����xv�'f�g��f�}]�E�g�Z��taα��^D����z�<E>*'q�٦��J�F�[�W���>�ޠA7W�??�=.-�R�җ��B_j�.e��_/�/b�.�pE��������H�(gWUS�a�u��kX����s�4k 1��({�x��b�������Y1���y�d���b��b���b�KW�(�v��?�j���<����]��:&c�w�@t�'Ւ$�y�3�A���о�0>|��4 u)1\&:���+�je�ˏ��V}ۑ���ysܮ^�v	P�͌���	ђ��J�=�*�aŬ[}��44��M�uxn�Ti��/�S@�ߜo��F*��EPX �!"g����Ƿۼ���'y%C@R-\9�p2�� ��# iiw��|rO��H܌���z!~:���tZg��)�x~�?E��
K�F�����nO����tb/n
�>�Y��<��p�֌����I�2z�f�\���ftOYZ��&D�Y���E�=�G��͗Gx�����N9�I�]^a��;@d�0�I�hԍ�[<��Ú��K�w�PdQX��B"�AI)QU=����{��~y�uX*�_"�RܢwLW�Ň���z�V�gv�������b�b�FìR�r5S����o�3!��� =�u�nQ���p~��Y�¥���� f���b�M}��9�����}{Q��c������]�&M	�tC�,��s����~�4�� ��fd���T����u�|�~[��վ�`C���}Y���WLR����U�r9'nYF��{ٮ�{�5��$��Ǆ�F�ܔ���s���D�D` ��D��N^DC��h#��J������Y��4ߎ�A:9��0D��+��.����Yj�<ZH++z�����>�o�������4��
���\JC�V�����e�z{A9]ٷ�Û����t-+���p����m�|	�����8�X�O�YJn��z�p�e_LC�ص��_Gy�c9z1�
�j�#�׽3�M=ˇH�f�%�1�j��q}�_~?j��P(ʵ� �%HVB�!Y-�S�;��~��뿿k�UaU���}�D�Ͻ��Ɇ��\j���_�=�8#�݈�a��u�{C�����z�x���ά^�C�ה;���Ff�E���-U�����..ޚb56/x�"��C�m{�Ƴ<���e�b�ePƕP���wۂhR%���W�Gm��G�ܯ-�[��c05!)��=�&�cS�3"���r��q��g�5��vnN�4��W�����e��USĵuވ�E���#��`��DdX,��U�"����2 �\Ҝ��2�x��	Y��ϙH�3OVĀ<1��
TX����� k�%�2�3V�6��ǒ�,��-����|��]�O�_��qL@�����5�V�j�7�U��2�O�e�s[md�p�Mu�^X𫨵7�Ŝu�՞�G��/�|��d�Nx	
���М,ۇٞ0jdOrn흄�����!����h�a��T289zv��,�<?n�rǶ�v�������b��+�p�z~�2�&�\ ��9tO�0����od�#���H�*��I���(V(��4E|G�����7��z+#kS�9�Nn.��Wp����+;����5Pu�����?�L�����W���ss�,K�N�o�3���vͥ?�A:z3�с��(Phǜ:��E�#@������� ��5��_��z�ﴣ�����G1�8-ʉ�.ʚ|9��~�13�l�S�4'�;�&(B�s��`��΃r��v9�����e�c��;��CX���Ҿb���Gz�WDHeʱM��n*7;�( �8׶�6ë�s��^i����D��Ƌ��G'�{ѽ���ײ�P��z��
=��֧���'�����*9��a�`��SvL�^�B:6��0C�yr�{ S���Sf��p�W�p�sq�u�Dx(�0>ҮG�7U�����9I�U�p07�K��6��370�^Y#t@2�)�Z9�S=���U�1��2�'�76��u+�T���ɩf��"]�՜2�v6����Y[Q��C��c+��.rjɇ��Z�xk��_���2EP�`d�������~��:�ԧٞ�k5���>����]�&��so�ϔ��G8��lxzӊ�ެ�zi�]vE��ryvN�=��,qYZ�	�1�V�v��~�pq:���Gq�o̩3�սq��1�d�h���G.�i��0�T���	2=:�k8f΍��������޽�Y�й�/�	�~? � �a,�H�#�{�������>޳�5��8�ZQ*hcv�6���|Do3?9d_<�>н�#�^�6�R��*���yU4JE�ٷ�{la��0�g���g�3��8�;¥�#Fp��e@������x������b�^s0�8;�7�d3`�~�DS��ѓ4���>6�ѳ��S8ƫU(x��+fN�3ʯ=ނ-|Vv4�c+�j��wnv{8Q�b+ C`N���r��sQ+��{��ì}������O��Ңl�s��7�'��Et�Ɖ�3�&���h��X�g�u�-�㄀eh���jn����O�(}�Y���W���
�[P�b1@F*�H
AHb�R,+$�B(����р�Ȩ "�"$EE"��������{����<��|���gx[�P�Rܝ>j��N�EYHW��ѕV��uP���7�c��&�8�5��&2��bޕ��@�}��; Ч�k5��v\���4��%ԅ	��I��n�k���퓴W	�mb��#=>����j�D���$Apk�ރ]�\����Bc�)�V!V��[Gw�xX|�oω�T�^�=wM%ǟ�+J�Z2/NI��>����,�Ś�!}ƨ��i�@`���"3F�A���^�3�8M0���!�$�d�
*b̗�;Q��.n�C����ބ�~D�Xټ��>/�;#�B��=�+Z�1�r� �T:e"���e�����X�H�ע2�q�̖��G��l/�X0��>?���{��B�] �Og���Cd��r�E�jd�gf�ӕУ&b�;�,<��|��>�,k�7אf�5���W{�X� ���d�R�%����}���#�1S\;�)��1��J��B�����oO޽��u�g,�}��e,Ÿ,�m`-�u�]�Eb4D�s��έ�:�.���[U%�8�U�&�4�������c����n���G��ɥ������?�5)l��$��bs�9�;S�y����hsd����>xKPZ)'}"O-�T5j��7�����&|�l����O i�.a�Aw���2~��D޿��'QɅO}p&s �ۺzN�R��D�`�ɰ�d�8xV��ve>D�6c��2��N�������w������폿��|���� N'7�;�z��%-纽�	NI2�AG��1���:̞X\�n$�V[����ɳ�2z:���!+�t~��7_ [���S_ve%b�ai�)�h�.�ܸb.z\N��`�+_��,c�Ώ� �����ͼZ�\�m_��[���o��G�
�/�s�w��B�۰����oy��f��x�o�L-�0u��:qjmCG^1�ɒ����)�0��Υr�������3�1hWi��x�?�Z)u���ۡM��YӐ���.ނ���.v>��h�n�K�^�~��
���	��+U��G��?v����cb��{;��ޔ�z���)9��E�U�;���!d�f��ӧ�9�����T�j4��-�w�G�=��" �j.����q�3RxL�@}N&�YȘ�^T0�������9��%q@
����
yQRF6�j�<�e�ƛ��az�[p���.��?)q
�3��[��6OG3#�a�x��SO$쎱bY�z��P?u�:L
�M�Zu��W��ѫ�P�����L��oK���x�5�{KE�CR9��*�e���1HG������;ʢ��"��Z�]=�`xH3���������d��qٶ�,���>�-�f���%�6D�.Z��jN��c�����Qhݸ31*t�+^v����8�ʄn����  )$Q`H,��;��o������.π���[���AH~�_"���!$�����y[��,�Z�*ɲn�E�:4eK�]@<�G�>"�ݦej��X��nA�m�G��+�
�������nmoۃz��Yq2],cq#,#M�x��U��4Dqڂ��� ��KV�u�C\��nb-����r����� ���b�ۧ"~'�EH�9���k�%�'N�܆;(<yGi��f8�a�t%���w��.X*�eP+���9�:3L��}����BЯY�-�3l��{��0w������X�,���p0SE4#M���8�t�����������5��ֵ�Y���GY�X#2���37M����Y7q2c�ʺ`�딦<O5�.��y߆��V�Di ��"|�e=B�W�ķb|�o�P�|�o@�j��4aCv�
:M�eɭ���$Q�<繷z �ٰ�Ö��6�1.%�G�T�u�野��4E8���y��aԩ��%��� �(��kdE��@�tI�F���q���s��DRޠ$�h��]|���4@t7�`�w*����k�y�
3������;�i�w	�ų��w4p���Q�=��Q��SF�f1��Y"VK�X	0U	�8�䩺CO>��24��dc+X�q&(��6�$�0����~"�X2���(�[�E>�n�^z_��)���/��T5X(G�u�A�9J˝	q�=x���S�}
��|!�؃��Vw%����m��jd��fw^�pj��..��S1��2��Z���K��bܾ�a����n����C��}������YV�n�m���^���v�.ϲN�@:.}�N\�\ݑ���O��e������Σ��d�__ũ�RfT�w����Ƚ�F�UrҴsb��˪ڤ���T�X[��"�
G\�l��o��(V��]�9��d茙ب��󶝱��O1wPY;�0�=*�Q�C�ڷqLi
�r�V���Ұs�%�v}���ur�����i��nR֒�8�j����[�c�5Y�N�3[�;�K�vv%_,�զY�ǒ��/�v�j�������"��p<b����us0�f��ؔ�<���f��eM����8^�1��R��x��Q=�I�p��}��j��_bۙsv8����]�����|� �Z��]Y$��[%fh����X�Vۙ�x�]ǻط�]������훵�\z�c�v�8���6m�7��j��iRh�U(�B�ڇm3��=ו�A*�����IT0۾����� ����B���/i���Ȗk�u����%3�J KL���Pb�l�U���5T��?����8mr@fB�p���U��xQ���HL����xX�:���<X���y�%h�[������WEM��P9����Y٫mްE|M��$��%�(���̆�ed�-b�����t��`�!P����+��~s��8оG��q�yzl�ҹ^n�UF����'$d�j�����D|A�F���/��Ǚ�A�k�G~>v��އH Ѳ�>?/ٯ���!���G�@��^<//��B���o:[�"�Y�w�Hg��AD!+�"b�R(��1o�Fr�!9b>A�/` ̈́�>�m�(�0�k�T)�Gf���<�"OvJ%�ݳ|�Ѻ�a���4�a�,����|#4>�����N����J�6e	�zJ��rzӫ#8�b�����<v�x��aS[�D{��٤G5���<[�Nz=w��`L���� Q�0"��7��f��Y�[l�s�엹�	��1�3��ao�7��0Щ3�tz��L��}�.����\��n���,���H��c}�:=Ί��9����>��eo^�������Q� ��y�d�Z:vE��{�θC&�u䲚=�V�=(ٔ��Zk0\�m��O]U����0��V�6�x0�ѽC���WX�T�!��>'*��{}��;LB>�	��/�7��������l���+�����=�����UF�[�[`�|�����~�^��q��Y�Ő9o��
T���){ʹ0���"_zk��3��.{�cl�,�n��r�Ĭ�P��\Ū���,��	|��^F7���?��G����u��r��ߍ��W��d�9`s%v`�(��5.󙻘6!�b��=LH3.��Փ�s*:�y�ɘ��T�Ș>�����숾/5� ��L�ҷ7Z�Q0;P�=�r��-�z`��'�30��_L��Dţ�Vy����[��>~�o~�~�X��~���@�P�.��e<�t�̼�?N��}_}��6�xƇR��gֳ�w�h6F�%L���(��.[��3� |A���'�H$�O���צ���n�T�%�YC��ﱼ6;,����v��͘%��l��>헢��f����]���͑��P��o������3\��x�tkJ�������y2"k�;�����$Es?��ww��W�v�KG[�yA��Y	<J���!��g���s�n���U&*=M�q��>��O�$��?�O߹����=������-�U�yJ�*�ҍ`�o>��D�,�Xmj@����ju0B�V�{�CjW��v�?f&�9�&��Ê��b`	�0,c/뿬'w40�YIy	�u���3a��:�Ex�ݣ���;ϳ�f�ϟ�����M0�"�}����߳0)��$�}@9�8��nӉ*�ن��&���K���k��
(z�S�</�����jV��'��� ���=b79�����Bra��F��x ���5��KV}J{��� ׼K	���v�p�J����H`A��L��އ	���Z����h���W.�~ zI!�	�HB�{�=�>n���^:��y��CSw����c.�<)�ic��l����Ir���0�ns�:�v3�ެ�����Z�v�rhO$�3<��|լk�&rKR���+��O��N`ǒ�v���S�*��>��*��(f�}����7Ѽn^1�^/�l��k��dy�A��zt�g"�:1�J�DP�
�U�U�sC.U����^�:+��{]�<Mr ���Q���]gV>K1/w�T��HCH�V��_��E�x����rŬ�Ř�4��DG��R���FF�~�����������3����u�q2v+qƧ��eG����UK��0@{ѷǇw'�P�w�"b"D �R��a	B �@  ���`��$�_��\/?#��������"��:P�O]}O��dBڧtҽ�1��&�� �e��5잡��'�m�o�i�,z�y��6��nmco=$C��w��A��ɺ��^E-��-�V�Q�
�m����
ѭA@T������,DR��b���l�Y�ed�X�Qbʪ2�(,cE���X,FĶY-#*�V%e�"?#�/�xٯ{*pB��NGΏJĞ��)�ܴ4WV��kfu��.T����l�:7�^1)�7�wfr|uu�C�*�+�����w�zӗ��̯q;/E�DP|%�Q�v^����+��x}��M\o� <���g�����9H{0���3���hX}�5�WW��<!����P�"�A��(o�#�G��Dvz��fי�wC�[��:�}Q�	[SI�=�t���� 
��'f����/7�3��sؐ�'����OTA���� ��>v��/����{�n�v}d��f%Y��IcT#�"�0��"!��J�rl_�r�ڎ��=�x�r�o�2�8� {� ����~|5e���y(�Ÿ����]����ׯ���w� t��� DN���P塖��@���z#a-�,w�jZr:��$6o��3�|���mXt5�u�??� ��˛�+PO9ӷ�hJ�h� ��Ԍ�1� ��{���w���5�؏�!�R (`(BAd"sf{�t���^�~�S�v��8�.�!��:���U��8�������^ͳ�{�ĭgvGDd����̔ul�j�9J����$��8��}��!4� �-8������Ê�`��];������Ȧ}�9��+#��;�sΑ[X�*���W���p }ǰ,���M��7�%�����4��!>%�_�\��������Ð3e�;n2z��WUb�OP�"�BCU�b:�B������p��-�U%�K�-�r'���\\K��5�6�a.��v��+�����V��R���#��t3�_��{�'�`T9�.�a��DHH,� �B
	A�򞙉|>�ꭿ\��oaUV��_ӈ-��)�z`WRyD7P���fv/y�����Z����5p����RݐˇG��)���Ss~�%}�s�%vP�L|i&�w�3���+� K��H���(z.$�tQќw��g��\��<�|n����3� ��/~W"zoƽֻ|������E�%b$��HVBV1�
 ,�Y%@��T"� �X�g�j���|�)-;zl����wS�ְ��NAX�,�0��L���ȣ�q�*fDϩ{g�=������C4om̽3+9��'k���A-ZG�Y%�j��%����(0��-L��OT�J�G����~"v�;�=�8k_�$�� �m�����w\}�2�a�/��Nz�2������}�ϴW�z�o����!?"���
BjzdLz"@���䷧�����6=��:<Z�gq�rI�썬�����/z�/D��!�[필���&P:<��\�Ӫ�:�~��O��p��G�5_C�E�ވ�@]d2]ЙEbRT9~h+���}���g����j�'7p���ټﳠ*A��Ȓ�UR	A�"��(+aQUE�UX2*@�H�@�e%�ܫg{߾hy�0u7�<�k�P7�Tt�X��4i����-.������7o�Ә��ʉp�Ĵ��G�n%���Y�M�X���V��D=�E�c���s�w��!m\Ĭ{��בym��+
ŭilX))({���+�Ӱ��]gA�3���e���>�VƬV�+������e�{��1��8U=M����S=�^����μ�OŔ��p�gmk��<y��a��D}�z#���֖��Bw6�oۿ;6�4���"��O���%��@X&%>��z���fF)��U{9\����U��(�<�zGH�航��S��$tw��o����OB�7�/��\*�
`59C���sӀQ�j�=j���d��}5
�����!N�L�.=�b`,�	��m��r����i�������ߔb秪�7��ޑ�v E�b��� �Jr2�4L2	ɇ�0syUg$\�R���v���Bc��[������vv.�[W�a[�R���]�w��P�^ϼN:u"����^�N'di �0�
��~�SB�=����}>�E�f>1G%XS+��u����~mz*��t�����HGvA���}U1o��<0�D�'F��05d�oy��A�\�%��[�s4�ݜ��q�O��:g,'tU�0mNV��#Xnp��;)b���wX���Υ��'1�N�	�y�t����T�7�ﾯ~��E?'�_̲��!I�(f\��!��.~�鲺t����8m�S#<�X�H���ͭ�4��:l~�%�Q��3%�艼qt|>�*�"����_�n�F��)��w[���вd��v6�^�*��do�ЧR��O�
}��Wc6 �l���$�2�,q+$�څ�[^6��^��9��b�b�h[���Z�f
��$�:�,10|���������1��r�����M�Y_f��!�Λ'B�`�*�/���6��ME��=8Ƣ�2y�	�9a���ޓ��8<;ί�l����"_aq�٢>#{�/�/&�qс���� #,��)Y�*Sp�\�a�4�;�5�Y	�11狐	�ӌ\;'�ޅl�MLd������EZ
#E�
��#�fZ#��̜)n�/*K�s�B�S���]RX5u�Qz�5bwąK�LT�w�+L��mp�R��5��9l���Øu�w$2����T���@���~[P�CΉ��o�R��q�s_*uӇ-t��3�&�N0F�t����AҸq�v}�~R�w���Ni�1;��Ǫ�U�֫G$C���BȨ�W�w:q7,�k�Ny>Gįd�\P}�*�p����y��7'�"�!��mF������ǹ٢_��{��N���'��&)���E����ό>p��Κ:ٌ�ry�E����n36�ɵY�����������~OY����sn����ʴ�cܬz��q6�L>��E�[��Й޿�y�?Di� ��:�HQ$PR,1��c��x��F��������1�7=�M�ԏ7u�װc��iy������R��ӊs��. �5�Ρ+}}Gv�����8�P~EKwU�9Lz�`�.x�W��_�L��=Q�J�B��-�X�<�.��|��o�Y���;�A�n�V���cDf}귘M�W��WƳU��k�7E���U��@����S��to���e�+jV���̨����)l�ZR�q�1���D�z���4�-���LF��]YI�9tZ�c�ַ�(eܭ��9����(���L��ա��MkMۈ�؃�F��/0���Wc��k��Rj��\�luf7vGku�ܮi/G���3��ܚ�[akE�T�*��b�.'�)����H%��9fl�m�B"j�K�g6ٶ[v3Lit�G/�5�am��'41�0X�h�ˍ�mߙ1���:��f�B�8�f�;��V����x���t9h3)���@���A3O�Mi\n���D'ĺ�4��l�_%��{�Lr�^fukR�
�����}P��~��,�]�2�p���6�o!����QK��>�y(�IP��")�
��FBF�ơq��V���(��ǕI�V���a��9�K�zT�4��W�u^�Z�%��J��Q�U�$I:q�8G=��t$��t�XK�������35�a[L�K������n��9�0=Ҍ�CY����m�|�B4
�\�V;]��U�N����I�:!��F���B��%�$[��()i&���H:�q�c���+k:%֩n��\;���&
o#�L�y�`��k��A9x'T��k�{=���=�6�T�ƿk��M��ܪ���pe�A���w�Ī�8�-<�$JB�'������N&��mG��7z���K��V�T�Pv2�]+�p�Z�Gwj4�ei%p�+�V��=���=���Ļq���ݗ�>�^3X�9�Gv��K>�H�6���ұ^\@�� �V
3m�et�3��[�o=|L��������*�/2��67��F����]a��E5$��H�n�܍Ѣ������s��A��o,���&����1���Q��P�HAz�htك�)J-vw��mN�hEA#d�Qw!�ƙS0C�E��pڡf͙;.��Ţ[�m�QKm�ɪ�-��F\Z$���h�����,d	�m�j4`\o:Tz��<�?_^�����ܘY�+���m�vk�Yw�6\�����t)�,�Թ��e��<2*yw"�̆�NV��S�d̩�ޥ�0�L�'mVU;DW�JRh���b��{��U���wc����.W'M��7��N�����l�ck�^��	ݮ�"RoN�s�jl��5N����V�=Itr��|P��G%�Z�]_��>Z�U��q��t�e���gn�n�D���VR�о�{��V( �l�Y&0����>�~��zTt>�����x>"�U�H�߱�3�^l;Ng�����S;^s1�U��U��T%�&�Dh��a�#�0M�~����?���Ks�Oc3 e��HR2aL�s�\�eR�I�^�{m�\!@�����sr�&�ݩ7�1�舏mW�K�s���&��׈��/����-��']�р�׶B0WN�`��^�U��}��S�e��/�}�̘��A1"zq��O�u(gw<ח�:iv�R]��w����7�#�B��H�����G��.[׻mv0U6�p��������.���Щg;��1���)���.l�R�_Y��&�l�&��,ZX����֟��.��xI�z�DF$
b���5�������qɦ�\�ӊ�"����P�l�%d���rFU�g��֋�޺�2�Y,|�.��H1��W��Bj���;�ꏽO|~��*r2,��|J�B��B�(k �J�}��r��M/�*�{ˍߤQ�H�� ����q�}��
(���Aa$�� �a&�=��{��7�ן���u��ڂ�v���'Z�6z"�ش�Q��N;��+|����iʋSK�5��#˂B�CG��43<����X�WϒLMÞ)��g�Uu��vt�x#g�����,���%V���^����dL��/A��{}�2��T��\W�ޏz;3�A������ۄ}� 7l¦�!��'�;�1�F�Ɋwz�W}P�S'��2v��r%J�����?�ϗ����d~T�_��ب���Q�f-pGH�-\o�5L׫��U=���,�  Қ�SÏ}6�������#}�~ &��<Z|�s3_]}����l"I4�T����UT�sY����bG�ve�#kE�mnP͹�>X�f�e2�+`���P�kC�G��K��sl����wt߹��|$ީ}[��;sOk�Y"CQU�"5ٕ�.�uV����:`� s�/-(���DFp>�G����;+c&�o7E���ȗ]�Jo{�z�r>P�kJ��O�Hu�<A�K0�F��c�dG��JA�Z����x�DDp�=>ŕ�@/����eӆ&\��aҒ�L�m%]a����-E��%�����lFL�f��`SE\���:i�4Z�1=��D]}���oꏣ��0xGOp�F�s�ŗXѧ�!S63����}ԷcQ����.Õ>�ۂWQ�V�Q��.?���� | ?�/ݢ{��v��G-RX�2sU���|�k#bM+��Gs��&��6�S�k�<�,�=6l�w΄T Ǧ�����>���G���w1u��w�L�
D��ix�ϔ�u��id�u�P<s|���>��"�D��(`@F�%Tm�%H�u�<�]o�1mmz�U��;�)��U}��VZޮ�5;:�J+�
�36�t曥�R��r�-s���8�fd��yҞEZ{�ol]N�,N\}��~c�vY��q���g�f%�}.�B���1�m�V~���#���k.>����	P!KY�'���x�Nc�cL̦^�M��u��з*�N<5�z�.\!�9����z"��VT}���0ߠ.j���Q/�k1��r��äB@H�lP#][ө�~xY^gs�����=u2w�{z���}s�2`+�k�L�Ϣ g���E=�=�	��ݻ��{���ùQWa���6�����7��)tCҵ��s�M`���V���ұ�p�BJ?D`?!Э���~�XN����u!+Dl�B��5�������.��iJ f;ۉ�߱f���]��@$�-Ɉ~���͂��s�����5{jr()Uj%�]��P�b��fz1�B�!.v��%��`O<���rMDFH�A RP�RE�������}�ｿ{��߻��ު{���'ݵ$����z���8�l���ٮˬ���,�
��{��4������혧|����*�~��yl���_��p~��Bs�[x��x���>u����yM�P�ճd(F�ڒ纁}!��Na��f:���y���gz&}�'髎��;B�ؠ�{��a�1c{!�L��Hf�83�>�ݸpc��¦s�����"�K4C=�&������؟�	����J�>�L?��3���:�0�U��F]���.�"�y�{���r�ҹ�jwx@=J�J�z��Kꌎ�s�_�j"w<��n8#r�R�
�ktץ�Lv�'�MMbt�e��c����X:����y��!�,�0�}�u�c���1�V>���4��Z�}Do����bf`�P̻�P�*���oo����u:<�:�n���y�/������@��a�!3�����.J�d���F�/�11���tj�E�$`�Q�JF( ��
�,dTH�`(���]�w;�����y�q	$�j{�<�4��Էԕ�ha�O���9�&��`�Ti�ͮt�X�{��k��6�so$g�[�g��\�2�e�걪��f�������if�[n�:���F����G�X�v.�,�t��4O�ǥ�'l9ʭ�k���+`��F��Ւzr,	S�{��)�1xW��  ��΂]���2�m?�����D�C��؁2�n��2��r�Bn:W�E�CjV��s�×=o���S:t���P���"\����]x����LU�k�@	=�B)��o�5y't|aeD9��g_FMF�f��!�u2���*s���g�و��w2��<�0�uί�1
��A�q��E�"^\w��'��0d�N ��HC�A�:.$OL u�y��v	0��X+�]�4�(`���[��Ia��@U����՗C�"{Ãu� 	J&UF�aS��������`���@�PG�IYR���}��39��Κ.Ͻ���꫑b��\7�4���n���7���e�..b
U��T����[��m5v��ظ�[��k��y�m��Eܬ��z:k��o��w_.-��}������I�����+o�P����2}US\�c�׆٣�v�E�c
��+�!��p��(O���l�xV�_W����b�����O��	#�z>ge��R���0ʢ5N�N�1]�ڳr���UL@�j��Rnh��p愄�r*9ڨ5�{jU���#��~j�w����  /�{�	��G��ݎ+'�Di�=��w �}W*��İ��MFc���K��ʛR����{Cѥv�mKN�D����ޕ��7�ѧ�rc&n0��yT��P��q$�ML�s�Ǻ,��[0�*XOC���*e��R��������e����>$|>   ��N���+�.�J�k_~1�.��O7�̉E����:Ob��vRLc��]�Qz�	��]�>��߯�k_^��H�9����\�\��Ys�uN��H����2wmo^����yK��Q���P�ՅI6
���%�p�������2ۮ�e�Ρ};�{�B����K��aF��Ϩr�7H2����c��/���j�z�^٭�0`�9#U%e�VLwP�Iީ�sވ�oފo���D}{�f]�$m�!�}(������ᴩN�s��"u�BB�G�4�S���/[�(�VH�J�C<�"E����G�<��%o{p��Q{st{7� �3Oվr�%Z��U��{��q����>K7<�0_f7�����r'gx$�u��kg7���&\���K��{���_1�k���e\���X��c�F�}S������3;�=�\�/u�⥌{c�A�:߆�u��q�11��+��!/R��z�^@�f�S�Fjņ����w��Q���΍D: ��������:�W
x��T]�?3�*@P �7�����W�i�~=�G��=�q���0��eaR �	'�5�����`��ѻRh���C���tJ��J�p֟�^��-t�Rt�`ż��|wunpd��@Fq�q&4=�̜�Z��*W�z��+����B'��0���9�Z��S��Rf�oHE�ӳ��T��~�|:
\�g�}[4����ʭ�H�ٙ�HKV~3���frW5��9��&o�w�Hq>�6ob#ދ�s����)�y��/�����|X.�P~U'/�pɎ	(�1��r�j�-�y���b��� DB8u��egK8]Ew��!�d�rQ��l>��D!Y{[��	�#l�0/G� �늙���L]�(���0�1;�5Ig�������~���CT�s���"�@Y"$Yϭ�s?h׽�Dx��g쯯zq!�mi��]9���g���\���l�����K�V�-FM-y
�+�^�q�{�ml���]�x�_u��y��23B3G�P�TA�T�����P�Cjl�iWS�U���H������������emx2jj7ԥ������O�Le`�Ծ����^���}f���$�|$�Zus���������m�[�4�B�5bJы�R�@b)F��&�S��l�@PFE�$�'�'�H ������.ۯ_���S��W�^����O�pF3�DWw�7Ρڧ��� �NԭĚ{]�y���;�a�z��j�_އF�$"���'K�`��}���nz�v�7D�%�G)w[4z��
'�0o�s�!	�Pq�֭��f��Fe����:����G��T���(LΝ�Қ��t��ERi�>}�����r�9�zg�a��}Kqȧ1<��x�K�%hM����s~ܱ�c&�߫?g����&dg��	�/:���19��0G�H(��C!�\�I�f1�P��Kh���/�1����pS,8���1��_E�F˓��<zQ��ޡ	I��.#���L�{��ڮS��{:^s�L�Jޫ�gЧj���w� �c�9]P���F�~B����@���0���2�ڠV3E}��L�~�Җ�)
��Tm����|��_��E; �~��� ��`�-�9�Sy��e�֞ݳ�v�!XK���:��:Pe�0/��Xn��V����]��Ff�n����fi�޷�(q���Zed�LYĭEC�vӛ��3���)�������n6��˪��e0Ec��րٳϯ7�p�ct�@��0��0cl�xs&��8�ɭ:b�E��ɥ~nj0AS�-�ю�Z��SG:��4�P|~?�Ub�Q���3j��yR�H�p�k��Ҍ�x��sz���z�F~�Xo�f��5�_
�4QB⭌I�?�$Ab�\S��T�v�׈�)GK5�3i{�e?��/,��d'�B���E�ܦ�r!HQʺ:h�1���J����dV��%U�md:ӹ�a�لot"5���y1N�۲Ѯ��	�*�����Ɩnj�([Q��1�-�"�M��a��xV`�7zci&{�w=���n��m��
��f>��N��w�����w�TΩ��٦�b5�K���֩F�TjL�{Wrc�rI5����&��%��1=m�t�e���v���=}�h�L:�V��Mti������FB���Z"̱$;�
&��A������,�wl�n��D�w02�h���,�Ju�-;ղd�8���4�ݺwZ�mX���$J$A���X��<�Y��B9���+�֓0�Q�z	S��;5v�Ǝ�����F���)���_M��T���Wc{���-�߶�y%����effj�fn>
�hQ���H��w��L���o3ˇM�+��x�&��ҕ̑ǜ��V��IMMB�ҙ�VZ�潝v��������t{^I	�Y��F�Va�NΡ^���AJ���`�5�5�(xنTλ!n�-"At�0�����N�ED��Z�Ev��l�Xtq�SR����05���5��S����70���s���tɝ���Pͽ�w�ѹ�;v��N�v#)Q�nK|�A\ �����2�<+�+즻�4����qا�Ֆ��hN�5�A�IUe/��yՐZ�k{Z���[�ئjo�^*vm����˜b�j��m�)��RL,Wr�6��I,�܇^i&f�����݆��u�KW�ؙ֫c��ݻ�]��p��;Nq1�Y۳��l^�v�� KpU��Ĉ0k:M�@=�nʴ���ß�5�r�aP?2y]��V�޼���la�FU帛]yS9�3����)����k+�ɏsbE��������> է? �ޜ������Gp,Ho%�ѭ���]2�e�PFT�bQaĨP�6�T�6e��Y��_� L$_}yc+�Ѯ~�j�Rg���a�#{J�XPbu�0���F#�َ�`��r��7�֪��,9��^sU�]�@����(C��痂�+��J��BO����r���;Т���(�巭�Ը�샍�ݕ���F����V��Q8�5����V�Ґ T��	��G�����5_T��L���Tކs#cf�o7���Z"�=�^S�)��n�`]�	�+�;�겕R���.�&REs4;@��_�z
0�~�x�~ך�]~�߱{���P��H���>Ke]Yu��|�����>���d�V�q�!\��b�wR�����T[dT9	Gk,����wl�����TS{C�ol�;v��قF$(-��S0�Apjzjs۶/f��l;��uL��v�B�U6��@�F�y_P@��Qse��ll��m'p:O����2��2��qZU�t���vΡV\Ǳ�l�>M�+�fX�~)�v���y{�x�a���x�zu�\��"R�Ϥ��V��i���X�������[��msW�(��_U���ӓ{�pR����<�O��up�;�U�ʡ~�e��W�e�5[�P�>s$e����UW�hȕ0w�eJ*x��1�G��M�)�����q8ng+h��w��=x�ݰSOU3�l�����a"��1&6q<��sz�����жm}^��^9��������QsV��C�O�O��mUta!qiw�1�v*���}�}���|'�+�  �>h%�""�)l)X�Q�э��
X���Bڰ�Z��K+#"��d+b"�X�,Ye�,���U*P�T��V�X���Nk�}M�r���#B�P̙ü˹���Z:�3����z���]4��Z|�'z4	h�
�P�F�ﹾ��sf�mN2�О���[n�)M%fy�O*-'������~$��#��r�K�1QH�Y�
�9��7��2n.��c���=V��e�6��:�轢n�{D��}��",�?||��,����Y�\!I��f�FK$��NtY��Ȏ\r%8C-U'I����{�41���S�T���n��8�'����=�/>�l?�%�D?u���2Y�9����	��έv��	ץs�r�%����>�zf�(�V��N/Aw�|˪.x�|���`���Gnr�B�tٱ�o{�(��:��µ��ߗ�OsǬo�Gv��
e�f�<��_d�8����?}o>��gR>;�h蚉�;&>��a
E/��"0B�1�I��߼����lA��b��t��ol���Ш�v.�cˁ�~��~ |I?H�B�������}�����3�Ηv�y�F��Z��gVeC��rs6]S���[��}��l��`�;�ɝ�3�H�p��)�tVs�jit^0��3q1��W�4F�����{x�{�����+-I�$��Ļ�AKA��՘�T�e��7��4��vƥ�N��F{��,>�*Q]F@�T��*�N�p�v�ʇ|��s@�*���}�=k|��W�����D�.�4�ډ�vzr
#z[}+�֧�� �QT��V�[��^2Z�k���.i�h��Cf6�Hgz/-?:��B,���>�o�>�_��;�f��|>����9�/��5GL�v_,Koq���~%�b6,:��n*���0��ʜ�P:Q�D��Vhz�[g�8���N��6��-ڷ�L)٥pU��t9�9V���:�m�\��G��d�-�B���Q��J��󟽵�9-���=G�b E�\��f#�~�yDdI$��"*I���Ɵt�����N���|���w��м'"��b�󝺭�@!�N<L�%�����h��+����(6��oLQj�Û��/\ݻ=���L��H)XH�n1�y鋍]�C��0�f�<�+Mh����������qL(+�܌����q�Ξ
�ǦJ���J;%+RfF��Y]��*�}�^���`�	  >����~�-M@}�d�@�_Ҽ�>��c������Vޱ,�|����U���@M{;ʳ�҈^����y���z䣍�|Z�? ����(N����y���]G,�4�6�>�b���y_�Ӻc����Vyz�/.���cå�Vz�� �͹@HYYN��F�A��z/b}�yLʶ������Dn�V�����)n�I�@I8Մ��	�|��5�f���lΑ.��`f�zc��)؂����{�������<o��;�cK��h^:^�_�艅�T�ht��/c]���9{�| vZ�eYe����ݏ>ߴ�,���v�\�CzVWV:�ΐ��mV廋��#�2�E��[/�h�Fe�x2#�l5O�V�|;���I�AݚE+W9��nD�̧�t.,D�7��u��AH�X,>��͛�W��a�K8W۶�����rpP�X&�Q�X��[���;#cʝи0"XaS���k�})�u�T��"�%�o���/��+��MHf������A����4�{p�:��sV�����g�j�;8�m�Ǯ[}��59̾q����Y�*�`�����0Y"�#"0RF(�"��1b*���ut�3��&���}.�\n�ɋ�v)O��D�٬������Qu�v�����2����84�:w���~[�,���1�7�����?/���c���@�)ו|KK9�=�k�����S��p��C�c��/b���Z�6v��K��B������q�O���-�4�Л��Ɖ���D�_�9L��!ޗf��j��t]���2u�#F�ԝ�SBK����Ϧ~N�5��~N�������d��=���-�%W�z�8wk��גK#��W�)��&0vv�A�U���)N7��x2��{'6\��u:4��<�:�^'�̇:�#p!�1B�HtB��tw ��4��-'=�yB�է?9�v��iGu��gd]��3��
��i$�tŹ�l����Q��^pɯr��w~�G��J�1�)ק�"ɆC�0�u��W�6N	��:�����"Ё5�&vl\R�g�{��*��W�����Օ���x�或�D[Ϊi�9Ն|؇�������֡��ɼ��v;�a�|ѿ��-bܴ)~ g�^�u���9~��7y���.Lys1q�톕o�V���寢�ˁ�I��O��^ƞ��<dGߝ�����~O���8�/�3����NH���ΐcAzh��)�\M(����DGKG<�.;[2\*�	�t�=��	է���G��/�����J��i<0���U;��/9I��$�F��nG����ՙ���E��V�-��E<@����i�ZU&;N��w��|��M �Q�~��+K����lե��l�A��vE;�2m�P�u�z�Я�
��.�ڇ{�m,��
:�B�Ξ����T�t�*��.�GV�X�����I�8o%�w�]��8�̕p��<ʤܸ��2#����UV�ە���.�x)z�T����@P�CDt��gd��w�A�ݥs��˺bBnnGU�s�2UM?�"��ϓ����7"�$�z���ПW�&�L)Oj�F涥H_J̡��٦?Rh��Y4	�񴛥��~�G'%��x��|hx%<����l88�9�C�}/X����u�|!4��6}�[�p=�v�G����TB<jy}ǁ�&�p�	D���z:��4���㷠�%�����6���=<��Vu] ����%j) � ,租o���z�^̔j۽����9wa���p8b���1����g�m	 �\�]@Mj?�Z�ј��q�(P7��rK��u�W�t.�c�Lhn@v��g����}��yu>Bq0Z\4-�$;w�DD{�Y�q�ח�Q��lFMؤ;��uK��b,�*$LSf�+�㽇��\(Y&�Y5&���5h0-�DM(2��+H� >y�!D�b�zg���شؤ��4��}TҬ����nˈ�nd��88rbQ�0�LG�}凭i"u`d�o]ap����ζ{ҍKM�RP�g���5�8¥9�6QP�0.&��%^m����&��3׺`�g�6��>��Vo��J�b3ݙ��7�\�;�hu����5��P]��.��Ϛ��<�����y�|�>� ���9�چ��2ۭjɱ
�+,Put�#���\�ޜ�(h� [�K;)T�À�"�,�8��Vr}oI}�OscO�����3`}��H�	u�U�f����{ܤ��ۤ�Bt;��mǪN:�3�Sz�9�W�9Y��;��0bp�&ٸ�����6�����]���:��2��Э��k��*F.���V0�I�OȺ���B=ڋK���x���`��\�MP�6�^%&�½�G��J�#%G�\?����q|�����+23Ț|����s�7�%�9���� �n���]�3�M�ƾ`3����5�8��y�c�E0�S�؅�P�5�ψ|�%xE����3R�����˽�<��+�M�I�}�S�( �߫~VN�;ݑPW�� ��3n��?g�� ��4����I�]3�����9��:�~n�^¹�>��;��ɐ&�e����΢�N�\,5c�g��*�VQ�L$Yz�-���7�x�疇b^Txj�Đ�~|;���xk�A﹧�n�	��ۢIei&W��	�qֹ/r����u��^�
�����%�K�X�/�E��K��%Ϸ3�o`��²�a|�,B�%Rdq�܄om�v�Bl椷�|X�@� r|�O��Y�~Zv�cњ�I4�Y)vjY|r�����V�B�*� �	�T���e\tc�#�⫌��(9����hk[˄����Z&�b��b�<��h��0D�\3V]��d4��U��Lcf)iLˋ9�4�TPV"��Ym��cr˚�-RLuR��3�{5��j���1��30SW��"A!<yAi��Z��$���c$t�Tr�"�Y��m�M�f�T�ۈ���	�$2A���1�k���h�������N歷w4Ե*�jh��6b�.LI<LLђ�a��\)�F(���������7op�MDܦ(,0��hNj�1חj�h`,Cu��V�\q5L馊M���bcT���&�TF������l֥��u�Þ�{7��0Q��g��ߔ���s*o��I�4sM=}3L�x���ӧ,Hg[��[ki�W�5����պD�G�^��n���-��k3FR�J���H,
Hm�i�­m�Τ@�p]]�$!f��ov��VV��I�k.�U �!�iSW��K�XsX[г�SH;	���]�xs��zk��$1#ud��Z�^h�s:󦹦�!�[�2J)
൷51Hr�IG)I�M����@Y�\����*O����@�/M��~�ѕP�{ҪPǂ�A}챢C��}�r�!��u0M��],�ͧ��k/�A\��bj����F�6�#;�ZV�L�\U���t�Tޒ�0��V��N����kbW�L͊!֬f�۴oۺ��y�4w)U�׍\���'GѶ�k�T����VrIRֶ��t�U�@r�<�*vg���b鮒SKv�dКO�K���7�+n�y���U+pN�7�M�m*�\,�0�w�T�ݗ""�:���@�-�kM��{���}��[կ�Ç'��$1՛y��:m�&T]gQ�h�x U���r�ݱ��	J8���=廹+v�Jb�ݹ�x�;�hC:�J�+
�}�G�TMk���f7Vͬ�E�m�ũ�,�d�Zzcܛ��&뙵�B�鏹A��wWH�[�,���r�k���I�Z�ba��^Sˍ����u�=�ǃ(�.E�GF�Pe�i&.��ó&MT֫��s�hs�\wz�.O	���V%X�>��=7]��a��8��B^�t�հ5����9��jO����Ż��]��m]<J�������d�����77��]ʻ��p޼̼Ĉ.�o��Q��;4`��m۽���\i�d f��)X���iR�U�V�;�2�e.�
;��vM*�Z�T.+,Tc�i�ַ"�'��q
���5c��
���м�i���K�J��霶j����7��y(s�8�"� ;�b���7�����1���L&���͂��H��;w�k�q��>��:��7GY=�N�Ģ�#·>��*BD�9�#J��
��׵� Uٵj(B7֬��o������{}�	t�[�)���¹#x��(��|눎H�s�(�͇V�mJ��l�$e48@���:J�L}���M*�&�3mC0@}JW��T�v��Σ|/P�H�b>������9��������֙�p��X�A$PE`�x>s�g3߾�~����߽�`��4w;)��N�>����U�t���{������������f��z'rE����f3�������&ˑ��W��f���	��Y����䭆MI��'JLE�]�>ɤ���&�V��w� �y���Ų�1N�'�i��so� }��r������b���T标�Pض�.�遦0x�v,쑸��.�	M��0�� ���}����B+F �~�n{8�#}�Su�1�ʘ��aMZ2�P�j �6�s{0x�{���
��(�e[a+"*��E"Q�d�HU`�1UE���IX*��E�)Y�F
DPUQcej¥DU����ĨEJ�2ڌ�X�F�U  �NVԚ��%�+/}�rj�meep�'��/V��.��d���'Q6 o��6;�hВ�0�<�J��-�wJU�wo�{r�=��Gx�w�����^K�_�s��gc���[}}�tY�v��E1��MZoA�����Q�Xs$w=ӓ
O�Io+&ڱ��� �M�ϠmT�����?!���a�R�� zn���.�=.nk��%��x�F�P2�����'s�����I! P!�5�َ�0�г���tM�`�u�_b�^�Iqp��)C��H슼��@B#�]:у�\�<����+�7�I0��ٟgHtɁ�yA��6H�����o�\#Cg�1�{���~��=��x�Ǧm�.�����~��ӭ3�!@���+�;��^�+=U"�Y�=nxF�GňLi[Xuo��V�q��N������3]:e����q��C8�~�y��wY���q ���>���|{�nx[��f(�+7�'v�w��sN��d��ݮ�6�n�h���-˓���a�v�@vs�I��Y�o�)]4���C5_�r��C������.U���
&7)ӱ�Z&�dJ�=S����}��K��r8o��q�0%�{!������RV�.!n�3��(�gW�q1@K�ć�uZ����ۙ�F���؄e��h"_���18�g������3{��k�a��\<I[z ��-� d�9����8����}�q���vou���7vy��(�.�G���@<�LB]%�W ������,��Hl�Ʒ���5��u��Jˤ��(S�^:Z������Kېh�O�}a������_�0�!F�z����v���gP��/X#�l� ��c5������{��� �ٯkRx>�ũ|�|>�x����C��4��w3���T�ޔ����*�I@R#@U$P�Ad Y"��-*�DY��y�/�y}����q��6ociX}�n�XF�#��%�\�����sT�x�U����k��i�P�N�ޘXrh�ո�5�lk	U�Z^��ܧ@�tzH/���f�@S�A�V��)�ٝN�������&�O� 9ODΤ����3[ć�if���ӗ[ȹ��0pbOI��sf����R2�ߖ�����}��}����"�����v\�=U=y���u�L6�.H�����wmi�]7��iA��H���?��DΉ}���}�8A��Iڮ�����C�/���V��/ώ:�y�)F��+����)�2����i��j���\�C�$#���������ƀϾ��?�ev���hγo޾����}�b�+'X%�	�e��s�Ӛu��%پjG�Jϩ3�u���_J�,�q/���,D�t��ݷ���y�Ӡ\rz����|X��67]�;K~���i��pE����`�:���B�2�����*)��nV�t�`�f�ܥ����zΎ�B+��
����2��������N��!|KZj���,)��,�L�ޫ�>�=u�/�����"S'�<��U�G^Nx�<8�SÖ�	�Q��T=����:t�8���-�J����f;B�2��֜�'L%�j6�I|Y��El�Xn�=�h�n�߲ }Wn�f��cT���yK|`D�Va�z"�1�KkӴU�H��DQR�H�%�;D������="{���L�v�j�C���<�͂3��G�z�f�r��"����$gT�)7~��
#�ۊ���礞@� ��^���#Ow�z}\K�\�[L��T���35cܣ=�s
���x��$XE�d�5�� ����v�B��p�}�b�	7��
b��v��0x�q��z䆥���[���L谦D��C{=��ߘ�z�����)��D���Ǆ��sw�$}Bݝ�X*��m�9�-��5r��!�_. q�F>A7��ݣ&Za��EZJ{-��a�%��1�./�m_��^>�\�O.�E����=>�_x�]Z)}�3�-���V*~�"&1H���&x�+s���lF��8�P��DDN!���l�.�-��s_r��E{a���LA�zW{1�f�\�1r����~�	{�+j���@_�b���
���޼s���yxzP4�4�3�gx�A��CUo��So�n���Gr�E^���@<ܓ� �;��q�������!QU/a����۱0��9I:�1�/����`�O���S\υ�Z]���%NO�p=����Uܧ�I��B�3������;ɂ�ZAFee.�CeFmU�tf�6�[��Cdp��ר��芛��7���9�5J�"w�DE�җ�b�-��9�q��C��{�3��?$B@A"��K�u���<�wrC��r�Fj�:P��h�n��݈�>�;6>�X ����u���E�ӄ��u]�.���p:�E�u:S�ܘ�5u�zPV@Cȣv�\pR���]o�^	A��ЙH@9�:zك���1*z'��j�N�.�����ʙ,��p��}ׯb�6��&w�����-�&ՒÒ;�kf�=�Z�R�"1C�a̤t�hV���)�k��A�:���V�z�Y���i���z��=���P���S"��Jd[q*�S�����q������u���az�
�L`����t�7R�xk���s'�kZ��Gqh3�Ķ��|�.��I8�ۈ����Sw����X���M��TJ*C�'D؀�4SP6fc����0�5Yy�7��Vv\��K;!�G�г��b�Ȏk7Զ�kأ픨�t[���;�����݄�Lx�Y���*�A��Ua���V@b�VB�Y ���,AX*(E�P��>#�l��D�����1fE1��oru���_uZ��:�]C^u������b����EM�jEu9���$�{kh�4�)��r`�L�:'�r.c3H:c��T9]	�����yI�rx���l���a�=p*��u�{`t��ɭ�{�!*��*�؎��,{]����}5!�u��z�p���Ǭl �u'Q0�`x6��vܾ�n%ij,.g,6��E�/C�Rh��,a1d6"�ޏD&�R;�:z��72�> |.���=V�~'Wz1[K��y�霚/��of�Zj�5�#f�bۦ�֬��lm����=���L������c�;��"���O�=q0�����t���tE��J5��S��T�5c�M�)h��P>6W����V���7���AB�EP`
�"���[����kp����yU���^ာ�����3r�be�k�i�މyB��k�����g��?��D����<u�Q��ŉ���ߞk;��`y!���"�>�����oݚBsnf��%Y����9���N
�k{�Df���5�\P�����k�������%3�㭤3Q�9Z�Z��X0��l-Fܖ��Q�?\7�J�R^=�$L:h�ٕ7���P�>���)S�V���M�ft��<�}^��3d�!�uG���R��T_G����9YN�[^�O���44Z�{�|-����qM��ן��[�FUk��c�)��y��I���<0u'{/�D>��3�\�؞��W���J�.2���^6�*��KϾ���V㨅�Ӭ ���u"��=ה-�42o��8"��o(�a�ǕH��n���Y�8����,Q�&���s1{8�������@���îʨ��X8��R�b{K�T���珤=��x\��{��ֺ���᝚�����7Ǻg�FE��{���)�f�P����q{p�����vpVx�TR��י�{|��j�}���)��ƒx�����\��/A���{τA�O�YuY�K�����t�ٯ_�Tf�ھ�$�̣��s{�7��x�A��o�6G��'{m�(d��<K��,�q�Lk���:>�@���u��^ՏN��A��]|�aW��2*�P�6�c��i�����ڠ���{�e�"��:s�ʻ�^wY=H�m��ο��7!�������:�4a��-˾M��Fq�ϖa_S���֗�=���b*:����cSP��uGP<�	�u�bp�`�r7Ӗ����+v�s��ɣ:^g���Ν��SF���zqfUY]f؋A�F}{�g�;1P�1=/�<���u�s=gs�,���+�>Ӱ9�.�ٗ�B�Ȣ%�0�ddo)q���x����KR�H_O0$���.�vq�x�n�L�Q�r����4�~���ݚ�,�BO�E|�ƚ�ښ�;whҦ"4m�H��Y���]��s���I���Ёe�yƜ�=zL��'���bG�k��u ��~�hVn�E�XkHb�(Qya�gq�k5���k�(Q8(�{�dPW,�\ug���Bh�(�S�QE����-��5���51/�lҵsv�lV W��Μ��Q��a�P��SEXJ�l�@�����0�(��o.�Bo���ek��ꙵ��aݷX��v��Kt��a[��n��陷�M�j��$C�#h���f}�;E	B�m$���!�]�����o
�S���u1T�	)dE��1*��B!�~DDJ�MT��I�bɌ�6Z�9��?()�EFW�*�]��6h��ۀ�A��1T�6	F����>:�?*���n�y2h��B�l�]���,�& UA<��P׉;���a�U��1i k�s\�p��ty��w8��L&�ެk/;����M��m*���g�yUL.���h�q*�p�"�U�c��ۛ�X�����:V	���劐Y'0�ۖb�Hq���l��WW�NK	` ~��[�h^��w��$�P	����6t��9�������`��%]z��	��^���E�g,6bٜѤ��n�ʠ��"Z�9��T+dۖ��2��,2Gė}ʺp�+3a[CU�2��Uwu���wW(J�k�h��� W|�M���Ϲ:�Z۟K��X�U�I��sFˀj�a��o���.o@�K�o+)���r���uς�r�_ΩJ|^��"Y�ܹ̬U��U0��C����X��y�k��eL���]�f���$�kfu�v��=���W�����cv���{h���wiT�6�tm�rSJ��E�WL���ǵSw� 68���$|;J�=�9��U��LuK��kT�w�Vw�c�Md��
��eCY�跻��%LrLb�I�(>{�oF��;?�]7���Ǵ�.��e�Tv�W$�6�drr"B]}$�U:�V�e�v�qޤ��eu94�����]��6<����wz���4k�K�۬���e��3��>���Q�a��L��xF����֓�E��v�Z��J2IyԈΛ������z����Z7^P�Q���#����Y�d�kMZ���=�Xju�7J�ƭ�M�K:���Z����Z��U���vT�MY{Wd���<zC��4O�<zv����e��n.����҇l��<7Ec�؞�n�BTfmꁃՄ�_t�;6漬�d�d��ky[���@�ڽ;5��ّ#����i����C�6J��ki֙Եud�V�d>R�zȗwò���+ξ���H��;S",(�W4�qX��������$V4�i��7�H��Z�]^`9�i�;��q斱q�:�<w]T����T�{��ܥx\�q��	V͂��+@�F��h�~�s����GS;E��c�S`h�س���S�m��Y/�����}9�}ԙdq�V����;�7B=�\�̐���XN�73OxJȣ�fGi�:�]q哺7�D�A���<��]�31� �7��x2�}�/�YsE���ʐ���Ë]�y�.q�p�� \�Nru�-�B��X����nn�̤�U(�+YsH(���������0�8E�.Hf&�r�Ď���l�3�4-�����t`)
k��om$a�x��\XC�/.pg{���(8�y������r��n4R\Ecc,��Ր���^UE�ڦW>y����U�^�CEzW.ޚ�5 ��v��[z�H��w��.��9P���,���O7����ٶ�����{fh6�j����.��(lu�u��D�(W��{�%d��v_��\��KH��f�,V-���� ���dK����p����o7:�2-���C9zi�I�y0���V������H,$'�]�7�{_�y��\���[�6�{#�)WX��tz�S�t�J��f�}���hm=���-�ݝ��,*�q�^p�q��y�"��*`�z"��z�\ ��nJ�/��4�q��T��-j&F&�S$ƹ�DDGӖ�{�#���>����Dj�Ȩ���r-{�(R~��A^*�f�'��sc'.D(���|�u
M�=u*�#r$�o��';Ǧԏ#1�X���	\>X��7{4:`�h���)eUg���q��e�A�9����D��� �P�M��؞>�:N����k�nk8�a�>u�(���ܻ���,798�T�D�wjl�z"i�u��CD�&0t���k &�t�[��c�D��'�5�}���s�aTLzoP�ˮ�:���9�ħ�9)�sQ��*��K���6�x�M\����Ltz=sK59�s��K�0*���
�zϱ��Myx��E�F̢4#� �ZUE-��P��!H�X� 6�d*�
����*�#V-J*�
1ly�Û���	�p����պ'n�ä���{��E�iv.]֬o��]kI�i�Q�R�ޮ�{�Q˵��%����}K��}�unf�U���(����7A�1c�U��O���,���q��-�u�]0�n�qu�/.kZ�D�iɓz���q�/���n�=vk��~:r�z����R�C�hv�rTG�7$������N�r�aKzoi:�=cì6W�������4��"+��V��C��[Qu4�e���y�8&��a�t/e�/��v�Y��x�8q\�V� �S��������Q�����w��Z�&宜^�K;%���V:�͗b,E��uQ��:o��z:��n:��Fq�ʓ���j'�(��F#���4�`e`��oC�1H������'���3���;�"d�Xj�p`(�ЫzyOT���kk�9}�Ҡ��*3z���Vf]:����^�t�u��m"2E��g�������\�p:zl�*�CoA�﹎o�j6m�q)�ty��3n�,�z�قt�}kv��.��gxG��x�i�7�P��Rw�>Äf��{��gUn��ˌ�D��1w�c�p9me|�<�\6�P�1����D��Y�"���)�2��A���q=�y�o�p���j��K�~���9ŏz]�u������ �YΖx{�\���m�:�M_kC�E�t{���}&�P�f�eP��y���V����d��	ۊ��[�7��X[q��ű�m�&�,�e��4��*�TP��Q0���{H>R8�W`�7l��(�\�g9�+�W6"brX9���إQ=Ɛ"p�S�Q�J�D�GbBo�y������d���|��nN�,��NT"��{�P��v�Ġ@g�����u9�!��Ab��)6�v��iw��4������M�����O�w����|�h�Qc!Pd�E#@X,"�AdA`�}Xv�Wy7 BU��]cL��svU���,��PK��ՓT6U7Hu��YQ&t��<��Ŷ6�w����s[׵����u]b>Ѭ�]���/oi�H��{��G���ևܭ����XXz�j����W�T����O�f1���$0Pb��(A@��H(��E�\s��A'mq�A/0�g����K���mH��c����:�~�f�\&t'���J�&\����\���[� ;E�8�f%vc5���US��q�QRDT1x�)y�`�"I��������t��3r���n�����_gvo#+���  �3�d�v��Z��ON&���*aa���E���%N`dq�����iJ)Q�Bu力,�]D�uH�-�o���F��5�3���k�7�1�8Q��wz�6>�l0�^#�lNf�{�U^�ܩA����59�z�ő��]�P����U��g����9)�z�v�P�>��@�I� �IU��:�}�F��Tz�cw�^�û;��'�g� ��� �c��YR�MYӅ͠�� �o��p�W5��Evm����s����[������d��'�SI{bI�:�ͫ�3���˭~�����ga,͡�ȋ����Oc�Av�N�"5੺�m��K�r)�6��8�{ >�B��������|+'�f�.� �+t7�[����w�?%�EQ�����,��+5]E�{��*�4z�(:�\�'oc����O������`q��mQ�ќ���K�@ѷ9��bAق�0����k4I�����U��4z�����.�Y��A���" b�EMu>�r�]��"sg�L\)hA᲼���1X�4:��J�Gf�/8�+�X7�B|f7Z�s-�D$�;�_��e�U��=5pd��d>����)C�vʼ�	C�&�g�*����3m��F�9�ѽ�՜���:���'AF�TD�DAX"����,"��Aa-�ČB�w����YW2/��t�G9�;���H2��J�'�����/O��[nge:۸�vab�]��ѫN��֞p�|�]ó�Q"������L)�C��?|==BΞ�trwM���BZ�B���q����ZFP�23`(aX�8�p��+�)��TW���J�@i,vPL��@p��!���h/ĉ �9L�<�2��Mt���Hz����/��1�f�r�T [���y��	$fj�R���;V��L�^E�����2��t�T[���ʧ��p��nS��P�q��ӢG�xE����NE�<hMʞ��z���[���7$�ፘ:�ͩ�"�(�I�\��7���/��}Z3x���:`*j�{�IYKX0��{��6.��<�@$����C3�%S������N6}�)��.Y&�_Z�]I�G"l�o53�9F��<zr\�1`8�S��x �n�FM���4=�1$�> ����������oĠ��»�=��E5�e��y�\��e�;��E��t����!�]�*!���r=�Ȥ�Ţ6e<y��q�ș����w�G�1��zwAB�xطIdj�V0�YĠzΈ!�CN
��d-.�\O�V��Pw��W����1��{O;�W��8�ˉ�ɞ�7K�#g­��[��ד���� ����ݙ;B��j�؆���O)�������bz�Ӛ��DU�\6Hz)9� J��+�h ��n��g�'��)B��s�M��A��IG��9�}es�_�K�^�{�X��̉_����ޣ%&�栵$��� }w�ͧ��D�n&/�Ĕ3��� *<r&"�Β���n�U�O]<�pW@SkO��!�:f����u.f&Wl�ƺ۳y�U�mAVF*�D �TB22)AdY"�Q�� �>��ȧ3t���^=���ߍ,����m�lАfW]=,"Ϻ&aF,X �,E�"���g����A@$޿z���sv�Jw���ea���4
�좕����śX��V�8Y��zmrZ�#>
�4����F+��p[��[�r��.'��N���,k����q)�Cta�8����;�5S���vO]�</�P�#	����m�*��ku!�Z��˝}��Ʒ_.��N���� ]��z�����t{��b�r|�Jp��'B�'�m ^���75�7ҡ�2˞�,R�s8�a��8%銪:f�:�GyU�
#'�5�*�m�1�{%�v�T��X���(��q���M�` 9F:��v���Ǹ�3%����^y",����6e�.����[Ύ��ȏDcZ��N\�D��[���U�C9�N^\Q�����LZ�����mF}�i��
��g�-/�zK)��ŏn��
�L\\u%��'�.�-.���Vyw/+�B/��G�;G��d:���!@FDb0�TQd,�m�D��*TD�Ԣ�#Z%d�� 4r:�wKj�����U���ٝtP��y7C��M�.��Җ�WQ�XpJ�';J\�0N8���g�ow�*|�9ׯ\�t��l㳴�- ��>��	0����wNHɍu%J��G)�J�
DΊ�g\��%����2�����X		��+|�vyv����{(��Fz��W�PK���Re�s�MV�Ec�K3A8J���oB!�^���y���q�|�ٓƱp< �
�������	(�rΎ�[i��U[������Wr��/����a	<eW�pI�S��ER͇.���b=��{�-�xcC��#D��h�o��sW�
��]	#=⽔�K�33[a�Nmy,��,F�dV�H������3p������rB�t�^�s��lb�l�Ki�B�>�-�J�J:fm��0�g��[y�[�:7a�,�)Q�!q�TQ�����i�ŝ��y���}4OÆ$�����W�Ҭt�|��n"<�nP���
��ۭ���ôc�F��m��+fV	�-5���n �E���p䨀��%�h� �y�qܱ¬<B(ri�@�!5�-KwqG)BT�R (,�RH8U�2�R�w[��Lĕ$.�5M�Ղ�g�^r�T2��u��os(Tf�d�c�$ὕ��Jl[a��iɧF��c��r:�FemM&a���\l��Ө\����"�E�ˆ�7Mb�d)8�q!7��՝��r�޵��t¬�q��fWY��J�I-�%���6��m)���^��iNb�R#7ۊ*:w�Zq!��4���4�� ��M �kvI�a�i6k�$��a0��J�̓U)h,1��HoZ0���dހ��b�!q��JA�@�aS�2���Ѡ�n��M;��0�Im6�a��M�����.�k��5�c��V`�j��m�\���m�u��7�@�(&�4���UZ���K҄m4�&֚���j��h�.�����tj#mc����P���Y#�y���l2��]k��W�dH��-�:l6�(PU�J�B�_�6F�]B�A���(��Y���8�F�,�� �T6���D�+M8���`,��ZIS��"���6)&�m2�L�+6���T�V����A_4
2�%5ٟD��:�X|����n�l��G��� �ݼ�loZ�;,�5Vb�	���A`�w���������)m޼���V��F�S���X��1�8��]�6T"�s�����[wvm�֖<ό}Z�H+�yׂ`������*^��2��u$y��s�k���۵i�x�LS�>��O[�5�e�}]o�ڱBd�޾�s)t��ڽ�K<n�0�3T���H�3�9@���R��׽�I���R�i�N��ɪ��Տ�����a"�C�,73���5���̚�SWh
Ī��>��ıۺ�r�r�F�����NT@� �C�e<�4��0������_���xZ�{G���27<�v�[�M�*��D#���:[�۴�)���wFrg��ݞ�[�ڢҰf[�z>��}2��a��YG�vi��s��TkE��q@�Vʑ�Fv�\�M,�zuT��Jێ��3j>{��Z��d���";�;���J����w�]��:�7GVV-�38%��}1�zI���ٍS˨U��4��KFv�Z�'v�<�i!�g�vJ�/�GT���os�@N2`�	޲$��7���N�;�.�4�%f�;�<�s����V˱x�%X�~�[�Yzzo7.n]u]��Hc�}���b�Qީf���PY��Rs�w��VU�(����6]��B�j����9�2����R5���'u����OT�dj��X�H�$o,;��82+M%���U�1�<O�Ŏ�2�w��O(m��f�Vv�bA�7�i'�v�])��sI,!v�h�����1���I�Ŋ�ۙ���9�=��U�&m)�Ͽ�d�ʤ����+��"[av�YC�JF�1��֑}�������n��;�~����q��bDT!�~�|�Y36�(W��W�Y[C�V�>�E�Չ��X䮄1HD.�]��Lu��TN��V=�+N��	s�3x�E��ʮ1:*�8&�^�QKk."�CavrI��W�9���V�^\��9
����_)���D�^v��Z�3ntL���z#���DG�mR�LD�==�j{$d��F�S�[Ԥ�FѤ�L?o���U����q}��Ft߅��$R��c�T��n��na��̍t,��VL�,z�ASG����D�>�[�Ϸ�/�RҼ^;H�E��j���P�Y����TE� �
��B�3�ӑg!���'{v��;��º�1ͼ����}�]}�fe�f�'�U���lYQih1���H�EQ	����`�J,d�2J0����AH0�0�A�Ae�R��T�%B�E�a��^�{��n�i���m� ���*�`v�z՗�i×YiAs1�r=:TW�ݾ�Q�����Ѽ��6\�s�nC���%uc"z2g��ԓٲ}ױ;�ƕ��}7�
��y�\A���v��pּ�����)�*2E:F2K�7=�y#�Ξ�N6�1�Jd0���T7�b\ð�S��y��p�NE�[3^�� n�!�F3���*��YJK�����$tNH/�sf� .�N�y�R0vO���%D���)��2!�0��^-+���}3�+
������J�e�#N5���y������J\z�C�9��b��xK.ϰ����w�L��G��i��jQ+w�X�ns.�.��ޛy��"�Z�:�șWpn-�j�r� 3��_f�u2���InP�zӬ��oF�Az��{��7�7�<R H}V���L���7*�ً��qݺ��Mv�1�Xt��{Й�j�)l��k��{��G,���3��捛N^D����f��Α���[��lw!�g]\���n�'6����P�/Ev]Jrw��L���݁��W���X�\�+Ʒ�����/�9�rup?Ojj��Z�cJ�{y�ZlE���W]�Û���G�"��6�lP�Yʽ�r�^7�*ߣ5��Rꍺ��ǷX��7�N�J�.�Ć��IU��]44nB!��)��;�T=�{\	Jw��-�Q���j�a���{:�>"�����Փ�W�`;�L�9�Q�w��� q�k
8�W�|_p]o>B�컂.�SؗW�>=��~���Q��
�2,��(�*��k��÷��u�U:~N�H�R�u�<尞tiЈ
�Q��FT��}/��9üQ��5�CM`���D�;i�ܶ��H=0�*J��p'��e�-Wyh��Z]^�c��ۣ.-���?C��A�(Q d��<�I��R 5Hy����i��jH�hb[(P=�Z�G�j�D���z�v��3��a!�q*}�MK����T��N�u�O��Jﺦ�o{�ϖS�{A��>�������D����~����h�'��2;�so�ͬ�j����ܔ�}<x�ㅫ��C|��>� ~�<r>��1����>3��3��p��݌xV�^Q��i�ʫ��wy.�� ��[�k�o`� �~�	�����\��>V��ݎ
/G���Ρ�˨'|� 7:��u��oyew{�2�dX{M����8�&YQ���L������}�.��}��I�un�Ee�R��-e�/ta�:�`��3S�J�����Pz��Zj�D�#;�y�Ļt{ 3ɬ���Y�*O�ʾ��/h�SMҩ��6���gt�������(YfT_a�G�=Z��P=�]ٵK4���AJ(h�w1ĐW�F1O&��8�±�T�'��o���xβ���7ަ���Մ;��jCsaD����>��VK���YJ���D���N�A�r'7_\򣊾�9��#�r�Sk���-��5�U;a�y�Hm��d���Ę����=��Z����˰��;εh=��+�0�1�o��^�T�̌�r��v�å�禩��i���D�fcޙ�� ��V@_J��dT}@P U@P{7�3��2U�t_��mi�ز��h����-��q��2U�m�4��fu��7�Ѓ��6��:�Y�R7�ۻ�­͊Tz�*�j���"/
��u�@nM�bu=z�@�|S+m�WZ��\�f�Q�P"�0�q�S�)��.�8ԗ޻\vSe�m���zu��sAX���t�`	-����绪vhP·�ЃYޕ
=����z"<�Y9��^N��х�$�E�5O{#�����o'M��7�=Ko~�˦u��L��������Āf2�d��_�υﻅes֧���'�1z�ڐپy��%����,�}Tq{�B#pG��{;^��ԤP[=!�)��-k=�̴^�*%f�8�D�z��j���Ȯ�}�/���oUo���<��&"f&&St<�hS���h�7W����i���}D���:*/�*`��:�޹X��"��8�wS����{c��ըԲǫ��R�<]�� �*5�c�9�J ^��"ӽY��њoy4����g����9�z#B_Ful�aj`��6&/�UZUsC3BM�O�ͣF�c����=�S��P�M;�G��R�W��	h��3֫�w��x���w�y	�-zy_<~�*\�kj)�4:c@FA,�X�A����hWrB.un���#��`j��K:�\�9:	%͊�㏲�
���T�=Y���?�<8�n��OA���x�2t��Q`��o��z����P�]��h���x('����V_�=�:|@�J�G,7��R�=�=���3.C�G��}`��1R���A+���	$XH,�%E""���C�B�=���I�}Pp���}�lc�	�+�5uJ�ƈ
]�*�uU�EO��.3U��&E���![w��(JB��B���Uw��V=�h.�W<F!���Y6W�i������3>�JJy;��)t>��n�0SԞ5���G�ޅ%m4v�:u�(ۤ��lN���*2��/�ȗ�Kox�p�g���;��a�q{*[�=���"�}��{�f!�������zYykfqF���d�PΖ��R!Z΋WG�=P�-�O�����{����V=7H�UYZ:�h�~HU7�W�q�0���h9W�yt%��4�w -�|�ob���rH�K:1՘�s;=��|�k�jw��;�{��I��� E�UU��[m�Q����X�P ��"��QBh)(�+(6�D-��ib�(���H���������J�"˞m��W=�=���;�m��������:�]�М�w���Kn_FWh	6H;|{J��K�y�������D�.}�3;���Z�r�0?���+��@xV�����������}��y�+b�e�p���{_=u���b�`�sJ����W�%�=����	�:͈�g;��鷑�+�x��ҲB
�S��}�QÂ�;�k_L���ԕ���\ٌ7�D<<�zy��r���r���B���<w�v/����H��M�g�ۤף���Z��gy��ڸ"U���ǑK�9Ϊ��8�t��Qy�AL�[g�<̈�����ߢ���{�*[u��:D�S�*g���{&�R�����.nCY*�eP��Wa\$�lp]�[��Ͼ�\���(, K��9�����<w�@���N�7]�����l��u�㙼 �$f\���) �r�����c(
��|�n&�Ncٷqb��'�f�K6l,�QxWuY�8b�?KJ6�UU���ُ7���-ټ���7�{�*�x1��f�pᮆ�p9;}A��)�A*������U_��r^Pw5����z��.�(�{}Y���/d����}�%��͢��e6D��~�c���&��dtc7�f�=�F*��9�7}B�g�cTtv�(ռ��Q��C8ӣ��M�.��9�A���+���}���N��S���Pʚlie�
�C��	۰��_��&z�jj���Sނ����T����<�Բp舏e�f���&tV!�;�ڷ)ʸt�@�Bc�}�1/K�:���-g��X�h|� A�V*a�[�i�/^�&�w��ڷ�mB��VW,�p]��苫����p�|m\�|�I�9�6����>�T��x~����$�(���yޛu�6P���%����f�p�UF�E�5()+eں��E��!�P(|�tDt�K/u��jZl��sF�N��f3`�A���*cA���*�dut;̩�[��Gw�P�����  �B雇��s��gH��q�]��(+[�b�����zm@��JCHEF-:���� '��=���͸�5���F�����PF����fY�Shtp�]y���+��Ix�B�i�B���	�ZJ]cpT��v/E��a����}�w6`�h6�pJ���<lV)��L2=�����a�v��iegS���u$R-�s]�9�/3N1������g�u�����8K������Y�5h��[@�i�u�0��:Զ,Ɖ#�l_l	�f��iGR��[MeO��H(�ܠ��8��Jb�ud�
�GK�Q�#.m����`+�ªI K�Ն��pN�;2�^nk0'�Mo{��@��]M�AQ+�\Fk�C�N5���VL�q��me�_!�RpE7�ni�V�v�@D�ƒ��� �����k��aN������ j��l9�;3��X<�mT�{)��U�K�����I���d\�����+m�&���d�6���PM^䬽�R�m�}�o�Xn�ce�t%G�Z6�,f`��UB>JLK2�M]����̮���چu�B=�w5�+�wv��룛Pl|���{|Z�M��T�;�
���=PV�N���A��]�XPĳ#A�oAy��X����ӕL�W�tKR�VX�b�J�3��7+�)���]��G��n���z�ʷ�4�y�%���nscUW�.��ѓ���FV���G�~@�֭� ��,�5�&W-C�y�s�ҭѽ��
�[��Dv��ϰ�wEZrZ&�r�:�`٪Iؔ�,�]
�23I<�F��U5��.yO���[=�j��L�4�̛OWh����Y�s�q�}7Lq���_U����沮�ĝJ`\��� �S��'%��Sk^*i���B�p��	j\�)��X��=n�s,Q�܈M;������-D���:���4�l��o��)���������ۺ[���o�+6�{q�m��Cx�n�t�v�!s^	��Ҩy�Ö���ش�:����s�ʆ�6�KZ�[Gv�
���-_.���t�:��t��O9�A�[N�Y���3�[�M��P�)�*FY�U�SB��M���Ѣi.}�Ӌ[wU˜n[V�n�T����9Ȇ4Q��K�izļoм��7�w��Y�˺��[8\���K`�X�7W�WA$7�^�>��w#��`�8=��x�����X�;��"<kZ:��z7��Wt�(5(Z��z��SM�b|c9�ns��C���2��J�R�I8���5�흁*ciL��U23!�vQa �>\�8��}��
�6�)VlDGE��*z�0���N��[�T�X�zߨ �Y��ʝ55vh���nO)�w҆?)]�Q�'�	�*���|�53���^��a�S||��პ�> W}��!ϨF ��MJCՍ}Iud�n�y�LQWbU�b9ڕ]dgkͻ�P���(�^u��^�tU��B
9"��ϋ��z�k`B��k)�mh�W�{�JZL3�l~��.�P}�\�^G6}��
���5T�O�)Q8_�g��V��^n�	�ڔ�)|��t��NG��kM^�5ͱz���#{���͌l���+o ����ݽ���گ��@Ȕ�z-�Z�ُ�͘ĺ��<ju���;�j{�YqM4E�Mgla�y|�c�V�C܅����O�>��a~�'�o/{�e7�����I��������Ӽ:5��r3�[s��t���|�H���Rv=r��tE;b���P .4�g�wܖ���(�#qd)�n`m]�"�BY�)>��WY��3 �ꞤR�Y�Ufp�U���@���_��#T�]��5��ǽ�x|~΅��KPcޏ��p��[xw��R7j�;�������Z��l�}\�+�I��snm��r8����YUX�#�������i�ɆY��.�{�kU���b��kKbVE�5����Q,ͼ�TS0��(@��w�O4_�C�9;��GV� ��lu�� � !(ġ���.�/etJ�Z����sSސN�}O�=�ZY��$;��� v�&,I���ڎ�ȱ�q�Y�}W
�\{�X'�^j�r��U���j��YMnL�o�m�9W ϣo���Lod��q��j�O;����fc��D	���y��=�W[�zB�
@	O�������7�J&�tg
��s:�ko���C{z.�nK�y�'q����.Bۺ�����np�*�j�`��K.�I�%z����壒�B����A\��/~�w��q�ߵ��@Y*2 �"!�X�� �H��
��H�ƶw)(��8�C��en�Ub�v��2���A�Xk�C�"~��x�5̞�J.Lڴ�a�L�Afuu]��u�	�IU��gk��Fa��	/"x�sS�Gn�W���Y4�v!r��@�S�E
��
��W���Q�%Pv��nMC�D���z*��lM+�<'�\�,�C7�z)�߼����ب�
����r`7���9Il�za��*�7mt���ێ�q�$[]1�9GLa��z��x����
��2��7�P/�Q�J�,󬀻"��z�B̫i]Q��ute�{�NP��|�G/����Z��8A��B�fu}���o����֕�s�u'��Fr�}�yl�k���[ʊ�v'T�����k�kɓ�g\έ�y�0�j���5�TK�B��y)�ù����x�ds=�.�o��y����'$RE�A���  H��^ٗ�Pwt�R�ήB�
�IzG�a�������[�J�N���Udfr�`��4/���y/Ec�q�̅NN��j_\��7���U�� ��3x�x�xh��ԧW�
T}�<�;"N�>��x\1��w���2%���U�>��6�pes�Y�6�n�7U7�f����?_�����N��M�������o$lvʞ�*:S.��<ʦ�n��T]�Ov��}�����j�(��c8��m��Ӏfu޺JU�WX�S��Z�]�V�S�ΙrM;y��l�xH��E�y��ǽ����Ej���E<���]U�'6�5�In=A��Qr��=��iۭ����r�n{>p�j�!C�-���9p���c���[n.�����ҊI��p�VF�*ӽ�V_uvSy�r�.�:�Q���`����ǽdɀ��LJ��^��ZX�﹌R��w#�3�N{��I���ko�X��ӫy��1�z��n���D.6�Bn�����p��L��\k�w�[4�v+� ��x:ӜK������sn'ڼ
2���3�
5�u1�+�p��KGL��TP��.������U}��Qd��V:}�D'�^Um,��:�9H�A�Z�������Y�ٙY%	��O�15�k��t�QT��yJ+����upY��(�B��
q(�v��V�r��Q-L={1S�C�8���z/�V�R"��T���M�eʧ�G�3E�_y��AE ��,��Z f���;ۭ��n�fK�O�Ի<X�������W\BŽ=�M�nԫ�B�VT�4�ur��Ѹl�P��z�{+r�xw|hxq�����'��j݋�+�������x>,p�;:/�mo�e�n[�j�B�k&.�CC�ei؈���hׯ�u�DG����a%�bmR������� �r&�woT'��\l����f!�g��dz����s�5H�]��tm�Yή��1�h�OVX��'����e���#P�^�i��U�����F��y��z-va���Q����{�R��[ƪ3p\v�w�.z����qt��kg����¯�eg]n[z\�Q1/K��ѳ^"1=}K8��F�/(��g�.������H��*�p�/ٽ}11$_�X��%eT"�E�0�Eb "��ETX���n-�fHIoj�L�(t:�ԡ_R�4���n^�!I�-����4�1�R��p'��s�:aT�b�zF\�<y�ސfw9en�"_�T�÷7��KB����Ǘ�m��W8�=Є�V�(���S�z�)�ZqK���.՞�V�ܛ4U2N��t�L:��	�L5hV'���9��l갧�^�_�п`߾ �̡��Erc��of��0Qɘ��P�(��e����̛K�}��fG���{�|G�����u
8���Ļ$V��FQ�3��;ʄ'92��56UD���6Cе&Oh���k��JV�y���:�WX��,'{���1��&��m���(�}���A��0أz�Mk7�q�(��3��	�כ^}y�]|{߷��>{�!�D�HE� 	�ý�.��%~m謮RoGU�p��0V�H9N�(h��U4�he��W����RbҐ:�I����6�eЪaNi1¯y&l���f�Y�z��=9���J���&�Wz�Ӗ$����x�٫��xN����ㅟ:�x����.ӎ�}c�ѝ}�`T�p��n�fZ
R;4o����U��iq���l�1�B���s���gF�8T�3w����q���i�~�&�so)M�D{�Yh�yKhl\�K��ns��;ٽ��um��q���Ĺ���qO3�R��:�x4�l{(H�G:��z�w:�����.6��w	{�xZK�u�c"�v�^�G����mr� H�@X�AI���-��u;��k}{��u�z��띱E�ԋ� ���B�G9X��(�$T����0�Q�
dE�b����maZ�UPUb
)"V��F�XDV�-�*
@��`�H��|�?/���	&�OZ��1�(n*�y�*��Q�pu�մ�3������]�����;gg+�6۩�n*�gr����m�cS��ՠ��z+b�.f�u�e�M:HJ��Z��o��7p���휉I��ڋ}ӝJ�+�fׯ%0jbb�ر��N�>|����鷫�;m<ݹ�vu*p��DI��1�hQ-�q�"<��>�0�Ν"���lIQ�;�J�e�r�6� �	�d�	�/�]s��U6#c����b�jmP����"uͱ����۸�  >�7����9ۍ��l�8j��-I.]�ٝ.g�Z���tw��s�2�r��s*�|&$!G!��P�H9�%��n���j쵗U9�Y���������V��h��w۽�
�
��**����R_(Tk2v�V�"��ebh*�JUP'��?��Z>b"�P(���>>u����x��S��������[��gh� ����:��A]l**�{�G ��z���**��?�����;>Ϯ��t2�bNB����EAs!PQ �
���`�b�vawwn-��邨 �Ï)���GCB����7�AYl3]�m̾ ]����=2@Dc-�R����c]���
v�	�8�}$P��H�E �APAWq����s����;?Z���HTUǗ��� ���RԈ-�Rȸ�V��\����TU��.�@cNϞ=��߆J���eu��Z��������ρ�1AY&SY�&} �P_�`P��  � 7'�`b �<��j�|	'C�R�`-k ) t� ��ºh�1( �i݀���4  �
�@h��)+[F��5J����٭AEJ
TJARf��LD��*U)J
�UYj�k
��4�*TT�CR�e�1�	!UEKkQJ��P  �U��m���٭L�&+1�������!EK��`   h P@�Pz
=v��P Z(zWN�	�/z���e�t���wNZ�6��.ݝҕ���Z�����9׬��wwzw�{:r�c�.�{�h�ɫ[z�Y��޷gsˤZ<��[;c=�o2�����v��t�����vj�֢�{n��(P��(=����h/zY�y�^�A� �K�w�U@��^5��n̍�6N(��8 tWv3y�� -�:k�h4��zj�s��jt�犉����� ����[ӹ�`47v� =����� R�^���5�(u��E
koZ�v:Ѫ��;���hg.�9( ;Z� p�1jE�*s�l�h0<�P�����

:s�Φ��h���ᢀkL�g��J�
PNyu��kA�9�i��t6e�eQ�c%�h�`�w�֧eB5lbU���l;���Z��Cq;��H([�r�h�	�o�
5�� hk[Q�V�9θT6���@�e��;z�v�D��A�RW�Ƶ�SXf��6���Y[ ���)�:]��y�m��3��
=: �c�դ�Ś���Q�q�T�vj�Jtvݷ]7C�4��W�(����� �E*���t4D�t�D:��;)�Q�Y�lu(l�-��=gF$wlc��R���s�QѕSYm肊�n��R����B��X �N���
魑[F�Fv��EU�R��y�wg���%w\9TO=����j��$T$K��mP*���R�,���k-�)X�A�w8� TMA�LEg�9lP3�7h�zw� �v���m6��D6� �yB�᮳�Ct��]��uK�T��h��c@�wV��g(�k���B�3Z֨[��DB�`{��:�R��L)EQ*Phm�	�n S��J�h   "��I)U   j��3B4FOBi�d�"��	IU@� 5<&�JU4�`����I��$�@   w�_���'�����g>��!�Fy���v��9f���5�^����>�v�(t�e�o}CxB"��{���CL������CX����P�[x�x�|��+�Y�o�f�ۃׄ=&��[���Y,�B��F�����5ɽ��3Y9��t��}��/��B�t���F�l Ǆ��"���K��b��T�4;h�ve&��^(;:q�V��ɍ�F����4���^	�rnqd�+5���գ�F�oR�rFU)D!Jgy��ּv�}Aνل��m����bR�K���K�Trk�fT���-�SJ�Y��z��Ђr����J�w�8�l!o�A 밖�!^�K,�!�q�#��<�R�Ѷe�{�]ЋA
�F�ڎ];/Z#�٨f���k���FL[12�K���jw)|�fȋ�4��`p�uY�hî�x�lLj�Cf6m�4�ˏ9�\@�ۜ��oLS[át�ۙ1ꈀ����N��-=����FDD׸{33xf����Cy���v���i�]�ю�a��v�ү]��sqo#V�O{^���V��ɴ7K×yE`�4�u������kbG:�k<ͲE�kkO���=�c *���`��(��@P2H�$TX��1`�
���@Y<��Ȫ(��b�S���WZڲf�ݜN<<�_*]YJ���E" Ā�1R(���]P�xp�]�:.�xe�����;w��}��+��f�|�o[�4�!�C���h���J�n�,�*��C�*.�+�7}�Nemջë��K�sOkrgfA:�A�Ǆ��fZrQ�և7�k��5䦛���Nh��d�����)�n���F���;9��L&��	��#D#Ňf��T�W�U��pŇ�!�H�R��8�pt�6*Zs�(�a*E��hz�eл�����0F�n�l��(D��$�~�{{�	ET$���g7��a�k�vMɱ�[9���B�|p� �I�FBP� *2��y�����ØZ]^g,��!����W�c�l�fN�[]0�
��m�lٛa�@Hi�<�Yۉ|o����f�K�Q����t!n�@�rGp���3	���{�Մ۽`�Rח�sσ8eMwv��S�î�����4�����U�%K�V���x�Y�Nv���ˀ���#�:W�3��"�H0H�E��6���l�,�������*@�hV((�)D�A�M0�1��b�3Bs�YCh
�:��j�-@X���*� (�*M2x�	�b�� �T���߷�1!^�( �|��+64����\�n�G��ѵbK��I�<�@�У	R)
��@ů���7�.�+p�w&���s �{^��I����E���I��Qqf=�K2m囑�����:n=�I5��}M�gmgq��k�o1�q�y�י;���]����|�6d;�-���P5�l���&= �5��w�����#�>1o!q�c���ُn0���_�͕,���u#��ᅽ|pJ�w�'^���ŝ��t��Ɔ��f�����ŵ��0�ݾ �����+��Q,G����������e|��ǉ'���#^wf��VY���A�V�RL"��F��K��^咍��ܒNa|�-^�ץZ�+X����n��8i����'=�4iOz\ȩؘI�� xB ����p^Յ���e'�u�CHC;�q#�]m��}w�d�ܙ%lh��㛶uB�ƫY�$�w�4�g��nv�3�����7N�KY������ Sgsh�o��O�*+C�D_�8�tbph&�9���A�&`�Ӵ��й� ��nf��Ǉ^;�����ٱR�aZ��NE���8��X����1fe�S�������{����a�[&�Z�l/�@I�F̸�b��w)��lΒv��h�A9}��3W.�=��X�Lǭ�ǃ�d���a��I�;� �F<��6�QAAb�TH��H��. �ɽ��qd���fR�R�#k�)2wn]���\�=��J���@X��V'�
�QH���#ԣ'��}�|<M#ٰ��ô�r׎N��6��&�<��\��b�k3���e@9�>�!,g�7��}�D:�z榭{b֡L=��K4�
�
Ql�:{Dᗱ֮odТ�e�&@�Bv����3^�.ۯ�V�Q͗P�
�<ӭ�Ŵu��[rd���J��G�h�ƭ�o��n�#�UM�rc���0��l靣��}7��ۂL�0�Xc�B��*f���/w^8p!SǕ	f ���^��Z�X�ه��<�]��#ssq{���MW���rS�E��T�����K�n��û�NL=����Zw.Ґl5��06s���M�f��UC�=`c!��,��j�
���N�*�"�a�QU��BV��n�]F�����Q(Jy&����F*�7{�I2컶���K;�{9���X�����.��B�j��MY#��n^׮���oSy�,�׵���[�Wfc�D�;��Ú�Y�bm�ZD;�*ͬ��N�r�,-��9�:���.o�;
R{r60%�t,q���[��$ �/�u2�&!�9�"��>�S�9R���R�/8ǧMK_o�vխ�H\-d�(�e�ɴ4��m�h��^��4�]�x�3�zǮnp��=5�����Y�i�Ʈ�0w�3S�e�Cӻ���ggQ���J����sǯ�7��m�L���B:�F���������I��Bu�����XT�N��<Ռ�Q0U����e���f�XT�IDU#-�D�Q'X�XUx��R�'��"�
�VA��8ʇ� #�q�1�tf�,�]uH.ك3qkE�"��`�ɦ<joh�Ŕ�7T�~6E'<!��3�B˼�}�#� Ci�Ԡ�D�U�V� �4��O �ɭ�5�W��F��r�A���JH�sr���	�u9�k�c
�y�A`cCV.R��Hc�L�� �E@�u�q��!�V3��^�IhX�.�TaR��A�F.� �2�Y�����
"�X�����2X��X��P���Vf���p�"�ٞ��,�L#�l��nb�ϖ�[Չ����&s`�:������{����	w5f���&R�{
;����0��B�Z��;�\,�7�@��  ���x" �#�Aͭ#"���\�Gac��R{�-�����K�/��ç�:-�f��+��UD�����ƽr��)��H���#��Yۈa�yr���d�z���X��K���ii
��M*��`�+�0t�!R[ώ�vܥi�Icdl݈h�J%� )��j��n8ݗg�>����}.0�H�ay�z'6w"�`�̽˺9����L���=�l�-���pvTb-��������eg��m�^��	�v�w�����n�^�N��1��#�A/bޤ�������ݥ��8<UM>�0��q���E@Eq~;�Z��M���Z�����T��3PĐ�ss"Ёi��5*�2�1<�9����x57{�о����O>��r��郴��sr��\�p���$���p��սo�%ii���hL����tf�x�!����
�SIb)��ۏB�73�`�l4P��^�u�^ڴ&�͖I�[�7z���$���d���xj��q���0BUm\��v�Y]��2��E����9݃x�gM>�i���[����r��^�0��mn�a��/3no&��� �M;�+m�d�!�6����%�Wm�H���\�)Y�V6�t�U��;$F��&6A�[��N����Ә��Rv�qc����Σ���LE2l3�	�%A�]K֩��K���:#���':.CлM�2��BRc�;�]k��u[ʎ���.$p$���1�"AbȈ-"&�b)��M QFAUb�Q����0FH�PFi�Q!�a8�T�� �ӹ�x��X01$�E��Cd�&�z����q [6xR%a�\���S�s�.�,kvQ0쇰��j�a���z29sw��9�痘|����2XB�FE� �A�mYE� )��ł1dRG�z�BR��٢	H9�yq�4^�r�`��h$"�ܝ�Į8�T�"�ufE��0k��Y�ȑі�Plx���[�|y���pd�D¡�&�J��q�:�DP'ԥ�
��e�б��U�[j�;O��zV�qMƌ����W2輷0�6k��FPx�Mg�0���c�{N��Z:L�a:�
�,F*o����5�y���d<�;{����c�lxԝ]���+w�t��'�\��Kǋv@|�S:���N�{�G.��=����1Y��Ŷ����"�	crL8i#�b��0�]�v�:��[ۻwr
�'$���8�EC3qk(P��TF�q7m�>ۣ@!�)�ȸ��^95�Zz"J�����+�_gP��ͦ�;;=s��	ݘ����oH�IN6w��P�1N�S��b"�4�����������`�D�l�1���[�%�gi!�p��܎HFxI4�A ��[;��m��=�Kځ
�g��R믢�rAvm��{KP哬���8A>��L������j47�ሲ�l�s����HaN&td/l���(�õ�UЦ2	6�M�S2D068��=�{8vH,�5�sT8n��.L�5h��y<��5��P��1���e�)���9��ǌ�n�eo���w�,M��?/�A���=��%4n%�i�յ��tK}�ս�Of�`��؅���J��$�ӳ'�&/L`�s�c��m�fb޻�j�!�ˢhҨ����16"�q �by�zE��=;��N�����R�@W�7��S��R�I�m9��v�]A��\%��%嚤���;�3z�k٫��`��X} ic���0A���}d��BK|�|�v���`�swH�<����������znYf��'5�cuʞTU�����+1f� ��2k����@]�F�h/DQ؍�x�=V�۝F��k���d\k垧{� U�r�١*V����w*��n�>���E���]��������7*9�:a�E��:�,\�>����b�/	��=U�a���� �Df��,"��'ft������%���rt�[��hJK0k��;z�8��.n5b��P�ʨ��͚|��˸Uʗ4�z��`M	�!q����T�����J��f]������}��'r[��k7��U�d�{�3��6r��`�z�W3`��b�����]�(�;��k�͈�>1n�+�ꑛ�_N��i݇rq5zB΅8^���	�<�u٘)،�Jǂ��f�a�f	#�����C��5%�жT�Ѝ[.W�=��l�
��Mˋs2�6�.��pzx���]ЈN̬�G;�8z�Ջ'6p�SN�\��&�1�!�)�`ص�U��xg��7�����0m��;�&0]i�!Z��04�4`w�^�0L���i��zs��e��ic��8C&�Q&���;P�wZ�Xt��/*�`ݑf	hd�3��Bb����x��x^6�v��ڴ����jp�R�y�6��=�tAk���S81�p��V �c�D��,�ۺP�a1G3��ɚ��j���Ɔ��d���M7L�9̖*}��B AD��#35jHdl��g;����ó]�^y�ĭ���y���P����� U��;�c��zB���݃�S�'��Q>{R�
�ӽ�g�����6��$7L
�u��N�o�*�������7AE��/]Ct�Sz۰t�V9�R}oi��B�<p�����*����O�N�n��W��h��rO�]�&��3��=�߆�Վ�*#ܠ�M��1ׂ��e��fK�:E\0~Y�a޵�X�4:����=��+���B����`P��̥c�S�s��oeҤ�z�p�+K�Q��oCR�NnwXϘ�*��c��if�i����|k�C��If�P��z���PM����V����m���9H�����%�~�{��а�`۶��U,�oCK�[�䊱��Qm��F$7�JX�=�Kz�dw���*o��F2+c�!A}<w9������ޮE��9�J�/r&�]��.3,�](��]���Εm©������G���8�2QG�+F�d�t�b�v��*�5��yG]����h
��}J0r����`�z8��,���K�ֺ��*�},Ie�L4�Q���qˠ���r���=�cxlu��Nh!�w�;Of���]1���l�y�f�����w���+���������;iG�Ј�Ŝ��Yη��Pf��M���f�A^Xm��UCv`��x8جY\�/(�4lV�{}X� �e�% �������7�m�>�j�'��[����E�L6/�(p�p�n��yde�tY��ם�`p�8LV�V�f�3:�M�e���Ȗ|��NrV�<so����q����Ε�*s"�_'N�ime�֥0��9�wWV�%,���P��b� �6��J�ُ�[�����Ď���P�q������p;ޫpއMJ��!Ly]�d���ۖŕь�\�f����ݡ}j����0xM�1G�0����뺴�|+h��݊��t��O�uy7'eˎZx�,���D�n�#HB��҆<�}�@��o/IF����Gn�7�3*��j�2%�^�e�F� :����]��蚫���`���3V���
CH&�,wWn�}�]sΆ�)}��ͷ��Ҙ������v(�b�1�%����n4���� Z�`����i��\��U������U(//�tPG7Wuh*'L:G޽}-Y�F�x�A�Ǻ֮�tQ�v�p�wH�E�X�7ho��c
\!��|�9n>�J�j�ŭy��B:��Wη�'�F�������ͻ�1�f�#䓴���ܮ����[6�s�<u ������K֤� �6:y��ݷݖ#��[�8:嫭�,�<�1�'�+���`��D�S�u"�Y��GW�sultv�o��N�b{��t���Vw�J�	��C���_�p��[ۂ?���Ht ��V�T�����a��@5=�㶈�7}����Av�4x� ]�����6٠�>z���$�U��ע�x7պWw1�XpU��d���[��.D:
�Oves�a��\�޳�l�uN���Y5�������E�/3��MWR�YC��o^�m�"��D{J=��wF	
��x�_]u��v@z��
��9.Q��}t�P8�v�d��3�d�2�o
���\`@vn�M۷��\R����S�\Gm�r�Y�h�]�F��ŚZ���3��Ηmf�[!7�%�y���R3)&Z���� �&��~��,�E�r�����v�hYʛ����%��vqWI�+�rtY�wA��AV�p`�v'����<4;�X�n��+�uK5�,�M<b�}�{$�SA�]�ڄL)d
ݤ3x�[��tT��<Gn]Jt�:���]g�t4=����e�H�;�~�;u7# C��1��7n���R�|i�K��&��5�*I{N���K9z�j��� �Τ�x;$۵Ea��%G��2��ORzkl��X�J	8�K��XJln�J���p����j�W�F9�V��TVi�Za�N\�;��az���,�R�[���,�&v9�Z��3��ʋJ*���S�[�	W�SHv���MY��/;��b��E9�Y�:�����f-gb�����HL�X*n܂�S�4�h�nweB�A֛?
�j���m+��W,v2 ��b,+="�5�E���ސ�Ž�&�fu�*���׻���y��:;�� �k/:�I�au��'5�F�v�;���j�7��2���-�3���m��c��W/��R��x֜��P��]m��<������T��ݭG]��[��Cs��E����|�uE�]l�6��Hgd]�F�]���CGJ�s:�.�[�U�*����X2Bo,��Kq�1�6U��cX��3��7���͙�� �}�m)�+/�z����`�@�ש���9W�r��Ft��s4��;e�����ٔ�G�S]��Iy�훜gila�o����&g!��]>nYG�)�6Jځ����4#ϙ4��r�b�<.G�������>��'�\���-�2�}0m�_�̱t݂�¾ԃ�3G�`֦vpUL�-v��m��Mq����ء֚�!�G�:��j� ���,'O�p���76org�`�+H�M�ˣ�@F�-yܱut�cZs�8�&3NSCn&�rP����b��v�B�s��6�|�<���*"�nb<�a$���/���z�e*���k�����w�7��J�d�II�,��\3G0���]��]w�=�u��Q���3q���\�u����vwe��j�4�qe���P��$���ܸ�=G���O�)�5�R�ʦ����{��_e��1�Q{՛����\�1��Q���)}[�Kͽ�/�]�Lu�w1�;;ȅ�����]��8�	\I)��ʋFU����z��O���j�m���q��3A쌌q6I�m٬��9(ݲS�i�˅���Dv�R��Ȅw�WgT`پ<�W9x�M̐GBв�괖��\Xv@��`�y�h�r7�u��i}���vY��\�Xu�;y�aű	��;/kiu�������9-Δ&�%`���p^�k��V��*���3���u݌�K�9��_k8��� (�0�-�P�lR�V�m�:M�Բ��/�����\��{�^ݜ� ٽJ%����q����N��7Yz��4OPVvO��b����1j��sfV��p'���+Z�th�qu�̵���ٛ|��3t���B1�N:�a��W�(����M��.�C]�*���k^0�~
�mq{t�,���A�!�q�v���̋�]��|
��:�]�
�(�@VSv8uĶF��/*�C�����/zVu�Waoh��.�z���S-en�e־{��2У|�vb�+�p�r'3C���f��i���\ꙅ���D!��p��қV$+[q)"³��`�h�X�V�X-�JJ\�֮H:�X�gI�V���Ҝ,������j��	� W,韶�b�]�f�)Prt�ܻ�& ����K����X��䝳Yj�e!R�γ��mv63�d�6RڗO�[��VE�@���R@U��fu�.�2!�;��B�u�:-��&à�o�jkm�yv1T�3����I}��p���hp9�����ga�:{K2���r��kI�(�������<�j˜�l�*�#���p���w¦�J�H�-���Oe�	�y�Ѩ�Q��]�0N:1ʮ�k)ȫ��
����:�/Yw���A�����`g����0�xX���������+���#��+]�����P|�k�P��3��ثc���3���c�p�Xl10�,���gu�����s��i=�}V�	]:W���v��Jݮ)����� ��Ig��;�c�'��Ҁoe�/���A3F������>��pZȚ������f��jV��c9T�ՑK�/7��"D�����Z�ܺMO���]u����tc���Ϟ�x�Ԓ��X\Y�&�`�.������3�R���6��nq��xE�������y�NǲX��^5K2�uݔ��N��}-�(���ٝ��>�|�i�^�	f`��.�->���7|K���u��E� j��g�m�
�+[K�1�Vs۽Ӌ��J�kV�9prӵ��Y�R���L��\�N�^՝5����	,��E�*�gA�+���3O�:��]�27�fKν�0.�	���Q[�{��d�q����W����|8l
nڊ!��o u�(�+��&ޮgw�F�IH�Լ�`N��&^)YOB`<�9�Ɯgh;Sj�	V�~���c_�E5��]F�Jg��:\�[����Լ���ɉi|��Q��8ΩY���[2M�avk��G&��[T�u%�_���
��C<��U8�@��+����j����h�G]�轳��vʣ�՚$�����i���RB}Z�]��6�v
�V���3�[��'"��������0Z�	��V��zޡ�sX�`Z��������V�]҄w��֑(߰����/vT��m���n��}[�c�Y�oT8�[˖��@9�r�(�̂L4���2�]���������,��fi�T(�t\TBmg۪1�,�z��G�p��_65'��)7�y:�LJ��y0���#U��1�j�V�v�19�j�b�`vB�ڴl��oW<#0U��1�?�u�)e�e��S�g��D���R:m����R/&��s���������!�CVX��Jm�5&ۍ���^1J��V)�\&����K��n��[l�MK
���ѦTP�w 0�n���E��]NK�D����]oG������՝5#z��wD��}ƷU��)J+߭�pU� �!��D�vc���)�PŒ� :tʮ�{̎�hDP84��������f�\n��Q*s��[�/�{j�o�{C�t�Au�{J�"�Uz�A�G�JQ�+�<�uv��Ҿ�X��>�gmv��	�Rle�NֲAy����c���bkp	�>��x�<��6Q6xJ��_#i1}u�q�l|���loU�E�!忇�.f'� =욎]�%�����k�:�J��﹯���]����U�zFo�e�J��璄�&#d�-̜���Weg,]1Z����(@����^P�d��� ���ε��wH��r��:�q3�]�w[��L]0���T8�n=n=�|�u���i�n=��B������n��U��>��mIC�'�r	=���s�M*�����l%�3��8rRfeᾸ�L��sM�U��ܦR����[�V���ic�5�0�0�X��>X�60��qǶ�m
ė:���{Huj����y�����xk[j�)�΋�����Q�}�v�K܉^�7N+��;���;�;r��ˬ��<r�
�"�����(/�dΩ���r��I\Mw�1jI�F퉓�S���"��ҖR����B.��P��m��)ԋ��%vX��{�U� �ۦ�[��z�>�a�Z�w�k*�%��S�b���ty�;���N�Nfh-Z����J�.�@uf[������Kk�c�3G�]a����tۺ{0�Щ�ُ��Z*�M��*�!��F�t�u�*T�J����4nt�/F6c�p������պ"��Z窮v>r4������%m��˼�G`�]s~r|~gF
�g7'yV��H<Xv�X)E�%^n�o��Y[rP���X�}�b�g���[�(Gc6˩�j�K뱴$�D���!u�za�4'Ԩ�H��LW��k�ΧQo�V8\R�e��c� ۛ7��z[(Z�Ҁǵx[�c17�r���jeWH8
)�Lg�0��Ʈ�LXӏ"rǋ7�+�R�Hjް�t���WwAb
t@D��;kb2�������a���F+ ԗ�F�Z���Gܫ�LA�]z^��E��ƖM�������\̶�CO��E�Vt}132��&����c�-��h�v:�*1
��/]��?	���8 �����Xk#}S�[%2��,�L�v�&EwQǠ��}G�Up#&�R�u.5i�)��9���p1rP�vk7hξd�y��f-��kpvj��n��j��]nò�)X/��,cv��):}WQ�Շ"<��rn��J�ս�B���kQ��6XE��Ŋ$��T��(�ʑ�3�\�S�&�6���H�W�0��N�G�E����bx�5����x�JS1�n>ц�v�]�.�./)uej i�h�(�n��Cr�A}�m1ƥI2��
�D��䩽�TfM�����{R�0���ꇉb�g 9�p���>+S�`���@�=����,�y⒵����{j�m�V�2��&��yj�p�xQ�<N0�n�tT=��ot�ڴ,�����X֑��ݸ�:{I���]�AtB�NjI��2��	�D�3; }��˄_te #�4]X싩�7MbP�ϸ��L����b�U�!N&��ӗ������I/�J�#;i=����TF;�J��G��su�q��S������Kl|)�}�����U�y%H�^��o�{
j)vQt1���qB�ĸ�uàv]�Y�؅���9����y�b���-�$�K�P�AҎN��F��5BV	ڃ�%l$���8�M\��2Հ��a7?	\B�(��(�v"�����6M]4UZ�쟳FR�z�W����F-����Y�sT��\� �&��bӶ�=>Z�ec`lb���}�yp��ÄwS���k�Eӎ~X-K�5^���X�#�"B1=�r�ٵ��]�YI|ʸ��xf(��W��/P١�k��� ӷ��,���*_�}u�x��d���z����J��P*7'`\��u��\���}�Ы��A��G7&��厌�7���8LnT�'�Z�z4Ѻ/��f��5����9���7�	*�t&�.7cs�5�8.^>&�?g��C�@9e�AJ�ʒ���߉)݊+�(��* )M� ��	!R��C����T�*��v���G���M$BB[dy	$�$� @�$�H� 4����l�!l�I��;�O$�q�bB�w���$���	�n�BV�l�,:��B� b@:�@4�1�����d!8�%�`wVʐ�Ad+$�dL��$�4�$$�l�I5�2�I��"��d
�Đ�I%`k� c&�Bc$�m!P�HE��@]�|�h9@U�IP�f�l�vq��3VIX�X��O��T0`C��$P�h�V\�Hu�����1���XI!�Hm!���&�c�s��f�`�����m�$���!���C��$��繽��E��i/h@�<��d�$�������i�3���++1��I�3*�}���C��B�CL:�CH��`Lݙ�/�3�6�0�,� 4��Лz��L�%aY]'���P�������]}g��cY��$�Ę�I6ɤ��b��%�W-Ú��nԐ�{̴�_F~�i� <���7(|�7�8Ϗ����'}g���	䩗s1�L�`A����)��儗y�M3l��`fޢ$�r�v��B}i�����o�^&�ud�Gn�P�
cp��:�1��N��ՙkˡ�+����g�͠{8萹g2�`> 2!V~� {B��6�!0弲I�|��s��R��_$(���X���~�=Ấ�\�!�kHq4��\��7ۧ׸I�X|�{������ȡ'o7�sܰ1��	�g���I����z 8�ila�{���X��Z���+�[6��5�w�ӭ��:_���(/L��с*�/0� }���ZZFO{5L`�{ێ!�xs;thJ�{��)*�d�wA	Ľ� ��Y =�γU`C�����k ֮֞B|��hu��4G����}��i���=�9nq�rHMo�N��޵}��N�^@x���5����qd��1x >���Y���kM���}�bj�`xj���x ڶ?{�~��0��醽�$=����Ih�j}6X-�=�1�ԑ��!;�o몛<͹��=Y`s<'��?{�E�G�sv����A��@�ʟ�S��w!��=��I��K�X��e�=��G���ۿ�'�L#N`���b:�I��<��w� �1$7s�Uћ���lц��;����q�{!8��GJ�nWNW�ƚ�U'"���gf}��|���; |�W�IX}��өN7�l)σwt������������-��#����4杻�Xi��^�I�-4Ǘ��W�������s�x%� pzOO����=�x}+�����@`�Jwɓ�|��O0�Eve��*]{���L.��q]�D��� �_O{s�deaǹ�|��>�l����|���g=�<���v��O,i"��~�˕��+���]�f7���p��(���N��S�{ozU�8)>$�.) �櫟mk!}[����M?������v�ّ�廦z�p����5p�
�|���*��0B���BG�b#�wݻ�_��pA�#>��g �0P{7pn��yt� ��Z,:Ӣ��4%Ӹ�u�<���G?]�|ނ����ˈ����4��F�
K Qh��'�m�w
o�'�E5A�D��|��#-j���I���
�l�#�F�çN�b����(�{Z��F2Q'�+U�7:��&p_�=pj۔m]�u�4�xu�6�u4Ŏ����0)gY]F�P@���︝�Eš'��A�g`��9v���of�u�/�B�3y�G�P�]Xm�F��z�]��ӹ�MWf�����W��DӜd�n���=7NB� e�r��Aƈ�w��Yc)�>�	N:^�Qn�>#����3�Db)�,��ٔ;;E��u-+�fY�1��\*�<�����m�=�Q{�@҂�j���Y8��u�KK�+���c9TY-_[�ZB~��u"��sniڶş!���>p������o`�:�2�NV_>�f�}.�I�̜��W.)��)��TÏ+���'�:T �&D�.�L�Z�T�����)�)�M��r��'Z��U��h�l@��Sz��=�7q��)K*�n�Di�X9�����e�$�&�B�$n�8l�vm"qۘ���	�51��:�m<WM7뮜Z���2v����CO�����<�3g�VK$_���>9E��
DR��W��X[��F��M0�b^�x�:���T�m��F-ˇd4
?�*�Ӽ�E�U����6^���4�(K4�Ɩ�fC��1Uj�Q�	AܬǏ$U���ưV"���Pʇ`!�w�*e���'�V$�ar�����-®�%J")�����ȬD���}��[��m�Aa�� q��<�xOGeC����q��)������9���p;��b����[��	�1k������A4�:��rQ���sr�������rW�n�Y6/Fnb��X��d�b���"L���~� �@=A�����Omh:�
�Wr���h;��p q'9V�&�},�P,B�|5)ע���1���un�Zf��{���Eo%����=��cp��l膷������Ȗ�ì�.��*,����gS�FgQ���Ԡ��-^��5�4���r(�1K�.6*(TնXm��n�����f`23�٧�Q���gq��!2r�ꑺi�ŷ������EA�9��B�dgE�a`M0�H;\��|�����fk���7���� I$	>���|�����ܯ�Й����O&��y�ް+�A�C���(�(I����:��s�r�YC��W��PkjV��2s6�S����KȈe"�U�8ҼRtmvt��j�.�ri�7aͼ%�������6��ݝF�$�-%A�v�q� �4�\�f"i۾z��z
����Zk� z�������y&n@�;+�L�	ϸ��9m֐����P�:�q�0�:;SX����L|�ŵ�ڽ��z���l���S��m�m�Mb� o򷗛t�� %�V�B�c_ǻ��V"��v�B�>���t <T�:ۮ��cj���u�p�8�:~�J��4��r�.9�^�{�����*3�����X�S#��i��0 eoU��J:�(w�+�WR���.���K�jT+�	3Kn���r�++�?Y�b��I�/��T����7���(��گ����5D8-��%��]KYr��,I7mNx�G���L�%̛��]Z��uu���ܬ�9�=�6o8T�%D9&��Z���m4�aoe�<�<�0gs�I�5�,8ǎ��{�u�V�P4�M��oj#�p�L��Lgu�I��,8��4�y��ogf�SM��NE-3fP��hٹK`=˫W8]��v�r���宰uȒSL�;�X��K3\���Շy��oK�U;��븭cX\�o`����ҏ}ɍ��s���=�uϳ�_}������O߫�Dc�kk��4���;(�&;3v���J�u�q_#�Cݝ�Os'�**.r����D�����-�눀�WW�������~������q�3�d	!���,��{y$��!6�	>BJ�'�ZY$�XO0�d�bHI���̓��3i�	��� ,}��	�������|�T!/�ɡ�`LHH���yJ�z��?o��ϳ��k��?F+"�"�U��h�*��R(1UTUUb*1X�r؊�DA(��TA��Ѩ��"�GM�QU"��*�T`�UX*+Z�1X���APEE���*�`����j�,b�,�X�EcX��c��* �**(��Z�9��s������U�cƢ��DQ*��,Q���A]R��(���
���TV]S*Qb�EA"����TE�.��kH�,�X�Tb#b�b���媨�UUEb*��"��F,U��+�QDJ��,Uݪ����R���ŌFi�����#*TAO�X�b�g�5����+"�?5H��eUH@b�F({;�"�E(�H�(+����"�)�TAp���E�q�󢉿���3]�!���)DyB�DW��TĬT���Ѷ&�A�S�V*"�Ve�ԱX�E�Ub��Ve��+r���� ���1պ��֕D�DDUDDT����]R�"�v��UUQ�9hǬ�DT��؉���d�E\k@QU5Ub��E�bJ� �EG����>���E]{z4�k�c�UV(#i�`�Y��Q��Wv��h[,F*� ��m��4�ƪ�~�J�k����TTA�aG֢�q�
�X�Q3��X�"""��5�b������i
*���R�+���E���QG�be���AF9옌cw3�dDWI�
&��iQc9eY?Y*Ĉ9C�1b��!�`�����YU�Y�Vnͦ,U|Z�H��d��2U]6uZ$�'� ���.`1��O���||P����1�X�WX��_�������R�����GM�,7�f�Z�k5�E����5�*�u���ƱX��+"%�>��T}Jq��E�Z��٨�Yl*�E��.���ģ7Ju��aGT+�EE�Q�
77�Q5m�=���PU�4`�X�;h��W�(�Q�0GV���E�3�b�jT��2���'��0MYD���^�dM!Ub"-b�s4���Ab�2�8����ٽ��AQ�^�o١z��ȳ�\����p7b�QUh��/�~�W�y���6���&�:IZ'S�hTt�-�pM���뗺��(�;�c|��`#R�?R�Z+�(x�ɡ��?s�7Â9F�Q��Z����4�H�kxٺ>�5�/֩�U%�sN~����8�n��-�/<k܈m���+���@�H�]��2�1�UU����GT�J�B��E���Ö�q)Q*_�,w��U�W/�B[���⪪�M7mU�J9k
�D�.ZL�e~�t�U���x����P�t�P��I'�5��ϵ5�X��r�����q+���f���m3%�뉥Ǚ��L�9.�R����v�%o�^~�E;(ڪ�CT��ԧ]8*+R�)`��0
��q�W͈�)���xv�A�*�S�i/� 4 ��s�׻U�w.6ݧ챂��g���߻��9�`�1�"0�auW���a^�z���9l^�Ϭ���̓J�$�!o�E�8����w!����4&�Y�Ӈ����d����ō�8��pG�S�����;2>���/��C�ӕ&m�P�>�A��/����۲��@�(Ƭ�ҹ����Rл�	E���z�0��Ҟ����q˕ɵ�t߾ՆR=�/�{\٦}B�y=�*�ajDI�LE��F1-�."E�Sxb&%/&���s)��X�O���N�b��0�B�r￳����ٟ�FQ/�Z
墈9K���Dxʃ�g���Z�q��_�NS�6 ;� 0R��j�	��,�c��|�u�&��h[UQYD3;�4�8"z����lTϩ����_��~Lx�����b~n��QTSL.]�f��θi"�Z��K��&�O�DLID��c�a^03�����y��ٚ�����������m۴��DE�y���.4�y�r��R���W��[Aa��*����V-B���.8���&�����i��.�NwxCH��L3��g�iO����5�}�����C�k��5���#��;� @թ�g���m����}���Z�Yi�0t�`�`����0*Qm�X_�K�8�Ƣ��_��g���UVX�-��թ�b��\��G�f
���r����T(��a@�p P�F��K|���bg�U7����~�����L��,A5/��c���T��c$��{���8�SI���ͳ���%��g�]��+���������QeF�s�H@b�����'���3�Fk�c����\��8k@��|Z_��5JSw��5�����9}�Q�뛻��Xmя3w�3E��Nc�f�K��_oX�{��R���4#��j�e�-��d�"Hu��;�tU��o�tf���A�YP�\,Z���7��Mcj��CZ��sZ[)r�'߳�X[d��D������ʔ�0��G�M2ߛ<�3E�m� �-�_�q/���o��l;�w�d{|��-֟��/�����̪'�>�e��p��E�[v8kW�����ͼ+�V�ϻ�-D�!m��]A~H�F*�(�>nw.X�R��h§��? AvXnx�G��L9Ͼ�2�!���Q��3N��ol\r�V_f=�ɩ�(ai>qq0-�
r�ZK���;�yƢ *���,D*���"��X��QE� � �#U@S��)�)�J|EO�@��sm�+��Gb�~��k�����K�l�N����1Q�a�U�a���I��Zb��~�eޮ�Ժ��E_PɉX��5�y�̴bs)��x�[�ʽك�̄֖�2~DJK$0�`��ˈ���]g��sӐS�\��<�<0Y���c�i�6�L�u�%��|J�:����i-
�Y�ӳ�&�tJgY�K��ޭ��!�m ����cd�a�3�����䥺z�e����8	O�E�����t�D ~����!���F-M�}�������'�$~pG��L�( a�^�ۼy��#��8���/ʠ��H!G�SMϲ��W�����w�~Qbt�R�}�q�%��E�$c�(}�|��0~![��U�!D.G����=�.�
�p���Z�D�q1,/�d��Ɠ J@�߯W��V#?q����`�2I��F	#cTAt,350ZH?��8�}���, �!�0����yNf����u�"���	�u �����D��2��px�~J~a��7�a�=�.4:�xC��n}�n�fLdmR�s=�Mi��a�����t9"���Ӫ�ϛ�Q�@�vzv6|
>���f�(��v����Oش����<�f�P�~>(��X��A'36`�J�ѯoJ0 �k��9��˥����6"��pf;'Ͱ���g� �(��D_F�`�h���	��H s^��Q�~1L�[�=�!��7`�'���Tj�R�l2ZZ~bP�ܔ� �����B� ����Z�$5k|fI���(���CK�ᚽs<���En������$�ǜb�����U ��߾��t�e~�~��do��ϵ�b@i�_�[�SmD����v@C�7�0��a���B-j HB �(p�'�e�z����`+��^$V�W%v,f�����ӍP��/޻4�����{�j���,@�h���|�� �+B	�!�NFJ�i^��Dxg��ޝu�=�§�IV��물�� ��l��|hZ� CQS�*I��|�O� �i��C!"쿬 �&�'��5Cڼ�ʑ��k�)@�j�S����AD$�x4$��fIy ^���X�g�fCH�	��XH��j`|��Ƕ.�+��-��-��yY����v�����xx���˛�6M�O�#�8����-XٝSj��h֯��l���1+)����u�ϼ�	ٖ��L���v.�~2�S�n��Y�+�a�C��;����B�t�����Ι�U�¶�.	v�7g�x�L������Dw}����ܷ
`"�\����Y��3B���;)iZP��z,/�W�֕U�"u��z��V��D�������H6�y~`"�c����o`!P�G��7��G|��r�e>����	���a"��������w�� ���:�*�L�J[��`Q?�m��Y`�Z�T�I���È4K>��]�0f��O߳N��`����7�4�O�>6�]ݽ���b��b$}B��瘒�!;JF����ہ ��u܉%�a�]#��i�w����ş�$��+��ٱ�����~ʦ!�Z�%a���|�ݜ~9�	;�8[
�ߐD�~�^3J�VlTqN��GR�c��p�/ה!w�,*b�Bӎ��HX�*���,����c�?rz����Ew�~5�$ࢍJ�L�Q�����F���¼~מ����<�-0��	j~�^{��tt}�tCkj�O��U��}3ռ��:n��A�bT�~�	�d����������6�e��.�S2g�����r��\�����!&�,`D������f(0}_B��)��P��_D�%;zVp�����T㕙��y��ߴ^V !�APb����(��R1"��sz�5��]9=��7㹹(X��@|�O�M��+SM�OIӫ|�����b�\[�ok��q2Μn��K��V� �8"kC����:�3
�s-O�-2��%h���OAe��ߚ���'�/w}b�$:Pa�Xkg��ۆ��{�OՎA�h����(�myV�66&������B ڝ��^�o�Y�Ȍ���Vћ�f.�pq�uz�^.g�;z�'(rwe��k"�}��[�����f� 7��)w��3m3'XF���o:�-;[\���c������Gm]_]ӊւ4�zq���ή�C��ק�vB�|K��Gƽ��w�ն��UpЅe6��h�zب> x�I�A�S��$���^4d�ߘp�g��u�� �]9�a�Ҧ��0����s3󘍴 d�����o�}�pZ�OzW��j��4k;���G$K���'Xx���?��͸�`?P�`�ln�?_���#ሢ	4A�r\(3�� =ɸk�I"B@FQ���*�6:*L!\�(
dCB���v�'(�^uJ�'�wb����+�G� ���R���G�0�KA��)��i��
F�'��j!E
��$|WZ��Q���;�Ϳ&e;�uvk�o_��
y5�њ�W�+Ji{��
ՍA������$��e��l�o�Ii�\3=���z����?��$�z�Q^�H<c:����Qf�s����� E����1�R׆v� `�J_��� �?U�ߨ��֫�d��9��Ƿ}+(|I<
�Q�������о���<Dz���.	�:(/�#Qr��M��SZ>��>>>�m�|K����x2"���߾��W����o�W��m�lx�_# �\���L��+ٮ�pl�>U��DP��-|��
U��P�r��K�_l�ڣ��H8����a�"�$��߮2���k���>���7ڧ��Ca'� �>�R	�� �K�5>����_y�^E&�=]2j��F�\�g�}"ؙG��P0�/a��/7����D ��g����=�!�Z�ǯ�ewe_�F����OcP��q8���������T� ��$��M�a 
BI����'�����HhBI]$��a�ٴ �۴�� m��?! iϩ�o{�Cl H~d���Bm��+C��'_�!�������0�$M�TIR>�LUb0$QH,�ԀQ/;�?)t�a˞�����[Y�=�_'Q*��u�ɧ�\��rG�6nv�C���Yy��IQ����C[ �t�����^�6�Cy�6s��<����F�� R� x�H�A7��	� �[^%�271��H?A�p���`���*��Z ��Tl氘J�j"�D.f��fH!%cml�� ��n�,�P��,X6<� 
��5�V��D����#!,�s�s{�y���YDBxTu��iK�<�T�ORp�o�vh�Tǜ@6��4�#	����cWw�z>_��H��7�g�C�_$GbD8���
V��f�pa�T��]���P���̥T��M׼X:��М�~~�M�h���*��Xu��m�!l��t�u�A�ܵ�4!VN�x�OgV�ׅ��w��S�W~@�\�:��.���4�3{2yY�a�@���p����H�Er��&6s&�Kԑd�A�No�Ȃ�s�V��3{�cm^AS��qu��>������|�h� (�FA�EEU)�W�Uu*Q�k��i8AM�Έl�U�<�-P$(����<�_��9Vyx��W��T�K�!���(��}�^Yk�5���pQ@s'���>0�=rs���a���\`#�I���WY��f\~!�ﾪ�X+k�(05����Dg4^��H�c�͡��]FiD���_=���߮n-.�4p���箽}ި�Fu&�������Ku�:B����,&xa���+��ibA���kU1u��a I�bC� ��sVd��� ��$1���މ��<�a�F{u|��]�י�= �ck� %`|}d��<r�˴����vk�w,$=�b�"A�.e1$�Z3-`T
��B�+$*�~�ϯ�kw��}�;a�v
g�6/+�jo#6ے�7K�
/�\M=�Ⱥ��۳���+/W�${����]9yVx��y�N�M,4����z�vY�KZ^ �6�$Zg5OH�[���,i���K]ͣ+�0���=����"5�ܚ^�� ������L��,A	��IaY�W0�i$}��q��@�
��� ����{�>���7U��ڠ���O��"����llq�ͷ�Gz}��jI��ޟ(K�u}��Nn*���$�1&/��b�sb�4[ҴF艀���Xm�g|fQ�dw�w�<���N��4�1 �o�0#=�d���];��%��.B>D�O��q�ؗ</�����R�g͔+��V�g냕`\��B�߻���_ۙ�a����۳bsFe ?x��������" �]Z���n_�T5�}�"������,%�^��)Z��?Wsu({�
�j�PzC,3:Dϥz�\n��3Oɿ�🿹�Nwx_@>� g����P�a�,�{P����j��Ӳ}�ꗻ��g"w��v)W{>�
�ǎ|��`Η�7fLA-N�q������u��-36���q���4~�46#���{	ao����6�|�ďՙ;4l��:ʺ!��^�O@�g��C�^����H��]���5�m32�Y�ҽ3E�7��y�^h3>N�)�	?�����C={�ް�ة�N��5��d!֙����-ᦸ������!M<�9�)�b��S窛�C�����|���]ݙ2jx'S���go%��@�Д$G��g}N~ۀb����-ߞn�ъA��DGL�s1:�G�� }�[��DS�xC&��1	4�rMj6���!Wgg�bVJTq[s8ص0"mu�wIuw��6e�"<���U����|J��H�x}"X5�6K�F�#]�C>
��&�LD0�oW����`v��6O#���v�Re�0���}y��"W���3��:�������G�կ���X�^����nS�~y���2�{�@E H�H�����P�;���߹�o�WW[]�\�^��[��"�
�t�ʈ�!�� a*�jBn�ةZ����_�]�BJ�.*Ѡ/{_�D#3�O�tFA*�m{|AT4��ut�_W���1/�)sL({琱T� ��J��-��^�H��8Fh����u�S��ԣf��1dE�wC��M5��/d-SF���č�,��?Q�Y�U�b�]u>�i�w�$�?R�!�Cﷇ.����^�\��[ҋ{��{Yn|�h��=��أF�u�@�c���5{t5��G��۝��^Dg��~��#ҙ4���7V��p�r��7�ҹ%u�^�V�Dp�î廮��
�����b�<�H� %�3_}qޝ�o�lW����Җ�JήV�*V�X��u�!0\5�=YS�������w�O]_���a�k+���״k�Yu;ZX�:����3��`2	�� _��]��ۓ$W�Ŀ�o��^��X�y`S�ư�7�{�M�a�Wجl4[�9kx�k�햭�\|�c*iͫT@�s�V��ϯ4W�����;5���*weݾ^����}lm��C\�ܯOI������IUTi����w��tjީ(K�^��2K&���5~�=�f�e�������Z�/��H,|��ڐ蚐XގM�>��޵�g�v�~ϑ�^'O�.��j��>�%�R����/g�z��'ά�6'������,���φ1��=����ʭ��X��w�O9ϻ�~���Ré�cn��?g0���%��gSU[��\�����`��M�ö͡�{4J�ag�{o�p5�qC�ǫ�vr�k�850���Lˁ�a�d1����Q�}��viђ��5z��o�;�"
�0��:5�d�����X�&W�<���\�~�6��k,�/.qj��4�^�Οkf��/Ɇ��~���w�9�{�4w�;�?@�p,~/k�W�~�,���NȺ  >fT�779�!=*����G�����d>�O{kp�@U�� �#lUUX��*�0U��}�=�]�O�w[��g!}M��8^n2��yzwJ/�7���,���j�#:�N`jK���|�tL�͖����7@���'i�Ǡ���=����쥠�҂��&Nx��dz��t��[��Z[��lnZ�0��m���h�������2	�5���ۋc�&�A*N��uY̓�U�Ђ��Cׄ�I�x��ЪY�:;�+:&�\ӱ�����pQ;���k��5�����lxU��uµ�������~�y��k$��BL�5����!�_{��;��o�}��T=������(�p���]}Qv���+Ѩ\�G"�,_U��Mב�8C:J�o�tZC�k�9����M���b��o�K��_���'��?g�|L�?*� ���}C�p�9�B�B�B�%�����L
����z�>��K�r0�J"��JZ�Vl}�r	 ����IX0�n�	wg_1���������4Ϳ
��5�k]5/���������V�sEN
ژ�M��Z@��x�Ks-��8~���D�{���[C�L��w�S���>���S��W�c@��sw��6�]e2<�]	^�m
,�3s$�b�n������ ^����ŉ�y��z��1�۸<r�4U�HĖ�%��8�%�nI�3���N8yȩr�a��:����6 ��ᙆ����*��)n@WU�+n�O0�[���yȁ)$q �9*L�tm꺻�v�B���[}vNEK5SNq(�Bn�����G��⣷2�,�N,y�dac��-V�v�@̦���.��:��oL$��yy�o����״�1�V{+T��s��Y�y4=<��e-!���n:-Ӿ��K�h�=*��fܽ�We��v��-s��X��G��vb³W�.��p�ұ���,қ�%b*�U��w(���[s�^����M�p��0)�����h(ٕY7�����[�m[�/�~���d��`#bϞA�j�I����Vw?k��R:�.�P�?�5d5$�/5�!�5�r��h�س��%� b�)�	���x��0yj���L�Fzنwh<�[h��EV�)\����Z���fV�KO�U�ӭd�~QG�zf����ɜ~K�������ջ\�}�����:�gY��pκ喗Ui�5�f������d��f�u1n�m�|+�J6���s'-���Wq�rFx�{W��z��檞}��2u|�;�-V_��i��f�U���V)�XS4���h�H�gc�z#S�N�r�e�mn�S?^�Ň���~ۊɱc���tR�<��j�B�V�5}!�"I�t�͎i����q�ozl�����m���mF�t�ʄ8��R\k�]�E�]�l5�Z��f��"Xʽ�M_�ֿu?|}�"^[��������2��s&X��j��N�jliȱV�m]C>|��-9���&!�}�|,>­r�U��^���	��;{SDu?�Ӧ[O������5�A0���r%�:�N�[Ӗ��k�^�U�5:A��v�i
�X:����3Y2�wCҢx1���;^R�'뎂Tf�
��W$v�5��@S�r���8����-e����S��\�E|��a�3�P)JC9��l�U���	*lka�����@��q�6�/�Ξ�͛�j������Ƭ՝
}ε�_E]������u殾G9){r��=�ŭ�#dn�>0c�Q��TW�c�5-\��8�+d��Ò�vk*f��ǥ�]���ﾬʬ�tF`�5Nj-i*�K�6�V��}+CŽ����wZ��+�j�_u$c�pz�>���eS���o܎�����C�m������G���4Ry'���?�9q%ݓ2�s���� ��ɚ((����Þ�����b�e�'�r������	8ɜ�Xß}�PPݲ|�������7��h�:5���˾�YA"��">i�3(�Н��4��C�����QG�OO����<�\)���������¿X^P�QUE��J1T��>g����6��oXM�i�RL�`���I�Yon���o�d��0�}e��a��I�7��T���!�?������ 9d�X����;�i���0��40��~�Ͽ_�C5N )�_`q6����Bb"O�I�מ�I,�c�oܯpI�����)|�2�������pg�? i���nXm+iS� ��-�0r�O�+';��F�YPX���������j����z��/Y6��g�N&�/�x�M~�/�~���k�ϯ�Αd�
��q~CHi5�ϳ�-������N�ßLfr�;M]�ě�+���ہ����߿�1H~w�ou
��h�O�n���-������sz�I���bύ��,��	4;ҥ�'o���<��09� ���?3y̆=d�a�Ҧը~kԹd�� ���O��*Tֵ��E�^�u!O[�S�wS��m�6�R�(1�������\�����;�1=�>�.��~��<}фt��0ߪ���| S�N��Z�����K�vC�MӺʛ@x��L��F�&���z�q�m�X'���Gȉ�oeֹ�	�G��z�[�Dgy��r8���	nG|:�
���~�o��R�/�1M�����U��FA[���� d�q�n���l�Җ����;2��f���x�g�L i؈Q���V��֥���g�G�r'e;�Dr���
홏/��0��>0��'��lL�G��9�A[K�9����,{ٮi�BJ��20���h�����d|vw;�������Ig���(k�'""�tΥK��i�*��W��:L$;>!���w��g�,_#=�	�Y� }tZhV;.u^{��������èo@`-g��t�T��HĤ~�i�'
$����ޔ�Ӄ��ir�DY��t|�C���<>#��ڔ9rmD�JϺ<��̂% ���� 1�$H,b@�=�ϝ�{q׷�J��ȃ�T��zc�^u��Un4(��w7=��g��ȓo+�#�{�t�~:�j��22�O��3��-�P>��A��o֙��C$�0,af��j,�1V��B�^�Fx��w��_ �/�\�V"`�%`o 5��D�C��7��yu������DC���;�G�Ut_���h �)��]��uGթ�g_7�04��^�{�e0H\Шxn�1�վ�.k>'0n��ő�H�_|��%�JQ��G�x��п��kI��9��@�^Q�'�]�>�a>�Fӎ9�=��!t�9H��*���p��D��B�ÈW�v�]�R�uT|nzN�#x=.<ЙV��?!z< ��ȳ�|���-�e��=O�6�S���3���B��I�C�#
R�e�k";E��"�Y���B��d�`b�A��8�F�蛣��
/�;�o�3��j���*�zbg6���HT���^�Їp7>�w���  ǥ����Fs�xP꭪8RS����s(�} ��
���Z�33��XW��s��s�Mn����*�\���D��"�����w�h��|��q+v�egub�*��1N�$�P��<$鯞��0K�8�c���J��lww�΃�G{��=~K�K��q�-����;���0H$N]׃�GK?=�?AZ��{�X(�����ё֏
x��(GomɹwFd��1Ր&���Ul�½Wj݋���}3Jq��| @�J)�.>�����6���^���Y��1߱���bq�G��T���]N�=C��D�^�ѻ�����,�Y��n�:����~������M��<*���|����߲��e�ߓ\�c�F ���"�HxB�@ � 6�j���S+�]2C�"�NsL�=�vr܄r˫�H�VD�@`�Z��ԭB��/��}T_\�Ο�F����Oz��ӱ��@����k��'��oý�͇�U�z�B�:7�w�c��!H#�./�_4f LQ���MD9A}F�ug�ʨ?wX~�=S]����!�K�����R����>��.�;UF}����@7�U"N�g�=�r�V�Ug��A:*u3�{�3�� {_ibT�#۞?�Y �A"y�ӫ�I%V�͗���G����9�Dw�ǛK�p�"���}Us-��{(�߸ۙ>��=�T7�S����E�P���^��#wS~��B�#�Ԙ��yD����|�o'.��~b;	>t�x�O���!���:��{>�^4�O	"zֺT��_�� �oO��<+�@��)����	�LwG9�7�N\��Շ��X����A��E����v�q�պ�О���9��*����j����@>�\�����U�\�Ow9D^�S��/T�v����a���F����&d�C�C�\T�!g��9����b�|�߭!��n�Lڞ�� A�����柏78��S����Gy����b�/�D,[��kEv�=�q���?3S=N��ꓴ���")�]����ކ4��{T�� �vztΨ��^*~���|����B����*#��̏lQ�G��V�ϔ���
���xb�2��}�.5����5D$�+�S��QúTv=�j+z�
[��Ts�5�� ߮r���3�u�]��n�a�l��rq�],����I��:����2�f�W��6�#6�����ph�S�f|�su���}C�>l���'��4B(�[� ��J*y�>v�<Z^sGP=n��T��Ho}	�n'2�x��26guޡ���ڔ "���;���&7;�f)�2����.0y2�Ҡ�y�M��(|�o�>־�#C�nD<>5�S�27<ݍ��iw�r�N�bPaB�c�m���4�k�ȟ���55YN����l�s����}�l��`���r�k2bv�����3Yމ�ۥU�?�o��jV�fH8�+�rB�����:�#<Ǩ���������{B�w�g�b��S�͔��n;��1B����}��f����;��^%lD\ә5sǎ�i�n���r��X�D�Y���R�Nc���8.�l�rd��,�����*�\�hH�_���![�[�{��]���+	���]�; }:MCyV����D� z��޸8��ө<�|�ﾐ~��Ɋ�k;��|<�	�A�Ǌ E�z����0V��^��det8Q||z�@V��{"���E���N��BF�1P�k���#�Wh���U1���ih�j�b��ask��LO?�!�x�&�r�7�_Խ��a�+��(�s���r��r7�_e�*Uy-�S#��!���9��CW�}�ٝH�*6Ǘ4o9Ͷ_�x��d�:�t�(��ѫ��_��?le;
b�`��̮
��	��4;��7�d՘tرE����i7�!�=��%������]���hǚ�W�tgyG��so=�Q��9_,��L���S�VJ��-\5��S_}[BT�S����c�����w7�Q��ɦ���8���IHQ�1I2<v)ۊQ��t�x���{�.�\�ܐOP��ni��fd]Gܼ;@���@"�4)@����j�J����sX*7_��N= �|ĸ������B1��zg�k���EO�hY�^���lY�s����.�.c�g�C]���H�d~�,9�!��;<�o����N�j�����P��~��k��RΈ���́�a �$8��z�w�~��K���z)����M�� �sJ{���s�f��e��')�@�9�����7�+8�׉;��Ϧ�����}��|�ِ�Y�qH;3Z�G:�����OT����,\�´9t�F�8��9������V9Գ���%@��s.�ؔ
�9�:��̖�c���-�Y�}�X0�B�T"9.��_��ɩ��0�;�����$��]��y�G܍V��8{���Ή�N�S�r��}@����C�ʤF��Q���B,G�ý}�w�A�!4�>�lP+�(������G.�Q-tUM$<�������5�"4�n�˽�'C~�@�п@|m����[#L����$�+�Ն�}��p�� � ���Y���b���G*����rA,~. ի~S�w:�J/ ����=TT9��:93�<�5��S7�lߏ��}U�0k���Ox����:bb�tҕY����.dR��+*�P� ��ҏ��/�&"V���^t�ߴEJ;�T��c/xh�L���ʗCz�i�_��ߥ���s��֞��@��f�t0e]�m#�����H������W]�"�]t\5)#0l
Ն�����"A����l{�#�1��\��aR(/Hϧ�Uzc��Ox��C�gh�1/���r	Y��Kx�ʣ�{����z�ۊ�dԩN����7���\#�qD�;{�	�5��� I ��\n:��}W3����W{[Gy~U�x���߽������6/�5��ݢ�Iy�o���}�^me�	�0�Y�x8�UlRlꦙ ���q�y�>��4kf�6#EAW��cmb�1EX�T7�u�z�gT�=ތd����샰��	�ݴ/�f/�V�}F�&��#�ʹH�>=�L�$���v�֮���Ve��Z��r���-�o���Q���Vmb#�t�I���H��Zޚ?Wi��yc��m �\2~}?�y�f�֝��>�=3���fJ �l��g�K�3�ޱ��F����!e�=�󐗏aRO]Y��!���^���ǳ^SY�2e���R�R�=
��3� ��3�x/��:��RM*z'�频���M���I}�9O������I&��{�X��:_
�M��*V�?��q؁�Y�;��������sts�G��6���Heg���5����p(�����_}�F01I�!�t����Ff��>�P�Q��B#�)�Eʘ�J��:�-)����׽9&���yCO;���U
�4�qcWD�$�ӄߣ���D7�0�*�W�*.������bZȟ<�5��{��#�w�{k#��9�C<�<Ő!j��(�B��H�?�~P160�s�"v��˝���0xRj�l�ǜ�=�@���fǑ� ��OW�{Q�m;)~�l�[��ɢ �0���޷}��y������"U�V/75_j��:~5��=�u'�&Z������7�#�Dh鸉�Ĝjwc� {�8J�]�<�
���_r�w�'�b��}oC�_�v�n�TU���e
6���jȶW<�Ǵ�b.T{�}[E,�ۓ�����~�U~�a��ӧ���Γk �$�H�]���AN�.m��A�u��SF�.)��FzMcF.�:9��teb�����sy\"�=54����yz�Y��y�x)um >����v�ԗ,1vߕ�	��\,ֳ��U@������d+�0'Gu��p�ɝS��Q�__b��L?��=�z�^�%��P��s[��ۨ<���@����h]zm<}y3h�B,}�	P���m���1�bj`?�f���\zl�DH�}#�������j�O�ۯ�!%��¹2�f.q��rȤ~\�b)
�G�,�q��O�s��Ӿ�Q޼�����dT��@�u\�z>��� |-RE�6�T�}foE��<
�Pݚ�u>�{D��y��{�K�"0vDI←�^R_?�ˣ	}�LXс֎��&�KY�r�b���!�(@�s���q�����}i�큐(�bF����Dmv
���ʼ���8����nj�9���=0�����|綤:h0"MG����ں�Ь�|+^o�f��w�7����kULg�P��Z#�1F|�o�i}v��o��t��	tD���5����20υ�*�	G�/g��.����	;��z��<:KYS9<ȍ�͚�=��AV6�V��S1|k=���Z������BI��ETb  �)>����_U��׻~��o��yzd���`y7x^4:��cP�%�����|<;1�|R�?��|���۳4��;l���<��,'�
��W%b"��T�``JІ��"�G��_wt��pmr�ߗ{m��˻fQ�J��Bb��]�)�S�\���H��u���-�uZ�C���8�
 �녭�h_Y��Q��cd�2\(e�@�t��X�A���)��16:���*�Z�T%,���N���7����ZQ�"�;��|�����-��xW޿Ni��/7Z�W�]�B.eGn��O�8A	����6��H\FuM��*����@�a�Q!�n<�܎�F���&�<.*#�C��wt�"Z�';�&÷��T��� �����tE	���hGd�l�@(�`�z}�M��=&�:f�ط���ۗH��g���	P��yb����.;My���ӭ�9F���B��za�43��Ԋ�-�X�2֥��u�|>��8��(��"{�#�J�����s���x��v>_��~حQ^'ѳ�j��߮(�I���k ,ylz�i�p4G����}���[��%��F�l{}Qw����#e|TNؚ��B1�@?��t�����9�s\�_�ݱ��+��U����t*O�t����?)��gf.�-����lpq�U�^��՟rB���f�h��DUk:co�G�W�ډg9�{!Q�]�����v�g,��sO�z['���YO�.?EeDx ����sPc\C�P�u��`�����ׂ*8^؁����TB�Y�6R"��v&r[z�Վrc�]�׾�O!玕,����ٶ��ü�lVh�q�ո��gc�Kv�8X�˖�2�3�
,����$��5��v[Ox��v��w+��0���1��>�!�U�o�R�,Ә]i��Ȗ��z<n�'�x at��2�2f��j�U~����(j��:(�E��>�>@���Ff	a�{����~
�^�lI%a��
�c~��m���ȩd{�\���q�ئ�q�hd]c�3�C,jj���N��wD�oG�|&.խ�a[��mk�������X��`����"9��]�s��`����@v`�[%�)���⺥;��������!��z`lD#S��L���F3��z1k����E����6� �j��_r&�2%"�ָDy�u��^�ȅ���qg�ʊa?zɓr���ՠ]�}Ep\��?��7y�+~�����Ȧ{$��p��m��d��ك�ю]��biC�o�o|>��o�Q�6<���Eвh�T������V�)���&�4��hm臲�Ҹn��yN<�t�%�p����0��ʧ����.s�����EET.��g��Q}��տ���4c|�H�R@��v'�Q�#>����a���P����{���H�G�O�ʠoz=NGF(�2Ъ�x���.�	���;/"Ҙ}"�(#F���Ft	���Y/b�y�\C�	��a�bf&U`�'���u�;/p!R���6�N��wV^��)K�Փ��&u��w;�(֔���Q��mU�uh�z����,�tjH*��&��ma�Mt�b�G��)�i�>x��qi7K��1�m����NV�eO��{7��c��:�p)�\�
ko>Ln���n��i��3���i�vv���"/���,��YN�_j,�S]��&�w��_f��.TX�D�*Y�|�W�T��]�8ٿ��j�34P�m2cUӓ�6BH	)D��,�W'������ �8���4���뽦�p٤���굲��G� �q��u���S��O�^n�����%1(.��X���Q��囊f�E��:�bV�(����jf���ѳ��-gZ�Ws+����ov��S���:Vy[͆���� 	}�����'r.��i�Xo�BҚ�ʤ1]-9	�]��dF^q�7"�瓡��:�c�Hn�p���E�7%J�9�A2���S���u�Fb˼ʎ��6"H�]wV:¾��:@k�\��I}ڜY�\d�N���E�m�*n����ut����3~�����ꗊ��_K	$�,k��	�e�%��������_$� � � �u�(6�Ϊ�4��Ε�r�,}ȝ��ޞ6]��:0{l�qP�7��!7��ڻ;�o�̈"��9��5� H��2�݌�|�!��,i��u��hI�h��:�5��q�t�	?֙����%�������yK$#���$s��[�����46���N���A�ϔ��N�����V�j�y��{6�2��F�kS���\x����J�vgwv.��\��ig;:�b֝��G+.Tf��qt1S�l�;��<��� EVJ�Q�f�Y0&YJ��}��;��s�{[��_d�n�ki�ï*>���f�vg O�6�X�<��������1���9a��N�Q�V��/oLr��Z��U�+�uj�e0�*�gQ���M��P:�Q�m��$B������n}3+Pw��:7�nފ���ۭ
�D�	o:�����w�7���#)�>�F����8�i\�oZ�.�5�����1Auk����o�<�#�^n�8�f��kb�`v��ǆ�<*�ê��&�ox�d���_�Mk�F�>ѝɖ�_-c 鲗D�p���D%�t����r�a�݄/�++*F��~���#2D�w�7�ת��8	���Lkn��zV�}ṟ�'n�]7�h�ն	�V���и_c�d�5���Z�ȳJ��� ��iMat/�q�[�o	�X�ٶӳݚD��w�#O-�5 �����.����/76LG�mi�n���Wl����;;i:���|`W;���'�g�����tp�]T]ZF��N6�:�c<H]�ؔ�`':�l��mr�O,9N�/�|> ���~{��IRqxe��H��b�v���{�b���ˆ��ژ
*֋���YEJ ���+fZ���ə�S���!m������5y��-�>���p���b�_�s�"�:�D�QOOtPr�0=zjp����-�j�"-���?+u����D�>s�o�"$�{�	���R�ϧ�b���̝[}4����#�zȘZ|�ѭ_����qGA�� N�����K�ƊH��S"�L�)Æ��NPO�%y�^�zf5.���!Ҽ��tH��\'�j�f��9+b����Q�y�]�~��\<|��q�¸��?YK�+�S)�k����&<tw�F�����z�-_�����K H7���wI��a�X��Ϲ��$3��j�<>ȓ�57���[���+�}�~��9$P!�� �u��r�g�[�e"�ĝ�Y�D~D�{�3�-J}�bۻ��j��-Y�Yg��َ��pn�KO{7Ǫ;Dn��h��b�� �tA\��e�{bG�}�a�Zs�[|5�[y��
�᳕��6R4;�b���{}(S��~ڵ�<K�t����U�2��[���5������w��q���yd3]����6����.d�����UM�����}��Q�_�F(�\�EW�ZQ���ˎ���1jMz!�ˮ�u��"˸���4��^�8q O� �>�������N�SӦ9��<-pFv��H�84��_���çQ��:��t�`A�N�啣1I�vW�
4��U����gm�%"���D��g8��S�+�_A �����#�	^�p�]٫_�\���SB�f�_S9X`Ek9Nh�SSc�]�g�y�{n}��9��sѰu��C��_��[��_�^���ܷ���TQ���eJcGx4rk��x����
ʪ��<��<#-wv�V4��L�9��a����`�J<u�.)�|��ޓi_�9+��O�\�h�����*�����5����Ӈj�xb���|q"�f#Z��J�����ɝlq����ȸ=����`ŖT�i�������5
��!;7�\�Ţ����z�P.���(O	q6�g1Zv�e��8\Y�XΚ��ob���6�3��LFº�o(�T=�>��~�=9_��t}خ_��Y=�
�)��O�}g~�B+��)�j��),s�"/�[�����]=��ۮ<���X[�D�Y�YW,�UhVZL6���g~�.g� �Q�:_�R��:'���ͳ�ջ$�q������2x��SJ���>�0�3�����l��
�MNBx�o�<�>��Wd�+�z����/��#\}�}�ckh��^ޤ�Q�U�����j��7�i���~:Ƚ�Y��4;C]�>�)	9�;Q�e�e��8X���,�q�1���e�.��>}vY�5֨�I1�/l^���F0�iY�"��߂�Z������|�οo���]��ğ>�Bt�y��δt�F��.r>�+��H��v����`��T������%V���Gh��C尭,�55�oO'�כ��ǚ��J]I�>Qg�]U*F�u	>c
L8K��,�Uq3��qNR���p��k�#`��%ڼ�2�WϸL8��A�9q�Y���"YE{���z��\�Ƥp^:d3!��b�Io�xFK�B�eKAbz�82�b�8����g������ᝋ�[��
���y��L��H�@)�����>s��&�?~�g4�;�I@4"������11q腃������E��mY2"�f�̯�u.�q�n��kҙ��e�oA�a��sh���顗J`�Bw=��HkI�a��v��î|nG�L�����a`G@���L���� �Dl>�Ԯ��WZU*|<ꗳ=��E\�I�	�����P:�y���,
ߐ�j���W�����;�ڟWݴ�'Y��}�3�9�K�]Ǔ��w�<c�Oā�|N����әEՁ���5]η�s���Y���ۮ��Y�U*	|0TF�k���o:a���e�V���Vy�AlVO�d	��˵��G2�?�><��������^�����RJ:�.�9z��Y]�؛U<s��\Z3
F^��G����]T�R���k�g
7�~"��]m���c��R�*U�흈�G[6*���R�yjk���=�Ʀr�jl7���}��b��`$����_�w���vz�����iN����[t��K�M�t�o	�|�f+�Hs=�P9�v��uK�qNmH-��t�7w�ꆵ,�ȓZa0M�dgo�@�`��(Tf����v!��	Dx`���x
?|i�f�|'NWW�H@��IM�5GT�tbQ��L=��r�p�K��g��Wz���Evf��S[����"(d@�Vb�O	2�K�����A?Ţ6r����?���z`��"2$5>k��[X��C��}/'vs*��a�뾥A~���HQ����]�S�U8�uZխm2�����l?��;��
C����cѝw�9�Z�x �}�	/!q8�������5���5�����X�z��'�L�!J{{�����
�ڤ�D_!�ׂI�bi����L��r����c�����G"cĎ��szj�˲�R�ᢋ�������&@���Uzu�!U�V.��S�<m�;�7�!Ga�wf����C#��O�ki_{yW��������d�V#�Q�9�y�>��5ͩS�:=WP�x�/y���MA�O*Me�ҫW9c���}4��yԻ��5.·��i'ú� ��AAc
�N��օ����dޝ�-Y�CΛY��G���Z*�
�Qb���aW �r7��u˩�AU���o���H�T/�Q�P.fԼl��aĆB��эM�� �0�7�N��>�{ry#�����e�3�N��١�O�-c�^D>~�LGZ��ymw�O���_ѣ*-������
��.�S��h=�9��=��_;���c��4U�D�p^,2'ZзB�C�>���Q�<fG؟|G�.�4��z��"|���o�ʙZ���DH���5�У�?|I����Dc/�e��;\����̞��S��[��&TB꘴�K�uQyXf�₿L@ܷWobv8?4<�H�ɳ��C�S#+�b醮��tq���|���鵮C�⒏m�-��6����x�X���zuE�x�e�\Q}�]�d@[Su�I�ۺg��A�!���0' j��d7꼩ʥN��:����%n]uey��%re�����Ge綗�L8����U� �g1����2BZ����6��F�)��mz��&	��| Eq�N�zR��Q\"v�X��כ;��^`�܊�aM��}�|�;�<����]���.=����7�*�kt��̜HM@�S��>z"���AQO��!��w�n ���Ǧw��ױg�9r�l\z0�&�!
�u�����ƃyG�c�6O8�i
��p�Փ��n1*B���@ ĉI IU@�g�_u-z�i���x:Y�f��1��J}c1S�z�jy���o;]hp���n�T�o��=�-zQΫ��s,T}R��u._u�X�v2>���H��Gؖ�^?vKi�a-a}���T�]�����~��������p<��r��M��g��A�������]�,'���R���ؐ�W>�G�Of|���1�~�n��מ�'T�����x����ļ��Ҙ�S�_S ��A��P�3񃲞��>;n��s���ۑEɗ-P�ɪo�,tܣ�F�yN�慞�g���3�u}�E� _t����>6�;�!��X�#%R^���(�H�L��>��<��{�~�vL�|�cW�dg �0�"/(gV��N��`��� �1��>!��!	���.a�Ks��f���7�����9z"K��7bn_��lsv��nK5�����$c�ޫ��+nC��l"
�Dqoz�0������N�p���nظ��`�tY�1t�3�Qk��W�3��������"���pxT�c���S���Bu-�2�N�{Ƣ��Ƙz�|֐eB��t�2�L�n7xP���}�}j���e]�����1�)�����Q��������֍�����ob��)�*wt��#9[K���nP��К<����9��̶��<'�� �$��Y���RoU�Ч�����ݾ0��$�M}~_=�8}�����T#lE�G=�#=��$�,���o+�z�E^35�Sm��6:�����ݎ@tq}�vM�&�!P��a�rV��hQ�D`i;-�jO}�����X9R!1�����El�҈1�}SJ;zW�:�5��UGT�}�+P��C&�oI���W3��R~���2W��p���X�HC�R�����:��]��H����ﵻ}�g}���L8�'��﫩1a�	�7(��j���ٌ�;wֱ���2:2���SB�7�j�-{%)q���=[�gTaa��'}��^_.s�<J�]�S�>ҁ�:9�	������ZL#2|�����}�?G�A�]�f=���E�u�u"���͞��H��Onf���[b_��zR��F��W��gĕ{����'JF{~��1��U[��O�j"&��þ�fQ�i��������n'b�����dB�]��&(�׶l2��Þ��>��ӓZ�12�-���6�*���^^�hЙ�:�K�������J�4k�=c�%�p>�s����T�S}�jD�B[�<���}K8�~�S�U%��\1�;OP�O�j��۹A�����~���C饧۟v|h��>��3c��R�� p�����@F1q����d-<5׫S�u�Ȼ��ҡ���Q�X�����2> .t��F�d\��lg��� ��)�v�v7NWM�|J��T h����
cA'���$XE���{��� -X�x�S3it�����%��Cꆜ�pČq����Eą�d�9A9\ޥLa��ݗ����;�B�{k8Xխ2_<�,��W��)l+Atas�jv5HÝ��v��(�{����;����L}gϸ��v�>�](��f�Q�Fv�zWϼ��=]]��tozsq��ޕW|�����g)>�����W-~ܗ2�~�틔	��=����u�r��>D��(�]�	������֦l�T�F̝��oJ��2WR{kh	��> �ߒȨ�M��[�S]r}�ݳ�:�\;�n;�ú)��9`�GnȦ����}�2�G��K����yx/a�'F�04�[�<t�ֺ�ҵ�;G��Q�[������Y�]��8J�Q��>4�;Il�#�����0��+�;�V=�������/��P?��7���r��D�+L@���)��iQDH�ݯ;��!��O�)��r:�D~�~Q�Dg�<,xp^���_�A=�!vl<S��-�Ѿ�7m�+ޗ7�M����6�t#R��cD˭] ơ��,u����B6b�A�8}���1p�G�/�똨�LV}��"N��QI�s�B'Mx�*3PKb<�{�N���F�T�u�˕�Ξ�m���3�O~%�y�;y�:�R|]��Ud\��[�.l�P;HV�O z$�İ>ָՊ�?e* �ɤ�P��F9���7f��_|5�Z�*l�Gj�h;ס_յ��7t��;/����y�U�w��О�>��ik]W�뤛�T���b
�z#㰅G礰s>w?i�s������|����6�������n���(C�F�
N�%lz}�x�����\]s΄^� �+�z����q鏮�*����;*��|���lЇu.��5�S� c��Ճ���g�}�Ap˯+������xG��{;"1����#�Z�)�HN��[���n�B�Rhu�0W\�"�0������j�,�P������������ݸ�w����7�n�3��|�x�GQ�g�b�]WP_?"��O4xs���(c٨���Y$cbWLr���Q�f��$z]�-��TdI�!d.M�>�ۋ��*�H��K�u�y��yP�:%u_�F�r�}�:�P�[/�5����~n�����vH�0="+� �� � �iI��F��#�Φ����8w�U� C��f*�ж��p�Z�ǅ��Ϲ���%��D��^�fE�!�D����;S�ҟy�� �Hs�
�������h�\g�WK�:��|_��,帢�>#�,��ND�`���-�]��W��_·����_�r�r�9p{��';�c2c�3��,� �ݤ�[�o�#6_A;�v�k�#����{�ӂeZ%�zn1ħ��|�ή��TY+����˶>c��՟~�p8��a-���'O�UR{d��׀�];�O�E�-NK��~��R���o��F���/��?T}0<Ǆk�Nr��0��~��_o�釯��;Y_}��9�e���*��1]���2�]��l����j�m7��w�:��w�H
�-`�}��z���y��7^����s���ü���k�����?�-�|�~��p��ٓ|���&=Ěze��5��1�rc������dA�YkBF�t�,��Vi�]"�G��ў8�{�=���G�+���Ц�ά�zwG�y.��~]��H�/�9O_����\��e�޿���Py�;삚�>R^�M��Z�F��6or&p���S��i/G�t���<F���{k�ރ�|i��	��W���Y1�L��!ײ�H�C&��VE��샗t�X�f���t����kk�o��۵�0P�	�LJǻL=^���U�E���\��C~Wo�޵#b�v���=��%K���҆���۾wz��U���}7!qLV����|�$ތdݺ0��T7U2",ዿ�. /#�b��w���[�5���4\ܵ#}j���c�ҹs���h���C��s�9i�r@��]�j��>n��6횾bT/U�Ȼ���M�c����X��F�Co�����
}��1��٭���4@?x�׍�������XZ�qI�4y��m�|��9�C�Uvي���^j8_0��*�ы��5oPG���)�
/\`�K��yaή7�wr�w� ����JYX���5)�W��bH����k1?
��������T&&$C�DZF��g�W#��Ӵ��{9��j&�_��Ptxn�o��|hNM�U��E���p����k�:%�����՗G��w*<f�[��:�ds����_g�9�GR�����2�f�d%~�t4��Y�}��a��hAi�]����nu2K�)�l��B��y9�Ha�����]v�)o1�zk�
��n��H��2+�3����7�������)�շ����� 2$i����;��2���T0�=�",��v��'
���"�>�ʃ�����ʂԵB�:ܦ-\��N�W�^��u-�jۗQq�V��jK���6�G7�Fv俟�c��J��P����ho�M>�h{*����%��Q��2������A�M�u���a,ܑ&� ���7�QW-G%M3�����$����]%it�c��KKLϲ�<niKqU��^$����H��"�6�of�����SN�]�b�MJ�n
��d�X��q>�Ώ^ss�kJӵ�;�6�=�:Jg\����(�P	�s5A'X��:^�_ �W&��Ԩ�WK[<���Q�Y��}��Wq�(1vu�J�ڟ�i��S��Z�dk�&���kG����v�4|^h��X�O�����y ���`Q:!ܷ)#N;ʼ�ĳW9��*cۧG��v���ţ��w����/*�M�pK��Y;���y8'��,*�qe�����m90++{{\C�y���!�'D,�e�s3dY�k�@��|�4� ��$A��QC��w�^M�8�ܱ�W�X�a�B�<`�����:��tə;dy�������,�'B45�iwo}vҫ7�c���k�m�4�-���wqfcc%����.�-�Gf_v�Bv�.&jEۣ�[�[�Vk�8��u�r	��d�m�T�L�dGǈ]Y�.� 7Ҳg5wj��6q�r��]a��.��j뾾a㷖nwt��w�&^'c��V�-+���r��ˣ��C�'X�[�`�v����mt��+t�;�`��-��I4��}uj��`���3b_u�{f�]�F�F��Ws�՞�8d��e��*Y]i�V��Ǉ�YN��+*��n��1��/�w3��o��n'EP�?]"�:q�5�Ӷ7N"V�Ԟ�0��Qk
�����j:�a��t�,������`kJ]�S2R�RV�J��oaF��5��突]���/'WW2F+f��9g΢�Гy2UW�ۇK�c�oq
T)��Cu۬�"m�^�+��^Ć��6׽�Cteo���/j.6;A����a͜�)�˹^��$!�K��W�e�	�^p ���5�ZP~�?^����n��Ly�d=�qZ��Ͼp����[�����H�����̳���|�x��R�N�a��P�_����.�{~��H���]�>W�0$��)�}�Q"󣐘k�q���v��Yi\F�ꪪ"���t9�2��ç&Z�4+\u��	A�6?Q�G|�M��)�kHP4��:�lA=��J�sU�	́�� 딻l�>ռyC�6���uX���2B��ܱ�o�~��-�]����5��A�W��f�=K��;�f}8��娜Ϣ;��L�1�pΫ���٪�6> >�}�2蛾���~� cտ�׵����~��½�Č��ħ�W�Hۊ�B���uAC�.���`�D�s��r��&�7Kz�r�=j�f��õ�ܾ_Um~����#+t8ڣv���
��\�|{5�n��ӣ��&~��컲$]nN��4ltnk�U>kٝ!üq�1}3�$��}�5���Im���)�A�ݫ��SHȎ�d�:�3��]�f��.��V��*U�kՌ.�o����uoS|���.�bR3..þ�[W%'��Wď);h�� ��Fr��0��|+  �����iP*u�(�W�$̌��T�lGlz�����ݙ+D�������5��5ЮB{�Fo�'�Vr�6{N������$u|����K���o�.�N��
[��=j�(�� Myw�M��+��a�Ը��r��:'�{9���w}U<�Ʃ@��؃��o����nvOt�.P���3�K�~��n�0n�q��T��RZ���(|�/UD�]��+�"��qK����� _:���dz��
Z��=��]�����#Wf�9o\9^��s)@������=y��=�t�h�U��<�I DZ��'õ;�Gz�;C�a^������ǏR�z�1��v���D��{��P8nC��3�P��y��i>RE�D��Pܜ1t�^����9��=�i;a>�Ӈ'.�fS�s��&�T!��Q����ڊCLyg����9�}��k~�qA�^���t}�SM�M\��[�u|�/O���Y�D�C�I�gԔ�u(�F)�ǄJ>���bv��$���?Bܖ)ۼӜ�]���r�uϴ�9GE7)=ib�z�4��C�C{֮�&1�R1�ܨ+��w�w���w�w=҇�JN
5:��7�|���BV���h�?g��4-���ˡ�o��f�����b�|�~�(�4�^����G3�'8�Ģ<���|/�?OKC��O]��<�_^}줦�Z���\�[пg>T.;]@�[�X|�{&;u=�҈��J^��C��{F��]ީ�T=ދ�{Q��i���ʽ�<���A�Se�%?
��� ���ӆw}jd���'�YlӞi���|r�F�o*x!q��p���X��W�H��*����!Y�
��%�'~qq)�Hg|�����3�|Ow�N��T�]��OW@�>����1*l��מhg���u"䒽T*Ɏv���ݖ�2c��M"`H�:���5t�ڊ��Y�-�7���O��Y���t�a)���P}��9[����vpL]������)u~�'h�t7�&~��Wq�A���i^fGW�DjxDn��K��x�h��]a5[Ly�f8^��M	���l�u����I/c͙��uS�S��TڳWѷ��"������v��#|�s�&=��B���<����sǬ��~�O|���^+]����[�&�a�lۤ����a�FK�c�	}�휨y���m�+��pHU}7���6a�z1�Kޙ+7��gzz�װ[_�|��CCj�Cک��sQ����'}�Z��� b��0��O�Ҿ����"���1Q��S�3�i�e�xS]�r��a��ڭ!�o�����������l˥E����Q�P�SS��B����h�L�J-�K*"m�zX�R�u������ ��b���چ�\�7���T}�8�.z�5��7��"��)W�+��p�F�r�n\V�nx�)`Q�r�ד[i{�Ks��z�F)������`E��ؑ�}YQ�<�ȞO=l��c^�k!�%��J��w[��6�{��zsm=�-X��#,j��=\Gg/^bFD�����x8�o6��3�k�O���o���mǘ��U��_WٱEʟn���zx����NyEp��E�`�;#�k���P���*Q[
ky��܆Pf��1�8c��|�����b#Sч�Sd%S�Ə$Q�qRo�6s��_>8��t�*��*���������i�ﾁ۵���Yw�dտ)�`N>\㸻Kf�7�ד�ԗ���P�׵D�_��7�?)�Jb��N���kd�ey�����O����~�����&��wNS���� 6U� ��f�dF��a���U�%�A�Eȑ�b�;
E�O�����X����9�������$��wzT@�i��T�[R�Ak9NVoA�aݜ� U�7ۦ��f���F���H%��6W��%C�T�b��]����n�j��w_}�X��� ���|0ϝ��W3c�s��)w��=���s;�`���:�^6xZ0w����p�V��CdѬE�����Ճ$�󦽴ו��D^�F���Gs�g�(��.�
7����� ڃh�QHw�dk���G���DTeA���/��ȇL`�g�T��wgӕ�҆����u�Q5\�)�Po6��U^�2���1>k�����׊7'=���g(����팂 ��o�$n}�L����&_���ڮ	y߭����`�+��5�ݎއ���ng?+���/�����cʵ�1TOOAxח���d�+�������9�|�.�=Vv�*s�l��\
�꧓�(? >Tߠ�؊��9I}-n[�^K���M�z���������r�m�)+w�)����g"#���bV�`#�-�����K0����1��ƬW�Y2��k��)���=]�c��""����?���8�͹��gt}o��)P�Kܟ���w-�����I9� �E;��EW���U��ޕ�Kf�@�>����M4k�`���Y����9�����b;5�y���$v�����Y/jg$M�b�Ug`�7^�6E�RS�\�v��P����"aU.�q6H�yu��D��f7�M��w�)���F�&(�s� T涥F�gD6�r�#�2#hd��pܮ�-��b�
|<����=��=�\�ܵہj�����w�Ӗ���v�z��Zs{S7��eE��.��L%ك=�����Om�r�tav�h�P4�T���o�%w� h=����1J�|�y8�k�R��M�n{v8������j���W�ɁgC���&��/
�� �ud�W7B�N@o�P�Ŭ7���=���|4l�{� �H~v+��0	�0-��0#�e�
*Pr���;�����*�7�7��v���>m$�.7u���5�����O���-��4�9��(9��b]HƑ���c��W�t��#��]3%e�ez����v#%��R�d�@�3�m�tU���lr��[�Dz��&Y��͢�O�kއ_�K��ӿ�������a��nJq�/��dEy�Z�� ���3^R 3��Δ��T�����,�����k+���OL�~��k���z�,ԇ���L�2�]Ow��T{q��1�$����+�7b5����Qȃ^Ϋ��n�p�U�嵕������w���!�g!7=$M���y��g5�����v�r=U�X�!��~]�mUs��{j^.y_-����NN^�x`�yp�D_$9����|x|�쓷�{N���og(^/K���h��5`mJ�HGv6��_s�R�Է목�U���]�5�^�6���B��Z7���߷�o�AC��VJԐ�%bŐ�<�k���y�������s����B}r��k{q�������9���'��R�A�j^6CN
Uלkz�i��F�����ˢ�L��@�0���ARx|��b'�*��?�Y|*|�&�|��'��ޫ7s�d�[4�-���C�5Y�nA*�S�#a��v2skZ�_������ڏ>�p�Ҫ�k2���v�7�5u�&r��,�|GfTG��V�\J[R�Ӱ��QN�6�+G��y����������&2o*Ϙa �Q��{����Q"~eH9ݵ��3�ס������}�󼊧\0m˿T�0����}����dZ*�sxU�[�L�e��T#���J�e�'����$_����T3<Ӯ��y�s<�F�O=�+lA�P����G�ǟ
�OWUN���#P�~�7ಔ��%���m�|F�B�5���.�k������ܽ���w��(1�PI |O�I}w�U��'isў����}cegU�^&�)�����ֺ%e�Ϊޱ�eɊ�9��R�"q�ʐ��v�]$qe�!4�,��V�|Lִ�<<�=���t�]Ă�w�R�>���^�v��1Mߧ��:�4Jdy)�^r�Y�*9���f��Z����ZF����1<q��O  ��Z�vȤ�j���u���V6JE���*�"��-*�ʉ��]�t���s�圫���|���o4�̨�]�G%��E�a�����-򼶨����P��x�F%TF�Ak���L!?RF�>wբ0Z�:�n �J]w�|vUbB&0J5{�Oll�j)������Dw=�`�G��ۖ�>8�a!y������Z�أ3}�w�M�KѢ2����zB﷘�s���k�GB�o7���^���oj��X�G��x,'&�z�"ϯŞy�q���R�	O���l+>ؘ�ZmNn��X�ݮ
��LѯV�'Ne8tv����0��tbBV�����ٵ���?s\a	�$~���=�j#С`C�|õ4��n_o�����a��g��W3�6`�3�u��.��{���.��Nb���iG�� �q�m����O�,�}�&>��Z�ظ9�Lvo��+v��^�Nuv��k�.��k)�Bؘ~�8�M[��䌎����N.�[��z��>����Qށ��&�Uv��,yGs ��ַz�s0��>���z��+d�w�����q��\�,m��F�?C�ʳ�:�����"����ٛD�1�u�Bq�15^�"�u�v|K��ka?0��'������ Y��ty���G�W({�ޘ���iv�K��j�'����PU�]���x�[�Fj����;��E�7J����}a��^��/����rDJsm��
��۴�!��tt�A�u�5ϸw0´5j��Zf�\իoV��;s�cq��q���f_G�{���Y��3o=����b��l��߼]_�x�N.�R늜7-]��~C�bc/ӥ>�[2g����'a��s{���b�1׎i����ym��@<�E!��_���D�|a�T��5�������,I�?�����yX�oXi��1�����G*�*W�V.�9��;'��lN���t;��U�f�oVHE-��	0���.��i՜��s�K$�Z�y{�)1�������H\v�kg�8c�zz���{��N��x/)G�'�P�wgK�V��S�m��y���_N�V�¢=f�/%L��G�G´��������z��ѷ�5n����G�H��v�Y�KK�=�#�gʽ	�aG(�!�e��'�C�
b2N��#6Kg;;�'������j��A��>W~݉�{��D��0���]p�>��l�-�gi7.v>;� �s^�4���YCvQ���9���)��5�l��ڋf&��3���_EG�gU4���Ńe����n�����@�w�~�|s�S����(�oD���3��CQW:F��#j���U������l���%�q\5���K��!���P�gi�����<�h�)U
�!��h��ރ.�v�]!�ؖ���0!9\�� �j:I|Ys��3��[(�s����ыަ�0kN\�����Ҍ౉�(YJ�n,���y����H���^��OϾ׿�uu4]�v��:��DW�|�N(�כ�{v�aw�C��RA�N*�}�7��g��WA�/���"�YP��x��N�클&=�4M`d$�i�i����J��)9޺���'bw.���ݹ�}�����B{�֬Mۙ�����!w����̹��g�:�`;��Bw.��Q����5�G�<���k�f[��nS��U�:[E����>�l���O̎3��o�(��3�^S�f/�!LoC;5z&_3{j:8���/c&F��k3d�����x��jj���1�y�ў��=[�D�X�p�mB��l�3�&��N��:+/�`��ܝ<�:��!���S'�p�]n14z1��G�ͧ�L��*�ح}qn��c6���SF�n��g��9��=�Hg(��(����r04Z��ڃ;8񙺤��~\�^ǰ���r=�����-�������>�L��1c	�;�oDns^�,3n(�$���mԀ�в�Z<��Y��'��Io��\����ݼ�ޭ�v�B��R��W^�_M̷n�3Y��
0�J�OZ��JQ�9���^`CJ>���T�P��t܁u�,�ݮ|��x�-����>{hV[=: 0�]9�����Y����S,r�n	(��{���g��,P��)oT�5���;5��Y}��
�v��pp�.kŇ��[�a��X�Ru�ڶ�M���}�c�B'I��<7��쫪�xX�KX���0~�4�dL��hDw�4h+���Ku��Z��,$��a��#��B���do�>A3ZЄܘ��H�xF1���6b��Ӯ3i,�[Y��e�Y���6i��T�\�X���4�νV�[�AEn�z�s�=F���z�2���ν<�|z�٨��}W�t_=:�� ��V�Y�߭���M��޸y]}'Q�WY�1�h6y Vy���P���4S�ÅӴô�i��@� �ݬ��އ/uu�v	A�]#b����}ԟq�y�ns�͝7�7%t�N��mg��&�͒��Z�]E�<�3���t�nb��`�D�)��(��0`��˸���S�V���̽�#g:��:��q۠��Q}�ApnA�@ϸ?�|6�O�PA[zs��*��������/t���V�[���q�Pc�3��G�[��_�sL|0�V���SV@��oe� 2��� Jn�8�a	� �,)�$x�4U�� >'s�D��W�9�����zFl��ŕ�H���3�~I7�o�*���M�/�Ky=}]�Ck�f����
vQГ=�9�/g_=ZK�{ݽӁ��h�.�9KeJ��V�G3�c+;����shs	�Ko�k�\�1n��B�J�»bf9*u5{�ǯL��m;���wzp�Q��t��Vk'����rd.,�d��Y��H]<{��/�v��R"t�r�b�1���ޅ����ȌQ��FQF��n�.�����0�IX�g
��e��YN��!���9墕����8�{}�&8ؽ����L+�����7��U�
�.��@�V�j�n���66:0�n�*�D�~��+Ԩ��"̦�����'kܬ/�Vt#�\}Ep�J+-��;�����yYl��4s=���޷�u{>hQmr�YV���t:u^��Vn�g�K��&����*EX���6�����0kt�6��F�~[�U�\�[ks%k��p��Єy���Wr��Le��:Ô2�i��V��]6�r��l�2ofiA�y�?��t9����/��:�����"�[ڛ�^Z���F%Ϲ)+�M���S���J���6�����9�]q���Y����y-���I����q��Vk묌��N�v��q�>^kƚ�����E�Uv�5�1�o5�X��p�$˦�0N�	eevM*��i�=�2q�`!�~�U_�~�%�x��+���,��r�Yw��J�&'PTI�	�'}H@�H��C{���eK廹��kP�\o4'�I�c�=�I��e�9Q�5������M+_��޼�V2jڮ�|�k{3�X=N��V�*>r�Б�̪yu�ȣs�h�3�ŭ�M��b��k<��З��}�4U����=�WVf���Kw�0$�#S����G^1�\T����7�ݫε��G���+��GU^��1b_��}���c���u�ɮ�4�刨�������S�Tsòg�uz��o�=�Q���1�}r�
�a�G�����=�	F��8GnI�;�7�ȧ�7H����TĊݒ���T�~��5���q"�e����h)�9Ø����Mc����9�x^�~�QrP����y����Z�z:Gy]����1|̬���4g���:�Q]U7�G�]��¸\-U>O/�;���wk��&)+v#��)r����ſ�װ�r�M�%i��\���.5�fќ�ղ
����~��S�Eߥ}�̒�X/��%OT����劳�pυ�V%�Ll;w/�/D�;#�W�����'�l�K>�w�}q���>��1���D��(�9�����X��otu�]�f��|qr!��@ �{D�t���!��ɘ�0����-w�����I�6:���0��͐H;/a�dh<8�\�c ʷ�g�dVX�i\�5J�������|��������/dm��c��\����j�*ܼ����=�Q�����9`)o��Ʀ:u ��NAP���������'RI��}w�H?��hB�op��|�s���v�lR�y瘯*`�]������Ak<��+�;&Y�Rc��5zc���kD�ofa�����-e#5�H���;ayS����79Ft=��&��=�Iw����|����50h{� ,��<��$���ob$5�Ý�����D�-�;b�D��X�ݐ��O6 b�N���}y1��u0P��ٽ��O��6{��J�J� ��b>�|�z��eG�}�袬q�� ;J�u�ڙz)����:F�&��8��}]澿l��F�b�o�u�}h��m�ό$/�s-�y�6y=69w)�{h{Π9\�6Cv���8���n袧��l����{�v�p�P��<��$b��K�ig!Q�'��#����}ʨ8���.T�=;2�S�7>�'��e�#�^����t�ɉ��"o�H���[�<A_R���&�1�N4�-�L�;J���T�Xc�[76+*oa{����aq�������{�5�\������M����W;!K�-r�bh�<���H;%�o-��Or��ZAWM��7z��'��D!�\�[yۘ�t������`ܝ��n�yz&ѽQ����T�.�z7s��s
,���������9�XR�f
��M�:�O�,���M���D����\�;z����_����;5Z�%�7;f'3l����F��g�yʣ�[��X[BӘY�z���^`�&V3v*4��D���}SҖ�;Rt=�� b��`��m�j�s|���V-��T���p�|�ì�D�|<^�yhtI�8�~�g�V����$���3�0�۞1"�Z�����s]:~�s�jYCg)�GbO�qlǼ�>N8�Q�}��^o�{!��b�u�x����ݮ����2˾�c$�@`��MUmE�8q]�n&]ʠz87��G�����Z���@�V1W���������cf�U�.��&��9��{1z�K��F�����u{*$�m�e�2J��!��9����i>���U���	-�ޖ�ć���d��Mӥj�{T���Y�������`Wj�O���s�I�2���=��Gt��n�L�>ճ��m�z��F����U���+�&�3wylw������>���6�.ؾuy`�mgK#+7p2°C��,G���^
/\�췖�9��:��ev8૱w�{�&����vtn�PC/etxxl�^T���;����Z�8{�s��L����K�𷑚�Fz_\:ĩ�B!�v��(�ⶾ�� l��I  ��:ŴЛY]�Ox�3t�/\�b-_�(e0��v�l��@�Y]Sp��X�`]d}ǵX���vDd�:�\���~~sk�4ͳё�Ja}��~KƏ�>��az�����\O�>9G���7�� ���yu'Du;��x����WW�ﾩsr�:+�u��쪢��Ė C��?{��G/��$o�~����k��!U!�w:c��H��C�>����_�3�$}�$ooW�:/D_T�����_����ܽb������}�{�>/�Y;��=SeX+��F���ʸ�nc�z"V�z�6j�ȎLقe��醹�yH4zz1yܕf�.��5���j��&
E���1ԉ�^.d*W��$GW�MR��ަf����CȌ����1�zD��sỷƯ���̫�>� �X�ǈ���b���q��E�pz=|�����Qq�1r���{�'��ތb�v�4C�ؘ����'sCr�Q���^�h/5c�[�)�~��ӓv���h��퐩f�w{'p���*h�k�_�N9V�Ni�{�H�|�fV|5�]MiJnga�E�1��`:��5���{}�����u ��N.�G�с�;2�=�6��u7w�v���JJ�{�%��\=)��κ��;}Q���01; ��#�`P?#�1�p+����{R��ő�Np(n��U�q�Z�s�waq2��:a`������%��˺�g���A����7�7oưv�@@��ު�*�z�^b7I�}��T���,u\��8�1F����N�G��=�������1��VQ�=ǉ�-�^�Q�����:���|�m��������0-�D^N�+�I��_]:C��$G�zW[���/"��5U��
2n�"��߱�yu�o��R �{��?�8?2xl�h ا�@�ٛ!���W��|}o�s���yG����y���Y��&��٣�t�.���l�r*ܺ�i��v����f�"o�F���ʁ�9�3pt��Iܨr��J��W�t#ۏ�\���st�7D*)�F�n0��:0�nz'���XI�t������e�p���>Jz�F�bg�}�,��{�o6פzHq�r�%����ϊ��\V*4Y�/��|<~�jO�ƚ9+c`�+Gv��N�K��{�bS��z�%+oS9�C�Ȯ�	]�>�b���r^a'(ѻK��S�0�m��PØ;sL
-����!*x��Ad�9׽�6���Z�rY�S��2�YQr[�|p�X�L�nN�F�Ǳ+�|��fֵ�ՁW,�o�M=�� ���.�N?@sJ�^�^�;�!�<�M���~�^K�%�a]ѻj Tk�v��̤*�1�e���|��y�ӟ�~��"�<��h@��qz�f���j/�.���d��ʣ���l4hp��2{��l=��P�r26��������W��~7X��M���T �S�Kj�*��*b�ڙކ·�Q���N9=���A���:��"{ #|ۘ[>�F�b-{}�c)3�c�ޞ�J9ݽu�P�Vo-Y=8L�l8L5��p���R~dk}�u	��V���O���|"�h�f��w�{~��vW�nC� �c��&�%	q�܌c4_�d��Q�=u~腧�8蔶ѭ���]?b*ʫ��^���I��зL���dlNXmz;��N��6���7#)]ƃ��x�F�_���9ׂ�<���h}���o����X��/N����h�����^�
����"�E	�=��/��۳S��G�8�C{ފ4U(Af*�[Al?z'u��F\���w����gC�����Ֆ{�s�D8���+\M��"�q��A�SB�-/E�n��Þb�"Zb�QrM彗��f��0�H�^�@0�-�3z��4�Q5r��ڨ;z�a}�hԶZ�f��W>�z��w�6Q�/���#e/���Ầ��tA��s�t�kF��>�� ��X�s���W@�"�؝�З���F�h����W����B��rd5ƶ��YJ�'j�('��%N�)���ac=�z�\�H�mb�4��]�O̸�q�E�
Ʊ�G>��s٪^�12��0�lB�K���+���S�|v�7��� �QԦ���]�:�3�,��B�,V(5u��z2�ҝ���Ͼ¼=��')ES��+4�Wd����4����臛Pltz���]M"��߶ޠ���`��+��8j�c���b�:�G��C�}�Ğ.�ԏ���XW��|�~�⣔mzOh�A��<' �M<��.���WGȟ����O]�a!W���N��:�x����b�9n��r�c%F¸�Pbg0@���a����*�Z�XE/*Gb~���~��ϩv���?��yH(LϪ�^��>&����ɉ1հ��$X��8��1�53��oďU뾹}�y���06�K?�2�a��l���S�q�����+��]�,F�!|$�|�����)�amF�w����_ʕ��Љ�w�����PR�C+�K��Ӻ�N�c��1�CU�Q��nQ��ׇW&z �!/;QL��]�33����Wl�y��8��s��39�PL�}z/T[u֘�S�{z��@��[� �xʸ�fj������/Vr+!��}�z�C����8�H.�|��R�l���^�VT���EJ���p��/p5 ^�K�$���E�\�u�b��p�l8�BPDC5î�(�����2f\{׏&Q�t7T\;��Ӛٱ��|���qd��P'�o�'��b��:!���&��^��zx쓥z��^�^��va��aߖ�	�Z�#�	5ݰN�-�����:�R�X���'��gL���#���q��j!,���P����P����u�߂�lϟ�c${�G��	^���jR;�Q�~�|?㵦C_Q�w=c^Q�c�a�r׊��b�.���5�f1W{c����;��.����1�+%�P��*!�E�XyK�gI�`g���Id]_U����g�N����\���](���/z�����}
���*�b�v�@^�����}��r�D�&F椷��|�|��]6W���CKEm�~\��c���%���G<��Ƌ���w�G����=�%��:o_m�gB�Y/${����؟��;�O�7��ګ�5��-�"����sJ�+.���G��FK�"
�a�![׺,�77�RgF��.%YYr({���qBvJ�b!wMc�N}YN�y�U;�?,\ͼ��ﷳ�Z�7u�%y!8���{��}����s8UW������qj�8����ާ����tp]26c�L�}h�N�������y�|���^nK;d�����G����(�y�E�Ob�Z׳]5�zP1�;���騅x�S�BO|]�26�y�x��Ǐ{�d�S���y(�zx�ͅ.�R��ʈ,`Q��}?1�LA����P�v5�D�昱*b�~�Sz{��>��p]�I����,�ti{Tr�-��
�xZE��ޕEg�T0gD}�x�\����}�U7���[Ȍ���z��#�Z�]�X[�z--�;��3��M��$��ʩQY��8*e�%໭�쏜�nW��)!T0�Ü,��z�f���E�!�pw�v��~]f�qQ�){���$���~~�4:_[�"�7��jح����z` fE�7s�%����CK����yvV~{�w_�^	����g��7f\7�������9�>�jX!��)���m\i�/s:�>Y+��v��7�1x��]�rs��Et���+`]��b�i�t��3ָlɔ�+_EJ�pqb�Q.�|���TF���t;�����㕛�Gw ���H���oßU>�t�/K艁_u�8,+&�6��mn�bNq�q)v�p��7�4ٴ���v�x�t�嶋�Q�=zj�A��u��m��eE���6\`�|g��.�#̾�� ������;ՆiV���Z{cc.a���^�ytW��sk�jJ��^�.���^[�;�����+�o&,�p��d���'�3�V���lO�Ù��0��"�<�9,F��["����Y���G��Y��βMB�9|W�WX�V*����+����\��~���B{����}^�5a�N�6�J�v�(m��K�8�%���������0^�3v0�>��>վ��>�3ٮ9���7}<t�d�z=�=���;�3C�ni�`��4z�w��U%=�9��C{o��{���3L�%Ǵ\��.���nսj�r�0i��
b��y(����v����>'���dw��ίq*�$�ON�"��|L�U�b��T�0Øq�[tX:y^�U�Dd��텪.|2uGyG����9��hW{&"m:�M���O����;�o�;�4Ʌ3�}s��z���չ��(�}.��*=@����>�V��^YD��m��S�-h�9^��=�.?0c�|kG�[���vJ���#��$���WJ�B��	��rJ�L����@	+��vˎ��5�"o�&r�����������>�9�ܫ�:v�n�o��e�����Z@/��6$v�.��w�X�p;F���\c�<H�놫�zh�.�]$�c΂��>Ƈt�XN����5�m��(���;�X���)cF%��oe��e�<)~O�'�j-�X������{��j�;�3n��ڐ��A
=��Kn>�7�E��ZG���I{AN�
qD�B2�M6�XE}���'I�n��Ӊ���1�:VIi$'�ya'X		����]HO���,�T�7)ƽM0̼��<��^34����ĒM�θ�(��Z�t�6��	�S�Rc�n��Ӻ��]=�2�nBu��P�d��nkZs;���5y��=~��6���X+�]φ�� ]�f�S�NSc���s^xR��a#I��q�o�JL�  �I�!e�&�`�Us�U�sĩz�����ϘԸ�S�_�ϵ���;���I�ͦ����@X V@6�<�=���>|����4/������=�d���G�,/~��l���<sၦM��{|��;��H��0K�Z�X{ە��^�x����t�[�r߮|͋�6|{�`Bd �c��s���,����a!��{��*>am�'̓�\H�$�>�Yh:��p�>��!Zg���0x{����n�s�Y�-ނ�LI�o��ڼOv��	9���e��W-�>���&j�N8��CO��.�������c����a#��z��f�B:B>u2�1�H�O����M3�s�������|�0�@�4�<��fP�B@�	 �fe�������.x�v�{۶��K�Ш�+��^R�y5;׳m�0�N�:�NP��
�*�!�#�¥
2�ơ�}R؁-$FD)�J#۪��~x�(/wv�3�_Qk���i�T6���߳]t�9h�QT�>ES.1 ��Y�a`�B4L�������-���Nb�^4���f�r�d��/�����oM����Rx�u�������z��r��ޒ�t��HE\��=�Z��'z�R_d�vJ��83g^AWWcj�Ǎ��+>]�oM�c�4�=�6�6>����45u�M}H��]�\���Rj}cF���Ŝ�������u'�؊��`����d����6���藒:k;��A�.(��i�	�7#{��Or��B��8��
�t��a�M�DT�@7Y��$�����	�h'��/�K��b�U��p�W��꯹���p
s����.P�)��x%ڮv��[�p�����;�.�%�m�H�����&O�gq�ס�H���w�d�:ð��ۀ��u��.�M���Z���Ezpu��1u�Q՜�3Ub��C��]� �E�3%�[�A,�>��;*�3΋����z�t������[X��R� ����rʏR�FoQo_b9y��[���.|?&�l�V��^X,[��\X�tE^�iG�%�I��&���u���K�%�[��s#�9]&\�����R�)}��賌���@E�����2����N.�0��됖��r�2V����,�ܧ]�e�ظ&���)Ȍ�!�9�|���ԯ��뱝�|��n踁P��%	m���F��.%oD�9{ ο}U�}_6�{�i���=܈�/�sw�������w���Y�m���vi���]���WuG՛r�-�u�oVPC�9ۓxf�]Q;�[<\L���t�_�DA/,���4�8<�ޜ�f�j����+}`�Z��|q�xs톴_ȋ�����	��8�kՊ��(''p�hsx>ܼ��0��\�Kkrwn�����ϞS�'�&n���x�X�$ד�O�\#��A�K�����9�|�s7�g�����T���W�6�}��e_��eE�=���(Nq��
��X�X�3���iܸ.�9|�Lv��`2�sk����I5V
��Šǵ�D�S�����LbV�b�)|=i^a��!��e��X_ߧ�kHL#����sG��0nW|>���,:�͙ڎ]hm�l�xϻ��>�>�3�5���+鮌A��WQDH=�j0��Z�86<r�#A�Ekʦ����(]_�Q�վ�m�}��vկuRq��];�Q>k���h=�=fz��4�p��&m_U���	�o��鞁X�x/�`]mz*����
N>�{��^���9�,\V;�WMu�1{^~n)4=�_�1��<�l�-��U���;�����+�����owP��.;in��%��R3��Sr�Wg
�f0�dJ��e_MWU�R�U\�,�E�؜5%�ɷz�u��y�3Rjwv-�X��A�R�񩉜��c�ݍ={�9��<��4z��3@6$\[f�^��ҥ?^w�kT�׉�⮩���L,Ky"�7�Aꌴ6�i�y̔\O�t�䂹�Y�kx�N�8��v�5�#�5
.����Di���{�7Kd��x�O���՗(r�Ob3pT
�Y����OQ��4l�>Z��nm{GVK
��Q�|b�OT�n���(lL��x{O,g�~?x~�ث�������r�v��x�9���Ⱦ���3!�t6~�N?-&)���	ҿ/Ș�dD2�r����:N�6������j��P�q6��dp�ó���/t)���X)�>�<�<f���>��8\�^���T�j�Xo�=�As^��z������"܇��}�S�>�#�!w*zW42�/��3x���@���s9(Jb��<��w�.C�+Zs�c�+כ<LrDꮖ!�Ɉ���7�^��eW�x��c]�*��G^�"�Y�d<s��r�R<��j�L�Q�n�޷���U��Sp��d�u�R$����tϳH۬;HF������z�������ҟg:ԯ���߻���{Ѐ�{�m�kěI+��޷~�x���#���χy�k�w����vC�V����� �Hx�����6��6�ێP��<��Z�A�v�#3��;���撹���M0�=j��z�&T����oNʰrf�t�����5�s��@�7�JÉ��RV{˾�Fv�D�켮�ms�VHR��肽��zj]�u3��� QS�4y�a��\1hKT���#W^�J.�Y�?c��
N�׃���lx�g�g�z���صhO��]���
k��n�ز�ޣ�눕9�ى�#���-l����*�*Ք=��1{�i�t��-|�����f/�w�E*��6�yE�"Dd���%��q��7!��������$jB/?.�J����X��N���Ռ�xb�F�:��\ݝ���FOMXD���:E	cz�v�����D��[�e�C�(�J�*`�:;�Μ�>�ּ�z5��g)�-�K@�,i[�Ұ���q�y9�&��SG��e�0Q�;��'ؚEv�_v��7�G"P«B��ft��ȞJN�W��8M����H��PG��w�uW���\F����'����p�җ�
�Q���׬�&����f����~נ�����6�����r���3�t��eփq�>��>c��ꘂ�J�EX^׭\��d�}J��]I��ޥ[�,����s9����w{y,���E$�!��=�g��|7����o�vԽ7���TWN�;;"��-:�8�;�G���;�sv�;�r���䮺<	*��1i:���/���j�9�99�u�yi��1�$�sP:���e��t������:-*Y�~�~�]lB�w���g��D �˟k�I$ł:��<<����t�V�N��z!�3R����-�ܿٙ�j�W�Y|�Ƒ�/}T��oum���0�(��8�|f���������I�I�(`>���]����A{�Fo� �z��5���w��Z��꽳RQ�S|�T燺��qzG�{:*��9�97�V_e����Nq�*LȆ�uH���Ũy���ƻ�%Z��{.P����}���`u��Z�T�kg���s>����]kD3����kct��Z79�67!T���)��]�cez��@�-!����ڎ�N�Qh�I�4�G�KU�fK�/b{�5�v0T��P^��q��2<�Gz7N'}�TUGo��T����{�C�E�����W2�����9���f)�j��|6���g����-�Hů1�k�e��}[�Y�n��
�T΅s$>S��P��\���V�|�����'�G���5جD�ݬw�� �8,��s���`��kw�Wd`����Yjd�F�2�C��#�"�2 �����Ͻ�W�w��#��z�wqB��7F�#Pv��)o+X�Y��r���<�%%*ޓ��2'.��j��D�t�?��?h}B�4�%�)�� ���O�er�����Þu�k�ԙ�Yv}��?�����OQ�&=£�^Z�GP���k�eɃ�x�{b����~��>=#�7�^��Wt��򳔟-P|��\B���7��<���[�T���'�QΜ�h����q��`<�.g�q��q�{2�r��;-�����g�7r�kQ�w�w@��EϥU�z��G�k����W'R6�����9D�ki
e�]�>��G��(��n�}�=�ذ��L�9�F�נH�^f`^�5�TMIHV�uŘ)%�|q�!��o)�tU��-B�7�ke P��P�L���8]�+�TS�B��u�^��q����>k�
��d��%�/��\���`q�զ捜�qt��ٶ������"��]���n���D\c:�4*R�_G6��To�dW��jl��FAێ��� �Gc�'�'�j�>�+ڨR������U���Fޘ���2w=�V�+�~-T���+��	=�]�cH^�]Ȑ��=-��>[6�+?��h����鴞Pn��ۅ�ـP�aU-w<8��1<���PIxܕ&��qj�x�;�������j���p���N�y��f�Mt�8>��%Im�x3;���خ�����A,=\~��V{Fq'g������L�w��o������a��vnF_���P��:(�!-����t��'�"ߟ�vz.�39��r�^��Q�T3�N\ԛ��I�ut���У탢�;ҝT�4���y+�рg�
�\f�~?`ɟ C?�����D�帴��3z����jj�U��Ϲ���K���'h����X>֩�`������ű�FͲG��Cqr�nm�b�1"�}�/�'�������]�ܻ�r�D%ན0s
�>����{5\Y�ж�eޙ��۽��p#"�"��眩���#�?X"�^ػ���.�Y�6��*�A�Qo�2��lt�5zb�A�<���:�\s��<�d��]T��������Gp�H�L��=��R��+�^:��9ܡr3N�D�g�b��~�����sK3".�`�>������j�b�:'C����,�g��C�!e�^,�𽍰��r��1�3�d�׹29�r:,Ǖ�����{�	�ɏu�q������UȇI¥9�&��\���ۺ��(�7�����P�^Č�K#*(�[ �TJ�x�a�����ك��x�*�����������K�U�v-�V7��˧mg3�2f���uүo(���W"�n��fWv���$�I��~�1~�V�#\���ś����E.R���L�׀���B.��TF�>�8��#��]=̯f��b�c�}����$��{��?��.�q��~�x��.�9��i.�>x�����"��G���ƣk��)�y�Y6C���xlJ1B� M����=і��g��E��]><pՏ^�&�Q�i�B"�5l%cW���a�۽�S���W��ۛ���z�K��ϼ�¦u�Y���P5.�?y�N�����}>��37w>�u���DU|�Lq+|m�qTm9K�Uጇ}r���gY3>���Ft�P���+���frl�Qdߊ�٪�\׫{��_��-G��Ӂo��]��tr�^Bĵ9ָ�A>�\��ó��`�FJ���8=��@�X�T�'L��1��ixJ�����ɟF��[s[y2�_dgm�z:#�N�C�Ё�A�ȯ���A���l���ueJ-e�8���첇�M��;A@�=owE7����&̫�s��j��jG-s"�=eu��H��ƈ38�VPHq��L����s��K�Gu
��|�8����c�q��`ᅏQ�2�rM��b$���v�9�\�V�.��=7tq�Aɞ�b��ծ�� ��Ɍ��D͞���\{
��_ӧm��6�m�Z��LOs�QT�������WZgb��F���>5��C�k�c�T#�ꈹ{鑕�r`j;�}P���O�r�7ԑ���j����c�cG�$�ƥ2i�ř9�՗�>~�<�(��9����s=��';ƾ���t�Y/��A���'9��������[~�����kj��>w�0�J1��(�WG�m�3R�FEO�e��G�����u�A�C�?9��+<��T\�]mz�׋=���zۏ��_]�_)�.���y�M�
�1���z������힡��"&�/3��dtcߣc+�y�{���sI�A��;��ñ��"�v���~��/�;şN�
���s4���el�V �߁����D1�5]�C����&�M��'Z��ӷ!�N(T�V74�����,w1��`֤�8Ŝ�(���������缥np{x�r��ྩ�Y�d�d�H!�m�n.���]D�/E���۴��ts�;�'�5�{�q!Y�����}�tOK<�h�o�G!q�:c� ��]�~�f�ˮg�t�m�����x\\3M�_��\��D�\��}��8+ՠ�;��7�7n����N�V�`�ǜ��W^�8����o�Qs���*NXi�:�:�}����4�/�������r�gU��~��Oy����;Bn�i�>��hZȞ{Kx{��'��
���u���]{�w��;����F5���s�����P�e�e!�#jA98s��Z��s�i4{f
�"�J�C�
s�~�������O�ѳ��G}�r����~�%^@�t�==>�v��Ua54��]2,wE`�{�ql��`]�������9��KN{���T���1��u�u���Ũ�+�uv�3�<��vJ#��3�BU��.�:da��$=n�'ym7=P�2��h�3OGv�%���V9�B�����B�l���Juʭ��X��*�}�opHP�~��W�e&:�fXy��:�`[[5��:�<���p̀u)���;{ں�r5u>fZ�
#��'n��4�bWc�1e	g#	��#����]�\3=	cJlj5�_w�;k޳r�{DV���Daŋ�=Y��8<7������|��|*�3>1z��*�>��T��.]l��4�N���}02i��	C�#�Nm�۾�?ckݰSSJ�:���C��8#����O�+�{��&�̹89ߪ�n�E	s��e�B*�~]�Z����IO�/20Z/�S<r�;�}�z���q��������27�G�}�YS����٭�{���Deeo����P�Q��[��:�[�o$ma���D�+����g��y�.G(c�c
'�ZJQ0�k�=�*�sڼ`�}!��,m\b7��Vp��y��&.d==S*=S��~��	�4F��}�:�dq�r����0~�|^�~��2�]���{��?�ߦ�Dפu���E�?�c��\u��y���n�jE��;��;D�9��MFx�#�Z&���.��L����6�.�l�cfM�7���$���& ��{�4zXL�Z���w�?eE�|���'�E'��`�f�ſSDCz�<vc�%��}j*s
겹�*CJ]t�5���G�dwWta���x��;[�e���IL��N"�U�j�k΋���q��<(Y���<�#I�j�#]XR�&�sKy]��HC"�s �/m���x`/B/ �a���&/\Q�16����!��K�|H�\�R���L�m��l�:�|����n�>`@�d��	5����2��cFG�����L���znw��Y�9.o>޵��$6ì��@�xd���L�odYϟۆwG6�op]-�7���x��<8�Zu�`%{��h X�Ko	}�yr	�����=�<�i���a��$ ۂdT0M���2�uz�7"����6𓚦|s��L�o�~p�6����w�h]��1���_�i˖(.���絹.��^���+4�ݎ�UTTG����gӴф]�m�<���ja�ݛ�䒤�!�\Ϯ�������Ú�3�{�-Mj�K��s�nd���ێx01f��[l���my���4�<|a�ܱ=�����܁��.�Calvs�y՞Yiu{���>�k���C]��.�߮��a��{�`	�g�1�r���O��-1��>#б��	��� �~�[�����	�Sa�����9f!���_#CD�Q	��) F
����hۺ�RbXӁC� �!�zӚ�q�s��q��)rb��"��ˎ)gr�b�Um�Q�֠�9c��P�(����|�ɰkL�|����5ۼZ�̸��̑�(��f���{y���M�TkJ~�:wUkS2#s"�n�5x��;����P��&d9I�1],����x�vŎzİ,.�g��<�����t1`\����8NR	�'n�Yҧ�V��Ec���l��"0Mݍ	�x���4�����!�͒|�O~���/
�ϙ_Qat\M]+تz�������i�'N�]Ũt.�t�싷���G��z�']SG*�<���y�pm�.�ܱvNˮW0�-��p�qUt�Y�q.5uC`�N!]S��C�o�Xe\'+_]��NiZ�%Qq�����t';N�R�H6�)]�B��m���[B�--�D�e����8����d]�|އ}vD�EJ#�Zo�n��qJ���ח8;�W1�P%i`\h�:�p�D�%��\�����:�P� ]�5[vOb�[2�s�i#ԃ=:xc�5�s6�>ksXv�mxt#��'X�cQ�ҰuξM`�31�R��;���`��|IXX�]:u���k�ajن�goMLe��G:��!k�c6�,{x����<�r�o���h�ˢuf�m@M��tt^�V���ʍ=�N��ko�ǡs�zyWH��u�+���f��SXt�(���1�We�B��f�&�A�=g*R��3y�Z�X�V��+y�u�$�s�fd"�\�%���tFaD�X�rsN�=��_s��w����$N9����~�Սywuo�I�w���fdrԮZ�9B��r�N��Eh��`}Y�%w!u�Q�K�G+��Jk�Ǘ�6���O�2��Eo}��QǮl�H1�~����U�z(�$�N�v����uě�u��u-�͜�m[��F�O$�>�~�A!��?U__�&�lK���7>����3Oe<�8���UW��b����_��'dM� |��}��C��w��AC�9���}]=�>U�Cab�ъ��W�O���J|��I��� ����wwFɌ�ޛ���_���Q=����7��������?�ݭz���Ƽi]N��UϲZ����/�d�^ԽTlp�w`P�r#��PC����G�a��}�ȯmn�:��dOBZ)��\��M��秉,�"R��Z�����#Υ�W�{uwPu�F���\#�/��!
H4^��ӆzI�^->��U�;����}{�+�B6�W��>�"#Xكt��a�<K��y�jfx�if�����f�߀�����y7���I�YΒ��m{N�ϒr��ݹ�� OȈ�.Z�ՔV�V�Kd}���L�T+�9y�u.�r��␂ ��J�v�:Ƈp�P}rS�Yϙ|��X�m_D9M/kAO��;3��WF���obr])u�W�O�	^���߿����\�6�|�,�nW�+�y�����x/^���t#��Ӆ�M��&�]�ُ���#d���I��iE�4{�$��ŕ��q�@��;;���N_-�Ŵ�n��qש��]6�gP���0c�-{��ar�+/��鏆�s&�Ϣ�~��@�\�Yַ���q�w�9VtP�[�s{[�fu]Y���&�%�Uq.�,X�w��\����u��dG{&�^���>gx����׆�A8۾�U׮�Xp�vd�ȹ��/��1�Y�~~���<-"�
|yP�/r�����3����Լp�w �| �>����o���م ��ܫ}9NQ��&�D'�e=��ۈS��SJ��=�1�+낽Z5�3�]Xrqh^���Fl�/��2 f�[�'�u�갣�R�h���J�|��AI���yzc����/��;⥴+��1{��}��	toٷ�%zp�h���<Ï�b�^*�q#�k�ol�x۝;��ʏ.����:Ʃ1�����m�5��k'��9���q=�#����S=�Bk�7Ilg�9n2ʺD���iWL�ʑ|v���n��CD�k�ɱ]��ԙ����|�u�����!+�sS�������bz�܉�yB6�ѐ��S�z|��y3��)�4��-]�̥�;P+|����O���u�$n"s��ã���A��\"�bi�������Gwfg�]A_ftoh�����X������L�m��7����}�:��${��G�������D6��mw���j���=��:�X#�<(Z~����&q�g{:��'�;�:�4�z{p�0����9ٍrT�t��H6=�-v���K�����+=/7����Q7lH,�6u�����{X�Dd?g��q�_��s��v���,/F��>D-�= �%�(��3+�TCC�����Si!�3�	条���y�;H�jKX�̡O����0a:��"B�O�{��w��;��ci���}W�_ 4r�Y� ��Ǜ��ʱ]�-�BCQՒ�us1��խ���-.���{4�q���fKo:$��ս��"�����WƠ؈�>Ԭ���rg���_Lk�Y��}��U���x~x�T]��\��`ݽ�u��x鮶�FA�'�ޯ��������ܗ�-.5{�\�&{чl2m�k� �!>��KֵϜ�k�v!z�{�>��g�у��ufgFA�z��U��G�(�#�u��Z���-#՞@~�oz����jS�t5��f׌�:1�H�P�^O�A��>B}�$�h��w��<�g��3{b8Wp[�b���f�&Tsw��9o>��$���;U���~���uwW��=�/�rZ�v��MB+4�j+c��2�;�����s{���܉��wr���T��EB|5o����c�3�����ӞKݯw^*�H����u�V6c��.������R�&k�0W�PVt�{c{���I��7�h�=���ĉ�o��<����ڒ�R���]d�w��q���t�'f�C%c� m�����kageǋ���s�grn��qV]�8{�S�g�L�*��"�ܳ�����s:�qY�Si�=�
������Y0I�z�v�ֈ�?�힧��9��
��۶��~�~�^��7���M�S����(W��?>���e�I� ��P��/�%knÙ�
�s}݂c�VO�����~>�dA}����X��(�֨ʗ��~�9x�u�؛��"g��~���z,��U�C��/.�z��|^zVg�*|D*������n��R�'H/�l���e�tw�6�ez�[��4�Yș�#g�l:ҲP���X�}Ⱦ��:+-�6�꽞��v��W6���O�?3��RY�Gʎ������~�/
K���+�H�)6D�@�X�[R�1�Q�6���f]��>k���V灠�і���j�$�����4D^=]靺���UE;4�M����O/uS�y��T�i��"�dn��h;���$��Z�����vo����k��M�6gsg�塃7tJ>�����]�z?��
��.5�h����gu޵���~�$��*��� �'o]��&���=ϓ���<=�ݩ�1�Dˍ2C}�a�7�t���&�u��4i���e�s��D�vrĂ�ƧK���?{H�o1s^�"�˲n��tIg����h��c�kG?p��些�<��w�p�嶏:�=.b@ ��TUG޳�FX;~����;#/	⽺4�r��þ�ٺ�JM(�P̚�������;�hB[1���ML����������ƶ-�	{�<�~����?����M�z��|��^E/�����=Ύ�r�8<6v0�>��v@��93l����A�����=b��T��q��q��_��욨�Q�s��|J7��Di3�*R`���[��>��1s�"w�1*NƏO(�-��/2	]Y0���vV_.��̣݊t��>�l�t��b�a�L�J$�j�5��`��=vd�ؾ��ؘ�=D!�"��Q��t\:>��b�W�f&������@��;b�-�*KM�|i,�X�u�D���W��Ƈ�R���Co2른�Ȼ7Aܨ[��'=�ur��0!��כ��;���q�ז�����h��<<�s94qym��0�������u&R˨��Qȭ����]��hRu
�����k���C�K,jB:�'r��c7tȧ݂���)���u56w�X���>��U0;�Z7�km��~7��W��]���S��)���ua�\�\�6�s�;�yyD���y�Xn�c���{lL�Qdg�����h]sہ]QƋ/o��b&{�����9s�L��zu�����K >f�a��7��Ϯ:�8�r�Ã�S�y���Fs�=i�U�N3vUV7W���|�Qx�����(���n���t+ò�U�����S��!�>���ct�G�in��+��o;-�7/.<���*>���k8z�Fς��*�c[;�%���M1
q�5��aO�O7��շ��:�u'�w���n�߼�hϮf�(1c�6.ǎz�}UU̷���1c�A8��Z\Cg3P
Q|U�ӻ{�� ����u��PD�m�U�2�k^�`���sBtv/s85��!�r��n���D'E����2�]{v��]!��N��NrR���W����7K�5��3��}��>�fl���������^���<G�"_AiF	z!Nm^w������Լ|{�7�
���X�[��׶��hN�rَ��7��B$9���F�`%���-�T�f
�ۗ�U�.�T��V�P�� ���v��iV=�u9�����(t��5���3���7Q�>'෢w=4��&"�o��q�}˲���ͪ������@��4G��r!W�o����m,�kHg�pїOs?uX�}����n�_=���l�kZ�.�a�.��S]X
�}x'���ie�f�F�{�9��>�L�<a�O�W���5�����Xw�Z�l���NY�%,z��7]&E!�O:���_�f��]�����
�1bq���;r�.��G� �>H�d�^U$��
$��ڂM�9ut�.cܬz'����9��<5��]>T'���d��n	,�������˭g�p��d�C��Wg6�TX��I(����P�%�b�}��#ჩ)����������;���(��v̼/:f#���aÐ�w���B+���W��Eӗ-bӻ���Kzuc�n�{����;l���Fu�@��:��ٿz�}�^�O`��R��M_e���ʶ�����O����ժ�����y���xx�|�<�X!ͳ�,c�"�5��?>�o���=��|=M}�ҫ�)��sC��t�}Q�Ybw��\���}L̽���!���:��>������� c����j�9�w��xoN�mb�c���b�=�
UxG��wa�2c�O�=�7���D����� |{r�����'����TO�/���s.�\2�}v�k��E���w����]�3B�T�h}�ޙ�w�,�}��G�(VT.9jc;���姧�P�%5xY����B<���|؍3W�*к|.3z]^���v��L��=���u�퉄����\�f�{;�c���@9�/Gp�|6�S�3��s|�;�(&�Wvux��΂�D����mE涜^�ȵ�`��9��A"ø)`�>ۼs��Up���H6��S�ǫU����E���M��}�W(̙�����U��ANQ��n�BUL|�_�]��T�-��Z�\�b�7�B�M�a��
�\_c���;�:�pg1�x��=�j��^��b|9^h��炜^�����gk��gu�Ԫ9xј>ۃM���a��t��>��O?O[�����[UUH�Xr\WS�B*�9�1��歙B���=� 뜉�2.�_#G6=�*����"��]��d?#EE$�ht�ڬ5�pay
��P{���9t�'���+�M�v�&er�����V#K�y�T����w�^�g(�dV~`uHqs�U��Yܻl�;z}7d�,fG��"l��UѨl�UP2MUzJ��y�_c��ϼ��d.0���t{ܫ��=�b�r�))��w�m�v��붺'!i��{���m	��"���zx��=~f �(Y��w�y�R`�䧻E����C��s�"/�:�K%��$�^�[��】[���s��y>���K|�ж�g�(����yL�.nٻV�g �a��ٵ�_ �y��p-�o�5|�e]���]�7],ek�G�7P�e��'�ТwR8k�f���"�����#�����1p�[ڤ�hs�n��h�m1,v����K׹�3���J���׏VL^�ӽJ��SfF��\E5FkU�F{��f;��	�n8�rh��X�q�>7����c�~7���MbT��A(��Rt_r�2%%%�bA�3~XN{Qc�`!��Lɡ���}�����2δ+X�u�xU7C=8̨M^b&�@�����ʮ�k8d�6���-v>����5j�z�@�1]�.�Ǒ�/M���[�� �o�\�}Y+�g�^��R�jn�ugJXy�M�.Q&�1��#3zmwF�f����;ui喛2�0���Cl�E����.�(�귄$E/�)�f�|��J$���$j@�����m]����l������n��4��]���}��G��BW@Ɖ-����F���Vn�Yw7p���l5u��Tw{iʂ�`�5Cw/ʜ�
͂<���G�x��=�
* �J1�)g�	�1U�̹�O�����:��G����ﶿ�m�
H�M5���\��۾��ׅ6�n_��^�Dߨ���E5�w����q�uP�5�JńU"ņ�~�A�`����c�̶� � 5�Y%(������e�S�t�CLwY�ǖ�"�\�Y�U��ۜe^Tl���e!��uvC�]N��G�u֧8�(Ʀ��.yG[�|��h�\`�1�8�Ƀ^�ȱ�	���39�{ӂ��4)s�9a2����n��XT�J���)v�v�Z�$�4T'�����s�x��GiU�C�T;0�J��z�Y={8b��a��yN�P����+�<�ԹLy�J8�T�52vzzK7�uy)2�-��D��[j�9�W:W^����/���#�ÉP7Mm�]]�1�7
�#��U�2�}Jh�MX�5B��n�$��k���ʄ#4�ϵ�ðLɥ>�j��=E�ղ��b<��Z�dW2w��0����v@�[t���A�ѐYzV��:r�
��oU��ɮ�ݝ��Xԝ�RL�)���c�{�12H[ЖL��s��,s�n�N>X-:�]Eu	ǯ4�&m"{^�v�'a��M��^�o,N�H�oǷcc���b��A�Jf�x�M��'QS�u�M��}���ޞʋ"K�6.x�m�ݙ��0�S�%�y�k�6�Թ(e�F�dy�o�p���=�N�¸�Yi݌<��ne]n����?��sq�Hā�|��. !g�h�`�b���k/˯�[|o^r+���W7�ML��nH�g�:l=p���h�G��_:0dTA	�Qçu�5�p0I�M!*�rr�]s��!���{�m�wY�� �	z^�=S��q8UMX%X��q�̶��Z�9��ɣ� �"�䫆&V���\�a�I��9ߍm�Ͽ1ڴ���tMu����`"[[��&l�u-��ʫ�ȉ��6F��B�u�^��;r]��-������ٖ�y��駓�wGY���r�LTؑ�/�&��H�T���,-�ê��{:w�bq=�]��s��+�:�Ne{sg�.+߱�>s�^�|�絜��MK�*Q��}����w�Ԡ_���..��t���}*VU��P�����7��̲�Ms�1���M�i�q���,���v�)���t�3�3W4Ε^}�;��"������>���
���UB\Bz\WR��w�x��-uw������J�p�\����~�Zt�)�>���5k�*^�{��������[CO��$��B�/q�F�<&�B����%�9�h��4�Ǌ�O��z}8t�lݪ5�,j�������fpB�&��HΧ�5�A"q�CὭ���F�|�y�z-��)�d�����J&=��-���FgK�#��K#�g.ht�=�J��"�U�3n;��{�uv�wX&��d4���]��;#2~v�k��R��9����c��5�ܞ��-�_@YQWݱ�\D䵶t���n9�[�@��5�i����*��V*�d{��|3+��4�r��"���T<��7��ƤE�$��Z�~���s
�i����wQ��u��rփ;�w�)�f�:L����g�{;�����R�Aҟ�v�y����$뎳>���r�*���BT��G�1����������T��D��x�~���1F�J�<=	$�63�5c/���8�=[�=N[E1k�s6׎�[�n���j�<yM�Z�����P��F1]�O�۽��#D�ͺ�+Y�B7[���HƄ��{�t8��_w���o�}KC��XjB��t�ڮX0j�(��@u�7+¶��I�'�fG�£}�׽;~�0�ZY�������S��wg����� Z>w{��e3�y��w��^i<�I�xq��|�B�	c��4��Z�cHUY7���'����} ���Om#n�/:�c�q�Nz"q��(\�;_�2B��Nn�Rd�.����R_wf���,�`w#كi��"��#���c�W}�xQ�����V������:9���49�hJU���ݗu�ǰ��H���N�eǷ�{~�9������a�����G.l��\�v{1��O`^x>�
U�u�rOݯ��u_����)�u+N㽡�!�ݟTF��fOz360<�|�*7z5q(��Y�O�v���g�����{q����[SR��ϒiX"�˙�ۓ�o|�ϝ:I<�Iy$#���ו� r�9����;��M�@{�|͋�T��ġ�nfnz�-��t{�`�q���iyF��}���E�k����>�*�!�8��(��ޢ�����ùz��{����)��⣙VC��WL{%
��?���|�桉�.����]��]Jv�_�=��cU4>j��&����c����I^�6���߱g@;�o/���<z��1����uz� ²�T+��k�k���vCD}D ��+:�D��'R�ؘ�͡�N���e�6�Z3%���4��+R���r���<b��ج�B�Y}��U��t�\a3��ˋLx�d��E�Y��nT:��7���MKY鬮j��n�����t+��3�m��������h.�9g��{�^ �v�[�"��<���Y^��E�������(�ElYT�^��*��8r��[�k>�c��s&0�������Ww�$ �buMy�<vX� �5/1z+�Ec���^tfxZ;�evw19}+�v+�u+<}��$�����������rg��y�d��#�klGh��2�
�VN+s�ˉQv��
�c�=�)%��_Ƨ��f���ϲJ\�}k	��Y��o
ݽ�LT�z����x�����}�$R���/�}/���0�������+�ߣ;�cs�v�9g	���<�t{f�U���F&��<��v}aŶO�{������m{b�r�����MݙK�vYX購� h�9ׁb]N�A_T�1tPbP`F3�C�2.�tN���3+{��^��1�S�P[���}����u��oc�ۻ8�q�Zu�e�w����l�o]��?dC:�&���\��1��-��<�{���'#���<j�0�a�ݷ}\�a2į��B0�=27��F��������^P�L��8_��������/�H�QEF+>��xV=�E�}=ʧx��d�5�4�n8u�\���{�/e��瞋q�6�]���	xE\�TM����fI�[�f�竘�މ�����"�c: x��c�k9�Q�t�����4�ײ�}�;��3s�^�����l�������:}UQQ2CW;y�>�@}�u'��ɭ΁���-'6���=֏����`�Z���"3t���Y�]'sZO��8͂��c^]l�7�{Yg�g�۞�|lx{�+F��.1hdW�Ѓ�(�K�1��o&G�z#��<������;6�0߸W�73�E�qC�_x�:�H����]�Y�+u-�������sW���՞��XA���;ﻖ9����������#�"f�f�6m�o貙�X��s����PU�	�D}��!�ɯD�S����m�p��!��DBV0��d�}؀W��ӗ%$�t��l�y���vr�O�ꊸ�s��hg$a�{�l��c��0�w|v��y}=׾�#9�76�=�U+��s�Ȋ�ݳ�@���iQ��}C�e_��a�4'��p��n*��c2ڡ�df����:�ї�����g�ï�[��@��n���"J^8�{Edy�9���
�]ڞХw���S-���<��4�O݊�G>�6��z���[}�J�ח]]��8�ɨ6"�q.nm�����ծ�Ҷ$��Y�ݷ�RP��c���[��������:z]A�/PD����TGJ�Y\2��8w���}J�⊙����\�u/[>����bw�n���˞7]��9Y|W���mz(�����VX�T��ӥ��3[�(u|�ؾ��k�k����T�#��o���^�|1�_�֞-���)�����+*��g���9�E{��R�լ���ND�n����.�tϾ����&���b¤I���ӛ��������븘ݷ>v��U�6�f��`�״�]u5�a��A%Yc����bU�*A��k����`���]eޘ��ep�C�Z������e>GK/1c��!���V����Rs���>���W{:��y]5�{lV�:��q�=[R��D^Fz��=�<�w
sﯲf���TC[�{���ާ��X��8�"-uF�E�����p�0r+@"��T�)���*���/�%Z��γ`��5|y��P�wo��0=�;�:^��d�x�i�PH�g/ӕ9�\���4'L�w����b�.P:|n`�y�	��iܽS y��M=�j���[�V9f��m߮�_��Fw�g���A�RsP5����{���}'���õ��a��Ǿ���'ү����FM]2��Ѫ%l#=���i�?�UX�s>N����/.�制��}qPk�N�7�c���*��4��\�v��Bϥ�N�
���3SP��J��c���=�zjK��{c����m��o]�Taw��'~n�n-xVՅ�Z{w�~�c���R��ǅ&;*����C�F��r!����޳I�y{�4��X�<�_����n��u�xMv>�Xk)F]�R��ݏ�%�\��f�m��z�)a�𠕅u��[��*�~+��Z�m������}ޢ�����7ӌQ�Uϻ�׸��D8w����8r"2h>/�v~i��09ճ~�b�E1���X%	�A�2�y�C�r��몙_P�����2du�g�ZNI0z��_L������ؼpŹ�%D���7��N��'K=ݔeT��Ӷ%E����~9��ٳn�%��������bc���b��~�S���;��*��(ȧ{���؏��cWl�E�`�^�ٮ���`������%�м����Ow���q�_IC7�|�*g%�}e����'�5%C2,0D�Py*7{<��=��2<1'���T�I��so��ͥ�}�}[�p������� ��bqÜףǖ�M�~�l���C�kW\�2,b� ExfW& ���Ш�#λp�܁�e�qr�+=�Ǜ�-~�Q���+�}ݶ�D�ikh�����8А4���]�L��V$�
d1+�W��*o���_.�`����,9�i>m����Q���m�G�Y:��Վ҉�Y|�k={��\�έw�c����e�C(7�{��mG�8!��x�#y�*>ܹ�o��#uޔ�r����m��cMi�=B��&�|���=���c/����nT	�8s2�LQ��!�C����٢o�l����OO�1�ZnPz+�}�g�̱�Ov�Sꝋ�WWLO��x"�Be���=�6������n	���P���i�WAS�דӍo�K9�L�_?z���k�ɀ|lq?��dw�j|M�yx2�M	��>�������A�|��w�#Ƃ��:YY}�.d_�9�Q}wk��V �?a�tZwRe&v�Xc{�e�vc��}�]-��ۜ᤮���X��/|��V������]x�l���0�S@��z&鱞�©�B�]����9ُ^Թ}}'Ċ�wpLZ�U"�X�s9��M
��U̞9n�K�0�����^|�'�?|�����2	���F�E`82�b~��I ����Q����5ͫ���� �u�pcj�;WV�ވ>�E"��**�Ĭ#i�{xyX�M5}�s���7�4u��Fۨ�0�JY����7v7t�dx�ih+�K�yY�M�
���uu����[;޼�{��߉���
�aCT�i{ө�Zyn�m�g/ђՊ5�ev"|==��O���e�)o8�vi�-eا�m%����2�J����%?��q�t����zOod������T\�ȩ����?Na*�N̥�/�����{��OTf;
�U��P�2�����Y��ט<��u���Uo]oL�j<�4����G[��Wl���c𪼙=�;+1k,F��s�g��w�Y�)�J��5F2.M%�k�v�D{Ҿ�ZO���jx;wZ�9͌_S陴�~:�0[��.��w?V�un{Ϋӕ�<���:���)}��OV���In������OF�5�-��~��:��7��ȶ��wA���
\s(��|��j�{s�\;���Ӝ}%�/S����J�mp߲x�����n?V|�8B$��Ǝ[�Lr�B�?VMz���ϟ�������ճ)��ʡ�>N�@)䫅U�>�鲣��J=1b޾�B��R��O��x�%pV%5If55�6m��ށ��������V̺pef[�t7���YڧJ�D7��"���pf6����|c��QS�,����F!������,�]�m���b×���!�o��F�%O!��v_`l,}�-g�!x�w_�����&E�LBuΔM��}\�|i~���D�'A��.�qy˴5��'L���H��I�E|�B�\��C�G��k�� q+b!�W�49r�m��[���=���6��ݻ
N�+�u���!{�,�.��I��*��{�V�����,�ָ���i�ګ�d�K]�vV�w�� �6B��R��UnVOc;$4��l��fD����j���1:�_�v��P��{��r����+]��dh��?� ݶ�&亜{H��{}צǎ+��;o�_�+�AY\K)�W���Op����.����9�]H޼Y���ڵ�M��WF�v:�h��I�J��8��.Lެ�-&/�1S2ixʺ傭��jt�pi�@���ޤ��6A��=ᑒ��]3v@�Hv4쒶c%��D�x C з�ul��.g�iI�a`MDl�HpA�����1�o��7�aQys��1����Z�4-���+G������Au >!�H~�Bd�4�B�bvL�d�(�u"	�-Mθk\���,�ה�����>��+�gMu h]+�	W`܊���١�V&&ﲰJ8�q��eKY\�fJ�wD��
0Чw��Q�ҫs8s|~�,b�S��Û}�3n]�t_]�JJ�!�bEu;��0�T\sW]�.+�y+�YH]�N�=s2��(���u6�jS������ j����i��G���4��0�Tm�\�h"w9��.�YH�\��î�J&�JT�K�씭�[9d�ԚEZ<e��J�t!Ե�K�h��;�ԡ����^\��+��Y�pm<p�z�JY��5 ��	>�V�\�d�*�1K��A�#�8�n	�&:�^um�`���iH��Gq���e��E�mŁ��O.9ǭ�}�B� ��H��{˿+�n_v��Ҍ������®-/��xv�*D�	.��]qu�C�s��oo�G�iCj�\�à�Yx`�*<T��hw9EmZ˧|�%��W�Z���PY�Y��\�}w�9�*�u�QS��)�
�c]s��%s�Xʩr�枑b��,OK�-?t�d���B�z��X�VY�BsRA��V��4�P�Hn~;��[�PKȬ�r��A�+�̧-NӦ�W0m*{��]C\z���	3t<�MM�8�vwM⳹��dڦ
�,���8�h�5�J�����Ro[�@��N(��yv�;�uޑ�wn�;Z�BKs:��3Q���P��1����|w���j�����*��_}UUS/��rw�߱��m����R7��:���Z������Ny�ϛ�έm�P�Q>U"5a�w��_J��uq�S����H'�A�,��˶�'��W�z�����e�|��Om���{鯜����-�/��,z���p���a��=S��'+`����mgmg��̬ߟ:��b� f�_���Q���]Dx�\���'<˫�ͮ����uO8竒��<���e:��wd��0�l���8ϓ��]ѵ>'~��vq�������^�q5&�<����?}�noV���^[�S���}Npx�����k�n�!8��Mx����̿"=�_ni�p��M�\�Kѱb���b�V�D!>�qA�Ps��^��u[~ca��b�V���9_����}�֮��R�	qj#���2�̟w�ʬ���G�]��_��$����qWb�o䊵�����{S�9�J�ا{:�Q^�%��VV{�|���H3�׆��e�lN����l��+���$�s�07y�LdwJ�#aE�*U`�C�UV"�F+O���Ё��״h�λ�u�s��Pr��Z͍��m����O,oN�_57��&�o7v�]mYoPӶ'![���O8��=�N��kp��e�Ȇ:���T�:���{7i��n�'����G�V�wշ�:vj��;��>[�˅v]ݛ��]���{5w����	����=g���fľ�h�{�5�9ȨX�5�(W��۱{�]z�|d�TTFV���~���c������@B4T��U��'*/az,p����'g'E�s�{�o�ؾ���gw�m�?s�;�gC��Q�a�
y�uǻ��ӗ����
c���q�靇 ������>�i�0ϝMH��L׍�W�Mq�q�[���|>G�P�q�&	���=뉑T6��s-�a;4mT�d�q�3<tϡ����B��2�M�=9��uz��V�\E�c7!`?ulǈ~S�2i�j�H9Q�8��f��ڏ<�8B���<�����<��B�kއ�d@�,��%���pB;,�:��><��:��%v鿻����v('�V�I4.r�Ea���)R�֭ a���� �&�]�o��_f��:�u:���WV�&�o*B;����{78��.L#��+ zrva�tY/u��ٲ�fk��8�+�&�Dm�}%wF�;��m���Oüʁ>ta���<U��V~}ފ����U�A�J/Lwp�̾�RS���1�[��[��nuyVG�JE��O�2�{*b�m{��y��{�b_���c�tŵꜚ�b<J��GU�B�B��V�:7*Z�i����7&��wy�b����"+�z}�=
�:B�s��Z��ˆV9G�1��f���Z�=]���C�M�j����v���ފ-��^��t����
��k��%���E7��D싔a{�.n(Y��ºa&̄w}����l���8n]LWUu��F���w�lYz���yρ�fT���X�|�I��ى�{�]�a��6�� ��j��֫�����{חX/`"���`O�@����� ��~6�]��1�ST�'Eع�fiG{�7��\@8���T�OE�X��� fz~^�Z��Df�4k؊ �{�7x3O�uj[����������Q)���޲���g|������'�������c��j��U<oke+�[�3+���/��\�'l�&��aۯ���R�jGX���1t���ob��#�K�l3Zl�[��J���ӭ��17wo];suN������n�wV��_G�PC�!�'Z�<E\���d{]�2<�����p3����9�ܨ�O5�����B���|0��6"�� $�x`����ʠ�u+����xDFϏ���]Ґ.�j�<��8�g맇ޗ���,Gxl.`=��}^eL��Eg��@O���mr�y���mL�����><yh��x4�^�<�|�?������GzG����0�-�Ş/���)L�-"H��'J>�ȳ�ݳ�oO�œ�Z�sY�ǕVN��?V�o_���J ���z�]{��z;}������G�UM�x�T4r����ܠ�ڮ����%i�>�J�]� ����ה��U��Vw-��p��aLE����>��+�\�wR���l�:A�ߕ�{����vG�
(N����ۋ�ݙa���?h*���5뗳~���ʊ��xt<=
i]�U�\o*����C}1}���Q��
',A �o�����Co$�C7��Y��	�� ��K3�;x���d{%S����c|�=k�Oa�V=�G���d��n�
άj��U�ʔx�E�т^=΁�.��;���i��Kq[ޗ�lZ�:&��-W:���ǽ4���7w�$��Oj�[�Ӝ����CHQt�|���}þ�!g�IN��F�~���G��B��~��N�%#d��Ǆ*��L��r �}�=&�.b�p�kR�GU��|�e�ֵPM��$�r��GN�8�m<i�>ow���q��]D�.lF��큷�!�Mߥ�/��	�l���4���dx����!�fA�gV� }U�k������3U�X���Ŏ}��ulE�6��~X6���H�>��J�~���M���ʧ<����$X4V
���b�l������z�k�
�ӑ>r�LJm]1�<":&n��Ƒ�C���W���^�"�L.�d�뼓Ɠ3����"�{K��9�i�c+t�kAS��A,b�/|}�O�4�stz�����A�I,Hak���6g�/�$�.U�l]�Bb����	�*���溟S�����������t3і��Ј�;��둹�g:�U�L�����v&+�v�����z<�ĝK����	��kH��״dh�Q+}�f$o��H�k���q{R<�,��vs5�8?��D-!�O���֮��\2�uvv:�twLMD��m����>�@�
���:�k���CE`�[�ލ�(/�S�y�j��\)����Oq��KO^�<�6���u%N9]m�B�gZ�+��/��*��h�Cg��3@�e�T^���53��O����0�>kE��C��~��.Un���J�Ϥq���ʶ�����a�Vy�!di�i1/)���E`S��zЊ�j1 MG�K��~V`���XV��T�Y"qM�吴�a����0<��������M�v,�чB�6~>�=l�sn�9�ճ>f`+�q�e-ubjF��O�ݾ �ԋ��(S=�}pt�T��9��k�����1/C��q�J�dע~��Q�.-ml@�W�^W=z�=�6��Ͱ�C�^:M��:����w�����z��1O�k�/�>&�gxN�N z�h�� k���Ƌȼ:���֗�;��m�++��_mme}�I}_{�o��2γ����U[��~9����0����6��^�Fi�:�M�O"�~�}}Z�zI�0��D��4�늽�\��PI��U;}��Ǡ��]s��o�z]{hI�ˌA�1У�+��>�\��(��
:lG�n㣐*w3{�w�]{}�r�.����Ek����xo�n劕c[-�E���j�=]C�;e��K^�Ƣl'V�����״�L�<�{\��u���u&������cw5V��w7�pm���i�x��K«�ͽ��N�fۙ���GA����G������{��<�g���	yM�l���x�׆�`����L<s^�g��`(��%�s�g>Ze!�/�զ7��OrS.����m7p���\5���of��$LX��Uht���0��۲����Uazb�8,3���ޑ.�~�-�1��x!��ϭ	}�f��&.�=*v�=j�B�$�y�+�*���7�}{�bU��x�=['�����>�
�O� 诰g�7�A�݅-�܁:�]�X�n�A�b��Bf鋞��陑�`c��ޘ�Q�@��K����a����th�}r����?����F�Y����,�p������Z7�V�S����1�eF;v�#�h|��$-Q���q�y(�v��2�@�c���B6eO�n����b�H��|>�8^W7�p��j}������-^Ƀ�Jb�����wP{zcu�a8��B7��n��s�>5<b�-�T�N�9CU��ݦ=\f1uc��vyDC{��}up�H`��)�����}aQkAP���Ͷ��{w�@�j�Y[���jG/�WF�q_~/9�NBp���3��sW���P�=&�[|3�}	���*����o����ZI���6l�1���}��1����|��H��t�Hj�9����e�I�̸0�V���_Em�?Kt,�/�-��/W�f6HѴW�Ʈ쇈O� �{7 g�⥁ƪ=����r/)P<�	|��B�2c��F.Z���?,�����\�ek装U���F\�"{�F��=�MAb��;��_w��z��t>�w錛���&<�&�(�Ju�z"�X�nN��������I-��	�M��+���y��t}{���fzz-&g����틈�n*����`��m/��(l�O6�,W(�����mfF�������֗����>wu0���+H�˽]
MT��8�q?�Ď�����mo'�?#��9��ʯ��<��2�w4W�]0�ލ=Uޓ�bU>>��7Lu�v`�팯K5A�z��.�;�PlAi�����s}u�����Ύ�~�&��;�w
���D-����Ҋ�o�g`�;�?W�YC��v��mG7��&�+9�6��ۻӯ��3���lJ�X��,AU�Z�A9}����l�:��|�ڬ�\�X�v�)�!�:�[3���W��L�<���NA�5�X]�k�WU�l�|8˃`ki����f���G���bx7ja;_���3���B1���L��4�"P�yK�F�*{��=����G��.U$���!��`��}�N��#�X�\W�·F�y�	�J��s���DOT@ö������g�ˤQ#^�����0�3���:��@1��&���KWyK�^�o/��)㸔d�������|x.��n<�NI�V�)�iy�0~=�+lKRuItk��De��=,�ű�����d�<�:6�ͱ�e�������a��XՃs)5��|��6���a��.%t���~�xR�Ӆw+���˷�����2��sN)��Cv�T:��7a�ک��q��cn���Ȯ��ɹ�����`��g��)��P��
{:;�ŋ;��`��Y�p��ML�Br���Ӗ&]*y�?�&M�8of2S���P&���C�÷��%�ڛ�L���۪NL��r���nDhPCI�q5��y ��h�`���]�43wv�/�i��&�jp��q����5W4���b�?��.�Yy{#�.K���'ބ>�S�
�=]��a����nڥ������R<̗0H+Y{��|2�Gu8;]�Z�^:�:�Շ}aT��:����*�z�n�k�۸�^��Gm���/��|kw>J��>����W�F{T/�'f��]ę��"]n{ƴ�|>t^M�-T��؉���'�R��[�Y	o�/�f�,��F�ʜ��۲5v���ˣ�W�;ƣ�=sj{Q+Up_�;�]-��9C����Y���i{��ٺS��zG�����y\�n]ַ��gf.�tרj�=E����������7#J�rp`+�S[m��9ڰv����A[��k�L�W#��c��V֗����kw�{j=򗲫(@�1�^_lu/X�T���~"_����{"Fv�:�[F&����n��ڋ�b�VHu�j`{��w#:�y+ݾ�Җ���Wd�P_����H��̂E�ؑ��т��U}���b��[�No͙G��X..�!Wf��_'�w��+�Vh��듂�Q�dMk�}5(��j��&��zF�z	�W�|�͂;�4����K���/�[����@� B)��V��@�յ݀��t.�{���p���'\�W1��s,���g%�T��<�S�����ŵzGa��8jU�e"�):��#p���}�k���du�[��h�NS7$D�VW�P<�	ns�p�����>�wη�-9�څ��5	}���곗�
}�i���� ��a�����:�.����l�ٜf�ȳ*��{׬��R�	�s�[zC"�?0�r��.��P��>(5h�J�xZ͒��0�m�4��`����K��
��1�޶��i4b�����o����9Z�B#B�2��Vo�N�N�ή7�֜du�l7�Uu���z�,��Δ
S;joL�ݽ����}�F9��U��.g`�u��t�Y�zv�a�?�.��C�#�_e�N�׻����>f�(5�Gw~홮t��H�_i-t������+�v��V�N̓�n+�����,a���N�E]&{)T��fѻ�CLM��:�q�>�N�y�44T�&K'�A�JD������b��7�a��	[�W_c��[��v|�<s[L��S�2#�㮼�$�U1e��;�O���I�@��zU���]�غ��5�N�A�>�����#�4��J�
��,���%�� ���u�piL�����˭�g�AǤ]6*
�k�r�ց;%s`���B"&�1�4�2���{`��"�-�ex�/�8<��&b2�*TQ�Uq�\�e��+�{f�ۻfW2����(A$��/�-�����~�慧F�"�#�}�
�G��֨��ˮ�C/t�Z���+P���/J��-��lj�L|2�{t��j9&�龔����;ft����_u>%�+����k��˚�_t(1X�fah#�z��g64���� f���#�wN�%]��ra�9�����O_WX���tf
��G6]_�J���K��0q�[R^*4az�[e����%��}���]��|��t�uv<Dv�y*����g&��ҁ��5�tu�H@�@�|�9�C-�����)Ѯ{u�3�B�w �זd���NV�`�54ԫ���xIz`ھ�O� �塽C�e�W��so�E%%]��|�b�M����7��xi�֫ԙ��mѣ�c�LvN��Z�V8��ݻ\�wr"�;[�YƲr���ہ[3a?�����-��qb���]��D�	��s��VY[˞]m���
��:w�e%��f�j[��(puIz�s�M7\�pe�OHC��;{8]t��������/E�ukR;�pK�Ť�K���4���vu����c�G��q���!�]}�x�infTo��˷�鰲�%��<��ߖ9�4������6�a��J�`�#��c�D�S��}IVU��[�ҭ���eq��w8�&�����+V-� :���w�Au:�,nl^�tܼo4�i�;����UU��m枢�֔�O��`���0!x�ޭ���t���i��������C�2ћ1I�"[��P����2�����u��8����Xw�Z�Uu{��*Pn9� |�~��S%T�z��u���'~{0N*�R8exzEl}&�Zޯp��k}����x�Q��Q}�csФ��\w;0!q�vR�}0���KQ�H�ST��,�ĭy����T��/D�[�̫�"3���Xi]r�N�J�3�2q�ڥ��c�o#r.󒞈����i���L�;9��=�,���l�ll{z#t۫���xQ�x�����w���X>���L�ؘ�Mj�;��:��q$߮������pu���[�~���<��B]r3uǜ��z�3�#O�sg�=��^�5��E�b�LM+w:*�f�|c�s��O }K�|"�V׊�+֔Y�����$�lk�@���0b�����{j�د�M��]s����c�>�*2��w�+��Nyz���كg�m���	�u:�b�	i��_��(�~����m�V��ZXy!��#�z8��FV�xU�}f2"���&f{��,�I������=��^��nI�Gn2��]��� JMvR�$V��y�S��q+<�����n��/H���Y�M�`׏�o3���7�W'��կcȼ�����x1Z��]$�}���]�@��@�H�#�u��S��o���TǎV��}��q�9���MpOo���9�}=J72��}/�-�rȚ���R���l�o���+���m=�Y)�����@���q��q�k�P��El�5���|��E`�sZ��Z�uC��V���?�=�<|v��p{���K��U�[<��W�vι�}�vX�\��sf~|t��Ng�.P[�s��*�L/&[���R�>��mE(��nRkw�@�kY�t��2f���WW@�1�WRev�v�һ!����{c�IɥwqP"	�s�{���&:<��7~�qpw)/�d�,�k��P�Ǣ��ӒN�9�՛��!;lT �Xo���Q������$G�0�c��Ea�'#b����V��~�Rxϳ�{��(��]��=�{T�9F��X���S|cdx������P;m����R������h�"tu�:�azD_��=�=�f$��i��+�~���r�N���5Թ�v�f\N{�T�%���#���n���<,0�YXn��8
�N���(��b����˪���u��ȏ��R*�n�nY��p+-�[��+6`}�o�榦]n_÷�<[���x(���\�ֶdU����nq����ʚE��"ni_[B=oA�Ҝh=��Eq�YF�xΎ�ʳ\�؏w&����t�+�Iŭ�EG�9����8wX��]u�GE������$:��.�����T=�xb��>���X]3�[�f�����\j9Ca�ʩH��1:P!�k�W�������2'��R��16m(��cڵ��	"�1���1�=!��3oѫ�v�����S�K������7�4l���v{*Fs�۵d�T�V�Z���w��xO"�b}�F���^�|H��"�ft�����=�##b�r��\��G+l�r�5�ȯ>���ȫ�tY��q�\�/)��4z����\}�����\k6A�s����\ʅ���-{W�H�_bx��67%틙��*x0Έ���V.n7��cOk�����)�;�w��yw�����9�_��$���0b>��c\�q�$�P��Ք��T1�Ծ�3��v����#V��<�p����j�z"Gd�Q�r�ɤ2�L���;4+�*�NZ[3F5�����K�6)b@9��Wbb�Q���[��Dj�w�^�-�v�����s�ӈ�X��ubuc�T�>���G���!�͒�|r��}�%��f�yԯ��֕b_	C�VT�|T�_�g�#O�|��Z�e���{��=�dl~��&c*�tx;0-��zV
����/��[��P
�����=��N�QYpܰ�wlﳢ�	�K2}�� �%A�^(��43733�ä�e?S�Xφ��/ww��q:�0��@!�3�z|�6�7h��q����y�]pF�-�{Qa~;���>�������86T��9,�*��o(��Bۯ</qٮ��c��)�R���@��;@��ߌJ�A�أ������{b3���R�纛;��>��눷��P�$�� �"��\U\�1��Z��˷�7�nK�&*�M!������˅����[o�7�㇭�ޜ"tϨT�<�)���\�D����^�M��Ym������O��>=���Nn�����g�ei�ޚ��?x�d��6����]� �=}.c����� 
'y�;U7U��Y���"}��c�х�'�����\!؃�>�������k+���󶵨A���h:��C�1͡��TV�|f��u��^w������.6z����z��<��O�2��Cb��-��k�W�3���O+[�� _bgZq���a�?�xɿQ���p�擥���
���d��!�T�b��g~��g�����<m�m
��:��<y�{� ��N���uF^��y-�t�:��B�R��r	uw5jRs��\�Z����8��zW��4�P�����(��7T�zUvŇ��.��Y���B,���œ�*�79�m�N#  �}�܊ɉ�l�kl=�1���Zgy�g��1��i�:�h<;�^dak`�������Q�J������bڽ�J����߽C�V�N*K6iO{xt���6�e�EO!ʝ�	��՚��gdM�\�$iӘ�~�qi�T�:;a�J{b[�7�bZ��P���7���>� }�Ç��Q��J覗>7���>�4�5*�[\=�)4xT�m�O|���ν	{v6���r�mO��d�w�/8���X)��/��GJ�nf'��FZ�WYkj���ֵ��"��ܻ��������]*Y���i}w��㆐Hwt����v�.[�
����FI6e�7��颫z���_�����+'cݜq�f���B��n���;����NS�wHG��0�ݙ���4;
�Ȣ�F���_�i�*�4LvP��G�8��B������\��V��>)��)NS����ލ>]�"��3�7F��|^�döX�X1>��Wf��P29��QBT��ݜ;Ǣ�	��<g�� 4}�����ltFp�@��jָ���<o����0E��x��p137�A�fN�BHsT�6��^xC�x�Uyռ!�i��G�8�荌�@�����s��Ϧ�cʆ����*�'�BF-���`�}t{�竃�
��P�ӻ3�X�w�K�!(�������]X:{+o�T��P�"�y|��ޙ[���_fL w5��2�b�-��{�C��%�{���7i@�f�'q��3��\{�3ޡ�	����b�k�E�]wo�����d\�ǔ3��m���.!�tWk�����QNıQ�{ɑ 
<'/d�⽲}�*���ٓ������'�\:H��C�)f�y�'��]�����3�Ux��k�2��]	=t;RvXzP�j�*��7)<��=���^�{8�S�r�~J��T���m���]Z9t�����8	�W�8��#����7{����d�<zӥ�>S���͡'aY�S����ߢ�h��t�.��$�h��F�1���nY�C<��Xr��8�I��K�:��^��y�rUZ�DR���`�*KY����7ܺ��ܭ�-;]��kJ�gl������o}���1�om�{P��6�$x?R�I��G�N硃�;6�։�k���r$��sL���0�*��Q���Q�\�����s��p_X�rd�y��mV�;�^r�TdPܹ+��'���/J��1��c�'���x<>������z��jvC9P<}!�a��"{�AWz8�@��#�_:��(��REcۊuZ�zY�`T���UUT�.�3خ���ʠ}��^P$LT�խ.O��C�w��t]J��3�┇j�[�Zlxc���Q��!=?v�K��1o�w`c$�]��^��k�SR���v��K�1;3��*+I]#����V�Enw���4E33 ���x/>j�����OrӾ����{�M��CQ�D+8���o�: �PߩJ��=I
i�y�������4����Ty�v��]���k|�Z��
�)�Q��f�;Zg'P��59��Y�+���R�83�nI����8�6�o�o�h�wƖ�:��=�2Zo���֝�Q-?e�VT��?_��J_�:�;��m�����+��;A{�4wZ3�i츑q�7%��E��=����'y ����Do��,p�؝�Uz�4fŻ��x��r�^�$hY�0��w�.$z�3d�J�L�S\��W	oJK�q0�A��һ��UЯ�JK���9/�+�y{�>�j�"z�1۝�R��xϾ�_�ՙ')+����Y�x,�8�g��`���zG�W����Ww�{ׂk����t{$h�2v���Jv:��[nn	x)y7�i$M�Z��R�w��Q0.�;(lƥ_p�����_�A�ӽ���Uz�o҂5h����ϺV<�q���O��k�!Yڛ��N��栽��؇۶8Sꎵ}��N����)��� ����8[�C�+ީ���(�w�z�V�DX;/�u��v��s�x��8���u�1\da������x�Gʾ�Y�qq�V�ƞ�3\���Xę��w|�Ӄ�?{E��;����R�lxT�2�f�M�3E�I��
�Uq�+p�������*ͷf��7:%�zN���_���L��R�Q�{��8����P�B�+�2�l7{�wp����M��9Z�<�� �F��u�W�=�kgZ��(�R��1����R�8����U1�uzx\_�G�A��wB��NЬ}�ƹ�����|,�_����M�~��*��:��v�K ���m
���4t�{ޝ�P��l.�������|��6����>b�ư��XW����s�O�{<�9G��k.���{C�~�.�}�Wؾ��E��,�!�`���Y���	�;�;�:	�o]OP���������0|Ы{AL��1�Wyb���V83�^>3��	�> ��@G���z�*Pl��^�o�,��<����l����}E��Wρ�0%�.��ؘ��K-��a�S�8��w�f��z��3ч'�ŜLN�2^4%oc�X�C�H�'E�����|pJ�����ʪ3�ҝ�5��ԳW/���r5��C����I4�����ck�X3!U]�y�j1����;FJ8׈�< z�ϩf�zrT�j�P�K4��t���r��0���ׅ�PL���zz/�0��0��fT��Ň�q�2��O��Xg!VG���0	�*��Y܊��)��3�G���>޾�ϵ�g{�|����"���H�T�TQm�PAa���i�\.cc��=v�Ɵ �Z�P���Dh~����+w�C��rȳ���)�P7�lz���=��{�5�����*�NV�VT�R���m�1K�轪��x��ym1�zf9���'e��3�ϰ�Rﵱ%ԏt駜�b�zoL���EFxC4y�=p7�2qK���O]����S?'��#�;*��>�?��zi��۞���󳫥My�^.�|�Q=&7��w���<|~Y,]i��|�Sr%��*�ƽ�w�zc��g�!�	f��s�M�}�s�א���Y��|F+'hqn��i���<�S��1��]^y>g�z�ɖ+>+�M�'��#m���,� �J��L,����n���Ҵ�OC�Ls|>����wt�s��.ʵG�gO}�d��dBy��P:z_��v[�g�����~5��j�v"�hԖ	�ζ/>`���l�,�ݩ\�I?������/�%5m�gŴ�>3o��� @���'_O���G�_����܁�"(pPR��w�
�Yvл�ӗ����jT8�Vx��Z����
�<{��J���NL�冤{0~�)�R�G�A0˩�tV��l5����$�k��'ܪ~[�:���r��ќ�["a�Μ�2v3�"�up<gs4y����^�bB�㙷V�2�{k �Y�W�+�{S%��һ�{���k���9"����L��	:n�G�[�`��˜��W�FYwo^M��"ۈ]�$oWB�zwL�v]vG|&ߴ�`�dN�bfA�[��mf�͹k�,Μ�u�ok�k��@���P(g� B^��T���@�R����}���(��	U&��B��ߟ_ԁC�́C��ֻ���@�����y�~��]�����^�پ�N7�Ƨ��X�A?�A�O^9��8�q=�ӝ�4��L)�+��BkK"m�h�{	��Cȉ��'������QflF^igA��*��Ȟ;��bRi��Ïf�p��b���J�<Ci��p�$���x6ng4XG'&/q{kg�R��Q̥mdX&�U��38������L�hH��[%��]��	��K;y�+������V=�[0\جYvw)�p�i�f����P\�&��%����r��:BWq��$����ʑ`B���Td�"����챢����5�x�2�fD�iʻDY9Z�%���i��M�Vv�4n��A+�˝���Y^$�Az�}��.��p�K:E_1�xN<�ЫD�5M�Ȣsq�ځ9�Fìjtv��IQ�Ƹ�̜{5`�����o$��!P�q�2ddfh������-��dG,i��{\ݦ�ږ���V�'�Ť���x1�z��J������o
*\E���:V 4n���AŪkkw:^��"7�	bd�Q�����FV�ԭ��@�<�U�(uP(m\�Im�����Kl�䵍I��2%���fI4�V�����4��$�̷��lz�8m�y�]�O%�6��PI���n�4*!��=���f���"�6�]z����NWH�u��R��O5�!x�چ������wWj炅i�vl
n+��ز�������#/d�d."��VH�6�tp0��6��s8��E͆���3S*��wM�B�t��{�7.��kFvuʚ4LZO�6LVֶ4Q�{6i��7)���7�d�7Z@�6h�[n#�Ѭ��y���tf�X�*������[{{��F�U���[�����8.@5����p-��mo̐�z��w`�޾J���Yl��g �V���X��ʹ"���S�i�7��^r�틱!6kgnhE��G=k���a��b�+!�{�uJ�kbxGpѽ��F�7�%3��S4Y��[N��V�f�L]ɏ1*X3!b^���+j0�
�I�B�2��"b��j-�n��
��5�<�f�,�VfRz�k�I+Y�8�~�6�����'d�����V����y-p��v	�y.��l}��CS�{{+���l;���)�wRW�/quȏl7u�̅�a,�5�C��L�Ӵ����yFT�'I�%}���k��N�����+QH�Cn��h�7�'$�Nē�V��ʥ`���y��ލ�n����h��d�ْ����y�$�s|Gl;��{��8�&��v�lmyM��3,�&,V-{ai�-������f�7���=�����&׊��n�����Ѩ�h�b+��%}&jݣ�,��,�a�e&�n�XɊ�P�7w�B���a�UT�8.�zy��\p�M�Sѣ�Y��](���5'Id>�c����YW	㵧���5��j35�s�q�͘��i���3mQ�b�n�!�%E�v�wH�EY�I2��,˲	z\ov{��7Zt������j��V^i�&ٸ��F��M,�A+"d�H\7��4�jH��x����O	<{�V���&qh�J�K�.�L�)NYŊ�yL��)֪okE+v����q4���B2����v�������E�^���Ρ3dy3�����,c;��G<H�ڪ0r9�g˛V5��D�ܻ/r���1c5"+p���5�̣�h�ڢ\�/	VEH��p՚�j-�Y� 7kFC:#�*X/FQ[�3�N����4�a��7��OtY���3�<��<C�!+F�;��Wu+��n��dT�&H����"
</�F4��M��ݗ�[�u��U�;F��O)��Y�I�v�F&��Ȣ��;a˶7[~�)�"�%SY� �¡�	��l���TKL���&EU��2�0�����~�
�/O7�y��.��ӯ�@��[��C��C��@����D
��Mj���M��{y�Y�v��z�� P��({;^-{��ov����3��x�x��H<-���.ݿ��e5�G^��m� ?�r 	 r}�$O�r^��ծ%Ϋ9��-m���,C�wsu�b�2�wgZ�cU�nq5�̴��u�j�#lT��m���p@  s)ɕU�i�kJfզ-%������m�V͆�m��jն�Z���[���U�5Z�e�l��`�UmK-f�	j���ڱ��jh�)��    @v��R]��� �C���h���Ѷ �&�۲�Tl�V�U�    � ��@�P���@t��4�����9i�4m��F��;��͍�ffŌ����{v�4k^�{¤��&�����^�
�e`��z��ybh�糣������Yڒ�����:�:�ًZn�e�۶l�I����P�P���Tt�}\PW�5�V�x�t�a�V��  zJ��LҚ�-;�J��;א�ܮZ�s�⎝:�@��G�ӻ�Y�u��V���fL҃�kwg]�k�m���X�M����.��=���6�u�QE��`s[z�ު��;w:�]�{��Z=�uV]ݥ5�����y�۸�F�7�����q�m�һ��6�[`�yyN�-�6�y���ֵӭ�^I��5X�&�Tn�.�,��U�T5�z�=f�V"۳ٺ��������kS�����f�\��u�km:kN�Tj:5V�{���s�#��8��CTq�c��v��=m�f��VacJ�)l��{���u�]݆���oZ���m�\z�xMm�/n<��u��l�zu׺�N���wx���ٯb�ݻZ�빷�.6��.�w^;{M���[�6դ���[�aAc�ճlm�Z���6����wm���6��s�G���{Ǽ�Q�sNJ�TkM��u�u�(�^u�QT;���Yv1��Y�^��wt"ܽ�y���w�Y����Un-WX�E����w>��+�3:�kN��[��R����k�]P�X��Q���scr{j�z�H��6�"���c:����N���.���;�ax���WOy֔�Z�n����5�U�ͪ{k�$�@�ܝ�F�ݳn�7\(��Z��{ox��{�E��<�f�^�I�=Ǽ�oq�[����zSl7n�o^��%֝���^�R�Ӫ�ݠ�l޻�=����SFm�i��T������*:�.���z� �e�󷻣�SvJ]T�����Lu*��%�<��-�'�����Օq�ܐ
��7uQܫf$�^�K��v���y�[3kR�Kl��-�m*��;k��M�\��ES�F;��(�]�-����)^��ǣ�U��n'V�vg6=��8b��룫c��z׼P^ǮC�캜��v�=m|3���SZ�F�f��Z�1�[V�-4�V�+kjm�p j��&*T��  ?h�IJ� 4 ���ҥOR<� � O����� )�Iꪠ   $�@��"�A���z��L��}}�����`�}�1����D1��F5A_Z��6R�y�iT9[�u� �� ���kt����@$� �!	� I ��H��?� �$���$�I1$$�I<�I ������H����"���/��d�����g�@�N�EY֠�I*��Y�
��[����s~;g4#������ˤ����%���y�ȋA���u6��3���A�D6k��[�m�֤If�I�RN�i�ܗE� &35�5��+b)�w�4�3-�-�E��*-Rѵ�2�#mQ3�aQF��].má�c]^\�u7n���@ɧ�b��mGVb�e-��m%��osic*���g��KB-��I�Y�������y�ڧ�3y�0,�B6�N��Od�CRu��رإ����v�N<�z���k@:��̃
�^��SOr���8p"h`rm<gr�z�ߞ�(`z�F}�5��K�u�i�5m�B��=z���i�*c`;r���[%�Bj#O-����1ҵ��^�.�M�V(Uè�
��M����Ӱ^P�����*-��`͖U������f�Z�i=��./i��.cI�Y6ºq��@�H�QT'4ۇ��/��!Q氊,
���`�QX����ER�1��E��"��(1��TE�Œ�ĕEQFc���=r��Ր37�l�q���*�R��T�(�!$Q��E��y�]L4Tt⩬��V-�0�nn�{�4
�Va���r�����!�C���h���J�n�,�*��C�*.�+�7}�Oc{���ǲ��!i���v���ݔ���4�5ۻ�u��gUC��k�0E�5���x��I������R؅0�8ƅb�g.��Շ0�)<�O/R�)��*KXCb ��Y2�+.J �N�������[S@w+\��l#O$��;�l�u���5
t$�(nt�9xl�2#{v-�dJg���R\n����@��eKױ���ab������M��պ���i��;e@<�u���#
�����a���w��ۖ���!b ��
�z�X�zU�vO�SJ����:�[��fLŪ��g� @�<����jȨ&�'�y{Gr�S�34�f4eehv���'�4����$�N-��0jXT�������$�m^T�r����r�6?�{k8��kUiIR����:.�M�7v�\��/6N��k�&0�EX�`�T�0*m+z�Y	Ӷ�'�T��ЬPQV*0R"��(���aRc+"Ŝf�箲��u+:ՆZ���!0U@QT4�d��h�,H��5�ohbB�XQL,e�� ��������7:�����)�ɔ
=
0�"���٠�(p�7�@���em�[ue0[�ܽBN�Goƍ��U�a8�b��1�w�Z  �^���q�vhEb�ϵ���P�Z�5��^��ʙRֹ��H��0d;��?��֒����"��7b�Y� ^�K�鼡�m�$�ܶ����'d]#��1��,cp�cį����Hm�y��P���	b�)�T�X�޸C�U��btw^~��X"0���oa��$5�i���Y����b��f�,T|��S=����)�(������%�x���!v��n�R.�F�-�*�i�"�Y�H��V�� 4�AWx�K�����AE��G%�e;�X:����kV�5n���a�V*������d�*��6��;��Ǆ��'��*I�)��=ș��e�ܙ%lh���bE�������&��i۳)d�sb	*8��V�jC��hmJcV�8��IwE���`P�jTw�E��˧F'�a�Ӑ�	+��u2�]��ݲ�0�-h�[1N(1EqXk{if��Tn�!�6p&�u��B��<�4�d�)�b��j�-]MřZ�����G�aj����˄�8T̖>ˡnkopB �*�y�.ʥX�\�J^P,�>��v29����F�V�B�rV�b5�P!�{(��	����J��U��H��Y��l݅9L��iDI#ܠ���U�cV-��4I{qP��x�[Y^��֥�3k%�7r�N��=����<��a�Rq�Pć5-���W/cUN�����<!���G� c�V/Rc%,�',���
�ׯ�hT1'��H�]��aD6�7
֢�Ƈ6A��s.�un�AD��m5�Ik2��LN*f���Th\Z� �6w6��� �Gf~���=��'��9��H�)1���6�\d9��Xr�Y���o\�:pT0���8�j�Se��$bp��"��T)]@˻	�#�n�l����%�1�w2�42�z�%^�,YOQ�{1R��⩭X���haC��RlZ�Dd�i�Uui,1f�����ط�k9J7�>��W�|��#��9fk���e�)aY���Ԧ��A4����MȊ�LbdYN�n �̒���᎚wI�H![�#N��pf9W0v�B�h��RǙRCT���YI�1ɧb&��OS��j(����ֵ��c��x��0R�LՎ�T�D�hm�9��u��B��Z��̿l��&.�!1���Yn��r�[M��++�>dʪ����k[��⌔55*��V�j�[�r�U���;f��z��DU�`��a�B��QXxέ�R�ﱬxk�ѹ��4Z�S�=�6�b��5{�If��͎�R�DA�Q%��6�B����ڭ��j�m�IFΉ-b��I��R9������Y5���ֻ����u!Ye$��y�X�V�ٔ��z��r^�r��в$��4�*�0�̫�E�bC/l�2ML�`�ɘ���Z��2mZ���(MD8#��R(sP!F�M��t����:[Y&^�P5����T�6E�))2��W3+�x��4+$mْ�+���*[�\���P�h�~��l�4���N��j�W�<pl��u�"T�X6f0�֩A�j�W�F��b:u���$�7dG+H�Q(Z�^P�Ui��<�,*/cUn�=.�Ȍ���!�\�l�J��ʋ)�� :u(�7��Ҹ/A�F܈ S�V�64e̎���2�Ip��톱eǗ#ے6 �(�I{S^~�P�vʨ��V���H�����۵�xZ��>���A��H�ERKC�f��o	�v�+)�[��B��J�
���ܙ�m��XFe�"�%7blSy���[ʵ�si4N��f&���Uv"zȖ����M��®��َԓ`80������$nn�N�C	]�N��X��7pan^�a!h��zp�2ƚ�n�F+ʭç&�C|��6�Y�UjoT��P�i��u$÷���u�/;���w���m�u��M����DDY"�gy��p�fo��XJ���3��	���K���c30�6=�뚽���o�)I8�<�u ��Z�Wm�kz�c�v�"�� �7��E��c�WJ��c������J5���["���M0�YcڬmQTr�;�S������$&Q�" �����d���))�0�h#D�ɴ,
�{�jf����E�D״0�ਊ�c�i�	V�]يd��i�w��T4���a��5mߍa��c��|O��5�p���$�
`����7��a��u�P�e��Cd"HwM@ӰWn�S\�,qQ�B���T��m��F&�5��t�[��X&�Lfv��e�,u�P���pg3.�&<F�6;oR��?ʛ�ԭ8R!\�^`�U�;p��"!�04P��Iy-��Pՠ���ɰ�*�4�ju��^q�&&��Q�sU�%����o1V��T;�H���v#c\���
��v�� �7�˩�� 16�7��"�S9V�	�m���5
���)�6���7Vdxi��-�8i����ڲ(wUu�Y{���n<C��� ��ͥ���a��c R��ل���{J��t��	DFp��ʚ�*Z.��w
�(�\u�H�(a�V
oNe*P���I�P�wx�$n�,��T�����!_Q#5T,�V�׮�c�W'�+��x�m�u%[����x]�4���,�b�CU���8����tn����L�{�f���>�=�>����QY�Rd�2@YWZ�JT��9���UX�#62J˷#�q��ʰsІ7Ѣ�mZ�PX*Q3�n�қlX,�����UM��[���WX�n�>
�^dxY�*�����E6V��:�;�ˏd���������m^J��1\�!����P>���U��H��]M�$����@�-�L3,^���L��Z)`�U1�w���B�A�шAOm�y
�eYS7�mnس�#��w/=z�ݦW���(塴C6$����)e��̑����T�E�J�FC�7Q�P9��C2�S2ٱ@Ǝ�A�L��ۈ�&4���%��Q�@����[[q,E�b��K+8�j�E�Ʒ-6���
7���XYXL96�neaE�r�d�M��1�fRj-��7k{
�c6��Ӵ1�uq�Y6%�����ӊ�勡R/L.�E�<�]<�1����K&���:m´*��R^;/LxR�&�Р)cJ���p�"97i��`�ݻǫ$�"ҴC�d,�z�`{�� ��*ҵ}��X�V��D�X̫̄M!k A�X��X;[T�1�ڞ�*�f��6��B��A<!]f�l�U�l�!j��j��ե+K���j�D!�4��]�1s8eL���h�ilڸqٓ$�6u߱in�2(i���H���� 4#̼2���%]����iR�Y2����Hi���bIҊz4�&��Y �F��Z��^I����G �H+	F�HJ�E���&s��-��q:Hh��I-�K�/C:����Z�+At#SVc��I�n$�&��WM2�EHV)��ePGiR(��ۑPa案UQ�`f4�%E4�1U"�f�$4�B<���bm��� �"��p�-����[:FeK������e;�,j�VA�4�����VP�C��n!"���,'���í�1�{�m뻤���2�Wo(d��+�l*c"*��F؏1֍��ZBZ�ŕ%[-m��H� k�5�Bхܙi��Tu���1]d�R�4�O6�<J>�w��L糝ㇷN��4�Ą�	����Y���t�q�Y1��3�$9�TN5f�@�X�-�a֑-(I��ʁƠ���D6�1t�ą@��X3�Y:�PR!�!�0cl�NұV��Hm�P��:������z���=�Zۮ��2���y5�'m!��,�*,�j�<���b�jE�H̲��
j�m��i�B�rتq*��B�,Q�����(��AQ�V!��*�(-B��JΡPuk�+�:�I�V"q����(��%C��B�D���+n��4�~|��O2Y�I��Ĭ`���R�8��x�APc�T�2�*0>���3(�ŋ�UB����`W�UA`��n�UP`�!��`gR�Z$v�dR)��D7�J��a�m��.�����(�AdX��J������m�n�=���I�����Br�Or���b���n�2>y�!|�Va�6:�B�	r�˭Ha~���
	��i:�xwsݚ��k�L�SN�C9諾�G]wNݵj����4hRܤ�>y0�����:���ŧ�<���3z`vxH7�,#��]�`�쥃*���el�*Y��$�5��4w�f�.� �J�������EH���QR�iem:�����Wn�B^f�7P�#\�s�b�)e/-��f6�q��Z+V�{y)�M��wu�/���NujS�V����*K�GX<e���Я������*��
AP�M��u���,},����g,dp=Q�m�S3K��H��� D�����R������X���Y�)�*Ve$�*�⮺4h�p�j���)��_�.8(��z�S�l�mICR��%ct���]an�Pܛ|:�	�V���c75�շw�ٳ�ذ�	'���;kz�Fhy�$볠�CU��>��}�s۱s�6�nT�'�X�9ٓI��P��`�g];53�֡�Sxl�"�`D.#��=��9�sm�ˮʔ���oGm�����[.����
BF��N��r^hG7[�`SSD۹ù�=���FnbA��6��@D�}�\L�:h#�m���f{�k>�1�	Yռ��k�ҽ�+�m�Ge�j'�T�)�;��Z��X�˗��Z:?#,��v]q���.��֤"�|���'�79eqf�.�� �PGq�=;�5ˬ��ݛ���⬉�-�m�G[x���s��s�:W��g�䩠P��_T�0Ȯ�eZ����Ӡ*F���+�.�ų�\R� ���JB0�\�v�`�YZi��ۦ��Ō�f�o����$���jh}^���]4�%�].�.�ҢЛ�
��ݳٹD&QO:�����P����A=�i�qxb�0�ޙ���4��c�'�����=��kk��|�`�e]��ӁU�Z7�0u�%4�K��ާ����`�3�uڅDh4v��Ɠ����{2:4��6�̕��3w��; �q�s�B�e�@:��֣nh��g��N�\�	W�0n�lܥ��<h1ίZ�;U�%�'u�w���ʱw#�m���5;;m�Y�Ȥ�N%7�����'rf"�+;�^��" U�����U_E��v�Re��D�C�e��u^�����jR״k�OL�L�9�L@���V�A����Țhe�tnZ���9�]Z��`��t���S����c}���9��yT$<�%�x�fe���wB�g��Dz���b��؃g^�R����E��; �*��9S���5]ge)�i�9��ޅ��쳛���h;�����Ψv���<f.yر_92�i{��}оS�^Օ�e�y�1��9*��2ok�>�Эch�}K"��Ǒ����*�>��⢁���g�s!���}`���4x�3�.S��@r���L<��v�Ԩ��'8#X��R��rc������Ayj�[OlW}��_ȶ��\��0'sD/�5|6RB����Ʊ�qWd#9#�kZ�3�]˙+@�oX�Jmt���r���͕9�:�=�ͦŉd��U�٘B���uq}��eL��q�ʂ�(���ݘe�*��>�}xL��q���J8�ԫ�(�.Q�f�Ἳj��u�NL���Z^�C���o5����FLF�N[o&:�RS��[Us�`�B	諁��B���I��ъ�u�gt���j�s���J0�r�ۮ�u��X2��t���z�ÃB�֥�n����ް��Injn� Hճ�-���o�����w�pzj|�g�����AP�m�����f'H��y��.s�<~�n;a�மX�:�t����*�6�e��;D�"�-�uܢ�
���r�b��Nę���.A��،2����{��z�A����s���������.9����@{��+��d3���ߎ�w�e:}�i��eմE�M��D'&us ��k�ak�jy���1��5�Ev.:K�6�	��tă[�e�n�f*��H���Τ�`�ۏ.�h��c�O�K�m+��_Y:�u�	\�r��mQc@[-�P�����ك.�La;.=�0S�]S��I���1ܼ:w����gGR�h�����o��P�&���a��ж��q���mK[Q�`)Vz�8Tr��\�Wo*b���`kb[�N�&ֵX�Z�q6���L���&3ZV���i���L�Υ܋U��\��b=ݒ�5�:�b��pM����	�6Y�V)b��T�����u�IJeI��,ʇ�VEyC�ư]��{Z�iT@���{�՜�?<Z��Õk�������P����t�o�h���(�wN�w�+W{�2��:мu����n����� ���a1�5Lᓋ���- �Z���t0f�F�\T�hZ塽\�5�2e\��	QYDc�2<���Vr�ym��'}��sr�Ց+';�Y,���#�1q�B6�*���'6
�[���d5tqN����!��8�|�V.����B)��h#����!�Ս
��]��x.HRʣ�k⹒��3zC����+3�(��Zc�ClʌfIg�/��d�α\��<\ u�F�b�Ђ���v�E�c�ћ78��ռ믘������L/{�r�i�g
�v!t8{BS{�s�l+ͱ����*l�&����'��M���)�ڪ���8Vډ5]�uo���{���*���U���2sx5gH��ސ�C/t���!�}�䆆I�F���6�/G�y�wU�_U/W����~eT�72�q=��L�:��q�:��B�s+�_
`JO�Y�4����������m�{i	�n�[U���}�(�\�r�ȷ7�n���qfj�8��SwO������s�r�MV+�q��)r��fV�
����dn${$�����u�ut䳠@�7���x��%\�s�I�W�#V�wd�b�IC�W��fB{0>�.�Ѷ�FA%�i;=4S�g]-��u ��,.�M�82��7������1-%\�:s=���Dq�K�!+[��#{s��iM�
�f���D���m��_�U�;�il�NXo7���;����`)�.��.�6�+A���,�Ԋu�B��"���XZ��j�/h��@!�aފ�=�(��ʡ��8�f���]��uU��= ug�Cua;�)R�$�XO�6��}�^Õ�-�a5`P%�g(�\��¤n92��������0�/���:Ʈ+b��W��(#��1�X�ky ��a��;xM��)t�r��U�v:#�pmn�E��{~�\M��찪v�F�m	J�48��e�y�U��nP<ɥk#m;�.���ZX�`�H�G8dd���O�KVyK��I4����E�$����t/���t���ܥ��-3y�[�}V�&�����C�\�x�a܇o:𵹩d�8wt�~r1wCީ7���SGN���5R�w�ZT�x
M����+ٜ�=��5nW��l���C��Z}˂���)e7��M�L%�gj�ǌ�U���8�)��ͣ��hT�
#Y�ݩ�;��_���ǫ��[�u�x�o����܍փ{�M�xGEU��"�#�^ V<��.��"��-C��tHs\2�hUX��0�3Mn�]2��2�xͣccؐx�N����aݡP���NRͰu����,�ddj����Y��'$���w������ʊ�t�����CHlCq���C.v�1��Sr�zI���X��W�-����%�Y�4u����7w��X����؍����Wv4B���)�Ō���.nvm�P��`�P�D��]�b4��K��������]���Y�(r;���[x[��H�Y�f�[���=\����^�m�c�ݢ�Sg&���h��rgj(n�n����\�����.�з��K-�T��ᕄWH�p��"z�r��[4�'����nj������P;B�8�tU��92�W4��b
���e,�:�\+E{��O��V�uԥU���l�����r������]�W@��u�-hF�$y�X�ݞ��IO����Vy�y�t���
m�Ӹ�>��L����W���F��`�L��D��^rQ�\�W�s_mt�D�t���<�3�-g4-��p귎��k��M��$�2�*|�P.�a�/��n&�ooD���<"��)���2�n��_TI��ғ�*�D�ۺ
{-׷��%c:��-��MX���%c��nG�%�d˙�������e�玶n�D}0̂b��\]�i�4�[}b���G�ۡF�3�9�U,3_ &Zǵ�(V$������\���Ǖ	��/���d����[s+�󺩺�6b�H����m����ZΩ�&xB̼��a�8氄�|�%l�/iT�n+����s�c|�]hg%�"����+��R�e�4(ɭ���\9���K '�whp��&��>�j�:,�X�;��,|,�z���zI����#�(�]/I�#{]�/.�Kz���
%=0꾩7���V家�nr8�D�Qk�.��o$�H���k@k�M����C��h�y�ث�=��f�ӵ�
Ѫ�e��5v�l����&��48J��xA��Mwn���a�%
-��s�4�S�=ŢA�:��1h�ջ;�!�juK�Ĵ�q>=�<kp���
���gl�����P+U��:>�~���<9���U�4�`�r�Ҡ�e��Z`�^��272�vwh.&h։{htMoi��!�mÖ��i��n�E��[т�t!CS��'sT�7�T�aY�"N=�\<f�������(���л���-�]WY�<%k�;4ݜM#4q��96�$��6�Dn�cw��	"������hܭ����ڇ2����AN�H�e���#�	�n.�6��t��1ٴ���dB(�ȇ1}%�z
��Z(ۚ�Wt����kcnm�"���{ֵ�hH4'V��-w���{��W]��3�&Lj�ҟǾ��ͱ�Sř��F��}��j[|�N������\�KF��m�bS.�Ф$�薎�3M�*�t��Z��a��6�Z�o�V��ůAVu�g\�˾"�����W�)@�Ԭ�����w��wD ���q��6e4.
���m\�A�έ��aYR�]-���*�+�6�޵��-���)u�\��q餐��W�:���ðFv�����7"�+�A:�cJZ���s ��-F����k2)y:�%ZN�m�gg<�ܔB[Yku�;v�_N�7n*ݹRqȮ�c��V��j�Φ/��oZHX�v�k��Ǖ��;�]OI�p,�).���EH Wj/��4��흩�&E[�@���Ul�D�� ��]S���p�r�S�b��=s���,�
��}c79i8%R��[�=�yc��M�3i�Ձ�"���-[5j�y�4���E4#嬍�JL0��t<�����)��fg+ا��)GnÖh�^:�Vt����;8�nsnnn��0|�h��$�]��C�����NɁZwf����G�A�C���ף(��A� W��3����w*j��q��q�2��7��_1D� �衻\a��*R2es���=�t(��F�<ʷ�/JC��Q�i�\�hhO�QbVG��*,�0dr7��p嵓&�Vni�j=�^[L�;�O%rc]҃�4C��y�����Mv����`�� ��C�fIAQ�����vΡ�ڪ��'�����ʙ��s�`�ޕ\�r�T�E69��D�q�os0��A.���P�)cgm���F�\0�����ۈ��r�\Aڊi^1p�#�.�7�b�N�Gkȫ�O�2�`{H�fp�vA�`�C��E5�_j&]�h�<.��]J��En!Y� K��R��T�1��^R�'V�i�J���A����gk���X���,�;5F�"�Q�+�100��M� C36��V�[�j�����f݁n�.\Iw[�P�K�9�wT�W)�nu�59^��eu�.���;I�a����&�A�e&�E�ܤye�b�ʲ�;/�ʸ��=T%�k���y�����A�]�֭a�̵c\�WIw�ɩ�Cj�������݅ީ�1�,��Y��m,.��ZX��F��b�e�a#�q9�h���l�k�Rt�Y��̸���0,)��mX[gja�5t�qa��=��(�ҙ؍N�Y����(�4�W8���j3JXv����N����_��ۢv" �	�F����дL�}�֕Ğ*����+��Sq������1N��˫;8�-�ܩ���|6�7u��vu��W�����l����G�o)�a꼧98j0�8���Fe�Y����Bg;Л�Q���ӻ���w3�V>۳�]�?�*o0wz��[2�PY�\�
����i��4�k�:�*d�c��yd��V8aK3AT�	c)u�J�ӡS� �e����J]���M�aO�,�]0
��M�2Ae�Yw9��F���^��t�e��>̽3f\%��FJ������#\��q�:�K(�i>���{"�Z��&���G�2�"��Clv��xhu�S�V�9�tY���	-"n��y	R��B]Qc�)3�,v��k/��C%�dG��\�n��9N���1����P�蓙@&2<�/��%�v�f
S����؇���!�î7��Ֆ�^@�c���@98���f%�s�*�n�o%
ë\��6��kja<��5�k�^s�nm~7�[�h���	 O��� P �!'���IHx$�0� VB@�I!0 |�!�B�$HBT!!��	�a&�X@YI��gi$�H���i!��2�`N2�4���	1$��$� i�6��	�����NMr�v� �J���'�$�$2N0�Ր1��B}��H�I�`C���I��o^ԁ7�`[a&�[	��� *<�����I6�����m�ZC��C�h�!IP���i�ul&Z�J�qu �$�/i ���u@����I�HN��d6�s�I�I�$��&�$��X"IX)r�?P����B���� V���XM�E��	S��I��B�>l&�i$�|ü�I9i�R^�!6'�"��6���5$�s��sy	������ u�@��i���Mv�''-��3HI��d#�\'�B8ɳ;���+7��A:�j���Y�BVk)�Cl<��!>�$�!���(�!�L�0�l>߭�R��H}�$�1���i*{�](�T�l.�8��CJ�,��K�8¤>I9�,�ba:�]�]�]���ēH4˪�&3��2w��f�f"�z�=����?v�2�N	8Ì����,�>`q�'P:��a�r�g�Em�Jʟ}a�X�C�]t�Nv�~��5��'^r��i��P�K�~��'P�ԛN�]��a�Sh�cƂ�.�^��#>gCV̡m�6���r�$�ow���8�|�r��e����|�03�=�4�l�z���٤�����m�a˂k�.J�I����}n[]�g}O'T�S�2kT�)>�6�5�g��`e�R����9u��N����x��ə�q7�u�w.��E�,��l3��2��Q#��vc��0A��٧g	4�$����X�q뵯�eÚ�2�@sW/{�}`m�hby���ϻs���1"���WiC8�ƫU���/��\k�'2q�SN']�y��|���y䫅ki�fu���A�c��Y�C	�)Zס�b6�(W��Mi�X&��T�ˮ���F�ȫ�)h�+��X{j�6�ג�Ed�H�XD���o����U�qX�퉶Eu��C���vN�P���
�!�\�d�m7x�yz�V�aj8ӵne9�lHi�5d��Rq����X�t���v6�`�x��;�}2.��60�olS�қ;Y{Ǔ8:����cJe$(6��=����V6���0�f.:,"|rfd˙�)�磇��OS#T��y�=�C�鶛��v���ЇAzQ)7���8i�y��]�c%]�F��`i��gE`�·�m���k�P��'W��U�J�O>f�f2��H2�����OZW.tIr�7�=��䷖R`<#>J)MպC�Xsu�]�댁dsCK���f�!��q��+*_�Zд�`�$�I�o�#y�9VfL�"n�h���6���z�uĔ@u��[�\�''ڍV�d�A���2]�����6���o�郭Y.p��m��
����,QN��:h��4>�ɫ�9���ݟT�if��}ݸ����_�1�G|�"��&���rS;wf�(��1f���[Օ��+t�4�A=G��Q`u��ь����V�G��kxXr❣��wض%��/�Xt9�V�0,%aܗ�M�:�PDVݧ@�R��ˆ�/�ƍ����U`֓z�։|.�.�R�!T�`�U��޷L#��,s(���ʎ��"W�Н	�.]j!F���9��C��k4�����D��ܣ@��=��.,:��J�^����h坠Z�Z Hд�$C.�s�pL�E�`��;;�l�V�̼Q�T9��::�:3n�[xh�����X��i�	*r��Ps�Us*��8�=��O"5usB�r�Z�T�d��*9�l���!O6k�a�؅�;~9/y�W)*�F�lsv�!��ū�`1f=8��X�<�ZiP���z�1>�P�Ի�^%DC}(S��)l�Y{��z�Sr8{��P��r��PP$ZYQU9c����r�E �"�Q/5⫲�a	\�ν��b�v���IY�0��t���p"8	LP�m��2Qf�ݨ��Hږ���L� �˨o�Z�2`{cq��(]&BͅG�-�V�TJ�&Ql���Њ�:+*=ע`���7v(�څ3V�f������*�o$��l��ۼ�(�Z��Q�.�(�%���7FU�#h���Q�l���vj�r�2�2Dm"�`e+���/t���l��{���rc�DCy�.�7�a:�����d��H�k�L:�m��E�if���Z�I�qL���f	��)��p�ԋU���5�u�Rf��S,L�z�7l��N��m#���7SZ������+9{�ŜaR�n=@JI"
Z�d�®ecS�ۇ�lV��!�Nm�o-E��繫5B��~i,D�k/�M�s%��)�#`7�'d[hC��}BD��m�6�ά�	��\�S��Zɴ3�D楺FAN"�e��*����f��*HYY�9k*d��yu^mdm�r�v�׭��P�DR �в���?�\:��-�5P%�!�Ę�L('no��
���"̴5�ɹy
r��T���V)��϶P7�;8�������D�4�un�M
0=�EL��쉅���W��A�@RDh�����^7[F��:V5"��edgP*,t��&�?9hmn�l��"�6ÉJ2��d�ZץՁL��+2�`zاV�P����b�.���І�!j��a�˗J�b$~8��Pm[!aa�ʹ[u�����v%Bƃ��8���� ��m�9n�n�0]E�T����A�-��u�6eS�� �Pغ%1O������ ,�A�ؚ��q��XM�u�kR�5�"&{{mDRۢ�V��hc���hVi��BH{.�!$�Uく�aU�F8�\Y����� .j-	fѬ��*�vЫ�Un6M��� �d�W3NM)�#Ja)7f�ݍ�NIvf��R��O��QݽDb�$2갌D��Ũ:v�����$XD&�⫨�
�r�o$Lb��
�AF��본�
�m�K0Pz1��V6�) ��T�ۺf�A6(5;8)ءb)GQ�ssA�݂�Gp�BV�:W���++HE%�9{(a�F���uo%{PMa[})GV�r5J�d�^bHk�)�����!=r���
�ղ��pj�W�f����| �ￏ��>����#��kН@M�e~���
��vqS{�%��z��Y����%�1ø�"Q�1j�`�!����#�]�]�l�f�d�7#���}����uu��P\H,��q�ʜ��
�IM�A]B��Q�]�E��gM���82��L�ӻyNQi���+�ܫ�����y������e
O�F=�T��fQ�2�K�Z�ܳr�.:Wj͌c���V���cZ^+宬�A�[ذ���\���DI�H�%1�[�>��Pt\f�雐N�
�َ,\�@��֍yr�KY�2���{˷�B�u���f�YC�BrȗRO�S �B�c*��1�]��,��NԆ���6�l�.�*��_Ρ��P�?�X��a�Կ�����ڼ=*S\k)zem��� ��#4 ���mj=��|�G	������ٸz�ń���*���o�l���kM� *�4.io9W�}#v��%��g� P�� ��3��}�eJܻ׼�=�]�o�J�A���ON��M�tÁe�4m�f�uk�R	�,u�:���8h��U�v�*���ʹ��S��Z�`P\������x�m�*Z��x�j�N�Q�P��Y�<=)�L�s\8d�N��I��Q$-�9޻��q ���wΆ���Ka	����7���\V�嚴�t {f���Y��E���Q\��n��ڇ��P��19\'׽��xx𽞱RJ�&e��^��m$F�é���몏/b�����b�U�q��Z�׭	�[̭���Z�p8Vd��P��S�w��^x�s~��ui���!�HC$��2l� �@�B	��l$��C��!�����*� T�� �G�ޡi$�l����u�$�uR�`�� T�w�M$62H��M�&2E� *��ǚn�������w��s�UV
�*���,ADb�(�++A|�b��E��b�V,V+U�,Xň�(<J�������*+"�F"�����1E��1H�DX���!�(�PU��PU*�"�E�� �1�Pb��A>�Tb� � "1���/�J�j�
�TE`��TAAD�V*�"��*+[X�Eb(�l����(�F
,P��ًG_��,UDDV
�����"�H�����#c"(�+Q���Et��C-b(1QES��($X:�pD����`��Uՠ(�*�c*����$E�E� �$U]�k�B��V1c���Eb�DTbE"��1�����������*�+b*�#AX�F"
�EF�TEF"�`���yh�r�G̨����������"͵E�"���F�UETX#8��ETc���Ŋ��0V#���cDQ�"�E��A���,V1QUf�``�TTUE��cF1�`�Chc1cQb(���]Պ�ŧ_g��\O3Da�>�5�?AG�EUAEDDQb
��yJ�TV"�E_�#?P�1DTtʢ"�?}��QAEUQ����QV$TH�+�T�F"""*;O�jTQU�݅UDQ;q*#X��"�U�y�4+�
�
,Pb(����]["
#�,��UE�
�*1r�
���D��EX8XV���Pb����E0PUT��Śh��6��]�𨈌��TAf�A��1AQ��P`�����1�~��QF(*���lU���UQ4`���Ebq��/�(�2��*�*O�
�`ZTT���(חCΰ�׃�/�v�_t�?2�3բ�*��娨��V:_kZH�H�EDq��Y"65���Q-(�"�E���f��#��C4�X���U-DTTDX"Ϲ�:j�|�b�/��b��b���Az�yh��P��Ϛ*EƱS?\��,Eՠ�M����E�U`��_�0�kR���#iA�j��Qsg�4�#�QY�X�b�Qb�_�q
�"1�JLZ^���A� Q�)Z�����֎�J�)s�_��?uF(�((�����V�r�b��h��V�������*(��(��T�EEM2�
��VT�����)m7n����T�i�Hߗ�4������bO�
��a�B�V*����Y˞��6V'�e�O�
���M~�EUT�w��RV*F+u�j$t���ŉ�US-G��骬EbJ�X���j�9��1���/�Q�/wB�k�~�DT@����;B�1"���41c�(�5EX�YU��7K���Q��E=K����QXn�j"1F *:=�j�b[,UD��ut��E�k4�Zc�U��,U�M���: �EAEFҚK֪���h�W�PV,E���kڛui��(�YU�?kZWIUUɝ51A"w�
�酥]mS�Ǟx4��d"�t^ZuuTV1r�T�TGW�*
�9�Ae�s������&?9{��TS��QEq�U`�ڠ�,D>�������]	z�;�}����tִb�b�����л�TR�Y��/mN�?sj"������[)�����v�Q�(�B��B=s�B	,��	�1��q�$�M ���L�(��Q�u��5b �~qAUTΧ�4 �r�4�1JWߵ�Db(�����V+o�(�(e�j�������ڻ�A44��H��DS������é.�~kfZ��P���]�B��k�]���r��8B$�� ����i��ݝ�f#�Y��׾��y���#Ӯ,����K�M��S�(��c�� ��((�j�H���>��h��j�w4�(�T�K�������Ĩ�'9��(���
���U����&�(���~�b9CxUt�bֽh}�h�����)֠��_j���<�ӿn�|�~~��бj�Q/�۳r0͗n�3�S�h�+b��+7d�浦j�A*Qn�ю��̨����ϳX�DF
��;k��Euo�,f+/o�&��ի��U��ʓ��;s9��<�]4u��?��W�GXA��+��=Ձ��t��#ʬ+Ǖ���îdO��]����xn�f�q}{����r�c6�=��.����n��K�%l�f@Y��Z>A\�վ4��MLs+D�h[����-��y�{�~���\j��~�;h���ֹ��PG�b�DEQA[w�A��*�KOa�5Z�"(��EC�*9_����;�QED-��X���3���D.�b�����>��-]�V*ѬK��ѫ+(S��٨��~֭,A85�QV��.)�-X�Q�"3�B�lԷ譛�>��4G���B�V�U�YQE�J�Y�V.:�}��z�(����*b�|�&�PR-�E>��m�Xg�!���Z���^�b�N0�*��9�Xb,QM7��񁂸_�j�C�V
�- ��o����������UTQt�1��w,1��Ga��ɾ�q�n���}�k�>��*�
�N~���È�f�U1bC����f 飖�,X����ޖڅK�Q"�(�ڠS߯vkd(�%UNڪe��f(��Հ�R_4Qf2�0��i�G�5�lQ>�e�v����b�E�Ң
�~�p���(�g�,��v�����ïJ���F��@zٴ������q�RV��"�hn��z��]��E+;�QΝѤUՠ�TPA��2��1�5�4���t�e_�M�Y�I�+U+|��xoB[QO�TE�1��m�UVX�(,.R��,��Lb0^��lO��B�!X9�E��Dcr� ��-W��u���|(/��\Lw}��LGv�(�R���j]��B��3�K�h�Ex�>�֪��Dy��h6�W��;�9����8͉q,�\�rǔ)�X���M'�T�VAr�wE55lXʒ����G�M{��3^��ض6��^�G���	 	��{�zdCm�[�yn�_߷�m�ɇ"�,����ì*#��F�]{
�߮.�Rq3)Z�,C-��SZ�8�
��O��8&R���MYU8oJ�,ެèV����
'������v�@lM{k��f��3����&�Do��j�R�����2��"��~���)��{N�c�C�13nw��4�D�������Ę��i���PD݇��8�*o�L�n�%ut�y<�3X�)Q7vk_�4+䧵L��r��g�ͩwfVo�4��	-?6�CA�놝[+S\��5�fQQ�5fa��c�o�8ͥA-%\��M�簩�R��n���S��+#�~p�.L��&��lK=h�l+�"�`�HG��	V�Q��t�yxz7�w�O��d $����BVj�_��+���D��Y;�����0���l�2�&X��G짘m�ehϹ���k+Y^8�kﵳmDDT;����f¦ͥ�EzY;��і��aD2K�nkw�/>�7x�������-�÷��+��/�T>�E�.Z��CI���2�V���h��s_e�h������̦0Tk=�����Ҩ��]0�޼�At�ݸ��+�yo��wJ!��S�(��ȡ�G}{<�����;}Y���,���~���c�_bZ�4Y��.Xs�\��E]��*�-�,�	�7u*RL�ҍ�2�`���k{)�jXWz�T'�*l�f�%�Z#/���`�y٣p����Pq3/"��{�J����.�h������>S*�����k_f�N���3�F��e�Q\s�^\I�E2��u��f�\Lws>I�IQOݼM��9�h59�M꛴>�/�fwE�CL� y�Ȣ4��/�F�=�UTݵ� ���
����&NȖ�[+�B�����TjTG^;�/Z�i�f*�0kaQ+��T�=�UEb5�[v)E��(fa��%f4E���1r�f"�[��F� ��L�<�o�uu�4���#F}�"1&@��L���`�ۚ�T �hK��d�r�9�}wƷ�pk�<����g�U�aXj�y�sT�k�%O���^��5�Ub[�
�.�C�Ξ
�G�Ѻ�ip�+nIelFcL�0|K��\O�Fk& b����h��[��l6�)��X(�ُ���ӛ��%J����y�T�Nl�x�-R�U/�1�8��ga�_���e��? hρ*�e�l�PC'�i��N'�vky\VV���M�n�n	�dH���ơ6�&!�5������-�V"s��ui?e��dJ)i��>��ܸ����Yu�������e��(�*�o{��h[h��6~&6EE�b��e
��j��k���a����&+m���<Q�Eg��M�_69���纩�~��5u76�S��.3�-�JD�
�a��w�����]~4�>��i%G�����sr�ut0�M��,�kZ���wE�n��Qʲ�ʯ/z�r?-�;�{+oQ�(�g�0�;>��V~g;t�w�ރs-|˖e�ۙ���[�O�����U�of�:�Q���j��m�p�z�C���wV��,kD��Ǣ2%GAB�Zs�8�r�{p��wG�`2A����X�k��拫V�{�lݫ~��c˚�DfaP��4:��Ko���Ҿ�0�쵹O�v�T�
���(������v��*bk]m�ϸ�@]��.�JЩ�*�\ʊw��������>�kH_^�4��^%�-U�8wV
��5�]X@���ou�s�8%]g���7�=�n1YO�.��ev�2��0�H�b��_��ԥ�+�^D���P2;A�
q�m�v���(n��^�;;&wG��'l��e��9��PO����u�ht�ڄ��;[NlY;op���L�o�d�-�x�v6��N��廢�S�R��7�HF��Q �Fwe���u_��m6�����Z�%ݬ���1����,�znT�&��V�{�?�QT"_6�4�W�LU���V0 �vhͷB6��e��������-Y�ֵ}�����q)��Im5-j>�ɇ�kH��j�w.��9w���٦s�é�r�����Z�R�BC~ 鬐|�s���=�Y�C��ƊH�y@�Ȍ�0 b	�B_"���1{0(�#[p�0�!^ʀ��P���4I9���� ��I�1E,0��B
�k͝�A,���	�9��m,��0�ͩ���SG��y��I���g64,�����:h�
ؙ?:@�9L�  +�)����JX�����6�*�R�*�����P��Α�W�p(N,�2Hn�}��d�C^��	ۯɮ�R����W-t�l�>�ͦ�N҈����Wk�Q{��ŕl���(��i�!����g��r�Q�Y�m̓{�Vy/�:�Ң��(���k��b��
�֗�MR�UI��d��n�%�X����)�̊
���C.*~�\9��4�g��<n;ؿ^��A���ow�:�&�� ���i"����_!X_��`��1@U�u�ġ�kaA
��>���G��y�QO��T>�S�
�xԔ�H�B��Z�7M-�S�f����4֡)y�j.�TU�sY��q7k�z��k+��Wv�.'�ti�֫�M7�\�g��7��,��tb�og����hZC�8$E�u㜽���|눑>���=[���C�V� 	�I���UY�.~��2hҵNZ��9�~fы8�j�l�<i�X:��
 ׊�V�"k�W*�J�D��jE�#k���V�٫���!ޯ ,j��U��t)����孢)&��U �@�O�ŵQp"1�C_ �`�F/�2�!�4��2��lD�/澺�{�w4��&�>�|��A�qq�&SgN1���ee�Y�������e�i�M�T#I[-�!���=�^`���+y��}[���S��<� <��}˯�����H��f>���
����yٝ7�d�\n��1��Lh���nNF��J ��3��T/���Y��[J���]&m(aY)d h�
�>U.W�_��$HD�b�9��F��Hu�(*�ƥ���hg�K���/R�����Ǵ��v�� ��)�U�h�D��AbU���6�_���N%Jƺ�����l�K.6-$�RJu�S��^����:z!�ӣp�v+�X*�'� �XXy�E5�w1UD?�M��8u�p<�����4@S}r�%�� F�t�<i�;e7uy^�����WL�'�	u��
()�ӯ*1�Z(�[wk������P�C�����E�T�kSA+L*�jB���Hѥb�nw%tn��+گ���J��0^m��E[_h���ʕ>_!��9�F����?KB�2����(�q))�R�C�)qAr���4��k�ŝ>J�����y�N�o�~5)��?/(��H����t~1�l}@q���Sv�-Z��Ҙ�ۃ0W�"۠U+��2B�-�\3
�%�y�Me�.[��G~Zf��Rzr�L�W�͵���Y�D�t���`,9G� ަ}GR.�T*����
%xT�_���I �Դ���k�=шyU�=7���w
����  F�< ��B��*��f�q�U�n�ݯ�A����(�Ɓ!���@�mk1%:+2f���{�K(U ο?u�]�x]΂�wE4 �:!m��~k�d H�l9�Co�?:"��#XdZ�ɝݚ�(�+Y���h�/��a��6*�:B�X{r��~W��>{�-��:{t����0ȥL�8����e�
�a�t[���z�63Ϊ��Q��w�,V>�	塼��֗���|(@l�oo�!�V�ܖ���J|���\�x]�����Msy�R������E-�$N0$�@ i$ۦ` �$��Hi�s�\I�HhBI]$��a�ٴ �۴�	�B�y	�Bo)d	<�I>{l�&$$����L�|S��?��I'�$��M��$ |�2�!$��$ m1�I�6�j�����I� ���'�B�$'�!$@����HH��{�������}���벝*���}���\�~PED;���3ssm�uD�����a��ԭӄ��;��av�s��|:��n�W��х�D﮶t]an�*��~֮T��u�����3�Ll�=��h���v�7P�ʔ >���_�Ty%a�(��������	����C�z��Ji�����#���Cm'Y��a�F�VB]�#{Sf��^�Z�)?�U���{��ڭ�^��z7w��"�#��=�Q=x&-��7��;���b�������xUl|��m�m�����_a�<��Oʐ���u��~����qч�nK-�.�߮��{s�ާi����݅��)�}��3��乞�@����S��9�T���>`Ѣ
�ҝb&���F=֕�^�Z=c��+��-�6�םm�@fjs/�uJ�,������U��Z��+.i�r�ƀbh�q(��?6G�C7Y~�݋Q,a�w��,�{�}���h(�mQ�0U�8�|0RO���!�z�T��,�N��ԯ��Eo����] ������'r���X��e��<1�qSm�\�'����2"�$�+H����x�ȝc�&X�O�DE�:��@ISj����B�I!=Hf[/$z�*d@�w�UP�[����* �,�u7�m�VUU�U�2h����b�eb��Id/l��2б5 �A	1�A {�k�]{��+�l���2�^�n�f≩���s
��ٱ>��?��d�Z�K!�{O$!T�l�@Q�k���𥏏Y!v�<�74B_�q��^���n�e��>`�A��_'��Azm<0EO��hC���� �"���+A�{xʔ<�Ë������.Uxo9ӹ��I9{��k�����@%a��֬4��~���!�����?5�'��'��C�8��q���s��r�;���{Bo�|��ܲM�m>@��o�ں����7I!�l$�?k^w���Y����M{���(��{l���)9\4b���{��.s{:��\�b
��)���}���hf���lS7��ݸ�Srn	r�+Ƅ6r�߶��]�F-�rAu{)x���_��j�"H������@�HU
��{�B���55�]�(�+<��RB�� �X��4����d�J(BCu�nK�u/LNMB*���Y��$�B�b��Ɲ���A��tH����{"L$
�����;�OV<TP�c�ʦ:��ks�è̂i�i���g2��z+�Y��h*!#K���
�e5�}�x9aa/Ɛ�������DRE�����hr$r�ʵſ�7*.��J$l�6�eH���@�O�0t��9�[ݞt�Gơ�lT���b骳��?&�7��̓�^!�]?���QN�hI
��L5�?�F恎�ܦ�W��ƫ�I'�z=��l!��D/_��ǽ��}�V)�I`H��yx2�#�[��y�)ʶ�R�o�Qh_��U{|��m�}J]C�R�����Hf�:|j[>v ���E��#�i����3�U>�
j��`�d"q�7	���<I~J�z��x�X�������rCݜ0h��R=��jΰ ���ؿ���)Y�6�4X�M`f�Юi���w-�hU�V��gY���]��R$�9�Mb����ƥn�`�����:�	M}.c��i~J���6:��� ���b� A��vbc���]��' u�^̢�u�7��*B�
��v�[�@�k
����QRo��y��]�L@��&��\��\��Q�}�"�t��o��q�?�x|=�jW��Jޖ1���!�'�%we�%d����jdqT����p=�1�ѵհ�
D��s)��'Ɍ6nZ�;��ɟ�� �3E�@���+�	�5��Y�Kx}�λǘ����H!1x����ѡ�##\M��Z�eL��ވ�#D���m�J�?Z�w��5��m�h��MO���l����1�J<��(��5�׺����H |M�^���t����q	@1Nj8%u�ewTv��ԊG�׷�yW_�ב����W��Q�^%н�ez�`|�T�9M|��J���|��Wi@��(hj��Wf���n��l���[�Q/�a�6�H�����D����-#饉Xt~�\�{R�Q�ǝ�~��/��:�f�ȵ��mL�K���sG�HTzkU���#(=�\��D�AC�(-���r_�!x���\�z�=Yvĵ��wP�?Ps:�Œ�A�-��.Z�%}'�s�WGŌ�ȇ��D���NJ��	���m+�91��qG�W_u�]�ש�ʺ.�[VG��Xl�c��,eT|E/�Ҩh�Z:k����yx}��>��#w��	-?N������|g d�R��V
���ۄ����~ -ƽ4�ԕ\�j^e���ҽ�^�}�6@�*�8~3�dN�d�u�ą��`{	^��%d&w�"7q70~rS���*vz���#�����G���>�=�O�맯V�H-�r��Ή+���;	��:��q��P�p�/����ë�7�^'�9b��N�ʽ�����#��*�e�t�Gc���V��u��n'}8��4�	�����Q�V�əY|�"R멄+qUey*XoP�B� �	+[7������[�u(�+��
 
�{׼���,U�+��T}��㱵�7�БB_6�}�Ka��a>�4Wq��ʬ�U��=~ϐ�_3�V<��X]��aߜ壓B�!��I!�9M�6c�uax
�k`�6�?x��#+[xrs���>��ݠ������Z>ޙ#�Rt�@l�5�HW����'�E-p�w�	;hP��~�� �j�^Uf�
� �O.���x��ֱ�}�0��bop{m16
�g����3��R)Y���{�n�f����i��[�8�~��,?R��@m&
��Q���裈ψ���4vwc���I��)�l1��/ٴ<��X�o�0�/������q�p�p�����M���N� ����@���,{خr��_��q���U�iZBp�����&8v1�)��#8AZS�4w���Q��߇���N��ANZ�΃&�R��+x�yC}G�a#I��ؙ�TB�WXD�l�����gRM1���U��W^�;`�Ĩ�a�ԩ����I�o��<�:g9ӥ�"�j<@�?Hy������p������V�d�ʖ����V]6�b��hL5��m�\��yՔ�2v�jU�T�gY�^ve�s�")�f8���{
R���X�ؒ���<7{���Ӛ��ˍ���:���ι�qq!'pݮ9�Bn;5ڋf���0q:B��@��5�.��ۺ�ޘ�;n.���À����\����E0�ن�
��{F�գ��+�=g� �}�pm�j�kr��DF�O�48եh��]� �l�ǩ�}м> �\AF�y��q���xCly�=��t1Eiߡ��*���C�A��xl>���|)@���t�mE�.Պ�C�]83�]�S'�;a���Go���X�p[$Q��jܩ`��vT�*��ge�;�Y[���sK��O>ǵ!��W�p����L�	,��X��V�|��Ym���/q�K�i:�0i~�"�_^�`i����J�sh���cB7]�"��� 7�Df]%s��0���#4�P���ÔU!�kjK���<�V)�9��ᾰ�����Vfh�+ؓ���UT�[�{�A���9�z�xt��04{U>F|���~�Ri�U��4�_����!��=y�2��7Mo7�QW�M�65qW���V0~~H�p� xj�z�V��-$��ϽV 9G��[�A[������pMdUMi2o�����=�$T�U�9����[�}AO�L��	$Yh�2�}�E��$�M���`���5t���IF�o&g͝��o�s`l�f�d���l����Q�J����Ě ��\��yȩr�a��:����6 ���J8��uϺ]��_Pޖ�'O0�[���yȁ)$q �9*L�tF;`C����u%���r*Y��s��G�udU��p�=�����d�qcJj�5L?�{�i.�#R�.�$����%��˝f�oa%@#}q�u�puh�z�`�����r�$��s�Y
l���yNJ����\�dH�d��Z��O!�/�=an[�~
��N���U�Ȩ��㦩�u8���p��̻�"z�nOF%,)���e�љCTN~�k�D����u<�?k�,�؍4VS*�d���^��m��I��l��˩YG5���G_0z.��OM��6�jV�MP�UM���Z���YČc�`�N�Wef�v�"��fX\P�jZ�mf��q��Ӹ�jա��b�		P{�]�&��WMS�2�K��j�ݵu��r�T�x�A���"ru��s{zKmRoaT��c�/"R���
@���}|���:�v���Ρ�;L��Qd��鴫�{swȡ��YRQ]@��'^N��������.��\��b��������Bk+$o���t��V('|'�店N����c{%�V(�DssB�s��Yk�g�3S�t���5�2�sjE;�����q�/9�eqE_s��C	�{2� M��9^��������OZ���;��>���ط��W`I�.�E���=�Q�e�B�$zIݚ�K���LEX��(c�0�L�gw,@*�IX�`�֭Qv���b)��X5��p%Sn�on�9��S}f]�̤�D��r9i�m+؅�us9[��)K�8�Lay��5��Φ��y��a���vu�J�}��!n���+�Hb8����m�M�o�F�x���^d�(�*�[YN��`����+��zY�%�v.Y1���q�;����[�w�A�8���F;��6�k}}F��~b,��C����b &p���q�ת��\_7YB���h�}YcxJGkG�y���Y�!�t��]��3�f<pz�j4���vTn�Ћ��M7@S�ۛ��Ճ��R����u��T��U��~��_��s�I7�"�3I�����V�8t�:B-;�z��S#�s�x�-����3y�+�J����/��d�����[��"�^޿Eڂ��w�9��"��G�l���$����|���~C�E=��h��=�����m?��M3Q'죽\�&5�?�)�"v��d��>J�a�o�����DO�i�f��Rɋ���/����DDDY�I�>ʘ��cP���g]�`�O���yC��d����A��"m�w2CI�TX"k�?�+7���Qf�4�7��{C��*V|�1%�=��a ;<.��tH�������Ǿ"�7t:����w�:�2w��;K�^Т�}��+7�T�5�嗔*#���g�0N�Oj�-�O&g���Ĩ�q��4Ȧ:C����`�G�8���pD�y&�6;;�3����w��X��!D�	��H(,�Mf	dDFa�g�Xm
���z�6�J7v(~B�c����07������d֨,MҌ��X,��d�����~��+XǬ��Vh���*�d��,�?�����OW9�I��ؽv��d�#��d�H�F�r�)���|�_��C�?�1=�d��d�7�T��e��+�$׾��?3�"Mn�iQ�ʂ�Ƞ�S�����'f	3�Lf1��H��-/��'q 0A#�@G�~��<w��uP��+%���������31�#�Ʀ��S�q�%Gvk���T�
(i�=��q���d�?�~N��t@ؗ�t��*�iV�T<�`�C�� |G%���W!���`d��ɍ��^���Q��J��8'�1�)_���`�,}u��.�Bzd� l[��N�4�E�F�!MLB3��J�O�;��̽9<���	���e�Sڶ2��eWU��Z>s��&~1�WQ]_d{�+4d�R2 ̩���i�m��ǁ���`���]]\�G����l_O�ږ#!E_��=sb7��M@8��@�U�>�&T��Q�"����or6����s|���jd^����!}+�Rqjpy�������v/L�y��aR�*���#בG�$=j�I�ԙ�^�z~�W婳u5���.zR����҇��V�lP�kĴ+��n�8So�| �����Tx6MS��j�֔8f�!o)��B��h���y����G*iYjtˮ\B�⥺��m��/��m��8q�-R��K�И������_�s G�����aG�ds�4~�7���ђ�����>�F_�F�x?X�'�T��fR��G���AKds��R]���k��]j?f':�NEz�66ɈgZ��ڳ��k�GZ%)��*}��\[U@�I츹^�3X��e�4�I�ls��|E�@/��������3W�HJ�z�*A���ޕ��Ny���ϵ����!i���ML�Z�1]����^v� �3�j�搃-k��]YAP�7?�.�yT}�-�	�l��f�+�&�G/o�8%���G���DAS.g\�v\�O����Ơ`�^��7���_Փ�7=��č�H[7���/S��A�(Fd�6�y~x5����TĔ�^�p�?��d�G���v�V!TL�T����L=ڞ��Zq'k�.G�h_�,���_#�����43�}�j�-S��2�Y�\l�g��<���͙+���P?Z�NoC[�芌�^��N�(��"aJ��ԫ
Q�>Atͻb�|�U%�6M��.���{n�7�Z��DV�	���B8���mN���lD�ck��y��!�>�m�����Ơ�Bھo�Q��|F&A���c���������IR�{��wj%M��9��7�����)����%�n���ca���u*�A �ԽU�������}1=�u���|�&�b��
*fQT!n�tp�4t�RӽK�u>�h(����wU�FN|�jJ��px��U1��19���;s��t���h���]��Tg�Ґ=&�λ��N�D��˺�"�tr�GZ35�YӝȞ$��@d�,��=����+�����[�Q!!���E������Y�#1	?B\v���#�}8=�oi�� ����Vǀ�ӹg�K����2|{�L8�9�&J���|�{D���v�ZB��� �f#���dD��]�%���V��R��kܗ<����E|j8��Jo
x�yG�@�c!�p.ciA��Q�뀣<��h�1I�2���Arķ�Ė�U ��bD�/�X%�w�_E��4��u��8X�=(x�dd��+��k�����z".9MTT�1�$!���祦�oB���
u�[�@� �zn�{�'�pg�8�H�w*��?B_{�"$��C/)�Y[O9Ҷ(b�s3�x@���X32-ǐ�����|�9:� Xފ�0��7S�+��!/N�jjv>���4�Ӭ������3ogC��=��-�e9v�g.���(<��N{�z�sF����N;}J5|��,�L�S�ZJ���X3eJ���D.Dn�
�x0����길vc��3�y�@�xu66u�����C��۱ʲȨ�0}�3c���\��,؅*�����,�����u��:�S���~`��:e1��?i3@�l�C��2�r&�$0��"~{��߉�o#L�,�3��?s`ڹ*gaL푹�Gng��+O����p#�*�#�Io������NX��Nҩc�g�zFi~g8B)��W&��F�V�,��;��W9�g(ׅ/k��ٝ�U��58̎]��	��
�)'.B{!���9jƥ\t�[��l�o�-WYu|VA7Y}�G����D�f�<���s,�k T@��]!�6�*�2܂��x#ծ��A�Z_	�ycid뻥y�I&:M�9��U�;��U�X��K��B~e��|Qfi:~���Ș����s�7]�8P���C�>�z�Wz�Rk��.�sO� ��쇄kc�L��}DJ�pZ����E4�1��_U�*#�:�8~�'�&M��jC΋sI�����e���[�"�:�M�v?R������j���o�#"�0	`��FϠ\����d�6"��ed<� ߦ&�=��z��~F��]6|B?e���	�_ؒ=+DO��v��1�%B�
U�W�fH�^��䖄/+^H�r	���>����Lc
�<$I!n�Ƨ{�6S0Yf�Jf�0��9#�6���HSމ5�Y�ܳ�*���>��8��127B���9�S`�J�c��DN���k ����#�ĕâ4߭O�sU띭�
���&�V#���Zg�yI��}5!y����<�#�Dp�<��"����>!(���
�z�O�p��#Dm��~���xsO8.v�W�_�D�V�J󯪣sfI2p6�tzDW��c��j}hI ���@���]nS7���.h�X[<��gγ�#��bM�<�Yv��:�uX���j���6O#���_`�L}3B�2�
�p)�S>T$H"H�vg�y��(�G6N�>�^�o�$�$7q9�N~��	7
��ލ�TA.��Pq�6-��pl^�:n��2P2Ǡ�o�o!��Gp���{�����ST��"��|�����`�����Q!�[z&@\��W0�wt�&�\q�%��v�yVl<�42���Y���s[��wE����F���5
g���:2�vW���� ��u�;8�.��t�{�I�їO��Wg&mC�#�g`k��9�K��v��ҽ�#�C�FyI�m���5�Y9՚(Q�{��K]��R\��3]l��\١ ���&�R����(���|��������`����ͩ4��۵?zS�I�3��},½�`d�m� #;y\�d�:	�ap��$���hŴ��Lx1��]@�w��HtbJX�,��|�bN��ad�C`sU�e����)�=ޓc��7���������^\����x��O���F[V/�WM��."fr3#���Et�r��>�����h���"�З��WL����(���[=3��@}�T@Dh9�f���l�Tp��I��y�"�[���F+�]'��l}�a�M�LПMr�"��:����`#��F�!�c�?r]�~���Pc���ɜ���̼�'�&�w1U���QM�i@�d��tt�[��܁���<�V�Ni����W>�����f����1�T�1E,�s"�Y�g0K��""Q��S���0�%��-���-,��xӜkC-��'X��p�"���Ѭ���1������y�*�'��N£S����v�^�Ll�[�ڍ���^ѤcŻ�-�K���(u	#҄�*��)ƂD�E��F��;6�4� ���Pca���b�+}|/˘֐��Dx��s;�S���ڄA[M��Fv�nSX��b7(i!e�5^X�$y����o>�A�Ul$���G�blR�V4�Go/���KD��,� �!Z�._ma���؆X�����4zv��6��(FD�sS�s�ө�`.T?I���g�\�d����E�I)�d�6�̋�����^�>̟x]�e���PJ�̸cqM�Y�r*��j~�A:�/fh�:ջ�/�-��(@�iR����y�:iӾ��l��Ϲ\�։�J��g�'u�S�0Ȟ�~
�p�M?~'�zj�ɳeyA~��f`z�F��u@!o��Ċ��H�ݛHh���N�
$��c% |�Y�3o�r{��7-tۮʳ0���K�������X�̡'N���HVR�����м	<��:I�L�5{���en������]�>�� VZ����`�ʿ_��q��g\����*c�Y\�D�c���(��K%�X`+��
��o���Fس�}���������Ր��$DX���6�:�78A�~E�w7��9#V��S�f�z�z�5������X?�����A��$_�v+�?�Ny��l=��b���0#��D��G��8��C2���ϧ���6s�i>.���������ѕ#;7 \f��?��u�|c�5�[�\'��S� �F�*��N��/R ��p7Lmك(��0d2E:���6�m]Y��c���,��џJ�C(�^c'�;;*�Q�ҋ�}�54�1/v��� #� �-����lR	=�=Tk�� ���zY�n�3r��Y�:�a땱5,Z�z0�
W���U
-Wh�Oh���ع�I�_�J˸ч����.��K��}������x�:�G1�ڵ��FU���rثM�(3�~��[�������n�H���P^�zSR>F�K[ǲ&��jU�.BS��w��oS�LN��;��[xs8�λ��������AS?��y��L�����Q�7D�Gf�����Q6����7K� ��UD���8�[���*�X1�Qf����WL�!Ep��6��+Z�@)�4���t"VnM�Nl9���^[�]�a�{���;��U^Lˁ�0媔�Ş�֚�i�9�X���HG�"�J�z&��:��}�w�C�6����4��N���D�zh�=_k�"�@e+��1v�qFj���$��3L���̒���y�dX+��7��Y�E��]K��o�FPAy���Ѻ�P^�z\@Йb�|*b�0��h�<�Pbb�*��N��.9��~_�*$:�au��h!5f,��ٜY�<!�����/7�2zb�y�}��=��:������O<~�̷j...����XC6Xڬ��ga���n��j���8�{�}�=��L�gtGz���q��!��"�6aC#	��g����Y�u+�\�Z���:m��X���<�����%�WOF�jH�䓯�>�)p�rc8���u��(.nw�q��}���|G��ndʹ�~X(��e_g`Qw�٥c��ΰ����|�J���v��d�&~��*�1�l��!�(��w\����dI��NG��2���[�\��u�ْ߳}f�1��l>Z��s��k�.�VV��0���԰aٺ���;b0������`�^�mg>�𭎟%!��S�U�<2�̓m#�E�2�M-%�]w,��&!�
wS{�Bq����Xokw�vf�U};geg�\qw��{��8��>�=�#h�Y]ٗ=���@��T������70k���S�;�� +�y��b=Tg��>qE�.�LK�sZ
����T���ߺ]+7QgA��O<����7�
$�Lt�O��_Y�s�^}aߦ�Q��;����߆�I*5V��y���r^�6M{t�˭��2.xH>�f���Ԛ�gl�ٶ���������E	Hmk�T��.#���lrވp���ɵ�EO9�ˌ<4fY�9E�UMfU�����y�;�s궭Kw��f�7S���uDg�7&das���ԡH�|��\*�fE0򏲐�O0E,�#[�w�Ъ�3Ut˙�Ԛ�c�[K�q��-����@������Z�|&/׻G����]ڪ�B 1��u���{���ѕ��n�q��V��B%�Lg��7��3=�UN�.�ǻĀ�e5��t���yH�y����w�ŗ��Gb�'���!�� �{�h���hF�;�!����m`�o�K�)tG 
&&��Dz�F�Ąڬ5�OL�����Yg�T`���3P+S��\��K���;��,�}�O�\}�3g��˵�&$P�ō�'8��$!��?U�=��lw��Pu�|Ȫ˨�D[ѷ��ɳ���޺{���Fk��4ו�Þ/W�k}����w^.Y��
�L��`�+C�\�SE-�ͦG-gWt4�U�������;Ύ�&k�V���'"F�;<�)�nL��Or�̻˱K�����+�ܔkb�@�P�^TF����SGd�)�^B&f��������,��i���VSQ�Ǜ3�l� �L��%�1�b��r�c�UIT=�vgn9{kgpv�{Kd�{P��q��
rO�9�ny��6	o��m�n��Y�3��^��o-����<n��<�6�ƹ�K۪6��,�^���3u�h-��l:ʺ|L�!2�r�% ��[o��[��v�;�9�|��;|~�e:�Ꙝ�:L\[�k��̯i>��xz�|:��1��p��P3͇��\�*�GdcЗ#;#��ef�E"�,.̪[o��F�U�>.��w�Y�0��s{U������C_�9~��߾��U�3~��k�vvW��E��hl�N����Nsf�g�������{��#B}I[pWau�\��/=�q;�U)ə��%e���}�̟�P �J�!��i:�|�׸_�28�:���V�9��l&:�8����
�v���ۑ��ju����%V[�ˮ��%�$�@�Mæ�]�"c�V*LQ��Ȫ��{iu*�K�}��e�ޡ�.��}u�7m����w�yf�7xݳ� ���^곗��q�}�;iK}�j*���Xp��1�nqA̎u�����Ok̛��/��U�n�?�~a4�n���[k�CcKj_��3�S���a]��!��r}�7��6E�1���Η	�.F����n*\Y]`���x�5�BFk@�P3]B,ۊ�b!�I���uFý��T����K��WL��gBb��<�=z�l+�a���	{��4L�Ѩ��*sd���3H+h�e�h���d(rǵ��]�p��d�W�^Q�dlD��ZB
6m�a���[u��w�(T��ˮ#3��-�c���`���:�	m���G?g�V»���
�xL#��z<��vC/.�;�l�7)_DߡhW�CB��`K������e&�G�	�3���xl)���0SW"�R��c��+�Kzz˺5�׭J�vB?���FF��(�� c����4M>}*V�S׸��b����-�#�qTS��L��툉^��~ꏏ�M�-�W��`"z��P���L\�=��=�\����q|���/B�ݮ���:�^�H>W�;H�zc�~���1{<*�E��D'��N�G����5�v���<���]N���F���*_WP��:�c��j��^&��;ޙܸ����^��=�������g������LňrKfo�w^9ApU�^��<5��G�TȔ�}�v0Z#����<�+��~Ϩ��\G�%�'Ұ
5p�@�7�~���N����g��JFv��~���8%A���6��p&�A鎞ڗ޻�����6ƿl8+Y{p&=d�7E>��yBɚ���W�n�G����.�;&��3s�6��J��&κ4�e��}7�ĝ�Wi��Y����T�9����d�;�o*PWg\�V��wpܛ���o%p�نI|YTL�j�'��d�r��k���D�Re`�w%����IY�!�ѻ�����[�Z�촎��`y���eSj�oC �U����YƘ�29���c�"��*rp})У�4�!�*�<����T;�u�����olf!Xy.�-.i��j���lX�ڹpJ��Vl�,Kn]��̴o:��^�ȣ����\OU���e��n�5�+`��K{����[A�N�4���P�����Wdɶ|V�r�w��5�h��0ѐb5���/I��Ul��6�}.��S��KY׭N��>1ʥh��q�x�q�URo�í�w�] b|��Y�>˼�w���bpǬsv���u���3]"�
�|w�0�̘9��,K[���Үf批O.�s�7dPܫ���s�+<�C����=x�_ìP��[�x���!8�����;ܛ��l�X)��U۽�`Ӌ5ݾBvP<�%��9�IK��܂6���EM2���ո�4���h�;���nK'ǎ��xlo3���V���$�Μ�Ր����YF�K�����S���ns�rŚov�#iSV�7c
����^mmj��c�� m����	��ʬ�`4 �df,�lގ�4y�p�B�1PWK��t-##�a�qM}���gcu��G�#%��Ŷo�w��[6�ӈB�ґV��.�+�Z��ڕ��g�E1PY�^�KB.����C�V�b��G8�Vv��c�cg���ٙ�����.���h;5�X�A��K{I�a����W��a�a�ovpO�j�\؂�Uuֺ�uXU�L��h9-��3�'܏�z��t'+)G�;T��3B۔�т���U��*Ÿ-��ɣ�6(fP\�޷a�2gz���Ĵd�Zre�z�%B��j�=s��E
uLP3c{s5d8�sSVsV�p����k
�Ҕ�ܥn5f�B��8	�ը��Er��ڋ5�I4:�g<
l��e⎖���!�!�׺7�W"z�Y�M)���i^f�N���B���O�a �������ekI��V����Z�t˷P@v~�)�Փ3.�V��ّe>F��(r憶6��'	)m��Et��pK{7f�7N�k�p;/���Vꢌ�{m�z"5b%!r-�,���\%3�q�d���v�d\B%
Y]��up�u�w3��c'=$MZ�kd��Y�p����I:WzX��ƶ�c�IU����ѱ�;��h���a�Z�!4wkA�06��������T�e�� Q�i�[�W:v�l�Ǻ�U�Ր�|���)���H�J�s%��-�vb���]ho��/�$��j"�byㅼ a���-��]�*d˹�����y0S�ؔ19�2"�eN\S�(yTK��  �y��;3h]*ԦN�����D��H.W_e>xŠm`6;�u\�8.���Zj��5u��|Oc�R:*�:�p�`��⺏zǌ��5+<��Q:��j�=�<�sbJ	�Ti�����^ޛ��Cy�5ޓ&;|��ӛY�/�ڐJ���'9��D�g�DvX"g�O��,I�RB� T��:�wqy��U�SѦ�g2�O�]$+4�V�&��vPi[\e�n������<6n���Z�~�}�)�4g��0�7>���r�B\68���~-��@�6����|�rVJ�>=��S�|ö�����?kE�1�>�O�knzl���yB�N��.*�uC(s���*;�ѧ��3�n���M>��w�l��/s�gr=�}R+,K�9��
�veQ�%�n�<��U�'�s�+��r����~K�LYzi����9u�=�\A���KCf�u�cL��
���i��\��<n���/֙G�N;S�֒��.�77B�����$>�ƃ�v#��jw�r��X��٭AO�b9T��F8t�y�i��¨��zÙ��fG�r �1��Gj!F�<�1j��2/����:k����P� ��� 6���w�$=eU�sܔWܻ@d���zx�@��_gj��z~�;W���\-�����t�۾	ӧW�*�9�u.�tf�T��˫��m���ǻ���m�qǵ�B�rx#��om��'��@�9���磻s��x�mG�/�����+B��"�
��*;}EiJN�e���t����4oN�R�ػ&���Rp��?�Y���{2l�7���y=���!�=S�	���AP������u���Y����Q��f*"<�刽^qb~��3񋘃d+�9s�5����.�0�l��+�9wN�%��L;˭�J�lt�xM4�Lt�+�:(��A|�����g'ȕ�3�ʅ��{��VK-j�Cb|ũ�9~�=��i��Dj��,B��"R~w�f�[n �l�#�W?]e6}۝ff6]������.�p��:t�4�Ѯ�O�C�����E�n��H���Ж�W�gG���]�[�{6�q���N��Ϧ�ë%�>X�����Ը���=w�ظ+S2Q�
F�7��������~s�[ƿxQ��������iN���E���V2��]�6����73�L�n��3"�-�s�x�)��{ʛQ���������{#�,�=&[�K��Y�(��2'˃�/$�f�����2���Ir샆u�(u�}k3'Ͻ�ȵ�UB��1�n�qG�g�\�WU��9"\O�a_a�ufW�R��wU���H=�;��Q��ܥ���ic��m{P��&ꢜl��t#z����G")V�,[�Q�|�FuD��A�{�P������BE�Tn������BB�ڦ�<��-���;�X{�n��\�X\��
lUj�=�Η�ي���p�}Y)�PU �!t������B��!ڗK�q
 �.5|�3r�#7������b�h�؋�ν�'sP��u�h��hWm^��Oa]�h�� �����w&
K������0H9�"l�W�;�kA��D�gz`��a9��~��|�Uek�r���-c
���W=��Q>w`�b|�Ҩ��NTVA�����Q�Yގ���~dq�4�&}ds���4T��k{����ֿC�e�Ǽn��c�͸V�n1p�4b1VG	�v_��	�k&��Myr�>*���G����{�0��E:���1҄��/޿f�T���Џ	����_gd�;�(�*�΍�\}��龩��se����%�N��uGJ:�b���R:��s��^����xE�Z��`yu֪.:����L�;�rKx�z�y�^�r�j�}��]Oy�B¤�;�V}��t.9�QL�Y���'Sネ�s_-�!�%,�{k�K��<1���&H��롟]�6W���5y|2�-���9��f(�)���"6/��huy�q� Ǧm��HJ��.}���싑�OI�Ñ��wU��^���ԔoG�G�޼��$�<�yA�{njw!狠N��$�Fʐ�7W�T}(s�n����ma��&G[/y�;g���@���.�˄�,}S(�dx�*&l�j��U�J�~1��=}��A��m+ܡ��8M�{�KeFV}=��o	��A�� 6��ý��ݛ�q��](�g�GY�ۧ/@����t�`�om�T\N�Iv;�Q<�;8�[�J�+:⳨�X��Jv���^���w=t\+�o;��C��ֹ���]���y!�T��|��t��
yo�en��� m�uIs�Z��AgҔD�������iD�k�筱���\�
�0㑟Fb|������ ����0���Fh��M��l8o&t����Z�z�y���*i>*�X=�f�Ly�,*�vl��ADչ��#�j*�U�.��<�"��Z�En�˧0�u�<q5�����	���b�������{��;��p��P-Tw�^�bae\*~R<�9�dX�}�x�xs�1�F�x����n�Z������~/���k�
�v��n��b��Κ��Dͯ40��&�Wċ>���X�d����>��fk({i�m@�&(K�	~'/�Fga�\��:���?�]UAv��������#�0p���S�b�����V.p���w��4��{\@,l&�����o�F1���{{�I��\��MEPYs5�ֲ=b�5��z�����,FUt��b��6ة�h/y��S=̅P -�U,C��{�H:������_.J��aAϞ���ʐ'>̮H�QI��^���Ƣae���A߲B�w6�=�;���ؙ�J�#��q��]��x��%�tG3~?0��O=2Aк$���9�������YU��qU2$��t�t��[
�3@��6WVS�^=�ڞ��v_��2d�� bV��%�dZYo���̏4c{Aq�%)�#����8e}�e	7�T[�+ԥ�E�T����4�N��n����xx^�=�y{����n�vpy���9�u�(W���Bb(�S��[?�n}vD�o�zx��l|�O��o
�V�e�ߣt�d#6R��=���.*��8��lmP1e߲���-zձ
�S�9���bQ�� w=Q���ty?�z���|�������ފ� ۬�/�R�F�0o��{;I@��W1�{�⹼�7���^眱B��lz�ZG���e���1z<\��TR��l�>6�KpKHX�z^s�&�NWG��J���Yr6��d&N�\�H�Q�3T�9�`�VY>��V�;EOg&zKT.H%��Hת��V_?��%Y�0R��|>���;?�l�G=!���O�����o94�j��߮�|�d�AIȫ�=F��%�Y�KM�cF�H��l��H���
�}���m���ǳS��2�0c���w3z�M�,2yN��Yq٢�'!}��!�s�ٳ_��&C�+؄����ǡh>ފ�������v�8���ll�����R�B��k�g����3�?P�9Snk�&ͣQ�_��0ES��FE�j`��K�n�J0X����L��CKӞ�g���mV��0�2��]��f�J��S��+{ y�{�t^�r��nr��EZ����YJ
�5:���l/0���ZV����Wb�|3,gTm�3'"�b ���U8˻N�g�lv���:2��T��z��]�d*�,U���Z��N�"���6�����N�-'6G^��׽�����"���9�3�-��U�O�
�=w�z��K!�E�ʹR������+�f���M��l��^"Z=��e�V�^��Z�li�p�'��z����g�+=X��I/0`����T?��6�{��{���+�:.p����Bv`[CXN��$m�˹���J��ʄZk_�%�Mi)�G�xVw	�BI�[�-d��}�!	�Z��__ʊ�)!�~����9�IoY���b�:�'T{/�|:\$��$�����a��W���E}�^��i��z3nIˬE��]�7��E��`&�|��v�S��YKi��I��[�Q��suyo���%�>z]���)��
���>d��Z0o�
�<m_PN>g��ex=�H$��	�|���TD�B�TE���瀈`�Ț�hтmǶ5I��8d�0��W�&V��1�i����C�ws�@릺ϟS����͎�o�K�J���a9��05�RE�ݽ��EFNWs'��8�,LL_��M\����D�9����9��ۻ�^*��p��Y�^5<�c�^�4큎Hɳlb�\h+���{��e���.�.�=�V]M�ݍ����Z���޾{67��B�U��w��G�F�	�þ�X ܓ,�1�	�xr�=S��-휫�(�KtR�`�+U�WCBw�;U"�wX�T�ލ�DN��r�v_ko���y�puL�������K:��c��v�	�:�i�̹�2��]��D?牢�0����	�wHN��/�,�s�v%�ޑ7u=׾Ou��R�|Q�yz��e�<���w@��a��p�ܑX��#�+	�3�ҋ�T ��<��½۝���eZ�D�a�uY�y�j����<c<�,�)��-��:Q�ӕw�MN�d�9	tz��.(��(��P���֘F�;���|r�T�{�0c�uv��{좞�߶����1��W�T��\u�
��4p�=&gG�O{�@/�.��[=R��ȥ!��c�w�`Q�vbRDX H�p���8O��ҡycb&a��kj��3j��zp��u�S�⊔�i�
���枉^�p\���e�^���}�M��Lg�,�?�;��V�z�ĽN
�\5�������o<pKX�@�3�G����f�B�d��ڀG
>LC+zOI�޸�@�މ�s�"i��e���>���}��E�Tn�/0��ρ��ݔ ���*����1z"Sȇ���n
�s,D1�\�q6W��`��sY��ԃ*��L���W.��p�l���FF�� �d5�HOy)��7C�UT�{m0�n���ÃX�����,`��d�v��n�z�vDj��욯$áE�݊����eR=��;Y)�[ދ��å�¬wjO"#:�-g�D���SH��o􇔵7;ϹT�|�Ǒ�LV���T�Ξ��wќ��9�޷��d d�z=��ě�8�;��7v�T��������t����c0���f[X�c�ګ��-C��҃���fb�ߑ�:gf3�u�����;5ןedy+�|̓�����]� p^�*�-�"n(�YG�h��kdM���[7�\g��mE���)�v
�q��9��V��ڳ��H�
}����+��j�.�r��b}�n�L4�K���m��j_t��p}�b_�	��{'m��N\a�k��M9�QorƯ���(-�X����\���}�ō��R��H�o�)�P9�#+��[ �Kۓ�ĸ��tbV��>����+�t�F��j��G�׮S7"ջ�@Ɣ�#e����t�ڼ�Wh�u)y\�`���zhKi���n<h��R�}/z6��*�Ц6�Q���M	�1^�_��6�}�~�}���T��nt�[��.3�%�;'m]Q.3A�Nɪ�[v��O-���~�0x봠�q=�>��Ӥ���P�X+��=�;����4\�А���:��X���"�if['�q7�P(���&bZ�S5=��R���4�tު	�ﱷ�����q���9N�')gD�w����s*�ROY��<U���⫴LN-���q���o{1;�I:��U��JS�<�����P�ѽ�:�LY��m����LGȼ&���WE�_d�Aj�B�Mœ��՟��>���(�)��,�n�곉������?VcS��|+������o���}/�J�#�W+�/h�U����E��)�n����}�7I��UA�N���V������_YY	�8�;O���t�L�Ɋ����Iq2,�g��Ժ3fp��]jc��JU0p�U=��9���9�I@���N�p�02��sqE^H�7�G�~痢C-��-�$;1���{U�rFhUH؈��ai�I���+�a�^�k�/��;FZ�E�
��k8l�>���;ʽaH{������Z��1|��=$������tXت��]+��}o�upuu}���ò���G*D�z!43b\0b;����j�6:}X�A8���(���T�6��x�p�&+p������zӫ����C��^?|7���J���G�l�Ǘ�:%��{�E,�1
��'���+c9k{s���6wz�2�Ak}|U-�wܺ��K�9������3�~��umɦ���B��f�?�������<=��+ۗ=2�n���O��� �a�	�ލ��خ��0x)`������e���;+�E}9�쬜;�B;��F�tG	r��-�+"R2��N�X�eL�CiSZr�Y"N�ׇ��r���^��#t��⎫*��t�9ԭ7�&��;���k/,��&q[�޹Ţ9��:,���a�C����e�%��Tt:S�[~���p�Z�ݸ~�H�u���ο���ɻ��K�7
_!QU=v9�u(>`j�������ۈ��7e׿^�����<}��(鬽��ߟ�ؿFiW��m�q��8�~���~:�{(l�Y���W��.�/������n�v�}���r6e�6K�l���b�:�<������^_gqYa���C�������w��l�i�'׻	��`��k���z�{F�����w�yaN�&��(8lm�)[r��k�X��]���չ*T�ke>�xM_���ǇN����伲�����D9<B�|y�=��_v��"�E���%�F#�q��o�ƽ><^�tb�*Q)�OWVe��0z��EF؜�1���{���6}ن��·�~��;;��� Ͳ���>�~����A5S�}�c�x46�H�gWwO��'�7��b�x`s3=���zc^:S��VTglU���)�( �ݢ#�����^W֤;��iY�PQ�B�g���n�Lm{;����<7�t���Q_Ma1���oɉ�Cޅ��s"c�ߞ��K���Aݤ\�6��kx�wgg]�X.It�q��X[J�VrM�8;��c�ҹs���h���C��s�9i�r@��]�j��>ddYDe[,��O��T��r�0�y��y�ș��gZ�0���H�����WzؾS)���x�!�Av>M"�p�j���b-��c;Ruْ��BѠ��v73����:
^��}ݪ�����>�m�e��~�2wb}t���q"�t�P��٩�K�̬�*�Qg6�{ػ]����K)̔���yɒ���قЂ��}�wE����5Y�����*V^ft�����)q8b]xj�g*�4�fj�W�,�˂�9�m9p̃"D��sB����S!��a���jT	�#���K��A��utxn�o��|hNM�U��E����9����D��u�!�q;�Y�N�G��0K`5�GZ��v�Z_���g:H�Q�ס�n�w8�k���1I��>�VѽU�p��w�Ef�.C�G+]�Co��ه�����.1��o�%�.&���\�󂃲�˩���U. bR�.��A��$}�3q�4���AA���-^k��=�&q�Ժ�ݻ�-l��H��0����#P@m3L���{/�<���8��%ƻy��+�[0	��iٽ0�u�#"6o��U����M�����*t�C�eMkB�_r����'\%m�#��M�(I�/���/�(y����G%��r_pf`,L�|ő�֠�
�?(����Q���Q	)�������ŀ�*�{l�n�!
�q��S<ś&�C,s(XƓ��Ƿ�}�؋(j��4Z���M5����i���:1���Aʬ�7e_$�R�;� }YM^u;��R�I�d����1�v��_@Ս�Rݻ)n�\��|y5}��V1�ˉ1Vn5��C�ƨ��C�si���b�lq{�ڊ�M/��h�7H������X��}��!wTĪ΋-d!s�e�X��YǨ@�޼��R�%N�yXp�`�+9h��:��+��P��#���F�* ��dR�Bro8Ұ�X�3�W@	��8�����N��Y<���Jv�y�fU� Т�>�3�%������Q}2��@��;j��+�����ۍ�}n3�pqZ�v;N�
����vk��!л�:6�P�W�Lc��k#sL��N��v����Mݨ���o�{iWra�xkR�b�d�Ļ�G�&��͚��vv��3s�͊5LV�����ܻr�x{0wz2a��JI��(��K�<��݆ˎ٘�.�N+�.Avjҙ��lT�Rx�k�7-RjT�L�mǯ�Mb�<�$t�W�!��]w����㷜�Lik��o�u�T�ۗ����`�r�͔������M=Hu�����ܾ��35(��.�'fmivmE�J�G1�Y;�g��{���>f�ԭb�|φ;���	��x���К������:�gP����sh�u��om(A|7�0��ps�rd��B��f>���s��?�G�����}w�lMm�>$x��eٱ���T=Fu�V��c���}������aS��}����m��I�7)�>��@��!�I��S�¬p.��-e�虇3��x���Yg��s���H�cGDu������e�+#}�c��J�Q��l�Rj����"b��Fy,�`3��+#oo�/e�ժR��_��s��n�ʝ��T��eF�����Vc�p(�tV��F	�8S~W�{V�[�Ih�����su�P3�>��tl��־wɳ�AP8�c�'Z<Iu������7N�X�OW��A�Bk"�����@�����8��u�0����<V®U0oaOn���w�w�FfB-�m3̃�˲�ů��CLЍ$#k}��t��N֊�sr��٫c��HZqW������K`�4�/���k��sЙj棉�,&�}u�����8r_�^U��������>ʍ݉�=�|1v*UJ7�n���3�K;�6�������۝�VZ��K�^h|���:v��JlZՑ�� (Y���� �Z���G7�k�S������uL�H��e��Ӽf�p�)�WֵL4Zɵ;B���P��U
�H�����F��ԙ>X�`����g�{�N���uica15~2��~ʎ=�U����MUy㤷���L/����8���g�i�(�x�nb�1=�8�V\i%ߪ@�����t��^rxmOb�:��5���O-�D�>�]$(	J��{֫4W������%?}j]o�I׫���_���q�\��ޗ.�ǖ���m�s����;:��ϐ��b5.�񞱰/˘�b=+���0t��f[����Ue<�K"w|��"����ӕvx���r��Q��v�����zaiV�轼���O^}��mGW{n�;��F.1R����w�n�ް�͉$�R,Z��3>��TL8���-Oqؚ����V�;��<�]�v�͵��:)�ڊ5o�� ���2��/!5���&֎�M,�M� dy�ܧ{ݱ�ў���i�P��Z �-0;t�Y���<�#U)��gͪ�u��}�T��^�ۃ�y�dl��h_��#�?�A������[gK�,
��Z�]Q��7GIp־�x����x+wZ๴��5�\½4.<�.g��:�d��5���8<�C��d��E�7�Y��82���Τɗ;���/-NM�����4�
���U��MˡU���.�?��:ؒ��e@�������+$S��|t*h��� �.ĕ~U�7��F@�t�'"&Bj3���F��)s �Ռ,F�B�TXsO���9�0OYU�=hw�3��t��F�����P�.r=�����FR�S�A]bt���t���uҧ'#�����d���N�N:�~(#�"�g�q��:c�'��_W���Y�rǩ����U�H�vwh^���4�.{W��:�f��l�~�!���6�j���3��������u<����F_�C��0i�|r�Fz���'rNz�!��~�b���7����E[�R0n�c��~]L�jBd�-�t��ő�V�b"0M�OD��ǯf g
E����VG�?WO�f����k��V%�!X�c��sz�H���T�3��w깇��6�bٕ�rQ�ę�p��혠^�R~wZ���+u7����J��)r^�箇N���/��P�o�d���潋m=�ߪ�y��5g����j��ϓ�]+̧�n�>3�t�����v8N1���k�L��R���K�����j�>��S���;�$72�j[8J5f �ՂN!Q]]m��M]��l��v���j8�D��'QM�)�;���/E�`��Z���"��]B��XC����Ι�����-�wq��N�^.�7~�E�ZVFܮA�����7���dnΐ�����&�������ݕc�%�o��=a��ُ�7�*�����\{֖E՟���X�ݾ�yڷ`�P��W�t�|�}yH(S��1%���h��s���0��ɍ�W�Z��Z�<��ʙ~_�{й���X�&�pT�`�ѿ?yl|kyG�2�*c���Dn�d�^s�pt�b�9zieCr`L7wf3���P�Pe�<�����W���8E�1�2��p+�U=qtgo����*�����h��z�r�1�7�uBD>\V���Vf�谶���&��d�w��ޛ�Wt�	���Q��R����,�ر��]X�Z#<`�I0��.���G&0FK^�w�4�������8�K���$q����Oy:z�gY��=����UD��StK畝������]��]d1h"�X\��U�cf8�h�ßewY�-���E��=���[�ׁ��*V�-v��ͥ�/��2�Nm�D��m�Tn��|}`��4����f�_�J�n�(5��w��]S��;[C��C���7m�Z�t��kuY�p�
�pw`JO�&��{��1$|�����BNjg9���\��.��q��y�o�M/O�¨�U�}O�J9v���_]�f(B�����`�w�!�a�J�a�����e�<X\r��_.����>"JX��.bڃ3�<�g��G�U���ڏ8;C�����=gv��Ve�W���N��.����G��!.�h�`�ftr��.ڼݐ�v�Ywo�������9��wX�~���P4�vn�P�ȅu��,R�Ao�\�d�w�fZ/ҕ8�n����*�#5D=KDP81+5���e{����q��{Ԑx�=`����s�e�bɯ�K�N���{z��5!�WS��LV��x���6L	�7\"^��%t��V�j	�(�����8�V��?Z1�"a�;P21���^:�;�ٚ��lvZ��ٞa���xXL�x���0���#������d)���"���9p�}���)�)�Q{x���'�W�k��̺ʓ�˿�/0#n�N.��3W�v��Q��}��:pQn�;f��f�u�xѝ���������캓qS�i�tCnGL�����V��eiz��'��}ݨˬ�ԧO�J�X�ؗ%�I1�1�p����ծ��mʏru�L8��`�=�i<Df�k��\u���#y[yb���c�mq}+��)���+�~�f:�Umds(\L>t4�ݬ�~b_f�Im��_s����E�����s��O:=��+Ζa�n)�߈N��Ǒ�)��=%����z�%����Pe����籷;�>�#�w6+��k���5P��A���s�:�r��G�7�p��L�"�-kJ�W˃ �-T�þ�9������_J�;c2Z���z���r7��=�����ͫ��.�������cC����~4A�����E"+D���v��/p��:b{��D.�a�5~(�U��|8'UUUYOӷ�q�1�>�J��ډlķgDY4�p5��<�dꑊ%L�v��=L(���~�|`q��p:y�_�lï�V�\�/�a������F��X����� ��C���q4}Uwzs��r�����&f��p����mu� К��Y��!�ez��U��Q��p�U�6{&���]U:��a{ZJuØ�z��2���pJ����/m�{��.Βt�sϛ�CZ7�ͩV$U�փ�]�5*���`w��D8�4�ݷ�x/ɳi�I!��ݾ���-��K�:��r��,�۝+�L]��U���4��>Wa<����]�ֺ�[�Z�pzMfo(iV���ﺽG���5�~����+�>?]o-d@��U�����Y����it�I��>��H�4.A��9r��xCx;�B��FOg9x���w�9NQ���=Ts�0ힿzf���^�!_rЫ�wp_P7�J��mh6��ϧ�gިh���27���[c�k�o�:jP�'v���~�7��J=*�������QJps��S�O�RD��uq�0fnN(4Oـ��dЕ^2�����w�Pʥ�Db�	���h�w�LY�4}}�c�79t�lբ/�	u
�-Թ�9��������P=���դ�s$0����[y�(h�S��r1C9WA<���H��J����T�lh���f�xmY��Eg����WWH�/6X����/oc���M�_/��c��U�S����Vu�8���OW�SF7��Y7��Y1ѳ}kV,����3��9�Qq7#�< ��YG�њ��D��^�*0��X�Y8����ݺ>1�v�a<��m�%*|��y;�Rrz&�V�$��ӓ�;��`�b�����ؙ`�.3r���J��<�%��\q�ʓT6��,g���k:�l�7� �3]�>ζDA2_Z�k�vm���l��&T�j����>��e(�y��g�4衙�eG����n�f}~[S���B�x��$fw�D=�{V����G�
Qή�c\vm�>nՉ-T�5�M�{|�Y���`��}�<��zٛ;��a��:dJ;�v�YuE�^��F����e��&C�^Ͼ����mR	���
oV���AG�;�&�CM�T�~p�����y�mfUN�jo���Ҡ���fЀFJ����c�iW��|5x�����ۃ_%��8k�D���<LKn�ϫg����Cvбq��(9��EM;�+|Ƿ��������������^@N#��}l�^\����V�>�V+K1s�"sj�7}�^t������5~z��g�W�.�ǫqx�
��뗞�Q��!���b����k7���-��Zpk��#�l��ƿ~�%CVQZ�)��ſ��Tl�G�5M5�9�.�S�����0���{�*�����7�+9�Z������0yu�l�]��UioLYJ�8��k硍.���a����B���kI�;���w�ڨ�aC;c��ۚW�bn��*�p}���Z'z4�q$�5.v
����Z^�vf��\h��҃9�f�W,IB��k7�w9��-�Y�&�N�qQ�t([������3I������1oV��	��4��������_�1﮺N��Q�H��z�p#�Nw��{3�L����D�\�=�o�C�GŊ	:��0�����Gch�m#0�9�l�B^Gk���}{���Z���FK���=|�z��s��,�bt�7�9r�z�OT�����pKM�^`����J��Ǜ��S�|����j/�2�,����S�L�t�=�\+�)Z�ٓ�Pg�C�o#�
�n�m>�.����;Alה+B�j
��w�&��`�QV
��&�ub���+��W{&4�zOA2d�ͅ��U���y{n��p�OU^����_L�#��HvN�z�GG-���G��o�M�J�;�
�������3Ѯ�q^�>Ϗ�T�1|g����S�^�ڄ�����Wp�S�1���(�C�9�0�B�+$_��d���X����W�T����6�{VU�����]z0��ǋ�T��p�R�>�"�E7��`�|hG��ڮNうk7k�6��s'E����Q̗��p�IK�Si�[E�� y?X<p7�����F<D�	��02$C�C&Wd��ȗ�
�(gc#���84���L@pݬ�5���������9\��F����G.tZ[�\/�4�N�������0ty���0��|�J�(k[\]�f_y�����+|ȼlx�^�N�+Y���ڌ��ͫ��_��N'-̨�zz�-)�,R�zM����*l'�[���<bOEBô�{Y��K��������[{�KUTƎ����f-���jW]g�)*~�g]+�P�$韈�ܠl���E�P��豗ȾN�+{��W��yX{�u�;�Yv���O=:͡m3�ķЅ���7l˵�^�6�&)%�ay��G	�n1G�ܮ{���g��o��NFW3|}{�Y�.�I0pIno����m�����6�y�-�zGf�>�<.�\f�\Q2��2���o�n���ޭ���<�����X���Ό�1S��5'%g��
�z���j<-&�PN��������2'p��9�oe	j3��h��P��<N*�26*��Г�[�pfB3.���t� +{/����gu.���Rb�Q�#��6�b��::�z{*�އ��XMQ+�6���������{�:�}�[���_b�).������n��f�Oza�����n���&s3�޼���}��Z�¡-u�}����v�[��]�����Ω��?���<4&MT����Y)�J����[����Xۭ���ⴶ�+y>(�r�8�B���=�K�aV��F�KK�1�N��4��t���J�b���u`�  *wX���6pz���ȭ�!��VwI��� ���F3���wUԬ/$J���iR#�X.б]�k�3��h�շ����ѳg���m�E 6h��x\Cf,g�Ҹ�w���j��Q�Σ-ꘞ����ؗ7�i:���,�	�ք&��N
D��1���a�}���D3/�!j�����3�,j/VN����{��˃�fvL��˖�I�mF/V1υ8��Yy�I]����i�������z�E�Ӡ��I� ��x�xj���9�7��X���f��y�-;�i8C�-n���\ˑL닋�f��۹3{�ȗR�a�K�ga��AX��x�*^t�;L�@�/zv{�����L��ϰB�z�L�8Ԑj��X�����V:�n�9B�Փ枤�Q'K�u�S���n�s�����������@ۛ��@a�Ήһ��q�f��/��������FWq��I��Z��;Cھbč�+Hl$���6�٬mY��bN�]�����oה��b�E�+��peL[����d��\���2���[�r󍚕�\�Q��Q�̓ѮvQ���BkF"�D�u��j�w鈳H"�U	y:���)7Pv��U�K��ʻ��"LZƴ]������}���j�=�V����0�}g���*�E�:3�j\���]H@�^l�5�%�޷!���sg��Uc�ev�
T�TΥc�z匭�j:�dz��Z�r�+jظ�U�au��2�s!�����@�sJTL�q@�PЂ咱p���n�?]��������m.��nأfȓ̙&^���iu
�j�w��U^�)֠f�G�\�^&/��ӹ�F@����º]��M�X�Jz�^sΫ��\%���c+�X[aM�Y����Q8�HY�1�bv�T�����>�3i�ec�z��2d޼���gm'�0k~��W�󜻜{VO5*��i ;y:��5���M_oJ̭G:�Nۭ1��i��Տ{��r���3���b�Ӗp��8��Y����fL�uu,g�<Ǵ*ψ��Q�n,��n�u������<-u�옅�\��S��p���o Y�.J+�m�k�*��m���T�R�hh��֮�m�j�8͞-��=�@�+��5��p��i��4SѪLW�5���W���R��O�黧�9)�[�Aʌ��&E\R�ob�vtW�Jϗ�n4'=�)�M�̄���[=''�׬^�+��B"�6��Ό�ǳd�	4wP�i&'����t��@�RO����j�IB�MV��K*ɦ���Z�n��v1������|a�γ}��x�q�W�X5L�1]q��R+R԰8Ϋ�+m�e�ϧ�$��q���^o�qE�h�3����77ˮ�Юh�05=SHa����
��������"��M��ʡg;��]ػ9տz��N�F��{6����lNc[���6�'���_]=�|$�)_�g��<���6n*"���N����
G����d�k�*��c�3]��\�4�L�+R�7a��]c<���(�K�Wz�Ș�6M���ܾꊖ����[{yA�Ṵ����\���1qm_������߅=�������R����j��'{|kw6"x�j9�W�_���{C`xLw�~2 ����]�'栳��d��纋������vsb/�����o&�9�{�9�{#i������m�� %�b)Xhi�9���z���>:�{~(�+���5�Wη��%"�����[ ߵv���$As�+^�T�������1#�~����vWֹmO9�W.{h�NÝ2�D�]��QQ�*�8�i`�H:��M v[cX*���]�~�؃[8�\u�`��XoTJaͭKYW]�ep�ӎi�h�t��)�^�ȓɄ-a���� �r+�틮�x�%��pQ̬�/�,�~�B�6]�ӵ�����`Vॆ�e�@�C���t$�CN��c^NE����U�eβ��Z�}~����6��=.N� ko��s��]�G5� 芊�ػ`�\S�D���/�$)�MO�ۏTl�xd�� o�c�s9����n��4��V���4��{�,�����ҭ^��{��=^���ͱ�(���c��](�k��[�1�t��E��T�'��Y���J��Y�rAH=Ɛ�g�`>�r,�G��F�!)���q66�f#g޷_x�?N�.=���L���˝��|qo'��w�Fz�(�}ҷ1���3i�(.���ܶ���Рή/y��������}��CB�D�f�S�>�P/�(��W����@�&�l��/a��1Q�V�����gg*�ՅxT7���j��\R����*'·��M��a"r=�$)[���^Y��(����	�����u)�97n���Yqz���zT��ɖ�Wxc��;�9�uu�*f H͝/bcq8�iŝ3q>x�AL�h]f�U��wUӑŅA[pq�}Ζ��"?,������V��C���fH��MY�&�:8�Bnz���,"L�t��^�{��,3��݌{Ϻ5������?�@�18UL�ɎDyva���k�"��4��:BX�=�K�=L��%mT<�J���ހ�_��䀹���ҽ��>)�LO�Y�P�)𲫬7�6p��obM�n�3�=�!�Q?�A���7�C��A�K�yQ����e�"�5�=랷Z��gވ�z&Gyh�{
mlXݺ����=�#v޻C3�7#$0��v�(S��1Z'ڄ�}��d���lI�K��#I�>��q��lV=����Ѱj���zOE�2.�q��튂�c���J�5I֗����Nc���*��U�(�I�w�o���"������H��:L$) �yu��`��$���.��>
'j�u�;�#gaQO6���{��N��{g��	���r#������� ����s���;jbm��L~�_���=�vuF�Z��}ਿS��j�Ժ���Y�	|�vy��.�S��� /q+�o����k���^�υ�f]kw�ȍ�=�d�o�|v1*sv��g�)��$(g�E*�默����\f���Z�Z�{�xHR�=��b���P�o.�oV�������ć���c�XK>�l,ꏨ��6ٸ�t����g����d�p�}�O6((�*#qM[鑢t/3�C�$B�Q�B�`I��|q��&����`A{��W8�����3Z1��pr���b�jMޓ#&�e6��d�`zO�{�1�����v�k�}��"{թ�|ϰ!Sy.���z&���HK��i�9V�Q,�x���'1�'�6�M�z7�:c�Pi�ރB,ը*��&*�w=�,�t��3�%����
�^���q��ɩ{��R�X{oP�����>�-��1�\�{�2�y	^�7S�,�WZ!꯻���U�qX��U��M+��� �B�W��~s��/�0-bkd�S�5;�c�*^�B��X�:��ax+&l�u㣃�TIEw�P�����O�C�ѻWK�)FIp����"�w������O�H��E'X7x{���b��_l��C37��������7�c�=ۂ�Ndb���n��t:���&HM��ѧv&���ۍ��>x<�᪽��{����o7b�[�S�S��s������]7%_o.i����z�.�bn7�¦..�!�ʋڊ��T�2R�%��c�"���P���>�!pW���K20��K5���f������{I��e������i��i ���fc�f�����VnP]Ү� jF���Ef��������pc�����tn+9�ސ�{ہ�����t:�Н�0���r�c�݂}ΉOv��N����풟S9gz�Yެ��)�����~��Z�U�U��Fzgj���EgB]ھG�s~�������O;�G�x+ȮS�s���<m��5�>d�����ߒjk1���N�2-~G�EG�J�T7����}Qd�O�P<%P���v��Q���z�X��U��!�n�8ś/^,���5mf���Mۈ�^��(�O׍��t*�{�	j��'P���z$/-�3�S��p�Tv��m���Q�c�Y�
�Dv1�Խ�P�b���t'����$4x{}뛁yd��B�,_�|<Ge=��U�΁ہLh�Sƻ�&�>�*F]׷	9qe���}�X}Ǟ΋�)FNz=9�>��$;�z����o������թ���i��}ͩgj:�4 ����{iFr��t�V�V�d6�`��Ǹj͹V^j�R�
���׉������֍|�,V����h�H^���Zup��-Ȳ�����!���d��ɡV�ih.�,��»>>�{�wˌ�����֍�q�	���y`ڷ��8��]�Wy�y�;���Q���n�/��H]��/��+r���a�W�:����_�Vn������^ު�>��(����4j���N�[~���W���u�bϱkOR0�&�����������"��e{+�Ȉ��f����ы��T2�l4���h�7�_�*�z�j}�����''���%"������ft�bѧ{(�`�'��*<;:/��K��`+3O�U�������{Qu�g������T�j�_���}����ݧ:�+ѣ$R��i���]�T�y;<J�ݪ��x�c���20~ܪ�tՙv��i���;Na����,�>�㻆=7��o3yg�xՇOЖ�|�Z:�op4���́@t>��:�[��l���_{xV����`����a���1��
^V��d$�#+	����-�M�6p Z�
�U�Q�����v�h�U�4�ֲ�s��0����K��v���!F��ʄ˷�$��9�_fǯ�5;:��W��bVW ��p8�g:��J]Y�͖s87F�z��ª[˦�4�2�J#x�=��wD�
���N���w��0�*B�_T�@��9�0W>�+9�p?{7�Lev��B7F��b���7�\�(�Ga!�1γ��O���ϭo5.�_
���i�mԏ[~�{y�6=�=�gm.�F����Pz�����O}�.0GR��0��3������&gv���&����e�H/#赔�U��0���]���B�O�#��.#��ii�o�}�����1C�v2K6lߦ��8��+
"��څ�=#�\#\Q؟�yQ���aQ�b�
WZ��@��}Q�G��3V+�����@��1��1��z��\��ߧ�����K��dݽUﲈ�G.�|�0�w�nW�;��ZC!@~�h��vj=X��V��+�W}�̅��ϣ��F��ZcӕC�D0lvo�:�T��vˍ�R���'��
�r=_P���Bo��֏v{uC�#�$�ڳhO�gf-_��3�#�`NZ`{���Њʟ�L�\P�Gn9�e�������K�V'|S6�ó�bE��I�w�j�v@ǖZw��I�S�A�1��CY��ڱoX [�3UY���=�.V�pwb�:MV�Ӷ��k;�D]�,,����m��pR0��vS�ɓ�.�e{>y��[��_��B.���O���â}�:5M���_Mn⩏p�A�Lgڙr�oCs���o�64uvQ�|��
�E�q.���52�U1�\����p�Xg����݈�ݭ�p��oDw8�e	�Ȩ ��*Dٿ`;۲��D���z�حT>>���']�����S��C�l�de���yKݻ@��p.C�W^�2q��Wǘ{��~��"c�LS GS��
�U|�W)�(�/����4��k~�}~���eWVP�6���įV�1������yPi��{��:�z*��`>��fĴv��J�Y?��Ν��6�d�Z�3�Rn4��vuN�F�g$�ƴW+Y��B)���Az&@���6�x�fy�^�����/�z������I����wG�KCtU�8vJ�ܫӟn��)����M.�8��U�����z5��E���vG	N����d�[�W/˞G���+ ��n�v�:mE���E��;Z8�Y:լ���4�Z���(�Uy����9:���V�3R\�g�f��3.�lδ�F:��]ЄV��w|H\c�����Q���	N-��G5�8�=vnne*��H��v7�p�W�֛�ڙ�ϵ��6����W���a�s�[�ݚx.���7V�v�"���o��)��ߥ�â�9�����y��yp= �ܱ.��ǂCt��� ��$��\W��	�z��@v׀S�5�l���îK�?(�{��׽��	0fz�\���<��ar���������u[�Sϛ�������-�m�! �`h�:uET�l�r0��.;4ye�Gkr6���>��z��'O��,ڥ����=S�h����2�|&���rg3��i���C�������y��o�D���$�X���yQnU��l��O�R�����7^��_R=O�b4�]��B�JS��f4V�4"�OUh��^����VHx�PU�O�A�K�[�qJ~���ہ���u���-5�n�<�ַ�YN�f�!�sd���`�W.�[��f�\��V��ȴ7ѻ�[��魾V}Q��ݹ	UT*�uH*8�:Uř뭌��P�/T毛��L�(�e�Z� jEz/C�VL�@��ڻ�x�In�N�8B[�� ȓ��&�[�1��7{'s��|�e`����P�M���o2�)c����/j��
&���Si��%��$�;��;����I�s��OUH�,��ʥ��rQ���PQs7�}�����������ڎ�^:^r錨��j�3i�}8����P�	���9yl&�z{�=�޻�)hZv��gaX͚�{0J�r%��T�zĲ��μ����1��$G�#�V
�{3jv��f�ne=�����wʔ�������t�̑��m���\����G>\��̋m�.+�<N.�V=O��o��7��e���������d�X���il�9U�ז��y0=��>9M���9"/b�++k�0+�)�,�O^>u�K�L�J�'rȫ���n(c.ت^!�TX�ppv@����n`z�D]�E�C���?D�gT���폼��n��9��V/	Ȩ]�#�5����u][	�~w�;hٲ�W���oS�<[����;�V屩|��t5�}s�<C�u,�]׏�F$��9�/2o����$L:�6�k�ޚ:�q/Uo����v5Y�*�O����m��)�_V:aq�T��W=��Zk�z�C����tff6����M���9K���5�"o��F6�N�W�E��;y�}�s�WDt���@�C�˹�%W��4��_-Va�;��
;��n���#G'�1e�i�HG�fp���L[}��&9��/:�����P��@�E��)�:�f�p����$���Z i�����@h0������F��e	/V�k�/����è(��J��������/��b���������fu��ں�)�.�58or��{]u�di�`i|�r<�(v��2Gj}���W�CdD� < ��>��@�l�U��*+�4�މ�o*�u4�w:&I���bf�=�;P�dӛUǳ(R�&Xx�0�2<	RBb C��m�P��Os�Ԅ��I"�%Hq�r�k����P�C���3M�l~�I$�,�R�!�E�wM�hqz���E<�&?v�~�;�}����.��!'YE	 �I!��浧3��z�sW�m�����l��H����\a�Ne<�B�
vح �V����w�o��ݸ� �Ci�ߵS�&�n�w��h���!�M����*��@NU��$;+��^Pd����V�fe*ޘ��������F� s٭ cש�u�Ǘ���3��?U%e˦N����޹;���y���Ciq$4�Cg����`l����ʕ\�GC�z����+��O��{����5N��5o��N����ܼ���o6��q���7�$;>�z�>�(9z�����&���Y���ʶ3�8�����#��S��X���=�ɷ�Yzޓ���P�H�(��IG�q#���@�2�뗼�O�@� ywL��H��Hy�a��H��>ef�e�q�r�GZ�i�!�p�$:�b<Ls����'X8��;��n%M���UZLͦY�"�C��n�=�0�n�@���$8��:�|���k	�q\:�I
���fV�)4�����m笓ڰ+"Ǎ���] ���P*>z�_nO!]-���X{���@��Z�c(�=������U ���}�	Yϣ��|�,�+VuSܵ�����8� ^+h�vg4:����b*��G.*X�����C�m�&�2, �SC�]<�����	 w�+4�t�M$ӥt�/��3��	' I� @�a!ĒB��,$�B�Hb�߾s�O��n�|��XծZ�6%��)�`�@cXJ�E̾��9��Y���8a�qes�wi�ݬ��LB�i������.�,Ѱ��:V(�˺�	���pT�G^p�a�/��\��ܯ�Riu�W�����f�r���*�C��*む���^mwy�9��}e���]\�q�(V������h�`���O�o�'j��-.���C�Ѹ��s��j�w���t��X �*�q�xf`	��k�6<�K�LK�b��E����i,*���.)���3�����k�:z��������b�E�AH4�c�Oe�ѽ&9���o��#�j�3z�=�^�t�5i���'�;!��33��z�Ֆ���q��m�5ұs�5{l��ө��.�F��
u0nhS����#�g1!.,6&;�ʼ��3����B���d�M*xV��V�]���R�Q����mb��s�M��h�++�|�Ã�\p��+��Ep�n����a~����h�:Hq�pw;y�*V���§��� �P�-]d\b��ϑ7��2����i�����8��b����Ln4'��}4�k8'�H�Yww��d�y�Ι)�`�,w&w ��4����'���n���fI����via��(32�x�U��
�m���wh�Q�����M�������l������
��'��Ţn�'�(��R�՚�����4B*�";�w1�Vy�"-=ʉ�r��#wYv�:�5v��r��=�)������x�R�ʳ��9�Za�i=!v�zcj|U)�|�弹2E�:���>.���l���L�-k$�r�>/о���1�gܜRz�jwF�T���2�s�G�!-@+�7�NO�ԯΔ+�`��,����`2�{:�r�~�q�W�G�{v
�8��@|��WK�w����d/��yӺ�}a���Hi��;&��0oQ���K���'��9���<��s���\g&^���:��W��T���gH{��ī��'��{yVhvnw.X�k�Y�u>�+�\F��v��v��:j�}G&S��9�*x��������Y�#G�Rt+��wo���zIGL��~�'�߅��9��lIй'�9�b���U���h���}P�π�mOeY6+k]H|�F�Z�)n+myd6�P�y_����YO�\�|���9!����Ps��q=m���U�N(ӧ�?x=!�9*���֟R�g��}�.�ށ�@Ʃ�h���l�g(�9o �B�-�|�.�7�h82�#Ӏr��	7��9gmËqJ��.��O+\���L�)�ó'rBI;��*^��[�Qt�7�Kg��܎���y��lR�1�e��[&;�?++V2��O!H�d9��}Y�&ɦ��$����eeh�����澛jz��z� =jr1ϳ:ٰ��.��W�Onx> ���T�83H_p��3!JN8��a�7�$;�*]8����y�m����ͻWd	��S�uV��nէ�O�w�O�1�v�m9��ŋ������C�*=J���f�u����v����7��<��=��U���{':'Gb})���핪��G�m/FfL�#e�뿐����'�~L4&t#�W\��|��A�;����[�b��0;'��H����Ҏ��e�IS7��<��u[<pcB1|�x�h�?X���i9=55�o���#G�p���!��7��̯�_Upރn��ˌ�
-G�oƵr�;d��2�ֹ���]V��Ͼ'Ǉg�c�v�1����v{D�I ���x�w��c���ѝ�8U��Vf�:�uxh�:�Ϻ�h�� �����f����pہ`㣉Kg�Tմ����B�urW�W�7��/�b���� �����<z@X�ykj�˓��@��$��+����K�z[���ꪭWX|at4d�%f�V۸%Mp����u�eC�:�\�ox>���Q޸�e�H�v�	���O�c��1��U�>���瘷:�[y۞����T�6V�i[��7Y���ۮy����D�Z�O:�6x^i�3���egj���<C����e �sRo++T���E�����g�1�����w~ǳZDOP�m�s,S�jdYxb����6_[z�q���1�V��Vo5�� ñ+F@�o�u?V���S���θG���Ʃ�y�:�����#��Q�Yt�Z��~���T���*�\:��5��&��A��Wڽ�FV.�!���aA�W�I����$�(�����=��9��h��E�i,�`zmh]�V&��y �.nMS�1���'nѤ"|�DXu)�+���uD�ݤ�D	�"�L��ޚs�r�iӞ��+�W�>����jz������}�5�PB��S���I��T��X.������}���Ɗ���0QM��h���bs$R�+BV62\L���%�%�5��)XH�V �����ғ����Y�&��A�#݇�MM.����̕��+3S������N�L�Y���m*W�ʸ�&�g���Ĳ��9ؑB5��٭q�Yb���^���!h���*h���Nez�u�Ƕ�_m��"`�[��Q�㦭{�<'��o�����+�=��#�O��f6�ę똑b��Q�}b��[���}hN�?L�X�v9YP=��䝝���wY�G����/E��2E���KU{�'ƵR��]���S��2�+Քޝ�SɸŮj����z��{c
CvhڛN���m��U<V�@��q�{�d��muz�3-�}9F�\bfS#���w�[;�C�w�Z=�c�ᮈ|,�1S���3ݜБ�m#�H�2,Z��;��(e)�&�T��*=�S�z k������{�v;R���9.C��h}�/�r���������e_JQ�rW�ۓ�w��מ��+�� :��J��
턆`Dn\kA�� ��q{7w�q*Ƣ|�W�����OP�;kϧR��Ӷ�L���;ϥs�i����*"�����&ڸ�{��������b�D�ave��t�4�"��$)��b6�����҂c�㽽P �9��%�ٷ�����i�ə��1��"�)AU�LSMw4cS��X�����^�ǷL����;�*����yE��H��G�?/LO��̳����I���k��܃�uF�����yT�3�q�,��r�&��J������L���^��G�F�l�j�7��	��ٶ�{��N�t�Q=匑u鄼eJ��G	���U����GM�0.�#E.c��x׺Y� �~+o���c��F�
;�)��.pWOR�T�V��t2L+"�FS���Z_]�U�7��A�e�&�j�b`���w���uV�1�N�����8\�9@��c�L������2�
��o!W��
=Oi�1�5ump����M�F�T��*P����אn�Q;�ix���b���ex���)b���tПv����U�mG�.����fJ�(��عdtq����cg�̳S�V6'�nuW47��
]��Q��끚��q4f�D{Wwa�ޏ=AS�W{�!Lc�2b��{�k@F=%��lo;��&����hͻ��R��gb�h�������Մk�.�]>��I��6��ĸB�iM�:�E�%�ڀ*]���dj髴��������*8�WZ�4˽�N�����`2�u��q�-�Mp&��ǀ��*�C굧�=�Ow]\VW�w�c�tW[Ek+V��W��,�_q�&�Fd���8)o��Ko��x�F�@٦���9ؙI����yμͣ�Cz㦊��y6�o� �)����tw����t㔪�W\���L�}�hdM��ԞCY�2���^�����}.�� ���J\��׼c(��G��}��V/'C�8˸�wJ��]{�1��[4j����]K��G��2-0Ϭ¢Y�0�ʮs���uL�WDkK�wvb�
����8K�툕;U_h j�@�Y��YK�b��K��xS�ʉ�TpB��ע�Tr�7o�ޠ�^oU��H�t}~�:G3�|6��G��!�x�����f_�8R�bP��߻qr���I�n��5[�*ںOc��^eە0�8gӠ�C��}k��3u�hB������snd�9�f����	���|JU�߆-/^J���t{�o�*�jM$}�����B�u��Z�v��s���h��vx�*��ߋh�ţ8q�g��I��r���Y�= ��m���ԱD�X�R�f��J�S/w�'��g-�u��E�U�ZS����'�b�w�;���\�c}5ʹ�f;U����+xg�j@�-��<e��'�͟f�2ACC�f)�8ت#��6�2U���~cm:�U}£\Wo�l!"��Ó�Z=0�GD����W�b�ix���l��d�^��zO��k�sQ�앶6 ��g�������4NA"|�o?l�']����Oz�E���3�{g���/.�D�%޷/T0��fb���B�绪�}�~�_^�9�7=#Y���>x^��j��3#bS�R��i:W[z��#o}�G�<΃�/b��wz�0Ęޯ���1���{e�����ۗOfi��ֹn���[�6��3�#A����N����M����:Q�����\�v���	�z�]��_GJ�A��'99q��0�Le�<j!��é���\��is ��꫰cf�a�=��hw-���D	�TW�M��q�}�u�Q�f~��;av��cF�`��+mlw\<H�YQoj.����D�١W7���U�ڸ ��ۉ��^қN9�]}�粃��DҎ57T1P�ZN�/��-{D#�B��\F�}v<"��F�*�J�������Q�[��\��A��Z�����2�ڶN��g����s���r�Y|'���E�?�d���1Qڻ�k���j��s�U���=e���;Rr��l�d5�p��N�����]��P�y�JGKoJ<W�p��Z�`ǋ�%Elz����f�9�kU�`��R�]r+�j>��A7Cl�^����D�)|�<��^cr1ۗ���q}|�K��Eˁ�r�:����)�o��v��:Џ�)ߞ�����]�f��������= �9��:�E�";�.s�vp�ެ�}C< SQ��V�����m	
�\�0�==ܓ���2�I��Q�x�6��*�uD5~�[h`��ds٦�H���H��������%��W�Ez�w�t����y3��b�I�\f<1�_�C��]�AA���j(����z��u�]��0J�;��+F�y���4s{�rϜ�R7��"�����n*�V����C��[�<b�;�X���~5q���ԉ�_��\F�_��ĳ`�8B��`�ҽ��O3W�>�7�0d4�.JMJQ���]|jw������ah�7����{৵��=7��a*Ū���S2׺��Mx�DNu��[�U;���,���͐:���p����z℘yth�w+
�W��@�ł �=Y��[��(XE�-�ʅ;&��y<����
JGd��hѦax�"e��d�}�{3;0�a��SU6C]a����HT���s^;;.�pK�L�/�0Z�V�UŊ��Iy�I7e�:����.�R����uJ�s5����I�Dޝ��j�{����D�`��#04OP��F�ל]�Sϗ��{WF��َ�f[Ӭ.�5}�&���p���60F���)�!w]2MzO����eا�E�K|$D�c���/Fr;�"}н��i	\�l���jZ��8��ڑ\��5�'��z��S"��-���
>��3���u�Q�3�����ӿ�o��pZ��y~��ݞh�)2�C;$���8�	�1�5"D���4��}�������n\�\�{^�U�������5WJ��\*$?V��0��z+,�xNi�8�7bTڪ��w��q�3�u���� ��%Z�l��S=۩��eo���'����6���.�AH���`�\�B]?l�����[�5u�QU))����:Lk=�1SJkR&�a�:��lJظ�f�x>���{��h�-4����ȟk�h�m��[�����d˃����2f�V��77�L����N���0֨�D>����5U�n*�_t��a�k\2�;1�n�T�ڭ9���h�]My�s���'���ī��!����{O.�Mn�ѫ�4����=�
��}i�8T1��Nv�����[�GWqO��e^�)��Gg�0+��J#��u���E��� rՒ�r���u�n��nܩ�E�&(Q݀s
�ܬY�B�� m쥦tXx��xXs6뻛)4^dШ�r��ۯ���m#Yiq�u{��}�q;ۺ���a]KsN��v�z� Ι��'ۃ}��=Ш���_g��ĥ���qߏ��Z`n�Y��!+�U��[���Pɚ����Ò�-p}�B��kxr�����
uۜ�n)��<_�Н�E:�,޽F��xˁG���ي�����iHd�X��gD�'k�<���u���C�}��LS��<��=�6=���\6�(>=��۔�H-�p�\��q���,@���ɾz��3����:|������O5���L>�z�H����[o3ѓ�4*�]8>�]7�����cwb�磜N#)��aL�
�W�=�S��罹>.~�Gۍ�C�k�n�o�6�pm>1Z�������ꃪo���~�����>t&�Dd�;��	�]�О��(k�D���=�����g��W/�}�*�P�=|�qk��k�3_c���Lׅ��CU<#1�'��)�Q�J���T�(z�UM�;5�sZ&��n�4t.���w{��Q����ʳ�uC�W���X2޷<��ݱ3'��r.מ�3���i#rS!TdTU���Dq�3�G��Mj�z������5�]Ԥ��\�ť^
�w8���������2�[��U��ꍱK�[2�ٓmM�F�p�"(Ie��'�sf�K	���^�Ã��Zɺ��Pb1	��`��	�wOA�Y�Q5a���u�����J�y�rN���� �{VX�
�U��+˗9�oXR9Ad45�E�<��E���FH0�\F�ֻt]X���n9W7"Ј��'j��QW�W%m�f��/_V�֛{�� ìo��bF�xu�^+����q���u0�3Aq�z`��^5d��V�K+D�@t)v����(�U�R��q~⡯�� ��+�v�� ��\�,\���A7�u��r*|뷳��'Wq�>�̵.��v�d��f�+i9l�{�χ���߀��8��@�g5�8%��o-���)����r_PW�OY(b���b�޳nr\�}�k;�Hm�Y	����i�:�G
¶5N\��T����E��d7��5Eb��A(��v0�[T��n� ,Z����꼹�G�Lo��+H�Gs�>�%�w.��"sS޼,f�y,?E!g���¹���K���4�q��'j�e�b�kVR���3�P]we���b���"�^4% ]��Ur>,P��s/��0]���NuH�z��u�����k�^SX%+���[ݤ�G���.�yXw��1�=�yu�Z\u}�3,ĭ�����_�\N�w|!�n`6 �i�[�*w	W�5�Z� �4>���X,V�����7�h��ǀ��wi(8��aȳ'u�u��B��Cs�t.+���1�P�-7ه�q��6�g8�92]�W����u��ܭ�V�'���U���'�#�d�f�Ǜ�&�w�%����bw�Ͼ��v�$'N2��'���ɶ@� R`	´f؀�ga��6�bӐB1l�����5ڒ��2<q����9t�`��%9w0BE��:P�0m'W�cv�-ѡs��Oa�F^ug/"���2�i=/^�]�=��j����Q��9�je"�b�{;����h��Nn��cvĨr�Fst�aΫ�*1Fl��kkӥ/����Fr�@��c�YUxQ��V�!�F���U�jEvX�U3f�e�׶bу�[t�i�������|��u�i��8خ�y�LJo(5�[��u�#�	����E���-I�Ug��N,��҈��	�1�[� `��v5��Z�/�}��8������Y�if�����?zSL�Ov,r�<ZT�S���Iv ��N����&P�g ��a�T��Mj+U>������T�f�\�d��L��S��o��M��r�GcFX=��D�9��!��O�qP�e:�Hv�J�ɍ��p��;͕�l)��1�*�U�TA�ϣ�-�Y�*�{	�U����%�J������[ݱ"h���e�z�;`Ӷi���m��v=��}w�@����&��"��X(L��]g�Tn�)ax�N��u��4�R�J�G�KVm����dT靤p��4o-N�`�|6Y8����5Q"=��Qq5��0��V�&�U����%wj>�!+�%XB�a(�*��X�< ���^�����0���`�����|;�V��-Y�Dv�/�WQ>d��Z��ı̉���f�O5˹����w7�7�0s�gF����:�[�n���SG;�Ѵ:A�����e���.�3�{ݧٳ#P�w�2�cʳ��сc�H�]�J'�F��;�tqD�Y�ћ6vsTe�ܽ�޷�<iZ2;e.\qA�5Xf0�&sX�=���s��U�N�xi�Zq�X�~��5Χu[�,Q)F�7{�lW��WSł�Y�R/.����x{��K��S���X��#��c��g*��{����s+�>k�xr�wW���H�Ѹ�;攱��1��S�w��21
	���\�|`\�(����GyX��x�O�޳|6�h�����ҫ�!X�	�}���J�E)ھ8K�}��&�mb����9�/} xt�?CͅօТ@�]�����7���,?�Ap��NF�mIB�����(�BG��*�/c7r��~�˷CLʃ�X/n�7y��foy��v2�*����3��ǘc!�-��4���~�Ӻ��3Մu{�s��=#T�8_�<��D�e��)dۻW�nl�7hB�;�̩Ԍ��op�B��.��X�;g��eAq�f#�8p&��%�.�6��s_e`�u,�y����a�H����'*��I�Z������!s�}k���&��p�P�q���y���mᬂ�i� ����f�K��\3A�������D�GA�.7��=���C��iR˵�v1f�s�W7���*�t�l�7�V�
��܊~��7�ށ7��f�L�J�2�	�����8.�l�ޫ׭�hȯ��NQ�z(��2U�ӊ��}Z��� �l��𺞿O�/��O{��΋���DU���#Q���(��8G)����i��u*m��,����s��廴<G�Q� ;|��~�0=�M����׎�f*��G�����<�Yg�YK��*����tҕ7ѝ�G"����0��&�"���A���p�Ok3s���)C�MF��;֧A�T�fwn��[������}nqvP�W�F�ڦFeO���a$I}ɣ�ى������^V=Lq�����������9��Z�Kvfo���mp*b�YR��{^ƥ)XH3����n*�\�����Z�l�T�[x{ 8�9ZnV��9�(3�&wB�LO�ʸ4�ω�1�å�Y����j�^�yYʯ�"n������0�~/O)����w����ٜ��H�;��L4V�ϻ����v���{�i�;\PtwV23]\U��"��½	��ML�*��Q���b�cE��8V�|g.&>z�܋��-61J�'t�!p:�D�;J5m��������Q�Mڋ���<�p	P�&��S=n�A0�t�'�۾Z�k��׮��s��1u*=6�f�j"vwgqA�ba�4�Ǻ�ҶNF�=��^�d{����E����N=�7�I�So�N�C���5���o�?z��B��j�x)���� I��B�ϱmg����+�nӹڽS�80�c�p�\�3�9d�׳�z�d�\�I��S][�6p.��P'<��^$�'V+q@S�9nsU"#У=��u�P9]���i�?a{��Z ؙ��r+ˤ�=쎰�h%�]mϭ����B�gֿl��W)��X:W"��7}�K��������m@8���׷^�y�c{+�^�Bq�Up(��y-a�j��s��+�Wvi�W]��/}:[���>/��v�3��
��y��@'i��_�*�#�K�Z�ڻ��끄ẏ�����oچV�
����q=�B�Ɍ�s+K�Sj�<����ѳ��u�X/e�7Ȥ}���֓y[v�t>��s5T��f�~��F�U�/qtz��8���ޘ�w����#�ɝu<t����V�����?��\5�A���c����a�.M��;5
�9Z�ta:�,�{�r�,Y�X�w�n7�"�۳��P"�b3�+s�I& d�䑉!\������
�^@�.�����8L���njA�Q�s�KҲ;���d�|��rw>�Ī���NCW1�OY5ӱ�E���1 ]n���0T@C��k6\�Sy�F3���l�/Ty
��u,{� {�.�1o�W޵[�w��2��N��J�W�&�WO�'��애�(B݀mc5��Aγ.���wP���Q��i��yQ�xx4�\&at罩z��pB�BX��:k�ŋ<��3�U��&`����4(�6��B�����O8:˛��]ӾP=��#b�̓�#<^��1%F{c�M����W��yrt�>�Sc׆�	��Q짊h*�[Y�Z��F�5�PD>~�FЍ����F��04��R�o�n��j�7�1Z�F�+3f�2:c�!%��D�2���C}�D���� �s���KU�x��V�_�3�i_��.#��_�#�'Flpc�r=J��=��z�o�-4Q�������Z��/�[����+�*��]T�ѷ�'�v�����{�ybrޟz7�Og�gSk�^��=^e�x�7�/1L�*Gu�y!,�A��F� �������~�M���eB[~�v�W��?%�]ahc�i�TX�{�����_�^���c�o���H�\������)vT:D��*��q)Cqb���foGV:��z�Obs"���r�yy���H�gY�gus��r��v��:d����*�t�R����s�g��yA����A��kL��p`w�&��H=w��a��@e�Mո�χ���ٓq���<�~�3w��\�-66���j=
�|��6����ϫ�p��/�ƃ���RpU{/ψ���fs�Ӄ,�|�q/=O��؈���E�T*�_���l���A8�]��:r���l��bכ���
;������
�pҤD�ɷ�f��}Y]��	�/.�o����7�G�����R*�d���F;��T�N��;�r�޾�'!*�q[��� ���`���I��G�NOr�~�)Uu��oO��mx�B��B��'۔�\i}f��0�-�K��.��y��jy��kz0(��k8���]�(ݩ�=kR���mrJ�q&ԓ>���s�W^�]~6���=��������O�����{����٣�U�ܲm��$~G�8<�D��]y�I�<��?B�vn�м|Ec��8Y3�d�����������#�s�YBHţ80J+���q���W���HA�t]�.i���Ӻ��S-�/W����<?]5�[��������U������gظ����5u5FJ第;��Dj�.�Mm�{\���AJ����.�9k+,�xR������l�6��t	�i/+*V���;S�&���� �sUu��BE������i���7Ne��i����o��镂�N�b�Ҋ�H��㌚!ij;#QW�p���3�8s��;�5<����K�²��lۦ��������o��gTX�:]�s��>o�x�|�}��v��+�`X�>�3�$�zkk�<��S��]�K������[��,�v��b��`�ݑ����_h�1��gǾ�"��}i���Dϵ�^Oۣ���5ׯjDl>T�Yߣh\�
*3ʢ�c*�G���S�8�1��%_�M�J��@�Kq��&`vlGH!��OyVX�$H��mFG��7��m�	.f�E�j�Rh����YKș~��kN����lZ��Æ�7����W��7(�m�Wm-4�8�����}��h<���^u,��"�a��u�ޫ�b6=�B�į�sf��^̿'��F��:ל�졫�U�Z�*$�c!�"���㠳Q�jJCطѽ��,�n����:f�}�~Ez��Mc���]��g;ۘ8���3�V�}�Ȑh�"^�>��0���+����˺E���RF]t��0.�xS]bb6��K�[=�<���8�J�5����xlj���~���V�5����kQ��5fB�0�;����G�w�e�'P�rT����]����hn�C�;p���P��o&`�ৈ��ߪ>�T�f�6�lBn&�%b��%S�%%�F
�����!��Ū�ga|��}��2���D?���1�F���u�F ��wß�+;��nV��'�f9����.�eQ[M 'ڬ���sSV�^"Oy��⢳,Uߦ�Α�.���h���}W63�}7�����ʧ7u�ڄ0[��ë}ٯL}�U
��h�������^Ӡˇ~�W9?p8�r���̣3��n�z����ov�Cezߖϲz���ߺu��wh��	3
S¡�v������˥��)A��B��^��5V��x����g���m��B�|IA��F+����3,\)\e�A��N_�l#X[�#�WE7�yz�v��A�����w���Nl����7�}X��~�����C*�֒�G����"sExV����Ng�c��]��]���\Y��O��ܮ��X�����3�^��X�D�X<����1�+TmB�����s�����Zݺg�	�g�,�~?9^�3;.��83W�d������!ϖf
�n1%<7��x�nz&59�����tb���ͪ[��O�{�.q�\����αru2�t>���ƲVTR=��x����;��s��yʮ�3u��y��m_6x;R31�*N�Oٜv���_1��f��	u>��]����Q����{���ӭk}9�кA[V�t�tc�+9b��f��dDv�Gn��+�p��y�|��|6�.�K�N�"x����zbc�﨩F<��t���%N�y}q�s6r��q��9f�:���O�-O�{w��}Z�G�e����k�K��F��x���!t>��z��q�!,�R�wE;��]��%wٓ�{ū�G����o&��'��?�V�-?��(���su%~�v�j�^��Z��Wvj���>YOӀ�`����ض%h�Kc�uQt`�ۑQ�KG��J]�!��Fz[�7�gG��u;�Qw6S9�:B�.�E�R�{�F�1G�f���
2��ቔ`2�8-$iQ<X�V��YU>X��c��|������d]��m����Q�!���I�)v�{7���m\6���9�=�����X�j�8���*��j���zQ���b��7�&��q�;�㙦�]��|o�7f�%�7��j;
����Y�!v�ir��w�g����{��]d��.O������~�i��= {�wvb��E�pg��I�
�J�Ln���^�_#�bb�{�l{OB�W`�o�M*�O�#)@ԍ��X�+=�T���-�T=�o���PW�=~����MBd�����ཆj�Sc����!�+��� �p��/o��}�>R����ݪw���
D���o��6'���9�+��F*����2��Z��u��![Ǻ�!��s'\�.	�:����_�X�Ϗ�+�=�	�8��ܡ�=��>eN���g.�W�J&�������^��K������~�5 {^�s������U�V��%Z{F��2+;��2c���
��|s�<W�(b��u��6]9js#�p�@��}���O�Nj�k(e�T����nɍ����08�����z,��H�K��5˙�<��d���ӆ�8~��f,S����6i� gǦ�����Ί�깁���f�=������o�YB�E
���������R�Y�Q��I��#8�*� '��5���$�ء4����U�bY���.ti�㑜���`8���gC��7����,ˬ��{
���G;�����C���}*�~I�˂g�O�N�ڑ-�8=7"��Lr�D�=J+������U�}I�*ǝJo���my�C���?%���ض����>��,:c"٫b�n��N�X=u��;����c�lg7�T���;ï(χ�������[�-������B�Z����S4�23 9�/��#�s�K�\��9K��X���c�)>�7X�A�n�C�0D|c�MΏdŮ��wXwj�((H{��a^�T��;�E`��q���e���r/J�ח*���%l��J�Z�Ɖ���.��c�����͊�{7�p�� 6����t���3�m,▷��+Z��=~�JW���r�Q6K���ޥYQ�y
���$�#��w7�Gu�vN���kmEtd��������'��@�m�>��k�y���s�虚G��W�J�~��	�7H������!Ěu�U�`�8*���(FA+��7]s��y�p�ԍ)1�-��Lq���iu��ɡ�� ����y�ѭ;6�lJl�&�kR�1���~Q|"ų�%���-flk6�����de�	����Z/�\y]GlϗF�3�Xo��h�mЈ�f�QҨq��UBD��J��(0�C��aL�>�7S|��]q9�9�%fg�v�s�Ɖ�	n�z}]���B�Ó&6��>��dI�}"7��U1LvC���u&v=Evx��fe�A\_�N;���L�Sj�eM�T�ҷE�(LGh2]e�k;!����n��%�L�U��og
 �DZ#&�t���pc�-�,Da��V=|�ɗD��_�{0r����4کPaf;����-��4�6n���ڭ�
]Hv�27ר�X��$��m7�g�� ܘ1��F�qe]2oN�Q���eKٛ�fd���Է�8]i�p����鯷����K_>���7�{6� ���¢�����W�P�$X�]waK,�]����D�;ʕw:���J�18�i�喑����4��0�LLz�uc+um���<�9:�#;@�+F^�5��v���pd�Qkw˧XX�AF�>]w���Η���46��[I�1�N�|N��H���ֱ�45�U��X[ٙm���uK�~�;���Y�P�1b��+�P�MRdSTs�|0�ZrKX���31&z�v��]��)y܁�D�N���y�엩
����h:��;�Ĕ���:x�D@\|#�#:�i��Ӽ�ݥ�u���]����O#ǡܨЭb�4I�I�eT���2�5y����T��YWlː�?)0���3,Z�}5�1�j�`�Ё�b��][�#�^�pd[��`%O����w[���l�E.��������R��m�R���1Q����c�����P60�JohV�;��`��T�r��J�/í,�i
e�R�0�̥�H0i(4�	f�x�/�7Vr[,�Lݮ�F��79v�ˇ��8�B�=�y���TN�݇�#mݰ��7�_9�v�\;��]ؐ��!q���1t�$�P;��\Z�(�ɚ�a�u���\�w0��@�j`O�zv�-��e�kcW[��VqX�z��ۻ��?e.{��F�롇b���ʛS��wW@���K��)�=�C!䠆�8:^W1)�x��9�#(WZŇ�c��X;��#\Y�����\Ô&���w'.�_t�նUp�ް�

�󥩠3�q�X��6��R�#"vy)�4d���e�'���J1sO-��ŊO+5�b�U���}�y�j�rү���tt*e��67fT�F�:��b��m�8@���|g8���|&P�$��3�O�S{
<5�n]����s�u���c��eT���p2�6��9��ĵU���ޛ�I��+R�/z�"��]�g��/���M(+�l��Zx���
2���!WHŘ�%c]�n��)��IVЭ+�L�Uuօ�]{��/�:��y���;�K{���BW]@��Xǲ�X�LK�u�ˬ}���E��u�K����s�Ryݙ89j��m,ؤe^�ؖ�b_�mٿ��ѣ����_E�wݤ�|��4��f+�M,w�%yU��{�"Te-`q��X��V�I�f� �x)&��"��9c���6c /y)��kf�r���R�ҫ��K%���P�ővu���+]��o���޽�r �����Y���M�2���66��\�������U��Gi�w/������; �N,���J�P�=:��!�P²f	O�����\/ �M2��*��Q��:R��]u�>}��)t۝��TZ������H%ۆ�|�$yl�v�A�;4E}��MQ�y��/X;a����<z�$C�>��>)A�P�wi2O� �c��=��ggr�vpз���NSm�:� ��=���V�{��hB7��YF�̵�`�\�GX��ز�s�	����=�`B���7�lq�M����J��u�K��nȂaG�n3܆��k�����ae}�\YYN���)T���N*#%h>'#�B:�z8����w=9Tg�KQX���<!��TՂ�Uq�Q���h�W6^�۰ژYS.pd����<6\yUgJ�c��w�}�F��Cef@س�&]N�˾�F�}�v҉>�P�C���SGw��mm@�9����\<�dLjK%����U;����Z�$yW���pěݵv.����e�5�a�5�n<\�|���؈pg:����r
h_��7��S
Ư\� z�l��LL��(e���Q�����Q>��}C��^s�e���<r:�XS"aXF���txei���"��Ը^�F(F�[�E*¾�v�2��׆�ԡ�����^1s�UDG����x:I����;e9������sɞ�Z=s�#!�F&�y�17�.�m]�U�z|*f.w:C��:{�{�S%��<NNE.�KE}�+�x���k�ՙ��4�S%��0\dXZ��ۭ��r}p��ټdhc@�p�dɑcC�'�0�9����68L��e��(=7s�٘ռ*�k�����<�_'�C{����1�j��(u!����D*���9{���2�"h�k�N@xd���y�����2�|R�֫�D�HY&ﺠ����� TΎ>�.��:�S���#��iݛ��b=5YQ�Z��S�蜰���zP��z��>�0b�=	k�ѣ+�=N��FWw���ɵ�7G�x��D\w����n�Y�1s���q�1V�Bv��S0}��=t~��ko���1ɞQ�x\g���^}wz��ͧ�xP���R�;P	'�.�m�A����~9�E�9{�|�]��}kg�շ.t���06�t�:��Ѹ׻M������|㡱.�Ϗ�t{aU�r<�W[r��VAd��sژ��p�bJ�!�����+���g3xK���U;�Q�Y��ި}���m���[��.���F��*A>anK��������m	8y>ܺ�OVS�_�-�aۡ���|���̯<P�����Xe��=[ZG�r\sN �T�6J<#R�
��+$�M�m��n]d��GW]�vk��'}F�U������x��'s:U��Q0��Ԉ��j|�ڣ�j��TO(�k$������idKC�<7F]��l�s�k�bQH'ݸ���p�����u��u��%ػ�\̔kvwokۮ`ߊ���պ�{ݖqu�V�N����UD�Z�^��6Ί��4%�ԸZ��x�c{\a�wm���١�w�C,=t%+�g3f�Q8���E�*����^o��Yv3Y��et%��"�j�C=:�lW��������W}3�o$t�N�*��a�/��e�C�(�f-6��իfFe�Llwr���_O
���:N��j�d����l{��2�k�E액�W4�eg�p� �з�~\Cx!Ƿ�N���)���Y�&���v2�t���
��1�kpӺlYk{OpM_�|]�z�i�ތ���+��z�^��)�Y�>�bQ3i�7�7��k�/�kK���&�ޠ�Q�n�'/�H]#"j�q�VO��X�$�v��\��@���"1V�'9�>��zT��jÅ�^t��-��S4�L�;�Ke���y�l��+6{��������]��Q|�Y����L�;��ӨN3lڐ�n/`���d����VR񫼴g���-w����ߨ��\�@��n���g<�	��UW^���j����Y�շw�I�J����5�����[2\0��x[��!�s�#��ו�6���n���HhpŞ�P4o�ꑾ�6s���.ղ�FZ��r��}۹�*r�����k����SP֭��-�4�ۢ�b�����/����ը�uț+��v�F=o��Ό�7k�B��9㵝��=
�2�PZ���.;Q[�Wd�e^����r]�H���r���G�jbE��e®n�j��{�Ǥ�^�=�8r��%"J�{�UlO�U4��bw�v!�1�����#y��LS���K%V�kwA��s���MU�Q:��t(�ދ��v��
�.;+�{�7��/y��F�_��H�y$iL4Э��͆K�>x�m��:���/]Ĵ����\�O\����ý.���o�4d٭�[��R�m��ٿE�4�t�zd�<뽷�R�,��dJ����*	�A��ʏj_���tl���}2:��JR�g o8hnw���r.���p��]��]�ӆ������޹ ��������dt�U��Cv��'W1Zp������=Y�P���*�Z�"mUpU�^U����B�k�/|F���1[`��ء��r�&����R.�S�&R�F��ﺴ�-*7���YNm��|��C�(��E�F��������1�9W�,��~�(ʃ��~�9V�D%լc<�b��q�����Ǚ�P�+ٯ.d�a���ƑO6JڹA��b�K�[Qy}�,���;\�jS{\�ŬJ#�d�/�-}�&�
���U[w=�_�֖BYj���մ��خ�Z�k6]%/U��U�jo1��N�ߩY�3Lh:��oo0��׆�Y�©�G���U�$�¨�V�l��xO2���;�mA�`��v"�!� ��n�V���,��lO.��cy\��씣� {���(�7�������^<�P8h4�;�S��<B�9�M������P����*�/��Y�����"�ϵ_��,��xaO�\Vq5<�Ϧv���q=�ݟ�wB�A�1��/F��Fe4�F0�<�N�[��xl�����V��<4����^���͹9l�ۑ����MNWK�����S�y�TvM��/�T��QK��U2��V�/�(�u���Ș���X�� tX͉0w2eێ��;~4�~3֣�忹}�<��b+�9�L����vۡw��5(�e�`����Ų�|��C��<�����T�!�8t\����)ޢ{!����>ˏ1�=eA�e��Wa������NC^�A8����3��t;6-j
�;A3A[��Xu�� *��1�f��Nz2n7�ꊓ��0��Pn���Q��Y=�u����M{v�mJ�㽇
�QSsS@�l�y���{r�>a����6�s��wKE��{w�k��{*�9��^���r6���4���}������TU�G�{F�%��|b�H񈙦3R[�nv�5�[x�]�����iD�C�5CMg<bT�Ԧp��7�hZ�kw^�ף�i�����N�ԖN�Ꮩg���KkGQu/�u+:iMp擱��cad�ѣ�qΦ{+�)�k�L�j��M���A�ˮ�T2{S��F䕭���/a�e��)>W�ٸ�����#Q<4&�8���Lk���1�^������ʻ��=�T�W7��l�!�Ѭ����PaO����-�!£��Q�9,�C�YPW�m�xk�%u��(�f�ݏm��m�r4��k�����9A�R�:p�� q��vz��亩5�>�':��H��,��x.���3ެ�@�\=���i�T���.I���n�:z*}��|D)Л2�A��0���k�|%�/?l9�[IpS�ouWz�zW@���S���X\�䫓Jk**\�M5h��.9�u�+���z��q^9&�4�/ёZ��R�;��VVՔ=!��ct2�e�WX�.���g"O���?z���x�s:!�0/-gw'1Cg��]��K^��<|.���f�"��[e�zXw��zcС���P�+�wՇ�잨�=��Gc�ߖ���}��Y���|�I�I�oz�����}��������}�#�~��<>�hs��@S�zu`BgJ�c�����ߒB�)��{��7s�������XT�5��w��ʤI��Y�N���,r��r����z"]ٴ�v� ����H�Z��8�}}O5�*�EtD��%9�Y�]�m�e	k�oq�����o�l��wGD��D���E�K��yW�Q��n[5�'.����1�b�ɉ�z�182{BS��oc�[1T��)�w�lB|��A�G�p��fq���:�od�L^���u�쨥G<}귛�������pX��㎾$��u�숥�#�.�(�G@��yb&����c&�wձ�.�K/ G@n���*,���)�[Ku�������S��9C
���kdvQ�yͬ3N=j-p��gƲ�bP���P�(xWd�I�_c�p���U��sӸ�}+U}�N�9֎/�*����kݛ�V�s���ke�oA��2��FЏ@�F����7��c��x3&�
�jW���^�dL�%�k=��
��>�s�`1��e؝w�B���Jӭ�kA9��?H�����ܫTΓW�0��Igs�Ij�x�nG����#��c�	�r��}�y��m�Q�^��2�	����1����l˂�Э��5n&y�n�	�OwE>biE�>]���z3}1�D����D*پ�B�0h��1�H^ᒺ%����+�����g��Rv�`�'�e�WW�0���F��M�h\��2X�3`U����,R#3�cՈ�k�r��bG����m��bZX�:o�q�-�zIa��ը�J��F�;nr�]�.�O�b:��+aW��x�d4E����YZb
�cѾ|)C�w3�=�=:m�����ei�ԫ¹x�U�
=�������
��Hj@�c�$����S�G�=0R1�}]ӬNG��;q�Ȏ�;b )U�v���+^z�N&֌n�G_��ߌ�0��'���7
��]�s�I��U�Є>r�[:��!D�ռ�O�{#�};Օ`��3F�8����9��y9���W�=*7Z?+��Y&)��vױv��F�k!�`i��r{+��~���c|�weR�[E\���|����ё�/=���֋+���8Ϥ�+`EV���c�%��`�S�f~�Nk��Om_���,�������̈e48�N{o�;��8�^�U��N_Y�����q4�����������ݡI�����Wٲ�(�3fiC��0�+��C�zb>��~���/O��it����[�P� 
�m<�Q�a^l�����Q9۔��H�=a��wI�����lN�p=Q��5��#�9�q�U6��j�����Wrui�.[9��ƳK�#t9�(��vQS���`���2�����N!'��(hԻ�٦�`�G���%
y�[���ޕ؇:�E6�uu��:��a�n�E\�c��ۋ���8��`��9Y�JEWe��,�\�f�q%�hO�f��˨9�W�=��
A|ø��ڃ{6맫�!%/�nq#I�o����]3�v1M��S�]��7��]mrft2F��R�Ve�tǴCF���+N�؜����z":����FT�>��0��б+�w��yӝ�x<<2p��҄{�8�������������MlWCb���mE��k����D��~��=���D�jj�y6Q}?B<��Kܴ��v��C�I;�Q����n2�n�x�z59ݭ�N���Ǧ�/E�+v%'�y�5z��� ��=�J�n�����i��jk��ޏZ�:�O�^qټX��97���P��C+'+�[�˥���M��\_����z�a��~�Uz��\�z�eY�V#h8�7�3�u1:���|/7�����x�<\�i3�(%���c��TmNX�F������H��9���ank�MYmS��<����[�Y��a�����yW��X�DWފ��n:���NY�y���>��5-.�ʙ���GK��\S]��F�D�^*�Y
��s������/r��GO<d��ƾڤ�fش5qݴ��aӍ��]d%1�|u".S�Z�c����tT)�g:�`,�����f��@Na���w:�vL���N;���^��
�j�΂�^��r\�O�]z�b��A^�{�t�`��sjnk�0}`�T�Q���bG#��ە�aѕ�u�Ǧ�����و�m^�#�{��}^�1{K�e�����I3��9���.;P��o�@h�F,~��u��{Kt�}Yٷ��v2�d�Ch�Jq�ɘ/�׬��	��z�o���=��������kgwP�F�FB�(˾�=���_Ƅ�^�j{s�k�'?*5�eTC��!�ю��z��[�GY�� �_gW����x�==�m\�����ɇɐ�T�R�}e�G��R�s^������'K���P翗�C�3N���S+Nv�7~!U>Ch�{:�͢	�z�j.��x��ӈ�+G��J��s�g�j��Pmz�i�^����O��=< ��t'U&�7p�Yt������.����7)�sq�=;=팢�}��`\/+)ukt��zq�ulj��{��(Y.@j}�r��a`w�(x�KWH�g��P/�.�3A�ս�0t�cPt���.׈�#2^W�*l�6r�wd(�Ё!m��eT�6+h�-<�ڜ�7��h���:��71i�[S���<�p�
���6TwC4�G�,[ÅY��fN�����%������bE���hpѾE�~1s+�<�����@˾U8о-�W�{� �m��[�6�����Nޏh��e<�\ND) �`[C�n�sI�|6�:E7�\�i
@S�E^���tp���;m�������'�Pr����w�d���S�#���*�q�����J�]p�2�%Ki�9[x�E+o%�μ�LE�;-��3�}�푕v<:��N՜�����\6z�*©n��*U�u,r)�[�1�[��tPG`����ki3u���'-f�Z8������:.���<��K�\��VCkDe_L���U���1������$��wZ�V61��j���q-w�O��{� �6B��R��UnVOc;$4�����fEB���)�q��ٽ��g�Τews���gu(�ϥ�㉊k�:9�3P��n�akK��^�h<T��;P��M#�n$vf�m��R�&�"�P���ud�o_TUxM�W���S���]�':n�_;N9��n�1����q�%�+�� u�{v����S����2�	���&���n���`��2᜶�O`ܡ�ġe�[�'�4�1sէ[�E�|�n��a�Ǫ'�����%�f��.�S��,�����Z)� +�fv\��Z�6HܳBɨ�c3K��v��:h�+�F���#H����X��#4�ֹ�{eO�h�-Wr̡o���֓��\F;��}�M�ܷܵ㟡A_'j�l���j�ۼ�N����VY�Rk/9g&�S�C�DQ���M������������7�z�F¨]�M8�tV�W^k�X�ɛ,�v��A�(M򂡭�J7��nJR��X�j�]+X�x�^bw�J-�b�NJ=���\�k��m{a���yX�(s%`U�T-��-<Z����{+4Ԥ����F�X
3�W�j�Yf�����N�٤��Aj_@D,���`E��,��r៝
G5���F���5Vy�fNSRR�#���b��;2��jB�/7��t���{�w��R��V���s���w.��!��f�l�S��[Y���+*��=:�tج���k7.��5f��pb��V��5����{(��d݂�N-VxVL}�u�BS�G�X�iX<9Y��9��e�*�7\����ښqҔ �|�̬{n�#b���|���C�GR�U�^���S0�v7"s9���n�<K�o[�8(�aZ�w�G�-��a]��ZjA}���gI����w�j�,ḟt�/���Ĭ�9F�a="�EM<�b�jQRY��O�Y�����o)ϱI9�h+���[}u+^�[]n^��f�BU�=��Ln6�wR�e�*�[�{��3��Zq�}��B�{�ڇ�nG��:�M��m��>P���V���j�5K����0�#ru"@>���p���<y��!���Ժ;��;�$��/�3�+�W��������Ϭa�:>R�f�t��1�_�o��t�����z����lE\g@���f�;����\^K,#�p�[��9�m�o���_G��i�^,��6^��fS���쬨��xtk}"H�>��"f��L2:��QgH�ӗqH��t�:p�WX�8��r��{�#���.en?��|�yQU��BL�<=�},�?-}���3[���uI�5��x�A���[��S�$�3��@��[����ݬ�|Э�������[�Т��[�d��컐�}�7�xW3���M�?'b��ެ���G��T53�(�_gN<���+��d%pȬ"�x6&�z	�[9
<�U�5����2k�E���c���Q��J6T�J#�EFNTT������ہ)�c���Dj̢[t�^䩅�j�_W��7q���<�eS�V�2/����q�e��\9���	'LE�3Y�R�4�_U�{��8�;��0u�!�CX�e>$=M���G�Eks���$F��4*|��9�&u��b��t�\�h������I��R�x��5�����[}1,�f�U5$��8�gc�N��W[����i�9fXJ����q=�A��m�,ۨ{DhY���k6�������zW��#wu)t�Wj|T_H�F���������ưi˰}��JK�{������L{I��]��J~�ٖde�VR�t{��ssղ�KA���M,�պL�z��>~�V��ޥE�+�l��;1\x�����cUi�}>���ݫq�ٺ�N�6�~�\3�34��q���{ޚ�������f���N�}�Cw-\�+�����]����v�����B��d��\���,���uWU��鹷�{�Jֹ�Z~o�d(���s�^�ۉ�1&�nx(����
n5�4��i�Cgi����t�����-��bQ^�iy�t<'�T�^K�!㣙~�nM��%կ@]�0���룔J�^M:>��
>�i�=��~{iձ�<C��U��U�h �zv��^Ź�W<{���/�羸�Ws��Oƈ��9+m���h���Y{��U���Ȉ���`n�n&2"��R����L���oѷ�>���еD�xHz�#�j{�\,i��������2���>���쐧է��[�����<��i}:���J�V���GG�Ѧd��p�F,�8���Ci5���
/��
K�sc�^@Ǳq��S����#Dwj��v�#���ܽk�v"�f�{ݖ2��A�]�WR��k8�{3�FΪY7�t�1�AV`P5�͌�y\6��i�r�v
�Ϻe2��9W�	U��FzlZ��ݑ��
v��8�DGCָ,|��|E%唢��x���I~ԟ�ۮ(tN�Yr&E筗�%nZ TS��xҨ<0����DlT����q�}xs[Q�K)�.F���q�S\+iR��C��f�9����=R���K���#�^6��nO��,A��$�Zj���#�;	��Q���0^����GR�Pxi�i��(C�Q�gE�p�����^;���7�$,I�oK[�&�9�u�o�>γ67�#����D�ɋ�� ���8�
ޅ�lJ�0+Ks�BO9��ӕ`����h����^tCxX.�
���nc�}����"HR�Uy{i2u�B����%*�>-���Eu�y�����,��O���׫���}n���6��//�ڋ�!U�͜�5�}����S8m���̠�����ޱ�]A���#���\��o�^�a�(�_e���KR1n�`�Ίycm�6��&��[��J��y�+QK���ƉT�F��Ҫ!|�U�� �	_5W��SF�ث�t���ٓ�{��Q�ݮ�O�5�����l��}v�#p���t^��oLǩ;x�D��n1�d���n�.-P�����m�?����D���v�,���,p�~�0���2G�M4z��^%�V�x���ݚ�!\����kn���(o����IG��73���R���^V�j&�k�y�mNL��fV>]�u����<��*7��f)�*���Ѹ�y���H�:{zo�.-��d%��੾ۧ��w�]b?<�'�"E�ȑ~�z��>ͣK*q���s�0-�����(ר�V<^��6n~���_���8�wˍ{���9Գ���w5�J����b-��5n4��B<���P>�a�~�\������2J9��G-R�P�1�'��8"�U������Ms�{9hkA���7k�����FrW�'##�T��2��usRw���tO8�'':m��71��2<b;`m��[���>��a�|�n�B�5�r��3�ǧr�4�"u.�O5H���"�ܭ��@��~��.�7<���6_kc��J�jpQi�vٟ_!f��Zh�n����z1G��z�����%����x�u�_��̿��
ԣ��/�k2dAB�]Y�Tz'յϴ���z;s�b��Ǭ�xA�6	ƍI�����9i3�����r;]��Xx^�
*a�Y�;
�WK�{�U,�]�L�c��+��Ps*��뭑@;֔;����{U����~��J��W�F�մ����̀M�rC�صpF-� ���2�e�̩�G�ʌ�U�y��x�����^N�4����~f�˲#te��Y<̽Y�����8�P+ޡru
��;�ȾX7^��z�aŉ�l� "��L���].�9�̉#Y��]>�F�AbVNI�7���w�dUu�-�9��lnǗz�+N�Dv���N-��!_�k0��ief�fUGt
�K���R��tÕ�iU�����|�n�]ׇ�כ	��^aN��}3>^8�ve<�X�ޝ��+inTW��DU�
�yrI������*5G�U��Y�y13s(�AQ˪�(���[�y�֪S�ݢ�f�L��|)�eR����{L;f�c�S�U�ם�B:��H�f^�Mܢ��(s��Nz�3[��c9�32rx���:9q�u�m�N�>��;�9E�b2�Up�d���ן�k�1�����F˨]���aQZ�n����]�˘�v)Ё؈4�����V���Wp�Z���fsoo�MG)ߡV�.�j� 2��6�e�7����ʑ�j��9��qΦ��f��Q�0m�'G"]b���j�e�i]v��d�U��nv�u�ڹ��^��x6x��ױ�6M����M��|�tt@�WcT�FKnIc��l�/7%mX��Q��)�x'k�{f9Rف��mD+�w���AfP�H��t�R���aJ���%y���wz����a�@8+E� �+=q'����ڮ�g���D&���&�|�URa���3n)�)����PV���|A\:�O�@��E�y���� :��>���u.y�s{��mw_HӍWױ���Op$��~��bu�.yWr�3S�+�8H�<��٨�� ��jW=cǮ:8ٳGϢg�D����odL�.��k�Ĩ�93�,ÎY��L��Ϯ�-�����0��=�D��ӡ���tr,�;DF�Mb:�SFc��n��7�.�rz
�W��+']�\V{Б��K�TÒ����k;2}�r��ǢB@�S$5H_{A���)6i��������J��h���T&cxs�w�2�I��f�L��˃<�����8������F�/8h�/gYg(�z���r�cqQӞD�>�ٯ��*h��y��T��Ǐ�R��{���|��n�k3�qv�9�2�\V<,�7y�+i7a�Cw����u��<�4���Ƿ�۶F
	��2_%��arȘg^�wNF,�pu,���J��X�Ϣ�l"��U�_:ml�2��%c�ҼW���7�/(gr\r(��ةԓ����@��=�ng��gq���~\6����u�R荎A���W��'��(��'�ױ������:�����^"��L���N���J�[	����[ʜD-��q�5D+oЇh��1<�̾�b�6zҘ�z3v��_P�/?�x��f�{�fjŤ���mC����i1��ϲ�`H�!�)��U+`.[��&{�����"�]�]w�FT �pf���ىo�L\���FF������IG��0֣���%��i����f[kё�T���}:{�O�5���}H�:��q0� ��=�z�~�ޮ��#E���E9�gZo�tq�9���D�jWs��r�����U����L������{'�k���{��JΊ���Q����d[��
��	��;P�>az��q�h��;w��
ꯝ��xܬ:���t	��!�c+njW�Uc��e*}�lp�Ga����m2��n��Į�=\*-
�7�Q�tV��9(9C�i�^�{�<��ix"奄��8����g(8A��bэ<���������{k�σ����A_P�T��!ؒ�*��B�sQ������8f�&̠{oUD����WN�.1�(�P��D��B9�$��[�$�S�*��B�[7f��u���Sp��<�É���q�|@���̛(��V(�>l��{�f9��g�^��u�k�b��LmD�w\ҟ^IPj+��B��n�V��~cv�^������e�1�<���[����>;Oخ�v{fԗ�[p��6s]��u|+��;�&-ޑ��$�w�+�Q�nR���v�Q
zi�a�zLd��[�_��W".pB.���W{�f.�О>�{���x�A
��3+.Џ��yH�!�a��@}�#���f�j�b7jT}԰pCY�Y9CS��u�!/iGlk{W�WFz�K��-�|W�������g����ۓ���j��w��;[wV��B��lչ�FP�����<����@��L�1���koʷa���t�~#��{�'��Otnz�73�e�;Xм�3x��/ߒ����1�>���s<���z�AѪ�C7���5�ӣF�g��������4����*\s΋T5_
�)"v��-��Rnx�d�z��"�O�#u�9����ݤ��>��y�l~����d�_W7v#&v��.^�g���]����k5N�3��'{�èu��+g�����Y��T�H�m�vw:��[��u�m5:v�pG�gqeͺ�X��*���y��z�G|�:��B*�[#����J�ڗQ���٨t�=�6M�� 9���
�[:J;�L�,��Ѝ�2m�#�-���\;���=�1��������]R�rY���n��1�'��O�Dk��8g��o�?��X=B��da�_{�9�ǫT�^�j�$DnD�{j��rL]P�*������F"�6�T�zO�`bٷ�{���&ת/:V���`�a��S%�u�O�戁����W��2\>���8�a�qE��ƺ�U��[����w!��(P�P���t8­x}�Enn>Ay��|iv1	���{���)���S�wŽ�Bu�>XB��Ш.t3f\��p+킫q>��f=J����˺�.+ʄ�,k��� r����Mu��^���_3��AO`�Ԅ��ye7�j
�x`�sUZ��8�� �
�A �Qz��=�+`Gd��̗�z�s�V��ve��(�=Ef��%��u
�W��$�]��fz��:Gk/G�\py�;���NxQ���">(�E@�����^���{-TηQ�7kQ�Ĕ��5j�A�9���"��3xֿE�HF�R����&L�1�u�ࣛfŮ/�=�f�J����ӅE���tYV}L]w�b��t��1P��TR@�^4�u���"���`��oX�;�M�b|6�w:���e��s�FZ�����un��l<�IR�-��h��w���B�g	�A{��G�q	�շ쵯s�]A
�9�,<{8�m#���30�sj@]�j����t���N�}�O��j�KG�شS}�8?ƌ_��)}�WC?v{t) �Y������!�X��hv	�y�6���Y�w��=/���|�fD��v�<7�)��[-P1�zz��u���I�*�����2 �5�G={�)�Tk<r9VW#��^���o���rV�)�.�P��
�+�i�\�k۞�P��բ��:s���w��9y&-��n==R7$�5�6r��S����OWt}0<�b
z	��x{W�]+�8A�3�^{�<��]��x@h��=##b��2����:��rO�2��}�h{ߝ]ɔ�ۅ~T�ݎ0 ��S�x@�u9ކz����-���v�Lą٠�Q ���$o�Y�U����*kЍص�^�ஒ�Tt�{=m@�]E?�(���H]�L-��n�����j�ue���y*�.
�Y�z�����{�r=�\����Iw��f'Ѱyҿ��T@WN�j3�u����W��G�[�Qx�>[�Ot��ױ9��n�o{ �v��~8��u���l��w���iͮ5�.3�]o1�ܤ��x�mw`:��]�%��ri�/ ���7��mp��/3���k�'�'���ϙ�/%(/�Y���e:�lu�F���hI��򐭕��0���N�7]���(��e�^nPW�^n�����]9�s2�SXw��=Y���>��8��s1,�N���+nN7�F�Ecۀ��4,ɪ�
M�GkI�u§�1��'&�c4��MAV��,Z1�t��|7�M�mZ�o�'7�5�����][3��ڀ����hGk�'�X�X���r��P�J��W��L��I�إm��eݝ���'�z�{ۗ��JX� �-\f7^�ve#7�UVr���F�
e���P�v��ޮ7�֜du�l7�Uu���z�,�x���U��{ҚamMhv�R�����QK2��8$��t�ف�?�.��C�&뤀�Gq����ͨ�q5L)td]ԧ\+4��cݧd뛹&,M�N:a'PȴfC�*E��W鲡�7�p����`�90b�r��n����h�)�������x�=!�q��[���5��A�y����pq�tRu�\u� I�`�Y��|�(EwG�n��Vį }ס^��i_zn���a���͖�0U��]��U_;��ʔd�ғ��-#�q��"έ��ճ�bn��� ���-�����*دzl���E�+C�<fڎ�S]�ع�0m����4�������
��\�m!�*�]7wsJB�_Q�$�S#bv�˄������O/���4$��G�\�gtUޜ�er��ă�m��l��"�Aړ��i闃���Nҷ݄���>���*H��^2.��b�.�0��0��C�1ם[,&�MN�k��bEe�Yֳ�J�x�HO��JWj�L]o=G_�f���+��#�B���/)g��̦ތקv��w�b��Gg.e�&�ʵ�'3;_r*�ض�8�*����7����SN�y�쇹��R͖�I���O��b�r����N�Vd�{��cS��=)MyM��d^����t��v@%`ŷx���Np7Su�`$D5*8e�L��v7��JW�����9�+�1�fu��U�����=X�w�սƳ�V�m.�6]�ͬէqgD�`�.�7���tc;��Wk8.�@f]��grl�����Y�V7��vH�oo3�J4���"���Z��U��}˂}���N�l,4j.�!���2����Sd�e�u��d�w/��`,̀u*tt�O�����:��[Xc���Ʉk1�$t��f�"�H���n�i�k���|��5c��é`:�K�Lː�$�&A-����ّ�me�ǔ(���-X��l�7�'~.�@�v��>y�h�|�l��"Y�Y�S����1�����v� fK�]����;R����V�'��_�W��z>~":e"F���2N��αL�GSiu:�n�}��{GNu�v�Ugmc�`���t��KY��ؕ�F�g3�����4�-�e�9��J��/ � )N<��na>��7��y���|�?^+NP�Au��;��v���e?$G���_�r�w��Ȏ�Ŧo��nT��p*2לj�iϯب}eE��>u�P��p�o��<��l1�ُ5��-��;Y���Cy>oP�砸x_���u��#*��p��<�S�x!>ua��#$CT'�}�f(�k/��xCwPc�KhWwp��g7��>���is^f�%[�ër}~�f�����IIbVh�v���0��n��RG�1������%��a��ޝ��$B+�)��F�Vb�)�׬��뉬���~ɯ�&ʹ��gz��Y`iច���U��1	0Z�s=��FggѮ��T׫���9��3L�x�hmz�hpr��wO��DUNΏ8�tb�u�&j{��E,|!c�e��8l�<�|=��v�f5����$8Zݪ��|c0�	d'b���y���h��O ���Ćc��n@���R�q�w��1�w<r�C�{�׈�;�>���V�L�gBO���>ۙekr�Wg��کc7�3�G=���Q�w�8���)Z}�{�f ��M.�tˮH\H6���d��V
�˵�\�
UZ.�	� ���Ɔ�5��P�_��;��j~ԕ9n���{c����xd7��9d!�p��]��Y��@�02[�ꑽ�oo�y~1�f�xR��/�)�����R���F������p�W$����5��M���U�>ބ��TjTp���[u�R�ݛ�P�er�@��5�?Jtþ%����i�WN�~�6�DS���UOpi/��f,�0��k���7�^e�H��WiW�6�!��������z][����`zK��M݄`vBq3���V!r������P�6�rY�ץ÷�{(R�}��f�8��K�z�������g�J�N�+w�p\9q'��ܥIU����݀Z��N;8�^�b���r��F���<4�a�,�qsY�w���c*�E��� �P��G8��y�Py��Ҏ�c�M��۽""ܷ����ay�z#j�:I�g��Υ���H���C�W�G��El�g%z� n.�9�O�$����xx�f2/����#�E�X���~2���V9�!�0�����#{l+6�*v�S�U�:"�8��}�m�VlTcǁ���)6\���Vg{�R~��ӻ����u���uu�yT�ɭHӛK�v,^�xŕ�Δ�WM2u�[�w�{Jӝ*���9�I�#��I�Ok+�ɸf�-�!����Am��,kB��~$�^d�66[���IH�4x�邶��������C�Ǔ�ܰuǯFw����ֲ����[�ʾ7�4�l���eJ��G���{�bo��S>����j�T��5�>X��o��c��K�#�n�1�^��?O
GY7u��1˄�]�p�tSbr4�=�
��/�%��׌�Dz��OE�u�q|�"�!��FÈž����\�DތaH�hlxf����W�+�|My⌝͊G@Jz5��L�E[�Cg5m+��jn�ε[e�@	����ձ���[��:��T#P���A:o� ꎓ�U]Z����Z����=�^�=�^�^�6�q���j���>��tPS`)}�[��W?����
7lB''k'<>���[s^"�b�W7W�.\z��t�㠕N.���f�۵�A�a����<�ԡ̧���Vl�7#���QV��2��4�K��Zġ�}o�)U:�QP�n��wo���_y]\uDw��v_�Ӿ�1O�ɵ�$|�!����tB�?du]xP�p8��W��x��m��ԽBbF�Z+�VJZv��;�@�X}j��22vǻr�R��XL�,�Qs�$��PZ]���nw]1��[����e�\������₍4mTVi��vʃr�e����pyH�OH*�K��s�>��MdΣ������p�����@��ֈw}��@��a�.�ޓ�����Ξ��#a�����u���Cخ�MI�
i	�Dǵ)!��gU]�@�nFEuāO�r[��\�9ծ�W+���`ٽB�z��ET1<)���܈�0AY��z�|v璻}�>��A��w�lF��[�p��]�1d1ë�a�)�8��;�Qt���غ���K�QEޗ�9�֗Op��ʽ���+.O���'g�
�R�0�������?���u�v�������J��]�^�|;����i=�zd��}j�d���F�:'�Bvׂ����6�ߟ��\y����]�������3��T�G�p�c�J�#�l#��@H��
���a����ɜ�ܙ]c�(�f8垐�n+Ƿ?D�:gL�p2��H���0���!{C�oQq�9�����8ܽjz'u�XFgN��Z�B�8�L!s��9�$�{����b�ge��|cˍ
6Ƙn�]鮼V�|T�#�z eԾc�r�lg��*W��7	s�}jh���r��D����9����8��jiS��xw:�F��2�Z�q�`�yچ�mbl�����|R�B�,; �YH����հy�E`�ԗrT�׼�D��Dגt�8^Q��,�WrbD  x���H�M����w7Cz���o�c��S+�M
�����sO'h�7�ⲏ:8�E8�r�A��T699�(p�<�ʹ��h|�ӂrO:�&N�,3�8yf����@�۟b�ΫǮ/��f���-�	�ty�7��z��K����;UV�1t\Q����u骮�_��%q��M ĭ�驔�O���G<�x@-Q ����5�b�ώc��L�]��<�'G�+;VV�5B��f�� ��oA���>D��������	[x_5Ahm]dtw*/�vO�����#	��t��G��']�O����\:��9����W�;�:����z
�/څ�=/tF�-0�)L�6�7>��*�����@�z��dw�CA�����^�{�7�^��G-��7j�B�u폯V���<�,��}�Zu����h_R��6>̞[]�{r'�o|����ν�������,��o(����q�1[T���3#]�`U)������r��*q�]�R�C�c�����x��S�aM.����F�q������fN�CSH�H$;�Ktu���8���Mɏub]|��Dݠ�!L�%%[��^6_	�{��ZH9�G�M��2�:�P�z��[�����u�K�6����Ԑ�q��Ν7M9����w�-GoA��~�ӹ�v�z�gEN:wu7��*�#�}��g�i�3���x�R�z��Ó�
�yW"<E�W��GA����d{ϻ>�dzn�I�]3=�o06��)��\�O.��w�c^���U5�0�<^�0�s̺��e��7�U�X-�P�&{�m��l��+������P�&��3l��:��(g��a�:�F��}�z�x�d�+�-�)d}��B��i+�C*+e�f!�i
˨�U���T�0��]�R)�;�+�g��q*#:\g��;T5�3��g�s�ř��׾����IZ�w�߶�ݏ�[�&̷3�W&�����M�C��w��/�ȁ˟Tp#)��Z�oˤ��u���5+.X��}�?��''��Q{����5`N������S�NsJ�Ef��U���|�>u<ӕT)Ń$F����]�׎��.��t1ә.z0�Ǯ\_T��K�S����c��&ЫWIF�d��6Bq �Ʒ��~�oM|��~ 1�4���[����4 ���j�R��0M(Q�OB���;Q�M��
��L�X��Q�K`Z;�hW�q�x�e��o2qH��wX1Έ��|��g�a��:�M�g�pFY��Q��&h��f�8$�X#$`O=��
i�ޞ
o���2�Զf릚1���=>[�(Dҧn�K1�{���;��He��a�0N������ܽ<*�o���Ͷ��pp���Gg���;F���s-�X�c!R���!��՗��p��q5��:t�72tp��'�Ot�W=������O"*��Tg�����F4�sB4���9�q*��u�>�خ�����	����a�w�&{J��,��@�)�����v? n����\ͨa|йW����v'�4�ϻ�IjVV���VZ{]g��<}��͌2)?'W�"5qUnΥ^�\��v�1������̐�{��@�li�}k���k�a-f�B7�h_1BRgh\ǎ���V�6=�%�Um����T�0Y��6ج�p�p�U�>޷3������j�rr�������Yb[�Ѫ�s�H���B�m܈4��P&3}K�끅1�1�䡇�或��>��a­'�ɘ1~����>O��S����s^����E�_�k�lc4�����'TK�B������MdE)ҽ�&���v���vx�8tj������;�h�aU�K@f1{![�-[�Tչ����L�G^���Y����e�J����q��߇1:	�x�t�Hwi�5�5[Q��Շۇ�%�Wo�3p���.�3��k��U��b~�)�D��Î��w�V�R�w�M�Ɂfr�',eU�;;��=1�sU���z<
��^��(��l�t�]aw��2������}kDέo�{y�g ���8��צ<�K���E�z��3��/�T�om3q2 ��!��r���âGU��:/5�Nj!���,�~1w=U����{"a�����$��.�y#���k�;(�+�ZN��[���]�ԅ�큾Z2��D�{oA˶���'{i%�k���5���7=P�<�����6�<#���^d]��o�m��7�\�R��+�g�d��s�^>�+6�`R��y铧�Lq�[��p��@�E�ݽ+��o�S�z.�(a:jy�,��'�'o�B�\&fj<!O]'t�]w��١��An$	��}C�{�I��|
����dv)ե,��᷀��g��^�������^�3^������¿jۖ.�=�7?
�`�����u���g��kѮ��
���[A��=ʗ�_�X/] 	�DPv�/%m���7�A�h���b�W�*��38Ճ�P8E4��*S�P���A������wOȋZz t���\�e�te.��C`����@�K9e)אi�@�kR��/gbL�{t�uT��iv��Z�����˅}p�w19/v�$NZ["|���Q��;�%�}p�MV�
c��<8G=F�u�"��P
�C1���Y����&Eb����{kl؊cx;7k�a�..����!�ؽJ�xp*O��{oF�NW����%D�{]�+�Ik���ǃ���}w�9�,�Z��23L�N��#�5@�n�`.�>�nS�6�O*�\�1js�w�`C��!��bk|�["ÿ#W�C̲��-���فo^�--�s>B���6����=�g����9��I-�"���ulk������B�̔�O1��G��N�G��4����yw�`P�b
���+P:���y^�=��9��C���	�'��ƪ���K���wl��S����x7���o��L����ܰ�9s�U���6d}�觾Z�����h�=ޛQU�5��=/;b/
��=��F�=S_\k�*�\ϱ�h7��`ԥݰ�{q,F�G.Ւ2�����X��������M���gE�u�"3<W�E#�Cº.��ґ�ڪ�-wXz�#9�mz�gŹ�A���;�:�AHt�'Gèk�5������s+�A��h��e�oN��P��a�Z&З�%�mrƹ���~Y�M,�4���}��C��D���[.j�V���&5a�Ρ��=w׷{v"��u��!��F�������4>��M6�;jf��;՞%V�罹yM	��Q��kf��pt�puT��$���z�,?(���:a3�9���sh�k���{�P�oz0���X�!��p�IW��:�u�<�<�~��g�NH�D�����b/�;벴�t���]H(�B=át(����Lu7������]�P�Y?��|��W�
�>~���J�Ӵ�(]��⮀���޻~��M��+��z׎��{9Ȇ�^݊�kOLA�)fk�q�}�X=����e,꺭�D��u�ͣ�-��k�!���V�yPv���}���*����K�C������}]&]��v<�;�Tn19�յ�����������e�h]5$��״N{�C����m �! 2����=�� ?��A�F�Q�݄+���o��=������J��_Է�}zl{lc	t�W�Ͳ�>m���2��ۺ(�33��{ıʦt�Y�'F�y
y4e��ײ���ݣ4RҳBG�A0˩�lV��l5����$�k��'ܪ~[�:���r��ќ�["a�Μ�2v3�"�up<gs4y��lqs��*=8!���x9j������k�D녶�M�ק����:.C!=�'<7��ớ��w�j�u/e��nhS��#7H��Z��7�oI�9�M�����T�JNV�Gt���6()h�v��i����������{v�$����s��uU!qt����:7B����e^l(��f.X����_�Lþ�r�=��;�y���$�I?�H��_�@�?���@	��I$�hd!BI �6H��$	$$_�! BC���������� �$��I! M��H����������� {� {ޟ�?��~���X�G�����*�����׿�劐X1٠���=e��Vy+@�n2�Xj� ��7���}E[L5��&�Tr���{�
�3mKb�F��RH,H`�d-�t]`�W�+&�Q&��`��v_�ES˽Yw��v��i�ް!Tu&wv��`��b2�K:�T��D���S�N6�{7K��nS���JPw-��R.�AK(�r�խˣb�R�d���f_����-�d�e������.?6m������S�L����4k�Ӕ�]]�2�Z֒�M\�m�1�0�sb�e�aܦuõ�����Bd���[x��N���{a;���(�5+FI#aI�"�������VHY��=��ؼ��;/@���@恱���E����Z����8�@gi���Ӌe��#(Ë��a�&�, ��1;�K��f�mj�Y��jx�&�Fj���D��$�s2��X�(���Wcq��^^^�X5�1����P�s%P��SF�����ѐIM���o�c 
9cN^K���7F֋�d+�9N�Q� �B�T����qR`+����0딩
�D^^5w�tL2j4Ui�[r�J��U)I�e�t}*L��cDٻr�֭l8.��V�V Q�X��:�6�P$�6�3[!8��-9-cR`L�m(�㙐�V�����4��$�̷��lz�8m�y�]�O%�6��PI���n�ڠ�l�	��H�q�b�D*h"i�n���r��ku���gLcr[ �����^]\���a3��eDD�1�J��i!-h��Y�l�ʸ�қj26�,�+��PW.6&��b�4���jo,"ڔ��[	!��.]�^���U�
F�+@:+\FȻ���� �le�.v�ɢ�"TY�,0X�{�1����u�H��"����
Y�E6nR����Uܶ�d���Yi�Z�k��g�5V��h�=3��4��η�4�ɕZmOf'[��Ec݋R3]РS�i*�r�r9
1�nF�q�*6iaDS��m�:q�@�V��IU��bg�E8�U`�J�l�����`&�8P̶ɴ����i7n���J՝R��2�4�HE�U�%J�j��-C
*��FX˳n�Aur��,+Y�Lz��FYѰL�-J�Ya]�	6��l��m�V,�tt��Rj�M̴�%r]�ͤӛ#ƩǠ^7@���mݩj���87MA<��e24e�)e����ZI���� ���;��1�q<��1�b�+Z1^L�X��
��e���bS�FMQVk�P��4,�Y �B��4݊	���25b��V'����0GV7m�����xѱ���z!;Q,F��Q����\w11s!�ۨ�ԈX�8���.���.�٧����N�X��F�IZ�DOe�2@��ȵ�g�P��(�5��r
V���*��3P�d�{�����g6 X˺jM#2�3l(*fKZ㌣kEX�̚M���3z��S�a��.�ټ�Z ӸQi���D�,�����JV��ml�7�tm$��7�n�m��N��h�r�]Ag�u�J݈	7A Y[VXR�͙��t=��"`�M��8�M��w[�V%Kx"���G��7��t�w�Q�qXbT�%]�w��&���
�K	�Βh�j��`V8�I`�甐���Mf�H�2�m[��(�m��'oo�#ݦMSB���!Wl2Tû���hۭ��P���x�+Ӡ��B�T��)&Ⴔ%j���&�HTt��3r�J���j�7E�8�WY��M%%��c �&�m��jR9t-X-�%jÇ��5t��U��6!B���״cKk"KV��Ҩ� ��
e�m�̙>���aͤ��gb�5hvUQ��Z�D��41f�4�0�!6�B��VQU	U���T�Z+1���I��pSwL����%�x3R�s �rH9�fM"U� �Ş��^E��}h��[���2�����?4��5rJ*"�R���@���f�[Nν��/���C)1�Ie7U��Jƅ����fK2��d�f5B�5�X�ܬR�*[�bm��h�6*������C��{��e�%�p��^�ƴ�WVr`�
�dKE�@ݹv�`��PYPfӮ���D��6 �e2j��f��	�eC�f�^���wE�`�Ջt5�mZ�IF��M��
}��쮑�����2��-±�ى 0�T�b��	�E6Qut*�W��A����F�b�Oq���I2*"<x��0P!�VӎU�C0B��s�^j"[JH�j�i�s@өh�F/.��˲�!h
�3R!r��
LMdk�Ҩ�ъ��[m;
-�ڬַ�D�J�m��,��[76<˴�16�E4)�]J֮hJۓV"��U�
�clL�i+�X�B�W=��s!!�[��J�8��2� �9E�F��A�{hM�"Sr�VT���m�"j�Ը����K
Y�ĚȔ��װ,�y��xKR��2�EN��t�RV-�+M7!�g/u�����Pa���%�b�;��wG��z!B@�@ �H�@���HB	�2I%�H ���� 0���@��		$ `HA��@����?�$I�-���S��$I��<��}�`@$����@$�I<$I���H���k @$���0��o��lѠ	 O��	 O�O��}�@@$��$I�������4o�� I �f��������I! O�Z�! No����
�2��de���Z� ���9 ��>�����(���S�U"Xd�-m�� �Xm��V�I�*��C��aUe�AX)JV�wi�  6U(R$U�jF�!i�IH�d�T�)��$�TQA��%"�Ah�P�Q
���%@U
�     	MP�R�*)٪��l�@�һ��D�"黀    � �   � h�0 @P($���\G��T�=���m���/@�^�vڢ��Õt��	Sі��c�7c�vPz������tj�wl�)��om�ol�{l�{�Mh F�;��嶊��k�_c��$*D�T/�P������ge�U6ޚ����Wt�ʣS+{of�v�]6��unáZ����7��ǵzTweS����ײ�u�ݵm]t���S������wr�o*3
�Ψ	�ʔRE!PR����u��:���uŶ��v���mZ��۝j�:7n�{Ǫ�owm�]�s�M֭�U[��Fٮ�Uu\���U{t�rU�����n����緵��۵�T�
Q$����TEJwOml�n���.y�jc�۝u3���ޯz�h��z/y�7{���2Gj�dٮ�ǷK�v��K��׻{W�]]=�s�۶�\�ۻ���^�^wv��:�uvK5[����#�BAH"�$�J�ں���v�j��m���ͣ�v<�.ՙ31�=3�즆n��m�4�vX:�g��:�ZS�'wv���z��n����4��h�D���^��Zc�Y��5#����B�(��S�4�Ժ���.�v���U-�cV�"]\I�w8ڴ㫝���w���x�)��۽*s�s��ne[luK�����u�^뵮����Y
+���}bJ�JIJ���������q�ӂ�uݴ��]�]SMn�b��r�k[��Y����S�U]�i��%��u�T�j��U�[wR��3ge��:�w#8����m�i��D�PE)9T���;��wQ�{�u�Ҭ�ӧA�]ԭ��V�����-�6�1tvJUn�nJ�.�����Q��ݎ�Y�Iݭ�ծsoO:<[u�1�(HT��$E*@$���5+#t��wa�����][�K�)b�����WT-�wu��ZU�U�kk���4�U��imM�s�����Ǝ��[H:v���UOl�*ٔ����z�Y�g\޷���%3�]�w,�`�y���0��w�����s.�(�9.�e����ݶ\ۦv֮�c;��UB��g;�%�$#����T�*�	BQRU*�(��' ��	��T� h S�0���F   ���'��@   O����@@ ��*�6!23F�&	4�$�#jb�1?��~_���+��R���Ra�ئ�˫�s������~���|�����	I�7O���rH$$?�����HK�� ���H�$�$	I��	I�"�����0R���Pm��?�1TȨȡ��o�pX�3\��NӚ��L�:�H�J�Y@J٢`.XB����͡&9�u�IL��Eh@ժn[�M�pfd�bN�i��u���c3^m
�'qL˼Z��nejA�@ŪZ�8sE�I�vicʂ˥v�Au(Ǒ�vi��MKI�(gʱ�?^P5��P}���Xm��?��4�Tv�����TD�m�tL#2�ӌ]1��/܁$U����i�ѧ��
�ژ��9�U���`���0�ŭb�J�E�d�(<���ޣwXi)�� �^��ژ��OS���T�tҦ��k��Ž86�І�����o$�������Й�l���&�9-�n���]�E̅l�Y31Xp�6�E4��kc�Z���m�'�"E��B�͖V�:me͔F��Ĉ����v)/�m�X�42�WQ]� HGhZ�$������|Ej
(V��,�()�$��E`*�5�aX�#���X�Ā�,
,�,��g��k\޻��q�{��{����{�l� b�y+�P�)Z�ƶ*%eE[h)DQ�U-��m�ʻ�Ƞ�-�2@F�kp��S;��vFS�Su��d�2nh�VbA`m���JʐR��E2��T�J�DJ�%C�+&%H,�޵ޚ�x�M���z�y�{ۇY6���y'��4m˄ܯ�=5T���I�Sjشn[͒*w3���ڥ��V/1���-�i������쭔T8�"�b�Ѝ��Ceb��)r�Q�/W�'��{�yku$"���B�gh�
���9��G&,�t���9^�h/��O�K�՟L�&�(};nTx=N�ь��M�JQ���ۻx��Y���Y��)L'C80�����Ķc�n���]�F�MW���ɂ
�[��
�+7u\)�[Lnh��5�zN������* nY6Xenݧ����U=�iվB�x͎�U
�R �.��R���T�����u����E*��WYHR��;B�Jց�u�ʷ3e���$�����BBu�I����8�^V9i�a	�$jcw.�e�R
+���Eja��"�S֍ɧdj逵[3ZP,.6^f&�re���u9M�Ǝ�;����#���x�-��ʔN�řmI���lX�"b�N]`L1��mdUy��8�	F*��
u�'�2-r��aޅV���Լb4ED[�3-��G47CK���fB��!ͬ Ŭ#2�k�i\�l����xB���I�mKm��w	��&��S�I� �fh�$Nf|��q�m�Z�1*�GWKk1RF�� u��&�d1�Ԉ��"2
EcA*�b�1Р����b�FA��V��E��PR)$Y�Vm��*��-���nⅺ��<ɅCDc
�°�"��V�.��/1P��~�}�h�]󾮡��d2N2+����2�6������wLi�S�YOq�V ��ڐJ�s.�$��|
c����X����T�X"�i����$b�)�PQU`�X����`���YFe��X��b�̖ �X�b�2�*��N��\E׳�ߑA`�fwtZ�
��,8+4ϝ�2��{(�=�R՛0��<`+�dV�H���)�MMM���J�	 ���z콧�-{d(�G�%d�	Ps��^��kE;.��i�F�U0#�`mm8�˻uk)!/Pۿ����7��vF-K�ʚ��a���vn�=�u�g{`Z��*��˟j���f*
X���� (��t��J�[�JV���Nj�ٹ%���#^�c[l�yDRP� 
Y�,�Dbj���UZ>�cke^qK� VPbj_B�nآ�K�:�V�I��)n27YC\�Twi5#�Z�Xv��	^by�Iw�(Tӻ� m ��2C{l'7��{�wۼ�,��v�cK9y@<g`9��a��7p$��a���VdVë��Bolm�j�[ػ܍�݅��u1P����w�B,��.]Im¦�Ԝ�2񱘤�uڗ|���WY������I�fQ��F����Y�"(�mS9��V]Æ��(zfkQ�ʵ.l��aK����nJ4�xE�ZU(�:�L������c��UG�Q �e�̙H�N����l��.�d���M��{F�� Kv�+m�3I�*R�rn|2M�F��c-���,SR�%�Drc�)�6�90cy�ÖT$t��U'��z#���(i$1�eBհ���v�h�mlr�Q����n�h5��2C��J�˫%�l����M'b��E*X*�M�J����C �[B���J�5U�թRC�r�:#�E�S�P�c%8�Р�X�4Kӭi6�guw��Ν��GX;�d�I1��X�FH�FE�2#�@����ł#��b�"H���XU@�M����V]YӶ��g^�.�r}�l���1��M��7k.呔��3e��d|��r���f7D(�8��F	�c3+���l����˹"�dXy�`q��Hwe7��Ö�;����y��u�1aM�k�hD�p�N�Fi��%"���dn�6�Ԃ�;��dwK2���R�EF�ԬV���]\�aDqMjĔ�Y�7@��5̩f��`���{��h;& Ԩ����<�}�Hm�I6�l�>�����lS�W����&m=�ݢ�*�&�F�1�,VӼ�k̒�?��4]�Lՙ[��܍F����w�ۅB�1RM��4�0�����{w����t�{u����z���
3k
�SqjXe��m۠覣�Ӕ�l�h(���P�x�f@�V���������h�ZRn;�	`J�7pށ�W)E�H@�z3,�:������+pQYq��DA-���ٌj�j���('`3B�Y���T�Qa�8m:SS-lՃ];�'	��jҺ��Ԯ]{�*R��L-�j�з3@xU��U�F���I1CrY�bR����{�hS� ��i'r�k]��I���{��o٭b���f����Lu-LA��OF��Qi�N�͠���û��$�@7�A��&ۢ2�	Csu��-
�$8#��ähQ�Q<4��Wz�˨�%^�A��*R�ʫ�.ڠ�)���*mMknʺ�TS6�9fK��Ȣ��2�;Ҳ� �����f�4ۦ�:r�����*pi�U�����#���R��4��H���D�5�M��iY�Z�	��ĨHnA���Y�Tij��F:�� �u�m��ɢ��<p㣢�:u*��siJ�*ƭ2��MI��
,�Ǭ�w��V�j��&�l�&�J�	ԑ���E�vʨ�õ(e�x�Ե>��+���?}X�[)Lᢨ�n�n��4��(�SF���Y��C-L[�n�V��A �(��F�U��Yʷ�"p��ҭ�)]���(�	ֈ�I�P��]���z��f��Ֆ0nn���1��ʦ,:���kM��>ܽj�7������2�',�j���6�:�z��$���"3DADU`�A�:3i�M���\��w����nm���2��E"�)$�k��ø�3���P��l+wC��o܆�g]��̆33soG��5���u�{��$�d�D�ku]����S����f::����nR�`�f��~D5z�X��v�p�c��IItBT�XHfġ�1ͫ�e䙥�L7CNeʋm���᎔0�hmnև{�[Kŕ1P�G��W15�ÀS�"�X��,�]ݘ���zo6��C̒|9��]̍����CZ�B{�6�߻�s3E/s����G�u*u�Y����3��8�<k[�_{��Pt��.�D^�T��j��l�۴bzS�ɍ�w̤��b��e�n�f���k'��kCˬ���L���H��Q��kI���H�����j�k����d�&�c!W�T��w��b/6��P�E�d<Vwt9�۲�Y
+G>A���,7񼡺�5���%Z���0K5{%����e �7������ͼˌ�2V����A,B�/`Fm�v*JR�2Ѭ����_Vm��FU�f��d4�9p�>b��;�&�c���ݹsW|�uLN�\��7��zÎq��t���`,��7�sN�,��/e�,e���JIC���hT�)�짗/E$̕������b��:}�ۨY�ZJ;�� ��}x�=]CU.��fP暑GE�B�6�s'oy�8׎���3��ٿ_n�y"�08�Iǚ��ܞ������.�ݽXi�V���Ge%gS`KN�M�J���̀;*n�.HU�+.ee[�,��`�������1�
�SU
�b�
�fQR;F��e��U!_P:�� w(�ւ�:�9i���4s��4�7����6p��ú�kƩ+2S
�����! 7C2BB�;,`	��/NM�0�t�j)�x�&"Q��
Q��^j^H�˸⧭�˯���/�x��X���p�i�A�Q��D3rV�T�K-��m�2�0�*����A�K,�a�-jw@TJfZ��dE��n ���f,;[[z�1F�%�g̭9�S��LJ!+m�v�a�
'm�5ț?
ۻ������q�=����MM��hP���P�wi����6��ӵ�M��5G7T��؛��k+I�]��0F0�B^-��
�c~Q@!�Z��X(����sJe�{�G�u���r8�7�R�7��	.������YJ��oFӚQ��X��ő�h]��t��Z{[GV����f���Ī��(�R�������
�44Y�t)��f���o���t�(�U���,�j;�Fn9�&J�Y��"�q�-�HE���z��N��Tl�[N� ��y,�h������� �+����=�lmC �RH-;����y�i�����w��级�B��Cb���GE!�pJ4����u�]�S`�5gؠ��Ui飃t�����{t̷LH�:�`�(EPF(
m��ȫ��Q��������d�%HE6�C�4��14vI��m�mZ�X�����L]*�m�X�5��L�V�Q��Pi$�dX��"�AI<�����)H�-G��ח3r�o34�t���N^�GR7[��@�҈l<U�䭷�;x҂1V>�]d�Z&Uّ--� �@^�*�l9�Sww\��B.$�s8�6�;��x�N���B(�!Y!�X��PgRB�
�Q*A��b�""I�*�PQq
2#$F0`�(��A��(Ŋ�*�#1!Q`3�t�3ٷ{';�{޶��N�.�|�N�u$�ݒ
,"� U��$cT
"��1	EX�T`��EDE]Z�(�`�� ����Y�%~IR*�`�`�PF(�jaY
�t��`1��*0X�F1T���0D���A�X�j��H�1b�R1 ��
��TU
��2M0��DE�LLH�GUT�̋X�T�Ec*E�@Qߙ��?~��2ӝ��r,*'.��u^:|��8xo]�b�����3k��q�Ŕ�;�b�%��ؚㇻ�׀s���cOm�S����9[�i����6Z������3�Np6�E�s��k*Ҕb{Y:��%eJ�����0GH��	�ݮ�%]�\�
��03�M�Fo���Ը5��Y/�|%�-��0�t��u�2 �gv�!�:T�N�^�ݹr�3�H��@�2,���1q*�k�+c�U��@蛼{�2�ma:&���}�8��po9:��+<�{�'Sw*����g;�uw{&��
��{Sy��9�s���p�ӝZ�_Q7N=MU���'Tޚ��W��-T�r�ْ�^�}OK�q��hU�}�m�%xg+��o{[ݦ�n�)Vm��נ�}�r��lJ�%��*�f�������:�cV�E�B��MJ�o��MP�7`�9)�{�{ݏ�z�m��VCٔ��KzP=�q�&�4��;�Fg	�����wLv�iM��[R�B+^ݚ��������c����*?.�-S�݄hewfK��6Vα�V
�F7�]9&`�z[��oN�D�V:������L�1A������Jr8oj�H	����՗���	�)o�����=�@���t�3�и�yi\�pӻr�WZ/=��0A�<�ZN�3�d���WBY��6R��ڜ��j%�˞��mMx�����ƻ)�k_h )}�px�oeJds����%���p�X����'z댕�>�:򇱳w�<-���X&]��1B;�k��q��R�A�l��VqT�u�-�+\�LX�����tBS y���9�f�,��+��V^����*���ژ�w,D]���lNJ&.����ǗM��S�fc�=B����1��<6���3+n���m�-��`.����A�d�!����w.���{�`A;X��;ﳬ�8��c6�sy���4����{jWbb�u:	il���+��W�I���+��
�J��t�Y����=�c��Δ\�6�|��P#��kǬ}w�=J�84�����Y�i���1J��������`��p�0�jS9�4tQgl@B�����R���ݢ��(XoM������%]�#��c֓�;;k��lv�j��9o[�20ŭ�y5��z.�%�:����]��x���s���|:[�Օ�Ʉ���ȸ�L+�Ԯ�s��ټ�D(l���N�Y�Bo��yxJv��g0��ثn#4S��ٽK;��G1�7w�OP��ӷC}�$�-�-2;o%Ţ���rP�7R4ҙ��V�#����yY���F�F����׼X�G����Y��v�};F��(.�%WG*Mt��&�M���Q��%9�����]��h(���3��m�́_Z�)735��v�Էl^��)�K=n����닂� �V<��k��.U�%�n�WS7z��=$攁3� ��V:�(���@���4���Шk�i�v٩FT�M����<��1�]n�l�F�_Q��}I�F�#\�H UcR�e��q��i�^D�F�9��W�V�wj��ݱ
!�RP
�f͒]i�W8�]�|Cb�]���z
�^`��BF�Ϸ,�RY�],�L�j�2@�1��t�t����}�����z]%J�ӽ�(���)�p5��f���o�4ղppPY���q��V�����ჹ|@9��_�+�".�ͣΑm�l7#�z9 |�gt�zU�K5��1gB�*�Ğ��r��ش#�߮�W �r��t�>k±�vl�����*�de�oI�[,���di�������4`��WӚ�l�u|���ed�E>�j�_�Z��Ǘ'7�ܗ�{y�}��ՓN�M+�q�+,=z7)V|�ċݎ$�Ve���3�MvWwj��O,n�Y�@C�D8zɷ�AN8�3Q�7�A8�6�	Si��*Ew�10����VUވ�ա�)�Gkon��Px�gFq� H����fiM�خ��ŕ�޹[O,�/ xrd<�����Ǝ�B�;7�	f�5*��\X)�[ڊ��<�f�ˊ�fh��;�)z�}����B)���V0���X���l{.i�+֡����7�a�}Mq���Āl���1�X-Vͭ{�k��:wY�.������Py\\��㻕ˡ�>ᮗ�[���]�5��v�.��+6Z;�nȒ8o���R*]С}K(A�f+q<N�������ߵr��2���1�=մ�&�J*��w����F3W�E�B��%(2��k �OY c��.ӦdʜfF����A�s{�^
��.�wpbdC��2�Vtz��,dv��P͐�bMvp��4���2�Q��j����E�@��;���_5ֹ`��meExM⩊$)�������T�1X6�J^M��hA���N� �s;V�(�y˫k͆��LVU���m3�X����^��}����� ������:Qk��N�oJ�I����w�Cĕ� h2(*xò��M���@���V�z�.H��롁ժ��
JY(��-�wr\�7E��#5m�.]oi�uH>�j��o!u�L��"`|�^uA��L���"��F�݅Gw7h�Y���Wy�;�%�8��X1�S5J1�{y+�t�U:�Z:�)�8P��f˽"�k#��ڲۃl�حc��a f�ˏ�m�M�\o{��C�4wְc�M��H=H����ڥ��]հ3,:��Lp����;vo_9h8�q�:V�s���4��m�[ҩ�M��7G.f<L���m�ZyKO��l��Vˌ5������e'���!���ٷ�BN �F�j�UN�\�x���/i�-�!��Jz����z�WF_fS�C�ݦ��_�sS�GoU^�P���Ԗ�x���/��b2����-.'�=�*�ǐ�M�<�#��8w�o�u��¼�J�>Go2�5v
�lWڹï�] �ؤ\���F�uG����:9s�%����\v�L=�i�U�TYi8v�� c��J _Uw2�E��Ž+J�Jr�U\�;��ng�h�2����+u���QsK�&d尐�2,��z�-9U������nڱJ%1�(�o�n>�1�C�k����f^ĭ�}Klf�*-�f�!c�*��G�YUs9RC�0m�67�@4� \�8�rz�f��U��k/%�9�L��pǁ��)�%�\�zo$U�����d9�W|��S����eg[8JY�v��d~Ok�ҿ(E��J#~+�k �x�).���=,^�v
����d�=r -�Y��?dX���ȅ�7���j(�9�md7]%�N�D�#���j���=���|����K� P�($����q]>\��"�p\\��6�-4��� ]��;Y&��"m��,��0u����عcaȪ�vgh
1�ѵ��S��Vͅ�W�h"�Ls�r�bK��� �d�啶V��Fc�3D�e���ae��Ύ����]�#��B^��Ť��y�h�7RI��pS%r��%5��9M-Vu6��.�M��N�W�ʹ���a2����ۣ�R��.�C��|̕5ҮY���:9�J������$�Aq��j^��#�UoR�Lbi6�j6�D��ê�XƭެY�Mܓ K4��`嬽{�Z��4j�6����]D��o�Q̽I��O��Ĵ.��P=&�;�.�j�MGZ4�\I�ɚ�Y� 5��CkgR����uy��n��Ʉg�-�F*j��x1�r������'�Kn���4�l`u�j��0#�{��]����}�gu�ک����Ŵ8jw.lۜ�LJ�F�� �����n��e��Fzؙx��B�.RN��,��Y��u����v�Aӑ�g� v�o�\����Zj��奀ք�do8r������P�1,�'��CI����7��{���G=�M�:R��edۮ�(	�eG���ZciMD��0�m8<��p����1AĎ��@�]��ܣk���cd�<��YwJ����Ǣ�	����=�+�$0g�.g�2���D_Ԅ���f�Q��=�ye==c��ݤ��)�eK� �SOU��u���{�Ր;�hAm^ Ь5��H��&WP��fg"�'BW�O##�S�ވ�ɕ̎7!��oNt&g[iw	��|9֡�yIkE]5BQ��97n�f��\۬o�[Д���
�;��;��W��y���cE�u�Z����[��˨�mé Ǣb�'*�3$���Û�diu٭3t�w��iֹ�G��dP-��i
��7{��)E�̫��sѰf�ۊ��y��Z����,��;�5�S�2z���#ӥ>v�K}{�q�&�a�ܯw��C�e��-�:ع��2��+W4MY��)$�m��m��i$�H��I�i6�m��m��m�K��m��iRm��i��m��m6�m��m��I$�M$�m��m��l6�I&�����m��i$�I&�M"�m��m��m��m��l�[m��m��m�RI��m��i$�M��"��J$�I��I��m��m��m��m��m�m��m��m��m��m��m��m��m��h��H�i2ZH��i4������ho��0P� �GeԼ�r��$����R�m�}��]�z�3��&r˽ɑ򏡽Ǝ����<�N�J5nd�[ࢺ�
"�`"���$�I]�q�;�����Yn�F-Zif
�� �fJ+d�[�m�[�6;j�[���w`��PA=�v�
�hI�F�ݔSf�Y3n��EH�Zy"�6hn�Z�R���W�m�Fu0�E��֍m���	���2��fn��$�ܶ<���g�A��++�*s�N�������FɭJ��wv���\�H�Nu���8�#�b�VZ]m�B��mg)!θ1޸�;��3(�7����+e,;��W��ϸD�.��7�9����#�d��]E�l�N|��ٻqb$�x�b�tW����4[6z��*n�^.� mdʳ8�$��q��]��Sޡ�E]�mZ�X�[�
���3o���A��d��[o�;�(#��4���3�ܧ3 %j��kL�%��)&â�I6h0� �
�!���L�h"o2k(�.��]�H]�XMr�t�D��o&�-gl�cK�ol�|��.ŧ�&��Z��֨�B��gB2b���ܳ*�e��oӖ�T��Ǆ�u�m`T�����/!ᝩ��;�ne��Ud0mmS,�nﬞ�j���m���N�xѢuoSe��Չ�+�����*������e��5���-l��$���v�k�[1�r����i��ʽ�u�6�o�H��4�O�2s�\]�uֹ�E3��Q��?ޙҙ#�p�{�f��vv]Aʚ���>��r/[ ���pԳ������q&}wj���,�	b���(<Ii��t��M�9�.h�&��In�mm�U��˩f�*�eq�����YWIp�Z�h��u ��@�oa.� ��M6��ۗY�f�,�kY�Į�,�M��G��;�eWlp[{�e�1�C�ľ]7���.*�x.�ك5�s`Dɦ�w!�p�����.�l�~u�5�uf.��6hT�]��܃1.�Mʔ,��r��f�%J���8�"���ϛ9�]p��;k�ќ6w_N3�r�,y(=���j�H�ZY�H(�rG�U�������p}e�g��;ԭC�����<Jd'Ǘ?��VR��[�kt��9��z�ۼ�r3"��wU	X���l�����p�t
�o�����y�=�4���3����+�#j��{���D��n��2���gh�1��7�<�;���TWM�]�q�p|D��׫���5rt��v��Pݍ=�}Ǡ�.���d�r��c/y�;�������f8�[ҫ�l�r���ƻt�|_P���!�� �qD��L��צ�nV�vv��q�u�@���n	Lhp�9�2��R&�l�`ٚ��}�����|Һ��͔�A��b�%��;���k�W}t�b��z��*L��R�ݭk��W[8&��/bHb�E3��NZ���L�"���x���S�Ź�S:ƾ�s�6�u�>�� K�0��mZ�uǍ�w;Eme�l��:a�~�(Y��r�~�X���e#�g��A��8�p�Β�`Y��.���H��CQ4��G!�g �7���K3g�f&5��pY��{o�B�)��\�uqpaY9 �M;"f
zw��Y|�hѝY�d1<�)QZS���Ў��[��A��V�2��+�v��t��\ԧ\Y����+���"�v*W0�Y���4���`�<aN���v�K��b5��U�5��Y����Z��X��ݵ׹��R{�gwTGj`���H�gz�`ػ��]����2�$F��������j�,H�e<V^5mT7��E�m^䩝.��2��WjS)J�[X��$[�t]��]n�胥bs�S�7tf���N���n]*��E��	8؛n�$��^�`̻�j� f\��ݸTw	B��̧�f,W��t��ю�`�V9����u�sp��@JV(���C� �=�W2�CVBv>V��]x�̊��ڸ���N�Ft�]iV�������m*o��PC:m���Ҋ�ÝL[�
&�@��%�_?�d��U��x�Yp�{��O7�륗q>���9ba�w4Xk1Zȶ�S��=m�ȳ�� ^����#�=CO��4uvh�N�V+u�*]Y��O�:,v늠�-M����h��V%��z���4�Lǘh�R��1WSǳ3�7�Ƴ��v��-&dxl�k����q>�� n�`:cS��8�Z5�W�tgdu��4*��*�z6�f�t�c���7��6�P	�*���t	��D�T�Y�5�$�1,ΰ�֪�F����<|&�}��C�& ~�����I �$��@�$�O�$ �?!$0O��	 >H1�d$?�@� H���z�B�	$�B�u �2�BV@�l�T	�BCL��$�`@� Y$��q$�H� ��@;�@3tb��i �	�%`E��!4�H��$�)$' �F@�@�HM[!j��E$�d�� XB�bI�2C\�$�$�!"�:�,��3�XI1�$:��s,$�� � �2^�H��i g���>�0�0�����Bq$�O�v��Aa���`OZ���L@P�c0IL��`i	�CH�ɭ�!�
���� �g(VM��4 ��CP��`u�q�u`m�BN2T
�,`�
���'R��N�XM$�%C�dXL�̇���>��C�
�<�D�fd���;CH}l��@<�u���#�A݆� q �Xm�T1��&��$���
M�ۡ:��q'��C�}�'�Cu	�VXG��6�'A�01�~���gRc�8��L���N�!Y&�eH����C�z�2��M����|Π/�fY�lC�N�&}|��1���(q*C��xv��J���>�E���}CL]��6��L�Mr�2fXV���I�~�������>��N���>�;�E�a�R�f�u�0�Ԭ�3l6�I���Q&��;��)19���+<��g�N�����:�K����z�@ǌG��La�tW.e-i�>g���x�=dǩ�R�h{��N���� �)̰�M&�5��m����m/���M��
�O�)��3o����eCw03zɷ�J�9�v�ת����z��k��Ϸ�a�6Ö��3��!�2i7���oH�{��{���>q�ߘ����X���y�jsW��n�wl�t�b�Mu�����7Ϸ��h|��j`�cEe��Z���U�GPQ���U��ԧ����oSx�i����3(��fs{ߵG-oh���y��DV�x�w;�D�ca��Q$��I�d�G%'�c�LJ����87��6�	�znU���;W�۳D���[��I��.��n�X�'t�&:��V,��d��U��8
��^��q�`��e��X>��H�Р��*�Ћi�����\�6��o*��n�s ���A�=y2���X*�è�@IB�6�ܖ�C�0�Ή�toon}`|�x���lJ���k�)��%"^S���ˁC����(�n�Gp���4�r�a�!W��
�IմJ.��A�_"��#2��7;�DV�θ��B ���Ҏ�E�m��� �-�pr�]x�`�!m�\t}� �f<��qj�+ .rP.�VQ���r��u��3q:đih�⼁io*�:!�Du��=�4�
��V�5�v�c���Dr���-7o8��[ÕLy��]l�EJ����=eH��݊(, �ƭm�)3�C�jd��&�a�^�H�F�ɸ'�s�}�t7;����HG�4=F2�.qF��Ͷ%_%X�6;2�Y��N��c���(?���›�#C8�.�F�̾��(�Y2�j�����$v�!�T7z�J�2�dGoi^s��� wӾ�vFY�Mu��pͱHu��;U �!+�n���ʂ��W)�Ő4x���xJ[�-�T����4e��8�5�Y@��h����%��$�L{��g=l:�NX0��h8�I�>j�$�
.�F���mf.鵠���mm�]�L�R��--���4,_2�R�fܮu���T�F��{]�Xk�W^ �3`hבV��-�ۚ)*�d��z5H|�hC��J�鐮e�uI�y�k�q�3�4�����1:5j��t��;���9ڱ�؅���iA�jq�/#���
���DR(�+��W{�:�T��p��(�M	WB�$"�1dqQ0a��e�\(��k(sY�sz�X����+h�I�����J�[�:�����Nv��q�M���p��0bΩ�U��:�h4r�i<��5�I�t��؊=ۺh(^��n����'�XԮ����FN:��z(����d��4RXme��=���c&����!R�������s�z�'uuHP�3J�kuI�
�;[V��O"yBVྜྷ�Z;��e�H�����ޘ/����Zt%5Ɩ���v[��Ƙ�P���WfV���a֔)�!����Ĝ)��U�CE+�JT���rї`������=�Q߳)d�(�_\hj�9h6��.2�Jb�\-sUor�b�֘ز�	n�#h^���7x��eLC��,*%d`S4aq�Ƹ
��oF=ٔ�ݲ�P��֕׮sM�DPr�c��f����5���$��2�:%�����R�O51`;{]O�}�&�m�Sz�D�/v��DsN���6��ɵM51�	W���uV9B�+�H�&r��Ԧ�Z��\e`���K�W����N:W�P ��$Չu�Z�ʔ)j��b���C�vF(���Y�yP�6��o�-6��β�Ӛa��+�UwCDۖEG[z,]��7���]!x���n��2i��R�baoEI>"
B0�PM�`��	�Эz���F�l$@!!zc6���C�咍+�a�d�[VkF}r�.��'�>�ˢu��#����)^N����pN�h���*;���X��
�a�����dsA�ЭF�P|9	%l6�M�],s.t%N��e6���i5�))HY���Z��+9�N:�̲��i/:\��&Yi$�hLQî��oiX �&ɐ�ݡBo��P�I��qҥm`���@i\T����jL;�ӫ	a��cImݼ�Ӷ�+��U�UN�^	y����EVab���1l�`���ڨ�n��`o	,G��%7Y�%��J��V,��Z-��P8%������5�:��Z��lcQ�1�[�8RY�sZ�)�Mt�A���a����jt4����i����%�mQ�Ѷ��I�˭�w>1�gu���$�?�� w��������g�5˼��\q�W[X�������2��<R���p�ԳY�?�7�
ƥ��
9�p3w8�7��-�)9q=�L��i�}6��V
�6"(;�j��#U��i�R|�h"^����4��m�}3�ɜb紬��<n{z@�vd`j�KWr�JS4� U���Ze7K�����_�^e�R�� ˺��
�Q�!
�0e�I�Z-�7dA�]���^*�LMwJp)���;e���ie��
��CF&�4[V�_p�5Zb!�2M�[ZX���3 j����<46X]�w��Lv|Bt3n�בv»1�؞3
�m�f���צ�d8��W1�fQ�w.�Yf���<Cy/������P��/�ӽ�k=����A4*��*#�,5�*�y�P�=L.�m����Yk�){��0Q��UӜ+�X �Ib��m��i6�L6�L��I&�M��m��M��m[m��m��m��I$��{��Y�vR�+%em"%ڗ��o&�i�Rۨz�*�V�/�,$L��0��*XZ��sT��T<��wJ�d�@�2E��6ng��{L��
Ϛ�ݜ�b�����#xv�yW��]�^��β�%�d:�w=��6P�pu]l�.�wbα�K|a��Z
��6��c�4��
뼼 5�sM��v�5����9:�ݱ���Үhܸ���n�%����U���ܻ�/��ǟ�~˚�}�k�?Ą�	�g����#���	�#/0���ց �}���J/U��;����s�	��m��ff���Ҷ6G
����]�@�֒��APп�y�Wx�7.r�x��� ��C����緰�0�6�!�'�bBC��r� C'̐����� �	 i �2@�i/u��+$��H(IĐ�$�@��$<�4���	�� g��m��@:�0���$�C7`I1!����\�|���߹�ܽ�pX"�D���,X�E!Ré`�F"� ��,�(�����Ux�j�D*��0DH�"6���,��j,PD"����*"�8�g�V(�Eb�EUX�3MEb���A��"�"����TA������b,EUX�(>�X�U"*��1�Db�E����X+F���+"/���`����"ł��YTUX�
��b�QV,U]R��*����"e���*+}j1X,h�E�V1c"��P̴F
(�
���#��R�X�H��@X�**k�bŭX���Db+DQ�*�H����d�Z*(�z�QQ`�1\�`�X+�Tb���X�\�Q�QA`�����%��3V��dDX�b����F~�DUV��X&%Pb �DX�g�Ң�7d��u�UX�����X��Q]2�Db�F,EUQE�3�d�V1DVR�0b��C�*�Qb���E}J�E �><!��׶ˠ1ZLӳ�u�3ݝ���b����Q`�X��X**"
,Q��?�b"�YU����>�ڨ��%H��Ǎ�T���Q�QW(VDDDTQE���R �*��DPF+
�`�E��1A�P����ҊδU�TX�X�%�Sv�"��
��]ڪ���Eb1E���jEDb#"+�1kX�Y���
��"��UU#"�E1���m���5TX�۶TQ�O�X(j�UT���"}L�u�S�UQ�""����(�
ł*�7pZ*1b"���M�Vł���ԣ�0�U��EĢ�EJ"�*�b�d���-j���|�������b���*(+#�X��ʪ��sR"*1E�׵�D@F,`��X��Dm(��(1��֦D���ۖ���Qb�UT}aUA��kO-Q�'̣ϰ�(��1Q簚E���b��փk�`��ܢ���
`��A�""�Z��*����~��*�"0F�#���N�u��F;�D���v�b��R�gɂ*��UA6�I��������xr�]�������]������f��QAC"����C�+�DAU���"��q#�w	QEO�i���YR�;ӆ
)գ�ATb3\��\�F���j���1�~�Q�DG���f��DFU-�b�:�e���4Dc�E娏�QX�*�?S*�ۦ *��b��_�n`��TESic��I������b�]YT4��)��w/�?.��������߳�}�g�UU�h����V"(������b;e��2,wJ����*��0`�2�R���3� ��̷V�
0`��U��"��}���W���5n�~�b�Z>J�Q2�"�����v�Qb����iQ{�٭�ݢ��#���{ߵ�ڏ�M�+"���*������*���u�c�k:>@TU���Q�xg��u�վ���KIX�Si���+�AY����ew��ܔA���s�h6�U��Օ������5Jh��U\h����Ԫjت~�&"�oԣ�G;�iZ�(�ը�=��M�Q�����G�}�dڈu��G��>��F���ݕL�v�x]������߹ߎ{_�p��"����YN5wj�sY�lwj(&[�)E���>�m�SM\�T\+ﵡTE��IUe�QT�.��TD@�Q?R���Tb�˟���UG,��C"��PJ�W@��CL�W���-�wxb�C�\jD���i�MZ~�1Z�PQ�\����{��ޔ�m�9/�+\�"}F鏅�j<����ohg-�*�P��R�����h��U���]k�cYE�PQ���P�U�V,��%~qu�.��ě��eETW��e�dv�TF���z�DU1��X�]&Drʞ�M%��A\����a�/�@��[��?�|��K��ƺ�Ù�}�?\��먎�+�\��u�(�{q[A�dL=�A�E��q1`���y�k1&YK?ar���.F/֡�\�ۚ����W��W��Uݿ�*ϭt���MclQci��޾sBĴq��:p���� hsT��� PL��.W7�o�4E2:A��v+�y��sn���R=r�u�|�)��ܽId�7������Z ���;���Z�@CY�4�'D0��/^�|%�=iN45œza5�����up�e,o���(�/}�}���3�1�6�r�e����ف���c���*���3wX���F��\��L����%T�a�>u�5��ӈ �Z%�H������т�*��j-j(��n�f�A�3~�&��.��&�-�����5�#������!U�-��d�{k1�AVT+ό�k�^�����.��]�����;���r[_Z�{0DX�c҉�U}�|��b�����¢�,��PEq�����X������}y��l��4�b�ZcG�*���J�F/�R`�]ۊ|��*�lF(�Q�ӺsB	����"�ƣ=��� *"�������'cx�ޑ���]�����d���B����?��/�&�N�2)�*��1'�W=eD���w(2�TGb��`�O~�֙U��j��)L��������G�����*=e2���TuB��+�\ۘ'[*Q\���N%A�{�ت��8�h8��~H �*UK�
�^�}γ[F��{���c���k�L��Qf��բ����5f����U����Vo��f^51��Qb���<�n�2m��qG��h�����D�_�������*u,q
**3��Oɴ�DQ�
��ƃ�{t��������xUT��&���/�qo�^QG�� �*nʊ9q1��}��)�TԬ�������Y컴S��_�I���9o�UGW�����h
�Z<�O�'�ܼg�9J(=����|�ݨ��(�>��6)?R�6�]j�?kzUf�T�|����$���r����]w�f������9LGv�N}ܛ".�w~x�m�7��&�*T@cIE���M��X���
��7+��1]$RYm�x�*�R��U;oŮ��U
��2�SV�Z�2���f~=��T��Pwx�|�B�����׵�ﴡ��w�3g`�����Q���1
�eEϵ�5E_�>M8��ȸX������~�z.��S���Es�?sf�EV�m��^�ۼ�+��1�?o@��wq�j����q��=��:�
TS�ڱM5�V(�P�n�t�$���;�#٢ϳ��x��W�Wx0U&~4� �D�+YO�U�ջl��:�3ق���k��X��Y�L�9M�͚��*"������3
�;w�?h�j��t��}�}�w��i�2�_�1�_�Cv�m/�M�d6�;�к�_�o�!��}w-j�����2�Z��a��j��Uv�v���A�����t�Q��f,�2��
����pS3F3�M;�����
i��
�ʉ��~�98�Vr��d�a���f4*��W޺��[>�;��P*�"��2�6�9�~�t�3�r�3����Y]f`y�'-���m�M<h�B�D�^&��ޕ+�&H"��f�a�M��b1�I�뎭��M+�q�ֱ;�q��]�Vr�?j��v�(P�|<���G�H���r�r�λ�k��a�����О/Ohĥ��ys��#i��/u��|J�9A�.�&���·�� �d����)���|�u�3�iB�=����.����M��ȴ�u��,�*��*�.�m,�eiuӕqԍjɌ���q�=bܠ{)��TȺ��U�[�DO���i��H�c,T���5����SN��T�:`V��c�/s1Jʯ�&9�ֳ>�.!��k��a��k.
�'L��{�W�wZ�%1�Q%h��ٍ���O��\�~�j����<̛~4�ޠ������C����f8-K�ϻ�yt����>2{��� �*x>-4h C��ϰ1�jw8�����M�)i~���өA���
W��Lj��4��e�}��c7����y�?~3�s��-����~�/�2cG�X��'��3O��~l�E�\k0�}���[�W-D��~��sbr�4b�������)&�Z���+��-K�_6}���V&��iε�?���yt�"�rU�����ы���Đ>-�o�n��LQ�i�;pR,1�p,��b��ti��l|�A�������:s�����-+�z�����aj�g�S�o���_�����*��$^v�[^�����u��ޣ	�f��"/�����ut�շx�H��
B�£,ѵ���Pp�����B"4�$j���*�����e���N�z��L�ߞ;��h�[=u��I�}^t�N����g�p�������d�����oiQ�h�� �Z����K�t�B(1��Q���@#^%��ND��-�A��>3.J���Ю����H*��y���󼽴t��U3y��t^��� |s��F�J�?��t�e��տ���N�r�֯�fw�\�4{�p����L�}��`
��GI���  ��V.D(
4C�F��`:�V�����a�/;%�
-���h�k���µ$���$}�-s��2�����s{>aU���]�A�5l�\z�m��a�Y�Y��*��!�Y�v��|�#@p�e���
����o�b5���q�˰��'V�z�����G�l%����(�q�l~lM���z�{6E���s��󆬬F��R��󘇲����^�th>_ �b�*���@i�������SA����|�K�������CԺJ}��4^7�&�}�ۧv����I��B��M������"y�����C2���k��ؾ���O�ϐ�?x}L-�D��`�p6ϲxi�fۧ|Bv�Ԉ��ǜ-��u�.��R�\��+����A� �qP�ms5�r�\/i��;�}�u˔]��o�N�4U�d��+��H�6�m6�7xm�Iպ�F���йOQub���eوJ7Š�Oq�nK.��ת�xis���!«!T����w���^Y�UsZ�:�6�q�9���6$ ��ӿZ?#LF�c�Ő1T�:��J�O�i������hW��*�]�C�:�N{��L���5��q��o^M�J6�^%�~����A��{=����.^7*�+��
aM*}��V�fO��9s��m�f������n�J���Si��o�o��*{=i�p+���}$"�z�j��Yi�M����J+���Sx;��@1�	 )3A�WJ�`U$�ɵ�R��Zm�$N�*f������>@�)(}��;
����d�Wun���Ձ���T��"�D*�~������Α���.5~y�*�P��f�?y�#4D�^٘~�����J��(K���ғ����o3mq�.����Ό!���E!�Ѯ+�t( G�@����	�i�X���~�H�!Lk� Ю�&4B���r �D�D�J���f�@h? i8�i�"�J�7~7��U��yn�~ě�ZY��wa��U�CSo�uX�Ȑ ]{����-��ܳ\=���������6�j>�^)��x:���e4�9Ԥ�����| `P�n0��w;4 Þ�e���) x��Pm�,j8wJ�����u珵�KxoX���^%H�e*(J܊��'�,��N�@s�T�EL0
A1H?��T����k��;'?n���I�f�H7�(�tT"� 24�P�bd�DM*��P:��T�
�K�k�x%Պ�*6H>�hxt 1��� *T\�$n���x{��}�j�����T��dbE�9Q;,���ϭ���J�iw<�}�񐺸�#����^X U�6���|WۤHK�2���Ř0�m�� Q��Ov������&|-R���Ѹ(�w��0�a���dӘ��8H�7�a\�J_BVj5����K8���IPv��!`�D�(�4j�ay�|(S
%�C�U����Y��{��t���0�����ϖE��mD�Bׅ���ن���&����i+e��7W5��4@�̼�W;s�|�S�YP�xm>��N;X8��\6�;�W#e��tp�7&4���m��o8���Zgx��:�z��sWiU͐9�z��IY���E{d������#h�B��1�k��e-���G�Gl�����<�/	�	F
Az�zW��),!��H�J���.�Ԙj~a�p��w��Br�y1TM
�m�:��Ib�v�BU��R�v��RIR�i�!@;���ł�x�wOC�v��P�K�܌h��x�A�{���Se������Ρyj��4�*���߭;�e�)B����� �\b3��^1'i�î(���Y3���B��������+�/��込�3gǷ�%�.�j��q�X��i�j�cA�@��)Ys̷g��>���P���;���<h��}h0�D� 4<��(�ɠ��R	�:��K9�7�D������P�eb1�pUg��
X��*^}p(�s�K�E4I�,���\KQ���>d��(�5��"ᯌ4�GH�Ǒg��^�E.�4J�b��Bg
�4FXJQ61�����a�pV�{@(
)*���N��d���3b�k�� C8��An��|���`����ǹw�UU�s�qh�����w*��I�:_�6U��p�`G�.��M�t��H�@�((K�Z��|iҍz���}�<��ύ���(���H>dP�#���.m��yr��ǆ��>��$N�6#UH����%���n�$ >[S׹�_��G�o�`�ŭ�^_@�i
������o�*��1@G�o���{B[oެ��g3�n��u�6�m!�<+�ʊc��?Ta�hΠ����v�Y���P�+�N��'{_]���B���T��;�eN�_n��:3ݸ��~"�Q`m6n � ZC~_�t�)���87���e�h����[Ƙ�@>���! ���lP�����=V+���a��G�������iW�A�\x{���O~��� c'7�	Y�<��xI	0�Hw|���!&Z�w�~�Hj�O��  � BC�C m{��HOk{�>��ΰ�hH��<j��}�����bBM�!��Hf{�Rm&��b����H`H~d���w����}���9{Ϻ�\#�V�9 �r͂�E�};Eb�k�_1�s�)���peqÍH'=:�ާT;w���/X7}�f�y���E����͊�@�L(!ʆ�a��	isAjf�#P}�`Zՙ��;�w@AO��x�lYۧD�I�L��1}N�t��w�P���>Tw�B�+A�Z4�f�d
���xִ�6P����k��Y�X���6�>XT*%l5���wƺ|)Ow���5۬�:uy�\*��w�:�P}M�O�p�k1-~�Ͼ	8W�Vq�BswCªǇ�k��D�5��u�i�-k���E5&/W^����n�p��uuKۺ��4�9������� BD�`� jt���?*_[ca5���yV+������S�	����y�|;��o�3��É� �{�ʴQ�^�>^[���Pb̽��C!�t��0�V-<��lE�ۻ�l����U�V
I�!�7����Y{�����t�bƧ�>��}\��˭�� y_���Q�^T�����(�G�<s3����m6:� |�+��,qu�kUr���[����� ��W��C�j�~�����Q���
tn�0Ǖ0�de��򥠑���B��c.���4�n{@���B��J'��E�c�պ}��T�G��+h��������U��,@��ɨW���l���� ��F}rVʸ�?6�  �¼��.y��c���7�Ii=K����s4�u���<�{&+ҡl:ڡ}��dL/���^�U
Y}��-qF�(ȑ �~u� �^�i��W�G�8h^?y��*~�-���p�E%�s���!�����H٘Hu!#���%�]�*W^�F�Xl��g���7����￤�מ�3=_��1�t`Nx��oz��w�����z������� oǴ�}_�wS}D��m���y}�T��X�;��}4J�7���]}�U��Uy�o����05�ۯ��ڴ�u67�b�\$�7f��:�|:[\�N����E�Tg$�jl6;
kn���F��l�g�~>Օȭbk��u�J��d��������N��Hyy���
ШVx�k���K��qz�����()�R��D9��廿��s���g���י�a�%�@UP�T���^�{3� �n��[��	�n�znN����
@����8��I5� h5�!I^��O�qA=���8����s��}��TbÁ֌�������79�%�f�9_�w+�.c����ͥ�q�j>mQ��4�q?_9�<<*�X?9�ExZ�WW��~�^+����C«w�AOVv��0y�z�_��������d�L�>�����D��e�b4?�C�A�KP��O�PwQv{H;���U�51���)��ѣ�u���v({Ýh��ꛦ>��^�+({]�<(�&���w��Vb����.�*���5��a�f�3�~���L���?4�
��P�����pit�O���ѵZ:�����_��զ=��#£(W�.V+v���R���F@���ЭAYT7`@�q+,P����c�׶m�1&;�.ļ���ۻ&�zM���h��4��
~u8�S�\n�
�H��"I�dCo�Q5�� �<�]�Pg�iTݏ�%��@�e �
�HF�����(������/�N*��~��eP
��p�,Wv��29!��R�݋J}��Ց�lv%χ���R���WKnQ���mVgUm���6�ԧ��>��7���*#;o�dZ�G��L��tg5�k�Ivn�����R�#��
:�	YJ�n�KTJ�����O��S��yy6i=G���z:�+��~W�N���t��M���H�j�I�AE��uۊ(|��:�����=�J��7ӽ���2���]��oM(�? H�=��P	��8+�X�s��Z-
�mӪc��g&��6tS=6s3a�bR z�IiU�E�W�O����_��+¦�փ�ۻ�Y _w�{�h��Z�-��+�����ڽ�QQhL��kB��&�#���� �h��<*�u����Uz��7�J���0�s�:{�K�K��ϳ�����Z<�b�s3
w.����k�Ti�AL
Ϥ{ན�s�O����b_o�TjN�j%��y�c�U�fO�^ªkP�y;C	i�J����Q���>�}��6+Lo�|�{�n
��҅�?��մ���Cؓy���*�=�Ϣ�^]��Lz�@i�7�o���B4M�l�\GRa<�T>xyS�F��̷�7��F�v���۔3�Omap���%P�Y8Ɖ�U��0�b's���M�LӤ*�����v�>������ޞ��9��+"4!�s;�b�Q��x>F`��Pq���/&i��*]�=^>�+k�I4�N�o�.�%���q'�֞�_֦��Y������}�1:|���Wۭ�#K��G�[�O��$�����_ݐ!n�'�q��&4�y�k����_u?+���ON�޹X&ơg7���>�@��X׆� uB��6�+4_����RsV9+�㚰̴��S����8-��m��
�g:��v�n�β��cu��O�WI6NU��KJ�x�VWvm�y�vw��{���1�Cq\\TcqN�7�u?�������5G�7쿇�{N\�R x`��8���ָ��z!�觲���ۙ������$mq���#3'�ښ�dt��d<��n>/��#�?UѶ)[z�`vU�}����L��knt��0�|�������,��{Ɛ���S�v�"���C��w�~ޕ&�u󥁃_Yc�laGP�����������Ж|epڸ�@�)����P
�T�e��������.�A.C)��o�+�|jm�8���Y�᫛����¨N�S�n�����S�J2G������z��/��d����Rb$��P���[��y��T|57��Uog�(R���V*U��+��U�����C�X�ZvO	ɟ��Wݐv�x}�]��V�u�^�'_z�̈́�p�=��<��/^��|U�7:��z�X`�4Ċ:�(��YO���Uz@�H�3�5ҕ�W�p���SAL*�~ؖ殖�5&�7�j�گ,�菰q��^�ī�^�}��tX���^T�,���U��i�kN�-F�aY����2�	)���'����׹G@>S9��[���N^s�*��J��1�\�Ӧ�:{�@j���]aū<����z��e�;��̐e�F�1���t�:�`9����F({V�%��JwNb�=����.�{2� ib�ؙ�y�����{$���b���W�&8�R"�h��Z�u�l�\�s��ɩ�ћL�;X�X����i���!��r�]���;�GO��7��%�gP�[�ŕ/y��(�������1\��%$�K�~ݢ�{�
�Z�u�9R_FU@�'1ɷ�M��/J&�x����%���z��T\�����\1H�:�%VP��^�B�Cu����*��ї����t����e�΃����rZ��#>�u����`��B�Zh}v��'(g���_oX��(�����-��������O��%�_,e�����o�}�-��<�<�ǻ�u%m� ک��C����RyX�-�1��8œ���zS��O"�8Ww��o�ڽħC�D�q�}<R�4�/k���N[�J��w��z�g({h"�����ӝ��{�N�"Dftń.����77�p#� B��q4�r����Ff��)U�G8op#|��/=j�w�*�⮸�v���>��˗^���M�'=�u^��!Ӭ�^b]��f��4�X 
��K�:f�G\���ՙ?$��׷�!��QZncB�7GFWo���a�m��E#�=�Yr�8m��Vr�l���T 1���U���?H�b�3��Z�fڪwUq�A��-cU,_f���e��a��v
�K@X�ܫ쯫�T	,�י'�_ea}�G`Oĝ�Ú��Xo[���J�1BG[�vuNo/bM _�U}��R��9_Sz�+�cP�}������N/���e�?�9��[���B�><<1��kל�r���ܦ}z�S;N��xe���xB��}�7w��udy���R���4����L�Y^�kzX�L���F��Hn�O/�~��oj{��ng�y����u���W�y:IB��hV.���i^Q�{�kj�m�q��W�Ϧsg ���-[��
h�L�d9F?��6�W{��
�������h�5���`�
j�aF�����@�C�Z���E+N�Y��u��e�#��t��龬�O8hWk�B|����ٹ9��~Ej�����y����H駎�����B�|fn��mZ��ա�wDH7II�����Ѥ����+�[L��x�g5Q��{{�nw�X�Z�wwWWy�9��݌N�0Z��J��xE��lz-��Ֆ���r1���ԬG2�>��}���%qY�JV/P���kג�Kz�Ĺ���e��bp�#��j����z�K�Uk�{Ӂ�Cs�W�e�~�cq߭ɻ���9ʗ
��+�_M��؆ �~��hܦOW]��4�}#����9}{{�K��ĬvDX�Nu�Q%��Ȯkmi�'���i
���7үc3FLʳ\�>����K6N�h��X��$�HX�p�f�a��v��5w�]��t��U��Z�ZG҅�lF:���{�+	�r���7%����1��."�"<��/�7#nՇt�Τ��7s�8���z��;���1g�@ᶄ��Vͽ��wC���2��>V��uf�	���w��Z���kɪ���.�VRI��ۅ<m��M�b�Z�e�E��j��wR���k��"�I�]�SfFNJ\�'}Y��D+�R�v��O&�
g]�r��]/�rh�J�Vk�:u��R<}e�ܧakڲ�>{0P�"�����q��cC��yHe�t�o��.sB�]�-q�W#l�/.ѻ�WQ�(��:"tkǹ�j�)8�V5�M���K��f#�_tYZ�]ns۳���;���f���.��hQU���H���� �����6�ͺ:1kD��8��7[�+ɉղ(h�� P�70�(�58��o�*�:K/�>H���|qO�ܧ4�j��F-����K�W��<7i�\�p'���S�� ��Nn&9���]D������=Zf���CPԮ��z��W���UJ%/yx%V�g�X��=[{�/�r�j|����][���&S�n��G��كt����M��ޗ:����1श�	vcW�y�ϩ
�s���vR?P_���-?g��q����}f��M!�������*�'r����C���)��e��浧L����b'�b�'����tu&�J�}����*"e'�c�Jw����뭍̨ʺ����� �IG�B��^��3mf�i�|a��*(��NO��iP�PS��k����&Ę󅆹eEL�3�+o1~C��g9��V��O��3��(�穇��ѭ��N s���{������1��m��vHB��A zs!G�'7�%a����_����+:�	�Ac��0��o�6���ϓD�P���~ֿ�{8���`����Ԭ��1'�8�I���:}�Q�Ong�<z\F�#�?~h�L�&��a�jg�g��j�0�,��w[�(:q~��f���6~шk�O��M}��fٜ)Ҍ��9�J�-�L�?w|����" �ֳ7��T�J������>����ų[�ߗ���L1B#��џq�����Ci�Y����C�3W���Mz�T�R�֎$��
�����?��ΰ�-��AUE벹�������K��/l�<e�"%A�����?��E�*J3���>������m���������T��?'�m�s�Qf�~��4��q�q*;q��9���aG�j��16ʕ?kXk��R(�J��X��� ���B2b G����9��$�_��;�~�9��7�135�k�_���-��a��X!���#4p�[t˕�y��S�����8���j���M*^��>�^~��9��!�A�E�5}m��y��-�X�����3TP���_� �<ɺ�'�����>��(}̉RE�ܨ��2�p�D�8���뫤�|����3�&KY�X�]���d�v)��**~n.1/0�oYѷ;����f0F{����Pp����(E�9����0`�����3DMɽ
5g�v�v�m,
ڏAů��Z����M�sj���f��g
m�-ˀoWLK�s-u�H�ݱ�����C*kss\�WF������V�4p��) Gv'C0�ut�Z�+**�'���LX�P(��!˔��2���,�İ��n4}��jncl���R��.����6;��G�]%�3ן�՝z�a�����`�_ru�����<*o������p�����{���1��J����9Ҩ�~�;�~�A
�*�Y(za���U�G�H'��׽S��	�0	�^	z�$��{,҅v~\ϑ���犼�7�Q���/*h�=�LǼ.~�4g/��ꔰ���������#��[�����v ��9��I�J��9}�L|`]�?!�|7��=����Q<gxt��u._�[@7/�s�1o;����y����W�C/�JR>f�4?e}B7w)�&�q���	f!�=�@ݫ�MXK׵����)�����W��cJ���#�&p��A�t!/��m�؉f2��u�5�iD�3�I����>#%yQ7Σ��������w8�J�����yQ����=����E6>b+5�9��f��|��)VwrW�f���;,�i��T���qB��
]��tv�;cF�� �L|��bX�v�.+7b�Ŭ�k۞��4��q�5���0U�2�Ulk�u�#��j�~��ף����$'���4�3�4�f���'D����TY�T롏1Q���׺�55��"����jfeF�����Lv��W�$��.^���s���4�m����)#�����������PG3��C�:K37fn������1�='�eeg�>	b"j��������=+����,U�m��~j%�G����►�X��U~uX�?����u�m�ʑ��������ʗ{���ձ��ޯn�<�vJw�]6;�y�c1튥q�*�I�H�l.W`b+3MUL������o��нTɩ�L�Dx�S��h�x�&!bub2�k��0����F�9uB�=�
&;B���8?�nnf�ȫ���� Aԇ�y,��Wy�qCD��Q��7��#x�+ͼ��
#s�ן�nZ����5���5�.Ѿc��M��1d���{>�1���G�_��-��{�`9_��꒜�ہ%��1[��M�~U���:(*!q�~9Ծ}+
����*�/�tmB������ZWθxW�9����G���$W��wS����=���"]NӴ��k��,W�?kqz.�t���q�t������u��(�C�{^�׏��7�Xfx�^�
V�&�`�ޙߕ�X��E�j`B2�2>��c�����|ޢ�P��b��땱�T���|�����~K���|xU�Kt�h�}}�.��C�
�� B�;����"C���#�;PO�F?���������R0��U݈���;9���~��{��yӥ��>�n[K�E�Zy����L7n��]o*v��VO*��oyWY��������������7[:[ƫ�KB��}w�t=��2�_+T�Q�N._ؓN�hj��"�W!�u�u�ƏnԢ
�3���2��F��󬵗'Kq��"��¾U��?n�F
��F/	���l���E@xCGN��ᡏA�>V+��r2"�yg �7_��{:��g�2���6�A�ŏ�$�-~�e�{,~��{"/ե#�_�a���{Z�v{~q%�&\�+��Z�S����nVD�n�1�;��� 8F"�3Ć���^S�%z����|�����E>?�P8��`�`��� �*���On"���ә���6/��c�ۋ���8z�v0 !L�kd_*��\"<>�G���P��}	w������w��*;�<&���f��U�i�b�=;i��kl���H���V8 V����'�xH,C����]i���G��37͇d���^�߲?k1z�v�k��f|�]2x�B�0����׺ -[v=f6t:���/�<�&���}�����m]��\'�f���Ypf��W��^˿-�}.�e>��E5Uh?<�����V�zw/,(�D�W�ܪpV�������j�#��b���0'(z�����h����p�=���it���Ǫ7�L�z3���;CD_M��"��>�hOUtT�;�[Q�U�X���O
��<�{�ё�_��O���tQ�{��\=���LU��#[9\�֚����9�su��}�'�X�i:A^��W���P��yu�٩�(��b*vf\W��ʷ6�6��t �V�^�遀�u�;P*g�ڶ����=��yl⑩C�X�yW�U��Le��0�l�Q��a���7*``�&�b��
jE[�J�ur�������޹�q�����������=�����#�4Z?n�!�G�=����Mo&-
#���H���[��|1��c�V�I�9Q�#@�*,�B�f�X"�
���+l��k��o�=9���nJ��m�N���[��\7|�]�n����~Wp�����Ĉb!`00�_EF�t�c dߦz�E|x���h�Y������$J���b���,>8`��r\�b�.�ѐ4}v�d`�3<'%�y=��e��wuH�U�eŧ �%��샕��Ɏ3}�60}��:����ޞ.~�u�X�� gƃ>��#�w��"�����ڛ��O�b<��N��>�VcG�<k�{�F��F�g��:~S}���b4T�һ��޻�*?��0�����I�6!��"���W.�/k����.�N��z1�>���C+�'�
U0�*�~}�5볱03��E�&�1&�w<�������O�+����g�
��/T��@K�]��K�K<:v:�ړќ���na�Ĩ-@vǖd��Fv�o+Av2��F�K�xqL�g��Բ=�Z6��Ub�C6�A��Sa}��,��=Ś!镊��+I��^�ۛ��9���dN%�(��2�}S�k��e�	�MKS����P���w.ݝb}��~z�͡��)��x4noUM���Uh�s���iX)Ǧ�ʩ0�b��}�^�k|�>�^�~7O߰Q�<�c��efo!��`�41
�0O1��+q�U�Y~����t���ZH���IS�5��}�qU�p���U�1���Գ��'KU�<>
Bu##�e���OFcZ�p�-��e�/���_?��n+�G���ç������_�*̦����L�`�1�s�ٜ�M]�R�we_�G��S���b��P#N�~w��2�ʼ��K�+��qJ$ky�f���-]c�7��{�rO9�<2v~#�s}e���0>BI!�@���}�|7����}�}_��Ӌ��O�+�/FݻH�?��^�h��~��o�U���w�1�Q�W��� ?{���V<�匝�s�;v��{*lꂃ�)rבB]�d���z��@Fu�9���4SYU���KB%�mZ��UxߣI�-��v�xHЉ��m��.��b�R�77T�h�E��t�~5���߫����g�
�����s�:m���3����ر��A�=����_j��6J�c�j�FtE���9��
�t���a��w�{G>��Ϥ3���R��'�h�e��N�e��-�1���vj��8�Q�1�u��cY�km̡o�����͖Tٺ��p@��4��؍C#�n���V��������ô�6���ޚ4�HEZx�q�t�Vf8��0����rVI9�/�aj��O�������+����L�X�!D|�V����C��؎~;���*�(�����x~����Nţ��P�/���|e�o'$�;��p�n�d���jDY���vH���+�9�O!r�f�O���Gj������1U!�\��g�Wp�����~��'���pUj�,�z��0M���~}��Ϯį�W2���V4*��O�"����yp���`����[��fcZ���ć:��\@t�-��]��3����x����#{'c�� B�f��3�u _�����Uyc�/�����Dҭ-w�뭕{6q��j}iN�.���P�Ǵԫ���R^�e�t'B����y�xԏ�w	{�JTT˘ �LB�9��eщ]w�5�kY��m�� ��T'(v�ϥ�䷪�G# �߽��*7�5���cO�+�b��*S��D��Q��&�g��\Y�L�է3���A�o����ߗ�vª
�&���c���jz.�էw�(�
�tVjv���l�Δ庂^�K�]B�y~�[4z�T�c����`ey8����G�x��%�?��7^���پ��g��*�'̩�]YL�v����ٕn��]���GmK]��`� ���(��s�"M\X0ٱ�:,`��y�:v�Nw�{��pk�����k�Vnc�o^�M��.�J�yO�Ǯ�|��6�����|�zb�B��<�#˽�ﶶ~M�-rG��f>	o�<N~���[)��1t`t#�G�����ߟNΚw���Q"��>հ�Șl��N�x�}427��w���X������2����E�g[�L�w8�,�OLd��K���$���<�৛���u����%u���kÌ9�v��S����#1�V<7O�;���c���φ�[ ���� ��<�����<���<�W���VnF)z�V�}{�"��p"$Msn�g�簞f|j����ϻk�/aΡ:s6BD��H���4��w�w>�V_���z�����������r�V;����;����u�H�ͦ�:�gkn���B����⚿�˗��b��<ۂ";���$sN� �2�mgF�-�|VTft����
�8���f[�"p��)��v��������i����!��/v�j�����B9'm,}.�!w }�<��9�k�4E�2�`xY?6{��^�=��NJ�/���亞���x~�TA��qMl(��I��3����s}[�Ϩȶ~�g��-Tح�g�ĺ�����i�r��t��Z��OW�ng5Y��y�.���Gm^gX�ӇX-�j���Q��ųL�\>ή�{w]P�����`U� ��9k��u�S�[����h�LPN���Ga�`����8�o$V�2�LB�Hҩ/�դ1�^��6��v��;���q�ԯ>r��)���V�Ml{�T�R�Q���Bˤ���Tx���j�峼s��9v8��FH��������W��K:�r����
�bY�c��*��{���Zt����;��;�\%N����g;1܃N�D���Tp����#ur�Q��;�sc� �x3�=;pb*����)�����-��Z�hA���H�TTV(�@�c4�vg�J�LX%K�WD�*v����)I�Ы8\o��^C�7q��o��bW�0sɅ��B��Lƞ�[�Euw�+��${��ˮLz�Vܫ��O��V���ܷ�����j;�#жthc�^u��'�0x@7����i>���ʙ�'l��:��!&ݤ�H��>�GN�OV�AfD�n+:)G�b��v�80�.�;�I���н����p�:��d�K.5���R*�_���T���&��̶�y�$�[���Ȳ�oс"�o�_m-�1��߸3פ��4�шy��b�z��ۍ�UV�-��l�û���b���j뺲�ycn�#��F� a |��*Ӄ��ۿ/���ҿ)e�绐��{�i4{J싃bb}��3k@�1S]�d��j�a���)؈br���	��T��le���Q�V�q�:Y;���=Nkɮ;�]�S������:�Rn�h�F=0���!�w^p��Y��3
M���L+���5�UfZ+�f���Pf�~~[�5U;̓������>s�S��yQǝP�U&iR����w
M@�,,�j'��Y�����2�{O������5�E���b�ߝ_��JzLTڃ;8�FDu���#.��RTEw#��ۚ�Lī{:S��)?�o���������u:���������]h�}��� �|��L���x�te�.`�a��j����1�^�!�3kc�����;�W@�ǯ|-v-Aw��^Fp�IJ��)���;�^��J;>u9����ʂ��I�a�9w�רV�9)Z����+�.*ǩ?X�q�5w���]hΦ������1pzvb�,������.�hB}������G-�DB����}�{���;r��r�ϖ��d�1剨��m������m^Wma���x]�\��bC^���G���/2�b�U�ӏHd����Z��w���W��eś��Fr(�ɾ�޷�C��29;��v9�S�i�̘�@b�)왠R������5���us�r]���4��a��˃4�)yר�T��B�Em|{�(!B�޷j��<��*�έ��NV�eO��׼6�U�T��8>K�]�cQ7ϴC�Z�<
n#݌.��Q�{M��Ctqo|��9r�q�#��+ޤ���;^
���j�U�x��wP楷O�b�[��u�F�P�b����u]�����W.J�6�BĶ�ݑ�,�p.'o��Ј�ڱ��N�N�Ǽ�t�L�ӏo�ވ0�l[J�vCn�#n�+t����_R�w/ws���u�������=�V/�m�._\�˾幣΋ƪ��{��=�>.SB���$���{�qf�[�{���T�U�ـ��,��������Y]�f�A��8�k<E�j;���}�d����KYAs��S{y�]Vۻ1Z.��c 
U�W�}��:@k�\��M��I�4�#8F r�}�	%�(+N$�'�'m]B�(<�b�,uhWB����a$�E���	k	� O)v����}R�v���&K4(���CJ�i�6������.8����BH�]��<��tF�a��钺��8d������%���w����re]Y]��3�+χ_���z{�����:�4�\b�*�&�m{d�@0�.��)�{Otm*j� f�aV�{�5NZ暙�w�MN�u��E����>5����L�fFbȦ����w�^�=�R�+��k��]DG��vt����K��r���̓´m�T=�N�ԅ2��n�S��X�e/bڱ㸝1V('~޾>�k�{�Đ{��k�m:D ��v�������W.�)Wʦ�J���9�z㠁�N.K�Wb�g��v;ދ��@O}�bV_ݍ�E��j��CQ�YZ{fo	&��{���I�\��WZ�H+�*쇹�K��GoHD����}@��}�q���m*9��*��ahM�g%b�A�;�����9���$��.̣�1�T�)��;!����k{Mͺ��7��L�;v���3�����L��3�Y��ց��O������,GNo���Mˡ:����X�WH78�yD�i�4[�Ws���o��6]Ѵe>]�4����&��}��]	������ݴ��)����� �}j��1�O���;����P'�Z��>�k�E�˱}�ͺm�M���C%fgEѴq`��QS���Ў��0�}��Y-<�ǵuy]���Ck���m��i$�m��I��m��m��m��H�[-��m��m��i&�t �J��)ps�����-Ԓ��}if7���v>�$@���%n�;-Z=Y�N�+ đE^�n�Vh�_D{jv������Q;M�uw;��זq��tx�];�/�}�dʶ��;�PN����&YN6��▜U�n���"�$�&�ض^��x�c#�wdc�@.����O\���k���-*|���B�뻇2�;�*�R�l�0���f�w���^#�kJ�A� t�ດ��{��tx��U�}_N�;u��z�y��'u[|]I�9��׈p���vLꩅ:w��ԉm$�m��w��s8�� B�L.$�b����q���z��eFEG.^2v=K?��I�g��]9��WG��	z~�i��_���&"a��o\��� `�Qc�w/c	��B=%�f~���M�s�쏫z�c߯ޘ����f�[z�
5��~]�d���a�w�ꁃ�*g:��q�އ9ɣ�4Ɓ�"��eĈd��+��l�s_g�ʹ�i�Soj�5����{hH�}�L@u{�v��+�z'g�Vyd3�w�,&l!�Oc>�ڐUp�k۽���W�hN")~$}���<��U�?S
�3o"793q,��#_a*��1���enTM��Ю7&7 Lt�]˞�0GUW�Ǚ`X�O�vD�����a�FLuy�����5[W��l���Q���Y��edn�1?|P�)q��Q�7P<��z69(ꙫɱta͆��W�cF�ߎ�O,��-rw|ו.�o�qG���q��^WY�����fbz�ē{�w�=�#��ݽ�"A^�l_��^������u�F��{Nʑ%]�M�-��'z��F�}���Y��!i�W�J������w���1�ɰԋ��~���(/:+���x0_A7Zw�{v�r��W�quR	�x��];�X���wq�P۽�ɪ�Q�X�G8��|*��Wl���y}�*�L]�kݹX5$ZS�����f3]w��Q؀_37%wV�t�����;����C({��`��s�ӊa~�3�g;��nG�2��Tf0t��&�1�m:Z|���G���p.�V^��"	S���.t?4A���b����Χ�?�׋b�.��*��޵_l#���^����䈛`DgMG��v�R!��e�=�t
���x�����T�bԯ�15�s����� ^�r;8�>�؝�Y�0\��J}�V�;��s�������_���¯k�<�8��`�A�u�n+V�ͥ7����_��ĺ�Ե��(�j�3L9��ÿ �	�5������I#�͒Θ������j\������;��*m�߷S�h��.\����~�����ٺ�&^x��Ý7�v�W߸����xS�����c�?�����SÞ�A��~���c"�U�S��mf,�Xs�G��rP
:�����w}����h�E��1����$���ᒫj~���߹��j�nH�s�������B:���?D�*ovʿ8=��8}��B�2}�f#;e�
�"|b�}��N˧Gݷh��}����ڰ�8�j=�(��z�+����wr�뷴��N�����&�ݫN�:�c���<�r`BDf��:3n ^E&�2w�����l�0E��`*�
����@q��i�`|���9v��쩕�W8�"Յ�5�7�C�����\!#�m^�(����/�:�8{��~з�B��ߣ���3k~����,.�y��R��azB~V�J$�MƋ�d}t���>�-���̥d9"_�ewÂسS7Ts���|<��k,��5�
ҡ+>~$����kt#'Ǹ�xA)���'`@Z�"�b]�z��@�D��]��h�4��'��{,��u��[��로k�������eu+9�A�=�x� }�rJ�U����ƾ�hn�O�{�ܹ���v��]h>�y���UD���uU��fA��^�uz��bl��9��^�^����W�2����OLή�\�|+�z��w*wr}�\O�zb<<ß��(�{���LI���?����ϕ��d�U��8R��=�0J<����ݔ�j�z�Ҟ��Z�T�>��z���I�}������׭0�}�v���UӋ+�K���r!4�S�O��Q�%��Q��S�ײ����u*:s�����FE��cB�9�J>�s6�{��]�����o���X��hX�s��:��߯�^˹W�#����1K�
��ia�����tM
ʳz�G%|�-X%��A���]��O6�)TkJ�:�dT�Go���QM��ŗÆ�8��ɠ�U��>��6��gs�좜j���Ֆ�¹��.ٙ��6&�]��d��A{��(�a��W���d��0P'�޴&�:��XΌ�ۦxU�r_�W\����Qۑ�����;�7�Js :"���y�י���1��e�~$5�k���@��]�3Hl���8�x�~��^�}�BN>r����.��Ɨ�@@�O[�Ҳl�o\�y]u!FH{p+�==�O���8������E�ۮz���	��O����:���[�2����;������7�����,}��y�~�poʺ�w�C�л�L��N���<�({�5ps��w*ꥨv��Q� ϩ�41�j�Ց���.�.�z��,�c��ې�	(G�F��11uo�"F�B�<\��LP����T�=��w�%���!��uϳ�/��D2v���d��yו�Cƅ�>��E�h��׵��R����V���̱�L��3j~���e'�S�J���1p¾��g��>B:�,���d	B� �b1��O9=�����81:�]���R<��vƌ�h�Iffa�.�N*�P�o:Ck�_Bt!דV��&Ol>��.S��<1��q������*]Wn�Vsy%����o �<��>��ƺ��ʬ�k�q��Y�WSBI�n:=5��I6�m��ȿ�;c6������ʥ��+K#<8t��*��Oߨ,r|s��F�Z��r�M�y�l�۸�W��z�>��y�᭞ǻ9e������W_{ s_��8���Y��2����_V"v_���ş���3�K���/\��t0q�W��T�^��1nks!ή�߯����)yI�m�
W1��ޥ���)p�����Ъa�]���*M�}y��1��nl������A��#��Erq��a������9쯱44��9�f����j�~��z9й9j�]�*<�g.dU���GT^�X�JJ���?'��H���3��S�����۰�8�3����4����,��ҫ#}���d%�ay�q ]�c�����]~�V�jx-J��Ţmg������|
DW���{���j�玕v��t�#����~2��.(��i鹰/NwvX��1nW?H/��{�@��d^H`U�?z��9�z�/mR�M-�x�>�I5�V���KU:�BB�aw���]W��:�m�{�VQ��c"���(��!���r��=����*s}��kxn\G+`���8����y�;B�Wo�e�ꍶ�a�W�	��b]Yzӕ �L�HWm�k����1��	�@�,�8��)<����ڸӼc*��}��8Ru��g�����+�ֲ�'x?.��N{ߧ��So�R�#�dH��5u�b�<�%V˄����*��ݘ��]0*73��}������-:a���]���]�0�Y�4�FŢ:����89��Wm`6*`�^�i�w3��4��)�VZ]ՌTb����q5w�z�{m~���S�&�ʺ�".��D�hE,�E�^���8�޳�;���HT�γ��������+���'�ݩղ���Yc�+]��T���I�&yor�����~�^��]��Ө[����/���~bH�/=�妡P.��(�8�55�Ink3y/7�hQ5}�\�U��3�1?�縂3�t�4ᭊ����5s�u�ݤo>?����q���0��uR��C��檬�Ѭ�OۇMFG�p;�z����}]3�%�І��x	�_fO�p�۵10�*�/3��	L�:�7
^��}��Ft�6��.�����C�g���T�;��vן���]�b��=�DKd�Cb�g�����P����G��,���IC������ d��/l0�iT+�\���,H��^pU�1��ms�]��.�kV́]�:Y�k���ưC�u�n�X.�m#͑�Ǉ�.���ѧ��z�nJ�RF��|339O��;�<�2 {yW�N��M�=\���HG�1�9�͝dW�J*}.�8GnީT�[��A0񩧱�[�y���l��i�ϴ���U������3U���!��ȹ�|��K����G��чkj�v��vce�;���gw6�1������壤L9 zL���^���������4�/7g�D��5����w-�mDY��6Dxm�Y�Z�~�LXS#��K�m�5(�TѺ�XN]�9v[j�;��ί�S}a!�����٩�R�N�d�e�=y��R�dU�^z�ԫ�Ϝ����L�g�iSܥP
Z�V��'�{����!��������_��ܻ�˔��%��8}y���G&D��2���&�{dLMQ^bۏf�&�w��D,�'�=#7`�xR�&l@�V���$	O�X��ǝQ��i�s��\������ ��	]��}�w���૝śp�pς�7���{����
�W[{��O��ѧ�a/�;��uM[q�V�y�����v7Nl�W EßZ�1��WU��i�<a�}�o�@���Y�>�@�>7�L�Skg>*��<��Sg�̝����k\�y���oF�����7���a��X���z�U�D2)2�]��vVQ��XF�ta�Æ�RG�WQ���ò� ��1h�\s�!��]^k��pa����v���+nN�C��dJ��ι??��_�����:��u
p�
g����iQgEv&�l)[��V%�Շ�ӱ^B=.w9���ʊ�C��V�~�Z={�X�l��k\ȇ�2�f��֓w=���=@�;��dÑ�|�ux�X���ok�;FZ{~N)J�����	�7��Nm�. z}��}��m�0�/���ގ�VN����>�����b���X0%4$\n����g>H��@w�V.������$����w�Џi�6^�FĔ-�ߺ����p���E$�����^��a����S��4v�!X��߭c���uc�/ޅN��b���N�������r^�N�A�x�y3��x�>ޕq�ޱ�:&�Q΁���U���Jn0�~?*� ���½#�_��q��6�)�3S�v�r�GJp��=~���Rh�7E�h�Y(�O�i��Hx�MD�3���텙��U�n��	���+G{5���Zr�ߙ3��w�ڿqW4��%#Mƪ5�?yRO�����_��n�ߛ��W����H4:�hj��7h��t셱'�%���pj72��2� V{c�CL�w�/i-��o�NC4	.�p��M��J����ǘ;wKN�q���� ��{��^���m��M���B^EA^:c"W �_b{R˾��Jo�絹͂��_׫=^=�{1	h/���~n�T\���b�;��W	d@7�B�.����売�!��;|-�ڏN��?e\�rR��*B)��`@��w�>J`/6�77{�/|| ck1�%®�҃&�H�}sq&���[T�Q���b�u�Gr�1�3�R�j�����N�Vt�;!�mn���ι��[G����D�Y!V׿W����H$���TUt�����~ɽ1p��x1N�t�g��Ǯ�aq|�Z�,&S�U��Dvfh�TY�7��6;�~�,luG���a�q�
C�
���e�A�O)���u��^dvPT��/������R��O���u��m��>��7kS��=�צ�=�Oz�j�d����]{ʮU�����5G��ї�i���GB����ds��&��V��O˱E�E��oy�5�~���ޛU"����{��hi��gn� K�����DaW�q'�	ԩ��³�Ut�]����c�v��9N��׶�f��}��������g\�{!�S�`�� 0�'�>C60�u�\�B��v�q�\�=��5����ۦ�S�6�(���a�3���>���ͼM�����N�rٲ�غ�1��}:�����t(b ������y�=O�Ҹ�9Y�j;�PƬ�;2X}�ܮ��o�A/c�8��XG����9��y�c�*+j�����!R�{���{�}֧%JQQՋb������c��|�-�c:�,�ş!�(��}9�$�꼟tt1`��v�{ԝQs^~���{�j�:�W�k{w)���e`��Z���hv�yo���E�E��߻��N�$Rb*K9�G���tM�l�f�(U+��
Sd���4�����=�u��!i�랙�WZ>���c7"��)�t5<|�
��rRIZ�N����]����~��m�u�wQ?�k,k������~�X�
�߳�,-��O#�7�}��e�h����y��Ѐ\(CzT����Ur���y[��y;�t�s�+ٔ�tg_�X�vლ"�G�'�6k���F�K��h�Wl�f�	Sr�Wy1J��(7���t�|��_�O�e���9e�zn
����A���_����M���N�cVܒ\�)�������s���t��<�����[��,�ٿ���{�g�*�ҳm=N3)W^Otu�=��7���D�;8&�6�:fF`'�ϯ��R�T��p:����
��OW���\�v5}0��Jlt�����Y|��)�Lt��_u�\�j�6��9��ٽV��ue�HL�E{�`/c5�N�ǲh�9�73-�8��<�ޝC�펮#,�w+�cz��S)ՖٽA�֫y��wXS�g��3jڵ���u1��7�F���
�U�t�0�ܔr�[ql�2Y���Ӛ)�F��S�r���s6ώ^7Ov��ꡡ�&s|�Ky%�Nc����u�çZ�=VW_/�R�+�J����G�:wZ����� �:��WC �2�3�ޚm�b�>��f �Bk�P�g`�l�/v�Z�n�`�����3�_��L��㞊*��S��j5m\h{u�+��v��O!:���B��y�Fv��E��s���M
��om �
]�&EyWwMI����Z���*���wU� d!����;��2�Ŵ�a{zDY��z��B�K��H�_*#�F�OG��j�ҕ�LZ�9>�y]D��N:y�`}R��VF�ye\U���-��tS�f�����(c#�ߔ����ϧ*�֧6��m��3�9K��B,-��ޖ�z��e\�	��"�w����w�U�`%2ެ��։���̰-B5�4�);T+�g�AȜi��]��ݕ�l��T{���+3;�N]�p/����� R��+Y�>���d����=Bc���ϫN,�\�':ݼ����xz��JG�����#��@9/�30&q��E7Rc�0|��ڌ���IM�����Lr�I��y���L2��-Py�
��Ez�Ĳ�a�v\���:;��y�lW�P��3�gE�Fֺ����h��srf���:*�Iv��z����sҟ=��+���2���2t�R�i�����S37V�C{.A��b"��\��>���
c5�+�q	��S��TMQ�h>]{��"s3z���0"�q{���ǀ��ʅ���+z��{Mq�����m����˜���뭽�z.�=�Ϲ���S��47���P����X�!�pfl{X��7��sYB���"-Ms:��<w�Q�h$O(t���3:��hK��X�R� �,�b��9��*�<���\ܖ��w�#���I���|���\���n�;���@����x�*�B.���A��D��i�w�ge=k1jYQ�������kcGk8)<���]Pv�ۇIXW�d���G 6V�kGw gh���g>8�QPc*˛{�ɝt����w��9z����}��/�^wcp��L"������*=7*ʥ`��^b�p�-��Δ�H�l='2�a�f�q���*3�ẳ7Of�� V�C N�;���7��oQ���#zFҵ7��z�9�*�w2���M�A�D	IZ�`������V�[w�R�d���tZ���O����}R-t�Z�M���W���WՂ�<��\�[+�G�7R9�ٛB���U�흝�)�Nv�T�w74b$J������9�j.�"�S3C���^i��0M���|͆Sr`�zG�}䢣|�d�.��]�&�=���[��MO��^���t]A�걖���X���
�*��a,�*b��じ����x�=`_]�^bG��U��Î��o,A`nh/_�B�Ŋ8�.f���-.�Xg&������)�
�>�h��,�F[�k-�����M���}u9�� vD��S�
A��0׆L^ê|у]�	���Ѽ���T<�����e@$g���w�E�^ʊ�k�fM>t2uZ��r�Uwad��&�	~�y���w��w����;�.㬧��x"S�����c����յ��/&'H�.�N4|`V�=�n�<O�ph��B���Y��S�`@əKtMC��ē��'��I;/oC�T0�����b�*�b�!K�0�ѷ
VT�ҥ�T�-�ag��)vA�?Ʈ!�6�z�GV��2�)��!�o3 ������	]�2�F�ՙ���M����1�[�k�JA�F��]P�U�Ђ�1�W�����d��q�b�z�����)'��V�!�VR�i��
+K׀C�n�����ܭ�Ò�l�Pj�,E�.��E�*�Qx/`���n��^�"�@��CYy�..�l$���lPL�]��r���o��Em>�{��o���0M�j���wM\���*�u8W�j"e� fIB>k�K�#��;N
�4��!�H����~�R�A���B�'�Lt��]躥�b��$瀞�
AN�"j�~�*q����q�����;�,ӻ��Ặ5��bE��U`�<�����`��X�tfM;�T�c+��_hB�7x���%����x�k�i e�����J��6�t���;.�{y@����uG�wܖx��Bk}��# x�ҙ�S����*ۨ	���A:�7A̓y�On^��������<	V��I���6�H���\�Ԣ�2�IN�(Ϝ������[�?�Į���%�:I��a�j��`^yS+~�Jj�ʋ�Y���u:i����_�"ok�|`:��lO7���F�}�<g�%��ɜ�#��>�2�	�Fa�ّ�Vkt7�;}�ϯ�En�[�C#h�;|�j���<�Y�����|�-]�cO��?��vm��>/�ơ^%�kW�w�w�TTjr��ꖼ��ʍB�j֣g���U~%f{�/ku�g���r
���iv��E���<T�c+�y_Z��F���jk�>�TV΁빍�� E��c����}~�)�������$�z=թ�^c����~5��_>���*8B'�p2yMMU�S6+�;+1��w�;�4�t���/U�ap��
X��f#[�d\�N��a^���e�w�{�ք�sD�Q{|l!�,��xm�U;�X9�WBm�4�m��M��������)�H���﮲��)��rK��X�@��\e[�9r|�L9=N�.�����7�jL�εGJ9R�|�푵�T�g�($��R{�ߍR
���Ď=�T�����&#�0��y-�>���N��J[ü��b�1`�6�|_�����S��Se��.p�uE�\g
s'�1��=ϕ�ݒ���1��"M�z��ˮf�z�1�]U -]"��6y��=�;.������GeBui��E�;� ߒӾ^^]Uk8q�B��3��y[*�ݍ��R���G-�$Ԇ#+E��Ue�?��~�{��p��7q�Q����D�@{��# I�OU�;�(�]y��Qܥ�a��p^��=E�����V
�k*���������6a�K��C�g�ǁY=^Ǡ��z�xz��͎ㆆ�$���p���}[.�0+*H��/��^FA8��pj������׵�5Jyz�)�?z�ϔ��:,{Pߤ�>���tDt)\�l�w���g��E�Oz�^��z�� �� ��R�wl����5/t��oR���<5�(P���:��3�`�&��o���X'���\w��al���u�3����|��&�@`�W��8�R�gL#:
Ӕh�5Sy.��"���a�2�Ռ��	�{��Rѯ����*��|yu�-N���gp���;I��wu��c:i����MS�=ͩ\��,�G�1�|��>SW]����t��_Z����� �f�?���-)�������ܹg�vfAvTj�~;F������U��,VM1Z�ާ�����5���x�A_����Տ�;k�o�~�ŕ�i���|z�^z�Ԫ.ݦ^�??�:bIW�/";o�����z
x��U�������2�]��{,ת �)5���i�������߯)�\㻒�?v5k嗖.�̮`$e��ތ�O�l����L���i^G��N�|6��'ǿ7�4��j}7ь*�� ++����Q�]e]�<>9��z��C#3/�߶b�/+���U��g��0x�E�����m�j^j��U4^;IY��َ�e��EB?*�N�_w���V�rVz7���������b1�M���
�F[�rg-�Z$;8���90�lz�璎SF�e���~ה�Ľu�4�(�2�li��z������m=�º����*�0����� ����V����l���]�'=팿W��yߢ� �go�Zƙ��sڝL�cw���I@U��3���w�$w!���>�K�b).~�ǵޏNj���ٱ !
Ffԥ�e��;���j��x�?b�@��ܢO����%8�ȳb�-~��s7V"��l:� Rz�^�ݡ��"��q>�r;V١�T7OEu
�L�pǙN�����%|�g�Ϯ�J��5)ܤ�؎֌��D-�tj*��;��Cʗ�o�7�����ZU�c���b�p�h�������:d�] IG��Uٕr���6��K�oQz�d�k7��쫯+��)�K���L��K4E-�K�\�J�cA*X����~���|�\}Cf^�J�^�2n򍩓��S�ޢ�NJ�S2�VD�� �A��.z`AI���دz�t�g��3�3.:(/�a�#��q����#ֲ��Z�)�+��J{^H�^��?a��J�����&�z�|.=r�%�}�4\���f��=�=��#�Vt�z�H~<����j��]vw�'~+?�4^EP5E��mJ�S���&5�2a�� �'��]�rF����	��s9����� �1����O��"ɕ��O'��U�^`�a�>xJ��'� G�+{P�v2�z�;[�����>5)��%��ז2�f�W�;ӵ]!���  mTJ;�ڀ#�6�|aix�,���dEK�P���Ǩ_+��I���m�ͮ �]{�[��ݒ
D�y�A�c�ֱ��v�w���iY����K}^1���e��Y~��V8:��+G�M��԰����Tm�[��-)��x�띭��TˑW{=ڲ:|C��6�([��b3��Ᵹ��n�Hz>຋����7�z�[hd��p����*�ǭR@,�G]�֕�^B{)��ڌ��-Jt�ʸ���5u���LyQ���2]�C���,fu�˴5����Ĺp�Z����s4m>]�����p8^��v�ayz�u(�2J�g;O|?ny�Os���4��;i�ӫuX�jj�;Ykq��5�
c����CFڱ�^V��O�u�|u�g?mY>����e5��X9$���H��;y�r�:�җ����w������p�Z��|�v��ᒷ��ǞB1�����Z�����Np�f7��=�q��;���%��a$ϹG`���z.�kT(|Ur~��[iȟ�}"�T;�o���nl�������7�3��Vޙx�5�3?</�
�����kC�W�k38��_��s��[j�G�vu���Ʈ`���,4����M��L��UH~��io�˹~\��Qm���?���W����PM�ҫ�Ë�!y�p3ł7�wZ�˽ji,�Z��ɪ-�,𩘌i�=�����{�[���u�Ӊ�Ե��5���{�'�����S�J�2���x\J*<����ݼqJ����i�\�z;0�
bV���d-{+��<j:OW��ZW�	�*�Y"�{����t� ��(�L���cG�qm������J5�6|��wC�W���Y�/��0eG�<;�����n�Z�y�;�3�.|qYh1+��[�d�>gyۛ��/\���U�>����uȶJ�|s�k��Ȭ�r!�i�F���x�G�Bɻ���b��T��5�5.�{+>Ɵ&ީ�t�B���#��DH���F�Kr"""a����d p�D���1��:1c�}���ȝ�3B[ӎ��,:酇�Wo�^ȹ8����=�FA�߬r��%�l����	?:pyОB��)��OZ��*������݃��R[��y"Y\��Ro;����	˿T���v�L���&�vO��o����[�,\l�m�+���
���̈S{q۰���� a�W3c�/+�.��z��~�Z6�۞�C|t�#�R�ׄ��W�1QK�Mpq�q	�H
�í��d�g�QOg�q۶~R��ED��;�y�1<��b�dY�c�W��^f%���[=��YV��Q�2��A��3uj�*�?�X�� g��6����3���+g�s��:b����R�QX��κ�Z��i�����0������EZ�t�u^�F!��z�*���=�Z]I��&�k��d�uݭ:S�W��S�����g_��i;y��y�Q��1\Wm�_��c��}�*P���e�Z��biǧ���~Iz�L�t-�Ž4�F���´��  W�3��\�E	ǉ\�f{��ٴ�m�a���䉮agv(\�H��I��UX�7nT�z:n�>�fx"�K�vX�lT�W���S嬭��;�Ԑ�qҕ����V:JE���*�!�k�b�Wwu�ݮG$���T�VF��Om��k������Yp*M�2 D�wv�;�����P�v��N!{�ަ�A�ACf�`��RaŸ���k'�'���*�dG�2D,���s?}>g��x��Nnx�g�3��YM՚�f�^�W1ЏQ���Ҫ���4}|}�-��7�jlO���Q��<���uX{�הXU�g�ܽ����~��m�.���z���ې���Z�g��i8ˬq}�x�Ѝ�n3�_���[��m�|�݃=�zL^ɚ�F���?6�><G�\�O���\C$u�z�͖��l˚9#U�c^���s�! �{�h�
��j,�A�Խ�������6d�D t�S��E�"�7�[��=Y՝��ׁ������&�u>5���	���'�r9y���|�?�
��n�gz�����_�#�D��@���'=�ĕ���{c����wqY�V%M�>�wxdX��'nޑћ ����%S�����{�h��ڭ<�#2u�x!��V�
٣m�)���E1��gk��q���(2�K[��ۉ������;�a�������YY=��y^�*@w�H�M������ �U��s��˓��7�W�ۜi�eY��#��Xul��p���;5e8��ͼ��̑�z�E��>t�j[���K�y���vΗZMѰ������t|��N�e̽��KlpwͰ���s���y�Hm�+�]�7M�s�Έ۔^�`tS�YX���F�a��Jă5�����:U���癫l;�)}82��F^�)Y�ǫV�g6�$�Kc}��g�D��h���o�퇋 !����b�/	�V��׎�:��V}��;��C�v0k���xuq���xo�*3�F�}����,���(.�M���1�E�����?"��VtҹQ�Y����t�N��V�"u܏\�-��a��G�u`�j�B�Y���gʗ bh
O��T��d��"I��Ƣ��x����
��6�czέ�vL����(_F�Y����q�U#���h)�"N� �@��J2���;��i��M{�p��{�o*Q�c�gU=���NP�k�{�»֛���
@���+ߩ{Ο��ť�����諸��*����p��0@�~��f{c2:�-η8��'���Sb*�Eu�1R�U�$�Yu�>La�K�ؼ��T<�f����C�j�S	�R��}��S�YׅA~�GWE���F�8���qy~��
�5�:���j��6m�2V�9\�m9S�2zH�^���=
7(	2�쒝���c�]mvNř�3�{���g�Ų�s��[k˫}	W�MwX[�e.��(��m�����%�Y^��~?����k!�F�V*ŁLEx���z���V�us;��Zc�^����<����\\p7�����F<W\*�k.J���B)���3��t�um,
T������6��������B��f��0�v��/��uB(�\+��;�Rɻ����oI�|f�� <�K�ѿI�.8�V�+��Vg�ރ~�[�/�~�³������^�����F�p��zfLRUP��l����C�ڔ��Jpް�~�t��߂ƃ?������rd24�,�*�+���%{���dQ�c�U���x�-L��9��8��{�V��4[���NM(�:�(��/�_�����ɢj��\�[�̚c���J���"l�E�����Zw�n^��=�E�X�(��>��9gr��G�\%������6��b�\6=[9�S��8H@��d��:蚍����/@]}��^��(�c��3!'��N魻J� ,|��Oz%n�L:�F~T�{�֮�z��Z��LZ���6���ww�ߒM�r�:��{�)�C�l��9މ#9Fëy�/�*Ŝ��GfqP[�����V՛)rޓĞF:LC���.J�]c8�=g� �Oի4����n/�2w�49h;*#�l�0����5'�UR�(k�DNO�ʀ����Ft� S���$���@T��sˬ[|̡�L�y�QK;F����N�c��V'�k��.���@�*�~�?GU��A�,�a��V��ML�K�,�ݮ|��x�-����>{hV_>@�s�#c��by�Vq<c�8M.M�u���#�O���N8��k�eI�c���S��b�U����ܓU'uݲ�2sq�.�X0ӣ�*��>SUM�φ�su����C*��N���<����o-�!5���y��Ox�ZĶ[�C]`���)xYa֌g7���㚺%�n2�JJtr�kZ�6��V�!4�^Z2��A������i\e;�ua5z�(�;]�H��/"��Q�Y ����f�P�K�����>�p��u��{��q=B<NU����^�ɼC�sN�3��)�h���wu5�}�>B^�؂GhG0ѱ�)\��a�Uվ�!}ԟq�y�ns�͏%v䮂�N��mg��K�;5��Ǵ�voKF��E4����8~��Z��=����ܣ
˜��K;[>��om�)�El��Q�v2�=��5���4�i�=�I��kv����>\�`�\\]��4e��ɛ��D�*��Z]�;(e�W�ա�r��@�D�-��9�AX6��}���oz�Ao�7)�[��oe�kr�;[RЬ��E�;� ��v���*{Ϫv���)}m!La�ʔ9=��n�+�AMˮGLط��3*��e�Fkq�����dk�w �=�0$����aG��w�KH�@X�:<9�+��@��Q�m���豠�v_+��{f�wK��o;�6��������r��=/=��*���u���`b�6H4�㭥�w�N��]a�����Ҿ����J��(/8E�5�vkp�c$V����Ygv1&vF7+��1���1�&�i�� 8y6��e��-�L�rB�E�m���u�2�mo�7W���Z��k�r���:�@�P`�fѮ_m�����i|�k^�Wm���J�c�r�j� l�s��*)+u�u��ӕ~[���Ţ�k_�|�}����t6��9V�@�Y|�Ҿ�Ғ&m����ڽ��e��΢�R`��wΠC�h�����q-��R�3q��GY����O��p��è蜝F�e�R���o��u*iM>S/7��G!56m�#��e��C�o8z�����E'N�ӌU���b�剷���\6�VJئ+��1Kq�2�G������)�{�#"�F�q���YE��ي�I$�V�I6�M��I&�i6�-&�I4�m��m��m��m��m��'�>ކ����&-!7������mhvo�\�twu�*R�𥤾�;h�������Λ�mgpx�2�4�i�48�B.A|Ms�ZRa�����DZ��eN\urH�S$VE�:�v�b5x_c|�ȕRjZK��:$���2(H0�����+�)�5b�m�m�:z�\���%��)���T�D����K�I ��[)Wo�J6&�`[��v����^�{)���͉_�}UU�Q˨%w��e�[C]����ưO;F(����}��A"��(Q��I4�m��-�0��]v���-�a+\�;r�#sAj�8�Ż��{�~��������F�_��4�Ntj;3qO�O.&�M)p$�M{�6=&������ߥ�Ò�GҘ���q�]u gy,l�n�:�o�8!l�m��`C��x8׬�Y��Fg/a�L��t$c��m���'�A��-Ư:g�P�p��W����D�M�F-�d_���t�mE����{߫����/���h&��7݅��b$<����Wc��\�,��H��f��Nϑ�Zz6�{/��`�I71o�����̬˓vz-�Cf/��?*�4�y����
۹�׸K|-j�؁�C��WȋG[C#\̙�������TG0�\��/|��]vZo��^��;��z��gXuĉ���d�zT.u�Uk��¥��.��B��5��551Ղ� ~�K�s��q[l����S�Q섯28�G��4	C�{�n��3���]Fļ��3��
��F��[�ד�h��	�f�ɭ��Q,j{�te���HƮ�zpH����T�W�~���f�$��xkp��}r:6~a��eG@(i�C!m/�/�z���y
�����]�M��u/%-+T��"4�r�[���v�p�1Ѱ�gt��;.��A٣v��7�zA8�Ј�=Q��;��*놺�H�!��J	���/��E�\�L\��c�܏$�B��r5�M��+�bTdY�7��uaxo�N;��[�C�&P�#>�z�<�Hs�jX��Ka�����B'�1��]"Ժ�S%I]O�}�ߖ�K����p7��=nZ��1&C��kW}obPGcۻ4
\^s
Գuֽ�	�b��G��܃�*����RIG������ߐ��r�oTq�E��E�u���j=����Vl��`:Y���������y�b��a�HH�]<"z��F�L�TN�W�ޕa��>�C.=�Kk	"}�KW�dL�oZ��yV�#B�T����2Y��ˌ���_S��(�o�Z�[0�������R���\���H�����Ǜ�<�/�^{;�o�}�A��=�g^��/ڨ����H*���8e�Jf����4�g�㾎7(�&`S�z:,Ff1�j��/J���Y[����Q�e0�/u��U�5(�9����H������z���#�E�^��g�%��	b���J�^�d��[(��2M�[��K���zh#{�}@)��_v�����,;�*�k��]mMH��U<Z�3Y@b+����w�8��$R^м���$�م�^_Y~�u��7���1l��ܓ����a��x3��ɧt����V�*���Ȟ��U��4�A�ֺh@�Igp
���yG�Fb��i��t�H9puonv�;�PB�/����zp�Fk�b��Lx[�������0��>����^�=�_��I��o7�	c^��T�W%�N�W�وd��%�j��|��^o@��S�Ó��Xc����ow�!�*� �2Ju7��Է���S�� �wƐO^yR7�{ܞ�v=3(��]�fv�f'�}�K����eN�LGV�#ju���V��fQ�������V-��/���rHy�Ъ��T�r�3�J��yw
���Ӌ��*�s�٘:]�)
O����כ`��5��'1�|��D�U��:�X딦~������z�C�%��M\��)ҙ��V�����p�z���g�4�Dogف��W+�NWn�{�!Q�z�=�lY���][��S�q5�F�j��Q����ڋ=�띧�|Gz���
��j�����k�9~g��˸Y]D�iпS���"��$�s^ej�7t����bwʮ���\��*�N#g�{+��%PY�n���ʩ��)�wL	����B1EQzj�� ��<I���|k��l+�`�Cr���pZ��z�tL�����V�
�}��A�@L�{���X(l<Ǘ��1z�����*��ï�b�Ц�Hgw�Ȍ����e�ǧO� e�)F�'�Ȓ)P�G���}��Y�͇��{���j��¨�sEeX�����<ˢ�u�쵮S0���/M�#w8��X%�9l���u�NW8�S<�G8%�A�Z�!B�ŽF�~�B��ذ�s�<���_2jc�FJ��t�<�8��:H~��S#�t�4��M�����H"�O�]ُT��܎v�bpp�TV<:J~��UfT�eS7Md�l�{��b�0��0K��=탚���fv��#�^����m�+�n&������
�SP�[Վw"Ap����D����Ե)�d��\��^`^������~{�r�J&Q�f)��|sd���t*�n�H��B��>�(�
��xHR������]O)�o�s�ʔﳍtj�S䣔��F=�g�f�a��I:�=ˣ�<sv�M�*��ۛW7�7ۥ�	Q���u�6F��� �@��\�^�P>������Dq'�޼l~���MW��c�)�q��ɱQ�~=��y9V�u�kέ�1A�<ϡ�{C^�ܹ{�V-�t��V	�9wSQ�6ǖ�ʾ��TOH�����z�<FTV]��=�d(���n�ga�f�Ad*v��`A܄�����=>��}=�׵�j'ƭ�%ד޻
d+�o�L^��fq�'��t�f��x��g���r�l9���hA4������z���q�ή��Ԩ{��	nӪ��q��k���n���#���ۜ(��mr/j+��-���Ro/��ᬓ��⭛0d��+�H5:+���TA�{��۫6+x�q��d��\��i$�m���ts���/{�.�;��r���J� �n�,���)��+��0$�ڠE.��ޚ��'�6�.���!�}�`��������zw/�8]MP�p�����[T�!� ��W6�hR6�y���	;�Lg���&:v�pU�!���GcSk��|B���;�P����k �T�@�̺#�FtW.)�Ij ��6��׷����W~���w�
�?N�E���`���P`��p#]߽3��{�чD���b��I(H}����{+N�:�|��DbI����/ĺT3�Y�w���v�e���]:�o	�V�Mc�OL��qt#zgi�n-k[�s6�W\bS���U{E�O�5����V�;�N`������rp�.��.���s��)�މɼ�TUHq8%�g&��H11ۇ=Gq�}0��D�N ��D�qT-���&l8�M�p�5Pn*�a3����6 M~Q�0�a~�,v��屼��xy-h {��qv.��D� �����/hzi�y�М�Uじ���Ւ[��c�&�o���m�����.������,�� �}ut�Q� ��Z.��?pذ��,��gaBQ�&+K���z@�7�S���2�Z0�!a���m��nU�F���e�5{}���M�btOQ���<��+�s�B-M���j){�4�+H���i֎'��B������J�=�]5����H�\��[���fxz��s=y�֌<7�F����ج���gf�_��=[���LV��\Lj�d?%W�y{�#���ps�~��ٚL�5o��:���p�ѻљ��:���ߎȒ���D����=��݄��ő��(�Mp��I���v�#���[#8w!�9�R���h/�zf�����sUķ�Q~��Ԗp�i%�a!N�f��_��_�B��9�m�>wj�[B�Y�f��}m�sg���,OT�!���z����<��Y��o���tR�l��x��o��?��ٟ����D��^-l����d���E�*�O����^��p��f_
���e:6�6+�G]��,=��LtX�~�<v~��z�]/�2�12�+�r;ݖ��pӞ��˹����b���c�nn��;rG��"�!��<���j��b*~}Gn��m�u�#`tL�������{O�I�61m�/�3ogq*�O��b;xw�{Ul����7��ܑuº�]�R�݊�[hR��&�U�f�7 �^�������`��,��_O�k6\^����wv���̧��n�[V��J��^D����Rj�e�� �M{��cb�����)��,0�8TW��s�M�&������=�.s��.�쬬��<1�nfvt*�2��t:#�V�\S湍 ����+ ��4�/�pm���g������\.,noR��<:s��!�_�c�{B���S���q��֎y��*䴐�z�~���I��h���Ư
N)�������}��7�P�g�o�;^آo5<{!��ֲ��O��<��W�r[�o�Qӵ��yK�z�ox-�����{Q���|��6�&^����f��s�n�v�����al�E�K�u�^,O���	+��k�d�R�{8u��K�!�}���#ٳw�&�d8���X��M���\�ά=�f��y�5j�U��V��S�C��Φ�z�'.iWs�^1�䭸���X�t��GE�`��������_a$[�IU^-�C�J� @��ݺE���=�P��3�xo�8F�{6�b��y=��2�qt�[�gP0����yV�[#/��rz;%�:o��x�Eu�-X����qw�Q�sh&K�i��ۮ�2�q���]����kL���v�c���WMS(N�����$)�+�]�X��Kk�#��ItR]s.��f�H���ǆ�����=f���B[�V���ccH�x�]3��0���������w�*��)v*Y��et�����5�鰉�w�����tE�o���c�'��[�A�-�Yi��hD�mm[�D�J��&^�nK�0 ٪f'��g^	H�ê�{sy�gSAPv�H��!v6`l��!*.4�����(d�7VLB߷m�O�:^��p��w�6�/"z�<ʃ�;��~����W9�{f�WZ���{��Hv%��K:Ong��+�X��4��u��p2IY+$E�	yl��9�������N����\������e|Y"O�� !���Zj}��S���Zy����:���O?5ܐ�³<A���?w��A�ꇲ�W��R\��w1@[�.�U�f���ږ��jD���W=j�wd��~�~�
��ԩn�1u��m���#�����MN2}4���JtϮ��Mh�#��k�I�~J��l�W�p���t\�;VxC��C�ll�J��"���熈�Fٰ�{�u(��{{�ܔ��[����=ی>ڕPNw��uz�f5c���ԟ�+`��ڥ�[⍫����"����c�R<��UVl��Ӗ\dt����ny��@�BJu�܌��-��<�w�~�����1F{/�Z�=C7�Y��r���a�]O�hG2\=Y�_i�?ӱ�~�(>P@��6\ȕlf����6���J�AT\�J'_L���]fM��qһ��]y��y�P`�P3r5��r�N`�6G���������4ڋ���G~L�����+k�Tm�G�̍p���K\@bcnYh�2p�/V�3RDК"��_�MX�vⓡ����"/��Y��0�onm��m�ƃ�T��'Lm�KM��l|VZٙ�j���}��u���vypK� ���*�[��Ÿg��Sٸ����)�p�-���������RTӓ�IO�J�4�:���op��p�~uP �	\[�����劇���S�l6y�F�[>�^�^��F����h.�`o*ؕ�f&w*��{�,S�(p���^J_SZ���Rl`=i<�Û�1X�yT�䝜��ѹ�����e.���������E�=����w4ḑ���k��YW�=h��z>����z����t�#ۍ��T<V����H�C�<�W���{����;��<kA���3�X����Y��V+����'�U $�*T�>�sʥ�X�ye<9�����V%��(�RR3���w��;F�v�Q�K�:�;�vvfQ���=]����>�[�89M���1~���綽�CM��G�<��ߦZ0j��@A5�hߛAn}vv|3fh�{�~� � 8���"r+ur�zQ�E����%s��9|�5�d����z5�k�嘫���웃X<l�,|��~�\!]�i����:���z�n���w�3zیfV#v"ˌ���~�ɣ	eaA�����UBs"�̽h	 5�vT�
�[�/Q�xX��8ؾ�5y#]�o[nm>�pp����oV��N�U�X�y��7Su�N�����ꕯ�s���ޅ�Ŗn�5�kI��Т�R�2��Wz:�7��]րͭ<so۩@
�	zr���snD(����96��y�b�jL�kT�h���j��F����/����V�K�g$N��d� 9sCC;,���W����/�D��܄�UI�E�Y*8���瞗R�n�b�������#ڎQ�� u-������S��{c�����]�wR+0U��)��:�O���Ƚ��Վ���� +G�,��u���j���Q.�FT^琢8�A��T�=Ƕ�:�Ʌ�MeE�Q=�G�����x����+����S�����l奔y%�P�B���w�` wj��M�?E�_niiB�������0[���P.�f�x����8g9���m��HSg���:��Uݫ�]�`���uہ�m��uz2���="V�^R�)�p8-����cΜ��A���k�*��3��Wb�Av�+@>�݂��X�����6V��W.fj����,�Pv3���en�HA�������8G-��u�k�+��4�l�Z���^�^Z�$������*�[&#"-�ߒ�jO�j~E.�m��w���t���F�(����+���\n�y�v�45�z���s�QZd�뿶ڂ��ON�1�r��l]nU檸�� ����v'�_;|P]H^r��$����WӏK���۾Q�Qsߺ��7]YE�LQ)�{.��"�r�nu.�)���cE�_^=���$]jxu2(4�MBp�C��{JɎ�Uun�fSK(�В�t��r��:p+]:����,�U���P:�I\)lE�ʻ�A�
�{V�-j�*�u�_��ۇ��+ՊӠ��⥷
�Ln�'I3zy��}&Ӓ�]����UW_��C�˽�\�ں�:�}�����7t[w:'�Nf�=�9M+6���M/����ָ�l�Iߜ�@<w}�Ԋ M�{�$�$��^����Zcs��JPuh�p�
N�Z�u�N��}�Q\%ژF�g9ӛZ�@.��+_Ľc��f��9x:�8�V�G�A�fh߾6������o���BBO0�g]����[-��k�-y�=��U_W�h��w���IR���괪D���t�O*1*P�ƍ�q��|!���w�y<�۟h����9����[N�0�Mm���r�Z_|>��Y�����/d�>,+r�Ǔݺ��3�i�z8�`{��]����]�O���V*U3�&w����P�)���:?o���|�B����x�w1&���=wVw*Sz�-��g[���$��֪�P�o�1��UUZKF%�]���#�������t��X ���!>`ϴHE�d|P��d3/��WZ�޾�$Ͷ7���"s/{w�u}_]�kc�@��
{m�{��nf�U��$��I��é�:o5�}�W�1�)�Z���u�
B|���ڲT��^nu��rs}�+$�=�]}�<�=t�"߻���I5�71��א[�e��U�a��W��C�>���������w]9�{P����
Oo~ޏg!�w_�wِ���u�.��{�Ih9�z�>ދ�x��w�5�oZa����u �r�@$� I1�@�'�/����?]��/��>߾�	դ܂���N��lu
����_7�O`{InVѸ�����mci�]���j���R?ud�&98-X��t��a�FAØ�'P�޽\#k���B�Xq��#y�va�fVe� �����G|���01�]�L���ʶN����[���G��$�o`.�C�t[엄5Y���Ѯιȩ��sx���o1��r���W�M\��Ez�p��=�ۣ (�}Ǡ,Ŋ�r�Op;�ݛm&�$9g%@Iד[�2��+�-H3Vi�Z��������\�A�O��܍���#b�;���b<��[Y��{|Ctkq(�	��r'��D�
$�J�d7�k\�u�Q�0ۮ�(�[�f]j0��ʊ�Q<����a�;rS�1!��΃��B0����K�����f��==�J5�ԗF���
�l��&s6��+UgX���9�Z��s�6��w�tmoe�6o��޻@�.��j����E�T	�VӨXp�X��Lgfl7��ݘ�u�%u�M�o�j�r��f���vw~])Ǻ�5t'�N���o����Q���-I�$�af��\� �vP��㻮ݍ	�R2S�p�W�
Z�.'����9��_R�]n�2��g{��`G�#x�P��2`����e5�f�Ќ����?�着���(��wq�g��mr.�v��͖	�)LL�w�Zlu��$,�r��c���v���J�PtZ)t
��r1rè.[*��W�U�LI�5���[ٖq�~L���^���l�u�!efn�7�Ό����̫�~94i��S� �G*�E��Bu�p�Ulɚ嶃��T��@��j��rϺ|z��aIM+��N�U��3D)\�����C���7��4V��'M�-���/���6�L����ҿPk����B�j$�"ykf�J틊�D�á!U��זs7NO���zW�6r��Mz��ھ�6���-O�'�Iy~@4�I�=ܶ�ʻ�;��!��ɸ�}��Ϣz��p>�uݗj\'9aY�Iߙ���v���ߨ��g����x�'�iފ�\���R�AY���`�ݵ�1%�u��f�r���C���kʏ TN���G����s]����3Z�u;l�T�"��3�	���}�z����/fS*4L *zˤ5������f������q~^} �2����\[ei�+�wc�?�)���w���NY�BVb�ʯI�ӽ��r��E�kLk�������,�Ƴ&' v���}cP�Y�s׶�9�K��qʌ��*���ͥ�
'�T�WB]v��V�ќ�"�\��#ۡ*Ѕ��^�����ͧQv��9�8ܺ篑�y��=��>�ZC7՛��w9��']�)�fK��VNE:ظ�R+�"��yq��[8���t����P�>=��4�a�y�z]���;*m�m!����/h�M��~�ߊEC���4�$\v�_�RlZ��t�����Rʓd�k�����T�����,���~��E^�\�.��Q�=����QSO$�dV�I�����t���xk[���3{�3^>������AJ��{v�j����*���9����_w����Ћ͘:�29c�Djc��F��z{a� ���e\wS��]!~�p'z6����'ڭYvc��!�<d;{�W��/Վ�bF��h�x�EN�3*yEg���`o}=�Xw� 
f�Ж9�2�c����'ӖoN�;���Vi�֮�z}�.�k�6��#yz@`��V��{�c���-�j���6mȴ�d�70�X�x�ߏi��x�1w�ǡ4���&���G�G��*�
�*��A�+�y\����l��,zø�)������v˴���{�m�LW�rnef+�0˻\��0�9��&�u���+��2ffwv}�py:��	۝��ch�k)�I�z�m��w��v��`�����z�Zބ(&v
��$a�\�S��;��Q��,�"����[彰��o�yAf5���̕��h[o���,=������,ǃu�ڋ.�T9:,Ǚ��]�gep�J�7��(��ȏbZ�@&�|�LJ�i6��n�[���g'���v9<���r.��>84�Oo�ֿ�K�=��x�~	^��F�+���*� ���	6)�ǻk'O!sΦd��v����8��97a3�hvm1���'%���l���⮀�<����7ݹ���� ���S�$��~�s_��)�oכ��+�~�]�g��7��XG�y�^z��~�&H��իF֔
]��5�Gfk�C�D��s��źw��|�n����7��<��ͻz���tq��+7�:#�)e���f�J�{���kc�3�T�ɹ�˦�Wê�T��έ�X*1a�&���?
�t���!5ʜ�����l,�E��ט�<!צ�9G��Y�S������1B���,G,���ho�������b�}�^#�w��Q�;Ɲcx=�Sw�Wō�U朸Eu��\{��W���X�O��H��}f8c�Z�Uxڱ4���.�m�ry��9>��K��'�	`���v�������t�w2n)��bMOP���K��a�[JşW1y��Ǒ�:c9�#�Ȟ��D)�µ�'�ދ}1��w4]��-���"��`]T�a���'�y^^��Uc�G��5�3�<DGhZ͕*@��%)���Xǹ�Q
��8l��FuGd�p�eoJA"��j7Ӵd�5�Ļ��P��O�o+p���Eou�-Gpb�8 ]�AwnAË3�o1��z/x�yu�r���'{���O)�Fh�����۝�8D��������5�~9�x����~;\y �]^,P�F}��)_*6g2=�zT7��N|4Ȧ�����GS.�M�=7+~��'scISn����>dճl�y&�1�ݑU]�=�Z��F�E�W��`ƺ��~ط�L�Bkz��b��K��y�R�K�E.�)̊�Z���W[�fB��y�ͨ�顉S����yǸg�$mM��&d�G�����_����>��|�u�/)��{��p���]8fKڌ�J��,��#�1oY��]j�&���q�늍M_����9�s�E`�6
�g��d����Zo�Wj�c���bC�蒲�kU�Y+f�i]Ǖβ#z=[X�F9�=Jj��瞼w"�P5�t��5���5�G�z�I��]�uE*�\�S�f�g]@`H� x�7�OSڰVW='���y���
mxߔUz�N�3{8�¸X�t6#����Ty܀��[劏���%���^�N�E�����;+yU�
]o���Wq�\z�CN�>�F�Y��
��""��ۺ$I�n]��Jʺ�t8�;�s�8wd��q��{��Zތ9��|	7�G��u3Ui��;�˚�܂J��u¡.�����dr��뺷��ϻ�)+����fRV>�5�$�St]gEAcs��#�^�k�ɒ�Z|�D����Q���'��wU��8��F5��`��dx��"�N�O�eZ��ܠ�v�
�h�o����s&s��
�vnC`��<�{���/'�{:���i��{th�]v?q���+y�c�Ӫ�����"�^pN�W"��DuC:o)��h�&${�1�0tr�9r�>�Ouܲ�U-����5�=#9�m	�Ȟ�:�T��Y��]���y��]���zdT���x��N��7=T=�ae1\d^��WmMM��ڹ�Fx��T��[�c%~q��~C�V�;�,�tު�0XUAԲ�����;�%+�b�q�s��n�;|�D����gn�iR J'�T��:�,����{��KϿ7����|�?��Ž,{��;���e��4�M2,�ԏZ�S�34{&F�T'��3�`V������Q�N�t�c=��0��G�OW����HJV}}X�H�Hf�w]�g�\X\eo��{��`N6=Ihι�t(�j�T���^�d���:�6����f�8�����Ap>�[�0������8�������I[e�W2^��.�}���{�柺d�r	��X�p��I�".�m�$�=�c}Z%ln��K�.���;�n�mkM�r�ztؙ�13� [gN���Z-W`Vv�u���8�V��M�����k��Gv�����lNx��1�s[X����οa���E��ri�؝D�cd����Wx�26%�P�(�P�E�U�/��M��2�2xԴ[.|��d��Azk�7�P`ɛ�7$���%��<�b{3��ݥ"&�q4�ʊ�}oĤ#��j�#����C��j2��#Մa�[������2��d�:�w�{����p���C�ET����ݟ�Ly�S��~��UpS�H�D8ޓՊ��pAN�QB�T�za����\�n��q�lw�"To��V�U|MD���P<��>��}V�)���=&w��cS{W�9�Lǒ��u�E�-�!_�Oeߥ�Dt<��W}���.��Q��������_����{��������y8Gx��oc��M�?z#�J9e��Ә�-?�1t�ꋶ�}�8�[�7�y�����~�ǡ���Xp�6�{�/�r9JU��5�7U\r��tf�ΛA���̘1{��f}�έ1��!��g"�\B���Tǹcto�tD�X��G}U�^�M>�[Fy�FT�Ru�e����^U�����j�;w+N,F�߳��=��V��bFB^�QFrةPE&���]���d�u�7��`0�<S��6[�����v��V�[�e,���f��I"7��īrmM���\щ�i$ۍ�e�,ymbū��k͗L�����ѡ�NY4x+����e=��Z������<���u����.��T����3���'��ܫ5��ô8d~�I�Q�e�J������Ƈ���m�U�n��E2,�O�l���i3��p!�-5���w7�ZT�.dK���א���C����=i/y^U�V�QZ��Q�.�OOr����*�e�;�^��4X7ь\j[�ݶ3W�Z��f��ה��Lo�/r<X��^8�iY=�&c�x$nM+f��ȕ'�Wd�T����l��wC�����{|�ϰ�s$�[�ԧS'˧�o�1k.D�����.6r��$wgC.�U�K~y~Jw�u	Z�81��G�4�����/�L�"��]^
�z���˽E���fa<d�|}������&_���$~�-�6<���UΜO
��g�m4���7�t �W��u�^5�S�ث�h���Ʃ��l�4/c'69�����#�k��ѵ�[����9� ��t*���v��#���
P�Z=A�z*�ˣs��e��������=]�%�,U��hD��߷8��%!]���5���j�ͷܩ����Tw�ڱ�O���tT��k�wE�F��d����V�iv��d}J�"9,�n�ٖ�S���ݺ��#)h�'���� �24+�X�c�ו:=�ى���,�p�;��Af&�q��@���eE���T����5��5w�ѯy�b��}n	ɽ��e�g���lG�ŝ�3��};:����)��F��]X^���f�$1S6���O(�風�	�noE׽;K��Ux?Ab����z�(鬢3FOq�4+���ʻ(ĩ���Sg:49�ŻӏҔzn(��O���V2>���;ѻz��K'���ْ���@�(��v�@�1��sr�f��OU{A�#:��R���Q�#��ɇ�e���A.Ovv�t%�"�X~��Iՙ�t��=fGqw�9��ڳ����6��W��᱕��Ĵ�~�8����B�Y��'���Ӆ��<io�u��V�=��߅#^������kh��ڹ�]���������66���9Ep�űRk^e�V�����#d��������{�;��qS�s��kӦ�T��i����i`utz4̍�p�4��t��b�&��fAN=S�T��rO�R���;W~eTړ���;�Yųz}����?tSBG	Xy^_�`ITY��P֩�K\[�q���6�f��x�a{�.�8�	�@5B�TW���*Y�A���Rt�*�n�� tuohI��o:�Bc��[���Z���@g��,�Q�vz,����~��K�,���e<}�Ԍ���oV��.
��]������~�����(�U�U'���|�/@�rDI�l
���-�"�g���b��xOM��z���(��W���i�����Q\�yٺp��>/�>� {���n���dn��`�f�%�\����ߗ賨Ie��t��������U�ya���ݛm7~�O=Fm��b���b�"����D�Җ���[���Tu�7�<�E心��K�6����-_o���<� ���54|��u&�#�ZUė:�4�W46���x��˶0����ôN����s��!ӱ�A�G��<��,�f�r��@��Mi��R�C�G�K�Z��%�s�rZ!���ǻ�w�]���಻���d���uw�wx�ǽ��,�K�禬�	.\������ ?@��<?m�bǫڟ�
?D�g-v�_-�z��\
B���}��2F6���k.�/f� �g�P�gyâ.��U��S��@�.��ϭhW��<2Qp�����y��0�)c�����c���,^v@�y�p�W��,$���P%&j��dץt����QQY�R2_���v���a��J�����]n�U����u2>Ʒ�e�Bx@�Qu�)|�����0�x�p��z�X�Q��z�eSZ�9�f�*�ݧ�nw+[OP}�xtz��-0L��϶M!v��q���S���p-�efd3q�z�o�8�ҫsهҸ�Kj��lW�N�tAP=��h�5���ݎ�Fj�ZJ��ډ݌^U*�t���P��w|�V��,�=#�l���Ԑ�B�g��3����mQ+q�BQ>'�8�����Ü
�����<U,�`##�ۻ�Y2�l&�GE#��۪�.�z|1��Y�Gd8b�8-��)���N����S�k]���u�w�(-c����p�P�<!��/w��8����o�.�,�q�Z{�GZC�v�'cw3δ�s���w�]�[��#�N��L)p��|/=Ѧ�F}�IKݐ��`㪽��^=���E��(�i�΀��V %�ٽ�����˕�录V�ý����y���v��վ������7Y%����oƧӃ�Q�3�ޱKI�S̜��s;oz|�E�ݩП�i*6T[�|�c���&߾��FU �����Ի��,�x�*sÏs�I�5���]	����=��g�S�]伦�Y���s���I�R2_%7=� +����/:-Ǌ�����/~�ϻZ�{��0U��M9Y�j��j�S�^�w�c&|��[��As�HiK��ǣ&���²7l��|�P����(�>�Y�X*{�Rp���>�B�,K�&�Q�ۜjݻ��hؚ�6�H������U��$:,O���2A�x]�����U��^¶j��W%muKq23S�~�y��F�Y:����V�coV �jG�)�����+��[ݥf�,g]������̮��$!�eT8b\6-R��iw]�WZ�W�K��Q����#k:�n<DիD�he�W+�>u�����,��9����P,7c��0���d���r�f�PL}U�+2ݹ��k;>ɵ�Q�ۆ �T�e�}N�n=���y�s�$3Oܺ�b�TE�Ұ(�f��`�r�c��UT����W�n�wi#_}Y���#ʪ���p��5�)aY1�͊PC��9��ۺ}���U�5�\���)�#�����1Q��h�wt�+�{j�N��Ke�T3\�ˀ����W��՘v0�~�.Gg*W\z�Nn��V:gr�r>n$r�*��{��ŵ��Et�.Q��>�W���F'.�����4e��<�Ϗ
���ufAå���X<)6���w`	�K�P�T�c-�����X����eRY�fҶ*�ep�]�{�Wbt�1z�����ƌQtV���dT���Q����������u6t3��7�X$'�ncS.����J��i��<;�0�<�\rd�tu
T�a����q�@幐�睊����S|�z$���䷻��:��^���	�G��Kou�5�*��*;����"fNB��N��.��p̝i<�����7k����������#1���k;�>!�uLX��n���-O�X���g5Ҧ�j�9b�wt2'�H/M;|���q�G�Obt��ܫ�)=V%���X��Z@L�m�5Ia�x�J�kv6t����P��A�l���;��x�&D+�q!t�+78q�7t--�,֗q��@Ry���c�Rϋ&�gz���`���b����5���QӜ�ۄ��ڥ]���h-��v*�Z�ש�wZ�&�ekCo8V�HO+�Ѳ-9]��<nM��WQշ>�1���B�;�XR=�E<��ٝG(�̽����J��q:�k
�������ݠ+%�㡝��ͺ ��p0R�����'��v����p�p;���g�vdZ��51�pԝ�)����<�Gs���^l��d��m$�I&�D��I��I6�m��i$�m��m�ڢX'{�z�.��(�����q�ho:<x	MMh�t��٧y״%4����vJ�t��!BBt�����j�<}0���:R/Ju��A[�Kc.�/M��D���"�Π�
���yd����Ya�`e��^Z��gH'���B����Ͼ���]���z�qv�����j��,�u+��y܃�w��Z�i���Vޙ�;�7��)��Z��\���+fWh�Q��Q_W:��OH��
G�e�&9M/���ꯏ+��z���;�﵇��#�"�y:A�M^�	.�lEIf�q����z���F�]x4�I6�I�ic�p�Ef���e��h4� `��}m�h5���� ���i�g��/���PS��x��Q+.����"Kr�i�e>=~ͳ��D߳�j��W� R����>V3���e��	*H�Y9�ƻ�L�:C�����$��/0F~��"˜�����;7u�[A��AH2���0�<��s��\_9#mX������M��CcY�>k���h�9W�c��4��g��.��h�mb�?e�h�?/z鳥�>��u���������\��b�&וξQU6QI��S��M[&ֶTp�2b�ܰ�
��Ѿ\Dd��
[H��k��}�]^ok�G��Y�����[N��Fǅ����*΃J*_��ب>"+ӱߓȧ��/�L2kȚ�]G�z�r��g� [��Z������&�����g��D>�$T3��� R�K�zG�)��ʴl����tfUP�\��	�פ�[��.��ET8���&�
o�*�P�ǐ�B�q�g/��e���ʺ�&4j��5W�3�5����@M�sQ {Ն��nxJ+��]��`�Ԃ���ͬމ�yw�ْ��l\U�Á۪��]r�JP;�|U�u�:�W<��i�0��QZz�������"������������8�ɡK�]�$��(���)�4oӒRE!�����n���VO<.څ�/�W3�����8�A�6�Fo�@z�u,��ʋ.Q.㧋�7p��/�׃%�y*&:^�n���`����p-�6��!�g��a�sFnQ33���`���5�g���^�'6�UXg;C �<A7����k}���G+����6��-���&��1I[1W��}�~>:77i9��5s�q(F��y)Q��w����nzົ�C_��*������|�D�^��vy��	U�N\/��*|g`L�!{��,ʛ����
\ިx�2�T�VhY-�UW�x�DD�C�e���Hz�A�r�T{��<f���z�w�������44����EvI�:kp?��=�8�z���A3C���D��W��y��3+E�W�鵿�w����a%�z�-s��r�	�ϩ#Q*c����zH�{TŴ�ɳ��w�׀����'�)ԥ/w����V<G[:��+=��U�9N��Pș�b�=�^����УY����V��m:��3���4}�\��=+���Y�����;r���=>��/�Y1o��Z#%dɲ&��a�����䊥�Xԕ�*������Wf��/'R��]⮭y)SS+J���F��ݙ[+,N�N���z�C.)-|�U�h!ډ�o氼�ݰMCm�XVa(Ω��=��=2^for���h3<�?�C�W��C-�dY��L���9�8\�������1����dYw�<��]ϡxo��x�%�P®�20�b��:�͵�OЩ��<"�����Q�A��hb���V�I?�S�7���=lT&��&��\�-��s���*
�����6�\�v�~�u񨟷��!���z�_������tOsͳ�+��p[33=�|r:��sWE��,�T|��o����^W�����w`l��<��{wd1�����'Ց�Ƽ��N�^�^O����^��'^R��N��a��ދF'0���w7�uϺ��j���D����y;��g�O�1<w���}��ߺ�Dr^�|+\��^�!|��woj�{o��x5]»�w+�_`#��TD@��i�k���#�\���8��~�:�,}]S}�z�H������c�wSE*U����+��D� �s/�|G�J�e��+��6j�A���33��Wx�c˭�#���8֍�g�ߖ[���v��������9������=�s�-��ZPq>W�	O.�����Cqd|��L��Q�,�^����ʸ�DƉ�znd{&!'$���NJ��1\���Xtl��nv��u��b����0[oR`;y)��[���.C������1q�G_�}��վ�)A��0J^ӭ7��$���c�3ݎo#�r|�p�c����s�ƸKC�Jm�R���t�S�fS��~�B�����R,�U�x��h߷�T��#�<��ң��/"hS�2B}̕��g@�c�->�7b��k��s�wP�]��|\�H�>j��6�<�&l��&&v��e���i��JϬ�G.��\�1�9i�UK��3���eJ�'�2��Q@&@�l*tG;�٠�N��b+�U�4�$��'w�T���..��Ԧ�mQ��﹗XM����s�+;��i��÷�4��灧UM�Vz�����O�Z�~-ɉǳ(��7w�5ܪh|y�4���I˺�Ч��f�1q:�iS��o11��:9����(j�]m1x�ycd\6�9�V4�_��v2]~���
=�κ�^
@B�Țز�{7U���G�j�0��}���qؒ&ed�Z�ߴ�+ތ�o�Cv*'�yN��*���C�v�gFd=�T�O��@�A�"��Cj�g�[PF���X�s�I�h8:�-8n�l�}�/I��P�3xh��\*l�c���r�ĥhZ�h�b��i�1Ԯ��v���\��b�O�j���\�d�ÿu.Fr6�I$�m���藹�:�+tf���7%	�xjj���t�򒳸���6����ߥ����Ym�J�8�R�X �p�F���t��ۿD����;f'O.�K�U��AeL;�3&�Q�~���H�j��^���~���ɸ��첛��a��8�[�龡%�+�|��K��qnf�g�����3i�c��s;�CZ6~�>�_�K.�j��N�U��*2�'�ɼӑm)�����g���BsT��6F���Y��T��2}s�~��vw]6+A�#��5}⑉g`�������* u �R~�쫾�{�×��OWN/�\�C�2um���qy�c ���;��g��2�_8�=\����
�;�f�6ۈ?��i��㫻ѽq�Q-�R�O
����~{�C�oS�%zq�������F�U�I��b�O���I�Ø��x���0���,�����[ڏ�_�:���/������/����}��\�1����=��\J�=2�y\�5C�1Z�S nZY1��x'u��7�����f��N�+,NOW��XO��0������ �k5����}��Ք�]Q7�+���7��nP����\mlneM�0)�KjAێ^ȜK�}V;4�W!/YK��\s^Y�"|ۣ�р��%�T3y���)v:��tg��-�ƗZ͜t�4����|7'H�/`�j�R�G�j˴�4�ك����2�U��<<v�(mݩb��u��ގ>K�:�m���޽���n%�ny�׶�MlZ�����Cc�� �F`�L����lv>�ǹ�Z��~>��%eEc��Aٱu�a�j|�]R��)�1�=S/�L���O�VJ�Sh�q�X!��9�/�J����]	���|O(���Q�S�����Q��ţ<�܉�Ti����Y����_v���tx	��U��=�q_UN��Z�Q+�;'�fJ��9v��bm�Ԗ݁�]�u ��<��zyߝn|�+��tK�p3	_�O�K����c��-�Z��4Q���X�N��F�~�a�;D2�N���^)�5e���'Q�3��%���C�ed�/�q�9��F��6�g���.m��&�
�wz�,���UTY���:�^�>�^j��Ğ%�[�l����T���s&^��P��{�<�r����ϥ�7�EUդ��e
~�z��A��c��:\e0�	�8���>͸Fh�>yÍ>��y.5͋G�kGvO��*��C��V��J����W�~#�b��RZK�hݚ��ם�Ǡ5Q�+g��'�;�2J�+w��R�>�����J�N&J'I]8S�Y�ue�0Ԕ
�m�Nw;@9�q�뵋�>h]�R��NY�Ozj�V�'��걔��;gN�/��{C��+��~'�.��+X3
�½[�c�f���p2�K�;�͞�txZ�)�
ǴMdJ��/ޖ,��QǻPƙد7sy�g�{]R�K�aNT���i�.KR��+��!��������v�x;��h���������k�3�g�l�yt��S<{Jί�pU��c�I�ٯw��W��oȟc�;���G_V9���<'	���U����~�hb���.Hc�!��V_��R#n��(�y$���"��hy��)�Q�k�`J�9۔u� �㦽\[�9�V�[4%x��SW+�?D����BJګcMS��# ������f;����B�z ��fN�,eQ<g��uo$�wu�k�Q�򭮛�Pa��R>w��;~�X˻n���n�<kflYp����P���6�rv�m�P���J5E�mdZ
8���<�|ES���>9L��TFGLM��l/�jv˙�vA��L5ʿ@4ӕ��䝭`��*Y��z���0n����w-�"���չu5��q��F��y]s�N�͝��u&���>�y��I�:�}6�kF� ���h��Mt�3�Ԭ�T�gV�{���NJ]k��S������J��Mh����H�4NWS�x�k�������Dhf�Rn�=t�ht�.9G�}��#;o!��l�K���=q������EP��բ�l���G���{۶;��Du<&I��L����P�5����Kǀ4}���}B������P�����@�*S�	>�V��iwWw^Ř��0<t��4=5ybn=J&�s9�F�C����ۺH}�g:�����B����/_|S�^��*udd������=S;���V	�k̃�kE�~H�U��g�������Z7]����'��w�(��:�S&��ժg�O#���ȸ�㼫�hWm���5�s��JN�����v��Q���W
��Y����0���,GvwO��D,�u��T���0��s��h�w��X|���=�YR�2	�k�_�%]U.����V>QP�Ѽq�˛�hR��p����9��}���UF��,^��J/�%�9ASP
��ʽ9��'n�c���F�K�D\��.�I_�Z��oH�ui�y8�#<|8L�	MX�FT��ef�Ǒ8��f��f�H����m]�(㋮�ӯa�H��W|4���v�&��İ˫N�Un{��̡YP��/٢���'�56?��[�_V�Cy�t��7�N��(w�=2����9%�T�3�@��Ss{V�N��s"����=廬�;"�3�n�sE���uY���v�m��i%��voeo.1�l�^��>U�R��j�pj`��ħuZ�%�U�tM�Gx��;j�t���
_k~�3�Ӄ��{O������+���G���,s���ϷN� �� ��Y�m��w��Mn�l�h^8�}]�ciWmV+��C�Q�s�� )�E���N��Wk��|�U�%��R�s�k�=叩T��%�b����k:�Py��^���p��6>�"0B���G��;�Le�땧#�n�\�r����۞�-s �X�����R68yzƗx���֋�y��p�*p��<��������]��ݽ����חg��Vh4�G{�{&���(�'<� ���uːw]��W����q�v�F,��BO��|��'�a_*|W�P~jES�(��p�a�8qK���Ow���q��g�]t�Z���k7c���$�x9���JTo7�f(<�Ef�����mVɴXۼ�t���u<�O��ܻ�_��Ag=�+^���[\���S���Qq9�
��%5]�:����vHs9��K܊�� .�8���.���f�G�n'��#K�*�ԏZ�}�5��??$���9�z`�V��	�-��F�_V�B;�¬J�ۼ����t�RI�)`��X��<o>�ku��lZ��1I\;�)V��*3���Z���ZJ� �x�����E�7cu�*��CF�.w:�b8�V5]��nsɨ�k���^���M)�+��
B�G��<��[Ocjۼ��[�߯(�q�g�a�.w(�b��V�����Wx���ײ�!nӿ���,���.*�p<���~6�Q��׬�{�x��^�fJ�7�j�4#�A�*ĸ�YG.��[�x'j%�bg�tǤ���y��G?Q���^¤�y�bܰc�G��enS�'0�����<wY���&��O3X5�Z;  S�"� Ef�Y������"d":��3���K�EwK���X���*��L��%SPj��՗X�?/yWw��1��˜�뇶��3��9�_Q�����^.a6��r�[�I�M~uas"H�^�^��ȓ|W�y{,�9Ǐt����JqRw&wl.���lr�W`I��9z���E�;�x�48\����
��lx�7�-1�n��)v�C�k.����L���!#'��P����eI@?�s�ݵ�~�3�?�OM��T��OL�<�o{G�P�;�բz-��P�kv]�D�\�;l�Q�GTh��i��-^�7x�Wv�]LU��T[+_el�C��~�(��q8d&����X�7֧�.h\-�_�u��C�SF.u��A:=��O^Lۋ�]�62/��j-r���J��w,��7�w���q�h9�u<c+v����h�Xj�_S(7Z��9����g1��崥��s�t3��;W26�P�(��C�~|N��H���ֱ�45�]&�)��/�B�f��s�Ws����3K�j����-nA��X�x�vؓL#sm&z�v��]��)y܁�lǛUR��w��Ͳ�d�Yݬ���K��t��<('8G�Fu����f,1^�:��JXy9�r�a�1�����#ى�ٰLý�-6e4Hy��}��sS�iGC.�G�YAa|�ϊo���VԄ�؋䶰qA�i㫽�Z6�@.��̈́�\�r���Avu=���	]�%�?!�H����r�j��:+.���܍����ʎ�m+�l7F�۵�.U�WY��ih��.,u�חH��{(�W>��맽t�jA�-+�1\����R����B����[�) 7�2���f����=ǟ&��
�D�q���7�[)���m�N��s�[�DA���<�����Ô���dm����,vkD�1�Ǿ���.;��ن.����s9�+�]`��3]�1.�1\��.��h���:vv6�]2޵��B������`������x�QSozl�ʛS��wW@���K��)�=�Cy���V�v!Ơ(ξ���ƶ\�|.L%ܣ������\����y�y��Ю��ZY3��Ј9��(�`���m]-l#�T�1%�v83��*��XR4]��/��T~��-��]v�咰�g�7�Etރ5���!����$L�-�3Q�'�#2ax��zz��2D�L�8����Er�m;�z˼��N�V���:p+q�fJ#����FV�	�[[;���d��K�(Wɕ����[�N�r��LJ�V�W�V�'j蝬�k�]�$��vL�6=���g�P�x�0os��S|)�yˌKrӬ"�m�x�>�eE�km��9W3f��|%[��@J��Ӿ�	{�vs�,ܮ�Y��t��HU�vM5��ժ"�@�Co�T�۷I���@J����+`?5ȧ[��L�2u�
�se� �f�UpX�8x���D��W��]��\���I�b�jIH�x���U�]o�]'�݈^C�#~�S����y��ά�'�xS\��n�ӂ���dvR��&�越��7�R^ 5L����x����"[����4�]s�^XRȔsq�]E!ۊ�]�h��gf:�[Բ�6ȗD�%K%5D�@����֊5n�-��lk�A��i>�os5��ud��e)�;��0)��u^#��vo=s��(q��:�tN�5Ʀ�U�������]yA��B��Wtx*d������X�-�4�l�Y�}M]�v2��ӊѸ6�CKf�������i��g����uz��;�|���×�`U:��q[e�e�;n�Ӥ$�.+��>�����7��{b����%���@>\ϔYC�#����6�2f��2�xf���1��q���'�_g\'|��Ǹ3�;��N�U8 ��Ҩ.���~=n�UϺ�^�J,�c��B�@�R}Grk/c��3�J��
t�I�j�<\�y^�1A��=[^�3w=�$�@�4����2}rOTz�y�Y�:�3=����o8����ooy�hX�p�Y1�w[��~���3zj���>Hp�TVh�"U(�����=+�@|���w���3��̖?Pmċ��sϳ���ׅY�x�	�Xz4�����]�k�=��-��7�FR�9uJ�5c(�E�6I{0�FJY�%N͞Gn�uu:E����\:��'V�ۜ�|3+7���^�뤶i��mw��Xo��6ޟm1+۔ft����k�^��ٽ�䤞{�%�|\)~��J�<+VVQΥɎ��9l�c����y��&<n�X�����$
��)��KY�Z`���!ݧ*j'���r�`c('T�n�GqtX�f�j�����Ta�����s�[x�X��H�f�r�+/5�`(lʹ�j]|�,PC+yH�΁r�Q�s0P��z]=y��9n���F)p�S�3�<�a�70�};.������5���UW��߯p�u���^�1�3�r�[�[��Q�O���sj���eJ�P�a<�̏{��
��8�M��\���<3�u��MڃT����\�����(H�vl]D�H��7k�=�7���U��n����L�'ޮ��mN\u.�fj�j�,)UՓ�y_YlM��>�S��ݍb�]N���t�J�	%������Pg 5�ћc��t�R�݊���� ��޷y����C���P�z��jCB󷾳TcpU��d��B?�xb>��^�y��(Ҥ�<�fn�qK�nt)��;�I���i�E{����L)�V����zF�S^Ε��B����nK�S8X��^z���<�۔�i�Tv�ɨ8���>��UW���	�`Ⴡ�#�ߧ�E��1<�u�5Xn����`/����h�^��15�:�00Y�;9w�>���ȁ5���מ�k��=�P�	W�%��?-��7�"�P.�s�*t3#�mO�C*Ba�fo�t�#��
Ȗ��|7q�E��s�t�}lB�lշC7`�t�[��v�q�Љ�v}�M�NRٛ��Iq��|�㖉�Mb���dukP�[�o^@��]���i�X��p��*���t�7���m��m���N:�geܐ��s:����w}�|�:��}� z��v����Y�dSI�}uy��W������|1q3��Q�[/��VW8��^��Mo����Pvo���Կ�/��6ev��3K��uu>2��[!�I����̝^�`895^�"7��^�JxPl���S${�״�w� ,���J�ٳ5+=S�Ѿ����R��@}�LK��U�aNo�����F(�T$~��7�XV�샴���\q��U�#�a˂�Aꑾ��D�u>Kw�zM��f�	���Z��M�N�1��Z>�ʸ�X���~��%�����y��Lfa��k&L�bm�z�T�ϝo�eyA�8���ᦚ��3�;GMx�xI���` ���ڑ^�J�P}x�}���X��^�=�P��l<�Bٿv{z2I.	;� ۆ��x��'=����ɇ�̨�~�W�;��}]���sC3]�<��jjA�#��&s�(,�WBgJ�,�p�^��4���{=�-ع�-�u����jUy'�!ub!8�k3����6�b�����ŭٓ�:N�R�w�<��+L���#"�呲�O�%��Gs��:=@��y�[rk�ֹ���BA����`
��<��ʰ�oWB7O�(IZ���t4wY�*EBs5��-],�7���W�r*֑�/[��4f5ݙ�*�gH�E7��V��_N�=<<�
�7��{U��}38	�Ż�ok��=,s��p�ϕFsA�u���#3:�3�>
t��W	���]؀�tI����o�&���1�<��//�
�^[&s��+�p�1/\>Oo��O��f����y_^X�ۅ�7��4��=g{�
�G@���'[w��_���o5�n��[t������v���<�:�n3#�gh���7�p�Yk���dj+%�EZ��s�o��
g�]���V��_���3^EKF�+Cj��{y��o�5.���tKԘ$rq��~���n.�؞�W��'\k�m�Gd��Y+�ia�5sP�����o�x�!=CG�}��S�����wP{<���짆�"y|2�X�V��Q��WMo�9;����Z:`��P�(F�
0%�W�s
3{��&T�z	f��ZVD��ף�����0� {��Ϻ�2-y�ĺ��_����c�QiǶ)jw��g���zJ��(�[1��O4+��'���\�����k�0���V�IZ��!f�\�;kUA(/+�]h���QqZ�*��=G���S|��ѐb4}u���֌̭�9��ԭ�����M4����6o
#]!4n�Z��Ҕ�AI.����@�{5�T�MSz���є�Q��>����S���1gi=ds}����C��2��%N�c�.@����xs0������p�>�c߱�t��k���K���c
��k�};Gm�f���ܹ,X���N(�@�R�5ڲ�/t
���f���'sK���V�l]����;���j�R�qT�$;}��uO��_��	����]��A���<G��g����g�x1��DqfW�ɸ�-��k����|��s|�̽�(��Ȫ����-�
��
�8�]���J{��d5�E`����ʌ���V@��̫xx�.�G�{EŷlҌ�����%^7ۑ�훵ϥ4.��g��x7�ӣ�f�g���*�}�j�M--G<�Nmb,V�f��d5w����yW��/���UO#?���G��X="skoc�2�����XW�R�k�v�`}S�(s�M�g�-9�V�L���
��g${�i1�ά5�u^J�� �2�J��;j�9������Z��L���k�]NRś��o�<�^�(s�)��ʁ)k&�\�yTd�;�8p�#���5��=u�0���)u��tZ��Q|�t�
�zO�u�7����\�n��~�^�}������)m�iw7ֻ��1�j�Keυ�5���ڹ��Ʒf�w+�]�ǹA��,�p�B�q9�'i�(�٭Zs����Y�G�\X�;v��d���k�g��1�E7����l����\teu���O �>��>.�ܣ�ov�:�����[���������Q���0���yh�׽m��_�.���������k��ttu�\�Y1q�/�K��a�<t�����^�N%���=��WF.�T���kzeh^�aMK��1'
��5O����t�j>U�Z��Y"���ʲ�w����I�+�7��<e�>���ˎ\��o�\`�ڬ��^���T�b\�f�)N.�r������#Ҷ�|�U�����7�����̢���U`_M��oa����AA�ӛ�&Uf���hW��jT�5}���S��t�>W<)!�4��ʤM8�C��<�`De߱��7r�!ݦ')�
�̇�����¬t��/��)�j�$�+��=�����2y_��:��;��yŞ���\�n.���u��ͯn���r��a7oy����bWt�J*W����h��V�_��v�It8-���Ĥ(˩>l@�ST�\���MG+��J����\�*w�v�s�ޥ��2"O���S�3;V�&4�=.cz�cN"���"�<
�;��C�i�G�E�S��/,��\���ޮ��Ս��z�g ���EjܻH�߶B{ie�gr�S;�*]�Ѻ�SUܶ6����m��mL��]cjd��W��-""�m���-ح�۽ �ڋ�ʷUU=��%ZVyO{F.�}繺3�mҍ�4��\����ȡ<�U����#���_��O��\��g�<W)�rܗt���s[t�j�-V�*[�-�}��X��'0���-c��ͩ�C��Ⱥ���=G�����ղy튕s�cP�M��G}p��q�E�*�T�-][P��:Y6�v(�#A�8���&*d��u��^ʆ,�}��Ļ��5�$���R������k���f�Pvx�G�_�ڱ���x��&�2W���f�����<1�^�⪨��=s�Q�]���y$��D{�9�]Ӟs�u��B��-8_޵k��\}���"��*
_2.X�u("�S�q��zv�:�|�%�<���3�A8W����Cկʐ�_������_~�ִ��[5��Η�T�N�:�J�	p@>��3��	��d+�⇩�^W����x�R�����.�
����.�DOk����f����M?S��>8h6�c��*Gy�>���6��><Ѿ^�1<��=]C��ފpS�1�M������a�m`���X(T�S�r�Fُc�h\��2X�1�]˗�j�nj��3���o�=������HnN�$�΃B}Wi�: ��p�\M|�U�cu�e�fI۔��|`y3f$�-��2+E��ǽ\K�b�T\l-���
M�w��Gq]��5)��doX����1C��p*�N��w�;�*�J�}�L���]�w=Y,*�l:kc8'e]���u�o,�G��U���nj��bʟH���#�UJj��7�XQ�|uW��4ӡ�\`�17'�=���>s}9����m��,!8霩�g�ũ�F\78�~'��>9s�+�~���xEQ��&C�����a�9也u8�j�2\
��9JλG�&��L�P�_�f�<*����=��_a�?T�gB�ͱ��.n9�g�U��jw-I}�
���I��B��M�0��Yǃ}��\n9,�`gZ�ə�6�j���X��/�r�~���Cg�
F��
�Z7����˄x��<��:v+=k��^;����8�j"�"��ҧ�������I���$@�tV��C.�Z��22\�w��5h�%̛�s��{�_:FUʁ=`�c7���at�Wc�:���t�\A�~s�����a�N��Z�TɆ��}�7��=nܳҰ���O$(%ث_
u��8�{�;�k7^�CF�� #��`�T(=�u(�b�{{����T��B��L��a�
`\�S���`��.��>7�Zy�<��7���9���;F���#a_��گ8D	CoJ�d�~�x�=��&���R�w��5����::|��K��<�������O2�9��H�s��J��>�_r1��U~��{���m��ڮ��� �x9ۦ�h�9�&���ȃ�:���D�Q�*�A��뜎�۲�+�z� l��l����&M���w)�_wފ��v��n���iQF�>3yy]����)�O��ց��'�'��f=�0C�B��wqן�s|���/8m5�_��g�����Uۯ~�~U0/G�F7��߆����b���s��7��4ߺ�b�8�/ފ��k�t���`�қX����þ��C��z�:[�s����CEFR����Wy�:W���V�#���vJ���S�:�P^ܧ���m�U�%���e�	i}�|^���s����㳣�:'��9�W���>�Q]�b����+e�7j=����t�J}�T42�xU�ĮtM��66cH{��3l�ޅ§�	,�M�![8���%���(yh�O;3g������X�Z�\�J^�T���[��WvZ�P9Bx8��/��|�I�ͱh��T:�}�)q%�D�pmv�}��%��i�9��]��xi�e�W`_E����jȬ����b���]�������	��b�:��=�72t�Ŕ�$�L��v[��o�m���JL&�P�{�s�9��+����[�' ���05ut��cQc0�8������9rĿ��t1{4�L��6���+��j�{���O)������gy�#�χq��qV1މ��Y��{B�)�sv_<��^h:�)��Q���*�Y�f\xM�rp���
�>k��3�����+к�3���/Tj��&�I�ke�7�<�r��2뺏x��b@��V���y��u��LqfXr>U��]����Av���*�.vl��'��n�&`�.K�T�b'���ˮ�|�nMf��G��W��ԫ?t�;Q�Hf�~ET~�$N9*�L;�|�eY�w����7���֭��e,��E8�\���kV���<0]�-Q�L���E�>F���+�/�]��:��A�cڱ���*Ƈ��>NCż%O����N�u��>1u�����]��T����QҠ㉪eR���6~���=>��^�e(�0��]�4�m����Ϯ +�_�a�P~�B�mԮ�/%t�wN`j��1#+v<�c��w"������9θ�l˧Q&e�wCrsj���ƕнٸ$��̆m��C�=����Vg���й����u�3����1��:d��(��(� ������g �9��;O�N��;gQT,��2� i}'��UsA�.�΂��!�$;�#����an#�t�)�Ũ9K�;��%府�i��2�҇��<��.��*�T��ǻ��Ԙ��(��[�we]"��]�e�6�s��o.�����~η�`�֭�i��E7�+z�j��]Ɔ�W�ԲI��n$o5��"��:�Y���]��M����37�k�����S��e��A�Ȉ�z��:�`G���gN�k�ا��&�@Euߕ����+�K
�K��^U���7�Ǯ��������o^,9:68p/j�-6�C]�����m&�*�t���3z�L�����hmL�
E��W�[��V�Sf��Rs���gu(�ϥ�㉊k�:9�3P��n�akK��Ô�gK�t ����������x��]�ķɧȻ�":�L��o_TV��aL��q�Ԇ�����y�.�.��&J�A�g��\��n^��j��˕;:�c-��<Bo�;���;`	_7v4��A�ؚ\��r뽬���l�(����pf���������훸Vr̳�� ��{:-����vl���z�dc�Y�h�Yc(�Iٗz���@{��`�Ym�Y�e���m��(i�+���\;+Ƣ���uso��X�8�}�g�
�|��f
��R7 ��2��R�^NO�S���kb�KU���{�\;��/B�淖�R�"i2�&��ڨ�eN����J�vâ��f��n�Q���|�ǚ��o��{��mm����(A}�mF�x�-���{XӾ,��	kF-�`�.�Q�o��[k����cQ]@ӷH^Qs�Ju%����WL;��љ��Y
�*��Û��MZk9Qp�Ǽ�ޡ�Y� �z^������N���TV�V��i	v�*4)� ��>M鮬��� [y��;rNX�՘;7���S��	�%�P����YF��[6��+�.Z�)����C�y%PU�6�1rS"�Ŋ6�K�v3[Q��i�a�i�ԇo.�v�x��q�l6��ނԢ
�jEj� u*=g�j��m��m��m��m��i&Ki4�i$�m����m��m��m��H�0^�)�Domv�����e�E�`�-���آBɤ��d�4�[���xtt	$ց��ؤ��ֳ��r�cHX�e-��Qu��>Bo:_�lR�':=}â�����0���4�n����0�1�:����4s��WHBvV�ڃAxX���P�����,C	�kM�6X�qwj����=��4�h�:�;��1Nt�Q�@��t�=����ݲ��1EQó�fHb���W�U}F�{˻4���u��A|��t��Vv�;�%�2��I�v�S��.�u�𒕶�I��)�C7��sO}�L���.���H��6>F���&�}ޯߑ���;�����sӯs�1?8��*����\�����|�4�ǘ��v";�1q*T��=3EZYto�s�*���5k��by8��Ԋ����럲�y�O�U���;���	�x��#�k+:�����G9fj7�Y@y�̂�^�+\_`>5:��.�{��S�7��
�ۼ����M�kf�d`Ȼ�E:���UX�*���2�c��VKs.��h�gtpv�Ce�Z�����VdW*�s;޼��M��"|@��A6�\�y�����O;��%ܽ�sw�w��
1@��\=�4����?%�j�nu�5�����Ov����d`Gr�"=:���E���V��$.�[����ߨp�ԟ�����c�ߘ}9�X���l�^�ߕ,���a�uφ�_��܎�
�TOe�w��Ƹ�˺��b�9|G��5��[�����RT2��G� �͞�~Wp���"UH��4o��np0�{�$aqp�z^�7�j��}KK1�"�.��6�Y��j(�u�{h73Q��>�c0����l̆�[V�����c\�Vn�x�3���5�����yd,��Ќ��kTi9J��om=��T��t���ѕк��,Y6��8�S���iQ�N����WA?/�n���m�8��obk��O�g֝#I79���1(u���5av��]'�z�P��6�½nk�я7#+�T(�06�+Q�;w7��^wq�Z�]��#{���`9����=Z�0�-;q9S%�o��=�/���Z�N���)]���F�j�U��{ޗ}o�ԅ١�k����~�,~��;��t��4��~Ã�~���^D?,��z3�LK7����o�yR��Rw������W����594�zw��;�R_�>V�^�/=Ʒ��;�&��q��cT	`�-�
�Q�ϑ�l�����0�|�/9�+�%�wk6H�k��M��$�*5�y�qV�S�^Ӓ�z�ٻ�]�R���~��k��[����IԮ����3�)�y�e_����'�8��s�9���4�f9���t�r.���#v�ީ���o���Ul��g�֐�ܥ��p홌[���],�5u*f��Y�;���:k]m��{T<%ܔ�@��녜eQ�x@��iړ�wY�ļ�0�,��<JAPtGt;��&�P��Ju�oWZ�`�%���u��5�q�`���V7��x�C���CMa�,)�����K�8��[�K��VxLj�%Ž4Tq�����}�۩}�z\B���B���*C���n�KT�Vh�å��J�W�b�6�iT���\�Y��(=�)y�^��U��.mI:Q����N9�#f�u�%v�M��R�=Ec�f���p������i�����۵ڡ^�1Y��
�o�	�Q�
�ZFw.�����O��t��8��^�����VW��3�|�{u`�9��\�������O�㻭�qw�}Ǵ�u=�E��G��I���7�� �e8{]~W}+�i�G��(���T�nW.��6z�t{c���nϮ�F��Ώ��=vs��
<�U����2Y�^�1yCe-�p�n����9���eM�wr<��5?l����[����K���GLTNk��D�h��g�p��r����Ɠ���tVg(:����:ӻ������yB
�dF�c�A�U>5z�Tk��9P�w��^m�����V�=�Ԕ��dc��1~���u����K��9=�2�_j�yANj��28\�oU�v�
�.\.$�g��� ���NA�m��R�����K�+#ͨ3>tg챶��U��P��Nz�4��ҡ��`MU�ûtl����%SA�J�\4��WW`8�D,[ݪ�)�����[+�,�tCf��ʊ�M����+����@82����uyӖiu-c�]L9�j���vJ�xs�i8F��?��7�:<�x��y�z�0�r��� |rO�:��xyޕ��u��p���V��+OwK��x��@W�1=�F�7���]�+l��^����}c��2NU��<>a�������tb����^�O��T*�|p~�����2}��-K�D��YTx{3o����/?�Kcv�����e���_��~��/fԅ9<ׁt�0�*�����=F�D���.�=���~O�?��a�L�wb�3H��3�1�Ǣs]��E���b�w� r��D��G�;?������Y�O���:�����_����=s����vpr����O�ġ���]�Gw+Ј�B�&UG���g�s�_���W;���`-�U��Ҍo�x߇� 9�i�8�S܄Zv�O� ��nq߈��Ϡ�ّ5�%�xd.�i;���̮������ܤ=y���by_�f���Ĵ?g�'߶�L_�"��ڸ�lsk��$�_�7������s�&?����5N�:�u��o�깕9�VK��p�L��@X�L(J��D��?7ӵ5�_�����yn!�4��&`{��v���j��\������R�8C%���.�ᝓ�n=dS�A��C;Rj�c���r�]�eh9�d{�+�8�W��YN-!5�߰�ICֶR9;m`��w`���1�I$���m̆EuK�hr9����.����U�V��مd��S��z�:�Sг��o(�����pB��ղ���\���Њ}YY��5�Q��j�+���9�DY�����>�B�4C!�o�!�VNFs�*m�_�3�2�,y�B1�\����ν�W��Ã���j��������U�d��g:>K���;�v7�+���cr���]qzCR߰�VA]1�!��ϸ!TL��>�G�nvU�[�OE�	��$��bX��땋��=��]C���u��0O?P�޵�.P�gI퉙S��j�#���c���*B�Η��uh�\̏HB)����3 ��zEP���PP{����:�ag�c��pGt�/:�aK��Kǅ���lעQ�ꡚ�j
G��^)����W����:�~�,���Ў��r?�U�/OG��&<�t o�'�u{�;\�^�C�q���^�XC�R�O
��[sy�x+Kz~u��Nf���v�{'{vj;;f����qIL{.��.�쨹����3N;��ŗ�g�y)j<�tA�j�ܹ��"*3{!�����;���G��-���^��%��m"�ӑ:+��Ä2�Z�\�;����-��)����F��3t^΋�:@��ZY
��'ѫ���f�<3a�Q�K_��l�ɝ8;x'`�|r�n��I�i���&3vOwl�޳4���i��ys���'g���W�Ac2'�i��=���}�ً���=�{Й)�]����>\��V;�/f|�a�r�|	G�Gk���B�8?p����[��j���?0�	\P��v/2��3�\�o�"���%��Y�hȒX�+Dʑw�o�ډ}<���	xXx������ݯx���w؃v�U��O�D�~��z߽gs�hWk�jK*��Oh�1ӕT;��!OaR�+'��w��W�/��>α��߭V�y$�1� ];��1&�So}��ٜ�pi��V�3�eA��		÷M�n2c���^W����l�,��D"�L�>��;�����eG�׉�Q�*Ǟ�~퍮���ه1�~�ⶨ�_\O(=S�����vP�-*ӻ�+>��>��j��6c͋W��ٜ��\+�8o��*�;&�ko�G�Y�����i��c�Qo���>�$w�`�]ɽ��<_�R��J�o7:�W~|�5݀T�;mܱ� ���ݚ؏dÒ���9`�kd� ���dۓEgY��]�[:��v;�{:��}��ҡZu�M"�L�ߺ
Ίjd�0��\k�6���;���:�ׯ%����ѳ��dDWw�ʰ���o:��C{��%#���ۋ�/2�ů�R�d�Hd�0�y���#�{���</�u|�zi������S��J����8����>�i{Pឦ�=Є�үA%�B�>�X��0�G�4m���%y���"d{��A��s��l�y�4Z��qk��=�՝��=��� )���V�=6���}��/`���Z
��m��q��0�< �����w[�)M{X:�#Lh,���~�#�`�Mf��M젭�St�O�x^��U/PG?w��Op�gp�;��9K���m�m�1��2�3G��$V��<P�ES�3lL�¸���,�P�I�~bMfT缣��VUr��*M�'�����2W��R����?[C��5#����VF���܀�3���P;S��qch~�z��]�F&:�c�]]�R��<��k-~�;0۳�/����ȳ.J����_J�s��2ߔ�WY�x�)8��Nh��z*����ʛ��*3mI��:�K�tcJ%�ԁ[C�����z�~����8@[kT�uٓ�ƬZ���_�0T ��tƌj����8�ו�PʣG@��(oqTJ��:��:�C�wE��~��8f�&̨yI��&��o#�����r=�isА���v�˜�Y���:}��*7Kv3r�_@	�|3��зyK�`�|�vۿ�3?M�`���ⱪEq�c�t�F�uÉ,`��w��Y�w5�]Q���%��~4l��K9l�J}�3�`��Mĩ�Ȏ*��\ᓬ�v߼����@�.�/�O&w�{',��q�y��a̞���9U�Rr�^�ثE�V�P ��w0�#�ȡ�E�@�nV	�T��s\d&�z�'��I��k H�AT��g-bs���ß;�J�ѝ��zu]ϤR���<g��F�z�鵮�*��.�z�&�7 z���]3�hn/u�U{��AV�����&7�@7/�=��r2o� �x���'U�åZb���'/W��e�"A��H=�)�%:�����*��ts�����I�;�緘��ǅ�W��nq���+O�%V�Ӄ^r�.��Og�CG=f�>�S�i��n�3��њ�~7k�9H&WX��=��^��o�(2c�2�(���91[���/l�����~Ho�)^y�_J��J����������ز�7��`�fh��z��(>g�׶潡]p�JP���M��ɮ�o����y����{i������4�R��4�Zӑ��\���;b#��tQS����[ܷ�%̠Bc,��x�o	�!��ۘ(1�<.}�1����W��4�m�I6�o�\ٿj�@�����/_z\�.��;m�ݠ�YHue��	��ػ���t�������!��M0��>�m��଻t�$�	�N�!��9�o�E4I�^Fu�>-���ؙD����<E`��mCϺ��}	xM�B/�П��'W?���]��TVu)&$�}�d�B�N��,�9�؜&X�(y��<���#5_^��S+��o��i�A�~^��Ы���̧)%X�y)d�8�%ζM�zs�q���)��Q�n�t�c��a1ߏ��r��Ŧ��G�����|����{�1�u���~bJ}G�K��@h�_{�][��L�ί�rɱ��
��9e�le�7�Y>�y[�AJ�i��/m1~R�
o^���&�=js�+{!vI3�cu�� ��)��nv�Z��Ts�����3�vn�Z��=�|�`�[�vY�F�������}Ns�7�瘟t��@�ҨجRC!j�qD���n��)����|n������OD������׫�z�w_����- �z��=޿PM$?V�/��9=������v����{w<���U�h�@��61S՜A�)}��{>x�-�f�[N�9= ����V�Zy��Dі��8����9RH�l�������cT�}�Z9���$ۼ�C�C��t��U�W���Q��<�0fn���y���5%2��}t��R���)I�����3�N�_��[I����#z�;�`(7x|�qZ<�x~��Nx�����!r��蕚��������g?y)����9%�H�X���Ozo�ED���F��6�w~���r����B�e��4\r��A���t{Ah��ׄJ,5�;�NO�#"w;٫8~BS�ţ�Դ~�K�"��#ջͅ^��r�\�d��ٙ�.��eH79��Ms��v?a���6wOڿ����7{w=�]�(?�1q!;鬝����(�����v����Z)U��UF���m�ߥO���ݹȮ����޹{}�n�x�<�w]�o � �L�x,n�AoR�z�5ޚ�됎x9��	nmJ���)ZOнvq�������t�(>ft�>ǝ�j*��{g�t�'�E���;��s��=s�r޺p�I[1R=.'b�Ȋ��ͻH9�S��?�ǯ���z֚�hF�eJvk'��*/I�9ꕘ�e��������`��'ԫ����yuL�����hOe��n�n�����.���B�VuKy�^��v�g�Evٯ���du���Y�1#"�nH��++��/BZ�xqoԷ���e)��4�M�Ů�gHz<=H.�9k��\+Uj@�\�;��Z�=WP���0��pwI��k�Vdi�/�����\f��wr�s@i-H<����yWֱP��&;w�ê;ZN+�>э�$90�[�Q|&SF�gø%�F7���WO��m�[��`8qRw�c��^jRzwL���¢�1�"(�\徭�W+�ni�]y��鵽Fq@���w��{����C
�:���<Jb0�S\-��q{,��@vm�e����T��΀nua�t��8�Kp�ٵ�a����m�lWt���\����9ҩ[N����ދJ�0�Ⱥ#]VT�;oy�GaÊjEYa����U��8%n]}�>�<�}���x���v:��JdG�{\�K��ܧ�3y���� ��)�
�<�w�q��#�mn�I���L$����t�H�\���6T:₆�n��+�k�������i���4tA!޶POV^ڻ���Z�g�	Ƴ%_s�<�}.�u��Bj�#���T@��:�]���P��t�S 9��Q��[J�c!���r�f8��+q�ע��2gX����;��ʔd�ғ��-#�q��"Χ�÷��U��0`�ݥ�e�A����CWR(��j>x�Q�`\7��j��u�>���Cs�U/��:EWk��N�iH]��#_�{ʖ�z�*���Zedf�ש.�c�}L(��s�l��i�`��w&�$�t3j�ū]��0��+��+���}Eκ�_U��Z/r�����n�pT:�r�\m�����݀�T�������sv���'W��P�Գ�ba�1r�X�ۻ��F�-�2*�z�󑀽[�D���f�䊊��D_n�F����hWZ9�+��tk��,��bƆӱF���˯p�n���4C+1�����p��Kg�\����*h�p�pҞ�ч�[һ\m�c5lT���T��hҳ�4:���i��pĸH��.!��:�ݸ��X�EM�q���VA�u��lT/sս�8�As�$���k����)�������7_cj���c�҆��X�vF�ƕm�[���+Okac� )ta�B�Q�.�f5y�N������mhД}[���U��Ș|#յ��yY�l��1U�D���opv/��;9Cp��4PޝÌPȹű�R�Y��B�K��"�Q'�L���HX���;Gr���<{��e�k}AMUE���׿i+i5����5�+��SjD�˫�p�b�����5(�;�!I�VI��{�Q�[[h'�_U��ǲ�k�I��W�-�H�&�j�C]:�7jhMG��'&�i�w��WM'��}_}U��ƌ�J��>ci%1E��V��g�=8@�:�u���u]�
�J���0jMx��X�u,)�������w�����Ꟶ���� i�W�~�U�{�÷��^^�y�)[����˽��_L��ǽ��zV���oy���y���"�r�ǔ��3(;�2��V��~@*4��d�§���B+�z�*r3�GN@��-u���B�Bf�'�
��uw�����oU�~J�Ol���@ޮ��T��	S��V����?O6c?�j�^s��\���xG��Ŧ=���W;ɪ��ص���*���� �������/PR3K���\��z��#��7Z���f?Ӽs�3�3.-u^7]�aTU��6�\�@��U�����Q����Ó�¡u+�� �=��_��(��������J�;�BR�#o���`��<󌲞���W�b�{��l�l{��Pt�݄��l���rN��mxXy����u;n5b#�g�"����>�n[���j��[��w�����P�<��_]й������]|�S-�z�n�dv�`����Jwl�d����E����?�,s�{@N����&����<��i�eƚ�����X6��-g�.�`t���^�4Ê�a)ס�Z��&�p�i�N.�a��p�ܔ���x�W^�1�﫨��NK��tx^wN��&���H���MW֘w���@0�v�!5Yk9�s��ۧ��Z7�o (\?V���]���3���deˀ��u��dQ�RJi�z��(W�|�qGNS��cs������)�Vx��bO�CTgw���M���O�9�%��9:�?��W�l^����Q~&)���yWq��B��+*�����d"�r��������O����Y��w��L簻�%�m*�
����/4é;9��d������o�r%��2�M���+:�;+��E������!f��&d���yS���x�<��ܖq�.Y	��NH�_��z��c�Ǎ��w\��tW㐉�5w�<���|O��ȥ���Ȫ~k$F�iN&燞:�d��{���%G�	��T&NY彷��}�8R0��X5�2��9R�,�\6F�1ܠ�K�p�m����P�S�D��/��oA���w��Nz�a��%wJEd�V����v��3m�,/y����p�t��"�y�c���:���.Z��V*vj�����&
�8#�+kjޛu�u'����cZΗ��X��\���sW �8�V����(M��[͜UB�{J�����P.n<c��#F3Em�Ͷ�m�����HR����zy�,�嗲qC��M���Z;#�ћ����`�ܛ���`J2�zrzDQ���c����Ǯ2�x�%V�e
誧c.}]��lƮP�<����� ��=X|�Չ�+��鎃���}.r�gg�MNu���n.M�k�D/���|��z-Ͻ�%�-�s��V�c���="^IR]��ʬ�Lvc�����?[�G������#&��в�w��,��N^J��܁��u]݁�w���%Yf}v�C�wD@p������{o�U�ߙ�-y���?b���w��zs��d�n�"�f�щ���⫥�c�-���������y>^y�G��(�'�|�\�?+pob�ך}vm�z�o��3��J�`�\=o��f���G�C�����^iV���C��nf5�v|��\�e��f5kS�<�=q{�bB��92� j�d^uh��a�GE@G���^��P��3�ڻ�2ϱpE�v��O��6�#�#U�}y�2[�m�딶�����Vfyv�WEkX��tQ�}G������&��V�}���%̙��d�1W)q�F�d=y�
�]em�!��!��Q
50j��[ڊ��ʤܕ�c�P�j�2��y���{��*�w�N<Q��^!R�@n�Mn+�}{�sbrv��l|Nweh�/�w,m�0h��X��G�f�O�gV�Tww"Q�k]���eue���M�e{šk�{W
�⽽ם�I�`הk�s�NkwN�ߑ'����8B)H��MPR�	�wNjgn��G�������v~�=�'c|�0ϗ�{gPs?%�$��罽*͕6��j�5���9�x�ȯfѶ���nu�s{r��4����_�_BM��ez���6���F�?GU<��J���0�&�>��&&��vF���,ۡ���.L�x8>É^/Ʀ�Q���ŞX�ڂ�;�̘ԕ��zE��}wiX��J�ZV���~�)W<]{(
c%#�D=�ap�9
���uG�ώ�?�hHiw��S٠������J������=R�A��bq�:�.p�pY�vi(�궣|E�.���X��c��y/���\�?`�T�Юk��;��_�h\�C�fwQ�J�����{�d�c�
��ç�Z�.[:p�%�_���^�"B����3�m�=f���HC�%�7�A����
�^L驲�cS��
�i�uHu�?�9o訯~�P8�R��YӂJ��eZ4>P��ۮ�!>ՅQXtޠ�*}�fK[��7}X�I�.m[�V੻����oa9��زn�fG��!	��g5v�d�Um����1n�o%�F><��ݭ:^R�<ڢ�T j��5qev�E�/f�j�3�x����#"�/O��J~���KS�eM0_����W�g/s
��z�h<L��:$[uw��}tfxIeWww�?L���V��܊�w���=��]<<޿X��g�G�ػ[�j{WA�tݼ��f�	�O�Q�>�+A��Ll֣ʖx���$�E��x,�q��8�w��ا�$򬮼��CN-oc�C4�u�v���=&T���W2�=(ӡ$���p��=8%#���U:,�.s��$�vlN��}�4��3�:0r8�����u�s�rji��l�%t����������`�5!�5���bVN/K(_�%���LR��J�aF�:��g
 Z'��D���' ����+�����_��젽��|�AN>�{n�eE@�!oPE�Ѥh��h�C��6YQ��Pf�H)]�z���z�E�w�w_��v@��z�uY������(����&�'���&�{�a�8~'|s��ݕx">T�`�V��_P�W���\\��˥K�N~�W7b-[����{Yg�c��%t���M�tM��n&T�ïc�j��Cn���Y[��	��D��܈ԭԂX�wث��5,>ɫ�L�J�e�\o�.EWYb�.c�f�3dV���,��X����ڸD�K�G~������Ar�3���¨w�${��Q���+{�sVV���LJ��õ�y5�b���e]�P�����Y����}zW����'c}�P�x��ց`��V��V�
�/�n�nlnNn&�������}�o!�3��S�|�C�<7�{��w\�\L��ȁ
�)ztd��gd��=�̲ugL��N0w���nd�s��x��or�	�= $�uE�djtI�#=�_�Gy��5^��w�<��:=�����z{�Wt�g��.�	��i��Qe����8˵=�K1�`��W��.m�m`
�����Q]�g�\�|m��k	rA�<|954Ö���՞�*2+iˆ8�a��7Yy�x�}>�U��\{�.��7��G�D�1X�۳>�jb��W�D؝f.n6ߓ���j�"͇�c���g�w�k����-�$g�%ȗ �L��ĔW�z�8��>}b2��2)G��es��	Η�T�\���;���*���	�������ױ�x1�w�
�	M���!������y`m9�M�B�V��j�K��r�K�;K�&�r�CS&N,r���Z�������&��Ck�e�����'Ҵ
��3j�i3U]`�BZ�$�m���m]]n�$�*m�6��{:i.�::��vI6��/��+�{>�]w�q���{!�R��x뚝xn�[>�,V�t�VybZ����eU���{ǌ���L��1hd仾]��Z�㞻@A7������٫�F=�IG$q8N�⊢'�ϟ<|ch�=��<����t��3�d<��S�4�xّ����?N%�t�Nm{ҹ�sg��}�����u{���{J$�C9�oD�(���7���7w�+�k"1곣�����q^�a��*|��p��5x�m���z}'��.���C���<dU$��u-�#�B+K�lZ��-��D����yZ���G�B,.1�>w��������U{8&�ה'�!�eVO��EI]����w����^���Cw���D��{:O<#Պ�XVN~�V�?�0����{9At�����vg{.�I*{K�Bg΢��͂�E�f�=�I]M������cۖ��k~�7�&:r_����U�O��z�,{-�X�*�C7�z�#�����៪Eg�e_�<�Ï14*6�3������q�2c&h^*����oIL2a=b��Ej�=3NVs��Y��y���������w��(^��,!�,A��mcE�"�Z!�����B㋩A��:�ὄ�u�f�]t��mM�a�|Q1�%����=0�rX��q-J��A�1��:������N�M��^��y�q-��RӺ�ƍ�X�����N�7)z�֍�{�ݵ{�B�E!�m����1�uG/V�[�(P�uV�ܣ��y� ���1(T�<g�ZTrM������r�;��'Y�k����'�*\j~��+���麻W�K�'���=�Lw�9[��T>��y����y����z����K2���Y*�����=�Ew��J�
�W�l�\�Fxn�|�\,���6�\Ԭ�韎����'��^���hI-���+l���	p��Ȫq�z���u�8[�:탸w�Hp�j,n�W˨��'DG�<�$��sҦgY��m�%�Wz?�<���V^�
>��M����m[����|V��5M��[��DulY�Wq>��'�.c��Ս�׼��d�Z�{���v�V���t�q���k�6^ᝉ��e�fWD�~�v�-��+�a�?��b=���s�O'*�]~\}��g���CC8�_�y��a?oe�9���i��}$�1V9�q ��z��P�G�����Aۥ�f<Y�P�0Lr�]�n�r��])��cޔ�,�e�&�-��gR�Yܦ�ƄV
��݊]��]NӋ�v�=mU�*�ٚ�]���{�۾EK������и�h܏����
����L�iyY5X �;���.EnR쌅̷�z��n=��7�r��+YJ^*Rt�q��
ű�Do��w�G}s��be$a�<���X}B����6��L��R7�מ)T��O���
�xv�ڮ����^Ì��\�}��]���$�p-w백%��ef���s`x���M�- ���M�h�8'\�]�S��\)���/��Ɲ��$ى��P��TQ5�i�#�6��\~�����Y#G�T���O�a��wmz竝��G!\��F��s'�uʮU�	����4��Ydd���M��y��{�ȱ�Ն���	>�
��9��I��}N��]l�R�̐�>J_we�`V�7]Dog���s��;�Jqu���D���S���j��]i��n<}��7}�Yy�aԦo۰0v��ُA�rT0)�� �3\�O�@^�������[���܃�\zs��wgkid���]<�T���p�CUky�n̐E��6���F�*墨���n/=� +��U����W������:fjz����w^ps����1�O#�X[�嬾�|��.�:j����j��_5 ]ʬ�}�/UY0�*ҚfwJ�c�ˍP|�4�\#�t��p��}��	Gu���K�M-�㎔�xX�aV�d��X_ފי���D�ڇ��]�k;&�����y41���x=�P ��t׫Ƭo%���]{:�Г̌�q@�}"�"\Z��6��ڳ��;��'��zM��7�f��\�j����W��QIue���ݝ)���V'�'*G8���5�7:� O-�D}���㶏W &���/d=7:.��w�Mr۩)���w��=� ����ʟ\�Tf���K���sc$�N8�������O����Q��c�c���o��:�M�k�ޯ:>+V��Зs}�},��r%N��ۡ�R$@��8�S��k$P�ݵ,�eɖ��k���gǑ�o��\�/N���ܠ��5=�:LbS8}�.+������yGU��+��^ׯtGUڒ���Y�0����3E��s���?�=�.���*f��4������=/�c�ެ�@��>�2$��n�����DW�<x���g�R�ӏ ��t	�^\4ަ�U�h�Dm����TY��HJ�!~NQ`p���Q���*�LPz���]9}�^�Z�<��h�C��T�l7b�m�}Ժ�V�,���$#r���:>�ը8qȸ/�@<W+���%tk*m���b�w�H!-͙MxR�z��MEs;���i�Jm����
��4�j�<��	k*����^��].J]�b�E�$�+&N�S#��V�o����+��M=Aq��×ݒ��I;V�ވP�V΋t���:���0e\�w

j��:��u3;Qr��ޟg����y��)�a �$���$�w�Y����$$�BŁ$�` ! IE��BI��@�k���ЀHO�?��$��� I?����?��O�� I?�?��/��,���O��%����r��?�B�*YB$�MY�I�?c�5(ڷV�T�1�;�*��!\����5(�Q�Ǵ��"Z`tj����I0����%eUښ��n��{�fꚗi�xha�B��71���Jٺ��d"�^^�!K�4�f�{&#!qڲE�����S�z����ڱF�	��})�(�@l�y�跘K�:A_l�1�E�F�2�����y����5X����Z��Ս�3a�-�"hV�yX(��I&DL^�d�iI*�,u7-@^XT�9t%Ӏ �r����W�[�����8.@5����p-��3��ݿ�yyZ���5�n�h$�X�e�f�FSɩ����Ꙫ�z!��̶��x�WS	��72�a��-Yt+ rd�c̭���Jt��Z��L��it�i���c.���0���bT�fBĽ��V4�aZ2�v&�DepEr�wVZ,�U�[j�P.��j[3%�e�0���"��-�d}q((�t-;ˬ���f�hԥg����3cJ��R8�m���&*YmS���6l�vI�d,�]��XڷX/+*�� l�4YWi�e������%��U�u�]	�YyH�
�^�j��4�ҭj6�ݗ�AHb�q��Hء2�3mX����y��y��Xh�
(��^6Y�LZ�fnb�Q�6�ڦ�r�F�5��.�e��6*�S4�c2�Dn��bsp�H8�W�%u%
֙��f}t��EfV0m���L�İٔ���Y�aށZ���;[�e��-��OP�����wY�x�t+j��j��&��J�k��Rh����	q��̨��@1��F���Ł���ȳ���hɹHʻ̬�g�Qú�J�bˉ(.6q{4�ysr�D6#�LЕ�9O�����7W��KVT�nP��҆e�,�"U�&��ύ�Ma�F�7q�t����A�Uak0�Uv���eK`�,�E0H�F�;2��(�/ݷYHc��%V�0Ԗo6+���'6FӋ@Ĩ ��ݩ�WP���W����t�2t�I���	��A޽�p!ĭ�������bSTd�S.ɳ,�@�[f9z����Kr�^*Ѷ���D7��ZX��b"��'bX����y�ݷOwF�h��[�Z��涪@ȥn��Ԃ��FA����IZ�DOe�2E�)���q�J!�����p�?7��6u��Ͳ\�p��7��-�8ȳ��[3&��c�yLޭ1�+�(���d�$C�Nڽ��Lu��Z�wu	J��m��f��.�����Od����u�-M���!t2���[��5M Y[V\��J���e�����S�qY��{(�M�֮�47�s]�V	Wo�l��^���R'k�*byv��Ă�ܔ -ظ��3jZv�z�gjL1�+f/*KN�=)P���SQ�F�-�t�];@��S���#�����ԼŊ%�n�щ
��6�-�Y(F� XwA���j�{cf�I4��X1������i�H��Yb���La��z�qVa�	����;Dc�쫍�n֥t0�TK�e�fV�ڱ��f�B�!���$l ��T׋(PI��\D�K�D��8v[�R�u�ue�)��1V��D�2L 7�i��OD.�I���h���ƢX����jd�%Z@
L}��8��r���� �t̲�3�6O�N֚�%yD)X`]�׳t$B�[g^���S�!��r���|):�h̶�e<��V�7�̷�:��PX�j����Qد+l�,#F	�U���]]ܤ�-H6	f�3r���7՜�>��`�2%�� �.�[7F�h�;�]Y�
�)02l v�);��2��fDM�&-ó������{a]X�C^�խT�kT�O���M���wyk]�y�rG��z��Ha��I˩7u�Rs*)[���a�p��� z��VjZ����R��srT{���8�<�,�jRo�Ae�I���^Ir�
ݻ��sPf�	�����n�8�w���[�Pڕ,�+3��&m⼰J����
��YYh+M\RY��ހA�-��j� 4�4<
�V�jm����6����ږ!̄��n&�*#�T9{z֍kf�0��0��D��f��#)T��D�۩q�+Sޖ���41�)���x�TgY��V�1�����K���A�pu�PS���(da�{�T8�J�2�kSj��������y$� �2��H �  2 @`B��! �I �$$�a		#	$���! A�$$�! 0����?���x@$	'�{?��t��A �$�������o�~�@$	&�7�� �ЀHO��� ���5��HO�_�f�������$�B I?�_�o�B I?�	I�����?��ۚ?���� �$���������$�B�	I����1AY&SY}]K��߀pP��  � 7'�`a�  z�  �     2 $  P   @          ��    �P@ �DQB@ 
    �H �              � c    ]0����>������`��
�����������[�.��;���� ���UT�h���$�ԫ��[�dZw�r��r�j��N�R�($�T�{���շ����T��N���v7� >>@ @  
ED�]�֯{ޯU^{�=f���������4ӞRB/s�4��ҽ#�s�ҵ�wz�R����X�{�(%w�*^库f��� ��^}�{U]���T���=���7zV���ޕmg��U<m��x��U�Wz��]�t���=��)x�*�　" 
�@  !Q �=^6��wIz��ʪ��wV�k�Z�x$g����ֲ�;��=��zS[�s׬���B-޴�[�R��w�R�M��Ji�i͕w��Kw�����W��.Z�`�:��[�S�x= �=)�W��=[]�=+K��OT��\Ꞷ�x�   D����){�t��7z��(Y޼����u:km��H%�T�[�t�W��ջ׽�ZڻםzV���B�U{n����wU�kW�w{��s��nx���Jj���ʵ���C-����k{ۇ�^x(	�^����W���mw�xP���P   )H%p:���y���w�������(��X�/a�gO@�ۧ�^{ ����k �a�`�=D���!����s :�_x�z]��ꛭ��< �~��*�P 2  5S�"b�*�	�L�&���mU*���A��dɦ��تTM2�   ��5Bf��F�   $�@��h��I���c�D����!�O���9�w��3���		�~����d�@ ��	!! �����?�$$$ �I		0�BB�����S�_�[�72?լ�wL����X�������0�me�3��т�+��&d���$�Z�+ЬB�Z�0X,�`�a�ĭF�q�ow�/l8ì?��XW����I�4���,aXsRϘu�a�8��ì<ì��vaXq��,}k-�ZS|�/wq���1�3�%I�7�CYJ<J���bc ��aϨhT~�0��пP��v��!�(y��8��aX|�����ق��q1һ����޹0J�J��*bwّ6����{��'�=���w�縷��<É��ƭo�fe�yj���e�_`�팼!���Ϟ7���=�'w`�c	����ˎ�o<c#����[Q�V��6�m��fe�m������Ls33
�(ԣZF�fa�3��L[q�-�kB������+��`�F��B���-*�YD-e-����`֫X9��`�JZ�����l��d�e�&9��	Z�KJ#��E�n3�e�Jб��B���ҥj��32V�F�J�.\L�.�3(W#l�)F��L�Wr��eua�ļy�LCC�E���������ʖTF�Q���-���Ђ�e��9�pt"-�Y�bn�3�Q�X�*�T��q��=�;�1�u�<�1�k8�L4�û��'�0������(Z�����X,:�Q��?����7�/xLR
�K���Ue��9�pCmd	�g�7L~
Ì0���aY�aXVa�Xu��q�u��0c��a�ez�c!Xs�a��u�X|�L:��0ң���L1�y��q�Rc
�l��m�ì<Û��0�aXc`�������V��c������aܡ�CyC���u�uc�
�a�
��6���`��i��c
ì�]��L>a�Y�a��i��Xq��1�Xc0�a��`q��4°�!�<���hg��߹�xr��jcC-��k+��m�j�`�
�,��`�*�YZ���YYZ�(��+X,��Xq���ed1��`�X,�LJ�`�X,�;fe��`�X,�5���`�X-e`�X>��`�X,��:�X,��`�D-�X,
!5�f���w�to�
�0��OXm��|���ݡ�a�Cz��;l>a�0��u�>tg��o_w{�~�����sj�L8��8ÏչJ!�Rbh���X(Q��\NZ�d��s0>a�
i�R�+1�&�r��R��bc*�U���5k$�0�:ì9�0�0�1�Ú����c$����c0Xq�Xw�a�a�d8��4��k!Xm��i��,8�%a�2��+0�0Xg�o�a�a�a��<Î3ް�0���X����rèq�=�x�ָw-����w�,<Ü����1���aRc�,+*)q�Xu�XV��N'5f��+�d�\f�}�sP�
0�e��s)��kX`�Y�Va���J�J�V°�a찬=��a쵕&��պbÙa���������y�m��ì`��'I��W�5�`����Z�p:���{��o!����.��g.-��V�݅�����S���8&�\��Z�ڙ�F�F��o�f:
ھp��Uְ��e��D�5L�0��V��-��m&�H��#�����I���ZIZY�>�ˉ��(N��n��aUj�� Ǵ�~K5ۈl�7l+D�����M^ecƚ�0̮%]5G�]����8�4�y̪">�ˤ�i�I���(��e�1���~�]���(u�ՅլĞa�Us[��8Ԩ�U�b�<� �RVI�ՇXi'Xm'�)��Q$�$�E��s!XfXq��y	�H���C)<�6��B)X�Hb[B�����Ќ7H��G�2�1�#��m�T�mMY�\M�)U��~�>/ZՅ`�`�
��
÷2����3,1��aX:��5s!X6°m��fXWr�e���57��W�T�>�wT.�%L�q+��B�������[0̰����Xq�����a���
0���>�9��Ùa��a����[S�[m����;���!��Rm�fXcn�k,8�z��J°̰��0ia��!�a��Y�q��aRV`���Xu�rV�4޳�]n���>�3,4���Wr�j�cV����d:�7aX6°uaX6��t/����{�{���\�E��e͵Ĩ��S-�9ar��
���l+[
��1.f0r�2�ܰ�C��B�iB�M�
��,*J°�̅`�
���l+�V�IXc�V�Z��
���l+�V��aXn�B�m�qp�\`�
����d+�V�N0r°m�k>��V��uK�[����;��ú�Q�q�'���,:���F�V��aX6°m�a�̅`�
���j���g�v��.�c�M"���ua�޲a̰��l6�2�<`�38�y����;����9���gX=�C�=�x��°�Xc�Xl�
Ùa��`��m���̂��0m��o,<���;�6;`�%��i-�ĩ�M����2���bͦ��>J����-����u�
b8�Jȣg����hx�S�&�V�YHy�U� 3+�
��z㨣8���A�ն˫qM3Z�1�3&>a�Xc�0�Xc�k���r��Y�,ݡrì=�a�3��Y���{��ֳYa������?j���UDťM0��wv��\q:��lf8��̯�16����*�*�m9�s{�hE�(�z4�����K�Ҧ!�2�败�YƺQZ��Wy�b�Z�iAt=�dĩ�f�oT5�Z�a�L<��ݼ���.Dy�hwVR�H{,6Ùa��!�a�;�d�m���5aXs,8�2��G12.Z�hV�She��_!U�ٙ���YkaXw,:��d9��V�0�0�oKo�AEmY��
Ù`��a��0׵��XwT5�,U�n�]�Ն�n�M�`�Oe��WX�5G)G�+�V�N�Oj�e���Ì̛z�ڰ�e�{/Y�SV�̮��m�0J9k;���V�
Ì͞ˉ����a�d�VC�̆�fXy����+����}�oP��u��ì3,8��2�y��LN��a̲l8�{�Cs,8��0�Xy�r�g5��e��6Ì3)����a�m�S�&<��c�������"�e�DXy%a�`�F�~�C��0��̰��$�Xm���e7������W+E7��^�c�̨֥,3ن&�{V��!��Ӗ��q�b�YL��fE��a��9a���V)��.Y9t9��Tr�5H�0V˂���!��0�S�����b����L�(�a��ֲ�YaXk,4�[���¦��YZ�]�m��x�{�Vq
1�=q]d�K�e�6g)\+�
�5�摶W�LN$�te�<�tQ8�4Xz��U7e5�
�晘i+�*<��s0C���r���;���Lա���7�d8�2ì7�Ҵ�(���3���7l*M0��Cl5���)����ڸ'V�^IXy����öì(��\i^Ҭ�S30��4���{B�Y��\��Y^�0.��j�:�kU��.Zֆ쮵��Q����*�ը�YuL��̴Wl��Q��׾��~�ηwɯU�R��mr�L3w�%��VC;�N߲��׷���_����P���V���R(
E�aUX��Uc���QF*��Q���i��kb�Z�[l@G\�:,*T��,�Z!Z7ِD�l
�aR
}��Z��XT
�ĕ�C�q���D��#s!Bb�"��J�+�EE$Y���c*բ*��jT��t�%���"�kam0�S�"��*������"1���Ujإ,i�YQ1�E-b�"VABDUUTE��Z��*EE��Y�(�F,���X�V@UP�ֱdR(
J�� �ZҬUT�����1�c�+-�f%�VX�ČH�"��%TX*12��QPPF�Y"@(�DQ`�"�1Aef2� ,PR
*�X*�1�Va�[\ �֥b,��F J�b�TY"�,\`-TE��¬2��1�R��BQ���1+
��ڮZ((�"��R
�B�\X��T�*I���FȪ(��Y1 ��)!��UF.$*E��s+2Օ(��V�K[l�!�L,eB%\L�ʂ�m(�*�Kb�Ls
V
�R�R"�f�$Qd�����-aATU[Lf
b�"�X�"�"9lU �UUT2��a"R�TX,q�1 �E!R�T\`V��C3j���(�j�h����(��-T�����fR�֖���DQHal��1*,A%s(���e*�Q���C��(�E U3,�1�iej�����T�T��TUSm%EҪ�1m��,ı��AE�֑f0�a���X"�Ad� U�K� �Eq���E��%CaE �
 �dXE�"�0�ư��*�`�Q\�+PY��`����T�X�-��Qb�cp�R����V��Hc)"�*$B��&2VJ�C
�b�
B�AH)�-��R) ���E��ąH)�C-�YR���C�R
B�3,��`��HaiH)%T@�UX��F	�H) "�
� �����C �2�
,��m����r �Sҍk)n.?ￅ���{�� ���p�� �p�<lpz��U' c�����` <� �i�T(���^VyvJ ���o'����m� ����=��7� โ�Zy��*�@�ͳ}��U� <    P�     3�x  m�����<@N��8@x x8=׷z�߻ѫ7�a������{X��Þ�w(�(;�ݗr�7\����^q��R-���v�oc����ל�v�ܜ\����{SU���v���z�e6v�à���Q�e����ɂy81s:���g�(`��3B0X�n�{tT�yOF+f�cf�ci��//k�<i����[b�q���yf[�i1����n��v.uT��:v۪9��Em����x��8^�=�H�B�;�zѝ��lڙ���Ǥ����l�p�m��riv���5�Uy29nY�s��+G��㍸�+
�wd��xx��˃�v�����[����Z b2v�r����u�&�skA0q���nn�u���Q9Ό�ak�ӻd˻A1�.`��e:�ns���<�;�^z�v냓n�<c�]�󛛶�FvN{��6�]��<���	��{cp��Kva������n�Cɮ:OH�*�n��k����vvb���{�����nۧ�ls����n����;lon�G��p�z�n�?o��e�c��s�y-�Ǟ�V��Sr�GG�Ӊn�U�Eh|�ݚ�]uZv��쐚w�W]���0=I��z��Ӻ�q���\n|��v�[��\�s=]$��i���[��;hh�--
����B�@U QT��UU
�  Y@U��@ `  
� +��� ��ڲ���� *���
�P���l *�   ��5~Zp��GZ�E��Ndcm֥�oUwl� @ \����޶���l��mm �     TN탤�1є����-�fU.� ���/`4�����J� Y׳����ݯ�q�a�*mp��T U  U �� 6�@@  [ �ʀ  S` Y@ �     ��x�h   �3r�VM�t�y���u��@  �@x Eꭓ��-t��k�B.J�u��R�K�;e
�Pt@)�����]5+��� ����p���    ` <  ��uA�� yYS�1�p��+)Tzڪ7s�U6�૫P �z�P�򓉵��ݷ5�� @�0N<�s����k�@w+(  ݶ���d�lQT7]�#�g�p�T9W����/fT򢙬��2ǧ���)yk�Y���0��˥W0z�n(!��� 
�7��־�  6��� ��c7j|M�(��)�Z6Uݴl�a{�KT�m�!T��k��@j�xصĳ�)�J�]! ���V�HUUN���*'*�b���P�6�ݨ��TyU꣺�۱Qlz�C��v�Ek�fꊨ:C�S��p����[   +(�q���� *�| �8w&h	mqʬ5�*����b�EUJ�T���j�R� U*� Y�U[̡TUPU �n���/*�m�J�R I K:!R�����+,*�@    �b�.ꪨ�R� *�T���d�@ �T  �n�we6� 
��  6��Qm�@N۱=�UT ��U p  ���9[Ume�  +�y
�v�wn�UG�@ P  >�� USo�ݶ�����h:��e[h*�6E�xu�U,eR�8���p�[  mP��^�*  Um� Pol��=Tz7H�~>�i)T�Y��Z2� �p  V]ЫW�Kf��ml��� <d�z�8NU{�}���heV�r�RlS�+�A�^ Nՠ8@  '
�u7���P@'�
 <U p0� [j�]YZ� D⩌Ԫ� v��Pp�z���5�� < 
Ƕ�5J��m�7쪰U�eU.�T��W�gU]ҥPP� `  ^OT`j��T�pT U < ��       �  N �   ��   ���     *��T @    �T       ��-�EJ��z�    p���	�      �     *�T �*U{7]f���m�QT  2���[v��",1�E�8O]��^�JL�&d		��'h�A]�0g�YTq����9�V*���6���[L�͔��& ��m�i�d��R��36���)���O��[�ę�ZU��5��� l�kmP�-��ڥ-���R����Z��cxYyƘ�{B�Y4E���GF����m��{V�lֳ�R�R]�3q�Ƀ��1�h������#k&�ݐ���%]m�qDoQ���M�M��J������cnx����=�8:�v�]�v}1��Q�2fv�]M#W�c���X����U4l0��֗bۑ�dJ��"x���h���N}�{6��J���ƃ���iR
:��Wml덐4��d��k-*�#��*c������q���q6['q��_Mn<;�5�����W�)eN���.X:]mmLL��B�,r6�0v]��B��� ���e�I殔vV	�JO(`�s;g̓$ʛD� 93�L0�es���K8y��˗j��  2�r�f�u��rP��,�T�G.eV�&B횶�VV�l�3F{�͆�&s�����|'�8�-S`q$��TT��Z�nj� RY`3�i,�W�w�U��r�:�4sS���X����U�jB��(��B�95NP.i�g�3؃k��pl��q���5n�2�=i6�k#�5vไ؀���*s��a���nx��`��n�Y��]�� !��\jNV���jx'mY��um����U�Zxu�1`�.9�[(��b "��fC��0UUT��d�J�"�v�v,;��s��H\`��Ů�;��r� �|                  VP       U �*��                     *�J��  *T   ��@       U 
��>     @    OTT�  U  
�     2�.aR�P*�*� �      U    R�    �  T    �|  �     *� �(  7v(�3j��U@m�
�6���}U�U*�P`    U �PP
�                   U      �    AT  ز�      _�}}� ,�@[%P   
�� P�    ��    �      
� @          �6@  �ʪ
���h  P"Ԧ�����Z��ګ6������           >�  T*�VQSmK�*�             *�    
               T      �@ 
� �>            wr��TP     
�ܪ*�
�T6�            U         
�     @ P  w<��CJ�             *�Ҡ     PP  m��  @          �     m���U�ݶ�R�n�k��J@��(�    �6ʀ  �5�T���z��۞�C��� U{'����e *�� ���eT �      @  8��,@       Ub�l�     *�TEm� *TP��� �����  �  T��U7[mU�                  T          P  � U�T             �fy�v��� �> �)�UU *�UU � {l`��  �*�uN�%@      �ʩ�;���ѵ�7�� U�� 8J�mE[���]w�;v    Y���[�� � T[j�(    T���� �Ÿ��録��n�ŝ���üT  ,2�@
�J��6��	YZ����b�vG�*     z��m����e �*�b���m��2�  �w�K�?n�X�� ���� ���wo֞[��^� '����{�@� w�k�;���z�1�p�� ���X�v�Y廵���ݨ [���P^x��z�.;j��\�,q����{��x��|�BB�Ԑ!$����_�`��I %������kZ��]j��TN{'�1�����7�B��M�� UUݹ� ������*g�^�y��x5B�`��U|��{gpN{;ٰ�]�mi�Ȼmַ��k��s�ݧ�g��bٛ�ݰ�Y'Qt&��c�6{"�)G�j�h5ۥ�c�3ݝ��];i����y��Ig�99A.�3h�0Um��U)� �@�]��;Wt��@6� ��aT�������bZ� +̀  yTg�s�<��՞�w*��v�n)�]X ���3��<5H��׉�<���(���KA�j����=�l��b�譌��mQEQ�򕴫�Y�y܂� T�w��lVJ�W�:+�6�� z PUʨ�A��T����OWs`���s�5+%@m�pa�텳���+*��r��l�U�r�Ψ8UO  'Uu����-@� < *� �PW� � W0 N   �*6��x V�۴�FM����7:Y+"Ԩ
�J����]����:��ֈp��by9;tl���tk"�Y����Cn�]�۬�wy��*�l<=
�\�q�s(kfk�p�7Y�2�e��.����p�eŝ��ƍɹ����.�; -�1٬�l�\��I�������ۮ��T   U VJ�       *�� xU  n!UT   �UP ٶ�U
�*�*�      U*��UR�P *�T� P
�Yn�=�� *��x�   �  
�2�@ `  
�   � ��n  � ��*� U �[j��@�F�0   J�l  � �UT         z�]� 
�V� *�e�����)� �z�ڭ��]v�@TU+�m�\��+��R���<嚭�nԄ˳��������� �vM�٤�p�#l9"���'Uţ\���w[`�v��z�:���D�[��wq�e��sp9�-w1��[���.�M�R�6�{��[E��U�x�TT
�����`�tWfr>�xR�Z�'ctBa�Qw8�p����#UP m�1Y@� 
l �J��7ت �m�OT�6�@U ;��SN��Z�΅�c�\������6����	����U���r *�+�l*�,jʤ��-���J���S���h'ڟ~����fe�mmf^���d����GE<k�3���ح�܎g�zb��2OT>ͭ#�8�d��%c�������!Ԯ���w�n���z�l�&�z�D�I&B��_�j��;���o�����5���ڢ��ۤ���	i&�e��7k^�g���܏z��ߗ.U���V���v�F�H)
�N������8��mJdB��Mm��JR����*Id�v6:e�$�Y~�^;6g�{f^�\�-�{��#}��֪H��'J�a0����˅�=^׃����y��_xvwWw�Uf��������ڬ��Wi	-� C��f]6����=�cyڭ�Oz�r?�-�kٛ�I�f(S)��d��e���^�V�¹+^VW�s��G�%8o��A�&�F8��ɃEmLޮ�.~#f���;6hǷ;n�� ��z�4�pe�B�)v��9ݛ�<���OKյUThW�l7NEz��I��OW*ѳ�̬��kf���z;ǃٸ�o:��T֤rDJD�$&6K�.���S'kB���2���ݙ�_v��k����$��ơ=�u�l(��/jwEf!�b'�y�8��#^bmo�٦�u)۷Q��\�&�e��S+?#���YX�<��lڽޕ���M��r�N4�AGu�{��9m��V�ӷ�+f���l��R��7���f�`���0US�v�km��&��v�U	V^P�C ZP F�-����#��ܫ��|������8)7�ԕ��(l��qw�H�etp��1!��\9������f�w=�2��v��+����-��6�$6�I��7�	�����-Z��f^K���Փ�C��&��ӉI"P"��έ���~��X���;�׈��dlUz��UCImܽ����R�RF�P��!��;4��;�v���ڙY�fg�*���_��#�DFNgh���*;hsLjd$:���e�� q�=l���&�p	��� Y�%M��v·�<�y��| �ݪ��*�a��I�#%ĤI���2�����Cna/|g�+��
�跫����V���t[�E"M��d�&���fݜ�*��o�͚5��u������eb��m'	��d�y2����W��{���8�L�/m����Z�ffm�l;Gm�TNM�U�oe)�^�Z�r�n��mmf��cfm�Kk*���R&����E��o�y�u9�w��.��\j�|KB�M��Nl����v�
��;�x��ums��t{�+7���
�g���U8�e@%m"�uUJ�J� �q[�3��{`�j*��A[�i���Vznj��7�   ;�� �    wm���*����U�wUw �� xm��T�@
����]�s��9[�O�ծ9�<�2]���Y�u��]��*�en�ש��RF�jF�,���.��~��n�VUxl��zr���J�ڛ]��d%E@[���t=��\�2�v�Ӻ֎�6ee��n�ܕ�⡑�1"L��m_�fL�YY28�<�g7f���f�V��)��MB!��0�$�fmމjkÃEeL6�];9F�խ3l�ٻ�I������H�!I&z�;�`C�v��W�
�k���86ϵG/�����v�ܗkRv)�U��*˔	ڪ@�\u��}j�Wj�P�e�"@�5a��f�D�#n6�8��{;���ss.�l�;��e?�>>#{��=)�q(c���$�"��Y��j�Sk<�_���I�C���x�ԙկ��^vyн�Y��(\H���\0&N�8n˘��|4qg�$��d�.���M������l���"RI)�f�K{��#���Y��/vo�۵땷6^_pl�a4�)��a�:v��mePU�vc/լ��㙤�\͙b�&'�"A�'��Sv���	�����6��9�x`����2B x�=�0.��-t����U��y���6z9����fv��fdYS��6�nc0$�A�7�X��Q��^�����V'/��-�g�V�)Sa�$�FcQ��OiӓwY+h��۳Ց��������[͚6*�M���-����I"74嫡�~zv���+fu��ޗ��n,#�=�̘Kl�P�ErD�R���u7g�чG��m�U�Wy��b��4�~h�"eA"Ĭt��H�����l�r��׭޴Uw
�����*��$�v0d��)mU�N��G��M{c'v����T��?d��{"-��qB`��=������{-��zwh�{��n:���)l�#q&�g�(�/n����f���v���`+o6޾�Q7$�2Zq�c`4��Y��y1f����og�\�޽�]Rb�8��>��٭&R��@�,M�K�;�ｽ�p���36�a���f�iK<�q64��x���ˬ�Us���V���UpV�1K�)p=�h��m�s�V�,���i�d�ê{�63���v�̑%�Ĥh���w�۫G��M�s��A����.5���)�$ی��1��)�ۓv���7�rλ�����o��c�D$_�n%R;�=hf�=х����Os;R��5h��l	$�e��~Nw_k����3*��~�ٴ|��o��t�����*�+m��U��c��kv�1�5���IȘ:I(!J���j�%(AB���;��ܸ@x�%��m���Vق�nک�VPe�]���nX+7Wnݺ�)�� *Y@�܎��3�eM2OR�g`N3CnvƮ�#�#j��v  �� � � s{`U�*��U� *�b���*�<aY@�P�㺞���G`X��t�7RU$M����T�� ����G�UwVd�-�\��()) ��>�]W�]ϵ���oq��z�w���&'[��%���l���7,}�K<8��gzN�|h���o�Q�I ���I%�nMf�n����skkߖ�����s�k��H�
���7p^C�x�䴕�7����o���2��ٸ��#q$������{2ޟ<�'v��4{+d���n�����+��)d�q�]�H�7mK��!nv�vIcgp��@�Uw�UFB�-�.�y���rm^w��eF�/$��\���6�#��ㅰ��3l��Ԡ��2�Q�gp�5���aѕ�"Mq��c�C,�fH��I��{F��W���������_��rl��&Kz�mH8���|����l��9��&E��t�"I�9����Vy�e�wo�֝5��/{Ʈ�x�ဗ01
���8ܑN5��"�آ���vG����
��UYm.��Lv�'),�$!F�a^wϿX;�Ury����xwh�cs&��m�YND�h���ҏxny��e{���������#l�i�i275�~��ץ��w}���$T�'P��$6�$��if3h� 1�� �g�O��N�H��p�ɲ�>J�}3~>ڱ�x�0����Ԝ˧��ٮ��ԝ@��#�m�\IP��a�fQf�<�O��Z��C�q��d��1 �4�I��0�*�HVB�C�0�+̐�������	����2!<�i$�B���>v���T1 ��+1O�	�ȳ�I!�B)$�wa���y&!���BbM2	�&�T��,��R��Ǯ�O�C_RN&3�X���g��N:`c��m ��a01&2~HB,���	$4��J�ֽ��o���fx�V�H��dD�5�0���-QռY�[ a���ǈ��G
�\B#K��i�G�r�Q��qڑ �%R#�"��3�B���h�#H=7Mx��G:��>��w�2V�@��GJ&#�0.�H@5 ���磆�n�Uf@wn%UNc2��ԊH���Lݝ�4�<8[����{�Q#HDq�t��Fr8�!K�`��9�P�"&$�8Aq(�,�|G����Ň�s<��KSHs�5�7=kշw�
hс2�N�
7�/i���_�P�[4���7�慬Q{�}ͪM�j(ڑ"�sն��g���KZ����Q~L[�E�z��v}y��_��h(�\"���Q�p^=�(��@���>�[���ߋ�0i��L�l��Y%c=Rn���Av^�s
�d��R�]�U��I��UUAm�t�{ 7nʭ��
MǕ����5S}�����ϼ(�����;yy7S)�=rن(�og_0��ߪR̈́5�O��;/�V\�ɉ-e��)�$ѹ+f�����x��8��&��"�9ǫΉdf��&��CXl�<B��`�6}ղ����<�{pB6t�5x���!hû�:HQ�KFF���Q�$����P��D��{�D!��sL��!���w���4�]=�ǯ��6�}�{�o}�m��'A֍�S��Ѕ��pS���k��������� 
��hn��'wqT�4��b1��UH��@uU�U��*�B��Y�Sb�m�W�)mm� *��UV
\�(��J\�'Y���g٥�k
�j�[�ͷu߭�   �  T T ��m��6�lU �j���VѰ6�Tm��Y�Ae�m�N6{[������&H�R�����lR��LR��A��54����v~UWf"e��`�����~��8��r�L�6|F�*�~�"+rWg���İ��E�6xr�"04�jD����G��!������څ~"����l"T��#N]�G�����Q�II&�NP�i�ã���!$wo�")�0ӣ�v@�Y�DR4G�ϛܨ��j�!�)���Q~v~���ƌ#M���Da���:^*��XS�Y�:Bk�{�oR��
��!aK%MZ^bώ#Kf��",�t��%�#H��M����Gv[�C�(�� Ov���FVr=�zv�rU{kڻ�w4��_� P�ʵ�6�|�ga��+�̕D�����B;��
#N:>4_�(�!⋏�$ɳ�+�e
:��䕧8�!�$��U�ƺՒ�4�8�)��O�	۳W�#(ߩ��4F�]4����ޗ҆5�dSY�|~H0�n)08��"��>�e��Y�6|-�$qE��;�oL�G��P��F�w�M���2EA�31Q"j0"0��<�7d�pJ#C��DaV��O�4ȸN�T0�|h���rY����%$��:oMy�5�����|��������(�0�穌!�<F?l�4äY��w�bF N�M�������5\���d�]h�]©�Uݔ�2����j�#@����F�g�C5�3��Ȧ,"0�����D������;�e�#H��zہӉ$�A�%q�4u�40��D񴬐��#(+~���qx3F��#u
��.�LI����p��(�Ύ;�8��D�vm�Zl��w�B��0�2�&d�^W~Z�_��Xh3�T�T��;SWW��g�b���̻��4M?��a�j3���쯗�_&��(�a��)&�#����/��v�o�v��YFL]�K<Q�<F����Da���O)�YP6�n��� !C�U)Yڤ�a�gr���v�S� +�)��r�0�2��"�q�i��E�s��C:h����DiE�m�#�:0V���#L3��l���&�1�d?�T4�E��:qa�,��}(�FqW}�⎗D��N��5�n�+�������Z�C��V�p8�(1�.�
:��=U�͎#y�fi��o�q�{=�K%����,���`�<`[�<�<B#T�S�c����:8��Dq;��J�A��Awi�6W�$�����ee"�td� �y�#�;�0i�8��+}8�0���׵bH�,�f�B#���+DI����b��#5n�d��jtr*��:J���R&�@��UU���֕�åر2MMY�y�~�$(���g��,�&��"j9D#Z���Y��s5*��ZF�	#wN��i��6������J��:E��}�8�#���H�˵/)��}TGT��7��W R�)#��kL#��<8W�\Q�kg�R���A#�U"8��0���GG�'-��Iڭ>>#y�ii��)Ɨ�[���7#�/"���D�N�VSP(�8g�0gbȖ��nE�)��G�|E�-�_��\>8x3fx�D"(��"(��[�粽x��.w���E	IA����A7����S����v6�SZ�f�;��:�\�ea�WsJ��f쓶�����}�|�m�������']�9��=qw}���벮����`U �gf,㮿WM��kr$�굳J�b:���1f���   ¨ �    ��s�6ø �����mTP�l;�lw)T��^��Z5�ge'v��OR��M��9YU�2�p;�w)�P��O�����U[j�o^f�Uyu���(���dx��4�4��7|l�4s��~��i���/鸚�",��3���E���d�Rv�(ڑ�%
�a|���=���+j,qa<���O�}��dN^�a{�U��m�
Bbf�$E
���E٬ٰ��*�j8Ւ�p�Iu-�.G��4g�Dq���I�%I��1H�"��ó��B�Y��g.���m�����(��I`����Eԙ�hU
�$%��>4~"͜��#CH�7�|n���CB�#��#Kf��B���S��f&�>�"T��#�P�J�F�q%��Fnفt�*��U���t��w�x��C�S��@��{k�i⸰�d�!�[��6E\G�b�#ɲ8mvJt��<=8��%���F���!O]M�0ɛ�-��U{��F��u�!� !3dx�-�g5�N5�2q�rfۈ`B4�Z�]�ڡ�22��^�?v�dG���k����8F��B,���@�g������brXr9K����Vg}�%�]=L���b�T� ��\��ap9��}�ٓo�Y��ڬ)�I#9(:@C�����<y'Z���'L�'�tS�!��U�F��,�TR�rRa�B�ՌT��T��f�l�-�fU���d�l�Y�p�S���J@Y*K�Ta����r���ޫ)yW��[Ȟ��r�@���D2�g7 V��m�e�����^ko�g-͒�[��ˉ���8�(K
��$3mKg=�a*���~ɳ��e�e}!*H�"�Q#�Gi#��d��"��0��i���:k7}���O]k#DWuM�!�#��wgs�Y���#`��[i$	$�ƨ�Ϧ�������G�S����s�C4Y��{�Ƴ��H"�Gg{�\�ա$�ȓ�������k}��~�0�p4��f|Q!�!L*N��1�ۓ>j8�EKk#r�H;T����w��뽍o9�Y]���U�T۹��FZn7qK�E�)q��B6QBE^�����A��Ƥ2�"���N�g�R��"�6�@��Q�Q��!��"8,4��F�"ݷ�%��S�%$gt����f�dY	o1�vB��@�� ��Z��<Ԯ8Y�+����,�َ
�Ւ�/�<C�����!�m�JAR8�m1j�Ѝ��7{>���"�0�-��0�DYe���b��P�Q����0յ��־w{k��Y�M��((�8�MUXDQ�9ɵvYd%J2��~�(�O-�#HE�G���$wF��Yp��v�6B�ȫ�J瑁bX��6]��g�ҭJ�J������L�sP�(R��-Ԣ>0��;��P��`��9 ��N�{�*Ӥx��T��w�o!�WW���l@f6�!5^��K6x0�E�!Pt�=�nb�	��\(��e��M�ٴ7-��>Q0LQh���K��&�og�n��dbR<B����:l�����k^�����"���~�$#��55h}������F�oJ�,��?qs�p5T��4�#����P�#��mB�.S#�;��8Y�ay}8W�+yȢ�ʲv��:�E��2���i��Y��E��![��� 4��'�X@��:�q�W�Cbd����Z���` =�O~ᕇ�$�iR�������{�M���5�l
�`T� ��q��i&�$�u$��<�6���ڷ6���ԝC��9�����N0	���j~v�ɧ߯�`�ì
�4È@�C���~���O�_���'a�Hn���'��O$0�f!��$��/�'�
����ݺ`����_�̆�@`@<��6�Cﵮ�˭kY�k(' `��{wl� ^�	�i��[�T ���@�quG=t���ְ�׫���]���Ok:+x763��α�6����{v�����9�`�Nm�u��}{�۰��le��ے��u^��^[:s�!Wn���r;;S����ܝ��=�Wk2WG^.ź�z�{���� � 
�  ���[ ]�mZe�+(U U�z�rP.ܿ2�2�`*�EP[ *�^�@�������_^��R�0�@ x8��T�[�\I� �UԹnK�_<�F�v��ɶ*9�U �lxx�Tf�wF3��<�mu�g����DeP=�����@U������-�6@ UU
�T*�Gn�U�[.�6%� ������;J  � ��j�T�e�T��ʴ;�*��� 婽��T�m ���uP��     ��  ��
�  �l�J��uf�VK���&A���-UecHM���y{�+1N��\��\�q�I�¸N%���\3�ʛn�L��ӵ�4/��H	nIh`.��I唱M�L-XFZ�t�11��q�8��Z�5��a�3ʕ��D���D�˺rz���[M˸�T3�      �   �� 
� *� 7  *�@ 
�      �Uk���     � T U � � *�T   QT��ܴ   6   �    .`   � �@      m�`  +(     ��YZ�x��}�n���p  +��P Y�m�W�   �  ^   UU��+�s*�@���+2�* UV� �����)W���r�?T�բ�̅m����{����*�����}�P�gY�F~���mUr��ج�i�8�7)���M�Y�?|}���|FKd)j����p�w�Q�ت��<-�����~��؀i��;wV�6��߇��VR�����U    �gZ��P�l�sF�N�t��Wd� �r!��UR�@� � ��۝	��Q�  � �`� 
�J�FØTЮ��X�vn/N�B-��G�����ր��'F�q���:6B�0�*� -�)1�v<7v�q����Hqxi��~#ŋu�"���r�.Ϻ
��o��E3�"�<�}A�䀠ZN�d0���#��+�xl��;���F��Y|���$��Ԡ�����1�����$�P)��a�⍕�m�G���|,��p(�'��$�QH�l��0�S��r{J�F�de�����k�EH�B��b�DaA3�"�S�K�6�߷�s��}�-Ÿ�%UUU$�;یp�؟k�K��Q9֞��������w�s���Å�1Ɣ,�x�H;UTq�
��u�*�*�-�8UJ��$���&�)i��$���{����,��g�ȋ���w�cx����,.~����%Z`HFJ�AFR�4w�rz�7P"o}7f��vT�/h���K�+��ۗ��]��&�P#qH�H��۬�
���	��{r�l}
5Nu+�R}Uͽ�Qg͂�MģqFܟT��2�kr�2�c{;��O}M��bϛ�W���Ѵ�����CLN�_��~~쫿g��*v���s���J���;�~���TA�hk��v+B��]C��ݖ�v�����Y��Y��z��J6ل��y{]��~�W�}+Y�?y����>&���\�o��<���H�K�SU3Fbb"�UUWΝ�yn�s���ŕ�|�/f7����~���s��0'TH��US ��]���0���f�m��<����ʉ�<�8wmǖ;��T�vz<�(�(U@�@mֽ�=�e2/ܡ����~����xzs���S�}���ߊ�Z2�%�K9��wzFt��QGu����(柩M#�yq�}�t���^���+���KA�Am���c8��j���lx��Z�J�d[kd��P���6��T	F�)v�ƽ�iF��<m��0�,*N�,���̈́Fl��}pY$�2,��{�53L�$I6�E��Ha�$o3Mb���^*�Q��N���҈m���8�MʳG_���� UȬ� I"��ہ�3���8�E��7�DHq���5����##��"¹n����~�[��K�m�����6H�%(|P���DYB|:k�G|��>��q>\+�x�ӳC���a��Q��G�!-��#*�Ər~,s�U�yv6X��<C4p������0���1U��n��.�S�j���tZ{#]A�/ n��d�ՅWp���J�+��u"�(8m�R�EAG�4��A~�n<|C:_��C"J��7��=�di+_�Y��d�q[�$���Y�kmd�y��'CN�l��.����x�����F�4�U��mj� �LD�D��"�MM�!�#����5YC
��Ѭ��U"4�ux�GT��&�Z^rk���|bq�T��D�t5��zH�H�K�l�F��ٸnF�͕����u�C��f�w��!�<Y�_|�)(�a��m���n��#�ȶ|t�8�ðm��:p�"��(���0���De�{�)	����'����j�F�٥Z@x����s�n�t�������vm�f�q�� *�m�sk�<�;�(����m�(G}_C����i�ж%�*��v���U�շ����W��0 ʠj��gZ��QV�9����S[��<ku�KZ�BPT<
���   ���*�l6� m���ն�� ��+��$dt��-�[mԑ�<��;d�K���;[&F�W*�Ŕ& 9X�<i�X*����EV�ʕl��U�7%�
>�!�<f�f�����ͲB4L�t4��t�66IcjQ!�<�D����h�$(��G_"����8~���!�C�^4B(�\61ŷ|C<_��{��2�����Ͼoq�XR&�VeU]̖E��c���:Sq�ȳ�!�B��E�Fl#�"6���F��B��F��-eiА��~|k��q�`q6�Q��M�Fo#š��{a��n�V��HD;�v�@������*bk����a�;�"|��IuD3��5��4B>8P�oջ̷��a>}��G���A���m�ܳ�M����ޯW���U�<*��J��%Mi歇3��'p�����;$#.Cz�e�DiMG��/�ä́]vg�o
#H�P���A�8�Q�iC�X���W�_��UC��ؽ�YX��w�(��\g6l#�O��}pt����5{��mB�	��)5��y����zךE*1D�E��YHnU��*�3��5��g{�\@�#e��$�l�bj��C���HdIҔZ���#HoU��*}^<���2,�l�}�jC,�!%��)�(a~�w�}����!f�W�X�Q����7�t4�|tߑ�?����+�D�gq��Kj�U�Tiw;�)�Z++�T�6@��T�)�������I��K��&j�j"�aSھ>���iA��|Y��9�!면QF��Q����iy��9Z�%	 ��=���Z~�[�n%��@C��:{�*��S���Ǖh�f����}Ѱ$ET
�F&�I#��Qa˜�]�X�,��٩L�yD3G��Ԩ�J��0��Ï�B2�FP2��d5*o�I�5-��q(��"ΥV�p��Dq�Y�-�������X��lC����}2�#�NKib��f���8��5{�1J���������-z��u"�b��~x߻�5��Ήs]pp�� ��U{z� �U�J�UZ`[{�<�v;E-�v�!JJў���N�9������vf{��=��oa�SO�D��I��m"߻��d>j�P�{�$f��k�C!z.��6z&�qG���k��糘ݪ�%$-���v8�E�+��Gu���x��<��(CQ�.$2%�<�n3(�$���q��7*���;k�+�.��	۞�E����8�p{��ݸ�kI�U�E{=vG=�'HU�L��(%1�Т0�pp��P�i�]���c����.8���IE�!�������\|�M�=$	��0�HQZ��څ��`*���1׫v .eU� w����(�?0+�XZF���Zkχ���T4�"�`���4wP���
�~,�]����\߾m�aڑ1Q��XdQ�Z���B#K�U�{��"̺s�@���4�1a0���b%��,m���ں~P<C�Hd"$�1��"ρ{��M���)_���u"������Fو�L�$�h�5ha�5�i'�����t8�V�t�Q�����f��G<�e�T��)B@j�P�d\iw�Gh�G�2�`��]���8D��\x���>�E=�~��p��Z��K��-��m�   5,����n^^��9ӻv"��?KݫX��N�pӲx;]��:����3��k���cF�&�n�p,�+++�����N���6QR�   #��Ӗ�β��24�j%
Q�E����kk���_ �p  -� �*� ����6ûl
�6�r��� ���^V{%���n��n��鄍�[\�@/(�y�PU�/;�p�|�ϻ���z̄�!UY0q�&ݖ����K�ܴ}��Gȷ�Dt���dN)���(�<���1G�;j�GZ��$9�T��lԪDx�x�Dw��m�HiT��\Ydx�R[�ņx�xu$q�Z��ӽ�^P@[q�")đ-�X�8�=��u|�idx�[���"U��+�!��th��Aܲ��2�����H6ۊFڂ8�i��·qw�����#N9\η�p���K����h�r}�M��+��G�(�,��t<E�5ho»)4�m���uƲ�����!%�LXDab�8��;��l����:��RG\�m��Xs���j�HN�*�UJ���T�cd'28Wl�����]z��ھx�F}�FOG�ļu���[�w�<z�w{�T?��F}�,F
I@�ȒQIV����{-�w��b;..�@��m�5��Gś�fy�@���ǌ=�a-�{�����j�&�q"���Q�E�X�0��C)�}p@p�Q*{V}p<~ತW(�/b��:Z�+#�RM�����zް�`ͬ�D�w�p��A����]����ͭ���>��!P��R����8��M˯j�.|V��L�43�|�RΏuc5��bgje�Cvd��h
���\LrvɮتUڥb��8�T{���z�Rf2f$�{X�|5{nffߧ�%Oi���Ń]\5���R�,�	�	F�(��	Eb�+*��CB�괫c�y&�}�;����_ـ��P��1C$��Tz7�m5�˧AD5������O~������3Y:����P]�&�k{�!�HN�6�$�%Ba$�+ �`�	'�'Rj�	!ē�HH�O���ܒ䄟!$���!Pc�* ̀�$'�h|���@6�4��$��@�~��!� ��BT����}���d5�{���t!���Ht���M�0����@0�O2I'R@<����Adq�$�`O3�$�'Ύ~�L7:ʁ$Y	��BIY q �!~B�H~d��|�� TH����<�dhI6ì>d
�?!	1��Hu �R��L�6��ϒm�'�N$1�0	�����C�Bq	��Y:��LAx��m������@�}��K(꾔mE����Z�����7X[F�CI$c���;�PY�t!���B�N��������EGq��,��Bj�BH�"RrV��li:>���J�[�װ9vEfF�x�l?M|͟=��z�v�6Q'8p>~($�����ڍ8�׻^�\'����Wn��ƀw
��d��.L�K�sv��*��k�:t�8g��S`I�!s{tC4Qt�Ұݡ��熼@���x�� [���D�%�"ύ�E��ݾ��~>"����1e:�ݓ웹�������A��Z�WM5�L׎Ǟ����vB���t�^�z�[E�j�u[��1A;hH xo���ufl�'y��&i����&��]�zm�je�٫�>[���9�{�uT�H	$������� ��7��ө��� ���Ջ<��{~���&�gSm�+h`PB�UBn*����a�>j�{���*���n��QV�B��$�΁�{�ѝZ�jf�~���uJ��(�<lφ�4������G��(�e��IIm��hR]�ǧ氆�-6�}wD4,%�#�g����fO�	;ˢ�s[FbLf蚪JI�I+��1�N~5� ;J�З{V���L��b>p4��'O�z�Id�%(�I"E\C#�º�U�~���\);����t��yQs�і>7�|@�"w�Im�U��J6ل䡄Q�g�Z���"͟q��h�� �~�G�HG
ӊ輾������bT��%%!I$I����ދ����y��9ls�Z����(�UR�@A4B켠:����n��׵�j��h�l�g�23*� �R�*�v�㾗���-�� )IUhr[nt�@';Uy$<�Ȗ@���s�ͭv���/w/#��l�  �  U 
�P �Pw�Cl  eP���r�uSn�*�P�K2vUZVvkZƙ:�S�K�qx���c�u�&��2��N�<K�Ɖ��^	U��&UU�� 쬬�]U�Ə�߷*��F�Nt�8)�a�����W�<E����#$(Ga���GGÓ�yC��v�X��W�R;Z�����U&��������<���KQ����]�|p��'�Վ8p���6}�gn����RF�ڙ�����,�:]���fh��)&�v7�S�w�﨑��]_���;s�h��FD�ڿ?5�^�wy�
Q�!i%�j1�_��%���B�A U���$�<�-��0��7�Dw+<Y���A?(��:-�sٸ�����ZjݗWz~��y��*��Oc 6�mw��5���8��I+�#N��A�m��Wb�E�J>-�F���Da��[�l�?���P�AJ��hk�m��=��5����>'~��yd��z�g`�,wV��A�<yӟE��BȆ���l��-���:M�5�ק�kv�2�QDZ㧣'�>tJȃD)\w|�ᆎN��S�H�d��%U"��>�!��2Y�,�gn*�>|+�`�|h�����:p���L0WIb	���!8kƈ����ZQ�4�����Pt��]j�e(��ۭ�:G5�s��[4G���ж�u*��E@UQ�ccV˸U<UwQ����t�W�R�
=�K����L�x�BgN+\D�F������`���:O�|���p(�mB#V�p��LYG�%���d�>:x3{z4�<n��-Urx�<h�L�H�!-$�p��:��y���@�\87��Fzjv#eϞMV��:!�(:|Fou�#L?r����Ӑd,vH@5��8��'Ϲ���Ɨrl�^Ŏ#=�27��`�Hr�:���ޫRI/�$��&��k�ܻ��?��E:v6��|�Y>/�֘s���^5�ܻ�,#��M��Q�[�v��u�X%	�꧂�^nѶ���	+�+�	*��d)��)��?���ƆC�U�f���ר�%0;o�{�J^5�v��m��ڟ�p�5UT�}7����7��Ǯ��^M���#/�v1vF{��Y��Ӓ"CL��0uzf��)�fddҩ�n���\e�_+j�Ֆ�&��BF�׻:���>�zn�\~B�꾜�y^7Z����'p��^6��d�^�b���%�h��G�A�ƑԭY#��?a�ŕx^��<y��E���p�=�F6[@��A��^���f��q�S���=gv첻�� �S��`Vֽw�ol�{!��FB��qGH����%��H�8���D�3?]G��'pC7�FO�o6r��hH�ԡ�:�X��Տ���<&�U�G�ᐨYG�{h��˫��9/}ܔ-�� Km�Sh�g�+�Nk�3ǈ]I؂%E��?q)���6~DaI��_���i�Jq6Km
q��9�>�n������'�+c�
&� �#�S��T����'�*��  [I&�Wb�g��g-�b4~�5F!n<j�(K�W�"O��t0����F�e�K��QH˨��%�"D�$�&���K��s���[u�k�\�q]�z5V��IhH	vy2-[jv
��\wx;������ܻ�u�6�Xm��z��Ԫ��ͺ�� Y챀  �������w���
F����[:����[=t�}�Ww��@ Px �`    ��;�Tc� *��ՕgZ�V�PÕ��.�D'�%%kc�7 ���ѫ&^��oP@�8�uuv�T��uU\�URZ� 6I.w���T�	�+M��a�h1��c�#: �ʔ�?A��~Yb���g�֮���}�x���Oa?Z�!d�+���8�5��&f���g����w�0Q�ȅfqB \Ǔ}��憺��o�K&���Z�4���Zv ��Ҧ>D�Of��1�gY��� i�FN�_��k�yZi4*�M�$�����	���<Vl� P,xvM=�W�"N�g��ԟ��t���F�p��x4�,ӈ���)�JÇ���l�<~&��U��0��i�_e��..?��wߜ���E�=ϒL�٬�K���Q,�M��Q8�kM��M��Cm�*�������s��˕��	���dq��i�ό#,L���f�Y�O�qJl������Z@�)b3dn����1� ��1�� �V���7�r�:Nd�4~�E-6�0�g��\E����+�|�Qw��\Dl�5 �ܒJT���=Q���>��6F���{c?\uR���M��̎'!2'e~�#�~�:��4�M��$b���F����G�#�L�zf�AƏ|�pS�+�?��])��'L��nH�6+Haѳ�W�i:l��d:��(��?
Zm Q�����~�������q�˳u2�(��;e�P;���wk�E� �=M�;�U^��6�T%$,8�ȱk�����^�s��{4v�~�6���0;�����	c�QTiAnD�iBs;Ӡ�\<}ަ3��6�ŧnӇ�;��6oPDq������M��v�H�к������R�6i�����F�+�+�4b'$����8j�ï��n �"~8�^��l����-��hHG�?�k���?ZɠA��!5n�!�(�����zt����3�}d�����IM��N4�I6%�+�gA��u���:Q�R�?�Y�����diÙi�ό?1}���w�uA�`$��E�(!E����s����^˸ִ���N��;��i�J"d�hJ��j��4|�Ҵ��H�X8�����ozW��,鳶-x_?=�'�5�����-��H�IcQ4m�0��r8q:����� ��[���'�'-u��t|��p��|�"g��e�#fd����6�Z�u}��1{��7%�8j�w��2`��ڣ>�bU�:��冐r�֎΂���{.�����,Cx6�s8l�u�tʍ�N%dD��ֺ{G�����o;�~��|/��մ��O,\�jm�R*O%��nX;v"!�IS-���e�|��hU*�Hm&Xͭ���ضJ�������j�+�e�'�=ؑ2��w�鶑�+��u�R�z�6�CA�m�(�e�`y���~̥S��u�U���'ZpyRZ���SUQ5UBDȚ� ��^������P��v��[��H��r;�J�3�n|LH�,U.2���BnJ����OP�������-����O\oM�v��;QS$� �cl�2�h�r�A�&�K{�x}9X����m��գ�K�u|����=�R��O&��j��|��P�*���Y�Xx_�9e{4ՏH&�i&�e�Ԭ]~���>��d:�p�"Ʊ�7u*���UK��uQ1�6*i��}N�	�� =���Y��V�T����T  ʯf�0��^]�=�Ӝ����c�]�Xa���l��#�a�rD�T��Ŋ$|&���'�w;���
��T{:945�Y�!) ˼3�u����o(�unj�.���h�EsnZ��V히18� <f�k���.���T   T;�QT
�u�{v�q��V2  *�]��e��7yeT U pU  �Psǎ¦�;:�u9vk�U8   �{�'V��n�3Ǐ��]iB�%�yVX9cmV�UTZ�P�b�t(��=E�y�	0���h�v���� U ݶ �UY��B�����P�fUE�PTP��l�� ��^�q�=��6U  �ں��J إS�k�dz�' cT�� ©8m��S͉�Y��d   	�   U  �P  �P[ �    �*U���mꉬʒ�
Me&��up�VR�[+~���g�7�͢�u4�;9|����"2k�h�����=�q1KIq�.��v ��eԯm�UZw5��!B�(΄� i���[b��ܻ<�f���+h6�x�KFV�ҵm�͖R�ؖ�e�v�vV�   @     � 
�   �   X�        6�T��R�P       �UB�*P    � �͕l�    �   �    N   � b�  � �@��  ���   Skez�m�Y:�r���  �x 
� �@*�Ue      U� � ��l�Y�k!J�`cUP�����҅Sl-����TS�%�YA�v��8����ȯ5m��*���9���km�UU[Ӕ�Prstd�7m�J6θ�1P!-Us�)Tm��iI+�K�x��ٌj��n��p����U[ ]�"0lM�wt�f��!����/Lw-S�J��)y���e6�9݆��Yس�v*�V� w
�  U �U 6��P*��M�[h.f�nmTT��)�wP ���c����'��,�9�2**u+�5R�D
V8��l�8Z�viV�� ���z]��[�D�Ѩ�"�T/��xKn�u����͞:F����x��G�+��#M�*�#VV7hHI?�I�:�wٚ��_IG��I���x�><��_�}{����!���Y���D-a%��1�M~�G�!d#��x@���~�{5�`��aguF�D�Ow�z7$0�d-���2�u�J0掵f���0�sz�x�Q�42(�P ���6� Q>�o9K	i$�Gb�[\Mi����"� O����K�(��dI���W]q����\��$WL%o�m%���Fa���%If����÷{�Uw
��j����kT�F�2�ca�>�fp��#s3�`�Dqv�� �>tH��Gە�-��SA(�b����6EU݉#:#L|�og1�#6T�CwS��B8<iE|3�QC����Y�C�����@Q��A�>�F܆G		�k�g����� �(��g�ܠ�DQ$� ��պ���	*��j�~��@7�}�K	��^�~�Zh�͚w�0/�#���>Tz�dg,?}؇��#I�	M7 ΑGD�v$�8Y�f'�Og���
�?�a����i��V��־d(p&�&a�@��]T�mm�u͖-�
�v�U	RX� �C�[n�����֢�{�~6���r(
,tx៧�m�������QY�M����$H�q$�NK� i:>��Pb/�kW�M}V��0�"^_��H�q8t�F|}㑢������V�̌6{g@�`�Jđ�{</t�����֝Μ�@E��Q�q�wql&�ViF�0�SW�G�d�a��l�g����Dk#��C���ζ N����n������]E�ؒ4�@�����G��v�V�q��&��B#
!2%���;����������A4�C A��[#�^��u�{�@;�OSd0Vڪߨ6		!lH�i�����C?���}��Dh����	�x7έ�J'���R9Ki��_��w��J��!�3&�F�"�4@�)�����ï�!�!������m��_���YG����@?(�ޕ��C8���3D)���ŷW���>tꉚ��%9��B"9P�,��Pj�vx���VP���ۻ�i+ >��۵�A=�;}�u绘3�b(I T�~^�.�S�>�0�hM$*B��[�{�M���!
�`[@B�t���W���l��v�\*]�d�[] V�w��ZIC��$�t�����������{���������[���"�=�LE#f2IN$�L0���ŗ����1���/a8�������^̭�(�⤎Q1Uv*��M� �5:9���Fc�x��n�k�}^���6
gࡒFKr D�4�yu���7�k)n�X*�9��Ӌ�{SѫHP���k�1��\n�Bũ22߫@V6�Ώ"um���f�˺��<^��/$����j���=�-�®tk8nE��s��u�]�FB�˲��p����Ԙw<���[�n���9��P���Zڻ��wR��z�J�� E��k��ݕ���Ξ!�y���T��N/7 ���D�'UP  <
�  � VڀWP�w�6ùTUM� �[�b�� <aYJ���P�YW��붽t�����pC�9$�*�we��n�췵�
�઄ԣ��k׵3���-�RS���{]Aқ۽9�D�:{w������be'��DwL^�T�7��$��і�M��!Pv��$i�y_i��3�T���������Fψ�S��I�NhA�X���A#~�� O��F}>Sq#�k�0�H6�I&�L?����yي���G�������F\|�˄�E�����}�<� JU���(�m�5��E!���G�>���f��
?*AȭJ~æ�cM�����{:[��2H5E���\��n�� ;�s��\�=�P;�S�d��UTc���8|�����v	�p��7�ߌ�|�����Yڎ�[�Wd" �"�]�����J&���h8V[��k�G�d�g��S�n�+�V��VAF�"OȺ��K�#�ga7�g�b���<}�������pH� ��������+�4w�	�P~����F�6��g�d���4��"�]����r�����VXG��A�)�z�{U��r�F�,MW�*�Ã�K��ZGs�e��#2�m���s9���Ji��t�К�+W�F��c�QQW�-v$�=��
Џ���%aWT��m()2���:�ׯVf�UxT��Ujl���4��18�-Ȕ����������>�b��Go_�DF��!�PQyD��:��K#K#7�(Ԏ0�fH�m�4jE�Yg���)�g�}�CŮ�")ua$Q	�wƦ>DY���XS8~���}`��2ѻl�'(?�h�7�8H�G�>�d�77�����RrkG�D�M'"�GJF�����t5��(D8ے�� �Pu*�#u���0��߭���ev��~u7Sq����G�vs�|׽�r�Z�R�$JTlo�
?$M��q��_��t���d+�V	e�BN�񋏸��O1��^���)v�����{ M�`��U3��ڊ���+D�� On;Rp�"R)�i{���`��=K���}K��u2i��|DFcdƓ�F�q:����>����'���>#Q|���|��a��#f�u��\\�ɶ�95l�[Dܥ�5%��ݳ����fߢ~H=�Z���"Ҥ�t���Պ!�"���\11-�
Y]��KaMu����ooٯ.�Q����KwQ"0�9��6O�w����^+�=;����BH��Mi`�?C��EIn�6�&Gw���F�:������z�<�?X�FFM��b9q�4p�c֠������;"�L �����4ݩѺN%��V��z�8���?X�Nz��HJ����gPJ�ݖ���6Y�¨?Q�G�h��m����\ӆ��#��c*~�b���&	�I$�ܕA��(Q�{����p�~
��?I��F|�˄Bf^͓��Z���k�2�ڡJ���'���%�յ?a�ź����v�|ͯX�}{��9WƼ;=�p~�6\�m�C-����ݽ��u��?�I�mX(�3��ҏ��:j�Ȉ�S	�"&��5a����]�v$�y~������Rw[�Q$Q��5",���4����L�sN�p�ۂ$���+.,"svx8��\�\�W]=\=��ӖU�S�n�L�m�T�Z���e�ݚW0v����V�b�U̬gX-���m�( ��� AY��㻺ӎ�jܻ�q��f�p>�U@
.L[qET�  �  ��  �  m���
��� 6�ڨ.�%�ͻ�fm��R� �ܩV2N,��.�Cq)��Qi	;B6+����L����T��J��[-u �V=״��ZF4�����#��Y����B<W5�>���z��쬩?#y���G���}�����$��X�k�de����h\�?A�kU���Ŗ�ؚDQ���x�wƾ�
<B;�z�ĉ�jf�*�&�_(�G:8]�~F���!8��`�x������7���u�����d(ӣ$QQ���V�(����=ybS4u䟠�)�HR��>!&jշ?Y�Mt'q�J����x���E��L�
UP}n���8���3��lUF��$.��u��f�~�X8�'���P�FU\³���Ny�UT���Uj�Б���	�I(� ���ͧ�����繇�����(�����5nI�	�{~���?c[y��9+�n��b(�����%�Q"��-�p}|	��"�����?K��~�y4���31�K����i����g��rFFRGlm�ic���g�[�YGf6`�[�����2l:�5�(��z'�b�*�DYDJ�bX���(܍Yu6ާ{���y���6�J�B2 <�ħ�#��u��g�o��{b�N,��z�.j��D�M2څ����5�����|~G��=7�_�F8d0�)ܟ�t}�y,qh����7T�j��R�b�(��D�a�T���ݕIj����@��v����V:+-���]g�᯻:��i��J@����㇈�-���"'r>Do�?�3_��>��I "F�j��4���d:�.w�Lt}���{��f��Q��ޏ6��g�qD�jL��-,��d�ZC^c����w~�{6obHDx�&����B0�o�Y������]����׷^�f�vZ�n�~��J������3���9u7K����V��.�ZȽB���u)��<����<��K�ݞ�ڸ<#��3rf�[�#5y�a�/:�?aGųOf����r���[��3�� aiaw�Ƽ�M?cy�w!�#He�f����P�B�X��&���I�B������&X5"��	��f�!LaB�qF�E�P �C�#\a�x�&�M��D\�Xa����!?�n���~p���dl��,RԦyM�k��z��ӽT
�
�m�@�Umz�jl��nRK���οY��_��ز�����U���[��7��q�&����#D�	��m�I(��;����9Կq���8ڟ��Qn�+�#��f׬AҊ����x�1�R� !�㯹z��8p��<k�C4{�	6��r��c#.y�}�!�~/G̋<��&�f�"�rD�m�����H�RY�6z!jg`7�(�h�{aK󫬊��&�w�� Q�n2o�VT�Zwy�D��2���V�7�nP����"�z�6HF\r��{R�g�E��=sIG�YG�9����G=��`�b�`�� �f���k<hT� �������-*�P�e� �:�~~���R��f�؂�?Y�_�6�2#�Fz#�d3%<%�im"��KC�+w=���k9�%�v8JH$V��6B"ʴ!�J>������t2��X������]Z3��#��`��5S�	��Mˡ�dq�ѣ����Y�7�S�4�r�k���玴4��v����k�ׯ{���V�$ %��C�[�>�`�͛:`�9�U��#�J�ƾg6��
Z�U�Ȳȗ�������@���Q�=d����OY��5��!���7�J��+7�)�u��;��7-��.{���� i�tͬ8�� ۲ڙv[\��z��컹 xn�ǥwPx-���r�@wdUԲ���F�&�w[v�̀m���3sY��[�C]�q�W��N UUUJf�՜ׂW��0>i� e5ql�2{۽�`EJ��T � T ����Gp EUPծ�TU `��Txxv����s�+�\�jq����n�d�T&�\�nٹ纴*�k2ƩU+Z�Z���B�m��)(|]fc���Ϥ�Q��I����<h���$3%j�0���4�Gl�_u�
)��	��
Si�d#�\m�"�P�B�X�6~�涯�\}�a���Pu��D~�q�U�B�����������x\:���i[t��0����G�t���4�2 ��RߜǦ"&$��܎QuUBڨ��x�ݗ���&F�⛳5�I���F|���yp�}��x����A�B�)Ib)�8��"2^M7Y�E{�����^�/ ;=b�N4�fJE�M�����y����[��"��K5���P]mU1q�� �MJ�§�[*�@�]uG[q���m�	��Ǝ����g�x���wf9�)O�C���mׅ��#H��#��N~�E�7��"*fjf`,8�&@�KXz��2/���@�-f�?�s�|#r>D{rxf�����M~�Y���]��xݮ��X��S��Y�[��ae����N|�r�G={��mF��p<�b��`�{��~0�VZ�]y�S�^r7�ӷ4�?#��u�EgȌ(�Hd:�p��_5�k:����${��-$r0vM�MM򏬄p�G�����ȼ��N�͐���ӷ���Θ��"�p�~��d�LR�0�0�EX�.��w�ڵ��ې�p��UCۻjw{^!%�Q���C_����ױ�������4S�M#���KS��r0��&Na8$>��>����WA�Y����Qe�?���>�l}�{c�Ɖ��x�"&�����Ca�Ӆ�L8�����-$�5H�$+hR�X�bC^�ړ�9�,5��<���iW������Ou��a��d�DU���&�L�+^#�̪~]&l��sI^;|s��<��/s�7��".L��SPI��W��8���!�l^r%��u�Xu41����_#<	��� �����f�H�8�@������e&��j��&��ĩ��	�<�QP"'aޥ�����u��=�<�)���[+c|����zĻu�m�r"(3�m��F��{�f^�0f�Q���^L���t���M�(!ٳ�[�;�`;-$�23L�v�����G�wݹ����:�$nvz�GgA[�6q�i�v�l�Pmd�W_h���}|�����C�V�e/H��G�Y[�=��Y�<�/��n����L;�5nB�x��ؗn��Ŕ�g���&X��W��H�~5�bf�Ε<�E`�ّ��^����n.�������6c�"��R��T� T��\�vw9��Vj�bd��߆6��V��r/zżult��o��u��8$��)@���}��BG����!������]e��0�"�u���@���;��_XH����M�B:e�ח�	����u��o��'��,l^Dx넉��+�>+�dv{�eH�8Km�
3U6H�Ŕ�O�"'L�G�F�ɥ5�s$Y*D��ǍqDg�h�_��n=�,��<~{q�ٿ�Q�Q����9Ak�.>E0��A@dC����Q"0����l�i�t�z�����o��Lws�N��?I q��$��Jv�݀�xAon�(�n���mf�.채YX%jU_-5�sp�d'5U��n��`�[& �`M��)Y�X���d�V� �l���J� *��Z�9�e@�q��O.��]����լ���Om�V�;q�@Ud*� m� 
��m탸6��`  �*��/j#l*������̪�ĻQ��Ge�{ee�l�-Ȑ.Q�n���U]T�J�݉Eev�U�iP�ȐJC:i�[4��&j{\}�#��QA.^�-���6r�ኄ|`��j�;�~%�1���~m髓$��V0n�Ѻ��P��Dn�:S;nl�̔��"V(�2�"0�J��N>�e��4�
"��r���BJY�i!tǭkJ��O�Xȧ�|r��#��W��2ϲ1[�1y�#&�w�H�:���dG8��s��,��I!"I}��q���zi���,i���U�ߞآ��#���Ze��G�oaAՄ�f�A"�b����>8Wp+�.�q�X_,;6��:v"��?x��B�bEB�d�w_|�YZ�����r��N	Y�x�崳:�w��=.��w��d��%e3����2Z������Q܁�mz����a�÷��\a���7P+���"0����i�����",׽�G�"۠��K��=<���'q{V��G�U]Y9vf���4�MY��!�,Y�Q΄O�bM�x����u�cJI%���������a�E�)dE�7�c�<�\X��C9o����}�H��.���a%1	r6ъ(�y~�:�<=ִϏ�>*�Ǔ��F)��"��ʊ��U�9��ǵO��;Vc}�|Ka�"JH[Ge�s_���{y幄k�6�'�阳�bٲ<B�H����!��;��~�����<�J�(�]D���iIv^�h�N6�3u�مW��EwPJ��f��ɝ���W�v����|F\
�^�kc�F�56#M�C,�M=��#�̎6Z�6H܉�J>�%z��T,�������_�ݞX�}ʴ�*���Q��DaT#�hc�x����_ʞ��8U�W�G�5Z12%�.6��&�?��Wd}X�{��u*��YG$6��c���^�6�W�6O\,��~��҂�M��C8j��"*(�Ji�m�ȡ���x���}@�?%g�0�Ƽ�]����;�"�p�������������߷���I�����C;��Q!;�R6B#�"e2��X�1�<Qg�ˏQEV@�瞱Dy���4���K»F;,$��9e���\AQY��B��߄Uw
����Ȥ��!�`I-�mP��Mr"4��z)��,*cƯ�Fp���F�Q�����Z/ #'"~ت��d`�	��V�'�>;��U��z��E(��C賩����U�ˎ!�7#-�8C,�O:*j����511$�D�2�|E���O�:$Y�{���(ɿE#f<�7�����>��D7kƑ�(�7��P"�#��-��0����6#-�V�m�ȏ��{�C!�,Nu7�eG2V��$;.�b�A�q���~���Z���#�3F�H���{0Q�%�m8�H��t��"M�^��s�����C�zW����_p�'�@�����q箝mLc��A�[-[�@*�f@wn��'b�+.zRU\�=���w�3�,!oMgȌ(��ɢF�YT�AG^�U�d�"�d��[Q���Kbg(��A�[R!�����ǮGVQB�Kd_���������sa课��Ҍ�������ȵ��(��"$�pC6[������l�(�˅9�}g��g���2N��fӛ+��U�z~km}��>B��V� �m�s�;�2u6=!��㆏,!OƯ�"��g�Mp�K�S]��4�vyN>�<����T$��$-��R�?i�gź�����
~��D;�,�d4E��f�>daA���!��8Vws�W�J�՝�f#J*�b���U3�VT��X�[3I�[�!�z�y�ҳ8w$Z��j�պt)�l�P̫����/��)�
�9jU��b��fU�Py37�}ji�N{41m�ےF�1�!�����Y�e`���RWt 
�=K�����T��}dއ�"���r��V�UT��By����x���H���:��{8d,qZۈ�ӬU�ng�`�.���������p�\�Wk�F���V��i�T�5��㖻4�n�S�5#v2�ڮ;�8;� *TU@�� �F�����X��iv* �\ʽ��%,��~�;�X�)�U���{7g�6� w*�^   �8@*�U/V��HUW^���z؛�s�$�mێ��q�p��f��)���E+mr�Sj���cg{u;V�*�*��y]��lJ�Uc=٦�l
�[ �*l��`�Q���
�� �cl7-��wUP *�U m��9j�g�B8Vˡl�@*�8T*��R�6�ͷ�W� �P �  �    @
� ]    -�h-l��ش!�ԑJ6ZE[8CT3�f �4%Q�w�qܰ���Ӵ�5AUVr�{6�m�@���gpٺ��PSm�v��P��n@��B6	��X�;3U$���]؎�U<kiev���%iթ�V��u�\ckD�a����K�m�ظ� �e z�:������r��m      �    @�`   �@*��    �    UE[�@ P       
�T��       *l��wk�  �l� P;�   �  �� *�    
� M�  .` �   ���mkh �U�m�m�P  U �l�m�         ��  �T�6­�0 *�]�TT�u��  
��w����2T�@wn�d�:��Qw[mm��T��ґ-Ekp��R�(�ڦ �T�ndѤٮmۇ������%������r/TU^��w.�wk��=�Ƨ�<�%��^y�C��ګ&v�QZUecu�����m A�� Ȫ�V�W�}��8r )�V��f���&ǋ)�vK������z��B�@ x 
�U�  ����m��� 
����EWp`�� <)Pm�VR׮ثP�,���H�=Z.��X�� 
�U�U.x�Y�maXتQ�uR�9f���<*AU�2*t�t/��<p��٢B/!:������}�;1&�©"�'\����D�"���?z{;�j��2ҲM2���M��4�C����z>�7��ؑO`Q�����F�q���b�8N8�9��n�n',��q6$����#����V�G�C:R��C�����Zq�(�h�Ofo���P!�uY"a���`P$Q��G���b���7�g�Ɣ�è8S�*�W�B�~�g���]�>bV|�#�|p��X����5NDT"H���G}Z�v	��0��.|fX�:�9Q�#s7"�X,��n�����b{�����A%E(��n�񟞷vU�v����wCJ�T��J�DK�d�:�m��l����3={?x�Oz/M����9�k0�:��g�=�q��S���e
!qŚ0{����n"�JF�	9q��q�����m;��G���,ט��||'sb����D#�R����7x����mՏ��3y�-��"; �[m�:MfG�C���""J<�7��(�h�F��U|r��#%fE"$�Qm<�3Z!9,q�Bo����5����������|Zޚ�d"/Ї?m_'?x�+�}%�48�<k��,���I�!0�*�f�"̙��h�4�����F�>Dkr`���d2��(ސ�̎�y.L#X�d�����$��i���� lv:�!�@�-��F��r�*�[ ;��*[>x�q�1E������a���7�d#��HC�dfO��c�v$�t��<D��*ǲ��4t����xX��Im��jёi�i��[��g������sD�p�#�,�4���� �m�wMa,�|ܓ�Bf�Ԁ
��,=��O>���|���X��ٿș�-z�������̲�\:^�7�"�8�N"ʈ�H���pG��c�,�7�ٽ��ah8���!�p��"H��P���I8[��wy�������HZJWS�_ϒo�e���qX�!;�W�8F�����(鳺�B���T
<a���������P:U�ɱ��ڪ�ggk=�=n�UxU<Ir̪;�3ų�Y.&N��V�qF�iMǍE�����8r�B�ގ�e_j�Xəs14����P��;婜���f�g����^��|�{�"v����>�8�1���<Q�P�z_u���xj�����f�C��E�w��f��^�j-�b4�E�[�L>�f��Wv	��D"�4��A�T�`���C���57=�o��홶���|k:cv�2B�+BKH"�0�*��9���#: ��Ǣ�db���w�-��#�	�J8�?'�\���>�Y*��G,�$Ns��/EJ��j�����#T���>���UTk4����ۉ!!m�J,8����"~T���u�#�nh��X������H��ޱg�c���W�#�yo���)Q�rDP��T͒4�%?i�e��M$YB��a�gJwhqFvHT�C3�9~��w�͍�&�rBJ]-Y�3�����#�:�
���s�ә�8�!�wqE8�H�C�Dqp�^�2&P���H0�o/�Cx����$;�;+~���;�YV\�w6E�Ԫ5���^�B�*&�id�p:�����p��f/�,���QEZQ����8�`]�}sO���Ok��]������P��a(
���N�Nݺ<���.���v�A�K��5RVq�S�l�.n`p��n�U��h��(�:�8*Gr��,����LQ),����c'   T��Qq���a:ǋ���d�;k���tm���SΌ��P  �   U T �l`��n�� ��o]U�F� 
bV��p�s2*{f��=�ێ͙�P�f��:�9��f����ѻ�]��ʁƪ�V�UKm�����5�I��j��t���noMd}����@����"�H�����C��̈́���-�">�ژ�H[i$n�]c���;��w���� G@�%�r�������c"�f�|��e�7]Se�[`�qo�����!v�^��=�����#�J�������9�Zq�F�,�3As1�P11E��47�֬�|���Z����aߕ
���<O}�l���­5���I�a4B�͸�n@�O>��,��U�q��D�Y��}� �/ _���?<�@ֹ�f)3#Q8�ҹJ�)B��F��յ#$c�N��2үP�J��eVW;c:�*�X�p�*�uh���1Ex��4xUz���,�D��O&Ƨ,�ێ#�y�	��٘}"�6�I��A�+Tm@���i����sv���f�7{oǒ6z�M���F���˄lE��#O�Ҵ����y��h$ܒ�ҍ���#Hㅱ���p9G�DxVW0}G����G��� ���~ߴ��\C
(㐵RUUp�G��{G�T�7^�����#4��e�i}�w��~Cu~�:��l� �F�Q�_��(�þ�����=J\q���)@�,�'��#t��u�2�#O������6 a6�!mm�j��ll�	9*���V&S��U	UTb��0m%�8�����ߜ>8C!�x�����e3�D��6掟�P���o�C"��	J>��3Z����H���RH��!�>����H���,����i��i��Bda����Xן�ٜ���ւ�7`���3&��J>�9�SQ�"0��r��}� �{��8]�ޥ5V����YFq��yr���]h��}�Z+e� YD'ۅz��,R�̽#��VxM��o�#�:k�è!=�eH��6��D3{m6�d���$�A�н�Y��pѿDzP�lIDwyW��o��������z½��d���"�љ��v�\)�[UId�ٺw��^ǰ�UY�OAs餮�H�ha/��,�ɮ1�>����nl�#Z[W�O>�dlAN4׏�Nt �r^����D9 �Y�4�i���E�<��o�7#�E.��|5Exu_p�yk<w�7ݾi������R8�Nzm�pP9xZ_q�3��c��b�M��=��_.��dЇ,��R�$�D��Y������/��8yQK��x�4��Κ��T��O�f����i�qj��i ���K�nt��U{�c��b�[������������`#H����z�ֆ������r��bac-�]-\����ɇ�ָ«©�}��U| �U����]�%�)Ӕ��&���?������p8�=�@�Q���2�F0�+!JGk�\��#� `�������pT|�������yC��´<,-6��ȋ#�<��������P�k��(��gFRJ!p��A�%'i��0��g�~�<��BpJ`a����G�F�!�ʭD"�[Ķ�!f3l�qC_��o<�X;����L72G����:x�=�@�Q���9=�9��:��;�K]�c2.j��I�da��W��>�1��Z�DOd
!��ůT_Ȍ"ϸv)�p�g�"0����So����g�%�Ǒw ���I�qޯZO^c�l���S�s�8M� lm������Twp��s;!s�ڷj�����'f��'6��=T��@ ��-�X��L�-�{]�	k�C:6�ڐ�-��;�"�N�����T�@  �P T  *����(w�6�� *�eP<n֛`� x*�-!2���`A�ΧV]�\����w%�MW�^8$m+m�TT%�5J�R�J��������&*b*��ET?���,��?d{��C!��48�>�΀��Pf.�!��j��q~�<y�&#J8�m(cn k����e�Q#��4�l�� �l�s�x�N�|x���=�Y��΢d-�c�"dl�F�Ό^ď}��G�����j�:�7Q���HD�@����[aG���w�)6a!�q�BG6H{[�D"7�d",��eZq����Y���{C��AŞ#MF�s�+�h�`I$��T.����5���c�D��g=S"(s�R.��h�����/�"0�%�>����Q���R�]]:E`��`���U�iJ��z��*�W)���٣c�B`yl?@��	��2$�	F�k�Đ�d[b�V�������I%뚪���2�HJ7 �|�͝]ׯ���T*7���>:��,��o���Oxy��]�O�6L԰�,(�)ukk5�o'��v/���"ye�W�G�U����Of�6�׳�NX�J�C)$l�nxB4�wG �y��	�;��8�t�)�X�e8����ܫ�ʏ��>Z�&����$ ͼ�u�O��f|M|�!�;�,�vgKq���5�����Wٜ7쟹�#��`�#�TT�eJy�ú���ݧ��b*��LdJҎ��R�k���g�ձ�{d;���#1�E�z_ۯ�9��x�'~Y�r�����+�RI-PeW��7�s)wWW��!05���k���w����fk5�{y��KHՔ�����X��l[@���]:C�.}g�����������R�Ju�W�e�h�.�z�sf���^9p�y��p^�M]�����^�������{�����*�}W�5�36���V�=Z���]hCۙ���%���]{7��F�	�1��
�$�U�k�����ۇ���[�w)��p���U|g6G��G��4f��A��&K��a�%"�d������D�ug�����(�9���G=�J�Ӻ�}��Bc+���8���Y<��)�m+$����J�T��U[J
�זW�wl�1&�fr�j�:t�C��*���G��0��<x��]�X�,��%�똪/�~�_=��ݖ�R[G�:Q��u9VӜ>!�-�����3��wL�M�e18��?�>��L�j�D	�Kv�(���)9,�^'O�f?XG5pp9;���LК$���535'�/d������>�J�sJ�R�)B���X���!Tݎ�4�:Qӏ-3 ��lnn�lE*��_2.5�k���^G/m\-���}�]�xԨY�w���q���������$)$m�	c��]� �˳F5R�UKmJ�qUl����?)܅e���N�5�r���<_�c�:TF��U�Es�+;?�҇����+]�g�0��MQ��I-�:�Z�E�������^ɒ�����d�l�!�}�h�6Yg����Qٚμ�}��2����CC����\�Y��0���8��@ã��W������Wg�l{�7}�)K$`�$�����^c���zQӊ1��+�1���
��U�EUl�XrY�Y���ψN�b`�DFА;)��i�����+�e�me�%,�Q��QĤ?.���ghbʽ2��=����m]tS��/��$�붕���rQ�;$���,�z惧���ң�J �]�fn�Yws�P�UPx���;y�ihr�^���-�%V�9�]��	�FUU�=M�� @����H�$�q�{X�%�s�]�`kl��&��  pP�� 
�Q]��`U�m��
�UP
��P;��U p������6��.�E�.X��	5�6%)@�9��)9�ڪs���k-�h�Wj���
���~f�v)���DY��5#�g���k�t�XF�2X�R)�4y@�
qMG�S��4�=�r��,���U�w Q&�I��A�F��<_�G3��C�Q�6t�G�s�����IG	B���"���l��R���!e�p��G�|p�Zq�4QWZr0�C.v_�c
(��P���$x˂a��4̙�$-����sW��<�(�:ֲc��M�x��=�)�l�)�~�9ͳ�:�����K�
U�%� ����'�<^��l��k��F�]�:_�m׹�{�Q�����Y0��!*�2�I�.�S��[e����UJ�P+@**KH�h[Yk���A�;H���/����mc6���^��%���w�=os��:��$���$�u�<׳Q�-��tߎ�d���Q��בd'���d�YZ'z*�,�'��]�:Ԣ���86�R&5(9#��|�|x}�ze���@g���E��x�R-�k��Q�_w���7ڶ�?���&ۀZp�6|:�H�G�/a+q�,3G�a�,�M>�����Ȍ�����]�F�I$d(����dIG6Oƃ4Q̆Z���k�����N�K ��+O�4O���?�	�rN�t�j�#�[hݸj�]��Q��%T%YP�*�AC�BC�7��qxqg�x�����?I~ڶ�O�݄����uY��;����>�l�����$�6R�{��8a�c��p�B��V���]F�	�Q��x��W���Ș���5LUDU"`[�Kd2�|�26��y�4�7���f����a��U�Y�zrP!ǎ�e��q�g��6�l�����<l�5A���XQ�x���$YC�r��i�¥k����Q�:�d��iF�Mj�kY��!���{��dxd��!~S>��yp��:{�_U[����*�N���"���U[�nv"�	��Wj��-�;�AUUݼ�^�,P�r@�6AZx�ϗ���/??~�Y��S!��A�,�	YY��G<yy�6U@ Z&8��^<|y�g�W�a��2�Y�^0�^���"��z_|�������h4R�# *(ETQ�!�3�п;�Ig�eZ��6���X���K��j���*/]�rX�����β�k2m�����w�\Z����,�ᖏ��'ݹ�Ջ�a��/q
��`����h�TT�ҍ�����7K������u�Oj�h�:u�m�d�,����.�Y%�	��-���%�����A�5��-m�{9�˸m�Umؕ��w1KU��-�V�I-V���%�,���~�dYElz�#��L�+�+�zd%Kc�:ff�y�0LdL�&D"d�EZ(��t�E�����8�.P�l�Di��B(�?B#*8�t��2�G�FSf&�Ia�Dv����^��la��t�˴]��Y㸸Y�Pqgyx����ݠZR'$�#�2x�����������6�<i����;p��ŷ��J#
��2%���&Q��"H�l�G�<R*ҁn�Ŏ0רg�R�#��ʴ��q��{`#gg�y�8���>��c�"��eW+v��''�b\����ݪ`խ]�骪�tV�������nU ~�V��S�c�y��y֪<J�d�Ql�[f6��ꡌ��  ���޻Q{��-
���z���?/���oTS�5�{���   <  � J����
��� 
����UUܪ��6¥@x*���{jy{��=���L�G=�,潔�j����Z3��8U�U���)�Z����Ѩ���BO�O�sa��l��C�w-���0�o�2�ݕ�<t��Ɉ�
[`7m�2���ޟ5�2�"��$k�W	j�SZ�/m��s�����pH�d�"jBr�L�"��<0W��7|��f�����=Y\�IF"I��=�O����[ǟ�~�]_G�%����ُL��I��#d�XNE�쿸Y�?Gu��Q��8���V�ǎ�x�0�D��Zzd�]�.�#��,��+[jM��
���M*�J�5cR�������.��T��2f��-G��/oVG��> �>�Um@��<[�Ǫ���Y���d4Zm��KmE�W#�;�e�+�C
ՅC8q��~�������?�Em?��.�i�v��`����i�e���7��"�f����H���x?0{�1��9�	Gs��M�fj�T�Id��<r⏙z�;^l�y�{����Th���(�ö����Ì����3ܨ��Y�0��AĥB(�~���t���˸�9�ӛ���i�:��G�� �X�b�׮q��5U]�l��@*��9���J�����qJk��E��yi	6F��k�|��>=DMR�4.�>��?����IU-�d��㒻���lϋ,��3�v8�G|Ew�K���ip��< Óq�,$�6�I�DE���!G��wԽ~gyQ�kg��OV��ķ���w���skRM�m�����*z��v�w�?p�E�A�g��;�2��gM�o�s�;�do�V��~�4��	�+�Α�A�ʴ��f*j4���@�7��<h��'z��ZE\E\����R�9sѳs��@�X
��c�]���R�T�UK�,�M]���e%����#8��gƸ��p*P{B�6S�B��b��2l�A���]���D��.6#\C8o�n�A��(��޹\e��s���N�9���U��~�u�J;)d�P�,C���u���j��4����?e[p�x뇗jv޲u��k�a��Qg7�Ѩ�n$���r0\�Wr��'�	�P�h��/$��,(�i���<l��1Y��6��a34F;�+�"��z�N6�04���]��>���cU����#�3�0�F�/���g/r���	�@�Q(y>�q8Ȋ�b�%������j�S4p<����T��T-�;��]m�JE�外X:�-nP�Zm���uy���2R����M��_��~ڻ[!�|[��q���o�,�M���*8��~�����b�SV�Y�d+�I`����4s6�AC�Q�'H�i���2I�$�h�i��Q��Ӿ_�f���"F��z�p��4�[9k���\�E?� d�Hڂ0�qdtׇ����Q�L��wW��na��qx蝞�}��R�Ww�����QH����YÞCxק�t�����VhDi�l���ګƋB3��U��s8V���,;��#&j��8�j<��>ٓ7e���痯׊ל0�E�����yO�]�Z��uY��,+{~t����>���uez���u�W:��v���j �J�   �=��+��=�TU8@  �.�p��aڼ<���w�a�r�gEs��<��񫍃Vf�v#2ӱ�Ѓ��mu˱;���quF8�' Z8!VŐ�N{�\�:5�q��{X�;'��N���NTiE�kr���n�G/.!�v�wYz�.9�����dU PU mQT 
����ok[ *�� �C�m�����P
�Pd�U �
�x�<5�U�n�m�S�UN@  gT
�ځY����8<<���w�}�nض���G�Iٕ�7*1�c��`��WT{��U �ʼm�I��U@�U�.KrEm�� ��Hn��l�*��@�EP�V���ꙗ��� �g�ں�u̪v�s���o}���b���{�1�p�@  c  �6扲 �F���      U*�@6 ���-U4�.�ї2��A�UH��T�5A��g22�*ʪʤ��E�K��B��յ9r�b�h���@J��緍����c��H�T�4\xx�����K��w2f#*��j�iI�vvn��N)N�f�6;l�ų:5�-�fKH@;��Y@�к1�Z1Z����[ck$>����   >�    
ʪ@  
�\�U T   @  PT-�   *��    U R�T�@ T    �6�C���   ;�   p    x   <UUY@    �  [[  � �    mwu`�n�)Y��j� \�P �6�� �      �  �P�   U  U��UwA�T;�<n��{$*���٨���G���q���R�$�[m�*�6�+f�l��
ϞX�qvyƕd譯�����[x���f�W8(		�ٴ�O9�<ӂ�����Y�$�K�MZ�6Ukh#�YH�YVB@U�VM�TSl�
�-�/-@�&݁8y��d�ó}}�gn�l(j����@     �  
�P��wl`�  ��6��*�t� � �m�PTp�(fř�{g�Q<v��� ���' %�&6��m7[���۹6�*��Am���A"����+�}�ko|�$*}Zh�����º�]9Hn�O��d{�M��I&Le�"'%q�@f�A�daÚL�@a�?l�}���L(���6H6�!�E������Ď�VfD�C4ק�^��d��;��y�Xt�4U��1 P@�Ek�4����v��r`�;k����M�#�4ry�k�̥G��[���~m�#�(�r�UO��dn���Z�r�f��E80M�R���A��b�{>���̕(�!DU�g�]�s�UimN�� � ܃!;T����gE+U@0�]Z۞V\L��{��"��Wj�M�TfMa�C4�H��Gƈ�ff��t����\!H�T��$�{B8x!�*�+�]��G}�+B<vm.��w��V�p���=���~��m`N&�0�&ҁ��3��V{���h�7u��V��gtRF|ս䫃�4��>���$�-�$p��!%4wf��S�8��Q��܁<l�EFap�{`�o �Lk�����0,����{����XDx�m9B�󊿦�)+�B�4R����5�R�,�<EsXS���(�.�W���jp�������u�
�����V�*�����Z�Ux����)��DI㾆W>��Y�D>�������سǹ9�w���R��j�3����+��H�;�2��f�t�:9�U��t�Q�����}q�UQ�m J�"j3R0�C��c��~���W�ߴ3�ߑ�'u^х�C�R����9t8�ܿo\i��n�2B[���>�l�X<]��Ǐ~ҏ �ÙL{{`�G�Ró�W�{�����/�j�`H�-Z�y����\�84�Po��_G4�-#Ŏ��'�ǐp�{\1*�$,P6�4��-!BY٭�+b�ߧ���ڻ�S�UW���4[7/N�V)B�����l�o��˟��ƈ�3|�{�x�Y(���VG@z,6~�䬴��`�TQ5B�4yG�Ġ��yu�%|{�<ys���C8s�쟸�-�*��F�n0[
H�I����@Y�0jL#M��J���㣫���=���0ÄY��HE\&ɆH�b'%o 8=�Y�Y�����?i��E��^���t�o����S�Z2=�<8��y4^e�-�<�p�I' -����+6��(p0�/�	e���G��}��<w��qP�l�-�{D���]�s*<ƍn͕V1��/j���kh݂��T�5U]&Y@�� �mϑ�عU'�4|a���q�@Y����ӧp�����G�f�<Y�@M��Б��Q��Q�p�86w�w)�~\�}�QÖ�i���a�Dn��b�g�3��&I�j"�1�?+����A���R�t�w��h�S�1�V��G��O'ܙ�ǌˮhHI��m �g�5�3������/nW���=,�:�3}a��捞��/�h��%V��^u��~ǗyN��E����� #e*�5�E�d#{_q�L#���B�����1�Z���UG&���8]����۫m�Û��{����@ W�HΗf�4�M�v0��s�lctՙջ?=�ꕵ��R�v7J�zˬ� �
� T =�{n�U;�ʔ�dtUFY�֎��sս��� T�T -� Ql�w+��l
���R� ��llT�T*�<
�Kk=
�+�ٿ��|s�Ď���H�I	臷NW3KR�UfŹ�x:Z�٥nX%UV�\�x�Unun�q$�n0��v�?����!i�4�Z4<�(p�����
ɝt�=k�fg�Y�H�9��B�d�
�)d�]�ⴿ�W�E�bٓ�x��{r�_��5t4��o�9nFۀ�"I��b8%G�f�5&}��n��,��0�r��^��Guk��ǲ<�r���K�@܄�%6\����ߪ͞���2�{��a��!���g�ε�P�]��UDX2F�`�J�!	�H��8_0Y�q��1��ސ��p����O�S\Q���q�@Y}�R�"f:��U�+j��Z*#!v��>xڪU�V�4�5���Q�,2�R�"!|al�u��}�ō3T���s(���(��^�;���w(
�6g梅��7dQ�^C/U�ں���=U%�y��2{��Ⱦ5��B��0�8*`Ⱥ�������MY1&�)Ēm8�>�G�@-�kƎG��}J	EIe'�tZ�iFJ6G����@v;HqP5��7/�^���F9��p�6s��pigu1����Y�(�n���A�JHXQ�[��>7�Kư�6r�K4ק��E�F��+��͜B��i��N���[��sen�8g,�@R&�*�-��N�*��kd��y4�f�.6���)$��h��ݺ_AC�/y�gD��Zl� �i<�r���>!�31�{��� ("�	.���ξ����g��U����ő�R̴��@C��3TRou3�6����L�f4ܯ>"�pO�V� ��,׈��F��[��g����Gy��4x��{�e�t����\M��k�^�:{��3�Ժ
��j �{ƴ�Ú�r}�:\�⣐�X���6a!��������:a�<�h�ڲ�]/�s� �h
�!�����&�"����t=
�T�����8�)vjM�t�m�X�����l��-���:�v�u���ل���@v��0��])t|O<�,�r�����9��F�?y,�0'	� ԉ5E������z��Yc/5�@C���辕���2��i���{���P�	%��ӯ]���ӥ�|�7�37���D�?ʃ��*��t �������S�Gh�p:����5�V���f�@�ޮ�܀ӽ~K4�y*{׋��{�[ꁶH�� ���k�X��{��w_3q*Kߨ��!�k�P/6�J�qf�{�}ߣ���e���M]:�$j>�#d۳�;+U]���Z�T��4B��B[����ݚ /h<fj�~z�7�=��u9!�O��kk�hs/y@A�#��#�[(V�,�;��ӕ�0�4��wP�g�#���+ya��̪䅉	$�i4B�����=��h�_���:�t�;����V�c+�P����V���QȘd)���ћ �Iƴ��G'��Ç4�X'���u�:l���hI5J$�i&�E��Ν{�!��0xl�6��az30�o�в����]�qԏ���)[�U]T ��ŵw6��U��
ݶ��{\>��+(��
��۰~4� wn!�]�wY�y�n.q�1������V���6�MtPm�h �+�  @l����ע��:�Z�����Q��γ�0hU�-SU@�z�
�
�� U < ;�Ta�  P +ն� U ;�E��������ݣa�.��"�j	�Vn�&ֲ3�Ʀ����gf�]������UTv��ތ���i ���_|�Ǚ�k�[C{J�~w�~�,�<��a��%�Měm�Cr12g����Ի�hw��������!W�+;�Q�HF���)U5�pS�*�{8���I��^~װ�fl��t$�2���$�GȎ��w�3�FG��m+����G68RV�4ȉHÌ�R3#�\���hO�Vc:�����p�ǃ�,οf�V}�x�$8�S�v3�*��Ytm�Q��K^wP§��8@�ע]����[ԠQ�n���,������hf�G}��?�A?5"R4���;�q���5nm�@Ѕ�Jc�rf����>��{8�esέ�um�P(EI6�f5����{��7�e���΋�� �����H�m�I�Ȕ��ge�������{���غ河���k�6�b�)Bcm�q��و՟�i���>?�;6�iH�jg�i�5�-��e�`)l��\�R�5���gv��P�^OU]̈́�e綉��}�����x�,���0 F��+83c^J���e�(�Qٱ&��	&!n$ˍ�!������|N�����:~�0�CpU�qt/��sM�P�2H�l��UŐ��f��(�>����|��:����1�h��׬%�MVU�~@�.��%,��E�Y���=����YgԘ��U㷈�Meײ���[���K3h�B���0�����b�2H��O�����������6?@͟�=�R���s�%�M���ґ��5��֨����_��,��)O Cߢ����*�A^�@2!��E�
RN$���p��p��:p��2��wɎy�x���ڞO:�|>����: �6��fJU�@X
����6�;��]T���DmL�*0��JFR_ Q�⟎��a5��Ͽf'�m����d��M���-���n%����#5�e�~`�#(��~�0�7��<x��E~�����Q��-���@�T5�D��:��F枡��}�٧���C��}s��g2�������J7Q�?i�B���4@gwB~,�<}�wnPG��ڞ�h��A��	��'��������i(�������+Hx�EFx��f����FF񔥕�f�;�6�f3uW[7\�/)���L��̓��j�ڥe�j�UeP:E��2=��?δ�CM��!��u���p=�F"|xh����5���I�*I��C!����9���$0�7��4@�`����a9���_�"ww�l�l�A��g�f�q��~���o���ԭ?��3Z�Y�f�3n��YDgu�.C#ԉ5	GXl�=6Y��Xx�gE��J��dB��_�Ü�o�4=K����i�Ȉ�L�$�ekHFi�?�پ[ݓ�ő�+n�����X?�v�JV���V-��÷i	�T�`�y��u�r3N�[]�K�r�{�I�K[��U7��.�g���U�vC��l8�p7n�{`�*�Se��"�ke{mq�UP *� <��v�]����v¼@���v��b�h1n��hۄ�u�<�@ U�*�^�   ����wU  U*���]�w6�[�B��VJ�e�Om������.�4���<�QA.�킷s6��vu2�^�D��져`FG)I�V��{kn��J������8x}�R��Fi�K?������n6��IM���W�##x�S�. C��Y�����S?��0k�_�2z��+�M �>j܍�ÐЇ����xh���s�i�¼|Gm���N�C�+��!�W"�/�e�#4�Q�i�Q'0��G߳���[���VA��W�ǼUD��H�Q3Xx�3L��Fp5�]���G�g�|3�(�v-��q����M�w7,؂ɘ�� ']�2��Wj�P�SgF`�2�����k�;���w�F/1�������qM"����F��?a�N���I�*�n$�2!$�4@�7B��	ѹ�~���jW�����������ӱ�l����m� ��v�>k���[U��x�S�=�H����Ka��Y�$��4\��,�X�t�����7�c���,���ť��!,��Jk�S�&�νV=��=q'�'�ߗ+���,^��6���7�8J��[`)V�\�`�Щ�d mUU{t��	Q�ܒb���&kPڻûu��x�C��sY��m��0�፹���ޣ;3�i�P�ԍ紽�s�;�1ُ���H�-3����3z���0:�xV�V{�y���1���[^��6�D"R6�if��f��Y3Z�^~����y]:��E�	i8�I4�e�<��M�W�yFez��k��x�{�]w��I�.�X�Hbf��M�,��|���j�]���Uݶ��w�v8�"��H�����V݋̩��Dn��Ds3�!�~���6ˀB䍴����>��0�� �(�g����Hh��FY�b�m���-
��)5L7*�i���D�8���iTp��Qc�J�9��AXG�z����	)m����n��^z��q�f�tb?�'��ʈ��Ϲ�I�va��Z;�g�C��oqM��\I$Q@�V�@�w*�����"�������&|f���Z싾Z����%�X��(�#P��J��uRT�s�]�UBUj��#$ OC�q����H�x�����F;��|e�8�"��_��0{E\��Y�ff�-�i6AmĒ�&��H�q{ƻ��?��w�B0ÚD/H"��>��!�Ug+l����q)(9(C�Q%�Q�+�/��۩����|w����0��م�����m�n$�i9Z}��YXgyY�@e����"0�~TF��q*S���Q�8��V�H���E��!G�?��g7���i��8+��
8nza��~Ex��=�����V�==<O�u�Ӑ�  +.xUsv��:��"b끍�=]vyn0j�ԭT�͵���5wQm�WH��^�����.�	[�mGwp��|�Sf�]�w7Wu� 3��aP �(��{85F����볏(\LТC�X6�W�޿\���  C�  U@   �e����U J� ���`m�@ d��M���<{��gC&��t��X�MJ�7a��=,UA�ڧUl���'<2��J쾙L��52�쩩������,��g����D�R�OW�"��f������	�&�m$cJXG	#�˪��u���׌�#4�١�#�"T��h�W�x	P�c���׏Z �{���|s��>|hi��L��'Y����u��_������n�HZl�x$�d���#�+n�>?�xOu��{���?وx���P�&TpF�-�6�6-́"����Yg����dG��n�FR@xq,�� cQ��&n3�P�j��r�ê�ݵniWj���BG2�*�6��&�-!���xß�x��7����
>�>|j�W�61Ӭ��Xwuӊ6�QD���,���3�+����w���(��w�#{�O�#ƈ܆��>?�̅t�ʘ���хl�А+�9K�5^�m�{�0<|-�@�V�{�j���3Z�(��{�m�&���q�J�\�_�P.�BFq�(8���?j����U������|h0��u���B[����vi�>=�y1:����&�wn�S���+��>?��M�P�%��R2$a�5�FA�(��M{.�����Ul�W�a	�b+�B��6-��� L�K��O�"���>?��%�
?�۵XY��oW4�D�d�m�����gp�ٔX%{�����K�H��V��v�3��q16À3�0[��#L?��5Ɖ�	c5�dЁ�u��珢���~�x��n�DG��������VRI ����'����N�i�dC�٩���+���*��{��741�i%-���]�͜�j���l�e",�0��F�������gH
�YԚ����mMٹ��XmPN�*��J`��*{,J�����k
��5}��	"��M�44�4g�hC��Fk������SSF��s�Z:�� h����a�n�[�(���y�U0��u���ȇ߷S��~�n�ñ#&�F�Ϗ�]�Xi��Fo/|�z�����GGq��!�C6iH�� ِ��m�a�$B`�ϥqssM�8�æ�B�#b��!�F�"wƮ���^Ɛj(�E(A�'��g9�W��J��+^�~^�wjf�VvD(��&���ٌ�;�1Lg��`�`LA%�2�����d&mUU:����dd8();�mo���^��o+;��u�}��Қ�1��Q'
!�����gv���{���-���f�>��E$j6LjD�$�rc�����f��p��z��g�G=���=(+JC!$br��=G����b�rݞ[����ʎ��mQ�P(�P���˔k�wg�fW��}�ٳ]�?}���{��9���y��		��$$ ����А��E$�	!֐�, �I$�h@���	 1���!!! ���B���!!! ���������������������?�H DH �! � H$��� �!��!$$!����!!! �����D��������>��		�7�2BBB�BBB��!!! ��5�BBB�������]͚4IIL�$�	��HH@?�������BBB�BBBB�c����;�?���$$$ ��x��~�$$ �h�o����e5����N͘ �s2}p���Q**��I* )%@J�**B���R�HU@�UJ����gcI%B�"�(Px          >   �            
    �  �  �  �     " J�wQ��n0�{������ s�
w�ХmB���݅9��*� 7U
����4�dR�C4��s�%OmO=�H�G� �R�-<����Q\�R�2US����RsǀނRLl�f����9%媥��$�-.ZE$��  � �     " �D��s�^L���9j�\������E(��ǀ�IH��G�J*���G�H�Y)$�i�;�RJ+�=@<�RK,��P(�b���T�-B��t�������$���ǀ�4iE�^̕T�ۢW�E/-"�r��w$��=�<M��J�+�Ҋ^��R*���JI��%*���@�  x     ��%S���R�{��픒�2�K��=�I$�� �QS,�6R�\��͒���]e�d��u���QJ*�[��iK<���P  �=�u�W-@:xx�z=��gB��\�J�b�Mi��7aC�����P�o^6�tR�s:����
[ lhx �     B �u
��P�,����ҫ֛�s�)E� �l�B�ZU
bj�����Kճg��)i�`U.�N���)� ,��Ҫ�M*�<x {ԡLMy6��M*U&&�k�6�mJY���J�Myj��{�W���%W-q�u�0h*� �      o
R���Ҕ�e+�e=�u*�{��Kim����JR����)I{��<���+�e�*JHxp �^�R�,u�!r�S�I�{�u$��m�)*.�<x w�^�R��{�d�',������RJ�ǈҊ*9���P�����R��Q2�R��U\mERD:�91T�K�����UA���hb)����hL�
T�d�z�D�@h�Њ���T)F  '�T�2e)� ������(0� ��\|�8�ν}I˧M�7]p�=�}7����:�k=���ￕI�g\}U$)�R@{*HuI����������<���9�:��ΰ%Z"`J���u)n��D';���n�t�id�5��N��s-LN�V�V���
�X<�+�Yڙ����CE��SA�v�!	Z�1t��U��Yv�+�y��d�c1���]n�9��^W�W�N�5rp�#�^KGL�oSA��Y�N��@D�ua�t����ʪ��eT�(�%�oH��Qi���0$��FfRtb/*�q�O�*4]X6�Ti�ܫ�M���(GU0�H�7CT���@Ԫ3����T.�pa�89}ʹ2�,i1НvqP��KR���Ӕ!�i�ĩ�IV�ۉ��4�"h��_=�Őɉ�+Fb�',��x���*sscnj�T�[$���[�	+��Z+@T�[�*ʊ�((Ie�=�E�9�:�˾]��d�^��홙[���:�X0���ڕ n��J�*>�1����Mbp*��ںN�T-���ɰ˱ej��p�&�cl{y��F���.e�AV���	�*�[̰w�x���˻ga��e7%-wY�����iP<�M
�Ķ��w5f]*�ئol�9ZVk��Pީ�/f�2�,X��6f��ɹ��%L���e�{�@���m�KV���wjC�hǡ�ç
��A��ұ�A�,m1KX��M��t�W�VQ�^�����2�e�$V�E�;Ol��詶CҮ3���+Ge�l(hM՛L9y�� .�AF[�Z�i���x6��e⛗R+N8��3i���Ք�FnZ�yl6l���v�5�F�U[3����ix�!U�q�y-#�j�W�PJ5H���b�����)ɳ�d�%������M��	l���n�Er*ل�&-��:��U�m�P�UHtު-Z�
@s��l�:Cw����ibv�\�"*�N�"C�\�L�T��j8V+���eZ@<��#.�/AHqcc�]�ނUpS����99�N��:��զL�Z���ȵ�c�/6Z�@�5p^un��bA�Niƙ�Sz�!Ժ�o�+|�ci��m[t,�ué>����m-;���<�W�/���'f�w��a�
A"����;��J]V�:����@�%t�&4��,�.�J�G�JzXTvP�i�6[� �����׎M�ӵ�5�*p�l�oq7��yn �2~FkU+!�f#Ǡe�-5�0�9�݅��Z�Q�Mʱ`*i�)���B�R�le�hU -[�Lx�e��:�j�� v�eT˗�kh'ko�0�X� �hV�V�{����DP�rᨩ�ַ-�6���=�n�ٲז��
,�6�M�e�,lj�%ڶ�t��Xf� �t�&�Pw.�7�x�'�s�:�YC��F������%.��Q��u,����V�]�{�X�FV�����d8�,Z�����<ں�8:��� ;���q88%�'7JS5c��;� �MSf%�l�bP�t�\�v� ��aQb��[I\�����(��u�)�rb4q4�Q"�o\
#[����%ۭ ��Q���ؐܨ�0G)ܰ�m"6�EI�2'��HY�Wg)l����/�EY�2E����Z�Pg�Bh��V��>�J�ڔ�A�''����=|T]�4��j�7�J'X�TQ�D5��4��T�%ZT�nXԮ'0Lt�&�)�M�Cu����V:9�+��Ym�6�iLj9����4����u�Q�S�)��4�Q�Z����ʱ+j4.�Z�$aOjI��r��*'a�Q��z�Q8�'�Ֆ�tY���&�tY6�𤃒���)���^��5�v�N��:i�<��^��E"w�z^Qv�[�Ieކ�F&�;�����8nc�B�%X�Hǚ�m��7V�H�%ݩY�EshE]�i����i8)n�ca�zc8���D�����#vB͑t=��z,��6�\��^��1QK�YLcU�5��ϳ7n�����h�W��vE�e��(GQE��
yN�K��R�F��dSn-��Z���gt�T�:u����v-+w�иq(m���eSc�����x��d�Ge�l�b���ڶ4ĳ1�#.�i]뢣qgU�ԩ��bCa�2���ŭ՘��5/n���7��;DTNeR��JB"TUH�JD,2�����͌�W�!6a�E{WR�VC�9�uo��歵�WUd��G�oi+�������6�7s6�,c�1ٺSn��Yq�7��[&�l��l"�Uw���`�QK*T�����٩c̷��W2�%Y�V�A��p=��Y5�ɩ�L�tI�@L��J����-����t���ɠ�c1푠ֽ0(�FIB�a���W����(���9D�DV�1�k�B̽�!�A�{Z�s!{
�SV���a�	�y��M��-�B��ԧ�|�����:�l��Y��Jφ�&�Ekڽ�bc"�T�΍Pe!�f)��&V�@jOb�Z��7pbTTts�a���z�GW�M�2�EQ"�k3 ��y��4��VF�"G���e�-MC�7^�fڑE�Z�������Qs�'�6��z��j�Q�Fe�K�� ��5F�R5�Kݽr)XԹ �Q7�E���J�Zu���1^4���M�D���<�o頝^�$��U��e��!�v��ĕ�ZUP�N��¶�+L�!�Ǘo(���2���bf}���њ[�L>]�V� �-νg,�rЏ�ء�])l��S6�bZ��}U~�[��݅ߩ���zU=�5v`�.f��_R��f�n`t!��_u���M�����Z8,�t�Y�&� s��;*�u,m�U�ڒ$D��{�]����T�[�71w9Z#.�I��S.�����P��e���t:��Kz~;V�W���i�KT
P�"v�[�ѭ=�Y�[�3M� p��3)b <�����݆Ej���X3`���ˉS{t�n��N5�f��~z��H��Sr5��݈f&jE��٨����tm�����QU�	E�w��Ô�Z�l�M�7�U\�*�`�VZ�[��ٰf�ɸ��p�5�X�L�S�y4[��,���j3����0�,e��4KنlhG�� ,�$Q.�=.�2��f=�����	�/HX�,�SW�n��F=<kp�t�t���i��IK�Y6�㸷����oudsq(������0�̽��ehi6� �������e'$XS�x��+t�3f��҉�v�Լ��cE*M�Q�7-�^�3Y	8%�9M�l8�k�
��vQW/-=����/M<�{�K	吅bВ��'{-6�׸�",�oV*�s5T�o�i�(j͓U6�ԑ�Ǝ�a,�/��q��e���C�W�)j
�E�K	f���]��"6nLt��`�%`��&H����6�fcW���r��3������ψ����� Y#ʣ�n����`����%��T#����;/�)OJHe[p=�ܟJ,�/�W��*�+7.I�QJ0�Eՙ&���Z��C2`��T�2����B��� UyZ"3�iڌ(��'�	���O يUɣ)Q�w�5������0L+4'	�5� ԄZ�j�M�����v
��m�[��Ӯ�YU#���8�{���R& �ᛡ��b�`�31�W@5E�ۥD����Oq�9��C{�P�8{��v',��}�a��5��)�	�
ˬe���]k�u���b���5�TsA����Lʴ��g�v�n!� �z^\r�˘��h,Df�!n�Rt�NM������P��z�h���0���\��% �Z�LeԽ&�zFc%%$��R���ƬGt]�WZ]����An˳ d=бͻXtPY�u�Ev��ʹj�8u��C\���0ĂAęֶ��hjh:��H�4�6�`y���Ũ'D\�1r�y�,��pX۴���c��20��ȵ��fA
+�ʳC��/��G���fҚ�Ŷ0fɷ�]`4!��Z��N;Ԉ�m0.XfKb=�A:b<���̕���(;�eZ����1V���Մ>i�5Zn1f�Z2+��[6������v���45�^�"���)w�1�b�4nJxi�y�e�.�MYZv����L�r�B*%.�se�fd�U�ntp	3 �xc
���\N؜v�:��s����"��&�;�a���#sF�S~ZZz6�غ�qR�����jسc"3h(uQ�Z�̃�����������R�j�n�+��I{�V4�or]9f���U�gU�z�݂�=�r��#r�h�E��7r�"���OpY��t��oÅt!yӪg8!���g<A�����^�O�i{ď`�Q�)c�E�d�0��
3
=�.	�	��������>� @�X��!�]ړ:�Y�,x�Xeb�b8eظ��ֽ	T���	YW��*ː�<�S��a%G3�ç�~�*؜�j
�8�(L�K������k�4c��L��]�gS͵*M"�5*E���ûo#t�9tZM���i��-ǥ�%S�������V�}�k>xo�6!����A!��6�*���U�-Hu�L���#d[Y�3Zw��:�	�^�`�f��i����W����5�b���^��$Z��p�pt�8-ҩ���t���*͈�����A�[	E�M������]���^�ۋX�VR�O䲮�Ǭl��U�0e�N^ml�,Z��B���Y�UA��ba�ʛ�eP�z7M�f��̕���i5�0�ɦZ��)ݔu,�e%f�N2V�i��n�b�N���KL]۷��a�30;�:��3M��q������c�~����ŧ��������`Pbc�R�V��X�eۻvT�D�sl��&읬4j���H2�D]��ɺt	�u�B̶��;2�Y�A��$Ǎ'GI�-�����XTƮ��7M�"[�Ô3a��n�DL�j��,:�f6S�@�82��$X�w�(�Xl�ˊ9[J�G5��-ͩ>i՜ij��vU�[c���*�f�ekJ�#R(�m�f��15��H��E��i�fۆ��D^��i�	,��n`����F�m[؞R8����ӂP��,�9��G�%���;���� ���hhg)������jѻ8�n��Ӳ��M-�k���g�5��.�hfk���On�ۣw��z�������|k�o�ݛ&��<�[@�=ͱ]弓�]��u�"0�FC�U�Up�+L��mn0�J����wT�݊`n��&"������&^�o(P$�"��;��������L
ݺэ���P�
������v���-�
T�=��8<��a�ps�����b������黵��^��\wH���b���k�.���X��e�ۙ�,DF��6�8EW7^Ղ:Re]��S&L�%�k+ �ͣ7 �CQ��w��nZ��L2r�e��y m���xʻ�o5�B�ګ۱�`K���R!�
�fݫ�[�Fk�+[�O��Y���W9o�7+�6,�j�&YK�H�Z������5��lL�%e�.
�͵Ww�nLwV��I)alǷk``�v�TAl���G"Te�;kkwsN��'������5���e
t��H�m�U�c�하ᚬ�6��ݼ���|�       p                ��                   $    6�   -�9 m�   6�      C�     -�v                 �Ć�Kh        M��m  $8�6�     m�   $                     ����                       � 6�                                           ��Ͷ            �o��y�u�_8�m��                          �q#� t�m�Z� $�                    �              �             ���  l     i��m���$ m���� �  ��  	��9�-�ڶ�����r� �(  m�                   h             �`        C�                          �                        �   m �    H�֛i0/Z H۱��                    m     �            �@ �P�6�      �6�'��zy�U,�oM��Xy���wGm��j���Hě�����=ֱ\�C�Kt:�	h؎Mny�<�i�6�1p]f�7n5��a캭^U��f��s؍CwR�q��Y��t\C���l��@m�����N��Gr�g;�xNN�+��\q�`�Tl.w+ŧ�9�vON۵��ǁ:��׷k۞�!���)w=�y(u����8	}��g�ҙm����}h��c�m�ݕ��SǷe.s�I����-�����;b�#�읖�u��r<��f��1)[�Z�vQ���V.�$���.v����sc�؍s����>Z�&ɛ�����לq��cS�v�yq�v4�r���/V����nN���ot]Ϡ�݊�ЅN���f��yF9��CQi�)t��s<�M�v7��7G&+p�Cr<{/]�^ø:v��u�v��#l]�)��p����-�����T�cjOos�I��s�n�;�j-�Tv����Ӹ���X�m1�F �CE�����rʩ0�qgs�.y �$u�ƙ۪s��I,�n��3���qe��v���Y{$�uQ�ǰ�0�2�q�"�՞6�`��W��6ul���Ӡ�=�ی]��L��S�n#��;�VC��ƍ��nZ�2���s�h8�����qu7 �.�p��v��u�;�ݹ햛��F�;��۩wlE�M�NhĶl����e�W��y��̱�mN;n�yL��q�pm�[)�#[y�n�usk��O>ϯ=	�V-�P���ZŎ��l�[�.L[��[p���P���V^��@�q��)�#�`S�����|��>�\;v웊���7��j�x����������)�q^������G�uۮ�Ǝ�e�)�uyX�^K�Re��R��9=����Xu�f�{A]<;�������^�ٺqWa۵��Og8���4F�`�۲��w�ζ]����c�sؖN�s�g��1Վ7gm�wb���؂yX$�d�v��Skl�^��n4�r�xG��4Y�F�M����[��5���wVי�	l�=����F���Aڇ�{���;=���Sj���]�%ǖ�
�x�\됀��u��v�Bi��8כe�lBxl�m�p����������jF)1��3���=!��"|�ѓ�v�bg��G�9��w[�	��GF�ګ���h7<xW/l�d��yvޥ;�/����c.�.z�v�v����d�h����`���c]>��v1�K��˴y9�,�`���z'.�8�Ŷz\�/�aLZ���Gn[k��4����vջ`��uۃ�r�#Xw\ݷc,65�N���T��=�F�v��y�:��6��%���Gtd��j^x��kv}�b�8�	��lcs�����m��[���cxޓon�<`X,s��5����(�<���6��M����vgu�`��u��vx��7�\vv��N���R:�v��6���rqj�Fkm�9����¼��i�^��I�n���H7�4a���mȷZ���)`�q�vۦ�[z:8��z1��ۉ�o���|�i�:���^xѹ����]�m���r�q��\C���=e�۶�+��Ź��q&�f��l<{dϐ�v��F�pn�'S���ڌn�oBu��zn�v\����������d���Tl=;g��<�c��7p��չ�qo^�9���չ-�
�o��s�v�58�Sj�!�痧��#��m��7��A�aس��GA��O��gn��=�����6�!��v۵/wLkvw$=��
��=����u��B�'�j-�8��67p`ևv��`ݵ�c��=��l���q��ӭ�4c�E�A�9���;�_��qU����^<��"Npk��kc���:6C3mg�m��Gn����s�v����������t�q���̏%��ۙ�����u��eL ��h0�m�ۛ�fMgY��)�uOaw\#�1Ml[]�up�kih�h�f�ˤ"��7&5ֹ�6�s�w=��9t4��m��=��o�8����8oUD����dݹ7��.� �և":�z��nuË��A�۰��'�$ɚ�6�]un��շ�����0f������)���I���2�B���&M��{ܸL)�]�)�[��;u����E.]zݘ^�X6T�z�7�����*ݑ�����]v9!B�t	�=n�wOc;��7<��y��ͲGT8�u�΍�ؼv��M=��<fp�'�����'ۢ�𜙡�:��ɛK����t��^���v7�8���ںs�s�i�xt�u���*�n5���M�zNM�C{L�qv�g��	yUlm{��,�ldB� ��
������4K�!��ۜ>w��/�fF���������}J�c�s����ʘ�F���9�7�8i�(v#Ǥ�n�2]��a��o����Q[Vݺ8��]�[�X�d��p�`��]�-��5s/Y5�m�6�G;/�<Z�nW�ɹ=�e�y���3���n���3��۱rjHgn�.ں�9�ܸr\��+�ݨyƉ�m�R��Γv�kr��=k���^0G[�÷Hm�C�O<q�}�۷���a<[��t�����ڑ�ۋ-��К�4�6EOVm��K��r:r��,�3��zB�\w1�@gT:.u�)=s�:�sq\����n��p��ն��z�#0��'T795��볃�g�-A�u�w��m������=�cT�`yv��t��#%�ŨN9�^]Kc�p�c\���V65i�ے(NR�$��N76 ��bŊ�i�t{.ظ2�9��M��e�ݹ�X���<��<k��ۚ�7[�5�<ް;Am��μ���eܜ��;X���7��x�6=q�ۮݮ1p��p�ʺ�M�չͽ�s�k]�E+�����v;[eWp��Qч��YޭǠ뵎:���V��
��:�3�cnd��iELwj+v퉱��v��n�{d������n�qǴ��[:z�8�.�}����΋<ٴ��.�g�#w���	��n=y�6��Ǝ����b۰�ۘ�:�0��c�뭸N��6ͻNl���9`�3z���x�mC�Ⱦ��������0��{��������q�K�k@]���$n}g�l��|�_p�v�'qI�|��y=���q�n][\�7�%N��O���1j�.3���v���Ŏ��i����1b9�cwu���ܺ��f�ay:6��]�݅v�ڭ���۸����[ٗ�\��&=�m�p���l{S�Q�0��Y�Uh�sk;�yrw)��-�\	q9���Rx���+�n��<T�기�H�c�N�nw�qr+Y��g��ѻV�qn�Y�9�Y�wj#.������y�������'n�;S����t�װWͬn�秷;b1�1�)a0���uNA�P����	�(ws���ur��S7�qn�+����<v�8�/v�q"�m�`z�.�箫u�E�ݼ��}�}�',��Hɣj�uk����g���L�����g��Y�Cz8e����p1�{Eq�Q�;;�rODi��4�[�ڭP0�v����U�2r��8�z]���s��45�q��q��_"/ sfn�gZ���mp��λ�<L/\�1���49�;n��k��Q�[��kQ]��S�{e���� �z��Ÿ7���E�WGo\�'Xm�r9��M^ZM�8۶��r{k�n������-��n�mAt�moe7XÊ���^wm��F��5�� ����W�n�:��vq��v4\`ѹ��s��d�`V9;=6�%K��稖$�m�(W\vݍ�;'g�6��y샻[g�۸�w]��';]m�"���O�.����Z1h�{=��gr=a�&�	�m�{�;8>�vᓜ��2n��K��2�xj��{Y���ݹ�'�́<�C�X��� Ar�����O;��wwx�㻻���}�    6�   `�c&� ��H    �)m8m�   ��   �        �l  �     ���m6�         �` ].�W�x�]\�         �`          m��2�   m�m� 6�f ��a�-ͬ��ۨ{!���f��^�+����(tY�����Jg����㒉L����v�4�]v��۰�GTg�� �g7f.�\q�xg���>
M���a����}V�gu�m��%�U�"q�%�X��n�vێ���[\s�S��ER���o;`:7=N�f���ղ9շ���R�vK���s�ࣶ� ۸�z��7Fw[�f��Yh9�>]�#�Zw��8�=�1�xj�y���9ps<����oPKƱvT�����9kKl�uֵ����y�D:���y+
�[���F̴��E�'P��K�q�=���m>�������c�k�<�����c��x����8n��D#�:zz�;�<�8i=���Cpy#m��֙d�>�lx����n�8l:Fx%�
Ld �v�]u϶��q�\�Q��ݰ����.�2��+4Ջ4qn�wg�g����9�Lg���$uو���+�^���j^�nM9zФxնk�-��S>�z�U+q��ˌA�;=���&��A�rU��ǅ7A�=\�m�h���Say��v����7b����x�����[g�k�{��h�S���;U��rk��[z:����)ƩC/=[5n�T���볱ηi;mݨ}�P��>����;n��\m�v�R{��c�b7 �����c�� ��lOm^M�<;�Unod�bA��q�Ö2�d�ʻ��ϗ'��n�t\hݱgI��m�<w�κٯ]tY��V��W!n�A:0=���΍����!6���ؒ�۬^���{����}��ԫ[@VĊ�m� �Ŵ�u� �d�� 6� �Cm���G(A���7�z�q��kmvE����]��m�f����;��GVz ��r�8���x���a���u��S�ؼ��*�n�}�&M`q��=���Ļ�E���d���n����Ÿm���!ݸx���[n�5].b�x�"������s9ջ>�zb�E��r��"�c�x����l��7;`<=��Nn��Cq�n�b.�/��_����(-��Y���K,�h~��O1��v�����	�KrR�O�m��}��F�K�㎘�m+\��&���vö������	��E^�m�7�d�����Vu�L��=��o�˛>��f�5�/�A� £��m��~�o��;{�mpc��g����V��r�Rfҽ��;~9�ޗ�'ye�nF\��_b_WM��ɇf��j�q^>C7�dq/?,���[$�L���=~�;��\,j�K�k�zź���[<D�tu%a�8�7M5sv���[qmzL�`aGN=5���������p�ev�&��\��@u�2��`ޛzܔN�_!3��B�z������½�6�x<��8<����ة�AǸ�SN�`I�,\��݀K{�r�v�y1���ʬ�U���1�㎽��@��sn_V�i}�NH�2
l;DF&.ዚ��f$@�h�v�TY��}�̮L��c��B���w�H��S��q�-FԌ�ڂݤ)��u�QV�P5u�i ��\���~�&T�(_`����]]3�Ao�G	)��Rs	����K�����p���p�Tnul5�t/$����MY�/��Qm"��d�A���6j)�[���睻I��eƝ�ng.z*�y���Z9z^:�S9`H�?\�E�؆ֈFox����Y�Oz�V9�=�A�g/
8 
��#0KO��˦mn�˛�g�z�l?j�<|�'y��2��&��|�ߵ�K����D��F�nN����}�쮙�-t��4o&�\���u����Y����hl���z��V�<O2�|K�V���Ӻ����:f\uܲ�6v�>��X����}��bp�⍥E�u77~�ͺ�0�	�OuH��,jq�Ox�E̫����[Yc[�'��.�De��1i����ّ̗O�*�PCP�'t�C:ƌ���B�o�j������vvو;k����Ctv͇\cU��RN���"���S;��M/&�N�+0|�����s���qd�j��~�fis�܎oi2d��Y�0�r6�%E;z��熉��)ܾ��6��4�Ǘy�p4����t��6���M'��@�N#�`�G������b�&�V:L����:����x)�a�S�� l��,� �/�=���d�~��J9<����5n���L�ݙ������/�\Ա�r�Qk�Ф�5��r��n��|�����*�T7vh��S�wy�������y����;��`I��m�䪾����X1�(1Y]�%j^	@��b���?"*	�2����h#�iU�ܐ��%��&MWZw��G�yv=���#Slք��v����5�?Y$P4@�	���M�^��a2 ��nfB@���}�I��AE��>ݏ~��|��`ƢI�Y�Kj�ب���u�8�RUn)������2ܳ;��'�jf�dVP?X��2�$t��x�!>��a�bտA����99G��b��������D�
�^Hp�C����xx�c�;�e�!��!�!��R� >��/����m-���"	R2�jx�l�O�Vd��������5�3�fy�zŇ�ណ-��aL�Gl�ڢ�-��p�f���8���(�]�1|,ډ	�q�v�g��ެ�f��=�{ !�lH���   6�t �����4�om�   8k� mb���[1㋛K�t"%��{<Ƙ��v��p�=���ö��Kg��Zݻ�4x�q�jN�z�nI,\JI��2S�1��c���A�N4co��N'<vc�sOG=�_T��6_l<�g�`���u�'�xw���M�4�Ǫ:����6'�Ʈ���+;D��͇�S%�U�m�+����h��˜�xx���+��ސ*�B]��g I� NZ�z�'�ާiw5ʕߥ&;�8�^���o����$w,Y�>�U��� � �DnV5�O2&�]*��,*#7R}�O��P-�6&�si��r�4���$��
��{����A6LK� ��3޿/���fd~��ei�������~wP�?"$��)�>� ��"��ǳ[�M��'n���x��i�RC��Gvv���1��о�U|��A�N	Q#�C2�K��<�y<�Fy3��+Q����9�/.mi����<}��SA6 ����h����[Qؑ�ln$4�u��5��9=�Qz�ג�割G,���߯ߦ���~w�^0\i�;�r� f;�v�k���ۛz-nZ>ƗŠY*F�ifF�(ٿ/O�H����m\+'�"�{�A�j�Y�m�Rg4��gݮ��/����X)�Z��kj���"�#{8�Vz��.I��%�aA�l�Ͼغf��(�7�QC����)���r�]�.H�+��>�����]�סasĉ�m��e��4�z��^$�A����v���ҕkg��%V�X<G���9��q����s��Ԙ��S����e���9d�	M��~D0����ܺ��E{�Y�ym1���"?-���r�r�x��x�d�M� f{WYy�vH��(c�`��p�5�mc�^�DGk�Fˎ	h�4ۓ/��5[���T�z~y�	����=�GW�����C�n^7���XV���|H�I pF��4�v�u�}閒���L���zͭ�#>��.�������+���:�#�� P�$��o0��!��%�s|<Ȍ�}�u��+���:s�j�"����rm��Z�N���A��d"5���ȭee` �V.��.��[�3�����}���U��Gk0�����D��H�S�O�����Ѯ�D3�r;�9�Q߯�ݼ����l$
Ʌ��ʾH���X�G�r%���e�6|��ܼ{�֚9�x�N.��|:�}�V����jS$ڷ\qնҌ<n��c�zwf��Қ|����S�FV�zs�hsS�S�rłF{������&L>����/Q~dqU�랿Ox->⦺��HR {�W�U��j�0�ݨ�y��gY�k�_��.���z1�A�{��tō˹8��y]T@�F	%�\��Ȉ�K��V�j��%�7�&�M4�4-��W~�JדWR��q>6�QHZjIe>���ws�h����j����p��d�W����b�2���]p��xl
�;^�Y�T|&b{������&��ﶦ�Y�H�������3��c�����5���&bj0ԓ;y�{����Y��Y�y����Ǳx���Tyc��Ӗ��C ���8A���V�����8��/k�snj9�<�N������ݞ��%�M��'j.%Y���������?|t�+���7��^�6���-�_n"��������db0�	���e�&���>�y���J��	���2Ӹ��"��~��W�ֶJ
�ɯ�@�T�"33 !��K���-�W��2�:u=�W~����!�v�C��n6�ty^��.�cL����k����4��;�����$^����b`�L[qT��|o�)jފG�i��7��_O���ǒL���X�<���c=���"��#WW��>ٗ�g��`�i -STq��N�-Q�j!0�����{�_�/�;�?<�= 8�6ؑ�h �`ڐ�( u��  ��`h�%�5�շ�_=Rw|R]��j�iu����70���w8��N���틤���Gv�4�T�:�Ɗy�:.��ǚ�9���b��&�ײv8��8d��5̜���F�ˤޱXv�v��zzf�z�5c��m�oZY��m��[��m�.�[�8�k��u�pm��c�"�횾�[�eZ۫7\�$���Sx�uf�5�y�eF�\\�!��@�a8��4�O�OQ���l�+o���m��ye� ��>7V��#�L��^�"���ni�&u�ݱ��5��m�]{;���
��]�b��=�<�鷛u����[Y��� �P(�Jdʧ�X|Fz�n��^���g�e���&)���\����0Ӻ�L̢
��fs�r�R��/��+qށu v3���u0訨{H��g���P�.�#��06X2$�/�c]�_�X���+�5������շ��F��>��'��q�$BRRC�����O,kc��܍˝����%������ۊ 4�2�Aܓ����{��D���6��$g�o>�삱z�^�y���o�xz����������`oL\�g�iF���2���
w�U��o�y�
�L͒�e�ޑ@�N��(0;P�t��%{N�ȌV�N�<;�Ң��3�B��l�nŋ͓��;�Y\:�le�Wc����>� �;�Nvǧ���}/}y`9��%���R��^��(|n�)$�f�;u�� ��ѥś���񸙾��X}��W�ez��;x��oh�){8E]�I�M�8IYI���d\ʙ���z�dj<�bG�N�/0B>�JX;���O	s5��U�j'8�Q��7Dnܶ�<bĩ�8{n;q۞��f��R�4�ʔ�$����+�{r�p�{���	zG�ͣ����^�-�|&�h{��d� �p�XKO:��_m�e�ca<�8��w�uL����ϫ[�3T�\�anE@�nL_a���L�g>���k&U\�C����8��&F2�+G#N9�0�R��l�#{fc��������X�#c%�/�C�i���Q�e��p�[7�d�i)��#�=��H)�m�����fB;o]������iZ�T���8� ]˰]b;�Y�y�J�n�=�|�T�Le��zk�]9VҒֵR��
�=�wu�t�mf�[�w
�B��ՎV(�ol_wV�ʶ���i��t�-�UvB�}�u�y}����>���%��ꁽΙq[�-U�k�/vL��Gޝ��6�ݕ�έ��*��b9�ӌV�%��vz	�uu/0��ܡ}�p��O9dؘ�˘/.�j�1%*73�R�]�B�+�]�VӪ�s6��)(�	f��ǵ8Z̘��6S9n'��cA�|f;8.��滓wm�8�Lݲ����',|�d�.2d�
�d��WZJud<㻼�O�f�>x9���h��S�n�*V˕�˥b䃖���S��^�ݻ��:U�j���W�Ɔ<vl��ޘh����������/w�no�w��z��ٖ�wXʭ2p򬗀X䥝̃�5�t�Z�p�D�+�V�5�d��{�����}���UǧrTf��fe��3Vrq�c*���>h�ב���}dR��#u��"(��]9nf�d�E�TrP�:���վ<�æP�eE�D�N�{�}�M��GbLd#�#�[	��;Ci\�2z{m�cz'/'o�_i<�5�/��0�i��0���4�y��"(����Ɵn0�����%�'��7��x�������g��!�=U���DV�"��1>�l�_>|�'�竬�HBsv�8�tv�=\�y�ge�_c�u�Mg�ڭ�wZQ�k]*�`�Ƣq��xj�><��~���K]��yR�¼���]�����H{ޚ�Cq��ݶ#��ؒ�q��y�e���OHF���=�&)Ĥ1�$rW0jF��m��.��i�,����(�(�ޥ�>d�H∣�~�c"ϩ[�)��E���Y�4P��K�lg0���y��k`�2�P@�M9(a$4�?{רϰ��da|ҷ�FQ�'�m�a���x�"�u�D\�����U�#F0��N���A&����p2S���B�;������]�4�FaoQpU�˕Ũ"��}���3�if��O��x(r�',\�"��q�.={m�ٟ�G	��Tj�1��>��e��Z��$"[��-"n�2&�"TV��#�*\օ|>5�z�E6[1�K���`M���E��g.�^�$�5�� f�b장��5<s|��x��BU_҇ujH��������p�a4GB{��3������M���a!�F�/K%RmE�uθ�vd�'N�@�:�_]v���Q��ݵ�wjT�y�|)s��!�_{e,�#�w��1�Y�%��$û�[�Ye�C���p��c>�&�n%̛![{���4��I�$�K�&�RP�!�0�G���Dɳ��u��5a��5p���C ���sDOo\H�Ĉ>�$�L�vD�>{�z5��\��
ؚRB�.�M��i�����FFc��QFM|�K~�Ҹu#+ؼ��<r�zPy�ˑ�&l���&�#�����ޛqpb:f2��ĜFőf��k�4��#�м����U�dA�Ӫ�d1���޻a�Ԣ`wM�l�$�"ޚ��Tj��}�#O+�i6EH�6�g�I 1���J�2}�XA�R�n���Sq�*[�Lm��k7w�+ȉ>� ��Ǩ#�!D��޸�a}dA�\P]d;=�@[���î�u�
��G��[]�ͰE杗[�E7����_�cͨ���ÁX[������z���} $H�zԛl   6�v�mp 5�m� ?�y ր�m]M�{a֚�B�n���Hmj��"ַ3W��d[Zw��}=��,�l�;��yk�����m��m����N�6{[��Okc�om������v�[��\ny���j�b*;L���s��g]�0woM]���"�v��t��m��uY[��������a�M��k+�U�g�Md�:���\��0f��%.C��#��ڍ[}�����HdeHb�I᧖F�A
">���,���'�2��Y�g��ؙ7�dS�e9h�?޷殉��f���G(5��4��C!M���M�|��<�B��o[o6e�����C������$�a1��4oS�Ia'�G_N9�a�/��O�G�J=<��^k�D�G
��n:AՄi�,��߽/�#-r�=�}���i�7va��2��Z,��qs��i}�v��G�E�fH}�3�*%$MFc-&�i�Tx�u�}:���b�葇H�����m���#�d=-�Sl�D]���b2��'�E�a�{�Q����`��e��q�� �}$S�7tW���F0�n�3N��˯��NXq�bO7�uw[Ϩ�0E�G���҉��#-B;Y�s3�&�n���6ԫ�k;��*ǘ�]�(wb�ZK"g�����Θ9�5m����Ͽ}]6y>�͑qRy��Ȳ;��i�o��jagȉ>���y%�vr2�da��>���aG���G��^��D��6ӈ�ӤH�ԅ�c����LB}�w�-�՘BE��cd����|�{��ֆM�ʄ��� �.���4��:�*ձ�t425J}��z:��"4�Gccbx�0sda�3��A6D#
4|�S��0�4酶��J���0BƲ;d���L�
�AQ�\�Tp�4�<��k�#&B>�+��'ݩő7g��y�\Uk�k72���v�����Q����%;F�Ri�%x#N���5���đJ�vk���d�$�[�S��Ekz�>ma1��!3ay�"{F��,��~W�C���<�M�?\%�4�Q�T���@�DB�^^O��6E���Y��?RS2W!�D����z���9�4���ޭF�Ef���7��Vҝ�Q��㐶��E$��\I�
�(�[77�}d.b�vۡ�㫪�����C� �Er�q�>!#�ߥs�#�"�=�U�B\�0���J�C���sV�1�aE>��Nf�!��m�C��ڼ��@�>�W4���[
2];�wTHE�#�!'�d3�������)�;"(�!B(�!Hg��Yn�߲[Yip;Q�A|ŋn#%�L��f�QUH�O�+�X���a����E�N��5tr3M�MqR��Z�a��D��rV��t�R����ٚ��6l_e��yG_�ja/�I�޶t�J��|�sda}/��2t�40��z�I$�K�6�����Q�UuD�ӈ1�fU��0E[�����L(�o%Ƥy<��ز*X8�c]7���W	�(�[W��
"�g�V6�$���c�@�����0��i��agXas�o^��Sh4i���ƅ(����!m����
�׌.:��u"�\�4�J��&�f�}AIY\�Q�jeW[�ֶ��OX�[=k�����;ɺ�z������U��%Dg���޽A�E�����q$9��2�z$q��ȗh2`�����ȫ޳Ӧ��xy�G�:�m�da!�J0�Wa��_���nH��IcO7Z�D{���E�4�g����嬥�҆8�T�2�ym�!I1�Ĝ"��������]=<��(><�6���{�r��n"}e��YDc��2,�u�I�Muu�����;��'��z��(;���B"n��]�P�!�ނ7�9���)�6T�<�0�RM$�ާx	��⽆e���q���=o#Sd�}Zºc"F!���L-�.�Gi5]ŗ�ݠv���v:��cj��=��G�ޠ3:Ŗs�_2��f��^!{�r��-UT�S4m���ɝf����%�WUe�o�*�.B��$�g�u+\�T��r��S^k� �z�G&&"��	�I��.7�h��0'�D�wESr"Α��#���_�$m�����uj[��]�źs���k�Ԥg)��Z|��ٽ�t��Pkr`��{����B,D�s���6U�c!3���OOc��X�����!eoGi��4�CGy�C,���Q	�W�mG"�(J,a�(�5!G�����hZa�޲+�z'ȉ �L$�V�葇�E�A=;�U��/C[=��~�J>��=E�4�a9
���fŞQy�߾�|�c�O�42\����vH�����!�i��=��̋L����äh�ydv�Gv�i��$NK="�e+L�q�Hb�%tO>�+H��֫}*���a���, �{Y��J�h�=^�\Z�.�*'M"��>e��]H"��$�nJyda�_(��ߑ�l�Q���_{�+M�w~u�us(�i�l�D�a���v}7��%�A}'
�&�7.���'�\O���3'�,8j�*��c����M�@�{o�HX|k�R9����V���I$�am������Zl6� 	f��   �� iԚn�Em6�O[6�TD͹Rq̝n۷+`{�rh�u���\�$G\vke�9�u�]�z��l�c:9j��n-�����o\s����E"7A���4F8��`b.3ݻ=g���Gc<���FPK&Ja�=S4�vK��xs+�����v�������=��)����䲍[V�\밍έ�Z,�<��jx�<k;���������w����<��wa��{����?����������m!�#Dw�~T0�4`A�"����2�L������6�G���i:Gms�|���̉�\bH��"���<��U�W0�{��t�|�Ǖ0��x���D�ߥ"�`�D���z�����r��Kv�i�&k���Q�!C9P�!RKzbV�G�B���=��	}n����<<[!-/RD�5)ב��GczH���!N[�E�^$W��p�,F�qICHd�8P����	��'�nZ��M�#z�9��7��>��e�{�oaK�y^��d�����:E#õ� Њ�"-���OM�N��q���CJYa�����W1Q>}aT��,�[ǲ(2a`���D�މ�G�p���=������j(��]zч�֙���p����;��\��;�i�zy�
��:)$�0���a�$B'�����<8I���ċ>���Oy�1���f����a$>����>�,�H���K~$"�8RI~#�{oH��i)I�	4�8��ݞ����ӗ�m5uԈL iE59�mAϨ����{e>� Tʁ;4�wJ��m��ES�/�%�B7W�6e+�oҹg��%�d�oV9���b,�<�Q>�&��^�8ϼ�'�iv%2D�qG���Yf�����gQ�N�����P��s�t2�asq���s���ls�3{'5��Mψ����4񑧐����m<f��I8����Q��ƃ�J)��G����f� �xޣ$�uD�s�$��0�����/c��(���c0Ft�b$��ߖ���R�8	r<ygA=h"H��~��梉(�.����s�Sq������*K1��	��h�M*"������<�0�j
�}��Ry4B��b@�]�n���OGB#S���li��v8&x��ԣt+$ֺ���д�,`��3�>��ȣ�����3�I�&������T��*���҉�W}-�4�y�m�/O�����mHY@��z�ӆ��W���Ɯ1�]������������dU�ȂN���K8-��@��$ɐd�R���Cz���b��a
��GĶ�rG$�5#4:	Һl󴅞7^��y�d��"�7�|��f;�2�w1��ͫ*f=�kj�]�-��}/�W���}�i���!�.�:;pY�/�S�+(e
�{�<L�!oa܊��I
�^��t���ߜ�<���|a8"��.��l��8m !;���F����0���B�-��(i��W)�}�^�a�ZaD��ióΘ�nz�by}DY�|���w�&
M��p�"r_:E�H��Z�Q#��>�Z���Fv;.Q<C�sD1#XQt���9��Y���'��(��3�:h�_���(O3bS�C$*յnz;jt�+s�-Zґۗ���0�kqf���ݜ.��{-�"+_��aX�D�z�Q���o���o"(�0�|�t�Qt�������N�z$_��!�i����%�>�adi���anĔ���@�
�_4�7g��}:y��k�q��X�S����-�(�e(�" �8P4`������X5l0����Ԙ�;�N{�"���(h�j�_H�&�\a���"�#M�D`�_�/�3�d�Y��5����ރ�5KD;�>r3�\OL�����qF���G�FA���� FFD���9/�p�����}�BȠcLm��Y����uuc��E���#DYBuR��\���rےpU�� ���Ga�0oeeZ���qn�+��u�q�`��#�r�S��Ʒ�6h��+�.�	-��1�d�c�������e�=/I�5���e��-vs��
��s#k�a���D��D��DI$a}��"Ϩ�<�O��/�9%�T�.9�Ei�h��[^;"�=�[r�f,[Wny�xKLnބ�W�i�B��dE��;�<t�爳D��]�4p�&�y��zw�|��d�"�+�\��]���,�:A�6M����h����ϟ��F ��2
q̌"I"Ξ4E1޻�N5���vc���[�qy��׻Q���Ν>�a�Վg�D�BȘ��w<�}�2k�<n�}D5����G�`NԒg4���5�QLף��ar	��"_�D��8�-�����ib�RsC�����Wu\�p�y�Z�,���Q�0ƣ����%�:��$X�ܬ:G���!�|D<�2Z��M�s���:�ޞ��]QA�'׌0fVq--��nב��e����#;k�6�Y��!RN)$�w��a���$S5��F9��.q>QTwg�}�B4�!���҇��Ya&����7�#e���Y�+�ۧ�\o-{�~l�u�tu��~YY��tiq�~a�����In5k����N>�9u�Ë8���Fºe�3i]���B��n��o&�U<�/u�v���%���ŎQe��f�|S+Mf�LJ^ќ��í�Z�݉\f�G�ggIܸ���wR��i��hP�qv�tv��B�^��T�G���k@�'�G�r��|�D��,[D� N���<�#��2q��7�B��W֕�:�W��r���i��"E]ݳK������d(���P����jS�"��P��镘���[�Z'sZ����]�y�9Z�,==�Bג�]fmuJ���t�<ru��͗/�Y[w��l�̆��u<']|��.��s�45b�+p-�ȝ(�b���-^Wn�iQ��ud̈́�sb����t�]�gn�͉�=�W+���|���cu`Ϋf�� nv�{����])QdT����!�՗�5��s����N���ᬳկ4�]J	Sx�-q>CtVM�3~w���Cn�Q����/{k{���w��w>� A��@�0}����[O怲	�%{�x��V>��ᰭ\���1X/0�3PB���VI��1�<E�4,�����W=�a":��n�8!���4{д7c���I$���      m�� m� �   i�����Z�7 ,0         m�        	6� �ѵl    '�\          m����6 5�l��ɛm�   l         l    ��`����0        ڶ ��6�z[�`<#��Ѵ�cx��`w]�m�9ܮ�a�C�mX8��!�2O�N�;lk�-��z��%�W���ȏ����]`�K����vڎ��1��s���㽩����1;�Լ����=���[�/[{>{��եR�G�#=����8�ӮGn-����N{u�8R�[a�8�ɫ9M�q n{#�n�`]��.��9+����&wl�x�g=��y�1;�L��Dݼv�O���d�8�BF]
<o���.��t�n�㶮m��|�<xr|�o��}�&/$��/nܺ���v��N�����اv��t�������]8�/��n�mb�y��t�;�.�'
���A��Zk��l�_Tn{q�cv�R������+x�ā[9���h��/c^|�앉�QCuy[Q�nEI����rQ�U�[�x���'C���i:�u�)���P,p���f���j�2�i1�n�s���;�\ra;;���O8�qs�=���B�n۝��v�n�p���z��!ٛNG��nS��4�[�Ź��ۇ4p����U�|���v;�ke� ��{uۇ���'7}��9���\tue6��ڢ牎9y;>2�2����[
�٪�qn�B2D�T��;�ϲ�g�6l� ��ՋM�ɠr���캃��`�6�n����a�۳�뇘[.=��t!�*�q��x��Fy^�ݵk���8��s;F!D8���D�p\�v!Wp�������������Ì.��p��ʊ�����n�:��F��}���}�<%�g����rvk�C��5\ H�lH��� 6� �� �Z  �oK�   N�j�U��y��AZp5	sz�.�ݺ��^�8;F玮֖+��hh��[k{p��M����@�{$:�8��C���B����n��ػq��v�n�=��h���q�7V���ym��n
��]���|����xm����/���kv��qm�&��F�˨���QQ׮��øj�]�Tյc=�%a�Lu����	l�ܗ��������-4q�Ԁ�����6F�Q
���\������Y��x�o,i�#H��1~Ͻ(G����leG�/Y0O9���I�M;���ơD���g�&c��!0"ܒ��A����몊Y8]J�g���d޲=���-BaY{�t�Yy�N�+�!�!\�P�|飚�r��?4D�$�I�xzD$���E3���sH��V�=1NdYh���$I[�q^�fI�r�����}J�D�0rx{��CME�'J(/��Q�Aߨ|;�0DV�l$�4�F�����r汄��ۤ�<�j�:���F���O�LޑX�"F��57��\��%�x&��$ND[�׎�cC��C�etW�I��
/|4��3h�>� ���B����cG�[��w_O�N������u��������MK���F{9�������ԛ=v�뭧c�sZNny��v��Pۉ��.��|t���h}K3�r$Q�L.����Z�{�}�Q�$�7��̃���q���#K��o���GԴ��<��܅6�E�܄��nKl��a��	#����#�

GF-��JHQ~��/`Wv,�9w3C�9f��{Ng�b�����)��R �����g���G�<�����j`���t���v\M(�0B"��f��Č6D��<�뀟�z>��E{t��%��#�9Ĥ������w����fu�Ԉ��Iv����8l�":β�,���r�^H�_vP��`0bPG��k�����M#��a�����)Ӽ=>�/b�:�D�����o={H�0ޡfR���P�o	6I�Ǜ �?zPýAb=�#��D�C��\n�ѥ��Gur�=���q!Q"NJt���,`�z{�F"���S�-p����HӤIsE���"�y�H��pp���/��>�8ۍ�Rd|��SK73�?���V�#سnsom���v�`��T�7a�]�n7ga/]��s�g,v˳�H���I��O�����"fݏ�6�>���2/�f��]�� ߎS�p���?f����ңY��Y:�����"X����2�q�3�;i/�󡆖�ˈ�G0��.��O��8F'Ӽz�C;�O���'ZȾ���#N�Rw6�s���&.}��^F4���S��ϗ,���E{��\�<��Z�E�,ߟ�*�g�������T�/�u7���JQ!K�Cx���r�3q��V9����w��^�"uJCx�ձ�Y���ܸ�T���n.h�$�
>i��X�#O(���	4���@���suCfsDȽ�<eƆ ��6�hi�;�,ƾ��*ȭAlB��������\�@�������I������y�+o"�
̙f��.#FHܒ$��t��;��,U��2(���D������l>��Ȝo1�Q��8��B�"Δu�M����ʣ����>:C�3՝��	���O$�ZڣV�=X�x8���ll�%��;{t��N.Ύ��v��K��'����l�$+f��s!&�(�L,k��'���f!4};=�!�O6��s�C�A�1���.��g��3OpC<��\Hn<�V4�!{�m�'�36�x�n���}!6��l�ʔ+[�E���^y[� �"���"���z�n��t�>ԍ�XX;G�'���F��&r_4�"y�(��ϯݔ:T0��H��pO��I�(�<���"���8E��A�'����l;�?��"�3����H�䡤_ʈޫ���A�y����Y�^�i��S>���2��Q�g7]7'�c
=4�M[ D�ebAk����\e�&ZaIN��bí`�蕌�s��׽c���guV�J<��iΛV�%^��?q��I�i�H�y�q���H�Ε���ׂu'��ƞcCO(�ǯT1a�4��|��o6���V�ȑg�l7��~މ�ĳ>�V�}��E���c۷�we�՘�i�YD�i� :�v_k��<��5���x�۩��쵮|G&���)QIq�zB�ZGL"���J����BZ�_��+j�6f�]t~��lPy��yl�zD�v�A}oC��8}i���}�]�ۑ(Z��+�|l�/�n7�8��ҌՖ5�	!�.��E
jf �	4D-�NhJoR`H���Wu�ɳ��*��k��l0��������nJA�okH�/�=#�Q�>��E��\��S����}�>�'��'N\�V��2m���(#�!#{�>ؒ�HC�H$ �%�m4[1IY���QSR�s4��A�'��'����L�����0�H�u�`r�)�;ky���Dp�D7��`'AF܎�t�K:x���tP,C&s%�b�`�s�3q�e���rEmr���,B(�7��S��H�M0k�e�;u�&����x���;$��wOY4��9-6UG[G�B�f�T]�.�$�D�
5+�e@![I$�vH m��&ٰ   ��� 'Y@ kx�   ���ua�y�Ps��rٓO����آƝ�O`͵ەq��d΋U���G2�nÇg\��M�[��vɒ�Aҩk�9셁�G]�P=N9"�{�k�!�G�c���6��o\���N��J�:u����n�ֱ��햜.wG;��N>���#m���ڦY`��4[*��'<\�\v�݂ۜΜ��b�N/�vӣ��n�k��P��_�~w�[������w�"񤹦0��ބ�}�A��2h��]�!����Q}E�\O��#�'�DCl�DM$i%#��C�5��R�}�'.x��{K�N07=�du'Dab�����q4{[H��4^m���딼�y,���Xd]gf^�n�K�$Pf"-����Q�z��hiu��;0EXa�A��zw�|��e�kZ�{�HaDw,�%#�CD/��)��I��:��?}X�҅��")8)�hV0�da���%�4{{"�S��:aFY�WO\P��8I���lOq��D"1��;�۞y�O��Y�S1Q���:�\'jI+���<�(���=���=�}&'uC���謉�$d)dD7v1����,�d����;/�h����z�W��S�F�2&[��$M����	���u����u1�]����g�j��/0����DdQ��N�!ך#�8E���3E�H��L(�[�B��cda��;�!﹈�"γ���\L>��Y�y��"M��	$��"�2w���U�ՂuTt�x���~���W�A"fh�#z�
�uh+��������Ԡ�ؚ�3H��j�&},W~ە�!� �@�\�W�(5��Ha�����#���L���>��e������ f8�f���t���7/�+�zl���������a��l%I}=qA��&�D��y�+��I��"� ��[�m�jH���ܙd�!�;�Ϗ�7Xc��W�4A:ޢ�-eoYBF�ri��Q^k��a�9�T�#m4kj���zDi�g�ƴ���y�8w%��BH�\�4�0���EO�+�Ea�U������]�f�k9b[�������y�Q�Ez��B�r��$�2����������՘���q�]	,F�"ˎ�gi���z� ��U��k�[�'rDƁp���X������?��ii"�r���y��Da$z�Wt�Ć�{9
<�����0Ȏx��a�#R���5�6�I�R�f�!�7�$پ�Q>���L��`���E�fC�r{z�0�$�a>x�瑇�]|q�y�Vڇ��mMt�NB�e�#�n��Nj�؇��l���	h\�Ϯ��qL~,�[1���	����ʮ�z�o�%EH�:ͱm�j&K=E�h��0�ͤ�)P�t��z�s�M.�s4N�޼��#�g_\N�88�L�5��9Ф8"rD�e�0t��xGOc���"7�F�Dq|S	2Iy��X޳Oo�����4}���M��l�ڳ�(t��P�d|=�̜�nF�l4�t�<��D��z�Ԉ�4�������m�>��\���|H�Q㯧z(a�ջ�F0cDv�'�GS'Z�O����"Y�$�K�!�9	m� -�/Eq(�g= ��g�<]]�Y����sՃ$�S�&L��҅�r>��s:EC��y�F�����=P�Wb�Y�1�a;=�"9k���"I�x�o<��f���N��Yw����0&KL!"RKzt��*�F�zP�����6�G@���3�l�!k9�e�!��CO3#A=u�;���*�Z���!����$W��8$)�FIcS2F�QQݑ^�MDn�sGuc�1��.�t4�G���N.����|�}Ht߯�*Z��Y��E�z�"Xp"�0)m3�L$�7���0��ф*�M��>�7i�k���3�>d�O�`��z�E�9x�V��Lv'�e�݅�V�ޱ}����dF;�0�����V��bu��f]�^��.�rz�O8�$�4�>� �=�o��Af�!��L�����.Т���4a�5-�l�D�M�8ID��?Q�>� �
��/��]��3��X�L�#�������K�Y�6���z^Ύ���iݩr5���z7NG��Z�.������ڃ�
NTq�H�,�G��/�/��%2���X�#:yD���>E;�e�-9��A#݋�X����cf��[W���m."!�Y�~1�F�(�$Y�M�ޞa��8�l�7kp�ZQ�x�rDu^��D1���d�mqʯE�Xт
!�QǮ2����:��}����E_��M6�E��(c�=�I�:d�jn޴�B>�f"K�N3	"$�z\�6F��Ƞ�ޒ��{��Q��iE<C��L\��'�n"�eIE�������1&X�`�Ȇ��~�$�c	.H2��ĆƲ�!̑�;�>�$�E-ݷ��_/Nf�hx��li��I�{�Tm�D�D3�E{
2|���讉U0<��bMY��bi����I����\���o<��˷}râ��p�E���EN�C�ϝ����t7Qd���K�71��lWA�gkT�RT��&��.�e.O��[�}]
� d�I�7�N��@   v�h6C� u��m�m� � �����/#E:7�m��=���g8ۑ�I���'n��Bi����Z��s��M���x���';]���s���v�s�c;]z-Ƈ;sayzEKq�ۇ�֫-����αy�'k�]�îwZn��=��<u�:���w_ZV�c�K,Mk�;WM��ci!�É7\L�^V���.�%+�s�y��o]jl�`{lCa����I	=9��B���h��3_����n��L{u�=y'ؙ���5��>��>�k����M]���f4}da��v�����C�E�#+��I��l)��F�2*=$��!Z��y��=�)��L��`��E��#�����'H��lc����k=!5�z�|�$:B��[c�������I��NH�	8�a҉4QӠ�"����w�H�HIb'��$k���Xh'Gլ3����H��CK""ky�a�ŸG�Q;����6ْ!I��Q����}�Oʞ`��8�CjQ�ѝm>��EK*`��7�����ޢ0����ѳ�AgvW:F���xyu�w�q�c���-�CH��'�#i_�Q�#N<��H��}e�E	��y�l�)�4�v�	Q^��"�.=}��M>�aK�3�~��H[rB�p�ې��5cm���uڸ:�g�����M�<����#��0(��7#R6��o<^+<��Pi����24�0�3Xq¦vꉓF����8l�깋��qt6�#�n#��#XF�	i��!���f�1�Jm��f�Maj�����ft��������Oٍ�Ѽ���3y���|hwf���,dAr�8I�n��0\��˶��m�(g����I��O���L�u"Vt��$���b�#�+���&:��Sab��k��k:�h���}�^Mw��Qi0ąI+�p����mOs�U�b�#�1LͽXƽ�A󷷝K��$:W�!�݈�0�Z莘�%��>�g4}}�Wk�A,#��X�E(�4���o^�(�e�5Yo����ޔ�A�e������;��}�N�1	�����72���FȚa�Q�}��"�S�`N"�q��XE��1���#s���M涎��2V�onn
��>�$����W"��x�bM=|g�D�#���졇�+���]R�,b��!�v�-YÍ-��GQsچ�N9ţS�`�<,�0t�:�s�t�HD�$F��D��.i�l�W]�#�\a����XƆI�'��2�GH�.){���<q!��Y����q $��χ�E��Ԇc�4��ښ�4h�B<a����k����ԭ�F$�k�G�\�����|i��B(�@�mÑ�28ՋL(!�&��=i��(�FDQ�d�����(�<��.ګ��M�Hy�b�+,�e�w˛ѝ]��n�a��},�A���ŊD��\��j̌���z�Ԑ[� �}۰k�k6/8�غ��+F�bL�Ydx���9Oi��ȏ�T�O���w꛻�����S*XH�E��mmj��7�Sxm��5guk�w�yEՎ�&'rl�j��j��3$Q2�c]��Zw����e�wG�J��d��`]Le`:����x����UwR�w���Ю�Zv ���e�p�v��]�1�r\��IV�o*U�#]��|J:%�bfZ-i����7�,3;*G�+DK�!�>�Q��-۵ �mhifoh�V�YYQ�܋�}�r��)�V�y���֮�WQ`5� ߎpw�=ue��aꔰ��m.}eK�N���o���%a�������s�K�i�Ӆ��b��J��GCn�sP&�Z�0�'2���\�Ov򊙦V\jb� rP�@��}��ZG9���`�s%sP�M}��5ٕ��!��kr��qq�wX�|�U�խ�2�S�x��b��nN���U�����e��:�N�|V�e�!���v��V�Zڈ뙅C��+��e�I;��hk���v�ۏo����l�(s&b�/嵔Sr�;� ��4��_@��R�0ce�,\�r�z�k�DԊ3"�8��M�w��X�:��oO-�i�pð�q������Ն�;������ä#i!w�ޟ-���_#C��;k�,ծ}<-��4�EHZ�����ӥ�his]A����ORެ<�0?��h����䡄t�d̙��,:;,�El�E�?fS����)��,����>�Q�!l(�Mn��t�D���U�Ѡy<\+��D�u��r�n�,�:���*b��g]�~?N��g�,��U�˹cNb�W�C�!�#b�L$�����"�]=CS��ڠ�/9�CO>hzw�dixȇ��_��Hb-HbS�	%>"�'U��������V�27��F� �*v�$rw'Z�}o]��ꘐz]E�>��Q6p�,V>��{4i�����my���D�m2��3추�|��>���z}Da�=��'��aFm#�d�Md.B�$iDIb�(�?�ƹ�:i#P��<3މ��2�A�P�ɨ�=���8{W�*�D4���<D�y���p��!��0���2!��`H�5ɣ��6��`�*⥤���T�Z�G_J����7՘���g�'��ڴv�r��a��Sv9�9�y荼y��[��FNo�e6ْ(�d���͞t�6Nt<��!9�	��/�ױ�|��!8�R8j����Z�C�����%�"����#�<Z���>�����dL����ղ������nYa<u�p��x;m���3�hU��d�l�1�ifǿ���s������&|�#�]���z��5q����P� �{)��5�H�$��.�b��1���Lv��N8�e�d���di�����F��i�.i���aI���]]�"'�oJ��o��v��.wg�3X�Q̉��>HՇ��;�.h�ȍ�#r:å8F�Y˟z��sHg�D,�7l�=�i���zw�&�����3�"J.`��m�k�8}$a�e����~�׉�"�i�#I�B�O�*ȣߍYv����p����ʊ�e�PoQkn��I�-_!�f����wg5v�t�ވ9H��!"Hs��^�ə�� �hH�t�
�|F'��sM��e���p]�����B>�4��������]�Q�t�Č>�a����W�e��u����n)E����v�rw�*$f��`��0���̢(�6&��t�Gz旎�vAYGE�ͤ�$���bE
�   [I Im  f��   @U+�.��:qJT��^N]�'&�e��R�a�p�u+�K�ru�mjݮ-O�X>�6g��%܎��g75�k�n����y�g���ݳ�;K�{s��|�ct��h�9�n��n�Ƿg�o]��v�p t'�����Spp�W-C�����{�=��t�:خ	�9v�f�h��*nCsnH��n�nr��ݓ�[,]��׸���9/u�F7����>n�~ha�L�ߝ�:��F�����>�$��g	��nX�y��1�y{�v�M��Ze`�A�.l�����k��J��9g}�����~s����w���e�zٶ�*�O��8E��ċ>��Ϡ�f��q��3�Q�.�$�gv��
��6,�*����f�hg$�JA��uH���h�N|=��"�X$ޢO<v	�F>"��o-m\F� ��s#3�Ռ��5{]��Ñg�=��������,�nԒz�O,�1W����uf�qCK8D�!�o<����s�qM�R�'����f��/4Ge_�lUD��4�0D3���~^	�0��.dr~=8D=�]"�����dRk.3}FU�g5�R��}�Ms"͘7��4�b\"�ý�tM(w:�6���0�q�fP����j�x���r�b��N��:�|�\r�Mn�k�9���ʠ����s;�����\��%�S���y����X��C��V7��>�9��H�;|�V�o4�6��s�X޽�Nd#��#��u�p��-��NI|Ӡ��B4�OLH�#��&��:.f��k/�ɯR=�n`�P���Eٗ�3x͸��\:��:��Ӝzm�1ǫ��Q ��'��w$���	�M7J�}�
,Iy�O"�w	h���'Ȇ�~f�}����G˟	�}H7D�!a�Pj��#ӑ!���Ş�$��Q4�!���E�2abJkV"6:�"��A�0���l�D�G�L��D3�}�&e�!*&Z���
!�]�˫���#�>������*�:��$Q7�0�8yG��>P_H���
�tb�}����;Y�&��l�#Sz���Y��8��
p��40������Rk~�L��A��SͶq�mHs�oE6E/���E	���`�j�&�u����#H�O�ߨ�����&I~��CP�$�ڴ�eWu�=����l\�"x�t���-G^a�^&:N8�r&-��)��ns��:#���!��L���Ns�g�H�@�\��Y��`�׬���c�A�4M�0��=0�{�+�"E�=��Q�Bc&�8�-�B�l�.�����u��g���{DTH�>�a��v�O"��e��zK���s"2��DY�U�hҏ�h���t�p�g��ě�H�2�iGY"���nƈ�f��s6{X9��&kz���7\�2͟�����0xN��oR۶��Yh[��NC��\�Uyg�d=SA3J�|��b��H���8`iV�PDY��A/L�&2�$@>�!��<�5����FD�t0�������ǁ�F��c7�}�̖#w\Y'O*o!:`����|f��(�$���ח��I̱GǺ�#�:h�cĳ��M��i9(Y�(�{�M�3%;�,�>����esҶ5�fO��"y[�"+�R��k6{��O��y>22y�����/�[4�r r�rB\���q]pe#[��!�ҹ.����d�r�.��qI ��&H��$z,���B����0�>X�O�vṁ�\��>0��葹0h��ۭ�
#�Cǳ6Q>��q� �"���~@�(�
D[N#��!E�Cqőf[k�B,�ݪ�`����v���D�!��"K�qz�r&ˠ�Iz`���܄�	�����zל�<3g^�Ċ6�9
e�͏�r�ӤQ���"���>�$�v;�D�$[f)3�,˰mt��d�L;��1M�G��F����^	=Q�BM����$Y���P�<��7�y��74�F�4z;���:qD^۝af�޺NdF[���'��;����.t՚��%�� ]�4��av��nh����.i�롆��X��tY���X]ʛ�n�؟Y��D�2Cγ[�3��È��������(�s��E�y���F1W8�>��9���V�f-����t�,�T�C�OX�s��8��b.w��>~�����4�M���	Mv���u��l���Oh���t����	�	7gl��0D��Ԇ8DqH>�O����օ�_ުs"Ϡ����l���&A��Ņ]WLH�G=�E����� vY���=���ZGJ=����>�[p��F ���q��,����ڨ0�=���#�p�d;�|�QX>��[ȩ�h�zo9��$T66x�"{�QT�Rc��wo�<�ĝ!?|��'m5#B[r_7�t�m"/�����m"y��4X�Ma3��Q�(K=��=�qs1����\��	��L�6\�u�>Do���<�o���D) h0�:�E�cQ�[C���D���#z�|��f"w��H���-����5�]��Dn0cѽ2�~�ڸ��O�c�2d�Ǽղ�(�J\p�t�GI:Ђ,�-瑆�%}%����5��0n��+�sjE�"0�gSȳ�8p�3:{�N�`�ǚC���>���ۏ� WYon�$��e�B�;hÕ%5���>�t�M7Z�d�����o@��zo'�����>@XӃm�   �khѦ� m�   h �kIْ䝎I��Y�Y�lu���ά�m̛�\ͼZ�O$3��Q��91�7"�R;�ݹ�p�(;�;��&����A�br�c�1'����t�[x�4���Uz���s@�'lѐ&�vT������7(�7[N؞��F��gsm�Oe�]�YpA�h		Ŝ�1Vwl�џTd��Ϟ�-��s��m]��K�W+�Jb˂'
�A�������h��۱>�����"�zbp�}Da����S�ȋC\�zrB#�"kH���k��5
�
,,��|>����a9
i�S��i�i,AT�d�`瓊���E�3 Y}f�_��Ď8EJ"H����M�h���=��>�%ĭ�]�e�a�Q���X)8d2�re�"#O,��޹c^��ϩ54D[�<�>�"�_0e?X��[qt���
�b1�)tф{p{]#}\���+���&��܆3RAXF�.�#o�7~�ڼ,G3EBNd^��C���7��4�lAd|p���{%5�ZF�ߵ������`��$�8EB��cC��	�
F�v4b���A_�t_>�yޡe����=����9�O-4���$9V���ޜs9n�}R�Hƍ�=_{�j�ʕ���㐶��E$��N�Nx����SM�b��Cv�̻u��8�랈�0h�S&�m	�h���g���bE8ޣO.��1�QF��Q^���KK"4ޑ��Ϩ��4$�d9�N��g�z��u$�r����!3A�`H��$a�cCM��۠�݀��}��N\�57\�����/e�R]u��&���՛�0Ӄh�.%�<���fP�>���w-�z樛L��1�&��$I� ��N��H�0���Fg��0�hrt����/�44"-��gO��y�,��/���T��w_H�;��O�� ��\�#㊆[�R��D9�:.xϬ�>���#bm��R�(@�I��5gH�XF����!>�wE����t��鋢y3�e�9.E��F�
'I�`Hˮ��Ǡ����:�-�q�ո��\0�2�1�$�MA	R
��Τ,��c��a�8k9��+d���4Fu�#<E�`��Ӿ���\�~�B�>�N�3�qVF��\�Q�{����P�j�v��B�N=��<9�{:D�x�T�n��j�'g�x�Ս���V�]*k"4�:]C�}��ާ_��F�I�6F3Z��Y͘�q/s�#a?��>�:�lH���"��(��u�����icA(���_y2��1�"j\n�J=�Α���޵�CO�j�5��1-�$g.��em�	����Ȭ��1q$0�i��gsHl��"ks��+H�X+��-Ĕ�G#��<�!�ʘN�`�a�rg4\�ۡ��#�,���&;��[M���D+��Zf���.\傡٠>`cCSdee:��J}r�:tv�m�j
�'���ؑQ���"�`�����[�к�Q���VB���a�A#�F��$�0����6�cH��YA"Ȅާa�tpME�������7O8hjqd��{01��ҴO��|���R,N0�;����ur���<k��(��-�U���W-�F��H��I߽���3�J"R�W�,i�b'J"���~<q���bm��H���	m�6�����ۇ��scZ�M���rr#���vY�s����j(�a����Ӈ�\��aV�o7�B�"ȼO�.H��B�Μ9p�4Fގ��4�!����ؘIl���5��0�:Y���D�LC���Q�(i�#5kB�7߽���.���O�&�r��76�z�D�X_�g;'�,���8DU�>�77�Tr��g�pw4�b�;݉��a�e��������l���c�p�"������uq�6��Dmw��=/ND �K!!b�L	�5{%|p�����MQ.'�u�$%�#
4��X�!�4���F�_{]	��l��"�s�@���8Ec9]עE]>�L�6��k��t����U�\�����q�W��`$c�;�
�˝�+yB�]�1	�B^e�j�d�0�|���N�H�aI
�����[�Ɯ
H(iҍ�iy�{ֺ;��1��O3�ɻSL3��]�\O�>�$�2��$\c�7a�����NH�oa�Թޟi;�|?
�9a9�I���k%��$^�h���.�2'L�88SsІ�q���6����C�|e�M���r0�Ɛ�p�#	"�TH�4�}$'��#h�[w,Ԉ���!�l}=�E�:x�"f�8k�g��J(L���rU��JuƸ��g6���(f3�\�F��&B�~�����v�'�i�~_�x�n��4�CH]XY��z+�a�G7��}|G�$yvEW�&`��&I1�""E�8�F"���B�F�$D�j�H��O������k��B���(�,X=3�g��%�ID!wV�j\*",����!���V���V��Z��(����y�����'ɓ�DQDQ���\P�oFۅ�υƛ���,�C:|]�\��~eFb04$2�j
�Di؉�����|��89���`�|�5��%>���K'��pP's�"���K��Zo��l���W7ogFm�x����̧�ͧ7�Y�)PO+7Oݻ��plfṀ�iW/RP��vuugK6�˔j�<�E�[zvA�sl#��]�N���©�2��W6�}:u�:��ܗ��sE-�Q���$Y����w���*Rʸ�76(�9���.���ޗɞ/{��L)�iY@���2e!�īa"�rQ��Z�|�P9�vm��ȑ��Ϛ���ܾ��˭oT�N��S_Z̪��;mp��>�9�Y�%ޫj#����M��v��6�>|�}��:� �:���v[F.�Xε/l�
;�6��C�� �r����^vE���+���F��v��zJ靈��:�ɐ��s�Д�N[&V.KN<��]ޭ��V�r�������|jn�l����H�ޅ�3u�p�Ay�e��q��.۱/�]�����I]t��U��J�
Q�6z:y����`q��gkh�+.�^��9�y^�*���X9�M��;�n�˓u�a��� �ճy.����R��y\��n8��]�b\�G����f�u��V%��r׿-��9�)m���X�p�h|�,b��"�sKK�ݭ�0�t�:�b�;��kw�hwf�e�B�k��ۅ��u�h��O�S����ϧ�������`      �lm��   �   4P /Z�n�$�m�        m�        �k  q��[l     v�����      l    4%�U& N5�l�m       �`      6�    -� &�kI�   ����  �@K���{;��j��/:s���,pDloV^�[��]�"�*�v�=�����ĝ`���<{*�a�=xH�dEZ,�/s��{��6��uȽ��r���Puv6��'��۴Qٸ�ghn{z�D�wΞ���9zM<���%�����q[ynϫ�Ͷ�gut=�0���GnuF7X㓓GOm�g.��7BlC���ܼmۅJ���E��c�g������8�I9�l���{�2������B\�w#���AN�z�h�ݩ�C�������}l����[�wm��[q�շ	ѩN�l�nu%/]�%�)[�v#���b��:뮎N5���Y���ջx��b�9n��]Z|���!�<W�K=���rca;qՉ6�&�6�%<v;���\75�A����s"+ۆ1q�&9v����8����>��v���'\�d�!gZ���;�t<�����6y2;g2p���t��mݗ\��ݱ�.[v�{1��f��FA'�m�aQ�S�:��T�I��O4��H�v��ێ2����v�q��ルtv���7�sɇ1�`����qc�v�d��s�vlby0!=�v�m��Wsi�Fܢ 7m�P<�y���6��1Չy�M��\n� �v�xws��}ca\��2��[�y���&��P9�{.��:y:��ssͫ�j�[t-���c�H1��K�z����K�q�6�9�2v���1vK���.�J3�b���W���\��/=Ͷ�.�n�ػz�˘��T5�b�qұ�Խۦ��n�٧&�ɶ ��[[��   �d0 ��  � *���E�U�Y㹎����:�nٷuÓXsq����ǃ����]���ҝ�n��g�zR���J8U�i�n3͚ݶ���{y�\rv���U�\Lm��nz3Nx�v,/	�8Ƣ_n�i�}���aޱ�f6��!i��y��l6�q]�_��VW%�j�g��Z�wN�}��M[<��+`�m�sw�n�9{c�ӭ�frA�����A&�~��\Qr$��ׂ0��<��$���o2��To3�Lk�g�)�>DWw�+4������,d�2����䌴�i�$�!#���{� �d꺲��DV�qG�Z�B|��$������,&�(�Ȓ����v�oN������Gua��L��fC��^I���0h����H�bD�8ޣF�������l&��7��`�0J:bB#cF[Y�oD��p޲$�7g�<�[� �QH�;Eua?{OoB����lWZ(P:h��Q��z�B��6\&���c1�H��DY��ŇR�n�s��b�AF,r;�8�Dh�DЊ8�����{�ő��d�CH�DjoQ�v�+��p�@�F��b�E�sȪ�wa�i�7�R�A�������Ȃ<~ֶU��l�n��m��ݻ:�YSua^�_;�Re�9��Cqɖ'r`��!��=>��柍�iI�6����0�5�w{"Bc<xl
c���`�S�g��0ޒ�1�	&J&H���"#H��]��.��L�S���N�^�l�rh$�a��8��ޝimn���_R�|	���r���RL]���Q����28_������'n�°�(�/�Y��~�CO+N�D�=|dI�aMe��ʽ�A�H�v�f����£���>��<�%��d�aQ����}���v�>�a��H�H�$a|Ӌ^I��"Ϡ���0�a���4���z�A�'���P�e�^dHF����l�:�בh��t��{�\��dNc�0yI
�;���}�x�ϓ�,�<>�u�$�%�T.&�nK����:yd{�OB0�l�l����։��OC��d73s
!�g�W�ٓ�.z��q��Z��#$Sy��z���4�\��&�rmp��ѱ����a3Qu�#����rq�;m��k�n��5ư�JN��8k��㇏�Y�{լ�-l)�V7�����X�cg���g\o{��!�Ƈr35	�a�<���F�>��z�O���6�v>��4:h��p���.�����A��	>�V�82A��ԻD�t�37X9��Rs1,��Tޥ8$�Λ��Vks������&��{�G��p���_�U�>V�e0r孷��	�-0�a]S��}*��;N�5����9>y��@��ubý���8�Ht�7��"�[��ȹ��x����UGz�Y��sȮ��`f
�I�z�	�k(���"0����ffd3�0�05#��<�in��-Q�.Or��~DI�%3�(w�9��d�>�'w�'�C�#Z��[;�)���[Ϥݕ�">=�:y�}^����$�	L�ZF��:��\A�E�o�;��P`�,�E����Ӗ���h�,d��~#!�{]��ce�&`���DYӇ��Vy�ܱ~^Ǎ��jHL��T9V���:3F�m���8��5�yɪ�1�y�GP����i-tg���(��]����n��Ə��z��a(C�7�d����N7������;�Gў���x�>�7��C�A��𯆴�4��I�zv�I{h�fz�a:��s�w�����DczOi	[����6p����Э\�hid�m
��d�p�m�Q���4�t�F��%�(p&̑�M���d�vB��D"$�^V����V�f�܃�3x&H�a'�"��z�F"�.��u;��b�9.9�Q�4Vm���S�m0�x���5���"˦\�����FP�������&���ot&n���٤e��l�w;�t�n��[x��`=�T�t5��F��p�鐰JfD"�9}�-{	m�l��L�#�!v}�x�"O�0�jV<fS��4�2�$e���"����`�Y�G�\��wS`�ɇO��0�1}���l��!9 m��VՈ�<;���>� �EV3&u�S�nM�>��0ٜk���3�ܻ.=�����}O���{6�bF�"�Nޒ::M���a�$��iu�"kdh�LEn�d�A�7g�dt���a�W�=��e8H�I�B�����=/��/�M�q�/N}4�]��	�q��.N;��Cm��(��,��2�F#6�s^�4ti�� �|�t�Y,�"��U�i4��Y���t7T��4�"$�{�
��!���}m��L�p�$boD���M���=�+S�#�QiE�z���É�"�£PX�C��Ô2��V�a�y�i�/Z���9=�6p�p��s��К6Q,��Q�vÃ)��v��z���B#��+�e6�
B�i�s5<�(l�1g������w�Qx\��(�'d��(�o��]����i�f�z�O����E"<<�&�n�`�2o%�zX0zK�:��v9��ig #�{�$��SEY��f\5ʦG��@�/��N������!m�$P��  � ��@  5V��  m��6�Ij6�M��t�N��4�P��t��E��v��u��$�;R�m�/9ħT����b�tu��ncy�j\nԡ�<���^97 lg�yް�:7����ی�;;<v.�b뀻y,6�\�q����m���7"&:����x:��Of&�"٪,g����*յd��vЉ�:v�s�y�B 0��U��c�(��ͷ6�e�d��)E
m�'ä|p�5�,�~�΋�/l�Й>z�瑇�Fc2GGv	�gfH�f�.8�ѳ�0�5.��z�_{��Iᑄ�J(T��#m"4u0��M�F� ��v�,�*%���F���a�`i�Q�p�D'Db�GB~BhѲ�f�<�^s��������C)��)�ۏM�:yDo��
�6h�MAN,�ˋ���_��e`�:�Ee�!�諀��ȹD9r��,��D4Gy�	񶛜ä/Sj��*�m�|Q"���!�i"�&��x'������s��0���)v�,��V����H�C�?��>�"/A�00��$����7���G�yO��d��E���51MBD�oN1O,�_}�,�B �h���i��!�#��Y�N�wZ_+.9�Hj	طYB�l�m�][���tF�<)���&���JN dQ�Pm�y�3�E4�瑆AC���_��O�DY�$�a\�q#���O37K=�Nmdd�)'H��=6ylz���)���B�mAC�tXa�2+w�+Ș�f�Q]U�����{��:��5��f�G�n����W��i�J�1pe��OH(V��Zi�ω�{���ے���e�>�a��y��A�h:A�.4�_[�M�t����9
"�#0J��a������"�4�F��9hY򌝅�'���bU��cG)��[h���D�8G�EGuD��`�--D9�#[�g�'!I�$��3di�z����q�D�/H$&��Y��&g1�V�>Q;��!R'�9
QcF""���^o5��L��#�G�#��h1����BˎA^#�N.�g�ޥ��Q��`1�۩5FD�����}݉}Dv0c,�o
�={�8�;ԣ�B>f�c�}W �l�¬���2$�r!MΣ��M�ݐ������]n��rt�9��z�:�40��A0��%}j��&�������fY��M�^��Ht��i���l���2��4�|�)�����:Q��`���d}�滭IN$*B�rX���������kn��P$#�Z[W`���AM�Q�Lu��>�,�2Gt�	p�}�����2E��a,�hhxbC@��NK<�oW(����_7R�΂,�A�R�C!�x���ߨ]�P���o8:�n�k{��8��ы�b$-ov�9i����Ů�=����)2"�Tk�+a���C!��d4�u�zU���B=s��`Ћ�@ӂR�ڣG���v}�?Z���:��C��B���E���
�&l��,��g�A��8D�|�,��3���#NG�hѲ/���\4�NB�(�:B0�6p���Ey����Y��=�#2&bF�Q����.�8$Y�$�(�����O<�'�byD|3�Gd�0����B�-P�ڸy��>vQ�޺}��ΰr�/#�[�i0��v��y�Å����{��}�m뙮�����&��dOGv��Fla��E�"���HMCy�8|W�F�6Q��l�t�D8Etw�{E��	��%��Yr�$K���ќØY�8DM"$�����޳�
�B�����`A�*z&����\FI�h�zQ���y0F��rzh�3S
>[��H�DIÅ�4X�޸�F[�!Ivn���i�;TH�oU��z��w�
�R�!��"�'�i���
|q�[1�#��F�Y�4��+�t��D����jaE�\WM�H��2l�4GGr�p�dB!/hn���;�	�(z�sG�I�k�Y(��Z�zN�����鼢�v�C�������siG��������qZe2�p8�2D�a�0�>�[q"Ϩ�8D��V�;�A��
��Hs�<d��"���t����p��~�V�>!�����D�v��=���jKSE��@P�r���5ʗc��5��)�מ��p��s�l�nXg�.��8���|�#�I
7�O���Zaf��g[H�)�%;bo^���	��z�nt��.^u�w�sm�<��da��.%p���pW4�F�!R2߼�i��de!�DoF!>t�9�(�jv�Df?��#���}��X��`&��l�Z�e��E�_;5�Р-��2�mAC�\��ӤT0��ȟ"��Ljw�$5����0���a5'�)��f}D9�,��DZ�uV�(�F���O+�Z~��Zf�D���D�J�iuel�������<�y
��@�Xu�0�]��Pܲ���#���򈙊��A"a�dQ��C���E�F��#�P�<p�������0בF,�Y�xt��:whu�O!�z����\�(ᢱ�,-�����v\"6�or�C����f���s��XçԅfwgY	������6,4At����pcՉ�"�}�={���_���>|� �m�(   ��jZl ���   Cm�t�W��^4l�v�&��i]m�W�ۣsn�w��t��Gk״\���E�{�Ѹ{^���@�� k��T��l���;V���s���:%ЦDv	G�t���K�h����uv���m�-Y���N�;8�+�%8�K��Y��ݷh;κ�ip,\q�ņ�Z��C�v�+��nmg�\v҆wm�<�	�$j��bi����ą�$�(dr���1g�ޥ���kKH���l�}��+��b��Gda�"'�$1W �~����9�7�Vgȍ�S�YIC�yvD\���j(M��"�loK�=��*�8�J�;���L��0E�uĎ���������$aDQ�4�;o�y�l:YV�N�x4���԰|�b ъ�E�/�|�!�2��0�FQ�J��C���mv��a%�|�O4T��1��#ݯtV4:B��"����$�$1��DD�#L�4)�}f��q�)_,�7�G͌$� �KX�g�GczH�ި�axki�#�4Z��kչ5�϶َӄ1��44"�F7������0�>O[��0�6�0�2L��S��.��|�./e�"��(f�M����`�#
ϑ�gˎ�����9M��ܻ�-��v����y��om�u�D�ʒ�ji�.t��L��L�(�Yf{Iw봎2CkqEtuD��>c�J"���l�\�Ξ[C��/��'�z��.�4����y��^B!f}$gp�����0@�I�/�/k]8y���CJ��kp����K/�%����Q[�^/fʰ՘�b��a�����.�Һ�iv�s�g��ߪ]+�n�s�^�(�PȊ1��tSX���0)��{�Q$�De�Vb��Q��A3�3%8.7nJC6F"���+Es�1�M�q��W��/�������W�'fБG�
/A�.j�9������C#M����1��l�������2�����YA�z�lCO��lQ�[�q>�����DTttH��\�����D���w�nL(W�5h?��7��,' "(��_�׺$�Z]�v�`x�(�����iMcR��Jj(��?WY��ݺ�VĀM�l���K�ܓu��2�'0���k��m{t��/=&�vI�O7�y��0Ϛ�w�u=�6c�ֻ�Mok�;iE����C�D�#JɅ�$�%�ο�衄�6��C)l��Xj΅��>zM����l��:���Y���ʿ�gѨL&B��X[�� a�૛�w��h荒Q��D]L�J}B�^G��A��b*�[��^��f��0� 3Tټ�&�(�D���{�s;v��ó41P�0�}.�����U�8�ܵ�x\v+oQ�(�m��W�Jc��,����g5���u۽J��'�>���V-ʀ1�ml�A�����ל�`B�g�u*z���avG8q��WXy�W6RXђB�2i»y�Q�.�����mk�k-�u�^�:+�[�9Vp9��7��^�9ە���ykK��;��� ��@:����	Z���`V�`Ug�Br��,����f�e�ÎFkz6G8[�Mv���e�b)0v���h�g*&�8�v��vd�:WN������v��X����K���\o6��
Y���K���^Sy��%U�u��]��q�w��%j�8�SZ/	��jG}z��Z`���.��:�!�^eHo�6�i�f[��'}��])\���@��B\��ƭb���>��ͦ1rs�aE�ݹ]��������ɇ�SA�����Chv��Q	�͙�:��q^��=!�;�p�{����x�����5&H��ӕ��ҵ՚���[|okv�YYY[���]g[5�a���Wֳ���(��c��~bB��l�>}���={-��."�aHc,`\���ʋ�T���sF�4=�]\`Ń������R5^���{ڋc�i��}�\���� �e�����>>����A���3�tVoy�5���/#6֭b��63���.yb�]�$�#A��٤�����=Z��s�m��vl����J#��x�=�ت�i~��uxmnuJ#w�.��8��.�r�
�YKVe���(�����*����!7��$���;٬޻F_X�I�opSs�G�ܺ���!��G�3��X),���40����(S���t`<DE�
4h�$D�HE?w�W �]}�&b�u"����>.����=����)Y����1�CL����ϡY����J~;K�kD�y�t�<��*�pA���x��i�>��v�RUR�^�K�N� ���k@ײ#WXð�ze��+��\x����k���-���j?��nC�����ݥ�/�F�Y7�dx8/׼���|`�Nwx㗎v�c�s��U	9QZ�(����۫�u�4��
�t�i^�!�u��p��sNൡ�5H��pC!H1nKu7�qzƳ���Z ��y�1A�����H��5;�6��R��?hi�N�����yx��N]���xS�|q늽��xm�г<5y�R�_s�z�� 2�Y�4 �C9�ޏ�B!�w�J��+ӹ-^��!;ǎ���9?J��f`ʼ�
' �I���~kg�U�t�W1hK�؞w�;�z%��դ���E!�$EX�אVk	�X�קS줳�PZ��	�����=�5���D�M�����vpIGn�D�8
�T�=�dw׷�8o8���Ѷ�RY��g*^�z���j*J��J�M�o� �l[�icP l ;m�@d� �l  m���P h�,�cV��I�ν�Gn�'N.Y䫄�od#��\o�xC���e�1��8pXk��n0D&��Zv�9s�4/k\��q��5��=��T�P�`�x�;c��;vz��z�g��H>�@p�)�Λv	6�{u�yn#���t���}t���1+�u���3Ͷ@��A�0������&��AӃ�'<s�շ\j;qk��Y�K=Y7b�c�k��7�͔�>��kx{kt�jߟ�z.���ޕo<��,c�=��61~];'������E�5d	pD���x�Em{��g{�ޮN�݄����AM�co�}��r}w2�ȟj(��M@�0��L��)Ő�{�%9g�X���<ќ2���8��X�#(��j� ���6��i�����foy�@x�[1���3����bFT�6ܖ٭�b�i��*��^6��u�u�Z�ߚh�m����z��ћZ�x(U2�_���n�߽\�L��x!&�9kj��6v:��%�^�U�\�Az��[Ѣu����W��k�s��ڮP�vyr/�U���{��<�k�Y�/=�O<��������j��d�`��r��K�oo��x�Z�d3[�Z�;J�`N[gRN��8�eL���~�g��w]9��,���,`��T�
��pӬ��vAۖ�b�G�
�̤��{jOs�x<�����>=	���2��d'"�)���G�UUW{ے�Z�w�����z�`l��9)73�fg�!�ί���N6CFr9F����sU������ޜ=�D0�-�[��Vbػa����"q�m�;3P�q��JEh��F������/��������V��mt�fP{�sp��W�&�mK�S_r r6ܐI��x�r��"4=Vn2��{
u�1ۭO*�nV�<���D#q �.$���~ћ��a��J�����7�]8�7P"׏C��R���'8�B7i$��-��R4�xK�xq��>��^���)3�^���D�"%��]�>
�ٗ��h��[R�
H�QA}Q�jo~��d�߾���n.��]�.�1y�� Iճ��s_Qܻ*�_A=W@��j�On���u�2+�=KiA�� s�mYS2��W��e������*C�4�ݫ�~wI�M�oȞ+���-���Z��]j�՘:�������r��`��&� �&CN�z�Ԃ�k~��G�V�S�s^�w>Ոyx��OxG�ʵн/ϳ0��	9F�Iٶ���A�a�<���Gg�qK�p��u�=\(WD���Tf�W;\�W%O�.Z���2�i�����)����7neoل/�$hG8Y�<(�/�߮nﾙ�2�2B׉�o0���gmJh6$\�0b��X�O��_��e�� �'`��|<b���z�׸{9쨟yaZ�%"�q�����8����I�P6,�&PR���+�o���v�t����>�!u��u����K]��x�R0ئw��0�H�0�s�:�����m^#����yv��$[���2��.C�{���t�؀R��V��bX�豽�#LAA6��k��/�Y�!��z�{��;]���b�<[��F%�Ÿa���?]�-���)��3jҝ���ܛn�()��Zkg�8.61[�g������Y�;	��h����!�e�q{�Kj|;+��N��Ǹ׺�P��ɬ>��8Mi��Y���C}�}��{��U��A�}����m%�. .Xh��f�m`�[@��m�yo,+7��2V�jk��,8���j�=wv$��S���t*�D3}�,`P�8N` My�p����u��F��!T����h����Q�3�㴮��ޖ�/Us��=T�`��5%����㱗�%�Գ�O5W'>���hx����J��{����J2�;����^"�^o7�8NfX��!ՙY@e�i'.�_}��m �Z�-]�CxN�їКؽ8�v�r�<���`	�[R    m���m��  [A�`   ր��dN�͸!�&94ź�v�&�*j���kuy�M���6���=������� M@L��൶��.3����q����9�=����`��t���SR�EäG:Io�m���,�9�4�mD�������xzzz�Y�����r!ɹ�/N�x�3YxnU��y{Q��έAjT��qa:[p�l���n^/`|k�,��D� e�$��m��9��Vİ{�si9�u#A�Vg.�^WB3���3د>�W����"(\,.$Ǜ�}���u���<��vY"fҎܥgWa��9�I�ⷷgvU��ˏN��S�Zm �6�FA[�h]���<�m?��~�o��*�C����'W�F
�ܵ�ףw4jN��#���)N6�T�#u�t>iX�7�+Nś��J���k�o_�l���3t<sK�QC4]�>�MX�r��S~	jN�e��<5�ιN�:��:P�R��N�+��u�}�|�I�!e�m�R���d�mcY�T;B�ݏg��N/8uֻv�����s�H���2G"m�&��]���^�����83��g�6��9�f���l�׏5?�)�������2�mIQ$�w7f�R��z�k^�>��y�q̸��v�d����7��.ْ��t��wZ[;E���f�gL�ԏ���C�g&H˰�1�t&��b�X2Kp���+�چ��bJ&ȒZr7#�����?���4(���>��U�:�ɓ�t�~�ݙ�qԞZ{��;t�3:���I���� �3t/J�X��q�!x�2����i=�;�R�9��tc"��h�;�$����?;޻�D���	Pb'%�ڈ���딷e�c=�k�Y���:���Ϛ#��������#���_���^_�O:K��Y���,MS��NxF�%:M�㥹��ݷ�֯0\�:뷟	��{ ��xWsyD��|��� �չ�ej���#�qk��f�礩�7겝��Q#C������_>����fVl����á����6�����ɻ�����}����ǻ\6�6�h�D���|Y. =����:��]:���&VUG�>UWGR�4�
ʆ��܎��ܥoE-I�A@��[[�����\������ʃ�~����Qw���0�9$�챒�O��u�n�kz���/cO�#pc�{\�F��siH�P����s��2��"��i���mn%�������N�tul��qw_�ײu���@��,y��כ�n��l$-�ɬ��dm�iz\v�m�lZ8�v�Rix���M �nڰ82�;˄�.z��_qS��[ӫ0:=�J�o卟��w=G�S�f>l���1P�)�>��;�U�.[�g6�f_��WN�ܿ/W��V,>~��v�?l���v��p���=G�Hb ��f`�����xmk�/Z}G�Z=[*|� M�x�{_DZFM��^�k(���a ����������Lo7�߁��z��K����8�GH:�t����͜} .��%X�s��o;�V:�fuf.=n���S&��/��͖K�:���h�*��ubg�^�1�bj؂8�"H-�d���̓�mZ#�z����e\�hu��==ّ{��1��r�ű����MM$]��"��JJ�j�v3�������Ȝa���n5���1GvLDiD���-�܇���k�^��W0ڷ��b/&�F�������gӻ������ȓ&�q�i�0[�z�t�Jڧ�u�}v&w��[�"^��͏�^>G���q�ײL����r�`�G�^��P;ѥ��q}�)��鳇��ƑG���ܺ�~[[�mA�>���>H'r6�΋�د��%���\r��?#�q/-�z/�q��Q^�2�+�/�Y�����J�o{H��	&��3��&���ٯ�d��cA�q:҆�P6c�-w̡�푶gq�Ӕ�RuU=�����V��w�ǈHX89=�"�Λ�Zxi#��n�y��=�=lZ�O����J}�֮w!X]`X듵�3�Y��__����ٔ5�)����E���V+*�#%�9��f<��6�]-8ST!��Z�;0l��>�6Ջ�/�6���f�G����q��/A��B��0�ȅY2/�C�U�W�F�l�+aA��NVI����ZBû���7.��uЋ5tdu��ٳ%���eϏs��
���� ��<��!5���8�S��,�z>*� b��7C_f�3�4/Y�:���̆�W!�1e^uɢC�{3Y�;8�=���e=��3���GR��qLev���aނR������v��piz�D�Y���8GL�������0��Z@��b�$�l�wh.Ã%�1�譾e	Tz��͔��j,�r2!L��x�	ޚsJ��ڙ;�]��
�{O�<#Zl`g.�ە4�-���J���r�]>��,�����n��!׫M��L9tw�u2֕�ѵ�;f+ogTcޭ��nf��0�b�3&��%��2i,��5Vv֚�ټDіpdk�h��C��|��8e����+�[ժ���"ɤ�H I$     �l-��   H   n�݀ҵ�`հ         �        �` ^�I���    :@���m�          �e��v�޽ڶ                    [Cl��f��    �  � �ft��w�M�XF�9��ݺ�F8�䮼vi�'h����u˦^��ѝ��=g���$����-��L�4�Rp���'j�W�]N�#{kG/���#����w=n�Z{*�釱�[�����uj�[��	����vN�!�����יLfJ�Ką����3����m��k�֧v9t.8����Y�ӽ�����:��9	t�CN�����	��s�a*���u���y�{�n�x��ً�v9-�䵌�����;pfqe{�M�Ğv;osõc=�ێ�d���=�3�]�ORvw(�γ/���YT���`�%ѷ�ƚؗ+��I3J�D%���y;ly�Hr��s[L�NT}e#�����|�6絊��uH�L��O[�����.�ݱ���&�ȼ����J���-���Q��֬O�c���vѶq@�7���W]ڍ�g�s��1��x<�>�.�X`ݰN��)�;������m�x��c��.�;N��'0��n{W��s�v8�h�v��ok$��%v;ji��^83s]���㭣��&jϳ����Z��7Y��Av5��m��9^���-�n+]Y"=^�6�1w0�8�������u�:ٴ��m']���(%n�����u�/^��<�j4m=[P/ћ9\�k���q��q케�v��=���q�=A1����j��f˞ 8�ۛk��}�|)<prq���[Bv;�n8��7�Ǎ�NSzĽ=��<��vüp�;�]&ϞŲH�:�Q�;t����k�ln�]V��ցm��@   m���� #lۛ`   sZ�m$�$��K�[O!vђ�(qp�+:7\=.u��+�5�Ș�ú����W9h卉�pl�։��Ʈ�ܹI�	�𽌖W\�vѡ�M��$8`�n-�(�mI�o8ζ�vța�'u;�1ղ��ޕg�'IN�G�޸8�uO<'4>!�rBy�̗K��� �)BL��˭uj���F�K1�q��u���Y���n(ܩH@��4���յ������mu�������Vy��u�L����A��x�ͽU�@�`R4̐2�pdݭ��'���4ƍ�[�~<��Vd v�>��zTۃ�?�t"jw��|2���"�a�$��%p�m����W�G�MF�U+sA��!�)[3���1�h�[���d8Sa�#��$;�����Ư�
V����3��S�%]^R�������Y��^�!W�����5�	'Ri�[�X����٢`��i63r����^��k�"�Am���EJ�Vbm�6�HN��]��nv�������L=�x���7m��Н���MÄ�jW<��\+�S�:k����׼��=���i�Ո<_�sj>��2����(��E��y�cb���׹O�IG�����nQt`Օ�N���X(���\6�h�=��lVS�+u�2pok�g}���Wz3��7S":]��{�Wwn�QVz���E�����>*퓐*8h�$�ss�J�3�Vm1�E{��jV���K�E�f�/���
����hVU�`f`����7W:l��k�<���S�m8������;C�$j�j̗�+Y#����!���2�w��!�Q����҅���L2�Z�z�#���EA�����d�o٣�3{� b�Ue
���.p�%�.%b�K�6���i{�`��H��)t����stC�D�h���Ţ_��>>9���R�7���хt�k��z���<�da�P��[KSl2
���nC�!��쯦��zH�Y-�Y���U~��xR���g�Ϳy���l
c#.�S�l��$�A��q7�%'+��c�u�𵸈]�	uO%���R�;���{G��	���P�v�q�vc�׷z6'	n�4�ס��}���/�2��@�]�Jۼ5�y�׎�.`�R�Ɠ�zf�.�h� �ַ5�{3��>���T�-�x�oMܰ�հ�r��2X�#;�KX���u���q%d1'r7#�*Ե��өK�Ȋ������_'%�j��m�un�e9h�E���VnRc:�.`cm�_r%r�f��ʊ�u[X3d���;�,(1ƛ��H�dͦ6�k�},����M\o�]t�5,��n����f��f�-��$>�,�(���4�>�E��Ҷ�R�~P��UGfT�tq�����5�<zq�)�[���>D&L
Fؒ[N�^]8��ݰ��:y�٫��蝆������.���f�ڀ��-��l�Q�$	�ѥ��[�����Ri�V�����$���(c�!-��9r^C��p[�����Ը�4_ ��<�GBƎ�7��&/Ȥ�=Q\���ń.�{�N(���M��V��`�B�a7tI7���]��x�m����}�I�/�O�<�-#6ݮ#lf�t֍�T�1���m��/P�i���Hӯ*�E�N�;1vS���<u�Ǝ�c�P���n�ܛ�/e��I��^�i�������xs4|���q��W�s�~�^0D��b#�|�)�D6�
�
�Ƣ���z6�������s}��M��P9R��O�|�h��h��v�_q��_(�,,�ab�x*�%Pk�yy��n������~R�Yِ�����]?=�M����W��Mͤ6�/��uD"��*��	w>v^W��0v�8W7o[޿bꕣu$s�1'���2�,3���k�<p�ch��M�)&;/����?��� sh�ӛ���Zr�R>.[�����{�_[(�.*�~��ۥX�����n�gע��ᑥw%t��ٌk.Ry��Ob�́��8����1�XR������$t���� �P �dր � 6ګq���@k�h�t�^{��CK����8=X�Y�;�{r�V�۲�z��S�����ԇ#���wl)���N*û7O=nm�!�kͻsc�/���=��y��b�q�t��HƺrqVr�6W:8N:m�;G������p=���D]�{RNV�V�v�˻"�g[z��v�L5AC�eZڶ��oF{xi�ݺ�kl�<Kf���vy����T�.݅NŮM ��_��OZ�_�a����������>��09ti�a� 7���mj�6�Ug���QM� �F6r�x*Wݯ��yᵢ�����ho�"���d��3޾M��ǆ1ڊ0�{�%w��i|�a� p�0ok��c0����Mj�O��IKp_�:�V%.��'SISSP�,d����γO�	&q��i�.�{UB�`�O8ﳶ��/J#��5bhT������Pix>�>�~�z�m?_��3v@9d�X&�]p�}^J�f��κ�Yb�׳��g�%ue/"�LI���mk�e�G�h��^V�A6`'Um[��l-��ˁݮ��c�m`�s���d�
�מ���;M1m͞6�Va����sw�O^�z����1����A��²=8�fW\]^N�֝Ծ>�,����38�' '\��yxʊ�{D�j���ЫI���=H��wx�ݮJ��D�чMћ/���%�Jc�_uy\R��D�n�>��&j�Qgj�z+�Р�b==��C���D6�B�rY/(��^ݶv̿W��X��^%�{�=�M�o�e3�r�`�vk	 &��`5Ǣ���כ�����W���:�����U�Ƥ��i�Bzg{)�_V�/��F���l9Q$	��y
�To<�ǵ^���K> }d�Lx.�a��5�;�R��o�u�L|ZE����d��];N��m�T��Q݈��eͺׇ#�n6�W�S���gsayћ�Mo�y���	�؎{�R�o�eOR[J�47��[��K��MA�YH|l%�I>����ko
��Y���o��nxoL��ͨ�j��x�-e)S3㹎���SY��I����`�w"�����j�������u�%2b�
���)�_v��=�`#LU`���]�d�ҳ����);�r�ݴ'A�A���jb]|�=֑�b�tb��� �Ju,Η��tJg�~�yi��|p8*bW�}�7%�vz}c�eIBw�c���3�D�E���I�};������>~ͺWYo<)st�g./�0����zz�V����"z�`���[*�ջm�Kn]�8t���n�1&��s����<].��]�ni��%6g�V�>w����+��y:;zsR��׆o��r���ӹ]yd7���:Aײ��&�F9iT��,�:�v��y��|݌�v�ǃ��h�2�p�v��;�X��,�և�&D��Sf��å6!@4@��Mj"����q`�|#w��l$1h-9ge�2b_v`�Jb���n4�6�I�7!����{ϟ�K��q���Z��W��J �ҵ�e�%���Wp���S+���ܼ2{6�,�Л�DѱӖv[8��c2b�2���4M�����qD�}�4�m�H�I�)ա��`ν�m�K���_x��f�!=n�_�ra�{T0�]�ٹ��t���B�Nӄ��)�ۢ^�K�ʔ�Nyc�گG*��
�7;^ϵ߲���Nq5q� ���}X1n@x��-Z5����Vl[��k=�����m �M��IH�!B-F��vsD�3�״��g�<�;�ִ�iy��N��ұ\]:Y���k�[PP��Xm�Ď \mɳ5�F����-�vPƣ*U��X�ܷdї
*�]:�"t���^��"��!�
��������'��m�U�>f�q�*Ž��[��ɭf���:�{�{F�4zq���L�S��c��^N����&U^U���r�K�����Q��O��TZ��i�0�S�]��O�����k&1,��:ۜć��fm���}f�bm��$��\bp��x�Ҧ�JT6E�T����z���ϯ� 	h��k6̀  �/C��K�� 2��   /Z .��5^�%��t���zF�7%�ӵ5�/��:�`�@�v�&t�]u����SW`]�Xݰ%ݮ7�6��`�+0���r��vvx��g73�6�7e�ֱ��,�6:R[]Oe�뮣b��z��������Np�.�c�D�U؅(�0Y����V�ul�6�s�7�Ѯ/n�4s�{N��\��������v"d���bR��18A87Eכ�]��ٹ)W��V��C=�Ǵ��5�z*l��/o(IZ+�?��!"9��o&����1�]ӗsZ��#L���6��>ЊR�v�f�6�އ�XK��XK��h�	NG�w�n��W�B���c[M(����@�K��3Ms���wP}��ؒ,�����������^��I|��1G�Z�%�k�PK[.VQՂ5.�5�6	G��ݟ��SO"<=={�j�	{2��ɀ�s�x�7"5�=^;Gw.����\��W�ɢ�m�[NBd�K��V����vɣek���9���a^���1��i��P��2I6�$�������Y�_����FM�H��Ӷ��xyT�OZ��[&	�� ^	6	�0����{��vȯR���BA�-���y�nU^��9V��(�]�hC`T,��W�wA���i���GPN$m+�ӎ����p�K���pG"^��[��A߹lZ�su�!Ơ�5Ĥ�g�o��&-�O[����.�����ˤ��{t��h�Տj���)��$&&p�_T_�L��;�&���G�K�}��[W+`!5S��NӫD{�e��Ҿ6g��kZm���I�sv�AF�'b�7'di�`����Z�oZmX�� �����帞U׽pie�dM��U�jgƇ&K]]]���9n+��n��zݞݫU��;Z�@�&_b�S���Q������ַ��B�Y�~��U��Y���?n�p��˚/jOg�fX6��bn2����g�����ՑJ����{%yT�gxD�3���Jط��~�7�.�������]���N(DA��$����
�珷׽��q���}��ɕ��꿼++�)��#���zbϕk:Z�ʧ��E#��MY0�,��o��3)�%S�2�i��,�9��"����Fg��]D�e;���*b\sY��t�J�ɝYZWAXbэ�Ef9ӥ^�a�htI[�t�t2
BY��H�K�x21�d��Ŷ�İ����ɀ�0�\Eͱ{�`Ćn�}���S����u���\6wj,x�*D������ڶ�����77wy��=��[�F�p1����]���A'Q�݀���v���f��g+�dk�C�W�ޠ�N�3�Ru_t�(m�����2�(�,���)=bP2鈒�����WUv�	IH��M��q�Gy�zw{xzp�[w`��)!��FųP�˜��]�Agp�F�M��M��g����X�$��:�]��M���T�c��n�Lһ;����7nn�\��r`|�s8�u�c�����]|��iZԍ^s`殟���ݖ���0���ُ5�LAU��)�(��u8�Y�jEI��
�Lu �;�5^d��T��}�������b�mn��rM�-�:gƗf� u��yS�4l̓�����P�����]���n�6�\}ľe��aȡ-(���^ݹ�`�:������{��nӈ݌�C�f[�\�{��ᣱ���Ԫ� ���!���_��i�bh��1'%�hnt�Gu^�9�V�N��	��
k�����e�nOZ��7���}&-�^��D6�_���kj(�U�qܭ`ݣ��'9�X$9�v��::8�ȝq��/l"�z`�3�q���;-�B����Ov�Ѵ�Uu����Ǟu��"{9�^wV��yWt=��R6���$.�n��ۤ7՛ͮ�a�2����F������=8�=X�������z�k�Q�&�כ��B8s�E2$@Ln��o�9�{���X��j8���ڛ�e#+Ck��}�q�]��ї�A-%&qH�ڼ������mi[�f�]�TF��G]�Įx2�gb~�4��x~ܐ��1OM}l������Ǻ\�\Zn�QI_#-�γ�N'fѽ|�N�w���B��>3+��i��2������=�߷2�&�d��r)2�\�;�ӑ�v�Oy����]�\-�X��f沆�y�Ig؀�ʵmP���:��eu�v�kqu�ه���8�1�ynn���a�W7V�5�����#��3��Etl{{#[v�Ҹ��&0��g�ԲX2A��n�����f0�
B�Ilv�F��{����Ai�e{I|�5�r)Tra�[�t897bg:;�Z�ƋɊ�q/�*��i�i�N̜�I�B�
�~���ܽ�Q���ta�l?j�_Cm����z��=�v�ٷW��M��r%#u����?�$4^9~����ù�
�JS��1qh�%�I���޴=N��y����tρ)��$&&r�tQ���yJ�Q��#��5��8uU"��;�v:C(����|��ˋe{F{C�]eJLf��ZU����pR�v�3-�2�XN���ja�q��b5���omuW�	ǹu�@��RxI$��vI  /[��  m�*m� �l��    ��޼��"�&q�v��/7���n͎y����@��H�m���E��	���<8MrF6⎇a �X湝�N�e6�7]����3e���:�=v�ӎ�~���p�g���MۖzȨÍmZLiӌܤ<�M
��0����=�Pq��U�s�������-���;[��5���*�j^�-:�cVz�n����6w<vu.��]���K!ƣm0�	I7�~�����fDܲs�xk/�S=w�`>��_=g�o_��u�~�0�I�5%I�նPѽ�U��w��;!6pR��vU����1�J�L�ݞ��h�G�3�OZ[y�+�]���(SB���<{����:�`��)��}��� �f`�L�Iǎp�_g���S���4[���y�Chxx�쑶�A�<2Zzo8O�Pӽ=�y6����.�c{hp��7Ũw|'�6n߬_'ڼ�e4�r(ZF8���=5?s��,�;�2.K�w!oCI��8��0�[n�U>eOݡ���m�X�������,@�dR�V�3�}����]�q�zh�]�tn��F�f�v�Ȉ�. �3�f��f��H���TPJ�p�B<3 ��aq}���^�G�b��n�[o�Y_y����Y�fyZ0'lD�E�\*pUS�����U����dP�\�s,@�澭�fE���+�m�vvR�N�ݙd���ݾ�fu(��I(�l������Q}�Js�9}w��%�I��Úa
l-��%w��h�p���A�;�Z�]���{���@��� �����/%L�=�z���}o�?wI��D�wvU��
~mB�.#������֩>ݽ�U��S*N"6;�Mx����r3�l���qU���;���A���"A!.){w���2'OV#G�۬�����Q��i�u����p�f�tZ]c֝�C�My�?m���?�Uڇ-mP��y�v�:}���m���v��8�#(c�m�Y<�91u�����"!�i��<9�Y��݋�S��[V�͜k��y�ybĆa���t�V����uAv��ƧL6�����1�2�w!�]���o0}�)��%�)�y�ӆ�a���hٱ� L*�"����=�_o{�O���p8
p��RG�!TY鷟3*�w�V���9��:�W��Oz��#5މi�p=�a�̓�w���У�ED�ƞ&#4u�u��*�0f�^b(�+$(/����O���tV��*wd�,��P�\e&$q��"m�۪���+ř��4�f(�i�Ղ�=�^��?�ۛ2��%�`"�ܷ7{�h��P�lؒm�[q��%:w�P�MP��p�v�}�K������WLmGD�]�̫���G��&۶}��$���T����5��l[T�չ��(ݗ��a���f��p�WW��G&n;;6��Hx����Fz�y�6m��f��y̱c)�pub5zq�5�����{��yC�y���������`������,gs�,���̋C`[dbÛ���Z���Th��x^�2�vGs�m)īQ8�l�~�g �>�e�$.�7�~��z����]ѱIe���|u�;z���>�(�Mv�n���mmA<��IP�Z��ڒ|eU��4� �q�ya5S�Q�i�l�J���g�7]�ޔ���-D�k�M��])�X��a\;����qa�ˢ�r���iKvĳӎm嫡W�O~�V�QP�ye53��_?Z�w_|t�jI�8~G(aw�]��~��:��6���.F���m.�5�@l�-���v-���.�1<�c�̫��2��Qo�+Z���B����k�	��`�n��5�I�#(q�����Ksj�8yŭ8�0���R�����O������Bt�d�t5ô�D7�E�3��Ui����=�Ar�C
�n��v��oJ�qa[�ɘ:�H=RW�y�̄� ʪ���w=3�}�l߇�����/,#q$(�[�=}�z� �^��U����!++mS�:}�[�71��eݝ;�Û��ߟ'��H�nTF8�!�P�9�PLD.nu	�z�kN�GS��1[_�E(���!��b6F��f\�����˱b|5�H�,8�d��U:�&WuFe&X`��X�ˮ��ŕ��-n5���z۝�M��ǭZ#��`�}�P7�L��#���Q�M���n�=-��j��yMټ��"R=� ��N�q{���h�f���$�I7e�6ؑM3   k�-�� 5���   6�6�m\��m����0���%��j���y܎�68]2au����B59RQ Ŏ{me�T��Gi��Vy���r\���;m�����m��n�8�l*���"B���\����^$�Z�n{E��`ptc�����ӷb�:��\�a��i��Ge������wӸ�Z8�5)�����8E�ku�NLv�x�\%�N{{��@sB5��z]�����l�������?8�� �WW1m\�3���7Zq�i"� Q�յ��jg��Őt�_��@�Rq�\�M:<tgr��	=z`ӆ0�$��+�+V�;p�N�����ç�iڥ�z D�/���R�����čGȜ�5��`V���=����]�\���<�t�[���вAds+�7����,�{�߾~�1@��Q�����������;d%���U����{)27�o�Oo[ТRQ�A+,F���_w���J�f�#e@�p��rnҺL�s��J����Ռ�0��Ӷ�5��5s]���4�WT�|���씱��3��>��93)`Q�!l'	m�'Wn��qXG���\�K>4%�<��[�ͮb�Usrr��i�[q��$'<���Po�g��Yݮ���{v�ү�S��va�*2�Hޞ��.�i$-K�ۈ��p���Y�P3qA�=�w��g���߸^c���̽���α��rP�i�hN�n0"8d����]��gi�Գ��b��)�[�H�J��a��,9�޶T����ӈ��l[��=O3�Z'Ƙ<������Ɇ�$@�"������6ٺ"���ڳ���m0�ۺ��n{��}=3<�d���稷�(4Ђ2�����b�hm��"G=��7)]��2k�2�2���b��WXsY���I�U/�:L���{�H�0ـ��rx��g�\^�k9Rf]�a�3α�5u�+v�EK�w����e����6���7a6t�g$`��o�H[rB�p��jף[��I���:��eI����v&�CK��^�u�r����t�F����������T�PR�⪃��'�u��"��}�>K����(d36��~�+�Bi�8�X��+
�����XQ��o�wc(tf��Q��T��<NS�Rm�Ô�<r��6�=�P����"d�C�B�����z��p¬����v���h���ð��ſ�A:ێ��zo��7�����l��rQ�R{y�y�6��t��$�g�|s{7�=�/��n�qw�ߑe��$�[�sg��������S1U�7}Q�܅�	[�T�w�"�&e���'���(����7��n.��>�v)
e�
��e��jn�>w������ƫ�mս�zv�E�OOi�u(X��V#�%C�S�N�c4�8���)������;Jd��[V݊�.��h7.u,.�3U�����ڸc]��2ɹf@K��g������ykm/}�F�1b�J	��vn;l7o����k��{{K�b�>M
��.)��ɯ	�#������ɱ�t2���̧��t�R�jn�c�%}AczL޼�L,nv��M�Ò9��zu.�����Wj�=��Ʀ�-����:�ʵ���ݿk��xӺ:o
<�r�n�G6�aܻ�7 �8�t����]� C�>>ɟ;0��Q�=��_���q�+)TȬދ_,�h/�����]���w!��vv�4��8�ӕ���sZ�E�!/6eq\hZOy,�[��?xf륻�{_�BFb�8�eG"�[{�1�y���Z������H҅�SPZ{�2O:V��׃��ܝ�����6���j9nIV�&����JaR�W$�ln�����9�NE ��"�t+�k�߿��;*�{X���h�ݐ��-9�㞷�[L���+Z�y�,�NEk�wgi'J"Q����޼����=�|��@����Z7�{~�B�&����mS�GS3�����~�k3;0 �����u�������c���,݋�Fcv��-��&cT��w��n�1c��=mu0� ���[���y٤/Y�b�`�����޼�p�	��i��QU��n�<ʻw)����AMEL�'Sbtu��&�L3Q2��2�=s�ozq`i�
���&ޞ<�2d6�o!@RV��zw�����P�����ȷ�M�!d�Ν��ME2�\��<ù��lf-����[�=��aS��{��s`�%�KP�:��b����*sC�tns&j�x�,TwR*`�q"�fg	��ٳ�*(^��kFBk{���m�т�e#�x��Tvk;�weA�m���tn�$[μ��d.oWOP�.����E��a�g�$f�|���nnj̽:���-Y�ԭH�J���r��qVݻ?j ��2n�4�N1��*P&Xd�2���l�U��[\���}�L3+;6z�'%.³#�����m�ް-���2�L���֒z���Mn�w���vu�V ����«��C�q9S��[u��S	fiAh뱈[��/DɹM����u�#��LI�*��VU��n����c�+��@w�uʹSNh�#���N�T�)�b��>�RG0����w|�O]�����$�ͺVmG��kE�x�w �:H�xՊ�7���-����b��Ggo�t'�!B�]�&_w�w�&%y��ǂ[���bGP�C�3�w0m�f��z{�#�v<H�S��쉸����n��8�IU�b��{I�:GM���J��=^�,�sk�|���߿ m�      ���   ְ  � 	�����l   m�   �        �� k:�6    Ďh�6�   m���y      ʖie٩Vݩ�[(�UU  �         �    h ]��� !�     �T��W�4���9���,\umb�͞n�v��w;����vnG�c�u�-i�v����r�g�9�#�������q��A�{Vi	��/����lb˃�c�׶
�d�-�]���τ����Y�s�\���J%���W=s�[ol�sh`�����i{��Z-/h:h9Q�f2+=�=:.ݢ_]��^N���p��foq�ט��s�d�ni筟[<��鬐��I�����pS���Pnn;p�i��N��e��1����N����7Q��q����ݶ�ax5�b��g�]�n�*���O=P�&���������:��nw)�����h��]m�f�������gm-��Rr��\���@8�cۧ�;�A�qɳ*�Z���fP�ύ�>�5�E=���s��gg�g�2�ڞ�6��˶��b1�lPlkq����� �����bq�p&u�4���n6�z�����ϥ�;=�A�Em�kl�����%�X��β�k����a�:m>L�^��v��V��y&k��;l�ݪ���<nÍ�6��w]s��6��E�Zv�,v:<��k�طu=@^s�݃���a^�.�荩<ö��ñ'<v�v7l�[[��r�''/]�5���*Z�	����ݟ`��z�^��G`��ɞ��(�ֵl��qp�7�.̊;�t�:1�.ά"k�xy��h3�5�5v� :�O��}�}k�'nd�{==�@���{]�"����5�l�؞l��Om�]�X�5�ᔷn�@s���r���Ws�nB�A�t����y��[�97�;1�����`#��$V�  m� β� u�l   UUq�b�mǘ�upEt�	8��۞s$k]�sƊ�mwi���O6fװ]ob8p&y����[+��f�;T�]�c���D���7O6}e6~��2s�����oT�a;��ƌrr�۬9|-i�4�l/J03힎�c�sڕ���u�]��Mƹه����%gsь�VV�SYF�V1�+n+��gk��m{s�ٞ�х�l��\�.����솘l�dm�?�-��ݾ~�zΗ�cuQn9���m2��4DF��2m�\�7S����-:0Ƨ�w�e��DDz �g/���)$��9���0S��/�QjG_�R�ɬg[�M��I���Zr/��^X1FW���3���M[�rHY��+�<�{m��ڼm�Zii���X���QPZy�F���3���VB�}���b���1�
r_ݬ{�5��3�VU�b)�����x�d�^eD��jV����p��m:��:������E�FFS1"�.t�{D��L�>eQ̚-2�0�N���[X�U1�љ3)߷��Aluv�Mx�}g����l?�S$ڳ��U���u���I�-͛�-��[�S��w>l�β��1�዗xs�|�=?]}�ʛ����|νͶ�ў5���g�El]�~�nC��zP���Z�W��I%�!J@K��o�}�љӡ����Q%�m�6d[S�����{֨v�tY|�yj��.ՏOt�K�iMCOeh��Y�:׎]�M�~���S����g\fT���ג�����f���m}�\)���&�I�h�ʪ�8z�zb*��ʫ�d����\�k������L���iZ��5=s0^��g�`�^b)�Xr)4���ם�6\u�2�5��d[Ԕ�\{�{�R����So?��<�􂙼5sQ�Ҷz��z����8���-�ʑ�Ż���/c{��wH��Tze��>�uB������.��]׮cH�̀�������W��n�Q�!� m�'R���m�U���^h)�D�ۺ���o:���0ԑ��bF�l�����}~��*�{β�����=%e�˯T�=�.7N�9��c ���7)6�ҙt��۝4a0�",��}�`��r�Ck��+�w��NϜU<��'N`*�Ǫm��i�-�����y�5��5���V�H�����m�Tfp�B����vL�>~���֒٭��S��W8L	�yz�[-�����r�B�2���1v�-u{e-l�^*�b����&���PD�Ơ�1�d�u�2�{sy�������ɸ����{�xb>��� ��I�̾ YL!�Ω�}������U�St=��̙
�ף��{����q���{o�|7T����հ��!���p^��ת���̩��-�]8��qus��c���UQgz��t�BR�Q�󝻚��{�|�=;���׵�ٿ�	 KL*���6{bC�e�6����,-�\���h����r&\���c>�c��ޝy�+��%�̺}�d̪c)S�F�S��iζ0J�/jRl0�N6��T2E�V��s|^�4��(�'�i�%pӽ6��e�U�,:1Y��e��G*�V��;�$�ڑ�M����������g��y�zם};��c޿g<��A�d�׬�6�K���zB��B�w�� �8[�;�M�#���^�=�:�����#��+�������i&�g$/2���˖�eJ^!I3�4�Y4Z��
!�1�y��
B�i2%��c�l��I�0�sB��v|�j ��F
I�aNL�l�h8��oOqu��WBu�a�t��=#��U?\w:AR���wI5��tF1�Qta�\��%�E���ֽzT�t^+u� ���=u��v[uÎ'�s������%��c�4�2�̵�攏��w��y	��;F2~���3'a��ĝ�Zʭ�'��F�O��7v�W�Z�!�	�B��� ����9t�c�|�Lʎ�x��~�L�Ln��~���+D���*�VC�60��;�z�CyZ<�	�Rcpgw��f��~_���� ��F��޶�~�Y IT�7v��1���Jkj#��6�o���T=K��6�"6"2���x�{`;l��L���5��̞�^d�s8�P3.��o�mU���(��O5�Ӻ�*p���e>�FH�rG>?t�;��`�����8K�:�����#�M羽�T�O��9�g%�h��k"(�5�EM��v��o���%Jƀ�K����Ŋ�G���\�Yz��;}9��*荺��5�/9��,a�p �BD�����   m�Ұ!� n��   � �yۯ4�k�̽z�<K���]�=� ��<>S\�2֢�@��F��tv��vn3�g�Y�A�(����%���{+؛h�y���:S�l�5۞+`�]���Ëg����}�\�WAgE���u��b1�6.�gX�yꔵ�qZI�kfΥstk���d�ꌽ.�H���2�[V�/]m�w\F�8-up��7�g�܇�8��Ĉ���W�n��(m���|�b]p��u@qs�,���J�-�<�xk��Z�x�'�mɧ7��s�u�zy.���,E�$Tr.���bE��7�ꄣB�viy8�`�Ѳ:����\Z�h��.��b�g�1#.A-�6!w�f+ޚ`���h��Q6��IX�O�w��E+)Ud�Zs�4���{5ζtDQ���n:|�����%i��|3Λ	��Q��FN������n8d����E�6�K��9�:7O��W<�JJ�!y�^z��GK__��(��o/���	2�FFT(#=�7^����'�c:�c�3����;�����K(8��!&�Vv2��mґqw �(e�p��z�˾�<��lHM6m�Pz��������$.n=����֖<s�A��ՔM�N�,�]�^�����F������/���{�c���'�ә���`��?_h��ϛ�_N�Dv���8����H�^"�j�ҳ#k��W�"x�n����K����Q���l��YXF*�.�x\}y�)MB�`�;��tj�᛺�|	�9�fT:��1ş��c����F4��iB +����;���eK)W��x~�P����	M�RF܃����.��oZr�
][7S��Il�E���+s���Ed�<�޷D
�㕍i[8��^/+֒I"
ّ�Nm���q|��k:�{j�h��fDVQ��F¾G^De��c��r"t�t�罄V�CQ@L���}��ju��ηo�#��IrVGG�{��;觟y>��{3gy�d�H�Q�w���g��!��HFx�����%n\s��j�{v6.�͸8�e�d���*�{ �������梅Tn������2����f
�����\�������^1\a��}�I���"Ä$���>ݾ���+-�斎�w�CVf�Eu����ֹ�1�:c��Af)��^nx*����I���m8
n�e��^����_�xV���g�1?7Ku�/�-m��X^2�4,\[$�_��QP����]զȽ!^�Y�.�T�G2�p������ҕA��VB�oK،�+�h۽c�{:�w�ɍ"�vt�X��_�P��P �5ը��w�<�Z�gBں��U<��oϚ������6�۔�>��f�OI)5�E�����lw=�vrb1xh��T/���
A(�uU�VZ��P��-k*�r�Onߛ�騄�q�����k��#|�׭v)$-��m�	ju�]���hJ��5�=�A�L[{۞:��Σ^����e�d1��q��w>�X~��٘W|���8�/sm���tk1���F��Wn꾻�j�&�M8pK�CUVc��?vE�#� �v��_m�E@�d�g���F�n�@5R���"q��|F\b�}mB�D�)#�e)���O����V���p��#\q�sهk���yF�������(2ǖ��"�L��nM�Z���2��k=�\����۷��d-�����7���N:�m�U�X?/�՟�0+���N5tt�*����e.�x��u
��i�U�LE�j��
�ٵb���/����}�`3���0����l&E��@J�b黗�}m�Ts��x��
�־�{]p�%,��wɕ��s1L%����Oރ�ߐEdM�ܒ$�q$�v�՛knҎ��t��p#�.�y��s���r�	B@�p��b1p�\P|}�=��k+�X��)�3S�<ԃ��&MF��)QC����E�a�lλ�&~�6e\w�yu4<0H�h��y�w���ƹ��#���7������;��v���;�˸���Z���z��,O���_��\K�sӝ8{c���2��cN[�}|�lq��e�R��_s*�5-w �hkI�x6��Y0��ꄧ�Z7(4W;��Dd#p������<qo+a~��G��u��&��j�ʉ�0U{ͷ����5Πb�����,�����߾��Ė�Ʌ��I"
ˑ7�r������EWt_i���S�š����� Go ����Jk����)E߀�|�Ҙ��v rh����E��ET�F�53�עѤ�yI"읢j�x��.�J'Q�������~��{ H[Cm�+`�` �HKh  �   	  I.$�����B��Y�ѓ�k�4�vC)Q�3Pc�E:�W:�V��6����Nw
�����F7Gu�瞻K��:�5�:��t�/��{fU-��z8�r�`#��kK�͚���k��b�F�翑��n퍥.�v��ΰP�	�$�m�@5�a�3k8V�S����eV��v��k-���cWZ��cE��ݶ�lk�f���،����l���R	q~υ���>v��v�����u�i�UP �su�/f /��F�+���i8T-������� ��|��&�:���Ge=�`��;�����J�y�Q�_ �u���ح�"��y�^�l(��/�\�������b;e9vk|�i&�	�Jz����c����B>�A*���0)S!��`Sq֥�&!�b��;�.=�5�� ��J<�o��{��
R@S�2ڂ���7f�a)�\0�^Xu�Ǒ�wD쇧�|R�1��1;��y�3��k��vn����d��LK�����)-�T��;m�s���9��!f>3I����c-�P��	5�i&v�$­���;_�*�x��̣H����w}`���[V��I<�ƻN�s�;7%ɞ��3��/��3�Ik�5�+[r=�����_��2o�iR��`���k��4�%s�Z>O��(��9��W=�Z���k呒w�0�g�%���������\��h߽�޵Z6��5i8���{�:���Aݴ��9a���Ŏ`��I7���Ĭ=V��CH`*!,t�R(Hs�����Md�t��Ko?Ƽ�K�V:h�M� �?�3������]L?�q�jHbqWln�D}�����tETks�BJos�޷�t�y��wzv�zQ�_z։�U-�̾]{�Tn��#)I�oGslwɏ�1M��+�~���j�ƴ�zY؊MwpZ��>e�*�`uKVU���V�A�s����-���x����6=7wb+<�0�B���0/I���v�w+��ϞJ�̻��|��لP�τ��K�w|�i��$��l�][ƉWwcd������H%,펝���7gP���0��r6�(1M�MO?i��gO�1���N��"4�/�a"��n��Fݵ��(K?�6�+.���"���gFb�	�)��`� �wc�����w`�Kw����B��Yu�s�˷I� ��V5��-J��w1���a���-��������s
i�A���M�n�Ɔ�qx�Δ�o �|�u��ݦ����Ӛ��rZ[�**��EczU{L�A�`�|b[iu��ч'LٗKx���ksj
�۬G:������J���������|wx��WY�ϱ���������on�����څ����s��v�b�HJT�f�It��	VFP��J/s9r��R���=�]��S\S�V�����\>����Օ�sz��WXhn��N���VȮR��It�]c�۽Ʉ_F�m�6�d��|4���T���K�D��ʓ�̭�y�d5�qn�ev۬�W'A<�5��<���%��X�r܏+/���k��݈��u�u��ܮ�鲸����WKci���b�b�ZX��ڰ������dw
��G�����]wY��Y[:�t�3���l��b"�U�)�[N�j���g�� ���ڸ�6��*ץ���k��S2���do�W}�=�eBO�D�\��r�Ė�Oe�h[�9c�Y�*Wf_i��v��	9�tGwZ��3n�����cJ�{3��9������x
��:�c�m�q,�X;0�`\�Vr7ssj�PSf�׷ʖX��ue'��$GX����ƭn��:R]�(�r��q�a��Y���+{絅b��93{5T�p�&���i~�w+�~W�Շ�u�]��.��;�X+�뉲�M9�6���ʽ�t���z�����͢���)���;fTz7g��J�K&��)��7��0�w�;4�}쉢�(�E�ӓ�;���]�=�z5^��y�j�^{?dQ�s�T_8�ƻl)o��=C��ٻD<7������!l,R���Z�j�n�,��.;>����=\��\�a��S��p�sT�@�*�����#i8�B�*O4����9�Q� ��G��0���	p��Ht�������&�C�"�|�A6�l���w;���u�2�Y��È��ӯ���2	H{��������!{�Ӟz|��*�z<7�*}���Ͷo��*A)Q$K�8y�f��>�?ob+�\8���X ez��"F��gdf=
8e� @�7 zjOc��G�;~,3��7��"h�'L��}��dv��r�vՂ-w`d���M�ʨ!l�4��v��O�q1�J)W�����E�yv�˓�d�<ٻz�}�*�)���ûM���£,��th�cTȆ:��<:��Y�0�M��.z�[;�~ }z8�&�u���N&�H�N$�.
7Ȼ��W��î|nt�W��6�G¦�e~
����/F��x��"�N"�y��-���o��|1��Ĥ���h$Ut3����+�]�s�F(�a�|���Ÿ��eM�n	0�J@Jn��}-\��������l��h V7���0��q�%D��7��3�'��<.s�m�G}�wb����r)������:ᅳ���,�3�ۼ��&XN�'�5L�1ƛ�9�D�q덮��w�����p1�!K��GͦW���r8�:;���o�7�9����9�l�z�:�뉤bۂ�7�0
Ƹ���o�oN�t����>3���q��RH�p���(�2(�vT$�Wh�4�v�3k#�M=qP�sbǙ�4�:}��w���}�iy����ӝ�]��Ᵽ�4�q�!2�q�H�=���.b	㟂��&V}��o���Ǭ�����^�TL�<�8@�\f;���������bD��mo�y�f����Pd��n�[��'Q5��&��z�C�W.�9c�w�y��̮�ښ��S�oi$�I6r�+i m�   m Җ� ݼV�   �����Vݍ�_h�&��l�65�x�>fb�7^�p���κ�۩����#���t��=4��5�=F�f90u��Mp
rZ�=v����x���8{-�c	��1��V8lw�KX�Ś�F���#�Ni�gz�bv�;+��m���f�8�Q�i�6,+ĵ��m[��y���U���>��sn[�w7�ё���g��ڔp9��Ʌ�	�[�x~�h~�����b5���UwT�9��)�����Sz�kq�$��͘	�l�M'�ߺ����Aпv6�H�M�QN��8=L�S	��yM�Mc�Q��l�4���kq��$$�Le�%�~�Zx�`���ݸ��>�<�A�����`�
����lOO���h^_߄�'h]pVP�߂�6�Mݱ��ס"_g+���aG�Q�c���w=��r�y�&.�y��2i�����]�L�:)���n��j5�1X1��!����	��F���D�g^'�A"���+� ��&i� *@�rC�ݧ��0V�2�Z�V�ۮ�5�Dj�|�U�?��z�C��h�
�6�D�W�@�Cr���H�<�����kGG�� �m���$���kq.�=�1�ȷf���SS�������|�O���[��Y�>(}�c�Wn��=�$#��TW=�+ԕ� B S����9�ȋ����Ζ��pXE���/vϧv30x�Df���U�}���~�U\lc��}�b�V�*�
lmT.�j��b\]�f�kz��K�����\H;6�rU"�.�*i�ay�v�-�M�R�z>�"ߖ���8�C�]�q����6Яw��q����
��"nH�B9#�WV�}4e>"���n�0�LwS�sM'��X�B��B S?lDN;���F^χMrc<��Fd[�w�4-�����n׌{�.����&�4��k>d�W�><�О��;��Ku���V!�D�#eS<�
��+H�s�[�bF�,Iē/mNq�u����0d��[gr*�Ӿ��v���S@<}O��y�*wf@��.z�[�o��<}�p�8�cU��z�\���T�q�dr([NH�l���\�i�6x�n6*z㨳l�i�z��n�����3"�����
p�Ypg2�&��Mp���O���@�E���D�(������m�G��n��Y����&sbj�y�����6Wk�_�qBYb$������:#��-��]Ĥڥ/@��D��	�ťf5��"
���bN�� �����>�i�J�ʷ�Aj���/� 9�O�l�0y��
q����lT�=m�oک|��LLH,��ZD��߫9�B*	F"lKP�9�E̙�{>�����p�ne�,�wǪ$���r�@�m�/V�^���2ǿYQS}�/�c�ᆪ�R�6�tL{sӌ0�'h��L�6��F�s��{���5_���[�8�h����io'��W��^b�Gnܷ���5�Y`�)�l5�W��y���}������������R4�9$�Xw�_0�E1�zt_H�B(t�"$�T�:��C���:%���!�#��v���T�����5�U�GH����>ۮ�����u���i�mq!��N��d�'��t:�ȸ.�pr��e�]�),�m�)��_��w��N�M��K�YcU�u}m�V>VC�r�1��\wR]ms<�:�i���¯�~	�ɂ#�
p�S�Ag0�R"��$��@+
W�����R���WU�s�} F}K���|��N���{s�������x����z��x"E��V���O,�����i đ6�E>��Ѕ�`�(�<���'����K���!"�ʀ�=�+8�"����	�^�Ap��0���1pϧ�ȁ�y���Ad�"m��/��)�;g�FD���ʇ�x��0��� ��y|aF��ꇏ@K�R�$��z�I��1���
�n���tM��DD�C�����tլ;���r�Mm��pT��{�`�߼@ͬ��5��������<s���68e��:s���:�i>`}���"�)�@�mV2�^\�z�Y�-�S�.{��mG��#���M>Dg�M����x�ユ�xx��䢊�ړv�nΟdI죎�N׮�]�Ŝ��$�a��õ�h���9�O�ߏ�[,N,���z�)@N4�,����{Q ��T{��E�\P����Iğf��d]s�R��Cz�#��no9.� ��p$$��>���9���@Q�غ;jX�m�IA��7ح5
	�>@�b^_y�� Q������5�O�d-w��D�����o��$��F�m��Cآ'��#.*w�4W��Ϗ����k��4�H��QԔ�Ok��&
*���YpH#���P�[`�M�04�ď;xB��r&��6L��s�A��8�/Ah0�t�Fϛ�[����>�x��=j������#Ց��[�;��0�n�E��堽�v��v�qw�:/�!@��ة�����D�̮qQ�c�,:r��ad7��"�+�G��hV��9�'<u ��W��c��~#�E��y�kO5(�օ�OU}]2��Mb�W��.�#�����' Wx#�Y��uYS��[)>Y�+�	�әr��I$�h��Ibtm@   v�I �P �6   mt  &�ӕ����p�[�sjfD�l���=�'���=�ey�������u�s�(�n{r�>��qɽf��3�N����m�l=�Q���m���v�˜]�gp
�nv6ɉf拷J\��ۛL�4�k�sՎ��՝�MO�x�����w����"�ۧa��ӻ:�ĵ���V�#v��n1�V�Z�&#/;�a��M˄�vW��H6$1��)3'����:kŉ��M7�<�"}��!�O��D?�*�8ϫɀ��' 7���<�;�d����5��p#�t���Yd�
>����`B����ؤ�b�I�\4� ���
>9�{3�p�d��4��q(�,�_ğy��<� ��?�d9 c
.F��^�[�i����p$ L��X4ߤ�p-���LC�Y*@J��٤1��8=�~r�xY��o1�x�l�%��F�*��X	�b���T@֗"�Te	(�Ǩёl0��~� z���d>ca�-�|��R#$)�#�a��oU�J�Q���}���L<���oa����~��❉�S�[��B>GGٷ>�D��lQi���������~Qq�R4ܝ�t�h�vA埋$�oE��� #�Q�>??Pa����T�u�|���%ϼ�N\��'Z������r�	ſ���0�O����'N���]��Im
�;n0��cs��h��$ӷa7d5������պ�K��Ȑ��ȣ��Q�ϒ`�!�5�8׆����L䁮Z�/�>`�|��|�����Ε^}�B�g����c���Mh�P�H��������N%"e1r��WOp�,�� Q�d�M�sπƸ�+S�y�ϻXOdc
�hҔ�(�/Ue^�ҷ�	�#ѣM�:�-4�z"��:X��O���K��.FN�o;�i'�{�~�4ΨC���2qpLy�!1�r��e��s�ߏ�񩞯W���!����v�]!��i��rD��� Q�c��	�}^�ݾ�aC>u���{�� (��
6e��c4���}r�[�$���7�px";Z�����4&�	�\�j���� .?�|�h�K�]�ً9�~Dx��A	����C���w�Sχ
#��!��.�2=�0�q��ǗQ�x=&Suk���H>l.�ⷆ��f`/U�����>/��|��D�xֆ�0�%�K�>���$�>�;I��6o4�i��Li��\뙕c�9���y�[�k�a�xiݏ���q�A�ލ�1p><G+�Gɞt'��0�0)�S��N�+��࣎B�-B�rB��t�\<�[���pmsɈe�9����q�n���)��I�@�h�őg�|�a��o9!�����l�$�=��ްHL=g�y�ӱ c�ؑ���)�Z��B�>1�:���y,H<D󫃤H�8c^�0[.H
q�D=fG�z�� �<��:�yL3�<}<!\���yΐ�	���u�1d�υ8N9�8Ȣ|Q�Eǈ��>���y��j�\e�G��[���Gqm|�%3��n$i�=������!�,=D=�K�q��|�I�����Ζ��2�?�:v�v��{a�ޣI(�Il>t��%�<ު������:��<iP�u�}7�Y��S��X���O�Ԉy߇,���^u��><��@>���Htv*	0@,���x���H8W��9 �%n6�u� H��a��:E����0$z.7p}��@����� ��c����@�O���;���J��'�t�jqs��F�j�} �s�9�69� ,<VF�� apt�����2�e�q��"��H�_��0o��"A�[xKm�܆�x�Wb{�sOǀQs�
�P�� ]:�d
!�0�����kW�g�G������@x�������qD��Eʵ�n��q��!�ɝbt]�.��.ސv5ϷU�/�#�����E?ww�}�{�Q�:gyW��-�dz���p.x�
�R���4��|b%���y�UQM&y������G$��8�o�r"@a��#�x:g,�Њ����l�g
m����z������.p�y�a�:�
���D�ͮ3�+�O>|G#�	��%���N[ �#� �d��ܫ�>�.6�E1��� t�#��y*H�J�E�\8,�d@�<�@�����n9#�@�A��(��đ秮yl�Q4.Xc�8~|=�<��xfU�g�=0���L����{΄'�a���r� ����x&jH(�
RT�����<�x�ǜ��&��b�|�|��O#d0�� d!�xt-�C�P#�C� Gޒ��6%k �p D �u��2u�7�
x7v0��T���*ܭO�$��q�m��k,2Of�ֵӾVr��G��O!HO�ǈ�D9$zH�\?F-�W��N(��#�;hs�1�?�xYI�g}���D.������>�r%��i��<�e<���s�,��}�>���+�� 
#��$�t��s�\���sO @�yHs�y�@a���uW��x��6�2&[��$�R�vϊ�pOq�ۄ,lH�f�����\ѱ���(��6JC#N9��0��xG��sO � m��\��l�xu (��#�]��y0�� I�� G�Q���[y6��R��Ȁ�<0�1� yr��,[0�>���>��,�
$�f���!�#2(�q�(�y�cC���y�!�8�GѢ�����2dqxb��#�#���n�9f�y�G��f�{�w�W����D>G��@�fďa�}����g6��|=�{ں��p����F8�s��N� :y�G���·80���9����#��y���<��y	>�^?���f%�cG��{�S^0���E��zu�>���x"<=${÷3Ƈ ��4�9�q� �8��C�&L�C06��� ��p3�9�������G���� ��#޳���| � |=���$a z��>��J�y�84�ixO9� p�>M$��2q�!�^7����ou��*�>����d�m��3o�<��`����MgǏҝ��L�������!���fG�dz�� �<���>���G��5q��d��=� �� ?�R@}�$
���R@bR@j��H�O�R@~$� ?*�� 8T�JHuI� =�$�R@|*H2��I�1AY&SYb)�ߎY�pP��3'� b�(����UR"�*�eD$��J���
�T���T)U)R%(i��H* (���J)M�R��    TR��(*�T 	R��ID�(D *  ���$���(���R���
IIP� �IHD(	 
RABEwJ�myhU�S�Δ+����*��k�m�;� �R�n{<�U.Z�)N�вҹj��\� =�e�O=�<)Kn6�aJ(
�()O=��[V�=�{ڶ�x��y�[m����x�4�;�,*�r�L�՜MҶѷ���Ym�\�¶�k���m8���kj^�%R�kJlSB� z�(HT%H�P
@���mYWݶ�ԶܹuSiWy�zZ��˧YjÏI �{m5�.����mźhl���z����yK,� Usޚ�Oy�xm������	�Mj�[q�:���vՖ��@���*����Y�e���m��m�7{k#[n-�JR�=
��[m{׽�+mm�{�O4���c%/z�R��"	��kW�= � E
 7^��ܵu�Z��g��Jsj\�m���J��J
�R�V3��oyB����ګ+o{u/*ڛ�����*��5K*��r�z��*�
дQ��H���z㢒P�w��I㢗�Gz�R(�Wu�Ex�I�;�IG��yeEnzE<�S�'u����$O(�6�K��	�Z��uti^4�����
H� ���t��8�{b�I��*�ĥ�q�J<�w��^]�EzH�Q���5�<�tU�i#�n�%f^1��It����R)c{e$z<sQKĨ��#%$�c�s���/.��:(ѹ��$�q)�B���$��y��(��z��Y�)*֮w��UJy�(���C�n����e縹�#A� 
�+[�= �J
QA@�"@ 7�ePs���Uto/pԲh���F�G�E��R"�=�Ǡ��]��I9�u��(Q�]ȩ%"\c*�����7]��<����Km$q�OLH�^�T�� 4�^���Bٶ�v��^��ފ7�R��q�]�=�O�\[Z�z��kgۼ��-��*���B��w-:y�٤��ay` :<���W`  5O��%T���$�J�41���a4��M0=��#"���@OȤ�%* �S����������?���?��<��yp/��gDpC���;#���8 �9�qh������9�88889�s��� �9���8 �9�s��s�s�������9���������_�q����RE��hhHdmd�k��Q������̓M����0V@��D���Lo]`��Ky��h���h}*c&�a�Ѳ�?^j���^ZR�F5&e�E{���ɻ4^��!�	k�jV`�X�׺�n�UbSh��kp5v���M�aݺյ����w@�8��Khə% �쥲ANBDӑ�J�^T��0�=}�m��R���SyO+�ѥ���lbZU�xct��ÿ�k�pv.�n��pe4��MՋ�&&6�8A{z�͛�E�An������)���,	���-�D�h��ܛXV�vm�j�Z�#�uww��3%�(�������2���5��t�;�.,5-W0k((�p[��[�����a��n��w�
ɉ�GRz�A��M�Y��p6we$qYn�eZ�g��*��^�rP�U���4��[voj)v���K�A�v��#�e+������otp�̥���	� ���,�v��F�L�#Ʈ��%�׈�R�eM�5���^�k��«�p��ơ�Ҽ�T(o�U��[0!�6�fj5��]��͊e)vq���5�q��sn�汔�73h�����Vثifa;�hQ,��-�M廥���XCUy1)���r}6��7�a�8F-�m�q64�+��7�a[d��N����5�S��MI�(L�<������,5a��s�OiV�Yh�&w�`��f`�y��x��t���$�*Y��)�ai�Y6�Q�X�v[6K����Tr-[��
�#�zz*�5���c%<a��.%uf�Ӊ��ۦ�/�˖,X[!w�a8.EWQ��Ֆ�����S��7�4.�j�V�����s���ɇ���[ū���*6f��*T���2r����u��(㦃7�֌b[Z1Џ�MuUua�u|�'�`�a�*hA�CI)`5X۷�Aص��5YP��+e�d��m偎yF=l	�*e-��:*f�@��c �4f��Q�]�
l�:�E��M�E�Ӣ�jѶj��r$�e�X�����N`���7ti��[Uy
�����������=�e ����,B]�Jﵓ��3���T�F�����5e(�����e�(V\���/m�(I�ҒW���)	�V�i�M� Q^̽��8���vFM{��R�����Z�(8�(ܺ/!�GSX�wN��b��zSZSuf�k�v���;�2VЕn�,���J��oF�O*���U4���;+tm��Nm[ƕ�X��S&iNH֖E�g6�[$S�rn;�mpd�o�Q��%X���-Y֒yw˭x�IV7I�a�@DJ-�h���;ae���vD�l�9`��t�E�Y�j��7�^{VdY2ވ4{��F_q_����Ɯ��W}��{���H�0k6��W���K�>��55���m���&DQK�)-3eTt��&T��LYi������R�h�zD�X�5�m��T{2�A�)��󔙈���m���FJ��7��5���u���Y��"��mY��$��k���Ɠ������jw��a=L�Y�ܖ��,��f��Aj����m��S1��� ݚoIw�Q���{��o0>�sD��W1#���F��`b��5�L��Nɳ�k]�&�8p&�j�L��R�ɧ�A�ۺJ+�lmhr]D�.�*	�u�2�Z�d��-��4鬭��͎i�=î�������d$�Z�dQ$�2�(d�C���PL�De�uW��.ɱ�uku��$Hőq�l^�`V��tؗ�oD�t�Ҏ]�ƍX��A*Q]o%��G&��	��,�����l�*$V�(�7.��"e�R6�b�د�Xq�9�����SX*���A�꛹��F�kB�4��&To&^�"�2ཛwU`��5iCwJS׹n�k�f���m�j]h�����9VP�*��\�+�0�:�	M�).�:'w%��n�J�Gn��{Ť�Щ�ɭ9-(e�D4�vE�Am��f�]�ȳuf�hc�w����b�m�l�k[[B�͹�p�M�;���ݒJ�2�	㊬7Y�Al��<���� $����(��Q]&�F!ւ[Eڥ2�w�6ʛ���ޜ�L��-e���w���e'���g���;�Љ����4%h����.�3��74�-T
�hB����7d_۸%�b	Z�ˊ&�(��^^�7�DJO/Y��+5�5�u�.�j�͍,sfkx�킬��3����#�7�[ʙRP��Պ�d�1���t��!�FH��Qf�N��f��5[���gI�6[q2Ϝ�EM�����-�F����%ܰ[Ú�D!5��W�q\ �C�Hn�FLI��1�l����Ӥ�7���C���!��.����R��Y��3���p�jm�#5b��6B����L��6���0�5s@�%��f
�Xcac�w�հG�����AcՖT��Z,;�YUmА����{e<īmZ�e��bW��3S🂷FXb���S�e���1�i�v �(���S[J�È�f�v�qe��{Bŉ6h8L'HYoi껱Z��Vêj�tۧMc�yt�0����n��/�H�d;�ufh�i�,l`2+m�j�DE�o�*�t2��C�2��Xli�ù�	��l��&b�7C�nf�����ܘ0��j�ɥ�S3r�'��kNmȦ�����*m��L�#��h�l�В�f؉�E���m�6=e���bcH*�Pj��s%�3>�wX��c���[�'D�4���vK��f�;�hҷ�p�+v�!l�x[-jpB�q���(f=��I�5r�Q��Вe�J��V6N�q��+r\Y!V����-,�T6�{u�F��8��i$�mk.l�zi���vv,�1`lb�^��ݔ�۩��ؐ�M��^�����5���f��M����Ćʹ�V��M�:*Lu�2�da�2卙Fms%���^�Kz5(��vܢ+~�X&���Q�ʒݼ�{���f��3��!/M�y."+)j��M)#O4��ǘ���m�:l��@�%��Y�������,�8);�S�摳+Zz&�t�V�j0��k ㎲\�[����`�����^�8� 1��OF�J�{����S�n�Z���.��/M�:���e�\���fQ�����d0�
��^��-4mꪥ���K*	�U���įg!����L9	��qY�f�t��9O'*���]��n�8�+t��v��t��B8��0����L=��qĆ\��9*S��ݰ�CZ�F�x� X�n� /\�ڶ�6�UC�]���p�H����Z^�7�B�4,,����3-��& OZ��.�n���F���9�S  f����oe�D�v�虝"J���Xf�ekz�MRƦ�va���%m����K}$��4_��]>y�a��9�)51�u�M"�4��\v݋�N�,�`ƶ�1�����׹��M1�1h��m�|�[TI;��cT�b�4��94H�n�[JMz�$�r=�h4�v���2��3�n;�
{�"��QJ�8�{vΙu̗B)�Ћi�ƭ���A72VC�aZ�id�h�xs�;��ł�Lm�q�z*(�DZ���ԫ) �+r�z��t�a�{��
���e�\ˡ�B��0��1(0SX��m��2V/W+)}[��z�kL�s�������ܜ;e���,ޞc���7W�w �,�"�Q��l�m[(���4[�J6��}Wu�n��&9�8{z�;P�G�F����F`3�MS$���Y2��otj����|;X{{J�{��3}H�y{��s�+c$��-��Z'�D������%���'pi���
<ۻ��xd3#�I�RkE�`�+B��a�SlS�ݬ�KݻV�C,�&mb�!Gf��4ڶ��LPL�ă�"�[䥬J���vX-�D-*�ed�^j�gtNm�H|n���)��껃NhPtQXm	�wV��̽,�BX:Eu�̨�1i�n�,J��(��!u��O�&T8l-�g4�#b*͐���XX6k�7��F̢�w��V�s�(e±�r�a�)�5b�ȕ��u��̓Q�C5��*44�z�BE
�)���f�o�
�(��u��^�t�w6�\�e(#�;�0Q��i�w��h���B�¦䚤V���+���D/L��q�0�\x^�ML�[�h��\�^�j�F�Sb\�okV�VDJeQ�RtM	�C)��/'!�s`�)!nͽf"�������S,�|;�M�ucNb��vƛ�Z�ȵwnn��K��a���b�8�Ue��v(�[MT���|k��b�L���6��m�E���vY��^�8����R��y���g,f���H�`+;2�	w���c30��5+�xt�l�!V��N�Qf�[��q7�i*�"�CL�cmԥ��ٻ8���ۚWy`��Rql���G����mg����[ܶ��EL'b�J�{3Z��ˣ|ԸmGʺVo&�ɜ���[d��/lR��M��e�5��F�Af�{+DD�.y��0)sn���Z��-�+ˡ�7*0>ᆫ��P�jb���X�-�;��K���Q��.\�8�ڻ�(�w!��0^����olT��|��0�Bx$��֊)]��]�j޽�T���pʾ2�N�"Gg&�M�e�;Of��(@7֦uE��՜�zr�zbd�W@�k�%�gn�;;�0l����#0��y�9���t���ذ�pv���a�Kve���嬵׎�/�D�+�]q���1Qq��+ t����[#����k�_�EZUt�c�E�tҹ�����+F�l�B�=���ܸQG)�P'�F
k��
K	3-�f+�]��)�E�5�$�R�䗕f`���R���E��]Q�[E� �ΩzyD�$��f��ɻ2�>tcn�LMP�cV���l�E��0-Z���k%d�N�1��vm�L��U�й�Z_,<������{d���[HY�8w�����-�lC���d3��N��w����c�{�Ltt�z� e�j;]��R�᫹��]�l��N�s!͐��a�#����dlj�T!�b�Okٱ��Mv�;��h&2�\�$���S�V.H�D��á�Ud���/`5�[s^e�P;	M�qP�NV��{��d[�)t�`��f۸�P��ٹds&f��f���ќo��W����֤ ֋"�f��F ��d�b�R�k>���@B��&�ʗ.�T<���U��`.Gf;��g�n��^E7sX�V�rU
2f��E���z�$&f^-��-�{Zq��rY�cV�ȭ�1�1���qF.fo]*������Օyh5s.�lL?]+6�[4lB�f���ݴ��R�V�x�R	�j��D=�`u&u�O*�F�ˈ�t.4�-�z$QR�^Л��d��4�kh�]ݜ6�u���ufI[��
�0  *ebu��+&\��bɼ��b׮��Q;2�4u�0i�P�ͻ��P%cC"ʶ�Tʖ,.���D��*�`Y�n���&�6��غ1�W�U��7�/c<6%����0��m�ӷ�xv%���N�Ɇ�����V��`%"M���
�%h��/��p彥kh��n
2��ػu)	��x�Y�_�M���s`I��a-��1RJ��b��Ja���3#Ut1�ȓ��5f̑֝��&7�B%U�b�+�T,��NRh��A��fʔ�3(�eb�U�L�E�R��w1DI�A��-}�ܝ��c iZ���PLm����y㼢��_js�o��[w����HUϤڻ��]u���f�@S�4��m �P{D+�v������2ZC^8s]l�ّ�3{�H��6)���6���TYHm�@��۬�w�4&���2�v��ĥ-���L�2�vB>�J�ر[�� ���\;3��YlV˫�:c��-R�In�Y�R�SJ,[[u�Ke� x�[7a-��mfMi��ݠ�*R�ڼ�Yu���*�+��[�L�K��%�V&ܱ�nl��ɩl�jlJH�KZF�l��m�CffV�6����
+I���9,����X|��
��{j�e+B�۲ֈ��z�Y���-Q�M�*Kx�y/0{(�Ue"���E�������_6\�BgD.�=�F�ڛseTM��wf���Րg;���멮��P�o�2Gq,��w�C:+�Cv9�u����%K2�8 �;�Yk�n�=�b�ApWM0������&�v��(��Bk���ݥ��Ze�z�u^��p��l,29nV�g�SY-��c8���m�R�c+mi�5#^f�"�*7�]�FnU����-uo]a��1�;�v;���r�a�M��F9G�Ű�u�������t�ga/��1���u�n���@60ʄ�Cb{�h�V2�e����tحl�YTt�)�toR�7^���M�j�U��sC�h�çw7V.O��}�UU_�_*����������������������������������������������������������������������������������������U���j�������ꪪ�������j�����
v�����v�ꮪ�U���k��55Um*�R�UUUUUUUUUUUUUUUUUUUUUUUUUUu]�����f�UT�UTUU]UUUW*��P���%������ UTUPu]*ҭUU!5UR��ۅ�H@�DP��T����+pMTPUR���#%]uU*���UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU]UUUUUUTJ�uUU�R��YL���uz��a��38�d3n��Ae�˶B��o:�}.�6�݄w+iB��51�"�S��9{��sk���6�nP���\[��ۍx9��m�%�=�.��l3������k
�B�Y�\jж@y��V�m�`��-��s��]��Yg��it�ef��
1��t�s�H�j�v��+��;r�+��kDZe�<��d���l��i�d������JF.�v|sWb�m���woc�xV�W��m��,\ř��3`�)PY�s-n��M��z.7\�I���ީ�P���9v�vT�)�0]3��[[(:�nd�΃��瞪��]�GGKp�k��aMqt1�P��,�Z;+�ß;�$[��:���<��nk���ۖ�F��s��8��lPq�f�ہ;<�ˣ��fcq=��n���r�M�s⭻3���t\5�#h[-e+2͍1)�X����;K��giL�̉l1�!WUl��-���=�J�.������.6�cc���q���s�9�a��g��a�@5�\F�Gn���M������䝺�����m�}9�Ng;Zz�:�{r'l7� 喴��L�rE�e�1��mm��o�ZS��BP&�`��OOgel]�uM��4Mt&�DԁXf2�f�V��<�/Wp1���;�r�G7�)�n�;���N��㝕�m�p���l�ړ=n���n�t�5�tv��ˏ'U:Ҽ�:������9gv��ۅ��t�P�^�2JG�qw���`g��BrH�(�E�Vݣe';
����������%������!;�tx�u�DD���w �v_�'����w��ve�����^n^2��N��5�r�����2`�>m5�����INwi��.����V��*)-,(�]`� 7-Y���[�-��y���q��K�Lq�[.^�Hhv���%��(^�t���;�vc�=p������W?m��qp��j�m�'B
��$�e���]WO=gM�����n�6��mg::�UN���i��f�mg�ܽ�k��v�v�Z�]���|�κ2続7jx���uz�����Ħ
������8T�r�n'�5�v"����g��ۗk!�ͼ����t^z�83���븴�]q�|]n�[��=pF���0$n�ӳvy�iLx�����2�g�݀�t�y[M�� �KH`#.s��B*ҿ�n���2�ܰ*!V�Q�Lܲi��,�W/
��dSm˚��e�-�'nl���b�n24��5�ۂ�k1��1U(�0�4�@���^�y�sd�o=�uʴ�$�'�>��
<�zp��k��w��.�VgXR-�K5����	�a3Yl�]abV�J�{<�]'/VH��e��2��h�G��uZճ˶�F�c�[Ǖ�����q��ȼ��-e�#�3��d5�:�]�^<(�ڛ�9⣝�08���vLW�NFb�6��lfL�ԛ*�-����B��"� D�{���v�.���ֺ��tYP���K�j�r4����Ǯ�"�� g�Y�t��r�s���� �Ŷ���R�]F f6�-&e���JP�������}������6�!/�;nw:�;�B�v	kƚ�C)�i\"h���e���\�N�o�ʵr��ZL�n:�t�g+k�9���붸 �9}������6x�φN��^��gz+��Vb6Zmi)��R,�3cfv���^jC^���Q5��`��XU���Y�G�b�ZS$hj�:��_k�zڗ����c
z�u��K�����c�+�eu�#�s�7���v3	����#�۴����ۦ�'=5�yꣳx�[/:���=Gm�h۩�γ���ى�Xp�=q�^=z�>=k�b�r�<�1��Ɠ�ی��jWZG�
p�LU˧u��4�r	���9�[�ݚ�Ѭ�����ܳ�{�^	:�n�@���hV䔛�&��X�X\̸[�n�]/��l�X�4h�p)	����c�1;X�-l��X��Yf���YX����������׭�+n���R�ӫ� �v̽'�i6`b��n�N8Z���͑P�����Ϊ�J�n�N9]y	&��w�i����="O=n�a���3�o�nTÌM�z��ϊ�N�zU�cn��]���V���.8�(saq�S�8�ݷI���,k���`���d�;1�[�u@���sָS;���U]v�����F��'���3j:��v�x�l:��u?)���#sL�Hc�XJkfȵD�R�j�C��v겸n-����cRt��e��4�)���`�����E�1�;/�7]��c�Rh��9�h�V&�pn��ς�x�`���� ��Ӥ�֞6ܦ�.��������A\��.Ss�4��7]x8�����<��b���K:wl9�+='i� 6�2#]3B4��m��u��nw3��M�<ǲ�P�6���5+;��Nv�p�a��*YHKivx����N�7v�ph�B�M�k����P�8,>w��*w�ݱ�z�hS`7n���(ٸ��֠�����ƯY�5x2�=���2�7�bB�A㩊������Y��W�;�Ӳ�mq����m���'�哧����E��.�p\�� A�ձ�	�Ś����0pZG`E*�� B�)���:-�zk�rdv�����8׵�Qc��A�1��iR���5�i�7 ����Hhb�]���3u��pq��nv�<�RH6�ܼ���^i�F����v;N6qP��M��C�aȏn.x�J���	��KFW�&��/b��ƶ��↕y��� hݐ��hP����K��FѴD��Y�0��n�gN��ol#,[�n2���Bi�I�D��\6�
�wo\u�lQ����;�3jʞ1���p�+���3b,��\�7��RHr�����3ۘt��
�01I���$t#l��x��z�Ѻ���y�<F���j!@\㗰-ڔ�
M�]kll1	�2�OM�wC�w��k���Ѝofq���p���:���zB�ɺT{p灰�O/^������x��'X@g9�8�`nu�f-	�]��g1V8��%`d������=��3`�=7�Llb�8�]s�vN,Lsc��b���R4H��n�i��n)�CZ����HK�4����F�=Q'n�u����wm08��ؠ�Ңp�� MZ4%Ԏ�P�+�kl!�M���pj:U������Q
&�8cy��h0[��)bn%(����xplb�h�e� qm�F0�Q᥀G7�#yV� )50CQ�Jٌţ����Z>j=v���㥞�۶6�w)���۩뇇E�7����,	��ܶ���Ht�е�-١�(�x\nCGb�q5�x�����W�m�㶩7�I���'GFUoqw;Orw��osb��V9��U�N�.��,M`��P�Wh��kq��ut�`��Xm��ݑ��]�3X�%��Nzć`����@J��(����U�^i-�L�(�KeTFcF�FΞ��+ks�
nv���.�谅�v���q%j,�v��Eij���h���ҳ��>>WXkc�����]�	u��v3u�vg���:ٷS�h�)��yh	�u�vn���x{n��.]��F��c�i�(sXWx�
��a���9 �ۄnى3fn�X���i�٨��̰���uےN+C�Wu�h�%�h(�l#
i�ˡ�������`7?�=��oF�Ӈ����؀��� �0Y[w	e�m�&nk
ҖX�4K�%ZJ��P���!��u��#ivvx�3IHR8lƩ�#�Ľ�5f��5��$�D�:�{�J�pb뱆�D]-���gڗ.�]f�u�����6��i�!�֨B�Xc[&#�Q�\�"I]�a�'��ֹoS��
G)�7�Iѱ��\j��벓�a�<�G���YɲOO���v�uȖ��5#
r��-y�kXI������M�n�u�-�ZMӛ7b�km���y�]�'U�Wf��ڶp�-�U^5Ӟ�;y(,�N6��M���	�)�ۃ�ROu���m��G�m I�C-�xu�����7b���W�#�=xx휱�s�nFW)���Ac6͍Մ�Vڎ֓ZM��l4u���d7[v^�K��P]�y'6v��
���)x����cb�7�W.���Ű��N��1�붢w^���:��Skv��r׶���<&�v�n�-�/��j������魺��[^�Ѡ85��;:vC/��췬�gBr�t���9z:ñ�v�nzV�y�u&N�XyV�V`(b�aF�7���f��.�Γc�ƫf�k�e�������픞�nx|c@"g�İ�(�̥M�4n�Il�٪��%Zbąyx:iykd���v�<B���n����C;��uo,�ahl�Yl1;��A/��=sه�g:�gc�=x�r>A��Cc��g� e�Fť���4`�X�ms�mj�	,I��gg{it�i���T�N5��pv�^��ua.�B�v�CJ��i. ��=�|���٫nu���ޚuHcGc�	�H�w&�:��+�.�\��7Q��r��3�Zx���g\W�9�lh�t�;
`�X<v��'@�vr�v�-equ�?{�889�s���8 �?��p�s���?�s��w��__�_�UUUUUUUUUUUUUUUUUUm@N����UUUUT�z��S<+�bNB�TpU��5UUUUUUUUUUUUUUUUUUUUUUUUUUU�eY�=�$�x����:{Q��lY癍s!�+bm���!�� �k-�h��cpUi11+�S��u5�)���K��w����:���ˬ���0�`��X�#Me��VC��]�b�r�;��$�y�8�`��K�Om�܉�m�-��dt#[�"�H-�R�P����Xnf1�}z��`��r��e��m;�]F��	c�����2�,A˙�"��e)ds�1v��v�m���Km�k��.��ݪc�z�b9��z�*�޸0T&��	�quχ	������M�J��I��$+����Э����Iq0\��1���[ Y`��	R�+ay�4�7��ִk�nZ�/P�����M���j��pY;4����ep���=K���'[�=�;����7'(���<�؀�i2�c
����7c��ɸ��g�n��/!t�;c�����:� Cx`p�n��{pr�ԋ��<��/T;�����8��cmW]��g^ol���i.��{v��Ov�NZ�{HL�SF��-=�^)�y�6�������YD!v5�L��� ��8Zd��mi��Id �����\������U�2{f1��d,��뱉�����r��-�nw@6Z�W�>X�q;�k��ur5�`�����/���0�uiF��v^w����C���I�e�7�i���O<OZ���M\(d�c������Um�Y����[������v�. �}uқёK�ȸ�q)�xqc�Ũ�5��U���k)��ݲ4q�SUӧ4�M��Kh�ʻ[8��x�i�8H.�6!.��%1�uu�t$;[�n��s�>�ӎ����m���F�����tVh���
ILV^���u�����$Ƹ��"�, s�q��s觋q��m,lۜT��۳C������w{ǽ��*���^ ��l�%j����Q���i�X;\z�%��C��zq��в�%-��M��A��!lY��l�ENcӍ�CAؖ�y��m�p\ө�v��g�c�dS�+��.���䱜���7	�s���;���5����:h�e)��V��X�t�^]�cf�u�#�=���O����퍁��r����d"��az{�ϡ�"�Co=��܍+�6#(��[P���U�s�Ȝ����;����w����~�xb��j�=�k����|q��{���c��;����$�����[�Ӝ1L��V��/x��'n3�L\��{��Wk�=���e�S��E6�� Ph(�ݬ�zڗ�wn�l^�&-ͭkG�ޯM^���Nλ&�-��(�R�b6�o=��Vu�߬��P��Y�H����X^�g�Ǹ9�E½WU�jh��S�880DP��Cs�1z�U���ݱ�uK���<��Ļs]���ٗ9j��h�Y��K=�mHZ�& �Ee��.
�Մؤq�Q�l$6����/68��1��e�\p���q��M�6��;�}���ی�&r���y��	p1�Ƨ����k0!�?f"�-���m�NG��0E7�ۍ�j���"�����/�����X��N�Q��&�GP��,��}!�Wص��(���'����ʳ�]Bv���K<2}�6GL2j��L�t１@�5�k-����`��\"G�7l�/�^��yg��W��tY�W52,�;]5'��X�v��L[�o&��X���7$��'U��T��nm�ف~<��=��3����z�0zؼ�oN��V׳Ų�[p��(�z.���ϻo��r
�b׎�Y�ܚ��,�3�;PI�׉v�<7���z��w����!>pܵ��3� Hc7ML�Y�S �4G,y���,���㗃�.Xm��/���]�6�#m%��ئ�z�gp�ٗC���xV'�s�<�ے?�A��T��0(�f�G��id<{�(�~�Xrp������}�(�����5Y�DfNB�Wo@��
$�=:κ�^x�{l���]�?��k:�k�.�/U���9J��>h����e�:z�K�B�,�z�Z�f\��2���OOj������d
P�n��d����]�zfZ���]��e^��p$KB�l2�B�K����9��3݇���l۵eU�������$GL�7��������_�i(#e'�`����{��mN�鱺o�\�U�{<�B������<�Y�mr�ݫ��v��i�����t��b/�,�����CMZF�i�n���5M�[�R*��I'�>�Q��,ɼk!�tM����8[�܈�;�ڃ��{����t�����q�(�	�%L���4��t�}�����d��ۏ %e�w�ʒ�ז�Y�Ź{�-���W_Zn&�',f��.fm��0Gd�6E��n3w�U��/�y`��lF��=��q�'٨W�Ld)�����H�e�5Q�d\��|$�Y��'���*�D�s4{�fk�����^�o[>h����^J*���+1�X⵭�Y6�ٓy���&��m$�,c�3�L�w���u�mw�;C�$M��`r�nf�,(�/{���7�N|Vk�gx��Z��#X"���Sn�c�ڱr�o2�{b�F��6�LG�e%)��j3���eRy<���Vr����9*N-qͣ	�$9�s��eߣ�;�;���jM���Z��ˣ욶�|飑r���3.����NCI��$�1o]n��ָ�V�Śjo#��Q��7�T�t���F�-�Y��}B�fF��vv�Ya&6�j#qH�g�L��ޏ2�ʧ6�����	�S���p�:,c��sn���0�[iyHq�nC�1�u�������[�sY�ݳ���Bd4�އsi��,�S]1��t>kO�ϔm���ڒMU�����a��{�_|Qٱ����;*v��w&��Y	��ɭŻ�=|r�����sz�IӇ�vou�z���D�:��c'�-�f��V��V�Cr�3��jjܡ�7a}k���!������ٍ�Q�c�Jb�������%��������l٣�8��K�H �=��<�q�n�eN蒸��-����u������Qo6�絘6�ȑ�\��2��lK���
�%4XD���b�S	{nvȷ�z⭜W'=s��+az:ܜ��W�`��3S���;f���5379���n�2�kp���[�=����\&�tZ+v�\�nS6�D�s|w/�G\�5ئ�NH���ۮw7�y�@D���x�#�) )%#���X��k�ڽ��iW{qE�t������Zާ�W�a�L�t�xWn���wAB�,	�"���j%�׶�WM}�񭺙q��q)�����Y����X~��
 i>�ۜ���$�07�;��uBo��+R*����NQ��j���|='����}5m�K�v��]
Wt���[�'��շ��|���{Iڷފ���{��1ޘU��̦�d�+}0�3T���T�k�+�B	l2�-��5�ڷ\,B�3\��1s|��=��v��֞=��w'ة"�/S|phݬ���$�9��Z�h^�^�l���t�+À��m�E��gM�ھ������5m%7����c���l�&��HzwW��d��ݷQz'�h� q��H����hW}/ڶ��Q.��_\�bB�雸r4smb���e�U�{���)۩����SpôOc߄�K*u�l�fs[�6��8K�՘��E���M��bs�ח{�`N4�ގ�#	\��<eog{���>ȣL�ۗu�3vϹ��#�S��9?�w�E�]tkB���^��
��2پB�¤��`M��q�v�n����w����Dw���n&�>��r���Y�{]��4�_��OB��7����&UJ�kދC�n���~{I�c$�Kϼ�����@��]�B���U^N�}�9pZE���Q؈2d�d�,��9�_v�0>,j�c�L�㣃�N��2bi�r>��%U)���I��u5�E��LŽ���k��m���'�U�e����
#q�(o�;�ٞx䠪��ռ)����&��=��v�eUl����|ڥ-n�S���&�4ۉ�
qÈL�܃;�}�OF���΅Y�揲����j��tI�$ۇ E�.�%.��t����y���y��.��WKnYȩ�5��\�����ġ���`�����y��\�֜�-�e�x���Xi��n1p�"�=�gq�Y$�M�~�-tJ�?��yw�:��v�(T�~om[��*/qaK^�F���a�׉`���$U������i�+��{[j�j��qO.Ͻ~�@����xz=jnd��\��.&0�b�b���۳�C�Z��6�t��щ]���C��\ʪfv�^��8͍֝�ڐ2��R��;��k�Y��fͮ}��m���nE���0�v�ײf����^��Њ 䄢�R<��;m�ղ-�PLc����^����Ō)��헳��{�+M���WM)�������������� p���:Dl�Oo/c���Ժ���v���h^�
]�JUr�/��O�S���G����L��>���ݩ�����tX��.�}���Dn:Ӑ4ɽ��ͥ��1nd�Wt6�j�X{w�D��n�	&+xR�܃�=O�]+1�`<(UᒺN�p7�{Q��묛�w���2�"��
$7q�"��:�K���(ܮ�}�y��|^�QQV�+�fC$���z�ҹ�a4'Sӕ�8�����RB�A�����c/s����Þ�A��`�׋�<�U/n�3�8\�¡F	l6�9�����g}���=���oE��SH�����u����i��ݱ�H�f�j�B`�Dc n��(�{ٌ�����Ͻ�Qs>{'��%eT�}�v���8am`�	��Q1�9.2��r�Z�<t���{ي��_j6)饽��G�����˧�9X1��m����	�����b�z~m���7�֟D�:��reeȡ�ɞ�{vU։��g:�>ڋԯ��s����@�.�Ȣ�;ұ���w�twoq{Lj�M��b�n{s¼�e�a��#&5�D�H���j�a���{Xtau �y�Oj�P;�(��R�&du�v���C������d
gu(�faV[�n7h<��vIӼ�2I$�I#����	#�(*I�����P�T7C�q��Y�l�EV�u�ɷm0G������ZKfViY ��q�B]--RN�]���+��t�]�:���n�͗<�.��E<v����W�:v��g���KIl�ҙc�g#�83����shzN�pM�L<N�0����q�;�\Ft���CAۀ��;d�s�=�cf�V���`���=�%�9cQ�T\㔕ӬG7N"��r�bQk�-�n��]�+uu]s����e��~�]e˧&�f�1O+c8��Cq�=�L�+��P�za��sз�B��<��a�6�M!nGydm
s�~���Q�wFQ�.$4��J�ӋGb���pl9�{Wo^��4t��ai�q��|���;����ڵ�;��wu�3������ķP�:�����<�6J4ܑ�
��&V�}M  1;�w�\�>��{o�E6�s��3�qhVU���;���+�w{<�A�-�D�Y����v%�n2ݓ�/:O^���_C���[^Ֆ@��a�!����
b\�n��Z?:Ŀ��p�:�$�k�˴��SL�3]5Dm��*�b��h��
�n�ӹsf��3	D������)���}�,���츷pڇb'8ԍ�c��vܰ�|�1�҆4diɺ�[��b�NY����;�D�[n=�v��=r,4sq�NYY�+l��K�ɂ��=��@+t�[�ݚ�ƭ����e<{����qw\���Љ�[��y��Ua��ܓ5s�3g��1[X�n�j@�z�#i�ooEnf������僽�8�|^{q���m�<���P�}�[������GX��*���@���Ba���л�w�0�_(ݷ�[g�+�j�����p�|9�t�+5��ƚ'~�k\^�����?Sx�+�2G$�hԛ =��ȫ����c�t��3P�j�:b��]�{w����Ij>��Ț���>�p���zǤ��c=�m6h�f�LZ�e�`&xx��R�D7k�у��[����]��)�E�IU���nR�[�9��0^��k�3p츆���q^֪X@D�Ϭ��F�	l4�:S����Ｓ������Rn�YmFo`�s6������wj���k.���P%
�	����H(Ç����-Z��_.V���}Eg�vjB�Ͳ]ݐ����=�36��Vf�C�z�#��9]Q,���T'�c��=�5{YIc�o��c�[1u�#c��k�4�A�׮����8�Z�pd�ݻ	��R�es5>TJ�z�u&@��&
���]�q���2�%�];{!��VOnn�*��z�9�E�f�m*j��͡E����r��X�7Cu��؋�ȳ}����9D=<�#���%��9��/1s�Z�!Gl�ٯP�5!�AQ��9h�ے�Y�Ķ�g!Ӆ	�w�g�❠P\�˘�n��e�5��*Xu.Ff�2<{Y��2j]��2�5h:㼨�vgK��wt��:V-�V�Odٶ�/7�Bq�n�_\
�V�� �Vwl#hu�`���_hNf(5n�H�sY���Z����̥[L���w�F��sE�Z�]k��#q*��Wd��t�}��r�W� �N�/�c�G5Ĭ<!�n��Ǆ��I�>�R]��wVz̥��̚�:��݄e�RY��t�5���{D�<C^��*��3
� :��\%mf�BN��}��N�Ϸo:F;Ҕh�<�v��R�P۲��/q�����8p�q�$i_0�bO]�p��ME[#̒��7"��(�_\�� b�2�w&&/��ga,v�w�J�@�b� �%�4١�N�c�d�%�� ��i�γݝRP%ǻ��8o��)�N'ӝ�݉��)�0-�C�G.3�H[�ٶ������Vl�I��PHq��Q��,��r�c<&
�m+�!��2�w��v�����=�Sx;!��U]WI�s��;y�+F�ؽ�GE0�p���{��X�w���Ӽ���Ua��g�9�'8|�������Gp�ɽ�T��[���ȏSJ�0�M��7c$.I�t��9F{�c��}mZx�{j���v�7��j��烻M�Oz�-Ƒf���{�3������鉃�ޒ�Vz��ی��E"IHPƜ[V���.������,��5;����9�
ｖ�Y��,Z���6}�6�a�h�+F�h�[;^���nC~�f�fs���^�$�ys��{��udI����=�D�m#!0G!كfVz*>{�ާ{�1�,���]�X�,B�]��w����	���se��yV佣3��rX�9�r+x�%��9�,�����m�
Τ�Qzt���iEDˊ���S/s�}И���!��[� HD�Q�
q�xm�>�eg�ϻcc��^��zz��7V�f�=u֙��;-��]zF<��!��^�7���Kqϣ�C�����SJF-��GY�m�
c��뎋n�=I�g�7[�}c��i�L��O�ϟ����	�ڱG���{njۗ�Tl)�ٹ"���P�����W�R,��@�$a�pb��Ϸ����'��n�{ص�Y�3އ p=�xkK��kn)A@`�>�<^�
d%9"26䘥��ޏ:Mt�^�ePsݣ>�^!]uc���(�ݘ��|)4bq��p���G�3�B�׮��Uo��M��ݯt8=ȹk�/|�Sf��ﻺ�S3���v�L��ns�}<�.m;����a��F���_J��]��n5�;s U�g{�9�r���.E{8w��tޥ�w�r�g��qXvr	�/Y�4����L��Y�l�`�u�:�i�7 0B8u��Cљ;v�ԇ^7.K�Z�˓ks"��*.���ڪ8���[h��������v���JL�ݹ�gx�fY�t�eki��R��M�[��)	u��Ŏ��E�͔f!6���]!���ؕ����F�+l=f�^Hc�1����X�:sGc�f-���u�8�t�cv�D��!�V��M���sj��h�y)��#���;������G6�лFV�vNNG�Şn�-�l/5�5nu&x[�<��f��(ٹ���u׉�ԡ[=���]\i^ՠ�M��̃�*˱6*�������Mz���S:wEWMt��ݷL���"���z�\*�a����{�"xX2IA�����[ڱ�3{�c��c>!Q�}��Z=ղù�	���R�.��D�m���x��=�%�h��P8ڀ�D�����Gip�/�yؑt$�{��õ��t����c]�G)�{��7��cn��(D"���$V0飣`�w�+MK��Ҵ$�s�j��T�s���t� p^b�o��.f�8^���JH�d�S��ʏ������Y}�z.am���}ULG��۔�CXNEM:�^7��V�dV!�k�9e�c�H�lh��N�K��#�V� �.��׍�I���ؓm�k �8�mHF94c�)s���XEwa�늘��Gn!oM��2p*B'h޳�{��C�ACG���7	, �p�������9T�a��� M!�
���Q�I���ț����$�ww��[�-��`4VuzNi˳ع�3e@i�\`�0p�R�+�\����l��{�����V��.���\�5c�eoGh�&���4��Qǝ���,��辄a/7�5�:��;�qf�Y�#g)麅z+�v��B���II����'l{�x]Źw���aޅg��*�z�����E<w�Zd�f��[~}���uY/�h���i�\P)pV�w�n�	�L��v����=���<Y���MO�]s �▗r�y�5S^}���o�m�`X�r��f֗�-���)nq�ݞhÜ�����]͘m��`�j����AI �Ƕe\�g���g��V����e/=)ʅRsm#[�i����~���6a���^�&b0��.$q��Ϝ�����,E�NK����x�yTlw`٬2y��iͳw3�˧�tP��a>��p��'����h���P��=��ʇ.�����
�
I�G.�<��qz-�gQ������і3C����Gs�ma��}���倽�f�0ŀw��z��6k=��ȧ��ցaHxÍ97Խ��y��Q���{�1]0b�>�M�-����0�,{�m�=dd�<����Ѿ7��U��l�ԉ��4����Ѻ_3û.9�"gL�؞���k���\M�zi�����:n��b�V5��P;2�Vۊ�H�	<Om��Ý�].G��������m-�6�-.oMŷZ�4(!B$i��m��T7���3���J�M����g��7�{VX�3����Eo/��d(�$0��rE�+Jda{��܃��!�Gnh�ٚ��;������}��٫�Y!��=HW�.���7~�u=�x��:0D	A�T���ƍ�`W���t���8��t(��/W3���m9��O�OW���i�S)�0��(�eHvo�^1Bs��Ͻ��w<�=���S;�7��B� rxgOj;��sE�3�>� ��r�s��O{9԰�e��j(tc���\�b�5�n@��z+�a���ݤ����v`V=��`p�c�HKa��:�o��]]�U����4zﺺ*���r_3z��tS�WXn~u�q�I��qx�3��ϡTA���PPF�Gk�g-�F��-�퓪
ݱ�g�]�4=@ݮ�n��`��Z\B��g���}Ɇl�ǡ�%�ԡ]&u2�V�(��9��w���&�ӄ�S�v��Uߧ�,ǿK��0�ǩ���u9�k�2���]L{�-{Հ^o`\.�hK�҂&3��7�q)fi��{�qgg{�+��5��Y�c���w��y0X�aDǪg��2���#<ϒbC���E9�={�Cg���"ֲ�;4D�nVo�5�)�b{�hx�t���J���L�ȷ6�J��LyJʌD����C����k�W� i s�ol�<쮺Dy��,N�w���+���vW�n_oa�L��^^���xN�����ehʹR������`�[zc�4�cr����s�"s�=�ʝ�d�I$�H�AU1c�UUUUU[S�N8c��.]O��[���s<;���p<��z����J۞��!�6��x�z�\-��<G��:G{��^H������|��>:�`f�L8@������Gi���B�����vwXO=��"���A��ѱϺj֕���o^��T���ݛ���v��綮5�N�ʳrk�����|�c��\�J��v�stk���vv�����S�X��ke�
�痣=�%���.�K)�*R-��
҆!n���/��Yl�.Q7��]Ȗ��E�����|"����Z��s���NI��*�r"���aH�4F^�~��y[���QڿF����8����s�]�����A��/�E��T�'���!�E��ާsMg�n�މw�]=�j����hY!�vQ�m,��^u��}vF߫i����2'!S;V�=u�%V�MQA��+��=�ʐQ���և��^W`��J�}�d�]�T���&[.C�F䗏6���SF�;��fqM�d�v��po[4�� ��� �6��l���/ͫ���A�����.ݮ���[��#��(�Кi�k�5F��]K��/S��eo1Q�'._v�&4�*�To+�H��=��j{�j=3�^isygWgp�V��q��a�a�#�R8��㺝�����Y�]���{�S�`�."d;11V����Ρ�CP�,�y���[�d
��:9�|m�]Uu�yŽƹڢ���MvGE�hɜt[�Y����}�"�-��Ȼ�.�^�A2V��3׳�����z�<<��4\rE�`y�n����gr� �>�O�l9!\r�ul�T?�.	���E��Y�Ta"x1(�`�	�^cX���\��{�y��t��{(
�Ot_Mg�y����d��?=���	t�:�8;���l�AJ �i(�10�p^����n� �����%Ƚ�ZotuЃ;�]�_3��}��­af�C��jur/m(�MߔR����;�k�!�4�����ëkv��Z��*R��6`��]r�Q��~������5�7���uCȱ����������n >�E���bЇC۷yY[[�2cJC\�P�j����x#�}�U̇w�������F�k'�7���G�R�^T.;<�pf��l�ty��E6q��E�<<��;����{'i��x��;�����,��N�^���D_=�/#]�e[N	O�)��ӵh�u�l��E�奩6u<`��a��D�;�K�[2����V^��\�g*xa^�� �D�"ӳۆhQ�Z >��/�ݕ��J�����`�+����c�F����*���כl;>�~�8PL��@�dw}����~�J�/��h�VB_es�h�*,[��tL��8,��V�DU__���9q�s��Mt���';�d����	r�����XxKM�T8sv�ݑ7n˫s)S+�Y�}��.�ﺩ��p�|���ն�R�ݭ���}�,a�6���g�E���E	e�`ME!���Ѹ�{à=�n_��>������NQ��9�h��C���v��A�G8lD͌��x�Le�#Q�i�sLk�]׳���I�wy�x���X^{=C��O��)i�z�%v�� \�.H*e7bH��6a���<��_M���3����QhKbP"���{��<�V|�k�]5�۫E�:%�7�o�����i�U{m����c�{:��K���ڛ$Y��&h�=�/�w�~�XY��-�^�(�'���1v��W����;A�+N�7�{����t:&/�_�L=�!u;�#���}��|߼K�ޠ0Z�LL�J�����[6�v��#8��n���I�qÖ���t�(�NI��I=�m����ڕ�G��u6gP;�E�g��P�*���+����V-��r��p��@�JH�ayS���T3�z�}�
9G���)�����*8��(ݙE���68��yJ�]3��GС�(�#�ǀY���ǫpִ2��I����ݢD�_	4�8��E��}1�+��!���Q����-F�qIU`�2J�݀p���� �����Uj��us��F֪��@�����������������FqF�za�}�R{���Ei���#4��w���+z�
:�ëV�xw��S��]���d�;�f�������������m,���[���L�X�N;�v�0'�͘�%w�	�O�¦���k���}�%rQ7J�NI��(tmj�[Xbx�C�T㕧ii�&��m��2v���Q�[�V���ծ����"o�)��G��d������V�@mK�ٶ��9�+�t�1������u�zբp����]�l ��hV�PP�k��u�M'X�ݬꊝ�*Y0�,p=�7x�eb���M����������}�f叭7�z�,�d����C�xTH��@��r���n\���n�w�ͻ���g6_^�X����qL����D�ô�b�\ph7��D���aZ��Vq����y��S3G*pb�l�:�n����#6�r��qu�Q�	aB��c�ڃ*֍n�ml�D��u�r��{��N�FwBj�.ݬ���/J�Es`|֟x��˫j.��+��`��D�y3�ZkS�t&v.�4Z��%Ů8�W:���;QPTu_b�o�U�V�U�EDk�/I��1�b�Va7)�;�Rd95̔;�5���H�`��fw���{E��A֞d����:�խޅ]jY�\a6k&��wox�Ʀ�"fj%er*p�W�n�����U��w�����!�)�W۾��M��f�ڰ�4�c]�.�Nk��\{f.'YY��΢�f�T���,rt���*݌\�P#�����^\9��%a���M�r�Z�I$�I$�I$�I$�UUUUUUUUUU*�U��Z��	�+UUUUTUJ�K����'�[�1v:8V�������������UUUUUUUUUUUUUUUUuUR��,m�u���Y��_I�3��Y �O/���`9n��(���뭙�iz&�y�i���k���k��KJ6mK��c�	�c��f.}vc��qг�����d4f%��X���{6݀�r��鼗7Ro�{ʣ�u�<v���i�y�/wH��n�u��a��ap&D�8���p�{{t67'Cs�I+F�t"Ci��3KIS�(�5��l�$޷��'%�<�@��:y87F��8ϫ�V�6hGr�.�!,ɪ��7Gi�<kv�՛�y}��kX ���נ��Z�:��Ln!���+���S�XG`�]�{y�n��z�zu�-�k�Pz�Gm�L����nB��f��i-�v���k�2�%�ΰ�s�H�i�����b�5`�X؏,Һa���4`t12	&/4�箝mOm�B�3a4�z�vےdx�����`x'��z΅�m�	���؎�X���9�7jz��/`tb��u��^V�]�iX�1�(!iMH���\�Sc�J�=��"�����4c�n&�
���B��m�2�ո 7�G��D�{�sYRڑлd58P��q���.Al.9'v���Ξ���[�7�U��X��03>wdݸxtlm��e��%c f�C#6r��`����{�Ɠ�ù�� �p%9��8ɥCh�֕aqT
�b�2�i��K��]��i8��,sl�7[���m�ݯ��eϮ��s� �v�u���,b�ۢn��c:\S:� ^B *�F�����{u��r���������/��g�V��ث��{��I
i"hGkMs����xvh�=��3G[j1�z
4���8���&�k���v�؇v��y�l�0:2WmY�h� �v�:5�Yv�9@���gcE۞fU� y&�d�+1�<\�ںx�e�+�5�F��e5�С9s�;]Y.܅�"GWb�ֱj�����Z��tL;�UUUU[!�օ.�b�Kit&^�9+Zy�]v�n2�������su:�<�s�^�V�%�x�b�d��])���;�ك���WGY��ʮ#�;]3��.4��l�X@���5�-/],�[���l�Tk.��bE[��F�jB�.��2�ۖ$tԏ,��=[����.K>ޑ� ��bTu
�sm,�9�RF�:��q�
l;�^�h�Dۄ�t���c.��j��Q� ����p>c���䘕���_��w&ȓ�z���ɢ*6�z�*�o��9�,�(ʾY.���kB�Ti����JH�����RO�xC�l}�I΄�WoD����n�̠���(�!\.��ͺ_oB�:L���Tٓ
�
,ڐ֚����w����&�[^�����y	O�VW�H����B�6�?6|�f�a�E�30�0:eB������y�;�;��k�^�5���}��^��� ^�+��【`0G�_w�Om{K<��e�	��=�<��yIA���֯�dC޺򩑢6�������{��1�պ�l�A�km�^WK]��R��;�%���뒆�d���;4n�k��N��8�����*��}�mEꫠ��
0��F;��ܷ��G�[��x��$�41���^R��P�[y�M==.�^�E�ȼz#�R��3u��p:2�?���$��ۦ��o]$b�w6m^��q�H��8{XQ�Qr��S1���W��_��k8�]�gC��tf�
��;�L�%��D]�0 �aa4��#_i��,�'"�|�G���`��*�׼M��p?��_t;��o��oo%��2���~24�L�����k�8�Yc���3������]�MV�Eq���Λ]�r0wki��|w���5��G{^:�LĤQ�r-�{�4�Uʅ�ȹ�,����'K�sޞ�W�R�>a.���a~��׆���j����+M�E��9"Hܒ
���s��L8�;��0��5,s��Ђ6�[XD�N"aJ$8;����������Kئ͉��[��vU�=�r������͂0�"��[ɵp0��ܢ{^�Bq���������ڮ��K.^`}+���0�9��z@��~�j˼�l��{<��e�32�S�gH����L�&�}j��N�Wk���h-��Mw��x!�k�Ϸ*����mQAJ�惚3�Yٴ,�jK��8�p]�X'ʼ(����_+O��u�.��ݪx�A�<�**�b2q��1m]&{��)���A���B�Y/���3�L^���ܐ������:����vM+��1�lO0�n�«�ґ%"�̶�&6Cr7�)dI)��t��	���\uAT�q��޺�\s��&d������wQ��� ��I��7��U ��n�]f獛u�k��9�%%Ƙ�ڣ��]0�c.2<f�n��}�}�gh:{�
+>��E�;�n���{�;��ip���݈76c���+�/���1��}�F�{&�QV����`T����d�1^��6&���{��\�qt�W>��ѥ}����G-p�@4��"�XB6T�eÞ�R���,[�L)�=k���^�;3 �����
���;������݁�ft��Q���Bf�j�חg�z�����x>hQ�K��Z�A�{��ב�ˍ���z�O+ܚ�3E�Ϙ�Bt�f��*�s��\U���=Y��}sr_Q�7m�X��$��+3oort:�J�����
��y��d/BD
D̐$������#��\vX�YU�}�#�X�թ�0F��f��U��8B��G���f�=C6�m�Q'#P� �\��ш�c`��4��֤��{n[�#�hn�/\Ȓ `0)��i[ب��܋wm,$��#x�;�O{��2��O�n�= f����(�QNG�@�Xg4y�6������LV� Y��>�Քbp��w���#%"��T�X~��(qO0��]
�hde��-�M�g�/l��������^xCmm(�/*��E$�w4H)/z;R��mN�rډ�
�P���C�Z�ы��u]Z&z_N�Zu8�Ԫ70:7��Ȼ&zv�I홹Uv��m�)1�Tb ���d[H�#��� Iφ�P�#Ww4\�|+�����p�Ñ�^��ۥ���чn�/���i��G��oeAzH[��f��gOQ��}�B��\��qu��V��X�2��7W.�n��v~����UUA��96l骪���j�����˰�[�����Wc����Yc����RdaHm
f�k̈́�8�@���m��b�V ���v�ԇ�7�5��jԭ�����/z��V����/HM�!MU�!.#��F��%�M͞��CQ�`��,HǮp4S��3��i���״�\��3�b�\�r^�)��B�ZQ�m�Wqx���eN:�;�9�c��~'|�uG��pv�����p���m���yܮ^n���v�M��M�h�~�����~�R�%��ؖ'w�����3���)��/z�����w��˧{3�P�~�Q%-C$�)�h���yP�ޮ�g��x�\h�{�j-
٨��)<!D� ���ӿ?x^,w�t�Ǵ��в�%�Zf2LnIu���0�����Q�&v��rá�Tt�����f��L�v_�{5��}�ʹx50�u�(�D)$W��cK+��n�4��w=Y��t�͢O��ּ�����V1���cq���b�[�[M��C'
�G�ZS]ݘo������)�T����L��F���B���R����EN媈g����-���&Z�`:붊C=
�N2�9�!��Ay����`p�dj!������˾��}�����m��O/%������*�u�i{�w����J8��`\A��Gz���lw/Yw�&٧��ѓ
���?2it���d�uv(�Hk7
\};���;ju��!V{�%+Of���tnxoNԧ�H�A��j�v�Ѥ3/��a�{���3_Q=�C[e�P�U�V�f�Aw��+m�^���L�W5ݼ'��νWA�8�>�wF��tW�J�HC���REY�Լ]��+l���Z�R����{�<�o��jh�V�C��������@Yd��W$�b�`P�Z���Qe�dw+�t7ن*���7�����5V��3�kBw[}�-�}r�VE�]�̎��3�$f��(��^́W�pG+�v^w3t���6���V��ָ��z���F�����*��`afN�>�.S��V���N�EGu�ۺ��g|�yׯ����j�E��e/��G#�9;�gk��ȶ:y���}dc�i׬ɮ.^z���{�qֵJ�lbFu{��7ퟌ	A)��r�n�����EE�fro�y��
�q�v� ��j���wn��� ^[s/;f�@&�Ʀ�OR��|�c]p���"�iܹb�;-�e{�E�f�R�ղa�
�����m�4z&��l�(ܔ0Z��J���8(�|�f�r1�%ʵ��|��1dOgFdY��l=./��&�Q�:��/�F�|�N8�n��%���*���C�yS����+��"��ui���]VT��o�;\p��z�GI8�&xk�ۻ=�c^�$n�ݎ�n�K\;��S�8Ϟ���Աi[m��-)�&F����1�_Eԙ���c7�5t�ݏ��v/H�<��w�������':o;y<ru q�8�n�og\#���Zos����Abk�-72UK�H�{�}]�w��g��g{�_�Le$�S�"��C���cE_r���K첯�וo�G��|k3}�IFL!r�,���VkͲ�Ŵ��L �m�b���b����V�h�d�A��
���
�{N]w�VU��+n��I��)_��yq�63i�/�\�\����&���7%�gc�=�â�Q���۽���y�݀e�{F֖�Q�v�T�\v�Mfl��x�I�q@c��r;�{����e4y��;��n�6�����>۞��{}6s���yc�ۼGC��=^ ����j�F%�pɅk��6�����tnv8�7dv���L@����lK��'�/{�A������f�C��r׺�1X��m���<��Y�ޑ�eS#��O�"�MF�mG&]Wsršy��84��lG8��e���;#ON����;��3jH���lS�gr0+5e��,��&�C�b+��	Q�����E�yTu�dݯ�{ne�2;�1q���:�ܙޫ2j���\�f�`�:�t���p3 r����P�Q�3b"�zx*��I���K��'r����Qo*FM׷n�8�^<��҈t
7ՙo����MH�lD�J6��j��5�atQ|�g	�#�����X����|�x{"�"����8U3Y{[�
�*�-$�׊�È�D��hi��nv@��s;6g*����$�����>��A��UUUt \��K��������'����D�a�3�WF[=���ڑ���,�	M�/�@�	u��j��c.�tlk��2�hI�n�5.�\5Z��j�����v筊:�^8ϫ����T�����m�[o.r�6U:���݀U�1q8�b�5��w!Q�䕑у��v8�70�q���+����
�5�S�.C��
#�4�ie��%�M&�ŷR�ڑ�R��b[K˞�!ׄ;`6�[��^)Z�Y�7ie�`��7{�:�ž�^U���
z�b;�.�0.04nr�����f�t�a�z9Z8�''q�\��l��[�x�ח�%����y��:�k���)��N������V�w垒�+E���� R'!�Kܽ#��_q��קl+w^�PЪi��_-;&WUM��s]?q�����"�.ڔ:0��A�Ċq1#tE���u�C:�{�wa�>羙|��]Muܛk�2�	���M�[�ޜ�����kSp P dm�ci#[�V�T�A�&gn��ng�����Q���u���s����8��R��-%��|:bܠ�g��B)F��cu�����wI�����v�D�n|[I�<�qv�}P�������#�C�0��Y7���3�L���3�.-sT�s�'h�r�(���|�;�6�DcJ�
"I�u,ٸC>��:a���Y.ѷ�qj���:��W�y�5h�pj��hoG��Z�Z���P���]N�[�Ӌ�z �����q�e����>�Ό5*;�!���k���l��f�B��oe9��Ȼ	Z�L�$m£q�����)ݿ:j��d�-7���n�ݼ�1��Xp���t΃Z>�x��9~c.����En�<ˇ+k�ݯc�1xG�]v�˥WnU����(a�6��>����e�qvS�v<�Xm�*%����z��<��i�>�|=��oS&�G;���is��7��S�R|������#�~��m�]��,m����L�v(݋N\yݝ�����.+�zs��$&8B��!�ѳ���;�sEh"��+zT]Q̺)�\��F�i3�(�v��u�y��"���,0�� CrE�y��!oףe�`^���f��C��Tq϶��yz�o�w��;�v(y��T`��v��M����5���j���ϗ�����Q���� �U\�~��6/x�Z��ځ���F�����|DX����T	%��5�q�+~B��%���եSiPf�À]yj�-�%�j���]H��޺5պw��0�J�G������1��X����-^TĬh��F�����u��ξ�HI0���ۘ�4�]�w���B=�ٽ�b���X�{���X�K�@
��@�rZ�)�ܶ��A�:�>T�v�'e8����{���+ �u)+3W:����	b�^uJ�<��W؛6	I�'0X�{wq�G�5cx��n�tu�ܓ�w�{x��K..����Z�1�U@cpQ�qD��`6L[hͧ��ۛ&)�dH�P��)��,�|/@г쿋�w�j*�_��*��뎎�{׈�D�ƠJ{Ub��g[5+�E���V�	��[�$�h3����?��\P��=���3;��#�%�!��6�xqD�L5)m(�B��@��́6b��ɗ���w%Y<(���Z�2�\N��^ .$억"s���z���CU}i�mN���E�s.������jX���ЏT�e�wׂ��"��YGN]�w[�=ֺt�\ẩ	�e;���u�խc���v�e�����\�Jg*��ͻUB��@���\�X�� ��Z9p�$Y)��:5�oI[�f�6Z��F4�DV���=��LAYEp��j��,�����VG.�6��\l��ý��c(ۨ�\���������V���`�K�U��Ǆe�Q�N;����cҶ5�:9��*��Z��{&R���b{/7Ԏ^�&�������^�I��1� fD��4���̨C�8�]��ՑN���6�s�<>�[�؆���5WM<Mջ����'o�����V���姬B�s���uڻ>��F��q�"%A�W<���t�\�E8�0�ԑWr�v�
�w�K�Fc{�������3]�S8�jO)����h>"mnmy��a<�%W��HY�# ��)���(N����*�����G�4y�Ʃ_�����'�i;���9n��>�2�[��[.eOBX�!iGĜ����*0ҿc~��%�
��4�2�Y�"9�f�ܗla�C�wϩ�tFw]���p�Ð�T�f2L1T����8}4�ךȐ����W�\5�w/vtBc�@���7fԮ���aW#˨+��En@A��l��8!ol8F���o2Y��xն�O�����"�F�2n!^�ھ����k���(D�9	�	R+ek|����8])�	S̋ݺ�buW[�޹8��F�$lu\��i������!XN��c�-j�-D��+mm���!�s\�O`�t
���n��8��l�t��1q�%����_C,muM��p�;y'{���ޫ�U-�����\B���lb��}���#�@�rG���yS}�b������rݫev{��5��S�~�pN�4'2�]���$�r����e��"`��L�H�7����׏�T��?h�l �(f�ˢ/���������0�Gl����>�K.�VKK�ƃ��#NE���� zOHA*�{��L�]|<�,�m.ƼC��� ]y��k�:<lD4��<rH�M��n�eS	�}�Y.A,���!/칉�-��RՕ*F�{^��bek�X��)!>7���~�������V�$��k��앝����kd�=�&ۭ9�ة�,S�f�n=sq�N�:���[骪���U��n��UW�U|�g:[έ[�]e�b��6������{k7f�n�n�񫝗��t��hh�;j�H�[���r�nx�#���N������fǧ�p��aE�n�s�	s�l�Z�۷:�vQq[��p޺h���рiI�"՚��yvt۝*7=�ڐ§k�ttZ[�u����G��98f�ō���O���K����4K�M����C�wg-�>���%�6zw]�x���N��8�b&k���	�u�����F����1�Ͻ�!j���_p%w��������o��.�	�q@T��z1����'�ta��&�8.��7W���{�����b������r�������lL{32�><�)��f�*�4�颱�i��ȼ��r��7�޳�^�LKLt�=[����5�R��Гp������ۺK�p��Y������د����r��g� ��bta�5�!|X�A��E��6�i��oƲ�R�MY�z���{5hO�xg%Ay��]ze�[UӺ9���� p���R���c/k��f��j:K�<��lu���t�x�k9���[��m,�8bnRlQ��6n�������.~ظ�H��]{e���^�ff�j�.̙u��1���_E� ��wc,�i�"݀���}5�G�d�ꋆ*LP��$�
�am�gX8�˪A�u�sn9��TJ5��C��>ԽKNe�07���oׅgm=���y�tӷ�5;��;�N�zv۽�tIݾ��ױ&s_IvyoQYƆ�#�y�D崃r4����NڏMm���>vAƧ��Y��9�.��l��U)^���yx��m�����&
qwwK���^8*��+�}Y�b�t��5M��[��<nl�񻵇���8���eЮ?X>e�8�(�d&$�7�gW]JwUR3/W�'��*��
ɱ/;�Dơ�<d��]E}��=�j�`����𧒣l�v��v8���rd�{q�.u�i����r��z�5�p=<����[jJ���Pn�i���F�{]�1z�S���h󶵡B���������jp�JQ�2��Df����ɴ8R1�ƭ�k8O.���E�c2j�:�>���'��%�h
� ����>e�Ei�UX��Yy��f)�LoO9O%�+���Π^������V��Ķ]?����n��&�ۣ܂4�ٳ��_]k�q,"��ѣ����s�VY�;��{�ۘ��{����w{�+1�6�e�;~�]�N�iMq���xS%w�ˇ՜�ɐn�P�j�gt�]�
��xr�k֫���n��/#��^L"��MfF��6�cN3zm��ӣ��&j*plw9��״�׃Ǐ��fr�z�;C͵�-Լ�GrLHdn*M��!\n�����g���;�՘utX휠�ݭ�-w�a�3���{c�^�蜺����Z:�.�mŒ$�d!3/�j�զW	�)���@d*(�V���/� ]���V��ƈw\T0��fW�eG���4�+�\*(V�@���q{%B!9��w7+v�n�d�������3{[dx���<�쾹r�i���紷�/vOf_��ɰ�|o�S�-�i�;���s�u7�ו�m��&3���^��%<���j���%v�}]�U��7d!�wp���e��L�,C�#�ԫ������
�hL֋$cYEl��f�x����;I{����9�=�s��@NmA�,W�
ۀ��m���V�U��7���I���������
�7�Sn|G�����o"+��@%^m�)J��WMb7 te�Um�W��z��@v(���\8�3ä�pvA�WT�D�f�?[�����?T8j
HR�ޙ<�cb9�n�#8��8��sٱ=��c�aH������4�9a���o��|h��9�&o{.��Ut�nR��,~	��v�sW�ݬ<�sa��G�+i7��-�L�J�ȭ��\[��VՔ��ں�w��(�}�wi�Z�8>*��ѿOPuɘG�+A�<ЂA )�(S�����݇�f�T�EC�=���{}�4�^����-�ǂv%��;o}�l+]N�f���eed�("�n"�rn8�� e��x�v��ۺ�ӖҮ��[\��|*ό��@kgT;����<�����y���Kx�s�t�x�f�h���*���4l��'K�p�����,�R�i\�Y��Vf�2�;]��$�I$r6qIBqj�����ێ���x�p^���o%˻^ױ2���غ۞��2kv�ٝb�v��$b�쌍�jqlf�c���GX�t�]�y��+㡏,�鍸M�n�S�qe�d����#�y�z���I� r]�nbAa��4�v�6��
����)v��mN��
O`p�y�F2��N��3N����lv��Du��j��.��s�S���щ�r����*��3�� c��s���_l)e�����E�H�lhմ�|:�;}�+��"Г�����!�q��oQ�i+5�&��B�ҝ�-���b)m8�LFJqn;9�����ʟY`c�Š�;ȯgwR��c����f��,��[�����E��o#A�m
����l�o�{���Ž�KQ���z�%�dޞ��Z&8�{\������/�(N4#p6�q��[��3�f�g{$�x���ܡW��p�1�M���-����V:�eq��k��� ��2����!,���x�=W����Q0�6����*�{S�ٷή]e��La�uK�V:����Hd��w%ur:�܀��k.&f6�]�F�#��%՝B^F[ev���-6�q��߬��;�u�GL��ŢR�s�DN\�8�nãs�ĺ�{����WW�U��e&arCߺE5�^��/ü]6��Q虈�^��Fl�u,|z^�j�#�}�C�*.g;��\t\���a�+(�T]%�n�Q�^����xL5}���:�� ��j�X�^�[�V������q�`�$1���`r����pg�9}[��RCI�_FR��������v�r|�*���Fu�\m�}aQQP�Ɏ1!-�ks�YӇU{����}Y���y�{	fDS]��&�.�MsG6��T��9�Yu�b�L�_�\)�@˕�y�vr�F*뫈�S(j]Q����^��֡��Aw�1�CS{ҏp�={\o�Ա��U[1t����Z.���b��ܶ�voG�hք�!�c����mL��Q�uѱOz�3�6���P��d������F����)��AB�]fF;���
$��.8�~�X�O{~4�� Vw�G�[��Ԙ�̏��C}�;sDm7��"r@��fm��O�v��RIG)�в����{Ӿ4=�|�����F�����ž��l�eQ�!ވ�鏳���;�{Fm!{�k���Cj`��B���K^N�y��Ѐ�e�)��g1"����w1�Rk����v][�ނ�)"2$E�����K/m�WџE�wU��zk"qG�k��-ڕ3y�,��ۖv�iUK<����䐧!�z>��+�*����^�C�{��-��>h��ά]#u�7����||�1jҋtR��"�n���qX��1X8㋢�f*wF�,;�X�ÑB�$�"I�'��}{ٛ�d�6��=}�'��~2�V-����k½1-�{���=^�}"(R����+0J��MǓ�v���Xp7A��8ߏ2�߲��qw4#�o�ʰ���.i	1}֙)5*B[;y=o��������l;}�z�������н�3������}������4=p�	���ou�A�L��}}EN�n�j~z}�t��^�E�7����ǔwf�'=�^~ ������-�WU�U|r�;�	8IR: �d����ތٙ�gCEf�����6J�7
���Tz��#X���u�/�"`h�0\,��,��ݕ�t}��;�]��E"��>y���u�齍c^�1��6�y-��V� ��~6��>�p�]�ǔ�����6�&g'u@sd۞YA�F�,k��,��m��Zp���X�Y�fã�v:�0�y�����MY�w*c
^z@�f4���#�y��j]Oҥ|7��*r��;�9'N�53S�ǫVֲ"����O�c݌¡B�����B%�=��;��Wnj�Y��@]" KA.�_��s:�ek���y�=�m�� ��<pƤrN��3%���On�ٓS�Ǭȹ����U��Ok��Y��޻~ȩ,p�d&8À�!�v���Aމ�G�9��n����x�ꖻ܊�+^�s�����>����y�U��M�b{�7j -5�f>���������דVT[/���d�xt�{���};A��(�76uKr8�n;wx��}.H71�M��`'Jޖ��cl�I�t1�V�9�c�\�����ų0*�3�͹���>�j�L�.�/w&[��=7F��p�Mb.ᒸ�f5�{��^@R�[n��t�r��t�B�PZ{QMјltB���)�l���sM��G����o�`��M�8�;���h��6qp����'o�\����o�I�4�3��YW{�f⡺�۷M�+�a�[�8V��ڔf�Sd�ۢ����	]Y#���Ϭv�s�S�^u��[P�����\���wj�G/i�΍��15���-��ˠ��ɛ�e��ʺ���V�G$Rk����z����oV���i��㭅��1��:�h��\���b�Y��w�Ԃ�.W�A�ޙ"��,5};��#J�}�^�l����\�VZ��f�B�C�o0�Db]��u�Ֆ�
sBO�Z���lWR��6�u�E�H+�!/�Z,wU�[iU`�_r���g�t�Α��0@�M=��dH�ҳL��m�l�[@�[ϖ�t�%V�����.��+V��1�j��5A*�����&l�ʜ%\v{�o
x8�V�dI�E�݀�6*�Y2v�&gq�j�<���c-昢ݙ����"�2mZ���nL�ꬼ5��Ѽ����I$�I$�I$�������������v�#%*��@�UUUUV�*ʉ�ٕ�.�J��ة�0�UUUUUUUUUUUUUUUUUUUUUUUUUUUWUU*�\v���L����j���չ�+�5��v�In����s�޸����K�X�
�Ɣ��34��|�u�'��]�E^�\�J\c'Z��x�k��I�8��h�t{M��#Wl��8�$�)�8�\r�[q�kh�w!j�[qj6)�ە;lg%ӓr9۩Ӯ5)�q�YP��#ucѺ�n-��5��\ˎra�᱘�^d��54�l���h�}2Ntsq�i��x�]!i��p��]����H�=\�9�؀��vq�u��yC͡��x�i���nڎ�v.r�nŝb��ӐK����1����e]�JV`ukd�0\��<���5��Ӱf+�g�I�l���V�a���J��q��8�dmY�a�v�G.d������yq���l�L�d���X��w[�n�)��C��+�.]�m�z�J�xާY�M{v�p���ϝ��ێ�˲�����-����\Rdone.Egs�a�kpn���˫�y�\�u�ɱ���ae���󸶦�I�:�9.�\�Ncb����.�e��t9uΠ�AY�����ۄR����e�9x��랍Hk���M���ͬb�� h�b#�b��q�U�';��݇ڛ��gi�;x��]t�۶�q���ĜP�;���鵹9�����&�8xqg�c���vop�jN]�7�����6Ҧh�hu{v���a�ی�=y�x�X�Lc��F����'8�.�<��h&�Mm��On�ό��C���ױ��M ���pe���(I�R�	v1n�2�	H�iH&�s�i��7�������nr�b�,�vy�s�b��v�p���r���ʸ61���Хu:��U�Vmfa]5&1�q#�����ݗ�g�y���n�,�Rsi�P.��7������l���l;UUU]UU�Fj����C��0=����qp���RhW�ٸ��eƩ�nَ�K����a	�t��q�@l4h���ͮ�L.� ��װ�Vf��*5#���jn���#����f���H
�q���֧��^"���r������;Y��l�����n2�����㱜F���v T2��Bz��V{����r�eݞ����T�뭵*����	��929yCGF�;��܋�ձq#9�[ V���:˞<7)��a��7�ǂ�)���=�k(���i�S��ۯy�&��D���21�َK��z��eͺ���[�F��ؤ��q��,=�t#�,X�0_�nևܱ�+�k0$I��1�}��,g��n�~n-����P~��+��G�6�=�H���ڏ\�'��A�IH�n,2��>$�Պ�3�v�W{q�
a�b�x=n�Sއ//�;xN�V���T#�H�0D��y��ͩ� tx�t����Gj��vfj־��۝�5���|&����6W;|���$��y6�)?�)R|-���}%��]k&K�$��\U�CF�E�`	!���)��)�0��J�V{|����$3�줎��~;��]��fa�B�Y���2�>�L�0�b������b����cV��e�9���qW-[�h�llM÷L�%���\%B��t�L��v�c�)� �}���Z�W�QJzc��r�z`���u�n	�v6z��q�z~q{�ItҾ��-q����%K��$Jm ,���l�`�������v{Q��37���_ǽ~=9v������hj,�jw��@0c.2"�5ز�t�;%�V>�)�����\���(�)z�����GX�M��K��5�����?8V��8R�W�����̓��u�5��'�����ke���y7�k�ŇdͶXF��?V��k��L7e�#i���Ԥ���Fj&َ��L�ۏH�[[�.����0�A��[L�7��G	�;U{�.R�[�jOt��a�g�6�t>��1����Gsr�}�"N�nĊ0amś2��o<Æ���,�N�\�ƌ ���[���Xb��}��Z&.�����r@�B4���"�u{~3.W���v��+ûT3��k7ԕ@E�vGh'QH!�*�P���35��.��4�tI���#��:�,�fa�}�қ��Vrj��4D���oN�v�ב��T��Z5��IxdA�"n�G�.)W�s�$�0z+����܊� mgyE�(rd�*�C�]���tC:���a��C&�M�G�ko�ߋtM���
T^z�(�Sz����rT���;؛�@�{��܁Ղ�a^�x獪����דr���ۢ��ٹ.�'�]*IaHȎ#����"��q�q����p��nD�F{�q|���w�F�nxͰE�u��%D&$'d}c3v��!����x���U�]GKc����}�<�a{�4�^�x�ќe��b�,�P��6p"�I�a���"��]wӓ:D���o��%��:L�6������l�L��6m�e1�|��H����$�u^�Jؙ�Ȍ�Uܻ��7��r��3�^�M�tF]�&2P"�A���w���sk3c悚B��U���-�Dl��g
���ѥ�̌\[�v{x����y�ﵔᑄYS�ڹ�}�On��X$�	$T�����^�Vɡ��ܦjb��p�</b7�X��~&����S���=o~��|���>{P��Rѷ(�iiXT�:n�,[������5�y�����ʒx����l ��H�bCE��OF[��<��x�ϖ����϶���N͌ݤ�_�F�.�3�iz[�r�V��P:e�AQ!M��ye�^��-������/�z��r��m�_�׽�3)Qm:��X%�����@Bj&�rf�t���}��c�l�����ؑ�=�Q��~��T�g�X���$���n<�n�����]�vdW΁�3��k�w�	�}���_�N,�\�Y�z�w�"��"HR2�Aޞ��E�8g:Um]���#��,�f槗���[}8�Kc�F�]ʴ2�mo���}\�Ղ�����ޗ`���'/�j=���W���wľ�ia�ʇ�0')�2�@�˶���׀*n��KUUUUT�v-�F��֭��9wfɠ-ْ����u�RQ0JpF�YxٯA�$J��%�6�,�2�5 �,����n�r�j�E���P��^; �Nq�g6Ś��!.����F�AKq7<v�꺍k�=F���8�������C��u��"���Ϝ2��D��2[D���wn4O�a1vx��r7N�!f�v��@�C�.ܭ-ډ2S!!n�:��-u�<S�lIfPp�\LH�M��Dq���U�μ���v)�2hy��B�o����7�P�{dt�_��Ow=�f�Ԍ��Pf��/�ȁ^>�P.����u�=�C��tY�am�U�[��~�.81�G�M�Z��l�M@�0a����]}�R���l�{�%E��U-�.��z�{*��ܯ<.�"��
=E$E��j��HhƢ�z�:W/'Uzg���;��K=�ץᨽλ&�����e�Yl�Z�$�Î��g�J�ޕY���}3��x���M����}���n��x�w�p�����w�5��HZc��z0qź����F��<!u�ll!z�Ri5���KŹ��(����o�K�b�e�c�H���?s[�;�e�w'R�ϝ'��#ޑŋ��*�Q�d"I#�{ܧ�1g}�F�_I�y�f���7��Z�b��7-Wx��{��ڱ�z7�P��m�Z/w���/[� ��n<���@o��Z}�vc/2{}�_Ow���{��O��s�ezR��ަQa�CoK�76�����-`.�3f��|����s1�ZV�������L�o�}��Ct��V4�,ҭ�S
"#�{+= <'�x*��^��T��G�=�����=W37ӚkMvƋ\�9E�*�RI���㎳�Գs�{�_[xU�Kj��_�۵K����<X������]��m�+V�c\����PY2fDK�1�M��aR7G��&W�o"1�q��-u&֛�3io5Ѭ]�-���O�ߏ���{�(WIV�GwE��+/Cm�S�<3���{�8SbB�m9���e��_{#T���;��7�b[�1��鼹Oc�q5w��ݻ���C�Sm��}��8�&;%Ch�n
̿L:��~�̎�2��{�,ޠ)��^�\�NeK5��Yt�ϣ�	n�3j[}�f�����X���W��Zjݱ��F����F�ޮ��/ʐȪ����jg6u �6�K1�M�$�W���_re/o9-�;p�U�{}�.�=�I�����:v��@�x�ِ�`ES!��K-�UW���rߚ��I��	�s����uB	�梷{&ҩ�W����qͥ��i�ޕ��ּc�^��x�����ބ� r@B; ��:�|{r|ֳڍ�z�]�Q9�ٺv��cZ����Et�2�WF�v��u1}T�7%$H{�9|�j9��()���u��Bm��Hۏz���Ľu7�Ch����:+,���l��w���uZ53�����=����G�)�*"6�G�a�P�}�+3uJ]�O�f
69��W��)0�r��m�@o;�h8���3<!>�2H�2##r-Uӓ]	�R5l�l>ѵ6�����2*��tc�{O��
�pS�'y�I��/v6�,K7�VS�2�ٙv�Xֱj�8�!�*��]���@Z�;�"�q$�>әZӭ��>�L�qޚ�Ǩ��ZZy���[c�.$Q�k�*:��;]��헃�"���T�E��w�ڬP4KZ��p�$F��.F���H�LWp��i���0�'']=/E�M�&s ��28b�wZ�mw��f�c=<��:����jv��At=�W\8��;��������1��y��m��L��Z3ZQ��1b!�#`'��棷N�Fw	���vRM�-�ڮɫ!&�v3��/vQ��CNI~޼�ds/��J��\çlw�kX=�u��L�Ӄ���M���3�P>�©s�+2��T$�
NC�u�z�kǻAN��*�5���	��<��n#igl6���B����W��)�k���;mx��f�37.ń�޹��w��m��VYk�,���a�=�e?��<9^m�0t��j� LuIu�*`!�Ы�G��������H.G�����8�݊�%+o�y|e�P^
5������Ul0�.�$�I#�(�rE&�c˚�j���������K�y�q��\@q9�9�l������� ��e�x��^ݞ�<9�뗇��b��l���
��1�^(<'y��ڋ)�����-T�̠S0 �7x�2�,ۂ����=�<T�����q�u\y�
0E�8�ֶς��GTm֝Ÿz�q�.:�/ey\��v͓�U4q�v����F�ܨp��ݺq��*�Q�t��&]�� �[�c��ݛv|�ugX��9���
F���'��\g��r�EC��{ŏb�z,E(�QR~f�#F7�SҲ&�a��|<oe����z��y՜�$�@�֕���r����W��Iæ��OM��"y�aԕ�����4�M��m�YT�o|�Z8�#]�����x��q�7V�G9���rm�WV/����T�ф�����\�6���uj�k�2i�����)�����&S���v�����sD�����J�\�o16�"�I8�e�/2���7O��1#�~WCL w�W=�����\z��?{]f���Y��R�	þ�Y�9�6$a�Ck��s0���.	�:<N&Ӻ7e{��/gn��#HN(��p�[��]L���Nk��[r��l^�7=�xձ���C���8�U��V/o4C�$�2T��A*$�X,�E��:+z�p�D@���m�Z{]�����#��o���Q�^�d��y}��*.�5�^wa��ٝ��=��T��_sBt�Q�vO8��ֽ,D�W '��y=�\{�v�ϵ~�o_!�mj�4FCEn�Э���~R��k��9w�C������brG�|o��u/��Qt�1���E��M��aH�uw����kj�$�c�(r�۞6f�,Y}د�=v/z��P#�mK�!
��K�%�0�k�)�?�y�|�0'�8��ȰoR4���� ���Y��ݨQJu��}(P�w45(С��q�����/�|�"��DJ�l�����i#���Q�W����#�j������qRtm���,v�,,u+�u�P!k��t�{1���P���'�#�k�/�҆��� �C���M˲A�$�d���y103TTwj�:8���4B�ޗDa��SX�;"5���2Q�FÂAC����dY^���wqx����<~�U#Ʃ'�,1͝:D�(�w^Lr�"�jF�|�7����'�������f���|m��	�2(䱀��VC=�B��z��1X��0!����<X�3� ���ωkD{���g�*ѐ�M�^����kr!���]�w��\�)�a�^��/�2,�s,�#S�.�hH�4�T�xf$��l�z7(K���xw1�����������.���v�s�MD]s�owY�k����\�\s+/�-s��n)��Vس٠��r���'h�eۜ��t$d�D�� ]����j�F��h�SN������S�X�3_D%d�J啚��n�����Wh�c.Ѐ(�釗+3Y�۫�z	�0��08\�۽�R��Vc����c�ű3Ω�w,�yܘ��I��M�]"��tq��#�T5f�͡�)V(�և�d��j��QeԢJ�ݷ���Ɗ
�_aw{ m
]��P�����Q
C�ຆL�!!�9ܣ|��������j��wa]W9)�ff����
�O9g�ۆ�2!ϹS�J��ݣy�V�md�_�l���T�7ޥ܍,�W�����
w{�:XǺ�d�9[�76��{;YT��Y!c�;�U��=y,�����s����,⛛�e��{\)�⨙h��&��&Ң=7I��)X{n]��)�FSzq��;�M��6��S�#@}\�#Sa4���{��;�:��oETں*A��qH�A�,a��?]�V��(��#C����a��g3c#���8jl9�^sUR^6��guncύ^��v�kK{���*��2�e�n��������-7�1�8ӵٹq�A��,?"���P����z:Fi������E��8YPC19%8E�s��$38(���wZ�q���!E�%����x��J���@�z}/�"OjB�}vp=��;q�9����>OH��>؊ZK/�؀�JnC\�K�̑�Q=V/�d�܋ ����s��q>��.�g�J�θ*},,CA�4�4Go���:B������c����ߟ��0ա�n��k<�>�9��k�ZuΒ�G���I���Yٷ���v^����&�8�4���CǊ����ҹ��Yk�̈́p�G�}Ɋ������H{�^,D�g���M���Ʊ}���5k��<��B�L%�i�$��:{K0�:E��K���_`��c|X��f�}���mrcL�P`�<D��ݿ*Qx��,�fȿ�ϥB;�'o-�"�m��;Ό^8a=��-���CF8�qU��	�0��ެ�gJ%���}��Z�>���<pI���p�ڗ�qr��G9#gy(Y���K��#c2!�au�ĭ�@�-��qŜ�y>ڬ_ml�t���=hx�ܥC��7h?Qщ�{=5�KP ��e.#����֯���U�ֹ٨s虹���}���e�G6��k���ma&�9�GfK���[FK�'M�y�'�R��NM[�!�ݳ\�6�����g�6�"�&6�0Hhf���i�!����;�u=\`�Z[��Ow���,>�A�f<�&>yi�v�jeL"G�>�~�l<Y2En;!`���4�����drHl��0���K�9ǆ��1jK�T1�4b\٬.`��E��US\&�Dp���w�)Q�L�H"vo��a��/�l�ޭ�z4�G��di�n�B<w�F/���`��������'��rB���9š%�m9,i�� o�g�Xå�p��h��Yݹbf�H�W�����z�]�Z�tY����+�*�������#O�Ix��+�%�� �ᯈԅ-�,�>��acNj����o�*u9诧U�(������3�P�e��z����;¯�k�L|F�a�����o��i2q�$h1�K�x�C���ֈ�2}}�:�Ҭ�d�,Rg�/Ɉ�dQ|d�.�X@�t�"�Z����x��ߩȼB��~��/>�Њ�H�,9N7"��>����e���}�����(����)=Ϣ�=�<����g��R�5aq���1#W�t�
�"�U��Mo��B����ˇQsii�f�G�Y���ӣ^��yq!u��p�˛F��H:i_gffF�K�U�'rR�[�-<�yPe`[�f�ZtsW{$�I$��m)$&���*�UV�tm�n[�ұ�ٜ��0M��H��2E�rU�k�2�[�+
j3LM�������\B�no\�sx�ϫ9C�0��f�-�LD�+��X6]\�}�2z�9�n���#�����Oq�c�HGc� �`Sn u�Y�M��SL[J�Ҳ��(0�^XBiv�qf��S�8$rH�c.y��Q�7;�[{R�i1@,ݔ��=���:51	f(�f�s4u�y5��B��4��v��\���vO������A"�9��!��dY�`����6{��G��>ۆ6���s:��YdQ�:����n�0��Ih#dKc�"�S@̂9��w�|�4�^��Ɠ|j�:�t���͐��^�\t
#�6����Aj��Aj���YvG� q�)CF����G亞��	F>#
0�p���]U-?��,Q�}�"���ސm,Zw׻,G-"�w��pT���x�X#ò�1q⌘�%�G莿�X��#O!�c�"�_q� ƣ�|��p_�~��D�9I
�g~\��V'"H�w���Ci#GH��P�X�t|�`a-�����U�zF��}��Y��3���L)J�`�.�/��A��}m_�c��l�7�D?z�-��t;GG<L@���k���P��,`6Bi��{�'��^&8��8�Di[�ߠym��֓Y�u��[��6B��G����N��Xe5e�gb�ZP�h	%DL����"B>�'Gޡ�X�b�D3*�"��C��dq�(�E7�KՆ�������4�:G�w_�a8L�es�Q��6�cEAP����C(�7��Ys����T�d(]U0\�t��h��}2F�8�Za]�(�u&���ٷv�f�n���kl�]�[���35XvB�kkB�(��g�D��������S��{ӔX���(�4����#�,�8F�=�&T]�AAi@�F|��LE$�i�#��ҾXy��"�N�j��23��<:�������LbPTN/^Q��g{u11p,�0�6Q������a}���__ z�#LA�P�⯏��HӚ�W�Tʯ,��!y����VX"}��?e�u8�R�H��&���"��D�E�6ff��o�]<I�D��#+�UAB�F�M�d����h�~<�v����7�0j�*�m����nv|��\�~,���8-�1����D�f�����#���Δl�>��^�����Ar@��]��b:��u��|�>|c�L�:(�n�#���q��,�yQ�b��߯���4GőD:���\�]���7�^�W��XӦ�ߐ}z��`�F7����KCA�b��6��v����>��HZe9+���G��a��g�*��d��J
�G�B6������i��2�>��Y��#谆��7��R�1��+������:I~����đ,�e�,Y������S��çƏǓ4d�U�C������NК�w��cϤ��u�B�Xù7WikVX��Xޝj�{5�WM[[���>t��vۺa�n�$Jg'�g,�}���,����cX^"�#�i���~��Ɵ��"����������I(!&8k�N�������^̗C��`���.�C#�y���C�t�."����p�f��:���.��U�C�بn�2��i��,���))H����#ǻ�i�~]�_74D7�ƛA�YQ�n'Ɉ���x���Ń�M�2�z���La��B���42��W��~���7%%���`J*�駮��ϵ˟l=xz�N���"�10��{j�r �r>�H��b���}�;�ӣ�a�}e�躏C���{���T0_�q�� �1T�ǟ|��H${��_�W=�=��5�3�>pÑ6��LD�4��d-X�&;պk�3}u2{����!�7 Fȭ�Tt������C�H�^"!G�?GUq\~���*} �����#+ݱ��	8��� fI#�:F{#0��,��خ��Vթ#j.�ab�����cJ�(�U컏r�*�H��S�X�K��0��	�Vx�ICH�����]��,�$�
1pޜ!��ª�+25�!�{����Շ	#ٛ~T-"��G��*�Ǔ���O�
�{ܧG5�X��:覲��Y�N�'>ޤ�#�Z\V�v�?(�k��V_D��-*3*桓��{�[N�ػ����ζ\��/�z�/�������&�-]������{��?=�,i��㇍��[^��cf��A��ܑK�����4�W�Bu�C?-=#�\D���0�z5"�"�}.+td�cXa��}h)R�8E�v�v����,����n�pD��_GH���g��'}��iK��(���,z��jΟ�P�mzX5���x̢4��i�c+Oזޞ6�(���x$~E���`0��"C�H�df�(���"�
za]z�@�x�_Q��9�p����`Ѫw"|�d]�|�vQ"��p������E}���r��ǧ~��8D�a�В�!A	BQB�
5(aDC�>���ɟ��Q�;\dE +��'}/�������!�^���KI��J����-4�&�C!�/�F8K�GsK���g:~�[ٝ1^aV�0�^�b��<C��3�ח� ����֗���f���O@$ ���I뺗a\i:��PC.³����CL�1�#
$�9���#�#;׾40�^4d��(ק�����p;Z�z��q���!��a�,�4��~���G�hv!Br0�Q�>���S�O�����7�W,ٹt������G��N��B���B;w�ΙP�Ă5��wފR%q�p�sr����ud�IT���;EȵUUUUZ�q;���dYڹ�D�M�T�I�)�6�
��aB&���ݩ7hq�,�Zz��l�ƞ��hNlI��4����1�G�{:wrNz��u�;���]�C8y9�i�vI�16ZZlZ�\�D%�+m�7 �����X6�R�R��*�,p`%��B��z���[��L����m�,t����c�3���b3���`&8ԙ [��ӄv���v,�&4)�1,ѳp��^vd0x+�� ��̡�@>u�7.g����x����ړd-^��&/��Dg/��U}^���$��Hg�E{Ɉ��:�bY�d�0N�$Oվ5�oR>�p�G�<̀��7m0	�0�a1�)�s�q�^:Gg�:�V���ݔ���x��d���,`?20��hG;�'���Lt��>(���n���b�}�2�)>/�q�/2,�H��bF 1��)�\����0��ϓ~dY��:�/���X,ؿr�<�j��?Q�]>��4�Þ���~���4�r�	mϞC�X��g+pk����.<����g�93G�_�~f���?zX�ԅhq��з�Y�ܻT;����6��Y���Bؒ ��c���g�ع�4Æ�Ǹhid�#%!x��a�[�>�_�Yk�Y������8�(a�C��<�C���G_��=�U��JP�}�X���i�ok��n���+x��J����)X3M*ͳ�����HsA�͌[����������xu����uQ���4�7�&"6,�<}���<��b�I�D�da�Ⱥ_*�t\"���'�ID
��E$@��2'�:^�<K�C�U�mW��[#A�뚪�Q��$Ŏk#va���%ډ���:}�ig��b_�G�x��#�vI@J�f�"_`�ԁۛ��G��¼,��|���}����c�Ax�1hLz�X�dYF,�W�/�GH�\��93\��2�b�����.r���}��#T� ��Vx�իaQ�g���,M���Z�M����y�؞����,�uG���*���W7ٰB����������m�Y��S&��5����!��o�#���/����g���]w�T�~��.)��Pz���"[��vd"}7���"�����ı�	B�L88>��Y�ƅ�/�|�9��-B�ί{�/A]���?3ğ����Ǔ�<�F������C~~�B��y�x�Cŉ�o�����?�����pW�N�1�b�õ�v�m� [1Y�`����Zw>D��V���a�G�b�p���v~t<GM�o��0��k|]���#q��]���7骯	����x���!;����)?a�DX>}�;�N�7$�&_$����#N5��>�Y���;4W��3>d#����3�.�x1����x�X����ǥi~��g��0��h�w�(�(,�x�(��$��!�q����7�>�7WM�Gށ�n����?2�zFȣ��?�d�?~�(+��a�jk(�J�� �֩�̱��q�6���9� Ħ�[`��h���ngY8����B"����z��Z��0�G̋>!�<��W�i��,�8��6ֆ��n�L)�Xt�)!Ȟ���s�����>�r���b� �������c�Da����~,i�`�:zDz>�mw=�u�-"ʄ0�	y�+�I)J��)�H�:{�,�_��:r����8R%�\ODm�_�ᯟ��HgǏ��d}hL#������	��6t����Ŀ�{�f�m��$X.Lp��1��v��U5mf���:P�%�Uw5I�.B�fЛG6�}�ߔO	�?�xO����g:b��܃$�M����&V}��$�o��]�dig:����Z�WW��.?`�4�8p����(#�)�i#$W�ߚh#�"���6�Ղߖ���H��d�'iO�_�FR!�O�a�M*�p�h��y�R���h���CX���Fq�!_@��	"��،5#V4��Dt�Aٙ�s���q�	I���|�i�ՔvϤ�d�a����ޗΑgQ�:E��{>5�$��:�:/�#��q9	-�-�|��l�L�h���u�����z�&ɤ������5D�́e�Yg�{r�>��x�}W>��
�ˁ ���YZ"^ɦ��4e	��s��v�%t͹Z�"����tTتw�eC�� �Mf�'cXlq�j,��*��4�s�s�a�x]��(�HD����E4m�|��<�W�}�Q��|��-UG07[��;O�Q��!�{҆�����a��;躓��Z`�dXzÍ��{�������J@.�k͍������ݪ��OǫS����z������3r�0�?Y~���5g>��j�j��D9��~.z|�t���N�x����2�0�=]���評���hi�'r�����4l�/�b�z�iq�F�B�%�g�#z��e�fcI
a^��FQ�ED2F�Nó�#F�����`�:h���_/w�Z�Ib��:T{����t���ߨb#���0ĉH�w�7�k��'_�t3�H�4d|�<�}���C+�g�Jc�j�gj,c�ŏ�E�|Mz�^:Q��ð�h�����]˚������>{���[�lC��_{ʌ$�B��ެ�T5�a��?^8�,Q�,��N�U�j��4�ݼ�GO�hajȹ��C�y)�	f(���0�����4�t#eYn�(��&��{�/�Є���Y5<���q��LY�>��x�=K�"ψ! =а^z3�f[�.ϯ�U�ɋ�AF�sh�0ik7�,i%�rsm��i�b��5�cn��E�,��[�����L�P��˅&4��ARm�3-����5��W�Gc;Ty��ܜۆ�ö��y�kuQo&:�.�M��g��/v.�͸k�=�c��e^�4�]̬m�Ƴ�gV7Y�[Nu򊁣6u^iX-ԝ��!��9F0�ZNn�ַI1u�mR�a�J�au��ԫ#���ne#-/��zU�W��Fm����^��gfuqӛdX�Zr<���Υ��?���p�^΃g��J�1�f���d���enZ������^\�f�6�S��^�=�T������i^�&�+ho�i�е���[�kP��놌�$�n����ӂ�L�L� �5i<;��V{]�9�r�Zw�q�}[�w{d��C��L�R�u�y��4���T,�"PZ�U����$u���ժ6�_my3��3y�uЛ-{��W���nD�D
Y�P�����o�COT�<�Xy�!�Tb�������I�M�y��R�����i�N'$�D�R��|�V����]�k(��j�u)��t���eɰ<�w��:ɥV�P�۫�;��=�����Iou%垵7��Wy��4���6�>M�/�+��o������)��=v��ٽi�pT���B�tq�8��RF�x��S�
;㪦��ܼ�/����Z�I$�I$�I$�UUUUUUUUUUUJ�mI��UY6)*��UUUS���UR�u��R�Ɯ[ZʛSq�ej��������������������������������6����Z9�#�C��;c��iP�l=��my��yĞ5c��T�.��L�\��rs���r��[a6%�UDJk�k+!	�X�;���7m���\pn�)��dGS��A�]������a���-6�ݯ+�^7=���CQϡ.��2Y��{mчp<�dG�q�l!�'=3��#�rsQ�����º��7���*"�7���׮MvS�=\�3�l�c�ly���x���y���_t��GK5���	�Fhh�d��!u����/m��Ţ�]���S<�ո��q¾���u�A��P���<n8���-�=�Obx�Y�nL��'�:lu�of���z�c�[c��ٺۅ)�Z��nֶۧTx1��S�ĵ]�l�F�,j�`.u���3q�6nM�ۭ���u�S�]���'�㖓��jy���2.K�5	�;q��WF�n`6��g`�0��2ŗ�зKi�v`����.HJ<���n:��yq�.��C�Xgr{7�svLݷ������;�i4����=���rj�x1x��7m=/�f�P�N�9M�x���6D�v6�I�(�0l���:�<�֞Yzy�k�1�͵������D��	���4��\J,Ζ�e1�a�-��6�m� .F��CX��d9C�z���oU��D�,)&�X6��@nnQeх#��6݂�fn0]G%�v�X	�f�yjCظ����f���,ħV9@Ev������ļ��l�-,4�aK�X¸�dL�u-������x��Hx��׶޴;�9�6��[�bšű��8�uve�P��aM�k�]�+4j��ԫ	`-q��B�I�Xˮ�^`Qۆ���m�&lX:)�X�B�(����,�M��lG��
;F'�8ݼTF�
�z�mj�c�ݻ�nv����Q�Y[Y��UULb��;i�b������ڛ+�e#u;� סW��i�J�ϵ����y�ݱ�u��5�|�8]^��Q�8�;m+��v���{&�ѱ�YBZg0ƫ+[xŪF@fٚj�a̖�m�I����-����uI��ϰsf�'\�<���M;t�a@�����\�F�K��-[������!\˩�DUi �t�F6�J�MtKe���,�v���B��j��xW����,pb���� ���-�{X�xKsZ�6����'�y^��|��$�]-鯨�?�]:d�U��l�H�N�S���B��5}�>~��!B�p,��G�-�wȎ_Y��i�C�� �G�&�M$�t��y�A�^oƇLh�f����#:>�/"��;�}������Q�����Lw/�:����M2:A�x���&�t«���/�5���F�F!�0���x�#2���h����T�WW�ç�3y�"!Z._��x��:�2X��IdiwD�bl���hi�Fȿ��J�CY��
jI���?fn�~�z�&=��̓��;�]^����#�ўC��{!���������-J�XC�^�?���q�6y�4���Apd�����#dt��D
��ɿ����ʶ����ˤǦ��^�"��'�<X�&cH�a���ة6�Wp0���W�R{����I �oTJ�ug���lp�G`��۶ˣ�i�/7E��쐝=��ru���.�=�;����Qպ�c�(A����kއ�jÇ�"�c�Ŏ��c�$F�v�,/~���/>#HI�t���g�
	I�2a��ێ��H�,#M�C�}w�_{��g*m��y'S�p��4�F�Uۥ�GB5Ԡ������9��ea����\�M�A]]�7�`�ЏF�0j'���F��+���-���p�?I{����`NEzyѼ�1��4�w6�:~U��1��{L��z�{0�a3�\.6[iF��Νk�x�F�e}�,i��6��I�W�fK�H���o<|`��=o!��Q�W�<�h��Ha�Dt�l�Y��n ��ؐDc�)�����}�=%,>��x�ތx�?.A�r��0������'�{-{e�6E �@涨E��_�=�Ժy���yD}��7ؤMƓ0�f9/�t����l�C�����t�~=<���Kə��0�D!�������x��"+}�iӣ���W��+�i�Q�]�y�]Ϫ�c��"]v㵸��k�NH-�'��rC�	��m�N;t�#MD�ZJ�y��c$z�g�E��׍o{%��O�^�ITh���#0��a��}���r��,�G���12@�Q$c���z����,�1��(a��������J%�'��E�sț=�eˆ�}v��C!"s9�$��p"*dw��(o������*�-q�B"':^G����dT{�/�>2~�3�C�1`��}�Ig���e�eƐ�kk���m�΢�nQ��ʾ�V����&��&�0k�����j�v�L)�ø킩\��^�<�5�~�!8���փ?a�G�{�X��oH�V�G�'����p�c0¤R;�4��s{�~��oG�E̽t,ǌYk��Ϩ��ZGJ'܏�YtP3���կ�jj�'�'���+|Gt��0��;�F�t��$��H% ���)Ǘ������TRC�*�ӭ����d2d����LY�r�_Y
߮��Q����N����є4�1C�|p�cǿaxѠ�{���Hq����m��v�շ���GI	s���l8���1l1XZY��t�{=���8~� ��u�Ŗ�"�<ayI�'u�_n!� YZ��$uU������o�Hi��0>#O�XPG���H����24f*!�$F�0�{���L�5i�yG�hi�&o��Z6��:M����D�2F�cH�����1j~�������ޞEJ���L�BLģ*IB���Vx�l�ߡ��*��F!��ߋ�p�={�����ob��^��m!�!E{ފ�C���y��Xx~�:�y$r��E$P�\E�v�����5V$�z=�_i5Џ�gAeO_��X��
���ȿw�XÚ�i���9�a�����}"��l�=L��!��S�ӯumm�ش\z)��
�v�z�����G�S�Xbo9!�h�pqL[���o�*�*�m�}־i����H���;�:}�=7�{%�Dk��r����H:�f4�+5n\׻�E
8��E����CھʸF���7���@�#W��?�k����wR��9x\4n-�[�XXAj�����B�Ԗxz<V����K��s����ݶnG4���2t{�g,!�!�{gv�8Y�j��6����G�Gr���ʜ���S�/o���YY��ퟭάM�<�cO0��%i|�&�"��4���Ȓ_���+#/����nt7/�~��^���#��F���5�����BFFM{��l�#Y}성�W�yU�<}$�أ&DbM��x�u�hC���(~�(�� ���������O�n��<Do�!�p�?Y�s��[��<�_1�!��|�a��[�2�@3f(aԋ�'�S�x0珴i���i�(�dؒ(�������-�,�캸~,F��k -BI���^}3�E}��\�>�|G�Z����al��N0�qGCH��0�+Pv�w�s�ma�Y�0�|+w���OEϯ%��b��ޞm!�~�8�YY�����p��Df f<?��h}�*�>��<��^^��,M:m��F���Tb�� ^@U\\����9\uQ���&)��r�xV�m�:�ܼ��6l�I$�H�26���+�j��������k`A�G�{sN�0y������vй�\>���2�ށn�p��9v�]g�Ȼ�U`�*F^8��ƶ�:#�-an7oDCQB�m�n؞.P����+K<������p�c"�[g=;'�^�R��˅���*ZD���ɮ\���nU�vM���$0����qͼ���=�����i��ֳт�n����H�c�vn�g]��ܯ/gWb��m��ۛ��l:�z����k<z+ j�i��<�$��'�����E�\�CM�DV!���/��O1G���0���Y;h�8a��,���p7��δK��ι�:7XG��<��e����|p�T���R��
,Ԇ�{�BΜ���?nL8A��&3W�t�DQ��:F����7p�|��t4�=��|�^�?�#���B�,8$)n�{��ֈ���?n�t0�!OZ"�3]އ�{��Cl���ly��#��w,O�� �!m��?�+_a��g��~}�FK!�_"7"�O��i!(����nߺ_޴(������`����8~�p+�>/�RD&��'H�������~��t�dLx�2��҉)��
E#�YUׇ�У��,�|�t���hk�95=V{��q���oq�8C�H�VCq�L1QG!�����c�~t�����^��O��J�S(+-֞�P	�mupE�״s����v:I��u��u�땔,m�Gf�MIrUn�g��z����cy�}��Bg�فe�@��V&!�|ȳ�R�ކ(iks�rM�w������?mv�6l���$���"s�'�fT[	��i��}=>�����G�;�&0���Y��r�Sɧ
1��)�����%ǐ��Y��bx'b����#�K!�W��p)ٝ����LVD�JMh���+���P<O��[����z<M��y3H;��E́���Z���]��>H�C}��_��R��Y���N�ߵ�_���f�l���H�����P��Q�'51���a�"W�yX���(*zO#o�U��������HM|���u\~�4��-#+-���SCnJzQ��ރhoэ�xp��r'=0�;Ab�K=�'�b�G�"��=�T+W�`�C���j�^��Y늭1�Em���g���I!�!�PI#��x�:IE���E}�t�p��D�B��Q;*󼘬�����"�>�cǈ��i�g뺯C^ZF�Hi2YZ+��Wr��Q�!�Y���ͳD����ķmT�N�Jt.�'�ٺ��p��Cn������85ȓ�ښc	"�d}F���\?��>�G�_�j]��f�W�;�z{�"ȳ�C��gN�=��,��]�c%4�7T4�R�4��D���a�S�:�N��?n ���b+#�4|�$ԡޯhb=qǋ*�@�+(F�>��Mv���^H��t�ƪ;��f��ɘ�f"�,Dщ�\��=zB=�\l�K�sT0�����xǶ��0�B����|1��{I�T
�3��Me�N��7JA�'"ݫYۜ�z9έ��Oc(eb�����9�&p��*�!aBxxF�WT����_zk؝��) ��p����׈�~��:C<1@D�����&⡤TrQ��o�0~��V�w���'�,��"���r����:~d'��a`�8e�^�xW�}o���Ͻ��[�ȳ �`��3�@��\�2�`�\�#����8ZT��X:ye�������z���õ���>�dI�,�8
*���\}R����ޟhxF��T}����?S�d*����bČ|TyT�ۊ�v��]���㵸���m���h����>��Ͱ�&�g���3�u����<%���4��a�da���=H��k�A���j����}�hJ}�w�:zDz��އ`����Ȣ�b{�H���2L��2�8NJ�a��f��{~T<O9���Ρ77z8�Z��}i�_6D_o:4A���X7�
Ր��I���MZ���������ͳ]gb	���aNJFaVt��,��~�#�adm�	������hLϹ�ɜ�8b�O�%�\�d����k�~L�g�"�&H���gE1��-�B?R���6�L��BHD�;�ŒD����釾�?�pXp�H�����zXx���^��F�B�4����F�7u�U��A�z��.0�1�3�r��$"�+�>�˱���y=\bt8�*x;[�[=G����%sH��Ο%g���cR��aRGC�d}�YAN��}�9�3��FG��aa0^�z���z�x����x�9˥ej��t0GuvJcǎc$���s,�<Iz��2)
ڶt�P7TS�;�l�B(P)c�ۣ�cs��m"#���i1�zԳ�����A�����0v��,i�����N+�?�V�"N�G��C��U�ΐ�o�C"�y
�����%���4�^\���R�@�0DS���B4�G}��5�;»LԪG�_���M�ܦ+W�T0�"k���0�И��f���1ӧ��F��.}��0c�Z|�E&"ER;�L��7� Du���΅�	�>�)W�zX�3�!���Y�r��<D���<7U�Ġ�Sp��w׾,�Ŗ���I�"��P�0��REbΖ��4��BU��*z	�_a�х��N��^r��@�f�?V�;�A����w��!��k��;��x����ߦx�����I�!��%�|l�|`�$�N��CN^1�,_Yxq�@��M�۬��A���t"׻%1��uP3PG�����>�\��O>RP���;!���_t��t�e�q��۾/���o=S�&l慷�f
=��3&&��:	��m��]H����FY�v��I$��2%
&Q�UUUUUm�;[�w����q=����:z�k�%�n�"4����4<���X�W.�[��x>#�i��T�cb���ݭ�G����spip�3D�ckl+�76�|��cK�s�ť�lö��g]�Z���/j���.���&w<���[�y�TG���[oF�FA��j�m{nc��5���Δ�9s�ۏc���7e.h1���"�ꇛc����]�����4���NO����A�Ȳ6~���}#�H�sl���D��z(^���8�2EJ^��h]v٘�pz��j`*	>�\���r�""����4&RD>c��P�M:|h���ީ����z����nu��3W�1*o��蓤Y��4	���t0�k'�B�>�<�d�!��GP�u/��;�����sp�`a��8�v,��#ul�����#ǰH�?Hw�,�~��*{Q��v��͋�����kB���8y�n�T4�ŧH�qf���t1�ʅ����<E�xYxV?u�F��l�6�2X���C�DDQ���B� ��#���1@�5�FY���s�s�r�BkH�F�<��*y�(L�qޞ�!Ht�,����f��e����`Y����W�7=)�ѳ28��O����Bψ�C�><��������:]i �.���&�E�;�cs텻9p�BH�Yx�s���ۄ�=��=��]/l�O(d{���w��EF���`����
���?z]��D�܆�L��VlP��!��q�#�L�"�9վ/�6y-}��O2��^�[�"G�P�	�a�42k}诳W,y��W�_����kc&7{u�B���7;oF��H6^�������{���J����A��̮d�e��o�ލZ�^���5|µ${����z�nЉ��P`��qYn����禥�!g%,�=>5ޟ�Q�( ��T�%��M�#���>��C��E	�������?t<y��w�yI-}>ݹLi�H�!�p�U�|��1�:5s�f.z��� �p8g�$���N��v��8�V��zt�~����G���H�_*��5�?Y9q��΁Y�ꚣz�k`q���(R� �U����b�����mLhEUw��#f�2V����O4g���P1�۔�R��,�_Y��13���.����p��"����Cn0�o J_Yl��ٳ�-�`AҍDU&3������*��췌���G���񞳍m5��2�^�,�V.�.ՠ��ݭ׋v�ǃz���(D���f}��t��<�zG���Cs_�f�^�g����r<}��"��>.�1��ܔŜ#.�L���ў�/�!H����"�:�4�����FB��MP�Y����\�A�ڄ=�Y�,��W�E���C~v�%�!����$|� ��83��,���ڵ�L�F�$㱄Y�C
"�1���
�M��zzQ�`�O����$��3���a�Qn�U��d����c�/����OAt޾��15�&�s��}��wݸl\ngu$�m�n�F-��V4���Ӗ1w�R�/s��w6�(vB��ͭ{��v�x���1T3���r�ma�\��C�fb��������}��N3�1g`�F����7u��ٍ�]��E�n��p��rm�����2u^}q�F�m���L,槽����2c�g�e:�F�&���lΔ�T�w����֔�q��z���>�ͳ�.�nvN�DQ�7��u�˖�.��t��7ǻ~�8��㬣��+��b�H60���P��}�s&t���0���Q�za���r���DtN���[��&��S@�0܆��;>՛�mК�H���3%Q�� �I��vv;���]��P�Z��)y2��wr�X��3����؞v��Lȶ�9��Wt�V�Q��GKRY�uc9|���:u���U	�b�I����B�<9+M���%]�*5/,����D�����@�U9�!h�<�۳Í�����G��!g-���{A�^M�u��ֳ�w@��d��"Y�`�j��sq<b������Xs��};X��
���;ޝi٥J���nE6)��׬Ru��;�Ol���ܪ������oӚA�Ȼ�ݠEn��G�����vPn�nM��i�]I}`hH�ޗv��~w:;��8@�^���0���y�3�`�S�nt��G�O�<�A��u�g�i��r�r�fDy���h�D�����`�وH����͑�f��S�GIy��x��v�hw�H�#��F_<�����+H��+Tl_C�G�F�3ZvՒ7�ꙣuuC��&2�\HA�b�+?)�YA�h(Q�ET4�ut��.�:�4�X~�SRI�2�c=+2Ƃ��,;_Qg�Y�)�{�B�RX6P!����D�1a"�#D����w������;5���xm���i�y� �>�=�v�i铘��>:��+[��OV�OaZQH#֠���8�,��!�������G܅���Dn�&=O"9`qZ��a�Dx6��_a~�A� �d����Y���FB��gO,��v�� �Q��|����5�zo�rrНPD�g����:��DE�����$�t�&���C3�Y�K��e����=k�!��>ɢCdh�
jC��Vyԅ�|�611�H�/�����	;�a�,������v������#F8�=z��]�i	��#�EVG�ͭJ�j#�ǟ!HSޞ��Ԛ�颌���M}�mQ�!�c�O�}Q�\��Fzs��C<F���uzb9E�IvL; 6hdb_�o����\F�m�Uݺ��{8�t;yL�v]�[��uf�����\]��U΅��1{��{5��#�_!}�,��|�-@�F6�n<�,��q}�Q�@��w���"������zו�ܺ�z���*��>�1&�#	�@ݫp�V�׻r`�����N�A}�������$����k�V�2�4ʽ�!������p�mX�j[[�K��<C�ծJ豶���D�3nG�>��4�y�����
t�G�B�>�^*�5q��OT	��C=޾�+m��Dq�0�wG�]~������g��qZO���Q(�0��9Ӂ�<��Y�_|�i��<O�c�_23�ޗ���&$��6JCՙp�G'�˹
�`���:�=<�􂁝�w����^h^:�j�(Hʘ�CH�L�r�F;=�1���'`Y�.�>���A�9���Z��>�dq>��xob��"(��H?:�z.�:y�ݖOP�H����!LDۑ��Q2��Q*����yr�q'р��=w����L�x��#����Z� �\�{���G�*<���v[S�0��#׻���'H�Z:jy}4�t��/b!1@L�%��7dMTY����E}��J4w�=�f�܆6���?<^�ȯT��ˈ�-!�]׮8x��#DWyz�G{�RY~	�hʽ!i���]wb�j�2�,	��t��(]�b^��Lǌ�1]r/����0�P��ʛJ���`��I$�I �%%Z��9\UUUUU���A���K[ ��]9휤�[���녱�kq�a����5"����ems�U�;d�h���-m+�S�u��g�es�ۊ����r0ua���L���4�@�Pt�����u��W61Ȫ��|�d��j5Ր!n��<�slu\�xݗg�z�bȸv�й�c���)�bދXJ�����r��,s�a[���ِ�=;v�7ns
��z���퓱��sGl�k�;����DZ�}�:l��(�}+t0��C�Y
���CQq���"�+��}/`�8��Օ�e� O!԰�J���S#�RPç�a�"~�r�a �%#��OM�k��1�=2�<k������OܶZ�C�;��j6cW�%�n�.��fu",/�{"��X~�niIO�o���$���O�H�0���Mkf���zuW��EZ�-�j���&�{��������^޼K`�=�<��0�/���]�2}�އ�g�Y�L�!���q����[�����t��|��w�P(����+cE����T�f���"����p�QB���P�,�4�8��͗����ϣ}����jlɛ>�d�N4c##�t�v�>4kb�i�(�14g��q��6�ޫ��<��F<� �
/��>���.'�ʩ�<��]hw�iE�*��§w���q���*dùMd�ut�#�g��Z�e��s]��H�泮�(�L�<��I@���1+Gj��2,�����F�'��?w!g�M��1Qq�"O�鎣�C�ʷñ�#O��v��A�xƞt������4	@7!I�c�ӿ��JE�fU�r`�G�
��L\��y�_ 3���u�%�7n��\6o�i��L�)���y:[�9���� ��̔l���������Ddz8|o+��Pf��(���I�d|�C�ٳ�m����^�Ǥr^4���p�̩J��������8t��Y�U�{���I6t� �q�h�V�qCgc�5�]�Pp��}�Gy������A�D�Bޮ�����@���/�a4�Ʉӂ��<��;﮽kF������X�-My����߶+��Y28�?Uy��������}Ѿ��FQ^7P������qu
�K�>6�b"�0�13gH欍:F�^�����d|��8o�Ʒ��CD�ݺW�Ҙ�y���w�T(%q�*� (�/��]��.<D��D�����F���.����~���D}8d�㨂��cuυS���l�=���g[q��\d�bUj����_v�(�9\C��8Q�?2�ކ0�(6G��feS���yq�x�L�7�K!{�+�9O��hq��|�'��B�hZH@\1��t0��h�Ia��ztP���m�fO{su"0�4F+[G�'V�Di�����`���(��m��9�]+�?n��A�*�T���>,��߁Z�-#�4�.E�z�1��!��,�8cK �ھg����Rǁ���K]
 ��>�q���y��yK7i֡X.`�U�ǯz�D�_0�àW\Wf9�u�iv��k&�[�߭�q<����������i��%dO����:E�Λ6�%X��PȠB@�	L��m���P~�O4���t�0P<t	+��T%H_�X�Y?2���ur�1��8����vMN�^�lz���粘�Bΐ��A�f"2ˑNJ果=#��C��=<�N��Y)�uϼ����D�x�لb���5r�w�qB�}_;�Gu��:k��eeӊ���?���*H[�����{=7.;�(T�k���q��r�Jv!M�uҫv竫��~����~�t�"����ӆΑ>�R.�:2��Zs��q���}�A˿K<h�`�S4����`�;sq1�Ȓ0��}��X�m���u��>��Y�?�>L�0Ȼ5�{ږ�#���1��ǎ��	��0�*�����\���8��}���!P�{�N��'�)f4�$���a
8�i�#ur�?#�_d����B�)_�;.�$�,e�+.N�<'��7��
��8Rp8��_@���E�Π�ߜ6y�_�j_0�"��FS*)%�[^}<�>�W>5d� mymzX��8^y�&�}����b�A���Ζn�ކ4�t��J0�E��~���u�u*)�ĞeF1wTi�_� ��/=�,D�\�)��M�LW�f��*��O	$�P;���F��~(�_���g��@�EDL$�g�PӄY�W�Ε�;</�ƌ����x.o���p�A`�i���w��3�D�CJ#����~���W��#}�Gnj>I�gc��k%HZ�)�O������nud�º�x�z!4��n����N�=R:f���l#e�8\�_��}0���@�j����OL�d-�da��W�X�Z`?-(^ �z�~seJ�W�j3�i(�li���t�� ��g�]L��7&'$n
D��6�hO����T�t/�؂2�p��]r��!~y�@=~^��(�tŨ")���D�Z6Z��;�;p���i|Qk�B�<n@[����G���%�'��b�T ZC!�d-�{�}����n�2+_��y3�2�8U	��y?Y	�z����W�*VF�a>^2DcN��J�0�~��d�?|sG���Z�P><-a�=�/�/+�a���"Mꃞ�l�h�"�t��0����Zv��Ė�����h�cﵦ�e2p�Ʉ����,"y��E.��ѡ��"�] k�GT����0W/^�?��@Dz�d�)�9a��`�*;"��^U���sJ燞��B�Zfg�<���z޻r��;q���h遭�szh����ݎw��=�3]ȓ5]c7Wh\�e����[�:˺��^���K�rI$�I �%$� �Uu��������Gc����7��8xz76���sX�zu�s���.�ۧ`-	c69��E��JB����wb �M\ck�Y��I�i�m�ې�7s:8�7����m�v�	9��:^̈@����M�4��uW�u<��	ucv�n��̋��l�"<�l8$\:[��\v=y�3ǥE�!��\��ֻ)-Z*��݂DH��ˮ�n0yu��]��t��,+YY�������=H�d~;�����_4��.t�<�>�t0񑇐���E���{Nƃ9��FF��?F��j�a�y}���㠛�KJLM䊰�>8y�,�o��=�����$l�ϲV�/d�5|�<#��:�4NFc�EС��0���������<Qp����c+���D;�$1F����$nH�t�d�03T#�����u#��Rh�H��F��!��Yﱨ��U���F.c�'V�G�QZ忾�Cu"6�,��VB��Jϓi�$���-����s=�'��W���C��SۑC�z`Q�,�1{~u�"Θ��?�}-й���h��.��	�w��)u!;�Hz�����ύ�c`(ib�S���p�x���j����\p�!��I���b�v]�ןe˲o_(��Hf��J��򯴊7Hl"r�ەއt��U�{�X:E���}����S�tG$Mj	ά#һ>��{ ɶ���ۮ7Rlk;/-���0ڭ�tq���������������$��qB�a������x?�D��q���^�� q~^�>�c~�FD�0���B��'�iӅ�£�;�%(�
,2�gO!R"��+�j�g0�b�H���p�s�.�B��G=n_vnɿ
B��}f��fg2V���z;g1ں�����ͻ�����7�6d�F�^����1�����yAB�|؊��_Tt	��C�F� x�C�a;�wf���'k�d��4F\��<A�)���e)s���i��%�n���a�$�?3B�\缫�"��3q�+�2�X�E����B�n��yY���E�?/��͇IFޡ#e��a	5C�VFP���2�n<`7��B��v�*xt���}��;<f�yL�>�運��"7e	��\���H���ꈤ5}�D;lt�-"]`è�������H�ѧN�KH�{La��[s������F�Ծ�f^9�i��=��Hix�)!/�Pa�$0��s�|�F���+<�턯��l�בp��H��i�A�mPk��tޮ���u��θ��I�=���3\h4���-��<'����?�l�����cd�{z��e�!�)|���GLv{Ɏ s�Щ����if�E�!��"�UD�!�`��K����ں3 �|������UҤ]/M�hsgx��4a���Q���Tl��xjg3�y,F����>j̓>��^�<Eo��ꪨ*Y���<�߳�/��EF��F�r7�O���L�l�οmo�`��#F_D�$�R��#�gQ��>�������K����={n"�_ǎ�KXϘp5MД,���15�ԭ$i�z16-F6T*��d�j�f�vÊc���'۸a�6t�Dj&�]�oU�)g[��Jפ=w�G��g��mDS�� �~�������{���yN��ő$%q�3��Ӂ���(�6p�V_�Ճ�u�1k�P�R��vnQ�g{�ʟ�}�;�Κ:Q�aM����$�)L�#j�ȓڸ����qC�g썆h���]^�կj+O�g���o�C�����Z��Db�?\9:~���`�,f9��x�΅��G��ؐ�W\b�n�z:�8b�t�cq������y�b��H�i0�������S]?���w�����@���Y꘡��dF���֨|t��tҏ���>�дλ�ј]��+�x��
P.�â��'���>��亹���(68څ��q��C��;���m���˧y���4�H��8D�����t�K~���;����3�Ё�o q~�{���j\���G�JI?X�����x�Ý$Fۅ��e�o��p�;H���~�՝7�4ѓ�*���?�C�lǨ�����R��fu��Ϙۣ�*פJ�}�GH_c�M��]h�'��D逮@đLD�6M��CN,���T��7���ش���4D���hi�6pj��P��|X��#�5E	��=�����[�Ez�k�8�����^\�I���}�囜kH��e���.���L���W4�d�N5@� T�ՙLw�]�v_�!�^��et�\�!j�Ώ#��e� -0c�<�H���Q��M���c
!���hΎ!Y��*�^{b��P�728�5(]]����x�����0z{����=6x�/��ڦ��H�r"��Xڢ�m;*g����[��P�͵n*C�um���a��%�f�[��s�`�c�ǧ:F"����*�MOә��3{�EP��F5}IAU�C���f��T�C���]<���#y��$�%a�>�}��M�9-�π�������a�d��+N�K����٢���L�N���,�6A�<_�X�}��V4I�HUQd:}�� ���yy�FbU�6j��:��֖��r
a��.�I"�2.P���E}Ʃd$F��#m���T܍�*�{^̤��B7�y44�2���BC��%�)��we��4���!����)��#%H/��<����ƺ}ܒ��'�H�s=��OP��D�Tg��O�"���P6�0��LN�����,..�I���&n�����a����������ujCC1�_<��=V������%�X�`!�}U��ݘ�5c�7��^������H�#������!�����~��F�X��#-�²/�El{�zd�*�(�@kpV)q*�� �5�R�k2�\0�FD�ի٧�8�C�R�6���O0���JVe�)��jr��f���Y��rWbZ7`s2�����_G�Ŷ����O.b�Mom^��2���ތ!���G�k�3�"�:lc��- �x3�[i#�m-Ձ'|�et���Ru�z�T��h�������;��M�/Kw��L�c�}���P��]���;� fT<rS�饕Y�ir9�g*�̏�H�1N?aS2����b�uL�m��!��Q�JS�A:���1v�o�5q�5�d Rw��a�̫�i�ۧ+��v��c���x�ogm����Yt{_,F�٨���#�,���k��:���f3�ٍ:�.�?��X�k����H��a齙��iI-T��l��XR�X�F�Z���4�=cw-�m*�ȨS`�6#��vh��{*I���b4������7fD�UG�T��xgEKu�ۜty.�Z������ s�����G�s�Moz�����Y��v���U>�N-�V�1��T��k���-��k�I��C�H��v������Y6q��eÏ�7���؝�fW:�F:�H��6pȻ��V��v��&2�z�N�,w৫��vU�y4��y\ �T+Lle�ce�Ka�(�B�U��!�-"Yc沃X5�ڟ:�nA�����O����֕Q��}�zk��I$�J���������������WcT�����	�ЕUUUU]Z�R@nA���6�-H=�k��J������������������������������C��f5���J�F�zr����و�.��,q�����A���M�N���杸G=�2�:�)�5�U+ƺ\C.{q�=�u�F��.d�N�]��\:N;�0��Ǡ�n��`����н`�t�s���r�]v��se�qmrF��vݺ�9��ī��u�vN�^9۲�VWM�;qi�,)����@�0[
��v�O9�і�;��������ˠ���)0��w�!��	��s���\S�E��spz��:��o[�@5��:��4AK2�ƍ�����V�|vv�̺��q�7 bϧ�<n(�m�4re�e���;KjA>m�6���W]��Z�l�ջ��6Ŏ���+�8r��nl[�{��x����W�^rY�v.��
rp�g��ǃ5���<N\��Ǝki,(��4	E1,gz��Pu\2v�ܛ�6����S��X'�n�NƠ. A�����i�[��^M�����P�/j� ��t���p�W��މon"�r������y�^3 ��۰�f�e�Pe�aL�.ת�<g�Jmт�G	RL�c�<�M�c�i�oX:��1��F5��a^}��rz�b�oc�(��1��ڠ6&��Y��#̬��j��%u���22�]�f��3l�I�˫]����w.��e瞱&�u��u��
��/7o[��5��Vx��t���s�3+rDAw6㗉���ۮJ��FM�1���Z7V�̼#�4��^�gJBh�����,su;����^�r�n������A:��zu�]b�}Z���Gu=�.��N�6i���%��)���]�H�V�b��*��� ��b0��������qӶ\ȝ)���j�ǝ$����X������dPm���I��!��;�'s��L��F�,�	g{���pY��C2�J(f��K5��UUT�SUN[n�e�����c��0gg�iH�6��A�.������y�3����{������Y��渱X[�-�Q�l�÷.�\^N�����yM�\z�d�b�x�ѲlӪ�_ƭ��ɇ=�y9d�p��q�#S],�}awHGGb΃Ilj���C��JMI�1�G0y�甊�#�3�p�n�]�s�h���ĻWJ�q&�F��8m�V�:;v�Z�cs��1\%�h���D�Z7'��6K�<C6Hͪc����Ŀ����a�~t0��0��|pٙP��~&�9�"(ˏL���C���'���lhGJ<Ak�N�����0���,��kŗE�C�]�|�yc|gғ�x7޽�����
�»�>��g@�]�c��UD�� ������W��ʆ����#L���O�xԝ"�ʥd�(t猸��bz�Y����W�j�]C!�oy��g�6,�����zO&Т/辜$,�z��TG��U��B�{WY�t���y�bSO� -A!w�Z+�x��l��.}4��"�1��Ȩi5�A��1w>OI�W��ȩ����|w�!�@�z^b�i�����A�{��J��7�"au"��=�T�@��o�}p�r8�=�Y7���ߺ��4>@�O.ܗ�{�����h�f��CNZF�Y�q}Y2�϶L:~�8l��O,���<��t�,0��گ�8O���{	?vB,�ѯOC>_5�O�J�#��"������nx��u��W(�A�K���f��q�uy.J]��t��Ѯ��="t�=>gD���EP#ʘA�f-��C�Q���Q�#}y[@����됃@�he�I��D�"��h���/�h�14�|H��t����y�4Ѻ	\z���ϱ
����-0.�,�f�h'z�/s�V$LE^Q�1�A�o)��Qe��z-����:^�_m�h��[U�hBH�y��d*�A�g�w���d4�P�Є���Ĭ�f��VC~��Ee��Gӧ�O;��#����^%�ChF�r8�Y�pR���+�"H��`�4n�����(d}mO�hV����AvT����4ѣ�i�}�m���uq�"�΋�D?(�i��l�$U���>������؂�L�����,�e��B��$��d�g�n�czƑ"�x�׾v-���4��Ϧ}�:�!��zF�3K�=ɟ��/E~3��պ�}'g���=>
��޽�xG��R:��ҹJ�4��S�F��gO�i�<�&/gt����"2��]�9�9�D�"��>�#��}�<��5J8%$�HI[�wα��ge�j�Ac�\K� �)��x�����A�	i�Ԓ?s�w�����%r�
wY	��.��������V��M�wP�]q~��9�"�z���z���3�j&�]�V�B"P�D�0S0��A�W���UȀu	{^���q�߽��\؃�#���2JOvV���:5��h?�g�a���V��b�'O�%�(ϻ}Ttdn�p�D4QS�77�gRqD�8J`�&Y:Vy�%Ae����CMpDal��W�?�F�e
�^�ЧK��)v��LS{s��%�.������7��u(���K�G�k%�Tף3���Q�*r�΂ �|�0���P� ܦD���*iQ����=h��՚�q9#F�.Ivt��aU՝�D���L�GbFi��E}|��F�!�Z*�6F܍�t�$إ_W��äQ�5�M4n&3��Cy�z|�$��(�p��ף�2�h0�'*d_��I�+�{B�Ǻj�ÇL(S��ϗ/[�9�e�8�C�ƍ�9�,Ml""���'
dM����z8��"���`2}����Ú,@��8箫vY�ud�X�z�p�pjηK�=gQ��[=��t�j�S���q�{Ät�o�_ҹ76Y'�~"H8Y"��yQ�D�h��V�0]��BhV�@�E�"�}�ݨN��?@]�N�<����~m�m��\m�~�:n�"N!�GT�,^+~�.86hz󎐵��Z\��KN�l��-"���L]w���d\��2o_��Ԇ����~mi"����z�9��@�(�S!#*�1_j�����dVs���K�f1e�7��u��K�dRGh
7���p������.����2��$�]��ΔF[Bv<H|�r$��a(�AR�N鯤6G�WWw�����W�ꛯ8b�!pb���h�}~�Cr=�Y��<�r �뗐�!�d�D`y��ġX��[�B�"��x<�S�u�gegf��F��k���|g�u��r�ӵ�,�]ż��Q�NXu�i��#�W�*��q���:~��a(�~MK6Z�u{���g���US��Y��K�!f�L�;�v�tO��?I��/�E̚��c��1"8��r���\<6��쁤S�aFlt�>��^��~�~�5%Z�V[�^j1���n�/h�݋�uh��+hd�jnQb���Q�����m���[M�Dw�i�_Jt�EF@D҃�}:�5idN�dљC��p����F���~�s���aw���z��rC"ײ��A�S&�q ��K�Ҏ�zEr*	0���h^�3���;���j=Nn����H�Ml	����}F,�"R�V��X�[�fT���+)�_ҡ�A���Ϙl���]��Aa7~e��cSM�IJ7�+����w�B���z�,���{,�J��]���<�i,�ьz6�ô��D��\�
�	�:t���`��x��(i��?+�I/�hF�r8�ΞYN�wUx��L؃������j�'T����9A�cg�H݂GhU?^�`�!��!C�.��w��	�/�0Q�-��"
�#D?Bɍ�	l�$Y�	a�`�=�y>ϥ���N�ߥ�*�~�Q�S�b�O�a`��Y�Oz�?U����9w�vF�&+>�j��V�{��=�w�QJ �ҵ�ޫ�ЕE��	'(ՃgFlǮKf��z�c�V�Wf^�t�e�*�j�y0�Miw$�I$�@L�	$�uUUUUU��9wsф�݁�ǖ��le[���<�mۊŋ<Hqn���O@+�)3(n˩R��M�p���K9�R+s���3���勍�q[�Ծ�Â��=m�ywY���
��[���\�����Ȱ�h;j����cd�rv��o�HA#	�s�-�,����m9�
�eeZD�c,�3j�q�<,�aݲ��)6����wlEʀ���G-��\��%&vm���v�{sp��ݎB���΄�7*k[�Ɓ����~B���db��}��z3�=��t���Z�7�F�O�\Aɡ�#e����P8�=ރ�Ά��K��0��̒�Us�1p0u	�T��C��tҶ���>�O������]y�n������f#>�$�]<���z�<�8f׈�P��P�_]L2`#����0t�,��� ���z��||��^ϯ���g�p8��]�UǠ-�� ǐ�Fooc<��Xxǔ6f����C{��ڞ!d��c�G��z{��v0��P�:����w|���V����o��䙐��4�mǺ����ʶ�?��)������l!P���3i�0}^z(Q��!4�iU�>�nB�0�E�@��}��7U}(�u�z�ьx��jd��K!1_,ϡp� �6�P2��,��f�R�������EY$�˘����3���~g<%�U�����H�~����c�<���#�)�]���X��L�FR��3�����_��g:d�"�����ݨ�G[�tp��[�=�FL��g
��^l�HMa��j[tiri�����l����C�[v�1(B;c�-�;�l1�0#өH!:~��a�"���λQD�,0L�{�V}�
Hl��':�S���O̦�$�4LAG#(a
ʲ�������X��u
_W_���E�SX��{���ru�o@+��d��Y�+�@1�a���l!wf�Z��.��2)f�)��V��C��d=��\���V�J鞇d����>���߸1r}�A���<Y��A���&������u:Ղ����D�Y����@�2Gs��=�G�y+*P�W.���B>�^��B��Ig���gq�"k����%�_j�J������]1���4�Þ-!�#!,LD�àq�TF\Oz�{$���p|KNh�#ю�/��)������w���Ou@u|��`jRO�	EL��߯�\x���GA���^�Z�E0�d�bj;�CH���FkТn��t9t,C!�6�=g>5�S���}(!�97Y��#�^�aV�F�2c樎���� ���>1������{w�S���'g���r�������q��d���8�0��sd��N��H:������&�l�[vO�h�#����M7�����tcԸ����V��B�z�f��B���vrO�@���řu.T�"u	&�C�Ib�����c����S��`-�|��VGK�h���:X�o�����d�qav����:��`�B��i�e�~r��'O(y	�/�%�{bCH�h�z`�R�R�2�Tg�#�a�1Q��"H�Q�%��0�&|��3g�=COء��͋7qC���?3b��n,�Q��-�Lq�I�of}b�]Ǖ�-{�d�`6inlP�ES����8��b�r���3�2V��݅�N"kc/u�U���9��c��r��\A#�}��iTYX�cEQX��u|J,l���&�p]�t�~ݙD{ޙ��}4h�9�UO8La�A� #fi>��n�#��F+�\d�N�q������uc���B#���ğ�/#O�h�X��)4l4�@�#��z�tht�p�^�ϝ���4�������]��=۰�?Q���Q{ӡ�YD�i�"�H ��W	�<\�b�
�XB��Ov:�Y�M�N�����wTƴy���늞�F*�B{]9�0E�F���g]<ID��w�^q�H��@�&�οo�h�?z���yAe*��L�$�fȓ�h�P���v��ʰ���"\�A�K&�^���i	����!���@�HG#r;�'VCP.�QԈ6����x�����&4���>#�9# %��Ld菑bP�x�D�*ӭv"t�b��1���8豫��_�;`��Š�h�����q��h�$S9dY���{0y,�p�([�6�q6m��K����[�����X���/^\P�t6�"F�	Jȁ���Yi�zT�R���G�[���m� �g��X�"q:u߶}qW�W�'����7j��L�Z/d�d�u�"A���PH���5F��C
��@'�Wn������j'�M)��)�Nm�4��3>n|��W)9�r@�;zu�j�4�\�X�2n V�6��̬�nm-��x3;��l�`#j�g�=���2%a�"��+�+�{��s��ס���d��Quf�c�ɼ�D���g�H���"�R�^͐��lt��"�jg�uz8�MEz�8ҡ/��ڧ��_�;i����:�v�YwlYuOWn��!��:m�xyd�]�^��va��hFbQ0Ā�$��^��I�KD
#q�yM<�%�#�QDC���������,"����P��{ޚ�FW�n�Ǔ�!��u��8�`�i"�P0�d��G��c
#q�\��ӆ&�����&;ݒ��HGw���bt��YZ��3���o1t�"�B�z��r�́��B5��o;�X���_>zw��eh^x���;o�պ�X��]|���=������Q���;y��Q��H���WXZ��T��D���~�"8�q��B��c�
�=��ة�$ݶt�]��.?Y?w�蚂B�n�0��m_n�.L8�:+(B��wD��<B2��0!�R=���f�ē�L#��O�rm	�N$J�?u��'I���زG��5OP�/��֣F�22�NH�����0�6v�~���<�&�#90�>�ꉁ)LU�ʾ�N��dRL����^�΅�]='W:�/f��U��pe1�LDٜ��y�Ӣvd�lˌ�&��w�L.���n�S�;�wSV�H���;��u���tm��A,��&�r�$��]��^��uUUW:�N�{	UUUUP��*��c��e��4�,Z؛��{׍*3�,fv��y�"0]p��ZZ��R�%�5�4� �׭���K2�	�3(�!s��.l���
�)��nT�Pp��'`�&�DǍu<Zy|���Nv֘� l]p�Hݗ���%��:��1�Zi^�&e�>���C�-�u��׶����\���,��rvG>��z� �)4+a���Ts���6����͞v�V��g�����	rЄ�hݙ�Yn��������|�Sdw�X'P|w���ߝ�6(Y
W`�iQS��!�D�i���'0�d�����%L_�'�9&P�D�k��ŤA��#Ǝ����",��28��&UY:��TC�:j8D���o�K���F�ÊӀ����:�l��/c��`m��r����45�"Α�+]�")碪
ĉ*�pD@�L�u{{Ĉ_.�w�~���c�d�mI��[Æ	0"��#��y��cU)'� 'b=՜�oP�o%�osi"E"�����A��\��A�D�+��֥����}�=<���$��a�j���f�aD�)�I�f���eI\{A�0\V���_�n�l�:�j���ϾubL�7ea�&I��N���F�ā:Q0(4(�O}z<v�2;e��lȲ(ޔ.��_�d���B�pg=��U$A��!e3�L���g�;(N�a�j���̿=�u�U��8r�H�p���DW]zhy����M�c5*h�W��]�F����'ީ8����2>͜��E�yV9,�5�����P[�rnY묙�퐳�U6GY0�E����4���r8��IM���|�]���j) F��G��3.��\�a0R���#;�H/��c�M�����[1��;�Zj���D�s
39����eD�A���;��Ĉ�B��7��&Y$b�r�r���W�6T�/CC�y{YL�;��7grm��~ņ�ﳅb�����	��*uc�C��J=\Pe*xem����:c}�(p ��N��M�t	ԋn~�"�2��~���"r���w�ȻϾ�zGN�'m���7_|*��6t���=�"Z8aB&��܎�!N�"uP	0ϳ��t�y��"�?@+�p��}�Z�E>k���P�	��C�7vfD�BQ��7=^��Hs�1��u��/�w�ZH�J8���d�='�W=���q罐������2U��s�d1��D�,��������'��A������w.d!|�8��zq9�#]�
�4�8F��LbDN�~�K*@Pf		Q��Δd���DB(?��ފ�4�������8�h��B�<;��٠�#�2;��"Nˀ��z�ǎ>��&~�E�[���'H|��+��C�	ho���I��
�]6�&Q�0qD�9맙�I�<L��Zn�ɍ&�0��� ����}�8���(@���yߚ�@�\ЛH���Fj9z�1f�[4��(䍝�A��l�
o��=���@���X~H:<�!��z�;���3�WZD���+��BenL<��N�d)��q�g����w��{��)p:`�[{�Xnu�0�c���`{�u�{�l̤4��"~�d�|��:�W/�գ#Ǚ�}�k��b��f]��HR"��$e� Ѡ�.�'�O���KZ�}S��*�Q�V4D�e���&(OD�#4�}�ׂE�)s��R�ݬM��v\
K�P�[�8��>Mƭ�셛V�]�8�T��he���׵�8:��v+1�^l�mq˨E�O��	��gKV��=�z
 ��f��v�d�?]��2h땅�Hr�ʼf�;�M]NB��A�E�p���U��#]𷒭-�9�r��*�2��g��Οci���k���p�ܧ������R������ϋ��qDO[G��N�F�>n��q�̮��v��v�9-m>��O�9���7�x�Y�8��ɕ�m[1p�v�xm��ƹ�r3{(�tط����Gֻ����󼬥��/h�P2����t�E/����ծkv2b�#C7T��)��n�eK����n�y.�V��C�m;;t�4�H=�J�ö녜��Zi,��+!�Ḹ�ŏy]�ufls�D������r�A���<}��1���x�<aه�Z�R��Wٖ�KS�N��H�b���� ݣ��M�ϐ!Q��H[[���5�S ns]�̍��/J� 7�2Iy��I��|ܳs7�C1p���޾�eGOy���+����*����\�l+g�^ǆi.][�#◻�o+�X7v��<��.h�h���u0̬�R��i��j��e]w<,�����]�wI뻻y|5��ٍ�55y��޴�c[t�Y��(��VMn��E&,;��얐��b�rw�;;y�䌏��2�'Q��Ory7�7�̶�*�n��D§B.�]�;9SϿ|�8�!��zm�|ϖ�n�C�B�x���4�(��>TY�I�4=*1�iFB ��Ɯ8Y�t��^,�w+4	C*��tI����@�M(��LGב�YO�L����A�Ș,Ƀ� bq��IEDs��D=�tC@�R0��uq�$`�&���m��g��?>�V���7C/_~��M�#U�DO/�����q�TFB1"dvʐ��ǌ��w/�^	P�VQ}��y
�Ԅ�5?=J��,��߯�����6Ƣ{�78�)�Dj#V��x��Fy^�
ϳ�o7S��t[�z��v�6҈��$�q{�V���Ն���A���W¾�v��@�ڠ���=q�Ak	?:w;��W�������"H������}r��c�AC�UHn������e���SS_'����~��EB&:�C�f�}�3蜣�H�=�a���D��g���}�����TC�ϕБ�c���,�L�	�{<*M�N�Z]�^�ŕ����eP5
�Gw��Z��	]v�;[����Vi�(>��*�����7���~�u(�'*k&��[!/�U�� ʽIj�)챱TN�� q:Rx�	&����|��J���;_�ϟǇ�7�̭^.�r^OR�!���}����K{�q tK�{kɎ2)i6B ��Y�{�|(P>���4��ٙ�K���CH�����S���@^��@�1��Z����""��(Ǆn9�A<U��Xf�2M�Tf�X��}�Ib@��NNH�ۑ;��wIo>gĿ{�Uo��'�C��>�|���5������],ac�g�T�v��OA��:�_.�WDT�l�T~�y�5�]9��
`c�X��2��U�"��|F�S��C��o�^���i[�qtsM�M�M�;���f7Y�'��F��3kZ�p�6�y�"L���������EB����Y��v糾U�����LXv�~�%� �����(�*�^x�r�N��2sƛ ٰdd�n:�/��2N�|Z빼���h�b���l�3�VΦÇ��v�^��1�͸/M�7t��a�ǯם������z4zY�D"i8���Y�i3�@p�-+�.�x��Z�\�C�tmȻ�۴	ɭ�Ư�¹v���M掄%h�
��Q�f�i�������W��r�Nc����c�	8�æ�Dt���ș]]���Rگ�L�u8�g?I�]Ϋ)���CHy�kţ$Q�X�C%�-k�����sl[\�nAtP>})v[0gy���cn��:~�˴�bgd!�Q�X���q�~?T�i6�WOi���Nuh+�+6��ÁE'DRh����gM�t����]X,��6>�7�ARv����J�I$�I7���mUUUUU[sM	X72�M�e��g�ݘ,�1�����7<���9�#�Q��N���V0r#f�]��B����Yu�L6MeJ����Q�Y���R�PzW,ֹ���w�.׌��A��UMQ�ۭδ��u��]��[����g�1=�fG7X�����i��+37Kt �PY�sv�`�g=�v��r��T3�7�e����6��{[���r��;[r�yG���̯1�ڐ��(D���U_�"iH�S��C��ZdQ��.}/+➡2�"q�j�M�ۈ$#v��RE5��?+{���ⵍh���Y䡀�8d-ɝ��a�@���q�Dx�u�{gH�F���0T����緍���a�F�WK�=�B~��BPH���V��(؜E�3�|�4�V��O��������d7�B'|�7nF7�Ө�W�i���[.�"r~%7����P��|��^��)�'�4�%� ����7���DGB�� �u��2��M5����e�����[u�T-Y���e���u�u"z5�99�O@ӳ��"�s�$-��!QǗ|( �>"��y{c�����v�c����Fu!�Q��Tj>��a�l��a�y��}��i|гw"����퉗�����I�t�.�gnb�d�G@�8]a읈����p��I�N\rݹ�]:��z��/3�:�ڏ�RA��Jar��wt�m�E�ʁ�0I��'֌��8[�Na�U��禍�;}|�_�zI1�q8k�O�=�ήi��r����*>S��W-��h=���k2���7�s�;����4�:��yyA�[0�A��:�];����s)�=�Xy�+�ٚ�pkSP�"�\c�=�J�C����A��\�9������g0�6(3�$���2fNߺ0�!k����dRB��j^�+�4�30dYzh�I�G��p��p����Հ�c
@�<@� ���~�5��]��>��:*͇[Pf�k�s������=�Ȉ�Nq���<�`�Ϧ
�Ξi�zwn*������{�
�HW�����G�&ϸ�i���&ں�ms�[�P���+�b�ڸ1>�L��AI�J��7�����ה#lr�����k��c���	X���(�#�����������L�3�AW��(�\�<�+q�������%�\p�=�9��5nf��֨�o�%�pS��<�,���R�[bȉ FvX�砰v����)�H��l���.�6�
�8���!F���7��e'G(2����t���b��Uf�da>�t7�ai�z���\P��ދ������7q�cu�:I�+Ǭ�N�2"I�G�[���|��g�N��-� j�RE>�X��y����f8A�tA:�˜�ݷ�-v�md9���o�Q�m�3r�]�G�{y)�p�{،��m>��9ԯjk�7&�(w^V�	��S�/�ҳ��jE�D4��\c�x�l���m��Q�!iI#w��仴�p�v�ojxwk�ύ���j���CvU�H��+G_�R�A���:l[ʝCN^�}�'?"i�H��}�(kLAȎE$::C���E���|lq�. ��(��P�j�7��K�v���v���'t��gJ3W��
�ݒ���XAw���\H��SJэ��<���s�u��2M-Dm0�)l���Bn��삦l�Z�N��0%!�Ŗgz����튽0
4`=����[,�$� MH��昶۫���Q�����&��v3w���3Í~_C�pa�R�&Gm�&$����˯Y=�f�b����_E���ⶆ���~�;�55�����Կ���Ͼ{�MIc�z��R��z�o���~��|�\#t\7K-��'��g�DړU|�"̣Y��������b
!��E�tG�D:}wr�hUk�;�� #�����#�0�i.'!%$���w ��x���ʴ󧔋��z{^K���E�r�OJ���+O-�޻�p_@��ӣ:�{���#���,S�	Qp��J�ـ!w��=}@"�Th�s+��vd����;z���nhPL��f���d�y��yA?|n�]�ꏕ>�f��$15��
B�q(c��6:�%����-etC�BB*�W�<��|���,�J��w�|�0��M��!P���1Y�xf��:B*���\�Å����~��V���c��b6b!��܁�U@��J7`�6���\�cq��a]y+��2�
&9:y,���y<��������m�3��Mvq��p�K��xX��XzL�	>�6~ Y�j�u���V��ui�����q5lE��:pf�A�A��W�V����o�P����C_��/%�����7�YU�ʢ�T"sW	k�ޢ{�:@S�'f�wε59x_�P�#P@�ECK�u�����@W��k��MŲ�|��f�k��5F�R�{~n��NS�J!��O{%QHB�>sv���d��U�.@Xq'&	��AO�Q5w^P��Y��l��ӹ�ea@�aﻍR����!Ґy�4����g,HP�07	yz�zw�Od��� :x�H`o�(a�c��ku7���D�Xx�y�n�\���b93z!�ݥ=��B��.Y�\9�x�fsH��H ��E��,n���0�"��s}��PyC�ڃ}���]�R�:�j�v�PgM���s	�֓R5;'Wm�[xؓh�S]�ݾ�����ܒI$�HҜi)$��-�ɪ����"���$�hZ�cCn)���fPl3b49y�D�uY%C�l��mv���������/:cZ7�r�ζЛ�H�^�g��繓mٚ�M�0r���;]��"S�W&*i��L!��M���b-z����cs�q���5qf��0m(�ҡiv�
,��ƞn��dM�J�6����c�åcs���� �5��R��^��٫a^Cm����g��מ|�i�n�g��k[�#"/J������QhQ�(
�g֨k��vyw��ܨ+&��W�4�<��|�_Y�.�c}��0��E�\zQ��%�C��fGU�S�M�0�.1��$�('1�q�%i�N�(��>!}���䱴006��Ow�$Z�A��g�r����H��!�_��`^�D>2���*��j��E��/�]0z�>��G������εI��9��:�X��!d"H��k5�ڣ �]�	w�G\�c9�����MuP���dY�,�0�?�D�1}.^��������呤
cq�	�0�c��b�s<�9�]�C�+w���uy�W�I���)ɓ�@weY��a��HlG���%���Yp�$�����[�S��@�B	�@b�#���c>d���9����J1W�W6����{M49eޡ�u�H�������8r� ����[��XD�<D��]��[��BE�4�A�ZD�h\��.4���FDU����+�{�]�-۪�M�f�y��������Y��q�a\e(S]����K=��~����&>@:�i�2�ڀI�B�� ��F�D5@��~�v/P'�X!��D�z�!�� 0���nI�z���sbYC�շ���{��t@��F���׀�-��,�s�t��O��7-?��r]_��
��#XMa��w`,��;�K[��g^����;�+:B�GU���jcl����m(���r a m���"��*�����\�*��v��̇8�k�E�+nr8�����vx4�4�Vt4Nl�hl��~:��æ�!�E����}���9�O�����bR�vm�	�r�U��VE�_�nQ/���'��Vh˕t��U������I^�esu ����<�K�G�|ĠI�!��i�l��T�����4n 4���`q���*�QW\�������~EG=�~ݱPy�75�7@rVG��Z��g
��@V����k��FI("������-Bw�6W:tJ@2q�s �y�COa�o���s���B�Z\�ay�CJ.t�Q�@���'=~�41�sHL�d��B�{������/p�m�L�eB�ѢV@%��s΋5��cbv9�땻�F��IҒ�u���������z ��?V�\��"#M�0x߼�_	��6���|'���6�=͟�����W��_4��ij�>�;�8��z�{�PvX2��_�8��,�#~��49�<�xqkK=�G�����wt��Y�hf����u\�D!�;b0��+#��`�]��m�z<sG6��Ǌ��yG���7#u�Ň�Q�>�5)�$��.����f/�����W���?M/����s����gUh����*{鍑v��{5Z�!w&h�\��}|`�;�۸��*�fm�רQ�����5A��~�h��\?� �!��f� 1��D��a��Ht��[�g.!d��~����e�5�c�K�n�# ���ͪ�3���V��'o`䋂�]~�f���kvg��9��_��pY�1�k�� ��8d)�nN�V_V�d�����HT|7P��b�}���e�4�6�k�>��S��Oz��`Ya��`f�s喵��hL�r�)�i��ת��X� )�t�U�`�X�m��X��O9�� �w�w�׀Y �i��;��G��\��?�����;}�������hR�4W��FH��۳r[Qۨ:�\g]��:c�p��M2�jkdŻ]Oy=��|[%$�s�b�8�K��쒹������>������l ��'��W(�I��pdu8�Ӛ�_2 F����M@X<Q��+��\��u ���i 3�gHm��h8D����3�(�|\����F�5���위㡧�Q�ۀi��D5ɷ�u��vq��#��G����@I����@��:x�<�9gs}Q���H��ܿx�Hq<��8�6+��f����P�ےJH�'��;�v��<��X��8p�� ��C%���P���a�<�5��ec|<�Y���γC�xi�0�<�us����csǝ,Uc���D8H�p��M�E"N���9��a���K8�NVV�0����+����YG�4�G�r�{�� �C��A t�2is��}����C���f�Ů�I��ŋ�lg���S,M>|<}$밸�.m?��e���x�]d�&!Ob�Ҥ�أ�s^=�������/V�*��G�
���9τ��ߑ�Q�>%2��\�s�����L�y�3˛罆�8v��y� �\BR�����'gM ��9� B9ޠ@�׼�r����/���<`�<�<絚��ès��\��$<Lm���M�B�)-Kf��=e���A=�qs���4�Z^N�Iێ!%��y�����R�`��r�S�����#��#1s��G�~��9ΞY�S�9ʥ]A��YD8�����4�9�4�3�`qm��s����k���4�W���iGO;�C\ds�#���ΐ3�z���A(�B6���x Q��y�H�W��p0�~��+ @}�3�̏��=���u| ~ Y��2z: i�x��q�������Gﾕ*��V��4��|��d����,Se��5�{9�{�p�  g����v���9�<��Α�0�^���9ޮpQ�9u� ����9 ���2@��p���9��p2s��~T @�2��0��<�OŲ�����f�up�����"�V]�G�&�\�Y�pY	 ,�y��
�+��J�I��<�����{�U�Z���D4�� r�ۤ�3ҹ�#��3ث���� �C�Q���0�9yб�6�E��[��8O9�y80�R�m@x���\ç��8��=<O�� �ي�H���j������U���_*�� �9���8 �9�s��� �9��s� s��8�9�9�s��s� s��9�9�9�s��� �9���p�s�������9��� �9��s� s��9�9�9�s�� �9�!�p�s��s�s��?�� �9�q�p�s���� �9�q�p�s���� �9���p�s���9� 9�s���p�s����PVI��{f������� ��� $ ���m��><z��HI)EJ�QUJ_f�@��S�%*����v%=��M�2R��!�[b��iUUEI�, �      9נdi��  $DR�
J��R�Z*�U��L�T$�(+ 
   =.���yi��\� �) (t���=���q65��f�*�k����{g#���J@ݞ7��}��nٳ^��Z��>���n��������m<�����ľ��9�w׻�{q� �R�� ��2:����������
4�tS� �w �|{�u� Ȼ� 7�晨7`2owv��0�!��R�* 7�<�� h ����g� 롗�>8��6f��w{8tz�8�� 1ݵ�@ �/�@ z��$*(R��`r��:��|{�p:���g`(�`�� ����^��/��`t�cwi����O{z�h��oZ=u�� < \�K�% � ��1���;���=�Ӯ�+<w���;��o�޸�Ϡw����>�W���zJ��!����6��t5�tB��jk@�C�G��M�x���������>���[w4���wN@<{÷��ѯ3"��Y}B�*���
�
����T��������0kz��\����o&����lk��mo��}����w-�������[��=�zn�S�j0��i��T�i �H{���}�}���=�rP�ֵ��v��{�Lf:����|=�V�{��Pu�篘��v�g4�>�:� [> 1�^ء 5�3]�
ױÃ�Vվ�n���o�{���͍s�"}w۾��ـ�=�w�9��Ƽ<����sו����EB�@
��������hk6�y�5ކ��N��i�w�<�,ԗg�zɝ�{�b����t׾�W[l޷י�.#m�>����[��+=h )�@JUA�� Oh�JU    �2T�3Bh@�1?7��)J��0&����!)J���0@`�P�%BE?*=OQ�dѵ<S���O�{�~������0���U☍��ޢ'w��9���� �I`f�� 	$�@ BI!�H I$�� �IQ� I$��@ �I-� I$�� �I��G���B� ,!�2�
r�
a�!���Ć�A~�@FP���`�f@��q<y"�(~}��^���GD�S���t�Z*h��h��N�{����Mџ0�a�3Tn`ߥ�c��J��nCC,�S�1���[�J�^(�f&�m�f�ڦ��FT͊�ď㪲�`��Q������E�l�R��,i%�7�4v������vv���n;�t�X�Cؚ�鋡��F&�mK��S��"���/s�=C�t�%$CƮا�{KY�6	y B�cA��q�&�G�0bOѝǰb,Sf���f�z1�$�p���e����V,�˱����d�$ \92z"�GK�����b����*p\�W61P�0\�~hZJ�,�^�HE1����ވwZI1��6bZN쑵aa��7�3N�J�ۮ$���`&7uA�fP��b��rZ�e��uiB1�e��NnE�fdӼ�c��r�Ѕ��tsN��zv�E�]Ip����H��ñ^�2�+s�%$�@�Y��{r ��kk�ͤ������<��_��|5��C������:��(J\�х��t����Z��{��w�Y���f��oV �Őb��ڧ�Y�NC�}��np�6�J0�%b����A;sdt�YÙ�-7`�0�Ywm�FI7ki+�f�KX��mo����SZ9�{�(��&�K� ��u�e+�b�2e�� �Z	���p��� �*�q���ME��"U�;s@w��{4��t��aa��]�e��W,Q�vSo���Z�z ��,���A7�����^f�syh����{�r����sX�����������
C�e1b��tm�7�I7IH�Z^	�vs�:2����ϖ�k��u���f��ڂ�V-���=ʉlz���v�F��@\)c�KQ �)+�6�hQS�~#���]	��V�#����8����:�A���[X�%��B��`D� �M�k�<�:^��UF�D���M�����BO(�p�	����P� ~�<��7�[u2��&�&��G;�����vӽ�G�C�?��&����'��Ȁ�2��t��K{KM��+��~E(�YU6��ek{BL�]-�P���i�oǹh"��h�d�g\���;hXM�A���T�����DBf���=���su��K�f�m��ݕ�\ޗ[o��Ŏ����m9�e�Ѱ��4v�:0��B����to2�RT��՛Lfe��gt�U�3wp��a��{+"�Ǘk}�N�����[��?�'��4�d��9ӷ��M�r�u�K������n����n܏��8�8WoL9ɉ$���%����C�#uÑ:�1��}+�5��HylXz`� ����+H/4�s�e��^�K[��l�e�vcYw3c�s8o<_;��N�rlS7u��N�7x��^R�X��w�8I�ҩ�U��@��;�釮U
Ek�����`��Z�P:�?�:�ܺ��
;�q,
�І�$�C��"aJ�P�w7 �͘�; %v(�nSI=��ݖ�@l��kHݻ���9�;N-J�A.��T�q0�S��&��9uU��m�7W�K�t<<
���a[+��K-7��\��G/KY�y��=4l�N]�뒺2� {��L�xl�x��{�T�cXIX����>k6	�Q�Bso	��46��Bb+���g �$��7��|ґ�DU�3\AN0QX�,���Sm������L��C /�h^|����a�fm�	L/6��P��#]�`�h�,���bKEa�{J�F+�Vٹ�>��޺^�5�"�Y���[���YJ��+���VҨUlg)�헦��w�+4�7#�2�@��(6��i�M
�i�H��n��VB���2�0�V���+�P]�`�)�.*MH��	�a�?���vn��?��s,֑*3�%H���9!3]4W�BC�At�r�s���A�1?�[����9e�$8�fr���J�]I��hPSC#���[&2�#T�	u�7ZQ9S!��k+\�p�J��9V^!3����F�KN1�RsW�ĩ�����}*���4�m&v��7E��ތ�]h������35κ�'j�5��u60�(I�*J��&�BDġ��m��3z�Kde��on�6աÕf�f��!�
�t>�ɨ�5%��d\*��wmf�t�E�������`]8��~��n@J���g7�N�\�;O�]�]��y64s��$��p�.w�qF�C����C�����n�0�3cb�5*,���㽹��U�}u]��hЌ����;e��nԄ+1��=̔.�	�D:��X"�F�l\)1pؘ�U����R!���8�3Z��s���Gu�ґ�^swr4ۗ��Mr�0m�yf�n$�����Ӹ��q�,��8���1:���=�3������5T�	�oHm[�_p�6R���_B!�c�a8y��ww���:r
Y2�zՊ7�Z>�N��Y!.��0�L4��1�_n��E����t�]NyiM߈A�$p�N�#NfV��l���f��f���4�3�cu�]bs�tk�a�}�#̏R�BPk��54;��KRM��y׷/���a=�s[-cv}����ɟK�ν�?����:�8%kוz7�n��n3q̻��R5���3��ݹx�ǆ�~P*Y�J߯h�� ���[{�[/y�[p*��F�J=J��8��(�望��Ǝ����6���ؐ
�2��w�
k���5C�(E��DʠQ4�J��"�C�gM��C�>��fg0�^�sB���4��M�����͋�$����Da榏8�$������5[t�����N�u��e�f�E�y���X�I]��5!�4l�b��5����k�'� �(�0�ݼCw�ѭM4�tsu��v�Wn�<i%Dzn���%��N�6f��VJ�fJa`2[\	�H����pA&�6��'�'oq$��h�i��3rG*S�T>�hj�#�)j���[��� ��5j5,�=��E��`V:����r�UQm0���r�i{��F 6,U��a��ݑ���?
7��G3�T�	?� �A+��!�A���Y5��6�ՌEH�SX�&f�d�Ӻsr�����;�݀��PEކ�d��(ъ��[�Z���n�J�B�e��U�A�~�M1u�0����tB��D�{��~і�/G�؆�v�7f�	�7!�Q���ǅ�w�{��Ǖu�#R�)�A��9\�<�{�l���#���q��n;7��N뛭�yR�gh�鳼S��:V\��&ص�B3ᛪTK�"���̌�CA�؎��`Nk���p�.���3�qmS�������׋q�d�&�z<R@��}5�q��s���dnofƖ�����E��7���1mbM�&]���-v�w�+��9Z��g�f"�6��(���-�p�-qk�<�>�,�%���Ff��L�o�VPj�h�p��'1�������9hm��-���Y%��&�]��v`����������%Vˑ��C���k��D���J�Nb��6ú��_��֚Z�rƱh�Vvn ɉ��mK�Ų���T�ƏiP�5�K3>i!��;5�����Avez���t��E�^%YluM���j�ܬd�z�72��߳Yj u���=J~�����Y<y��0U�l�F^�6�V��+��Q��j�8L�����F;��w�]�� ��pfbOJ1�����v��):�|�S��6�KShJw}�k�3�Y.�K��aɷT\��=\R7d!'��x�+4ĆU$�PB۠r�t��4��a0�m#�!�����$+�x*�VQvs/{7����i�F!(�9t�z*�0*����b��G���P�nʕe��ֳxΪ������b�i�W������F���yL��y�����61�0�5u
I���2�%	��6���k��H	�H7������=W4觾��$��`�~����RDռ�\]2���@^���8n��V𺩄պx]�˫�ܼ�mH��ԣ{.X�QcU��EQ�5ַ���N��֎���-��U�E
�M:aM�.Z=��ocE��qγ�>B�*��O�,C�Ff�3Y�!��c���HA�Q�Ʉq�;F���>�D�Ao�"���D�F�`�@!�(J�&nB�ݧ��L������ʭ]��i0�Eh`�I(J{Xbets�^\i��;�MM;4ow9R�˭��T�v��^�MT��lF�r�b�:!1ѫ�\��p��F��8����k�%tLƮ���b�r��sUwStf������tKhb%s����4�]gve����s��f��5���(uɚ��w~��>���F;�E%:���f֛��Rs6�����[{��{�i���Hm�Y�4B�Q�m�t�uD�ڤ�K B�F�0�c)+��Ct���L�Yu�:`a�چ�UY�~&�F��r}��g���κ�4"2�����ι�u�e���� a�fP8\�����4�b��0AV&�]#�d�F�b�'��:�S���/oe͓�w��.��Xn^&n��e��Pp�b�+S�V��
�s���.���4�C�zN�2�C`��,�&NϞ�q�a`��%ogԽѭZ��6E�ʼ�5��j���W$��+�ܪ�9�%��-)��`GI{�en������vi�ʟ���D�C>�'���vgq�� �6�D��f�Q�7���Y��y��k6M��Ӻpe[�a���&���s�Sz��ക��@Ҡ�y���,D4QAbj�9R�S�$:x���m�
5L ������^�ܝ��p�M�3`{��hY�Úb�K�9LN�w�%���ݗwkh�=�b�z1�!�/d�:U^
��U��ϓK��՟�.��Fт\y��A˃��h��t�����KU6�BKL�-.�\RڪW�+j9��b��:N阝i��B��6q6993#��L]�d=��c;�lA�.�ɲ��ݵ5p�BQ��Xfh�"��1J����"���#+N�eܓ��eir�Sp�S!�Z̆�ث�@~��ڤ��x$̖2��:ڰ)�[GF���±��5@JE��nق虎��\�9P��S�ٵce�7Zf�z6���9Jop�x�x��u��V�%�t�Q��Cw��W�^�:�/y���F<�*�<�=m˽!�B��E��5q�o��l�.o�K�Ц�e	/��8f�V���31'��K�޵6��A����qm�Ly��D̒���n�F�[ݧ16����J��a2J�4�B�X9F�P���B�B�a���0��9P����d
d���a
dUZ� i�ר������> m~/֟��4{}�x����@���n+�u��q�;JvD�o#)���Xbk!8Y��VP�ܻB5C! t�mMiv̾	N����f�V`TVU��ݻ��sy���W��La��u��7��9���\��7��Cm�z���m{9��-Z�M&s,��d.��P���|߰�Cک�!��w$�!�� i�8�-�8��HaBd��2�ad����
d��{���;���ޞg������	�U%���<��B�X�4�ad�}�i�y������d0=2���p��y�og����]���V�9y�m��d�l!����ABdUBd��,���0��6oC��l����f��0��hC�!�@�i�@6���ʄ:�6�a�P��B�� ������w��V��_]�Cg�׀                             H       ۭ�[��/,˄�K�    3      H��                                     I                    ���@  f]�d� �v��-��$�J	$]�( ��ٙ��I$ � �  $��  I  P         �      �                                           f%��  I��,�  f               �-�I l4  �He̩    H   &b                      �  `     v    I                 	$  A�                                     �/��ٺ_��?�S��j�S�� Xế������U����)�6�vʔVa��\����s���5�|=���3�]�1��oJ�����-H82&�;�ie��9�6jť�ufn�.1��h�b��f��8މF���]�|9�w�8�n�C[IC�����)E�fmi;�:=���Ǧ�����)[�©5V�Z�^���<��G,jw�m���ݬǔ�&љI�;�2�r�k^�"JEbK��r�a��ʖ��qc��V��3��R}Ρꃒ��К��'W�.��MR2��m��V���>W�^Gѹ�g���<�+#���_lf�iژ'QrVl]Z]_�s�
��8���*���������:ե�oK̚�
�)�B�m!�K9�������ċx���T*s5֤��t�
��Nɋw9Cr�.�z{�yT���,ʺ4�nr�"�c��yv�$�
�Ռ�Xl�,z�s���9x��h�m��M4��G�)t[���:��������ɤ,�܊zr�X,&l+���,�зS��լ�A��i�Ue�q�$�6L��/�'fvz4o���Չ`Y��3�@��(4�l#���;fD�v��������M�V�Ga5r�ދ,���8S�g`��qܮ��{Ϻ��;�-��&L�=��/�R�eG���)�络|6:wt! Z�O�OZ}�D����C�\jٛ~#Y�0)���z���r�e0\sz�'�dx��b�t6=��F�;��o�߽�(m���M�`�>���Lܛ+5��h+�^����uvz6���~K<H����Ы�q�ibݾY�+D	��Ţ��@n�vPTs�w=��ͷ'Rd5m�8��m�svwgY,�_7$�Ʉ����e�k����Wp�qs���}\Ιʚ*�]w)]�.��V��"�o��9QIRH�MS�>��e���r�#K�O�r�&��m�m�\Kf�؆J�֟*���mf�J���UjR�����$��UǨ�ff�q�}�Vd��ݬ�*qTT���}ӪIM�ί�|�'��R��W%�N(�4>�;MK��O�+;d��ey�g�����5��>��z����Q��%�;ZT�>���V����Դԝ:��x��9q��t��l�@o��IŤ�m���i"g1k5�2Is�n�� 3$�I{JgI#K�I.�D�I����d���-�4��#��1)֘kN=�D�w�b_�E�#ٻ �Γw��Ť�d�6�]u�D�w:oE�Im�y�w1��6�t;�ޕ�4z<[�Џ
�l�=�vd��Ɋ6)���rF��b�o�ܫ�DN�(�m�Ի�����1j��e��t�8(��hbP��� ��A�[���(i�����]��fY=6�q/�$,�p�����ך�V����wDu�E�a���Bj��x����٥w�D�'1�7�{��eNv�3�ټK�Q��Θ��(�tpfO%�0��fk��S��滎ZǙ��^���!㮯�s9�{N�Ś�f��qw��|40��ݙ`!�i�5F���o�Q�����	'ӽw�2��C7C��P��3֠��r7���ӧ1�.���H��V�H1�7ݲ�w�*ݭ�i-J�ޫ�oc�����1�z����ξ���o	 E�
#G�:L��Ii.Y�Ќi��F�{��~x��]�*<{��U����ӝ�ˢ���&	���� &'�6�u}}�<Z�\����Ybףm�i�k�dP��)þ��|��d��V���3;�'�r��k�ལמ����C����L������i��J�|:�_0��b�ܣطk��n�@���;��d��:��3�ss���:{�-�}�ŝv-9)k`m'�����1>wbaX(��_S���8�j�^<��u���d�ʹ��v{�\���}`�EDSv�~����a�K�B��G�%�Υ��δ�)�Kwv��P`�=��O��͎��z�g�rGx������f�o����5�|t�j��b��V��jtN�6�s�ٓf{���є� Jo�J�{ڏ��5��#,���� ������&^Z�Ƌ$e��_!�"�_�J�B�Ms��[$|sJ����%iĮ
�w�=�|�y�}3ޱ��n�9�ɪz���������gY�	E����Ix���#����35ӻ�z�|^����(Ь�mb��˓m��&0Q�o���B�V�a���4��ٛ��\*�>�����7��,=�V)�aЦ���b`��ו5dX�����L!�R�DX���]��G�n���ZY����Uy���'>8�u�p*�Ռ��p�&s��N��|I�[=��g������3�y�w�u_q۵��'0,�/B-�h�R��]��K:�q�
D`=ڶ��w��zvt�4�n<���q�111�f��a����酌NZ��bS��3�.�]s#.�!�ś<��Q�$��I+ꌴf������uqԐ^�Lfn�뚽7}����T�_KR���uayj�Py�ȏl�ּ��(�]F篗���~����<�A�dA��\���Gq�=�,e==Z����D��4������Q����T���q�v��&Z�zh�tK~^]�+�����zl;�r8�N�kz�ݭ�L�C�5��E��_y�_*���x`:�����l��%5��h�,J�%_@NU��fJ����;wV� �����vm��:���ːY��1�XX{;1<�٘�#ۗ]�k���.�������$�����ͼ�{hR��Qh��V�B�>2���+���i7}A4�`��:���#����'��Ԭ_/�t���e&���ۻ����x+p<V��o3�Z��}�m�v'BS0�x����smaȹ9Y]�F�H-��Covnl�Ծ�Au����=mn�l�ϙ-n=;�<)��&L|��UԾn�]û|��F%c\���u�S�)�7�i��&��ߍ�l�y9��=��ue�J
��ޖ=���e����������"�󾬧E�d��vx{3���2�^`�WOm�;��Ӷ��9��� d��}ʝ���FV`�tu�F&+�w���IG=$[7�̭��e�>�<3[;���}�M�=l=�q�������z��rvJb6�����S'�mn��rݏ��x���Ka���4e_ɻ+
=�N��49T�9K1�+AlZ[Ǟ�컊XG����N�7t�{���{���{�Ճ��͝X�� (JS���p�T��,�3&�<1ea�g�S.��ûv�:�!8���S[kz�ĬG8D;<U�����r�T8���:��X7�2�S�Fe*O\ͳ�U��y�&��uzoFE8�=8��B�ֺʜ��ј��p^`t��O6u��ee>���܃��K�}���U��2y�zZ:��Z9݂�;�ܗ�͝un���00W������ć���gE�nL!��- ơT	���� N�f�FlD��W�W@��)-�%��Z��f�R;�α6�5ZykE�\�XcW��]�s.�ʇ��:�fs���؂w}`��r��:��]X܁��ӻ��Ż;_��2ےy97f���^�����ҟf�S1G����w��vZ�V��`�������ї�;³t�ѹah��z�Q9䋞Y�Z��30�;K.jj��M;B��;g%��ޒ��h$�3$���c���{����{;lu��t���Y�$����X9"L����H��a�u��1��=<�zk�K��!n��T!	��V\�7##�-�]�^ef5-��$nl��z��%v@f��n\N��2��z7s1�·m�x����vqzC�D�������=��ث�5�}�yC1���͝F{�B��V����8��.�W3GNŤ̳�ͣ�/}ZE�_L�d�x�~<H�?��5`��m{��0=�]�|��vwss7���َt�wϊC�0 ��E�lX1
�HeݜDF2B�U/����v��ў57|�D�N Km��0F�
�.r	���6i\���hc@�$y��N^�y��8��(_�$���d\�u�5�c���"L���v��9޳z�u����d�h�2�\cvK	�i��h��������x��#�J�e%�{#�z����y���l��s�D�u��h�sL���~j��1�!Z�X2wj雺m!f�����t^��
E>�6I�&���*�x��^�B���$��&��M,.�t����ȗ�]Ě������F#�V�K1��n@������[R�C�4ű�VaPH�SQ!l61������a���"3���5��F1�}��\L��O�@���B�L]�N�"�'����Ĉ��ش��6���8�xF'ܐX'łeok��7��?r^���n@�@��Ǎ�d'�(#0�KY��(��)M����L�k�/�G�j�
 yyd�X���a�[���H��H�h�7����c�a7�R�T��p=���Ry۪;��x` �A�K4��K��Hv�C�}��n���������\�c�K�T$�K\2Y3���������1D���I����-'�ܝs^�k)�
0�Z����Y7c�
��5��M4�Ss=��T�֎��%$��M�ܼ�g2�͢Xs��>3�������P��� I�����O4^�����ۛu��#?A�z�鰜\Y"F�J'��Ό.�dP�10��8��%���D~S�އ3��Q�@�O�)�
�l��x��
e��j	hD��k�/>:�+̇�F�sYZ�9���I�B_&�����&��t$C��m��������";�H��E� y{�A�������&�1�W.O��bm��^�cN8n9'�ni�����h����7/�a�I���]Fxz9�<Şe�^K���Eaj�Q�C�6#Sq��{�D��CĖ�^.�̅��+�A*|�p�
�~�B+d�I�"�| ��Kt�dl��F�0�7��L�Q��ӒŘ�iUke��Yg1�tZ��imh�dB���.m'=�}����t���MO+��B,/���'u�r%�L�7�g�^�fn��̾*_u��b�D	���UW��Vݏ�%N,�����(5�C
�+p�+��0ڟ!��o��!�F�)��.�8z&�1���4�3���Bb��dy������ �����A������#�zUi���l�jL��[;�j(�2�R�u2�/
˾�:<!��-�8ы��b,#���������-U��ίhᚵ�W��ONћ�#T��f�!�Ђ:����@G��{�A!/�f��_,�[���{kI��Ufq��gs�UQ��a�&H4�HV��,�9Jo��ئ�u��Ø�)'�8: #B���H�$�w��pӣ��X.z|�|9u�~��✡b(��X�&�>��y�o/�(&�|`(z�ʷ2���r�;Is��a]d��.�˻�X�E/p���y/�9Y@t�-s7K��*}��|X�=w).Ҥ�O,���h��Q��0%j�Nb�
�ݒZ���g�@ս��(��y���5H�l5�>�v���xj����.E�1�3����,��\�ҹ�B�_oi�#��묦��:�z��SF�޴����V]��/�$)��>;p���\b����1� �C�IZ�,]"�03|}�{����Q���Hu�ν��	��@�N^RWx�с!�V��T��}��Ic�uHcs�f�r��&T�ۗ�R�wqqݩb�فX��CǷ���0���ۿ���P�9wC��Tc�S��WV.���A���ea4��snjCO �	ŝ���+�͕�k]���k�k;�����Ѐ�I�� �I���� �a` $������~���U�����V�x      �izfM	$$�          IfU�&&1 �L�@$�   �        H�@ �@ &"I-��@      �H   	$       ?����[��?�V�MΊ�kT�'x�tX쮩���T�XwO�/��,(r�I�7�v<�y���h��Ǌ_>�7��z�w����:˜�ӱg��d�y��Ͷ��V3����	�k������s:-�g3��rK�f-�>z���}�D/X@5d$wf�.كs\�s��vDǽR�wM�+,b�5s�M��\̤_h�� ��5%�qg�����v��M��{*���o�/"/�k��g%�M�޷~��MS�OM|h��c�(_��j�+2�88
^rNNo�NIpw�W�E�|9���g��ӛu�H�����ǟo��9 ��9y��s�<�c���ݝ��5E�ܟ��Tm���缶����|�>�-(�\3�vh#��it�v�F�$vh8�Y���#��+�������8�b���p�i,C��Q���<���,��
����w�م%�d
��)���UJ?�ċEl"=Dyoef�6��y�&淽�5+|F��P(���l��d�4L��bb6������:9�~�+P�BV!>�%L<���O8&&f�eԁ��6B�*H42�rj�J�V �Z�	�WH��Wʓ,�p���h'���DZX���
5D$'�C��@��ۨda��+���q%�d��r[U�?�R6�Ar�IR�������ouQ�m5w�T�:��^w||�Rnz<^OS�fs~Ĳ�;���D�W����~��_�����    $�$�I  �  $�����߹�Of��a��7P��{�B�Wr�|S���_J�Bpd�B����+����ò��ZSH��O�0 �!Dp X��]*���03�8uE+,���/g� 9��m��_m��Xl�2b��-�H�� ��s��!��׫�Ǐj�Wl�Z�LM��5�oᯫO����֗մ�zﾲ��GRs8�~����M������x`}�~�4��]��ݢ�q�8�*+�rc1�;�M+��&�U���+���v\5k�Hz����6I�~!ꦑ{]L�����[N���u�	��F�e*�^ս�zϚ��V\��n����5�5#�>���A�����9Dp�a%�f��g��~"Ϙ�}�i�
�CuB���0?���^~c����쓎S��Е�S�#!K�R�W�$0�`�b8C8��xi�%�Ӱ�@Ҹ}�����z�1"���[������4�,
��x���_rKDE��Di��m$�I&�)+�޽����v�..-y�e���R�/Z��=9;0��t3Oۇ���G�NI7X�?c?�G{�>&���ƓM���<~	!H%?+̩��2���w���/�{���٬��W5{���g�vS*����ַ��}�e�/ۍ�Q�l�XO�X�����㞞{�������CP9��4(�&f��aV]]k5��޸�ⵂ�e}��������+�>�}�����,�z�w���[�朽s׷����
Bd ����9w�>
O:�]v��<����� )ľ�8�#��ܖi��WF��)�ޙE��Yܥ뼯4�r�)Yfc�	K�XQ�&�rD�1���HO_^>~�;I�r�e4�)��`����H~K�������:�4��5��b�"���|�ɔ��\�F�]N���ﷅ��St�fM�ł� QdY�g��L���ާڣ�wV-��(˯�����m^�^|�"��Ş�G�@[m��lp���%UUE�R����O.�9Oa�ܾ���`y�S�11u#�	?| :���џy��k|�gݫ|���<V>��oR�~�+�jb4D��a��OG��~����D%p`C��B��R�_�a��]��Z�dU ����b	`�Ȃ�(��
*����b$`���R*� �`��,��C�n�w�_*q���:˷4��t�L��ۅ1���u��%��>Gui�bX�:��v�Y�f!��IGr��¶��M���ݴF(m�y�ۦ���n�r2�jn�qryD���V����M%�y%ҽU4������L��z��� Ms�� H��$s�[�`h�q�#�ё�5�v��w8�z�v���U����(�ش�D�^_&؇�����=�7����ޓ̤��m���o^��Vj���v@����R��<�}U�W�K9�e��@�"l�Ӈ��_ʸ�c�?<}>sZ(��(��(��rڃ��qf ����*sS7�g�j��yY�����.���1핽z�$�v��kBق8}��L`V`�Ώ�z
���S�C�;��O�����"3?�Ec��ß�l�~���x�<���4��2i�V���ѺS��u�i.�����\$�Y�g�ӽ��>~��r�Z��b�g�b���s>�������<�����q���5�Ϫ���ǌ!m
<˧5E^����پ�B�T7�:������n�Jo���&�*�}��A6��Xd} �1i��P���F�;�	#D+=��L��i>�}�Q�zB��W5w{ϻ�w�����΢T�����"HFE"��(�d�
J��D���䯯��f�|�n����<�͛��=6u��S]f=jR�g53oY�4,�8Oд��!u��i0"85���{�_�����n ���d]7�q�u���+�b#k�p��
z�Fq�l�퍐=�?�|><Q�����#m�#m�#��vF��
/�B��]�,�µ��Qj�U�f�ݬ�m��a����~����x�?�1v�ɘf��Y�lT��E�1�D���3G����|�����$'�l�4���2�l$���ٽ}��o_�>i�k�i\�ۇ5�V:נ�
`	�Z�?C�xƉ&�{0b�)���u����GF�X��S�'D>�B�u���9a����3��I�L����:1��eA�����x	�xڍe����k��u�O���i��D�n���s�mO������W���1AE�D��@bEAb�$XE�E�� ��Ab�Eˢ���8���m��Ò��%s�6:��Z{�M����+]����9Rf�A�8b$O�O��VYb�s՜�L���~X��.��� s�Q�SlSmj�k���Nҵ��r���s/7�9�h�w��H���7]ޭ����  �   ��	$ I  .��ڽ�r��{��s}��3�/KkS�ıqz.�-����-5R �Lq��
mQ�-kb�X��6ߢ�+Q<�b-T�*D`eHS����]�]�
Y�D��6ܒc�ԑ�+�O�ND�%��	$p#��-!r�X�_���_���dSK,����Z��:��>��������k�:|�!�!��vv��U�����{{��]L�Us 4%d���cc�2�@c>�,]i��z>b��h��bRYmȺ���+U�-��o��-���u2�v�� �
_RF�b��*b)��+�y4�U����֟*k�Y��*:�]��]���:�c�!b$EB�^M�d(B�e(K��.J5Q~�S�WЀ�D�{_w�Z��a�z�sm��kZ��ʣ���|�B���+���pD�zR6��+�E�X���.�����YW��G��#���Ƚ_Hf�IoN8����r�_V��<v>�5�0կ� ��f�G�����mʃ(a?t��JI-��m���y���1&�F8&1��a����LN���ilީ��5_X����u�kU���$���{4����j�������j�7��2b�M�C�$�0i���j��su�M?i�W#�0�������f�7t���׳=�"TT���o��q�3��t���	�--����V�]�Fvl�
�� ��1��T�y�I֕=�	!�"Ϟ��q/�ˣ��8���xx���q_�/ER�/�t�ai����z����6��kt(w��&=u�		�ں�n�l���ޏ�P/�n��_V(*�"�]�Ԑ#N��+�ڮoW��h�g����ʚt�n�{���w���M�>�W�(�]$��zv�<i�)�z��~B��>(��~>#w����ۤ}S{���[l�u�Iw����\�y��v�!�v|�O���p����������t�%��ΑH���~�~���r�
G��<A�M��H 1쒷�ޯ+.�_2����9�֋��Lx�Q�D��#�P@EX$ �c�_�/ݢ��ӻ�2RblM�a4�8�\�gΟ�����Q��$G���#4���,����N <:��w�u��;|�,�=�y�ˉ�Zg\%
��K���H��t4�:����z,����4m����~�}�i]�G� 8��a3���谵��(u�e
�J�Q��,��`�BU� R������Uj�����.��h�*���MZn�+�G3 �X7}EQ��Ќ|���y!݇i�u:��5���u��,��r
W�T��m��e�+�	7a�}�)���9����r��ܮw�u����W�!�]�;�q�ύ3V�W]uʹ�6sqy�W��?^������xm=�FO��j>��U]���\����u���P#>����Q!g̤��c����B�*��׵�ӎـ� ���= vW�{���8{�5���x%��(w^K%�'y<�ej����rp莈�շ:���.�E�jHM,ؚߢ��o���q�uY,&�4���\G��d{ﾀ ~���l�����-�2�Rt{��K�撦;ޭ.�ƳRt�~^4�I�I�jhh���l_p�w=$K�������;=��1����F("���ʠ�"R*�)�B�h��
X�bR֣��T[��ܯg�K�s26��������+Au�kiWUo���R�@nG���<�>6� ��Vmin]�b
�۱���$���ӎ�-�����#���/ ��}qC��M�熿�&*O�@`�d��BI����y$�ݥ1YP�� ��peFV�'T�[�Y��h�;�o��*�5^Ra��gK֏�݊jȋ6��JȠ��i���y t=�k���6�:�<�vn�R�\𻭯&�4��VB2(�D� *��"�`�y��H�y�M4�s����2�Amh�A��c�B���(�s��]S�Jz��|7&�����c�dΙ_}_Uvspyt��x{-l�D[�K3��d���è{c�+�#΢hf^�Z�;��gU$�/;^ճ��}�(�>���3����(����V�p;�&����5S�����w��VQ����$�őB*� �Y$�B/7�ouSf^]�} �$  3 	$ f I    d&�z�iu�F�^�fn�ا7N�<Zs���ꆮ<��^���3���_s�$`Jrjx�v���$e2���ֲ�K,Q�D�eߎy�V��n��ѩ���$�v�L�Fے0���9P��p�f�-̈��ӄ]�����Sb=�{�1��55+6�|�Y�a��w�m���ײx,ϋ<�� 0������
��G�gc�I���G�O����K���t���|������Z=��圔>�U^;��f*3�_��T��3�{нO)���W`:�c�G�}L�-}����"��4ޖ����eE^�9�x�Ժ�{= f�U��85Ms{��vĻ�]b>���}_|�v���[I��Ȼ6��S�d�c�k�ٛrǺf�]R^F�}��룔Lu���&K�g[d��m��,߳N������mX�s*�n�Zs�$�_WX��
�n�T��^`��2�x�h��^��@��3Z�����6�It��}�}��{J�����a)�&Z}F��bU���% ���TV(���(����E�b1Q�,EX�,�("*�X�Y|����Qќ��Ֆ���.2�F۔��S��eDxnZ�Fo��@�]ҸN�`_g�o_p��JTwiw��J���dOA�gMŬɱA�.�]�5��e���[fy�)߼ �S�ﲺ�`,��[�:�'nv2�񬉙A�B[��'�/�{�
:���e1�u�F4qWj���;��K�X(1� E@X��B0�D`�D.�����f�87�e+��#)��b�7�ԇ6�3مsmR�ۣ�q�#ئq��e��,��Qy� 5�D�m�Z�3 &�9��jj���	�oט�L&�^�<�dmб�⬓w��G�P�BK�՗���w{y����w$��'Ԫt���u� ��N���/М�j�9�}���ЮꜧIA�}��Ak���)�t�#1���kh0{��ǫaþ�:R��D;���D�i�cq���#��7�mk��d{�o����owl�7�/{�	}�j����/%���h�Y��.M����ՍS�[A8�	�(� 2�A�n�w^�(��j��U���ow�䵻9�YI{��n��yU(��7����[�=�h�f��9_���FT\Y~%��������Ν�;�x딉���OoZҳl2��i��L!H1��-$��YV�
�"Ze{)�W+YH�TJ�P��5Fc��(�Te����\�K�\����*Z@KJ)
R�(a)�]���`�T�ނ� ������`q���7p͕���E-�����Ke�AhJIl��ݚCwNT�����V�Mi6r���9��=ì�`"�jB�]Q
V�e5E]@���-D�w�֗R��Mtj�-B�VJ�.�JJd��eBѲ���K�QF�H�iJÖhm����y�{U����AC;q�R�����6�Gc�6��s�l]���v�����ч�O ׇ��f�疫�4��]Z.��y��%����߹��[�(�O���^���3�n^�$�ʗ5ڦ��1"�u��n�*�j��Hp*E̩:���W�5Ŷ3���>��\~�-��J6�g>�6��m���IM�ǻ\v��p	��;��ٜJ��Lٔ�#䫨n� pZ�����yё����RX̘3)��V�/�J���*`�S�&>��N�<��=}�j�������F��Z�ʃ��7L��2�L�+�⺷�7��j�-��n��c;�؋��A�i#z����1[VO{�j���*¨��i)����� ��ݗ�@�O2�y��3Ws����
)>�]}�f���q�=��>�b��S�@�睷�Pe����мm��D)�&�$;��Lݪ�+fJ!<��	]�|�.���>U�>
��%wC[�7v�=����ԧ�IKC����k�]� ��'V�gqT)>�Ι�y{|�y��<�S�³�m�eV'�v�k��u������e�;� �tF�K3L헻����{����Pq	�z��h�Hu>Bm�i0a��$XChOj�}P�HE1�d��!��rM�ē��o}��˽�@u��Suo~�!�Y�su�l�x2H(K���C���I��ް6�S�'��	��ٔ+(!I8�!0��u����w�$ʠ�B~A@� ���?a�l�IHB�P��~v�����I���ܢ�Nk5��޷��i����Hq$�!&�J���?f�Hm�d�20��A@����I�HNf���U���\�$�!��P?0<�8��CYD8�ʢhm�������)8� E��/*i�	��O�"�fk+���b�e�bo�s��dVb��%���Vڙ	'�o_�	�[&�4�W�
h�[�I�]���1$�[�	8�*I�2�@-'��$� �-��>C��i�������/����o�g�7�4�)��0��'�>����I��P1$�<�0�g�18�2#ʁ����/��@<�_H��\]MO����k;�p� ]%��@�1Ip��Ҕ3���X��9�/��}<��X;�z���mW�E��C������1ny^��Qo�%>C�`�ʳ�ь>G���>�n�M@F�g��O3�Y�D��πʝ�\�fϾ�z>�"������f�!3ݫ�d���>��,|4�������GQ����cy���F����@�s�{""� ���y�DE�
1˞A�I���6`|
{ܯ2K���ޠ�Н�5�S�1}}����/ �ؗ�.����G�DU����(q�ݗ�T���VG��'�Gh���н���T2�F,�7
�k�s>� ��Bd��K�J�ۙp�PL��Q%	-ԩ�v�ʝ��1�e��Y�D�H"(�T��PX$��a`�( ���+b�5��0:8+.\��%��KJ������ ��gb�Ә��͵2ɔ�P4^2�z�;X�F̕�����z|��Um}��Dy��M��6�J蕣��.��v��UH��u�\o�q�]��,B���*e��Ax�J��~Z�����8������xe��n���(���5�j�"�T����4�!���*�
b�U
U  ����]��y}s@�]�x���f?/#�
8z��M���=NAɳn�EL��|g�B�fI�CL�̭�p� i��}$z">�;�9\��P;�_�oZ�bLh�����Bf�qk6�Xgx^����!{���~��ֽv�_�e˙~O��J�,��4e���wӫ���DD?_d!
����׷��ϴa�����-��X�KE@�����RQ��h�����e�    )�2@   $Ā$�  J�8��{y�s*okw���c̷c@��hEA�a��/x��<���C�F5aq+.MF�?�Z&�	N6����Z �|��(V�*�s� _����NI }��k}�9��ͯ2�x�oR&ona��.=B�q\����vN���x9����hI����!�:�Ğ##n�N��Ή����~V�z�A�f/�{���}�u���������U%XF���O��W�4+:�ҷ��-�:����	�lz�a5�-�m�Z-GF�ս�3w�_ky?%����޻\!:Ȉ��F
 �X�U�PU���,�E��+$b,�` )AD�go_}�׾��9}sl�ب��=�?y�y����~X�&bw�8�G�:N�{q�pz09����]f�W�40���8^X�B��t������{��l�}D(�.��ױ�^:��E�gv�q?wi�\����K�ÕXGw�O����9�g_����2�bfU�R�S��7qy;S}@�E
~*H��~�""�[��E���W���xʉ&��j��'=��$	$.f���5����S)l*����v�Wʇ�3���sG�+�_u�N(c���<�����:w+�^Ď�\�l(��k���^v�R��M�9t�E[ZE�D���y�mb�G�	WVk�ʬ�︱�5��5�_�>{���g�>�"G�{�ꏊ1��C�~�5�N��&m�)D�+y�w���c��b��J�9�OO�=�O����J��2����ϫ�������}�>����dU�X�"��aH����޳_}ʷ0��]���y��k_�Ŀ)����r���������n�x�fz{�y�G��q�9�)������R������'1֢_G�}�;97z�<�~�L��N�f��RhйO�T��b��&q��/ԡ��n᡺;�b��L�y����&E��x�ȸB��UY�O��*���bo$��u33�'?{���V�rcz��
���Q��T��z	��$�Q��	� �r��>��%��m�҇eP���-2J�`3$�>���9���ا��������Z�F�U�}�|#Y
��1\Ů�ެ�הMlX��� �ai<s��G�V�`�V�}P��H��R�U�w�	bFh���>|�8�|^#�;�~.�[�}�|숎�B�����V�����y��8�[�;��n"�w�s�*H��ԦY=�b�&eV�.�sz����I�V�P�!�p4^�1�.>��o����j��$(�+�*�m�n�bb2��b��^.��f�4�r6�d�vs4#S�)�r����[��˟_��9���)$ ��w_��������%�1=~�$�M9���wU���`���އB���m	�U�y��z��Q7ϑ����S>���s��Vj������ל�\�U$����c�}<�L��t���玚Wfk���%`_e��u�۹�^U��"%�0N��ׁ1�:���C��3|�]gΟ�˲f��ޭm��m��n)9+Φ<"݀f"e��@�YL��ut���;�r3���o�J��C�ޙ�֝)�_U�h���t�Y�K�G��|������"c�͔_	u�t7�8�ԙ�qYfǴv���}}��|º�wu�ޅ��ʤ��
1d���$l�u^ϴ�8/�!��ʂ#�ʸk�9MN8Ϛ������S�uH��O����uއ��W�}�VcZ.��Y�jj��]�.��%x�D=K�o�[~YT���9����h��u��K9��ҫ}E�C��������Ù&Ռ� �$d��7n�_��WM}���}�]��Cb(��*��A`'m��1It��������9�] ��=ۃ!�D��S��	�J�{~��J:�d[����)�R.�οG����'|�������%�D��r�GtҮ�����9k!��7�mdxT�ջ�Q��:��>��Z�+&tC'm}�Ђugkg�BúWD�v���-&�M����΀��"m�#I�	Q8���~7��=/��U����NӣS������ޮ���VB�&�6��؞p��%/<���{M1DD���ޯ!S.Kc��V�rR�gAw�w�"7I���(���"j��h3㝫�g<�NQ�4��P��Mh�����×^B���ψM�9���Ɂ1���F{����E�4w��j(���gY��?9�̑���&m��僭��u�?�G���nf��kn�]@�?DG�ݾ�Gۼ�W� A�\���[��b�c_#S�^�"-�
q��k���s�D8=��o��0��%c�WU�W�Մ��YH���DJ��m<-:��QY�T��E]fC�9���/���!c~7yU�?c�_�]�c���P XK���ǖ|	�)�TUA��UPX�U��)�E(�
�`�b�,D� Qd ���
�$0b����g�wy� L�  i$I  �B[ 	$  55�=�=�;�zn_ez���.�;��q��$��Np��}��Gٓ�n�q7��p`t�"L��(TW�\��l����T"i�
c��3���I4d<P�~�`;5-��	$%�:.���5y$�Y.2�%4�E�����:�'��,EQ<r���v��?^��}����WͶ���QO@^��_�}�Б�5�^�ݻ
=����*�|�$�������ޕ����n�f������]/%P�ʖ/��f���ԸF���}�u�vw�LtV�\d�33$���9>qD��Ů���G��:!+J ��tިԟ�<��F�^s�/��D{ՃӤ��ad��\}^�i��T�&�8v��\}�[�8�9�i��.Z��.Q���J2٢�_$qP�z��S��DB�{��
9��qH�r����z�`��S��Q�1}����;��rŘ�[����f�f��o�JM�i�7�i�-���À���q���E9��u9+/����f` �O���V�RHA�I��M��iR�2d������������!�1X�b0Q�� X��_=�ey��Y�z����;4���~���z����7���a��jcϝN�`��se�� O������>��O����m����(},!`�d�;�����Э�Pss���7�m�H��1��F\m�09�}�7�r�+0�T��1q�tc��.�ײ�)^��*M�������1T��_}�yz�c��w��9�χB��;�V.�	K�����൯��-�	��p�:N��֞��OJ;�12�gS�]�lx���#���f'�K"}��!u�G��GS��SJ�6%�����*����n�i���J}R�ٽ��!W��L������Yz��w��X`A,�LץO+��<ɹ���x���G��^�������
�5���Jq[e9Y2	�R7�j�.��r���J��/w=d��W��(R}��+�6tGÔ��+'OT����t*��?|E�~�W�~����I�o�f2fn� 0!���0�}2ˑ}�}w%����4g}}�q��m�o5}���`ؔu�]aݍ��}�N"�s9�J���PD���d��������e��3��+��Y>񏢄}��*H�f���>ɭS�f�+�6VIXw�Ö�:���+�T|�s'i��g8{2�	U'������M�cx�?k�;��K�Xg�mn�O;�7r0U
DD"�"@A�#E"�s[���DMz@]����r�m���|�Da���b�!L����$�,�
Ad"��
��t��>�w\2�Z��Yy:�q����I:�gW�r�u`C�kw �L;�{g���c���c��aW�ߏ<p~B�q=�8Ψa[aGן~��t�d���7���UeS,:�g����?gAwTն��ᛟ}��q�7�1�=���y�$��Y��ϩ���K�g�i��H>���L?m�84�ّ�H7�\c��S�ݑ��7nt���\������$&�͐����\�f���6�z�ܷ�|2�b	���L_��~�ʗz�<�ieԩ�g�Ӓ���8U�FQZ"��4w�^ e���R]h�����|���.O�V�֨��(�ܗ���P6v�s���M"z�T�|͗�=7cIGy�.�~��N�V�4s+��R)V�91�>gN.:���8l�н�o7&']��#ĝ������l�֚�z�O՚�^���	"*H�20� �� � ��WS"=�
��X=t�R���=�k�L�Ğ��E	�)Ot6	��ؚ^���RG���φg���6�@,���Y,�;��o�U|��&�Q�Y�mo�H�>���P��ג5��m��	췙�JZ�U=�;�E:~��Q���~� KT�Q)a(AdB��n����3��_U��޳6��۹l��FI}H�yݹ�\v�Y������d�zfuD�^�}S$�㾥y���:�G_T4�,��꺝&y%Nc���^�B7}���x.K_��������3~ni���	�C3^ّn[��j�Xx��R��B�o<��&��$�� ���K�$���1��k�Za�)��	�O�X}�"��5D����ע~ᴥ<`�</%/��x�C���;�̪���>�gޙq�a��{jr���ޘN�x��i'qahNݽH��M�/)����Ka��9���t��6�>%_��C2�}Mp�6d����u�>�x��{yO/�ɾv.�h�§�t�fkڕQ��s��
����I� 7Yr<g)Sѵ�C�.�gt��*��-��k: ��?�{��U_u�|A:S�G*S��1&�i2���a��׫��+�l���:�mwO����g;��*�@��fKܝN�.N�\�|�ΩQћw|%�P^ 1�
z����a�	�ȫ��T��EV$���e}��q���w3�Vg.�Gc�rs�ﾏ�����NZ5���y4�X��V[�衃��������(�:G��c�G���眃�*�2��V).���2��s��h��G6�:�h��#��f�(�uok�V;ޫ�/��0��2m(�# <{3+������j�R��aT+�X�s��%
uutAk��8@��R�|v�&P��yI+#���Y���x��m��?���&*�!&ᆦh���}��p��Ny��1�b�,�-cNT��NTL�G3Vˎ5Z�fe�:hL:�K�VR�WB�̘��J ��Ƙ�V��-l�q�V��HPÔVc�U�MU$��3e�(�AJ�өs(�*�+�����N��Rj薫]Q���o2�����%+��NZ;�J��T�f;���R����������TT��o*����U^�-�Jӯ�E��3҃��������0�A�rb#J?��<�Ǟ�is���!lv�g��=�R��<�"��E��=�'p�]���Y�U|�W}�9��]��s�����      �              	$$�L��3&D��BI$�	$ H      ��  $�$��   ��� �@    I 	$	$           �e;�+{����?;%��)E�K绱���o�p��;�0W�p��yi�X}z�|W���g|�}�ge֋Y�pWzJd��i�2���w�֗�*�(�Ùz����	!�+�Y��;3����+�zʡm[�xDM�s�w5��@M��R��\��ulw�(��`�j�r��{9;Ak�����S�������[��;�y�G6=��>͔r�E6��g�@{x��������"=�g�}w�����(h:����;joj������N���Sx�e�ˑt΂�^��ۛf-U4�B���u.yyg+\�;w�]'<��{2��)8�%Ή�?�z*�ʽ�O�+��E��>��f/"��W<p81vz�&d(�3%�'n���R��PV��9آV��i�s�nH�
�ClՓ�5����Tl���?&ʁM��1�N����e.�c̭?��d+Q�A@�z�FC���d�D�Rp9:����R}x�X�#ɆG����UI/tw0�d	����H�BH�m��!�^%�ݑ��5���p��&�1%u��jC"('!ƥ?"����S8ALI�B[{¹���t%<���T�ޙ
(�6*��	~T�!�9���*E|MY�Rʣk���ns�D(FY��%a�_9U,�Y���E�3r���=6
V)���Nl�^NE*8�c�Fu�'{�S� ��o� ���v�g�+���lI$� ,̉  $�$�   O�������k�o[�u~��]��<�����@�]�MEX�������=�71��$c�"�3A�0b�Ae@�Q��BRBG�Amz�eJ�Y52g��5���W{�/jUc��n4�Hl7���ğ�T�4p�8�3�^�T>�>T��]��F��x�!_�Y�(;�N�v�}�T�sk!��uyz�gW�J4O�U��D�D��>�ϊV϶M䵉U���9Z�C\f-�g>�[�a��T}�FR%�7n�.��봠ʀj{�%��VoO\�Ep��;�yܹu�@��׸��ۭA�j�NYg_l�1ԡ#���R>wW��D|j��>�LE�'^f�A"qs�ѣ��ڇ�T���"��n0W�ъ�ջ�JD��%�r&W^�KV�E��Q�b��=ddL쉏gI�_O���j�)�DH�D�a"{����.�v}}��z��(��k����=��KRѯ�Y]'��y��#H��hA=��p����V-�R���˜b~҅5��hkD'b��>�N�>��Y1���t[I&�m��~��w�6	�U�eJ�M�)2��jPp;�1^�P���xة��+���_n;����>�&2w��Y�O��Z��Z�S���n�~�>d��h75����"�G�}�N]g�����.�%�Ww����n��������(�JX��UQYV�v��X]J���.��YF���r4fw�iF�6��w�S���N�޺E���u���|g���{�ӺJ�Q�q��%�G�F`Y[i�� t�-��C���T�����8M4\�ض��K#��֞�ԯ�0�Jh_�^����Ǧ����sM׼��>�9f����=QZ�.�@C�ζ�hc��@�Z �����P��K�a]s�)�~4�w���ٸyD}���ã�q0yd7�o���/]:�-�;)(l�H��磻���P�̆{�1����ui��Ζ헦א��c��^��F
g�7B9�X�����dĽ���ƣV��Fe:0ov���o��/K�I��--Q���U1Wd�@)��S	4�ש@�ꕢ���0��:�ǫ��z0����[v��T����H�����o��&�����@�����/ɏU�p|��9���~)��7���"�-����z�{l��ٳ]��1�]$��W���l9g��zfw�x�ŕv��'r}�S}�8>3�ٸx�r*�Mu���Pp�o�K�{���)�K\�Еq�^t��Uܠ�5�@4
j*�T��y\zЭ�:�l��Ŏ�R�g=��]�����2#&z�^�43U5u�$'�5��+0�v�[���w�O�2�Ǻ�I���FDG�i���V_|7s�*��d�����Hܵ���|���h��ՠ6�c�hG{w�k��\��'F�b��U���L���b�O9��Z�"1v�8E�&�<�]!U���1M�E�g 4A�D�kv���p2�D��GN������ȮK�M˽�sW���U�CI�L�)�ށ�33/��F6Qg/Y����_����e�~��F*��@(��n����h�l��{�����ĝ���3�[�DX�9̈́×rse5-�n��oDx�D��;�Q��OK�S�9��t9k����V� ܄���Oo�����\v7�gY��ĸL��dd(6��V��9c�g����jUxwI���vU�.�n��*<�Q����͗	��~���w=NQ�5�8+Ϫ�C�����)n��>'ĩ#�nP?e¦��]+˵wP#]�I&�0c-����Lʅ�N+�h�w�iuF	�]?�޾������t|�PdQX��@EO�~�6mz}��fs�����Ը^f�fVEA�Jk��gBUKŷ�-��58��-�W��d-���e&(����-��k�Ɉ������&��F�CD�O�����]7���1��;�w���g3\��WK�\_@�9���ixl�X<PP�������ᶒM�ӂ*b�P��(*�$�e��m-;����z��Z����T��ou9�8�P`�K�[�ޤ�n��N�F��OKk���9�kt�2&���6�3ݛ1B��ޖ�	����!�fk��5������߮����"�|@F�gNϠK�d�x^.�����W���K�C�ꉘ���ꦱCqq�Ln��o���L��}7������w=�1Jwq�}�ت����I&�>�����������~��-���`S�y,DǒBl�a%`�^�6ټ��]{l<�0
�/�t�P�Ofù�W�Q��6oA]���@Ev��T�%�b�~�4/��֯O��D^��)��r�x��k"�hL�2���JҎ���r�Y��j����\�����Цj�{���R����UH�(�ZF� d��$(����=���+V�|�\yM�Q���1 ��>� �>�]���_���%s3z���u�� �@  $�  	$��̒@ �v��׽�ޅ6�>O��_X{���:�-�i�\;.,��;��;gh�5)��*�i���ZZeTL��������]��	�%GFL�Cp��_'b���j�4� �#q%$���]�ߦ��4ऋ$�(i9�B�;����R\efU@�P�m�M-@�ZeN|fژb�����qF�h��
  �{D��7�d�ENm�ʾ���g��f@�v G�����֋�E�y�p�wx{Q���8�u�P��ZI�U����d��1M�w�xr����k���.Mp�8�ON[�L�~V
;	��V1�G���cVB#"�d" ^}N�u�.���n�L��D����`eB�����<QHR�ʁ�5K^3}F����K��HC�c���OY�y��Q��V���1�({��չA��3]�Կ�s���Q,K�S*m~���F.�޹"]�zP�֥yܚf3;�������R����<�ޡ]��^bS����[�J����V���ػ�7�U���BG�o���^8�ݳ�J�[�;9�
�����zݭ�{��I6�m��}+ڐ��\!��p�[m$϶�9�a��>�R"{��>�����y�êl}�ي�iP�|���}�dĆe�{�z����S�0(O���&�c��.f�����*� �.�{Z�~w���Q�� |>cH�EK�DF��w+�F�[�,j����ܜڧ�ʳ9.K�Jtw�v��rB�c��2#�s�T��ͤ��-����ɞ������������w�LV���7�� V���7��I�w~���3���_�tWk[����RrJ�b�k���3�`�SYm�F'{m��`�=�ހ���	��ԡ��T��V<�4؆����i�Փ�@]!AW��]m�vF}C٬���ñ}NY̮����.��[Pt5V�=��*Ĺ�s�as��k*L�*����n����M���K��Z9P�����>���@w�ɥk5���#��tz7�D��qº
���,kUofv���5�um�X~F�*�,�&��q\Il ��1�r��Ix�0ffa�l��Ӕ>��IG� m�����SS�P#聡V��k��n��4��<����Nn��^WmnS��cf��ߤ4�>r��t�*R��.-(�FC�T��#u\DM�����@�|��}*s���T���3�$��xGO�4�]��nA��~[n�ewޣ�9�u$�_������T�q&cȪ��0�c~�0���P9�$_�87w�0�	gO�����i׮��*��� �$X@�[2̮n�R�{z�|��a�yk��:����#��a'_;y�u#��]i�.a0�<}5q	�h��j�,W����v~�o#9S��S���PSc1*�?{�O=�͹
o���>���Ǽ4����s=:#J"�
�1�YQ��p���3u}m��%�_�m�K���GN;�([� �I�s���U����]ӣ�j��|1!Nz%����D������`�j�;f�1R1<��a=��:�E����l����x��}7ۥ�o���I ���s�+u9zA��-�>0�D!ޏ��½tIil2���^�h~�tf{�>�aϔl�^���v�'x�OLS~�Zb@�n��ԭ;�%a����i�Q�]�+��v#�(�&�u*Y�}
q���Ћ�=��IU��,E��f�{�Y)=�����L8,���x��YMoyETo��	�9�т��s.���8Hg���<�"g���	�/)*�;���>�gG.<_Tk`@��S��3nz
�/άFfd�p�G�c2VjV�I����i#x+�]!�n�[^,ThhdyoB����9�~��>����k�WvߡEG�JUp�$`*���!�DP��E@R�RX�T����j��7Y����+M����3�1�ِ�оcl�����[��[�稒���&4���x�fV�9��D�	k��K��=AA�S�2Z��
�H��m��+.��X�L0������z)$�^��KD _�UK믖>y,����o����Y�9_�+������ ���v��7rߥ�p�2�a�Z�
�ךɊƧ3=㸾�%�����{ZCt?�>_~�b��g�^a��`�8lli�3�eG�#��B�>�y'�����3�Ę��0݌�k��c��*6����Og���\��3VW��V��a�J}K������o� ��Zsz����4��Ώ��tmL�S̃S�߳U�c�:�U���w�ļ�dM�ǳ�\JK�;�r^����������zfmF�i��̷ZW���P舋��Ѓ�#M�2_���؈z�5Afqmezf_\��\��|ɉ��LG�򺿸��xA~�-V�`�W�ߢ���5dş� �c��q�+�E��9������Ǿ�2)��[�[��NĜ�U-��^JG��=8!T���-���>��ڔ�0��@�@����ww�*�{u��59�fs�   Ēa$  �@��I  <���f�������~���2b��������V�;B�;�;^j�r�+.�(�v�VZү��FT�IBeL�5�7�3*�(����j
�G$mF�b~���3 W��^Md��V�*���L�f�)�m��T�N�{��>�*�f��X9���x��� z�xr��p��$���kw�s_T��7���(y�}t[L�\�v�����z�5{��M̈آa�5���IQś"��lw�離L����ir~�~x��8�4m�#����!�:O��kE紐$,^�2f�`�S�.Px��.��1�� ����_Xt�4zKK�wЫn5.o�*�^1�����&�����4���ɯ���]�c;l��HR��}���D`���Әw�K��wV$�Y!8���G��j(��~��<�L���jf�I���UQaGCw�<w��ل�	�ig���IW�����v�y�������Y�㛙U��q`m/\Ӝ Nr��[��w����6&�!��}���Im��M�c�(9ULȻJR�4H�4`nI�z�%j��#���M�}��37�Ьq{�ϽP��EI��w���Koo�ǳ����Eg�_̎�p����~���/�Y�B�y�T�G�*���4�e��Gd�}�4�����TR\6����Q�wb5��N�l��+e��$��NRqv��d^F��]�Q�*a>�ݛ����p�xT�z�m�ߝ��gӧ؟�貽��ޞ�ٚ�>�*�w���,�J����(	Z)���9Ii��M)V �������_�k�Nz�"��!?����~>���f��9Df��D#�]~GNI۵�km�̡�K���IoES��wE[Ez�%5����F�h&j��~�|��Y��*��/���n��B۽]�y�>�	�S��Ą�X�^��j�W��X-�U�x�G�ù9U
�Dc>��n��ܦin�|v<8��w�Bq��Ǐ�>��1Sl��i$۔�ޫ�$�-�f.N\�39�NQ^�X0]�S�j�1��:�e6�k�6)o5��Ɣ#�܎����1�[��q�hV
��>�N��K-��ڙE���B����P�g*á: ^^�^�zx��g)9dϱ�r}�V34���/�zF?���#׎�E�[Ȱe���re�&�_.v��k��.=�>�~w��H�"""��EW�<���~��kݽj� ����"��©��wCl�(��0�Ľ}2�	y��D�?�ޠ�b�X�<����㽸�x� �'�Sy��MA� �A��=%��P=%��Y��>����Lo�K�R��uQ��<�_"���!$��+�������2[��Ȇ�I��h�ݠ��`��v���	�%���ˋ����q�C�r��w��eïVl3�z:��qBq2]Z�jF`F�a�_Qs���#�+��R,��ʫ+.�3y�5-�4�e�uQ�˖YM�z�Vr�ww�ܥ��5i��S{+*�-�-��U�8q�H[��ۺ&s4[m���*3��ۭ$���*��(�j�ɽ�Gc9��+X���*��2��^٦Rr��ٛݎ�q�D�T��*���BM0$B���[p�u�딽Lh ��cx�*	�H H Q8�YvYwH�$r��2�؍��/Ti�eJ̹���oM��W7E�;�����C�_�]�I����f[W�12�CP��Zi��V���@ǟ��!��/��}O�Z(�SV5hQt1�i���'5\�s�}M9�]��w�$�G/EWm��d,��9%��:�o��}L�q��[�X�捛�aɞa�\�]�g�<}�/�k���;a�����<��EK�"xv�����+����7̅o��Pf6�,Ҽׯ{��jٗ�ڼ%fL��gd�2�[�-�|����ɷ��I�3m�6ۈ��;��\J��o�'a����Eψ#rIc�7+�E�}�.�]��sC*x+�v�����zN^�=�N��"��u}� %`������eD:��峺͖{H�^��oRj�М���*�9O5��Dћ+��&�:�ܥa���d��iV���s\����b�j��5��j�X��� !�c�AE󡖮L��}�@�Mf[��gN�5Ս&o�Q
�hh����&�Z}e�H7�	�뱼~�wd,&m2zl׽D��˂�(;D-,WsK����FV��VNo:����&��׮�*p��G0�dEJ !���f3}��dre��b6ݢy]��+��l����a�@jW�_�ז%<�o��])ɽ
M��Ga��c�ET&�#�7�ƽ\�$�٫���q(��<%���`'F����[it:ٿkq�6��_��*�x���C��Vmn˧v3H�A|z�fc�l�����jLQ��B<aƑiE�*����F�xp�6L��T-9��M�{�/Mܤ)G>̒=K��V�ĝ��S�5�s�߷�ճO��Z�s�܁��
" �Y�X��c�U}]�W����5`ߑQi%L��M�^$��M��yB�[R�P�Y3(����$������ƌ��b��K���w�o���*.8�ڝ.-)�g����;u�s���Pi��ϧ��Ī"���i�lB�@^�5����8;�=~��[�X�3�:�����P.N�^;�lFnɖ#����h�Q��|}�T/>�cU���Eg��$�	�6K)]+��K�W�h�p_�l�7G��8��S����{౉�yc��F5��f��k���ԉ��4�mX��ׯ���>3m-�=�o ���x�9m�s�c��w�3�z�����h��3v��v�_0 ��!��9��]rr
n��c{��^���n�t��A�#嚨īK���0Y[&����u��7\�mq^�v>��K	&C���yz��i���=B=��p�'5y�V��+>�y�Y�z;I�imt͈��hyoU~v�37����lD��ٵ�=��i$�I&��S3=�B�Lb���$A���T����<��D}P,J�N(�G-�r.�E���>z،������f�z�Ѕ�N[��� ��u�=�R'=A�f^̠eOrXc��YA{:�������Azu7����GE���1����(D�{*q}�}�+�Ao�ui�ꑯƅ�:�c�h*�>��FTf6���*�N!�՟{���0�y˾����l�k�K��۞��e�%���7��j=��}T���2>��՗P5�Cg�S�����եc�ZL!$��يEoB�{�Y��)*��n�r`����Q�vC���Mc����I &|~��̬��k�fx���t��XzWzj��Ȇ�U�>�cJ3��+��{ƫ��S�/��a�w��l��xgh�r�C�}��ij�G뫯�W��%��޿Ww���  	.�2@  �@�   k��+�fo�3��H�	f�}��UzAk��5�Ɩ�4���o��s�� U�x�A��O�z�B6	&B$��&� �L�!E'�X\���L*)��>[*�mWRFe�Sm���$���1!E\�s$Ai�m6[a����>���/V�eOo�Of�ӏ㸛EN<qS<�
�=Y��E=���u�*x������d���H1���٪�5t6H�:g�r��y�}8`s�Gi����� �]D�U�&OE�/<�E�i*-b��Dꙉp8�zN�l{K�u��*^l�eU�z��(rI�L�J�兑�x%3�;�Q�;�W�W�5�;�c'��5�#�z�yz����=���i��t�"����+���P�;��.�䚜V=��U���ݚ�`	���Qmp+/߯�{�p�I$�C_����n߳}�ϡ��8Xrg��7��d���=S��>˗,G���mՓ'�G��w���S�\�����Q�>�Vme�I����x���#bD^3�ʹKI$�oVC�EZj�[��_�KPz�K`�_5wa�!��5:.���W����y|ᝳ��	��l���^�ʤ�˺5��g޹:P�[N}�ط ��nk��؅��z��������g��9O7��1	!�$X7�~9��[�WJ���+��{��u��q_V�*o+�$!c���W �}[°��'V�jYT�h3��\�/$s�꜒(�����-F�g��]��,��C�v%k�}��*����KW�|Q)�Кf3=y/��3�D��E�C�n�h��=�IG��grv/Nz+��Y������C�*�8��b5{/X=��p�dJc�v����|��m��Ug=i�=����=���^�+��~2߸Vt�p��p�6t?�Q��xl��\�n�O�8���s0�m)<v�.��5g�^�����yH弝�*�uλ��|}��w<q�G:�C��Ŕk-d*����+Sau���l��m$�ex���IE/�)�SrP�"yY�������Xu�Y��)��6M�X�-0��9+��]���ܭu'�HB�$��~��y����W�����}qंU{keH�j7Ҹo5xf,>�סR��!�~k^�Ǘ٘���}t>�:u
0�5���7����=�D+W�$�Y���ٿ`��>�TǗ���J�U��ē̈́��ّT��߲���?]���E*��2�F�DQ��$Z�Eh�J
��H(
��"4T*(,(����P�`�*�TZ�(PQR�)+���Q�=�m�w����/��_i�E�B�����/��b�L�t��QEb�}Ǎ���[�9A�����>&���i�j;I���zX���y�~� g�CE��������'�m����ހ����eN�Z��EB�G� ^+����/g,��{m �$��v$V�Ǧ5[7�W��=o6e�(׼{�`̂DĈ�Bݪ�bH�Fi{��Ǘ����0��M�.�Џl1�;��Ř$��ְ��"+�|������� �u��u�\(Z	3fT˟L�Q�"�x�1D�=����(@��+j�O��l~�z�w
꘻\'^��G��61��1�>�q��x7�i�>�����i��uz$x��A:����ko�ne��$:�� ��@ȱ�@�}�{UGw;��x��/F��^���ѥ�"������w2�IϬ�f�M�.Է�Oi�h^�{Z۴�(�Ȉ��Q�+�2k=���Ι�4f}���jϾʙ0qs9�o/{#���6p2�S������Ҹc�f�oڕ\�BLRZ)�:g[��_�����|�T�ز�L>��
���G�B ��@�`B,�����|�_vj���<<H�Ň�q{�6y��#&�?.-bR-�i]�_b�t0�b���-�.�ujK:�u�W��
�@:'�W��F]�F�YV�U:�G�½�zꍅ�T�p1���fWh���v��qyHF.��)-��|����)�'򪲛rInF_ސ���J���ca0�C	8M�@�DO��K5�8��\��r-(�����AZ�b��jٵxD�������'g�
�}#N��<g��&�w)� �D��N_V�D{(
��0�5nl١V������n�T<v���io:��y�0��<9Nc1�����.�/!)Z6�w�gD��k������O߸A �� )b���72�J;鏢 �/�i;�~������	q�]��lt����N�C� �/PF&<@���p�ѳ��猿K=�O�J~y-��S���>��pF֨���~�ז�X�3��Jo��4̱(|s�<������2E�R�ܕ����/Cߔ�P�߱������ei��i����%;��G��/��u��Vw��UY[���sy���H��� �RU���d��@�G�A��xb,_��3X���d��$�H  I � 	$ �ޜ�\!�s-�(�|_����j̖�n`ԡ᪶���mB��5���TTH�$���G�*�q�<��4h$��_�V�u�" m�,�w��kBII���o3��fe]H���ny9�Ae�P�u� YrFu��C+�R�Z���1��I_���xT���WE<��e����6����T�MP�5�c�U����+9;�k��%�뛲�5||} �Y�1J'�aN�HE%��`k��[�"}}��P�u��	�Y�a ���w���/�>�J��"�-e�~���T�'E�Ö�UB%m%�dof=gYU���/�O�������r�$�o���m�A��Fo|D�����Y��'m�%>����DA�]��qآ�(��.���z'{]���0��K�t�y߸��Se���󎱣�޵�z��2Z�b��$��T�AB1H��F

������UW������g�h���7�g��(�	����bN�k7٫��f �L�_ī�J��-�L��m�N����i14�Ε������yULK����a�V/�ne1'�:��նaK�q��t����V��VZD�2"m�hҳM�+kE��/�/���v��cڪ���aLZj��s�sE����ѧ���[��u�b�;t��c��4��+�M�W���rg��]��f9!��kil^ �h�^V���!$'oy��{�{��;�g��>��������SX
h��s)�o*��i�E���Tx[�sf%*�����ur�ʆ6T{m&r�v��$(d�^�����H�������C^���x�x�����R��KA���O�/	��3>vm��~kqV�җUv�y��|�K2/Y�A��[�0��D'�@#3����g<:�W˃��a�:�u�����F�D_��w�A��n{�@�<.c�=yU����z�y�$ ��Zn𻼂���v2��EP��7�Y����T�W��6-e�G��o�9`��b,hܐ�nu�x@UO.�������+C;vHF@�K}	ɴ;f��/�eІ9j�.��}�EٌO���M"��#V��"=Q��1�6+p�I��L��ox��b�o��	����]�鎺�h��)������R��[��g|�ِV%�����n��k

���j�n���M^u*�vS��+��U�l�i�v$������B�&WX����P�p蓺�u�S��/��U���Lʞ�?N���r��[�F_�o�p|�ǖΣ�'�yB�����͕�W��ƛ\
;ׯ�+��0��t�)M�}��'7��s��5���4-Rn�#�A�9l�$��
�q�[A��1yXTKɟy����%/u�v@7�
����R��*.I��>�f�,�Ͻ|�I&�I&�Ra�
��)'��F�jH<�Gj ֡lǜ�O�l��F��Iٚ��ygnWU�]�-�Wt�Sߨxd<������t!}7])&�C3
�Dq߾�>/�8L���{O�*���$�����̳��u��@��@&aWpt�NT��e.Yb4xnv�O�ɜ��B��IU���=�E��ۛ���E�R�y�1�p�W���x��D$n�pE+L�ɴӒ棙����z༗X��c�7I�r�����"h�}���т�R�φ��{߯����%^�e�
#E�� A�$zLMHԜ�;�b+oN�B�*���\ڹ��ا�����`YΫ��� d�܆�32�U��-9�Q�V�Z;�=T�U_�Smj�D����TK�����vodG��ro"�C���R����I<]��}�.<�oa��vJ֕���I �j34��bV�2i��ʤ5I��H]yd�@z��
���F}�����D���؊�k���'+������Y��5f���@$Y#�8���Af�Vi�=�խ�B���=��Wڙ<��ǝ��K�k���_X�b��$d<H��W��J-҃�ss�����q��M��O���q�m����Yf��⾗3�j-��7c�p�yR_��`*����oC&+~=ǆ�Z�7���q�S�5��.�����̄�3l�~ֳ^�n�}����ު�GR��M�����GgN��}�8�I�䚀�]ו�t�����W�Mߺ�{;�$�l�c�?�<3AGozh�s�v�s0�����]c�`�"��+�D�ξ�&�z<�����Zh��x̢�%���rMa��a�N(_]���إ+��͹�/".��-q���
]�e^��\�L���䗊�ස�S�$�G�~�]Z�'y�.MvS5^�]U�t��en��G���#��9��ɏ�K�3�+��m/�pd�;`:
[��i�;`ӯ�	�m�\�3�V4A 3�ȶU(�������B��K�#�}EƪUA��M��MUJr��aT�1����1B�R����scb<j(����Zr�-��M4`V�E4�kXX�e�V�KJU��z�z�I�Tћ�hr����P��k-9t�%pwn����ReT��U4-!I)]\��7�yAH���c/IJ-{y�2�s���T�2���jm����-5Z�h�N�CV�c��ߤ���c�	 ,J	D�U�(PH�M_`�<e9wi��`�"m��0/+M1/G4�t/��E8o��^�h�=2(���H�      Yl�  I            ��y��2�"H�I@           L�f@�@   L�$�܀I    $�I ���@           ���})�.W�>S�yFn��2@��x�}r�Ɓ4#�
�"�\(�W/T�^U��X
3�՜o�e�鶍��,�Ls�������x������~��`���]b:�$۩$D�SM��%+u~��ƻ��{��J5��]W�.m�{Lǻ�b�zԙ�:� 猚�O��M�ʙ�g��lV���3�o�w��0\qyMd�s��W%�=
b q��j^e��]=�c89���Ǩ�F�M�|�dֵ��q,�a<7��&� B�ߡ�P}��bt��PN��/v����Z��>���a���~����Q��p@��m)�BWC_R��>�z��3����B���7�!a��y�:'&:�O����c2��u}0���3e���fE�vL<"ϼ�4G30zMBKn�Ox�+V�������K�ڴ��큖��s3;)[�>��Τ��u)=E�Uh�mF0���2�����X��ό��Ć�4�*�)��F��ImR�rT(��`��*-4�Xũi6hD5T�^b
2�gU/1���]$�I-�n�e!?�!��DXB,M���"L�*�O�5#{e2��NhiyF��p�.v�´�08p��MoW0�-����/���(,:Ϣ�n���5��A@�A�[�BLl�T�`D�{F�˧�qN�Z��aL�O�n�s�a�������˄~9�m1�L�#����j�3   I��   ��I ��g ����}�s3e�����s�}O�2�%��o��fu�zxI���]���x�ѥ�}�윰eٖD�ь��M$���m�u�۔Q���SDSlL�ȲIRH�rM�i�VPB�*J5Fy+,�E�WP��?���/i����l��p ��C1|�"&����q]s?}8NPۢd:}ƝB�=Ҿ�8]eWI�m��xW]��c�.̻h��jՖ#=��ȳ=T�C���*����>��]��D��|�]t?wY=�z�h�2��7ƨbhD�汬m(��y�Wr\"�G�u}g���L;wͷ��k4���X�DW�}�yEþŮ���EȚޔ#�}��JⲔ�h�sӂ|�]GX�d�?1R|qC=�}\�Ŧ��z���Vxݳ_|i']$B>A�-�[�Q���=��ǔ�-����)]�伃��x�����P�-�uS�_j1s��
o�������>a"I�Y{�ɣ�2��H�Ű�p��_��8>>���E�\I��T�x��sd�a�4qgq6#��"Ȅ!�r�ۏ;R];9���M$
�_)�qI��ic^�>����>���Ă�c�u��n�$kk.0܁���׷��kQ�Ck��=,���k���+�g9PA��c��oot���zt��Q[��Gg/q���_�̰󺌫2�6�[�;u�bE���Ȇ�[����GF{\^��>�'������.��~���
(��� >;RC��s
����{�y=]�Y��6���1T���D
��D�K���/&}t��PW�Dt�����؏<�1H����Cmh�r��}�:nN�9佺��{OEU��^�`���θ�ʃ;1��vv\�����%؛6kq8���.L2��JuvLOYO۩���r"��xou��DG��1�Ci�ܑ��0cp�$��dIHu�0{|3������6lQ�1ؘ\��C�DK9)R���Y��4vF�NuO%ˍ@8��c,aQ莪�6�*���Qt 겹R���l'�<3h=��R�[��0lY�P�Ӄ��F��V|��O��H�����o�Q[и����o�H��C�����y�&��ړ�U��/�����fQ�}�w�=%� �1!V*���#���v$�d�[|��im�΢v�JʽQ�D�e@d��HC��"z����Tc9�~^�Քҏ
������<ݞ�k�w���D��i����:fF�*0�¼�ԋ�~��/��w�X#l��ްu�st�0��]��5k�F��Ƭ���B'�d�8y���S�v���4">� q��q�����D���"Ͼ����}���(��D�~���MS�z�@
�����3 '�SU�k�3[��cP�H�Zh/%x���4l�LV�F,FU��cz!�e����}lvU���{��jz��P���ՑV��'L?f����=$wk�5��</���U`K�g��r�l�/ �}�����)�WT��i�Ѯ{;�~7i:2AAa���Wg皯���L�`�Ӫϻ�V�˷�x��eپz�s�������V-J �{j��ˊ��<�s��7*�91u�z��>Wx_۠E� ���fc`�u5s��xXf��Qq��ư�T�mzs�ϯ+;�60�Y"Ed` #U!EQku��/��Y�^{���E�v<��Ī=��z{�o-A��fu�RΎ����b���ɳ��9��b6�n�{�e5�)��a���#���@'�q	ш�$��^�T}�������[�`B�-SX�2����NQS��Xmʌ�A{����m�N�(S2�4
�Q�����?�c�g��������v�"��+��W����k?z�c�8���>b2V�=%;4�=$re��S�_C�gLo(�0G�}�����З�J�{�g~�׫�������{$��k��쾞��>|M%�#��h�N�X<�)��g��kLˑR>#(�1�/�'wά�~�ǈş�#6���&+0mt-��bի�m�O�i�e���m9�K�T]�%AM�S�Y�Knv;�[?Q�lw�������O޻����wr�@�������" ��1O%�=^��S4�7�`�~�%�~PU����iʕ쎱P�ʼ8 C;eޫHa�X][|�z�{=�z?����?V��Dd�$�!����oƸ�����\ �  WrH    �@   
{������k�&]�u�����
��]펝)s9���ƛ�$e��H����]� ��	|�v�!�`���M�R��T���+꾀�T�kSWz�fT]���\Ӂ$�P5C���!4#��-��/�џ&�9��>ebxjc�+�a�ޝ��ޘ�`�^�׵�������D�9�/���Uk��-.&]��h�3*���������G�Ccfq�cֳfwb��q�#����Y�EfR�Ŏ�t5mgq�]�'x�>�V�U�i�0��6B�@�;mr�Q��U�p��E�fR�vE�CӍ �QF.�x�Yh�� �u$������[�_��^T�P���dJ=~�op����c;G��j�_���}�L�,�C���n�5��^3$I����P9Gݦ��u��d�R�����i�8���ь�{���?@����L��'Y��?SI-�V���s*^�$Ĕ�K�eH_9���:��଄��M�?�;��ƴ�"�F�d�(1���y�`��-_=�,�-�Ӈ���� Ab0��/���/�[�H�t��l8��I��X]�G��j�>_��+[����$4�T,ib�"�
0d���B���EǍ��~1o}淽]Ӭە���z��=��y#����XO���L�۹������ޣ��[珻)Z}�F?~�����A��2j�no�{}��=�c�<�w���h�؋|7�+�t�<Y��r�^�^�Z(&S�A'��9PGP6({�nW1,������%��������w}3法�g$��~������g�]O�����JªT����Q�֌��2�L���~�
��c��GUq��&�ʥX'��"D%˗��uC"9-�����sY�Z���Q�(�)tRR8]�GF��?E��51fG��� /�s�U��s)W�s/�e�e��Z��߉�Q<c��X��&�<W��!��٦]}?��!���g�]�խ�[���8��DKΓZz��`��ݕp��6�qW^S���2��;u�Ǥ��}���.�g�a���Ǭ@;X�9�4A�1�������Q�iD� ����s�8"��u�7���w,�����������5���z���Ô44S� I��s`E���U��7�v]}�E�%%ܮl��&5��q5�X1��^T�o�]���u�̓�.��պ��wm?��&�l�| ��g�y����FR��m@���RD����Fq��)T�eƩ�oe��`&��x�ɷ ��d�J%�������b�wr������wЗ��/�λӰ�N�˰�xl��K3Wݮ�_>�?q�A�J���~E8b'v#��m�m�'0��٫�e�l�V�q!�F��o�D�C�S�����}Q�8#��rs��1�rc�e�L���`ucѝ*���WW�faM����wd3jי���%�E]�|�m�_ug��o���KE�f���]xj�0�ll�{�� �C25�����>�&�K�V����׀EM���X��͑�35C�q��r�הh��(B
	�o\�����ek���Y��#K��au�V"�_�	�f��䰺; �U"tD�Q�5�ؓ��#�^�4����*hRV��<�яĚΧ}z�qE��l����5����y���}^��}�����Gy>����BΡS�P����8�*��.:A�^����V����a�����DJ��J,,U��8^`[�/	m���(]����e���X�B6�F��	�f���!W���Dh��#��{�d��%$����y�M�0�r��Ql����]X/�X!io�ė��x��8#d���m^�o%�u�|��ڎ9p�
����DO�-ӝw�U$���q�򋮑N��,��T9*U���FQ��qey��}�+t����Ykя��6mEP�zI�$|����l��"�]���i|���=�1��B����u:�7�DA��{��x1����q�w.�Yέ�:��S�'���rͶ4xo'݊&Jt�.J�x҂K8w�r��Y�]e_@?Lu��޶}�q+&�q���AB��Y^�a����U21���7�.������,��⯊ܹ��9�{Q˼?3�)����Q���s��?;4��n�ҹ�׍��nͰ�2�S
k���ӿ;��/W�d�$f  +� f   $� ��r�=+]�����1��E�4������&.�l>{!���=�ۈN�@{yslX P#���E7��*[c $��r������$$�|��j��d8q�Ꙏ�RI$����H�7<D����ld��cc��"j�t�d}Q]�;8�s-'ד�+D@S7&����"�8>��N��5����0<��8�5�e��>`tN+9>���]FǪ���n/l�Yza�`"��[������}�0v���p�~����h.a�+�^G�qP�tl�x�b��5�b���թqGw]$�l�H� FU�6k/p���L��0j�çB�S��u=ETڝ�����P�7�لO��$1#5�k�.4��K��,�6C�EĞ��ϴ��d���ܺ�M�
��y���"� ��UZ/�&#��^�*��U��x�.}G�g���͘�#��>�8#�f��m$�m��4�%MBCI�*Xi��`&'Ɔ�Z�z� �V*o�\�b���{����L8S���0.6$�;րx�����S���V�U�M$�Eϔc.�{��x#�=M�� |LH����U@��h�֏�[Zߵ�WKnu=��i�e]�]ʵr��`�M�����7C�ϛP�e��������ճWf!zq���7���sڽ��
ȣ 
#]�^>�����h��p�lm�n�����C�.�&�'P�����/��Tyڀ�q�
�Sw�)�蔓ϼ�X�F����nV�l��O� a�]K�Bl���ڱ�h�8��#�/)��-Pke�t/
�dF��מ3J������k�j��bx�~| 7����Ώ~Q�t�<]��[�z �w��n�ڇ8��h-y�;7ĕ
'����O��NsI��m��J�QqbL�9�Bh!-�&�L��-��D{��m�KB�4�q��x��~����|�\����@Ns�:�PcVRc�33��T�%URH�	Tq�"�f��C���f�u�/U��G�Nӹ�(���b,N�WButߏ�)_=�*DM�:E|�L�A��j��������!�R&v��J��|�D3(u(�G]�A D�P��yY���L�g��n8Io��5�7�y;�Y���&/o������u�`B���f)ffp�%������2�i�͎ثg���C6!�7���S�/r��M]u��&��q���N�⠭f���u3����\ `�/Oj��Y�h5o��7�0JS�9���n�~�L#]��b�iQCզY��:�$*!�Jˡ�9�hpa@���XV�&Y�Ѡ��Q���Xo�#
�NR���e�.��֨P�+�ì�S%%�iM"�HX/RVn64o��C���l�Vq�*5O.�YM���b+Ϝ�4h�սo�Y-�p�a¾a[�
Xƪ����&��s-��n�[�Ň�=�_a@Hᾄ��!� �ڳq�5��d}0٩����oϝ�3᷷�g��h�*yP�P��-��eU���B!�{�WFXo&�N�CX��'�
��1}�F���t����6{Ӝp<+����%f���;7Hn#�c�)ca���%�^�ϕ}��c���Lü%�g3���4Z�iP�7i�̓_Do�I�m[voigh7�.�ĖU+MY�-
ά�0t�WaĴ�l�Q��3&͊a���<p�����oݵ0k��޼_�	_	|��n���.ŏ/-NZn��5H����2u��Ժ��ͷ��Rmn�3GP�m�Z��=Б��=|N)��
`sL����&R٥Kɤ�cܳ�.vK�����f�-Z�Ls&�Y+&.�,�,d���]Ab�̈�{�h���[��k�%�|bS<��+O�JHM�9Fk����x�ӽ�vF��d�/w7i���8�4V���N�ڀ��b
먯�>w���]��fp+=�T� �_x�2��ܵ����
�<�T���܈_a��6�ܺ�h�(�W��[B�ov�EC4��ǻ���'1M��9;����z���f�s=1'Vͪ[�zKA�����:���e!�(�����q�͊(#}�C\z�a���A�+U��<�7�#$f�/�/n
uF^����FW�@���Ge��sԸyG�� ��^�F�w�Ւ7��q5O9T��֨��A���щr�y,p�G�Jp/�:@���y��>/J���u6�, s�V��W����W��V�]d�Vnj&��#���*�Uu/��E6�<K��ٻ%r�2S�6�~[p��,�;6^��y{�����i���G��@P��W�޵�ߵ�;��W~ޫEH|�o*42�'}�ob�*+XR�r��j����OR|�ﻲ�h�Ga.��Un�n!J1C}��c��0bn�P�H��#��O��gn����M� z�[���oV�e䰽��%�8�*dއ�<؏��Z��k��p���&����DC�pQ�uڡ��{������m�s������5F SHC��u꿹��6�a{4�r��w9JR�[w����(�l,�� N=4m˼����(x�ͅ���Dnּ���Ź���M���dfk�َZ�huS"',�F��9Ƒ3N�5芛g'U�]�
��U !gb�w
��̮��Km��{�����(h���́�-��T�H����tQr��t�����8�1:���ݘ�m�DF�s������
�i��?x���;��P�S'kH���$�:h7G��A3c26vzb�ë��9'0��8��E�#���K=��K�C}Y�ga<n=j���flE��@����a��5Ԥ0wB�$�UD���9��y)c&�"T"��M
S7�-D	�k0��uK��5�
">v����<฽>��J�-�j��& ��}	şUL��/��.�|2�����M�u�w!/��ّ�dWLU$o���4s���k�P���羕1�b�3�M����0D1���0��JU���N9����p�������o�ͯE��4	P�"("��P���H��F���R	T�QHUR�R��4 �UuwW�I���[ߵ���@�  3 H�	$$��   ��g[�7_W�v��f���o��i��y"}��Mx����_��������[&�v_��5֊��2D�jD�j(�q)s$�����%�%����G윔���W5[f �&Mrk�3F��K��r�Ak�K���־�%$�
�QV���n�t5壙�a��U�M$�kc�m¼uճ9�Z&�T��6�6��X�?m�E1M�|ȇ{�=}#t�L}XbÒ���&w����#��+7�O����Vo��3$���i.r�l��L'!j��l6�BjT(5�x ~L^�Bڀ�<J�Vj~�A��}��u���F,�B�O��f�*VpF�Q�ـ��\j�Nirt�����uW��}k�ƨ�  ��Oqpܫ�ث:�kv�i�z��Ͳ���F}7=v�bO��+�yw�M��/nx���p����W�1�@V�M�-�]u/��}��տ^�ػ fk�u\�ZM&�a�!\�̣0���|��Q=�|dMj�.|�R-�ӷ�.3Ψ��hF"0��n�Ѹ�5�}�8hP�^�;��aX�n�CHe�71)��}�ɉ�>�y��{y^�����IhEXBE
H��Y���w�8�^��o\��y-oQOjDM:����;��;.>��J�Nnշs~KPd벮k��[��ҟ��>wg7\h5QS��{�xV�g�}ۆ9 ��q�p���^#`@���Hu.}\���Ĺ���p���Q��ʪ6mH�1)	�#G���:�(2�on��c.�/9�������D]�c4.L����	gd��l]�6%��R��&3��ӔX��\�-�w�ႃ�^{O�J�ˠ�/���|�!��9X�'5X��N�.�`�:�������y�U/k�yg���M���� j��kY�&��j�c&K[d�䶎Ł$�@db��%��F���]�� H�{�TN,��|8կ�P;�n����
�n�t�~ۜ�m����]���z��k���Xy2P�Nͱ'[ڬt#�PN����9��5��^û�Y����ĝGt��UW������浬���z��7�~��}�7FAT�RAAH,�"��o��k�[E�W
v�u=OIz�_t�p<���-r�}w�)c���ݱEs�>�Y��J�_���,|]����5Y�-CDݭ_��Wq���Z���{җ�z���6��˔fs� ׈A�*���.�J��� �+X4S��[;ِj�@����|���V���	��)�j���3������S�Cq�3��  ��V�k[�6U�K��]8%&aK�s7�ǣs�� �EV�ϖ]����<�ܽ

��~f6ͬk�顑�K���0�y���kBj.'sC���w��J��L��������1�} <��b�<^�nX&&��pbQ�7�i9Zi�v{z���Չ<�Y�zY��}3v���BA'�l�V}��K~�ZUÙpߜ�'PB��ٴ018mfx�sں���kz�.U)L�Ej���W��v�o��@��\ݩ(uerV!�X�w���/�y��d�Ͼ�W�8�8>ǲ������7\�:-�i�|��f�u�Z=�����E	��.�w�+�)��e�U�'�=5Q5*R��뺇޼횊���"��Ii�m����+nD�$끠�[�7 �}s�=���*=���Ҁ�e�p�j���;��pw웇S�������b��iL�����SZ��o7�|��;�.�I�*�`�����0Y"�0b3��Bp|w�k���s3�/���zx� �\�-'���,�w�����U&u����B�վC��l{�߶�a�j����3D(�Tnh��Q��X��y��¢{qV[�#�uh��]TV9 z=~�}}�}
�T�h���D�"��;ӫ��Nc���bp9H�Ȥ26�|��̨熣���[�Q�%�ab�}w=y?>�=��US���s�m��   ˙    �    _�9��	��`䶁L�'�Պ��g�k�֎D`����̖iԑ{��+�AAJ8�	�Y�9z�Ƙ������K�N��cu��)iS�"��w
��d��#m�$B�-	�-jL�����f�%9(]]󽉻�oEE�]|��^?pև[<x�2�Ӕ#����������y�ƾ�ܿ00��{���.���}�Hɴ2b�cҴ�P�SU�f ;���&���z�Cܳ�&��[�&��P�����hA����y��+�~���UY��G���-���2���/�,A�v �J�S����LwNgs��DW��{3{�q�B��m��w�d���%�rݔR3*�3�
�e;ѝ�ԋ��ȷzmBʭ�ɭ�k�5�}�]�n[��I6��8��.(�ZmÀX!�ų2T�K���}6K�w= q�H�c�'���W��T,�88��ʼ�������?"�Xo�,������s�;5�`���H��~ �Sˋj�5����5���o��V��J�=m�i<ds�=�Y݁�#�Om�: �HlݱöX#��v��\�;�zxR�ܪ0\l�V��lA��#�Mdz�����cr1�WojgY�kY�r�ƶe��$�3ٻA�t�r�uUU��9���E�l����{d�����o�wI��
�S��+l���Q��[p4��b{�g�ݳ��(Vw�ǉ*WP�+����|��'�/\���=����$� 
���0�A�a���pe�xOv���.���3~f?��)_T*����f�=Zk��KԂ�Ql\��p,�;f�G��Me�w*NC�ry>�\LX�t��j����8��P��t�Mp�Y���˪prW=ډ�먎{�>��v�5g�@�9}��(�P��E��j��h����b��ת�*�!VT���i!:e���W�W{���ʃ2"q��N]5V�c�;� ڏ��������;꽗p�tG�}�4�ξ�zQ��e�g�4�G�xx��D�A���\��E�O+}*t��sܫl�iڸ��Yk�����J4�H�gst�
�nV	���Ղ�5^��vi�+���ԇV���9�~��I$N6ےH?)MM�K�Ru��`�VU��A�1F���>��|����ʣ���ە<<V{\M���c���U�2��C}�ϧw� �\ʥ��R��T�o�u���	7I:��ӄY&���k�Ȧ���S��k���{I6y����9vF��| '��*��#�n��x�o>�g�"��z��2�Y}����fs�+ch)l�J�-� 륎w���Ý��*��H�@���}X��nPl�;â����T�4�Vͮ&{�����R�z�BiԜ�3Ө&���!\����Co��2-��Gt[��՘��t����y��3
��x�������>���x\}�K��m�ے?!)+%�J���.��i�,��7 �ՓG"�:!1�^U% �@Xh���.w%��\��M0�(,�|#`��VD��(dR��{�u�8�K|,]Dߩ.Y�$�s�[�Q�)Y�B3���O������[�9�B>�b�����.=c�2���嗵�]�W�wy�Y������bN홢a3=Pݳz'���v%��6+����3U���c;���w}QSp5��l��#z؝�vBg>9 r�ӿV���7����B��+��@L�,��>��&!�W��]�<i�1�p�7�!.����S��w�˦,�W�Hx��ޒ#��Ӯ.��w{�ո�թ���$8R]��x�4�ٜ�fq��p��XV���.�ߜ\uuЍ��TM�	2DK@���,O��"��S,a��g������p��R�0�UL���G{�y�B���PB�x�h�DO��� ?"d�oJ7x�i��R�)np�>���6�I
�Y�HdS���wdn��[d�,�oWV�Т˪�]Y*�4��P���
���F�z�*�(u��A�eYyR�X�%�۫JYM�[��QE�Z���TPV"��Ԫ�ں�ye�)%�IT[u��[5�.��cK
.�EA��2K���ۥ����Eu�z�wx���S�yH�Jn�YUCUv.5�L���T����	�$vA�������EQզ����UV��JS�&�3E��\���ix\��`KeYG��
�j�����ԇcZyem2 F��PXYT	���s��r`�X���qV���L��f�c��}���y����
kJ�S�b7J=�6�x�ڏ�=>�V�5�w�n��*�H�����1]�/�������_�{Z�pѤ�<���oV������^�+�~�      �� HI       H    ��fFd�s$��A$�I �         ,H	$   $��	��        ���@           �W<ǹ������������W�mn:Z�7��g��6�)�?Q2P��h��bY1�j�cKp�,�C��#f�{4ru�<���{;} ���k���iVI%�:>��MrJ����ky$��QҝX]�=�*v���Ʊj�]$��Q���@��S}�TI��eT��
���9ͻ록����D�vXx9�i���o��Ѻ�{+to+T"AǸ"��L��Bގӷ�"N�� �\EZ�Ia�
jFx��Hن��^蕱h����%�Ky�#��T�Jp�-�&u�+uJu��ɒ���.��ӥw�d�5�6���W���䣲����z���Fo���i�]�ݡ0��˧�>}{|�#���A��6�1�,�>w:�U��MM�R	�G���Yp�d�q��Ԟ{=�e3I�]T	�:ǂ�}�4�އ�;'p�]9�7%3X�eP�^�\�t���}A�c���OjiI�)S���Yנ׌�������ͅ�K>~�5�1h|�&~�p��e8��}�jY�=�x�DIk�~�OH�ڄح4��l����I*4DԨ��K-�aBSB�^=�x5������7��wHTKj�]����4��V9t�:�5�I66�>�.6�Ȫ�2CV[�3>0�1�W��u0���ނ�q'yz�ǫ���I�������?B��:��.��1^���{rE�e���r��2�����Vj��W�.p3  //   ��@H  �y�ou�ggk���~�^F�q(n�Zf1`�o���-!��H�{Dx�l�j	6"~�j��h4L�-`�q��P��!)�,�!���M�!C����;n���f �V�7��Sr�a�TN(�-���Ǳwl�yt���n�I�#`�̛�T��RCG�S��/Z�s.;ٖ��>P.�dP{�&6�����?o]����l�^�/�釻~�,V ��"0���WTڽ�����<���r��=v�vqu�N�U:2��Y���z������-Ӕ�9��j�z�ʇ���˗�����6'Z\��@٧�m�<�[�1���6�Ҋ�X�$��Ѽ��;��ﾉ��\a�7���WM2�\�{��j��V�k_I�$ �5��p�
țp��p�l�K�������p�w�h�C�5Ҥ��ySK��T�o3H�ɕ�DTJ�e5g����������b7_{m�����i��P�Ȋ��QH�dYaI
V
�UTQ�@X,P�Q%0UY�1����P/�絲 w�Mh�J)��wu������Av�}+uI1 8�ꭝHG�$���F[�!�ژ�֚��S��}�ѧei��b3NJ�����+�ɷM�M&�VZۮ5B�%=�鴱w]��	%)��co����0v��4_EQ�I6�leC&]Jf�St��K���ޱR{/1wc��^�sz�۪��H)$Fn��S�������,
�7��uHJt+��י��E��ze�m��d�_���j��e�h���	����5�����o+9�e��\&KE%b��ڳ����+�i������2�$L,Y��R*ڂ�8f�#Z��n�]|�^/�I}�@'�|;�v�y�'#���Q�d�OXOOEw7��J�b쳴�e<����}��r"�_����+:sܫ޽��A@"�;f9d����v聽�=�e�������}%t��;�l�,����v��3����6r�.⑺��E��\���(�|⳶����~�菗�B�C�J&�WަeG�e-ޗ�"�f�ʌ���<��H?6�|=�Q�˦0��p�[�a%�w@I�r�%{r�p!>�!B���ț���),]"�΍�f�Ӂ7�+�e�M���¥_R�<fZs+o�ԫo��ј4����2�V�R�F\��X�Ζ�=��n���+Mv�:I�L���-�ئ��0�=�'�{�W㵑�Ō��)<�t�g�������k쮜R�8̸o2�ه=�>T������]�������XQʊ�g�-��}N�w�]"(��$AH�AT�d�E�a{�^�Wyv�7��u�v��գ;��I�';��[ T�Dے�lgx��,@*�Y��ٖ�u销i�_T��'�	�ӛml!����ܕ��l�&��z�:L朝�GB:��=�kw�$�� R�w|��5�sp� (g&�)�[eU���{��Ój�XC0�k�W�W�V]�����#�#�/������m�$�Ny�*Ww��6��K���j������Tz�W����,�eA,���a�IM����6'4t)ǫ޻�6�6�����t�0�ޓbr�To�E�>��l ��)�n�N������o�kOkf�_o]@�����iG�n2��?P<L��yO�U��lQv�q\k�[4�%2t]`Ǥ�oV�
_�g{v 3;�˰Ԯ4����^�
��	��O~���ޒI$m�$  2�&d    �@  +ݍee��* CʱV���%�W����~���==f��fL�L9�FV0�&d�l'J�q�{ȉk����@r��L�C���JD�ŋ��"Ʋ��f��[��M�$�$���u��������a
"�m�)��ԧw?_Ԛ���ih�j����Z̖�%�gi�Rp!�3��d���ӧ%YXv�w\���x�]������R�d�~�R�:}��J��)Q�g0qq�k�]D|@�?olP�ܳ�",o�zϢ�a�D�l��(կ�<�o��SU��,-�N#LlK�A��o9)�Ew%�jj����N\���ڴOm8.�к� �Ք�O�%,`��J{s��ݹ˯���ک$Y=�t�����y�� L�R�.kB�˵�ԊSM�71,.*��jsb3sqצjʔ�T2k`�Gn���xG:��h�7B:V���B��.�U0�+'S�P&R��s<��:ƹ꯫��8����˴t�i��*DUu>욂w��w$��0���$�o�=�����������>��+WR5wX�#2{k�����D'[�Dty_N�;G}�;9OWY�G�0�p��
��[�3��RCz1�|���頹��3T�(��)\����G=/�9;+��T$Rk@.����d����_v#�!q;��+'��q�C������������hOkjc[<ߛnInH��?�j&`�|B.��Vg<Y�_���>�ێ Y]�Irf-�4����}��[FjM.���q'XgQ��tj9TH\[��FrnP�������y��ȳI�Zq_}̨�VC7���z��YS��בhZ��-:�5X(�B?^�g(���>>�9�w���{uwsę����0�s�»h��ͼ<�ݮi�
��Z���sV���iO/2m����3�]��*_x�\v=���ŭ�� sJ�J��sW�WQ\�#O쿷�G|ϸ�>��<�-�@ӕ}�=j����
�����s�	F]������Ƶ]��w���8��d",�BЌM`�& HF�RI$s�oH����U���K�q�Y���s�(?c�o���x��y�~}E�*��1�t"�OFI��k\6*�ƥ�]�j���6�����Wۣ;Q�]n2�]�
���r�)�q�^Gq�$x�B k	�w�����1l���k�
��l�Qx�=�1�ny�!�n���3�[��9�A�L��p��Vͧ~�՛��R[R("�x�
V�
�"���b��+I �A~�����3kuɢ7@f�6ާ\ۜ�t����Q�s�[3��}r��Vך�g�^6yf�Ǿ�Q̟Y��Ż��jg8L��֪i���j|� ��p;���rǐ�������Wi�g�b����,����M�M��"�ɇpRpdL9#�k79�1��-����f�NY�������������8�e{�+�`�Sy�κ�ѽkT!�=$��U�^�� )���ϒ�1�@)�/�+���3U&�+>�����.��}�8����'�-u藞�P�2�fG=J�e�˃��3Ҷ��NyGw
9ծ�\�zY��U��;�$Ȩhɥ�  �("��" 1�;^��=��A�*Uf[�.�mw<ӕ)^f��7[׳]yR���ټ"ծ�X�;vC'��x����{�O{�I@�ew{�y�g�$�  	$    HfI  op�n�]jT���ܙ}�}ڄ��\F����ԓ\8�f��J��6���V:�sg ��+��G�
%i���j>cJ6�GN*�	P��:����	/�z��$r@ ������T�ܬ���VJl��g&N�`ڲ_n"��@[�:�!;�*u2r��6�I��d���U|.��l�U�,�K��v]ir���X�\�N����ǨA	a,KB��=~�}�V(u�3{�^���<N����B	���Y���>�}�p.�K���۸0��!4y�Վ������=UVp�5=�}���Q��C��H~]o�� �Q�r�J�c��L��Q�{"��F�jĢ��#8Q�TW���=+L���6+���??]�$���WI�b8:�șe�i��Z���\]r[o�����9�b�D}�}1��F��2V���t����H�i�hs<vԭ�%��%�C�� 5np�?�88p��!�to#�s��R��+���{�O��,ҷ�o`��R8�r�f�WX�u�G�ʻU=�}-M���s�R���㚞A�˞��o��������;/g���j��8VP�/j��Os-s67�d�e�2#ﾏ���4W[9="��h�K��[�SV��)�W�ßWa��|૧e����Y;��&��{`��ȣ���W����	�%�������1��)Q�#|V�{e�6�I�	L4ۄ�l5c+��k>��C�b��ꈸ0f�h�KQ���}F��*�ĥP�D�v}��'��1�"V�5v��r����frHu��7��[���F�.he[�"6;2���f�uh��K;=ύ>���69��L�T{@��6���훇��t��j��bG]�v�'7Ý�|ri�M�<(M�����;���w��}e�}�J:A��=e�K�Ow{Ʃ\���$��Q !�pq���S�y��F��F�`!�p߽磗����罰i'�K����k�����fb|���阾({s�\';G/��"ZJ-�Tt�K[�5Y��%������0�!,vl�;:���Yך�x]ONtz��Y-FJNB�AʬZ�Yh�0�-+�ъ�ު�4+ )�9/���*�k-�Yxa�����keV��GB��X�v^(��ӺӐ�ۭ[wM=�px��i6,9���1�$�b�U��E��(�*Bhn�(�t�@��C�FѼ�9wv��4f�cwUT�jt`Zj��b��"y?j�ɪ�В�L��j���eh�=`��4��cJ�yTN0�,�ɣES(o4i����Y_`��3'ѳH�6�(e�Z�4�$1jČa�����GT]T�.a��<ͥl����h�7�7���j�`���f�R��1;�����a��������g�����l�Fv,���U(��d�F�t��b:w�|:����e�̡b��S�Ku�6��YP��N��ZU�#PΦ�¯�����zy��sO>
��"q���"34{��e�t�g�y\>�`��97����k�믲���N����:Ӓ���(�G-�*��6�9)�H��p.�H�.3U	��vc�̝RG��}*4Ω��ۥ�u�h�Q�J����]���X[{n�zMre����KG�}�Yp��N*`�X�zi).$�݈�iTX�{/��@�0��E���l�w�� J��N�3d+x�˾�	��p	�'R=�Q��G�>�ԬUi���V�ս�����V]1��T/F�=�:m�}t��hї���[���K���b�ٔ� �D'�����"��.Y�|��	��T�2'gV�Ă�O�y#����'�����b��$�3no^��]�5��5��a��lG+{c�n�YV��NӾCx��U�ܮ�J��bv�$�a�Tfa����B�T�B�߯f�[�b3{/�1�C�8��Y����)��w_j�Oβ.�qa��1��4�l�r:�I��H���l��/���wOl�H����~Gd0�3����x�F�q#�]=���9�˹�����./�MU.����e��t��S���ãy�+��W��'0�6b�L%��f'7z�w�L�6�m$�����GQ�-��'"1�[Se�g�|8��1�4鷙�p^u��]R&T(����5w�#�fCvd�J)R|�����'۳u@<=�'��,2�k
�E�(ݬf�&j:�����m5�� ���맛�{�#��I	wM�Y�ܗ�jq���m�m�AaP��/�;M�����<��k�*��L;�[���x_�2^��l��������u5�·%��w�k��=�.Q	����	1���Tpu�<On�v>��ܹ�R$aL�͍��^�a:ET>���֎}��\�~"p)���jꪾ�{|=Y/��}�r{��s���zH ���H̋x��4Z�8)�a7ڗMu�a�O+�bs��޵�[:��o�[�xb�t�t�>���tܥ��}V�
�<;�Ț�;����^�W-5��՜�n;~���sY�Ob��|�P��s�Q�w����8�����H�ؚeݺ�_a�C\V����jjf��-�w���)Ɛ�8���o�i�[�Ԉ롆��e��&�1c��]�U�$�㝄�1Ah�����~���`������5��О�bvk>"/��"{2桽�q�EE*)UR��#)�(��UR�0T@��������s\�5� I   e�I  f� H ������^�����(�=���(y��Qg�ڗ�M<}���>�a�9ē̌ۏ���4a�JT�`(7	!��T��9�N*�<Y�Go��DV8�p�a@����r����� g����k���5#��܉ͶZ�WS��t��~��v�榦�U��+A�r����^���B�y�Ht��O>n��f7�z�Q�i����Kv�ʝ�������Z#����'��ʠÑ�X�{6S��L`��V�*�b5OknrM��-��ȷ��3���\6��=�, � �@�1a��Q��=��Qzg���҆\8tT�V��W���n�,q�t��z7�rS���4V\G�}O�S�c����P�8�O-�AM�ǹƲ�KM��mOsh�T��D#Dn7R�M�Σ{����|9��51�V����6z����q�;����\�ey���Çg�L�{z�����R� ��@'�@~�}q�%%"�a�L������|[�
�ws�>���G������oo/A�2(6Ը����vnn���D(�¦�q�Wi���_7��V�-!S�z�d�e�ي1|:�u�ٮ�S�m�#��Ķ*n��9ږ��[����IvKl�y્쨚�yyj;>�O~3u�yK3�� ������ f>�+nEW'܍؋A�iQ0�2��z���-X�b������G�ڔy�.{"�]�|�e��m$w+Ѷ�d���Re9��+�^�=�+�8ϋ�:�7����̶s7J+�AiA�C����s3�xƸ;��>���DjW���2�d����w�w�U]�.�h�҄���'���N��� �M��u�.����ܠI<��o��+yx�2UH�R1����И�VnkӠ�mW���4)�DO5�)c5ЛdiȧBp���a��qm��6�nB�oT��kQ���P!iLUsu05�vH�*�e������cZ�o�u�Rf�k��ٟWۯi��1 c ����F
X!]�h�]��E5�{�H���_%�M��a7L��2�t�g�aW�ۓX̉	8WJ�vZ-hq�+&\�q�y����L�I 	YN{m�x�IL���b��1�ab=*�c�p~�꾯��n<����ԍY�6:D�?���+3�����sy�|j��]�Ig�X�\Tv��
ҍ�__}g�z��J� �\�=x�rUU0�P��ȩgb�v�xv��q�p�/��un �����zk���kX%���P|��cz����7t�`�����t_{�i�|�Մ���\�;4�@$��U�r(Go�����L<�70û'S��G�\]v����ܪƓEI���<u��Ӓ>DVd��E���&�ʓF��0�h�ˆ��ڑ[�yS�2���Q���������<!s�-%)$�I6ڲ��W|�2���L���h��evFC2{Z'���:������v� )
��q������\>(�-bP�S!�R��)���s���\$^�x�7�����>8µ�<���ⵤ�Z>}�׉J]k�gj<
�rclo�`!Rq��Gb#MV��������R����h� >P��[Խ����:%�(�|F	g�9籎er�)V���܎��T�E�	˜���� �`�ɘAg��4Ovl�w�]59�0	�>����'�ͻ˲X(�H�"���EY2#�Xt�;�����| 	$  ��@ � I    ��9���oY�U�9魻��v=U����]<)��9�k
S����7������
%`l��'�zQ��/g��	%"mSQ��dƁ�)TTg�Hs��	����IY$�I"{�\ҾiZL0�X�)$���2̭�v������p޳}�Ir��e27>����eP�z���uu�p����-��ѺW�3�"s��ܰ�	K<�|-�;��>j��J�lɬntˎKoUv�eZ��D���rNL�T��n?��.�����Q}ji�q8�f$�,�3��R��ٛ9�*��_��3a���>)QCQs)��)�ȳ�똲cj�)p�[9�+#oCձ**w<ü���1_�Wꮽ��K��3}�Y� ���YkX�(TE�D.'?Ym5��jq�{�yfb�e����kl�y`�Z���>;�WWe�I���et��")�:o��4�� $��$�[bz����f�@��u	2���ڍp���|����+��E^'Î�h�9��NI%�t;�E	z�&�<U��+]��w� i�ӫ�ol��� Jotuc�B9��[5�+j5|��}�v�1�WӹC�ڸ�&���錷����@��ٲ�n�y�ͺ����Pɉy��]R�ԋۊ���M.*�r��ks(GQ��-xsK��#�V<�Q������S�kz&�5���m� �J�Kѕ̚���~�H��(��FQjzab�t����d	;&E��	>��K^X���X����I1wp�x��$��m�+#0>�7���Y�Y�����@��*��V���FFE�,�o9|�r�繾=��
�k���M-hA�g+�� <ܾ��º؊(ŋ ��> ����8ܞ���+��ʳ����6C�N}7=S<wfmL6�o}�q��]�mۦyb��gl�!�
��D�u^��̿2J�[�3wm�-=,u�?]ہN{����� O|x�st�bi��Us�%K[�������F�ʪ�r��wM.ޭK�"he2�I���퓻��/s�sB� -K�#��CdY��.R�i���x���7|���9�lO��×����틅V\��4�g�+����X�����t'�����F_�������{xFV��Z�!u�}�*	�Xט��0�fF����j�+�f���4Լ�D^qb�M��U�5���'$��{��tF��d{lkv��S�ܿ���3A�|�9}�m���>�	�AU��EQE�X�PH �� Qۗ���أ�ي=͙�r�硦��(�[7+���(����N��SCI����(]�Sׯ���쯩U�q���st��\�0�Q� S蒹]�9�8ҝ����p�b��bv�+�M���Ԕ�I$�}�.�N����\��O��-CL=:q��be^�s�Y�	X���3��Jhry�Hܧ8&�x�+i�/N(y��| 6W���¦ewfE�I9�i"юfvF�`s�\V���+{��CYLfk���ɝ��"��{�Y'f�c�NN���4��r�T�_16.*�q�1y�Pe,[U+�2�K�@���'���5�:mS��=&�Ws��ˆ�ᲅMs���bhe���3q�Z3S!���Qع�R�z�:�#�0"�j�[v)��b'=����I˳����n��Z�K�ֻ9�5^�y��K��tEB�H�Jӝ�q ��HPe��g�pEq_|��M�W�wW0��B�X`�F��w�%�'���>ʯ:����Dy��b/UZ�2�޼�HG4Y�8�)FmC��T+;�ma����9�;,@`e�ʃxj�t��:�`��X���:��5Q*�[u*�V�tPJ@)��@�d��A����	 ��)kT��4i)$+WyF�eAK/n��+{����*[���j]#5F�r�m&�h�^�(еP���s2e5$�q�)t�&����U� �UB��V02kP�A:*�*�$5FZj�M��HMh�2�*o�z�훛q�,�m�+��˶��%1Un���s��J�u�f]�y�7��w��i}yW�j��v���r�EGYuF�!�$&��j6�(q�B��U$�Y�bh�Z��H��e��J^]ɔ�FA�j���k01��˚�-,��*�%-A�@�aIaX�(�ұ�ۗ����e+X]��s."[��n���e�4���e�ޕ��T�)[��26��S�E�)=�����E,Z�G_��`#���@�[�4�g����W�$�H    $�w��              $�yR�2�2db$�"H $� I          [	1!$�  HI��      I$�$�f`  �        ��3��vw:.����ݜ�K��t���e_;�W���10�,�hH��W'���͝}�lՠ6����.��a�^�m���c�g�S�������$��27]#�݇{PX���C���3����qO�����S�ҍմwK�Փit�iřy���A���^��F͆�x��j���z^r�*\W��*��i����gE㻽HR>��r�'����H��r�]p�Z�eA��i��%��� <ϭ~8��݅����o��o�wďx�f�VP:��ۘ瑴����Zq�������ɐ�u���"��,ԗ� ��D�ab Yz訑�\���;�_ނ���I�RݧD�^��j��<��6�M�7s%лP�ߍ�oq7mtTq���3��[i&K �:T0��<��o�K��k��$!\6�JGY���J�Y�w*�M��tpm�d`�j�haT=�G��[�d��T�M~�#d.���Ju	�0��!�U-�������Fn}��{��F�#��m�*�������C!P����"vӜs5G��ʌ��]3��*��U6"L�ۑ���$X���MXI���~l�>!H���ZX�8r��q@ܟO�n�3$朰��
H�21��ŉ�("=m��r3�8QM�ɤ�Ƒ�$C��(��5(rV�'���5��a\�a��-Ҳ���`�C8r��iAK&R��Wy��U2k/��$�  T�  $�� 	$ ��;��̵�'ivz��vع\v�Lm&��氃p�Mn�`v�P���ͱ�|"Кs��[	�M�X�l��)��>Aʚ,ߛ,����0�u2c,�� 	$aԦfG�ٕ�!." J8\Q�u���]�MvC���]����+��)3ۧ&�w�37�s����"ç>�i"�W�rƱQw��˯oM���+'>ML���j=������'lH�a��N�:�e�nP+��E����d>�M:?#�7X�$�}�����+=_{�􄆟srI+����%� ᵹg椞`yv ���x�%ɺ��M<�C8E��|l�یf��^�c7�m;�T��*���#�G%!r���{�f	$�����ܮ9u+Wf�@�r�`$�N����3gX�&�<T�lL��>���́òU�\�
0���	�è'va�yZ�I���8 
+�ϯ����ᛇ �b&�j,�Z*��ER@*�EQ	����`�% ���� ,A`��U
dZOomͩ���]�uN\u��\�Ȩ&)����6�;TbL�1��v�a>1�WG_$��w^�b;�����C/)*���=�E�E���^ݍ|���=,8gn����Ž
=�j���u���eod�eO4/�׊d�z]��
r����x/4�ƣ���ҧ`ѐ�d�ț3܃	�ƌ24>���R�)OMv�26+/�mmgs��7`����U�fG�DG�ݭ��M���FW��Ѩk�i�3 �P�"��&�L���LI��}U�vߟ=p��n���m��(��C�+��!��s0�x��]w3�'*g4WY@Z�+�w�䡨]J޼�[=�n�������Sm�1z�F���v�hޟ�l�@$�x8{��r�*\��8'nP[�͹8�̂5P�œ���5x�{qțXx<gއg�4{ז�%�Q�ئ�R���~�P�ܓy��@Z��v�Hl\=�"�.����Z��-���R�$v+�cت�*_u�s%�7,��`<O�����q�8�����Sڍ���#79%�Ou۾i�P��&"I#m�5�^5���I�:�Q�ܨ*�V�
���/F-퍊��_��y��yI�30)�Kc���A[9*ٕ�f��'�ϋj��y�G]����i�z��E�[�"o��#��n�� 슙Y�[��0!DDh��uZ���_*,�I�*�:�l�]��&��f�m����I�#!N<]��<7���֯��>�uw�{T�Y诎A ��DFU�E3ݟ^��9�^������-҇�mfZ���D���g!}�&��ֳJMM��O�LK�Ͳ{�{�b<t�*žݣۂƤ�����f0N�ې5N:8�{�Ean��r*���^� ���c�� ��&�j��%�3%2J�?5Z�\&��U�p��١�.2���*:�%2]�'��s�]uh�.�|}gV��n�� �=��W��j�BfL�M����^�׻��9���I!2�z�7G��{��P=�.���H%���!Svo����)=�QA����尪��r����痫sݭ���&�S�����21@�='�f�[� ��d��¥��9Ld�=�l��.^�]��ܘР@@ |џ�*=�e�����P����:���m��x�>8�@��!�ֻx���I  �0�  ��K`$� 3q�]f�&�H����ǜX�i�rc=��>˗ίc�xW��}�f�w�������ʅ��Ykr`I�IBE>aF~&MHaBC
B��L�ze���*]�仛jkR�ƒjf I$�W���Ϡe�\%�s��%(X�J����� ��7�ޘ7=�eq;OUm�5���FD��Y!ȺQ��;�X>�e�.����)^:e,��>���.$�D>�rDN���[�$l(m�������%_Qt�Gm��vM%��4��u�d��3��Y�h��}��[�p����Y͕��)�)��ҽ%����UP���I���aU|�8�Xe�"��y��wz��9}m36U��̻�̨&�#���ӭ�V�`6�I��>�tQ5V�D�pIBl���r;�6�Ċ:�5��Rz�==��I~� 3�K�������~�qXI�#���Ϲ��OV�F�x��/~����"�d �*�P�0F�;�S���H��}4�{t���z9����֕����碱�pp����ɘ�۩f�x�D���m�h�gb���꺶�K�}]�o���]Ak6������}x�[�ڠ��%��Y���q���re�h�۳�&���c�#��mx����w����#���hXi�=�nK��xxz���v�M\�{�Vј��3L���R�dw���������,V��gՒMu�&�`.���Y�[�.�(%�^K�Ht���օ��ыbҥ؄�s�e�V�-��6j�I�+Y��&����=V0Ε���W�+��cv��d4�̅Qt�\�[ �1dv���m��M�
��-J��ci�w=\nM���Y�3I��� �{A���'2�$Z���޶!�n��l�z_N��*��v�<\�����|G��v2�Q�՗�Ac�}B��y�	�̘����i<��#����"��r�3�}|�4� c�u�*F�I��3|l�n�M]2sS��;2W�)*�$wU�.�sQ�eeY�R�v�QԠ�w_7؅-K�VIm��M�c�h9<a\0���!�Na��z%��1ۋ��d�_w�{_wZ~�������^���x*�$���S�s_{{��s���\��+�Rِ@��r�gf�
@�}��sp)5��V���\�|�Thij��+��j�u��I�ګ].gG�`�����{g�g
e�2W�O=����;����7������ٕx��|�9Mu�#q��z1�����J��0�E��`���D`-U5)]�A�qZ讒��y�)�>�9�&1^�Y�}� ��^����鹾����z�G1��oq~�IL�P�]���*}����`�TJ�sU�vf�^�����	� T�H������Ґ$��}ٺ��r��J̫���~�-�*{��w;��]��~}�!�ү�hB�8P��7v�g��R^�'4���7�-�����ҽ<.,`�Ƙ����9l��or>x��t\A����N�zf��f�3O%�o�o+!�<*�Q����Ň�`� ��1��ś��T�dTc}�U��)7�{T	P�-��]�dbf*�+q:Y���Y͆|���E���{.\i�L�_�f���cK��Lf7r�r�;<��[�Mf�V����f�}{�6ۚ=���b쪡j�UYER�UU%EE�Ă��X��!B�h	�Z�U��)��3ܮ_%�}�RH  %LH  �v  I!��l�P9�vv��Q[�O�l�$��ͅ�hS�tC�}����EsAR�2�ʸ�ɯ�����$b�Y+D��	2ߞ�w̳hr��T�B��ݽ��D��(�Go7{����Ќ�&d�kF���U����<9\b���]�T۰�g��u�1N1�r4T�c�z�\oM�l��r�f{��+v��n�j�g�ͧ+#Nн�\g���AR�<��̼�����[N�h�K
�5��q���F��Omdu}�U�}��:gq����@��:!a�L�ӤwS61�=���p�G�?��Z����YNp���E��k�����mu�r͕��6�.�&z갈�M���Ff,������I�:?��_|o�����$��$D�{$���-3%�'ؓ�ն�z*��/��o�٧�Mu���ʮ׶�8n`u��]�E�������K	���I��3�dP$X�k]�4��~�yf���e��F:�`R�����κ�bíYa�za��uk�Ӳ�\,�,��U��"뉇Ώ�W�|ǳG�5��d��:3��APc��CL�ǌ�ϫ＀]����~#$;�6{{D�n������:+@�P���LM�Y�����X�4փ�k�zmfw73H>�o^Tٌc\N���)R��ZX���<7�cb�g�`R��{��5G&v/Z�s��J�FC�����Mv��-&�M�B������Q0@b�YbtyMT�������>�wv��S�ະ͘�(۞�ȫ���'k�sM6X�8��)���#��@�]���]U�{6տ{��m�¯�&ctg%�)�;��!��SS�u�/�]�5|DR�?}a:�����&��ձ��mH�jr���d����.�J�sz�����x��ui���3�Y��F�||��0��#vM��7�U�#��u"�;t�1�f�NV��y�sy��w]�M�����eS]�v��fE-u�^�Z�P�)��
����a��#.o��0o=~8�B�$�Cu�2�S�(1���֫����θ��ʪ��wi���5|�2��+-ī(���֣uSL�.��Q��R,Q���(&WLŗ2AQ��C��C�PR�ۗMY��ѱ)o^8�*���`��2�R[@�d�j���]�]f�Va�[t�����2�����>�<@��Gt�Р�5���w�aEk.�����:��zr�����&�X�1�*��l�h�MUQT�зE-�IH	#6��D)Ac4Ζ�h��~@�^���F4���[�'�P$c)�Hڦ�	���pQ`2H��8���j�?L�>��>t�1U��R�uU����=�=���Ά)iΨ���^t�&?����6�0(���X��;zsa:��5'Q]��,�gb(1wӮ�Am+��p�6�3�֍y!5eS�:�VkL#�E}>�z2R�	Y.����,4�үӮ[��
g��յ�n� nxseT�:�*���I5��n�[��
��`�N�+�ld�7�^����8��s�FG}�4Գ#���gTx}"@���W=zmvWf&�n^n�L@fi8�hf���ܭ}�)�/�}����<4��1���66�gK�-���=/�2��D��1͞
LJ���i�'��e�H~�7�����\������B��Qdh�5�r�|�#xV�����u�ы�G��.�[���Dv04O+��d��!V�Ƴ�)�k Ũw-��ʍ#:ڣ�I��<74%�9|Y��Qx�1�Ɂ k��Z��$�\)���d|���� ƺ�]3*�g��w��S	n� ����'�NI����F���.K��D�s����0ZC4��̣���R���+��W4b�U�E8g6��k<�L�C�������/��^����]�I{=�cb�q񣶦�;����Z+��L��D��4�����=�2L�k
��J� }�p^���� ��G�����0�+�WY6��Us.A�WG�v�[�˛����|�(�
4]�Z�(Ɏ��}����z�]7��٫�����������`NL�+R7�/n����9ОR�W��ͨǸ���	3��ˮ3�nD��}5L�|���Ԡut��j��Y�u�;��xʽts7�hh75AK�T�����Ҏ�s�j�r 럻d>z�����3
���q�&	��RT�J��<�n�k7�?B�nno�����x���
��I�r�Q�{��eÍ�6��ὥ�G;���_E�#�>F-uҞh��e��w���X�'��V���aʍ��kU"U��FT��+smK&@�7�O��˨.�>�M)力b��@�oyб�H"�^oF�w����٭%u�6Ҩe� ���(C,ˑ��]o6�NI$�I\��Ps�m�D����4e�e��&!F����U�@�}���N�x�Gi�ߟ�~��/�n��3��?0l؆;���т����a����b�~���9����{z>bu�����u�O�؝0k�Ũ�1"D��^ӊ$++A&9�5=��zY{wJ�nf�W!�X`ZNN�:V��[�"���$p�1�F)p0oJ�3�M�G=c#a���KWj�B����T�����ːj,1'����;t���w���z�!�r���ϼ@��I�z�uOj����Q�ן�{U�H�����nO"ƀ�2!$o���>)�r�5�~�~��;_B-��`3��Mf�Q�绣M��[f=ު��1̨5w������@���y�/i�����%7���   |7�񵳶�m�IL�� 2�0  �@	$ H ���Z�3�;�z�K'������d�O�Sr��y�g�v՝	���샥#O�H� ���C̱�E$A����d~b2���R�j��P�YLJ
��K�!/..�I�rom��H]n�}{�}���
B��J���� f���&z�ȣ���;QG:X8!���ש~v� �5߷k���r���_m%�}��wn��f�%��9�sUD���F�S�(I�`���wf�8UZ�	b���k�Z1�����rk�ƞ��f۷|��m�V���J�6;���!��W�4���A��q��=�VOmC��].M�?�A�+�dn+0u�B�\�-�ѵ�y���殃�}��e/��ϩקϾ �$"�n�C9�)1�z���)N�U���WSȮ��5�V[�+u���wy��ۃ�@��/7�:C/u�G��H��aU��:�ۡ���/�1/u���k��}�3�x�U�苙G��QZ�l�=q�~rb��?��(X�(=卶Ҏ6ܐ~/T�(�Vi�^��efUzu뉷�j���9�m�O�w��m���X � EF@DA@�#���1O��/�G_w�j�G����8柫H���!4TF�;�	4e6a��W�Fn"!�]��te������ß�o��-��p��"�'�OӇ|�1W��_��٣ش�O�={��B���O]���!�����o[�Ƒ�^M���xK��FM�GO������o��B�Kn5�5�-�����~ܒEi��������H���4��Ǭ���/|�^���9z���Z�%��O&�B��۴�B@4��7�t���ݭm�]bT���=E�g0����<#�pbɃ����
{U6��T��o��v���[�V{���MDL�0�Gm\�r%ME�������
��#d�4`�����4p�i�:^���Rܨ
=�u0��쌩q���������I����߉�H��w[͙[�̽��cYF�0����Ӊ^�~���s�HA^��u�{U�j�g��v����շ>7M>��q7�:�5R�Ŝfc]C���ϯ++48l�pg�X�%������nBΉ�����(�~��1�a���#F	\�����.� ��hx7ˏ}Yu\�xDu����f:~x��k׋��۸j�{�-+2ξ�3U��V��o�}�r�;��9"�,~������r��u�>�2
e�5�y��0_)?mt�nv��wn2��b���q��Ӎ^I�ͪ� �>��7聁#��T��Η�j���i���ϱ�ohW �QȒJ�3˪�#0��G���u��QO��rZ��uue�K�N7z۽�Ogv֪s�c8��eU��s��x��N&�4�0�=1�-u2"�X?X��=�Gb�-س��!��k�i�S���Ě�C��{g~�z�����v [־��\˭M�ʹ30�-�r�v5g�Bh�2���gj$ŋ��� ��o��X��8ޛ�N��{����C�����r��j��j�ۼk��}�FҾ�ί��4�Z�b���"��E(�8c1�S������ϛyUxa9��ʀVRT�Df=����GV����`� �˧c�����G����&���n�ۧ�R����e=�i5�]'_4ڻP�Jq��S#is��Z�1��b/C_vB"I�x`f G3cE���(W��]T]��h�n�]9�ɐ��X���Zr��zپ'qLI�rE@���{������sP=���B�,��:Sɱ�1�0���hh��#�\�rB��~$�U�-��HF{G��sw��h�6�3�M��a�:y��7>�<�+���߽�m��UE7U�w�-�_N|30 /z�^�����7!�L(L"�M����^�8�0�M�.����Uڲ������u��Ѯ���&3߈�����|z٤v���e�G���L	������a�V���da�J��C` t��@�u҅��3Q�B��b0�"0F���X�:^��G{�  g�q������p$�"��b)�ņ"����
�}P#t�Z#��ƘY� !�r.?fD�� ��9&dS���A���"D�]��0�b��Hڃ���4��R$L:P0���fw\[����lB'/5ŋ��H��{�I��$�C��E=��x�!�-Z?kj#��Q�ޯ�=ث��P��2��! h�\��S�˪-��j��f_x����V28Ȼ��Q}T�*�]�8���ݫ����$�  �� �a II$�Is�w��{�a��n��&�T*m��A2膸V�q��0f@�6��� J����Hy��4e?�e��Y)E�&⊤]]�j�[�z�|�m &$���3�J%̉Lb����O����%>P(��0�Gql�B!{	��jF��h^vJzO|�L�@�f0���?_�����\!�I�qCFԸ��yw0x���$p�sZ��Y�kp�;v��hN1+����'x'+���	TN(i@W-�r��C|��|��M���|�wtm1�W�i��	_��sT���W�nHBhsZF�~Wj���u�P͸2��__1�˽�-!B��a��"��𰧩�\�F�����C���u|��Ĉ��ʘ�?wjM7�����;�K�ޘu:��	+n������E.�۳0"����d����Y���wYZv`���H 3"��8Rl,�����K��_��4ȥ���s�33y�_L޳r&@Ȁ7 2(`�m����4��~�G��
�ƈ������ی��ił ��p�ZO!)^�S�E쪘>���;��Y�i90J6@B����9�O=����9�t���$_0���AAIL�B(DX�B0E��n�?�ٝ�u"�z�W�i��>u	�gq�}��k�&�a8F�l��*c�6�l�H�����_٤���$<|G���ų"�}'��Z�Ԅ9��/b���"F���]ƥ�g��q$R7� �(E=����d��N�<��4���SN�>?!
��F����H��[��}�qV�?�S��=��P{�I!lF���P������7����^v�k��^$��Pi4��U�:�j�������i�N�+���sX,���f^e^��y��JO��ǚE�JD���NK'�A�J)(X�b�3�a���A@�b 6a����-���_3���i$�o���dr/�E�)��c�DS��,K�q� �r�,�Jl�m6��ꨱ��'G��}�._nu	�o�UrDp�p@ㄡ�tC��m�R������}w����6ۉ��Y�>u����������\uEr�<��\���\�v��I�ח�i����9ۛ'k{;Lر�׊�S�+��$F��d:��q{X�����դ�59��&%�g��_ޭo�9|u��h��� ��{6nM�����/M�-l�[͎m�5wc����xz�Z�N�����L\ty=�G�v{�q­��{�m�+��k)Nz�������7tUU9����y�Ey�ɕ������\G�3I�l��i	���X�J�	D�
|�C��7bxF�p�٪�BKߐ��~�}}#��2:/ d��C����t�&���3���b� uL���xT���P�����F���#`����%��-"��<l���U&I�r�Q���$�É�uPG
�`����X`��M��l���NP���wU�j��ꭧhR�vq�p�u�_Ͳ�=���YFni�`��H��M-x�2r6�1�up�>n���T��y6�o���<���=��U�x���₳�}��\QJ�h��t8(�XNnt��dX����iG�6"�l���NCCG��E2U�J�ˣ������߁Aa$Vn�bT��#B�`����B�*��>C�+W� _B'�ʯ/��qv�~��j��z��2J����__y�:�a�*�tP4�(E*QU0Y#1 ��AdY,A�
��T`��*��)�(�@�dX
����z���>��5��|�[�&��N��ӽs�0�2f�7�z��O]���}���ᝒ��=3xa1� ���UR��.�#k�"�]�Ƈ&:��	!Q��h�ާ�YHZ��#}��la��z���}�uD!�Â0D��i5Y��$��6�!E1V�V�L-�,Ģ�L���]��t����6����6� C��@�x��m��������i��]�2�w]�ՃZy9�sIǌ��N;u�����SC0�"6�GS�aμ�f���"�ŀ8W%"�c�,0p����"6IG�'�W r$F����?%G��m�I�H���*�bg`J�� `�Q�&�F�#>K�J�Yw�[r�	;����/.��q3T7�]��>�W��.�A<���Fp�I`��yD��� ��
%����uF���u�V�}S\��Q�s�Y���|?��Ҁ!iF@Ѳl�>��,����}����y�k�_W�]b�J�=����W����q��M�j���]�׫+����>�-����?� $�O� �I����?��	��U@?����@��$���!-�BI���BB$I g?�^ I$���@ �I5�I$$�~���?��� I'��������'�~��$�I�@���dIo��� I'����L�I!$����?x�?��rI$$�kƿ� �I� $�O��@ �I9�FX I'�W��5�Z�r�a�I$$� I$�s���� $�O��I!$�����_����?�w$�BI%�����/�߀ �I?�� I$�����b��L��]�}D�� � ���@  nO���>w�         ��(P� @��MwL  �     �  4*� HJ��h�J ��Ф�����QKlR�
��H��"�               w�RT��  ���G�U���}���w�������*���}ކ����鯵��vʌ�ۇ`^��w����j6��>{���� W��kw�z*(�sZ�� A��y��}�>�u�_|��υ˧���}�r[퓍��Ӣ�����vm�|3�|�=���=P��0;�u����**����Y��S����   2|�/�&��e룈Y�ҋ}�z�Μ���|k��ݟf��ЋM�nt�o;^ڕ�����}����3#�g��m�ܩn
D*���`����=������&�^�J��0�M��N�Nڗ�ѝ�|�{�ܹ�ne;w9Wh��F���ע�z[x�ʆ�  ���]�}���6WcS��u���8�{��k�g����۲-������Ͼ����Ыg���Q����-6���*G�!ZٟvtѾ>�����os�E���wK���3���/]���u���}=�+V#^�>m�٥���������JIJJ�  ����}�����[V���r]��ͱn��mvצ�_|��i_grUm���q}oj���fTz��>�pU]k��5���=�:G{��R"�2�K*̵6V���{��Y�m{����P��g�U|)6��W��}{�Kg��Gj�O��.Cl[8������A��R�m>   H9��=����]i��:����]�g���֩�W�n=��w��d�����#G���|��y�w3kL����/��@w�o��6���8�o��=�{�������UO�Os�U����[}}�^�U�W�7���m�l̵/H�8m�ox S�)J� 2h S�R�� A��S�"R��ddh�UO�ڪ�JJ�� @hT�)��J�   	4��%B)���4�'���������������s�{3�6��-{�����7{�$� Jy�$$� I '�!$ h@��섐 ��!$ b ��	 @���^���	���Kv�w3�4sўL|7�'�`�vA�t�s��~�*߰W�l��w�MBd���ܻ� ���~o�n��҈��4�*�!r�z1��L�v�K�\�a�gCּ����ιb��U/[�3y�kI	���˯vpB#*{���(,ʖm�8)5�ݲ���fC����]�R�;�.+����=E��N�t�`{��	��B�gL�{���H*,�󰚮e�_dl7M���Zz����JE�8B�X�F��psx�u�x�p5e�2 ۈ7_L��n����fP�r�aw�#m����tf����YKk�f�|wSS�y�&�}���U`"OE5U9B���-3'�&��,:�ặv�Ș'"�(ޝz왷Pr�f�	;�9Rɼ�-&7<K{�ټ��7`d���u5$':@"XԌdճzڴ>6t�v�Ք��֤ӓoH��tY�+X�vf�	&����!]�����vc���`�M;�_(�wWEޅ��F��C�ū�j�i")BS�,h��,:8.�8}��`B, 
�##�,X�b�
@�$�PDPTX��$V
2,X �"�P�a 2�
!iED�`6��m��Ȩʱ�����H�(�P�mU�QJ��H(�DR"(�*"1H,Z�+J5�FJRTE�"�Z��P����A`-a*eUPQ��ŃcZԭJ�V�(FҪ����E ��A��X1�,6�E�(AE#��j�E��UU)H�-*��,hX5�6U+m�FZ6H6������`�((���"�P+Q X����$�d�I���
AH) ���PH) ����
��
�R
B�*AH) �E�i�+Z�
B����!R���VjDI"���XAA@*AH,���� ��`�XQ��(*��-@� ���YXAJ�-E�d�R
�H) ҁR
AH)
¡XT��R
AH,���-h*5�B�-�V����R$��)Y+�%(�+#+@ )
4RP�QH��VE,V�PA�0Z��X�mP-�)
����� ����Ae�
�m �`T�HT��R
AH)�m ���R
AH)
�� ���R
AH) ���R
AJ�+�AH)�m+%H)H) ���R
AH)H) ���R
AH)H) ���R
AH)i ���Y*T��R"""��b[b�PmYJ����R
AJ�PiF�QR�QD���V�*4Yi�X*��X(�UUb�(* ��UQEKJȊ�YKE��ԊA@UVH��`�eDJ�$UR
D��REP���)`�*(�F*����*(E�>��Nu�,�4s���y�"!�\�j�8,�n��i�`JVk)��.Q�>|�A�d' �Rx�9ɬ�1�x~ݬ"�KpS�%Mǖ,!-[���w&��
j�(h3/5�Ӊ{e����@=�b8� ��
�(Ù�f_�ᇜX����-�JP�`��A:ˣ7uq�����V^.�FvLG9cA��4ڒ�K�G�o,�>Pex�\`�>Ü�b����
�5mlL��2� ሜl�N�՚2P2k�5�@Pƞ�n
L�m����-��M���oN�d�p^Y�s�i�rK�N�]��,М�}�h���,��
�VR��j�NS�3�.�n��&�PGL(�fs�шp}�8~�Է��O��,<��9'�D��6ڒR��� �Z�Ca��x�}[O|ZZ�����.'�j����7�/0W�.�C����*����
DO��t�������>���k� �O�
�Z�����$��X��M?&�b_�� �ɬ���������N1�+���6�)���Gx~�E� `,[;�`����IY�sc���[i�&�r���:u�p��Q�Q�7�3s��æk�3��J�!���L7{�o�o7�2߶���b��޲�]~�y׏4Ƀ0`��^�����)ñ=��wsN���!�YRQ�-� ��w|�s�\8�� _vgm�'�"�G�b٪����ҫ��6F�6�c̙]�mds�f���$L��L\_��r�0��f�T��cx"�^4p�w�����t���')qۭ5˻�Y��x��4��	��vt%���-�3�P�+�N���%+݋,c1�]&)�%�1�ND03��p�{DQL�ʢ8wn]$���.�D�\W<�4P����M�O˹d?q�F�r�Q��c�����G�|�y��9>`՗L=L�<�!�3��_KM}r-�	��2w`Ő�n-�<���-��\����08��^7lh��=]>��F;tm;���[<�h�I�,
k΃����3�G�B�EV4�YyEwy�d�W
jj����P������,��5���4�hѱ���''��B��m!c�dΥ��*�}ʒww�kO;~�>�\�����k��S�n&�+gcU���f�m��R�(N{b\�������\��xs�SA�z#`C�s��>ܗ�a�Q*\9Q�g��<�0������\A�4�\�� �M��X��ӕ��$0=���g%�MRΘ��Ntt�֚ kx1��5��$3��#pfS�,�VX��ۺ'R��$��UIw.u44�>Sz�jK/m�Qj/�Ns�f���+b�`Mi"�ɳv�1pĶ��NZ�/s���ۺE�/+Z:V� ZoB��y%f�4�i�Q��F��q��:R�X&F#T��vNA��}��ca�ow� -�d�֘mV��7m������&���&3;h�r��LRIǲ�����.I!Z]�u�$|..A��6��Z�C��G]�x��t��M��x�z8��u@�rK�����ː^�59�/�v-ݗ_*ք�rk(�)K�:�TN}��Ґ��4�l+����7N�xT�F�ݽ�`��%���d������w3#ry�[�F�"Y��A���v*���x��_)
˃l=")���wTI�zm�^E�^{˫����Ɍ��-]���u���qs���]	vA��4�T>avՋ��;~K�i���{���qI ������K�hkp�n7�7������{1fӽ�ϊ�=X�eܹD���:2s���ѳ�)P���1*��	�p	�  �4��\53AܺnA�_�]u�61E��u����ʧG��TK���Z���5�r�x��v��5��T{��]��b �DdD+(����s��-���j}�l�$�%��Bzi!�Ϡ-���&0�j�{f)Dp,�`��h{������iO�x1#Ӝ����9��!v��.��i��Mϋ=�LTK.+�����㻍�q���z�q��q����MM���v�.H*OT�RB�\�t����hF���.0)������!J�������x��vR�0`Ǹ�:��{u��g�ǎ$��)���X6 ͠�ۑ�.���z�{8�$7!�N���IZ�ע��A��&���7����{��. <N=2�ѝ
ޟB�8�Ao+��]R��}!0]cݞqqg�wm��.L��3y�<AHg	�e�J�>�(�-|&���/�޻1i�i�+&#�i�:.�h��N���wj�����X��6�7^��קF[΅I�[;+8�7�k���ceY9��:�H�7ѬU���"%������b\V��^�����S��5�)�{#C-�m���o%�n7F�%��K	j�<h,��X�1Ȼ��� ��wTj%�eL�3,�f�Ӻ�e]]�9�VS!��0�[x`�d�%~�v��x��Xp��f"!��d�tXY�;OuGsF��Bs�Ω�Q {!�9��	N㶇{gI1�NK��YB�3)D)�Ơ7��;F�k��Z�I�V���w:#\��y/�����y�>��p�.��F8�ռ�7����"0��?o�x2>Z$�yP�9���x�w�^;�:h�uĳ�l�,x�L��Uy��]�@gs�䁝���r;1g>fK���ֲ�n��JCW)�6@�`�S��7���ݲ�����3�5�*A��"�	�� d��7Fj��X9Ǆӷ���1�@���<�do-�v���>ɂ�
`�y؞�^�_G)�P�}���`�UYt��;�j�7��FF�����")B�FS�_n������i�%�$�K�0�;s���b|;���#��Bm��B�t&�����!xt���gn���0'P㻢Ep�v�F�|�ٓ#u��z-ߺ�9L��Nl�׭|�.X0�#���	kt$c;*΃mv�6s���,2���CD�˶A�{.(�*Y���o�M3/�n��j�7?�p����k�ƽ�R�#_/�dcX�"��J��lʦ���\���8���xICN�2g,
� Ո<9����� C6��
��tJ;6�w��s	��y3���E�{ooi�Vp��{n�7\cqC��Xhа��M�����F��۩��qi:4n�D�-�<QLdl��g{��;�im��p��jM;4�ӻ��b���՝�0`}��L_F�}x�7�F�����;c����y(qД��B��vvb�8;1S���i�7�[N�t�1��VT"�Ӄ���;7%'��~* u��<'H���GMf��ρ׻{n�=��n��tj��6��+wǷװk����}&�>��l�z%�#�;W`�nʓ7�w�gd�e�R5R%�\�e��A}y]��*���P,Ӗ�\%z��>��~HY;̘AO@��9氮o�v^9)�7^���e���	c_
a� �e��&%O�_�8��i�-Nl��b�wN�=�D��$��DJ$�W)�NŃ5P.�o�iհnS%Ž�d��x�K[�ks���������]^���i�5ϫ��M$� ��o�n��n�v�N9��Z�T~rk!�����Vބ���s��:�-b��� »"n�s����Ue����b�nN�0����w�wof���K:�Il%�p���֎���'��0M�X�"���;��rCɝ�F�sN�Fs��	��܃:�n��+�I^�DvG�����M'�k��,���[_�w��9Ѓ��])5����ڡ˼�Ղ������;�pUǃrb�Z:�=Kӹq��w�T�[ϗV��x-7]��.�VD� (�5@uB�}��wz(��ʃ ��R�����E���:��F<he�H���y9����͞𞞭�σCn�^�ohx�i���{^�@s�����	4eH,g�]�/IKGd.�9zY�^;�,�veĬlx��&Hf;6*�&T�����왁�w��/$��5�ѻ K��;ykʾuP��T�&X2�Z���3��u�?��oL�>�p��_�u;8F��`��է����Y��H����6��w���!#�Iԕ/��El��A�ۊ�f��j8�ɀ��Ջ��Y�q�V�1�05P��a��g 6>;���L�fC`,��{%�[n��Va�ruN�Ǳh2��L��1�8Η��(ҭW�:��*�s��q���­q��6o.oK��v�h�B�w�w�d���),iW���F�����w-���c) K紷V�Εn�T��M�(��>��B�<z��ĳ��5ם�$%����)�O��gg��`H��Z7Ě����MM���*Dq��V����Wo�Ӿ��\�_pPj��95h���{ժs�g�?{tk�����!"9}l�-�����s�1�w�=�����/�z�����!ض�<��]�m����d�y������"y\�����X덂��דy�=�������VS:rmS3�ܥZ��� t������8#ߙ8��T�j�G�߰o{�/yl�ul��]"��I�4��ڮ]���^{ڦv�76��Y&�>�Y�H�<���<IG���������$�xLgƇX����]�.��|�`ޮ}2���X��*��UXSF5�W:�}$|r]Uj�y�K���Ҿ��O[u���m���U�ۛ�wh��\�[yr�g�O8p����1d�$\FV1q�*���5lԚ7��1/�l��@�3��͛���u(������N����}�I��̹'sNŇ��Nx�������Yx2��_R�F�# l�O��k�v����G%N�%���t�:�]�`�3�Y��ǝ�{���I9}g�&P�V������wNMb��r�;��Z��t��;���gtS��Y����t��b�;�.��k[^1���J^��ėD��--�+(f����m$��۷tc\�i�E�����%�gs�i-7�0��b�=�xD�r/ý�{=��0<o8lER��퇒�MFj[���r��(���q�݌����yI��_ܙ�+ޑ���b�����7V+�Rlf^QS[ײ�%�<�]��ŚuFs3v���l��l�<�o���nOn��%=}ʫ�~!?m�Ǥ�-�l����@��L��v`ҒK�I:I���ݳ�M�m�o���I�R��Ĳ���g)/��ث��K]���ivf���,g�>�<]}�־��t��_G؋���|W7����^�^.A���[잝@ܦ��(��'�N�纳A�U���Ӷ�	G�s�Ú毿Y���y��eC{M٩Hx\���~����{��c�W	��I���5���ӝ��w�Q���y�&���y׭�k�[�^����9��5��Y3sy;/�c&qut����&��vfl��E���M{�ޚ�)-���P)�'K�l��v�YrT��ro�����;��Dҭ�x��7R�U��P����]�V�orfs�jB�a��rt%k�ldz�r��H)���b[�wq�*�b��C�D�UW�V��no�5$gڮ�O��Ö(ƫ2_8�e�3�2�������Lw�%��v���ċ�W/x��@ɒ�}D�fy��F�wm�k�e��S��ڈ�V�^�,�zR�;�.��'\����R7��o�E$��Q�yg^�*���ǵ�3n�b}�Q��F^����e�]14� �h�t�*���
0jj�{���˃�O�&�\wQ���
U�H38=ޙ��8�s.���oyr�t 8�N�,��c�-z�	��Av�gS���Яy�4L��U+�_ ��u;���y�+�<��&wH�x��x>#��)k8#�ͨ�_Lu�LR�Al�����mb̮9�l2��G�}�q�+F�/,n�䯹}(����_#��Pv�ţ(�[1�(s.�� �M��A��X�	��������z�'{�=ר������^����/���l�Օg�\X��ޓn=�s��(�s�i��-����#oYGs����Dk"�u<Z\}<0̤����JN�З�����R*�o������*W�A��Z"��
1�L��
��S���$��K&Jo�Gj��}������듆��m%�+��2NtV�K�0�1wC�h\zY§Emܬa��.&�K��ٗ���J�j�hy��Ґ�|oph����.�K���'o�s�	��n[��wgZ��b�5���x��]�A��Y:��l<�+��s��:��Y!$h͋&R�c�vG� +�\_1�α�"@\�e�۞�_j�5�A���������i����<A̝�NOi"y16=����x�$V�yL�����j����C	���뙖�u�z���^�e�G:w���^��sۇp^�Z�]��۫Y/����C��<��4��t�GN��������y\ç���Ƭ���S#:�\�mK�GGmZ%�
p�m]�� n�E�B�(�� h�/��
��w2eݼՈ�.4iL!T��b��U����v��	�K]�Vۅ9ܡЎ�У��Ж�Rh�V�E{WX�&VY�,�z�,L��v,���К�n��A�߻�	֠gNx/�[�h-4 H�+xw+UY���	�UI�����R���^k����u}	ٙ���i�J��ou�����ޒζ�׹��������'�{���(�o����~��M�ʴ��[@fCK�8�u-5$�!vӮ��f!�K���s���T���5 �F��xcc�q�5ծ?{��2����X��<�����{��F���}I�k�)�y���{���b��Ûy��3����Uƽ(}�׶�r����iq�<:�=�^����=�U-����l��38R�z%�Ej ��5S"�`�o�2c�9�s��nn=�$�ȷ^�]��^��/:ۺ��;2mٻ�x	3��f>[�I�:�3���$��V.:(ݥ�E�NI:+8�^�K��kz�(2�"�cE��Щ�s��:���)���c���	�H�eԻ�I\�w����is}��#;�;ɽ�����wm��ݯܬ��f�pP�0���隮���d;���K�/��ש�0cB�\R�c#3�H��z��w�����������6qd*f
;ר�1�����Gu0Im=2��9��a�Y��ʂ��]���@�V0�b����ͥv0�}�\��O�N���3�b.���'=������^,D�6��OfV�P��>�;3���5���[�sF���fO6�e$�yP��x���FTUbEP�p^OVIz�I3D3�k�9e�ƳB�ْ *RI^˺
�m�ic��w��\�N�N�#���+˝�2���(��~m3���w�b_r g����A�m3L�^���;$����)��I6�ߦ�a��+�u۹v����B8�e�\���=�į�r��}�^�Y[82����#���g�{��b��`�]��"=kr��r�`7˳^Q�'s�ayrF;��n�oD����z&��t gf���.:�Y�c���i�{3ܵ���Q�Մ��$]�"f�Vj�VA�x�M����}�倏c�/K ��q ��j]���L5y�F�D'n�3[�B���5�us�ԝ���@��W�D��3ݶ�gZ[J���\>�����8�*w�:�\�o�=�yGL����&	;�\,A���vo.�����x�kkqV���r�^��&Z���78�z6U���S�rY�P���2E���Z�j{��s�ܧ�e��D��7ݚ+ELWZ:���^*�s��)�ߑu���Ӗչ��ts]#�d-�Q	�f��K�P�h9*6:Msw ���䂎��s$`ՙ�X�{��S�{݀hW7��Nu6�>ޱ���i"r��܂�v��/0���Z"�X�=;cL�ؽ�$����6�h���:�-b��WOtGL�kF�\�0@��6��b�x��Jbs$<S͍I��]�E.�A��۸�υ<�J����]��T�/u�Y�wZ���Y����\bM6��G��"��嫪>ܡ6��O7s펼�bm0��KSˊ�/)m�n�֭��|q$:%/K��^��ޗW;��'��C�hT��힘����07H�VͺN�ݾB�ǕJ�T��t�/#u7l�/Nڛ�N�%V۶^ޠ���Rr�{�Y�W���t�tp�j�=3v��k]�$���xr%'WcS֖�u<�gY�ZL�av�d1m�S+ay6P{�i�G���Ɣ�\n�	N'���*>��*��9��.n�6T�����h�\o\v,0�*�<�N��6{��ҫ�Nj�%n�{���� ��LJκ���Os$|{����6	�풬A�ŢkΧ��(ޥ�^|���(��y�L�����#y�����P�zI�_%����x���yFz|u����f��_��]�w)��5� �m;$r��J.m,Ѻ�a��u�W�C![����wj��N7ղ=�)��������՝$p�-]��Iw�k�9�����+Cx�/l�l�M�  �ªx
� ' c ����U��D
�%t@x*� ' c ��=��p0h6/;"�0��*^��1���/T
� ���p�� �p0��xb�ׂ�7;qJ��R�����U����v�m��U�s�V�z��,aWD�l�
��LeS�e�
�7������ŕ8�u < < ��6�*<��]M�
�,�  N ���{��k�gT"�@��t� :y�=T�&��QonU�
�燭��ڭ�� � ��Puh  N ����	���p�� �p0 �	�*�� .���AsV�vwK���=m�   6*���S�1�p�� �p0  N ��yTN�z�����=��>w�#@�   ��	� �w��]ܻi ������;ݽx ��8@x x=�*� <G�n�b�ګ'7�u�mmV.�
���l� �@d� wp���� ���
�   �m���y�� �R�m�uTv� 
���U��<*���1�N  Nr�=N/ C�e����ح� cT�����iHw�-��bz��n]�J���T1�]U 8*� ��}U)�8.�݊�7����T+#�V�+��^���m���ͱ��   U    ['=O��Y��Ԟ�V���T�6u�@��s���Ъ��m��u۶�
��*��T[@ U�*��n�P�U�ʫ�����m|��G7*���v:���׬��;��T-�� ���W��73m�  �Ա� [%UQ�}�K�  ��^��f������gn�u��n�kw��;+���^���^$�R �M @H�P�ƚP�R`�l��o/m��R���r�ͷn��׷���\�'n�Qwsy�緵T lm�s���dY����{�k�#v�(�P�*�  U6�C m��'�����ځ�-�f� T���T v��   *��lP  U u�o[��m{���ܗgowon��F��z�cN�  �      ��                       VR� �      <T      '  %W�*�l���  ��   � I�    *�       T�� ,��@       � � U�T� � P   `     P*�      �@e�*�AT T    ����
� 	�P U��^� <� *��GE8�eWp1T!�C�` ��|  *����V� �           
�                             -� �   ���>                                               �    �U��T      T���Yٶ���{�q��{j�V�;˚7�k?�	 @�a$� ��B��H ����ӟ���~C�I`B��L[��������f�)��Z�bO��4Ye+���}q,u������{qN���̇�(v�r'�VPN[���Eջw��8y�~<|Y����
5<{6�I�5="뼭��./z{��q5��_w�F��">��J��A'ni���v�a�ߧ+��WpO+*IӉת��Ş3jY��� /������_fZ�i`4�0قmM�[�[���Z����Z
!��vݨ��bOs�D�W��w���ߤ�wq=��R�AC�����'�R��� 	ZD�wx�ǁ�լZ��V{$f�ӂW��rS;6L�O��ǡ�p�;W�7�L��n��X}:�V���L�K��Wr�r9r(�<��������S�$�����s����I��軆����{�	s�z�W�L��w�Һ��3ؓ+�.]ܤ�c�,��`����[w�-a��}��ﻸ�
� U��c-�i��a�v��{�m��p���
��U9��Z�컗�֪x� ' c ��  w��1�3�� ����\�֛:����T��=T�����)��sg�d�ݽ��A�筀������ ��leR�]� UQ��s_^z�J�.7wkWo=��@��jM���GYn�VU�UV�9��ꪠ      
�  x  ��`U ڲ�   U  P  �' ���5�)�J�(         P�          ;b ;�5������׽��}U�URy���\��˂d�t��+�h�'�g���%��殆r�wz����{,���~���rFc���RIm۷� )�kM�m��N=u�=W����/-�=���E�v� *U� ]�[` @I$���L��n�3
L�l�����%$ID�Aē�T��-��u0A V�,�B����~���:,�)�/�-���n 4L�����g��}����g�<��~[������}ld��`�w���LC�����5��P:��'�p 2�-�NfX�g�堡�5:��� {�}!�.�ܾ����_Ny'�o]t4D[|��K�H�e� ���Ϻ2��&�N��+=��x<>l��Z�eyz��]�����Θ������[�5+��5��t<4�}©����R�NBb�ν�u+�k]H��w /tM��;���|9�ﾪ����cܓe��
H�c����1�MM��z�n����[/��۹�+ ��h�Ѱ�[f��к���e��R��2���]��OH�I ���wC������W������M���_Y��M�=��@%H�9�w����\����<a��Ө�V���C~����:��ݴ��Or��U��n&Ś��!�U�q��:~T��$��_��CǞ���~lQʦ>a���$�zu��� |>7�Y6�;÷vU���64C�99$�Xw�-��՚+B���E�{�<�c�z�؊�M2����p����#��㙚?e���Tݐ� y.��m��%dYR�C1��2�C�j_�9�kB�x�y�����5i׿	��'���w<�����]��]��o�8A�.#��9G����(���(u:��wM.���<�z�sn[h���xW� h��^e��>>���Q7�^0��ﾃySŋt^��E��nD�١71�I��%U�h��)��W0������hzF��Rm��]ݣ�[��@��9q=5;�l���)
A�X�,D*���"��X��QE� � �#U@_�7�I��JZ���}YѮ��ݑDi0�ZDl�O��U�K*n�"xy�&���Mv~�r�� +:�SR��-Z��-:�u��j�ĕЛa���� ��[r��;�U�����6&G��L�u(��#Ka�|�q���S�M�d�C<��f�bQ)}�"�B�0��^�pޠ�=��կ�>g�2����wk��:�V��:��в��B���}�{*���>�̅�\m�m�߬4��q4k�.����#=��&�s=�zY�Bғ[՞ke��6��H�#���\܅k�U�k�|������5��6���	����ޑ��nA±ˬ���r�Á�߾E��8<#��3ǮB���Tˣ䇷5G�}��Q7����_��������-�i�hx���`}�����]��� .C�rVd�(����>��*}֩��z0K�����-,{���B�
��9*�2c���1`��U��^�F�^Cwz�s���F��4Y�	˱L<;�8w۬�Z�}<���u�~$���!Y!K`UR)e�R���-��9a�&%e>�k�o�;>��ײ^^�zi��@�>ԟ;r�V+%�����	6[��n�bgRŉ�v)��F��;lGoN�6L�O����j�}Öb��s��##�v��i+� X�7�⁂�F?�>�����%.{�����~�G�n��f�w	$�(Ap��/x>^��;�H`���[Fi$m@��<ʵ��7��� p��iH�r[���9y��[�_���?q㧖�l����n��mn;9�\v�4��Ceח�%��OQ������č�9�tU�R���4!R��u������.눍8����ξ�m�U�������Q1�*3�s�X�I�0�tFkO�UQmⓙ2K�/}��E�wo��T�b�@�E �1T��QQ@b��g������g3|�n��=��T�w��퀫o3�1�Q�0���'�Ex�����	���2$�fŤn�D<�����[�(�������X�CBp"���U��Rt˫���
���>	dN�Z�ķt�݂��v�D���~�_�o2E"���O*�l��^TpV�:����z�R��*��T�cz�k������� d  6ʠ   ���������~�}�6��ێ�*��S�I
16����h�C-O|ј�'u����N�c�Fw�}_nZa�����UW���x�w�;|��R�>��]�$Y qӣ���q�8�Y}��[=�j��qW�Ey��z)Q+ơ-ѧz#�f�^�~����(��Xe��a/�g���U�)����z���_�ͤ�ؽ�O��ظ7�|���	��$W����d�I��y}�}��B��|vo�S�M�l����x��Y��`t!<>z��ST� K��J7�Ħ���))�9@�F�i�u[��+���^���|>C���>.�q���k�w���Gx� a� H�ۆܶ)����3]n���d����IyC���$	m)$im��(8
ECH�$~�녬��;�z���~C�!')<�������UU_e��Z��)3E�04r��F�[ĲF�̷g�W������p~t�W:�`�R+q�|���tL^L�(���&^=�Qa�uޕ⣥������;���px�e'� |a�����q��K���d�F&K�xo�{!���46q�?$pn8�ٹt4b!n�c%�}U��/d����3~�כ��u ��Q �ˀ|�(����3���!ON�WG�h��p<b���L^��������u���>�V�/ض�i�.F�]�����[��eG�K�Nˍ���<`�%� �[؏rq���Ơ�/�oE%{q�Zۧ�MWF�6��۞��m�k���n�m��RI$�H�m�2FS��D�p#��� ,�
#�PdEQEUF
@�z�%�:�kZ~O������AV�	(�:K���Tj�D��z����
h{�y�c��!���6�7,L��P���G��	MZ@����۹�t�8{���M���6�]�:g}�������z�9��HM�	!�䀊��Q@b�VE��Ub��M��r�Q�4�Պĉ�e�`
!�H~�}F�N<+��X���ؕ�1�+]���Ί�)�fƱծ}Jt���u�����>����ᓝ�Wtn���������=��{� �W�M�7��d�a�}��}Rj���}�����;c7��8���|2Ԃ[�oF�Iµ&��/��]/U}�����{m;����q��nm�t���Fۏ `0�m$�i&�Ȅ��l���K��z���m���j�\��ޏ�}��������m�/s����3]���;r$	�}7i����w�l1y#���KY��(����}��� �Z]��߻N����S����E���/NT:e��9�ӄ��{N��"K{��В��/���3>9����d�ČHȋ"�`��*�`� 3�S}뼈��m�{�)i�v�$3DkA=�.��ܧ�iW�6�A�v��H�ƽMP���_-�o23��c�l �3����Mj�_W�M������S�po�fܳ�;��%z�e�M���7�Y@�$��$��� �R4��Zz�v��pݜ�k!�jؼ����� �����T20z��B��Q>A񻙲lF�#����7����n�`��@(��$@'���A{*z�4U��Z��&������Φ�B��X�<��:y5��S�{��� �F�J|�O�#��۞�^�|�s���2��w�;R�b	���kr� 31��Jo=�W�S�UU2RɈ���w5���9�a�����u��;�9��Ă��XD�)$�?�SǨ^�:��_������,�[��9}�����os]��Z���q�S��J��m��m��8K�ڮ������|����]�*(�u�ث��*m]*�ٽ�ݹs]Һ  ` ��  
� ���������������+���]ʡT�*�����k>|��R��=���FS�ک�GeuS���ў, ��삪��ULӖou�]��[����'^�G�|�#�u��[�����6$��9��ݵ�|Ϯg����{[��_y�|�ʧ着����o��/�)��l���3$��{�'!
�r��p�R�9Ptwc}}���/�w�绤�Ē)�u�!��U34J�P�����-�tΓdv�����;<�_��-XӋ��9�;7%�m��Mݰ��?x�ɪJ�� 1��^����׳�Xק����u$�.ۍ'C�6�j��p̸m߼>������TdQb*��VH��H���3�*VV(��c�T��UU�*���c
�>��>k�;rp�eG�z��O��mf��[�J�o)i�C�ؾ�m��'��nm榳�f�_����P��O��
�K�$��ds�߾�����FnV���飨���.
u���Oxk�4.`B�*��rH������{��0Y �!��*���_}�9��������IW'La�
o9"�UL�o4�k�ɺ��%����r��Ӄ�^����� ����S�3ooRwm6'LC1|ԑ��m����E�G:{��8��x=�tӅ��hO��ڏ�$Yo�ѧ����
�}�������pw}m��-��I���Dě��],g����xk�gP՞����-)��v�h�W�f}��^y�������D���٦|���46��]]sE]�#-�U[��-1Cn��YY�t�������� m؊���_1UQ-��UA�ыj�J�a�kw6nc ���J8R�X����m�٦�y�֪5"��0-l��&	J��(q�J,�T�\��ׂo[�kT��3)h��1�� ��O�dr���'�>��c0�d�2ۉ��4�bգ�x���=�����hS`84iCZx>!���i���/�c+]5X��uQ����r�Ն�oz֪��\ټ�Zi3I��y�|38w^r��FG���,�Gݶ
 �3�*�s4M���f<�~�{\|5f�֙��s]�azP�G�7�~�g���G(�&������s(]\#��Ǩi�q�G�O:��B�h�����x�g�08xo�<��jm��FkY��UETAv��-�Y���۫u�[M���i��J�w��.v����b�"� ȳ8�(c�S�!����J��+�1���u����Dզ!Z�V��m1ո����ƣmMj�u�Fc�N[%���7���p8#��LKJ�^{p�ؤ'm:�&S��K׏�tI�OM�jK�=��!�!�����2u�]�����_����`��LB��C *��UF������l0��d�4�H�@�ܜ�������=�g= )�r�N�L�	�.�#*Z*�2K�`FGw�I̘��X���N����߉}����7���\/(�7��[V��D�U��ʏ`uʻ(�I>0��T�k���ӽо�^-}��;q[�{Z�+c3������ر�J��CxK��n�T�7W�M ��e����9���R-���������pl\��6/1�M�B(��f1�.h�S�q��0��ɱTߍ:�����̖��\`�P�s��9�̛�+��ޚ*��* ���jڵ�����j9�j6�v��]��G7R<ò�.ݧ\���ç�����Z3�U��E��je:�;y=��V,���K7�)�\)4�4N�S����Z���3"�%N��L�s9�{�������XNZO�3�:�}�?0�$4�$��݇�R�~AT�I4�'N���v���\�K���aw<����o߹߉w�S�	.��&�xɌ�HN�d�c��	�$�!����:�Ԃ���v�O��E*��y��o߾��u��gl:ΰ�M2]�1$�ֲ��}GZ��ϩ&ߘN=Iē�>N%a�ϴ� ��z�2Vx��`H/���~���~���'��C�N��ˌ���Oq��'~�q'�X,��߾`�d�|ͤ�'Y��0�������?{���w��M�m�ݸ�wW��f��~�<d�i��l��c	��S���i�ԓ9N��0�P=w�	�ޤ���I�'��	#<N���H{����!>�ߵ��������C�OU:�8��C�ĩ!�x��S�Ǖb8}������}�g>=�=��x�&�l��^�X�!�<��
}��B�N��7^��]���q�bn���B��G�{��&�f���}ꤢy)�P�S5_�{? »�?�|�q���Z>��Լ��]NU��\r�k�{z=8S�Q���q�֪�Z��H��m�PY3U��Fi��y���\� E4�`��N݂�f�MТ�)�������w�}��}
����'�콈>z�OM���P3Z�Sw��7~�����=�Q>���%6��v�}P��Nk=�g����^���? BE
H'����0F9��u��{G��{�ݗ�W=ޭ�/u�uxL
�D��b^M�]y���֮�}�D2����f��{�F���~��-�l?������n���K���~�w��{ԟ��*JF��
!R�#X�@��Ѵl�V�)aTb%)Fu��{h���>��#��a���zaL�������96W �4p�G��W�ÛuY3�ps��>���{ԼO���D�,�u��O+LM	~�(�n�
Rck �<-��#b�`J1_��wG�w�@-�!��]H�B�(�[T#)kPi ��/n����գ�o��i���Fp�"�;���͇ٲ>}����dی���>}�_�_5�˞��r���{��UT6�'����k�6kw*��bջw�n�۝�  ��T*�[j�   �:��ߟ����Ͽ�^�&�$7$m�fF���Lp��{]��G��6s�Ӣږ� ��0� o��ߙ�C	F����.�q[N���>��Yk���������A�U���%߽;
D�6J&jX���"��n��+���n<`�"r��OΔ,'N�F�*���Vy���=��y���PPUEQX,��PX*��DPA�,��M�1X�URB�V(��M�r�;����P{wӉ�����Ѱ3�鞙�"�ޗ�z���K̳|�Ϳ�̤�>X�.��y�_���O�=�'Ƽe��N����\�>S��u���9�_{0�D�Y򍳄_�C!�d`�ow����4��D����}}���b�5%nOl�]�Μ�0���������QrT�yq
�4�^%�!`��>��N���q���c�8,��]S�{-�MY!dП�?I5騖��&w�2I+�5^�xU�n�`2�?y^�eק���K1,U�����]�l��\���{1{��%B���M�4��)�����[Eߦ�0^I�u��E��>q����p�>��=�|�w�O��!XA��>?| bX3�Ə����y�����
B&����3��������﹟#Ó��ѪJ����ܓ6WQFH�ޓG��>��r��my�[&��Ա�m�=��[?l�dE*}⨾�ۏ��mv��5Nk���%�q�n��.,�!�ϒ��,�����79���
��vy5oUҺ G0c�DQ`-��9{wS�����a%����i������k��u�:«©��>;�}����+8�Y��g
khz#ﾘ���a/_~�/�[%�?xj��d�X.�F"����H*��u�lk��=�夻��Kt�Δ%�1�D�tJ��>�.�#�}2!�Tj�\�r8PWKԛ��I�n�t;kDh���ݪ4s�Ty�c\B��Q�_>�0G��E�gv��5S�ݖ\h@K�A�[t���0�;S���N�2�u�,�;���]"^Ag29V�u����P>�Z���z�x�������J��RY�������^�2���~�+����=9��w}xBx��  G��}��D{���8����=�v��7u�9n�s��l�'�;N�bj�P2r0�\<�R�x�B2(�m+���:n��l�J{m�����W��MY"@�G�}B�#��_:�W��$�|�C.�9< 66�;��ʝb�	�����~�q�>�ìْ7~�|w1�N��@�}�r׎q�>������}7�vL��?w�����6�2s�ϰƏF5���޵�K'��%�LԒ0qrlk,����z��Kq棦����  ��hyw����&B��Ԡ�bBe�c��[w5��An!���'~^�	�"P�Sg����{f��}�5��w���
�
H!!!����u����B�
*�də~���~�7��Β?n�:�o,+�O/��v�NB�d�h�ڸ�u�0ru���5���+�;�j\�h���7����5<J{2�jK3��t$Z/
��ZQR�p�{������;�b�����}[|��E�k�� �UYF��4�~�nb�\{n?z��^Hg%J�9ؘ�G9�u]x�&��o����X{��������f����H��ɘ@�5f�����m�]��S00�h�i�3�e9J�Jv��1���IZ�y?_y�n��(g�2wB?�|~�k�g���S�kz�Y���j1v��Z,ZS#��)��@��lz틐jhh[X2~�#C�+��۹��g�����  O����y����ٯ�!��ט�.�^����h�I˨��':���F2G}韅d��w�ݵ��}ﾏ� �.�1 �������:M-�ޮi=�f{}����"AV ��İV1# �ETDH�PDQ���QP���� �E��U��`������o�w|����Cs޼9	�ؽww��o��[�K��{�q��r\��w��RL��a={�N2�Tu��Ŋ�|�>Uk�J�8�fVe]���m�T�z׀�1����T� � w����w�w�ɶW�uv�w
n!$1�#��~�������Ikg���~חu&�6��b��w���|��x�w�>��e��(q���=��b��H�MI�U0�jY�a��i�xjH1��7
�"L
��dBF���}�}��m��?e+r}�1Ts��00����%tR\���A�,��yns��9fςV��W|�1L�v���t��u�� l�����:�c6�섛>�u�����ݸ�s�RpFI���=k)�.���N��sI���$�k�1<H:zp������F����{��M�
��#;�y%���\�z\��g?[��>����Ǎ���M���eOW���}$1By݋w{��^^e�ӎ��������y{��>߹'�H���""�$3����������W��*�c�}�}��OS�9ȫ��z@P�D��s"=E��>$I����1~sY�7�vB�!o���k~矼�o���9����r��Z�����g�^�{ l6�޻�q�;��I/م����nz#������6S;��Ϥ`��.��o\.'N�q�d��隙��,:���L�e4r��KT߇�G����� =#2Fd�"#�7�}�^������v��s�����BH[�cu�Z7�S�k�t�1�
��������ުf C��u/	Ǹ���O����G���j��Q3f���"����E��vb{�=�p]�}�+}���5f4n}�T˜^��*e29.���Xu���?���+s�{Վ6�M�TQ�aP��bI$���z����~����*m�@����4�q��l�w7	�l�	\�C��O�iKL�S�U5�
�����}*�Zr��)�׎��S�(H��~�����k��gX8dw��+[�(�_J7e��hQ�G�/<～�l�. �4Č�c$�M�������7� &@���(�TAQPPE��0b*�I�����~y���q � ("'��������b"��T�d$��<���w�os9�ꕂW'JI�4�ή@�T:���A[Cz��/�L]�ص��9��3t���r��]��ZV��� T�Uc�% զ�v�z�,�L�,��l��Ͼ�>��z|�zjhT��̞��w��=Ǚ�҉j�f���JQ�mY�a  ��\��Gj�<��|ġ0�ۛ�����> �ߛ�R��z�"i1^g�v�K�������]}v�S��y�䏷���OWm�B��ט�k���΅enH�����mʙd!gbFx�UlǾ�" O�ա�[y�`��"�W�Ԅ�W��s_�V���*L��/�lj.m�h�=r�Z��=,_�&z�f��T}z4<Q��� ? >|>����dB1�@/�~}ש��ݷu����<Mvѩ�~[���V�b2�H'h�.���n�Z:K��D��c�1�&��u˖�c��G���pr��P��=�ޯ��~-rW�+�@:IT�---
�d�Yz�w�o�����g)�����Y��m�:�8��ݼ�-(�|�9r,w���
���p��Hi+�D2�h�!QS#Я��7&�U�ߣ�",q�{}���>��$x#�nJ��S�D������5�v�:����ﷴײ6�*d���I>
IBH�x�y&}
�e�ؗ��\�&#qK�V�}��}IQ�.�Sk��(��ګD-{5	������a!5�`��(����-f�|��+.�)�Ν)�s��!�D}��0������~�=�S��ʸ��'!3H͹�.�t�]�~��-��	dT��q�#w�,�7]�0��H��i�!z>���U�"��2F��U�v�s�우w����tg���Ω��/��-2�zc�}fN���2��e���Vz��
�	8ҭ'���j�Dcm@X*20V ��?I�=W'N�%�j�lJ�ϼ>�|>w��pY�ͧdg�=��ԧsT���}��q���>w��]9����\Q�\�Z���ݦ��x�uWIq��]eĦYG-R��e�\�iMZ���.YUq���2�7$��a��`��Y���;� ��{q,D��+��kro.U)�]l�<u���pZ!Fo;��m(��c
j֗ڜյ�i��s|;��Wɢ��-TFڪ[ˈ����f%E40�-uL�m̴0�@�(��Gf}�đx��hS~hб���[.�¥�ʴn��������5�Y�ǀ@�I�!h;B7"&x�pz�MlyQ��l`Ŕ1��7�>P;�x��۩Kdj^/���᝸
YL�61c�[�I;����cG'ܳ�%��z&GZ��vg�������V�s"���E��#F /)�is�q]#�l�b�T188+sY���em((�T�o�ox]��u���V�T�� ��ҊaY�V��Ȼn�\�B���OS.�5�o�ym���L����-�K]�%r�b��J�)���e)SWY���)��UEuE%jA�k����r׷��$��y���V�G�-p��n��6Z���A!�
6�o^�v��̦;ttk܆�6��3�M�y|v���؊�5�!�����pU�G`�n��x�ǐ/T��]�{ыڱ��.�b���]5滯\פ�x=��.����B[�o*k~�S�SL8)�k�M;ׇo<��-�;��@����*2��o�B��.��j�{�E�������2���M��f� #�Ε�
��_פ$�{SE.{_k��P��S�ҧ��ǩ�����v����|������
��o	�ɜ<�;LӪl
�"�g%O�
�л	t��V�z)锍�s�����O:^*����a u�Q�1������O�v��6�x���c
#�we�/��[�{�Sar��~�l$�G�E��9LW�4����^�q�ʺjb�b���M���}	/���WJ��.w���y-�����l� �< �-��8@x x��$��﮻Ϭ�	w�.���U۴m� g;n���*��p�  �t��nN�W� ;��U@ s�x]��^��U��|���6�Y@ m�Nՠx8kj��U�D����w<*j .�vy��Uw�����ŵ�[�w�]zҲ�E�[h��z�ۻܯ/V���Ν�P��݋�@��||�<-��N�=ޅ��       x  �> 8EP    *�UK(    U �����UV��PUm�       TP        P���]f�ͯ���ޕ�{9~�Xm�W��嶂��ӛL�A�kU���8�jb�k���vn���ϻko�۰�mj��m{a���'�n�T�G�Vw^���6ն��׺��K����      [  @ x��_�?��}�yZ�����I26�D=�<�MW��ʈ���9��DD���z��MF��t[6�WXU|�5�3�u��O�fm�
[���\Q\�=l3|��\�� ��Y7�a�m�: ze]�}���v�w[��ܯ�<z�++؛�i�dz���4&Dl"=l�b~��M3V���J�6Ἔ��y8�芛szO�Y+����d.�CUt�L����	�h��o����2��*�r�:��eܳ2f�J^�{����!H�2F$	���s��^[�]N`��+�b�z!<HN�oB�[	����w�����n��L*���d��_�}��T��m�$n$�P���6�2Fۄ��b7���ٷ,�WV�뷎�m�dc�\�A}��D�Z35ݫĻ�!���������G�|r�]��c�(�V�"-�����Y�2�:������U�fMtn,e�k�;�o_T�v��&��o]ܕ��h���4u,o��\�Ĩ��f��ƽ��?V�L삩y��F���{����)Nux���ιg%-�5�W����yoG@�t����ǕF熮w�Ҭʼ�Է��O���̈�O*�VO���УQ���yh�f��u�Zg,�}�[��ˬ��h)�\����S?W�h}���r2�����_jf�f��s��i"MR��v޻ݛw�V�=��M�θJ5�+:���)�t�� �%n�^�[-�>��?}K߇��x�1��2r\�P|�����=���oMH.�����K��9`C�+a[��j6��b�}C���x��<L��iV���zl�O�8>�g��=ԾD:Y��[��C��-��{�͡O���L�aPt��<:2�����7?OC��݃��T�*˕�qF�&.X�D|}��E�z���{ѽ�W�a����[Q��z�>e�b^��b+�p�F��`f�d|L�̭@r���"4�#�)��5��}34�m(C(,W��l�F�ޙ^DH��6���ԐJ9q�aH�J�I$�H�l�$�I}���G���J��F�\�ޞ��'�
�$I����)l�q��A���i�dU=�]pq�K�4�V��	q%L�/�:YTC�W�:���6���4Г����G���É�%_�����\��Pm�Gd-�Wҝ1v���L�#�����-��nHU��|����������S�}��}�8��yB��'6=�C �UBI��F������ u-���X�R��vW��R�f�L��"�����RE�AUA,`����x���kxg���e\�(�։ZjI)8{ya����>B�����WQ�n��^��h&�Y����E/z5��
��x�ȑ�+���W��2}����W���84�ݛg\�����3�(�[����ﾎ���+���o^��%o;�m��*q�v��jX �;=�{C��4[=�����=�{����&�eoS�H)'��(5af	?]�B"#�,�t�[�s�����b1�*����?��_�� �U"���h����'�<�{ f0��dgn��lļ�[7=�x�r��[2��Bݸh�rI�߇�pd���]��X)K> ��ǢI���FԈ�8���sL��ZVO>\���.��q���<����'���O����{0l��P9O���3�RW��L�h��ɍU>G�u����e��T�uLLb{�;'�ty�EŪ�� ��>�#�L��������e+�oHx�
G��>��������pv�L;�񇀝TPS8���!�f��{�C������	v)�i�m�[NH���\�{� VS�յ��f���<y�e+=A�}u[l��+���0T ��`��   ������ߏ�ݳrk��z��*�*��3\��/�,$eD�ӂӝ��a�/�W�</l�	�Y�N�@�fC�6$f*���|�K�e��������[��Vug.l��_	S�x��id־��CY%�J�:�~��k}��r���/�[mp�ߨ��ݿ~� U� 3��>��½UO��>퟇��\���Y�y�{\�ne���Nqc�ۮ'ޢc�#�s**�(״�l���9�a6�+�����|�ٱ����ם�0Ny��&q�u���
|7���q��dZH@d]���Nrf�0�_US���m���w������6Qk�)���m��s|��n"|f�{O9��&ĒF�<m�����
�ݧ�\���wM�D�sl�y�hVA,F�T�\�: ��������w�耬���36|��(��]��ۍ+z����!�����@QV��Ai WĚ�|U �=<�G�*���n̜۹�W�HJ�c�c �����;j<WVfy*�O��`ߤMN[����/"WA�	�v*]�K7����_���}�GFc���W�t�7�!xGLɓ�Qyw�5
Av�״�v�[.�ݸ�[m 72fḒ��0�e�|#|��K���#H�����\�Ñ��ֽɎ-�?f�������^�t`Ó��[Sb�sx�x9�tp ��	��I;U&MȄ"��+���#����G|=o�|V8� ���7�{\����93[�)f�mw$w��ac�[O�ok9=����)V%R@�BF�eD�
Iq�ܢ��RFI�pFyqӺ��{NR�T�a��DA(޹�����g3�v�'�r�����K<Kg��~c{��%��b�!v���mR��ut�����ڹ�ܜ�xU��M��z�:Na�~���Pz��g;�sh]�A{��.P;/�,$����R'�<P~
��i�q��,a\�3������w���/��Tp_M�3�������`�6ԥ5�$�����.Lޜ�^�,��,�����7JE����UL~�Y��B̆MQ�9fo'ɼ�}��nO�v��'!�=jQ��>@�n���<��	 D�R0&k�y��9��Z��m�Ne�}��8N�F�	mA�Y_CŒ�ձ]xZ	���.9]��j����-z�mw6�p*�*����2G��Y�9�lZ>�FX�7~m�Y�-�d�{����݋|xkh&x"����p���Dg���2X�>�w;�=�o4����ю� R���>���Ѳ����'�X�'��ۚM�V��$�'+$ٲ�����P�KT�χ��*n�<�l(�G�ĄK��&Q��(�._���
��i�k|���4�^��P���Y!�3����߾�뛳�P$<`E)"2���+��U�+ �Z��0�aE�@j>������5T{fѨ�fc�%�7+���γw��H_[��9##e��R�o�s�^���b��}%���4�q�N�i�|��<v� �9���+?gLoO��m�ˏ�������� .p�T{�< ��x�{�vyL\T�����ݺ� 𪾷o^}U\"L�wl�\���T����'��]���h�Z���}��|�d���,3�� ���ܺ�>��]��?��Ƴ�z�ϲ��Lgm��tP7��҂s1(�yba�,�eD��5��AEo;-ӗ�����$��g?|H���{�g;ɟN�d�&7'��N����fI�.	Ŗ��<L��zy������:� i1q�������� ���DQ_}3^��.�^0AE���F��s:m<�����k<њ�5!l��:V�L ccN2�}���9�},�Ć���9�C�$cd��G�fB� {`N�R*
�^k�|{�Ǚ����á��u༛;;Ƅ��,����Cjd������7�j���o32�f`3z��ʪxW��*��yų�@z
{{�mf[eU��wn��ZЪ�벼   wQT
�    <����������U��ܮ�R�z𛍦�P2d�/�[N/U1��8&���������߸W��vI�S�舏Mϲj>��W�q�}3����`vK§&�8��@�(מ4�ϲ��:}��S��Г�b��Y��h:�#	�}�l���)���3�g�
��7��+��/��EZG8�#vYR�X������R�N��g����.~��+~��T�{�y�RO����%�U~��k�����`2�u�����,ƀ�S+rdۛ�{�NӮG��0c�6b���c�E���SFz2ct���wvpa[���l��U\y��aӌ�rp�,|rצ!��������m��GR�Wu��odV�U?wΠn̂���롯���#�r��:Ӣ|'�3&N@�s1)�yѦ���o�-a��Zl]�JjF��;�:#C
f{`��`ug�:���zgl��Y���s�b����O�T�w�,=�a�'u����|�[9�=����'�>30��Z�ؤˡ\�D�4[x���2�S����L9N��3q�[��THXb��>�]�O7�G�|}D���<�^��l\B��0�%����+�
��GLl�����<�+Y���iخ���"����Ut+�ġ��|��k5�,�E�
��ba�R�����9>��ӓǮ�{��:��;��������됄���~�߻��~�����Z�d&H ��x�H�I.EHAƲ��w�Vse�R���Av�:��Η+毢c3Q�rf�O:�3oi���<q(Ǐ7��#�����$��Ŏ^4����<�*�an�%&?Lz)wXs3���۾}�~���HO� �9��_̪����}?�$�R��0�,�c�6���������y�*k=��]�7��U5�r�t����! p,�=�[�#�0AU��4i�u����SF���5�]@9y㚃�8f��@�0`��h�I��z"�M��N��Sg${l!�`�ƙg4[{��[v�\����Al5�r�>Q�j^��z�~��効q�(���:�,[���ߗ�F�:�`�r)㩜=ff�w˚����a�4s`�&A�n <^�=:���W��n�7 ;�O�m��Lx K U��5�۹����[�JJ!@�<�bX����z_><��r�lg�����x>�����5|�h�9y�Z�E,!/�E#�����3M[Jð�^�H�M�$?a�"ŭV���<=�g���UZZk�Z_�um�e�A �[���~]��I~/!m2Jl��85\��G�0����X��
#"d�-�Q2�qV&Q!�}���A�uҾ��5��5�N�����w+e>�.��懼	ݺ&Rf��_j3Ծ.�j�6t�;މ���^��6��p�Ie�,͑�������,���s�ygq�칋���]�HY�X��e��lgg-���3ڦ���J	��;�H��+�S�g�ͳJ��̳ڼ�����rE�] JҫZ�b��J oW���w��G�����|TǞi����ι����`��rܛ۽�p'hO�_*�B��M���~�ë;�H�7�n�K�N�gvo-kFۑ��8̐\Z�3qe.�a�A=S:�g2���&���C��!o��:3��F����t��Fq�]q�i�b/����CE[���v��h��5�t��"�6��2��Z�e��Fm�mQ��vN�9�x���GP�������G�ފV�5���6��7�VT�q��V:��ޒ��;z�G�yr��[�uj+5^�v�ɪ�|\�:��Eq�.�ڃ��w�a���O�u��߉R�2I��^�_br"x��P����J��׳J7�4�*s�0x�r�/���Φ�W�G�el��5u&�QR�3}[ԛ˗��#�yO�]�a�j�k�i���
@�ȸ��aO�2���:1��kW?C��$�"�E�V
A��+����3���7U_n���v�R���+U���z����)�*	�L���ڣ��6wܛ�iVk8JS��p���:8Zr%�ޞOM<�~ų�����lz�}ޙ��<38jL��T	t�2m�#Z�\󪓞m�H��GE��t����lt)���G�ԝ�f��DDGӞ��Q�뺇*�����F�Sq��n�yض[:�Ճ��e�W: c,b�[���;T4+�����Ԡ��#H���S�U���j���\��>�y Ŕ�'���SrWb4�r�L�C�}_^|\ز/;S>EM�X��]�䎻fA԰�g����˽j����s]�W~�~��9$&�D�>f���, Om��3�;����oY������7+�m�2D��4�)��(��$��I&6��l����z~���x\;,�I>��R0��۞��g��:��3��3UH�tc���z�1�1Ȋ�9Y3w*ԁ���;|�S�
N����xkg����X�-��C�G�~>͔9?gd�w��uL~n>���ԽvE�����6+n���X�S̉�;�a�ך�x��r�@��X�1���uz�>^��{g:��UP�6��;�ε�d[��z�;�o���q�H���Z5�?/n��zs�����Wqv�y������G���I����0}h��~|�ϻ[���_���O'�So�Aɥn�_��-�|�G��<�F�b�F��e�  O��TQH(�b*
��=�;��=����صԨ�
ܮz�5\6kFC)�z�����!�F���O7v�Q��rI$W��sn�NoY<hIW��2
�-={��[|��v�vܑꞻ-���0 ��P0     y9����߿����y�9�e�v��TL���"8�~��DO� �~�9�n@b3I��E���-��<�_tI>8�K��h�طY��t�KR}*�}��o�iO�W�{�;����A't�t|O�1^���T�-��4�2�8���9������	����IL!Zy�6g��7�L�%u!�߾�^r����&�Ѷ������S*�͔���� |wK��s1��+�n$N)L�zq��sRs&c��<B>e����G��[=��w&�0�ih�N���F*��;?[tV;�n\f�]��"s��Oc�*�H��tQJ[�>Ya>�l+�?}G���VD�sU�U��H�I�#��mݦ�*;=x-�|�;�����$)�nsg�,��.'���=8mfӾm�͠�mщg%Hg�À$��| ��p?��Ѵ��wnZ�K���f������XC� s>����;�����
S�@H�{�����)Z����mf�Š��GD�Y,��x���L��]�	f:rc X��K�0�+��"�a]gW=Q�2mun�L�0��l$W��2��h%���dÍ<�F��ζ�$GW��}�y��9������M ��H7+,��>�r�R��nm+;��Ƣs�:�S�Lbŷ���"=Op����5��Fj�`G�ܤ�Z2F]�K���M&�]��	[�u���Μ����+��?8?A�C����=�-!r'�Y���QU�J(㑤�)�?D�m�d��I]X����&����>��@�r��TĽ�"��Gяq������I!?�L<�[����������<T�w�3$}X�*��N̢���sgj���:�I�.��5/F������,a((ڙ�L�������Ju�Z���U س�f��7���=���9�qz���U�0�,icE�#(2�(,cV���Dlm���K`ʬU���V�e��Qkkkd�J�lPU���N�Բ�N�&V�y�D�Q�8�8�ר��u,}[��.���������"i�4��e/Om?e�c�����s���?���xj!�t�:��VΕ5�)��U٪�(ã���Mͱm<i��[ޞ^~��q�%z��WtB��@̠l|� z#�I�/�}��jֻV�!���1�$����R�j�{�*=�[�K���7#t�b"������<��O��.��������M��a��o}�{w��S����{�I5\��S�0���\@0)��OMo��7������Ě�� ��ڛ�<'�����{���V�,�T�ĭ$誆T-����si�Z�&ܚ���n%�rEm_��*���������6=#�߂����D�.Ĭq{:�yj�zK&yQ}֞^��1�F�0}G�@>�~������ي������X�y)��E}�N
��K���&Ï^MQJ'�糷a.O�s�#��O��؍���M��2�ڼ����	PB������Sw������o\�24���3j^��v�p�ه�3q�E�Jyϝ�~U�-Т�]��m���STC���s��}��L7�l�/S�0�Tsvu[0�W��g�z��t6�o<���D3�u
kKA��ҭ��~9.�}'�
�/�y�~��I5�9�f�I=Fk&Q`�=�9�?j�SlO��W�z��~��[�W�ݳ$1���zA3������~�������� |��/���}-���i9�d�u��Ɇ��!�"�H���윪�&��H���}N�.�+�/���R>�?U]��\��d�yqm.W2#z���������p@���>n�3J	&V�C����s�Vu��� `8o�6ę,ĊE�>3��}�7��U�^s5�ڧ}�$@b���,
������?> ���7��:1�oU����P�R�\ϱ��:��
�����, Ի��7���[m�	m B��I6-\�\ʧ��5UUU,:����������iom׷}Z�[��� 1�Q� VR�*�   ���o��?~/ݳrkݻӮ��T~q�ϓo����u�հ<��-��B�"l7���<p�UXt�%]9��Ĳ�Ӽ����Qsi�y��"��t6�Č�'8�j!q��gd�͜�&��-���I;r�p4'�Uk��=��g6��WYOj�}����j�r�o��?}u��/���vPXnh��2��f�<N��ͼ��iN�kt�/W�i��έ=�L��Y���]�LW,O��aن�O�&����1�}S0�d�Sn�N&�f�1C�[���O
�����ψgK��qZ���Ͻ��`�EQdH��*�A��X���E���}�9�|7�~��1H���1�r�(���(�\]�x��U.�j2�)�I�RbDi'#m�$��������Q�Ќ&O�5T��t�`����{=v���J�Ў;<�U"��������yh��}�fv�+�_\� S@w�w�?l��&ʶ�<�jU�M�̜��En�:u<��&����i-TI���X	7_H��8p!��u�bT����DYQ��ɍ�����4��lʤUN�ҎP=\4O˅�-�����a�C9��Xҵ9������a�� P���3Ⱦ��/Gފ�c�>�cO��.���@e�ne:Y�{1�-zc��/���8�g_�g\�s��J����m�s爵�y�7��u��xvyX�HA�){�f�p�.��}τjb���3�%��]��x^�x��\c�=�+sܒ��6Ғ6�)���I	mF�$7I��x:W.VZ��߾��i���gW�ӏ�\��<�
�-fNo���Ҽ�k�R.���{#$|��Q����:����p�}��=�I�v���+@��rN����n��fcH��/]��{��bHI�awt����T��4dW��fŝ��s���.����z.7-PU���w�WD�=}�;P���)ӟ�F?�n	��������rr�����H��h�]m��*tEMe���F��L��h7s6Ga��l	w��\��EH������ezϮ�pMU	&؎:PB�i˄��w2�c���>zI��U��3ԥ���L��p�ѳ�<�o����{w�d�񴜆H�`�Ӊ�c�6ؒ6܌�T�di�l��N�V�^j�LB�gk���D�-�g�}���m��9�$Z����x22��HF{�Z�}j��>�w%�=-c�7^H�j�ev[�2�f>.[��6fc���V^5����Z��*T�*����v�z'�p��Y�iwj�ٕꮼ��Ώ'��s�=��^^V���}m�m�{�6�E:��ls�Dn����R�~������dr��+Bҥ��ndZ�\J��ۡݰSSA��;�,ǩ)57)I3�-��e�h���n[{��s|3ZX6����^��]��5jUX��������R�9ށ��vΧ�7���x�T7jܴ��ɡ'���n�On��S�g%5'���m���֕��h�lk���t~���l׮�������@}�n����W z+� a��;�:�Cu���Z�;7!<��Qx5�
w�Yz����2��>ktq�l�t�Tf`w���3%;foN�����;�^q��������t�{u�3{@0)�s֏�G�E"���f�}����;���￺z���s�͕=n�1�*��yGMp=��Mt=*b�,y�������W%:վ���S1�ٝт�w�s�f�,HBmh���ۆ&�ߙ����A]%TPZ[�]��[q[n8`f	�4.��v>V��K�������1\��e
($�<�AVqf�����F�h�Y�橎�����Yr�շP�/�7�e�/0��4Z~ �~ƀ�9KҴɇ�E�e�х����^�, ���EI�4�!����QK�I��5��i�1��K5���a5|�X#5��̏�����^(n 8ŀ�p��(��	�=��E�q@��!͚�sL����j�>�r�O7ߑ3⾸9zN7r玥����R�x<`T���I�H� ��9h-��:�)M7����p�uM.|�c����[��b��$�w�[��Y�CwGH]��E�������{�M=u��glg�P&��U@�;z᫁����ܰgj��Ѡb4	�vJ�w)��n3y���Q��6n�ݑ7,_ͨ���pѴ�G�/C�]�	sv���t�q����H�ݺPN6X٪�f�\�_W>ٟ�^��B:��q��2��"- p��3�ѳ���ɗ����z�3��ݱG"��=pc>�[���oXʆ$
^t�=���KIeM���i�U̽�ů���ී�<���v(��I����F�q����M۶����BϞ+<_���V3(��l�QN�f�W*�����I��0�v�@��꬚�ƽ��SQ�L\5��*�Õ6-"Vʘ��o,��y��f���&�V��O:t�B��[:����g{E��ղ�Y�=�뢕����7�Z��5+e!�Ghd�c��x2�h��{"J$��I$�8�c ��u�TE���޷-�w��8\�0�@ �ջ�	U�d[kw��� �p0� UwȪ�N ����wiU@���ǧ�Q�;;il�d+*ps����j�� 9���ڣڤ�S��wvVUU<��-�` w[zs����;l@65S���l�m� ŗ��t�[�Ƕ�W���6Pۛ�����^���VUl��]�׫��      �� U Ų�     3� ��    *��@�Y�7nn: �                     �  �:���{�g���~v�Z�췓bV Yb�ȅŽCE�Yș3���(�n{�e���W����m��7s^�T�[&	6<h��=���ݭU^+k{�T[l�2��;�  ��  y�    �������������Y�[ͩ�lרUw�UW	�pf�Z�2V��v[�V�+�U~�6}%��Oձ9����e�����	�����QɌ����g�]X}PESfr���:�˷Ԭ؇��̵]��B�z�Ͻ}S����ΒV��
���Qq35$�^�� t��c�˖�ib�,��(���|����꘮�LM��lG�_}C��`�3n�7&I*b�[�%r�tu��������oٮ���]��'�;��i���	^vE�N�cz�Ws��Y��� �5��#_�GL�p!zv�*�����No�S�9Rl�	��p��Y�-�������3~������w���kν���W�+\)�!=�#OrМ��������b���;X��!����Wa�z����%��.�|�q|���t�&H��wNz��_^ݾ�~�!6��1H1�Ӿ�yA����r�ꚥ�K�H���;��Pf�r��u��$���b�ם}��Y�a��Ƈ���U]*O�� �W����)e;�f�۽x�B� o9�q�C4�2YB��gd��-~쐟�"�����t�ֽx���L�@��q���<hiZ�\1�e�Ie�7����qC-�Cz4V n�s������=�v-t�S��*�e{{	�bcu�̽q���݁��wGDa٤l0�mG�߸��6��R �����
��ϣ���&,[��Vw�}DV�﫯j�_�@�`�	`2K��d�O�O�(��qS�qk�����x�xL�S������	�$�z�λ�,Ɏw6.�Ɓ��vW��2F�ܑ���5���)vv4�VVۭ�'���P�W<���+��9~N�������׺Y�Ib�jl4Z�~��}Ƥy[��}RE��s����o{��w�^�\�NT� ��Xõ����f^�Z�d����M�56�9��Av_t^��8^��7�>���~��ak��xz.�c7�W��NG�c�u�I����|�#
�.����u���dGA�غ���� u<�+���'�#��DW+�~�yddצ^���I�}n���/���S��zݻ��8Ib(�{W��彽�!��:��q�,�|��5���w�#�j�S�'c�2j�*�8�nR�d7�+5M�@��u��%�
��f[Ν������|> |�ͬ�����,m�I0^��{s$�]��3K z�Y���=��~s5�-7<*w����
˻"��`��rD���/O������Ɍ��� �����D	mc�SÙ�w߽�`%�����w*QB�A�!��W�[�����yf�܏��x�y��IxԤܜ�Iծ�n�uURH����¸�B}�$��]����n��ל���{��S�<�o�z��X��V+��0��������xB/	M$l��i$UL��Q�_Q�1���[{��Q��ib}���~��5���ݍJ�MLu	�'b۾� UP�u���q3�N>������q9�$^]��EO?%UU_g�3�{���r9�C�'�;}�6�L���k�R������M=��_{k��&�t�Bd=Y��ӝ������LЪ![sw��w/k�����j���bln����s��R�I��9(�N��DM��k�R*�3��D�8��8��]��zs�W�;�s�x���� c$$D����	�E�u����^�3��1mU�xBU����.�x��t��lk���ۿ��|�|��S� d�����<J�<�ܭ�5 w{�I�*��z�s��� �  ƪ�P   w��������~��zֵ�f��m��©��Ҧ�[b�o	b's�7�j;��ټ�镴�0W��	jo80E�!]ۛ͘�#�*=��~�:�}���[�҉;����(u;����N��t.MM+���Y��k;K��+���p�V���Â���ߛs��+"V[#��q�u��Y�9����3�?����~��~Y��L�G��AE�r=��Y�o^���a���]�-m���B��/�`�Ԃ|ԬUo{Jz��*-�ۭ����PS[<������3&�!�ZRj�UL�����T��3��DDG�D}6x�}�3c�Fo�s��`�",���Ċ�*�Q<�(��+E�Li��z���Z���e{U����#��5hb<�HqX���ʽ{N=�Y���y���n]��ZVm�	Z�n2��r��@�Owӑ���	B�2՝�Q_��w��́71ʧ/1��*�3�}�3u��{hI�l|>s�/ʻz���}���E�T�\�w�zyk���^9�/v�����N$�����l�z��K�����ϸ�v+���H3�ȫ��i��=��Ң[�܂H�xJh��4�I i$�L�HG���.j��譝�Ř��rC�*���wy*wݘ�<ڽ颜H����j�@]ϔ�`E�ܔpVF����|�{�z��ݻ�~ӇT٨��d��2ryP%������_F��#�"��On�wlwbr�Z�dZ����=Z"Gx��;��M7L��&�&�ٚ��iIn�_N��S�yz=��D@x�oK�`�T��v��>�w3��׺�8��^uw�����ϫ�~R�����q�!iܵ��%($���ٙ1P�}��v9O^{��kl�le-�Z��}�R�qW��`?}������������vD�6�>�ewxU9�C�	$��!�����>�}�����:x﫽��)��r�i)�+��Cx��0��R�s��,7<^�-��QYPJ�>���s�y&�)�]~�N�4Ù*����ߟ��~����Hfk��Π�s�t������j��H,���b�^3/�\���LӍ��G^�z�(���'4f#O��ݢk9�w����ݷw�Uވ��9g�j&��������9���bO9��i.<���n�aO��f�i�~���%��*;vp�zg��"��;W�.D�ĵnS�}ߔ=��Yɒ0�:�G�᳘b>����ݭ�?���-�n���]�(rFܦ�'�����z����=��#�WV,�����SN��E����|.@-+�G��B��']B��|��I�t�_sz����e��}ݭj�֪y���I&��]����+V?A�K�C�����{u��������O{��:�������* �֪�:n���`uF<����$~��3�3�o��U�{��[��^V��hP��"ۥ�^�s��|i�G����O% �{o9ӭ��� Y'Q����5��s��y�ܽ���AV|(�>$��r�E��,�������n{��v���Q�b!����̻�:��������l(�m�E��ƒe��޶�����<��
�0Zg�^;��M9�:[m�FݓǔPc ǅP��   ��v����~����R��lY�tV��U�S�yX��1B�`��ՊNم;m>�j/P��]��-�30���{�D?zǕx��UI1޽鲮�����!��G!��\�:f^F�Êf)��|�L���eҡ�z.eD�6fH����c��;vv�75KA��6�t��b�L�gB�#nvrm�@��5'Zc*V4�>[<�q�`<�y0q�_r}(��-��ԍ��U���qNMo���q{8��~~ ��}�����_/{+�V(��;�[����	�;�OB5�5].���1�6�۟^���gp��Y�������:��6�uC��E�������p��"�
���'���(�����Z��7߮�$ąV�����=<��y��X�����GA�V޿(߅��l���9iO���KS3t�ٍ��u��~����p��(E����"#�~������]�<Y�����w	g��Qa'��^[��W'^1_^��+=3��<��Ӿ�gѾ܅�^�H�}�72w$�=���z���<��`p�2�]j�;��R�j>���u�Q���b����.5rR����ș���}Y�]�7Zr�����t�#UT�U��ө��*}wu⻾�c���|r3��,x簳���W�k3)�;Ӎ���w\��:CA�|܍}���~�����{���X��}�϶��_��6L���h|nu�֦����OomU��[����z�s(�Ԗm��	`� X���Xj+ , ���~�#��a�l@�$}~0�Qcc@�r0AQ�
W*��đCE����{Co;�;�6��R��a�4Ǎ���2i���8O�h�?eg=��R��}���*��1T��L/����`�E����%���.�w�<�����slVHX�q3Sg!�c���>7�@�2���e���y�Ȏ���B8�<͖�(�f���:���w�|;k}�5OyVDy����mw����ڱ�6���ާgI�EP��ћ��MZZ
�c�-*��Z��U�&&u��en���N��Z'yT�gƓ�������]�������"�וIں6��6ĭa�Ff�o!�,���X��[�K��0VU��3��-��`��}��/uͥ�ۊ�1w�f����oyb:b��5�A���Q�y�{W���o�L̕�u�@���L׳�x����A,S��zW	r���na2��I�[������j�R�������qb��l��|�$������yC�1�ű���#Eȡ���Gk3���T0V��X�V�u�ǬE'sp2�㍥����,c	�"�d�@U^?�8`�[C�����ϧjٯ>)��_D��2V+ޣln�yҳ2�Y��n��;]�2�����t�"���d�{���2,�[�w�����RFͺ�m�Y�����j��Z7X;�U��:գ����+�(�J*H���,�	6���T�r�2d��o�b{60*Z�r v6y�{��w/Zn�l�[��5c�毨�2���9�f�3�ND��5�/J�y�0,L��OWb候m�pO::�n�x���q��E����B�������'�P����NU�7���]���Y[���*M��.d^�y�}�������sm*�$�08܍Ģ��$��䍷��6)?^]-�O�j�fOpa��3�ɮ�x��$�)�{VOjx�05�n�fhLG�}Fϗ^O��(�D| |}Q�^ǭv��;�6h��^v�	��uvtacԻ�m�������?s�����*��i'�/.w��D���m�m��9ݺe����$fe�*s��k�_�^�T�'�ea�E}V�'�z�;�w:^[��">G���/����dN���V+�"�+.�Hk3U<M�Ӌy48T���]���٭[���n�B��ѕ2d�ƺ./���갵#��\���Z�6�z$�Iz��[�GQ�t�~�-��oO^�S�oY��B�������G�ð;�<V]q���øs�s���3��x��I[հ=(n�|�
���Gx:�J�k�Y�6�L����x�9;�K8{ٽ-�6�3~�y���H}�D��UP�TŸ	Y-�*Y52�8S�S�7�!�oͧ=r��.��e�����@��é;ʻ�ӓ��m^(���(����������|�$`�x6�7�D�Q�TML�Te��^u1��y �-�r�Pg�Φ����7��X�ꔣ���W�(�P�U,�lDZ�E�,����R�*UVV�U���P��B�UZ"T�� ��s���J�"o�j�ve��ރn�#��T��fd�Β�nvmo[�������~m_�]U��z����l0P�x.;���k�k=o���^������ssR�P *�;� b� ��I$�I$>k2��tLF��$�"�H�e �i$�J�H��!��ϭT�ɼ	Ǧ ����U���}��}�Z�k�+Xy����=�yv�T���޵������|��N��C�;L[��E�]���<W(�f���[*�b��"ha~�h[�,Y�Ewmܿg���M�k��ӑ�=��q�}}�G�xⓧ�?�;w��7_�������%C;/���˔�Kr�=[n�M[�k�j�3j�][��M�RF�s5L��}��X�y�"p�=|�<�p?h���|�r�,�s�;��%RG#�E�B��U=���]���/��������,�W�У��V
Y�{V��f*�r�^�eg]�{p�8��"��/��s~��$�$2@X9������������BSS�rr���s%��Z����/	���wg.���%y����*�:ۉO�w5<��7�fi��u�����1��URD���J�Kދ{�*�	��g�����.���]�^�	�	;�9-��hg���$v���ֵF�n٩���~eq��&�%�<=�-j�9�雴|QrC������ �m���Gv��Z[��k:ܙa�����C~������G���3��4�}��ě#���yw�u��8��
�^���n��~�:�5���{�^����
��ֶ������粏��3���>�sW�+2ww6��c�ՔB�����oQ.�pc�X��d�0o�UUڝ~w���'���I�C*D~��uO��q0�_������9�����HE �QAH���$�}w�o������}޵�uŀ����h�[[shXL�*0�SFt]yQ�����[�x��u�w!IѶp`#[�8�ے�gI�=�4��a��=Z�dɝi���T�[���E���U���'O�t&���[��'.@��-+
�N��wX�.m�y� �z��[��$$�_w[��}�{���}C�˂�G�3�n�(05NON�O
��]���#^��ݛ�&�RH�rIu]�l@
��no������6�ʙ�b��	�T2�K1��i˾Jw�֢�1����)��ٕ2Dc(�M����0�&��P\�Wn����O=2��H@r��`�n����~,*�����ny�+/�޶��l���t������KK���ob�?F2������VE,��d'`h�R����ڽ��H��MH�;�8P��^ge��>���w�%9����;�%���ƽ�\XE�/�ץ 	E ��`���=|1`w�ta�w��,$�\�������*x�y�9�E{F�x��������קc���A�M�>u�s~� �0�������ǐ�| 	�9���Zb�J��/ka��0қ[1�M=tfgZ��u,@J�{���4㑴�
F̈�Q��nCS��0�M��������weײ���z�Y�\��Y���ؐ��`��^G?����̦�s��N�en�7�KM�m���^e����H�DT�#"�,R?�?}������n�S�=���u�z��V]$��y�X���m�5p	�P�{�m��:��	y�<eۧ�m����j����u�g,�w?j�5e@{�����^L�_��[�{�^�gFa<a�J�.Iۙ�$�hŃ�nl����}ٗ��[�p| x�gF8ܕ�M��]��ơ�z�A��,`2_w��POa�i��XKw �1-�b�7�<.�J��/�q﯏�޿����t�{�%�y�x���Z+p���8�J��r�$�.t؈Θz�`�����u��0�{{S�K0u�ʩlT"��}*�ʩSns�����R�Tݫ�h   �� ����  ��}*�76�즛	C����&�D�$e�m�Dq�M���I8{2Gd��Tb�L�,3��]?,  0��|syZk���*�g ����nZS"r<��Y�/9�>Gω	=�)$�O<�~�����f��ޗ������S;�ßLjyTT�s�Y�����<R����-��th�e�&���Ey86��h3�i�����2$�1[����c�==��b9����|R�x�"��>�v�@�P�/Vbu�Q#`�2�GPH��@ ��<�j�n/Ly-��b���m����;���օg6j;��!�,l�[!�鯃sy*��B���uu���od�a��9�`ؘ��@�`�2��˛��A)$*7 i
-D�H$m�hF}���~^/��{}�;OY�ƽ��l�t[�I�Ҵ���?c�UA��N��e-v�F�v�?&x�=����VTΝ��S�zX���������;�6��X��l���٣����E�!q��sґm�\�-���=�,/�i#h����]m���h>�(�xQrh����n�eY�
��UF���\��F�glGϰ.=9���Ē����<q!��-��1��U�d���#��Ք䁺��]5��>��G6)�ɍ�s29H���/3sZlh`�ܢ��B<�wX��cKڡԥ��7�0(�a�Q��]?[�8L��O������
�F�+�AG��3o�����G.�sfe��!v�,���r��T�N�Z�T�QV�V$��m�vX3E����[3�����.T��mɝq�%�D�ց���:�!+�S��w�אm!�pbx͗���^�Ѕ'!0���rto�D3��|����ګs�_\��X0*A��<#:Xl[�j.J�"}���g��}�g�fu��I��$x~�R�W*�L;���=����j����QˁT�v�n�|1���gE
㲕S;e��t��e���>���~��=E��%}m��>��s��������ԯ��^�:9��tt���e�Ы�T�o2A�|p@]uc�.=:j�bi�����ʨ���S0]�Z��j��CD^+K�7�8|���K��G�[9U���.�4��9`�c�Q�m������ �D����b.�����:���5��{Ț�%' g�.mo,k�'I��t^�=��|e�V�^}�4o��	4s�u7W��:���D#�<�Q�0�GL��ULň�K�ltu�ı���ON�z�&8Z]~0��(+]x�j]�3���y2���!�pm^�����g��M��Ef�E�ݎ�2�1�'�pɱ��� ��<}�;〪�d�͊����u�̤⎎�ܬ�(�O��H G�=��!�w�:��V�1[8Y�����Q��c��=�a�}4�'��)S���nwxy��0V�f
�eI@̰vi#C�
��'ur�-Ng�N��U���!�{�	,1��&��M����߇ݢ�v~��j;i	�fڻ�o+g �U?�^���_�}t煶�L���5��t��CE�i�cb��^7��x�G�p�N�OK9�0�5�R�����m�5�m��ىf�_��i�8zb�ظ����4��v{)g��)Q4��Snu$ʧ��:ِn5lM��#�c��{m���Ɖ�<����0���y-�M24t*c�Š��~�؁�p�.�m��6����K�ᏻ�7�]߶��Y1�5'�i���+�Y4�a̓��^��䯫Sog��f�
K��>f�]�����46Nӈ��0�����a�Y�����<>�������4lxxGx����!�W���_�h$� ��q���I��^�bfc5��jWX9Q.��R�MQ@��*EE2b�d`�C%�N\��j\k�Xs>Ѩp�����y�M"�������N���i��M��CSI��$0lj���Mar�-�$�=;��[� �ˍfah��R�#��YU̄��$Z�PFrIC}�pnYnp~���}�<˛7)�>��(Gm�!0�K�Yj�/<9�7|Ɋ�//�NEM �&ʊ�w����8y�r��!`?SJ�Eܼ&��"�+�<�ί��s�7�n�V���(� Dy�$熄r
��9~�=��g��%��7�̈́H�����aܥgUk7�f��s<s���/�����C{A�/�W�͑��nO������hK>py�op]]��&!e�>
��Bh�-��Ǉ��̥͗Ɋ*1Tn\qK<ˡ��U�YF�AX���
�馛4i��q�n�b��Q�&(
+�T���21����H��|睠�-˪>8�*�ͽ�ik�ΰ�%b�;�\t�&�%�k�E�N�fG�����l�5ay�.��Z����}�5�w���Y���Y��Nԫ�sdy4��.e��b����<�k��0�䇏]���V_W�I�＋T�`7���sdh��[��D�x;��[ů�m�}���ߋ��d�k��i��7�/_[�9�8���3�w�Z���SVx����z������v )+�{%��\��M�8��V9d�A9t�ڭݧ�Pa�Y$�k�l����ظ� >R�{brW۹]�:"�^�߶��+��+�h���^BZ7���}XQ]Zwv�����o;B�0,-m~o��B�k�^�<_=�[:��y����"�1�z��E랑��5|o\��|��F�Q#s�U�ㄇ�O��uo����MդUĖIh$[m�J�U ��,�Ez����Uny���޽���[/<ol0nW��ĜT�������C ��� ;��M��� ���n� ��z��x�[<���`P U
���V�*�ܛi�P���������guKy@k���V9��Ek�����)�;s�֔�mlUUU��<��zڭ�{�mmjm���}l�5� VV���m��l�=o6��� �    @�p0 ʠ  �     �e*�@*�UYF��l�K(  U     P*�         a-��m�@8��A!������LPJ�:P78��(i�25��\��-N�<���g��15��%!Ͷ� ���F��l�X�G��+%�7�{s�^b^oj��y����.c���8 �UP�m�   s=�ߟ�t�����)1�0�d0�m$��6܄�Tp�����P�X��#N��$��Y��b��n*����xݤ�n�f&�};'�:��0Q{��2��	�0'>6H#sem�e���j������Xjh�B`�f]��=f6x���� �X)?XR1����߽���������ˊ�Á��d�J?08�=ƸĹ��|�+n�]�O����-e�m�w|T#rx0�".���	��G���_�5x����JP�R�����Nd�(���0�������u��R6 Д��Y*�G0��A�[s �nu�t%��;���'R����ưh3�]���^S��I��1�́�R������Z���i)�y��]�m��	�Tp�k�s�#mn��o\Q��>^��<3�Py��2�sƤ���;�W!�����9��I��}�{�\�*��ؼ>�A?� ��0R"�����-��i+U�P,�6�Kj2�b�
�PDcV6�+lD��_|	�WS3������/<.��M�5�g#��Tt���!ߤ��S����ι�Z����6��ս��Q}�d �s���G�t��,�$��1`M��]��]��;e�P�UZh.��H�0�@��CZ�W��4Ζ��1g����[lWgS��a�-�f%������\�'>FR~���lޥ�͋�,���=��wW���
f��Wy����4��g����~��2�ͻ=�:)D_�EW*#�/�yp� g'?kc(�5�~���3��%�QzU��
Q�uڞ.��߽޿"���w�g �*�-GL����/��Z�I�ڑ�I,� Ʃ��[�������29��)������L���4��r+�WH��_� �?k���{����3�۷����00!�����i��L���֩�U�`\;f���1<�Q�xHa���Έ�����DG���DFS�hޯ�5D
�t�Ғ�
��:�fw4��W�r0�ࢉ��2;8��0=a<���1����5�SDX��m�lF���1#pVb�ք����<j�é.��W<�|��SD�:���~��y󆽷���ewi^�OF�J˜%��\^L�q�a�7IndwT�R�[J6�w��.	+��j�3�w8���@��5��;o��%X�JCI�D�	�bHۜd��*IK�%fJ�b�	b�!���A�	�&b)�\���V ��wsr�kv��z!��y�?�ha���x!�=dDW�sq�N�2��
���W;wv�s���ձ;��׭󡖤��h
��p`���3�%��	���`25ݾT޺˛����B��C�*�'Fiz~K�
���q�D��n��ݨך�J��l>.�1�%:,X�>���+�H�� ,�I���������
�+��w�~QK0�Z�cqK]d ��S\�F�h �k%��ǫ_`(�qs����L��/[�/a"4j4OR�Д��L-�tan
�|��nz_���Q�
�;>��+���y�MWI��f�W';��\�=��'��ww`��ҾV��ċ!w�KZ@��'�Z��ㄷ���a�bE��Dο�"#��*ջ�-�٠E<��|#I��[�M�{ݾ�19�-l�&%���!���r삺�Fk�(���}�08�/ž�{�o�*\J����H_����x��.�>���L(�͓�Z`�D��KN�e�ב��\��/s�m|��Bo�BT���_���j<Y�������7�զ���z&r�9�ȶJu\�
�Eu�5\�?U�ٛ��k�H]��{C&"T�I3�1����a	�*b���F��|񧾚^��yr�__��{�(�l����8:x&���B��\n���r�I�;����ˌ嶫%�ۧ�v{���k-����d�u�/�m�m�Zm+B�C� �S��V-�m�6����D�s��]ݳ����6�@�@w  ��P   ��_}���������e}����U�v� wLb@�y���8Q���C��\¼G����:\�wJw�US�|��E���"�����'��f�T��#rz�1q:w��n?��I߼��T>h���«q��Ja���f���B�1:��^G?���
r����gL7���<���;nʳC>�-���ؚd�c��}է��ik��X�&�]���K��=gP�U����=j�lp�.�EBԎS�Q���/K�;��|�<;���E�8w�o�Q�]�l!ƵB3k,ý��X낾'Iʘ�1�{iЫ��o+�}7������z8Ȥz��
����G�����I8c�B�A�F�Fۚ}�W�Q��T�\��□����-��]
�X�����7)P���ysReR��+4lvL��kO�ע�O�Gb">���o�Y~yV���Vb�7	�,����m܁n��9;��O-ײs �]�\K�w���%����i�]�E�P\{�wb��h���)�GNF�v{�@�N�]&���=%�#D<1�}��S��[�'�Z��oϳ�M�_�z�7�-�9ɒ��3���r�$k�{�;��3LT�0��V���V�a���ۭ�4��<"q:S4�d8�a;I����'Y<i���UWS)�~q��oǨ$wA�����ߏ���=��~ÍFj�#��?f��9�ѶZ	I�J�"䐶���Í0d)�t\\y��V^hF�BI��[0�M�s���Ǎ기ٵꃰ���Q���^��>�$��!��w$R��K��kH<t$n���Ν�Ch+:y��M-��/�Nr���^���"�~x����p��ֽ����b�g$G�=�܏���� �W����L��y�-�B��b�k�v����*�6���+5�Yu�¼�L�s��zuz�h5$���ܰ3��ǵyӇ��c��l�oJ�F��쩮��{i�B��Z7�ԭ_x�.�����w�й\��j��vP�<$��m ��1�LX�S�2�M
�b�ﾄ4b�ȡ��t���8\�MK���,e7L��V�gj���I�m�4#iȔND�{��*�Ul�2���������c5���6I�����oP�瞩ֺ�U^�(m�E�d�N���c�[�a�#��dy#��_ճ!�O"������)+�j��W�ﾦ�L��~������{_���&}�fZ'U獻��j��X�S��j�׭�{���`W/�]+O$/ƹ܏�s�q8g�uaII��o:]y�����&����0�z�WT'3�$�a8_��s� Ad���+E�P�í`
�Z�`�	G�S�]7ꍙ��]զ  ���m���XAt��lG۸��[����{�J�6��jw��B��k��i�<��Q���LI���PЇ�g�kך�>����Fu	�B�V�i�\2��K���,ۊ���]�}�\Τ��%#��$m��EWp�{pW�}��{>��d]M��n�B�;�g`m�Dn�u�O[�\�]]���l4H�X��ʂv�J����ej4P��c��7}�}��� ��U�R�&���$���T�a�E���-X�����%��k�j9�İ��[Ӷ�-�]�������/8܉�M�OEL$Nz�*BF���ީ�䮴:�H$� ��l�2
H���O�9��&llụa!;�r�~�o<�h$�$P""�(��<~�_�V�{����΃ٽdv���~A*��@�����83�l�߄��a��z�Z�ǜ4��$[�B�H�������f�1��;�w�Y�t;�عb&m��Ner�ge:헜��lK�ի1c�l��[xU��uUu��ڞ 
��kʠ�9+�O>�y固N_Y��u�KxڀU �  z�T   �$�e��g�d���7��>i$��đ��F"�M��r���ec��<�^}�A�Xa�_��%���gD8��tޭ�H�h��C꽕��xѯ|  d���
��4a�K��OI�:�y������u�4)��"��͛�7�xn();��ON$r�bX�3;IEiA8<c�w�=�G}smO�J4��
m�}-�b�vl`Rs/����a��0�*fbXZ(��o���v���Ǐ9��.Ы��}��o�������(��+q:��e��lPB��<4��s���E���R��˄�N�!Z�qͧ�M�(:��L�<�cF�&�#}.T���w�k��h�[wn[�� �U������=�y<E*f��S[ֻ�,r��\�V9�)��&�U��}B�U�V�ޚ���G�q��NKA��xeZEIk=c���㇮|}��,����T�����������DƤ�/"5���Y�ר�"�9���C�4d�Ƿ��J�����oy� �e>�g���;3�´T�ݧq�ۜ���g����C�ZL���]�O���[hq$�����ѫ�Q��-/����x�R�q:|�3�t&/	2I�����H�4�9���2�*tg���������͇њ�GI��2�Z������i��J�3�mJ%3�-�:�_$j��c��$hn���!�f��s�sm�|}ʑݻ�5��܎6�rާ�d[w%S����\����}��F���!��@@�%_Qq�����uԘ�wT�`���K\#{��9˜�^}�Ѡ���Lfԃ�:L�@a�u��ci�,]��Lf�V���H�����7Ҽd��{#��'���3��ɤ��3�:��w�/-�Rf��õ�Ti:#`X�$~P�!pKȋkG����v��3T6.�9�j����[�\sTiQ�qߗk��ᖅ>�8o.���,�$UUP�lv�hUb2�@2���l��tQ�-�0�Cz�|�F��^5t��Q�1�����9��s�gZ�i\��)S�
�,���2��3 ��Θ�m:�ßFM�'���|�kՈo��4 �|�Ҕ+x�ݜ��,�Fȁk5!�Y�x4����5��+�<�� i����X��5�1��(x� ���g|-�X�π
w�Qn�w���#7ç\ys���;����ހ3�Wq�sÕ�75��a���9���BZǃX�ϣ�<��AU��s��<u֣�z���_i�
H�P#30�c�@L��e߶_A����@��Wp�� ��i�-j�hDfQ�b�*�b¦�{��7���r��ѣj��Q`q�Xi�fVb<�ɡ�Z�D1�ܺa�wnG�U#ƃo�ӭ��dݝ��us�|\�ά���72�輪��(B*fGF�/�򚷄�
&�׽!���w��%wjM7�.;�ˮ�eJc�'Y�d��kJ=����3�F64���;��|}�:�S+$o�����e��&��&V�<�8�q+#�2�6�/_m����y�)F���+Vݽǵk��7�+s�ί-{)�K�%����㭧��%WE;�ڨ�6^�:�����-�����[V5�Q�@r���B�scKa�"o�Xƺ����EVwn��5z8lm�Ǔѳ�Ⱦ������ˈ(�+��}%�ڇ��rnŗ<�U�L,�b�7��9J�7��ھ��:��N�Ts�ݩzx΁�|�����RK���8���9!��S9�bt���m��|���H=��o�����:AoCâ�r�k����~�M_��ܛ�1G[s���wy�bi�R��}��y��<{lL.23���wa�����9U���&g=�I�&�Eԗ�i@u!q5�}c��W��rD�������e�Gj�q���t��<���Y�\�Y��QK%���t���q�&��x�����޳i�'�4��p�+�a:�+��j�b���8J��[��C2��P�Ķa�mq���z�����I�!�8���!Ff4đ��l�F�����}�@��8}#O������K�Q�9E4g���{���K�IJ}<��WsF�}^o��#�HWuL2zKIߎ:ݞ�D�Oi�(��ɏ=3�O�M!�D�:.#{u���୦J;ה<���x���E�yo��k
�x�V:<#]�ݪ�������3{�{WM�k��l&H��]~#�&�����|���3��kخ�oΒ�͚pE\�@�>6\���舀#��3�=-�7�	�5�+�m�d.�}α����r5�O1.t]�"g.ĭ��$LzY��i�g��*	��2R^L=�P�C��A�'e�绥��~^sP��ܮԋ�/�ۓ>�����x`��>����m��zM�㐘�R8I�I$�#m�H���l�p&*�/%��.��~��Yl#�"��u�{\��N��ѨGG�U��^_����o�\O� �	�2(F�bd՜���Mz��W|^�׿X�2��S6��<a�졻���͈?Dcmr��i�t�F;'j�5P�z0���xr���qXz��ϼ��M�k�k�<p:��t��*�fC��uΒ�]|h"d�����
mg=�ΫZ��K8��}�z|Oc���LeO}vkS�|F~���o���ft͖�W�t!z�����7*�;Y.�w��}W�sZz�}1,]����0���?kö����ʆ!ָ׀�?| �W�Edc`*�Ԣ���X0�U,b��
��N�}��ϼ�5�.lj����|��
�y�Z���^ͽ�G���{��a}��	�F���^>�mW��{{F����t�J��J�������wg���;��+   �  6�   ]��Y'�k��U�n��-��!���m�d��
/�r��6����$2pHX��k��w�jq���)褏v��Ni�Zٚ(8zt064�T��s�x[���a
{��M���/�xx=�rMƴs�!ȳ��I�JZ� ���:��_�|"=ҳ�W�}���;�̎GZ6rݨGd��p0���Y,tU��=`gY���W�`��jP�(!C��tgL�_!�ӳmJ��4�2��f�}uwWs�p��#xGC���[ޤ8�rm�>N&��<,h=�P�i�c���m�5��u׶�j�K���|/���'��A�2,�=��N������&c�G���vr꥞&#�7��]��Eo*��l���^b��*j͓kz��$�k$3�6�mv'<�7ڕ�w	&B��/�t��rZ���?{)���a0Ιt�P|����׺�e/z�44oc����Zn)hs|��Ȧ5� e�\EM�*��)6D���K`��<��9�ާ�r�E��Cb�}��Of6��6�q�Qu�3ن��t�r�JY,B%�+cS7��R��I�^�;b�h
ķ�T\��(]{�d5cݬrz�3k.����a�n(^m昢[��м�3�ə�}7����r�Q�i Q;3UZ����&RE�^�LtV��*��iB%����[�1�N3�P�o_Z�^�f�j	<�d\I$N��������~��ՑwZ�z��6�$G�6���8�&sbY�rr��8��.N���]���S����dþvm�������[�z���1�D| ��GнD/q����6���4��u2Ȩ�X "';F�!H	��׌ݯ�u�8x��)�#1$i�a�TH�9t�{�UYG�����*�Y�Yb2$���=�����<�3ׇ��~�QAk!#�@{�.���[N��'����5�l�kԻ�m];ή4C;-��O�8�"��H�"�D��Ub�]�x:'�Ϋ����m������$�� ��H�
(��c$�y�}�=�U~2/`J��}�j�Q����'o�4��6#�z���L͐4ObC�>y�q�x�{YO]��3�s��W"�C]m��K��f�IF�jH�R)D6�Ib���[���94\�+x����71U	)P�N���|�Vt�n~�_q����=o�+�{2pEE_�.�/Ȝ����M{Sz���vr���_oU`�a�pxB5�[viѽ�3UgYL�Y�	#��5����X�C3��c�͐���=���I���*��W�H�����z2��˽��������y������9���XCҺ�c5 eEq�E�r����\�0=j �a>�h�>8���x�u3(��E*�؇���}���0��\xU[���6}�<�$�!�'�JjD�C�nv,/N>�CЈ`���/ͮ�N?i�~���˳��!�4gXR�,�J�s͞����T옌q�ۀ�	e����ɒ6ܚa��m���Y��Op$X�I!�+�ȵ�b�w�ֵdZ��x+������,���
��7�h � �UB�{����_J��)�5pҪ���n�7�aI�*�"Eu{�[�|��ۓ�
W�v��I��`q�ٖxcs4X�k{�*�m2Og�y�4>W�/}�e�f����34����t�-��?M>�������n����v���xK(X Y��>=�V�^L���9��_��hmvV3�V�wvy�ٷ������2i��~�g����)��G����| ��"�ńP��b"�l�fH�9s��1�F.Σ��Z��5��A���ދ�<Y�w!��:!z�g3|����5~�V�Qu*��M�YUOUx�@������k=o�7k�u�}qy���@ w P P ��m�W�u��އ�D1,)�.�}Q�W���|�e���~��w>�� >�|	�}2����Q8����=*�	�9���uƝ�5�w&�l�����p����������WN۽\���]<��S!��l{3O3������fk[i�%���Њ�9�o��쐵Jd��g��FP#C@@�j��7�Y��6,�ꆀf��֪L��&HY��*8z�z﷫y��2P��+�i�;%d@�W&�A��������<v�5���z�[#L܂��#��!(n�ng%n��0/�ejt��X3J����?�">��H�ݥ��͇��:�rH��"JH�g/5��W7j�p�۷ ���6������59�ޔ3M�vM9��;�f�sz�H�9LH��f��]���e�়��~�U�}T *� ����B���:k�9���/D3�нh�\EGJ�$����x�͍ W��� ���h�x=n�tМyU�0���;��3˛�s�c���A�$��;9�_R�T����T�̌-�br��m'c6f��ޙC0��c���6@J&�jFhXXjY�Uf-Y(Es�7.˳�z��7+�,{�z�=<2�N���N`B9g����1�q��jЦ��]^`���{��^�*�����p=@ဣ!|Ζxj��j\�wkn�֒�����Q��I �I& ��/���/W?3�+5������
zoP�ߪ���憉��ǘ8*���V�g.��{��#X�Pܨ�f�D�? �=�n���ϫ�.�������U���>',�QD"�AUAU2,b	qߝ�y�{v��c����',]�3g�͜/j��.a��<ˁ�1d�B1H�J(0TT���D�@'ࣶw��緼���Q�<��F���ŝ�+cz����6�ݶ-7�wXԸ�.��<h�Vge�(k�w��w�Jt��G#.Jn���{������6�f����ܞ	)e1X2�S�+M�l9�J�p�b�˛i���#�d�K0{e�Æ��̼��}��o��4�����Fn�o��}���;<��Hƈ�q�h�G�YQ�$��#m�i�xKj���~+�B�/:6�գ���y�:)?\ݳ��inW_9��oM�[�:�%�0�[��=wՌ&�����=e����3�˥ّE\�Kb�aπ��'[kװoY�x ݋:��H�Z��o��7����w<4fL�ӕ�G�J`�7�QW�A�Yb���6���X���\��Ρ�Q�_�7ҙv�o�۽W��S�0�m�:=|�u�~!JuP,�}eY߾�*"�Db��
DX	���1X�J,�5�VJ���E"�VT��H��8����L�aK�^n�6�QLPΠ�iQ�5�D�e�<l�[���iE-l��W���el�����ϰ��.�M�7e��c�:��.r��O)Q�*
��^z��;L�.��<�|x��I�۽y��%�h@�e� �[m��6Io�L� �H?�$.>	�z�Y,�`��l�#�C���^.�n��ɱ��++��=��TT<��R/D��Y��Z�i��| 
�vc��:�:�Mq0�D�Lq��nL���J�)|�O7=;nah��#HS5�40>�^�ق·7�:Xµ~ի}��i����x�9���G=��$�n�'� ��Z��v.�[!�S����:�V��v�&�����}�>�N������Ww�d��d�ǝŋ7����I��B������s����2e��[ɍA豃��2^jᲴ˽�������{~c�rO��&���=�����V�ɅknT�m�����Խ�����ܼ��6���5wR�m}&>`ܕ��LXc\�)���.�k��O5�c��Vaɬі�c`�O7�����&�ɛ���]�2M��3Ff\��\kML�Tl�m�F���ѡ��	޷F�6�;\�_ak>X�ı�p�
 ϱ�7�+b �`��;#�Y'v׃�i �2j�޻6�Vd���^�Љ��x2������9��],f+A4Z{�L���iޛu짮p�~ e�E�p��Ć86?���ɅH@������[���΀�7�T��ݍ�}0�S�)�۫���=q�LY�����5�� ,�y4�,�]���0f��gg��2���y<�_)
�Y�E���F���a�e�b�QE�-rkkv�vŊ�@9�zo=���<��"���@K��p���Sڷw0�ъ��e��ҩ�Վ��)P���[#gzs7Z[J[X���ǵ�vA��ꓳ��.�m�r�t,�~'��
���&]_u�i��\�I�r�ҕz���b}�0�w��i�:p�7��G5M{g�(�.<#f���P��uav� Ӌ�Z��m8�m8�}�z��ⵋ���-7,���k
�6�k�钑�k0ً&)Y=�)m�Pr�u�;ϒŦ��7�T\�����_�')��O(<��c���G��ϳ0�C���V����$
�zۙR�ž��X�WF��Xz��X�Ÿ+b�x��~�ࠗ�x{�e�~A^"�ű�X-C)�Uh6��n���)�zz�Z�C-���ѱ:-S�pi-�ؕ�����+���{�?=�������͋��a}kP�T���@m쾺
7�V�s�V@��1����:�i�] ڮ�=Y��.��*�j�	�;qG�V��b�P˸k'�U����l
�k�@ p����t ՞�m��0v��P� �.�yUꪧ��"�]�K{7om�:�=Yݙ��w�N�*�����i�������]�jW����n!��^�Ϋ���9��]�T��م���v@+)��w�W��@�7�v�w7o�  �  ��@  p*��    �[` p
��  �   ڨ[*��� �*�       P          s� m�^�w�����W�I��q�9�'Q�4LF�n_]�=O2��O�᥉ݹ�:���Z�r�ӄ�k��e�z���iÂ��m:���ے7-�a���y�5�wl  8C �ب    �*�Kj�Fו�J#�D�I �%E�M��F�@����޵v�*ձx]͉{6*nX�{�$9Vac�F�|1���U�'����.�,Fp���}Օ^Й&�1k)m�Z�~�FK�I�}��y��P����;L�	<�������=XuZk�Ma��czd��K)q���z(sV�p���#-�*��S.��n�V CV�)΂C�!ٳ���6�e5<��J��}�g���3��3��	|ׁ	�2C��|���]k�����V���+.��-��[hQ��WK�;��p4v:K��)<w�-l��Q�|�S�|*���/*h�x"���"ɡL��	-�e�,w�S6UUH�I�yoo�[.�Um�����\���S�����xl�(^.��li5?}�G϶u�Sk���
0�m ������V@�����l���Q�a`�0���ZXʔIY�YJ�#aE�*U`�H��EQ��
�HO�ߥ3���ɡ�����Q���A��@�S6S��8&���Zy��Z��3fYR'�Ol2e���&�kt��`U�UB�	!��3:w��M�mƘ7��T�o,s��Į�>��+gp�
r�M�k�-�ϛ= FoK�W��hd��;�ν1�=���9x�PzV]��u�;����5�7Q#�����[|_+�OٖN7�7wC"���4�Nm��C����~gE�'�R���b�!R��%9�V�38XAt!N4���|R6}5��zz|  P;��j%ͤ��j6Y!�	E�$���I�~x�!gRܗ�w���w�G�(��sڰmL�� �u�շ=����5��8�K+��۔��P���&A�y�.]Tcz�'h���,4��p�ί*Z�{�ΦI6���\����=��n�8 UT��B-)�h۰��Y�9%�P�D5=����4��8{c�sp�AW�*c7	/灼���us����%��j}����� �)Z����?,Mv��:R⪕�:,��񦡓[�6�qN��o�[����jcb�0h��L'u�&�+��=3�<�cND�UV;=%[���mZf"!���7u}��)zc��δ�ƑB�b�s΍bIm��_}��C��w���m�ۮ��n뾯Y}XZ�
�05$g8�T|�;"�:r'Ͳ2��l��_u��0��ͮM��s��Xiن����9�&�t��v�}���H�i�ti�� P��R�zBf
@�
y�.Wl�sݼ���'�1��U��3��LL����U�¤2�����0*��\c��Z������ڴ��h�M�)����v��;\�̞8%wmHAab�	^�X�:כo��<S��H���
�Nw�\�5�}ΕX��nK�:�r͊)�-i=�X����	�a�:J��쎶��+��o�|x��'e�m�S���t	�"Z�}�,��y�M��?8�{wu�����e*8���sR�9�[�B��/�E��-���uV�&�Q9��� �m�d���0&��ǣ9#gy<��s�b�X:mA������e����"���]���Y���drVCʑ��J,S�|�O|K�b.Rs����:��CP�^#���L�"����$�/�w~��ߟ{�e�|�4�d����ҫX�N�3�K�(��G8���>a'ϝF�VL�bbx���]?nĥ�t��i��G_ܦ�篛�#:�P:4��R쬷8�a��#������+���m|��(�$�;�"���s����Tꔇָ�$�$ݹ����KνMbV��P��fb��c�f�j
.=����5���~�]�$76���U��Ư�Y�ىNW��L��EY׶F������������R�w���m�V�y�eW��{��;��׶���Gp� �P*��  m��m�l���?w_���+Dn�U��{�Gg�ܖ��y[��~��8[W������h�����[��,i� >Ǘw��GYz:�H�������#�ⶱ�}D��ؾ>t��t�c4��ܠΛl������D�[�Bo��i���`V&��S�Ah(�iOkx�^5������R*��|�x�>N�Ea8B0��/n?/r�W����n��P��QR�;Zx� 5!�c�8D�!g*�n��K4��<-��c���:O����Y��mc��1���� e��-�����-��x|.�X�o;_bz�i�S�k8��\c(X�JbL��rw.P�;p{zow{q�lm�SqD��ĉ9#L�$m����'xn�:��St�_ɹ�Cf��
eu[]�I۾'���T��=��0�J�qH�9r���9��U���(�,��QT�U�Ϲ���~wyxR�i�o0B�ӵ�P�x0���vn����Û�r�`'���E9!�1.�1eC��-#��1����;��Ӷ���[��|�J��·��2p\j�gY��bXP(HCK�v�ɡ���X��Uu�I��a�+u��}2$Y%���jjj�YVk�%�ܡ�'n�Έ�ҕ��އT#�9���k�"���}�Bv�6�s�Be8�6���xg6��K�i�G��\�����Y֧��d@�F���X1q�Nv���TZ��h�,����|q5(��^n��Tv�mޑU�*��s���js#ĝ�m��Jh���0��#��1��=j�P3kZ�窙��0���x��K��*h�Gg̾����CR������e뗏׉n��mU���h�a�i��3<B۽x�W萌\=U;kL��a��T�Ҁ��d�����$�H$�o�'r�fڍ��J܇��9%	Һ��zf�X�.-
`���ꎞ@8m;�r����ݍ.���2�<9L��c�U�vX=�ؿu8@n������K���3��l-����	�5����yF������{A���6ȣc��
����.���V孔�W�M��2iմ��;��
�a��@C������4�����U�������-�Fm�]ݷ$Sб�0���R�s��?=FIp�����k�e�s�nM��$P��,�C�����f�Ӽߺ�%����ZU[lYd���B�o��^�+
9�yFW �����^�4pHWr�=�5�{��ř�N�5BF<|�O��!�d�;J���GM���WwU�Ig��g��k�LpƝ�KV7F���b�k'�}_T4$ϕ��k�xd�k��8�G��xƵ��zD��< E>RQ DX"#��Q@@�
�x+]�e�戎멶=���1T�u��<��e��S+�f�c��L.�>d����-
��#��b0�����d��0��Ҵ����0Էlu�Y˹GO,�x|���_`^�}�Rh&I�F���K	��@6�I��X��}ӗ�금׃��+ıu������'h=�Q������/�f�߇�,�1�Xwm����<<4p^�����$�$@<D$�댤V���Q�y���J�]�6S���TM��x��B���nwK�}!9��=\�k[��:sI.`��S"�֟�2Og�v�UT�m	��i.y�սO���z�8Fj���T�tGFj��כ����ʞ���Y�U �۩X@�#���`�n�9��W�٫���J�
ï�I�pE�E����]�АA�(�PȌAAQ�b��6�ʌ��,��ؕ*(��b
�E�V�5`G�Y=\|&� �.1�N�y�r�V~�W�_�-��Ͻ��{7���mw��}�w~W�< ��Om�z��h@�Oa�mT�
�g^�T��n�'�i�T��R�P  �T 
�   ��_��������~����{���]��Wp����7��7���X�� �es�K.��5eQ���_��*���gWvU��Q����b�d�i��T�'>VHL�s�O��oVq�<t����h����+�L��R�5������N�nJ{���	���B���x�r�$��,�:���k��N�R��3���@�j����5qg��̾�lm���ۃw-�`�y��6.���wzP#�$i�k�[oGdγ��~�̦��Q�3,�T4�[vy���k���oޙ�Ì����eBm[G��S�-����)a}C��<����~�q#$�qݳ�UmĪw
�w��]��6�FX�3a���o�gq8i2�����JS�N��3��� �C���}j7�h�'�y[����~���vU��f��:�$�uk|�R
C@j��U��v~f����C�Y�Y�B���ԓ�ƹ;���i�O�s)�\�70�1�F_v�MY�v$P����#q�ͧ������9�]�#�Ax�7sX�8��oZ޸�&�:�]�zq��ϵ���P�0Vh���uЛ���m�.CD���΄�e����i�ˤ�˝�3?b%���o>u�<$"kU�x��e��|-<鳧�t[�#��/+ݻ��^l���^��&����G	�О�(j/��u�\���Ѥ��q�k��n�N�^G�>y7�3��k�γW��zs
м�6I�P������w�ݼ',Յ�8{؟e`8E���#;]�bG�g(-鏳�~�s����-��F3���$+:YӠ��}�\S��f>���5o�� �|�b���b[1�6�=�:��ci�}���F�"�=a�}J#��Tˁ��b[�5��y�.�7PKJ�EyB�&54[�AeJ�CY�tc4�1M��� �5Ī��"�b�L	��EX���Z��N�iea_���H�+m�r����TvYA܃��|��%��Q[���v����7��X�^@� e��щbR<��3�v?��8QG�-�12�Ǒ<5�e/K1����TVe��҂�w�7��S��L����N�c��>9��Aɿ:��M��1[��_:�+�o��a�p�M�{��4��۲�|t]��g�(2�h���6��>�(�)2�>�#���ĤP�Hb�b`�l��(�y�f�����Y�cu�7n�i����y��C�F2�9[��y-�5���1U�̨�i��k"f#*��E�UWE�cr�k��j�ul��X���aƘ g�������s�������2��D��]����tӪ��6�'8B1^mE�7��Ϸx����*����W}�i�3��/ ���+M{#��=�,�,�]�.{
����&�Z�2��$�1S�{�,���5r
��q<�6Έ��w�K��¦uH��C԰maΤ$��eHi�.���i��������ŜN����Sj��=56�����c��t�GwY���£���k�[na�i˶�^�E���8��Y���5N�v�ShT� ��k�r�x9�{����
�'k�zy�٫����Y�v�&�5�[�e_��d�g���HV�<~KV��Y�Yw)=�株t�҃�m������l�)�U�ɝ�S��[���`5�.�*Iejbȴ�rީ���Z�i(-I\tAm\���2�m)�ZB$�W�[�+2B�i�ו�~�H{�\͞���:�¬vۖ�X�'ڻ%a��X��g�)�]����IK�TYoR�^ɻ#w�� �, \*�ŏ �½u��`b9�Sxqyn�m쎱�"/K�H-=�&Qh�`�͎����{�����x}ˬ��p�d��`�A��!Yu�1�g>��k~��'��rا��vF��r�v�����o�Y��U\�a�q�.﫹ޑU�*������'�Ϳ�럍��|��n~�SsY�Oa�8s˷'>����xb!���}�ܯ�`f�Sq�q�/�r��F��>ر{.��I�o*£�i`}f����B���K�(��ԅyK[�rM�L�4	��+�� �7[P�,o�g��V����uk�"�����L��oɝ:���,�x8)5% o�'��1<9 ��6K(-saۺ�TX�N�U�}� (
�w�y��w'%}vJ[q��ʛ��V�,�����;�Ju��z�c��;�s�^D�}U�G;�dYM��#Y��ük�[��|���wO_���YCO���<E�l�<۩A�(�[�^��w��ۦ�p�Y�8�Q2I#m�ی��2�Ϲ#X�+��b�˭��^a�GA>��zd��X+�ح�7d�uM�#��'�'qF�<O�þ��	������ٲb_6gk8&�d&`F���zy�y����b��[��V��`TЁh`xXsS�����`q�$A��m5K�ѹ�0�}mU;�5Y
�3M1�:dљ"s �%��+�̷��c�T��\���U��Ƒ����	z�ۋz���V԰> +W��;����3j�>�
�1�5&;/Mфʭ�z[���V�2}$QO1�}���Ko�:����ߟ����$���(#6�v�#���˻�����܊�Qmw8�e���i[�X�6Y��?;_���c ����z����C��GR�m�*V�P�^�.'p��[9�\ҹ�뺠� Ͱ   *�I$�Bdu����}M����L$8�)����I>S�4����t���\��>��"��]��?[��>��&3�cZ]�U(��0�\r�q���:DtW��*X����C�s�-�4�N�'7eɤP��3ft��B(UT�j�Ya����ݭi�#�}�e�I�'��=�a� �6�c������np�[?+ �$u9�o�fDo3s�_�h�}��}��i�'�  �\o�W�w Ӊ{���s}��c��2����1';X��a��f������kq�=���../��+������<��f`+TNL<1�	�^��c'�
w��j��V~�I�m���]ª���Dv\J��$^A!,��7�0g&]t�� 2�)����QTFH}�����xy߼�}���㨶E��dD��,��x',�2�2�0��ي���YX.n&�:�4!g������ي��/�<���[��l����Sk�;��q�S�yG;���,���.�b����0Wa^������9�w	�&�09��� [0sr�����ܑ�;ĭI�|��ۓo��4��ݛ��}�|ptW�݁�d��F�L�
�X���wHN�1�a���⇡
��ǅ��<M*tjCs\��2���s��LL��Xl��Lʓo�8TWB,�l��;gm���W��/��Ōf��z�D���u*�w�b��\j����A)#m��n��T�<}�-�����Kڃ����JtpL��V��s��O�><}]�/��Z��5w�q����7��s�.�VgWf�r�2��sP�28�`aR0�s �A��SX��4�?��Bh� ܓ�k��c�X�#ʿ<-����Œ((
 ��aG�p'��y����O�K�����Jy6��t�Z�ڕ��qB�݌��AwS�>�'�%,0��Gn�X3�5��1F�s27�w���bDѷs���̇���EgX8�{g9�����tDe���9yd�:����!��@^0`���x�-�7�� 6H��LT�?s�
஝&S����^�����JI�H�a2�d�$m�d��>PHDl��w�F����� �A��޽������)��+T�,�7VA�b��
����i�@�`iv�\�R�׃�5��F��.�<tXr��Q� ���]�w�Lm��7��l����:�a�B;m�Q}y��Q�ӮF/���`�����8�����1��fňcv���UP����{�7ZS#qC��#�<�+-Փ�X���>鉛�;|�^Q�[��rNŹw{v��&�{$��ns��/z�A�<#F���'j�}s���nguAi�
�`�dX�<bCG۳��њEr����Ij��R��2��Q�����u�����a)mk���{��Wp�W�|��m���*����Ƹ�i���q�;�f��u���z�
�U�F�8��B�L����>�Q5�6�g^Z\��>���F1���/�U��[=�@�m>���X� |�T��F�6�!g.�,[[���N� �a�O�z�Zִ0懾�C����	F���FE���4��g���v4.烳�-��]gc�!<�ܱ�Ƭr�^[#���N��H�To��j��3;�L��b9Y���c�n ��C[۷}�Nev.�lO;h����c�E݊,�	�ª�,��m��R��4wz��j�������qzE�Q�i&���Su�5�cǅ��tx������F��Ƚó*z���ӏ�2��k��Z��ĝl���k��9�  ��@
�    w	�=�7�K$�P����^H��I$��5�	�F.Q�A{�nN9k����#(�o�].��7�[��p"�Je�����jYe�GxB[1���V��>X℁��8$pJ�;-Ib(6n��S	[F�_�DG��7�{�mpتЭ���)��6 b&@�&�F�O%�����i��.l�D��\}����B��PnXXl�.�p#�D��D�y�7�V}�!�?Hy���Mz���K~8��>)=ܾ�Y�g1����^}������'9*��c���7ם׽I��[?m�C�-3vk�[޶0T��'C6B��gs~X�m��IL$"Jc�6�2Fۚ_��L��R�q�+|�=w^�w�ݘ��V0m�b�jN��=��y&|d���aӼ���d����{nw����i�r0X��Q �U1"�)�(�H������s��|��>ْ�d�y�>�v���~	m��K��mp]>��:��a�Cܦ-v������Y����8��s�4LHi��s�6��K�5.M̍,vI�2D�aǅ��z(s3f(!��|�$���(�yK�!S�Ja��|w:X/E�Z�JdV���3:�����������!�-�[�'�R�ͽOG�|���� 2�oww�TZ�4My�Jc4ܐ���\W?=�m]&x$ާ����'��,*R�,XL������>�c{�����oxeLI�d���p$��㑶ɒ6�(��$�5��;v�fM�L�}�ƜkW2em�凭z��%ۍ�Օ�{&A�1bW�\���ET$���ץp}�,�m���vd�ϙIX�,��9m���`�Hx!�qK���1��i�����Dɪ27pJ�Z�������VaT߷,����4�>����;�/�n:|�w�Q�d��Q�{���2�P��(ˬ����f�ua!����K!�e���T�R�59�S���cI�s�+��ǧ~ |���jl�a騰�ڢ�Ӱc`��&]�1����u�v��[w|<�i�3F�>��Y��e`ذ�J�[�.����$�X{FT�sb42n,�5E���{ם�V�Qm��m�"�Z��$��#n|IbF�[���֠�-�gk���^x^�ȑ������ﾮ�D{�l�|,5Yh��(lA�;OMQ"�$�ɋg�[���iÓq�@	�	�g��?����,z'�ڛ���k�.t�&�GX<n�U�=�����y��{s���2�'���fz���f�ޗ�S�ӝ�d�����	�*H׆��k�J�򷡭��t�;�CE�/�(��C�����9�DX�����')$�`�d
��,�V���"���H�T����X�" �%��Z������7q\���(�ݜJ����I�Z�61�X[��+GVWf4RзX����C`6���`@�731�L���	=3ɨZ9��i��}�� �,��䮴v����/g�I)n6�1�[ۑ$$�����Q�KX������\]�P����Vk��]�4�g9a�(K�\��ǌh$ѳ֥#�P��[>\��9Ɏ=-�����{�7M_eX��� �l�a�6*x�j���>�[�����F��_+<F�r�z�HҬG�u�iC����O�V�xG���z~��
ӱ2�D6u
�I����,�?Nz�׎�;Sa>
�ZF����8)�;�?c��>�ַ���3P,X���m��\}�أe޹�v�F�/����ߚ^�$1	����(#,\��杫��� I �� ���H@��?��͒I$'���!($bH@ 6�$	���B�/����!��Ik��߰$� ���	 @�H �?���'�����I ��������\?���!BBHI �H�@�@I!$��d!H��~�`$� ������ ?�}������@��7�`I �$ _��� ��5�$� ��0����6hԒBB`H@�?�@� ?d���	 @��$� �������?��́$ a���o����	 @�-`I ������)��{����8(���sn�_��0�� �7f�� 4�PM$4 � H             >    �UT	TUP�J
�U*��$�RT(                      �    4�%�w/aXt{��=<�������1��mtz�G����{u�V�;�O�����}���R7��l>�p�@(���{�<��gf�}��}�w��.ٯ.��z����+���o[�<������+p觾܏OVw&��}�ukt5���n����� ||    �}�7���λ����o��m8�S{s��#�;k��U���'���n�i��tz����K�����w�A���y�t���o{�q��{�w���� u��� U*�i�}�oU�ݷؽ=����N����z�z'�]o�{o��}�;mzu����ײ���rWZ�N�޽�^>�����U����۽�w��{o�{��]�<P     �v.���y��N^�|�;���z�{m��w���SS���^��Wm��;5���ֹ�u�n��i���mj��֎��t�mw�H��@� �P�+�}ݥ���t/n���iǀg׽�J�w#}��﷽�=eۼ�x�7���T+���}��}���q�`|ﻹ�������N��]��`ݎ�     4�]�c�#v����9��o��Y��z�ۻׂ�٤��Pk}�{��x�s��v���t���)�=k�f�������t��Ws���>��x < >�PT�����ӮO��(3��=�{8������{���-}ju{ooN�n����2h��[�m��x>��k�ɗygݽ�}��m�w[=�Wjo��à �   w��{�����yO���f�|���ꔫ��{���V��[�;���3�\��ןJ�����K��n�٩N��=u�-{�����=�})B^�>�yB����x� Q

�xO_Wm+Zg*=��7�;�'F;;�8��=����z��^���F��.'x�����!����s=�>����/wv�ەΛ�  ��	��* 4  �  EO���U%  �    "��	��@h 2h��Om��P"T ɠ �� ��
�P@h    �D��=4)���������h���?O��	�?��쟺�{�}��=�_�����q��� ���������$ �X{$H%! ~�@! �����y!�� ! �z�� $ ��d+ BB ~���$�$'��� ��BH@̀B���!?��HT��
�  �� ��d$́$��d�!�I r@�HI�I����%fd�%B��B��I	́!2f@!* r �$%@�P��$	P � �IPB�$	
��%aP�$�3$��2 ���$�@�$	�HL���*I P 3d s́��9��(�$P r	 T !P���+ �09�
I"�d��d ,��  J��� +X �$� �I�C I+$*@����HVI+B��Nd�d ̐	%`K����7����o���b׬~'��9�Tj�W����+Y:pVT�Co��P��}�![&;Gs��/NnV�&a�"�~��O^���氕	 ?O/�>�}�����,-eK�WN���,����|D*��2a3��^*�~%`�g˙I~ݑ$/h��y���5� '(-������y`x��!�C�AI�����q*����9��ZÒ�si��fJ�X��~�;����d��}:�� �I��bnZ��[�K�1�f/�B�2C�C�C2�{_7|��ͳ��7;�[46��ȵoe�P��ށ6��vf�.�b뉊3X�J~���	� �B�9�0٦�DXv��&.�.�6���ׇ���^�Y;'�_Wo#?+ k4cl:��kk7�ڲ��L]+�C{����:��%�������74�.���ٷ�������3��QE�N�I+fq�����x�t����oVt�P�m#�]��2m��7d�d�{1?œ��fPw���S{6QB�$�����T�58�l�X;7��S�t����-Kթ
F�m�u¿W�(�D��u˚º:*��p��7$p.��(`G�ᦪ��X(f�:�2�\4���K��W�t�e(-0�ǓY[����z w�%n�;��+-M[ӁGb�k�Kf�ɚ%I��P�o��g��`�;!SVwf�	�6S6�ԬX�P���0,��SZk�N�(���u��y��}�����F�:��ǹ&�6ŵf��K�k�Uo��F�.Z�n^m���N�Q ������(��u�i� �h�3�:�8��h;t�X,of,�����Ճ�cJ��{��6��G��%_i���B�/�*�w��G����$�>$=� ��$>2��=�ZOI�C�C�AH}H}d*C2�R�R!�!�!�����'z���N�7���M��m�լ�2��]�w{b�R��NX[�ޝ��̾�q�د)6������,�EWi�fdPeM)��Z^���q�N��֕G���&n�u[�K�d�iY�Y,nTY���ӱ���#0���G��H�>WbC;P��-MyV*٤��s?7�ꚗ-��&�Z�I�.KMfˣ�Y;aڷ֫qɏ�G�e�#Ȯ�Xh1�+7�Y�e�k�ré�]��\5� Ω{�T�%�E�׌�:lռ�ysRX���4e��Fܭ��j�9ݣ!邹�d{q��^�9`��W��mbz�&4�� *^���lk���B��v�_də�"��D�4��wI\�����9���cm���&�eB��(�E��e�Oͽ��uLt�B�̊�����{<YS����;MU���L�77�ԭʼV\��/��r�hX��Ӓ~q�����i֬G5���}��WV����̖�L�%�pИ�Hx{g
���+��9��޼�\���ë��NU��w\f��p��5|#���ۏ�%�NL�l��ʝx�z�3���t� ǺkB�X3o�]$�*Ċ����/+��c:�Ge�n�P��ً(��]�(��xfV)�W����0�5�}�^�CX�ӳ���)��Y
�U���f��>� v�3op�Z��-5�����Ւ�ͽn�N{SMv_=���h��=}���z�Em����ǟh
B��W�"���qtb4t��,f�Y)�����`�)仩Y��q�X�*떻�;�_8���7�^�o>o��/Ă���d2CĆH|H,�}}�˯��}�p�sS�&�I��_$w���l��v%Yn�����6��c)1.�WgE���"�,�[b�6	R�V�r��Ox��P�5vג�(G�c�c^�f�@&K	����0T,n1�X�)UYv�����ܭݫ��ݧZ��{��h5�*����1[�4(��-��\��LF�F�=g4б\�ٰlPb�Dp3r]fK�a�3T*#A�3��6���nj&�����7iL�3n�Nv{{B�el���wW�$�-Jܚ��2���web���;5MD���S%��n�7�x즄���fd2��+{���]e�2Zq��k�4��XNڵ{1�r��ۥH�
"�n���H�֠�F��d|�;Q���9�hI��o�IZ)u�oE�[��W�%�f�F��[e��b�r�3E^V�h�kd#K��'A�U6FG�,��j^�b8�i
n���y��a��W{�����L(^L	���z3Z[�n^�^6��Dua�!�'F&P{{�jԻ�� ��U��E� ş��ca�(,o-���f�E��Ѕm]qU�V�`���*nJF��IK�a^>��5�<�j�r��5TA�upc������L+M`��de��?Eu�Q�ܨH�q/�L��Ij�w���m	��]��=���x����x�(�.��U�W]�Vʫ�%*u��2�ہ�9W(=6��^�$N��F�R]1$�aZN�t�h�z�6��9�j�ڶBnagFa2uO�X}N@�������
��l���C�B���!�!RR�R�R!S�(|H|Hx$����4U�J����QAeZ T$��7���@���7�Q��Z&��
���>$��O�RR�R$>$>'�I
������!P�����מ������z�����H,!� ���S�����$��R!R
���B����8�d
�R
C'��� �2AHT�HrB�>"��v��V#A��^�σT<H)*HzH{HrB�>�>$<H{Hd�� ��
��=$>$9�Զ}��������!�
�R
C�d�R
A~�T=,j�L�(��3*J�R
AH(V �@��B��*AjH6�� �� ���
AH) ���6���]As�TP�¤fJʒ�RT��R
AaP�i��b�OL�d��Hd��R
AH)>�U=�qX��0��RT�$��g0��x�����ciz����ԅEa�
����!��*VOi̙����Id�R��T�KJ,����0��W��*��ښ)nLZEd`�'�i�Xs�K �=�L��>��R{OH!�iXd�$2C�C�B�=���=$<}�d��� R�I���H)U'2����YP����!�!�/��2�O��	�4W�K-*OL���{H}a��da�L �=$=�<I�'�􉓜䝨�g WƠ�Ҋ��
>Bf@�!�!�B�>!釤�ć��O2AHx��iiHzC��Z��w������Hd���H,!�鞘�����4=�P+%Ǥ���������HrAHd��������!P�!�!�!�!�q�'ć����rC�I�'�����糽ϑ����>$<H)!R���¡�+I��-`����,U�|C"���{��㪾�Y=$*C���s'�I�Ͷ�� �92��䂐ə���C����������!��zHV���Ù`�!�<����,���=Z�|�Rx����/�J��Z��m�<��߯qOam!�!�OhT����
��!�z(�9'�����R
C�C��M�H,!�4��@�X
E�!�1�du��ӑJ�zjE�ʂ#������K��JG�y}�y'��$<r���Y�AE��C!�����۷��o{�c��E+#Nn��2�zO:q��c�,S�J2�\�>�W�m��u�DC��F�M,Ա��a�m1�
AH).�]eA-;VlQJ�Y�ɒ
Bە��³&��aR
AH,*
¤YP�X-H)&F�*T*:�u�m��渶ͷ����1D��*T�����6�0��{o�H) ���l*��R�Z�M�IYP�����2��R��+%�� ���R
AEH)&5΁RVT�g��R
AH)P/���
�eAjAH)ҐP
�`V
��m<J�kT
[EQ-
¢ȂZ�!m�@�bP�A�k����\l�3�Z�
т�`������ZR-H) ���DB��� �YE-�B�XT+
�RP*AaX�AE
ʐP+PچH) �5H,�.�
*��!�B�><��C�&Oi!S�*
C�C�L&�W�?t2����DYm��zCz�!�C֡���)>�}Z��|L�0�+F!R
C��9P�����F|Oh�y$Y"��Ϭ(��ԇ��+	� ��2����$=�>�.Cۆ"������J���>[֒����̟_5�
�G݆L���=�=2ac����E���t��X�>$�ć�1��B���3�5�߸�LQh����Hx�����x�=[$2��ߖT^i<�iX��!�!�<H|O����w�Q�$+��R��[����V�aP�o��ϭ��}HT��\=�2}Hd��"�I�!�	�~�6��y�"fTAX��+"�@�
V!ȴ��y�p"�\wF�_EO�ȧ!�+}O���F #�>R���ʨT*��`�P�=��II ���d�����,�[PD�X�Z��Ւ����*�ڂ���A�QB���6����°�m�B�U
��R
AH) ���Q@��35�Q����HrC�	�����$<@�׶���������篆�~Sߞ$E9!�!�!RR��9!�x�@�*+'�-����C�|H}@�����!�B�=�2B�>$*C����!����C���!�!�!�!�!�
C���OhR$���������$�Oh!�!�C����*����Hzai!铽vNF����(?�ɝ���M�a쑟F�h
�n�y���@m�""(�mef(d+0h�3�!n�e���_�e!���;���������+Lp0��p �`!  ' c �� &�` </��� S�  �     �N@     � 3�[!��v�8zU�p0��m�f�М�o[^^�ŷp  [}��� N �    ' c ���    �   l@     0 �          .�5O  ��0��x� �   ��m�n6� p         ��r���\-0��         
�               @ Tܫ�ɶWu��J�   �  lùT   x    < <
� �@xx�	��8@x�m�8@x  N �۹��W].��K�̵�i��K܅���f�U��]S�o#{���u�];��{���z��z��6�۬���z��;��6�qy�j��Z=�DxN9���tn�ܽDh�w��綶�WVnz���mvlz�]�g!��^r�Lc*Ӟݰ��Sn>���w+�^]u���핳9k��^սٜ�m;�9/Q귛�sݷy�p��m��z�k7����3ڮ�A�Zu�^1̯���5�޽���[��Ŷ��^�<�z�Ogo���j�R׶n�z>�[��ם�ҹܷgm7�o����;��]���m[y�:��ݽۻv�n����2��+ßc����v�������]N�#�s�]����D����s���8{TӷYu޻�t��uݧ*���ݱ{�׷��o6�ץ.�z�k��v�����1����;�]��4ݭ�s���ݽ�^2��˸���v]^^ܹu��u�W�ot��]Ys\nw����O;����x�Sv�.�+���^���w�T�nyݞ���e�;��m���{{1�y�����v���%N��i���r���j�ޞzݶ��ݻ�x��\�ϻr[��q�۝�Vv�V�]õ��ٮ�������gZCm�^�[Nn�M�婵�mԝ5����uʺ�ץ�Φ��jZ\�7u�wsu�c�'l�^���Y޺�i�x�O%�[睎G���6�u/=��ƶ٫��Z]�ӭ���;{7W{:��v��޾5�o&���ׯl]����v�n]�ݽշ�`�����]}S6���{���ջͳ^J6�MK���&�l;��/v��g�j�ϵoy���kݽYl��t��V��n;jZܷ����嫷z>���K��5'�e��;<�v;�}�ss�{�����Lw^z{��y�;�ɞu��>+g����v���ۂ�f�םƔ�=���Mӻ�{u��w�����]{����wc���T���6��-]�.�{כ{�����[�{g�:Z�l�p�{����Y�[^wbu����x��uqeꎺ�.-��������\��4��ۼ����W�z�u��q�����v�ܵ��w>��^s]v��{��;�5�����gR����v�{t���������K�m{w�=�Oge��wn��k�n��w����{�z�V�+���d���n��Ze����G^k�ۣk���ݥ��ܫ\w{zn��S�um��ku�7g���2rQ��)yئ�R歘i�ױ�S/
ui����G���^��v�/K˰�{)K��6^;m۸^om6;ݵ����lֳ�GZ^�S��^[��v'u׷uqV�����ٽ���l��fsy���(�mɮ6����u���{v�i�p�R�/rU���������Y���3ok�������qN*��E�^k��n�6�ܧr��]�F���y��s�5z�M^��u����<cG�a�^K+�vܽJ��jZ^���N�m���w��4�'ֳ�շ�M�]|��w�[oG;�=�ת/���%���jq���	������}����7��]�����R��u5�N��U*p�r�h����l�m{����f��皬�kz���z��ݽ��;ɞ;���m6�v����o��m�k������-��oe����yӹ�3��w��;����+�ٸ���]ŷ���h�a��wl�����z����EC[��r�{N�y����=ط�����63u󻵹�o=ɷ��ww���V뾮��Om*e���gwU9}��S{U��h��x�{v�����x��v�m�w&�����n1���L�������z�����/3��Y�f[�y]�����vg����s��z�Y�R�%+��.����sn�.���Ӟ��{w�����������^�ڜ<��od5�5�e�J;W�u޼׫�w�-w]������M9D��x���T��Q���y�G\��Wu�_N�����o�N�ok�gZ;�N��z��eݞ�R��]��qsh�ջv�8i��V��[���;;Dr�g�Wu[���;[�\�ۻ�t��r"�p��^:�[GX��u�λ�\ӻ��[/o;�m�kowwv�i빭osoK}v�.���sm��׷����]ݫ��x���z+��o{y�w��mv-1�a�y�gR���Zl[��n����n��k��k��?�����  U  @                  lR�iUϋ��֕8}���:������r�*���i��t]�֎�y�w{u����߷߿dS�eU����ݳ����s���W^�W=eu�g��u����*���틘   6�lVP�    ~�?U� �N�\��� ]� ��:��[v��o����    �*� *��P  
����_��m�ώ� P   ��   U�T*��   � � @nrJͳeP ���b�*T   *��U    *�� m� ��*��@  U  
� ?�/�� ��     �2   
�  U   �   62�fڪؕ �   �}���  p['�� ���l �   � ��  s���́s��
�eyY@���Z�36�@   T � �a�T @       PUU�{�Z�UUv@  
�*�  ��ͱ�*TU �T�+�*T<�;���]kd����@          U@W�u�V�*� *�ǭ���R� ]���[                *T��      �?     �� @           �TU UU U        T�   �0~                                                            �          ʟ2��ڶ��ov�C�v�.[ݽzwz�V����V��;�>�w�t{n��7�jT����T�vݥ�s��ݕ��
�6ܺʭ������[>�u{��`on��Gv*��Ve����)� zƽ���Y* ���*�{j<k�v�q�U;���k��{z�R��mv�dw��mUUe�����n��u����g���6�� �Wm�[�x�M���wax��=��lU���s%kq�ʦ�披�纭��ڧ7��+��sR���
�*����ݻ0           �~        � �{�                  �mS��                   
�  �     ��         
�	�6�&¨     
�    �` U T                 u� .eP�@ U �
�l�     W�M��*P            ��Cl  *R� �  ml�
�             � � *�    rV�ĩR��£mT��  J���P             @ *�� AUT *�T *U�l    �l�� wU@�  l�             �j��        �              {l
�U           
�    �                   *�         w lP  T*�             
�x-�����7��~�߀l��@      *� 
�p  -�     �P           `� 6   U  U ��+( YAR��P   ?��          � U      �l�   @  *�P ��,�^�۩[w6�ٶ�    �Ov�m�( T� 6�2w^븰lK^�$��[[ �B��m�p        �   =���UJ��Vڪ            �ݐl*����m [�  
�e įP � ��6�ހ 
�ս�  6¨  P 
ʳ-w��
�wQ�{j���P   ��*���;������|B ~�� ~��'�BHo�?����������_��@=�HI?w�~��+��*I#��~��DBh��I$�I  ��n�]�k�{U�m�l�^�m�6CՔJ���Y��Ѐ����m��6��Tea�qT� @ UU U  �ex�*
�Vn��m� �T {en�WU^�m�@  p��]@    �
�   @P*�            ��s��Z��ٽҭϯF�n^����2�ʯ;{z�y�W;.�늺�t���ۖdn�*� T �    �    .`U  [j� U    m��d�  ֠*�  
� ث��(    m�f�e[    n�    @       � �P  ةUP      ,ʨ
��� P P���s���
�U� ����  ;ܷ��p< *���9�#Y������?Ԑ�H���(I������~C�=ӽսW��8,��
ʹ��ȪR���T�-���  �q���wWuU�YV�A��� *�`�*�C�
�P�.j�m�R�<�QR�j��9���u�m�U�]�խ���j�� �(P@�9���d��n�w��>sa��)׋w"(��_ZYHQi��L�z��PI�z�b����kD���`��HHr�ۂ�q�����yԔ����$��vcC�x��2�z������\����S�{]�J���˧���(�I.�^w�;x>^w5�r�Ӧtm �\' �_76�[[#vfj������F��{�N��D�n�fvm `�`��s�ѳ�i$�e@<=y���-���,C�{F����Z���T��x���0[�*eED������ ��)�Y���l[���-��Nj��T�
�{leK���d��L��!�I��a��"�p1v��`4�M׽o����"�U��fޡ�83aLs��g9�閑qݧ���v���ՠ`���ݽ�3�՝��6��]s�ǻ�soU�w1���η=���ͽ�}���ؗ����/Nx��e���nwZ<�#��v����ǭ���ov�+���T�|�c�gfU��ə݂���e����WOx��B�Q-í�h����Y��zy��nx`�{�����^k��#���҄&�!���a��D(Ns�r�_׎��	B!@E L��I�B%��J�-��D7�C��K�v��yxxr�F؜n�/V�WEeP��kZ4�y�3eA��Zq�?	�K^����� ��|���y���T;����;s�{�=���%5ew�:��T�uh*�I"D KH�i2+Da���v/N��>���u�.���ٙ��.f� ���2���	4�#�l@eI��k�7C�(�*�G�{H���^�<�ͮ�se&Z�rA���)�Hu�}5{Ȑ2���X/r�����U�*���C����u|{�P�V�;�>gИ�'��~G���:�`���Ǉm0�I�:��Z_qu2J P�wp�:���tn���=7@�=��N9D��<*�Z�k8�b�wR%�'���$�$��%7��ޮ��[���;��Aכ�1f :fE�<�=FJ%z�]稝��"��ĒI�6�hwo�j�Vج��w)4�-��	��̩�{Ķ���Z��Z=��<�r��I=�N��c�4�O&U�CXR�� ��m� hf����(�If�+.�����m���;:��;�Le�i@�^׹m��s���D��e�<�ܹ����{z�R����G뙇l�&�nl+l�
�xS�_b`I$������6�;Ukj�vŜ�J��,6�$ I�=��Cw_��\�Q���� ������?Cs�Ě�����5���2_��X�@�݉+�����l�u�P$�Ԉe���wJ{1����|�@�宬�yً{�eI���&J'i��}B�eȀ�y�ki[`�W�f�c�Um�ڽz֘������?����>�5,�f�s��޽9�1P���xd��A����U6c��ǀ��m������{�g"�݄؜������v���� �s��@��{J��N�֒B�~��ӓ�Ġ }���G;��o���1S�����\5�R(�3Yx�0���yT��.<���T �a�M��h�M�T��I�o���l�'�N\� ��K�w�w�G��E[������kZ[D�]�t��N�L��{�H����lt�x'�z�7���x�m�O2�� K�B�an�(�����ka]�;!a��C����w |mPW���v��Vٮ����pP   �ow��o#ֻ�]�k�@U�U�TU���T��Sl *�aT]� w��F�Z6ۙ��/J���;��n p�U���jWt�d����|��[��prK���!�;�߶��k��� ^��\#�8��-��U�]�*���	�ĕįA��kT���Y01��k�ؽZ�L�\=��'��\�EkD�	�o����>J�� ��S�����O4�ݽJ#l<����Z`�{�_�(%$�"3hU���e8P���DC!��.d"��́��i���S��P��@y�ݔJ�'�y��&�x]���xM���X�ɺ�C��fȂq��Y�Ɲݘķ��78Q���nW���Ho��e�����Zӱ�.��mU+�,�JT�(�[i2ZI&����ᛝd�G%�4��b��%��4�;�C��$���O�m�Su��-�P��׫@�*�����"���x���i�ˬp��im*I$�	�m��{ߟ��lCom���Nܣv��Gn�[5������V^�ڴ����ov|��z����e��K����S6���{���v����u���鷰�@m��T0J�̐f3a�"R�~��}FX�:�U�Ƴ�)ivr�l��d�H)���\���#ծ�w}�M�`fib��
�.3\6,�1�rH��>��+���kı��m�;�]_�(5@�%DP �,�,��$R?A�a��C���<k'�17�95�#�4����ޞ����t��s��;�,@&�,lٽG�31�wy�St�(����� 9f��5��]�-�λ�uג̾l`ڇ�@�R$ѭH��k��6Pm���Se���u�d�Hb�vdS�i+�1�"��٘54���
>�u�^8�*�}+)pI:5��x=ʲ�'�2�9;ʯ#~�:�{��媷��Q�����f�y/�(p*ސ�H���n���!�'�E��nÓyrVa:l����%F,�Te;��ֶ:�&1�F��Y4�+!���Ì�Lg� [}��^ݭ���i�ߥ����T�$�T(Sj�"��Z@��0[m={�r
�w��'e��s�C9�8d:*��X��aٯkc-�I6M76ڏ57�;>����W�k�N9��s�������f�&{ AN��n�'����Z�&�m�k��ݺ�P� U*���,:B�綕�vs�_]�R�܁�[���ov��-o�ƛ�mFn�ԑ(�6��ו��<��~vA��1o��STo6u�ݝ�<�3��6]���zT3a�i"[I$h�q�繾Wg($Aa*ˇ7��מ+/ �� �&�f��U0�I?b\Y�6߿�r��h�O[K�l���;4�b����h�A�ݲ|��=�N�-tR:�aEFj��/(Fܕ�K��X�(�H�:V��A���e��x%cD��=;tx�>����_���xL��Ozy1^���H��zn���b�BI2Jm������M�b�X�F��E?��7x�W����+'��٪��������>YH�M�2�	��o�-тXУ�*�,�����r�%��8+�:�m�C! ��{,���_/t��ͼY��o����v����@>a���v�M�i$�By��ةV�;;]�f��������GwD����x���:�x�]}p������(�I��S�qH��L��)}��mnn`�y5pc��0�H�\��oބDs|�Io]w��P����ʱ;d�ӳ޸5��Ե�+m��=���m]�Ԫ�Pl��:��V�����*�   n��W^ܻ�<�7X6��
�� *����B�Tx
���@ x��K�s7alr�۔-����cv֥S�@m�w{u��m{���_�����I�e��Q���~��Ĝ��;y��#�/L�B �ම{$�H�J�,*W�ݍ�H��i�jfP�<"��3�ݙ ���!�oD��N+�yxS�&�Q6�e�*�ۡ�窞X�4|��;�͓B�S����ES{��oN�Sm�����d&�H�B��&�� e" ��Lӂ�&	���`��r6�f_~�> s�r-�9L�%���n�$mIA�׳)e�4y	�=��o�=�ȑ:��\�f����E�!�+R`0�L�e2W�p:����UWp %I"� Ci�noV�/,�ElG�lG��:sx���F��!"[���c1��ZM2G�)�]�5氩��x�
��l7V�:�o)�82�㞷��?��v�j���� w{x ���M]��f�=ʍ���G�^��ko
�9�vkn�r={���Ƙ�]��ΧV�qN,y��Mz�r=����[��������F��v��@�(""���W�^�$���}�gNŜ���,U�wAZFM@	��\��y'ޛ�w>�P�x�N�>��9d�U�nlɋ07��Ԁ��zR Yf��A�I8v�=�@�L��ACD�m�p�*�o�n�U*�9�ʬG߲�hت7PZ����d���V����XbH�m�%�����8�w͒$���i��u=Һ�	=�\�K��5f��X	$UզŶ�z�eT;�f$�H��I"�>{uY���Dfޔ�{��S���f�����$����,������%��L��}\ں�Q���vL7	�֕��=��D8��1Ƿ/70�A��I�y�0�A���ύo�����O��FEEU���/}#I)����ݯL�?}�~�F�����S�ɗ�/cT�`[)���x�=ˤ�)]����t�ڽshr���-Ո�1�Yu��af�/�:����pe.�-�(��Eɹgcn��S�@f���%�j&��t1�
�������wOGV�abu���7��2b��[�Dͫ�*.��l_V�/�/VM�͟A�LD�0n���nbE�v�Vh v�y�kq|��������>��/S�Z)E׌��9�S��'��|���M~i�J�O:��������P=������d������<Ǥ/�C�3�Y��B�ߘ�9����B{gϖ̄$	  @X@�� �O�	?�9�Oh�O�$�H0����O�2'Ē x��� �`r ��!� �!P�>�����{�������={��������	� w ���1�ouomwBvڣ�1�   �  w;�0N g�j�� .c�     
�/v�
�1�@c�����{�����;���v�ۼ����v������^s�p����n�M[oQ��x��*���׷�z��\ �eW��[�����wySv
�ig��S�KrVgmxz���RןT��g�۷v�l�]��u��on�h޻�E��ל׭n�k���/w'�_{w��{��.����q������ݷc�w�^�\�c�ٹ۸������3܅��s�;g���{9���Ӿ�|��/ki��on�ۺ��_8�����v�|�s�[�׵զE�;Qih�ݶ�]��^����wۗ�nn�yy}�>�Gt����\��wS���K��]�꺾��of5�z��;�s���ηw�־�[om��i�֮�v�{{<Խ^�;ݝ��o;��nwz�{���ze��;��8�zT�;3��.�;��9������{5��)�Z{U榌j%&C� wI��\aosq~�֋~`�7J�#�"�,NiT~ۻ~���w��������P���M�(8ǽ%uFj�nW	��z֓�����QQ�}�ȡ��)��F�k"�57qm�l)�т$��K��[�����Z�T�+�1r�Z��/�U�npE.���q�fќV^;���M���(6�-�)��J�6nls�"B@���s�F�|7�>»4��Lj�cC_{E`�U��]գ��m�d�ۆ�M\u�%n��{&
GT�E���~�.M�c�����P�~�Jo�0M��h`ō��q�Ǜ��i��ĔټU+�/Ρ&8�,�đuK�Ov���1��TP�T��	��<��q�ĭ��~?N�)�Q��Ie?r����b��AF�"�#�j7�uz�m��W���{]�n�ow�	���M��kd8��U�1��:�YJ�ѢE��0�*"�㕥8+�G�1uNM�lΧ����N]�x�^:�rV��ٌ�p�P��)"��<8`�����Ke��)�L��e��P61o#c�X�$E���<�n�#��}<��CG(�J��n�7���* ^�ߪw	WO	*6��	6� �"�M�]� 
�oy[;���������1���l����,#�9bo`����(��"��:�g�hz�A1R�B���w�t��=��J�,<]iQ"3j�@�yit��0���N���	8v�{)u.�[2:�
�#��}��u
{G(�4� @#I�I߆��)ZM�rT�����˘ya{ƽ^j�z�M�� w��a.}�	 WOҏ�mR�`�E�É��B��lō�-���z��zQ;����f�{�Ʊ�����&Q��c�I.��	"��o#�D�Ţ/�v�6��	^���1*�%�xwE\t�A6�*��~C�&�)���� ���;k9�ն*��ͭ��cB�윦��������H�Ȼ~�W��*Zɞ�zty�3e]��\3pK��K_	��b~*���JEL���u6����l
�����w��V鴪]� �   ��j��y�M���m��;�  � .`P�*�@କ�� *�M��CYw����~������5Ӻ����)[m�H�l��w�d�#�P�����H�L�o��}�7"T.�x����e�¶Zd�4؋=y@�qd��)����5\��a�����L�ZN���TǨGYn�r�Qs�"���F؝�`�H��H3n
���Ľ8���I$S�A�xdWl�J
h����;</�%N�\i@-X���7��y�mK���D�Ԅ��%7	�'��H��:�22�[V��(  ~a1����E����I�.�|h�����h����\��$�C>C\�B����19��ձ"$6��T�&Ki$Bb����lek�%6+9Ft5�y�Gfpx0��4"�Z��D�����V_���o���T��/q������n���x:�F��e���ȭt������������d��]@$��;Ձ(>MX��MD��՜#4�
8��I^!7`>����
��Z��"P�d�7q���lF��/�dX�&ߩ��lw<ɼ����C��.�mv�μ�v������.[lt�$L�I��m�(S�ՠj���<�O"��v����_=n]ogrs��ݥn�X���J�n�����M������w��n����n�����w�4�gy�Q�o]�ݹ���B���i�o ��#�E`�V�b�V��A���,d��Ӯ/�tn�,Ꝙ���I6�l�_e�[:��*D� ���K���w&�巡u�]���tFq��{̠
x��\s�v�e,H�Pc*!��Ծ��ԡm�fw�R�Krk+��k�w([��~���En�.�B��-(l��;�G�`��U�>&�����q��b$k0�Tx����F�: �U������pn؜~.�f0�gm�b��TM-z���W�Ժ�-�A�3��<���6�D"�&��ll�� UW�۽��RA��*	�4-�p���v����2$lb�A�~���K��:�CF�J�<���H�Ď��QSpl��	��.��y�aT��z(�ǉݜy��W:tEc�g�����=�/T�8X('hS����vp����n�N�&�AG0�:c�<��s�[b�6\��~hg�С���ߋ7�������5}����~�+�xP��B��|�-�-�խ��L�k��`����B>6(Kh0�,$�b�T�&*	�Q��-W�����-�K����ߦIyrȍ�R�Z�i��]�ym�]o ���7��ʏxm�7�	���uڱ�q�o��4��Q�}`o�0��vk�u.�k��C�k�)v��PH�r��*]����$*`k6���qEn��n���I�BE�Hn��C�xL7,�j��� ��aޡ�����7�gY�,����T�u�g�Kk�`=fю��7.sIu�B\*x5p���"��_:C�	1h�y���n��\ �Y�e���jE��&�	̬@4��-"�A�d�K�^���(B�&Os}����)���X�)%ȇ57I� �:�c�r�nc��.թBhm����� ����%D
 ��/�� &�I���˃����	A�0�$�%�{��Ѣ���>�3��	�����I�_=p�eFc��ߚ*��*5 9�s�Ve��md�\lR)d!�%�6�R-&�H�9�z���W1��<>�w����R �"E�d�ʸ�	��WA��]�4��t?Zŕ�Ʉ��D"�Im�S��a�-���u���qm�w����|#F��\ 0��.j��R;�r����:ȑi�s6�1�'t�ň��J��%"�p�A����[&.z`��6q�_b��'v���7��#�'��#c�̞O+4�(�:��nH��K�K�u-��m"�@�t,`�h��T����v	�����ܦ.�.��Sw�P\L	D�lv�6R~��)�pSv��	��c���;�nvMKH� �P�0B$��($�Nh89��l��#-]���ٽ��GL�2��A�.,v���k��;��Rz$��$.{va*��m�$�d�`�QL�w�x��w�Q�'�,��"z
�iBf��x�u@#��>q1j��98���`�F�*1�˺�7�H�m���RT!3Qq����S.�tҺ��������W�wwv�Gp�O�` �g^���?b�WV�m�]�P   �|������]�� ��*���B� �*m�@� 
��T� < �[kr�nǵ���y��͗��w ʵ��9�7�w U��ou$C*��n�O��W����� ��0��������A�ц0$s�^�Ʉ`�!��Lїl��I'�BV+&E��B�j'f&#+��&��dFQ�ф��r�T{�$l�V�a<�bo+4Tt�q�d��)9���OWo �c�Ƿ8+bk�/�;:����	������ƽ�! ۲?0�e���$����=��_l�b|}��ײ��Kx��'f�V��V�P���(Y�ኲ�sU����Cbōl��:5mߥ��{e�p3`71X`I�5��l�	���8C$���CY�z�mF�UP<#A���\�åe��cF}����Ȕ���]�z��* X6�Kl�ۂ�! ��EUzUp�tMmݵ��LTp��c�Է������;[�<����G��ٿz�fgC\�����I�9Y�t�F���}�)yw�����^Ł��V54-���l훚��n��炏�����T�R������Uݷ�U_wz�����x��nuˎg��呠��z�s�w6{s��sܯ�n�7��ooj���R�⽩���P�<�b�甩�r�[�[���y���vϏ�(q�8o�)����Y"�2��Ԏ�|%J=A��fs������j��P�e�͢��0+��^4ZU����	�)J���H�ᾃ�ׯ���CkP��*���8Y*Z%5P�wn����.��^�ocU�L��N[����m�l�����	E�: �X���S�ҧ�ݶyʅ*}-�c���=�7E4��h��ә%����I&Q�Rk�]�鮘n���o�b���&���n��
����,�I�s���
�y|���5�4��6V�--&�l��@�T���`�l$���l���0�~d�	lDU��IU�Eq��طћ��1W��R�Ui��x�%��!1S[��<#,�=|4�9��:���$b�Դ�����&V6U��⏸�|b�g�kkx����^���ם���i$�(O}��TX�k��ɞ&��*��T	h�?y{�z���ߪbS�K:�HZ�k�V�SoW��Z���V*Lp��N���c
��{z&��rF9�cK�-&KI �v
����W�u��w{��u�q����y�y��#���5J�Q�j� �Ԅ�x�lE�g�8.��hӐ��O�=���b޹��fHQi&�l|#r���(f��B4\ǃ��.#�r�й)8X��ױ����坳�j8���F��_���% H�i&C��� +����ը�!��Q7�o��Cx��<��߂�z͋��&����������F�D��K���<!{l�HG�i%�9�p�e��O9Q᙮b��*��|���'�}Ʀmy�
�L�����a�N�qw�~f�'y�I��!��Q�%�pu�yfŋӗi켡F��WC��T����6=�x֚��aF�_�PwPA���D�&Il��t���޼�=: ��!�FC`���%2 CL�.y��$��-�_��5�DCC���� Ӕ������O1�ZO�c�S�7k	�	��BS�#y��"��&�lX0��GI�h2m-(����5�Il�wSM�u�h��1�!�\��mlY�Meq��PB�s�j�� FY��v��3��n�jlآ�khI�� �h��-�W�=� �j��-09��M��91���h����K���n�P��q�Lq٣�	9�����m#F��d��8!��@�+�nw\��YV�p�K�V�~��H����M�R+�y��LR*�Y����E��U�SNUzD�L��\Ԑ�=k�6�q{گk|,��
�uYN��_P��Ah��9�<����[���q�|��J��I>�wi{�L�Ҝ.�o6�kS��n�.^�����Ʊ^ia<$p��u*�}}6:^�<�P��r��������Bz����g��IPJI������7�م��>�b�W�M�&��p���\�(�#׫�ybUw��h���b0Tڨ��?}5ן<�~��%��F:�k��o[��;6:�&:�k+5d�,t�,<=6^~[�D$��S�U�]=}A��(��wd��ޭF�o*w[vb}��ےj�&IY�"*��F
�sJ���H�e������3}�/93WTF���L|_F���Vv�ڮk.EڟXs�����I�gU�T$���5u!��m�ݠ�uD��؅q��9�,��O�{voui��nI{s*M��[�u�EI�X�Ưgfv�>�QЮ�u�[Y^��'�wu���*��Pi�tϦT<��;Շ�"���y$}_L�3�xY!��zAI�?��'0���I�X zO�
�~%d��s!9'��Bd��� (���H+������z���[�:�V�`h7g�$�I$�I$�H �^��5�ζ��J�{=UJ�]��� me[�����s��� @`����  �
�PAT�  2W��EUP*�F�u�� z�@T�� zuPc��   �am   �                     T���p�%�m)ݸ���mݻw�]��[�Swf�m�v�;��L�.k�^�xe.�Ѯ��u<�    �   �    \�  
�PP*�   *�UP 
�  \�UU�   
�Y��*��� ��U �@U+m@   ;v 
� �� C�   U � �  8[.� ;�T   
��U �    *�P�s���M��~�gnn{ �*���  �e���F��գ�;��Q�����;���%���yg��6���fu A��z��?l[{*+ �   ˷�s[r�/�f����Cl C�sU�P� P+�   w ����uuع��m�V�[`�s��_�u��Sg�W�-8܆Nq�[�	���Dn���#^�v���Z(�{�U�wg��3�6����rIV�~�T��d�r��$�%<�5FxlL]quW��b��ł�h��:�b[� ��C�������E�;�Omp����:��	15�����g����/����ՆH0����#*6	ҵ��ZOY�R��*�\lt6�����U���C$&'GY��G�����Q[���n�ӑï<��DAWa��}9$9"�}6-p��ռE��%��������w]����:L�O�nCFw�O5�&u��m&PTj8P��[]3�j��"-�gzǇ��X2a{GBo�(h��~%�ތ�K#p6x�P/a��T��U����z��EwUP�m�@�(��i$Z7�lp�=M��H�ޛ#t�=y�æ~�*�v�p�8C f�;��7-��v�[�WSn�"8�>�ۊ Y�a�<x�볕��){<6]ֻ�,�>��1�e�9�K�s`�r�Y}�f�[�k�^�l�)Y��� wn�T�׷��z���{�ok��y�7Δ�+��Vw����㮝��׷��u�׍or�[�ų^�]�Kv:�[ͧ]��iFP�0ʆ�. ' �2�FB�c�W�#j��Ļ��(<7M�uF;늍`�#N<N�U�v!�`�rD2��Qa��Os�-�:iPǪ6=���w{eݑ1�S�1���h'	�I ����{�JE���CLt7��]�@K�[,��s�ԝ�;�c� �A�	H����`�I���X��n�Z��"@�iy"s�E#��WV�������)����-��0D%���8�l��D��L��2���tF�msG�Nŗ'��2��8�\�T$���0f��$�����3 W��w���U�~�����7j*���U*���ݷ�-W���w�ӆ4`�xOwTC����Z�88S�"/�;��V1\f�n��"����w[�2[��#|��gi�6�-݋�����6��}��ݔ���,U[1͕�G֭cY"Nb��F��=�K��j� $�ĺ�Ki�]�kx.�]%A�V���C��70��IV�����y�\�d|�vk�髵�dqj(��;ׄӁ����2�թֶEU��1┋|����w���Ǻv��1eI-6�Q������GBMCD�p� pQH�!C_ �`fakFJ�t�9(M��P��?�W$��]!8����oX��4Rt��+93�a�����IN���H�7�s(x��ץ�
=gE�Վ��L잺W��u��i��}J�-s]#�G���&���NDb̉��X�~���(&�$��P,H�[m�:ܲ�p6�^��V�2ar���"<�^:�X�>�:#��͕x="5Q��1�z�!b{oBP2`E�O�m�dU4�I�j�Fu���pLz�Oh4/��(ƤsB�2O 7L/|��=�����}"ý���a
�k��f�f	Ѝ���5�t�|$E��i`z>���@�Z����;A�$�h�T��s�\�^�Fp(Ş_�j�Z��I$�M	�M���{mC� �@P���,|�E��H&`Aq����&
�lNʷ�	#Tp#D
�%���ŋ���}P[��W�k��0��Vh&*ҍ�/"�/X��7xߚb��8ZN�����oףD6�-��,Nf%�f��L�m�$��;}��.+�L�Y�1����	�Gk�܀y�۰(#<[���7�5I*I7@;{��;�
��Ѓ4�D��e�=��.��5-t���y��b����"�wF�M����4�}�	l&�ð��wUS�-"��g`H�<\�H�Ӓ��և���cIt�{�Q�-�8s=6�խNY��o8�g��L��V�I>2P��?7�f�c����X��}=��ԡ3կyV�[�cW�0��|�Z����.̛�cÄ�'JCKi L��@��ݵ���#��s����͹�H������4�C�Y���m�G���k0��cA�0�_Ν�P�V�x�T�AI���$�9$��M]Z�C�KL��^l�l�DQ�}��n˹�:^G��co�Iv#Ñ�=��=s�d wpc��b9������I�޵J���X�z�rgF��9V��@&S%�ݥ.��6��ug��~���v��l�U@   9�vm=ݒ�=��ڞ;��Pm�� �T ;� �M��pT
� ��f�-�+�w��*`mM���ܢ��@*�zD���A[5لԬ#
�}2_�4�\��#�N�!�=v�܃]�de/�LK訚���!5�o��f�M�
�a���Ќ �;��W+z/}o"Q�3���00��[�y���wf��Q��1�kxB!�����њ}�QE})��1#oy�>����*�4�:�nc[+�*(r�K=�]rgo9з�8l���otaA+���f���JIi�RQ�ƕ����,	Af��*!7�?>)��$~rڌ��{W��e�z�G�Ư|��sf,B0_Nr<�Mj�pX���zaױ�<�ّp�i\U�Úo���0�1e���v�]�S{%�((�v3�.�2���$k��̮�� H��"�v��H��y{�pM�eyZ�����@���m�M���N�P�e*���z��")�I(]�~Y�'Bs1�q(����7p�fwR޸�����{��)x��}} ���T����a� ��.���Nis"a(rh	f���#�w�1�aA~?�+!���دc��/����#�wg�ݽ7h {�o7�@6�x�������۫7��=�Q��۽z�y�������V�7�����y�g���{�N�m��׶���aBh��&
Ѓ�$a� a��Ci�9�b�%�r�Y�:�%kS!h��`����&v���[��쎹���v�0��'��Hr��ZhWr�N�8w�Gr�5w�B�_H���|#E��Rs��S���"�A�h���6�J�)$uY�]�Ǣﻦ�lr��[m���2r�<q׎���F�#��!���Ƨ|i�u�r�ҘޕzT���E��qm�W�?1�1c���@�(�&',�a��{��y5�t5D�Qc��K�eZ03��ѪS'Fɍo��y ����"������Y�Y�rɆ�I m��m/;�� p����o-��$Be42�v��=d)�ͷ��M����($��'uB���1�5;Y���6�wͩ��e����Y�:�єH��M��beX�?3Sލ��-[S���#A�8>����qS�"�SѢ�'��Yl0[�6��,$6v�K�]U�[%� Y�V���4�ϳѱ�@�۔5IZ�<���s���&skT)���Ҁ�1�D�%��O��\�.�Lb�&���\5oo�{[)����^R.5ީ�C�LSf׌����{��ww��ou��=n����A�^JJ���'���^a�v�%��Ջ�PI�em���t4���� �a>�1������e���3�L�����f:�u��]h�d�5Gz1h��[��P2c�)�|�7p�$Qz���Ww'��/�_c҄�S-��$�n��6�m�J�n��&�m$�w��F�K��ި�0^N9kdU<�a�����fn,�d���Lf�$f��44yjX�6�J�{S=ڄ��}R�N���[:Ó�7}/h_�t�g�!iE9]�_��V�n� �hm�ځ�x=��xd���$�������#*;��.tι���'8:v�ӕ]���LFzH��]�4þCF��})6g	� �x��Dr������9b%�98`�J% �e���4I)U��bJ�����cd��wMk�ښo,�>ŋZ�r/C*N�~cǯw����m�?B�yi���]����ӵ��z8!;�h���X�&QS5�ʢY��83Ld�]�:«���o+�5�*���3�Z��'.��3Va���QX:��*��aJR_&�-�D>d4�I#�[U}}^�Wto�����ҡG77��/Y�0Z��0wb���������Yͨ':MjC�D�)�p�z��6�e�ZV�(O����eh��jj��]=��\�k�]�����qm-�,�o�5�=:|0-�^�rC�w��T�Jj�y��f�o(�����9lGqU'ws���I���\��r<��f���4f,B=^*����I%I���*����r� ���Dq�@�V�.N�St��3�0I�4�W۲a��xJ?`���r"�黒����E��!>߰X[�׉&$e�I���\0��<|eyB�l�ȱ��&c/ܲ��;��3��*>��n6
W�N�W����{��g��Hi��ͼ��{�5N5� z0��6���v�	�m�)PI0E6�1w�6�Tζ���Sm�o�E_�`��   v�m��yx�7��6��`  � �*��� *�
��
��n�UV�Y��w�M�ݶ�����p $� �Se� 4�A1��?���)��ދ���V8��[��~��c�V�Rö�T�i�����)��#����!&I�Cb_����V��[1��x�c6g\��	j{�1$b���C��a�a6�4�ʨ(q���=m'��B^�	Q �U_[�'�p@��g�̅p��_���e���:���}�H�������JHJn!�]�޲&/��$DKd��ゾ2� u���۽O6�wOƮ�����ǲ%�
�4,!"�ޛhBZ����Ay}��{���j���v�s-M ���`�b�4��*�?����O���uZ�ĩp疞氌�pI�\D˞ E���23�O�1wWt��_�{�^��muwV6��^����P
�U�Zn��]��1��nl��.��h[J�f]/|j�����$�֓��=P���%n�z$���zP���Y�Jm�и4pܗ�W�z��ۼU���qUgw����T�8�=6�kk���nP-W����` �<�wU ����M�=��=�s������>�ws�sݶ��q��������mOT��\<�G�;t���m���n�];ݽ���*�w}]{{���t�y���Ͽ�~d�����*;�3�4x~��/Ț&y-�ޒ����;�c�wpLO��b��[!���O+��*V��Z��=��W�m��y���Pb��!(�;i�k����M�Ҡ��܌��H�B9{m��V�< Ĕ��xV���m�,=����{����j��fq[�oX'����:~�t^��)�6�]	�1�zI��s{6�ua�Q��Z��[w�L"����b�����h�-M���[�'n�t�W���<�T�cef���ǎ�H�T>��=ް��x��9��`1���he$�H�%��]u@�T�m���d`��C��\�y�r�5[��X�mj&~~��r��޿[��3�c�syFY��GԒ-KrzxHk2;D����z��M����eO{ŋ �w�@�oU�4�ck��Tp����Jil����oC)��o]��6�-��4�!�T>�\��x'�xV�?����5T*����r�z�9�lW�b-�,Nܮѭ���a�i�A��B��u[=D1�@nL�)ue�ӔRy��=��Q�����8�u������ct˜��9cB�Q���O��i������U�r��2I5��ɗ��[���t��o�]9�1^9.���2�h�,�YZ���Y��fP`�l�9^vv]W�M^N���졸�YP.�}�oG']������ga:�!e��3���]-+]�17��ݹ��-����;��8 ��p�m3?T��.�,��%���S�o>��n��[�G}�~�����o�>��	��C���H��BBT$� I>$'�!���,���V��9	$��}aL�� ��I� E=!�C�! =$���$?	�rC0�VI!�Y��@����!!��$9OI	'� C�'�"�$�'�O���>0�� V!=!>�$�0���
�>X�G�>���	'菑?@���8�C;�l/�Ҽk�5$�-��m��m��-�� � 8��T�o&sX �p��  �   ���N �JT0�&�     G���  !�z�e[�o���;����T�]��7�=��om��w_>v�������^�w>��v������u{L��x����i�8�֍�*��-uG���+�7m�].�^�Q�;�xj�l�dN+�v�������v�n�w�׫lR�w��un�=�<�|�y�rU�w�Kz���oY�j]v��.��n��Vݧu�W������oomW[׹����+�{ᴮ�ݼgz���۾�ݳm_Cg����^�vv�קG�e��/9ε����ގ�ש�\v�^���ɋ��v��]�z��[�;�v���g��]W���w��z��tm���x{��׭�5vx�T�������j��m�^{7���Zx���4J�)����{���o�����v����޽{5�z�Z�ݍ��o;۲��G��]�˽�n���[\>:���v�`��}���g�c�J�2(Y/1qS!n{`l$S�N]+Bǝ�4<	)!!�O_����h�V>�F<�/-���D�A"/��p �Ÿ8�v��Δ���=�y/2�x|�7�=������<�.&Q�>x,m�-�ǉR��tM$����鄣�V��Gm/|<P瓵�����6L+��B8Yh��j���w##}*;/L&��9h�2��z������j�*��$��D�m�A��I���;���РF��\êK%�7�7�<z����\͸���^�vŏ��d"0�h�S�ئ�+�E���'Yu�*a�gtcR���8�hj���3/r��4� ��x�烱dC�{v�h3���E�Km��LO�ي#��J��l]{�_'�[sօ���P���b�d>���f�2s����Ux�@�m�(L`|B̚�(X� (j��M��1I� �>"I̯�ؙ���[˾+K��w�ZwZ��z��OvF��BE�Ѧ�E]���ʔ2;�>T�41yi&{|62�N}��s����cOY ��A�!m���z�b�6"�U䧲���:IKp������x@�-oon�S%nZ#u���5��� �JY�d��,@�Um(-��Y����V�Ϣ+v�Ϸ����L��26[%*�˱}�	�S�hn�x�_�UsF'wr0�	;�*���JP�L��:���o<�#Nb�e�����f��l�txvɽ`�P�P�>ya�7x1�J�-�2^M_Nɉ/ac���N�P�7d����/��m&^���T<��v&*�koѥȂ:ɖ���Lo���3�
��!���)߃\�r�S��[�`�1CM��"	FBT4��a%���-��>"�nr<�Ξz������1U�$�\y���(��T��0E���!#m$��;�"��< �w8�uV�=#mML�L��Ǳ���M=F/uGrN�\�m��7���ٝ���:k*������ʊ�f̮3d��m�ꙥ��`�m������g�*�]��J��UT   *�^�����ޛ�-�˺��6��`  � �P*T6�UEP+�[ Q��ĜwAWGu�'���߬ ���c�@©T����)˟���ܠq�(/J2р�囓�:�[+l�Ɂ�����57�.�����/��4��n8�s(z��M���f�d��{�VT�ۼ���Ћ��A��1���1�G�^�z�\�ײ��I7qվڎV{kwn���D���ÉY-6�Q޻9�����'uTq�cF�7�D8�4�K�O��[#6��l ,��=������p?�{|�*��H�R����?��>yL���%3�uu�n�"dLǧ�z��*���IjF����-T���zl?�����r�k�3���`�ְFo*�#�� ��Bt(��Қ�|Ą%�95'���岅ڗ+��[N��"Eg�b'}��� TD`b���މ� �$�����Nni�slb@@�a�($�I�j-�of�T)
�kҥ}jkV��*4Z���yeS> ��]����Ȋ��� ��0]�J�$̴P-Nf^��#Q#�A���uN�u������<���4q��-Y]O��1�'�i�m�D����n� wm�ު��;��5�뵭:�+�_�re�|�w���^n��w�Bޞ�f��ջ�˭z�%-^{=��S��w}oB�����ݼ�w�w�w7��%�e�nM�E8����:b?c�����9��+���K�X�� @�˭^��EV���
�I�J	�a������Q*r�1��U��xM�mZ�z�<xH�
Ǥ��;b�ti	;�~Hn���)�i�btn��b"o��	0t)I0*�hAi` �L��P�=f��{^���3>U�j���\,X�n&%{Q���\�n�Ї^�S6�~RK%4J	��}k�Φ�Q}��"=�ݬVB!�)�Âx�U)\��/� ���G���i�\I�AI,�[&K�CZ
���6�W�� 6I�H�q]�O]��Sf��Fz�����H�US�1��&8\�`e���@�9`��\ݶ��r&pbQ$|�1>�J��;�-�J%�ѪY����#K���b����a�	=�����baQ%F�~�`:Fwy�q��Y����������ق��f	��r��ڸ(�hݎӮ٫��b���iP�7e��$�Ќ�@Hc�� )$Q�x4TlT;�ǿž��u;�:쫣�<*��� ���N�C�l�ґskZٙ�V/ Ɠ��х�V�~�w���_��H������`I�
u��Ä^����'K�T뽶�EŸc�CyJ�Ď�p-��&�7<	I;#DPr	�n���d�$4�M?� A%��B��U-�]z�?~�����ߎ�h�C+�Ta�y�*�[]a��"8-�N��@�Gj�>���V*Kn���i�H�#�ț�[E��jtv�w��jU����G�"Ǟ� ����靍��6#B�G�_g��E"��m��˸���eVWdDmW���=j�����?^߉�al�5r+Gl��xe�Y�crL���vzun�l&���	��08gB��~��/�j��V��k�G5q^1���H.�x��WFxȁ��Ũ��犑����T�����\�BΕ�P�V=2��zv�q�6h躹�>~���1��ٱ�z����ȔW�%�/�g�x�EV# EG*��3@�=�d��|�+BE�^/'3���!=Ɣ�&���b�i�ZH�M lknΛ x ��ݽ�{hRA�n3q@�Tv�&����uU��W�3����|"˶f���"N���W��}�4��T�Q�<l;�H��lAs!�^��ɾ�ǖ����b�VQ��C&��
���D��:��덁��I�L����B������8 $����{L�ܯ2w�z,�$k�6!�v�&��6۩+��Ks�ߦ9�����M���6�@
���%<�y!�g*��]��� �0� :��h��Bd�D��܎���a�xg�Ё�S���U�;p���<�]/���u���͔=�z�q��	f`H�Im�)�����a�C�^Q��S�.���0Ud�9f#��]ƸR�4°3�n�] 7��*�_�����N�`�{a���ļ�9��Z��W�)ɽ�[i$4�i&�%�U;��YA���mkf�{_�
l�   u{=�o��u�n�wx����`m�� 
�P �  `T��Tg�
�`��C��7�ۻXڛv�@�U�R�Z���i��%ߣD�i07?��ծͽ"�߁̝	�$X�:Ă���+���")N�{�O&��~j���8�@$2�����Z_L׈�*�cQ��ޟ�'�b�Ls���R�vy�-a�]�2O���0
�����I&�p���7lV��1`w(�^�=m�S��K�������^i1���'bN�R���Q�H�V[���풪��& P-  P��a�`�\Æ�0��u��9QR�.u�nǛ�e�驊{���DQ^
�����p��l���$��4,9�a�R��P+v��hv2��UlA�V��u�6�.o�B�cf���иGa̞�)Z.�!<y�����A��%d��!�u]©T��n�wA���r��g���4�`��6r���N�X"��)
Pp�s (��PL[�Y	���d�2�i$��7���Ϩ��D����.'��^��Ab�~or)�s#���Λ�yj�Ǚͺ�m��4� �w7���<�q����}-�ݻ�{{s�&�V���kn�n��mg�{Vr��v�=���/	ͩ����\nN�H�HޑW��{��j��"؄ ن����cAV��䵲:X�(4@��0y��U󰝨���u�WLu�&fא��R�� ���)C�2O�b���X0<�;�\Y�E�ȽR+�3�����fl	71�E���9h�M2f&0H^�/��[E���j�k�j;���6D��������<!r~��@ Y37)bo���o��	�>}�����|+#4ZF��pa3%��"v�DƗ�������X>ݒ�.�K��)�u�пs��T�m�>��g�$�J��tX�H��P�u��Z@$ۦ�;��[ wB��Z��owj-$�g(�(��*�Cǵ����DC~cɸ�՚pk~pm�����Q�$���{0wC{ʖ��Ùs�D���Bw86{�y���~�4�ތ�~��G�ӹ7K�cy�8��pðQiJka�D�5��i�����;�#��`�b�T���g�cmō̮~���=[�T�%C�����a%/��V�
�u��p�u�֗H������#`P��OQ&���Wcj�q�
o�H �I� ���-&����e����w�gD�W��
;cJ����K��!��o��5�,�Л�K�pv�[�I$$IM��|Y�F��rc����n����D��6C(�W�,\+�u��9���܅���8F�7jy��"�-�L��{�9�J���U*���m"[D��b뎈�Ѧ*QF�8b{���*��1��p������Ѝ��yr��� �.���-�q�!"Q%$���ly�<�.�8�dv�lF��W����>����Z*�P�,*��,��=��za@�+��� ه���j;Y��mt�f�5G���q�f�#p�7���p>�b�����Egw��G���J������5�vG;l���u(�-���T������^U>�����;M
�󂠼�@3�Ύ��Yn{�bZ_�[=v�ܳ��d�gDe�ܜ"F�
�����m$�U� F�yA�����')X�a��|p�V/iqsb�}̞
��b�	�P���H��2Q� D��vE���M$�i2�8*��ʩz��m���BD�Ga���;����c��4��Qzr�"42�r�CU^^C��]����젡FNش)�NҾ,�y�r�i��i$
���2��ޕ�V��{y�9��Z-1X<O�0��Oi�9�.c;cĖ����p���a�s��Hm¿Y��f�
�7�*nE
�9§�\�^N0a炅~!��f��U@j/u��{�H����n����b����,t���.�@w����{��U͵�yu�޼���x�R�8��^ݸK�Z:#ۋZ���^(q�HS�-ϳw�31XP�;/�:H$�J6���=Ջ�y?
c|dF�C�m�~"�=lrfW���c��B���65�܌g^(ȏ��.��n��\��h�e���l��d�\D2̔"���'[%q�p�L��a��޵��K�w���=������#s �7(��1x�Z��ٵh�ڍL@�����.���%��"��R�k�f�N�Um"^�5�*�u��@9u+'}�喫�mn$�9w��wn��t��޲�z�D�p��,��Du�j��`�Ȇq�g���+^㫺��6%�#��r�u�a��|fn)��Aivu�c��e9�9;5�6�0�]��2�.�ҡ��0>t���v��V���0Ԯ�c:�f!v�ʠ  �Zb�ݽ*����ϰw
�T;������*�@�lY@w
�z��T�
�*�� �Pz� Q�J�t1n��  6m�Mj؁R�� �ջPqT�m�T   �ե��  
� T  �� �              ���/owz��I��^ۻ�z��f�ڴڻf��̻M{{5��Uj����<�]��zn����<Uݮ�n�   6   ;�   U�     T@   ��  r�  ��    `<U �U  �@� U
�P  ;�   �@ *�     � �  ���
� x    [J �Uw@  U  
�P�y�ny���3j�T;�M�   �Ͳ�;�9�K�����]E~_~��᷷��޻�w]�.�� U(�{b�^�����   z��u�onw��;��Q� lP�Sb�P� @ �*�p p�Un�f[c�����?wuUV�~���]�q�qRm��P�(%�Qe���>��D\(ډ�>"���u�E���mL���c��ֺg�y����Hާ>Wpc bj�D�Ye�@~-�zh':u�	Gc�
Hj؀8��-�75�`-R".�rt�N� � ���^���̷J��R���)RH���u���A$�B��+)��}v�������y%����Ȥ���"�L���bD������`��[�B!@ *$Ɓ��T 
�LRM2à�<�NS�CUhĜ�ݣ=*۸��z=���4��5�q��iIp��V�P�yPd�e�Flh������+�����e�����]��-I2Mr�9�0*��[6�X �6�;�ڭ��n�!8(U����e�~�^<�=�n��V���Ww	�l�)�^ŷ;;L�n�ug�v1�+��\m�13�����,ѓL�r�
�5�w^,�I6�((� ��sZuj����z��zu��IӺ��>͝���m��vg��]��tڭ���綼�kWv�{y��xʥ�����#��k]�r�6� 4�m��P� �����M��*�W�A��{9��{�����%�TQvi9i��i��cu���gNU�w�p:�Dۮ�.��槜p]�Q�OTޕ=�<�I&B��ۼf��j�ٝ��[���^Z��ޏ[�٨��rw{�=:��tծ"GwU�[�*�[ץE��|3.}�/N�ـ�^��+#��G��xD�g���&�i�����U0���#
I�n�xrھf�<A�|�E&
d��z�׶�PlVfe�u�� �)�T�:�v���I�;���:�Rޮ�6�T����.�mZD��ݍ�+��:5D�f���V{��c��;�@�ڀ+`����9�݄�7��M�S����b��E̎E��}�53U�7�`�z�x�zq��Y�@�Wea�����.��+b^�L�WL���F��y�1�&��An�� @1B�R ��n��J1d�\�I���}��w{l��볦g�#�"���ݜꍜ���R���o�z~ɵ�c�x�ϼ�:K�E��_E�m���X�.�"�M6ӛ���<*)�U��'�O,D�U낺]����l�;��&`���^�t�N�E���5t�8ʒ(��I[m���%������W�^�kvy��Ə�Ηέ�rWJ%%g��I��[x<��y��#���)TU��'p,�;b��	$�5z?e�����<k�|����U:Ҙ�|e�ֺf4}p�1�}��z�	���w-�QѠ.'F@���Y^�� ]��*2Rba���*0�+�׊ �K�\�Vv��/��8_�<Q)�J,O�6���IT 6�@4Pa�M�@�PH_"����D�v��!쎶��B���o`�9lٗ���3��܀6G�b5�ܙ�v�
(���9 ���^��Ř���cӤL�`,��.Ozp1��7V�eP���,/D��7�'J�F�ځ��2��u�������L�X&Km������J���(KM ��G3�����~��ݜ�^�u���z�{�l�
X r̴�pKI$���,�ݾ���S/��5� L�׫1(Z&V�����^��Jo5�7��뻭~���H�0�9}U���c=^��\��]���Ծ�h�����F�xI�sI)���W!N�izY,��H���j������+��a�_0�	40�V܎n��_^-7�x\0�>��{�܋�l"��%�H�{�H�� 3���{��y�.��\v۾2���O�$] w�@8��{zD�VNZ�W�<gZ�k�&�����+r�[*�.������3����WOw���UVȪCȭ�����U6�@ ]g[�{�]so;��wU��AT6��`�֠����m���z���;�R�˥��UܛXq[2�!RI$2Sm�C�ݶ�YM�Y�C{�ԺhOvc��L��T-�&;r}��(���͡\>���a��d�?Y��N�.���y)[��ߑ�4�u���q�4owmIn���R�G}�M)��$����� ����c�`�{�֦hm�ȏ��W���{��X�iY4xe�QD�)�e�$��z5XPw.+�{�� �DPR�P���@�P�D8i [ ��;69'9�
T!/����vv�ܫG�lO>B%I��>��ڜQW09��0M\1�c*���J M�J��H�c�
����;�v�=�%]"ܸ� ؅�#�S��]���a�'^F���m�H�V�����n���㿋ʶ��6��Y�i$�-#$@4[L��
��n�\���>d�����K�e� N��k+�\g��'���v��7�Y��l��ęL{l|��+�h���`��~��Uq�7&�fkaXL��Ђ��.������D��F�B�JΩ�P����P��;�Ǹu�����_w]��{�ƭ���z��y�'�����<ޗ���g=or���m�v{�����g��A������u=�((�-�-!`� ��+�B��������bѧ>�ɚ��Qb
��R>g�6:6-wx����m*G���uQ��7Bz"ʻ<6�âa;���2l��}�MMs�F�$��X����h����Koj.���F�&�6�e����0}	"`
R�j�� h*L6��(1M�k9�.kv�7�	w��#gږiZ6bՋ0^˖�FVѐ�x���G�hܖQ)"D���wR7�,�>
���,�Ǝɳ��̫cb�3�Q��k����w�/xbf{�qe�*yX����lp�
@~�����{P��e6�I4��  )�HN�Kt���;��e[\>��+�p��yP��2kL���3�H��u\�����V͕�C��,�rl�JI&��'����^���1Ỏ��f���,h��⛍&�X��	Y1W�I�
ʪ��rި!`� �+{^���0A���31�9��N�<�&���$Qf��a��kojsd�NT!����(��N�z�f��U�N����jc�'9U]D��M(M6f3[�,���{1p���+����ݷ��ý��8���|�&{W>-��M/�YG1����z���;W�,��:�0��WMy�D��l����!n�ͻӮ։����!�[F#]n̡`��?p�f��U�c����,ݟ����ee ��(I6�p
%6� ;PUm����wy�U����ɣ�_�n�;6<hb%V�#t��,���9*4�}ce��Xȯ���v��i��]9\iɨ����}l��C�d�~���߫�@�>��ǅr
7~���Rtr��lҬ�S�٧��$�)��cHk5e>\�H���$�/,�"d�<��Wڢ��p�D�%��R��%"Qv�UN,]�~��tWM0�-7��b��;���d�XH���ַ�U�v�y�}��z�o���H�:��֕)8,b��^�O��&�n�`�dg�,U4���Y�=:ٻO�Y7���G��{W����H�I;nl�	��n��I��@ho�VN��r��&�`��i�F�(�a+kdJ�<�I�/3���� �-�/�"dd+W���HE"H���m K{ m����V�]�l�/��Tc�|*7C���<�k���&8F�7���NF*m��"��a��Ĩd�H�W�) y��h:��Q"�$���OƖU(���+�e����kdVƃZ�k{�%w���!'1���v�f����vJ6�HkF�����[�5&4�N;w���Ƚ%@W�_���C%�Y�{�<�&�ݻ<��J�V�$�U��G	���T %Z�0_�P@	 *I�� �r>����<�o�=5�����q{N�2�m$9���:e�m:Wbl���m��Ja:�b���F���<N��g�I��*Ʀ���L$����`�sQ�(v�w6e��8��:pta��yW\΃Nָ�_�U�7�z�]��ⶡ�7�ߝ̹�h��m$�0��N�'J��p��
�T{f�U*��r`[[ �   ��t��z�g��o`6�l�� T� �!T � 
�/Tؕ��R�fɛ`��]�l}��oP6+�l�l-�z�U*�H��M�Z�� ��[�;���\XVt�tΩoǸ�=�����3��ӟT�s�09)��*U�A��i�a�=��Rը$�$���U(�ն|i��)�P��&7D2�L\�r4^�k
&����Ny�����	�H���I>��X���H)�q�0w�T$_Y9<>a��p�&�`�Mly�Ғ��S��,o��tJ��(��$������4�J-"PLN�6�F���7wWwlַZ{99������!8p�\��a���Be-�`�QÀ�D�������B�qF���)�h�:�q1��GU�Ē���/:���}o�bcm:��/s���9�@���n@������������v��\X �IM���гͶUA�+7EbI�Ki4�	1���L�ޏ[n��&c��ie�'U�(���Z��^�K1b��D�YĴ}�+���Ѽ�f9s�a�� �0�i�7o���[����r��J,�=��f��N6�ϊ�팇�&�\Q^[l$�2�`4�m���۹��j`<��W]�p�oo3����z���_g�^��y{s�Vݛu����{ݻ���޽����wj������������	���u�$��" �F)l�$N^��k���m�Y������f�B��<W��4W�(��'��g���A�&�f�W�>L�w�X|�%���v�C����9�'	�F9Ĝ[6��1 �T@�m$#���gBБ����J`D "L|Sd$�2o,[靡�I�8Ǯ��sn�o<Y�F�d���A�02�@,��վ>H"��b�h�3**�A$�qQ��n��Of�,ܘ��5i�F؞��Ǽ�����Tɉ����ȏV���,�*�X��GR��XP�P	�����{�AM��E��]�R��I��_q���ms�Be���M�VY7�yblg%����u�Ly+c��}�3^���LY� �$�Hۂ��
�Fɂ'��{��蹋��Zu�;hL�����fu�m�Zq�#9&"���k� Kn|%N��D���FK[m6�71�P�&�xwbU�ޔ{mF���O3'�#-��m/O21���ob5'���fv^7�3�9}��k�,�,�]�z��Ρz[]��eC݆�&5�į�,G�[�*���t��ͱ!��vU�$
kv��VV�6���P	eЮ(�V��!��Y@;/j&�D�;%ާ"ε:B�-=*I4���D�V�-�̸N1H�y���ۂ�cbua&:�K3u#��ƃջ#�w{k��:^;��G*�w������OL�}�*+т�-��C8m��'b��P�� {�+�.�����Ȯ
�N;��v���ݻ�r�9�nc����	k��I:m��m�q���J� � x8@r�[c��  p�8B�    ��*�@�� ��U 
�   �Q� �`p0��xw�/\��[oY����ooonVx�vu:�z�79�/-��{���v��N箹���ǜn�v��U���y��<֞ù��u�=������q���x�XU3���{��ݍnڶ�稵ɍ���;ݹ�;�]d�ޗ���m۝��8��Ŷ�Nܺ�R�θ�n�۫}�m\w�y�W���w���Gl,���6��ݷwU\ݼp�m޶�������oqצ��/�s����s�������s�G��荦�{U�.zr��w1����닻��������s���癬�}�֯7ۯ�v���ө�V;��i�Ju]��N�]w�ѻ���W��g[��^�qڳ���W��v����޼����6���ӻ��7w^�3��Ϳo߿~�����[Kר��<��l&;ye�뻛Em��$�vs�M(  D��~��|���*�n���9��gA���1�.�x,�R�i��GA�F�݆`�" ǻ�7N�[���2<]������.O0�eU��qFƙzu^Q�\�V����aɍ�=����m�w��&Z�5z����.+Pe,�q:�l��0<�|v���Ҷ/�#v�x˞z_H��bx�z��q�5�'�������;߸����)�nƵZ�Uwe�W���w3��-����lߏD�GbQ#�"qF��8W��wج�圧ס5���<�Ⓚ�Ђd��b͛��H��Q8;�9���\��7�:`ک���ҽ6R�)�˝V���:�z����z��&�d�I�,�Ή�F065�9�3N�p�Y���0xĭ瀡���Qu���cG��_4ju�r\��B뎌C�+��`٠��S*B��I$���6�����C��f2��l��!B@�$� E�Ȟw�Q�⦎X�TwyC@��8��gN��o�]�pڿvT�E�Pc�H�D�*J�#rϽz7d\�78,f�A'�2H�WV��A�`&*����|x[�y���`�*�=]������Ŭ<�WԤ��@��N��q	�>*{���z���-$�`6{Cݝ��T;�fm�ݶk�L�)���QcE�=L�P�i�����z`7mp���cXXz'UGxǆ MF�Y��jfb�ɬ�sT�7���i�M	�/�Z'��/�A�;3�R�Um� ���g� )��X�5�B1_EgN��ږxio���I&Ә�b=�|�H���!�Z0��vԫ5��.
8V�8��-��.�qP~�� �8�!�:0CK��}��U���R�^�]iu�T'?��:�{�ʸ�1CY���4�Mi��ޘp�#ش��T{	83��X�'.��e�h��ٗ=��f������[�b��r_y�����	�^���▷=��6�����W�;.�S�J�+�M��vdm�Ҧh1I:i.�m�K
��L�Ju�[[U�QT�T   ^��W-��u7��H`�P�  �PeJ��6��UG��^� ܋m[o6V=w��޶��ߍ�<=�2��J��wWu�,,��{�2���J'�h�p
�J���*.�g	پ�F/ ͧYŹ�Y<8�v
J�<"� :@H�R}��n2�Un.�c#*�hh�}Ֆbx����:9Q��)v�F|���[�AT[��Ω�[��~vFCG�II��<.���\F�=�s���ňҵdǺ�+n�G���,���-[Ҩ�1�!Sx�U�� $��?Er�2���*�u��JT��[�[	�$��"�!&�it����j�35���c&�RdU"N�7�+,�U�	ԢM<�f�����n�j'���'l�>�&���G4_�3���&�xve8�õ��m�O��e^�f{�jV�CPN�i��Ӥ��E�5g,��q]��茍2a��K@$�)�kP��
�V۽�$(&�I�j�:6�W;R¨�Q��8����י�5Ϛ�Fn�΋ƶ��W6�繸G!<���)x��Í*G�M<�Zr��s��K=~A�>����ł�o:����c��7�[�sf���U�*I$[a�Sm��������P�w{9�umv;���m�9f^�97�o��m^�y�[�u�{zuf�ޝ��v{]w��שmݶ�^6�#�#�����3�oiBi��I�H' }xF�~e?�Wv�X�G{V�������M��w_b��zU�[!=� �D�����l��&L=��b��MI��/a�ƃ��ȋ�7��V�MN���E&h��7k[ y"I��Lq�i�o����[wu�5�t��oz�z�0�a�M���*E��^�Ƀ^L+��+I����mꦽ"��5�J�MJ�t�h�B5($O<	mGxEs&��1�J�ƾ�3�h5;�ѡ�d��4�N�~�{u[Q����Qg�{{�8�x�~L6�H�����7����m���%�m&Ki$�h`�\=�@���\\Y��vv�<5�Q���Mr՘�1�[�y�װ�-A�_hp)*��HI�l���v(�6e
R�X/{ٮ�+�}�Fȁ��F��`b�1z�\��JQ��ʁt.�%6sk*��%PI���Q0��fz�M뻍�7���8��9�"�2��4��y5v*���0�Um9�! ����� ��a��#-��1.5��K@��$�(��p�&��z�w{��z9]=��z�� �@N�ci�۪���0���PGf����lz*���Ѷ7P�)0wr*�sp�a����\����v϶N�'�ҧ��w���רU{EC^�$�a����*�9��r.�H��I6˄��'T�*UX�ݽ���R ��|��GX����Q+���}�}�K�{��ftP.�����Tƚ�a.	$�we���������J��ZR����~}}�þ��4!��Q��^��ZW�jڷ�YA��)�K��xj�F�j:��˪���u��Y�8��,%�����	�ن�=�t	�IBP�(�2`6[d�����RL�-�ï�@�o2咜�\�oPѲI�c}��,��Y��u�UC\��:�;��m�kt����h� �K{b�݊�4�!�-NlmVள�\��׮��[�w̢�gH�n��M02��VWx���n�\��T�L���0�,�m�X��f�]H[-�s���	��HvV�[��t8���n�!vr�p��u�]K�U����tzi������={2�XɄ�g@��.Ƭ27}�N������kdK'�'��[>cje��*b �`�㨷�8��M %�>L���bQ"��vG�<K��tߙ��4g8��'c�#Nh����Ύ�"b�Ƽ&Ƈz�H��E�bc�1�x9��£Z ((DЂ0�2��A�#$��J�]3��&�Œ�7�5[�D�.p 7���+�F&F�Ve�w�Mdn�8�' �C��/&ɲ[i76����T�)r�+�}�RDi�.�t�F�LdT��6�22�5S�SJ�F�B���o
�#��򱜣c�yM(��	���u��w�M赌�9Ѡ�4'6nM�%��w���۹{7#��Um�b�;���ʥ6�ҨP
�   ���n�]Ǎ�A��*�0 
��P\�J� � P+�w
��U�^�;��\�[��[m�v6�o7[m�J��n�<����r���b�cvy�ɥ�_�ٳ�tN�Q�񊕃���h��l�oQ�#���^|6��O(�)�ͭ_���ia�SH��s�blƏ��0����.<]��b�
:��K`ǹ+M���qxtL�rs0C�&�;�5�L\M�Y�%��@&�B�xĎ~V6��O���7b�lt�Tb\GAy�\q��ǘ@�Y�<8Z&7�I���u$��R=�9�yU(�`6R��dؚ�	yHJ����mr����oc[kw)֏����o�j�^�X��1b+���4#�E1ӦU߭>'�l_t$Y�]ӽU�ӥ��E#V'�C�1�6Y�����b�)�3���LTD��*��	�BbĊ�$�-6wt��%��R��.3�+MVi���1}W	Sh�h��f5�*�U*Tm�uM�i��a�������#<�H��1C�ح�m$ g��>��&��]�zXd֐DgmP�pf=���P��N�`����iRW�S�<�:5sޚۣo7����R�wLT��7$(4E���/��DŻ�����T�H��e"�m$����-���ܱ��.��/M��o)�����{�5�z�m^h��^����s&�m�zZ���U׻{��]�s�s����z��V��K�����B.
�4� 
���ww��J�Mh7f'���P�Y���9v��`/6ǣ0�����]U���+z�a�QN��^<��t1<i��ę�7���F����a��a��qs\��6�3�:i�UA�4̙{2�l�e7}g��.qS��l���&� �3�0�p�!��p�č����8��<�k�T�8H��V����ֶ�E�&66��AP[�# U
�BF�I	���ю4+�t8˳"��n'+v��Et9�r���F_�$���T�(	�:!l�\d�C�U�v��#�n�g��%sh��n�
��^�\��@*�U]�挔�O@��8�[�t�O$R�����ͷ�>�0�.�^^t�[�k���}�y�����T
{V-���j.E���A`��+�<��?%����c71�9@	P��� �sY�sڢ�q����׽c-?p�������q���@*m��Uqwj��$��c��<8A�bt}�j�6�n�B*�ǭ5ɔ*-�m���30�c�^k$L`}��0u��v�H�OQ7���5G`A(�m����s��c*P��޲��׳��݂�Z���R�s1���[��­�Vԍgt��ɘ'aw�Pb
���4��orp�6F�1CX��D��)���亩{��FF��j�N��&Vt����D�B��!�;�Y���#lOg��I�H�\;�o2�"@$��0[%6���ǫ*ثlV����z���i���Ux���3��H5��j1�rDX�P��bF�Q�7��i�e<Oe�^�:	�U�Wd�!~�&̩Jm��j�1ƔX������������ꆘ#aϼ��^n�;�PB]�;�d�
V��>Q�'oԒpH��3�a� 4f�X�8���{1k�`�+-^p&c�K|���MяQ�<&|%�ã��O�=�kz�(��l�F�[<�P��-	
F��(�I�0���D!�v�<�����@]���*�p�?$�H�1��et <a���l��dz�$-d����U�J�����z�����H��}$wy9��ٝ�$0S$�����4� �~���ꃳ���.0M�'�.	�9���(L(7�E[FPs��	�w��@jn���$���m2]�on��+�E[�%0�I$�H����-B)��)��B�*��Jϼ���G��N��HH�m��]��e<�+~�َgflkQ)���g����F�X���s^z �"��&R�N�d���6
gc��"vL�^�)���4�e{h�+<��PLX�H@"`َ�^)�R�M��7��E7�fA�żc��9����He]��7%	�E��A��>(Hv�eqq�>d�=&�$N�]���^�n�e]�mO�'�T��B[�^���m����g(��b�b��(w�V�YÌ�S{l�%��(��D�x��vd7�cH���h�"����Ɏ8)��NЭ�}�����4$`�;|V6�Jd�Ԇ{�`�q�����xF�5���"s^���T�.�����yF���wo��f(��㙭��K&��;M��,�PI����^Čⲳ9a��ܮ�C����d�|�V��z/oWZYa��H�8SJ�����˒�Ln]�^�n��W���	+/�y�����&ni�Aw�;z��S
�G�ހ�b�ު�E6�(U-�j,.���YB\�YT� /X�7^�)V��� n�:�ˋοؖ��7N��+�)��G;�����92�/�3�It�������0��"2����N�œٴ��n��|(�U�
�0Fɻv�m��m��m� x�}�]ݽ׻��{Y�b�ֽ���qT 2�k��� S�e6  �wl>[j��6�U@UP U@mݫ�ol
��  ^�[&�|�P n  ���  -�_Se��@  
̦�Uw   �  �  
�                 �g�ݽm^�{���v�oomn��I.-��6l���n�����ٞ�2�%�oV�;�g{�*n�   �  �h    6�  +(  �   @ *�[   �EP@    6z*�l�@ *T� m��*�   �    @        Y@   Y��  �   T��  <  T �PU
����� N�*=Pl;�յ  |5���¥F��z��
�����T��P�����AI�Cd�%QT{e˷ U���V�P   n��ז�z�;��zն]�a���T �U VJ�T� *�^��*���[fRٸ�wQ�K�[C���N�wsR��� V���2�P	A���<;Ni�:�p��L���r<����i��b��	���;�UP�;!G��<��Am�1�1���X:	��!��d���=�=�m��J=����F�,�mʄ3/�S2.-D�U��&��������A�zI�#�$ٳiSI���`YHq�&�H��V�=1Û��J�C��lģ�ڦ�(�=��zx�F;eh9���M�+?[�;�����	�Px)+3�*(L��@$MQl6R@���X
�����oP���1��Q����X�ݬ_'#��}1��8w��"���i�t'͞}Y;�ӆ�oT60q�h��o xUZׇBq�N�(h�'�lo�rQ(��W62~Gak�t6yE��V�߽��|SBb���W�,�B$i -�M�z��+��6�R���CH��E�1q�{��q`�A��q����^6C���tE�#�~�������G�k����\�1u��F��Ǭ� ��Bs��1U��%��?y�D��u�D,¡P�PY�>���_���ڥ�ӻz ������j�����m�ݼ��{����˚�woovz{2�ou��=��̩��w������ۧ�o��7k��w����wם�u���w��ݽ������;{s��Ƞ�&˾,�����G����lH��,�jf�$�\tb�Q[ O��b�5+��m�I��iTPݵ�j��*�Ȍ+�{B�z�N�V��@�ܺ'���RNy)#Nӻ��IM��>�6|5�Ǥm�ioW�m�[u�w��nw�Y�tכ&��'hCH<6���Zh������m�1J�P˥��zX�:w�x�$��oZ��ZE��	�fc{Z��ޥ��:�)9�L�1U�_U��LR��Qxc�m��pS��D�\2ͳGp~��АmO#%'J�Y�e�Z�[��ݷ�ɒ���X��d�)�JL"l���hVL�[�-�t�P�D)�t�H�\�W�D��\Wd�9c����:$.j�M��9S	-V�M$��#�$t��v�}3W�8h�h���'�Y�C�'IQ�����e��ǏC)<�J{�C�ʷ�~�I�I�Hbz�@]���"�xo*dP�����1�I�5*~Q!�~I[�sacv�̭����qT�4%���~pL��;���*���
y���c���ҵrD2�b��~_|Oj]�e�kh�v~&s�H�ۆ�PЄ˿W�\��\�wP��f�1�do��"X��,%V�Dx����Btdǆ].|��Z[D AR�ט�1]��~� d<>=C�Y�#�SX�riu.�Gx�Lߒ���n�L��y�;�+� �Q�2 `�u���{������U��f��P;�
��u�Y��a���������\���80V�8�b;W\M!¯ۨy]�1P�~u�I�eP����j�ffQ�i$&;"�����-.�Y1��(}�ܹ�݋��jĞ�5b�lZD�Y��H�$�(8Otuf������up7��`'|�N�'�;5����g�%R��" ��n���R�h&Z���p�|�1X{��@�� v��oK�{}��<�ݯ5٫�?��o��0�w�rt��gN�3CE1����{0~��%�1-���uԄ��a����W�r�v������ȶ���4ckb�&%�S`���1����4�x ���#�V�#��<u�V��4)'OI�9n���Id��#Q�^5~�
$�A$Jl��dZUm�\�]ۢ\Wu�LMw�ɦ���7R�dhzJ�5&G������p�)A��1\2c;<Bk#5-,�D�X��O�3ʆƒ��Bf�|3Q��G�Q��@�E�r�Io�k�S<8��M���5:��A����zn3�GB@L�\U`x��KU�����7^W܆�Y�psNI���#��Y�/=�È�p��
��8���nusL�wc@8Ov$�Đ6A�M%�$�T�_qVk�;��;�9�	ʯqzw#�u�u�����xs���Dئj�&g �!���!�EkZ�O�\�x
�wà��Ic�8�-�I`2RI&f��ph�HG~d�̖�<H�(�E����-��*'���N��Z�|g Ӯ5s1��f�� n�|�j����h�+I��fZ<�
���۠Ѫ-����T�*��jnoc �p
�P�   ��w��Ǯ:�=|�P��*�ڨT� `*��� @QT x +�Ql��r^�uN����`�+%Sc)T%�Ca2m���	�6]s���k��yTlJ�x��^�x#Y4 0���j�c{��u?vs�i�]�ҲO9ậ2HVSD�\pP<#η�9���:��`��ց`�:a�WHDDJ�n��'��o��4b��gj1c�(��,�L�ʎe�iU]�rj�0`��/|~���t�}�`�� "��u�ؼ�H�����9G���w�#�T�:��qb9Z��$���(��T��Ld�L	q��Ѽ�Tt��c;�8�9;���V�4E�S�#@�ck*4��d���x�e��d�H��#���+ i7�j~����RJ{9�V�=bq��h4(�{G�z�p4���P�b�jl���_�����V��wP�w�l���m��I$@P` Yd2�jr���y��Z�p�-"�é�]��ȍV��]���7E�̛2x�R���A^ĉ�$p�=~�(�S)���j��Q��,��z2���2�����y�q�f��b(~�z^N[{�w�+��W��۫���]zخ��m�c���3���w3��Nwz�w�ܷ�:�����z�N^�^�=�%��\����w��{v���]����y��^�����z�s��re���y{%��P����檀�oZ�e[��;���&b���'{�o�G�>1Յ�,�'ZL���F�!������WCp�4�`C$E[��C�-*�]6���񥷜���'�ۃ@��)Jh��w�pW3tE/��i�����H���!\ ./)j&zz$LU-���\���%�b��Y[��IS���E7: ���7�<���&y�(�r!r^�o��&�@�GL�r���i�}�U܏Lp�88�s5�Y��ЂM��Lx�;��	� f��o�u��mM�}wewm��m�� �!�PM�<�˕��= ����4AQ��#�Χ4S��7�1h��k���4�;�a*���5�Lb>�,I�@)h�b�P���F���xH���!i���V�q&<��'a-$+3�=��m������Zo���4�[W��tH��f"A$�!]e��q8ł4\�d���]�G�/�z㩳��
V�3>=F��*7����ngc�Z���>�Q�<Y[;|�׷�B�e�r@�*�(�-���s�ݚ�Iin�AE�I�0H,�Z6M��O[�*8�:"7�I���1��p�权ek���;�ᰐ'>�R�%a��-��IBN�W���O@��{.�:͓w}�	�԰B)J�j9F=o�0>=cw�0��:"��ǵ:�i&�I$�%��Nj�*�@m�.���2����9����0��K��י4����j|�kn�a���< Y�6ĸc wF����&�ݤ[m�J�8}=D�hf�>1�n�-�'x��k�$@�6L��Q&�hݳ��yyW;��E��d��cw7qt�.�M��z�u���S�c�orx�%_F޸e�nOm�ڿ<�Ir�i �F6�]sm ���(a�0YP�@�\7���;�\��R�S�v��S� 0��5��t�S��Q���k�j������;b��B�J��x$�x����B��I��V@�3~�yǺQ��N��-:�0�U�"���L^����@xn
$)�'�䓅1��6��NLƒ�F@$��l��3���� m����X\Ǥ@�/��5��&�LP�}���MP<��Z����FI�Fh��.��#K���8D'&q|ƃ&P�h�Y%4������r����;r�+/ze����@�?�>�J����F��&�	��r��vDQ��k��#Z%��	��n}��(��7\���������O4S����)�B��ry���q�', zl��/٠q��rI �f��R7f=J6����,zt� ���2�H�e>Z�Xԏ�0�����������jC�Y����̴n6*-F��d5	RG�;t,^6�p�Ev�":F�!�h\ً�囕.r������t,I��^�L�����B�4ҺǺ�T�ot<8L��I����⽜8ej���}7gv��5���̬���j�`�];����y@�����o3l���,�@*�   Z�����ޗ۷�C�dP��6�
�6�T� �` �����W�?f�튪�qݸ���^�߶���S`�󺨪�m �e�I�Z-����~m� ������5F?_j%�<��<`z[��EL�t�{�<�}\��������UŽu|��H�eg�K���4�p��%�IẠr��W��Ӯ�qK��#4�èr���BI�җ]��~(����rX��L_ <7ǳ͹
�f-}��n�a�mųV�a�f��l��G�3'9s�W����.b����k xn��D��U��H��hm� f���\��۔ݽ^v�IA�H�=1BA��/)nx�cv��ݎA��_d��ٽ~��Ezw}�`��扱*�U<g�	&!�b�EWs�Fi�0���f:�@�S�X�Bw�Z1ct��NqkN���IOa�Fީt�Hh�t�A	�Km� ض)Q�|�ޝP79j��k�0��p�	�J2��(�ܾ��9���T��.���s�}$�-�7J�U6I%	���]h�� DԜ�X��<wU�xQmLw���w��v�V؉�p����m*����P m�Usx{��������:��h2�m� #d�aCP�B�4��c�U����v�g��U{�o����[�\�9ڔۅ^gZ;�è��Uu��׋�9�k�;Vq߃�q�Ic9~�O}���&w[��:�a:�QI��]g�v�ڪP�ɔ�E��z�k�㑣
��U��6U����l@���k�]��	�q{`�-���w��}tHl������2{3%$I Q�A�"I��D�8�w���]z�&��qvF�����$Fa� ���Bׯۅ�)�l�w�)ʘX�$�IѸ�ń 2x�fwH���4X�k<7ڰ#F��H�:ЙW�_]�3�����KtߒJ�K��;�[[ڿ�ν�d�q��m��H�A�d�a�O*������˅��%}�3�x�!�{��F��A	��ü��
$�$�h���@��(������f��I��tv.�>0�uI;B.�
�	6���-�V �H�Qf���A��ݚ�cE��`;LO�UQ��7N��'��{z��l;��p?S��,����ëTέ7U/�Ϋڽ%�J��jΊ�G\v�2���̻��U�� c)<����Y�.�w/�-�5�1���0��h�Vˬw[�\�3��e\��l֭˷����o8S����o��k�v����w�Z�+�Yc6��{��ɪ2�tT�tm�{��s�:œ3sOT�CR��%GS&����V��se���V�V�`Ĉ]�ul���.��BAf�n�^\�I��癵����rP�cjs�$\B�#]������o�޲]�(�/]u^P���'T�;�*���׿5�������U����� � ���\�5zwz��\�  	� *�8@  ���K^��  ��8P     v綢�z� <�@]��Z��؏^}]n���ﻷ;�ܪ������[�ڬ���M�����/�u���:�*��n����w<���b�s�<�������!ɫ��sM��5�k[n0�����Of���ǳ]��w�r��/[��;y��7}s�m�o:�����<v�Hی�ۭ㗦���5�V�n�����Ty���7V��^�mE�㵬zw��ǳL�{�K�ww;�jw���R���*�K^��^�u_7yj�{��~�ھgn�/{{S��ܪ����f��ݶ�wZ�]ǹ=�{��n�q�c��m�y�{v���{Ov���^���v�^˶��^]V�v��鵫����hŦ;���غS�]�{vS��f���g��ݷ��4{�:N�dӋwS[��KN��S��ljV�Z��)�n�wsG'n�k>�b�m��Z���%��ϵ؋��{���ν�l���8���zh{��{4u�BE�1!d]���e�&�l�~�$���݀+h� �
!�b0RMҀ`&	,��!^�8����K��E9��8P9:Ť�t�z����1�q�'Dp��"�ZJ M������cC�Ƚ�/|2�`2|�&�^�v��ۭ1����NF'F7L`���G@�	M�{U��{�b��9p�CE2JL�	ު*��@*�z��lYE�H6��TL����6Y�Ɂ��L(���cĮ��Dnӕ�T��5��:�͌	A|�(w[�)9���O��&rn�[l����*���_�w����87��|��:�{J[�q�eo[qq���X�1��}�a�l��E�d�pJ����Լ���L`���7��xc��;������o��m�e���i;�'�5j����M���l��������ܱ�J�+�4���R�;�"̌��b�c�'���݈������t��M��4s'+�u��i^����vˑd�59>��%$�l�";�T��L��SVO�jS�1ō���q�5����l���ǧx�s[ш�&�)Qb�Ḧ�?����[�j��_F�:��P��~������:�h������#���<�� �+�?5;��%��8۩ph�ե�*c�LyѨ�����Ko=��
%�%NK�`m[xm��$��X�F;�����
���n���רA*.�\ ֕�%�u�ݞ��+6���)7�m�PT; *m�ZdV���j9������w"�q'	�狅�l�n;�%�<��7E������[�'��WLP�%w��]�-��N�u���>����rjj �����t�_���홢2%D����Y��.$ pJxK�0s���ޒx7���-m��h�Rs�t)R�m�B.c<$9s��;��ī^�:����A���]���U�
;4�H�K|�o;��<$����T�+G/�`�')i�!�݇x�깖ޫΗ���$B$
T)&`��݊���.����*�ez�.P   z�%��d��=ݶ��l6���Pm��@[j� ���z�e U�*�?�����W[��y�Kewl�U]�ٵ��۹ �I4�@"Hj:��ѓH�~��O�p1�0�Շ���m��۔��j�=x�k�7聤�6��q	���^�V[�u m��!���6���"�cy�� �\���n���n������~�D�.�C�i�\:+޸���P����D��e��G�^��&�=q�B�Q/P�jRB�F���7ѡW�=�IS��z ��1p�x:�>E��)���m��4�����M��ך\�7�w��r�R��n`A�VkQ�����M�(�1"��(h�{��L��u���H������!��gm�l l$�>��zL(����'#��vk��<�y�8Վ��d==^'��k2}´\��! S��ɮ6�nN�p	8�"����w(��m �+�st�A��2j�{�8!���i{�\�z���Ei������C�Mŋu���T���ۡ�YH@M�뽞��y��j��=s�ni��>�WHE�d��������Z�?�۵J�;��Wׂ�@6(��ܻ[w/m��_�v��߽]�o{V�]�Ӵs��u�swoUw{>��;7�n��5�>����{�z����:����8;�ͫy���,�	��`��-����%?д!��Џ����5�j�i4��P=A'u ���^7kv�(Kν���χ�T[�K���緄c$��p�ΉA�a8������w�^�0Q�X{�f�����mK,��8¼�(6���@$o7�e�,��a(,�C �/� �I`���h�IS���t`�����!�}�=V�o�4TG+P�{K������Mf(�F�ʓC%(GE�,|�q���.�Ң���cz9�����z���Xu	�ԇCa����ݽ�ED����6����T�QRP�q��3dE��;Ԓ�'����02ZZ~�5eh�47Ðs�W�=Xc����Ed��oA)4� �7��u>dIL��D��n =|�@�9�Θ1 bRcI��
#Xq��{O����w�sS%7
��}��.>nr���JI������`|Ũ�r,.��<��¨=Od������mLd�ww���{]ݣoswI��wXݯVgĎr���Z�fGW��� T���:��b4ҦKh�,N�@z�kx��E|P�I  %g�0à�D2�S-��ˉ�I�3wN���0p��������T�jlyh���3u�@���s�~˼p�&m��jdm����-
�FF��/ۚ"�(ֈ��՚6\�3^'x\dtg�I+�;���6�I �@P��֛ w  ��w�6���,�ܯu�1����Ŏ���"���=���ɠc���J0��`��Ⱦ��H�7��*&��$���$آa�W.b�H�- xmMCj��Msm�܉���6~)i�O1�d^�v�OB9+3��a�	X�M�BI��b ��}[ȯO��QB����u�����z+�޸�]�0���7��i�-)\�9��tS��2/� p�I0�b�,��i6 Ł��
/-�֪���G^�����~��v�7�Qa��*�����t@��<�>"�$�*�#�GP�-���X�m�O�F:X0f�Wl�@�Q	;�����}f�$�؞*Z����������'2�Ss/M�^�ҏ�X��|hw������8��p��X���.�S%��m$��������Uml�[X�! X-$�-�Y�P1٨�3v|��"*�M̳y����1^<4���S���[��w�mj:q���]h��	�*�V�B�m����k0ׄAb��h���A�-��4�7�Qa��1I*��մ.TX!��b��VF�D�����q�}:��D��Jc0������Q�P�+`3�Yw�-U����Z7q{-�(Of(���^5�x&��lu��^�y�n�H
�e�DƆ�O��0h�V��E�P�L��A0	�.e%��͈]�sZ�3+hi����2ǐz<'A�Mug�@�1@i�L�w�<�Ǿ�+�$�.�Nׄ�d�X��aZ&N�8P�p��T��Ր��Ϯѫ#�dA#{Ψ��n\�CA�:vZ+�� ��,2wsX���+���*�xJfykw7U�u�;F��*h���]vݶ�� E$��7��f� ["�mM��5P[iU�U   =��ֳc��w��
���T � m�T;���*�Q� q�l�˺����vw~�,������eT;�R������%��f:�p�6zGA@VV8�(p6E �I݂k٘�[���aY0?�Y�&�@�Ȟ�]���z}y����J����`��$�c�ʉ�)� _r�m���GuYB����vr*�Mlf%P�.��ت��7)2Zh�NZG����ގ�0N��R����ٽ�c֦t��c�ϓ��.P�F�,�����q͒ibFPD�I�{\]�Ɣn�{�W����ݷ�ӽk+�{d�j���SZ�0㪲��
�6f�{P����*�4/6m�*$9�����)��&�l�y�Z jBčE�;�9���b��,���F�!���bm���G	)\�:�U���D Z2��wm��tw4�� $��PM��%$�,��ďq����'����y��0<5� �ud��͎OI�ʚ.�C`^����D�(�X�9:X1��)$% ���748���b\��_}��$���j��}w��0��%��M%��xT�mV
b���z������S[�v�� k�^� ��{���y��<[�n��ؿf�m�:�c-�;�=՞+��{t��5.����q�V��v��yMi�����)݆�<W��\�7

�x��t�
DX�t�*Ŕ���E��]E���Oo�Q7���^xH$�n�'Fd�B{N�DgL5�r^�_f�
S>%p�#弯[�������Ҕpn�,��m�c+�[1P \���
��{���޹zm<��f��M���EuF��Z����N:��腃\y��_��w$�we-M��"��T\�ǃ��RH��T0E��=]�2�;ų�qO�O)��[�9˶�hۏ	9 �ZŕSy�A�!:3z�,��+ƫz�o绿Ϳ��\5�[CR��Um�J�[7u��UI~�?�}�>�y��hp�70p}�嵡�'p��~t�@�~�Y���4<V�SI!��iA&u$���A$IZt�e7}ո�+��N�b�Y���D��؊ۭ�J(
}I�ʹN�T.�i����S�+��.N����0���QI �fz��RB�Q��.�Ri���Ӣ��G\�V����j�T'��c`e�c���Z嫋�n�g�}/������w�Gt
�	�J����䇩}=��kJv5��Z*V��N���S��!��՛s���L��{$�P�ݾJ1~�#��\=� 8)s�!$����~BoZ�O�L��D�� ��<�����u�-�5<�mŒh��y�Vx��N��9��CR3�{	��zL�ns	��/\��nㅲʨ�#�-!�t��u(�b�U$�,�2�6�B-i�Y���8��J�����m#��E���s�<��˙+)m����6�U�-���ф&�� �5��Y���đC<�Q��Hg{�G�3�����<�����rQ2d�x��J������Ȩ	�؋Jm��`=���I!��Lm�5Q���o��Qj�x�pr4!�b��֢���`��SAI~#N	�Zr������f����z�z|e��Q�T�5�kz�q����aD�̾�`��6>#t�F�.3Ň�;�΋X,>��|0��_�a����)�W�7�r^^��݁>��k�70���kbI^48UZJ�u	6�
sM��.��&xA���7�w}�;�.*Vt�.����^�h]�����^�FW�*!���o'-�Mc��%%�U�A�cd� D�"�i�Ii$c,X�n6�����+���G�UW�qh�Т�t�LqX�שp�����gI���=����N$�4V�Uw|��"R Q�J��Z�.s���Un��Y�cx�(�p���Pb�����;�c�����%�qinHL�H��װ�	�1QZiR`���{r0۰������h�ʅl�os�ʂMJ��g,� -��g���"�p�3�n�E4� �K`�[B(��0�'�0�M;��Ĺ����X �#@�\1������ �q�;`un"���.��`��Ӝ�ZU�n�$�YL�z>sׇ���O�o��*Ď�ϲ�3�t%�T"������� t%oTq� J&3�9;�1p O�=��IR�p7e����-�A�5@�Z�fQ|���#]�)u�nv彮�e�Ne]��К5�n�k��(6�9��ܗ];����2��a�x�����HF�;m�;	�����rчb�#Fd-Y��t���Ț��wwư�q�vH�+�V�W]0�.�WؙF^�:Z�qѕ���I�=ׯs9��8��ڻ��T����[��7x���U�Z��jcU�*u�^%��
��:��6���ub�8�O�oT��݉F�Ecr��ӽk.��GW��$�7@CƮb�\��=�{����b�+��b�:��   �N�N��巗��=��^����� � 
��wjm��P �mQ� *�;�;v\�� U    PP2�6�Tm� *�b�گw�@ {l j *�m�+kj�� mN%�(      T  @                 �^뽈坶����y������:�]��oҭ���ޭwk#�u�m=ӻ�غ��e��w��2���r    �   s    �   �       �B� m� ��     U [l߹߿_��   �   � �  /T    +(        [j   Vڂ�0W
�� R���d    Cl :�ll��Wv���N ��ٲ�  u����x����vq�����^���[v��b�*����~��
�6̮�z��k�b��@   .�wg����N}���z�6�����ꢨ U   x *���  ت�p���=�K���;3�U�mo5��v�b�E������`qRe�����\5�@��75Il�˴bIA'L{M���<�- 7��K���^*�p�4`�hF��Ilʉea"��p����ş]�pzb��[��1B9�����F�?�K��7&�q��
�z��F$:�$�m��A֕�81�t�A��@�+�E,���{5O�����4o[� ����*&3����I���-Ht�ZF��bk�H��F��;��d��_w�w����������w�V�/ �X�G���srXS�y/jxp��������s�Y��E%��U��ǂ�� �j� ��.�i�ɪm���Pb+�zG�t5��[??i]���v|�N ��-�T銳&������4Csp26UV��gvE�0@hm�ޮn� 62�FۆKHY!�������W�dr�95�,j�`sq1�Ev�)�0,Fg�[�E7�]@t"��a���Z���q �eU�6�GQ�(�LL1���5<�~�CPa�n�ÇO-#�K(��}1]�ޖ[J�I4n�� ��=�T�q���W�{r�w=��ٺ���N}���T��˷z���z��O;�y>t�>r۝ӷ���n����ݻ�����|�۽ޟ�A/���d$��'�Fa�jOG#�����f���ng��3�Ayn'�;�j&������^�ݮ"�x^&V�m���`MY\u�S<xC��#����}��:�l>ڳP����Ѯ��ItUfh�N�!�$f���ȷ��f�J��=�Y�2�T_�+֩�k;k�w3���L�U�$�f�� J^i��1F7��j�� ��:a��VK��S��W�#E���6r���"�-
7��� �gy�Q��1��t�u\���T�(�#
\�D�� �u�s����3x��M�V�#�z�M�T�VLQG6�6��.�*� m$IA  �i��I�v�Б�T�h]CC����&hps�8�4�H�h$��O�=��;�"o�%5~���:���BQus=v!��Ia�z��43�9�:���Q�:5��`�1F'�P��9����&��#�wT7�l��L��$�,�'��v+|S�Kĕ�$q����W�3��#�zl�QRQ.�p�B^J�*L�:PJ}j:�A#X���ݍH4� 7
mo��+-6�62�c�����sh� �h�D&i!M*L'	�j[~��-���F��#9+�!&'L]y"nctZT�9�RG�������v�ps��I�ґ &�J&��F;��L��ݒ*�p�>��&�7�!^ ���D(�}'��r[��1���S8����T�'`�6w������c`z���
��h�{zs�kب۝��]�����799&�o�sX�t��z�9�b�Ǽ�&q�ȓ��دc�DtQ��Sxj;-G��R�ibD2�QQ#�⤧���z�F�V��R<���~h���Ç�,,�/�W��j�tz-���/X���T�G+�Z��I4��Ɖ�>�ژE8,ia H��Kb�P�[��o�p���AL
�!֘�Md4'���g8w׷4��FL�G i"Ӯ�H쬻���
�AL�i�C �H|���I!%"Y�a5�,�����En��s}�T��(��ld]q��X��A�`���5# Gv�Eu_�����Hn�FY.���/��287K�E��-��}�
M�a�"I �1.��Q�@�F���D���v6�<����Ǽ6�kLy[(ž'^d.�j��.V�ǽ%!b���OPT(J4��{f�7y�� m��KM��E�Ii'2;��(�Ĳ�ҋV�\r�s{�^��+���2P��ĵ,BS����w�:uzpB9Y�9R-� >�[��F�D�a�X����y��r�şz�l�Qva���?p��򞢦Fo(�<n��U/k|���W���c.=y�=�É�4�$E�c��`���`�� ?y)�~�&���@z���G���2�O�W}D�g�=��	��e
ˊ�dxQ5�$�B�ð^hI1@ `P�ʠS����Z	jqO��T�TǞ���%�u������\)gA���\�c���Eu�rC�:Tq�@ƽ�E�h��T!g�l݆��¤��Y��ۻ��Y� zΎ�3u+�V� Q��Խ�ޔ�u�:Pې�E顡e�:ͯ��8���t�LéE]��4��>K�)*-�-�YE�����2.��+\U���f���   ���b���n)��al��m� U*���  �EP+� US�{��m���W�ݿMot���z�+�+�;{���� �UU][o$�I$�w��c��Ƥ���3�E}:H����E��-ڎ7�tI��w,P2���W)ǭl�o�Y-o��l��G����������{�g��hP��8Z���N/L!X`�c�_���_�:���B��a�5r�e6�-��	�{~U���xX04�'t+�y�C�@�>C��NR}"/�ؚ��r��y'��q��6[�>��n��Z �I$�rŝ�P�� ����T�wgoO���Vou�Ԝ%lV^d��߁��EVہg!Ā3�t�d�i!Ԕh�vd{��yݿw@�7q�B7�?+��	D�4�����_��"u:O�5*�\zb����9��*�ܫu��鮲�]�ŗ���4��ܑ���L,+ix�i$)�����
���7
�q��CI$1���K꣧n���=��Q�.�#*��m�ā�����k�췝�q�x$���Q�f}Y� "`!6=G�vsJS�7���Ռe���MX~R��\Q��ͲĢeM��U��w }�6�@:��zז�w.�o/�����������e]����znz�m�{�������z�e�.^��n/�;�{��G��g{/�����<���Y���A%A?�G��4��'��Bէ�y�w-	\Tx�T��ў�]W|�xn�n�@8�
di�IRR1Qk�������Щ鞡U=D�Q�����3�*�=]�E
�а��������71"4�Vޚ�k-l�=�Xp� D�1�E.�*��zr� (�Q��$B�t�&(�U4@��t�9����KF��ˡ
�����������7�L��S7�i����%�]K�m��ob��F/�?]R��A6kq*;�hK�8���r���H����%�݀�&�CEp�"m�?�1��!#TwSM�{̩�7( -&�	2Km��y}H�U-��Z*���tc�6���w�r��]#k��dj�Y'�^�e/I�\pN�q	۟��֦M��,�J�j�C&�G��VԻ�؃/�b�gj��������l5�*��Uv�hת��p;��Ɠj�rgwOA��i�`j(�O=�ĭL�3?s �����X���9K�vW�{c�]#Ǟ�T�C�x6o/m5>�uQ$eQ>���P��E<������2D<��vwC$Vǲ`�l{�2vT^x�d++>%٬��xP�(L�(��E&�*D6T�Czû��2��#Ԑ`���z?r�9��u��sQYC�!b	�a,�q��8�{�A�ͬ��a�e��i��b@&�)���� ���	���;�)G/q�|�6�%Ζ�Z@_s�
	�N�(l�D��콡w�G|���E�߮|o(:E�I�J��yM�8�
��������aڋ&�8�n(��j���$ �����;��&��n8����Hޑ��� #�v��J/�ކ�{ct�a��W� 0&:-些�*�%5U  i_0.���0i�����$�%�$m4��H�k��$ "�*2�_5�*��1й$��$�^y10Ц��I$�R˪@�n7�;��04+c��� .*�w�2\���:�#Ó�� �3���֏?���A��*�{�I�{1G� �nHDX&Z$�3|�2%\G��*p��t��` ���f^�a���u��?Ͽo� aS v��xN�ڂ$�@0{��g�k�޵4�lFq���~��86q5gq���F����zz�l˪쁑�$��|>�"
ޕ�h4�l�JD'7����@�vˀ#:�ȖՉ$E�" ��W=�@�"i(��",|z��%�G:�?���S70ڮ����	mu������[V�����<��6$������ڛ�^�ֶ��P�	�H��M�Hld`�fKSD�S�\%�m�P�����@H�8 Y?-T��9�2��v��j���qB�iå�Ө�F1 v�{u-Z�d��J*��h�>T(� s?t˞���&
�ޥf��Iq��>d���~&"�x>��,�I{�F���P� ��ə��C[)�����g��Ԁd�⮢���RM���R�D|E����ǒ�P6�EB8���Sm�}��b|�+�[�� k�_U�& d�#�G�5��s{�gA	:�Q�n/��#�ⅿ�:�o�R!��Ȁ# |D<5W7�Ò ���i���{��aܫm��ۄ��&#e�	�\b�D�<�ɱrc7[��,u��T%|ტW�D���ܵ�܁u��	Ȑ�Z�R1D6�S'�@���FD� ������"���Ԭ�����d.#k���8DH��~�b,F�&5,qLK?n�-(}����:����f.")�Uc����ԡ�qҝk-�7�^�)��A�m��$GĢJ���*e�n��m��n �cU�B�l�   �_wlmכ�u�`6�Ta� 
�� ;�� �U*��UT�G��wVSl;��3��|���t�m�m.�mU��UJ��w���i"������j������
#�0G�au�\�3Tu���Q�T�|�=1Sy]�8������ Guq�;[��<@��5��<�|u}����<��ЈCtŋD�p}%o\��%��c�dm;g���E_�\V(�}Vd@"=��}��1u�р�n"/��k+�f/��$��Kl�s��>T�8}��W�G/�~^�VÉ�" �&A�!��6�ֶGTh�*�wr#�£�ZK���
s �"�(���h[(��jb7O�0w�f/�A �CPH�Q)(,�A��N+���nP�V,cD��:LwL�>aEi�b4D%�>�R���f��B$Ae����=�.���T1?H2o����g
֤I�p����}�O)E��1]��1yM���🾑�gB��'��c�������}9�c����?X�𛻞ӎ�#<�[�����!�d��0��l��Ul�^���e�����=|�f��zϟ,?V|a�iDb?`�rӼt��yZĢ
��H�sj,���"0z�p�1�b�ƒ��B�1�A� �K��
_���nSZ�Z�sE��śͦ��x�no]��������'�Xjչ�n�]z�uh�'�ܷY���<�޳�-^}��v׫���[U���x���糪%��q����fV���^��{�Z&9�;���|��v��؎��g^�|���	?�PAկD ٍ���0P��X���ݸ<��"$V�����f=�̈́P-�F c���"2}nQh$�F`L|��`U�N��g���X��;�6�_!S&T�Ⴧ��B;��^/j<�n��e��p�P�,RH�+m$L��d�qi��H��I@ �(2Z, I,��B/�|#�h�1���ᆎ�� `3����Mi�8v��{�~}��jW�KЯކ���e$�,�1�y(�/?!uP{�݇��ācDtN����b���Mc��5�����f�E��{�WBQ�I $�&Km���J��@*�۳����t���s�� } f%"խ�[E���`I!�US��$_%�Ę2w�\�>�n��E�����S�b;�1���b����M �`2�]�<�Um�B{[s�%�r7s������|��Yn"���Y��VqP��u�4���_q�Oc`劲�U����i�I^`�m�3�>�R1�n����F��d�����Ƒb��C~�g�2�᭩u)���܉�T�*.���q=�^3�V�ʟ�)G3�U]��T#)l�	xO:�߹3y/1��x�L9D崜⓽��+�y��;��a�wȷ����ة���N4	�os�v���2V�(t/Q1�u���c(����x�u��h�3a"���m�Zt.z��of"�1/���8 �kp��YX����f����CEU�вgLl[����m^edQq0��8�N)F����|�1� k�w�h]�"�jv����M7g*[��P���Y�y[���6�Y�q۔�ԍ���S�Cn�dd�u�������󿭷����W� ` �zxP ��f} �^����M�  �     8Ow���'�  ]V��    U�n2 U` < �׃�7�K=r���2��S��w�nw��N��.��ɻz�ˮ��^�i��[�uV������m�ώ{���Kݥ�W�r)�ɯm�-��W=<v���s���r���l�qr�F��ni�ۻ'<�v�����z���Z4㻒����l����wp��w|��;o{os����L^�����m��^��7�w��ny���/on]�ݷy���u�����u���������#im�6*�n�ږ��]֜{v�7�nkOI����n8�J��{w7wj�1��7׼>��{�N�]׷��u�;��>��}�smk�����s��Y���yݓ��}��v�Yy�s�۵���z�KR�;��k�ݛ2������^��9襷ӭ9ϫm��[,u;Wi��x��v���]ƨ�v�W7v�;��n�i�޺����ŵm�=�T^�t^q���g�'/�P�C��m��N�0�s�4/��P�ue��i(U�VbL���'�P��m�(!�	����4�p�`�}��t��G[&��_I2�I����/��ET�1;�M'=zN�ʕQ;��-slz��*@Z[I6���qT|�^��Q`I�o�H�Ǧ�نi0j��آbG�r�|�Вse�Zl4�6a�@��$�-�[%6�����Y�Gu��[efo>�Oïӛ@K<r$Ų�VM��u�EY�z��!t�COZ��M�Ț
׹�!��.��*�n�Z(�I��M+
���M���ߺ+�]��Q}�X�c����$U�s���ƛ�K�K����v^{�|��Y4|3��M�Sw�ȧ�p��G�<�#HƧc'�;/�U|"|�^lأF_h�/ç��`�ލ/w�H���!� ��M�"6a��Z�_�2b��uHh `�` �2�h��L\¼�r��-�Yƴ��۪��< ����x�9��ET(v^����?Fj|�
�)�rF����xZ�b�T݁~w�˗~Y��6N�|hg��ֵ��@ԑH:��i�9'�2gF\\"��A�'�����U��&�k _���6�3LXv�W"_�ҩ�����͗Rk��( ���[T�;l wB���Ea��H'�%�H�샫�Ֆ(��q�;���kYb��ښ�X��������6�$������!��߷�k5����3,Ѥ�M��b�q��M��4�p�.4䢎��6�J�8
\�V6s� ���`�fw7X�ͅxG|S���n�0��6�*'�8���,� ��;�ĥ L w
��<��O�JB<:��ʑ�0�sU��*  ͽ��#���;���9c����-ZF干h55��c�i �� P`�%�i�0��I�Q�{F*�N��x� f�'Y�������u�Ƒȣ~���w�ޙ���ۘ:���7��`)��$�I[yY|S��@Gw�<�ƍ#�"��d@�8�1'��~�~E����^�L$��=`��f�4G��%e�J$M�3�{�	hk��o>7*�$����m�6�k׺��GqT=��U 
��*.���um�u���@   '��w]���w�����qT6���
��AwTU@U   x [!T�N5M����ۙ�n��*lWr����
��PU*��Uw�-����}��-ex?�08�1�DQ��
\�}�$���.��7li'J�p�������O]�`�O6��x�̒�I$�j�w�C�i)��U2�l9��KyB�_!�Pߕ�H ;��*�Rej,j,Q��N��@����f�Ⱥ#�s��� Jm$�hOy�p�s�V[t�G5;�Y���F�F�����_p�Y���Z�o�@��!��T:gk�@$�e��,!��2��I�2"��T�m�tYu�N�Et�n�,�ذ��> a����Lj�oH����zg{-l��N�t�N�����18�m"�zO��X%�_53Q�h��Tl��$�o�y-���t"�g��Z�7�O��q1��,\���o� X�I6 I��1��֠ج̣��H���=> ��"�������uu<���8�T	���a��[]�#؞�W�O�k}�{�$'���d"��ȻWL�N�L�1tz/�+j`����_aF�_h�W������%y ��B�9���u��u�Ҥ�M �$�l ����� ���o��������n�v��ݯu�����ޮ��립��vF��-�^��n.��qݿm���귞�k3r�|^�-����_e��C(0`�b���B����s��jmL�&�;�K��{׍
~�ް9�i'�RH����bc��4��kv�ܬx��U5y��W�c64u����.���0F�oa	�	4>O��0��%�ws���ˍ�lye� !��J&�oW;c����.�U��wC�v��fu7�[���bW!����c=y�xb�Wv �0/ԉ���~�Y缶VX��+�����ƊˍԮ
�P�P+�?z�z����@\���s�i0�3���:��hM%m��� w Umd!&�i�[K>ݹy��Nv����'䭌s��uW�5rw"�����\I(��!�z�Y )m�!�;�8G�YT'T���٤��᪽�J_N�i�vw�p��2/�:6
87��3���5ɈV ������^��u��/tN�R'�Ǣ\�P���n,*��Fm���f�l؊yr����i�?\&�~�����y�jE�������Ͳ�A ������KƮ�w�ݺ�8┦E�8l��Y�]V�^��of
���fV��|g���y�ۻ���/jQ�{E�� 
$��q=��Ӝ`mvA�T<�ߧ��-q�n�>�N����GNr6���:E�u�X��Ǘ�ǹ6�ew��uB�$)��M$�,B �)�P�T^�S���=�X��2pW[q"��>��96�xUq�n�˼�pO��lddhIm|N,PV��'2Ym��i$�sZF�W����8��W_� �4�Y�JL�$g�qz�k_n�����K%�:��\w0�2�����I�����%"\�} P<luse�ƣr��1ǖ���ڱ�����V�Њ�1�;�!l�t�؝��O�D��YM����m&Ki4	L_���'N�7�:k���j�\���]����s�[ɻ�lwH�"�(��Qz�j�� @'u�O�t�8�V���u��ĉ�W%hi�A�#��y��НV�=Ѭ�1���QM�l��3��S�P�6�m&�V���y���p4M.n���Ã��JM���{�#	�s�d�"4�Gv�O��j��@w3���ۋ��*�rm��� m���m$���i��0ʳ��5bc5B�PJ��w�@3H�(�}����#xoI�j�n+`��f���Ǩ�,c�p|I%$B��r"�N`8����	��Y���%���3H�b�]�0ô��� y��ʙ�hBI�D�sչ��?YX֬�HZE��*�="�e�߲��p�I˗6�x.u����y�kk�@ʹ�4(����VLb=��`F�r����1)He�A%�$��$�L�h��D @%"Hg�!�?0,Aa&Q���N�5fx����m���QZr��]�L�׮��w8�Y������-.ŜXKl��*LH�����5�λ�k�tU�1:�L-�,�t��;K���@6���,��]� �D�T{}��̤b�&TRUosL;��gn�{n{��û�V_��ߪ�6�`\�گUBةUT   ��ޗ�o��뮻���P�  � �@���*�<   <�S�een��ݧuڵ��6��ڻfl��*�Mݲ�v�5���߉ܿ: o��J}��k��s��r�Z�L�0 �x��^����谞X�	lz��+W�Ƈ3('G�j(���f�69^o@CY����F����J6 �Uu?j�E� gb��F�����E� $�����׸����*��(��9XOG��-���6}ej��2�
හ؊�]��a�ښ�{�̉���(�C����OC���1��(3H�i���l��I��J�n뻿�n-�o]�V����]f�8{7JNI�K�ObvG-q�2K�w�� h.�,}O�+"���8��lxO��B����㈰�I%tH5���a+	S�F� 4	�u���I\��$f��B�R�4c��]�*BTv�aGXT��<g�S:�����E����lwv-�����w��)�Hyx
k:Teo414�,R���q��8�d^	���������E��%�6�25�	l��a�@�~�QA��@���$��
 ���˳h�3ʰ�j$��^�ujf!T��ܱ3Ff�%��PI"�$�l6�m���' ;�;��3z�v�om�n�i���]�;�kO{���}g��u�sڞ�[Q��Ǔ��v��[w�y�Gj�+ݹ�of[vٍ��}�ݓ��<��#(J ���#�Tz���wG*lp�0�&f�5g4��d߫*v�� ��"ȁ��)"��
���D�Ȱ�� �K�Ly/���_j��7jYip�|:�Pzm;e:�k�י��ysݕ)�h���o[x#���dl�wf�h����ը��Ӧ����l�9*YYN6�v�����
��=!����r�b����+W���ӿ��*i\��T�I�}���~�q(�88��ϷK�~�*�8r�\�4r���ϝv�+�I�"�u�H�\4�V6`$�c�]� ���2���&�$[m_h2ʏ-3�t����?���hJ�����1�<ZhN��D�Y����S�'��O�}m���M��d�&�5A"�>��jEEn�v�W�Ć��EB��ٍ�� `�>o'^T�N�);j%{�'h�̒�% )q�;'ۋͼ�`遝�q��R���+B}~۸Q�L�Q�v&fר[�&*�n��+O�D!��Hq�������D)پY��xŵ�t���M5tzI}�N��x�Q64�r�M�v����^M{���������q�C{�/��g��KLP���s^v�f�&-O�����C�j�1@AM��ϴC�¸:�OmS5��ŋ�x����>Ǣ8hǧ�$3�����\<��$�<i�[�J(��-���`�qlT[�u�n��Us����q^N�����b�7�S��9��D�8,���C�(�j�f��H��i��Lxe;t�|d�� i*n�8��h)#���W��LZ]Ve��Z�X�
��zs�۹�t���m���Һ�MYb��p���&�����: �f�L��t�ǊF��Qf�^��G�;���:����A��	�Q�I��&Q�6�Fg��ŭG)W�r{��Qͻb�]���v2U�u$�2�zx��'x{�y.�j�T��A�P��JKJF�E�X�7�u��\�m�+���7w��{z���e	c.�s���#Y!GG�V������PO�'wf�y�8�vMƮGx)uVF-E&_�*�s� +�&�$�M%M�Im�]����fۻ�ݷV�HA�Qct`;.l�ܭ���G~�@�9�����$5m���)$�������-��H�n���<$��_c=H�����)lNF^&�z1EɏH(�iц�67#7P��^�aHE��Z��2��g�7�'��]FW�J�k0�qI%E=��yܧ���~g�(+������ε�綼ۚ{��*�k���+4h ���e����X�(|�R��͔�m�%��H��hT�����ʿ���������m�y�ϭ�ױ������������ $ ����� ����� I!$���!Lx�1$��Մ� {��}Xj�Y		���  @( �� ���HBH��BC�! O�پc�׿������$	��?��~��7������~��?�O������?��?�����X B@�������� ���F �O�a?��oʓ��=ړ�����_���� ! ����o��_�~���?����=���O}��������2�E�B ��   @a$ �� �?�|������ ,�?3�o�O�����^���O�����O��� ���=���7�~?��տ�����O�O�=������� H���?/���/��?��ń O�BI?x B@_�!��?́B c��}�� x	��l���J��O'�|����7�@ ?����~�� �������������~��?��'����t�� H �?��%�_��� ����~�����=
`����C~���>����~y���χ���3��� ! ��?�?����??�~�������~?3�	�?��#�����|��	�}����~�����d�Mg�d	̋~�Ad����v@��������\  N�         ��(�P       ��       �)@   	
%(D 
�U

( 
 
 (  �ɦ�'Q��R�Bl�U�%Iт�K�j�9EwS,!U]��UY��Pk
��e  �� <E D���
)ӓR��v�
CX�X�gW3R�Mb�32�(֥%SwtH��N�$�eQkU(�Ѥ  f�Ѫvy�0�*ڄ����Rt�ER��9:�ERsjU�J�F�⽙S��y�\Ԋ@  �    ���J�ݸH�ͪ)�T�rU�SZ*�M2��F�J���֢�u:l�J��ݹ
ڥ  R����ywn���w���ڎ��	�:z҇F�s�С��E&������J�Zs���к  �Ĩ� 
<�{�hWG;�<�s u݁<<�׭6sgAJu�����4e�9ǔq�o{���trQG{u�f���B� �K�����s���B�`��5���G.��B�Z�s��{=��^�d�*vw`iA��N��\焽�Ӡ4  ��@R�*�V+��ԓӗB��J���W���mU:h��B�vn�N���.�9ǅ9�vzꁚ�� ���
:8 J����7�p%�P/1�(7��
=w���:2:�<=�t��Jz2 A��FOTz�p � � p �( �W� ��=���V���QK�=!�K���=���[����K0zt]���Y�Yѻz�I�ݰ�iJ	kF    E?	JR�20FaMd`O�JT�4`0` 	�4��F��`  a<z��4�� �� #	�S���UHi��ɠd`CF� h<��hI��4�ɚ�?Tzjz���mM�S�Ԏ>��~��W��G��̍�>�0��º��_}�����[�<}gt������?ϟˤ���I�t�:t��}�N���N��w9��I��N�t�����I���'�I	8$�Г�iӻ�t������;�wwt��I�;��wt��ߣ��1���������;��ww��rO���,��C��������X_u��C���1>|�GȈ��c��3+���g~��!��KvUX�5��S�l��h��?X�2E�JD�o1h,]���:,�DWf�(�L�َf=U���el�y��J	�4�����J�>�%�!����[���3.�=���zs7�4q�޼��eݻn囬�Y�7U�ۣ�[u.��ƠG�*ق�"�DT�������˼��P[ѧL܏N%�e�+o6G��7F1x��ҳ�҅���Nf����i-���MB:X�̻"�!�SU�4��X����qƶ���5&X�ˀ�HFU��v+qk.]y&��u^Vj|��x���Y�Zҥ�H�W���V�Y�fU��VY'u�,:�:2�*9�;��nY[
�b�w�j��O��wVU�",��ef�%���'j�:p��!LcZ��T��v��sZtS0֐%�ًKϕ����a[wpf,"�� Н�ְ�"-��N�֩�m�h�Z䘍cZ�ML����nY4A+}�R��W��I��Ê<��}_Y4K�6\5��
Xh�[��,Wԓ�|��֎��Iz��N�+E�N��RV��E�φWO"N��'I��'I�������z���g�,�V#D�Ȧ������6��0A7S͹򀼭�M�dv��R�a�E[�J��p�W� ��Pn�ť�e��/~���
��揄h��`�	\Ё���NM����!�>7��9�N��5�	OJ�Z�A��o+Mnf���N�e� l��t�aP$Q�W���yCmڱ�P��ӈ����:�=ξ�����t��*GC�(�fb*�n�6��%ٍ*8�1�%a����k�S6:�i��'�4�kQ+��kh ��c�	���j	e��5���6�5uw!ܩeQ��*f]����dʘU�z/v2�/4�Q��f(sv^L��Pj��X(C�ޭ���k#`�K.ɺ���#u�7p��IUCr������v�}e7�����h����.��4��#k�9v�hK/AH5�������
Uw���m�!3Eۻ˩���.��K�����9�2!����޴w�,o��ViٛZ6n�%^���C.Lܠ�˺Y�g���G5�N��9�ّaޗ6����9��R���MmǢ�׻�q�#j�è�nn��U�җ�����6�m]
�tf��`�˼Oo	V7�"��w���uk%�w��&h��Yʽ��'tf�gh��0g��P��0Kͣ��m9&c©e1yjn��Sj)���o�,��sn�7�=�T��\3����֛F���=R�hx���[YOw���opV�X3q�:�+
�O
{i��Rm��Pdo/�X�'b��h�����^�r�AO�����l))b�̧d�L
�dU.�6�k)�N��Y���ںv�����a�Rw7r�Q&U�1�&[�!�k�t*�]e�
���.�y�z��3+6���Z�B&�t6=n�Q_UW�>����/����2�o1Ԭ��a�fA� �2X'�!��X�V����*�fû�1��$��f�e�Lgم[Ǐ�xĭL��c4�tn[rkF�^F������H�5��t-+u�]��9Y� �i���]Q!�,׹i�{d�(Mr�cv1�����^�՚o(MHCm���ֱeXW��,YQ�b�����'��ܽ�@�<6�W1�b���@;���A�I�i�����T%�u���J�0���5�j�9����*�O+n�F9s��F��5�
U�Ƙ��[�
�����]6A��).�b�*I�=���������mc�Y�^4�I����BV���2i�.�QvQM�Zѭ{7ie�H�GI��F�k�E4v����M]���e$t��_;V��e�zHŌ��@�Z�m�n#��dr�<���G�(�����Xu���%�����@�������Gn�񕪯L��^!��l�^TD�	���40�YX�ͷL�8��k�� ����5��9���coh�J���AON�XO$
zn뙦�^Gb�<��d��e�Y{$����+Eĩ�[��P��PVV�]�j�e`�w0�.���SA<Y=�E�©��f%�SZ$U4&W[����ma�ZʱJ������,ݫ�Øu%t�t�>��]Ů)���V��
��J£�:�dT�D�k3Fh+Tn^^H	��IQ[Ll%��R���UM�E��ZtK�wwfV�x�A�vd��&�k-J(a���iu��m�.�e�Akl	�<�)@<�M�e]b�Qm:z/v���X�VT��s6�k�Nܣ���@NV�$�#i��9f;2]�w��¼���n�32+wnRG4=�s%,�"�+*+�ֳxk,-Pֈ7��ڽÒn���N�)4��uh	�Y�TV3Nl�^P�]��f*w��@O�hɗ��0��R���H�o#sh	F�3����;G�u�nY˾�A�jsBZFGV��^�{y�Z�v��Y�U�d�.�L[�]���7]��e+:�vY�毣�r���S�U1A�f�m͙y��Qi����n�ˆ�l
S^,��,����j�I�L�5���7
*Q��N��X�?ql��)�X��b�7mُ^��B�m�'w���]Y��m���j��+n�8�P��4}�W�:���p���,��Ѵ��e�C�*�D�}���������nL���OUU<���i�*t{ �3#�8f�˻��ܥ?��#J�l �(.2�d�M�c*+;9t�o�%ru���vn�1#��|��AV�aJ*�z�m�,��K���7�����eN&\��p,���`͎�l��EǕxt�-�vװ�tt\�Hkv.恣;v疎x��&sH[؋ʼ*�ڣW�6ؘ���^X��%�"l����4�&���`�ˑj]+-NRIȓ17bS�O'�/t�3�r�&͑��:�[�$骱�+�)W6e+�R��p�8��X��\v�Ч�@Wt�x;��x���r����Ť��F��;���|�A�dOr��v1�+^SV-��Ť�t����O��%K�W�h��`�ѷ��S3r��q���Z��2(��k�q}�dZ�r��]��Uڭ഑�6�Em�fn˿�^l���Ѻ����)ܗx7+m�Ba9W ��e,",�4\X�]�L�U*���ZnYw�w0(F�f�f�F�b�MK֭�7��9!�M�ܪw��Rä	��, #DY>�`����m����(!�L4k�T�9Qh�eL]��R�̸.�10W�P��٪U{��Ê�oM���M�W�;��iI�5�MҰ��)�3VQ�Ol�AZ�Y]��e?�C�y�&�w��Zm����`���k�.D�T��7�
�O�J�l�
��.nȠ���Q�@?1t�
���̖}Ϻ�It�e���a4w-]n�/�ܑ����d�0���n�؂�1j����-�B��*�VP=�������6���UN9�VT��-��*f�IR�� ��lYu�os���X�]�ueI�V��
�S�ۨX'zs�WZ�WɊ��<yr��.�n��^<���G��MB�;�f+����+M�����Ô�դ�v��BI1�rn�����T]@�؆a����a��י��S�/Qx?�[!�l�
����[2���a�T�'b�u�-	��pS�L�͛��n+WySVM��X7P+�cB�/rc�١K.�^�3j̔�[V �D�;Go0醚��3�s��$?��ɮ�˽��\�I=Kwe㿍%-��6�]mF�.*[sr�
��)Q��[D,�Q�wR9VR�s=}V�P�}4b��EVX�}��4v���bnV-q�X�I��$-OC7uG��p��-
��+R��{B�o�A�r�-�R��"^�3K�]��>u1�I�fHU��M��t�
�cjxI-`4�ZW��7�x��E�{�.4��༦1I�&����:�݇��X��ݢ����v�mnG�L�;��24Z�F<�sES]+����uħۊA\�Z�	=�VP���@��o�6��U��PD��0,Xuaú�olx*��ШZ/\Z�E<Ε�[����i\���(;����jb��B��Ƿ�c�q��1�
�����F7dO �f,֢����
�by}����%=�I
1n����i%�,��f-{��+�ݺ�ݭ�YX[�G�s(��*�d��L�w&�u��Gk�3�'0��������r��	�v���d�Ұ�j�<�]k�N�Q�7Gw8��p�����]i7[��u�l|j*�����A=��X4�;W�:�䯫���?RG����mwJ���
c���^�� {*�����vv�7P��b�;��X�<c!��o/":�B�MQ��F���һ�I3�Qf��t���nL�)|-k�F=���[iW��P*[����Cd4ͽ Vܶ�F��%�7U�Ҷ/;���y�;1y�#K�m�I̦�;(9�QX�#���^K�t�j�N��d �\�r<��}���܏��{�������݉ӺObt���h��}�O_����U�]�V�%f��!˸,�Ŧ�b8�l���o`�TK��;8��W#�~���}J���'������$�=���y���<;�������O��t�Ow�w��{=ӻVO^������d<kވYc��������9��֝'�6��ԟ�� ����N�,��}�;ܒq���Ϭ�3뾾g�}g�������o�              6�   f�ݶ�� m��jA��`k           l                        h              �`�` dHm�Í�                        m� �`[�-� 5�����n��-��l��     �]�0Zlm�������mm�2���r�m lN�4l��!���Yg[��5�R                                      �6��Lk"��� l   �`                  6�         � �m�l�i6څm��e�6�6� ���m    l                         ��l��l-�m       ��� ڑ���              � �`    �                             �[ �]��Rc�!�[��YL�+6��vt�Kf�¼i�C�-�\)4İui�f\h�y�6����Gg6Դ�[�+F�E)��Sp]q��gN��i���e\�^�ڛ'T�[l�3K�]�C�X[5��q���Z���XJ#�b86kQ`ڙ62��5��;6�/&��P�%M�����5\�˰K{�HFD�9tj�v��+�֕+��fZL�]4�$�:9!�����!��8&�m���cK��G]�A"it�YL�,�
G��ڈ�6Xm�!K[�"{v�����:m8'!�ݎȷL�M�ڕp�jι
ie�fc��� #e�qme��	a�UU*rZm`h��a�J��uԉ���Tc�4�����K��m)h��M�f�\�m	�U43,���%i���3��5SCT�4�K0AH#���KB G36��A͸��գ��.%����č�+�]k\K�])��u���k�tP�#<�,�h`�0Ћm�"R�D�m)]�k��pF���][�eԼÄv(��3Y���b˱
�Lf��5q��Mbj�Sr׈lۅy�����T��UÀ���FS���u�p��H�ݲ(���m���J�m�]��vt-����p��qC5S�l6�-{f)h���Rh���f[�7h�A����hl�I�#K
�����%�Wf�J�]�\�+��a��Te.���ѩ�G^4ɥ��]Qe���u�],��.s�M]3��,ݨ�V��ۅ���J%[�,2!������&)Y���Sm���%�C*�idX�i��5�]t��6�.fcp���BZ�W[4���b �a����Ԍ&ekEHE��d3Uu���4�E��ѷU��f���G0�LtI:k�u��鹛�yu��[Z$���fi�LZmp2��ihc@Z�5��-����)1^+�mkdVJ����Й.�U+,.��wk4�X��O�t��E��,z&9ˑ�]9�9'7�t�D��mf��,
i��5�kE+6\8�����[���l�f���Y��-�-J�l���lA��
�su
�c��V҇���v�:�z[j�+Z��Y��4�:��m��&��Д��+�ю��I�KXL�=lL�h@&� ؉+v�)\]����]V�D��og6,dY��9��v��:��6dm���Y��r�Ͳ2����i9�1��R���r�[�l��PuѺ����:/��a�t�aCV˱JK��9�Rᚚ�:k.ЮU��1n��9{^��H���7-R��vK�F6J�i�]u��J8Hml��m7f٢⧍����]-�MD�{sqj�]���+T�4bWm��%�V���mfu��\6a�K+3t)G'W[���;�^t��İ׊8P ��щ�Z�u-�MXSm+u��"-�m"k�[f��6�Yv����jɎ�sk�����^�e��j�"Y�g
�U�ׄ�BR���ȇm�e�5� ��ʷ]+�f�E�g%X_fݫ���䛍f6��K7C�ޭ�F��^ȶ7�ؽw9bv��N[�s�Eܭ!n�V�e�������bU�#C:�˴aΎ��!P͛M���l��c��̗%�Nn�7Q)	�Y�m��.T��-�Z=f�M���tց��j�ʍv�hA����8�t��7p�cih<fʣ붗����)l!JK���H��FФ�˭���V�Ʊq,%&KH1�����3�L@�ct�
l��Q�ͩ�҆m[�H�T���k�����Iu�ڱ�@ht�n���t�f��H��[�cFB�ۖ����lY�zh�7	�c��Rٮ�Q����h�2��ɹ��n֫���gm'T�7YY]
p�K6�riK0����SG[n��^Թ���b�:M|�<�r^�MfDT�;^�X6��fhC:i������p�RL��Xt��\�<��zfvb]������ P�2ͩ^%ģK2
l�X�56m-��x �V�P���X.IE�]q�[Y�$#L�hJ�$����0��E�J��g/:˃��3���H��\MaZ����2�I\�6Ĳ�<f[)��[(���f�xż�q
)�홑�-z�%W6�R3T�k�]V٥űy������9٬v�n�kVؑ͠,�,��].�mBZZ^��&�GA������\�n6�e��n)%�b� \f�[4My�&�m9�kMɴ�`+����kz�CG[c� K[�-�p��MdvZ��� �l�Ԩp�ǆзj�IoRj]c.!��eXu��Q#��^�Am.���ݣn%[h���T�L�j��]VG/b:�Y�;X�EgK���mz�@�rYs�͵�U,tZF�X�u�9,ڧ2��Pe�[�Vh���a��l-��Q�S��\D-�Kk�E�t*�C`�%��7ًs��Z�]kt0A�
T��	�]i�EM ٌ����t��h�hY�[�.�Y^)�#�m.�ZH�-�gD��K�Yݖ��Ke-�rlǈ�����W[�K2�h��8��
˄����فjAn��f���[A�-ohGj�*�kQ��5�1c���n�T�"]s�ңqn���ہ��;V�2;�3�f�]��l$sQ.��3n�&/��\in�+�ݷS�Й&"J�u�)��51f�6�mAM4,3r�	Z��Ms3i������j�˥˫���3`eA:[��bٮ��Z�%P�ŮT։7:s7k$�v��\ٍku)�&��h9h�q���h�N1��!f�n��uڮv�+2il�t���]WZ8X�pԅ9j���w5m���M�� L�;m^�M5͕y����K�100���#5�-�e3�Y��ۂl�k+��m��5FbVʖ���]i����d7��f�ڮ[�m.�4LF�i�.��6�kf��K�z��r�D�a�T�;m.���Ds*f]X"d�&����f��E�雈U��X�A�X5�J�]�kWP�%o0�1l"�<��h�XS�ڋ���0�Ҧ.�[�V���0����e�x�uЉ��ka-�K���U�G�h��jXښl�B`�f�҄,�Ҧ2�1&�6bbSky�BhF6�jj]���eT+1eĩ�c`mck/a3�S;5N�J��#�P��:i�v�J���Zl�^`��I��`��.&�l��X��[�jc&�u�KF[������f���[5l��lAuF�
�D�5�450�v愁���c�Ŷ�����7T�svH�f"�/-l�ʤc��U(V�i�����-�^Ew-s-��-!<��'�_>�Yw��������'|�����'~=�Ϥ�O������>��?)�|��O���t�OGN��'t{���;��Bw�βK�|0dN����$���1���t���;�I�I'pt�;�t��O�	!>�_�?A�>��~��P�����TpHҒ���ڹ���х]�l��Cd@?�1LΪ�!����ƺ��h.0��ƘYp�%�ԩ��a�\P��=֫89;�U.Oo�X&�Q?�z�jԭ�05�����o��j�&�>5�80o�{t� {��`�4얗;�3z��4g���n����m��P������\�B�A4Je���j�JL���lڅ�Q���0ʂ�-���ә�t��Rc �>*�Ǵ)��&&8��~JL��"���[�y0&�L���.ޫ�P�P�V�f���zK7�;�rZ���ׂ�X�$�wGLpH��L�k<�;ݴI��l�ᇈt�M؛�ײ�&�
 өs˅ю��ު"�P/N���o�N#^4e�B�w�&р�4�S �����n�O�|����~�Y���t�֦a}�Ha���ʍZ�D]����MF�U�6T�C�� A�kU�{��:@e�����`mo�
Im�ր�`Z�   #h_/�^E�MmӧKے����ɭ�f�Ja�m�������)�⟏��on�̳e�m�=ab�]t�ڴ�d뙗;kydk�vU�kY25;k�3@�\�p�L�ZpF��=I�����ԬԶ�L��)�Ԛa���gwk�1&B�a��Q��uj4O��z�9-l���JQ�#z¸q�;�kSz�!�is�ኄzO
7#�2��B����o.3Ӕ5&��9��q >ࣣ3�
!� �	�;Q�F�r-$�0F���I%I$�m�1t��%\Ț�YΛmQ�;%� A�E��0����B,vJ&'q[�b�C	x�
|@t
�A��y1���7�i�P�fQc]s�Ձ�to
���z��AK�ܽ%���Z^���=��� Ƹ-8ϴ���wM�YL#Z6�H�Օ2�\,E�D�$]�Gi�q�J�O{ovD�<>�R�Rf�;������4�rL�>E[I����i�
�Q����V꾇LK�<��vyc��l�>���_c�,�
Q�&L�Ǭ���71׹\��6s5�J�^~�L�}� Y�*Z���N.�*�+/����9m��ݩs8�gU`ۜ��#�Y�/�u������T���A�a"�Ng*[�-�[�e4t��dS�*AD�P���R�	8�8�i$�eCD2�v�ܱv���rN#�9]?����`�],��C���ns���4ej�Y�I�'':$�D-3M;�̅b�ZKa��,��;���7%���v��,`�|N]ӭ�~��� �:+��.��0��9��Nh*l�`R,������#��&4�J��u`�4�h�3Đx<5o�z���RhP���rS/;j��\U�u)�%�D�qB�q��O��X6 ^>�T��za����n? M�O�h�7����6q�:�S=H���$�N$ڍ(�"88��j�@,�3�5�.)0�YM�w`��!( 'M�@"{����Ocu��h�6�4�c~�Ee�˻Ap��Ru�YGp�`��v�[h^q���e�pD�[ts�h�ڼ�����������?h�Xdr���,^_��W�zmE���'2��k��t��@�r�h��[�d1#|,m4s2Z�Cz��X`4�_��x�*��^��hd�;�)\=n�/<�З��o.g���K�� �yghװ�9����P�7��
I����h<�Rv?���;,x�o15��W�s|�gF#Ĩ}�<��^��ᛏϡ�3;:'b�J���2te�8�N6"��Į��3K��;���˃{� ���xX;�.w���tFvr�i��;P&Ԫ����Zr�X��UȁÝ/?���dֹ�䲣,/C�co=f^� Q��}~ȷ�ma��1Z8D�
K�NE+��zE�À�I6�I�`���P�"����z�mn4��9v�����Ɏ����pP�61F�D2,�{�v�����c6��	U�i\�7sAM�T8mȾuE��'F���o�������,�3=�K~#h�|9�>*4-�{�=�x?X�^��e��dRg��Te�IN��{F8_�Ǻuh�}���xj�����}.mfW��h`��/Uv�5s�A����w�KV���=1�`�(p֗i�ʕS3y��yDq�vz�7�ӊ��⸰Y% Њ�bG;�Q���g�Z1�D��**�f�|PBW3U��>�Y�>
���.����� �a8N3�[�k9ۊ�D.�s$%E	㓵��u<��L��}.��7�'e�"q�q��X�0:�ƧzɴE2�� �|�U�ugO[�4�'Tf��|��_6���[n��7��R5�Y�(��Z3$��v���8��r{AΉ��;|���"	�).>8-ةBV+�0bM���6[3]�dq�wf�64ŵ�#��E�.6�� 5ysN�
�Θ":���Χ#n�Q�B��؂!��L:�w<�R>�pn�M��5b�9��LX�ghV�xT��<�If3�2��4d(\��M_��:a�`؈�4��:wH��8����\��Zp`]�N
k�{s:k��fp��F��r���xٝ׉]Fo��:|v:i$� �S�v&mW0�l �` lְ:�X��c(�W0f�Cǉ��H������I�J��\l�T�W�t��:Fٯ٤�ݮ�Uér�с,f��"m#
keס��s��f�e	MԕP1�*��Jr�ee�]ͱn�t�7t�=*h�%�mM����S߼���hJ�'�W���}�6���{�p4�)�X���S���?�O'VJ�nvX��xԥl֞JT�Oe�4�`r��s�G�(�Ac��<b[|��[�4�4CA�6{�TFMT�o����=j��)���	W:ݶa�E�X��,irT�gK�\��mH(�Ih
���y�,l�+����flG'L�Xc,��;R�nhL4�/����
v����Q�7V�C��	uv�:@�[��lX�x�q%��9����:��{Cl�a8�@DJZ�}�j� o���rw���t�ڳ��*B�i���X�Ax[0u�M�*��3RM邅��ɸ��y=6-�%k7�g�)Yk72��w��j(!͌1���G�VyTTov6�0�+^�Q��->�hv���S�0�=�Ҙw{�0���A))ZM��v��F(ޠ�:�ѽY�#b��N��˞�к��w3�Z��*l]:���Om���-E0<���S�׫'�ͫ�/�FOϿ�c6�5�g]�su�7��Y��KcP��d���ҋ���������y��[�5ß3ʏo'�}�fל����6�Tk��u�������^���\�zt�V+��R�X2֋�0aS��r������[����=θ���ip��1�6�����\d^� Ƶ�An=�`�h�:8<:U�]����e�Se�k6x:�^������ff�]��E�#_���_��e�6����a�x���߯z	N�SD�^,V��'u�����?q�/���_%w&Lu��]˺�`r���qSQ�x�X)�G�q�7u�9�4uft������gȧ�Mm�`�b1��46b�YI{uQ,q�[�c���հ�y�۫U���u���伽q��Y���,��;����oe�t�p�X�X�jg,�S�Z�9%e��cEl�YG�Ց��ϕ��R����l6�����yN�=^����D(B++��%\.�wn*�s�b�n���+D�G��d3D��w0���r*^������l~d���x�NF�n�����O
�2{o����;��w�Z��s%�@2�
��~�vn���(�'���,]M\.������Z���q����{-�l�a���v񻰟g�7����@�x���.��n/����M�/�ڜ�1������������k&���ɵ��sJWm`��4�m� L�n��������P��|a&Cf.՚��\ޚ�p���B��vg�/n�q.��E�<���y�˛�T�	&�8X��A�J�eҝ����*l�@þ�T�^��}X/ʠ�6�oN	��!�t2Ŭ<wn�*+Xx^`ўǮ����n=i��T0���eV��8�Clk�9ZZz�u�s�<%�5)�M{��y�s��f����l)��[pbj��Ʒ2�Ggd�pX-7=/�ܵ��}鯮�ey�����㓗��{(���|+z�:������M@0�1��e�ڸ�r�J������HV�{e�ތ�8��;wҶ6�)��-�`K����+!j�w���x�u�^�	}	�[$����&~in��;3*X�ZWK�gqb���K�O8��D�	��9�5p�=r�]���=sb%��*��Oݘ�-��rs=�T]�����0yN���D�z��w�9'E宽���$�hy��ݫ�M��b>��N��Б���M���tY��U����0������=L4�4�������U����v)�\�gg����He�N]"?4�`w��7��2�V,H#>}�)RC�X�i%�	k�MCS�W���m�  ��nF�-� �h 6��� l�741wΔ�Erx��W��ڭ�2��qe�i�Q�In��-���pV̡jd�u�7K����PM�X�.� L�K1(:2�:��:Y[Mm5;A��ٸ�[���W5���n�hն6���� �&Ќ����{��|L��z�^�5.�{_t���]A؞�<��`�n��;Y��Wwh���۾ʥw�Ū�_�cG��{���}�I��D��-�ż�������1<����'N/.�F�䞒%�j��Pm��h@J0�*U[����%!o^�:�[�ߛ��z{j���Z\���u��U��ف{0������IZTM��ԗ��]�����[��[�zfjZ��>N-���e���JQf�m���\�A�]8��E�I���}[�~Y�j��)�TrNj7���1;�Jf74��҃L�3�����}}5���g�q9�{7�0���7�us㺇��=�j

p%�8��m��uK{�od�+�%��6\G����4.�<S����y#^���·��Wژ����kZ�s�������a��ϭ"�[����^�<�Mطfl]z#����H�=�t���E57l.��]hˑݣ�ll�侫�H�yE��/\�*�.�47�E�� ܰ����Ἦ�E�IP`�W���V��@��ĸ�]�}�7r���e��.����eLV�8�^�wV'��` Fyj��ힼ�Q3����8o���ҵ�e��U�x�]�	tx^V�y7v�Fi�M=D�ÎlǞ~�I�a��|��S�
^��=0<4�`N�Ǻw6���ʸ���s�@���;R�r�����ӆ[v[S��
�1�LV��v�Cb>gq�MXAC;���ܴP�HQ��&͢C�D� n�Z�!�0-�K�h�԰�-�G9n���]mC>Yv��A�ytܘ�ͬ߸-ՙ�T%��P��!�y�R� ��ⵒ�M.�]oj���[ؕz팓jflh������1�W��m��m� �\`�6�      �  m�4�v     �f�z�� ������m�N����      -��m�      &�m�kX     ,6� ��`  6�m�     �Ye�4��9Ӭ�4����ׯ���M�p�6Yf�^G%��kn��ڑ�c���֤1�IIVʭ�h��Z�9t��$� �5���ƻ!e�
2���J�Wh&�Դ#l*�p�\�{@�fLӶ���Kx��	cf� )M�Ү�֓SR��T�*B���(�R�S[�h@i�Y�ۛY�����^��I�0��kmI�g��چ�^����&06�ɴ����	��c�QQ�Is�k)���廌�Z,ū��V��Z���˹pi�h��$��lM�2ڥ�[@��f�\5\��G�f�nШ�Si�"&���f�@b�[�Z��8%��ͩ����c-u�Z�q��cn�X��M��4 ��kͻk��%��F[SWm��ֻТ4��g\m����ZF�U���m�^�h�4)t(˝K�-�ݬv��(Yq�k��Sf4�pYi�vcu9X��N�Y�6�t2]K6�7T����b���ZL�We��l�1��nR�ܮ���m�7m�l�F5�i�*��,2�̭���ؗn�oYet������9].B:Fb�)��Ѧ�;2m��k]���Օ��6�ͻ3I��]s 	"I��ڦ��*ޞ��%��f�����pE��g4���tK�^���Y�]Ne`]����&�EQ]4ԕic�M+�1.<�Ǣ?�:|���R{��>�>>���x;�N��q�:��Ĕ�>�u;����Ν�>���~u��w�ؘ�>	=�;�;��gc���{��|މN��=ȓ��	7:�j�ܺ�*(%��-�H�6Z�`�w7n��k��dhCM����H���L|D|l��#�>�LI;���>޷D���w���w�=�n���W�|���@�DDxxG��{�W��}����]�?�������/L}r��>B>���츏�Y3�������z��wS����޽i�����"H�8G������E�C=^���<����#�c�G�?G�8}�������� ��ޓA`��_���Dv_��0��p�@_������}����1{�{���B#�} C������窱�$	ғ�v=���D�&�g�'��c��s~����IP�}#�G���>�1s��
1v|@��'Dp� �����p��۟�G�]�@\J��"����>�"''t�I��t��xӶd����t�I}����W�:���Fwu�j��
��[s��I�/��4���ýCa�hI���b̛�_�nЖ'���#�U��[����Q���.N��E
]]��QЃL���;���yk��1z��`w���������l��:�ӥr��h�v�Ա�V�m5'N��I 3c5f.:{�ʑ��k#p���91�LTG�x@��_�˪��s��קX�Zs�lv+V�WŊ��ާ1,Z�QR"���u�W�=Л"���&��+r{�Pm/Z^~JA�G.��C���2H�G/nj+�0[$�S���6v�OD�����==*i��<Kv���V��W]}�w�ͣO';���V^���M6Q	3בz[�����{}�c�:����W����]���=��K;����\���	0z2jww�X�������O���\����V�v{�P��L�UNΊ�u�&�� i)�h�.��o1�Wc]�oǺp{��޹cn��v� �fH�˶��'C[��^��Kz�k�o���U����]ܐ�up���U�n���4���ή����7B����� �eI}������,U�2Q��
̫7���2>���ܞy�x���i�E&I-�:��v�r�J� >t'��`�kld���g.tf�Ko�9���|�]�]�\����`̻��V~�L܊���쩃/����Fu�z,W����
�e��ck�����+JH6�LLl5G�z<|��Q�fy����V1��S�qVT�n_a���?���t�wI�~�΁fl����$���B]�&�;ny�L�������rbt��ö&ngRqr�A��U����Ŝ����Q.1����F����wFQS��5��� ����D�s��[ndh^]�"�Y4�4_ 	���'��m��Ƶ��5�d^2�����d�TXl���^�^W���^�Es�5���[��O�>��c�lg{v����o4�N&��59V�+sL-9,}��؇�C�i���'����<a��9|�*��ݡ�)4�#GLYΕ��6=��ί�O�ᱞ~�!��N�D?*�gt/�ܐЄ)����rHFg!d%L��^�P�m��m�i�r����Xv���h � ��;�|�z)uf����]�h�l�팹��+��Bh�2L�r0���J����DR׫�s��L��Mbf� ��l�-V�f���6CcCv��h��3�h�Ժh㱂�4Ș�:��
�)�$#�M���yG��7��K4r�7���7%J��9ܛH��i�\��.��g�->R�a����e�BfI�s7�;!�	�;��^�X'�̭����@������cv�'�c�>$�����.`'o^�t�f�{4],�˱5�N��4�W2Z��]���J�C�Yr\�i�䝱8���/����.or���o�"[	�Ў�{\��1;��8���Į^�ݞ�X��$}|����^�w�&�9��cv� WR� ��2�G+.6�f��6���;:`h�ݯز���rY~���ۧ�J���W�	k��b)v��{�$|T��U�z�:�N��w{�|9�f��t]�&���a�`96q*���'[E.�{m�9���[:�WC늞�������<��<�w&1]{�՗-�y5�/Ns�R��1%s8��a��c	Ԭ�m�dˣ\����ʱ���U�֢�$<�o'����ݾ'a8I�\����Uol�1|�%���$�d���ѣ��KćCN��������G�E����q�hb�Guw[ӪoM�G-��>���v//ٟM�A(��E��w�f���i�ݛ��vŉ����N�/tܯ�ך�I���N�@PXE2�1{|EӨ�/���^�`�=�=NVW_4;%��kY|��2vw�=��u������$�F�p{w�5�|z���pW9��卍��N�n]�.R���ɥR{<��̖�d�O�D�'����ڑYcg�3|��2_�K��q�C֙�^%m�����N!�h��QBK�ɍ���{��r��7�_�z���i��%�tv�s�K��ם:.���Z�&�����T=2�'�7L��}+wk����c����c����3�7���hHŇ�p�^��6�,�kx�"���.��uj�J��z��s��{���=) ��m�VK�Hc�T���l��Aj�VAa�0�y����٭�M�ǆs��Mk�V/��l6��]�v�\�^�W��}�V�+�vo��~[������{����K��h˨b���N	[-Bp��ڨ;���P����X����L˞7-E��ơ<���Z�����L�Ǉ�ڼ�K���Vྕ�8C�ъ�rR���,u�_N���C�vn�T�m��- K�=1X&�������z��CH�I�ut���6��۳�IMl�C0�p���p�Αݳ:��:ҽ�8p;6*H��;�V���і���&�Э�`6P�=�;�ڧ�ur��6����dY{��c���d'��JT�9��u��귆�8c��v��N�p���oU̙w.���q��N1>��r�N�z�F�b��w�n��(oW>�_h��r�U�ڻ�������L�q�vىގ�f�N�r{ڑ�����1Y�8��H�Q+]�)�~�SϺ��Ʈ��I^��_�N�S�:7���v�T*L�a��vدX"+.]DW1m����墻�F�4k��o�)�������yu����R}"f�f�M7�SJ�cf����al%W �1"�[~~�K�m���I��i��m��X���������n�;ǽw��y��o���e&/��]�鞣�0��[4E��5}ܘp
e&�{+F���9A5��hk;�l`G7C*�,��q��;�8�������>���K����=�"~;6�L���v�G��֤MV=Χ�V��C&⠈`�tݹya�p�a�0�X���+�$� ���4,�vx����sK2����X��9,1��6
WDͣhw;M�`�.�[�,���3j�|M��}�|�v� oP
kj���`�  �a���6�c���y��"z2�if
l%6���i�7�[i��KIcu�N��3�4�Qf%��;U%�5���`�\j��V�F�M�c4���N���V���q�N�-]#�YsQ�͠X����[1���si�۫��bs�g���5�߿f䘠�H���$mC5�ug2�tu�)e�ʌSx��7;�bC��κ�����������7���c��r�b���:Wgo�p�-�o6�5q5�K�`�L+є�i&�E�	ԻVڻL�/i۰�n�/n$��l�0Pb����n�pqy�ƪ�#���f:��0z�uw8��R���5t���:St�t��cʟ?s��e�(|
�N���EgzҮ�F�மiƼQC;�@��\�`��p�ش�W�T��]��,J��h����_p!��#nu�Ό�c�W��3J%�M�#jb�;�fat�p����P�.��y=J�*6�t�;�,��!���<�,
�k�gm�s"ɾ4#�y���HLe�ds���/oXi�����|�ޔ���	�=�gq�DՍ�~O)���e]423��Y����iwv����j�-zUQ�/�N��[s;lNC��7���D���GМ�g\�.��\��ƎϮ�v�$ⶕէ&�_<f��gm���Y���oj�����iO-�#&������3Ѣ��Y76.D���G%3��B��5*���N��cz��ʁ��K7�R7� ��xyu�����i���$���߽�����-^�ƅh��ذVS����1��~�U<��²��D���Lg_i2�e���z/z�W.쬮�7�^�}fΉ�M��B�=N�W7�Z�Z}�
��h��:`�0��p$]'Y�o݋3s1�H�3Zۉ�%劯�r��Ժ�<���8M/���}�גhR����`��Џ0It�oh��&�/�rj�3��:��(VN�K�Fٲs����'Xi�e۝\�H�����H_�pL)�����lU����q������{�����+�Rw�z
I�.#::~�*r�yM������ĳ������"Х��ӎ囜��^Ϡw��\&H^�)Fn=Ϻ�:�����S*�0V�wfϓo���l�){�a�eLW���Ay��.�ۀ�癚��y[R �;+�D���c��� �z:)#��W����S�β�{�M�*n��]�S�W�T:u��,K?l�[�z��1��=��4u�5�y�ɰcQ���WN�A�܏646t\�{�$;��Jp�Nf���D����3b��vi��Tn��W��_�O�	ܿg�Z��]f>��;$�<Ki� �"��0�dѺO#����F����V��`N��.�㯧mk�$���[(����+j�q�]h\��'y!��]u��$����]�{3y�;����	;��Ӹ달(����n�Vk|~���<��P�!�Pw�9˞���_'1[��,8!�v��C�\86o2S���G�J��DO~��0���Y�]���u�=��(W3�5�P�Ӈ*;K�Ղa���"�u��^rZ��Nڋ��2��[G��s�o\��mrw!|h=h��L�%���c����\a�0,Y��Mݦ���6�6��f5���ّ�Ec��o'��R�O��ĕ�G:'�U�\ߖ��w���x�B�
�E �zo�:����\��]$:�-]�YeK;Q�xt�R�r��[������!���+��ѹ"�\��8�atN��X��zhm��r=bv���Y��,�w�]Z�۔�op�����+#�Z dױ{L��ُv���v:���[>���vWJ������텙��r�o7	 �(����#������t�u��.*�t��Xvټ�r�޺t�Ƿ�b��AHT�Ɨ"�g^.�+8��ĥ��;Q�z����î�U�,���n.��_rՖ���5x�zi�Oz�K< �b�IX᜗�Wb�ڰ"�ru��J�ɚ���F/{ss���7�"��A��@�q�����/����1�/�ʃ1s}j7�잹�+��=��QpQiw�do^m�����U��O�W:G��p�~�h.�1(�1L�O'�3� o�!5�x�Jp��N�$��C���a=�]f$�5�o�0�Ƣ{z��uF�wHb�u)�v)�G���2mn��)Bpn�CZ��\�*�vu��`� �P��) a�e�mK��Jm�U�fҫ@�	@�pT;��]��E���o����]=Sg�l�Y��,v�u��D���њ�"F�F:�5	�щ���~{�V��|�t91o�Vyp����V Dh����5�J�Q�Æ��u��s���Ptl���~����V��g��.�p��pċ���#�t��./�f�[(��n���w)����}���B�&(��6�6[;C�^��.c7�ۖ�^�o%���
B����c��*����d�ǝ��+�m��&�e� �d� �l X`m�� z�΢��3/i��cVgak��+vlIe�c-u�3Vi�`M�el�M��L�Qή��j��Ʋ�ʵwK�m�jD�Kl�75��6I��j�wY\�\d#�2m�b�Z�%���D.�iv,�mp)���AӠh�+�[�Y��:̷=+)�<��*w�)��oeY��t%�Lb�ѴsE�K�����Z;m��X-�(���߼0|��1�]~������lWD��z�2�m pj�V�{:�*��zx��M���Sg�i$ڶ�i]��H��N��.�Ӡf"�A��l$�^w}.�NG!*tm�Zf�gu t��5V�W�eÓ�kۢ*G��M�W��/-w�x}�O��X3v���Ov��<hD遼���yIo����WQ+�;Rm8m�ӋƯY\��DMӢ���n�+8U����r}p�jڱS�#���b�}8�GD=����^n�TXL6�<y���Wr��~����eګ�Q���]`ו��=�ѻo��&0t���'��	6��Z���C����]����}j�ne���1ĳ2��:0�"�R�}ЧZ'��9�F�$�ʄ)YN�2��+sBQq{��$n�:�J�&�v�=�U�'Cu���7|p@+�M��]n��jiH�zvr���'Z`��L��f7񫱎hMpY��[{X6Թ֕EYlgI�z��Y��v#y,���	�s�h�z#.��#�[��D4�{��x/e'����[���GK�"��t[�r�z��]u>���5*c�_9�$�n��qg��
�B�I|��ǅ�=��	�GE��C�rʁ�)⮝�'8'
�uV�j��1�,�G��.-~��Ug�\>[Soۏ;���ý�sW.����X�+A�W{�����(C0�"��6+��k������<������i��o�{Ʀ��~��bd��w&�>�W����T�	ƚ�W7�''��詀8C�b�T�!��.T ��%$�$AN5����٭����)��JBPY�5{�)��EI�;۰�ю�L17ԩ_	��N�������)���0��HRW3�� f�ՋW36���;
�P���5�fߜ�%!����Y�wT��9�WP�(}�(=E֛˃�[�n�M�==�j�}4OB��O���\�2�M[h���9&��������g��]�hSPp��}m�p�u�+wE�+�
�/�҉�=���n�V�Z#v�uͻ�q2�3�����w/n�g���Y>��	罛5]�GTq�R�7`f��d ��͙-&��G^=S��=���������d�A[~E�vi�d��{ჸ��O��F��k����ԑe�e��`�anU�Y=�wOV�tV�?�-��m���*�hX��<�43aA��A�i�0����WL��'�16����%(�SZT�7ydhULU����a�M:uޫ��|��� �����3ܢz����+�M��ݲ�wK�_Hۊ�!�r���N���e��(�7DuXo<��O2�#��O$b��V�}���[k �U���;�猻��ӈMd]o��@�C�>n��Ҁ/���{�I��oP�Ƚ�v(t�u����)�e��ltj��X�1"��o^[�u�<�rψC��AkDW�\���u��ǥ��}�;S-���Ϩ��7�YMi��O��H_�ؕ�oR}�
x��y˘]t��x�@Te�ٝOt��jzh=����#dJ�xm�ȯ�fL���+n�ƠI�k�Mstcu��.�cz�����p�h�$�Ѓw���G�Zـkw�v�2g�X+��֜��6f��*};K*�{�.	D��I�%^��98]Z�.�����Cs�p�b�R���z/y�~w��j/.��ʾ[񃩁D�Ld���F�S����@����a�t&k]�[��;�xu�y���~��FȄ&m��O5b���nA6ɉyx^`�mޓt�ng�=K�E7�_M�b�o�u˦\f�h��nv��tW_ְw[�{j�^�
�{��0�p[������:~|��88 	4������- �� [@ �ͷk��Y�Ӧ�Ks�ܐ�,�چz��[3�,��.�+4�K�"�֌���ez�$�Y��-h`�֚8�Yu��-���iZ�C[e��֠9�\����m͹�&�%&&�\��m�mk�&nS�vXY��a�3��A}�ӕ�^t�����\_Ne�#�bMu��`&�	�5�E^���kfn5�����y��E;�"����(��w���e*IH��xi�j'�-����m�n6��WT����pSގ2��;*h4SIQ��s�:/KE�]�n�v����A�~=��n�M������V��츲P�w���8��U���t^*n
!�f��1s2gQR&ޓ�����䆣y��A�����U�y�6��]�8	�j��g!�I��aL��YIj�0/}������s�]��2��G��c����㺡y�[���%4a��}�$�b����i���GgGy}n�tp��86����9 %5h�\��I�+��y��@6(u5^��^��ty.gC����$���ƦaR�ƻ�Q���7<_$}���`v�qf �����D�#�{�ۮ�,'j�Vt�ʿޯO�wp.$-\�y=Uw�S(6�i=��W�3&CbI�ّ}���l���@�[�Ṷ�f�f��j\�x�b�k������{��<�J�w�ٚ�����Do:���}qp�s���#�N@��ʇ��!,�3;�?F��ɯ�x�7�f�A�y��)�oU�����D>�vz�.{�&[6�z-�<�N�Y��A���^��ju����2���v{�xv:z����绣hs5����3pz�Ot�H
**@G����n-�B�Q���͊�}��8LRs|r�L6rR���/�;O�ܪ�;� r%CI��4:��n���Ǹ8��
���.�sGgu��-����¬;]u�\Ne[��ʯ��7�2�- �ޝ������{��̋�L敩�����tgk��kf�:ζ-oc�� " $�l�m�@���iݨ�մ���a�]n�Io����U�ӦVX��@��߲��-Z�I��e3�p	�N��5���R����UYF�w2�M��i�F�T��5��Xף�+º��L����4\3'atY�o4mj駏�}��,8)�_z�ۭ��:�����w����������{��^���{;�=�S3|�$�-"��0`5��W7�p#�K��1m�u��V����1`��;�����6T�_MNJ�v�wi�+�ow�rPy��l�Gw8f��k˿|�=�\�^�A��Y���ݞ5�h����2����ש��tJ�}廝<Y-i%N����%O�߬I߿����~����mk��ZK]*l̎6�\h���6u�T���<󷈚�TX��sV�p�\)+�����²X��f�u=7E:�C,���DX7�f���}�3n�8
���Y�״���U�ZG�'u��1�ù a���\N���LB׃a�s��Ջq�me-���@�TWl���F�����u郛"f�"GYP|w���xQ�ɑ��%��W81ղ��.�;�l��N_g�!�T
��h�*�/:U�u���W9�}=4fO��tm�03����8}{�������AӅ	��B(�eoT�\<�}ON��g��,g���J�!o��
�>�^�}���r�8oj�SFe�/��r+��ɵ7{V゜�4D���m$�c�	�5mMa5J��һY��7�n�RC M�ў�8��赽�s�����O�W>y֢���V*��2�]�=�[sS�/	�ngM4T�v�.���}� ���{b����S{b�T#��$���eU�lF������e�No��R3��y��"c�}��@��c_v�3��9��C<�E��u�Ա�i�n_v�����l�FD�3E���+������ha�4�J�L��^���*�눍�YF&3%��utE������۷m� �*�.�yd\ m�@ l��v�[t��1+��9�#�b\�Kf�Qi]��FYi���ԺG&��`���vPnclPH�Y�i�,K�z����-a����˳�RR%]z�1e`$���̣n٬Z�E`�3\D�[V�Z�d�i�b�mzG\����8�_��o`�f�60��D��7j7������o.�b-ڷ�K��h=�^��t��|��%*�gt	ItJ�{�N�K`0j��\f!��z�L�P�m�I���m���[n��=��X�bՋ�즡 l�&��n�T�E^i�;��=�y��2N7�n��e�=3\����e�I�S�U319�h�(ѷO��o:w��Yy�U��LU�{ޙ��*�g��T��${��ˮhAg=�f3�jjʫ������U.���Ҍ�ɣӂ��������ͨ�Q��	�f/�1m .\�M��c3jn�¢���,@�b���TP�7����뮿X���a!��P�E�YZ���=��[y�CA�@��'���Jb�����~���~���fUԬ��B�7Qڦ���xo�˭�KX�j�Y�8o]fu.��%�y`�5�E�p�ަ�t9�u����Pv�cPk�J���h��S�*N=�m��܊ŭXB9�{��7Ym]ػǯ~2�bwf����NM����9������f�6�'|�c���>s2-T�n�b�ckj��)�*��r�����3Z�@�f��]���⺹W�mo��WWS� �Ε�E��c��-��-:���^����n7O��@D��`�F,z���:���9j�#��o��|�:ˇ���`4�Wy�v�]d��ۚ.��]_,R���U��ܕ,̝%�yGp�n�4�+���������T��]E�+ 6j�:��&]5E=F�kL�C�K7�.޽�,Rܽ��rѽ�W����\��v�*{`�v;338�w�nNx�f�e�-�8��Ks���0�\IT������P�S=Z���x���1W�+2�Լ�kc7+(��m��m��m�f�iK@         m�^��    �E��"� H�j���n�����+      ml�ٶ�  �  j��       ��l �-�   m�     ��Y�5R���) ��ó4Vւ����-v��qu���el�@aWj�.`2ƕ4��eh���4�ql�\gݥQ-n�"��k��� �j��,�k���2����.fҒ$�:宎����:�ׂ%l8J\%u�[Y�38��m�Z��7M&[YKv��.�6�vۇc�-���7Y��V�A�n�˦v�v��/,+fݸ2�n��s)-�q�XItT�3M5	V��W1����P[D�Y��\]��Y��s��;jv�u)�v�4,�Iu%M����j��[�i��-�vwє�l�\�hn���jMMH���j�c�W�2��Җ���Z���J�)��k�Ys��sc�-��t�pĭ��[7kŶ̮F\:�&�j�um`P�n�:el��Sb䴦crY�4�5���A��B�ʦm���m6��c�jK���ie�!m��`�t1fB�4��XX�S
�\J���4Kf�l֖��՘����4���̠��$tK.q��fፘt��Y�a��.KC¤�6�j�-�Х��m��&2Z]F#� b3e^��Y7`����Զ��Z���A�iw^��gF�M*�J�S7^�;����	Lh�6� ���s����[)-0]��ͻLHX^��i�P�{:�<�����?�������&'�s�}���v�͔�$��7t��,��2��z��뵺�m�nT�)��%I͇R+[����M.�iI����}���٘Rvi��"�n�C��wH)ƕ���!�d�+Y��]p�~�����
��'6�X}ף޳�����5J��9�m��װJ��NqS���n����F[�hOt.q��/�5���^����J���)��=��Se0�I�qqFp"�\�;���s��c���f��W��e!ϑy��Ew�兺�o�� �7`�rd��Ponm�[S��p/;�^r�#�SjgW<��;���!Y��E�Q�\�*�PE��\�tu\V�;7h��\D*�{��[���2Qi��u��;ͤ�%��-�6ih���
-�C�ǯ�����S<#7:3�(!����gawT`�xC��Ta�Z��X6J�)E.��oV����	WoqHWU��ޛ��V﷿1ίߡ4mz���P<�nndW[n�����=�6�g}��{�mE��"s�sݽ���tr3N��h�I�s(����R����5Q}�j�ؒd����z��t_yd�Z%7G�x^�̍R햳�l����s���r�j1j_I�ɽY��d󢽓�3��V�O̯p�6"uUs�x�o��,uon����	��L��nN���}�x��jo{;pn!�k�k���\^����G�s�'l�H��3�g��cv�wpՁh����m��l]'"M�;[�S�g^$�;q�Z�u�l����p�|��]R�{�چV7��e�{�T>ǽ٪ĉ�S1ۺ	;�t����7�x���.��fo=�a��������:����L���{���l2�&5��P�xy����W��(s��p���}�=�a�������]]���"+Yx^�.:��6���۳�*f��*��������}���N<!���=�oݢ�s��C���M�dF�b��������V���'ƴg������<���p�B��5<�O:��E�a�p[ ��b,a C�pqWE���{k�w���:Ņ���Ri��{"�m	��鞎�:�}�%0Jh]��q����`/X&lwt$�I�II�)�Ћ��]5�F���M6�;]ʆHq�/x�-d^^�n����oZC�)���|��2���+��h0�7�*�?3�:/ע��|�.��u�9ggj������薔�ϜOu��vG8:�f�N���t+ۻv��g�ے��[���U��w���Tq��s�f7�qQ��`Oj��==�0�7 ��w*�Z��-�gy�ꆎ�f��ٗi3+sj�J܅�\ʷ��8���+�^���vв+����h��Ϻe�m��T~�m�6 e�k�w� &�  ��` ڦ�H�k�fYN]z���ZRP�]uR��{�b�YB�S�^��ٺ��Wt�׵ugX��=p�;l�9�kvtt[�:��ͮ]m�I��p�Q\Jy��$Y��ۤ���z+�aԅ�e�й��:��e�Q- a�a��n!���]�[�&��x��S�ɒ�m�S���&]�S��K:8GnѸ}�JSgx�k��~�kދj	^Tr ���`^U��}}=|�t�S�����6��\;:��y��2�_8�w��p�T RF8��d��"eSk�j2��;��ݨe6�0J������C���Z���(]��fbz����t-rV�Ջ״y`-2��:;t�#��s��i�ǶE�!C1|f&����p�K�pGV��^nv�o.��f�!��hw���ї���=�����=��V0z�H���K�k�޲r��M��z	�k/��Ws������.�\;ޣXw6mW쪧�ڵ5�a�m{�U�a�T���Df����{�Y��ȇ�k��&WY���L
�^tT�����}���(���:�k!u�X�՗�I����
���]c����'�K��츝��{K����)�-�S�:��fm���e�!hL+S	$��ZNػ�1i6�ukMk��X�/Ȕ���C���Df�s��R�+�Ξ6,��^��Ӽ_^w&�N�� ���p��|{�r�$����7s;�db��������Y��z�a�K���s?;�ӡ��}wu�.���,�s�����z�V��R:Dr���;�\�@�b�a�7N1޿@u�ޫ��+��z�q���ԬHg0t��=1��'�����!��4�.�����G��o��X���W^ֶxʿ�����eN��s[��b��Rϳ��Y�/ p�
�!�Zt�gr�$���"�l��	$�L��z�iv���1�2�&��Bʫ��e2˄`iWݷw�]@��\ͮ�Tj�lI���n.�h�����Q�`�Bж�#7�V�6�BY9��fe�#_f7�q�}�����kӨYI�M��%ի9}��`ґƺ���B�[�5ߧ�o�{���o*���ݗ7�:�%8C��
���M� ��MY��9�j�C�췽r�+�M�c_1vl�5��.��0J`A׆$"c��P�Q�ٳ���˼=H��|9ܷ��|��~o��ݓ�%5��#ɖ)E�1����ֽz�Q�c���@�γq�%͛ܞ���ظ,�o8w��i���{�12	�e��.���-'
����&%�t�߼.F�ݺX�f�N9��4��ek���220�����­o��6J뺎�_[�N�OH�9P���u���E)��lE�0�i=���˦��}��Q�ݮ�x
z7;�~�]�Ϻ�:�b<����:�!�):>~wݹ��Bg7����up"R����vWw*:���P4-��L�'3i7I�ޫ���%��/�4�P�;���ɝ�^��e�_���:�艝k{8���$���;4�D�����mӸ�1���(Q��������y�0^�	�Pe�{s]���DNK�ĭ�N9���O�^b=�]��C&�:�uu���T��d0�>>>�s=���.�U�s��$�L$�	�m�rS���ou��1^��0�	`4���`('�x���n$���1��������{ڄ�~V���p�����̀������S�z̝��s���Giո����CV�I��؎v=ʙ�a&�l%]~��j��q�o�x�_�G��򚟽\�V�?1{�fg=ީ�;U�p���	��n���>��1P����:W��OC殂pIr�Yofm��뱕}U��٠hU��u�N��������8H @��" � *m��� :�ʺ.�Z��hh�x#��e�Kݴq�G��'%�{V�e���YX�������$kV�e5Bb�l�& V�J�^h��6�;�Zk��3j�Q��e�˂F��˳G[vk-9��ـjk�5�-��; �Cbs�{$em����Z��`i�R7F� ���I�1�`�V��ՠ��]��=�&����y�;h���o��K���>9���`�� �ky�a�wW8vV�Nv��فCM���I�Ziܕe��9%3�����H2h��*$+�g��Uǹ:��P���x�=�[E���w�3
�3O�!R!�I���Clޚ=]
�8<�4�1� W!���a���kV��ů�M���Ra8n���-Uļ֢����JV.$���b�K�^{;ǖ.�t/qo}p}WG�SI(0Si�0i����G�7�λ^��ê��;Hu�ݕ���)]�S���eᤧ��o��v�m^���}n�,�@��b�㧎�`�w�1L��c��:�6���+�f(1�;i�m�}����sH�ЩV�]vG|�ۓV��j��A�M'�_�3�<�-��n����'�%��c����5ޥ�����w�Cv�v[�ڦ�V].+�SYN��x�۽��2�y�'���@O��֭�(t�{�K�N{7�H�D��-S~p�%��z�����%x�p���vla۞
����8���pÆ�)[��3UOY�3{��^�+ǽ��|_{=�dc�*LŽ�~;�(�s��a��t�3]�j��d�w^�zJ@2�;�z�ܬ���(ۥ}Y2�����$d���.�_A��pu�k7����C8�y;�����te*��οfh��[��)�3`-����;M4��a��������B>��+`�6���ۮ��i �L�N&�ݝr�V�1���E�7[u�Q{���9��԰载5䈝^Źfǌ��vl_f<��kVc�h �K��vw �Iq�L�%�;��ҡ�J�L&�:o#w�Pe�)�novJ{���}P�z�g���=�dv%�2�m�(h��pk4����g[%Áө�s:n���ե�@��{���֫��õG��F��V!�/�/�=�辽�9s�Jh()2�[�����7Q/o����vD>�5�et����|{aA{wki�h"źؓp���V��7�=S�uOr
��e����Q�f�Ee��T��6;��p���-�aݦBRȻ�*j;���`4�-&ۆ�p�T�MSa��sT��Y�\�lR��H�Hɼ�U������#��Kr`�Ʈg�M�r��C�K�Suض�2���k�%�y���94=ϰ�.Ge����R:��GB�������r��c�"�z�k7@�:ӎ^�=��uӋ �6�� �Y�6j�Y&&	�/f&4ʒR M��e��T�)ǁ�h��<�Y�e���L�:��}�^����9Z���*e���>�s���^;�^	yW�E�V��QD�Kj���W�%�ҨEm�Í�hø�n�os���/zƬ��ض�2��M���e��������*Ⲏ�sz�E��2�]{�;��������4�n%��[�H�y%��h9�2mP�R�{7%�g�|�pv^u^8�Hڬw]W�s�9W�ܮ�U&9�r�I�&���K�7嫥dڳ�mU�&X��X��v� te�]
yd�F4@��{��g�9�b���Y�oT�gya�4���$��Hk�\�e<�J=ݤ�XP�E���3z�$K�rmu��yi�R�5���:�#����P�I��r,9]�Y����;�R�uWMSir���3H<X��]�Vr��W �2�� �����������nT����3`^e��|?����d�uW?�*��_��K�sg���\�˔��,�%��*NE�����2��ҵ߆��H�g9^Iˣ��	�^>]��g��ej��=�ǪdN�iMQ)���[�p����ڋ���E=C�>o�3	ܽ�oS��WiZjh]�o{6a�[3��n4zO(�[)��!F��W
���v���1���v�l:���Ln,I�`Bi!�*fLɈA�\
�~w������2S�������bDb���7.��'���0�a0�=���wF�Ň.X{k^f�ȑ�7��ҏ���Ez�x;+�/K��4��qc�)9n}�ܛ���\QƖ`:_��7~�fv��Z0���2����4�8mߩ	�F�Эg͍/g$r��N����T��;�IAl.�gbuP�E�x�m{��(u�kf���Y{�K�*�\N�k73j��b�{i��Bꛚ�9�h��u�Krn�ՒTۄB)�� ����.z��v�� [[lm���wl�u��%���m�V��M��Ѷ;K�&�`(�p�ه96uK^�t�s�7l�t�&]t�m.bBj+��cJJ�2�@�³D�ukI�5�n��۴�8��4`��i� un��e]ڭ�0ڬ���	$��5�c���8�b��g���<q�=<+�=���T�����;c�Bb@�*���[�5q�۩�ǌ�� XM�e���Q�F�kla^/��⬜{|lfJ^F��j�MHLU�����n$��JHY�MU����Q�����o�O��fuh�`��/��un�V[�5��6HҺ˥����wGzb��L���{ĺ����X,[�k������Vb��7�6�(M��G�u���f:Nk��}g���*ap$mTv4#~~�UO�;Luf}&�z�8:6��*w��E�
-��_���TݯU�ªo	�]>�I��l;�b��B�֝t�1�9�t�z;��������e
���%C.
e��W��/w�)��V�i���JD_������5��ʉ�C�4J+7��>d('������8I����bj������F��|P�_������]�'iϹS�p���K�y�q����oƁ{�f���(	p�Ҋ��̮�v.��:/&�Fc��W_���]m'�8��g���kW2J]�N	OP��=G�����~������ ���l�m�n��%�r�חtڭٺv�ئA$������}ܘ��(( w�.cCǇOR�c�&n����l��`�UU��{��� �åҮ0���'(���]x&G��� _u��_�u����E�|�Q�Dg(�/vԁpX�I��߼�g�!���sa�%�W����w'Z4A��%�|@/4%A /}Z��gx؏2w')��8lF����b�O���]���	0��	���C�k�f�ޱ�n>Y���䤹Bq�n�J*z^۝C�*�񅽂�ζWi�8��ٝ�r6S���-�/B���ad��].�l�����xvv�q`�D^�V����]^U��Y�\�%���Z��j�\Am��2܁�|+�Iw�.舑;�����1IM&��Z�f�c�/Ky7f�yҦ�|Sa�H����"ۂR��}£�G��[��=�tsL5#��T��A0{����b���OŖ���~<\��y+KtְE�cy����~��N��n�0�L�ӓFԧΟ�n�'�G#�}uRI��z|�)���NS����gt;ʼ�*���/����(;�a4\B-�U�5��t��f�S�����>��}���k��=.��!��/�j;E�e��"������zW��{�no�5�!��.7�E��g]]ȡH���MJ���b�{^,`�ޞ��8]{8:WwvZ^t���I�J���M0�4 T?������K�w$�{�@�'���뼝�o6G�m�c�h�$�*�Th�E��uK��)h-d7Ү3L/]���NEx����I��M��~� &����O^�����&KP��f�b���[@G���Ō��+��m���>Lz���F� ^G�i�����lAa��"�I��tt� k[��G)��Ø0�4�P�B��7��4TRǀ�<����c��͵8Md�^N*�)�}{��Ge>��L��B�[��)^� �;y{��*���K�r��B=Z�b�T�:��z��#�9��M ȵ�1>ʰld��-�ǉ0�)8�׌M�\�/<IA)��]ǔL���}������� ��o.��˯Ls�ݲH�dw�)���|j%C�9�ړgڎ{X���MY��)��4�u�601����T>�2r>��Q�cÓ�9�EcT%����=	"@P����*�!1i`4�~ݸ�� �žSm`��0qv4i\iTu�h� �4�e(	�b9{��S�z�S�p��4�$ԝ��P�W��C�O^�z��fS��$��
=>��ކ'��Wr3���n7i����b��+G=��tgM p"wW�����0[��˓��뇓Q.xlO|638G�ܦ�I��|^�SX�y}u��Pvج�O:��&�&�G����!�r���כ��!0�G,8�2��ܹ�Vzk�3&��S��#�� S"n�4��g0��CoMfpSE�60��HW	v/w�UZ�\yɔ1sn�A`m�m��"˹� �� H �  W&A��Lݝ4�8`6&J�髬Fb��Cf��� �d�k�S]�
�k��9�+�klۘ�A�iC��֪Kp��q
!u.ѣ�S�v��� �і��ɵ���7���Q������Xj9
]�g�V/h�����v����
���1⧳x�B�Yh&ش=�烦+��c�+�>����W#��cx�|��CW��E�{w�~7�+x`ʝO����N�߽7-�2��L	(w��C<<�n���4S1�ݷ�f$\�m��aL	��ͭ��1˭�v��uVbB(�:7wx��p�g�����<���}�͊�����{���	U3�\��p��[f@�V<���E�����r��=���%�5G3x���V՘1���S�R<+ɭ�༸"��Nr���znʛW9�Ϡ~D����<����3G�q��S��=�)�*������WNxж7����i��26j1#�AnN���ǀ�v� h����w�z)Eg�n|�� �~k�\�3�D�Yޙo�qsN_˅�#�݇k}�g��NmW�#���N�^�4��P�>w�p������T��
��ԷR��l�����9S�fh�Q�C�r�Bl��thc����n���Y��x���[�gyr%	�	F 4��W��I ďoE��J��fҤ
$�n
�2ʆ@���r�ťa2u��՚��d���7��9A��D��{�B|�p��T�v����#�W�_�k׽Ĥ0�<yD�w��k���~8=�93Fã�tT7v
μM�>�x����^.���nkۘ����|�a�D��)�Tr��F�qT�"�-�+yBژ��wA�+g���P|��~�>]މ`z�<�B}˦y��q�,��%Q��PC���R}���k�jy�#T�4�(w��B�� 1�O
x���<NO��>��m �ihMS#�򋋧>�>�ɞ\΄�{NU�ھ��� �pf0�b5%L�+�2 �C�b����D��7}�y&������]ixnO'B���;<�A$��I��A��&�t��F;�݈�jb0�e���A�#��63Ń8�ܻ�iB<*s)sq[�ų��ǐ�U�o���n27-+�M�h��7=��F�%��+e[<}s��}'��e2�a%�X�ˆ	���c�r�,�Xj8��K$�ј���r�l��^�6xW�x��0h�o�����x��&7�r�������k뮣׽)1��h��H��쩜�`��,Mc�ˡm�wV=�qFIНs�%�̹50D���h�stl�Ԡ�{�|s>��쉑x�,s�]v���m_�h<�zY������r��l0`��~7C&�4�!v�ڕ��OS�_�y�������t���EϞ���vU���^��A�K��Nf6o�<g�O�wHP[J`�a��Rǥ�B.��1) P��Wm���ΉͲ���5��`�00�HD8m�>,��is#esbI�R�S��A�f��L���^Ĉ�H�坹Uz�W��B%�	�!\wyVf���^-��t)i�@|�{�b�y�e "t���L��Ǝ�A��f�#8�-�Bǐ���G��a�� "����yQ�ؼ
7�X�4UdJ�+��O^����P�Y*�A�)gL�����(?=�cݱ,^�#Vm�-zcc|�,-Gӱ\�>^fS]��WB&��ؐ��9[�!���y�$Ҽ�fչv�𬧝ÄZB�xq�KR!��wIϷ�0H��c�eׯ�k��a�_��5�{k*=�¬�ۯ&&���ד���r�J�hz�a��Z.=N��ꦘ��Ǹ��:n=�=�,�MH;�A�K��/6c��a`����}uV���M���_;��ϛ3v�����*K͸ �L�h��p-"�������͢�R�;�6��8SQբެ��?*S�i�ww���ާ��
m	��.+�t-�)�Z�^��.��F=Ǉ:v�bf����Ȯ�هܚ;5�a�l�:�x�\ �d%O&EM�M����ȱ����l�ݨ�q��#�w^s���:�p��5�-��h�6�p�z���w��P�6�m�1�B>W�Ow*J������j��wLT�\w'm���?$yH�M�Ӊop�ϗJv�����5b���r�4�d������1�Z�|�ߣ�� �7��˫\�a� m� �Igv�\Z�rw.&��,�
�-.�&h�m	hM�����iK��"B޶��H�z�bM	sR�̮��l�Z�r�8��敼���2����t�B�az���b�@/+k�*�]�Y4����kf�Z��E+�=�H���œ��O^p��(
X�i:�O'�0�4Xd�q�ztz�5���Җܮ�՛�%Fx�4��&B��`�I�ě������%&'�i����ܡ6�S
@�b�����P�*�4=����3χ�͂e�.�[D5���$k���0�[fw)b�1	�#���R `�ީcs�����雠+M����]_Z�2k�ts�i8P�*cʝ�y�p��v��zX�p���oV�U�8g���Cj|���B�^��;=�ȓ0�A8E尸�p�fsuf�N��;�1ف�*����oM�<{���bj�ۯq�+<�ݱ�ғ-Cp�t�x���n��8/M]e�'���f�/����|�M��!w$��!�:U���UC�=#{�(��I���~C�5Y���3E��x�F�OK������^]\뙳����V����k��s���0<zl�gZ3]�ڻ�Cd]XsQ�L7�v��(�xK|T]�G�>�f���kX;z�,e3�dRٰ0+^�6������a�k/F�p���� ^���M�Oz@l�U>�����{^�Z��n��p4p��@���e�Nq��񌰉}���\�`TY����8�׳f��X��w ܗ�uz��2�|�3�"˹gr�7u 9S��ΟI�t^���)�]�XwU���Z%v]�w�q)e.&��O���dP	ăd��ۙ��k�9���n�����`�s��ԴEg���}�z��Uy��ݙ�w�W��z �'
G9M����k^n��f�;;s��u�n;��`�(l0}��	"K'�%m��U7}y�:��Y��v;��t���6q����[�;����j��d�8��͌��k�:$T���:� ��N&�ݺ��@L�c]�/1��Yo.��8����({��שn]�����Vu���+l���Vi{2A���є�y�h�o� ���7knɶ� m�  �   �gmՀ   ��n)KV. �M��X��t�R��n��      ��wM�       k�-��       V�l ��  �6Ͱ     i۴F��7:�Y=�RXe�ަ4f����[ ��Kc��ۋY��w-�C����[�&�O�fM��������Ɩ���n�:7fݹa�2�	z�2��V�^hæ0FMmīe�m�t�0mɲ�l�'T�[�CSr�[aq�k��-ĭ.4��:����6VI��H��GJnt��%��])�Z���m1	��u�z��i����s��+�R���[��`���g0��i�b.��k�b:m�X�[JcM[�H�f��]6�d��tm3ƍ�[��ƚ۳�e�ےf:����1�n�;;Hl�M�y�s�-�b�tlpU���.4�g�-�;-�����.;jDV���G6�P�8�V�76M]K	�)�X4�:R�4Y�ST�k�F��HǛR�ۦi2�.Zp�R�F�m�Ŏ,��Kje̥�Y\�5�v(�ci-�zљ���\�6�
0 (k��14Ah�&+�]�k�f�iÂ�s�C2�b[Sn�L�]�,d�X��2�\�!u6�3*�ke�q5Q�1%�2�Km����h�$SC��Y�ڸmy[�L�i�C7;pG[:i�s	i{r\�i֝	μ�ï$n�[9y��t��tْ�:�5�W\vٗ,�&�ӛv��|��^��Y�ɜjƕ��Ya�lv��i.l�t�[�}}���;�{�?w�q� ,ȟ�	��^x��a�l��C�Z|�C��Z:sՐH[	�(6�J�%msIeja��e�SM�l�M��K��2�~��~~~qw�[n��Q�4�_�z�������W�m��`by,*l;���`(e��.)��v�U�$�����ըA���p'P�{��&~��1`���G�^(|���*�����0��ȘN
n;#Ok�l�-�Ax���k�Åv�,����G��h�v_���B�������Sn/7U���:��r�8r�n�'�p��T����(XZlv�p�~�gOW������~��<.4��}.�4�6�Q�ԙ��I^0j	�q1�����m��v�bz���G�w�yWt���q���̧=h��f���~�^�C���F�gV�w)z��T�����ՔY����T0�-4_�C�����K�m�e��e�БW^�"_�4�)��7�
]�~��~�rO��;�|}��V�x��i��'���t��	�BDXۋ��&it�Nb"�9�jgn�X͝��5Mב������:��cLfBj/S�ɢã�=�p6o˼�:˜�Q���Q�xжm��[�Z�R�{-Fħ�䬦��`/6����^��J	�h,"�?��^��y����BgS�k��FaM����ln�ö4����K�ǳ=�v�ו�7z�#��.��Ց� �0~%�q�V���j'{���3' 0ö��]��Q��0{��B�If.����(]G���rq������'������-]�(�s�{u 7���X<U�ݮ�1VP��B�4ߴ?L3'���6�)���͇�F����۫��9��M��-�z�_���V�˷`�b=����u|�ǵ�-:ݶ��&�"�]v{K�ժŸ%����|K�<��,3O�^Zkl�B��34��I�>��W,���t/sE�a��E�/D�Σ7֦�ќ���^��B����GgC�;�i-�<�GH�z������dW��c�Oo"�	2�-�y@r��;��I������"����.qV�`v�#�3�e�N�Z7���ٺ4�Slw1]b�~�79��<dP~}�lx*>���O��{�U���(.�j�{_�J�,g�I�W���c3ܹ����K	+�zx	'oZ/�"�},O�����mu&������x2<({O1e-��8zy��C�	�kz�U�כh#�׷Nχ�Q�z�[��4o<*�o�8�2{	T3{���i_]�,NܨO��Ն�o��!�%1e��*��Ӹ��li!�[�1� m��m������m��Z\L��:�r8AP���-��(��!ݞ�><f�����"�#�a�h�| �2���y���=�M�¢٬����^�~�(C5�U�W)R��앦�^eH�F��z<��~�',���c�4��E�X�-��SlNR}��Y�PpiɆ8y��7���UQ=J[�V�﫲N��o�'��θ��ŎE����c�}��5��B
mB�.29<$��<���E�����W���2t�J�btm��'?���2���!v�On&W�0u�2����K�-V�eŧ �D-�W�n�o�k5� [d �[�ľ��6�� [[lm�T�NۧE��n�-ї�-�� �b��M��mJX�b܋min`�кi
�1iL� p�b����Kf�Ue�;iq�� ����3i�qX\;LjV��B�,I�K�E�����`E��M5�b���4k0)��8#�1�t�ǅ������Щڭ4;��J99�"#=	4��e��;x^�����%)��܀S���&Ϛ\�)'��d�wq��ϭ���c��%�u�����a8�^yuͰ�V\��{N=�H�G$�I�I����u�5�KZ-&�8�|���Hڻ�s�V�y3:,0�^��������l��~�!�O�m^�˒��ov�â�|/9e{�0x���j���=fo�o7:�LOÆ� �V�S�6�{�AI7�-��cY5u�z0�&:�/���,Ub�u��V0x^�=s�!Ӻ+���k����j)��!�_I�1Zp	�M�,{<��O�&<�̯�Чcl��Z���nL[�'h;�2X�UvX�M�p�x���h�w�p��f��=��5t8X���k��Z�ʖ=��l���ݨWJu6�F��ܷr�;Eem�[IϵE�����7��d��d��1�iL�=�M Ϗm'�~S����	�K�����v�g+[�G�������̀�}��bl�v�����v��
饣I]D>����jP���w*���~�&ǆ��~5J~���C|Ѯ�|9��8m���E������ȇfF�r����ǽ���f�p�1�d`kv��zf��Y^����ۭBnE4�������hn�/Fv�
y��:�d ��.��g���n��3�T��RS�~[K�Ǽn	��Gp�м��n�<hh۹�4�z��y&9d�`eI���ǄOo'6��sb+�Msq[���uw��ɖa�	r���c��_�]z�B���3y��H��tڃ�w5�b���:��QU-��I���g�7۪9��L�S�dz�Q�qN�`p׼����G\O���i��m��A@&Q��8�є���uF��$��Gy���A��;�5?�2+Kd�*�No�"Ҵ�舩D�;�����<�}Mi�WR�^/�Z�G�Z���;U3W���A����Cg��3*����ɶ�����OSG��ȩ�F�n�ev9����G.���C�|o5^t���vc���
S�=U�NvƸd�8KΣT^9Y!�To���hzv���Z�4XD#ἅl�H�τ{��nN��h�p:<��ߧ���JL����&@�2������~鷵e���2� s�.�3��g��ޜN'����}޹~��f���a&�DE��'��F�,��M<��W8O"졄�����ّ�d�#w6�p�N��������,�	t��U��qD&�-60��,0b�	�)�;�iY'&I�ͦWli[���S&H�[����0�d����,Aa�z��=*�F�G�ݹyM�e�����6qΧ�HyDƇ/�t����|K,��6��y$��^d��<�3�&�}����}�󨤯���f\�����#�{y�s<�X�o�>���@��P��^�����Ļx���{+]&�Yk�s
��R��Y+Z"n��gl�[u�Զ�3��"6��u��'�g���|�W�� �S��gɏO��T����/&eGm��e3���i�m�y��2N؏���T�MVi�L+h=����{�늓DϽ�:��h�c��M�)=�[��m��뾰�����ɠ~f�h��ۍ�V)S<5�Z�0B��󞑄C��ʳ����������q�_�t�S)���N��g8�&lW�����<W��)��m��_�+V�tr,��R���cM&����d�������F�*���`�ï&�=6��I�����kz�[�ow����F=M��Ƣ�i�ep"G��O�8���%��ܯ��W��8��q����=������n��w�l�pڸ�=�����f��̚�T-��~O����w�V2(y���G(��ǊL�2"n��V��E���>���0+|���:IFo�'H��n�ss��(���v~#+,�v�Y-���9�n�a�������	��VԴ1,�陮�l�`�-�s� -��Z�l  [.�oe�4�$�&�k+u���179�ˠ���cS3:&�[���%L�i�]鳫ّ}�hk����U�gM41r�l+���Z�hA,#HVee�I[�ˊ�$���f葴%#��󖚶,|ӄ�h��nNtѱf�oOL��W��p�,`���_{ÈL��h�U27IC�{���SV{���/\ҋ:D��>k�Q,�lS������{E���e��z�)�HJ�h(.�Mx���xݘ�����Gz��_Q�����>v�6�]�n�ZyѪ���썖����ћ�&�����v��}E���ug�VS�T������V�8w��k}�з�j�����?��P�]�sr�����R��O�0��eݡ3�=�;�(�Ah���]R/�3��ꛯP������p�p釫�2R�`�]�v�bTk �4�]��v��:nPl[���W�0���_�/x��`���܄H\g�̦r7�������Q��slR�x=i뮖=�;�k�{����#���h�6#�m맢�³�c�rm|�dw��U�幢Z3�]}�R��{:ʑ>1q{	G���t�z�{d�O���1tɣr�T��� �gb����a�&VΙq��P��+yi��
���$��ç�T����A�B!�����s�{U���>ԥ��,Eæcz�<��d�`�*�`��5��hU�`|�8	��Pv=y��H�9��5�E��P�{�fzEt���:�4���Ⱦ�^�i�xz=�&�a��F+K�2�x��i���m�E]��ǆ��r�\Q9[.���di����U�G�a�7~�f�l0�n��O����U�]���}��G�������]�Fk��<�|�(��9�=�^"�|w9Ψ���LB	��0#	g�n�8�4����w�T��w4l����׼�1y��݃^f�)�H�#G��⛦�>[�fDLTPʁ���n��X�����H
�������863l��-�剂:��uV�ѻC��wM��"`&�j\=�y��e��2���{��U�|$�GF�fM��,NU`�S- �����l�ynҥv�m�b
��@e��-C&v���Q�xh�m���|0n(ꍪ{ob�H�٧�|�Q���!P���b6��5�+g�2�uwn��FT��4��7ko���	\���g\	��
�e��8��1�!�v0���sc7�������83�>�+��+3[㣻��4p�~|_�ՙ���mCP���}q�r��>�n/�_�i�ƇYι�C}ISɘK�ފ^�����<e_������Kp/�m�IB.�Be������.�Gu�3Oӳ�a@��K�-SjۛB��
]�᛿L]Jzp��٥`{R>$nz�k{�[�l�nxN������z�V�[�g	|ߩF
��,c	Ui�\��ۯr��u�� եF8z����&z=��,C,�w�|<NRB�]�'�Zo��n�x���P�m��I���6VV�����Ҕ��h�Lh6	c�x@Y��X�6�z�GNO����MY��qx�a:Ϊ��Qy
ww���@��/�E��]<�W=r���\����LZP'0���}1�1����ʱ��n�\�G\�8�jU��镯�Ooj�[��-�e,�B6k&}^������%d��Z��(L�Q�ҳ�8Ɍ�s3,���g&�بu\�.�'�{�܆���B�����q�4C��r��f뙽@�Ƿ%"z��WU�R�ۧ�a�%ˀGXY�E�kg
�묬Gk.⠻��0�k��"]J+�+��oVF��F;$[�6���Y�ͣQKB��H)�\YYc���r�=��/T�8�:a.ҷ]yh�ٝfuZ<b�����N~|ݜ��J�-��Q`�s��/01%���%�pYm�)KP{��:�J���K��DEg;{��RvA�.���4�t�n������oKćP�Zj��{u�n��7Em4F�w�c��YnI�$�͠�K�=Y����[P�oـ�]�o�t�V&z���.ӳ�a�#� ֭��q>�݅0�}�+ 6��.��c�̨U�Jf9J��M��΀�J��b���4rFt���-ı�^�[�&b�Е�WVj��m�ۃ+������I$:�w34��BE�Y~�Q!6�?t��+�r��5���VԳ�.�]Tz��ʨl���Pk��d�/'of��}H
��+����zv�f���M�8�`b������bEEg������i��J���<ONi��2�����>$p������i�)�߰�~�C�s�g��ߑ�P���y�,�B��~�*f�������"��T�;h���I�Ntܵe㑴�:�&���0Zd(m��^��C��s�[	{��{ćv��og�Kfl4�/��Q��k��+_H/�Š�pP� �[»����$���x���N.~��r<op�zڊ�H	����ɩ`����?z�U�t�)���鄼��ooFn|�5U^�������j&/؎���U�h�: �Wݘ��=���#�V< Q��s��\�m�+6-��Vm�|64O������"�ց��,�>*iR��v�
��8LT�9:��+6}0�����O�����~>�@ $�mc��(  ��cm�&v�Mv�Izn�v�1��c�tu�l��*u؂����F�:YR�+���#B6f&�ܻǂi��Mv5�`a;A�h�k�B�bd�Y�Նkh�1��B���b�9�HѸ���T��Z=QҺ���i��[�R1,��!�4�x��3��f�����/�q1�s��},P�=��:'��C! �_rL�����E]~~b��fY�іfI�M��>�8��U�=�����3�Y����K���>�-L"b�6:���~ه�$��va H5D�n�7,i�w^r�#K�g���A���H&X�������0^nE�H�v�M,��<�&ߧޖ�������rMy�cOWu�����&�0���<'�͹F��-HT4W�R��!<,1�|����[ji	O�m�9��O�ܣG�g��l}�0f;�^�;>�h�O�eF�١�-{�r܁�����;|J��ł{HU�U@���ǽm+F7\d�#h��3�B�@�hA�}��D;��؄v�<����h�-�[�~ѡp�β��=�P^�π���NI5l��l"}�&���c��T/<�����<T��B�uT�p�J�nɛ��~"��ݬs�Z�*�V�+j����	?�}]DMP>�vz�z=�[J�Ju��P�l�~5>(Ṕ'��~!�m$�i`�)�+)���\�͜�I`$�	@�#��怣#G��x�R��޽�#�c
+�_g*�G�V���q	�`���h�7������cйne7�J�d�x���S�̋L;����R�qJ��½��y���6���T Mߛ�l"�jf�l�
b��Xa����������{ST���D�&S�̗�	��v���T��n\��݉Z�2�D��A]���
�z<�_K�>��� W�D������Sly�::i~�c&ԋ��z�lU�w�$͇'xš.NqD�{5:�2ȁ�r�u\!�K;޾N_'
��~������"D��Du�9W]����a��pDTYZ��U�%��փN�[ci����I�S+ u���[%ɢ�Xb��h\	�����M��'kb=F�m��o�U�:P#oӺy��/�@���E��9�b�_����;^�����sV��J��aWƗ3wW��V,�q���/k�g�L�/D4�&�>F)��1�>S��0������a���l����*e���	B���R(:���p���Y��"҆�5%�S B�ST!��Y~��;��"���Ra�����N7o��36�5�����X��nsg���u�HJ�෦,x���B�ُu��p�CN���c��I�~�����f:s�� v���վ�����LVh]]�yٖd�J����	+ʖj�ffK�6<ey$o��<.<��-�e�����j��{���(���zӗ�k��e�T`W��{��7� ���d;�ǝ�V;.�MSe�hǙF�en��"M�軳�bv�wP�>�桵ܢ���1�'|�F�nl�x�ג�~��Ī��������Jd4�vH>�#��sn��R00�4�+b�,V ���nR;|i�=��>[w(vQ���3�뗞�0SP�,�ɂ�9ք7&]^���(�?L��ٷ�n�܃3�#���w՚�r'Ob\��Vu,���wcr�������
��ӭ�68�h
/��{e
�Hqk��8ԕ�ٓ��3�]�h[��ƫV��H��a0�7c'y�gsV�t4�)Ep���ȸ�ǲ�]��:j�<X#�aw���`��\�������"�%��h"��=w�w���]כF�54V�CM{�x� ILϥ�^4f)�\b�|0�L�P��_����>~k�7��\�Y
n�:�̉���w.�N��k�ݗ�M�yt��.�٦�B$��[q�L.�t�ʮ�/Q�#3t�MV��X���ǈ7�n�p��gug��OOwemڮͮIl0Zj�)%8�*oΤW�^3'��E�����۝��Uu#�&9&�\ܲ���^�k�~΃��	��0��)b(Tq*�6w�C�Z-U��{z���#�N�Uq�^�E	�A��U܈�d��|��WJ�j�Sd��C�4Jӽ��tLh��Wu�G�tFa�T��ץ)[�����
�ʸv���陛�?m��;y�V�t�3��w�fڼ���ߟ>~}�}�Y�m��@�l�s m&���m�lm����ɤ���Kf��+��3��X�F&v�u�V��٭%�/Y���LA�����#5���FT�f[Rj��Yu��f�ThiF����h�+f!	Bd��9y�������tL7j��`��]u���Ͱ�e�ib�i��O����aR��*�Dʥ�n���~������6���0���;�h��wk���᥂s���oW�l����X���?V��WH�����Ʉ0H�~�Pw�ǛjM$݄I��zT
�	�љ䟇H�8Ij�y�]��H˼��+^պs�[u�!,���kJ�\�������ƻ�+qC�Ψ�`��a۸�H"+��l��޻�/�On���)��/�(�-VC���)�`tρm��'%X�٥���ʒ����'�d�,U���t����{܁e$���K��ur��Q!��,�Sӻ�eݰ<�vc�E9�t���l��4v���E3><;^^Z7���*�MD��O�$���s�f`u`4<[�@~�77J�UY��d]� >��b�k��i�a��k���K<m��޾�t}�P���&�����!���Ҵp�2!�|��t���v�ά�N�X�W9Th�O��SɄۭ��[���h�|���;w-�ⰲ�u�=�h���$��#<�V̯B<}U;Ѥ���i�]A�>~gj�b��$E�6�o'�6a�I��e�˗`�b@n��6���A0؇ �8�^{Ҥ�D\y4���&��WVt�o� ��Ǳ���|����!�rC�X�Lϓ��s8�I�����}��_�TᘚJ}�r��Ǐ��|�O_m�\�%<7�}o�+����J3���P�M,�c�<�G��X�c}�:;�)��ή�]M�4��ޒ�gu0|�,UBj \���:¨��uQ9��L(!�P�p+O�ڨ�K=9���4O=բ�ydC1~�o[���伬#J�4�jVs#�tv�|��'�_�$�7=.��s��a0����U|���mH�a��{��X�=Չ�vw�zZͺw[	� �?a�ǻ��`0�K�٘�W)C*Z�Ը��Crp���J-��mZ荒�l��ZuŶiu��9�aA`�a�E��ų���bLJ�R5�k�2���f��'f'��X���]l��O�3��?�,tK&��ئ����í�2��F�t;�/9���/4-�Y$7��Pm"L���Z*x����%�ƈ(2tW]�j�u���\}<��rU/0��&�����_�p@��mCd��ŏI��Wj��C+ݬ��6bW���Ms��4zx�n�ZX�%=�e�|p�f��~>�<iL��~�!&0S��=�(�$���2OB����cW����&��Y6Ո�ć��}���ҹ���b�������v�!��j$�Y���W졶k/�_�|��c�j.�����������4%:�e��1)zߝUx䛼x��M��t3�O� ���j_�z��7Ŀ$�m$�m(��d����nj�\���T�����$�^@�u)�2����S
��૓��e�����v:��졻����d���ƾU�F�k��W�1����.ޞV���߷�7y���!z6r�1��LP7T��W�͙�{�[�i�s�4j`כ��tpԴ��S�וKv���lf߫U1i����!����h�cfiI�]?�C�Kb���f�n�Y�:+M<m�������޵a�5��6#���t��$ݤX�0M9g�~fy�]kL���Ϳ
K��ӻ��>�'+�9S���_{F�l��4�{����Ϋ�q�`�P_؅0��l�1u;:�sU�0�.QꝩЬ��-v׭�[G;[�*bl��<ͬ��lLʏ_�}Z��>[	B��������*��1�t�����p�E����[���5��#q)tn@A��!�\�&Ƚ�,{�8�;��zN�	spuUI� a��vtL������ѽ	��6�q�k<w���T1>���Ҳ�)5�=~�޺��n�1�KAI̒sg��{D"i!��x��>�Қ���Qp\T�q��K~~�����Y�1� �#�+��?yFP/I.�E,�ó\Jv��*�6:�]�yz���s�v�HH [�T��^\!�� xg[�UW��yX�ڻ�6&��*a��!�d��y�K��o�j�J��<��\��'�tۦ�`� 
km�����n� l�` u�Ml~��S�dCcM�㶙q�q����7T�W]�ʨݣ��4�`�cG3[�fn�&�!e:���Z�t��F���m�ܓk�y��0�e�rv�^�����H�`�X��[n�iX:�� �N& p����Ҡ?��~V2��G�yz�0,��;g=�����$�M"�N�31Az1�"�OM	�Y�W��FlV�5�9����g��Nj�=#���&�Q���$	w-m��n�I6�N%Wi*���N*CǪ�p��ASu"g�(�m$�l@A�Rr�u�2�4	lG:����l��;s�7>Z"J�O@nd�
���ߗ��z��E�G)�*����c��n�N��&X4�.B9iC��3����TM�;�մ��y� �o{"f�s�h�/9�#���#ִyZ�M6������K��ck�\�P�2����Z�{��8���d4���FF�w����c�a]f*G���'b��m1���5�ǀ��	5Q�3��=x�8���G
��J�C�g(�$IQ6�m�.>k�ٕ�T�&P�	�z��A�R���:3G06���M����Bc;O���]����)ǐ���UnX����������k�2a��n68ӊ7�ٞ����pt:�u� �Cھo�ev:��%��{��w݈�e3ZݳPd�Z(b˛�d,ʅe0kW�S�ն`�|�t��#z�-�}Ϛ��G}��&�VZ��ʽ�����2h��fA��a��w9�2����"��!�n��n���+�x�x���Z�4L�}R�fvmguŗٙy��b9�M̨r�H��]0�Nbo�=z�iE��R��T�2*���R�H�WMlh@�j'7f�����!� dWX�X��;B��6��eR�θGc!s�#q�:y!Օ��"�-GdO/VO7���#HJ���~��U����i�c=�,���ϥ뾟u_<�µ��'j*�!F�P�fԘ��$��
-��.�O��6��5X��fcX���L�F�X e"���]�_ܧ��4潱|�eg��ފvW2�Z45�_f���r��*��q�1�ufm�{���6�dK ��,)1���6�f��W1xº�S���sm��m�[BK�         m�k��    
��e�hm���zU�&�[@      I���v       /YWf���       ���P   f�     u�[j��&Vi-�z���γ5�+l�H�`LJ�MaJ� �]�e���rl�jU��4ZM��R6�i-�R����P��Y���Cc�iX���*�Qaa�]�7���n���-�7&�v��sT5�:��*֌va��\Sj�K�Mk,)�)�m7
�]mݻfN�݈�q�t�u��y�K,Ĩ�Ef%�
�������;Gs�D���\��l�rʓhsX9F�m��׬Ҏv�X:�Z�::��y�Z�t��u�XE,�5��Ķ�D��c04���5]��.rG;Z�k���y�隳f��LA��`�kj��.��{vү�ڕdİWL�f,�H�ڰ�r8�7�χǈfx,�4l���T��� M��SI��\;a�Qqˋ8G[62��-��b��&ع�[5��-��[�jh�k��RR=��E�am*5�Rɫ�tnr�U&�k--#�s��4Y�,\�5����{f��k,�Gi�	(�Z,H���	���v�r눝tn�;v�hQR9�[�Х�d-JЖrm�0�v5��ޗ��u��2�m/I�6��-�J]u�[�J�M�&��T1s��;K�l�nՕ#*��f�0z�����/��:gitm���yWt��qt����M�3)()-�Mt,eBmq�D���-������?��fk�~Q��~�a����l�e����;���n'G`ڑ)_ܡ�XM)-�Kl8D�@�Jiu����] �������C��-��ܯg�,g�Q�uE��Nŉ��mv���h~��4a)��=�(���	]'7�<�9;$�_���qs\\����͂��,�i!����xu6+6<�|�.�)��]����8-�An�7���
=�DLp�aY(�3/ގ�
;=*��q�,��z6�U�!J��T�,*�}�U�z<�%�I�Q�I����6*Da��i�g�Nd �(S{2�I��=�[vd�/�=PrEz�&}c��M��`���)�Ӗ��j���-O��.��
��%w��W����`ݹG�4ً��f3E�$K�5�����Q������q#}AD;�M���]�gG���;�μM��m���	-��"��Y�)���l��L�0�L80,����z�uޱ����O�.rn �#����(��w���r����WoCy����;��y]RY����Z�tw��ܚ����PN1�$TY�f����7�E��=ӌ��oQ m'rn��.��Hǳ��Xw��[O����@LT�o,�zC�g���KL��}��}�3�F���Zi�,�@�^���_-�M���:C��
��6��u��2ǅ�T�ם�:._z�d�6o�H���2��WUy;���ttw�R�6��{`�l$��]%8B.�M�����:�L��*�ڑ6a�.'y��f�`+��_�P���2B.�Y�v�!���m�V�����?w�PY	���߹H�]1Ԩ���ʢ�V���2�{z��8	i�RP6��|��8�U.�V�6��]/�������}Lϑ�P:{�oQ�`�M�蔶�vò�e;�lI���K��^������¼T�޾O�n۞��Y�ݟ���俐�`��tr��^G*^/k��p��J�x`(ʑ� sV�Ɲn�V�O��;؍6�����-��Ӿ�l��=�ں/���I!e��X�$p��f�Tr����=��F���΃<���
�N�ٻCA�ۀ
=D���G��y����7�i�W�;ń�ɣ�,xzM�kj=K�*�oWi��@y����$1�
]�&qv/Ivdo��mw���	�)<������#��S��7���mβ,.�S�>�To��>�t�b�n�����.W������K�Z(����������%��#d����:�u~�g�7�3�扥���M� 2^�z��`�e����B`��'hf��~;�����Wޕ1th �MN�O��f(�WC��~v���S*�(I�>KϛN��d�_�g�r��44v׶�=~o��^���P���,���8�˾�BM�	&��+�I���g=�����t#
�<��Ut�u�8l�r `��;��'v»ΨN8�b����;�P�ڹ�C��Nߩ{��z��V$�ȸG�j��{�c���M{���b����˥S^X�I~��]�^���V��f�p�B��g2Px�m��m�hʷL`���m� �  /J�3���K)5l.K,��%���-�х������b��5k���출0ʫ�Z�v���a^SSEy�3h���hi�]��m�8�ٷ��ub ����L�%%�m�0�6�he�J��V�r��pB� �%�6?v�(�\�@�4e#��]���N�t�-��{{ Ӵ}�	3K��#�]!-,~�C��
������uLyy��ƝWu���@����g��_��l��A��#D-sq�v�ab|hg�,t2ɻ�W([��m��ڜ�����fD�E6�/�p��.�v�m��u���{&��τ;~�N�$@�u>�V�`�����6�j��"�(��x��Y�m���:������א������eS&�Ka.�h��,}���gBP����}n�F*�0�;��S}�L�nxx@�VU⼩{<��_1>��=Y7�䣥�ǐ'�S�Z��;��,�����+��f#�5||�R�s�0�b)0Y�5]J�~u�!��h������/�7֢���>z%.ޭ�0?�O\��
泮9��>N}>��)��d�l@M����=~G�����@q�{�d�$h�=b|���"���&R�����g޻�J�*���wSA�T�h�Ρ�'AWנYU���徻����t�k����Oi@x��1^�i�iqvO%��uoV�$�2�n��-@��)n�:�b����Mɳ�	p���0��A0Bd���������� k(�~�hò~��'��˻�����MU�W3>՚T.��T�{v�] �W0%{g�Y�5P^��h�x�d-�aGy�R��c�Ƶ�/ׂ�.�s�E�EW��̰�p�.����ƣ=�n������"/4A�/��y-1[�yG����x� ��C���}��q?����<O��O�z�v=q2SpA!�'ň[�l�nԎ�.p���^m��i���A�H>�eyӭL{ҽ�Ω1� x=���@�Dz,��p�p9L�y�/N�g�>�[s�,P��.q�!O�&������~9oU�w��Į;뾞����*�D;��j;��O���;�Uȯ7y«8��f��i&��a�!�K��im��k���o\ٴ�3I(@"	�d�1*h�����Ǻ��0G9M�s\�:5��<�J�<,8R'!JʔK�AM���6]�D�3p"�z�h��,�9�^�!caj�<��u�Ǔ��a=5ȵ�q�PXn�?Z�������bM)�ûݣ��C�������FL��l+��n잙���uY��7����M��s�z�|��ܸ��u��叡�
��ꪌ��;̗�DK���$ȀxRk�׽�c4?aݪO)�Z��r�4��7YhC�Yyz���;��g��'�m2��A��J<�8�E��xtz}��ӣ�$+;��O�A�����A��;@�Ub���6��[ X����<3���-�o�f,��j=��1�g��A��d��7�ކ`��)2��f��WflM������V?O��#�I�i6�0��l�lź�st�kt��h*�� �[�y]h���S�g�v���d@�2���P4��G�;a{GntOX���A��s,ʝq��X�.�d�!w�����_�	4�V�I�'i�j�~��^���_	��h��uK��ނ@A�Qf�<D�g�}W�B{�s�4.-x�����ʻ����Z�s��Տ+�v��]\�	&�n|�<�9�ݭ���#^��i��9Q�FbVA���I8�J9��{�p�9%�}}BnǗ@*"�j4O|��W�'�95 @��k,:�&.e�����	S{5�c��W�.��&-��b�8;<�^�uξ��[B���y�x�k��� l�W���?9�)́�;�Ù`	b:0{k�>Uu������P}��4��e9}p��&Y-"�g�M3������@&I>h���p�<Q��F*r�l�rk��#�F�^�2d$�?��l	�Re�
7ә�H��znJͮ�/�+!�&b礩3QǮ�nJ�tz���t�}���mz�#��	��nO��>���ucؔ����3�^q���x���leh"�P�ǌ�����m���r]����,���<.�\4���IF߻t0l*�G�`�/���t<����I�m��X�r�u'F{lA��dӎ.K:�㭖a�H߬�&�u�� ���[��S���#ޏ�ڙ�U��;��5�l�x�{+y ���NOs5�F�ԋ�kr%���^���������;]0 � ��L  �-�� kl�m�ʕ�Hv���%�ٰe%سSgu�v��"�7�����׍p�ڭ@�\]+���K���eD�^Ƌ-��̫1�,kaf�Nn����u�n��4v���b�F��,��itM՗^%��Zڱ)�tD��n�3����|\��v���@����I��vu_�Uq�%:c���j�Y������J+��C"���Y�1$�/�+���[�N�;�^V
�\�������˩��%�L/�pZ�)a��$���s#H��$Mzj�ѵlݶ�u�<����L��tl�цXp��� a�5����8�P���-����W�iW-�sM�]�_��7��f�xp�'QN�`6r?���� �vv��2�
�o��p
&�b�B��=����;5TW@1YV���q��&}�u��$XFl��Q4Kr�rh�z.�X�W���XT��Ȑ�����νV:Md�+�D�[���UD(߶��Yf������PpR#9"l"!k��m��Tj����nꭲy�Mj��������\>BM���_M�될z�9$�m8m�K7[�Ч���%�9��,���7��^�9p���g8��`z3S��Q_cy_��:2d��Z�ȯh�t��g&�0�(%0��6n��l�/j��Nu�7��v�~(�?~��q{�6�S ��v�T�$/�1X鷪4oX�����K�Ѷ�:E��ӫI�:;2�Llۭ�
�s��U����@��EQ1�564��XO�tצ��6�Bd:���n̟xtw_��wzp˂�4D�w��Y��S�����'/��7n߂B:����k�^v���i�yu\!EZ�3ĿO�}�É-Bm�e��"��g'2TT���Iu��P�̼�!w(�}�h��O�O\2{��5ꤺ���n������=�u[�=≀� ��{V
�w�r�_��rD������$}!�a���/s��e�����J���Ɩ{ӺkČ��dn��2�����lz��zX=�q=�Qd� ���T<��9��V��]N�
-M��o�Ut�n��+|�
�Du5�/���H�M�Ӊ�h�$�K2�
��ܩ�6/ـ��$�i���Zi�]���P�эSF.��M��.Fo��������R�2{Hf�d��tϮ��L.;ef뚘��q��h�d��{5��j���l�Ng[Q�,ιgJ#y�
;�ݩ������h�l@��{��*E�5�^��n�<)��}����2���$ΣM.�x}i�������*���(&�f�<dh�T���=w|�0��T���=������D������.����*,�H+��u��a�l�����`�Y�;��4r�S��y�S�SC�zH�+-����x��,���F�L��1�����f� 4j�꬛��D��s�1���׷j���{v�8�h�at��l�x���ʾq�b)����KҔg+s��߸�{]�D�o�@LO�����M@��7N��K�u䂔/�$Fe��8l�5�� �E�������1�K���SP
*{��롂�3�-�|�؜�䄖��>Y�� {�+v��j��U4��f�A����+<���˘7������|�r9���@�-:�t8��?�w���i��Z�T�J�T}��X����̍@�%�g��w� %I�P��Z}b](��*H+�RjSy�9sKRz�`92�S%���=	����CJ�}I䩈n0�t݊�o�-n�?�lmwxk��g��^m����a�c�XOu�YG��g\�^�k����\a!H�ɝR�m�쒺��H"|S]��c�x}�<�\᜸<�.-��v5�Ӊq|�2��L����9�{f,T�݋iJ(�U�^s	����c���s[�V�J�ǭ�7���
hŷ�l�Dff�{�(i�'G:�Bry�>�]豵yu�y ��TL9Z�o��ڕ���\/n�i�UK�9���Z��Ow�k+r���ݷtv�4x��@j��\����ـ�\ 9���Zt��w �E<�2��-��5�;Zau�n�]����Wt���w~ɸ����2���#�*����2�f`k�t�"�/����nd�������e.�k�|���/`1m�*^�S	<r]-��4����\��uQ��=v�*UB�+�����@�����U����X�y^n�S���'�wړ��ɮ���|��f�s|̈́�컋��<���b��Jf�Û�;~��#'��y�ő�\껺���'v�HBr	0G��'�Y0$��D�vo �,��qF�>�{2���m���xݵx��ެ�SP���ҙkd%!�ۄ�,`E�j�d��׫2��Gf��0�zz^�q���&-Q�!E���4�훸��립�6=�?'��[�m�M�T�%�I(��q�m]�5���ʹ9Y��O*�<}�M��l^
�E����q���?S�>�ug���z3���-6�)�PT�.4��O���ˍ���A���+��D���a�
V}�U����װ}�l�ͯz�PC��B�
9���Wo���m&�x��O�g�M�V߲�-�ŉ�l�"wU���邥yfG�S��Bϱ�� 199��C�Q��,� w�B�<��vy�M��A�'������s�yMwz��]�'n�^�0��yM;�&��n0Q��9�i�y�E5g:Mx+�<ʹ���ϯ��������  [x5��� m&���   I��'$����:nmnft��u��l0\����oP���4KfyM�E,���aaMD���Сn�Q�5v��(CK�.]�Pin��f3u#�C�%�͙�T6}��N�{7�u��{3BRn��!.���- �?ߡ6�����Fp�N��R&��L�~I�/���ިl�o�9�Q����x���,
X���h��,t����˟�^<�����P.K�:#ۧ�4�
9T��O�c���ɺ��@AÀ��@P<H��H�=�|weV7]�;���=?l�۶Vےlշ�޺V����ju�֦����dC�+�p�z�[O̱+s��e�
�D������͊���i+�Y� ��N=7�cNYN�9�Ʌ$_��g�S��W/2���=ӝ��E�X���u�Bp��@P��.e����E�@*���b��c˷����Ƹ�M\����v�[����L��9�)y�
{qv��_1vo��^~7� Whv��_}��&�E8���|��u�ֵ�S�]�|�%��Z֪���"�t�� ����h������3��VˠՎ�b�SIhw>-����b�oLh�Aajy�����k#u��6n�B����O�?=���c�y�cA�N���I��}f~Н�������9}��3��x��<+I��g�@C��:�6]X'5av:/�3�8�-��D�q��q���S����y�di��{�BA>�.T�$�e�@	0�ᥬ%.Ѷ�l�2k��J-6GE����.�С??�I	�ۭC�<$;�����
$μ��ܻ��YY�5]��8�0���H�aEU� w(@$�?I�j�l*�9�k�׬b����D�o_T��sRLw��U]�=e_G��s[���M���\JF[C���2�W�%V)��r�ZX�X�]�<U;a`�ct�.�*`O�;��O�#�}���7�50�<�f�\SDQ�"<��g�'fUeS,�"��������Xe�S7����� \����@U�Iz�N�x��- ����{�a�[�I��3�\
��x�/�y7H���ϧնP=W�ގJu�qU��s/�=^�3��8���	�?a�r�u1���γQw�	wƶųe�hBޢF��m�����פ�cN���um�*���X��b�B���g�<� ����y��='��U�I���i+w�Kj-ni�yS���:����o����Z-U%�^l���jz�a��P������<=�w�j)"�_Y�4=���,V���ɝ�Q��FA�,���^�D�G?uQ��w1 ��"�9.��,�Xo>��y=]��j,zJ�F9�;G�s����L����ӓB����z��*�h:��da!��>����H8l&�lȺ���''v����-H[�]2�~�[�@2���{���͏3(y>jDRP��+��<k�3����2��M#�+��j;=��\�8�N�H
��;�`崓
��e�w���cIOwҖ!2x͉����W�o���S`D�>�W@h�i���^^�����>n�kn���'=�r�'9�Ԇ�C/��	���9��e=џ�~n��ҋ7�Ѹ���RM� ��F7���z�Od��u����ｈe'���x0�Lt�����p��5�>�d�@ x�*0��	����s�1 �^8W��l*� H;&4���w�]�&�
#�hi�Xb��݈Q���?��S �e���^��h�"C ���M�zl�c߼32��-����O�Z8��kzg� f{�P�9�s�Hk�99=�榀�j�v9��y/2RbLNϸ��|���ʯu1&At��)ߨP'js�E1�)��~�����3}��)(:WO����
��l:�������i��f��ߴ�#gΕ[�=�Ό
k�8ڣ��whJ�U�<<MT˃I��'�K��f��$a$�1�O�ď��DЙ$txa�:	�g�l��a�m�ګu����X&�6j�Yn���.!?��� uu��]�u(�<|�m
��_)��\S5���PO��<o��y�.{��-MPrƖI�����=G
�J�=�H�e����~����f��ӘP���P�`�����N�p�C��p׬#!�nm��?�5����]/z��C<uڟ�z���g��ȴ
�C��9��W���{��`9����i6��~��&s�UIkJI�����:��BL�W�'M����@�u�8½�׷��� S)r�7�ps���Ď�i��� �j���Ma�-�����  =:'6u�[�]m��f�e*˹,��.�,��r���])���][����S#m���+�6h�Up;k�YNj󵆚�[of�.�X�T"Ii�����e%�`V�ը�L�F۬�-��8�s�V:�#cٚW��x_5^�S_��n+J��H?\~]魔<iW��eϧz�$�L�A9|nh�bR��7DmS�S���wkN݉ �N&����q�{��c6�*��H�s��z�]�~�&�y�O#��D�]TQϽܼɄ�z(ⲄF�x0�iOTjB�3w���8�	 �Ji4� 	e���hmoT�0�*��k�ib��7��n��5Fx�����8��wkޗ'(��v[�I@��m��[�3|Ę��A������`�PORQ��ݘlPJ�0�w�ٰٖ�yj4/y�_o�)�^I�>��`
p���5��9">�Ι�8�k�#��y0@-�V�< �3U�]O��m���`���G����?�A�&��(������a����T�v�(e=��o�4c�������Ⴚ���Jt�Z��j� XexT�7G��5�.Y����d	�7d�B�(���L����Y�cI՗׾�b�׎�?��'�_%��D���z%�o���ׇ�6�I�Y�)���7�8�b_����  ��o�df��T�EW:�G�˺��]���uwbyې�� �4-�Le��0���7�'UB�N����.�oM�,����Wl�A��ؑJ �y��f*n&}c���8m$椑�؂�c\�"<o6X��3���B($ZM ˈ뼳v�Ĝ�Yt�HOL����ʆHq��Κ����QľTU��:��䉂�Ԉ1���r���`U�%�!/`�j��y^�-ף���i�B�1b<�G̟�Jy2�)��ߣa�4���k�3�׿�>Ȯ�>�a�F�{n=�����໛�G�v�|��Ә>?j0�r&ms�d�#�z�����P�2�3 �>��X�3��_���}ձ��X�� G�ov�V��oȫ���uԱ��$~�<HX��US}43wY��DJ�T����v]�A8�~D������"��G�}]�b�FZ����>��Ǚ��k���������b$B|��dg��9��󃩺#�W΂�7��o�f$P�a(�)6��ާiE{�~�(n���I�D�u��pŏ��'�;�SR�;F�?!˔f}U$J8 ݅�c?BΏ��#���Gװ�Gh��˓W��3�6*���|>"8j3�DF�	���~��p�Bl��AO̟�[Lx|�eN�������c�?Wj<��z��P�l��mB B|�Nn�
�[L+labˣ���!S�����Ǝ�TZ0&�ǔ��b� �E��`Q�_4�a	�7���;��>�J��q��85��s^����[wY8��d�3*�pMWB�	�a"���{�-e����]q6*��Ʈ�
E��;M�р}��U���JM�hiRh�~�,A,���Ϻ��� �X��Б���1ZU�}yF����L��"�O���_���J7����G�ez�T�m#Ɣ���c;��b�F��>��iQ��G��2�!� ���H���+�����B ��� �y$}M�f܏�Dbjc�#f[�Dޯn_��G�Lp#�G��P���N"vz����	�"����D%��N�f��l��d�1�1#�ki8c�	1��s��&CB2��e���)�:@*'��������<!�l�,1�#��>���K� ��~�4Z:�6L���<c��z%C��a�Z�"�N�X�/�N� *�U���>��R&���s6�Z_�[=i)j̥�����~p���m�G����$A�^�`
�_C�3�z�b#��5o�o:r�}@�~�q�2�@��׮~�݃y [	$ʻ��":����>�D!�Թ1�~�"G"<�E�T�[�l�[D%
ٷI�����<�WK�z��uPC)��A0�5#��!�?{�M�`	"���	'��a1�=럪LdO���}�:������G���(�>a�y�/�*���j��w{�(��è�GC�0E��Q�;��r��F���Q���y�������c���x��G��v;yp7=��y"D!O��"4!��]�1@y*|D��4#����T\��y	��p\�P" ��;�_�h�/M������D ��/#bt��O��}+���I#%���i�sg7y�m�����Q+;�l˚����z���j�a������Fnv]������k��o���Fו�W�>O� B iB(p�f�b"g�?`PbG�5Qb<4G�M6��#� "/f�hCۡ#� �m��XBDx&c�F0���C� h��ī��BC�{&�"8�����~�lp�DzDb�n�bE������ۆ>¡F�>����$H�³� ���`�(��>���a�{�8�����S'p	�i�4����'D���#�.�1���M���B�!�M������c�`���
!
ĺ�Bk�U�~B��_޷�"�!ZY��! ��C��b]w{Ћ` p.��`�" ��̻pe����Ap�ܥ}|�:�ol����me�F���/��Y��^��6��-��������^�<�������#c�f�
���G�F�1B%r�ɈG���&:	�
�`�zL� ߅�1�r�Y[��t�-�&�U��}#IDǑ���u�(ANa�"OmX�a�0�{&e|������} �c�7�:�ϟ��"t�y1����p���C�&��j��G�>M��5DV{	��?:5,����'�"H�:yYH�[8�ک���F�G�a��Y��F!h��G�x����Q���x�S��9j �8|�F�g�>Z�I�-ѽ�z������M5�N%��[��o���^��h�w�x��E����4yP��٤~h��Gg��
�@k����E|�,Y� :+ܩ��0�Y���j�q]��fE�%���#�Ss�uqLn�����Yb��� m� � kX �
�0�E����0c�؄t�iSC!���%���Bg^�)+��]�qd� �Ԕ�h��əR`�͊��3u�4��l�4�l*n��3�`lJ�ĵ%)��-�`�Y�kuh)qk�u녲�#u��@K4����E,u���/���|_'J_o^q#�f/�Q!����`����j ��~��w����Q�T�C���M�O��W�L�dѣ��uO��_����A߱��وm��*�Ծ�U��H�!�
Q����m�`��d�p""�<�Di�8�&����X�#Ɨ�D1�d������ypm�a����#,�$�>�1,��yf�Tϸ����c�$}擬�x�>�M��I&�H5	���-�qK��s�K�q�~A�#
Fы��O�>���-̹��>�\��,d �)�u}!��0�G]�L�������=���(�s0cw��P�	6f,Q�a�J�T�o\m�Z�g�\��$B����������" �V{���;N��8Db>�wk�F�(�޺5H@ }LoK�s�S����Ĵ
l0n�/��C�*n�f�a�`!��
T%�!)��6��G� ����0O(�<MU�6�\�v>��ɳ�{"0E�}N��¸�	U�Ru��O	�2U.9���2G�.�f�G�z�������Ty/��{����l��&;��"�8!�r_H�(&�^���Ǩ�`��\���̗O���5�'a"]`��{���䳲�N8�K�>����g>h�B��:
؄u\�>��#���ޮ��(���n���Z�45Bk�ilo*�n���A��4n;wnn�l]#�N�(�ϦVW!3�U����MYʚ*�dۻ���β�^�u".�w`WS0=441������)�n�!�L+	!ѽ�����wl�����۫��r�H�2�P��"H2e�)�$8�cb����k����Q��s1ōKZ��\.`��H�4���Ф]h
m-�}Ku��ь�[�͑�:��C�6L���y�e����,�뫎;�`�o�HWwom�o~�l>�N���s��
��˞��I��:_w��on�wH�w���%N���z�aq�lS����s7�����n�ћ�MM�A�퐃o]6��{Q֜�N��v����V:���օ]�-�̯m��۔�U�N#��h�8�;0�Unt8�K�8Զs�;�7���Ulmeu��߱Lg��ޗ��+.��
�1Z䈆-�/2��Jį��`⛝sz.�'k�mA��Y��E�gM0�*��Sol|Sm�   �h-��\       �` �l�m&     �f͎d-�@3:]m�k�9"f      mn�      �m%�m��a��m�    �6� ��    m�     �7Y,u4��T��uv�:%�m�V�,0�p�����MuK�Z�<V�n+ZP�;+
X�KH[F�jU������;0���v�	4�f�B[�4Y���ńh��3W��m,'j�Mں-�{\7j��V]�Jkwm����F�c��Jʌc�i�֭5�O+���n����[%H�ڙ�	�ix���%6��:�R�`E�#vb�ʽ��M����S��V��o`��il,4�A&4d�mU���f��q^K�).uk2Pu)-��vr�*&,L���+�l5[D�g2˥f�k��P�kn�
�Tlu��k���ͣ�Y��h74�M���M���̻Q`MKlR��cq��"�9,1�Y�[�r��4��$�e+�,��4pb �s7h꒥�A˰��e1��o\�;P&X��WRis4ܘ�P9GZ��0ܻ�j�륆El�)��i���]���!S[�x��խݷ���lc29.׬�Z�r��Z.�����Y��Jˢ�����J�����զkx�ZK4齺��jC��5��p�JXܔ.:L(��P���іsW�,ԛ���.����`f3]�[�t�@M�Y�-S���Jr�u�T�7Mw=4�y3k�5��lݥ�Y�H7�m�E�M��i'vn�bd��Ԇ���
�}���l��~���D�C�Ş���r��<7�(0�X�54�I��/��5�T���)DQ?|�Ϻ=�q'���NA��m�~ ��WMVj;������2p��z�}B1��5$�,���w�d{�#	��T�|q.�ގJ"��۪�u���zi��@V`y�A��v�����0&�D�0�`�O�����ϥ�	�����v��!��ŏy�4�GU�I���f<�*�Bp@#2k�B�<�͂Q��p+r wY�:������ج9c?�����+�1�c�޵"@#�:�!�G$.����L����,��Yʙ���ȡ��wW�{�$`ň�y�������@E8T;U�� �1wt�$.�����J�-g�MUc Ցf�Q~S�M;��.	����'�~��&+�X)�R[�츠��Ѽ�(&V�
�^tv���x{)�C�u��|��F�"���-Ljk�7����#�L�t#!�p0������ǫn��2���꩎F!�����y�\'r+��$Ѫ���7��M���\ �i�|�e� ��H#��sK8�s�)/M�,�J��e�&>dC�(�2s7������H������ƕ`��y;��d�EEJK�k:Fw^zV�ț4Q���;r���-n]�.a}��4[w�W{�,}�^�T�ս�?�E�d���cH �VP�+�h<O�ix���HC��Er���;0j�8�vK�"�5�WڭCW�%D-*��Bk��J����,2��[����K�^[OLZT��kԇ��ؽo�ٹuD�����6Wz�=�h%wK�2�歇���T��%8\,��S��o���E5���W��"[�t������}>�Y�O9f5���Eۑ8��lС�\GwT�P`�+�3k��;�ٝ�(*8*��9
v��#�#��&x?p>M8�����jN�nV�d\ S4f�×��F�b�_0�2J>���z��M �7���j�)/obw ��O�(��y��PM*l��I�3��х[�ˋ
2�~���Z�ʊd�Ʉ��7�/��~?��`�Qo�=w�Y0�X|�l��3�g	�=˹��ݧw��vj&ȑi�7C���]9�JlG��$�u������F�9������b�4 �p�]~��N�Xvy��~�L5�L�� ��,ù��O�6�)&��ǔ�>1l�ǣ8���zm�1����Wm@����;����`��e*E�77�ncF�:ǃ#���H�~�k�U%����,�CY})/�{.bF���Q)šQ/\jI�Y4+��L�����!B=�A���dc�ao%)<�(�}Q$kǌ�M�^��I0M:h������z�&~Wj����Q�+�YUY���%xzH���ֽ��c\���o�,~~w���]%�f���� ᖙqլ�I&y��w��x�Y~3�(��Q�-��^q26�6�M��uXsI�n���h�Խci.�i�֪�?����}q��7�K){�bY�<�PG��� 4����۞J����Sx5���N`��f	�o���grrI�aD��x�~V�2��3��C'6�Y��;���nbC�׽��=�c6�c��c`f��$��p�A���L���<{����TáD �y���u�t�P����\ғ�ط<#2+j0�0�]��;��������jq>�S�	2�^U�фu]T��{9����j�==s�U.VA#/�Ӥrr��g�+&�Lc֟Һw4�w3��f��7��� �`&�3m��v��`  �>N���m�.�y'[�[&�1(M50��a����Ȓ�vt�۞�U�J:N�t��:��VkݣW^�)]a�"�ҍ�]��ѩY��\�#�lm�śB8BG�]���`+u!r�GK�Mu\�%6�U��/8���F�������G�J�9(h(/w��i�"сC����f������$��k;�xq���~�3TL
č�켃���j�iz|a�H�@�9n;W��̫�$0� ?]���	t���C���Q��Zs��^��U%�"�u��:K�mY���$ۤ���E����˃]�z�_Y|���Q�'R�C��;��p�A#�F$��S��R�H|�����nPΙ3{�̔�`"�N����|����TH�X�=��sC֖�t�E���7�;Խ{� #M���p���@�{��Rew�Mҿox��4�M�9 	5�w&�M5���}�~�7����J<\'m8N���jШWVTH�+�V��y{�D�a�E�'f��|JI���i��0|Tͱt�Mh'��;�Y�D*����ڑ�|>53�<�Q5}s�(�yL]R���x�zj_M���������o,:4�8V_1u�&�F#��GS��˺�d�I�'��6�O��b����Y�Aj��X�+?w^;ɉq�,�:\ݧ&�8QEm���]lV�tҌ�K2���.�OMz�g�p�z-���~4ݞp�s3��?#C%��f{�_���6����mt��N��U��7c��mgY��&�[�㬳w|pՁ��:p{.[ؠes���3-dF�j��C�+��~��jl7DJ)�zf�6L5�<�x{*�M�Zb7wT0���n�@� ����usج6p`�F��;�T]:dnX��rs�*���a���$X6Nd�w�t�>#4G*�V��ѻ��I:��?[�|:G�B���L��ܾ���R-'	���܆�fח:�����u=g�{��j�L�-AI:��p(�6��]�S0��x�9�ōOn��ىh�P��#*-��&���qU]r,�?+�-FנK��8& �[͡�Id��y�������><G!;�Oh��A �n��Y��L.���ZG��0������mmyt %�Y��u*[�q�&�,�I.���n�5hw�]M�� ����zm�p�F��ʺP�	����O(��`�������63��C�M���Y=�����թa��t^q5YRz�7�'ұ�!��2a��!��.i\ܻ�+I�og>�}�T�81����Dz�W�.]��
���*&<�ѽ�ӣ\z����m��'
I���hq�Џd���. 6��h�E�d�A�z��;.eF���R�=ދ�i�)�ޅu뼽)yG��#)��w���y��l�S��+	�2du��X���Q���xp�^ɠ�v�ߧ	{�L[�U�'L�L�j炦�n�w�8('��FJp4���2'&�ី]|���ޜ�
=�w�+�I*z��~�F�(c͸S^'����f���l4J`Z�s�k���-#��nD#��PI?���"(!��l�,i�'6v�Φ����י�>�߬wzzM"d�@�3��3��q������x(��4;w{�CU��f�N�>�tr���s��5�ʯ�Gw�B��2ե2�L���9��ܷ8��ia������p�ڟ]���v�������W�&WS.�瞓�B��G?N�S�w	���16��7� �vҺ��
��������2���T>:3�V.A�]T���R�Gf�{.&ܭ2�RGz�~T���}��i�p�.|��}n�ۙ��`Җ�X�W�fym��#]h"
�j�`ab���Ϫ��W	q�W�0�W��2�`���V��J}b H�Ǯ�]W�ov]���`�#�JyܤR�fI��wY^ �Gk�T��͑ĸ)�Բ��l��&���I����";a���{��6�I$ˀ��y��mg2�^�����CH� &X��`��gG#�9��S����ޔ�X���`3���O�s{T"�I�nR0�4o6*+����+��֏�]���;U�!_�0l�6B�U l�|��+��Ga�|�v/��`�e��q�iy���z&�)�`�O�7U�h�p=�։���t|$2{�i��fe{��حR�B�14oz7�CMBL�#�-+�ӹ[�1t$/p_��"����L���ʜ�_�˲,A�X�ـ�b.�ᡊ�l����;S�݅G����p��l�y����,�����n��n 8  m� $���:[e�kkU���JƷm��[�΀��kػJ:RɈA4����0�.��hJ�R�"YqMV���K�)Jj2���$b.��vP�چ�8aK�֚�i�ٕ�7��mnZi�X̦���-̀�m��?��|xO�'<U���,�XX��S/5����k[~��&���t5���6z#�h�r���dZ�Q��FW��z� �/���X�#��yU��t����E����vh��
e+!E��QW9`N�P���������W����k"��`���^tQu����ّ]Hh�\��j@4\n�����v��5�L �kBjt�>g|�I�Ut;�כ�^��^!	�G]w�G��]ޤƚ�4R�o����>�ѓzq�V��_���(��&�|�.H����j_^x�-�ʄ��\���q���~�U��[�?����k'�m
�hK��R#��!�]����(qIǼK�sn�_��&S`M7�����='[�Y�1Q��\�f�҇eM�.��<�D�6pl����H��{�g�L�f=|`s%��o|/�
���t�t��7	"h�y�.����z���S�-*����3÷lsի�࣒�2���{&}���Ũ�N����w>�ݼr((R�^2�L��D��Iεޖn���g�����>�b���c��@�nu�m)z�"��2���:�63Wm��m}��_�w��dٞ0}�kc6lw�U�.Hy���S4f�K�&��L(8*�`������T��E�fn=g&W���yn��b^0g����ۺ�72{
�L��y��e%����d$!���[A�A�%�-&��<V;+g�LJ?V���7�<<g��SW<G��B���sIM���(��j�]b|#�^F�̧cR�P��2H8	:nuQ*��QյԪG�Q��Y��3^��	�h&�q>썗W��Ή
�zg�&]���mH���%,M�U�3^��8�?����W�����r�;��Al��F��b�ŵ�FE�EW]�V��Q��-��m��d$�ċh3-�HƱ�������CH�	��?r����o���{�
��Od�ƶ���'0򳑪Վ��a�)kk�)��[Zș�+5w��rE�n�H����K�,A��D��m9��$C���fAj�ev̐�+��}r�qy���T���~�k�S^Y ��o<ث�AܮT��z��Ym��p7Wb촳a���61��L��m�b����yVɢ&E�!�A�Ԭ����T�wq�m@i��x��^m"E���Ȯ��� =:2�+�C祾������UWGwx_�2�,Mx��]��2���: �F��|�>LdiAK��|��pv����G~��χ��M8��������4����޼��r���F�l02�rE�I6�%��N2v"���/l#s�����_k:���g�&'x�5�+R%lZ�e���~K�8ox�P
�������0[i��6̣
ݽ��B���!ڥq��Ö���u�&uy�\.V��gnT�0��f����e}���z���o���ߜ�'����   ��;����{�wN�'~���<�I�|���:wwN���y;ĝ��	:I�;���:�������C�����gG���wO#FNzN�t�t�����w��<���g�w����;t�'2O�t���I��N�;����������ww�<�t�oRw�|JO���Iĝ�;���<���|����ۧ�y������ӻ�wI;�n�������N��;�'t��ӻ�t����	:{����N������;�ߝ?w}�|��'~��H|I�o���{��oRw��������;����N��	;��t�Iۣ�t�N��������w^������ӹ����w���2w�?���O��N�� ?����sw��?#���ĝ;��G��I�;�:t���'FN�N�t��i;��N�O2v�����y��;�o姉?���O���;�wN�'|O��x$��<�����������'|I�I�$��|Y:����;��S�?��������w���!�;�wI;�'�w�'���=������oh.�&������$��_��'O�?�wO2N�);��?/���O�I�3�;�wI;�}���~�pI���O���'{{I�$���D����$���;�wI;�Iߏt���$��g����g��D�~ӢNzs$�S�H���;��Y�?��>#�$��v>�q=��c�O�wO�=:N��'2N�I;�'i�œIݻ�w^��ᄜw����N��ĝ�ӺIާ�?�����O�:wt�w����};��}��������O���������sӺ�S�I�w�O�ӻ�Oϧ��Ν�gN��N���'���?w�I��N��N���'i�?������|��'~��w|I㻾��N��ĝ?2t{���N���~��|�x��ӿg�o�=�ӣ:wt�w�t�3������?�~���'}�N��a'~�Y������t�ӻۧ}a:C�wt�w���t����u�����O����;�wI;��v��w��l��Nޏ2s��<{t�w~3�OoR���"�(H\�wx 