BZh91AY&SY�{ �߀Px����������`�8�� p��ATP�Hi4�	�	<�lP�<�Q�C#LjOF��P       �& �4d40	�11�O�!�h      R	���20L�i�0��4LS##Se0#5'��=C� 2z���Q A Y�$ �   I�O5��~���`�"�I&����R _$ 4sG{i0���+���۩|HA�! PdbQ�PDAfBaXYaQA��Ӛ${B�T��y��e�O��ݟ���K�^����<���TK63��k�����.a�c��{��mFlƒf�n�<�Qs1C����7��d��c�G
� ��bA�:M)�k�!b�����D��߈t�����4$�m�3�(w������%���m�ȰɉE�z��>���ac��	Fk��F�!=ʓ*�;u�J��(������$�A  O8	�w5��mpY�$l��9F��Ix��fu|��S��t��"��6�=���e��M�*�`P����\�\,Ox��� �p�I�J�sa^5"�΋bj�o����56� (t��лP+{�3�D���v�)��v5fn�aoR_��aبi9X��/�����2�%�=ݚ2��R���m@,^&�g-
&��r2Ye�<��������fg &-Ca�.N��a�-k���Z�wV	|�d4nY9�V�-a4j�U�(F�4���P���#)�5��$������`�|��Tb)��w~�n�Ӊ=ae�E�R���7�L�Se��ȝB��|	e93��Ж�/�r�L����m�Z�c��mB���t�B7na�>f��۰���k���;BzO���eT��,\]����
�P�m�\ �����ߍ  � DJQ( ���R��h@���*�b�
v�,�g��ͮ@Pg�E��)^�I'0BD��V��ą�@�UYGu"��b��F-W�jg0� Ř�'��>��_m8'�c���S�)i��oC�$�(�� c�,R�s�A�8��3��y�ZL��&!����z! �RX9~���M1bKH��U��p�[�8�[Q�1d3!$�ӄ9xt�31�ñث��֙�ZܡG��y��^#�@i���~p�lj��g��tb���K���<T�	������>|����6�`���f}zqw�fo���ǩ�:��-��4�DG@�tI� �<�u����� U�MNE�u&^]�G�C����=%��0^�*���?:/���r&I%2�Hj�#u܊�M�A�'��=��\y�U��<��U�yp�`a|$*c����^�������<�yX��7�~�1$S�',`���^j�P�l�л}q0����,T�A��-EBt��4@�%:��������L��U(.��8}��7U#@�UUqUiMnQ,�v<� B�;��j4��b	�f��	%��YG!�T�b^w���3�|R��w9����8��B�GQ�}qb��hI'M���i��]]H5�I'-�Dunt��f/̨Jr0�"i�C�e@�7�� �7�}[�Y�~����l�"��o��3&���YE5X.&�9=�!$���=���6B�d`Yg�� ӯ*��2�^���A��+2��j"&���2z��>eB�Ⱥ��t�L�G��U�/����da)�4���ڃ�]��BC�T	�