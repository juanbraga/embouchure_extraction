BZh91AY&SY@ܥ�0_�`p���2� ����a��7H�R�U*��������cJ�AE��i�"֩TR�,4�1EҡRP�Սm5�������U����JH)$�*B��(�� J����J�P�(J*PP�JQ�
��*�!UTQIRUJ��(��RE"��HN� ��՛-��������n!�Q���J�]7Yt��k����[q�%�v�np�Svべ9seRۻ� .�R@�UGMb��ܫl�Ӗ�8Gu�h+��N�;�tPpv:h�6vd�p9�
ѮIΜ�+J��s]�Y���rJ�i�\p��̪����U�ds�,N�����e�)A-�.!�lt�Ӛ�
�sS�N�Ӄ�ҙP]u�� ���-ei���GA��U
'��u[.�S���\�M��f��lWf��sJѹ�WJ��LwN�wF�\�nۉP�[i@����]�m� )��R��U$\�٨��;�(Rۊ�):�n[��fswkV0WQ�S�ASw:mU�juRi\��K�u��b���� T�*@
�R��r���u�m�5��@.kv��S�:ӻ�6�g5��sU6��	P�s����ۺ4�.�q*Ui�v h ���
Q"�Uۖvj8���tu���)���mj�w;w����Y�P)�we�d��i�[.wwG9�ml���ٕM�p5R)��J�UH��B�ӻ�)E�t�;�u�l����re�&�imBۘj�J%fB�\����I�㶬-�t� P-E
���:��p;Wi�֢�(��g*ݲu�wur����&s��8;�V�0r[ĠP�; �%)J��]5��5��t�ld֜ܮ�;�$��5kPwWU�  5<�j��      "��Ĕ�T�0     �&�Mi��M)�y4���z�=OM��"��	JU            &���@�@#4�e�Q��Қ�ZgJP��u�MW_}*V�a�.�_l+Kj6��
�B�5��"
������ ��� �!�c�1*���#� w �^y�U�'�D����
E��(G�o����`�*�)!U�l�r72ʫ����y��2������M�yDY�H�B���.ƺ��H���h ]�I^V�+��w+]�u�k�ec+MY�M��L��w�7�;ٟiMj/�W!GFZE�WDP7(�N�	0E+t�=s^ap��W%� 8��^0�6��)ͽ	�J�Yt*���WF���I�
�Pʷ�7�,J�36SOr�E�%���S)�ڒZ�����&�䑳Un��0`u��;���{�lV���n�K�tpPq�Ti��	H3%-�y��9F�qArd�Z#�p�7a�pe�o1)B$�-�ƒ^��t�Ɩ��`WB�Z.�<)r��9�����y�bIX�̭�
��Q�����N�\��*Y���+Z�E�C���t����2�l50�6���%��M�$�V%]aCn!R��;�k�.�ed%�U�����2�F]���{6�&�9I:��wp8$��Y������c���o1�JbZ]4Cu��V���Ų�xc�k���F��M4�65�m� �ܩ�n�YN�8^ӽb&o2@��4��L�ܴ��AI�N��U����OUjǃlނAح^�f�����5��� ;D°T0� ���nLl�X$�*�B^�(:٩�`������-k���lґ
���ԥ�YP�U�wT챃Z%�`����lV�4��sX���[����e�[�xH��mH,�2	@'Ma��M���w�*�k�	b���̥ch6���ƴˤȳdͬM��a͕ f�:7.c�tƪm��CqJ�:Y{���uci� /���Wvf鲁�'��h���m<�5�Q`,wDCxv��n��� �u����t��#6�h�+f82�p˖�!ټ�F�X�s0ۢ�Q�l�'��!}pC��P�9BD�M�4c�lnI[Z4^�Gɍ�]KR�:�f�3UD��b��S&�#�X$!qꁌ���d��6(V�U��j��M-��y��v��6�v��aw�r
�0+�ES�BsF�	�Q��	�9���3_�h`�{5MX�*����M߫��(o�nܢ�\֋S����]���UG��.�����ܘ��W용�yQk�*�E��(\/EY��d�+��cXm3>�B�5�<�k��*��(��,��q
0�V����4�0YBc2���ܻQ;f���7W}��:v��B�;p�!5�=����NY1:0� ����Y�~��k�-R�kA񠉯TvNR���͚"h5�kEL����}LV�(v�UЇYD���ꁂl�DD�Q��"(��﷭��No����B�C���o"����%)m�������J��6+��J�
��::�sSA���#c��ٚз^�Ǜ��N��Rv��YDG�^�V<�]=��(��>�Da�4d���4� Ј�(��.ji���]��#J��*�!S )���l���`�(|�B��WM��6&�cKh��R�:��DDimÐupT��ͳ�*�F)nb���LT҅�]GX4;0�X�cuz��N7�:�4�6X�sqc�rL�v���I��#
I/��O).�nH�m��0"e�vT$]E�"^	T�~M�cA�@�n���s+�,6���|���*������Z�F��T���({��xՊ���?9#aV�@P^�a���h8�1ީQ�c��`�v�W )O�2��ST�̛��p��W�k%C-'�t৴��g40��M6H�����Ra
ݣF����U����-�ژ��r�dZ��oQ#
��K ���]�m2l�NϠڟ�O��è�^Iy�²�Dv�<T�o_�T��p��E�m��6��.Yx�;C@ϔ
���gו�$È)�ݍ��9Y/9�[p*�-��V�`������Z4�Q�o-�.9OI����낦m���3��\�h߽rl�YDZ�5h(�t-;��*o3f{��߇�-<���)\�T�-:a���ec%�]����[z `��)�W���@����
ڃI���x��ݚ4��۟2XAGhX�U��`5u���,CK��JD M53���h�4i9�P�n������/���x��c֡���*4�EѐڼU�B`LzrH(��.��60;���6��j+t���t� �2fKd� NCh�f�X��ԦqP���C�9R�+ÿ���n�����<�͞i����"-�l��=���T ��
�ƍ4�5�`f� Ȋ��Q���=Ԏ��V��ĕ��kf�}LP(PrQ�*��iRh��v3�g�*@P�P��*5�:��m�v�ۧv�]�v*���R*���1�f��D���+kb�ٳv0��j�-n�%m�[F�V*��������+5��X�JߵԦ�<sv��U�AR�sZ��m��uTvq�oh��)��*�U��ο��^f55u�-�@���צ>��f��1�ض�B;_%��{֩!��Ck6���wZi��������ܷJ�	ť�'!���up�esS��:�12���ܮJF�c)dW��J�ELK�X�nK$m���eM7���qd��+ft��+�KP��%�i<�ƉϜUǵ�WyB�b��Iti
D�)S�s$�;�̴���5�B��C�j��jF�5+R��9ڴ�L��)jƬ��f����:I�1e��3r�/d�B�f�欎��F��s>�r��m�4q(<Tbn��������]Y�E+�>ef bA6�eJZ��[�B�MSQ2�f&3E���aOu�>��D�8իe��S4���%�u.謕hi�9u�#�\v2ٽ4�I|�5�4��f8�Z4v�,Q�kz��d$B�b	T��X��]�3Z��;x�ۆ�,1�l�l��U�����v-c
�����!]�]]C��S��ʹ�^@��m	�IYj�2�CT���	?Kξj�z�߆(�AN�L˫�5���HZ�L�p��`�r��C_,5����v�0Ӄ3��[V
ѹ�@�A��D�Z�\J�a�M;�lQ+㶬�� d��BܩB�L��wW2��);�7�yu-��R1stkd��g��2���;��ni��OXx`T"j����n�o:en�[�`#v����Y��W~ݏ^<�¨�C�Yp̜�sAY�&;�Ӛ(��7ԥ�D�j+�
��͠I&��
޷��|CL+�`�Q2�7JnXQ4ʚ�N���kMw<s2�we��M@SIBZ�fP仔����ʃ~���5�4��3�*�f]�&�f�Xp�pLZI��WV]�Jl`N���v�w{����Ys^ɚ��Ȋ��84ɂ�E�7h��iQV��thhsL��(n!�aT� �"����R�6�	#W��{�-5*8]| �m�ti�ث����1;��;eް����i�5#n�he�+1bX��B�:Ķ���А*F�)�bc(�d�u�%������ �v 2h��MEhdāT��G��Px��i���k�͞�c����֭u���>��U��ƋF�2 �5G`o���KDaܽ9�)]�ɹR��6���d��ӣ.��%�.�ַ�D֛�)��/�������Y�k{�^w9�xLh�K�i�(|Ϊ��^�5Y�B�hA�Z>��(�4&|�v�SϢ�?�����V�̨Qd�(����V0��1@
��cf˻0E��U��G����kUS�c�e
�y�9�k�[��S���nԥw-�IS`n��f˔n�GXJ�:�A�$�P���M��TE��)Me'B�mZ������%�n|(e�@��uU��[U+S�,r�V;�j��h;4�P�b��QJ��Z" �Y"Jo(��n킟�w�[Rv�B��:6㡭y<�&`,�ͬ #���J��0��޹�:ƙGq�[5��	w>���m2��������B���#S%f�D��F��r�7�g1�-ُn�#��e�3^�.���Pb
�ֻ�P3lA�i�ǃ2U�P����]��+wJ�V֗�AX��K��/G� )������붩�VP�
�,Q�4fY�4Q܊�� �Jĩ����]i���+��J��9����D^���0V�6���ۈ/�C
�c�f/��,T�j�0j�i�`T�ul�"Z��V,��tcF:�*�*3�r�b��z"�_�*�Z{R3l�E���-m"��dϚ�w�k��uܷՙ��cMB�-��t5����Y����)P�(K��̵�j������w7��;aFu_kGR�-�����"1mc��يU�Л��@qm_q��e޵��Z�1�PM�V�8�k~y�����ȅ_ΎD�(n`r��eX��)ދ�WW���ȅPg��Z���e0l��9W�D�T��*�Ҫ�PP�� Պ^G�R�bo��V���Z����pV�K�U\�(�#aO�.�V��\���nH1	P�/U`��̽�C�V�mc�߃5���z.Hh
�%L�*�sG����{�u����<kz�3$��R�m�����n��;���p�4R��d�h�=2�Z�Uyt(P$fʣr�9��v���w*�N"�$�u��j�pH��o����1��}fiNJ��S�I�v��vf�i�'�Rt����s�|*���b�<�P�*�O���4jJWO�(:<l��&Q:�3�Q��EX���^�����(���. �˽���h���-�x��d*pO�	y&�6����ә2�rܠ.�n����2�Q���f���:ӥ�8�wxe�.�A�.GN鋩WZimPfU�p��`�ŗ�-��~;���L���Ed�L}`&�?��D|��b�5T1Ҭ&��o/*��蛪����kAJU�6RIDu�U*nХ��9q:�f+{�۫��])���nЗ1�3ﮯZ[>��.��Z&!�2�9Z���I	�x;s[���G�5�=�X2�^� j� 2A�a6���iJ�J^Q[)�e�����U�4���"e\���JR��o ��542�f�����݆ж�Q��'�����ʅU�ڢװ��B�Ǩ��jᗕ����#S5,��a^h�(���m��WPԠu{��Z5��S�j��67�t��Yt�+�Ӳm-��o����E�T�_=r�>�)8,�0����qL�h�a��;��^J4oc��-""ҭ��n�]��Cj�h��t���6h="Ք�� P�C���n�k(16���ň�e�eA/.; ݒ)���&��杸�h�z���R�GC�4.�v�J�u1���Z���khˢYX��Q�`�ړ���R[T���kkl1�C�D�N�7+
njl�XCtX�F�4��#�����1C�^���þ����L[7V[���r �i9#�1M�&G
X^˗z^��ۂSl��Z^�KtIJ�l�u�Z0�d����=kz���h��
h\t�q*;���wdM4��.��7$W0i�ܶ�@P���i�@�ںuv(l�i�h�>�sE�̘V�ŁQ��KE0�a��L�c>��l�-�l`�6ΗlM0��,˔�tɢ%�\�d��"�
�*3��[�~ڱf�<��=�����#n�����8�e�eZ��t��O��_]
m�F �sw?�;V�1P:�0/33+]�o5�G��[�rPi:�.�yx�LX��E�Ay�e�k2/��e��GV��h�l	�l��^@��s�$���j{K��n�Tb}x��Yb�\2���n�Յn,�7���7&mRl��9'�IAc%))ҺD�ّ���MJ�5%:2Ֆ<�����Ξ�鸩�E_q�T��A�H]�C1�`�MՕb�â�����M�"h�{��u�{��E���]J��tMdY5$�l3r6+(��I>ze3�@����gv�*�%Ub�!��aZ (_I�^�"V6]�����ܶ�ԨW�XO�C��@�	���f�\L�YA�EK	��Ŗ7q`��ʐe���јSѻ�	%Z䠐T�%l���A�I�3I�J��n|Y�k@�z,�ԕ!���P7Y�hVY�d�ֶ�c�SK����k����.�.���5q ��4ke�-Uwyal<�KL�k����/�PZ�{c.��Cp`�
��<��72���͔n8��t��H:�t���凭��B�o3E�/41��@�;&��H)	�բ�"7������z,�s,�V�eJtfA�hF��I������";�EJ�Mb��g̡`�I��;kw��Bj�;k:[e�%��X�(����Vt]干���I)j�������ɣA�t�%�����,k��%#���HIi��4��+j�c�y�v��7��n	����;Ma�*ݶ�k�G�
�ܘ�#�R�K,Vn+�!פ�qQ��5��ʁ���Hޘ�;{t>��c��۲�G�LK�v�.�N�-N�N����	�/kq`��֕��b��x�/(�U��6,�J��VEoY�Z�o9�iryk�P�V��"J�r��ӡ�.�So*$u� f�?�Sn��֞�ֆk�n)mU+��j8q���3EL����Q�(Yn���fW���Z1L�7L;q�����x�L�3Z�pc�Gkq��Ò�9z�r���3M��L������G�E�Z��_�+���������@eN�]����\۫���;j�5��_Low;S#m���>T���-⾌�봥�i	�+J�	����0r�[��\�n6�Y(�ήj@ky����p���t�z-IξBԃ���dw0�Vǘ'+�N�=�����(um�:���rY��«�ֽ=;Pa�U}�q�{�$d9n��1x�L�)E�!����u���X"�j9�ҳkXnga:�V�0�LTu;V��ê=���D���ގ���,*#)�=li��ίU^;�n����8�Җ���׆�(m�ʖ:#J,�]�o</&�{���uG�4�bo紃�W;,tݩ�V�e��_\��wW7g'��4d�wF��4��/�uj� +%�S4�v����:k�k[N�"uk��E՚�Mh�/>��)9�`���	i��\��աV�~�f���E����V�n�N)Fva7S�"3����j{	�<┴a�c��ئ�f��iQc)�DV�8�s�
�U��Ǜ��ʥ��)W@��U��NGDSr;a�nѸ��x8�� z�Y�N�1���҂	s����z�-�zxfNʏ$���Qƭ5.�%q�����r�닖�LV
�ck�8mU�\�q�D���9��}g���L��xvc8N��c��)��Ei�BiZ�ew^�E�7���P��DN�U�Cd����)��u�bTE���*�����;��J<�U���9��b��:�����M�ݾҎ��k"�|D�cn�5����!�ܮ�]��j�<6ܥgYI5�mI�Qo{Q��T�)|��R���\HWJC��WN��\Ψ��u�z���5d���'��5��+�G�%��+GV5`�����H5��SսL^&���-��V ����Ī<C�XU�`y���zn:t�<�ۦ�4�w�S|�.�%PA��wnsI!��h,��3�jLr�IP`�R�ŭcod	� ���Ϥ���*��݉.m��M�=ܔpٹ�K�1��t��Z:�T[�w\6��Fk�Z�U��WF�s�_�)}�9�	�hU�eZ��K��:o9�V�(eܛ���=��{��9nN��5m�;z����s'^���|ܐ�1����&�'���Z@���ˊ&̻�O�w<s��z�Ry�D��j!�/�N�Zk�Rҹ־��W=͜��Ux�J�Ի����gTZ�o��9QIRH�MS�>��z�ww9W�������}|���	�Q��r杆��H�ף��2�5F��i��np��u�r�ޭ�a9��V����L���ǩʝ��J�o[�RJm�u|��|y�S���)�&�ѧi�v��纏d�\�V�<oN�����H����=�=+vaǋme�w��U�IS�J:�5fbY�'N�8YI9v�q:o:��A��	����m���i-�۱M��$�w\�3} ɋw^R����Ϸ�K���$�Kd[���wRޭm��-ƹo%��ؔ�L5�^{�]�^�/֢:cə ��7n���i<�f6�]u��zgE�Im��[��f�g$�X�ѓzˋ'�26�$�w-�IF��%ϒ[�.�;wl]�]�4K&�RK$3��mo9�.��9�����V�>���V2���M��X��Y���Ұ]�1�e��K���R9}�*Nq����^�[WѠR�S�SF���y�a��5��@;3+��"ow�T=��iY�1N�y��ݶ�<Nط��E�D�j��6o<��1	��v�H( ��VU�ᙉt�F�{9n�C�RHH�=��ҵ:��	,.',�!3�eFQ�V�N��;j�Ore"��h
�--X��z�r�Y�J�A�v��$�e]��R��՛!�e�ۄ��i��(riv9�0����74�\(��uk�c���98�8���}����s�B:��1��B��Jc	S�t�O�Uؾm�r@�]��3'k����l�n����5��,�ΩҢ�0,{#����u�=.���r��6uXwm�%�1s��ɺ�!mڔ�g]ugP�}�,wp��Y��:�g\�����|�tT�s����g���],� ]�S7Rك���w;nN�{-%:�:#U��|B}�Z	��gRi-�]ܨh�CqP�$�.�o���ww.�I$����֒��$wweV=m6 D�=s��E��u� ذ���.�t�s�b�����9
�n���3q�S�@=��6<������ٹ��+��X����v:^mc̑R,�E%��`����Ac���O={o<ԉ���`kdP�Pf�>4��I�56Ey�gy;¹���&������S��%r����
3���z+Z�ōp5c+X���hpko�����p�
q�)��^���S��Y�U��ex��X�����E���;5+�̘�̜���h��tt�C���p}/t5��"v�i�˴<�77��ʷ�b������2�96e�i<�G_&K����Z��jn��xS�ۘN;��+u����!�T�j5GG\;�5���"�Ӛ!z�{o�c =�O���^v!(�9ec]Z]��ՋQ�s�HB�S�v3na���M�9�Ґ�����*3�{�)�R�Z{�>4�p���DS{��{g�mU����ε�h����ݨ���-'3��oq5&��N���9�vYK9�����X�aRE$��&�ڮ��R��f)PWp�X	0�-�KSwe�M�����,��K9ѡX�M��:P3�K�u���}t��5؈pu �u�N-=ؤ���MӘ
+:�l�Jfk�V)F��e�2��
k�3u}����([γ� ph�h.���H"��k�ӈ>�Ϋմ��Ws���n�az�PG\�\a�d�U�G�sP�ל�
V�%+����ge�_��`}�:LU�۴�t�WU�q��fZ;*l3z�Y	�w/�]�����dK��z,��D�2\˭J�i<��T�5�s��l>!���#���}�ٍZ��$�KX0�Pz����48�q�G9r� F^jx9�N�p�F�����S��0`L����@��Ky��&�
�Y�vg-�i=��M\�����ՄY����_4%v��2�a�t�'�5���nAbd���d�
`բU�A���LF"��h ��j�sH��0��5��J�9t���^��WXb"�r�<X]$��^f-�w�V;gQz:�� B��2v8�ۺ=�MǺ�����K4�$8��p�f��'5��-b����ݶu.什T@k���sr��7I��kl��Ԯ�W|:n��÷8)��ز�Jvph�x����3r��)w�kbbw5���لtD밪�r.EP�K�м�qR��/�W��=�2�L�K�V�e1V��gL|^+{�e^#9Z/EId��Tdnζ>�W���z'[M�A�a�Z�����}ӏ��L}�7��.�Һ�R�}-K�NI�u�U��=�p��or���)u��P	t{��l�ΉQ���s��V�����պe����V�M�ڶ��T��Ƣ˗j���;�;��+	
��j}������n4
�Ι�n��9�,����i���N]k��Z�q�82�;�����ּ��;o(��z�SN���n3�p�rp��yWjS�R��nj��`=ۻ4��swk	;�E�ܛ�W܍�[�D�6��
��É���clJ�7-HJLf^bZ�SWf���l�:u׬����;��e�Un�M��q�&�%1��`��%e�j��7Z}S1%�-���kkP\��vv:\�w':�J�����`N����I��j��;+��J��R�849��՚�ܳ!��o����c�����S9y	d-����:[�K�'c�#��;e2���5~��?S�Q@r&��\~��7gk�9��>IGC6���o-�/lq=V'0��.�z5c#�"p�(��+t�V���}����.�@nv���s���c�0�:uun6���k+f�hV�N\t�.�	��z�J��,	��Ւ�X�r�m;��1@Њ^��w8��w�3�J�k"��U���)2�����w�[���I�#(��v�+s'!݋l�����h��\�3+�����9F�2�em��@�T�������m̜���S*^r6w��k��PA]f�H0�8e�I����2���:��X{�#�gf��bѵNY��R�x�
�W679,�j�U��ưѲS��ͽT�d�=W5|���fTl�*�I�*�=>T��ԸK=������n<�ѝӹ��|iժ�#�Y}&Kv7{V���L�W��.��%f�r�*T��nc��}���A$D�X�{����fq����<�h���� Ʈ���,	�\�:�@(��ky�Jy�u���B=D�7\�5�1\�vv\7v-vf�U���i4��
{xC�2tv�2n�vfk��ъ}��N�r�t,�d[��R��p� Kh�����n2��bT���gROO�M��*7"N���g>{U
/b��3'e�V����Ѭp]s�쮩��=6+*![Ehh����ʻϓx$Zk��;\�vn��M>a�yyb�o7��	�h�\�h�+ �ku�4�lZY��q��X[�Z3h7yzD�h5s��5���hK�/{AD��Ï�4�K�J�3#]�S�Ͼ��K�'o�
��T�N.,��.�w;���.q�|
k�ܛ��|r�9��Q�ղ��k��B�*X��� A�/�kӶ�i����Q㹑�lS��h�ۋ��}Xk�}�]����"O@�߲��%��=��L�Á�m^T�}�Svq
�ً]��lt��&��ǵ|h=��r���Z���;$U�8�<� ڷP����TM�m��t͘Y�nہ\�b�Y��V%�y���3n$:Y����}��Q��:��ːsN#��f�tAf��kn�*9�v�^9�)��[ҏNRQw"0�T��ƞ���������P�#�&����\�b�$]�'E݊魙���Cq�6N[�K�0榪��[R��7p���Qa���5��R1�:p!�]�P�l-�z�RY�KH����ʥ����}�t�[���Y-�+���V��ͫ�ξ�IvK��a��gq�ű��h�Ȃyt-�|u����ܛN��g�Ы�\,h �ME�N
2ێU�o#]]-
���2�/37<��F��Kz�v�8��p��s�ҟ��*3�d��|���YC�$�5���Z��7��1!of��)�ѭ���Ɠqh9ph6�I��G�f�F���|�^� ��ćѕ�Eu5U�:$�׮bj��J�nP��j��j����>��[��Q�N;��1�Z��V�o��N�2���j-x�J� ��o���&v�ANʸk	�<j�v6�kv�]��Qۑ� ���Ҝo�-�c����܀i�w�j:H�Z�v54:�gۻ��bm2��ݹcyYm
�rK�U�� nն�[9'L۽�L]��zCv8}ݗm�g� �vH������A&+V�(-4֌�E��bW�h]�&9����c,VK$
`����12wp�r�v�E��=W�:��
;	�s㺰�g�y��������0����kμ�/A{\v���G#n�"��oVus&�9��;Ө4��a��k�����m�;�o
����IJ���aBc�e���]q�n�t5w���;7������$}N��Wb ��j%Q՚��S�k�S����;ę��G�gfo��Nש��R�2�R�(��9bߕ��blL�D
���b����,��4lQyy}hY��:F;�{A�sT�w�S�q��pX-�ү����u�]�T�W\��02!%�u�4$bCb��k#ћ#�|x4�qѣ��V1y��P7�Ȫ3���uv_��kp�z%\ǦP�2�j���."�oK��O��J��6ޫ�H���f��G3��6&eY;�TdnS�-&h�w���e�֧������\n`*Y͔�!�l��ݢȲ��!��%V~@�&]�-�:�������Ou��Q�E�ѝ
�q+��k�aW�9_Cɂ����S��х��������"`(6^�G{�(�Gd�4O[V���90��Kae�Y;-f��]����P����s�`}�{�sg02�[�E�(�k��6湗zz��^!��R�9"K���8��]�u���x�]��%�RbM]�3�T{ܳ������ҍ�z��Xa������[��W]��jL^�߇�8܀{ۥJ8�7=j�qf�����E+��u�ΐǰ�\��!����6=�o�=��ʛ����WL�Ov��0P��|��
�k�|Lk.��
V*�*����o}x�XR�jI��r�����q�������0�'�2:�YwѤ�DŐ@���s8�D(�]�w2%nJZ[W��\#$pe,�����o��kp[��n�@�g �c�U�9�Z��)������AA}*{�4�%�PW�k{N�7Hn�tQJܴ+���ͷ�j�d݋M�����Fo�=SS۵nR���]�k�x��c%觹}Y���>�ٻ�/�\]pR�UI�f��/��L�u�SV��nt��[���T�_h*=��0_�4^�>�d��|6��G��k���YL(�mC'fRݫ��v�u�j�X��3���,]4�\��FĹWlg˺����� B�+>�Lp?��i״�Q�(*�ŕ��N�}X�=����Vz4rp�
����z���nHzt�B��r� ���������3��R�gq�5������2	.�"�'�u�k���8�����a4OQ�U�d�Ak�^�L�S+5�9w]�o;�yv��ܵ�p�k 8�y\8Le5���@�Pc8t`B�0V�7F��u|�06�:찫Sl��sH�1���Eq�8\�E^�ؐ�FuƤ��Od2�nZl4kJ1XY��pz�GR�b���*}�.:w�닉[�iz��o��jMqu�v���7�uhMy�c�V.�r��;*sf�`{�n�������N��p.��y+gK�Ƈp�Lt��v�9�r��AWmwPTDu_ x��Z  ��xxsEv3���ޠ�I5�ݟ]i�`�a�O�.���Y�oK���T��h��n��w�u�n`D3�!6�}2�A��t�dǲ�`Xm��PCԖܔ w���^���wɌ���o+��'#���ۥ��ڷ�K�K:�=<fMt�`�7����;��Ԕ-�V�Ps~�c��m�s{&Ԗ�sWK��M*qq���f�[׌��of
��]��
]�6�A�9,ɓ���:�8����-c*�VV��{��ԁ:�f!��Z���_pPy�#��_�K._�_�Q=�JhE�b����nz�X�ʿڮ�罝t�geB\2��'ռjJ��6��0A�*�V*t�J�[��8��Ƥٺ��}�K�_�W�2�M�Ql_J�� Y���f̒���`���`�2�Ȋp��?qU��]S+Q�Dnf�S%���\z��&�o�a'����;�u�o�s0��8��j���,���\h��K�*^����Ч��QΎ�b�h�M�64F.�V��6Wr熎�u�ɬ����t0�ˡpCp�A����0ÃGkg[���W;=8t%����8������[�K��LS,�[ǻw��B��F^:%c0mbX $H�p^�RR���ʅ�qf�<�j�I�I�}6ʺXU�'i�ȅި�Y�2`��5"̘Z�\m�Ýv[��՜^�ִ�*J͇Z�l��6y
X6=���t�/��r�R�;w�2b}&��n��Y��o�y޼<T�BI6R�����>Π|��s�=�vFS��u�v�is�`��2>�pY��S��a8�v��Z,�N��;t�΋3��Ȝ�ǏNuCUy�F�Iծ�(c�e���
fF�Vˆ�l��P��{4��Ǣ����S��U��_��W��{}X7��u�u��3�.ug���B�R��d�����y���+�*����3�=�U9Y��_��{�z��G�ٔ���@a�[����|�@�B�wp��5��	��\ux�E�f�]3�q���}�}�ڌlkT>��ԁ4ŀ`���'�F\�3�
"�:9ъ,�"2�M�V���� �ul���=��o����{6ר2T���o��qMY�[-�8}�[��p����Ж�0wM*���Y]�P�z�*,{Ï������:���z���x}{�*� ��]���j��qj�;՛xY����PQluňufFoK';�ܴ���٨���Dj}8��u�m�޳A9����"����&��T^�=YЦ���}U�'u�T$W[��2]Y7�z�s7c��s����!��R �������[����\�"��c�.5#���<�C{��ݲ#�=��b2&�F�}�d��gm�زGt�� �s���d�E �򽨚'�+��w^���"�mg;h'jN�4�tuvFV�t�޸�O��@R
B)�r��y��7w���B�J�P�_e-P��)�\�|G�Z̠��)�}Џ��(�3����rM��W��<=�"����/�;���Y�qX3��72�Z�ŋp��]G���SZ��Dͱ���3T:;������UQ�A �APEUAEQ0Qb�D�1
EV"��d� �
E��B1b�AI���b d��=� u8���;]:/��p��[k�p�޴���n��u�U��]Uӻ�*	nr��/�$�+�k[y�)�`�|���G�㷛���|���a�"��vWKr��8��f��Mot�&$����ޘ�u��|hr�� N�ΓNO��T��͈SyƆ�r�GZ�Ṛ�g�⺐'��Wmm�S�&��X�/� ��w[☌��>��0��
�bM��r�}�׹�����l�N�K4��1xĞ��#��cwVÙnvh893����VY��U���o��,�J� Iy0bw�\��TQ�2ɜ��m�f��0���]E鍞��b�Y%�J�3�6r	�Cz�m���筅�WvѨ�]��^
��U�/p���� H��eL�s�4_��d�Z
���׳73�V��O��]�rٞ�͚������~����b�UJ�Q�(�!T�)J����d�[ Z�����ԩJV1o���9�o�����̕�*�9:��p(��&�Us�+��[�
[]��w}�w����W�m7p�O�xu��RQ_	B��y�Q1��֕����s��} �)�����Z���{3�Ǉ���Z^��o6F]�m�P�\�܁,t~��~�u�
r���:�<$xBjQ��e�;]mFA#�g������L@���g�{�S��VE�����=ѻRl[��+��a�!�]W���%��GM����r3�m����y�y���fyC�����j/G���QS�İ���&�BD��C�f�en��GL����~N��?" �(�"���HH�,Q�� H�A��" �1  *H�F0Q�Ab�{�^�g�g�w�f�k�����q�ۊ�v��a�}(-Mcͨ�T�Q�yEl}ܫVNÌYN��}�����d��خ�
��6�k�HG�����b���L��k�䐶�7����يg�V��ʕ�4��.�C�4_={l1}�׵��FnT '8=���þ��v��z����;��m�ti�9�g���D��skqn���À H�M�l��i���ӽj];O"�k7��W�����u��W��V���u��u��;	���&��  ��͂aHK�n%�pBy�c�wp�̔�Q�;(���]:Om��.�0��IB�f� <=�]� =�І�bz��ޮV��MH������?L����A���t;�*R��t��t�j�00 ��T��ty<N�]��T�خ����A��D2��X�&iu��Ӛ:�=������g�,~�ÅB4�'���n�B5�����7�~���Ur�̍'�������Kw�S#w��{�O�>b���s�իzb�:l���'S� aKn��I�wJP�Nk� ��X���7�h:��;�����9B�9]����',WY�*u�W���p�����q'y�oI�&ޓ��{E�\��Ɨl�/X�=ܜ�y�U&D���ﾪǕ�l>�k�m.U�2NTn��AT��	c�� A��8�=��ެ��ڵef'S�`z���R̽��h�U�;��x�39�:w[ַ�c��6��Ã=���[�.pA������"6嘐UYwu��_���/ƚ�{���sۼ�a��|%���B,Dab@D�#A PY`��H�� X�DDU`�� ����g�����^�����܇R]���=�%,�,Gǐu�M�t<��C�kU�+�k�}�iZ�f��x���V�ccq�99=Q�3"L�<7լ�t��J^*<�O�ɳ�C��\>�}�񄐇5����饂�(m�(*�*I,"��1`�@DX#Ҡ�
��V
� "�����(ł�VV+Ub�V!UR�L�(�#�mF���<��v���3i,e�u�]0r�+�V>�k��Ο��L=�A�<�ۙ���j�`��0R���lp[��94�͉��
��<�üͤ���.e�X��]�o{����X	a��C�q�h`/'�p��j�E���xx[���M-��{Td�������9��|�>w���=��tU���+�TM�zA�GF?x{ެ�y�-���y=����Է�5�U��|�5)׾���A+��]W�{e�W��gv����7�!��>�ďUe��uz����rp�r-5	�s��=#X
��x�f�����}��<�5�f�T�:�v��m`����1� x=���Kv�z��s81�r�����$��Y�}aR�}[��Jr��؆D+��<=��	��m�G�\�PuV��b� ���ДD�U�VV��B�B, �E�HČ����X(+$�-uH3e*�u�+�Vɍ���ִ�>~G^�R�,����J�/S��u�̾��wӖ}V$1k����V�u�D�D�Qa����j�շem��!,K�v���SS����=�tG*˹�Ȭ wx�fGU��n9,�W� Ԇ�贲��B}��.ʕ���fH�v�{�Ws��|���9f��U�gT��^�&�g��Y~��҆�1I2��z���Tw.�>79C�F,XEȢ�1��
,"ċ T #UX�G���}�����t���y��U,��s5k�؀��}�Y�t�=���)&��B}zk���"4�/� >���g����-ݬ�scy��b�k+����ڽ�uV�w�:b�go0���c*�3+JL{���)[��ѳUN���X�Ҹv00aɤV�_��s�߿}�=�����V$�őB*� �Y "�H7��W��ݓ�r/���c���ǊqjF��������5X��̷��5ͨ�;�FCB�MM�AG��+�GU�:X�}gu���7�K:H�CSq5��H�����zF�:�����S$NV�wN���6�f�t�O��'����#�o@.&{�z'��V�p�:�� z{c������&�����ªU�QJ��хw�����~����r��lY[�1�'o�(g^B�Ǉ���X�]l�/z�.<}Yϥ ���!�u�z̒3tF�a��!K�[t짆c��wƍ���<��$	�$S?�w\]wƿ6k������OD�r(�٧7Z�l��9i�muMZ��6�p��k��+tY��To�vW�xz2�sǉs�0�$�ӷX*��;͇}ے$��]Q�o�2�[��ݳ�OF�㜥y_g�� <ǽA�
�,A���Acc-%AE���QE�QQ��"�b�X �*�PYiA" �Ȣ�*��VH��R��H�FEDe��VJ�����f��������V�R㡮�7��g_P処��y���]`���E�������B��/��X������[3];�ڸ����z7�B+�Q���ި�qޏ�vXJ���������tk0I.|t��k8uwN�c���o����b�{�I�V��H�"3��]�N�k�cHv<���[�q	;����D>�rZ��p}���E��"T��# A��D� �@�0$��A2�r��0=�2Ҡ�����^�����7L:g]z.����񽷯7O�N����7��W+~�����͠F����2���Ov̛�Qbƥ��Xed�2�pS�U>���3�Q��m2�rd�#�f$��  ���3�&{�oR�9�+����b��L��թy�\U�o��a��o1��޳�����쮈!K������CmΪ����P��d��[��p�#:�[N\��=I_��jE.����W������]y)����N/#B��C��p��׉@�OR���ٚ6�v�i�A8
����՜a���+YY+T
1�`�$���aw�LM_�\7��UZK)D2�֝
����n��29fO;��WC��b��Vb@LJT*��E���M!t2�lsa�C��/���̽N��C\,m��F�;��9�nc(��1	Rc;�y����WVR�ym7���Nâ��xf��<�0���Q�i
�%�)�t�`h��AQ ���.�r����r"�[�%��*VH�Ȧ�1,��Ab)�X�#N�ÉU�rRi�J�.kn�6nBh���>�>��;��KJ�`35���c����B��w�f�K�Q�pA���ѧX��+�^��kf4a���տL�ڢ{���xo6x�W���G3��5ϯx��1�Q*��Z5��Bպ5��E.!�o��vw\L�FE9ۚ�,0|nQ�6��ub��U���I55�1�F�7"��N[�&H�?W��LD�^���߆��f����1�>�(�9����]�L�ׄI�;;2Q	*I��p��;Ǭunۭհ��k�sjG�u�m���Z)�ަB����h�o��M�k�ngiu���t3�^�@;HokR'w�ea&w=���IL�/2�r��p	���̃9��{uM��[���>s4�Q�����u��N��0�kB��SS"�1�49jRu�T�DN�j�f�wQ�)�[�53&�-�G;���t:�s|C�ޗD���7�lc�����ݣha��	{ΗY�S@�U7����3-nV�yo+�xh�B�v>�
HoNCv��(���+;e����m��V��C<]�pbذ��o���N��Fh���b��6�\�6쾈V�ɼ���ˮ��u[=��VŽOc�5�Fެ�շ�6t�Ѽ���t2IYv�yV���`db=�=�)3Ae*]�y��@N8ְ$J_#�J������Du�bλ>������^7v�[�ݵ;H�qC�-��0��1e�&m�ʘju��7�s�߇IR��/�q�0�821��rnk�Uɦj��3�΢8=w&]r1vƙ&�\���Ǡ��5J����9���}}Fd2�ܬ֊�s�Ug����	M�J���z�^�r|��u0卢�/9̭���4�̀Gt�zj8O.H��F�������e-t�h�:�!�p��G�Kp�W�����p��Or�;�U�]���8�Y6��S��fv6�܆\��/z���F0j;�ՌR������hd�C�V0��ծ\�`g���A�Zod�ƍ���?���]�F�»'�dA��9���c�Dm놌xN?�  M�R�:��,�'B���`a\�쁈����a9x���
�o����"��^*�t�fns�oM\��7�����$�H���!���ڵ,}��7�ii��R(����@��&T�����G�kTg{��;F--�QS�$��Fd�&�~5�P��	l����z�/�u����ݾ�P[���s6��o�
��C<n�!I8n�5h�6����H�(��n��BOp@�nt��OPG�������<o�>�Z{�7ߵh;�\�-��h��^�S4-jK�>�
l|9�������3�Z!i[�ǵ���Z���Fxe��&�z�� Q��f>3.w��~��z�I:Ryj���<!�Nԥ�8p�Ѱ�eJ��h��[h\z�}S�
 m�����=A���$#Z��ڴF�M��XS&����k����gЕ���)+(�pݽ�[``]���;�Hu����§�5}���>TE�˨����6 �/W�{c���JE������P�Z\���X��� ���=���L��KS�����xx��R*�@`�2E�P�IR"�A�~��ԡ��j��l��gv�1:^^����oF�n�W�������2"گ�g�D�/
E�[j��-uSz
�G��D�����W�}���l�3��?~�k��81�8�Y�n���Z�?9˧�c�b�s$ሴc`[Z�ɆtT�*�mAzH�/v�o1��[`��Q�Q�FڑjY�*�A�$iQ���b�l*�,%#R�U("1��
�[FѲ�6�s�����ꂾ�#�GGu�߅��OqGC��/gD���|�����isU;�E;���[P�Wb�ӛ:��|  ������������eF�@VC[�Z�Z�D��i�y���;u0�{�-�6.��ZY�>������RB��_�����^	!�{�2�Zj�,A�K#,dRJ5�T��Bڠ��P����s/9�z'�7�s��k�;۳qЪ�fLOuef��9��'��y�3�=e,�[� tiF�>��ɣ�c�#]D�
��W��gw_M��z�\�@��άk9bU9Պqпa�m4�����7S3)�zb�%��'�+�qk��X!OG�=�a�� �iQ��׹�o�ţw�G�(�ea��2��FH8�W�/g򹡙������YrI����za����b�n|�#�qǇ�2"(�Q��$)dTb���AE� �b����!	A@
��+� �1Q�TH�D������PQ?}������5��r�+�e�AViT4�������Ox��5/3M
=�a�����d�>��=��+<��E�pZ\U��������������F��ǭ�?��2�o,k��}�V��wF;�P��K���3r���j$#��#�Ů����k��Y���Ѯʽ�7�u"<���ص�1,�߄}�~u1+B�i�q;�[���=T�Y׆�`�����hԾ��-@�q��;ba�'6�{R�1g4&�χ������S2��?��_��4���Wߥ��\|��lZ�U�j����/x �"�+�f捸�୒%���` k1�Mf�3��^G+��l-������7�d�Wz�r�L|q�1"z_z�	s�ˌҵ���:���7��0�%��d�o����໦{u�KNY�#��2*ȬŊd`0��E�A�YaTPD����3�������t������P+�{�18�0�,F����Ωܙ�+/�/�#6�Bn>���Q���&:�Z�B9�� yG}�?���g���9���Z��#<�B�Y*�qtJ���m���co����7�&y@Fr��J����]1nb��u�i� y�<���s�f��r���)�߳yE�ߌj!��Q�!I�cl�=��\�M+#y|u�օ�G�g�'E�х��e��0���#H/��\#���C��F>��I�ͽ,m}��lL6U�p�|�irRŜ%�F���=7ə+i�g^S;�%�r��g/#̚�P��+���{����f>;�D}�*0{~�T����Y��ic��Iy�������/N2�jχC`d�n�����-F3��~�ɋ�^����]�՚}�d �e���\��[$T�L�9w]<��wJ����쮐փ��:Cs�����o:_}sG�;����������� �H(��Cib_:S��Bߐ���"Z��-l����V��02���k�Or�WfT�D=��w�� #���cMUJ������#a{�58��{�_{�#���v�q��E���b�����3�t���Lƾ7s�	B�XOW�b	�C~/�A�����ꬪ��I�=��o;�<�h]��{��f�K����+n-���}?Gm���¹�Z���r�֫��Gr�}�WOd2ŅFp��މiB:�!g# {1��[���������$�D�;�͏i��-/�9F��p��up,�#oG
���7����#�H:�ތ{wp;�S뮹EL�glI�� {Q\��Ԙ�),?Y[�F}X1C�|���ވ#�^<�ظ��w���{����ŉ�G_+'f����������E��Y2
FH��AH�U��>�~�﮼x6"����@� �$-� @DyC9}�kWzr/R�����V�}�ţ������ٶc�Щ�h�ܭe@)�f\�,Rf̫`�y�o�ywRٹxr}G�6��sԆ�Z��E$#�^��̌1��qG��}�X3o�Wdu�#C:At�}�t')����c�W������z �����e��9d�4���^
��L�����'���=�B�{��r�L��SUw�h�Y��{�ޯ�a���y�|�J1G��q�m��M�㠠(#����"5E�K
���W*Ss�����ʒ�v���q1Kջ+"��}1���ǾΑZ���z��SF��؊����uГ�~�}Jv�������G�W��"~Xl;����N��{=���ⱈj�,�x{�H �	 }�ģ"�X����)b��'�qG�4$ƺ�.��t�S��^�f\.�J�Bg��y�uu#��TN[��]/W���<O�>�����[��Y�����-����)��|0�*� P��(��*��"��P{J�"�Y`0V1F" � (�RAAd�$`
*X+��c"�A�X"�1U�* O�ks߾�T�[T�'s�pF�1��2���
�I�s�����vŝGTy��h�q��^;��.]>���.����{�h�e����J_L���~���kx����#	S��D��<x퟼=�FŮ�lב'�B<���/���m	����C�8�9o`��7��*����\����Pв��xx4���>���L1َ%�W�^��+��B4�G�f�^���_$wj��οfg�ߘrGyEe�*%L`x@�]�p��F�� �tu����������q�՘�NU��g���$�'�3p4Z��8X���f�oV<f�-�R	�n�1�"�Ѕ��s06-@Ͻ���R�9�\z:`�y8:��Ǹ��ƚ~M(���~��l=�K:��oĎ��}Y��*5��'q�X"q]�L�)~��w0!��E��#I�	EEX���/���/蟧&����<=.s����}���{��/���dXh��߹���~�ɨm�XB(�b�(�I�q������?wW�5�)h=�N@.X����p�ra���6Wm��v���2G5X��q��`'5�{J�����m�[z �kwu�	+{ `e�<�z�\k�}�W�G������bԈZp0���Ɍ��B��P�Ķ�Fs�P�[�1U�
�&��������\�پ������!�}����3���s���f�WM3b#�n�5uSX�Y���A&�,���Ժ��d�L�9��B���n�y�y��l���~�,���B���j;]!��nC�;#��=�ُ�a\�*�jdap��N����1�������߹��ٜdD$��>���uq��Y������O���[�,�{�Ic��	�(��W=�	��+��a�M����p3+6�s�&7��쇫<l��Kn�x||<O�*���y���<��]pb�)˱B��p�����Acs��FⳔ���}X��%wZ���i�����3��,��o�V��$�H�T`)��H�I�H1��Q���AU�TX���Ǝ��}�v��E�Ŭ�d�T�$Q`��R ��� D�PDKJ���E@UD`�y����z���n���יac�Ք��s�8��Ձ>��������颙�'8-%0�ڴ�J���n	��%���㷖�7[�gj=�N��\:{�bV��Gt��ߙ"��G�ׯ��C]c}�F�����ݥ�Iud�sB�@�Q�2w��� '=P�	_�*F�O�p���I�n��tdx �����x�u/�H�B�w���6�usbV�T�&����%�-�@�~���������s+�?���<B���#��)-k0y�7��.o�\��L�nH8�;j�#��W�7�k�Gts1�Z�ձ܋C���{n,��߭�l�³�QDbpM�v�������@��b��LmaC=�	YXg���{�,3�8�����;жYY0x�DT�Dda"$@Ad�22,Q��ˏTlW�ZU� |�ç���c۔q]\�v���Q����h����H��u{�P]��9�Z;.���z����ޤ��c���U_W#��,?ߊ��L�ܳ���5���.�߻����݅Ejږī	D	U�J�aiihV��5���^����0�R�m��{�N�+���rs|�rJ���^���W�)�c&�eG!��eqG'5�\���O@��7��op�i�����OE��g:an�)>� � � '���ȫ=�����'��L�&�몉�^G��V吴K�y�����:�� p<lv�X�^�m��@�`� Up<}
���](��{�d����εL/�1�H�[�FQ�[=N���`"Ŧ.s�|�{
�,o�s�.9ԃG���<-�[�4ϴ�f����q,�#Q��J�7���ʻj��Ǝ4*���YX�-�Q羀/5��&WzˏH�Ɔ���*1��:�]�>�@�$���>��ڽ~-~����5���z� �U�o��Kgcyu���`��Z�x�c媛�K]��Y�b�
��i�E�D�>Yb0U"�*�����g�dF-j�Q��� ��'�I�Bh��qg��B������Դ���;��N�����/f������*�t�i���C���Ih�4+�(P���0�}N�ОKD۹G��p m!V�m��n���������
�HAMم��U�P��Y�?qv�4U����tbhCL�i�"�5Օ�8mՉ���[�dt۹�kXQ�DС�lͅж^\���M',� ���f���£�e�WMB�+GZ;K�:�˾v�mv���k�R�
[���5Mas��{�oNi:�ZRo)1V�F�& M���q� H��B�N�$QT�2�~�9̱V�o1,T������]ۚ.G3�Cf�a��b���0I�z� k�Ҡ��Ɲ��L�K�=w��X#7ܙZ�o�����'T���sB�ɡN���A|e4j���jR����ps��-���=�Sbk�kC1�z���;�sgn���J�f��������S[�F��Z��(�H�R���z�դ(���5�G��̹��L�T鸠w��t��۴�܂�������@��I39�J�+nВnի�br���(�g�0�q�5���&���w6k_�\��b�SYn����̝�T_�M/d�}�Vp����I��{&n]ݕ7uO �-V���*߁���뺦�V=�*�9ȕ̾�%�fj.oD��;�/\�Mz��V�͘7��S�U�(�U�@ٵ��̪���Zk��{w�u�˸�%��F8IG��<�:�sp�vJ�j�e�2�N:e�7w��	�:��h����zƶ[��E��-(k����u��^��k:|0�6�>�m��9��.:����c���u-sD�~�*�=ֳ]�.����rw��jޕQ���@��(v�8Z#b$�WΏV,�3�8a���9:L�+jS�Pv�Y�Y�rp�N�b	��ڇ2�4�Vv���H�Ta�D,���f+�N�����T��z�."��-�~%v�we�O�L�W9���Š+�uNo�[T���85�����J�i����-�S'M��D-I��S?��:��D�b�m+á�*�G�DˇJb�^L��J�H2	\��e���a�E嚟3��g)4T�\חhJb��/��ځr7���}p�3.�w5�&�81QʹRP������� ��Iz��Ya�'�9�Kquj /c	Ωy�&l��r6�(�,}sreO����*��Zhǅќ��Ր����m18�$:VS���r�SOQ��hV\X�z*J�Pb+�PK��j�\��������X3#�U�pgt�6��nm�0k����׵��Y�ztz�����1|�&�ddT��L̒z�sF�Տi��c}gv��7 �6�1��_un]�i��N�f"�M�t)��/����(ֹ|�X;�5���3=�l��8��ƛ�,��N�E^�Q5�wY�U��[H���@����+)�t�����Հ
�����<�����yD��V}�3K�D%X���o���Vcj��a+���/2�,�-�%
�e��o�ܓ��*��W�`k�SQ�i쏺�.xe�EfF��wd�]�ں�����÷=_bꖦZςf*�V�S.����֞kڷ�'����+"�",$H�"�W�
��?��e�s��e_��N���k�j�s(��irţ]�9��Ycx�ۖէ��{lIh�\<����M�~���T��\��58��sS12����{4x�4��7���.5x�e�8'f
�~	�<$��=�/���ȰFw�ߎ~���������l�QYiU*��EP�����V�"��?�������o?��X&`Ŷod'���Q��.��~�H"��ۚ��e�(��%����F���nd������q�kԀ�8�<��آ�Yr�¶d-����,�R�$_X�f�m����c�W�{�JY��A3]0C�
Y��}�"9�ݙ��.9��t9�qE�:b��j]�\jp�`-��l��勗���Y\qVN�!W�x
��Fhb�8��x|60���QaÝ��K6V���7^^4��x~�k ��>d~���H�_r�W�v����i	qd<���PQd�9�ٯ�S���<�{���b�C�O<��qP:6�Q��4N�H��
S)ṙMic�;�{�֊��{Y�߹�����
@��!˯�I�=����ga���b~�^{Ļ�w�Mk�ћIȦ�4ҰT�g|���tA�[�n/O���庪�nkx�����
�'f�H�ޠA7W�><~�=7+u�!t��GB}�D�A//.����Ь3L������(xoq0�$\��S���h�PV͉��֡V�OD���ٳ�n�V�FK&ge��_k�9k�Ѕ���ôƕ}]=��T��iM��:�����,;�&�ԣ��k*a���O=�+�BM���&�Q�&Ǉ}�|����-2���u�z�t��]�9byq�款ܔ�b>ͯ��ޢ�'J#��q4�W4P�0c�4�4����+���i:	b|�W�MU��fH��d�B��4ט�� �UD )���@�BeA`�{�=�w�n�}<�T1$�t>�ukA�u!;HD4�և@F��/�7�w��8�=�kd53�uc;��V������z~���)/�0����3�����
Q�B�u7˘6:�1�.���:�s�!�@_Ucu����^�>�8��vwD�����Y�=�׆��������:>ͷ��^`��(c$�
�xW����&?<�C֯;�~K�w�PdQX��B"�AI)QU>�}��{�~߽Ԥʎ�9|B���f�8pu:ޡ���+;�;{}O�����b�@۬.n)�H�Q��Iw�1�ޥ�t;(��ܣ\"Ӹ>��f�I�~ ��K1	��~ߣ2���piXۏVH��[������M��w�daXk�/*���,zH�C��=� ��frf��]�L6
���6�廢4�Z�l�>j�.�'��^<ފ|�^��;��zxyr�a�K͋�0�.,Ď���&n�bg�[g�S�-�?q$@�.\��Nt�(�ߐ�Gʳ�+q�����y�HȯF��b�8!�jt�
��y�a^�b�AY[տ <���ߦ:���� �C�k��i��<5ț,n����hvC�����ك;�Æ�`�+��u �#q�8k��0Rĳ?me)��1�q���B=1_��ka�=�Fڬ�^�U���$\Fg^��2�w2�Y��T���nN/3^��W�J
2�F� *�R��VKh��}s����X�w��_�>T�VA��xO��s9���퉬��C�]l)���ֆ�v!Y�̋��ھb�IK�2v^�N���]d0f�U����"�:��6���A�E=�C��b���(��΂).�9(��,��㌧R�֧B����lv:�؈��/��=;����|<=�WL�{��.�⻍VLoÛ��&n�9r�,ڿQ��<+�`�Y���ʙ��#3St.�*�d��}R� �}�x��`��DdX,��U�"� �<�'�x>�*C�j�h�E*]���Q̾�y8
K���#�
U+��	�I��X�i�^vV��1[��T.ȺC�l��=p�#O��ճr�B�a�|?c��M���Q��߼_C3��ͳ�j�'&v�����T��֙��N�c�#����������Sy������[��"IGw��q��js������N!�?���cS/#$Mi��0�u��.��`e� ��R�=��1h�����lP��M��W��{���od�F1���H�*��I���(V(�������_���uW_�"��Z���T���D��w_	g��s�,8c8�u�@�O�ʿ�CaxݨE�nxbŉu��K�ent��iO�N��z���)@��
�ǝ}\ ���,�6<<H� �3L�����ץ�RV^���Ūg�1UGz��<�MT��g�L���o�E3\ҽ��%`�v�a�S=��>>��>?Oz~lL �x"o�C7]��7��́HA�R���{�xB�Ǖܢ�sW�u�
��I�s9�H���
������V��~q�иF��p]mq����}�K��)�������Y��D5�#�K3�.�d�������=ƢK7�֊�47jD}�<�B�#���EEL��q����usX�V���ݍ#�,����!���Y�%��H.���$�s��L�F���B	�Q�L_����x:r��Z|�0Y�LZ#�fu��Л��,pEGd� ��m\�SP͙�Y�\u���~}����c$UIO<<	 �N;:�jj;1��D,ؙI��2�I�]t���Lع��z	����8�=���T�a���Mb�E���O	�S�Gb�D-iZW��1���̭����r��v0��`��6sh|D�Ƨ~~�V�W�AQ���A�I��(��;�/�ɽQN'���-����{=X�I�bo�D� � �dbE��g����~O��.~���������BA�*ۦ�)Ef�<��\)�����W�d�mm�}�/иN?K�ӄ��6�?m�
/�����_0�a�/b�)Fj���
�z�V�Aྷ+��qk��]�CW�C[�.`pz�cv���"�[4n������ K����&{����S��"�j�qmgE􅎠;��k���q���w�3��ͷ�ȶ��г��UL���12Л6�ǵ �ќ��L�B~ܗ��_Z���=��=���_U�G���
�wx����E�@ˁG�ɆWo
J�*4[nl��l\BP{�P�I��?{��c�W�r����W���
�[P�b1@F*�H
AHb�R,+$�B(����р�Ȩ "�"$EE"������]�}�����������fuZ�������9�����Y%�#�{�_>�[٭Z"��+k��w^�z�ط���̝�fs�`�,
%K��q:�yy��uP��g�_/�rWo����cǗ��ĜE��y�/E�d�����|�q���\����!�禲2/�@D惊���<��M�PVzYhn�c����~|����{��]BK�C�+J�Z2S�II�z���rbˁ�8�P�퉘�m��#����G�M�;}��>u��z�ad�1�Č�@�^ǽE���w��+��C;�{�M~N���r~Q��R�V��?�·
�C��_.�]_��HJ���;�)1���{r�WRz8��.tےL4�h�������Ý��������g��㽥G���<�>X`զz�W*�b-��,��g��kKS�#�q���@�^H�b\S3\�1�> >:g哜�AXI���{�?m�M���A��Wr ��#KJ�T�Z�+.��_f�����Eo��gC�z�;V��[}�l�����.�Y�q1\�Af��Y/`7��~s������7	"w�+4��Ƴ�Eb�0:E��t$ZB�zEd鎷>�����-�����XN~�:K˯��/�����'�е�����ڌB�h���e(ˉ�CQ���7���/���Շ�Ɲ̍��r��r��xz%�?x����ű�dpY�M؀�^De�=R��KC�3�V�,;����'w/z#�a�A=s ��Zٌ9�>����{ǏӘ��2����@�.��Mg\	�-߶}���b ��tl�P5=^b�޸gg/�������F�F@��g&G�!�}�x���6��;��~QU��KmvF�.�+E�S,4(�`�'pu�+a��,��  <�\��m!�X�!x+��k��UO�-�����'�U�O�[6�WF�E%,����xC6[`�b�g�9f�u�V/,��B�Gc `j	@��jY�lfgR��2z�c{-����w\#��%<��.��aڇ�eǽ�E���N��l���x\�GOFt
�@�wzo�0�M�(+�> ���_DA1�#��Z��*`�=��9�8�N��J'!��V���ttaC����%��FG��)2<<:^��ST�ZC�{�� F��r��t3�cQ1�����f��`���5��U�x�gD�&�b;c�SP�/�1��agy^s��.�70��/�T��֓�(%��7_�Ng�:,v�,x�ʞ5,CH��=��u�y�eؚ �]��=�V��+F��͕��������Hf���������bMa��TgEd�*�'�wE�r:VZ%���@�Rƻ��~�;����ho��
-|B�*j'����ELT�a�Cy]�g�c��|065�4�`�)w6
�	�k(df�9w����T�9�Ӌ�m��.%D�Bb+���  RH���X�w��o������]�5������g;����6V��.Q-���ۙ3I�:�nK�M"�(�_Yʱ����U�E����|Ei���Ks�-���ذK=jY��X�&Ćǎ�ټnV���㢙@(qV�.�Wy���6o��<j��]�Qe���.��(k�ލ�E�5���[]/�*!p�.c/I(���`q
�%2�p��Z� �c	q�Ӯ�!��Q�k�َ9r�	c;�3�%�
��T
�na��cN��;��n���P�+�d�s��*v������#�-%��=zF�n\`�M@9,@1 �p,*���#J���^�Ҋ ֯3Z�]ffTSIfA`T�ˌGy��m�՗Zɻ������Jc�����W�;Ͻ}槐KJ��k���V�l&%�k�&�.�7�f�
�`�F0Awk�����5����!�ѷ�;�{��<] �9���C��͢LK�B���0�h�a�}�4E8�����R��ԗ�̂ mބ��15fz�m�����}NJ?W/�(U	��o�}�is��Ժ���:Tk~�U�n]<��<�2 媋C_���|�Z(ElGn�f��w4p���Q�=��Q��SF�bU���8�7E�m���)�i�X㐌���w�j����LE�x(���@��Q`�c�W�p��T	��^(���׃�C��4Z��y�AS*SY.q�ZZp�O�	�c����0{�S��W|e��c/Yq��G�;�x�Zh]��g��8�Z�<�;Q��mۆk;��Q��Mw]#�S�e���sܪ�_�Y��Q��Z^�I��Q���$�1�����d�9sd_�}R�a�b�K�0jtlgP��m/���R���9���-ckenɲ3Y�[˓d��@ Sue��+fE�jG\�l�(��j>P+���Y�9^޻xĝ�;.J^v�j��"�=Ҏ>�*���DKGMq�N�����F���zW-t��Ç���J��yW�=��`�B(L��F�9�ę��Ө�w8�Bi�U�t�G��0|rvYA<8�=ؾE	�m�Y4����+O�U�U�����N*Z�'q�sn����6�!M���M�y}gM���R-���`3����ϊ�{��c������������V!�}˱�
�da����Kw�d�ͺjȈ�yH��ns	�Nw:�g��uٗ}:l�%q�8)�3���y2$��u�^5�c2V��٩��e|��Q�gl|�j��X���8���������k#�WP�wso-4�A�hPL�D����9_b2��oB�^�%w�ס��[�q�����S���ɑ`U�TԖ���{��c��@����0�����ĺ�.���7/�Xקm^�>^� 7]�-�n�1�� /2�N�b��#7��4v�e��Ū�iٖ�2�E+antB���$J�=����+z�1�����PLŕf�;kJ̆ i�(�j����A�5ף�..,�ޓ�h�	e�Q�3��lu���p�h_*�3e�e������tF(Ya^��?Hg��AD!+�"b�R(��1o����t���
�$�R�{6�#�qK�n�c���GT�[�Hѱ�k��zȦ�D�&���om'ϭi_i�}To���2��ϔ�����o�J!�}�c��\�[�C��̎/j�Q���k�e�t)#g2G =��z�Ǧ�w�m��ξ����J�=d����	ލ	f�{aA�����m�tE�����VC���z�z��d��fBp�>R`�F(u��>�wׅ�늢�.u	)�0xR��?va
a���c�S�i���{ ���=�X�v�˪5�����7�z;��0��q�>/����n��&�j�� OBJM�Z+2�-$�p��4�>�z��Dr%:�w��u������G�[cE��o���i��#��@�I�{~w8��s=�~�1�Yn2�y1Π��zFN�Ѵ�S�\<�[�~��>��MZXְ�����Z��
jh��)7`yԫ���~љ�ў����*�j�V咙s ��sҩ9p�Et�Kª<�A1ȫTј�\�z�!;�3�}��2�n<O���"��Iy
����]������ǥ�5��A#_��F	b�':�����pGXVH���-�"� UmiN�
�v�����'Z�Ge�>*As����i��W%O�� ��G��=�d�L|x]���F�n+.;��-����ڭ�����}኉	AE	"����)��e.e���;���_����q>8Y�Gsr�W��WP�j�N<uty�A�v�yVp��C婢2�EQa�g�������5��]f}�U����
����7��`����	 ��j�mM\&�Kt�n�������S^��oU�qP���\��עv*�7F>�j��? -����D���Y�ɑdW@���u�w{nz����d�u�ZV#����d�P��:��<�Z�>�u�6"�V���*�
I���T��A?bDn��ڼ�0��zlՍ��J;����N潒�b���jvql�ڔ&���(�����R�5�wW���:�v��	�H�9m1*�:pH��T��u�WԹ�
X�O﨤��f�h�y�H:A ����U;߳�3Y����o���L$�_����w�v���zs�JL�$6]�%�J0��@A�2j"LuX�خ�ft9K��;��c�,j���Wg翿���N�z�����F�uj�z&[�Τ�4>^��_��/�ףE���KǽS^�9q0��VȜP�"HFsRJ{��	����g���f��z�u���$��$XHq!�i���������y�>�󬛋B�q��qG�Q��-�X<��x|4#tՑ p���e�F���s��՛����εd5E5�wn7 ��m `y��/�r6qF�8��=�*w##��."�[��2Qy��Vu̴� c���(Z�6>A���][����ݙ��Ő�jFJ�#zzf�G� �
�G��.��E��7qPC/�xӵ�������~�V�#ņ��h�_��7� zƜ\Na>�0a��ĕ]��U�pz�j=�*\�z�(j�&!؉����O��!b�}����}k8!9L}�`;q�M4_���\�'�.�p��S{���K�[�w��r�t=� ��!H��A@  �������H����\�Q�Az�"�W� �)�>������|i�!���`�D�a�`�4o�F�]�{k��Y�=�� �IAv\�5S��u���g��5qp��5>[�Km`�DaU�eB�[j+A@k*��kPPbDiab�bŅ+K�����b� eF�YY+V1TX�2�����im`��-���KHʬU��Y~4E��r�'����d}N��9�����r�mN�5�X$�N�N@�������fP��]�����W��J#��/yf��8����,/tB���G@�P�C����9���&uq��� q��+>�܏�ó��կ<W)��Y��6�x֯T���j%��!�HlB�T�����&9k̘�G��rhlw�Ӄ�+�Z���:~�5�6=�X0w�C�>݁$�V�p�F�<���^k�o�<Ha�(�8�Q�PFtF|<��d�#*#��L|�{�vf���+!ۂTiC��k8td�Z�z�t ��=��R?R� *:��{� a�xJ9|�˲{�
$<~��������M�"e� g;��f�u�2gJ�׋� v��;i�:w���W]r1,9�ECs�n���V�@�x���?��ɤ�c��6��T|�HE�5wF���\�\����w�X��L�l�|8�2̇��]���s^����8�@,H,��No�g�7O�?z�+��N������<Ӥ�һ:����L��w3�(��2��H�����tV3$�E����ї4j�/�uhc�d$�(�ni��[O0!�UT:��ф�l�l~*�]�!���Ilz�yg{qVx��S�r�r�cx�yB�F'5�|*�0l�p {�`Y#��6�Y	|��*��E?�4�m�-���:�E2ڮg�T>�tYNz�k���p�Ŭ��h��E>�z�1������}�T��y	�N��D[e`�)#ǂd�|'+��C�+غ� �|�������]Z�̿5A���^dpo���5V3�o�����X�d�!@P�Z?�O���I��Trݽ���%�د��7˲`[C�/ )��s	��Q��8+5��8;���	���.)lz�In�%E�>[��ߔ�"��������*��p��B�ל[�8�T��#[���'�q$I�GFq܉f�Ɯ]�	p���KB�_t�
���W2�M�����~�=$1F,���D�R�*�A��2A@��$����TD�w�}�W~x�6�KF��/rA���u3|V�M�:u0�9`�<���b����R�eC�~dvMOgmB9������<�ƿ1|U�b�*Q:tW�8ݏi��{�od87���VW;bN{���qڿ�}��ڈ��]{i�&�S ΐW;s�]������C��0U�f1o!	A�Rq)a�E^��q��tV�p�ϳ�[w�>t��E�լ$�"�x�G�)���O���s�iz�5��i�W�v�sGldމ�T�iC͘ϙ^#`Ի\�(��ǂJ�ova��9�F�Ig�y�ѸFz�f~G/�O��X���K��8�R����1��z�F�e���6��o�v������5u�yߧ@T��$X����E0PV$,���� ��dT��HĀ�
Kw�V�7���;n�}BA���V��T�Z+��=�<��]��t�S�w+2�|n��a�Xh���f�Ǚ��Yk���-�޳�F�S�U(7r�P��GG>�^@$-��\MǾ��z/-��eaX��-�!(��G��;|����6�y��λ
��r���5z�h.T3-��7q����L�Sh`T�6w�ܺ��H�&2�g^j��r�DW!�ur��~��K�I�����=�yT�7	G/+�>����PO�w��)*<� f�-��K�y�R��U�t��6����0���Tu+LCN4�) &~p8��*���37�h�r��/�×ʼ�T�u� Ö��=n��<�0'�L���5�#39��]��D.8l��c��"�$X# _����\�}���9}�v~�uI��;3��X���t/E��|�RƦ_NBK�u� 8P��׾������5,qv��k�W�j�{X���k<�Z6��V���Ꮮ��S�F������,X��q�r��D��4�S�����j���tRM����
�L�	�=K���?(�Law��Dڗ��˦t�M]�2�>fH�j�Vu\gtA�s��ȗ@voy5�4���D�Ld�O4_ ��o��Xu��h}�nԾ!��@ɴ�i���WN�o�.��!��N-�_U�|7�A{�lk��n�|�z�9�����e��V~6l�S� �]�mb�`�o��/=s�<���n���B��4�!}�Ǝ����O\G-5���+����|3]���xV�l9H|�̎�1+P�(#�b��2�V��F��E˿wZsϧ�i6HZ]=w�����5.���ݳ<��~��}ʯ��qI/����#C��&�����\ͣ�k�gݚgZ��t�m���N��2K�qL�sRZ��D{�G�x�{��_b�|�� �-u��g��/uP�XxO�85)U�F�&���"�Y^6�t<��7���P�A�ݓZm%�J�yFG���EB/n��L/�f�]�p�Dѷ0���݂�Aqf��Ɛ������#qϻ�f���s�A��e(���j��� �}���x�H��}�M��Q���1�X0��:�a�>�6��\��:�U�|@��ޙ�9+]Rk���.h��Į��멊�R�$�@�sgU�q��:,)���O�$V�����v����b�l�(��_z6H[��)φ�9{:/B����V�ҫ?xFGj��{��]�W��QZ_"�*}���ä���k��Bs� ���D��,���N4D�Q%<�U���U��g߾��y����"�H�����D��lh�+���W�X��?������CΧ|��K�)E_
TWP:�ԅ����5��V7�&�OcǬyJN+��u����>�X9��I<W���'xV]����_�:�E1���P��R=��5�����b�W��l^dL��u���
H��Xc���e�+ڽho�9ȧA�`�c�4iU�����R٬�S^�����)y�^��(.<}���s���X��e� l�d�����r���>���L�L�^�D-�v<�W覡��Fap
�|z�.7���b���w4'{��+7}�w+*TJ�#F�.aM��]��v���q��NZ��Aِ	��R�����uS�c�tSՕz!�BVԭK�̨����)l�ZR�q�1���D�z�ԧ4�-���LF��]YI�9tZ�c�ַ�(eܭ��s���=lQ�ܘ%qk�C��֚�M�ތ�3^aE1*��W��7��յ����(��n�46�.���\�^�1��g9k�5l��֋P�Uw�ŉ�\�
���kLͥQh�٭=�1ץ�m�CTJ\8ٶͰZ۱�cK�289}s[�k��q3@��E���q�1��LG�0���
Ns3^B�8�f�;���Su8B����)����}B�(�A�W��x\��8�?�RSc�TI���K��F���, �*Q�h��TQ�_J>����\��єۆ��	��y�o7��\ޅ}�x��@b)�8��YV�l
ҕi�h���Bٶ@�ECHH�V�V��%���t?oJ�/A}������a��:z�Νe���6�6�>�r��7)�2�=aQ=�o���qۣj�x���A�x�t�{|ҌLW����-����N��`Kx���N���ou63r��S����6H|0(,k��Q��E�ʲ�B�m��[�[��Y�c�n���t���KwvR����̺o#�D%���.dRX����n�j�ן���x���Q�U�ڙUe":47$����ee�4٢i��S�-��/*�%Ȕ��M���b���	Zв�
�鵫!=���tK�[ʭWf�Ս�d��5�Z W��un�k��W���{�Ό���<��nғTC�e���rݖ�]aHT(t�]fU+�G�	%�X*�p��Kr\���M/]�JW��պ�g��pb;�Mt��>AQ���KVV��ǰ�����n�8�6v��܁�Ah��>�����V�%�nXo5�*4��� �U�kB��٬w:����,P��[�f��� ����z%L˃��9���UY'a��ض�t�r�	igd�y-��t�	Y�u��W΂4���B��U1f�y�tx^s�j��E��ש��f�.Ld����-�dWN!�7�8��Tf��_]X��I4��.EO	�Zf@^NE=��;`L���K�;us7@ҫU;n#�JRm��a�,c[��7�҅��&�hۥ-�{egR��F�`�_kb�]l�w��WA�)7�D��*l���5N�����l���Y\�
��!��̭n���|�N��Ƴ��K�$"u��d��!+�|s�fh��9^�Y��pSY3����  �O��a��J*b��G�!{V�ڵ�*���&C�*���IW�sN?Q�7��`��l��Yu͕ҋ��J�㯡b��\MB��]�_G���zc�ۺX�l�}������-�.*���Z��v��ۙ�������O���v�,��]N���d&���� =�� ����tRoVׅ_�?V��������,	�H�%�#N�%�N�^���)U��sf)Ֆ��A�Ｎ�!?��G�!D��w�>kej��I<���T����g�z���^��;��8��ѧ!v�M=�=WE�y��m��TB=����u\����]�F�M�[�����s�v�j)q�+jJB�l;r8t*���gQ^#[�^��o�z��#��1Z��Mf��k=���K^����ˤSL��J���vL���G{��;��h:��]Ҧ�!���ݼm�/=�{�#�et���΍쏼$3�|j�8رQ���#��C���Z<���������w�B���d>��w��c4�h��.�pn�x_�@�`��	��RH� i���߿t���?����A]펠�ՏP j9b�0)���N�0�s�'���օ�7�	"r�j�t�8R�h��G��ړG���\kO�n6~{���sO�A5�ƭ�����aK�9��[����1u׬�����Ի�a��p��a�sH����=b}j8����=�t(��w�`��ZI,ʁ��O,���:�;�^Lx�@�U�G�%쇇�Fۊ�(��r�Q�����_.>_���
�b@�������be����|
���3�=\w�8j�����T�ӆ�  )��X��=�:	����"��UE._�_f����_�`}��6�� ēL�@���H 3�˙ا��n�N��m�̺���ܫ�3������%�0�"�-����Q���x-�ؔҲ+������>�&e�}b�oT=[��2�׾ \��:m�e֙۹�\�ٜZ{t-"�'������\�A\mH�����J��V�Ӽ�
���:��w9��u�]ӬV��z�B������zd���e���Y�n�i����rcc;T3�զ������K�럴(d�(��n���g����-�wt�&�j��t�y,>.7�"���Ɉ����)�������}�+疾 T��0TW�>��y��4�Ή9{һa�6�E�خ�5��duz��֪�^�,��2?�6�9�7�B�h�ߏ��������������g���v������w&�ƕ1�x� ���Ǥ�b�g5z��c��tcMEDZ�		5�[zV%�y[|�}����j�k��o0R%��63�y�@�z`�ιE�o������DVH�YL ���Ad���� ��s��[��vl��fR�[ꋫ�3�ιa�͔'g�Av��]�i]Ӛn�EJJ3��p5���*��33!ï:SȫGp�틙���Ǉ�>kʻ�]�7����f%�~.�B>��b$	��R~��5B��~��Ot���<���Q�����ey���ޛ2ƑO�����K.h#n�s�q��B��-�̉A�vE}�)3r>�}*ZMg�v��vwx����tnn��J�j���I˒:��8YLFs���� �'��޽�9%��VB�\��c 꿀
�=�/>�Be]?�/ۤ�pd=�%s��T6��$o+Ω*>ؐ���w-R�4���Z��us{r�==}����G�Z��+���b
�?>��rB�4=-wR�[q�ͅ��<+=�vC/ډ�i�}Ưh�ٱޔ�$^i�D@\����U  �M����>��V�ៗ4-X>�Օ�Į=5���vBb8<"�'Pt-h'p)ˋ�Y��mC�u1�p��߿3�j"2E�������,�TE?g>��v��[w���˽P;(�k[Ewlm�vk��֩��X�WǻH�=/�*η��,�u�EQ��/,�u}��:�o{�]��|3��Yh{܃?��2�b��p	, �v�E�:㻸��5;�R��
��
Hӓ,���},z��R2������}��%�)�'�o?��K��CV����}�@�:���y�o�3E8��?z�Ǻ;t�{�y�^���C;����d���D���|�H�¾�|������Z���Y���gN 1���dU����=7\��vBW.�S�Ā�U��I�ޑ��E�ދ�O�i| ��w;.(j袑�Q%�RUvdO�+��)5�щ3|�ҺWN�n�0���[)'\kQ�1�8T;@�������}p>���������_�΢'��xw�!��,�m*���4��[�+e��_�R�s�9�L2�����迱����� Ab0����0���C1���E����7 ���T:5b�"�
0d���B�# UdE2*$E�0En���߻������y�b�$ܼ=�O+�,�*ԑ�j�u���f_5�әu��8+�.��^�������Nm�uB�Y�P��^bɣ��s6�M��!1ٵ �Ԯ��:�)���C�C;���ꆴ:U9u�v��q?�2�@���.vo����ΠBS(g$�g:�i�I#[������V��  �)Α7m����f������ŶH��9��'U�S:�ӽh�ܷ=A��X�d�ĸڀ�;Oz�])�r2<���bE��eG���ڷ���jkS��yQ(O/�#����՘�_@�'m�=dc	u�;����{�{�>[<�M8V�!Wy[ɫ�r$1eι�Q�~���a��N
.�o���������Ť�cS�A��yP#���1�;��h�\K�֧eUlˎ(`�<Z�l`��$���7 ���o}��U�y��Dm�EM��${�=#�5���F�\x[V�ϥ@�4G��#�B$ �����E���!P|��0�*��V�bt2���Z�x譶{-��)��E�=�E�㨙�Qf�n��.�d���c��Z�ɕ�>�N�__v���u�Ž��q���$��x��z�1ҳG���� 6�z���l�!���"�R��nDۀ�}Ɨ1�9�C���Mξ��5^b�a�s#R�7r}M����x|�/��dC�]s0��os��SU�{���-��}qp'�30��.�q��k���z�>=V0B�dq0vz*��#�!�����F�c�[��؛;H���{u$ܪ٣����/`���"� i�}�����3Y-)Ҍ�c�"F U�������Ä�`��}x��f~U��X9���,�|�������'��sP�A+��a�T>��7;}#���Z��x���  ��zwW[7����Q��k�(4���!N-�k��闊�o!�I@Ȱ滦h��H���.�������}�Z�zk�E��Y�8��}��7WӇQŷ4���yǳU�fN���]Yg)q��E*�`RM��:���K
b�W�f�D�4l��Zsx��1��|C�@��Fhlz��h4��m~v+0��8�V9�j��g&�H8QegOuC��!k�B��r���ϼ%���x����wx���B�c����N��֬���q��ܪv,j��-l�y�md<K�A�*1�R��BX�Z�~���F���Ԯ:��om�����Αfi}7�ߛ�N�:�R�f�-�P
��w����)Wىhb�_s�eXޢJ���p�|=�T�[�_"��᳹?5��O⋷���˭�-N��l�|�,�$��Z��xX�p��Ԟ�.�9V��D�Y��v�\1������x��@#_Z]����57�aN��,y�M���\�j5 =㷲�H {�r�B���;5£!
�[���IP����������i�������Ϯ�x���*2�XT��U Ɖ���wx:s��v[ڗ��k�Ū�PyO��-14|���0ꆥ^U�ù��_�Iq�=�/7����;�{��:З�fwڕ#�:���ӖP�:P>�����{�Gq�GA�T�Ս�/}=���M�I��H����Ny�޹�����&Gr/�'���.��&�`P�n��#H}��!X�Җ��*�;��yVo������np1�a�s��H&.�r���ܠ�;`o"'r�]�W}%�5;Y�%FTq����R�=��E*�?:#{�O���;�)��Ͼ���YPX�a,Nv8�M�WEV�tCʽ#�h+�,LHNyudm���_P���ܭ/��s��d�H�Cs��.g�����=��s�f��Al����MK9{0�o�S�o�	<#�ny�C�M�hucpt��
A!�u�[�N��&�� ���0�&/6Л�7Wީd="��?�P5��Ǯ賨f���E��@�� ,�߅�w���3&�R="�n�9Pmr�
���Y+U�w�D�%콭��%��)�&��nC�O(�n׊�v���2&�t����:���c�������~O���:����1�H" ������y���ZS��v���ڇ�;�j7�5hc��P[��D���#�A�:�:�xl6c#$�_s瓷1���q��l]D=���G���Tee�bT�����^{�a��R�&R�u�]N��b�"+`k������o���D��]�Y�Ykf� {��8x�����FH]l�5=R�/D�>g^�i����2��s���{�/C��K 뇡�}ݸ�";؉�^�� G�˯��J�3�y�j�~����W>^u=���{4K��+QQ]`[��7�d�7K�`�D�{��'g�m��`��c���d^�O®Fc�&64�j4<�KM0	Qm3��v��D2��m+3��{ԯ_:Ag-҇���xly���S����Gl���Y�7�\��6%(U�ao$e�@~��0�m:	�t�S_��i�7����e0w���s���߯~�A��G��_s�i�7��fZ-i��0ݰwi!bՄ��:���c��_rb&��kݛ
�t޻˽��ӣ�m�Sp��"�{��E"�~�L��)�8���(q���sw��aӿ�3cY�����t���׹yu\Y̦�s_�h�=��|�&0�N�D���)�`�Ù4u9��Mi�b(���M+����OYm&�t"�\�1$sT��Qu��}Cx��j����_�P��~�X�e5�ϩFm<��sz�"�1ޘ�[
��ؙ�~��
{P�f�M�+�$�
��t�V�v���m��\��i������ԙ����_!�X{��QB���&�HT�q+f��2\%�*��T�����q9*�V�A�3%��l� ���S
4ÜiVbVE�j���ηya\��_wssN*�h��˴Kg�9X�m�"Ї]f^h'Dm$�p�禵Z���}XX.q���只����\dWR�J����lD�a(�⥍�֩F�T*L�{Dɏ���km���.���ζ���Zpe����`�F�Y�Ǻ����q!�$^��AK�5��!=��i��mŘnH7�] B�<��3XI)ƈck�d�j��M�s��v��7K�ɔ��L��2IY��J�6]3Z�J6m1s�$��k!�\+Idot��j��kI�6(����˾�B�McCFV���{[����2�ma��t#*p�[�y�U�[s��/��L��t�a��xq��+yeM����"�	3�i��a�]���ö7m'�8;�쨥^�0/�9W�Ve�IMM@�ҙ�v��Z��w��I#ڠ�X�!̙�y��f�:LVt���t9Pc�e��3D�_+��/Pp"	S8�kpo`v@��x���~�!�4Ad��N��ug67m"�K����v�jU�󼄶�.Mj-�;����ӵ]�9V��/���35�Y��L�#�ޛRU�#��q����nB���]w}�s�u�(����S]� ��4H�=WQf��9������0�d~�Z�VK+�V��3u&�k�L��]T�-��ȉw�g�5Z�	��RL��u�t6)��Wv�s7L�	:�B˚���A�5�KW^�lLkU��q�$��g/���qH�v����NT�in]S;�ȭج�7]��T�e��!��h��.����ݜ�Rj���#w���K��;e�/||�ۋt�m?(��=�SM@}&S�"t�a�7���Zs�l|��m�VwĆ�49F��j�}��rw7��yQ���F��&	l�������\G%װ�#�;����͵���S��<�C���a�z���j߉�]�B(�����5z�8��T'�ӧd%T��o�y�W�w>���P������3*�	�P> {�I�{.����`���[�Ү;z������\,뜐�5ᜮ���������+�e��RDQ\���#��#a��?Ik>^'��Kx�]�Sm�@�Hզ��
3���T�%��h#!s�M@��n�+�{g_�OwGk�[�Oޟ��<#�q?��?����_�{��� |� XHG�����"��駕q�]ON�ݷ\�R�m0�q���0s���&�����:q�$*1�6aÎRs8w]���������ۨ^�jv�{�D�����ĸB�:��b$�v�U0vj�]X6����g����2ص��l�Ͽ?�g�o�$SD��mxE�!Oh2{���g̞!��|�C�mj�]=ucEK����a<Zȯ�\���◲?fX���3w �̦���xD���9
�%�â/�5��{��y��3^]kUz���t[	f�Rv�z޴<�������������l�|�N1�U���!�i��]�d�~�¡�ud�rY�Ð��>dº�#�L�.�`���<z8�.@�|k�/��ԾY|��.�DX�iC�L�t��W���:�fˁ��n���_;<+Y���`�?O?p��{kԾ�t��0'�X��9t�d��"WH�	�.6�f�؅Q�>s�'��L�!٣�I@�����DPE#-�+*"#��1����KQH[V�TQiedb�U,�lDZ�E�,�����ʥJ*��Օ��KZYB��u�3�t[�Ӝ"U����yo�VS$J�tnW3V:v�X]���K��b�;{w
�ZT�4Os}v�I�����H���+r����8^�s<E���n[�s5�0�a��i~�_�w������ D$����F���f�Y���������֘V��M���()E讕���f���RNPh�'~�xQX���=xB,rb>�7�E��m]s8�	�I�7�,al'�cb2!Jo#�%��x{�ቡ}[�M���航ع`fО� |@�'�=	�/�l͗(}�r�6q�๠r`1/�ɋ��ظÁs�A�غ�-G'(1�t{B��d�ƺ���V(t#�|����v
z�~�|O3��o\�*�(�2�{���u1؄��x}�}Řjx�rm�фQ���W�#�<<����W۳��x�da��.�p��ﺜ��
���ӣ>�+��w.\���ri�{�:M�=H�hwa����K��w�}�U| �B��)	�$��z^Z[�߁�[ֳٙ�%Id�ڍ^�Z���VeAZ��|�̓�T��]eѱɾɉU�m���ɝ�yܤR9v���=�|z�rYڶ��e
q�^����Ej�t.����nr�C*6s��-�؇^g9q|�4f�z��|T����}N����̪�~ދ(��ϩ�=�#�)��Tu+8-:/sI���]NF��`x�֫�w�k�����?rM��:�Ө"�t�+ؒ\��_�"(P�������<$;�Ȯ�t��2���X��d��)�hV��χ������|���9��RilV���:�]�n	�.оH9
��΋1����ݡ�ߕ�j)��޷��E���v��6ؽ�GG-�R^����P�q�[}@�=��d�_Cu���8ឪ]��	j��4�z����^�^ݗp�p��2��@ī28�<�����-���F�|D�Y0��u�P�x�(��� ����Y$EI"�Y"�X��M~�Ư�:�k������]L��/nn-w�zKY�@X�%��13d!j��T"���AH���8����^d��c5N�m�c+�I�C�q��U�q�O��L\(��"y�ӧo9h��5���ئ�Eԑ�I���Q��溁�w����TP��o<9�zrew��\`����K�Q۴�%���Q��j�@ c9��ű�L)���d�@�_�^g�_�c���_wy�嵻�Dy����c(U�׳��<�(Z���c���g�^%������P��n?�o� ٟ��o�4�WP�
���c� .�[Y#�)�w���a���F۾���{BYr%��'MF�wa�\���衊1
��+������������� ��˲�:�j��(Y �!�����zx��Ru������V@Ԅt�8��V�������R#d�ߵW#9wݦX�mR�)��Va�":�8��i��:���Q��R7�?~;-R����F��x�ݏ?o�<XE���qsv�zVWV:�Β�r�V�f.Tu�!�2���R-��j��+2�YX�ߵ��euw!k�����Ӡ��1�߳c>K�~�]?�����R)������+���uK��~̇�0�0+,�vE)�ի�
=�"�0��rsji�].a��c�z4�E�����Y���|���b�;��2R�2э>���D�r^�̝�5%A9�i35�!�ldT��gy����Mz�
or�s7u�m3�8
�f*�`�����0Y"�#"0RF(�"��1b*A����m�zD@ga��{�s���F�Qu����%��,>��䵽[� ����A� xX{]H�F�娮��������W��b�|�!m������\4�DSו|L%�I�6�3|eKƘ�y����(}�ѭ�t�,l> �;�S-�짻v�aw�>~� {ݖ����߄�R�@vWQ�/��W�X�;j]r��V����L�X��:��PV\램>�*ڊ�Up�E�<�"�Ǹ7Kj�Q�:�87k��㛺��/�w�bou�3z.�4R5��)N7��yy[B=��`麝^� $1��I�:�#7�A���N:d����Pn:� ��#0��g�Y��$���Fb�۾�J3Qx��6E�	ի��g��+����I���g�$���(�ӯ�w�pʁ__�η�tۈU';�ل�#����ÞQ�!���Ku\�3�`u��=QQ���>�G��?��5����t,j,��G �"��B�ٮdˍ�ٸ>mjpF= O��<�^�v��%Wx0M
�o꯰���-v\*�~y�ע�|�6�z��V�oGj�B�pHk�h��lvɥZ�+�.���!��xu[�
�A�z��Z`32��,�p"0J-W�92.�G`C��-ۏb��6UNM�
�!�J[=�K"��	9�g&a.������Xۅ�L1Ӆs�����N�9�J]���_�o�r�%J�4�0���U;�<8)�M��'�«r<m�?lެ�.l�W}[86���X�ѽ��hT�������W<��=4XN��d��6�]�f�Z���aj��8�t<Մ���~yS8���}ıown^:W��×G��Ҧ�E��L\�w{%&��p:B�T�8�_V��/��;��uzZ2Q�/�u�f����|} bF5`{ޠn�zf��yG�����uY����a]u4�ĸtH}K����vM�WyڴZJFwbX�&����\�0�����No���b��� 3�DT<J��q��Ϩ܁ǞL�,��._9�+=�.^���@J�Ȅ�)2 �x�Q3C��F%}ƃ I�s���C4���ȰpBd=/�����(��3�xVK���~��n��� �}���v�I�(Ld)k�x��5K�xĔܿ17�Zp{�ɫj9E�~�z�i�Y��G��MOL�p]P@BJ�R
@YϏ~�����x��B�gl���0�ۄ�w��[�,���lF�o�ˍ��v�ol�g9|y��&t�p|e�͂����m-ݪ���]�k:���߰j� �Ya:H�q��u��x����"+��ipз"d:u� ��P)�WWR/x�!fSMO-��*�{nV�4*-����۬_���`<�6d�lu(����
���-A��RI���b;�L�¶�j]�E�$+�נ�g�(�3��4��`U6L\W9�lEŐz�PE��=��덮Ȅs�(������K�~���ζ{҅B�^��1��>i�7�c�3F*:8pM*Aj�7�k��WL>�S�Pz�L�x�S�˕G���F�#�S��vfb�A��ۮ�ev��T���O�B�Ύ�q��Ce�����|   ����},N����&)�=Pԥu5=)2��$2�:Ȳ#�*�J���۞�X]6)t8�4�k�v��WZ�c�ܕh�~�߿D.��*�f7���7����ﾺ���;v����i�-��y�R�P�ػ(�gp�QS�Y�ȭ`��psȨV�Ke.��O�Ρ�,�=����{z��.ګ����n���)R�e�T����}��u_'����&�w!;ѦeJY\#.��S�O���������t��u
�4��[�6�X�B���pq�43���av�e��� y�*��N�Զ��^�_��>]�g�ҫv+��ߴ��Ӂ/Ga��)�Go�
\Z �������U���f�Y<����o:gT�}�*t� ��ß+?O\�}��+�� ���^F7���� ��%�~
�W�/�?*��)3��N�2�������8�����h��� 9�}B��� ��H��Kp!~߮�莦�)��oq����LˠOez��hW0<6��G����S:2+GS�/�9�'yR�ۢfl�$�8� z��>T9�>�{����]��0E�\��z2������j����Y��g�Q�B�T~8N�@P�����uW(��ȷi�L*�
��(1N��jA�-Fc��[vRM6J]��k=�χ�k�嶛�����!��5�7�qя0�[��2V,����<B�e��o.���h������h�wE��;��v�p�Yt,c����<w�VW1����3.,��QAX��e��	��.k�I1�KLr��W��[��
f,2�ƣ$�p�M^;\4�R�s�/���߯��P):�>�j��Q2�-�n`�n�5����u�*`Z���7Yi
�-V�������<�̬�bw5m�����T�SEfٳ�rbI���.V`Le4b�*��o�c�Wr���/Q7)�-aZ��Lu�u40!��t�+V�8��t�E&���11�EEۓK*���jd�n�6kR�}u�ßk{7��0Q���nS~�_k02��ԝCG4���4ͱ׃S_SZt��r5Kmm6��F�Pֳ��H���k���5�e�ۍfah�X)^���h�(*�M�E�E
Tf���3�N��Ԫ]Хi|Fa2iʥO] �|��a��!�DQ��D�
7�r:'ج9�-�Yȩ���Q[.��9�k�5�s���J�-g/4f��y�W��a�PV75*ӫ;oJ�k�n��2�U�,������� ��a�1���Ԅ}M`�hs@�u�vn��.�4��Ve�"����ˢT���&�;�sK<��򷪆�T{��t����QH���K�ֹ��X���7VmK'kJ�6�{ؑ�f��F�{���ۺ���\hnR�+^4e�mM�:>���\�������I*Z���� U�(��eN�Dq�t�I)���d�M'�-f �+�S|n��=9ߞ7��n\闾M�I&k�V7!J���)+��"�s����b�ִ�Z��=+>�2�կ�A�']�7�^: ��[n�rI��f49r�ga뜠d�˦-)C����w%n��N��0�O��*��Q$vѵWlQĳUZ�	�Mճk;��	Ya�1�W�� ��N)q`��
Ŷ��:c�R�wn��v��ys���³Y��)!�KV�Nڋ��xw1c�p�T��8��d��nJ0C����
Iق��`ٓ&�kQ�� 3�m�vz����v�^2uKPS��������ɋ���Y0�MSp�j\ї����o�Fh�jE�£�Uj��9��b�
4�*Z��d�S��[n�o�&Q0��^fą�`�_E�$h�����:+��^�3W:�P��<P��ú5'φs�;,�7+��wxj�T���:k#	�
�U�Pr��au�ù�t4��1Ρ�Z�A=ͅ|d۷������z��b��ȧx+�읟/ B���qʌ�-J;n;�s��F���ˠQH>�;w�+��co�h�c��*���#�T�(��Z���ݱT�\�3\"����˯f�:3�e���!R�	�Y��P�<c�[���H���bD�+�6j�j+ˉ����5�ʵF�^����Oz'd�=�
��V��B8����q�����#\I�����4§j�Vt�zk*�S\�/���~_�_�?~i��O���EV
�ǃ�s������o�=���s+��%�V
�l=^�!��8��K�on�TYCk�vg�f��+��*�^z+��ar���lPʽ����9�S_~�<n�8~ל�v��8 �k@d#S�#����`E&Ԩ��(n'�f(��� 0�y�߾���c���r@xq9]�gtFGBъ�
U�X��n'�+�(� �p6��v���zAV�v�Ɯ�#�PʅΪ�Z�1�N+I�}!dQ���+=��S���q�a�3]�J�\<k�f��ԫ`�����(�e[a+"*��E"Q�d�HU`�1UE���IX*��E�)Y�F
DPUQcej¥DU����ĨEJ�2ڌ�X�F�U  wY���^_��m�M�=�=��ٓ'We]>��ޝ�Nn�X�,S�s�)�+MX���$ܣ�]
70]�tj�fCw^),��wѨ�ӝ+ě������M&��]��=�'��عw��7У�����ז�B��E�=��Pn
��y�g��9��<��l��_�bZ�I|")�,�<g��ڏ��٫�Yގ�J0�KE�����G�6י����>
�de�>��{ݿi;�oG����
B
 �C�k��PC>{�D��h�U:��������c��=���+�0��3��bj\�}6��bu�3�=���Os\�Y8O���ZJT��X���W��k�bH����7�,�6�Ԟ�sx�24�ە���i��r�zz�	
 {�0 �U��8��+T��`�q,LZt<�%ͤZ��}f�Z=·93$���20�g������,j�Y��ǿ��s���wa�(O�����~>Ћ�J�s4g;{�Z+���p�.���[cv��6�n�Pq���o���1�.��/��a�Z?DʠR<.�t��`�C5[J&�H䤼�p�v�oM�o�FZq�]+3��V=S�*}�=�G�/���^���ѳ&�9���S���qpo�:jP���N�	H�M�v�q��a㜦L��v.�q�k���8"� G+� σ���G/�2��p�&�ۅN
���KasJHQ�u�י��1J�1@���h�:����D�N�%�ݦ�f����Q���*�_\��������X�_-�������<�A�xl\q�jn���S���<
�?Z�Ǉ��c��-�w�V�Z�����mM�."��ddvDΝ����ЉQ���]�5=���F.������])d�B�ü���9�~�Ow�Ҝ>��AEUI"
Db
��(,�$PP��UH�4w�߽߯~����q]�P�9�]�pg=�:���ܓ�i��i&�c��Aê����Ѕ>� � mM�ۓn�E�t�Hq��	U�ha���ܨ�C�$��f�O
H�:F����R�gy����][J�")��w%�uŝ�wWو�^BX�ʄ3����Ñx8�j�_i�Bg�|"h>���s=>�0u}��UP�=2y�WOv����]��~9Z*�h��b%㻀���7B��q�]ڼ�c��g�n���tߦX��v���X0�ӕ�����A�_�X��c�Bu���[��\ X}�t��B��.�[�Lw*詬����q9��Q�+��9���]s�RHG�������[���Wy�ߒ��,��Qu�Bq�ǯ�0�Md`�
{��Ƽ��t_���yR�c�ȶ�{�2lz9���	�%	�{�1u
�44�/2�t3��/�:�ap��qt�;��67]�;C]r��i��pE�����v����ߍ`�JNul��K��љ�ڄWn+%>��9j\�S7VZ�@ə���Ȟ��O��������Q篜6���k��S�F���:ڏ6R��)(��Nʷ�W�j�xl�\/������A��e;���4��&�.K��D��n:z{�h�\���Ǫ���U�k�a�z�C�'�����NR��?}�V�F7�f������I@�V�zX��qo` bGZ�L�
� \d7�91�d�^�UR�"Z�Fˀ2�[�gE�wwC���=31!״�<�D3	m�8��'�vw������_VׯvO��a���v�g��@hQ�P�7�mP�"��?� �C7�ˈ�A�1��	�ռ�����م.��jC�dY>�~�p��	���:�E_�ц��f~u�|���K/���#��8���dޠ^s8
�GMobc��Z�W��4G�}/D��>���Q܅F�8��_J�Q��p����Ʊf@[�n��ǖ��hҾ]w|:������P���:�[�@W�ab��䴽�iً��}rNչ �I���b�.�J�D^�}0��휏�ﾷ_`�;S�JO�a/����n"�������[C!a[%�� "p46�n ���F��aH��w h?#�ˬ1�KɊ��лَ����r�FlG�·�I���+�N3�c�n�*����x�hRĻj�*�;��F�ڌԁ�Q�k�t�=����ݙ�Qܨ�T�E�T��ɟ{��n���Ƅ����J��Y2^���xU"8n�{���בz���6��z".bL�*}�p�k��gTm�^�rs��#�K�3�ġS�Z��7��sP��p�Kt���Ry�h�a�I�?z��+
ի�c�KȌBM <�k؍���ON�����T�QS��@��E�f����s���_�R���:��R�Q`Y�r��ר����9��_I��;�ϳi�sm�i�%V�i�sd�Wu�S�j���(4�uή7Q-BK��r�f���)��&=�\zA=*� X��)f���Xw����chgyD� �����ױQ ��t�ad��s��|�6X�����́䔽&�/%Ԯf�|@��Ĉ��K�D ~[*M��
r�u���'_	��B�3M2x����VtqJGv{�x>����'�V[�w�.���+y2/ٔ)�?K�@�JZ�)�Gc2x�M��3��T�V��#-T󸬮���௥�|7�� �ʪ{��^	���q���#��b�p�ư��}_R6]�"!)�4����wƫq쨗,������9���1q� ��R�,$��3�{Ƶ�9�󅷛��;��l�F����*��M=B����Z���`�
���v]�D����`xb8ɧ\�ϺCLH�����XB,-�U��U���H*!���V
�a�k*��Y`gJ ��=��ȑLj��ܜY膚=�5k\+��v��^q�Ept��E��*�9,�
�z�Yl�|�muc���J��GR���L��g�n�.N>�I�Y�~���J�C�K�3��Y�@��N�':�4�5϶�n��4V��H���zn�z��������qi�.u �U�*5(�g��z���956���Y�F]n��k���G�t3���v����i��q�A�B��<6Z�+u����Ёr�uZtr�E�C'W9�[#���2���^C�=�y����?"%+�p�S�~��: γX���������\㻳Yڼ���@uQ`�K�~��8��}��K�3���K���Ʒ#6�7�6��pR�S�k%/
�<,j'���[��E���
��*��� P͇��o�W�����zʇ����ִhv�z�v�8B�������ڛ�4r��X^�m�H*�\*�W�����<�+ض�a��C�*"1X�7v�;���η�a�^26�-��̠3;�s�Z{o5c$��}@^'��t�iN�>]�N��;��k�Z6�vgp�(=��b��Ja�y��ѿ\$
pZ�͇�G��W�� �����i%+%Hr�n5�D��@�n�T�|F�B��x{�\��5,���\2'y+�Ξ���&Aa�]���5��HH]��`\����dȯM�����x6�h��ô��ؓ�_�
ķ����j���݁ɪM�������	��#k����u��	�i�Q#zn!G�w���1>���;����YԴy�}��U��m5��C��9�bx/��2���o�k
�������c�d0��ޒ��LfA<�Y�9o��<Чs׽3\�W�g �.�o+��]vg�롋�e �M�	zb�R�h1,����!���!�܍��/�xxgf����2`k=Ӟ���"���_���b��>U`a���r��3Y��Y����������Q��rţϕӽ�yb�9,�;"mJ�7�ا�pi�*����Yt��+2�WM�3�ݛ����.�n�on7���XLf1ް6�J���O#S0�\>����]�l{���z���=Lw�`�j�q�����L6k+�mz[�X�D���޼>پp�z8.����mo#����Z�{8Df�x ��dY���磕w��� u!A��8�ӥ���᫺DK{ε5\��x�\�OEǺC�)�~��
�v΅ŭ��N)���$F��V�|�s��2�FʍK�5�n`�MA�V[�e�G���D�Nnv�������8�3���G�(�+3}�������ɳ�}Y�tm�J�4z�tZ}����y��e���G
,�$�dD�˷ٖܕ�Dܲ�Ǚ0F�	`����Ԅ�I�n�O)m��8:��pbt��ze1J��2��Z|����PPd� �HQUQ�.[u�^P�^��j�b�D�i*�)�2���ei���h�՛���v��刳�Nh���ZG@����v_,ܭ?V+� �j٨F�أ�5�<�V�5�u���ТX��x�"�\��޸菻�*��*��2T�Q`(:�Kj,�i�4MLK��iZ��w6+ +��gNfN�wz�h�4h����ky[��㘎�,ln9�iD��yv�|w�s+_k}��Z��u��7i(�D�Oܦ����)���z��֨j�E()�Bj�bI��6NTa"I7<01e�h	����u�����(��S;EN^�2��U@|EUAR��U8��u���c&͖��kf���L
��Ի7v�i*B�t
uR�"�)SE�Rᩁ�
��Z���w[ɓF�
3f��"ȲbT�2��N�w1�hUb2�Z@�\�;�6���{��{��&hoV5����Sw�k���6� Q�1�����9��s9S\ջ��J�^�q4}sp+���"{5����Ku�g�J�ܰ˶���$�U\�z-�*L���'  ��:��Ն��沀���RX�lbƃK��WT���tXT7DνZ�)��5��oz��]�r�f-��N	�꜒�
 
d�3��pʚ�۵�/ p.�R� +�3�U�9���Zle@��TLQ�V��2�V�;]kAg�%��|�M�/{ls�N��B�ϡ���Ъ� S�3oa�z����mvC7���x�"}[��r#.��]FZpK�H\\�v��,ewO&�C"��a�T�G,�Ԙ��S�Sw����+�b#
0 S[3�Wjc�xh�d����A]/{h-9��J�y��mӒ�T�j,!t�[+\{U7z�]�q^��$}}�ңOqNv�J�i�T7�ڶ�J�u*��(�.D��=��:��L�6�n�@S�ӼY�3���u���'g��{���u��.�})VX�̩ĪĕLi�"�O�|�h�Zf�˓����J�,.�&����]��9C�o/cŹ2�))�]�8&h�����k7VgQt�AӪ�E�T��yཻLM�V�׶\�&��Z��J0 yԅ�M�:�Z�|aW�D-��/jA���ca��I86i�j��R�:a
��R��ҵ��CM�K:���y/���%�bo(��/�_eI�Qh�,��liT����ţl�-il!�6ց���c��W���Ac5�=��<iƃ���P�F~���m�Y2�n�IA�������9f�l��:6kM��d�1�["&V��:���E�r��H��:����Qx�Xϔ�+X�I�쬣�k�=];��7��S-њ.˴)l�G%��d�蔄{�g[EK�q�ˠ�6�!�3�i^8r��]/
7)��P�У��ݚ�8ouf99������c��z>�hPH}y��/f[}Lm��ʛ-�/�g'�Χu��ʲH�ǜ�Ӑ�g��_h��t�L���t�;kfHv`�N73Oz�dQ�"FSλ�K�p哺7�nj4~7�뫆�z���P4N� ���r���P��V�6�b�o��KK6Ӌ���T|��9���r�~�����ƍT+���3�p���=ӹ��s�� 3z�t5��>T��ܳՇ�EiG�g��F)����q�Tw7'�1q6��톹k��kn����8�Ec���'-^��Ɔ)哰�cX.�]���`��Lŕ�a꽑��<`;{�,1n�!�����
޿�$���Z�Rg��|k�	8&��7�,5��O7�W6��^7ާ\�ym��,����v��"���[)���؂ ��O��=�z#���%g�z���.�>���!x2����*4-�t8P{��<;�g����^ȓfekN]I�Nt����o�/���Aa!?=vt�y�h�|�:��5��s9����U�!��{rf1���`�Do"'�p^��:�_V$J�vt�;º�6�9���+��#��U}5$E��We�K��l�(�u�;-ķ��]�0��̂���� �t��+�[��}8l�ηl&������Ĭ��LB
͙�cD+�q/y�8L�E���	��ˊ֧eO{�ƶ1�w*"�!��{?#�>
��p?r���[#����N)03����pஏ.D�\�ߕ[z�N�5ˌ� +���P�c��7��D�;<��U}N��Vy����f��΀!�{��EԾg���61l@�z��u\jx������ �h��+6&��י�vᒱK c���#������*1�^{��YK�S�8~;�/���)���̋����#K,7�a�n,����l��=y̌dcd�~%};�<�yJ���b��	��wP�5�m�R�J���T*��)+�B��B2V���1Ub*ũE[aF-�8z��~'}-6�<��K����4�0hu��Gq�,S���C6a5��&��T����[��Ǟ�(�+;n҉m��}\oOR����3|���&�ZW
Y�O5}ok��#ʼ_��9�="�9��t��Q|���|yGգ=�NIF��]w�w���aa��:r�F��̐�^!�B�"��2�q����ws�7'�+'���L��6��"b������4��ێ��Ee��ݔ�n���S!x����xP%��z`��SNr$��a��<��W*ե��j8��(��܍O�X)ON��i5��,�7]����\a���1�u-�ׅ�� \���F�dtk��Zk�x{�d뼷4�wA��x�kړ �.7�_G��!�si�Z��ǡ��8TW���O��.x�л~��j�^P��Sq2mN��Z:sN��<�Y�ۑ��WtKR/6Q�C����u��K�}��ҁ�T���
Y�X��xؿ	|��3sFV@*j ��\�����|�P �c�Nc��7��kR�gT�2�Lg��79����^�8n2qc�+6����U��ϙd8r}�z�g-@��8X�4�Di�*�:�[Ñ�$�6Ů�^��j�/���'�k�k�Ǽ=v�I&X5�b��7�jbbO0�p�S57[.a�<����Us��J�ͦ� ��,�����jK�F���X}��yA�}_W���M����y�Wu�����Т��i5ue�ʑΘ�z6���u3V��
���l^��`��J�q,帞�Ht�n���W `�������NrQ̋��nu�z���Γ�m���].g�u�!�Z2����X��p��^�Wܧ��d���}Oa��ۻ��{����r�ev��rVQ8���j�:���o9ȱ\{��.�U-
��+]`4�� Y�>�����z�o�ζ�2UH�R1 D��(�AAdwՃjKj�ɹ-\�ۡq���7e9Cz���D�U�\�$�r%uԢ���<;�^8�v�M�@����ے_ky|������:�b��XD���q��ڎ)<Sj4��ACkDw+�[le��g�q"Z���4���k�~������V	(1`@ �Db$X�"��\s���7�8x�'ʋ�往ޓ�2s���W(<>����0:��Zy�K9YZ�����i�	:�|�L5�\�X��YjfM���a	U���5�=�n�ZfXs�҄P*�Łƽ��qF���w'c��7��ȳ�� Bi�5dN�aP�Bri��O-��rƛқ��®���v�-��,荌�JPJ�r����A��%��|�w'�ԝv�M:���xO�ZΓ|,��s6y�0D�ަ�+���h�����+�7�G�8����
L_ϧ6�/�c�������=Zj'V����{դ���Z��e#4�@�DQ$C2��'����~F�q%���7�A�~��z	�Ƭ� �LwOX��+.jΝub!�V��r�/��g��-Ցf��:�nv����=�.5���ߧ���(v��^�&"�6��:�%7/�\���ep}� �V��(QӔ����:q��Y��t�9`�7�9��d�8c޵u�MmG��ZU&ީ��&�9*���r��[�+De�쟒�"�����唴%f�Pq���6���/��#I�[��=��ӻ�W<� �E�qbqWDi����OoHX��^�z�Dt��h���� �z�{mб#"��t#(�S�]E�W:�w��A&��>�3��S/UJ�b7�^�C��#V�"	�֦���\�����	��W������qÔA��鋺}����Z��E`�!���J�u v:8ǩ𵾦��d��Ew*�d����W��m�6�����A��0toau����En�#^'AF�TD�DAX"����,"��Aa-�ČA*�\*u"5XX�z�<w�h���本9�X�mt��y�t�tp�ۦ��#s;)֓�fta96th�Z�����K��gN�,���V�L	�ޡ��>�r�Y�ۑG'�wP1������p��Nij\�X0݄�uxv���x��A8��)j�Ό���nWGu>�}�i�o��"z�_�e�"�~��.;��9[�:{��Ҟ$L`WȪ���@�L��d�����]�#^c�6h��*�����'!��>�-sZO��LOc����j�9w�)�� I�����E�f�c.X;K$0o��y\������+7m��Cc����)��k�LN/RW�c1�a�0���P8>�r�\˦�h��|��uh��e]-�r��}+��u�cP:�� E*�����B�
�;ݍqa�C��ƴ��V��><��}���v��8�)���uSw��O0�EW@���6YP��+�\>�2��(��6%��pg�uP�
�P�������X��4�i�{���e��}�c��o�m��Ya����]��8H0WvJ����G��)7�m�ī�ÛLw\���P&���G�;���d�v�x���ލԸ�*�O_pQOb��|�q�V�]�)���	��R9��)���`a���f{f���ӿU�x��g�d;��ntEл�
�gsֱ7�kM����$��&����w��^����\�i|o��&�{VO�2�G����R_$�=���n�H6�#�r�]�z.��Ś��+�
���r)��x	������Y������o��k�9�#�c�+w\[�$ҔY����F�q��Y�P�$�E8�E{���ƪ�֒鍋	���%z�Y��W�=t��֍]�kG�ܸ/8�nJ#��l�Y �ؖ���r�o?e]�Ddb�B
ED##"�$E�,E��$�}�kv��@��=����һ�D4:�l�he_N����:Z�q���X�@X�!Ea"ȉ�$D���s��Xo�������f��<�ep���\��KW
wg�l�n���[(``�k ��jĄ��lRg�^=�F�Mt�f�����.�Jܹ�r�c������U2�s�E�B7��u�7�7�&�B\b���F�y�W��7�7@�H���}�ܶ�9�̹��$ۉ��B��Qp�;�9�S!u�cա�{Y=��Xs����c��N��xUB��A`F�y'�'�q��j��ҵ��{�_��>V�+#ة��=�Z�F�V?$&s��o�x4��v��h��L�\}*�W	�F׹�K���Y���P��_=pa�Q�ܔF�4��������ˡ2*5*ފ:!�<���̲t9��9�O��\�A��\��s�S��gb�j��t�4=��zoc�C��x�'��n�F����M���E
=�����h��i�3�V�k�5b=bT�m�������C�
("TdF#	EAb�`,��XTKH"�AAX�J,�5�VJ������}cvǸ^����{ၶ�n,���6�:����������+\��P�S.pĜ�+>z���RT��'[�9��׾��W4 %UU�W�9�08����R���rc�,�{�/hp�p awG�g�9�z���2��Tl��v��Oh[�;���ҸT�V��4:{��7�M�V�`�0������ƽǗ��I�Q=����8�\�2�`-��}s�1�O2Y�\ <
��jBц�/s�@�!�Θ�ÖڈX�f�@��Ԯ݁;�"�E�2�#�ז�Q����r\Re�ay4;`�n<W�p���x������V��z<w�xe����
8�m{��"$�L<���g���v\s�Z��B�C�#|k��n_�~�nH@;����{�Xs���]F�p���ְ�e�����]#�n�=O� ��x�+K�@�`��G�i�����׈�\�gW�+��3I?P�o�b�O��#����{X���m�h��~�x���!9[E{S]1�]�Q߲Tv.�`�%;�Lc��] �@�ͬ-ֻ̱��iη�w&�c�u����%�1�-���	P
�H �H�AI �V�`HH��nj�,M3T����7�V
a�w�Iy�5P�1ַ��̡Q���������Vf�)�m�3Y�&����E����4P���3Iq�
[N�r��`jop�A;.[��0�4!�Sy���Ą�ˣVv�i�szװ��dS�5{2��lP�V*�����f�ٱ��N�n�M4�-��6Ҝ�X�Fo�Tt���CR`i!7i��C��A�&�Ɇ٤٬[\�E��X")*�2MT�d����m!�h4�3G5�z	�Ѕƒ�)!m�L���+\GF���a4���)%�ۥ�wq6fTR���i��{\6;�Uf&������!{���^��{$2bE�u�l�^�&��K�2p|�4�*�B��ȅF��W8�E�th��܄�[�Qk���.���3��rRT�B�	���o�B�0�G(զ�m�jj��[����odiQ�Ud
4�)�He8�k��FƍP@ƪ�dʌY����t��'!�( �˄��f�+��b�������*V��u�����[��{���(ا�vP���'�<7N�}���b�E��Y��;��a���w�V9�G;ɪ�U�c{Z��NRBGihV��v��y�͚˩ym�\����]��g+�eAuu��v����$���<τ}[`�J��.<�2��U�w��B�Y�eo6�H�3&�b���SIG��,��v���܀��p�W>�/����37�J3)t��'h�@�K�5JkOh��>#*�k��j��:����J�W�'S�Xw�Y5K��(X���z��ˇ��V������v���<%�h
wu������:In4�e� M�̮��[`�������kee Շ��@���?ļ|:��~�^�˶/s�FW�`�ɹAt�5��@�t�Od�9F���i����h�w!YtFPc�Z�g�8��v�@�*�>�2�٢o�ޒQ�D)��+���d!;G.}��d:5T�뒴�[���mG�v�]�k��@kn��;���J�����l��쾥�і�Չ���]�1��ׂ�FTӛ��%xF��,.D����������L��u�q]��Y�P�I�7�����L��!��t��ҧs�үDRVmc9���q���X5l&�Zd7.������{�;{�:\	X�*���[)�u҆�B*.�eZ�C"��%z9���:�
�& +]ڟm�OK5I��o6��׻����2�szJZ^���>lY�)���Yt0n`eec9�̰hN���wJ�����k����>��qd����卙��4D�`� u>�uҟ�4 �Y.B�����f=H���7u�WH���������r�o6�˿�[|��*���P���Nh�K�8�AW��]@�����=��������w���ߡ�P�XO�<�Y9�k���f�Ԭ��ӕ�On�v��5��(5<�힇A��`�i����uͼ�����\C:���CQ��N�8����3*�ttwd�X����Ŝ���2&�J���V�Mrm9�X4/�x���/�<�_K����A�q������� {��zԴ��o`�����y���r��x.=zJC���;�@�n/`�郦ء��T��o.�5�g�3�Mǎ,Ə0��cɡW��F"2��Col: ���[�|����񔀤b�����pB�L8��E��)�Z�w����Xzt47�%A�I#�ux1�y����~�οo��o�h��*�X��6,����QPU$�"���AAA`�V�2A%BQ`
H
 �D � Ā���)ic*Q��U"԰�믿u���W�E���knI.?�8"ӻ�6�zѵ�e1�2�Q�[R۫��ou+]�!9���@�K�/6@�a��,��X��Ǟ�6[~�n��^� ݵZ�1*�_N��I�9. �7���.��f���8����c=�iY� �3�Z��zwk������)r�]�bDA��!�u��y�<��̪/��~sƅ�k��2���`\f3'���!��D-ʇ�f�X�NF,w�%Z�>�M�P�
V��9��aX���x=Wk����k�fxE�� �=뙧ط��'����q�{^谄���re֘`�ۿI^�#�M��)� �p�y��Y��s�)�'�;2������7���n�
��;b~��A�w�PQ=T"�<B�L��H'Ov�=���Z`���˕*��z�,���7��o��)$=V��\TL��t�#�����dT��y}9�y�e:A��(�R�!����1�!ۗ�gq��{6�9�+�c���|�н�S�~ ��yy�c�,�t���l�	��t�ۈX4f�5o���Av�l����Ԯ�Yڹ�N\dU�O��8���jܝ]c��Mx�N[X�;=��W#M
�Ӯjtv�ΞC��
�����֔A�p�Ewf����q
�;�/�eI��yS|��V��<�7��)��>Y�{���GW�P�(Ԇ�����0�q�z�]�ݘGT�cg�\M,ÝV�WOpgvǇ���룒<�[|�;tP���5YZ�w�m��7�9~G�x>�\^[VF�&\]^��.�p�}�����Ȣ"0�DdY$QDT?��������u�Ȣ�L$Y"Hv)��,�PE)���Ƅ���zz��B�U��Ee���"Z�i��-�J�Jވ/B�Ǎ�&�z��u�Yc�ъb.�0�X{�n��[����'+R����$>{Ѯg��RI�qN��T��V�wj�7u������z��EC|"�Ot��;����)!p9N�y}��LD�������K\jr��ג�<7_������lYk*$'���{�J�Uy�d�"j�5��$}�}�A�z%d�w91t��sk;ڦ��w%2����04L��i��3�\gt�'7s�f<�'� O�F;<#�3}�]�t�����0�,��?'m����3�{Y<u��^뿳�}����UU��w�o���ϑ���۱˫�yu���FK�� ���Y^/�Fd�t,�ݠ����,���:6p`���h����!��jJ�i��]&�ջx�C5C��k
��o�Y�z�8&�.�w|]���q�ND��=�^�; �si-S���F�,��ʓ�2�V����k���k�31�̂Oe�E�0����<+n3��zs���xx_n�L�����^r���)�]�aG{J����o+���y�R4��h_!��8���K�z�θ�cf�:���ܲ�p1�5�׫��p.l�W;�s������fh�
b��Ǳ<�b���3_$=NUڛ\߽1i칯_H�������2��5=��[F&�fϝ��D�}�}�N�n�&"���|���T�.���&��`�yW&�.�YT^@n��s���w��?a ��=�}�d �*���$Y~�( *��(d�ѿzC�Ḥ���8֊}�+�ͳp%��1��2Q�l�K}��ۢ�ޖi�H"J�]��CK7�K�s�w{�蹱J�Q��-e�$W#MNG�o�;|��c��������N8͚;����!3�(�X��m�]OjC�%p�eM�鷺ǻ1�Ǐq�]KX.�F�.]u���W���;�'�W�޾BU��i���}�J{�ڭ�.��
XI�[|s<��,j^Sx�:l�@te�Դ�ސkэT�4��b�&���("��gC`�|�����+��<��O*�x�T�3e<��s��6:(��t��w��捣V���z�<��J�:S��z��ڨ/��1��丷�k#k�o;/��ݪ��E��Z޶{U��/ @$O`�0J՝�it��eB�v�/)G�'n�.�+��\��r�ʇ6�E�ebR��AQ���O�����vr����ٛSˡ��t�J�8cݶ��d�pK�� �u�b�ۓ[����v��{�tX:ެC.Ǣ�p�|D]�j�Z:L�t£*�sv�訮��5��\;;�f%Љ�N�=:�t6;�ml�����۱:l;b����W;;ձo]�d���M
{94pXĐ�F!,�Fx��7���܅��u�"Ǝ��igK˞����zs�������mMNŽ�7^@���f7g�%�)���2�}Q ��"g'��*���y�弬wy�;��;��h�8ݜ;V�s�b�p�׀��1��J��I[�v �9��e�65���;�y[�`� |��iea ���AU��,$m��"�H���W�+��m%;C�_T���u�Y�w��,����K��*jU��X�K1�����A4$��o��i��6����w���x3M�����A��5�6w+���FtNևy���s���l���0�=�v��W�|<
��}%�b�w;}�]���c�SX�<���LS��0�Gnx�J`��Qx�6�ak��e*��<͛i�^ʅ�r*w�B��k�í�=�rJ����t^�Ɏ�o�0^�����CL�'�]z+�c{a�H�*fπpt�Wզ��;��c���EO@���Ų���~�S-�5���!�;]�.kE]J/���_9����]�^���L��F!��f2pRA�s]�z�-���s����,��[���	!mUUe-V�l�b(�,V$,"�D�EjA�Z�A�1J��l��ZX�%J""�R ((,cik*2ҤH����W>�>ͼ����?q��c��G;�����5Ğ��х�v�`X�ô-���c���V�"�>ݙ�Ȍ͹im�ɼp����+�zA���q�����DI���6j��T�W:�Ռpx��^9�NQj����*�ۥ�OV�^����\��8�*����Nv�ӱ�kz����r��\�3���gw惘��6�}3o�1��RG�<����u�g;�=/*u�8_{o��J2��T��A�=4�fJC��dy��yosf�1Waps�ܺ�6��]s�j���֦b>�%fL�Sx��O�u�@ȼ�w�W�<=�==�7��d)f��q熈��z�lon�Q�oq���j:V��ɪ]C�������r�6�����"�"����z���߼�ݰP��Ë�X
�r�\����L���p�!��s��V�Ck`��6���V�M�;�v�ӡHAW;��q���.��q۲���j�ɏ��
�w� ��a�n����)�U���5o7�MVjh��+��Z�ʵ�N"�V�sZ8ΐJ�]���UV��y&�w;7���3_y�t��o�64�!�==0��iaY��T�e6.V��k7�ӆ��c����V�2�瀾�nƼ��3Ҩa���6�GDӺ����I�&�ؖ��pu����[w��#���=�l��t��o��Bٶs����۲��FX��ò�]^X����"ЛW�<$E=gy�wY����*�=ȇ�&�nΧ��3��AUr#z�,5�9�o�g�y{�ם���� ��X���o٧��xj(���7�jޓHX(L6U�*ӫ���*��bf��h��υ�lP��Q&���,Qui�ۡ!�K���2���M�B�R���yޛu�6P���%���c�Ͳ����
�jP��r�gB�R�TTƜ�`�㎲�KM���h�i�Yl�`,�3�c0eLh2�q�Tc���y�2�wxh���Qc*�J�������٩ώ>C������e��R�b�}�K�f]����<��m�����b�=���͸�5���F�����PF����fY�Shtp�]{[��Vegƀa�����KM?���������v�^2���5n���l�8�mZ��Qb,xجSA4�d{k�t+X�9=۷E���Lz�ޣ�"��m�5��2�4���x�!�y.��W�q�	z��U�]k6�wi_V��s�:(: ���u�j�4@��?k�������"Z� �Z(�&��Qܔ�f&@�����YtZUM��.� UQ�������(�|�\1.	��fY+��f�[��U}Tj����%)�;d:a�-S��8�G�ǖF�L*+G,��
t˨4^�:�ݪ o�ф@���يM:@����3;N���-?l��o�P�ǻr������ծ"Vi����k	OkX(U����Y�~�J@�,s�U�zV��B�5��3v"B�yl�g2���@��r�i��v��u��od���[wm��ۓ�G�k�����a�������k�;��\��ʋ��nuľ���S�6U8��H��&^�u���p}�������j�dj�v�������|l�ND�N˿��X���2�������R���G�	�>'V�D���8�sWs��Ua�%�'����5�Yڀ0��9�9r�f��n[��c�S4���qc����*t�AJ/��ۊ�v���`z�yh�Py���}�r�T��)�4j�xH�$�
R�*k)�.yO���nސU�2�SW�6���/k�mf����a�t�;�3��"5d>�-7ħ�5�Jؓ�N��Qj��ww���'!G.�ּUbh!��	1����B����]Iv9�n�s�SnEsF�,�W��߬��ڗS�k�1J�µi�9]>Yj�m=}mV�Kv雦�b ���������F��:]tLR�]d������Wt��`�w|�d��s�ʂ�6���C[Cv�K �\m���йū��I����\�����41��ހ]-��B��m2���4����S�y� �]�ς;w'M'j���)���������yE]Ծ6-'bo"��%TZ�iin�$��>����ο;��iGt.�$2]�}[HnFx�.����}�=�?�ƱU�S6D8S8%v��eN�8%��e@2ȯ�|���ܶE����f��ht�w<fOfq仹���uZ�#�cp�G���y�=.�y;s
�r]�����[���-m\u3]a�wM� h�UǎȻ���yײdt��/�c�/v�f�����X�UF뽫�z��L^r'[���λ�S����ڱ*u��a�ф�  �͞�p�"��Ybr�.��;ՙV�����c����hk�<&v�^㼪|��Z��W����
��y�QV�D��װ��f�X�C�d>�q�S�X:�׺h'@u�:�Z�\�n㒗0�N[�;�[�0H#�|R �3�ލ�Վ�x�;Fv���:�-93(�����(�'���-˷��ٲ�K9EJ��;��o3(vlw�����k�%;�{�4�@x:q6��^���y�E�l�v���oj2�I�b��|�L�����9��V>�n�~�dZ[�4=s0ҹX��7X5�ۺљO���ݔ7(V
׃u�j����b�!�@��,��|�HsνNԝ�o�WW��]�m�pAvļï�n�b�ˆ�Y}c�[c��|��4��u��r;��x�j�[��z復�A"�aVg_����J��}����E!�M�j�2!������|��T^(���= �Weޣw]�i���@ڒ�l�Q�����\k�+Tۑ��/g\oV)�b/(���ej���0�VDD,��3��~���g��y0B ����f
֫5)�w� 7BT������$�a��R2��	+k(����.R�DWss;��9}\U��6��p�N{����qx��m��r;n��xzo��]�w��/yF�1]ז�)�!�\ZKq�@�My&}�R��
���Jlͮ·����[]��f�*�G_Mfڢ�:�7/�G�V7´�j�W]�����}.c{%�E���1����{�o�\�� ��O�}�{W[�|B�
@	O���e܎`��(����z�>�WY��dS囚*�e�i��9n���m��|���O\~�Gcs�x"�T�.�w�<�3<�D�Z����e�Y]������ODu�g�}��~8����`� ,� A��X,XE�A��X>(�P
����M��3Vy��g['��ҫ�Ĝ�˥SҞ��q>2�>���W�x7Z�?u1�B�,�Y�^[�ȝ]D��q��IQU8��Sx^;�6�1<��Ft��+	�q�F��s�Y���Nu�.*�)_W�t��c���������C�j+�9�����\��Q��
U��R�E1�>ͧ�U)�VI���Z����=�&{��y��Ht��S�;�L��cqO���4����;yٵq��sGTT��r�j*�'u��_��\�]�+[q�r��w4��fgFv��癒� �=߯ksW?����	d:b�}_P �{����+gt�+*����1��/zb�Doa�}��9�w"g��0���y׺y?+�3K���S�@y#�5���Q�k�tg\��5�<<��8q��o�|��j{;���NH���1�� �H�"����Ԏ�U6�uw����#��\H~5�bC�̧/4G�*�u�!�����Av��w�u�]�Kf@�''M�͊��̿���U�z�C���Y��!Ѵ�w�w�VGW�QW�
T\��ҰE�3����rf&C��}�X,B�;�8��_���ڜv���x�s��*d�r��!���?W�9zӮӏ2����3���ZҎy��[:㥸���FTK̐�{u��u\>���e���$��'%��s�z�N�ގini��
��agc�;���t�&�8�]W������#���c9	���
�w��m���F�e�v[�ML�^�.4ĺs�3Y7G(��z�J��V�{3�;�9p�H���dMa�[1[��f#G_"JQI;9�F�*����B��]��j�����jP�Hmw;�
_8�����S��B�\ݓ����as%N�][/�k��ݞ7�P�����e���C�2<s�Ӽ���J�����q�"����F�+�rcq��� �b�1�T���t]�ws�J��܄82+��]/u�'ڽah��N�t+��w�u9S�z�n���_ �웾���;������}6���!�aU����L�ѼV�����c=ˆ5M�6����'�^#mhV�=�hή�7\dn�t�ۛs�]{����E�k=�SmXC����FT�7OM8L���<xD�x9Ⱦ�q^��۞�:�T�s=�rA��z]��/�~4�X��" /mR

X1U�@�]�w�[��n�Ů����J��j���ؕo,ukGro{����5��+���-�WUI]p����-sq�x7|%xp�������~*]��{�t�c����uw�l�c|�o�[���􅲗�U]� UZ��=����sa�O�`m  ��=��}��Ojs����|E�T_>��͑�!衄+�8�ήU3�ˌE��X��h�]��R�Os4��2��g9��C�h�+c�g8x�1���O�2ʙ���j�P��]燼+���;�^����Y�%��ٱ2/-P���t��ٰ�-�b����6�O*�5�nojr��VC4�^C=y�د��R���P�����Ź��{Qe'/T.$t�aÇ����	�V������P��F"(�@Q �����/v�ݲ$���:��ۢ:����)
zhf��.�WI�-����4j�R�:姶�[ٝ0*�k�n��_$�w��^gs�-�����8ts�F�ށ`��k�fvV�����Nk��NN�q��{r��.LOlFs��οI��4b�c��Fwf԰`9is�C���7�b%\ÝK����^�mmx7� %��P��*�r&�{1�%jb�'v$5<+�ۦ6��2b��7ދ�dy|][��'����n3��I����?;\k�ћ����]�D���GH8on����7)�<��f���r�z���h����8k�������v>����O����{"�ta��w{�����a<���.�jy?^k��ߏ��{9��߰�"$RB,�@���<���J�Dh��S;�[;��MeM�jN�}�mt�F��%e��/���*7��%�R�(��Ηm%��*EE�%WT��P�d�h1Y�1oN췣>�4�-�w�l\��-��r}UU�<D�FV��:'g�u��ڵ��<\���DL{��&�T��t���T����]��<O,9��c>�P�'v���z�M<�L�ӥ��ў�K�{����Ssx�;��7���٥lN�g�xM�C�앂����
u��9��к�ҖE���p̱s�b�cޥ.^{�Y�m?~ʹgrީ�Έ���^M�}������]��^�����2S��y'rC�/��Z�$,�,�RC�u�����S��ַ׻�eM�cFk�S"�;��J�=C�8�X��(�$T����0�Q�
dE�b����maZ�UPUb
)"V��F�XDV�-�*
@��`�H��CD|~�@o�߬��x�S�[�H��N�!�n�J^u��贷3W��Ⲯ��62T�g޵̬̭��s�f��}4�Ƨ�ǫl>�8�N�j�C&qm4id�\r!wQ����8�=�#2�6�^�{�VFH��oE�K
��w�PN(;b�M��Hx{�=����O;|r�C:�2Tgt��0�#y�;
&#����j�t��W==2��}��W�h�U�/o)O$���{gR�W9b�u�`�4�y�Nt	՜�J��RU�rȫ��"�1��7UU_|�y�g
�C�[h��]��7��_vwwm����fz���q�Cz���锕����=$�W)���h&;�zTX�,�y~�Z���g�E�ػT�'/�ó��]����Z*j�����9b������
���~<辰(*�B����HEU[��U �AU@�"
(�Ԗ��"* n�AE�}>~�ym���Ϝ[�6����zffzv����˙�U�Ҙ{�5"�
�\�AX���s�m1���}ܳ�*���#˥�$hk�'d��
�*��AD)����*�������C���?֪*��Nd�E�;��vE}�<EA\7�<1оA\�A^:0m@Dc� "
�+8����)�5�]#�%M��c+J��
�do���t�TU�.$Տ�t�VEA]��A]��jDA=���8�9]y^VƠ��	��AZZ"�������c:�+�H���F��L��**�{{+�q�'�b��L������ � ���@  nO���A��TR�M�1�X��T�$���(U��'Z�(����PҔS��35�����D��UJ�����U)�4�*�(���TD�"���)AB!!-�֊��RR)(���HHD��[[%���k�   �P�kjֆR�D���$
���w����     = t�Al P\1Ӡ�@(�i�[h���s�m�e�i��ws�j����Wr�kd�v��-�{������;ܽ��8�z]��G;����^����֛x��E��Q4{���{{�{5��r\x+����ڼ�PRu�{�5����ĸ�P����������S���ޜ9v�uJ/Z�рw`%�R��K��{o)@UM�M���J���Z�d(���w�ǀ�*W`׏.�IK���q�mv�AH��DI@��ڹʩ/Z
]モ�g��g���P���օ�z��P�:z��{�7�����˽��x�JJ��y��
B�;�V�Uzh�5��(��R���Ut5
qP�Ekw-�)@R�t�U�D���<��%�of{�
�A03JB���w��eSYxΩOL�y`�j�*��9�U��Q����jT�6�N��hiJJW9ν��J	�w�V�mw��u�Ow��i%[���ʄ�:�N�9�wT��P�;�V�SA���<&l�{�%U)^��
QR�9�6�{eNu��C��{�������z^�@�M�S� �� t�8��J�`����3�0���*��ԙ[[@ R�9��A^뼯4*�\v��$z��ljPV��V�h�����qq\]n�8=T]۬��B����UU7Pk%ҥ��Q))%�zKEݜ4F�k���Ef�9p誤�m��֦К�����l��i�c��Ҥ���{^�M����mU�`F�z��#�0TR�5\�����ײ�(^곤.���˂"E ��[�rt1D7K�	�.�n�¤w�ު�L��r�PW�7�R�0XP��R��޸Gzoxk����Ըt ��^z���Me,�gq;��C�nNu*"�n�8z�]�ޏRQC�x�^ؕ#����� )'���
T�!"��O T�A1R�   �F�U@�� Q��  Ѡ "���T � S�MRU    �HJ���&��j=O���×�?��S�W�?�>��!�Fy���v��8�=��w7��{��HI$	'�'o��$��D���I I?�BI I,C��II���I$	&  �u!$�$��/��������X�N���6o��zM_�ߖ�A�.�FK=hY�k�5<��V�Bu��^��d��;[�^K�B�t���#w���1�+,H�=3a�!�xʦ-ю��L��EKٔ`�wۄ�P{:q��+]Sd��#K�~�F��Y%��w&�8�W7u�����j5z��2�ISEmѻnd��Xk*�tnEVb���"���ۨ��U�Y[z�֯�CJܒ����	W���o��M9�@������Lʖ@BӃl���[�밖�!_y��1��h�&C���)�H��Ah*�I�*�� ��kM��Ӳ��=6j�� CZ�D��S��CL�÷v3��ʲ�"�͑�i��`p�uY�jy4U�u�&�L��6�i����,�Vf`�V�F��n��̊"�ه/�F���ҩ��$}�N6�5�I�z���\.HS�0��)���R��Fr�fS�Gw�,8h�h������n�kU�<z�"��ݜ�0Sw��ph[[5ܥ-�^E�,1YH,�o�������r�]\S}X��
� �#%J(����R,EI �A�X,��,F,�O$��*�0c��i�ֶ����wg�1WʗV@Ҡ(�DA�1 *�T�,��r��ܩGjЄ�3V�[��
T���&7=�~�:�PZ2�+����(QӞ��Hi��(�*(咦��6ʢ$P�J��J��a���������4�S�}�ɞ
6̂z�A��7yN����p:�pf�f���o։8Q����6�[��Ь]qm�{<�n�s}�m�da�DB>,;5U=R�\̫��xb���fR,ԣ;c�.L�b��70�2�F��X���F�N��b®��g/C���+�u�Nf`͓!9�W����C\��l��L5�{;�k��u���z�W�7��89�l��N�0��aQ����7����{r�q�x�`��B'�~9����'���1U���pW�Cm��c����� H��?|�eQ�d/�3�f�K�Q����t!n�@����3F9�Fa?11n����&���(mK^_�����C���ʁ��T���Z&ǋܽ���O�C�y6��]��G6M�s�Ͻ��sc���:�d=�d��bA�ER,4�����dQd'N�o�4�aR{B�AEX��H�'���i�I���q����@TaԬ�Vj��P�TDQP�i��(M�dXH� "�������
�@XaDM0���� �������p�T�R�R��O$�ҁ�F�C �[ke�(Yb�w�mIBVǡ#z�x2�ՓTN5��x��������Ed��}�.,ǡ։fM�Y��0�J���߽$�$�7"��k-��h<))�2��s1�'r��n�`�	g�rv�C�_0B�;�^eZ�ʫ.Ibc�	B��#̤�;��;{�����,��v��6��{q�O^b�y������g*�j�p�޿��"d���fF,�'�5�)��&�*[�`�IdÚm�k�Vn=9�6-	�aV��9�"�ED�/qM�Ed�� i,�����VY���A�}T��#�Q�=Ӓ4�����2@ �7�U�7R�a,�b��/�n��۞F�h!���f�)�K�;	6��x���e���e�Ҍ̶٬�]�1iU�V���x����r&k&�{�7&I[6�8��P�q��lI4��R��̸5D�skv��3|ez�;%��Mf�`ٱ26{ͣ��6~�=J��>"/p9t����L7�r�%p��L���i]Y�r!���T/ �8N�w1���ٱR�aZ��NE���8��X��|��,̸"�q`[���F<n�5�4�!�Ƿ��ݚT��!�-�~j�i�����A9~�#��˹�yՈ�z��n=��{�ﻆc��{�����<��6�QAAb�TH����"R"�ۇ\m�"��t��%X�7ksM˦��:��de9�7X�D@��L˩t(Aq���!U"�A�)�QDz�d�d��u��ˡ���Z��7d>�~�Y4�)�B緣.�Y��ɧ\�v�[�N��Q�v�-q�yU���c�lZ�)��LԳO�T@R�g�t?|�e,�u����"��bB�9f��xʼI<��g�Yz���&p�y�p����knL��_��+W��0������y���p������ɺ��6��z=�c�0<���u�[�
�����Co-챥���h�"�l�]���������d�6ۅ�w2Й�|T�����������\���R�1��+��
I�<[m���Y�nyiܸ#JA��P�����}���O%T:���2`m�޻�w��UQ2��U�Elò��)8�2�p�꺍�^'	'-T�P��M��[cܤ�rT�Ҟ�ҽ̲@0���=��b�f毶]qh��չ�?MY#��/�륨���o��^����H����@ًB�����h��w���ʳk+<N�r�,-����f
�	�R/�m큻�w2�5�ǧp�V�6g��g0��Y��������z���,~~�S��T����u��]7�^�^�䭵.���x�.�h�r2���[ö�4e�-�+]�������#e[Ȭ�_+&m�A�S�����RVL%��+wv��&co/gQ���%]�i ��1���^l:��i��W(GWH�=t��0�`w�Q�5ۈN�wT�W��
�I�����J �
�V�W̱wL�Z�
�`)(��e���J$��
���QD�UY\�X*�1�gP�Xsx��n���!�I�4K!�W,��`�ɦ<jo�P��N�n���I��g����w���<�򒳨��E�{`u(+6�A:Ճ+H,$:��;�k~�e��z'n���6J �{C�$[���Px���M"���T��R�±r��C:d��"*��4����d��*KB�9t�(��
�X,���J1wiX)���>f�Qb�ԨlT1��`����D��5T�{�q^���`�]$ֻ�x�� ��,8����i��^�ڊ��3�}�Q�rl���	Lz���y��l[�54�{{h�)+X$�dt����;�o��!�x�VM�) �w���skC�d^�_Hmr!��q��������j����HK�1�:~ر�qm�5&qX\��U"}i9�Z��w���=֜g{C��HR>�����ȣ��3�G�v=m��|�����SY--!RR���Wʖ.��{���E �-�*�K�6^e>̑ZqCxߑ$�w��j��n8ݗg�O�B482����#$�o���ײ���h�T�M��,��C�0���>�z�&Ke�|����y�1���-&���4(�f_��oޫ�~~��{͠���X8��v�2�6��m:�ǡ�wzQ�JE-��jI8�Ab�����CK&.��Bb�b` ���w����[D�g[��ц���0�3^]��d"��(�҄�[0�f^c1I��v��2=�u�Y�m	@�i�촥*�,�BR&��܈�v3{L�m��*�KޭX�1�t2�qdwn������Y�nT�ADSIb)���ǡx�����E	~��=U�m(�t0+/V�ͤ���eO`:`�ɗVT�WF���KT_��[W!������OTˊ��X�Z�97=��4o޶2ݫ��tԇܗ�[X�ʹ��ɔ1���P�����������|�w�P�P�@�J�J[�ث��L$M�ٮY���I�t�*�p��#MԻ�˫$8⭕��fM�2���v�+ �d�s�Y�Þ��:��L���c���z]K֩��K���:#���vb�v��%j*+K��7NL�O�ۨ��T���sGT�j�;�``��" ���e��Db*�4�EU�DEDb��(�"�A�D���!R ,�N�����:�y"��!��i�n=@�i�<�l��J�Z����S�s�˲Kݔi�p��Wf�6��X�9��z�ay�7|��O�@Q@�Q�Ȣ�d"M�(��c"�TX�F,���gki)D׆�% �BI��4^�r�`���	�1���%x�x<W�e�s"��5���,�dH�ı���Eل��~��܁;��M��u��Ul��x��o�5Z,�lD.�Zj��7�QZ�t�u6 �������^J�W57��;�n4d����^e�|�0�5�$�)��Yx<�������Z=&	�0�Ka#3�A�5��Ϯw3!�DQ���<�w��o�X��2�"n�V���YV�^U����3�w�I;��Q�J`{.ܛP�$-9��i�5��tC@[�gt�N��%�J��uO��eDv���n���*����[0x�EC3qk(P��TF�8������ǐ�6�6��ͥ�Ó[ŧ�U�ͤƴ'O!��]A/Z�����&�����~����
�	���:1�S�Jy=�"*�J�a�O�;�W�73ٸ��(���1���[�%��Hy�����g�I�0�	%"�e�ᴊ��.Jw�
�	�\�w�R��L9 �6�(��jY=`?3�<p�~��L��厄E����f)D^^6�b1c�G �c4e��^ٛ��D�����1�I��2n;{�(�eJ��)�*��yk)�M�*S7^b��CV�����ɭ=B"T��-��#f#�ٕ�/SI�����(r��Yc�|r�Rw,��J��p!(>��/յ��tK~�j�j�����(l��V�	 {wN̟L_L`�9�X�X�F`�-�߮߱�h�4�-6�;d�M���B�$a�I��,zwE
�����۩L"�"�5Ǚ�1�ܭ`;Wj�VI�5�V��W3%jb#���N�qe헏X7�OIy�dݬ �YR���<=��~�e��-��Io���s�7݂���|����1;K��Ү��e�LSt��%���V��
zP�w2��Y������Ի�� .�#T4�(�F�u�� ����K�5�EL�/���q��$^Tc\��hJ���.%��J��Mخ9�"߭~˲������Ff�enTs.za�E��:�,\���/��������7!�7�蠚�y�D[}�� ��3A�Yx�ٞ��>Bb�kg~K��rzz���$���H����PL��^n5b�̓����	�����<c�6c��E��i��i���?�!q����T��ʋa񒇌ۤ	OnCtM,���5i�gR�F�=�50���1�a��`T�
QR��eE+4�&�fB7U^;l�����&��Y�VK�z�ס�����Ȳl��M[{l�C۷��l��Vס2G�����N�d�V<-�X����0I�g�2D��
�t��Ѝ[.W�>�	H�c_'Sr�d��M`��͒�ܶ*	6�nޔΔs��p��Ջ'�8L)�f�:|$���
�.)��6�[E[>��2�^�h��a��p�u{M(���Ӏ�"�fB��`ih����aQ�*7+]�])�l�2�Gj�YMX����1�p�M6�M�+^xbymM�� �n��v�c�	ǂZ%���Bb����x���/|z/�A�V�R��f`�hKV"^T�9l������K��pb9��0�A�c�n����wJL&(�{(̙��V�LhaMn&H�Tѓt�}Q�2X�i�52� ����#35jHdl���N�%���vk����S�+op\!�6�5
���vdO��ަ��[��'�e�&}�=�r��e�u�	����b�	Vb'ٙr.��;���\U+'��xޞ��8�-M�T8^{���,x���f���n>�0����*����O�;��s�_�&�[�$���ra��;xWP����JW�̡v�n����ג���l~=�.��(����'���=�ڸ�0��J<�s�����
���<�������q�:{
�*�(a��x�`��0+���QSn��o�u���]f>��j��K��ƸT9�d�V�Z�����L����;��^��^Ն�t�9H����~I{Oi>���U�>Z�����q�Y�ͧO�y���u����,{�%�u��	;�k'pV�v*9t�*i��m����:ڒ��moW"���s\�,^�M*�U�\fY�6�P3sv:���ٝ*ۅS�ݫ�_z<s�m��lo�.r��ݮ�c��z�T�����x���s�8�8����R�L�j���!^�:o���X��>��^����ƑS���\��m���+�7�H�g/��ptn��j]=�ylgp|���e�x�WLo�f3h��0m����h`^C(����!)��=���Ј�ŝX�q��*2<�pN�F�M���en�]�G���3����uX�]�1�(M÷Չ �_BP̼�k�c}�uϠ��I�h����p.)�y���}}a�{���f�E����#,pO^s.]����K)�=*�|E�9�B�g�cz�� �3��5�}x�ίJ�c�`�ôR���qG��4L[��%S����uuk"R�iou	�o.�˽QW0�^͝���\z�ۓ�w��Ya����w�V���4�C˭?��,�Mr���O��'.a{�9��V�a�@sk6�X�ъ<���� ��]զ��[Fw{�WuN�a|H/�������t*ŗ����W�`B��҆<�}�@��o/IF����Gn�7�3*��yN�Y\�����d�Ǧ7��J�ۺ�47�Y���h�q��v��gp�{�>���!"o�Vf�����l���6�ג�y�q)�˥@����L�a~{�i�{��b,�9�Z,<�<L�8�������M}��<SˣV���ׯ��=�ݶ�H>X�Z�N�:m;p�wH�E�c������y=Me��Uս[��6�ͣ����/5�~�W:�2p��j�
�ntۇ}i�w`��9��r��2��:���W}'<��P����t�jMb�c��X�}�q���b:]u�6����"[�y��Õ���n�+�Ҧ���H��EX2�)Ԏ�*����Jû�*{RX�ܓ������r��>�>�mط��s� ��l/eH��1�۱�X/9������f�[�՟lS�"q�_zyʆT��ǵ�2�!n��y�w9	�  ��$e�N�ޯy>�a��i��H\q+&d/�g/�� w7]�+هQ�yNG�ٖ�K���k�����o�ܸk|����y�N����TF��k��;9!��`�%�$bu������;3c��2Ǒ���侪u���qi�_����d�2��x+�C��q�]�n�Z䡧
huΫޣ[4���w�r� &�(��s6�HT7�־�;s]�����ۊ<��c)�3oZ�}���� dæ����}{���mܼ#�!�F��ݴ�Fr�����%��vqWI�+�rtY�wA��AV�p4���Ϧ��ׁw�]� �yzI|ph�-�O�ƇGGf��9��r�F �6�
Y�i��<��rT0��#��j�mf7�`�mS��{��>�l������mLe9� ƄnR7sr��d�x��LR]��I6ङ��RK�w`E2Y��+P�t/�fu$C��&ݪ+�q*=V���z��Q*���a�x:(ؗ{6�7�,�\��P�@�M�h0b{�y�q��pnK��$��Z�6�oR��,ս��bˢga����5��
C9>�70�iY�r���k^�1s���d�^I��!Ye�v5LV���4�8/�ݍ�\�]��D8jVP���-,wFDM��ۭ��d2��:#	�ځ][�fR�zb���W�E���x�D�MA.{�=���:�qot���|ʵ:w��t�|��g��߻$p׸���'h�6�98�T���i��N.�l��K����/�	�j�+�\�e�웯l��7�!�wB1t�Ӊ>�=���`�o)+�^��������3��d�8�E�9�3�	
y>�lV{�f,���|}�i6? |{fG3z�!����r�1���G�s;�{��߶hr���i\��ٚ��3���͙�ۘ���o��e{q�>�B�D��3v�ޭ4�GD���qS4��;e�����ٔ�G�S]��Iy�훜gila�o����&g!��U��P��^{4�O��_��i�~�	~:�C�yq��]���,���E��� �=�mb�Y�/M�)�R�SK�t4�i�PCN�K',�/����Q�MY�C�4��ڳ�6�ʌ�`A-�XN�{���]O����t6Fb�
����v]������W�+�Pޅ 4!8Fr�Ggj��G�Pw���j��^ɶS�i��niQ#s�k�'n���}�V;׋)Ue�oc]ԥd���ٽ��V'�f��2q�η/���*����6����ݷ�Ϙ�N�Q�l�r�����w>죛�MRf��,�}�p[�}��Y*�r�Q���8{0�:�B�
P�TҗػOqaq�K�S�>�/z�tvx���=X�#��wE/�{�bY��e��1SI����:'cc��f��A�[��*W� �6YQj`�s^�˾�������j�m���q��3A쌌q6I�m٬�(�gv�[}���>7�>�C��I���ᐪ�O��O�]s�۹� 5���u�兛ϔ2�n�½�}3�6f/)������K��Yf�� ��v�Ëb��.v^����53i��k��r[�(MJ(�ź3p��b{�w�M�S��_A����>I[[YǴ��oM��̐��,�N�{�ئ��4.R���2�*�j�qpSWQ�={vs\�f�(�ƴH^z��܊�n�{��MM}rX�:��vo�kyN���Ǟ�&]�:���hw�.�:���B��s��k8�|�]�C�� �Rx�z��9���R�ts�jk&��ȗ\���i��5�\<�����:YU�փbCz�0�E!t��%�o[�2[�ϟh���xg�H0ݎDq-��x�ʹ����uu�jq�F��9X_�ǟ��}�Ho}���B�h����yd+�$����FX�l�/�j���NivB���:��q�X9�;��<�;P��/aI��m�7ul�FB��J����IK����Cqk�3F1r�u�e�3M��3R�g���z��
�3�u��.���\�9:il��wv���͑7מ�޻{<5�{�Ӹ��� {��:=��cc8�LSe-�t�U�����"s]�
�L��J��Gx�j�f��"������vzzkm�yv1T�3����I}��p���hp9�����ga�:{K{����?bK��14��{K~$<�Ε�rM���(���I¦"��;
�u*i#ʌ�ަA=�|'��
;�@��B�Nr�֏1q���F��s-�]����:�/Yw���A�����`g����0�xX���������+���#��+]�����P|�k�P��3��ثc���3���c�p�Xl10�,���>�슸t���3�ϑ��m�c�� w�Q���\��Jݮ)����� ��Ig�wj�_;�6_3Ʈ�X�������o�J�S�Yt�CZ8-dMX��x���3V�5+jl���sjȥ�EK���$K�Ov�*�Ȼ}�#��D��z�u��fg=���Ԓ��X^,��s��1�z��i����W�˭So8D#+2�m��n�n�VS����v=��,����Y�S��y]��V���I]�,J�OLr]d~�f�#O2��K3�iv9i������^�Y�\��vD��7�J׻˻�i��o'���<���=o���n���6Yf3��N�n��fK�0K��&%�6V��h��--�ʻ���HE�*�gA�+���3O���m'%"w1�ӪbƦ��٬��fJ�w�u(�Ay���E��]p�<}��C}}S�l�ng�AH�=�e��;{$��
f���e�
wg^u��n��#�t�*m�Ȑ�S�`	&2�9���e���è��	1��5�S<3`�˘}'�2�lyv���1,o�s��3�/8ΩY���[2M�avk��G&��[�a`����x�y�x�	�����
��}��;���j����h�G]�轳��ӹFA���qrwt{v����s���;�=Yqk�tNT�Z�I}�o��|ND�������kx�-E����h�9l˜�>w�{GX��7�L �	5P���Mi��;�<) ����'��uî���x�VƴD���a����Ɩ������pR�eY�3Py6��8��Xp�[�}f��6m�Ze]U�IF^E��Z�$۪Őu�y`J�Z��f��u�n0Y��yU����y0���#U��1�j�V�v�19�j�;����zX��t콯h�|���l�YjYl���Y�Ѿ!-@U�V�ɻ=u<7G�z�zV�æ5s0CX���eZ��8jM�u!��b��S\�L1�#ܗ�T-��!<gq�7����������Gh��9|�\���4K�X���y��E�Wޖ�Fww�Ҷw3c��RVÊye�X}yOY�,�ݖsh��GM��X:�)$� ��Ê_tG��8�+O�S&9=��]Z
��
���;�%Nu�k}�/m]d���*ݒ�r�'�VT�'^R�b�=����=H��;�M���ױ
������]��Bf��}����'׸�<��qu�nGv}w�ͷ���F��(��^���m�x����{z�tY�\H��g�珢�>�L�ny���範gZ\!��O���Z�;{y�>���Z��T���V{�y�&�nd뇼������y�~kr�Ax�e�"��
�$NY�
$���}�_t����gw+����c;��u�;���S
��eC������޷��^N��ך�{��#���k����t�s�8"�����9���{�����sv^	Kn����m9)32��\]&Y˹����nS)Ekd��F�wS��8�<�{y&�����mȈ���)�{�p@��������U�^��ͽ��k�����xk[j�)�΋�����Q�zw*562QʩT�L����;�	��$�N�>��cf�{�y	}���R�/����!�._E[w}�zy�W{m���R��i���;n�]��y�aVA��?2|�_m��Y��G�P�ٺk���%]�{�tU�ܑ�=ǫ��fU��yV���QY�9���%�db��t#O5��5��wD<�0�f��ݬ��uӽ�&z�#�q�f��l5��������S����X��T���N�a[h�j�N��R�<�(�8;�j
�a}�|vE��,E�I���!Jީ�^躹�hnv̫����>��r';s,'�f�k����]sy�Ǚт�Y���/�Ei�R��5%4����7D��c�,�GU �1R��V,�!��p�Kp'���b�:g���i�9�]L�Y���՞>.ueٗj� MK3h���6�Ec��,�^f>��x�������({W���3|� ;jk��P�t�������p�
��j���Ňg��V�Y�@��,�CV������'ϕ����d��^������K������"��&�x�������Ī>�]Jb�����z,��4�lt��]�]ݝ��e���x��Z- ��{�鉙�ݹ7�Salw�G]`�� ��cĝAnOt͚U��/G�Ln-$��e�f�KՏPܓ�q$��(���w��Dw��/R�ྴ{_,O�J�Ըզ��2�<���)���C�٬ݣ:�U����嘶su����NM���ạ��U&&�S��앲!	k8�L�k�|w�w91߷���%�=��"��H)!mB�e�nB5���KБ��f�f���U���OT6�"�^���N�:��q��^�Վk��b��W6S��"�Ys��On{	�4�q]��/%IySZ�8��{�P�\ɕ�2��
�D��䩽�TfM������i���b��ዒ�{�̞��O>�����W�B��X�*ƷSB��5C�JD���,ǣv�Y�-Y��r8]<(�=l����[��w]��Q�;��SO�k/b�d��q��U�O���Ԓ��e-����fv@�������@G�h���S�n	|���ӹa�sqم@��g�j� �8��*�/�}?$���+��+����EDc���{{�6�U���B�KЦ	m�k3׵�Y�n1����ì��cK����.��mH�ܦZ�k|���a�K+��)���ݝ3���n���ɜ��%K}#��E�֞w���;=2��&σG	��;�fZ��0���� QӖQ�V�fi�j颪�d�`�h�[S
�>|�Ŵ\�#�h%�aD�|�vo�3zZ���@}�pec`lb���}�yp��ÄwS���k�Eӎy`�.�{N�=cl���uD���ʋf��5w�d1%�d7)���o��k%��'�q�ص�H<	�ʩ��}L-¥�_]f�;���',$^����R���
���>7�k�%����sX5�`Hۉfm	ԛϊ�#r��&�9��3���N��pIu��.

��Obӑ!�j�s:�M/=ۊ�dI�K�����j����n��?�U�{��W�?�I$�����I� �?�$��?��	 �B )M� ��	!R��C�$��$Tl��,�sTM��� I���HKl�O!$�d�@h��i��1�Y m��!� m�I1��r��`N2LHT��Q$�Ba ���HJ���PHT$HY��200@6���"��l��Ra,�d�a��i�T�����āĒm� �i&�C�B�i60$R��P��I$�v�d�Ld��*�"���H��m(
�I*L� m���C�6q�jÉ+8� 6��I�j�{�d�� �J���I���Xf7�u�I$6�)�3�P���uNv���lY���BM�u�����3�V(q�ܤ�|�C|�7�H�:�%�hg��L�������0&u�ef5���"�e] o�u��q�HTi�Shi�CL	��2���z��咠�:�oSBi����++���w޳>��+���	&5�2@�I�4�l�HM& k��^Y!�q��9�F��ZI&9l1�k��^}B�r˜û�� 4߮0�>>�fj����v�0'��]��y35�_kGܦv�]�u4ͳ�u�q�z��:=�5�:�	��7�H7ｿ�x�AՒM��C�)�	ï����;�$wVe�.�H��+�Oϵ� @�t���8�9����14�s��&�S��˙sL9o,�l�;t��ԁ�{���MCv�P�yc�Z����A��uI���S�*i	ֹn5 o�O�p�Z�� �o}�)�7�BN�of�`c���ϟ������� q�Ӝ��9<��pyc־�館f�/����s^�'y�:�I3���`��ϝ=�����n\u�5��P�}�������$=�yӥ���9N'N^s��S�ѥݲ@ǛK$���j�{{���dz����Bo�u����H�8��q�2�{���'-�:nI	������֢o��w�B]��/�b�p����Jp�UUr�º�^׽���kU^��nB0q�;y�fo\�2��I�~��0��醽�$=����Ih�j}6X-�=�1�ԑ��!;�o몛 �]��y܄�9����U���O�9��]/}�og����P��5!�o}��!�۵�{w��o+�8�כu�]�UH�X�P�����i��xF�؎��I�-�-b�UZ�)������Aƶ�ܟg}��!���<�d'_v�l���g;��FD��39�׎( ��=������u����1��ջdsCN�<o�l)�	�zjhqɟ����zKYq�WX�i��+gU��C�3��c��uW�����{������:��!�kx�p�k;���e+�f���� y$��2p^3S�?�̢�K�{��&�o��-ov 4W��۞%����g*4�l�NXE���tY��z�Wn+;��� ��eI���n��{%���J�u��Nl�� R7CC|l�,��h�C���$W�_&َ�ϼ=b���Vʭ���V����g�d,�Yn鞩�$c)v�\&���:�Ʀ��妶�"��H��":��ۼW��<y����d�;�J��6C�i����i�kr��O��or|����;1Ճ�r���ˈ�kg4�J�B%�(�[�I���wp����G�j0��̈́����v��wW��n �Vɒ:dnl:t�(���R�w}�D���v�\4d�W���X|0�B����&�ݽ�t����C�Ž�@�H{�>
���g������e�!��hâ��$����Gl]R���̀\���x��Նڤk�=�B'H����v�p&V��Ϝ�2�"&��Q�պL�w����eH��A�|ׅP�I�Gr�t�.�ݿ?��qdg��1�tQFZPY۠��+M_en�E�g��A�	�}�y)��?�
�˶�͝�|�r���+�b�ϊv��rx�I���Y-_[�ZB{{ԋ��.�h<���+�?8V��y~����ȑ�ug4�]�F9�x�4K�,�k�\���ҟ*�uL8�>X]�xӥB
bdM�T���#�u�i�f�h  Y�c�nE�{��>>� �c=��ݎG��+c��7����v�eYnJsI�ē�����$n�<6G=�H�;s��>�S����t�z�־�b�=�����CW�0�;`����|�ܩ�
4j�~9���B��g��|B���G_�Q�鐃b^�x�:���T�m��F-ˇd4
>�\XT�'N��Q��+��&���D�1μ�ʤ�!�|��ś��A���3.ٳs�o��#Z�P���Aы�Q����"���8���đ�.C�=�]np��*QL��M�Y%�X���}�n����&�B8�D��d?D5ڞg���y�l�`]��$�(hT�����Ip*��/�JM��_��/|���76�L8`f�я��wu�DR�U��߼�����"f����f�)<}c������� zd� ���k&y��ta+'cs���=$x����I�NxܱQ���4�T��&�~+\@�XB�R�mz+�~Q�Dcu�&"���N��#;w��{ۆ�2k٢��������Ȗ�a�F��"T�w�n�W)�1SH�+:�ڗ2�k�t�?S�.E���rB1�xc*;"�I�b%[�ۥ�f`23�٧�Q����L���T ��!˳�#tӧŷ������EA��~д���,,	�	k�1����>^�3\�W)��7?؄�@���?�,��V~�x�?Y�<��A�TpaҶ@���u�(w{����w�	2��P�Nu�WK(u�J���mJ�fNf��|1��)b9�X���W�N��ΓA֭X��M"���9���PR�Zp��"��{8*���7�klq�vG��[�]�j�4��=xWL�\�O'D��P@��]����3rNm�]b`��t��N}Əm1�n������׋�A���ښ�]%gX�c�6-�����F�Sdt�ڜL�m�h�kH~V��n�� �n���D>�.�+ZzӼ��P�ga����L�z���Y#����j�y.^_n|$A��m�����mwy�6j琳pа���^R���Q��jh����×�];�ث�OS�yKܗԨW
f��e�t(�^VWD6zͫ%Ni|R��m���8����Oy޷TqNg�����3���u�,���ēv���4{%Ne����=���cm������oǲf��
�d��$�`+R��Auͦ�L-������&�}�i>&�������otn�j�*��+v��N�/�1�_o��}�y�Rl�!r�0b>���ٹ��}�3I³BXw*�W�4���Ϧ)v�]+c�:�m;�Nfaa�F���!�K3\���V�צ9�.�T�r�����S��=�6��x�s��l榴�N{ϳ�_}�������O߫�]��ߵ�����ߞ�� �J�y�+֙�|�Ivw��2{���+
�1��J�:�j�k�R�n���u{�:W���yyϷ�s?��$�2H�B}��Є�$$�	*�aid�a<�y��q!'HO2N2ͧ�$>B` �!��&2�N�0	�IP��Xc&�Hu�1!"�~��M*I�x��{�>�fa��{\�����V"�Ԫ��H��UQTEU���Qc�b*�X��6�QQ��F���41ET��(�Q�1U`��j �b���A""��DU�*��a�`�����cE�Eb�4Q�b�(��(���*�j(��dE�\b+V+1V,E��1UD`�~��F:j�uK�(��J�*"#QYuL�E�QU�$Z�
�QDb(�舘"(�icAQ��A��U�*�v˖��UU��#X�*�A�TV*��Z�DE+("�Uv��T~�(}KF*+1��*�c�T�Q?Yc�(9�d�D;Kw쬈"��"*�U! DA������PQ#��2�"(��iQQ��˯}���o7�Ժ~ﻭ�C1EG�*�TEyJ�ELJ�A]o�]bj�5?5b�(0UfZK�^�V(��fZ
��'.!�j(�*(�[�ߝiTM4DEQDEIl,|��(�/�h~�UUQ�#��zʤEH�-����6M�DUưTP�UV(�A1��Q��!��"DT|ܿ���*,TU׷�J����;eUb�6�fE��U\.�q�iY����b��^v5���Ѝ��.�nʙ�w"�� TA�aG֢�q�
�X�Q3��X�"""��5�b������i
*���R�+���E���QG�be���AF9옌cw3�dDWI�
&��iQc9eY?Y*Ĉ9C�1b��!�`�����YU�Y�Vnͦ,U|Z�H��d��2U]6uZ�Y�b�H�yLҲ>���[�����V�,q+��UV/�LQX���`�ĩF��F�Z����3G-Q���բ���O���F:�~tcX�E�R���ޟws@�>�8ӍU����-L���v�,�`����VUf��Q��:�O���բ�ĭ����2��BB� ��/s~R�0Q:
�~U�3����{����cuk���X3=f)��J�1�.]aQX�|�ՔA��\���D�V" ��-�3J��a$*#-ӊ	�~������\��&�r����&�ܕT�BbZ?x�~/��jS��2rb��,�DG�"V���U5�o\l�����Fj���CN���?kX�T�OԪ������?rhq}O������Q�Tb�֪�/)M*R,Z�6n���m���bU#���/�W�Y�AA/��P�h�h�]�8§�Z$D�7�f0�hc쪫3�a����|�2�A"�[�a�-�:�*&R�T��X�Y��~�_�F&������UU"�nګĔr����\�.�r� ���4�e-���Y��i����uӚ��7j���Zɑ��SX%���({��'�X=��j�LV�2_޸�\y�X����0�/����7h�V��U���QQ������5La��Juӂ��,r�ϳ ��>W�|؜��9����ה8�������$�$~E��=گD��q��?e�_[>��>����S���A������Lg�3
�[֗���b��}u"��`�ک{���e5q{�f�ߩ�4��f�=��n�'�]��y�s��kf�V��� ,~+�)E9�i�� �]�X���@e�E�@��2��9��0-�.@hd��j�-+��}q�u-���X)�ׯsm)�%�5t��N��M�����W^�P�u5۟P��Oj��ŘZ�fSf9��Kmˈ�a��X��K�ɭ*��G(�V&�����ӱX�M60���ί�2Uy�"@�A�-r�D�����M�<eA�3��Wc��-N9�yo�{^��T� �� 0R��j�	�D~D(�(*t	��!��TEQ��M3����m}�{[3�b�v������<Ch��8����jTU��o��4s�H�V��R��I�S�QQ=��b_i�߲����n~>>ɚO�S ���m۴��DE�y���.4�y�r��R���W��[Aa��*����V-B���.8���&�����i��.�"�1���|�~�:��D� ������}t8v��3Z�|�b<N�s��2Z�f}~M�ڛ�����`�)E�����M
V(����F�Ņ�0Ļps�\j.����~M��Ue�rܰmMZ��+e�lf`������{�w/�<ӛs|�<J)�=�Sk��a��5T��oCi�«��52;󁈵/�Z�1��g�/��Pv2K�=�~��8��}�3l��vw��pWv�J��2}�b�i��YQ����R�t:}����A��:��{��<���w0k�
C����i~��A2�������7;�؛C��/﵊7]swp�1�fn�fh�����}
Ӳ2�bf������Q�2���_�]��9����Ѻ*��7�:3jgp���	���LX�}g�o�|�������[�洶R�O�f;B���/ﮐ�ن�׳�����`ļ�z|���?4���PL�f[d�0Ke�\K+�ߵ�$�iݨ1X��)�����(�QE)*_5g�G�TO&}N.�5��&@����Be	�Ւ$�_M�9��JB���W~�����A�@ ��'�����Q�MT�,m�J+ޚ1�������y���<��Q��3N��ol\r�V_f=�ɩ�(ai>qq0-�
r�ZK���;�yƢ *���,D*���"��X��QE� � �#U@S��)�)��nT�6P%}jJ�Te�Gȣi�n�d�}����̺c�T.�#�f��O�d��Ғ>�QGR������(?�"���dĬZ�ۼ�fZ19��v�<K���^���fD���D?"%%�S0PQe�^ˬ��!�<������L�����w=[�CDm�B�Jќ���u�Wî�Z�$�/��g M��γ��]�[q�C��Ac���+'M;A��m�ח%-���x�-`|�����f���#j�ei.>�	�Y_n����8"J:������T˂�-+~pG��L�( a�^�ۼy��O=��;�4��ʠ��H!G��S�c:j���ּy����O�,N��ﻚ�ȹlKCZ�F���]3a��ư~J�l2�%T�
!r8~�J/�{�Y &6��-�ε`���b]X��di2�����zob3��7�ER '��&?	$��aQ�Xfj`�}���-�p�rn��8R�B3@`?}���͚55��b�e%�@2�$jA��<�̩�F���!��7�a��G}�eƆ���bϵ�ݴc�Ɍ��TNg��i�7{l74�:��$Q�|�uˎ������
��{?����N{4\D�?~�L��Oش����<�f�Pm~(��X��A'36`�J��BA�f5�c����e���
ŉ�F�q}��`D���o,�	�F��쐋6�I{4u�YW�அ�0�d��b�|��~�m�8�/�bD�-�KKO1(RnJFB��/l�J���k��?Z)�����t���� Bn0��ߊt7�V)�rz�o��9Ǟ1A\���*�A�����_#l�ߏ��l�-�c9����:�sm\�M�	q����!�-�D�6�$�kPB�C�1?=���˓���.���G��d��w!��(� ���,��ovd$�MQ�_�X��h/�.�q3��Z�w4T����L
�g�V��q�t�\��
��PY$i[7s����ں��>ω��1�c�!K"Y���|O�AJ:�E/C!"�R�8�!�ީ@�ץzD�T�1���C$�Ü���dI��f
H����'-;0K�!��P$��?2D�L<R�@e/��S�>@�t�;�y�FV�k~�t<�i���)���tw4�4���ď���.ocd�d�fN��<5��p�;�ev�ł�y���ر�#���#�B?!�׎�+}�fO3m��I��\'r�:��uĪ�%}�<(`Rwgvt�?!s�M��L=���v��q�m+Z�*�_�J(�� �+��╴�A�D7���~�C���0�	?G*l��o�R~��"b*SeF��E#��Ru	��g��l\	a ڸ�q��d#�c�B����Ce�Tx��!�f
�cN��s���������@��=����K�Ul*R��D=i鎒��],�t��4���������T)��J�bE�S� �8�nI�c�b~R&�w`?�B����<pBp�W��Nn�g�n��Zۛ O�1KK��KphC�9����	']ȒY�
.j��;��f�b�ڒ���������xck?eS�g���������g#����p[
�o�)/���A��Z���0��P�{��8�	��!{��K������� ʦ?Ad�/�u$o��cm��KO?o�C$y�0��>n�@�0@ IFϯ��S�}�&������p��X@�/XK�BAZ��^}Ւ����~���	����oG��X��)Q���_���wF������)�ԺdQLɟ�w����s�v�u�r�����,L9��̇�	���㦙���pF�N}3Y-�ns�"��`�A��N9Y��W�=��E�UbH�*�**"�U#)��(0�zk�<��ܔ,g��~P���	�"�4����:��� �neU�Vh��`�����`,���2;2�(�x���$Oε!�PaʰwkS� ���I���{�ı!����HAB�3U�ܚ�s�g��ƂHuCe��g�n5����'�c�"��ȟ�D(k�Zd��2����Q��a�݊�D��x����8ۅm�&b�7�W���x�$KA�-Q��{������ś�T�t�ē��Ї�{�頋3�j�o��A��+��Z�֜g���3Rzf.���Wtⵠ�<`�h>�3����Vn�`��l&���8��;MC޵��E���'Mk5M�����m���+�SO
�	kߏ��8Po�8�g�)� 2x�^�hA�G�t���L;�p�[�[ �����2>,�s�y�l�����HF:�����k�m�A�vWB�S��7��ہ�`>��H�_�d��~)F��ޠ���h��+H���(3&���	5���! #(���Zi.��0d�s̠)��:�۱WC�Ω]����^1��|���z�S[(�Z�6���b�8�}���2F�����e"�$#��ɖ֧��L	���R⃅[�*�j�l��(�5�њ�W���
Қ_y?�c��䈯��xP�ePjYt1þw3H3O2���fk���v_f���w{��f�5����,�����:���$I��)���8ë�D���2
Z��`��R��8@F���h:|���k*����  �A������Q5���dOD�,�-a9}rʁ�A�o>�Kk5��5�`M1�'��Ez���O�.���	}ʹ*��Xߖ���۴��F�dmp��X��SO�xbR�6~��%/��?�УV2��ēW45w_�]7V$7;H8����a�eBI�\d�̢{X>4���>���T���l$��8���/g�A�&2j}Ye+� }���-��Xu��	�*P�~HZD�L�8����L=��@���^��A_�Έ�(�I�!�_a�}|c�W��~(a6ڃ�>ơBdS���pQTX"������$��@�I�L"�HI1���$��� �~ImI+����,;�6���v�u��\��$9�<��ym�	̀Bu9�M�q�`Hu?$���?0 �X�@���	�
�I*Agߩ��F�)�:�J���_��*�������<��#v�T`�<|�D�V��;&��r�=�4��Ꮶ���u�M2�������	�b�f�E�������IU"��>m��I�lo� h2�a�E~A;��:@G(�ׅ���?w8v���p���`���*��Z �$¥~��l�?_D=���wr�����J� 0�7��|(��4h:<� ��f�M[;er������͖�dF�\���k�}�E��z$���D�S΂y����-lC�c&F�{���ԇ[����]磁�l�� ���F�3����#ؚ3�?a��D8�B�{w��S����@�R��a5��-�r��#��ڭ`�vp�[{H[>��] kh���DU���΃ ���갬I/���$aQ�����m�����P�l:;�ofO+9l1(���ٜI���X�����d�iz�!�9	���VNcU@��>�oplm��*b`�Lf��������|�h� (�FA�EEU)ݤ������?G�$=2/����$���zHQ����<*tEvb�&�6��v3�0�ӥTyY�i�YDL~��O���8��z�
�/���a��C�������V_cݹ?#�� 0i��#^)�����Խd��}�~K6�c�Y�Ncϯ兵��#!E�1��n��ױ�Y�%���X�3����"�j-+��z����?j��]d 6H`�~�����Ѿ~�3z�?{�|������.j�Ն�����'�Id/?��~k�O'Xq�Q���_8�{�s��wOH����@	XY;��2�*k/5ݚ�$��	{-X�H�~ˆ�LI-���X�"���_���ޡuI>�_�}�Dx��Ӷw`�xsb��Ʀ�3m�(����ˡ�-���`�K�Hx��5����=��}���/�g�N����)���=��������A�m H��j�:Xh7�4_�S��T��T��S|��@���<��P��N�M/RրR�Pr�yάp�K�*�mp�~�wzϷ�]��O����@T,�xo�8����A�8��7U��j�G�>���5��!�L��)|� Z�d��g�P�����=��B��w�V�3�$����(%=�hO4E"����"`>�l��ҩ{T�^4�n��ػ.��Jҁ3{I&��}vK-�{g�$�����F��I�#��=r1<���&��m��~�u�w0��nؿH��8yJ��y���b�����^s$���V]z��|�t{��U��mW_�����v��c7kwl��x�+�T5�~�H�&2��"L-������k� �?��љ$Ȳ<d�F���2�3��L�W����l�p�ՠ����';�/�K���f�k~rR����*����s�'�9�;�z@̚uC�z~�E~X���v�t��ܥ2C�'L�?t,�����T�us�k��9��y_�3I��O��ڵ�@�%�_���~��Φ�'Z���*���5��M�<!���EM�5��MT��>#|!M�]�썛��	~F랼�f|�� ,S�F+��?|���������*�����5��d!֙����-ᦸ������!M<�9�)�b��S窛�C�r*�ݼe�*ꪃv𫗰�?:�Q��=z��2�4F��"<�S;�s��u���7w����Ӣ#�l�ɟ�~c �5o�6�N���clĤ��\ϊ>j��Wh�W���,��;�y%�U2iY	X3V�ש�-i�p�¬�TP�M��V�`rE+������^z5�1�*��hU�4��%�L������0;P�'��_����xb

!I�C�ڼ��.8�T �}C�Q-T|�:Qk�O�q����q(	����~Ρ���� B(EE�>��������{����﷜�I�;�^�R�e��?H�7i'�ЉyW�R�t��H��|~�;[sT��p��5�����ꅦ5��ʶ(�����X�#}�(8O��� 2%�`�.i�|�*����^9�8�)�`QG�߰׮���[�k�TJ��f'��â8d��G'a��+�Զ��r���C���u��+�ѩ�w�$�?R�!�Cﷇ.�������>3��k��|t`#E�.'&:g�t��)�2f&�e��b��d��(j쇔��D�V��H��O8@A��ͻ�����c�AV��rJ�"��Z��/,�5j��d�rp@����`$|A$x�� 2 �w&r��ק���Җ�JήV�*V�X��u�!0\5�=YS�������w�O]_���a�k+���״k�;�~_^S����{��Y�a�ш�"+���g�{Q�nۘ���/�s����6Tq�/�D1�7��x�s�p��_dۉ��B:;G��Q��x/"�LF�}9L}�)����^��k�OFh;���/�:�:'f3��n����x+k��� !^����d�����L�4Lazf�|�(
���/���+�$���f_>>��)����V�͝O������߶���X{,F�ىbU�nN��Q��n	��BE,�L[���?K��EU�A�Vh����|r��^l�a�&&3����s\+Gan��f2Mm���g�K�c��!��,�ߴ����(����Ɩ������I��N��V��*gز�dشbob�դ�CZ�*�OG#��.`G2��R��,��.�`�!}lFj-]�td����^�F�?{��
��qF�:o�'� 2.G��z����ۙҳ4J��k����mL氦��8�,�'��bU�_$�����^r9 ��h����]���X�^�ҽ���d1����	$��Y��3���<��/.�]���g��l�ѿk㙯}�ݸ�0�A�b���QTH ��$� ?W��;Z���a�f��A�q����K����˹ק��>��(-�x���%S�ev]q�+(t�z�ܗf<��՚��boQ�3��j�����⶛�2ԃb'<X�=Z�:	�\�D���--�B67-QKʈ6��a�^nzlyfl����H��ű�t��'NA:��Iʪ��hAA�b���J$�<Q��bia91X t���9ۚ��}Ǿj�;�Q;�Tʵ�����f��˵��g�(��>c߶���߯<b~�d�� c  �({�n�mg�=�)����$����H��F)�t�!`�U�o�yX%����+Ѫ��Wژ<��Qj�}u��}+)���5Kf��˩yw��WK7v�B�E��/�玒N}us�dܻ�u���/;��������s�����O}�2�A"�ɏ�+�����5��I_�E���ެ���<@K�S�꒤`��xh	^ʋ�U{�o���wN�/��-��ב�u���ˉ�\H�9�g��ػ6���[SӡɠwUH�͒���p|GW���#t��+b����)x'`�ճ�d����%A���ʉ77y��o��S#�r�J��z�Y�3~�x�_f�z��\�;�mu��9�X�������#}���.sEX��)m<-�N4Ig�k���Iw�����.W,1zgT]���"���:�30�x6�E]��-�
��mЀA�zo'�o4N��K�3f�@��A!��{!\�RZ���'"����8��y!7VEYZ����qQۙh�J�<�20���[�w6���0��M�I>]ϴu�ޘI�����5��i�c֬�V�oT癒�n�K�;`t��\���{,���{'�7;��=�r�U]�[}�O,��+�b�}��f,+5qo2�1�
�+n��;"�Ǐ��=��6\�9u����_�5I�<
շf��1��CB���ܛ������6����?G�z��d�ss�>��:NM��A�d~�15ڤup]̡T})� �o��
�gÈ`�{���2�,�yK{J:��j�n�Zs1��u�[%톓n�2�����y��ћ��.�PR�isεMj̭N����{����mͮ,�ry�rD��M�ʿ��T��m��TM�[�}�=�4贶���s����C�n�T������L.}�u�Ż5�9�}(�[��̝`���o���Jw����W��y�{��Γ�1j��r�>�5\,w��&��ذP��9{��mi���k g&��mCA��l~�i������tw���rlX�f!��/�*깔j���Wn.:�ڳ��%���ð�L��]�^�+qa]U-!L3���CK^����O0tF���fY�
��(镍;Ap,�t���_�Փ~�߼>��ϲN�w]B�W@Z��ʍ�,i�5��'U��64�X�v��s���MŸs2rnJw�5��w����U�(��[(z�3_�!{}�4xO�y`t��a��E-���@�ڊ �1/a�Ri�+zrݘ-s��;2�B�|���.�d{���]Z�����.����0�^���i8�u��\t��YBAFh��r{yM�57�L7B����������Շge
�cMK���gy�'4<�h/�������	*lka�����@��q�:w�-=0V#t�/T '*l��N=�{��y��ӱ���ɛ�\�|�rR��9�{3�[�F��p|`Ǻ�)ų�n�jZ8�Kxq�V�Kw�$0��T�+�J7x����^������;��U嚿��{��Ӯ���`�����o��3�^;�:������Ը=Cpb�2��D��b����e�a�f�s��8�'�O��h��N3g����ėvL����O�[3&h���['�{xO�N"������9�Oڦ��V|$�&r�c}��ACv��J~�����v��������}s���q尩2�������V
����ʊ>�z}���!�:��LN�n̜DM������,�Q�����;��ld�/h{z�m�LH��{?��?}'�d�1�K�q�g�����%yJ"0;�4��ԓXo}ܩש�C�}���h@r�X�AE'xw$�ANaM�ha���C�~��j�@S�>���m�ɷ�4��*m�h_��ѩ%�l}�1�����	5�<>��#�Ϛ!�T����ן�.�v��3�����`m*}s�:���P��%d�h��*ԟ�;?XmR6�sW����"��=���'�/
�R�5�c�Ty�.�Y+��\E���Mj�s��i?��?&����œ����Wxq&��
�����m&-����LR��[�B�Z$S䛻�h)�c�a����޿�B�4�dX�繾m�@I�ޕ(|98[}���� ?T�A�O�~f�z���}�M�P�שr�{�0A�+"���T��k%d"�&��h�B��|�7��s����ꍠ�1˯���Ҥ[>�� ��n������f�i�^\�����QJa�U��� ����@�9I�=?RQ;*3��"y�O�'~͢�?'��D't�o{О�Kh=��?.��>DM�{.���HD=]s�J�z#;�KƬ�5����Â�>��xz#��H{p�8�6�.���!V��o�.o��	�3���T
ղtOJ[�L��|�wsU��e0��b AF
�EZ��Z���G�H�~n="'5�|���^�ޕXA]�1���� ���t�z#c�r�t��m.��3����d�
�i��ؗ���.���[v����w��ח�zK<��gC]�����0�Tc���֭5޸���dHw�?�?.���p%��g�b1+=Q ��M��eΡ���wR5�#q��u�l��B}"Ξ���)���J� �݌5��T	[E9�� 0`�A�A:�b��v�]u�k��D��}c��}O��>�C{���PAc�q����jf{,�����[���1��/:�٪�f�����*�z/���)+�H���w\�'�q3�����gK�[h$4�}��K�߭33l(�H4`X�͸7�.�YDb�ײ��|�ʌ�����D�A�^=���D��dJ��@k�l�J�-�o��녂4ׅ��,I�]Ox�Uy^V(��@3�S_$�/�ꏫS�ξov`iG޽���4�`���P�,��c�}s|�/��c~�W��K
�)J0h�o�����i=�t�������ω�x��>�%D��^4�Wڐ�{B$w�#���:�|�E��EB�3�-��*�;���sЈ�t���q�ʵPv�����vE����߹mA�����'aE'|�w����"/q+�F!ő�)]��5���gL����� ���%
LnOg�	��U%�� -�T��A�v����Y����Ӊ!R.Fez�B����9�g� �~���m���C����IM��P����&��I #�cS�Sw�*���Y���;t��A�|��Y��9�ŀp|B(�J���g~�ُ��3�2�Wegub��_e��d�I�CP�t��IK�%�j��K�%vr6;��lښ���Pg�hd�A���mI"?~,�iS���-�꣥m��F���m��70\�[�6�'��2b�{���ٺ��c�+ժv#�$R#�=��k�,ر~�>��p��4�����Ԣ����(Z}c`=a:����N�����e=0f1�a����z��>�����G��n&t����"��HD���oM�x�dP��N"ϑ�)E�s�>�++���a̢���k����(�cTDQIV(���?^�=��W��d�7E�R��{�8���V7��^�����L���;�XAɏ��9
�naN?%w��R�*{��F��gzg>G��xУ^&�<���=�1>�Eg�!J�YhI�	OG}�xF8��R��>r��,�Fb���0$�C��lgVz����u��s�5�@F^��!�S�S^������_y鋮��Q�x�z=��H���÷m�ܣՇ>UY�>�N��L�^���D�$����E�0��OǦVL��ga{�$���㮍���B����S𽙀x_]Ay���<�;���S�S�bw.��/�I�J&'8�/$���x#�J�A�RH�w�#�R�EZ�*,%��|>^�)ӕ��\���V�\4\���'�a9�GT��gЫƖI�$OZ�,H�u����&�_�]�5>$]$ICs;1d����ɝ���غ�緃n�Ú������9�__�ɐ�v
��)h��3����~���^�^�&q��þ׺�ޠ��\S	�9�o<j{M�~��2\ל��gD$Wd�ύ�5���y3'�Ђ�i�8^�5���^~�Z�*���T�d/�p=��?}� @����P<����T�q���t�6|�W�lQ�h��|�1Mh�ڇ��6|Z��jg��_�Rv��ࠄE<t���VB��ƞ!�/j�v���N��Ck�EO��?��^�Y��c-�r���YSzО\�3�qm�|��5@e?�~՗��e��Q	:*?,����bڊޱB�V�7��u0�7뜪0��2��v�om��m�(8�t�K>��~⎨.z'3����C��Ͷ�ͶCx��G�f\(��ٟ%��pj��P�O��nd��q��"V�0~Ҋ�fϝ�O����[���1rR�Bq��̠�;��̍��D7�h�;6� ��n��l=	���Y�kL�d�K�Z�<�OQ�5���.&ij��OQ��h��������#�؊>��Sy��ȝ|Ġ&&�x�y�iJ�ّ?H7c�jj��`��9��%��u�˜>F&�����Ƒ.S�W>���)u����Y4*�����8-J�"����z�eE�^��'"o������_o	�Y����׾���e���P�S�/-V�&ք.3��G�:�40�}��q8U�a	*�c<pw��6�o �}��՚�\ɡ���ҩM�1��ٜi�w�2JW\���]�c��y�$o��N�i��荭�=�Ӯ��p����b��(@p�U��V|9��YB7v��N�����A��s�&*����$m�(������Z��{W	����E�q��}Z����˙J���;�1Yh�@[�;KW@�P�hտ��?{s9=�\�<����:����O��Y I }ԭ����i\܈�$(�~��{��"uw����L����]U{2Z��/Q��8|G2�y�~ar\Ѽ�6�~!������帠���ʂ}ұK�4
�.�q�����C��i�����j�:�4B��l�$z�q)� ��!�rc�"�6��^ԶG2����&���Ψ�w�bn8�c�Gt��u��F���\5��S_}[BT�S����c���D�,�׍����"�1G�ט�v�RL��v�`�,+��2^���7�$�/���a��Q�/ǐ9����M
P&}'&ڱ��twz���
����S�_�~1.궰h�Fe�cy���H��Is�g�Y0y�+��|w�`�Z�oA�ru0%ģ��;�6=�g��-�T�^��t�Ř���8{���q��щ���pQ������}�9������z��צ�oU�S2�Q/�v�wW**�\˘Rr�Q�}�����$oaY�7^$�ӝ4l�H��p�z�lY7��&U��{�KaMV���Q�yYE��V�V�.���φI���ڟ�&p�3��ۼݝ1�!룏m�怣"�R{��Z*`a�'�J�K��j�}-�*U�K�9W�vErj}*L<��ekoqI;}CA9m�]���F��յm�mUFm�����Q$����r���Th'�Ћ���Vb�궙�&̤#O�C��
y�$[ᷳ6G�v|=�&G�S�#�^�jf��]:ۺ���g��ߦ�>t/�k䩁懖��#�g=�/J��a�}� R*!�)ðY���T�Z3Tw0E�{�	c�p@�[�+����Qy ��Ω�z���tA�ɝ ��Q�H���f�~�sꮹ�^�G�xc�/N��;����Έ���)s"��ԡYU���f��Lz<·�����<�΅LN��7s���.S&{6���I�"l�k��^w�/y#���Hț���10`�)5S�n�.�=�P
���>���C��]�JH��a�����>Ȑ}�>������t��>C=XD�/fas�V�z@��l2:dM��d��Ue�q|$��Sc@Za�CzQ��D�Ԏ�T ^�Jv����Ǖ�*���&a��POp��oG�I �}pz�i�9��k[��+��������}Q?`�(�U
^�w���9�8ϵ�ʩΟw��t6���~?}��p2y{�g����ҫb�gU4����S�w�ٰ���� ���1��U��`�	���۽���ow�w�m�v��\ߙ�cY�҅��E�j������w�W#@��ǵ���̺����%�����]a�\��������rϤ�K��T�e�ۓ;y!�X.�T݂���:��ΥM�����	7�����g��y����@RBG۸��O��>bbx!4g�#C~�z�?��FR�Y��s�T^35q�o��%	Z潿��bQ�1��h���2�YN�N�w���^�� ��x�^��RDѩ&�=�Ftԁ=}�4N�\a��\x<�o�>���MFb�MK�eA�b���`Q�r�������-e���ޏv㛣���h�^7`\��@��[��\��c��5���ʌ`b��C���}��͙�}R�J��j�GH&R'�3�1����u�ZS{�5Y�z"rL/C�	v��w�>��i��Ʈ�|I��	�Go�Ȉ�^!�9Q?��γk>����������u��=պ��=��k˞� �ǚ��4���0��5�f�������K T�Z�d���:����=0Q��)��>�9�ǎ�)�-9��y�����N)7�='��%���N���� �ERHo[��f<����r�ٻ����2j���3�t�k��{�OL�>�D�O:��:��<�'����y���	�U0�����U�>R���ü�T\g�GyR���v���_q�t(ۺdG�a�"�A\�͏i`�\��+T���.X=ͷ's5/ޯF*�<+ծ�8Ԍ'�t�Xq$E���()�ͷ�8�8�h�4�e�:����I�h�كG0�Ό�^���	b9�S�C6�br�Ϛ�.�����0�B8)um >����v�ԗ,1vߕ�	��\,ֳ��U@������d+�0'Gu��p�ɝS��Q�__b��L?��=�z�^�%��P��s[��ۨ�P:��m{���5շ�ՎB,}�	P���m���1�bj`?�f���\zl�DH�}#�����*V�|���Y>x!Bd����2_5oK=��O�Ŵ�EE�K��+��<·_N��Gz�ts���S��1�s���ӣ�h�H��S���I��H�H*�Cvh`tv�����m�i�-�/L@���'�C�P�m�lz�;��K�rNMʌ�ũ�>�[��f�i�B�P��>�Ņ�2�'%���#��ӕ� .Q�čQ}�����X��7�x5Q�|qy��*���*�!������v���^����������W\ z���o�i��P'>��o����֪��� ������7���n��k��+�^UY�B%/����|�Q��|/�U�J>�{<�pXw���T�����YrF�z�f+���#��P+I2���a���y���CY��w����I0�����DA����#�NۏZ��87����
�w��C��v5
�^I�y]z���1����eR�6Yc.ӹ����Η��,b�|�WHa^! A���XEPb�� �������P*>hfhr���[�k�.��om�vywb�1)P��L[���]m�⋖�`����R�a˫XK԰�EY����JΩP�1�k(����by��z�
�2�sG�dr
�z �BE�k��X��g�]*�A��z'Y��C��pt-(�]�g>Y�������R<+�_���c���^+� �ڋ�2��U�'��� ��V�o�n�M�.#:��U}b�iz ^��ؤ�"bma�y!5�u��hЩ��G9/{�e�#8{�	�++]����;�πwDP���F�vK6���F��$ގ���n#�o��{�{��4c-��D���c+$B�L����{6i�LÊ�B�.ͧ��(��U�R+ж�`R<�Z��}�0}���d�s�+�'�ig����H��x��ңWKT��-�S���f���x��X��Cw�"F�x����[�Zz,\GB�'l|O�6�-ܷ3�Sar��]�����S��n���� � �!�> s�,iS�
�QV�Gݱ��+��U����t*O�t����?)��gf.�-����lpq�U�^��՟rB���f�h��DUk:co�G�W�ډg9�{!Q�]�����v�g�����2b��|�O6��>�hi�YQ)j�i���7�H�((O�S�Z���7ؿi
@E�Q{�M�a}�-��\>{3�E���8r{���ƘI�K\y�º���Iw1
i�3#�7އ��fIW�,k��X�A�A���}�N��΅%'�ݝ�����h���>�n�oSZ噰b�%�0w��
0yp�,^7[μ�0�_qf�3Pv��@���$@T�+�І�V_e(��N�W�Q��X~�;;z_��׵[F�XDl=B�X߼Acnq4�*Y�(��B��&(��4H�WZPo��Ɏ��=O�=�������CWb�Z0,�.$q�ƪFT>K�J[�b�{!�F0����w��R�zW�كel���^=+�0��˔�W�P2���b��Z�I	���L���F3��z1k����E����6� �j��_r&�2%"�ָDy�u����!��0��#}��Qb��[�Y[Z�j�.��Q\,����|��*�r�� �=MLL�g�H�W�6ܟvO�л�=�ZY����N�9]����p�qM�*y}Qt,�4�(��gkvչ�d�扸`�%*�z!�t�����S�5�8�Iyg\#20h�7��r���gfK���.��QU�lD�Yb�4A>��j����Ӛ1�$X*�����τ�Lo�2Nt4to���m�a�=1�@���X���,���BE�"�	��
H`y��q��:��;RUR���4��C���g�@�{�ZF� �,ي�0�j6�a�>�G����ɘq&����7{������je۬*����3�ދ��ܹF���(� ����j����F��%]�g���IY�!���U�3�Of���ia�-�[N���^
���H)�X����{h���^	h��A�s����h�kpf'��f�y�J���8Nf�4T+фV�)�q.��ֈ{��k�`a.��A�{�BdG�G�Ǌ^�f��6TX�D�*Y�|�W�eR���+<\�Wq���ki����k1-��R�'�,�W����^�d�
�^��r|���=p�76�Υ��(��wz���b�iy�V9�]�^��B�bP]�9����ޣ���7�t���������^8<����d��e��7)�E�a�s���u9>s�g���iY�{" ��ыX�h�nтw"��������-)�̪�x�%���s�x����{h"q��x���w[]6�eɫH���k("h��ͺ	�v{�]/�d���d�=��,�4�rT����^�]�94�^�/�S�K"�k����1����M�������%��5���f����P��t���⭷{ծ7�g/J�=%���ۂZ_¿$� � �f��fg��M �3ҹ�]��'3� ����}��8���A���{=����DS�Nb��zb)>�)��k��b\�5Ҏ���	3�1GYF��n6�
��]�4}	D�>��@�ax�S��pYC�����ѓnr�r���SU�������f���]0r�s��r�r޵��Y��[�<]Ft銥k�����]��B��r1kN�H���*3K킸���f�v�C�u�7w�)�VW]�C;��K)[[����D�zM���`��n�{r�q�{ssW��`�-�(����R�L��d{'u��^��Ko�[LÛǫF�ML��x��nX����Uf��u�Z�L:J��d�8�Sx1��|o�$B�'���U��u2��=������vK��4����f?����}��}��u�胧��L!�6�@)�WxF���qCz�8PFĝZ��}9[��+�ג:Ӣ�-�{�9	�=�r����"���t�,���[{	]c��^�ܛS�}�:�-�Z*�A�e.���-�x�K��5����
�j�_PVVT�e.��	�AȚ���rf��T<ð��;�^�I�����P*�v���y6�=[`��`>�o=��>HE;��k��{���t�g�<�z��q�[�v��MbņͶ��{4��a��LS9n��w4���v0e3�2ӎ�v�ܷf��	v�[b롲�}-r�e�-x��ɧ�5�Y8�F��_dWu
�J|<��i��_o�$M���%�@��8��yh�ۂ�����^���L����>�`�	\�{�1:ؒ(t�5��+�}ɭ��{�:]J����|l��PT�K�yb�b���D���L�3d���7���X�z3�/����?}��Aڌ\V��NrDYbGV��*)��QF�MN8�e��U$E�7����m�Q9��/ c�5�0���С�\|"�?6��Žۯ�_�D哸�#�zȘZ|�ѭ_����qGA��Z�H��Y@�]��7�d�H�7��br�~�+�B���1�w��^��0���p��x���4p��v�+�K�A��`�ݗ�ݽ����<g=L+��}����R���2�f����S+'��Asr͹�1E�ez�=�:-�s2�ABV�ˊ�����k+ve\􎥪��Ԃ^�[S2�'�rV��>���|_�|NIH�?~��s��?�S(�N$�ઑ�M5��%��z�ʐ���{M����΋�	j͚�<pDp��u��c�+t�Z{پ=P��#w�kEG v���
�͛/��=#���ӟ*�᯺��WPW�����������L�o����N�n��H�et碏�1�="��u":3 LH�����w��2t���S5�����cha9)ϒ�Kw~���~}��^K�}�K������
��^=hiS��r�m�m�FU�4�;p-�n��3/g׻2���}�3��q OȐ~*��mf�����:�͓�sG�wZ��#;oq��N
}�/�H���Ө�{}�H��:d۳}�L�v<n��)�|g�r��«�5����۸JE���l<�M��qg6�4WB��Ac�A���F.9�"�*�O����#Yd�B��d%N<�C9X`Ek9Nh�SSc�]�g�y�{n+;�����e�j��ؼ�by�q��1'���˥�tb���1��H�ㅞ��ǧq+�/���|j#�(���]ݵU�.{�3�k�Xc��}}�'�ŏx��׏�_f9�/(#<Jx�H���0�ӕNJ�~��w�q�õN�1^�ʾ8�e3�H]�V���b�ζ8�v�ʥ����';ƍ�S��|":g��HV�xC�|Yc�:,<�1v���.���(O���j3��;[��pf�ׄ�c:j75�����p�?Q1
�L1��mP�����/@��|ù��}{���y���/z��_��:ɬCU�}�MV��Ic�x9|��t�ݯ򅝹�������J�ڹ;F'%����-&}����F��e����po��l,�~K��0�jү6�V�h���b�k'��=���LU*Jwt������F�c1��+�\q59	�dm���*��KuZPZ:�fLq��Gt��6���+	X�>�Ʀ�|�5B���-;�'���"�7s �uwT�7Ĥ$�/�����j�#-=��P�����=�c{���>}vY�5֨�I1�/U�=:���t�(_�Ts׼X���7�:jTl��{]�f.h��!����Ө}-a$g�h餍��\�} W�ޑ����1`��ȩs����$J>�����9h��aX�4�=>�%��;Ǿ@3Nj����=���R0���I�sRa�^�A3R*��~�����A�
-�G4��嫔��%ڼ�2�WϸL8��A�9q�Y���"YE{���z��\�Ƥp^:d3!��b�Io�xFK�B�eKAbz�82�b�8����g������῵�~�����������^n$����R�gG�����@ ��7a|ީ(
�Ө�I۔լHl{ҟ��܀�V���\$Cfo�����eh�␱���.;zp��~�F��M�S�B���jCZLc�w��~��s�r>�gLǗ��l;8:e?Zd�mgI2#a��f�u�����ҩS��B����=C�	7�2�#�]��u���I� u�����Q���~�߀�c��O���a�{r��Ci�'X;�J�S��,��@���4ωޓ16b�s(��6e��dY��=>���ܝz�w����R�`��Dl6�����;���Zuk��au`��D��d��@��K&�.�Kr6���o��uڝ�����Q�f<eg�n������lM�0�F;1n���f�]s��`(ȇ���w�1��L���8o�]׊��o�=��7�F
{;Z1�R0�Ex���^�����:%\{��L�|ф.��������jd���s;����d��'������ȟ����z��L���W'Λ�����J�W0�:�{D�s��E.��QJ�	$��T���s��fFD��	�l#;~� ||)B�4����%z	dl("��"�力&n������ �)������J1�)�'��nX�Ic�q���XJ�]w����Ȯ���kw3�=E���P��&U�{�^��"�ḴF�S�����������Ʀ?KS���h��9�#�tL�����9�G�0���R���t�w�$)��?~|3{i	��[�Ey����!5ZJ�h��J���iD!��j䱋�λɜ��a���<�Ή�������A�s	���뛖���!I��S��9�ߴ�Pf���O�4½v�9GQ�mu��k��c/���(z��q5p���C๤>�Q�Ș�#�v������춇T�X�	�� ����&@���Uz~Ϙ��쥋�{T�Oz���M�Q�y)
�2=]b�Ra?^OR3; Q͌�ln��4����?���G�lw�]�����6�NP��\qB�9�,���}		6������w9�+���{<��z�z�cy߽�\��nU���F�d6�wN��喳����g�9/����:�����������
�B�����gU�\3�b�9F\���]�c3�'�P'w!���aQ�n�S�t�?xbƦ��w͘]��'I�}a�=�<��^��Ì�F2�ۧx��gi]�{;X㈙�C�1.��ks�>�!�X�W���VGt+�>��������5Kf����aߪ��W�ec�;*='���ִ-ЮP�O��Cj�{�l���>�G�lae�_�H�_�%������3��٦ܚ�BM]Cr+I15�����\�s��+w2{W��O3-n��L	SV
�{[.�j�^4���]�O����a����_8;I��p�[���x�5��=����{"��} �jKn����}/���<iƖ+c%���QGf�z�_eu���l�}vn��Mj��|W�b�Tp�P3�^T���R�L�X�n�j���������ʫ�3{�n��<�a�������;���_s!	��-��=�����ۂH��3B�pͯP{��27��;�)�oJT�+�N�5��`gu3N��^O���o�σ^�XY�s]���.=����7�*�kt���z:Q�>�uBF.Wg� ��My"�3{�)LwG�O��{=+(�ד�Y�q��4���*�׽�}3^��P����92�̺�����c/m	q��@9��{)��#�T��T�����,r3C���+A��<F;��[�7F�N��{��i�j�7�GfU����z��sJ͙q�>���}R��u._�����.ۮ��P� d_'��gN{ZD��RN"�ͷ���O���ڎ�OƯ[Q�pp6��C���F��R�8v��ج��k(�������'<����O�l�M嚜��s5�V{�F�z�%�_H�WτA��^H�iLt�����G� �H(`����O[��@�������j�.YdT>�TO�n<�B5*L^2<��g=)�&�rkl����^A�g���g}D1����d�K�{����ڧ�:��o~��ɟo�Lj���dE����H�7�=T�2�`�ﰑ�)����~�}[��a����-�o3���z�p8�A^���$�؁[����ݵ3���k��x	������ې�����Q[ޣ� `��)�ѥn��FEYD�-�L� 賜b�+�gR�����g��M����EEI����ǘ=��{l�~�*"|Ƌ/۲=KǻdXz�|֐eB��t�2�L�n7xP���}�}j���e]�����1�)�ގ�-��Z0�\<Nو�D�X��UQ�T��	�Fr�2�	��N.��KЩ����2�Y�ۛ���쥪v�I����at�/��/3�/PD��복x09CN*IĚ���{�p��{�u�m��b������Y��{+3�GP�W&�fkz����lu'K�s�t��op�f7e�d����:��׻x�
5Ȍ'e�MI���������d�ï*b�u����N��zW�:�5��UGT�}�+P��C&�oI���W3��R~�ߔ���0�p���`�;(�E�s�(>��� ���wdJ^�;��̦{��sw�ԁ�����fk5W^yl�g��Zb`�e?,���ĳ٘���]��Ǉr+��Q>�H��Rمp'x�mq�]]Y~�T+	hx{</��MRts~�H���C�P��ϭ�-���q`PxWp�ُh(�}�u]H�f�g��#�9q��ۙ�k��ؗ�G<ƞ�ԣ{Ѧ�U�����%^�ib�ґ�ߤ��|�EW.�@�a&u���en����ns��U��Ԅ�|�q��^�p���F�&�]Y��J�2>ͅ�����>��W�&Z�:X���tV�9^�M7�y84�ۺ�UH-���\d*��������_|Uϧ���R�M�թA	n��i�,��YO8MT�Z�pƤ�<YC>᪪�n�;��
������M��>��%�%��ǯ.ڥ�� �WGb�/H�Zxk"�LŪ�D��2�=�Y�\���| ���:'M���Htw�ˌC����h�5����>�7e^ҲI�@�4Qz�@H�E�Xi*I>aP�U�8i-^*����pT�3�h}PӔn��1�br�H����7'//u>�(��<X��Q��F��o����8�j���kf=<�!b��y�>\l�����c�<F���o�&>���u{;R�\���l�Æ3v(�#;]=+��p힮��x��7�9��`�J��	K��UT3��D�dnܫ��A�nK�q�{v���}�̾��K(Y�ohg�Ә������d�oA�7Z���yS�2w�ͽ*�D�]I��'���0 tf�~K"�]7+9nUMu���v�X�p�V�h�L#�${!'�1{���}��n��hC������yx/a�'F�04�Tuy�=s9��5Dr�wR�i�+�}Ѵ�v��f'v��Tǁ�`y���^�9�1�'��a�vY������`z�1�}�9U${�J[�|N��yD���;�YNǳJ�"D��x�ܮ`!r}�O�3�x~K���-��Kq��*�#�1�Ù��g��N����a��=�D� �f2��4N�VW�۩ЍJ��.�t��N��d��O���ي�(��3Cô��]h�7X3�b�1Y��8�8:7eE'����5���A-��m�tQ;���&���=��k�����Տ��S�'�~�>S��h�ؤ���S�q�w9�t��R�^�l.%v7<��3�!H����$�v;��R���C<��L���4�����ᯪ��Se�;W;A޽
�έ��ѻ������yH�e��'5�v|a-e�y$~$U��RM�*S֤�4�E�B�/���_�L��;/�RUa�@/� � ���˫�����^Ϯ�g��bX�Or
<�D�<E@�x�����\]s΄^� �+�z����q鏮�*����;*��|���Ρ�P�݃��{� ؑVǩS]�Ӟ'����M�|F�x�|��8G��{;"1�����j �d����u��v�T-�&�\�u�2-SX]>6�"�E��B��������5wIN\��4C�h;�Mǌ�>i�ࣨȳ�1t
����/��H�'�<9�	�I1��@G��^����+�x`��|*[3P�9G\Nc7bI1�*dI�!d.M�>�ۋ��*�H��K�zħ{�G�N�	y1��lofU��1Bl������{������7�u�'oz=�\���_�4��e�]{n�I�<�W:�oc����WXlo՘T��Bڣ��=k�7�>�:��0��d!2v�fl�ˋď2&����4��g��.�B��#î������|FW�U�获1���s�9n(����=~S�g�1Cpm�d�����/m_��{;؞.���������D���Ɏl<�[����v��o1��<��}��ڸ9�����^�t���V�{����q)�2�$s��sf�&�6�aM{#
���p8��a-���'O�UR{d��ג�Y�����2�U +6�����}�N}�<���q�����G��xF���*��_�'�7s����/���{��V�%���������v����yw�4�:�w�C�ԈO7鮥Zo\��wzc������k�|�sY�G@ǫ��ѳH��)�1)x����c�~�����Q��&��sL{�4�>���k~�c���3�C�{~Ȃ!�4�ք�~�|Y��\��Q�8�|�'�rt��ZOر�{^���u��է�W�������e�G#����p ����,�����
1�}�SQ��K��i���T�:�o;�M����+ b�}��'��=��������u��}}��,�VLx��=1Hu칒<�ĉ��Ց~�� ���=V+ٮgq�]6�������C���x�9�}S���W��{j~d�W �qߕ��w�H؄wݵĳ=rG{�R�-��t����6��ޫ�b:e2_M��\S������G���7�7n��4����UL�E�0��)�%Z>�
���v�TUA��-��++X�srԍ����M�J�κW�do4pW�)���dL�]�:�w5��p@��(v۶j��PX�V�"�E6鎔;��bWl��..�'�]�˭�9�՜7EN�� �z��&��D}���O������x�T���X��$u�WD+���o^�N�/�~�Z���] ܾ�j�P�/w�L�L�����Y� �H$�R��c�0�Q���qIq4�&��W�#v|#��n�L" LH�����;��ge^k�����=��ИǚA���ny��Ry�&�4'&�*�Т�]]�i�����YG:���帆����r��n%�裭FG;o-/��p�t�ԣk�B'j�ك��	^�t4��Y�}��a��hAi�]����nu2K�)�l��Bם��1!�C�s|�rX�d�s��v3��A,ɀYeI�^A�]}�1�o�����L��;W���I�m�����qe��n�����"͌Wm�bp�K��R)#�|�8�F08���y�B"�j4��w��Aү@躖�5m˨��+iaJ&�XwBͫ�<�FW��f��B�SV�P���h47�SOӴ=�y��VU��!�V&XZ��aL���-C	`_y"97I��oH��-G%M3�%)��I,k`bF�
L`��iii��_���6�w���,I����H��"�0�������SN�]�b�MJ�n	 �̒~!!#�<��=�v̳%e�ͼ�Om����#���<T|*\�PI�:Eu�N����mL��ao������]	�`:�F�S/l�wwW���:L��L�	[�\e0*LP嫦F��ji�ִq��N�m�^h��,i�a�a�\٘I�˝���#Zk0V�N�gl٫���U(@���9N}=�OX�bzX���;e�]�ɴc.	y}+'v�ҵ��޵�l�\���^�q���M��х�U�1ɷ�:�P��aBtB�/fX'36E�&�d
�A�γ@�b�����s��`��֌��S0��:5}�8S�z�jց��<�4w0K�Ŗ�C�}_�¡��/��r<:��=�֧'�x�ʗj�SK���r!we;��e��vC�?�%��w���i���3�ᯒ�6��u�uu~�8���Gr�9��=���/����Ⱦُ��2vń��ϹX�ӻ3�ʵ���S�(3�y�<{V�:�m��Ӌ�޻�e�v9�qm�Ђ����)/L�:;4>Ru�i屎F�ok�_f�Kmq�L�v�bݜ��sIW��Q�.깽v̍S6%�^XG�n���dj!ti�Ew9MY�s�ML�ZKʖWZz��/nq��YN�"������2=]�7�������a͡�o.��������@�bͤ&f��n�gm��c���z�TE�[{ �o$�D�S�S9�iK�jfJX�J�iX��(�܃af�Y<�P+��������fH�l��w1j��ɒ���:]��{�R�M�uR��j�3g��8���8-�S]����]��dʌ�]�A��3����$���lglG�'0#�O�^��%��&N�k�A��|<��Ȟ�U*���n��0�.{�^��ϛϊY��c3.���	S�l#.�t}$�>o<zy)}�T��l�b/�M{�}=�x��$|��.�+�Ns��>ڨ�y��L5˸�V�]¬��#`uUUl�:�6/ב筑�DW�= )�J}L�ۈsn�KCȹ0�6������w�������c�
u�]�hj�<�ܛC��:��]u�!J���#��G�(���0�ZW��{��b�0#{P����=/M��	����c�2��f�pΫ���٪�6> >�}�2蛾���~� cտ�׵����~��½�Č��ħ�W�Hۊ�B����$�U̾����5s�.T$H�V���4��z���-=�k��}\S��)K��#+t8ڣv��X�Ar����٭ku_,Ɲ��0�s�Ώeݑ"��yʃ��yv��U��C�9�8��g�$�ƻ}5���$-�~W:d�u�v�7M#":�9��`����-vu��\��O��[�@�W�ɛ1��3�tW�ә=�=�N(���m��u�$���j��}��ڵ�`s���%�*�ќ�'8�+z���� H#�>��ZT
��{
/��I3#6��+[ڲ�Bي�o�7��c���O�a����t�^�ٕ1�l��)�U�����nI�kk��H~�hM��|��:��)n������ԁ5��Y6����(�W���]�jg���v}f��O��5J�n����|G���Cs�{�Qr��p����]C�Žst��w���J.<vvC����#����Ԛq�3)�o�}�u��Y]ݪ#ԶRו���-��N������5��z���f�˙J�F�X�EI���9�k��E��,��
I"�}W9>�߲;��{
�;ghE�hX�<z��#հ��೵D� w���6�r�y���G�Ϟ�I�.'�2���mz�����2��U)!?������W���s��&�T!��Q����ڊCLyg����9�}��k~�qA�^��|�t1��42�C�YG@U��9�T�"yI!�O���JB��j#�c�%CO�h��q5��׎!�v��j[t�$WG*�r�uϴ�9GE7)=ib�z�4��C�C{֮���~�*�~>:� ��=�7_����_�㽉7У���c��#O��N���5��g��4-���ˡ�o��f��������j�!�0WL��r �w�x�����-���~:q��60c{3��f(q}�Uz!���vϝ��M�9�q��F8C�#g
��k^�&�����A�G�=�g�wz��P�gz.�xL�;�~1�o�8\�p�7�Ix�6& E`�� ���ӆw}jd���'�YlӞi���|r�F�o*x!q��p���X��W�H��*����!Y�
��$���*�0#}�*+b�<�>�p}���{�J�?W�:�N��`֒0�#o�{��]e�mט"��v���n�Z���\�:*#�����$e\PP�=3v���Y����:mz�z0����>�Ȝ�����|�8&.�Zy]���o���W��C��?p�~+�� g��������vawL�¯���"�
��Ԕc!O"ô�#��%z@"$n�3��|a�##�7$��6f���Lg�O�Z�Sj�_Fߌk<���?tN5����~���x�ur3��k޳S�b�.s/��V5��cj��d�9����B����|��&n,KY�c�	}�휨y���m�+��pH��g��.�������9�o7C>��?_`�����a�d%�������}�ޗw�>�ӿ�ݺ��� ��Q&�P���]%�Ѥ^�=S��6w����Z}e�xS]��s���:v�ř|ru�l��C^��K�x�uB�0�*�Շ1��C��w6��� �GdjQoYQh_k�ǔJ�[�gt�o�aOpZ��?�p�ȷ*oMx���V��+��0(�}�#�5k�<DP�xW{H��>�6 ܸ��߶v��!:����SUܢ��yr� i���)>��e�v${�VTf�!2'��[5s�׫�g�aD8���(���zͯ^�{D^��Or�V-�H��9��X�T�*�J��H�6�[�Q�,�	Վ�U�;
ۏ1Sf������b��>��v��㹛؜�᛾��.��8vG�ף��u�T����G�����c�p�32�)�n	�'\�F6��h��J���H��
�6�ߞl�-�|qY�T3_�U-���/������}�k��β8�zɫ~S�0��|<W�&��IvY�O�o'��2t${+�ǖ39�>/SK���O�mF��5�yUA2��P����f��Gcwa׌��7t�1�����@l(�ﶬ|��C�#}ְ�\�*��P Ǣ�H�1N�������Pv�,ETe��Ɏ2����<m��m�x���K�~9�}��,s�ԃ\.�7���RJ�����f9;�E�����`�aS��	'�rzw{�^�w@���g�^�u�x�ϥg���EN����yn���lɥ��{n�����w��������AZ+��F��s}Z�������#:��arܗ KjlOn\����>G���(�w(OWo�� Kj�QE!޹���4U[�}Pu�S'�sn�7,R���{�=�Ƃoہi�W^�U�jҚ��k�EU�#(a[���ߠq�Xx�rsѻ��r�8�N��",��j����π�5s>:.��b���ύ����+�E�H�K�ٸW���<������xz��+q�Tϟ�ý#_���g��bOG�������Y�L�΁�*�p+7����)�">N)�T�)��Gm�c ΀_8�e���kbu���<k�z��`7�3�4`�7�/eK�ĦH�'_�E�6m٪��Ӱ}��?��j��|���*�V�{R�X9���8uzz�L$���d�װ����i�=�"�mF!�~oqƚ��w-�����I9� �E;��EW���U��ޕ�Kf�@�>����M4k�`���Y����9�����b;5�y���$v�����Y/jg$M�b�Ug`�7^�6E�������h�h\ϳ�ja�T<�H�9�/n�'S�2���nj�d����;6���]�t{rT�Ӭ�܎_u�Dm��n��Ac�ۯz���.�U�����c��̖�p-Yc�ғ#|n�:rұ���/T��Nojf�w������S鄻0cǵ�wZ�I�ٮY.�!������_����E[��]�}�<�o�R��*�N7B��Ŕ�-��c���ݎ;b0���x��=+k9Qs��]y!�L��+�ڡ0{:�T���n' 7�(b��r���|>6}=� z�?;�����}k�B˖%m@T�q�{X�0�V��\�r{��LHJ�;˺�����gt���Mb�w�������ih��G�mAxn��J�k5�F�yT����>�|B>���V�0)�5�ȉ�d4X
%�yF�{���*�=?W/y�h��Vd9P���bD�?i��W����w}c]�3��72�
��_+�Ȋ�ȴ'�� W��.f��@f>��)���5P3�#��Yw5yB<�W-����$�y�4�+%�j�\Y�c�*�|eF�������=5c�I�_�W�n�k]��3����WW��*᮫Ճ�k�r`��o�hB6���9�{�GE�-a�Y�!*�������9���M��.������0����/il�Sa�6sk�p�+��#щ_$9����|x|�쓷�{N���og(^/K���h��"�����O�v�̽�0�2<�� g�@���n����a��M���'dT���͈o�AC��VJԐ�%bŐ˪�U�?��.�Z�U�~��粮u�"�<��[s"q����)�q�O��x��2��n�
8��8h���!ܸ�Ea�t3���2��X�� �<?�hx�胕ng���ά�>]��H>s�ד���U���o��\��]�!����h� �[��ۍ���J�9��Y���xB����G�n8}�Uq5�rz�;x\�9s�G>#�*#��+h.�-�s��cc��Dx��Ļډ�ȗ��x�ɼ�>`���y�|�?}����Rp�2N��[7{��X�o�ta�ǎU�F���_�{�������.f/`�l�D�-��Y�ʷ���cWx�mm��*� �1y�"-{�_�E�
�|��C3�:�g��3�ToD��5�6=�M��C	z��`yb+��'���[W��m?L��YJb�ǒ܂��6�>#o�G�O�w��t{�����/w����gJDb�B,��~�Z��v�=���H[
������+��4\zkr�]8��]�pVەJ���Tp�Mm�8{��Q�,�$&����jۏ��֒g�����vzn�K�x�A���*X��7��.�B=��)���ҧPƁ�L�%:�Y�1EG6�ڬښKQ��Fj����z�'�6��� �&��˝�Ǚα��}�f�K�ف�8Z+(���ok]�%g8%���>���;�ڊI��2���]v���Ha�e�R�W_l���ڣ�����hk��_-Ī�ڈ-w���)�'�A�g���F\�Q��)K���ʬHD�	F�|y*��.yԊ�s�Jb��@�ڰb���m�]�d0���`tK��s�]r�V��:�گ�� 1t-��Y�c�ﻘ�s���k�GB�o7���^���oj��X�G��x,'&��D�KkTWh�b�������+��#��.s�c�i�9�"�b_v�+;�3F�[8�9����7cî\���щ	Pf0���|{'�k�!8�����8g�{u�j��S�|õ4��n_o�����a��g��W3�6`�3�u��.��{���.��{��=�쀲�&t��������$��s�l�^��y���c�'f/���wS7#=�{�K�!�:\�&���w"�uS̸}�0h��#�dO��/��S��R�(��'Z�{����m�H&|��ހs\�#�41���
�&����s@�;W%o%Q����2��N��/���r�:�f��.�n�G6МnMW�H�@�s�]�����O����=������?`�Sjv��Ƕ' v�[��&Jw7l����,��Wk��s�v���,�]��{��`~��\G{�}�|u�q�d)�_u�)w�Ð�"S�n^hU7ݤ��`룦rk�q�}�������hc�����M;��ƟN������NӅz:��>Yq����77�U���54}� oR�
+�+�RZ��WC��^�]T���;1eM�=p��,8{��a�\��58�B�j+�2�F�}/���P�� ͞ܬ��
���p�����\�0õ���g1�qmv�g}��+��44��9��{�qǈ����z��S�^�#�p�v��|�WE��T�]��[1���Df�Y�0��oI���3I)�b=�ɸ>|�Le��H\v��Ms��W�����ř�zyN�ؽ��z�E�vt��m�5<!(����e����Nr~��!�W"oG� q
�^�QT������R��uo�5B�v��U)��c'��_	x+!4L(��?l��d�Hp�LF@��[�f�l�gz$���"R�ލT�h4A�����۱0xy蟓��3��1	��c����
rsM�HQ�wQꗂ=j=%�ސ���+�L1�i��5�l��$+2�����^���K�D�=�ˈY1�ݵ���!�򶳜�S�>�N_��(�oD�����k&Q�.>�P�أ�? N�Qۼ�y�WE6�zK��!����N��,m�{|I�1t	�pF�>!g�j���6�e��5�r�@�WG�:Ꚏ�_\�=3��[(�s����ыަ�0kN\�.�j�̼=�j[\�\���测W>�{�u�f�8��I�W�����+^N[�=��l몳g=l�]�EJ�S�(õ���ݸX]��aT�m��2�z�M�{���UƐkK��p*����DT1���4Ű��`m	�fč
aɣ���u��
�9S ��������n�4��鏾�`Ⱥpb�.�oHz<k��~��2�K;Q�����ԁ�js�M,���\I��c������-=����بuw$� �ΨI߳ ���#�p�7si�lDr����Z
�#<��>3}ayJ*ߛ8"�kq�`��-fl���b���:mMS6f9�0|��<;�L�G��HE$(�y��/�Meޝ��tV_�$�=�b�R�)kkQU�:΁<#f��(ŧ�)g���{�t��
�m����z�3hH�4j����{��s�����ڤ�r��2�\p��l${�݁� �=:e�P-�.S/c�M�΍9aB��wyj����{JpgC&Cs����ⷊ�79��o��}^Cf6��U�i5t�=�5zC�m�y�p�OpŰwN�L�����tU���g�oz6t�m��{У��$��p�t�Q3��;ט�ҏ���U8T.7�7 ]} K+�k�$�.�c��;5:O����N�2�NFǚ����Y����S,r�O��2�L���Q��j�,��k���փ�e�gL*ۏm��f乯��o�(}u��'X���ф'�gz���K�U�O��m��ъ�u��:g�ች������F�Ѡ���(--֮�kW���v���1�	�)�<�#|[Q~e�=Įf�0����ù|)�c��F��Ak�`s�.��QoL86�e�Q�MJP0wM'��U����Q[����5�Q�=@�/��L���3�Olw��cf��L�g�����i����0��6���d�t3z &6���J�k[�f����<U3&�W5ڹ�0���k�y8p�v��v��9�%��ؙ%;�}�݋dS�}xv�>+�\(ޜ����>����Y�:oVnJ�<�u�[h�<0���4vl����֠���pC�"6�ӊ������f�ꜟ]�B6�=��3M��f�N��j6��}���U3��W%���p ��A��\�f3�d��<P?�<8G����zX7���ɲ�Ycc���ӫ�n�}�x�_��3��Q�[�����0�U�9��Ր"2��1��bb/�g-��������Gt�i����zѵ#i��4+-�x��@�(oK�@Q|g��&f������,��͹0���Bw|�ܑȕ������\˝�tfpS�����,꺣l��ffó�wg�!����>�ǚ������j�=O�a8im��v���-Ý�!t�}a���=�i�ݜfyuDtM�v�30�Q��t��Vk'����rd.,�d��Y��H]<{��/�v��fSi��FH�\^[���`FS��qxv$p�n-���:V�:4�b",��{.^�D��3ؾ�ޛZn�
�L�29={�p��dٞ�L+���������E��	|&#Nt��y�͍��3[�J��Q4�Ӑ%}J�e0��˺マ��/r��]YЎ�q��q(��kd�^�֝�[b�{|z.�^i%����>��#��W�3���p��0UA���I�þ9��\+�')�.���W�I�#�NE��=�{�X(�G�Xlo�o__p��Єy���Wr��Lbt/7��u{W���8��	���xW���>[+��ٚF�yzϺ�t9����u𗧖��=q�	�򛲌w�(�r�Q���"�u�ܿk�fBE*2���*R�C�Yt	��)�8)��NL[��R��{�50L��U���`\'e�}N�އ�/���X_���J��f��V�^���	8�I����BYY]�J��Zj�s̜}`!߽���%�|�B�!����vN^+.�^�Wb$��
�"R�5���X�oww̩|�w6�-j����	;�q���7�"��0Х_Y������V$�?ýy<�d>յ]�b���y�c(��\dq�S���ǐ��S˨�mFE�KE��-mЂn����Y�|愼���f�0A�:��7�.�I����T������}�צ2P�k������{�yּ!���z�bv�h���:f,C��wo���,q��A��\v��B��T��`��v%��F�S�9��3ԇ�:�~��X��Ũ��x�>�rz������E��R�#�$���dS���w`��*bEn�~�Ȫ@�u���{8����>O�E�;�\�/��F؍}|��OM��)�304�7��ļnV�Y��`o?Y¾��Y�GH�+��� =/��������YgR�+���h��xW�������{
�}ճO��U1]�xd�e����g���{G��1�� Ͷ�w���fќ�ղ
����~�4=�Sg|9��̎�'{h�gFh����jٌh>R2}u#:�sg��YZb��C�e�,���@I�Ǽ>�H�GLsZ�x�d���ٹr*NE!f�J��K���Y�qy��/�$���4B���E��ssv��e�K7L�i����c���!#_�����F�Ï��Ζ0�q�B�/�[ں�SJ��U}���(GǓ��߭o��g.�y{#nO�sv��@nϻP�IV��D��I�,-�2�18//HU2].kh�����C�P�e�;�2fLp}Ԓw��]����d����o5�=�߮�:���o6�.W�y��E�>��~�z�ˡ{R�c�a՝u&:,�W�<oIv�M���f�������R3YĈ���c���;�-s�gC�rnL���t�x;�
���ȸ�[�S�d��sx������d	G�b��!{W�I����h�i�b&���V�Ty��t��d��ɍ�S����}���Bt�����
Wx:V� G�������Q��y�(�j4�Ҡ]c��^�u������I�=���Wy���멦/v��Z��@���0��L�?1������ܧ���:�1�T�EGm}���W9�0��x܆��Ǽ��J{��[��[��y�,�#�6"$�}�p6���Uv<R�ʂ9�f^jwF��$�v�Dzk���;��10cDM��  �|S��|6ǈ"��^��$�&#�b�Ɛe�Usf`P�����u�f��eM�/{���%�K^������v�씫���:nH��}���
^�k��Fq�uozA�,�yod�"{�gj�
�n�1�חh8�,E�!�B����3�4�w��/��;���2��L�z�q�Y�b]��=�׶K-(n�W�r>�V�͢�0TL�nq���|�f��n�ϲ'�v&����n/�b�w���Vm��q�D;}r��\�]�����[�|)`��uǖд�n޹�{ט!���݊�D�"��,�>T�����ԝE�� �د��X*��y#ڷ��+|��d-U-t�\3�0p�;�1��n&�4��W�5�~<u�0�=�a����2T/ҜX��9yn��~�wҸ��Z^���f3��M*�E���0��C�����of!磻]����>d�}��I���ޚ�ڋ~p�|�L0��@�po.�z%�鬵1�80��z�b�k�m�������ʹ�h]I�f�����D�j�l2�uK�P��F�\2Ps�K]Ѱۊ��j7��N�F���i>���U���	-�ޖ�ć���d��Mӥj�{T���Y�������`Wj�O���s�I�2���=��Gt��n�L�>��w2okM_������?�����L��{�/�l�>?C�����e�:�X$E�def�XVa~�~?S�|_��2'�@�َ��Qs❇N �*�]�i��Ɇ��]��#���]'��*%2Nƻ���{�H���5� ���P�S������>[����%O�C��9FP�_���gO�H E!��-�����B{Ǳ���H �z��j�YC)��S�����ʟ;'ֽ諑d��@�#�,�c��5��*x��n������]���H�r,W�����������Z�xFm��A��s6o=��c��X$]9өA�|��}�
�NEtA����w�T��]��:��vUQ]ObK!�v����#���7�U�SU�ѵ����쎎;�1�[$s�U�-�Ο�������#{z�0�^�j�M��=|bl��C�/�x�gB�~S�~�'q����l�p-�j��_��ss{�����T�Drf�/p���4G�,&�n?-mȹ����e=��98[؂��@����f:�1��̅CJ�������QY{���\9zy��x�=OH�v.o9�8��-9�4|}ɀ7 �Yf��#��駺�n�S���ڌW`k�!EƘ�˟�z��p4���Gz1��N��+bb23PVܝ����#,�;�0:�ܩ=��_�t�.���s�Cz&��{��|��b�u��Ƨ�z�4�=�ޮǃo9��M�3Ѽ�������.|��#�%Mp�r��m��{�~��_f9�\�١kv��ݵ�l�p�'�铯y)+��ȗc5p��+s:���e���x,f�Vr������Ol����{R��ő�Np(n��U�q�Z�s�waq2��:a`�Qv�}3n��#��n�B�鸝̛��X;`  }doUw�G�q�1���>�f�N��R�:�]��	�#D{�T�m���È��IV��T���+(՞���d�Y�	{��{�_��>1�B�O��vC'o���
�p%�N���������ᄮ�ȃ~�Q@琭�����H�uқ�[!��g#�n=qp�5E�@l��ə0�	�+1�ˡ Q����:o$e��M�9R�U��N�,Я2�2���^[��H�6{���FGl�o���G�7�D[�s���gN�퉛��\�\9R�r�\�cy(�7��`��yF�ɣ|7P�v7=���,$�:QLLW":F�⏩�o�)YJ��0�������{�o6פzHq�r�%����ϊ��\V*4Y�/��|<~�jO�ƚ9+c`�+Gv��N#t�~�R�lv���XP��*�٪w.7j~γ��<���@�������sn����ﮋ��iJ����P��N	 �I��wN��9�z��w7�h���7G1�8s�$�����e�`�l�rvj4�=�^[�EK6���
�d}*'�v0���r�k�S�ӑ�3:�R�{jǣ�����{�6��%�a]ѻj Tk�v��̤*�1�|ci3s/�	���3�请OS�pםB��R=�.��Ȭ���+C���vmB"ةRsrg648Hܙ=��6�g{(M�B�ryk���������?�{n��VԿ�g�_�_�*7�ݔ@�=�4jgz
ߵF�W�]8��+��T��Ӟ�\?j�7�KC�E���o�b�&s�,{�܉G;������㥫'�	���	��ޮ�r
Co̎'���ƌ�]_%cC�@�~�x�^J<3�m���(ێi&�)����[�bZ��+LTt^SsG�.��WW�>�Z}c�>�Km�����"����ŗ�'(��T{޾q���#��6'k�K�蛑���A���X��ѱ�;2�^U�ӭ*������o����^6zy�Q{�gEG����Ğ�n3q�\��ECn}�D���$���)R��P9��@�1U��
==��#^ENNo�p�v���A�iWْ��>̹�"{kt��	&�őJ�2��!݊hC5E�赍ٛ�s�Ah�p�	�����¥�.eL.Ļ�#W��<v>]�8��Ŏf����v�v�.�{��ִj[-
U	3orH��U�t�Y���c�8���SLW-"��o~�D��<WA/�ml#� ?��79���Yq�r,}��	yo��toF��^���z[}�t*ầ&C\kl���PՔ�Ђv��}�BT�^X�Ǔ��0������/�=[X�
 V\���۶��X�H�뀢��0�|�+ǝP�-6{Pm.HGtj�����?O��"���T���
:���=79���Dh���,����,^Pݾ�f/�ʇJv�hc>�
������OT���]��;�b���:(V�VO�mA���dJ|J�u4��~�z��q�S,�^�`���o]�4T�L	�E��W�g�Tf�q�{x߮�/�:�f����K�ϴ@Ѳ����jf��o'b���?{/D���B�MV!�}x1���G��2��QU��X\��ʆ&s�oz�O໹B�0e��R�v'�?}�'�^\��o�����N�wk�Ay�a�J)���d���FLI����!"Ŧ!�������c~H�EeMf���WB�Șt<�ceN������='�;��C({!�]����Q{w��}X6e9L-��c.�Jy�����c���u(��?0^R1`�x�����9��X�#�nP�v|����y��'�����n��,����R]�y%��2;a^�]�̛t���wz<szί��N	�w�#NIa�[� �xʸ�fj������/VsN�[�����c7˔�j�sP��8��g�g8c�YS�'/}(pb����5�ԁ{I�9�r+茑$�������`'��!�"�"�w!D'n7��2����y2�m�����ގ����͌�h4s��ˈs&/j�>�}Q<$��a�ח$�14�2�(����d�54b�ǮkI�Y3���Vv�B�,�ԯ4$�v�:|��������J�c���lM�2�ĲvV��b�@m�x)�	��<������M�n^z�h�a�,��C��U���.r�z�/��J��^�F+.~��B�ȡր"�\ƼW�A�7�.���5�f1W{c����;��.����1�+%�P��*!�E�XyK�gI�`g���Id]_U����g	b�`�!z:K���h&G��fV�&p��J�8dXZ.'��N�Fu��g\�Q>����-����6��.�@�M�ꡳ���[f��/|X�5�`}���<�q��zo���}��q��n�Λ��3��E~�9Ƥ�����$��1ߥc���U��5���R-'F��TaYw'�D}�HÉ|� ��7��P�da����r)3�\�����=�v�w��8�;%\1����Ƿ�։ߥlgp3����������-�2�ah���C5��=ߣ��>���EUf-�Bzc�u��}Ex�h�S���}:8%������7��2>Pt���k*���䳶I����x�"��R��<�z�u�Z4,b%/A{�ް$��B�@"�Ͼ�c���Y42��&8ɒ�5�9��Q��`���
]�P���%&6�)�o�0ҕ
0ؿ�eWcX�O1�i��+�z��ֲ+X��ֈ�g�v���^����p�^����R�H��[Ң����聟mO�b�z;j�o1�w�:��u-^���A�F�\������Z[(w\�3��ǶφN�0�p����h��Ycھ.3��/�9�H��G���(n��YR�|pw`�7�R�1,/A��59��q�)r藒��I�W��~ �1]�$�1�����wov][��e���A���&4�Ŋ\�ݜ��������/�lǣ����ŁtxU7��<��q�R�ƹL�7Kh��N({�ԉ��^V3�W����fr�X����+�M̱[���M3�\Y���~b�(�G�E,tk�Qr��G�{Z#JxЋ=�/se���rѾ�G���� �����<�T�gK���DL�T�]HLV}�<=��ng+.7��8����,���u]�:�-�E�z#��:vX�xq	��Y'*g�+����;.0]>3��R�_X��H���N`���4�Fno�=����0�T����`򬑅�v=����=n(3�bށ�7n~G�_�y1f��d&��}.���k�Α��H�����w&#��G%����dPu�۵��.���VnF�32=5��Y�\A���E78W�ͬ�G��;j#���q�!��������f�F��`"N?Ew�3T�ɕ����c&��w��Q[bf�a�}�<�s�b�/8F��^1�^����ִ�{�{�e�w�Jf����|�Ih��b*�/]��J{.s�����_������ ����-��չs뒖�v���;hT���
b��y(����v����>'���dw��ίq*�$�ON�"��|L�U�b��T�0Øq�[tX:y^�U�Dd��텪.|2uGyG����9��hW{&"m:�M���O����;�o�;�fPm��}Q+�F�SH�y;����#-P}7����׆���]x�5��KZ:!�W���D�#��S�^"�+U����(�q<t�s�Z.[c��5&o0�ںV�U�M+�Tjg�<��%us��q޷f��M�a}��۩�j�辱�gN�{�﷽�\pA�2��;�f��M�\��n�b�lH�
]+:��Ũ+��4��:�w.蘍��=4z��b�ˤ�y�*^�;c=�ޱB�f�<�ƒ��/Ur� ]ګ�,qJXф�y4[�|�k�cO
^O��]���b�N�z*7�1ͦ����6����jPB�v�Rۅon�s���>�	�RK�:�)��4�Z�a؁1LNt�8s#���7)����Ұ�HCI!<�C��i:��HN'����B}�$�d��8�N5�i�e�u!�����?^$�o�uǩF�P"׻�ٴ8�=`H}��b��t�F��>�����[r���"��c$�garB��!�*�=kw���,P�̾���v�mYP����1�d�#�|�1_a#I�ڼfk��#��>E[�����ậ�:��!�R�[L���cR�$:����mS�i�D�8��o�y���dl����j�̐>a��{�����}���Pum����kU5)u_����~�{Ю��j�f��`i��b�o��=>Jz%�)�P�˧�+�γ׿sc�_xS����� 6��}��s�� m$"�XH{=^�7
���O�@�`I�$����[u�����r����i�IJ�ˏ��|�d'����gsS�#�ֹ��B�LI�o	7EH��0���3K��̅K��&ǩ3W�q�ݒx��w���$�6��}��+�˶Nj�.<x��Vg.5��YĜO����M3�s�������|�0�@�4�<��fP�B@�	 �fe�^O�x�2���an�4�TI.^�nP��hh��J<�inc�>ب�!}!]�}�w���B����a��[%��ȅ"��0�Q"g�Ʈ��ݿ���Z���t��U�y�0�*@�B�<I��(���p����C��2�ʗ(#l��H%�Feux�Ǚ����5�\͵�����=�{���A�/N������[Z��@�\y.Y�[�_N���
��TŞ�L��p�g�U���hZw\=W���9f.��ۏ#F,�\#湫rvW��;ˇx��ǁܹ���ެ>K0�#Nf��	��O����I�E%���ȧ����N1�2�}�;���������@���71:w�s�]� 
�d.3�9�=��5{��䑏�,5�<�xZm:"�J�̮�'���6��Փr��W������X��tgy�`���@=��N���S��8��p*�&)N�[�ޔ��6l�0{p�rg��j��}��$A��;�W�ĸ����9��=E<�C��%1��6�wM����ُ���ܺ�:�y���C��}z<��>ٻ�5ׇ�3�>'�[���%�[�A,�>��;*�3΋����z�t������[X��R� ����rʏR�FoQo_b9y��[���.|<���!Z�I0Cj��ۭFӻ��=/�SpV�%�I��-����=q᪗��/ٚv�Zr<n:ӕ�e�Z@o`��u*��yN�8�|.��1$X�m�\�,/:����D�c{��%�li�L��oAE��k.1��<�3ו�J}0Lưr1�i��js1v|��"�]w��YB��x�N�1o���`���|&��zT&�/�U��{wm����ʗ��["ZwR�8�ᜓ+D�X�c�W�M[�&u�D0\�^vr�;9J��ڳn\Ž ��c���fu�W�L���&P�	\	�P�>�	L����h��`�cޣ67�O��ͥ��*�r}�o2K>X�	�19{��Ld�)�!���L♜�&�ȋ?n^@�w�-��ڧ��t�^�E7�h��S�����x��H�'t�h�G�{҃^����s��:�o��O?K����)Ǖy^�D��Uf�ꆷG�Ϧj��j��B��E*�";��c1u5&�8��ɛ�x��R5_�qc<ۆ,��3�A�k\��GA'��ĭh˯Zj�/a 2���w�[E߾�u�p	����sG��0nW|>���,:�͙ڎ]hm�l�xϻ��>�>�3�5���+鮌A��II��ް�b��#�=�Y;]��q*�L-�a�XP����{�}>��'"�^��[�v/��|��l/.�{T.(z��3��xi2��L�$p9��|��b�e��v
�;�Ȟx@5Պ���b�<�Rq��h���`�U�9�qb��B�YR����+���]|�=�D�&Iq�6���B�X Zq�)7���=~ˎ�[�7	F����S�z��Þ�Vn/;b��)�(@u�o"�lN��i�d۽V:�@�w^�癩5;��AG��)ox���Kr���ƞ��d���bn���h`�a;ɑR4������8�`F�u^��p��)��~1�w��|NTe��sO��d��}C�/$΢�S[�̚u��m.C�����Qp����0�Nֿ/��t9ʞ��(�[Õ��FyQ���*p��
e�裡�Q6z��-q��P76���	��fm�ɾ1V��jaO7U{��6&LN<=��B�Y[����\�5h����x%Z��s����W�}ׄ��B��6�/��U�ǋ�� ��t���w[�b������:M]w]mM�k�R΂s�n�Z�L9h�r�7B��M5���!s�P�#ͳ�vo+�=s�����(x�J��p����t5�j��[�Q]ϼ��Y�5I{���t8�8�ٽ�8�_��������e���������P�����p��ZӞ��^���c�'Ut�vLE��j��g�(��.cĝ�Z${�)<�z�&U�2��~eG.��#����Υ�F��{j��\%���Z��N�l{�����u��!vW�{ޮ�fvY��q��4B����x��,:��ꪝ��{m[_m$�o��w���7�8�/�]�U�3g>{���Z"T�����u}��4v�j�M��t����֟�WZ+'�k7����g3��e��:�æ�u�Z�=tC	�*DDun�7�eX93_:l�ӄ}���������V8�<jɗ��UCv����(={/+��\�����m|)-�e׬�P�:�{[V�f�L�f���������#�	j�w�dj���Eأ �;��vk����VY����P�=��hO��.�����-����Ðz�G֓y�7)�%��Oią����X1�n'���g��
U	U@N�ŋ�9�^�v~1��\DD4�j�*�0Z��=p�gb�����������d,	�`��|n�c߲�gqt�� :�J|��ZH��V�˛���NTd�:t��~"���qT�vh�n�~"E��2��!�g%Q�0{��gN{�R�^|���ϳ�ז�%��i�4��}�Xc���<��yFrF���|��(��œ�M"�v��Qw壑(aU�r�:F��O%'L���&����]$Ny�(#�u;�:���yV�#pd�T�_Z�Z;�� �F�R�KbgՈn�2�%>P�4�j�Œ89�ڎ��5O��-ӳ�f<���˭�}C�|�]��1����Z�}N���cI�4�`�w��c5�p��3.[4i�#oo%��BT��d!�~��������58ΓL;�|���%7ޯ�a��J�/N�;;"��-:�8�;��թ�ʞeE�Ɯ!q��kW$��,�*��|у�oK푬�UA��.w�Jj+M�r� �!G��Lw�g���sjK���ɢ`�'��fc'ٶ�����$�s�c��$��GV�Ǉ�Rۮ�J�)�[�oD1���jQQ��F�a��yt�J�\2��]��|���=6{�X�\7el�����v'o1�����h(;%��+��ד�(/a�����WyF��x#���Q�]W�jJ=
a�5����Q��/H�Y��gEZ��<W�&�j��pwz�� ��I�ގ��c��:8F�����$��<�Ǡ�}|��3�u6֧�=����	��~�βb |fÈ�T4N$�d��Udq�Jh{o��w��^��P=Bo��"|6����TA�1�cM/�R�F<��D��X��f݌;���kb��E�<�ލӉ�_c�AQ���'�G��=à٩<z�^�5k%�p���y�:���
:��_5�����q;4s������9�~���/��'�����t{��|#��Z=��Y�"<������әtm�J�Y����$ 	 x#�I1��2���O)	ܱ�U֪�wW�ߵ����w�6{�H����?| =�M���:I���6����u=�2�2\��F�i�2r��՚��.��Q�˳�bRR��:�� r��F��]L��;_�=5!pFM�]Ҝp�����fP')/۹:�������quC��.��	��}{K��4\�p�藇ֳ��,-{�Z�r`��>^ج�.�_����H����z"�z�����U�ԣU��~�5�s��a '��������z���I��~̒!�5��sz\o^̣�����x m��{DY�jܲZ�s]��4��s�UdE޿'����!��Iԍ�{c�tt�GQ"Z�B�sqϻ2��o�+����`~W�L\U62x�&ѬP��c3��Y�Z�jJB��,�I.��Y��yH=���(n�j�F��Ji�������ٌ�	�4���0>��%z2�yuI�|ע��~5�K�j_gF�-UV�㳫L'�9z���-�m=�-I=�E*���Z�3�:#�t���uXhT����m#p��Hȯwt�ك���\>A֎��OFO�Ք}�W�P�y刣�ch����X����Y�f<��iƨ�-��Uu.���;�L\|��U%�f�%g���7�M�s��A�I�w��A�����j�gC�h��re�dpD�2�b91v���a�Ѷu�������_e�;��۹��#��xγ�l7�ӻ�s�	���7ӻ��l���� �[k=~����63��0�z��? ������1��X"�E�̕>�~�C��<u";�}���Ky��r�^��Q�T3�N\ԛ��I�ut���У탢�;ҝT�4���y+�рg�
�\f�vy��ԥ\���6����#I��
ܙ��'���}3SWB���}�Om="]�y;@��X��
���>�N���f����}�-������S�����v_���ߺ ��L��œ<�1\s�N-1�͡l�H왃��TБ��3٨���z�m�V����.�ȵ�n��N�C
7/��(�j�$O�z�G��D��w%]t]*��mI�U��<�ߴe�����Lj��@��y���uƸ�C�y(�����a/�ק�@�ᴑD�=�{�_�WF�uK( s�B�f�ډ��D�u��A��(Y��f:D]N��0}��=+rm��$�`��4?I�������zD,�kł�`^��{R��:{,�#��&G!�[�GE�����{�51�8��[��y�n�P��u��:�����*��8��t��fe���ؑ��deE�b��%k�y0����óg0�&�ܷ�W�U��Ύ�eF_JYKH�#�.����[�ɚ�q�J��� %wYz�p���c�jx�� a����Hb����F����713#N�\���r��}���]5ꨍ6}<q�Gb�{�^����&$��>�W!���ٲ8��8Y V�4j��Vzj���*��yn��z����+�f���{Jq�~�M�����P��@�|��nte����f2�O�5c׆t���n�ZyP��� ��[	X���l�|��}��n�Uê����"��<wr��[�y�3��#�b�K�6���uw>�l��-��y��ݽi*����צGdٶ��r�N��������f}�<�>��?W@W[0��٢��y"Ƿ��n��ގ���~'#���]���3�����%��>��2	�������u���2W���!��f�r�9覦g����F���C^�:�G��'����L���{�^���S���� kP~2+��G�nq#�y��dYR�YpN877;,��M��;A@�=owE7���I�*����E�Z��\ȮOY]t��1���Ǝ=���b�oNg��v���G���y�����:xY�GO,z�����w�D����G>q�����>�Z�2tlĦ�T�-���}�&v��?z&l�l2��(Wue�7���쀖�y./6�(U�K*b}ϝER�#��Q���:�;��7Ϳq���l
}�\�
�u������k�ܨ�=�`�1�����]L�B3|��αx�l�9���q�l����Nm��eh����h^>�\F2�K����`��\_��s��Ud�=3�4��{û�{g3�z�j�!W\?
�r�Ya���H�_,�u�K�FEO�e��G�������*�x��U�2���<�emB�Q�9������i������xu{����n��G�Q��@o�t�>�^0yg@K�0�-�����-=�嵑w谎���
RI��s�gU:�]�ߧmj�"O�w��]s�}Ox!�c$�Bi���ݺ�E���W�$C�SU�%�s�;�
xg9@M��"^��tmՍ�-c(�B���l�5�31g5� �"��u4�Dy��V���w*=�u��NHd�nv�F��ld�� �j��#�j�)��4���s�k�Z�0�B�=��e��f螖yѰ߸�B�*t��}&s.�ʖf�[~��[�=��s~�qp�7~��s���rw;�:���������w~��v�fzkM0�c�w[q�+�{OSn��ި>ˡ�P��WW�6t�;��Gz�z�o��"m>���a�؟���ki���%�C�ɢ��؆���紷��0Rz�F/�t0�vVLv��m��4=7g,+	��G��e��F���A^���	�x3j��8T���["�H�u��R�)��R�+�W�߁�k�v�Dg������Ob�z��I^U]����z��я�/=��
ٚtk
PMtȱ�����Ų��H��.r\9���������I�DW���1��u�u���Ũ�+�uv�3�<��vJ#��3�BU��.�:da��$=n�'ym7=P�2��h�3NAF��7�h+ȡ���2�����V����9�	�S{f
�v����T�t�?}��l5�}OW��e�\�`[[5��:�<���p̀u)���;{ں�r5u>fZ�
#��'n��4�bWc�1e	g#	��#�����ߗ��NĦƣP���{s���7*G�@Uo �qy��FX��՛���xښ�]�1���z}�Uϧ��J�8��U}�z��!m�[#n�,Ӷ���_L�E��(�]���ͻ���_v�MM+d�G-��8�x`8�>^��2j[�89ߪ�n�E	s��e�B*�~]�]{����rúvGwy��+�?P�[6�*�[�/ur|s�y��<��!���z���W�����mmv�u8��;U6�,�_���o\ul��Q��^EF$�����r���v�b�D�IJ&mwG�ETn{W�����<�zE���F�vj��O30շ���YO{Ό����wQ>�.��D���G}���� �������8��T̟�����g�)֕􎵾��/G����խ^ɻ)o�Y�mp&���_#�ܾ�����[P_,�T]]�넂�M�0D�s���>��\3����82���ǹ�G����u�`a��o-wys�Qzvn�S�w���'��q�+�4D7��l�'T�O���u>>�3��P�,�Dw1.�$.#rQhX�x���7;4�#���%2��(e\�t����Ouw �S$��g�W;�W��b�
��&�sKy]��HC"�&�Q����^�_ �a�������#h�xM3=szb�Nl�;�J뚗U2��k
Wi�@�	��́5ozx����W�I��oM�+18�4d}��	�|�I�O�Y�~O3��Y޲Cl:�M$�O��߻����A�3���sZ�JJR7L�+�ǎ�NcÁJ�Q*Fw��$�nVD���Mf~U�8q�:5�L�lk��H )�Ȩ`�!��sޯU��]{٠m��S8箽L�o�{6�ZKem�g�0Ry���016��4�e�Ti�js��6��*g0q7��n�O��r��V��^��i��y�l��{.�����䒤�!	w����ބR��d�<kV�ȳ;'>�+M�o�f�G��j�e-sa-�T�k=[N+W����}�b
z7OoZm�i�]���̨f�-E����9d�2�k/s���!��{������@8���o���Ƒ�柮�;��ˇ��X�N�f�g{�9Ȉ�����멢���g+[~�s�=0+sG�/���)Bh��A@@���x5�o�m�_T���4�P�D!�O��9���F���q泤�A?���"��ˎ)gr�b�Um�Q�֠�9c��P�(����|�ɀP`�C�=~<�d��m2)�#Q>�}����g^#N�W������s�q�V�3"72+f�q=~��j�����©9��C�'H�Q�c�,p���%�atK=/�eoN�T�.b��
=5	p���Nݰ��N-R�3��ǝ�ke�С�n�hN��\@��n��]P7�n��׻��Y�,M1JR�o�e��Qat\M]+ت}q�;~��y�1��t���Z�Ar�N�Ȼx��z]7��u�1Dr����ךw����d��s��\WuWHE���SWT6	t��<D�C�o�Xe\'+_]��NiZ�%Qq�����t';N�R�H6�)]�B��m���[B�--À&����fPy���u,�J]�/W]�;�R���ք���ۧ0R��8�����n�	ZFX1���;nP�:�J%�q����x{̇�_{�	��eΧs�t�R�t�c�5�s6�>ksXv�m|:�F�	нü �}W���=>gwd�i����z�����V6�N�l!:+�ajن�goMLe��G:��!k�c6�,{x����E�ִ��v�{���X;���9[jm4������'vvTi�*p�we����{`ٝG-�9�:4�%���C����<����L$�/�������U:���Z��>��iv��)եw
�w�l�6\�m�.�i�e=y�	�-�W�37�}��;p�V�}Ϟ�
=޲&���8翪�ޯV5���߈I�w��}��29jW-x��|ԹC�\}��K}0>������ޥގW��ח�/NmI/��>���	�.�}��`Z���*z�lq���bP�r��8u9?v�=�c1r��y<5��E�o�\tU�<�x����*��~���_�&��%�7:M�>��.J�+>#9aI��UU�,�\(�:�bx�9�P�ó� ~�~�$��#}���_���7��Ǹ�}]=�>U�Cab�ъ��W�O���J|��I��� ����wwFɌ�ޛ���_���Q=����7��ý"��䒅hVo��1��\�3s3�-�9B�^���5�3�ʩ��tOr��gR�&2��?g59���la��"���gH�
�=	h��Qp��=u��3s�+¶{ƃޛ��+lx��{uwPu�F���\#�/��!
H4^��ӆzI�^->��U�;����}>��lB�B�Js�!%�, �܌�x��oHѷu��P��u>�������\�q\�ݝ87�o�m{N�g%�㬿{��8���Ɉ��.Z�����D��K�?s�������2Ɛrg`�lcݤ�bX����IK�X����J|k9�/��k�5M��)��h)���fv����]{�O1�܊ك=��w����{�3��;`z���o��tYh�&�Xlˬ��R=��^��5=2�GoI�H�c�M�[�m}F�+�h�1zҋ�fh�nI��	(F���(�����v����Z�ϪoqT�����u��N��_���1Ӗ��Ű�U���Q���i��Ug�q�A~ |.z,�[��}8�����:({��A����3:����~Γ^�*��i\\.7��[�Uv�|E�j^�u}�����ή��^��n��]T^��`���[�V�bz���J�S.o1��<-"�
|yP�/r�����3����Լp�w �| �>����o���ل�">�Ybϒ{E�K"�˛ބ
y�G�y{qJ~<�b)Qѧ�&;}pW�F���=[:�tR:�-�蓛��oV��?M��UJa��g.�:�lNܑ����ɠ�˄^
w^{��Ю�\0b�Ǌ��4���^x��}���e]7V�*�����ً�����6�N��˨��α�Lz.s�|�"n���3�f|�����5z��~�o۵���&70m"�u1M�O�;�nQN��R[�jcﾎ>��u}��[���Q�j"�d�s,����D��f�>�k�J�C��0�;�>�|%*��e՗�څ�K�A���g�/�j�NX��Z�*�W�+�z�W`��;�>�%׮������W��;��p�݉���ڛ��=���#�sy�-e̗��ݾ���սLua;�~�}%a�����8�H���3HV]���L*̵�ޥ��ͽrDQ��[sލ��PՂ=c��̼��gVw��Iѯ�}3�c��OW����x/N���%NgJԃc�"�`�Q�*��Ի�����{X��vĂ��f=��k�ʡ��~�h��G#�[�v���,/F��>D-�= �%�(����g�a�~��6Ϟ��N���,�=;z�]�\����k��w��0>c`�H�|������4��m��{�}W�_ 4r�Y� ��Ǜ��ʱ]�-�BCQՒ�us1��խ���-.���{4�q���fxݼ�Uv��ӳ(v�Y�_�b#t�R�ӝ�\������zB�%m��Wj��+M�
��:���w_a5�td�������d��d�;�JVI�������W�̑Rg�q�� ����@bc��Խk\�Ϧ�Gb�׿S��y�8.gVftdhǩ�qt::V�MM]	+ɨ1"Rɪ{��{/o��z�:�����"'B&=�����<2�<�|�9q�Ό�>��w3�o{��I��@��UFR�7^i�T�N%�ח��e�1S���]J�� ������׃0vvZ���^d��,e�s^Qu�AO�eM�}���ޟ�ws�~�̬E59wv�ΐ�g�ʐ>��P32�[¯Q΃��a{�p��:+�&��&���5�>C��5r�>M��ԏFK�
F����{���I��7�h�=���ĉ�'�ፎo�,�p����=0s[Z�w@.1�>����ҨI����wy��7I���^�B){�rk�B���vA����ajiVm��M����b�-J�c�H���,�o��\Υ�Vt�k�c��-m-��Y0I�?���S_V�Gi�~��+mʸ��R�w������K�nҿޫ���^�5���݉��޿��+s;�`��P
�W���J���Wx�����|Mϫط�����r�{/"�dר�v�g�¥������G_]��_r&{���
����Y�9�u�6��4��^t#�B�Џ��������5J�l� �����ݗ]���l�ѕ��oTҍg"fP��%��M?��L6k�܋��!�X�������{>��;Uǫ�R�֟�<���RY�#��:�l:��/
K���+�5?n��U~V1VԳLz�Tq����Y�k�dϚ�}�1ۑ5�K O�x�ә�b��]	^ɞ����LrsZ*����&�X��r'������*K4ڇu~2���L�o��s�533�x�J��N+�vo���'x��w��s}���؍���U�E���������!Yb�z�	��4_>��3޻�Zk��u~(���$�N޻��(M���{�'���`,x{]�S(c���d��
î.o���!��Mj��hӷ�[{u�˲�b���:�YY#����)�w�;��\ׯȻ�웡��GY��?r�&,��n��Ƈ�:��.���O>����ym�ξ�K�� �}�FQ���іߣ:#;uN���x�n�/\�g0��n��J%3&��GD�{6�;��Z��{��z���Q������ �S/�N��snI���g�����Hl��N� |7�7uR���n��#���*Ӄ�gc��x{�dXc�C6�_`P�������I��ї=O3�y�K���v{]R�+hu�O�F�s��&{�JL��`����}�b�z�a��%0��]�`�<�ӻ�.��WVL*�u��˼vwb�(��}����~�(d��E�l ��"�5��`��=vd�ؾ��ؘ�<��㪠��ϼ�������6Sqh�߄�":T���	���W��ou���c��<]�W��axo�f��ڮ+N�g9�b4)-˩��l��� �hQQc���T��/9_	SZ٩�ǭoK�_f�c��hf_I����).i1��b�f��`�?�����?/>��f�'P���.��k��;d�Ƥ#��Rw(H�3wA����hz.;��)�����*��ϹuUL�֍���~�a�A���;�����٧-����دyW��+^���\�6�s�;�`����/ǽ9pM�^ߧ�}f��IHչ.c�g�E׏Z����5&O^gE�o�ewf���S��\n��\��4�8���D��Tf�}�N�뎮�=�ef���W�5�HŞ����O���쪬n�e������i��� 2PC�3������W�eƫ�#����+(C�}Y�����>��Y�V(.��鸋ˤD��ӞW+d������#}Z<��ލ��Q�#�O,�rC����^S��)8��]^�Y^~
���n0����~�S%֯pj���NR�X��	MT�_�����џVھ4l�w	iq��I_��Uۤ�xcI��{�����C��*���d5�t�׽v����k��`����sU�2�F��n���D'E����2�]{v��]!��N��NrR���W����7K�5��'I�^G���+"B����s��l�q�.��/��g�Ha��`&TI�yݙ�ٺ����V-�>����;gޱ�J_���L�Y6�*��ʩ�7q�2s���N��W8^��6k&�j��󡢜ʐtl��+�����F�C��ɬ��W�r��^.�5���;���x��@v-���q�}˲���ͪ����/XQ��ޅ�9ڐ�̟�-"@��!��2��g���жu����Q�-��k_e�C�0��VJk�U���s-,���u�OyG9X��I��#G�"h���|�����"q�W7�lX�&}޿������ovw�y��E!�z^�����~3�j� �1�+ŉ�"s!!���ؿ]?�,z���޽�� =�I���r��\ǹX�O��G?9{�}�a���Rx g[��KeI�$�x.��҇.�����N�FU�l�H9N��B󤒎<��u�9�q��_v>��`�Ja�����.�j����g'A�97��3/�Ι��c�Xp���������L��b���קN)r��틹�ps^Ɯ���ÀٌS���]�z�:ʠ}s�[�\v��먊٨��)�qY/_�1W����-ڲ3c�}�§��g���`��j�<��U�<O>Z�O����1�E�^O^z�=9��~S_��zU}R�����+�4���t��h�����ϙ޾�9ha�K$&�A����9IF�W�O}�^�q��sӹ�X���y5X��m^�����3+Eɣ�j��x�I�t׳���>=�LMuwc��V�LY�*'���W��
�.c��w����"�~�;�z�i䃮��M*b�>��L�
�ʀ�w>�^��+*�1�Ԏ�i�����g�R�d\�.[U�!>7����^(�B�y���uz�^O�d͂b�ǽ^zj�����e�=G>ȝ����w��M��s�^���m�{�t�,>��;� U�ln��z��,���������m8��ȵ�`��9�����GwXQ^�n��8����	j^�n]�vp��v}��=���A��?9���Op0�^aY��+��T%T�Υ�N��Ej�M�Ď��y��~�X�p0�YFg./���z����u�3���5��Ց�&�Z�f������ʏ<��t��T3;]�{;�tP�����\�r�]�,ExeҸ�~>ʵ����f�f�{����� S�����F�U�m�H�ՙb-��7�'��ٍW]�����[r�LX��NF��Y����"��[4:_mV�80��S�(=�t���	��np����;q2��X�Gg�։����g��K�{���!�g��D"/��*�@�U³�v��v�㻙~eN�7���/!^\#����s5U�(^f5�Q}�3O>�[06����G=��Y���R�ݶ49��Sg뱷�]��9Mt�ݔ�;hxOW/����-	�ᔤ`Cw%w�wާ*z�`��9���j:���+�>�̝�L�,Z5����H��X�q������G��NB�}�7�����k��/�qFD��o2ӆM��t�y����O�9�s̊`^�%	�E�Gj�G9�KZ�Q���9YG��'�ТwR8k�f�����w��:�j��)�
u��@�6�>��M����m�}=)Ը6ld_0{���U���Of0�me<�[���R�U��0��Ƭ��;�޶�S��{Vx�Z�}�j!B�g����`.	�і׆3�MbT��A(��I�ʟ� dJJK�
�f��s�E�F�CC�7s�u��᧡��;W�#��cIz4��{�.�Y�u�1�U�c�,��v����+��]�����:�Z��:��W}��q�z��c.�r=�ĩ��X����o){��Π���GVt���O$�r�a���37��tms�}:t�}%�՛����1%:igO{���4�}�2_���]U���;��O�өD����čH3�uJ��Ġ��TY/��Ӳr�t��[}����;�/p8���e�_3�fB��sy�W	�uK���fə!��$y��w�3�ф�a�HnS��f�i��r��Lşb��/�@AlGJY�A3��*S�=�w��y3���~O�����k�Hvݠ��"!G��xK��,��
m�n^å}�Dޢ�x��MF5\Ǥ�b��$:�n��aH�a���wt��f�Z�.�?�mA? 5�Y'�Zʚt�9rlq��Z�(��7�-�E�0��{�v�|zh����x=����6�SΛ&�^~�é�bu��n����y�e�-c��GX��ܾ�+��m���sf�N�s�z4wy�֯Ovqb��C�{���ջ�W���N��)v�v�Z�$�4T'�����sԞ_���)����۩�t��ÝK�����Fv��kSD�A�/y��#��������2��D�52v}>���]_%&P�%}�1�Cv:�gh��:�x����x�|s��Zf6
�?��F��}��S>̃=�*ӹ�9؉g<�y��e�w�wv"k�D
�nZ�O=��6[0f�ubN��į?e�ۭtz��DtK�����~U8n��&���̴�^;���xj��&�:sS�A�]��ݝ��Xԝ�RL�)���c�{�12H[ЖL���z�Z���\��Mph|�s�]�`��3����m�vD�[e�K��<ڄ�ڞ!ݾ{��K�,#X\��]&���F����zS���u
#�y�c鳳Ԯ��J���p3��n,���$3;0���S,�l.��3q�}�K�r+
�,�ӻy��70Q�u�~�!>�̓�bG[+3c��S߯$�9����`�b���k/.�>�m�yȮ�;DT\ޭ52ڥ�"�y�0�Dvأ��y5���z�"�N;�c��ri�%Fo��h����&�wø�*^�m�wY��UU^���T�{i�NSV	V<2�J��ٺ{�j��o&��H �����[���r͆�'���x��<��v�0n�,L�7�hiG�U6����=�U~Z����\s�;�:q��ꞷ.��R����D����U<�H����;����w�9V&*lH�ԗ�ȓ^�$u�cu����y�=�;҆�8��.���a��B�k'2���9��ɭ����H����W��EUdH�щ(�|>����;��P/���sU�:M�@��#jӿT-�U��M��d��ƥ��,=A�߆��Z����l�j��*�m�z0�۫i�pu�P�nN�F��Gz.�G��{�9�'"����
���3�r�2/Eg*٤�̣X3�Eߡm��r8m�Åof@϶1�V���U\f1E1>��eyC�rc������IZ%΅�^�ʍ�xMj4�9q�K�s�ѽ�i��p�{��p��w$А��ѡ���[u��C��+����<>�)"q�C��ky�xF���LSw���:�hH�qEO՚��X�7�5��뤻�:�T�9�r�H۴�pY�*�]Q�6㽜w�wP�m��QшJwX�����dfO�ԭt�J]'6�~��v}��ۓ�"����**��2눜��Ο��M�#�{�]f��1Y_�X�7*�UL�q�sφeq���n_T��&�37�)s�Q�7Hp�� ��All9�b��	X}�;�ɋ�:�]�9kA�ӻД߳m�&|�Tw�f�=�C����t�x^�����^/H=�f2}�=��\CHW�$ż�����k��~Os�#����`�eX|�{�&�W--T�L\?F  >��uq��{�d_ٝ-������m���[�7[_}�T��%��*S��(��=����t8��u������j�3e�p3Vj��&�UǇg����z���B�W�'Nk��r��U�t�܋k�dJ�Gc�5^�zg:��,�]�]wf�H�ݿ֖uE�᳼��}ju�{��g�MUZ9����e3�>h���E.fr��|^=����j-/���!��ĢHQ�$*�
,���q�o}�����p�d��6�2��=���'b�ɓ��l�$.N��$8K'�7��0f^�J�&e�K��6��n�Sw T��V?-�'�_>}�o� ���Q��y �]�D0+�ϯݗu�ǰ��H���N�eǷ�{~�9������a�����G.l��\�v{1��O`^x>�
U�u�߽�/��l�#ƳSUSW9r�o1}7s��/�[�z360<�|�*7z5q(��Y�O�v���g�����{q����[SR��ϒiX"�˙�ۓ�o|�ϝ:I<�Iz����"�^��(�Jw���n�\[����|͋��d�bP�Ig�|���Ώv��9z�M/(����~Ȱ�}���G�E\$0��U�#ۢj8�(�w�U/�w
~"�d^f�j1,\�j����~���{���]zb{��뾢�z�+�U��E`p�)�z�{F�Tw;-,����f���S�M�޹��J�+�?.��������fQr��b|�r�M]y{و#�E�	tS�yc�_�N�ɱ1�C:�cN�.m�fKwu�i��fV�i�����,v���=�{���~x�]���s������]��l����6�u��o�w�𚖳�Y\��+��x88'����Wx=<gj
�)�u{[=Z�]�r$�W�,���A�r��~E��y�=P;:��렪��w��ݺ�\��W"�͚�6�At�'Y+r�gجp��d�A���۽���D���lN��6G��@f��/Et�z�Z�Ό�Gr̮��ߘ��Vm����t܋Y	�A��w/-���{��"��O�Gz�؎�jX�Ep��E����Wa�T�i�#���s���=��r=W�K���Q7ְ����kD���Wu��T��~�edxOvzq>������8� ڱ�bal;-?S���V=�FwT��j�r�/�9Ǹyp��uQV�񊘩N�v�p*g1�R���X�ƾ������M��Μ�=9"}����:<��ٔ�we������B�>Z^��Vg�G�*:����M癣�2.�tN���3+{���������!X@��L�^�{e�N�i�$�`���ɻ��V�z��si׼O���!�Ow���.
r�vB޿�s����0T����נ+.F�
8d2(Y�n�VƟX�wR��b2ԟ�<��f��Tl��i��jd��T9�4���~�FAE�d���_��w^�ݝ��1�a���e�
7��m���{�/e��瞋q�6�]���	x*� �Rv۟��s�wU�ܯϱ5�����9^�/&3���v1^�������C�]Z`WJ�Ϳvzw��[����z	�9�g��57=?+1�T�70E���@ ��:��}d��@�v6(n'՘5����ΖՕj�ol{k�rs�ou�����߾�1��_��6
�m�fad띬�n��ۛ��97�k��v��2+�hA�^�{%Ә��wQ]���|z������{RQ�!�y�ݔ���g�j�O�ʵ����n�u�n���.�,����xz#]H�ZW�^����[�a�L[��-]ݏK��륦JkC3إ�jYB�'8��7Z��7�@��o���*[��gd��&��N�����vć�-	X���݈{�9rRO'K����ʧ�z_Wg*��Q��:mf��"7v̤!�4�YRm���
f��[^�ƣ����cR1�j����m���W����>��F���}�����#���`L9���K�U*n����ݟX3�ʪs���@�oO���}\:���_�,����$���ǴVG�s��|��Ѭ��ǳrez���v<w��6�����v�5w�C��w�����k��gxVۭQ�����GXڬ��]�Ҷ$��$�ݓw�
�\�)����s�Y�V�bZ�{�=��
ns��QIy�����G��v{��PO�Uک�(��mW�e��8�o� gy��	�u�\���@~���>SU��-���A�O4�no\��M,Y��Պ��==�g�DJ��w巷R�^�t���t՚F:�k=}����:�5;79��U�;�c�k�g��T�L�z�	�p�{�/O�R���ݚυ�S�n>�=�\�{�q�ݺ|L�Ln۟;L_�ڛB����߮�󣣮���	�0�y������I��� �Ŕ����ޛ9zNԧ^9�g��69{���?t�G}�漢��`�D��9&,�k_0��OG���T���]�����t֕�[��k��Lt�mK�uz�,�����Qy��[�#�t�"9Z�}�u9�z�6�ëS���z�ZW���lU�ȭ ��^�+�����ϊ�n�P�w_Xq�=w�WǞn�Wv�����s�s��/fM�W����YVr�9S������Bt�y��z~v,����go�ƨ��3�h|�Q���5`�m����KܓgI�:{4gz6z��E'0�Yo��7�{�����:J�F���ΰ0��yԼc=�;sG	���.Hν�V�R3���JTNa���� ������M��/�gr�y���z���'j��1��p_�m��}^�w�WG�g̢N�:̓.�#�Ut�^pZȟG�}�������=��)ٓ畊$ipԝ��\�T�VEIj�VUe�6��֞QOˈp����gb�F��y�0ɗ)Ů��
��o,��}�ƕ��t�f��y���Q[X��џlJF�v>�!rT7�e�ŷ���8��(WV�_h}lF�(�Y�W���� `f��nh��j3	>��A�D�\�k�^5�k���K]A��˳�cO�^��έ����)�/���(M�����:��wO]1�y`̾ζ�.�����:���@n�~��a�Gb�Y��p��l�oy8noP��>����uy`ن�MP�p��-�+;�ڪK��ć_�0ڟG�*�w��j�}��|ʺEm�2)��=v#���1�~:�ס�k�{qX=W�;q�?mz*��N�I�ow��-�V�9��?;�J��g�Y~g�I��IP̋,ȃ�.�n�Y�c��Ui�Old�f�s+�����^={lz6���n�20�A�y���;�1d�w'o�e�}F���-�F ��X�Ew���O��ْ�f^I�O(ܱ���SAb�L����n�J(#� ��O�׷2��D`����|Ƅ���W*i�<׳�����W���L�[�cӊ�r�`�~PTT���浚�Zֽ�������}�rU�:&�5���c���d��&�=ד�s	��=빊�l�C(7�{��mG�8!��K�-�_-�r��y�[���zRu��G�i���1�5���_8���>��>�����r�ޅ�P&8����1F�������f�������=>|�ai�A�G%o�l(=�0�+��l�U���eK�gNµ���#��FТW�����3���fw�h� �}�V���=�;f0Ï_tUev(��9��S�.K�y3~ocQ��P���^T�򺟧��ZlQ�y/�r��p*y�a�%ѝQ�[qy4_�E�ݮ�yX 
4����i�mI����!pc����1J۪����2�)dsy��*�;�
"�f��v��������g�_m���f�h���,���Ic�YB�]����9ُ^Թ}}'Ċ�wp,<�a\z-�KhoMEf9؜9�ϒ���0����M|��O:{��t��5v�s_����s������Ȣ� ����Q����5��k��{]����=�Ο�ggy�;~�E"��**�Ĭ#i����{����ٹ4���Λ�ޔ��6�n�|��)g�3H����}��q����.��ga�>Z}ÆXj��Zu�Ӌ(��w�����<��7n���6,�t�vŶIgo�.*kKb|n���'zr��ܹ�R�oN����z� �+ddU��f�dgݓ�"��n�Ǥ��I��;U+b�S�S�H��n��4���������ݦ:}Q��+�W�%F��/�<��+ }���z���N��?p���tX1lt�ɰ{�^��صQ>��<��U����X��Yb5߳��=�;�mn���1��ΪV�s@iu�u����+蕤�-��u����:�y��^G5D�7�o �q����E�]���׮�x+G��u���R���>���%O`��W�� /�:��k�[:/&�ONu۰oCבm[��U���QYˮ�Sw�K*q�S1s�3������t_g�׹���G?l�q�پ7������"<����z��	��ɯV��g?��dx���=jٔ�u�T<3��"S���h�d?c^U<��8f�~��TA4^q�js�<	\�MRY�\��6�Aiw��z��NK98���x�Zm� ����=���^>�xҺ�7�]��sv���л�85��ހsI�֖U��փZ[�Mܖy��7����x�^}�Y�{j�ܓB���]��`l,v���B�g�!~=E~�r���Z��8��v�;ׇ=? ֞�������#@?��6� L!rtϘE�D&�L0�+�hB�ɿ�!��ע� q����xJڽ�D� NZ͠�q�qӛǲt]6fݼ��aI÷#erμ���/w%�%���:�[�c*ޜ<�<r@z� ^��p��S�V፹��wFc��z����
�J�QU�Y>�vH:it=}��l��\Z��/imp�������j	���ZZ���&&�-ay�����,b91��18�Q�]���e�"6�����+�AY\K)�W���Op���c�7����u#z�dZ:68p/j�-6�C]�����m&�*�t���3z�L�����hmL��w9&�Z|{�����5�5�u��KQ��d@�O�)utEj'bFS���͉I�a'�I,���Q���Ir�}��JH�+;�ǌ����/]�d�E%޼�_W��~�Sm՗٬{�c7{�-A��eh��AJ�3�)E���S'��ތ��˽9��^޷��y�=�]2��놵�Y�bϭyK��m����u]�g���һ0�vȩ�n@u
�q^+/$��N���gU�<�Gh�~�"�X��
w|oa�*�_n���7�H�󶟏I;ݛ떦�o[����8fr������Ft���u������w�vf�ͬTJwD��7A�D.E�(���:O���5\��0Y��<&w�N�����ө���o^Qb�s�:��Ŕ����:鴢h$�O�{%+k�Y$�&�KXm"���x/�2e�5�̿!b0(�ͭB�:hhdk��j6R*�&It4����"���R�x�ڃ�"�<�����"	�&����y��lǽ%e�`�{����k��&ۋ;Of�\s�[b�%���w���K���y_Kr������du-w�enqi|7cõ�R$�H�u%*닭:s�>{{}�>�JWz�Nj���Q�ךv�e��F��<�|�X�׻�q�L���T�Fg[�zE�כ� �h��|S�:�}�:=���f^��ُ]�kC�<��[��.�o���a���s��҃��^�rڵ�bmz�<�x���ކ2�ʂ^D���kG
�!>4L�;���
���_F!ˁ�8n���r^��]ٸe��q����gsm�ɵLY���q�фk��uӁ9�޷܁�Qm����d���]}�%^���=�}�,��A��fZ�/n_5��9V⛕2����Wc2��W�UUE��Γ�p����m��)��[�ɏ��,���j�1���v�pŁ���U�S�wW/d�o`㷂��0gG���O���g��4r�{o(���U�C^�%��l�m�)��NU�����V������~�l��Z�����+�⿿l�=b�×���0�-�Cs�"�����ڀDDk>:��1��5z ͚��g�/��� ��.qn�<˫�ͮ����uO?%FU%��v�H�ȸ�/JF��V��;�OF�^�p��S��}�#��Z�^Wd���.&��g�`�� S������9^�+p���yE�d�?y�`#��i S���K��\<��#�E��'\��e��D��/oג��:�����+��f^���Vߘ�~iض�����W�U���]��W{Y�X����]�C�n~����A���s ����	?|'e��(?G�N��B�Q+�ڌ���C���To�D���RX��eg���i�Kt�-�-t({�p)���zF�weU!���+�T�Gt�aR6[�V�8�Ub-�`���Aa����j�C��Q���Y�,�}�r�z\;�8dW]]Qf�s��ۓz,rl���wn5�FՖ�;br������o��%v�Y{2!���e'�VN�u�����W��Xʞ�����)=:vj��;��?-���]�wf�����{#��]yl�\9ˣg��'3C������������ |{:k���� ��*�i�,|�Wu����y��/Щ-��m�{Nv{ñ��y`�{ !*TԪ�v���b��-��S�g���k�=ۚ�\k؀����it9����V��l��l�QO;���{{�r�]zB��Lw_��9=3��Q;�k���G�GK�Fpӧw��&���\c�f��hA���Q�T=�xɂp"x��Oz�dU�&��F���N�U172"tF�q�-s��x��>^��������vZ:�jz+k."�r1�����c�?)�4�5T��͜Hj�f`�G�F�!Bef}Kl���w~�����C� v�yr��pHߗ�c2Ń�/^�o�M֤��i5Q��._�G��Hn3s��#WgX�l0���'U�|V��왳:5��9pk���g�4*e��|���U���I��P��k��X���1�e�<��v�C&���<;���c��3ޖ\P`:�3{��b�f0���H�;Tr=�#!C�R�������X�*���b�w��ڿh5)E����9��JJz��2�y0e!�3��+W�	2�@�!�;,�驁J�P���]vS<�{c�YO&���R��Q�bо�Ф�����M�
�֦Zp��*�ɧu��n��q0G)���G�B�N������ᕎQ�o/���֢���7!a^�
#�==��d��+)/��k�s�s��M}�Q���2)��v��2/D���⅝�|+��`�Gw�K+9���m�����uWPh��m��z�} �ŗ�HK���`�eK;�Q�7�$�M���U�N���a�zB>�6�L�j�q��Iw�yu��!=N���t@I��< ,�W�gb�>R����fa�T_+st�ֻ�z�(�
��1�\�iٚ���
7q�2��.�����"bos���7���ww/��vr�^[���1;]˻�\Y��ty��EA���ʈ2��0�=ޑ7{_�k4t��o��0�e'<�*e��<OĐ��j-j�V�]Ks��E�(F4�x�ff#jX��8�ٛ�&��⋧nn��6��S-ӍR��ˎ��E�ٝl�;F�1OZwRf3�֙���C̸��^tݜ�nTX���J���@�ez�>DTr��2RNV:
io��n H����eʏt��D���a�+}yr퉻�"�����0��������̣i�:I���.3vrDnF��J�B�9�1�8Z���F��~=(țq�_V�.���N�0���m`[����nY�P�A�o�tØ�F���TdY���鷧�����L
�����ʫ'�k��+Z7���	O��}��j����=��	�Kf ��'����='AL��N��n�6����u�����j+�(��܅�2I��X�%gr��w�j�\>�Q���ɧu-�l�ϓ���[Ǹ1��;iwdxТ��z-�����ِE��d�=☃�D���|�ʭ��f8���;>Aл�U�\o*����C}1}���Q��
',A �o�����Co&3~�P��),��K^�n��?iV� ��J����D�&;Yc=G�N�v���P&NNK�P����� ���5Z��G��\�%�����Nꃱʺ�&� �t���q9���Ӡ)�5��LX�;����*��HXd�W���L�a�*��Z{z���W��4W`Z|��u��l!��N¬[$TǱ�"V���GD'3S�	H�>Gx1�
������$�n�I����=�԰Q�{u5Y~��T~8	8�wQӥ�>�Os���6�\c�!WQ>��;�bѤ7{`m�dSw�t��D{��o�=� ?}��>�t=�Dq��{�ՠ��Ub��誶�yL�nV47=�c��l>][d��{_���z{�"ρ���߯�'�遛�br,ȸ�#��ٹɋ��c^�47��9p������P�~z�Xi�E�Ԯ��Q�3uGt�4���8|�O�`��L�rat%�]�4����L5�3�\�A�{L3[�[Z���ߍU"	c�{��R~Y�;��cև�&���US�Nn�Aa��{�`�D�J�Wi b�T� ʄ�\�R�]O��N�R|��}qT�u^{����I��Dl��u���3�v��ɦu{��t;�;`�x�o�SbN���puE�ЄՈ�5�y]�����.c�g�q�F"��FE�o����H���q���w'��L hW���l�r�b�x�`Ѯ�|���D9敞V3M���I���#��<0��]9��2�ӻ�#�e�������(r��U=������)�靝4������/�z�o;�WRTᓕ�8=5m�y����`�+u��=���Q&.O�������X_�3]�c��36X�ri,؟d%��Ab���1�D���l���r���p��D'�fHYnE��LF��~=��X��"���9 M�]�w#��#��Dj�2�T�Y"qM�吴�a����0<��������M�v,�чB�6~>�=l�sn�9�ճ>f`+�q�e-ubjF��O�ݾ �ԋ��(S=�}jzs�S��U�[��`}�#S��=0nH5��?��нl�\�	��8���vH�O!V+ʔ����)��=c0t��Bfށ��d�?�ȿ�����y�s,�dmp��6�����ճӱ�9u��؅CA��ұ�n�?G��+�rn�!�r#�fG"�w=�E�(o�P1Pm��8���Pu�>��E��������:a��i�a��Ey�W��ѱB����o�r}�d7ƽ.�=�$��� ��QƎ��v�w��*�^<Ʌ{]R=����;�w�q���S��N�V�{��6��۹b�X��znm3� :6^���3��f�uK�U�w�.w�I͂����|�Y7��NTw��]X�x�g1�H̩m��{)$�x^j�O��zj��Ց>���s1�<��h�4}�����|p�z��ǜ7���/)��� ͛�|���l5Ѳ	�'�k،�{l����rL��L�:������&����Jeտ���������<��כ$�����~��8�vQ6�>s
�/LX����t�W=�;�"����j����&u��e��¡PjnϴF0��"��؇/p���Z��2pV����TY'�kg���o�ϵ�&���h3��{�
^�)n^�	֚��;t��3>@ʓ�[�mm������r���xd�_F��huGUn]4#'g&^W�F3��sn�>��=y�v�A�aԓ��"�F������Fc>ʌv�FG��>��aE�HZ�yy���P��=e^�oԄl<ʟf�%����֑����}�p��o�~ᣌ�'y*�_	J��Yo���':6I�=�1�İ�a�]�8��.�y4�*���rLH�]�j�/z��7W��+����8/vL�?Qq$���Dtu�8�@��D� ����n�v���q����:�#�ɫ�g8��^sl�Y�7�,�o��gZ���U�Lۨ��[����♲�3K������������R f6�o�@��9_ַ���i�N����&M�>�ۆ�më�<	kB=G�i(���̓q�kAZ�_U�^w��v�A@;hU�[��Foj�x�`q��p� ��܋�T)�_)�P�L��2�ˀV�h�O�+xus�W4�Z�(�UA�.7�9���fOi�PX�s���|�����q��F�v���*5����л�|oq+�b��;�o���֬.u$�r��'��=�v"��^���T:	�����{�����*%� �11�� ��@G
=ͯK�+=bV���~�~�U�p�A�ulzb��,�����"�#��.�t)5S�#������: z� :3�����������*�����a�����^%tËz4�WzOy�T��7�(�11��قk�2�,��뫪T�,�z�A������8	�m��ҾCO�::����/�,��*�{�Y����z�\N��_oi���|>Aޤ�r�����Ya�}��*Hl�N�����Fy�*TQc�WkVꮐ�%uHiYW�q]5Yx�ر,��S\B�u0�g%IZ��A�e��Wr����av��]V����.����K�f���7����<�0���Qi�m`=�N�ŁW9�D�dذ�`	>��yc�<�h�g�+b�4����ʐ�d0pv��'e���,t�+7"���;���^9�#��~��gmSG��~��G�H2�F��GNivd�d7�	[�)D�EN;{WU�<��oW���Ԝ�p�*��:Q�k���>�bN��ຖa��8	K�D[�qI�K���g Q��Whprjk8�%�ϡ�df-��\d �~��yѵ�m�\�-Lt�u5�K�Ƭ�H���\K������W�q+�@�6[���<�+�q]�إ^]��~����mLC�qO�:�z��81���N�����u%&Eu�00G��M�d_/��#��=UAM���P��S���.,Y�XGK�"ȯ���lp�jdRry�asB&��A�~k�@a� �"�c-�ȱo:���2w��ع�'c&�n&Z��d��W+�����F�0D��Yi'��kƍ��x���C6"���ȐS�I��ڜ6<�bf�mn>�U�<�6G8X���.�Yx�ܕ��'�g~�>$
~���
�g��{�Vnڥ��F�W�H�2\� �Qe�s�5�\�����w]jԞ�ʴgS2vNR�3̩�<=��-���Z��n�xjs��+�_�����X}��*�n\�s'�/^�}�P�P������tf�t�u���!��Y�y4kt�Rb'#�p}J��o�d%�j0�����OI�*s��	��z���Y��sZ�/��ʘ"0���=�N�D.zX�]����R3���`v��>Z�y�O�]w������k|�`e�WytFTpB2��
��7.�9��+�i].Np�km�T|G;V۾߾H+c\��r�钪�c� ��rtJ������k�l���K>����d��28�.:��^�\�5=��D�C�Y��N7�a�$Jvn��I5�)wR�f��C�sS�g}��S�^��Δ�ׄ�o»$R���etZE�Fd,�č}f�κ� ����%=�(�s~l�>& r�piu!
�7l?��8�+�_!]�G�\�ꏍ�k"k]�UO�o�Br�Lw�ϼ/��X#���H�;ެ@���rY�!Z�����"�o�l�t=[]����B��w�ri�/ ���7��mp��/3���k�'�'���>gp�����[�͍S���<�g��3zǇ��|'a�j��c\�(�!��0޵/2>���[�W�vGn�SMʜO�3FM4Xo1�Y{.�$N���5�wA�P �5����:�/]sq��8�'�,�>~���I�=�k�ay�Hėh׫��]]"�?0�r��.��SwA��ZqA�DbT���l��!$	1&+&�q6R���5LF;eɆ~�@ɜ���sg�P176�\!��S���t����[��C'/1զ�t�a�"ﯝ(:��SL-�����W�1���M�q�P藄��49g{�n��|��C��ɏӶѝ�G_{d�{��h2�P��}��7Q�][��(l�7s҄����>�[�*�q�k�uAg�#)�;�z��EC��Q�=����&��f8��g'h
s�N��t퓺�H���Ӿ��@��P����Ǟ�75s��{/��vr�J��][XY���'��(�k7)���U��%�N$�b����W{�!�JF���t�/��#� i(��2Y<����P�Hj�CuS8b?PB��a��)��2N����AX��y�[�Zнָo����u�*j�j����Ѿ^��{`��"�-�ex�/�8<��&b2�*TQ�Uq�\�e��+�{f�ۻfW2����GZ
*����S�%��5�|�l���iѡ���37��bs��\HnN\���2�L�����8I���;�e�DMۙa]�n��,c#*ɘ2M1�})w_��a�0[�����Ĳ�swX�b������q?^=�X����ͪ�q�+6scHH�h"m�mp�uZU��ü�NzK/�g/@����ٽ\���.��A��:��8U.�iw�YSM�e���%�P���ٷ�՘���$�bs7��Ї<�;ڌ��y븺7�_����ݜ��kJ�`�y�׈1!E%�0�=`��o7��d�F��ք�9M��^Y��99Z�����R�#�gQ�%�j��>�����a�9^��;���v�3y�Պ6�F�l����SZ�Rg�ۣG~c�LvN��Z�V8��ݻ\�wr"�;[�YƲr�~t^/m�h%���>��f�h�sŋ���w�XJiq�3��I�O��m�d�r�Q�&NP2\MvlF��/"�Q*d���q>����g����x���ɍ�Ξ--^*Y3.����������qB�&���αuڬp���=T]��=+����o֭-�ʁ�m�tv�]6_��S�@��,�%�����:E�T���L��ca(�2#ƾ�����&.��t���*IƖ��:���;��R��}1`ҝ60I���^�Ë�@p����=���ו˲o��$Y�9�UU^����T�V���C��,�����]�'l��{;�q=��"̴f��RtȖ��$�ڝ��uj��[Y��R0�OjW���[���^�(
7�>y����d�2��fS��^V)�>��M�������^�[I�EV���6�q���z6,��8r���_gX��)/`�ǌx�9a�[1p_���� ��|��~@�o����۲	P>�p�8n�o2� ���G��`X�u��;�*ϐ��8cj�/9�M��Ȼ�Jz"���I����2D��B����.ɳ鱱���n���;�)/Tƣ:u}ں�;��Ի{��8P��S�WQ�t#@���S���x�=����ƺ���o��Ԓ����׳k�w��^�]9���S�i�|nk��V�G��,t�=��훉�a�Z��<��.���Q[^+�ZQg����8����Mhv�{����v��}��b�y]�/�=`�uk��2k�4����;�<�O{�l���dG��S1��i#ܺ(�v6�e0EǨIzx�$g3�4=@��\:a{�/LȰ��Q�?we��N�-�a'�"��΄��lx>ۧ������#Ø�=͝<B$
K���٘�>�Y���zvJ1ٸ�p��V�[eApk����V�s^���[��nM��n�f��,jq	��&�8Ƌ`���xy��~�����;����S�ߵ��35Nsվ�ú�S9Z���Pwǔ�G�!5�<1�
G�|�I��(�ʛ��з���"j�-J߲/�Q��T�����d��G_�%�2��������!��Ү:�w>.ۊض]q���Z�uC��V���?�<�lꑐ�ʱ>�B��Թ|گ�l��z��x��sSPu)�O�h�x��D&�
rX��v�R�Y���q�;�A��5<ͨ�Q]�"]wlMb��#p��Zݣ��WPs�ʫ�2��n;Vi]��E�Q��Ф�һ���Ž�]�}n��?g��;���
~�a5���p��[��ə�#���m�����b��*�����P�����$G�0�c��Ea�'#b����V��~�Rxϳ�}�5QB/�����Q��z������W8���d���P;m����R������h�"tu�:�azD_��=�=�f$��i����8��h����7νC�f�xn�{��Y�a(?���#���m��ظ��A�*���c	�ף/e��(��b������G��s�Zs
顧��׾�n�8�>��n�F�p���3�r�3p�Q�_N/^Ng7XX(���\�֧����a�g^�s�ιGR��74�������N4�@��ͬ�	�z�gGMeY��lG��zP�Q�:t�ޤ���"���zg~;�_v.�գ����R�ŒuqC�l��P[�a�>�)��n�7�ΰf���\'hl8�U �Z&'J?{��y_����]��fD�ך�_{&ͥt�{V���$@q�51��6��"�W�m�5{�ځ1��
w)`���Tp���c捕�Wn�eH�c��v��ʁ��ًX^�� >�	�T�O�H���� c�Ё�WLΞ՚�����dc�A�^�띞��m�nZ��y��^S�`�.�"P�=7�E�?�V�����Y+�f�"�c�{]7?5b�L�Z��n���ɣ�e��]��Ŷ���t@�X�8`���p3s&3&b0�h��U1˩L��U��Y2�z��K�������QTFH{����_�}��w�(pI��J����n}��d}��(���u5Ӂ�]Ö�K���I�>�oǜ��i�81:,�C��q,j�ٚ1��o��.�إ� 8�;�Ge]��!F��n��DNB3}�e��z����ڄ˞5�׽�����b��J�ԖtH�7�Gp��T�")�G���~};|���{��2��5�:q�́����٧�T��s���t�\���R;V���O�k�v���p�%�=�gH�D��%��+w]�� �X�=xg�!�)���� �".����tW!6�fO�x }�D�9�$L(�sQ�ۻ�w�|��4����{����+�D���9=PkL��$�ͨ��<`<\dz�0o�j|�w^��{F���Ɔ��=�Z��}�&4{���&8�K)J��[�.~�����vk�:��%��aԄ�f�+k�&}w���b�(��~;'�i�؁T��K�c�iNN��ճHOf&B_}�G����$`�6����q��%Z�`��]���r\1WZi(��D��~\/�D*؃z�)aD�G���{0��@�5�q�� _]�ɤM���v���4R�e���	1�����<�ɔ���wٞo؄mt���dUP+�d�����sw��n`�zw��ҾuR8%�T��1�t�ک���j��3���^.�0�̘s�Ҽb�A�IUTc�us���i�Jy�Z� ��x4\h��N�Ўz����W�F�x�"b�콫�ثg�#K���%P�#@�˹�u���zA�N9Cb��-��k�W�3���Z�nڝ���!������F��47�@��C�%2�]~`��ȡ�Mr%N��)��w�ZF{jp��)ϐ���F�7ِ2�3+�ͳ0fgr�H
v��[}���W�qm!z�|�������9�I-Oy�
`�	zy�������p��QљS��SS��jǎ��3x�ϡgL3s���:cO��T<��41�Ɓ8�t  g���r+&&��y���j����i�损G�ǎ�1��꽠���y����~��x:��G�+�g��&���Tkj�!*�c�{~�4	Z�8�,٥>��y��n��7kn���o���3T�쉰ːd�:s�ò�-5
�5Gl5�OlB�f�lKY������'�@�P�p��
"�>�]�����u�����cf�\kk��!�XD��~��w��Q���Ϥ7fR�p������d�w�/8���X)��/��GJ��i�ʞն=b�q�:'��]��R�:�ktuC��/��u~�AA�x��c�|"�Z�-��̰.��g�U�Up�݈�&̺&���U�P��O/�ZRV
{A�����8�3J��w!fq>&�	�wc�ڜ���e�"<t�&o)gr�>����A�8og�Bo�y������&uq�^��Bϫ�!ݻ��A�3����0z)�sT��{Ѡ����Ϧ.o|gB�&���|�u-K�XRux9]!��#�� �@^�a`��üz*@���s�~1��Gٍo���Dg	�	���k��C����ޜ�[�A����3zT6d��$���:������2��u�=&���,�+���-x����p���/�i�D
��av��Z+��|KG�hNN��L��}Z��2�FČY�a���g6�xˁ?Oٲ�=�v.u�̌��̠u��R`oa��W��x�B'���>�����b͟3�U����q,%�W�2|i/fI��{e��䷾C=������}���s�3��������5	�j�oG�ɛIl��ҕ��F�ԏq��1���<��J+F`3
"*}G�kOE����AY��#�)�Aj�}�Ѡ��:"�l�x�e�Y��\��i缪�&�5�e��z�v����F��DZ\b������z���:Kw¤	��	"���zF�x�����s#�&_��u&wo�t��:�W�h��N���h}N�.+6���g!Nb:	�{�RWM���5��d95>��cZ���M�5B7	�@���OGt�!�)�'b��gw\�V���+1EX;�ʒF���&c���.Fomu����f��Sԩ���?d��no�D�{m�ڇ�!�#����M�z=w=QٵV�H�cM�b��S��>����$�b���鴣4�<;ύ����ྱ0�����FȮ�9�iS~�R�,�KUGm�lg�.}h�uw�=1��q�q��2��{����P�!�ϫ2òC�v�d�C����D�����qv���Gھt3�+P:;��6��Ƿ�EǷ�A�����1� �Ve��h�N�eP>��/(Sn�t�?Qp�g�R�+�Em)�;IR��S�q�M�r�vj3��'���viy��"��W.�d�˽Qx��=�t�L���{b��\����]�Ү�q����V�Enw���4E33 ���x/>j�����OrӾ����{�M��CQ�D+8���o�: �P� C��cS�������V�<�.���vɪxՎL����!E"�
0R,�~�׸<�������Nh�VbJ�wwT��웒gl�9�:�ͻ�ì��Z6�b;�E�<v�YO�����w��c�:4�:�Z3�5���g�ӽ7U��:�;��m�����+��;A{�4wZ3�i츑q�7%��E��=����'y ����Do��,p�؝�Uz�4fŻ��d�b�1�1�7���&{)���6O�Ԯ*��E5˽up����w	��+�m�]
�Ԥ����������'�c�݊�=�wt_���5T}f�ϊSm�4�E���k�i�u^.7�]��^	���[�쑣x�ۿ�7�(]��.�m��%��ޑ��6j�%JU���uD���졳�}�W�0C�=~��F��黵N�����G�x�|�ޕ����<����7\l�=N��W��
�:܌|��B�z�WG��"�ݏ�)��� �����h�E�X��+2��m �M�<i��Q`쾹׸v����ύ��\�j���Tx�q��F������pMk*�-f���]Mt��.uJ_H�X���6��L��[{��Y0��#^M/�t��]	�9Tg���Y$�tUq�+p���ŷ����t�ٕG޶�{���~���d�r��Ҏ#ܬ�Ǥ�e��(Z�cuFU��zN��;)�9+Z����޺��jⵇ�ml�Q݅�Z��5|�=)jUڗ�\K+�?U��L4|�	't!����
��<k����o�C��	�������_������F��}7d��Y�"�J�4t�{ޝ�P��l.��������ڀ��-K�s9!�V�G�us�F��^�+|T�F�Zz��WE�L�|����Z(��XQ� �^;�39��<gsW����L�Y�O�	�ɮV�Q�<�6�V�P��ޣ_t��ҥ����y��:��v������+�uB����q���Oym�vʥ�^��.��r�>�R�2p{�{�I+l�B�����1�i�C��L�F�[pm0y;�P�xЕ���c��#�ĝ��c�N���(jS�k�+*�ΣJur���� ��-�Nca\�����t&����AB-LϢ�ٻ���ݏ50͓kP�(�^#�� Q��>�����S���CM,���7S��Z ��C�^!A3l~�5��RD��`�[�S�d_����|n�����C�s��<�����A?	PN��Ȩ�n5L�h�s����Oy��}�[K+d�V�Q "�R1QE��A����w��s��;�����;CcO�y�s(C�D"4=�;[\V�R�yr�gw;�Sv�o`�8�[͆{k�6k���2+i�!�~�VT�R���m�1K�轪��x��ym1�zf9���'e��3�ϰ�P��L94�<�h�j�ab
s��j��R܄f��z}j;%k��=(aX�%"Ҩ(��\>��;8����Aɼ��tD��ۉ_�{��y�XT��]�w�ǣ����NU>?,�.��a�E)��t��a�1Ǒ����5�o��luˠ�q�'��A+d�܁�!�����f�yj6�ƪZG������&�����@�%��L�U�Z�����Ţ:G��5�KKf���vȈ��|��^G�AQ��7FYriZ]'�Ί&9��fu}�;�zED9�yeZ�賧��c�XѲ!<��(�3���z�'+qJ�]�+�^�xk��6rp�r��1�Z���s�U�Lxo�]gD_Jj�2ϋi�|f���cT(�K����lN��?_j���C���N󸎨U��7H������������gע���ݺ
�<{��J�9�3���A�fq9�s�.��L�2F�9vC�z�#PҔ~�<�@QӔ �0��9p�6�t�$�ީ�B]�Z hy�x�ή���h��w���$˨��,�ر�f�u.��հf�t��I�d��=��N���T�<�s1�<ж�Y��]��1��ke�}KtV��^M��"ۈ]�$oWB�zwL�v'Ka�u:��w��� ȝ�bfA�o�S/
��}���hϜ���$$���$$���/�Y$�����@��$�I$���1�!�Մ��	B� 	_�@��?�a!	k����$�����I I7��	$�$��������!$�$���Mj��$`n��5e�ȣi,����aan�|s�8�q=����dM$<	�={/�ZYm�m��9f�ȉ��#(L�Js �M�y���D�SC"x�橉I�o=���l7)��񊔠�[��6��u*mn�oL�OY3�;R��8�e�0)�KlY*�Yt����5�L�0��êQ��d��6���;��sMi�I^[PX`������>Ȭe�0\جYvw)�p�i�f����6�ku�� ApQ;��nm��(ԭ$�m�&T��y���d^8�V�V�nȭ84��K�z��zt��]�,��o�EH���&� �;LU��[.���FXg�� P`*�b�O7��Vz�� �вe<r�\Ǌ�h�f��YNn2A�P'3(�u�B��ہv78<YfOf���>��o��H17fB6�f��w.�t����٢���@rƜ�����n:��h�H�0�k6�`!�"j)�Ƕ�f���J����v�<��E@ˈ����b'��0�d1iE<�f�H�6E5e��$U����G�/�MX7}J�J�
0��X��TAD��aM���d���n��˽�g2V���I�l�z�O]2KqL�{)Vǯ1C����ٴ�\�`Y{��� L��]�
������V/,a�����c��݁;����[�I�[�����5�����:��sqx��L4�%l��/hk!�ւ�,S�5��e옌��P;j����j�b^�d�ܔ��X.l5���L��	�{�tФ�$e�[ں2�Esk��b�SBf��C��цɊ��Ɗ6q��g|�935��y�œl�i<lѤ*��G7Ѭ��y���z3|�2ʡl/|B�N �Q�2R���7
ݼ&��G��r �Uu-�lŹ��N���O M��� �1ˋR�jFr	�na+��L�B(�y58���ཽS5T��!6kgnhE��G���48�~x.��eЬ�ɒ �2���)ӌ^�j��2J���٦�2�u����4�b�Ly�R���6�AX�Q�hT�Mؚ�5��wJ����$��-ucHG�´V�p��Y�I�!�1$�db��끦+,c�i��[���>_*�\��	�Z=p��v	�p�ce�B�YXr+��f䘶���t&߀�[%$ SE�"#���M�ِ�,%�F�3�?n���������;���^t��:�Y	c�q��OE^��^j)Hm�խ���<�?�ē�V��͉�~�[y�L����v\r��l�����\��Ve�4�!�v�;��&d��m�F�P�C%�t�������M���n�+�[x�u-��|&-~������ͩWn�&��kT�Zx���9�7
��]C��l����ڷh�!A���0XkAI����7�����o~������Ԫ��p]��y��.8w&�)�с謏?K�=M�Rt�C����=���YW	����>���u�B-Ff��x��n{5�$ �挀2YAu�v���h�DQu�]�)�@�lL�yK1=��5����`��hU�����H5Z�P+/�hɶn Au��~y������&L��ᾢ��i�"V���Aq��eɅ`�ޭ�/��AZ�x��i�e%�|q�N汸YtKM��4R�h�1`�#�����}���F~^ݡ׃cߛh[��Q����/nz�͑�`�6��d�=7۩����nQ�����Սo�(�7h��Nl~�@P؍������8Rbn����Q�4imQ.M������d�E!Lz�f����L�����e`�DylwD�n���{If0����o��˼�-��y%ˬ+v�:nb3/Bl���nӱ�V�Ѫ^�4<aIQ�x�r1�G�4b�v_<�p륔��;F��O��E�+qk��'wn{��5��s���u�Y��p!	$�	! D� �	$ I$ 2H ��!$��ђI$�$AB	�$ ��" H�I �������$���-�������I$	'�������}�8II���BI I<BI I?��d �,����5�$��������k��F�I$	'���@�d����BI I?��@�~�'��������d	$�$�o����?�߈I$	'�-`I$	'?�����d�Md
��σ~�A@���@ ܟ}���<�ER��h��e�l!"�b�R�Z�h��2���PF��1%�J�=t� �"�-�0  ����E(�H�
�#�UJMd�A�U		��D�H����H@ �	u���6eT@�%G�    JE	P�
T��"T���  U}�9JU�Ͳ)=�    P �@ ����  �@A�
�aX�6��Ze�k}uty9sV�+��E�1�Һ�:�[��L �h���E�%���t�K�]�� K1��k�ݫlچ���6ݸ��gw'kl��
RGmJWY��
��47��yv�ݫ]2��F��۫BAAѮ�*� !8��d�s'gdwQ��r���C�i����]k5��wl�����t�\�-�IQ��D� ��t
�wr�htt]���S�YRtNs��s0�˘i��tꈬ�U��h���d��ͪ빭�m�N큡]ٹ��v:��9�ET�5��AT�m��3�������7sQ!�Gu���p3�)������ֻh�blkY���'QU&뭜�]�
�qUR�\��M��g�I]�
$R�U��x���a�+�W]V�v���)��w�ݶ�X�gd�f:��TF�΍��]�n)�i��iکb�qU��V�E�pU�ԗom����;w `��	*�X�V����u�8������93����t�wl�c���n��d�3��k�F�w �βU)�U�U�N��InQ�u�E\�UJ�[$��dDT!)t�ʪQt�85֝;��h�J�����Р�kZ��9N*E�[�U�UD�v�.␝iU�Mæ���7&�!l�s.wt���u�ґU�� J�X�(�N�ΈRJ����5;tC�hi]�1��:�%�Z�sm%�vI�aܓn�U���M�٩J�S:��N�.��GN�P�+t!W;S�k�E
�H�UHSZ���@M�nU;a@�C����R�]��a�9�N�Xr �':�ܝ�R�����������((����Tw*�亩��j�A��#��)J%%Q�*U&��]�gt�(�w!�tj�*���Υ.�.::�5��S����&ݸ�,û�	U�;v����ã���RB�2htW:Q��ϯR�T�U((֨�B�*U"�m��%%RI� ���b�R � Oh�JJ� 4 4�I=F��驵=L��S�A)*� d  j��4����   $�@�T�&4Fdɶ�c]���Ŧ;�;�3�d�1M#�0Mt�����]p�}ݚ��u|��뗿?�$��I7�m�x�*�EDS���+�P�����
�B�+ZI	 O2HH��e�W�R(�'�eH�+*� ��J()�,V��Y:�gZ�$�[%f0*�L�x)���v�hG���=sɗ�J�YAZ�L��B�����r;N�Ϯ�{XEh@��7��Y�mn�e$���[m�t[@c3\�YY"�"��ycKC2���4[
��b�-'h�P���*{2�]J�b���dkFT�+!V�fc�B0���j g�Qr��Y�!��3M���{�KT�c|v謳��n�%�/L֭�{B+͆�<���d��(Zt�*{%AV,��r�-�5�T^�T�W`b֡��U��G+�i �bw2*�x]b����5Vp�D����x��$�?�qpХE���;����Ϧ�Pw-5�E�V���f�i���u���ʵ����/XrQylt�Y���D��d�v�nb�B�F�U*n�GN����ԾwiQo琻l����	[M��{��n�iwY7�aKJcI�Y6ºq��@�H�QT'4����/��!Q氊,
���`�QX����ER�1��E��"��(1��TE�Œ�ĕEQFc���=r��Ր37�l�q���*�R��T�(�!$Q��E��y�]5w*Qڴ!h�չEV�a��*��	�{�8�tay���>ۮ��Ԧ���ORd:�,Ɗ�9d����Ͳ��:��钺Cw�t�7���|{��m��q&��i �=�w���P^S�%+:��\�-٭䦛���Nh��d�����)�i�4+�����V¨��e<�HT�+�[�e��KP7-چ.��r�[�ZmMܭr���<�^t��K�:��)В,@��U�6,��C7c��LJ�"
�ȒE=ղ/���  ���*��T��π�Nެ��<k2�{�V����=�<� �I�FBP� *2��y�������n[�f�v���Kb��Z�L���05"@}#���WZ��V�l]�ݼj�����
�����k
v��6���V����D��5w��V��4���D���L����$�N-��0jXT���%e��0Iڼ��IQ;��l|^���u�Z�JJ�0���4�бw�n!�����)y�u6�{\�1�"*ă��Xi�SiX+�Ȣ�N��ߨi<¤ ��b���Q��O!D��
�Y,�4'=u�6��éY֬2��1�1��"�����'�P�F  Ȱ�`
@EH/y��{C���:�ac�^��!�Q�1|7�N�+%*���@�e�B�%H�+��vh3�'�/v���f����Pr��R,���2��_�)�n��Ģ7n�R�@A��3#J��Њ�şkon��Z�5��^��ʙRֹ���v�l�0V�Y� �S!�/�!m�ȯ2��KeU�$�1��Pԑ�RH��a�����rpE�;Q�SOfc�+%^'��Cm[͎Ȋ�t.&K�Nҥz�8���j��+���ה�FW�-�0P$��a�6��՛�NnM�Bl�U�E��6�_*4TL�ܔVAZI� ƒͼn�ᐻX�۷����ч6�n
�c��`[X��T�  f��*���c��U�yH(�Ay�䶌�tk�WXٍ=t�sxg\��x�Ws2C�CH�9�('W�`Hfd����6ܺD�wre<T�T�ǹ5�L�қ�$��YsvΨU��k6$�N�t��\�F9��N��@޲�j�Y����"�t^=Ԉ��-�5Tkl;A��]:184朇`I\ �S/ء(��-�b֌5�4�W��G���l�F�bSgm�X��*��AS�cN�fIr��!:������Y��--pHq��q���4��DC[*�j�i�����S���e���V7��R��� jG#�Jx�4n�m*�w%n�#Y�5�x�z���BiV�2��$h��Pѻ`�nf�4�X^� �{�i�$��;s)��Wn��Rcɢ�m�F�XC�_]ˤ�ٗ%�y�e�men�2�*������ݾ��'uHqR�nv��g}�[��׵���3D<ɠeI�z���*Ld��咳V�R��m
�$�SIk�1!�(�qi2���(ӣ���b̡����ւ�ɴ�%����18��sƵ�iQ�qk��@��۠J�� 7����fW��]�8�w�͗ 
EI��!�
�!����Ö����{z�yۂ����'��3T��/�#�n�f�4�6��*rMٯs)H1}b�Hİ�1��@f]�`�To\d��E����ew�*:�(�*�Չ)����d'Z�b�Z#$�L�ʫ�Ia�7p�h\�l�ž{Y�Q�A�����>�����_P�7&ۥ�j�����"��R�SQ�zӻ�7"*�1��ee;���/2Jz��tӺN*A
�t�v7�1ʹ���z�EB�<ʒ�*��H��dv���Z:^�HǷ�n�C|Z֖�f��j��K�y3R�j��wq �*U)����`��VN��}����Ij�������v�FZң�;�7-�c�(l��Bmc���f�FJ��[��s5P���9q��KA��De=xd�*ŰJ��7��V(#B�٢��t�=[��+ī4nC0�����f����H�Ԥ�E���t�J" �(���^��кs4�_�mV��j�m�IFΉ-b��I��R9���߅+`	��n�w(sZ�Xԅd=���Y箪3�^\Xf����RЖ��ȓ8wlӌ�H�k2�5su��� �4Y2͂>LŴ052�\)�kj�^c�С5���H��@�Q4>�}����d�q���i0j�R�a�����e�R�K{�T���mٺԼ4Ь��fK��^@�tmn5r��R���f;D���f�Ѧ��
t��m=oqZ��8��[�{�N$kQ��u%&���a"*⭆7�5�W%��"�D�jyCYU��d8�t��=�U�T���"1�wA��d(BT����TYO8��`өF�W6��zb6�A �����	��.dcji�pj�%Қ^Qի!Y!y$&�b�N�����>�P�vʨ��V���ږ���c
'��Rf�C��:7j�VA������W��&���x��nFk-!,�x��D�Wnʼ���EPJn�ئ�qѸ2�;�kj��h�9m��LiQ���D��-L	����[��b���|ެ$�a�y��n#����A;9,%vU:bl,����}�zՄ��E�����[
��dkVNX�{����^�T��ɩ�R�eC�y�/�	ԓ�foQ�t��{��k�Y��B)6�*#dP� =��f�ú}��3�a+�RV����o�&�C�.�r�	���\��{��j�����T�$����$Eku]���=�u�l=�`���U����}�0�6i(���p�w�����v
�X�]c��J;�DZ����C"̡��9�uN��3NMv&Q�" �����d���))�0�h#D�ɴ,
�{�jf����E�D״0�ਊ�c��,�л�^�}��7��5N�a�!8�sE;��F��w�6Bc�l��~�u�k[)v8�1�����iXu1�q&�{i�g�B��j8�>̾2��}N�	\E�Щ=f�)y�tE�nщ�Mf�Ɲ!��k	��ݧb�u�A����pg3.�&<F�6;oR��?�P� v�v�r+��#{�[�t��N�����*I�aZ�K�U�U(�嫼��,��e�W��n	��8�Tm��u	m�!Eh�@�E��U��7��@ӻ��fT&��JVj�K��e�.�A�o-�S	z* bm$o)�Eb�r�fәb��X���N�ˑ��u�&��뉉�C7v��u7���wUu�Y{���n<C��� �si`�1Xe�y���`�va*l�_`z~�d5�N�[U@1[��Vw$�������FtGk�	5l4��54�0��J��z4
̶w��%C�B��Fj�Y�j4�ϯr�c�W'�+��x�m�u%[���@�.�t�x��^1l��*�Z�8����tn����L�{�f���O�$����s{o��5}�{:SWjUF�G���lP�N��i���*�`�Sv .)weP��T��򲋼)�,��ͷf�M�,q

�|�B��(ࡒY�tQ�q��e���!_}�n�"�QM��*������|�8��$�ZF"��6���s�$���|���F��W�5�}H}O5�@	(j�I
�-v��%h�|i��j*��`Z��r���j���������(P����!��}_<����6��R@�_fiG-��%hlGN�K-��d�,�`R�*-ZV�2�Y��2���0\��ҙ�͊4u��fe�T;n"��ң�L��1G��eFj�Zp���RfQ[w6��p^:՚
�m�nZl�6���(�/����aɴ�s+
,c�-c&jm^Q�+2�QmDY�X��U���֝����V���t��M��-e`�&�ww)�"��E.�S�`���K&��ӷy���|v��+¯tl�7[*�Q��s%��mF��e���b:�K�-+D:vB���.�
�b��+Wُ�j��HŌ�Lʴ��S����j��	��0�ը�ZM8R�h�T)�� h'�+��M�j����*�,�AS؞�c7`vj�����T��CVi!L��b:�pʘ-U;:њ[�´\Cv�l�2/���Q��`C�̊�[�@g ��^Z �w�� ���iR�Y2����Hi���5$�-;����*;SY���-�j�^I����G �H+	F�HJ�)
��.�t�٥����eitwuM�e��FޫWIf�͂��"���#5�&-��L�LB�]4D8ʩ!X���A�H��CnE@U���!UF`y���,8����T��d8��M��I��bt���f����0"�/��a�3*]�6�EV+)�RƠ�%dCN*�ظ�.��`5d:��b+ X��"�J˯��D0��*�U3�7Kۚr��R�^��Si}���bآ�aJ�wVWXpSy�gt�#�ہ�V*�Y1��r�E�i��3QD�����}�e��Z��S��;���M�3���&s����ۧ^�a �Bq	�
��C��,�aa�N8Ԭ��g�Ć��*'��v�i,E�ذ�H��$�Ne@�PQ{h"e�`bB�a�,Ԭ�j()��1�U'iX�Z�Τ6�(@�`�HW�۽I�����m�zw�v_j�<�퓶��o�C��m��FHbb�N5"�fYI�5J����4ɡb9lU8�Xe�m
(�ET�DE�y���+�
�C��Fq%gP�:�����f$ݫ8��H|�`�X�P�D@���`|�b?>Lb'�,�$���V0X��b�E�D��Kk�d��1�*O�DZ�E��
cb��*�R�AB�+�*��QV7j*�0b��y�3�b�-;h�)�Ď��%U`��6��IU֌YmX��,by%G��{����o��h*t�q��j�М��ܾfb1ea�7]����y+0��v+'TɎ��J�ӎ�V����&mh��{��w�w36;k*
\]�[G�����nڵI�M�4)nRc<�P��`��Q�Э���ߞp���!�%>Ѫ��ٔ�].CU!�Mn#�9W�*Y��$�5��4w�f�.� �J�������EH���QR�ia 'eB�guFv7B�fwh�:�:&�;�Wnh0j����D�h��k��D����&��Z�;���hӝZ��ծ��
����|�{t+��j��V0Sݣ�)�X�����v�Jj�������G%�iL�/��] 6Q��R���&��U�V֗���L�����B�fRO���*렳F�g^D�d�FTwK����tA�鎛�}���%J���Қz8Mu���Crm�� $smZ�O9��֛V��kf���;+wJ�\�0�V�m�EK2M�;:�5X��>��}�s۱s�6�nT�'�X�9ٓI��P��`�g];53�֡�Sxl�"�`D."B��=��9�sm�ˮʔ��"ގ�7CMx�]K�Ӱ���ǧ;��1:�MP�&�خlu+����W=���FnbA��6��@D�}�\Nuee����}ƞOv��S7b;|��k�ҽ�+�m�Ge�j'�T݀�mQ�=ۈ#��dɸ�v��~��V{	�v]q���.��֤"�|���[������KKѐR�#�螝Κ��Udn����qVD��r��#��p
�͹�g��+�����T�(Q�/�70Ȯ�eZ����Ӡ*F���+�.�ų�\R� ���JB0�\�v�`�YZi��ۦ��Ō�f��`���$��M��G��3˘ގ�3Z���_Wk��[�Y��s�J��!2�yկ��<b��%fJ	�SN�=�ኄëzf�`;����ŎԞ�֯{���k%qW�ןwkYt��*��4���$o�`��Jiܗ�ݽS��d��(f��aC����udTƓ����{2:4��6�̕��3w��; �q�s�B�e�@:��֣n1���<����V��`,��ٹKm�x�c�^>��v��KNN��Օb�G�>�Ajvv�4�7�I�Jײ����'rf"�+;�^��" U��b����Λ	W�i�2l�&�SN:0"������U���������V9�N�Q,sl�y#-����F����X�S�Բ����n�*����gP#���}F��U�d�3蜼N�*Cʲ]�FfZ\p4,�{�TG��
 ���r�D�β�R�y��8ާ��0qU�Yʘǵɪ�+;)Nx3N=���zㇲ�n�C��'D=�^�:����(��b�|����� s��I9�u+���S��^�W�����	7��V�V��F�����Stc��ֹP�:�/�׵0e����[p���}`���4x�3�.S��@r���L<��v�Ԩ��'8#X��R��rc������Ayj�[Ol�}��_ȶ��\��0'sD/�5|6RB����Ʊ�qWd#9#�kZ�3�]˙+@�oX�Jmt����7�R�ۥ-�A�e�R0��]��%V/fa�w#tA���]�\I3��BP����]����wh�ۣG��/�	�t�1��Gڕ`:�E�7�6�h��(��T3%@,3?,ׂe�޷�i��xc�159m����-�O�xJ�wt��M��g�{Z���`I6�:1_.�,�ۼ�C�Nb8]�)C��NQ�u����P[��5�(h��x#�����.O��}o�,9�[����5l���{3���������@�O�����s�*�ʺ�9pk��Y`�ߦg7�p�}�w��pWW,j���:{m`�v׍L�},�Y�u�$hdc�]��nqnM ���m��6/~X�5,N�X�����m*�wMg������4j;V �h��Oi�xS��o�8l9��b��W~;��������I�V��6�����̀6����U�U3_r��YoQ�)�JѴ ��,9uO��V�d�HFdK�ag+�wv�Z��I����Ƌ��|)�Is-�u6k�'@���BA+��]��TX�V�xT/�7�'m��`ˮAˏG\r���zuYe±�gUŪ���۾heqj&|��s4՛GF �s�h�yG�'Z�s�\������ιW��������Ȭf"�s��G\�x�2mkU�U�'`��_T�ξ�c1;6�h;�Y.��a�ɋn:���ٯ8������l՟���^��.�������"��ܪ�B��ݵ��i�φ4(��=�k��w��v�D]�����Y�C���xr�r]�^�x�<�*[8.����t��G-�P��ݼ�M��n���Z��0�v��c�R���"f4��S8d�����q�}���3i�C�*x�-r�ޮ��2���u�A����1��X�f�9�vE�i�]�F42�S9�ݦ�[̋�YF����R�f�'6
�`y���AD[ެ���z8��dON�X�N����\4�REC�������C��Tᣩ�t]�;^N� Q���7�;.�Pyb�8�����fTc2K=}��'^u�叹��x��0vk�x�:.�3n�ٹ�^���]|�mP,�Mu�*Տ��l�wOC�@ʖEu]�,�@�fn�'���Wr�h��y����'��M���)�ڪ���8Vډ5]�޾�?7��V��.�*܄ݩ�d9����h�oHw!��w\�m�o����rCC$ɣ	�X�b���C}��u��K���&4_�U(��^8��y&L�x�l8�DV�V9�ևQ�Z\�P�#pfb���dU�ͧ�).Ƕ�=��·J-���}�(�\�s�5n���9�sҵ��F�:�̗O������s�r�MV+�q��)r��fV�
����dn${$�����u�ut䳠@�7���y��O��z9�$ܫ�#V�wd�b�IC�W��fB{0>�.�Ѷ�FA%�4���)�3���Y:�`��vS&��Ig�H`}[՘���^9����8�%����z���̴���X�R�Vt"Q�s6����K���۴�`
',7���S��R���.��.�6�+A���,�Ԋu�B�b"���XZ��j�/h��@!�a�փ�^̝,�����;�m^J��5/�U�@�`��`fS{���m,'ۛ[�>�a���0��(�ͳ�wO��Ji�R7�@�UK����0�/���:Ʈ+b��W��*�����¬Y���L�0�D��&�\���A�V�*�;�6�A���]�=�A�&��Q�XU;��a#:�����X��X����n�
|0r��M+Yh�ئ�uw�z��)����s�FA��є�<d�g���&��wz�O�2�PV.��[����M��+�fhk����0�΅��ܢ�[A㫍s���6T[��^=�p����bRo=׸���)Qrj���+ƴ����Qwm�W�9�2�v��?p�C�jZulgc����.��YM೓kS	uYڻq�.�k�xo��]�&6d�y�a��ݺOX7��3i��{vs���fr�pM�g�hf�]��#�u�k���u]��U7Ay�����It7��V9h:go�����Q�d�)��������� �Q�K6��U�bA�5;�K39�v�聽�f�x�c��-��f�
����a	�2�I�q�0��^]w!6�t�����CHlCq���C.v�ۑ(w-:� �Gʉ�+�Ӥ�ʘ�N�լ�:��nm����]��I찲�s�3�q�}�����w�2�M��Сɂ�P�܉��x�i��|>\^m%kܮ}����w�Ms��m���y=�i٧��3OW(�*ݻ�ׂ��u�;�Z*l��"�9���!�s��j�����4l�ʵ�a*ڀҜ�֡'D����uY�G�Y�wdO]�]Z�bc"�$�Pv��R�cܾ}�*h^gN����&T���i��fT.U����}ݷ%���%m�]JU[��]�6�z;xw;�J�y�苬��!�y�s��d�1�uc�vz�%<�
��mY��Da�� )�+N�Xxj��2�;k�_o_m��V�2�c���!y�M�x�*�:���J�����y�>s<��k��\T��^ֱ@�=&Jv�o*��ϙ�����#Ě��If�O�.��.=�/zC �����D���|�J)8��Lݻ��������ךګwݪRoY�R�ߛ�ڮ�Y�0,�!�.f3�,b6�G-�b�:ٺ	��2	��iqw��$4ҡm�����-��
7�1��͒�a��2�=��B�&�4�>�ϸ}:�EG9��e�>t�����^D;O� ���nh��W����{!"�;��N�p��e��$��5�'��+d�r���".]�xS��U/C*������r�p��.�&\�B��ݮ�/�Ø.ᔰ{�v���n�P���V�C����������G�y�g���`}{ûrEK���<Dok���}K���%������{4/�f-�Gȝj-u�����c4�c({����B����t���o7;rG��TL�v���!Z5\�,�ڃWlf�h���l�@���̌�k�u`�f�CM!(Qot`��ޤP��N���q@�0Ţ�V��d�����/3�Q�����[�6N�T�)ޮrN|��핹���:�~�9j]��GT*�n�u9I�P̲�W����]�M˲����t�� �jćD���{Q���9o��*��dY|��})B5<����w5I�{�I��S7L.
��}[F���9)(���л���-�]WY�<%k�;4ݜM#4q��96�$��6�Dn�i��j���W�Ưᮚ���������z�U�
m��N�1*v���t�^.���rcI�\�.��72!�_Inނ��֊6淕�!쮃0���A�oH�n��^��x�)�ղ�KE�(8��e��gw��I��4��﹦�3lrT�fv󑡢�Axe�ږ�9�S�',kjt�3�Ѧ��yX���ˇ5�)	!:%����z.�Sa��Pk�7"����M):F��V��]^���F�u�>j��J�PZ����6{S|�b+	ous�,��E�	�)��9pVnh�+j�"�%'�x�|�%��H������Ħ��r� ��:�pl^�UǦ�B��^�;K���^�f�܋���	ԃ�P���/�3�\Ij7]�L1h�P�3"���rU��� l�睻��Kk-n��b.�_k�ݦ��[�*N9.�89�np栍\�b��������o���y^�3��%���g�mWv�%��vȩ��J�E�T�r�aw�بQR `���`��\�D �gyuNV�m��N���P��C0l�A:�Cur��炕u6ul�ycN�<��������P�ꖭ�
�y�4���E4#嬍�JL0��у�}f���)��fg+ا�fSآ���]
����������nnn��0|�h��$�]��C�����NɁZwf����G⃒�&��^���"�5� 5_cXϣcc��ܩ�����I�t�|k���a}�����Cv��ۮT�d��K��<{v�Q�֍by�o�^��%ң�����П}E�Y����p���ޗ]Ö�L��Y�����Qym2�<�aɍwJ��{涆!4a�xO[⥃�Rx��c!�%F������:�oj�
��[ǳ���*f�=�Py�����0kJ�.���7�>��4^jt�h����A�i���Q��CW+/&-kv�(�\���Q@m+�.�b���f�,@����yt��z�^i,�n�4���wY�6���n��T����5�$��:E�B$���5�Vf��9tt@�Ž��gER�_d]���о��%Ԩ� �;�q�Ӷ�U�:�º��ff�vB
��}\����LSc{���s3�m"q]A�.᪝��5A�ηƧ+�U�������Gi5l9o0ɇ�Pw�I��Qn�=�{]j��N����g�e��֫�0Y���1�Ѵ�h;+���լ9�����+��]�rjtھ���e`~d7aw�nLx�"�V|�K�얖;i�mF%���u`��Oy��f�q��.������ۙq*{,`X0S��p�x�����PZ�T��i��\���z�I��{rGv�']�+۩\v1����7x�	#k�2�D�[���]\� _�04���WZWx��+_|�J�MƂ˾f��FWd�:�zg.���Էor�����;(������`I^�8�4rV��i�څJ}��W�3��Ѱq�������؄�w�6�]G��KwN�*���YX�n�)v��laSy��3���ٕ��ΰz�@Uvަù�x]��u�]�iZe�U�a��R%���e+�N�N(p|��p*R�|�t�FT���˦]�ݵq	��H,�ګ.�"����c�K�x.�l��Gٗ�l˄�h�]j�_�����h�Bn�C��	�g�.��ʒi�Az�)B)�6�l���Y%>�`�s�gE������b�1;
���j$J�.��:�Wc�0���b���$�ov���Pp�+9N���1����P�蓙D&2<�/��%�v�f
S�������d}!�î7��Ֆ�^@�c���@98��l�K��BU�ݨ�J;�V�UfmG����y[�dk�5ϯ9߷6�����4{��@$���BH���D	!	�@�C��
�H!O���d ;�@4�%B��!?�I�Bc �I:���z$�HE$?�Y	0'��M$$�BLI%��8�a� bBm m$�ӄ�\�@ݰ(�$:��	<����'�d`fP�n���?RC�X� m�i!�׵ M�X�I�C��Da+"�
�$� q �M�C�"!!�B)֐�7��$�C�E�T&!��`@�	�����@�@8�hK�H)11��P=C�}�u��<�����m�q	=�I���%`V�V
\���1�� m&Ь��uC��&"�v�f�BT�=�{vE���	�I4�0�;�NZbԗ��M������+��{�I1����\�Bm�#�!�Hg�6�h`�u�]���I�@��L�u/��	�P��2l��1 �
���N�ڡ�8��E�;���u���!�HO�I;�!��g�9��Hi�9�d���~Ԁ�C��n�I<�`|�$�J����J�9�� y��ұ�/,��0��Nr�E�r��N��t�l�ir��q$��2�;I��6�̝��Y�Y��ް�o�l+�ݡ��S�N0�"���>�:�O�`����Xc�ę��EgR���Xw�/��]9���ߩ;�oF�Iל�w�p5�<��ߵ4��*u&ӽ�s@i��{���s|ލz�}�O��q�6�ް�Nr���6���r�$�ow���8�|�r��e����|�03�=�4�l�z���٤�����m�a˂k�.J�I����}n[]�g}O'T�S�2kT�)>�6�5�g��`e�R����`�.&�j��?h��X���jw.��E�,��l3�v��Ee;�gf?�--�vp�H�aJ��T�����U��
CK���G1�06�1<��u�ݹ�Y�ט6oGU�P�?1��j�<K�f�3EZ��0�`�'ƫ�*����<��v��@1���r��A�k	�)Zס�b6�(W��Mi�X&��T�ˮ���F�ȫ�)n�t��т���c��ElS!�Cy\�QY0�)�#�F��> wG�z��t�[ʏ.�c��u�R��G)�	b�Z�n���p
�A9�U���Ml��;V�S�&Ć��VJHE'�9L��Ձ�]�Nϸ�ci���˙Vۿ���rSw���q��ؑ���u�G��	�X]^��4s1�G���*��|�f���@�e�N������?�eZ
��4�
�qK�C�鶛��v���ЇAzQ)7��f��S��|)��e�2U�$j<6 ���tV	�+z���i��;:��$7�N��ʫ����|�*�e�֐e7g�j&��Mvv�JnwØ��V唘ϒ�Sun��cV�u�r:� C��R�`��Hkł2\wt�ʗ���-8�$�(�z���b�U��:H���)-���!�^��Z��U��].:���S�]���}��5�Р�K���н|�&�^⳴���E\�[�[Y6��9z���Qb�ju4���E����M\y�n�!��	���[��N��t���m���.a�&[mn2������^�q�f���[Օ��+t�4�A=G��Q`u��ь����V�G��kxXr❣��wض%��/�Xt9�V�0,%aܗ�M�:�PDTK6�7YN�b(�}�k���R�7Y�%#���.����L�+�b������a�c�Dg�Tt�I����L	r�P�A
4h�6!̥�OKY����6j$����_]�v��F��x���c��D��tVk@	���e�.r��	��L��gs���ٗ�6
�2�'G[GFmӋo�Yk?M5%NQ�xV�H�Z =b���qֳ��(�b�/^Hَ�pB �l��9th�2�rTR���=��Z���nA�']*J���C��ڏxF�����w0["3�cɕ��Z����3��K��\��Tl�Ʈ���kA�j:iM���e��r]���Br{F��ݝd�c����r�E �"�Q/5⫲�aV�e�6h=��l�%Zkn#o��.G)����t̔Y�7jk���`(����@	L���e�s&�k9ʈ]&BͅG�Z%��
����{d�߰�hA�l�̙[ti��TK-�S5nYFaK(X\�ΰ��F�"N8>�m=��b�%�j���Yn�Cw�TeZB6�
�E��_L]J��z"Ak��;+6�&+�9�f�+ϵ��jԀd�tcOc"�Xe�<B�@D]�V��C�)�%m(�F�\�aףh4��(ǓK7��n�d�MC�e@% ��0L�YLGE��^�Z�f�P٬c�b�4��)`�e׎�KE�+h+�ܽ��@2ER�mC[�B��hZ̥H\�Z��.ap��j�6D�,7�ɫ�\�Ʀ?�r_���/��i+6k߳����Ȥ��ır嬼V7�̖�B0�0UѺ
�8�)h����[�䊭Hh(��u��lђ����f��$\�v�d�ٺӃ5�饰�*���
���YY�=�V�0![N��a��,Ǐ0�%�TE"
��*�Y��RKsMT�{��b�&&S
	ۛ�����fZ��ܼ�9D
T*Y�Z+׺���ܸ�;��������Ton�X5u֬T�P�E�ز��&m�"�y�4$F�(i/��u�hܳ�cR(�VFu���J��bnC�rA�
_��L<�@�M�H��nek%[�iU(�ǘk(]��i�P|�iX��:�kE<{6B�ҽ����=�TV�XXd�sm�`�.9f*�]�P���`+��wv &l�uC���:AQsU�js�P|b��cm��F3�A����6.�LSĀF&�u��,h� �9�b�&��8��@轖gd��Լ�{��^��Q��6襕�p���c)�В˰HI*x�c�XUfQ�$��n|�b�VЛ�GZ�`�e�ۢ��:)@�ca�ٛ-��I�s4�Ҙ"4���q&i=�����Gfhи�,ݔ�:[A��F-BC.��J�Z��a]���͒@��Bn�*�� p��.&�@�+^J��n�dh�x>�;����Fѭ1���caQ"���@�`=��oTa"�S����J��l]��^&�dtE�w�P5v�wqD~���
a�b���V�ƕ�T1f���ڂh�r��J:��s��VL�w.�u�n�C[��X�2i����f1Jɉ*�o�m@��9$�(
���}�]��G�_�ס:��P��z� nϓ��c�:#�;.a��݌.Kn��і�;����WK�O��f�:����&��l!F@�3r1�o{��]qNyB��j��ێ=�S���Wi)�bH+�Q<�=����1��׵���at�t�};���������o/�s3o7���X��I�h�,���^�h4:�Zʬ�����m��t��p\����0kK�|�ՙ�pQV�9�땜�4�h�;�a���ZK��k��|s��@c6{��ZB8�r�.��S/�{���������T�W_P-���!��H(�Vc���@e�ˉd�b��(q���o;��<$�3����h3��ckV���궾�c�1�;R�3'��'j���Mu�7�HV��ګk`PU�:���p�=��|�G	������ٸz�ń�ޗq�d �o�)"h̓�`ɽio9W�}#v��%��g� P�� ��}���U��e�5�ݸ�4h���]������]`Ѝ�7Yw}��ծ�HD&t����Ze�1ǹ6غ�Yf�;l x�ŝ�`P\������x�m�*Z��x�y)[=H4��y�2�xzSv�������r��'���9��͢�q�s)ڵ�uvУ�wS]/�3�Q�u����O5�j�g,դs��4p,�ü�>ׁu�IT�+�M�2�}��Z�^���c6�^43���!�WjFs���)Y�Z^�u�&�Dl�:�^_!θ���|�xf�
�*Q�+rl��#��Z�4��[��4�b�p���¡m֚�3^^x�s~��ui��|!�HC$��2l� �@�B	��l$��C��!�����*� T�� �G�ޡi$�l����u�$�uR�`�� T�w�M$62H��M�&2E� *���PT�)��V�z�p��I'�I �I#PX���PQ@VV��*�T��bł�X�V* �X*��Px�AUueTVE�
"�EUQEEb�grb�H��ECQ��&%G�*��,U�E�(�PAb)�����"}h��,A@Db**1X+�0_ԕTլF*"���`����"1T�UPEADTV�"��
*��Q��AQDQH�X�)��

��kZX�����1Y�1E*�9K�F(�DQV"�1X��*+�Z*�Pb���uLPH�u��( �1AX�WL��@QU�
"�**T##5UDH��AH��=��F��b�ib#�(���ĊEUcES)AQ�cU�V�UV&4F
*�(�"
�D�(��-
��"*�E
��"�ъ娏�Qo1QETE�j"�EQU��?Z����F,q�����1QU�)�`�F1W�"(��E"�#�mUF**,X*�b�(��d���*������ �b+��|���b�*(�"�QEF�Z�&/�}V�/Z��U����H:PUTTDE ��G��Eb+U��b3�
�EGL�",�ًUUU鿚�bED����A
�b"""�����EQ�1]�UTEC��b�1��Qb*EX���B�]P����"�*�iUձAb �0^R�MeTQ��`�*"�W-`�_�DH,TU���`�!o5*��kPcQ5J��Y����l,�o
���=�Dj����`��
��(��g���b��
���]}qQ�UU�F��$V'�b�B��(�b���T��`�6�EA(���t����E�|kr��Vd߆����uh�����ą9j*"�����քR1,Qu�cDEF��b�0TKJ*��Q`�z��*���z���51�kDEE�Q��a����E5������X���,*#^�Z"%�*�3抃q�T��""uh0Sm"���r�X+"�L?Z�T�� ���Pf���T\���*��DVz�<h��X���B���f�������(�ӭ��;:7#���מ�����{ �(�((�����V�r�b��h��V�������*(��(��T�EEM2�
��VT�����)m7n����T�i�Hߗ�4������bO�
��a�B�V*����Y˞��6V'�e�O�
���M~�EUT�w��RV*F+u�j$t���ŉ�US-G��骬EbJ�X���j�9��1���:�_�|��������WxU<��/��1"���41c�(�5EX�YU��7K���Q��E=K����QXn�j"1F *:=�j�b[,UD��ut��E�k4�Zc�U��,U�M���: �EAEFҚK֪���h�W�PV,E���kڛui��(�YU�?kZWIUUɝ51E7��С9�ZU��8�y�K*��@���0/-:��+��d�u�#����D� �2�9��UWIU������e*)�F(����*�0f�Pr�"YQLK�MҮ��j����{�uJ:kZ1F1DS��jh]Ҫ)�,����Y����VZTYC-��~�zʻJ���!C��w�Y���c+.�|I$�A'A�@��Q�u��5b �~qAUTΧ�4 �r�4�1JWߵ�Db(�����V+o�(�(e�j�������ڻ�A44��H��DS������é.�~kfZ��P���]�B��k�]���r���U$�H-#�sjG�7gw�و���q_�.�?MDF;�\Y]5Yԗ��Q�\��Q/��MDAPQ�1>Ղ�}�>�Uvպ�iPQf�F6�7C[�.5�1ǉQTNs�Q5K��V�)��MQM}L���r���(ŭz���ѩ�%W�S�Ec}����<�ӿn�|�~~��t©
�TK���܌3e��������4����J��-9�i��PJ�A[��c�}s*"�+s��%Q���N���Q][������ɯoF�j�q�E�|�@���ƺ\ J�x]�� 4GU'����+� ����o����o�:{{�V����K��2'�N�����}M��X�W<j���:����$9مt!X64.@n��'uW��c{�GH�V����l��׸����EƠ�<ܧ쳶�;�jMk��|�.�TDU�yDY�a���T���a�Pժ"���T8£���ڛc�TBڪE�
��;ۿ4Ab��(/YQQ�1y���Y2��%b�Ŀl���r�8�횋>��j����Xq�a�^r⛡rՎ[RWW���o3�����w��x��5,U�Uc�TQE#R��Vj�����{���J*?�*����8��T�QO�p�m�}h#֪#3׹�ةS�1���h��z��SM���``��ں�������H*0[�a���?h���U]2�h,��Ab_n�����ʸ׷[Y[��5�}�@DQX)�����q��*�,Hc�ތ�4rޥ��}����P�a��$\e�T
{���l�Ī�)�UL����]Z�*K�,�T���1��F���'ւ�l�n�6#ur,X��ZTAPo�n�B��e���#�{S~G}����o�U�@>7B�'-kq��X����E|�����6)�T�Vw(��;�H��A����e_�b�k�i�ݪ�:ʿv��*�2�V�V�1��ބ�������c?0۸���.PX\���Yۤ��`�q�؟%b�~B��Z2���1�bS��ݺ�x|> �#�&;��R�#�PP�Q�YR�.�f!FS���u�ߴM"�j�[�UDբ<��4d�����^w�fĸ�i.x\�c��,EX��ك����m+ �p�;����,eIi~jy���&���_~��������~�Wک��!m5��ޙ�g���[�W���[A��aƈ��?562��
��ѡ�^º�닫�L�V��P�a�ֻ�N%B����~�	��wxSVUF�҆r�7�0�����{ƨ��9ur{�����yf³6,��4R��US,4�`i����J��Z;��֔��%����ҽ�;��1��͹߷��E,R�7��Gbp~I�_��Avʈ�쩿�2)�̕�����h�`ZX`�ED�S~&� 4Q�f�#x9Wh�WfVo�4��	-?6� 0~A�놝[+S\��5�fQQ�5fa��c�o�8ͥA-%\��M�簩�R��n���S��+#�~p�.L��&��lK=i��� �i�A!�\%[��F�����~���w���b�P�\O�֨*�Z���t}q������'uc0�_������fZ��|��������3SMek+��}��m����'}�W����Tٴ�h�\_ߎ��b_}��B��� �b��}aw�ۼ~��gp���a��g�C�*R�(�Xg�M'̨)�µ~�3G�Ú�/SFW����GM6e1��Y﵎��F�D]R�8~����n��O�][�~~˺Q�ϲ��b�>��(O(}�a�B��S;�7�1��P��CK1�g��-L,�W,9®i�"���a���y\����)&l�F�U�`��C򵽔Ƶ,+�[*�6D�Y�f�	�v�%3����[x����qb��ܧ 3���-�tCG��Gw'q�T��<)���i�PUFbUH߰̾�+�`T�ˁ�1��R�ΰ�,��뉎�`��3)*)����6"�9��c�a	HK�v�	��'���C"�L�$/�����1USv�����5z��k6���ya�1������n�F�Du����֝�b�3kN��V��:�\�S���8�,�ݡC3�y+1�,��1��c1�3?�
�+W�oA��e����kH�I�=�:~B!�X57�� ��M	z�l� ����PG�:��s��M��y1U^������5J�RT��Le�YUV%�p`���8��઴{��^_�k���;��־:O��F��\f���|�3Y1,�~�E��߷�a�9MU��G��~v�]f��68�*W�6`����bsf��ǑC>�����>����l9�����>ա��Ao0�-z��&,^S��N'�vky\VV���M�n�{��oՐ	"B���8�DRD��,D�u��E���Ns2.�'�}�m7[%-|��k7.,i-m�]D�hj�y��	�6]^R�������6���x�cV"��1a�C2�cw5tf�ɐX+�@W��R gGbŁCA�������$��C!b�JQ���ڽN0_���x�0)0+!�!")���vh��tן\T4����r��湆�v��b&�e{5��X��ZD��H��?$��jI������쭽G���l�	]�4D��v���Z��,˿�3u+\�	��]k�و��<���uh�SY>�$�ů�ـ@�n^�Z(����z�3���
�(Q͡~�rDsۄ?;�>���*l����~e6?4]Z�3��f�[��\��&H($�0�DK-|Iq���ZVZܧ�;t*uӅvg�3ML>���z����u��>�G�=��XV�NW��TP���f�'�\e)���Qӎ�1�̋~�$ �3ѣ�'錘b������_!����p� 1�E�kq��x�)pݼ�+�	���e��zFS̮��ή�,�]��$�or���XS��3n��2_�.�̾ܺ��.�a���;���e��9��PO����$���;w�_ki͋'m�՗	��E��.��Z���ܷtWj{�_�itk«чH�+��:��T�3*�{Z�mEos&ֵ>K�Yi��cYVj�xy׽7*m@�D=Ɵƨ� �/��0���m)c�9�����ݚ3mЍ�~~#�Adl�"0�#������������c�O��Ki�h�P��'��	4Q�(�]��R��,�g>�:�g/�kh�խ�+���� �Md���|ֹ�-��2�uE�^L�#'fwZF�P0	���8�ـ(@(� �ۄ1�a:�Te�w�޹�Hi�_`���f�O�� �$��J=6A:<X���Y���:���ڑ�(@iQ �?_��K�WZH���^�9�]d��|����@�����3�Ȁ �O�%��&Aޱ��Fp��1�(ª�I++u,�p�{����S!4����L�Q&Ka5����I��R����W-t�l�>�ͦ�N҈����Wk�Q{�����U�t)
&��eeo���eܢTsVm�s$��՞K�FΆ�t����#�3�Ct@X��B����T�URfr�)w���PG�⼓���+2bJ�I�
��"��W�P���㯲�;Ng��=G���%��
&���/nOY����&
yQ,�]<J�m=��&�]�g]X7��wz}����6 ϰ���6��7�Ep�j_�k����x%�������h��T~7��%QV��f���ݯ�K���ۢ]\5ۈ���Ѧ�3Z��-4�?!s��f�޳4��шs�὞O��uG����]׎r��g��"D��t����8���%--�^��a���.fMV��\�_'2���3;�Ѭ5���6+�\�D�\�ܐ�M`�J��EP�I\3���H�$ms�~jܠ;5c7�[�;���_
�_΅2�!���膈n �Z�f<`@�'�bڨ��!��m0A#�xd�Dd?�X�C�"E��_]z7�C{��A�j��o�9Å�[h<˸m-�ee�Y�������e�i�M�T#I[-�!���=��M��dM�[�v�ț��N7��\���lsޅ�.�*>�j�� f�)��j#ad�)>�����z�VL����X4ӝ�������chP������a �T��
0�g�D�A�AHA�d<��бU@�n�7?0�Rd�D��Ep�6�;�P�(�:�ULL����tj�V�W�k�kbQ��)K����_i*�8|�b�q�wG��T���KT����T�k������ɑԲ�Ǚ���RJu�S��^����:z!�ӣr���,��/��K(�e�a�7p�")��U�%6vd0�Y#+"���4y3�S�h����J)� �"�|x��v�n���z=���쮙�O���P:S��^Tc
�Q����+?sI3��F�A[�
#Ƌ��B֦�V�U�ԅ-E0��V&7��Ѻ�^�~0����Pу�)��稫k�9� �R���>��g=,X�4�iY��tc�~̞j���r�)�?H{��y���_n,���0��m�^v��[�_�Ji�O��� t�4\�G�����HP��7i�ǌ;85��}��`�otuu���mMDZ+�&�IK��5�4�}6,�D�6�/w�{4+��9A�1~���E�9+_Qp���e��oS>�q��	*H|�	L��*n/�z�̤�DjZh�Z�5����������v��s���� #d� E��]ň	Z�! qPcwު�"���T�a�@��J�e q�������3DK��S�P��~~�>���v�Ѧ:��H[aŽ���"f�����Έ�������gwf��O�S�.?}6���Ά;���b�Ӥ*�����8�W��ǯA�D�ＴK@R�"�4u2$��
	�F�,0�x�S��("���7�L��
<sr苌�R�CyA}�/�'���P�����HC���-9����w�ֹ<��f�&���yO�	�T��"����?�N0$�@ i$ۦ` �$��Hi�s�\I�HhBI]$��a�ٴ �۴�	�B�y	�Bo)d	<�I>{l�&$$����L�|S��?�@�O�I$�H)�H@��d�BI�$H@�c �m �3ׯ묓�A�	�N2�!RHO�BH,�I I��U��荒��i|Ә��{)ҫ A:-7�}K��Q�>��L���GC�]Q*��D%v�D���+t�:;�Wa�y��٫~=^V�6P�'H�Z�����4���-ݕ�T����"�v71ADiy|�\��{� ����n��( }ͳ�
��v��.v��;� :�q����r����ُ��F-7"��N��E	bHE���<�d^\L������	��@V!G�ߘ`1�۾�v��oj6( @3:="�Ca2
��s*bb�������xUl|��m�m�����_a�<��Oʐ���u���߈���Fy�,�ܺ#~���=�̻���GӷD���@�/?��1�S�L!��,%�@����S��9�T���>`Ѣ
�ҝb&���F=֕�^�Z=c��+��-�6�םm�B��͵�F!*��ө�����ȋ��"�xB��qʟ��)Ģx��xR��E�/v,UD������Y����=� 9>0�?���̣dR
���I�pYd6�\��b�!�)�R���8�~���TB@k�<_4�� @D�Z�G�X��e��<1�qSm�\�'����2"�$�+H����x�ȝc�&X�O�DE�:��@ISj�������o��Ws��5�Mm �yUC!o��訃4����A�!�`R�3FB��?=LV��,S	,��GZ*�-PA$�Q ���N�~�|e׸�����<c-5�ܶ�%>�?�7�Q'�d�Y��Z'�X��Z�d<oi�*�����H`P�R�Ǭ��L�[��!/�8֌�H��7}���0m��ʯ���]�W"��X�!�~�UipFF|��;85~������{�CZۘQ�j�'O;�$����mֽ]?��V^}Mj�L�{�� O̒�^}��^2y:�~"����J�u�y1Fߐx���C�W�-jf� �����?}$a V�w!F��I$�a$��Z�}�~��_����{v������?CЌ���.1R�ܽ�Η9��[ʍ.O1Nf��U���n�Ŵ3Uy��6)�����w������}�Z~�!g�	�dD1���

�b�/��3k�t9�A$I<�&�����	
�P}�}a�R1�e���Y`�q����h��_i�i����!'��$���l��$K��D����=Vd��$P�Ddب�q�j$F��}���??7=ȓ)�#Eh{`��*(}��eS�}�����F��k�(U_��+@�fzwe��w�̇_i����B�C,C�Yox9aa/Ɛ�������DRE�����hr$r�ʵſ�7-�e��(m�ʑGA~����`�B��(��Οh��>M��S0�]5V~g����_ْ}��4����_*]�s��*w0���v��;cr�Sm^<#��I$����c1��O�	��h�g�E��X�$!�#P/����"�]��wz�m��e?
;X&���t��k_R�P�(Խ��k�_���um>5-�;W�����4��~�N˹��SU�3 �P!���Dx��O?���H�[�Vs�߫�e�ą��8�~�˒��D ڑ���P�r�&�ے����y��+�*�$w,R� S�
暹a��r��]5iہ'J<p��UB�'I�Rk��5+v��>�,������HJk�s�{K�T�h�����/�M��n;@�+�?=�l������U��k�]�e^�x�-���go��	f��	��**Aʻ�fV(sZ��[՚��]������%Dgm��]����n����y��{�ԯ=���,c�7����zT�ݔ/�+%��u�S#��No>��9����]R�H���e5�d�1����W'qX�3�A���h�(_0E{�!�@{�ݖ����c�z��|���L�ˤH!1x����ѡ�##\M��Z�eL��ވ�#D���m�J�#Rj���|�y@�,ݖ����)�t��{��,-J#��o5��}qRz�|�0++,�BPS��;]S�2�;�;OsjE#�k��<���泪����~d-��@5�~��3��Ę	+��P�y��>[V���@45c�]RAX�;r(��;�)��P+�(	[q$	k}M	Rޢa�������]4�+��뚏j^�?�T�gK��N�Y��-rv�S+���V,�}��ս��az�F�����>b��&9©��6��!��ϔ9�u���2mx�x�f�|��K�з�Թk������ϱ]3S"lHJk�x�@t4�
(y�u�8�[k���>�
�����S�tZg2�.�-�0�قǕ�Xʨ��_-�%��A^���U�7_���_3�zJroךBKOӺ�oo+�9��+Ԩ�Ȳ$��Ƕ�'�4G��q�M `5%F�#S/�4ڻĩf(�==��B�&��S3�dN�d�u�ą��`{	^��%d&w�"7q70~rS�ך����1�G2=)����K�5�{����~W]=z��Am땅ntI]g+��U�'/l�xǦ� eB��6�+%��ӫ�:'��X��]�{��Z])Ӵ�����r��.���KB���J�n/g_N��wӊ��J`�0�]�u�n������%.��B�\�q�C�
��$�l�^�*�HB�QP؊���у��Nʡ}�K�և�aQ������ ߈OBDYe} ��o����0�K�+����Vc*�_�g�n�������u�.�w/�{�:�ɡ��}��Ȝ��	1�W�:��x5�i�_�TH���W9P�����h#j�|��qV���H�{LƆ�_T�~�Nݲ~$R��p<`���%�7�!�f�e�Vm���
���Y���@:�kp�MWޓ��&���`0�ަ~�O�h˓:��"���W���Fj˩���Z��ӏ'�{���*D�`����=~�8�����LGgv0�H�4����V��~^�kc��F`��x6�W�<,����_;����b���әb�N[���c��p{���_��G�Z�]zǮ�3U���p��ϖ WddN �)�;�OqX(��o���]r�\v�נ�-��إG�c����F6��3B��j�����OѨ;�q�$��ȵZ�%u�S�F����J����ğ���S��s�;.��W6�������	Y���@>^�a�D�L�B3ӑs:˷�9�x��Xrт�޾�Gqu*˓w��Ҩ�e���,�3�m���)#6��R��_]��ĕ�����A���*�����wչF����ȵk8�����]tu���̃�G�OHὔ�NT}��q�m��ڲ�m���8�iz�;��ܮ��S}�i૩���h-Z>\b���x��gۧߒ,�h��J��~˽I��B_u���DJܕl�A�Z�aBHT�a�j�=��8��6ǝC��GCV���yR?i2���:}+N�n��ZC��qo���Y�WK���&Ճ��4��v�ս;�T`��:<f�uy���V  ��a��*X=��ݕ�5W�dnT���<�.��
�g�٦P~$z�*�N �z��Щ�!%�7*ݒ�X���z���5������g�Ll����<��}{u���C·�o�+m�+�(�X�����ԑ ���#2�+����9�f�i���~�������<&jǠ�I溱LQ������/�ʳ3l��<����ʪ�r:Sݗ�iD��icç�y��ک�3��;�j���y�ɑ�h2�g�9����?���z"Dcxe{�߳cWy�[�c��]�mU���<�8Q�%/�BM�bC���~�ո��λ��\_/D��wr�7���wV
Cq�T�	�*P��T+֪u��>���`�_��:��E��� ��@TX��L��hwh�A�����
����K�ϛ;aN /�6
��'	���ۣe�(%҈/�T�O.�$��>��.����+��3�.��hL�`�N�h<}"����u\��@ �7��ۏ_"�����39��P��|�_!Ԗ�o��ȩf�i�"�HMՑVV����:�Tv�Z%��ŏ0̀�8~�@�\�]�F��]@I3SňKu#G�U�����v�i�w����UԌ���K�v��n�:ʤG�n�8C�uY��a�])nt-����j<�,�$���oQ�*��:�^;��EG��5H�éƏ����2����=����K-��FeQ9��XR%����{��y�]�f���i�9e�s&H)Њ���3le�M�(f�"f�J�9�62:���vV��x��Y}��Ԭ&-R���T}6���jV�m^��ur�;��.��o ��P�W�7^��㝝Ǭ>���,X;�[!!* �#Orˠ�d�#j�~�Y� '�[�ɍ���X6�ֲ3�ױ��"ru��s{zKmRoaT��c�/"R���
@���}}�r&�,��7Ņ�C�v�T��Z���k�][�+��E�ʒ��>��:���wj�5�JW�'F�F�ڷ�'����Bk+$o���t��V(#�S���T:�X���3uGBͽz�nhB�.|yAk-}��jv.�6�&�Z�m���U�8Q)��u�.��C	�{2� M��9^��������OZ���;��>���ط��W`I�.�E���=�Q�e�@X��m�<�u�$AZf�IEw�r�q�t�ٶkv����Z�mEۧ/ሦ6�`׃9��MS���p� �Y�}3)9�$Ei\�Zy[@��Gv!b\�V�6C�R�w��:��c\�����h�]��0_�vj��}Dj���n�H[�n=�ꇒŵ34��ͻ�7�s�	S�Օ�X��(�*�[YN��`����WYV�͉&*��om�����p���v�`��6��V����J�Z�#w�����k�g�E��hu1��Au�@��`�N>W��\�+���(^8�O�,o	H�a���1���E���L-Ant>-�ǎoV�F��Y!nʍ�)�e���4�NWnnr�Vw�JJV>	�C��R��TC���W��Qnyi&�T�i=�x�T���agHE�r�S�*dunvo�q��&o8�q�W�ޅ�ެ���v��q���]���Z=�L�sg"E��(��l��\IY?����8�S�$�(h����Dt����׎�i��ɦj!���w��`�ưG�
b��z�<3����ҤXk���r��"���� �n_u,��:�b�=���"",�I�>ʘ��cP���6"λd�����c��#&'�wz�&�l(۹��M*��]����{���5kG�#��4��h{����Jϝ&$����]P!��e��xP�bk.dk���#��Hs��w�:�2w�2v�,��D?����Y�R�P1�,��Q?�1"���&	ߩ�RE������6�� �y���HbO�g� �?Y�����&�5Q���<9~�w� ����L�AA`�jh�0H�""3�=��hT<�sԩ��Q���C��h�`�x���h翲kT&�F	�s,D2st�~п{안�c�_�Vh��Р�}�$�A?|k�,z��'��Ǥ���^�~�2F��2@$W�)�H(����~�E��I��k&'�&ٽҦ�._�&������Akw;J��TVE2���܆�8s0I���c�i��N�?!�q 0A#�@G�~��<w���B��"����fd\FO�$}�}�dA�H$\nIQݚ����q4ʊ�H����2|��~N��t@ؗ��YUҭ��y�a��}��O�>�_�=葴G�({b<�:���hڷ�݄�G�AX�����U��n�$���W�:�d)�Bh�����ծ�a��SS��=���M����ƻ�RKk���Dt	��c�V�ves~�Ov�(�F)�|��ԉ��d��FH�# 2ʘ�P~�֜F˱UԻ�)3����){##=hݣ�br~~԰�(b�nȅ���ZjŵR�����2��B���'�{���|�^ӛ�f�S"�����qޱDEzqjpy�����w�v/L�߅�y�C�_�n�뺏�_�
�6���i=����!�Sf�km�f\���##�br�z8ɔ���^�I�tzMjn`��&�8�Q�-��ި�l��u+���8f�!o)��B��h���y�s���4��:e�.!DqR�p��\7����E�pD�Ť1V����������ʐ%��y6���Cg�\X��_�����~�QB�N��}���Z����"yUH^�e/�Dx���H~�yϫIw�Q��u���T���;�"lm�ε��g��t��JS�"U9�r�)�2��%z���E�5��V��'!��\/Lq�� �T��R��c->��(���
��׵-��?<�=3|�}�D�F�L�'zjdz�ɷT~G|ب@����0�~E�Mk��][`�� �J	�Le�f����>�/��[(Lr��)�(��HG_��zI���uV`���*bE��K��˒��o��B%�#X|��Y0��s�M�+ߪжo+9b^�yꃼP�Ɉm4� ����v�u�k�}��(r�z�D#�:�
�f���f�Uð����p�+o���A����}f���B���&���{�kT�j�w9�R���f�<D��0�W�l�]���A�ֲsy��^�o��P�%��Fb��ԫ
Q�>Atͻb�|�U%�6z���{n�7�Z��DV�	��̯:��f)ţ���TD+�e�/K[��$n�u�W�N���5j��\+
X��%�.Z�����lȸn������i���J�/�s�0ow�ڮ��A{�ъR[���PJ�6����7hPN��^����\��ņ~xS��s-�K�{<�l[8�n@BS���B��L�CN��wx3�������W;�I�=���fP������Lv��Ne�N���n<��!{�.Ws8U���I�s�ǲ�S���*�Fr�H�]��֌�j�t�i[�mV��R���j��9h���ِX�?�( ��>ݹ�H�1�Y�CΡ���C|��A�'�������έy�oN��	�԰�T'W���`��~E#wϦ��`4�N�c���ߌ��敏���v�ZB��� �f�̋(D�]T���c�!�÷N)t���ܩɨQGƣ�>Ԧ�W��}$V27�6������
3�?��@���*�$,Kx�Ih5R^�$Mr�U�XGp(��[YOI@ wPAS��@tC�b�{R$Qq�"����� P�"b9����W�ع��Jkۋ
u�[�@� �zn�{�'�pg�8�H�w*��?B_{�"$��C/)�Y[O9Ҷ(b�s3�x@���X32-ǐ�����|�9:� Xފ�0��7S�+��!/N�jjv>�Վ�s?d-����;u��t8�5ϣ�\$}�\�����K��!uFf��U��0D\X�W�q��Q��.�Agzd��T�Ԓ��*UUB!r#v W�c��ܞ��U�ó�ɜ��J�é���E����<v݈�U�EDk���A�?.�ʚ�p�С����3��x���#\׮�:�S���~`��:e1��?i&����몟��>��Q��}u��'���2���w �̓j䩝�3�F���Yu^�V���./�m�|]ڽԮ4��,Is�iT��3�=#����)��W&��F�V�,��;���6��Q�
^���ٝ�U��5:������LԀU�I9r����B�wu�N��M�Ζ��Ѕu�W��du�ݴy+j��MvoS��'1�˖�D
���smR�#-�/�}[r��9
�
S�ջ[ԭV{�
���!�I��5���^���UY�)���6�`�=��U������P��W��2��#�٤̪��\m��Rk��.�sO� ��쇄kc�L��}DJ�pZ����E4�1��_U�*#�:�8~�'�&M��jC΋sI�����e���[�"�:�M�v-��|_�?"�Lf��*Ɩ�|	S �	�l� E�]�\�Lcb(_VC���boގg�zg�a
˵�g�#�_Z� ���m� 3ұtD�Q�Wj�!�0 �T(�XU{Vd�K�語IhB�� ��a�~��A������0���D���|jw�#e3�i@�h�n�:�m����=�\����<����^�3���ϣ#t*	ڃ�%6��;�D��ɶ�
y���=�I\:#M���G0�^���P��y1�`�eb=~�զyw��j��Qr����>#�b0�DG
s���/��I#�����W������4F��.�{_)TO^��D�s�&��a1sM�s{:�}�2I���c��"�G�=SS�BHF"w���r��_D�sDz��ιvw��-�<U���ee8gc٣�D@�,L�RZ������δ���5	 q䁦�&��(@���]a���]�^B����6Uz�!���}_G� �tě�H�oF� �kr�8��c86�v�7`�W(c�a7�7��?����^,��G��z�KX��#啧��o�Ix�U��d��us�WwKn�u��]q�E�f��6g�@zv��Tw��������s���F���5
g�ϔt
wθnp/{8��iִ��0�����&�!����.�e
��Lچ$G*�×��\��G��\�����z�k���dɶ�FΚ��,���(轍��%����.T���j��lАGn���g�O@�:�dA�]Z�����А�N��#ƞ��v��Jx�i!|�p�/��W���go+�̔gA2"M�U*�[q��1'��Ŕ�0l����	y�d�F$��"Ⱥ@Ї�F$�!��I�65^�]a��.�����6��)=N3=9{WM�d��g��ˬ��/�??�pJ�0��x?g��a!�蛒tfG���'�;Y����\��1��u^$C�:���陞�����B�kg��]�- �J�z)R��_TSn�i�d���b�39{�[F�f=��T�~x��o�f��k�P�Į!Мk�:&M�~{�T���+f�L
_cy���"���vW} ������`���,����󸦆ഠA2JR�:c����BL�ߜ���ӷ�Q���}c}#��d�zzV{���a����:Hu+�K��`Mm�}O��(q=�3��Ԕ"vw��s��he���B���DA��\�:5�0�Cf>[�R��:%^���-��8?�֍���ٷ#S˾�3h̼�Ř�	e��z�]��X����Pn���F�H�x)��*�'��ĩ=�Z�=����+��'���w�ƴ�κ#�N���*��~>�"
�ows��f�nSX��b7(i!e�5^X�$y���m�)�sr��a�����ͱ6)Q�K�����v��gr;;��ޛ�l�
�&����f�3�9��Ҝ�{��]�O��KN�8��P�L4+?5φH	�I�_i"�*���V�n��!@�O���g
�P�������L<ˀV6#��]!�<�tH��m7~��&�E���}1o���BJ���4����P"�'.���Ϲ\�։�J��g�'u�S��guF�&��'�F�X�Ϻj�ɳ`�ao�
eԑ������t(�LWY��6�у�@��:Ik$�J �"��f�R��z'�nZ�]�f`!m���'�+������o=�BN���Y�����/=`�]�$�, �5{���hL����e�\��]�$(�̱@����C��6H���e���5���N�r{��0�G�	�^�1+�����
��o���Fس�}���������Ր��$DX���6�+w˜�zBί5�̼�q��q㚷����]pMj�g�?n��}�cG�PA�O���j���Ӟi�[y�����{n��/�y�=2����'|�̢g����s��I��AO�����������90ϊ���h^r�=�w�:�jڡO�4���W�b��b՛⃮+?0��r,�Ei��!�H(i>˳a{�3��AgmWU�����OR=��W��|}�Q�h��OD
4vvUx�ե3�.�.<j:izb^�N-�@0"&"G\A�[#d/<ؤ{Xz�ׁ�"g�r������'��e�tmSU�}`��>��S�Q顃nh!-Wh�Oh���ع�I�_�,��p<eE�����_pf��+�����'Iץ�K��㔲-,�ŝ[6�V�zW;���g����z���+u��������&|�ꖷ�dM�ԫ�\��/�ﳈާ���v'�Rwwn���q͝w��'#�A��肦~�K���S'�*����k��%٥�D/�M�1�F{M��"�UQ"xt�?DV�f�J��xY�<�&�@O&�!<="b��O��"�5\J�ɾ�͇"�ݾ��q��6O`�[~��ɀ�p4��R�8��؃z�\��2' V�ל���D@�Ð�w����Yی�͎����O�$�b�����u�,P���(�g�t�9KG�0�;3U���$�Q�dm��6d�`��[s��G�2�O�H^X�t-9��^n��4n�Tׅl�ޗ4&X���
��$ǣZ#Ï+����UN��\s����THu������F������Ӽe�\�n~�1��ՙ^�A����Z�{Օ"p(�4|$�e<����2ݨ��p�w��-aP�cj��e����?���U��2���H�/2i���ڟiǘ�8�D�5��3���T��Xut��:�����[�M���_�6�Z�V��r����t>裿ӣk5$xrI��A�t91�D����I�7;�8���g�ތ�t�#�V�2e\��?,li����(��Xlұ��U���l��'������WstT��ֈcdL��F�/{���^� �M��r=�!�L����S�����?7��f��['+}qu�q���A_s�+\��͙W-��Wh��Q��=7�ln�݃ � *����Ḣ���Q���;UX��-��"�B� �q��ii,B��el1'#{�Y��Bq����Xokw�vf�U};^��Fҽ���t�7��9w�o[�v�.�]��g����t���:PR}�w��,��޲L�zX�����u1F]��#��2x8�<�B��Co�YE\omX&�6��7cҩ�ͱ�@�tFɊ�v�:qM����/�,Ϲ���W�ϯn��2�6�fȻ�*���{03�]w�c�d���= ��L�@��X�2e�YH,�F�
WL d�T=B(JCh{_*�@]�q� ��c��C��n�M�uz*y�^\a�2͑�.��k2��NX��s�υd��۟U�j[�gw�0���ڝ� ,�� �=�3#��
G��W��W(32(�}��rxY�(1e��>󾾅W����\���3�]�$.���[P��p��^�e�����:4(�.�B�����p��4ܧ�>�}��&U���Tg�[����0�؈�maQU��q'��[���9C�����w���	G~;����z#�D��HtyӉ�AV�j�'����7v��maq~}�k��ՒX ���Z>�c=�يsjq��GÉ�b���D0�|�3E���Fr�k��t\w��ϳ���K��Fl�<Yv��Ċ�����G��a��5�g��������?J���Yu�bȋz6���̷���ON�3]_y�����)z���sJ�r�5w}i�4̚�A�p�r5mS����eI�N>��������VPw� L�z�_l}F9��"�8��;����3.��R�w+>��w%Zئ�=��pU�٠�U�jh�#����DI�σӮ4�=Hf�#�ݖ�!I�.uo��͓)��D�<,WUT�v�#ʇ�=.���/ml�nӏc)l��jN>��NCI��7��7F�-�-���@�:�`�+ݹ����Y����wG���x�1�{uF¸��Q@���J����2r�ED�^^�LZBe<�M��~��Z�L��y���U�־v��?�y��� �R�$O���̯i>��xz�|:��1��p��P3͇��\�*�GdcЗ#;#��ee7�!y���׹?tu��n|<�7�����ӌ�m*�]��ǎk���K�B�w8�'{�M���9��Ǉl)@,D�Cj$��5�rۡj��xu���^�U��y�Jۂ��U:��Iy�s��*Y�Ɖ;5��R�F`�=ڪ?䊐؉E��i:�|�׸_�2+�p��[�Ƚ%3a0)�~�ŭ��]a<c�����m � ��v���ؒ�-�e�y��\ْz�B���p���1���V���Ȫ��{iu*�K�~��b7�kw�I=���)�g\ϙ���5,PԂN�5{��^DeƝ�h�-�A��
�Aa�'�����29��$s�_�hG��U��5�ƈ��u/��n��k���:�ƖԿ}�f- ��-��*����Cwj��n!��<l�=pb'ʬ�d�Nir5��3qR�r��(�@����3Z2����G�D1	9_v.��w�J��0�Ip�Nuq}-�/�;��6l�
��l>�B^��M+��j+*ʜ�%8�D��gd̒��r��g�c����?��N[�s��|}+ͺ<���i�0b��WD�4�/k�ǰE�#Â]�n����A�w���-��8z{ή�e���~��(/}�1�hf�I������vC/.�;�l�7)_DߥC#|���z��O�[�f�j	�R=Q�Bc���b�
g��0��ȷ��k�����Rޞ��|���R�ݐ�į'i��+�8����'��MO�J���Ô��o8X��b2�s�U���#��b"Cױ������k��(���K��y�YT�rF�])lI����[u:�vdۡ[���~�T�B<�2"�|��&v�.2�ǈ2�}}�b�8xUj����O�܏=�s:kf��<y�3]D0��v'�-l��UQ쌄|;PȒ)K�����nzs:o	����d�J�L�K�Z����<�*�8^�w�@��o����fc]B�/F�lM�}�k�9h�.��("�n8�4�`�GQ[
�NZSZ��˅q��y��M��Eѐ��7�~���N����g��K"z���3�6pJ���>m/�Mփ�=�.�wCqC��UNm�~�pV��B#e��a�ۜ�;����n}�2�SZ8�B��ɬ>���eM�'�R��~	��a*�-���$�2�N�B����|5_0�fM���B�q�u���=�MF�]� ���\�:�軈˔kJob��
(�궪�I��i�BPUܖ}tjH*��H���4U��s���u�.f�j�j����� i,#�]��`ʣV�|��8��G5�R;�p�^ۃENN�:x�d2�\ǃ;M�d�Ⱥ"vg*����/���ؼ�+%ܥ��m>�m]�����W.	Q��͐��m˻#0Y��\7�/f�Q��d��.'��U�
s��Mv
�!�����l���m��dl�L�èf����&$�(ɑ��zƘ+�)ܙ��:[Ε���������2���	�NԸ{�sw�#޻�kg�KL,ޫ[(˔x`�Y�[Gxxme���I�o擠�Ġ�{�c�كTK�Zj�<����v3"���]f�k]6��;����h���"��9�vEʺ��9ҳ��x�S,��Ҿ�WV^[�=��]���v:�gs��=Z��n�ڗ�[��`Ӌ5ݾBvP<�%��9�IK��܂6���EM2���ո�4�GW[��o�]�}nB�S����Wm��E̎�\h�Noj�Vq�s��K%��@��S���ns�rŚov�#iSV�7c
����^m0�]��E�Em^SU��v�) ��L�̌őM�����6��R�*j�`��.���dr,4�)���<`.D�h�9��������b�![6�әdm,�r�,��9᮶�+�_���E1PY�^�KB.����C�V�b��G8�Vv��c�cf����r��Y�z�uԋ|�� {rV�0r�[زN�P��h
�Ns��{��xf;U���Z���Н;�^Tf��K���];�q�����}�����}s�%M^��#4-�JM)��[]Ҷ�ε2J���٪���b9ER0;�{�ݩ
��l)��C��	L��%Xp��΢�ޅs�s1�SVsV�p����k
䋶�{;��Ƭ�(A���;ڵ��B������{/M����&8�Yka��z/L�3+:�����<����ڻ��f].�f�J7�p��K�ө�sM�is�xT�JoV+&P@v}Rͫ&f]��;ݵ�"�|��*4P��lm��NR��:CB8%�����]�Ϻ�j�[��z/n>/	��ۧ�k$Y&�f��)�{��%�n#�k"�*���r��Q$�.��l�p�_6OP9�D��6��t�L�$�}2�t�����{�!ʺb��t�62gv�C��/M�c2��rA�v��i��J1��l�,�IZ 5V�u��s�n����{��[]Y��x�Қ k���Ŵg�jг��0	���vQ|C)�5�:
��[�\Wh��
�D�����Թ�_.��K�ɂ�%ĥq��4(�9�gn�&֪!��]��  ���Н��.��jS'`��	Qv"b{$+��gb1�]�`<���cz�JQMd�`���9���ά�+
T��[^F��=q�l��<�ꊓ��N��<�٣��6$� ��UF��.��Jz�~�ɯ	o���ED����o�\�s6���d���vuQ�������à��A�{�����&Lt@�5�O�f��[��U<�ٗЃiY�r�y7����J��.�u�,���'5��p`����;���M��=Ǳ���W^�������nv�a����;i�V��3�㧷�7\�+�5j��Ͷyd?Fn'c8G8~�����$�P�S���K����]P�J�v�e
�N��i�0���D�/�O�.DD��v[,e���܏v�T���N`�AB�ݙTsD�e��G�6�@�&	��\Ө��3�6-���aDK�q����^3�u���6m�^�4�L0�|{�>_Q�Phl�Tx�NN
�Z��ȭ,F���=�zrf�S]9�%��_+��G7����J�/�(��3�Z��f�r�?"0�p����C�Qը�&/�2��v^�"	7Wf)�>���9��P��/�<m��S��@|Ӷ
f@m�kk���0H,zʫ��(��v��+-ͬ��v������Q@���3�{Q�eD��3(�w0B��?3޽^���=�����v�p�^��������m���ǻ���m�qǵ�B�rj��z����.��s�;����k��8!����Z�Q0��ӺŖ�u���W�u+,Qا�7��3PZ�>խwGA��7/m��޽,��p�(����7���nȣM�F�SYYO'���=�c��1U��*�^Q�ڜ�A��.�ё�;��L[���;�(�8WDV?p�_j����A�����m��Q�w6dw��{��u&��ɥJ6:��<&�W�:~��yL砌>y�`fX��G|����܇�?^o�����.x���Cv��a���4�	o�5}���!VP�)?;�3}-�c�r��+����>���#�Y��P��ft��{�����Ř�e8�uMR���wt��/�&�*�%�f�Jrbb��\3�5lU��s�s;�JQ�ٯ�ά�=���]��>�9:�as���;jfJ3J����������~s�[ƾ>���G���y8nOG�:	�UH�
�̂P���Ԧvō7dᙊ{��f�s��M������Q���Í=�ΐ����).V^������$�^I���><=Ͼ!ey%~����
P���fO�{=�kf���Fc�������B�̮�=��rD�~�O�R�J�ˁ��3}Bݝ�l�zz��%e���σ���Տ٤nPTfkI�Vț�(���Bƈc�ݿY���y@��eiw<�Ȭ���ֽ�_����1�*_ށQ�����cK=��_|���c���M%�!e��^����V���K�Y}v�����u �ޙ��;�ch�T������B��!ڗK�q
&n�w��7+B3{�-�xf!V�}�����rw5�G]p�ƉO��������z:�%8�?3��w:����L�A��ys��&�~�p���S�M
�^s7�E,]v=ƟE�����QU��.������+ޏe\@���Dt�L�o�y�7"�z.D�P�m|>ƪ�^��^(�28�V�W>�29��Z�*J҇�&EQ��Ѳ�iF9wU(�7/n����C��|o�ꜳ�����ނ~ɯ.[���Q� S��S�z&r?3YF%!��uL�{��/�����c�]�ʇ�z2����$ӤœT���H���:�6Y;�Y��(�Tt����+���5#��;��e�����L������=��+����q6j��T�D�����^���֨��L�
� \�p]�W�⇏rn�*�.�񙘍k�G��[�6B!�FJY���X�ǌxcwS�L�r> �C>�pl�-�㔥�������<��UK�lLdؾ~����� �����!z0��V���b��3O�#�:u�~��|#w=���g�?LK<��Ȩ���0��*�rx����N�l�
uuG҇;F�N��F��"du����c�{-�d�8�����O�B��2��G���&^�M%������'���m��ʮAwѴs�c��[�/��Pgo~�-�UC�&��7��W��U�ξ���>�	�](�g�GY�ۧ/@����t�;)lYot���V��w�y�vqJ�-���]qY�X�gn%;Usk�yo����.뷝�����k\�Kk���v�^����*|G>Xe�o�
yo�en���N�B[���k�kA��V�o	��ZG#� CL_���J��&���r3�B�q�+/2�,�[�aeN�ި�A�I�����Ζ����B��^S�<\YEM'�_���|L�	�?��B��͞��(��5��{ER�*�����n�A�:ܦ:j��sY��{��CO�Mf��w0B|������:���`�����6�L��F��61�^����]|h5;��B������Z��s�1�F�x����n�Z�������5�?��5ȉ�d�_Ƿ��B1H׻����Dͯ40��&�Wċ>���X��W�}��dRd�BM�:�Mς��J�%����#3��߮aw�G�	z���.���]}�W���C��Ƙ8u�k��1M��Z��8��@���}J�f�q ���S����7ͣ��t��O!���O�h��=�_�>B�*�#㢵��t��,FUt��b��6ة�h/y��S=̅P -�U,C��{�H:��-����YL�Cº�a�����"��ލn�m��`�ò�4��9;~>�.��+���]��#�,�s�7AZ���]��R���l�ܪ�R6%e���1)�� ��I�.�#�/�ĸ�L_�YU��qU2$��t�t��[
�3@��6WVS�^=�ڞ��v7��p,��η�y�n���B�f[���fG�1���Œ����uڃ�C�pG�M����)q�|n�)c&���x���:��g��!62lJci7o;8<��i��:�+��޲��n�̶n��(8�!��Z������3��l�a�F�|�F}!�Tr{sS�R\Uw�p8?z(
�޲�/��5JS�.~�\C�\i��28�N�D����c��>�ꬓ��o}�΍�i�؀}訒�ɒ��,�k���:f��?<��[׊DguJ2����r�]W���i��9�6Thc�4���pO[�QJ�]�D�۝-�-!c1���[�x��x�cX������������uʔQ�3T�9�`�VY>��V�;EOg&zKT.H%��Hת��V_N�I������.��٪ɑ�y�B��}�1�C�Z�~?m���r&h5uވxgf&�ު/C����QëG�н����A%��@1�v$HV6D��TJ�������1s�[O�����کW_Kª����h��a��u�ˎ�8��Jho��~�K�:��kC�s͚I�=gS���C�M�?��7(���[&7����~�؊]�(S� �vL�#�Tq�&����5�b����>p/���*�HX���2/�S��^�w"P��ɂ��z�+�̢]k��9/]��<�_���u/s�f���r��\��F�ģ��Qz1�CY���iUk��M�փ{BT;8 1G++����d��
���c:�m��A9��jz'U�os�f_7�ϲir�t��P+[ᦧ��"n�;�C.�"ξ�K���vx����?އ|�U�w�yi9�:�cZ��/g�3t��O��8�|� �s�riTH:?*|��a��x5,��>��W-7<$f^�?8~� �,�éaIO�B�y����/ʶ����������`�*���Gnv<=u�#�w��$�"N9�O��C�1.shW�9�pw���򺓢�
�_\D'f��T5��rF����t��̨E���1R[֒��xs��$��#qs>ȃ���F�l_��X��a�fw��Q˸�Ϲ�٪�<��{g�I�h$�¥�񝎥$��$�����a��W���E}�\i��=+o��"�t�\o)��Qa�Q�a	��F�,ꝣT���R�g{�o�wkzj4{nn�-��߁/����w��M6R�B�3\�"�MBj5����j�`�`pSP�,��/v� <˩៍�B��B�TE���瀈`�Ț�hтmǶ5I��8d�0��W�&V��1��!�>�/e�ʪ��ez<���.����X��%ťL�]{0�����)"�n��Z"�'+�����v&&/�Y�&�ZD^�P"|��f������٭�J��>dVw��O%X�W��;`=$�Tsc*��XX�a�ji��_S��|�o�:P��A�i���K�v��v��#S�̅��g�cm��)^�I�$��%�Gvk��OT甭��U��p�W%�)`�A���+��NK��E{SU�f����t���p�5L�,�I��7~&W�{z�?N�T���v:�h��q����˝Ӑw�$A���XoC�z ِ�t��=��B�w97a�Z��wS�{��TƙSU�=.z�]ssy	��[�}�Q��ꟄdF��(+����o�aIXLr��r��muA��z��L��.Ϸ��!���#9p��a�U8���O�q�ԁdiLt�oU��Aҏ�������jw�'�K��]qD=	F>��E�C��;��oY\�G���;�i,����x�?Ύ��»$�˽�u�
��4p�=&gG�O{�@/�.��x9�u�ĸ=����U�+�nۄ'A|s}»��<3�J��i���{��0ͪ�!������L;G�*S���*�ʷ�z%z�rzf	�3=x2{�֜��`�>)dq���܀~��[��8�S*�p�+�k�׆�r�A���-b�5��Yn:�cٛU
�ߣj(�1��=&Wz��z'5�^<���E�_�#|����}v�Q�W���[�>�vP��>ԫ��bL��O"�v)�r���C�f�ߴ��/��n�luOmL�Y|�5J�^�.&��ϣ��>Ku���>���[�Zct?UUHG����L�85������I_Q��.�X�B���Q�C#��NSl|����O^0���W7d��s,�1d��ioz.\3~,vc�Ry�Yk>�J��0T����/HyI�]5��v��%���N�N�;��+�FsG`�Sz�;�������A��vqdM�M�(G�W��]�Ǝl�0���f[X�c�ګ��-C���iP���hGs��xOGګ������;5ןedy+�|̓����zT[*�`I�G��(���S3b���8V�D�ةu��Q�x%�pok��)���� ���y���oܬ81v��</{��"��t�r|ⶄJ�2�ȓވ�ט)�+3¥b��������\�Y~��"���]m`#��C�H���ӣ3�w2+����o:&�bJ��mr�����4br)Hs��G7��(����e��|���Տb\^ɺ1+To����mа��B��ӝWcW8S�ʀ&ӃN���5R��~8v����b��8U�/]Hz�A�H��=4%��_I�7�p{�8~�90����ey43�L�1�}~���p�>���>����a*yB{�:L�����������(����d�H��QE'�����?G�<u�PD�8��K���L��(F,ƃ����G\`�.NhHAьϝNh�H��f5�=���J`tY[ک@���b`1ױ�c��t�՞6
�y�Km�΄B����Hd')gD�w����s*�ROY��<U���⫴LN-���q��ۼ|�����j6�&Xƻ�-���NYt�E{.ۧ�N"��f�mj���1"ԃ�n��L9oew���Z��>���i��N�GQM��g�t/U�H��_VH�U���.��P��|&bx��9Tj9o�|�Ǵ\u�6�~��*�y*^�X�����>w��t��p�Q�0$����I�I(�N� N%�i����	��1WQ�^W��.&B%�u��:�Fl�s��Lp��J�
��XG<�>�1	(�C�IՎ�@�S�n(��&��O����e��B�Ŷ$�f4�>�j��NH�
�t�-1�����<ʮ5U�j�S���m�e�+&*s�9|��/�]�ex���(�v얡��_,��I>��kwuG;]6*���WJ�y_[�\]_CF���f�0줼�:e�ʑ.�M؁����s�of��͞�z�LF��>�q���-"��/W?�t�t���53��r}�++brwѴ�w����}\Pn���^�{��\|�u��.cؿz)f	��W�1=�H��[�[�ß.>���ׁ�0�[�������{!\���g�f3��;��B�����u���.�M��~y��>�s|r�{���p��bf�c ��{�B/� ��oF�@lW����<�u�/�[ϭ�g��}�~����N�㺻�jj�~����zϱ��!'�ҫ>���S�Y]�u's�د��WV��*Yu{6��̈́3J84��z�� w��q̎%��<�Z\�o��qk�Z#�Y�S��A}|6�8_h=v^�"\��A�C�?%�讼�u�ۇ�B�{��7�#��b���>���~�4�L�G��**���#q��lU���Y��t��$6��ӞFO�	�O_�%:����f8����W޹2F�6���7c�����g�ǲ�ʥ�9n��}�"�b��>8������`�g�l,��#j�D`$���Z
�jq��+E/@�M"r������VXn�s��.k0���f]�)�,�hI���|�9>�>���=d=�
N{�w�𼰧p�uoS$��3�.3s�3{�������8ln�S������xt뾫���z�X��z�K8��~Y�����p��[�E���85jK��G �qz�O�hU��ٗ����[��!��l�����=�7>�9Fb#GUR�1�!zl��+�x��t����f�6�w��U��#èPsb��Ha�[C�+T�wS����y��ؽ^��~�/Lk�Jv�
����N8��
+.& ��	�� ��l=�,�a��o=�f�AGu�3y�VTr��̈��ާ"q�1����Qަck�%$f�RC[������
��{5;+/Fʲ.�vOW�0�o������MVI0�c\��cE��R7֫��68+�:�\�����_,�:9�3��w$@�e�֪��FMB���PAb�� �0�<�j�R�{ܩd좵3��δ%"0a1V=���������L��̆uXy��4�mÉ�j^u�����I�fJO]R��6r�fj��6]��Q��7���;��(�*:���-���U��̝؟]*x�E霡/��Sؗ��YrU���J'g<�[�-�s�'5�Yu��K��|����ۤ�h��:��k�>U>����Tr}_F�@�%��N�o���9;ޘm�}������B�i��CA�C4���b.,'�J!�#��Q�I�Σ��Ӵ��{9��j&�_��˺�<7f7�f�4'&�*�Т�"��8\���5ѝ��M��j˛�Y�N�G��0K`5�GZ��v�Z_��p�t�ԣk�B'jݠ�q��y b<�-}���z�X����z���H\�Z�V��88��f:)�_M\3��
\c#�ߔ����ϧ*巜m�A��1�@�)�Q*��W��0nc�w������U���9+�x�y����kWAN��Je�Y����&l ڻXE̼����<��B���x��ƟpA.5�͍�X��ـEG�ۏ���p�ʍ�� .3:��Ρ{`.��4%��f�Fbr�<���@Y��Y�u��@�ˮ�	={R'Y���/�(y�{38�K] ����X���%�#��A�4|��ڌ�;���D$��l;r�w���;qE �G(\�oPf�����M][��hVR;�-9ɦ,�*j��m�Y���X���ئ��C�jot��cvU�J*c�BՔ��S��}�W�$�H�#����n�.c�;N5Yl7��u��MNS�9ƺ��j���ˉ1Vn5��C�ƨ��C�8Ӭ-�K�c�؜V�Tzi|%�:Z� ��X;���w�qj�uj����.pାkk8�[ɧWF�%N�yXp�`�+9h��:��+��P��#���F�* ��dR�Bro8Ұ�X�3�W@����)Ǌ��bާ�޻����.Um� VUj�Y}׌�V	jаj������
7�&@���v�2�bcm鮹5e=�2��g:���v�i�������B����yC�gGp�T��P��w;�S�\sfţ��؆�wRN�16{��J]>��k��-�Dm�s��d݁���[n��t��G��p�LV�����ܻr�xz������ĺ��1m�ua�r�`8{��q�3i�w�.�C�S6򭊖JO�yf�MCJ�ɕp\ޜ5��8A��[�Mn�!��;���y�e�o9��ץ��N����-)��]c���l����Lzh��^�-�Z�fn��{ufR]N!�pD��`z-"V����'�}�UW����G��k��|1�7.PH�n`��o�P�����q�;:�ݥ%��@�����c{iB�ـ�V���$�j��k�y{q��a�(�ؘ�b/�7��\ǳ�#ǿe�Gf�voiPL�Y�QZ�_���y:$�C���ϳ�g&�3n�rM��N��<b��r^]ǎ).o����J�t_�@苮{��_�r(�V�τi&`��}��}>b�wQ�G=��hm�u����&�me�@��4W���B�-�Q����?nK���E
�,ꗗ�6��~��u���#d���=Y��Y����[�&4��"5�W�pC~I8��~�Z�� �m>�VGFȽ]k�|�9D�р�Ek�㨙�ou�Tȑ	d��fI��k��������,�~y�Ҧ����l8���r��{
{u����C��32hxիh�d>]�-}�f�h�![�Ou3� �fzv�W#���z*=x��N*�v��yI{t�?Y��|��W%��k�������
&`gT��RZ��,O·���x�I���teF����>�;*��7a��y�U.Gzk�i�������k�4���W��4>J́��;Uj�6-j����W���	�����cKt�]T�ћ�i��qʬ�r�G�1������4�d���e�Yi�K�!1��%n��m{�M��L�,l0ON�\��=ǧL�W�����3L9y�ۜ���쥱����q3>��o<<���7h���4�8���g�i�(�x�nb�Ǯ�=U��WIw�=�@�+� 4ל�SؤΣE��a|�S�KvQ9��7�,��<��9�3�և���1y�g�[�u����^q���%g����_�s�Č�RV�Jզ�����}=�}eb��n�1��hx�X���`1�Mt�E[D�M:�R��5�׀C���{�lq��"����ӕvx��s����1���<?L�����
ʱ̫�m_ޝ���6w�S7���3�-���꯷3�����BJ���LMʈ�M�J�[�����*,ޕn������U�Wln��м�[^���ݨ�V�ۂ
A�����%�W��&k�p�NӬ�l{�e�Vn���~����s��gi.d�W4�F奂�_���]Z��e�����Tj�/�ia��&-��!;LE��b8�$�/o�:[��%�,��;0��N��9�[=�6S�h��c�[��ͤ�Q����q�;1}�􎻓��e+�:��KW*��o(=���Bv9ۢ�_@���Yԙ2�t0�4��ɻc�{��Q��B�NY�3E�qG�+L�N�W�tf�*n��ׯ��Y"�p�4�L*S'ux��Y��0g_��O���	^�
��N�hs���!%~ȮT�MU#N��NxVc�dӾ��g�f`�k�:�Z�/xWQ�D*�|09�}^��ǆ/26�9D�~���c*�>-��AuW_a�!5�jD<K������cw�����sW��j���|��p=q�U|�$�-����n*DȊo#¼P�A��Lփ��m��߄0���׭W����r��b|B��x/�Ά�r�+({�zZ�yڮT��DXO'��{j5㠴2���D�W�ٱM։���R0n�c��~]L�jBd�-�t��ő�V�b"0M�OD��ǯf g
��>���O%�xk�:ŧ����hWf��nN���9YW]�^@2��5�x��v�!ꋆ��^�5�7 I]�r��aĭn�`6�q�=�)%@Z�����D�����'��2�b�d��b�O{8R��+��V}�L��l�9�ҼU�� /��](��}�v8N1���k����A��Q��zN���)	��ǗQ��Xy1j}�@����̆��00R1 g.�q
����m|����H
V�wk[ύG �Z�_��Sy�
xN�3���h�;=�%����P�;N�I���Ι�����-�wq��N�B5�b�&�}�j��4�0������\l���-�c<
�v~ �:���,A��c[���Ǭ7ܻ1�f���n~��,�^�Qӟzv� ����˜{2�^��X�]N4�J�5{P��ȺS�h��s���0��ɍ�W�Z��n�?=��2�_��oz=�����nieZ����Ʒ�|�*r�8��F���L��>�Lv(�w��T7&�suT��x5�J�2�r�F&9���"=��sli�A���_
��닣;}�7�9Vg�/ �G����A�9���!��^�r�6/E��P�Hy7׃&c��1�A��Y#(ӆ�>AC�C�|vRB��ub�h��=$��l��v����-{�[���"v'(/|�/��t�m��jb�m=����f���Gb�>�2'`��
��_<���V�=�`�+!�CAz�奊�1�P:8r2��)m���/� f���2�>���)R�Ak�NVm.�|F���{��܏�hp����B�.
�v�e�9|0>�9+5��t\��jv�޷�U�o[�v,��U����n���h��u���b������ ��Mi����S_^v�p���:ξ2�w���rC�6��6�_۞�R���s5n���4�]��p�iه�
�c+����<p?��X����RW�粒h^���{�m��kƐ�=E�j�֢ !^HQ�Q��zF�?k^ɛˬ�yLz�"BoP���+�Y�\7ߩ;�K�t�F���܄��q����}˦��@/vC�ێ�eݿTs�f�����s������)@�ٻYBK"�J��K��M��3~���mM?{]E����w�9� ��Z"���Y��,{+��μ.��z�G���q���Y5��z�֨]�<�9�EQ����lnj���6L	�7\"^��%t��V�j�?}��f�ӱ|D�e���4=�C�Z�����_����=շ�ң�N�n����
����`��'3�E�6y8�#�L�9 X4�Ww�G"n*�n!U+�U^s7�@bgxb>�&=�s�����Ix���S��3�M��Tc)�Ek/��[��ټ�n٤c4gv>�)b}���.��T�u�ۑ�S/>��rg�+Z�B��L>��e�AjS�Υ\
�ZlK��
$��vV��8������Xﶀ�G�:¦K��0t؞ݵ��[���ɶ���sN�&�������[Y��म�[4�2$�<Rȩ����P��|�>i�Y�6��3\�6��7t��X����)�_��qr_Ώ�l��r+�Q��u}�:��׺~�Ǒ�*�l:��C:��T'����˗���m{�eF_����?k�W9ۇ����n����	�{�0}_��7�p��L�"�-kJ�Wˇ'IV��5g������}�G����Y-N��=E�
�9�`��i�Wf����Cu��|�6�|��{��qp"�]3�CDx�m~^�UK�9�4\��wq�??e�m9b��T�;���$�K�����tLrO������C �K�%y�T��_�;�pm�q��h|'=C�8��cs$ur/8M�E��.F\�/�a������F��X��K;:�1y�Ʊ7�MU]ޜ�܆�o1��	���\/m<"[]x4��)��X*��1*p��;٩��V�8���E��x�W��"MyJ�{�VГ���vE}�^����TH@�y�v(kF�y�*Ċ�z�u+�ƣ�C"�����ը�����{��6m �	$3���д�ź ���@�\��	�mΕϦ.��)t�f��N��+��c ��g��kr���z���rRO�e])[��}���><�J�����+�>?���� pe��x���w���}Z_�	3�ϼw��mS5uoz��.)ߗ�7���(9�d�s�wTnoK�=v�a������`��f���^�!_rЫ�wp_P7�J��mh8��N�N��Q��9lP�r�/�A���B���j�m���^e(���"6���qgz�C��>�-��fa�7w''��\f�hJ�	Q�M�I;�(eRܢ1z���O��&,��>�ͱ����6j��w�����"�2�$�l��~�Z^��l�x"���ݠ���oum甡��O��������ͦ��[�l�dL";�SN�z���QY���tU��<K�ƍ�!�u:R�l���5�.6��o�<>q韶z����E�;��Ϣϐ�h����f��d�F���X���'���tn��6�E�܏d��[Ie�Fj�Y�Ii
Ecx���n��r*���ع~����R��ɷ��E''�a{eP"�����v�9$�vҥ2�Z4�ֻ���+2Yt�F�
jۍx�n�6�5ʓT6��,g���k:�l�
v��]�>ζDA2_Z�k�u�����(�Jw�Ȕ9/�{h�nm�_�#:�"׼椂��'�ʊXfb�)�>��pF^!_<]ْ3;آ�=�K��v�#����Wv��;6��7jĖ�l��%�??���<�վ��³��_��px�{��a��:dJ;�v�YuE�P6<�o^e�yOp�Qy��u2<��{dc�AB���D\`��{��	B"i��18Q���i<���*�c�7��z��2�h@#%UL�H1鴫��>�C��}vm����{5֢}WY�&%�qgճ�V_Vqˡ��hX��������t��^?�������=���͈hzg&l����v����� $��}ƬW�&�'6�x�wѺE�LK��m�W�o"3|\��P��.aѫf�Q��<ġ�H�#���&����>���E��^+9ے2�A�9}�;�w��c��_��]/�K�>���Q�o#0�����N^l0���{�*�����7�+9�Z���z��hGοL{�{�X7��Z�,ef�."��3�̧ �]�ҡ{���iX��|�Iu��E.�YEj�6�v�Q!�4�-t6��7�U\�s�5�u:�t����'*���/U�3HS.4f��A�ĳh+�$�V�5�һ�����o'J���:-��o���rv��r1u��M�ԡ�gtjd)�)E�g�]�鹾��4���t�dz[׃�@���a�{�&b&&~�����yx�o��R.!`�}�Y��Z���T�`1���Ͻ��I���(l7�v����GF��=߰Q���u��bJ��g{P�G�c�U�Dk����5�������7B25/���d��v:3��]���$V����v^�
aƓU�Y���p��k;fOEA�!���2Aݿ{5�ڤ�C][jb�8 8O�B�"v}.��ӽ��*�Xd��P��Ev���dƜ�I�&L�y��S���`Q�_�26��5�y����uT��߲���A^�!�đ�k����g׶�*.]-L�3)�;����D��2���D{T��G��S(gz�ŷ3�[�Û;էT:���vZk��CY�V�k�/�v�I�o,Dz
Y���*MJ؊�N=�*ɁRb��y�
c�K����4���C7�$Ѭػ�3���=��rw3Y�\��g2p�Z�p�.��y�WD���6�մZ��&���b���m*n+�t��Q�����R�r��;���2�����m�Y���@]]�����Y;���8no+I���,�`�ڎk�Htr�E��>��!���7������|��3�*ϱ�β� g.F�@�F�����_H��#VS��󬝌�tQ�g>yLX��ɭ���wӊ��]�|�g
�"�.�g�ѽ�A��19��z��Ϝ�c�$�T,;H���������x�}շ�/ԵULh�q��&`y�VTE��DɯMMa���z5�y,I�?�N7�@��1���o��c,y�8�:E�}U�˚�y����Ży/��yp����TȲFO/�Gv�k�rԣ�J:���\S[M��}�<4�Wp�=�P���K�����VT�~w����=�-��Z�A�����;/���ػؚ3j�B���q�Fo����E�mu�*���N����9�����\_��i4+�{y�;k�]b���p�Ô|]�sQ�i4`�tW�'��Ug�;��a�+{(KQ���G�:�}��qVr�b"^\"��]ӥT<���9=Ma\ +{/����gu.���Rb�Q�#�ύ�I1 ��W==���C�ά&���lry~R[��W=�w>����sP��T�e%�װ�s-ۼ��i�B�2���ֱ�mҔqD�f|w�0!��k{V�p�K]s_mb��)]��{���n��n=��=�ԫ�#��u'��ɪ����VJ`R�n+9V�.�F�U�x�%Ŭ�0*�Y|(��5�_>/�44���+���2�4�%b��l�R�X�+��X+� 
���0p͜�f�2+x��k���ap/ +,:ь��9]�u+��$>�{&�t�D�Q�o"Ὣ�*�W�ը�AoɊ�n�U8�7ՓiŨ�9�q��%Մ����;�F[�1=^EKn\ޥ��˺��[�WpH��&kZ��8)/�2^Ն�Q�
�鮮�U�f�)�mf�K�٧�V=S�r�`jt�{:�X/�n�����CX�J��f�����^�s�	��f��!�^��|��8&Rf0�3�*�Nr��!�٬�A�N���N�[�nfWA��S�����٣,v�L���%�T��z����yC7OgT�p�O���՚/EمN#��i�t�F�)�s������o$��n�(9�������mKB������i3�ց���������J�h�HSj�Ob{����Sr��6)Ήһ���Ӻ_oSݡskf��i���e���qʎ�Ʋ�'z���f�V����}y+
\*ۉ��Eu5u��оV_+��{�K }%�ۀ#*b�OF3&V:�u�_q�f��S�Z�7�m>�F���ѮvQ���BkF"�D�u��j�wڮd��B^N���
M��d�|�f`�@Sj�o˘-��֑�����q�k�(S�q�ǅJ�'!ұ��z3�q�'�s���.��k�A�S�{xɒ��q7�몀#�èU��?���t"�J�m�L�,B;2�;�o�k�:F�.��8��a��W�/a�)Q3��}CB�J�ë�%���v����ʹ���}"��	���%�r�<�:��`�FT���������X�嫨j�����w7�� �qT=�WK�@����+i[44�_R{�"�}�:���j�elh����ku����pS���n'�R��3_3���ͧ����"ɓx$]�Y�I�߽��<�.�Ճ���J�t��,�H0��N�x�mb,�W�ҳ+QΩ��Lif�z3uc��/���y����X��t�:���5������IE7l����b�_�@ֽ�����ȯx���6���>H��ds\��S�>��734� ��\�܎����ͧ/s�=_ uGe�<}&��ta���Q�k��l�,�䷍e��ǜ(eg���j��nw>U�>CQ)Kݧ�t��眔���F`�um���6I���ց��~_ �:ޙx	�]w�����;�d�b�P�EM��N�s�[�9�+t��5�G.��l��	C��S����$�*mf�d��.����	e +v����a��n��)7�u\����B[��[Wf�ݽ���x�ou�0���z��X��m���I_�4��Tg^z"ث�5J<q��VC���=��U�f��i?`���AQ�`��]�[��T?��9T,�p]��g:��P�I���=�f�\B����k{{׾�&����c����[~(��خe�['�ϧ��4~ߌ�ٍ�� i���]W����2J�s��e��3�[�'�V��o5�f���g0�|�z�Lʤ�=�3�k�dLwB�>[��yYW'���H.ady�>���\FƛW�{�>�k���+?G�2"���(����q�|��$�o�n��O�G;c����u�hl	�螟z�����O�zDI{$��cw������vsb/�����o&�9�{�9�{#i������m�� %�b)Xhi�9���z���>:�{~(���˞�}��yXn*��Kfzoq���~E�,5�"�+�������N�s�{�~��}���XѾu.�{j�)�|;��C�s
�.�X!R��S@����
��Wb�v ��1�h���FR�skR�U�;�\u�q�2�8]�3n�;�5��L�k,�1Ð[C{�Esb��uҧG$��9D��	l>�vU>��H�H�.�i�����S�+pR�w��T�j��b�ۘE��w�7-��4'�]茶x�(��ΐ_���G���_�A�rvq][�ͥ��{1vu<׌�*++b��qOA|�ntY"�AF��d��T�[���"/�c�s9����n��4��V��́Vr|!8@���6*���/݀�2��'ü=\l�)ntO��̜�>��u�s7L��[ɥJ��y��b6�I�d;������,�� ��*��Ѿ�Jc�iD���Y�����M�KV�ӻ��^ÅǷ9Zi�y�9s����|7����;�#={}���[���^7���]���mCq��A�\^�R����ח���1��������"��}��_nXY��7��{~�]y@ƿ`�s;�#1��+O��F�����c�¼*�Cg�if��w����/A۝�Ӯ����!Hj����2��qD}66�M�v�#�N��ɻv6ǈ"ˈ{�pG�y9����
�u޷���Q����v*f IR��)^W�ӚV��W��˱.ڂ�l4sD�o1n��9��Sg<�ʶ�)Y������-�A�5n>D2i������9��1���G�M�A���VJ�s��:x�k=����'�A��>B�=�H˷����򩭃u\�c�]�f+�0Z�ȁu|2qε�W`�ĿA��0o,qn���'Lx�:u�;z�����Sgq�^�ϟ�&�]�hG��YU���8{	J��&�DU��l�+�"�J{D�¦���O��,з���{�O3�3��qJ|�}�د�}�W�dw��7���ōۨ
/.�ܢ7m�3=�r2C��nqB�:�����H-��Q1���Q�N�+0���J�x�o%�h;���ц�J�o��/�8�S���X��mz�>���*8��y�.53�݋:�����95�$G������v��}v;�YV�b�U!K%M���%J�UX�+;�sf5����ڹn�����TSͥk�^�'S�;^��1�s<p���+k��0H'��p�/���dژ�d���A��nk�L������6+<1��\s���nGnPK�۳�H>�p7��^^({��XG�<f-�g�3%{O>�tI�}��"4C�<�i������ĩ�=�g����8���{�ti�^#��b�ڏ]p��@q�G�gp����C]�X9����F�a�}]�Y��|Hz�!�z��s���F�Ψ���Ca ���]�[�ي��4��;�mî��wm���3�TF⚷�#D�^g���H��&���,������o�8M��˼���M�q�����f�b=2�����8ԛ�&FU�m#�r!���:�ݟmlwz^�n4=�/��1>5�g9�/(3G���w@q��DǽJ^'�����i~I.Q����ǀ� ��o�ѽ����OF�L��L&��L�e����lw��(���[tm/xo{����Խ��)k,=7�cՑ�}�[W\c�Ys���e��HY��c:�Cu8Gc���ݪBNT^�X��!��Q���J�B+�޿9�g������@�[��*���}$Ft�s�K2��D��# n���;ND&��0'jq��&�ݣ��̚��&����hWst��fƲ37�.#R^�����l{�-��@��w��l�!����^�58`gW��`P�#w,���n!+�}'i�i���^�Gw`��H��a�g�v���U{���g{gɼ݋Mn�N�"�NW���+O�D��*�ysMǼt[���u�q��1qwI�T^�W�&���n�舾��t�,����\u�>�A;{�n���qK8�"!�;�W������tڹM;\� uٹs:%�,����O�JS��(C���Ef��������pc���w}DVyJo���n�.�p�R6���:-���v��|�w�۶c�ґ9[��۽ق=[���"�v����{@����/������M���3ʗ��Q�B�s�9��>�y>�ϕ���Fh�^�|k�+�4�w���fc��
�*z$�����ߒjk1���N�2-~G�EG�J�T7����}Qd���xaɑP#�������\,�۞�5՜z��UA�y�n�>#Ɣ�;�u�X�%�e��1��et]
���BC��>�� ?<^��{L��7B)��eśf�`�b���sB�Q��w����@vx}���];|Ć�o�sp��a�5��G�۞�ڧ>��{�O�J�5�17��m�R2Iȋ�/g������<�t_�J2p���͹���&(7�j~je���wGW�V���m��Y�6���4�0Ѓ��b�)�I�4v���ZmXk���ڝ��1�B*���Wb
US�2��0�w�t�r�s�J9[���֦+���������d^�"��+�wt��>��Ku96$)��z-��H���Q�{W��:��wY��&�;����.|�Ȩ�ۡW����qbs�͸�{5b�����|��<��g�P�3r�qu]AO��FN�8���:Md7[�
g��4���N�]�8�v�/�W�v�N{��7��A�x:|G],���#�E�ewT�[�.�#˩�`��v}s�j�h��7o7�F�^�:��{a��8dh�F�cx��|b<� D��f����&[�Y�Ropw{q���!�vg�8{$lc��15ĸ�EZ���?��ۊθej��W�M�G]� �v~�D���h��5��&�8�ձ^�"��O�G:�Ͳ�+���W��Us�#������0��Lm+������@����UӢ^��<wpǦ����&o,����{�+��Ma^;��K�b��'Gmw`و�s\���f���{�w��L$�P�b���:~t�d�m�j�/
B��⶛�0l� ��h�8�Mek���l�D�Zi��e����a9���wv���a
0�Ee�T&]��%e��J&�к�fN���ն���mΝmn��]� ��Y)ufw6Y�����v�kC: �ђ�t�b����+g����#�=^�}�1Q�ｾ���0mm�} Z��+�_���8������hF���]�_�q�F��tTeH�dO+�ud:mR�߱I��|Ojϳ����f0��e�x�Gޕ��]`o%����ߨ���p�g��^�O����
C#�F��x*����Y�ɻ�r�ɭ�w2o��-e,UGF���+�;q��iCYQ,�/�,h��K�Q������i�P�]��̓���ԫ߰8��+
"��څ�=#�\#\Q�u���*H���{���y�l��C��'��ə����lg [ژ��՝�����=����/����� �uﭣ�Z�J�˵�,�3�:�$�FU��ɐ���DNӳP�����ڰ���^J�����j�Ny9��]����<��(�S��[��K�.dh��׋���˿�U]R�X����c�_�eX�״MkX�O�gf-_��3�#�`NZ`��ᛡ�>U3�qB��橔2v��Ҟm/��;�ʙ���.�O���(�V[�<�ӽ��Nr�B�{�i*B�W�Ջz��Q���n.�9�[|�݈K��5[��CN�7�!���"��af�'��h=�ゑ��.ò�̫���f����q�%�fu�:&]p���4ߦ���:��.���{M�{����c>�˗sz��n����΅��{Yt~8�y�S���6ָ����C���*��FN���D��l{���z#�ǳ(LVE@���R$�֦6e�{ZAwU]�����&���QB�\�����j0� �A�F��T!~ِk1{����ĒS�s�un��9���``�:���8Pt⨓�^�n��<k4K�5v�\��q�G���rEWVP�6���įV�1������yPi��{��:�z*��`>��fĴv��J�Y?��Ν��6�d�Z�/��\8�7�/���^�����g 2'�-z�~���_�>OyW��T�N�,�R���N���aĔ6t5��7^���^p앋�W�?��u�T�OB�&�Q�y�*��J�H=�b��u��;#��U��vǲ	?Y������!��� ���]�����^����?�ֆ�(N�k3��X5z�*��@a�*��e�����cdԗ%Y�sٹ4L˾[3�#ю���� :����B�g(gF M�:����[?��k�<q�z����U"�\�s��o�X�y�7o�3;���_E���;�p����=�Cv���ī=�k������qEnwi�R(�Q�&�~"����Z�:(3�n�}���7�����}\x$7LO�K2�RO<e�}����ՋLb�M�x����]ş�0������6q�.����D��Y�jjF���{W�T����2��}3����ْ?{�?�W�o{h�q�Gi�cJ�0�T�a��\vh�ˊ�&��l(w}�����N���Y�K}Y�"z���yq��,en�M'�� �gw��/~��*#w˗�2�7|��D���$�X���yQC�{&j3���*�x���¢Nq�72��>�z��b4�]��B��d1��i�z�D���߮��C�e��~2*]z�ˊS���f��w����˞���q}׾��c��B[��$����uR���4"�t��(6(FE�����ް�Mm��w���Hr��V;�AQƙҮ,�]le的�x{.�[��L�(�e�Z� jEz/"�3�Sj���%�}:��	oQ�� dI�m�J���@�����٦�Tl^�3e��ە�_^�9FD���v5�h`&*H�i��V�M^�V��m�i��E�����}p�Pu\�`�U/h5��o-򂋘�ݶ���e�Ϸ�CU���t���T��\���ߢ߶���4��������R�;������?z�(h��i��a��c,�ݪ0���[�__��.�U�3������<6W���3X2"�e(�ʵ塒ѧ�9�Ǒ�-�u��_�]MU��5ض���M��`�#�.U�fE���Mk����jǩ�����a����N�j��{3�SL.��{�o=���m���7��Y6�w7�䈽�T4���#A϶� p�]�5~��.�������~�M���2��Fȣ��4�#���1�!ہ9�!Vl�]s��Tۅ�1���}t��P�zx�~/L=�پFL�r���%	Mc�{dd,���oS�<[����;�V屩|��t���+Ѯ�WJ.�-��:I�e^�uQ��_U�m�EϮ�v�ÿtq/R���޿o��lm�f��V�NLJ����ҥf��,��]{���]g�n�J�<�c��WW:��vk�D�f،m��v���6t�׽.�{����I�؆�4�Ro��h1 �Z�&�7�w-`w�89��v��]:�)ū��t{���שugb�&9U�՚�<��nu.�;���B�(��x3'T���NY]Ĕ+�S 4�f�n�4x���t�Ӗ��C�Y*d6+��+����,�L��q<�εX� ����V��v��8Q�^H�͹�Xjُ��J��������*l�of������W�c��0��r�7��{�;�U�����'���(�(��.R ����`v�!4b^��$���bf�=�;P�7`�o���.��{���T8�hq���@��!���!8���k�	�ԒE�J����8ש����ԇ�7��f����x�I�Y��B@�^�f����!��y�L~���w\�K���]m�BN��H}��}S�M��f-5�ͪ�F�Tnm[l�W ���@�2�h�+��a���j?(	p��+ gp�s���|���/~�N��y����s~v�SfP���@Si�^l��-/A#(wgn!F����}[��$4>�v7������k>ѶH�kD��q�v���9��끴�IYr铬�~���N���湞jb/��BI$<�1�r�����Ϛ"�����	yt�c8�]?']�����;{�վWhm:�^�?r�,:'����a�IY�n�����m����Տ�i���ڭg'[�*��H�{C����B��۩��0���ԕz�R�s6M\/��s�I�L��ޯ��O�u��Iu��Y	'� q�<��}a$P�$<�0�ۤLg�2�n��8��}��@4А߸g�d1&9���O��mx��������.�\ֶ��nئn���C��HO�M�y�j@�d>d��5��8�f$�]�{3+D�IԄRI�6��I�X�c���yC���Āsw�=sY��'����܂��=�`u i��q1�~���^����uj��<���\z�5���P�W j�"�_�E�a���dPŔG�U�3�}��ó�\�t�_:��3�w@�l�6�q��`�:�����.�>�I��Y���i&�+��|�u i�� I8�H|�1�	$���da$�<�� 
 ��av�����/C��eC��.��MKR�WJ.e�YΖB��A�C�+���N��empbb�HtE��&���w�f��</�1�ywX�6�Q� *����L;��x�pGOr��I���^����[0nÔ�T��+��CsM��g브_.ηo��Գ+���=E
�b�{}v^�����Y�����d�Yx���|�K�+�4N�gxw3{�}:7z^� �YC�=��>B^�y��X������j�a���7;�U�is�uE�!����v�tq��M{GORk�軋�/�)��x)��7�1��M�s�\o\�k�Μ�f�6f-2��r_e.��u1�X�8�t����{�]+8�W���i�̼�@�.�F��
u0nhS����#�g1!~\XlLw[�yx�g�ko��-XX�ܚT�	�6�R�k���7��ONY�ո)ʔ�U�Nu$�<�wϗ8p}�����w������)+M�6@7s�I����v�T�]���OK��d(:穣z�k�t���kn���̮���8P�*�p[�]P����{��Yq��l���;�s0
0�Ig5W��"�t�N+�c�3����u����7x�e��n���fI����vk��p�n������\ݾ[��|�x>�]N���Il��\޶^o���W�T�Pλ���-_�h7>����Vkw��T��������ai�TL�����˷9�8ɨ��<[��i�)OT�>��-��U/�V{?����I����S�L���-�ə��ख़��ͩ��e�|���$�]=�u��|}���Y���_܄�#�_^�&^���z(�r����{��ȯΔ+�`��,����`2�md�c��G�T������V�u$��<�c�w��Ay�!v��;ј��G�8��Y����Է;j�3��h�{��<+O��9���<��s���\g&\]\�>�����7�������*�������z*�K�u'�s��:`����Ճ#Hn�"�MS��re1�Xι��V��W>X7W����<B��X=��7���c�J:g�-�$�o�|/y�ua��[�ؽ�����UjҥǨ��{��A�/���ׯ������g��m����Ci�����j��U����_��בI:m͜|��k�1�K9;a!Zgѧ�?x=!�9*���֟R�g�Ϻ)_~�}D������kY�Ĳ"�2��}�vm���5���Y��R^]#��Wm>F�:�%�5ں�-k[j�b������^4�B�\;0w$$�����5���H�zĶ{��U�\ӫ�qe�C(���u���K��"���=Zy�Gh�!������q6d]ա0m�S]��ՠ��x:<�湋���F�X=����z�k�%���L�ink��;b�v1���=��ƈR��J�3�{C�¥Ӌ����������;Wd	��S�uV��nէ�O���3�ӻB��?��eb�σ���������9�<)'Q�\�y�z��>�����W�?,fK^7^~�1��T����*�#��+U	��`�^�̙pF�}�z��-?.{�z����BgB8%u����\���~
5��(��p]���9+�1�=(�f]��1y��ɳ��gU��7�#˗�������煉��S.q��0��5z7C.�#��έ�'�Q��9�WN�uк��1�*�z�"���*��X1�#�]�^�:��=��N�>�Y.�h��$``ӯ��Nc��.��`��_�fjaìWW�]{js����[P�i%s~w��tU�:�ǆ��J[<ꦭ�t.��ë�r���ɽ�|cm�'0u����b-孫|W.N����uIձ�mr��㯵j���BIN�鵀�M�aK�z&2a����nwZ���*�<wF�k��auЇ��<�
f���(O`���|3��-�_r����,�]`AƵޞ���E�>�ow6V�i[��7Y���ۮy����D�Z�O:�6x^i�3���egj����k)��A�(��VV�{��Eԭ���q���a��z�S��]bm$"�8QF�E��-�{!�O�e���w�N�]еozEf�Z:2;r�d�غS��n��s:乣��פ�5�6/���ڎ�˦:�<��^���3�#�<&/7�Y^]�_j�IX����/Յ^�'w�⤒�`�w�NR��*$�zţ�����o%�}kٰ#Ҍ���%ֽ���uq�b;d��4�O����?z!ݐ.��;�i-m��
�r?��-M��(�s��~�� G�s��OS������t��'r�z�7�rͧd;5���m�$j���m� �z�V�]V) �f�����J��]֜��f�P>�j��ɒ��ޔ�$U� ��vz��I�p��,��QwR�����&��o>Zc0oF���I;ǹ�#<o�]`����Fҥy���bmu��Wn�oAͶ�#;�FD�b臅�u�#˽h�\�" ÉF,�%{n���c�O�����0J�����(�q�V��1\�F'��x������{4�p	�YbL��H�L֨���GI����B>�'|�z�P�����Y�rN��k�J;���#��}g����"�c���Ͻ�����k��~]�{f��������ڞM�-sW����]�R�F�تt���mvz��z�����k�ְ��&�Uذ3k�ձ�n���0��݈Fː�73rj��WٝO�wn��D>\���WS��hH�P6��_�K��wgm�ɸ��t�ml�[_�4щs#ʫ<e�OJ[���&�Y�I�t��N���_"�_�������Ja���(��+�ɶ��I׌���55���T�o���lݖ�]�{�t�]̫7�gD������c�����3�d+k��R�ӧm<��ݶw�J�)��)���F���v�m\B����Yz�UR:yK ^skc�z������w�V\�pg҂c�㽽P �9��$�1v :
�Yx�μ�����M�V���-ì�/h˂9op�c��*t�}׶1���1����J��{�^+Ϡ��(�t���i�}1ٖtt>>i?u8�U~��ck.�ʖ땷f�xB�qwl>��h�=*��h�������LǞڏ������vo�"�ճmt5�s�����5"7��#S��CN\�)���7��S+g�6"F^l�Y�:�?��\�H���H�1�f#sU��b8+���s�+V�&�Z�)�Qޭ/�ʪ��w[X_�ǲГn��{3&tt-��gb�vU�/n�΢�����%k�䭒h<*�|�Rs{U�_p2.�¦�B��U��0S�d�q�][\0l���d���,�ʔ*�{����TN�Z^$�����x�t^(���E�z�hO�L�w=d�Q�f���"��Q��r��㣙���љn�J�2��2�1B�ٮA�or�Z.v��f���CM�����{w��PT�U��l��T�����z6A�uK�y���k�k�����ۺ/�V�l�F
cxm�v�Aj�5�r.�e�$�'��բV�뜑�K�������@���]5v����P��EG;�n�d��^���%p��)t[	6�}@)��]�iU�>)���'�l]++�oN��X+nQNJk����f�|%����9$؈̟sQ-����'�ڼM��șٳ�5���>�Q�Fu�J����8lJ{���I����,�?�O�����M�N9J���uȸ�]C�C"h襬`~���єO��k��^g�p�5ש7��R��./�����p�x^NߟI�E������`�[Yz�K�6/}9�z/t0lW<��b�^�n��b:�G��?_L�r�y����1e�{��wsB%��v�J�����5^�Y�,�s,�ޱU�na�O��DXr^�fG�Մ������h�n����py`����r���4ǰO�~�B�g��ݿ�e���,V%,]��+Z<�v�̓U�����=L��]�S#�}:�<.��}���u�hB������snd�9�f����	����ob1�>��d؊\GK�����F�4���[b�5��k�j��S�j����7=����s~-�+���f_;�'Lm��&[W�RλÍ�AKLe��.��l�؄�U2�zv�`��#�-bU�{���"߷h:����-keu�[·c�;GG����t���	[�8�[R�o�/��/��=�{4���
wu��1L���Q�A�ْ�%���i�j���}�aT��OUh��y��\WA����N_[<|Y=ׂ�tޓ�?Z�����W�>{�kX����D�D'�F���bu��Y�����Z��3:G�|�����$A�P=]�p��C��f/������Z�z_������9&�k<y�u9`QG����T7Fda�Jr�^@�׏K��ck$X��f#�r_7�s�#ڛ�y�$��|��A�oO��/�_/8Ξܺ{0kO�x^���to^��wu�p	�'������p݅'xzt]��r�Έ픳w8'�{�|��E�{v��]}+�q˄dT����¸ú�1� �lB��GWr�1�̂d{������,�nv	�uܶSuo��W�$۔��)��]Dt_���`��U}Z����vS6��Y[kc���G���Wd��0[��JD�����S�]N����ۉ��^қN9�]}�粃��DҎ57T1P�ZN�/��-{D#�B��\F�}v<"��F�*�J�������Q�[��\��A��Z���#~��������Y���\����C���C��s�5����1<�pTv��Z�-ڧy���vD8r�Ykf���=��8��q�&rӽ|0v�oqT$�r����ҏ��;���7�1��IQ[�wr�Y��Nm��{+'T��W\��Z���M��W��b��7�/ʿ.�ߎ��>X���6�pk����g��w.m�Τ�C�׼�J�r%۫��B>��~z�Fx{k��wE�fzow�X�h���{�����HT�d�5�Çz�5���MD"w\}[6&�|w��$+!s��t��rN(g[����.2��1�o���&f�l�νt�P�f�&��D�4^#��]�A__w��=�;�֒�J+�}��mӃ�U���|���������g~,��O�$q����r}�B����qK�:��&	Z�x\�h��0=�ޑ�o{�Y�F���<zNwIj��s����%L�z�s;5�8r`Fʹf v�Y�]M�M�?y7�|F�_��ĳ`�8B��`�ҽ��O�����)~�U1A�ʂQ�gWc�����O�����.�o��s�mzh�d����ظ�6���.&"9�dl��*-���i�� ����iw�:V��2���Fde���Fw��D"�T��0«���Ey�ά4Y�B72~fJ�j��U�q�����]u�.�p�Ҡ�aeʕ�f,��ٻX;c̜�䢶K5Sd0���|/��K8�>�a㳲�(��Z�˂�� �u�pҥf��JLJ����m힛]Y��U�eKH�o���m*���o��oN�a�5e=��ol�v0uu�3�$Ϣ�M�ř�V��N�>���7�>�u�2ޝavɨ3�4�0�����E���6hm��Nq��k�}�p��Fx�]g�ʢ��5/��fm�x���t/g�BW1[5�/t���˩6�7p⧲��ƴ@he�B���em/O���ˀ\��g=�����t�t�ow�9!Ǒ��]a�]��r�Q�P*��M�*"���*}��,-\��6�{:����u&<�u^_ZQ5�j:�3R����"zq]0:���n�޴���:\UqNftWPZk�w~�t��'&_0�rU��g�QL�n�W�t~�Ź>�~�`��v9w�
E%�]��s�It������X}o�������j����;+�~�b\M�pb��9��6	�+b��5������ͣĴ�b'�"|�u���[�n7�Ok��;.bt�6��@��IÏՕ��mP�[�\`[��Sj�tC��qnn�SU[��E�s	z)ߜ_|��=Є��E����-f������6����z-��Q,���u>��멬S�{c��f�Q�A�>9ؘ��C=��k�
+�$uw�c}"��yM&J;=��^~ZQ�����n7_���VJ��ևi��E�r��K���,��Gv�+�r�g4Fg� 6�R�:,<Jv�<,9�u��㲔u���}h���=�udvՌ}e�ǥ��+�i�t}��n�6'�u-�=:KE۽��:dk_T�����{
��ÏX%xS�W����V�D���%}�ʵ��u7=�3Z~�?q�T�>աbc��9r����:��X���H�/��N���f	�^�#TU<e���y����~VawV�����2u�,u���}����v}w��X̡�>�R
�m�_�?8��y�����$�8�l�ܦrAh=ۅ���ӌO�abS�&��~�4κ�H����0V{��=2���>�sW��F��&i{J���Z(�0�A�຾��3Y�;��>Wv'��g���m."t��G����q+��Ӆ_z��?jO�`��{�!�Ƥ��J�iܡw��5��(�����X���\��v|�M�
�ɐw�b�|��#�<11�P�&Y�Q`����{��=Y�L������d�S�ɘFףd^�_�T�_[݊��C��CN��xF.cfO��S��ԕ���P�9��56��vk�2�M��'�dh�]S����7���N���]P��/��0����(�Sr�/y��y�V�*Ƣ��ycWAu2FEE\���G�<�{h�֬��M2��5�]Ԥ��\�ť^
�w:��#%�.�P�lS˺
�2RN����)��6���oW�"�蘯	<{�4zXL�Z���w����V��4�Wt�uo��C��f1Y���y��ں��m��
�+��:�g@l��q�Yc <+uV�x�.\���r��hk�c4�<yd	���*&؜��,��:�Nִ��)��+k�[�������ͩ"��#_V�֛{�� ìo����H��10U����W}�ZwS
�31K7ӝ邲xՒF�XR�,��Х�3�,S���5W5J����}_�����_R�M�%ڹ(X��wH�m![���ȩ����̝]��G2Ի}�f���m���ۭ�6�CO���	�ok�ʪ����G�z��cs�]KA��DCk�/�+ꧬ�1|�x�
�A��7�oZ���a�Bi m }�n����p�3&s7�nkYIIBjF鐶�樬X(%tn�j�W��ր�T���W� �H���Ӕe�B�����6+-���SLz_b�I�T�?M��Y}�B��W�j���-G��\77GmTT��4[���qp]we���b���"�^4% ]��U{���Aig}���p��8I��
����
���WVa5��ï)����r�hKT�w`��UEK62�|q��页�.��K���Afe���p1V��+���N�=�-��� #�x�N�*���b�WD��>�k���X�>=eJX����
��+0�]�	�2w[�_X$)�d71��B�_=�5*e��0�=����'&KGQ��e֝�L�棠�H��l�b��GO�G�6�n��k�7�M��^Ks���:��)�}����HN$�d	��O3�!��l�� �8�P�'�*�.W�v1xS��J��R��*����#]�*̣#�	}#�R���.��Ȫ]�cw]].�Li���R[�B��q���6����^2M� �ƞ��d��T�Ip`�F��QأY&s���EZ�	�|�w)N�r�ͼ��ca���o*	j^��	].n��9�q%Cf(̓���ma�t��q���]H�,p+*�
9[�Ӥ9����&��en�%�e�M�JR�F_{f-:E�I�X]��MQ����7�P2�mv�Tyt����=���9]z���Bj,�i"�\�B�N���]*������DEV���-� 0Nr���X��>�k�upԷ;5������y?C�~��� ��k%x��ʧe��p��1���0:[[s{uQ]�iQ��<R��mj+U>������T�f�\�d��L��S��o��M��r�GcFX=��D�9��!��O�qP�e:�Hv�Jmjƫ��5²(�6VU�x�^@�<������\z������ʝ,�wP�U����%�J������[ݱ"h���e�z�;`Ӷi���m��v=+U.Kb�t���"7rv��e���Bf���?b�u�Hs[��u�{�u��T�B��W�a�;���2�Н`�����
KO{�Fuf�-�o_�D�p�K�]E��+���3�Z]xp�*��rr���m����!F0�~�,V }���^����~f�A&��<�]����y��:�x��d>i]D��+-j{��2'�_u�m<|w��^����wm�E�Xט����]o�c]M�'F���2˽�[$K�RN����#�z��x���qI���+Ϊh:	i�n�$�1�׆-�OG�FQ8�{A�f͝��gw/M��]s��Pw!�&8"�����6�v)A��;d`�\酫�w��^p�1��ޮ�9я�gOWI��*�����Y��x�T1�E��R��N-���qܽ���]4��Gծ�K�stq�n�Y箠!>��?(ӯxH�����:z7g|Җ=��2*|�&F!C��"���1��sp�>ϙo�wΌ���y��U�$�4�*+Z�4%C�����{�ae�u�`�Xs�b�!˶��..+Я=#�r�Ж�6;GU��HТ@�]������M��Ap�s�NF�mIB�����(�BG��*�/c7r��~�˷CLʃ�X/n�7y��foy��v2�*����3��ǘc!�-��4���~�Ӻ��3Մu{�s��=#T�8_�<��D�e��)dۻW�nl�7hB�;�̩Ԍ��op�B��{����l=} ��;��G��c�Ѥ�܆����k⬬ t����:�Z{=�V�}D�]�[	>�2U���T�di�X�Y�j�7Zm.7 @<W�l�����+���[ۋ6o���E��40��k��y�MQ�t��~�#ޱ�/D1*�&�,�[�a�jG;�s}�lb�@�t�e�����J'6��ں�g�yo��������e�<e���b�@�y����1���Gץ��*mC�C7"�N+�tpq�jw�X������{6}*������蹋���E[��a�֯�*��@*Q�ؽ��ڃW<*#U>��x<u*m��,����s��廴<Gc�R v�ͬ��`{<��#닕�T/4U���u���y"��@��+�U����*o�;��E�küa[�M�E^��0��:��{Y���kd��+}�U�;֧A�T�fwn��[������}nqvP�W�F�ڦFeO�������ީ�C����ئsn�R3��'n�::�߾y��is|�⧤����6�1F��O�=�cR��$[����Dߤ߈���{���}[d����9�V�����l���G	��Ы벮$s�{�xp�wx9>�ڼc����l6�E����_����b��]��s��m�9���w�:�h���9r������>����a��][z��)���!�v�h���B��q1c-��TV�><�lVLh��§
ԯ�����P��r���F�)VD�D.A聶�iF���t3w7�����\qI��V����F��+&wq#�q5�M������e����zcfG�̹�������]3z�;;���ͱ0�]c�
��Ri['#S�G�a2=�Mw��EI�:���Q�ۗ؜Wl8Ǭ�5�]��Z��s����-����)���)�B��T,<��q�������5�>�?!�Vpnj+K�����>[9'��KU�4���5ջ3g�괿&�����JC�9lF���0&te
3ݰ��Y��ۏZ������T��(��k���c�V��]8n�j� ������B�3�	k_�qp���V�k�bU�ﾉr:��/�T�ͨ��ٝ���(����Ȱ�$p���e����V&�*���[�3H�Fd�xƛO<�dY?.��z�]�{���y�5B 0b	bB�j/��1���]ʻfKjF�a�������oچV�
����q=�B�Ɍ�s+K�Sj�<����ѳ��u�X/e�7Ȥ}���֓y[v��v �{;6�T�-�Yv��/�s�)9ꪝ�7{y�:�<L��S��K�<�O��������fPgg�X��2�e��t��~���B�qV��N���3�ܦc�(��ۍ��D�	��P"�b3�+s�I& d��ۻ5֩�֚�l*-9j���"���8L���njA�Q�s�KҲ;���d�|��rw>�ěu��x���c��k�b+��oP�tM`�����V�I6z��)pŇ�Y��������B��F�K逺򔅡r�ɿ}���zi\�� To�7����5TM��fO���+A0P�� ��q��T.7��T)ۻ�ˍ]|���~�op^�����S�Rz����0��\��#X��,Y�Ϥu�ڭ��0{?�1�Gq�V"�OTw�xษ��\�X�������D��d����9�(j3�:l�=�����˓�Y����7�hLn���e<SAU�آ��֨�}ҏ`��M0�ϬO�_ҳ��IT�G��s'�9ͅ��A�����;�_wGL{d$����Vz�o�h�3����e�xz���xs���,�ضrg���ܑ���681�9��lh��Ŧr�o�-4Q���}����up������+�*��]T�ѷ�'�v�����{�[�����W���b�#�n�;�9�.�'��9��z���AY��Q^�@K������
��p9�J�^�=���ܘg��ݬ���"��zXZ�z�U&WkS�ۭל�"�	9��dߓ�� :���J�T�N!4/Pu4Z�Nō��ĥňF�%��X�����f�6�q���=��3\V.*��&��.<��]��v��To�:��+$
�hX�yPfä�������#=D���W>ͬT������{"n���z�F��T^�D�[�Q��yOk��7�������f�,=,��Zlm2/����qW��sl]���g,"�<h9����'W����9��aW<�81��7�a�4��b;0L�N��F�r\�}z2�����2������4_d�Z/�m�^`q�n�����#Ux�C�7-�<���f��}Y]��	�/.�o�1;��y�ǉ�[�7��;��{�(o�j���wT��}bNBUN��=)U�����������r��R��>�s2k�+�=N��Ӗc��B˽�|�o����";-�Y��D{sv�<1��p���X�}N�=�iug�J�pv���V8�M�&}!]�ʮ��C��'��s|,�f:@��8���=t8�c;�o_��c�Ϫ&\�s1�`\p"$OT���ay�6k���uFZ���0�^�qOT���� �Y���tc\���B[T��튁��x!`�w����U�=`�k�~ˇ�k6������r��}�l�ď�Mv��g}�a3|�z,=��w~Y��[�~�QQ�STd�z�ûtF���D��M�ً�
+�b��p嬬���K��\s^Y�"|ۣ��0'٤��:p��r���˗p� �g�U\��]��=��!�l5pn��C4�W|�w���w�V5;���J(=72�q�M��������9:�L���Ü����w��]��\?{f�{�h?l�Lv��!VuE�ӥ�؇:_��V���7�˧��Q'k}r�v����1\bNנ������U=�e�T�ɩ��
�����GjLF)v}�)�������:�w��1�y�E��S�"���~��8A�u�ڑ�?w��7��o�T�'�nk�F�͙�
���;4�����d�ITԷ��ff�t�o: 湺#�5�y�cܼ�z�{�Im�)�SU~�����;1Q��g�uE��+�?n	]ص���ouC1Я#.nP=�r�~��Ziqk��%O����y���Q^�0�?Wvfg�w!>�6�ɛ��� Q�j�]ן]k����M�"�p졫�U�Z�*$�c!�"���㠳Q�jJCطѽ��,�n����:LE�Ux��L�󉾔�>��	���ʀ����oV�k��tOX�� �7V~��W(�c?Y>x��K]�%����9�2�xS]bb6��K�[=�<nGX��+�:k%�h��վg�~:�ߍ���@� �>X~��Aw�EÃ!]J{�P�ʞ|+f�����l�+ �ަ�]���:g"��Mf�ӛB�G��vKB���U�U�m�9y��� C���Ysʗy4�[�����BU=R\t`��L{��άZ���_-��of���ø�y�Lj�������n�s��gyߍ�׷����l�ݎ�.e<<�1�t�@�p*k�~F���M�bn��W����5^��<'��c�^V�#��ЯڞZ۵Y�+K��!���[��>�zc�B�T�SF/�����ͿG�R��p��m}�4��#_	]w*#@���to����0�C�s>��Շn`0��ӭ@�C�F���I�R�k��w�O��].�D�J,�"<�Om�0EC��G)��{՛�&��s;�o�P�3Pp'ъ�-b9��
Wh�w�Z��&/a/�������.�4���?|3�mʭT���d6�q�s�ܨ�����k�\!�n�m@6�ߵ��7�LO��ORn�Zi]��l,ꇡv�
�{˂�;:	��{��}r��1Fs�ն+t�����r�gP�>3�]�\����߼�	˙���긗OMOZў�T:�a��uh��隽�$4wΖYw�Vgk�[n4������4@��/-�s5҄���WW�ߴEc{>ܑ&�_��O=�6���>��1�yMù��v�R��I都޷9;����7Z�x'��ю���g��#0c¤�t�3��VR+��;l��.��9+�Zؘ*4�#4�/w�}Zu�o�<H+jݎ���ٲ��,�Vj��D@�G`��v�K�z_V��:>�$�X���U��{�#P9v����oҜ4<�a��}��0T�W����3g+��Z.S�j#�����b��G�x��իq�f^�n�����h޸��܏2C�Hׯk����.tS��ء[2W}�9��Z�9�rM��z����kr����yV��y&GuTE�ԍ���	�:�%è�5O�S��3�)+���-�Z"�����>�q��<�%���ތ�c�ɕ({������w�.�Êg2GB(W	Ί�7�ٓ(��BW��v{��.c�-�����\�R��\GM9�M��:��c��|������d]��m����Q�!���I�)v�{7���m\6����l{�����X�j�8���*��`���ޔb������v����y����x�i���WF�����ټ	CwM�2��`bc���iǁ��]���\�n�,�Y�u�%^�Y<-3���7Y�^W�׶'؎��}��j}Bꐛ����g��I�
�J�Ln���^�N>
���x{A��Z�v��>X����6�H��1e�r���L�=B��C�f��:5}s��j�D� �L�NȬq����Z*lys�el��;;���cC�H��{}L��a�����S����pR'/�f|��< tOn�z�T�s��ye�N��-ff���������	}�ƹ����h����`C#��>���u�wŢY���;�n5н��Ol��Me����Cz� ��ܚ���:�ydV�>l�ץ\�Gn�{v:�i�;�V�т�'���Tb�Yk6La��b+���t���;U7�#���]�����-z��!�O��U�e����b��1�8;9�^��qV�E����	x_�s{聽R`sOOz�ӏGؙ�bTq�gM;��q�^L��#�}u�� �I
�{�g=.C�
c����l_���q�bdOF|=5/e�����'�H��P���C�ew�b�Fj)L͈F=��W�KG��]h|m[��B��i�r\'�ŋ�s����C�z��u��a\=�H��wG5�b�9��a�&'.	�]?e;wjD��<��<����1��p4�r��6��c���We�&$�u)���1�������g���eK��gWx�p+Cg^!u캅e\��{\��qa��q�	�ށR�"dd�O��>��v�6uo��.PFr[���j'�c�L\��n�U�c��7�,yQZ���>u�~>;1I�&h)��h�X���k����y��\�Y�/��­WY���[.�EY���?�J�r�Ŗ�ҝ�G��m�z+�d���)��٘(�ε��ge�]���sk$/]���o*�� m�5�umC��m,▷��+Z��=~�JW����=�&�vc:a�;ԫ*:o!A3�d���=B�jѻA�%��fS�bt\{ul}��7�<f��n����^��\VΝ��W��%��b~�:�g�1^ñ���)����l�x'S��r����l��|�D���q�6�#JLi�D7�Srr�s{Hj�\I3%�%���z�dh�}J��>�i*���Ⱦ��B���(�-��۸�c/�Ub�ϖ�է�lP�ԍ���:�}����{��;f|�6�q��R�}�3G#n�G�5:��C��ڪ'��V��9@�����
fA�	����B��ؾ���i9_r�7���<)𤤜�w�^o�(P�91��co<����D��W�#}=5QP��d8�ݗRgc��WV��i��L��"�;���|V٘�r�ɪg��i[��&#�.��X�VP��G\���m����r'`+�Ǫ�;�8G	ڐ��G�^�A�|8�pL�"��ddˢ��/߽�9`�S�hܭPaf;����-��4�6n���ڭ�
]dw�E<��L�TEzo֔�yc��EH����j�7��;Uݻ��dz-Ԭ���h�3M�2�V�ޣ�-�k�|�rޗ7lݫC��E0�Q�c2 ^���fJ�b�I�F�B�	�E���)e���6��(�'hA����y����7lrЍ������nQ�rbcԫ��X3�ogN)���Y� �H�Z2�i��G+��o���Dv6.}��۫� ���,����й��Ch_%������ω�5i�z�:&��j�ska»3-�P��%ث��p̈f�]�]�xu��&E5G1���=է$��:�33g�lgm�Uںr����M���o�vKԅX�qq�osǝ�bJow%�v��=Ñ��λ�}B4Ks��BG���/���}����r�h�u�xU7C=8̨M^b&�@�c
,��e�x���Wu~��c�����5j�z�@�1]�.�Ǒ�/M��2-�����Eb�f���yK��fu��7��W����fD�bl3V���U�
�@X�����׼8m�[���]�ҽS�H;<+�M����T1�(-�f9J<��2�� �Vay��kכ��9��u�}�+%᥹|Ƥ�Z��:����#Ok�yu�%�)wa���wl=4�X움wm�þy���.;��ن.����s9�+�]`��3]�1.�1\��.��h�L	��Nׅ��L��lj�c����+oPٛwp���K����:�aا"jr���D����#�{��
tn��y(!��Z���J�.opޔ�[h�u*�M$��t=��O��X:�5y��������)"�������9^��������Y�2%b3�t�εJ������)7�c��v��6�݆�;�}�F���!-F��T��t���;Y����⦩���E�fm�7�E�]����շ��w#���W|i�B�>��</%M�(��a�vz��3s�ʨ����G�ċ¦��t��c�W��+zn�&�l�HV����	B-u��s�Uk�� !�t��$�A�3n�ކ����d������4��*���`��s
�G)����ӳʈ�ծ�*�Qɗd�Eh��;Lī��ӹ�m�bZ�.���{]6���-./����Z�N�^Đ�Ꚛk��kݩ�VbU���1^Aq �X�._m��}v���@�H�N³�;��<�*��=�*���8�~X��V�I����I5�i��I����=콺�KECťu�
K2��̀�K{�̡U�"��O9�V�ef�ucT�V���KϺ}�>�f��Q�)��	�]O��&�v�o�7Z��1�37JR���;k�b
����{l����}�u|"4,��C
ɘ%>k�D}e�nA�L�e�U�&��t��P��/p�}��)t۝��TZ������Yy��a-���G���`q�o���DW��4���B���ʏyǨrӮ������I�n�.���Z�Gt]��ggr�vpз���NSm����c��V�f��{4!�O,�6%k�����t�����e�8��T���+�N�1�]D
��=��Os5�˟^T�ą���E ǫ(_�����ɂ����ae}�\YYN���)T���jngh�CQ���=jܙS�D���ݗ��ꍋ�Q�㘛.��
tx��ݐs��s�ȳ+�K��|��w���=����9S.pd����<6\yUgJ�c��w�}�F��Cef@س�&]N��>�E������d���%E3�;�"��:�[P8Nt{}B0�:k����F�/��	Nz�<��u�bw�2��v;wI��Pb��HPkA��X�YF]F���gȈ���s�y\_G ���3�p�m����'`H���/�j��,nH�	�#�0�u)VӾ�;�[��{.wEY�׺
�4������+M��i�����|21B7J�h�E���p�^�U^�;�=�`��_m�DyA�ߙw����Qk�s�S����<���գ�="2�b`�釙�3}���޸�\��¦b�s�=��c���7��2Q[{�#����R�ԴWE1ߞ1s6���:� B�&��d�3�k��]�V[u�Z�O���7��h���2,ht���ttG15�4���	��,�{e��r�3��R�w0Q=Yg�����orwS��9\�,�p��
S���v�����;˰�;��쓐�>��3�s>��;�z��ɼ�t؋��$��d.�^�qû"�tq�qw]P��򟤷xd;]2�"�mlL܏t�S7r�=�.���AtG��t�bo�'�GO����_$ lD�6Xf���ۋə��}���ܕȇXy7ܩ��@w��+����^��ѫեP�WZ�*k^�������zk�/��V<y��/
}⛫>� �q-�����ݝ�9��4^t�C�2/Wl�f��d���E��muUڥwF���L�F�{f�E {��Q��Ļw>>����MW���\M]m��[*,.IaSq~�Ɨ�sl�O(��u�� ��Κs{ʭ. ��#�^9�x��Y�ި}���m����v]��f���*A>anK��������m	V��ܺ�OVS�_�-�aۡ���|��sFey�,��&B�,�y���=���qb��P����T��Y'rl�}W���Q���~ɝ�n�bKn��������x��'s:U��Q0��Ԉ��j|�ڣ�j��TO(�k$���l�a�c̗��\�ҹ�w7A�:s�v�ټ�k�C`�z	�E2�}5��%ػ�\̔kvwokۮ`���۫u���,��ޭb*�,N�t �T��9�q4it��v�V=ެ���nѧ��G;��cn�tr�:��p.�J\�WT�k7Am��b���Q�.�k<L���x�S�X�g�]��9��r#Wbv�T*�pM䎃�0IڥQ�l?㔼���{E�Ŧ����l�̠�)���W#���R���Iۆ���@��ϫ�ǽ��/ֽ1�^�=Y�\�Q����'Bߝ�pa��ޡ:�?LL��s��f���r9����O�0*;ƹ��N�dI��Q<��,��M�������F�SN��ޛ��R�F�����BQO��*�9�ꟹ��p�[�Z�ǻ�����-�0A�פ.��5[8�+'����q;T}�;�r	��׾(\ns��a^�ƶw}��p�q�Û<H^&9��f�ݘ����g�'�+N��x"�:�;ݜ&��+y�/{i��8�#�u�zC�yQ��]����;�YKƮ�ў.�ʟ+�����
{a�ؒ�����α��*n��U׽+���,!�VyumƝ�Rj�p76~Mi�~��V̗-�^�t�d���H�c��wͬp�۹���1g��麤o�����q��l�nZ��Sr�^�O��w?NQ3?][}�Xs
jվ�f��t]LUaqc��ٻ:���c�v�.�Ǖauή"����N�(���J���I�B�Ս��	qغ��"�&�*�݁%=w%�4� ^�0�)���{&�[��G2^�ofn$O[�oe��w��s�~(�䌋WR�$�I��g�8#ݳ<��+�B�$s�=�j�͙]Tڻ����r5����e��n�����(�Qn:}�E�׻WSA���=Ī�|K�C�����o�+�IB�o�(�o`U�OL���3�ֆHo��lȎ|Pb�d�CImEfdY\�ub��Q�KI���ȿ}I6��jJk��S5oHp��HǦH��λ�qٵ/ ��K#"l��y��e�W�Y��|�X#��?g�P�n�	�6ddl�r���O|�c'��.�u�tn��H�u隼=�_���%'��_��:���"�a�����Q�N�b��=)���H3&z�f�y$���>>ٕ�����s�Y��r��n�g���聽B;���7&	>�Ά.%w��FZ����7���y�i�ZTo���.����&�%��
Q���،6)ϧ�ہVExc�r��Y!��<Q�c���Nr�ވK�X�y��Ǌ/�}'ޡ�Wl0�dO��Z-L+�S͒�6�Px8�R�����K�9/;�P�Dy���x�VN��Nۙ�{Ք��mz��W���^��:䗚>��kK!,��}G	��l��lWS�yN���.����[
\*�57� ����Oo�P�G����I��.,mZ�
�ݔ��{�EQ�� 5K�$��K^[},);&as�w"�J҄˱��^�p>b�+ԲK��]������)G�@�[:Q��o�KY\���2�I���r��xz����&N7<�SDv������؁Y���X�}�]�Pg�W��?E��O ��OWq5<�Ϧv���q=�ݟ�wB�.C���2{K�.�_L�h���Y�]�E��.���ط�N'��X��J�uz��w6�@峓nGg4`J�V�4j0�
��i��f̅�V�s<	M��	̉7]�3�o�qF��<�"b4z�-c܁�}c6$��ɗq1W��
z? ���Q���ܾ�S�-ޱ�Bd�}׳����!�Fs,S>zM	Gc���`��=����-��CC�NW��h�ِVx�v�S��}r[��VT�\19uv�-l�it�1u���-<��?x�C�b֠����K������AsgX����݋𸡛�_=�wf�=�J��*2zn6�Nr��M{v�mJ�㽇
�QSsS@�l�y���{r�>a����6�s��dT+~���	��U�s!6�y��^P+n5��i���!ف��̏_��c��Af>1�$x�L��-�;S�-�m.���u�r4�Z�ciCS�m�N���뛠�{�ue"�jеV�;�F%�Ӂ5I=�3�,���2�G���֎��_L�VtҚ��'cU(��ɵ�Gr�L�W�)�k�]��Ul�J��L�0�.�}r�-�ƶ2�nIZَ���Y���y훈ʭ�oIB5�Bk��>�ƾ�]a�.#g��=��]ssU���q8�2�*�ER�>g]57�ö���c�rN�]�.�J����g�rʂ��n��^a+�laG�@s7F�{h�>Ch�k���u]�o�h��H$�ðS����������̾~���W���OE.��ޅµ��{Ւh���B�[B��!�k���4��e��;����m��gOEO�=O��#�c&\7v�^��tO�����a�7�b).
uM��A��J�ޖ���cQ)�芸u
XG�Ȑl��.'��͜�:�1���s���:2#]+y����؜�X%�;�oNԺ=��!��ct2�e�WX�.���g"O�R�ށFd�9^?\Έi��Y��Gu��al��g���E�>R��s#�Os�<�l{/���b�xt�Te]�s�z����b���1� �,��=>��B5��9{w[޲|�)=6_s(�W���Fl����xzN=�A��zv�`BgJ�c�����ߒB�)��{�c	��'.WWLc	�܏����W�H�N=��-��Yy`X�mR�|/w��D��i��*A��E
��yVq����k�UX��=ZJs\��3�������O���(����h;pAT���X������l�;��ܶk|N]���c�Ş��"��Y��-ǋ�;���~q�R}/���a>{� ��8dt38؍Dr[�����1x7�߅�۲������n忂���pX��㎾$��u�숥�#�.�(�G@��yb&����c&�g��d�S-%��R��:������-����QLTzFنz)��h���P�Y��;(�������l}��"3
��'�v2�9�}á�^�7r�q �V���N�9֎/�W�Ί^5��Ыy�Ȉ��5��7���Pvi�hG�{�R�����1�`ؼ�>���9�狖�R�K�"v/_�ԕr>|+���c��˱:��D�Ϋ���n�N��+����3�w��<n�VmS]t#x�Ėn�PI���Ūm��xk�9�<�= �')8�ۗ�yrݞ���Ly�}�����;i��Ȏ	�39�>�\ wu��yj��f+ѻ�k��ؚQoς�f�2���ELdF�&�ф9ȭ�.�:���3�/�H�i��w~N�7V(7�ܧ����#��F)�G�����EeՏ�
Lh�Wׯq3��͎Y%��6Yݝ�E�DfrCq��Ie�k�r��bG����m��b]��Λ�C�Ke�Xu�Euj8�R����с����ۜ���{K�S��,iK��Ξ��ja#�U��s��L��uxy�e`̪��x-�*��ga��/R�
��WL(��^�6"�j
�Q57�V�/���%5dX��ӎ�q3#���:��xO��p1���3�"�Zll�B��pD�mh���ݔ���\sԽ�W�ȵA�H�i=���U禳$�~�|+�;�,�F��K�����]���ʰze��aPP�qNCm�Nc����J�֏��{/�@��vױv��F�k!�`i��r{+�'}^���Ny��7;�2Ƽ��a_/3�d�����y��`�wp�>�ִY\E�y��f}$[*��gTc�,�D�ղf~�Nk��'������,�>��ι�"@�3S����29�&W��g�m��a>���\M(��è`�:�g$((���hRt��+0���l��1�=�ԥ@�j���d��>�/[�w��Mk.,m�FAxOR�GO�F���dWs�;�JE���Ŭ5�"/r�ă4��hq{%��� ��۝�F-L��p����a�':.3�j���-Wk"�����Z�ut�ٱ�	��C\�j0��G[b���D��9sN!'צPѩw �M��֎t��J�n�ra�+�u��m���С���d�w�*�e3��X����MsN����7��R*�,�fvv��i&R"+��"�X��8����nYpWo�k$ ϯ*v6v�m�n��'��U��ϕt���}��7Pk���vk�P�r#�'_(���;�Vˌu��c�!�~���^lNw���a=)��zE�B^�ϐc�Lчe�u	ʦZ�;��xxd�å��\q��	q��	1���?,�خ���j.��L�-��\.�x�==���m�g�3�M�_OЏ=��-2>]��0����܂��xuX�,��q��kvc�[ѩ��l�t]-��=5z.[�)?�\V�z���'�iY���wu�@��X+�R��G�Ct'�8�l�,zX�����^T������-����gx�&΋[K$W�a�]tv;��Lw�L�5��;{U��b6���yS<��S���'�����4��ժ���tE�Q���VV����ʨڜ>�~�9�
={��+\�׶s_2���8��ڧs�y�%�η���!��2IO5��#������uI��6.���3�}�VjZ]�3t�]V��������S#U"v/B,^P��|y|��z��]��烌�"�X���ef�qZ˙�E����s��ILn��H���֫���b
C��[@�[%���)vA!l�&l�������Qe�j�˕�N���m�>d*Q�:�}{���sU>�u���̏[у30�K�9S���A���(�������HWm��0���Ժ���OE��N�l�@�6�S��=�y��p�����2�I��K��������a�g 4o#?L�:�̽��H�>���y��74�u�F�Z�mT�5��Ԝn�U��T�P|����v���/����31�sU�X{��Qՠ�HC!�P-�ҶL�{��z�v�̬|�����5�du��rU�dl����ݏF�95g&4�C��=X�t��|��Ʌ�o�{﫧�t{�߷s5������J����j�9��� ���mOa�S���A</^�E�>'/�ո`^�FyZ=�zWO�>�z֬�zj�[�7������	��'��l���ӓk
9�d�J��]���9!���7��"�i��v�C휮���r��Q6�L-Qǧ���QёVƫ��A�nM��:	��W'� ��X�����p�������� ����:b��:|owk�b��/+ѕ6E4���u�c�)���t���FoS:�b�|mڀ�B�j6�����L��m�
y*�Dm��:l��i��'_]!uv�vh'���x�+�����bE���hpѾE�|*b�W&y�tYm5�z8��|�q�|[��Q���۹n��ZK��q83{q�OT�yj���R,A��mŻ��$r�]��O��UsA�)L^�{'S�û�<���0JwO0�EA�^Gk�Y����NL4�s{�v��q�����J�]p�2�%Ki�*�KR��_*Y���P����3n�Mv;y�U����ى�z,g:ˮ�}p�ꘫ
���ʰ�W�Աɱ�n$o5��"��:�Y���]�:ƛ���h��h-p��t���M��m 0���nd���k��d6�A&P�Ruv
�;�6U�8y@x��� �U4�+�nޙ\��nw	o�yO �d*�U*}EV�d�3�A�K���3��3"�Nzׇ���8��l���3��Uͮ��{}Z���y��q1MugG:fjC}��L-i}6=��ñ-��UݻsP�[x%���y7m��1K�X��4�r�D���&3���EW�ދ�x_o59��e�s��U�s��n��&J�A�g��\��nw�'�j��˕;:�c-��<Bo�`x��;`	_7v4��A�ؚ\��]|���2k�*9�R�h���|�n��õ�TOCCchK�v��]>���Y-�r�S@W���21ݬ�&���bw�$�˽N�٠gM%u(���:�i:�1�f�aN,y}�1�{�tb��u�iP��VokI�k�#���&�nZ�[��ߡA_'j�l���j�ۼ�N����VY�Rk/9g&�S��o9xsꎮ�R]-�N�J��=������*qN9f U�Uך�V1rf����au݃ ֔&�yAP։f�3�nJR��X�j�]+X�x�^bw�J-�b�NJ=���\�k��m{a���yX�(s%`U�T-��-<Z����{+4Ԥ����F�Y7�bVj��@c�k ,ӗ�Z�I�y�+� �/�"�P�0"������>t)�OW練�Y�6�,�MIHPv��.ⅈ�,�0��4��^o-Z��sx��#�2��έ+�52�gM��]�ZC���v�ħei[�		`VU��zt�v�-�Ya*�r�@p�6�����!�V�ʼ�}c�z��\β3k�T%�{�:�sp]w�����2�VV`tNe���oJ��>�f��t� +�_(r�լP�aV�;�-�w��k:0����;y����m��/��Ȝ�y��;��n�0�Zu�T�l[�+2YOo��e��a]��ZjA}���gI������ Y�q>46�v_�2�8S.v��r����t��Ӕ�f������"�]�ܣM�9�)'1mw�e�f
��Z�:���r���k4���]�SM4I�R��6�>C+u��/S"Ν�����|�����NX�S�����}�ϔ)2�镲Ed�Z���R�-�qT=F�nN��Hֳ���r��Ǜ�r�z�Açu�z$�>E�'ڕ �7�����96�ו�>��6�ʁ�ӕ���T�^�?F�q��^L�Nt^]Fn�;:\U����;�����U������!�8�{r���Qߊw���d���ڊ��ez�}Z�_v$r�K�B�3 �Ѧ]�(��K驑*Da?p����΋�:�m����X2iUjaO��SBY�7��b�@uR=\=�},�?-}���3[���uI�5��x�A���[��S�$�BȊ���Kr��9�������{a���Z�«c]�_^b�x̔6��r�z�:�"q�͉�Wz�j�5�����յu���Z�Y6s��klk�Ȋ."BW��.7�ba{���峐���]�[�Ak�&�˴^,�v=}�U��n�8UMd�<�Td�EL��Z��H�8��ITF��!��N��J�YF�`U�p�,�w��ΆU<�a�@�T�÷;��5���>�͑�<��>M���̙���mA/�����=��k3:�ᣳ$	�GM���x�$�^�57�g;����H�=��arey��Ș5�m�k1�%rm�^j2�ux�&B�K1�s�X\���:a�E���̬�335o��{6�X��Q��p�[H5�2�Ud�����a;uf�P�쭢�  �:VGxzw	�s���zW�^F6��R�ή��U��T��1�A���y���+�+��i?{}�ϫ\�S����j�g� m)�{fXy���YJ=�5��~���Vʹ�0�1jY"R�m6MO
�grvp�r$M��*/!]�e^��������+VFk��&�{f�c�S73S��fg}�%F����5�O��zjz��s�<C���K�;�|hm�uܵs0�r^n��te��gk��w�q��,�H���m�]�I�~u3S:�J��y߯�[b��i����α{�Gn'�Ě=�ࢸ,>�L4R�)��0���e��1�������/�<.��E{��t}�,�R�y.Ї��e���6&�x\�ϢLǐ�+��n �w�%�QW�1`�����X�綝[s�8��Y��^ƂW�i��[��sǼ��
��{�Uw:����h�C����;v��}嗻��Qm�)��hF����c"(�U)���n����z�F�}��=p�j�TK������;Q0&�5� �;�~/��.��ou�3Rr�9Ize���n�:�ph�Ndӫ�-T�Ek o4t|�fK�eM�b����6��Xk(����n�G6>���{O�8�I��4/�b��X:ͤ;u7;k���f�唅k��{���sY�V�����݊�����Ze��`�R%���:r�.M�[
O���R�k�'���qN�o*��{��M�^^��3 ZAN��a���z����������Z�/��ɚ���.�qC�u�ˑ2/=l��+r���>�;�.B�j��=�B#��7x?A��������~�S�\�c=�㸊�[J�lߪ�4�͌����FgX_�ݗ	���sr~��b菉 Y�,[��̏��'�1Dv�;��{7ϔ\���صS��v��,I���2��p�_��B��w�U)��!bM�zZ����NӾ�u�{J(��6��O�Ng��3B�mNe39�Di(^͜B��H�,@}�4LtY	<�0J��N�N����F�>�5�D7�����^Ly�{�~u�<(TF�m��*#�P"H�3�1:	�)U���ln�)ש���k׋β�v��~"߂��BgQ�~���G�}�-�Q�:碊�����/s)�G���Yv�^}��ϼ���ny�:G�ըeE��V���M	\�Dx^��QH�1��>tS�o�n�46��[��J��y�+QK���ƉT�F��Ҫ!|�U�� �	_5AgoSF�ث�t���ٓ��S2���t�|٬%h�(^#e�S뵸���ˢ�.xszf=I�Ě$<[q��9�^����3��>]7�F_F_��Q!a�ݫ�&9vK1ߧL-��̑��=+�*h���7>�W�Wc��R��]XOO5�rdg7�A\դ��M���o�Y��)WB�/+xL5`���&wmNL��fV>]�u����<��*7��f)�*���Ѹ�y���H�^X��4���TL���Bg]���M�.�鑩��Wz��k P�M�FJ��Ŝ���i��t��w3�У^�9X8L|�=z��ٹ�~�Y��b&�����q��x�tzn+�fLV�æ=�=��[c<j�i�y����8}T��n�O@5�o�s�4�m�N�����	�.���}���{J^ȁ����1�M�塬-nS�ݯ{s���_���5S��;��	I�\j:q�<�8��鶳���(��큶��]l_ܬ��O��u�d�v�q���ف���i�D�]|�j����:6E���)q*��<Ƈ�W�b�r�g0�V�=���wm���fk�2�=�Er�v�^�Q�;e�����1��c5DS��n���*�/�uaZ�q���U�0VѥԊD��8���|2�P��옴�q�"�j��q�Rf���z.�w8�g9��f5oC:�좫{?��{`�|��<{A��˃��˻����ζ:�r�=�2�����i@T���z�#"�W�k6�F���t��m)#����`o���6-D\�d�0v��G���os*a��2�;nGb�y`|�+�����8�s�_��s���7[�ƞ���x�7k%����=b�m��E��[3����n%�P������W��Z�w��a����^`|���p�����|���5<��TOy��]��;iڳ��Y8��\kb��u�S�����{dpj"�Q�mY��~�+�ҫ3/9����<�cV���/s�>�^7~�Oa'}��cfL��+;ӽ:%a�-�*��]����\��.I5wא�EF��j�=��;�&&cnac�E�*!yu^�\=kx�<��?vd��y����v��h��f��:6/(��88��H���@�+)z��ǣ���z�4/r�C8����9�\�oO����Y���մN�ѭggd��ܮ-,���������#�(����{X��1�����F˨]���aQZ�n����]�wPܩ�X-X��`E�.�~�t:���5A�s�;�����#M'���6�ߚ� 2��6�e�7����ʑ�j��9��qΦ��f��Q�0m�^TȇWX�}d�Y`�W]��.�F�p-s���n�w�aM��؍�N�����3���<YV	��{J��]6�-̧��ۺS	�euhDծvSP1�2�@�3
|�	ƚ��َT�`i�Q�=Ai�%�]ܙ�k|F�\��{��s�����Q9Q�Ow�A�Jq�eQ9���p�k�n����p�;����{l���Uz_k�2za����(^P��pi�6��}%��N�*�SӴf=d�d]G�o��-�����.UԹ�w��]��}#N5_^ǧE=��K�:vlu�j��\�C��}*�-#6�ą�q��AݐԮzǏ\tq�f��D����{��<ș�y\)%��׉Q�ǈ�Hp�w��#x�y]Uv���6�tFm��"u�����uк9i��#B&�\��1ބK�dt��W�=�[E��;^Y�)�nI�̡t���xt.����eQ��Q��4�$��x��B��'j����wA������2�c�/Z</��D�ķ;_MA>�,ZY�_"�Y�7AF�*M�{�m�W����O�i2�B�u�r��'/�79�Ls��]��n<2��|���P�����
P�wV�⏃a�����b���]�{#���'�i��M�o��G8*w3{�v5�(+{*p����*�ӏ)k�U�����O���Q�9���l}Բ��U*�b�>�P,B`JO~+5h��;�bٔ6$,��W���7�/(gr\r(��ةԓ����@��=�ng��gq���~\6�����qԺ#c�Bpl���v2	��#����ƶ5�xy}9�c#κ��W���&|Fͧ[@v[�g������-�NϦ�J��!̜I��U���9�9���֔ǣћ�6�B���x��53ϳ*=x}�tDMm��aS2��{Z7���фx�Ħ�e�xח�b#~�]�u�7T��PSpnA<2��nS܁	=��.]\p�#]\M��o�aF����%kkQ����ڒ�k4��GO������\�����t�N��j	=9V��Fu���a�A��({��!(�;�];D(E{��s�δ߲���lsl{Έ#ݍ�Fw�\���������PP��Eϩt�z���5�}���z��i�gEC��v�_.�n�p�!�CL
�53j=���Fk�´d����ÅuW��r�nVt����X�����5+Ҫ��}��>�t�k*�)S:���fvU[u,�_
�B��Tb]�8�JB��tW�uܟp^x�Ȫ���{Q}+����+�i�mE� $�^����_�>c���|@{mR��	ĕWM��΃��輿��4'�$ٔmjv�\:wmd4����fulӱAQ�y'6��I%B����W]/B�ٻ��Z�r�w,t؁�ӫ�*�V[]P�j&�(�g^F�T��nh�8�ܢ�_R�r)Q �;н�������:�`�<��>����WU��UD�F2�|N�\�?5�ʶ%��Hb��׮��/��mza�Vٟ�b�{<�`(�������_tN��1h��ױ$ý�_J�Kr���b�Ps�Lc��c$t��B�/ڹs�p�^/:��ϫ0�w莄��uܜ����ZP<�n��aǩ=[f5�#�R���uLq�����WlF�J���k5K'(jc�]ξ�#�(�oj�J��^qIw�%����}�2�v����\��Wrt�u���P�L�>�yU4�c���Mtm ��cm�ֹ@Y��
�U.D�O�^�2�g��w����&ϾW�������ꆾ��޼�P�lR��d�p#�U/Z�����<�����>G��Bc����7��֝4C=�/(t�}�i�č����'i�a��M�
�**�]UѨ��$U���7]s����]�IH���ٝ�ឌ��&A���q�wb2gj*r��F}^���l_&�T��9�rw���?,�ym��C�[��Ї
[[x������UG���!A8���KhB9��,��Y@��EZӑ�3Y�^s��=]�������R�tlڏV��^X�j+jM�d�@bu��ΐ���=#+������%�{C��\;���=�1������3z��������\���+?ވ�{�p�j�/ ~�Q`�
�9�y�e~��s��V�aG�\d��ȕ�mT��îI�˪<0�A��u#N�k�e	阭�/�o"�I���D�?H��x�^ʮ9EL�02�J��%�u�O�戁����W��2X�=��OG�΋b��_=a�N�bI8���w!��(P�P���t8­ys�"T��7����/VT�ۉ���7`G	��z�B7�^�|����ч��{�tL_p3��-��I�=,'�^?,�]�yq^T'Qc\�M���dzk�<���F���}
{T��'���)��[PT{�����h��HŰ��^^���}|�#���97$����^����dG5�]�4�ӷZ#��l�f氉6t7�����Α�����b��=�Ӟk�;��=�P"%,���������e����"�&�j4��W��xmK�L�:H
w?�u_��}[7�����i0�eُ��$G�6-q~Y�#6RW?/w��*/o���ˢʳ��y�!���wJړ̵E$%�l��pT�re�]g3@�[��UsO\$�κ�EwYzz�Dі��8��un��l<�IR�-��h��w���	C���� ���#�8�����Z׫�]A
�9�,<{8�m#���30�sj@]�j����!a�3�de���J=g�5�m���˜1�)}NAH�����ۡI2ȍ����Ԭ��5�����Y���E��G�V�;}��Zػ��繸�WgN��Y�=L˺���̇�ѕ~��ux) K��#�����5�9	�+�z�rzP}����g�w�4^���¬��Z`W*Z���FT(�uh�|��z΄�y[�����X뇣f\,�Y�d�����i��kS��L(؂��P�=���JF|oHX�7�ݞG�~�e�w��i.V�xUs��و�#f��	z'<�m�3�9^�:~���W^s��GP!v�!>��D�<6U{���.��{�c"!�S1!vh1���v��c�bbZo3����:���j�Ӻ�ۖga�6-�F�0w�u"{�Q۾@�5[0d�����쩘�w]�D7!G򝎑�-�	��&��[�u��]멭����߹��qyҿ�̨��� �g���-��:���T�n�E���n==�˻^��6��.�� �栫��ͳ��>�FȾ�}����Y��9�����I��[1J�V�v�o5и2]��@�;�� 9:�򹍮�e�vS9-r��A���nT��ų����e�FL���hI��򐭕��0���N�7\�e����6֞C�&����&&�QK{��s�e���7�z�Mg��+����Q�u#Zt˶�ԃ�:�Ƚ��Ƿ�hY�U���֓��O�c{�NL=��i��2���t�{�X�cx*�Et�o*��ڵ��vNofk95�K4��gٵ����Ў�dO����G*�u}B�+�b��-jf�׽���%I�
F&I������4���~^�4��0 ڂ��6cu�7fR3yUg+YhDhP�_P*��	�iع����ӌ��M��ꮴR]�C5�B��+b�^ƅ4��[SC�����a�3�hz��E��}Mŵ����}�������<2n�H$w��o�ڏ�PdFE�Ju³@�<7�f=�vN���b��T�q��Fd:b�X�ep�*qACy7
�y���v��W6<�z��9�mP���X���6�;�x�o�.�9qn�o��:�ծ)q걄��0��CH�:�$�0N��h�j�"���7T�[W�;�S��K!ˍ�;sm񕆸póe�Ll�WFf�����{eJ2LiIي���8�ea�gV�m���Mnc�`�B/��(��`�f�����Tu�"��V�>x͵@���sr`�}��i�gIS���*b��ūi�U��ӻ�Rj���$���_oV�X�$�uk���ܦ�%[,�����*�N�2�jfbA�6�@o6_f
�ؓ�[�]�X����S�����g� �w^���`U��"�{nȄԩ��������a7�jv�]�S�$��f=@�������b�`|^�=}���7S�Vb5.�;�,B�x�8\�m��zwa��Wq�S����v���#K:�4��{�eH��\�g�8�.Mʏ��6�ǃu�K���K6X[]&�->Z]��ʒxJI;YY�����@{B�Q�Jk�o�"�D����EÝ+-��բs���#�� Y" ��Q�-�g�s���2R�.�6	�	\y��0C��u����N���ū�[Kc�|�MŹ���J�B�2�t��L30�i�e�Wn�i�Mk�ౌ�e��L)k�w &�i;� [5�����y̜v&�h�~4+��[@=jW�V.��.	�BZZ�:ǔ�gm�uֱϔ�	��i�n�e�u��d�w/��`,̀u*ʌ�O��;Ouٺ���o����*c���%�p�%"{�Q�9�X���y_�9�ܮ�뫆��k�.�s!AI*ɐKf}��|�dF��Yl�3?e��kt�o瓾.�@�v�^[Ϟu�<�.:���n�g������a���@��ݸ��ْ�r�2�7�jX�;��D������z>~"8�D��Mzd��ӝb������u���f>��=��':ㇻi�����0wvB��:cs%��o�J�#X�3��WS�ښs���t�Y͗��{���-�'�v���<�{/�G��i��.�P�y�n����O�	�Y�*����7��Dt�-3x_yt�"�Dc�dX1>�z�G����I���r�L�D����󻠷��A��Z3}�B�Y���б/{47����z���]l�_�W�C����B�k�	��\�RF��rbѩ�%f��ڟV�N�{)m
������g�u\,��):���ǫ�9L��Eu�nw&�|�����j�$~3�~g�_�K=����c�;�7�TH�W�S���碫Ҕt\l����}���F>X��~���gz��Y`iច���U��1	0Z�s=��FggѮ��T���&�SuUPLs�ֳ��6J���K��i"*�gG�F�1Q:��5=�_��>��2��6_S��w;^�3�BY�r-n�TI>1�i��Y�����ye���e�ƄCv�1T1/K��+��[�uU�`�&x{dvO������oNm<�ɄFn���cR��@��_I/���X6��-g�.�Q�������wr4��\ܫ�fwj�dmٛ����i��怾����m�"�E+�G���;�{d�#hn���;��j}�*r�O{���?vW����2�O�޸j��m��o z-��H�ѷ�莼��3e<)vIgӔ���v�)N��#H���hp8l+�F{FG����uI*�؟�B@j*5*8hq�y�-��
�Tn��sR9y�}����:a��}�l����}�nx�)�b����84��K�F�M��5ˋ]��/2��p򀫴��W3]T��f^e^�Qj��D�^\d��x:A���Fd'=��b(k�t��8�ӭ���&��W�d3.3�ӱ�龎>��ް�8@zy������Ӥ�@�����\I���w)RUkw|�f��޾z��7_���Y�Ҩl���o�1X{'\�E*��~ʯ�~.$H<�&���;^lT}�4�����S|6v�H��-���E��^k]�s1{	�ynkw��b��>�Y����QF[#�^�����bS�<穎��%��->W���o��GwN����~2���V9�!�0�����#{l+6�*v�S�U�:"�8�9���vߵf�F1�xܶ9I����%��wf�����ͷ}lR��L+%����c���H�R�c��8� ��N�Z�7��;�k����7e�I&�oq&Q=���&��x�\�<
GA�>icZN3�K@��A{ce��$���G��?L��.wfo\�0�n<�v僨X>=z3�^6'�Ƶ��}�z��U���ɤ�eOc*UF=��yY�zmC�@r�>6.�%1#\.�W��Yz�Se��mi��U�S~�s�xR8�ɻ��A�\%Z��ۢ����P��(l�B��^�=x��G�ɴ�_WY��r+��tl8�[鉜�ΤA�����ǀ��l͠}M5bGWr~Y��l\e�����Fq�b��BI�h�y�l步{�a�C�ع֫m�Kg��;85+蜷�Տ���#�C��t�lA�&#":���7װサ���&{��/{^���m�疏O)[���=���)���)x�h=��W?����
7lB''k'<>���[s^"�b�W7W�.\z��t�㠕N.���f�۵�A�a����<��xtC�x9����:��O�]׊��\���3�a�����˙��X��;�PN�ݿSk	}�uq��7��|�Dϑ'p�����Ӝ͝5ޯF
7�Og��S��$"�o;�nhnP�=>z�Č/�$�V'����#Bw,�
���:Rdd�v�����Be�l�*���	�*坦9%
��!WLu���)#�wY}W$+x�hr1���MU�}eݲ��\�Y}/6�`�
k��P���ڏf�uE���ܮ�o�۳�fuT,�r�M��T��D[�1�.�,W��ȹ�׎��]�t
�l_��Nz�<;���Iq,�kH?$"Q��#,꫾���Ȯ��#)��^��=N�/��g�<��R�6��:6+�"���\rnDT�� �̅��=A�;s�]�ޟG�n����ܶ#Dx-Ÿ|�.꘲���0��T�𨍺P`L[~�){�(����<�����9?g�S`�7P����}K��7��)d��<)fϽٝyNo<��6��;���@�^�|;�}��i=�zd�ݾ�E�i���o��yb���>�|�FA�i�z8�*��#����U�d�Y1}3,���
�~s�i]�`���xh	�Q�;��N�^��X����;�aܨ۾��z��=��'��8�f#����G����F���{z��ˎ�)�5�������G��ѻش��o;�i%|�j0����y%Sݶ�[;-��\hQ�4�u
�Muⵐ�����.��+�s��*Ď	'�YD���2�ES�E�����n������b�Nd�6��%���}��U�����oY\��t��"�$��_�P���:�R+w�\ڶ>��:��J���%�-h5�$�}rK9�ܘ� �;�6R1�v��;����Pޤ��n[���>�*���r��]b�����C��y��
)Ǖ3�������̡C���m�kC�n��yա0�pձ`�����7�תh����u^;�;d�9A�Y��ĸ�Fs�Aq����*R�p4Dh��U�L]c���zj������	\u�H1+b��je9�77�/TH3���kB+ئNcyn��B��x0N�xVv&��j�u��h-A��ރ���|��eF���`��a�9������ԞPto/�vO�����#	��t��G���uH��ޡ�h����go��c�k�3�ɯ(�g�����_c��Dm�г�x��=�ȵ�u?CG�����`)�}�#�2��G�E�׿����z�.#t�[��n�h����^��;�x'�Y���4b���g\�7�ƽ2�R~�Mw�"p٦�Ȟ����j����[.l���2=y+�`NL�\���Pm�S�&e��*�nhOC��e����c��4�q��g�.cT��SK�8<�uу/\E�z 髇pwٓ��Ŕ�0�	��|c⁮v�-�{��rc�i.�>ZX�n�x�B��-�u/9�[��&���bJ��[ ���\�H�:)����:��U5���/����R�RB�Ʋ�:t�4�>�[I�t34e�zoП���I��M�Y6��GL�����d�{^�S�3��҆sp�i8��91�p�וr#�^�z{ttn�ln�&�k�~�fP�d�Uw�3G@��s���C�n5�.��"��cN��O�Ł��Ax���L7��,!�Y�;sf�݌xچ)3߻lx�f���\��|(~��:Uf��W�ǺDԦO�K�kQ����|�<�cgr��o�VMaZ�>��~���Ct��������崅e�X*n�1���zj��O�M,��x̝Q��8��.3�����Ή��9��7���}����IZ�w�߶�ݏ�[�!	��	О/$c��>3͝+�;��/�ȁ˟Tp#)��Z�oˤ��u���5+.X��}�?��''��jobC��]~l�V��k��^�>?Q��4���Pvn^X���������>��&xQC�ͮn�Uvu�j��Γ�k��|pS�c�<' �X�f��ܜ�u���a�ÖK�ގ��(�(*h?%�|�ι=�N��'
�5uk� �fK�M %.����fT��&�JmS�P����n�y�B���'9w�pn�k��η8d)}m,3��Y�:�]�V����tE?���8$��,^�[)p���V��̗��򻎂��!�&�#y�F8SH���S}>���)�����1��c5i�^����t�:Xy��ݏ���s�Q A������7�WoW�zxU��FmL/�m	d��E��ϻՌv���4�Z"yv�B�g CWk�/����k�-�t��:nd��XO��騮{#'�w��DU�D
��eQ�� �i�T�iw�s��Uk��X}��]��~�Y��*N#i5�A�&���6�8UGP�V>@�]3�P��йW����^x��wsre�*i��t�����҇�ӱB�e^nP��x�<M��\���j��.��s$)���P+[|� �Z�2Z�KY�Ѝ�Z�P���1�(m!����g�y �[{熲��`�-O_��(��=>�N#d[���w�@~Ҝ_)����^���ON�7F;��R�o��m�Z��0����o��9)
��j��ǈ�"ӣ�Oc{���ֺ�d�89ļi(W��h�Q=���F�`����îk�w�����MuM�f��\w��x�'rhF"��Z���-�ݬ-e����F�e�I�ݴ���^��_r`vxm*��hXod+vūa�J��6�:]I�H�ԛ}�82��)_W�;|���CΆj���<�6�a"J��O\ŷ�ɋ}�p\�_v��7�a��w<x?	�/����S�WC�����,����X�;+�������~���9��Lxxx���T4_t�f�{@���2������}kDέq�.��u�=�e8��S�B�"7Ժ�̎3��/�T�om3q2 ��!��r���âGU��:/5�Nj!���,�~1w=U����{"a�����%cL]��G���t��;(�+�-'@��S�C<+�Z��{}�7�F^��H�r.	�v�c-�ъ��w�rvNu�(���s��c�
>H�#`��s�;
�u�E�Q�,of��ػ�}���+�袻xfI]G<���B�kf ��מ�:|0D�e�Y��1�4\��҄�sR��G���{��L�X�7���
��>�]�A鈈��mK��az�~�F�R�n�%�R{�='���/��v���v�A����:���<6��,㾁����ݝV�Cs[~�֦kՐ�wٸ��ڶ勯Oz��º*�wF��i;7��8E�k�"B�����C�r��Ǘ�.V��GG�@o����8�on]�Rډ��'f���L��38Ճ�P8E4��*S�P��6�u/r�;��:#-��#���`b�s喥���^TGeY��B�iJ������`�4dzhs՛��f!�3
t�{gnL�#s�<�}k`e�9�'ڂʙ��_h�ႅn���CLd���`�\'�U��B��q��E��e�������aj�V}�30I�������d�*"O���:�&�/��|��d���������l��{ɰ���TAZ��߲�T��Ɍλ
��$��C\����:�!]�'X�����Y7v�0v�}��)��s'�GaG�P��59�;�!�Y��]�1{ا����k�����M	�h�Fb��Ȭ�������ncA�o�؆z�!�����ؑ�,�wVƪ�#;�]߼��w&���������:��^ޙao.��
,A]��5ek+�تt���ӿQ؞2�"{L�n&��b|nF�b�N���n�o�X�1�g=�=�^ާF�~��<ڰ�����z��+�:#�T��"qo"{Ϸ��ʖ��������y�xT_(� B6`����]��V��}�{A�F��.���ۉb0�B9v����FǠ8�ֲ�؍,/��x=1��ynrJ�'u�w"�ݜ�}G��]��;���ȍ�Z��|B�YƱnnm��-�ε�L�Κ���u}��w�SԎer�3OT�Q;��x��K)�&��Tν�Nc��JK��j�ٙi��Ş��S��A�^n�x��5I�u�	�0�gP�{����۽��pA:�d���ߞjɺ���}o�0z*��S�IU�����SBz;Tel�ٹx!U�y�=�����.$��L�NmK���m�z<]�}�U�F���+$;}n�*���P.�����/oDn��;Q��!r�����0]:�}�nR
-P�Op�]
7p��=�Lu7����j;Wo�9�O��|8�W�
�>~���J�Ӵ�(]��⮀���޻~��M��+��z׎��{9Ȇ�^݊�kOLA�)fk�q�}�X=����e,꺭�D��u�ͣ�-�����������\�ab�=����]nỺ�B�Y3G����L�-��y�Xw���bs�=�k��n�[�!+�����M��rкjH#(/�_�h���q�/L��	��v~�}��	A|F/A�:7����!X���kx |��͸'/�P�ml����|���>`�7}��v�l�O�u;;���6�;����^�,~(�X��pb��
Y�Yʰ�����vސ�۴f�ZVhC"�&u0M�ں����<�Ē�r�$��Bo�r�R��T�Z3��dL:�ӖfN�qdQ����f�0-�.u�G�5\����Vf�Hج��]�\* �\-��m.�=N.W��r�	��9�dXo�ؠlm+�#V��{/ �;sB�ĵ��"��O�2�;w��m �W�Mg�ERA)9Z��4r�[xؠ����ЮCM4�Ǝ�_vK۶)$�X�z!C[:-��۴뫛�����O{�JT47Q�y������`#�;{QF
��t��q�\�/��gz��+�TP���
�!۴ �ւ��#!@��H�HI#� H)AATZS�
��Q	�ݴ T{} *�� Tu��5�=�\��u����Sy���ԡ��Ҷ���y�N����.l�$���U+jC�Օ��Tj��!\����5(�Q��ć���JEؠa�u7N$�B�KT�47��mӶ��Fމ�!�L��he�t`�]�ub��]kJZ�� FӷcH����
��3��X�K0ޫ��Y�odJ�42'��j���q���ٺ\&�r����T�rވ �5,��tݑ�j��$�B�#Ҫ�E[�f_��M�[b�V˥��� !��eه�o�F��U��`��J���;m9NU��C/H8e�i)��ϖ�1aa�6+]��g\;Zk�/6��˫�m�kI:F�����SL`�(ԭ$�m�&T��|�FJ�-f�4�(c��[b�K��������]�,��o�EH���&� �;LU��[.���FXg�V(0.��
߳�T�-&kf֪śOF�J�h�f��YNn2A�P'3(�u�B��ہv78%���˅�[�\�c��w�ҧ������hT�W�Jn�f�� Q�r�^�7i��6���!_a�t��8
���E�ofj�6�WgJa�)Rz���j�[4n���AŪkkw:^��g���2tӨ�y�zɣ+�ԭ��@�<�U�(uP(m\�Im���Bq%�ZrZƤ����Q��3$� ���/U�i�In)�oe*���(p����6�K�l/v�����݋�AVټ��B��������N����<V��4��B7O/-�4Զj5Ad+qҼ��	3\�gM^uL�U+�����*�fM��*�b��Q��7P�g1]�"��q�0�6{٥�������-�Ik�����m���e�.̥P�p��m��`�9�'I���Z�Ӂe7�U�ݻ٩��5f��U,�e�)�3Hh��E�!�	V�N*�lܥE���Uܶ�d���Yi�Z�k�Q���[�Y�
��F���\Xs9N�:v�@;͟%�5y%7)Wy��E#0��
;ƒ��!��#���c ��ow�3f�E9j�أ��bf��sk�̎�(�٘�"X�T���@R2���g
��Y6�X7��M۽a�(R�gT��̫9ֻA���@�Yi��:��5���Wvb����!n�B�#�k>)�oUD�2�kl�ON�)��C[�R���+n۬�Y���%V�� ��i�J�[�I�6G�S�@�n�����R�U�%c�Mؕ>32T�ӥ�t5
Bn�&֒j�A!@*�*�N���aEx�e%��l[*��[J�a2��=�e�)�&��5�ݨi�[��2�hV�f��A0җF�P��
��U�CZ&���q\ö�o60c�oD'j%���
:Cy��6�ˎ�Km�Q�#��6)�\P�=DḼ�[f�dlbC]8j�Ebc�%j�=����S"֩��C������m����Z�L�u&����"F̸Һm�؁c.�4���lͰ���-k;F֊��4,��f�i������l��Ĉu)�W�t�x��r��h���T%+{A��I��`�6�InZ��=�R�^*�P���v��C3+v 0$�emXYaK�6fjB��{I2D�����q�V��J��Ea���3Oo��҅�F��]a�Sܕw0 e�ܛW�`+),'�E�V����ǒK�_<�����k5 BF�kjܭ�aF�h�3-ͩ&+��l�0c�%�:�ҕ ح�������m���״輱�٠�S���B�T��)&Ⴔ%j����F$*:`ۙ��o%���5Y�-\lb�, f�޽����!kI5)���Ւ�aÊ�Xv��Z���k�Gh�p��q�7��zӡ�
�X˼(M�մ
k2d�j��S�%FK�S�8�(�-Z"�,��&^�&�a�V���*� �A�)��1V��Fi+ue@�\��A��a���/jT�`nA�2�sH�i )1g�3בaE��Z)&���e�grl�4��5rJ*"�R��@���f�[Nν��/���C���k�v��JVcFe��)�06��GA(�f��V��66�GO
Y���T�3!�ʚu�� #x�P�RQ��8`����!{+�q]YɃ�V ��"Z.� ^�˶��
�ʖ��ug�*$��ɰ{)�W�}{4G�MK*�7�����D֛�.��X�C^�խT�kT�O���M���Z9�[�o-n��+=���IU��w2��C�H�*�^�R�j�B7/�U�=��f
I��Q�Ƿ��U�{�t�)��K ���On��*RF�T#OS��H�G4�"1yug7.�܅�(lF�X�H���)17@ׅ�Q��ض�v[i�Y�oΤj���q�RY�[��nly�i�bmn<�(hS����\�0��&�E���U���ke*PҨ��1?���s!!�[��J�8��2� �9E��Z٠�=�&�)�Y�*H�U6�5v�\o
��w��,��MdJO&k�S���<%�`ϙY"�P텺_ŵJ��Ӭ���n�-X�C#����W/�5��{V��i�c��*!0�B  �$�D� D��BB`H�$�X@�2@ $�d$��F� $J�DJ(������(
�X�|�� T}(wd���P��� Tr �
�耨
�bj��
�GJԷݳ8��$P�@ J�TQ;_UQ@W��+�y�%|yY�+�P��kp�� Tx To���d�Mg��|�IY~�A@���@ ܟ}��o�{�SA�[�i�H�([m���+��l�U��(N�*��,��w�ٻ�+�B��m���  6UڅXm�f-b�FƪfͲfL��}ι3ed[5l2heb$�TQ[�1+ ���X���X[f�T5��l�R�mm2���     	�::dM*B�QUI(+lJ �v�[J�.�`      h   @ >��O<� @P($i����U��J����.ڻ��]5 �u���2�(� ��zvh�4{�n���ѶP�� ^��-ݜ�[i�(P�Z�cY*/��h���1�[
���G��Cl>��������sƪv�۶�g=�{ƴY;�������WJ��/sz��v�m[q�;�����ww��<xٗm�u�[=��]m��ݻ�ާ{��.����z���wj;7��`/'u��������42zf�{�JM��޷^�٩�ݷ������V����y���{3�Wn���o��]kn�N{�{�V��o,v�kmW1��tyZ�m�����sU�jj��ޚ��ܶ��ݴ��f���6��km��U�=�OfVڨg�w^�Uc�땨w.�u�V��{;���com;�;��j�GKyJ2J�U��ݝN�v��0��뻰�e����h{�l���r�P����2����i�Ƶ��[q�;�;��^۱���/o=ml�ݝS�׮=�sYiu��N�\���կgu��cM��u�[�]��ݲ�F۵N�u�������s�M�n4����k�f�Mg}��r�=������QEx��5|^޻n�=�w�wv��v^;�r�gw�^�/{����n���ks��wnE��s��չgVݼm��7k�����{mamvI]��-���Ǯ�z��Z:��m��m7�.�6"�=�l��5���뫴9��;�����n��e���Vm�ڍ)���w�[T۝���[ރ�Z���ޝ��κ�׫��os�i�������cvSs�{�۱���gzSKUl�%B��6�S7�w�ٽ�ۺ���ہ�����m��^ݳ��ޚ{'����;�R���:ht#��6������$���έ�ºФ�y�o5�gWXY��[���w7v���z9�F�ѫYF�kiR���z����j��Y�M�u��7������Nr�-��۝sd{����77N�#�z6��ս���mݗ��xQK��uև.�C�tV�뵪(�V�m�4�II��{��z��v�c�w���-���e��첺����Z ���ܫ� wIN�]t���{�s=�m�m��z���[kn��z�M�^��o0�=셯�c�H(�J��T�J"�H�$�$N O�&eR� @ ��FJU    �=6&UIH�@� *�	)U   T����UH   &���iM��Lj4�l���߷���������|~Rg�~ѴR��V���/7s��{-���������h@$	'��>�0 HM� @���  HO�H�$��� I?���HLB@�$�݄@��~�(
� ((�0E�Y,C�Ɉ����EFE�4�����5����sB<�1w�ك}�7�bL]�)�����c��wY�JeM�+B�Sr� �97fI�$���ZܗZڻ&35�Щ"w̻����oF�V�TZ��Ӈ4Y��f�<�,�WkR�yf�$Դ���~U���y@��1A�1c2��m,��4�Tv���r�"i6��&�x��.��	���@�*����i�ѧ��
�ژ����*�me0U\�^bֱU�K"˲r�XՊXoQ��4��y j�MrmLfv��\Ft�>��.�0�3ݒ�І�����o$�������Й�l���&�9-�n���]�E̅n�kRV	���u��kx-�VS��ޓ�H�o��^��ڇC����������N�%�Fވ�%��C-�u3��_3y�}m�μ_c�eG��(�UXw�#�(��TO0��IU�� ֨E�PQb��V#mb�ȰX(�H�"���y�sz�o=Ǧ��{����u�Y�x����:�Ch�jب��m��ER�[�ܫ���ݓ$i�Npף�/0�9>��-����ty+1 �6��q%eH)U�i�"�B�*J�h�%h�����N�Z�Mg�{��e��{��=�ì�y��
��<��^�6�v���{Ue�s��FR�Yz�Z�S�����,�y��o�.�˦�v^��[(�q`E��Y�Ѣ����)r�Q�/W�'��{�ykuN���u���"-Qf���{���,X7��9��9^�h/�ا�M��3ug���6�ѣ��G�c��m�ܲh � �R�$m�.���wz̽��e�W�Fr"�AQǛ�pv�f�����
6rj���LV��-8n4�P��p��m1��J��]�:��V6�vt���d�Aa��/v���K�{3N����ltʨT��Y �~��(��%�2�ŷ�El�����2)V�@���B��	��V�{ܫs0�Z��]�RI�y�-�$'Y4���k�)�X�b��L�L9#[�ܻ��H(�����Њ1N4nM;#WL�ٚҁap���0!w&Q+?��l�.4v���\�������(�Y�2ړ��lX�"b�N]`L1��mdUy��8�F*��
u�'�2-r��aޅV���Լb4ED[�3-��G47CK���fB��!ͬ Ŭ#2�y�ZW.�(���Am^�n�Ra[R�lk��n�	�a�Rz@7��(	����n4�kVF%\���mf*H޹@�y�\���DUE�"�� �b�T�hPYXV �R1X�# �H�cl��UR�)�,�+6��v���ʙ�PW���t�&]�*�
�ȋ۩Z̺���B�-�K��GM���un�� y�q�AX��İA���On�����^+�X�b�I	S�ӵ�j�����$�I!U��Q	ԩ �Ed�5!�,H*�"ST���2*�H�#`*�E���AD�E��g�,A�*���H
e�U/j��r���g��"��d����֠UU�a�Y�~v��/i�T�4��KVl�"��a�[i .�K��MMM���J�	 ���z콧�-M�8�A$��l%A�z�z7�4S��^�v��nS9V��Ì�n�Me$%�
w��
�Cy�db�o��*js��g�ٻ��=���Mk�&T��˟�E@Y�,F�H� lA�U�B��%+^�Pa'5e�ܒ���Hס���2�Q�:��i�+Ø��y��G�6�U�G�* e&���v���^�ժ��N�Kq�����QݤԎ�j�a�J`d%y��{u%�T�Sk�� m ��2C{l'7��{�wۼ�8pd;m1����3� �ՃK��e��X�0�
��Z+2+a��F!7�6�5z-�l]�F����N����ZHPͻš^��˗R[p���'�0�{�es��ٺ�u
K�Gh��i;,�5���r�4�0�E��g7Ue�l8k�a@;�3Z��U�sdWl�
^o�	�(�Z,]�iT�x�e2f�R�+�ߨ�UG�Q �e�̙H�N���Z6]ɗW�]]m&�j�=�[w�%�rR������m)i97?�iQ��le�?~Yb���/2#��Om)��Ƀ�����ۑ���T�J	莮�~P�Hcʅݰ���v�h�mlr�Q����n�!���؀��ĺt@���{�Rv* R����۔�l��j�2
hV[٢	Pf����*A�wNX�Dvi�Z�85	v2S��
Ŋ�D�:�M����]��s�g�}����'�Lx0)�)�`���(�.% ��`��b���(("VF�*i ���J˫:v�Ӭ��EюO�fə\3:aAd�8v��YLNS6^�_�K��YWg+]�ɤ�"���K2��j��/��l��)E��P+��vS{��9n�������G] 9�
hf��\���ò�;u�M�(��vC#tɷ������#��˶�f�\ouKyR�Z��uq�
#�kV$�2ȇ-ɺ�ٮeK7le�j��X�"U��R���΃ϱ�ݤ�ؤ�mv�����������^k砍J��!2؆C����o	,VӼ�k̒�?��.�j̭�N^nF�vuoܻ�m�K�&�c\�6f_�2�0�O*���C|�޴���²��\Bǚ�uy[v�:)��4�+�5Z
.�-�?���j������QY�kJM�{�,	_�w�Mr�Y4�ǣ2ȣ�����B���TD�{n��Յ�b�%,��NJ"�J�1]M�W��iҚ�kf���i8H��[V�����r�;���R�DBah�i�2�B���WCmV��{��$��g�H�V��-N�jɤ�r�k]��I���{��o٭b�����?���R��nD�k�5�$�ٴq�xwv؄���h0���tF^�(nc.����e�Y��q��:F�E��n
��H�]GY*��\ce'T�--ʼ��/vD0�3r$�ڢ��)��2]DFE@����+/)@
���?^[6@Ѧ�4)ӗ�O[�K�T�4���u!uGQd�Q�i��H���D�5�M��i��-e��bT$7 ��լժ4�Hr#]ŐC��6�[d��pʋ8q��x:�MṴ�BcV�Z�Rm��*��:��ڦ�N6S�v�c��H�Yg��p���-Aڔ2ӼcjZ��� ��_����c�5n���EQ*�'4�[�iݴQx��Q���"2�Z�6 �1�ݢ��"*�A�DQ�����eJ��oJD��Z&&�[�R�=dQp&�������]�yi�`�I�j�77Bvr�WeSbm`���`�/Z�A�AA�Kօ�,��2sJ7��s}��^�k������+��u�i��HBh��g4:旝����sl�m�Xq�U��)AI'�\�N�ٜ��ꄯ;a[��s~�5[8���^d1��k�z=�٭v���sؔ��y$�$�$c[���֎��G��l�tu����7)~�8�٤����CW���l�a�AX��;�4��D,�0��C6%�Ɏm]S/$�/T8�p�A9�*-�NV��:P�U���Z�lQ/T�CSI\X�ףN��b�L�Juwvb�V�%��w�2Hq���w27xn��	j�	�4۷~�}���q�c{۽6�ԩ�d6����{��T���o}��y#hѷ-�[�Ѧ/=	�D=�2щ�O7&7De�/2�Ӊ�E�-�����k'��5���dam&l�xM�_�D�m��Z�v;��7�%�����*;{Y*I�aŁ��U�U(�,��J�'[��&G�0����9���-�B����8Y�ņ���X+.�U��̣�W�X �zɖR�x˩�^�&m�\`�Q�ʶ�=��
	b�86 tf�kwb��/ɖ�e��w��Vm	��FU��MV2M�J�����_��K�/kpYS2�`�`���szމǬ8�k'Ok���i�{��5������cm�kr�<�M[i�iv��pS��O.^�H�+cQ����Q�:�~�u:�IGu{��/�'�4f�����3t����L` �{2v��Ӎx�{�s<�-����w�,��Ĝy�o;}��!�La{�������Ն��Uh��DvRVu6��T�d��^l�Sv rB�]h�Ys+*��eK\g6ؔ^�01�PW���W�8(7�EH������?U!_�Cw�;�SkAtpݜ��~�9���a��no�8{���g5�T���ºƿA���j2t3$$+�����r�����h㥃QLK�y1�f�R�X����R�G]�o=mV]~���/��mb�ted8I�ʠ��(�ݢ�+b*l���ֶЙ{r�]C�Zݠ���m���5;�*%3-U�2"�aDG7s`�������Q��	t��3+Na��S�J�{B�ڬ8�D�ƹg𭻻
0X'༛�i����2jl�SB���ʇS�M<�^���֝�zn��9���7bn�լ�&~���`�a�X��b�+)����C���ڰP0;ee/�sJe�{�G�u���r8�7�R�7��	.�����-b,�`l7�i�(��V r�dz`�Gs-=���+U�VóF��bUL�U�ԭ�A~z 4�!]f��5[B�0*V`hٚ���akN@<Ҏ�X�"�6���f㙢d����4�9h�B/-����n�;��Q��z��$ �
�Y��7�Ճ{`�+����=�lmC �RH-;��|�x�w�Ab�=y���{y��ЫF��BK�m�����ݸ%P�sZ�F�D6��6]��7De,�(;4�����{t̷LH�:�`�(EPF(
m��ȫ��Q��������d�%HE6�C�4��14vSp"�R�a�J
�@��B*���aW+h�Bĩ�(�H�eR�b�����4�n2�Ed�Y ��HM����!����x�`�ys7*�3H�AX�����u#u�X�=(���X%m����#Ɣ���!u�h�V�il���h�W�a�����c�Z�hEĚ�g��g}����׻�@�Eq$+$6� `�����H^�Q�"�H1,R$DI=eX

.!FDb���2e�R"�QDf$*, �u�n�{6�d�}�{��]��e������N����AE�T`
�b�D�bJ�DPU�!(�*��5h������Q�Tb�A�X"��"��$��*EX� ����B,+!X��X�0�%A`�h�*�b0T`��P�1�MXb"���,X�F$AT1
���QUcI�cTH��i���"�J����k*��(��eH��
#����ܻ�Zs��nE�D���WU�s������F+��>�C6�qL_W�YJùv)p�[�}��8{�x=|�o�4��i�8����V�Q]-�8��R�ӗVy�{��ڨ�.u��e^)F'���*�VT��9Q��t���Zx@��1k� Q<��=�r�9�Fo���Ը5��Y/���Z��^�W_���,�3��n\�4=�v����-#�Q�ȲT~s��ī�L��5W�G]�n��0ʡ����Y������ru��Vyv��'S��t`B�3��:���^�V�m�!��d�w����em��	`��5V:����Szk7I^�(,�R��tt\���h3��"�x�w��cC�	D��39����i�۳�U�agu�#bܲ7[R�IlኸY��`�7w�rN�Xծ�e���R��#ST9��,�Jn��1��c�c����l�U��e'G:jޔal��M3�o���닼�]j��t��2͂P#HEk۳Vw20���Lqc3��1%G��2�>�unp.�#C+�2_vѲ�u�
�V�1���3 �;����z[�,�x@z���W6���P]ʍ����,p��.�/WZ%7��/3��R�a{�{@�-w��ge�q@�ҹ��v媮�^
{5l`��y����gR�;)"����fl��[׵95��Ks�=tښ�.)�U���vS*־�@R��px�oeJds�����ʷȞ=�2ޭ#pU 3�}�v���l��|}t	�r:LP�������yz��W�7����*�n�E�k�ɋ�tP�.�Jd:ؽ�2��Ŝ�TEpܳJ��Sx��Yz^�S��n�i������z{�q�Ӵ�%�Uww��=��g�ܱ_b�š�[uo�#l�mocu�u����M� �b�_iܺP"�=���c(>��gY�Zqon�mV��BE�iYa��Ԯ����t$�ٗ��*Wq�.�r�G;PV)���4�M�\�.�Gڮ��j��.���SBy�`׏X�w�=J�84�����Y�i���Ԙ�ll�y}|K԰dk��c��5)��ښ:(�� !}��ߣ�9ҁ�l^u����[�t3[�r��n�-����N���4[��Z�1R�[���1ks�Mu�ދ��b����Wp!!�{\�/ݯ�Kx ���u��K+��܋�$¸�J�Әdd���j!Cf���:�f�	�Vv�q��A)����*sTR-�����O���]�� �ޒR����Ud�o{wO-�e�Gm临Rvu�JF�F�S3�
�Ŝ��qM��Hn��-V�X��vvw$�Q�x�~+0�N�o�h��%�4=�ǻ�F���<SӤ�L=lI45��<�K�����FsM�Y���S&�f���x�ß�Kv����L8:Y�u%`]�P'\\0J���2=B�]�Yv�u3w� S�NiH?<�ժ���E�f���9��mI�2�ad�!� ��;Σ�W�q����ČD4y�tyfa�Ms�̄k��
�j[,�2��4�M2+ȓ�j�Εt�}�9�m��S�u�w@h*��6Iu�Cq\�_vy�y��w�rc-�+�	y��H��ß�,�RYb�Y����d�(4b1���:����|˶#f��a�9�["g���������=�3�B{�V���Ag/#��eZ;�r�����E� ����h�̈���6�:E�t�\܎�K�ףϸ�>4����
~�|F�`��z���ۣbЏ]Ю��7��/�~k±�vl���Vb�q�2�N7�$�-�G_Y24�HM�\����v:�uS�	���i>�P��͗����q����[��Oo7Ͽ!�Y4��һ�"���ףr�g�$^�ջ��fiK��P�m�h���{=Ksr�6�j�p�3�oz��q�S2f(��n-6�qfm,��0T��2btN2T��C �n�Wh�B��!X��7[k�<H3�8�$NUYK34���WY��ʋOo\���S��<92P�	��o��A�8�4j^��lk��X)�[ڊ��<�f�ˊ�fh��;�)z�}����B)���V0���,ZGn�=�4ƕ�P�nsAwsY1��GC/�S\f~����P�6K�ٵ�z�usgN� ��%ա���]�*����I{m��.���m�F���3��p)٧���i���cF�#�p�GZ-.�T��B��P�L�V�y��SH]���ǈV��\�8���<��e�O{�oum-���EW�.��t��dc5�/i)@x��CY#:��v�3&T�26ұ2��jG��;쩲-�qrܤ�\�Q����Y~gD��n��s��<��fR�7��]\��TP>��oC�J�e�]k�
��V�TW��*��B������:=%Oc�C`�����v����g�S�z�K:��Hv�F�����b���WŴ, H��z�gQ�ʽ����KG�C{y�+^*t���ҝvޕ��1-���+4 �dS�y*�3!݆
;�{�Y�3gw$���9U��YE���a@e�Fnd�hH�T�0cxF���<W��`/�K>�2U���B렘1�\D��Ҽ����wh���v�ݣ|9gc�Q]�����;q`<�AL�(�i�䯵ӉT�h뼦��@j�U�C.�=��Oj�n��b��M���.u��=Xm�+�:}~Ǿ޵�/o{��7�l=�l��ma�xD+w�`c�'/PY۳z��AŃ��qҵ��x� ����o*ޕN�m7��.�c����V�5����(e�`nw�̸�[:OՍ��(�8���&n;�p�5�P���TI;�se��ʼ�:՜�@���(J���>A�9ٔ�P�i����nj|����*Z���׋^lB��F 3.��q���x��ҭ�y��S�R;��y���W.��9XW�)]����Sf��U-�sI֮W�����R۾�2B2��vI�i�ͼ��.��
�z�zDU�TYi8v�� c��J _Uw2�E��Ž+J�Jr�U\�;��R랝�př΄mh����S��y3'-������eܳՠ�iʭe��t�{vՊQ)��F|;q����\U�n2�%o��[c6Qn�5	AT�L�=zʫ�!ʒуn3a{�O��ڳ��'�Vk+%\���_c�t�ɇxY���]����EZ�_`;�VC����\�����8���R�S�g��=��J��玝(���q� 
x9�䤻�נ��6��Tof'S%��oZ����ȱ�i��oog^�Qpsj��n�K��v��0Gk[�Փ�~=���~FNp]�%� (^�Ha��8��.UdW��..A�c��RWQ�.����mo��,��0u����عcaȪ�vgh
1�ѵ��S��Vͅ�W�4"�Ls�r�bK��� �d�啶V��Fc�3D�e���ae��Ύ�%��]�#��B^��Ť��y�h�7RI�ߎ�8)���V�	G�k��g)��΢fݢ �e�i����j�Y��:y,&B��^S�t{j_�e��hzY�����U�7s��GG1�R0�věh.2�MK�{�uʢm�Q	�M%,ڍ�.30귅�1�w�qSw$@%�]D0r�^�����q�5a{u���Q+s��s/Rx��S�kq&�i(�f��I�x̦���!Rr��e�f��n�m�����T�u�t�^Al� ����ra�e�� ��M[��;RS7rVq��)m�/G8�$�[rڨ`��^�kz)Iy���w�V:�i�8w�e�.�L�����Y�!��ǩ�#b�χ'c����2񑴅�\����Y9�|�m3��"�Aӑ�g�;z7ήC�Qp�5}����kBm27�|�j�j�T5C�I���Dat��݊S��LǮe0x�<�H�3���T���m�7x�K��Vz��V/�KW��a
9ꗨ4(���۔mv7�6�l���ZK.�Wc�u��R�6p��ǹyĆ�"�zc/h>�E�-HJ�/Vj�%��g�S��?>��%��H��*]p��x������~����WV@�xB��Ʊ"+��]B����d���	W��G��+���"W.�/�^h�R1wVN��F�"nZ�nþ��C�kWIefw���5�j���\V-찫3����>Ux�'���&4P_����fǺ��]G�nH�=�9V�%e�6�s#K��i��&K���>��Z/�9�}9	q�$,�}�u{��L^�r�NyN�#Z;�Ov��U;���3���S[�9#'�m>�/cVX:�=�:��!�T�&ʽ�C�e��-�:ع��2��+R<jͤII&�m��m��I&�E��M��I��m��m��m�]&�m��H��m�KM��m�i��m$�m��I$Zi&�m��m��a��I6�m��m��m��I&�I4�i�m��m��m��m$�e��m��m��l��M��m��I$�m����Q%M��M��m��m��m��m��n�m$�m��m��m��m��m��m��m��D��E�I��F�I��l�=��;C|�)��02;.����I%��'�K�����V�>�s�|�aٳ��bü�$��5�|�2fť��N�g'�B�B��r	0RWkj��/g����{�FYA��(;<o)fL@�s�i�y��l�Vԝ��]ȣ�ٳx��^�
�hI�F�ݔSf�Y3n��EH�Zy"�6h�r?֮���3�ű��*jc��d$筽��:�_U���3����ǔ��~
��X�^1S�*u& �]����'6I���w��t�6�K�J�ǹ7ק$�A�׋���`^cn����nA����ؔ�>��G(i���iZia�eZ�7n~�tk,�l7��0��/��#y��>�u	�c�U9�mm�v��IT��"ŀ:��3i9��56z��*n�^.� mdʳ8�$��U��S�ƏU�Ų����R���3o���A��d��[o�;�("�bq��r���j�NMZd�`!��L�%��)&â�I6h0� �
�!���L�h"o2k(�.����.�,&�a�:r"Nw��w�,�cK�ol�|��.ŧ�&��Z��+TO�}Ƴ�1Vee�Y�`�����݊������ͬ
��y��%�7:�>��`V撸z[<�r�� �̼nﬞ�j���m���N�xѢ!�����<]p^��a��ЈݨΆ��e��5���-l��$���v�k�[1�r���@���r�{m���i��L��.#':��ܷ]k��S9���&�Δ�+�S��13��#0$=�B����$����=��x��K;QZ{j��a��v���ـM�k�J� :�����*�b�]�}��ړ �#�����'�B�B��ﲜ׳x1�p����̙N��0��]��(h�$m�ӷ.����Y�NֳY�]�Y֚a�Hu��]��Um�՗Dƕ�S�| �o,ᡧ.*�x.�ك5�s`Dɦn���QCZq��z/v�쮇-���]�6hT�]��܃1.�d&�Jw{��Y3J�Qr��3Sc�U�>����%�͓�����gu��8/Bǒ���l���-����d���w$z�Y������N�W�YVy�ӽJ�8�z�����B|;i���ppզB{'�E��ßI[�@fdSR!��+ Ø����2�F,\,���.�x8ws�7��lL����J�Ķڸ/C����C���bK�KJ��3-޳,y�fV���O0���w��SEe�q�u�/��n�7�T2K��8���<L��VZ��"�fOӕ^��#{̱�em�U�1ǚޕ]CeÔ��5�%�����e�C��A�≳��Uu�M89[���֙ǆ��I�c��$Y1��˺�H�����fk�]�����u{��)D����/K��;��Q�3�/�o�z#}F�*rh��6ov��:�2]l���P��!�I�3��NZ�Mj�V�I�f<Q��)�b�� quy�yR�A����^sw=�׵nm#�U�{%��dnPe�o�{�4��P�M����d�n��G8��� �y�w�EgIY�0,�@P�ǤUx���Sn#��3�z������s<�k�^��еJ���ή �#�'$��dL�ON��/��Vc�O��TV��,<4#�oV������+[W�
�nݻn��k���<�X9eb�1>�D^��J�+7����}�������&��	�jĽ�������X?��T7��W�X@Ǌ��{͝�u��-򶅾�v)��7�3�vİl]�y���j~�N�#+j�@��}�Z��:YOU��[U�z�B���m���(-R�������X��$[�t]��]n�胥b*�f�Ǘz�PƇ�2c�pNcB+Y�q�6�^I������w�>�eѐ3.Z�n�*���W��S̳��e�\J��o0b��Q�պȹ��we�%+����.�u�̫Ր�ݏ�A��}����S��W1V���/m�����2I1�sc:m���Ҋ�ÝL[��c uXe��/���uO�.�/p<i���~�Yw�)����&/�sGm��k"ڱN������"�[� yz��us���ؙ�����;`�x��LT�g�$KW�i�6��1S���9�r4����R�vΥ�J�����V(��7o^�{Ǒk������Ո��ʷ��/p���5=�U�)��r2p�����8��.Y�f��Y����NaW�h�à�����l�djIbY�aY�������|���U�W�H����9��I ��B$	'��I C�� O�I� I���@���@�!!��B� b@���Ւ�I&� ���a'P�-$%d	6�%@�d$4�LBI�$�yBN$��7`@���HuHn�B RBm !8���!��&�ICz���$�� B��I	�d!�RVH��l�� Q�LI!�!�Hk����d$Y'RE�z�&}@�	&2ćP1e��}���a�BK�	�m$���'���AՐ8�b�N$�I�!���,1��,	�@4�XI�
`La�� i�;`,!<�i ��Y5�$6�S��|��dRL�
ɱ�ƀa��`��x��0���I�J�RE�,ՁXy T$�B�xIԋ	��t��{,��	��y��B����G�as!X��a�̓P�hi����(�ζv�wH;�ݤ ��|ʆ!��$�Y��B�AI�{t'Y<�$�y���(c�:����²ޤ�!�;�1Bo�w�,�*Lx��i��3)��+$֬����pa�Y�^P�I�������>M�x@�	ܤϯ�&!��:�%Hq8��<�Rq�[��!���TuC�i��:�Ӛ�铩�Y�L�
��1/�b�� ��<�����ԗ�ڧwH��=�_o�Ѯ���:����m�Ӊ4��[
$�>c�x�&'<��g��L���c<���gS�}�ڟr�T�����	�4n��̥�8����8�G���5�]�}t�I��>���9����渚Cm�����t�ͥ�sw��:�SI�E=��m�t���n�oY6�c�)]g3��Z�_����[�Ms��b��L=f�r�t�s�d>C�M&�����Owa~�tv���9��}ۙk_}o7�Nj�T����� b�� �_�ە\Z��N&��wL�SS+,��jj_����0��<����Su}��`&K('����jfQo����)�j�Z��g{��׍[A�k��w(�B����Q$��I�d������1�%Y���;�*�Bu����o63�����(r�:�� ��ܗr�U,yM��P
��t�R3��6ct�C�f�-t��*�v�(=�w0��As���#����:Nt��7i�����#W0�
��(at�ד*q�*��e��,:�P� _����R��t�eѽ�U�����x���lJ��N���҂Œ��/)��������]`cz27[�Q�*ģi�2ܮ�g�*��P�"ڶ�E����v��&�߹[�:�Õ N�_�X��$�q5"V[L�劺�P�+2 B۸���� �3J���X�9(}+(�TsùR�:�m���bH��sL?�8� A[ʣΈn�n��n�1CF�^�v0즣�ko2��Ա|�D����Q.]�M���!w�{OYR'p�b� ,q�Ff
L�x��9�v�����b�R ��r<�l9Ύ��~�鳱6��ͷ��C`^e�#(��y�ī���f[�:"ѣi�xq�U��
�N\�<a�wb6Ne�VAE:ɖ֫�^$:bd�1���?��n���e��
��Ҽ.�Y*@�~�vFY�Mu��pͱHu��;U �!+��#}w�m��SA� h(�|�:��d[��u%8h���q@k���U�у[��K�Iʘ6�d�z4�t%Ҝ�a���q`:�~j�$�
.�F���Ҷ�t��z�x���.�L�R��--���4,_2�R�fܮu���T�F��{]�Xk�W^ �3`hבV��-�ۚ)*�d��z5H~X4!��%ut�W2�:�ͼ�5�8���r1�m��v����-���o���*��YN�Y�q��9g;��E�s7��Q��(�E�rB*�Ҷ͚Õ�hMb�ubQF�ˬ�)�0��#���\{.Z�F.YC��S�М��
˔�Y��&k���ʕj��u�/���
';^�8�-Ef>�0-L��d�k%�����'�2�	;���қG�w@-��۬�� �I�5+�,��ѓ����=YYQʲFY),6�����pb��c&������WIAm��wr��=}����(L� �Ե��ąn����SȞP��/�v֎�n��i�X�{���a�9kN�����cF;<d����1�;T%~@0j��ܣ6,:҅67Qc����71��J��*an�e�-9q��-�Ǳ
;�2�L����@V��A����q��S
�k��{��Zcb�8%�܌-�z�G����pʘ���,*%d`S4aq�Ƹ
��oF=ٔ�ݲ�P��֕׮sM�DPr�c��f����5���$��2�:%��n�AЩT��������ʿh	�88nB7���1���τRd`��<!a`����|��HUi��#H��Xb�R�)k"�q�����.�_�'SCP�t��? ��$Չu�Z�ʔ)j��b��k!�;#xւ��D��T7�Q��ݳm��@R�hl�-=9��^�uWt4M�dTu����Z�qٜ�u���Z��-�&��ѥ.�*(�&�T��RJ�Ef�`� �ѧ�٦)R6�a j	��.��w7,�i-�vJ5�f�g딙u�=Q��]����L�&�H��t�4��pvkDV1Q����ŀ�XV�T��CVG4-
�iU('Ð�V�n�К\���e΄�ӓ̦��7U�&�E%)86�KTZeg?�T�;\�!�Z�"�͑�e��LV���Ѽ:�@�v���["l�
m� ��*��*�4���*V��ۈ� ֕�N.q�i���ø]:����4��-"�fV�;���7�.�x���D%i����gM�&�V!��?Z%#n�f�Gx�(�X�q�Jn�^(J5J�d1��Y �Z"�\:�pK������5�:��Z��lcQ�1�[�8RY�sZ�)�Mt�`�ЇC����׵�Fd{u4�BQْζ��4m�{c`��w]��9�! �$���?�;�������泿�5˼��h�8ƫ��Mm���NIq��B�)c���8�jY�����f�B�Գ]aG:�n�����'.'�ɗ[�8�����S&�E{�P��j���>�O��K���F�\�ݾ�-�-����X�%��Mڊ������}�{E��׵z�d�A����<�#nd��,n�׍�_s��q @g.��+uF�<�*���9&�h��ݐY9vb�x�A15�)��Rl햺٤A��*ƭD���'^�v�XA�<��ry%Oz�쁪6c����y`Iv!��c������f��_=]�"�vc�*�<f�>��͏���Mt�q�c�fQ�w.�Yf���<Cy/������P��/�ӽ�k=��W� �K��z��ʮ�o.�S��[jĭ?�K-t�/{yf
=}j�s�a�]��,^\m��-&�I��I�[i$�I��m��I��m��m��m��m��I$�'�p�@U�we+ҲVQv�"]�{X��n6�E-���B��`���"�D�A�I�����G�<F��kX��̳Y�Q t"�ޛ7	��`��]�?�wn�x�P��	K^�;q<���.�N`��p��������Ze}�œ�����ۯnz�3��>O�LX!�fV<�M�.�����X�1�(;�P7icQ;�̌3��-�A�y�*�ķ��*F�$=A�gU�{�n��fs��ڿe�g>�5�Ԅ�	�g����ʊ�ڄ����I��k@�Y�?e���iE���Gruս�r!!xZM��Y����qt���£}�#�q�"���y�n���=���s_{���k�a��H��	Y'�oaa m�ClO�Ą��-��@�2O�!%݁*`�@�d�P�^�! VI1��P��!�I4�!�Hy�i 1���!�@>�wP���u$a�I��n��bB=߷�ڹ���g�s��{��E�X���
(,B��R���DAEPYQQU�1X��
,�(�$UEP`���Dm*1Q�Y�h�X��"E5�TEDq(�֬Qb"��b(��"
�f�����EE"#E���#�1Z�X*���P}j
*��DUAVc(�ł�A�'԰V
�1QGHVD_6)���EUE�U�"���T9J**((*�(��X���QDUEUEPD�E}J,TV(��b�X:ј�"�b�,EF���h�QTQbF+
1V�b�"�"��TTT��ŋZ�M%b(��V*(��,U�*�EUQ2�\�TQ���(�� �Db�����V
1���Ub�H�B�5����

1S�QJ)�Tf�AXȈ�b ŃT*1b��j����LJ��A�**��\ϵ�ERn�Wt늪*��j1��E"� �e���b�X����g0Ɉ�b���D`�S��U�`��AQX�"����* �~<!��׶ˠ1ZLӳ�u�3ݙ����%U"**(����S��TTDX�2�EL��w�}w�QQ\J�UA�?Z�A��"��P��������?e��AU6���V9����Tb�>�g?���h���X�FKB��E������U��*��b�1E2Ԋ��FDV#bֱb*�ߵ�EEeh��FE��cAQ&�~j���l��*�R�P�*
��#D����1V"�Z��DE3YTQ�U&n���Tb�EW���h��F1[j*�Ga��b��E*�(�ETU�"�x�~��Z��"�51��f�뇯.ءv
"����8��U�����LG0� �""�_�{X1TDb�F	U�,dFҊ�"���jdH��-�h���QE.[QEG�T]}�����|�0L�b���{	�X�ަ*�эh1f��]=�(��`�����""*E�~�� �?kZ��.����#aib:j�T�Q_�1Tc�TH��WmF*
E+�|�"��k%TiT�i Q�j��ׇ.��?~���5�|�mO�AFj�1�)�X�)T0˂��TDQ�(�X�,A�7b>�p�T�v���,c�8`��MZ:�F#5��5�D`���z6��X�1g�U�Dk�kD`�R�V(��f^���DF?4^Z���U�R�3�1b�}�b�XV(�A�����
n�DU6�?�t��i��)]}�(�ՕCIH��-��r���������=�}�9��f~UY���<�b"�����6#�^^3"�t��J����S
c,�*����=r
}l�ul`�	neX�")�'�)�Qe8���V��W�(����)b/0�}�
,wlE*�_�v�׾����� �"9i�w��[����b�+�ܲ����⮿\�YV>���� �E]^��g�{nw^�][���� ���j��DW��IE���&+��(�),�>�mګ[�+�����j�:�Ub����k�TձT��LE4ߩF9h�w����N*Qb+�Q{�ښ9T�(e-�(�,��ɵ�3*��)2}����5k�*.�T�
�9����k��s���r�hEQ�c����j��^�X���PL��R**�;�}��!榚�j��W�kB"��f��",ˬ���]�Ԩ����~���.�ŉ�?SC��Yo�EA���7�:�����E"&[���;��;j�������b���pb�����������˭-�N�[��ǰgfF]��?"� #�+�\��r�2�k�(���v��EX
��־�5�\��5Z5b��2W�^���I��fTUEw��]GiEDjX�!g�dES�Չ��dG,��T�X����P?fx��hP�X�_�������Y>9��f��������^��颱���?w\b�w��fD�ߴQ:�?'=�w��e���(����b�j��ݹ�<q�j�yKw�y�]������M>d�6�6��]��4,K@��)�޻����)C���/�A2v<�\�ᾬ���-�� �e�w�Uͺ��H�L���ׯ���s;��7�g� ����vZ���3�W��|=��Ú�$�Fb]��ۏ����)Ɔ��oL&�����{W	6R���ƈ�D�x��s�<>���)�I���,t�U~�\�C=���ATUWٛ��PEM8�0DUZ��`�ְ�/�*�����a�M&�A2�-*E����o�AW|���QkQE�[w�4(������4Չv��49lTE�癬(��� �m�Fi
�9o?S&��Y��
��^|f�\��~�w�iu������O���ݰے���sـ�"Ńn�MR������6�?�(���9eO��(����7����<�M�3�̦�gɦ#2�?YTO��Ub18ʓr��S�QT�b1E��F�ӚO���A�5��_� T4EW-U���~	��?��5��˽���Y?<���;��O�8��ɴӦ��bJ���I�U��YQ;�~����X��X(S߮��Ub&ڪ��S-o﷽�/iQ媠��ʁOYL����P�2��6�	�ʔW,��S�P}��*����#�9}��` +�ҡA�T� UZ���u��7,�?s��|~A�z��J,�ـ��X�C�@���=����U{j����,��Ʀ3��,V �2�§��٦M�t�!����mQs3"��+������ޅN��!EEFs���6�h�4�Z���t¯n�#Z?Z ܹ5DUA)�{�I���"���[�הQ�� �*nʊ9q1��}��)�TԬ�������Y컴S��_�I���9o�UGW�����h
�Z<�O�'�ܼg�9J(=����|�ݨ��(�>��6)?R�6�]j�?kzUf�T�~a
��i?�����V2�+���X�=d��Sݦ��w&ȋ�]ߞ3[j���ɠJ���Qg~�i9�*���'������WI�[z�5��T���N��k�v�B�5̹Tի����*+Y��~�����(
��u?&P�|� B������ :��b�����u�_����T\�Y3TU���ӈ=L���*�������7��8��4W?s�6n�Q�ea���}����b���s���7w��*+���S�8��p�E<���[b�*M�.���rK�(�Q�q�}��t�7��
��Y��3��4hy?8�J�S�U~�n�*`ΥL�`������V/-fS/NS{3f�>ʈ�?n�cD5L �����;ڇ�x�!os�t����y*�����A���Pݨ�K�Sg���N� ��/��?v5]�Z���agc�L�f45j���"��%U�Mڗ����S��1F����ʯ�*;�Ld�M|��4�2���X)�
T+�*&~�����QY�_}�����Ъ�q_z���l���>k�[� ]Y����t�痖*��tt0/_�C�+��5D����ͳi��hP� W��D���J㉅Aȩ����1��VLF5�>�qշ{ɥun3��'uN:�+���^'�R��� ��(L����G�H���r�r�λ�k��a�����О/Ohĥ��<��m����:�tg>%q���^�G�yp����F�:F�&ea%�Ƃt�نO�+]u��ZP��El��t�� ��i����α�%�e^�`]����\,�T[@��ˡ�>��[�e1�
�[���~�����}��Lo�#��R_�d֚�K5M:t)ST�Xv�U�����E+*�8��Z��(��b�ߴi�⩬�*|�2���h1_��kX��ID���f6�ޱ?79ru�E���y�6�iޠ��
�G��(�j�َR�����^]8����@?=�` ��*ʀ^�M?2��3-N��y�U��e-/�޵Zu(3�5�J�ZɍU5f�L��!��f�`w���>���{x���*8���%5� V��	�}1ns4�����G�δQ��Ƴ�ٙ��張r�Oɇ�g6'.sF*�����hr��m5�1����?RԸ��g�~���bm����X#�+<��H�Q�J��T��4�1p��| �I�[Rߎ�}���Pӆv�XcT�r���F����l~x �����}e}J�9�E�AX���rh`��0��t߳��7��S/�k��[Dj��$^v�[^�����u���Q�	�f��"/�����ut�շy��;T�?&�uK��sY��~y�E �_����!
b�5N��PW��e���N�z��L�ߞ;��h�[=u�=��>�:H'WRHU3�8~ /v:p�{\�_d7��ƴR��G-q��1K���Hd"���5�
�(����o��_�sۮ���b=�7��/��]�	�T)/* �o��󼽞7��TK�7����Wu���T��J�?��t�e��տ���N�r�֯�fw�\�4{�p����L�}�ӥOٽhr���jUT^n�s�{� h
��F��`:�V����ް�����r�4P5߼?xV�Ğw?]"G�e�`3�fZ"�9;�og��*�v��h6&��K�\�L7k1+?|�Pf��ⳬ�����F��J˥ͺC]����b5���q�˰��'V���}����+�al�s�Y�M�h��؛s%L���l4�������YX���M	�1d1�9�?~��(��|� �b�*���@i���v���T�I��cޕ1$��d(�>�|P� u.��o0M��Gɡ_av�ݪ�p��$���P��b���2~5������Uo���`�Ͻ�&}܇��>d�f~C����L-�D��`�p6ϲxi�fۧ|Bv�Ԉ��ǜ-���^�裓~ys�q�ʺ�u@��//�z?yV�N���yu;������8l�W��v� �ݜ�bl`�mvn��ؓ�t	��i��Q�r���Ũ)˳�o�An�4�ܖ]���U�����RC�V
B��A7}ރ�qyfaU�kX�(������ G޽Y�x� V��W�̨@�m14w��zvlV�Y��/�����������T��(2�3�
��c��b�q��o^M�J6�^%�~����A��{=����.^7*�+��J�0s,
�Z_���"��T�F�{�g4Y��*S;q�M�
������*{=i�p+���}$"�z�j��P�-yit5HP�p� A����KGy���HHy���V��%�M�Z�"�n�"w�S5F����x!�l���E$vO���d�Wun���Ձ���*b��q�P�F����:43�u���Ư�1�]
�����6df��}+�3�AY���H�T�B\��azR}��S��m��!r��3��9�AX�l�)�q\S�A=�@�o�HH&#H�ƭc�����Ƒ�B��2����7����_��:�yj����9���� "�p��4E����7��U��yn�~ě�ZY��w3�&�ֆ��4�Ȑ ]s����r�p�b:���ҧ�d�� C����NP�U����m�Ҥ�R�����| `P�n0��w;4 Þ�f,�G��ՓCh�t)$���EדGJ�����u珵�KxoX���^%h�e*(J܊��'�,��N�B����n�cU@�*�����"l���e������|RB�&���a TPݿ~�\�u\�O�����\J�ҩ����@
 ��#^��.�TIPy�A����iЀƪ��<�Qr������z���tK���4�#�<���lm�����^Į�R&�D׻�H�~�2Wdq��|��� 
�&�zA��~� "B^�-$,���on0��ߪ{���\�u�ݑ3����F�e��0¹�c�=�Nc[�~6߳!�_�kv�[ך��J����䒠?v��!`�D�(�4j�ay�~)���P�yvy�}�w}�zĝ;55L'�kkz���~_��K4!}x_\�=�i�N�o�8�6��[�Cus����2�2\��%�-N���t��}���v�q5��mZw��,F�Qbtp�7&4���m��o8���Zsx��:�z��sWiU͐9�z��IY�����{R��FѨ�x*rט�5�ݲ��M[����F�������a0a(�H"U�J��a�����(��䬟ޙv��Pػ����V�ߘ����wt����F�:=e�HK��	V
�K=�3�I%J�4a�,0� L�c�G
��U�=R���C�.[r0A��9�����ǘ��;�ۃ?:���,Ӭ��bc~�\a���ܢ��4O�t�g�GsUAֈT��-�4k&w�=�SրP� �7�B�,~b���yhf��o�K�]���?u�C��K���uB�T�@�
s-��a��P�֛[grUG��������懟�%�Y4�JB�4GR�	g6�㸈������ ��F#Ua�
����K@k�cO���ߕ4A?��F�h�̦q�_����\Q�j!+XE�_�4�GH�Ǒg�k/@��p�%E1r�!3��m�#,%(������|���Ð
�J�g�S��Y2s��ت�� ��zꚡT(�����N��yz��Ԩ�� ~�]���߮�2yv���4�/6��ܪ$
��~8�VK��x��}�J�H�z#�uuO����4�F�|��Cߺç����؉�*�Q��E�;ʟB��L��+/9��h�C뉢A����U#����Yݝ��@�ڞ������	��k�)y~(�d���H1[AGX߼U]�b��v�I�����߽Yݬ�g��^�$+�ϒI$Mx���^��oF����KƁa~[����ʩ +��_���:kh��}v6U
�b�V	PK�����ve{���~B��E=��֕�a�A]�����w
���L0�'X@����c��1N�:|���&B4@'�ؠ+s3�Pz�WSI
�S|$�O������iW�A�\��̄�ߠ��$���@�w3{�BC�$��0!;��I�������	[	�x� ���Hw(c ��u�		�oz'�� ~�	|�@�'�XO�B>���HI��$1�il�wJM��a@�C� �	 �	̐'����~�����9{Ϻ�\#�V�9 -r͂�E�~���p�ԯ����������R�L�8e�V�f�/X7}�f�y����Se��� �J��(Z�w�!���#G�9����kVd�
w��m��׃�ՁXJ�(.�ZZ�I�7j��m��z�ď��P��J�u�� ٥C��0A�^5�6��+�'qy��6�dD*�D7Ͳ���
�@}�t�����/��k��J{��EQ��g�ӫκ�ۼ����m2|c�sY�k�f}�x1EgT'7t<*�x~�#X�Fz'�<#��L1k]~/�Ԙ�LM\���1��V���uu�X����/�+�����2@�{MR|U��u+�g�%\�<|�Y�o*�{W�Ȇ�b���S��!����i��=������{�5^��yV�;������pױ*Y����d?�L��ʱi�/3`,v���C��+�w뼠I4�6�Rd��fｯ��{3X������W5�2�|�� W�c��>Kʖ�W�W��5H���fw�25m��Y�DρB��H��w[6�W.���
ݕ�4/�o�i,�ZT���W����U(P�C�v��<���s#/̮��-�DT �3)u6��(��}�s�����(�3�m�wV��>�7}R���V�!w��q�0e�B�c`X�Wiק�{�(P3��/�{-{�@?�T� i�^WO�<����}՛Ť_�R���;��6]ng=O=G�Ɋ�,�W�t������LY�wugsگ�G��^/\�@P��Q4G���]{�M��v��4��O�e�W0�H���0��.$ ��uo��#�0��BGa�Y�Kʺ	�T��\�
����knh�?�}�}��O^{����s�c$���������w�����z���������~�����Q7�%x���v��4��d��m-����Q��F���U���7�������{u��[V�Φ��lSk��F���Y�å����@��	(q �Q��FrK���c���̱;Qc�},�����pyT�H�T뼕9~�t+K}g�+���N��Hyy���
ШVx�k���K��qz�����()�R��D��d����6
���?-p�^I`T<j�3��~��fxQ-ѷ�K��v�����x~ Rm�LQŷ*I�A���*J���~K��=���4�P�Wj�w�A�^���3FP�
�hx�K�ś��D�a
�ҽ㟉��*������-�H�u��>
�_9�<<*�X?��"�-L���V?l�/��be!�U�� ��;W���r��T:�K�)+���Y4I��&+�~
�蠰�1P2�O���E���:��e�L{�.�
tEx�0|�Ԇ��2 $:�E�0>�{���;�W�J��a�
(DI�j���zҼo�{���Q��
�������zL�?f�A�Ǧ\����8�S�*��]��.���	^=U��Xkޛ|U�>�ZcگR<*2�y"�b�i/�2�&L�[Q�yf���0|GuEBYP/qYb�8���{5^��n�1޹v%�W.��0�{�o��X�Dlq��|�P��ǲ�>��t(U�E��L{"8;5D׏����uw	A��Sv?�Kʿ@�e �
�HF�T�[�Ā��>5m�E��K���EZ�/�����'	B�wo�#�-5.�mذd��܍�Y��b\�x,q��)k{�t��V�dny�7h�=h2�A�f{����7���*#;o�dZ�������ʝ��^$ߘw4e�麂G���%e+�����	��3:�(38�Cl��l�z�*?���I��B>W��kVX��	ׇ��[XZ>��B�p�
5Z�P���:������%r�H����}[�M�Z.�[���X��$u�t(�w��,@9�c	���Q6��1��3��~H:)��
9���1) =Y����W��+ҧ�d/'���z�xT�Z�aݻ�ᵐaU��yW��:֏�h��ՙo]�<�^�Wv�n���"��BeKZ7�0�x�K��άU��t���L
�F��U��
o*��-��a4�t�*���bs��&�i�֏7��\�ˁ�Z�q��UF�����#�쟁�]?{��Ŀo�TjN�j%��y�c�K¤?�ghK
o!�R�G ����AR����R�T#M�)��B]�b,DP���3�����]�{o6�%]�&�/�z�&��T�޻a]�v�Z���mӼL�"��Ԁ�O �*uHח8��EM�sѮݴ�v@�����.���|Ə]X�Xy���)W�U,�O�u�h�D��þ"xTGh��dw��Hn���aÝ{%dG�+1��C*��Er3v⃍p-֙y3O��R�d��y���+k�I4�N�o�.�%���q5�u���W���{�q1>�~{�fN���_Fv�U�iWQP����A$�W���U���v�>�ձ1�C�D#]������]t��zu�����65�m��0.R��޼6�����Y��_oWʓ���X6/Ն+I>;x8S����� ���s���'mf�<�.��v7[�D�5qD�d���)iQ��j��ͰO=���'����r���ճ3V/�q�V{���a�+I$j��7��ؽ�.\) <0pU8���ָ��z!�觲���ۙ���3�Q����Ag��ݽaq�Gzg�u�u�����ݧ����Ugnj�e^���Z��T�n�6��L��Gʪ���+�ɋ��i]/�;�p��ԼZ�8,,�߻��u�g���B�`�+홍�Gon�o#O���>�TU�+�1ʲ@�O���m�`0}f��*�Pg������.�A.C)��o�+�|jm�8���,�����p�OaT'Q���7V�T�xR��#�M�ͮiz� �Kౙ���}j��Ԙ� z�4u���,�~�f���M��[��J�!�Պ�k�J�k�~�+�1ި0<8���]��trb����G��Jڎ�Kפ���B?A��N���^ \c����G�]�s����ei�$Q�IEp�"�|�;9U��#��@�JW=^u®��M���U<��-�]-VjM�o0ա�^Y���q��^�ī�^�}��tX���^T�,��`����i�S��L+;�ܻfS�%;������(��0s�U��]���<������z��N��<������vg+ӓ����Q�aT�&�2A��������9��nR�*Gz���-��U81�ڇ6�7��]_]�ǐ��q��]�6V؍[�[w��+�[�n�mg&�u�l�\�s��ɩ�ћL�;X�X����i���!��r�]��������f̋�ItY�+���eK�s�x}�b�k�Tb��J=$�Kz�ܬ]gNѴ.�^M{7��b[R�Ɇm�S~��҉��9?pUd�V�!a�g��~
�EΟ�;������Q�EeĚ������_	U����n����w&�,vt��m�竒����޾�?v�C�XkƇ�a)�r�qSJ�)��zǦ�FWƗDvL���N"���?W`��|���
+������/\�Y�Ow��J�� �T�B�C�e1�!N�h9��cs`�9Y�G:�xh��J+�����~��q)��7�g���PƁ��R���~�9n�*��5��u�8��9���9C�;���܉����F׌{=���!pDq4�r�����3_l���#����C�/=j�w�*�⮸�v���>��˗^���M�'=�u^��!Ӭ�^�.�g�fpr�U��3U#�`X��=
?��s���M.�?W�g7OU�x���+��ux��6����Ǟ�,�9t�6�p�9}�|^U� �����x%?H�b�3��Z�fڪwUq�A��-cU,_f���2׌s�����p%�,GnU�W��Y�2O*����9�o�'�N�Gp楃���{��P�*��9n�Wfn{�$���,e��ljT�P��C���o�sS8��N�n��w�΀��h�ns�i
����CoU�^r���>�?r���L�:'^~nl1���_y����w�Yx{�T��\._oc��j�0[���vx���Hn�O/�~��oj{��3�<�{\̺�s�{�+�<�$�Al�+L�\Ѵ�(���5�X����s+���9�i� ���V�CB�6S>��Q����U��|���� j "|�4Ml�K�E}��ݧ^���fյ�����P��鵞^�7[�vY�9k��gM�*ޛ�l־�x�u����K�q���������W���K���#��:��t`JR{��3w��jԼn���"A�J�o}w�8��{'�Et=�/]�ۅ~Y�Th���[��V1֭�����u�{3wc���L��R���~~��}+�e�3w�o�s�+̷O��_�jꀒ���╋�=Jj�[y+iaͰ1.b�>�yaqX�;H�{ڴ{x������Z���F!������Yf_�����rn��T9R�]]�cU���)݈`�	���ƍ�d�u��|�K��;�h����r�L%.�y����j�7�����O��!��U9�J��H~��4,�a����ш^C�뷺cz��"W5�%cs�ԐZhm!c��ͮ�)��u�$j��鍾�锵���҅�n��8�]�"�Ȗ����/]铓���pc?�."�"<��/�7#nՇt�gRy{����]XT�{֝���i���8m�2�ճot0��d���������N���"�ܮ�<{��l�漚�����%e$��͸S��mq�W�_,�裕ӍZ���_���ɱ�\V1��N����22rR�I;�ɜj!]��ӴxA6`S:��P󗶷jt+�}�4o�yU[��ď�Cj�x�K��Ǩ�jD��+n,�a�Ɔ-]��ˮ���7\�@�.,Z�ڮF�x^$]�w�8��0�V��ѯ��Ĥ�G%X�	7���wv����o�Cr��B'S�{���z��CN�C]4(����fX��Ò���v���6��E�Z�0�N,�M����rbDul�+r fM�9J1�Nf����J�΅ҟ$bks?S�۔�mY[�Ŵ>����=§�<�E�7����U���)r���c��E�Q%�.��)9n�ͱ��#��:�i^����U(��U���[��c7L�m�쾥�!���W�	uo�N��<�Nm���fӳ�[+y6��z\�W�<Xǂ��%ٍ_���W9�R`#�`g=�l�e#����է��`i'>��w�i}d����hx®Rw,>�bLLO�}���֝0R?�
;J�O�ŊO����tu&�J�+���	#�aE��F�or�4�wevnZ�L�����䏨�޽��f��$ӂ�|a��*(��NO��iP�PS��k����&Ę󅆹eEL���7��?!������oFՆ�t��~���u
3��x��Q�t�W¿X�������.�r��{34�{�DP��  �A����'7�%a����_�����΢�r�X���1������QT��b�j!�j����������k?`i���>�OR��SHbO�q6�����a�!F�?\�x<4��� #�?!D�g�4�+3S?�i�;M��aDY���	P�:q~��f���6~шk�O�i&��?l�3�#�Q���=IX%�I���Ϭ�"A�k3y�L���)<=���]n��2��ޮ3�+W�1B#E��>��U���M�Ϳe?&����^f�u5�!SiJkZ8�O�*/����Xw
��9�UQAAz�{�z>��|m�:~������`�e����hG���^̞�W}�o�\~��i�I�I�;���h��-b�5s��o��R)ĩ�v�1�s)3>��j��16ʕ?kXk�t�U��Z�,_�()���1���� ��~�[���<�s��ϋ�&f�-b����R�J�Q_��2��f��}V�2�l�
�� X���CՁ�ǞV���m�SJ��{�^��T͜��B%��\��x��0�70��H���Bc���������|8�y�&�ܞ��oޞ�����2%I#3�Q� e��#���q=�����^>T�N̙�{�%�,Ƭf�����Eg@���6$gw�p�S{[3���}fcf�B,1�*l�FF�"��*��0Dp�V^��3�&�߂��V{�n�oV�����Z����mt�g6��&nݦp��8�S����,��]5VxE<X+��0�Tf{��W�P�:C�ǟ:N�]�y[����:��؝õ��k�ڬ��螮�0Ib��QCC�(1��e}�_{>������/MM��6\�DtD�>E���\ϧ�遘�mD��ν�m��T���%�'X(��}���{Z���BȠ�k���Vء+ݸ3�MVzU�~�ΕF+�c��܈!R�X+#_�1�j�h�x�~A�:ݩ���qLu��^��6s�^���]�.g����ү#[�(�X�/*h�=�L���������,b?�Wƃ���)��x*������}@�g#�wҪ����>0.숟����p�_���TO�����\
��8�*
�n_*�b�wd�9]����\ ����(qH�����+ꁻ�NM\"+�d�砘��v���Ǡ�2�c��������VZ}(|b�c� ���ӝY�B^��嶶�K#)�J���#8d����k���^T@���T�������qb���"m�F�4zI�O�r(q��Y�Ū���ǣiLVE�����XF��|�e��18J�w�<��P�?!K���:�}>1D�U~�Kw�_�c�~�y��xz�dc\ �nv���~��u֌ك�Cj��2�Rb����ԳG��\(�|�챚_�⻆>/l�k
�")Qd{�S��<�F�^�s^����x��`e��S3*7֞��c��b������zJ���w�d|�I�G7pf�w�M&xA�,�,��ub+���3����SG�m��#�{6�K��������|�D�C�לi�WLzWsU��Wu�����J?f�a����-u
���U|�/d_6í�oM�T����_=�8�����陜bו����{��N�;������걑�*�c`U'%#�\����Vg�UL����w����-���Ԧ`"4�S�����Y�:�~^x:���G�G���]P�բ��Э�~��nnf�ȫ����T8�P"�cD���L��h��PޠmJ�5`Eso>,�W�ȿ��-Ԍ~��D׳�7�6ↁ�;���O��l|Œ
q��ь��
4��5��8����j���ꡧ3�3�ݡ�5�'W�x��sp.c.�?B~����m:&o��m~��g�U|�UP<5xj�9�
��1��ǀ�#�oa+�˻�݉��.2"����1x-q�_+#fѩ&�3�劜�b�љ�M�h:6� ������2��׸���|7�Xfx�^�
V�M��˶g�+��X��E�j`B2�2>����������Eb�>����+c�0��������tnP�L�JF"�g���]���X��Ȇ=�1 �N}��V�"C���#�;PO��<~��O�/�/U]؏X�<���u��}M����N�:���m/=-i��޻��0ݺ#u��1��7�Y7B7p�tW��1�ޱ9�<{�"��)����5\"Z�Upk�۠q�d�u��Z�r���jqpB�bM:����oч���\�ڂ�����ӂt�C��#UN��-e����f�ȸ�wa_*�Z����@���*'N#��U}6a��QC`
<!���B�gh�c`߭+��y��������κ����҃b,c�Wx�X���NR�3��D	�����& C{�&�i�*�!�7��Y���ؽ�m� �e�X�:cDf�b=��H@�A�ϰN��,��\
�ǈ�q1Kظ��82W�n����yy�|X�uZ��9�u�]z�,T����5w��ʬx�눱0,��d�h7�͋ߌ[���ūk�Y�K*������'y�d|*�~Z���=�Dp���ɬ},h{&zy�"�w�xM��}��W���<����b<� ���f�#8,��3��$C���ߗZf5�w#�H���3a�>Ff�^�߲?k1z�v�k�T3?|��"�L��������clƂuQ��-o�VQ9�Sڼ�I��q�O�f���Ypf����^�uz,��3�)��R)���A�Ȩ�Uc~�����_�K$,�wt����4�W[�-C��}�;QuV&���3ޏ���g�Ҹb���ִ��z��εl�}�Z">�ڍ�jh���׏�͋���D��(D|���U����[�z�{=�h��/��O���qQ�{��\=���LU��#[*��{�5ywu0s���W���Oh�!�t��o�N����ݐ�덳S Q`!��4T�̸���ʷ6�6��� �V�^�遀�u�;P*g��^{`����Y�6���f��$t��B��۾�Y��<��c�VR�����b����^�BL� 45���Γ��`�6ֆ��S�{�?�ǢQ�h��!��o�5?W��&-G��^���N���cU��H~"���ʎ	!Qe���0���P���M���9��j��Ͻ��q}5����Mu����wȐ5�&��yO�=v߶����H� �AC��Z0u㥦2A��Z�����M�3u�V��Y��C瘢�f�0G��!��鋣�d�]�Y#Y��E�O}�2�k���H���qi��7�o���+���ͮ�h��G�Fuͥ.��E�܏���o��t�gG���u��0E��wO�j�M�q�Lb<��N��>�����k�]�6�p5�()�gc���o�=�c�F��zWv��2��^S�M�@��O4A�b�!��jDt��/�7��ؖ=��;�v~܊]`�?h���@�ϰ&���̧bp�P��� j
��ru~����^��+��g�g�
��/Tտc�.�x����g�O�ï��=�.����<J��lyfI� �gk��c j��lt���V{]=K#�C��[	:w7-��ݳ`+3(~�m��Zggj�b��y[�DǖK��c�A+�fD�X�9�,��;f����C-�N�jZ����2����ܻvu�o�M��^z�@K�)��4noʦ�I�*�*���|"ZE�
q�l�ʩ1"=)�K7#j������L1�t�� ��;ɝwٚ��Kl�u�Wiֳ8;^���/ˤ����D���J�9�ص��л��K���_=����J�BZ)I�j���B��H��EYB$C�5�i��G�h8�n'�{��=��b�������$x=]@h��u��FF޼U�M������*e�G{���K�m���Ν�g�0�;.��|�q6��|��&�E��ס���mu���7��"���:e��w���rI�2��Nψ���!���0>BI!�@������gR3Ix����b?N/��>��7v�"4�:����^�#�z|��U���v�c���W�ɂ 8|9����c���X���s{Ц�&�r�ϔ�X�K��E	w���{��m��@Fu�9��4SYPݭĴ �^խ�ʯ�a�6彖yT`�<<ݏ\���f,.���+��(\��K!F�{jc��ڧ1�ʽ�ʞ�6�P}Y���Q~�߫�֓�x��Y�U~Е"�Um��W�<�UΝ7���w�k�.�28~hC��I�d�^�c>��:�J�������Ӂy��q2)���V�^���|f��⸉���z�����Yi��0�9�u����՞i�C��G� �ӹ�/U�i�v&;wj�ı��{���O��U���ywNfc�Ѕ&��<#���Y$�d�A����?O_x�Լ)]5��T���(��ehx8P�>������P������ovE��6>#$��Ѓ`�X���#�/�y9&��#1�����/^E�f2��u-9��Y���.�P�w�n����oO�����1�
x.Sw���rg�߮�����:�J8#"�Lm�HWǫ���>}｟�į� �e7el�hUM蟼D������x��`����h�1�slO�L)�gN!8UzcX)���k���-G��l�Ƭ�
����͋�3�Ȫ�Y��T��\m94���#��>x�k�������q�#��J|�]7�`�Q�i�W��)Izɗ��N��_{��.�Vb���C�gtp1U�@���l韝���22n^ӌ�W���5����n�%�P�
8>��o�F�f���mX�E�ו�1rt*S 	҉��G`}�5�|o�Wu�(ui�����u�#]m�ٿ/,�������������~�Ӻ�BCj��<�P�uC�״sy�J�qN�p�Jr�A/y%ꮡK����h�Q�v�����+��`�Ƿ�?���r^c��F����{7�\`,��S��Y�F�
4r/��N�/���h�ʤ�3��GmK]��`� ��t\�9�-ˋ66E�د9GB��)��+6�3��t�]�HP^��8�|;���,�/l[>�x�yux��x�;:�FW����z���yv��������n�y���1�K|��s껠�U��\3AF�2=0%���}����N�۩߼2�ې�P�Z=x�����o!�MMFR4w�u
�G˩���e���֋��oK�N.3��^=aB����_w(S!ěȸz���7w=� o�z�eM��kÌ9�v��S����#1��xfx�_���c�#dTC:==lt��e_C�)}��>~���\����c����·�����w&����*
m������O3>5�ʽX��s��u��s��x�N�����zT�K�w}�鶵ػ�d���:��� ��T��v:�ޡ�DU���prD^m7���;[u�mB����⚿�W-��Euy�";���H�|��kk:0�os�X�3�,���P���~v�2���j�)\�����T�r��B{.H�:j:����Ý�܄r.N�.X�.�Bk�u|���w��,��#�����pU�C�t䫡����^��S�[�3c� @�n�#��N�2L����'�pM���l��g��?NI~����'������<�l������J��j�&�]	P�ڼαM��[\t3�ڇ���q:}�n}�[q�D;��:2�
����-q}����	J�����fҰ���e�2����	}Nq��H��e蘅N��R_	�Hc��]|4mG�v��;���fD�}6F�������2U?�TC0Kb�P�r�5�3~Bw�tr�����]�"+��3��Ehzh�R�W���b�ܴ�$dZ�,��s�gկ�����t����;��;�\%N����g}w Ӽ���>�#�[5��\�g�>b\M%UOӕ�����+:�ߊG<�ƽ����gb��P����#qQQX����x�vg�J�LX%K�&��dT��􍢶��7ѧ:�Ly_�NC���v�y_E؎�fRy���Et�"���e��G����E=�[��&=Q��nU��&~�e�Z��+�zX�H<F��ca�F�	�:�r'���
o]{R7����Ȍ���}g�o��\�	0=v�CjG��~>,��AfD�n+:)F��������]Z
v�&j��B�/���x�> ɪ�\k���R*�^�!%Kʽ�np���3-��{�$C��ys�,�(׾�	#���Խ�c����g�ĝ1�<~h�<�^ X�[@�޸�����81����C�k��ݫW]՗)�q��&6�Ddn���J#��{Wi_���fs��\�f=Ҵ�=싃bb}��3k@�1S]�d��j�a���)؈br���	��T��g�	,K��F7j�r~�:5��GHE2k�텗xT滴��bΪ���,g#�GED�;�/8SS�,�y�g[%]L�5��!���M�7�>�^A�����X٨ҩ�l�V/Wu��a�=�<`}וy��3J��@��=
���:��i���:yfTv�����+si���8}�&�Ȱ�����W�|i�Ҥ������x0n��,;�Tĕ]���s\I��ogJss�'���s��?�4t���V�`��٣��~~���x>�h�� w>	Jx&^���f|n:��p/������(oRt�#�"�ۺ�î:�}�ͅ�4�����9G6t󘼌�T��H���}�[i�}:�T�ֲ.���LI��A��׾�����Vw��� 9�y%�X�Olb8�����^�#h]lb��ϵk^D��`��2o�_u�V�ymuG��R��Y��0=^T���iJ�+B����a�����{�W���^D�e�<�nz�Z��;;t{t]�\��Ć�:�>~.�E��/2��@*�i��d��������^���ň�n�/�Gۓh5��T)��ay�5n��g�r�I�?���.�3����F6�Y�Js�]TR��綋�^Z^^��ee��k����p*[a!A"�|{�(!B�޷j��<��*�Ψ��	/ �wa� �{AYs.����cQ7ϴC�Z�<
n#݌.����=��|��8���Q��k8��G�oRC�@~�ׂ�1G{Z��s��9��9�m�����[i�!8���U�+�رi�r��3l�,Kn]����arv���M�o��`���{ɇH�ͭ8���]�vŰ���d6��26��#48���_G]������x��cq6V�������gg�Uh�SFpon+��ٞ^�}=�G����j$Eޥ޸�F-�=���*V*�l�R�ROU�]���,��^3|
����s����󝀋]^�+�o}1��ImIQM��tq[n�\�h�/Y��)WD.W��k���V�R�i}=������1����I,yAZq'���'m]B�(<�b�,uhWB��o���}��%�'�<��/�7U�֔�ٳf!�<�O���<
ޅ��N����CG5	#Iw{8�6��7��L��q�%��.>�-�OP��wג䮥\��Y��^�<=��9��Hj�v�g��(��py��U8M����ހa�]/,SN*>����Tզ}�&w�?���.Vz&���9��!�ڮv���@z�ޡ0 y��"�7���ލzHp�!J��լ�]tiG9�����/�ʇ�_��6]hۘ�{N�ԅ2��n�S��X�e/bڱ㸝1V('~޾>�k�{�ĐyEX�B�t�A=���ف��˗W�+�SuF%C���=q�@�%�+�R���;�E�v����q*���,���z]���+p]�s���I���&�v�;<U֧�
�]��5�prbh���Rܽ��W���6�XM�G?�^⫹����vrV+�c���\����Hj����Y�;��S�Q.�JE�{���xK��%F:ķ|�:|qY3��6��L��3�Y��ց��O��xx�{�#�7��l��Ё�Yxb�	Q+��
Y4�-�k+�����{��tmO�s�%��<qI��u߳xˡ3qc��:����ve1T�����׈�����S�o���r�=�j��ٮ��.���6��6+����F�b�j���Wp;�gNa�����Zy[�j�����Ck���m��i$�m��I��m��m��m��H�[-��m��m��i&�t �J��)ps�����-Ԓ��}if7���.�8����d���6�����đE^�n�Vh�_D{jv������Q;M�uw;��זq��v��"�wL��{��#ٸ�;ǘbwv�,�C��x��a۫�v����a���e�l7�\2>�vF8��d "�o{
���X���rҧ�/�� .��s/S�¯.۪�s�(�h�}�h=���ZV���o�n2�uW%E+���> |>Z�=�G���t��-m�u&��#^!�c��a�q3���4U���gR%��m���}m3�nې.���K&(���g�0��ǫ{&TdQr�� 7cԳ�?�^�h�|�2yo!�o�d�qْ���&"a��o\��� ���*�^χ��5��ٟ�@|�i6!��`��W�~���}��u� �g�a�ϲo�� .�/���;�~�z*g2���A� ɣ�4ǀِ"��eĈd��W�>��)�ߢfc�fg''`�:�՜��lΫ�+z�|�^2�U;Q��3k�;Uw�,&l!�'����H*�^��{�:�#�����7�j䈖H�k���1�8�^f���͉e���}������F�I�nY<�H܁�*�|�'��]"J�ʸN�Tԡ��
*b��:�M
�\���������7��"f;頮�}�3u�ѷU�*-�f��p2����� �=��69(ꙫɱta͆�lV�Ǉ������0E�N��K�=���������=<uV����}��Y�ΰ�z�F��j���W���c׿b���?R�!�&ey�r��̭�}=��8�b��&�ny7�W����lx=�2ܟ������]���R���Qد�3z��I��S�h]���sۢ��ԻFp�r&`�k�+s�w1����#��!j��6"�X��Z��5^�m��-��^��«��`��^����"ҝ�5��|+sjZ�	8�>S��Dë�.Hl�Qܝ��D"C݆�ge����G-�.�mbr7Cq_*��R���_�o�fӡ��{<�}G��ayf�$A*w;���`˟���#4�+��`{���������عK�;����{�Wބb�0BA���l}��$@�T(#�m��Ǯ��k&�ڣGr��}$�>�l��Ke�})h�5���iߗ��8�9��v ��j��3�n�x`���)�^���w���·�VOt�g&>�*����s��?P}�Er[�թ�wD����Gxr��Rɠ�n��;c�j�3LsOJ�S�pN�5<��n�IFl��tŕ�����R�����e���u����z������ϲ��ӻ¡��"e᧋��9�z�K�?>#��WEY��8��>��E��:��yy��>����SU򁀍�s��c�Z�YV�缎9��u9�K�]��k���<>�c�bF:�{ᦉ,|���U��3`���˨C+;'S�u�,����ؼ�Π�A���sԕ7��e_���?r�!q��� ���Ϭ��^"'LQBJ��G��Xj*
�̓�h�)}�^vϏU�Mپ�n�������p���k�0QZ76��.����xaTn뽲�<�r`BDf��:3n ^E&�2w�����l�0E��`*�
��m��2���=w���n]��fQݕ2��s��-X[�Y��D8Ɋ��U��j�G�_*mr���9������{\�'~ޛ���*����.r�y�����Bz��(�7���M�ʞ�]~[���̥d9"_}�߇�f�n���1G\�y��8�Y*k�<�BV~~$������FN�q��8�S��::�� j����w��g*R'³Z����i��O��{,��u��[���<k���R�W�eu+9�A�=�x� ~�9%z�h��8~���V��]?�}����wK��:�A�{�G}�T@{ι�q�z�>ρ5������&���rk����������[���\����^���Z��^r����R�v'�#F��틅"�yeĒ�I����/���-���"f�$�^}�����`�x-[5vG�)��,�m�Hw�݃��ؿt�K�c7���A˻��z���m���WN,��\׸�Y�	��)��J�^�Ë����>��Vy�9��J���y��1�����O@1�ke��m�*����o��]/!q�2��Ҽ|���(ڨ��N�o��eܫё�oy
���R�B����Xh��f"B��ިC��_7Jf	v��{�E�괗c�E̓��U���c��EA~�8�}߄s�eE7c_�L�8rG&��WSX�NZ���m�.��s�\/s�����7vcbo�]�AY�T��2���z�_���un�YP��Ό�m�<*.���	�Y�&�Z��]Gvا��\�U��Ȉ�;�DO��qZ���#Jss���5�@�� m��}C��.�@�N#m=��[P�&�<�|�j2cU'x�Q����Dt��7"�������#(u�\]=�E`����l��պ���V�%|��I����D�^����~��*�f��2���ޝf���g^U�_�s�'aVò8U)���F�[R38�~�$��^��eí��9���8U�KP���>5Qz��Q��aVWh]�${Y�Y����B$��.�5��2�(Ei�ۖ���<��/.�������k����nԄ;s�}��z�S'�`�f7&�]j�xxС��Ḁ�h��-`P�{^�*[�<w�����{vЊ��q�#�s*�7_E�.�i��چ.W��l�[Î�s�`�wR�J��lU�VC:ע�.{K5��ގ��ȴ~>B{z��dz�;�ȸIffa�.�N*�P�o:Ck�_Bt!דV��&Ol>��.S��<1��q������*]Wn�Hwy!���O,�ԧ��5�C��1����mk��6�úpUF�M$�m�_"���ڞ�_W��ʥ��+K#<8t��*��O��������ywlnb�c[��L���"�{2k��aQmQ�V���&,�q��<����kw,e_����O��8�������� ��F,�)�S94�>/mm��o����2��KU��-�{2�{O<S\5�sy�2��P�����r���]t���_Y�hcC���؜�(��}y��1�B�zx[�:���`���+k"9��4W'!\������=��k������1ns����J9��y:v���al��^U��{m7;b�@�,^%�I�}N���H�>�T��Z�(�\έ�	��9��tf��|Vju��d{r���	l���8��.�㲡��wg_�GU���R��h�Y����Wb��2D%�*�sw8|b�GL�OC��#��s����|���������9�e��9�r��������!c��Um���~��z�/mR�M-�x�<�$=t��$�����n�oxk��y�$�i�:�eޯ%���6����>���U܇�t��+�f�2��6[��6⧤ӫuۛy 8�bk���+8�
����)C"���Vʻ�@��'����9�{���F�:_K7=�z}�w�O:�;����|��?��o�=��v�X�ε��!;���������{�m�T�~$}�
���F��O�i�q����ý{=�nȘʥ"(nbKB���6�2��Q�:�;�+���p9t����h�����'a��&*�k�S��V�J�w�@��>-�XÓܑ�Dg r���������2���qvi�À(d�
���ЊY��{~=V��m�7���i�1u����OmZ��ܵ���'�ݩղ���Yc�+]���\'o�'�?<�ܧ��G7Z{X�{w�N�o>��py}�d��"��zX^��P�x�}%MMz��#��=�mV�Dx��!r�V�RT�(���=�}	LD��(�k���7��W�v�o>/q~�x��U=������p���ʦ����?n_ȓ<�`�s��=2 4P�p�oB�=�'�E|u�q>9�bo>Z(S�{Mh��}?(��j8�i��,w���b����հ�Jje�M�����̍��ȧ���Td�~�N%�~�ع�⫹uxT>�~�Q��!�b9�P�7;?C��H<�s��8�r�~{Z��;{w�����Z����Dt�e�,��3�����eC}�u�n�X.�m#͑�Ǉ�.�(9Q�OQ<��ܔ)�*�����339O�q����!L��U�Ӯ��	��ǫ���)���;3y����R��(*r��y�A���a��/B��η����G�-8����}ʲu��o�j������+l��w��-T����|M�v��\'n�}�Wf6XO�*�]��su��B��_������P�(�r�~�$����x�˘o&,�q�t��5���c;����Qj�M�=�<kRϻ������[r�J>��e�����r��)˲�V(p�޶�uxl[7����I{��<��.����OfYe^q���2*�/=TjU�g�m�Z�����ҧ�P
^n�����w�S�!�G~}��E�}[�}yr��䢷]ӱc�(��f�y�����g�w�<ؕ�&���Kcٸy�����;7�Ҫ�QY�.��K�T�� g��4+ȱ�$	O�X�\	��L�>z�ȃ������; X="g؁+�]N����૟b�\&\2��7����+1�?�"����?x-~,%�N��SV�{��D {6{G��{�=;��"����1��+�ި���a�}�7�@�Ӧ�u�����N��
����	�i�R�p�_ٓ����c˘� ��M����\�������-gB���T$�f����˾����=���K�2N�:p֊��u���-"�n�@�1<k.6o���V��a8)l��5t;�GrZ
���ټ���ƣ�h�n.:�����v#��u��k�Yب�;x��q��8��qo������mw��]x�u�Yき�b�v���03�>|���%�/5��&E�OX��յ�T����d�U=�#�Jhd�z|)le���┠m߅�z.(h�c����n*. z~����c�L?���������x�}�d�2�O�|.s��=��:�SF�)�qP�^P6U��_G�˝W��p??{����MG�J�׽T��p���E$~97����^��a���c�,[�A���}gL��l_�����N��b��ܟ�u�����-ܟ-�^���:��I���U_�g�%����j�e]�M@!��g����{�O
����<9Ǽ�6�)�3S�"�>����덺�+�CǇh���M�s��r���<�����A`�rT���Q������}3��'�����>�0����?N�߽W�U�)��H�q�F�P%�RO�����_��n�ߛ��W��/q ��E���pݢ+9Ӳğ��q�uv�i���󗹷x�-9{InfC|�rѠH	v��lVscz��on��WzIdu_Uu���ף�^���m��M���B^EA0錉\�}��K.�?�)�����n�S�fϔ#�9�{�.�T�qcf�].�8��uig��;��W	d@7��v]�������WŠ:�?p�E=Z�bS�qu�R�B!�l� Hz}��J`%���x&i���gƸR���,>�H�}sq&�����\�'"� ��a.�aX����ލ��s-Q���[���?z�W)%���w#���������8R	1��]"'����d�ȸfz�1O��C�u���B��D�:��������;�/�N�mP+�'](�"ǣ�5����8�!��dq��6������g���&�f���z��U�\/SC�f�l��u�T\D5j־ߖ.nד�X{��ƒ=�g�m���r)#�B�r�d4e�8��/���4e��6�z��/W����q�MEL�!�i�v(���H��M�7ƻ�#��g��GYʀ�O޹��ױhxΝ)���� �_C���pxT�o��Y�%rF��1��{�3�ܧe�f�6��g������g\�{!�����	 �Ğ���la���|���8���C���H$7�e�8;�Â�/y�JG��Q�D����`f^m�l<}��Rw�͐�v��4�����ח|� �W]�ʸe�����^��kW�8�W'+8MBy
՗�fK��+��s��8}b�n��~Q�-g��(g�n<Zo|f%�S1�v��Oޏ,���]:2:;��h8��kN�z�W�!����,�ş!�(��}9�I��y;���`�d;w]R{��N���>���{�j��:��L��2���;>�~��yE^[�u	�"��l]���Mf��H��4|n��I�9��c�_��y�I�1�M��aa�C�[õ"�.�2��s:��_]�ՙ���I�w���:��CS����R��JC�+V�֑0�k��>T�Sݶ�:�;���k,k�����q��f��Ti�+T����t���\{3~>���e�h��f�w���Ѐ\(@|T����Ur��y<��D��g�;�t�s�+s)�νyb	��<"�F�!^7e����_��Tٙuo��Q7�J+���h���e|t�|��_��f���9e�zn
��������'�77-_aw~uZ7�rIrb|�΋��N����t��<�����[��YG�~doީޚy��p�M��͞��X�<T�$�)S���s�a��D�U��ȏ1� ���C��t��w������:�{`L'���[w�t;��`ץ6:P�PX�V�"�E6鎔;��bU3&��t��y���ޔ=[}��s�/��2�^�k����d��Tr$7��jC-E}�ة>ޢ�b���&�.�N�	Κ��I�z%$��8��T)�sVլ4@���̹��5/�(*aV5�l�crP]˹m�!���wNh�Q:ΤQN����76��/��Gv�P��9�a����'1��Rwb��Raӭ^��+���ԨJ�R�:j7�(��wu�9+�F�Yy��'��=�L�����C���k��	��CA�i���۵j��у��3���%~7�L��㞊*��S��j5m\h{u�+��v��O!:���B���#;Z͢�K9�N�&�v䷶�x.ʓ"�������K��x�`l
`���wU� d!����;��2���GޑF+�ޡ8P��"�>�X�F��4�;D�)�{���c�+�)�G�sHW����hOM�~���kAw�pqnvc���0��0d�)C�~?93uԆ�+�������uMkt�.b���;'z[q��l��6�]R)�{�qo
w|]�S-�8����ƛ6��s/.�h�$�P��y�5"q��K�v�cvV1���a[�Ӭx���"�33o�QY��� R��+Y�>���d����Fc�����h��邟$�>���xz��JG���fg�k����8��"��1܌?(���*����Q	)�ڀx�����p��c��S�*Tt��}�^���,�j]�,�nN��ur� ���%$���w�Q���|�u6��ܙ�������3���ǯ��<�of�����O),��0��IswN�<j?���k�`ܮgy�J��b��xJ�ħ�Bn��-Tx�^���NsM˗�������o��@���aD]�,�J�ܴ�v������3-�x���-��Ɍ��N�z�M�v��M�7�|àh���čͫW*�1�'���x�zg5�.a�-�X�jk�Օi歺��CA"yC�fX] ���sB]wWxA3(��;���[��{8�"�k������0�+�<y�>L�ug��%rZn��(���<�wK;:��|=���g��}��woa��
Ǉ�LZ�T`�{ ��`5�Z���ϖ�>���xQ=Ig")z��q+-�(� l��֎(�  �с���|s68ǻ�1t8c��1)p3�QM��=�n=6�r�����,���x�]�	�^̿�G�_��v�B]X3��{mN5�9ҝ�I-���^L:,��2��㫎<ƒ����
�2r�{.�K`	�G|{�s���pjB7�D�V��/V�8ceT���^C�4���Y%%kU�֏۹������h��ղ)O�4RҾl��#ǲ���Z�M���W����~���&���^9���W�&��ŕ��0�W�.FC	��ʝ���D�Z�S�� �f�R�,30�:�{u��C���3a�ܘ._�ܝԢ���ɲ])�\Y���V>�Un��ؾ���9r+O�t]A�걖����}�
�*��a,�*b��じ�����	Vz���\"�++6k=�ӞQ+ǈ<&oz�}9��״�d��r��7��S�2vdx�1\�X،���[Q}�w"��_/�t�-���As�F�9�p^���>��:->�bJܫ����}s��z������m�uG]��BK){��+r��u�ɣ�]�+Ss�]#j����N�x�5���� N|���	����U��S|�z�U�V�3~�5_V?�m�7ެG%�y1>"ĺ�8���F1����~��,`C#��gwy]QT(ZK��`��Ls�������{gi�Ʋ�{����*��@B�*a�Ǯ����|:`�[�%���G5؎3gE�^q#�ʻ�^�y3c���%.�~���WtφNEj����3��7Q�]�1�=����bT����dr9����ݩ���]{¤@Y!��G�2�z/����y	��&wUOfn��c��M͙%�UC�I�N|*�Б�㗁��]��{�*u���"S��X�Dv�>���L4i��:�o��w7?oq�+�M!ivU󰏺��Op��7���9���eՕ��v.��C�k/���]{��xdtK����sH�P������H�4��ӂ�j������}�N}��b�T+=1p*>J$�4:୞W=��b%5�.����&�7>^W�N�v���K�g<}�,ӻ��G��k<,H��r���ˌ���ꐫA3q\�Ǳ�O�Y����ǭ/��^�����g�V�:l��Hu�]��҄���	e:ApB��N�=��Sދ~�uG�w�L�j()��׷��# i���G
���h�*����蠝V��I�kΞ��\`���yj�k�<	V��I���7��T�-N�m�n���w���Ϙ��<b���s���lJ��I}��s>0�W+�U:��iu{�א�{���n��Vk��A�L��{�.�tυV�D����)�����q)���k�+�3�� l3��E�x#>�OP�5[3Uf���jv�����l5[j���u�~�iO��ۆd�8���vV'ӹ���9$"��'i�{<j�^>�.�w�}�**<���!�뽉��m;;��sG�L�3��H����Q���� ����o\�[u���L2�v��\�`}��^{�Ml�����s�� ��A��3���AOw�
_;B��3ޏ@�ji��ee�pʳֲO>7��ꍻ�ު���0")�ѝ����;�V��S�X��WY��*؆��Ny,SO3��d\�N��a^���e�w�sZ]�dEE��`�����aT��9`�a]	���I��I6�����BL�/�M"�3����0<�s5�/wyb�ВnR��U�3�'�I!�1��e���ٝM�mI��~��T��Hw�z����{��s�GT���oMR
���Ď?
s�*��o��2o6��e�=��w"8e"���LNi�b�G��������/9L�:M��:�ʶ�q�S�c:��Ӭ�~϶S����@�K}wC��AnO�*�5��o5��J�D{|�+p�/F�k}eq��SM�*�P����͝��P�e�fi��SK`rQud��S�Fec��F���J$�>né��n������ǹ��=�n�W��i!D�@ogfF@�[=W�}�(�֚�G�K�ԃ�&G������Y^�6xg�gf�Z7s�l�3f����t>����VOcڶj���U�6�@�Е�׷v�
��V��H���ٲ#�����F�;4#���z.YR�Ñ�!/m,S�k,��/9+C�����I����
@W?*���B�{�"ϓǛy������/k�"v�)A��z|�{Kǝ>G��)p{ޞ��3��:��3��zFkU7�cV	�0�W�+r�c�U�η��_&s�{X�mD������˥�~P�²�-�.���H�͊��N�pF�^Un�\u ̣�m��Ý*Z5��2�\��.��0�ju���;�4���M�����Q&�S��峎�'s���&+�n��!1X��1�u����h쳤������P�G�]0�7I�_�;�R�5ܗ׬e�:'�2�������q��n�V;رY4�j�z��=���oI��
���}���wכ�N�����XAML�q��<���+vt�J��,�LI*�KȎ����,�ނ�;;�Q~���Rڏ�jR^�w�C�M��oI�<�=�����U�č�{b;�KRx�V���qfW02���FR��l����L���i^G��N�|6��O�|�@ӯd|�L�u���۫�٧)[��t��$�WYWw����z��C#3/��ޅ4+���QYJ��^���*�#�s���i{}Z���cM ׎�V}�l�b��q�@����&/kҒ����;+�v���!��c��|�b1�M��wZgc%��c%�N�ӛ�.mm��ϡ�䣔ѵrr��|�y��{&��FS�G��=kn��>[5`j^��F�U�'�@��«�M� Y/��o>����+��罱���ߞw�z�c���ޮ��n\Ё�b_˨��g�\�;Q&�NN!ߖ�s9[�~�z8��ܭj).{��~9�*e�b B��U��2�};����ך�~���D��Gﭹ)�E�9k�_�[��2����`�	��� �<rw��$+M�H	��l������f&x�8c̬��9�_'��9s�ҥ�MJw)j�#��,`z����=N봐����"-�;�J��r�X�����D�9 z �L�ˤ	(���e]�������m��K��E띒<y�5g�[�����iN�]|O�ξ��#DR�镱�jf�CAqx.Z=>`������=ҽ����3&�(ڙ;��==�T)�\jb�[jȝFy"�s����PRB�Fg�=�j�R3�\�3&:S����7E�ך��"��u��iN���9]W:S��G���M3�4�۱A��(SH\�P߮�L)��=�z2�j����и�ql��а�L��������yu���8����$i���ow�Z�\0�|Y�~s"�����dU�ד�[��)�ܺ�K*�Uʘ�SZ��6��1W�%��do����I+_f�O�*����V|���'� G�V���U;g�j��d�{�"�������f�s&t���:�m`��B��x��H��T2�e�w�;m��,��}�/MB�7�>=B�]�JL���|�k�'�C���á���AH��7H5�z��1������Vx8�>�%��J����!�>R7������B�����mK��_Sj���~�E�>���9d+����;�e�	>]���u�5q7�G���jj>S�%�i�a;���u�tKw�o����{�߁��*��֩ A�#��kJ�/!=����F]d�:|�\U��a����&<��X�.���qP�3:����D�i<\�Y-PJ�׹�6�.�Yv�j�/@L�]���v:��%m3���_���v�]��^�[]���7\$���
_Q���.`�	,ex��7(��V=+��9��]>:�3�mY>����ʀk|�\�y�a�{�o�f�ә�qP��;�G�~��p�Zu������%oֳy�ڻC/�jHR��>s[�����P��5)�������{�w �mu�X�,iy�-ͭ���'����ZG�r'�;"�T;�oףמÍ�-� ��w�����/k��/ƳЎ^M�ϑ�x�h���?]���\`%�f<r���{Ʀ��`YW��gd��8cذ�c�f�*o�fV�T��>f�~ܻ��˽���jS�}Y��#�|��d�=*�(��H^n�3ł7�{�c�g�A��꺝��;6�-�D�i�7�`
��z��[�A��y�x�j��z�5���t	As&u1~���G}p�Du��tnջ�Pݜ`���מ����I=�n1+T�W2�ۇ���ܞ5'�l�ZW�~	�*ԲE8�b�L\!,�
��@�Ywѣl8^;����@��E�a�F�a��'��R�X>�����Tj���y(�N6�)�S޲f^#K�(�!��Wb���u����'���;st���|݊���ߛ��ǫ�E�:Tp�;^Eg+�3OO�FVc㜏f���yh%�����R�����ɷ�`�*P��;0�N��;<9�W��{�I'\�i�yk7Ūd�x���X���M,��#4%�8��E�]0��j��gb�(R�P�Y�m��s��ir���GZp� ]�����9�f��Z���0��wv��M�ந���[o�ϓ6�k9��߾����yix�zpKP�s=���o,���r�y��u��l��u�����}�@��t:z3>�Yit��j�,�(���{'�_aAQ�KoԈLU��v�hrʠ:��3ʳM��l z�ݼ��G��j���c�3�:��.
�e�����`9ʮ�9��1��n�VE�#a�|5��ĺ{�����x��a�}��{+3��Ej�����S}�"�s2�z)��k�k�h��`wS�'M��N8�lA�fV�v
��2}�Ղ�J�8��|�
7�A}"�-`�c��]�����ΐ_|�����
�x�o:�x�7kh%�4&���7��z�Vzݴ���w��(��1\Wm�_�-��߹�l���=v6w��X�q��3�l��uؘ@��+׆:��a��L�����}W5�Bq�W9lY���si��c��Z���
�nu;���t �����q����4v(�3x��1Vޑwt�ɱS)_�;)O�Y[wV4w7� J�+�s���t��}C�U�C ���U�I]���v��w;iR�X-j�=�7�����(r�e��60���ڤ����"��r�U�8�B�i�M������^����Ëq�l�B�N���X2U��qC��r���.zY��{1�Я��������X)��BxL�kiU�t#ǔac�ԚUB��3Gb�àB�8�|�@�D����Tz�f�TM��=�kTXU�g�*^����A��`��=Qp�ې����ز��)���J����,��[��yo7�m3�.��C�b�Lю�޺��L��G�v�����9ӻ�7{�x���o�c�0oc&z1�o�Hs��=Z�����b��f�:�~��4��Yy�}wfsR�p��X���^�(�3|u��Q�:���7�>��h{�ɴ�N��}c�߯���r9y����~�+�w�;�l�|����q�y�C7�	�|�1%eC������~뱷]-z��}���|V����/�cL��yNI[מ��k��j����<dVc�v�>~�c�+��^�6�r��1����3���}q����W%���ۋ{�{b���0�vn����YY=��Y�ɡ��������
�nO�����˓��7�2��8�eY��#��X|�&j\)�<n���:���ty�M*���_!�1.�� �r;I�:]i7F�K"��a��c�˙{�+�����a1qT�jEs�Q!�4�-t6��7�U� g:#nP�z��N�e``t2�����XI��+�zOi�1Y���,�������{�ȵ̲��\��}�MpmJqe��g6�$Ԗ��ž�Z�e�ѿ�M��nEmy�UNںu3Z�W3��jN��)�0��^����BRv�z8b��VLj�U��s��7�)P���]m��ח ܸ�����Q�n��(��U�W���Q�UgM+�U�k0\�s] o���ճH�;��"�G-��<�w��]���];����ӽUpQ������|���[wv5ʳS׌+dC�[I�ܾ�o]�oѱq�mGy��4>�w�y`�;�PR0<�0DI��	�	�]�ío����Tӏ<� ��e�η���pӊZţ���g/�Q��H��&eEQ�`9ޢϼ�9.��<')Wn:+3�ɕ[�/�pK��l ҽ���o�2:�-ϛ�ni�k��Sb	���9w1�sM�`�ےc5@]a�K�ؼ��T<�f����C�j�R��R� �+�N1g^�lutY������ƪ�Q����jí9��~����I�zm�+W,�C�T�̞�=�c�g�e&Z�I)�~��J���>�3Z�a�6[->`����]^�J�<k���E��������W�9~�Kv�,���G�浐ѣB��	b��"���ƽ[n�i:����i-1�/x��F�mX�PO��w>���яᘻ�ܐO������W|&��xbާV��m:7�Ր��3/��5
������Na��
_U��Q<�W3�w�Rɻ����oI�|f�� <������
�W����-V�g����D�L�ɼ��J>�j/�r���w���92�fLRUP��l����!��JvuZ��a�>��� S3~�,h3��yB�ycB�yO��\�ִo3X=�s�L�?,~
���b/e��+N|}�Z}|��G�W*���N埄;^��cd���u�qW���h��zW;m��:(fM1�z��ߌzH�>4���F�c�\��*���Q'w��G^ξ��V2orUU*��wz(t�UCU4��J�����S��(���vJ��]CV��;�=��-���}��_�Q��F|fBO��F흙�UT�Ԯ-V���m�pm�P�R�r��l�1�X����SƤm�����W|�o#�Y՞k��NB{e@7';bH�Q�uc^l��ҕb�IW�ٜT�u|�y<յf�\���'�����.�2�۬g���E��I�yg��1Cj[���̟m�^�R�1��@�3 �C7ҼQ֤�
�V%;tD��yP���0����N�_��$�׫];�-����!����䴷F!�����v�Zp~��:�;ѣ �9�K"���b�Ӈ��kùPs�;�{1Մ��ML�K�,�ݮ|��x�-����>{hV_>@�s�#c�]}1<�+8�1�&�&Һ�M�ؑ�'�9���$?m`�,�: c�}:��r^,U(Q��l�䐰��9y���;J���T���MU4k8_>�M͛`f
�#}��;�{��4�Js�ְW]�*wX���6p|��Ck$�u���L. ��e�Z1���+��V�j�a�ʉ))��q�jT�'�Z���u��4�eߠ�R��n���+��y.�&�XeB�k���e�T��3� A����itw�<��Q� �G_�G���#��[ۻ��,��;0�9<R��y8p�wS]'�s��n�;B9����9J�f�L`λ|$]h}j����gl쮂�N��mg��K�;5��Ǵ��oKF��E4����?��ּyOl��^Q�`�Ys�p)gk`��X��%:(��9�7��X���f��y�-;翴�!��`�̮��Ȧ��Ų����˥��ݹ�=';����ɜJ&
s�K����U�yO�
������d3{�z}a�Or�nPs{/C[���ږ�eG�-i�9�S���wA�Ьʧf�uxA�w���]�sa�Yػj�ƫ�@a�Ήһ��tFkq�����dk�w �=�0$�N�zf*�8.�'#D'I+��+��Gp��6�
�j�X�]���9~mN�9���㉨8����Ǹ.Qu�����6�\6;���s�V01g�$�q����ӻ��Xs��t����3���<钦�
��`�E8ݚ�5���"!�VY݌I���u˯�ۼ�� �P8��û�fB�Y,��%���HV��m�]Crn��\V͡������U{�V��a�uR�t�Q�P�(�l�5�����1�m���f��[Z���o�G
C׏{��`���	�����Ԅ�Z��ʍ�-�y���	]���?9ߵ7�ٮ��u�*�(��/�W�ZRD͠p�:����;_	��(%&�7|��͢��b*{���+IJ���/uf�Y?*6"=���}k��Q�9:�E��2�esMYg�S����5f@�q�Sfݢ:VYOp��8f�0hj��dRt�=8�\/�\&(�X�y+M��a�d��b�]s4��(TyȻ���)ҝw��2)�n'_-�^N�혨4�I%m��i$�m��i�m"�m��I&�m��m��m��m��I"zc��i��o)�a)����+b}ᘲא���PA�?
ZK�s��]߈E��6-�;�ǹ�9�+O)�ǂr�k�C���/gcF��)	ʜ���8���'�մ�J��Rcy���g2�/��ŠnΉ>z9��A)u�&����D��X�t�{N���W<ƹ~����Lu���J'����
\�H���J�xjPa�7{��{�ج�,�Ѿ��w����^�o��@���o����i��mwCSʟ�`�v�QAo�}��A"��(Q��I4�m���L§=u�.?�[H�V>�
v�.F���q#�wӂ�����Ǽ7Ý��ǫ���l� ӟ#雊}�yq7jh�Nt��3���VWMR�x!~�\�9+�})�l\'+���K8[�O��n��[f6� >�C��Vn�<fr�x���Y�@RF0+!��]z���=�^�h.5y�<ڇs�NEm>���#f��ܮ�Y���3���}�f�R����x��|l{A5��}�\��D�����{*�j�˞e��x��5�c֝�G�x�	���x����9$܋k*���9rn�E��l�����YH���y�j�<�+ϲ�����2�v���?������������X�͡�j���=�C�Q{����}�0��ݯ��v�9�uĉ���ղ�s�«�o0�.�yb�i�!�1���Eq��l�����#�U��h{g�_D����{ט.�*�6�j���wŲ��gƖOoI!��Ͼ �Qn�m�tk~��u���"z,g�p��^����vҖ����C(��YX��(������+{=|<����[��W0����̠�F���{k��ޭ�y�B�a�jx�~�t��:������ZuS9j-�~7݂1�,LtG3�S@��X�
��ѻ���z���A�}�D,�Ajt���Ek��=T��=Κ��^�]%����=�:���N$.�{� �P��T܎椾cj�JO����;3n}qr�s�%u����(d����z�<�Hs�jX�n������D�N����E�u�3%I]O�}�-�g֤i�ޟ��nE��E�<�/4�/�莮���5Y����f�nX$�EV�s'����*�������sw|;3��~Bs�����z��^ǹ�/������׊/��I����/Ľ���<nvO4�_��o�hT���Ʃd{v�R0<��s��X@��8��!��KՄ�;�K�OdL�g-�y�VV�����h�����};��a���N�@��z��ܐg��i*��>�~�K�_Li��V���f��^{��6��$�V�څ�X�z�Cˉ�@Ȯ��D��m\��Lڙ�_t��^����\r�f�G�ޣ��m$��c�k@�(��|w;Q<�NW�18KV��W\ԣ��#�
rKw�#��y׺�[�����Tޕ/���p�n�Xc+��~�d��^��;���uV⨒�*[����k��}���!'�H���X}�*�k}��ښ�Q��x�
f��fޫ��0���񻣺�Z���T�X^���/�_���w���d�[�|��n�*:h6b}��[�k\V�S���V�*���Ȟ�����{��l �k]4 b���]��<��1vq`6]5�\[�۝�����#�P��Q��x({7���齫�k�)~�sVjU���^�=�_9j����P�\k�w�8�{���UDj��d����ڣ���oK�B-���B�
zΞ�Q�V*������L�ǣiy�fRI!юWU<>����z��z�	Թ�5�) ow{���t�����o���C����>����#�>w4�����8�F�^^�����n��$!O�V�I;N�T�׻��dj������M�;ON.�YV����Т�(j���UT�z��MS\�s��4:%�����c�R�}'=of'Q��v��K~�4}s��J��N6��"sqw�l��򸩭 m�w08�jc#�er�t�q���H�e{.&��v�	2�U�H��u��O�}�:�=����Qg�}s�����C����W�D��W�����yA^.]�Ȣ�$�N��>��=��v��q%;��QƧ����fz��f��~� �Ĭ�u�2q:粻|bU���~�ʩ��)%+�`N}�P�QTD���AĹ�6��$��{~5�d6�0y�졵^����\�������yD���U�A��|�P"�1+���=�U=�������ù��g��v�&���Q����~D`�T���-�=:xְ(��H*6�8�vD�J��<n�+�����L�z�׹�M����G��+*��ww-Yk/+��-��M�>y��T-�Oۣ}2?Vfo������ף�#G8%�A�Z�!B�ŽF�}���aa�+��J��MH�FO���N����>b�nt�}b��&���Ӳ*mE��}�A�G��O(���:�'^8�ˉ�BYQX�����
�*̩�*��nYM�i_'v~o~t��-G��D�����k/��y���h��{tO3����!=��Z�>3L�,T�>q}mU��</~�FO�D����Ե)�d��\��^`[Mo�Wx���޹t�(�3�?���yb�|Ç�;��>�+�h:��ʣ[�S�TWC�a�G����<���o�s��VP����p],��ǳ�"l�L<���y��9��=��Uq)nm\�kt�Q>��b�U��f7m��y�A��As9x�@��_g�[�=Ĝ/z���A�D�yI�;�=�*~����N>��iV<�2��^#�,���N�:��^~c�!��T�o���'�9wSCvn��Ǘ��
�����z�^�c(V]C�\J�`�駰n�ذ��n�Y
��>�;����>�ӳ�/���3Q>5o�.����S!\�}�b��L�ͺ�-c\Ν�v[��wt5�+�G˾٧	bڞ�v_�{j_Z	UjWւ㙝\���R��nt%�N����Z�k�\���ů�:Gap9��8P3Q�Ek��#�	L�4��ܳ}�G���oS�X��fٽ�����������^�Y�[����fP�; ��sm��m��wI��sL��B����PW�˯8"�+$����:�Ot�W�V�%>5�F̠:[��'L���������8�q���u�(\z6
�ӹ~���j�ۄ���='���Nb@4��X�����`�f#��l���Kܥ��ƳɎ���}���GcSk��~E��|�:Fj���`�5P8�.����\t����ɽUյ��u=�S�N�t�Oc���;V`��Q�Y��	^3�>w{�?|'�z0�J/w�V}Ԉ4�v-��,��p�xlvxt��~TF$�/��K�C8��z}�V�s^Ӌ��G�M�~^��f���f8;t�1���Q���x$ɽ�K�Ț��4��v�!UY�55��M_���.�$l]\y�����,T�����BroוRN	{��3�V�W$��aͣ�{;0��D��'X���[�>�L�qʛ���Nj��U`�g���Nz NZ�Q���%�׹�|�7�أ~��%�x��.���7����g�/ ]���ʅ���+1�TvFc{7w�W�c�&�~�i���z[�Lzĺ��O/`�ʊ��WK� �5�p��?pذ��,��3��(�����z@�7�S���2�ZQ�B�����5fܫ�/5]�������羆>	P�x��������ЋSb�s��^��.��>�9ju���{�R�!�7w���WaǺMp;TФW�(��w=Q}��6��ٚRy�n��Y]�}��Yw�m�\����{|"W	��{��c�U��*�g���Xkp�p�}Q���Ifm�`}-^Ӎ�a �n�fz��μ=��$�A�B)�|��g�6��GOő��f �8�1�elu��k�����[\}�.]`?i��;��Ǆ|���o���N��V�$ws��6v��7Qq�E�Uc��r��%�HX7�1/Y��v����mg��Y�;m�sg���	�'�X�����Ho�C9��W��mj5/b�v+�.�m�*����*K�Co�7^�3$��jv�q;�uǙ8���y�����'oڙ�l�껜�M�}�3ʲ�V�_o��ɓ�W��}u�\Em��m��2�+D�v�ZBpa�<'��s�둋����˃�=���>c��7բ*��/fDaڴ;���Qۮ��l]b�Mh�"�ȝ�U��~���L�-���O�e�εi��
���Cs��!�)��ܑuº�]�R�݊�[hR��&Gu|���_}�ryg�В���rm�*ޔ�y~�Y��qz[���� cC2��Ѹv�ImZ��9(V^�y�oKdTII��C��U4i��͍��[H��Ȱ��Q\KdNa�M7D�K�N2��<��H@�������<�ṙ�Ы�ʣ�ӺҌ�Q[����s��ל�L{���wQ��f9�;��]�ܔ����p����R��4�-A�X�c�yZ����^���}�wS��ک�11�:H����DM#�����ǖ�N)�SE_o��{��7�	p�no�;��(��'��x�y�r{ӑ:�D�W�L��<�4����t�p�0����]�پ8ڜսb����:���"�(2Y�a��7o�����4/L/J��R��ǯ'�}�	+��k�j�|��V*Sjr:�K[>J�{6&si�}��j��k�'*"7��嬮��]<��N<ūsg'3&�C��<�(x30��US	XX��dLC�SC�Ձ	Y�QcyC/#��a$[�IU^/^�Ǯ��<��n��g������P��3�xo�8F�{6�bߜ�{�3te���5�Rg}1���տ�e��rPY/L�۔�^�*\[�]��/')[����d�.-��W�����f}=w�?��^2�[U�{i}<���f���׌e_3O�n��~Ô�����6{O�[�{�=�dz]b��%�я/y	��ת6��!-���o*X�x��Ǖ�td��ل��)�u�׺��Ȉ���L��H\4/_8[\o�/��&Uޒ�\V*lQb;�w�$]�4�7qnQ��dye�{(�I���n-�+ΧZL��ܖr`�T<�Ou�
μ��ê�{sy�gSAPv�H��!v�S����kJ�r��2�c}��IS4G۶�'�:�k4��$�O�m��Ury�\w/\�_�_��\��=]jw�t��D��Ke��t��Ϟ��^����iU����8����"�
��z}��7]|�6w5	ؾ���"���{G㲊�,\H��j�΂���5;�+��O�U|����:���O>k�!��fx���JZsgLO\L�C�Q�M�ID�ۦ��T��EWq���W�Z���˃��m�<�Ga���5ĥ=�[՜��H�oγnqg�&��jp� '�餅������������T���bd^�Rq�M�Zq5q�n�V.���j�s`8�|-�@��U�&����4xGb6͇�߷�F�+����0]z���PCݸ���A9ۗ��VԌƬvq>p����z��&�]o�6�r�w�x��O�y�-H�Ks�Vl�P�,��HÁ�g79�vk�wN�;���峒g���χ�ׁR__�8g�W��Ƴ} Sɺl�\�4�V��ʡG~(|��Ȩ����'~���j~�"�E�M�(l��'��%��I�/h��>'Z���L�]�fM��
|�a�\��<�T"��G�/�.<sq�4�߭�N�}^��M���dw��~7,�V�,�۾�k��;AT�����e�8��vܼ[p�IBh��a|�5c�ۊN�������Mf���a���m��QP�\���-6�m�����3(�ɗ��f����vypK� ���*�[������0��w#~���y.)6j��Q�Ǌ;@��_�E�臻���v=�Z4˷�5;8O=uP �	\[�W��<\�P��B<&�c�ȇr=�J���kq�Q�~��>��p�ܫ�+:�L�*��~߫,S� �JI�%��Ư:�w�60��va�o��V9�f�O�+;=[�w�����wv����(+r��!;g��~�\R��2fS���k��YW�=h��z>������1?��8�n7�����7�׊@��=�ʥp)�S�f������g�|�frð2�q���D���ub�ٙl�{�R@=1ҥJ��.yT��k5�S���~��s�ĺ~���*JF|���v���W޾���>g��Hy�~�E����o!�}�p��|��b򘾮������m^<�N�)�Eח�^�|1��}���Z/e��^�] GT�yH���\�6Q�>��j=��-[aw�ݝ���=;Z�5���U���웃X<l�,|����6� 7ٗ�n)��Q� �u���s���g�R��P�ma��O�g<ڰjDA����䪄�D'�
5�z� kd�b,���^���7x:q�}�j܍vU�m���u��ޣy�I[w�0J���;�uѺ��"u\5��T�x�0`�8�k�uv�.F,�t٬�Z��o,���z�N�� a�w%7��={�% *�%��/c��9� J,+5�&��ZϘ�^I��yJ���R���ub�|5��O���Śr�|����8�2a���ϥ��Z�yj�hxK��R�����
)u����m�s��Z��.(=�*sa�����9EL��)�"���k��Y�gGh�>yh5Ru!�[�Ĵf}��Ly���E��>d����#5{� �T�vm�_��y�T0���to+�7���y��+Zx�*��]���&�/�z�l^yV�KחVƯ������jt���w��7�$��:��ʵ�u^�>�.a?	�+sm������9�6�;k��;M.>�M8�1yq�����W@����t�X�����0B�z:���m��|�2���="W��)G��e��0rV����əP$,����wi��Wb�Av�j���s*}Zh��{~����(| 3�^qQ9�1TFu��7r��<}�����1�J���T9�*�<�r��Io�Te����'�}
�t⹈ǈ����ԟz����nV8;�g���@�J���ѩ�6�t<J�c��g��e���v\ǫV��ώs�Ȅ8��*��&`J5���ܫ�UqK�Mud�O��v�����偢IEV3{����|*6��Q�Qs��u߻��×VQu�Jb��OVw�|7:�p��MX1��/���M��Z8�WH�r�MSk(���"�t0�p;�=XğmY�j�N��i��tp꧴6�4��Vǹ@8�6�R؋�w�����Z�JU2�P���ۇ��+ՊӠ��⥷
�Ln���}gj��H��C{�1}C�
>��C�˽�\�ں�:�}�����7t-��݂�'3o����v`T$��[��k\a�q$��a ;��[�E &���m�Xq��^o���1~Z�h5��茰��s�+��hr���=�z��>�APMг�p��xÝ�1
a֔�,=ʨ���6��7.~�[aM^}y�Ì	o���¡!'�@3��\�u������@�˞�9���~�GVk���JJ���e�iT��S9]W�V�ޓe�ϫ�c��Yj��_���7z��́͹�����a����^o��s�us���~����w�Ǆ�I��]���^<4� |XV�'�'�u�*�΂:���|G�t��U�-,����O���V*U3�&w�u��\�n����t~�7�����y�����bM=7�����;��d�\��T��:�-ҨR�ݘ�]Y���%�Ю�c��������t��X ���!>`ϴHE�d|P��d3/��WZ�޾�$Ͷ7���"s/{w�w?W�-lw@��Om�/v��ܪ�8�oy'�Hd�H|��y���ь!M��(�4ì�R�o���Ւ����s��ː����IY$��j����!릹��=�d�I�y�����9Yi��i�y���@��?���!�7_[����=�t���C�
�sX)=��z=����|;��fC���װ��q��$������z/��B޴�5�i��k��a�I�a ����$�H��

!%����ÂDli௑�HN�&��rt/+c�T�.R��=��%�[F⒓�{�����AwC��v.�H�<�ɴLrpZ���+��H���1PN���z�F�wn���<��F�����̬ˮ&5	-厎����`c��3�����l.�71ю�Kݺ��Ib��]�"� ��엄5��J�h�g\�T�݋��K��o1��r���W�M\��E{�8jݞ��рo>��b�c9r�����Ͷ�K����$�ɭ�v�˖��4ŭvsrm
��f�.N�§���F�ee���p��w^�V���p�+���ǜE�"�pnG��	�eG�>�4���mb��W���8�u�e�kq�˭F�l��u��6ӷ%8C��t�c�¤kuq9��,[���)���9�Cvwh�N�<z`!�m��_�&X۞]�����x��n��ݨ����|�0�/s�S��-*��*��+i�,8G,In&3�6���q$��Ӿ�|�F�<G�7�>ځFBA�E^�[�f97Ώ�ܢ's=�Z��I���<+]�����7���w]�1ޤ&d���V�h��\O'%G.s�\���]n�%�6��ה���#x�P��2`�����w�(��\a/���� 5�{��m����h΂�����D����&c;ˋ�6:�
cxN�9`�1˷0��2��j�=c>�0����y�9�w�zB��g�Ҥd/����b_�cZ��}e�ι�zoEn�x��.�Y��^̫�=94i��NlA��sU	�MU�ɚ��A��k�a} uh��b�7�;\��{/wA�[=�Yn���@]s04�bXr����oç<+�\<2|n�n����Ɩ�aٚ4�uouÁR��Fm�fDl�zH�N��a{��7����������a���*��[+{=9u�wK&��S�}�ڷu�Z�\�^y%�� ��#��m̫��Y�z`��M���޹�*��5��.ԸNr³j��fڝ�Ӷ�(7f�3��t�^ߖ��O�G��T?X+YrV�Y����`�{Ց1%���g�M����c��}�[� ���_��絫��&���������['r��ڼ����7�/�M�B��eG�����CY�SQ���Lf�
���i(E��x��љ���r!�r�$;\>�P�>u=�2`�>���ۉ@���cS�˾���0u�^���xe�x��P�}�8r���am�C�/�����|%�6��SL��O�.��'�2��S#!�oR�ySܶ�M��� ��7�`U�?ǯ^m:��'��q���=|�����y�û��Ύ�]V�x��wt�}�/tv	Y9�b�lH�6p�į�:�t���%���ڽ ����E�שEm�˔�U�s����gc`�����if*5wc���^m�����A�*��^sDMh�$���˿�����1�b���-�J���n����/�v�W�FW�IJ��	�ȉW��QSO$�dV�����o��lF!��ֶ�^�7�s5���yD Ƿ~R�9߮�6�VS�~¯r2�5k�w�����g}�E��L
��1�Dj��2�wr�T-�*��I�2,�X��ܗ}���JЅT;�j˳ݢ�,�b��q3�s%sg7l��o���m����qz�|AuU���٧**���!c��i�����Z�'���f}3>L�+<|z�¢������9l���0�Ϥ�Ekx׼�9�}��S��r��B�X8�U�Gҽm��\���_Py�ݪ��W��u0/�G̏V��j���Ӕ��=���#�b� �N�+q�Ӱ���A��=�7l���Ru��EpՇ3�x��|O��>�V5�M������*W��ə���;����;8'n}
*Ǩ�k)�I�~o=C#2���!~�����X8/_ַ�
	���q�g'��VZ���z�Ly�F-P�Ϲ��1\�f��{�ϩM�XaD1�h~6���y�����{$7[�o`�"�c������n���Ë.S�T9�KZH�o�i�X� ��p^�ñKv�uc���3ߐwc��y�\�9���������y��߽92��xT%~]����sJV+���X�����$���'Nȱ�>�G�E�#���G����=y5���K/�]n���jrul4��]Dg�gkz�6����z9nlͩ$���\%R���RNi��Y69g�˽l��M�n,#���=	��}�L�ɫV��(�Îkr����ϧ�wl�d�z�.tzkeu�VEEϥ��_�o��l�'�,m�ô���1�8��{&�{׾vk��j��;t�g�S�&�o.�M_��R�}�^�X*1a��C��~��?|��*r���]�c��G���{���fm�-
��Q�8f����E����3v�v�ޮ�^{�ág��;zR�s�8�g������8�O�Jn�y|X��W�9p�.�1Y�8޽ʼt����r� Բ���r��UV�V&�7\%�-�.O3��'jn�=D�����u+�'ۼ[2s�u�
���Q}Qw��R��]v�(���{�Sh��h�<�bw�<�J����(��lZx}����7sEٟ%���bLw0.�Y0�]׉ܼ���⪱�#g�1�3�<DGhZ͕*@��%)���Y�;\�C��ņ���ؗL�Ǔ6R	f�3P��.��%��v%ܴ
����X�MN�zY��"��{������kp*Y�3x��[�{���ˮ��Y8�؝�l��$f��mp�ۣ�J?*��ܦ�_���t�}���Z�V��!���aF�ʻݞ�O<d/1�a�Յ�^�G�蝋N�����Z�������&^U��򡑨3�5�o=��|s�]0	-����^��������U)�����|<�'��ߢ�Ƅ׺�#h@U�j/}I�]KE.dTj)w�NdU��+b۟oK�v+Rm���\f�x*s��#�=�>�F��}�̕��D2�G�7/��p��fp>`���/)���ӭ£KiN���uO�J,�؀�qoY��]y\�Cd�q��M^�g�����������=������Q�ﭤJ�ڰ���:�tr�R}��v�;Z��������-��u�G���?n�vX瞼w"�P5�t��5���5�G�^�lÙ�t��M�6�J��mVu���������Օ�I��f��{xέ��z��r�l���#7��Z+���5�}�b���rt�9[(�-�6��*K#%�ol��/�W���r����O���XϪ����k"��#K��.�(�=��D�6��mt���C��c��>�vIJW('�h���Ú����z�|��S5V����\־�Ut��*� X�Y�@+���y<�������k�a�%c��\�I�7M�tT7:(��1�����,�.����jzɚ��uB6䕮)��vV|���u�Q�|�CS�5�t6V�f�Pk;ׂ�k�w�7��2�d�a����\���l�4^��l
��=�VV�"��{�:,kȊS]p�i�����7:��Jۺ5�g����TPB�yL�{G�1#߼�~`��\r�}I?yܲ�U-��\��5�#9��	���c�G*nj,�x����e�����f�&i[SV�?X�O�إ}/)ýf�h���Ț�.�X��~�j��Aކ��sf��)��MnŌ��O����ߥ�|�y�ˡv �c�>�}��o���O�h��f��n�Q;ja17��԰�vǲ���r�U۾5����Ųx�6�|ߗ�F�������v-�cܧ1�%N���5�q�]�̪rE)ҋ� �20���<&a�����V.����U������"|��5=^��!)Y��bq ~�C5��?qaq��^�����MJ��z��2�������nz_j[�c�u�ڢ�^��:q3B��u�M��֣�5�Eq]��0��ij��kcos������/`V�S?~�wOy\���Nkw ���u���T�R"A�����]�yD�"$R�7�&X�Vʺ4ᵭ4:Eˉ�]�bg4��<�m�};K�h�5]�Y�Yج�/U�!�w���Yn+���dwxzn�zJۚ��u�ck���4��z�u���[ȧ&��w��,zJ�:%���r��P���~g�]�>���8*z�<&��{X���{m�	��f`m:f��������3s�S��o��y��ΩgtTz�M����ͯ�s�p_Q�݀�K>i���F0ѭ��P�b�f��F�Y�~��+�չ�Q���#a�x��J�,7�����s�-OLW���%U�OzG�Y��'�)��+��|�}�gHjz�L���󰣎�����Q�}^l������(����i�_�궹OGW��3�Ou�M�^�sL��%��j��-�~2B:��=�~�����Lq]�%?X]頣���/��3|W�>���:�G�`Tr�p4A�����~���6���d��_��9��x����#�.��M���j�Uq���ٓa��M�X���fv�륻���_��r��)hL�Vt�Uq�^���S��i��f@�;��=7��v��1ԴN���I��v^�;���V�M]���G�U�_�&�d/Q�fQ�3ԝ`�F:��)�j�s�����Y�����/����S�L�j�:�$d%�Ug-��ROnx�pY�H��&X���J���TN �w�T�vve�ѝ�xh{cU/R�o�m�EQ�vd��I�i$ۍ�e�,ymbū��k�.�]c��K�C���h�W�?��W�c��0� 9�����]�0V��N� ;�x�{D����*�c+��2?q��(�2�L�U�z����C�Yp��r�A9��S"�T�-�Z�� /4vr�����l�[$9�����*�y�z�O5�)nՓ��[S2���1�ghV���}K���ܻu���[̽'�+j2��M�cK�w�c0�y5��`Yi]j�}�Ƕ��������ま����f4��ɥl��%I�+�]�V�[�"5W������k�=�P�p�s$�ijS����@��b�.D�����|�����H
�Ά]�l�����䢷��S��p9�_Mpz(�ʪ ʝ8�,�9G�R"�Ld϶��ў�xɌ��{�8r����P�6q#��÷5�u��2�*''�ϛ��f�����}]7[�kMn)��U̴Ty����+2�"ż��3�t�\��S��U�k!��~�i|CcXe~��s�����eݥ��ׂd��(b����`�������擙'�B�z�
KY5��hD���ۜwh�����;|{r�l���T����Tw��X����A��-s��(���L`-�0�ڻ�k���j��Gԫ�!Ò���=�mޫV\wt�IG�����Y�=3<g����h��+�YS����}�m=�.�&����Aǳq�b���R�/�D׋�j[������'$l��-�8`�^�b?LYރ<�1ow�3���o~�0C�׳k������!������jyEWMD�L��[��\=}U��q�(��^��9GƲ�����4+���UvQ�S��M�T��;��pƆ�!0j�zƴ�����ո�n��_�Y<t,�~�c�\��;����n���vݩyk6��1��L;�J������Qm�L<�/`�Q ("��K�!�c�G.K�$�5f`i�>��P&�w[����mk�z����7��᱕��Ĵ�|)6q)^9=���Y(Ood�
!W x���L9Z����~�{��%���[D^V���褨�X<���8�^�_<�F��Z^'(����I�<�b�5y���#�|}�r�6'�w�4Z[��3��V}gĺy�_o��d2ݸ�8)���d�}􍣹�ϖ��]&����uN�S1��k��9��>ə�Cz}eY~��[7�ؾx1��`�H�++����Ue�5�Gr���B&����ff<C���\O�� �!K�+�|�,��m�z�):M�u7E�::��$�FJ��w�1�t���ŭTej 3�gfs��s?�=Y��%~��K�,���e<}�Ԍ�����w���ӎ��{��x����QR�UT����Q~��'<�U�,Bۉ��Pea��R�Q*o}�*��ݭ��9�;mV��x*e���u�=i����T>�Rn���%�X���F��V��Ձ����^�����u�,��n��g�Ѯjs�����.6s�vm���g�u<�����W�.r*b���-�����[�ϐ���oxyT��~?�_A�o|>�ū��q2�3�$�YM3��,}��dh��9����<��¹��ܗS��.���g_�G�U��77��Nǽ�W姹e�7k�����Ӿ��+O��B��qc����]w<'%�x>������iz0x,�󯓬���a��\&g77r��v�Jǂ�a���j� ��uʻ�q^�zD�G��lX�������2Y�]�W�ُ�jˁHR ׊��c$cnb�km[��-����S;��Ə�1�^d*�u�e�wEXG�}k�_���E�/;�h}`��<^��IK'�읏l_��åϠA�9:��>fT �帠JL���d���)o@#�EEgJ2_ɓ��m{zÕؕ�e�ݔ��l�mU���d}�or�܄��1t��R������0�x�p��z�X�Q�zhs��d�n,�c:ҵ�3��P}�xtz��-0L����&��_cq���S���p-�efd3q�>dJW�����Y�����h��.��~P肠n�ޛE�7뉻Ќ�,�����D�ыUJ������qn�J�:L�ͧ�5C�M��tq�HT!A3�S�3��js�TJ�9�J'I�N)#:��Ü
���Uv4�Yh�FG��v~Td��0���'��}�*�;ֳZ�����+�����8fph�tYO��ʞ�g��ޣ]��.�@�q�ƪU[�M�{���S�2tI��|I8��Z~��^�֐��{ٚ��G8'ڕ�5� Jr:qd����aK��~�y�7�guRFR����	0q�_��kO{@r�Qjx�9As�:-���v�;��Z��7=k.1�� n����*��{��3���Y�?9����B���d�ǧe�zjvpu�5F}@]��^'J�d�73�޿t��2.W�S�����N���yv�D�?uC�뻖���ٱ��vz��R�\=�XJ�z*sG�<$Ț�u���������Og1Ù򅝬�9��v�
Ys��W��1X_%7~{� WG!^t[�9-*�Vڟ�?�7)?]��t�ゴ�9kVR\�V�}P���ld��U��Τ3��CJ]t�=0�v��gM��炄���f�D	�Mf�`�-�-I��V�����X��Mޣ��8ջwSR8ѱ5�mj��!�ϝ��� HtX�>Q�d��_����U��^¶j��W%muKq23S�i<�m�x,��Z�Zm�T����Ո=���bv1v���q�|�=,.������꽶��\��-�BUC�%�b�!�O�L�.���\j�t����U���#k:�nf��<ijُۓ��$}xSv�zQje>�̵~�@��U��cL����M~���S��*��_�Y���<�Y��&ֽF�nPuR��.��:�������XHf�ܺ�b�TE�Ұ(�Ү���#�{w��`	� ��P�>wi#_�Vm�l�򪪿X����B���lإ9����+M���O���V��-rk'$�x�Nz��V��F�q$�^_*DGg���l��MC'�ŗ+/����Z�����vr�uǯt���(�c�w/w#��G-����7���1�����6@��ܪ��th��]��ž�֩����AS}p1���&��K��԰x.Rm	i<���*��f�[���_���<��ָl�K3,�V���Xb��W%����r���P�ռ_pu7f4b�뢴�W;5��̫��s���q{�Ɗ;��,���R�!8�Cs�t.P?��5*e��0���â0�mqɒ���)R4�o��.�-̅p�US�PW��މ7��y-���α8����9y�L�-�����k ,(U�>Tw�����"fNB��N��.��p̝i<����񛵊�����T���hs��V��s}����D:�,A�T�v��-O�X���g5Ҧ�j�9b�wU��Ic���X���P��H�z�7*�
OU�p<"V-�V�&[t��ɞ���<�y��ޒ�2�&����A�l���;��x�&D+�q"�T�Mq�JDY���˾��+t��<��E��F�g�ɻ��ޮ��4v��[�?%�g��.��Ԅ�uu�p���YV��Mb�e��z�ga�}�˄;���(Ki�L~ǥם����n��g'׽�|\�<�8��6Ŷ�ꊣ�����wb=��)���Π��������Y.7���m�����0lgw)=�õ���P`��ܧ�<��"ז�T�i�RvL��W���p��͐�l��M��i$�(��I6�I&�m��M$�m��m��TK�wo^��<��yX�F��#��ǀ��<Ә�؇f�#�s锴�n�O�I
�m&6�p�T9��_l��ґzS�F�
��[u	zl��'�_Y�u�T�vs�$�twb�#-����0�R+�=1��W_Щ}��]���=p8�J�j}y��vth���߳^w �]�֨�b0mշ�sN�C}�'���څ����O{}���,yF�E}\�:N�="�|)U���%4���U~�����s���Na��~�j��V������5{�h$�m�%��ǫ�/�O�eiu�\�M$�I&٤�S� B(�5��/x��A�5X��o�A�Too�TO�H�c?�|���PS6+}x�����Z����'�Q�>,�ǯٶq�H��`��B��i��TvaVr�[5��v����7i�v�9�ƻ�&V�C�����$����g՚DYs�}9D6y���@���w�AH2����s���s�ܸ�rG�X������M��C~Ƴd|�_��F@�UzLv����ҴJ�h�mb�
~�<��|��Δz����У����^V.o���bi�}�V�;80�8����V+Y*��x��yg�j�#'u�KԀ��V���W��[�4_�;��A�=jزFWՈ�
?(p�4���/�[�Ezv;�c9��ye�i�Mj&�WQ�[P9Mq3Ӑ�?k츍6�^G�7�/.��<�!��A�b����
Z��[#l)��eZ<�I{�fj�P�qW꫼���n�`]V��qk�dMd�z*�P�ƪ��;�b����d�{eqS����m��&���0�>���ٚ�}�PP�k��QZ]��l�6
}H(�W�=Y�y]d�g�A>j�k�/�[��ۙ�P;�|U�u�:�W<��i�0��QZz�������"������������8�ɡK�]�$��(��t�ӒRE!�����n���VO<.څ�/�W3��r}ٜW���7�Q{��f��P��Ļ
Qj��nv���d�o%D�K��zy}�P���p,�7�[��e.ۇۘ���&fpx�bb6�0�^�<\
ܧ�sj�U�s��>�:N?c�(�����gW�sN�C�E�Sט.v���wqF��j�>��77O8��4WA�^b:�PHZ��tpܧ{�)zr<w="ٙ�կ�[qӮ�S=S�9㶛05������ON
�302��_s*tϠL�B���Y�7o����O�<�N�i��㞭���ϴ�ï�c�7_��_:ú��8������d�Uf���z�w�����?����_IG�]R#�}��sv;�u_�hO���k]����"Gy+��<�l�������ߦ������5$�X���N�^۳���j%Lv8;y�$i~���*�l�c��.u�&jZ��)ԥ/w����V<G_׽WW�<���0���!u��kb��B�'�B�26.O�^�ͥ�u5�g��֦�ڊ@��P��Z��1��8y�C_�9?a�|>���ݴ�;`E���3;޾�~H�Z�IPOb����{�O1t�J�<?L�b��悜���a�3A�{�z\����̭Q�qH�k�2���h#A�L����r�<Wv�5��aY��:�
���zd�����g����l��Ҽ�2ߝ�f�ș+�X���<�.+��{�����]�.�G�y#���/���sz�aWz�TV�>
xLg�v�����⨑>w5}�����v��j�O����#@.��g�� ,�Lb���s�<�W��f����+�#ݷ��9s�$������Q?o��C�7ò�`�{0�#ҕ�f���m�S��|�l�̠��^.�%D\f0P��Xm���󙍟�W꼮����;�6n8��n�Gq}=�7s�����U-���V�U���v/���E���>yJK�>��a���E�'0��Xw5:W<��F�Fp������w��ϔy>�����}�������@G%��y�O�D/�<N�����_q�y]»�w+f��F�	�TD@��w�땛����1�{u6�J5>�m�*'��7���)�XY,n����*~�p.�_-��8j'�
G2���>��[w��/@3>7�7a����������w]z1m��W���L��`��n��e���e�X���ٙVh�l;�	ެ���iA�D����]u�ɣ�����cr��)��Y��	O��ʲ�DƉ�znd{&!'$���NJ��1\���Xtl��nv��u��b����0[oR`;y)��[�v�!�VX�Iʘ���}��վ�)A��0J^ӭ7��$��T�vf�9��8��뇑����s�Mp���)�9K���6��LZU��e
�_eo�K�E�j��������/k���\y[�Q���4)�!>�J�~g>(#X����7b��5���{.�0K�U��=�-Έ5��V�p�6z}5�b#fCb�.w_>������7N���GO�|}�q�Sy��|�cuw�R��ܙA�P	�)�[����x4����ת�W�}�����������Ey)�'ͪ<}����u�яH$�+�AY�p�K�c��2i���A�UM�Vz��Q銝��K�ܑ8�g�M���M%ꚏ�eƛ�1�~ȼ�(U�E�`�r3z�ۘ��qs��G=[��%+��c�o,zEǷ�"w0ٞ�^��۽n$d�P�y]\-
@B�Ț�YJ�=�{HmF�����ot�F�{�^.�@� n��2׮{gz3Ϳeب�C��:hsث�4=j_f!����G�V�ue�/V�e�jڂ4P��R�s��NX[A�ו�Rӆ��;��A���q�U#7��ɕ¦ˁ�9J�-�JV��F�!�9V�ʃJ��s���ƚ�v�Z}�uz��D���c�^�����w"4�N����&"���Of,��:���J�$��ՙ����%gp7>��m���w��.��}e�F�*��K��Y��6k�K=+����R�.�m�U�Q��\�~��"�`\�ېё�wu��x�-�����&��_e���uw����K��D��S6|�{Ō���ys7�=^��<��O+g�3�T5�gñ��k�A�e���V���a��^�FL�]Y�x%�E3�w��K�~b�w�qBl�}���':�x�2v���#�֊��n�F��P�;�j��2�2T��/pP@�Vy'��w÷wo�-~Ξ4��^��σ�>^��4�\F�Zin��V]}7|9Q�|x ���v��fٕI�iF�8��2��˳{�m�^{-<>�����޸�Q-��)h��^Q[C�{�C�oS�%zq�������G�*�I��J�c˚�>Ø�R4�MS���xF꿡2��ˤ���w��_Y��^|8 �p�ٺ�2�A�zk\���D�0s�}�s�5Q�8�S nZY1��x'u��o]5�����<VX���3ܰ�k�a�c���u� A��ks#;��-߫)8��ozW-G�ogvܡ�%���\mlneM�0+0�� ��/dN%�L���s����%�ծ9�/,�>m����_f�����׉���wx@س�8�0T��8 �Fi����8nN��^���R�G�j˴�4�ك����2�VX�#�VdnfM���#��K�uu�/��[-�"�zw-C]�ݳ,>x%�١5�1����!��z ?���@�zNI˗]��D��<3�|��'�w�q��4����:�О���s�Z�X)*����>	X9*aM�Ǻ�C0sh�q*���mЙ+pΓ�-�0
=�}_4p��?/qh�-w"~�G�m��g!о7���lZY]�;���5Vn謣��U:��~�B|�Jə>GdO]�',�׼�K�m��˪��tb\v�R+���N����E-�nĵ,C�G�|$󄼏�<�}3Kk�`�|C�;�3��ǆ�O�:n�Mӷf7��ʳ9�.��V��'�ߌ⺉tF�A>�r��e�\wNx(б�ڌ�Cp;%͡޲i`����n슊N�17M��Ԧjn����zi���{s*\9wr31e�wl�Nn�'��'��%u�ֱ��5S�@)z��"���yg2�=�=wC��r�|nr\wdN�2�{�%i�ul��lx��!��]f�,�T�q�&�mzw�݁�޵o�mZ���Ǖ��W�~#�b��RZK�hݚ��ם�Ǡ5Q����n�֓��J�Ci�b��kʔ����,�<yK�YV��$��#c�Rՙ���uo{hF������1`|l.dz4����G�2�{{�G�Pg�B�͎��ݫ�哻��@b3��}��"�����N�_�m���3}S��*��f������u6��8��<g�Z���1�a�:�-��G�E���<��}[C��:h�is�e���|\�5gد˶{���G��V&�ݭ��|1��ε����yt�u�)�=��S�kFv�]���y?���Lk��������;WΘ��8Ǎ\��ҡ�jj{4�<�鋷�mUrWE��}D9�v����Q�"6���s}b�!������� ṢX�́+�s��|� h�㦶��`<s((�3^������W�~�6��6j/��u�K�J�UJ±NFau��Th_O@{,��匪'���~�:���2wl���ӆ_(��,?_�����]�əl��������5wl�Dfuޡ	��{�>���*!uV4}뛳Y ���Y6W���}o�@�Jl���Ӕʁ��Ddt���v�ӝ�N�s>��e�Sr��i���rNְL�ʖt�[[��7|�Z�c;��Ȯ�t�{ے`�3��Z+kgwz�t�ףyf�KF��z��[��r$��M��v5�{�clc4r�&�~��+)6�պoz �>��K�q[�t�wQ6�щYga�,�'���������AGDj�/������Dhf�Rn�=t�>��w�+�NR:E�6+י�|����R4y/�S�VT�p&��omL�=u��u����;��Du<�$��L�3�����kq{U<�,� h�<���P��@�O�T7��������BN�W�h}���KE�����}^�95�Q7s�τa���>���j��t��λD�,`b��>V��/~��S�^���dd����+�z�$v�~Ȭ��W�cFp���0��Q:�z|jmJ'33�~���f��9�������-k��*��=-\��+��H���ľ:�Kv�����Q�w:�Ĥ��)�|�����s��?�¹��b.��*�e@~����������k��T�n2�s�s�Y�h. �^�(v^׺JU�Nӳ'�E��$|�WUK�q�ݬ4uEC��qǓ.o�Ф/���~禎�<���<~�k�Ti�R��_�Q|X�\#�t1� �:yV�z�C�zH�gM�x�]�rpR�tJJ���4cT¡0�}����ь�ТA�c�SV&Q�'�Y��j'w�5:�4G���J&�ޅquִ�p�$^E+��RB�]�'��z�,2�ө�^��=��k*�a��h��+}��M���c�t���ś=�l�-�)��:�5r�rx�wU��L�ه�Fx��
t�c���E���{�wX%�vE�f3:�v�y��uY���v�m��i$˾�n�]S��!��c���F5R�4]�]+��z7Cˮb���4xZ��-
_y��3�����[���~�6���u�#�J[�9����ϷN� )i� ���ܳW��T�H�0e���y��ZNt�yA�}x�:N�T�u�w�����9��MPŀ�zS�h�9ޚ��Տ�T��Km�G���?�����zǰl3�-;i���~L�+���q:�H}1�߮V��ٺ�r�ں�~���r�`�ڻ̋��y�wͭ�G��@֭���Y��μ/�	 ��^�1�8���~�Uw��޺���5ݯ.�U�Y��e�~�M��Ʈ�*��4*�ںrW.�%m�G��Q�!z��,��!'i�u��#��Sⶥ�H�����L?S����v�f�����X螝��3'9T�lu�{I9Z���%*7����1QY���?/UzM�Ǯ�
yҪ�	�yp��#>�؅���ͤs�b��A���c��,y��*��T�}���<�����f�.}b�$9���%�EN� ww��x�pT{/�j�vM���cKWW��>Uc��_{�l�b���X�A��	�-��F�_V�B;�¬J�ۼ���@�|)$��
wu,Jk��7�-�C�Fq뗼�!r�s��i����������mi*����n��������ݍר���)����͈H�YX�vlgq��&������yJ`�/�'��]z�T�[6��xhr��/F�nr��+����%�ϧ�V�������E���N�J��Ә�%���W��L{v��YY��F!Ө�W3��jC�g�mQ�5�u�`�v�Lϖó%S�������9e1��e���^W��D���1� k3�x(�Ϩ���-���j����\q�(U�}�á��*	���O����5�B�<�0kaxv@ �H��H����%�)����R�	��j����yY�#�%.�T�g��gڪ��m�d�*��Wf����`�X׼����1�'��9��m���</xg���M[>���h.g*u��4�Ǯ�.dIŽkf.�$��5nY��<��uc��N��Fq�1q�5�-9t�һO{���^�"��<X�.z�a�;}����[�O:Y.c���[!��˻;��̲��!#'�D�N��)j�RP��n��?T��	�N	؄�����d�ͅ���5��U�uh��|E}�2�ݗ|=�=��"T�.sU��g��<;噽�ZIhQ��tB1Ql�}�y�uVQ��Q���p�M
'u#��-�o�O�.h\-�_�.X��9��u��gMJ��9�w�6ld_1��$Z�q���7��Yݾo��G���s�x�V�ә��
��\��Pn���s������c}��iJG �|�gK�v�dm��QM�b�N�|N��H���ֱ�45�]&�)��/�B�f��s�Ws�p̈>l셝�\�9=��҃·��,I����=c;lr��Ӕ��@�!N� �k���g�b�K�m<��f�h��xPNp�h�뽧�#@��G�<2�ު�z��2�F������#ى�ٰLý�-6e4H�D0v�E����w�E �qaͩ����7���+jBolE�-�PxZx��&G��͡��sw�K���3ۛz��
�u����ޟ�o_�7��WMY�Ee��ó���֒9Q��4�Ѻ��m��q��htA�Z/�ˋeu��"��&���T�t����H2�J�LW- ��T�A6�hCtV]�6�jͫ�_rUo��4�y��i���u!\H�<|��f�Ke1Y��kG\��Qi�{�.�$��p�.�9������V5|���mp��5wbC����t:�0�Ҵ��@�g<eqk��w�&k��%�+�s����2���P2gN���k�[֣7Xa�Vq�z��L�^ʯ�����6��ʕ��,^�e��4B��}����ʒ<o.!��u��<��.n\�2���y�\�9�3��ԁ��}};t�W[hW}�-,����D�uєM�wfuZ6����*k���;��e[s,).���N*?�<-l�E�]�9d�8��,��]7��p:�;y|�(g>�Dv`���@��0;H���:ק���$N��ӋZ.�zdW/���ٵ�e�����l�L�Q��p�GN���Z�z\n����������eo`8���S���ha�������Iں'k?M}˽d�����g��t�,�8������)��{����Ls�\b[��akl�����E��8i��c@L�\͛�nR�!(K��N��%����Lp�r�EgW��6U!W�4�_oV��YXm��R�n�&n�+ö������0�"�n��3T��,*�͖ �7ګ��!��v&�r'J�eb쬅�5�������0<Dp �!��b�}J�>��B�e8Y�𦂝����`@�nudI=�O�w�����(J1���R�}�>�ɾ ���:��]�b 3�Kq�VtF���<���{�m��G�r��kG�=��W�
�s9h���bcޝ�7�.����-��{�j�b[���ג�n3n�}�*��,km ��d��e)�m�p֘�X���gp;7����y��
���n��aX����}���<����|�+�<2L��J�w,yDl�OQJa�����/w��V��0m̆���G���Ӷ�/Z��=��[^���]�:���×��*�H��@�+l���|��Кt����:��c��^��ي��6�b�p;�I ��*n}�#��$O�hɛW�����o�c���z��u�wʺt��#=����Ykۊ�/�w��߻i����}�'TK��C����r�H\�
N��Me�;e��l��,������y�N|V�V��߃9�l�sǣ�*E�u��o�AY�=EZ�1�=rJ����Ś�H���یL�7�O@\Ʒ����q8G%!Q�"�n��j��3zj���z^q�x��iھ�}��uὁ�'��â]~Pp��>=�%��6�E��c9�����
���6;2���]��6����g�O���]���u�p�(�T�.�C��G�2�u��$����կz�s�=㑇���\2JRp��O��z�3���\ˉ��
�(�R1!�R���ӛM@8a��^����h�nQ�Ҟz{٬xz�wf���y����p��>j:�3¼�:��u(vLtL���{d�/	��X�]��{�0H'�)��KY�Z`���!ݧ*j'��gf�X���&[���]�Y���si��j8w�_2�m*�{^Rp(�f�r�+/5�`(lʹ�j]|�,
����^��F��D^�W�����9�[����(�.j{�rg��4���σ95#z�s}��$��S�]3x��V�Ǚ������ױ�0i�0�mTS�@��j�O'3#w��P�Z8�M���]��ќ ���>rn�������I2��v��*ܫ�&7UL�zv��c�a�W���O��׮-�9qԻ<����
XR��'$�؛���l��7$���ٞ�����`"|N֞�:�Mm�g�w��Ou!��v+���!�����޶��<^*jª�����M�q�*�;��#��GЛ֏#�>�4�/�@�7|8��ڷ:������i�E{��j��)�W�MG�l�+S�Ε�ˣ��DwX�3f�����J�{��x(lӚ��(ɨ8���8N��ʋ+n��	���z��g~�B(�ř��k����v�z�;3~�^G�ym���^��ݿ��{fK�x� ��y�Ӝ{������:{ء����C\�o�q��
��s����o��v�t�f]M}�,���t��%���o�x���ޝ���[����f�n��s���4"��������-��_d���O���N��E�o"���^��א:�y"�3Z}�  �3�
����]-�m��m��ml�����Y�Q�ߴ�h�/!&�fRr��{���r���R���fm����9�OA>7��ƣ��T�o��vhC���/G�&��my���(;7��ϩ|>Y|OI��+���Y�\e;�#��q��,-y5�՟�Ȓ��ߋ����o���v�ݺ��Sd�0�pz�#ަ��#�(�e�WRW�͙�Y�>;��Yܕ(��i]8����Dzszz��������^u���*�OW�(���sʺ	�U�G,×�#۾��<�t5-�t���6�羊^Nb��܁Lb����.U�*�ԥ����1-_v4{͝�c3�sY2gm����S;>u���j4�Xq����ƚ�y����Zz�I��T�AuC3�[�+�����i�g��Ѱ�Q쪄o��b��f��$��'t�6�y���،�������՘B���}vg&��#�{��ѡ8
�f����>����^SRL攠�=~WBg�TB8Z���iS8�=���UR�3�pf�f���w59�������fٿl���1t��n̜��Y�;�m�j���G�E��M�`�'���-�ג�a���D���n��<��������Dl��Аy03�����O:/{��rQW�v��bBm�*j�[�ʕ"�9��h��E���+�� �H����3���H��w"��E+]ǯ�u�z�u���{U��}38	�Ż�ok��=,s����Z��R����x�gR]P�����������uwbA�'/�\��o�Kl���<��//�/d��L��W��b^�| "��1e�~%hͱ���[=9Wn�Tw��-��uS��ѓ~� F�:�yk��Uf�-	@��ҽ���n�]�%�ד��:g
�P}�z��l���N�#�9�o��=~�Y��ʲ\��5����]s�^D����3Z���fV>�Ճ2�y��ozj]FV�+�!�}.�sչ�����sD(�{qx��ǟ��I�,^d��KDH��C'���x���M�	�>�����}Z:���	��y�S�p<�Q�S;.UѳJ̗������'x�K��U�kAF��Ӝ�c��I�%�	f�;�_�f$5v5�g���J��@�h �z�2-j��u��.�{������o�����<Vj��K�Vp6�Fُ��y�]�<Wx%C���/����<����Y�`�Q?��V:,p[v(|��V��^j�N?y�<�B��nƌ����ܞ�fe}ӥ���@D<�,(4�͋jDbˣd&��+Y�X�R�()%��ݙ_����ƈ<9���e((<��_��v|{�O�%Oü�����/^�m`l�y�70�*t��_h�Ù���t��7
3����A/�:��}T�N�,aZ��v��O���_�;4^v�e�bǧU>�qFR��,����8Gח��EsO��2�D�ia�Tȭ��]��1^�;��P��Ԫ�U<��z�]S�%�����La��.�x����x�4����w	�����Uŉ\\V�M���P�^���g���{0W�,��j�aܯfEW`}]�n��W%@���i�\�3�z�?��=��S~��V��wN��@�6j�R��g��z�%�vv2}H�9�t����B�.�w�h]��g���os�G*�d�C>��i�I��^-G<���b,W��R��5w��Z�쇻�^�ו�F��d�z���x���^(��e�<������9J�;z��ޘ���P�L�њix�ʵ��u�?#_{�-�z^���GjW��k�`fU	C}��U	�U�;��k'6d���΅t99K{3�ljel	C�L�̨��6*�}ʣ%I�4��ďd⵬���[��.��X�!�@5��E�@�����(�nM�+ιp�E���^�}������)m�iw7ֻ��1�j�Ke�X��얷ɵ��ε�;k�Eݪ�=s�zVD���R��R���]<���-���Y�G�\X�;v��d���k�g��c~�o5ioɰ̬u�+���2z��)���}n\���߽3ƙSb^��[������W�ƣQk�÷�:Y墛^�9����Qt/잏���b�~��hM�sK�e���l�sm������Wo��#��X���H�Rn$�u�&^���V�]h!�e�n�������U���~gl�mUi4�qS��wt��d�'ϕe�;���r�����(˿)W����Dx�>�2)i9>3Qo/��5��Jh0�����9t�|z���#ez�ڎU����ޮ���+�g�<hc���"��E�oCZ��𾮷�Fj�sDg*�G��ُLSW�o�:��U�
Hzf�l�XN�Yk�p�묙�9{ջ�k�-�OWl�0�a���QW
O��Nn�+�kl��~Gg�/��@�b���i���}^qg�j��2ۋ�(}��_ͯn�ʬr��Л��{��t1+�W%+p����\V�V�����L��p^�ك�HQ�E��(թ���c�C롢���"CZ\�s������@���׽*��fgj�$Ƃ|6g��`�_�4�)�ڒU��R�\'u��*�&�4{1d]8.�����ڥ�*@_���.�Y���כ8�J+V��F���	�rU-x��v�3�Ǉ1k3��ysm$�m��S!8iWXڙ7w��e�V��gt�ge��<��}�Dv�yƪ��`2�IV��ڧ��{ϵ�=�����l�����_��6"�Bg���JX��q|SRv�H�^%/L�{�Ź,^�]�`�N�������;�6��6jj/D�`=����x�]��Tu�RH��n!�G�����0[�]���\�#z���o9�
��t�f�7��4�D��vL�������w˲����4�k�C;ש���84:��-ʆ,�U>ڛAX��J��٬����U�!A�L�k=P죈v��_{jソeD+Jɽ̕�Z�g�����<1�_�x⪡;RU�s�F�:��.=�<�y��C�2\'t�����q�Y<�_Oޞ����ZV��ԉ��Z;��d��b�|}J��ՐeN�5��gA�鼒-��xW����Cկʐ�_������_
~�ִ��[5�ߝ/h���>���9+�%� ����N�O��B��(m6+U��zuB��fs��t�Tʍ�5�[[n+���-{�{��.���H�/���߯,�nv�k����Z8Z��;P,+�(�=�{� �ٔ2'*p�n�Tp�UKv�Is�G����6�G�Ь�+k��&\��c��C�69d�;��gvv~������ ����#�ќok�rCp�v�&�t�M�y�E�Ʋ��5�Vō�u�}�'nP3�[����͘��.�Ȭ1�����]���нS�+�������g�jS��d{�b{w$b�,�U�>N��;�ϹeB[��N���q~��輛���`�Vc��FpN�;w�ݵ�����s��v���r�_�Wx�#�*��5h�u��XQ�t�V��,�N�������=2�:��9�9�z��=o�M��t�T��b���.�)߉�{���+�~���xEQ��_v^.՝�$�8ϔ�Q]b��g&:Y.��-�R��a��Dۺɖj��Y�gO
�:B�q��_a�{R�
^�c{���s^g�U���-Iw\*ܿ�Yҁ�q��3QZ9@����=��)���K�u�_��L�9�+�V�����FF�^꽿��R��N�к�\��.Ѿ'/~Z̸G��y��o��b�ֺkU���ˮ냈���.�)o�T�ހB�?xʭױ4�
�8�����;d��K�[��A��i.d�[��=�i�2�T	�P��tF��s�Uv1�n�0�,+
Q����P�J�~6{&�������5
u6T�s��+�r���Ȇn���GSp�Q�e�C���2��K� G���֨:P{2�Q&����%�a*�2�-ҙe_a�
`\�S��ݰ^�|Aǟ�-�5z��p���U"�
vY���?7�[*��m��O�j��~�gڹE#�{%�M_W�%׽��<k�P���G�.�|��ƻ�olV�<������s�[J����_r1ٵ4���|���76n��.4�Z!�5]K��d�N�M�9�&���"p�>7�=G\�m�=���yW��X���@���zL���&M��t��@Ǽ��W}�U�ݝۿb��TQ�����.��L|��'����U���ҳ�� ��F�}�t�����Q�^p�k�;��=��V�F�`U[%:[�'=�����՞f��=�X��gEl�w��o��7�ٳC7�)A�~�U�lJO2�V���٣��B���%quk�5M=R��mˑ�]�p3v2(�2�d�u�q�=s��t�_����y݊���'�uiAo��W�Ko�Y�^p��콁-/����I��P6�ck�HB�I���7���;����F+�!,��2gv҃�	�� 4��{Y0Uӛ�=Bb�7^��f��.�{�z��Eݻ�&]�˼b���E�<�u'������_Er�ݭO�Z�/V*X��-��*��Q�(Aۃ��"��k��N�m�@�nڡ���ZIsA-�"ﭙO`��+�}���g��)X�&U���[�'zňk.�-0X�(��d>��E��<�z���N��=�=�>&��e:���"��-�������Ra5�K��s�9��+����͉ȍ(p"7ʔ�4�|\fg�뿛��9rĿ��t1{4�L��%{69lWA�$���sc��S�>'a^�(�Ntw�K����&ҡg�֋�
��N�f�x��`Nm^�����D��)V���e�af��}N�,B�G����K������ǳ����?9N.�H���}�\����f�\ݣ�gz=�L6�Zz�l��N�J��A��?���+k���]�h.�P/�T�s��T��;vk̂r]O�����^��u���k��O�}�����o�vYk���J�*��	"q�@Tba���p�*M��;=3������8��M�"��yC}�8v������S��p_U�I��"����>M{���/`*E v���l֓��U���:����%N׹J��'Ӫ�����V�9��Q3����M�6��@���gGԓ|���´o_G��j�����.w�g��;�g��3��wK��n�k��F�6�Wr���Q��05yz����u��i;�w,/d��Ŵ�E�k>L�=�.f�2l���重+�{�pIљ��-������2xaY�W�C�B�2���n����&bkTPƫl�\<jq�:X�,�����ۆ���h����<[�;�Gd�EP����@��N��5���?f�m��~�H��N�3�v�[��)�<
n�jR�E��,�Gyn�&G��̻t��p��=�<�j녁�I*Z����I�LBuΔM�軲���rI��2�U��V��Hf~��_���X5��~�j�QM��ީ��5Wq��U�u,�lx��m~d^�N�(љU�ބMB�4ع�g��zj)�ݲ�V �dDd�=SN��F��YӠ�)��	��P]w�bߕ{�t�a\�vY�ʵsV��;\z�oϚ�F��Ó�c���b�kDS��.�Ȃ�H|�O%�����4ђe���#Cjf@R/xʾX*ܾ궒�6�:����V��;�E�}.�LS]Y�Ι����cw�Z_M�,���/M�k�[L#�8b��m����o�O�w(Dtę1�޾��$�aL��q�Ԇ�����y�.� ��BOx�{`>k.��y�v̒
rzש�ڲ��NκF��|&6������6�� �+�wcN� �dV���4+�]�e�CfiF��d[�4��v&��pZǶn�Y�2·�	�"��t�h�V^;���.ٻ���H��v��Ѧ��Q�4��.�;Gf��4d�ԣ�@Nn�V!v4s]�n��Μ/��Sy�)�����<���
�}���L6��U��mf�nA�=�f�R�^NO�S���kb�KU�����Ӿ�=���ux.����2n�]���T�Q�[�7l:,�6F����'��n�S�\�W9Ϸ|������B�/�-�(ۏcŰ>|okwŕ��-hſ���uv��հ&�l=65�;t��8d�P�L�0��]���L������4D~��sp3��Mg*.����28��K��~��L����:��Z�Ȏ�Ɛ�nb�B�����oMue.V�m���9bWV`��nR�OW '��_eB��(.1e1l�V��GЕ�M����rK�*��Y���L�+(۸-,���emF�e�1���R������xxY�]��nG�zR�+��1���Ԩ���=�6�m��m$�m��m��I2[I��I&�m��m��m��m��m��F1��n�L:#{k���|�]/ �.B(��lu/���M'�3&i��ݬ��ã�I&�͸6�$-�����@Z��3)mGʋ��Y�5��y�إ�\Ntz��D5�:)7)Z2a���i��@/q[�ac�wAl��.��8}xs_x?&=.���4�5�K�u��M�ڲ�0�ִ�F�.�Qr;[Ƿ�ƑM�]�b.�]��p�$nz儍 ���U�<�E๺�g���R���>9{ؔ����u��A|��t��Vv�;�%�2��I�v�S��.�u�𒕶�I��)�C7��sO~�&T�}���ٽ��v��ݖX��$p������v!����8�^�����⼫�F��t��l�LN<�+�ig�.�%J��.OL�V�]��ʦ�t5km�Nzw�6�F^������1�^9v���v��� �7�?"8F���|���A/����}6��7}�IQ�Ϗ��1�Y�O���5��wN㍵�}�q��f����n)�mzm�F���S�i�ګ3J�GlM�L�Em�Cq�Pn���*s�A��-]Y\��+2+�J9��x�7�
�D��|�mع����q<�Ӈ%ܷ��"��;��b�m�~�4����~K������k&-O+�A?-��9��鑁eXDl��z�E���V��{& ˥�C����P�W�mb�[ѐ�%:�V������j|)9���� �+�їS\�!�@�>�R�d��T��;��Z��*�TM�q����'�>��vr�d���!�7�^�<�oO�N\�]�ˢ��@����������������_���j��}KŘ�\vEY,��5�h:�~���ՙ�>�c0����l̆�[V�����c\�Vn�x�3�Tx������t�&���}�*Ίb���S� �)r�g+}��>#mȑ�!W���?y���au�;m*<IӜ�{���'��/7���+w�i���_`�{'���w~�]B'��P��(�j}
{ٞs��=a�FݸW���c�deu*����ogvv�L���59�1��J�<��7C.��[v���N�iD#�բ�iۉ�
��[��F����k�|}>ӚQJ�i>�-5��٥^�cweĝ����C�_s�Ac�f�9�'�ǁ�>��p}�R�sވ/"�B�=��f�J*,��*X��N�j�`���U����594�~>�w���L�/�+qЯ���^�-�C�\l�1���s���@�*2�BY�E�:=�1���G��*��[�{�E��ʪ����v/c�v�i����_��^|��	Υޅ!��o޵b�t���r�u+�{-�G8��
y^A�YG��ω�'�1�����T�Y����J]lu����R~ꛁ��e`/f��qymW�H���0��^�^��zf1{��H�X6L�ԩ�.��4Idf\��+h�^u��~�%ܔ�@��nq�G��o@�%�Y�#�~L�3w	�ϔ��Q{]��d=�,�����q��.ĸ͑��Yˀ3^�V(�@��cyы7�4;��4�������3��5�$�ۥg�Ʈ�\[�EG�z�4uݤ��]�fG��pxm
H$F*�+?-�	j����t���Y
�X�p\�*�����4�3=��)K]�� ̊�"�z\(�I>(��i�~~ѳ'ᑳE+'�_M��Q���{PvnJp���������/�k�B��9EfR�*e�xM���Ťg�t�ҽ��n�r7��:��y��ϵX����?,�9�V���s���.��b1p�A]��HIKE[��+[rQz�%�������ݺo�
�p���]����Nz?��1�����܅҇�X7*����I�;��{�:47ca{Ӛ. ��U[!�nϑ����/(zR�ˇ^�lGp��3�މ&�S�a�Ǒ��/WDҙ¨��KԠTG{�Bs]
4K��Ѓ(��L<�~gX��$��v���ϤeV4��I�⏨�yB
�dG�1�A�:�x�����!I���n�Hc�y���i����=9���su�W���B�51�~�9�j����d��*p֌��gUQ���o��s��+��p��\_��)�� ���<󍰞�@u]��߿It�b�`ٵg�F}�6ڟ�X�%��v���q�C{v�����v��K���4J��7�^�P�i�2���q��Iov�̧�fbG]l�|�-���**�7�+�L�� c�� �|�{�^+G$q��NY�mԵ�	t0�%�b]��V��+��I�6W����y��W��O!��3'/Ɛ��$�g]���l�:���^��	^=�.�q�+2��`����=��' w^v�Y/�J�v������9V�|���>w��߮��F/x/Y���M`eB�\w��~�Y7L��|KR�bP|,�<73״�s�/���Kcv�����e���_��}��j�Z0s�V��eý%��.��檅�f���N�3Oݪ�!*�ִ�O��λ��!��N�_?(��+U��v�e������J$�j>���ۍ��ի"\���Z'P�f�m|Z�����=k"��Qvr�I}�O7��|�F�RUGw+a��&UG���g�s�ޏE�W>���`/H����F7�V�8ϣO����"ӷb|2��"��7�'`�ّ5�%�xd]^i;���̮�����1�Hz�>�݉�}S4L�-f%��<�>�j����_��[W��ms��A5����=����9�����5N��S���m;�6c{ߍ`��˞!l�'A`
]0x�+nj%�x!�}>�����V����q���3�C���W�<:����&�@�j���,?�躷�vLZy���O5�A�I�)�F=�XB���O=�OG���ᛔ��������%�P����N�X$x]�&��Lx�I-m��s!�]R��G�9�K��}j�c��n�aY-���u�t])�Y����:���dF�!t���A@�.D����E;Y�g�!G�}�V�K��|���9�׵��Zhɢ�Ti�3*���z�;+��L�vЌg�y�{�οR���p�� ڛ�)��^��; ^U����V;��t|�)�v6�����:�e�����K{���
�Өt�umwЦ�ֱU�����;��q~|&��#Üı3�+�Bx����iUװ��sή����u�U1�2�I���S��բF+ү���洉Ri����w�^V�3#d��w����.�(�H����J
����]F�g�c�X8#�{��e�����Kϱ��q.��y�C��^���77�p����'>2��
�|�����==���1�^� ;|�>��������<K���qn:�b�2xV�e�7��/"����YT�d5�~5�:�f�ų
��E帤�7.��.��T\��h�;.9U�f������{	�p���`�˝��"�7�o�����-.�=\�m����,�kh�֜����Feˋ�`{�X�
_^�!���wo�?\����Xc�l��c{��'���YO3n���%��=�"�gN�	��Q���4�:��ɤݞ�wُ�b��O��Yk!޲6T9����.3�*��^x�3ֶ�"
ww���]w�7/�ϰ���X�|V�_�u��i�A�$]eV��1����X�x&"�^{W�p*c���7f}�S��}�6��)ڪ�^a�}�2�K:�xL�}���TK��T�K���6����z�K��u�]/IQw5�����K��-�=>�K*�p���1ӕT;��!OЩ����v$,����t�T�>��`�;=ܯ�e ]>ˉ� �I�����x6g6��4��וӍeAŴ��M�n2c��Ҷ[���/��	�y
��Ԑï�:�L,^�W�ς2�^yڣ=�ǜ"�h�R��Ø�=��z�辸�Pz�	=�B�A�z����aMD��=�7�sx>�ߛ���h/��mo3�K���U}&�k׳G�Y����4�i���U��S}�����{`U=�s;�M�{HX���^F�_�J������	�w���]�Js����K��٭��Fr\�t�X)Z��"�&j��Y6��Y�d}w�gSxn�v�`�R����T(��a^���~��lq$&�������5ݛZQ��GFL�ג���1xtl�Y����V�}-��R9*���R1j��P~�\�y�V-|�mv�q�X�w	�#��z}��Y��JW�����8�,�zAR�ý��q��=���io��M�oB�[��˗��ݹ0�x����9�<iI��Vr=��3�:kb�[�����3E��s��<����=�m�r�p Fk1)�m�B+dKz�����P�3�-���3�l�3����!�Ϻ�����Jh+ۀ뀍1����ߕ�̎xe�-4Q�O	�߆����%�>�5T�k�I�koy*D��vqW��������#��碼���w�������C4�Hͱ3��FFj̥d��A�i�ʜ�Q�j�+*�Z댕&̇�Wfdt��3�f����>��;
jGk_��VF���܀�3���P;S��qch}���
�n*11��*��R�H}i�sYh8xa��vC�����/�1dr|"�~���[N|-���̷�/���|^)�~c��nvH=�W�v�eM紌��Rk�:οIw�F<Q,�
�W|^����~�޼b�m`J��N�2 �q��+)��* In�cF5y���8�ו�PʣG@��(oqTJ��:��:�C�wE��?�hN�I�)z�M�%>�]�d�{ޙ-i����HH�͏�ue�i��m��?g*�F�a��n^��6/�~��w���o���w��Ϧ��0A��ⱪGȫ�# �t�Ƥ�1%�B��ynbʏe$�iD)o��	��77�cs�lGwOn̯H/�kblO��&`#�׊��ga�~�+˫��,�G�<�ߢ�NY�k��Z��d�@�'|�Vⓗ����Z/,·"��#���8� {"��/| �#�X&�R���!5�!?7u&zU�#�R�3=���拇�tX���՝�s{fBw*���aK�qW�םBU�4���l�8܁��(r�/P�-��Un��[w >�k8����U[M����*�����W{�ٿ�J�
�>����_G�P�"$�~�ޤ)�Yى�y��ntts���i*�Fw��b��i^ߺ���f�|��
�щF�s���9XQ�����͉3��߅C�v��̠PYF�1��rl�gx�:�cv����Ҿ⟺�ؾ�1ՙxd|�91[��>Kn*�/#v��DNyU,��53ֆ��cte��YM���ٞ�ߟ�F����yb�c�\T�65ѧ>�����s�]��cg���V�b=���t��t�T)Eb�	� ����.z�C���ۺ(����9@�÷-��s(��:x�'��w��$;:�s8'�ï�x{�U{�sM��-$�nJ���͛�T"����z����At��o&���C�-O�N����?�s�g��/��}���.�X�!E\��b�&Yzw[�o]9���h]�w��ly�j۩0'�2���גx��(%�,چ&��;��З���"��	����������W�*+:��K;�!йS�%��=���6_���N�3�ƃ�����7�#KB5{gO�Q��/ƍ���fD��B�Y5�@�$Is��ɸ̀��}��AH�g����l�w۷f��Ǜ�u��I�$}>�����(�3��G��l�O��,�-�GC5��)��.ǵ��^4�z7؄QJ�=C}W���[HE��8v���k%��w��k��u}ǆ�b.`!��o���*�������Ι���Fڜ�J�d.�&qL{��@�qN5>�����\69��Q��N�rsr@{�;&��eq�C9��e���i���M�|X�J�?�7���}��|4������U�I^����/޼���/i{�jQ��H��|:�z�P��k�){=���Ǩ*3����C����9�J�]/�9|�,���$�
��]�G���XY����\1K�� �����!��m;����7��Q[�i�o�FZ�����v�vyʒE#e�p56������
��~�)&��j��E��=V�^rkUFZ8�X<���OU�b��Ԕ�`���3�>ʖ���JOXݽ�GQ�<:}~S¥z�7G��#m�;f�Pn�U9kr�N�F"r��P&�,B���6D�յa�*���U����
�K���y�mg�_v����:Ǵ�+U�ԅW����]�?fc����+��J,5�>�NN�FD�;s�8�"Ϧ����sft?zg��6�!F�S
��U��sm�L{	�3ڻ�� ��)����?N�~�j!��l��|n2��Й����4��o:��x�C/������Ǯo���w�ӛi��]7.fPбΡ2�A�׷Us¹H~�̹=�ժ{i�Xk�US�UX��޼���¿y��J��LyߍTu�G49��	nmJ���)ZOam��X�Ίnݜ-`7Lb��lύ��y�����۝6��LY�����'P�:�a���t%zb�l��EV�+/�0m�AȞ����~=~�F�ִДk@�7��)٬t���T^(�sjVb��=����S��)L���DNҭ��c˨
d;W�u!<��ѻ���7ܺ7/
81=�gl�q��y|�t���r�Δ�9f$dT��~���
���%���0��R�+���;�i⛗�]�Egj��?f���E�,��Ʌ���Y�z��D����;��O�`j<5fF�R����b�56ۻ��$� �N�KCq�_Z�Bv�����v��W\*~э�$90�[�Q~)�t����ţ�WJ+��yT�6խ���8�;Ǳ�z�/5) �=;�hgi�Qs�r�w�x���} Z����t�ޣ8�to�;��=�vzi!�v\Wo%1I����8��j�U�;��2�M�E*WAg@7:���:�l�c��sl��0�A�ضʷ�l�wK���O� 1��s�s��W���E�겤q�{κ;PKR*�U���<�+pj��y�t޻�G�s�0E��˱�m�:S"<mrpY/��Ƴr�T��;��� kC:��$�Y}vv�N$v$z�k��T�q��Fd:b�X�ep�*qACy7
�y���5��M[�yPe��]�P�����sǤ#x�!v�fJ��<yB�]��HT�j�#���T@��:�]���P��8��w���[�a��h��2��|ea�<Tz�Z�2�L�5?��v^7�T�$Ɣ���Ai#��Vue����v[�[(�a�W��L���^ҵ<m��0.�hx5pN:ƟWIS����UKūi�U��ӻ�Rj�����޻J���֙Y�5�K����_S
v�\�}�hQN��4�miIY&����oO�l1�?L���e�:�`U}VN�h�˓/c[���P�%˱q��'s�x�n�e{xB�Z�gBC����:��s�]9Y�S���wK � W)�ݣ"����r0�4Np�~vhnC�2?Q��#�B�ZӭˮX�]q�_)e��46���4N]{� �t��,T���'Gַmïg1�}k���H�7�:]e�)���$�v�;�v,���j
ة��ek����ѥg�4:���i��pĸMu,x�5�Nќlf'���vm�J�7{+�dwZ-f�%B�1�[���<�I��\�q�8�B��O�/݄�����[{��{J����
�+�*۲����+Okac� )ta�B�Q�.�f5y�N������mhД}[���U��Ș|#յ��yY�l��1U�D���opv/�R����gR�(oN��(d\���P)Q���P��j�H��TI�� ��=�)�#�zNd���_^3N��&��4S�:�����Z�ٚ�^B��u6�I5ur.B5�yàb9�ƥxd+{^eJ���e�A晐��g_Y��:���CY�ḹ�vF��R��Z��B-	��V$��M4��ܕtѲr��|>��"�ʋ��U&f�nz6c���+/��m��}�ȼ�}����_KNx%n<���T �57��_�o�˸;ai�>�o[/ ��y_E�r�;'��w�Aqu�cg
V�b�jQ���D�_��h$��pW��O	�UCeƹY8dXn]���fcE~c.���	W���&6�wEN3�F�Z\�l��F-�"�ozjf��j��:���ば�]�P��{�����J�OzzN�� oWs�^�G[��ʭQ;�h�����՜��ʚ��bg{|����P�V�gm�`Z��\����۩�~���H�V�>�{Ϟɷ��� _��3׬1왺��}�1�;�;�;��W���zc��t�+���=���Я^N{8�';3��':O
�ԯ��̂�B�ک���Rڞ�u}캽��w�	J 0��K�ۙ�C��3�2�z���V*��K�gf���UK��O�8��V��qw�&�v�T��!�6���,og],���JJ^��OK�u59�c���g�f�E�{����ï2lg�A�8���h���[�>�~��Gz��ߓv/���6Y*����r>�����,s�{~��#��'�Pl��ǣ#t�W	���hv�tL����qk?\����o8C�){YY����� ظ`n�P�:���R�uh�O�)���A^�8��|b�1���خ�{;�1돭U�<��'dW�Ū����p�@�T	q�5�'�	��O�rݵu�ʉx+�?\=���Ф]�J\�<#r�7y]e�ز(�C�Ji�ۇ��_��5qG�)��X�w]Ñ�$J|U�+=,I�P����:T�N*�xqt���6ĸ�QG'C��������:�;��^����O�������{�+*���\����Z�9���ԧo���Y��w�}�9�]�O��6��e
�����0�O�2��%{|^#Kx�|�/�<��n�y��1�Z��\�;�G�o�y/�3'�/g�8���+� a7%�c˖Bn��$^/���1�|ǝ�9Qީ�=��,ӽ�yw���8�x�M@����[o���ESֲD{�Jq7<5�%���{���L_<�P�9dv�w������UH³�`�Def��J�º�+Qt�|{�!��ڦ��>/�>��=�ٍ�T��Cl&��"�{�{N����JEd�V�����v�ͷ�an�m�l��{���� ����v;xN8ӣ~��r�5���b�f�^(m�`���|��B��1�M�B�Ӛ�����D�V9��5w:\��,�!գ$_Q��j��*ak�w��C��D�ۏ�2��ь�[@�sm��mff��)~��$����b:9e�Pǃ��E|y:r����f��p�w�ɾ�ؑ�0�gNJ�f������l���W;8���g������_Z�x+7���nK�����n����)�]˥��:\�q��y�i}�����\����^5�1������[���%
�an_�r/G/[ �50��1/7y���vF�3��ꗅ�.����Y;��wHɁ,�t,�>�'/$՟{ z�����0.�(���U�gn�(~tD�MA���徾W�zȿV�q��Ƴg}��K��gf��{�ȯL�1"W��>*�\:2�^�Z���8�O��=H�E���%5 σ+pob�ך}vm�z�o��f��*u��p�M���5v?">t<��H�q��*�C}P�[��o��+�7�lds^jq殍��m�1!y�L�HP�#���E�W�$+�:*:l��en��߯�<���{�,�['`[�h��z���p�j��ǯ3�%���=�)z���`�+3;�z)
���qn���Tx7�bp��ɥq�ᏰY��\ɞ�#&��\��i]���(�u�q�L�6�b�Q���TE���UwNU&����sWy��o�櫣�.�u��8t�F��x�J���5�����m͉��b�ݱ�9ݕ�8��X�8`>3ܰ=���ms�������o0�;<k��;�/L��v	"50fp��H����^������[�+-8.�b�m��ߺ����c���PMt3�e9,='|wo���=�jno�Ԫ3wX�ϱ�|�g�u3�ĸD������X���C}u�^X�ns�֞��6��\V�_�70�,�sO�9����O��p2���b�`��F�=��y=�%����D�t�}WV=/yS���۹�5�zرܩŪ�N�jȍ���7�Y�	<�U���{4�V`�n�Q�:-��mݥb&q*�4����2�n�s���Ld�y�ЍH�!�����+�G��t���^�BCK��U?M ����j+jP��}ìmJE+���e\�c/V�z���^Ǖԍ��`��ӓ��-,�n�+
3��k�vT�Юk��;���vй�.�3������ƞ��
Q�6�˃�B�åuo��{8Y�߾(���!lS�*���zឳT\�HC�%᎛� ���4V;_ZXZ��~o�V@op�|߇A���[�TW��P8�R��YӂJ��eZ4?(H���u�j¨�:�PL���3%��b��u�$�6��ς+�T��t��`7����vlY7m�#�����t���h2}���Z|n��Y���mIn֝/�EmQ�� �w�\Y]��aٻچ�L�9aeX��I���/�M�=Y�iQ��c�$%]G}�+�_�Dh��q{��x�j�v&-��P�j�fxIgԒ]0�gc�ܭ	�r+��A	NnW��xk~{b�����ä��)��4��C��[Ϣ V�Y�a=��(����+A��Lzk��R��r������w�����`Ƀ���k��E��N'�t���X��f������큲eJ+�s(3ҍ:O��bz�����rE�*��]M9�w�\;6'Lb���~�̟�!{Q�p��9�954Κ�l���X]R�]fx�}�f����z}v%d��e�d�������XQ��N�F�3� -�\D���' ���]vo''�m�[�ge�F�C�8�!��	�ʊ��!{�"��x���(v��K!�9�j�x����-5Kk�\wo{�zĿk��,Ⓕ�Vp��:����Kykɣ��'y�ɷ��X`N�9�W�݁[��=��Ǵ�j�nˋ�=����ϲ�t�b)Ϩ��؋V� 髇�=���^1�Y�n��&̺&�tX7*vV�ױ�zA�5
���
d!.���Y[��	��D��܈ԭԅ�`��U�V���d�Ҧc�K2��7܌"���f�1�3���+ms���S�XC��Y�3�a5L���1d.�9[��p���=�t��Z����Օ��{���p�~M}�Vjy2��f�7kI�׷�i�Z�UqR}uBeg��7��x��w�����my*9��W�
�/�nD76=�ӛ���6���G��Zׇ5z1L��S�y�h��r���� oC7w����M�^�{��d,�Ι��8�ާ#!����]V����.����M�T^FG��N�3�����3�ƫ�ҁ��g�:gG�#t�ǳO�{�+�R3O�A�N���f(��L�f�eځ��K1�`��+��.m����������ό�4���>���\�`�:954Ö��e�=V&TdVӖ#�(�<�e�ݲ��S��U��"﯃zHb5K�]�L��S֨�(M;�����c�mN�SsO)c���g�w�k뫿������.T��������Zg_X��`�^�{���A8���8���$*t1~w�z�IU&��B޻>6؉+�Lk]�	M���!����]b���s����ڬ!1Tլ��!��r�KE�ݧG�Bl�Wz�}�X^�xZ������&�\!��T��wV�v�W��ZZ홵c4������{�-D�m��LG����7l�t�6ٛFj=��4�]�g��;$�i���+�{>�]w����r~��^T��A#Z|��9rv%��Gڸ4qnn�X��s�5↶c#�������K]�%��\e��9�xP~>�}�����c���D�:R>>���i�Dm���y<��t��3J�y�~ҟ����GfG�j�Fݢk��$�z£pR�>��u8���W���1*�髾�ٯ��0���7���7w�+�k"1곣�%?Q�q[;��T����� ��)����~;��Yo|f��R���'�ޔ�n��"�]�bМ��������87��ԝ��>
aq�ztq�q��3'RJέzl��}Ys	��K��{ت��KR%�_���i� ��߽v#�1׏G�^Γ��b����S�z�L>�=���PG];<ٜ�]�ۗL$�?R^��4��uyS�<�%s��[��]3�郢�}1��Z�����*���@�@O��Jޥ^$����ǲ�U�B�t'|G�b;�B|�y�3�Y��W�1�s����3�ұ�G�r��p#&G�X�*�,�{��\��<a�Jќ�bn^`�dl�y0;�JW�-�{��a�[X�B�ȶֈo�t�z�f�vѫ9|r��%�z�&oOE�I����v���b[z9��
�%��wԫ�$�Y���X]סg���~�Ykn�<�8��vN�����8Ѷ���=����/W�Ѿ�w��W�a
�)~��R���%��mxl��4k�.I�e��V&���+63v4��Vl��s@�'Ve5xn���yԻگP����K�O�-J���n�����ue��Lw�9[��T>��N�?^4]�"޴G���:d�̿���J�����4���v�:vT�T������b4o���.�bǰj�y�h��\��::g�yxI�c���^���В[#<V�g���C7�T�^�8"-^2뺘���Z/r���*�Mn�er7[�w�#M<�$��sҦg���m�%���@��t�Ҳ�XQ�/�ܬj�"�0�0珷�T�k}��V�:�U���x�~��^�*�S˼�;b�d�ͯ?�j}.�*�^�.�n9Z���vSv�.4D��ۓ�P�o�w�+�_D�>Ы���ĳ�=�=W:��r�%�ˏ�Z��]#��hϣW]dt@��Y;.�U�:��7b����]�tf��������X�/F�] -qZ��K�8�=�u:1gv.)�퍐��}}��!��zP3��5���`���K�gr�2�X+��kv(qv��u;N.��8��W0���5��I]J�)�|��}���=W��q�ѹwF�`Px~��ލU�[7d�U"�u>y"���ddo;o^�J�����hWS��^w�8�^�3�aX�TG���qL�}�:�L�b�:z�)W�:S=�%IW�ݞO	���<ҕL,t���� T�����eE��a�*�L�Qv���Q���]��/�V`?S��NlW���FH-S�M�h�8'�U.詋bd.��/�~�?Ys�M���5�ư-�{v}cJ�#k;�`��մ�j�Y1��ꚼ(��T�?T�C�{n~R8�y�y#�<�s'J�\�%�D1�G��f�+��S��7,یȚ���.��Fv(
T�u&^U�:�����H7x;2C�ԥ�vQ�ds�` �u��kǄ�u"}�2��뱺j$�*�,$�`��u�x.P]�x���7=C�,Ku%�y�ռ�+w^�ﾳ+��a{$�k����w���;l�V�����c�	�_���m{$�ԡ]G��<�����������&^�ChWqHע����q�.&��|`b��7�>�1l�FC���Y1�껱�Y��c��]ל�{�duLpS���yk/��,f˩Κ���pE�Z���@r��_p���VL �����ҹX�EEr�T*�)����U���^�(�{�	y	��q҂��:Th�o����X_�+^f�M��w��vMs9��A����^��n? ��\
*�׻w����-�١|�m�ַ�^媿�'���/qx�K렳m}��=&��zݛ�г{_�o�w��c��-�9��폲�'x�ŀ[�r�#�m��ʑ�.i�q�gW ���4G٢p=x���	����?�����I�^����La����L��O�p�̩ۚ�������*_gV��62Jd�9^E���i��}/|2��B1��yM�s��SxZߍgޯ:>+V��Зs}�},7��Q���4z�a�5��Q]~A��OdQ���úN�\7S�(>��ϭuȌ6��\�{�;�|�-�Լ�mѩJ��q��e�0z{iMϛ�-�3�;��>z};������ٛ�����ڟS��z�O׫��dʙ�ܚB`z�MV�����ޘ���z�#>O���I)�7G�k�;�Q�_�F��r�y/�m!![���w��cŞw����]L�z]��"��鉙J/�/ҭt������a��� �n�D���m���XͳO��]���E�X�म7 oq�c��}Z�s�\����b�B�]�݁+�YSm\(uKM;��	 \��6d5�J-�)5��V�q��)�ok�p+�6�84ӽ�|�K�%��o�N�z��t�(awy�̓Ԭ�;�L��9[��lPR�{*!\��i��.�엷lRIڰ%�*��3錍����-��%'���u&�fv�8�%Y�?�w���������$�(@$	'��� !���XBB@��@� �@!� B ��_�HI C�� Mw�7�@$	'�� ���@�_��?�����	I��W��_��������?��F{����j����3�nx�_\ِI"��R����1mmYY*5F����M�~!�Dʏ=�W����P��Ɔ�I�W��Y+*���ޛˬ/
b��ј#�j]��ᡆ����L�&A+f��5���yzl�,S�5��e옌��P;j�����O������45�b��-,�)�(�@l�y�跘K�:A_�d��̣b�SBf��C��цɊ����A<x#����5cmL�c�y����V
6q�I��-ZRJ�������
���.��p�A��?�%pn�xM1�C�� 3Z��[�ًs09l���ț���-̑�Kv�A �*�c/c6Њ2�MN&�p�/oT�U#��^e�]Ɗ���kyI�KT�gm�ii�ջd��J��n��N1zū�p@4�+�Kf�0�i�2��L�	��1�%Kd,K� �cMF�S)7bhTFP�W.ue��e]嶭�Ḏ&��2[�]��I�!�1b�h�G�ADc�k��-&4ѳ�+j����m���K4��#���NRb���:?�d��
h�f���)�w��w�N��t�1�*d�/A�T�'r��Ds[AV���td$Pf�e�#p*�{�l���4�ҭj6�ݗ려1S��M��lP�i���KC�{m^ir�e3�7��%-��	�]��R�9ԻT�sQhڦ���eӌ���I��"��L���.;؜�9oC�,�U�	]IB��f2�����wh�ec���4�0K��I9Y5�a�g��a=��������nL=B���e�4�
ڽ���{	�zR����Ԛ-+B*;�\GC��3*14Pzg�ѽ4��`n��2,���vm7)Wy��,�4�8w[I\QYqb��g��LW�7*T@�b:��	X˔�n&��ٺ��JX0
���+r��(���Δ3.�ei�i7u�$�~7�u����Ǯ��Ҩ���U���5U�f�c�a�-�oX�fe�"��ٔ�8�9D�x6��C��*��i���y�]��Q9�6�Z%@���M����f���e�<��Q���N�XƈO&*�죁�%lD7/oV[��$ڙvM�if�س1�ԚlPL4� ���ҭh`��dCq\5��X�v")h�v%���������=���mn�k$#�S�ک"��屩I���kI���L����2E�)��c8�%��}I�8U���`l̈́�f3�l�W3)3��JZ�t�%ҵ��/�jӭ
dk�{e��l��Ĉu)�W�v�.�u�k@4n)[���L�{Ѵ��h+x��%,c/F(Shj;H]�m�V�@`MS@@VՅ�.�R�t7E�mnA�ã"��n+2�/ei��Z�҆��w�k����*��-�ܓa�
(�Վ��E�ұ~יkkrP��b�#ͨt1i��E�Ra�A[00	yRZvi�iJ�m��b���Z7�n�������YN��S�FES�Y���y�Kf�I�0m�[��P��@��U������*z	$�R]`x�22j��]��#�B�5�ڲV�8q^��WIJF�k��D���W�zݭJ�a¨�P˼Xa[�j��e�xm
 �+_�H�A00�UF��j����V�ip�1\:�0��nJ���eՖ��T�Z+1���I��pR��v`�uJ�Ӭ�S���c7K�9�I�H�i )09���q��372Ax�e�grl��N֚�%yD)X`]�׳t$B�Z����/�S�!��r���~�e�f[j��Sk+q���f[݌�Lƨ^=��ڨ�i9�v+��"тlUww�;D�WF�)(�R�Y�܅�����"�i�`��۶Em�Cb]�YKB����$i�a��]�
���Z'w�C,�6`tD�rbѬ;8܁*W�Ջt5�mZ�IF��M��
}���'p7���ך7$yǯvbC�JH�]I��B�;�QH��pՖ�Gt]\��ݭ�FJ�R��.��m^S�����X��I��r�R�M�y&[G����v71MA��&�=G1L�`.q��C7��Pڕ,�+3��&m⼰J����
�򬬴��),�AQ�o@ �-��j� 4�4<
�V�jm����6����mK�BC@�B����&^ޅCu�Z٠�=�&�)�Y�*H�U6�5v�\o
��w��,��MdJb'��*��u��U��F2r�C���j�G�Yu0��Z�b�F�����jTY�{Z�T]�n�������I 	 @�!H�@�@		 �'�2� BBH� F��0�H!		"BBH�HI?����� ��[?��S��@��?�?���	I����BHtI		�@$	'��R@$	'�k	 �$���0��o��lѨ@$	'�� ������ ��� �$����3���sG��.d �6��������@$	'���HNo����
�2��.c�P%�������9 ��>��� �@       h P  �   
           < #@   B� 
(H E   @ (      (       J ,�(    ��HF���N�����ޱ�;��*�twXk [�EwXjH%����;�_@�;�w��q�qF�������z缵a޻�U^��uJ��*u��*��n��V��g��S{���R�9�+O� ||� �  ����YUo{w�ּ��7�:�Ѯ��^�ӞRB.�Jh\��ig�y��U�wW��o{z���% �w�5���J�� p��n�k�n�ʴ����綛]��f�底#��IO=�꙲�W:�J��R&���n-֪�Y�j< @  *(�^ƭ�n��Ex�USy�^Է��*��E3�^�{{�U�z�J���绥P�=D��ީMw��Jhw�u=D֜�u=[5�gGl.�R	n�S��wzR��=Ԟ�ް��Դ����^�K��)OT���m����{jiM�nz���7<J    II�:�,�:��nP���^8^���OMl��H%ޗ�S��m�+��x�Yoz�����{ҩzn��U{ew��i����V�y�E=n��^��s�HJ�J���rZ�޷z�m9���m���ꩻ���{�-n�ν�[���o;��	�ݙ o< �     �$� ��=\� ���Z�=����(����z�4���=n��z�`��("��g=���� 1����=D�����C@�� ���ް;v�9�T� T�6U*� d  j��I�)U   S�ڪUI�ɓM'�T�eP�h2!�S�ʦ�UT   �HTM�����L�)��"~?��C����?����j��D����??�HH@0�@�BxBB�$����?�HHH@?�d����BBĐ����S�_�[�72?լ�wL����X�������0�me�3��т�+��&d���$�Z�+ЬB�Z�0X,�`�a�ĭF�q�ow�/l8ì?��XW����I�4���,aXsRϘu�a�8��ì<ì��vaXq��,}k-�ZS|�/wq���1�3�%I�7�CYJ<J���bc ��aϨhT~�0��пP��v��!�(y��8��aX|�����ق��q1һ����޹0J�J��*bwّ6����{��'�=���w�縷��<É��ƭo�fe�yj���e�_`�팼!���Ϟ7���=�'w`�c	����ˎ�o<c#����[Q�V��6�m��fe�m������Ls33
�(ԣZF�fa�3��L[q�-�kB������+��`�F��B���-*�YD-e-����`֫X9��`�JZ�����l��d�e�&9��	Z�KJ#��E�n3�e�Jб��B���ҥj��32V�F�J�.\L�.�3(W#l�)F��L�Wr��eua�ļy�LCC�E���������ʖTF�Q���-���Ђ�e��9�pt"-�Y�bn�3�Q�X�*�T��q��=�;�1�u�<�1�k8�L4�û��'�0������(Z�����X,:�Q��?����7��ؘ��J�)*�U��sF���d	�2�>�??�a���y�z°���0�+0߬:�l8Ì:����1�Xc0�2�k1��9�0���:ì>a�t�e��iQ��ɉ��<�L8é1�a�CL6�a�a��y��u�0�1�0Xi��a�
�L+
��1��m����P~��P�!���
��:ú��`���a�LN�0F�4�l1�a�a��a�0Ǭ���i4��,8��ì1��c0�o08��aXu��@���3�~����<9I�1�!��`����l6�5B�Fl��`�F��m��eem,��J�ek��YX,8�_]2��`�X,`�%`�X,����2�`�X,����`�X,��X,Xy�0X,��`�P���`�X"�,��E���7�i�a��}�'�6��>a��n����!�XV�0��q�a�i�g�=gO���I�,�f�q��q��r�C��������P�����7��m�`|�lӬ�N2VcL��'��a���U`�+&j�I�aXu�X(sVa�H"a�c�1�5C�+��I�a�0�`����l:�L:�L6�q��i���B����0Xq>J��>d1��Va�`��P�,:�l<�L<ì1*y�g�a�a�C��k!��P��{���p�[s����fXy�9a�a�c�C�4¤�M�3XVTR,����+{Y'��XsV��Ͳk.3l>���y�i����9������0w���+0�Xm%x%a�aXx�0�XV��[0�ZʓV�j�1a̰��`�
���A`�<6��a��Xi�����+�Ն0m��ۉS-]8B�B�ˎ0Qt�h�浜���[j�ˁ�a���ö��ar������+�N	�-eV���e�D�ѣb[�َ����0x�u�1}q��W)Gz�q6�w�s��]Z>I�R)]�i���&��u��^�^����'Rm�7T^����M[c�E���%���6Z���ZTk����2��M]fW���Ԯ�Euh�h�l<�U]e�]�ʤ�P��}K2՘��ʿZ.�Qt�:�����bO0֪�9���q�jTm*�؊�b�z�f�+$��ì4��6���I(�m��i"�w���3,8�I<��$X^�!��q�J�!�a�1-�RV
M0Ri<�tr�q;�����	�g��ƕ�6���d^��E#��t���ׇ-j°r°m�`�aۙ
�ya���\��XV���aX6�L3,+��C2�WY���d+�p�vٟa;�U�Z�8��T�\��qLand����fXu�e�X{,8���m�r°�Xm�i�r��g��{a̰��0�X|�-��ҭ���Ug���u��ré6Ì3,1��a�5�a�Xy%aXfXy�e��4��e�������8��+0m�X{,:�9+_�oY���]�՟n�and+��d5l1��
��
��2a���aX:��aXj�B�uaX9aP�&�er�4�2�ڊbTmk���l��B�`�
�����`�
��39L�enX\��k!X4�Y��pK�%aXn�B�m�`�
���l+[��1�l+v-`�H�
���l+�V��7s!X6�8��\�0m�`�
�W2�l+٧9aX6µ�fd+�V��%�-�w�+�w�;�t#����xOt���J�iaX6°m�`�
����2�l+�V�R�����瘻��-4�C�Ն�sz�u�2�����<�t��a��0�TN'S�������`�Y0�Xi�7�
��a�7�a�,+e�w,1�l:��k2�w,8��a���J°��탖�+-�����4>jg�h�r���6�f �*V��T�7�t0�T#h)��^"��5Y~1��,�R�L.�y4��'�o-TVa�	_��F��E����6��][�i����i��1�j�w,1���6�\�4h�.۔���)f��a��c���:�8%Uc��V���&��d�t��UL�b�&-*i����z����c1�&e}������W�V;ị�޳B-iE��a�5�d<�^��1��E�.��5Ҋ׭2��#����J��S&%N�04�z��P�����a����W/)r ����C��Xr��C�a����Y[a��$;lǬ9�
Ùa�����9��r�{B�Ǎ2�C-(���
�>�ȏև�X#
ùa��!�fB��Xi�i�3x
[~��+j�0�XV��[��Xy����ú��X9b�;u�����6�w0�m�c*{,��q�9J<a\B�}�bu*{W��.XoV`�d��Շk,8��z�J��etn�n��Q�Y�_2��Vfl�\O8������ �8���d6�2��=�IX,5l6��{z�X6ì7�a�aĕ	���>�bu&0�e��a��2Ùa��q����;��9��Xs,<��a�M����l��ǔ�2,�n��:�,�<,��"��+���0���0�Xy�m�e��w,1&��l=�)��G�0�¹Z)�̚�hcV�.eA`���16�ڰX~��m�����#�+��`�_k2/}������(]X`°iLLar�ˡ�R����G)���\��=�0�Xq���E�����l�*`�Gm��e�0��
�Ya�݇w�4����b�(;h]Wƫ�Xb��Q��a���%�\�-1�9J�Xv�W��4����bq&0ۣ.�棢���y����j��)�XT�4��I\�Q����e8��{���)߯��f���a�k!��a��.���Eݡ�p�Ɖ�aRi��f�a����M'���P���8�:���J��5�d�aFB�H���gZ���y��a�D�K���R�ݠ���y�t�{V9�Z�7�rִ7eu��b�oX�E�V��G˪`�%e��e���G�������u��Mz�j�L��k��a���q/�*���v��v�������/(C�R
d"�1A`�P�6ª�V)P��t11���UZ��L-R����(�؀��LtXT�YhX5J(�B�os ���
¤
�3�������+
�2�-,l�h*F�B��HEЕV#��
H�-k�T-�DUJԩiJ��0J+kDE����
a���2E�1�U1�F)-3Dc[m@�ձJX��
 �(�,c��Z(ł0D�
(����(�
��*%F�iXT��1���Q �Y1�������)�bȤP�+ A*��X���Uq((c0�#$V[b�J��*����*Eb1LJ��Tb*e)
� ���R�,D�Q���"�E�b���d1�@X
��U��U�c
�"���AA�J(�X"!+�@���"��(E�X��Z����Xe�bcH�1%��UABbVX%�\�PQEU��L��(��J	P�#VT�9Q��TQ�2�bAaPR
C- ��\HT�+X6�Ve�*Qm�����bC2�$X��J������QU�Ţ���`�j�EB�\H��-q�+Z�*� ���ŴEH�TE�Drت
AH��0�e,�D����X�HbAj�B�3
�(���Q��f�+Q�R�[V1WQkZ�+K+@̤)��--������HbTX�J�Q�+��U��Ɔ5-(,QT� �fY�"cB���m�em����I\,���2�J��UTb�1�Y�c����"�a
�!X`�Eb��-� �,�(�2,��E���J�2�,��A�Ȱ�Ea*)�`EU��T"*�*0�pV(��(1U*�S)P�+�P[k��"��V�33Z�j9���R
E�2TH,"�ILd���2"ń����R[@ �.R
AH)��3,!�
�R��[�(�)���1H��HfY��H)
����RJ�*���((�f!V*�*2�R
@E$*AH)i��$*AHe�Y1 �`9IX�A�-��R�ut���{�������wc������c�� ��8@��  ' c ��g��L�D\���˲P^��#y=��m��`<�	� ���8@x x�r�� <T� 6�m���ʯ��    *�6�    �c� l~~9�uP����	��8@y֖�޷Vn9(��-��������=r�<Q�Pv>-�.�,n�q{�<����Xi���1���Zі���fQ4a�8��Ѣ-��������9�X,�v"�l�A��D����)�c�m��pb�us�P��f�`:��ݼ����V͂�����q�^:^�h6xӵ���.��r�A���̷�
�c'	�ݥ��\�q�t�Ts���۳�	���u8p��{.�p�(v���;k>ٵ3y;C�I����<�,�H*�E���<��=��k֪�drܳ��HV�m��qpV����������n��ً�طK���@�d����7W���M:�ւ`�۶#���V����s���I�vɗv�c�\���u��6�EŶy�8wl���6��&ݞx����77m���W\mN:�n:;Ly�ɸ[����iĖ����R-�Ň��1؇�\t��:U��H'��z3s������}���Ѻ-ѝ�H6ݷO�8��a1���Յ�U�v:��ݞ�g
�p���j~�s�>��2�k��F8�[��=n�Sp�帎��k�ݮ�����5�5���g�!4�#��k�`z��;:�q��tN������9�,�>�!�8�z�I'd�a��Uv�њZUUU���P*�� 
��K(��@  ���mT*� 6�  @ W��� M��eQTP U )��@
�mwU�UV� U    =i,j���R�#�A"�P��2A��R淪�;�@ 
� .ZV�n�[Vva�Um���U      � �v��d��h��HVQ'l��K�� �*���*+n�mR�u��y���wk��uXp
�\+mU @ @�Al��PP  ��r�  �  VP  �     <x�;Z   *�ܫU�a�8~y��f��  �P Qz�d�z�]
�k�B.J�u��R�K�;e
�P�@)�����]5+��� ����p���    ` <  ��uA�� yYS�1�p��+)Tzڪ7s�U6�૫P �傩V�:Y�0'	����p�U<�8�ϟ{���m�mܬ� v��^�]���EP@�wh�՟�aùP�^�2��`��U�E3Y\\e�N3å�eyk�Y���0��˥W0z�n(!��� 
�7��־�  6��� ��c7j|M�(����������*x���� ێB��h�]���,�k�g:S��j�L�F��ݬ��m� \���TNU�W
��m��Q�+����Gu��b���,���=N��0��Pt������=]E@�@  VPV�m 75@ U �> 5��;�4���V��J��A�J���@�}f|�P�M�*�@ ,�*���P�*��*��7Eom��Um��YjD	 	gA�*U�BUU�eeb��    �)���* �J�+m6Kd l�@ 
��GvSl  �Q�  l
�ڡTT��%P@
�P w   -��S��V�[� �'���n�v��TyT  U  ��.j� UU6���m�`=^�Y�U���Sd['�]�R�U-��:�g e�  �� *���R� V�  U����AW�t������H�J�-J�7b�i��Z�  ���V�r�ͭ���W9� x�T<��p�����s� j%PKHҳ-�/�Ux8V��  < �*���檽@U ��(p��T 	��`m��uek� < <U��0WR�x xۻ�uA©ꊧ�֫@p�� +�l�*�5�0�7���Wu�T��PVR�^��UwJ�AC  1�  Ux=P1�q�S�	�PT � 
�      � 8   ?�>    
� N      � 
�P U     �P       86J���*���   �� '      �     � P �T�U��u�[u��EP  ˒�t7H��9BDXc�6p���ʽ��� dL�UJN���N`�
���#e�:s
�U��<m�F��W�)y�L0A
�"Ӷ�M���'�fm��3�SkaH��	��3̴�m*d��d���m��C��*j���n\GuJٖ��Z��cxYyƘ�{B�Y4E���GF����m��{V�lֳ�R�R]�3q�Ƀ��1�h������#k&�ݐ���%]m�qDoQ���M�M��J������cnx����=�8:�v�]�v}1��Q�2fv�]M#W�c���X����U4l0��֗bۑ�dJ��"x���h���N}�{6��J���ƃ���iR
:��Wml덐4��d��k-*�#��*c������q���q6['q��_Mn<;�5�����W�)Z�pww,.���(��B�,r6�0v]��B��� ���e�I殔vV	�JO(`�s;g̓$ʛD� 93�L0�es���K8y��˗j��  2�r�f�u��rP��,�T�7��m�:��wC�*T�l�3F{�͆�&s������'�8�-S`q$��f�*Uۭg�5U Q,�݂��x�+һɪ��d�w@�9��{pY�NLqu��5�[v�T}!p��(����A����6Rs�8�N��n^����c�����p\�l@HJB9�k��vL�V7<Nꇰ[G��,�®�v] ��5'+_��_5<���Ҁ�:���Vu��-<:���gҭ�a�Le�!��*��Rm�2J�b�x��m���J�9�Pv�.�I�Ů�;��r� �|                  VP       U �*��                     *�J��  *T   ��@       U 
��>     @    OTT�  U  
�     2�.aR�P*�*� �      U    R�    �  T    �|  �     *� �(  7v(�3j��U@m�
�6���}U�U*�P`    U �PP
�                   U      �    AT  ز�      _�}}� ,�@[%P   
�� P�    ��    �      
� @          �6@  �ʪ
���h  QSH��U*�աGTm׵�[k(           |   �U ���ڗ�U              U     0               �      %6� @ ?�|            ���"�
�     ��TU B�m�            �         N     *� 
�  �xmV��@             U��@     
�
�  �+�T  *�         T     � Ͱ�c�mJ���ʹx7�T�V�T    �6ʀ  �5�T���z��۞�C��� U{'����e *�� ���eT �      @  8��,@       Ub�l�     *�TEm� *TP��� �����  �  T��U7[mU�                  T          P  � U�T             �fy�v��� �> �)�UU *�UU � {l`��  �*�uN�%@      �ʩ�;���ѵ�7�� U�� 8J�mE[���]w�;v    Y���[�� � T[j�(    T���� �Ÿ��t�Yvx�\����na�	 U  ���R���w,�X��u��1h��#�*T     �U@�U�W���U
���T�eP  ��f�z~�f�m�y�7o�U׶�߭<�]��  N3ӗ��,*�� � 6�nwO-���c ��׻̱��γ�wk;��P �S�P
�*�������v�G�h>��X�v-�N����� �$$��i� BI�			�� ��H/�_���kZ��b�WU�G^���|���|�M�P�wSk6�@Uwny <����J����ןnw�T.��a�W�g�w糽�u��֞|���kq�Nƺɧ=��{vxk�-����5�uB`z�v:�g�/;ۂ��x�v�փ]�^�9�=��ەӶ���g�m��y񳓔��j�f�T.`��@�S` +2�ֻ��v�黶�.m� 7F¨g)3�"ĵU 
�`  U�����.�g��ʷ=ݲ��pV  y���L����R�8u�z�7q��
;]�\�f����
�/ui�@[�,Ί�ȫ��UQǔ��]�����@�;�mkb�T*� ��]Q�d� �� *���UE��ڥ^7�z�� -����q�Y*l;�� ol-��YU�;��kgZ�@�FuAªx x:�k�=U�m�j ^��T 0*��@ m�� ���p   �Q�n��@��h%d��R9Y%�nt�VE�P@�3iG��SoG\u�e׭�g��rv�����EN�mQm
�݌�9�Y0��5vUJ�xzظ*�f�P6����n��e�ˇ�]O���ˋ;���sE��
76]�v@[jc�Y*���s��)7��;�n��%P  TY*        �� �T ��UP  �T@ fکT*T� �      T�*�UJ�@ �R� @*�e����  �*m�   w   *�\ʕ  m�  *�   
����� �̪�T =m� [�lU��   * � ��UP       x  �TUw  *�[h �tM�b� [[ �� om�j��=u�� QT���s7x�w]Js��T��5[^ݩ	�g��}�{���y���Ԛ �P�2b
�Ll�K`u\Z5ȩ�u�Wn���c��J�MQu�!HWC��[-�C���9k��V���w�w�h�
�Pٴ�ܶj�-�R� #�D
�
�W/f�oGc��]���q�Juj䝍�	�E����g<�UU 6����U 6 rإAT�lU U6�
��Tj�*��m��\�Z�΅�c�\������6����	����U���r *�+�l*�aL�	(���?��������~�����+��fx�skk3��B�d����GE<k����[��V��G2�\�w��.�����28Í�Kq(�P�;�^�[.�Hu+�^m���+h���,�i�IS�$�
�w�^�k|v͘���F�&��ި��{����	i&�e��7k^��gu�}#������ʷv�jӢ��'hdl����dD��un�ĵ�jS"`n:km�jR��6שP�%���X�q� �k�~�^r��fY/|g���:[�۽|,���{��Xх��S��y�^f�N^��m}��'�M�#Y�ԕ��t_����̒���J�L�I���)�+0:�Gv�or��~U������G���^f�$���q�*k��q����i+���ea�}�94zS��aH7�bh�c�0�L�4V������ݑ�e_�vlя};}[��'t��f��l��HP.�F������m�Wp�z�&����B��a�r+ջKm��ʴl�3++1�ٳ���g�ۿ��}�oG�;*��-��dC1�k=���г�-L��㛳,��3{ú���\�%$Q8��"�Quw{հ�7��p����!z�N�e�ǵ�5lM��^i���Jv�8�p@K�$�l���*eg�o3,,�SQ�
�m{w�vطM���DH�Q'@���;�����۵��zwڲ�j�Y��7g��8.��n-�vu�G�:�`��λn5���SJ�T���/(	z����dU#���ޙ�y~�����v�����;����ݝ�UY���,���F"�;;��>��:�y�����Ǿ3++wa�N�]ݜ�"�.�lBCn$�K�p��3�A��j՞������u��B���8E��D���y_a��gp�^ߧ�Ç�Y�6w�6*��^CUP�D�Omn{��K�0������C��vi��wY��N�{�2��7���V7�+�(ŉ`�"2ёͲTv�2���MW^߻l�8� �6ǭ��M��F#�� ��*n��&X/|�}���y�n�Mɕ�j0Rj�q)i�1L����(o��̺���B�t[���v~ŕ��@jմ
0�W{w��5>s�<�3l�٣^�c�����̼�T�m��!�\���&y��p��u�z��x&X/|�}����Y�����$q�܅D�ٵZ��)L����p랡�Kˋkk4祉��Z��U7w��>��l{t�-7Kx�{�΃���w=��Ƭgı�*�� �R�Nl����v�
��;�x��ums��t{�+7���
�g�;�U8�e@%m"�uR�@�@ 
˹S�3��{`�j*��A[Ui���Vznj��7�   ;�� �    wm���*����U�wUw �� xm��Sr�UR�F^����iN�-<gwV�禨l���v��� Ygq�F�v������[���x��КMH�e�r�EÂ�M�u���r���ͳ���+�ҮmM��d%E@[���t=��\�2�vt��壼f̬�^�f��f䫖T26�"�I��▭�]Lɕ�+&Gǚ|svm���men�z��m+1��m�f*m�z��՚���YS����}�����ٳw}I������H�!I&]{:��C�w��E�u�c5�f��Q�[�����ٹ.֤�Sv�gU�(���=��{����UA*��D�,j�.� mIq�X�ž��w�˖��z�l�;��e;���ܧ����1ġ�BR`���k%f�զ��Xr�~&B]'���ƶ�έw��oǝl�f�\�p5"BBIp��E8zt�=1���4qf�I��d�=[[�}Sk7oW��&�-Ȕ�C
g�������uj����ٷW�W�[�����o�4�)��a�:v���ʠ�4��6z�Y�{�f���͙��	�I�� ��F�ڛ�un�L��^�*�� �;�[ ��"���s��J���~���;O86�fˎd�k��v���2,��ƛE71�H�ܛ{X�ˣ6�{��l��V'=t�<�]eʬ2R�ÒI�ƣ����NM�d���k������֭7�{TC�o6hثnl�5m�?FXrIa��<�C3���	�;�+fw�l�˼�XGz�2a-��B%I�	H{++8w�n�ˌ:=�[��<�����ڱZ�4�~h�"eA"ġBQ�$\��UL�q�Sq;�h��OUWpU[���ab��d�V��y�������ݢ�pVi�Tm;Ɂ��D[I���=~=���꽔�y���;�_�������[r�Z���h	?��}��E~��͙bz����ɀ��o���Q7$�2Zq�c`4��Y~�y1f��qⷲ�z[�o{p�T��K��ٚ��D�lrյK�e��N}�i���+y����xe������C��"�M�"�Hr9�.��.�LS��w�W������ѱ;R� �ڦ���P
�s�V�s��Ŵ�2b��/�>�����!�$IG"q)!96�����h����|�A�ӧ�q���(�D�n2Kd�J$�nM�Br��{�w��9W����]��D$_�n%R:�_�ͮ{�
5�2�+�|����檐�J@L�$��3��meu�G�ꙕ�7]���6�h�Ր�[��������Vbu�n1�ڸ�o��w�l?v�`놳��CU)B
`��Yݢ����q,�o6Ƹ���v�Hm2��-*��V傳uv�۠����^���iu0�T�$�,�v�1�6�lj�>��6��] ��( �
� *� *� w7�P���*�[`⮖+�-�������;��ȵ��X��t�7RU$M����T�� ����G��*���[�rd�R$q)$JQ�cC��Vq���Ǩg^��U_I��Ă+��BD�"�헧���ŏ���e�(�ջ.��>:��js�a[mp,(�hV�|3we��6�����g�fMγ]̚E�P��$Q�ۃ�q�3��Wp��Ι�G����zv��.+����6'��<�����~sE�l��R��{�����`���c��7mK��!nv�vI`-§�U�U�Lmy�#J2�q��R:�z���^�%e����I�b��^�6�#��ㅰ��3|WWjPR�^�||w[x^�:2�H�\k�x��/Y��i�_䮯F��U�[OM���Fo��vrl�f&Kz�mH8������"�~���[�sq�L���Ҡ�$g��JF�?�YYou�{��^Zt֬7|^�����I=ϲAጪ�(����6�OW��<�n*�]�URA����,��ض� $k���|��<�9��u\�n������/�nd��M��)Ȕ�S��iG�ny��ʾ��nC����{���|��I�B�hZL�|�����������$�
���a������"Ì�m ud2u ����<��I RQç&˼�+�����j��T��>�x�ޚI̺}����o�d�����3l:�J�?0��2�6��'������@��$ɉ >I�BN0� i���P��B���q�aXd��ͧ���O���?���Y	�I$�����a�??2���!Xy�|�O�@�E���Hio�Hi$��>C�1T'i��O�q6§_�g�:�6���=t�|����q1�b�,��=��q�d�i ]�+i��1��Bd��$�I!���T޵�o�����zF;��1��P��&'�����dY��d��<D��T�Dx����B#K��i�E����m��!�"A�FJ�G8E�g]
#~X8�xF�4\�5g��9����D"����cI2,j���?�#-���jA-�%�GR�5U�ݸ�U9��I֑I�C)�x�!�����ե�#>V{�Q#HDq�t��Fr8�!K�`��s���"&$�8Aq(�,��"��I�Ň�s<��KSHs�5�7=�o��o�4`L�ӄ��{��v_�P�[4���7�慬Q{�}����j���(G.�άL��ۤ�����E�05oE��STa���=~����Mp�"[�F�Q��{�Q�v���n�γ�O;/����g��Ր�$M���&�8�e�ؗ0��`�O.�*Uڥ[����5UT�N��v쪪	Uޟ_t���s+�vUukOE��Ow��޾���InC,�`�F��n�����R�l!��}���y�~�}��k&$��c �$�K��[6{_{����x��8��&�ƇG��n�df��&��CX|FpB��0d�>��FǏ��E��!<X�d0��B��;���@ʎ2Z24��2�Y�$�ʆ�$gC�� a�g4�?R>'_��#L5��ύe��o���ܚڸزH*����j{Z6�L/�WB���N��{��_}��_U�T�mۻ����*� Ɲ�t�ۈ�]��x�QV������[n�*�YKknTm�
\�(��J\�'Y���g٥�k
�j�'k6��~�P  �  P P ww�
���T 
V�`Ph*�*�h pVwPYt�y��͊q���O���l݉2D�u؇���b��B`*��Z�0��^����0	(\M����7��ʝ28��w�������\Y�W��?��lix���pT��4l5"M@Jq�"��!�\h���mB�q{	^�6*҆����Ȳ;���TDD`RD�I�S�!Y��3�%�	vŌ"����ts�D"���D�������R0di��"��"&�dvl�k�qCM�#���Da���:^*��XS�Y�:B#H��הZ
�A�J�i��3�<�L>F�͒9�DY��A�K8F�e���!������C�n� Ov����2����ӷ���
������� �m����eZ�g�~>_�������uU�!;�3�BF��ő���l��(�!⋏�$ɳ�+�e
<��I�����V��#3s<��&}~�Z|{����x��2����i���;��Y�GH�oOt��|Y�o{��ۆT#�I�&jg&w���q|�Kj�GD$,���!��cy�;9���<�{e�5	�����������8ݒ�(�!w�b��&��Ԟ�i�p�Ԩa٣u��&�Z�Rq$�P��#��(��]�|���wU��Qa��SCHY�f��#�V�Q@��0Č@���25֑^^�f���y,�k#3EWp�x-�we�[&Wq;;m[bZ���0�Ρ���hdSx��i��2��:l�:��#H��{BC͸�8�I�rW��G^��ψ�Mr�B6x�,�����Y���8Q�Uu���bH�-�����GM�wdqP,���4ۜ6��=��Ȉݸ�_`��o�]�j�w��A�8���;SWW��g�b���̻��4M���ר�󳻲�W+ܚ'�e��P��DGDY�1�9�Dq͎��FƑ�(�����x��Y7��
#�����_�R��d$#*�j��ER���K��w!���Wj�;2�2��75��#h��. �(ݑG��!��t�i�Ύ;�8�"ȏ�T:,�0p���(�0Λɲb*�d�a��-P�#ft�4äx���J#�8�(}�⎗D��N��5�n�f[kS��MI�������Pg{s������	��Y,��0��<->�&vjrg���^R�ؑ�T���dx��8x3�x�F�ҧb����tqݐ��w;�ރY^���\l�S���$F�[,Ъ��L��<�hql�F��T�F��Bz�Pdiw�3�4�,'��&[m8$b��#5n�d��jtu����,-��VdUm�T��m٭+q�K�m��h`��������!DE��>(�g�5ԁCQ�!�68�"Ξy��I��JD�.�.��|�x�ç�+^8t��}�8�#���H�
�jV����QiS�C޿��HLRD��B��0�:|xp����D.��~��<D�:�R#�#
)޺�q_&|�
$� �i$Kj�ٲ7���L�68��8���~�!��a��W���ӡ��j���"&�@�3F�j�T�FWBo�#�Qnb�*�q����3�
!�F(��e+t����s�εkU�	IA񪪁7����S����v6�SZ�f�;��:�\�e��G��E^��=�]����}�|�m������	:�d��U �닻�Uw]�u <�̠c� �;1gu����[�'GU���U;ɣ��,߶z��  �U  U    =�.`��w @U Sy�m��� xm�pm��RYZ�Nt�㳋���NK��Uڦ����登h;�w)�P��O�����5T��.㞈�*���ET���Ƙ��Ǝzo��>�3��7^�E�=fu"���6��L��O�����P���z��B"H\L����=�t�"���,��Z|D�����Q���@�m�
A��"DP�i�!�]�͛�"���Y!7
D��Rڰ��qx3Fx�B#����/���6�&)��C���Wd"@�̠��9p8�,p��n�t���Ɛ���-����e�`�IB��j��l�0��-Ub�{2�7qh�C!�qN���O���d�k!(g�/߾�re������m�BQ(k��\Ic=��`]!4��*��U[�Vc��̪�.Q��2��=���fy;�s�y����d鰈�*�j8Փ!�FN��d���ǈ�����I1"Q��rF���!O]M�0ɛ�-��U{��F��u�!� !3dx�-�Oo�����o����Iq��̈���|C#=lw����(x��eՆ�Qz���R��]��:�z*��Q��ԉH�E8�H��cﷶ�����!��R
��@�68�"��K�?w�S�<����[��Em�مA�/�ǒu����t��|hۢ�������4F�g����\��z�б�cU*mU$mٴ[<�vY�m�U2 �6T��w�������d��Ģ��8}��4�,�F���`��dOVuZ9S Y�p�"�i
,�,�2Q.��5756�[�$'��1�ś�qP�'Hfږ�{��:Ug=���g_���L��%I$\�$|h�!�8mvJ��(�������[��v�[7%���aN�C�GO::��焲��?fFUܑ��JD�I�5x��4|~/�W�����B"rt���m{���}��BD,��w�B�%B�&�b��C"B�T`�|�Mo���/�F��<,ϊ#�<�)�I��<�z���,���6J@k(M�ڪ�i�qBu�
K�
�p���w7��E��p7d���x�H_��Dq��Y	{/<wc�4g��,���k^NL����=��j�rX6�2�����#��H���ay�-�p��Y���8�QFwH\�L�lE��6t\���ڠR��񹹚�����db��R�c���f8+[VHN0�N�a����<��Wj��S+=Ѝ��7{>���"�0�-��0�DYe���b��P�Q����0յ���>�e���zg{���Z*�1�\(��E#��We�BP4�,Ng�"��4��r4�^�}.|QGtm�%���ݴ����2*�ҹ�`X�V8u͗k`촫R���2�,���<��&łB�[�D|a�DwWt�Q#���9 ��N�{�*ӤY�7���w�o!�W<���9�"L���_ۄ��w;��Y�EO���V+�������P~�T�}�A�rؙ�U��5f�Yd�Bn���x���F%#�)a��?#��/�n����5�;nG�V�-���ve�y�����O�Gu�P<F"�+�G(\U5���gH���#*rB[m�`���!��!Rk��"�a��V�D#g�d�#u�<�}pe�1p	�d`�@_�?��d>HV��4�2@�	�!�4�8��㘽�Cbd��B<����� ����8�&�J����h��v�߲m&�?0��4�`T��� }����I4��&ө$<�橷��չ������`g9�7Ԇ�q�L@���S�VM8��x�3 ��`T	�@��|�@���`_R~��f�a8��CwW'-�>�2y y��1��$��!? VH�̐6�� `_�����d4� c䄁��B}�wX�]kZ�3Y��i8Sۻg8�@NOvJ� 
�Ww�z���9뫫���aW�W;w�]����tV�nlgh9�-�c� m����B��G'��;:s�����V��^��ѷa����mݷ%���2�����t�B��1g�:�vv�+7-�չ:�{r��d���]�s۟׺z� 
� �  
���E� u�vզ^*���P[���%���.�)��TU�� �������*�{������/s�� ��1�.�OU��Ĝa�*���r]
���7 ��M�Q�� n�c�ǝ�:�6˺1�w�=�k�<w��z �*����<�\ ���U�p�Al��� ��U
�V�;v
��ui�,� 5ԭ�U��P PfP�T���.�ǦU�8@y�T�^-M�^�
�[h6���e   �   �   -��U  PdTo�V`ed��
�ra��ȰqJ�VV4�t�`+��ח�r���ʬ�7d�,+��]�J5�@�:������ ݝ;^�B� є��䑶� ���M��YK����Մe�GNC�'�À��%��X�v�<�]M$@/l�H���'8�z��r�7�      *�   �> � 
� �  
�P �      lF�     *� U @6�*�
�U   TU8A��-   M�   �    �   6�eP      f�  
�     e��V�( ��}[�;o5A�  
�`T  Vw[hU�   *� W�  UCb���\ʶ� ���J̶ʀAU� �w;g��5HR��}���8~���[(�DԠһ:��uEQ�����w{��gY�F~���mUr��ج�i�8�7)���M��+����u�u���  ]Ԩ���j���+��ھ�}�G�ͭ���s�q�n�aP����|ue+�����P   
�u�8A8�Í���h����=Uw[�m�5ֶ�xT �T ;� PK�:�l
��  ` �� @
�����TЮ��X�vn/N�B-��G�����ր��'F�q���:6B�0�*�5Pql�I���Ỷ{�Іԋ�RG�0�O�a�n�C��ĹQ�g��Q�Ǌ7�~"��F�Ͻq�(�K��d �ew�53�˨���ǆ����ʸ�h�e��]Z7P8�����DnoQ��\$��%��NC(����ΉF�C�G�8�Q,NO`I���ٱ�aq�:�Pe�L-#JD����H�4y���.Q�*�F�<B!y8���m[w�3�u�oU����y���)$�$�;یp�؟k�K��Q9֞�nz���S_j}�7�)�����׊At��UG��qk��
�
��dR���܍+rB��-�ż�\��^h���yt��n�,a��<��%����/pI�2D�10�#w��7:�Q�U&��qFo�aweMb����đQ��^綳�y|�4����E
E̯��dpxT�xL-Kە�c�Q�s�_������|��z(6�������j�nZ^�og`�2)勺W,Y�{э�&��n�I!1;�g�_���U{<�M�S�hu-����2W=n�!��|ZYQQ������
�Iu۫vZUڥU���f^�g���]֪����D�MD�:֥%ﭷW�V�s�ˠ��w�urտ{�p󫻩#.�MT�����UU_:w������7V��p������8m�^�y�kD��Q"fMUL�*�vz0ûO=���g����*'���d,�ݷX�O�SY���nj*�`������}��t{^��\�7��;���Ѓ�ӝ���"���v�+�A�@�[d��ig:�Wu�Ζt�(�l�M"�i���8ծ#�/��sSs]��w֒Ƃ�q@�+����%�ڬj�['����U	�U	�j�uG-��c�&
ѐ���;3����0�p8�(K
��&K-�f��a�2��\I7� ���MDL�T�jD�m�ZqxJCZG�8��5���^*�Q��N���҈m����~IL��&y7��MS*��E�m1�[p4�|_ҢGh����� �60��V��i;��M#������@�?�* %�73S~�f��q�"�=�Y�­=<GG���o!�ާ�?�'˅_�����#�ya갣!&��B[��FUR#��<~,w��H�@E���&�O�(�)z����2|wG�B8����,?��z̄�",)tZ{#]A�/ n��u2w�«�Ud݉Z���:�{6کP#	���E� ��U�>!�/�q!�%z
R��ў�d�4������,�M��p=��6���R�ٚ��u;��ױ68���#1e�(ʁ�u3��#Ǉ�s��$G�"k��@�4���(�5568���lf�\�ada*�%q�S$�E�D��i����44�t�j��E�f�l%I#�GƏ}d�����f�Da\=���i�_J��P��<<&l7{��ŝ �L_V[Q�Quɽxnrg�\�ޭ��yǶ�o��DaӇ����F(D���B#.;�u�HMtE�����j�F�٥Z@x����s�n�t�߻����vm�hF��� U�b��Px;�wVP	�w�7d۱A�}�[����Bؖ���v���U�շ����W��0 ʠj�;���<TU��Nu���T��n��GfR�ִ��M@P�*�
�    ��`��� �6�/wV�lWp����mf�dt��-�[mԑ�<��;d�K���;[&F�W*�Ŕ& 9X�<i�%J��l�QU�2�[.偀Y,�m	Y�T��\fv};��ٱ�a�Fl�sl��?�!��*�9��Ɖ?�l$qx�{�>��L1	�T���ee)�G��t����3Ƽh�Q¸lc�n8��x�����#=�̳Բ����q���W����|d�,��_�Yқ�ضE�����B,"3a)��G�4e@�R1"L�ڭ���'�9'����v�8C)�F��a����hc��p0��U�9���&g&ff"P��"�GN�<P��Sc���iuD3��5��4B>8P�oո����u�O��d���r�إ����إ��Jl7n&�z��Omz��Ul�U��F&
�H$�9U�K�K���z\���!�yW
2�"4���s�0��.�;3�7��a�W����\fK�F 5����Fk�3ٜ�W�U�_b��dabÉ�@��!q�ٰ��<s`6m����TC'cH��rj���%!$8�Ug���a�~/H�8��Q�&�-"�Cr��mAP4�����ɚ���r
���Q�n�����t����,����Ǖ|k q��W�'q���!�)=¬I$d�c�}3S�59��߼�|a������"1<�!F�u�CO�ΟZ?G�|�~u(��d�ƛ�i-�mV�Q���
sV���=M�:����%&�/?|滂�ȲT����dqPf�`�e�z�mE��p�T`�e(G�^�S�I��U�(�a;;3���/��7�i
�?�ĄD�=�cvI)�da�ʴb3NX�ž��"�Q�Q1M$�nWDa�=9����<~�|c�w�C4{��}J���{�
�8��#!���aa�)8CP"��$�3S3FZq(��#�R�!�=�H�"�
!q��}Y=����m�}�>U~��ZH�I�[�	2}_}^����J����oc��qjxw{�vi���1�o����gD����8VƝ����۵��l\UZ`[{�<�v;ojj�J8�r]O�3~�m}u����
�"���x6�דǱ��m�;�i�H�D�N6Ђ-���C!�U�C��)�B��vHd/@�%�X��D�(��u�;3�9;���L���Y"����9�W����B�v�S�HIg��s|!�����P��1���[N6�F�Q#��#���Y�!�k���["�f�@�ًF8=�������������ʢ4����:{�a�(%1�Т0�pp��P�i�-�W鱄a�yrWpB$�͐��u|g#73�鬓��o�q,U@mG��mB�U�T����� ��V��[]8�b��,�[A�-���&r{9�z⡤x�9��B4��B�X&٬�^��M�O9��������r2�T}5x�Ɩ��tE����|^�ȳ.���:l�l�?LXG�,�|�41f,Q�K$�����Nr��:�B"O��~R,�������Kև�}ԈC#3��f#2D�I�[��אäk��O�γ���"�{��Ql�чK5�f!E���2)k�[Va"/���ff�w�Y�}��u��YwG���i�ʾ9q���N��tl�<2�������}��ͥ2V۵UUU�M���r7//Dn�ݻu�m�3�լP['q�i�<�6{i���9�w�����cF�&�n�p,�+++�����N���))R�   #��#i��'b�b$�M�T�h)G1������wuW� ��  d *�� .�;������� ܶp��l � �W���{�w[��/Q�yza#q��4��'^r�TUmK��\+<�����z̄�!UZݷ�F�2�#dB0�?�f3�[ˢ:nl�@�'����FtO��p�#��(Ypח��XABAc�%ISW2n���,��H�9�ȸ��YR^�qe��Io����mԐ��:P��{-Z�ۍ!N$�h��F�'��N��,�B�qq�J��Ez�6�����#{�U��@��`L�@ �W7;<��7���ɭ|�3�iÇ+����4|�x�y!�5외�����#9
^��G�(�,��t,�5�7�]��C>d����i�CO��TSQ����ߦ,"0�1y�4���㶌ݱ�g׮8��
�a�we��!;T�]U*��UR��8�	���-��fny�9�>��ǿy�&���^:��i�-�;�E�=p׷G�#�g���0RJ �D��I_W����[&�w��v\]�s�ۻ;1����>�f[T4���G�{��=<��a�G��4I�E"M��!���;�^E�#��2���E�O�Q��C���ҏ��K�>M����*EH��K�<a�Gt��B6�f�k"v?k�%��oe�X]���{6�{�܍�
����T~�3��T��^����U̙Xhgz�����k���5SR�!�	��][��@Us�&9;d�lU*�R�*��j�V�k�,�wf�I�����j�����ˬ�/MoԾ,���:���Z���Q���QX��Jʇ�s�иz�*��ߪ�p�~~�g|��5߾�aJ�+#X�.2�z7�m5�˧AD5������}ᇼu6_��?��N�1���9�jɿ����m���	1�	P��Id
�&��BI�IԚ�BHq$���S��{�$��!'�I*?2HT��
�� <�		�$�!$���2 m�I$6��'���Hq ?$���'�m��~j����c (�$?$�hCL$?!!PL$Ą�̒IԐ2@��!8�Y`I'X��I4�󣟽�β�IB~f��VH@<�E������$� �0�8���$?2O0Y �M����O�BL|��R@!Ԅ�>@�!�q3�d	�E�d�|�}`C�����BCi8�N�q�^?r�C�2 i� |>�}%�u_J6���D�ڋ���g�̍�JB"I$a�'+�w����t!���B�N컕���_����"0����OC�D�-Ȕ�������E�E�q��r��mZ�"�
#j<t���fϞ��=F׏b����}��OOe�mŅqR���\�{+.��j�Kĸ�@;�SŲ{�V���[r��bH�IE�s���8g��S`I�!s{tC4Qt۫��C
6s����f�]��pDp��(����<l�[�y�~�	g�dzpxx���S���>ɻ��/o�_/�4����bA�c�^��vw�6�f�,���I������\f�WU���0��Un#:���o7�w�u��c��u$�]k��M�ML�W{5~��}uכ�ּ�H��H�IF�qvo��*��>ޝL���M��άY��F+�Iy���~{m��;u�j�&ҪqU ��t���T��A��kJV�ޕml�0b"���g�5T�����i�;U􂃥r��0�8����:ޔ8�t턾w�-l�����-5���ɚ��b�ڽ��0а����#���R���<wP���P���h����D�P�"RH�jIX|F�J9٭��W�B~�����L��b>p4��'J:~�պK'�)DPrIb*�׏m}��8��'pC6Q���խ�#������ٙ�ɾy� �]0PD��"ώ�!W���0��mx�6@w �����4 �:3ر��>���Z1���,�ՙ1U�R-u���/C[���r6���h���ݞQ���)���nf���m�sw�f���T�[@7k`��<!��V��ڔ��U���K�UV��T d������Nv��&Hy͑,�U��;�Z�ݪ�r�=���     P �e  n�pm�T6� �U
��*wU6�©�Ud� +��iY٭kd�N�/U��C���0���U<�{)����J�*�l��8�UV�7$�������#��I_�nU�8�Μ�p6R/b�#)����0x�#�!2'Rad��>?�4t|9='�6x����0��7�Gb�寏�}UQU���77>�N�J�c��h��sS�8P�{V8���p�U�����B�I�\�^D��iF�?W���ۅ$و���PL�;.��ֻ$3G��.���c���~"i�_�#L�'w��*#5Ҷe�?s���鄺�/� J���rtC#N���g���}���.�!?^�Ok���nÞ�ŕ�&��V�9wOպ�6��P��dڪ�@wk�V�����Wq�J��ӆΏ�Z�h�	��h��E�J>-�F���Da��[�l�Gܵ���QmYa /�����M�9ɯ�}�o���;�vCȃ%W��$3;@	c��wb�Μ��,��D7�333�� %�%��93ɹ��fk�����d*�������O���s\wm0������Q�(J�Dq��>�!��2Y�,�gn*�>|+�hil�����:p�6��`��0�)#a�Bp՚ C�u�ҏ��C�5"����r�VK(�D��nq�8�5�;3���+
�`(Q\qm�ZX(��
�8Llc2��R��T��- ���8���-�W����s���nf5��ӊƗ%�E�*�2@�G���Ӥ���a����xp��\;$91e �[��8����ڇU�Κ�D��L��}��𐖒e�bl�����B�ߌ�_��5Ã~�Da���b6\���oIӢ�8��df�z�a��?�wƜ��$h�"*""�������x�q���A��X�3��S#q���F�4�+������I'�H�R���G��i��4S�ᵽH�r���}�ZaϽ����罰x#��&�p(�-āM1����@��;]T�[��6�xZCa%x%`��%DZ��6����	�����5��V��~;[^�������)~�iw�ѩM���
�UUO��{���{׹�Ǯ��^M���#/�v1vFy>�4IM9"$4̍�U��ue<��/9���n��M�������wBC_�$DP(Q��^V��!����h�.�������u���P!�@�w��H�F���b���%�h��G�ˍ#�Z�G<~�݋*��x�q�G���H{68�<l����1�����y��ʧm� z���ewS�V@§�� ���t�[��eMdB��qGH���t����H�i܃����uN@^��ߡ?5�*�JpՒ~|�&n3[��Ͻ���<&�U�G�ᐨYG�,��Ȟ������E
��� ˓m����|��}�b8��;D����%7�Y��Ȍ)8܋�W8R~�Sa)��-�)�_���[�aC�U�~ҏ�=j{���	kGNjDB4�.�La7�����e���������R8�����s����Q�[��@F��������|2(��������
��y-��i��-l��[��@B�7`���gv���n�d��j����$6А��d.Z���UTڶ��;���,w��r�u�(۵` U��%�n�R��w6�Ҡg��   �Ƿ��޽�����F����[:����As��������  *��P�     w6��
�� Tm���:�m��ʀ�T�p�z[/ ��	���h�GC�F��z�9�@!,�j�����R���UpTw���H@l�8\�5+6������F6��kv>�3�|�M�>!w�(��6x��j�����G�[� ��V��RQ;�K?L���2=����g����w�0Q�ȅfqB \Ǒ=����w��Z[��+P27�×r.���AѥL|�f�ͣ�c�#If���td�J��/,4k����hH�SFf	""o�m�{����[7���O}������5'�<k�!7�`�� d�2K4� ��JG#�����0�-�7Ǐ��<8Rʿ�F-2-�$�������9���E�=ϒL����x�X�%�	�z�
�ԘF8��(���ڥZUVW8P.a��X9r���U��#����0����ƹQ���긥6~DYR^@� yE����fn�Q��!)%~����Z<���/זr�:Nd�4~�E-6�0�g��\E�h�g�O�s�|~�?����Y�ے���]]�!�*�~�J���Äq}�Ƕ1��U.�@���Ȍ��r"���/�x��G{�A܉���ČV��h��jt20���`tXh�i��G<o����r���O�M18�eGrT�"��Ə��l�#O<��u�6Q�~��6@���=9~"��ݾ�p�ܻ7S)�]3�Yej;���wk�E� �ܰMU�T����X�,8�ȱk��޺���s���m�~�6���0;�����	c�QTj(Tr%#H���:
U�������1i�y8C�����z�#��3���C-Ē"HK�֘ayk}J�i�������L�"U���4b'$����>5Ca��l�F���f/g�6}��D�@��[T�\k<����wճ���1���V����]^G�O�.x���㚓�ry9����h@%ն̉�fj��F�de��<~��+���
�~'�����g��0�ǁ:�q˷TvL�T\҂[A)w1�0ZUꐝ��j�Hlw�[)�4҈�%��#Z��>�Za��UG�;�^ a�+���F8{B�⎧[�ٟs�/W��U��K2��F��G'T֗� ����r�[����v������������2[�F�	5U+ʐ�/+g��Y�߱`�jٹ<�|����2`��څEo�lJ�~GS���^W:���^�����U�}/����g��]�'L��11Q3$TN���n�v����y"_�t_��.um%k�(ڛsԁ����+3�ܰv�DC���[,S�x
˴��4��U��*�L��[���l���DMUSW�^s/�<�ĉ������LA���ʼ�����������|�F@�J6�D��u��w�J��]�u�p��u�9��t�����k�H�p��� ��^������P��v��[��H��r;�J�3�n|LH�,U	FjLz��Wz��Z�Ǵw���gOx�n�v>��Ⱥz�zhfs�Iڊ�&��cl�3�4|9`���&�O=�,}7�-���6�[��ݥ��o��Tj|�񺱩KM�W�ݵ��B����:�E��߃��U�ƚ���$�f{������7�d:�p�E�cfn�U���UOe[uQ1oplTӯ^�?I$B�00 {]=���2���=�X�  �^��`;���[�z=�9mc���l�ó����Gn�v���ɋH�MI��O�6$wm�s���trhkd��BR�xg�Wg���Q�����]��ѐ��ܵS�t8��=bp#v@x��v�^��]ݗ�*�   *�p�*�T n��n��7v���@ S��B̸���,��
� �
� �x��xT�Gg]n�.�x*� c ���oaz���u-��x��sΔ.RQM�e��1���mUUE���-�B����X��@��/L���4�� U ݶ �UY��B�����P�fUE�PTP��l�� ��^�q�=��6U  �ں��J إS�k�dz�' cT�� ©8m��S͉�Y��d   	�   U  �P  �P[ �    �*U���mꉮ�isͅ&��j\:�KU),�R�v��r5cq���.�SKӱ3��@n�b#&���<`��-#ۇ��"ꛗ`Ѡ�]J��U�sXMr-���I����1�a��U�)�˳��i�B��h�灍@�eh�+V۝:���vP�]����T�   @     � 
�   �   X�        6�T��R�P       �UB�*P    � �͕l�    �   �    N   � b�  � �@��  ���   Skez�m�Y:�r���  �x 
� �@*�Ue      U� � ��l�Y�k!J�`cUP�����҅Sl-����TS�%�YA�{��8����ȯ5m��*���9���km�UU[Ӕ�Prstd�7m�J6θ�1P!*��ZR���<�:ґW�/e⮛f1�5�3h��ۿH[!Ul�wl���6���M�PNT� k�0�1�AF�R�n
^in��M��{ݡN��vu���P p�  P
�P �l�U�m��U���ov�6�EJ�aR��u ���;x���{�z��箔Ȩ�ԯ �J�)X��q���j�٥Z��8@��������sT5$Q���د	m֎�иz��H�6�o|(�r�di��\�����	nD�i%�(�O�ﾪF%ᓓ���|y�ڿ��,�M��C���zA�-� c2���,��4B?{��pp����E↲l�?�wPda�H�	����%n%!�|@Ҍ9���hx��7��9i�CJ8FT!"�M��O�c����5q$�E����=�������b�6D���uu����w����I�q�K�d���Bб��7V���h	sq���c��*��Q��weR�#��[���%nvjs�Rdnf|���.�U���(��m ��!g'.T�J5�(c�	�*��I�c�|�{9��������~���J+�b����"�t�G_ܗ˙���]�	3�T�2ey����h �Fyx��[��h�wi�#��'�5n�<@��J�G$���e�$II�}��.�Q|4W}_��<G|hϫ����O������r�d�����b$�M�Ji��t�6���#�~���S��@��g���C�h���_��KH�?�k_2�	
���8�A�k����n��Ź�R��*�*K�  �p+m��v0���w}�G���n`q�pW"���G��|��>�����P�0�>?�����2H�06�I���f"��w�bEG�7���wl�#
!2%����$�w�Hg��9S&a1�di0�U��#�l�8�}�$�����{��-\�ƴ�t�z �,�P(�8ᇻ��h�Q��$�+��G�d�a��l�g����Dk#��@C����l �#wu&�"-9$�����Il�@�x���#��G;~�v8��I�!����F��L}�Fv���շE۫Du�����@��Gp�Mn�:�2�w
���.`��U�P�W�$L$d��#��gG�S��ώ�ˠ(��#D�W��O���uh��EBBW��$S��D#��.��t��<ClfM���Ezh��S������rf3�^o��Ơ T�����8l�����w�a�c�wVJ���w��;��٩���^��Z�E�F���B8����|�Y�VP�;�}�U�+ 7)Ϸk-�����o�c���[m�L��>�rN�q������Bi!P����
ޫ�h��������ƩZ�����zl��n�¡UܶOU��n�{�%6��@35Q@�3Q�.�I�J��v)w�����ޗ=Yi��11���%8�m0�rX��,����]ExN,��I�q��̭�dqRG!*J�Wwbn)�����|Ϫ3H�ǡ8��u/�����&�L�2H�n$DD���֠d3�lߐe�|��yb�En�v��K����⑳rO��+��օ�Rde�V*��l%ٝD�vv?��=꬟<V+"^I!�Ȥ#mUuV�E�8U΍gȽS��v�y��K�H�R�.����/R`V��rӮ�!CV3r�;�� UU6k[WvP.�Wt�P	Yz������wZ;����9��;O:�R�J������kj���̽�r��   <
�  � VڀWP�w�6ùTUM� �[�b�� <aYJ���P�YW���~yn���ո!園a�V�-�몒�sbN*�]�UBjQ�@5�kڙ��NT�Jw[|�Pt���Ny�Q<h����˱�5�D�2&�N%��>wCU(��I�6�e��x��T�v	w���dz�︴I]��rH�����"
t���?I�6�?p�($s���&��F}>Sq#�k�0�H6�I&�L?�3&�ي��z�#������F\|�˄�E����Dr\�1j�T��ٖ�|��L�r3��v��G�>���f��
?*AȭJ~æ�cM�����{:[��2H5F�U�\��n�� ;�s��\�=�P;�S�d�UF1�/+S��Y����v����Cz����Ȍ=��W��ͨ�%�2��!#�"�T?��_�FN��~.6eH�ȳ�����9�ޏye�{���f��+Cj+ �n�'�]@�đ�3�0����{لa>�pDˣ"`��U@5SY�O�ME_�ٳ�Ca���1��ͦo�!+0�5�4��|���Q� �ȤJ����Nw3�[ڬ]����5�bj�YPdo��T��߷s9���b6$��db���s�dwU)����_Bk��_�p��d� ��
Z�I{c�"�Ab��+
����i@Ie�t��v�z�6B��jU	T���Ɔ35Q@ɉ�g*>DY\�E�,�p������DoJ"�ug�IDؾd�&n>�*U�V�&ZQ��x��"�~Gڤ<Z�"�VE��|jc�E�h_�Ņ3��=�^��R5�2l�(�����}$�}�צ�h�G�l����_>�:*NMc(�h�ɝ��(�6{��g�����^���	8ے�� �Pu*�#u~��0�ƾ�����E�ۯ���x4�M�����)��j�C���d�18ܑ) P9�AG䉷5�>���P�n�?q�̅}J�,��HI۾1q�p�� ��2(���k�;X'� 5��
�ܫ&PZUڠ	X r$D8{qړ�Wi�& Ċȍ�W#OãOiWǌ%C<�/����d�}�l���FcdƓ�I�Q6����1K�!?V�:`��E�3��<s��s���<E�i�_ȉb�|�O�Z��)�)��!'H��v��!Y�ͿD(��{"���LD#�I�3�5�'��B9NE33��bbIڪ���Ш��/��MMNw�f�2����w��_Ȍ(�f�M���p�����N�7�;G�.��ZX#��飑@�fh�q��2?{��F�:������b�D�8�b]QE7oՈ����7p�'e�3_M��{�`�(6Ԥky=���[�M��p��8���?X�Nz��-�����gPJ�ݖ�ǿ[�,�B�T���4k��6��~��i�O�fnOosM띟�5��k�C�,���Us5WbHN(�d&�ڽ�Ο����*���'|<u�#.	�{6Oǝ]ҏ�f�����
&X,V��[&r~�d�M[S�}[���k�������Y���5��Ͻߣ��jp�bL \��᫕G�ĸT,�����\��K�C&rpZQ���MZyjb`�2$D���F�3�7����Ĝ/"��|S�w�S��#
N�s�$�=�Zf��FE��$u:��w�ӹ%���"d�TV\XD���4q��B�8,��z�{(ϧ,�UTNm��2�=��S�Ol��D��+��;V�kV�b�U̬gX-���m�( ��� AY��㻺���P�tV����6k6����� Qrbۈ�*�Z� ;� +u� *� m�w�6�p �����gsnꙛh�T�A��K-ʕc$�͍`��7�;e��#�#`��ۮ�+u���«�U�	�U*�T���#!�( f8����/�#_q�~#�G�é�q��<{���WeeI���؂�����0ab��,��7�����_���3���_ȋ<Ym���"͝���g1y��wYg&Y�w�*��,A�T�5"�G�B8y���3�6�7�lQ	şUH�[�h����)�=V �o��ڌ�1�.�iI������ז%3G^I�r���)�#��Bf�M[s��$�BwT�����W�E"&F�r2S5�Ty��ӣ�8��$��c�ÛQ�bI����cg�d�?�V8��gU&,v�7�f��\�m�սzw�V�`x%V��	(=U�d���$m��E8~�9Ç
���㻝����Ҍ,�޿X�V� �!5��7�fjw���H]AmUR�8y�����%�Q"��-�p}|	��"�����?K��~�y4���31�K��U���vry5��۩m����
����=oO�� ���l�h��G+g�d"4�uk�Q��O��U�������L��M����CN���in�{�߸��1��ע	P�FD�X���qӎ��,����7�lQ	ş��[E�Q�����31Fb"����e'lM��U��c�C"����G�G������H�����LLF��ݢ5���n��\ίo˽�Y@8≪�jR�5�.NnL�)X�󼿙�n�w���N��/5s���G�"�h��(�����43�^��O��y�ԑV��6̃��s�T�V2A;զ:>�Uc=���3	Y�i(���G�p�3�8�i�&$LD7P�T�B��~ev�������Dx�&����B0�o�Y�f&3/4���������vyU���̺�����a�t�s�7K��V����=�d{P�>��3�e��G�=��t��7}�wW�v@�fnL߫{�f�?��0��T`G�(��i��8Y��Q��Kq�&bvM�P�%Mr{3���9�;���L�gc6�u0�d���#dMA9Г}|n���,�﨤��)@����)�(Rn(ސ��j��yk�:�����Y��K3V���#��c~��^�2�Ѵ�8U�.�
XrYny��r�T�����j�;�[^��wPD�)Ě������5�Z{�B�f��B��W�+c�ElBo��B�G��~�,�u}R �0O�H#m�1UVN�h�B�sJ��Dd��6��![����&����t��>�/��bFZ�W&��y}�����s;���̆h��0m�#�员�F\�2/9}2��;����<����0V�e����	�O���8�w�n�o�lQ��0��WY�'�MJ�ML@���d�Z��0���3L�!�erzh�VK+Y+$$��~��N������1q�>��K�)��w���%YeQ���*�e�?|�s4N�@�K�^�=��Ɓ�UI 
ݮڮ�n�Ү�U	V^P�ë����(L*�ƚ�CQ��2�ߦ�FD|��Bd{"��d�����U�-�Q�	`�w3����<ﺖ���ѵVۀ������
�!�J>������t2��X������]Z3��#��`��5U��31d͆d�t���ѿ�Q�қ$igҷk���rδ4�=D�9ڿQ7<�=�k
�V�WO3s��{9�k�Hf͝0Bߪ�ˏ��q�_3��c�-p*�dYdK�E���1D�ETQ�1W#n��h�6�m��/�(8��1��:V?IX��=�LS�����%�=��l����U\�1���Ë�p�-��e��6���n�˻� W���zWu�ۚ�*�v0�Y]�Y�#[�[;���v��&���4F��cRv�k��6��UI� T�k�]Y��x%q�/H��SW�#!q�e�U*P 
� P w;��`U� UU@gV�mQT m�
�Q���ꆫ�z��W\��.��h	q#�4ݢ�p�M:*�ݳs�eWt�Y�5J�Z���$L j����o����<<)3W�����s��d��G�S]���S�w��K(6L.8��qY��WbȲ�,�з� ����9���qx#�d�����km�mY��ܙ�ɛ�yz���i[t��0����G�t�{;�ǎve��{ý������\��fn���,�t�"��:ű{G⛳5�I���F|���~�#L7��Y��� �B�)Ib)��<rDA�Kɦ��>(�t���0��e�ag�Y	Ɵ��H��Q�"4���5�����m9�4�W[UA�\m��@:�R��4�Ke]HK���ꓟ��&�p�a��|G:6w�J���X`�Hd;�3锧�!�C����摳=�֯���#;=�k}�m�Cd�Flz"�<V&�I�f��PY��y�_�վ�"=�9<3_Q\M'Q�3��ѹ���v@�dīj�̲��a��J~�:�i��d��yG�}��_+j6������;l��ܝLT�����!<�ח��}�s������i�Y�#
8R�F�'G��>ws���Ͷ}�w�A�[�g��7�>�.��2;"�y;C6CdG<n�N���G�:bk��Q���,��k�jCڼ��"ӂ��cj��onB�ª�Un�m���x���@�mG)��l��;���_�ý�4S�M#���KS��r0���]+�C�b�9�qD[�TQBTj��*�,����yBק�폸�lc6x� q���D��#q�hl:p��q��$F�I�@��d���:����jLy�r6z�a�ͣ�/���^�g�����w��]�{��޹.�m�[2j��r��9ʧ���f�=�4����=���̞r�8cxߢ"�����51U���|���}b���"[�w^�q��Q�C�ɑZ�3���p5h3���کg��=��v�m�Y w׳ ĩ��	�<�AG;�,�f��V�����M�J�[��X��%۬�h��@ј�5S3TЬ�#��1�z���W�4�|]&�lS~�vl�����b"f�T���"Ե����,��Ks���!�u~H���֎΂�bl�z�I�Ț�1F�j���v�p�{	�y�}e�֫V�2����z��z�����v_��}�����w�y�vJa��h>�݉v�9YMVx/a��e���{Y����^&n��S���V-�*����3myT
l7uz�B����wM���+�U<P�*�7-B"䬌l��Z^y�5�K�m�cm�a�j�g"��[�V§�7��뾜�M�q�}Xs�}9	�
j� ���V����u��l��=�K�7���!�;���x$Zm��M&�n���;��Hߕ�#����F�+|8�����G��H�~5#�켿|�����	W&1 
�<�{b�n'��z��#JdҚ�9�,��An�Ƹ�3�4w��·�G,�jY�w_"1�X�J�眚���GLkb�P�!:��T_Ȍ(℆è!�-��|]!���c "0�Wn$O�i�SC�U�
2H�*�an�l< ��k�R�[z�6�X�vX�,��*�����T��@2���H�Z�0P-�V�0&�e���R�X�v2T�T@����J� *�
\�'3l��5vi��z�{!�ڵ� @Z�pi�g��*���@ 6� UP6���`U�  m�@���AT���mfUyvN�j2Q�w^�Y{6�r$�x[���UAWU9�ҁw7bQY]�UyZT6�$ҐΚqV� ��f��a�ᆔPDK�W�K|�b���8b�-�ڸAN㟉g�ib�Z$�om;Ο�%d�2C(�y��=�ҙ�sd�d�i�Eq��2U�Zq��-�i���Q�k��˸��KV5PS��<��&vy;3ɝ�Ǿ��.>�0nEq�,�#�q��2<鯖��1}��^K~_���<P󄲨��Ɋ����3�~a���k;������,i���U�ߞآ�Ǝ�}r��/�E����f�A"�ȴKd3�	�o�{��Tx�`�S��؊6���7�
��!
|a��rۏ�#�/��Ç�9��F$S�F���:�4�$Y5mU�T\��k��wW� ��T��l��XV*�\M�y9=�f׬A�n,;~�h���܏3u�{��#	ȹ+F����<� lť�l��$����&���'{{3����m�dxQ�UՓ�fk��#OpA�Ց�~��ŚQA�%�@���$�fdjf��p��icm
����s5:�1��C,�����E�l�qbߦ��S�?9�M#$",�\fA�LH��h�u��x�����L�ه�
����ző��p0�ȧ鲢�<B1�Na���S�4�՘�}��y$���Rfh�L�120�����N0�x�Lşc͑��D�M7a��x�,�rk��?����.R1ʿ�C�L�JK���FRq����!aU�lQ]�UW�6
$-�%��S�_<�3��Ϧj"�V��#["7ѩ�o�e"i�*di��G���"��.���}����Q��,�޹NL�y���z���r�x�x�Ta�QU�2��,�dx���뎷��2~�g��qM��%��R$�G�1��<GՎ�w�gR��G��6��c���^�6�W�6O\,��~��҂�M��C8j��"*(�LLLH���E�Y��s�%��O������tnG�F���dI���vM�Ty��ܞ�Oc�s]�2
�[?j��'G�N�����H�L��V6x�Y�2�ƔDE�<9�Q�Dy2o�.SԀ����m�J`�p�E�V`*��8��j��UN�0ffOmu���+m �$�Mw��k3�=�3^�D2<�
����+�C�2x��_���*�q��qg�w�e���d�[Va�g���������g`s�U@��X�E�NG��<�N\q����y٩�����;��\��%hA4k>da{J
�l���wO�yFM�)1�命X׵~q���z!��7G�噽7"��7	nF��"0��bda������@�yHd3������B"̨�Jݢ�d�fqȽPZ�Di�z�Y��yBa��F]"�hZ%��GĔ~����"�F��G��6yzC�ΰHf�#-{V����3�{������8�(	m0�[S�â��m�ʩ�@*�f@wn��˻$�e��+H��\L���ϡЅ�5�"0���{&��eR�iz�W)�$�)�ەmG�B:m-���b& 8�jD"P��!�V�q�@�᪏�\il��qx#���l=�Em�����U���E�D��EĒL�pC6[������l�(�˅9�}g��g���2N��fӛ+��C793S>޻��j
�`5k.
�Vx|��L�M�Hc0��ƋS�����¦�I�ܩ���E�Z�o�qW���em���Q<�o�'ggӽcƂ,��肟�(Q��<Yo�٬��Pgn+�D&#N�����������fb4���S7��L��*]��[3I�[�!��l�3J� �ܑhXkٚ׽u�t)�|nP̯d��J���)�
�s�W���,ح��W��y36�ߔ�]Ͻ�y=3A�
�H��QUx-ty��iX(p��ԕ� �Uw,J��JX��M�{Pb(x��-���`1jUUHx�'�ϛ�g��A���#��糆B�u����:�^zv�z�
B�K�jɺ�Ol���up6�lm��l�6�eMa�P�͎9k��M��8�R7c/]��Uv#� T��*�T�l��w��L6�ݰ6��TT��{sfJYOl��wP��S`�P=���n��l	� �U�� <  1�p�U �^�͊�׭���&�q\�	4�ӎ������+l��w�v��Վ�z�' c%)An2�PVURUZ��4f�
�<��{�M��@�ATT� ;��T
��-��m�T6��n[� U �m����uK��5��:�-��^�' *��S�*^��9��
�cd�    <    �T  ��    �����/bІ�RE(8�il�PΑ� TЕFI��1�r÷N���UYʌ9��ݷIJ���f�#�AM�ka۫mC/����'���b8��T��Ywb:�T񭥕�tDc�J8��V��Z�U�p=��I��[K�Q/E��b�Td%�t�� �\�^ߞw/=��     
�   T
��    .�
�   
�   UTU�AT  U        �@*�*�      ��l�v��  +&�  U�       �@�     �  T�  �  *�   m���ֶ���^*F�f�U  P `�V�P        
� �5@�l*�As ���UEJgZ�  ��'z��%Kd v�v@*����eu��w�z
�����{[wi���Q�L �
�j�ɣI�\۷^guk�K���^n�+�z�*��\ùws�\ǁ��5?T�f:�y�(qvrj��(Ɗ�Ҩ�({�UO6�shomm�p0)V�W�}��8r )�V��f���&ǋ)�vK�qm�מ�U��T�  T��@  U�^���]�� U�UU��l]���*���Z��*��,���H�=Z.��X�� 
�U�U.x�Y�l�Sw`�q�<��@U�xT��(dT�����w����f����~�'��E���Ě#
��8�p#Hs�8���QJ��e�Q2 ��ȏ�c3����=��b�x���G�F�?[)�
!P����q�|t��N�N*j��y�Qg�8�e����$Uܮ��,���}r���Δ�4��.2x�9�m
!�,�CDO�����H�4�����(BE��|�/v.n�i�q|�iHl:��8ҩ�}�*7�}�ٍ�Hy���C&{3��o�ƃmfƍ��E�x�B;���k�O��is�2����ʏ�{�����e��tw>D{9���/�wvd��	dmFU��ɱ+��j�I��N�iWj�UiP �H�y�Um�
24�d ��ɝ���g�i�E���?mf'_q�G�n8��*ab����D"�8�F
O<$B@l�-�h��#������v}<Q�|�Y[0�^b���͊7��9��Hl;�K7��}�:N۶M�!�~���ށZ\l*��̃|�o�L��K��(���آ��BB�U�ʏ��<����E���Q"���)4Q)Ƚ���g����+����q?x���5f�D_�~ھN~�a��'�E5���[��I�!0�$m�fL�C4Y|KD[��#{"5�0t�\`2CYoHdfGX�<�è9ٝ������e&G
�$m�K��Ԅv�,�����Nh�u��UY�~2��q�Ym��|�<���s���P�� �C����=�t�=*݉8��,��,cʱ���>��d����K<{sɝ�=�ܗ��_�7�k�|X�9�D8G�b�FTFzz�Ӄ;���x�nIʡ3bj"��"��I�ώ{�.��f�!��4�oƲ&gK^�,�g�>>8,�,�t�Y��|Eyi�[�$��IC��DM�#������;f����S���y�G��#/�BZ�$x�n��ؚI�D P[�_0����{n��C'x!�hBu�_��}�!U�Q�㺑B޹بx�E�?'�P8��urlF�'�����{�z�h��x*��2����[�md��:��ێ"�ٍ)�񠈢�ԡУ��#�V�\[���,��Q�3"nf&jb�"�fH�U:{���{��b�4s��=��-����Nٻ���ȜI�NG(�I�=�G�Ƭj�����3p!���cw���S���ڭE��#N\����x������>/��Y�H�MVq�A�T�`���C���57=�g֖=Ԏ��Ofwod	omB8h6e��#�((c����3��Lz/ �F(�W|2�ʎ��=0�Ȕ����>����߭������n��<��¥�8v�z��n�]~���UF�K+��.U�	m�Qa��Dn��!�G�����#�"0�Xڱuq����S۽bϏ�û2�ixݭ����(�Q���S6H�<��������4D�e{��}�ŝ)�i��Q�!Pr�������1��L�b�[Z̢y�ٝ���1�G�u�q
�}�3�q�C���q���+f��.ᆽ�dL����JC���y~���!,�Cq�r�g�(�#�5�a�̑�sd_=BE^�ۜ�j*��䀠%�m���i��Ή�8H�3�,���QD:>�z���g��>Vh
�PyN}��$�����k�珞�d����?+n��vGr^�Ilͻy��u���l�]��BqM��������߰�m�.��1���
�ܠ$K*�*�JK,8��H�8   �7f��3	�u�olɶv�M+�ۭ٪�Y�m��  �   � � �.�6��`�iT]�޺��*�� ĭ��*�<�ci����{e�;�3F�Lͫ�u�s�Wm;A�na�{��j��Uk5R�T���e�J�J��" >"[��Yx���<||'���8����y}_�>�ܴ�"��%���$J6�Iю�0?����n��iѤ ��"K^�bQ@�wF�E�����{�B�e�
�\	s[�~���s<�+�i�����?i۳H�e����M������C\��͠����@SP����������C?GF��4yŋ��8����0��~��W3tu1��wȰ�"3陨���"'͹G]ŻF��-
�J>����^@�k�~y�w�m�~�F�ՙ�;i�z���յ#$c�N��2үP�J��eVW;c:�s�I4*)i�$�Q~����d"�
�Q��E��<)����q�q��^��&߾�8��h�*��_[���(�L�խS���w34a��~<������qa��7K�q��~�,��+Jퟤ�}�yur�U� PMg&{3��C����i�Y\h�q�xtOt}G��� ��������QG�����A�&�?�7uxr�~���	��f����p�#��:���Cu~���G�m��H�J9~�E�w�w�.#O�(z���AdR��.YO<Gq\��g�#O�nr�|~�M�
P�v���A���$�Cg�XM�/�6�Vʪ�1Y��dJŷ,F�K$V\?�O��2��(����1�S94HNnh��%
��]���>!�>����._|��H���RH��!�7hvߺ�"bGH�w�i�_��ա�20�W���U��O�w���wD���� d��B��}�sܦ�DaC��_8�N����fp�ӽJj"�C7g����-���NL���{�~�H�ڥ�,�2��7'�2.����J0�]�o�#�3E/�#��_1�M�>�i���m �"I��!���x�G!8hߢ=�]�$���;�<��y���������I�n��
օ�&f���9p�5mU%��F]��W�� wVdU�։Ϧ��m 4����{�x�ɮ1�7���3s`'���h��Q>���6F��Mx�t�B
7%�P���pB��$�FAGO��0��{�u�W�����gQ��_)�en����,��co��a!q��q)h'.�=��r��Jg���˶�.�m{]U~]�{|q��`��o{�������tǂ��)NTR���^3��:�}�Β�U�~7%f/�F�:�� �mĤ���5lx��:�=r9����$Y�N�Dk�����dx�q��{=o�!��_�9��BYV"�2 �qZ�2l5�q�pT��T�>�諭[*��v�Sd(������,�-�h�/��%���6�q{��<��!(e��adVB/����)��#gp(��$y'�(TIX}K�8~s��z?�"�ìӣ",�/��$#G���2�B��w�8�ٜn2�Q����9+�_��CShx�3�FFr�!8%00���|�K���^�s�rE����-���,�bm�An(k���+[��i��H���'O��(�>����e��Ļ���������-P3���C<YCtq�񺏸�r�����~�p1k��#���l�(�J �#-���>Jo�?�\��شd���'��z�i=y�u���5Oe�\�6� ���v����;�uQ��=���gjݏ�o�������b0 4�R�k�z�U�wl�T)�hJ�2�MRx��@����3�iM�B�{c����޷���/k���   �  *� UP�����x Sl�����l 6�P�-�U�#]l<���˸+���]�)���+�d��m�*�����W�P�iP�R"]��S��u	!Tfb*��6Ge���#؜}��a��Y�Ftǲ�1p�da�U~3�������iG��m�q�dq�ýQ��0�>#KV�O�f�7<G��C�l�{G ���!U�D�[H��j�O�l"$��o�
o�bH`�E��>�V�����]8'��#�=�θ�ٞ�d�w�{�hFL���⇒g}�-����X�P沭8��d(K�".o��A냋<F�0�޻�2�"!�$�B���/�Gֻ��:Qj~���M���Q�AHl����}d=�/�"0�%�6	���(�eHKR*�U�ӠTV�Xƪ���崥S�V�Hl��U���ڳ�Ϲ�?@��	��2$�	F�k�Đ�d[b�V�������I%뚪������Q�$�N��0u�h��g����t5���>:��,��o���Oxy���V�x��t��J�J������c���y=7��}����,J��>
�����_{�2��m10��8�&(�!E�J�?a�T��<{�Jo� �N=�`�"�*�r��#����&2�*ڪ�r�S�N��/${�|���@�
�l�p;3����~ܚ�s8cy�{�v���l�:��Z���j�]t�[+u���a���۱]¦2*���f*
X䠓��k�;����A������s�y�ޗ����sU�����I�D�iĒl(d�s�7�s)wWW��!05���k�˻{����w{��M�CN)('&���B8'�ض��� �t��e<;��ym?/m핛�yd�V��y�����nl�vr��zO6����Bk�q�3+5_����g!����0�B���צ�-�ͦ���+Z���z�!w�-��Ӓ���Ʈ���n#Ƅ̘Ș5A�"JF�W|����?q�)�Q�ֆiܤB6Q��-U��G�/�a#�w˻2h-��C ��g&3z���쳁�3�4�Y�l�f�#�8y
#���q��W���!1�`D���5��ͮ����T��L;s�M*�R��Ҫ��T�C�T����UM]�gN���r1�Z�܀������(����Q��lBjE�*(�s���z�
VJ�Q�2�����v��*�s��3%�����fs3�闉���'��2'�RI��Q��?In���E�֥'%�����!�����yۛ�|�{�s�d��$�"O��U��\��e�㹥S�G��B���j�q��n�V�M�(�ǖ��QFf����-�Ў1��f�B��sM"�8y{j�l�,��R�cƥ@�͸�]���ML��^]���b�r*2m��u���4cU!�T�[jU;��d_�;��%�
�:%.T��k����?g��i�,�QxRށVQ΄���7J���"�v͞P0�o�5U"�T�&���w�Q7��/���q;}����CL�*��l�Ξ:�q�|s�N��jX��cY+%�+Fǈ��x�jEd�R<l��4��!�c>�J�B��g��)�QӶ�U��(�$d-)M4ԔG{����Q��@Di_a�8d�p�Tw��"(��C���٩;<������u𥅶逶*�Q���貈�H8�̜!�8��-�Fw QG����$3e�!��*��@�/�]�wE���/:�_EI( &5���rQ�;$���,�z惧���ң�KUP%�����ܲ<�皡^���݌=zv����z�ӝ�[�*J��]s�*�)*ڌ(��+\��� @���K��Ĝ�!��k����.u�,�m��d�UUU �T �� ��Wu���A�j��UT��T�*�@�*�e%��m��]���\���k�lJR��s��RsM�\�;����ۘUw
���Z��� �B�)8($IF�pD>��IՑ
�ب|G�{��R�L���S�j=ʝ���^ʮ����/�jD�nDP֑G����s��`�j0�Μqh�nx�; ��bx(��(_T�D\w��K�G�P�?"$,��nh�/��Ͼ�h�0���aچ\쿰�8Q������>�l��L޻ܖ�@!F�
0*j��m�2�x�b�$[�}T�jo���	�L�fyN;�y�m��ㄝ뼖��,+����������R6In5Ǐg�]�.�/���qj���7��{[u#�J�1���ERdK���A��G�����R�T��
�
��Ī�BO֍��3 7��g]9��|��=��9	�ҟ�W~��{��z�DDA��5j!���v��lc�n��ތ��5z��,���̐�+�-��#�y;O���P�)Ew,#�pl?R&5(9#��|����}s<s�<��Q�H����Z�[��z����n�7����	��@$b�'��������"������а�Q�G�j,�T�~�!>�G����"(�H�!F~���(��i��f�9��BVճY��BءӤ��&ٕ���&��ľQ3䝦0�n�vG:�h���Wz��Z�ƀ�*ʀ��W:
]��ޗ��qX��r�7�SK:~>K���-���7a#�*n�F@�s������t��b�m��$D�sZ��fla�c��p�B��V���]F�	��t2��|]���0����4�m��jH��$L}	l�Q���F�"�7Ƃq��"��������"�^ʴk!�O�yk�997�}�1#�h���U�x���Fj�K弰���M��Ȳ���_(���J4�G��<��d��ㄩS.U}_W���=�`�2Gc!v�}5�u���������Ůr*�N���"���U[�nv"�	��Wj�z�d�PUUwo3W��P���"b���e��3gÏ��q�S!��A�,�	YY��G<vu�aA�H�+�?���O�ʾXp����yAŝ�f�k�Y�(���e��k�~p�N��M\,�-������l��϶B��>�%�"��jo��p#N��#O�K������]������������^�}3O3]��ˋP<RVŐ�2��9��$��0ڱS+��~�%�Q��������m�N%#)%|}K���
K#N����F�t�0ۊ��Y��)P�Ȟ}���%rJ�"�RИ�.�٬�Ykm���i�����P�2����F�T�m|�{O�t�O�߽3�"�+`x;�a5jd�_)^��k!(;��g^�3����t�]Pr�e���QV�&�)Q~�~,�N4��-�4Q{��)E��+�Јʎ;�8���>�"���MT�0�ƈ��J��^���D	�&�p�B���!��PE��dw���~@��NI

GZY�U��g���_(^��q�q�H��(���㥺c�o��O�ψ���[�"h�d5$I�����EZP-�>8�����Qdy�V���|�6��lp�m�����<Ϟ�2��8�b̒*��K̜�g���r��2��=�oݷ����� �ZR��G���]�T�e[��N1�����Z��*Y��E��m��w`��2�  �6�Tkz�E�������6;�~_�8�w��OwS�@  �  U  �P sp6�Ta� T� p�����@U ;��T��Ꚃ�k�n�ў�ID��V�,E�k�Ihx�1��S��hΞ��iV�T6��r$�5jn�L[Z(dГ����D��A<��f�8�;Р�0�v7}i�gM��;�P��\"������Nr�3ǽ����k�W	j�SZ�/m��s���t&h8$m�\�5!9�S*ǈ���rL�����S�|�l�s���qI$��UDD�ё0;�n}�?F澾EKE�j�|��˛������$�
���U{�ha�_��:w��SH���{�Ǐ="� Ñ�i�A�F�%˷H��.�1��ړk:��T���U�R����T�*����C��T��������Q�������a�G��&�����[P4��q꿤�x�zd��)�f2[j(Ԓ���/u`�l0�XT3�9���1�;y����}��v:֝�g���n2z���-C�@��xJ�<p��FlQkvY޹�g�y�8��>!(�nq�ɣ�L�Q���"��ǎ\Q�/]�k͑/#�.���t(�n���H�O��oȅq�Ì���ߙ�Tpꋼk�?����Y���>G�=��+.����]~�nL��,	�TWm�b�N�s��]��U�6�*���[Ӛ�ݶ�F� m@e�>v^���s<���Gxd%�@�dWEg� �J<D�rY���>��%� b�pE�{����lϋ,��3�v8�G|E-�3�O��p�1�x A�&�-XIpmēP����!G���\���Dd;���+.]m��yy�.l���mf�ԓ~��Ñ]%C�\�}���;��E�A�g��wlʚ���Z�ޭs�;k�o��7`a��ي�ȭ֡73�����ӌ#�y����\~�]��+l�:�K��(��(��,�ڐ�#m�Ñ�=7=m�
E��m�:��j�5*�H5T���Z��F ����6c3[��p�lk��Q�(���,3e8d&~�U>H�f��'��q�'o��%��q�����Cw���eZ.�+����5�t��&m�_��ݵţ
%��ڥ��9��������{�700�O�V��:��ƚ��w�OL�W{�s{.5-ĔQ�[nF�
�W�$����(x�4ph��+�
9�k�+O�;�^1 �B��W�3Dc��q��x���D�m�R%#����Q.<_��"N���
Ti�4Q���j��ܯ��l�!J܎Ǝ�K���ܰ�S�Wj�S4p<����T��*Ԅ�[�U�9 ̳OXj$JD�)ȼ(���M}ʇy@��z����/���m]���>-�i�s�o&�w���w�Y*'���v"G�g[������/�a��[�qW�8h�m.����N�;�ɖ�M�RI5U��7�ψ��I�̳o�e�#c�L=t�8Y�r�����6O��$R6��!\Y5���ՑW�6h��5A����vy�4p�+:'e��j�Ԭ�{��@Tq� j)1C��8r��5s�:Y�m���+��!Y�,ѱc*�0���w���w��d�p�9	�ma�x��3V���~Q��*8,�̙�k<��'-_�ؼ��
Dx����,�,'K޹��uY��<���*����o����o*�_�n��z1{���{�U���UUUW�ǵ�Cu <6��J��  ��SU]X^��&�r��8nY,�q����5q�j��c��fZv9�{>-��v'u�6�#n��D�G�*ز��r+��F�n9�r�k�d�|��{[iʍ(��nT=w`�M�����;���/Y��3�6�5ml�� �
�ͪ*�YB�����kdU6  �Hwm��c^�wjT�l�J��!^���j�m�-��uj��¨  �T�P+:b�5ԧ��Ӄ�}�����׷�T���V]Ԯi�Q�[5K�rǻ�P^�����<�UUT[`�-�F� ��Cw^`,�T���*�J���T̸&�P w �=v�ջ�eP۵���^ {�>��^��Ɍ��   ��8@ 	�4M� <�5�0     �T � )�  �@
��SJ��s*��%T�ʜUJ�PT*�s#!;R����@9�X���� a� 4(�[S�/�,v���1m ���N{x�;�v8���H�CEǇ�_�~�Ը�)gs&a22�[�����ggf��t��i�c���\[3�\�ٶaıĀT�������[{�����6ټ�(    ��     ���T   ��P @  T   U B�   ��    P U*�JT  @    xn�AT=�N[   �    w    �  �PU�    
� ��  8@ -�    6�p@V
��ڲ��*ƪ � U  �l
� �@      �  <U m�  P P��WtNC���N��B�-�*횀:���)T{x��n�JV䖫m��Q�\f�iڵ[%ųB��:�]�q�Y:+k��v� �w�.u�j�����
BeB	l�s�x;�wUQ��Re�g�d8-ݬ������Vgu*��mU�<6EPM��+��)�/-@�&݁8y��d�ó}}�gn�l(j���ր     -�  J��W���6�� U�m��U��;�T��
���� V�wLY�G�}u�i�P-�
��rpYBcj�v�`��`��M�
���[w:�iZ�p0�C(��籛�O��O�M#�`��� <w��Z�(��Cw�~gK"����I2c.)!9+�������i3l�9�f�0�x��D��Cd��aȒ,�ܕ��V$u��E���W?2��O{L�b��U�8Q�����S	H��$$�e�(|F���wn��P�Ty��*N�>8E���=�޽��Qlݭ���v�FGQ��:������ޕ�y~������G�	�e��`�T��߯�ϻ�{���%FX�2-���K�nt
�-�ѕ�D�����]ª�U\�EV�4e��	Q7�����һW�h��0�ky�Y"�f��#��u�ԇ���.�H�FbBD�ocG1�U�w�˱H����G�ͥ�P������g4ryt���n��'l�	H�i@����v�{���h�7w�q�-hx�A�ςZ��*��>?g��2D����ۄ$��������|�x�<7oһ�'��tTfG�����t�3v���"T(d�#�' �>���Z<Bäq��c�*���`���J>�2�֙K��x�氦1 Q�aL���jp�������u�
�����V�UU[Z�Q�*
� eɅ����O�|�"$��C+�PN,ɢYW�^��ٻ���o�oZjѶQ���̸�q��DZ�
�f�(an�G�������?}��-5�>Y��$r@�H����ԃ�<}�;Mv1Z}K�B��7�C:���wW��,\=jT",�N]0�/�ލ6�M�HKrӂ�Æ�{!��/�x��(��9���lh��C8v\g.�r��6�}a�d��p!\Y|{|�s48|pi��ߔ;��G4�ZE�;����y�
��V!`����ɑ"�j��%��ڢ� �;��wkm]©�*��/w��A�č �k�I�{l�����x��0�7�b���^!a�4l<����/�P@J-E�����>f%��ˬ(�)��%c���.s��gb����>>"���L��[m�r������~ϳw0�>9�J���gGW1{�[C�g�5o�e�L��T/������af��f���L/R-���ج>��n���C��֌�K�<8�d��C��zX1Q��rY�O���Y�k���ü�h%��5��G4/���<w�����-�V�"�I�g0��h���Uc�(��os=��v
��Ul���2�̰Kn|��~*�?q�f�=ޕ�Ԁ�����ӧp�V�L������,�&�m�hH�q��a(�8G��r��п.H����(��!�o���t��m��a̶�޴�$�Q5M�۟���q����X(GJWp�XF��?%i�6|E�y>���<fz��!&��������r�C����0�����>��n��F�p��a�j�>=]\_�"4��b�&R����%���]�ng��1�ھp6R��^Y��@�7��<h�����癯;�{�B¬�"�����W�d�v�:�pWn�Xss��s�yz� �Y�m��]ж婘���*�k`(�0�YL^���+k
�F�n*����Y��P@ � {����YU��keJV�:��,�k����oomy� U �U d T[ ����6�mT� +m@[pU
��R��B��ʄ~�����S5���H�I	臷NW3KR��ӳ����*��UV�\�x�Unun��-�NH;տ�����#ME�C�I@C��3�_�VL�R0�����5�H�9�~�B�d�
�)d�]�ⴿ�W�E��7�'�(���]=w���3ss߷@�[h���p���5A�3y���ae����[+�~������"���ϕ�/�H܊�&))����O�^>=��1\g�{�g�GC쎀g�����(Y�.���DX2F�`�J�!	�\e-0�|�f�Ǐ��b�zC3dI���U|�k�#�{}+������D�A۠���mQC��EDd.����UJ�*ڦ�A���ּ�=��V�[�G{�#��i>����x���j�ڡ�@M~�EU�"��r�s�YR���
�6g梅��>�tա����WS;ts�j��o5٣�Oq�9Ʋ ��ȍ>#Ɓ�SE�g�RӇ��)5�bM�S�$�qH(}J�܀ZY�4p�84r}��(%$q�D�=�9j��(���ET��լ�+��^꟟8�M�yp�daӘO���(����5�������<�igH�պd7�	H��������l�����(��K4��٪�0��6ج3������B|Uiհ�T �6V��r�T"i�-���͡�l˸U[ *	�@��F���8)$��h��_AC�/y�gD�f���A�y>�=��|C8fc���*��������������sOu������ő�R��SC�!��L����L�ͯ4��$�@�cM���J8'�n guk�\��|T��؈}py�;�f�x���7L�c<O�G+��8�$#$(?�� �tt>�bP�H�Υ�W�sP�5���\�9˙��<��C. ��$�?x��劾F=�K��^�ˏ��pAߐ�Cc4:>$M�Ew"H�Ь�I���\�*B�h[�ݕ�owwc��UUmR2�dc6n�j��� ���;h��� Xޮ�ڿ�*�5\��=�;b�����K,M�&�A�j"�q�yF�����x���bP��]�ҿ3���^�9����@�[�"��̄�|�Oۛ�㉁gֆf��\����Pu��R�< a��i������Ě1D��g��Z���������e�,oWJ�@i����d���.�����|�Ϫو��RF�mԑJ��a�����3�
J�QVE��CV� �a�y��W�E���j�ￜ�^����*p��=Yf���i6M�;#����-��U��M��]���!-��AH}�Dz���g?=L>�/{��rC�݌����{y@A�#��#�[(V�<w	��W���9��9�����e�d�ޕ�����*�!�!!�M&�Q3@Y�To�j��ٞ��2�o�.:'+�{�1��2���4sw��q��
9�"��3�3`�8֚ X���0��"���w�:|Y��$��L4�n"�	��N��!��0X��6��az30�m��eg�����qԏɒ9M�n�UuP���/��ۃ��qV�8+v�su�p����/s��v���6U[��]��Z���qs�)�����,
���ɱ2�5�A��� k��P  U���ww^����h.�R��%Fs�K�u���5W��  R�@@M� � <x w�6�l  
� W�l� � w
�����K^��6h2�[�)1v���f��a�k#;,jn��X[vvjUڤ� 6�J���9�ˬ�!���A�%�����9�34�]m�+���ۼ����n�m�^�I�ل7#&_�=�].�Z��Vp?���C$*�����A�IԒ!�*���
wEWW�P�j�lMe�?k�s36{�����`*�g�g6����k|n����6����犣�)+odTET���R3#������畘ξ/wpt�:����3�y���VZ�&���<��)eѶF~�-y�@
��@�UR�L�/NY{��o��\�dgl<��+0^������qO�PO�H��$�&���|�7E����L_zL��|�f��^q���[��m�P(EI6�f5����^7�x}s�w�i�E߷�}���t��ې��)���g�����MǸ��杒��<��lJ&8KY58�P�و׏��z�2͟�;6�iH�+O�{<���y�`X��%�����j� ��i�U���l�*������	�;r*�bp$�%&���W�#6w�yL�������`�d�?��Qނ�!E/6$�a��$�-ęq��4!���Or��l�!�����:~�0�CpW���� �6���(\2H�l��UŐ��f��(�7�1?��~�x�w3�=v�9��ۯXJ�Zj����l�m䔲�Qsuf7�]�e��8����j������U�e{�c�w���Xd�Fj�����Ю��${���S��7�k=(�>����|`�ꕄ#��-�m�������?�ʉ8:�������e)g���p�9j�U��g"�)'IH�e�k�8@�8P��8@�/e����;kg�#��w�L{N��M��ْ�@e��8�6�N�iWU*��.��S%��;$`�'���g��_��[r���ى�1QY��� ư�C�46�i�a���NJ����3��M�f�~�0�7��,���������QݽD����
��`�~�a=�s�s���|^��ׄ�x@�/������̮%��oѶ�F�7'�#4�C����Dwt'e�E��w}(
"奵.�FY�b~8N���?�. {�
lj6S)��JPF���R�����Te��a�������2��\��n��hƊ.	W[7\�/)���L��t�e�r��*Sd����"�sP����.��GC��(D7xu���p=�F"l���S���f��M��RH��"֟�|Iͮ��!��'���x,�����snU�~ �o��!#i�LM(Lm��5@�p�{6|xn�J���#5�g��E��p��#;��\�F	�j"����=6x��Xx�gG�Mʳ��B��5�%�9~�5Th]+?�wSMFDF"d�&�(�Z@�3Hf|~Çr^����}���,�p��"~�oZܷT�G�}w�_��n)H�z�r���[j�v�f�궺9��d�z�9���b�MHwaT�B��͞Zځk]��8e#���v��0��M��[������ƨyT@ �  �˺�۶ewwW�s;a^ z�r�WV1]����Jm�m�d��Y��� ��@ �P   j�pm�l;�� *�@m��;�`��ۢ��������kmk��<]NiQ�y���]��B�s6��vu2�^�D��져`Fn�#�DAH����x��rc9C���O&p�����^��E<xѽUOj�m��$�m�eʯ�FF񔥄������>��)�Ĉo0k�_�2]iWKp	�Y@�<�{?{��>�O�p��p�0�6Go�?iӦ�J��Do��lѲ��D�����(��MwJ������<�lܬ���V@�F=����%8��DB�����#4��~�0������$�B+��lfd�(�v-��q�f~
nù�f�L�@�H:��J�T����83�;S.�ۛ[�-��v��W�k���$w'�����4�.�}@�0�����;HVN	&�T)��I&dBI\h�n���'F��M��Py{[���x�_v�Sh�D���e�m	$��3Z�uq��[U��x�S�_�"��\�-��Ed.H�N@�rb���X�t�����oN�^��<L�Ye���!,��Jk�R�M�S�]x^PC�D�<����{�/�X�� �h1��cyS������m���
�
��@ 6�UW�N�`��N�$�x;�g��C��a��ed�.��~��z1q� �cn~'k�Q��xiܡ˩e�{���wbc�{��H�-3����3z�����_���ۚy��B���n���wNL�F"
�)`4�f�����Y3Z�wxv�^�쮝��`�ZN$�M(�mKw�O��`��2��`��2ƽ��}�u���ź3��Ǭ�$Vk�NY���c��J�T�HJ�Ҭ��j0�JBu]�g�}��ʟ���TF��H��fqbad2=y�q��l�.H�I
qP���穇�� �r�>?�������lTg���<k|�DZ-BRj�nU~���D�@F�iTp�F(��^J�4s!ނ��(���j���KY,���ַ�8���������ʈ�٢��I��ò�h��B?���)��@d�E@�id�r�?�p-�!鿟+ذ�]2af���[ZB#+_�y�|ra3��8�F�61*�0�IPcUϖev�U	U����=&W����H�Y�z{�H�4wW�|g�F~ҽkH/EzP�<p���%���d�I)"a�ha�Q�/x�r������B��!z@�=yQ�f�XX��Ϲt��T%�|�}3�!�G��0��wΦ���d��ϓH���,��^��Q��Ќ6�I6������++�^3H��=�H�4]�#x�pqT�G?j��q�^[$H�m"�e���W�����Ɓ�4�B�F�?��0�l�����{zX|qP}yyx߳~mV̖���U\`C(���gmծ�\ly���q�W.�j�Nm�������o=��@��e�����Е�v�[mQ��O��,Q;1�jIvB`v��*  �����*\kc���<�q3B�M]`�<1^��Ά�vw  P�  EP   =YGp���;�@R� *���eP ��{mSm�.ڛ%����ٹ�%s&�h���z�*�)�WUl���'<2[J�v_L�^e�b�L���#�6*�`�����
k�7IK*��"���L6S��D8L4Si#S�$��]U�_z~�D�� 23Oo�8B0��%A��ȣGz�$�J��lά��C�^��4��V^���CH���3����Bg��ׇ)~�6�hZq�E�Ln%!�Mi��$�d���#�+}B?�xK0��,�{�����q�\eŴ�A�?�3sS���B>"�{�u���#u�3�E���B0�7HA�ĳ�4��FSl�B,��9Z�9�Em�ꮷlw��Uw�[-t�Ul+uPM�Z
C���;�����,f���?��Q��o�z�����;Ƈya��ާm��'!-�Yu��Hg�U�|���Uk�(��w�#{�O�E�#r���d+�T�����22b-Ȕ��
q�ϊ$��A�f�巐"ן��ڭ,�t�ּe���{I�$l2\D�҆�(����H�>�?��ڬ��ޯJ��چ�l�ύ�םE��%tP��l��4!��Fk�a�̫ x��?Ya���!���T�)u�P�Y#"@�S:ݎ# �T�Xx��]�UBU������F�r+CB�Yi�֣3��ߴ��!�٩�f�����ڬ,��7��J�L�[�6�	�Y��gp�ٔX%{��?��ڕ� Xݬ7?kZ2��r�H�0s��2y��0��x�'P%�ׅ�kB��볡�7�����*�F�TDYapE�$`E��I)#
J"�8�.�\@]��r��������~+�ي|v*����N6�RV�lC6s�^ 3�w#g�)�4�3�����w��M����&�+fG+aZ���G �Iİ ڠ*��U4�f`��*{-�[k�$���hp�_71�g�ߴ��i��8����3\G?������S�R+naI%G(��FGr���>�����)d���;��`Y6�^n���B�rPf��]�Xi��Fo+0�~�,�����qa�J��"�JD�̅�cn k��	��>����>|q厛�]
����\���z���Ɛj(�E(A�'��g9wWx��O2��j�N�L�egdA���$�2aq(�IӺ��xy�6�ݛ,�TUpS�-�p���e��[���\�]��f�/׻gs7��뽇�Ɵen���nq�TInf=�������������L���G|��f��5R�"U�d������s}Y��U���E�z^쳰��_m��Lb����}����K�����vZܕG^�Tv�^�h���	��l�F�'qf[�ʱ+����F��~�_۞��s�s�����B�HHH@?��?� ��$�$�	!�H@P$�@4 BI?��H��$$$ ����BBB�o��$$ �xBBB�����������w�_�����|?���@�@'��� P! $�� H�d���BB���?�HHH@>�����ڄ$$ �?x�O�����o�����Ą����RBBB��k			�_��7�;���4j���?B�'����������~����?���h���HH@3i��?�����HH@?�����s�o��PVI��B�ӵ ��V` �����{�>�P(��AJR� )%@(�  
(��   �� �sgcE@�J          �       
   E  ( ((PP
  
T��� �   P H���� ��@�C� /s�����T�0 &�`� �Ю� @z  y$���EW�SŔ��s���)!�yr�F�ԗ��]�8���W�Õ"O<xOzQIWs:��QJ��t^Z����S�Ƕ��  )�   P@UBOzP���gW���T����o]��J<�s��J��� �ޤ�T�s�֩w��G�E.6)$姼�II �����	).Y<�JI�g%^ ��T��r�����g@*�=@SǊ�Q��W��U�꧴l�o0�r��X�E/8x��"��/z�^F�R���E����0���\�9*$�@    @�( ��"�R�׈j*���W��.{t�S�S�q�H��)稥��^l�$���͔�J�sc���Q���)O= ��f�g�J (  � 7X����s� ڽ(���;���),����t w0=wp 4 � U � �� 0 ��� stJ���qB��@��@q���z��B�)��T��9 h=��@e;��zՌ�t�����^�(S����A�3�-%Oy���%=�w��4� =)T�;�-Tky��x�n���Ʒ�T� (��@�  
 A()�

w3�-)��r�ղ��u)�Z{��m��G��*s҂��<���޳�y��;�Jr7�p���ꠗ�JS��g���7��<   ���gQ)�Z��ʋm�y@����]�#Ԓ��:J�j)޻��Lw��)@y���� PwMА�ɠ�� �=� 8��ޱ�A_ ��h�T�F�"��h���hL�
T�	�" ����TR�� '�T�C=Rh 4 jxD�z����M5�n��Æ�����Ƕ�g�<k�٬�w�~z�Hfv��) 5�.Ғ�R@wT� � � �����?��$���F㮫?�&U�`-�џn��=ҙƉ	�@��	ov�"ܶ�����0(=ڷ�fTB��t�,g*wL(��������fV��n�n��[)F�V%}��ڵ�Fb/��<���;�r�1�_}_Ud=��"���^��֩N�^3��v�VR�w�LnWPUyYW�M.ꪩU''����W��Ǚ�U�@���I.г�Qt*h�/*��h�+c�.�Y���jX�����Xu8(���'�P�84C�投� p@�/��C��c	����F��X�~9��(��ݍ�[m�VU�^�G�&/��*W��ٷ#A��3M��4�<���]��Yu�F���)��I�����������+�0^N*;���T�&,,侮�,�W�UT-��>̔�RW�s%vZ��r��[��B�Mڕ	̾U��ˤ�t@c3' U�2��*;WO*�E��2�b�f��w��d�j��7�cZR�#A�.v� �+�-�S�:��U�g;u{��:~��3꽚m2Rv+�7�X��4e�����*5p��h�w�5�t�Va�W��d�8(n��8�\�/f�R�a��`M������ʂ:�,����Y[]K,��wjCҰC�e�ە)�^��C��(�WYZɧ�t��bˬ��z�"�M�&^�KJ��������*ʗ��;�l^i���jw1i��.��n^�������BM�HiK�]mb����<_T��H�8�D�R%;o�)��R�[�b���&�y�V۬{T�����9��V�fAb�7oN"k"�.KmX�R�Q�D.�n�k���)ɓ�F��Z$R2�I�7DɻSAR0�ϋ�%�U��G[M���ַ�'v6�(k��R7��V���{7�Hf�̸�*U��&b��\�oPH
�+�v�8:'p�z�L;=��&�V�9�9r2뽾����c�^��UpS����y�YJ�-kD�ժ@k�֍��d"��vh�*���Ũ��rj�<R:�֢/������A�s f6s��ڼ�6U��Õ'�����~����6�z�K?UB+�
�[	�6�
ZJ��,N�{Q��GEF7���+H���wRg.�cw�1Ae�ݱ3[����[(���ˣ�e�V8�=�U{�2M��-�xĎ�+��I;z`�#�%��|��u(E���$^�
��8���a����I���Vl�F�'�0e�4E8��YG�&��A������%S&���$�b���oh����@�P(�$ݝ�ku;�9�65pe�6�\U`[�E�d�V��6�[j�X�0��k	��hI���e�3��QݫÛY���XSu"�t�&�Pw.�ֺ��R~�9��e�{Wԫ�}|�ǃ�o��9���R�!����/r��Ϝ�g٫H��7L9f5��=YV&�v��ܫ�s��� 9�O  s���s���9�/����q���e˄ܬu���,�b*̣�tù��$��	��S�n��.T7(VH��6�`S 4��4z�X(�`�W����wwB���֢���7v6tT95�VR�,��Gotԛ�G��
$HdX�U��E���K>�ժ�$X*����A�Yv�!�V��>�N�m�����L��]f��*.�U@�j�%�WY
�9�CY,�Md:��N۬Ӣηq���4�X/V��W@��I5��v���#���w5<:�$n�ٌ�jm����9Py+7lcx)n,pdSq�Ы2��3t��q"ͩ У�'Y�)�B�ZN4m$�k�t�4)�� 'ii����9%ͻ
�V`.�k7m����s1+�b��f��$h�(��Ό���v�[�Iv�^#J��ӛQ�
- ���1�2i�ܚ���Y�w[.��֜�Hb�H .���L,YgR��;�bZy{I1�ݤ�'.�ԅ+�;3k6��cwU�7&�oei��o�<#n��E�܄���E����i*)b�b�n���-a%�`�X+,j��z�t�m�F�2=��[�2�$�*��u Z��������=8����n̍��2Vd��du�#3Wo�+�OP�=	�14���N9�W�J�G&,�� 34��'�Շ�ZkY@�W�c6u�%�o
�af�� ]^J�W�R"�s�qJ5)�QU#�)�.v񝻦V͘���ٛF��{WR�q\�l�w�|�m�Ѹ:�pwYw� �YW�����Y�v�Ϧ�<˃bǭd�3r�t�݄#��0��M����xZq:��jTrӕ/1a`�,�[5��^�*�mЍH�J��7�l�#p��Q��I#`��0�äS�����=;�.h��cl��`�n]m[Ӷ�#�Q'Xl���To4�֒�ŗ�C)ݦ.����N�;�VZ�˥oEN�6��Ρ)��CX��R��ۼ c��s
��C�R�a���$�i&�-��Y�F����q��q�ۛW�6<"9�
���H�E2�惙P�Z�����H���z���"�R�T�ڛ�+Nh��ɷy�bcu�W%P)��N�5Y4Gh��D��ԙ��,sY�����jm�{��-Ͷ3A�cFJY�R��{�^����)Y��IN=�`��k%Snޕ�9C�	��W����J�zQ��a1_ZJw3�����X��I���A:����r:j����f-��p�B�7M^�-�[V�k�`5z�+Q�1��oе-m�`z�%1����m��9z�]>�$ά�3�.��#�(u��/M��g6#�ܬ� ���5�b�v,�V�=��f�N9���=uk ���?�Tƀr�A������J�?%��ٕ���93�rgX���U���f�W�$m{�4'w�;^8�{�h�%i�H���3[�:n�4��%̙��n�YJPR;~�xM�ۄj��:)��/�[P^ii�y�P����,���"R��BPS���`-�]�Eb���]�/3u��u�����e��c�X���s(�T©�c׊�c <U#��*��̥y�r����Mcܰ�8�!X[ܩ��f+W�]\�:�a��Y[�%Ⲧ�CHD��Y�ufRRZx����Z�++jb�n:������i��)��7Xtɵ��ie`�Yu1f�S6o��m��n�Ka��4&�P��Kv�{P��F�0�8�t06ȷ�����\Z�Èl�t���f�&��e*�ѭ��/o���y��J�w�0@)䑄�&�=���X5�j�[�y�,��tS�140輺�P��$�J2v����9��ˬ�1d�v��BjX-��l�����P��4��f�`9�"�N�b���Tp61MQ%f��Æ���k���䙬cZ K	����36���LE���^�OYt�Y0��6iVٽR��CGf�m��(Uؕ�D�B�f��NHE�c�d���X��c��o�|�f�/���UU�$cw�y�U���ʐ{��U%��T,L����`�/�M�Jl���sc�J21ne?��Ծ�n&4\�I��֛�RM�Y�HX��Ym޹j
fE�1m�!ub�Ơyyo-�.;l<�L�v��UɤS�7/Tǳ3l\�cKȔ��
*�"՛V�xn�B�j��*��]f�c��U#���D<�����)�St�1�bZØU�f�',��N�%�n.�FiB=9��{3f�� ���v',��~�a��5�U�f�x�묵�m�za�5�e�N�so�0;�V����p
��<�3.���f�D���\+2X����B��(#WCw�����9� 8��Uv���q^�#ov�� %Y�I �Ƴn�Gn�5)0���Z�
w��0�n���u�/.����/v]�N#����v��E�۠�y�-ɸ-囗�7P�S����4i*H��x��Ȋ6β����i��k(�IFnJ�`�@��Ytjг�3MwQgn�܇��4#�q�8��&���G�ܖ�d�q�V��w�Z�SR܊�Ѣ�[�n��x��2�
�F�&x�qIxfl^V��\���fᣗ5J��UM���Z�W�VY����L6�'�mH�2Sխ���r��Y�`#,
�ZM��,� 6ꍁxrJ��A��kbf[2��Ŏ�YO�+VѢ�,�5���������KX��U�nxp	;�9�,�9�9� ,��������P�w��:��"��&�9�!���#�����ߞ�y�kr��ˎ�y��e�EU�dF��qk�y[�2X���lhs(������v��{��%躳�5z%�KU����C#��ֳv����V為ٛ[\����n�X��D���Y��p��gÅx!}��;�x;�d�<�p��r�o�����9�89�+ӏVRǠ �F0ɼau(<f{�\PYg)����}$ (�8�5�C*�� ��Y1�1�(963�"�f�`%��x���I]�+�r���"�0��:�$���v>���U�9�>�*�q�(L�F[�"�m�cg9�|q����P����I�ݍn�ƾ1�[��
;�.�7��,mf7b�f�'Ymb,��Q�W�~���+��etu���	]���@��;G�U�,r-f:d�&\�h�hL�
n<�X"ܘ^]^���)���		굗g6��Ëa{m���	*�k�wX4w�PK����:�
��gZ�y�%�U�R�N��$��-���[Yo1��ꭸ�F�Ƽ��WKfn�����Z˫��^�HA�B�:y�(Q"m�j��)i+���-7K3kv�T_֤��Ú��r!5Kq�D��5��ec)+5�=d�,���e�o�Aܴ��(�Տ���C[��^����,�5Y�{�৒�e� 3Z��vnSW'G�VV�7�C���.�M�9N;{��1Aw�yi�4���M��a�e޹Fn�����b�3oQ��]Z��Ŋ^<�fZ����b�J`��12�,��V�T�K(';�eM�tQ����=���=��fYDN�xi�K��+V�P���VXo.�2U�� ��J�tjd֛&���R}�*�����p�r,{g���b w�+q���%^��f�Ǡ��Mbq��cV�0�JD�m��,��,�)�;���WVq�V�/#ѯ�c����*����oͼ�)3K&�'{����I��l�:q
��0e`�o�J���1V�Öέ��c{�ܷ�5N#��ܽز�h��5�)��C�J�#Y��UX���f�?Wʸ��}�dЅ�%�oZ��O��%�ܣCt�HZ��Q�����YQ�
���f�u�P����ۺ���p�s.�J5�{SギI�­��Ib+0Ý��E�'�!w�	��/+H�s]b�(����t��_In�uePR�a�� 9�A�s��尧�w#i�6;U�E��L�7v��7�{�-�n���f��	Pp�e>e��٣�D�� m����1��H5\�yVH�H9ڻ�m�d���cɴ�����t���ǘ��aW�� �$"A1w�ؐ�bx0<��ⱸ6/^ݑJ�:�a�h�Ȝ��ڻ@�75J���|�r� �<��|���]�6,��E�-7�d�G��hӕ`����V`�I�&\56"6�]ދ�]^Z��r��3n�`(�^\���oN;�p�#t���ǵ��V���7u)��q܏�eJ5��b��r��L���Ȧ�@�m�޾�߾�       8                ��                   �    l   Ԝ���   l      A�     �                 q��Kh        M��m  $8�6�     m�   $                     �m��                       � 6�                                           ��Ͷ            �o7m&6��kξ�l8�a                           ��G  ���� I�                    l              l             ���  l     i��m���$ m���� �  ��  	��9�-�ڶ�����r� �(  m�                   h             �`        ��                          �                        �   m �    H�֛i0/Z H۱��                    m     �            �@ K(m�`      pM�מ�z��,�ޚ9c��8��/q���۞k���<y�,���["��f7.��2zLu�Lk�����Tw.�Xe�n97nM�f⍱�WUm��lP�p�ٷv����Z)c��sf��i��^3����ݸ��G���\�#���kO-�j �s�%��˶A�:�q�9�����@q����=��r{x�x��n#��S�G\ut��.RNa`�W�W����MIX&��^ogI��v�=
ηu��ms�wDq�����8>!��)D�&9�x��=�c���o5��:��:�ع��XP�{aQ�A�tk��D�y{�X{�rn�7k������VBKup���oC��md�8�n����4LWok��c�[�t�{9����F��;lve�G/;�[�����p.m��bTv�/��X�ֺ� �	�)���n%:n|=��Wr��n"6G8�]6q�OiM���.w=��a�gv��.�|{�&��ύѠ��8�g�^����vpW�VIui��%�nȽr��qe��.* �뗓�UN�Ws�^������M�v�l0	��u�k��ml/�q\N��cm���#D�v��hq�rYy�.��im!��;�e�n_#���Z�sO���գ����ݥ92r�V�kS�״Y1ɕg�6�aގwmnVEݳ��Y���`�u���+kvt�f��gN6�%R�yo2+=l��X��l\���]q��{6�g���p�ԋ{�r��P�8)�M�z�N2��g8ܯ��{z�ϣa�%(��,la��>K8��8��`�Lr��.�g�]���mnK�ԝ��ai��Wo'��g����sA';x�r���cm�睷5�c�	\�Y�G�㬽��n4��7�<&{H�(����ganޝ���IF;R`�O����7�v�v�s���p,�x	�^0�ۆW��Z���7Cۋ8ެ&r	e0R�h��Q*t`��c�r<[�Zx��ծ{a��';���H�X�<9u�e��$�Ƶ�n�0m��Ԝ�y�]o3v�S8����e�g��ڱ6Ǣ��w=��E,�C��t�M��l�^6a-��Ap/�Cn����$�}Ys�5Cr��.W�0���m��u�u�m	�`�Շ3����f�sk,n�yB_}��2��i������7Ts�)vl�^��#ۂ��\ɉ�X�����}��� m��Z��e:��Ep)�	��]@{jx}��P/�a(]�Qv��q�;��Ӹ2m���"��:���.����{�.�g��ϧ��uh[.�uλ(�Q��r�8�˺��.Dic=<���;,�U��1���L p(��q��z�ra�ܹ��a7��<�i�<%NK�1n�;F��x�4��vs�h�쓽k���u=8�����z9��[fݶw[^ �͸���<��;r+j���L��9��jm��^:l1�W�/mnk�N)(-�E�l6�����m�r���ں*�4=�rq�`@ۮH\����[ˢӸ��Ś�N�h��SHd��{xg)��]�	�m���clF���|B�;Y�;`�{<��WdFx5:Ϗ����{g���[��ɓ�7Bn/ �9A�J맓l�7`ۡ�+���n�8��Nt�ط(�7>	/K���۲ܧn�W���z�q�'aOf{p��/>��8�v�/aR���]<ܳRA/%��M.vu]�&���'sX������箢�V��ǅ�Ky�m��n��n�hORc��gu����&���C��9�[�-� m�ݞ����rb�F�H�k(�Ƕ����8ڹ�v�c����ٮ�:׮�	�<v�4�O:���<Bg��w(�3oKaNH=��QwV���9]��j4c�QL�:kӔ�!k�c����ǡ��̠�;y��i0�OB�t�PJ`{v+�	KX1sV ����-�@�q�Wl`�,']�Ҵ��s�5ݫ���ٸ�ًr���J����l�c=pnp�ZLF.�=��k���ٛ͜;[�m��k˜u��1#b�ֱ|&Ifї;��N�7cu܇\�ݢC��Q���2vm�� �e�{&<г΀�����m�g��q�{]9�w-u��p�=���q[�s�uCq­�[��I֒ۆ�-�8��l���E�x��f���:7RN]�n=��T�[ݽ$����P��=G=�/�鍷]��wQ��,�i�(T�v�[�ۗ]C;c��+�헷�M�iv��g�������!5���6��:�	�&�y���F.#!��L�ǵv���7%�0���_gן����׎�9K���́�-gbK���c��b��:8O���]9�s�i�x�\�y#�T15[���:A�i�:%<k.ܯ;��=r����v��Ӕeۉm=sP��/��v�9�gW.Q��r�\t7��x�"Y�m��^ݧ��&�]{j�#�X�w.���T�鱫���tܜ�l�mK¤��I���'q��7���v�g6plvy�1qA�;ug��w2�\�]�e�On��j�I��X�砯F�CX:����Ƃ�p�@�p�`a�.T+tZ�*�һXj����;/ei�1;����7BgF,�Wti8�[\�뱽n�5ȹ�p�/iU����}s�m��{n��3���G��0��\m69�n�wfM�m�#[�.E���K�vd��EM��c�Z�ּ��ϴ��C�g���7m�����ڝv뮍��=�ۥ�Gҷ��p�9�mK��[�x\�5��������[Ҧ�N;rG/9�g([�O��\���ֲm�L��*p�N��=I��q�<��1\�ݵa��(�7UQ�P�A64t�J]�Ҟ�	��в�J<��,��m$��m;Eۀ4��z�W���v���|��7��pu�g1n�[&}oaW�<e�t��ðIGO\Ʒa����'�v<��>�s�n8܎�h�c�ATnt��c�Ǆz�c�<�ڮ&�v�x7P<=�Qͺ�l�F�|��ls콺X�]]eiz�q9Ӯs;xC�:�&����gc�X@9r��9��7N��w<��Ո�c�?�1����Fp���,k�]���f��v��?S���/�z�CLg�=��X�88a��D{t�{t7n���2�4X���=Yu�[؞��#��	�^��[�<]	o�����9��x5���N��2��r���ܳ{P;��}���2��v���p�Қ�EJ�79Nu���u�s��M��k�]�G=���rF.�c�xҞ p�6$֬tf���9��b���'Q�zn�{!�۷�1����,w9͓nx�q���t���!����h꛶Fq��v�c!E�@�u�Ou"8'P���x݋��8���:W;u�ê\+]ڏ��n�N�%�����E�d�c�·s�v���I�l䣊��oWB�w��$��}w�i�^6����=¼o�>,a;��� �G�	�u�����[�y��q�8-��pwE����ۨ�5%���soC���[�\��=����s�Wc��Yn�FѦ��':]h��}w���
i��q�m&d'8�,��zo.�t���7�n�+��z�p);�nW��ͫ-���g��;+���4��r�dy%���O 6�f��hr�li�H�^�8�e��F�v�m�y��y�wW�k�zŭ��1��[�sN��nѮu�+�-�ds�3�vKf/<���J���Y1<n�!N�h� u��^Om��9O*u��um�<{r���wO-���z]�t��f]��O9�87=��cq�ky߭���U���@�86]�Yx��#��y���uÓ���l{)�r�O	r��y���m�G��8L�E2u�;t�$�Z���������*ۊ�Z��R�۞��x��fn+�%�0f��ܽ��<�v�4�@�^v�Aۍ��3θ���Z:n�nη#<�2,������uAͧ���I8��Pׄ��m�m��їu��XY�8�J뭉zMq�3��@��U{JH;��w��wwy��������   ��   ��6� �@   � �Ki�hm�   �    6�        �`       �WX�i��        � �tj��̵��         �          �K3.�   6�6� mf`;p6nˎ����q�7��n��#���u�]��8mo*m6�7[R\�0q��gJ�ՠ7X�I�Tn6��p�9�^7a[��Y�s��-�k�}�yv��ǋ2�Ȏ�<�����ذJ��3ϵ�N��9���3������]OT$�;��*�������8Ű��b6�N�1��^]�����뱅�ݒ;)l�v+e��N�=���%;E����Ǜm�u������]\���ݭ�F\�w;8��:�-yz�5`[qF�c���g�g1��v-Wlq���صm@�$�eѳu�jrq�APײEr1�����&�/���v��lH�ݗϚi=^P�m�m�˞���]����Cm>
S�Ӑ;���Ƶi輶��[�rkpg�i�˫�v�%��] �n��w<��v��s[������Ix:�mm��8���Z�J.:ܯ]i����rxX�n;x�]����]�ӟ&�[p��nԗ����m��[�z�r�<\.�2ȶ�$K��;`��s�k9l�n;$DY��y)���=�3s�ݼ�8sv�Af��W�\�����L�ԍ�{<V����[��=��;�H.��mJW]�[e٬q&mn=����x�f������n�nM�Z�pf݈;T뇫�NV7�{m������p��zO"��v2�lu�H6r�R�s���d��z����^�y�g=n�vw&N F�<���y�7f8����ŹV��FY�p��:2wdB�n}����.�:w6�k�ý�{������{��;��ڶ$P��m� �-�7[� �$ �� /Zl���z�)��xT��z"H��"nf+B�;Z����t�-ݯ%�/Wr��up�;���t5�`�7v.�O ;���Sq�^��	ҝM�p�':���t7�8X�٣����W����{�nzݽ��q:�)F�Qxv�s���n"�+�;[��������4TLSWL�p��x��Tf�*t�n*y|q҈s̝�9��/�c�>����@�{�E��+�
X�y��N�a�����&���*��J�/$��<p�-���^�N�GqF%��X{�N�?����wݱm���@�$i��ic�xm�f{-,�+^���_�v�,�	�W���[o�[�p�Z���EIKg�ȼ/����6���ㆭ{	��wJ���%�r�{S|���RTŽ,z�~D�6$�l�[���^^�^�@v:����y���&F��bW�m�S��n���}[�A���Ʈ������%�ӝ��ɺ�r��.tҷY�a��on�:�x���Q�� vދ>�8���|q^Q���ܛg�s��'+�
�\��{�%˾�� m|Y R�:$Y���b��1ɀ��s-�>{x�v���ȇ�r�6歛�ɺlܮ�/4)ϱm�0uj��k
d�C+ڪ��aֽ͹}Z���9#$�)��������4��is��g=�[������̂���<=�Y�`;��|ڽܔ�u,@�R�d"BF͒a�)�[�ζ�:�Nw^��/���Z�,��H���X��o��nyV����JUvB���D[��C6�j��}o2i܈cˏ��%a��5�5p��x���W��]��f���q6�Ʌ3v�-��u�q�\9(M��Qr�m��f�E�^w.�i�)�z��1��i���!��;�z]��5�Ժ�M��.���HI&���"),y�L��mn�7����ɞ�V�x��3���`���a�^����=��Q����DP%.�z���^��;���3N��f�]!쨏�/|s;q���l�vrc/6����n��q�T9�f붤��yu��c��:s+���p��{����zU�Uݔ *B�G&Tѻ���۩p)�9I��+���{��Y^ﮦŘŝ��x7��z�P�h]�$��*�􈨱��<��V�fN�C���t�<q�=�zd��]{����l�v&�ee�ͻ-��7":vܫ����о�������Z:�v��n��H"�
+�y����Ȱod��~���xY<���JA9f�{�%��m�J��x�{��D�gJw/�%�~�q�ys�bW6��:�M��~k�4�jQ8�v�ȏ���o�}Q��%pP�x���3�ub���siD_���D�B��B�H���A'�����@��!<ά~�:�i��A}� �W�7e���ŭlf{�ڏr�o4nb���W�'�v��7�|�WG�OO�ttep�\��w`px�%��s����w@�����i�U~�/�Ժ!ؙ�B�jJ��[��ܣ���g�5���յu�<�JJ�]�JW{nƎKs��,c<����hܜZm�����}<l�ݼW%X7k�I*�%#D�gf������0��{ D����}����"��k+ۨ���Зy�ʴj� Qsx���)=�u��}O{k;�kc]�!�[�[v�՘��5�n�כ)�0x�p��j�H�1���"^���X�׿C�-��<y�懼��.�����F��
H�B3��i�J>>\���yAq�����H�h�S�$�D�k:�k�{i��Ҥ�	6HUj^^1ș���p�H������ڞ�oK���x�L�P䥃l�ܿ+��CQ���f�MY��@4��ڈa�/+q�9h�_������7��'�O�5�m�u\   �N�� �a���OV��   ��`��.�V��<��L�����ɬ�lq���k��<��`;��]��8�����&�Od}�'N�;�N�}����x���<9G�"^pGm<��Ϟ�k��9�����b���:d	��;u���c���l�S'>�=��� �<��M�W��u��Xo���#�������'��g�;D���s����vIoHs�.�ݜ�	6D	�KR#�z'�v����+�&����V�:F��|���L�rͮ��d��U#H�
�E#3%~��#7=t��4��h��I�q>#E@8��ؚ}ͧ�.>[s{����S˞�v\DP&�QJ�%%���_�7�wn(�B��j����[���e�[�挕�����{�QF��R��s������|�3_�w���)6Ͻ�Z���k���4�3|tz����e�E]
��YH�u#��{"�=�L+��jO�ևw�yw�,6�M�M��>^��NE+$���h����[Qؑ�k[�)���^��G#O�2޳u�9bl��+��7���o�k=��~>P�4�����@�ܻ�^i�sٸ�6�l�N��*��H�d 
Gb��_���ۨ��{Ff;�J�4L�z6��:���iOm�ϻr��X?7\�����7��{Uxct�e5{9P��N�x\^�k2��ap�;$K��:ւ��u��ӱ]���4	�AAB�]�Hܑد?Y¼b��=�Q�sK'�3Q�#�<�*v}Y��V ?]ZWj�@�{����^�7�|����y��8n�*3'�yySs�C�����=-@�(�H��̋ݞh��E��w.��1�szV��^<>]�b3<�gף�HT�X>IZH�vI�b�v%���=��z�t�!�7��pa����<<LΩ5���]����˓ׯ������j��f�B����=^��_���!;��Cg��]���TU"
B�)M���ė���|=��>����E�kmI������/l#_b�{}�s���"hդ����y#g}�6K)��#1���2WW�:�ǎ�F�?d�˼�1�lr�������r�v�H�6B�Eh���l}+p�H���9�{�y�~���L�/�|�A�L���9!Ǟ�Nؽ��WJ���"���A30,X�}Oe�g��M��p(&S��|���8X�	��sI�������^L�?.�U�����^G�/�Ǭ��w���z�\6�U����׉$mq�9�1`y[�qm��jMzN�zmV�}��b�]vՄ��)��SG{�TȔ�{���{���{����=~��z������L�$��V	�WiU���q��ykŸ�[�5�*��"ʙozaáw�e�N��rr�"n�uR&�!QA$����~>h�[z�~���nǨ}������i�O��=1h���Đ�	Y$�<���i���i���[�~�{y��,K_��?ES�;$S���;�67p+&�����
Ng���K�(�r�w�Sl�L21eKp���#�)B�����JJ� @�h��욷��h��*бLl��$f���p~H{�N`��لt筄b����AR�hU[`ۗ��Y��W�����K�%��7y��.���fSvy���������>z���T2���c�s�����]]�D���o���u�sq���Aj�WiXQ�JZ7�Ft��[�!���f�{p�wV���d*�{�"OՃI�2��"�݄�@ �sOk~9�<�m���.VVT�u]����{�E�ڹ�~S2fe>�+�!�A�B�]�(��y/W�[z�M���f���	�8�d8`2j�n:�|W���-��b��$��H�B�<����AG�Wn��\�'���=����-�����[K��~�Ë³q�M��)���Y��a�-Q�j!:xD�@�_��_�/�[�_}z=�8�6ؑ�h �`ڐ�( u��  ��`h�K�k�o������M]ˤ�j��%�u��;���Dt8M���dv�ޖ&�t�1��^q,Sv�^Wuϭ�b�m�<Xw�v�lv�f7���ͧ��M֞��F2{uOa�`R�q����F�v��>�e絶n,*��խPV:�#c���G�
�>T݃�ܐ�n��MSm�6q�
���-۬��J�%�Ry��{bڤٷE�	Sn��ukJc9��M@�@��)yE������F=�/%�����Wnj�y�hjRomxj7e��h J�DAJq������qR�W�������#�r׃��=�{<Y�e�Q-��������N(
G$�Vvn�G�V�̘��5Y�.��)C�(���y����]@"hՒ�V@	2p�BS� �o�=���-�NY���TMGGڌ��=y\f��/u���,
�u��׾��#9b�ڕ�;��F�0g{q��{���|����䟧�=\��%�E����N^Y�VL<Z�6� �{[8"Ñ ���v@�
h�P�JK��$7��vk�^��ɓm��j{��Ҽ!��p�u`��z�/;���j�Т��%�Q�ŋ�9��<�ِY���5���׽��8�s�6J_]�4U��.����5�,����X����֠W���OS�/z�>9Q�^d{�T�;�N���j�=J�6��J��(^�O{:	�o;/����}/}b�^���%�^��S����$�k�H�h�E��M���� ��l*iՑ������_{�,�zh����^��N�R�+�I~� �]��+A��G��#p��'o}���u���(��ջ��Qk�9L��y;E����[`���M�b�g'X�\�Rm<���v�B�F�v���۪vT�����8#���\y���դ��}�m!{��*��鰷�n;g�ym#H����Q��aZ���f�m
;u�b<|��妷���F����p}[�aMps�u�%]�B£`�����w�c.{�p�)U]��3��g=}G��+O50NC�i�+%;ę��j��`�9!a`�:F�K�^5�,�&�N5��̰,��#K0��`J��6^����i�˜���ݾ[��m�X��K�^�0��ԥ�vm��t	}ρ�n�j��T�gn�.�|�T�m�����}��!C	`�v0Վ��n��_ۂi�%�b��t&C��F����ܺ�ث��ko�*t�7��]��H����`�����
�Жv�X�3N�Aq��n[�����݉% z���WW�J�r�Ep����4&h�Ɇ��X{���f�9�u,�F�7���vKJ��pyZ�ada�)�`c˧FĽ��D���*m�#Q��[u^�ͩ��e����Z]=�:T��Z�;����<˼ά�F�M�k&�9�얯�H'aL�=�w�|r�'�h�5�.�AY�F�g`<�`B䎴��Ւ��GN�d�*];7$<�Y��|���aU��sv�Z�Ju�������EC^X��V�o.�S�ӕy�7z�����姳\:�z����Rqs�,g���z�伧��l��M2�����'q�����mݞ�Ư�[`��j�Stj6fPoM35g'62�����zu�z�t��ݕ�}�<�x�v�Z���e�Q�C�y���y�H�eE�D�N�{�}�M��GbLd#�#�[	��;Ci\�2z{m�cz+;����ǘG�:F?��>&�e8��"7�"d��1z��c�XDx��2�q��n9M�����,x��$mm?D���#fODUuu�"�����O����o�^������u�$!9�a6{<v����x{n4��m���jb��MQ�C��~��启��(aı����Kc�hB�v��x���ZCw��n"�����v�;S6C��<�Y����w{a2�JCrG%s��d��s�]m�"�jY�ב�QQӽKb|Ʉ��G����E�R��S$��v�Y��(xf%�lw�8��u�k-dRji�%���!��Y�v��a�D<U����6(�OY�y�gG(�#��n-뭦�l�ь$���o�� �Q��R8)�|įD��}wTtHӤY��E�V~������?��V��3�0�`
��+��+��++��c"r�:w	��?A2%s1:UafA�}Yڹ�n�n]d4I���n2KH����z���kH�.cB�>�Q��-��%Ǒcda��y;�˦��>�a&@�x�&��횚{���4��BU_҇�bH��J\_|z'OOH�<�'��ퟴ�sn���Hkѫ���T�Qts�:ݙ:�ӥ�9�4um��o!g<gH�Ӥ�I3�V/�.x�D3k��C"��<��;z���2X�"L;����%�^d;�'/V0��"j&�\ɲ��18}#H�� ۄ��p��jJD4GNdov�"d���Ѻ��e���peq�!�a��D9�'��$rbDaQ&c�"F<����1s�{��4��\ěN#\ÿ+#��"���t0�0��|�K{����,���k��x�R�A�ϕ�6E��ēe��DQ��M��14�e)�8��"͑�kha��V��W�VE��N�E�����Dcz�R���7�d1� �0�zk�uQ����:yZ��dT���m6t	$8RI|`�!�߷�eX��Zp��Γ>�6�f���y'�D#���}D#����!Ϭ�>1���g�(u�Ix��n�E>�MtZ��U�l�cV˭�G7���)����6�]�3Ǌag��{���������"@��֤�`  �˶`k���l �� ^� ];j�m�u��5�f]�n�CŴ����U;0𮹮ȍ<^�{\`ƭO ��wk�n%���v[�湰�h�Xl�c�î0#��xo�P0q�ڄ�:��,9�<kM���uFm�(�ǵ��;l�S���u������n�W
��K�!Gq��d�Vb��Dꭰ]c[���]��fE-ǒv�^�G=��l�ǯ����=lth�ʐ��FYm(����f�e>�$��V��>�,�!��[&���v��"��"����2p�ֲ�����6��Sp(�r_>"�<Ї�l�[o6e�����C������$�a1��4oS�Ia'�G_N3\���p����
><ۤ���1*2�E��aHÄY~��|����,�"��U��Cwfސ�o�Օ��"Nu�#����H�,��u��Q)"j3i7smQ�u�}�I<F,Ήt�!I:��Ϟ�1�0�6C��y0F�E�A˖#/��s�Y�H��t�#f��d�[p2�I8�a�0�z�e��ɈoV�F|~?X^��4-�4�D�\����]r�f�(��l�p����G��k��M��m���Plb8���}g=A�َ�'cN&K�^략��$k/[��
�lVw ������6l����],�#عf�V��W>�<�y_Z��
����i��Α��D�gҹ�(�8k�n�E�i�JP8#m8�8A��HY7v�s�!>˽�/&��E�����K*��懻���W�����\�6T�]�IAf���,������)��e�
��<Da���q��#��.��2	� �Q��z�硄Y�L-��bTO��5��$�Ěe8T��J�qQ�ay��<�8�Q������v�Dݞ�ƭ�y�w�=���=�c�
7�oes�3�>4x�����E)	4ے�#���L�obH�C;5���2|�f�ѩ��"��f�6���萙��<�*L�&.m����J$#�"Ϡ���j	A9 �)d$�wP6���Oq�l�#�\�u�{IN�WP�C�?*?��bbd���<�7�F�"�;��������G�;��QJ� �I+��t�K��2˻�޺�%�grp�N{n�˸�nM;�k,�6%���ߧY�w��{�\�H���ު�B�Q<������C���sV�1�aE>��Nf�!#�D����j`)��Ԓ��(oe��%ӽ�uD�YB:�}�C9�(O�N2�C�"���y�"��h���ΐk��g��_/|GN��a�E�FK�$�q��.QH��l�ac'��oGS�}:ۀ����64Y!��s!h�H���w�Թ+iiZ�T�!�+8ñM����Ks�Ez)#u[����)V\O�l�"O���U<��V wv�I$�K�6��^�i��*��w�����*�F"���l����&Q�7��R<�D��Y,k1����p���M-��}k��U��D��c� ANDRpS�hZaz�F��E��[װ�>��G}e4q�J&�Dkz�G�A8~裂��A�qK���u"�\�y���ɽ�M�!Bm����C6�D��X�
���-�Z�v7]���Nފ�n�V�TM�Ѷ
���F�z�E�z�B')Đ��`ʝ��"]�ɂ�c���s"�z�WƋ�4j"��y�e�dt�ÅB+���/A��nH��Ic3�,\�7�*�
8mWO6o�%���{O+��v�2�ym�!I1�Ĝ"��������}�kTaR�i<�9nq�%s�<����_S4:y_!��t{{�|8� �Fh��O�{ۙ���lz���v!wYBh�FSzT����f�"�8�e@Kq���#�ҐXi$��u`�nn�+�fY���>����50FHGլ+�2$a��Ht��ڂ�tv�U�]������4�n̫L���m�ۂ��+�Hf�!��ee�W-��a���(�詙��g2i��"ә4���8�)��i0�՚QP�!r�E�%>+�Z缠=(�[��`�w>a�Z坛�L����"����\o<�D1�`O���ݕM�:E�#�L#�'�B�4�m�mނmq�6tu�����T�Z.�ln�mNH��[���xڝqJ�lt�Z�=��%�DQ��v_0���#C���[[��8�E<�=��C�l�u�B>4D!G}����#؄4G�Bk+ImG"�(J,t�Y���^�]�4-:d�7���މ�"H&�	>���$a�g�FON�Ut�F��V�h�ߨ���1�Y}M2NB�h��g�GO!������}I�ْ���(��ޣ�E�h�<FU�C�~AZ��@�������C��#״s!�&����2D䱧�YR�ɷ84�/rWD��"���8�j��h��,�GH{k ��9��z�ݎ	��b�Z�uyQ:h�m�$��.�e�@�����m�C��GMZ������5��6yX�+��
��b�޺�8�e�>�a[;�"}:`�]��M��s��E�I¦���˭�	Ǽ�f�����0��ȝ��h���^gM���xٳ����D샫oy�o�$��[E�wA� m��֛M� Fٷ6�   浀���[���3sO��,	S2X�Z{uX[��ę��m��llNs۞-����p7F�]���g����6��Np0�-۱0c۞�L
i�N�s��[9r�"��从.�ջ�w3]v��M�gN�n�+�󵭭ۉݧn��TV5��l� NkK�uv������)�kb�j�\$'X�.��+b���!������s狇{Mr������}��k��4p�~{�;�k�~��?_��y�#�0�h�ooU��F"(�_�#(T���м��l�i�F���=k�+凚�G{	D�đ�N:"��FY�{+�.^|~�}�O�,�D�>r,����#�D88�'�|[[����r����ݾ�>$x��:HP�@T$HT��O�J���_Wkw�Ǎ�H��G�mu�H�8�Y	iz�$��N��>�;�D�oD��r��Q����E4�6�\RP�'��G*^�$=���a�+<Ⱦ=0���F�ޢ0�HS���"ὄE/u�z����
!��8DI�8)\��CA,p�m8��>6y<���w��P"�{a�Jn���m\�D���SN��$=��rX^C���(�~�es�Μ4x���z�����[Q!J�\9f܋-��kY�5��J\��웧�c�5ݷ]���I��faI'�8�GH�$B'۷+�?xp!G�����O,ø�nlk����8�B6�I������>�'c�[%�$"�8RIzG�z�f?��JOdHI�$)��>��@�������]u4^U8漟,�gR�"��טb~��T�@��Y��df��{�QT�*��D�H�Fcq&�KW^lO��D�$h��m�4.":y�Z��s�U��<]��gu�<O5��,�Q�RJydt�֋#�w�F�<�W��ǐ�⹺�\��,��g)�狹�>��f�&Nkqys�0�+�;�Cy��kM��a)���9+�"�7/�vQO
<̽�f�a�	��4N�ܮa�؅EMމ}I��i���ȔGEf��#�o1F��^�ңHS�$�%��,��|�G�i�az����:Z���k0!M�26�ֿ��,��'��$9�4�q⊋�f�40����5�+����&��]��$!8u�v�^B7e���Ѯ�
	�;<��!mM�5et�cv�����iF-�b�.�{(adYÇ�l���5�y
<� mkD��k�}DKdz���8Q5���B<�2�ωOK��mHY@��x���Fȫ����0�.��x�y}D����lJ�2*�dA'T�7I���{*���(Ѡh��>v�nP�.v}�Auc�ΐ�Z�t��H䐆�f��8W��z����u�<��Qѽ�FS1ޑ�������.m]�6��ձwt�NbΖY� �Z'&���v��w��"�.��-�m|/�
j+(e
�{�<L�!oa܊��I�V�x��	���M�t&�Nh�b�f�Qs���h�$k	����i��?D,����y�Ab�4��9�ɭ0�HD4���Lf�=k1<�>�,��_ ��9�&
M��p�"r_<E���Z�Q#��>�Z���Fv;.Q:C�f�D���������t�"���{(��3Μ4B/��6&�bS�C��		ۗ�.�n�&��m��js�Wl��#;&<�ܽ���4mnݺ�]3TE����N����z�����"��ǚ�a=*/C�����P�^�/�Ln�b�E������b���Yh�/�V�%"p�#�9¤��>���O�3��̍8��,f����h����o��O�E�(0C�WTP�,�}FA��H�=�'7��QY|��"��6
P�0≆S�őd��Ȣ:/ov_<g�����.��;,<\��W~�F�O�ݕ��O�0�y�,�{��Qy��V�"ddA(H������0/�4�iwݔ,�1d��:�E�(���WV1�a,(�Qo��0E��'U)���`�g�!Y�$��_\%�fKb��)V'npU;�evs��ѕ�Fa�N6l�9J)��c[��4F�ɋ�s	-��1�d�cǐ��������/	��+Q���3X*6�̍�Y�=0�"���Aux�$�"�#��C��GO!ù����%�T�.9�Ej�&�{v90o<Mv�	�u�p�ێ��<�5��fzf�-8�@�QA�����G<F�6y�Y�Aw{���D���,�5���爣�NG���A�iѮY8A�l����Da�g�kWO>{~b0aN@ѐY�̌"I"Ξ4E1޻�N5���vc���[�qy��׻Q���Ν>�a�Վg�D�BȘ��w<�}�2k�<n�	���w��s���5�}�}�k���>����t0�	��E=����1�-�����ib�RsC�����Wm�R=8EaƺE�[��vcQ��q�d��\V�,h��N�z��o�0��x�����|yg汮V����a�"�;�`̼�U)|_|��CJ�C\�3~�i���%I
�qI%��OWL|Q"Xq���20��f��As�򊣻=�"��&O��4b呆i wv����Gm���m��.7���?6]��:�
��P�ܹ]1�A���?K�єތv�쩛�Y3�}p���+	wf��]ь\0m;�������Y[���eBeV
��s{��<�)u�ϴ1�S�Q��jl���=T�*��)�6H�-̸�ݙ\��&�'s�i���Eʢ��qQ���J���~��=z/c�jf�p���J�]�E��2�j�xҰIbu���̆�b�'):��tM���۴�Z�{ڏ>m.�F�}��뻶j�C:�]dwZ.g^]�65�dv�f�hv�76�00�F�i����}�2>׼�uNv����H�]bR�4!b�]"�!CZ7�6Y���%�[-T�d��@���{Ie��yU��Z�<������;۵ڜ�خ�)�+�m�Q^\Ȯ�V>��d�4lx�t6Z|��gq�7�2��GU⠆tv��ژ� �]9q��˫��H�v�d�*ᓒ���Nَq�X���@�S�T�T�yŌ��f�e��}����a4pś�[ݚ�^_v!ݝ���]�ޓ���]�;ci�`V4�!���޻���u�`�]Z�S�4b�^ a�f��c%���K.�q��YTmdgT���c!#2�d���T�n�5�c7�m�5��I$�8      m�� m� �   i�����Z�7 ,0         m�        	6� �ѵl    '�\          m����6 5�l��ɛm�   l         l    ��`����0        ڶ ��m��^�y_3v�솳�y1�;q`�GT-�a�]l�s��N	N-:�tr8x�']�y���w�q�(to]3z�&=���mF`��xm�g������[���]۞��į���Gn6��\��z��ƺ�z���y�1����n���\m2�ۡ����q�u�W��q۷CN��1:zM���y�ҧ\Ld8�-�%v�N�on	���z�Sh���u�����Z��uS'x��6::�im�C��ٜ�f������n��h���x6�]��ss�'���>�5���N��G5�F@�ݍ*n}F�v��os�i��b;Pm��|]���*�xw��<��Yc���5���J[������^�'\r��ktWg.�v�[���]�-�<\�2!��M���Nîz��vޫ1��h�^ۢ[õ,�dX8�8I|���Н�	��l/o%':�-g�ڸ���;sm�)\�H�kt;x���nzFx��w��w]M��)6��ptvx8׎l=x�a��k:&�X5�����Z\q��X�A�[<�M��cc��������^�j�<v㛀�-����ug����&�����;�u�z�x��v��isS`M�s����ד�T�]j�U�΃rYt�����!b����kte�f�n�W��e�˽H�2��"�����ۛ��(Q������y���ղ]Wm��cw-�\���@�Z�i����\�gr��9�9��Oxx7����z��F�</3�֩��/]��n�;1�:�ٹ���1?\��K���{D�mĮ�ܚ� $H�$SZ� l [R Y-  n���    h6��Fӷeyݱ�m�;��أ���v�fk�yz,�׎��N_5E�릤�,\s[�絏 :��o���^z�N.��K˶�\�y8��wn|y��lf�d���v��c�zݱ�xA�Վ�˶���^�]z��U����S�1�l;�M�8�;J��k:��U�;hY��qE�y-����i0��Wn;:�����#�4�.�N�ӹ�̰�d1�ڶ^r�m5 %��|E#(�Z�es�����0����{���Fb�W^�H��z����t��ʄ�G&�Ooo��[h|���(��Y�1�`��nI\� �Ȃ����E,�.�I3��D7�,����W!:EC���\�:y�O}+RC�¹�P�|��\=�3^�4D�$�I�}>"C��"��n��G��C�;R١�4���D+ޫ��2O3�EWG\H��V�"$ك��|�d4�Q�"p�����ʕ��F�ǁv��	<�:E����E����\�:A��t�g�����|y�5�֞%���"�VD�jo6)��$R=К�Bԑ9n3Zz<�և�,�=u�^�a'׌(��� gd�HDi�4�L��,�
��<Q��o]�^/���߯��β}���>�i�t؝6,���z�f�y��6��p�tn��{��4����b&�)���\1��|p􏏸B�>��鬔,�&/�e2���aG����ޚ�2J��aƳ׌4�.C	���$aR�<t��mw;
m��%�	i��E6\Ӱ�i�����O��#���=�6�,�ީ{	����҇>�Tz�1�ˈ����ͱ��l77�:i�b�.Ҥ��5d�>{�Ǒ��'i��cQ�q4x�0��.I���0�U|�e<v����=�vᙡ� ��x���h��$����kA�0�]�21$E�|yE��w�*��dM��zӨ�`����ԁ������Px�=#wmxS#؃<X��x�zB�Тl�3
F���a�xгi�
%�'sy��E��x��H_�w%
��I�N>����9�Q�	�N49+��y�4����.Ygܟu�N$ J"$I�B�2`���OOtHÄQq�}����79�5	t�.h��]�\o<���>�%��'�gq��L����Jif��_d1Rm�����N�'��u�wWI�Z�X6�t�1���s؁���;���$Vx(.��",i`���"kg�+ș�c�M�ϯj���5Շ�^�[(��{K�ӧH��z�{ba��z���Gt�DKW@�n#\�!�~C֑��yii����q�>��zqD���a};Ǫ$3�d�N"u�����4��w,��>��:���ֵ�JZJ@aN3C�.Y(�ݭ��3R<+�E�����s�OET��H�i��/5���r�.]�;��h[ْ�SF��d��&�N޳�4���1[�Zu�Q�՛~���1����K6Q$���*���Q#(���i<# �8	���b��sDȽ�<eƆ ��6�hi�;�)���VEb�"_��q����	�Wn�'�rLE�\d7��[y Vd����fX���}��=޿�}�t�,U��2(���D������l>��Ȝo1�Q��8��B�"Δu�M��������c1�������fjh���-��Aa$��V�u�]B���`��a��1��]�Y��5��.vh���ag�,	
ٺ{�I��"�����<%�G�6y_V䠗�W�Ȋ� ���Jm������n���=qeL�:͛�}�l�����98�~ܼ$�/s���⥙g�7�	�c&�ԡ8ނ,�52��މ�m��i�����*�ja;��jӆ���C?f���rAd�CnK�DO<E��{�A(�>�5t���D5
.�=i�&H�}/#Ndad����[��"ȲŎ��a�Bb�I��0��Q��[h9�60u�6+�m6J`�����C�zJ8Q����D�,aG��i�bbKc��L�H-u�\�����L))ݍQ����i�1k/GK繽g�p��꠯����u��j6�����}��r����V�/<>ַ�4dr@�@�`�x��<D3�Z�7]X�δ0�uj�,7&��O�M��bJ��,�����"�����"R<�}]<����ߌ��߾]��Vbm��e���[x'M��|\�wl�mbz.V�`�Nx��ל��P�H�H[����/�x�,ѹ��\Ρ7�KP��ڕ�X�����B���4$<��Q�"M�� ����s�>�6�b􏾇S^�ۑ(Z��+�t��_8�odqY��,kC4]uJ���A�h�[\�Дޤ��'��뉓gU���43��ar.;r�6
n�E�(a}yXG�|Y�=g�\�4$G��V��;ݷV^.t��(��"z+�t�E͕l�&ވ1zz�Ǐ=8B4F{p�D�RB�A!H��&�h�b������(����h#�#�����w|ä���پ�0��:�09{������|���"�q��b�N ���i�).�p�ZS��C
,l��̔,L6A�]�m�\H�a�M��nY���(Rl.l����ΩNg��"�D94������׸�{�7+�����(��;$��{�4�]b[�N�V���l�gS������F��f��vT&'��I$�WiH��h�f�  ںl �e  A��`   ր��m��N�ݲ�GV-&�k\��&�v�<�X7T=�ؖ�3��>�{=j��0���2s�<�/ē��L���nl�ĸXӞy�k/+�_d��NwZ��Kݗ-�����8@o`��7D�����y{F�:E���Qh
�#����u<��
�6���L-�d�e��b�U�W	��wDnx��p��8vu<�:�84d^A���r�h��뵼J?�g�O�;N��ٿ��qQf�C,���<�s��8h�s��C�V#{��$�����YG"�+~"�"f"i cH�(aR��3�TO�����oir���̎��,Q��3ܮ&�ki}��ͼW�쥫ǒ˯c�ՆE�}:EmndD�bE`R"�q|E{ʉ�]��A"�0�N �c=;�>DI�׵�	�?{�C�����GL�CD/��F&� �F�D��u�J
����0��x�OH�s���g~ܖ,���<~B�$�oe�<���B7��ZAČ>!�gد^��Β|��Ϻ����Y��p@��$�gQ6y�Q�_hܔ(��0��1;��]�EdO�� �!K""��ha�:G�7j�s�xO���d�L>���U��)�#i�-�H�&��Yܝ���^;rqۋv�Y�ۇ�Y����F��2[�E�c w����Y���'���~����A�&`����B�1�0�H������CgY��}Y��&AG
Y�j-��D��%"I+�Ev�s���F1��L<�_5�]خ��W�3�<�8��Z
�.�{<P�Y���(���⚉�0����:E{�\��$	���ݔ�ʤ:y$.�8&�� mi�>�`���a����E#�@�q�� ��x��go{+�|h���������a��l%I}=qA���!�+k'�޳tp���$E�S����
8ԑ)�;d�!�9��a��e^D��z�|o4���e	wYɦ��DAy�瑆���R��Ѭy��Z�����#��oL	���ܖv2$��E�C�X�DP����G�"J��،��Hnr�s4+Yȣ�|�Wnܮ{�C�"�+kvP�\�0�I"��������������՘���pg�7fug&��<��h7k��
���l]�0�B�:�N4䉅��9�������EPS��t0���}\�6��B��$m$���$5���Q���A�Dsŧ�#ma���kX�lD�q� JFn��+!�z{�o�s����4��(���0�4�0�3l����(aDIN�
4|��#���󎭵!����&�
M�!F2��3ާ1blC���rP�-G�(��S]qN�,�Y:�|�执����ʮ���ߨJ���<nu��y�5�%����i����s��T+B�8�;^����K�����7�$�������A3'�{���R9"M�ܝ#;O�x�8Q6��#qoDi�tG'�0�$���y��4��}`���yQ�G�\����H����
h�Ą|���
4F���M�1Cr4�a�%s�Q�O�O۷���$E��-p���;Xzs"}Z��D0�睝衇�V�	����P�iL4���O��iZ5�A$�_I��Kn�+�m]��y��mij��\��m���0��;��R�`݊�..u[_˿����Oq�*u��ϕ�6p�兟]i�B�s��!�+�ܔ&��;�"���\u��3b�r�'Ƭ�=���0&KL!"RK|p��*�F���C�n��P[�`b:?��[gEQY���,(��u����1�Qn�]�H�\-h�������I�E���#$����#O����ȯa&�"7\9�#��̋�El:U��lp�\P�t�<d}Hx���T�������wo"%�(3��0_0�O;�,��	o�:A�֪m�a���M3\lG)�y�&|����,�ȳź�vJc�=3-��-eL��Ƴ����u*�!h㺖�R�B�",�5���μB.��bmj�.�󬝓�N+� �"O��"�l��p�Y��Q�L�����.Т{���0����c�D��$�Mg����aQ�M�ݏS.����
B,A�c����>����i.�mf���Bu�zݞ�ͼ�MGQ6�[��v��nv1u6+u��ڱ�0����%Gx�"�}�ő~Ii�G�qt�#ΞQ>(�FϑF��Yn�Nd5�H��b��$�1:X٢���y/�FR�"y��7� �a�ӂE�:t�d,\�CV��k�a�}�i�ZQ�x�rDu^��D1���d�mqʯE�Xт
!�QǮ2����:�~�ۃt.Q{^��kC���Ep��"O��%�Sv��2��1X�utMq�I%#��A�5u^E��������F��l�*�:�6�?[q#*H�-�]�;S�,^�z�	��+�!�n�_��>X�K��=q!���#s$uN�ϰ�<FKwm��6��ә������c�A$6w|�Fّ�$IDBrK�<�y[/e�ZP>H�f¼��e[��Q�r�b5�l��������y�CgwUa��G���g����z����h��f"��񆗤nu`f�a���� ���b����6.��>y�%Z�tO�'I%q [IѺ(   �am�a���[Ͱm�  p �j������gh���z��.�҈׳�m��$�gd���5��Y�61^X�mb^�Bk�[���h�d��]����v:�B���Zɘ��5��jqȰsueq��XJ�]�hýb���7q�7Gc0�7=p+`[��Ol����ݾƫ5�58��cx�v�h�!�6�0�9gs�lW9�Ç^����6�'n�v�n�� ����p�6ә�h��;R��'�[~w�~!I�on��"$�02{f�<t����>><�^����{���ԍ�t�<�������H~H�dv��D�.Fv�Г�!��IA��o<�1�
F�o��V
����ɻ�ŕ^E"��c��(g��]L���H��j����|]e��7�����ؐI��NH�	8�t�D�(��E�{���� i"1�Ib'��$k���Xh'Gլ3����H��CK""ky�a�ŸG�Q;��^	�̑�M�n�g����	�S�<�՟�,i�!�>Y�ٛ�\����T�Ϙou'5G��D:a5��f��,��\�K�}�����%�`�#I�[���.�O�F�{x�Qzl��2�d��@�Q���bSi��r0�$�3E�\z�O(�:}R��R�yg�m�Rܐ��%��&I��Y'VM.��u���ɻ���^�r�jZ��yQ�j��-�ND��IH��_U�n�A�N��s#Oc
#5�*a�n��4oXQ飆Ⱦ���
pWCla�0���:m���%�G�����k6���P��nGC��5��M!n�z,Yþ�w��|��1����{7:�#{2T>T{��|��eEX�U�͢�D���]�ك��ޫ�'�������D�(��w���0�p��DQ�ζ�!4[S�0M�bc���U6�.����v����A��ܥ��p�J-&��%sI"0�G�]n��x��"���i/���S���u."��^<��v"��5k�:b��B6d�1�����]�Xx�9(�,a�IQ8���c���w����x�D�E�N��20�,׬��&�w�2vY�Lļmđ���.
6D�"�H>ݿ�-58Pf�-�������(���l�{�Cǵ��H..��߰�Zٽ��+۬ �����[�\H�oIㅉ4X�m�al�6^�۲�ܯ��Y����,�BkV'+�^��F!�ոV�6w\l�C��\��75�^�/n�������I�$�߾���ce�0b���b*��sk�6B>�#{+��;��[���AK�^u�I#ORyE��Z:ޙ�n"�� �Yѫ��G�C���g"Fئ1�`�A`����z0F�!c{���HÄ�mv(���[]q^�����!y�_ {�6�a�ӂ�Za@���6F��LdYE0B"ΐ�ٮ��,r��Qަy�]^�W��j�_�-�Z���F�Yo/�fi]2���n�g9��gK*q���F�.�\뛝5��LC���z�5�^�;��w<��f����}]vݵS�`WK�\�^���U�R�1WI��r��6�Nyl�fd#D&�,境1�b��ׯB䨝v	�����D�r�`2��e���&�6�Z9$;Wٜ����8����Ӗ@xKgC�l�8���C��Xs�}XED诇<hv$G �@���0��"���V]]�6�V��c�n���3���I�}���-��{w�5�^��Kk�82��3�Y�[*L ֘�6�Un}٧Z��o/-�z^='6��{!n�LT�Z#��mܥ7S�.��V�����.;��T.C�!�/��ʴ���(��0���o��9`<������;L���L��֣!�:!�K��cʺȲ�V��w�ne�@���VS�u�4N�ܿ�r]��9EL�+.51^�9(H�E�F���]�G�	O7����[w5����]��>�.�!���D��c)�|�e�˟d��������X1r��G�;2N��1;-��^�W݋7.�����Y��V���;Wop��d�j5� N!E�5Ċ�'�Z�y}\m��[}�i}�6�v�ٗ����¸?��{B�̔�"��H����
ȕ,�6X��͗>���$ׂ��fE"q_H�M�{����:��oO-�i�pð�q��Ϸ���t�G5":y{6�t��C^ޤy��$U���
�ȹ�olp�g���T���8Y�C����B����5�D0��39S�X+$Uċ!,��1ŇGe����#H����j���
C1r�;�߽�>��Q�!l(a���gN�JI�e]�-���ݎμv�u@v��:���*b��g]��~�����>aWw�r�����7�cB�L$�����"�]=CS��ڠ�/=i�k��[�h�"���>e��� �Z�ħJ:EN+,#ksM(��̇M����9J��I��ֲ[�l.��$�DQD"�ϧ��M�>���r��0�Q�Ϧ������D�m2���3����yN��v0����Y߫�O6�G����\��H҈���(�wMst�F!g�h��H$�)�R�j�LD��_-[Cǧ�y����s��P�[���r�Yv�	�>	x�h�E#{�5����K�i;��5	����I���4a��.�� ���kn�;<�P���/�l�;v�}�>�:�#XX����G��)�̑D�%�,t6y�,�6�����G�M��xg����p����~H��!;��5b��)[8K]"���XG�4x�/��}�GFC�H�I;�8�*ѝ�w+��:�f|�:a�],sr�o[���b�כ�d�l�1�if������<�6A�Gv��k�:h�5�mw��^.t�.25��(O �w��[1�H�$��.�b��1���Lv��ē�8�r"i9�k�t�#�e���Z��Yڵ��b��Y���W0�A8FR�z�e�|����,��o�����-2&�f��#V�5�!p��D6Dl)��Nl�<�7�>���g�"G��t�;�ڥ�Iv�Q=���+�k�G��j�۝k��QhJ�r��֓E��lF�����"���m}���G�h�ܨ�\�XQ�ջ7��/����DH����qr�y`��D�;��HGH���GװD�d�nA�"Б���7��"M�5�8M�,B�=;��_>����4<y��>��PӄQ�TZB�/k{(a�b�!.�V�W�F�C���fG)fA���#ږ%ܨ;��v:�a�%��#�w�yKE�:nR޹�UХ��ٓi���6ؑB�   �@[@ ٵ�    � ����JmF�y�'�OI��X�sv�J6���nm:v��I�P��5�p�1!k���u0�mnm��nqc���{D�t*����n�5�5�:�L^��;D�[=���۬���㋋�l:�Y�;�NU^��y�c�׵'/5�nkVي3��{�|<}�wFn]tE��m%M�nm���.`9�9a��ي8�Eb���p�os�=�D�.{sd��޳�k�3>v`�����$ad��?F	�'[8L,�#r�[�Į�k�ߓ�$jm��+�se�E�OR�X�F�P��L���AR),�I������ޥ�tz��y�C�w��(t�=<��}�Z5�].�#���ۯXI���a#x0lYU5M���2AND���{�\�P�G�{��y�$A`�z�<��'��`��ټ<��q`��q̌�V0G�h��tJ^��<����G��M�(��1�RI���*�b:�`�7.�خ"�i`���<�瑳�B.x�)�@�Z��CSQs��t�����͊��:F���|��+ϖ���Kq�29�?�
Ȟ�X�\���2)5���>�*�3���b�Q>�a&���f���}1.h���:&�;�fl��f}��3(m��A�հ��.�[���ó�����ްnz�����s��(�X��4�]�D1x�B��l.Jg��)���B���Q��Q�,m����<�5��P�~�3�ڭ��im���p��{��G	2FI��|"e�ӌ��!9%�G��==1"̏,6���n`蹛�����4��R���V�޺4tg-d�R��^G}�����u]�r���.
"�DD�&9ܓDZ�<&�4�+`a��(�%�<����8$Y�67��"n��4��g��#[�!c�`�����Pj�#�a�B�B����g��<�i&��0]֜Ȼ`�L,CiC�j��F���i�GֹVܭ><V��,�	�wv$�l��%D�P�|�!D>���������pG�P0�E[_w�'��L3��y����|����{���q�;Y�&��l�#Sz���Y��8���)�����d/*��V}�/�Dja%<�g�ԇ=��P�dQ������P�q�
�Ff�ig[�>�0�$�|�%"ً-����h3�m��2�Qۅ��Py�wD�<�t���-G^a�^&:N�D�0�l7!M4[po:~6y��l��ق(��K	�q�:�zԌ��e��6R���hewz�g�}�H��QF_,��"!��&���΂aÆw�ƑnJ�Cdat��7�_�y4^��ED���\�j��,�6\�7��ޞ�!�2#)��E�uX�(�F��������w~:�%$�&ҴP "��"�#Z6G�Kw)��ߐf���K�~�>��_��k�k3Td����t<{z���J�f�E�t��\�ub�ctr�<���ו�o{:ײ�y�J���"�5��	z`��1�A"Α>��F�Ym���dM�C��GLD�C\�8>V{�f�tW4��D}��Y'O*o!:`����|f��(�$���ח��I̱GǺ�#�:h�cĦM6���g����:A7��e9�,�>����esҶ5�fO��"��k�/;t�Mt���pW>#��.�n{��i��m��V����$�����R�nR���9�v���r���8۫"��H��9d��BG��<�,;�H��bx�����4�C�/w�(}����fi�<D<y;���\��	�*^�רÀ��H�i�{�u��!�E�m�y��v�|Pe��4#A�6#tUp��p�/i���ț.�9%�>�8?r�D&&�BΉ�^dY�<�$Q����S-�l}��F"���9�t���'ӱ�&�a"�0aI�̑f]��k�X�GH�$baܟ�=V�Y#��´$�F�	7PA0�$Y���P�<��7�y��74�F�4z;���:qD^۝af�޺NdF[���'��;����.t՚��X�!%���X*,�*��i6rS�o���ǽtB���Et�mK}�Yp^f���'�Gl��&������᠆��mI%!�#Q���k>�a��6fz������Ͻ�t/��Xx��t�,�T�C�OX�s��8�᳾N��������~�_�L�ۮm��eM�sjoC۰n�'nۃ\g���(>'�"��q\v��N:;R2s)߼����o����{���2,��`��ˎȟ2`�O�XQ�E�tĊ@�sٔ\�hx��e��a0��\,N�L�#��9���y��$h"�t0�$�8�֪���sa�\.��_-E��!��*q�6l�\dk�pP�����,��|ۗl�LSz��7��x �'g�k������4 ��%�:���&�"���B���N�0��wj����Ő���~���\�l�h3W)�Baf�9b�͗=�hW<F}O��ʆ��bG
H2��<QcX�D;V����7=��+�޵�""����l$czKl:>��u�D�(�>ÇQ��oL�_�6�6���X�̙6D��ղ�(�J\p�p�G	8� �1Ky�a�	EIx�D�Gy�ki��Dn
��ڑgȌ>����,��!��mnு�>(�#��`��F���2W��Y�w��H�LZ�j�^5�+Y���}d�ŷ�E�K�P�@��2����}�����_~� �-��   ����M� $���   -��'fK`����wœb��B�7FĀu��{�y��ӛFܭ3C��Z${f�4�m1��:�Cv^�c��β�e��n��9��Q��<�9l��n��㵹��<��u۶��v:������+�ݕX��1y�ۈe9y����8u��y�����#�M�y6Y��u����c�Dv��؎x�{l�[��qڰ𻢭���\�Sn�0��2��£Po��<���C��~�2'ҙcYb10�D_OLN��>��w�p�hk��C��HDqDMc�t�����F!^AE���߇��0�l'!M7%�{LcIb
��$�<�U��:,��s�7�W�$q�(�QD��M�l� ͐�rȭ��\�)���@��u��`�??'�FQnN��!�0�ȩ�oi��{O/��6D��]<�B�_0e?X��[qt���
�b1�>^4a����.[�@������ J	Z�h�6T��۳�]nt��)wk��s4T$�E�Zad:oY�}�q#Lf�
#A�˗5��1���Ƒ��Ǆ�����`��$�8EB��cCM����m�cW:F�w�a}z��{u�$��� u��!f6��Ri=1�Hr��!gϽ8�r����
#�(m}�n(�R�z�N9iȤ�!����u�ɳ���l�ۓ6�=j��q�H��gY��Z�K�[��^-{��'�ߠ����	1"��oQ��[ҘϨ�#JL(�/[\�%�%�oH�ag�GZ�H��'���6���H7��"-	!���L�$B��0�1���w��_���c�6H��r�T��5�i��?2e켕%�Z�IT`p�4aÏ!�G�[��yy%,̡�}D9���[���Q6�9�0cDMo\H��A��
>��葄a�ٰ��L�a����3I�p^	vh�R"�qp�O<E�8e���x�0���GuV���Z���$aqP�y
S�A�4GE���'�Q��l��e)
Q� R$�q���_WH��[l򎐟r���v�I�c	:El���=���O̖E��ܳ�b��(� H���t1�$��w���y}5n0�4L���I�����=��$,�{cz�t�7�3e�_�g��mI�پ5�wB���w��K����PG���!!�w�/�aK��</>μ[J��7h)$-��l$�ཝ"Z���T�\�k1u��t����7h^�ճ�J�ȍ&ΗP��������G۴pWHď����|��lS�k����FQ}6$j�Q�ZCGa:�>uשu��p�k�=��2��1�"j\n�>������k��.1��1-�$g.��em�	����Ȭ�����Ht�i�힊��ϼD�&w�V�
�+W�[�)�Fr;y�C=hW�x+�FD��&l�ݱ��Lo\��4H��gm6'R�Ii��r�!63{*����|������2Y������/)��䒜�o[1X���"�`�����[�к�Q���t�}ν������8�kr���2|���f�,i㻫"�#�Y���7��	�h�4B��0���N ��\/f3p�zV��#!�"O��_F�R,N0�;����qr���tϳQ�2[t�-ͱ�*�[D�#L��Ȣ+�oesg�
"R�V챇��NE��|xu��)��m��H���	n������!�ƽ��c6{M�cv9:����@qZ�C�# (�Z�(�e(`�0��k���u�޺�>#�w<����~���#��d}߆��N����=�g���\g�E�!4`��W��K8�b3�hv�#����aE�-��1T�����9�F��q�r�E�/�3�����ΖB|��n�"*�H����9Sٳ�����lV�{"a��jF�l���|����������<p�"�����v�q�6��Dmw��=/ND �K!!b���͚����=>#4u�SK��{ؑ�E�,a�O�hQ��'{	��l��"�s�@���8Ec9]עE]>�L�6��k��t����d͹OkG�ʕ^�T	�&ȷ�5��;V�һxb"�8���Մɒ"a��M	؝���$�wT3;�̅�i����(��G���tx�h������}V�l_{���n!�$I�=�"�a�(�p�~�Bp�FJ�>K���'4*�£�B�NE"�`���b�3��
g�Cs��-3˝eա�擷9������6�lo�����w���1y���,aӍ!��FEv���i�0�HO��F���Y�GAC?���ׂ�<t�;��M}����[IE	��J�>IO8��l�k�{Q"��Z6W�2C����6+��>�N(���Y�ߩ�E��l�d�\�U`��O�=ϻ����ڑ��_$��N0�$Ö"Ȝi#�e�l��^�f�af�v�
I*�-��1}��;�e�|EJ(;L�[{����#�����AƠ% r"�.
|D<�>��<Z�ѓ�S����o5��P��2th�(�>������p�����`��n�p�!�:]�\��zʌ�`hHd-��;�Daȉ��ӫ��|�F	���@�n�j�U��Q�O�����8(�9�YO���-7��q	�6C�z�����6żH��jt�S�fӆ���i�x(n��t:9���q\ojw/[p�7N���,����J����؏oV�x!�Z��_u�]�H֮���j ��ή�p�N�`e^|tK��i�/6�6�Wu��Ws��؝�	���5� *<��Ygz�w������r��g��`�O��e�w���!��U��b|�vbǹ��N��)�lK��]���f_}�3�
��:�����XR�q:����Y�;���y��.��8З�&�ƅ����5�v�ggay�]g
��Wq¹wƣ�2u����Ɩ왏/�sV�'Z�/�c�z��R�Z:)_+�7sR}���od��U�+y/�62�.uu�w�n��U��se�8�=Zxg���p�!#��L#w.��O����U�zZ�}����t�ɡ[e�i�۬�=�0�-�k�VĀ<�90��[[K���ջҲ�7��[0��IN�2j���t��ɻ����&�{7��.�#��
���ѓ�v(7�#]8�8Z<%���@�ʳ.O����wi��M����3"�ӝ�X�iF�v60K��Rݖ.�B�����'��ڴ3g.��y�IV+Q�i��c����w���={{��u���       m��cm,�   m�  ��z��wm�&�m�        l        kX �7j�`    �Wn�      �`   �,ʩ0q�e�h      �      ��   m 5kZM�   ��  � �]7L��ݷKV�yӜ�ת[��U��	�t'W����]j�g���yیG1�t�Y�u>|T�:	�3��g#�3M�g��usۮ���x�ł:;t�/Ա<���p�1Y��>��88����m�Ɯ���r�v�Ⱥ:z�I��'���r��ps�z���ŀ;�vnY�H��/
9�l��y��3���Q�ۮÑ�����8�b<��s�G#ėG`^ח*�]:Yze�����jS�)q��fw\0�Lu��e���n�)��q�l���x�y+�c;��{/���=[��+g=r��s^Xmx�5L�M��.�����������!^ݻvzy7[�q֭a��y�G���"�еFƽ{�/Js�/0����tvT��g��{a�+���s�ݮ��*u��/[�wi�L��6Gs��JG�ס���f���$nv��m��Nt�c1�9f��;7+�p�n�]$�x"���� ��(����n���F�Վ\Y:�Żn3ig^�<�Sn��,^"\�X�V�m�7b��Zs�8�Ǥ9�6G���ɷ
�<����'��<w]#z�u=<wns�� N@Aat�.��� ۮ���d:��{<ۀ|��n���'�����l:��������ʯizk��[�^�E۳�W[�u��g!����e����k��in��۲-���T��k��ۧ(�=�ݍ�tpݭ��猆t������'t/Xxh=����G/�Z=W`O�tW%u�`6 ;��ۤ�Ɏ��lyv�Y�{�M:�׳NM�3�l 	���E   �m �` �   �  k�k�n�#��{���ڽ�.��=�����I�-��\�n����xo;kq�g�[�=�宓�������5�i�櫝ma^�%�-��m�X����秅�v��T���}"v�q�d�����E�D���lqq���i�ޤc�GŐ���iq�lSg�7`-�/;qڼ�g��*'�nծ)ݍ��;C7�ᶺM��7Y�m��[��f�nr��+�[��䃿�i}���4k��
⋑%������'�'�FKy�u6
�y��`�_+=�N<x��fܮ�Ay��?���v����i��RI�!#Ǖ��]����ue舭>�8�/Ե��'�I�����Z(XM�Q�$#;}q8�nޝ��:BƲ�S9`�sa�Aw���*6y��t��ׅ�H�+,ѥ�q>�a;	�D�M�3/�����X����Gw�,B"7��>�����q$�)2Gc�.������Y��Ϝp��u����8EL1��$*,�e�oZh�3���tE�!��Xu-���:X�(q��a��#����@�H�hENK�B>�b���{;(ah�M�7��#euRn("H�[��yT���0�6F�JB��0�� ���J�M&�Z܄�܄�In8AN� (v8�3gq��������v��i(���͚����9:<A;���>��?<�(�&�u��s����(�lW�nJF����Nq��2&�Q�a�$7Gp$�(�"l"TPW0�p�"�{t��9����g1]��͏V�݋�7��eeM�����`YR����f���WU��Mớ�r�s16�w17��F�$��tWH��<��nP�ƊÅE�wM
9�'ֺ^��_>"*�|�LB��B�Q�ht��U���D�}���!��ɛ8C��vX������t��WS!#I"��I�N-y'��>�7~�ĘI��E@�M�|�B� �í������Ȑ�#�*ٺuq�"$�]��4�V���Ȝ�`�*$-Ψ��D޳�E��8��I.�P��e�,wŵ�<ydn�>��t�h��l����։��OC��d73s!��p_0���v�>�޺+�>�x�w���sO�ɮbm�&�		�j{n���d��q&n���ɹ���ю�nMɆ�(�q��J(S���_�?!g��X�la]B���#�}�+���Q�|����m����^�{�r1�܌�MBu�a-�>6h�����I�a�܎��\�CƏ�#EV�ajh��q˧����(�j�[����#�X2R�	�$�0�`���I�Ĳ>�Sz�T���:n��Y��i#2#1ɜ��y����{iv�bh��)��-m���M�i�s
�ߐ���n��D��c1�1I�;n[�թ�	{�R�+���o.�		�~M�jHVv��fe��/�Dv�.��~\����G�����.�z��<Fn7L�ga�`jG^8y��g�Z��B.Or��~DI�%3�(w�9��d�>�'w�'�C�#Z��[;�)�����I�+D|}�<y�>�����$�	L�XF%�<�D. �"̷��Pè0Di"�^��x��}��4E�2GL��޽��z�1��	0F�v	�:p���g�Y��z������C��m�c��l�@*�#rbu�&�<س�1�9��l���n׳��٧�}��QF�:V��}���%�f����X	��{|>�gw���3�|��;���B�㝾�#�����+�_i�0 ӆ'&H,a��Q$I��O7��u�qGuN�޶ʇ��	��!=�$in[�==<���hV.`�0�A6�}��T=�u�h���0�y�ť|	|��	����(�:l�>�&��Z,� �'�򷞆H-��4h0�F�\0��2G3	=8��׳�0�Fv�C��fPc�QG!e� �x�6F
�X8lQ���h����Ķ?�ɭ޸�`(�]0��WOtHdޒ0��V�����L���xUrB������-��l٣�We���WY�v���8�9����p"��(�T�=2	LÈ��_�!���^B[qD.31�C�����lO�I�&mJǌ�s�撆C�D���q�t�����|���,�qn��C|����:B�_|D��6\M��6�A������:ԫ��䖫���	i#��I�׷Y�]fq�j;\λr���������a8�of�lH�dQ	��GGI�>� �8D�v.��Ml�Ɉ�����H:F�&�D3K��(��k�h�v�]�<'rP�A{��<�e��ӆ�8�K�yV�w�Ki8�X8yX���lu��EΑg�ї0��;�����
0t�5��X�.<40b�"��K�E����]��zFv"O��EQu��duW>��s�K�Y17�XBf&��~�����(���"�v-&��'
�Ac��M�-����ꫣ�Xw�y/�w�ms�����+�
"�C5a3���Y��������N�{�o�>�h�q{q6Sl0�)&�pW;�Y�j��3����B;A��4���j/!�Y�E��̐y�m����ޒ0�6l�o\I��Q|��$G��$����M�OKG�eΰ��d�ci�d̢��6��SMZ�3qZ�����U�c]]�HՀ���۽���z� H[Cm�+`  �Ā5��  U�m�   �cmͫ�Z���⨍v�W�w;6˱��٘��'8�V���'e�Շ����tC���#]�r�g��������	�ԽM�K�Ikj��PHxv�=��FO+�u���Fx��r�v�����=8R@��t�W7ܜ���3#ٮ�k�����۞�S�,�t��`�jY��M���		��Gfz�h7h���]��ʌ�Sl`�{s��X:��T�2In��6ӓ��>=#Z�o�h����#�������a员�4F��1��̑���\q�g*$aj]�������Iᑄ�J(T��#-"0y����#�Ff�V�f�E�Z�cyD�H�0�4ި�T"�1C�#�!?	�4h�
�3q�d/9�����ά���(S�&S��GH&�<�3��
�6h�MAN,�ˋ���_��e`�:�Ee�!�諀��ȹD9e_Ժ+�:�D�#��������M�Y�	��Ds�e���>(�|�F�4�E�vp��p�[Sm��y}DY�t��e�`VWX�B!��DwH�ԐjD�2DeI(t��xޞ�vV��������E���+�b ��kﷲ��HC��T���}Xa'B!F��}�u's�������m��v)qX.P��۶:�<�g!��r�VN�z]:Kr�*��]2ݷgy�v��}"O�V��� �!��y�/�V'��,�a0�~����t�����ا���2c}D���<��g���Z�0�pH[N��F���.dV�dW�1,4�袿fxv_��Y���Wdss3i@_
]�w/mB���\tPv��� ���=�t�7j�:�1��<����5�vP�W,����)	�Y�փ�2�K������WJ�x�/Ð�(�3�Nφ�������"�0�F�_J=�,�}&N���~�1*�v�S1���ۭ�3�KX��sv�s؇���d3tG�J��'!I�$��3da�m�~�J�V�<^�HMĳAbL�8c��|�wY�8B>�ONr(�ƌ68DEm��>�1��L��#�Y��#���cE�����=<^B��.�6����bc�Rj���!�%���,���`�Y���z��q�w�G��|͔��ڹ�&��e>�LȓI�L���<cη	Ĺ���8�۱۬�OkY]�7m��\�NqD
HQ���.t���m����!�c�D�i�s'�x|!#�zČ��:F"
m#o��N�}b��~l��zױ� i�ąHSNKQ�/G۶�O�/�$a���J�@���im]��W�XA6�G�1��,���8���$Y��[��4�C���a����rX��#<�D?O��:��O<��{K�C�O08{9�P��+j���7��	tU�mos{H3$�����^���c������ǹO�f4��,�"+%F��*�$1��B��]n�><)<�mφ�\J��_2�<�&�'����ч����q���'m��B�	��<t�>���qr8E@�>).mxf3�b����6l���QpӅ9�@�PP��0��$[��v�JJaf�X���ș�}F
>�`�`��g�8�6j��Z�	<��a��．I`=8>�9q;1[m��6t=z
m���{%���֮��]��]m#[A�m���`kw���|h�_�A:�ګ�]8yM
�|��w�|�60��"ˑ]��$&���>+�#O(��܉�!ȃdI�F�fb��,"%nK<�0��$K߷�y�ޖj��*Α�I
�뮒1s�<X���+��II�`�⧢`�_E�d���F��{����0�P��X�FK�10��,��4D�8X�E�-��e���f�o)�zF�����D���]�:G��_
Z����G�t�C��
|q�[1�#�$�H��0���W�:p�e���k	>�Ƹ����G�d�h���'��4ȄB^���ݦw.P�oY����}Nŝ7jf��sk� �`5�)1;r"��M��羙�N`����ǝ#�<��e��q�d��\���D�K���g�E�"N�+vݠ�eb}�9��2PvQ��:Bfd��8h��94��B1G�ρW�n��glml��+�ty�v=\r��w[r<�d�X)�7���N�lVW�vWqhtB|�#�I
7�O���Zaf��g[H�)�%;bo^���	��z�nt��.]|�w�s-�<�!�dt���u��X�H�l8+�C#�ou���d\�!�DoF!>t�9�(�jv�Df?��#���}��X��`&��l�Z�e��GO/����P�	�m6���.SD��*V�dO�|�a&
5;���wu!���!WG��b��t�,�a#�֑;��Z��C4G�<���IE�`�L�_<~�O=��4�)]�"�.�J|�M����;�U�
�bìa��z�B���ȱU���D�UĢ	:Ee�>[H�H�r�rJ#OK5,(������0h�d��+åӸC��y��FM����(YG��al��\HGӲ���c{�2@��{�gc�ݒ�Vl�gS4p�E��%b0S5�ņ�.��#=X�az�6&�5�uy�c��l��I$��i$I$�   �H�-� [vMv   !���n���y2rPdd-Ԛ��WL��rە���k�;p^�EvճH��<�UӦNn7���,ՂUv�s�`R�#���%��G=���bwf�f���SWT��7Ng#r��,�v�n��v	�qt�a��v�"��s��ppq��z7cq�[+�X�ڕ.l]6$u�6�n�q�1y���#��r���ӓb�Vu�R��&�bBʒI29��!�ǿ1g�v�
e�-"S�!�����w<�ݎȳdDOLH6b�A02�//ňsdo ��<F[��.�F��zD\���j(M�Vp�:B��h����]�����Ӧ�θ�ԟ�p��a����(�<F�'m��=M��K#�؉Øa��3�荾����;h��w��n���D�A��葇 0�0��]�P�h�0���Ck���	.C�ry��_ٍE��7վև�T��Y⿻�D��!�0>-,�0GЦ�����K��|�W�ߍ60����-bE�A��"wz�}�9᭧H���k�p5�V��K>�H�=!���C,�cq�QH8+�~0}�I�z�ǡ�Y�a�1�f�ml��\�/��Q���,�D_m��ɘ�<�9��M��g����|�j�`�����Q8�m�֭�F��
�;a�lvp*��p�d�u���M��k\i����Hmn"�����a��p�DT������,��=�/���6��.�Iy��|��|�x��0��у{m�0@�I�/�/��1��vn�P´�cp����K��Iigp^b+>@��ٲ���v/p����6���wG�Yx4��wy�z�ӿ��>�'�E*F98n�k�&0�w�/z�$������B�{J4|�#axfE��
�7%!�#��>
�\���&��D��y��ÍV�lg����hH�Ʌ��5l�O\HG�"F:~Ǭ��,H���r
�6y��M��v�^ �w,c��#��ѭ޸�raHDQ�*::$a�.Xak�q���}=!p����x0Fi��0!�ȯ���%���f׺6��}�v��|�����ٴ�����%c�?s��ڝ���u�VĀM�l���K�ܓu��2�'0����Xy�dT�9�(�\���iE�I�fs>��ފ)�:�;�O�asf1�]k�Ѱ��ƺӶ�X�q�>ˣ� �I"�nՐP���{�Իt�7�DS��¨^-,{ؽ���Ն�Kf�1�h�%��E�;A0LAaT	��F`D��x���kyJ����kCDX�ٿ�tG�c�����:5�F�r������x����W̑�l�t I�i�w_]��۷���N��8��t���"�VY�<�o�q�n��޴	����n�_�yͰ3 t�ne%����ާc�K�ι���z*�����%=[@'X�a�HE��쮧Y���n��C�)��u��7vbm�jH�� MA>��u3C��˨��a��{���eo�
Zk�z:s�ĩ���X&�q*��bR�c91��S*��'*<��-�F�zɭ\dծ���\	�H�9�c�섋4�1V�:pl�8�]�}��]-e����c�=�s���1�n�k`�'J�՚���(:�ۘ��øJ|)�������e6m]��3ɑ;�������֕ƨnX$���t�:�鰑�[S�}{����gVc�}\:�3�X"��V𜚎]l��G�ڨ�+���̾�g`��o�Θu�\��Q��ᵄ>y9 ���ە�v'w�����Ռ��S��dm��=���3ɰj�Π���e�.�s�Yq�3�f���oLhЦ9�v�Q|�=Or�T��y��kv�B�
�+�Ym�`qu�sr�[맅;�c�m��γ�qg�ȱyLW����\;N�a�e�	Z6H%����Q��|f>Hi��g�ŕs
��Vm<��%Rc������޷�n���1!w@�H!ue*qڎ/w�E��u$�U��3�+m�c{٦�Wt�}2?56޽�~�+#���%��f����D��8��d�vi,k�����5m�2��k��5���/j�ۯ��(�^՞ux�hꔈ]�1e
��7�YBs��B��,�g(�Sw��B��@�Q����f�̋.����8-gT�ٷ��d���]^{�����vf�����
K!:��&�s4J�5�	]#wF�*VR1��#Y����r7���6h�����o/,�ǵ�0=���t4�߆TIB�h�5v
Su^��V$$�7ڞym?9����mt�\�]�cu��v1|b��y�������X��P�W]JEZN���]9d�8�� �jCs�h�C&�/I��+kk>�AU���4(XH��'����1f�|r��9�{�;�C%���Ⱥ���6��40z�(�i*)]��s��ƽ7Zt��Ѯ�n�ҝF�hy�s�[���]'j�lr��ֹȲu;����zo�?Y�]�=������K��zL�Kk�k[ͦ:�_��6� U���I�>��bmd���N�>y܎���x���b�:������!�[�"R"��AQ&�U�zg��b��J����sz|S���kP�o.[ޯ`瞕(& "��4�$���7=�g�t ɕ����4�ȝ�3�}�W�_��Z����o�9�F:��b*	��U�)W�Vp�Ǽ�/0��;)W��Ȉ}}�&jnwF�k��J;w�
7�`���ғ/�oh��ɁHK�ӷ�����0Խ[����n:n����~��f� ��ŽV�5 ���ۤ �J  ɶ�  6�;k5  6���v5it����*��mךWlݨ�Ĺ���͸ne�r�WU�6��lr.s'h����k�n��s������m�)xr��� dz.غ.�r�ҹײ�^m���8] %�c-��gU��� ���,����/�����r�]`%[rm��	Iɯ�3d�9������={���&��y��glIù���q���V����Vx��>��B����y��u-Q��W��-�Z�2�w����ن��p�����@���J�JYm��w���SYjۋ���M�����e��g?mB7J^�S'hܺ^�b�*�
��V@IA�h��db.�y	Y-�h`(�}�N" ;��ȃ'�fyIU�ViR*�eV���Pǅ1�N��M�5�������{MI@�h��,��l��Cv<���#J��IZVH$*��ｋ!'��L���
��^۬����r�H��m{����~����{~�qs�X��4R�!-�\�K��'UmoK�b*��q��H���9u�m��]]�m�E�t�A%N(��>k�J������b�6��6��{I��{y�c�1L0Ktv�O j�����I$�Vo}�ܼ�r���n�lr�w{�y�[yEx��A�M}���.�vZ�8-1�̰z��w
�V�T5|]�YB.��o�kbzS2
n�����a���[��)漺���h$��R��J�0�e�m�{�%hi�ew���ٽi�;4�JxT���<=GJ)|M��Q����d���:5�?zOz�����/��+�{h7۽� �;��ᴞ���W�F�VAE�)`w������]e�iΖ�wB�y�{]5�Q)���dO}���ֲ� ��QJ�TR$��lN�nxz���m��Ź(ы�������꥓��]D�D#q �.$�?�Q��`�I���1+ڦ�ލ_���خ�k�E���JC>_"{���I$$���l���.����{hz�����~���l�ض��"�x̋���i.BT	TF� �8#ZB��(JU���{�ZWx]�ϟhQ��$�9Rul�j���]Qi�t	MR	QӘUI	��q��.����t���;V���W�l�~"H �J�V����o�0v-j��.O���=#}�2�<�]k����'ڼ�y��� �	RD�	%"���ާ�!��ۙ�X���xEf�������Xg���J��3G:ܣz����M�)�S��d"we,v���ӳ��9ڽ�74vsLn����iʷ�m%�,�jJ������~-��{�:����Ch�2�X̨�ͻ!���v���$AE�����\��}�-R�$X���j����9�U�)�z��rv���g��"�$PB�
[X���ٓ��0j}eYb��D�:������^���F.�(Ր���f�J:7��3!=Wk7ö�+6�S5�^�"ʌ�趝�x���wr^"�6)�]騌9�0�9��Z�n�n��4Wm���ےH�P�,�ad�u�嘴�����j��3��f���H�J�*4�V	�����YŞ2�9�G�W�r|�[�3�$��*�
���u�ګ���m�s�|��%�Y�ms!^����[t��jW�%&�ka�C��]�#��8���8�秶. PJ���~��H��y%-VG��=���\pb[�Nq;�����C�iP6~*�B��T����`�;��y��=[&25T-��K�[q���� �a��q��U��m�����l+7��;+]�ዘA�r�ю���ݙ�u����K��do�A&Q��@J)W�k���L�ԅ��Uj�.�U�P�j��ز~�1��ym;��:��ՙ�z벯Q�S\�
�� ��(�L����1={�*����X�-�-|�W�Үz�t�/	JVV\��;��������D�v�$Z��3"�T�K�7�i�s.s��s���-�s6���z�<�-�d�>���}Ϗ� $h��    �e��kh  ��Z�   � g^ȝ��ٗ�u��Y�mG�kk�/�y��5�2޻�ds����5Ɣ�s-�cI�Y2iY&מ\`
�;��XU��x�-���')�K�F���Hmm��Fw0ֺ�t��5�ֲ��� Ŝ:!�h�κ�77k�ۚ���l��&^��-sF�uJ��M��m��y�B��t�ը-J��rc�,c��`��S�W;��L:6��n�$$]��j�ݰ�g��xe����O ���,���9��tf-��`����O�~>)$,U�*��$�����YSr���2��X��i6���N־ʴji�{�����~��3P_rX;�[H)M�Q�Vc��t����F}�����wBW|,$N�4�5=���[�k@,���K�JT�
&���E��/cj,:��������Eo)õ���y���^*���7I����I������ɰJ(E>����m{[�ݖ��k�es���y��qB���/N�k��Ⲻ�{��@@y%f͕D����pؓ80���x�-nn�N/8uֻv�����s��{b]�k�z������{�=�S�bpg+�3�mAs|ͻ��ف��ч�3y���˸�6$$� R��2����~�oXX��×�x`Or�g�/4�Į����>�%�))�������7���x/�WLtz��{�転ԲF]�����5fc�����[���Ή�5�˯j  M�J��)��U�ţ�BVx`��vg��/]�U�Yr	�e?_���T�z���[u� u�������n��^� ���ȵ�*�,�z��O4R��;��r��jnb�u���z��,���$Ii ܀�f �qb����M�~�OvY�#���U���2��|;;>Qav���iY4���[�{���}�~�=i.�6�W[DX�&v�����.���X�պ���5�����^ݸ��ٞ*��T�%P�d���wf
I�x��������V�3{��{3#ܥ�l������3겝��Q#C�����tv��yJ�� �����9GǗ�<v���3kD���׼T������ϸ9\v�VM�6��.�H?8���dd�������U��F��˴�h�U�o��¶�hZqQ6���xh�y���՛�!��)���oQ-�Y��,t��ë��~<��T�b��z͚?$h�J�I%����wB�/���{V��Ǟ1���ے�:.�����m҅w�I�B(�E$�c�gW��kC{Oo��x.�|�+�[]�*�{�d}���:���D�����{����Y��\��d�s�������<	c<P3�'�I���`d��[�+��)��/�OR���Nw���Z��Q������c1|ɽ[�Խ�</w�j��Ud��R^���a�Ň�vfgL�]8,�~~�w.���x����������c��ʺ�:��RV�Ք��? ��Ҷe_���ܬ�0�^��>��>�	y�~^�����6�ٱ������B8m�T����>>O�+у�������S�/\w��/-4��!�V���7�0KV�t�eH	�dD>��ƙ* �-l�3J�h��P-�pY�k+�e�8{#�w���׽~��r��!~�@�tM*EWI*�%�KݞR%�k�g�z���o\���Q����8sv��zC<v>5���?o�� ��~������61@v�-�E
�ac�L�7S��Ɍ���; 
b �J&�Em��;�R�mOE�U�6��bq��ɷѳ�0; �4#���.�b���o@��(�� ��fx/z���%mVu��v`�.S��hF~��3�?/42Ü���"����P���5����jT9f[T���?�Mc�n�Ay{�MvX~ۗS��kx�j�yu��T� �IFud�i�a̾�vu̗��z+<ד��ߣ�ެ���I�)�z���^�ϗF��m�$* iR6�ҰRإx��~��z�i����G�y���x�ܭ?yץ�n^j৕U=��' �:���W.E�e�7m
tْ�j��ӡgm�;�������[��ۓJ���w3Ae�W<��ccr�s���]���T1�)����ȴq��t�]�􌖥�gLS|�˧�'�:�L@v�r��;;7b!O�8U�{�;Iô.�����]�F���M�S)�Y�N�܌գ�Ef�
N�Վ�Q�)��DQh���ǒ��o�Zn��l�ݬ�E�]�]�WG8L�<^͂Z��p����x��޳�p��]�3Z��/�G��gV`cM��:�J�kB�;�4���f�(r�n�v#���?�b�uɦE�x ũ��+��{9p��i�:=Q�s8hpb����zC*U���E<U�[�W[��˾&���:a�V��#�l�P�YD�L�Nu���=,�L��G{]ؾ���ۗ�/8e���K���[7�Zޚ��kI#j{.��oYN]�gS���� �A^J������ʽ�6N���Ω�m,�֭�^��z����e�Ԯc���~���H�#��he;�\&f�m���43�@g9C�	�]�%�4�	�b��u��Uݳy�Y�ċGp��mu�Df��|�fN"�w�i�#+�^n�ms�R���$�$��     �l-��   H   n�݀ҵ�`հ         �        �` ^�I���    :@���m�          �e��v�޽ڶ                    [Cl��f��    �  � �ft��w�M̎N��3���c���g���v�<�1�5��t���v�j�j�6�݈zS6瑕��3+#]֮���e��X�m��������\�FѺrx1������5x��gc\T���f���s����M�1�º��6�x�)W)�GQ�jD���t��N��RY:vkR�E�籼�6��45<���bܚ<D䮛q���z]F�gL�:u���u�];u%������Rǭ��8�O=�pY�[��n�a+�} U���ZR��`$�>���\����=��G�mq�E���O���!\�lO	gNo6N8P�Σ!�ۄ����*;ti�Zڬ����M��>���F��E�kC��T��9㶎ͅ�^�X�;g�F�j$��g��ڸݞûn8[�	=�k��v�y�q��8�e���v6s�A�q��@�eV.Nm9�m۸�,Z� -d�-r��u�/c�5��N����6)�˱��^ͳ��rj�=�yܻ�xўj0�r٧ю��۱=wg�NL�q�<�{E��䝸x6����男Y��Ty�G����vk0�ɤK6�a9�ɣuU��%�Ju�m�F��H��H�j����ysqd��GY���n]��;9�㮈�7o+�,jp�cO1@ؕ=-,�v�O\nX�%�����׃d�k���\��X��:q{�'#�>+�g�9�|Gk���}��#p�����*��q�����Ӯyzy6�V3<<8�9��ݬ����	g�=�Wk��]� ��n�6ݤ/\8%�ι�[l��;Wd�W37d�	,�u�m� -h�m�   �Hj݀ 6͹�   5� 6�K�K�t�k��'c�y��j�d��mv��7O#�d�9&G�c���k��>ۢ�z��y^B�"�*2%�v�N�m[�u���p���ˢ�&ny̜��3�K͗�nq�St���z0�&@cΎ�=u��)�cګ]b{N�݌�����v���3���Azs>�Kْ�r4\��(I�F&ݴG�,%��*�mS)'#�7b�+DٗoC���	U�J�t@)3��>���J��ל����5k�<�����ިB��Yssi��U��A"��� ��u��IyC0]<xt��nyq~��`DO�qb�w�M�|�|7KJ�{�+�^�"ѻ!]��D�n⹙���.M�}�}�fLu+@b��/+`�g���&����T>7EX&��E����=C��]_`4rV��l��[���VN����9J��	�U�_�.9���j�����DՕJ�	%��g�כLf�.���%��a)@k�οk��V?��#�{�;��+����ۮm���c���۠֗���e鲜�č��W��=g��=n�� �_iR��I*��+�>5�+!76r�Qu�:��yc�&��5�pY�\ڙ�O��	B$F��E7d�#ʁ�˧�sE`^\t��nf�j��Ep�����CRݺ��.;��l֞��՜�B�i=��ā��h�u��u]�9�n�Fe>Ӗ=�+��s�t=Kv�ڥ��xV�ڽM<�w�XEU�.�I;�=�$��<���?CH׻�6�i�8�d��ăx���6�B`�|G�ThU�(�~%� ��uw�Vb�*ܐy�R�������}��dۋh���Cj�mB����+#���!���2u��E�:��)y{�F�gn��R�[�z�5���F��f�׆A7s<4��x�6�o�mr�B6�]y�n�SNù�s�6p�[W
��:۴�S�AnSvZ�=n���U�dl��,�h���s�wx9_w>7��+ǋ����0��dt�(Z�aA&�ՅV��JW�+�s��֥��"������j:�j�.4�)�c�����͵����f7?v^ D�(�H ���ñ��Y[z/�ž��Y[^u+�K���n��[�̏���3_^����%�K��{�q�᰽S3�}@U޸^'۩=�
������y���K�{1�����&�%d�e*�ɹu�=|��v)Y�S�t�~��U�)w�1�M*�ؿg[��ĭ��5��]<@	�4�Ĕ�H�O�˧����jY8:|*���׬P�{k��h���ڒ��YT4S�:�g˘�`���9�f�x�[l���aK�T<�=:�Kg�Xk���xI,k!��x�ZG��'M|��et�u�{������>�%�f���Q�c�XA�/F�w�mk�}�qV�/UL�*P�'�y{=���1�˧-�����M�u��tڠ�&�Tl�UJش�e���)Lū�׊�fU�[�w{u�+>Y0�O��u��C��I� �ZJ��Oס／�����&��������)�䥬�(c�!-��9r^C��p[��Y��=��.T��u]0\�E�O�;�L�@�J1���
/����K���ډ�[�^o��>/�ØHI+ю�>���W��@�>�7�O�o<g"�1Cm��1F�jMhۥLc]n�����oP�i���Hӯ*��q�����qOmcW7=���6�������w��|���h���� �P���N���cf&d+y���{ W�*m��yB�2(4{�7Vh�$�AR)$��!7޼�֝���xx�����T�F�g�(T��Ku�pX��5=,�[|�ͦ"L�p"��6
VY):8�p���خG���^@�Vy��"~��y�V{7��J��F�y��k��=�7�
AD���P)-]ϲ�
� ��dO�/73z�T�;��=�ή?d�Ë׫<�-���D��Q�J���ҧ�#�u��Q�KN���Ȟ�[��/,���W��3w�u�h�qמzk'n�P��yu�O2ŏ�M]�
Ln�J�v/`ø�S��͝AU����W��d�6��8t������:@ �`ڐ�( u�k@ m�� [lr6ާ���m��^�5u�s��3m_�}�������{��:���q�f���.��6��\D�[�跦����-�<�8�k��X.s`�u�:��+۲\�u���.��N�r&�^��lE>B�3�����|흶{9�g[�1��*�]�CV�a�`8�EL�#�l\P�#m����U�l�����ˌ�:s�I1۫d�/K]�]����G;��O0&�IH/�M����)���������eg�A�t�.�d�u����Y6�uk���;����j�Q����?-,��4(a#���!�}�I��=��O�h�4��n�O�]�M�TU� ��k��d��<sV�z�K���Ջ�Z
ģE���i*jjŌ�F��g�@B�)d�<�mTWW��j�r���8oSG��u�������j�p��~%���]��z���_�hn�(ZVJ6R�ܮ<��Ԙ�;�8�+͋4-�y�x��WP���F�mx=���/�gR�2��y�TE���		�A���/M�in���aL��a'n]���Ӷ�#������"��?z���j����ַ8�,Ly��;V�yEƄ�A�������z�[�z|��@�
@�V�%-�5���*;��0V;��Z��֥cr 3�k�b��v���6v�Z�n����'rY��!+�zr�4����{fd�}�j1��=�X��Σ��D?��1�Ci �-"�%���+۷�mK�yʔE@��>��k�d���E����Eڠ�$�T,Ur��m����{s_����\mj����í�˵n�=xVLYճ%�~��+&�@*�T�UL�Ħ��yv��/}�m��?ZE^���ƏyJrRy��R�k�����k`��Sm�A��� �U;�����Qc���Ń����Ѷ���mգ�5ђ�v���f�����J_���9�}�T�7��+u���n�>�c�!W6z�V�I/L�gw�mm��8���ۂo��nx�A�Y��w5��~E�b��Պ|���u`רY�&���IV�Я��Tf�|�3���:���x"��`!Cb�����̠��M�]s�[}�U��*�3��H���a���%�Ѻu%�����Ft��.�p7��Vi��h��Q�6Q|	KҲ�����&��x�3=~�ի��!��+�mI�[ܵ��!��X�.�P�}�߂�YT�Gvyv�<�a�/g��;�x<i�e:�ϖy�-a���/4�z�\(�ц#�`�s�l[� =8:�cUx��Y�d��W<M�����rÙ���յ����	-�ge��ked`�N�}^yKoP��zc���.]�A��]b������yL�|��$�H�!m ��}��gOW�/�W�ٖE˲���>9�2��ŕ�r�v����evCf�#h����kV���ұDڤM]�Y����-^�$?/�[0M��&-�"�졃_LK���}�9a�� $ѫ��Z ��5�*�o��iX�M�ѕ��6�絇��)B%��j{�B�~�"��aΕ�
�6�#E�^%�ms�^ekJ������ڊb�0ȳ�{-&%i��o��j�@~I`�/+ݾr�W6��{�Y�]����������xY^Y�Էc���G+v��VM�넄�)�ۢ^�K�ʔ �=�����^��[	�o�_�)�v
��@�m%Z����~؃'˼�קs��c".5Cc�S=�)}�w|�Ȳ�S���$�N��P����o�i���������%�V/J��8��f�ee1�F�n{�4O�4x٢H�(U�IKT�֥��Ň&���і������p[,���XC�x�#��_y܅�A�ZND+e�(�>l�غ���5ˍV!����V��G����{�+{N�4�u��аP �4,Y*��q~ŞJ7��":�+�Mg��p2�^g5�&�Ɔն+L��*�j}�Ԅ�Y1��J<Z����;���jm�L�3�Qxfٝ�����r�M����)����}�n��������B�-��ͳ`  �����z��� ��`   ր�l�W����N��ln�N+��+�Z��meͥv�M��h��v����j�n��݄�Y�ոܞ҇Ga@�Y��<�U��n ���"�h쇖�R�V�ܭk��[#����Y�qd�]UsrS�Oօ�c���4sn�oUi5�:Uڗ�-�M���ݪ�N����vlsã&�x�ɞ��4��Gj�q�m��:8s�;�Y�P(p�a���	��.���2gS��^�d{�3i��ƫ���j#x��Y�$��R>7EX諴���6�Ɂ)�b�Ll�t��֥�H�%���{�쥜�_�ny�_���b���h�	|��!)���������x0���c���r���eo�V{v�V>�,��5^W��@� Y�eZ���Si�����6z��M�^|�(�yV�x��ל��>
�\���j".]�h� e �٠����I������s_����Q�q(TW;���SDj���in�o(��eA�{�{���ZTI)Y �	;��la\b.)��!V�<js{7i�W���̩$E"i�$ZI-u >m�x�������>�Dۦ��-Ν�M�H���������"l* ����	)��2\��{��#�o�wm����Sͺ�N̕W��Ыv���]��b��tm>�w��B-�j�ek�KY09#���P���r7Ǽ�����=�̑�Rݭ垒��a��n� ���T�#��ҧ�/(��n�O^l�Y�Mڻ�{zy���Rط^5�L�N�|Y�C�a�]�?���x��g{�D/ţ����]�r��%U<����ǋ[��yk��#H$٫���D���Щ����^��^��\%�:'T���s�{6�^��~�S�/��x*�޸T����V&�j�a!��Mf�㎝vE����׮���k���B�ˤDطu�ͼ��J�����w�ּ[[�y0�C�=���������{2$'bɦ���� YVU�h��e*���y}w^r�El|"
�tk�����sa���S���R��6|N�w�dCn�����T���!���u-�]��/o�xvY�i��p�����AC"�~K]��B�xE��0�ճ�����Ҫ��u8����ks2�
�"�ŀ�rq��R�F`�4Īp�E�Z����H��u�ȟo������i���t*��y�t֓���Z�CAFo��i���J�u�G�n���n�
Yln1W�uQ^Z/���d噘`l�f`��@R�������d�:��dW�}p>�Z�$����wu`�f⵻Q�����.��f)�x�^Ü��W7w{��frof��	Tk�[,���A��_feP9�N[����*!]���N��k�ٗ���-N(�I�}��\�p�۠��2l����D�e�Ÿ�I���LD�[ԁʫPL�]U��%5/Uf;�shgC�;w�_\��s2�_ V�i�Of� ��o��V-KT��9��C�Ba1��ptے�k�w��m!zu�y�2�z���Ã������&�u��3$@��9�k�'^���k<�����n޶��f5���G$;���r�WK�d{��iN�/Ec�K�ϦT�$n�`�r:x��wP�8�.��`Ko�N��钶K6��ow�n˒m�xyj�*|7���ٻ��s��Ӱl=����&e~�yq�_�Ճ:^d�!q��|�m�ÑBZQŞ���c���'�ɮO[�����7c*��Y����^��8h�}��5*�>fM�!�����D4�14Qb����2Ѹ��5�s*�̝]��&
�ݙקֺ=�MO��w���-�9�?DA������$)Rm���^�-8ȞX�DX�.�����G���g�#�5��fWCe6"��ӡ�Ϯ��s��(z�̧����ih��-�<�O>D�s���7��]���)E�Yh7k�˦ӛͮ�a�2����F������=8�=X�������z�k�Q�&�כ��B8s񲀰n��J��*����3�~Y���ۏ�؎",m����@�����o�\sV��|;{H%���E	��\R?z���z|���F֕��am��uD`�̤u߰,^�~�����������;!9�1M������uy��n����Ǫ�M��☷�I �յ{��N��������~PW_�m�����6E�	u���X2C�ܹ�G�Y��i�ǻT���]�s.�.�E�3sYCB<夳��U��lf����\Stn�86s���v�C�"=un�a�u��mٺ�ݱ�Gd���QѼ�9aZ�:��DWF�W��5�7l�+�ڂc~��z�K!U�$1f[���z�f0�
B�I�z�Fg����cl���%���qȥQɆ�o5���݉���AkL//&+�Ŀ]z���e�Ӆ3'"�w�+�V��v"��\UDo|�ц�����}�^��׼��˛יC�����QM��r �4,%��~���c%�>'�ǟ����ʫ^����t�E�Z"�dx��7�U����|��]3���C9|�k�w�R��g!��t��UH������xݎ��*�#�'32��^ў���NS�6��ۭ������3��b��AW,����V�W�2$�A��ʾ;�+}U�`��u�I��rx��I+�v�m��n�6   ��`��  F��ll    6�U��,��Hsc�3�+�'��9����=����T�n�W�T{8�0�>m���Mӑ�v{03��[u����R�v��M&�y���{lk�����/��<nn��C�7I�V�SfƑ4hKu9I�����.v���6v�0��]�ӷ'Iκ;���p.s8�s�lW6ԡ:�w<^��v��ʛf�5�׶B:�ڃ��ƴl6K!ƣm0�	I7�;�迮>�ț�N{�e�g���ԡ�n��Y���RW^Ęm����C�][eш�[n�gx�#�g*.'e\l�q3�T���}��ƌ�|S?�[Բ�� WؽiGP��5�i��`�TH�׃5�O�{�gX���3e�N<s���=HoV"�\Fq��L���c��;C��Gd����	���y�x�B����̋ɷ��E!u��C�1�*ǳD�̙��/��Z�e4�r(ZF<2�V������c��%�;��7���֜~٘U-����2������w7�}�������������Mv�6�[de�`��ϷC˽����g���d�9��m��Ւ�@��	q�#7'{6f2Ee�"��UK�J��c�����>�4kvb�55���%�M�1|ŋ������b��8*��t^k����F@�=O{��a}�s�w-H�S6�uͻ̵��� ��-#��<ǻ}�^����yUU�ٝI�
���F+���Y�7w{݇Y.2Ov��Sam��+�Gulw_CDl'	�\���V��vn����P5�a��<Fc�k��v��Ӛka�.���g��{2U��Z)�j�q$ƈ
�$7Z��gv��V�\r�L�8���F�5�Woç���-�{`k��V��ຯ:`'pi��0� ���t���`\N��F��O�Y��%��^6���f�'�J�nͪ贺ǭ;^���I徥�.�m���bAwu&k�;��k��M�x�,�mr�Nn�R�n�y����#�q�����"!�i��<9�Y��݋�S��[V�͜k��y�ybĆa���x��W�a�Z��㉆�R�c�_��;T�M܆Uv����xD���g��8ˣ�ߞ�Vm������*k�n���6�������%EU��P�h�~J�E��y�2�*�y�i�ͣ�Nf�
�ׇ�bz�����=<XG��؄s�F:A���Ba��a�h�c�y��F3G�1n�����ڧ�/�w°���iwr����)1 ��I3(WQ�_�JXE������K�_���"z���*���6��*i�3=єp��|2dI6�-��Q���9�PL*��������/H�oo=Wڎ����W1�؏-�M�l���Im鐩��������MR[D�ܶ٧XCjm�t����=�Sk:����v����y�InVx��L; d�gQ���u͛k6��3�s,X�l�X�^�f�f��4pn�P�K�gx�{�(G� ѫ�,��*�T��h��fE��-�1a͇�{�-``�4t�/S�t;#�����U��N6N?D�m��"�����*������a�U<�F�%�v�M�ָ���k����-5�ٲ�;����&��RFT-��.6�F���b܆�`n4/,&�|�1�;͖;��Y!0~û�gzV<���iy�D�����;��(#uǹ9*��B���R�����y�/f�l,d�^B��z0�&���,�������S�p�h �A|E!D"�Kz�����=����|
�B�#A�I��k���6Y���d��e	�~��R��fU��i�m�/��bmp�dY�v�%y#'&�B�-ڇkc��ڗ�m�ۥ6��:����5�b�Co��7
��/���3�'7�wVLwC\;N��C{t^��J38�UW�E�f�&�\��D�¤��3�wb+=�Q�o�_&`X�A �I^��2��������f���Z�'M��Z0'AE����{Ͻ���g���e�=����9çٵ��3s;�`FQ��x�=s6�>|��E#a�Q�,�x
�P�ˌ���7:��=]��[#��O����N"�`�N��1#y�݋�����fVR�i�4l�B�%WiDJ�K+��2��,0Wd,oe�uq�������t�e�m���mcֈ-�}�=���v�y+i�8!X��k����٥G��v���+2Ձڤg%5��n���9f뽲�n�{�$�����)�`  mp�P �;   F��T�( 7!��Y��᝞,=�6ӵY���k-���4n��f���s-����L�U=p�v��l.3Ƹ흋��\ʝ;��p���:��9��������[L�m��;��Q�t㱇�����#�\m����n��;n�#�5�Q�+W?���i�s��<�a�ԓ��m�������=#��F�wD�ǆ�n�m�]q֩5nm#t�x鐼<C�*�������N"�#U��[W;���n�֜n�H��A$umj�ڙ�{n3�+����+��N8��I���-]�q�z���aIOlW:V��v�:��)�Y��OJӵKD�@��_�{���Ƀ�#-���9(c����V���W^޽e���I��S˗J�{8�}$F�{�`�o!�(�8��7_���<0)8T`�#��zM�p�U��v�{慶���ߚ�U<]�oB�IF���|G�aW����«{��P0�07��Fd����g=\�����-X�S
�M;oSX�1CW5��=sN%qeJ���{m��ݧ�~�5�g��HĠ�)Y4
�'a�Nr՜�K��]<�lv�j��T�n�sru��](v�p��	��-��Q����j��7}�QG2V�>̦�iޘݷ�z0sC��cz{�h:ܻ���/7n#�1��w�L%1'S}�y>��.=^����v�q�;m���e����F�u��Q���фƁɉV}�2,�=��6v�x��dN�8��t�į) �N�nvÞt��J����:q�-�s���z�D������=�0�$���[�rh�P�l�v� �mY��~6�Rm�|�=�}��ѳ��c�/=���ob`��B�����xs�Zl�ȑ�|s�Wv8��猪̭n��%hU��v{���z� �jc��h21*s��4C��(�R�}�'��~���iI�گ6���4]���n�h�c[���x�l�ub5��졙	�kų9#��z���$-�
m���ǬΌS��ʷ>*t5��;p�3r�j�v��.[x�.�(ߟ��~��oU:������D�F	���x{�H��Ǜۃ���ۢ�`��r��{�WǡBi�1�c���zʵ���
�0��P��9�;L���x��̤���)
x����ҵ�Q�Dw1�?������,���*�̞�Nwap̜l�N��#�T[>���������m��gD޵��U�m����cM���]�M���Q��I��37�o�ٵ�/ߎ�r��s.D1a�.��9*ż�����UC�M�Ttw!b�V�U3��JMm�>U�C�?����]�"���褌���E!L�!Q�,��L�G]��}ҽ��W�z���S��z'p���1�J-qՈ��P�T����9�+5v�}��ޯ��\6�R�!'Jrһ��S���(��6��m�+,-��P6�ɸ�z�Z�B��m*�(�����U�����Ƀp7ob7��PONS�vm�a�|�t�����z��Ŷu4L*���z3�q���ӈ�
��w�d�Ⱥ]�hfS���A�R�7M�������&o^]�7;�h�gx"4��3*�y;��U>o�>��L����W��nU�m�������N��(�Zi��Y�D9���M�!N<';�>����>s���N�%4F�fO`���|E�\d��X�jy���,�C�t;)f݈�:���8v�T��A�j3�/�
h=͑�����>Tm��ls���3�#wfoWwĄ��q�ʎE�Yy�1�dȲv_��iW�y˿f<V��k<�S�~��+�FՄ�.�G;���ب�U��X�\U��b�H�퍷N��;��a�%���.��9��j�[!����߷<}��R�۹N�f[�y��˫��~ڑ���7�0R̤�V�1m��N�D�'��+�}�}�����W=�7m]j��$jѸ'l���b�0�d,�v#j�*:���f/V[�f+Y��6L�G��f[=3�^�]zڻ��+�v.�A��\j�����S���zϻ�S<�F�^L6"�m�?_Ta�bآ=8%�w�.�=�~nZw�Um�[�O2���nl~m@�QS8��]���=�6�a�"��$}�_v��i�G�p���\��m���s&Cn��%hL�}������yk(̋x�џ�.�ee�?�8�.Y�x�=���d�Fa6X �^@6މ3z����֚w���f/),,�f\�u��E�tX��7G��W;���y�:[����q��;�R%b�θ�3z���5"U��mp���A�5��ь��T8,nʄ)��n)���$oX;��ⲷ�_
�cK^����"h\zo�I���ehm�M��Z�[�S�!:t0^��N����-}�������M&S�g%��	��hL�%j����{\�7JW3��8�����IF�Yv��z��d���7	qf(��R�x���U�.�y}5j���
�8u!���;_K��*��p�����YY�[t%�X[S/O]���|��0M��}�ج�%�9]xY�����:�g皮X'!C>u�!HN����.0w,1��ȻA����`&�.��]v�Z�2%՜$�Lt�[���kM�`����+R6W�í�>�N��9ش��W.���+��鞐_wٻ�t n�e��J�Mp�4�j�QЧ�+q3j�J��/I�rGa"�L�Y���޺��n�ɔ7n���g.�;�.��א�i7�w�K#����~k�����       m��`H   k   h� �n���Zm��   6�    �`        :�  v��#`    H��m�  ���C�      6\%�P[j�q�b�j��   �`         �`    �� e�kJ�  ��    m �;��7X�����l��Vw=�a�.�q�ts��+���źn��ϱ��c\n6�w[ru\�IY�盦��/[�H�y.6-��M�zx���G/�����q��g�۾��̕{��p��ם��G6��wD,�nv�$�
��As�I�|[Wv��[8��^����1���زNٻ����[x雵۵��r�M�ŭ�=�޳�����O��k��{ˍ0������q���u�����-�aV�)��nɮ�l���c���')�Fy^oc�v�l��y����qdk��Vv�p\e�9-ƚ�z�v�����q����E�{v�[��'�A)�Q��e,-���(���չ;��@f��=���p�X}���q��Kn9�	�ʨ���&ml3yg�T���I�l�q��/"yR�.:�6��g���@v�Ñ6�Aqls�f4UP��\��ϵm���Y#
[S��[5�tӽۗo;O�ڷ\<��F���0�^�[��s��-h�qm�<<'V�p0�^�Ʈ�����aN���'mlmrܜ0�j��۷F��·;�cAƬ��a��^e7;��ew��/��(5q-�9�5�`6,a���<s@�������]�ڮ��mΝ1/1������o��.�6�	]�ی�xI.��M�cq۝�Snrd�����o'qɻ-��n8��#rn�ۆ�ʯa]s��}�.^��t-���|]�ͽi��K����6k�����b�î�z
|�{q�		�y�8�l�G$5�z�g�����{�jۓ�!������s���9�gy��m�YN�0 ��m�`  �� gY@ :�6    �h �iz2��N�e�o^:�9�k^���ޝ���'&7Eɝ�w�u��6�-cx]ٸ��Y.�X� $�tyS:�A��6�{\�/*$����H_}��$������m���-/�h��MBdzz�q�b��ƹS]`k�-�[^����n�ڮ"����V�Iɺ7iTx��&uf��e��I�bmq-%��s�9S�n=u��ۋ]�25ۉZr�����t�L�a�����?~Y��|���g񡘨��l
¶�MN"#y�6�.M���[Ɩ�cS�;���""=`���g�l��ki݈Z�)���(�#��)Md�3���ݤ����9�|�]A����|�c�"�:"h��3�B��+�<�{m��ڼm�Zii���X���QPZy�F���3���VB�|���l�XC�b\��Dx��6vɝa�z���H,eU Ğ��3&�* t^�R��@�h?�3�Ciԧ9�}}�>�~�;��ш��f$Qe����T�;ϙTs&�L�-�<ӳ����#A�t�fE��w��G-[F]�$S^7����?�ė{6�U���5m�N��F�m����-[�[���s����m�z��ъ�����w�91���3���<���zޗ����om�X�-V}�V�ڇ���=���+��#�k�Z1쑂[2����Vlҳљӡ����Q%�m�6d[SĻ��t��t{ye,Y�{�]���X�]�e>u�㊳eT��P�zߐ���U��T��oF9�Ɨ�=q���l�G�:f��e}�\�Ǜԛ&�I��UV�\�A�E\UyL�^��K��-v�Z|�9 I��}+U�Qf���΋�^�Y/���r�L>�y�ڔ6\u�2�5��d[Ԕ�\{�{�R����So?��<�􂙼5sQ�Ҷ{"��=�s�> �)Y ��U�	�')��]��b�7�m^�*�p��!n�G�[]s��T*z{��B���z�4���G~�������a�t@�)ZJ�TNÍ�u�v��q�uZ��[cw�'��n�C��#A�č(�A)#����긻Sq��-ai+x���VZl��N��2�t��:|F0��}�p��n�)�L���F�0�KQn?{��N_T6����R����󊧔� ���S��M�{�"e��[��<ƲV�P�
����Z��M����R|~I�s�W��fcIl��A)�j+�&�<�D-��X3��w��)n0>�r�m4���y�mx�������c%Ac�'�)v�wQؔc�.ϴo4���5���ݿ>���NOU�9���Ħ�!'*Hr�2��d50�:�y���[QW�M��w2d+o^��GE��w�ƈKe����=�a�%�l6�$�d)����=UlOFeM�4Al���mS����{|]���;Ԝ�b������g7�'w߿'�z��{���7�B� v��r9��.�K�jl;�k�tNō�a�1ȓ���r&\��ݱ߾]ctv���ez�y�d�Y�O����Le*p����[3>����*�n% PF��jP��[C�q��z��6l���vŧT��SN���9��V���]f���l�M��VM+�s�I�)�#r*�g2{�܂Spۻl��/9oZ�'`Н��{���0��6�":���i���vH���,�6Wt���E�t�}7�룟����}R:�����#��+�������i&�g$/2���˖�eJ^!I�5]�,f�m��KOgŗ��X���dK%��,�/7d4�Ta<� ��d�q��RA#$�0�'{�3��状M���[c��D�9�ޗ����
�@e�F�I�%n;�0�j���s���'sKZ��Ssy��*���y.ݏGAX��<��ۏ@���9Ւ��;ƝӦX�����ґ��BN�4o!0�'h�O�ۦ`�d�L3�8���YU���ョ����̫U�ƽm�cP���d�r-��D��?�vJ�Tʕ�����ؾvq�YKGEY���\�]�01�
�c�|�ﻰ}������L8
�U;{]�*G��=�=r�L��.����J���_U��'��S[Q�������z����o[P	qH�Mc-��w�3�x�G;2z�y�q��(U@̺[�͵W+�Ģy<�CN�X���ϟu���:$c�!�N��Q�A�����dK.������|�(�O}���L�����rZ���F�b"�s\ k�~���9ړNU�L�J�
H�w��ָp��a�Y��er���Wt�W���n[X;:�,!0�8D�����   m�Ұ!� n��   � �yۯ4�k�̽y�o:�<Gm��ۯ7�7X�[8�-�+�6��<up=� عû�)��i��\�;n�u�ڮa��f���\,jy�Okn:��`]-�#�9�������INZ�+��伎��e�^�+�&�e�7�'N�j�ؓڢݓtF��:=�J�G,�16�l$#���h��Ӝ��<�ݷ2�壴%ڎ��/;���7P�wܸfݛ��s_ ��ĺ��}����`Y�;=��[�y����^�3��zO�ۓNnW����u�lԼ�0�
4�QȽ�j�H�&��P�hQN�/',S�6GVq��K�Wm��Բ�Y���$c�%j����y�LX�0��M�C�Du%b�?������U��i�Dҋ����:��5F��ݸ|@��C��;���EՈ�|��˰-c��c�+
��7M�����(���Wiv]�!ڧF���
眉IU�/4k�V8��k��\�&w���	�&Y(�ʅ$g�&cˮ����Xέ��L��d���*�@��7���;tHI����mt�\]�:�~�|s���wYw��B���m�	�͹����@�x�sCx��q�Y�^Ƭ��-�r���Ø�����Lo�9thn��*�����V0:��2{�9��,Q��fγ�����컝���*K�S����˰x�^"�j�ҳ#k��W�"x�n�Z��g��Y}|2f#C���u>}J�x͉���V�6�Uշy-nc1|	�9�fT:��1ş��c����F4��iB +����;���eK'���~^u��%d-R	"JU�}��wv�7�9S.���މ�ɢ��q��U�"�b�`o[�v��ƴ��W��Ӆm���H��6dnE�̼ϟr����Y�(+�USGg�2"��ob6�:�#,>���k���S�o=�#6�R�n�AU�J����>�^�K���h~��'w��b�Φg�ي�3gy�d�H�Q�w���gbR�a!���n�*��F{!�����펱�ˮm95^yo�*�n���n;�{��Tn������2����f
�����\�������^1\a��~ԓIIE�I3!�}�~CٌMӷsKGC���s^!�3o���@�t�k\�L̝1�u���ۯ7<�BH�W�Ry��N6�7
R2�j�����WtV!��g�:��K1��������cj���d�k�����e�V�F�{���
�)T��=pݭ3o�WJ���+!T7��FL�e�mޱ�=��MU]���̄V8�	�!���h�L;��V��u���j=�j�+%T����>jR�s#���3#nR0����G�}=$,��9�Jnki���;@!��Jв�FgeM���՝]�3ٟ�K��<c=KZʁ�\��S۷��1�j! �m�O��������٤r	%d�(�RA;��KFS3��;ͱb⌾Y��=�\tl��|n��M�g	���q�������m`�E�d�:2��)M��"q�^�$�O7�|>Lo�����U뺯���GF&�
8KR+��yW�w'G�m���~��Om�E@�d�g���F�n�@5R���"qi���(>�h~mB�D�(�{FR�+���ϙ>l1��w
AZ�5�;�=�v�Y-g�k��{j��A��{/o^�cd@�)�mɘ����̰��wW:7z36����zư#"��M�4իQ��h d�?=YP�-���EVǓ;�a�V�g,W���h����6�:E���Վ,�S��[�Y�����z]vyLt/0'z�8v���.�@J�b黗�}m�Ts��x��
�־�{]p�%,��wɕ��s1LQN�l����@L؛i�$I���kHN&H��k�I�iwY�������B/g���^:ْ]�ssL��W~���ߣ��v����M���5>��H9�d�hq��U8Zl�4Y0���rg��SfU���9�&v��C��x�w�cqu�W	~�q��ȇ���˴6�q�<�w;��A�fc�6�����Gj^����͜���>�&L4Dˈ���Ӗ�_'�kF�tET�2��ʩ�K]�6�e^���FVLn���\�����\�n�# �����m��<qo+a~��G��u��&��j�ʉ�0U{ͷ����5Πb�����,�R��Z7�w��IpE�Ŗ-���!$�d�H���꣗^����mg3�'b��=�C��t?e<@��A=�6?���[!rTR����%	�16(�@��MW$2	d�-��4�jg��E�H;��E�;D�2�y6]��N+�|��O��~|���!m�$P��m� i 	-�      $  $���]-ѳW1a��m��h+f�^��-����v�R1:�!�9����9�MsH���r�w&��ntm8�yW���lk�97j'y����N����w]��G�8�5 X��� ݋�;�q�M�~d�>;�N��tavUI��t��+ld�k��$�n���E�M�m�����l���ںXrd����	��-�[���rJ��������A"�/��/��,�����{)��x�	>��A����ql^� ^2=ټ ��W!a\�p�[���ɡ$B�/�$���v;(���R/u�%U�[!�	�N������{���i�[
71��W>�6����e�9vk5&�M��.y�=��4��4�}F�U�`R�*CMt�$��J+�LC��c�2w�\{Hk{�A!��N;��v�)R���e�e!$fMX�S6�`$���Y�#L��O����b{�0bwM(��gu.�7����������P^�?�
HX4��]�Ueu�u���D�#�7��:�Ӡ;�ї��[^�w�j=8�$L�@I�[��v�"U �)��F���	;P����#�]�m�i�B��Ѭu��n��]��Z����ɭK��?�ǭv�ĝ��U�7آj���}KJ��Wp��_Q�)+�y��I�n"N�s�C�x[����v�����XA3�����|o���ٜ������vikp���xDd�P�Y�fU�}F�Y�9���@1�e��I��WG��|�<��C`*!.�gq5"��8�z��D�N�JqK4����]����{x���}�zf�[���u<�&��q�jHbqW�f	D}��Y<芨�稄��繽o�����y����^"Ʃ���E�il�^��k	��1�$c)#���{�cژ���)���x�v�O���|�{9I�/˽�*>��IS�]�FT�eX�[:Ua���=�L��\1g��I�Sc�wv"��
�/�o3�����oWr�q���<˺��wg�&�t��%�+�廿�$� �m�Um�L꣸Bq��`h)��ՠ�w/#n#f�5�N����/ne׮�u����
�����`#'�����)K��XH�i�D[��y葷mf����ͥ�ˆ�?%��8Oqs���	�SA�	��f@�9̇��3�ֲ��f���C	1 Qyǎqv�8���ƴ��V�.�#��zT:�s�>�s�����{Қa�d1����,ݭ�z��)T�A����{�M��mI�43s>䴷�TU21X���:��o��C�j������w�!:���#w�X�mCF������Ve=��*��=�e����yn���W>��UG��u#5���uF^5�HpV�;�3�V�֕[}���)xi��vEmwf����&�@�ϬeK���d�#�ݨ�83�9�֗��4:��,��d_P�s����]Gw��Z��Y�kdw)�޶�iX���͊]gV��iV���#������W��u�ȹ��KT� +A���h�<��{�v�P�W'-e�:�u�\\ޑa,U�C8��0P��S/���_opi���Bf^��YY��_�έ�D��r�٭}Z��H�GpP�q:8�y��$�t����u���G��x��Fƻ��^=��5��k�a$��+���|��b�nj�ٜ���ԾΛ-�.︜��Q%�#&;��\9,��ݏ6_1��'��T �+�����Ȓ!��{��ܯ�t����ݘ�^���h��'L^��g��e�f<�؇p��}d��V�̹�j�Qsf����LY���y�8���.�^�|�"0n�� sT��>O��U�Z�,U�y�"��͠�z�H�H7���2(��{���?׹r��^����^��.��=�X+�3n&�lR*$��O6�j���LK��/���g��;�����w��Q�ݞBi*Q-�~�)�}�o����A֝���4[%�(�rx��D���1�o"k{�tW<N�}ݧ[�^�ɭ+��+1w���Rk)�2��S�ku�dx�xx��\R���J:��Քݮ�ג��� t��۪惷Y�:�����m���Z�_��58�N;�����;u���d�eD;{�c�%�%�B1��)�7�$�Fc�d!�H�:�A6�l���{���UU�2�Y��È��ӯ���2	H}�}C2H
��`z��ų����]U���n1LT�=���l�&���QD�/�D㡘�Xae�{�珰{<Xb� ��+�o�5�k;#1�Q�,����G[�X7�.�u��gp��E�8�fO+�{�#�������S,���Ϲ4�*����L�W1��!>tU�Ǚ(�^�ϸ�E��Y�_.NY�i�7oI�y�GR�)��M��k1v���e\��HumfТhb2�Q�&��y��ϳs��߫�'����4������`R S�2˂���/z,�����z���A���]��jF�jm<O�S��g�㒛,d8`�U8���j�Ea�Щb����,ҿ�	�$��"��n͡��n<��Wn;pw]�#��\���G�(�3b�mvsv�+�ݒӤ�;������ަ�����E�#+e��׈�@�o#U@a�f�hJ��1�oU�g�O��x\� ص~�,̬BG�|�B�T
)��*��0�a�±%� fz;w��ù��	���#Ʃ�f8�`�G!�����.=q����G[� �c B������_C���i��z]��x;̵��ΐ{#��뫮&��;nd�<�+��2�7��89�/=;�>3[�-@�i¤���EfEʄ�����Fmd{)���b.*�lX�=s��O��N�!�zO��/=��>�s�+�b�<�SDi��nBd(����A�.uP0����(}��f{<R��׭�ݵ5�n"gy�A��1���<�|�(�{(?3k6�]�����gz+���+�Τ��>J�^�Y�����We�h��]w�5���k�ԒI$�X�@�`   6�@�-  -�y[   ��� 3�;	�k��p�6�,\�gYf�l�j�\�kY����u۲�/h�\�a֑*k�g��F��]���7[d3anϛ��BK="��^�nV��n�K�$��i��a�^�����3��n�Vy��4]8���[d��tL[O[F�=���c0TWw iӓoYp���L�.۫f
��c������n�X�x��:��:���d�Gظݜ�gccu�&g^����������}�#Xl�EWuK3��}�;�`Y�7�F��M_8�فЙ���ן~���|�kt/}M$X�&�`�Ўy�F����<���&���(�h�zD�	�T�
5���ui&2�������90i��C��nr?���x4w�S`�d�D�FAC�&Ͼ��Y3ߌ�'i}pУ�fm���g߸���TK����i�><��ɍ�����.�#��s���5����
��ۃ�{��UL�:)���n��j5�1X1��!����	��F���D�g^y��$P����F�nD�M3$H��C�ݧ��0V�2�Z�V�ۮ�5�Dj�|�U�?��z�C��h�
�6���[* s����"�����]Z�g��|�A��a!<�I��Km�������Mn-�)�ɵ��\n�^w~?Z'�����vx��h�U۽7�|m	���(��s��%o �����k��"��w��󥦱io��ݳ��݌�"�V
G�vO��|��U����߾�<�L�����m�δñ��c޿{����N]#u��jj��"�.�*i�ay�v�-�M�R�z>�"ߖ���8�C�]�q��j�`j��S��H��{�����ȫ� �ҟ���f_:y*�3���O���iJ�@�~�%ca����O��j���z3���5C��6�ZE!"$)�|̭0y�t��>*`����{����xU^���B{[�l�,]�sϪ�X�%xH��o�Z���k��ԙbF�,Iē.|{��M!�v��R����l�ET:w�`�.� V��h�����=(��� �����x����6�Pb��V׫��(\r�Ӓ&��=���M��-�mv�q`�c]��у��/WI3���.K���<�﬉�~�NL����O���@�E���D�(������m�G��n��Y����&sbj��C��lf(���яIqBYb$���	[�s�8����E�JM�R��@<m���ZVc\?� �h�V$��2}��M���s;+�U�����N�{�O��N�y��
q����O2��=m�oک|��LLH,��ZD�oo7��xK���]�t�|��*����m��{3G�p_!}�Fk��.�r^�^L�2^�{{`�S~�~�@�����=�j�.ClWDǱ�=8��"��~i3���5#���w��:��瞙n��1���sy�����^�Uy�����ۖ���MaX<�?�������no�7��H�������lt8�8cNI$Vn��KQ�=�</�t�ł#ȉ)�"�c�a+y��x��E��0�����~GW2��,���M�XC�
8D�������~WX�!:���M�$#� �6��4��j3��ݨ���늛iӓK��%���E:]��(�>K��Q/��@d�)���5\Wַ���Y���b+�Uq�Iu�������F���|���M�L S�b���A�A�[�v�H`�O���g����fT��ǎq��d&��9.N��;�n(��t|y���>��]nC�mA���q�<q���m��bH�e���{>�B���E�	ꏻ�����o`$����.ܨ�޲���/�X@�����i�G�S���!�����x,��i�jY2�D�����>w�z�pv$�uP��>i&+4H���t�6O.9�=�;~��Fu
;��7\����V-�7f	�ਈ�}�:�JE�����l-��
�g��a�w:}3>�r���5��Ie,0=<s�1�l0p(�M�,x���@NI��y-�N2��j��:��k֚�Im"�As�M�h"=604Gm�i�#<o}'��0�C�&�jR��k:wgMɭݪ�y��on)�7�E�C:܍������M��ڱI��bqg�׳֩Jq�e�7�c�����ݽ�/��e�gL�N$�k5p�N޻������N.�����[0��D3�F��yJl��d4P�m�IA��7ح5
	�>@��t���u��t�C=�{��	�O|���2'�� 鿓ȒrAQ��m��,��"��ˈ�g����<<����v<�� c��GRS5=�g��z]���,�1�\��`���8�篤/��D�q�ɑ��#��@[Q�����T�O#g��-��\�Np�����:�DO>#�������`��:��7��}��*n��/K|���D(�ު@��$%4D8�s��*<h�R6{w����!r��W�����+qtNv��$�Cǎ����] X��E���dsu�k1(�ƅ�O}^2��m5�f��yY�]X�֞q�!w3��3!��6n�Nv��e<�:}��z��}k�I$�T��m�:6�   ;m���( o   ��  lM*�&��yU��qɺ�ִ��P9���zݽ��1WG����;�cyb6]��:���َzOb�.Kָ��][��́�d��r����Â9Z���$uk4����N��pu�iD��ޭ�l=�+� �M�=s�[�n�1���[�9'4�yXӦ�m���\[er<����NDZ�����9+��ͬƻ�u��l�!8�lHc%�8RfO��}k�5�����_���\�s�>�\�	>��Mr��|��; \c�u�7�Z�מu@��;��qc�tv��$�Q���7 x�O��h-�E n8���L�ࡄXTx1���5p�f�hֽ�`J��iY�y���΀�����YH��ǭW�/��G���p"�y�	3<�V7�#po�>���d�*Ho�wc��Bpld��+��W�<\$�(�y����g:�Wl^�o޲ʙq]��B�}9f���d��� ۺ�z�0�|�È[d��H�������|׊ɥ(�',��i�}�g�8��s���m��@S3�v'�}Nn��!gݭ�D��(�0�H�*(g��e=Qq�R4ܞ�<x0�쁐yg���7����B�D�BΟ��Pt�p��T�y�|���%ϵМ�-�ΔO���N��8;I�:�� �W����S����:��YwӶ�%�H)���ۑ:���u�:Κ��ץ<�(�j��';5uݚq6A���N�<�;����r�|�4���8�#Ȟ
��>e^��g���O�z�89ҫϷ�@���@�4������X+���8�"��`�R�`�۫��H�LA�&�U����ix���&���&���;��y�k���t�H;c�C�iJh�K��kҷ�	�#ѣM�:�-4�z"��:X��O���K��.FN�o;�i'�߾W�y�tB8Gg��]r��.qt�dg��5�x��V�/�e܋���z�^!�P��m�\ Q�u�G���>��}|�aC����|���;��(K�Y��gW]�TO��y�B��z�X��� kD_ϕ�޺Bd`�E�w��� �����E2\���)����p��y{Nn8kL���H?k�����da� �����C��� |G �|yu��d�7V��@\A��at�G�4TK3z�u�|��>/��|��D����0�%�J2
�_	$��cC�zƱ�j�ψ�Ǜ�mi��|�W�5m}Yn����c�y8> u���߳O}c��#�O�`|x�Q+�#�vw]	Ä�Ξ 5T�9㏊��У�B�-B�rC�Ճ����`�df��nP�t�m]��*{k\�<ksqh8�)��I���`�őg�x����u�� H= 
,���ްHL=g�y�ӱ c�ؑ���-}�KP��]���#��wR�@��'�\"@�������䀧A���C��9�� �8�߆���TO�:vh�s���,�!����u�X�������4вx|x<X�ǌ��mGSȏ l�T
�,z=&�ܿv0�4�#Օ����2i�����V �O>!���yMn��\�����#ǖX��{�J�,�|��6��IƵvo_P��#I(ωl>x��R鏹�\�^4��>3T�ϕ:<n�/Mꖫ��jŵt��y"}��quq��·!��|DΞ¢��nzǼ8�D� E��R6x�OJ�{�$��m�܎��
 �Y��#�o�:Ǒ��#���5��^ #��DO7�m�PD@Q�d�G0�m �����t���t���L60�4�m���߄�0��� �x��I�@�px����"e��F8�qt"���sψ��f�
7���@�YupR���,�~��En��� ��*����ֺA@��� 0�� �[i�q�6}�q�8<C�"��e��cv�Q'm�ggVٮ���&۟(Nnޒ0����9��i`���Æ�\�њut��r���G��g���<C���}|�WH�|^ Y��7�\
P8!��\� o��C���]=w-Q�Ux����	 �y�;��� �:x�&��O���qp�"�R��l�g
m����x�����.p�k�:a�<�
��2���@}]���=Ђ $��ψ�vA;8.In�:y���<�D�۾�><ጱ�w���. ��� ^�L�"Q(K�YpP��!� x8(�ow]p{�d�|@����@c���n�����r�����0x4�s��2�����>0���L����n����.@��r� ��߾Й� d��)H	RC����y�p!Ϗ9Ϙ(U�`�� ������m����y�� Hp�yP����������Ǹ͉Z�|� � 2�r���i��M݌(:e�0+��+S�k��\�̺�*������.W[��zLe�q��%j�B��y���rH���~�[d�'�8�p7�� z��O81 ����8$=ޜ��a$pY S@�� ��}����M⺫z�9��pv��O8�9��Y��� X#ǀx�G<@F�9Ϯm��s @�yHs�y�@t�p�:�ǥiO�6�2&[�NsJm����!ַu�^�̸A�-��v��l�OiIf΍��Hk���w|�w{�g���8>k�x�h-�x+��C�� ������9��� <�W>�\�r]uD����>#��<D.Tye�fG�6�G�|��D��I@��!�#2(�q���y�<�:��4��8ΐ"��@sǓ�q=�}�2�i::�8���/�-�,���y�8*�Ĺ��᯶�|��9d<�� D
 �k��0�<�=���W �ǃ�G9���~�S06�h��x�	���8(�U��C� ",�v���p�83v���<x8(��O_æRъs�G8>��!�
Y:�s���<����9��w�hp<�G@ H�uP�&D���M�\ t��w�`?]�G���� ��#޳���| � x9��]0�9��y��n��80�axO9� p�>L$��;8 .�۠�� r� � (�� ���ڨ�h�K���	C2� ���G�sG8(�r�s������ �� e�f�:�x4uY��Y�8�:G<y�Y�>�ԧO7��̮��s�����Ĥ��$�R@i) <�H
��) <�H��JH���� 1���$uI�R@wT�$�I�R@p� ?�(+$�k?�4�`�G0
 ?��d��A���UJ�DT��R��RT}����
�T�钨R�R�
JP�EJAP�4QBJP)Jhl�$�                     P              �         o�����_^=r��7�m]���R�v����g����w��]��W��徤7ۯ��y�{�{�w�w��V���  �����ݾ78ھ��x۾��E U��ow�w{�}����������Ϡ 󾭴���_V�:}�������[�wM����|��_}�����w>������=l6�<mJ������{��s����ӡW� }       �yn�������u�����/U�i^}�z�w���|�����yޟ  �w���|��}�}�s��՟]Ӿ�g}}���۾6�)m�< ݯv���o�{ݵw�{�m�N���6�X�xޝzZg<y�+˙� �Ǖ^�o>����R�>u�[g��|_{z�So����>���� �{my�;ϭv�{�7}��w{�|��}�%������1�%
ͻ�         C���w��e}w�{��ҷ����_��ϯ{�w^�� �_v���毽�k����o��o��ޟO5���W�ϭ�s� �W�o���ϕ�m�E�>��}6d� ,�5Ux��4S�)�)Ep 瑬�h��׬�W�(��=�::4yt��(���ۀ f�=18���v2G��W�U{e�nQ��]�;�&�+�������         �ϒ�H�e�*����*�b��tyh�=4D�{� oI��w�o6���tU�i#��)9�q�W�RK�� \�e*��5�{�kŪ)x�� ���Nx����c�9ݲ�$� �F���t������Dy�:�Q�c���i�J{� ����Z��ze*�w��cOF����v�Dy���6�B�kf5��   }     �tQlEs���tuZ/9��:k�ttTy�/=�.�D�7� �{kX�';��I�[.RM2.6�kl���x�U�`��� {��8���J���$%� �(H��<��aE4�ӷ��W�Ӛ�� .���vv�x��
��O�5U8ڻ^�wW;���J�� �*�h
ܰyzt4��d^���΀�4���/�5��  ����@ �{FR�i�42�oL�5US@22 ��U*'�U6� 0��~� R�@jxATI� 1O���/���n�e<���tP3�8!�v����ֿ�s� s��8�����p�s���9���9�9�s���s�s��?��8 �9�p󃃃���8?g��ߗ�.��<3�35
H��m	����c�#��6��U���i��3z�
��h��ɍ�W	o>�-W׸-�Ld�L7z6Y��V�^��B
U��F�̳H�/yX197f�אd1ba-{�J�k:�\�٪�Jm!�Mn��yB�ɷB�l;�Z��tq}n�ݧv�	m3$�ݔ�H)�H�r5)Q�ʐ�&Y���-�;JT���o)�c�4����KJ�on���w����\��۽+\M7Cb�ub񄉉��^޽sf�n�[���p�'Joaw�Fb+%�`�*�*0w&����bÚ������]�����C��# -���/�-1�Mbm�w�ˋKAU���
'A���젪��dx[���²bF��Ԟ��Po`kVf&���IV[�l�V���J�;����&o9e��*��ݛڊ]�z�;���h]�2H���J���6vv��33)gj��BiH�(h*ݼn��Q��1�a�r��8T�YSjbh����Z�`��0���60��dt�9�
�Uz1��lٚ͢�A,3�Fb�l3b�J]�cj8�b�F�wǛ�9�e(��� "�'5Հ�*�Y�N�p�FK/4�j�yn�c-p��^LJnnŧ�E��Mŀ�XsN�mCqF�B�*
�g��E��)�rө�`*r��,nSRa�7,b�{Cj�KXx�\Ǵ�G �U��Z2ɂ���(�٘&^dz-^53�-��,�0J�jn�r�Zd@M��l�|ݖ͒��9#8��E����*¬��� ޅ���m�(��Om�ˉ]EY���kr6���2��]�N�U�fz�e�:�&����dM������i�� �9�G����82a�l0�j�<k9�����GY�e�@�J�2C0o̜�4��abJ8���5�ؖ֌t#�z�]U]Xi]_;��n�;Xy抚A��JXF�6��Cv-f�VT4�6J�A`�,�y`c�^Q�[m��F�G05�E���P:�:���!�ļr{��7N��f�{nr���m���e��1YrV)�&�(Ә4Gg0CM�naV�^B�am���D�v@�:�r�H/��÷��w��d����hU"Q���x��YD�:)G��G/,Yy
�-h"�b�|����2�EGJBj���ySpHW�/bz�#s3]��^�T����i薃��2
7.��rQ��5ӫŬX�k^�֔�Y������'*�����%[��G3>6R����ѷ��ʸ>��M<�������q��ӛV�EaV*��ɚS�R5��nŸ́��É�\���GjE([á�`�IV*��KVu��]��^9�RFՅ�naP�@c"e�!�utY��w-���Y&r��� 鴋B�*ջ�Vo&�8��Ȳe�4h������<���QU}O�9b����{4�p`�mԯὮ�L}[pjk]_��U�L��0�R.RZfʨ��JL�v`���	�3�J�X�b�2�Tk�I��eރS;��)3x/n%��Eތ�I(o3Fk�%�R�Qk$"�VE��ڳa�I�!��'s#9��.�w6�z�V��-��X.5Gn���h� �5nì�yX�c7�
A�4�
�2�Ң����W04�`}l����bG������i�kڙ�ҝ�glֻ�Mp8p�.M �ԙ�
�m�Ol���t4�W���争n]*66T�eµ*�5!D[��h�Y[EǛ�{�]dd-9�s�j�Il�ZȢIPe4P�J�3YW���Јˊ� �c�]�c���i�H��"�6ؽ����3��/މ0����w���T���KV�La�4	ӀY�=�˥�٪TH��Q�6n]��vD�-R�mf2Ň�^-X��s!UU7L�2�U�-����;�7sC��օ�h+tL�2�L�+JE�e�{6����j҆�r�B�( ͭ���Ժ�5�7"/Tr�:��U���
W�a�u���R]JtN�Km�ݺ� �݉���I5�S��Zr*ZP˲�$i$�$��	5���[�f��? ��.�o`;r7.��dې٨ֶ��H1�sj��r�8w+5�$�-^e�$�X0n0�\6��C6x;�k�� [l5��q��c:�|��� �@�.ZN���Sr��ӻӗ��WcT�������Y`����R��,�<�v�1�F���� �%�fc��f�f�E��T�[�`Ґ�wf��w����A+[9qD�e�+�����p�I��4�Ef���n�eۍPy���l�o��U���uz��DwF��yS*J���Wl�f<w�R׎�:$9��8
,�I�[L��ƫwWl�:��n&C��H����>�e���aY���xsS(�&��V4ъ��+�b  �h{i��ɉ1w&=��Y��Zt�����Ք�c7��73eܛB�^0"0�43�b6v�-M�$f�R�&�^ܹ�i��F���F�b�d���ÁT�l l|�����v�ֽ�,z�ʒ��E�u*���!��qYOl���m�S켺�J�9fjc^�V��X;A�t��v&3m9���r�jkiAr�q �����N,���hX�&�	�`$�-�=Wv+T�
�uMUn�t�w�.����ؚ��a{��i��v.���1���EcAͼ�Ph����[�[�\��p�_�+� �w0�6�퓻$�Z��p����W�T��u{�XmAx�4��fn]$�sMi͹ջ���#�%M��	�dr��͝:UL�=h��r�Ͳ�Ǡ̰pX�BLiP�S;d��g����}�z:��s�ᨛ��A����t�L��p�V��en�$-���e�NHQ�4��%ǻ�I7&�NV�9Z�L��PA��f��.0u�nK�$*��3{%�����On�(ӳG�b�$��e͙o@�:��u��Ř&,�U�ۣ�{���u0^� 飵+��F�V��ӗi�����x�ٶ�*�^�EI���Y��2�\��(ͮd��S"K�IcOC�{���[�Eo���R0�"T�R[��/w��3&r�D%᩺o%�Ee �\��$i摵�����gB��hd��+1;��"R=��G'tJr��6ekOD�xN��ݭF`�`q�K�KvV_W��Rr����=�c��کB��t29z�p&�&���5s�g>�E��F�d͒�fQ�����d0�
��^��-4mꪥ���K*	�U���įg!���EU紑���q�jB'P��"����UQͮ�n7g�yT��VT�Ui:A�!l�^]�UT��f���C.SR��)����K!�ޣڼv�,W�y��mm[oy��!�Z.��j8o$Y�i�/i��U�oMek����Y '�-Su�l7r�^��}����䩐 3O]�^�7��"{;btLΑ%
Y�n,3X2��V&�)cSa;��]Ma�����P�s���F�/�a.�<���v������&�Y�f�;nŊU�pǖa0c[g���{Nm���N&�Ø�Y|��>d-�$��v��w�V�ge��$V7E��&�Xd��Q4d;z�	v[�[k�7�=�ji(�n�e��gL���K��hE���V�]Q ����+	��ư�U4�r�]�9���l��{�6�8�h"-e�mjU��h��n=P\:p�����P��A���e�ݡuj�Zg�)��k6��+�������MýG5�i9�M�dj�snN��U}oO1�nv�廐^QX(�жI���\؁g-�%QI�����}��=�y��R���Q#RTP�0
�f&��TGq��n�o7�5�r��>�=��W��c���q<��z����F��h-�J�Zh������x��4�A��m���<2�դ̩5��0R��Ir��)�)�Zn�C���nݫH!�v̓6�T���rfm[z�(&EbA�aM��rR�%AN
w�,¢��r�� ��5t��'6��>7yoi���u]��4(:��6�ڻ�W�Lf^��S�,����Tf����U%T�s�b��˧�K�*6�o���t�f�P��,,5މ��́b��QH���+k9�2�X�I0��˚�YdJ�T���fI�������q=s!"�`�KI3V��}�Wi�È�/S�j;�C.C��ȝܘ(�U��;��4Vf�!q�SrMR+UOk�U�
��^i8�t��</k&�^�̴\v.X/rQ�x#r���.`7��]ؗJ�A�� ��F�������a\�$�H[�oFÙ��2p��x2ŽT��_��{XӘ�!���V�Ĳ-]ۛ�+ Œ�Xb�jĘ��-�Yt�]�$��U%�=_���(`��Dͭ�v[{hn=G�pkW� �fT��p�p<�qY��*a�p
�̳B]Ų�y;X���L1q�J����]3�;U������GY�V�;�M�J�H�P�7�u)ed6n�!u����X >Ԝ[������[Y�m����w-���S	عR���օa���5.Q�2���ɹ�rg$/��/&���9�e�t�f�ѪPDY�^��-�C��3
\۸�}jֶ��wJ��gMʂ��a��2�6�� w���z��ǆ����d��j&K�/:���{���7��wf��a!b��;t_'q�;О	#����Wv{��n���f�+�;G\2�����Ӷȑ�ɷCSvrCN�٢�J���QA'b�g�Cޜ��ޘ�&��5��	e�۳����,)�=��+2�C.�d=�]0:Ǡ�,4G]���f�ݙyF�#yk-u�a�Ƕ� ��W\p��LT\ff
�0c7�V�H�8q�����z즞�\�;�n;I���*Ol�B�=���ܸQG)�P'�F
k��
K	3-�f+�]��)�E�5�$�R�䗕f`���R���E��]Q�[E� �ΩzyD�$��f��ɻ2�>tcn�LMP�cV���l�E��0-Z���k%d�N�1��vm�L��U�й�Z_,<������{d���[HY�8w�����-�lC���d3��N��w����c�{�Ltt�z� e�j;]��R�᫹��]�l��N�s!͐��a�#����dlj�T!�b�Okٱ��Mv�;��h&2�\�$���S�V.H�D��á�Ud���/`5�[s^e�P;	M�qP�NV��{��d[�)t�`��f۸�P��ٹds&f��f���ќo��W����֤ ֋"�f��F ��d�b�R�k>���@B��&�ʗ2�'[r
�Y���,/G�k22g��J�/"����\+M�*�3EB"��˽p3/�E�˖�=�8�F9,�1�[dV���
�u��37��ky�BƃM�	jʼ���I�&����Q��6!Q�Ac{n�[N�a�rT<l)�5Jע��0:�:�'�O�Me�v:n�۽(�`/hM�ֲB�
�5�X.��Q���[:�$�Պf�a� 2�:�H�.M˱d�S
n�k�z����A�:��4Ԩi���r�(���e[n*eK�r��q�Y�Nn��,�۷uz�j�[X�]�+Ӫ���ԗ����moke���iۏV�;�{w�wd��sAu���+uA	k0�&�`�HK��V�ˏR�r�ҵ�`�7�Yq��]����C�P,�/�&��v�f��0$�㰖�v��%`ڱL�%0�Yr�����I�㚳fH�N����ۡ�ȱAͪ	I�')	�^m���3eJ	䙔K2�R*Ҧj"�)^ufLAb$�P��뢍���p`�V��q}�-��x�(���G�ڇ�����{oV���-rRs�6���]e�!م��P�M9v�@=�
�ݭ8uD+)�L��׎�[-�dlL���.�͊y�4��e%��Ra�.�v�%���M	��d̨��kq)Knk�� L�ݐ��R�rED�,V�e�.lx�����[ղ����T�R[�ǂ�jԪTÒ���a��a�;V��Kh�[Y�ZB�m7h;���v�#�]ht�J�J�~V�7R��u	sU��,h[�#�rj[,Z��m����˄	&�����\\�ffⰂ��z��ƷNG�0e�:�".��m��ڷ��p���з6쵢9�*^��e,:Tu��h���)K���J8�YH�t�b�wsp,͗4���OnQ�����Unj�٬-r��dĎ�z��:�k����&[���E��o�PΊ�ݎvcjvs�R̮ 8N�VZ뛪�tX�P\�L(�-f�+����]�r� ��3��7r��ib$֙x�^��W�;��9�%f[�[���Y���Kr��'��h��X��ZpMHŗ�ـ������WdQ��D*(e!D�[�Xs���t�����w���C�y�S`��Q�Q�l<qw�����](��XK�'�g2<��t[�B,��2�7؞�Z+���cm2�6+[%VU0�yh]ԁ(�ס��Stڡ�cu��0�����Ջ���O�����U�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUJ�UUmUUUUUUV�UUUU�rUUmU@UUUUAN�5UUW]n�]U�UJ�VҭuVƦ���Z�U��������������������������*����UUUlڪ��j����������_R�UT���U�UUӠ
�������ZU���&��U���p�É�� `�z����z�n	���
�V]����d����Z��}UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUWUUUUUUUR�]UUuT�=S2�;��G��u��v2�ͭ�/v��;v�9�sQ�e��qs�8g��ysmP��Gr���zu�m��n����q�G��v�\���=����<����6�A�e�[C�	kOf�Cˠv��i.��\r���n�X۲���`{V������km[0�9m��+�����<�)��͎pc�r�qs�s�l9�xM�ڻv��Oy�8=�K���=mی�j!��힕M7��v1VQ7IH���ώj�lV-�s�n���cTO
ܪ�Ø����Y��|]��6��t�[�<lG��tz.D^���:�m����a�=�'Nv1I�m��l�=l�֝�mlx���q���:w��z���yw-ñ�7�5�Z;n0��9��[iß;�$[��:���<��nk���ۖ�F��s��8��lPq�f�ہ;<�ˣ��fcq=��n���r�M�s⭻3���t\i�p�/)�N��]nw�u��{m���v���lfEȝuF� ��鬍bre���c��˧"繹6��X��p-f&x��Nv�is��puu���ۦ;�p�}����v��c�������9��i����ȝ��ܘ��s=��;���s�c����L>�we����nv�5m�.����ػF�u�h��u���q�v��8�a�����<�/Wp1���;�r�G7�)�n�;���N��㝕�m�p���l�ړ=n���n�t�5�tv��ˏ'U:Ҽ�:������9gv��ۅ��t�P�^�2JG�qw���`g��BrH�(�E�Vݣe';
����������%������!;�tx�u�DD���w �v_�����ø�9wf[�,pu���)�k�lC]Q�.�m�L�&�ёs]�q �:��1��������z{.d{l!��7.{8�3خ�kǁ����s��������f��%��G�>mݮ�vs�nM�݅�n�]��c��p'��s������m��qp��λvEnD���N$CXE!c�X�t��t۪�Xx��sn}v�s��5T��=v�8^6oF�p�y-�����]��h�h�u�u����y��.{i�v��.^�W����Ja��h����ӅKG)&�y�X'b*�z	{[m�v�,��ظ���A��zs�:�n���JU�g���Au��@�n���sF�˝;7g���Ǌ�\O���s����]	�]M��cW.�m��"�ڸv�'�)��m���;t0vɍ�Ps�7,�br�*U�²x��r�pwu�ۛ*y�ط��;rfB�೚ͨ8 �2kp�m�-���ם�6N����\�M�Kbp���p��g�\��.�^;h���pd���z��J����n��	��s=�6dn�]��u����$v���r�J��j��j���a0�k`㗶x�q�j�'ׇ�ݑyN>��\�d�Cu�ת��qv�]x�p�jn����w\\�����1^�9�Y�¦�x��ܰ���۲�q:{7g[��0cm��0v����7k��_.�k�H�'E��t�v��#OA��=z��*��y�{u��wI�9�)=�nAb,[n޳��8��]�h�jݹ�(.�#��=�h$���Í�K�۝ή��Ő�]m�xu�-�h5�䱍��F�v[�����[��Z�V�-&K��˺}�������ru�\k������g�<Vg�'M¯V賽�t� u�yuvWs�gpv�R�Ϛ�Xӳ*3�X�|jC��Sn��1c��x�ť2F��Q��� ���ǭ�z�]�;v0���ZZ乐KX��:60�R��WY�>tc��9e݌�k�5������=tx�v���MF�z���<��άu��Q�p�6�y�s��vrvbqV<�\pW�^��=k��D�y�c��'�;Ԯ����ژ��N�mli,�8A��s���5q�X7#W��˹gl"�\�u�ݐ�k׮�#�דu����.��[���K��6�1`�8����;�]��zx��qا��ڭtkA�z켼��;Wn��HH���6����%m�utcJ^zup@خٗ��&�Z�zm�i��Z^�Y�*<x��X�ZM�	�"�!$�v[���1�3���I���=��q�x�㺭ʘq��O^=�y�V�֏J��m�֋���J��<����l.4jr;��6ҷe�x�;L�yl�Gf7ku���Pnz�
guc�\vʫ�.��՞]v��Ӕ���T&mGQ�n�Om�Q���~��#sO/m��ާ�:^��C=i8��m;uY\7�|�[��M�e�'?JU��]�{gtZ;T��v��5�e�ކ槎8��u�w<G=qۓ�BA���>
)����^W�OGN�w/Zx�;r���_k���Nv	rN��M�tӶ�7L�u��#�׷ ��Q��bz,�ݰ�����V�G���0�C���*ݵ�b�Cd��g<��&y�eġ�<m ��jVw<�넱v��7�wn{ 涟hmo�i�ݷB�"к�A�E���!�4��zJ�Ƨ�ls^��ۇf-F�mjt�%6(�vŋq���j���W�+���=����k[�<�'Y0�Dڲ�ڊ��B�-dǊe��kok�ۉ�7LOE�'O�Aͨ�6#4]�๩���cc̏cC����í�7�;7���`�1�vݚ�j;�2��i���\��rtA�y�G�N5�t��X��;��Ó6�n.5�z�m�rs��7k�������C\G���a���q$�=�N��;����z��<s���q�����l��[D{qs�BU]H�6rZ2�i6�{��5�dm�4��w&�P �F�=�b���l�w|j�;f�q�� u`㌶2�|[�~{b1��m-ۃq�]y�F�q�UA����aZ��냎���6u�gs�mYS�4 ��n�es<9�lE�[k���jIP���{s�{V�����K�q��q�1͓�<o<�\v�z7T��b�<���}�D(�r�04�v�w^&Qx{[�F4�zl��������]$�քk{3�8�v���7Nx������Mңۇ<���yz��ew���wc�vY:�9�9�ػs���1k��ڈ�,��;h��}��{g�b�L�;EOM�C��S�m�N3��\���ƶ�C����:8ݛ�'��Zx�w�aָ6�>R�;�b���TI��y�:��L�"����Óۭ�n��v�s;�gknNץ�k�QŞݵ�{	��2�kqϬ��Ʈ���7`�]���9��㭹�`xz��j�s\;�ݷ�z�8�gv�s�k��q�n �۶��:۴����-t]��z����Q���e�,��H>ݰ񴫹L����O\<:,�uG9;n��������n�ka�G�;A��1���k�ugm��Px�����W�m�㶩7�I���'GFUoqw;Orw��osb��V9��U�N�.�ݷ�x��ݛ�`+��"6�n:�Q0M֬6�qn���.��y�`�=bC�w����c�NCs�q�����<��[�����/ ck���FΞ��+ks�
nv���.�谅�v���q%j,�v��Eij���h���ҳ��>>WXkc�����]�	u��v3u�vg���:ٷS�h�)��yh	�u�vn���x{n���vq���o:w;z݃����WU�=��cG$�p�Q��z�q�ƻ����n�S2��#�,q�nI8�nؒ�b�13�v�����`įn;:��7n�l�a�O�v���z�n7��K�����	�ջm��V؞�y��Aon��9�=��n�\g���ZJ��P���!��u���.�Q�u����qa�I��~�������uZ�;t���x���b+u����mt���6q�j\��u�5��)���`]�Y�vx�����[=��b�1����+�l=��ݢw:�-�s�H�<&�i:62Ë�[�!�]vR{7g�"CH��v�96I���z��.�ֻЛ������lҝ��;��qA�y�F�u[�]u�KgV�t��ظ��f(�s��{	�uUٺ뵶��*�dUW�t窎�J=��3�f�u���g
a����ԓ�x�>vpm���Hz��u�g"�m�M��ذ�9����^;g,Ck�۱�9 ��ݻ��T<2v�ڶ�v���n��{a�����!�۲�]�\<:��;�9���ָT�}qK����Q�7��w76�-��:t�Q�_]������]��Vz�X۵�ۖ���A�5��sun9}�М[V͍�'�Mm�p���F����9���}��e�dP:�8����%�����#�ss��;�S�2v���
��m����ɣ���6���#�����9�ls8�b��mu�l�=<X�}��������]��G�n{u����MW�·ܽ�=!v���v��g�ڼ�4���J��U;	�!kck7[nj塝�R�_=n;.�^��E��c��u��{0�`L�[�c4G��G�6�(lr�9�������sоq��=���R�ښv�5��X���Te��;�S�8���ڥz�3'ngq�Q��On8w6�vlOn<��<vj۝e��7��R����B|&]�I�N�r��K�&�M�G&���nL���::����uծ��-�1X6ۇ[/=��z��!��]�KY\]��w�9�p>s��� ���s�s��89���p{���~�_�_�������������������ڀ�	��	�������UR�xV'Ĝ�Ԩ� �Yb"j���������������������������Tʳ�b{XI����tt���س�1�Gv�#���f�\mnl[�ڞY�n���n�.�OgM��8��c�/[�f��j���z�H,�Wk��kkՃ�[�ݺyr⬇5��dŎ�tw[I���qn���t�^��ɹ�S��F�lsv���1���<��fM�����z8�9�������]��ٴl^�3�1�۞,���9�GS��=��{s�E�����ڕ�:�9-����X�h7'v��yꍈ�c�!밫�z��P��T'9��>&�ޛ�96�+n7GM��U�{'�vF�����m��=n�B���=�<�۴��{rfyϮu�:�t�֍sm�]����8ɳ��Q�N'f�tլ�26`�q�:��x��gc�4����cc�]ǂa�����r�� �l�@Osv89�����y6뮂�wNñv1�\�<���1��&���Ƿ-�H������C�x�[�#�ݦ0�u��m!vu���[�����p�׷nJ|T�n4�G���e1�o	�r�ۥ�уպ���=�����5���nձ���btv�]��h�Mm:H� ����j�G��I���1��h� ew]�He4&p<n���n�s���M�5���Ř#�ܓ^6���q�+=�f���|����ۨ�H�5G��ܜd:��zM�/A� �M��by�zח��j�C&�P�N�R�l�Ώ ��b�݅��\<]˶�q�뮔�ތ�\nE�c�OcË�-pmғvd-��[n6��p��ݲ4q�SUӧ4�M��Kh�ʻ[8��x�i�67`�Z�nk6�ε��h.��φ7mq���d��P��^��h���#WWO�E��\lsڰn�Y9�[��஻\z�֛#ѵ���l��	��O㣶�Xٷ8��'�f��{��{����x~����u�
*vɒV�����N ѫ��5�#�EǪ�[k�=��7�m��rݣ:�[��ce��ݲ�9�N7�b[��+շX}�pN�-��}���]�N�Pnt�\v�3��s�/��&�0q�'�n�Ƿki�IO]p;n�gYȡ�['	����vŇ��1μ$ug����Qz�u��5��\8l�\XL/A�w��9D@3�c��ۑrx���p�<9۳�;2<�yy�"x^�����[�9�����~���oZ;mSG�yc6�կ�=|�y�{�~��rQ��Đ���S�}:s��m����ֆH�OV��j4�;#"q�9�0'dN/��ysMvm�B����D�Yg9��{P��^�浼w �W�����9(94�>.X��λ&�-��(�R�b6�o=��Vu�����s�Z3u�E�����������˸�͓sfg��������"���r���:��mn��]��pq�Ė%ۚ���^̹�W��7t�L7�kP��Њ�U(����Zړ�Vw��vՍں;]�{>�v-j�����2,�UJ:�K4^].j��˽�����Z%���=�G�����k�^Xd7�-�7=��yD��AR�[,{̳S}���ˡX�X�+�H:����z����l�ux"�ۗ��}�X:qҌ]m�pi:/z�:�'o��t��!��dt�&��ɇN���]���ȩ�6�Xe�$v,�!��7�<��~Rp:r\��\�����vC�Чo�EHm��i��1���nI5fN��2�����ͳ�qvo��K�[�C�8��4���Ѻ���x�CWn 1%�E�b>uY�m��AUZ��+>[�PP%�F{�j	<�.�ǆ�� �/WZԹ��'#i����Dۥ�m�7^��ֆ�i��Փ[����#�<���]��q���	�6�Fn�|V��g�����Ss=s4mIw��H[���y��0;�}���A��T��0(�f�G��id\��]/A+Sw�m��%m��Q��E=���b�&�1�����W����B�ǧY�^v���m�#�~�a��6��gU-zEץ�v]�g/�BU����]7��OR�}�(Z���Z�]��˗}�S0��i��T��������J��ܬ���k�0/L�\�Y��ﯻs\�޻��J��*�	r�A�V	rSپ�=Q���{���]��v�:	7�}:����U�@�^ĥ�on�M����=N��K{W��DVYT����l�U���:�K��`8����u^��-��;(�W!���g��-��9Q��<���;}���;W��N�暦�-ũasF�������+����Mp��=��Ae���Ӂ���s{Pt��u������~��cn1!��!䩙:�f��@N��cV}��L��q����Sn��RB����+0x�/ze�X�*���M�ۂ��ܕ�ìͿ{��Fȱ?-�n�ʰv���,���sӧ��a�7��5
�	��6TR0Qi�̿f�6싑�O��k5�#d�3�e]h�Nf�{�mz��3qKԭ�g�����;����ES2�Ef;�V���p�K"����2o4�0d��-����q`F{B	�c���{N���ghvĉ�ݶ�B�bvM�T�=ŕ�6U��|���}a��8}�5�*Y��6��:ݫ�.�7�M�c��(:�}BBB++�L��=Y�Fz����O'����_۞��%Iţ�:�x�Ə�'�>Vx�Ch�@���z�I���9�^ܹt}�V֯�4r.\\^3���tPm{����  Y��kw��vr���t���$�g�����Ou��5�n�͕��27����:�	0i�P��F�=Ze^�y�NU9�!DSW�f�ڮO`��0�ʵ>������0�[iyHq�nC�1�u�������[�sY�ݳ���Bd4��a���[�SBJwX5{r��|G_�� �Kc���9�ә{oF���_�Qs������r�S��9/U��^Mn-݈���]�nP����zN�=#�{��ث��'�&��G(��<al�36^J��"�8r����#SV��a�k�]�HnIwn�����h����SUUUUmn�������#�bnV��xIv#���@B��ac#n9-����WuE��=x�vpv��#�-��<�zڭэ�l���9����͸���^3��la��=gm�	{nvȷ�z⭜W'=s��+az:ܜ��W�`��3S���;f���5379���n�2�kp���[�=����\&�tZ+v�\�nS6�D�s|w/�G\�5ئ�NH���ۮw7�y�@D���x�#�) )%#���X��k�ڽ��iWCy��鞆���c�z���BѼi�a7��s;Nyw��Q���R��M�<��^�y]5�ƶ�e�39ħ�����dw�+XT</�`	�N�p(��<��nr�R�0���rH�1�2��n�A7�c���H�Q�|���I�x�y�M[r�ݹs�B��=�,V�Ĥ�}�m��+�x���v��������8w�iw�)��7�
�L8��$��f^�z�u�V��9]7����se��ܬh�����H�z�qbqsQ1��v�w;���f,��M�A5wd���W�rV��M�/\�ݶ[��l:���[n�umQ8-�4]X)??�Ö���S�<��!�ަ8��5t���6�M��N�@�wV��p{6 Q8d�9�6�w���i�������$*Ι��#G6�-Q;�6[�Z'v4]�;u#v7��
nv��{�	eN�-���kvf�:�	xڳۈ��vɽ�x�Bnv`@���z,	�&�x{�؄a+�������sԴ'�i��p����ռ�� ��u�����}����k�ׄf�㵐�I����$e�n&㎳��pm}��ؼ��$k�B�Rǎ�T�q_�|��!����NU;�Ѧ:��D���*"Iz73DL���׽�X�r5�2���\�I���yQ}���o<���!�����M��%�Z<�$TQ���Y=�89�z�]�L�����3�����Ӽ�x�\t��d�w�6�%;}�y�.p��^"��b��xl���6��L�Z�U�e����
#q�(o�;�ٞx䠪��ռ)����&��=��iZʪ��MӬ��JZ�z�n��M�i�
��{�w��ޞ�����
��Y�e'I�Ձ|蓖I�@��]�`J\1c�9w1g&�-����]�n��ܳ�S�kk��{���ӉC���ɋ�	L�7����9tZ7�¹�[3Ǒ�C�rX���m7���v�ߒJ�OV�p�yۙ�N,��΋T}�c�*k?7���}�����T#z��l5�X&F�mIem��3���2E`T��km_`�X^.)�����h�a��ۓ���xn݂���","�u��,1�h "�I���EP����C��\ʪfv�^��8͍֝�ڐ2��R��l�ۯn5`���ܰk���]�R�,���WQ雮^_����]��F�Q$%���y�o���n��cw�b^{ҳW�0�lb�g�^�nK��Vټ�z�`��˽�bJ6�
�|P˭��R	�3�4Fɔ����;Ɋ�K�9/~;n���p�ދ�W,ß^��UR�*���9�/s�#�i;�N�,�3��Ue�4򼤗;�}Wڳ��fN>I��iόeL��AF�In�����{�K(���P��Bb��-�n���|x���Y�3�B���v���{S帬���u�<��xY�Q!�ۍIn���2\��	F�v�cg=f&M�K7(�,��.�n��Í���j�4�+�q�;�g��!H�:(�u����^*�u�7aه=������ny��^�gfp�#�B�$�mHs{+[�������=���oE��SH�����u�����O�{�c���'��8������$0Q��UF����{b��|x�< ᅅ$�T�M�[�є�≈�I��q��;��h"�~Y�q�Iw�^����L���5�Ň�=2����V{w�~x��`Ƃm&�<`�����Hy)�+��ތ)g�d�I̹;y3�Onʺ�2Rl�Aއ�Qz��i��ǧe�dw�!�� r(����ݪ&�b�H�=ɚ`��I]~�zn��w~Ij��-�y&���#n+n)'�;�ƚ�n�Ӽ;`����jZ�̎��4��}b���Y��@�wR��f�e����v�˟���������uUUSs�&�D$�UUUU�S*��8�Ƭ�6Z��O:�d۶��x��=��˹�=c��'v����5	t�d�I:}tj:�n���v��v�꣞�ú����{6\���E��Y��|_m�zS�k=�x��4����)�<Fr;��;�N;�6��$��T�s���=�܏�s���gKڝ�4�|�HW=��6muin�vѨ�s��_C�5EE�9I]:�st�)M�+�!0��[��2����]��·WU�8+�V?{����Ҏ�[���1vO\��t �x׫<z� �c+WeΜ��ݚ�#�d��!r���d�kzk��_k^��p�5[���_��ϱ� ���K4�<Gj���:T�fS��t�o6YY �i�q��|���;����ڵ�VoNdwu+�[ǹ�;z�a�I����^���^�����Y��Q��8T���ll��(�<�+���Q\O^Iϥۙ�ר�	�a�YV� �?4����༚Han0�r'"�w����.����V��۳�]t�v����5y��Zl;�<���:�LK����E�q��i�lV'��)a���������������h��
�n�ӹsf���`Y>�j��*)sۋkM/R~N��O����j���R7}��,g��r�=��cJё�&�og}�]9g/��u1�J'B�q��V��a����"r���[g&J]L�Xa�&�[�J�n���5mn�N�)��6����9����rwjf����T1eZ��ۺ�s�3g��1[X�n�j@�z�#i�Y�n� �ʏ��M�7yV��X�5���3t-�'UlkN���4��,��)�w�~��#��t�^��+��6��F�r�=�\�W����;���9��k,��*�?<,�n���W��p����G��j	z�tp��#�z�=��i��;2\�BT�K�On���x�-GҝyUy�=��㇧f�=&/S�ki�F{6�b��,�3��7:�r!�]n��X���_�^)-� c��t��ì���n�ש��L�{.!���\W���/;��ݨ�`�"m���JwW�^���{ ��:��9���(��6ŝ�bD]W?n�ڼ��u�˾�=	B���c)n�R
0���n?+����V��W˕�屟QY�ݚ���l�wd`:���c�ͷuՙ���޽�(�WTK&�,�	Ź��q��j�^�RX�[�a���S�����i͉�	8ة�Z��"��_n�{�a2�j_l��f�ʉU�Z����Wt�+��5w]FR�����3���d���R�H�w���5Z�l�Ҧ����[��w,�t7^.͈�\�7�m���C��8ٛ�ZC��"�95�v���-���Y�ʏ.�țE�ܐ݊θ��ќ�N&��͜w{�v�YAr/.b9�n����k�aԹ�d���f��ɩwGά�8ՠP��ٝ,RO1��W��X�EXG�=�f�(��g	�.E��}p+�Z���Yݰ���1�x6�!|e�9��\ջ�"��Yf�uk�6���v�2�@5l3����}���13me��WQ�v�oh��g���w�弯Jʝb_bǺ�nD�<!�n��Ǆ��I�>�R]��wS��K�	w�5r6uoV?��h��]L�h�d����t�zw0���<�7� u��*�J��B��I �^�7�!�n�t�v+�(��xj�]��b��e_f^�g�=(p���0HҾt�bO]�p��ME[#̒��75KY�z��ug 1\�[���B����o;���E�u1d�oŚl��!�y��t�Z�1����7Hq@�����ʘ��8l�Nwv'�����Y����!n�f������o��na:<�*�K,�����ŝy�X�g��V�~�0|�Y��5n��yϺҎ}{-a��n��50��MM�\�罳ܥ�"�J�m���b�2����iŕ�����+���2���y}�n{��22on�#�ǁ�ß�o�?���\��nغ��h݋�f7H����Í{�c��}mZx�{j���>6m��9~';�{�dշ���bk����k�{W�ش�g�;��b]�&C�Mw��p7ih�ev��Nw�KK(^���_��`�OY�ݏ����9�D����%���-
ˇrl��`F�H��7dsM�P�/W�W�y��:j��٠.�"�tĩc�Z���4T%�R@v�U��]�]��L~��ޙ���-~>�X�EV���A7Ȥ��o�F L|lk�.��ʷ%���{��S�'!r��arY�Ñ��ʋ],�D���0Eg����In�U�. �{����7�Y�z�a h&��8S��n���+=~}��:����Qj��
s�������#Kǐ�^/o��{ӥ��g�ȡ�[=��ݷ:�q��d���\�:-θ��SԞVy�u���9�*��tˮ�d�>��?p��Vg���X��O�=�5m��*6�TrH�$0в��@8���htX GJ��H�1���y�o��5TO�¢�e�xX����5XC65t�u��VsT���Z����dh/֎�%��^�]���WL���U=�3뱥�/��wd�!wn��f����a(�> 6M�[��|��x���u�`��k�r.Z��(�ٽ����mݳ�2����O'G�N嶹��P��(�I�"c[ʦ:�v�6нs�������çlþ�wlδ��A��[7}�/&x���g ����3N�<�d��Q�U����&�Z3�f��r#�^M=��jMHu��۾�7;�F���!��On��$����Qm���Z�������v7=)3v��������R�N����j�bj!85Z��;wng�qg��p8:�n�Jp�%�7n�ہ��+	[����,V8�y��>�7kZ��gre��t�.�Z�[`�
q2�z�<5pcq9ݨȅn5�]p�\���+l�w+�JyrH���N��uuF�tͰ�.ѕ�]����qg���n��x�ƍ[�I���7<ٮy��6nd��u�vu(V�ncgWW�h;Sq�7cѱ]��VB���o���n��徛�e�w�}!VVeUѮ�}"6�Y끐�+I�'"�Sh"x`2IA�����[ڱ�3{�c��c>!UN}Z��GuF�k�հ��gL�u�'so�u{���i-�E����f��iLR\�+��:4�>�**DP��ķ�8b74b��ж]���w���B!�l�"��M�>�ם�+b�>�(0f��������5�}��T<�5�.�<�D��Le8/̨��h۾���7�����R�f*��2Nd'Ԇ��xqgA��˜#�ү�,����vT[lh��N�K��#�V� ����ui��;���:�uQ�(I�a6�#�1ǔ���h�"���}��ѻgH�mw�X(�
�sB�oYҽ�ࡇwK����F���p�T�;y�^�u�$�G�AP��bZ��X 4�6j;�6S3�}��d�����t������.�I�9v{4�l�7K�F��C<�zK����v-��/y��ޝ��y��uY����|����{�'�m�RR
�Yf���ش�/辄a/7�5�:��;�qf�Y�+gm�˅�_[xGe�A
"B�%$%nf�ˠ����w��/M�z��d�κs�6*�0�[��gc��fn�c�q���$�R��J���;��+<*�7B�+0�{�/A|x���%������A��-.�&��j�����|?�UGl����v���تlR�����9Ϛ��نٱ�6���@�k������Ӄ��}�-��GB�Ȁ�OkVV=��X���۳��u�����_y�O�#��Y+�Ul���Q3 T�yU�gJh.N���_\�\s|}R�W{y��x"�h�yL'�["N�pd�V�C���݀�S;�m�r�˥*-�k��lQ˺.AcG�oY�lb��s{te���w�����A�C���d0b�`/x�������t�:X���p'����t	��VlY;��ǲp��ކ�����(f���jM{B�y1;(���B�\�篽�ލ��Z�V[e��M��)����9k�|=�ƨ�m'K��z=�X�n(��o��M�vy�w�k^��y���w�M�$�LTi���.l9����zoK�Y.-�&���#l2����[qũM�
�P�rw�b����;�Y������;�ږz�3|���e�#81�yDV��
�B�BCMG$Zr��F�}�5�6�a���3w{��r� ���۳��DI�HWV]��3���u=�x��:0D	A�T���1�~�����];��y��g]
:7w�9���i���*�S'�n�y��V4¢08�a�!�=��x�	�c�>����D�x����붔�YYwPW��Ξ�wk^�tg`}�A5x�3���g���Xb2��:1��v�l1C��ՙ'rPuE�I�&��]���v=��`p�c�HKa��:�o��]^W+�ݑ�6{3��.�#Τ�Qƅ�ݖQ~K{�^��3�w:�]p<7�i��Q���AA-����9xzx�W�N�+v��U��<\]v��� Cv��gj
��]݂���B���T(�Oi�MF\�}&Z�)�����(��;��w���&�ӄ�S�v��Uߧ�G�K��0�ǩ���u9�k�2���]k{�-{Հ^o`\.�hK�҂&3��7�q)fi��{�qgg{�+ٖ�I�f���6�<����'���]��㹼��k~������A���鴂�����D�mج6D��+_m5�)�b{�hx�t���J���k�ȷ6�J��LyJʌD���������t�u�y�V �a���﮻Ոy��,N�w���+���vW�n_oa�k3vc3�	:��;���nMʸ�:4�77&�8*j��Ԛ�A�,F�/;r'8޸����0VN�I$��uTptŏAUUUUUmN�8�z�t�u>�n:�����۝��CY��zޱ+nz�l���^�R���]p�����amy#n^�Z�e��\�뭁�V:����fb�|2���������vwXO=��"���A��ѱϺj֕���o^��T���ݛ���v��綮5�N�ʳrk�����|�c��\�J��v�stk���vv�����S�X��ke�
�痣=�%�Y���������E&B�13-ς��\��z;��I�Op��ɡL9T�[����=�&w4)m�������IdV"�^m�[j��_��|�g�9���`��T���`L�>�2��7�;���9f_�u\��M��
�@���"��oS���ڷn�D�o�C/f�06O��Oޤ�n{�B������5v�썿V�E-7�8dNC{���~��ے�+w&���E��x�eH(���kC�ۯ+�}إ]��xW��*ge�yE-�!�@�rKǛ]�.a�4KP��㠷�eί(v�5�t�`=�p��'�^rn�;W͎ȇ7��?���N��mav�unݻ>��x��UŜ��u�	�5F��]K��/S������;;�]�5Pf	Y-C哉"xR�P2:��L������d�Z�7׻��S+�"�ǘ�w��N^��<`��m��"�+Qq!ٗ��=Yk�CJ���Y��%'V��Cт�6�I�X��l1�v���{��y׮����Dy��'��bلS�"�:Y��y&n�����3��!7�g�}��h��v�r�i�g̣u�w��;��Y��|�a��
�6��\W�2	�ϲ�a�Z���D�(�`�	�^cX���\��{�o��t��{(
�Ot_Mg�y����d���G�b�E`aGjMB��^��߱�,u�(�m�8�?k^�͂�8�c�K�{����w��>�g��t8���lѷ4.�����{�P2OJ�Ξl��܆l�r�:�����7�}k\6x����+�(Z�UI�wך�;��K帖��๖��Y����jz�ܲ{�K�W��-v��V��/HKA!L�Ґ�7T#Z�2y�x�^��|sYn3G��8v�*�bo�]�tz��锇eו���O!���[=]j8���d{�	6�B5PM�y�.>R�����<Y��]��\�t�ۧV/Ov��"/�×����˲���Ɣ���ڴT���6U�"���ԛ:�0Q[���`�A���%�-�N��z+9��i��<0�F㌐Y"A�i���V{X�SD�{������u!R�0]��c����#E�{g�	�x��6�v}F��6
p����R:Ȱ�:�I�zn�'=��V��`����R`:=Ѣ6��o�c�g���D��w�r�5��]6��!��Nw��=A�ی��ˋ��𖛦�p����"nݗV��9�(��{^�����=����C/:��:���4NK���l;k��.�=�-��(K-Cj)�]���A�^�m�Q����d*{J�Y����u���#f��?(�%Y��d�v��録�j6�M7i�-wB"\r������� o*��C����W6�N��ג�V�J`d~^H+bnđ9l�{�zy]�#3����C����6�	C�i�X"c.n�{��<�V|�k�]5�۫E��ꛎU7�IUK�4�*�
=���jw�V���xƗ8v�ٻ��mk��N�-wz�r{�ۏ����A��TT	�7l��c+m�>�P�{x6��e���=�c�{{:�/�𐺅�������&��9�&�0���TP�)��Ӟ�l��\Fq��ݹ�Ԓ)b�-;5�qF�rN(rI�kn��׽��ԨΛ?vw\QhA�-�,�Y�=������W��ܬ[�3��b%��*�$$:~���p�M�r�l�[ >k��-ʡyp7Z�칡��F�`���9돕vy�}�����y�a>�4�D�N<ό����6=[����mvzK����:��(���:�<����#��C6;a��M{��Z���,���l���Ay��|D�k�*��^+w����piڽ���������p�8�y�B��hV'e,���}s����P����u�J�����E^t��H����[�Ftgv��fމ�,���rv�!������5A�zm���qK|��:�����r��Ò��#ٳd��Ӂ5I��T�57�u~�/���G����mͼ��W��#���^o�u*�r��-8$��B��� �N�W��3{!���غ��p^:��M��gXo�Z=��s&�VoǇ2��j^�ʹv�͹X�+���MElG\;��F�ˇ�p�����'S`�3B�p%	1���]��u���Ψ��b��n���w�6V*�����[�k=���nX��y��"�PfNΎJћ�<�w�D�t	;w*ʝf�Ϙ{��y�۹�H�se�ꥋ!��@�GʛnLTN<;J�)���{k1TM�z��F��5g��퇜�e34p2�/	�F�#�����o8�3j)��^�p�)8�9ݨ2�hѦ����ؓ��*�gm��QP��2�T�����q`�����W6�i����������Vn�DNG�9���:�Bgb�#E��R\Z�ep��)�b��.c�ʝ�=1�)�o����;\pf8A�\*�&�>�z�L�g&���uf�;��]�����/h�?i�I)��}Z��U֥�e�f&�m�v���jm"&f��VW"�eq���K�X]eYZ�p���k�ݞ�R��q0ݻ�T�|fk}�
�Kv5��"�d滯uǶb�Ru��.\�����U%�xlK�]1zz�
�V�c�����r�.�^����M�ÃA�]ԋ^I$�I$�I$�I$�J����������Wb����/ �LYZ�����*�U�X���A8��Q���´�UUUUUUUUU_ʯ���������������������Y`�l[�����Ǯ2�Mq�n7
��y|\]��tu�D��G]l�K�7Us�f����N��#]lm����s��ͺ�ݎ8N�n�c��f.}vc��qг�����d4f%��X���{6݀�r��鼗7Ro�{ʣ�u�<v��4J���Q)�&��M�s)*	dg��[ȥ��2&���&k�s�sۡ���:�w#�8�q�WT�u˹7�g��N�vo[��ʓ��w AE�<��r�g��(��=v�����F��i ���w �ݷuf�_l��� 0�>5�8��ְΩ���n�.�$v�������^�l��X.��m��<��[��v���۞�aG��܅wB�76�Z+��;���$e�K��a��z���m������m���<<c�\�X\�C�;l��n�������v۞�u�=�m̈́���q�nI����C���C��:Ŷ,t'�k�b:�b�����ݩ뗬��ы%փw>D魰��x�=���:w<�}��9�����k�q��������ۧ ��|l[�dM[n�m�#lv�a�q�����,q��ʛ��Q��ggi�v�ɰg6ۻ��whQ�l��9+u��{EY�u�Q��3�vMۇ���[v�r[���U�1�K�]�7��c��N;�o��m�ؽ�;սشk�j��\�f�m��g\sn������wl{��ͳl�n��ɶ�v�C��>���PX1�!�z����sn����h���L��t��`�����[��X��/�\���NN.�R�<]�{%kn݊�;�}�λ���n)t�]nKóF����:�Q�c�V������{b�x;R�4�ݴ�읅��!ݷp�z[#����Vz�8�>��΍b��]��P+�qY��v癅�n I��#��x�<v��9�m
�pQ���Md�(N\�N�VK�!a���غ��Z�����V����5UUUUV�xc5�9�g��W+��A�˸���i�Ut�	��p�r�<v���������	z�[<g�=�K�u���E�nۊ۾�u��>�K�����-ǈ����=�XW���l�R�Ml��0\�m���<�b�67O7[�q���n;f�wf;2��A�,n.�Ǭ��=[����.K>ޑ��la�l��]�W=\C
HۧZ�n9�M�sË��n�����]�z��9��M����\͎���;HZI����קљ'��쳖#ofȸw��2rS�����V|�=�B[��Ecr@������%����S=�:���-�^����M�*��
��Z2�����w�a�&y{½��}���rX1�!�53-��}7�M���x-eg���%W\��"�Mȸ��\²9�'�~����)m�{۬�#���՘��w�.�ǎ�oM���uj�oCl����l/W��r����}m���$ƤW����@���=x���6Vࢧ����!�("�Z������dh���f�b憯��Q?z�U��;mm�c���k�x
B�Y�b�9$��\]rP�l�]��gf���tk������~N�S!���Jv[ហ��
0��F;��ܷ��G�[��z�G�&�YQWd��f��s��ű���5�iW�W�]3�=Y)�,��v�n����nbm�XX���0Fw6m^��q�H��8{XQ�Qr�/6�S�R�	�'�����^���}�fr�������g�.?Te�ms�������ӎ<h�}��|�,�\���=�g�������^�6K��6�}�����kf��]�+<Oq�#H��lF6|������6g��fyGzk;�5[����:mt~Y��ݭ�3U������w|w;�|D���iet�Ӝ�?��4�_+E�:h���8Uk��M��܅eڌfv�=��M�h�^�ng{ݞ�q��q�K-#V�-���O���vh�*a�	ܷ)��)�c��8���ؚ�=��8��(d�����[�so�w҅/j�8'��6-˕�Ov䪮l�7�u�m��qo�R�k���y�� (����������ڮ��K.^`}+��z��_6e�ќ���'���]�%�G{.���Z�{:E�X���`E)"�n���}�����7*`7�;뗮x!�k�Ϸ*����mQAJ��h�gfгͩ.w8�	�v-`�o*����]|�<b�e�h��Cv��-�i�fۻ��&��:K-Q��ɆScN�-I���^?]W�gh��7J~��P��+l�u9��Yq��Y�xl�3�z�*�k��^	C���"�̶�&6Cr7�)dI)��t��	��t�e��±\��]`��������9�ٻ.�;���B�|�i2^�Rʠ�������nn�wb.7;�]n���s'ctB�џ
��e����I�d3Ox�Eg�H��x���S��Po{'b�7�S�	QD�n�̿\9=~�����60�����d�
*�5��zl
��S���4+C���:6(�O�Q�U���cU}���6]e����蜉0"����.�e��~�Yb�ħ��E��{}{����b2`x+��M{G3��S���qaQ`J�V��'^]���rV_Tg�����G��-.�j�u�w�hk^FW.7׸�Y<�rj��f�>cy	�m��d��2�qT�pJt�gPO����}F�̜,�Pwt��f�LbV����ǡ����i�#��ڍ���H�m��ˎz�3���6�c�9=�.�X��`0F����0���y�0�
�(��x��o��ži)$�B[
��i����ш�c`��4��֤��{n[�#�hn�/\�
�u:�Il�p��1�����mg0�O{R7�P��������3+a=l(�G=��3�h�z�"���|0D
qe�sG��jy���:�4�h�����[f'M�˲6P�1�m���������uШq��FZ�Q(�ݼ����wd\c���;�W��}~��b���.�%�Gj]���[Z"��R��R��g���uLΜW~��k[-{.U�����Df�휓�3r��K(�^Rc��A#�#)"!���x�o�ëS\��h�f�V	��ῇ#�)ͷY�uq�"��cO��5O��.�Vz�G�!n����]�=F���u
oMp6WQ��;W5[�Qc��{`�\���S��9���UTmS�fΚ��������<ܻu�lޞL%v0�n8n%��0q�9]ͧtc��Wgl�.Ս�e�X[�m�/(��X��n�ڗR��lZxׯ=�Pۋ�o����L����ӻu��nΐ��6��%ÑDKʛ�<��2��d�N7X��\�h�=�g���c��O�i�0���g��ι�佰S'���������$�iʜu�wJs�`�m�����Txm�n�OX`�G\����.�����8��iq��aHN��ږ��������������.v�ı;��o��)�O��O�WY,KN���s}k��;�(��T��I�&fd�F��9ܨhm5��֪K��T��!`���m�U�"H��+=
�������o�;f��C�����.�1�crK���х�oΆҕXL��奊���:9{�^y:b`�k��kٮw;�U����ۨ\)Db!I"�n�X�\�ct٤n���ȼŒ�4�����#��������{�h阹)V�/�l#��¸�����wn��BW�j��5��R�Z�\8&'����h�hVz���z��4�w�(����R�9-��iT�����u�m�z�e�Ns�C�g��<�S=Gn��Q�l��nJ����.�璵�k��^h���ll�yy,�}U�=��T���NM��_N���Q����@\j8�®_�c�z˾0��=����WG7A��@�hj������t����9��<o!�P�M!
��q)Z{5��h��g'��w*��B��;Η��dQ�=S�`�{W�k�'���kl�a���蛲sV�0gH�&(��RG�T�t�:Q���ypyK�ڬ)y���^]Y���Zԩ�$-�o���'ղ��zlIk�K��C��\�a�/a������	����.��͛kD^Ix����0�!����B��W��o�+r���}g��HB�N	Gr�<#��m��(�@?Vy�k�Żp�ؠ/�Wl/f@���#��;/;��:x�y؛P�f+z�k\pl=E�N#]D��p_������e�j�	�9KgBu��#�]Pӳ�>W��׎�~CL�o"����B�	#���������[�N�#y���/J,��^�dg6�{~��GpL�gh����z��$�NrNz� �؊�yӗ���Ynn�	K賆z��\xݰ�7����1rۡ��������ٺ�P	����vSԳ:�_׫�iD8��#�/�(L86���"ܳO)v��0�WR�y���E���ɠrC2��7%�fR���v����+`�nKZG��{n(���Oo����(சy�gyyY�z��/�F�|�N8�n��%���*����Y��-��p�A�V���"��u�|���f��}�{/s�\f/V�[+�J8Vxk�ۻ=�c^�$n�ݎ�n�K\;��S�8Ϟ����#�L��i\�;Td����U�teɜ���u�E�m�ݖ�c#�)vXD�1U�ݹW=�y�e��ި��Ĝq�
�Ʒ����]�7�щ��}PX��g�M̕R���>����w��g��g{�_�Le$�S�"��'��Zn�Գ��n�����6�˓_���f�J���B��LY�	�b��景9y�!Id�[vo~�4�*�MI��B8-�cE�Lg��-f��_���5g�!9H[�פ�gղ/c;�(���ɂ.N�Z�цbw�avћ��ų���a�g(�`Ŏ���vs<jۀf�i���Q�1c""K��;�&�6_T�<q$͸�1��	������Z$ӂ��*�����os��P��L2B�ç�ۜ-�;9ww�{j�1J���ڂ:H��7b�u�N��Q��W��s���#�G\m��P�v��2��ձ�-�'�/{�A������f�C��r׺��ǒϏe���+�r}7Y�5����e?��5��u]����{�:�g(G:���&���zZ��H���RFD�uP����hXo!Y�h!�1�˄��q�}}�꼮���9��|��V���P�h����J^̾�vo �����h��;,t���p3 r����P�Q�3b"�]�2��*�'w��w��w�I��ܪ#�Hw�|�/��6��R���c�������؉�"mw�.�\��7�Z�^RM'z�.�oζPcM�H֞�$E� ���A�s7����J��I2E5⮰�7�"go;[���'1\�͙ʻk575	1�����}�~���UUU] W<�Rꪪ���j?�����D�a�3�WF[=���ڑ��G��c:�τ��ulv�z(kuւ��n�������t`l;ۧ7X-�Nħ�F��8-]�nzأ�%����ت��I�ۋ���1����+�eS�0����^��,�\>wr�IY;n[�c�s
W�����n��C]5<Ar�:��g���yِ�e#]56-��nԈu���l�nW>c�;�Ƿo��[�yh�m^)Z�Y�7ie�`��7}ڨ�&q�~�+��d��7�e�)�g���4.0{�돮2��E��6OG+G����n2˒^t͕��u��ђ�[�{�<�Av�g��n�˔��OFF�c{�C���IK�с�Bã@�d�Ú�}\&���[��x�O�j)�U��2����z*o��"wv*��/q��C��,H�����X���C-�n*w~G�{`��T����:~�w��V>�Rn$P��Nd���y5��
(26㱴���P�}�9pp��yqG*�v��7�7~��ty���	O�-��ဪS��	]~�{ힲ���=<ls�p�^��]Qe����k횉x�����y:�����jG�O(���¯ư]d4�7��a{A��aI/~�V�Cf�ݞ�&�WϦ�����z�tvp�+j�,�K6nϺ?�v����K�m��Z���:��u��^c�Z&\�(����V�V���T<��G��V����ވ'(���\iYyw|w���J���fs>1����/���8lD&�O�2�f��f�-R&b6�Q����GO���ߝe��W�0�N2[u�~w�D�/��}c�T��|��]2:r��]��/�q�I"�7m�eÕ����ױᘼ#�nyd��\����\�>��] ���e�j��︻)�;E��6�r�BSF���' [3s����	,7�D��,�uh��ߝ�����V�0�ţ���eC,'�P��r�l����7]�7bӗ�wgC8<��m�㋊����su	��*Ho�l�:�{����G��J}*2���O�b\C�<e�e�h�w]W��",��y���pHR7	-�e�b��mi^�����9�Ub�oC�Q��*:��e��!�����8Ry��T`��v��M����5���j���ϗ�����Q���� �U\�~�F�d�/���Z���cl��5t��������J!�[Nk��VV����K�۫J
�Ҡ��� 3�;�{�\����v�̖E&j~��}+���Nw;0��c[[kL�yPLC��4J�� r��ֳ�:zu!$L�r��'nb���t^eޗ/��;f�)�㛙ca�.n�cm.� *�u fA�j,�FWrں�����Sy�X��▲��gd�)ԤX��\�o��t%��y�+p��Q_bl�%'4��c����ƍ{�Ս��Q���֣rLwM�]���2�,d�l�Z��qp`�(Ԣr�+Zs�
��*��2A�U���p��j���4��F�.ileV���*��?VjM��	��nƤ}��뎎�{׈�D�ƠJ{Ub��g[5+�E���V�	��[��h3����?��\P��=���3;��#�%�!��6�xqD�R��N�F�!Yn�Q�]p��1��5��J�xPoc���ep
��+P� 0\I�-jD�7���[C����Ӿ����3J���]��-u��Ա�;�B=PN9���^
R����Ie9f�1K%6m�ե�֦lZ�j�Qi�=Z�:ڽ�o�_l���$�r�'����+��� na�ɘQ[Q� S��Z9p�$Y)��:5�oI[e�,�pMM*�Ј�LV,˧�!�1e®	�t_P��*�W�Y:ٶ�b�d�/�V�F�Dz�n�>��v�ؚ��g��]���w��<#(6����q��woL����Q��P\�W�bХ��2����y��qHd�^ݹ�ݢ���I w��f0���	My�^+|�&T��l�f�*��yy��qڗ�I��c��y^���>���ȝ�;�~��V���姬B�s���uڻ>��F��q�"%A�W<���t��$�q�am�"��.�Vﾗb�ʦ��dN�pf���:�ܞS��f��&��ך��q�Ux�􅘢2�1B�N���y�� �^�0LN�EdF�o+=;�Ğ��)��{�OΟL�j��k-�2��,k����N2/7w�Ta�~��K�
�=�e�e��@Ds����.��V�\�S*��.���ቇ!P�:�d�e�T����8}4�ךȐ����W�\�Ѳ��U�S��B�~~o�^�:�yuw�h��<z���X�-��6���K5������ᖵ8��'��mgnb�
�+Ӷ��a�"�@�`�T����Zş?h�z�J1	]n�7��BZ��8}�v�C�$8��]�!���t/v,
!`UbR0S�KZ��KQ<���[l�i�o�8�=��������y[<]-`�\v�k���w��kʻ&;J�d�����%��]1��r��ںv'�q�[<]hvڛ^�X���P&����!�T�o��X�!*�O8l��9ܮ��ƆLgl�Z��*���+=�]"2 ���a��0Fdm&L$D��`�����ن�JM�S�����E9j�#$��Bf#�����>�K.�VKK�ƃ��#NE�5�� zOHA*�{��L�]|<�,�m.ƼC��� ]y��k�:=v�m�9$R&�˷u2�����w�4�^���tQ_k6ny(d�]3p���5!z����7]�n�|�(/&/j���������IE*<&���+;{5�>���z%�M�Zs&:�s6hR�Ͱ��NC�ѳ.��F'��UUW]*��Hj���*��g:[έ[�n���a�-m���m�l��ۛ�{k7f�n�n�񫝗��t��hh�;j�H�[���r�nx�#���N������fǧ�p��aE�n�s�	s�l�Z�۷:�vQq[��p޺�.;�q�k�э��Og�d���Cnt����jC
�����h<]n��\f�"NS���-�<s6��?��c���AUP�i�DQ�]����q� i�u͞��o5q�Ӱ��5�X�����O�����B7�^X�a��}��P���l�����U�����W=��2$.$ !��c�O��U�XO��ç�M�p]u�.n4�g�R���������9�5���mCk=�r�ؘ�fe��<�)��f�*�4�颱�i��d^BI�t��M�Yޯc�%�:{������5�R��Гp������ۺK�p��Y������د��th�XED��ƐWC�,i[��<X�A��E��6�i��oƲ�R�<�4}�,��\ٔ23�_�n���[M����@��J&bQ�k��f��j:K�<��lu���t�x�k9���[�񪢊��w�ծ1Yj��w�t�L�`��b�Oe"|/�Qu헓mz�m�իh�2e�ߠ���}^4����,�i�"݀���}5�G�d��y�T,NBg���<ˠuܻB::湷��*%�ic!��j^�+2��q�s7�³��ĎGz�<�iۉj���W��O=;m�ۺ$�L�E�q&u�I�<�Q{�ÂFԚ��Q9m ܍8 f&S�6��[s�xO�.��^��������'�-�	�痎�pV�8��,/B`1�FM��-�W�
��/J��Ak؄(]/v�Sdv���O�*�n�a�x{�/b��`�]
����_����FBbN�y6ty����|=v.��u����Jk�3�z&5��'���+�Y�T{Uwv��S�Q�f�Lg;La�92s
=���:�4��FչWl=m��8�o��]�Q���j��ܯ��mm���f�z�wR�"?</�j�dw>n�ŇdN!i@��7&X>���V���0T��籡�f�0L#-�U�q��v�Dv����З�5�*�0�J��>e�Ei�UX��Yy��f)�t1��x�uJߗ�^]^K�\S�ݹq�n�i˝�ga/��Q�W{i �5���a��h�����B��v��u��Y��!�l�m�>�9���2���Vb2	l9��n,v�лޝ�Қ:����^�J�]��9�� �b����C{�8a��7�;�7��*��/?��0QsG��=(AK턴�5�PW�T��uj#g{�/�\�ߡ��4�׃Ǐ��fr�z�;C͵�-Լ��[�7[dݣc�ɺ�.6H�{c���73�v�0���9A�%�[�Z��6�c�1x=ol{��}�Uv�y�G�kо�S�D aI+�.�*+�_Jr��S����xrs���=�w<��v����`����Q����n(���]k�"��@�������V����N:���9�=��f(���Omi���γ�=Vjt�7�zhN&f_��ɰ�|o�S�-�i�Fw������o��+��b.�Lg���[�яG�P�;�o�ý�b��iF;!��˅�.s(���f�bv�_24<������*Ƣ+uu;��Ec���eb�����$�A�����d<�	ͨ:Ŋ�a@�p����yW{ݳ�Ġ⒩v�7ݭ�ڈ+z{3��(���/Me�`�DW_��J��ܥ!�W�
��F���*����p�Z�h��;�YK��xt�n�6����Ct'�󭏔3-+U��Y���I�գhF�$�Fu:2uE�u9�<�cHh{
Dh�,�d������C�����g3���eע��
��m�C4��6��B�j�����l>���=�}�j���b�ae��3͞��$��Y�Y�9�GJSsr�Ỵ�-C�V��ߧ��:��#��v'�H$>E
pV]X�[�����K7׋5M�L����x���E��	ؗ� ��9��ti;��K�Օ�������1ɸ����Y�Y�ڣ�D��r,7���E�y��4uh3�)�G5�;�ގ�rik׭o�U���3{����_�Y�T7Z,0��G��:^���vv�<ifڗ{J�͠ufk�*c�ۻ�I$�G#aG�D�Ū�����n:�Ӷ��u�{�W`��.�{^���s�b�nz:pɭ�/fu�8y�1��R�wl;���a�V>�:Ÿ#�����va_x�g�Lm�l[vڝ��/'�N��s�;��<ZL��;s��Q�c��]gu`�'n:�9��n;c�x)=�Ñ�Y˃q8f�<�;�k�1��'D]֣t	�N�h�/\i�ҝ>�܍��w/l�/���ns:��9.�:��U��Z��ٞK�]��vƍ[B�>h��+��c������!�y<}����뚷�X&��⼲hE�b)m8�LFJqn;9�������Y`c�Š�;ȯgwR��c����|��EnΒ����ChU��f�d+x����p&-��Z������-�&���r��1�����5��te��	Ƅnӎ=ܫ{��z�r��Ԟ���Y�d�]��|�t���Z��X�ݕ�|f��;�w8O!�E>A	d��Ġ���֪����}���{�+.�
�2[���,f�Y����7T�Ec�o��T�H� $�{�H��^��=��:�Q.�J�[���Ρ/M��B�\�Z�BWýహ�vZ/"�(w�y��Φ�W���ɵ�fEd��(���9��wV���arCߺE5�^��/ü]6�rQ虈�^��Fl�u,|z^�j�#�}�C�*.g;��\t\���a�*FX�s�3{��������u���d0�ڱ����v�C��;C�m ��@�!�E$���Vw���#�վ�u$4���e+->]�y<,��kj�;Vd���|��N:�w\*͓bB[���5�����A[��������ѣ2�qc����⫞+9��u�s������l�'b2�SncY������dx���^�L������蜽j�Q�zcd57�(���!]�`�$���*ХVKeB�t����嶃�z8�F�&��l=u�k�/�Wv���H2(\5�:���R�/$�,�c��������;(f�Eճ|�eLm�+r�[=��
Nw^y�i�+�ޣ�-��jLCfG��!������|斻@*b���r4c�VR�� ���_Q�䙫����<^�O�=tGLT��1L�2���մ�k����鏳���;�{Fm!{�k���C#rﲮ��/iq͗$3��U�s��.�j��E3��r�>����E�׉�.�髮u1mx��֭��,��V�4�r��u��I�[��t{��g'����*g7�h�l_=�����G��A0>I
pbǣ��B���œڃ�3�^+N�牘w��[��<}�˄[5�A2xA8�T	���^-�ݺ�+�"�qt[��N��%�z+��r(S���I5$���{3|sL��߻{=Ӓ�v�[Y���yY��PT��;/��؅��r։��������rvi�{ �U�����n��q�qsX��|
��U��xn:<��i߂�#JMDʐ�Ą��O[�9~9z6<��p�,�����
�Lna���&6�w|��g�e�2���\<*b$���A�L��}}EN�n�j~z}�t��{�;��zc^R��"tޥrvG OK��j�KoU�{��_�N��NT��^]M�Z�'S�ܽ}YP�sO:|]q&�Z&�ATt��ʏR:Dkʯzz,�>1��28�ee�k�N��A�z��B�/{��q�u�齍c^�1��6�y-��V���\�%�/�-���R�~>��ce�6�&g'u@sd۞^v+�cxKGgC�=�0W+�)�!0���5�Ʊ���͇G��y��zD(Ξ�t'�Ï�6A��3֢���e�nk|y�X�s��§qfud���,��s7:������O�=�f��g��w��d!$���f��{0���a��_��Ԫ�P�$�Ӧ�էr�B�[��k7V�_l�8cR9'pN�K����{'���M�8�=�FN�L`7����Ti.�~՞��슒�	fBc�8
r�h8���zӛ�V�OJ7��ިm󺾪��W�a�O�s+~ �4���o�u���~X��ڈMn����w9w@�s6u�Օ���;l^#��:�<E&�N�ku��͝R�܎%ێ��.�c/E_K��f�h�	҅w��m���$�Fc�j@Յ���X�+W/�r�l�
�L�nw5{��gZ��0˨�ɖ�9�Mѩ�5�FX��d�0Y�m������۽���6��  �.Ь����Stf��{Jk�=����F�a��Q�;I�M��]�'(��n�I�Z%FY�V��Sk��1g	�;�O2fs��u�I�	��ʻ�S7զݺo��\�Z߉·�M�ԣ6R�&���\60J��]�n}c����Z�պڄ��0D�*�Ľ��V�9{H>�tl�+r��Ѧ�p�VRB�ɘ���}tU�]�R��9 �z�]0\f��}�Kz�e>�M=7l-U���h���@tE����L��ȯ����r�[�� �Ͳ�WӹxB4�p�Q��#�g�W-���ٴ��P��"�q�]w�e�4�B���Г�}V��1[ԫ4͆�]ioR
�F喋�g�UC7܆5z����;3�h��)�Oe)Y:4��3��v���hky����޶���e���r�ڛ��ք�*��V�8L@ִ�M��AA���s�w���P�M���L���ə�yZ�O(>��y*(�ff�G/9 ��L�V� 7��6�����>^Ǹ���$�I$�I$�I$�UUUUUUUUUU*�JFJU�!ځj������U���*�]��͗�S�aj������������������������������UZ6����<��k�ՠ9S��s�V%�k���ڒ�u!8�m�qo9y엎<�l��qÝ�ݣ�v��`g��Мz+qv�{]r)p=��uk#�㭬vJ�'\�Z����7��]�L��x����Aq�m�ͭ�-܅��mŨئ�nT�u��NM�h�n�N�ԧ���d-C��ՏF�ݸ�j|��Is.9ɇ�����gѺ���Ơ�ꂎ��$�G7搸�Ag�����x.����.����s����-�
�ۗg�Y��1l��a��F�!�m�j����`2���)��Y�-n�m9���zo#�-U�ĥ`�V�H u�:sˏnI�Xi�;b�fxĜ���ek��j�a�4���w�c�vF՛��n4r�K���1�g�kk6���VAлmq�Սm�u�����$9�r�r��>��g�ԪW��u��׷i'Oo<��띸��,n��[���i��&F��R�dVw<�p��ALܺ��ju��P;\�<�^��_;�jm�������E�T��;wnm���A��űv�1PZ���upvvB��)wX�pFŲ眂�uru�F�5�pL&�bwf�1^��[mq��bc���-FC���;��݇ڛ��gi�;x��]t�۶�q���ĜP�;���鵹9�����&�8xqg�c���vop�jOm��v�n9�=��rhv%F����=���g�z������;���=�+�Nql]�y�f�Mʚ�]r��[�5���ù�cK<6�ʜD[Aϕ86�&wsZ�x�q�;nw�wcQ�z��8��b��c��ً���V�SŞtbÎ�3�{�l\�C����y�\���W�R7�u���\��I�z;%Ӻֱ�w-��۝ύ�yfy�k�v����'6���9��p���h��f��n�fñUUUU�U[�f�����:Jcۭ��
!�]u!օ|=��:I�-G��m�=�Gn� ��s�㮀�hх�;-�]l�]�`(AS��a��'\TjGr�=��9�Gy��^���<9˭OO��Ec>���a��=Q6v�]v�;B-ٍ��eW]�;a��c8�)g��@�e��2�����g���˻=	��&���[j.U��ю��rdr򆎌=�w����b�F(s�@�ۃ$u�<xn.=�$�<}	��V�v�cWh��ަ��d��i��y���4�2� ��ύ�u�'&71}�<;�����ˬ��Mڲjw�o��u\��:���Yᛵ��,iJ�Z�	c���q_z�w����{�����b(zz��چb-�nvf��i�e���*���`i�ۺ޳��ߜS�5x��;vD+���0k��W���J��U�����U���?5�$��$���L��:�M[>C�^�O�mC���;Hq��KT{�A�l���N}�}��׻rl<H	�X&�Z��s�ù�p��=u��.L��qV��]�������R�IV۞�k߷;��w/0\�噈���6�W��K[jn
�WUY���2�>�L�0�b������b����cV��e�9���qW�WY,Z��;5�g+oH�/x˳�*vu�'�(o�X��Jp�2�sǦ-��R��꩜�G^�5����~[�sM����tޟ�^Ǿ]4����\}���%K��$Jm ,���yWV$����W�*�˻2����I�{8��x��j���e�'��o�tc.2"�5ز�t�;%�V>�Ǐj�A^z+=�
�=:2�o�g�F��na7ה5ވ蒴'�JB2�^>7d�ͳ�d�\Ǉ\��E� �Q��#��3��^ӎ���M��P���������w��{��[��n۪8��<lhxn="p=l\ql<��k�U�W�l����.˞�u1��@<;��j̆���zf�-F��Vٔs�w7/�٢$��LH��Y�/n_z�N��Y�m��^nNL1� ������b��"�6�8�]O.�F&db��~'���f��xT;3O).��������%P|����	�R|F�C
��/����}�� ˄ou3]o��H�vN��K`Y�j_lt��1�\���M)�~�ӆ�]���g��ꕃs�F��i/�9$M�����f�U�\�;o��빼��"��Y�QhJ�;ʰ���l)7 PΡ�cņXa��Ʌ8��fQ���7�D�k�>�E�B��0w�o=^�%LL�}/�!��	����h/� ��U)y���&�@��E/n-�r]�N�(�IRH
FDp�0%$>�W��s�&��<�%��ǋ�����D9>��[7<f�"���2��vO��5E�Ƿ�9���E6:����_����0i[<T��/����WOOqg���-�=���v'��-�H�*�_ft��"u��s�zM�,��b��}<��Jy���Z��t��nQ�l���m9�\��Ew�}Gm �{|\�Y����㥜�z��}~F�U��������c�v|EB���]���F��&p�h��P˼��Ž�g����W����Y@>E������
{w}�'��I"�l��Y[�]�8�+L2p����e�O��e�W�%\��`k���[?v��ׯn��7�`�d�]�F��pvY�tp�b�vw&�1��ͭt���T��7'Mf;`�IlH`h�"�	��s{�=���h��s�w�W�_�h� ��N��i���լ�5Y(m�q
L�T�*P2���[u�~�я�P��{�~�(��iqݵݚ�do')Ԛ���/HL��m]{�A�E�SD)%��8ry�	��d��o+VƋ�����bD��mD^x.A�YS��b�{�I	���y����g%���ȯ�H�o�Yu���-�qt=/Sܿ����k���e@ʩQh�j�kӺڏ���:��v�{a��
:�m�{���蘛�.7>����zq|�Փ�݉��F�[�x�W65`�5B�v��7��'�tI��GZ�x8�{��e�|��/��Xz��L	�G�L��$Gr�ݪ��^ ��6�	-UUUUP�ض�;Z�(�ݛ&��fK��"��,�s�m��0�����n�\n2s��b�\�\&�q��:�-�.VP��s�
�U��d��:��س=�1�o]�Sp��`�n��U�k^Y�6�a��]�x���2�w�qgȏ�|��$�A��%�oC�q�x�;	���k��wa�5��:z�p����tgXwn��n�r�����h���QK��=�ĖeM>"�4I�Ӵ��罳;��o��p3�M�Ċ"�|�v�����#�����{��4�d�G������Y+��j�R��9�������Dyt���׷Stp�3��t�/�N�x���X���d�wǮ��)y�v�6s�㒢�殺�P�B�"��\�2sW=6淺c��0i�y�$4cQE�x+����3�i�}i&��d�Z��κ����q�J��,��IQ�1�+"�P�'�*��L�6�Ĺ+�j���1z�B=.x�w�p�����w�5��HZp���qn�4�2qр���]m�^��ԚMl!6R�nD�;��&�_����������2�	�8�9��~�4w��5��N�5ן:N9��G�#�/PUdFa��$��}�r�lŝ�\Yg���vN9a�R����WF
ܥ��B���׍�jSj�]��]Bz]�rahc3-�/t�3�]�V��r��\�*Gm�w��3ݳ���ߍ��>{��ٕ�MH3үz�E���	.܆/Q������6n-�����3u��<��˛f+na�7n�Q��i�X3�[^�DF8�Vz@xO�A������м��07�O{)��g:u���p�.J�Ff�4�q)$�L��q�YՇjY��=�/��*�o�U�_���edPG;�k�������]�l�n)�=��:H���)m�.����X�Ѹ��vw`�{��#���Rmi���j�>��lrS�x�{�O�.Ӻ���d>rKt��u�u$��J<3���{�8SbB�m9��v��zS�z�u�gݟ�+mꇴ�w���:�LL�9�q�{S�ff&X��fv�Sl+��v�f��]���nM��K���yMx���E���2�%��s��Tg���}��-�γqf�z�U,j�h��ͭ5n��h�D@w�Q�WV��HdUy��[���^�4�<�td�$-�y��3��gyfC�w�P�kk+C�JOU�ۚf�W��=F���"��R]>��/q4�:��UMV������ާ���o�	{S�S��̊˱񩸶�g�&�w�=zk ~4�tچ���Xz=B��^��x�����ބ� r@B; ��:�|{r|ֳڍ�z�]�Q9�ٺv��m��"UЫ5��^
d�ܝ���nf,���$=��|��t���a��_nZ$�����Y��o��k/6z�m�@��؄h���a>�S������.�#s-[΄�m�g+E3ȣҔ�1t	�o�󊠬�l��AC��[��QQ��C�*wt�wt���R�wpl��O�̒(��܋Ut��BHp�ӭN���BI���{x�I/V��h�A��c+(���L�0�㛦�,K7�VS�2�ٙv�Xֱj�8�!�*��]���@Z�;�"�q$콿i̭wH\���E�Y&d�8�M��Q�--<�]
쭱�(�5�M&H1:�Z����mIw��+�k�b���ֵ��fʠ�8Ki�mj����H�y��n�[�n�ю�WI�a�NN�z^��&��L�{�28b�wZ�mw��f�c=<�����N�	ܸS���a�O%e��y3�坻ɹ�c��|��My��"�2�c]%}J���Sȝ97߸��r�3Sp���&�~�g��헁;(��F!��$�o^w29��:���0���Z�o�a+�4t�����sy�9����p�\�,
̼��[cL%�}��}�>�{y��y����BC�7����G�K!m{6۸j�w%=U�s5�b�m��b2�u�%���W�hCӗ�I_U�4���.^\s׬4�@���W���m�W�y0o&U�]�EL"�v/�f����i�z��#�gyX�U�n�m���
��ټ�2�(/�gu��1������m��l�XIm-n,ys[MUUUUV���<{iv�<�8\qˈ'6G6�מbճ�����̼�O�࣋۳�'�2�r��B��]z��ctua[�v�2�����1��Qe7v�Y�eN�vΎ۶��a�^#�̧6�x#�On�>*��jF�zu�'u��ஹ�u�qn�\`K����^W,eݳd��Mvݶ�q�����*2��n�p���TpF�{���v�Y}k[u�vm��M՝c����68)�7	�~W��\�P�e��Ǳc؀[�<��(�yG.�����\�Z��C���Ye) nE���jı^ug*-����ҽ�nQup����	8t�Χ��r�<��0�J��}�U��VE݋��I�myoKn�1Hywq�n<P���B����~�6��+�W�U�`*B�h�Xpkw�ҮbyQ�M9|�x^�f(q��j��kv�"6��ʉZv�@t,�۾9�:���n��~^�&O���M}��c��1g�zC�^�Fn�rm�oX{ՙM�,��;��#���bF�����W`�$Z��8�N�ݕ�w3�����+`+�P�m��n9-�3��~��q��Vs!�]>�HȌ�5V��V�PT}��ު�W�kL�	3 ̕ ��J�;�Ь�p��ź�)�D�]��Ok�:��\��p�m�3�8K�l�[O/��BԦ����5���q����=����vd$%�h�0j�Ƿ~��b'���>�c���p��I�j��W����֡�a�Dd4T��(��6�n��s�y��gAz��s��brG�|o��u/��Qt�1��O��/�ƛ-����M{.���B�U�
��fy���O�MX]C����*��v�
��m���k��D�#isJf?����ҧQ,(J;d���A�XF�bA�7�\æ�=�,�;A�|�B}��ԣB�c��F�J�ľ��t�<�..�}+㧒��4�
�"�|_m�����
�!�&��ӵ�T��q�����FJ��t�G�=��c=��U���'�#�k�/�҆��� �C�NߦJ�A���D�c�ϾT#�����X㫠,�ӌՑ�E/��[K�"5���2Q�FÂAC����dY��Ei��{���{����7hyW9�B8YdIҏ
��˶x�0��5k�9�M����<]Ͻ�F0��k�p�4Ih����m>�F����?<�����������޽�e���>&�C���G���`�_<��;�Z܁j+�W`೗-�G��^�v�ٮa�ڪ��:��3_B@�������1%-�e�Ѹq@�]̿�M�õ+Ms۴*72��b�,CĂ�Q@\����t��x1:W:�����\�[�a��,�h!1��u�NC�4����T�X�gm�=A��#�6\�Y�ji�V��cV�{dbP�}���+�Vj��A��ï#]]�1��B ���\��f7n�)@Mل7с�����ׂ��"����WَK��k:�)ܳLdY�rb��H��bm����ӣ�����5nU��)V(�և�d��j��QeԢJ�ݷ���Ɗ
�_aw{ m
]��P�����Q
C�ຆL�!!�9ܣ|��������j��wa]W9)�ff����
�O9g�ۆ�2!ϹS�J��ݣy�V�md�_�l���T�7ޥ܍,�W�����
w{�:XǺ�d�9[�76��{;YT��Y!c�;�U��=y,�����s����,⛛�e��{\)�⨙h��&��&Ң=7I��)X{n]���M��K8��7�Dۛ�O��KxCWCgj�bk"[fV�fˉ{b�x�ʐc`dZ:��M-�G�?a[V��(��#C����a��g3c#���8jl9�^sUR^6��guncύ^��v�kK{���*��2�e�n��������-7�1�8ӵٹp�ߚy����TCHR��S��ւ:Fi������E��8YPC19%:E��w��$Q�VGxV[V8�~�Y�d�O�Uc5s"Y]6'�O�rȇ�B�}�tS�ʗ�����Rp�	�%��}���_��܆���U�C"ș����*�o$a�}�����I�s�[�j�~*/��;s�Aj�dI�8uW�z�,���z֟�{m�߽�j��PV
��yJ��q��-:�Ii��\��n���ۅ�nwn;/Hp�qND����i*(;�J柭f.F�GJz_�P�q��t�iz/ƄA���^2�G�?�ξ��K�6���h���
~M���a*�و|}�o�5���]�z�3�Fn�F������|�3#�#�6�DUeyXˌ��H�&͑~�zjHm	w��T;���ߘ��#�E�x޲�h�n*�z�6F�����,�i|ȣ�lD�b���#�=�3�D��5| {�\��22B�~��$p�AJ~����!��U���tEp�[!�s��j�s��{�Uպ=�x�{j�t� ����w�鿺i@�����VO�x�_e��%b[w�a�ٺ����_N�]FE�\s���V�U�����Y�.��mr�5�K9�k�:��&�a;7��EAn�sH�_z�j�=�X8ڌ��ڄ�!���j�Ȅvg�G\�Q��q�ɤ�VwH����Ю�>����H�77�&����"��%}r�<Y2En;!`���4�����drHv]ŘGul%����up�Ssl��Î3Of;�TX�U5�hdG?������2M��s��cO�p֯��޷�c�g
=uF����6#��c��`n{�`:Y�HU��[ނx�`�Ha@����qhFIf@[NKBńi����V,ׇ�8���YYSBg!�&񨦾f�׳VG	���ѝ���o�n�����'��F�O��4�
9.X�%�� �ᯈԅ-�,�>��a�δ(����s�+���_��(��uW}�#�x"n)����_�2<�2;���۪c�6���mC~��3I��#A���͌�8�˿]h��Ez��`�l�"��f��>��*��4���:k<h t�,�"�iC��^<vt?��f�P��:�mυ�t"�R7D�ǚGIZ~��DkM�}��Y��/�O~�T{|��|w Q�/�G�Bj:s�$5��Y&#W��M�!��>:E���ę�f�G�aȻ�e�N�g"�B��Ꮧ6��ĐtҾ��̍ޗ«�N��.ZyF����:�2b_��~�߿�������s�*������*�UV�tm�n[���{]��;�u�T��X6����V�����n'gN:�u�n��v-�s���sz瓛�m�}Y�!��m�Cn6�q�vK���q��ϱ�OS�=-��z�v|qzC��n9,v���y۱��;gW���y�:���u�ȣ��;����{v��zz��`�n�6�n8��1�J9��c��oj]-&(����]�3G�v�'Fu�s�q�v�uĦ}���6p_�")mj��[���\k����A"�;�CK"���20�0MzE��G���8��)�Ƞ�oEL�!�������ʫ���=&�G�C�2�{	)� fA��g�燾B�y�w�A��oհY	yB���~�j:��i�/�վ�a5�r�J���p��;U�",0�Zȣ���.�'���R)T�����N�֖;��ϰ�?{��je��ɑg����q��A�G��~T���򆈳��b���F�B7�ǘE���R8A�G%��p_�~��D�9I
�g~\��W["H}Y�_sA�F�#iC��B=��L��"j��}d��]�)��X�g�a����Obp&�%��0i_�t�� �xWe,�Lp�N�6�A3���Q���tuj��a8����}�顠�
��{�g���f�p�jd�"o}�oҮ�����f���۵����z��S���;�-�	�'<�n�����n�Q%���h���ؓ�#�X�41{"��Y~������8�,Ѳ��頽zq|�w���ޭ�Ȃ����zG��=Y\�y�����QPF�,&$qP��#j>XD��=7�*c�_���2���"�BVP�ᵯ���H��g�L+��Z�;��/�lIffZ�&g_R^Q�ûW�C%��+(ge���F��<DB<b���z�
|?A���h��~�|o�i�#M�>�	�AAt��տ���� ��e����m���<@�ŝU{.��Ȣ7�����_ʺF{=(���ƥD���m���mP��rD�(�����GP_6��_g Z,�1aB���>#	#Nk�^�Sn���y��?�|O�T�g���C��e-Ԉ�Bq���dYr�"}#8ff��?d՞<I�D�D���*����e�"�i�<���O'ݾ��z��0��
�~/��۝�?vW,�x�>�Q��Cq}��4��~5����<�F�#�i��?y�$	����3�<]��ns�u��!��6�]���Y0��q<�+�Wie�ʎ��V��;��kw��(�_~�뙫��"��&���J���:d�A��U�,遮N���$���?8Ǌ�-!�2��>��
�$-2����A����0�����M�%tس�E��-��mQ�!�G�"�}��a^�с#�bs��9:c�h_��v}WDI�i�5��H�a�2ܖ,��\T�O}���i����F̑W~�P�/��g�y�]���~X��/�}к�0�M��E�Ֆ3�V7�Z���v�V�ť�"�.�]�v�yۻ���I���4�~���+���h:�YDw&|�+�ب3����)L�G��|$L8IA	1�_t�Vy�
���٫|`��ư�(�?Y�Ssފ�AY�\E����CH�diwI�ޚ�^���H��P�#qq�!����e%#!	q^��x�q�"�o˿K�ↈ��X�o�>�*#�Q>T#�>�ǈ�:FUg���6\���u�u���?P�0�8�Cn:���۫m�2QƤ����&�`��������s퇯@�iø��P�!���mZ`�((�����g��:�!��v��a�}��z2��A��dy�=�c�\P5�|D���<`W6���!O�	��7��+���ΚŇ��ӟ8	ațPģrh2;���F1޶����ẽ~󇶾���=�E�7e�����nǽ�_2/���߫��|W�}y�>�yy��������xA(�!Q�m��Z�5�0d�в.mʺ�����!�mJs��9�~���������Y[�0��\�4 Z������������g.�W��`����oNڢ4����FC�фU���Ӝ��mi�H���+ɑfz#��A��� �����c�R�7�z��]YT��ۣ���'>ޤ�#�Z\V�v�?(�k��V_D��-*3*桓��{�[N̵ֺQ]��56����Zɐ��@Ftj�]n@��y�&��ض����~4��㧍��N��olÛ5ă�Q�ܑk��4�l���B�������ޟ�6�"�~��8�=��9J�d�cXa��}h)R�8E�v�v����,��&q�Q�/�5}"�M��#H��fCY�#m}܅�V@1W��_<XY��~��b�7l�~d3�}ym��hB�,g�G�[lf)�H��p�e"9W�]h���_�tĞ1K�.};��뀵|�7u�'��#1��[�H�:Ge8�8�_|5�y}����>�äB_4�::M��	4���,ܡ�A�	�G� �t˾2"���Mp�g8�;/�֑≤�`�>^�Zb�?IåDP��E�� H�	pH�i}X{�A��O��WfY��o���;�Y��S_#-{7#�B�?q�y���5Xo�l�B�.H�f\���i�Q���1���b0�IÝ><�<pѲ7���cI��fH�B��z;����\=cO(���̴}�:p�=��H�^����!���=�X�􏬋��KiҞ�|0<O~��
�f�ˠ>�ODn�<lMJ�6��v��{p�՘�WBK7o���F`�9�ܮ�E��]G�$�I$ψ$��.E������p8�ܴ��"��ϲ&۫r��.u�R{'����j�s�v�ݡƴ�i��M��{#)�9�&*����7d�/	����9��=�8\�O�Guvy���٦����]YMsm̓s�V۞n1�m����m�m�v���m�;9���r�
��=nz�2npvk����ι�<�z{M��c����RdnSGNU���v+<��]�[��z�[\���`�Wa��C��|�n\*4����ߘ��{��[MzߵP�tbA��é^u�k�Г�I"�ދ���Ylj[����%�$O�|kHޤ}X�$�,4y���n�0LI�3
����:����x�;}��QzG�fr��͞#���"g���F�X�udyW��}0h�Ҥ��a�$���T���}�6�)>5ռl�݌#�Z+�H�1e9+�>4y���9���#G(.��5��(�_F�pg�
-�<�n	k�U�Cs}>��ӧ��B�o�dm��cKSRJkI�X����z`DMunG�q:p��*6~��x���K�(WW�4<ZB�RG=ϡo���v�wW(CHmY�c����$A#$�sϟ�s�i���p���$=\FJB����3�}��#�a��a��=�B�N4�m!*�i~�`�,��@�G������	CQ�;f:zvÚ�7�l�r>8zr;	ֳ���\�[=�/\nD��4��ź{�EҼCO�Fiuޛ��՟��iӞ����ܾz���̟OY�#O�FZ�^�P���E$N�`�/�#�-�qJ;If�����v*�3=�b��~�=�C�n�mF�lI�Ka��s[0�j'82������-�.�a�E|rY��/��I�%+����ѧ��7s����xY	����#��ۡ���/����ӄaF�4o�ޚ�G�%_ ,N��o��F�_z-m��\r�!)��s�� 5�3O�^�w��֬�G��f���i8��������%�=3s�Y���{Uۡ��o�`���gݱ��)=mۄ�$�2laf�#�t�*
���~��f�!(�񏮓7ٞ����G�E��sʃ�0����DV{�!�5dixȇ����%���J"a�����C��,���E|�b'�Q�k��c��Wm\P��$�6��YU��4C!�G��[���4��P�]��CƄ�UuI�[��y�瓐�)̝fc�Z�k�����n �b�v�o/�ƴ�|�q����_�~��h��_�����·��-��F_�oƬ�hY	�EZ9=�;��Țy���M��Ld��_i
�V�$�0���`�����;�ܒ8�|�G�ǐ�8�M�}طƾ�.,1~�f|���՚3�2����(���	�{�Cҙ~g��u�4�����w�Q�P[i�8����Ğ��`"���4�<�]8E�zӖ�H�����A"Λ6����sq,3mMe���Q:$Z�8�!� ���;�;�u'3�	�V�&�Z.�(i��N%��9��y�M��4�C*+��.���>"���Y�W�i��,�8��6ֆ��nˍL���"�����TU3��D]u��I�Z��k��D{|�il�<�$����h�="=_��=�vpͼ�� ��@�.�k�8_J�R*8"��4�#��B��_:ç)	hK��jD��D�C���o��3$Q����B�c�B`ip������k�<p��������x�`�a1§$N�MN�U@*���=�=��;Q�� /I�����QI%�_�zk����^���s�;"y
$��i�A���&-�d�&m��b�j�@�!�;Ѓ?x��/���)����A�Ν7��Z��b!$d���{�M|�$Z��ѡ��e|������t��$�C�wM|��@�$Q�H+��Pӄ�W��	����z�Ǟ�Q������O�����JE��jF�iʈ�,��3�<�I?b���#�����ɫ(�I���ä�?e��/�"Σ�t�e"$�|j8I��urt_~G�"�r[
[��Ӏ��P�j�"�F$���гi��ȃ�V�n�;�c4E��z��
.+��'��~[�%VO���1j�M5,٣(H����w�&�]3nV��}/6�6*���P��)�ބ�k�:E��օC9a���+�#+����G
@�$4㱤]#�S�'��;~W�"��У�|�eU��n��>YG,���J��|C#O��~��:`������T9�Yk���M6�ôq�����F�-���҇Drmun�d��թ�J�r�p�����h��Lp�da��<՜<�+q����Y������~A:���#�ܨ�Ci��9s�s)�w�H2(�%�dw������E�N��Q::�%zA4F����s5��HS}Dm�G�. ْ�qXYٳ��:{|h��+�
����X��Z���e��z��#�P�G���a��H�o<�e�N.<�|�gV��h���y���C��CH+W�o�Jc׋!o4<hc����#g�ɣŔf��\VM���W{[lQK��Jb�U�[m_��w�pX�++׆����H#�?Oz�!Xt�HĤ��m@���г�a��,z�#y�d6�b���bDb�2r�P�F
��,��`��0�#��z|rƜ�0�r��9~�ppؓu����BO̊4C��T0�U0�t�3��C#־�,����?e�r���eY���!�Q�z���6��&���y��f�{����dۇja�j0g��"��S7�:��I�#��T�v��o�r�&�`����Q����}37'ff٭wѮ����7���*𑰆k8�gI{�u^m�\!��d+*��*�ecl^5�8ⱺ���s��Tv�k"�FU�mT�Tgl��#J���ں��& ��M�[;@�Y�.�:�.�;9�6�R2��P��P�1{��f��l,
e�X�vgW9�E���ŧ#�{��\.S���5{:���+��!�co����浕�kS��2Nyys���h4څN�}{���9S��S�o^� ��M�[����ϡ4'm=�m'O�NЭb���t���ׯU��j[��'�x_��k��;WkN�n3o�z��l��(p�ɚ�Vιco5�yd�.�U0E��T��h8A=��a�p�s��p���������5/p9���mȖH�K5�arբ��Э�Hi�b'�k=$6�]�a�ھ����);�I��3��jTRѵ7XP�>����h�*S�o�r*���wK��}�3%��\.�;�n�3�,��� a.r҄�P�m�[G0I�S��ev�y$������Z��n+���E	ǆ�B�&�ϕ�Wn7�^���h�n��zRl޴��*F�ԡW�8�i�)#K�xk)ޅ��RH��u�G8'Ǹm�$�I$�I$�I5UUUUUUUUUUR�[Rb)UVM�J��UUUT�UT�l�CԵ��ֲ���aYZ������������������������������"�M�g���uH������ZT2l%�^r8^q'�X��1�����0W' B��=���x�{un[ �t���ݻ��>v1Ѷn�q����ݸS��Ȏ�=ax�b�-�Ý�#��9՞Zm�u�^V14�n{C�<)Ȇ��B]��d�G��ۣ�y�ȏP���CJNzg= G8��=���;�uCpnm�TErn���\��<z"�4g���n���ۨ9�$�]��yH��1<��O`'m���F:�qv��x��]3g�^�AˋEV*�mwl�y�I�qw<:�}k���΃�ʡ+��x�q���n[�{V��񞳄,ܙ��Ot��"��U[\���9Z��%�u�
S���5�ݭm�N��b7mԧ)�j� =�p��s�u�byܜ8{7�f�ݭ���]7^�1 �e�<�b|!�9i8{v����c"�cP��[�tm�� Snnfv	���-�|We�]��#�ln�cq(�B{�����ƈt�y=a�������3v�zڸz�����=��r���<���9ɫ��8T��K�ݴ��훎�B:��6��,#K<���ە'�����g{`��Zx8e�筮Ƕ�U���@u�n^,j݇��x�m��E˻����i��8F�ͱ��m�����9P�& YP�޺�$=�ԣ7�kgw]Oa��*����0sq��qq���+[=�:��'��m�'lo\/k���=��<��n���Juc�Wl���������ln=�lvsnN;&2�<Ku��,0��{v�%xR9�q���x獩a��رhqlz7�%@��v�;:�SsŚ�i
���5*�X\q�k�����trq���z�1^�:�7<hx;�'�v
�N�v���k���q\q�q���躢7PT��h�T00ؓh����kp[�]t'�ʎ����͆���cE��N{�UUUUV��^;)�ݱ�
��O:P�.}��g��\.�K�O������Nz�1���i]LS�..��7���˷.��iD_n;u�Q�N�a�;z2��n�'��
B��Km�:��jg�9�W�W�RI��&���{;kc����"\=9��`�c7tY6�+�u6@kp ��N.���j����2���<g����b�bvM��Jټ+�e��81NV�m�z�u��Ƚ�g<�)�`��?���k�i>�5�zO�������fNw~q@��g���W����� �w����/��
k a�>9U�Y�G�0��:^!��!�[L)��.I\��P�R�x��ߍ�0��F�����#z>�5��ӽ��h�m"3��?��P�_N�Z����M������M`�V7���_~kS�%"����c0��#�#̯�W�$���ɵk`]��֖~�9��� r�Mx�O��^n�x�4C#Ց�L����;CM6E��"P�6��@SR��'��Y ؓ��صP�TE'W�[p��_8Α�{�7�qdc�ء6��$�XQ1�Q}N�H���s�z|�Ӈ�cI�~DfI!q����6GOAЯ����2~dQYU�M�f��ͯ��VF�O�|hF�0ȓia}��V���<o2���=Z���tU��@�oTJ�ug���lp�G`��۶ˣ�i�/7E��쐝=��ru���.��������y"��_�:G�Pg�֟��:嵧Ő6A��b�c�$Cq�頼h��/{�k~!��T�Y���

	I�2a��ێ��H�,#M�C�}����z�Cqk>���
���d�U|ȶ�]�[Dt#]J��?���H�V�yZ2�ቛ&�SN�����B,l���N���h�A�%x6+�(*��E0x�&����ف;�[��
1��^�آY�_�هpǙ�b���E��n��(<���m(ԓ9ӭa���l���A������M��{vk�D�珅�ӛ���}s�A��A�v�y,vk��v�0<V|i���$*6$51CH�Di��͟D�����xx��V�������(����΅2�r��Y<�P�n/9����:ꕈ�Tw>����_��C����=v��X2"����L<N���4<��|��M�g���*W�V�7�vF�D3�(��a<�c��"3PÄE�z+�YcP��?r�i�Y1;N��x�B����}V�|^�����{X�Rp�Am�=.[�OF��m���"��QG���҄:E�}�X����40�Da�qx��l�ϙ��}�U�"�b�n�,�E(���� ��h!���xA�C�$
5F8k�w��~c��{��1�>в*��_,�NU�MB�ώ���P�ɨ�M�و0��H�}G}7d�F#����]¢��8�.<�PE_�e�>(A�DᡧK����>8Eǽs_i���D�@W血��>�Ig���e�eƐ�kk���m��E�ܣ	�*�}�.�����M��L�`�YA���X�ܘS��q۫�s.1�V�7���Bv��}؅������V*b��4հő��	����%�0���,�\�矠�����s/]1�G��:s�>�V�҉�7#�j�{|kM�������GI��?�-�^��C�`���� �$H��"�c/K?+A��E$=��*�e�E����dQ2k-{ȥ�����S��!e{"�"�Ǆd�_v^z6�?f(t��,x��/4/wbܐ�Y��ov�ؼ�`ɍ[x�tt��9J��6Î���6�Clb�:���*�U�������D�~40�-0FU��^Rsʲ�[7��6��h(RG]碅௺��w���A�����Eq��q��OѴ�G`��r8��
X鋭N�k�cS=��ϸ\��,kL����)~ٜ�мC�GB�.�w���$a�4���D�o�S�b
$��������ǽ<0��g�o�0�Ƃ:2ۋM���?�-=8w�|����#L�D��Y�_h"N��Gc�[q�ϵZ����8��F�Q~���Pe����/�a��,�I��Tjr!����2Pe�f�(��w�H��ǜ�̛�G������Ƭޯ��ȭ_a���:�T��Ar'_�~�8~ߤ^���tʍ�:]:�V�ݝ�EǢ�/`��h7�z�L�{a0�ņ&�nΪ��c*'����������dAx�]��_4�e�|�$BSr�>ߞ��٢��Q��MPx��_Q�r�֊ʚ�����ŝ	�W̋?M�_�ǚ�o 2�!;�*�"�iA����?���|d_��a�enZ����5K����F�m�K<=+mer��x����`n�7#�t�)�Ǽ���(y#�[ɱ��4~M
��U�(>���A~06�Y�aT�۬O:=�������s�T�����p�4��Y�V���i1b)sON�D�^�E+csEE,:9eK���?i
�_���C�ȳ~q�6�Uk��7�{f��C�]턶�^}�W�����~N�\���:K4�׻$Ы�j	���вώCPl���"��_Q>pnU�8���	�,��K+�t��
���������	��0&bƖ���~w*}�
<|�?e����Rp�n$�#:��dQ��?{r�+Ƅ8��	�
��\:o��/H�et�0���閹pz�[-(�0�Q�� 0�,���]����Xx�v2�
��y6��s��C�<�س�����H=��E<F!�6~s��U	�����a�ݗp���^�n���W���h��o��F-�� ��U�˫A=,���U��b��:a�(����x�n��]���t��d�I$�G�������e������NN��LU;Q�(�k"bg�Ϣ��s8�}m�5�e��ݸ��	�r픺�[�v;c�;�m��>-,�8E�����X[����GP��s��'��=Ţ��
����0�1��<\6�Ⱥ���N�����g!���l��2�7qǓ\���ܫ��W[(HaÔ���y��{;c&ө�g�������0�&�ݎλI1�^6^ή�wV�y#�7'��u�������x�V ���vy�\��ğ���ϾB��s]6Ez���w����螡g���i�C�ڶ(E�L0��{��8���Z%���\��#�d�z�2�H���8L*IC�����B��I�z,agFj2�ܟ��t��T5����"�@W��6<Y��z"��9���������8F��z,�zp��^��
����
E�n�/gZ"TcHd����ä�=h�0��z+H�!��E⇃ԫ|G��9Y4'�v��N��W�d,_i����t�>أ%��/��~��t�}����hQz7�o=�_{��N�G�O��@���6t�1\��ǩ"-����gC��+ϣ�?H�F�~�&<A�{�D��L�"��,����hQ�v�{>t:k�R�N��E����e�}��"�9�"�7ʅ����8�޻�x���~�ʵ�O+�_gMQs��)""�֞�P	�mupE�״s����v:I��u��u��ȣq"���ƥY����7	����o���H�G�sg@��V�WQ~�B+��a����J�Mg:#ؾ�8���Q�4��I�0Q��"w֏b�����u[4������Ǧ>7Y>T4�a�4z�y䫕[7P�hl��_�k\�@Z��ef�Q��������ȸ�3e�ը5W���2�,�L^��%
&ع�/\�Gu��>U��oM}��x�B�y3hVDߢ���v`{<���w����H?m�u�-`̮߰+�#X�yڎD*A[Jiq�ƶx����_;�~$�P��A�}n��"%z7����b����6�UX�]��X����/�s�Yq���!�/ɑ���A��2(����\}c��Sй���ӤSS�;豦�!X����=�*��3g�E�p{�5X����6=u�1��/}�v�zGo}�äy�JI!�!�PI#��x�:IE������z}4��-�ݐ�aY��P���4��E�|懏g�g��.����ֿ:�Z���ݧ�y��I�u��8� ���4JH��LKv�Md봧B�Bzp]�sb�l����v�a�������8R��I��T�i$A포�1����g���,�����a��pA�#�g���0�<DWx��,�����?P�Mg�&2SN(#q�CH�+#M��I��J�����"Z͓��(� �^T"�>�gԑ&�����<h�������vʥϦζF�͙�j�c��d`��F< �[e��18�~G�HG���i}�7cO�`ߜ}��yڨ���1
��ᐻ��&�P+pϋ�5�u:/\�)���nլ��p=�V�s'��2�Yh�f��8R�y��C���<<#V]�f��k�M�Ua:�"�Aj1Α[�M��g�h�ȡ��TH�JI��M�CH��3Q�
߾`�)�B�o�Y'�4~�B���璨3��Y��U�说�0F3RW�f���k���g8x�{�U+zydl8Fw�����SL˕�t�V�w'J�}�O,����eA�X=����Ýw�荟@�$�c���*쏮P�_Y��V��C�>g�y�?]g��������Ԍ|TyT��ۊ�v��]���㵸���m���h����>������sE�y!=2{�����[���0jm{�_i��i���SH�Mߢ�5�5}r�yК��P��,�Y�5ފ�t���eB{����f��d0�e9+�Y������}��P�<��xho{z���1�{�w�U��TDg>�6A��4:�j�ńWm�x��ל�@�����;�:zy�k��@� 0�8L)�CH�*Ζye����}W�t�,���12�d��C��'ެ��|G��R>͚ҹxɳ���^TA����$1臭a�fD�p�J�7��=$ZlB5�dT0�!
��K���xx-:D�ȳ�D�z�4+P�~PY��wY� ��Mא;.��kn�/KYW�2�Z����<�xnY���T�v'�9v1�'��N��Okya��?m/�W4��\��Vx��5!��FP�$t0�6Gڥ��}��3�s:�dz�F��I�M{�ΉX�P�#��V|D#ޭ�;˥�4!��Gu�ʡǎc$���s,�<Iz��2)
&[:\�����6s�(��P��狱��@���vN{���=
�Y�������:�t:(�f�n�x�##z~�It��E}�3�IdY�.{�B�0��WU��YE������4�:rT�D]�rҤ���`��<�i�(����k�{�|�ܫG�g�g��o%P����� �!��΁�zF��)��(�]�*��N�Tp��t���K(��6�Rg�J!��-����O�wv����~�1iݠH]���J�W��g�6Ej���a�;}�߈g�m�*ӗAE�(�1�(��~4H�F��4����#�BQ

�E$V,�iCM��%[�ҧ���������F�F�Y���:6h�z2�=��8x�#�J|�G�3�|���.�-��<�7�)�~j0�m�b2ItF�<�0�<ӫ�Pӗ�aW�kN�$|���^^����{z}}�/ݲ�>_U�h#�Fy�+6�q�ޮCG��)�M�ם��w/�q��#e�q��۾/���o=S�&l�u�(�f�̘��`�'���b�u s�(f��g��w�I$�&XdȔ(��Ϊ������띭ֻ�����8���{y�=i5���vW�7\�Vfs�nN��۬qƫ��b���<#�ӹܩ���+mٻ[�
�Og]������f�����8W��gnm\��C�Ɨ�秋K�هm5�λ�zW�^�u�8-^]N3v	dL�ywY�<�1m�ɻ�<��q���;�F{T�k�s�nQ�읇^t�y�Ý��{�N��)s@��.�n�gT<�V8]u���`l5��m�kDI���?h!�YF��~��x�	��00�H��_��0��gi$\��g��_<32a<t��0J�O���L�p���]j��G��\D`5>ܣj�Bd�e�?u�8ԃ퇲�3����ו�)����1*s�⬒��	dQ�l}u�B7����z+}�!�T<%tu�R��󺍯* i'7
n#�Gb�-B7PF�ј~Ͼ��<{���#����x��=��6��5������c�-hY���G>�܊����n!��<~C��&2�P��R;爳�kJ��d�9Gӊ�f�4G�GM�ݟ�u�igbh����аy/jF�(�|���SٓXA!Rdi�G�<��J�dJ p��w���R81"������p����G�3?H��
�zU���8�D*��W٨a�P�Ǖ�:�t�ZyGK� ����m7�v=����v:r�1�����s�	�{#h{=��^�0&�P��-O�[��O�E�f��E0{�v
�
J�ޚ�=�H�]�i�nd_��Ōw�Q�'ky����0��oƼ!��!C�b��(K酸�1�$q9 �Fm!�oދ�Z嵭V��{�	;��l��)��մ7��H��4-P��jТl�xh��:>(�YG��?���1�/���2��b(�z�ձs{���^��I�ءCW�q�C9�D�Nz,P,��8�4Ge_��R��_���$B�J4aY���?tuҪ�ʣ��}�קƻ�v�'��z�DX��f���k�����Ջ�c��H����y*�?IDR������v���ѫ�#1sז����8�bfhf��������5��k:Q����g�r�"��`��z(Rn~�w!��zﳮn�0��3n5CP�k�������.Q���A���]�y&��YF꣄�k�mi�w�����J�%�I�4K_a��1��}
�c���\�<1��,��W=�S�r����Bx}�8Y	�0 ���D]��SQr9�Z�ݖ�_��^<3�q�m���FPk�ŕ�����ڴ�6���n��h��"�@<����y��N|�5g�E�G���Cs_�f�^�g����r<~�m���>5t�|�{*�#s L�Ma�=V_NB�%1lEudi�����#a��{f�3{�����h��4 ���Z�M٣�=~�h�>!����0�X���]���"�#ꐂG��p�߻��T��6j�3�D���f�(�(����/�sU���Ҏ�
�8�VK_I �cxЕ}��FU���y������c�/����OAt޾���Óo9�@>����6.�3��x��7X�wV�#��F�\i����)c����뻛k�;!F��ֹ��v�x���1T3���r�ma�\�&b*N��/f0���o6r*7jӷց��dE��2�w�o3]���^�5P�j&��!����bd��k
9�m��#�Y0������ɏ��1�y��ih�˛��:PN�R��f���ZSLU��5����76�^����ƈ��o	$�Ǘ-<]U�Գ7ǻ~�8��㬣��+��b�H60���P��}�s&t���0���Q�za���r���DtN���[��&��S@�0܆��;>՛�mК�H���3%Q�� �I��vv;���]��P�Z��)y2��wr�X��3����؞v��Lȶ�9��Wt�V�Q��GKRY�uc9|���;x��E؛b�[RuD�'`���z�j6�����9;��U��B�R��.O��J��ً�
�S���̽�<8���q=�<3h�55~|r\B.�xD ��r��=,�:�K3�Q8�n'�Wcv}Uykv�O�`�S|�B�=sD�N��ZviR����[�M�gy5��i!����$F�w*�.�� �x:V�9����-�V�ܤyxJ��7e�V�ڹ!&��ԗ���@]�wj�'�q����c�U����Sj�7�C8&	U:��@����z�}���57���,��!v�.W�U,ȏ ����h��_��lb"�1	Q1�qÄis�x�����kY<��7��R4�����ճ_=!��#
dxj��8Ί�G�C<f�x���5wF�^]�1��P|ZB�W�a�O��*�Q��F9qP��}���,������ui����L)�n6�p7ҷp0k=�B�}f����V�诽�!�mh(Y^�U4H�� J��rz!m�ނ�1�f�Z^�/�\t��4o>��gۧ�n�=2s����Y:�kx}����k���%�=�ܼ�j(3@�#ڃ1��cB��{��>���UD�lG-�ADyYU��H��j`��'��B̄G"2�:yd=[��z��;��Y�m���}�����dOF�(V���M�De���zhY$Q`�B�����(�F���5���q���=��"=�>ɢCdh�
jC��Vyԅ���j��H���ً��K�4ɚ=Q��,鳀�n��Vp�mCQ�u�ߝv!�'�8�6yY/6�(-�`�G|t�m uLcz{S�Rj���0ff�o��Α�#��}�Zz�>���}����a�<C#����r�'��s0�١�e�~ݾ��'�q�VN	-S�O0'.�#	�973�9q6@2.	���*�B��wYR��w�����0�5��B�|Ȳ�$ciF��#GW�E�lȾ��g��Z�A�=��=��z�z.ȶ}~�&�#I�@n�ۏ�����_��k�Y6�p8�����\��HyBW����M�����}���-�MKkp�uX�w:��]6�no��$ ���r?a��X=٤3ʹ?v�xP��<��h����U�����x�؛��P���wYO+�G#H�t}������k�s網k��n�	GS�L�G����t��,گ�t4��'��`�����������&�<`�)^�EY����nd��0\��V�-"z+|��@����Y�ϯ4/N5p$a@b��a�-Q��D��W��X~�.Q/���	�"��� �<�W�K�8���&V���H�;M��UϾyd<���'�C�x}�ِ�"m��h�%su8��v�G��|�N��GN���V~(�$f�"������B�1�:F�=�Q�Vz�Q�,�A��nP�\=A%�G�wuN�д>t���i���^�Bb���K�,nȚ��d1/���f��(�~��b�tDsؠ쯬���j����憏.#�B�̿dQ:~�.�гt{�=�<��B
�ʄ-9��ˮ�X�W&UŁ3�Ε1���,K�������+�E�vX��-:,������n�I$��RI5mPr������kyƃ������v�s�9I�:��=[3�c���.�=OW<jEwef�6�箫�v
�N����Z�W��Z�;����1���7�����ŬC��t[��ۥ���*�#u�7;��8j��9^�qw��cZ�ud[�q�;�\�A)�7e��޶�.�.�.b���Jk�����={f9�<���V�:+;Evd2�Nݵ��ۜ¼h�����'��{d�y;\��<Z����<"-H>�6y�y>���y�!�W,�sފ�CHQ��<E�_���4���9k�m��Ё<�Z�M+�=�#�RPï���_��KZ)ڪ��[|}za�z2F�����
<o��̜�Wy'�Nbx��^�h0hᆾ�(t��C-20�A�˽�j����YIO�s�{#@~?�D!p�{���[1��jG|��N����;�=ʊo"�N(���P������^}���$�B�s�B�����J5��nw��p��?3&�G'�y9]`����,��������K��1@�X�^ۆ0x����n�8G��{��h����Y=豞[�3Dq#��i����ߡ��W?Iha�&p�|`���h�FG\��,<��|lۋ�PfȲ�4ٟ�vF�<d�z��W[��e���A�5�B�'��mn9�۸	
yF���b��Ȳ0��zt�*t�j�)_귨:2�$�V%
XUH���t����Yb��b�R,��뫊:��!�-l�3*bSЬVEr�0���k���'��?w!��Nz�(\d}DI��1�}���y[��DA�g�R�Rk�V�m~dv���0�ѠJ�
NK��.�z!�a���Pӳ �<t\7錚U�,�h��0�:�ʽ�D��l�.vh�rfuL���I�l�U��n���1�0�B��4�n�gg_xFǠ#��6�����#H���Ū(l}I"�\��ʯzg�i���ּ�0��|sv�!U������8t��Y�U�{�����,Ơ�q�l�Y^Ȱ���o��r,�P��}�Gz��c�m�qs�&Ѓ�������@���/�a4�Ʉ�H������;޺�Z5��S��w&M�|����љ�u�<�����߫�B�3k�JU�t?z|#l�~9q_q�?oL��1"
��|>m�E�ab911�YKe��&�������Rp�#�nﲆ��t&�	�1t�#��}�a,�:h���YE��}��j9x��-��!ȁ��B�v�f��E2;���%,��p�u�Q'Gp��
�Pv��{E�5Zζ�qָ�8Ī�?����}�!d!�"+�Zt�(�?Q
�w�����da�h��z*�n}ǝj�2��h��@�L�ۯE{�ƚ���'��,N@*���Kf-�>'������K0��A3'�����$��;>�-2,�~�p���(�4��t��뎯MZ���~� ͕�\���~4B��&r���9if��E��]�j�Y#з=QA� ��}G�#/�sC����CˡDzg��/��T�nS����u�V˘,�z��޺����3���َu�GF�_�]�x�ɴ������'���G���'�x�t�4!,"{kC�X<�irU�ak��$	0a)�zN ���J�-��k6F鮾����@�i��Ҵ��J�g(��6Q��^�,�Ҽ�m�;fǥ�~�8���#��m��C!aa
��D$fL��%5��p�8D�"����:��O	Hk~�}B�|�8|~8a�;���\��P��W���D�(���řYt�>�O��'
��E>��7��r�N҅N`�Ƹ۪']�.��b�7Ud�T�U��8�-�\kk�>�"$_q�_���ȟX����8�w��v�d�}Y �g��6|��s6��_x��sת�8D��`7H�]�ԤbH#"�y��XQw�8p�~Tw23�zOy�Ƒ���:Ln����:�#W:F�@�߲P���[Bg8k����������"̝?(�dL���q��TF��~Gھ�/�g�:G�CZϭV�p�47+r�'��V{E��2t�P8��_@��΋ÝA�8l���ԾahE ��*T��ͭ��~ꏋ��}�d�y��ߦ�1#��ؚ�7��>��#L���Eh�_��-E��=>�����?���QO�$�*1���O*��d� ��x1�b'���M�*u^�+��$�TՃ.�큕�]l�[F��~(�_���g��@�EDL�IDŋ?F����y�����?q�̊���֌�����#"M�D�Wޚ�gމiQDV��/={7Ա���.��X����?��>��#e���t��;}�>�:�b�]Y<p=�`g�K��\u�'h���TN8X(��dRTV�����mx�H#ڳs�,�0�������������׈7�ȡ#��8T����q�E$0�pᐽ<��h��sy����_�q"brFࡤ@h�Ӊq�B|�ʾeI��B��/;PFk�'J����%Yz�,�'��lg��A"����E�z*�����	z�j���8y�IjrY�u�������R}������F���/��N�G"�v��^�o�fv`n�G�:��!ǘB��|F��W=Z��F��+43$F4�*$��C�ꮖA�S��4|D�8�Ջǆ-?G�j���qCO�s�q�;����,�ȉ����o��P�.��Ě�͊����D�(����m2�8\d�
I�\Ӗ<���"�E+�1CS�r2�7�$#������|`�^��_m��\F���Z���	��+���Z��4�>xy���_�����+q���T�f���&EĈGL�[1��Ѳ&����Ķ���Nn�1�U�3q�v�ϖ]poj���j�5��a��n[m��m��-�����CUUUUTۣ������Ǥ��<=�@Gz��q=:�9��u�p��Ӱe۞:��B09��<Fwd,p禎���h"�X���X|�H�+Om�h�p�܆����A�u��Vsh���=�I�dP�����dB�^�*oY��ۨʽ���D�K��u��Nd\	η���[�b۸,\��7j����m��=(j-�=��wn��Ij�We�t���"F �v]v{q�ˮA�ݱ�.�z�;"rtg:�NG߉�F#��|�H�������s�Y�����#��=�&V��gf���*�2�uz�塮!F���h_>:	���D��H��㇝"͚�<��,�8����틽���0�R�U�v��b�D�$n׶2ņ��CH��V߽�`D�F������)�cU�lm�T
��Kl�֫�i��@�:o�W��H���)�Wz�	�"�1{ﶔMu��l����m=j���}�B�o�P�H���#xՐ���7���m����Jk��G/?KOg���{8z�0�ر�0,�i,�1{~u�"Θ��?�}-й��Ǡ1h�]<;���}��k���
�r��І�����~#���n���<[IӦ�I��K=�_c\t�"�z$�{�q�;���ϲ��7��d�$3s�%zj�r�p��_=��VZ��Xă���Zڦ>��}���2`����qUa���U��M�^x���q��cY�yn�`칆�m�Q]��c��Q��/��9���5���^E�դQ�9��=�_x�!B����2(@�^^�>�a�ލ��aq�׾U�2ΔC5
��=Y�JQ1 ��rK�����DM��|��t �L$i~�8j���B�h꣞�/�fɿ
B��}f��fg2V���z9^c�t)��_[�1�wM1;9�onl������c����򂅲���5}q�':}7އ���x�y�CZ�]�95�6F��վ �)"()JA\���G�zp�kۿ.�|D���la�f����,�C^�<E�Cb��A�0��v2�O!/=������Y����\�t�m�6_&�T4���i��-{�kч�
�͋x��y�O�Q�Ͻ��c����O)���}4P�pȃuP�=}��sr���u�R��"�:Q���.�a�A��@�EC$qhӧ@��Q=�0�^���҇M.��dY���_G�sj}l���p�"��0����A����0!���i4k�1~4��� �p���g�+nJd�N�$q�������M���9WY�l�lD����$�G2ʄ�"M��dy�K#���J{ޯx�$#Ϡa�B�s�����e���� u`�.`�qT����9Hx�6Ee}�f��8Ep�.jK��$�P��U���6�|�5c�}*FZ���Uǘ�f)}d⍿tW�������tP���lІ��4���,2L��ű���X����wwMa�����x%�}h��ێF�i�<n�����]y���|Z������kޛ5aZ/u�Z��V���n+q]�V��]���{%�g���Dؔ0��B�M�nS$37Lj��I�*�mA���\r+(T]��G��7�(3��2���Ȣ#/�MbAr�:�]"V�!뿚?K=@�j"�y�C��ay�}�Q~T���^R�vhq�!	c�ǟ�颾#��#��N��e�b����`&�����r��-��O�>���M(������\r��)L͆C��"O5őU��E�,�?l8�f'l8���n�ų�a��$���2~�~W]�
{+�Y�0�xv��q�4!�v����<,(��(�<�*C=]q�������)�ٌuǧs�,su�=�s�8��V��2*I-��W��������=ZŤ .^�q���(���!z}���J8GA}(�ى	s�L���<,�x蚅(���n��V�������O��b�A=�!\V[,ž��A�bF��|�SWY��J�τ��A�&���=�;48���;�4=��7�Ё�s`q~�{��ݴ�}kޏK)$�b<h3�>���t�ne�2m�Z'�`��EY�rt��fQM+���\���g^>�}�����!�����˿>cn���^�+����!}��7k�u�H�߈a��EL�g	ʋ�գ���p�'A,�w���i���4D�ײhi�M���
L�?5��Ǎ�Ba#��"�̸ʏE���Ƶ�9��s�7���9�n��k_C�9f��Z�0lY}v��o��',9��n�C��m�*Lj̦;�.ۻ/���|�2�y�d�5a	gG�ϋm2��1�s�K\�(��&���Dz\l�B���W>��q_���c��r�^gM9�܅������>A`��1E���;T�InDY`�TY�eL�t��t������Hs���4ی#�:RUH�%��DL%��}c\6E�s��W�6	?N�8`�?z.��0�֔~��P��^詛�"�X��-�ї[cHG5�P�(Jӆ|�k�-N��ml���m��������2W҆��p���cil�DQ�&O�z��o �/�,P���r+$����au�T4�ǽ��Ԫ�Ĭp��W����n��-n�!�L]kZ�kY���C��/�7ka"(Y�Wz(z�$0N���x�۶��C�f͆IK~�y!!�̒���j叻��g�Y^�����L��⑒��i�vl����w$��	��4N�U�M �,����|�|Ȳ2�� �V{ʄ�����B�#��YLu�9"g0��x��?CM����>9K4�tE�kI�Y�)B8Q�W�k��,�#A}�ۏ����x<��+Ɯ��6prDa�[�K")P	�����j�,yf���8XF}��=2}�(݀��R#"R�*���ᦗ���s&la��ʜ}��)uǛR��'�U����2̔�J�9w�v�]`���f9+�-�9�[YWBޅ���X��a����'�1w�&���K�W�L�F�}�#㵎p���S��61�n��i<�-���ζ�����r��H[G):�=K�X�4	Cv�|�Tǝ�[�ɗ��wB6ƣ���{ab��_:�Ae� fT<rS�饕Y�ir9�g*�̏�H�1N?aS2����b�uL�m��!��Q�JS�A:���1v�o�5q�5�d Rw��a�̫�i��jdP�ָW{lcL�b�eÓqW�����X��1�Q�ˎG�Y!����EA��\���yx7.�( ��c��㓴:Q#��e���fR9�$L�SE��aK�c�k���:v��*uڼ4E3�5|�[�G�`��RN >���������iN�vdJ�T}�K���tT�]��w����6̥���rqK5х��FtS�y���K�F'츄��&\;Q�q8�	[|�W%S�q�334�xZѮ=&�9M"��M��+�s�d�ǎ��>����bv�\���=#��:l�w+�Od�NLe���X�k+��=Xw�c��;ɤ�K��Z�]x�V��X��p�Z"�ۡ�����:�eZ�jd�7�6�=O:ΐ�Ø=�qKl�Ǖ�Գ|��$�I$�UUUUUUUUUUUUUUJ��e%�P�HM��������2�r����jA�]��UUUUUUUUUUUUUUUUUUUUUUUUUUUU]UH
&�1�ϝ��ZUr5sӕ��^�Gan�[<Z^{h�s����Þ��R)��Z�ӷ�WÇ^��#YF�ʥx�K�he�n8g�λA��`�"�̐	ݔk�^ˇI�v&x�tm�s�ݛ\���n��t����Z��ܜnl��-�H�9N۷\0Yؕp�s������;v^
��n-���oY��lݺ�v�g�v�O9�і�;��������ˠ���R`1�ӽYpM����❪.x�ۛ��ݹԜ�z�-�i�$In��3�;Z������+O>;;V�]lg�ӎ��1g��7F5®��:&�	�/���1�L�o�o�:�룷��Y���z�q��رՕץx�Uܭ͋q/rq����*�Y��n@+"�N���A@.Nl�S�ø�f�|:���u�,*.�`����ۜ%��\����Nһ�r&�p�>}�wY�mݩ���mض8l3q��]�/ �<�;�����n^ղA���7W<�B2�m˽��E�����/;��\�f���a�t��X�v9�����-�z�3�xT�v��-dp��$�V:�̈́�1�;f�.6���ccP����ڬ'!�6*��9�l����M�bn^�9܂<�s��L\�v2JuGq��om���ͳ�&w.�w��yܻWU��zěq֛���\*sȼݽo;�H��UY��E�h^����,̭��ێ^'�3n�*��64ǧc�h�Z�2����Åyۮ��;�����!��E�\���c��+tvx��v�	�^�Ӯ�����gO:8��wO-�t��P��׷/6u�����v�m�;���yxq�<v��ݷbN�j�v���Ȋ���ŴqӶ\ȝ)���j�ǝ$����X������dPm���I��!��;�'qN��UH��I��Y�,1�n*�q�r������X����������r�v;-UUUU[�Ƀ;=�JFѷoZ�tmlu�u��h��ȴ������F��p�J�/5Ŋ�܁nڎ�f��v��u��48�s�m�ի%�=k��n��f�W}���q�v<�a�v�NYC�G�=l\n���K;�XA����س��[�1�����n�ғRrLr��|��"��L�\&���n���#v{q.�Ҵ�I�ѹy��kU��ݷ����򆹭�FW	v�+�&0����<�����͒3j�����������N�t���a��aP��2���4�N$u���5�7������R�>�"�<A��A����bF���M}X�P���n�Uٚo��4.8֚���c�����Y��
��_�qts�3�ʻ&!����w�u�+�0�ɼ_D����0��XH��N��Gp�~��+��@� E�vRg�}�a�D#Z��z)�ʩ#>���A�F7�ޛ�8�hm��H?j�k��ҟ8u����W��@Mt����z<���ԍ�4l���g �*8GEIl�*C�v�fs�]�ϓ�{U��*v�>X<���DR�0G��U�3u�(��	}��@��yEiV�����	�Vz��WL@�ξ'�]�X�8�=�a�����G� `'��nK玽�a�z��4`3]롧-#O,ψ8���R�	��&
?g�6GQ�'��ao쎆�L��OJ� �^{U���C]��9�,�ѯOC>_5�O�J�#��"���[�utm��7���
�7iz��p۬ݝ�n8���ZJ�U���S˭�׺V�$Mvw�.�rT�֨�bg�;ڣ���G �	�m��D�ʾB�=Hnk�=���t�,��#d*��/�h�14�|H��t����y�4��	d{&(i�=��B�z4u���+^��RE�s�ĉ���6f<H;��u�'W2u,�ʛ@���X���Z��-��&�4����p�c�2H,��򯸊"�օ��''ފ�HC�a^��E혀ȏ����=Y�l�c�3��� ���4���=�pO�R�E�Ȓ0���6r����gll}����-�z���eʃ���VC6l��Ҿ��d�q-v� ٢�x�)B4�d�Q�*��w�y���htol3C�T����w�6kA>E��mI1��1�Xޱ�H�E�9uz�q#e�:b��M��2�6�g�Q�=A2�b��T+-�����mu���o]����#���r:ԅ�\�L���*����ag��Gս�C5q[6<���-H���Me�OEK��I�/���Mz�g��]fB�YQSAm�ڠBۥwα��ge�j�Ac�\K� �)��x�����eA�	i�Ԓ?s�w������wgN40��_:da�Y�ߥt����g���\W�Yڌ�T���E��?2#�1^#�!G�h�:E��O"��&����B�B����� �&����g��{��nN>�4�p,̒�S�k
��YGF�?\!�z"��F,��,�����E�g�
��g��v+z6���"��^�K�#}	JR����鮝+<���ʋ�w󡦸�0�6a~�1_Ce(^���@��P�*�~�b��� �Ǳ-�u,<�tN��&�G7��W�^��=KX	.*������5������;�D��n
��CL������WIY����{?\Vk���S�%�Ҏ%�iWVzՓ��3�;R3t��_��pt3dW(:f�[y�TC�4Y�I�j
οMY�ȳ:B6Y��1�w'�Uo���H���*k�Ƿ\���ђADZ�%��#>�BL}��VQ�鼞p�N�`�@��l��>\��w��*YEj��κ�%	}h�� �&�DL��'Y��>#���-AO��q��Sf�(+�8箫vY�ud�X�z�p�pjηK�=gQ��[=��t�j�S����v!�g겉���k�܈6`��8� �+b�����cQ"����b�����&žH(��3ކ�\��9Xƴ��/���!���c��e8���H�:��au]zhf���\t9���,��&Hf���jhi-#��dY2≌��X����!�̃o��[��ȇws�ZH��x���m��&D
$�#*�P�����f��/z��`gK1K�`Y�C}>{0� �H�F��Y��:LN���4�C�e}I���]�(��:��x��V�Ig�8�P'  ��80��k�&��i���Vu�+��L��нHc-�!ꄓe�}:u��(�D!ed��J�CNOvC�[�{�!{Y�Q��ݑ��|�]v�]G��'��Y٦/�Q� ��y��8]E����t�fK9Wqo>��i��L�s#��w��V��(��e�	DA6�qZ�Xg_>ok�Z�u�-�%��!��T`��^�E~��_(��7/�f��rjDqӒ���dV�K���d]z4���:L��z��g4�`�j4�न��1wպL���v/գL���My���u��u�F��d�r{�<V�v��Bu�҆�"����P{����CL��2l̡���,�c��pܮ�=��D!���c�XFu�:�"�g���6\R$N$q�xzQ�ѯH�EA!�]�΋'����!��S�~_o�Dr��L�wE����n��{&��p��2�� s�e"��T7� SZ��� uW��8����#m�?G	.�����d2�"TY��hQ�y�T,����h�J��k=^7dO(�EM���}�̏
E"o6�nŲ	�,�'"�s��4Ġ��H�Q���Ē�0XXB4c��vt���w�����>}3i�gM}�],$�AZl@ެ�튓A��Hn	]!w^�,^�zP<���<P�����=�tv�*�^	`��\x�"
�#D?Bɍ�	l�$Y�	a�`�=�y>ϥ���N�ߥ�N��~�ȑ�p���3CϠi�h�0���Oה}"����'s=�2ɋ����yu+`�=��û�(�% G�fVf@����uw]v�]`Uj�9�#�٭�������խ�ٗ�]7YG*B��]��k����I$�I &I�H��UUUUUm+N]��a77`l��<�[V��5�=[v�b�[����1Ѱ�v���re��S��n�*Y�Z�[�$L��=�w,\n[��v�����]���nS�s��ݮhU-��u�N��f(w��@E�SA�U�,;%k�����>ݻ���1gv�<$��=�qA�yq�<s�I���xY�ûe1�Rm���؋�����[���U�JL�8�g7��t���_-��s��	�nT�8�A�p#�7'߉�
6GI���N������x���=!���x�_���ٳ�i���PG
1��*�p8�=ރ�ފK��|F/q�$��\ŧ�\Bya2���Ae���UP��Z�>���^�؈^_�(ĩ���%D�t���$���{���<>B����0�����}\ˌt� ��c���q�g��A	�^�; �ҽ�b���T_���J�en -���=;�"y6g8�,�8��-?@����}(oa|���S�,��,{h�uOw~.����R2;�N��X#W*��4�-�|��2�qƓ���G6~�?U�|EB�ݿE�9A���@�8�������gPh�Hej�	���+�8�lh���f�M�d��m]�08�j�R �&+��.F�*S�����
T�HMg��/	%�ɍ?O�E5�w]z��M0�����	8�"8��W��Վ��C�Ԏx�Iw[�cPF�3�J� Ϯ�����z���<-�܈�==Mڎdu��G �l���S�4d�϶p�ы���*MX��P��TG(ܵ{�zeg��PdT�y�p�3��#�}��⳼↝�
L�?KH� �W^�ءF�α���_4C"LL7���5�$6q8IΧ�����)�%�#QǶ4��aGO�E�8�z0Yiu�__g��hVL��}��݄�u��z�s�Kcw)շ�e�K��QV�4&��.�o���"̊Y��qu�����lY}�W2��/�B�3�XH�"x��|�C���2O��Q��!�FF���B�?a j�S�X(�ξ�K��]@�����	�$q�:|p��!dy7����r�A�G���L���5ZA��<׷��B��α�
���j��yl���ȭu�2.>�A��R�~8�E��V8�PU�di7�}���aѤVf�W����&��m@�BF���P������S�{�^uE0�h�(U��$�K��>w���#�
�A|��_6���7GHY�6��q�uo�jD���,r�Z��%4 ����ۛ��;O�b��(����G
��]�b����R�;���:"-q|cW�6��˟e��f��uKkr)A��th�<5\c�Y9y��5�/��).�=��n96�9��Q�]�l��������kmUw���WF=K��Q���n��+���a��d/g�ΰ�?V��Ά4�j(l��!.��uf��|�Z:B6E����L�[��Ӛ����-{/�t4���;_qϷ�H��\ �������u���b�G�0��ˀ��E�N�P��g�MS��z�dE&��3֘��������y�Tm&H�8rIc54D�ߒF�����ڡɕ�Cd@Q^�Pg�80>��l��9��N�b_d�F�g�-aU�yXRװ^N�f�����ATU8L�}����,w+�fuF�yN���"m��uy�>$��Φ���. �־���RWF��B�Y�؅=����-P����%Z�e�G��Q��\z>�6X�:�.�3h"+68f�v��|�@�8�b�L{%
w���-���W;�k\������^$�Qx�}�G�����I�a�!13L�;2vnz/�x!�z a^Qyk�:sq\����\@}�b���D��E�x�}~��W���lV�\kUX)�§W�>)��i�dV�c6u��֏": ��=qS؈�^�Ok�=��(��c��막"ȃ1�w~c��{R �d�w�����?zԃ�yAbW�來$��`��ѳd;u�X�w��zHs[z55#�1il�B���ZC!FN��c��߁Q=�DYYl��-hO�U��	���lG_��}�l���0�~OO��C���	?d�,G���>�<���ʴ�]��!E����ɺ��}>����#|50u6B�,�'m���� �m.��Zs������[�N�(e6q"�Ô��ϥs���ȷ�����z���4�r,G��U����@���{3���#������'%�+L��6�����ƧU]\
�9�E��5W��3�4s��QҘ� �{f�[���!����)�8�4�x�|��g����X�{� %2�ݔ"4�ͳF�U�fg�����j�#g3��HgoCA��]杸Q��ukFM�
���:���-�A��xQ���,�`#�(ά2{x-�LȔq����x���uόF�Y:��@�0���f��^��ǳ7�9�/�=�E�B�x��mʠ��B��t��"�jg�uz8�MEz�8ҁ����b�?�V�:*;6�W;s֬��,����`����6�<<�x��/Qk�0�Ҳv
�B�Ejn[t�ָ�ʆ�:�Yk��l3�rZB<E�DUϽ���is�D���ƍ#����~��<�P\�!�_EB�Ӏ��#P0�d��G��c
#q�\��ӆ'���@���T8��쨛�Ui0�^�i�|f��+���Ŝ�^����!��n:ɡZ�i�CCH������x����}=�V�珐o��m���(�DYf���}�>��[�=Y������ȳ"�H�]z/�&�
��,K��N@�?M�'�g4X��#o�B���~�v*FƤI7m�(m���O���&����D��$��G;��ӿ��2|��=+O�F$0A6T�t��40�8�u	�ZӧF��w���!�D�D���X}<�d��tZ�k���o��Q���9VF;c��Ճ�(1�al�%����Y�|�&�#|�Z��_[�D�����dUd��)&|x��į{�B�.����h��3Y��*�zD82��&"l�ph����;2|6e�u�z�;٦tV�зZ��r�g���mő��C
[k[���Yo�M �lH#���;4�����UUUs� T�簐�UUUU	@Z�k&9�f
�%c�D�w���>#��Y]���xȌ\ ��֖�����IeMc�+�/u�x��=m�N�p{vc����6Uwgq�tO�*q�8x듰U�v"	�ƺ�-<�wmq�;kLp6.�w�n���v��[[��4�I2�D�m���:����f{lvԮ]���KG�9;#�ig=m�t����\�9��sěb�k�v��
;Q�F�3��qay��nݹ��4tvygh�f�������7��+���9����e!J�q+*_yݑS�$�@���(!�>���y�S�D���e�H�b�֦D���4t�^w��g��A��$nExKBp�"��n("D�o��GK���g2����E!^�%���������#�B6��Sa��0�8���E��.�H��PODD���_�x���;�?_�q1�2q6��n���	�0"Ј#������jǔ��q��=׼(X8в>K���i-8�/t򘄶}y-��Qhn������"òA�K"��>�M�I�8�Iv4�E�Iu�_q�+�0y�>s��[��!�����os�X��´�$�_���YF�ԁ,�`X���T��x��ؤ�G�7�FF�Ū�����v�5%B���o�t�f$A��!e3�L���g�;(N�au�и��ש��6�"�9�$Iȯ!���~��?\��45�R�� ���Mc�`�����N��6>�;5�F��B��g��nLv�:�P��r�]d�7l��:��r:Ɇx�-=u��ɠ�=XdݦG�I#i�"0��+�W4�E$�����eպ��#f
P�do��\��]~�eY���lV����զ���]1�@��0�3�xi�TNDiH��(�H��(��?�e�F��-�,�~��NÕ(�1@Ȩ��w�DT��p�r�r�@�j�`����L9�'X��	��*uc�C��J=\Pe*yzʭ��T`�Af�Y
*�"�^�sZI����H�T��n��}��z�'*&Q�*��w��E��.���u�«��gO�?Cߒ%��"m��ɋ�t�.0�j�Ha�>�c�"ٚ�a����؏���Ȫ�Zf�i?]�!@��|�`��;�VB"� A���\65 IϬd	�&D�#�߭$`L$��e�$1��8��켦�=���*�fMY<�|�HB��$�s�Ȭ#E�H�\F�MVz�YP;�W�g!TN��dh���zC"N�ү(��8h�ʐ�BTq���*�Z��E
�o��!�������RB���^��ý��lV�}fG{bz�$�S�i���J�1�s!�}��c��!�`��Q�%��sW�m$RxM�y��=���a��g�s�O3v��dx����c�M@`)-Yb��������0�=�a�V}K�5z�����%���b��8
�2<��8_H�c�br���^�h\v��GG��={o]t�Gyx��r��H�^��}��C���bA-Ƀ����P�
v��}����w����-��# -�qXn\Ih�k�Y�#{ފ`��s2�f�`x���$�wʮA\��[���\�#������o�.��J��$e� Ѡ�.�'�O���KZ�~�����"7{H�\jN׾T,��:C��@��Z$b�K�O�M ��љ���4��1&�ηlqwL|���[�q��l�2hTd!�H�P)��eIfD������+b1��f[�#iю�%on�8�Z�.��[�Q�K6���'q���1�G\�/"C�fU�4���j�r7b�/{�Ww4R�ط�im��[���V��8�<e�t�M�\`������<����ҕ@��P�Xܬ�|]6ۊ"z�<��v�6�)�v^8;�vev��F��I�ki�m�|�φ{Ĳ�ƷNL�[h*و3�c���l��5�;���G�����m�6�>6�I?;��y�S��r�ЫAz`��ʩB���I�o.\�^@j�8�T��wT�˪��J���`�tf��t�r���=��W�4��;n�Y�Z`U����܂�>��o'l����{�
UWc�p��4i�OD��k��'�va���T��:��e���Ǡӥ'FR2X�z&�x7h��gs�Tj�Œ��j�}����a3#E�xKҺ��h'����{�2{�����l���v� 귯�Q���g�����
��Ct�V.z��3¯c�4�.�ݑ��K��7��,��W]|�4\�{y�Ya:�fVS�`p��� �P򲮻�Q����t��F�'	%)w�{	�c� jj�I��iTƶ�N��2Q�-����of�LXw��-!���%���:vv�;�uheDN�W8���oo$7�m:U��m艅N�]��v|u��~�"q<C����&��-��Ї��|~u����b#���yY�	%�c螵"�(�Dq�Ӈ+ �����ž��Z�0��6��9d�x����3U% �m�f�ۅWҨ��D��)���0hɃ� bv�gd���:��DS~�@��FA�O��<�����B�]REam6�ߎ��5���n�́�f�rs	g)6D��p�@�:\���dh�#R&G9R¨x�;~��ܾ��$�k
5ﳲ���*\�u+�a�*�~���_����R@��l�!��cV��x��Fy^�
ϳ�o7S��t[�z��v�6�n�dH"1H����$!���
� �?{����b�A?5D���DU�(�KI?U��/{ʸ��.Fh�"��Ȓ�#�^�W�T����CHq]�fg_�~r�Q�kc�K>����r�E�b&U���a�5��>��:�Ao��Q:��H�v�o�G�(����ڰ�Y>YbF�9ȞAh�eN{��rl��̱ɚʕ�z��twp��Z�]�0�!�j[e-�[{bu���B{ʮP;��B2���KJR���ݚ��!���m�H2��� Ҹ
{p8�%�� uU�<F
BIɮ����!�7T�bs��z~h�� |Jꈉ��Iio�Ȃ�+�J�pK_���{���q�i��"�PFQ���ŀw�L��Z������
�[\�d\٪=�ԲU�/<Ψ��-ڲ`�"���DF:�kH{R�
�!e�u�fl$��Fme����Ė$nf���H���[&�MQ�5�v���x��4�i=��[ޟ�B���]�"�-��0{ 9�,jw�.(7�"��;9�.�F�D\��՟��f��N�d�@��,>̯$jH�r��T�W=&�f��#�أDn��E#���B�j�og#��f̜b�c]�ͭj������*\�Qn�}\GZ��^W~n��Q�;s��*���}|�,;~�I�x�:a���,��0���b��KC�s�6A�`��&8�u�_�d���i{2f�h�XǺ�d`�}�篳��p�9��+��A{�2������p, ������>��F�B�2H�M'Y�K5�#�p���ze� /m�WQ���39sv	ٷA��¹v���M掄%h�
��Q�f�j�$]��f�qب,��烼ݠ$�b��v����͑�G�s\�_���f)mW¦c��t���ݮ�U���gi7�Smx�d�8��d��e��~b�p��c�m�k���.�Ϡ�.ˢ�|�r���̸�ag��UU!���w��%�@ ��g����#g(���mSgy���W�&*Vl$-���lR�aD�`��ݓ��˧4�!�6��|�b0X����Z��m��]@���A���������uۓ��z]vݝs��,��7f;oLa�.���,���s���TA=�S�0����٬g�P�`q;��q���<�;kg�q��O�︥Ԡ��Y�s-/$��]���`�0=�	ڪ���1�[�i��F뱮�-��;q[ۮ�db{T�b���T�ƺ:;���Kt �PY�sv�`�g=�v��r��T3�7�e����6��{[���r��;[r�yG���̯1�ڭ�TV�����g�`��y7�~�'��=��o�<}�/��f��J�0N�d�s�7�Zn!��+�uG����7�S��7஦J4�]�Kwݬ�b��\�q�v�"ͪ���q����F���0T����緍���a�=!�����8���?].��m!�M���
�'nL����'ս����v{�Ge�������9�ۑ��f���O��S/�v�����^[�_�}b�_��O���څl�	T�BQ��nQ��vh":��7x�Ji��Ύ�,� -G�BۯJ�k/hE���m]\�F�u4vw������5���ȷU�E
&�DYf�����g�P5�/l}>Y]X���|�V=��VC�;<g�]�|��(P�����!��\��y�\#��C�d�g�O���ŧ�Q�3n�����Q��'�=���<N��4�ˎ[�#�=K�]\�TԼ�x��j>YI�(e��<B��f���~Ҭߢ��wo|�����%n�3Әk�y w��q�_;��u��F�`�C�N���h�n3��C��^Y�+�eG�\�+��UT�<��F�a+�s{uG���xM4o{L�M��Cn��\uEl�U��l�qt��޼;gE̤F�,ya献�fjy��MB̋�q�\�}(Xu3lk��'�UsL��b�F'U�Àأ�X�\����P1�;~��腮B.�β͑I<�sN9gN ��� ��f��9��i���)�1S�^�P����E���h٢9#��؋b���ۘ���e��:�ͮ׶��k�_#{����BX�'�Pf -���\q���,��U3o%e��\ΐ�Sn�HM�q���nM�u��瘶���q�+�b�ڸ1>�L��AI�J�R�O.��(F��1O��!��9[^�C #��/�QGU6/\+s���6��3��^��r��8��^�O@[�\�mq���:�4չ����X��@�;~��/���7|��e��z���DI0�[���w=��ܭ�aL�:E�]�f���v���W��d9
0�܆����):9A������2�5�Ld�*��4F� Ev�P�C兤\}�nCqpaB�/z/�/���?<��pi��t�'�P��a; ȉ&5T2�oi��}��;�����j�.�h��IV��_W�"� �_e�t����X���wb7�¨۶���Z.ᣇ@�����v��FCʤc���Y���(�Τf�W��;
.���6��4��ї�l6���t<|�I����(������Ӏ�n�4�}�#y79�ӏ��܍��9�7eY�"�u�L�*�æ�V�h3���+��$���&�bD�Mw|�֘�-��Htt�w��,����׎=C AB̧j)��6�"���T�|�S���͓�A��3����+��u]n�xC�, �;�so�$q<��Jэ��<���s�u�����r��X�]b6.r����p�f�d3d
й�,2 D� L0e����^2�F���Fh�Q�@B��. �ڿR��UW����,��}�C�'+4���&���,�5����0�#/���7��D~�e׬��3w1}݂LS���!�j�A�횠C?L�no��2���ޟ���g���&����=P�)u�=_7�ď���d�+%QI,{Z}�?�zs7y�T��\���0Х;{�C7�� ��Y���;�G0�W^l�Nr�hUk�;�� #�����#�0�i.'!%$���w ��x���ʴ󧔋��z{^K���E�r�OJ���+O-�޻�p_@��ӣ��JL���ى�:�,%F$��h�l���ޞ��F*4r���xq�W�%���eN�Dīհ����Ou�;��J����Qw�>;�Zy}�-��%E�P�����{}���s^�;�T3M#�ژd\ܞW3����G,��˻�H��l���*Ks��V^p͍�����_a��/>��(G9d��[U��*��5��:J��:�F����y{+��n3�L+�/%t��p T(���䲃�=�4����Q��-6/P�.��Pe�t6���՚ha�t)��+�U�*.!��!���/`��F ֐ �tp."&%B�[G#wΜ��n�|��앵t�����r�����:�a�١��4�����
�d�Uz���H�XG=6�������A;6C�u��������1!H�*���u�n e�@WgQ�p��[,��@Ꞷif�,��-�Tn{� \w����t�U8���T��U4�,S�7k�H�a%^2��p"`�ޜ���Wu�A���Z��o:^fYXP�D��B�cjD~#H�PVz�#��$W7|�!cLc�K�н�ӼB{'/���؊C~�C���3[�	�O�'
��#�ku�
�7��3ɛ���)�(j�yr�����c3�E]:A �7�"2���mdd�A~ܜ��uA����7���uٵ*C�֨�ot�˺��5��jF�d���oc��k���һܝ"���I$�IS�%$�7�o���j����H�m��m��N^���x���a�F�� �;��Ѯ�$�vM�ջM���p]�x��v��Ce�LkF��CyY��viK�pl�7�2cm�3W	�fP7Q��k�=�Jwj�Y5�^Mcj���i�z����cs�q��ۂ4��Wh:ڹ�W&˛lN�cO7\�&�vM�y�rX1��ұ��udDaF s�B)Ek/Xxlհ�!��u\{g�����>g��7j3�\5�ʑ���3�2�� AD��՞�Cc�ӳ˽��AY7Ƹz�%��H��Nk�<���qw����y�,��ҏ'�a-"�2:����li�1q��y&aA8��ȃ�I+M�u�G�i�Y���͚Ɗ��M�$�@a�H?9�\�wr8c�-*�s��mX�Q��èIu�w���@i�tf��cc$�޷��۪��Q�i����`l�`B�D����k��F�"�ގ�0�0�s]���>���34;������0�?�}C:�ր�p�+���F�)��O�H'��7������v]ȭ�
 g��\�$>r�$t�x3&Oyݕg��|E���y!��x��
��d��v��]���絚D��A����0�W3�}��0Q�`n8�w������1(�^�\��>S	�4��z���w��^`{5��	Ӱ*Ԃ2++�H���O$�W@u�m��i�h/�����U|��U\��}=؁�2�[����^3�u�Rݺ���jǛ{n�P�{��=u����tN�q�촶��5u>^��x��/�{���qk��>^�f��:5
 A������z�=����&���<F����3rNs�H�������@[� ���$*6؎%���ile��7h/���i�&�[���~@V�Q�k׼S�g'ݘ�Z�}C:��.�C��Y��:�V�Scd�plw;�<��@�H����2�B��.�}�
�P�<��Vd9��\�,�[s���W����A�Z���sg+@�`�p�	����:ʬ�N�0�<�������&/=sN�0�����&� �=���ξbܢ_���O;|�ї*�i�U�O͜��l���񩋚y@�0�n�-�@�&Cp6Ӑ��G�s��{����s/�8���h^���W�
�� 4�Z|�]d��Py�75�7@rVG��Z��g
��@V����k��FI("������-Bw�6W:tJ@2q�s �y�COa�o���s���B�Z\�ay�CJ.t�Q�@���'=~�41�sHL�d��B�{������/p�����vρÌ�������:,�']�u��`�c�V�=J�m'JK��3�g=�?o��Q�~�f�7URDF�<`�;�y��5smit�O){�(m�}��PD�  ?��\@d|ݦ���\k��.���X�h&("�4���8@�����װ���z��ŭ,��(�/�}L�.y�c���~�CZ�+� ���V	��YB4���#���*�P�ch����9�~<P�,�8f����,<�	�1�M)*�Jj��\�\#��ul���K\��缰�{��lF��d=��ÐNB��j�B�L���Y�����fw	��l��]m�閅cU�R�T������6Qt�+�$�>�4r �* o��g8ZC�*� �9q�8Ϭ�3�FD��@`�9i`�vi��mW,���^�4��;{$\���k5�.[�<�F��,�����4���\6x�q�!L�p*t��7:��� ��	6����4�(a̉�B��T����l��kp�h�w�XGFg�X��9e�}<�7\�n�iZC�u�ꆸ0�,�
k�<v>�8��f� ���a�H<� x����@<yŤ�k�Q�r�0�ݥ�Ux�N�n''@R7�U$W�ђ%�v�ܖ�v�����meN��6�G�L�.��	�[��{��B;I��<�9�q�/+�%s�uk�|]#�u
'� (����k�"	 ���d�4 q��5оd@�O ���x,���W7ι�\�@:��� gvΐ�	x6�p�n3\ g (Q���k��s�6�k5	�9	�CO�� �˰�k�o���^���:G38��]Mf����ㆁ��t�y6r������#ΐ1!�~�8=���<y1pq�lgx
<�AB��ۉq�%|��w��s�x�V��Np��A��0�K@%���;����xk�M����:y����+}�f�0�� �>a�:y���g��\��:X<��W�p����8�%��D�$#��9�s�ib!�4v����l����g84 �_B��8�!�p"8�s��ގ��x:���3K���(,�@��*��zv
X8,z��'r�I����O��I:�.+��A�O�0Yx��"�:WY,	�Sحt�hv(���+�٪[��ps��]tXy�8���8��m$%ݣ�b���襔������87S<�sL����a�N�<�`t�3���<�F�t=����@x�r��w��.u�:�x4�� (�O"�9�9�f��p��.�4�T�KO��5���G�X�r�q֞���n��ո���k�n-/'X$����w<�OQ��)u�L�f����������������x�ʿV��O,��Y�R����,�"^�T��y�K��C�xް8��n���]���hs�x+���4�
#����ߡ�29��[C��H�}�߱	�{�
&+ K4���(����,�����\�a���V 6��H���G�3����m|�� Y�2z: i�x��q����{epz��+Y�}ht���R�@����@�		
S�i.��� y��(z�iP�C����~|�8����hs����]r��s��
��c$k��� y�(��W Q�8�w�@�3-s���~��[*�@�I�h 7W  Y���Pn/�e�9�xiE�5���������y��pr��d�9��3�
<�Y��5Z���< TCH�,�m�J�=+��89�=��x�� 
�8q�<���m�dQ8Le�s�t�'��8� U.pv����u��:y�#��� (����������pt�	k�f��-�_�L�a�[������p�s�������9����p�s�����p�s��� �9���p�s���� �9���� �9���p�s����s�s��?�� �9��s� s��9�9�9�s��9�9�s�s� s��9`s� s��9��9�9�s��s� s��9��9�9�s��s� s��9�G9�9�s���8 �9�s9�9�s��1AY&SYp��P[R_�`P��  � 7'�`a�����T��$��ER�٤%(T�F�F�`T�;M$ْ 
(�(H6�PEUEIR��0 8      :�4)l��  AE-�J*Z*�U)D�DE�(*�     �4��� �IPP �G�����`��lXX,�ؓ�k�gwנ�Sa���;���g�v��;{�}���ӵ���wm��|�oo>>+������.{���}ۋ�� \�*���� =Nl��:���o�t����}�@��!�: x�J =x|}���y������<���>�8{�>�����H| 6UTR  ���O=��� �ݚO@��g�ր����y��z��)�4 �{���>c�m�������-���@>�笏�@�(T�x��tf�)�t|{�p:��zf� �p��}r����^����;�#�ޗ[�u��u�M�h��c�h�wu]݃�%P� �DU��-�]�l��q˻7�9�����t믐Ҽ����7w}m}�*�>���n��j������@����xw�/o�ѹ���im����*T�*����oA��V��d=�����c�G�n�h����g�����_]}{������uֹ�c=4}g�} ]�(m��!^��	��h ō�|�o{�������}�w���c����_^췛���:w���Uۗrۻ������[�/w{��籶���0��N�|R$[H�
�P��\�{ݼ��I�y��ƽ�,k�ٷf�\��n�����|f=jo�=��w]�un�־z����S����ik=:�=A:| cB����f�;�]Mp�ﳮ���qK���ݜ�7��{1�c������u���f_}�7���{�m�sח��u�tz%R��D [=��n���G��6����|���9�vu��}v���}�w����J)���W��}��/���aw�U����j��omh��+���|� E?	J�   "�ф��@   dL�SRzLa	����D%)J  25< RU    �H!*!2 ѣ'ߏ����������aX0�N��_��濺kZ�?� $�L\}� 	$�` BI!�$ $�O� �Ib� I$�� I$�H$�,�I	$��)��B� !���
ud
�d!����6�< ���V�(7�?��F:��J=�H�a�.)qЛ�l��fb�I���.4*`�kf�@^\3b4��,��sњ�s�.���RP���rd2�!�����@�Wj�Dk0a6l�6H��7�b2�lU�$U���[=H�F6H�����(y��7�4v������vv���nef�9u
b�Џ3[f�pSY�.�MNGX�7 ��R$�
��P���b�m�E-dG��%�����e�RĘxm6��;�Cr+�7zt㳃eb��:uMxr�b,�� r�f&�=Y%�  �EV�R(�yL�Ѝ�w�TXvj�h��v%R�aJ֎��e�wc]�u�d��B)�T`��V�C��I�T��s$���5f�rf�f"�ӹ�$͂��P�PY�t)�l�6f��e�j�ń1�X�k�܊Ļ��4+3j�cO���4!f2�i�P�C4�:�X���-f�K�b�*e^V�xJI�.� �!���A�l��-ֲ�P7����Q�V�򕇆<�hn�4�/�U��"^䠔4-,�hY�ێ�5�KV�oc�Z���4�,�wM�� ��B=�A� ;T��I^�p�@F��0�^��T�(�P�v�( ��	ۛ#�j��h��фZ˻h���*2I�[I\�6b[�d5`�7�huV�k��v�F�$�Q����; ��B�W���d�;,A.�[{.�	f+1�@7�U ��3(��-,D�Zv��Kf�8i;4�T��f�=p��wR��t�Es%8�m��֛�)�d�	��t��^$���u�v�b�{uid�*)���wM՗H,O*�VSyB��X,R6����&�)+K�A2����c/5�#^z���R�ͺ~��f���Ak��db��D�=[MR;o#��.�ݥ�����X�(��r���h��=�`r=�VS������R��ڜz��p;�Mi�d#q����	���a�L;�
�+fb��e�%wzo �=��yG��L����B����d1�Ieb,]��#&,�C]f0h����j<J��	3EU[Ѫ&��ܪ���5�V���7�6�ܓ�R�&U��aSY��^�t[�(ET��x��R8m̙,��W��m	�t6�%))é��DBf�˺O%jWB�c".�=)r����{��K��X�vkb��Kf:����[NZV�6S��#cd*�yy�k+�WK�mY���fZɶwIe\�7w	8E�13�L�N���WF���"yES{��	�g����q޺9[F�n����:]�Ԟ#tͅW�v�r=��1�����y��.��}8�:-�37�1T�K%��j���HZ�+;,m�LJ��j����4��ݐ)kr�͖l�.�k.�n�D8)�њ�y��Лb�dR�1�M�[f�f�.�h�J�15��@6I�Ҥ��62�]�[>�{p�6��D��*�`�u{P��A��U�}uo+,L�wB0�X%�)DIƆW�DV���n��1�v@J�Q�ܦ�{�5��-Ԁٰ)�2֑�w���ojպ�k�4	pG���Za�'7p4L
��r�R�M6욳t�ax����Z��dz�È�Zo��mkG+F���t��gN�:ēV�8�B���B^w�斓9:�$�x��v��yͤc����0Z�Y��x�P�\�F{9%����e�攏-j"���
q��řd+W���l8i�Y��OX^{[�c>T#d0nX{g�f�S͡"T!��j�;% �90|����Xk^Ҵ�Z�6�]��c���/*xaH�u5���e��������m*�V�r��=3YJ��@6�VV�G`�CB��Pm;T&<�P�d� �˼�U���e�aP�wlWF��`�zV *��@�0�DdVi��xk&eQ�4�f��Q�*F^0��	�Ql�O`��)⦠�4��^�2���2<V�[�VԐ۹w�"G� #*Q&Y7��aZ$��f2i�`�6��e�Y�v�v�CI�7W}��:v��B�;p�!5�h�6ӖLN�4�)2��B��U�˗�"B��� ��*;')AD���W~4��O}����i<�c|�5�pa�Q'id��`��(��4�a���8�E���8t�̺E%�cyt��m���EB-���n�4��$���A�O6�ʗ=���~F|c���4,�#����������J��6���9G�[�VT�N�@�r�@�d�A��Lѓ��#���įn��j�*�)f획��1)Ee�2)�zin�%
;�Ȥl��,H7iY��K�ބNҼ��h�5����upT���bc�Vv�#yHӪp��́b�æZ��!���^�$MWyY��+�l󻶸������0m�yf�n$�����Ӹ��qj�(*&Ѭ�2Ӥ��-��{��dZJ���I�2�d5K0c��̓%���D Q&;g^���2����%f�N��(Q�*�B�v�Itop�0�g�c2��K�B�0��Pg���lk������Hі,=�^UNfV��l���f��f���4����ch�boF�j�a�{�㻙�Q!(5�H՚���ͥ��,�+0n(cFR�/E�÷q�O2�,�=���yܓ��+��6�<���ALJׯ*�
o��QN�f�wu�kz��Q�!��f㠩)��b�W�x�($È)����^����rAV�
��{���Z)077V�iZh�kZ�W�5�%�l3�7G� �e��j�hߞ\�7GVQ�MZ
'L��N�������{2��zP��XW[���25�ҳ���R��5�zI5�v��w���4	>:Q> �E
Vh����F�5d̎�.�B�����Z������B�(U=�CH?!�2I�Z'��A6P7pA�p�n�
�QF���֢	&�����rܨ��T�<��놹�oU�Lӛ��t�ԇ��������4 �jyF���dӍ夭ɖ�����7 r�<�C�qƆ����E�1ו�b�U(juf�:P��X �� ��G�(ijAD1�ISi�T�`���K��B0�b�v+�쌔����Q��9��ؒ��K<!2	[�tCA���W1ݜ�mE�� �HI�R���30�^w�N�0S:��y��ۡ�oCD�
2f�h�D�	�-ƭ]�H�F%m�F��V*�W�ލ?K���{x��47�Q8ș+t<U�P�[�+m+X�.fL���1��1]M���9X�u��*�XF�SV���r>��yj�Xٖ-��Gk�ek�v�ѵ��J$��5	4X�S��8U���U=SЋ��)��sٶ̌���3m���N)�= �"�XN��P��wKj����i���[͹�LB�;R@�C�ot�.z�������ͱ�L�P&�ʎ�Hbжդ�؂]d���kq��lC��a�n�yK�wh���1
� �ՔV�r�ŏ�ދ�V�,�jJ����B�K�g�+�iM�͓W��W)�
��i�)�����Ko0Y:�=RkK-F���&�(����J�ˑ��A�kԱ��"ek�iP�i�nZ���c6M:~q���0w4�'qIf��Y�=w�W.$;��z�i����*f�����$68��4mT���n��cd�L�"�.Ҧ[���wtV�����OS��Z��6Z�vhء�/'�@O����X[��N�]ڥ�Z��2�,[6eV	�*�ݨ����b͆S5_���u7�@�#qU��B��Bѽi���ֹH�3E�me���݅�˹y�J9�k)貙�+Q`��,��Q����iHK̐���۵wLщ�$�(��Wb�9���d&��8R����2@ҺW���U`c�s��4��g��
�MRQ�P��H/S��P�� � �3m�F�1V�ǯaaTz!�,�fN޹����f�H\k��
B4F��,��i�Z
I+sĂ$��/�d|���
!�Q��B��
&�S]�]m�Ǣ�U�b5��$#l�j��P��wA�2�Â����Iٱ��
����s"�f��˦�B���O]A�1Ex�Eb�	��tU�k.k̙��l���%9��L�,a�DT{J�����O]OZ�n2�8v�	'�Q�������w�m��6��z�
���'M����fK"��\���y��Q�70�C2	!� �W,�1GT37�� E1��ߩ"ETyHК�Y�����BV93rf�8�݂e�I�2玭�c^�&�)�Px����������l��i��6��6(]�b�
5b�$�5��Y;��T��lF�r�b�:!1ѫ�\��r�*�b*�ٰp�W�	�rJt!M��	��m�}��^�%U ����@��l� �-b�MM��;3w�'��k�x��(���kw��q3��Sё5A�H�[X(���l����Ȍ��"Il���m]ڣOY0�m�+�y�����B��4�[TL��(�3]Z�,�b蕻�6�f'V�Zt2%�I�pm,5^&�#h�=�����n�k�E�66�'��ef�� �� /.�x��s48&j -U e��R�&�V��(���Q\љ������2�6�n�N�Q$V@�Tf^&n��e��Pp�b�+S�V���soez-�U�R!�<'�^!�j;�����煛v�D":�Y��◺5�U6FȴBW����mR4�w[�sN��AӰC���`GI{�en������vi��߫���*�=8�K�n�L������wE��DTߦ3�uf�a�~yLԘ%b�Øl],�T4ʠ�:I!J�кw?q�7��l�I[m�*띸��wQ�Eh q�8n��S��<q�̶�� Y�ֆ�m�`9����7��2����B���a.�*�ͥ����()P��V/wGQ�k��f7�1�!���n�*��y��T|�ɥ�m�ψ˗K	�F�X�n���7V5�&�u�4�G�bZ��bZf�hit���R��[Q��>Q�wL��N��H��A��U�r n]�"9���ۇ$;l�b�F�A�+��vEF3*�U`��(�u�f�2,��Z��B(H���#d���Q�Ĭ�{{`�{L޳!�6*�P�9��36�	3%�����
f��ѻwr��e�MP�a�[j"�^���y�Rnz�A6����hlm��x2lͷ5J5�&:Ef�Yz��?i��
L�;��87	�&k�wۏN�
�f14n�
��zU���Y�B��/)5V巰U,�n���t��
j�P��n��k�El-\�3p͏t�m�S`�ʴZ�j����ǘ���L�(�j��y�n�ߜN�4�O}}�Լ��!�IuM���CT��!� x�1�+ ,!� z�4�dv�d
���+%a4�@�V@waBd����L�PЏ��XW�����Q�>���8�Ve�� o�dn+�u��q�;JvD�o#)���Xbk!8Y��VP�ܻB5C! t�mManK�	�V�e�^GJ�*ʭ�t;f�eeͽ�x�C����j�K��4��dRm?xR��~��s,�{�{����&�]� u�l�]@�
�u3��D�awd���{�$���=d��P�2XC�l���� q�+ b�c x�� x�+$�]�G�x����1m��T'P�_O7jcq���ˤ!�@�4�2<�m�=݇�;�3����T�t�D�o��g|��o~S<�o��Y'�!�O\`z�<aYABd�x�$�����RGl{�@1�5��8nI�q�8�<a��<@8�adj�!2XC�@�m�1�:� :�������ٝ�龽�����                             �@       ����s��V�&��n�    $      [jH                                      [h                   �8�  n�m&�iE��7WPūmc�[� .�t�$�1m�� �  ���  m          �      ��                                           `,��H  -�H &�   Y              n���[ht8  ��M�-    [h   �(                      �  �      �    -�                �� ��                                     ���{�w�;�@�@mN�]�NKc����n�ڰ2��W�['x����9�*QY�[�{q��n�"�U�s��Ӝ::�Nr�o�.˘�F7�L�Nu������Y@����m��il�Y���8��W��ܛ�(��K��3n�gM�t�ki(v�ճ{(�lͭ'cԧG�]�Zx������e#�1Xݖ^7�L0��`�ʗ���
ٽ�Y�)VM�2��v%ve���ֽ�D��ėg^�Èk�-u��ǝ�|�[�\g|���C�%}�c�54*!�8N��]���d=���;( ���uFO*�#ѹ�_�5��VG}�о��ӵ0N��غ�����/~�p)9��Uݒ	7ySd]tx��NSv��xɪr�=�#~�Y�܍'��P�DN$[�׀6�S��jJ���I`�t옰�s�1w*��ǧ���K[�R̫��O*+���,"(v;aj2Apa� �=X��͓��Y3iQٜ���u�y��J3]�7z�G�)t[���:��������ɤ,�܊zr�X,&l+���,<�����^=�f:َV��r�t�2�"PSSS� �YZ��"0�4MA��Ci`�%�����g��E��+f|L+
����ݾ�֗�)�����"�Nŝ��-�r��Y�>�۶s�Q�Ъ���/��>H��Qt�Q��쮪�:9�^��H3���U�M�5�oy!�j�^W��`�
vvcx>�{V3(�V�m'���R��8۝l�q�^^uV{���A�ڡGF,g=��Eb�1͕�����/r��V_��=[�^?%�	�$slf|hUŸ�4�n��앢�Mb�XA�7I;(*9�;��l�ۓ�2��zf6���;���I/��fd�a�u�x�Ե��T�+�R8��}M��gL�MW�����rt��[�Q��G���$i���D�2�ww9W��'�9WA�6�6��%�]lC%~kO�{��6�g�wsl��
�)V�A���I_w*��d33{�վ�+2Q���S�8�*Wse���$���Wɾk��Nk��ݧ\�F����]��̕��ur2��쳆�������^�x�x��=�L�ר�ے읊�*J�n�{+�jen�ZjN�Np�Ib���q:oz�� 7�s$��J6�\�4�3�����$��7[} �j$��3���Ϗ$�w"y$�FDw��IH���k��j��L5���]���/֢Ñ�ݐ\gI�����{2yL.�բs;�7��$���<�wI���om:�ll�����G
u�[0N�9.C�Ɋ�ﻭ��ELg)�K�DNj��[��j]���H����Rs��B:u�j�41(ju�a�V� ���Δ4������t�,��S8�ƒp8y�l�n��y�mlxw��:�"�0��|F��@G�tn���һ�#c��A�Mn���I����6�L�X�GdwK�o��'CC2q�\��J�@K4��-kt�e�wxc��i)�\������	�:d/he�Vi����၄�#u.�!�h�Q������٘']�БQ=�՛��t�%�u&v�5.F��;6n̙u��mJ@<.���
A����;�@�qV�l;Ih�T���\�{�F�����է'�Fu�G�KxH-�U�Q�e7P��Z���Q��l�f��
��R�ǻK�5Z*_l�9��+.�P2`��{;bb}#hW��)��n��d̪e����m�a~�,С��S�}YN���ɽ¬5i�� f#n*��_fj�'uu�cY�2nB��	�_Tg�{}��< ����A�����X��{�s�� \]gp},���RY�c�nr��Ouŵo�"���ŧ%-l��`��s���&'��L+���q`sU'�V�0���mȷNik��sH���DX E�Qݬ߫,�@�y��������gs�cm3�>�C�R�ݠ"���yӀ�]͍���-f�[rGR�-�ŞYf'/�kU�e�8z�+[�N��ݹݶ��:���Վ��{%��;�>ƌ��Sv3����襈�na�`�W� Kr��B��/,a�B����+��H�u��ҕ��S	�a�n�u9V��;�v��:��zN����6���ꎩ��`7œJuu��P�NV�Bd�����L�A6]�0D�
GH�xuy31���:�<�^����(Ь�mb��˓m��&0Q�o���B�V�a���4��ٛ��\*�>�����7��,=�V)�aЦ���b`��ו5dX�����N�׉f�*(�S�͊�:�,G�.v�k�15ܪ��N|q��;��*U�3�|� L�wd��=�����q�Σ��^f����(��h
u�}�n����X����J��wá,���x)��j���h"��D�Ӑӵ��R���(��Ƒ�8݆SKe�-9T��D��Z3�[�m]��HH���2��Fؓ�$��2љ�8�0�KN$��ph�[30���葻�8��Ez�r�Z������U��Ϋ\��q�g%
khe�r�T���>�s]��r�ooZ��Ύ��wnTe<;XՋ�r�D�δ���k7����:/�����%WzL����BTa��H�Z�K���������;�낷v�52m��6%"{��r�&�â���j�3��M�����-e�[d��	ʵ;,�V�#ٜa�`N�����r��Ͱv�R���r1[�;gf'�{3c{r뻍r��;�ܣ�8���:��t4�v���/m
Y�
!�����VG�_vЂv2��&�&�lܧ\u�dh���S��t�E���ͬ��վ���wp��\/n��B�bO.����g��{N�t�d[��
� �m�9'++���#(�Iŷ�(m��͑���( ���82bg���͗9�5�J���1\��^vA���"v���inV���[�b��kM�N0���V�d��*��:߸�8��l]��*;� �j�Ӛ/Vw�;�y��x\��,a��oR�����ӵ"r�0Y�����������E�e 2M�־�N���#+0`::䉣ΧN�Y%�"ɖ(*���x{ �x�v��8;3�)��$�v�7 ��s�ʝ�z,�6���F]�Y��^�,v����S�t���-����<��T�2\�#��t�N�Z�m�Ǣ�ť�y�˸��y�Y�SwZd��l�;��W�i�����E����sNp��W��<,L;�-�!rd�"�Ô�8�]��v4�uB,q���>�* &���׉X�p�vx�[6w.NR�@���w��j�zK�
w#.����*Z�V�6�<Ҥ��].����pQ+g-+��f�_Kۭ���68/0:Zl��:��2��t��nA�8����B�[³����Ua�f��x�nK��΀��uf�+����l�k���uM��˖C�H�5
�M,hԾiw;7�:3b&��e��qIo!,5"ևK7��޶u��Ѫ��X�-X���+�.���vfT8gvi�c3�|GV���V�t��:��-�2�n ��nh1fM����e\���Ʉ��]%��o�g8U�w��ku`-a�<��8���mf��F������%���h�ݓb�g�.�y�/ug��av�\���*�v���v�Kw�!r����w ̎��oΓ��WP���ܨ���XXac,�	;��T�%�s�\[�P�J8��1��}9��{�\u�uoP�%�h���2�#zUUӡm5̫����OČ��S�D|�]��}ۗ�yn�4���Wv��ÕY+O�luM/h�� �t�n�5�.�6�F�"��Ө{$�cm	)̛B�s��Mgw-�lR�ګ�6�.�S�C�.�4�,*���dݤ8�2�t�~�9���EU<��Lu�o��&&]�����"�vc�4��!�G	�E�lT�=� ���u4��#��AV��9��BZH��JI:ye��'r��E?\ɄT��Bi4�"	A�ۣu�4v�N�^"�zA��\L�_{F�h�lj� H�8�_�uH�M�T��Z]1Ĭb"Y0�1��6֘�IP �n�m ;�Ի��:���0�I(c)��Y|��>�����z>zD91��"F6�ꦊ�xg,u�(0�i� #"��b��-�����2S�-�)�l] -픊{��I�&�U�[�U_.�B!�����ڕ��+z��;-�}� P,7"^*�f�i�E���������%��m� L��ͻ�URVh:7�,��T�0��`��B�l4cn���r�ݐ�7�d�m���1�g���w�ZT�lH���+o�W���CN�x�A�0��$D��E���	�o�Y���b{R
��`�M�>���k��ڗT�b"ې!�q���MT����.ʠ�X�$�YD%JD��Y��~Zz�U�p�h �XYd�6q�2�Uھ�#+�"�E�BD �v�.��pu�\!/*A�p@QH!�͚N%':�Q����� "X!�{�]
Đ��*����]a$ch�9Z�b��E�M�	 R��L�D\�,p�٧]V��
�h�Rn@��2�J�{7S����f�LQ����٘K&�>�N���4�I�2�T�Mh��D��Tu��
���OO^���D��$��|��UcGe�B�'��N��͗{P�u�������/+���n8R0��1.�2kK$H�iD�zk�e�#"��i��C��Q���AG�s��P�H��@�O�2SF.�C�v��
e��j	hD��:�4��������Hѽj鮷7X�A�D%�����Rc]`M���a�Zm�����w6WU�#|qZI5H��p���.�]����&�1�V�O��TM���q��q�8�^��E/�@������u�!i	2��H���Ne�.K�皊�j�(�!��j�u ���y�$�R���\.�y��*��#��T�Y g:�I��BX+fk#%��f�,	����eB���of�j�Hd$�a��d+����B�"�T�j�򉾾{w�A���(@�4��� �!���'1���Dܾ8%ȃ�h����ՖE�@]Y�(R�}n����]�,2'Jd즁A��0�UYrS��0ڞ.Cm���H��7H����-wJ�&���0Q���kB��%�KmG8yn������`���D�~L�,�9.���X~�m�-Iw�El"���2� X��	 D�gr�cN4b�e�E�n�l:��(����I�W���`��aO

)����F�٠��C#amD�����#5��,�y2`�Gƞ0�/ӿ7eQ�Ra[�6jIx�\&� L�i���=9LY�r ���Ȧ!t�ճ,ݠ
I��Z�V�P4Da%sy�pm�ΞuU	���g��✠�Sa+]MO��9��"PL��2�e�qsm���%β]�u�w�H#.�N\yf�Zc�ͮ���0�]�wq\n46����x�jue�.��!S���/�ޣW` JՔ��˻$�_���K7]]��z�5Idb��l5�=�e��Z�SR�qdLhL���,��\�ҹ�B�_oi�#��묦��:�z��SF�޴����V��/P$)��<r���H���ê��A���tPD�l����q��(�4C�)F��!��!�[y���"�e-Ͷ�5�4��~��<�=�Or�i+xk�0���iە�Ж7�:|�1wuf�7��j�6�s�����ǭL=ih���d�&N]��&U�;�+t��Ջ�(�a��XI�!)���x1m��SsH��� �f��X;���Jǲ�����m��  """?�I'��?� ���?��I	?����}����������ٯ'��      ��x��[hm           �Lؖ,E��d-�@   [h       m�m m  �[n�-�      �-�   �       ����������=��v�Lw��A�.�꛻\�lJ��<A{;�B��Mٜ3#�gQK
�r�FͻR��\���i>��Tݽ��[׷\+A�u�a8�ä���	�k������s:-�g3U�%k�k6O<@�⮄m#�
ڄJ�#v��]���o{׷�Wn鰥e�]&�zɾы�����D�����,�26��n��ባ�s��s�Yu�f��.DW"8��86����	��9��UcX���K5P�[��/�T��w]z.rMNgl��:��O���k��8T���5�N�D�J���K�~νV���{����֡��ɶ�Y��h�1��ÜT2�t��r�{��PG�g��g��;4��4�I�x�#f�.`6�+����G_!N&�C�;�'G��H�D�1Vt4���xP�Va�Ms��
��<!U��0fv�aIjW��a��RQ�^$U
l":�wU�R�Mqr���]ݑ^W��AP�3)�=�@�#'�Dʜ�#l��q����	���X������J��У	i���H^C�T�QQ �e���)Jci�*��"�U���-���*f�]Z�0�	����;ZE��		�!�U�{�s��%L0S�aU�m%id�>A�UJ���*FЈ#�U:%E�	������)��G�i�ӛx��j�;\�'}w���t�ݡ��g��g�g�_����|�   ��m��  � m�������O��ϧ�uy���kޠZb���✼������YU��S]����ig.cl��4��
~h��$G�a)t�2>�D�Θ��h�TY��R]z2� ,�L6�m�[�T������FLU�%V�"J`A����dC��r�0�ԅ-bJ��E�?W��|������4�yY���xP�=����Ҥ�2}�h�o�� H�١�\�u-�nF�Ӥ`�6S��0��x�h(������|��Z�Aeq�Vic�x����$
P����[|Mv�>���1�7��x���B���A�����|V�"�ȋV��!�H�L��2>;>��@�DY�Y����@f�C	+91$n��@q����C��*/lXl¸!�����`|Bʱ6j��γGs���:n��	��C� hu7]:w�4a�4���c_6D��9 N����T�Q�$^�>َ�M'�}ߵ6�`�o��>����m�s;���~�n}>k�m-�F3n��=�Z�e��)$�t�R�/Z��=9;0��t3Oۇ���G�I3�>�~wn�x�u���Sny^Z��$�@)�W�{�=<x�EaLg��LÙ�7����7z�c��v�(t�l#ᄒ���)Uyw{S%@��m���d��'�T}Qɴi��˭���^�����AG�32g.�//����:p_B��ob~���^�� ,@�w��?Q���08^`wn�}�8����HC�B�y1�����G�����c=�
)h;@Q��vm�E��W*a�f����Eq���T���j��5}ju��iJ�3 HZ\b�53�$ٍϤ���__�C�y�ጭx�ֶ���a�%��溡C�6��80Mr�X� ��4{32e?�'�|O<�{��щ����֧b�T�(�,���u��S]�z��>�=o��q������w߹��'_K}}g���%�=|�$���m���;ILJ��j¢���R��۳q���"����c;֠-b`m�R��6l��  }���Z�1q���CO���;�3^��m{u=���T,�Y�)��:��V�yȄ�v�h\a�"���=t�L�GY�����\EQb���� �F
���("�*����(�V"F	�"�A`��
�b�A(�<×��S;gP�_�4GYv㆙`B����\	���p�8{�mm��<���i�f�#O���C�e?�l�Ml2�����}�i%�3��h�Pۄ�{�M�L*ݮ�ef�ݸ�����ȭ�����K��K�f�f�~Ƈ���5�����+$	�����4h����T��<x���|tp5��>�����f�0�@R퀟}�A[k�H�"��lC���U�1��_9��zʟz^3�|�o�����䄃��Dw��TO��}������gwqHf�����:Eb�_<UO;�a��|����G�.���F�꺪A�[q( ���˔ݼ���U��q�)$p�G�d�za]s�{��6o���D��L:y!���ظ�;��hu���X�>"}�v��E���"��h��/��N��>���h��2S�����g*���3i��u9���Y	 T�N Q�C�8x�����0R�����b���s>�������<�����Ӆ����=K�6@��v��!G���t���3�s��S�BV���8l��6Y�F��/B,��m�V\�Ϭ������GwxL��Ǎ�h�G�^���|�*����6wLJ#۱TXÎ��w�!U^u�y��C����RQB2(�R�Y*K[,O9���~�6�y�9�dY���S��6n��6�f�tѳy2��h齗��i�Ή���M�bZꖓ#�Y.ܕ��/����#-c�Ȭ5�4��}�y)#��`d���!\B�}hq�r}� v`t~ {��J l���H�rH�rH��[{q�b�!�R��H�P*��d���Ï�v�	���0,N������qhq~tb���ٙdWS�����=�ő�f����gy� s>��O{��S�	��f������� }X�`�vE*cj��)`'ʩ}��4I4A۱j�Q�����'dnV}Qd����C�S�������xk�"�Q��f���ʋ��a�h$�����b�H� �#z\j��^>�c}wf�t�rEH��" +#��1�L����y����Y/o��rDAQF0E�"*��PX�	 �b�@D$b ( �PX��&R��z�����X9�xg���Y�,��dw��E�VYx�W����rt�ːeq���$������k,�e���u�v���?,Ea{b	@3'����1N7v]���kĻ�m�C�dp�x�ePݽ�G��$�w=�5�xH  	   �Am�m  M�$�7��ϼ���y�~>IQ�/KkS�ıqz.�-����-%QF��ȇ��5J �e�lTE���U^���w숵I�*D`eHS�o[�Y��
�WrD��6ܒ[���r����ND�%��	$p#ǹaVU1x�8~�~���"�Y���8���$�C�Ǽm밵Vi�� C�!�t/.��G��_)��g#{S]D��́��6v}>�y˴�Ӿ�P���ugCmd\i��.��䋽�4.�wz�<���:������D�����"  �.E^�j�p��&fHCE�Q�$"WZ��h'�.ȋ���ՇE_� aԇ��9!ȹs���)�����z�R⚪��l�n�Ѐ��H>_�����Mg�̜s�_|��⽴�zϟ6ٷ�:��x��W/��+\���� 0��#�ki�&>x*R�rQ��#�>v�������-��a��ڪ���@�/C��g��D*ʎ�������FcT�������)$��M��O��HF��lěq�d�����7d$24�z����su�^����Ɍ�˘k� @��kS�V���N��,�<w6O0a!�կ
2�1�@m>n��o1�ˣ�o�u���aXQ�Vdy�s3S��h�{kٞ�**r��3�"m�3�	�o�;'0���_s׏je��!٢I:|!䆕v��8�<j���I�>|{��g�SYOW�m��Ì
����uQtQ�+��M�GÁ��t�#qU�H� �>��0Hc]*�=y�:�Xi�����RS/���5����n�H\P���l$�g�>a��m��l�#>\��>B"h�e�tj�:h�c]K�¾B�E�(�H|x���FWr�D^��3�,���{���v��〹@s�	
�lC8a�������|#�2�r�t���<�C�d�|��F<gܟb�?�`B���A�}����[��{͙7no�]+����j��z�CCb�F F $H�1T�V	H0� �������6�'��P̐z���'Ə�EU�X(�LN#�i��o���_Ce
���ŧ IL�Ѝ��j��w�\D[�r��W��Kr����;�.RG�á��׼�w�e�v(ǹ�n�>o�Uݍ*�< @���L�|��6`b�`�<j

���K�1E�X1������2B�kU����"_��6���Am�\�i�M�p�w��)V�QTj4�4#>.{c^Hwe�q�CN����r��9�]nj�**܂���%g[u5�v���M�h_i�u4��[�`��\;ni�̽����e�;�q�ύ3V�W]uʹ�6sis}N>=��of�㔘˷f��x�=���~����oٙͽ�ݟ���/�0��D;L�D�~e `�6S��	ɡ{D�k��i�l�t�HLj���3���h�e�Cs+G���|< $���dÉ�O:�YZ�x{~ܜ:#�;9mθj�|9���uZ�K6&��g��}��$���󖦕 �<�c ���  ���SDy�;�Ŗ��J'{v��~i*l�����ы,k5'L���B�u6��}K���" F����޾�徜3�c�nC	ׅi6 �|HEYYhJ"R*�+�+IX�V!�n��5�n���}�ꗪ�dm�%���τ�ZV���Ү��9���܏���y�|m�uN�����2Ʋ��<8��)z�tӜKu��� c�q�t�]� <7ޫE�vxW\���ܵD�*;��/���e�{����Kr�SR(q1��k�#}�{���Z�
�5��ZÍA),�jW���p vꚲ"ͤ� Ҳ()�Zo##�Hz�窱��N�n�)�����T��<^/g06��VB2(�D� *��"�`����$k�ޜM4�s�W��U4Y��!X�P�Aj��;���T�iҞ�f���7�ޘ߬z��!����n N���e����a�|�fr�쒳���xultw�y�M��K^gw���uT�^�[x��:����r�������V�p;�&����5S����޻���T������ubH�Y! ��P	�I"���9l�ڻ7}�m�  I m ȡm�   >����9��Wg>��;�����q�O�����;��֘��k��ѵ�z¢E���uI�t��S��L�,(A�P)]EDN,��w6y�Nͷ��y�K�gΎ���nH©-&n���l�f�-˔�����Y1O�}Lؘ���8�F���1�}{���h)E)���3��/y-H+n;�~>w¾&Q���D���-��ꯪ�R�y1�=c���?=��c� ֏iFe�g%��W��j����W��&g����/S�}��U���Ȉ��m���Ǐ��}�NiJ�Nur3,ʊ��s���u�.�z �V��+��\��z������ H؊�勷����zM�fEٴО��s$c]�X�5N�ۖ=�7B��73�foZ9D�Q���rd�u�Im��iaB��F��p�J�4�^2'53J�π�~~^voޱ�ޥj�7�����e����Gz����ٚ�ըu���I��� F���Zo{;��3��M恵dX�b��"�v�����TV(���(����E�b1Q�,EX�,������0gw�J:3����QT��_h�r��Sv*tWl���[h­��h˺W	����qm���iJ��.�ITܿVA���p��Z̛��ܳXI��[{|����Z�\@ �>�׹[T�$O$b�v������u+�*��O�2_��2uE-��c�뜌h�Շ~�^��'�B,�"�,d`���"0Q"��=��t�>63��+�Ћ���"�o�R�ў�+�j���돹�3�;.���}V� ���$�촞�6>�I ^r��z��3���V��J�a4��@)�S#n��d��<�=A���ަ ~�9�n�o������*�(>���D��*k�|7�';ڥM����PU����Eps=�ՏJ�N����_WMџ��ໍ�ǫaþ�:R��D;���D�Y��[O\��U��6�֣w��3�c��owl�7�/{�	}�j����/%���h�Y��.M����ՍS�[A8�	�(� 2�A�n�J�<H �RHRpx.�<�%���"*͙Eݢ`�r�y �m�
l_0��@�R��t���Ġs�R��v7�4m��p�p�	::ꨓ�>�i�����*҂0Z�W��eP�tE�~U���Bt�kN�PQuh7Xb�'��2���(�حm՘��
��FaE<�aɤ.�UM�l0bcQ�������d5��ѭ�jӸ[ӛ��2��C�&3���meue*���x�[���:.�zw�n{��x�L@[吣2�XKVS��r�љ���Y��]��#%o�r"�[�%��*VH�Ȧ�1,��Ab)�X�#N�ÉU�p�ㅽvk�.�&n�O@��h�(��A����ep¹�.ֆm��K�ski��Ε������syjV�b��V��p�X��й��%O����k?u＠4G`>��z� #���z�M�;0�Ś��ŻcHᴊ�c��9��\ʓ���x3\[c;
���G�gvm�}����L�[����'�F�Skq���p�m�����vg���sX��:�pR�M��;����#7)����0fS�9V�	H_h����P7c��ra#�ى���^w��j�������F��Z�ʃ��7��9����b�+6�9�gblժe���.Y]o�!x�˫|���ݥ[4��ڰ�{�KT6VG.CIL�L�6h�����y�[�Wt���>�ZԐX6QI��k��fV�KL������C�!��t�|��*��;�:��׃����9�D�w�)��C�%l�D'��+��՘^��?g+9�v��B9�A[]ȣ:���ݤ���!��zk�î�N kc��I��3��
'����]��sX9s�³�m�eV'�v�k��u����r�w6.���]-���*�S�Z��q�.��C;C�O����RC��	���è�H����0�a6��i��C�q���d��4�|2~�9段�͆2@w� V�����wXy���w����$&=�?B��j)8��{�ĚaX0����	�T�]P�I�@Yz�i'/�~�͡&�R�
�hL������m%B턬��	��	��`@�5HT�wz߿���\�퐟�{d:�L�l%��:l��I3�M��!�!$ ���~t�H��Bw[����zy�@<a&���A@��� u���Hu���@XC�~@=C�k��*u>@�	�f�ۈ��'�@5����ߵ�ֵ���\�?��ت`�a��&��BI������	1�ha/�'���XfB��4��@���G�I�2݀bN�ܤ����	��0�!0�����������$6��u���M�
�q���q	��>`q<I? v�I6�Y���f���� �=�!���o5�s[!<@�l��DD..�������5��8I�.��� X��]Z�J�x,z�ٗ��>��[��D�H6��"���wd��r��<�M�(�ƒ�!�0c�Y�h�#��\�[7}��#X���ɬ�|��g�eNϮV3g�G�}Q��\�o��͚��c��%����<0��5S�ْ#��Gg�#�M�m濲�=��l3�}Q��숋����;}�K� �(�W.yu&��Lف�)�r��/w;��dkz�O3Bw$�tNAN����M0w�M
��AH�n>����_]�P�-�/Ҩ<3-o���p=fO܎��7�{I%�e�$Y�n	^���xx2]���$mF��B�WPN�hTP%�sA��R�M��ߪ�P�#��fg��� ��R*�@`�2E�P�`���|EXk�8>����Yr䷑/޺ZT��vP�`�C;���ćNm���7l��j�S���b��I��|���UV��}�G�9�۬3mԮ�Z:"�_�`�T��GP������ڭ��+�Yp}t�t��寻|�yӈ��`�(�ɬ��Q��F�/�1��FڑjY�*�A�$iQ���b�l*�@I�LDI��w<����Y��ϼ}�g����=Z�&�r잉� �ٷL����S�3ܡT�$�!�d��fV�8K4�㾒=D��_x�Яз�tձ&4`�NK}!3S���r�3�/g�Mɐ����?B^k^�s��2嶾��3�3�e����=���̀��HB�ퟵ�y�u��4~��=�;�Xň5i`Db��E��Bԧ��fs������M�|    16�@   �-m� ���7��gS�+:��rE�Fn�ܘx��*Ȱ�B7�^i����]H���5�eĪ4\(�� �B� M	N6�S�Uf��*v���m�VY�J@�N[F[m �s<�}��3�:�5��M���Щ��ݯ�^;��������x9����hI����!�:�Ğ##n�N��Ή����~V�z�A�dg�D\�6��Y`=�io�>?~_�ݲ�#`��k���+�?���Ni[�Ֆ�V������=R�����-��n�:̐V�_U�~!�����Vi�� �X�H,R*Ȩ*�EA���A"�c�1B0� �y�y�������u�:��>kb�;,����5����c��H��$�:}�ǢI����2fEu��_(���FD�ybdi
��ӛ3��K��^�Q�}�l�$f�^��x�ҡ��7=��ݦ�poK�[�/�Tya��>��RL�ѝ~���ɉ�VeJ�OD{�����uM��)�h�""�舊o�)���^��-�*$��;���s�����B�M����o;���e��3h����;D+�C���	d乣���L�'1��w[}��w;��/bG_/��{��ɳ!ZgҦ���?:��q�9t�E[ZE�D���y�mb�G�	W>K�X��|? 4
s2�}���!�$}2�t�ͤx��;��!��Vkd�1��L�HR�LV�D�S���ۺ���s|���{�B������Y�w�y�}�}{�܋����W]}��t�DdU�X�"��aH����������u�5�9���熵��K򘉫Yw,�J^��̰�ΟyF�W��g��G�>4qO�W�R�?o���,��jM�sj%�}����w���ɇ�Tɏ+��p���o�e&����uM�f-�g�Z2�Jx�����,�H��g�J�dXΫ��l��*�%V%��]T =�b�$�c�����+u91�~�F�W(���*w�=�}�w˨�y��O9\`�[l��I6��C��L�d�%Y�0�[�U�9���ا��������Z�#w*�>�>���X}��b�G�oVzk�&�,yi{�rB���9�Σ��wŰf�y>�P�$[j
�Q�����#4[�a�>Y|>/Ɲ��-��>vDGk�\b�^q�Ui�R|b<�[	[�-���C��9ʕ$_W�S,��3�����}��5�������Iz�ǐ��>��Xj�˩�;x��6th_)Wknsw����;�P*�u]Jt���+��w:�#6-�Ӫ�W�R(]�k�ZW���~">� �" �NO�6K�/�P�RX����NDӘn�u_�P٩��^��t*�|(jЛUP]w�M���5|��A�1�菾8�%:��걳'e0sd���D@'��zffS��<�<tһ3^ti+�/�S�����b��A,ɂv׾�	�ҕ|��	�Bt��B��>qSm��.w�[i$�i$ۊNJ��`���N(�S����	�R��������Q4h`U��3�ӥ;K�����|��/i8:��7Ko����6Q|%�s���Rf=�d}���k��}�s���
�tE�׮�z�G*���<(,�\�j�䑳��{>�8�p��/*<��*�H�58�p[>k��0RuO�#��>��3��z��_���2�yY�Ih�"�Uf����wt�g�x���L�.i�b]m�eRb+`<��s9�^�׏M,�/�wJ����G�{˘�ӛ��wRqXȱ�"FA@�����[��������~g�y��}�8"����P*H,g�����H���`M=�\����}��*�۔�k�eX�xeocC��v�ZQ�k"�����H]��vnu�<�ߧ\�;��n�5�G�-�'s�;���u���Y�)�[k#¤�έ��)�������9Y3�A;kﾄ�;[>�Һ%��Ͷ�i4�m�u�%u"m�#I�	Q8�π��R�=/��U����NӣS������ޮ���VB�&�6��؞p��%/<�L�ic��ܮ�vs���JR_s������M�:�#��H�p���E��uA�P7��{A��^C9�zr�ѤԺ�/��kE�O�n��~7�|Bm)�V�L	�_}���3ގ/d�*.��X�sQEV.�:�Mg���vd�0�<�3o�,n�^㮩�b=���s0��K[u
�a�"=���*8���*��y��0}|>�sH���:�)h�HS��]=�c�!���Ȝ�}~Y��a+b��r�.�%}��@���"USi��i�E���V�*�2��u�Q�ȉj�e�*p��a��nc���j��X��\<�<���LyO�à����0P`������1A�J�"�Y`0V1F" � (�RAAd�1s�vϧ�{���E  �m[h �K� [h �ɷ�~}�~�׷}���eva��ՔH�%'8�s�W��^��ve#i�ޕbâ$�2�P.
(R+�U�Q�4U�)A0aBcS;s:k��A�@0��G���R� -��<�ns��se���ڛ\$Ji&��O���u�O��X��x��;k#�9U����E]ӌ�#���^��_�}�Б�5�^�ݻ
=����*�|�$�������ޕ������򬗍���I���+���较���S�R��}�h7��a�9��I1�[�p��p�̒�T�����nO��w3��(脭(�1�z�R~��M�!y�h���VN����=���D}q�{��_9S`�G����q�C)n��<0罦@�j��G��TE(�f��Y|��Ca꾭O�FIT9q�˞�(t�+�|i�#��N*��邓-NϑG4,�}��S�X�f��c�)nk�S�i���!�a)6u���A�8�&��ֳ��ǻD.u�eܾ\����w�H ������IT�$ �$�L&�yU4�o�2_��~矯��~疄4�E��#I��:��w�\�W�߷�ݧ#h��?}�_�5�^������ �XE�,ژ��S�/7 ǼƆYj���{9�������2�7�n=�ﾊ��E X,Y �^	�_/z�y|L�6��5"U�7�����`s���o^�^Va,��b���+V]�eRR�c�T���o}b�{r�����|ǫ��,s���S�w�]<�=O��k^=�[�A��Bt���=i���w�beNΧ����Si�G�G�!��O��D�L���K4<<g���?R��w�B7?<�n���x�;�鶛�4��/ݛ��rxo�ϯ�OYڵ��h{�1�%���(D�zT�o��̛�K^�W��]�zߵ��J���zx�X�|ĭ��f��u(
�~�F���%���%���Y!s���J�x����n��ͮ1��<�sK����s0*
���>�@���?sI�UUI[�	��b����S0��.E�}�}ܖ�#W�$ѝ��U�"+��@=�m���{pE�bQ�Eu�v7�1��8����*33]@O�5��?c�;��a��L�Ǽ�V/1d��>��� �"ݛ3��&�N�P��D�Y%a�({[8�|V�P��Q�Q̝�I���l@�4%T�Fׯ|%̛b.��Wj�<�	n��V���w�k�=ys$`�0��E�D��$F$�D1O5�y�2	^�t�}윩�hB�}(`��ص������$�,�
Ad"��
��v�;�^o��D
�,��J��I�c椝\���\�s��!��e�޽��C��a�����c��aW�ߏ<p~B�q=�<�a[aGן~��t�d����㶰�YT���輇�:���]ŕ5m�<ixf��D!��q��zOn�{�G�z�+#V`~��v������Zi��������S�x�"�dC��������a�di��۝>�n=�,r�����D@�yb}��r~1_\������5���4H����7�_�&]y� ˩S$��%�;p�ڌ��E�h�f� �5��>���Q1�@�_��YV\�h�^;�Q��Q��/��}�l���i�J�D���h��/�zn(ƒ��]����\��h�W���R�<�r2c�|Μ\u���p٥�{J�nLN��*8G�;��/�5Ѿ����k������s}�@��$EI TFF"@ PD� �������`��P)}�՞�w\��냦nbOY��������lM/m��#��s��3��nJ�`�~��[��O7Ώ��Y�m(�,�6�ڤ}|A�i�*�v�.�dC&u)�B�rt_7�s�Wjb��4��ک��/AZ���*�Q�
x>fw���ݠx��ˇS(������륺x�>�;s�������/i������=�^�}S$�㾥y���:�G_T4�,��꺝&y%Nc���^�B7}���x.K_��������3~ni���	�C3^ّn[��j�Xx��R��e�{>}����-�� ���7p��z#F?(���*�1E:�o����H���Q.�-5�蟸m)O:��K��.7��e����*��ϼ(Y��\q�qx�ڜ�>(7��=�58�I�XZ�oB7:S}��r��|�:R�k�Ny�7�./Ͷ�W�vP̮�S\>�NT@U��3���Z�w���d����O��l�׵*���s�]�8� n��x�R��k��J]F����T����k: ��?�{��U_u�|A:S�G*S��1&�i2���a��׫��+�l���:�mwO����g;��*�@��fKܝN�.N�\�|�ΩQћw|%�P^ 1�
z����c�I�ȫ��T���	$���s"��}��g{d����;����}�}G��:rѭ�F�ɥ�cT�c��\�Ν����t���:�Pp�B��;�w������r�Vf^�K���;\��<|�;�Qͬι�-r��6Y�
+C��Վ���K�:>�/��J?�����=�<2�j82��`�*Ƨ������{wB �՗Nh��}Iszr���-z��%[d[�-�U �U��}�m�x����JjX|,�f�����M���3�׮�Mi�b�0�[��yb����ϟ�)W�0���С�6f��[/.QuA�UAW�X�x��b�Q�2�+
  |@�1!�ګ�� E$G��,0��dBR�y�!O<�c��0�HH�4<�%i ��d"m��P�I���6�	l	����^wmx��JI+!��!$q$QRN�[b����"��L�z�}&���[�j0�A��b#E��9���͈�{�������q���y�a2E�Eb��ust
f���\*{fo�sw߼�f{��|���߹�      X��             �[m�$�K*ԅ���h� -�      ���  -��H   �PYm�    ����           7�p������_���3�^l�^���{��zV��S�[p`���W,0���hw��V1L�/Dα�@�X�j���Y�Q�pCۦ��\
�y�83�Z_$�4�iW2m	չ�	!�)�o������eu�ϸ]��U�jݻ�"os�ù��㠖�y%�?Y�گ��1�Evʚ������k�M^W�q��mbȼZ�3�$r���lS����}�惇�$�_:��V��-wك:�'�"=�g�}w�����(h:����;joj������N���Sx�e�gv�_j3L��C���ܱ��J��s��9Z�Q۸��9�D�ٗG\�IŁ.tM	���U�U�R|��X���.�V���b�Ȫ}J������IwAU��'j�7lsDiӦ�L��o;ۺ���;��3F�E�U��J�I�+�������9X>M����-�&����e-�[�����d*�Q�A@ѭ�(\6i��%�$0�ɵ�	�F�{Zn�8��#���Ҋ*RJݎ��@�m0��n2ErG�ڨ�W��.���ףV}9U�-DӶ$�M5RA9�(�F�,�
�.�8AL$�ڠ�鷚)�VGQ�J�wP�p�sz\(�N;ȩ��%yQ���P���^&��
,�NK�M���uD(E�L�uRS�y�TY�f2�tEK���U^��ja���l�]�F┍���{[t�u�3ԞPtA	Ro�@5i�=��\���w�w�s��m� I*�  [h[h   ���}�/���翻��z߯�˱��7�H�뾉���s4�z�^�ٰ�V፵ !#q��h&`�!��ʁ��	���������L�o%m�}��9�$ ��}w.���Ħn-�v6�O�g����2����đ�B�����R�>�77��%�
�"�&YA�m�t(8k�D3��X������n�:�Q�|�l�%�$^a��|R�}�o%�J�|����j�1l{9�rߣZ�� �0��.xٻw�w��]�T 0�S�),Wj�zz�r+���W�[�&�˯���ŷ��j�P��r�:�g����]�7J���#�U�I���b,);�7�	�+���;���<z�������h6�V����R%��/�2���Z��. �*��gq�#"gdL{:H������a+���+"�",D"*����>�g3��=9�o�Q������ֺ��K=�����<�tc���[�F�4 ����8X}�}�َ�^�ce�1?iB��k�5����|�M'YG�,��h�-��m��m�Cs;�Ī��2�J&���BxQ�(8��k(N��<lT�I��v/��h{�M;�R�ӧ�z-]j�R)���s�~?M�i�4o���a>��@�˯������|!7��Δ�}�T� 3����*��1���e�Zf�R�K��i�*�Q� CFg|֔`��h�7z�1��L�d�A��DY��W���O���T�wzwIW
<N0x�a����+m?4����>�~}���2�`�{�	���[ֻ�dpR ��Ӛ���F�M��پ��@������ni������G,�w�2�9`��#�C>e��y9��mu�(KD�_��Y	v�+�qe=/ƃ7��]�7/菶>ܸtx.&,�����t�P��^ž'c�%�I��wc���c�����a�&"����.�1���������:,tu��u��L���HG9�>��>�,�����\#��j���̧F�ٟ0���rI6�E��5�:j�*온8@�!��a&�:�(=R�P��v�B��tЏF\��Kn�{������gd�;������>���ϵ�B<����/ɏU�p|��9���~)��7���"�-����z�{l��ٳ]��1�]$��W���l9g��zfw�x�ŕv��'r}�S}�8>3�ٸx�r*�Mu���Pp�o�K�{���)�K\�Еq�^t��Uܠ�5�AA �^��bٺ�:���xk��V.�R�g=��]�����2#&z�7�ML�M@]y�	�z 0��/]�D�� v���S�̮���n�t��7ȴ<��}�ݿ@���	������Hܵ���|���h��ՠ6�c�hG{w�k��\��'F�b��U���L���b�O9��Z�"1v�8E�&�<�]!U���1M�E�g 4A�D�kv���p2�D��GN���HI�������v�y2�Y��4�t�⚝��30��p�ceqK��;����j~�'xD  ��)�S쫖����o���=�>��N��x���ꃢ,D���aˋ��9����yyз�<\"b�w��G��X'�ϩ��U������q?�nBT�৷�|��WUt�;�������\&Lz�2QëQi��ܳ�Q\t��*�;�Ɂkn;*�g�U^h(�s���Y�S��_�V��vK�҃;���mb��jÅ"�����x�$r,��ہ�+5��w�-��<�t�M�$��|#���2�l�
�F�(�o�]Q)�Y_���߳{�Nϓb��+(����Ӈy��/�ֻ��CR�y�y�Yu)��ѝ	Q��o([��jq9�Z^�ݨ:�[7WT�LQ��;�[�z-$�1�k���RJ��Q8,�9������y�F��O�)��'���C���9��"�_j��BP��Mפ�K�e�b���w��/���H$��$�����M�f� �T2�e�����x�߽�Em@�\n�`y�I��0P �Uv�B{�@z�᜿T�nmT����a���ַL�"i8��hS=ٰ�# �_��n@���Bva��N�Q~�zh@�z����Kّ�,G�D�lvt���FM7���P0�+���x��[��4>����j��k7$��&��.T�qQ�0�Q��yk����:gs�XC�w��}�%�� DD!�28Ӯ�>��ӧyV�`�Lϰ)�<�"c�!6w���S�z�z/#�^�7���K�m�k�T�ٰ�q��a�͛�Whu3DGQC�]�E,B�8	hج߄{M�7u���u����
f@�\��1u�Ⱥ�"L��1Ҵ��.���e��ڦbF8����>�݊kw��g/�1��f�l�EV�U d�
���sg}�{��g��Z��q�7�FcC�����  A��O���=UĮ�綿]I$���  ��  -�ŠI-� �vg�w>�Ц�'��t��{��'X���>ˇeŗ��z�SGl�f�<r}e[�3Wf�t���(¢d�.�ضH�CEn8i�-�J����Y-���E���˖e��v�ͅ� [��v���pӂ�,�d|���
�P��#�}Hq��UyB}�Ζ�4�E�i�9�j`�ޟO?m�٢��( 5�ר�bѓ�9��*�"*=��)�E؁k��;'�Z.�}�e���G��w�����BIi&�TҠV�u���=7��]ߝ��.��I��W��5���}=9o}2!�X(�''�X�Gןl#���FE��D@�}E]0�V]$��v�v5���ӌ�ʅ�Q�Vx���W�j�.�f��b���K��HC�c���OY�y��Q��V���1�({��չA��3]��/�\�pBK�ʛ_�s�Q��w	"]�zP�֥yܚf3;�������R����<�ޡ]��^bS����[�J����V���ػ�7�U���BG�o���^8�ݳ�J�[�;9�
�����zݭ�{��I6�m��}+ڐ��\!��p�[m$϶�9�a��>�R"{��>�����y�êl}�٘�iP�|���}�dĆe�{�z����)�'�R�s1�c�3F�ӎxEO�o�]�V��r�;����~>1��H�*��Iߵ毚�9U,.X<դ��9�9�NS�fr\� ���(���8�T�/"dG��J��ћIM�[5Y�=�9�ϩ�>*��Y��x�ژ�5	ho), �0	�=�$�>��{��Y5���)|�������NIV�T�y]xf`���k-�����m���'�����3����<ۊ�Ҫǝƛ�8��t-9Z�w��/�#��ѐa���.�Ϩ{5��Sxv/��9��38����pj����g�\�X�"1}�.w�-eI�e]>������)����s�kG*};G�{h�94�f�Y���}��F�ȑ�A�8WAX��C�e�j����^��N�������_%�D�x.+� ;m��ݏ�.ł	$��혚�r�����(�$��>9��jjsj}4*�4Mu��^���{����#�K���qS�l؛�����[^Ζ�JB�Eťh�~ʃѲ�n���������O�Nz���b"��b"�]O������c���5uO�m���{�}'7�����qT8ʗ�$�y^x��oцT��"j��Ӧ�����-�E�3����H��,,�a��5{�}��;��Sת����q�����vu�[�U�<�|��Ԍr�!u�p��������&1��,!�4�^�����u��9S��S���PSc1*�?{�O=�͹
o���>���Ǽ4����s=:#J"�
�1�YQ��p���3u}m��%�_�m�K���GN;�([�D���;;��T��W�`����5@}�	���=�`YB�L���܃C0�P�U��~t0����~�"�m�c��Vq�M�UY>����������@W}��m�L�_��l��m��G�Fa^�����	�b���n�?g:3	�ΟB0��6�/O��S�[�է�)�Y�1 ^7UKjV�����z��4ɉ��.����l�>���������k��ǧ�OT�YO��Z.jW�e����a��ٛ!dÂ��׍M������PUF�z��Vs6ղ�Kjx�J@od��l�r���?GШ��NAyIU9�>�Q�.�:9p�y���[:���s�V9x�l*�Ib�1�>�)d'T(fg�G�LUM�(Ut����mx�P<=����E
�K���1��l�'���=]�~��8�i #TNZ�#A��1V��
@R
@���`�YD����N4r�^�Ъ�&�g�9��oK�=��SZ�>8v�ګ����W<D��R[KN`ko���G1q�c�-py�s���(#Ъr�KSwa])�-�եe޳���Q��~T �B�"ă���[ih� ���UT���c��z�z�Q�����c��7-�Km��m�\*�+�A������8�]�������7��9?2���kC�n������3�\#����`K�9�l���;�{���dDDP�3§���m*5H�NK#+��v2��;����`��c��Y=��s�%r{x�Y_$]Z3I�1(Q�M.����r�U�x�i��f4V��sc:>��ѵ3�L#2N~�W�����3�W���7�Őy7�Uq).t��z���¤B�Z7�陵է_�2�Ui^��@G�"/��B���7��~�| ���e���{����J�R���>
����&���]_�x�< �yGO��N0u��o�GF{�b�֏�X1���Ԣ���QC�����}��-�-��Z�bNy*���ů%#����X�o�Q��zi�Jh�q| | H"<I>@���vSͤ���I$�@  �m��� [h]@�@ >^_7�S�3�R�[�իP��՚��+�X�S�읯5Y���+.�(�v�e֮o�-���j�e��iߴ�
J%���59Q�Q�؟J�V��͜��y-�Y�Fl˿��ɖk���>��N엽/C��r�ק膃���H4���5nx
!bA�&D��k�� Oe�׸D��QS>W-]��}����^��Ss"6(�w�f�qTqf�ȱ�[�;���8��8\��߆^.�N5l��+'�t��S焪��{�������=���˔+�K�`Li�zd�95����6������*ۍK��ʄ�׌y}���oJă���Է\������S1���W��	�da>�vb"0{��i�;̥�v;�@���KNO���5sA�?x�S�M��53P����W*��0�����;����i��
����w������x��;E���ya���Ϭ���̪�W����6��i�'9xv����r~��6u� =���H��H�rB��,�v-"E�e�*��RVR���mۦ����y)�{}�L��t+^�s�T9=�R|c���FutR���1����@QY���3#��32�y_�(��VeP�Bu�&DQ�k�8YC����/�lEC��8lw3��eE��C��j�؍q�ӧ[;!w
�b��efӔ�]���xi�����v�̘����	�*S�G���ߝWk��֟�\���ޞ�ٚ�>�*�w���,�J����(	Z)���9Ii��M)V �������_�k�Nz�"��!?����~>���q�A�ʜeb�5<+GT�Y��{��fP�c%�Z������`;����o�����t{�#u4��5{��?r�p�,��}�D����J�`t!mޮ���N����DbB},^�g��5R��j,�*�<G���ܜ�*�v�1�D�7MF��S4�m>;�	E_��8�b���{ޭ�rD��6ܒ�'���$�-�f.N\�39�NQ^�X0]�S�j�1��:�e6�k�6)o5��Ɣ#�܎����1�[��q�hV
��>�N��K-��ڙE���B����P�g*á: ^^�^�zx��g)9dϱ�r}�V34���/�zF?���#׎�E�[Ȱe���re�&�_.v��k��.=�>�~w��H�""HdU9�ܾ~��]����ow�}��8���kp�d4��9
*��-q;ϦV�/6vH����;��V����3{�w�}�����jo0���%�H9�%`�P<%�ȳ���g.1Ѿi�㲺�ĠpV"J4z'c��L2 h��f	x��n	�1v��&��i1�X,��/h���NAH|��u4Ģ�𼗹quY�};(r�WT���a̸u�͆u�GS��# N&K��n$e�i��~�"8�A`�� �$�I�`�PW�����$��n��"��n�)��n���^��&�t�9���k�%�'N�܆;(<yGi��f8�a�t%���w��.X*�eP+���9�:3L��}����BЯY�-�3l��{��0w������X�,��	4�`�
hF�%eY�q���/'+*7oR�NZAA ���5���0̨��:̂�����m�՗Zɻ��U�W\��)�'熈�V�Di ��"y��z�"%@�2�@(�L	�f��}�GZ*�|�l����X��een�)�c}ۏ����n��z�s��:��3�I��]-ʷ¤,���%DAY���:��4��M�*��ɜ�7/�yϖ>�ެ��f�t���ve=��{Cr�ٜ��©s��QQu�'g+�+�2���k�
��r�(m�����k�{o��T��ظJw�:��+�.V�Kr_+�=u�m�vRp��uͶ�8��fW������lk�w�s�ܒX����`�u��ėʯ*pU���쫲vM]�t}�]>��4���@ �+ ��OM��w[*!�F�-��l��DZ��x�t4:X�ڧݳ��@��Lc��Զ'4u�d؇]" c���:"_Y윢���*���L.�巡�"�oS��Z�f�ԱK��0 B=��,���C-\�a�����̷+�Ν\k�L�ҢCM�Y5�Tz�k�i�3��7o�;�6�=6kޢh�e�C���ժ���4o9#)�!�s[��7���#���zt��Z��vR���DE�$�3��f3}��dre��b6��ϋǠ=%���S)�{78S���)5�O4��WJroB�r�Q�t���U	��ý�1�W���8vmn0��%<�����}����r�m.�[7�n<#Fܣޫ�C��[�QHw�*ͭ�t��i�/�Q��x��x���(ֳ��5��9���n�0�w��'M��99UNg6Su^�K�w)
Qϳ$�R�U���1'Fn����}���y��m���~{ÿ~��4( ��Ad#b�1�;o��M}}�~�@�5`ߑQi%L��M�^$��M�)�a�����y�%T�mb��&w�sДXў��Z�i~�|N�M��eE��S�ť>����~Sn�.r�_j;��!����P�Ad^�|��4m�W(���8����×#^+|k�z�W���j��+�{m���2�wRR�6-�"">�������ތj��>�����D��9��e+�b}x����;�ٍ����}Cgbt*x]�CO|1?c�,cھvƷ_l�y�zu�Z�1���f�M�k���^}��b㍥��Z'�-��|!�t�-��ulz<��f~�^>ޟM5�n�|�Ӌ�@DP��kyc��u,�NMAL�n�[�Oz���Sv��ނ�,�F%�{�����k^\ܗ[q��u�:����c�����d9Xn���x����@��'��<8��3��|������G`�2m-���m-꣏���p&f��Vw͈�6�糛m$�i%$[j]�~B��-TbDnA�MT|<督sh���R)���Eި�?}G�[�q�z�^�ՏS����~x��N�6��
@D�6�ٔ��KpU�(/g^����B}�%ӗ9;\ ���`{>{�/{�O�J�_{*_lJ�P[�Zi���k�|EN��Z
���E��Y����6ʴ�!�՟{���0�y˾����l̺�R��1��+�{�i������l�R���9��#UyaH���W
�3ݽ�ұ��-&�N�l�"��o�ά���U�Of�b'�#��S�ě�M�c��`�D��I Y5��߼֮��{�g�ې�I�5��w���;��mE]�V4�:��=��j��<��xF�~�f�@�w�v��.�<'�|v�� fnnfo��.��w���g� �� n��  ��@   �����;쫯N�
�g+:�/�R�S��1�Ɩ�4���o��s�� U�����O��˄dK�I:���AB��!E'ҘZ���L*)�tOӦo�Y�mC�����dU����{U����\�� ��6�-��N����z���h�����'�Q����M��8��f\��|����Ϻ�<VZ�Tj��2U�դ�^Wl�L�$	K3�d�<�g��09�#��x@�} ���U*�'��՗�Z"�4��v�$:�b\5ޓ����{�ʆ[!�UC<n޼���{�+�q9c$y�	L��TsCN�U����w��YS�]���=M<�Ju@�FyN���h���J�|�Q��z��F�˗jrMN+�J��Y�n�X0�\�(�9XU�W�ܓ�!Ȉ����m��~U>�� �aɟ�/`�{������O3D�.\��6J��VL����
raNuss���!Gp�uY��F�-&�ֲ�i�����x�g6�-$�m�Xi��H�#`�T�H<V%T��Vd?��`p�����^^<sӹ��v�� '4y��r)z�*��.��J��z��B*��M
 h���o��㾦���{�S�>[A`� 7�:��(�_�RD>�>�/3��ԙ�Z��WC�s�S@ӊ���Sy]	!�VZ����1�5V):��Rʧ+A��R�Qy#��wT�F7efn�j5�=W��%I`���+\��UGYU����2Z���M6��1���~&���%�z-:�uKG�1�*H
=��;��yzs�^��� ���G�&*�V����k��z��[��"P������p�����l�b�9�NI����%�&U�e�wç��[�C'�uÀ��<��F�g�9Ზqr�Y>��z���-���ڔ��0՟!z�~��{��#��tG����:�b��q��������]g{Q���|�n��(�M�Uׯlz�Km��m��<�%�p ��M�Bd��f�#�Rb�a��f(S��:�@�6ec��®\���|��������@D �R��I1<������o��混����$��[*D�3Q���y��0i`����
����X*�&<��ē�����ӨQ�ٯ���_7V��@�!Z�,I �2�mU�^���s߱�J�<���J�S¦\��ζ��rgǪ�.�ݗ=���3��Km`�DaU�eB�[j+A@k*��kPPbDiab�bŅ+K�����b� e �"B�!f~5^3����{'K�<�7�`pХA$�m�`�f�X�;] j�QX��q�l�s���Pf���F#��r}�׵��^߽,z�{��V?��3ӡ��t}{��j�l}�6�z�x�@UJEg�� �-S�"�s#� /�c`�r���`轶�wO}�+H�����+�B���2�k�=�0fA"bDw�n�m�$n�4��tc���}�G�&�r�G���wb�O�^kX}X�;��w��|�$ �=}���x@2�I�s2�\�f���%%�韩�U��W C}�G�3�r7_����{���6h#�u�Կb[���� ^r'׻_T��7uN�D���h 'U�W\�m��¡��=$�T���h=�H�/j���b0=oܥ��]Q��y�A�4�\���=V>�Xi9���݉��:��S��>v���/k[v����
<�r�Mg�5���<�w}�o=���Z��o�G|�~׭{��8E����ol�i\1γS7�J�|�?�)-��3��g������q\�y�`�YI�zw�Ezr�� G�
Xd��]_%y�w<�y|o�/mY閻�l��"�eQO��R-�i]�_b�t0�b���-�%�P��+�}G�髌�Yn�.ѣ[��^��T#�a^�=uF��*}����x3��Dp�;xB��S�h�[~����`l�u�">�����6܌�t����4�	�!$�4Z��>��,���r�Mȴ���c zykY�Gݫf��
}Ɵ��f�[�#|���({9�:6��KЛ�ܦD��L9}[1�*�XÒ@չ�f�[[�o�6��)P�u�:�u���s�Ie�����]��Y!�{V��JA֍����>��ᢇz���V�~�DHH,� ��0���ut���@ �+��tZT�}=�ј��Q2���7ҝ��/�A&
^��Lx���]��ףgl��~�{ڟ�(���Z:=~|����}�����P;_�3x��Iw�-ر�g5<��m�h)�bP��ry�=A�3���Jd��R�ܕ����/Cߔ�P�߱���������_}��Jw��
��_�=.��~.��[���^N����p �Œ/�D�R�*�A��2AOxQ��#Ԗj~͕w��$�$� [h�� �m��@ K���E�g4�'F�/;9���BZJ��U\ɇ���#�
�X����QPa"\�N��0T!d��ŤѠI)�����t��" m�Y05�d�8-�-������*jI���!�۞NiPC�f�����a�\�ѝy8��T����{�~�RW�x���&�Fd�O$kYw���͢;=��.@�T=�x.X�x�m��Ŋ�GNŹ�n�@����_H7lG�R��S��In���<$��ȟ_b��0_>sN����	�d�y��:��O����KYb�=�7��kp帕P��[InُY�Um������!۷�6�ffH�iL�S�����ߤNp��5�J2v��S�,�D��*��W�+Ҏy���!��Ǣw��ߠ(xs0ht��A�������6\_�����O=������t������$X����E0PT��8~��ns�_}k_S���7�g��(�	����bN�k�7��������7ys�a��ɐ��-��ܳޕ�m&&��ҸRf_	��`m�kV��O������1f{��1��[f��Q��0�H]��i��e�J3"&چ�}+4��_����~�}l���RH/�|�(�
�T�Y�<.Mx>0Iպ��Z��)3�j挎3���]�k*�ow%�P;�l#1��p�Ō�[Kb��DZ��hG�=V��p����5�ȝ�l�W��%M`)��̧���}�����PE�n�͘��_cs��˳*�Q��5ڧ�<���){��o���k�"Z��_��{+�1�a���3�J��-�+�o�>�'t��ٶF����l])uWalǟq��pĳ"���u�絆��!? @��	����4sé�|�8�V�#��^]>��}�l$E���x�[�f�t{S���=��͙�|��g���-� 7��wa��D���R�Iۘ�ļ�<Q�0���E��#�}7ꜰfi14nHS�u�x@UO.�������+C;vHS�z�Brm٦b���t!�Z�˳�{�f!�|`]9[P��W�� ?X���e��N�Nⷊ�fg�p���s���~��.т��]q�4CN���`HG)Q���3�Q��+�O�s�7K�zʺ��+���o8�S\݄�����<�"��0�nn�J�2e(�a�u�*>;�u��;�g_%>�C=�ʶ;^	�Sܳ������Tu`�����-���X���p��o(V1�������՘�k�Gz���p�Af:Ο�)�/�#�s�$���}�&�XF��M֤c��3�-�b���A[��4Kh:]�/+
�y3�5Y���������^��!�jUV%E�6}G�2�օ�����i$�i$؊L#!��F�tI���&���ټDF�y�D�f�߄o�4���,��v�u_����UwK�=���C�Z*n�IWB�uҒl�430�DG����YS�Ώ/��W��Ҫ�l!"O,�l��<�:�7_݄��fwH��I��R�#G���k���l���4+���_`J~�DY>����~�_-g���e{1�w����B@�����gPQ�ˬ�N�)��F�Q�Z�^j���T���rq���/&���;_mf%�`�'���<���}��){��isf���"�|�!4>�Rty�[s/!�ˬ�����0�����Cp銺�>���'j�#Ӫ����ˎ�r��?z�H���9��z��z�h#V�'^/����\�G'��{"=�ӓy��H},T�2I���+�e�q�{�+��9�O�Ct��<��8ݟE�d��A�����Q!mj�W@u�	��T�#>�M��h|��{DtlE���_�$a����>�)Wc��>� #��A����5p��Mq�V�l��/3�۵]���������;��e:¥���-#!�G�2��ZQn�������C��*nn�}�G+�m�m�n��4��5'�����Qm_��;�[ʒ�^[T`�V;x�1[��<7(���_r���>�jr�^��;���� D1s��6��2s�n�V�2,���2mH��:;:p|��!�zE���jw^V����*�Y\Z�m7}����A G�fs�!��
;{�F۞˷{���md�t��d� ���ě����:�5#k:����q��r'�Oqņ�nk�E�
pJǹ�\��y��Թ�Cךp��S��ӥ���b�������v�.�2�TH.K�"�b�ԗQت��1�H|O��z76����>�ݦ�h۱��xñ�3=귘M�W���J�w�+k(���M������ko��{�`O�U�ik��*�ʕ�A 3�"�Ke2җ��D-*&X#�}�9��l�v�b5����M9j�@��d� >$�ȥ5���`���<s;��-uhc1�Z�Av�)� �{у�FcK�(�%U�b�.�=�(K�(A�̪^�d�*21���iB�F�藒P���*F�]�bsW5B�o2�>tB$��r�37ʊK�A ����6q�m�`��c4ƗI�hb�����P������7�ބ������f�a�
	�u���S��Gr�5u�I5Y{�ʨщts��x��3�t��hPO�)e<�R       2j[@ -�            �M�,��-�h�m[@          dI([h   ,�[��m    ��mH�           ���Q�֪�����5fa� ra<e��cc@�Ћ�t[�K�E����/*�{,���7�̲�t�F�/;I�}]%u��qG���-��:)�^�]���uI�RH��[V�$�k�$JV��ב�w���wN�kz%غ�>�\ۦ�8��w Ő��;�v�?�vg-�6qc_֬>�C.m����}C<���n.S"D�׆�=0dW��.�����;�&��Mv��Ǩ�F�M�|�dֵ��q&�:2��m�+$@�Z�BP{������9����{��n��A����� ���.O�v6�* ���b��(�}��z	J��'��A�� �� �O2v�b��1�%i<��Si��=X�,`�A�8.�/�v��jT׮���:Y������9wc��$��N��SU\�E����-�i��,	ut�fvR�9�}Օ��Z�R6�
�U4ye#I��J[i�E2K4��[����f��.��M�b0e�%�E@�(B�X�y)���K� A�A�);�*
2������e�اD��"e��b�(����Xl"AY�2�PuDI�N$��Iܔe�MhawF�h8Z{�,�9�!�Y��E�S@��-��=veæz,��� ��7�H(h1c�HI���AҲHgpd,�;sJt�c(eB)K��ֳ���� 4�lXje�?�����W�d�Vf�۵@@  �[@  Ԁ�������}/�fl������юt�Q�xgJ	^�L�Y�{Pf�i=��&��z�:w���#��"��Adh�Tp��qJa6�Z���.��������79����I��Vh�����Q�ԪT�BX��&$���zK�~~�~�&0� �=��� ��tV_#�O�z'+v�Y�q�P��t���{�)�U�}�la^��s��K�.�4:Z�e��jrr,�U;Ǭ$�J�19:���F/Ew9"�_#�]��Oaޫ�f�p���<��k ��J+g�p�ܗ���]_Y�'4��m����KvJ8G�/����,����\���jQ�ޔ#�}��JⲔ�h�sӂ|�]GX�d�?1R|qC=�}\�Ŧ��z���Vxݳ_|i']$B>A�-�[�Q���=��ǔ�-����)]�伃��x�����P�-�uS�_j1s����Ŭ�ٙ����$-[i�����:9b�08i [�-�ۀ�̅�4MG��zh�:ˉ=~V"j���nl���7��,�&�sӂ�Y�1nVA�q�xB˧g7��i��U��� ?#i?ޭ=����߽�5t�t�4"1 �X����edI�ˌ7 ind�����qi�]�-�Jop��Ķ;9�hիQ�5�o���8o���Tz!Dmo��-��ǖk��|>�2���2�˜�eo@�תщS�s"�o׃���gvy���=Ǝ������x�y��(��B,�,���ޞ�E���/�~槷��^Fѿ;�*��[(��Vzh��h1�Kɟ]0����9����v#�1�-����3���1m�?�7��YK�����T��i誷�����\���Pgo�=���˞��C�QV��b&�n'"��X� NdK�X{=YQo��� '�,T�I���C� ���H�T�I��JBz����sI�&�%�h����L�Ǜ�G�ٱG��bar��,�Jz�Mf�l���9�e<�#.5 �Ռ��G�:���D��&}EЀ#���K��9��8�͠�UJ�o�D��gB+Ng�K�Y�q<;����>v��*+zz|�9��I��uۂ<3�|W�6@�Ж�Ruj���P&eI�Lق�B����G����E�d6��
s�&��M�z��uԘ��ӝD*�z�Ɖ.ʀ
�:)����=��D�Aat��s����VSJ<(^�ۻ�6l�vxw��!�g[�n�m�Οg���h��+
�+R.��/�*uߩ`���K��z�������k�w��կm���f���S
u� X����aN��k�Ј�����s׊ws�b���>��7s��wC�����'�(b�5Nm� +�_��H ^^g�r3�';��D�"�i�\<����.�dѲ�1Z��WoՍ�M�������W�v��G٩�#1B;�VEZ��0��L8Z�jt��ݮ�������MU�,���˅�輂����ϴ��]R��G�����$�d���=9������w�wW�K&U�Q��g��+N�ۏY<m�W�$�����V��?#|r��0P�҅@�;�ڡnr�</O:\�|�Mʿ�L]z^��ϕ����o�3txG���5�M\���}�\p6��=1�^�>־�]y�O�(��"�
� � ����C���\�{O��s�l����w8S�%P�렷�r���e�3:�k�gG\`��1T��d��v��@R�b6�n�{�e5�)��a�������@'�z��b I3�s�t��
�Gg�J9om�gt�Mb����58mDYO��a�*3�E�cl܍�!9���Р�D\q��T�B%)����?�c�g��������v�"��+��W����k?z�c�8���~b2V�=%;4�=$re��S��k��^��B�DD1{x�ۖ����>�Ύ�������D@�Ǎ���Lσɤ��v9�	Ӌ��6��󓢍a�r*G�eF=E���Ք���X���لfԾ��f���:�C�{�C���3@��4��9�r*�r	PSfT�VFo��۝�����b���}E�[��]����;�N�`AR��Z~� ������Nn���M�+��E�_�ߔk3�B��r�vGX�Fe^!���U��0۬.�����g4W�����6������NDFH�A RX

?y����o�<�   3v�@   �   ���{��o9�|�f�����{��
��]펝)s9���ƛ�$e��H��92�Y�@Մ��S�-�DV�5
"���T�N�+ԽL�!�s�����+w|g���q�[h �y���\e�}��"�)��7�I��F��χ�X����Xd��p�7�8X6��5�h��(C�q8�f鯤Z�lK��jeZ8Lʫ=����������G�Ccfq�cֳfwE39�5�ld�U�j��L�yҁޡ����n�:N��}X�)�� �ta��l<���tv�厣���N������6���:��A"��]��P��	�l�H��=)A���MN���&�|~tdJ<}zݠ,�Ç|1����)Ƹ�{ݯ�귶�����z�^3$I����P9Gݦ��u��d�R�����i�8���ь�{��ov����C:���0B��UO�H���ϼ�w�[b�D��2�|�۽��13��pU!5��� �Aս��i�E.��ɺPb)u���b���Z�}��w����|���X� ���5;���yI�-�^�3���:�Q�>'�7�9v��� I��(�, ��H���*�� �x�p�E�%��]�hԳ܌ͻ��Kzo�.Lr�!۾��C�k��\���/bz�"��W���gj���������9�[U�/9�gl�r�e���;���i�Z'�"��J���/Ok�\���W�֊	���I�u�T���[��K6tD�f:	p���%Gu[z'�L[�=�����}Q�L���C�Ⱁ�iXUJ��T*6r��6m���������ͅsw\�[��̢��������\u��C 䶦�wg�g�j�g��F�L��IH�ts)�4���TǺ
��v�m ��>��'3Ɍ�6͏�R��m�U�o��(�1�x�mj�W+��?��s��.����T������.�[�j���qь�I�"%�I�=Ri�rx�ʄ8`ڛq���)�p�ٙJx�����P�>�j�e��0�nzc� �w�� И��s�}�OI��4�uə*�|l-55�TcAG럙;��,�����N�E�4�0�"H3u�O��(߄Mb�A�۰xZ�蠕Ĥ�U^N��c.�Ci�À�Z�ayS�u�rw����72N̰L�-�l������{� �}9�Ë��E���Dm��#�jQY���T<,[��R��RŽ��>����T��VM���&RQ,���8�nk&*�w-�	X��p]	~Q����L�;��,�	G��.ĳ5}������3����]�W�S�"wb>h�6�-6�/��������\�]�OҦڭ��(w
y2>�{�<�� Dw��N}�7�"p�Lv���<�@c#�z3�B�������)���n�k֭y�L�ir_dUه�v���V~�.�z���Z,{6nX�r��Wi�;cf������uo��G9�Y5�_���G���KN��W�~Q��G���&��eN�/)�=B&@�d	��eo���x��B4�fY�b-�� �FkINK���Q�'DI��[=�1��2=����H	Y�⦅%`�*c�=�I�>�<|a:�"���L�g�n�|�g��.�S���ft���F�z!�[#��ΡS�P����8�*��.:A�]�3�y,������:�XS2����V%�ѝ�n��m�pe�S�+�Q�n��n���9I4��Xk���
��<�#DG�w���$��)$ǽ]�g5{x�]�n�M`�5>��`�}��H�}&$�x��Ÿ���'��vsj��y,;�S�?H�q˅xT_f""}Yh��뽪�'�Os��]t�u�ag�b���R�|t��2��Ӌ+��c��QXs�t�^�}ՙ�j*�+�M�#�o�6�eM��6v�H��v���f���	�g1p;������ *A��3�e��~�+� `����0��o��Y=�4��m���y>�Q2S��p�V�ƔX��ý� }E��u�} �1���z���ĬX�U�_q��f�8�`�M���dc�x;n"]�I_W�Y/��_�sˌs
�R�������EX=׏�S^����Ϗ���<x��O��WǮm���ql�&��������=��o�K�-H  Ȋ  ,�  m }}י���=���[S�v3��l>���E�M�վ�&T�����Л���լq�P@�(GM��fӅ*-�l�P�9J��E�@ےE�t�qH޲6�b{�ux$����s��K_n�"��0`&�K��6=�r&��NG��C�c�G2�}y?b�A3rn�H��yB.H����D�X^sQ�mޙ�sΝ�.K�]�Z_q��Dⳓ�i/��ly3����0�^�d�v���Ǫ��M�`�d�{X���Ӟ_B,v�s\�nW�������h(���cj; ���d'����XO����wV�C�q��o��2[����
�9N�5���;�3/g��o��L�XHf����0rGY������Dg��>ӫ��� K��r��6�+���P��d�D�vg�h M#���E\�વ^/^�Ϩ����<]���y�'��wl���m��m�]R��I2a��&��N��7���HW�g�Z�z� �V*o�\�b���{����L8S���0.6$�;րx�����S���V�U�M6�h��eݯp�v'���ҏ��E��H[`{�̻�����z�[s��=�N��*�Z�U��w�;
o_u�8��A��|ڇ;/����6v3V�]�\��1ǜ��0�'�����
ȣ 
#|�}:����[�v������V蹩^ߤ1}"��mBu��Qy�~@�G��H�6�{n����Wm�����X��]-�խ�>�	� 4��}�M�^�V=2M<�vE�be9��l�΅�'�!�r�N*���N�\��W�P�Vjθ 	{}��S�x��NFF�.�ĭ�=I��	ƷxT�C�D�4������J��IO����'��'9��I��i%s¨���&f��3VY��%�37�o���~�ܒf�B4��'%[�k�>�����=S����'9�Pw�(1�)1�����v+�4��t��-��W#����"X�ԫv+k" �{k#�9#%���R���~�J��iR"l!�+�bf��+T����s���s���K�A�ts��\��S�Aܨ �*u̇�Պܭ���}yX�f3�]7$��@jcf���+73�>Lt�-vt4۱���^�+n�6b�fg	[OZ�\"P˂��0×��v�6t���fB�1�k�D#d~Cb�5���m�aeRmQ�@�f��^bg��)h��������9^A��� C`��bQN�,��,���&"�[w��)� �@��۶a�`��B�#�	u�u[��C
�rb&��kݛ
�t޻˽��ӣ�m�Sp��"�{��E"�}�L��)�8���(q���sw��aӾ��3cY�����0�0�R8ը�'��`�O��) c�m�С0H@�m���Q�̚:��c�c���ݼ�����Y@Hᮄ��C� �د-�1�n�=�jbj��ws�]S����᫳�h�*yP�P��-��eU�F��u�ۗ��5k��pg,�9ݨ��J�����h�T;�l�l����
��@ル.IY���G�)7��[�(���Y����~T��&\t6�	�w����cw�1X��T�m*&�3Y�k��I4m���n��'�,�9��oU����c�/=�Ar�NÉi��|�MnfL	���!�1ڮ6BM^s��nR`ӛ}�Z_:	W	\���ױT�iQ��Y��I����L�c'Q���K�a�l�{@u Fц�S4u������	����⛿�4�Q����y2e-�T��@X�f=�<���d�n�n.��nfaN�ծ��2o%��b��!Rɲ�K�le�^*;w��;��ګ�H<\�T��%/���TzD���z-��bYu��f����V�Ot�#�Z���ǘq���:w.�OKW]E|)�,��w՚�tWz
��_Th�9N�\�Q|JM�3����� 7����}�N��r뢨A����^Z%m�}������3;���6�P�����y��ӦU�}���ll�u[6�lb���,��ۗT��c��������ģV�zi0���l���ӭ��/j��Ư�95��UŘߋS�'.�N�G�z���>��������p�.�y��X����*��g���z���1T��1.Q�%�H�	N�[�H����=����Q��^�7�ܐ <�����>��q�͜뚜܉)�sQ4��F���W���|,)���]t���1+���)����ۄ7�{���ֶ�$��n���;�RL�>�
��s{����G�������d�o*42�'}�ob�*+XG:ňּ�lH>����F��Fs�V�	tR�t�q
Q���q�t�G�'b}��;uTN�Jl� �����x��[/%��ܩ-�řS&�>1�f�}�R���CX�Nӆ�O)7O�n�"k�*�����DL���|�o�s��k�zn�< V(���(z��c�ͺ�^��-��)3]�R��Vb�ζ�[i�����R���J��h�.3afC�����+=@ﲚW��M���dfk�َZ�huS"�cN�8O���/�H�,C���ߌ*>=T�����+۪;2�b+I-�$�I�]��'�Xb�E��6d�T�e�?A�0�=s]\��]�{}?l=O{\�����*�˰ͧ�}��±xi��?x���;��P�S'kH��� ]�<�5���rW>4�A���9'0��8��E�#���K=��K�C}Y�ga<n=j���flE��@����a��5Ԥ0wB�$�UD��7����7�%�M-��S&�s ������[M�w� Bʘ�^�+O�01��ŋd��9��=e_Bqg�S2�E�������w�}�n��K�vdE���I�)���"��T=f��Lqغ��Sj��+Lckr9�c��x��ӎ}�xEk�"�D��������j�q|�ƂXR"("�����m�PKP���(�-�	U�#DBciv�p]�U�ڒI$II$  $�m�E��Ջ@  ���{B9#QR[�z�a��R�w�\��	�ޤ�]�\��f܇C��P���ɠ�%{��:h���'R&�QE�Lm���7�]It�6nZ��ˎvf��y��$� �-��Z�Z�Ѹߌ�S�*?��oG��ړm�7�����}ՙ��B�Ϗ�TB��­�O�?�d6X��!��i�B�E�q�ɰ&&���l�)�m�D;�������bc����Q3�(Ϩ�Ip�Y�
}���b�}��&�O[Is�U�cd�
`�9T�.�`��K��ʨ� /��.g���v��γϣ�	�����>��[��~�p����v�Y�U�G�f3pA�y9����x"Ҏ�e�_�L6���C�� 4���=��r�#b��^���]���6˟O���x�5��_{˼*n��s\Z�X�Ÿ~�EU+֘� +p��ծ���ӊ>��=M�m��nɝ�6��i�E�
�j�p�����OQ=�|dMj�.|�R-�ӷ�.3Ψ��hF"0��n�Ѹ�5�}�8hP�^�;��aX�n�CHe�71)��}�ɉ������|�_~���~�bV�B��,$@봨�߮�o�/7�K͖����"&�BTvr�p���ٕ�v�;��e���@��1���ǖ�`4��1Bϝ���TT�.���i��w,�$.�N7�"�}�d�ȟMS�\�x�!������m	ƣ_5�T(&lڑ�bR�F�[%0u>Pe���:',�]t^(s�#�f�+�����P3�Y�T�0ha��g�.語��}�*t�&Y��M�а��r&[��$#�������%5�A�^-w%���C#tr��Nj�	\��]��?��>����ǢD����w��=rԐ <����'���s�̲%�A�6K.Kh�X2L�F.�YN�i����l�׻�D��[ÍZ�����A*a�}���GHG��6�/jG����f^혞�X��ZF8�z�oj�Ў�\mA8z���x����|x_�f�N�wu�2AU^���0,k5�[^�sO�H�ߟ�(vh.&"dH�*�
H()�DV���a8l��,��S�f���zKך��s�� ܜ1hC�c��K�N�+���&Y��J�_���,|]����4�jZ���Z��[��㯮µKx��/P��1��zm��(��A���Uը�.�J��� �+X4S��[;ّx]�'�����|�>�� E�����S���c7����*x�n<�}��  ����9�<�2�	I��R����D�����+�5�U�3�~�����'�/B������k,r�zhdv��뻶L/^ke�]0�����������R��+�>���/�!��3n�8o���M��HV_�ZQp�Ѵ��4��;=�BQ��ĞH.Gt��-�^�:f�}wꄂO�ٞ��ۂ��.���2�9�N����h`bqB����F�9n�*	�`�ҡl�����v�o��@��\ݩ(uerEmv�n���оv[�����=�\u���{+�OK9��u�Ӣ�Ƙ7�n�kzw�v{�3>��E	�3y�٣�S%��ЫOzj�jT�=��u
?u�l�U�%���KH��m��~b�$J�'� �܉���{!��
�yh{v4�&C�F��9Z���N��\�&����ev=a�ث��S5#�{l��6�e�љ,"(| � �����0Y"�0b?z1М���a������4�2HW�V��ܛ�����=+��S��*�:�n~�yj�!�b�=�o�Z0ȵz[�院h*74\L���,t����Q=��-�U:�]�.�+	��=�G����>�y�*g4p����[�Zq�����'1�m��8�d
dRW�gyI�Ts�Q�bk�٨��갱K>�������}������y�����#m�  bm��   [h   �����wi�9-�S+���b�t���1���"ә�.�L8�/2�IN���J8�	�Y�5u_����I�S%�A'@����=��B�J�ˈ��tReInFےH�RA>�E�I��EA��t)�L���3�f��Uk_/`׏�5��ŏ6̯4��ʖ��bbp����I�`�+f 0 D���x���$d�1B��Zr�{)��5�]�˻/e['	Fk�삮��ɩ��&���}��}ꮾ}}AJ�ߪf{UGq��Q�c��5Kz����)���Kh��3�T�#n��ә��������{P�hC{r]��5vWq%��� :N�s���̲�^��"�S���n�� ��[ۓ[p�t
k�=��:���)��UUI%�h6,��E�n�&-�����]�D��6;�9��*D�)==g�^��g���7(fU�F�Ї� 6����~�av��^3�.|#�����a� T奵kMv���_5��skޭ�̕vz �d�x��n0{.��\G���tA*�:ٻb1�l�G�B�5%��V2w�𥻹T`��<��
B��1]2>�W���V�ל;F�����qE���՝!!�kfX�BJ�C=���J�-WUU]m3��~��^Ȇ�y=O���K�P�.���wt���P�SO����ʽD6[}m�ӌ6��Y��כ�}[;35��a�x;�F�{��y���������-�n�k�ʙ`�f���0��m�	2�<'�\ZT�(��#�r��I�5�G�'jv&��]�.&���عk$�Y�v�&x���]'r��:�'����Dň�L\�L��\�	��N4�U��{���%sݨ��n������o�SV~d?n�<��R(I�E���9�/eM
��^�0�T�YS+hU��闏���z�w�߭\�3" Wx���Uh�0�S����!o�������w��%����vpŦ��e�G�H���bi9c�O��/]k��î�J�+z��*�9v�7��Z�#��ҍ'=����<��ª��~���`��W�=ݚn��sq�!գ"�Nf���M�m����I�iqTN7`3,FeX.��aO-���pW�@�/^��=l.=�S��g����Xjv:n.�]�*�$7ю\�w{�b�u̪Z��)�%O��]_Np�t���8E�n]�6�Lĉ���Ȥ�a��t�l/L\tn��.������ �[%]�adt�ԹC���A����UtOV\&S+/��V8��w�lm-���X�`t����z=�s�z�R�� �1�����-�2V��r���(�01�h+9,��g�p�Y��H��)7�t&�I�=6�6��	
��\U�x�,9��l��:Ⱦ�J�\Vrf�QB����5���}����}�����=���䍷$*|�`��J��%@]D��˙	��ɨ#p�]Y4r-c���RP	����}=B�r[k������Z	��D��8/���T;�Ƀ1t�oz`��	o�����%�=$��.vkyJ3%+4(Fp��	����{~�q'=�G�l_ٟ��Ǭ{fQU�����K�J��"�K?u��LIݳ4L&g��ol�b��3:���^����JRE���Kbi�fg�.�#׎H�e��d5��E#�  �;��,���^Z���plK��RϪ��n�b�p�O ��c��l�p� ��K�g=��0]���ڥ�I<Xޒ#��Î-��uf7�+qS�S���Hp��h%P��i��9.<����'6��U%�"]9�9}Qm`F�r�*&���%�K��X�^)�.��;ٜ�{���l���,�U&G��F���`]&�jKqAŊ�T"'�;��A�ȃY5�ҍ�$�l-��JQ�=�:I�i$)���A!�*�5�7�qя0�[��2V,�����a���H�DU��� $��h�wE��;��v�p�Yt,c����<w�VW1����3.,��QAX��e���My8�H��3	Z��%��Y.���b�)`�j2L����I�E.w;���~���sJ�R4t�D�����H�«=ArL��bA3$m�|��|}�4BCIE�}q6F8�T�(��D�)4Vm�1M&$�&&h�r��c.��U��~]��]�y��^&�nSZ´'5f��˵u40!��t�+V�8��t�
��ok���Ɩ]�D�|H���Gk�|y�#��V	1�s�(ӭw*�H�����1]�/����"$�jٳC	�,s��Ǟ�<�N���ϼ�=���       e��m�-�      m�    ]܉*Kf�m���m� -�         ��[h  m�R��        ���          �y�>�����߹>=n�sp�g3p�	��i)M)T��k:���v�8�D�+ɍKW�[��۲wHلp���#p�,ԲV��߷hf���K�h�Y$L�����6�5�*F�VM�䒤Z4yGJu`w�8�d��kgū�t���FN��pW|M�1Q'筕R��+�� �6ﮆw�{�1��a��I��kſpcF�xM�IѼ�P����2��z;Nޘ�:��qqhM%��)��Wy#f��{�VŢ�;�^�=ɼ�ֺe���֦N3��L��,:����Vvgci�iһ��i�J�yxv����-5�����Y���I�tK�v�d�GtK.�S�y�nr@�Zi!�zŻ���6�un���B���t��3$��V�q8�
'1'}}��%��N�ҁ7&�v)��l:	�4ѳ�l�Xj����5a#h��.��J��x,Ȭi�~>���Ϳ)I��sÌ��i�7Wv.��eȍ�.
,���H�p��bg�-�ѵ���J�e֛��-v׹JS�h�!2*�E��6�)�d��DLJ�S�-�aBH�M���p�8M�J�Lgk.2h� /�O�ٓ�E�PPƏ��٦Y$�m{hU�6�ȩUFHj����3��: �^`�N������Uh�7�V;x�Y{(��y�Fn1g��l�B��#=�A��c�y�������@V��
��|�^L���7�| Y  6l   �Ҁ�� �>�{�j{}ϼ�}o�X�6�P�t��$b�R�u�pZC�ou��ڱ�tYH$؉�:�KSE��0QT*�(�l8T�<��j��e��qt�Z�P�(:H��	Sr����� e�I�J�{wl;��Q.&[	[M�b�"���㗢�P�:F��7�o ����<�K�^�F�\w�-"|.�]�Ƞ�)&Lm;3��:�t��b��_c��k��O�>�$DL� x��q��J�r��ǮIJP^z
���G��bC��_1:t����O��n����n�n�f�n��)ΐ�KW�6T>��\���i�:���R�?{n��P��y��1���V��9'P��S[g}�" 9;�9�6-��\��<����>�7�|�\�?[���nJ�L�7��&�()1�JJTb����<���'�yF��:�]*H�7�4�OЅKf�4���[dE@$�&SVz��>�հm�� ��YcД(�	(�-���QX��(Ȳ¤*�T������b�m$�VE"�im�=�U@��i��E"�0�^��7h.�B�n�& �U������^;>�eʹ�c3U*���:���@Ӳ��ѱ�%\rgfp��ۦͦ�j+-m��y��t�X���u�����������;_Y/��Ԥ�g�2��.�3qU���]�����oX�=����ꖹv�������{���x��[��^uWܹ`T�����BS�\�F�͎Z-��L�������W�Z�L�Ms=	 �)�����|���Y4n�iF�ih��Va��{Vs �za�M>_]����J=�A��1�l��r���W}��/Q��g=�\ F�V`��<��u�5*7�����	����p�PBݖv�l��[<�Xo��iΙ��s�v�þ��7��1 �H��r.�#w����z#T{����T���ۣ�c��ay���u.g���v���c�s����T��F�n.%k��Rw5�S��B���+��1#��o�����҉�����Q�Kw��Ѹ���H�w~\��4�)ͬ��)����e���8I�����Ż����UH�NRN��t��BCm�/�ț���),]"�΍�f�Ӂ7�K�2��td�R��p^3-9���jALm��Hʦu����kY}S�S�U����h��Y���r��h㤞�O1r�͊i�cے|��~;Y�X�/2�ʧNq�_=��O�f����.E�Tn��BW�w��+S@ܟf�򅳷�C��6�O�:w����UT� ��F ���x�{ď�o��n6F���[ڸ��tgt��7��}��d
�h�rR��7e�^�<Z;2�VN�2�Wv��=�rN�m�6��C�����ևN��}�蓻�y�;8[����O�g;��߭� &3����v�"ۄPC90e�L��*�n`����rmY+f�q�����˷3[\U^�|��|����=]�U��D��)�=J���Wuo��\�6oM��Ѓ3�<�'Fh��w_�r5�(pxS�Y�e�hi��;9�9��N=X���i�ɷ�>ߦ릶���R�[x�w�,�{(�e��';{��}�&�uf����Ŭ~�5W.T�P
�kv���Q�e¢��/�ɡ3"Yg����]J٧�)��� �=&Cx"�K�L�n�gv�v�Ɛ�2v���!`�A$�E��u���ޒI$m�  &��P   m   >���g�ʀ�U�<f�h��v��F��m>��S,���˻K��FSi	w3��c6��]h�D�������� �L�C��T����-Zՙsnrc�����x�������~���\!\�M��Y$�NC�R��w]= �}�kKG�P���L�RЖd�1.�;]ܘ���D��\Ͷ[+�ˀ�V�;c��G��<].��qo�N��|�v�n�e����vm��m�sM�`W,�`����h����X~�ءO�g]U1���>�ц=]��ȣV���m�]*�p�'.��M����]׳!�ܗũ�Wo7��9s��sj�=����֑V��~Y)`s�O*Sۘ5P�A�=}3���H��������0�)P� >r퍼�۷u�{n�IJi��f�%��P�NlFnn:���YR�j�Ml4(���O�\�-�\Η��t/SG�'FCr�a��� J+�n_2w1�u*�y���|����GM&�Y2�EWS�ɨ'y(�pbNYW{oX��^��q����X�>�/�r��ߕ����\�=��|��n�"�У<>�竎���6u���a�0 A�9]��0U���*�d�l��f�ʊ,����[5Jb��2�e̬����dpS�������ja�B@u&� 2�j�*fKaY�_*Q��`">��M��hVm��\:��xx^�.��{iH�Ե$�m$�dS2�MɴL���d2Kb�S3]��ck���)>�ێ Y]�Irf-�4����]{���&Qjwbzvm;��l��N���GJK���s_q`��\́;�ڦ�����	M��)ׂ9�]��R]K*ts���"mU��P&�.Tf�wc���׷��vye+����f#�s�Õ�k
���6��Hwv���*��k�S��Z2����K�T�}ٵ���J�7un����1kt�ҵ��7\����W(�Ê�_��#�g�oOB�@�� iʈ��ȷ<�O<X�r"#)f�������к�)T4�ٱm7�����d��	�{9��s&���K����y�zD��d�����j];���޸6���A�[~����5Cϋ��($1GJ�GA�� Z�d�d����V��b�͗�����R4sN�V/xzD����T�����t٭K%�'�1%����Nn���Da0.���t=�-�^c��Q\m�j/��F2��6�5�t�ǅ캨�s]�	�Q�
�F�Y2��r��f�[&0U"�*'����am"���b��V�����/Ǥr��ͬ�&���d4�z�snsy��JÊ]Gu��lϓQ���LA�SW�.59^V�ΊP�OT���̾���~5@�;�@`4�G9�Z���w-I��!7Sϛ����,�J�go\X=-�M$�d�}PEU���4�(ȘrG*
�f�P�:.�,����5�r�e�%gW��7o�o��i>�vp�BR3K�=/Ϙ��'%O�[�eY��"  3��Ὥ����"�P��C5Rkb�����m���ڰܪ/h�ȫ`���U����iK/:���q�M:g�mU���s�^!�#�}Kr��	eͅE�����PE
D@c��g7�٫��Ӈ�Vg9{�-�iØ��Qk�u�{5ו)>��-Z�qՎ�g��t,O��i2�u�}s�W�I����{�;>���@  ��   m�I-� ��9;���r�����{q	�.q{�5�)oQ&�6���+���G�eX�͜x���|�BD��3#�X�F݈�I�N@��)�ԗ��($����ж� ����ɖwnI�fw�T3-�Z����VK��^Yht�Vx^O[�h��Gs�c�Y�+�a�T�6���x[z���1�8+t�]'v����� �����%�XFN��}�V(u�3{�^���<N����B	���Y���>�}�p.�K���۸0��!4y�Վ������=UVp�*}�� @�ן.���3׳�g<d��j<r�1q��Cw�Ӟ@��Jh8�1(�9��qU�*�i�J�2{�M��G��ϫ$��$m�)B
�<bV�����P)��n�5�:8����%����}���<�Sb@�����.k�w"^�.3o����	���x�Z&'�I�^ْ��HX@��@Yz%���88p��!�to#�s��R��7�9��8<Fԩ�g%�b��$$q9�_f�WX�u�G�ʻU=�}-M���s�R���㚞A�˞��o��������;/g���j��8VP�7��h��������2m2���G�@�H�+����Wd4n%����)�U��+��ϫ��p�pUӲ�v�����P�e�D���M�dQɍ�Hu�5�`H.�(o�g|����M=��H����7�a��B�kh����R@�,p����7�|�3�P�k�ݫ۪nq��d�nK!��f��J���P� ��#�El�������@&Q��_C�{av���9$:��I����[�*�/W*�Y���܍�_(�'{uh��K;=ύ>���69��L�T{@��6���훇��t��j��b��Yۑ	�����70�&�c �*!i���G}�ڡW�^G����#;R�EQy��f�)��7�8C!@sǖ4��6��9ۻF�1�#lD6��{������Nv�܃	>$��t Yf�q�+O^�,���=FOK��e�Ud����ȕD�и�#��VB��!��n;���=ok4�BP����f����^=�|�{;���h�b��:eX
��ڋ#ZiMS���+W7n��`y������N�X�e
~�Jh�	S-�h��Ly�3J%l�˷P���Z���z�mjpXwm�:4ݤ���>�R�%B�L���T�����cm���P�*�H߫��dj�@- �V:�b�d�S0%u���xk|��T�e@�J�MT��I�bɌ�6Z�9��eѼҊ��X��wsѳDU&����HѰHb4�D�a��	�"�>%Qm)O��@|	XrY
�=�h�PX��b��]�y[q`��U�IT��I�<Z�Xo�:�*b9>���,`��[)����z��%i�b+�ΛK�Q9���2V�2%�7�2��{(	NA-�d�޵eB��;[�iWL�C:�[
�x����ӝ�:�79�UnQ�"q�|J����ܹˬU��<G*���5�iާ�L��l�٤q�oT{����ϓ�nJ"���A������t䦕"j-��m#(��T'�Uَ+2uI_m���:�;�n�Y�Q��G�*��]w�3�al	�Xy�5ɖT�_a9u۝�p��F�%�}�$	;��b8ZU0���z�P<oL1q�s0��-��a���S�L�
�!r�Bf"\e�ԏA��`n���O���+G�i��s�uod |5��"�^9.�1K����{a�x��H�F_CGn�G�.Z�i�gfSh��1A<ZOLP9�/l�ʝ�󂓥!6Y
�R�u6��!�����%S�u�OTK�o���p�4͹�{��DK�Ks&�+3��4N��[%�`�������!Usw+�iҴ9%�xm��[�lV�[�i�6�1��s�f�[�b3{/�1�C�8��Y����)��w_j�Oβ.�qa��1��4�l�r:�I��H���l��/���wOl�H����~Gd0�3�_�u���Čhb	t�N�����.�^��~�>���*���6�R�C�ޅ;zl:7����p9=rs�f.��[mfbsw���|�@cm��H�(�R:DN!d��A9�Bڙ+����csN�y�9��Y���"`�B�s)����'*��w�-�M���=�`ë��ك�������E5�i*�nߑ��vN���Z��%J����u��>������vY=�BHL��y�l�׎�;��4)dvY<���aŬ�nv�sN6
;���y���UIT�v=��*r��>�����P 9�=v+٣��������i=�0-DvI�tR�t�$Ɗ��Q�פ�=�����cr�H��y3�67��{���P�78��u�}=>ќϴ�N�� @oW��ᕱ0�i*���I$����Q�4��B5a�B��������gP|��p\�
]O6(a�i��)]�^�E�u�:nR���Ծ�x��ӈ�MA���{\/o�����j�R�y{��v>A�c�Q��L.$�$o��UF��6:�r���kί��"�bi�b����׵{SS4n�����N4���F����}�L��&�G]X3t��{��T��0�̩k{�-�2rw�0�8��=���w�ѵ��H�*��B��WGB{I�٬����܉�˞�4�f�AA��TR�*����l!VA��.�f��כ��;���<���m  4��@ $�u m  ����|�>��ʵ��G9�� )@��R�=.�3na�ٹZ��y��$��f���2sF$�E�A�I���H׷4�|���W�T��46�p�a2��3���g:7@}���_s�F�8Ԏ&�r'2�U6bx6��dݮ9���c�/��w��(qǻ)�҅@�ސ�5f�|����o��t�92r��>��-)ޱ��֤����l��b �{��]ʔ眮��Z&�4��R��u!v���-����Yݏ3٤[�B��1�|�$T���l�F�e8�1�LXtwTc�Oz�^��z���=���U��w�Kb�9�5F�|7�`M�S��^�r�~�" �]��OE�}��q6�[Ƃ�ӏs�e�h�䍨ڝ��T���ʄ#B7
�ҴM�Σ{����|9��51�V����6z����q�;����\�eyޥ)M�u�+lm���՚�'œ� ��O�I A���l�(���f��N���3�W�e�n��z�Y�C�`�V%�vݏ�K�Hw[W|��+����n�� (k�|��_i�Թ�Km�[���Y�a2e2�l��D:������m�#��Ķ*n��9ږ��[����ބkwF[���:�EEs����\��ϺVe
~)��� V��\&s�GхmȪ����{h2#�&�W3~�����V%X�Cb!�æ������:��dVB��c����m���`�6��NX2J<S!�ܜj���֙�~gW���2�;ٖ�f�E`��.�W
�V,<{�wlc�m�|���<cU���t�w�N΅���Ϝ�ü��r�Qv3Dn�%H�Xy?`���j����b�Y�����y�}����٣}��i*,d"��H�a��z��r[�d��t厫�2��W���7�k�w��ȏ-,֢����u��|���[����;v��r�e��$�)��n��n©�Y��v\^apC~�t�\d+��j\zι����� �,Ea ����H̣v/��oY�#)|x��7ׅ��2�Tˁҍ���^�nMc2$$�]*�h���l��s�i�E�w[[E2�@ �1��w��qq!�����0����N��bX�Vw6�o3qt빦n�/���xk D�U�ٚ��� ����9b���v��,���������8�Ϟ�5���ֹ�z�xÉ-�����tu5~�{,���{�0�|O�p�u����]��{c�*��(��
���R�7��{�x7X^�G�U�.�q�ذ�<�b����Z��A 
�oilˊ��M��>�o�3�0����n��]�-�+w*���Rc�;d$�䗵"�%��,<�)5�T�6p-ل�G\4��Ԋ�{ʝ!���Ƃ���]'Чp\<�}���\pyi)I&�H2��<M�M��dX�kH���F��#!�=�-�s`H����:�UZk/2z߷���C���E�d�&:��IL-�>��"����t���o��A�+YAs�+Ϟ+ZN�������x��ֹvv���w!v6��'=dv"4�m]nA�]�ڟ A**���������K��]Os��YR�'�`�}Þ{�W.b���v�R���v�y�t˛��=�WaA`�-�0��ifh��ٖ�&6�js�b�}L����6���<�a0xYQE`��0dF#���{��[�o�� m  �[h �@-�   ���ϳ�s��}��y��^�[��V��Yt�j��e�)N�S�Gju�N��:�!@�Ue��I=9��m��*q�@�R ��4���#&49EP�g��&�pX'ګ)���/�L��|��d�7Z�ۋ 5��h��9����[���Ý�u]XR�����'=qYT �^�=��]r>m��<+[W�t�.,
:g0D��u,D� C��["g�1����8aZWfMcs�\r[x���s*�P�ZA �}��'%�T_�e�;#tVmE�^��+�������g�{;�*���,6�ٛ9�*��_��3a���>7a�渗�r��5�rн�m�z��<;��́Y#z��QS�1���������W���[���I$�-�˦,��1<�QA����Ue7xSN;`�$�/��[�R9w.md,��[��A��x����6� ����d������0�p@I���ʊ��䭝\�7�ƫ�I�nw`��k��}+��_�*�>�K��4:���Io���B^�I��O|r���x�]ýs4��G(��+mi��I$tV�;�"q��=�;eq��36�E};�9���Bo�뾘�q:{�m�d}�!���'��ۨ{�lu���Z��,H����\D���-/qƷ2�u�A�ѷ�0$��!q)�r<%c���9?]�u:���m�^�=�n���1�xL�^f��rZ�RtKr�#(�=0�1Z:N��s����������g����a7� =��l���H<A�{M�ʕ��T�I�s^w������� �#X"R*!H�x滝�F�w��y�B����~=SKZyY��'�7����=�/���X�@X�$x�>h�rv]ޙN�lut�������׳/�3�,fRa��ϰ�4�k�ͻt�,S5,흔�>u!Vh�Ϋ��y��IX�c�fn��8姥��G�p)�y9>:�	���7Ov&�ˡϕW9RT����aˈR���nL���)�Wt���ԽR&�S��d�oR��;�{}��� k %%�* �͖�p�N���:��:�>>��C���^���N�S�;�p�˕�Ɨ,�v���@�Bk{�;�[�}������5<��췊i�f�V+��o4I7�U�q�1���r���X{����_v����b���pT���� NH/�c�,Ƽ�^kw'�.�U�ɹ��hq*���Y/�~�<�3u+�7UWuwT�EP��$UY��H � ��u���Z��KQ��{��zj���r��R��(-��Xe44�K\=/b��u1mz�y>���*w�l�7MNu�S
�P>�+�ݳ��)���z��v(�'i½T��7�x��I$�O]]c�9X(���d�O��-CL=:q��be^�s�Y�	X���3��Jhry�H�9V&v}�Ԧ�LV�(s*���OY��3+�2.�H���H��p�3�5��Zz�ͨD�'���/D{p�����;��E���\�N��7�	��ui�i�M��J��<�bl\UV�c=�R�x�T\h��]� ן)}0" Me��T�I�����2�xl�S\�8ؚ`�*�L�r���Eh�$�v.u��ެN���L����݊b.�ў�VAˤ���T�uM�Ji�c�%у�]��q�Z���%��"�`�Q%i�Ҹ�U�(2�u3ݸ"����Y�&ѫ��;��]s�k,0U#nu�%�O��W�Z���+q�&�	b����d?[�yX��h��q�R�`�a��)��e
�l!�ZN]�J��YPf�R��g��*���F����`�����R��`� P$Y ��p�e�
$�	V�5Z&��*H]�"��*�����`�I�7B�7M�&q'���Sb�f�NM:55[$���*3+jh�3�f��d��B�wt�����,v\0�5 a�hC��!I��	��F��Ӕ���0��dS�g�1��H�|I$���3t,�ڑ�\�.\�Pd=8�[$�Df�qEGN��N$5!��pf�@:ɤ�`Bn�<L6�&�b�䐲,&�IW��j�# ��6�i�A��9����LV�.4�iH1Cl*`(CE�,�4�?@�p�75K���ť�?C:Y ��v��"�!P��n��u<4JV���������t*�Q;�������������G_(�Lj"�j��f�E����I     [hv6�              ��̻�mIeE[Vմ [h ��         �-�Km   ��ٳm     �m���   ��       �l���� ��!��ݰ�ɽ��D���N��&U�zn�sے�v��_�r{������V�Zk Iؐ�b�������x�����E4��p� �Tw	3����H�wa��.��P�,���nj�S���@v8�T���um���d�]8qf^f�8�b�gs�pQ�a��=�ڳ���a^��������1֕$�ǔzr�;\�q�͢�/�@�ܹ	�a5Ɔ>*�ܮW\-íPEd���Ggu�a�@�D{|ǭPȯ�̔�g��b�B����w^vo�e���M��yN.��~��O��o��wY��>")��I}r��ADM� �����ș����oA��9�G׉fQ�.��`(��L�x&������]�U���7�����*8��]��dx-��^��s�C
ˣ�*��ԺY6���B�i4�u��9T�a��gqr��۹�E�r�[l�-�Z��!��}w)�Y <�j��4��F�[���Q�'mh�k�JY¨����������v���GI�m�� �.+��d2�� �*�"uToM�(�0��,�-��eJQTqEI�e܈F��"�(P&�ؘ���P>lО!H��jU+��˫�6�'�Ϸ��9���+��� ��\�ێէp��ꪬ�7�(��
m2h�4�UIDr��g��?7�k�pa�f>xUt�(��U�]d��X�!ڵAy�����)R̫���*�5��@m  -�  m�h ��I$�k*wmM͹��5�+pU���E���ci0](n�5����kw+���Bvv��G��E�4�%2[	�F���M��E4�Q��9I��y�wvkf�
��X�d� �6w|���~���n��d�ڋ ��nǕv�5�B�kv�k׼��$�j���湟wZ���!R"� �?��/4�u���cX���;����e׷���Bd��&������Z}��a`��6$}0��'W�v2�7(�y��z�_2������FC'y����Z�Z{sv D;�1�rߐp�ܳ�RO�<� Ka�<Y�37]�	��hg�=o��[q���+���}P�ӹEI�b���k��9�rP�+k7yU^��-��m���z�݈Q 6�@�r�`$�N����3gT�2*|{z�"w�OOy�T�+�FP�a>�u��l;+V�1�=� �/k>���߹�\�`�b'(ز���bEAT�l��)��Z�X�d�a	D�(, "��(S"�r{{nmN��
��br����EA1M6�</!��ڣ�f鍎��	�nr�8r�'�K���+��N��yIT�Ǒ�Z-hE0�o.��9z`7����1<�)Sܚ��
�\tS�Z:�DB���L����g�a"����ީxen������np�ƣ���ҧ`ѐ�d�ț3܃	�ƌ24>���R�)OMv�26+/�mm{�;`�I�62�_<.b �ڒUUISnI#+�m`�1�4n���JdR&��][.��*��*��!q��:���='\�����QO��(W)�"C�Ӥ��������&ɣ��"gZ�v����Җ^dDFAnєh:y۾��ʚ6�c8��Ku9�3V*6o����i�[>�٤@$��p��bլRZ�Ś��
�Y���oV��a0��q�����nDڳ��=�����Փ�sQ�ئ�R���~�P�ܓy��	��b6�)��ٛ\�v�;���r/��MY�W=Zz����2G�����	�e��}'n^Î��v7wz���z����ߓ;�}z @��������/l�yrw�o���1y���(�7)Kqd�V���Z��إS�w����Oi��N�[ݴz
��P[��<y���\���r8l.�:۸�9�E�˺��n`�� :؎`_���S��n��Τ���`��f���:�)Qg�OW��[gB�=�7��5�m����O�
p����	���|��]-�OT諍� �0�DdQM{��9���W\O��sA��(i�S-�����wR7���r�Bm�}k4��۾���Ĺ,gw��N�z.[���h�6iPeQTP���Ѽ���K���F�I�C�{��V��"�߭5� =�v=�H �^e�����[����U9��Z��:����d+F�yd%2]�'��s�]uh�.�|}gV��n�� �=��W��j�BfL�M�LxfS2��]#��D@�WN��9���T��z�qL7�|�u�j����+���ގZ\�[
�=�*z��>yz�0���{�j�;h�k�9�#�s:�0gb݉��%�P-�1�c&i�se'apj���wN��΅ � �NyUD�C7��ךj�lҗp�]>������#E*� �
Q��F�� -�  �l-� $���������y�F�����*%t�1�9Z|:ؾ�垺��K��8S�C��Sof�V����o�x�Yk.`I�$�"�aF|L(4�0�����2kFO7n@Ʉ�K�N���Tn�Q�o���2��濙vٵ�7.�홇)BǪToWק�6�����+���z�h@x�)�ז*2$vJ�EҎ��;�X>�e�.����)^:e]�0"�RĐ ]���{�o�[�
d.���.�-IW�],��s�]��SIld�>y�|�8s��mVjE���/�� �sN�y[�9����5e50�W���7�s���Y�i>�B��*��"g��l��U�o:y��Qy��D�͕c�s.�l�*	��%>��y����m��]MU�."\C�%0�n܎�ͻ1"�N�DMv���P'��}�/Ԁy�q�S2����O��+	5dx^�y�8_����ޏ��}�g��G�1RE��"AdU����0F�;�S���H��}4�{t���z9����֕����碱�pp����ɘ�۩f�x�D���m�j��v��Czs�i��7�|���]Ak6������}x�[�ڠ��%
���>u���*�ڹ��z���t���Zi�i-�Tu��0����aH��{��<Uڅ���� ��=*}��X7��)��ucխ*(]9g{<r�3�{x~&=N/\���n�W�7r��� ���z��'.v�܆%�^K�Ht���օ��ыbҪ�P!,�'�O݋�����I����e�*]����&���q#��g��2l^�q6CL��Q�K�Α��#Gi�ʦ�����ɒԩq��6��s���2c_x�w�a8��  ����t3r�$Z���޶!�n��l�z_N��*��v�<\�����|G��v2�D���� ��S��!VZ<��fLI��w���wLY�D`�NR���Gk�o��Sʔ�I��˿qy���T��'5<`ɣ�%}��Gu_r�s�㱽��xq��&vn]����	v!KR䕒[m��p�OW L&h�F�c�"��ƣh}���Ǔ<��v{&G�3J3�*k� ��G��xy��\���:��Mk5��� ���l� fs9d���V r��u�������c�wR�S.M�i�(I�<��uÒx��w�o�>��U�<NF�pr�;���"C��ܬ��]������;����7������ٕys��<�S]x��b�Bތq:d@��ZYXH"�`�PUA"2����ˠ븁�tWIE�<�j��_S9j�8�N�V��mw��`9Bg]���Y�I���Pa�[)]�nCnP�]���*}����`�TJ�sKɰU[�δ||r�Awz��6y��v���o������6��3kk.rBܐB�m<qW�b������ˉ�}��By������C<�&�z��i9����Yh>���f���qc�4ĥ�?q�g�+{���f���(<�Rw��7�6	�y/+~CyY�Y�T"��X�],8�.��fq���,�gr�S"��ҭ]IHh��{���*O��/0n�q���r��G�ܐ�ڽ�(޾W���ҭ�}"�;(Gccf�@��v�H�W�Y�w�y^�j�5�%�Ӽ��e�=	������Z���(�QDX�H(XE��`��(�!�	�[UVTI^�׽������-�  \�h  �� [rI$���Ͳ�yuu�����^�Co�SMpntKtgUE�	�*�9[f[h*)��.Y����L}����נ���RSD��	2�;�uk̳T)�wnr3��ns����{�z$��F��Vl�n�u$q6�-�ڒ�J��@���b�u���m�L&Pq~�}T.�-n��ݝ0��H�o�G3=�g��\o7m�qP��Gfӕ�������w���bCه�FG���9�[N�h�K
�5��q���F��^�Y_y�zf�u<m��a�~+*oΈXC��'�� ��͌xOpa�\�������ڥ:��7����(E��e��N�i6��f���f_=uP]e��j{#3S��m��$���z���ݶܒ6ܑWˮK
�����VK�KW�[	����Vk�M�J7�����&�����eWk�M�70:��.���҆����}�%��w�S���݆�	;�ߙ�i�ǥ��5��ˁ��.u@6��op#2�t�]@1a֬��M�0�ú����V.�J�*������G٫�>g�n�C�����Ϋ�-A�N���YX̞�d��${Ӵ���y��Ǫ��dv1�N�{�W$�y�B\jm16�glnn>;]bh�Z9��鵙��� �J��ySf1�q::N,�KC�Q��}��:Kc�����6.�ʬ�&v/Z�s��J�FC�����Mv��-&�M�B������Q0@a\�X�SU0Ddh�+��O��ݣ�-+מP+�����E������_L�l��q}SMtGot�
�oQu}w�<����D@�o�Gbw >S���au�RM�5;�WXb���SW�E0� �K���u!(�_Gφ�䎍�u32+���K����ޤ�j}��-��г��-���3��oO,ޖK�
�̓8j�������DAr�ؽ�#�^#MÑ���f��j-���
�L5k|�<E��QD�.���V�A��S5���e�n��"���,f�;^6�B�I��c�˛F�P[��T��x}���I om�@e���ۭa��D��.�F'��[6ˆ`b�7,*,Q�AH��[.��܂-.���C�'DGNd�R��Y[����	PW4o4�,�c0tȱ�2�4Y8�1�GWC�ʙu��4wx�
��"@"�f��7w����҃���e��R�b�}�K�6�x�%!�"���{N�� '����"c6�8��KY.R���	"��"@�X�3eRƏ�g�$��d,ж��Q�ޡ=V�Ҁ��X�;��݋�QA�X`bf�0GVƖqkmU����á9����
���_4u۽O4�׾ʋ{L�b���Le�K�c�a����P�|���ˑb�H��̈́t�Br�D�+��Ő��E.�u��H-�q�{kT�QL{�@Ռи�e�im��l1=��Z��q�۷��K	�g���^'AK���mwf$ np��8F�g�F�l$���7u-��tg�Y'X�ܶ2^��z�xofF�9ģ#��jY���j�3�<>� `�wG���6�+�vW7/7v& 34�T43W����V���Y�ԗ�>���E�2��Kb<wP�ڭ���u]���:WMeɔDî�̜��n��&�����NH�q5�� ��7V�ⱑU5�(R���Q�*,�ƾ�To�Q�o�؞�;N��1wh��իp X�T�����q�,��d*�x�r�3-d��{9Q�g[Ts);�g�悄��!o�<^�/׆9�0$u�KC�;D�K�1�Wl��#�:���_K�e@�ズYn��Ja-�DxY�D����5�3ٻ���v���x0T�fHf��9�sx^JWr]ep���Yʲ(���|�g����qmvﰕ�;t{�8�]�㥞 r���Vnu
��S��w˸�@�z�}T�=�6iMgU�&5r{*d���ʹ�fxˀ>�z�/D�v�`�J�#�\��C��1���//{ؙ:lrƇ�Xם��y}(�y�b�d��̮��]P�@oWa�;�P�2
��%��m�-�e"��}B1*��R���	sUS~�G:�P���Y���?a&l�&����z�1ms�����*뭃���xx3�}T�֝�cj�L��D���)vꃴ�w�޺QۮcU-ZZ� u�ݲ=QQ�q��}@@�� U��;#ҵu�!�[����OХ��>S�3��4a�1W���mv�TFEN�^b՝oɭ�\���߆A���F-uҞh��e��w���O/�im'ĳ��m��Mu�wF��7�����}g5ۃMV�Ty�����S�t�R�U��0����c,��F���x��o�ɟU�� ,�K;��$��^|�gJQT����B�@}�y��s7�ݶ��7�o�L�ʌE�q�C#�y����F�C�+W�٫C���6���>�W|u��F^���
ńC����O���?Q޿��Oe�S2縿���m����z�9x�y�H7��P���:c<F�b��� �Eg��ǌ_mv��)�f[�;w�/(�V�q�KHй=>gG�E5#H�0c2�R:>�`ޕHgv��5���Աi�b��,��s(�|NM��,�����7��;�.�G���~�a�A���< ���0m#��gbk�º�x{�
���WOb4�D�B/��,H�� گq�E��镕�4�y(���y�]���(Ą!q��RT0�g�/��D,�5����H��`V�Q�{�O�@$�|LY�M��vI$�[|�  ��  �m��@ {���s�&Λ�\�Z��䖞�Uʒ�<"�[��j��V.�:�5-�JF�ґ�Z518�̱�E$A�Q�F�ט�����!�&(��*�������6�n[�<��iKm4Y���e�j�Tt`�HB��	R2|���,���- �C��d}-���חI�oڿ<P�|���g���|}c�v����Dza�帜6I*�g����س �t��6@�q���rH+y�X=�C���4��H��}���؇��R7��kF����g-�J���EN�:�X�~�CO\$a��ă�#�d�#�.{\��ڇ׸�0\�t~-(���J;5���D��+2AF������h��;q @�����^�Ͽc�B�݌��SN�ܧ�(���L�GR�8�M!�Ղ�gLV���m��^U��|Ek~'e�0����$j}`%���ٳ@�x���k�஭1����8PKA�A2!��*^g�s��^���/"�j$Y�De3;�HҎ6ܐ|]���(�U�i�]�H�{N�E��^�ؽ�4Q�dןf��#�2U`� ,� A " ���}b�w�3ͣ���OG����8柫H���!4TF�;�	4e6a��W�Fn"!�]�����c���k�v1Wu��Urqc��K<�1S��ǥ�]���wʈ��K�48���/]���<�ݮz랜�;�v_S�R��&}g�����8B�+��ן@(�-��`)�b�#��w�rH�����a|:��� P�FY���G�
^��= ,��tɘR�oFGX�<��dN���k�j�O>��HjՍ���Y�Qn��h����Ă���>!�gR��>�HC�Y��i{��)څ�R	�����a�nD���.c�--t�M�S�p��d�n�6|Gi|4��i�de�swSf_=q��x�b�	OH�8<x����z^��� �;���gd�zҙ�s�H�z��B���GVϼ=��I�F�l�����~�dU�yC�Vg��G��a�i')y�a�iO�۟8�s�z\ ���;Iif�#�q����U���8�N/Y�C������F�����.ΆfEx��@���װ*@���*]�*�d�����@`���I?m��*��+7�wϽ�iy�@ȉ�'����v�3*`U�J�C+�ٜ��z��|���ҩ���ݸ�K%���vɣ9ly��w����/�F�Kh�/P>sC�� g�d]����]\#��P�Z)�;gt�K����^F�8��#�v�2,��a�!����ޒ:m�Kى��.עN�?i��/���t�U�NC�1�q�p�a���s��4�ዙ |t�G�^��^��]{��Ro��fq�N{}.n����$��$�I!U�X1N�`���
��U��x� 3�#U?�I�D���Haϐ��#��y4���XJz�ݮ+�nK�r�U@����$+�j���l�Ht��I��1���G�vFة�iǢ�>>%�Ŧƚ�4�us��@��W�_�����,W��lѩ��[vv@ӐJ����>`|cn9 {���#��{E����>yd�ޤohH� E�Q���2"nQ�A�gE,�n��t>#��0��/q��h�3�~�Vd
K㚁�,>�[���(W��]T]��h�n�]9�ɐ��X���Zr��zپ'qLI�rE@���s�[���M�׷iR�b�>'���j�d�O&�tHƔ�6BI��� ���#�^��Ėa�[Ű,�ζ����[�Bqfd½n�A4r�\���m_S�o���c�S��9oY���WͲKm��m��"{��i'�n-H\�ϼK�s�`�@��}ɑ	��|�KS奚4p�J!Z�=TU�E�:��2e؈B��	Q�VF�5�0�Hf/���2��U�+�Ah3����xW*>�H4>�a��L�rP�ūX�-��}��(���U���  �4��j<�$���	,Ƚ��[G�0�/�9�)
���������+�0����}�h���>�_t��3"�|h~�eikh�� d��f��]O�A���0�Ȣ(Ж�դ@a��߾��O�qɝ�0#���ڼ�>*�L{��B>Wᜌ܃��7��0VQ�J�튰��~;;����σ���A���C �>�O�٤���k�H�/�et�s�+d+QD@��V{��돼��������m  tm�m�!h�@ 3����c�}������s�y2W���mZȥ��M���f��5q"�P>ҝ ��a �	@��1Aʠє
~��G 2�)E�*&�NHnn�s.i��Ӌ@bٜm��0eJ-�$��I�U*��h?!|~ф���f��-��D"�H*P�'�J$�|l���U}���J�|��v|���dD�Hi=�*!-�����f0x��5.z@N�B}՛���0*��؝b^���:�t�a��?�fe�V�@]l���t�J�C����4]6Dϋm"�Q��	O��s��J^3.BCZ�u���SM��3��W����9�̠�6sUn��dgy蚡u����tڒ4�����0d*#�L�1v���ydۛ�_<�;��|Ͱ�<Nu�����G�
U�(�vI��;�=�b_b��1c�ՙ{|��UI���h�b��m���/>�Lv����|�|��N����۶=@I�?Y�N�a� n dP��USйy4ό��>���a��'������܉Å��'�;oy}��Ī�Z,�H��6�`k^k���|z+�H$��C#�>��Yj׾���Nu�7��H���%j

JʨE�HF�2z�=[5��k���Ů��S�|�����.�[���M��p����h��x^u�P�W��Bլ'~��@F���0��T�G��Z*f0���)ԣ��\��񈑇���V[R�+��IFw�v�E�`jBv���8��1�o�0�4p���D!T~�ۧ��0� 4��\s�!�5T|+���-�mX=��Eh=G'����Y3Nv��ߟ_^���/�ھ�@m������wbs	�vGFD�(H�E��P�%H�N��\U�DH�+%؈�	H�U��I�d��8)E#�:p�ؾ'W�퀙Xa�ę��.��G]/��Z���m����29�G(����*DS�jJ�w���z־�v3�\9x�^�����Ƨ��i:�)}��$s�TMU�É�����5��q��k��oϳǛ����3�E:}f|k�����-G���*�X���+&Ξ(����dSϺ��}CD�ogi��#��_JrE}��{�{�uC�	�ǹQ
�n���������|�Y�{�1"�b 1 F�,��q֪���ǳG��OsYu�H�٢������8*�7f�$��昫�9<���6���eUJDc�� ���i#90�#�[ ���u��-�V��+)+uQ;Fb�;.�+�&�㔆�o�A�b`d�&���v��I����z^1���BK�@:�`�ut�|푱q��������+��ZG�s�*�9�hQ��g�Vċ�'�Ř��}���e{�|���N϶H��F�m0S��52�6ʢa���17*�#{g�B�&,!�1A*L1��S�C�a�0�.T�8�(� G���/]~�h�dO͌9X���+�rϗþ��D}#��#�"�4�	�f���������>O��|�쫻�qS>�Y��uE/�R'�iCW�ڂ��d{��8Yr�h��t8(�XNnt��dX���4[B������7Z!ƽ�!�@�Vu/xe;T㛡둜������ӥY����=f����5�|���
�ס��U�݋-n*>�v�t��>���|m�<�3:��
��(5�QH�Kc$a"�#�,� ň1AUR�µ�����RD�b��(�,{���3�s3c��>��5��|�[�&��N��Ӽw���2^#3�uft�Y;�����V��s�z0(f��c�A�Ԫ�)*]|F�*E��S�Lu��B���ѹ�\�^�H��c�����g�Hft\>��e�9���4ͤ�gsl�m�3��NZ��s9��78ͩ
9"��	��F|��>���cB�^������<��Q��5��>���ꭐFskk�Ts����� W�l� HΩ�edi��i�-)���FnL�/�X�rQ�!>B���:(`B#d�~�qP���r����%C�*��D�ĉ W �OЉk�ش�-��؁:G�X�����H��<^Uo�,���n�,�|�8�(�"R��#�:\
��^q^�2�ܤqO6��P�f�
U��Sx�{L͒�L�zt����r%s�Em,����(�$3�lh<z�$Ϻ�̵Rv8�����8�V��]KO�B��e���~�y���4��ԇ�i4߷W���o��iqo�i� $���I	$����$!��HH@��K`�a	���!I	$6$	 Bb@��?�$�$�>aBل��&��~}$�BI'�� I&�� ""#��:�?��h������~�������?���!$� HHI!?���'������HI$�g��?�@ I$��>�������$�o�� I$�I$��O��0 $�N�cY I$��9���~k��F� �I?�@ �I?d��� I'��$�}����?��74?�� I$�o�������� I'�-@ �I9��?�1AY&SY�O�3��߀`P��  � 7'�`a�;�   �      TJ � �P$Ƙ            J�
R�!J�R�����%% E$��R��"��H$IUx               ��T�*�  fQק��}�n���on�۞W�}�Q�������޽�z��v�O�[>�vrt��`��u�,(ӣN�8zwn+^Z�x ����!H8 >�����Ǳ����}���=��=�m��l��O[�\����n�6���>��/��n�s�O�z �/�v�;ss�"�@��:����   o�޶�;��0����/�w���n��t��۟��{/g�}�:}������ּ\�����:���_/��j�<��(mT�C������_w���^ӟ�+�3�s�|��{��G֊{o����sw�u=��ﳼ��w<��=>���gA��(%�}��   ����.��o]�����
�^�t2���}��x����vw��v�ۡG���A��ymQӧ�J*^$���݁����=���[��1E��z�����g�����g��OO�<�T}��=̥�p�����P{�$��6�����  ���O�ݻû���랏&��d.�s��C������K����۶v۷��X|��ӻS{};|qA���}���f����� �ov٠EI�����މW6P+��y�Q��q���_s��;�ܘP�w�^t}��vSݮN��x��ux�Gop���@*xR���  	���C����}�i�/�q��7|۞��^�+�ץ<��p��H>�{}�ν����V�x��U��|��Uۣ���ZJ�5@5V��ֺ&�Zѽ���p�����n��O}����u��/�|�	}=u��t)���/��Kױ���ܦ����'�RU@�@ "��b��P` �L"����{E4 h 
���UR	IP4` �~�*�   &�D�4I�=@ ��������������f��I��H۷ص﯒��^�\����$� Jy��I ��$��	$ R@���	 @��� ��H ��� ?�_��|�_�Md��[����y���ތ�)�φ�d�L��0.�nv�/�E[�
������XɨL��4�~��:O��ђZQ�b�Ƙ�W�.\�@f1Q�i����z�2L�zח��@p�� B,Qj��q �o<�i";�ܙu��DeOwswa��Rͳg&���\����p�Pҵ˽�]��se�p���}Ǩ�ui�ΜwA4��U��owwp�E��vU̳+썀���KOP9[��H�g^�w�H�0�oλ� a�N�����Dq����ÖP���l��TL.�`ͼ^ӳ����ݰ���)m}ۏ���jr/9dѯ�s�v�I親��(ZBz���d�d�c`"4�E�[�7V��y�Y%ӯA��6�^R��'{�#�Y7�%����ou�7�p��&��=������HK����o[V��Ν��ڲ��ZԚrm�u=�;�k��ځ$��zd+��ڡ���3N�y�]�lɧvk����в�\�����}R��q�Y$E(Jb��C�G�Փק���P�����(,X��%I!D""���� *Ȥ$XH�B�ZQQ*A�*[le�*2�ej(6��"
*��T*�UD`TR�iR
)T��,���R��
�ER�jQ���E"��d �Ab��XXJ�YEUTb�1`�ֵ+R�����D��������A�(�b1b���d�QH�)#�e�`)UF
AR*�J��E�l��J�k���R�,m*#*AEX"

"�1H�
�@) �*I!Y$�E"�*��R
AH) � R
AH) �*B�*B����
�R
AH)�`�Ad
ֲ�� �jAHT�d ��Z�QH�+D��PP
�R!D �*AH)!X(Vb�
���P*AH) �ER�QdY*T�¡R
AH4�T��R
AB��V ���R(��Z
�aP�h��m ���%���
VJ���F��
#
��
��
B���+R%`ՑK�+@����+V5Th
B�d�%eH-m�j�YkB�A[H)�!R ���R
A`[H) ���R
B�*AH) ���R
AH) ���R�
�aR
A`[J�R
A
AH) ���R
A
AH) ���R
A
AH) ���R
B�AH) �J� ��Ȉ���ؖشTVAR�m@� ���R�TQ�TT�TQ*�-�U�e
�ZAa
� ��
,UUX��
�*0UTEQEҲ"�R�e�F�"�P@U�#$X1�YQ��T�� ������`�PP��FR
�EI`E�"�
��|���HY�h�	Sv�DB9<���pYn�d%.�*����S��\��|�n���NƤ��s�Y�c�,��XE���"J��,XBZ��2�L/{T՜P(�f^kZ"��2�a؀{��qn�7��Q�3p̿�8�b/�vZ%������"�u�Fn��93n-�	ج�]B�옎rƃo,h/�%����Y�|������
}�9�B�͓��Fj�ؘ9S^d��8�n��4d�d��,k�.���=�����Y�[�蛙��ޝ��2༳�����^�ܻ�Y�9�����gLX0��\�����×)˙�f�{�z(#�B�9�����C��k�Kq�����2�ϛOm��W�o��Z�/ho5� (9J�$`���;մ��š��,p�����pn6��Y@*�{��sy���0j��M�2��Ͱ�D�kwK�*�ḥ�<��0d���ݏ/M-×ru
/��{�`�س0"pfMd,�d��5�Bq�\�A�YLm�r8���gz,�b�ݣ�  ��J����vr�N5�sgo1Ӭ;�]���Ҏ9�y��&3\�/T�h�Fa��s|�y��-�m�}�(z��/%�`w�G�x�A̘3E��h"�,;��ww<��74��eIF�T���Fy��vs��~������DS��L[5S{�u�:UcX^&��f߬y�+��̎w,�82$��U������8N^Af;��*� RoXR+ƨo��L|�y�b`������֚処�@!���i$���J�p1�[�g^��W8�ӏ�JW�X�cʺLS�,Kpc���`g���&�����Dp�ܺI�>9^]�*�ظ�yvh��Y\����r�~㌍�="�9`�3a=����a�r|
��.0�z�Xx7�C0gEܾ����[��&d���!��[by]1^[�ܹݳ��z`q�5��n��;��&,z�}<�v��:w!�<�kg���:e��My�w��w��y�7��A��;�^Q]�^|`���ob��610}�B�#,F/�A��Z4lh�����k���HX�Y3�kvJ�3���r�������߀����:|�fl������	�����kCǹ�Y��v�F��^Ę�;{@��904�W��|��s����\�1Ϸ%�yXhTJ�Ta��� v�7y���t�s�C��/(�%�fj�"�4�h�q|�?��rDDT��,득&�����u��x'	师��T�E:��,��<Gv�Ԩ�I.t�R]˄@�3��޻ڒ��eTZ��Ӝ�Y��gh{��JعXZH�rlݻ&L\1-�-���B��#��y��֎��H�к�I@E��=Zn�s�Q�&\x8����	����9���S�np_h�����{���J�i��aK�#v��Cє�����C���gm#bB�\�pi�I8�\�z3�E�$+K���D����6���XKR`htx����/:b�Wi�^a��G����T�Ia� �C�ܹr��6#e���%����ZИ���Meb������D�ۿ-)?sJ��½�.�P�������o
�hۀ۷�3��é�5���`Z�������4a�@�D:^C�U�߫� ��HV\�a�	Om�+��M@����m��,J��]_�m�����Lf��j���W�s��위��I֊N����^<�][<����z��Y��ց�m$�J�4_ϓ_],壖�#��o@4oV/kp={���bͧ{��Pz�D˹r�A��ztd�	ӽ�Zx����4�����qQE]�J�����f;�ξf���/���9���\�c4_9��^^��,,|6U:=EZ�_%��j�m�!��O{ٮݚ��u�u�k���D�� ���e"}�|�w�e��w{�.�\I>K�&���C��@[F>La��;J��R��Y�X���K�u뇆ҟn�bG�9G�!�s:B��]�Q���+���z����\W��#_��w�	�*�9���5�4�;W]5���"\�T��Z����,�w+nЍak�\`S9�Ǔ�� B�_o���z�:�&(�8�0`��q�u�!L�<��	�H�Sw��.lA�Ao�#"]e�$���q�HnCНU���Q�E/��Q\M39�oa���w\@x:�zd'�:�>�q��W9V���^�B`�ǝL�g-�ݸ�آwM�� Rx�)!�&Q�k�*��P����wx�sz�Ŧ��t���!�gd��g:��ݪHr^ZV�b��2��z��^�o:=&�l�㊌��/��1��d�8�9#|�F�W�l����H\[��ՉqZ�az��ޯO�4ְ��������9��9��#8��E,%��񠳳�cP�"�Vg x��Q���2t̳��'N�y�uwL�YL�s ��n�x��ю���V���w �;q<8�1`�DB;%��d谲�v���:��J5�SZ�@�B#br3)���m�Βc ����9�fR�S;�@o1tv���q����2�!`9c�tF�o�_c��p}E��]���q)�y.&oC�߸D�a~�-��d|�It�Js����&�-v�w�tѰ�g`�X���錪�kr�؀����;w3d�vb�|̗+��y�d3@݄ڔ0��S�l:�����+Xo1��ey;ucZ�g�k�T�<��ER" *ɴ4n���԰s�	�oQ��cl�eU�y:��[����}� �|�<:�#p��Sd�(�k#4����鏸w��oK���d3����DR�H�����!Iٳ����lK�I8�p``v$.�1'^��wclGքە慪�M��ӶB��=-9�����N`N�	�wD���4�Z�U�&2F�o��[�u�r�@5�`����Z�h\�a�G_J��(H�vU�.���l牄-�XXeӝ���՗l�8�\Q�T���A�ߠ�f_��!l. բn�p����k�ƽ�R�#_/�dcX�"��J��lʦ���\���8���xICN�2g,
� Ո<9����� C6��
��tJ;6�w��s	��y3���E�{ooi�Vp��{n�7\cqC��Xhа��M�����F��۩��qi:4n�D�-�<QLdl��g{��;�im��p��jM;4�ӻ��b���՝�0`}��L_F�}x�7�F�����;c����y(qД��B��vvb�8;1S���i�7�[N�t�1��VT"�Ӄ���;7%'��~* u��<'H���GMf��ρ׻{n�=��n��tj��6��+wǷװk����}&�>��l�z%�#�;W`�nʓ7�w�gd�e�R5R%�\�e��A}y]��*���P,Ӗ�]��gk����BsF2�����xw��XW�7ϻ/�����q��|�����0� q2�Lܓ��.eȚŜN"�h�_�v��f,`������羈�xd�s�(�CD�
�#�i���`�f���!�m:��d������kq�-n|�|;�6e���Y�V)��#�М�q�̽����R	6����F�iDმ�寅G�&�k;0��m�Hkx�>��+|?" �+�&��g?�jO�V^AY�)���3�J�7x�v�hj�$��t��['�n�h�ʘ�z�� ��!5��*b/���m�$<��Tk�4�g1�p��	��3�f�-��!���U��Gd{�H�4�p8f����L����z��s�=�ғ[�m����mX+�xk�^#�g\x7&)5��#Խ;�޷q��O��uo�ׂ�uћ�b�UdLb�q�TT.W�
�w���<�0�% �^�j<]�������cƆZ����'��oo���	��܌�41V���F���f�;�\w��9�ɹ�FQ���q�����4��vB�X����e�2�gf\JĲ�����hܷ���H|�yNh��d�$#��x�'HdY����_�Q��^U�����2����x�ɜ��@q�7czf��B�ߧu;8F��`��է����Y��H����6��w���!#�Iԕ/�vԢ�ve���m�w�s�d��Od�fnj���,�8�+dĘ�[��U3����u�l�!�C�=��-�7M�0�9:�n�شZ݋�Eq�gK�oiV��_m�R9�_����zFaV��c��7�7��P;W�e!]��
�ȲKF�Δ�����bm#]��m�f���GM���%��[�lgJ�
y�\���JkkwaE�!g=Y��Y�m�����l�)�O��gg��`H��Z7Ě����MM���*Dq��R�u�,=w���e�}Kt�������95h���{ժs�g�?yh�QWZ!)�BDr��B[ͭ��Ⱦp���`��O�C��0��γ_{$ӱm�x*4e��
�א�� ��M�;i��D��5b-#e`��"��&��{}�}�G2��t�ڦgy�J:�OM@�3�W7�"pG�2q߆���@�9�`���^�����ר�E0#��iq�\�����W�нT�h4`��	=O��;���Z{���%��x>��;�sO�<���1�sbk���v���]��]s�_w.��7	V1�����
ty����uU�6�I�.z��J�OY=m֖�M�ΠoUW�H7nn���C�.���*φ�p�ŗ�b�$8H���b��U��j٩4oS�b_L�5�ngac�7ӄ�QwE�����w՛���$����rN杋eڜ�;]#wax��e�	�&��܌$F>@ٖ�'y������
�J��Kku��|u��V�JgH�6]�;)�&���޻�?炝���%��X;�rk�c��ݶ���Ӥ����%�;��ݺ�H���@�3��Kuy��ܻ�lP]�mxƢ;�){޻]�"�ؒ��n[��Ik��wF5;H�J/vϟ��.�;��Ii�I��k��s�$+��~�+�����y��umK�w�J�5�n��M��x�6�M�Cv2��6��&�{1|krfH�zGO�[=�[T_w��X�1I��yEMo^���x�v
�i����z�q�_M���Y�s�u�=��T���xC���!�u1���zX��]ݻ:I�t��s������$�$�t�����OY6ٶپ�wI'yK��c�,LBcy���&wb��-vZ��٘o���,g�>�<]}�־��t��_G؋���|W7����^�^.A���[잝@ܦ��(��'�N�纳A�+噧m��2
�s�5�_~�sk�}�o�)�hvq���m�^��w6�-��1�+��a��^Q��l�����ĻǨ��Xռ�L]r<����5��۲o��ð��}ӈ�㨟G.�/�c&qut����&��vfl��E���M{�ޚ�)-���P)�'E��7���
���]���z�'3����Dҭ�x��7R�U��P����]�V�orfs�jB�a��rt%k�ldz�r��H)���b[�wq�*�b��B쉲�����-���
jHϵ]Z�>�Ö(ƫ2_8�e�3�2�������Lw�%��v���ċ�W/x��@ɒ�}D�fy��F�wm�k�e��S��ڈ�V�^�,�zR�;�.��'\����R7��o�F�EK(�<��]� ��t��ᙃ7v�>���#/\v`Y�򮘚Cr4G�k�L��55U��������'�S�;���ȅ*�$��L�拜X�4�Fi�����& 2���uE��-z�	��Av�gS���Яy�4L��U+�_ ��u;���y�+�<��&wH�x��x>#��)k8#�ͨ�_Lu�LR�Al�����mb̮9�l2��G�}�q�+F�/,n�䯹}(����_#��Pv�ţ(�[1�(s.�� �M��A��X�	��������z�'{�=OQAiK#�̽�_c@_K���]�)!q`��zM����o��Q�9�_�ѡ�\/�26��w8I��tF�-�Wb����e'�.�Ru،�`���{z�()���YS�R5*�v�Q�g�]_@V���gwa%��w�Y2S}B;T����]5�ζ�\�v�\B��S$�Auot��
�t8��ǥ�*tW�ѭ��yr�m����m�{��t���f����)	W���Y봹�mrv�G>�\6�j�s��Y�lQf����O5K�(>�+=P��
�;F痫�B3vt��Dy�d�[Lp����ds+��49�Ȅ�A�-�{6繗گw�r���>�&<Zm=�:oOs'z�ST�<���|`I<q+g<�rfcj�Kǵg�T�n!��
|t����y:�=C��/]2�#�;�|Oq/]�.��sﻭ�*̨��'(F�]�f�Q��s�w��Јox�e���<��a��{��cV��H���y��Y6�У�����8K���m�7@���E�V�� 4]���m�ǻ�2��j�R4��*Rt�Wk�*��WW�]p��+m�P�Gz�Q�ۍ�Kb�	�V�g"���L��
+,��o�a�&i�;n��o�&�����o7��u�Ӟ�����M7
�����Vzi<�r��zRp��4�Ԭ(uW��%o:T������l�4�%��7��wׂ�s�goIg[ak��C	R��W�u�˽�x�T��~����wЉ?@��ߕhf&��̆� q��ZjIBB�] �C�SN;�Z�=���1���5 �F��xcc�q�5ծ?{��2����X��<�����{��F���}I�k�)�y���{���b���6�w$g݁�/v��zP�s�m�o�hacE\<�MUtI��<tHw9���=��xs3�*��[�V�x�UqV1�_���av�|,�]��f�z����2�Z��x	���1ٓn�ܳ�I���1��2N��i�Ǉ�$���q�F�(}",�p"I�Yǂ�jv�%��D�˔�-�o;tcB���`���/�Lx��׽�O��G�.��jJ�ӾWhw�K����q�żΎ9�1kk�ۍ���ju}��Bh�+�O�j�V�o1���r�-�}��O����s� �D�嘳ո{���&�OOoa��4��(�^��ƺ�BSU�xH�%��ʆ|�.�@]fN�*�B�v���X`�z-�
���36���1��s��>}82�g��e���#�h���N��,9x�d��=�X>C�\����uziɠ�7̜���rڷx��m�IV��񵗀���Ċ�r:O7�b��3�����s�B��K.��"�$�컠�f�&�:��xOK�	���y_��ys�&^�����}�­�s�\.�lK�D����X��!�-�i���Y�d�7w��!t�3�!f�{��l5��rn�w.�մ�됎%�{�-�sz1+�\�v+�`c���4+�k�qw���0*-����@�s��k���G�n@�8nZ��vk�1��a�l/.A��w��׭�=qݸ`OD�.���"w���Bx�?ls�1�8�`&{���v�1��sd��$L�j�\
�4��i�u�@S����u��d�� ]�K��q���2H�h����kt(WV�B�N�vړ��yh|��薶&{��l�KiQ�݋��p�w�g�N�gVk������O(�=8��'}���06�L��r&�{�9�L���^ܚ6\�=��p^d�-r���z=*��ک�X��P���2E���Z�j{��s�ܧٖ�P��`�vh�1\h�s��x�a�S�Xp��~E�n[ON[V����t����D&ś(B�.Cq����pY5��c��
;�-̐9�Vg=cq�=N]�v�l\�J+�׳�5���ڟn�/%��V0��~w�h��Mb���2�b�T����C�m&�ѣ��Xu�,ZŮ�v�{��_ggV~�ǇӘ�'&�ؽ1�Ҙ���cR~��}�K��t:��.��O$R����{u��9��q�g��֭+;wzup�M�{k�Ħ�Ȩ��jꏷ(M���GS����{c�6؛L3w���n�[j�5�{/�_I�K�������K������!��*E���LY�u�KM�m+f�'Pn�!F�ʧ=�4w]?��H�M�&�K�Ӷ��S�	U�헷�8~�T��E��r��5h�86Z��Lݮ���mI%5�^�Rq�v51�Mik�S�vu�դ��h�C�u2��e����z� Ggq�,W�BS���ʏ��J��hm�zp˛���"��kp)���:J�g>S��͞��<Uc�i�\��oqu��d�Y�UF�������Fyz���c�d��شMy���uԲ�ϔ�ؠ�V�^j�8�38燸��(��jw�F�#�4ށ�h��i0d=�+�7Q��m�C��٥<�W�|�u��G/��x@9��d�.^!w	Eͥ�7[�4.�j�(d+s�u��]�������G��05�2�ۜ�����������KWp�v������
6��^6��p)� ��8UOU��` < < U
�8@U⨁\���Q��` =T���N ��m��dT��=�K�p0��^��1�N  N ��c��[z�]��n)T�_]q���@�����N��7*�nuJ��[���*��-��[�Ɍ�pl�^��W��7�X��u`�����1�݅G�������Vŗ��	�÷��w=�vLꃄU� �VΝ��O=���D�ݪ-�ʺ��^�����{U�cw�@�3����	��8@x x80  N ��  x8QT e�6�ب.j����sX����  �UUT�p0  N ����	��8O*����Z�<��sǷ�g���b� U    x x8  ���ۋ��m  ��_>v]�{�� ��]�  '�S����M��]�Ud��βͭ����U��͐  U��l� �Tؠ[  |��T    {sl軞m��5Ԫ�hU���' cy�
���eS����\�S������t��2�+w��.�2���R�Kx�؞�rۗkҷ<�k�aWD�@ N
� 9�UJlN��b�Ǯ� <U��ꕦ
�Az�W�++�[j� zslw   �   �9�}v����uV��µ�튦ٳ� ��=���UemUc�ݴ UAT6ʠ�� ��U��u��2��U_��w^{k�ֲ9�T�n��wo.�eom� �V��m� �v��q��n� �����*�����_  V�����6�Nxwϟ={;u�O;u�[�wi�^�wZ�wG��m��mm����y���붽��N⷗���[Wy�{f۷]Y����O.k��O(����s�ڪ  �6������,��j�^�ݵݑ��e�T� �_  *�`��6�n��z�mm@���Y  �^�v� �WԀ  EP6(  *�:ܷ�ˊ붽�ud�K�����wm�w{�u��Z  ��       � �                       +)T �
�       �    ��� ��@�@��  m�p   x 
��    @        ��T z�
�       U p�*��*T U �   �     �@      n ��@
��  �    a�s�P �� *��m�M�p�UJ��"�M������!۰ �_>  @�h �
�d T           P                             � m�  Y}�                                               U    d���       ������IO{�۸�m��W+W��ֵ��BH ���� 6�H@�@��$� ��X=9�/���K��b�﷯��EOH�7�OV���}g����)Xu��c���\�f�ۊt?o]0�d=�C���>8��r�v�r.�۽����S�����|��Q�)�3ٴ�Oɩ�]�l��q{�ާÉ�}����7�Q�V�U�2	;p+H�_�ث���v�9_�j��yYRN�N�W�n,�R�oh� �}�޾��2�s2�#K�Y�n�jn�ܺ�v�edNB�QoӶ�G^s{�'*�;���n�' C������
�.��Y<��o6�y H0��&��N<v�b���j�� 5���X�����ٲgr|4=S��m򾡼�d`��ut����2�8��:f��_�R���;�ˑD��U>��|_���'�oF����.f:M��E�7�5�w;�HK�E��ھbe��^��^H٘ę]�r���'K�gH�;L���۽�k�����o}���W����Al�O ' c���ا�lU�u��@xT�b����r�oeܽn�S�Px8  ;� ��y�Ơ ��'� ���m�<,b���ՕN AN�ۛ=+ V��ׄ��7=l }o7w��7 ���c*�����*��{����rW�q��Z�y�zU�RlM�:�p�²������w_UU       U  � ��c� 6Ք   �  *� Q8V���)M�UY@         *�P         ��q�g���׾���������p�z��\$[��d�^SF�=�<=�y,x�W5t3�s��E>y;G��w�I$�m����L�ݷnޔ ���6ٶ�U8��\�^lO;�l�������]��  �W� UwUm� U �m�ϳ^��{�J	b)IRD�JDI1IU@�Lb�WSjb͔/M�x^���Nk�S���2��؜�xf�D��Ͱ|,xg�}_}V~�z��]<�I`w��I{�{i��;�l�~�[�u�ݒy��)��$�e��phNZ
�S�>�����������m߯5��p� F��CDE����D���Z�Azc�l�u �2h��ӥ��֒���v!�]>ӹJ�8����6��������͚��M��K:@>��)��U����GF���Q}�kԏ��r�DߩC�~}�Ù����(�f0=�6X(��]�;1-]=s��-������5���_ݻ���
�v��u�k��ف-�_�� �L�*~���t�t�
Y�wt;LÏG�����R��������F�Ɨ�� �q*F	�{��w�r睷d؝O���^�G������4տ9Է�
{��2�=��q6,��qgt�\���qۡc�C�c��n'��+��=$�n����c�� �PK��E�PtF����4�f���y�!Μ��e�;������
��T �?$?.X�%�(�3~(���/5,�A��g���YI�UM��b��a�f��L=rVE��/�3lM�#(�=����)��d,w�7�����V�{� �nB|��A��s�ٮ�����Eݜ��c���?@C�z�(�@�z�EGd<�׶�!;%L��T��[�r�EWO<�¿  �Foj�-���4�)�����{ރySŋt^��E��nD�١+� 1���	BpxA�4I��}��p�4=#^I�6��.��­����뜸����ʈ�Ad� �b,E��

��D�AaPH�,A��(��T�Y�*�/ݛ���-f��|>���s~nȢ4�Ut�b�ba�k=v� z��=�(�{�]���� 
α�ԭu�V�a�N�]G9v���%t&�A�{ki� 5r�ܣq��b���y͉��om�,m��q:�^a�ā�˼��]}�s4�7��+����JG`ȳ�5���,W�:|�Mk�aθP�p���w;��Zf��jr� �A�Y|s�^�����_}B�m�fB��	6ض���h󊸚5Ɨm��t���gI��۽N�����}2\ع�͢�B3���wg}sr�W����w[��t<MS�z���˖���!3w2�e_��+���o*�!�8���Y.+#��7/��W\B"YQT��H4�i���eD�v��~����w{g���t	�	���X8Ge���"�K]v��h �nY�j"!�v8yw��>�)�ǽ%���N�ؖ�=�}_!T}��'����,�Ҡ�G���)M̳����^|޹�۹��5�9v)��}�g�u��S����s=N��Ēwp�d+$)l��E �l�*R�c���,2$Ĭ�٭}��w�g�y:�C��OM>���gړ�n\��d��78�QA&�w�-٬L�X�8��<v��<�Z�4�K�Ӽ�z?�/7������0셏��D:nL�R�pW( �doO�
5��z}|��=����w?pZ#׷v�׳@;��{ �W◼�G��$0i�R�� YPcN ����\d�|P�)Kb<�g/2�!�~���?>�_r��r�|��k��e����Q�o�v��bgt�'3O$�O���
������eԁ7�,�q��xn��R���D&�7Ioh�C��oM�{�ͼ0*������>�&5�Fz.|K)0�6N��i���-�Rs#�Iz���Yh����>V*�,B�H�*�**"�U#,��ݳ_Ww��o��ך��R���Zݰm��`�Y�<�:fv�ä��ޘ�ݴ>�0�:�D�����jm�M����T��Ol�R �TD�}hhO�U^W����7
N�u}=��[��'�,��kQ8�����`-N��Q8�d��˻o0�����Y<���'yQ�[H�v�v��J�����Px��������
� -�  �*�   xw��Ͽ����U�X,�ӷn;���N�P;�-)G8�,V>ˊ0�-Ѳ�����f����ܴÍ�g�ꪯ��f��d�3ޙ�$U�b�>˦ɠN�t��ja�~�5�_E�=�ŏuڡ9\U��^g5ފTJ�Ktiވ�Y�E�׻�����q�/��ib�K���7��r�ei�k���}��si&�/a��j6.��3�~�iv	 U�bWhU2I��=������G��n���6OB��<
�h���0:�=^�~��� 4�;�o�MG(RS:�"�mV��)����~���<������N0X-u����Q�4c�%�6�-�bi��a��[�Ƭ�\�����0��6�O �X	�h�i%�8�#����\��Ik��=�w�p�9���tBN0$Ry���ߣ������i��I�,Rf� `h |jn]�V�y�l��~�mZg-'8W�W�}�ϳ�󦊹�SҐ1[���|�N㠺b�e�E�NQ2��M�����.��]輔A�~��ƓXf�8��xP�f0�(�)���L�u_F&K�xo�{!���46q�?$pn8�ٹt4b!n�c%�}U��/d����3~�כ��u ��QA�� ��_k�{��I�]�������t�+�ɴT��¸1W��/^��V�H��`:�W�n+I�[s4���F�g�gҽP�@�ÿ���КLo��+Ib5��#ܜ|x8*q�4R��r��X�f.�;}���+�
���l�o��4��	4�ĒI p�m��I$�m��2~Ͽ`Ͼ`� X�F#�Ȋ"��������K~u�ִ��'�3gs�肭�Q�t�;��������F2L[f�
B��h���F���5x�$��z#��	MZ@����۹�t�8{���M���6�]�:g}�������z�9��HM�	!�䀊��Q@b�VE��Ub��M��r�Q�4�Պĉ�e�`
",P��N>yu��χ�/s^�{���\�����w��gEH��3cX��>�:sKz�:���_F�E�A�p��� ��7M��tr���n��W=�j�����w2v԰Ǿ�ﾩ5LZ��o|P�����M���jA-��7�Z��aZ�sa���.�����~����i{i�~�c���'.�`ʺ˻�x��i$�I7�fD lw;gow"^GkՏU>�;l>^kW��f��} [��w�$��o��v�n9{�޶���vwaۑ M[�O��9�Y�yV��o����>��|�]\��$_}� D�.��o݇'\{�f�����X"���g�*2����[b��m�%��w�I}�����]��`2@bF$dE�`�PT|0F��ǩ����Dj�\���=׃����m�Y��5��ЗtznS�4��h�ɻ|V$[�^��{�n��eػ���y]zEUU_,z�>��j�_W�M������S�po�fܳ�;���/o�K	��I��8m�����͢j�@9�Lr��ɓxP���t�ǝ�~����������t:��B��Q>A񻙲lF�#����7����n�`��@(��TPW�!���V@rW/l�r���9mM]V%!�M`�Iڱ�yQ�u=Joj�2ij�t?DDy��@�4��Fv����B�����h�7��۾�ڔ[M�/��[�����/2Sy諭�������L@|LS��um1�|3v��{�gy�}��_$���$H(UT���pҔī�.���wN��}n�p����]��v�j37�ǶN��++m��	��,�/j������ew`T���׶�b��詵t��f�7v��wJ� m� 
��  *� w���������k�<�:��Uw*�S������Ŭ��nqJcl,�ޏDa�9����vWU:�\���
��*�]ET�9f�]��5���Ip��9w�/ވ�a2�
)ॻ�J�|�y�bHop��n��Y����{޼���������'�L�~������\v�=����]���#0�L_7��r��+JWQ�)c�A�v7���~k�r��}�{�HI"��_��q�S3D�˰uΝO�b��L�6Go�M��oӳ� �U�}Ս8�>����r^��.����
��S���3T�V8�DD�o,��lL���v��j�R���e�mƓ��ӛi5\Y�f\6��HI߈|l�U�*2(�@b�$E`$X
�P�++PX1�H*�b���QTH1�Q�i��5睹8u2�G���W���V�6�K�-�%g���⡁��_H6���N76�SY�3z�/��h�Z�\�'���S��_�29�o�}�UzWw�7+T�����B���:��l'�5֚�!}��|�9$waj�{�W=�_	��,�A�� �@C��
��˜��yn��_{$�+��0���7����B��s7�qٵ���]��krrĹi���֯UU}E�k}^ͩ�}������XN,)�V 1~E��@6�K ��"�#�=�M�Z����i��e4'�_mG�d�,���Oh��W�z#+����eY+&��l̙,���T�E�7*�X�/#�?X��9(Ρ�=����ZSy�� 6�<����1�&���(��W������_b|���&>v��]]sE]�#-�U[��-1Cn��YY�t��������!6�EUSԯ������QV*���hŀ�E�%V��5��71�XM�%)k�,ny~�6�l�Y<�kU�L�a�̓�S�wKR�ݥ�{�o{k�7��5�it��]f���f�պՠ�:��b}f'�ֶc���1�U2c�m��u�s1j��<Gw�o����k�4)��4���<��޴���}���1����uj�:���Qj�R��{7�kUB�.l�G-4���߼��;�9MC� ��f�P}}��� A�m9�&�Lɳm�I=�>�_kL��9��0�(D���߆?|3�y�#�f��R�7����e���x�8�8?���>Ry����G�o����y�������&��H��f��<�TUDn���5�-����Ye�ڸl��N�ԫ�|�2�n+1Z�a�=�BS�Q�agt�
zrk

�ԬQ������Xk �YTMZb�uj���[�����j6�֩�X�f1XJr�-D䙼�V+��g*bZW���ۆ��!;i��2��]2^�x,��NP������܀\R����<�'^�� �>���+����-t2 ¯/:�Ti�]w����kN�^�"��rs�3��l�e�����傝���]�FT�Uld����Gw�I̘��X���N����߉}-�cgf�Tw��U��䭫I�"e*�i��G��:�]�m$�
�z�z5��i�ދ�_vC���H��ʏ=�w������|L��X��r�%�~�A�Y��æ�|�2������{)���b�z��e��6.w��M��Lv�{Њ-���c�8��t��_T�=����������k~@$n�>T<&���A�r3&�l
����E]��Dܝm[V�����C'>�F���:K��H�f�G�vB��۴�7�xt�1��#Fv�S�<�mL�Y'o'��Œu)f�e<�+�&�F�i��wvй+R���b�^��_zgK�������M0�'2�r��!ԓ�)���!�1%d��? z���
��I��8�u���ֲ� x�_l8�|�3������~���Hk�ʟ�Iu�A6��Ld�Bu�&�u(OXi&��4�!Ԟ��X~C��|�)P���Ͼ�~��~��|�C;a�u�Ri�'~��?|�;�:ְv}I6��q�N$�a�q+f}������i�����A|��;��~����e�>N��Bu��\d7�p�xÌa;���<`z�d���� =k'�m$�8��'�}���w�y��m��æǶ���@;�����kX��x�P�'��������3y ��&r�a>a|�z�V��I�'���OS�Fx��Đ�)���B}��k�����!S��P��u�q,�Y�RC���$�{���Y�p4�	��4�������u����5�gw*�j�1�]8S���S�їf��y��}.��Ku �%�j>j>��N)*MD�U��~��(�D�y�;�r;�_}��ٟ�\�����ʏ{ވ�y5/(|�k�ʹ�k�Y�w����d�NX5F�hV��Z��j�m#�	�EAd�V���j���Ws����ɂ��v�����(4^�FḤV�L���{��*�y'�O��^�����ooi�D�̽k�����}�}G�ר�URL��V�v�}P��Nk=�g���9{�o �DI(	 ��z#��:*a�'S�|�Eĸ��o��.{�[񫿗�G~���D���'.�h�
���uֵw��DC/��]O35��
�W�KR����(����lw�.o;=��}߾���R~��)
��(�J�Eb��KFѲ�[d��Q���ך�u��^�y�Ӭ!c)\�V�㶜��%��g�ۧ�Y��ႜX���N�Y�6�f9�:���z#hc��Ծ��l�}�kcu&�
i5)k�bbݻ<)I�����H�P����E�(���}���;� 쐄oﮤ��!UP-�����(4�� ��ۻ�s=5h���D4�y�+��W��}�f���>��V̲m�_[������~��|��.{��k� ʧ��9�UP�p��{�=��٭ܪWU�V��u��7nw  �;�P�m�   ��n�~����>�{�D���ޡU��W����w'w���.�ѣ�s��Ct趥��#�*  ���w��Q�0q~3ˤV�Ҕ��UP��K����{`zP�1?�en��aH���D�K٢X�Q9-���p����ORu���5����k�Zr�Ϋ<�|֞��<���((*������F(,PA"( �@V&���b*��)!D+` �ϸu��xCD�(=���j3rt�tl̡��L�ZoK�]Y�%�Y�`����RW,p^`m���}�է���Oƾ2��'ea����kx�:���eڝ�k�ࠁUBOx�̎�
���
>6 ��N�&�u�٦i��A{�3�D{�?W��C�ԕ�=�1wS:p���/��������*��ˈU��Ix����h�:�(c���ޟ �����eN��{�n�j��L4{�o�y��Dk�<iGz��J""*����p:*T����g.�Ӷ���5�׹&����Xxi�Cɷ�!I��ަ9*wn!���O�NnG�:|�c��d�5
��^潆�ϫ������;���b}'�"�H�# �s����治<��k�ټ��u�Ф �h{]�C8�/Jl�������9�x׵J�/-GA����գ�
"&��4x����S3ͣ���7^�1mKޣ�@Ių�L��eO�E�>�}mcJ�R0 �0�K�1Z'jx���&�=r��q=�DG�6������<�5oUҺ G0c�DQ`-��9{�S�����a%����i��������n��XUxU?���|�/��P�
�#��`s��D{ޘ�u��__~�/�[%�?xj��d�X.�F"����H*��u�lk��=�夻��Kt�Δ%�1�D�tJ���=�Ȏ!�ȇQ��s��p���ԛ��I�n��EI�x�Ӄ6�C�u%�8Y8�z&x@�Eb�L*�ru$�&�<d����U?g��w��ʛ�'s�u�:�Q����r.�/ ���z��w}興��9���x���U��N%i����^�~���/~�om?~C;k��M�z��I��6ﻇuUUU���7�}�Z/b�v�XS�����Ƞ��H������ܞ`�;ŉ�e@���p�KI�ȣ���7����=��)��ނ��U_�15d� 8u���)�>��y�}_ I�~S!�d�w����N�M��f�ng�Yvƫ�y32�k��� N��G@{���G����#�X-��sێ���0�7�z�u��_�5�5v�{�������i���RÜ�|X�2�|;	��"kU�����_.���x:$�
{[R�dq�	�%�v�m��3�A}��Ëd��z�'�ByM�7�߮}�~Q���k}��~D#*() ����?����di
�(�V�c&e���Ν�|ߞs�:H����i���Y<�*���9�%��j��p���ޞX�^��8�c�	Wk��%� � ��IL�.�Ĩ�:Sٖ�RY�tX�s�"�xU�RҊ�#���G�� <2'xLT��wҁ����#����w�⪱;�=o�;��.ۇ�-��밐l�<x`~f�׊����(2+�Wޓ��bS:>�z<�=�r��o�UJ��Ƞ��Gy>��z�V�Vr�QȂZɡ�לS�Vu��m�R��3����{o���#f2:��@Ȑ���ރ�l�u�~o)���˅��?��Ei�-)���7%72��Qf��l\�S@�@�����Dhw�v�;w7x"���=�=�!����o�PT��\�5��y.��#a�/TS_Z�r�$��pq�v��#�����²C����n������ޏx "��bAW-1#Mi�t�[9�\�{������1�D��Ag�`�bFA��������Q��"#EAT�mb�1EX�T�|3����ߜ���˟���xrU�z��e����=���6��7����g����z�+�`�e�8��������>|��^�q��<�ʻ-}V���z�� ' cpe�T -� <>��������ߓl(�H���*��DB����z�s����5�r�w��m.̐��g��>zm}_}UO�UU�x�w��˔'VP��}��1K��S$\�&�Ī�@�,�����!�6.I]'F���n�}�>�������w�6Qt�e�]K�+4zQ��ӑ�0���U��ǃ���۬�̓�l��}�]��3���3m�
��?��s�;h�����l����� 7/v��qH9�'#���� �Ǘi:�Ә�M���%;]��A�ӄG7�Ȕoo+Gޏ{���r¼3���/�Z�`�5�PG��9fq��};G���S�%9a��@�U���7�]U
4O;�n�w�«̽��q���۽�9��/y}G��$�IA@PA�U$�x?w��{��9�j��EW�>���맩��U�� (x"uU�oA����P�q�7��}��d�'��2
B�<5������?y�<���s5��7���}��1׍�e���L��@�mk�wX�vwy��_�
9I�#����#��C�7~�6S;����0KF|差�޸�MM���L�81i��:��qe<�4���fi��������#2~�����Fm}��GdX�:L|:�~����U	�;	L�(Lu>���L�p���]�Ÿ�z���f C��u/	Ǹ���O����G����w�}�&�"'I>���s�G;�sJ�s:4�Y��a�2�[6�H2!����O&����ǣށ�>�{]�~��^M#���,��`��Mcm��m$���2'���ϾϾ�_��ɷ���#H�3��g��]� V\�C��O�iKL�S�U5�
�����}*�Zr��)�׎��S�(H�p���j�}��qx&pE��Gq��b��B�u�F쿉ƅ$}9y��>�l�. �4Č�c$�M�������7� &@���(�TAQPPE��0b*�I�����~y���q � ("'��������b"��T�d$��<���w�os9�ꕂW'JI�4�ή@�T:���A[Cz��/�L]w���%ʷ�������8:AaiZ638�SUU�_h�V�I�E�8�i0^��x S���F�?{����c驡R��=\���=Ǚ�҉j�f���JQ�mY�a  ��\��Gj�<��|ġ0�ۛ����{��36��q�'L�%C�?^g���?���
/P]u��7n?���*j�ZfY�e�k#&)�61���O:�y�#͗�p��nT�!;(��""ݽ������]&����:m.�E|�HHux��5��iK)������������6���.���q������~g���>8��=:g�Y��� �1���0�c$�_|���S��?�n����&�h��>[���V�b2�H'h�.���n�Z:K��D��c�1�&��u˖�c��G�ˤi���M��)�IU�y9�}�W37��̹"�XZZZ
�-T���=����О�K9N^>��r̨�Koa�9�Vf���iG�+�ˑc�l��W.����y��.���[!S��G�6��_�z��o��DX���G�=��$}�}˫:����VL�3u/IB���7ۻ���sI"i4�F?�����C����a�8v�h�A0��_\����{ޤ��J���V�"��Lk��%F2�<��l*��0Yx^\��͖�g���+.�)�Ν)�s��!��=�-� a�������]����VUD��C�M�F�<��F�N1���c�����0��{n�ә�뷦}I�m0�/��"#��U|�7�A�`�����f)K~s����w>���ў/��:���_��-2�zc�?Y��,錣GQn�j��SL�:�+R�|��RȌm�FF
���
�Y��Z�_}Myw���s��{$$zuV��h��'DwĂT�D�s�)�^����Ǜ�|�&1�*�s�_Sָ��h���-�-��Ln�ꮒ�E�SB�ˉL��Z�k\ˬ��Қ����\���G{�6ennI #��E4�A����wf�&��X�dWX���\�S���x�����B��wSX�Q���խ/�9�k����w[b��E84Z���T��uK��J�haPZ�rۙi�aF�f52�'��۵O;{�xS~hб���[.�¥�ʴn��������5�Y�ǀ@�G�4�Ӎ&�$���_��h̸3����"��qf�#7'�va�[u)l�K���5�3�K"I���,x�u	'vUt�h�Àd��aqi�#g���L�;����<81�g�Q��j�0b(�MtZ4b�v�9��:����)�C���5�M��V҂��I������w[�Faշ��k�����Hv-UU��vݸ�b�K���\)�k\�%f��Me2���ݮ[���LJ��q��S-���R���Ks.S����J�
�1<�_}��o_�Iuj�[v�ԏ�Z4�Ǵ݃vl$���B-�.m޽�)G�Lv��׹nm�g��L������tk2Ci_5ૌ�>���;F�)� ^����\���c��]H���ܺk�w^��I��{w`]+��]��	h���(ë���c��t�TU�÷�cΖ��ΠrKv�\�k�ء}�v�^=������D��Q��&�o3u��Jօs{/��I=���=���f�^o��iS�����Q�QwK�h���o��S�pl����U�7�����h�i�6N�b3���H�]��X�V���F���E���ʧ�/m�x���:�(��qx�eg'��`}�f<t|�����;��������r��^�� �C�ۅ�N��R�fwҭˆ\f�ژ����%:A�SqD,v_BK��g�҄}5���q�Km�"��. �  z� 'h�� 9���=�;���=�]����uUv��o ��۪{���`  �6�]-�[��U����9�P �y����A���>7|M� VP eS�uh N �Zڷ��y�( ����
���l ]�{z�]�en!�qmsV���W^����lV�;o��޽���+�սvs��{T<��b�Pf{_;��uOm�ӽ�w�n�          |�T    
�UR�    @ p���*��U��T[`        UT        T+( �Y��k�|:��~��_�Vt��F�m���4��=�u�o�)�<��Z�19ݛ��}������v�#�Z��^�p+(	�q���)Q��׻��8��m�n�5�wR�;kv�@     � P =������_u^V��s����m������H2$�7���hǧ�S�ވ����H��3�~�.�?��m�����fkNgv�>�9��tj4(	n��&��j�bF�,�����O��Y9]���G�x!mL�Y�8�Gڌ2
ڏV�^��7��ý���^
˗c�r��߸d1� s��j,	�fI�f�}�4<�͇�����#íʔ1eWA�D����8cm}-�_�����7 <���u��@���8�R��zO�D�A" ��'H{��ϻ�|�=u9��>V2:�H��Bx��oB�[	��ng��8��|Z���i�C興�!�o:�7�>�Jwp��xA	|DD:H�I0M,i1���=;��{��}�u��X��21�.[ ����|Z35ݫĻ�!��������G�㖂� �@ݲ�m�D�
Ϲ����?@��v�j����2k�q`�.�_)ݫz��C��94Ǜz�䬭E4����c|��%E�5h�~9l���&�Tf�j�ha��/u7��Ф]9��'W��\���ʚ��+�IZr�-����#ힽ�yQ���j�{�*̫�=Kx���z3"7��_Ed��F8�S%����"�����2�Y��ַ]C�Y���S̹!��[�&�~�����eO/�����L��ػ�p��$I�*A�^���{�n��UVG���y�	B��aZ�c�8n�}�V%٩eVϣ���{��OJc�����rA��]O�X{���ޚ�]��w;��7Nr���V·�=��muv�߾f��}��E�`:v'v.��[甠jQ>���PU����WR��f�Ins�3�<�:���6�>r�`Y0jՅA��<����d����=�vǮ�bU�+:�LL\��Dx��z.;���M�F��_<��I��a�F��^=���e�b_c��8}���03@2�&MfV�9XC舍8��y|��m'�3Jf�b�2���y;��̈́i�]��D�w{-�^$�-6Ri�� `��m�m$�#ga/�����b��n��i5ιm�ﹲ~��D���X��ԥ�f�ǽ�!���KO�"��hh���zB��乮x�)%4�貨��vu7�e�m�/��i�&,-%)�?G����VJ08�4!����ޠ�g��`��.�
�u��G¢�y�pwґ�5e��ےDG���K[Ai�}CJ
�\��?{���8��yB����}�d*�I3x"��t��^��c$�%�S���μ��:q���9=�e��,��,R���`#��NK����[�?w�;(���E^�J�RIHa���N�&�����4�2��wܲ�\�@�62�WDz)}�k�ȄSK&�Q ��.,���\�n���������:�M]LX�Ha�����Q�&'J���SBo�qX�zd�νe�J�w`�۸T�����d԰A�v}�}����a��^'�Oqt_T��C��u�$�~��Յ�$�v)�4�����]n=γ�_�=���w�Y�G�e~'4�eT�PW�}�}��Q?��4��1�\�#;u�E#��1zX�NA�`���>�?�[406�2�/��C��DD��t��֞'���j��\:lK�ӥ��tf�֕�ϗ.�B7���f�;�`&Ԕb9�9��̟��r��oъ�r����3�RW��L�h��ɍU?#���|��{/��c��bc7�%e>i�g��F���0�����"�`#h�`~�ÙJ���$���
@�ɝ�1|��pv�L;�񇀝TPS8���!�f��{�C���|;�:p�H�ҍI&)��ƵG.l�� +)����YM��`�k���ǞVR��w�U����|}c @ �<�
l    <!��~��}����7 ��ݷ�k���¨��5� }� ���/NNw{��\�U_���l���'೘�,�̇�lH�9U4>�DmV
\��2z����x&d<�Y˛!oW���<Pд�k_
�w!��ߎ�x��u�RI5��|9K�s�歶��m��HHn߿v *���{��|+����>)��˩���y�{\�ne���Nqc�ۮ'ޢc�!��죞�Rm;05���W|��j�??��Q���e��w~7�iu�n��L�n뻝��o��o�?�IfE��E��q;D�&m3E�U1Z�Z��J�i��w����{�ʰ@*m���?�fB���,縁�������ki<m�����
�ݧ�\���wM��^9�{�u�C�%��j���gD�5U=�����=��~�3g�fƵ�hJ4k�1��-�zi����<@�`�����#I�$� +�*�����<�W�X�kvd���R�JBU�l�~�t�أQ⺳3�W}�u��"jr��7Ly��LñR쨲Y�8G��T����Dz#�1��}���&��/�t̙8��z#Q�Gh�}{M�hձ r�}ۉ5��s&`^�(.svZw�6H�(�Ù�%	��&M�Q�ز��Z��[}�N�DV[�B�x_9уN�MmM�d>I��M�����[(&<�Iک2nD!��_G��=��x0�߇����X�X��$[|�=�sS;� �c����p�����<�.�t�֮s��݇Oj
��r"�ƈw�t@�1$�i:�Co���?���N�<:�ڦ;_��z��G���g3�v�'�r�����K<Kg��~c{��%��b�!v���mR��ut�����u�sӹ9@0�*���M��}U'�b��nK9��h��ɍ��Z�dMd/�,$����R'�<P~
��i�q��,a\�3������w���/��Tp_M�3�������`�6ԥ5�$�����.Lޜ�^�,��-O��KY]��m�v�2u7�̆MQ�9fo'ɼ�}��ܟ�;G�}�"r�֥ �����Kw�]g9羀H �"��3]��߹�xܺ��}��9���R� p��.�f6ڃB�8���%��b�&�a�\r�}��ٹ��Z����mv�UxU8�@��|�YO^��:z4U)V-��6�fȷ]�_U����v-��=���x�rj���ҀF�z#>�z� U���s����V�F82X�1K�dr��+D6�F˛df��=`���V@40��X ��2���H��WߨO��>s��;�r��S�xv�q|E��j@�E��mO��)����{gi�k|���4�^��P���Y!�3����߾�뛳�P$<`E)"2���+��U�+ �Z��0�aE� ""T����W�d���,Gk���ٹ]vu��� *B��e�ș,�J�;}��Xw��k3�/��Q����Ag��=��^.FKYs�]����P�5%nOmKoj;:�Ƨ?DE���g
�G����&�N�$�򘸩�%-'���u��U}n޼�:*��Q�wn��"�J�*ul�wTs�G2�z��:o�,�1ÑŃc9�!�����:�S�d���{�9�o^WY�+���v��jAgEy9=('3��&"�TM��Yi�V��<N�w%[��f�a����^�lV���K����t���O�gGF���_0b�W��&hc=<މ�pw �D��s�4����������H8�/��(�z2f:���.�_ ������D�9�6�N�����.�=A�)�v`��c	�li�S/�{t�5���5���˜,�
��G�n�njC�7���޺^���J��EW������w�wxp�d�x/&����?9�� ks�Pڙ9�|6����ڪg���̼�޹����졅ʧ�ql�P^�����Y��Un�]۷uִ*�n��   �TU��   �}�}���~����m���+�Ի^�$�E$�m�^K42՞�jx�~��{g޷�W~�^�y�$?�1OhX,DD}7?d�{�|��ߩzgeŲ�업NMN:q�/���0P?ן[g���O� yjt��{�V��6�Sa?G�!��#��^5צ~��4l�UUF�<qZ��7ȫH��n�*U+!��Rb���R�� 6`,�^s�eϽ�>V���-S����'���_��������Fo���]k��Ʀ�q:�1�<��ܙ���^䓴���]U�+v����4��(���������ңn��|H�U�g�6���C����n��d�SJ#��F�)Kf[����Z����{"�©��uvd���]xghx��c�,֝�3&N@�s1)�yѦ�6i��*bY�����h5Rl��˜��3=�f�0���MwZ�3�_uņ,�����9ı{|�ϧ�*S�������]����dt�n��Ӟ�W�����||-z�ReЮX"z�-�0�Z1�:S&����1۟zfTq-b���THXb��������}�z#�?G�yx̗�}�)ݮ����X �'��	ڱ��G,C����w7�������c�]i<%�E4#��Ԫ�WىC��yR��k�Y�� ��ba�R�����9>��ӓǮ�{��:��;�����H|s��Bl��?s����}��is-h�$~I�i$m$�"� �Y�Q]�ӏ+9�ީ`�꠻v�l��K��W�1����3y'�p�7����8�cǛ�L��{��zfu�b�/x��~c�yb0�s����=��9���r��>�\��a$'�c��߯�o=��˭�k�(����~氦8��=so�!�j;���l7�r���>;޳y�5SZ�.�I�.��������0MaC[
3F��[+j�e4m�+�s]����9�:�i�S
]V����w�)�ߚ���8�6rG���	|i�sE��_5�l��.�D����Z�.3�ƥ�?�7��N�X����>̬ 	f�ҿ��I��$qYn���x�gY������E�0�y�y��)	�Pv���ON��"U�[����pa �xsMc6�k���rV𒒈G3=�,:�;�^�σ�*"������$��dn�l��_3�7�^`���D��Z�ę�S߮��}y�[�[��	�w�&���]]�J���Umk�m�J����\J���3�n�---.[�������q����ˊ��ִ��r�i2��
[�b�t(�X����D�m�X�q�1:�u��9䟶��p�F�aT�i��Gr�S���XNh{�`�ۢe&iq{���=K��V�#gN��蟽n5��iw�Zr��ݝ��n�MΗ<'�w�˘�ʸE��t������[�&�&vr�ͼ�=�j�������4��"���=vzl�4�i�0ݫ�i� �/�$^���*���.9|T��{nAX�q,�TqP�`̋O,f��q�ʙx)���O���O�Y�y�۱�Y+1����]���t,L��y,�7�l:��ԁ��{�4�$��wf�ִm�ۃ��ů)��7R����3��s+��k1��D;�������;�᡾Dj/p_�L}�g���v"�{��4U�o�A7h�6��n[�Y�Iɀb,�n_,�(e��^M�f�v�Q�wd�#�g�otu	8N�Q���dz��i�Y�̰�slᡬ#z�eKG�1ec����*8���dqMw�)]��V��U�m\��g�̳��$P��ͨ1n�q�{�N}$�WY\���.�$�[9xD�1è��켇,���'aS��٥�o9�<R9y��lr�Sy+���el����F(��߫z�yr��H�&{%��☡�Rd�9ZgϜ�AH9tX�)��]_Y�F0����j��~�d�dR(���H0����fw鏁�����J�����>ϕ�Z�6�+ץ���I�/ 6�'��G��$=?���
S��p���:8Zr%�ޞOM<�~���|�^�I^�2����C��}P8%�(ɶh�k�sΪNy�F�"4c%�5��j��ФgG����'}��,���Ͻ�Q�뺇*�����~�l�7�,��`ճ�-X9j&^us�0��.����'j��w�qx�ζ���qF�;YOhMVKSe�.\Wmr����ST��UM�]��5�10s^�}y�Ysbȼ�L�4�c��v�:�R�=�cG+.���S�s��w�]����L䐚`��B��_,X@����g�;����oY����N�nW*ۡD@<DC��q�	;�Ia��Ll,��K7:���C��8vY��~�|R0��m�U���b���-:{5T��F8;9������3���7r�Ha�L���ϵ>p���7��{i\����Q�Dzo��l���������	�1��4��R������+�9�[wNO2�ʞdM�S^����N8#�Z��(��G����p����}��P窨@�Bق��Zò-�ŽQ��\7�Y��8�$Xo����u��9ʜ�7�؝������{���=��1�����֎�������������i�T�|q�6���V����!�ݡ��R�s��yu����+�gy� (�EQE ����+������ϼ�\v/��b�R�$+r����p٭�ݫ$�mf	�f�0��"�Feݬ���W��sn�NoY<hIW��2
�-={��[|��v�vܑꞻ-���0 ��P0     y9����߿����y�9�e�v��TUL̈SF*}��(��l��?O:\��x��x�+���#.��g	d��p�,Q��>΋j4����s̾��3_j{M�}���@������CG��=P��p�d-�v�LG�=�s����iY�p��� �$��fq���e��99�����Y���#�:6����K��2����u�7�2��t��>[���)_��8�3���CS��I̙����%����r��}t����F�-i�{��Ug`��n��mˌ�K�p�Nv���}�W�}.�)KcQ��,'ݍ�u'�}���F>�������m�	IcM�16��`£�ׂݷ���?߲D �1�26��q��6�h�37�P�k6��nVm�h��K9*C=&'�|��3}����ԛ��8v=�ō�"����Z��NHC�!� ��}�fs��I�w�Qμ��JQȋ�g�Nt4:�v9ٺ1h'�Q�)�K;p�7:w�=A�#�q�Y����:<R��0F��H��WY��Tc��G][�����")	�z��-�Z?L8���i���n�Dtq�ؓ�[1ss94UL��i�R�
�%8�l9]�Z�Ʒ6���rcQ9��n)Ʀ �b��kX�S�)�义)jFd���5]�D�UR'P%���M&�]�����i�9�8o�"+���<7�v��S�^{�Ս��8Jv�k;z��� ���pvH��i$m$�x�m���?zB�}3f�
偮��{(E�̏F=��3߻�y$��I0�]o����g����<�s��632��͂��6�p4�ʎgj���:�I�.��5/F������,a((ڙ�L��x����Ju���O�U س�f��7��{��s���M��.��a�>X�(
�*�FPePXƭ-�-����,���X�%e)R��[*�����`�
ؠ��u�t���e�nL�(󄉮��q�p7��Qm��X����*\9{p13CSmI^D�'�h'���^��~:�J὘Q�B��I�����uvO���n�>j�Ҧ�/�Je�vj�B
0�᫯�sl[Ow}�����is	^���Ɲ���3(L>��A���韾?sV�ڷ)�)�Y$u�j�Y]oh�t{+���]jP��p����;7{[w��U?�|��˛�o�[�6�݆�������'ʦ>��q��DGƞǽ�MG�5�����G�)���
a'��[�n:����mdgq&��D������	�璘؍�W:��dҧ�%i'ET2�lM�os�3L��!6��W�kq/k�+j�iW�TE}�?���􏍿����G�/��"K�+^ά�Z��^�ɞT_u����y���G����}�̬��������9�pnf<��pV��ۧ]A���f�aǯ&�(��s�۰�'¹�k��"3��������4�w�(�//�l��*@B��ܽ�n��3�O�)�s�ӿ��3j^��v�p�ه�3q苼��;���~[�E�g�ۻ�T���!K�y����#�����=����k����ل"�4\���o���<��#�Ha#%	1+K��2N,+O�K�I�!Z�/�w�0nrI��λ7�"I�0�Y2����ι���6����-'�~��������T*H��� 
���V�^��׶�>�B�@�u������Z++��4���R�]���d�F���|�@L@vNUI�~�H���}N�.�+�/���R>�?U]��\����|���+��{J��}Z�Oh� UT�n�3J	&V�C��]�]{Y=��T�'�'��pΣN�|>49��޾�W�y���j��� �Y ��DB<�* 
�x�#�	��~+a��͔u]M�]D�Z�v��c#Fu{Su9�XA�w��o��(��l�@����lZ�@��Ocj���XuK��W���>|��-�z��S�b6�0 0�;�
�SeP   �߿����������nAm{�zu�QU�*��6��m��=c��j�b��r!m�6�b{�8W������;_X�X��w�qܡ�L�f^f`ȫ����#=	�&��\s�Y�:3g:≰��f$pRNܢ\
]Vb��=m�tg9�oN=H4kbb=�~�a�B�u��u����ܗ���vPXnh��2��f�<N��ͼ�ђi���XkQ�Y0	�x��Rg$d��ot��+�'��;0�I��6��+��i��a���ݮ�MV,͘b�Z��@qD�H����!	�r�*f;�g��H�c"�(�
�ddR �F,AAT"���������p��S��3�����+�E��>�R�9�����Ϊ:��t;�߁� v��$��Hm��z�)G�5��،&O�5T��������D�}v��6��4#���H�b�:��st��uw>�3;~�/�s����-�;�;���t�e[k�f�*�&��Nu�q"�{:��b�H���鴖�$� ��,��H��8p!��u�bT����DYQ�D7&7������U��3����:Q�����Yp��RvB�L>(g7R�V�7���\��5<`
�(��N�xtn���Fh���Ѭ�:~����Clo��vu��Y��t�P"�3��Fu�vu���994�K��ۙ��O^������o�;<��$�){F�vE�wO���LR[[�{�˳�yOӂo �]ˌxry��Oğ$jH��H�Pl, �m�E���$�c��׮��o���������gW����W+7�4B��Y��쾷x���*e���KO�@�Dz'����f!��G�>���T��$��I��;r�m��Of�'~sˏ�m7^�32������e�U@قۭ�/g�t�u�h���͋;���-{]_���\nZ��5�#&�<��lz�2v��3�;RS�?V�����w�?��;����]0/:�01�"Ѹ���L>T�>���%(=%��C��d�n�l��^Q�%�o=r�芑y=Ǡn�TzOL�� ���<��}Z��ʸI�1�s(�1�k��礘h�Y]=J[1L��T�|wa=?z3�+~������������[G
׺֚�r^�����A�4�A��� $���&!y����n�R�ˋ3�Y������ �ޒ-L�L�h�� �xv$
��ސ1O�Ӿ���=�6Mʎ�������-ڧ]�댣��K��1����u=U��r�r��֠+ʕ3
�-��F���D�.| �d}���Շ�+ꮼ��Ώ'��s�=��^^V���}o�[b�ͮ�N��� G����q��U+����u�B�[>�b�ZT�PF��GW��6�wl��{�,������1�JMM��RL�K`��{Z60�����f��֖��rױ�Wf&�Z�V*t�7s9uA��ԻNw�6�n����^ދ�B��V奷]fM	����n�On��S�g%T�#/Sɷpz$2�cZVCHU�9����Qu7�ib�*r���{��@�#��n���.��E}2ߙ��Q����w��ٹ	�Z����S�:��W��q�/i�[��}���MQ���kq�fJv�ޝs�3?vw8��/3��-?"��ҍ�I����a ����Z>��|!�.k�y���{��<�w�'�������9�fʞ�S�ݕn�<������|���1t<��h������N�o�+t��nvgt`��~ٹ�@Ǩ���ۆ&�ߙ����A]%TPZ[�]��[q[n8`f	�4.��v>V��K�������1\��e
($�<�AVqf�����F�h�Y�橎�����Yr�շP�/�7�e�/0��4[~ �~ƀ�9KҴɇ�E�e�х����^�, ���DI�4�!����QK�I��5��i�a8��Md68.M_#V�`ds#��d$�#�e��1`�����I�x�d�ؽ=�9�ŝ�,c6hT#u�0f������>��u<�~Dϊ����8�˞:�*\8>�?gM�M��ʞ�w�\e����5���f�X���R�ap�e����3��� ��)�@��I�����Y�CwGH]��E�������{�M=u��glg�P&��U@�;z᫁����ܰgj��Ѡb4	�vJ�w)��n3y���Q��6n�ݑ7,_ͨ���pѴ�G�/C�]�	sv���t�q����H�ݺPN6X٪�f�\�_W>ٟ�^��L-*Sr��2�����w��$úɂdˏ����=[��n؉��E�ۋ��!8_{��uygV8	��J��9�ii,��qrBM?j���ص����y=#��gb�,��O�Odm��]��ݻa}/���,��ҳ������q<��:w�+�rѶx̝}t�[��n~~�ɩLk��5;bb�51Wv��i�T�5cye�����7�5���*x�Ӡ��Z�ח/`�8;�z(8�O��I��]����:Ԧɩ[)�;C%��R�����B ���%�^6�m��N*��8@z�hUj1�sw��w]�x� �1�/P {`un��Uz����w< < ���6�]Ų*��1�sq���UP �w<����Tp��[*��ʜǀ7���8�  s��۵G�Il� =��쬪�ym�[�� ���{m�v�*�
l:j�u��ٮ�8 ;�/W^�޷��m�>����l��7wy�+'\�w�U���W/d      QT � �e8     gT �T    UU*�	��(n��t@                    �6�m��a��M��h�%��Zn�;-�ؕ�X��!qoP�mVr&J��3�-����}xvU�%-i��m��w5�J��`�c�ᶋJ��)ݽ��U⶷��E��C+/AӼ� 8;� �`    ;����~~|�����U�ښ��z�W{�S���3w�W+NOݖ�U����_�M���@����ϳ����6�ϧ�2&ͨ#K⣓�33t-�Gu`E�AM����s.�R�b�2�v��B������ꟓ��t����T��2����&��N���f:̹l��-!2�{2�Lz/��W�"��S�鉲̦�����о�lw
�F#�Gi.8'U\{
��gΧ;�9�%�7�q�k�XD��y�t�2�A+�Ƚ��c�S
�a���5�x`
�Q�H�5�2:f�����;�S�9�z�Aʓe�M�󄆲�)o�G'��ٛ�}O�?���嵁g^�N{���<B�d&!�ܱ���o�?�Z�8KA��E��=��Z�#u�nQ���f&�1Vs�u
_#��9SO@%BnFi�^yk�۷���$&�F"� i�W���uwExV9{uMR�%Ȥzbu���3M9�j��e�F`]1N������1��k��^���P���E�}ď��y��q���n��Ί�f�ey�讃UXH�MP�t�[�Wu8��d����,U�&�DC�'Z�����L�@��q����ϔI:r��SU"m �QI�w�풌'RA�s�= �+zX�93*~��@yU�+��'����L�z�'R2%�����.��óH�`	�:�OC�q�mP� {��;��*��!6��a�w<u���5����������׻��׽wt�Uw��-]�*�i��&�1Ks2�� 	ޜsD�59��|�����M���\�2̶Η�1�֖�*<�X����wD7�X6�.�ƚj��u����z!��{s�ߊ򹎜�'Y�_}Ly�k�,夺X�6��sH?�b�C�ԏ�������_|�@}�Y����%������D�M0p[%�;[���;�e�U�FK����CSoc����e�E�}Ӆ�-�z�� �����xv����w��v3~�}NZr>��tI���穭��|�#
�.����u���dGC��.�o}�D@�y�W=��OdG��� r�X��~�dd��/SZl��>�P��uR�{p[�N���v�  h��S�apȲ�j�L�)���9=�_.�Mr���8�s@��=�v:�&��Ë&�-C}��Q���	�7Y["_`��;�e���q{�����xxDzq���|�|����I3Uɍ[]T�Xf� �\�o9.{+��8���s§q�X�^𬻲-=�l�$My.�x�x�'���G&Le�`w� {ޔ��E" Kk��ϻ�����D��lổ(�u Ȑ�ݫ��G���{gd��knG�er�H<�{$�r�nNN���T7F:���$Y�z�a\{ޏ<���|"""�~�8�f:nb��r��'<�o�z��X��V+��0�����������`��=�����������2k�hLgm�V��;�v��C�O��_+��k+%gݍJ�MLu	�'b۾� UP�u���q3�N=�Ue6����Ik�c�V�W۱�q��ǝ���!Ɠ���㏛`�pzõ�)V��`w�&��w/����}:]��<�}ݺs�a�Z�w�J$�
�5�7z��7q"���x1�ʺ���V&�뮎<�9��*t��5?8��m:�4.o�:�j�U4g-�.��qW0qs����Ӟz���3����|O� 1 �)��}TW�R�y�O��n�W�-�:�K���m��v��ӧ�c]:�>��k|���[��� �eS���x� y-�[4:j �<�r�T+=�V����cu�@  < �UR�   <&￿�ߟ����%���k�����a�W�SC颵Cز��X���M�&���vo��Y;�}d�i����)U�O*�no��b��N����E�V>�w%o�E�w>q]�P�wU��ܜ9���\��Wuٴ�[��v�?\����p�ǜV�q����ù�6�%vVD�$�,E"��E֊mg(磦���ϼ�������Ǯ�{SFAR1Q�N�Tpo�5�����j�I^��2�ۛ
(�S�lڐO�����o�OR<q%Ae�=���k^� U5��ݭ����q�5���Z�T�e8�/p��N�\����ff���o�L=~�wh��}��o��,$E�X�VEX
'�eQ"�h���I�=�GE�Խ��קn{+گ�u��^����yʐ��ۭ�z��{:�%��si!�ܻ�ܴ��X���e-���7���/��r�ȑ0%�C�Űw��N�T��&�9T��!�b��;!�&��[u�Z�Q��yfe}�}_z�sӏz���=�SQr�i�O����l
��ޚ��^uiVT��$Тhk`6N�x�%��gg}��~������_GQ�ru��� �ڙ����f	M1�i$m$�)�C���|�K���'�+gcqf=+�ܐ��A�^��Z�y�����ۜ��W^2��"��MX˹�,����
�Ӛ������w��������NSf�f
��$/�d.��K�\+9ms�ܽD1�( (P��gv��v')%�qE�ˍm���բ$w�[ӱ�����t�[��Rj�j��8�������{!u=E�7��|Л�fK����DC�������mc���r^gpf����-3�T��g��?)yac~�8���Z�}�vAq�F�fLT9��\�c������d[f�c)n��c�*�S��/+���yz���~�:�=ͶϬY]�Sb!L�DD	H�m�.B������˿Gt�߫����h�\��Jt�뮃��+cL21ԃ&\�qK���m;VT����\3��~$٥3˯����9���m�m���w�����y�f��w�g��=���l���!�� g;��S�Z�̿��	L��3�������
QK+�Nh�F�7���D�s��G� |=�wq��]舍��zƢkʻ{��am��w�gy���u�X+)�L܍>������A���Gn����DZۧj�Eȗ����z/�[���6�x�����[��7�9Q�}�~[�|����]v���fk$�d��y�S�*�8�Cy�`��#�WV,�����SN��E����|.@-+�#�ᐴ>��{�rHUVO�yt�WNe�1����}f]\7��֬=j��|�;d�j���<ݎҵc�R_�=�����s�ZR�?��˜����:�����pO9��2�8�e�w[�I�<$�y5/:H��_^g�3��}�j�Os�)-��R�FF�	�#fp�6���;�N�=]m��RW���:�{��D�:��w��w������刺2
�� �"���g��*�:8k��,w�S��v���Q�b!����̻�:��������l(�m�E��ƒe��޶�����<��
�0Zg�^;��M9�:[m�FݓǔPc ǅP��   ��v����~����R��lY�tV��U�S�y|誡3+�=MX��S��������;+oUB��7�"n��{c�IzR��&;��Λ*�NMOb�tr(��P���^q�����W�c�oj^k�W��.eD�3$By��}u�cn����h4����7lWI��C�m��M�cHUF��LeJƟ����Í[��Y��a�i}���w,���R7c)V�P�Ѧd�f�t������@�=_������No�Q�PS�qx�Do�ZC�2��Y��Z�u�M
��553Q��׷p���*��sw~|�>��Y֛i:��W�es?3V���
�r+�T%�<��ǩ@�u$Ȭ�����+�I1!U�)����O<.y��w��'�j�/��̮��˽�S\̘S�Ӗ���Y�37N��ިam�[����sߵ�:�" �"

`��E��y��]vz����>���p�VpLu�z��_�ru���zyҳ�:����;�[?F��
>�_T�$`����;�[��l�=z�z�Huðz��@�k�U��t�*UMG����ȣ3Q<�'o��\j�s�ϑ3;2.��̻n�層'o)���F��"f���u3@;�O��Ww���y��r3��?`�Ԗ¸�;Y�N�ޜo]��u�.��1D7���͛���˛�5�\�`o���>��>����`lvC@��5׋Z�S�{�i<��V�n꺓��E̠}�Jcm ���K�ĆR�QX`V�f�:ְ�s2��a��Ry�LUF0F47#��pB�}LI4Qi����6��kslNE!KL�3Lx�o�7፡�8O�h�?eg=��R��}���*��1T��L/����`�E����%���.�w�<�����UͰMXI!bI�D�M�� q�ά�ޝ 0<2l0˻��u�{"87Kp\Ni��6[t����γ;�]����t�S�U�e�*�"���?�?���x��A�_o����EP��ћ��MZZ
�c�-*��Z��U�&&u��en���)ӱ�D�*���sty�^����ۑjw2�f���hݕ���ΗM373y�gFj����r_$i����ٝ!mEP�f���x��m]?n*h��7����T~�m����T8֡zv�G5�]�^��[I��1�XgPܔX�D�{:�	�Y��:<�p�-�9��*iT����<��\�Y{��Y�,^�M�8���	/��pGoh�P�F�lCvu�H��CF�(D�������*��8� ��c��I��\�8��Z�^���0�+vK�Q���A��<P���N};V�y�YH<���$D^~Ǫ\+��9�cm-G���<=gZs+���8QN1�H�*�;i�N'�{=��E��}��>��]�HٷC���]o�1ݣ�}�yiX�f����q�Z�{C�Л@��|��EI��e�&���ʗ�^SqL�xm�Of���h
�����1�s��ll�i����=lj�<TՎ\c��� ��k���,]�L��9�x�~P<\�+��UH��bg��bz��',�mK�y��v���w�'|3�7{���!g�Ŋ��=���dI�K�Y{n�*��`�.�ii�����v&��.d^�|��o}�?������?��6�[h�ٞ�$�i$�ě���e*o	��Ưߏ��d�KS;ܚ�w�)bJZ7�d����[�f��{ޏ�G�g�����>F"#����W�����'w&�ڋ����=5b�N��N�,z�c[�&*@� 2{guk����;S�_tf�����˝�i�#e,��C1[x��wn�j�}�I�f�����Z��藦&g2���^�V���>��}Ws��o"#Ѕ|�Um?U>��xm@6���ʬ��+.�Hk3U<M�Ӌy48T�������x�=;W{R-��hSAjd�U�t\_kcu�ajGt7��m7n�vmb�$�I}t銭��e���A��+����7��i)����U�S*Lؿ��d[p�'\U�یbue�����������Z�%oV��P�(��
���G|U��f���{�uv�'/��N�R��oG�wͿ��ܷ�5;ߔ�؄KU	L[����"��S-Ӆ=�:�yrV�<�s�-�#s�p�c�*�j=�
�U\<3��|�zrvܢ����v��[�޴!��6�$��O���h��2ꉩ����ܙB+�S�������ʠ�|��r@8�Ύ��ǀƜ(��Oޏ@��" DU,�lDZ�E�,����R�*UVV�U���P��B�UZ"T���g�ο�M+�T��Ѩ/Yٗ'#z	w�mGr���[3&�t�Ss�kz���7��+���j�Z�įk���sa��S��q� �P��^�Y�}%�R�-����뛚��T�  �� @�m����G���{O�m�HG
 YH&�I<l��ć�$D�w�w�R�&�'L@!%��ߏ�lw}o��[�kV�Z���l�8y�e�]�5U�gd��c�n�gw.������N��q�F5����&��}-Vʬ�Fh�_���iG]�w/��������V��]9�؉��G�ވޏ|�Ѫu���Ψ�隀~v�T]K����{l��N��+Cն�4ջ6���36��ոz�ە!tiW3T�m'�H��Y� �S��0����X~���з����`������Ii�m6�!��T*��S��ϥ�o�������������|�=*�R��ڵ�u�����{Q��v��T�;@�[`�SU���$��H �?yy����<�7�����	MLr��ʺo=̖�j�J�'�k��u���H��ogsK,����|�W�s;S�t�w<⬪w�K�r�X�Y��"b�t�\��E��j�����~�z#�ۺE�e쐞����k�����x��Gl-OMkTk횝OX��g.�lbY���|Z.�#�xs�雴~(�������� �m���Gv��Z[��k:ܙa�����CE����y�ߌ��6��}�1&Ĉ�B�e�^]�B���Z�U�ߖ�w��o��}��f�s=�{K�|B�YaP�z��W9{y���P{��Or:��碖{�C�U;��v�1�j�!Ofg`}����X81�b�D��(S����e�?cɜ5�L���VU�߶�s'�SF�m�D���o�s����'̐�A`�������!i`8-X�lya]WY�
�AϦ�U��6���2�
�4gH�*3w�+w/6 n���):6��
e�0�mV���
-�I9A���Y�V��2gE�B>���U,V��W�����%Y�{iQ"t���>Z�|�����Q��"���Ǌ9��%��I�Ž}�BO5�u�}��w�z���$?!�_�x�1!�svA��rzu�xV�~"��o���y���[m�m�*�b U]�p������7��92�n�����n�(��`��r浨�Fd�{�:�J|��ʙ"1�f��a��by�\�.z��S��	o'��B �$ 9CwA�N�`�������ߋ
���&���o��ⷭ�7�@{�w&a�d72J I/GK��Fp�8�Z�o3޷=Y�c<-����AJFӫGj��k�"����2wp�y^ge��>���w�%9����;�"����r������T�7筠R�����2�3g���V��	LVĥs��un��uEF�s�{���y�+�4#�8���'x-�;��6�����y��x��k�g�� 	���l�r]�1b�Vr�����iM��Ħ��33��sa�� %�߿~��|%SM�J8[X�CH��ML�
2k�Y.`�Nږ�n>|>s�.�ʗ�1����\��Y����2,;`mk��16X
�5FhQ�:�X	�t��f���m[}�,���h����RF(�"���Qb����ߢ�K��p;��F`a�|�:�=c���.�K�<߬v�[N���{�)^��c�Ϋ���^l�v7�m����5R���:��4�ρ5E���=�SRN��/&x��q-��;��-U�O���.�@!v�(җ*�3�7����u��0�=舞�p5�;��7f�iaU`�Vo_eF`T�)Ng�֠��,h�Y[Ot�Π��*��o톃��L�}|��O�1R���B�Ľ�:��D1p��q���I�\��0���[w���Foojx`if�yU-��^ׯ�P�U*m�uwWwu�[���r�   0 w5P   m��;���Q�u��&�I?�Dm�i����2l���~> p�܇d��Tb�L�,3���|4���²����i����\�%��ˍ�iL���~��f\���>$$����>8]<�X�}�Gٚ�_}/W3�;��w��>����+��#M�x�'���l���G3/A5<tZ+���',3A��L���$4mQ�&)��}��U���;4��>.^��K��T�n��K�u���S'RȪދ��[*kbx}`��A�z�����"���;x���]Y�v�ޞ4ܡ̽1��FT�2���Ue�-��Kd8�5���J�8fP��{�]brz[�8�b��|clq��N�����ׯ�H���-&�e6�oI%�4����{t�N���١ƽ��l�t[�I�Ҵ���?c���۽i�m��g�_7IGCC�\���y��:lЅf��	���Y>���@�'Nĳͬ�V9��&��u�������"�����H�Ň�B	�bg���4��{��v���v��Y4l�[<(�4pi�t�벬냕�Q�3%X�hMT</���̬3
�'�S���^V�Mk��<�L��ŒB�h3UQ3�c��7�G@�G6)�ɍ�s29H������640��Qhd�s»�ud���P�R�O��w0Ł���X=��(|�����sv�Q�J��Qyҙ��cgh�#�T9�2�Ő�w�[�r��T�N�Z�T��h���>�N%ԏ�����p}�9s1ϻ�Z���O}SnL�u�,�G�¼��0���NWMޟ^A����[�ĝ\=�Mڵ��p-n�t��F��tC9;������{j��mz���:��R������b�3P�1rPL����}�|F}����d{�&�|�c���۾ǻEA�����W��_Rj�9G.R��-��p��tKɝ+��UL햏�W	��=������L+ "�Lv<���!B瘜��2^���J�Huﱣ���GGIn�7B�;�R���a��uՏ�\}:j�bi����{2�#`w�bF�+T��V��dRe�T�2���=@�\�I���_��u�Y�;'\�'��qC��6�H�Iqh m�G~ދa��K�?3^�dL�:V����hDr}8 �<�skycX\98�L�gE�C۪�b�g6a�y�I�%���s�&sy��A��3�B?�Fx�)3�<(���V��ltu�ı���ON�z�J�\�B�Cuᑡ�fc�̞����s �;�j������_����(k4�/��p�)����=3�M�gi�<i��q�8
���@�����c0�k|o_?x��\*����(q�?�C��:��V�1[8Y����Q��c��=�a�}4�'��/d�w;���r�L�����RP3,�H����|�I�\��S�0�{67�j��KF2-ɦ~�ȏDE��C^�5\��,��&*��Nm��v�pS�����y�Ӟ۹3�߈�O�Ӵ3=��a��;xާ���:y�%;M=,�l��IJ�"n*~�(k�m��ىf�_�_4��=1y��\N��S�a[;o����Ʉ�ߴf^�ԓ�g�2:ِn5lM��#�c��}��JNcD����-2�q����E�=<B�2�۱�@�Nn�Q���6]���t�ɩ��}��uxc��M��w��q&0&���3��2�œ@i�d����xfvw���M��$�1�uT�/����G�ٰ�46Nӈ�� �+[�5��!f�I��f���c����Q�/&���y�o�y���g!����bR�{��3z��5s+�`,L�b��`:�J�*%�3
WI�(��H��LY��d�	˔ѭK�r�g�5�0Q�o5)�W����6^I�4sM>}3I�:�ji3rĆ�R�[I�.B�e�D�G�u��z��q��-�
W�r�k*����$�X��I#�o�n�-��}[/�'�sf�5g�|�$8���u��r�Ú�w̘�2���T��l���{��� �U��iVh���Ӕ�Pes����Yx�����=J� R6��� CF�?ekG^�:켈��ʨ��0f򹰉"T�}t}��;������y��Z�`�=��`��'�f�����2s[�{����ܮ̥�LZU��<���/vm�?RV0���x�,f$G<�T��/{����nR����7.8��e��X�۬�s �m�\	�[t�M���M��7W1Dq��e��(P���R�����K���f�i#���1e�uG�%Z����-ay3�)�X�N��7ɱ�a��Qo�Y����<�z�:iMX^uˬ6��̐\n>Њ�i���w,����J�Nԫ�sdy4��.e��b����<�k��0�䇏]��v����c��"�'���g���'x��C��b�2���V�k�?[xǽ�Q�
����:�H���ƛ��y�����)c�k0;�<Gq%��u5e����9OQ�؂��u.�%z/g4���Xɷg�^�§,�h'.��U����0�$�-c�C��arxz����2�.��'%}���� �)��^��/i\���\�F'�b�ѿ??��ӻ�~^.��y��akk��p�d*F�����۵���>G��/k2(c�Z^��+�W��Z`O�ח(Ҋ$nwj�\p��I�ݫ}0͆�n�"�$�KA"�m��J�U ��,�Ez����Uny���޽���[/<ol0nW��ĜT�������C ��� ;��M��� ���n� ��z��x�[<���`P U
���V�*�ܛi�P���������guK( �w����2^��qT����;�nzzқm�������g���[U��v���M���/����@
��y���������]  x    � N ��  yT   U     � ��R�P*�(؛m� �e  
�     �P          ol�m��d�	$o�9������h�@��fH��;���gapc;Yj�&y�Gr�M�bj��JC�m�Amܞ�6�Se��*<�@yY,��3۞J��{VV�������s� I�p*���l    ;�����������>�.�n��'\nu���$�`&L|��~�X��Խ���Sē�f�I�f��nNE�v�Y�阛���=׉��(�*1/�O�9�d�76V�vQ��v��i�!��u�<$�:�Gt��3�5��c-SK�`�'�
F<�������{���������S���J���>��3��w9򔭻�wY<7
:���r_L᭤����tn;�ey��,�>��߯��_ ���)J�P�9X:�̑�AӔ� P�s��u⎸��F@��%[�8;Knd�μ���^�G}_}��S���}�X�S.�K�{�)�}��ʘ��f@שt��??��m��J{m�w{Wp�wa�D<%�vu7;v�+suV��>���{���g�Py��2�sƤ���������l 3i�ۻ"��2K�S�}��<ֽ�v있�>@�E��TX�Ym@E[IX
�J�dQ���[Q�+(UJ���#���Q[eP ��K�9��3��Ƌ��%��4Z���3��f�:Uz�!ߤ��S����:�mj�3��w?V�;�E�����W��=���d�'5�I� �6.�wO�j���v�ġ����]�1��Va2�Z�ʼv!�t����=�ߞb��̬������y�K���]���9�������Ȃ��ۺ^b�Y*ث>���se����&�я�|�
�ܙ|�4��~���۵��h<�!��h���X���������u�4k;�=���N�d,J5�����r�����.A��{fp��r���x�a�\�s򽠩�,�cT�ӭ��kmf�
�����zml��Pq. ���4an����z@���H��^wk����ɝ���f�:J+J [�vY��eMM��T�*��.�TE옞s(�$0�n{�gDuX�>yXQ����|=��3{�f��YΑc:RT�Yg]���z��F\Q1��Ggqf�'�$�1����5�SDX��m�lB��=1U3Q�ǚ���M�Xc7��$�y\����M��������y�G}�ݥ}����<��8KFp����`�n����<����<m�*�m�p�I]0��Ui����2w~Xfv����^�'ZD��D �d �xSM%����� [t��'C
�����C����  $L�R=ܹm��6�A����N��}�}��8���{�-1�w�Y��fS�l�㨏Q@L���I^?_Y�J�B��|���t2ԁ���W�����q�<!a;�X�F��ʛ�Ysc]�b^��z�V���/O�����ԉ�[Il�7͢2��{�'p�&.}�ƒ�
,@X�J�P��PY H���VAc`�@��
�������R�<V�X��R�Y 7�"�|�Q��7Z�I|q����
=\\��G�:AS2;��A^��݉48�K��q��գ��=(JK��*o�����:��tB��g�]2�<lg�Bj�O�l�rs�����ꪚ��ȓ�ǻ��Uw?�_+ok��"�p�&�_Q�
N�eV=���ċg�~���V|�V��-�٠E����
قSܙ�S�V�b����l���y���|�B�vA]@+��(���~��6K����ym�ҥĬ�\�Lr�'��ڄ�`��zw����r�Lȗ٩cIء���:�4��g��6�S�!7��*VH{��~�o���T''��O�o��Ms��L�p<sA�l��B���fj,�<}[�Z�I�2�MGa���uduq �Q�3�1��߃��Bk�LP�<"�߻��u���ȇ��*���p�Zg�r���:P�3������� Aq-ML�`a�]FjRv�빺�2�9m��y��򝑫����������L�R���m=�h^�}U�{z�ŵ�����;=��uѫ��wP�X�Ө T�� ��*   �1��>}�~l��a���j��۠���2��uεB�k��PS|��ɱo���16gK��t�zEU;����_�0�_ߺ���^(f��.���nT?��q�M����;����ʇ�=B���k#��c&eY�m��P��N�sב��

EC�9RF�೦�ߑ<���;nʳC=�Ooobh9��o��R�sS��u��0�*�	�w�	u�j��W|܃֪p�f�b�$T �H�>j6^�E�u�u�O�gù���֩bއw�T��tWIn�r�ƇVT��fGF�o�:௉�r�6�f�t(�N䍣�.�����#у�=.�W5W��Z�=p����!8�C�$�6�I�H�����p�m_��.>[=/��l�r�V��hE���f�����˚�(�����Y�c�d�3Z|}Z~���&�����Z���3�L�f��� khF�tfa��e�2yn��� X}2��]����,� �4.+N��-2����8;�~�Fg8��H4Z:r0�f��m���U�m�1�\>Y��2�F�xc��{�˿+}��V7m��q	����Y��+��3 Nzk�h�����K�nHL،ѡ�T���F�d�����]d�������'�A�'Jf�,���'i5u���d�'�?3��e6��3������*t1	��������Y0���jFi���ǳN�Y�0��ƈh��vI�'�l$Sm$�4V�Af��~^P
�քn$���ذw:�����WG��&��/2���X�x&�?X�����N�F�f�F��،-n�=0q�֩�E={v��9p��(�x�k��\�E��&:��S@cM���KW�Ʌ��O
y�1-�ݳ$#���(��-�^B��{Gн���Z�ݺ�{��,q��c��d�5?z+���"�}�z�E9I��c���%�v���i���6dL�@���}��7Y�� AA�i�Mb>�d�*�`oN�h\�yi5k�vP�<$��z�T�j��a�/T�L��B�X���h�ݑCD�B) p�r��7��X�n���[��i&��F����x���M�Y�⪶Z�k}?���~{�sɎRg��*� l"����'�����k�uU�҆��X6H��N��:�.`f�>�ݶG��9pY��[2��)xRnO��ZV�P^N�&H����w��������'-�~N�\����h�W�7j�nR1�J��Z��i�	,l�|aM�4�٣t��l��ٍ��H�1�)vJ��8�*��p$�T�ČNp��kZs&����0�z�WT'3�$�a8Z<��80�H(��TY�,:� ���VP���~˦�Q�9�k��� �r���`k.�-��w�ktq{я{	P��try�N��hW���z��<��5�^TĚ�9�}�8-_^k��^:ޏz��Z��d7
n�k��)1�h�����_,r'n�����j�fhV�]©��^I�������ߣ����vm��V�pL��ȁ�ι��kyCk������Bc1͆���L�F�<��, a{諭�^w�M�}��33}sW�E@�+�� ZumJ���_��Ջ��o��K�
�!��,�}[l6rw|;D��R�6K�7"wv���S	�P�EHHפ>7�l|�ևX���:�"F@�IM_���A���oB��p֏W ��^��<����d��DXE������>j�Ͼ��K�:f���P��~A*��@�����83�l��I��w�7;�����9��Q�H�2�r�ꯇ�� s��<�<�xc�;�w�Y�t;�عb&m��Ner����<���ˇ�7&��� �]��n��U]s7������Z�-�J�SϥGyf�m�]GlR�6�@ x  ��   ��v�z{:{Ͷ�8�i4� ��8[l$V6�KKX�%&��h���^^��<kϵ�7�>��ۃ$�������O�@���ȉy���X��$e�""#��EP�4���*�d\�@*����������hSuHE#ћ7�o���,J�d,���t��Xq�h���*;�%���0�}����\�S�)F���M�o���Pan͌
Ne�B:b@P4,!�FEL�KEy-����ڴ��k��3s����%���$fOvK�8�ov�2�y6(!|F�H7s�sۧ�!T뻪��ƛ���	U�!Z�qͧ�M�(:��L�<cc�#���AWSBk)4�¦�EU�[wn[�� �U������w�MB�p�%�B�'N�˗���Ln%_{ޏB�U�V�ޚ��NEþt��n�gx�l�DAd�e�㇮|}��,����Tu�Ξ�Җ���{k*吲f%7]�M=N��0_����~����?b������b�w9�$gd�:-��T3�<<+EA���w���X��p?/Y���ВdGQ���O'd�0�5H=u;�W�;�Z_wq�/\����2����Y��Vo m�k��}��I4{��HiY:����������͇њ�GI��2�Z������Y��J�3�mJ%3�-�:�_Hս��=VH���7O"C����w�`OƑ�n��ZM"�m4�oS۲-������|�Y���~`��כ�1Y��.1�;}���L�>�k�ot�G9s���p�h*#f� ��4Plw��s�`�S�գ��R0�s?|�}+����^���9���U��O��"y�,��^4t�M�,N���M�*�Oď�띍���2>ȃ)ًJ�1:L�5x��֭�.9�4���˵��p�B�O�7�`taE�*�*�Y6;p4*�A \��6mo�(�W�M��X��y�Oy���J��(����z��z9�3��k4�EŔ��rb�R|FT�f`ܙ�ͧ[8s��)���������z�������y;w�2SRE�^ y�p�<6p����ъ�pC옎f	���V��?z�D�� �eÇ�L9k�c!<P��Aϫ���Z0�� �3���@�g7 Fo�N�����v;��;#�� gl����+Fnk�t�3�s-#�����	�G�y5���+_����<u֣�z���_i�
H�q�30�c�@L��e߶_A����@��Wp�� ��i�-j�hDfQ�g���E�
�9�7L��n%�˚sF�u�+QE�i��a�9�Y��w&�AkƱ�r醱ݸd�F5��5ۧ[wɻ;��!��r�\#:��4��k���qBS1BN�0_y�5o	`LѯzC-��r����&�Ɨ���k��1���s��)&�U�
"�B���R`ʧV�~�>�f)��7��Z�͍2���{�i>�o6}O�{ucx��ͩ� '�Iƞd�Q�9Ŵ
շoq�Z�vM�\���s��E��|��n��x���J{���*l�+G9�����~��ϫ|�G^وN�}��궎�64��&�e�k�p_{�TUgv�9P����ڌy1�=̋��j�������X}�z��&�Ys�"�I���LS&�^�)P��b�WݜgQ�)�J�r{�/O�<��|s�Is[}��g$9YJg3�N����lo`C�ޞ�A�Gs|�}��qӁ\�bW
�Js��k��9hʐZ�O��u�=��k�w�&��//!�ڻ'�?CǶ���#8]�'v`=|��Us18ə�{RF扼�u%�6ZPH\M_�X�/�Ţ�܀�;y�it�D�gFv��$,�,D���λ��þ6�����% �����R��?nM����-����f��7�����j�1-N���^�:c%K`��W��y�P�Ķaٙ?�_��+W���uh�a��x��F�W1�\5�ff[�:���J��6��<����Z�a��Ir���F{0�Q�7�{��zi)O���j�a�K7��~�V5q�N_߫��oI[+��ՌI�a�OQ���e&�dXf���[t)�����K`Y4�˭���5��JvU�O�zOgN"�ڪ�ꭍ.�<�7���t�f����eQ�!�x��``�9{�,�ɗ��[G5�WN�7�gIAf�8"�P�|�˘8S���D@�{Hθ�[�o喺皆N��6�2j��X�rP�t9����:.�3�bV�k�&=,�s�i�g��*	��2R^L=�Q,��2j�Vy��ؽ�ޝ���w����/�ۓ=���W�u��|)�9�^>�j���Tװ��i��d��`�m���� ccA!~����Qm�.��~��Yl#�"��u�yz�rL'J���#��U��^_�Y���W+ �	�#P12j�K}�^&�������~��e#�F�m��x��ف-��lA�F6�)|��Ndc�v�L��u1;����T$��k��x���F�,x�u]J�c�U�̆$!Փ��	q�X� UT�Bh�r,�)�y�5�H�[���׀}*��c�1�V+z�����F~���o��z�Y�3e�T�d!z�����7*�;Y.�w��^��9�=I���.��u�퉘}SB&���ˎ�����^��_�lA�V���1��QjQV�`,E��1`ąQE'y�����w\���9���w����d+�窰5j[�M{6��~���3=��3��&!m����m���/oh�VP>���P�Qqsۻ`��q���8]�w���d   ;� �    +��׾|�ms}�M�RE��$6�6���i$m$�OL/���,�+��8�	ޫ�.z_XP��Z�ԓ݀�;S�t��f���7�"�����6�B���S}6z��|C�]%C�C���0 Q�����Lӌ�S�z(��9��}�0vE;:*��q��j�����-�&&e�Kt�,OXāpf��Ľ�7�ڔ&�P�� ��vt��R���8�:8�O����w�0do�`X[��i�k�6�'ji�4�(s52v�T��-�2హ�Z�ȶO����Mn�|���
��X�9�&�Iޘ�z��:��=�.$ۮ�:��J�!���ww�����%�o���P�o׉$'o!� �;N�n4yz6��j��J���!�U�(`���B!3����B���f�䙙��+� �ֽ�;){����{x��֒УqKC��nE01�(�/j�*l�W��I�'��[L�hzۨ�DMY4�hv�"Y�0�õ.��؞�m��m�㢢�p"g����*����X�K�2VƦo��Z�3��b����1P4b[�.pv�.��Y Qrv-��eOw,�e�=�k�����4u7�b�o,CcB����&f}�޶>����=DF ���9'5Q]��-�tt�΃��@����mt��R�zs�ќ���ˮ�� E5X�����~��ՑwZ�z��T�SF*�d�n����/��4�!�����qrttJ�^��$�m�H��X��Ѩ�M�:CM���a�q����� �x�/�����\sk��xP�R����"��`�����l� &p7�}�ͯ9�p�,��
�vGt8HE
cJ�@�)ˤ��r���b=����U �
 �(�dI���zgE��u�Z��k����?v(�����=�NWG-�}֓�I���K�q����O��¬LW�V�<-
O��Hi��eF'x�����������5�^���o߭�I""AE`�dQQ��I����{���q���{���j�Q����'o�4��6#�z���L͐4ObC�>y�q�x�{YO]��3�s��W"�п�!v=���I-"�m��e�H��X�m����m}��C�,�3��v�.�MI.T5k����k��9��I}���z=�[��q��'�**����|�����7'����H�9jls/���0r0ø<!ڭ�4��֕8y�W>�Y���f\�����o�PcgIp�	�!OS{+|�N:>�E)d^H(l�w���˔�::�N�{&"�.R_����W�W0����aJ�����
�C�r�������i����7��9�y�̢9��b<Ǎ���(òÝq�\��39Z�藠���;�r w�\�b�h����Aq%��ݸ���f��Ή0�<
3Fu�-����[�{�~��CM"�x` ��I i$߃$H��ߎ�4���+�~���*#y�#>�E�7����N�_y� ��p{z�w���%�v�a^]�f�  ʨY�/w�����P�9��U\���&�s�)6%AzdH�S��b}��]
fj�t
e�����b��{�e���-��J��L���y�4>W�/}�e�f����34�����������gr�� ���td]��<�O�YB� �����|.�fDf�s7tti���A�p���w��1{6��|��:fM"�$��ۆ?.���[�=��w/�ξ|a�,"�֫kg�c0��q˞�I��1vu�ׅ?Q����w�_m��]���}�N�w��y�W�<n�R���(�T�W��Yz���{����sv���]W��[�@*� p U  U  ��%{G]�=�}Cma �Ϫ< ���|o�L�ߛo���������z"�z �z�0��4hrS7WUF�꜍�m�׺�N��u����m׹z����x�=���"���Q�nC�3롇��Jd6~F��y�y�e�M��0�0�X��N��,t���Tș��xF�d��Pk%�s<���2���&�#�$�F�H�)d�!��$a�ʮ������5�4j{�<�hm��(E=���u�G�#Uɳ''�/77�5N����<��^�*�L��S�pq`��d �����޹e�l�N��iV#�P�舏gx�/j�z}�qy���{�i.m�[k�k;�
�
n��n��n���1�f�:|^�|�]Ƨ=҆i�nɧ7�gvl��oS �pg)�P\̡C]=�ᳬ�\א[��j����]�]xhBܝ�y'M}�4�61�tC:�֌��Tt�OxY���˹���ub\�S��O��mԮ��*��7=�z�&ys{�w�q�rm������Oٕ�ƿ?~ì��U�#~�br��m'c6f��ޙC0��c���6@J&�jFhXXjY�Uf-X��3�y~��m�"��|4�P�1��<2�N���N`B9g����2�q�54�N��,W�0=�Wm��Z�*�����p=@ဣ!|Γچ,���_{��M$��i���� �C ��@6�I������l�i��li�eyf�Ru���]�T��<��9C<X�X��>��l��^��*´mʃ�7'"����۱���|���{�����w^c���YdY"��E`����0dX*�*�;��:���s�����T���*��J:�t�K�A�g˾���$��"D�QA���D� U
�>���O4�l���R�;ͻA�Ѵq��gw�J�ެ�(�ͻ7m�M�]�5.&˅r��(���`��2���ҁ��N20uH�����3��a,.�m͢�51��w'�JYLV������{�iҫ�rX�����7�<+`��źًņW׍?6�����(MEK�#�u2�uK�~�4gd�{����D�_	�i��`6�Ir+$��}t����w������uhᢥ�z��O�7l��4�+���{7��-ÝE�ًn.t�c�{�ѳ��>��/:7��x!||�8��1��;��U=�X/UBzoDDE�<�/@�1��b*�e�鳈���2eޜ�\H�=�S1�j��i-�v��!�8v����߂�lc�W�#/݅����k�=��Go�e0=io*?o��<��T]V�<�	����A�DA�U�H�!���A+�E�F�J�X��Q`��ʕ�"<	���&nR�fn����5r��b�u;J���j'u�/q�f:�TM;J)kgGڼ�g�(�e�_x�.W}�đu*o��ɻ..ؙ�&�g(��z�`ֈB��sN�eYS���ó�uOZOyNL�5U3&*h���m�l�߂�& h�HH��\=n,�t0b�k����6�n^w@Z��`��Eq�@lݐ<�7D�0�ɇ�da�{�>�m,u�
u���a2�И�-\ܙ7�-�R�6�:nzv���'"F�*�k2h`|7B�%��o�t��j����~�X��Uт��4h�i^h��`0��V�Bz@=pu��m'b��>�Σ�Ui�A�jbk_��{y���G�S)v7n���]\�y�1���^^�5U(W1�{\�ny���@����+y1�=0q<&K��\6V�{������{~c�rO��&���=�����V�ɅknT�m����@���_�a
5�fbd|kǌ3k�1��&Zb��QL��t�X-�zy��*�Mf���Zy�4݄%A7�L�ff���mա�32����ZjdB�esn�4]F�M�N��5�����
�|.�Y�b	�0A�b�opV�6A8���vGF �N���na!���oI�4�;�0��׸�4"f2�����p ��N}�C���F���'�a�w��@��)�2��eQw�-*q!�N��42aR+$:4��DV�,%s�(�üU"$7c{,�L$�&�
f���m;��\|d�E%��_��7�������ز!w�hG���nvy��+{�
���U򐪥�tZkTkni���YV,U]2�&��4���� 4ѡUU�)[qY�9Em�؀�=��d91�6��n�au���7��S�)�i�.R�}Y|�F��&�n�����,3a�k$�Ь�>���y^��S�����̄�iB�{�8��W�@�m��1mܷ��)���}��G����=
�W��r�橯l�e�Ǆl�<
#^���ri��
�Y�6�I��C>˽V�x�b�F�G��M�+}��¿M�����H�5�	�œ�����9o:���b�I��ת.B�`VpT�')��O(<��c���G��ϱ��sO�[��TH�*��neJ�-N����"�7Ǫ��G�ǆ-�[%3��K�7�U����/-��
�E��>t��9-����]�)�u�p����Z-�-���btZ����r��lJɎ�`���Ԏн�����Wrzlf��������f�|��Y�6���_]�+v9�j� nfe�*<^��V�U����՞����z��֨���p��h�-u���z�Z` < <6����T  �z��@�Y��xc �l�e *  �R징^��x9R.E�T��v���C՝ٙO 'z�좨.����mN *��J�ٶ�{^��n��Ou�����s�����J���_]�Jwd��m�{�Uz����z�kwsv�P    �>T   '��    e�  ' �*�  n    m������ 
��        U           W; ���w~�w������&�)�8��G��U1�}w(�<�[�>[��'v���{��jq˻X3��m�\m꧀;	�
����z6�nHܷ�y��oY�l�Mݰ  �` �b�   Fѵ{��%�(x� v �H��)�m��<(8�?ɧt�o����A/f�M��zć*�,s(��r���cI��m0��K� ��=�G�{�]Y�z$��-e#��0�W�ר��rI��~<��ٓBq�"�L4*��X�f�ZqO�qSg�{G��)0i;�;�ň�Pthr+��P���فY�m&]���"� ���
S��FC�ge��&�5dK ��|�7��HN�'�%�^'��w���Ͼyu����/|���G�V]��[=�[hQ��WK�;��p4v:K��)<w�-l�ڣ��f���U��
^T��Ei4<E�B�Ar[���X�v�l���5A'�彾�l��U����w������0�P�$0��<4>4'�[���j}�Dy�ι�mv=!F�4Vt��\�����6p�A���!ힸ�zQ�a`�0���ZXʔIY�YJ�#aE�*U`�H��EQ��
�(P�>�{�YO�=y*�����+sG��2�͔�4	�h�V�qxV��7�ٖT�����n�g������ް*�*�a��r�;��&�7�F�^�Ds2�0h~���nG����xX)�u69�t��>l0��=1���hd��;�ν1�=���9x�`zV]��u�;����5�7Q!�뺳�l�|��?fY8߼�Y���c@�(���x(UP�t��њ.x5*(�.�*M�S��n#3��A���L�HCr]Jf����UUWP�o�����m�^z�����ݺA]��<c�DJDBu���t�򝸁5�����Q%�`ژ;`A��U�nz����5��8�K+��۔��P���.��y�.]Tcz�'h���Xi}0��J4:q��z�M@�3�u�M�?0�g����US�FY���nîGYdd�!C���t��,ӽ�p��`�ἂ��T�n_�y�Ǯ��94�ӦJ+%����;)3v���Z�q(yV��^�O�P6J*�EX貞;ƚ�Mn��A�:9�1n��fX1���(��'90��D�p�d�v n�ᬦx�������/	��Pc�g�ۿ��:c��"�b
Ak�|��Ľ*���}�|Х�����kv�sۺ��_V�©ȓUR9��dd��2�dGc�C��'mW���ne��&�tH��֬4�����c���]��e�n���f$N��4Њ� (a�B�"x�!H�O3e��.{���d�}�����-���֡1�`�:.�����]_=���0��;�q�0�LWZt��
�ɪ�w>�i�t��Fd��+�jBH���� hUn��s�"�(�$��S���=�ƽo�ҫ-�y!�U�Y�E;e�'��3�1�3L9'I[�����;�t���X��M��z݀��*���d�,eq�c5Ϝ{{wu����kD��X[�Bx��x����Rx2��t�8�������	c,��E�i$m$�!�E��^��H���'�[�b��jfh�pwX�-t�I���$����3���7���P;ϥ)�G'�%�1)9�p�������z����� ��O�A�AϾ�I���w�������Zw�HCLAcٔ�&�W��v��u�D�j�)U�������>t9�Y0;LV�����r?%�{�܉:� ��^%�_7�Fu�
�ti1ĥ�Ynq�9�G[1+gW=���2�;�,Q($I:w^ E��`�w1Ω�*�zXt�@����{̛����36a`41T�8
�4`h���U0�n���~�_�Wk�͵:���qAr����][���߈�����ێ����eu��������R�w���m�V�y�eW��{��;��׶���Gp� �P*��   6�m�l���?w_���+D�o@�
��Y�-��~��+�B�8�:�@�2l8���G�=r �|��E�9����������"�C��UIVu9>8B,노���n	;�2'�ۮT&5��9��j���{�C��h�:�u(M�#yk16��It,CX�<'��1;��x��GF:A�H�B1�i�x�8P
����0��YzwǑR��YW�w׌�
�L*^gkO@�:�rG�$,�T#"�ј	f�S���zlw��`t�'/�ȓk����'�
c���& ���[x3�-��xx]����v���f�R�1^�q�)���P��ę}6��\�5�=�����ܽ|�H��,��k%6�Acm$�>8�H�������֥V�B|��6o�6P�U��a.ԝ�`~�D��[��&3���y-�o���������T��IEX(�V*Ł������;���y�i�o0B�ӵ�P�x0���vn����Û�r�`'���E9!����T��5��#�
�˺w2��q\y=;m�y�O�iS����fA��\L�6 :,K
	i{NY4#�v�KA��j��)3�,;n�qϦD�$��<6MMMU�*�ab����>d��Y�R�����p`a�82��{�HC}�������2)��L̎�C�s$F6!Ȼ��p.Jd���S���2 i#@�f���n�;]z�TZ��h�,����|q5(��Bo7j�;u��H��Oڟa"���@�F�搎�(��w���9�gt�Z��֫��`�L)s�p�(J�(�t!��K��C3������{1�x���d�~�Ղ���h�a�i��3<B۽x�W萌m{UC���"��n��9�4�,�2/'G82  ��qM�
����7`��7�rJ+�uv'��;��\Z�����<�p�w"�g;�1�,�-K���x���]��D����6/�N����*<h���3L��Y��U���d���FqO�ep`щ���t��[I(j�ֿ�ú�Ip��e'��&�Й4��Y��U��G��w !�F��wu��WPE�i*���_9l23m���
��,pL-0=C��D����`C$�PpF�s����e�s�nM�D��B
H�)7�oǉ��N�~����s'�OtWHX:'�]9������J�������^ �8l��iI�̿��|O^y^!�|m�H�N��'�m�/�LƁ�:NM��SQ�΅����Y��$�-H��r�ǅ=��1����������?�wN{gb��'��!�=�&�\�]Όz6 E>RQ DX"#��T ���9�(�L��|��"K�E��쑊�+�����M�c,���Y]�0eCOBaw�i�$��f�h� fe�k2�C^f,܈�>Z.�==���ن��c�n���_�����/'\�}�m�m�R�*��j�����$Ԭ`&�I �I&zabF��N^�w��&����5au��7��|��� {��m)����^_��Y��Yaݷ��T��ᣀZ�_��8�[�8��d"M�s��t�oe]eR��?V��)�����o,/���J,`����t�������Ͷ��ۆ"ʰP��7S뺝���s��v�UT�m	��i.y�սOէ����x)Ê���f1R�xd���+���t�'2������C#H5v�V$Hर�7��j��j���zf�B���ua�a�B�qBAt�1@X"1DEFD��k*2�Ȳ#+bT���5�*��P{䀺�)8�±d�˅������rނ�b��ov.}��ټ�͛k������_���U=�����<�͵Rp*��{��S�{���զ�S��]K��@  �P *�  �m�n����{�K�'���x	���Uw
�Y�C����y�3=P?�UVq=�@��h��7p��t�d�λ�7ٮ�eH�$�U`�'#MgT�:�A9�d���t)����˞��nT�� D���k��b*@3Ƶ6�z�	܍�C�wq��3��L:�lKʱ0;A� -����9ǻ���mv� ���*[��q��mP�"vPB F�,�39��}[oy�s����fr��16�+cr*���P��qY�k�[oGdγ��}��MC��EUI�Tu����)�4��1��ͪuG�*ʄڶ��Ƨ�[���b����������v#32�f��UmĪw
�w��]����FX�3a���o�gq8i2�bD�)Oy: �:3��K$`c19u1&�n�\��Y��֬ȏDF�z!A`V	J��C��_vfg�͡��AHhPs�����ב��}k=K1hU-gv����c7�b��$hLU"�a���pp��te�j�՞�bE��^�3.�������F*Z�F�GL÷5�#�������ns�u��:�>ׯ "iC��Y�G��BlS���kmIr&�ai�O&[�X V��OL�ٳ3�D�ֵ��γ'��Mi�g�ʎ�*�I�rd!�]t�E3(���[I�s" ��5٪R�z��:�EE�νk�Rz:4�z�6�]v����U�Ts��_X��+��S���p6b4�� *+���뺌��m��#�w&��2�:1�&���C	DC������5,q�:�|�y��b�������!���$+:YӠ���U�:�fc�����c� 5:#��|��jͨ�矻�m7���}��DU�3�Dq�J�p1�lKu���6��f�	i[h�(UcƠ��wh,�Q�k3N�f�F*��M�1��%TDQ#�`LL2*�DF��0�u�K+
��ևRE![o3�nhm�b�����;�0�/�4ʊ��ܛ�]�	�f���ZE��	Q���� �!�89QGc�/�Å{bѺ�!z\y�PR���%Ef_�F[����PjsYɔ�S<	����>���V�}0c&��ǀM7KX�oD3�|뢌�Y�S���q��7�w7׬"X��io
�|��N"�U��[�a�ﲌ�(��:�,!g�c�1e7�hyF�̸1\�v,K.���:�xE�+;���tkZ�rY�7��{��Rg#�pQ�%:3Z;��AcU[Lʌ�f�&b2�*TQ�Uq�\7.V�_-f��V̮e�.fh( �c8K���;/���O�y�J'Nb�`��-��ޝW��a4Ƒ��j/Y�t}o�6}���f�V�=��1x��"O�CC�`\����=Zw+q�Ӓ����p�L���F���2nu�lc+�2L�>��r�����\��x\O �ͳ�"��ĹR��ʙ�"�R���:�T��M�!��v�*���,�UQ�@�y<a�$(U-6��+��Sn=����8��A��wp���@�^�*8�q�����F���n���]�M�����P\T�lq�6�IB
zF�pg-��p7�o��@W�8�X������~�]�/�8��õA7y���[*��$�%=�UjC�x ���鞲+p��R"{K�AU���Aދ����p��R��Ǫ���ԩ�}��Ky0�y$��1dZc�oT��֭U4���: ��vn��[���-!W��-��M4���Ϳ\�=�.f�{��ݝN�V;m�n��w��]����V,nꁳΔخ��Xs���*,��V�/dݑ���v� �
�W-��V<W7/]e��u��Kb��d�wM6t�����0�i��d�lvN(6�u���u��NK��]g�����wE�T����i�S�7+����+[���<��8`���s�4M#��oKK��Z6��뢫�ݝ݁���� �&�I i%��Ri��/���|��n}���@��4p"�]*ʍμJ�ج�q2NGU�Q�ꣲf��F���s��#�Tx�nm�
�U�G ����Sc�
{3]/�p�_'R�-o��4j�0;�&��\�a�څic|P�<�`B�t\�s�v�Ae����"2t�yjѥ֐Եqnh^�bY�0�T�O��ؙ� � ��YAk����j�2tB��cޑ�[.�~�4\��㤯����N�*o��qZĳ�_����y)֓=ڒc��;�s�^D�}U�G;�dYM��#Y��ük�[��|���wO-Z�yPxze�GEh���&m��uZtr��W�������ڕI��a�xG  6�i$�I�N�A{D�H�E��s"���ӳT]�`�)�)Uj�@��*�	 ����
��Y�
�˺�$0.r*bu�� ���yջ�U�1xr�{��Rywu�2k1�v#��/��,�V+ͅ�ʵm�M��M���9hxy�)�4Lm�F��zzdxx,��5���
yt��!�tt�&�q=RX�3�}�㺐p޳\|�ǳ�Vl�SC�{ޑz�mqOe3��elG� ����|�B�24��zhw;f��e�0�U�OKu� ��ü�KJ(��ž��R�ȃХ���tƍ��������|��"�F(1��6���2Gs�1��wu�!)�����v��n���RwE���,J,�{���߷�@=�շԧ��:�#l�R�:�׺�t�q;�7Z��R��/]� '  �m� x T m��h������R\�M"V��`�Icm$�)�A	�}�{ʓs�랾��pPT+�����w�W�r��r�kK�J���������6U8D::�r&6(�MՃrE�Ɣ�Ѥ��4�T�lΑ=HE
��\�,2s"�֠���3#��_hڕx@u�oQj1b��)�Q
#&p��m='��$Vϕ�vT�:��7ѳ"7��9���h�{����>W�6��DDE�}���f�j�&�)�2�L_9��!0y,��x�s�������+��^��J�414X� N�d����w�Ol�A�a��Q90�T39t�"_HdJO��5:ؙ�&R{�oy�Wp��:�Y��eĬ,BE�Ɏ�|Sre�L]Dxa���DPDH, ��� h��67��+j�r-�g�.�=w�!>�	��̃��̼�0p�b��B,�7[�R�H�����ي��/�<���[��_KǅM�gh�M�%O@���F�x�y!1��W)k��#(�S�����9�w	�&�09��� [0sr�����ܑ�;ĭI�|��;�R��kp=&_��G�[(��FI8�o���q��O8�kgt��؂�r���0�h���fFa�7��biS�R��61��^k��bfط��q�N��&ߨp���Y$���*v��GYWW�f�x>9��NY����Uw{?~���!4X��a�[i$�I&	+ ���d��}�}�?×�9�^bYiN�	� P���nw�I���a��sZ��iS:d"�d���i��%�gs���<#���94�8�`aR0�s �A��SX��4�?(P.��"�-u����tM١�����k0�\�<`,Y"���$C
?[�=[̎�X��
%�^�����dP]*SɷWk�z��Ԯ�eK��bUɮ�7��_y��	�GL+e�P�6��Ww8�C�U0��]��e8�6�t5�C��󺼑B��V0�7^��{��,!�n�kEl�N^Y<M�`�8�fsH�����o9��"��4��#���pWN��>ϳ���{K�T��i7���4"��U>��y]�����ߛ��ڽ�p��J��^�B���w��^�iB�����3�AQ�`]�6���K���j�n�!�U"5�u��jR£^�+9���<��wN5ɹSy������í�#�މ��E��O�^��"���ޮp]V�ܹ���S�]p�lX�7j� UU� �=])(g2!qa�qSƬ�0��VO\ Qb����ϵ���-��$�[�w�ko'��J�}�dw�F�&Kޭ�sѲwE��ڶ�]�����S�lKQ/��P���]�!G����J�B1����N���� ]��[.V��Qu�=���;�Bw�Ł��&�I �$��8L�����R�Dt�#$�N�pN�i��b�{�_�B�Aj�h�'�H>��M5��wSP9�zg^4�p+��x%�%;�	��L�g��&f�^��z������s3>�1�Fo�6��N�Z���j�S��-�v�F^����+'�q&;����1Z8/�M92q�70��]������nx��*O*�,p�������~�#�,R8�w�j���&fx���>��3����uM-֤Ӎ�_�<v�3�����f��YυUU�,��m��R��4wz��h�5���)�\^�r�TyZI��(�՝�^�v<x^�G��Q�Y=�ntm�"�̩��8�N<{(�����j��u�K1���� � U *�   �KO{�M��>T4�m'� ���0�۪�����Rf��El��Ը31�]8�9E#|X��t	�H��m���5�	�>{t��>F��H�5���|R�����P�0��� I^��RX���ꆔ�Vѹ�DG���i�Z\*9�1`p%�"^B��P�&�F�O%�����i��.l� ^[��]�5z�!Zz�*5E�32��<4JoTOg��~�g�R�􇙘��&��l��pr��ta��[���<c�jTaR�}�b��eӬ�Rkn1�n�Y����ޤ�tL-�m���N�0�g�7<(B��c�H��|�|߻j���m{o6�nB��S3HM݂(ș�E�,&@�Hf��^��Vj��X{o3�Rw��컇I�b�L�L�{���5�1��μ�f��#�I
AQc(��}B��<��|}�=������d��>�s���5<߂[y�R���\O����(�iP�)�]�z{�~�yl�醉LMTO�zHL!�����.PԹ724��&��-�S,o��W�5+�w��@�,*�9�e�O)t�*s)L6C8/��K��Ңj��$F# ��{}M>qXjc�������):�	(ʏ{�cq�s^���M�a�$.|��6���=����j�3�&�?M�G��=EIaR��b�d��tL؍��پs	���\�l����Ъ����ED��M������ �/���ᓺ�"$Z�:J.@�[N	�����n6�VV���ŉ^��.�m��u��N�:��h?D׷����/���u��r͹�.���Ɗ�Z�ŗ��W+M�Pt@mZ&MQ���U�Gg��wF���7���y��{��B=a{�/ý2�����z�z6M�U7�ܽ3+5	p�2���o��j�Qۻ���6X��ELe)cS��L��m����x�	�U}U��56`���XmmQhi�1�0{L.�������;f�뭻�y4��x��,�粂�lXo�l�ݗy�R��t2[+����ָ%������ǅ���߽�ZH�X�,f0�)��`6�O�����?-�=�[4�
�-#��𽹑#���G� }����s-�=���-٥�:s��TH��<�b��������Zp��� �;!2���G��؂q��D��S~x%Ιd���+���c�QXa3��ˋn�7��W�99jc(���ϳ=~W�3^�K���i·X�Aa%��$k�l�5ڥcy[����:B:i�Z�Ǩ3�Bn]�1�0��L�,AE�E`���B�b2d	m�P�iel�J�J$X�*DTQm�PA�|š���y}x���W+7��8�V ��j�;��wC���y#���+GVWf4RзX���܆�l���4�<nfc��5"zg�P�s����h�]ZA��'v���X�0���߿�ϓm��V�n��ި�y���uA��թ�O�E��E7�}�G�W�Y\��0�o ���J���Y�GOL( `����hQ��\ѣ��և�����]Ox�=ɋ����E�c�G�vX0��<O�M��G��l��hB���Ά!3;k/g as�g�4((0'9��<C㳭���z"=)}aX�[�]lu5rIDBpڻK���_���'jc�'�V�B����'�"��y���g�����=S5ŏ�{7��fjj̖-F�`�BOi�N52#E������w旫�B~;ţ�
�y|w�v�>i�@� ?�H �����!��vI$����4� ���!  ��&�BICHHH��!C� $�ן�`I ��P$� ��� ����O�?��$ ����������������A�� ! �$��BI'�d!H����	 @�?���5H ���O����0$� �o�� ;H ��	 @��kI ��a���u�lѨ@���	 @�O��[� I �$ }�����h��ߙH �o��������$� �H �����(+$�k*�آ�����
 �������9��  b٢�@  ��K@@ ,d�  h         (  ��    :%U@�%EU
�T���R�*�AJU%B�                      >�   @[Ǘcyu�Pm��zy>����(=k]���}N�@5���wf����=�(�>��o����H�
��s=Ãg/����;�4���^��zz��}��w��s�n���owG=��1�m����w���k���׺��;u�i6�{m������`� �  �����/����ﾏf�����;j]�׻#�6��r^����zz�+v�`F�m�^��[�������w�A��}y�8��=Ǹ����ݞ�_ {�*�Fo�|�}ת�N=��6��=꓾��_]��}N}���]���{���w�_N�o����w�y���]�w{z�\z�j���V���{g�/�Wm���4���G�    �xW���ܸ}�}vܽ��oofz�{ӗmk�J/[{�z�w�Q��ׯzU�kv��K��u�m�a���lx�;���{��z��N���z��{���x  *��m���׵���ޮ��j��9�ٗ�U�{�}���¼���׎�oc�=w�����x9=��>�`���ϭ^��v��as�]��{�C� �    �׼�����n�q�n۪��םo�.�w}�D����᷻x���gw/{���W�F���ލ�N�5��כ4c���=ۧ��s���}���h���J%E{���׸9>���{��;��zZ���z�>������-}jw^�5v���{΃&��1��t����|��ܙq��}���g#ow��ϸ��Mowq�� �   w���yn޺��=�>����0���^��U�ݽ���mZ�� �]K�L��.���������I�y���)�{�C�u�of>�&��'�O�Қ����8�^�]���x� Q

��>��u�ܮ��{<��E�� v���ϳ��y���Ͼ�w��j��}�u�+��=^�s�� ��^�uMj�!����s�ݳ��ӺK�ܽ����   "��&*T��  44  ���$�R �    4)�2	����4h�� 44*{mUJ�� ɠ   )�Dª��� �i�&�SB�h����=F���zi4yO����`O���__�~��s޴}��4�}}}}���1�ߧ� $ �O��ǝ���B@��� @�)�� P?��/������$ _�_�� B@��B�H@��.�O͒B~�,!	P��d$��+ I���	
��Y$�3  �̄�� ���VBL�9	$` VI	3	2BrV@��̐$�VHT�	!9�$&L�%@@����*$�* � �	* HVC$�!S2@��*$��d�r@�Vs$�($�3		�s%I 
 āa� V�0��C!$
�*2C�B`� g0I$P�!��3 $	P��0�k $��0	2Hd	%d�H2��	
�%`HT s!	̐���$�	�ߺ��1���T�,߿�*��r}�����"
W5�!�k}�ÖN��2���9E��7t�VɎ��\�eKӛ��	�f���ߴ�߾� |��$������;����]Ѫ���T��t��B�?}G�B�jS&;u�b����VVq������B���q9W�k��Y�r�"�|L��)i�`zHzHzH{H)7��~���T�h��n��J�a�Y���v��G�[y?��f��FSW2S۾�\]n��N�
�-Xᭌ�%��7�!R!�!�!�i����-��Y��h�����|OdZ���(�eo@�y�d;3L�J�u���L�?ng��p!C՘l�n�,;Lٓ�G���Tu��B�c��jޓ�=����K뚘�.�-�����'v�RS7J����e�η�IgeE�n�1���,����vm������qL���Qxk���Jٜ{6��u�8b �*c�w�՝:T H�Wb�̛{�M�*�-��O�d��s�Y��.�T�͔P�I6�����+MN�=��vT���wFu;�R�jB��:[vp����
%�2ĩ���r氮���l�=k����z���i��r�
�������(橒︕��*�JL;1��V�0-���	[����
�SV��QØ����Rٷrf�Rf��0����}X;�T՝ٳ�BwM�ͣ�+<�*�3��C�֚�S�J9��,]v�af�o�{G?Ez�Ѹ��1�AI�ͱmY��-R�D���[�0Q������t�zC�����S���H"m=�52F
!2�cZe -Z&��ν�"�� N�=ً- �~�+�`�FҮ�F�츍�}Q�kl	W�r�i��zJ���o���)'0!�!�X d�$9!��������I�zHx�� �>�>�!�H)H)
�������{HzI�}���o���Ϧ�m�լ�2��]�w{b�R��NX[�ޝ��̾�q�د)6������,�EWi�fdPeM)��Z^���q�N��֕G���&n�u[�K�d�iY�Y,nTY���ӱ���#0���G��H�>N�.v�+5-
.�չ������wWXԹl^�7J�BNrXZk6]���m�վ�[�Lx�
?��(nEwn�E��^�l�j^��H�gr�[W�.�5��kNA�R�0��KH����t٫yV��"�1^"h˼9V��[��նs�FC�s����Mr�tr����1�����Li+n@T�u�$��G9T�����ɓ3�E�5�in{i���swC�ۑ�fQ�m�M�BQx������ziӾ���Ù���=�<x��wS1vv����-ҙ�no+�[�x���^-� �9�б���$��7+se�ӭX�k�2�5L��[C�-ؙ8K� �1����.����V=Cs᝽y���ׇW+p��6��:ͱ��-�j�G����;K�4������5�:���.gs-�A�tօ��0f�ܺI�U��˩�^Vy�N�u����N�YӳQ���(Q���̬S�"�3e�9�a�kn�������s���:i���B���y���Kr�n��;W��7�n-[S���^vej�x�ޅ�t�=���/���y�B�}�w��>�����ｏ_h
B�$�+�B��8�:1:Ry�3Q���\G`аQ�]Ԭ�w��ЬOu����{��_~q��������~$�$3!��!� �}���>]|�w����jrd�)>����?m���ĆR���[8��LFexmШl�m;�H��*�ش�T�թ\�9S�#i0]�u䭊�熘׷Y����v����Iӗu/&�gf�֖��vV�n�_W6�:֎���sA��T��A��١G�~�l��~x�b6��0�@a�9���*�N̓`"��#����2]Xɘ��P���N��l<CsQ4�X����JfI�ku*ph[�k���+f`�k���%h�V��-U	����+�e�٪j'&^ҙ/6�u����e4$]K3!��1[�WD2�,��г���X�Ё�VZ�vիُT˔P��*E�P�{u�QH��J"$��M�'�&v�f�?�b��'_A���%h��ս!o-_�H�y�U�tb�m����-���y[�]�!���.㰝�T����Y�{�Y�♤)�R��-�^dY�3�]�.�Tn�0�y0\&�H2���in	�{Yxګ����� ��A��i�R����W��- ~ō��8��e��w{5��k�B�t�VZ��O(T��)N�%.݅x��Wtք,�E������Qi����{390T�5��I��[P�։F�r�#5ĿLu2�lA%�I�:ک�&�%w;0��oU��ۗ����FԸF3��V�\w�[*��l,d���nʋn��\�0\8��n�YxS���u:�s-ND-ItĒ9�i:��a�r��7f���0��Q�TNf��=���RR$*B�2C�>$������}H}HT�ԇ$���ԆHT����BOG��uh���b-�Y��Z��ʴ �Iz*oCu|�9W�Vs�@�pa�D�C�*B�T��S�}`r}@�����!�!�!�!�!�<@�!R$>�������nn�$�YWL�Gd}H) ����C�C�
AH)
����9�U\�µl�R
AHd��I!�
B�2C�!�{�6ұ}��9�5C�AH)P*Cć��$*C�C�C�C�C'�
}@�=!�C�C�<��￾��R �9!R
AHx�$��_�5�Kja��%H) �+
�S T��!YF ��`T��S�H) ���R
AH)��z��T� ���Ң�H(f �2VT������R
��L�k*x̆HzHrC$��R
AH)����������ڒ�9&g[9��C�w�|d8����=��C�R�>�*Cć����R�{NḋԆHx��O
Y[J��iE��1f?
���ER�{SE-���H���"9+}�d���əYG�c*Oi�HoM+��Hx����l'�$=>�2Aj[�)P��PR����R{`_VT5��#9 �<Hd����V)�=��SE}2YiRx�x²Oi�3�>�@������iI!�<d�<D��rN�G3�+�,����aG�D&dI�I
����<H|H{Hd�
C�C$=�=�9!����.�`��R$=�*C$<HT���3�)!�C�~�d�� �=�9> x�
C$9 �2Cć�����B��*C$*C$*C�C��0O�n<J���'���{￞��>G�XC�́�!� ��H{HrC��X�L��k5��Ab�PMg�2)�!Y���:��+'�
�䇉a9��I�l<�Ă��ʀrC�
C&dS�H��!�i�iI�T"!�B�F���䇌��zd��'�E'���=���Q}%��m�g��=��)�-�<HrC���!�!�!R�!����<H|O� �>$=��xߔ��O��
�u��YR�#�����U�Ƥ_PDw��|���*X��HrC$-)���=z��/���*NH|E�>0�Y<Hd3�,d���w���1��^����7J�i<O]8�汌��)�%OW"O�U��b�]eQ�irQ�vK5,tv�r�B�d��R
AK�WYPKNՃ�R�s2d����a�0�ɨ��T��R
�B��T*VR
AI��J�
��]d�b���-�m�=y�Q-*��*�5�m����+������R
AH) �
������ֆ��j��VT(%k-����T��
�ejH) ���Q@R
AI�s�T��'Y�H) ���"�¡YPZ�R
A@�����B���OIY�`ʁKh�%�XTYKXd-���lJ(1�sA�[Xˍ���at�+R�Z0[l[`T��Q�KJE� �����T�ђ�k(���T+
�aR
AjH,+H(�YR
jP� ���%ڡB�UV�=$*C���Y2{H)
�2��=�>��kE}��C,��L��J"�lI��R�j>�!�!���QA�O���f%h�*AHzL���0��P�ω�ߞ��$Tu���0���̒�� d� {Hx��2C�C�r�=�b ao���X�T��~[�i* {Hx����[`��}�d�O���C�L,|�}aQ~����0y�>$��	�!�d�����Mh��+E*y��}R���HC�`d�X�ʋ�'����>�I�C�C�|@��aA�{�!\������n*[KEZ��C��__[�����h�
{vd���E><��C��T9��ڒ��X��Qc����@��P��E��oK̋���7T��*}�E8A�X��|LR1t�)�EOvUB�T5� ���a�=�x��!�!RzHs''Ĭ�"ʅ�J����mY+P*AJ�-��m�*[jT�+P*AK#l�j,+
��T-�P��) ���R
AH)l3[H)Hd�$>���=�<HrC��{o����ߏ�=y����{����Y䇉�
��������XC��aP�Y>��z��5�za�!�!��Ru	�*C�B�=�2B�>$*C����$=$2Cć0��������������!��B���I!�AHx����$�Oh!�!�!�ih�O�����Hx��
C�N�dk���E��H�޸�i�z$�ѹ-Z����0Y�h�$DE`�����f��q�-���%�%�+�0���߯��}���Z`�1�p��Ӏ ' c �� x8�x6 c ��x <p�� ��  @     :r      � �b�`s����ү@�1�p��=�m[7n���z���@-��  b���@�p0  x 8      '    `�      1�           �  Ytq�x xn�1��P�T�    m�5�mq�� �   x      n;�����i��l�         U                �  
���]�M���n�jT   P  `ʠ  ��   ���U  ��� N ��ųmy��� �p��� ':��v�*]Ne�[N��J^�(�u�N�4��]��;yݽ�m�k�j��7;�>w��^S�.X����g�O;׵�ޗ��ۋ�cV�Z��r#�q��ws�p�����#Es��U�=��z��s���[k�c�j�9p��b�cV���纛q���;�]���޷_l���\m�������i�9�z�U��Ӟ��뇵smW��[Y�������wZ-�ӯr�ex�ן9����o.��^�-�^��y����{;xt��;Wz���w���������n����;i��}���=�ܷ����Kj����w����۶�uO�]��/y^��֞۷mu�ݥ��u6��w9�Ý������%�wd�9�ڦ��ˮ��c��{��9W�m�v��޽�\�y�޽)v���]�s���wmwm9��ݰ���z�m���m�����������]��\�۲����˯v[�r��{�g=z�˚�s���Zy��W.K�꛷	u9]M���-M��n�{s����^h��,i�^�m�w��ُl�η�^��;�u�g��*w7+Mץ�g�W=�����^��;���h��v}ے��s�m��������n��v�7v�nw�:�ob���su�n7-M�shޤ�^��[�U�޽,�u5ֻR��ɻ���ۛ�3y8�f�������ףN���y-��<�r=^�	�˩y�Lv5��_.���n�n��Y�ٺ���O3����y5���{b��^����r�v�{����b�ꙷ�^������m��Pٷ�j]/f96�a�ͩ{���>�W��}�{Ϸ�k^���eƳ������q�R���0�ͧ-]�����=���\Wi�<�/uwY��{�ݻ�{��;�u���c����^��y��L�/i�[=�׽����M���5n��4���--�n�ݻۨ��{�]l=�b��=���L�R���q�^�j�8�w�޼�ޖv������=���{g��kާ7�z������6���n+��/Tu֙qlw�޶�^w��Q��^��޷ڽs���ی��m�%泶��W���n:��oe����ީ���w��:�W��s�Kۥ�ϭ���g�^ck۽y�{;/m]�K�pp��;\��p��{��=��ܫ��]/v['eh��sw'b�/w&G�:�]��_v�v�-n��Z���u�Z���o&;[�i�<'v1���/)K��55l�Nֽ�:��x�S�M���2=Emz���)z^]�3�J\�����n���{i���on�[f���:���������n;��;�������ovw����}{foS3��ί)E�nMq��of��u�+۴{L�Ç���{������f7��jϭ�]��{]�Mt�&��qV�j/j�^su����;��z��5�o;η{�����j�N˭ݝ���=��Y^{���V�0�R��w�w�o�f��a��>��ޭ�roj��w{���z9�q�޽Qx�]Թ,�m�S��n�Mx�o<ow����u�y����\֏^�������rw��S�+��G���5�f�k���g�7ow<�g��[׵�+�^v���y�L�m�^��i�s��N�{|>�ok]�}͵��ow[{/��l�Ν�y�o��eY�]���]��ť�r�-�]][D{l��e���v�E�w*ޯm����wk��omG��Ž6����ٱ���ݭ�m�y�M��m����纷]�uϚ{iS.v޻;����纛گm�.�Fos�p�۵�n�u��w���;��n;�7W�-��;q����g����F7[מ�wN�y�g��s2�����_8�o��<η{�ms�2�ڗa(9]��u��v{�w�wM��.���]�ۼ�����h��u����z�mn���=�{!�	�]�/ZQڼ���]�yk��W^ϵ�ji�%�s�v׺�����/[Κ:�gJ����w�v�u��}Zu�{]{:���wot]ݣ���.��r��j����G��۷9�Lm��6��ui��#�{=ڻ����y��:���݋��d���{����J�:��k��u�j�����{y�Sm�[{���;O]�k{�z[��u�廛owv���Ww���^�[��ܶ��]��{��۽�Sk�i�S\kͻ:�W�z�b��f ��m��B� �0�_/��I� 
� �                  �[�*��wy�ҧ����^�u7r��^e[�]�6�����;��n��������l�q ��������z�_��.ws�*�۪笮���μݘ[%QUU��s   �m�� �@    ����  T����ؠ��wGU�nԜ�m�;���    UP QT�  Y~�~��͹���� �    ��  
��*�UP    �P  [ ��IY�l� ��6\l[%J�  P�
�   U6 � X�PU�  
� R�����  U6�    B�@  T  
�  @  �Ql�U[��   �ww   Nd� �qm� U   @�? U   .w=��.`=�aT��+(����^ff�(    *� U  :�;���        �
��ovKY
����  TP  3��;�J�� U
�z�J��Gp3�k�l��1�U�          �����j�P S8��U��U  k�]��d               J��       ?�    0 �            U *��
��
�        *�U    ?��                                                           @         S�Z�[V�]M�רy��e�{��N�\��vۻ�
�6�w�ñn�Ώm݃;���J�zz�j�q�۴�nw=۲��[fۗYU�����Z�T�b�ݵ��su����v���U[j̱����6�X׽�k%@��UomG�un��;��v�Һ�w�ob�[j]:m��l��|�z�m������[;�m���6�`�l�9���  �sJ���{o鶀/��7��/�A综m����csT.d�n6�T�\�U}��U�T�T���ev�n`*T��R�Wԛ�{�f            ~�       @�t@                 `m�z�                   T   ;�     ��         T8ڤ�U     T    Cl 
� *�                 n� ̪�( 
� UT-�     
�)�~�@�            p�hm� JT  6� ��T             @ U P     �J�ؕ*T��Tm���6� �V�ڪ  b�          � PU �*��P*�J�m�   �-�T �ꢨ U   -�             @�Wt�        U              m�^��          R�   �                  P         � m��   *�P             T�t�UU�w����� -�[(      P T�  �     @�           l�  ��  
� 
� Vڅe  +(*Vۢ�   ��         `
�      U-�   �  P �  wb�E�kۛu+b����6�q     6���M�e 
� �fN��w�kݵ��ܫk`�U����           ��7�
��Y[`*�U@           ܷ�� m�Wu��� +r� T����� @w�fۻ� T��  �U   � YVe��UR��=�omR9ު   �EUPGu߯�?�=�B ~�$ ����	ć�� HI���� z���3�����		'���2�/�4G�L~۪��HÖ�m��m��  0��w��^�گn�dr�sn����Ul�Z�v�� EU��lU�
�+���@ � ���  7[+��l�PU�u�5{nh � �+u���ڪ�m�  �0�    PU    � *�T             �;�������n}z6�r�m�&𸹔�Uy��ջ���u�\U�˧���ܳ#u��P  
�P   �   s� �T �   m� [ 6�  n�T   U �^��@   l[6�+*�    ;v     �   �     ��  ��J�� �    fU@UT�@ *� *��n;���إPxT��� m���.` �录P��;��W��q����}�}����HI$X@�P$�X���f��?�����ޫ�sP�f�wm�U)u��*T�Vڀ 
������;���Ѭ�m
��[` M�Tm��R��5P6ީQk��T5X�@tm�n�v]�����n�hE@�	( aHL��c���L��7{;�uG9���v���Ż�SaM|/�,�$(��I�W�tl�$�}�Ir?�{��S�y�Zb$$9P��e8��ً�t��JRJ�iZA��1��GXP�Y_ml^j�E���)�=n��%b�u�e��p�tMu��7^w�]���棕�WZt΍�H.� P/���^kdn��z��0�s��v����Q;���@%X;wX�X�bM$�,��f�*�Էt0�Hm�ѽ୩���s��.A����������5��߻��m_�n��í��ض*-U��m$�sV�j���V�؋c*]���&`Ղf.��N�?+�)ہ��6K��n��~^��@Y
���6�Q���
`X۟�9ηL��m�����~�y�uh��=�wok�gyuͮ��\����\��i��}����F����ooom{�%�g���9�ݖs����h�l�����{��W��K���t���?�91��ٕj���fw`�k��l}(�����#��KA��e7~�`Є�8�io��D�����:ZȻ/���+2t� I�Hkbl�h4�
�򜨗��iBP�PH?2d��e"R�Kl����㹒�F;��!^���'�Kբ�YT&a�֍6�B�n��Ev�{��y�Ă}�׽��2(�� l_)�'^u����� x��N����h1��M�+�6�׷��C�AT�H� �6�B̊�}z������xݹ�� ��_�o}E7��l{�2���	4�#�l@eI��k�7C�(�*�G�{H���^�<�ͮ�se&Z�rA���)�Hu�}5{Ȑ2���X/r�����U�*���C����u|{�P�V�;�>gИ�'��~G���:�`���Ǉm0�I�:��Z_qu2J UN���n�W��n��1_�g��~��=��N9D��<*�Z�k8�b�wR%�'���$�$��%7��ޮ��[���;��Aכ�1f :fE�<�=FJ%z�]稝��"��ĒI������ڪU�+3u���&�%��!1�ٕ7�x��:��]�4kG����.[��'�	��{��I���(k
][ �����wX��,��Ee�[y��-��'g_��'t����H�2���lw���6J%$�-��.��G��]�سՠ
���d�8\�>��4�sa[e�WMcb� bI!^��̴�� �@T�����
��,6�$ I�=��Cw_��\�Q���� ������?Cs�Ě�����5���2_��X�@�݉+�����l�u�P$�Ԉe���q9�+�j�ոwf�3��j���ʓ��L�N�	�����ˑ��ki[`�W�f�c�$�0�)B�QL��M�Vɽ�a�gB��K+Y�y����N{T72r&p�pfa�EM���2�� ��E�f�=+!�Ȯ�a6';=y~���]�r�x 3\ᴐ-��Ү�$��u���߽3t���(@a�s������4�T��:���rԊ,L�^0#,��U=���ˏ)ġ(D�  Xd�h�$m ��-��x�/+[5	��"�.w�����������V�@���z;a�֖��c�,���S=�^��$��G�9�[8�	�n^�0M䨠�#�CpS̮��HCÙ��+�*q��{���=ݫ�\o���M��p� �ڠ
������^��]m�Z�
�   ���[��G�w������;��b��mT2�YJ�� U <6¨�� �+�����m�3��,^�)��w�� �R�m۶Ԯ�l�R�]C��w�}�N@�`��<�0�v{��z�a�C]^�k�9�{'�ţP�J�K�C^��a>B����>��j�c4�b�&2�-s��YI����߄��:cˀ���h��<M����P� �rZ��ҩ�{��Dm���W�L/z��C����Fm���0� "�L�
_8H�d6�i�E�,�V;�(Q�;<m5q�*}��5!�;��W���y+�ɴ^nv��E ��h��7rn�P�wF� �z6V`1�wf1+�y��j!�%[��orR��u~�X�mkN�л({m�T���$�M�e��%��i��؞��Lr]�A�ۖ(�2QX�Ns��>��I��4�fܥ0�[��e��:�i'=�B*=w}2o�o׋n<u��C�a�-�I$�6Am��m���ߟ��lCom���N�F��݌�k�=���톽W���'y=v�ݟ<��޷{z��u���q{���ͼ{����g6]�l��owz�m�%��0IeC�� �Vc0a��,B�x[���[�0z���J�Pn5���KK��dce��%�ALn��Տa�w���h�K3KݠT9q��eq���E7���]�v�^%���l��*���A�a*"��e�d$�"��F!�`Ca��x�\��T�X�wT�Ѧ�?N������L��חyހqb4�cf��8�ᙌ˻�\��L�G�ݞ� �7���W��qm&uܛ���e�c�=�r"�&�jD��T}�eت[%6^[%��ݙ��J�LsH���fM����]eW�yʣ�J�\N�{E�r��	���N��߼N���s9j��>�b|���٣�E����
��2�!�w[���jA6��i4[���\��FΛ(�8���Q�4�N���ٺ��*�wSZ7I9^VJ��E�Xq���� �o�R4ً۵�B֒�m2����u�J���J�
mQ�A ?�H�&m��vA^n�<����~�g;��E^9��3�! �5�le�2�I&ɦ��Q���g�v���=���bR�m�WG���۞���'����f�}��l娀�l�e/Oov�C�T��ۮ�a�h�'=��˳�J������Kq`c���:�����pBm�˺�v�%E�w욍oF����hg���j5F�gQl-��Cȓ9`yce�P%N'�C66�%��F��W�{�嵆r�D��sx��y��Ҳ�����ۢ�J�i"��C�K�7A;���]�u���i{m�ֺ�d�b����h�A�ݲ|��=�N�-u)N���QQ��lQ�rV�,C�>�`ol�3-"��[���闲�%��������}���_W�_S�|cWh�0ru=��|�{��"K�黫O]�5 e$H,4�)�������M�b�X�F�I�;o��M_p0
F�0n����wgf��VDc�h>�S�(�e"a8LH�'�����F	cB��,H<�"V��`=�vh�g RD�<�p�I�A��c������|��8(o��6�dfVI�+{��	�Ӭ^�i �?f[��"m[I$·f�H�����b��L�u�Q5����BH�Y�ޯ�����ROK����޲s6�%I6�
xN ��I��E/�������&�v7f��r�Ј�No�w�-�����2����w^yV'l��v`���{ږ�CE��绺����^� m���_�*�@0^�ژP   ��*�ۗ|����AT6�UWp T�U*�TU x�  U��s.f�-�Q�r���նn�Ԫp�m��m�Ih"�)"T��;:۱�r�����a�b_��()��]���#�/L�B �ම{$�H�J�,*g�ݍ�H��i�jfP�<"��3��� ���!�oD��N+�yxS�&�Q6�e�*�ۡ�窞X�4|��;�͓B�S����ES{��oN�Sm�����d&�H�B��&A �DA?�!��pL���
�cD�m�̿�1z�Z| �70�[<(r��$KmOzݠH���	�fR�^h��{ݬ߼{�"u�����Y�cЊ;�ClV$��`�* �d����l�UU� J�E&@(�Ӡ�ޭ�^Y�r�؏8�:6�/ft���{����BD�[���c3��d��S��Zk�aS+���E��5������B�-5�y����U��t� ۻ�� ��zj�ϻ7���ڙ�m4q�������Þ�f��#׸��li�u�aݜ�uk��ǐ]��שw"����[��������F��v���(""���W�^�$���}�g����ޅ"�K�{�jF�P	��\��y'ޛ�w>�P�x�N�>��yd�U�nlɋ07��Ԁ��vR Yf��A�I8v�=�@�L��ASD�m�t�*��N���Us�X�9�e:ѱTn������M�����İđ&�%J;9m��bqV4�%�$Iw!�
�9�{�u{�X�ݼj���,�H�ui�m�^��U�Y��H��I"�>{uY���Dfޔ�{��S���g�z=��W����Y��ad���h�Ut��B�m]`�݊Gݻ&��kJ�G��z�RU��ۗ��j �i$�w��z���|����<���j(Ȩ��TYr0��<
Q�,�^��~��H���{�)+����/,^Ʃ���SMSB��{�I,R�Q���z�.��g�<([�
cZ��O��2^�t9Ǚ����]�ZFP/7n��r��=��S��Q���u�I��]��xe�
�������wOGV�abu���7��2b��[�Dͫ�*.��l_V�/�/VM�͟A�LD�0n���nbE�v�Vh v�y�kq|��������>��/S�Z)E׌��9�S��U'�)}R�t&�4�%a'������|��C��r�9�!̒jza� �׬x�����x��{`�P���[���2\�C�����3!	H��@�� �$������ ���OL�|a$2@��{߃>���H�	�0�$� >!hC�2B�9}HI�����������z�����  '�� � ���c������G c      �w`� �n�'  \�=�     �^� �c *��=��]����M���]Å�j7���]��ᾷz�ל�v����{�v�g���n���k�n��9��A�8ʯ5�c��{��N�0��:��v�������3���}R�ݟon��lu��v�yֲ���ݣz����^p7^��m��ot�ܞ�}��w�����ܖ�Q�׃u�J�[[�.M�p��������7�7����/ok���<�n��͸�w�����i{[M��x�w^��g��Ǹ��o�e��滜z�f���d]ӵ����jQۊ�^�ڽ��r�����//���h�ټ9랻��sr�Iw��k��WW۽��ƻoW�gy�zۙ����z��km��>���N�/og���ܧ{��|��w����C�o|��c�L�׺gsvtu�*[��ӗV��{���O'w���<��t��i�W��0l!������&��q��Q�u��3Z-��0|�*P�
���9�Q�n�e{�o�붢6�p3��w.��cޏ���5[7+�ׇǽ��ΚXx�r�8���m�Q�f�>�dѰ�Ȅ6�M�[E�� �
bt`�iF=B��.V�b����U���E\������f����K���"�`ٴg������f�e 
�Km�A4U ��U�sc��eFa���KZ]L����!Ҕb�cC_{E`�U��]գ��m�d�ۆ�M\u�%n��{&
GT�E���~�.M�c�����P�~�J}f0M��h`ō��q�Ǜ��i��ĔټU+�/Ρ&8�,�đuK�Ov���1��TP�T��	��<��q�ĭ��~?N�)�Q��Ie?r����b��AF�"�#�j7�W����U~ow�ٶ���y1Ӝ�m<$�n��C�uZ�M#�5���$^-cY�.>9ZS��Ytq�S����&��?ۏ���'yj�yے���gˇ�n�I݌���LET%j[-$�O�
gt�-�*���x�������7GP[|�
��S���]t4r�a��\���yH\�����p�t�`:i �l��)�EwP +ս�l��������c[�~��xXF�r<����Vi�vl�ַ�)�pM�D�K�d wh�@�>�=��A	$��å�J��U�K�K�Y�7�<
w����xH�÷;�Hөu�ّ�`W!��D�]B���?M9c �a�w��1Ct�+I�nJ�~�ys ��/`8׫�\�U�r`���%ϻ�$
��Q���T�H��q1�hR�͘����՛}ӟow����^n��X�=�1�����&Q��c�I.��	"��o#�D�Ţ/�v�6��	^���1��m�W;hPM�J�~����Ji>68@'m����~�m�ʫa{��sk�8LhSA}����ۼ��`��#�|)�oت��KY3�oN�0�l��խ��N���#.��=�m�M�L�~�m=�u �[��������iT��T   ��6�}��z�i���lw  � \�
��U*��Y*S� Uz� �g����wu~��k�uEU[6H2�m�E0�e��#��&�p!2�Xm�RDBd8#~�]c�y��3��x��X=ҏ�Mx��<`�<&��Œ�D������r�1�b�;NI02ͤ硫Z�}F:庣�b�/J�m�����j$�6��:�<KӉ,(9$�E<���Ev˄����܁�S����T�ƔՋ�CMw��Ա�=�J}HA�,RSp��|���ӡ]�#+ձejZ� �� �0J�[i /������_߼ƈ
lU��
�O$0��8պ藹���{��Sh1$�yU*��m$�LW�СM��~���g(Ά�!�(���&�]�k[]R�#��y����� a���^��9���պ��q��� jM"�m�_̈́a��i���'q�=�!d�P	2���`J�V.e.�D�g�1���$�W�M����v��{<�i2ZI����k���W?1b8v��-��o�7�o�{�+�WX�U�؊�Yf�ۂ�C��=�~���ݞv�ݽ �y����Q��M��wIyN;S������.���9�^�ҷc�Vy{�w�j�w��ʦ�y��}�߻��7{��S�{u���Κs������N	D ێ�����~R>�4V	`���+I7�ܯ:�[�t��:�f$�:�M��1W�YbζzJ�7�� 0xmu��G�<(�ɦ�m�]`�s1�t�x��^�(�wqW�	�s	��$C(1���j_LM�P�J3;�y�%�5��q�ջ�ߍ,�N��+t��w�^�iC`����9�-ؘgI�W^1��!nN�#Y�B��E��0�� �j����S�B��+A��©�]gD[�:�A��Z�����u[�W4�I�V��[i$B) m�����;�
���w�÷j��Yޚ�8Kaj;FɌU�Z�61P��ѿyu�%��Or|!�Y�{Urd$f�Gq�����6Ia���K�Լ�0��E޽j����<�d���:"�1�3��bh�×�	��,�)� ��tɻ8ID�H7y�E�\ ��O�1�Ye9ͭ�w\,q�o����8|�+s���ĩ�e"a�2q��_w��Rq,웰xP��H��8���PQ%����Z	��x�L=�:a�hG��� Ime��AJP��Å0#�W�6Z�Fb�Y�o]��'�� ����Ln�ժ��B���n��xi�~��F6T{��l�π��2�'��ܕ��H���|i��C�]��t�\4B#_!K=+�A"�ʜd#�H�vãXD�J`k6���qEn��n�J�&�	Y!��1%�m0ܳ�����h���g����nHγ�Y�1c�Z���bϖ��9>�zͣ[�n\�$�D�6�T�j����E��t�
b���8;;0�%Ը��ˋ��ԋejM2��X"�iMX>ZE$�@�n� ��,(1��P��P����g��&��;*��Be�P�hOut��u��i�E���v�E��Buxr`�9\���@�B��%�0D�	6�pa�3]z�(7� Ѥ��q�4A�9zۦy�4{���	�_=p�2�1�m��^J�̹�2��G�6�����w)�i$S�ҽV�uҋ+���J�������V�"�2A�\L�ى�+��^��sp��b��d�l	E"�$��)��m�ͱlTs��g[�nӿ�����>�^a. u�5Hw])��˺zy,���=������B� �x�ň��J��%"�p�A����[&<8D��.q�,>.�Z���';\xč���I��H��t��'���:J)Άz�ے.�R�R��KbE��H�P5 �2Zs��>(m�݂d�?d��)���/ĝ�Q������{�hݸEb�i X�=���۝�R�$��0�"��?#
	(��f�k["n��WF4{1vomL�s��wͭӈa5;Lxq7>L��!���3�	�ݘJ�%�fI'Y%(�D��vk�<��I�'�N�P�
�iBf��x�u@#��>q1j��rp7�Mp��Tc��t!oL�U-���RTaI���;WqN]��J�A������:�ۻ���;�2}�� S:�w��꺶�m*�*�   =s�wn�7�z���wT6�*@qSm�� U <
�P� ���[��v=���Ϳ~l�o+�U����ٿC� ���{{�X2��������e~���L�MC_NݯY��1��-cG0P)�FqR�(�4�v�m4�p[�%b�d[|�-���vbb2�K["m�]fD`�<z0��`�Pj�p$����P�'�M�f����N 6,��e'5|�i�����L`����lMa�E���gT?ZP�;]ؼ=ܠ�׽d vG�/YF�"�bI ���}��W�:X�{��ײ��Kx��'f�V��^�(H��,�P��Yn�9����q���bƶf�������=���]��qZ`3�k@4I"JyǄP�������
��ڍl��xF������J�7�ƌ�	s{�)m�b�,�w�T$ �m$�"�)��B�r������ۻk۞�Q�GQ�GRޞ�sK��o$��{��zO ��� ��w����Ck�d�q��S��wO諴m�A[m ���AB��q1IN���K{�%�XlecSB٩ض�ٹ�,�H�x(��,�I$��;�1�w�{`<��o������{���t�ͮ���]��#Ayj�����x�'J���k[��(�R�b׬oqK������^�R���[�� �P�%� ��`���$��%#���E0W���$T�Y��z��'�G�2� l�~��עV{[A���Y�S3�|b5c��ƋJ�v�a5�)U�8��<7�~:��]#��B�mj0EY�p���%KD�����T�wߗm��t����u�-���ۄ�	���"��t@��k}F�{���P��]c���3�}��覒�m�rs$��0��)$�.%������%�l��y�!G�R$Б��ۡR1��);.s[[!^{��D��`�	����h�i6�m�]� تU��`�l$���l���0�~d�	lDU��IU�Eq��طћ��1W��R�Ui��x�%��!1N�� `������.�U�૧Q����R��[�⼙X�W>��C~g�kkx����V+j5��;	��I�P��Od���D�!�<MzW��T	h�?y{�z���ߪbS�K:�HZ�k�V�SoW��Z���PT����o/0�����MD�s>Ɨ�ZL��A&*�go�-H�^�o�j��=^��v�o7O���	n�	�W���{P�dX&�'��[��(�73�ޤK]�NB�w�N��-뛘�d���m���0G.^�}B�j�#E�x0���:�*��2�Q���;��{�x����Y�>�Q�fg*6����R ��m��d0�@� ]���v�K�!�(�B���|VȪ�(p����$�M�l]_y�0D_��C� ƕ���l$K�T�h���
��ZB,��PUC�9N[�S<�b,���)�{G0�Q����8*�2������!8�����Rxb'��	��YHQ+�ݒߜb�Y�b���{/(Q�*��ㇸ�,&:vM�i�5��xXQ�����A�&�7	�[)��>�ox��.�GN�!&l Q��P�.!�IL���K� ^C�l�Fi	1���o�湊�Ra�¤���i��G��{�觘�-'�1ة�����g�)������z�G�,I����$�46����x�H���$�z ���&��g[]!l����<�^E�u/��|c�A�΁�"ߤf�����:��F��7�EV��
���I�[h�-_���XQ�Ҕ���A6v��ƶSe���=/dOS�ջ�CD_�^�0�f�H$��'�n����m�����k]\�M��s�$]e[��9/=[-���#�$N��6�H�a�b�i1H��f�n�j	�-T\/XqL=9U�M52Cup{RB���T۩��j��`!�/[*�}e:�}B�0p]�˒4�8���%n��K5�u�މ*'$<�~�ݥ�)3�Jv�y�kZ���v�r�׏wD8�+�,'� D��\N�C����K��*.W�֗r3�@�OP#���
�5�ǪʢRH�\3�+�vaAA��&���F���S|I�~"�2�5�8������Fؕ]�8��504X��j>�S������^Z醅�wz�uh�n��{�vltvLu��VjɰX�Xxzl�����Iئ-��7L�z���Q+D��#�/ٽZ8� �T����+/�$4.�$L��xDUm������֑���ۛՁ�f�:^rf���o�ʘ�:��W%�.��M�\,�\��>��Q����DΫҨH1���j�CA���A��qٱ
�{�s�Y[�*������Ә/ܒ��T�#��h�����9��^����}���]|�v����zO,����U\*2�8��_v�ya�$S��$^I/��3ӽH~5� ��$�?�I�'0���I�X x�$�2J�!�s!9'�B�2����x��H+����k蟆y�{��q�y��<V��m��m��m��`U��s[��kMT�7��T��ݯ x f�U����*�+w;�M�T� �m�Z  
���TAl�  �!�Ux*�UU�TlwQ�� �T 5Iz��U V9:�  ��р  
�                     @�θQ6���X�u��v�=Ի���r�������vw�/l��\�v����]c�\;���y�   8   �    ��  ��
�U    U
�� @  ����l   @�#�UQT ��l��Vڀ   v� @ ]@ *��   � ��  p�]� w�   3 � )�    U
��繷�����~���� �UE�  ��Ӈ�����G�w���q	Ž�w���K�}<��]�m����� *�9�n���~ض�TV6T   �on���_V��=���*�� *�p�֡� 
�W�   � 6%}Cv��s���2�����}��@�1P�Ϙ�	i�.�2s�
�PL�?#t���uh��xC�=-^B�D�ݺ�D��>������c�J�����oT�$ӕ-��I�߈�C�@�W#�q뾗fߢ��[
�'L`��oLg�ob{O#�$ ��=���\vB$�L$�׽7�p�_vI�D^w+���"A�=�M9Q�N������z�r��1W�c��lDVw:���d�"!1::�P�Q�>캔V�}�[���Gp��h2QU�Gw���NIH��M�\<�(4�o|�A�dƤ���(n]�EE�����̀S�R7����5��m&PTj8P��[]3�j��"-�gzǇ��X2a{GBo�(h��{2�oFrBK#p�::U�7���R����wP�]�J����6�H��Qi��H�o4��z�;3>��6,F��z�	�L��U��p�@�*w�n[��l��4��ݲDq^}׷@��$�x���g+yA�����sf\�>��1�e�ե�9�m9g,�ճt-�կu�h��{�=m �۽�� U �u��k^�o=�������^wM�7
�m՝�{�s{�l��{�u����v��[ܲ��qlר�dRݎ���i�~�M�@B,�*h��� K0�m�����U���%ޗ	A�hG3�1�\Tk �aq�w:�Gm�C{�!���_bx[��m�q�J�=Q����K��.쉍:�a�U�#A8M�HϴWs�
R,7�2c��~:�Z_2�d�S�f��I�� Zl JD���0�O�(l���FkwD��	 �kK��2)�&���(�υ�'3��WBI�ޘ�	n�1�pX6j�ɢXM�Su�HI�:#J�����'bˌ�ybo�O�^*��^�PL^I��-�(��7d���]�oo�u_���{{Mڊ��J�w37m��U������w�1��{��$�����H���}y�&����ͺݞ&�_H���l{�l�V�P�E�C�3��,m�[�-PG�`6ɴ�k���|fqb�َl�>�k�s@��4�Y��\�Tq&f%�[OU��s[�v��(�@b�m�=�����jJ�τn'�͔�fG�f��v�������]ē��`�p=t|"�V��:�Ȫ�[�<R����ʽ�0q|/O�{��j�sT��l�X��(����t$�D4@�� ��5�6f�d�WK������@]s��ErOy���D�����5~G9����?s���b�d��Jt��E	�;�C��޽.�xP��:->�te*gd�ҿs�0�MT��Vk���8.�^�5�zpB#dN^��S��$�A6�%6ʀ�a qllU�x�r�m��Zb�TѬ�AC����6[z���L�A��3��3�-��Ѩzcp�nĞA����d���,�b.�vȪi4�)�\�$���C����<���h_5�Q�H�\d� n�^��4{��-���E�{��!v�<6׻�&2͖��a'NkX��H������}��-��J�k��v�@I�:�4;d疹�K���
Q�<�4լ�i �I0�8�+����ڇ�$��I�@6X�2�1��L���5{L8\؝�o�tF��F��K�;6�������Eʮ	�:�)�a�ܬ
�vs[���V�H칧w�[�����GIܳ=|�M��h���Z%���ĳ���>I�m�$��b�o�{e�z	�]��=�;�����"<4A��{{�2�vg�wZ�q�f�f�I%I&逩��l�� UU���%�I���V��O\Ե��Xn��:I���4�8Xt�|0�14#��
>�t�)��%�����֟]UL0���J�� �s]"wNK�Zݍ%�0Q�5Dwx�F(����KV�9f�	��I�92,Gd�v�;>�(ģOŋ�sd��x-b�X��}=��ԡ3կyV�[�cW�0��|�Z����.̛�cÄ�'JCKi L��@��ݵ��� u��=�s�,��=�����il��#۶�67���a�0+�ǁ�4�o��`�W���TN�f/��$�0��m5uj�y-2�y����!F��oi�.�O`8�yM�Ώ�E��T{�$^=�"@��$pBÓb0y����5��$�^�J����*V�����Q��NU��	��Æ�^��R�
�ml�Vz����owo߶ͱUT   �Wf���,��޽���U�m� m�@�  �T� ;�@��	��m��b��z���;{��*�t�W��р�("K`��0���DaT�K���k���y���$>'����k�l�����}]p��&����L�	���n��/�������G���J=��sY!��k}��;�^n�hn%��h���ߦo����h�QDCJ|6�H��b��$�1J��*Ω�����ʃ����@��G����t-�� �w�PJ��&ٯ��iI-6�C�8XҴ�X^%�(,�P�%D&���6D��[Q���j����V����.lňF��G���\�;��L:�>g��2.M+��טsM���F,�Cq9�.�˹b�od�6�N�v�b�&_�čbR29��:`	#$Wn�9��O!v�	��L�+R�ݟ����ZM�B)�pw�Ҫ��UW��[=r!��D��Ј��t'3��h�w��gu!��mn|���,`�����A	�%M�`���*	I"ᚈ{t�>��r&� V��l�R:G}s����������9��~�?��v���۷�� v���z���[�y�s��uf�6Ƕ�7v{w�W/3��7v�ѓ�y������7wo>vl���tiލ�w����۽e�zX]���u���z�o:��.|
��r��~K��'T�zuJ֦B�C,�'g�#�L��#�����s1��aOK ��&�Ю��'Dp�&-,���j�V�������F�þ��M����65E,���!բm��RH$�J�K�E�wM���I �0�]�"d��4x�7^-�g�7�/	X4����5;�H�ìӔ�����ҧ�w�,�K�nb���	���P}��	⍠�b�a�?��~��ɨ����'o�:���FW���֦�R�:6Lk~gX��`t�d�'xϯ.��͒��L6�I �l�iC��
�����m�D&SC(wj��B�,�p����8�_r�O�wT-M��S���9�3`��q�ڞ��Y	�ȕ����D�n0��&U���5=������5�0�p��4Ӄ�o,G;�".�=-}}���Ck�r�Cgot���\൲Z�%�k�o(ູ�NL�1]��CT�����>;.�a76�B�\>w�L�GҦ��JnO��vl����%�ɯ%o� M[�����d�a�W���V&|��JI1�ZlF�����3w��޼l]�������wOms,�����!�Nm�Î�J0+]�8��:��$	�Ò�i1�WQ����N�{�m�рlB-��#���/�_W�%��QׯMu���,��Ţ;&�<f��k��ԑE�f"�k3�nlu1-/�L�Kl��n��6�m�J�n��M0�I��E4��c�5�PZ&`�z��1T�f�;f{�n��V�p��PQ1�|�-������c�p�e:��1L��j�����:�#4�Ѭ�{f����;N�l�$-(�+����J��M�����P3��B2���1$�p�߹X���eGs���Ι�8�^a�]�c�**�������v-v���E��ٜ&D��v<�L8N��O/�列d���(,�D�[ "h�A$�ATJ`"��*��_�����5��ji����-j�]Ƚ�;������k5���
��UM����9���ӵ��0����$w��;��L��j�0;�D
<��pf�ɼ�Tu�W#׶�W.k$U�v�g����N&]{�f���;���u[�U���M�[l�(|�i��M�-�����s+�
�������;��Q������j����ؽ:�7~���d�Vsj	ΓZ���4��{�Cpަk� YF,�����x�b�wDYZ'dZ����OGB���8��u�1�:\[K`K?[��t�N�a���%��E�ƅ�p�-��f5��[���(p:b���[�UI����Ƶ�ep�(W%u��1=٣�(���W��n-$�IRg��J��1>�ܵ�)(�Qg�Z+v��'n)�Q�f#�`�`i���d�K��~�Q��E�w$'5�����!�B}�`��W�6LH����#�\0��<l6(ʵ��W�gDx͌Q�9~�I�Q�^i�7 �Py���q�R��t���U�[�G���E!�?�6��5�p�8�\���\ڻx/��'1��A$��`(b�0m���m����ۖ��eP   �t��\��zn#��m�T6� T ;�UWp U <���@
�j����On��K�m�Cs�;��d� 	$I�-8�J	����~�N��.�É+xO��8���H8kڵR�}�V6s�:0������0,��I&��~?`:��Z[�lǚ{�㕌ٝs��%���pX��K��$@s�6�q�u��\�o*�8��_��KsvÆ�6�h����z͎�B'��{��Wم��.Yv[�Lӫh����>�Q?d�������m�"b�]�DD�H9�8+�,�w\�u���w���n��x���R޿��]����v�@oM�4!�L�s|PZ�xp1�y�MeM�S ��覐Mkq0Q1b	�L�W���G�_'�FN��ubT�s�OsXFu�$�־�I��� �,�p����l�������{k�����6
��EUz�U*���v���wn�<#�y�������1�m+ݘit��T}�܁&ƴ�o� tЉ+v���%�gC҅�j͒Sm������Ҽ���� E���;�w.wb�.i�Y��[]��6Wt�kr�k8�Us����y��uh#���z{��{��=���<}���v�m���ӭ���˻�ڞ���yޏrv����U����N�w�{w=�U������{'����g���~?~���ˋ�"Tw,gh��s�_�4L�[��%#Y��
w��N����_�;/��CG	,0�W��T��ɜ{G.(���}�����k�BQ�v�:�M_�O�A31�	E����rݶ_=ZI�'A,��X~����s,�1����{����j��fq[�o[��P���?L:/u��W.������$�o9��]:��(�U�`�-��&e��b1Gk���i�Z	����
�@�Ɠ�p:R�Ԁ�`�F�j1��IEcժ&�crh}��{��o��1)���C���V42�i$l��f�.�@�T�m���d v���s��}���n6!b}�U����ޓ�<����N|��,^T�>���I��9=<$5��Q։�x=_S&�sy�2����ōr;Π}���r���c�8T��g%4�gw�m7���k7��ݛo���h�٪Q.Nb<�<+��ȉA̚�UT~}�a�_��+ͱ�'nWh��pz0�H4��Y�]H�������7&P�����i��<�i�|(���we�O���q�ot��e�N򜱡U��^i'�D�4�n���KQ�*�ld$��u�ˎ��խ����A�ͷ�.����~mw[4Si��XFf,�b�(0r�q��;;��妯'm��vP�W,�e>�7����nvs�|�3��X��������L�.������C������W�f��iI��pܶ���*Im�XdK%a���}[���޷2�����>}��}w|���!7�H~�!� ���HJ��x�O�	�Ad$�	HC�,	�@�$��@	��<dh��O�)�>�>�ā��@�2��3NHf�
�$<` V@�r>�$��H|d��BĄ��!�	��I3	����>0�� V!<B}`I�`$<@>�+��`G�>���	'菑?@���8�C;�l_����������k]���8@x-�� � 8��T�o&sX �p��  �   ���N �JT0�&�     G���  !�z�e[�o���;����T�]��7�=��om��w_>v������6�����-w[K�-ۮ]�3�Q����٧\8��Z7d�v����ܯݷt��xx;uG������8����WsϞ�g��%���w^��K����ջ����m�e���Wyޝ-��7��g5�u��������5[v���^�o/��o9���]o^����쯹�һ{v��[��n��v͵}y���wtsK�J�;r�ӣ۲�{�^s�k����ׯSz�h����ܘ���a���M^�ר��wV��v/d�m���u���:+\��W�.���m����#�^���E��S�o[���=�۽��y�����i�'<�+̦���wu�U���۾n��^�[ׯf��]KY���u��{v]�����k��w�m�ݞ+k��Wv��׌�P�W��Ϧz�:d��"���2��E=D�Ҵ,y��C����i����|�Z3����7��{�s�a���k�bc� �6;N��Jm��=�y/2�x|�7�=������<�.&Q�>x,m�-�ǉR��tM$����鄣�V��Gm/|,��ղ���p����B8aRqVj���7##|I�����a��!I�z������j�*��I%�(6�NI ��ۧ<0E����3O4��5ɼ:*�������,�G3�D��x��.(^x�)b>S��Da�$�{�M0V3���N���T��� Ƥ1qb�շ�\V^�{\iz@	 �	�bȇZ��H�g�봋d��!����4GOB�!�غ�*&�Oƶ���&�ً��p�}Ϫ��d�+yҪ����lP�����5`P� 
P�B�%Db�:�|D��_[�d�Z!o.��/�B�1i�j�1�K`wdm��JY=7`�۰�yA��`�(�س��o}���;�6�W�i53s��@)$�F���Cm�=^�������Gy)�e���D��.� �(�x^;�[�۩��[���n��q�Mc��n�:��C(�%�� ��UV҂ؽ���Z�%n��En�y��W"�p���F��d�A���v/�A1*w�õ�`��j�h���F'xe^rB2�IJ��Y�@!��m�p�i�WL�����?,�R�_�����u�0x�B�Ez�
ۓ�0�$�H�E��
|*�`P�~�e��I��E�vK| �X"�	�e��^C�}gbb�����\�#��k�c�&��(�<`�	2�m"��5���ENLw�n邀�6�P�%E	�DIP� Cm��lVn4��@�����:y��7�:|P�V�`n�qq�{���hYPw��&H3h����2�`��q��I�Zt�53�a3'��N���m4�m��-k>��a$�� �������a�+��*+Hu�72�͓�m�S�3Kۺ6��*�UUm���ϨU��ݶ�ER��   U�{���׽7z[��u�m�T6� � j�T�m����W��@
��ۉ8�*����nOϿX]M�:�r�;�R�-�ۺS�?��xq�(/J2р�囓�:�[+l�Ɂo�ٕ�jo�]�e��3�^7K�i���8�s(z��M���f�d��{�VT�ۼ���Ћ��A��1���1�G�^�z�\�ײ��I7qվڎV{kwn���D���ÉY-6�Q޻9�����'uTq�cF�7�D8�4�K�O��[#6��l ,��=������p?�{|�*��H�R�ӿ��G���L���%3�uu�A��Dș�O����>U+T0�ԍcUlZ���1��������N�lgb�����`��T7�GY�KD��Q�ݥ5T��(J3�rjO�x/}��FEܴ��*��b�+sd����: �DF*ɛ]蛀� 2K���9���ͰU�����I&Q��]�e��PL�T+1�J����Z'l��j
�Ls�����J|�T{=��5�WI+$�2�@�8	�z6��D�"7	�:5�[�<��+��f��eu>�6��ȞQ�%���.�i�� wm�ު���i��]�i�y^���ɗ���>�k}y��u��z{M���U�\.]k�y)j���<R�ګ57wc!�vv�qɯr���%�e�nM�E8����:b?c�����9��+���K�X�� @�˭^��EV���
�I�J	�a������Q*r�1��U��xM�mZ�z�<xH�
Ǥ��;b�ti	;�~Hn���)�i�btn��b"o��	0t)I0*�hAi` �L��P�=f��{^���3>U�j���\,X�n&%{���y.M7DhC�J��m�)%��%	A�>��$�b�����ddo�[6B!�)�Âx�U)\��/� ���G���i�\I�AI,�[&Kf��ւ����U�u���)4	�#+��뾽
l��m�]7*�5T��7<a�f$���mm��	�d;��L��i6����F��#�O������r���e�j�iv�&��!5�q��zk�Op8#/�؇�A�IQ���.���S<�07�lm�~RM�z*��e�mP��g_����	7*Kcl�h��ޱ��ⴿ�B�����	L	Xj��g�$��Me\<r��<?_�����u;�:쫣�<*���@@�܇�^	�"�ֵ�3Z�^A�'ï���>.�V�vAF�m��)��)��&��L�G��O�+��"N����{m\�7�pǄ�8��ɉ��[�pLTnx�vF�����P!��RHi�� �K(�Wp�[j���~�o�u�9�e��96$ToL,b�,�8���$G����((�]�'����I`���-=�$xv�h�-N��N�W�-J�ڹ�����c�X��@��a}3�����h]��#���(�]пM��w��bL��숍�
�_���T�#5<����� 0,-��Eh���!k7nB)��=g�V�(��h�L��N�t+�7阛���_��՞��\W�t��E��R�^$��ў2 m.qj&c��D-ž���6�Aq����3���D�o�N+�r~�;|���4t]\�]��?vZ�o�������I�]�dJ+���#a��FkN�c`EGMy+n��^�d��|�+BE�^/'3���!=���&���b�i�ZH�M lnΛ x ��ݽ�{k�) �7��q�;K�hs�b:��M+���Mw>e�3K|�'d�a��y����Y�G��6�
$II6 ��ݯJ���j�c�V��U1C�(ǋӡ�cхq��}�l�mt���A�Ғ� �����W�\q�KĔ�I�ъ���1}���!�zW�͢F�P��;�,"i ���Hq\�r[��n�1͗W�\m`Έ��J V�I)�{�;9P��"�f��Q��� ��D�b%�p�$��u�SC�=H�Z�<�
�Qۅ5-���|'ӯ��nl��ԛ�UpK3E�Km��LN�Pv�urR�P������z��\�W��La��\i�њaXηt.��H���/��cy
�[�E
�l-qچ:�5w�-I�4��)����m$��-$�$�j�pw+(2X�R��l��k��M�U    �g�m�λ-�����Cl�� T�   l *��R�*�l�Z��l����f�[wkS`��whj� �U�_2�-6�d���h��&�'�{�������9��0D�	ìH)A]�<"�[�\R"��g��a$�l�7�OL�Q;dC!</�,a����x�Nkh�=84���q,�Z���#�s=凗t��X �o�viiD��6�E��"�v����{X�;׬D��[}�Ʃ;�����&�p�~��Le��Iؓ��Ŕ�C��sR����q�;d��:I�@T()�Xa�!���0�,2]gkS�PB,kzݟ7�j���B)�wW�!Ex*�ޟ�����z�T�pг"��7L�ZI2�eŃ�l����6d��+Q���;TW7��p#E��ѥp���=�R"*�]�$Bx�'�K7�|04�!-�J 6�m�B)6껅R�W:ݬ�O�����%*ib��fl�[G�V�E:R���� Q$83ؠ���%;�?pɤd"=�IoOk��QC��5υ�/��������\r_���Yi�*_e�FDgM꼵n����@��HL� ݻ��� ��{����쾖����=���W�sv�5�k�uϽ�9wd�[���i�����f��7'Q�y$oH�یw=�r�PNlB l�l�m����TgrZ�,y zo<��*��N�_rM:����:�3k�Y�)I�	� H�c��'�a�M�l�u�����d^�����c�6
����"��J��^&��$/HƮ[E���j�k�j;���6D��������<!r~��@ Y37)bo���o��	�>}�����t�����3�)�Vm ��F'��G"cK�W��va�n�q�P����:�h߹��J�êhm�3Ϗ�~�$�J��tX�H��P�u��Z@$ۦ�;��[ wB��Z��owj-$�g(�(��*�Cǵ����DC~cɸ�՚pk~pm�����Q�$���{0wC{ʖ��Ùs�D���Bw86{�y���~�4�ތ�~��G�ӹ7K�cy�8��pðQiJka�D�5��i�����;�#��`�b�T���g�cmō̮~���=[�T�%C�����a%/��V�
�u��p�u�֗H������#`P��OQ&���Wcj�q�
o�H �I� ���-&����e����w�gD�W��
;cJ͈����%�o��5�,�Л�K�pv�[�I$$IM��|Y�F��rc����n����D��6C(�W�,\+�u��9���܅���8F�7jy��"�-�L��{�9�J���U*���m"[D��b뎈�Ѧ*QF�8b{���*��1��p������Ѝ��9���sY)3�A���3~i\�0�M"�b��6<���L�o�;y6#Hp���`�s�l��р�f(n�qo�_t���=0�sʕ��ۀl���m�����6�ySU3xM��E�y���s���V�A��I�{�J��m�$��Vxؽ1������f~@b��.�}f��ds��\n��R�r���%N�OX��9z����P!��Ϙ�Xc�Э�8*�T>����.U��V%��E��aP��8��Mfq�F[`����b$k0�iXh�L�] �4k����1�r��F/���m�b��6*g���>6+0�
�ޔ�-�%�BI�gd\����M��-������l����Vڻ�ȶ�$���l�]u�_	v~b��q��k�R�r˓\�<�Q�W���=Wc`p���젡FNش)�NҾ,�y�r�i��i$
���2��ޕ�V��y~��j�<6�׎��/3�Z����Gb�j�����%�>A{+:�/�5�v��<�[p��d1� B����C�\Ƽ510��B�Ii'�;>P��D����}����+�m$؂�0��#o���(������Usm|�]F�7�8q�^#��"/W�7n�����֦f�ׇ�
b�s���AL�V-����k)#)2�*,|Guy����Rs�Dod=`��G�!S��&ex؊&8�)�<ccPL���vpe⌈�{��*���U��00�6d<�/eksQ�����Fՠ��DfR]vm��+j��^�_z���.m��{l�bG�C�"���ܠ.����k���fգ�j51ƌr��Go���H�MJ	��9$���}qg~y��◄ؼ'}�喫�mn$�9w��wn��t��޲�z�D�p��,��Du�j��`�Ȇq�g���+^㫺˦X�`��
�%�"�qE巧*�r�	��י���L�����(ۼpvg\��@��J�����m��{�ڶq[+/��R�1�`�U����*�  mi���v��W��z�>��@*�P���z� �U ol�e�+%�wySd*��7�A� Fu+��\Ż;  ٶU5�bJ� oV�@	�R��P  �V�ڠ  *� P  
�� 
�              nn������wU'�k�{���n�]��-�;j�j��72�5��ַaU�һ�[�v��ww{��Tv�ݻ@   �   \��  T`     PU   �� �P l
�lP    m��T�T  
� 6�T*�@  �    �  �      `�  [w+d*��    m(�U�  T  *�B��y���6�ͨ P�7�   W;6������U/Tvn7�u�}�o߆����z�Q�v��
�T��E트Uz�*��6�   -�{}�)���נ��F��B�M�@� U �� ��7
UU�u�m����߼���U[m��+�w=���I��IB$��6E�Hn;���qq1ꇬ�b2� j=��h[>}Д�8g8wE�oZ�u���zU#z��]��8���IQe�u E��q頜��\%�� )!�b �p�d�֙��H������;����M{/;�2�+ǱJ,F��Ĥ	I"�3�֦R��cE7L��/m��2ho{�'��\
<n3�"�3�8n��q3ǇY���+����V�l�@5�  ���	P *1I4��T�98U8J!W&��6�L�6��{s��GA�.��Hˍ�CJK�u�f �����ʃ&�/�0�cF�f�v�f]ܿdO�+/��h��0����ajI�k��ι�UWtٴ��� �	�H)߆�n�uw�	�B�w.��-C�z����p�:��6�p���H��`4IM��-���f�j:oLu���u�n2ĨĪ���1�6�ɦn�N�^��;�Ҥ�`�I�]z��� ��P�m�u{�:��ڤ��[|�f��]y��ͻ3�k���:mV�^���^wM\t����^���x5�*������kɭw%˶��, �M�
C�@&6ƅ6�x�^�wm��@B���F���}QE٤�A�Ke��-����jV�9^�@ލ����v0��W49��*5D�z����I�
I2xG`���0`�3��gn���9���r7�����I��&w]����'�d��wud��iU޽*-��s��zp� �e���D�Y52=�[�&�;=>v)4�Le�'�B��E���qRN��p��Ö��4Y�#�)0S%6�5޽�ڀb�3-˭gt4ά�}S���^k;	&7@�YKz�@c��IRN�̻�u�Yi$�o22��7�4��86�Z����ݕ�ǌ���a0b��H����K+�`&�)�w�Uۇ�J�"�G"��������ӛ�0_=B<H=8���  ܫ����k`�ww�V@�/|&qV��,l�}��k4<d���H( 1B�R ��n��J1d�\�I���}��w{l��볦g�#��lXۻ����s�J�)������hrKAg7�oD�W!xg��tb8��hŋB��(�m9�=ܣ B�E\��x���Oau^�+�Џ�z��S�~�f`�]щ��gAH$�P9�h�WO���!��h��%��
A"P;�ʫom�{u�ַg���h����|��g%t�RQV}^�a�����g��b<!��B�E]�P�w���*1a� �M#W��Y��|�ƾ����,����C9��U>S�Ǉ�)�7���0�z�Wrћ��t`4	�]����B�
��� �&&���b�k���x������eg`�.b�i1#����E�D���#oaȡ �D�@ i�AU�S/���{�b��a�;qޖ�y
�籽�T�a�f^W�/��zwr �����rg=��(�3o��&zuz����L�{Ӌ �$�)����tLqQ��B2�W^��th��w#Lm@��OW�����AYi&[,�%���z�U^�
�U��%��M�#������D���[�/a��fw�J��6
�, 9fZI8%��I��d��Wxb)��x�&p�՘�-+V_T�W/\ͥ7��������ֿ]Hl�L�e����qƱ��e�.\T.�M��_d�����e�q�$�����z⫐�~��,�Ji$Bs�j5M��C��@F�m���/�p���p+nG7Zf�����|�ry��{<�.��%!�3����9&�	&@g�1��#��,]u��|e�%�!z�zH� �^�q_F��!X2�u꾈����[](d�D����[���V�t�5׌��LGI���z�{����ت��EREn�m��gT���  
�:�;�j�y�<{���
��P� 6�n�d�UClEP+�@��*��],�Ү��`�Êِ��
�I �)��mB���m����f��B{��drf���n�1ۓ��~EFwE�m����&S0F�&	�ʹ��w�wf_E�|}aJ�߶���ѥ��pu>؛�Ѡ�{�h"KtG�%J�4
;�ZiO$�%��,����ߓ�Py�)n��p^�}��;W�:����+&���
(���1����D��OF�
���v}~` �� �Tjp*ȇ `���f�$�9AJ�%���Y���{�h�-���D�8;���q{S�*��1]�i���<LeP�~I@	�	Uw)Lp�a\w<#7�2�_{s�wML���
�<�u���*lݞ�_a:�7�@�CnbD*�Lt\O�w���^U�"͐0I&�iA" A��d�Wϻwh���G�1�'܀�T��\�,�p=�X�^��=~`h�=�0��������̇0�+dH��$�c�c�h��t�}�/�ه�%��8�U�i�Zl+)�x�Uue�~�5����H�HS)Y�7`�{x>��x{�����޽��뻽wս{^oT�O>��y^�9g���Ӻ���]�x���v�^����H<1���z��e�E�"B�E|��W�_<�{;Z4��93Q��,AV�jG����F�e��s�|�ͥH��\N��6Y��a�B/DYWg��xtAl'q:FM���)��|������QB������xY	m�E�6��$�@&�,��]�Ց&�$L !@*SMS�� I��4�)�Mg3�e�n�F��.��l�R�+F�Z�cf�r�H��:2OY����M��%$C�ZN�F�e�G�W��şx��6q���llR�c}j6�Ma�ӂ5���L�x`�,��O+#��ޭ��H����`�jU��I&�P %6�	ւ�n���tS�̫k��b0�}n{/*��B��i��X�v���7c����ٲ��t[�.M��I$�w����?|k�p@��ކ<7q�Ԍء����ōv�Sq��+��+&*�	<�YUC�s?N[�,Z$�ob��qy�5�R�f6`�#T{��G�D�Q�Ԃ��,�!֩t����x�!�9y>���Դ9��R��
��״XCmLxD�*��h��I�	���kpㅕ��/`&. �wes�ݜ�;��^�w�wV������j��E�@�����(� 1���A�^z9G`j��x�P����<h��"�m���"��$-�9�zu��1ԣ�߄"��h�k�ٔ,'����J��ty���e����\�,��E)&�D��4�@'j
����2��#wj����;y4y����GfǍD�Фn�4�%�T;�%BF�Ϭb�ӫ��5���T-"C�>���+�95�<د��ܔ�rL��н;��z�'�tX�B�F��JN�R�͚U�Jv[4�\�%"X��if��˚�c��A���d�e�dL����*�TVR�V���}��*W�$�J.��ŋ�O׸n��ɦE���Qa��y|��K	�����ʽnܯ=O�}�o_���R��Q5Zҥ'�^��\)�=��c������l�������z�0�>'�[7i��&�u2H�ڏj�A�~�?	�'m͛6�M�q�1٨����b;Q���>3���,"eml�6�>��8Fn�c����J�8��
��k�$�H�A,%��@��b�j�ս�C�[.��(U�
���3�c-��e���s}���
�f:�H����sv� �.�W�%� bI�*��b�$���OƖU(���+�e����kdVƃZ�k{�%w���!'1���v�f����vJ6�HkF�����[�5&4�N;w���Ƚ%@W�_���C%�Y�{�<�&�ݻ<��J�V�$�U��G	���T %Z�0_�P@	 *I�� �r>����<�o�=5�����q{N�2�m$9���:e�m:Wbl���m��Ja:�b���F���<N��g�I��*Ʀ���L$����`�sQ�(v�w6e��8��:pta��yW\Ι�k\S��5p���S��c޼V�5�����F�.mEZ96�I!L �ӡIҠ)�+=B�UٵJ��ܘ��*�   ol��9���Y�u����lw  U*�5HU ;���6%A�;�T�ٲf�*��l�s��[���y�e^�J�!� "S`�� 0iV���6��;]3�[����a�j:4�����?���NJf�
�s�q�e�F�@�)Եj	>I$%3UD�+�m�}2�p�69EI����*����Á�	�Z0�|�5�*;���;��I>��X���H)�q�0w�T$_Y9<>a��p�&�`�Mly�Ғ��S��,o��tJ��(��$������4�J-"PLN�6�F���7wWwlַZ{99������!8p�\��a���Be-�`�QÀ�D�������B�qF���)�h�:�q1��GU�Ē���/:���r�S��Uq�9����w@�ƿ!��4W�-(�ͭ�O�۵>��"Jm�v6��m���Y�+He�[I��I�}�f^�z�u�13�K(�Q:��D�����02��Y�$�R'
�%���]��֍�;1˜�&���3Oٻ}T��57+�ȶ�>��aʏ@m�3IZ
�M������4
I�e��i��m���s����ym�������g[yͶ���޾��'$���:��6�qWw��w�u白{oq����yk�ۻ�ͽ۫��ה�I�xD(A0�&R�&,H��������۶���c�## �P8��3�x4
x$�_Fh��QcfOE&�)A2��L1Vr��E��@��*f�}7o7�\V׃�`�t�'�8�ql0�N/�� ���`�0%3 q�;�ٖt-	(-� �B ���6DȔ�D������P��/+��IV� k1�0�M򉽘9_A�<"���$NB1b4\��u ��A���J�Ty��jnLHq���lOWcC2mGk��LSf��G<OI^���,�*�X��GR��XP�P	�����{�AM��E��]�R��I��_q���ms�Be���M�VY7�yblg%����u�Ly+c��}�3^���LY� �$�H	IA���	���0C��^�p�d[��3^>U���Th��a��9%����Ҙ��|��p�-��;�o[�m-m��0��qB@���݈W'zQ��\���_*@/�UE����c��rT��߳{�1<�gk3��Y����f3Xt�`�YgZ���mvu���;*�5�1��%}�b<��aU�e۠4��m��\+�� S[����ٷ���K.�qG��`ڷ�1Ԓ��_ee�ָ+�v��8�f��tl�L$����9�R;��Wy�]˨�E��\���W���:��^%�����cA�ݑ�;���l�/�ͣ�g�;����h{��m�͕��K���L!�6�R�^���0(ݡ\�w�u8�efEpVBq�^����D�ܣ�eq�3s�ef�KX��I�m��n�����6�x � �p��.�ǁ8  � p�P   ��Up�n-� 	�V� @  z�l ���`#ǀ��n^�嶶޳W]9����ܬ����u���nr5�^[q��+=��׮��]s�}�Ϗ8�����/)�n�n�y�=�s����{wW�ݵ�㙞y9��L�9���Dp�c[�����-rcc�h��we�;�]d�ޗ���m۝��8��Ŷ�Nܺ�R�͸�n�۫}�m\w�y�W���w���Gl,���6��ݷwU\ݼp�m޶�������oqצ��/�s����s�����7#��8�WwDm7sگ\�kӗ-f{��w��W\]��ݶ�^g/k�\��<�d��޵y��x�˵��v�N��ޞ;N�S�췺v�뾾����:���8���"�5��՝��򾾻�u��v��̷�y��n>���x�2 P�e�ۂ2ffJ!�6�{�앴�z�:����c��^[N���V�.�Owg;�i@ � �e���s�H��1Tc0�g!��a�{�����Na�&|l��R�i��GA�F�݆`�" '��7N�[���2<]������\�a�ʫ3⍍2�4꼢/N�Э��k8Ó�{�����:�z;@L�xj�[�\V��6Y��t0ك� `y���f�l^F�*�<���1����%�6�j�1(O��������{��v�S��7cZ�T����l��w{����̺G�ٿ�
�ĢF�D�'"h���YK�9O�Bk/��y��'��ɦ7L ś7% �	��pw�`�b���<&)�Q�	=�����n�i�J4�K�\�ňë���LO���h]5�&�M�fH�tM�1�����)<ҧ�9\��s�Z�&߂����<H��9�P#�+��5�\tb�]��ڙR��I ��;�Ԏy�^0��\(DHI ��%��P���0I-�pr'��j�vx���(�@P� ��N$5�}�_d�<����j0;6�5VbS$�*J�#rϽz7d\�78,f�A'�2H�WV��A�`&*����|x[�y���`�*�=]������Ŭ<�WԤ��@��N��q	�:,T�ˤ=t�)u�D ZI��l$·�;m��w
��S�l�ͤ�,SܢƋz�����G������0n��&ư��N��� ���s������Y��boI�p�,_�O7x_��18vg����2�5Jϴ@S���k�>�b����Í�,��ߦW��M�1��{�����;�f4C�a�;7�ԫ5��.
8V�8��-��.�qP~�� �8�!�:0CJo����mW[K�K�zQu��<uP�������S*��gok�x�l95�2�z`1�b� X[qQ�$��o�1b ��.ג!�K��^�f\�>/�Lw��,�S�Un�}�� ��S� 3�7i�{��-n{��m=�Si�Tv]�&��Wj������	�L�b�t�(6]2�d��QT�k%:ҭ�����U �   �^ݫ��o���ۤ�U�U  ڨ��Cl`U*���sU �P nE����+�����[]wo��� �[%Q^����fIe=�W�~oz�Ҵb8w%LN�f3����n��fӂ,��Ŭ�
&7���\b�2I�4�m"���Rcv���U[����ʼ�5�ue�؞�p�> N�Tm��]���9��F��U��s�f��������A�b����.�gOzi\���1b4�Y1��
۬Q�4��!��V��4�7�e�T�3m`�	$8O�\�����J��c{��D� @� ���f	%�H��I�]#/y��̺�P�P� ��,U!�{R��b�5F��Q&�I�^��KQ7w�5 �ʂJy���]�O�L��B��/Ǚ���R�;2�na���6��'�c��i�=�5+㡈�'X��ti�Ry����:�\Wiq:##L�D�m�	"Jm��
�� �Um��r��i#Q��V�GF�\��jC�U 8zM�f.��rvr�>c���o��0�Ͳy�n�AO=)n�C�1�{p�J��O'�V������r��_�D>Ϸ:!��`��θ8��X�`���ٶ�"7�cJ�I�d�iP�^�]Z����g0umv;���m�9f^�90�x]7kj�;�Zݫ���ӫ6����[���g���Kn�����w��v鞳{T&�H4�O�q A1�ׄj��vS��q'jՌ�w�j�JX�����)�u�,���\5�ؐ	�Jj��>v͝�`�Q���Q��,ntԚ(B��h<����c|�m���xa�0��Rf�p8Cv�Ų�$�(��PV�1f��?�+n��f�n�����S�Xm�ɦ�zt���Y�/Td���&������MI���S^�^���)�
Dԩ���*�JszR�q�b��'�1cv���`o�x�~�(��2{̚V'\�i����ď^��G���
��̜z��p?&a$JL��v���EJ��fn��L��I�����{��]d�������0xk�
��;���!�1�c��l�a�Z�n��"�RUv(����)W�Qb$l����^��\W�����M�����"b�T,�\0��단>��Мʼ��>�[I��I���Q0��fz�M뻍�7���;<g��A���l��㙻r�0T�����V)N�C�WP��F���6d���ĸ֫�-N��D����4P�J��w{��z9]=��z��<L 'o�����wTvtZ�Y�{���hF��lz*�����;��)3;�k�8��0�OыϮ_�}c�g�'E��iS��̻��kk�*����ob�0���vJ��~�܋���!"RM��%�	�uAM��U�����@����[��¶��^�%qޔo��@��z��?Y��d+)��1���F˂I-��kC&��n�gp����a�����j�_�_a0ﺫ:�d�(��ׂ���+�ܵm[�,��M����¼5�#W�b�e�|���O:�����^V���̉D�Hۂ���{�˅��$�(D��0-�G�XP�)&a����ڠw��r�Nt.b��h�$������"B��r�y��ufa뤝]5ֲ�i��s���QJ&�����Y�A)[�b4�!�-NlmVள�\��׮��[�w̢�gH�n��M02��VWx���n�\��T�L���0�,�m�[k{�n�ԅ��w;��w&�!!�[�9lO���G�������w�����^[����E���I�����g����%c&�q������jr��z��)��zű�zxR}m%�Ѧ0Ʀ_iR�"b��U\����$�P��c�Μ���f%.�dx�ɞOk��,�����!�ѯ|)3>�3���Ș���	��ރ��)$�l���l}zp�ր

4
�SS�ҽ;���W�/���)r�g/^M�%�o�j�J��\�@o3ˤV�L���������+�q"N&�F^^M�d��nl=���@�9R�Wl�����]�����ȩDm�de�Nj����荌��%�8�
�#��򱜣c�yM(��	���u��w�M赌�9Ѡ�4'6nM�%�Ż�Km�ܽ����*���s�w{eR�U�T�P   �v|�v̮��� ��K� Vڨ.j�J�m���;�P�*�c/M��݋�^����;B7���ʥ[b�Ewmwn9UL���,����K�4��g�^�*����~r����oT����=l秔d��f֯��´��)�Bh��16cG�Wx�}f��.��1h�D�%�cܕ��{����:&|9��!ГU��.��,��@ E�Q�bG?+|٧��I�1v�:X*1.#����8�		���� z,�-�$�U�:�N�)Ҝ�_<��	I�)Tv�2lM܄��%|A��m"�d��D�"I0!��z���F����x.�"���AR;�*OP�����\��}��)�3�MýU�ӥ��E#V'�C�1�6Y�����b�)�3���LTD��*��	�BbĊ�$�-6wt��%��R��.3�+MVi���1}W	Sh�h��f
͕ �*�*6˺��$���c�qg������;����i =����t�0g�j� ���&�� X[;hℓ�1�(gr�x"v(�&�{	�4�J��4��h��W>λ�
#�J��1S�ܐ���d�����swiRI"�m��m��m��z�e��,kn˺���sy��gg�;���Mj޴�W�<�ק��7�ɺ��mޖ��6�u����k����U��y֭���e�;k{v1pP��	 PD�c�þޒWzkA�1=�FZ�z�(w�!˶7�y�=����'��t���u��[����sX�����w롈!�LT$�8���+.=�z�	�1'���N�n��nH.;lt�d5BH��Z�s����)��=t�s���cd�$�0 !���H0 �������v$n��F��q�k]"��(��FN´�Ov��|r(��1��}�
�ߤP��U�4�H8LNw .�p��\{��]����)�[�����M�r�-%��ʨ���H7�0���q�R3Ƣ��	�6G��HϺ�J��- �6�]���K���R�������O@��8�[�t�O$R��ۻ�ͷ�ς�]����޷��2tu��Յ����Sڱl��Qr,�m2��^�6���/��>����� J� �Fq _S������3��]��ν�+i����@u&�n㍧f�Sm$b���P�w	$-�G	������(T�a�kt��W�9i��L�Qmn�!���[���]bc�@F����Ӿ�#�!=D����i�I�W�Daϣ��@4;�z˫�^���v
�k۶w{��{��N/��H�o���k;�.�L�;���pT�U'��ɤ��{����6��*Ō�%6�MD�w%�K�Ȟ%S@��­�׿X[��s'����~j'�VI=�x�N�yb{<0�MZF�b��ky�a$�I��)�KǷ��b��[�/���ۙI �=cN��}G�gk �k���c��b}f=F4c15��<��M����V���8t2�$�`���B�JM�R�&�!9��vc�(�]�Eeɹ�-�XUuCL���Rί7Q�(!��@����9n��h���u$� �)&��u���V%(@꾞�Z�>
Ɔ�W�	����*{>�tc�gO	�	C��p����qz��^�% �!�[+Ѿ��-#�KBF�����
 ���`��&�p��vݳ�móg�����g:xw�L��9��nz a[˱��0�c.ȹ�����U�J�����z�����J��}$wy9��ٝ�$0S$�����i,%�����s��lK�"���@��!;G<4`3e	���h�}��!;��{(M�¹�b��?�m�KP6���Ӳ�c[B��m �L"�I2�1~�)�P�
s��f�a��xp�	��g�kmg�#�S'�>�%m�Wn�YO8�ߴ�vc�ٛ Z�Je�b����z�Q��/`=��܀(1}{���ϑ�U��v�7�Q�;&��/t�A�P2��t��Lm(&,rM$ 0l�a��_)r���c��y���3 �b�1�U��s���$����}���"�� �q�$;D2�8�ݟ2r��X�$�@b� ��IA)8l@O�T��B[�^���m����g(��b�b��(w�V�YÌ�S{l�%��(��D�x��vd7�cH���h�"����Ɏ8)��NЭ�}�����4$`�;|V6�Jd�Ԇ{�`�q�����xF�5���"s^���T�.�����yF���wo��f(��㙭��K&��;M��,�PI����^Čⲳ9a��ܮ�C����d�|�V��z/oWZYa��H�8SJ���O2(]7T�u(&:�I�}�7����3sM�z�������V�=.�}s��Tr)��B�m �Qau}����:ʤ� �x��P���qJ�ؖ� wI�5p.\^u�ĵ�ɺw6�]IM�
9�X%e_0�ɖx�q�JK�t��/����&q���V�jpe�,�ͧ��w��Gr�@Wul�Q�6C�i��m��m��l <n��������=���wk^ώ\�8� �m���u@ ��  ���-�ATj��*�� *�� ����7�vv�  �e-�l>k� 7 n�l  �/���m�  fSl*��  d  U  P                 {��n޶�m=��o;U7���v��$��q6m�m�t��uu��vWW�ܷ�F���3��z�7v�   uP  δ    `  �  T   
� @-�  ["�
�    
�=@�J� *U 6�l�@   �    
�         ��   ,�Z� �    �UU     � U�*�{yv�� '[
�����ڀ >����SaR�lx �N��S��-�U-��8pa86�PRh�(��=��ې*��B�l�   �lgk�c�{��=j�.����lx� U*�+%@�� @�Ql�AVu��)l�J����-��Wu�{���TWu �w}������1Txv�Ӣu��1B,����<á«g�D���fjV9g��Ud(�7�b����-��=&75\�
C!��jc�.�ŎJ��b��ze/^*����)��yX�ڤ;�L���R�W34�K/gSo<>���'lx���fͤIM&�7Q�e!�8��}"{�[�p��n�!+�����{j��@�����할��vB%7�8�o��[��s�Rƌ'Aब�@���>=ȻZ=u�j���t���T��x7f:}
0paz;�������r�O�8?��zDV�b��:΁��#��Ef�p�����A%�'���U�xt'��b��{���G%���sc'�v��Cg�X��nM�ـlw�4&/LP�5}���"@6�"����ܢ���me*���D��.�� +��;��(\��dV��J�gG+�(������f�T�=]�t"�I��Dr7V�_��
Z$'1,�]�BQ���[�]���*ۢbhT'J�
�ޜ����ݪ]m;�����֠;��-�V�m�˻׻��nܹ�gv��g��-��]����lʞ.�{��q�ݾ�{v��v�iw{o<��}yݷZʛ�x�����|��s��=�z����wŜ��Ba~���h�Wc�M���L��B뎌ZJ+`	���V��x���-��I7>�*���#��C��cY��xhQ"�@"�5��5*�}�D�^C:�I�#$i�wa����)�[��&φ���M-��uV�w]��۝��n�5��t���!�xvr-4\���c7zgmLR��2�e�-^�V%���	�jb7�T߭"�H�m31���	���,�)�)�*�?�����y^�[c~�c�4��l�Q���t$S���Iҳ�r��A{�-[���`���d�T��-�m�Y�%&	6��t4+&y��� �T[:V(z"ߺ{�h.a��LH�+�2y��wņS�5~��霩���@&�E@�ō:w[�r�w��7��<2�4 v3ͣZ�N���!o7x�K���Ry���F��n-���� $�l�����[׾E���TȡE��;�cR��jT�ډ��J�s���`�em�M�����--���`�>�l��W�w�S�dU����}����!�KO��Ϥ���6]����g�g9I[p�j�w�J���}1��k�N���sF;���^�K<"�����2wA�N���˥ϔ�!`k@kmQLLo��zMw-�m�p������W�#�SX�riu.�Gx�Lߒ���nL��y�;�+� �Q�2 `�u������ʽ��ݽԪpUWn��3�?���o���.UȽ���l3�xf#�u��+ou^�=�k�Z����B��{�P���"�m$���d]^�R�e��2+�b=%t�1��&Wr�'v,�Gy�"{��u�S��h�x]f�#ؒd��<�՛��zF���d�����y;��(��ַ��ȕK����U��KE��k������a%0[�	�Y��k��8$�YK��k~�]ل�0�Ðs��8�w���)���ك��,�m�ϛ��'V�]��ھː�k��|����>E��(f��X�Q1-"� ��G@�<�{���������_&U���
I��F�[�p:E�&���@ᗄ_���&�I�$����UV�U�Uݺ%�wYX��q�,�n�Q�cu*fF���CRh��i�.	�2�MN��q����Y�ie�&��H>�}y�T64�M7cᘪ��r<����Z/#�K|�]J����*mm�A��F��um#�q��: �`42�ƸnbZ�(E$��eѺ��0�����rL_!d����ݎC�k�p��o1�-ήi���h	�ēX��3i�d���j���*�xGt}�s'5a" ����l@`�~)��	 �b��.�≱L՞L�@8C+O:C�ֵ�\��z���A퀒�'~qR��K��I0�3�=f����d�̖�<H�(�E����-��*'���N��Z�|g Ӯ5s1��f�� n�|�j����h�+I��fZ<�
���۠Ѫ-�=��T�*��jnoc �p
�P�   ��w��Ǯ:�=|�P��*�ڨT� `*��� @QT x +�Ql��r^�uN����`�+%Sc)TŠCa2m���	�6]s���k��Z�ؕC���{]<��F�j�T1�/���w�I�	�1�ҲO9ậ2HVSD�\pP<#ηvs�<��4u�����ѭ�PtÜ��������'HO#z�_xh�F\��b�@QI&YF&��1���Ҫ�\���$$`���^��Q����2����z D���u�yܑE��k�r�i���*
G�	�u���r�iBI!(Qa�("�Q�,��㳛�y���4$	��w qXrwe1^�p h����F����TiW�*$���N�^˃���%���]-��]*
�s�RJ{9�V�=bq��h4(�{G�z�p4���P�b�jl���S{��l�m껨y;�6@�6�m��H��� ��e$��q(�Q��*�`ZE��S2���w�� �u�2b��������7c�.R�=��:���H�6z��2Q$�SU��#w1�v��ѷ�^l�2�˛�ێ�5�{AC����r�ܫ��_�J���_�W;m ���]YP�P�{7�g=���gsz����7q��k�o:u;�]ϝ���9z�z������r��9w}���hO�u�ݏo��o��Q(����=����Î���_�CqJy���U@`�7�-}��˂`�F�1~�l��Ʒ�����rI�&]M�#C�|�U�}n���S�n0!�"���얕n.�@W�u�����	n�����@F��4RI��.
�cÎ��E��� ��4X6�I�P ����#�D�OD�b�o�tL�����|�)-`��2�`��u2J���)�����ɿ�)0�̸�F[���{x]��5J:gӕf���Lp��*��zc�!�œ��Z��^�n��c���� Ou`�v��;jl�(��m�� D4�	�aǝyr�����c�cF�*3��|�z���r����-=��r����Gt%\?&��ɌG�ŉ>H-�W
�Q݁��ܙ��	0r�-7��
�.$ǖ7�%�����vxA�����T��\z]NW��Y= �^ݴ�I$f�DWyM�F(�F������q�������\u6b��aJ�FgǨ���F�7yba�����~��kQ85ת8G�+go����h]�B.H]�a���B}\�.t��Y�--�(�0�0��	��@&�)��)�{eGgDF�@�	>�C�4�B�Ӱl�rV��||6���Wd�4�E��I(I���ל����`��p�Y�n�co�A7�z�C)BR�G(ǭ�f�Ǭn�F�gDC��8��C-$�I$�$��I�P�T�l�u�-�7|x�P]��a)OM�̜v�e(^U`�`5>K��k0�w^^.�b\1�;�Hm�~��N��-��%s>��"o�3k��b����݆�Y5� h&t�(�C4n��	Y<������٢�I�J������WG��w�J:��]׌�)�1�7�<J��o\2߷'��m_�W$�r4�J��.���IB��0�
,�@ ~.�AP��ծMd)|�΋;cv��ft��Ⱥ~��|������[�Z+r�[��t��h����>-��99�&�P����Ą�m���4GaO���8�?p#z��η��5uJY���+�v>��H�D�3��|�p�3=o���0�ɘ�R��m��}��_�� +m]�wZ�ఠ�=" �)�����7�b�3�7X��Eso��F5�~]�Q7�g�OP�/sG�������Bݢ�d��W3�k5˾�W��6D����s�0����*z+Gq�0�<./��E�F�t-�㨍h���&�-��T�{T0�rF
"o˽<�N�{�dH�6yK���b�����5 [�g�x~���C�I�7>��1�Q��-�cӠ���D0�a�Ђ@�8�C(���Ƥp���ߟ����'�>����;R��7 ��&e�q�Qj0%'+ �J�8FYۡb�	�˄�+���
4�KB�w�=��7*\�3۰Us��xI�b���f����ᦕ�=�(r�S{���d��OOO�ho����+Wph�V+�;�X�i��-�Vef�ݜ�T���ak��f�QwWun�fٝ��YրU    ��q��;�/�o���
���m�@m��PT6�T���
��~ͯ�U��q����u�muW~����uQUV�E��&�h��n
�A��#��oh��}������ڠ��oky2��E��o��r�;��w�T3���z� m��	/����0<�xm�{���'��y�"�ӏg]Z�K�FiчP�q��8��W�.�u��Q�ᇮ�!H�� xo�g�r8��Z�G����Tۋf�nØ��#��OL��fNr�&�c5.!2\ő��	��@��%6�)��c�4�X3R�ۄ -k�����{�)�z�휒���������7-'��8=���X9{a}�{wf��ö������.륥����h�M��IFaI���|�=&s�,�UHJ|c�N��C�,n��)�-i����)�!�H��.�3i���!6Im��i 6űJ������H�嫛Q�$t��4=$nm(�G��`0��=�J�w���q>v6�`��E���]J��i$�6v7�=�M
|U�����6����)=ٚ{�~.�o�m����p�\;�ҥU���o`����;�ͥU�g��u�Է�\�)�L��I�a�Bg�҂Ɂ:�����s=�j���}�ݤ���;�v�6�W�֎���#f������}z��un�����8�$�1��u_'���yw�;���c��a���Z�.�λFmU(^d�m"�k={�����i�QZ�������]�\�ͱ÷ٮ�v��'���ȶ��ު���!��$��f���̔�	$G�"��'����f��u�td�;���.�Grk��Q���2�^�n�����<�*abؒm$CF� ��ə� :?`�����Y�Ձ�5�D1քʽJ��Z`ݎ`���[���UR]�wj���~��{��T��m��D" %����yW���7~�\(��Y+�ș���!��U0�p��Od����w�Q ��$�E���W�-�Ewt�NF�7�}X�L�[��)uq�êI�bu�U�I��u�mr� ?bD2�6�u�^z�N���:n�ɒ�2>���%����qu�A��f��JX��NvL�:hf�S�S:��T�c:�j��+�s�e�:*p]ڴ�2�2��WDb ���k{�gX��� �<�,�T�:j�����i[.��nir�δlV��s��Z�.�v�gm��O�g�FJ	��ۋ�k���j��ee��O���7&�˥�R�ѷ��C5�sL�L��=RK���L�3���v%Z�.�͖��[�ZŃ!v�ղ`B�,�޽q���ys�&ko�f�go;��C����@�pM
؍wgKKwx[;z�v44��yu�yC��T�R��������7���?���0�  ��ӻ׏��  N T�  w�*Z� <   ��y    �=�C�@�z ��x
�Wn�z���v��}ݹ�V嶛E�8]�e�^.�u���ں�wi�wZ�n��[W]�z���1wݹ�_[{�������L�4�ݳZ�Ƶ����{'�{��ٮ�K�͹z嗭�k���y��ݶǷ�mu���;W�m�wm����m{S��U7S^Zwn�<��y��JW�v6��q��=;�L���3��om.�������۪�W��W�Z��e��������{��{����;u�{�ڜ�/uL��V�V�7v��[��z�=�q����t����m��w��N�]�m��ƥ:�s�v�Z+˪�����6�{���m���z����e�}��n仼���g��{wv�wp�����S�iŻ���奧[܎)�n�5+v-up�׷^������wS��s��u���-z�[i������E��=�N��^��W�ُ�N1�q��������h�>��.bBȻNEV˰M��N��I�{�� V�!�HB��6`��!� �LY��B��q��5ŀ,����s��@��3 *�i��\Y�p!�U�@I:#�d�*�Pm�L�w0=�E�i{�c��5��������h@񌅅Jr1:1�cm�^�:�Jn��¯w�܃׹��)�Rd��TUݶ�U*�m��2�$�m�/0��+i%�l�=�e>�QW�5�ǉ]	F.�ݧ+�y�k]�u�����P�xRs��vL �ݒ��l3W$,'�zU��$*�;��(po��u����,�����2��%1� ��c3.���(�i@�<���4�s]��x�Q���f��~oW$��i�wc�݀1-B�U���i%��w�O\"j���Q�nJ�oe9�:����d�"��#M�mu,��b,��|�+�8�z;�؈_���{c�N�nV����9_����H
��� ���+�\�$����)$�`�A�r�gd���wƥ>�X۾^��#_z+����? �zw�W5��BnR�(N�hS���R)-~M�[l/ͦ�I���~������:�h����������X܀T�����M�z�mԸ4tBj��1�&<�h�V�nmy�����.K��<$M��s#��ZI(Jv�:Qܔ`��0�
��70���魡���p<d�ZW��j=ִ_v{��L�ڞ�1��AP쀨I��i�^�#Z�P,N�ġ�Gor�*k�:M?<\,{g+q�q-y��A�,n��-�bܡ=��ںb�y+��*�l�t���0�v��ص 䀀�3��PCPa��h����[�b����l��*&�O����q  ;��S�@�^q��T�&������<�kox�3Gj��[�J�Sl�s���!˘�U �ܭ�%Z��צ�b�$f���v����4`b���Q���EZ[�y��	�'�_wb�Z��0�9KdD�D�v]�ê�[z�:^&�t��)P���[�v+(6�Ⱥ�Swp�]��d�P@   -꼖/m��8�v�Ol��l6mA��Um�  p6����Tw �l�{���©]n����-�ݲ�UwP[f֛+n� 
�$�i �!���FM#���?�}�Ǥ��V��a�tF+onRb��Z�}�r�NY`�W�3S�ȶ�x��x�1,�d��I$HA��,K9��܊ٍ�3��x1r�+��:�S����o �Y�����1)�Up�ˋ��,ȳ�����PqQǁ�����g�8HW�%���JHP�Ҟ���<&���g��2��� Je��}���C�"�d��W]6�x�[d��n���k�.u���ǹC��u�0 �+5�����n&��]�|h�4x=�O&qt����$I���	mu��ߎ��Ķ 	�W�Z�aH=&`nd����NO�5�N�jUlf�c`m�ù��<�Ugh�)r! S��ɮ6�nN�p	8�"����w(��m �+�st�A��2j�{�8!���i{�\�z���Ei������C�Mŋu���T���ۡ�YH@M�뽞��y��'}<r_[�6�5�p?]]H��l{���W��~��#�j��wo@����lQ巹v��^۷�������z�����޻��h�m�����:���}��vn&��g�k�}�����.�뽃�Du����<pwg�V�5�Y,��-�[�.�MUzJ�hC�oy3<kp��>�im�z�N�A}+��n��bP��{m2d#�����8����=�o�IǼ�v)����q�%mC#��"�h`�7������;+ږYټq�yZPm��H�H�o�˜Y%��PY0�AB_ (	� �D2?Ѻ���������I�C��Jz�6�h��V�����-׳�	D'���Q`��&�JP�$�<X�#����0]U�E=���s'u�7@�.Z�n�����Ú�<7O��{ ��U[k�m���7J�;��$����)�
fȊ�w�%�FO)��`d��6��j���*ho� �*�xz��|/�֊ɽ�ނRiP�o"�|�"$������7��@z�@�zsٝ0b �

�Ɠ3JF�����IOU4�.4�Jn6q.���\|��c	���m%��y�����Q��X\/E"0y���Pz��/��rw��ژɈ��1)����F����y�^:|�G�O���:�� �dG�@��Q�u[6�i�L��4X��(��c���&� �@@J��a�A�*�eR�ZM�=В�f*�Q�`�*411�sw-�ܩ�>����UcPf�l���x=@����x�$L&�I����5ד�Z���J����F8�^0!�վi�n��p����	��W�JwK�,7>m$�$����6@� U��m�)�YO�^��cw5���b<-�+�Ec�{Ո�@�Oڥ&�j�B)��f�s�����$���$آa�W.b�H�- xmMCj��Msm�܉���6~)i�O1�d^�v�OB9+3��a�	X�M�BI��b ��}[ȯO��QB����u�����z+�޸�]�0���7��i�-)\�9��tS��2/� p�I0�b�,��i6 Ł��
/-�֪���G^�����~��v�7�Qa��*�����t@��<�>"�$�*�#�GP�-���X�m�O�F:X0f�Wl�@�Q	;�����}f�$�؞*Z����������'2�Ss/M�^����Z	�|hvF�v3#���P�aʱ�8ߢ�2^�&�M��{jl^-EV�ʅ�U�"��I2۵�����37g�N"�T��7�z�^����N,��1�Z�}e���{�֠3�����ր�n���+pen$(&�)��xAt*	f�����"�^O{uZc���}[B�E��HF,>�a�doIM�^�-�9ӬoJ[�!��31�l8��	��=U�pOB��\N<U�w�ݢ��b�Y��\�n�f�a7ZO��7���	d���ZdLhn��Z��a(,$\	��� ���P"Y�|؅٧5��2���;Q��?`3,y��t��VpJd��4�K�y��{�r�"Jr���xMvNu�F�aD�c�
@�I�Y��������;��VD7��x��ʔ4zc�e����\��'w5��Z���=�:�����g��suX�[C�a*�r������m�m�(�RN����n �+6����sU U��[eP  ���k69�;wq�
���m�@ m�� C� *�
��U �͑l�������gw���8`��nvUC�U-��ܡ �I[m&c�G
g�tec���dR
4�� V�����8f���U�Bo4�L��ژ��ѷ��%$��u�x�/|U{�H�r\�@�4���ވ�21�C����E^	��Īe�r{T��&KM�)�B��w}���f	�R�\��ԕ7��z�΁���u��|������\==��-%O͠�I$��K�b�.15wU��ڿ�^����Y^k�&Px�Ǆ�Қ��U��TI�7�څ>�w�T�y��o�Q!͕m �ILm�5Kg���R$j.A�ȝ%G�&�d��r5I������s쁝Bn�G�����z�h�����wm��tw4�� $��PM��%$�,��ďq����'����y��0<5� �ud��͎OI�ʚ.�C`^����S5
8�6�'K6QR�D$T����=/}93��k��`���Ϋ�]�%�4�	x��Ie��2��U����^����=:�T�띻t �׃�@6�8���ziu{O����/ٵ�wN���e�q��ug��{^�;s�K��7��iյ����^SZk�7uq�wa���':�� CA� n(�:c��<&�� ��e(c�`�Dy~Qx9�S��TD�s0��I&[�#I��;P�Ӄt��ESi\��W٦��O�\4H�o+���9k�fo���� e��f���V�T  h0�w^��w�^�O-z�Y���_뷑]Q�tV��n��ӎ��=z!`�e���]�I)��KSm�Ȩ�$q�Ԓ,�-U|r�OWy̩��l���S��f���Nr�6��D�N@.V�eT�`PrN�޸�62J�ޣ�����o��v��Խ�EU[hR�V��n�UR_߿��_aO��m�\&��`ymhi��:7_��%��_�`#3��T�Hus�PI�@�(�:�IV�6�M�C�n/
��S��h�p8��"��{�&�Rl�Cfj���>�cw�P��h����ggðLb�e�D��H4����Ԑ��Gt8��T�ss;��^��;�:��o�*�D|wZ�e��lq]��\�qp�L��������2�V8.���Va:IR{9�A���/�b��ҝ�rv����<S���d�5Hb��f���s9S �z��5�0wo��_��yWq�
\��I$��d_��֯��� �Q7� 9:&�2�oh��R��T9�\Ť�[���U�WG�7<��U"�����K��8����	��D^�g@��e�Q@G�ZC��;��Q 6�R�I2X@e�m��Z��C��q!N&���E#��G���_yh��yם�2&VR�#Ոm(�d[���L'0A�k�ȳ��"�x!��<���Ə�gi	���yG_3�Y5�`�.�d�*�z�1#�#5!��P.0./I�2(��%�%�{��<�COX��5j�Y�V�q�:��3�&�L��&hC���ۭE=���I�����F�"��	i%Mt����#������|�F�S�k2����q�y�$��}����l|F�%P��\4n�	�\谹����f�x�M�Z ���}�yw!�������MF�#s�&�$��C�U���P�m�4�Q��Q��Bg��*�#p��wۃ�B�gI���y*�鶅��_K U�ex���A���r۔�=�A�R]�]��6@� TIB)��d��A&2Ŏ���h�ZkR�X.�d{UUy��
)7I����z����q�t���ذ:-,��HEo%Ww�m%" u䡎pXŪ��:Z(EV�텛7��Wh;E/O�<�C���:
NpJz�^h'��d��t�L]{��Y#��&o�����#�yOP�_[]�V��V�v�1�<�$ԯ�(�rː����~��R(W	�:�� �SH�	�	e� ��I
Ӹ�K��� ���B4��ct͙�D�++�a��'�<ԕK}b��>�9V���ݠI���t.���^OW��O����j�=�ʗ#��K 2�E�M��	�@�Jި� �Lg\(rw�b"�@�*{_l��<�n���}�RZ���j�赮̢�%��*F��R�N���{]h�t�ʻI��4k����JPm sCݹ.�m��z��;�9�����F)x�m��&?�E6�vj24�BӲ�o����%�D��[��5�p𳍃�F�]µ����vҾ��2����ӈv����oJN��{���	�_n��إj��ȿv��ݠɻ�.nR�:�%�SB�S���,�`8W���Q�-�&����J|�z����J7�(`���4.��Yv�::�Ή$�5s���5x����_��+�\��q��@   7Zw�wnW-��T����ow<���p U�Sm좀P[j��T�۰��@�    *�*�Y���
�l T���{�=� �` QT+m@y[[U�  jq/Y@      
�  �                 ��]�P�����	?6 �!B�)1\�;�[o3��Z��G����{�w;�uo���v�M�em�/v�   8   �    0  T       J�P �  mT     � �ٿs�~�'    0  �T  ^�    VP        ��<   ��N`
�P-� 
�UP�,�    *�� 6u���5J�핷�� a��e�  �m��c�6�Wy����uu�զ���?��۶�NUտ�����@m�]��u6�7n�k�*�   ]���mݽ���s����m�l;�`�EP �   � US� <�U^��[�{��19��vg(*����ks���N���������˟ߔ�-Ϣ�k*���nj���h�&��N���5��y�<Z oG��"�U&�h���"���$�ٕ�EyiP�Rя�7�x�wcK�W���h��V&`1��3i,��� �w�}�^�+�u����@4��e��ZVX���9�d{�ܮ�<�,�7�Nz*�w��k`T޷�A7���TLgw5V �/�/LZ�����i���y��50wd$�����n�[����۵�Ӻ�d��^A򱺏C��X� 䰧��^���#k�]M�b��J��}(�KӰ�Q���7�A�� 3�]��/�T�)%�/���>W��(�kSƶ~~"Һ'!�$��@�AYt[ة�f4M���ݻ�h���dl� �7���"`�$2��C�\�� le*����,�CE	�Ǉ��T��rkZX��*����b���HL�������i��WPf�Um(�:��x�^trD���k���Ԏb�Z�*�JI�Ĥƈ�m�a�!����7zaç��å��n�����K-�I$��L� ����8����=�w;��wl�{]�'>���*\��۽U�^�Uۍ��ǂ��:w�9m������ݷv�f�s���u[���z�Wm��OŠ��@d�C���#0�5'���~�cyP�j��73��Ӡ�<���:���G��-������3F+R6�LO0&��:�<!��E�T���l�>��ٝz6mY��WJ������$�*�4�'N��3L���[�Q3�[�_G����u�/��T��û��^�
�*�C
��NW��%/4�i���p�5Uc�{U�0��T�%��)���+���f��y%����S[���S�(Y�c��j�Lj�F��9�W2 e8��Lu�E�)�n� �=f��;o�f��Л(��G�����������m�mU�
]6U^ �H��@A��I��	z�s�#:��к���=��VL���q8ij���IU@�({s�w�f<D��Jj:��	�w��-qu`uى酹$|��z��43�9�:���Q�:5��`�1F'�P��9����&��#�wT7�l��L��$�,�'��v+|S�Kĕ�$q����W�3���^�%TFP(��22]��*L�:PJ}j:�A#X���ݍH4� 7
mo��+-6�62�c�����sh� �h�D&i!M*L'	�j[~��-���F��#9+�!&'L]y"nctZT�9�RG%5{�����spf�����Zj�6�	����,GQ��{�3qwd��:�����ż(�F�W�#~'�
9I��y�����a���(�~��;��q͝�u�mm7����k���l^ޜ���*6����<M�NI����V(�<,f����B$X�(̞�8�l3��hVC���(�k)�5����B�Z4�"m(���qL��^�}b�ϫʘ�1��Ru�a��Ç�,,�/�W��j�tz-���/X���T�G+�Z��I4��Ɖ�>�ژE8,ia H��Kb�P�[��o�p���AL
�!֘�Md4'���g8w׷4��FL�G i"Ӯ�H쬻���
�AL�i�C �H|���I!%"Y�a5�,�����En��s}�T��(��ld]q��X��A�`���5# Gv�Eu_�����-�˙w��+I��6A��./}��o>��P�hn���II�w@�Z���6��&(Ews��1�o��L��Ӕ��Q�ҙ=o4���}{�F�r�&=�a)���bz��BQ�(V��6Ѹ��wlU"Zm�0�-"KI9�ܖ�Ev%���Z��㔣������A]�@)��`ݾ�h3	,q�����0�+6*E��׋x܈��H�l4K���O4��^س�Q��{�.�7��u��ҞS�T���'��[|�*��o�7�Ǫ�o:ߥLK]~��O$��B(�`���W�����L��5�6"AQy�O�̼u<ĥ��x�z�q��&#=�쯈M5(3(V\U�#�1$
���@� x�H1� C 2�6U� �4�2�KS�|ʤ�<�p��)(�k���l�T�K:��2�V��%�WdoL�H������^�(� �D���=�`��6��'�d��ǳ1������-�9�+�(�j^��Jn���	(m�\���в�f��ޜT~D:P&aԢ��s�	fs�%�����,��`��FE�V��*�UQ�jTU   v��g1y�׎�����E�6� *�U@m� �
��� *���
�������^�ߦ��Yvs�m�ݕ���YUw [*�����I$�l;��1���Rqg~�¢�
����r���F�1d�y�z}��X�$d+]ǎ�S�Z��?f�Z�B�{F�a���M�+;K~�2�W�С_�p�En	��^�B���v�/V�ISV��pu^%*����j���m�[I"���Qc��`h$N�V=��H2��R|�Y.,���D_[�5k��G�O1�.�9l�@}���_��6�I"�;�8�Ѽ*0�ϭ�����ޟ=�y���.�O�8Jج��ٕ�㠊���C� g�&�l�C�(�!\���#��~��&
n㨄oJ~W����iC	11��-�4D�t�NjU~����+$s�U�Y�V����]d3ĻN�/�
i�/��#MsژX0V��D�H$SM�;�XUw@n��B@��H4cˏ���GN�ţ�{���,]h,F:U�'F�1��=K$�K�o;�($�I�6�t���� D�Blz��$�攧�o+��ˣﾚ���Ⴘ�w#�e�D.ʚ4/�;v�=��8@6�x6m@*�u����-��]t�_�{����y��O��ʻ7���h����۶�s7Omw����ˎ\����^)�wV�9F�q�:��^7�1뛻�yk���w��J�D�Q�ig~O�n��OJ�^�Z���yţ<����`��#W3;��f. �ƒa6��ߕ�������O��Q�J��R�
�/���w%*�B�w�b�zƫ��ĉ�Ryx��W��Aw'f`��$Iif�ڢ�RFr�9d�
P(�D!D:B�@*� �H@�R���R��L�eЅx������QQׁ̉�&��{������~�®��6�BD7�t{��䟮�
�JI��5���4%�}B�X��9Y��$UF�k��Y��;365+�E������p)�'����ǽ�T훔 ��H�%��[����*��{�wF�Lz�X�1�wOI�EÊ�q���9sJy�����rV�25�,�Ư{2����.8'wԸ��m�ڎNkS&��JB	%U�|��d#�ī�]��A��I�{3�PB�~�DD�sj6�ZH��r4k�LP8��cI�qX93�����j���05T'����V�9UR��(��s�hE�;Li(ܞb{�]��olqk��q�U(�<://m5>�uQ$eQ>���P��E<�����x�&��]]}�)���M����;*/<M2����^h�(H�HMM"��f�"�E!���΃a�vu�H0c�nj=��y��c��<UH������	i����w�<e^� �y3k)`�o�j����l�X�	��b���-i@&�|��Blsġ�Q��q_*��IG���V�Ɯ���z�
%'=;/h]���$��F�Q@�7���D��i �����Sd5B���wy�i�-$Xv�ɽN �ۊ'{��!G �{����	����8�X���Hޑ��� #�v��J/�ކ�{ct�a��W� 0&:-些�*�%5U  i_0.���0i�����$�%�$m4��H�k��$ "�*2�_5�*��1й$��$�^y10Ц��I$�R˪@�n7�;��04+c��� .*�w�2\���:�#Ǔ��bpȃ���֧��0���(��E_�qI5�bF(�@����D��fo�fD�����N@.��L {����,;��ß������*`.ҡ�	��PD�(qC���}�֦���0�;��Uݡ��.\�5�q%�7���ǻî��u]�29������$A[ҽWm�m��H��� ��rP�h��pgV�ڱ$���@��h$M%8�E��T�T��G*�?���S70ڮ����	mu������[V�����<��6$������ڛ�^�ֶ�D�� f%"�i Y����ύ���˄����/f�^�H>��B œ�B�J3��/��i{樫p�7/�:[-:� p�a�i��Pթ&Kh�������eB�� �o�m>���&̩݉�A��"=U\����?��QL���!���0l�\"� }<�L�v��Ov��U�?t~�$7u���h0�����#�:.��wv<��ꁷ*(����mr�m����_mZ�n\Z���0`��1%!
?��G��#:I��q|�QP�-�QՓ~Z��%�D� a᪹�������n]ױi͆ʶޝn[�����&=q��@�Nk&�Ɍ�o�V�P���_�"�
�r�kr֯�'"@NUj�Hp�F��e��O*�i&
{YC��g�C�a�V
�_F��g�	���zD�"$H�?q1#@��8��%��A�>�Z���G��芳�*�� ��|"5(e�t�Z�mGƍ��t�bb�n�l3	��(��-��J�mn��m��n �cU�B�l�   �_wlmכ�u�`6�Ta� 
�� ;�� �U*��UT�G��wVSl;��3��|���t�m�m.�mU��UJ��w��Ii"������j������
#�0G�au�\�3Tu���Q�Pa����u�s���7��.��z���3X~�[���}�xr��)=�,5�u��d��B���+	��@v�y1q[0'�>�H�i��F�k�]ot`)���d��� Y����]�ZH�O�#t��T�p��o�\���^h��*4���D�L��C�m}�l����U��GӅG�K���
s �"�(���h[(��jb7O�0w�f/�A �CPH�Q)(,�A��N+���nP�V,cD��:LwL�>aEi�b4D%�>�R���f��B$Ae�����>���d� �`�x~�F���n|�	$\W�����q<�"d�v/���7_kW�~�Gќa
'�R蟣���#��7��李��N�D�b��n�{N:���=n6��L�Rm�[lµ�d�gZ��m�6����T����0��G������g�F4E������N�9Ҿ��k�*�s]"uͨ��Nǘ���1ä�銸{J��W��[�G`�5/��(]~�=�2��t��拕��7�Ms��:�޻ϟ�~����<��V�λt �׃�@6�8���϶�y�.���j���{��]ݽ�֮8佋�/^�=�Q-������̭1���9��p�Ls^w��Υ��R�ݻ���^������� ����עl��o�(G�<>�?7n0�h���:qq~��o�ar���E�����[��Z	$��8&�G�Ӥ����^X� ��ͧ�*dÊ�0p�\�Gx?��z�1۾8e��#�$�8J�I:�1�ZgrA�`$�P $��� K0�(������Z<B4��.�8a���w��l��Zt������eu����+����# ��I2K!;��L`�J"����E@�T����6����	��}��c����
���w�5�����f���׽���(�$�H�%���iJ��@*�۳����t�����@�H�ko��l��HA8�T�d�I�q1&��B�;O�&��q�Dv..=��☎�i>v���41SH0X�`-�U[GrP����{\���m�fơ�_(&�[��A����$sG-�T �/F&�2�}W�G$S��9b���b<c���W��:�m��C����e@ۿ,���ф���)��1@bq�X���PߢDY�cd!p��ts���#�ES������U���x�Z)Z�*~��-Uv�)P���%�<�PZ~����m��0���s�N��P�A���w���"�ުs�b��XW�8�&���ڳs��Z���\�D�Y�{�U���z�Bi�׿��(̈́�3���miй��ݼY��|ľÿ�����U�>�eb��{,=X�~[��S��ݮUնa�z�`�j�+"����IƺqJ6EE�P��Y��'\S��F�m6�щY4�0Sv�����
� kśw��]q��lś���z���x�{��RnN	7Xl���������������� 0[=<� z�>�o/[���� �     '��� ��T  .�OP    �۷ ��0 A��՛ۥ��{yo�su����;���O^�z��ݽoe�kv�u�����}f��m�6�����N�/v�^�Ȧ�&��w��֫��;_t�9�zܹz�"8٪�������)�vNy:�G������q��i�w%�;+xٱ����F���{Ӷ���=���Q���o{�m��\q���cz�y��ᗞ���b�������w���w[o���]Q޽��oq�m���[tM���ۻ���s�u�{۶��{sZzN�/7�q�ezUl�۹��W��wy����x����Zv��ۯ9�ݧ�����k_v�.{��:ͽu��읧c�;�z��[��ݢ��^��Խ��u��f̭gWOq��ow��R��֜�ն�/4�X�v�ӫ��Ŧ��Mޗq�3����ݽ��r���M��.�{����n�ܖ�w3��9��s�&��B�\Fi��|3Y�[���|b��(�&KI@b�n��g��=Ј��El��AN �%��A�����k��:���4O��I��Lp@f�g\|dx:*���i9��wX�T��ܟLk�c��R��I����+����_P��N�}�x�Dv=7�.�3I�+P�,,��=C�<�����-(�z�a�鰻�$Ym�)��'�ڀ;�feַ%m�Q��0~�~x�� 5;�a��dmk�>��
*̋�4��bzמBhxl>D�V��ly-�@�p.N�Wt�w�E�L$�iXW�}�,�oG����u| �^��E���
�;�7ܩ"�#�>�4x�sZ	N�"�����ж�5Ћ&��q<�	��n��.@1���'��$`)��d�'e􊯄O��͛h��mc%�t��l;ѡ���	��!�B Vɿ�F� 6�J���fLS;�����W�a|I�C"� �P�W��Y��k8֘�[uPW'�ԢC�}/�5H����]��G��O��a\��=N@h�sOTL[ʛ�/��r��3:�I�O��7zֳzH�)_�8L�m��d�� ��bQYUp|���@㵲�������ȗú4�E=���p��eԚ���r� %m��l��;��UV�"�0�D��c��$P�vA��j�Nи�������et�MuO�]�NZ���y_G[��Kj�\o��5��h�Q��h�@&�H1T8��&�_p�n��QGWΛj�H.l+9�y`�0B3;��kf���)��g�aNŎ�S��dRB�E��ĝ�bR�&;�D�ĻȎ�bO��ܱ�Ā�TO!^*  �[]zצ��;���ȓ��Z6�bdZ-���G����ڴ�hB (0q�4��jD$�(Æ�=��x�DY<`�3F���sP��Q�p��:���H�Q��^��ʏoL�^P��	pIu���
�QI$�J[��1ڐ���O�ƍIΪ��E\/jD@�:%R���j?a?"�}� ���&E���~�o2<"��;F�O�0��P[��t	hk��o>7*�$����m�6�w�u����{{� E�T]ש���z�+u�*�   Ow��������w[z��m�l;�@+���*���   � �B��*�j�U�ӷ3�ݕ�Tخ�6m+�U젪U{���t[v?����
�����`�����Df�@)p��t���u#��ރğ��/���L�7a���08���m]��)�%�I��X�j�.�S]��e,�s3���C���*��@w*UB(���X�X�7���Y��)�����t<Gr竕�@��I О���璬�2�@�j$w �i{�<�j���ˑ��ᠲ-gm���߲���B7���t��$�I$�u|XCW�d"2!"��K�uq�y���w��?>�I�v wR\�,(�i�������ޑ%G5~���Z�O4��(�35#Qbq��E�.�����K��jf�7���T|g{c	������t"�g��Z�7�O��q1��,\���o� X�I6 I�����Z�b�2�$�e�,z|A1�EZ93q#�s��8�4x/U�q������/2��bF1�=.���h����HO���Eik�v��`�$�Nb��_,V��7	q��ʾ�n��(鹠J�A�΄�s]���Wd�-�I$�&It�n��GuPP<p�k�N{���l��[���n�����ޮ��립��vF��-�^��n.��qݿm���귞�k3r�|^�-����_��C(0`�b���B����s��jmL�&�;�K��{׍
w��`r5b�0N$��mɥ���3�i���6�X�]6�j��⯎�lh�/�ߠ2]���`����%>h|��`+��K�烩�v��ˢ@C�4�a�s�:�n/r���(����;�U�3������+�oŮ���k�6,Uwh���nfAZ(�o�|�lW`3����T�ۏ�WB�S�韽O=~�Az�.	�yS��4�o��˝r�m�&�m��� w Um!&�i�[K>ݹy��Nv����'䭌s��uW�5rw"�����\I(��!�z�Y )m�!�;�8G�YT'T���٤��᪽�J_N�i�vw�p��2/�:6
87��3���5ɈV ������^��u��/tO����R������>�'��j���y�ʬۍb�Xw�b�}�	�_���Sټ�ĵ"��t�s�pif�m�����|��KƮ�w��u�q�)M	��p6Y�{�Ʈ�f�Sd��n�y3+XX>3�M�<�m���E�(�]��3�D�I$L���>��Pr�УΎ�9��┾Us5�x�#�d+0t�R���F���C(����s�����q�M��]����P�$�E6�I���@%6��*���}�47ۖ.}�^��J�>(�-��^\u����*� ��u[_���6	̖[m$�I"�֑���򁺽x� á���3;�bғ.	�\^�Z�۱��|w�	w����.L��q�)�u~��)�IH�$_A�\�G8������q��+��a< �"է4"�zN�(ۓ�6�q%'�q�\��㩼nRd��@����Ȉ�t��}�� Wwm^��}��w��ns�y7q̓��dS��
/T-Q���$���g�yE��Z�Z��a�SV��4�E�k��܌z�V�=Ѯl�e{�Sw ���7T�<3Ͷ�I���-��\�&�����n������V6�����5�bY�2~h�Wv�O��j��@w3���ۋ��Ut��C�{wd �[h��I!4�i`1�g�j<��j����*5��r�f��Q���Qk�F�ޓ8���<V�E����.N���EL'��m��ؐb��q�K�N�j�kP�Sg� 7��Iw(��� ��wC*f��-	'A��V�$�ecZ�U Aij��<�MA��e�\�p�J��Z���ok�]�E��6��У�Gk�Y1����-ʾ<,{{ĥ!����w�3�xH9 ��!���(�(:`6X��L��Nw;>b�ムhj���*+qEi�K�tg�A0d#^�/}��Bqf�C(:�'�Ĵ�vt�JH�\�1c���<0�~u� �k]#��A��Zao!f�[�|��_u|}��B�&�n)dZ�Xz���O+�����g��u���NU{��������;����Y�?~���m�s j�Ub�UP   k�z^��箺��wdCl  d� 
�w�� �   ��N-���ڻv�m�jֺ���j홲تU7v�u�t��̿߉ܿ: o��J}��k��s��r�Z�L�0 �x��^����谞X�	lz��+W�Ƈ3('G�j(���f�69^o@CY����F����J6 �Uu?j�E� gb��F�����E� $�����׸����*��(��9XOG��-���6}ej��2�
හ؊�]��a�ښ�{�ր6"c�Gu��OB�)^y�?�`�4i m�"x{cQ�rt^�&�W{w]��kqo;z�j��<����ٺRrM�_8�{�9k���\o�ޘ%Q}�I�����+8+nv�4���i
�LH:V_�"�M$�M� @���.�v�.0S'	>����o�ce!���Hjя1v�	Q��aR�b��6�L�B&R��i�6�`�v�wb�^��ݷ}��%6�/MgJ��� F���Zآ��"������?�����S�Ub�F߆F�-�7�o�V*(4�H�T��=�a@�vm�&yV�A�D����n��L�$!
�^[�&h�����	$\���m��o�������O;w���c4��g.��5����{���{���O]��������;k魻�<�w��w���޷�-�l���>�n��ݞwy�a�	B�;�|${�
�Y��.���M��d��<�撂y���eN����Y2�%$]���V�(��@d�zɏ%�����Q4F�K-.χB�*M��l�gPms��5�b&b۲�"�m���ouV،��1wvk��q�z�mZ���:n�oQ���3�����n�hy���A���i��q�( 6+[a��R�x:M;�⦕Ͱ��M$�hW��,'�Wr�����\�t��A�� ��u�0#G*�٫,��m����!��,�]T�-e�HЀ%c`6L��{�u@mm�̻��$�@$�m��AYQ�t�����[��~�	]y��#QG�M�)�2(�y#K7����yd�Z�������)��l���F�"Y���-H���ê䙼0�<�Q���l�c�ܠ���Iוx�Ӆ#�p��ډ^���8d	�H�U��t&�/t~��WV��N�����(��r�'��������afmz��Bb��|��tBn����\�i�{�A���k��[[wKKi$�WG����l��%a"%�St]��{7�ד^�/{������q�C{�/��g��KLP���s^v�f�&-O�������5e� ��Mg�!��\_��S5��ŋ�x����>Ǣ8hǧ�$3�����\<��$�<a�����A��ES%��0X<��[�]w[�{\髭���4��\���,�}�;HC�~K$J��Z��:��6�Fi���������ǆS�J��A�I0���3��&��9+��~��DŠ%�f]��ŋ��ק<�����O
�{Z���M�+��Ֆ/�W	8yri�Yk��3�&m��
'J�x�ku`N������q����Zc��9��)�@�E����e�m�fxh�Z�4r�p��'��u۶-eݭ��a%Q{�RN3*'��ۢw�����ƮEAޙ�/�<J�R�Rґ��~���r�k�Ͷ�q����� �oWW�L�~�B�wVR1��
:-�k�wfF��wvn��d�j�w��Udb�Re���g<b�j�M$�T�d���\-�� Vm����uh�!E�р칳�#r�s0a]���,W�# ���n�Ҵ��%�=wo��+�-x��މ�����mv3ԉ���Җ��e�m�\��6�mn�cr3u�U���Q��ů
:�.��}y�|���ex$�AV�
'`��TSܭ7��zx.��}R�wt�����ּ��כsOr�J�F�����>�<�kg!��=�!��{��e:f[w�c&�%�31����j��o�{G���np�xeϭ�籧��F�����������X B@�!B o���������;��O^�KB���bI'�U�� {��|�$&�	�H	 	8@ �P��		�P �I!	!��	h��?�߆��˯��H@� ���=������?_���o��������������G���'����>��$ ���_��� H@���� B@?��	���„ғ����~���� ! ������������������Y��G�~��������$P		 @D    !$ �� �?�����?�I $ Y~G���=����g�?/�z'��O�����~� ��_�ݿ�����?a�~���������{��߮�  z�؇���������� ~� ���R2B� ��X~���	 =_�&+_EJ��_��y?#��1�= H ������ H��p���|�^�����a�O�w���/� B@�������� ! ?��~�������O�����������}�o����ԟ�ߐ{>����g��{ H����O��?"|Oǣ����y�������ϡ H@������w��R$ ~Ͽ�XI����(+$�k)�M��$� �������5���  �         ��(�P       �� Ҩ
  �                       {��M
O8��Jf��Q9IR��R��j��9Ya*��d*��D�Z��wn9�q�w)  ���   �_A@zS�ΥUL��!�R��9ՙ�J&�J�T�kR�&LH� �M2R�������H�Ph��8։US�����	��*�Ƥ����(�Lڕ"٥J�6*%M4�����H P     ��FXP��T*VYR9�wfJ��2��2��F�$֠q�s��T��$�B���@ ��8	 &@42 �� 3�t 2 ��Q� h���@  p�    8�: :2 ���s�p(��� 4�D(	h9�p�  ѣ@����4Х���@�4�@$d��c�� Г@�� vr�@����   � �    b��� H�2 h�p���А� v �� �S�P�  h � e�@ �ɠ ɐU� �a��P �� P��   1 #� w��6��@ � 8    (��@��C s�pv`h
24 ��ҩ@i�� k�tdJ� ���J�Z��   �!1R���d 2i�S����)�    `)!&��zLSi��?T�mM=@4m5?SԅU?�ڪ�I)&  �L�` 5<�F�C4     =��&(�   4�@ ^8�,Y2�Ej"lX��
ES�mIR�k���N[�W*�W�k�P�D�G�R�ze~hĊ��3_��f,&��`afVbҥ5��VT���2�T-���.�^[z[v,�\�R��z|�c���c��7:��{kی����^����JR�  ���M3R��Z0T�����+	M�Uc�ވL[�����@�c$�A)1�ŠD�X9vn�8�]�Т�2�f9��V�͕�����(&�V�����+`��H��ҳ-n��̺���xr���8��4��F;z���v�n�%f��W�n��YmԺ�K�m��f
���]Sw�6���.�3qAoF�3r=8�m��h���f���q�{�J�KJ�+Y9��pR٤��[��	5�b�2�X��MVLҶ�`WW���ۗwXԙc�. �!V�5حŬ�t���yY��a��GYgMkJ�A"i^��[�f��VK�Yd��X��t��Ԩ�0�n�%�el+i�i�W����2�</a�!YVDX0��TQ��h��K����T��*(�1�j�1R�a�v�-�hm�L�Z@�sf-/>VF�z��m�����Zgd�Bw�Z�����-:�Z���u�%k�b5�j�52�����d����J�?U^��U$k��(����}d�a/��p���(Ua��n���_RL1�GZ:V)%�1; ��;OXuIZb�>_V+�����ꯖ����g�s���پYܬF�Y�MC	Oe.m��`�n��s�y[@����Œ��ä��P��j�W� ���7Nb��^�e��_UUP}�Q�wL S�+�=�ô)ɶ1W9'��Q�5��V�a�)�Y�U(3]���i����q��ݔ�`�3n��*�9*��o"�m��V8��:q�@�Q�Xǹ��ܽ�;���e@��t�q��EZ-ѦÓq�1�Gf6Ĭ4�;ۭyjf�V�7pD�ƕ�j%ya�m��y0�v�A,��f��F�f����;�,�:z�L˲�6�z��S
�v/E��]P���0Y��n�ɓ*Zy+p�յ�X�dl)e�7V��Dn���y�*�nT�^�S��/ﬦ��`R�m}Z��eќ����mc�g.ލ	e�)�1>�w��J��{�!�&h�wyu6�@��۩r�31Tg6�D7V���ւ��෢J�;3kF����u�eɛ��wK2����(���un��f̋���Tn')�
�n�2kn=��ܛ�(aW�EcstT:����X�� v6�+j�8T{�0��[�]�{xJ����V�o/K�Y/���3E62�U����;�6c;D�Q�>GT�ma�^m��i�3K)��Suf�QO���mܹeTӛw�ɽY�mڠ����E5P^޴�4�ǔqꔳC�6�:��{�/(��{��5j��C�Y�yXVRxS�Mժ�oN��#yx�����;�h�Dw����k�z
x5mmռ�aIK�e;$@��`W�"�wi�vYMRt���7�Ӷ������`���J�2�ɍ�2�IK\��Wt��.�U��pf�͘�֮ٙY��-��r6𻡱�u:��������}�I}���ua��y��dԫ�2����)?�ު�:�Hx�YVk0f�)�1$�;7�/Zc>�*�<x�k�%jf ���أ�rۓZ6��4$p����EY��/�i[�����!��H�O�7���f��O� t�Bh��������^�w��] F��yBjBX�o/Fֵ�*�Ȱ�ibʎKd�G�<���"q�⹌��ͺ�v�Ŕr�N�L��V��.��VRP��n����+Va�|~WdiP��y[t�1˝_j5N���R�.4Ɨت��� U�`���
�Ѳ�Iv�k�ROi�M�%X5�����wsk��X��L�ͬ2���ɓN1ub����oJ֍kٻK/"F��8�MX]�b7�XZ)��W�j��`�)#����ڶ�/�F,`�^���3n�q�'[#���f^؊=YG&FV�Rì�O5Q,�6.X�Z0�` -ЀtE����;p\��Ux2e�"�իg��$�L�w0��聆b��m�g1��`�X5����h�1�w	̥�+{@��T,�2
zuR�y �S�w\�5b�;a��h�$��.���&f��aZ.%N��ݲ�������J�;W3+ػ��iu��z�	��1�2,�H5U�1/���"��2����lU�kp��U�P4ح�T��f�^fé+���8�E��Z�-qL��
��V��V��� ��Z&�Y�3AZ�r��@N�J��ca-T��<4��lZ-�w�У�^c��2�cŸ�ͣ��%}�7�X)hP�C�N�K���omv�(�R[`M�h�H���l*�j�i��{�P���ǂ��u{��m3X�v��W�r�pY'qLT��1ْ��l6��f�pޙ��Xӻr�9��;�)fQ�YQXu����Yah2�v�@�������vW�tiI���@L͢���sdB� r�(ԓ1S�oL�|3FL�D��^��d��F�y�@(J6�M���8v��r�]��sS��2:���C��2��۶"�ҬK&Yw�b��셤���m)Y���̧5}���/u�7r�2��+0�nl��j�M����tn\7�`R��ff�d��_�W�:O*d ��.֫�QR� ���uu
�4Y����g�p�b݋Pݷf={Oq����޺[YugO}�~\z��������uB����^������t.���F�,;�I\��]�#��W�*�.E�2�Vu=UT�vlZ;Q�����0̎L��.��r����F���@()@P\z�zn&��1����u7Ⓓ:�K�;7s�����~1U��R��^/e�E�2Ib�ٹf���p�ӷ��˝Yn�ybV��ТM�y(���ŷN�Z�.���	c�n���4b'b�������ni{yW�U�Tj���A�^k�]�$�DA풶f���@6����r-K�e��$��3r%=�b{"�N�9�-�l�}p�+幢N��B�p�ҕsfR�U.�����ŏ�U�o
|(�$wL�烽~��4��m��\/���v- ,ExAj��K����}1�=�L,;Y�ƌ�yMX������[�G��5<F���/E^9���m�F��L��=ǳej�LȢ$Ů����j�A�#\tϱT_j���F�۔E����.�9y���oF�ʺoh�r]�ܬY��	��\�fє|XDY�4\X�]�L�8U*���ZnYw�w0(F�f�f�F�b�MK֭�7��9!�M�ܪw��Rä	��, #DY>�`����m����(!�L4k�T�9Qh�eL]��R�̸.�10W�P��٪U{��Ê�oM���M�W�;��iI�5�MҰ��)�3VQ�Ol�AZ�Y]��e?�C�y�&�w��Zm����`���k�.D�T��7�
�O�J�l�
��.nȠ���Q�@?1t�
���̖}Ϻ�It�e���a4w-]n�/�ܑ����d�0���n�؂�1j����-�B��*�VP=�������6���UN9�VT��-��*f�IR�� ��lYu�os���X�]�ueI�V��
�S�ۨX'zs�WZ�WɊ��<yr��.�n��^<���G��MB�;�f+����+M�����Ô�դ�v��BI1�rn�����T]@�؆a����a��י��S�/Qx?�[!�l�
����[2���a�T�'b�u�-	��pS�L�͛��n+WySVM��X7P+�cB�/rc�١K.�^�3j̔�[V �D�;Go0醚��3�s��$?��ɮ�˽��\�I=Kwe㿍%-��6�]mF�.*[sr�
��)Q��[D,�Q�wR9VR�s=}V�P�}4b��EVX�}��4v���bnV-q�X�I��$-OC7uG��p��-
��+R��{B�o�A�r�-�R��"^�3K�]��>u1�I�fHU��M��t�
�cjxI-`4�ZW��7�x��E�{�.4��༦1I�&����:�݇��X��ݢ����v�mnG�L�;��24Z�F<�sES]+����uħۊA\�Z�	=�VP���@��o�6��U��PD��0,Xuaú�olx*��ШZ/\Z�E<Ε�[����i\���(;����jb��B��Ƿ�c�q��1�
�����F7dO �f,֢����
�by}����%=�I
1n����i%�,��f-{��+�ݺ�ݭ�YX[�G�s(��*�d��L�w&�u��Gk�3�'0��������r��	�v���d�Ұ�j�<�]k�N�Q�7Gw8��p�����]i7[��u�l|j*�����A=��X4�;W�:�䯫���?RG����mwJ���
c���^�� {*�����vv�7P��b�;��X�<c!��o/":�B�MQ��F���һ�I3�Qf��t���nL�)|-k�F=���[iW��P*[����Cd4ͽ Vܶ�F��%�7U�Ҷ/;���y�;1y�#K�m�I̦�;(9�QX�#���^K�t�j�N��d �\�r<�Թ��:�ƺ5�:���Rq��ģ�"l>��>�wS��tU{W}��	Y�x�r�+�i�؎:32����:���,���ꀭ����a_R�Ʊ�'6m���s�t�˖�q��n��kN�8��jq�2�몺s�+}�t髍rڭtќo���f���UY�̥�]:n�9m��m���fc��1�V͛)�����ëOw���<sz�N�鮰              P   *T�V�x 
����w2�� �@          P                        6�             �*� T�qUC�s�                        � @�� ���Mi��� r�*����m�     �W�U�UQ�T�f��^<�@m�w����ڽuZ��X)1�� ��                                    UR���9��V�#U P  �                  
�         *��R�l.ʥQUPJDK��� �Pm�   P                        m�N�e� m�      6ͷp 6��vh               U �  � p                             `{l�Ӥ��x{�nZvǶvNtԘ7]u�՛�u�v��p<Ͷ����$w�9��ώ\s˵\Q
�s��X�G	��::�:������uӝ�]�'([qe�{��s;`K�l�x��z{8Ò�hN��������1mBq��`�)�V�ۺ�	���mj�<i���7;պ�:��B&��m��l��w���6\&�cpK�%�㭷.�I��s�\F��i���ڴ�[�����Kֹ�z�i7cq�nxt7=k���.�S�����k4�V��v+�7n˺�u�6�oF��u[m��,J�Ll�vx��v{=kGob^��m�<�YS��-۞Ӳ 7�����n��krX���4��1Ń\�[�nk�u��ˁ�u#�p�]������]ӓ���tv�5�!��na�Fz۰n�$����;q��:�ѱn��8�v͹fxN�:����pȒ�lFxgf�R��6�Y�L���ю<s�=]���Gk���3�7�87e+��׶-�wg7L���s㷱��v�Y��y�<��]hBSIkq���H�'�j�xQ99.�u�-�bway�;�v�i��m��m�Nw��cW9Ƴ�rx��^Vh�+�����9l��շC��t����ˍ��;�<�-����p8�n�W��[�ctv0�����<�P�ɺk�c[$p����c��rŻ\&�n'���(�2`��nyA.y�<ط�7\[3tP;��-8�}W�!<��2v{F�P	���]طY��.��j�F��x���ݵ8J肄�f�n�<)�1��cqZ�(\��Ϯ'�1����NӧN�G"qnv�4l{B+��n�ۍp:���d!��|��j�#��k���<%�vzg�^��((�t�oF�x�[�˩�9����z���l�K���H]��d�J�D{�!܊r[�'�������l�>�b�L�tkM�z������5�f��m2��u�O��8��^��1�`��t�%�5��82u�ů�h;����K�]����Yk�22�{p��[`9a��q��lK��X��\���{ �<��Vzz�\�O����2Eۜ�@Mq��l���ݩ�МyxѺ�vۯ�V�r4㜖i��ِNn�g�t�i�g<(�7Xz0��t��z���v�]�MMk�ي-�z'��,��j�t�u�q1�G�g�ٻ���#�g;�v��9�ӧ�]<�d�ݵ�鱆����]!�g��&��͋���Z��	�Fqm��nԼ� �8h^�-�y۴]��%Y#����sv��!�q�q�K �˭�X��2�=� [0���y:8������[e��1�l������>�,m�muqƻe+y�ۍ'gU���q���i���u6&GF��[\�]�e���]:S�쐶��I`@q���v�%�IF6�\��i�ݶ�zA4 ���9볠���/%�,�����)�US�������>L��=W3�=u�5�pM�[�EF�;��#:{c�qN�])�q���môL[oq��ĝ�nɴ=Z��K����v����z3to�.��gv�����0�\����Q�;��]�;x␞L8��GlO4Y�u�oau��c�CD�ϙ�"�;�^ݜ�d b��y��vw\�/'<��i�=��wc�k��x�I����Bp�έ�!9��S�Ý�A�7�CJ�vݵ��l�ʛ���;��Rqm�a۷kXu݅e����嵌,����61ݔVvx�]+Ff;:ݞ�us\<D�^��}+�ã�]�^=����"�WGRܻqn3�&����\�G�s�6Wi�\J�rϧ0�v8&v.�Rz;z)��Rf֋fܜ�vK�:��.�(�.Kk��f�V����k����#�%f�ڵ�5�m����S�ۛs�=VE��	�\�B�m�2vnv�[��^ɓ�vm�s�fm�:,n�:vÈ�[b�$]�V/M�\K��<O6��c�E>�7��"��=�!��n9w$����v=���>G�kr[=[�k/�m��9�1Qх�O6ې![;��l6�d�l�;	��y�T5�@�	%����[�ͽf�^�n\���rƢ1v����;[�8�����!��f��K:��[g�]�Y
z˵�l��۷M/�v���Ŷܣ�吱�x���Lr>֣`�'&��{��ܾwNg�mڀq�v��H1��N5�7I��nA�u�)�cu��8tl�oQ��q�ĝ������-5�/
y�v��B3�^Щh<\㳓��ko�I�r����`�냵����`{v�	��z���l�n�R7c�7d9ݫg��n��u�YbM�^Rs(ݭ��[927m�4ˮ�]������s��U����y=�]��h�8R'mm`֦�cu���w �]r�F��n
�[n�`� ���z�շ�^�탛,e;bI��݁���V���l��&Q�ۊK@l��c�n�8z���܀e7S1�0�n
U[a�<R9㸼�;g�t��X��Lf��-�k>�������ej�v6Ko]�7[��8���͎�g�����vu��ۑ:���v�Ge�����%��ێ��M��[�K�Q#��6�P]B���t�&�g��S�Fs��]��v p7�Ooj�ݍ�hێݞ�ۮ��l�v��:5�ɛ�6��rK��M��8ա//E�^�6�cEv"�=���6-]t��x�6�e{s'[��݋�;��N�;,�h�'@��u	�=5v� �1��y2�1[e��i5��k��tg��B�{uspuƷ맳+��u>Q�4�axy��=���բˮW�B�1�9����;s�����]��pKt6�n2v6ݧa��#�!�+�D,�ё��v���6ǌu�p��ލ�N	횻�j��ne�@r�X;m��^h=�&�ƺ����3=����k��<���P��[9:�s�g�\�����G��{��ۮ�p����u�����nM��S�ƏS��7��arwq�iێz.�䭌���&�s˨���q���h7U8�U>m���IÚ�#vӭ���\r�<m����ҧ=e��c;t���`�7d�'�1ö�N�=��;wmS�VU��z;pɧѸ�G;�8W��7N@�Ȯ�n.��� ��%a&�%^��&DՂ[q��]QP�˖�D^ʻ��;v�������#���x��)E5M�R��Vg�[�����U'LQُم%/�JC2AY�)G1�0c����lϫ<��n�\8��� ?��cAQ�$����ʹ�������l,�����B�3���C<cr�i~koof��	�>f0���T���Spâ���v%�V4hrsn�\����M��~���jԫ�>Z�3s2��0����`�6�
����u =��0Q�vKK�����4gT��N�L��	�R(H�h�tP�.e!t��%2�i~�\�6�킝��a��	�TAn&��{�U&�ǆ��=*���p)��&&4��~JL��"<�EqV��LI�S&��(����#�b���t�N�a��F�票J
�~$�� � ,�1�#72)�~د��$�a6Rp��0Gv&����ܣ��Du.uh�1��XX[�[J���x�`���	�k�F��(W�4�m	�H�2�^�72vtE�ִ {ɇ�0�f�D��q�jfިC�vTjպ"�X���j4R����*�P�Z�cݘ���(�����V߬�mŰ �Pl�  UUiu�<u�� ;�c���rf�^=6�X��3���K�JgPY���~u���:���U�c�=���n�8d���7(tm#p�YS�0��zd�]��^�]����x�W�[>h�g'NU�]<�u�!�������u$�Tl<��4?f,F�i�oF������C*<|tA�nÌq�k�Ł��T#�tP���Z��5F�8�Zgg�5&��>�Ht(��� �0p���%14n��"Ѱ=$����J�I�ۂb�L-�f�E&벩k�scL8B-���G�11&�X�J&')[�b�C	x�
|@t
�A��y1����4�M3L�����j��67�\{�=``����s�^����怭/CO������c\�g�]g|;�&�,��~R#1z�W���,�&"�";M�3��U�xs�{�&a��
�- ��a�̤�Q���3�z�(��h?��3��[����Ї�}N����/^yEl���3�٢,|�޾��Y��L�N����71���^���f���W��։�CO��D9�Bk_x�	�����+/����9m��ݩs8�gU`ۜ��#�Y�/�u������T���A�a"�\��f��d2a���FY�OW�T$���������Gv�q��U��LjܸХ��n�v+�qs�:�K�U��=d8O���9`{-Q�@VV��ĝ��p2s�L�B�t!�ӹ�vd+��Y��d84���H\ܖx�`y�c����8lQwN�i�����t`p�7�W�s��c�9�h(l�`B�*��a���Α\Y2I�u��gk4uI�X�	�I��~X3�w�R�B�x��H{��yݘ'Rү��0SPK��J⅍�W���(�l@�}֩(��y`cP1���	�	���|��F���X��L�#���a8�j0|�D��l�!9:��Y�g2kj\Ra���H�AQ�B"P {��� =�xs}'���t4z�TA��X"���ݠ�^Z�:����j�P.
�U�|[��ӯ���[q�n$[��q
������������EN�u��e��/LTA�PK��v�^�QcDe8	̾�Z��/�Pzb\�6�V��@�H�M̖�Pޡm7WƮ�/J�0W��=��
W[��K��t%�!�˙�o1���ǀ:^Y��5�/f�*4�(M��&B�p9��:G���c��~41.vvX�L�bk���<�,��ΌG�P��y/Z�s=�7�CDft�^E޲�4i8d���>V�͈��t���fik0��7��1���<23@5��r�x^X h��Dgg.(��(I�LP�mJ�
�<���r�T�D�y�m�g&���%�az�y�0����v����E��kV���$��PBZ�}�Z� h#�,싟�������J�qe9�y�*4�qt�N���u�B��Pu1���Y.
�ǔbTC"�gt��{04Ȍ=�'<%V�p�����pۑzb�/<'��oQ��)��Wb6X87�*f{ޖ�F�,�s8|T4h[��{��~�\��	�Ȥ��4�
˺���l��p���t���
�{�����Ø/l�\�̯-���[`^���j纃�?�	Z�/,��vcA�Pэ-��S=�ם�8R�<.�Y�ZqR��W$�X�H�p
53Rl�F0}��H��h�"<�D�9�AS�1쓹1�g��d�o�����kewPM�i0�'Ӷ�m���qYh��W2BTP�>�[��aǑ8�Z����GƯ'%ԙ"q�q��X�0:�ƧzɴE2�
b`=P��:��m�e�=��~��@>�U�����y��퍧h�=8��N���};l����A�	���XLn�ؔ���v*P��v�I�:�a��f`+��F�#�-��@���ԍ��� \e%�@j�sN�����fR{g����j4�YXw�"êG=�X�#��tݮ�V >3�^Ŋ�{����hz���:�H�1�ʛ���@�}l��ʹtâ��xhe �� yn״���|� �X�8>2��Mt�ongMwp��(ӝCC�]c|/3��+���/�O��M$�m�v!{�GJ� 
�P 
���u펳y�G%���O��|���4��m���r��z��n�ݷi:�m+'Ue��-7����<t��Ʈ㳥�}�3��4�s�v�^w m��6�v;=�0�����=ة��V�@�
A�>)�,�Ϩ? |,T���^�ۡ���F���a�x0�)�X���S���?�O'VJ�nvX����|r��s���Ys/�@�^*AhW2\�cL/52����\�b�^ �H�T���Q5R�V;�d����`�����B%�;q��������dި��b3�q]�Sv�zK@P��]s��cg�X�6(О�7�"4�8g�a�Y�9R�.�&@��h���9wylh(Λ�Q��b��[�0Vf��k�'NX́#P)X(�뭭���*d�[	��* �<�����Ֆ@�&#ŀ��y���/�g~T�xQ��+��4���[��҉��!��.(LN�ҹٯ,lط����m�d�e���'q��?Q���6<cs}�G�VuTTf�D�u��e����_�;}Mr�Ҙj�e��L;�������J�m4�rn*1F�i�f��Ͱ�w2wU�\����K���ǤISb��h�V�w/p6h�)��~��v�XY=&m\�~�0~?1�U�B��=#<�g� �xM���6��s�����X˹8/َU��Z5�:��jyW�n.my�8yz�i�A&��X�^�?9+�ڵ���κ��M�b��*u�-h��=���e���'����g���%�	0w]i�����^T��ͨ3sw>+L���ƾ(,�ȶ{�h��h��[Wio�k|e�Se�k�:Po#���Yx�33n.�w�����v���k[YFSb<pߖ�9���)�0�h�+�E��VW��ò�W����2e��|<r��Ԯ�zd�؟yn�۹��+^��MFA�`�]1ƴh��H�l�ՙһn~���}`�K�Z�A�X�95�p�l�]�;�^C��e��{�ul2�x���k3��v9}�//\o�Vo{�K:<�������[�y�:�9V&V7��7���ŎIYt���[8VQ�ude�s�t{o���$"�[�~l�{�S��W��</7�
����G��[�����Y��u��8�>�h��5ގEK�p��}���̕���������z^���Y�Om��Z[vS��k[:Nd��SW����{2�;�� ��=��
^[M\-���~ ���V#��"\f�m�������l73�.�7v����{�=�/����?e�ݳ���s����%�{S��<��9���}��A��b�Md���y6����ƴ�nW���P0�m�؀ c,ca�^�f�h"�Vن�+�	20�n/c��5�Vx��ͅ^��d^���]Z��y}���՗7��	&�8^V��g��])ɡ]�"��4�;��J���gՂ��Ysa������I�7C,Z��v�������z�(�X��֜��C	^���Vb?3�Rc9�ai���-���dԧ�Q5�Q�-��9���3��h�31mщ�s�c�g�V�}������e�;��To�5�ݬ�2�"���rr���O%a\��f�G�35�}�����#���~��J�������V�w%�͏@�9���쬌��sq哃	q5v�z����{me��}�����~}�����cl�^��ߥw{�c��b���eڒ���y���K}�\V�֢wD��ٟ{-a�]ѫ����0��.lD��S`��������Nc�����|3�^�)ֺ�h�O]c�����$輵׽5BU:d�mo=���{�v����Gݲ})ޞx3�(D�f*�Nnş=����g�l��S�+���0�t�g+�{[�Wlf߶��ئ�r���3/ޭ!��9tt��ӽ�޻�,�;���X� ���\�I�b=�T� %��55O^��� m�^r�6� �� @U�� �8a���\���퇕�9KN�g��rcmnL���^U�X�y�n7N�䙆��;h��Ƭ�0p6)6�tv��qs�qθ�ld6.yJ�޻:^�����$#���U�������*��8�����R�gq���9���۳� l&	�����f��[��#=��{�w�Ū�_�cG��{���}�I��D��-��ڔ�n���1:����'N/�kc7=������ͼ� .�W�y5��d��ݗϫ���G͂ko==�u�W�	�-.Yz��*�y�����tz�Z����*
&�t�jK�W�ܮ��|]���__��=35-]X�'Ïnr����%(�L��J��[ Ů�~�ߤ������ܿ,����-Jcʂ�I�Fn헦'2iL�{h0�M(0���܃9������ףe��>8�s��oxa}ovob���u5��v���2Kj=>FB�cgD��өf��I�r��^�SaE�X\A��B�s�<}|~��1����<�x��}�������G=1�z�i��h=����-ռ�O]u��1s��t݋vf�ע:�č��G@*��tSSv��NU֌��96�ϮK���[�R��r�ڑQ�Cp�dQK�p�
��{���h�Ql��y���i�$
��K�u���]��w*����_I��+:�Q�T�n������ua`xh� n�*���x����P�;Ji
���/�;�+]�\��[7������G��iw�q�mf��t��O�8��y����fz]��0e=� ��/3��K���{�so.\��,�;4�83�,/���8e�e�1:M��s4�j|7kT6#�wTՄ3��]]�E	��nbl�$?R$800�!	�n�]C@�)oR9�u�e��h��˰���*{˦��e�mf����W���v#a�b�w,�2�wS��K�4Dx�u��{K��l;bU����������������g��o}��~��   ��:�      P P.��    �齛� y[k���m��w�v�      `�P      �l�P�@    ���l�@  U
�     ��n��v���w4����SqǍ�+/=�ڃ��|b3��[���p��;�)�Z]�s����vp�� �v7<n�t��h�絳�W��ə+��:r���C��!_]�tvn�z�r7r�1nxzm�`λgr(�9�\���ш+/\��:�,n�vî�\��9zS+���4G�l�����g�urn9*�'i�s��Z�]�5v��l��ѱ�j�x�1��Fw1^�wh�6�`������(H'#��Bz�a�C�Nc:�sb�w<U���e�]�qێ����+�vЍz�ut��5M�:�.���+�1���1�=N��uni㔛�M�k@'y�=�n.�����ز��S�uy�i�*i*��yJλ8ûc�j�C�9˸FB�ƴ�O��\v�g7g��5�������ͭ�v�!����l��6���w�q����Fg=N�ɸ�q���OX�#���a9���j:��u��,�x��n�U���p��çrL`��r=���氼l��.ޚ8�bv��v .cn.��Ό2���GuC;��(A��rv[�9��u�n���v�����5� �❵N�f�d'a�l5Z<�T��s�:�I�m;q�>�B�g3�rv�UkQۯW9�]t�A���%��&+�����G~?G��A���9}#��>B#�>">�#�1b!"?�~���>��ӏ�����i���2�>b�#DF��G�^Q���<q�F����>���0$��٪yr�(���Kd�� B@�j��&/�M�x3�hCM����$}�^�L|D|l��#�>�F�.�9c�~}7��v���]���1�f��q�G��Ä}!x�����t�#ﵼCxE�����Cd(n*�!��Dܦ>����D`��9.#�J�L��}��>�����������ؾ�DD�>����P��_��t-�샮�|;E��r���lN�u�b�Ͽ-�Ͼ�v1x}�c�"#����q���ĘN��b �������}��k���;X��B#�} C�A���v����� �>�#� �cP��,C�"4}��Ss}_@q$}B,}����G�X�l�ξ��Q����N"|b#G��>�� c�}묹�$}����8���!���>#�W���ö���W�>��Ղ�oW�eUw��<��f;MS�®&�\�Rl�1EM=+f�s`�l2�a�	4qP�Y�u�������}��=�|�t|���3پ�p}9cN)mnEF�2�=�s�U�ּ"b�L��?~w�|w����jE6N�w�ݞg���u�s��5�%U�[��@f2Ǳ{�N�r�z�dg�=[�Szb�;Ӣ(��}]W�O�]8Ăӝ3c�Z�B�,P��f�9�`��
��'C��%w��:aS��� T�5��nOvJ��K�©H<h�%���sz���I�����Eu&d�
r��{'-�$�O��Bn�쩧w��-���]Z��]u���<6�<��DLj��^�ա6�l�go�xY�����{}�c�:����W����]��򝃵y%��>��\�!&Ǧ��y剺J�ꡜ]����o��]_���C��R���fv�rpV������`�Y����Y�yӘV��ĳ�>��A�ʳ^ا�p$k�s�v�;㊎������?t�i��YkwR�W	��+�YF�^̃O�n,���+��H�t*^.>��T��{i������Qس%�}0�ʳx���#�͊;����s�'��ЊL�[FuK�������~@|�O?�<���Ʌ;e��\�ͮ��rs����λ޻�$�(5�����w�~��iY��S_탣����X��ѕ�����c+v����p���Q��:5�{ٞc���Ռg���\U�qۗ�q�C�����/�s_�s�Y��"=�[��^�S�Ku�߽�s��d�X;-mԭ���Bș����N�+�٩��>����Q.<��e�#{��M;�(��E��B-*�c����GY fӨ�Rr�,��F/��2I�ze��Sֺ�f�P�����VW�Y�5l��J��]>�֋���s���u��y�}y�|�����üT��{͌�a�ї2���4�Bl ]�S�)[�jai�`C�/f�=��H=]��=�no=������W�����I��:b�x�G�l?<�î�O��h��_A�}N�D?*�gt/�ܐЄ)���ߧ��o���_~�/�������υ��w��+[ڙ ^���� P x�������8;E	3��|��:ԋ�uՠ�W�8�[�m�Ѷ΂����<v��3�-ȧ��.3�O$�V�ѳ��t�vD<�
Pק��j�k�v��<��۵����z��gI���}��S0HG������ʣ6D�Gձ��vܕ*s|}��H��i�\��
�^���)j����O���3$Ϲ���=uA6F�Y����wl�ʁ^Ɛ�������i>��a�� ��=�������n|v��,�·�B�N���vvR�_��[���%t!�\�5�n5'lO�;7��t���y�{	�L��l���I�߯�ŝ|�%r������.`k���*�y�5�(���*���āYHRL��x����}�.�ۆk����Ph�����qtz�J��!y�w0�\)1�{y�Ke(KrƬ��(��RW�T=��:7]����潘
Y�w����u�����ĪO���mD��ܶd����Y8���ۊ��������<��<�w&1]{�՗-�y5�/Ns�R��1%s8��a��c	Ԭ�m�dˣ\����ʱ���U�֢�$<�/Ӫ��lf^���$��٭W�U[�*�F�b��rܒΆJE�M�~H��:�m�յv�qqq����je�=�<�1d#��m��7��#��{�IIU���Ϧ���
f�l��р���3a{g4����W;b��G�v\�'n��nW�l��P�$�v�󓛰L�<f//H�u��������!�r�����.>3Z����������Ht�)$�4���۽���㵶'#B��
��s�N�n]�.R���ɥR{<��̖�d�O�D�'����ڑYcg�3|��2_�K��q�C֙�^%m�����N!�h��QBK�ɍ���{��r���U��%��Wհ�랽p��ͮ:���!%��yy�P<ve�'�7L��{+3+m���c�����	P��3�.o�E�>�����޽��^mYN��E�ۖ]a|���5��U��)��I��zR@'���/K�Hy�T���l�Aj��Aa�0�y����٭�M���>��X�U��i�����n]�2W�U�:�fU���o���m�_��Dx{�9�<.���;=R���2��id��E��P�+an*�~��V�k��4ļ��f\�j-֯��Y:v�c�s7��`M3�{j�}.n�[��V��ǕfzR�ب�,m���(��C�vn���m����%���	�h����"��`�^5h�E��N�%�f�NR[y��CC0�p���p����ɌF ��δ�{͊�%*N�dte�3|	��++A���6��}��2��-_x�j��vE��0�9�B~��J�o�X���xkÆ>~'`Ȑ�t�7	��Fm\ɗr�,ln�����˝:i�;)���ޭ�`_ܡ�\�}���˅VLj��:�7���2����f'66ћ�9���z|2�q#cz��1^�)����J�wJuƟ�*y�S�����׽�+��������
u�Wz�k��R��&��i�Y�VM���[B�5}�墻�F�4k��o�)���j`�j:����m��OdL�`��p�1�f2jߜ�Wy!*�Y�����ҭN(��k�$u�1��ӼqZƺ�r�����ӛ3R����3���T&'O�2�=[ x��Y0EօꚊ��L82�r���ol`���o�5��60#����}������Y��t{}NVM�	�%�GG|Ӟ�d?�|�^�^̹�?�q�U��{Ui��=7Cwf���lx��� �p6a��չ�W�IZA+�hY�����ۢ�
�e�����1�:rXc�l���F��v���@]���.Ym1fՔ���}~|}=T �������� *� U)V�/&�<:HM��1������ֻ������۵�;p�w<3�;��Eۮ�1��.��Cr�ڰ	�;��hnD����ݳ�:��X�-n���a8�ɼ�(]���&6m����E�:�ka�B�d��&�7�㿬���:����I�D���rF�3_n׵���coAH�,�TyM��ns2D���κ�����������7���cVdj�b��̜+}���c���!3WXT�f�a^P���M���P��s��s����!�l��M��A�J����*������*������(3{N;j6�\m�R���5t���:St�t��cʟ?s��e�(|
�N���Egz���#�b�+kZq��({wT��֛���ŧ8�{S�3il_�׬Jݻ��D��Rϼcl
�n�p����EÙ����o�ʘ�N���[8�+��(�pK�h/N��\�� H�33�2������<�	�l5�����"ɽ4#fu���HLe�dk�����	��[x��l�i��S�cD��gq�DՍ�~O)���e]423��Y����iwv����j�-zVa�/UN۬Ys9lO�эO[́���)Ӣ�Wu���'{'����1~�up����UUUm��qq;��z�2땹[��9+<�/��ϽS�5C�zk6�x]���S;(��鹱r �.oM]�>L��2�)�jU�i�����mW������Kٺ)��f�_����^p�涟��/���~�
�o�{'�;�wb�X=Oޫ/��������T�C�g
��f�}�u1��e��i���^m�V��W�@����&ǰ�]-*���-cuq�%�������� 3fi�+@a"�:̳~�Y����@�����M�/,U}3��)��Y�ix�x������@��w�K]��y�K��{G���10'ھ���$f'3TmŝP��0��Ĭ��rc�n59�����`�J(��l'���ة��Sb��p��ی<��d{�gm����_����GAI1��c���b����~�2�v�%�pކ��0A�/�.�w,����y=t\f��	0@B��z��}ո9׎G��b�UႴ{�6|�}�ngt�Kޫ�(:b�g_��:;̦Qt]��~f�j[��b�ּ�$T���^y���I�b���G�*�~u�3�:n�Pu���ڜ:�x�ڠ�ӯV�bY�d�܃�w)����w���)����c�`�"el��"�㺎�06p\�<���n�E���S���w��"7�ݿ��.Nf���Ff�uyoU�t�����yu�<��c�~c�N#Ķ�
b/��o���~�X3g|���>��D��Un�oP���ۗNN�P�$`�P��@%��4���YVkO��յ9�ת�n@�1's��Mn����&s�Јe��p��J�i�m��T�@��^+5�?_t�W�Z��n�(;�����xF���VhF4�s�(P����ҟ�GD~gן���9�CA����n�w�<���%
�v�J�p�Gib�Z�L31�dS����KC�8I�Qq��V�kh�Wb��뗰��c�B��/����#��Ĳ�4�lp�a�K�8��:�)��Ե}��f�"�ƳCW�{26��c:������[i�vX��h�D�J�˛�Բ��^� �URȠ�/M�V�Q�˓���Y嫶a�,�gj2���Y�%LU�J��d^��m�
�ܑW.@��	a��'[I�p�46�	t9�1;Qto,�Y�[�쮭x����7�{KJ�x�ܭ2k؈��N�q�ǻ\�f;F�a��w]vh;+�v�{�{[Gv����9]���� f�wo��ڑ�qn���m:Z:̀�I:\̬;l���9x�o]:jc��1Gᠤ*G�K�U��S��}pbR�P���=Mc�Z
R��M*�E�_l�cv�/�j�x�eq���rʽ4̉��y%�|1a��p�K�٫�emXv9:�|%nd�F�VZ�Y:lߍwg3�{j��Բ��J���P��6��a�`�zf<�z��T���Q�^�v��2V��<�܄QpQiss$f߮m{}��f*��'뫝#�g�z?L4cJ3LS9S���n���ZsJd�
4��"K	��n	�P��1$��9z��&1��&�j3L��C�-ԧ�S���7�=6����87B!��Ue�S���R�LDJ�%$4�s �s��=��P!C�P�\��|N�-E�{ f�&B�ژ����{<�/;{�׷Q1�!�f�����(�����L@&s��"�}�+�ۡɈ�xg��˅o�5X���w�j���+F8����K�S09AѲj�u��v.%[[�l;�]��5:�	�Qo(F��k�./l{-�[I7[ ����q�1�̃Op���}9��'/ƇF�q�n��S'�s��ܵ��[y,��PZ�Wo4	WO7&�$V<�G�\�m��	6�ݼ@6�b �P��U�  �[�{v�����]��	7\XW�����Z�v4u���y:뇶��۴��U׶ɠ�$�=&�O	͞A��^��ُ^nNX���ɍ;O-��F�Y�u\<�w.�[����k<�R�h���t�(��V�Vl~��-�J�aO<�
��J}.��Vo=�z�؀w�m�}�Ĭ�s=����n��	y��}h��D��Y;��LK�*a�[?U���i��I���X����U��xt��M���g�i$�2�N.up�{b��[0�۶��E�I��Ib�n�.�O�P�8�;~�7����2��Y��Q�ݺrd�m��r0�e`�^r�u+7=���zު��eぐ�e)6t/`Dၚ���uIot���WQ+sۉ6�6�O��W���u"&��R�]7m��*��~���'��f��`�O��}q�^�r�+ך��iAa0������Fb��~����eګ�Q���]`ו��=�`̷��:rv��=!&��@mt���Ggjl�|_EZ���bm�ĳ2�N\:0�Q�h_=�S�	��k]�GK$��HbҞ�m^�Z&�E��󺨑�p�LM ��wj�Bp1�э�M�^�k	�km�P�M)����~|}�������7�vک��G�X�o�6�] ���=�s�EYlgI�z��Y��v#y,���Br��� �����Dl�a��(��!���r�����>�ӫp7|��p��7[�nS/m㭧�0��Lj# ��>��5 ���p�g�:��*5
�%��������d�ƣ��bz��>��G�e?*��}�8W�#��#a�&�ez=>�qk��� �>j��ڛ~�y�״.�ۚ�v��x�ߒǜ�y\��m�e�RD��,���lW�Bħk������<������i��o�{Ʀ��~��bd��w&�>�W���Q*�f+�����s{0�{s�VJ��2\�%ʁ �$����)�O=��"�.��۝	����Ad|C�d�攦Ǆ��Zss!��!{17��^���O�������90',S��va�����g�@��:4��*gֽ��L~������^�Qb 8p�/1�@����d�N-��8P� Pv��7냏�.RM�;;�j߾�'aLӧ�{�-e�h&���}D�M{ִ�6��L�U,��&o�%c#�F���m�wl)Y�>�$V��^��Xw!�2�,��L�FeD�w�q���A��5y]�ۥ��+�O��y��^W��J��㘭��8�!�\�тo��u��>�c�NN�i)n=/�J����_�f�vA�K7�;�}��Diᶶu���IY�[(W�h�=WIzwf��د�?�-��m���p��㲑�z�gc�ݠ����>R�`��?	���VД� AMaRlfj�`ULU�ө�a�M:uޫ��|��� �����7�Q;TF@��ٓF�n�����2�Ecڪ����V0l��9��yTGU�����a4�*�;���A�v)��kݯ�U���[]�㰰ٮx˾U�!5�Ώ> �瞷_yl��br��m��Eh�Y�T7r/�̊&�z6�٬"�IQ9[��,����� �����]��A',��=���tE{٭�|��й� hv[݇��q2�
l���}�֛�t�� d��݉Z��ݨS�Ӯ\�ۥt���Q�7&pI;��Q�٠�|4!7�FH��xm�ȯ�fL���+n�ƠI�iUc9�4���O�T�k��� I)��AŦ���� �f��6(zgA^�B�Nu�����;
��R�U��E�(�؉3�����g���i{}c��>���H������g<�Z��j7�<�fV�ʉ��1�w3��Ot7��a��G�5�=Й�v]lwڄ�������á��ҍ�Lۙ��j�n���6�m��t_�2�D�G3d�(˙�N���M�+٘,[���tˌ�x����.������{�mV�aV�v����s6����;�����x ��g镴�� U ����^N�8wgkră��Χh�g�^��r�Av�v�.e��B8王��ɻw$'������=���x�6��r'[����yk>iM�͵�qG�,,8���\pGWp�q�Ɔ�h;=v��]�����}>���L�#���J��}�0F��Mm�Q`&�	���^���ٛ�G6�������~|�N�ȱ��8���#��u]�13�J�R&���y��׫*�m�y��F�������O64ˋl�E��M$ID6ň�]�G`�釦���L�a�	��?�}���Sv�*�ᵱ~��m��ˋ%�W}�n��]�_n��E⩦��s�S�$��U�����Wg�p���o9�9��޸���O?F���wg��֩N׵p�O��
`��:�%�<��������V]��w���>��e�xg�����nN����_���\���ڽ��>�����3�D���e㟓�} %5`�Z��>�W���O�lP�j�1ν���乜�;�IM�ML¥�Mn�����՛�/�>�xI�;w�� Ownbm�u�ֽ���[�|+:v�_����-�ą�].O]��e�-'���ǽ2N�̋ܠ%5�ka�X+��(c7��3�g5�k���_�����n��}��^����Յ�#y��}[닇+���Ď5>�Y��-�7`B^�37i?F��ɯ�x�7�f�A�y��)׀���<�w��pCݗgn��wBe�i���S�!4�U�ܔY:���N��[fW��n�r��OW�X�z���Xu�a����wf6@QP�P��w]y��[��N�g����_z p���|f��l�J�w,`�6,{��S�Y�7O�>��P�j1����Y�����uV»�պ�h��7ve��V=�U㕷XE���nv����f�8e4ZA5�:##����/Q����+S	 j%�ݦ��졟j�ph'�y� " $�l�m�@��y���nb�[t��0�.�	$���� `jj�t镖%�P:�w�;KV��j��g.�L�� �D�ySQ9~U��H���U�2�u�Zl6�Lt`�eI��[�ƽ�^դ�d_T���!��;���~���f����7XXpSؽ0$�7��[/ u	��P%��W��'/E�ջ��y>�'o��w�{n�f��IZE��0`5��W7����n��2��+}�dh�������*w��'ҷ�ڭ�6�o��4F�Yh�˄r�i���ϳصɵ�d��z����Z&���+�+/��}z�>�D�G�[��Œ�f�T�N}p����T���ĕ�����~��nU	��t�]�[Ttb�����G��D���p��_�4����E�{w1�k�U���~���]<+%�\�n+�S��tS�2���4E�~�`Pp��������6�3��<e�K�{Nl��]u�}�w[����X�qd�y1�C:���jŸ�6����n�{�+�j�w�	4���r�`ߐI��=7��a��9�装�#;l��~5Z���J0��s"�;�N��Am�*�I⇔n�N�*�:��ث��V>��3'����6��NDm�>��GU�Z�r���ʂ�!V2�jwn��Ó�d�#Pe��w��Y�#��|[��+�Ϡ�\+v�U{Fn)E4a�\���"��M��ʷ� �I^&�-��m��&()��I�k�rS����u�c��!I a6�ǻ4z|���赛�}��z�9�1���ů_��VѶ��^�Pۆ[k����{�nj}�c��<u�����.�E�^���" ����3nR����m��&{;�V���	��ە{=����q�B1WP�y����m�}�>�χ��3���SׯR�姵�}������4_��R�/^,�A��CNT��ɸ���b�����Mu�bc2[{WWDZ���y��z�@ m3@k6�w4 U ;� U
Z�[�˵�'Dvݎ1ǫ��6��v�c\��.�1�.��sw��籒��(��A���9��r�]q���8�v���̶;8˞h�w;�;���.5�N����J9�����p�t%��I�wM4o.��������q�'8>q��9�5^^A�D�G�<Q�"Zj���6}8��ۏ"ݫ{4�^����0���7�M�R���`JKbU�úJp"[�P�m����C3m�1� =�e�I���m��� ����ѭ�h#G�<� l�&��n�T��_���m��<�Vn'�7L�2���O�xy2��)Ƌ*���mZ>�2��[S��{���̊���b�S���_V;=`�z����� ��k���]sB9� c5<�VU\�P�fJڱT�7ӫe��Gg£ga����R�To�d&E&���g�kH�u����f�^��p�ǣ{=��:�2M�u�����;��Hb-�;�yVV9q��;1��蟴Bǲ�0���۵Jy\�Ftu��g�O�e]J�Lt+Su�n1/�����!ܺ�Ա%�f�՚���gR��X'�^�_���kC��G\-�=%iv5������[�:��ذ��њpmȬZՄ#�׺L�u���m��z��)v'vm�<<��ۺˋ3�l�PNi]1��i�n�w˦<�^�s�3"�Lv�*�.�6���2��2�+�W.�ر���5���mΥ���.+��}F�6�����uu;�0��[�Yͦ;8��/�ӫk���^l��V�t�=TL
V	�bǯ/����ɺ�83��6&p`����Ê���0�Sy�v�]d��ۚ.��]_,R���U��ܕ,̝%�yGp�n�4�+���������T��]E�+ 6j�:��&]5E=F�kL�C�K7�.޽�,Rܽ��rѽ�W����\��v�*{`�v;338�w�nNx�f�e�-�8��Ks���0�\IT������P�S=Z���x���1W�+2����������|�w���   �M�l         �
�ײ    ���w9���e���鶷�^��s       6�xʥP  T  x�m�      � Q�   �     ܹ۽ζ�/��;��ݱ�X��G`9"�6{�f�ܽ��e�d����;v�R$����\��ع�Ha�����c�\�2����n^R�]PQ�J[n�t�޻Ls�slGus�����0%�נ��=�Jݧ�q���g63�y����h�9�]�	�>���-9��R^�kqF^{
�涸g�[�6�ח�ź܎�/]�e�r�[�#��״x;w7��:�ېwZ:�..���.5�:�x,׋���\�;ն�Q��V�ngrj�]v�I���[r#����M�/iqΜ=v�]�m-t�;��a㝽�\��y1Ύ��ST��ݗK�θ�KI�J�!���Av�lX�#`��z���^��sbx�WH̊v��a�b����1�:8�c=x�6��&�N�˞C[n�c�Ʈ��N�8�m�)���s�m�[�Ϋg�v�ѳ�\��r��=bM`-�I���/P/K�\�u�mq�;Så�h�G;F��<Ũ3Cc��\��z��{X1l���X=��t(�;��]��m֌��v-Żm��� �Mg����6-NW#�O(����a�wy�ut\.��
���g�E���m�ָHR0[c>��f�yܺٯ�P����g��]�dD�<mpe����T����nOg�Uĵ����B�F��}��A�q��Y`�R"L�U���g�X��q;�F����k�ֹ�[m������|�d,��'&��b-VeT1�6�� ��V���8(4C��/62V3W�[p�6vVz�2�*X�ڌea�^�z�
�O=hb�S}�m��c�%CI'���;a�gr��aі��	݅�6w%�{^ϥmM�h��k �^��[~�)��a$�ڮ�F�כ}��M���y�p�����}>�R�U[h���5!^,E����(�7O��e���m�6�'�_�f_�	kQͩ�
������wo*�쥂-ҍ��QW��('�myj>�ڸ��rn�cn��Ul���SO4��6�ֺ]����AʇP�ĔOg�f�������|v,�S:#��o��ju�r�G�wD>an�F%�,��d���R��f�`�k��0�uv��u_<��{�n�{����Fר Ho��V��Eu��A��~ޣكo�w��� ����Y��(ֽ��;��-�C���i�h4���aFZ�Z�W�y�����,�3�z���>��Y9�։M����#T�e��94���m��d���ڌZ��l�oVd�<�d���ղ��+�$�8���?-����Y����5�z���=1Cۓ�z��c�������ۈ{����gy� ����*�����K�d�%��ٿ/7ks3ƬGY9+��U���ֶxnA��,�um�s��A��n����D��JU�*����ec|n�V_���fS�y��V$MZ����I�`8�����/_r��]��]����{��#9o�ձ����9~��S�Q��ћE���I�bo�6�C*8���U�����4�����5��y�[�ث�����Ek/ޅ�Z�fִb{v|�L��]_�6�_<϶׻�ǁb� �?��籃M��4ֺ.�=��M$�I�Dd��6�w'A�����~O�h�e�Û��yM��ܤ=��5:��g]Rob�F0�8-�UJ�<@�l�*سW��o-nfj�[�)ac=kԚ|lis �ȯ�Bb��g���^�	CL�b3�5��d���x���|�o���UV�8�Ӹ8n��v3���a�us�7����;˸Ƭd_�%�I�,w��Hf%#�=w���f_��%t":M���V��vGE��]{����n��,��,Z����Ĵ��z�woN��}���E:?oUЯn�ۻ���nK�o�3=[ᗶ��͍��C6�W�f3]iQ��0'q[x��~�m�8M�+����Z�Tr��� <P���2�&enm\�[��+�9V�s�2��x���N�Eq�5q�6��L����?��ލ��@�oKyk��V� �� u7q*v�ts��O�4v��nfd3�i��gY:yٔ�d�R��k��K���nm���[v�Mp�k�3o'iz�%\���6pb�8ݶ��ء���u�bwg���A����\��pd��Ap �p���,M�8W���;L�)�ޕ<=܂e�I�y?zRS��^�ô����o�s9���M��E��*9 {�y�/*�Q>���,[+�v�v��8+F�j[��#:ʱz�<�=�|}���(4�-�H�D�aH�:q���V�k���F�TX4n�E1Q���+�����}��O^��3�.��J�Z�z����T6�Ç{�W^)F�R:Ƽ��ƚzw$Y3�bl��ov'�}/a�XZ>���sw�ŚLR,��=��e޷�;F__S4�Ϟ���s���OqX��H��^%�5��>������/"r�e��*�{�~�>����{�k������U=04�U����(k������R����#7����z��p�D<��n�2�����`XU8��P�s�����yF�7��Y#��Ǥn���N�d����Sh����)��TX��B�����Gar�.33JjeǞ�kη��^�V���&���H�-&�y:˺�o":R{��+� �����'���C���b�W;Z�)@��l�f�b���i{~�M��@�z�ERN�
�^�=�9J�J��}������ve�W�Z������T�	������u	����a��]>���@��u9�}v��=\+nWi"5V�	[�Ж��-إ^1�t��m� s�.�\��]>ػ���Яw��b�a�'�\��\	�>[C��^�)��4�.�����G��o��X���W���:e_�@�XQ}S�1��l�^TA��^�۴��� �6#"B`���z���s/Ⱥ��'|�$�I��m���k���m�m�M��<�q��.�Pm�u^�]�iukR�s6�ڨ�Jȓj��v0F��RMM*�ȅ��`F�.]d��	K��3-��1�����=w��^�@�e'7� D�V���=� ґ�26�^�;ʷRk�OZ�b�N?{�U���w�7�6�%8C}r�U�ަ�Z�n�f��eEڭP���y�*R�k�h����f<�b�]��&`�����$"cf�P�Q��ɈS{�9r��i�]�O9����3k�;s���+ٕ�u�j�p�L�H�.��$�.P_.���׊���^���@��ӵ~K͝�~�!�-b೙�����Y�N.��x��L&�e�F̻w�}{��'
�Yԓ�&%�:d�N�ҭR����M�W\z�s��(���81  �00 7~�Xީ,d��u����N�N��9P���q�`�E)��"�Z�Y��J�>���t��o�]J=����OF�v��K�h8�#FJ�u��k�H� ����9ۛ��&s}��GW%)���ewq����|B������s6�t����8R\@����Mus�����|\�ޥ�&]e�.γ����ַ���������N�N[��[[��];�	�-Ǻ�F�J87+c,o�Vkv�/5�(2�>��@X��E��CĮ�N9���O�^b=�]��C&�8�md��ߔ�M&C�ç}��Ǵ�m���%[z,Iv�I��I3���>k�y}���[X^��Ҭ8p#A?3�H�n��NWQ�����z�M�jE�o֔��p�����̀�Y�Ǯ�*}�l�͝8ƻ��v��[�nj�=�5md�}���cܩ�жh&�U���������e��p*>��)���˵oS�Ǻfs��_��B���f6�$68W�nq���+��B���X�^�=��	�%�ae����g��U�-W;�f��W���/�n�|}}|�ﯗ�p ��m�� *��T ��{��5�l�껞��>ۊl<������-gu���ES��9%���#'m���v5ě�D:M��u��������>�]q{r:f�v�u'c�<�ͷq۝���8��`N]�m�Q�i�GO0=q[.^�b}�����U;�K��Y�#0f�8l�3A{�ʭ׋^𭥢��&����y�;h���o��[���?�	�z0YE�]5�k�3���9+3gۆ�r`A�m�fh��r�C��q���^�v��T% $�e_��؟;�d�d/wXV-=OF�V�md(���¥���&�T�u�~�*��7���¬��7Lx�
�=z�r��2�b�g�=�7��vI��Fvn\�W��Eۋ���V��gD���w�ӯ=���s�:����>�3գ0���J��z*�m?<��o(T~Sy���1y�:��c��X}�Y����ޕ90�a6^Jz����/��U���w�Y�"���ӇN_�c;ט�mj��vq�v�ֳ���북��>�tu��9�shT�o.�#�tmɫrg5ez�Ǧ���ΙݞL�ͷAR�q����YW��R�O�a�P��=ł��bzw������'	�XH��$|�"cw3kʽ�2w�D��v��z{=�]ҧ����d�ql�H)��7�z�S'^?�cv���W�7F(�{�c�.t+��gB��
��-���R�~ۙ>��r���6׸J��hy���zY劓1oe_��-��<�i4�'EL�y��3Y'�ׯޒ���^��+9zw�6�_VL����-�E�K���j�\iC����u�=�N���f{ŝJ�6��ٚ6��V�Je�i�e'�NSM:5� ����;A�Y(R�薫���^�!]��tl�ۭ���0G"�῟_϶.5��y���̆�!�F��%���ƤD��-�6<g��b�1巓Z�|3A�\,˳�
K��gy,��V�
-�P�`�5�ٿFf� ��0St(��d��ȍ�{P�6�gU��;�=��W�]҆������mL����l@��$jE�ậs�V����&廭W���j���ox�C�_�_�{5�~ܥ>��

L��Ve*�Gc/M�K���"�ݑgư̭�{��5��r�wv��H�A-�D���	Y7����NU�<�<e�9��Q�{,"�kkU-o��yZ/ٺ��"۴�J@^���SQ�Y��̀�L��n�H����Ջa/i`瞂j�)R`$S$d�G*���^�͑�{Գ�����7��`���)\�e���אK<���*rh{�a�aH��ӭc�X�f�8���������r��c�"�z�k7@�:ӎ^�=��uӋ �6�� �Y�6j�g��	ݗ�eI)&���꒙j�E8�7bm�G��7�L�镧R�/��S �ק+VvueL�p"Q��.w]���a��/*�1��
(�Im^:�J�D��U��q���w�߭�u2Ԡ��X՜����f]u�i��6L�9ؘp���\VQ�NoVh�7�\��`��r�����wrƕMĵ�kw��/$�c�7�9fM��*U�f䴬�o���Î���	U���Anc�*���
��G;W);"��>��v���t��Vs������������B�,�Hƈ WO{����;,Q6[�:��,�,<F�ta|���7ix�짗b�G���+
H�]|&oT$�t�M��Z�"�4��[��c�}�@�Y�wr�t�Bu�	7].E�+��0��U�y��\����m.ZX{�i����j�V�*�]��X|�v�v�ٰ���"�%�Fl��8Q�>��o��f��_�Y�h��z�#:�Y[~�fm�Yդ�-�Rr-�4���E7^���5lBE�8���N]ghL����;=�zg(>��{N�Ȝ�,�Sa�гl�����m�;ފz�.|ߨf�{�ާʮҴ�л���l�ضg���h��U�[)��!F/Y+E_�3��c�Lfl>Q�Z��ۗ4��I�8�I�S2`�LB"�P%#��p:|9*��%=�����#�����>��3�}ܟ{7����	�ئ<�o3=.=J(r�ýStd�2�ldy�);�ه���wx���\���t�r����4��⏚^�8_a�n������2a���e���a��4e�R9�B��lay>��۝>	��TV�S�Ѻ�H2am�9���,��^��,`�������*ow�zL�[Wܱ��ڱ}���wu;��к��NcAc ��v��M��x�%M�D"�m��6��6ݧ�i W�T �*��;{��ި^	�X:ɮ^j'����:�x�xⱥ����j:��-ō	Ƈ07=C<��tv�&���8ݺv�$g�q�\�N8杲���5�L����^��j�]q���;�V�#N����ԇpv�Y��pp�B1��D�<ȡ$Y�+��>�N�ׯ(��q*O��<����!1 \Urt���\k6�y�Ӧ�ـ	�5��.K���3����=���a�v�t�ǒ��K"zP���{���Im����MU���j��6����տ�ś�ҭV�c�Ɖ�,�u�$�s�#�9�zb���کw�u��M���K�B���&n���¦�]����Ja�Q��j7-�X�����ֶ�'����}S@�#*�|�t���T��፣,�I�^.O��9�5"��Q/���Tݮ���T߉�"$S��_*L�|3��f��O<O�z��zϏ�c2�[���y��a���	�a�E�L�c7J���m6=Ul@�;D˕2Eo��vnP���4T��c`xJ+١Ξd('Om�=����&�PZ�N<�����e��c��҆"����.�S��S�>!�z	rf�q����oƁ{�f���(	p�Ҋ��̮�v.��:/&�Fc��W[���o)?ѧE��:�;/�X��RߊpJx��ؓ�u�َ�\@Ϫ{6]ȉ܀ ~¨���c6�84�=��g�=A��U��������u1+LPP �}.c�F����&n���l�oxv�U��7A�� �å��<cÀ�<��pr�ۮ	��1Z�3������~#�.q���Gڣ�v�H��><��w���h7���q��]{�S���;�Ixg_��4h��ӳ�{�'֭�'}��>�F��uk��aބ�`���Nd!�5ڳLoX��,���rR\�8�Ӂ]V�X����6m�Xb}�������5-�l�oj6S���-֭��^	΋<N�]@w�~Z=������|]y�U6<@[\��ֽµϥ��I���Wz��l�����\T�y����[����m$�	3%�r��:�2��ő~)��$[P�p�m�)zA���Q�#��-���t}�����U領;���߇1\�u����Sp�k?.K�s<���kX"�񱼃�a���?{\N�z3�i�JiɣbSΟ@��'�F��z&ꤓ����>S���NS����bW/d���jeщ��K�T����q�WI�e���mOW�u\dQ�k6��۝T�xu'e�1$6�*K��QlYFj�H��N�y�D�+�ޕy���h���(�44�g��uw"�I�>ǰ%��+�����w��=٫��2����sUUG�A�Š�G�����4��
A�����\\ד�.H����4�{w�.���m�$w�_����'uW��,P{3�^g����!��.�q�0��en�r+�i}\4R{����ժ���l>]�o��tg�6����Y�qR���῞�lX�)X�=�`pA<�ꭇ�:2Q�����3@m���i$J�S����p�f�.�xR� ��1�]�%�zE&ݏ��8�(�o�r7Z�PӄפZ��!�W>���I�69)��(Bf/*1
�o�L�{x 2����s��
�:-.��V���[�R(� l>Z=��$�c8���08���m�4.�_L��a�R.&|��14^�s�_���R	n�Q2{&���������_����=Q��.��H�(f�)��{Q݅�b	P�c�Rl�#��%r�&��g)��4�u�6<�j�i�T=�d�>���R�O�Β+�P�}�~3�vD��5�	��U�Bb��4�}�qsA?�z�'����Ś�K\�&���	P�M�R��H�#Wv�S�v�S�p��4��Ԝr�(h?���C��>]X�>&�ަ;�ڒ.p(t����}^��>s�ꐼ5�0
���j�{�N���vuˣ8i���]����s�ZI�\���p�5�FD��#����LZ;Z�NW�J�<#��{�����GWpw����%��v���H���܉���C%��L���`��0�h�ZUgf��d�z*`���a�Y�ț�M ���8�c��Y��}͌/�U�]���UEV�WFre\ۦPI�Q��u�ݯ/ �`� � �Z�m۱ۓ�������td�I<c��s�[GI#Ѷ��ȓ�M=�<Vx����k��J�c�v�v��r��V���vg5Ë��X������q����ݟOQ�T�S�������Xj5
[�'��/h�����v����
���1⧳x�Р�Z	��-����^�c2y\x����~��G�w���u�}�_���͌������O�=��s}�r�G��{	��%�X�gG:�s|
f8���mX3R-m��H0�&��1K��A-��5ٝ��nلP!�lffi���Y�K�;+�����Lo�:ث.�/���R�*�{�� �$�ِ*ՎRG������LJ>��{�6�G�3�\����р/���t�1�� iC�rk'4.ZiD'�C��tݕ6�}��|��ɓ�rV�O��:<;L^:������g�I����ޭ�q�lf�ax߰�u��FBmA`&$YD�{���r�͚ �]]@h��7{�8f�(�s�(�X�k��:gh�3�2��ykN_˅�#M݇k;�gh���Uȑ�[�'.�i��@3������5;�5O
��Գ��6Gny�蜩��34u\��!ֹN�6���~�?��̥����OKw��Z�@Bi�Q�8U�U)$�ٱ}��~�����p�V������c����x'�rv��n��I�Pl�ߞS~��q�gNd�u��"x	}1�=ƃ�QG&��������J@3��)#���.�>s\z�O��{'�4l:;�Cw`�y�y����t��C��-���nk��Rf��9�HZfzT�nLs/޹h*r}|�9BʘЄn��+'a�Pxky��;�,�ڨOjٝo+��JL���Ш!���Ԟ�1���5:�Q�`��#��Nd8��p>�6|�zT�8�O;�{ ^siSH;Bj��T\]r܃�v�Nq�1�6�k����+�X���7%�)g:8�<"��P�zşW��C�7{�u&�������[ip�N�B��o�ڂI%�m��m�N.K��+r��Z�ܳ&[I�D<E{����Gjޛ�"45v�;���
��4f��3@��:ی��J�S`�*�M�`�Q���u4J��V�\��_I��L��Id�&��k�������<�����e��"�{��^�.�@�xN�ݡ͝��x�`���#[ �I���L��~����h��8G�)�9^�3��UI������)J��6=��w��*��T2��y�@����ȵ 8E�y�}��y���'8��ne��r\سy^瞎�©���8$1���@Є`�	�l9C3r�IM�7C�sL���J�w'��������`���r�f
�t+g�K�;���B�w���v]O�9��PY���!=�!Am(I�nE�'���:Q0|/M�v���I�&�N�n�"�x^cu�-�x���Y��BB��m�aM�Ӌ�I�lY;�]ץ>:�H1L�v�F�׏"DͤI���U^7����'�q�h!���@.)���m�0����޸�H?y�P'#�;S#`1�}�=ꙮ�&d�s#�84Q���6��U1Z�a'1\��d_���Qk�#W�V i^GJz���uj�Z�WZ�K:d���P��oz�U�B�^�G��Y5 ��S�=ϥ����V��.fS[��[@L3��H�
߼&F���K��M�W����S!���Z�P�'��9��;y�e�_!���S�}%��v���ש��Q!��z��[�M(X���Y�CE�S�Fd�SLI�c��o:n;4v(�!4M �-)-]1~ɍS�S�O0�۪��Zm$���w��Y��Mq�b��{!��p�.�2ZEa������QBܠ3�؛0>���]�2 �l�P62����=���������(p�
b�B��B�yL��B����[�qtc���B@�lL�<+�ۜ�{���ƴ�3�<�w���A4�J�&EM�M���v����X|;����2��Oyst��4uԇ�{<9�'M�/���E�nH���h��+������� q�h��eU��'�.7S�.p�͟�<�n&��ķ�Y�˥;nrl�n���Vl�9x�T�^\���D��$>>o��� ���۵��k� �@ *�UUU9v7r�[n�t1����]˛�48]]�v��b�m1g�+\�k�u�|�vƈ�3�n�0�9$�ڍܦ�@��ݶݰC���%q���_%�vi�طc�v���#v��
q�� W!�r)����u(kӃ'�~d���p�{���ě;G&�3��OӻXGZ,2Z���8:�5�e��/���՛�%Ft�4�,L�{̓{&��7V:��I+�(�bye:��wT&� JaH�kx����_Ƈw������{��x�K���n��:��z/l`��!1dof'�/sjX�iV1�3ta��T���UfMlf`3'
E@��r�t�����������G���1�Y�Wd����υ��'8<�/jgsډ3��_���C��}��՚�:+��L�f�����i�4w�:wNT���d9�]�T�sH[v�m��j�C�=�d�q�ι���SWG�{	�^����z��M�	�&�ᐷR6[�*��5�P�#7�Q�8i'�/�I���gxG��xL����;n{ǜ�h�G}�PN�Tn6"�B�CU�6��Z��%���;�����0�V��n����EV�r�����5^�`Q�ϯ���(�ޡL���l��פͫ�$4�u�Z�ѵ�)�ó~��q=�p�ސ!��O�Au�.����׻$��t۳w�"��*��Yf�f�<c,"_F��|W=X`"�:N6��ٻo�f�'1]�7%�%]^�x1��uL��r�Yܺ+M�@T�tzs��g��yJn�u��m�fV�]�|�\JYK���:��g���q �39��e�Z�b�>ۥg�ACnnX:��u-Y�>�v���U^u�7fe]��U�ވ#	�SEF�Ǻ;r��כ����ٲN����p�]d[���X0
f�H�����[i��M�^v�p�m.���f_�7v��y�*�V�N���aZ��&N$�sc9.���Ή �����!Ž���wn�l�a��v�cuV[˽n� �e;7J�u�[�v�Gff�o,r��0r��D̐}d�te9/u��  *�R���U T  ��   �w��    
�b�b45U]6TDӀ��l�{�      m��Հ      ߮�        
ʪ wP  
�J�  
����w<�N|����T7=��ε�Od��r=�=��ᅳ�OUl����|L�����1��p����uv�枚pp#���n�̼�j��sU�LF�6؟Iӭ��ֶ�V܃� �������3�����RS�t�ٵ�MrYm��؇'c��؜�y�v�P��T��l��μ\�瓶K���5���˚ջn8�	է2uM�1O,�s��og�i1�n(L:G����kquX獸:�H��8� ��w)�]�lz�=�2��ێ+EG8�����ċ�<�Zܳ���B]z���^k4�=��A�N�z=�]��*f���n��ް���rv��V�v�.���6�b�r#=�N{unu�v�9�]�Y���)�����g<+t;��6s���Y��c��SA�L)�t����0Ճ.�ryq�:��^c����۶��η\l �d�*D���w�l����vnT��l�<ƨ��&����ٝ���: *^yźC���w*�aݰu�^\?+|�v����%�<��]�<W��q/m��n��Lv��=a����V뎋���i�Ctu�#�G,ؚ�KHq�+0�5���K��w�|��:��T��-'M��9�v^�Ŧ�Eq	�	�a8p�}���Dt�A�����Ƥ��!!�����!�p�$�P�kw�q\��uz	!?"�m���7"���<��>��5�vݹ���z�6�������}o��%��<��2F��]g q�Me��>
ہ}���^*l;��� (e��.)��G���#vsHF��r��� �6G��O~����SF,�������]
�@zyt��v<@��L'7�ø�'�	͠��nxc�
�LY����Q��_)�҅^�+��K�;uM��f+/K�q�z}[�����k	���8-n��2(O��gD���1��?�w�F���^1��^���SI!C,��-���r%q��PO���Â=U�}���܉�&ߞ��[�]�ԛ�V�z��i�_�4m��b�:�>�a�"]��uR�����5�2^��-�ڝ��C�<�l�}���ܱ&��j��,Tv][D'>I$�H��p�4�`(Ao�������:=֐߅��O��^i�a�÷Ԟ3��a����HOl$E���.�f�ψ"}�E`r+j���D��;7,j��#IgG{�o�t��Ƙ̄�^�M�E�Gl{�X�5�� �q�ve��zD��+����G��V��h�^C#bS�rW��zu�6�OK5y���PNAx�����큚G?OL�}X��tf���Ƕػ�7"ɝY�tG���V�{����gQ�B�z���ʀv?��3����a{3|��v�]35S��ʌ�1��.D,�b�nj�^Z�B�8:�C�>��xk�~�y	���3T4CE�|W=/.���xޜ%��Y��ަ*��г�o�>�&fN��m�S��{�F���n�K��{ٰM��-�u�_O���;�`�b;��������.�KU��a�!�m����<B�8nx_]s~�����W��a��
�5�xB�+���d<<�^��Z+W�}��WB��Z,��R.�pP0M��3{jk��ח:���^j�9��l=��c	n��t"���&EuWX�ù���L��s09H�A��5�b��co�+�)J��N+6mr9�>x�^Tꕣ~�}ϝ��KE0���s�.g�s����E�ߩ��Q�:8���U���P[������T�c�6O�]�����j��h�#5,$��ӠI9xСzu,��bt��5���+i6�0l�6�oG
�X��U[��~�u�pa8Mx{�;�~�A{yt��а�8�ګr^#F����6���x���{�{l�FR��lX���OmWW��g��ŖN���N�'	����fzc �I6�m��P�p��@��#���g���k�`�ACG�n����*9J�ϵ�'��َQ�\jH߀$��0�w�E��{i�h���k(q�������B�Ҭ�\�J��$�7���"a3Q��W���Ϩ��|��.�Y��M�>� �yGAfA��&���I��=R���Rݚ��:��|_2|���?\��Fo����\O�ю9�O��٨AaCM�VEǣS�&y�r�	���?�^�ϸ�ҵ*%��Q�+Ĝ�
�ˣw؅ڸ!=��9\{`�֌���/ �[�������Z����~=n� ۸�^�;~�@@ ��iV��X6������v[�m�쭝�l��G�um�uv�9�e�
�X�p]����Ί�c��Om*�xt<H��c�6�E�� �x���-��'f�u�"G7nأ����v��{n����^�C��'[�.�m������67N�,/�����Щڬ47�ʔ}>�Q��~#�D�+��
��/r��Q���[޸z�
���K��Hq2*�,���{|�X��]�i���	l0���r�3��W�\ov<�M�H#Ri$�$�Cb7^y�0�sĎu�n2dA���oH����aV~��8O�^�ɬ0�z�#�i��Z}��9��A�ѕ�ujRW̦�pW�^��U�?�V�t{�������&�^��,�GVm�eh�$�ȷ�q�9^͋6�Q���]�e�.�Gu��V<8^b�x粚�N��>7�[./n7M�n6�M���'%7�t��临��9�+�p��#,�܇>�0e�F+��GW�G��
^Y�}.n����H�l��6���{�����.��B������� [\7��}`W~��,>W���O �Y3s�+��=s���څ�"�]P�ϛ�N��r��]O�z�)����Ѳ�ܤ�/�罼�A0�p��3;]��L���(�t�o�Q�w��� ��U��d�KXoX��+��c�6K�\;��\l���u��J ����XZ�;�߅��u���R��|cr�g4k`^�i�Nf�t�c&���ޙ���S�_r�Pxpݽ��ݷ������>��8�7�-Z��ﭿf�5	�a�VG�Ü,홡�z�<�,�{�t�q��-��.Β)!��d�T��>5%;�唷w�n��"�.�E7T40e�ښf��������I��WCD,�O*�r��l������]�8u]��^�52�4�.U�U�pz�خ��B�I�fk��mT�0!�:ٵv�;�5�Φ�fZ����Gs��5��5��L�S�duQ�qN� hǚ⻇Olm��Zm��l�jP	�Q�sX�u�;�[#y1��D4���;4s�>dV�z̶���"�j{�DCRH���y����"�J�B�����Au���V ޕj�j��:�4b�s�(b��{Ff`03su6��a�<S��Q�j�T�#4�7g}[� �Z�`$j�ܞA`w����|�Go3���Y��m=s�X$�r1�%���\�1A����ި��١�a�|2\�,��Y�a�����{��nN��h�p:<��ߧ���JL����&@�2������~鷵e��t/TJ ֚��Ϗx�S��z|�O�i�KA��ѽ��2�$�T���Pͅ��O�=����.�%���.ř'Ѝ�ۉ����y�si��,t%��U[��v�Bh��bȜ1C���	�rF��6=~�$�D���
��ǞC�F���qv
@�e��J
�A��~�V�3�4�=���6pm�σy����Oܐ�M����n�#Ĳ�L�j�G$�����Ӽ~���ng��h[I��΢��g�y�r��Џ�����Ѣ�	���63؁	��CR�b�{�������l���1 s����S4�_���F�d�h���f%���m��R���m�˂]�NC�O�"�G�4-��]}@�a�Lt��ڒc��Z(�)rfTnP�,�S98�e7�|9��2O��#���ǒ����7O��H�Sӻ�f�xT�&{�bb��XMlumo����xy�f����~���/�@.����g�\eʰ�J���l`@�r�1�
�vG������Y�o ��������i8���:w���|]'H�3�k��6+�ψk��2{��5�E��@��m���|�E�ݮ�lαG����;!C7͒��#s3fxω�����u���4\�&{���/�U5��{�T(e�1�љZ�b.f��V�'Df���4��m%�ŹYT_o8�l��W���Gd�I�7w�D����-��6�/�����`�W�Ӿ�5��[1�|��'�3۽j��4�����>�2��)3�ȉ�75YP/؋E�zNo)�Y���AЂH=��8�Fϻ0˛���En�S���Yf;�b�lL�Q��us�f�P�0�o@L�ⶥ��e�L�h 6����4� m�l�*� (0�|��8��:�rr3�f��^��9��cj6��i��q��d;hw&�;]t��-��m곩&��E.��f-�얫�e��݌��ݓ����G�Y�ȸ��oV���v�qoa4���Y��8M&�)�����mnl���!��y^ּ�:$��m�5{�4��M6��Q�#0�T9��O�MY�08�^��(�����9�0��4!�[����=���n�ݎȽy��$%z�4
zMq!a��ݘ������������o���+T�P�<�봐nm-yp�+��.��ۂt�%�z�����UYOFSGC�sW$Ⱑ�{�Mgk�Y��l���s��Æ�@���@�g�M]�jT��~=���b���z�Й�ybsG��A`��ޭ��3ÇT�u_w �0�4\:a��S/�uYbS��#����]�C�{�7(6-���U��>�����W|	�|�$B�oo�q���Kpj*r���X��I��,mֶ:�3H�c�o���Ć�a��7Ƅm��T�C�XVy�����_4�]��ϯ�t���3�p�e`Z}�˗��L\^BQ�s��t�v�w��;�����d��O�]cqM�C3���Cr��+gL�1�Ƨ�Uⳍg`�gwΡ"I�86t�K��f��.F���1^��V����%,�Yb.3��P��$�ێ��p��|==�[]vI �C��M a�#��=B����[ȸ�
�kL�ȭ�8�N��>�wXc�U�M=��&�a�A����8�ʇ�_�L�,�ax'^/�:6���݈1�PS�Ly^�'h�n���	��a�Bx`���^lW�Q�K|h���X�h���dtq�]��d�F����&��f�eFߞ�E��<s��\nB�LB	��0#ĳ�n�>P�s{î�S�+�X��''ѡM��M�����~�_��H�#G}J��>�=��	!
0x)�y����"��z�s����k�'B��F�s�c�e_�gO�L�W�j��3(k�n���&�o�R���	�p�6F��2�V��9=�6�p�9U�QL�����mq��:ŋ��x�LA@�����d�P��5���$Wt���Ǯcy��u��ZHoʞ��������!P��+�yj@��ʥY�̥�]ۻ��-�M1�M���u��W/�3���{��m#0�K���z���T�iP��޹����L����8�0��o���[P�������{��-Cj�^�댃���{-���f�1:hm�m�Jԕ?L��ZH��:�<�NEaS[}����ϬN��5�u�P��m��ig�-�d˷�ݹ�4�ravP%9��AKڶ�к;��3w�R��ri@��$g��+7s�l�ntNo%�+I�@��C�FǸ�=���,4}���o�ˋܺ�QqN�z�5iQ�|�ʃ&v;�X�Yd��p�}I
�w~N;a���>ϟ���ﯞ�����
�Wm����{q�V����6u�Wb���: /g�K��?����u?x�t|6j*毻��l_����&������m�(����l��Z��O��e���O�TVͽ���{��r�<�;�wR�*8�a�R�L�̬{rw7�6�h7S){MɯL�_�]�W�z�mɩ&mp�~�2���k�o20�����32ɚ�}�rk]���gU�r��}׸��h\Δ,�;-��D:��*�6n����{rR'��uu^u-��z�b\�u���D^v��p�޺��v��*�;�ƺ��%Ԣ�r�o��5diYtc�AU�oh՚��5�&�g�!�YU#��jd�jW�_��M�Z��+uז�͙�gU��!���@q>����w���/���X��1���X��^w�ܢ��G��3��l���DVs���'dB�.�I�@���ݝ�����Hu����q��Y6�h�tV�Dk�yv>�Ŗ��K��Կ��՘޼��Q�V��U�&�WN�ub`!�-\��;?:��<0j��7�=�Sa7݂��m�0Pr��<�ʅP�4�c��K4�M\�
t��]v)̌�G$gN���Ke赻bf*�	^�eu`&�v��}�2��_ȆWI!�c�9��V�.Ȋ����x���e��[CP�|f��U�YR�Qp��ڣ���UC`��m�E��5������A@Τt�T�j�`�7*���M�4�Pb=}�w�(b+ݼ�h�bM2	U�_'g�CݴL�8X�z؞$h���fc�o
s��>������Y����l�/���s\"�$(lGZ!{ʯ�hh�|&<�z*��L�����$�pP���F:����k5�tق�!Ch�Dyv����2�K�<�i!ݭ���)l͆�%���Q��k{�3��[��M:*y@q-½������W�U���v��7o<r:ڊ�H	����SR�[+��>�WمAL� �u%��f��x�s��UUз8�q�{�j&/����USh�: �Wݘ��=���#�V< Q��s��Z�m�+6-��W��\xd2h�<����(3޲H���]J/�v�
��8LT�9:��+6}0�����w�����"p �/U���v  USJ�UY�׳�����doUn�e�0\O8y�|�[�p�:�8kn�L��.�@��z8��_>n�e�kO����v=��tݶn�j��='hE�q�`��҄����n6fct���8�b䙱���F�[;�3�1kn��J����3��T��7�$|_a�c{jzzX����W���C! ����3Bp��7�Q��C�������3$�Z&��=��xnJ��S��/NH��1^"�X��ZԹ]�A�E�	�C�H���2��;�c�Q ��n����ӻ���i��y:�$�D2�c��	�*Eg�x����Pz�蘩<ț��ʩh� ]���6�{���/��_� �!Gн5̣8�(�gY5<�dh�g*�%цZ��`�>�uԄh�a�稻������p�輖��s�Ovx,�>5�����c{+��ڍ�	�L�ɻ43��e��g�d��?w���`��1@�� �Wm�ѕ���t�I�{���@n.�39�B3B��/|(� ��d~�#����N�SE�l�����Vv2��̱;�2��y]q��hI;�p��g�P�rx=\k���O��B�qT��h%u7d��r?�wq�bY�UeW�x��VU�w��fum4z���}�#��^�i@pIN��ܔ2��o�O({�$�Y�7� SM��M ðu�Ntv۝�PLe�)i L�!( ���;�E��(���w%�\r	)k~'lo^XO#�#���}��ە�>�n��A�	o����f�9*j΍:�����V�$�;�y{�~�z,lQ0�HG.蔧R��<WgC�w�t6���T M�6'�d"�jf;d�S�B�'�05�u���+�Z��7�*&Q2��/��N.��q���T���.Y���F7� Q� �Wu�4±���=���]�'�W{Gض�L9�����H��=6�^�w]e��n����$��Z��(�ˊ&ɩ�d��"�ʘ>ڸB/�K9�z�� O���}�u�ln�ՔD�����9W[�wu�a��pDTYX�ƗU��%�kW�.�R'I��L�So5����pq=��w͂��%6FT�-��u���i�򪐼d�����k�  X���@<>�q���4ghv��z���y�Z�*�I�\_\��^�)X��r[���3=�`�(	tCM�i���" ���:�)��0����[�#�W�d����T�ggL�+{wΤPuKז��of��ЋJp�/K�L�
�MP�y5e��x�ɱ".|ߨy\���'�Zq�1�>���ս>���j˱���+��郀h��0�,ً�ށ<(P�1�{��`b�୾Li~t�'��Z!�َ��gH�C�<nuo�.�)0�W{^ve�5��43BJ򥚿x���K�68�䑽���q�:��0���]]�/g�H��u�/�֕0ˆ���,g̦ٸ4,���Gd₫����;�nz���F7Q���Rq���/�hE�֡�����zcx��1w���4�ֺ����&Z�z{ɋ~�א�$�i��{L�9�P"����t��A�K<ȓG!w)������v���.���74������`���X%e�s�nL���}DQf~�s/�o4�ѹg:G�����5��N�Ĺ˼��Yh#������OEw�Kj�٧Y�li~h
/�W�vJ�����w���׺�G�H#���r�z�4�	������֭4�a"R�ѻ�S"�`Dk�w�����T�����}^���D���n>S|"���e�M�w���q.�F�54V;#��p� 3�j�	�ʇ�u>}��"`6����g��漻�{86˂�KЦ�Cm\ș
t�r�l��Z,�����qZ�V��g%[V� Iz��P���.u�*H^�{0��<z�0^���x���^����Ozo}��,̷�y~x%��i��I(��S|�Eh+���xN�'�������o��<x(ɞ��Y�</9c�}탣�m$a���P��U�6slC�X-U��:�mU<��N�i�]V�#��:���Fc%��D�P��� �'2�ɸgL��MA���ݖY�27N���ץ)[�����
�ʸv���陛�?m��;y�V�t�3��w�fڼ��w��������u�P۸�6鴀+��� Jʴ�UGh�i���i���ͬ�F�����`�+ݼԝ�����S���֍ݒɭ�q?���q��n}Fqɦ�T�!���u���0�s�;����n���#��۝�7Z������(���[t4��=�M3/!��^�t�<8i����m�_5Pk�9KZ?��z&U-���'�|��{4���6G�n�;�h��wk���᥂s����ӯ�c6��l �v�oN��rlf�����'oPw��[jM$݄I�b�T
�	�`��'�d`�$�Q:�(�KV��^q'$��VP
,�� �����u�3b��ż�>,1����ā�[5#%f��;�^�N�h��)��^�(�-W����ST�ٞ��(�J�Q�J1}��7꒕���'��;NX�Q0=���g�7=ݨRNM�4��n�Z��"�9������;9���c2���l[�)����+g��G�Y��L�Zpg���M]�gD�h��{�	<�w�٘�X������UW�̋���;�Z�7p�[�i��d��^ܺ=�P���&�N��GME	��g�x���&�Y��-˝nj\��Zp.#<o�檍)�r��	�[�ַ//bѴ�;��v�[i�ae��)�{����I��Fy讻]��͌'�:\6� �������VdWq�	i����M�@��m������cv7l7^݅�0pJb�b���wJ����"�g�s
	V��.�X�
1�����@w<����&B-��~^}L�'��s>J$��IS�=ז����M%;�n��Ɲ=Y��Vz��yN=f��S�J�LE	�%ꃽ�P�M/c��������c;2tsSI��[�mR�����>�0/1�;���a8� ����rF-����n�0��	@.)�~;f�Ƶ��K����O�NoD��G�^���ţv�����o�?ƥ���A��_,������6�7M�M�j4\�'�͞�*�Q���f��=� �v��wg6K^˧u��]�؟x�c��N@`4����05��R�T���*������J-��m$_{�u�w�+�2�!�,l3��p��b��_LI�\�$=��o܈��\]q����n�q79�O��뭐ԩ��q���Ŏ�dڛ�Xқ�˘u��(��n��h"��n71~��d��6�A��3S/-`���\ʨ��� ���[w�>�ն�=����:+�J��$�����g��Ӟ3x6��Sj��I{��q_�����qj1+��Κ�Q�h?t*�{2��H��NL��Λ�N� ��w�+N�8ҙy�v`�� �O�w)G�J�ה�:!
=��]T�N�5tJ��V#uU̍���,����U��&�_��:R���JU�}�5}�f�{r�ģ���X�1mE�\�nh 4lnir���\1ԇ���[�U\}&����)�[N��zx���'�P�i|K����~}w�~�J+ݷG6��q髁�Tc\��qb㙖��0]r��S6e)>��S
�!�V��ɗ�����r6��ޡ���zd���ƾU�F�k��W�1����.ޞV���߷�7y���!z6r�#���n��+R��l�wo�-��O�F� �y��[�pԡ�r��^Te-�6�]��~�!TŦ'K��λ�ڢM�9���'ζ~=�.����1/�;̛��%{tVq��v����ښk��zC����26�&�d��0M9g�|��ֶ�K}��=Kh�ӻ�ؘ=�NV�r�Ɋ�_v�ɤ&ixv�+��8�{OAf	���)�롐o(���㡭VxƭQ�9S�Yc`Z(宷[mn6+hT�ٵ���L�lLʎ����PpA吔 ��a�.^�F�p�^ t{��$�6�m�iZL#
�D�VOGZ�Պ=j�D/�`�&	�/=�Ŏ��&�F��^��Z�C���А<|7/���ͯ{�)�tf�l1�\s5�9Û��y=��#
�(Rk����mՕѶ��`)9�O�{\��"h�M$=�S�	��76SY�ܷ��\ \g��o�f�}�];�3&7�×�e��g��f-��$��^�f���|�H����݋��C�������	b=5A^A��۳��8� �����GL��\�Nl��mʘe��jY)i�a��������������oϏW�����~  �;�b�i� V� ^� �U ۋ����|�!��=�k�G����m�{[�׳ɶ�����0���;�;l�h�GK��v�h�<�$�9���{6��W�z�MO/���jXá�*�r�\GW�mX{�	�r+y�'b����5�ɀ$�����'4��?w~2��G�yz�0,��;g=������)�X	�&a����(�>��d���%�Z3b�������;�x߄���F�g���gN��]K���I���0�m��J�"�U~��O�!�j�|JX8~>�o�?L �Z���e�)r��Xz
���0�l�eH��l���Wl��O���~T&�h>�^ꫡaSjU�F�"ƻ���9�<�a�� ��҇��3����TM�7w�(9QH�86�މ�1�dM�o�k�#�>Q�#�`�k�4��x�+>i��7ͮ��z���^X�7A�>`t�d4���##w��S���ߏ�x�m���s(�Y�3n?�v!���*��:'�I���<]�_���J�>(
�T�F}Fi"H�Dۜ�^Z
z��{ձT�&P�*5��(���Ʒ�}����d#sq6�*�i	�n�:�>�r��*���4�!j�ծz��c�2a��n24ӊ7���pt:�u� �Cھo�ev:��%��{��w݈�e3ZݳPd�Z(b˛�d,ʅe0kW�S�ն`�|�t��#z�-�}Ϛ��G}��&�VZ��ʽ�����2h��fA��a��w9�2����"��!�n��n���+�x�x���Z�4L�}R�fvmguŗٙy��b9�M̨r�H��]0�Nbo�=z�iE��R��T�2*���R�H�WMlh@�j'7f�����!� dWX�X��;B��6��eR�θGc!s�#q�:y!Օ��"�-GdO/VO7���#HJ���~��U����i�c=�,���ϥ뾟u_<�µ��'j*�!F�P�fԘ��$��
-��.�O��6��5X��fcX���L�F�X e"���]�_ܧ��4潱|�eg��ފvW2�Z45�_f���r��*��q�1�ufm�{���6�dK ��,)1���z�{L+�����T���w��m��m��m��sр         U*��     �*�6�
����ݛ�uն       ��3j       7�f��U       P
�0   
�     l�5G\x՘��9�8�f��t'�"���m�m��Og!�lz
'�qq��NC������ݸ��]��9}�\��=f��õ�qcN�+�5�g�����|��t��f�]���OY�����O\Hc�v�#�(�p=�:�nnۥ9��s��u���J޽Gk�׭�׷���3ל�kpg��&�u�٫d�v������^#�m�b�g0�oWQ��ɺ�x���iB|��"��ؔ�e�����B�-�,;k������\iu=�ܽ��1�����n�m8R�ig���/k���פ;2L�л;�/:ۃJ�nO<ͮ^�Cٲ�wS�e�=���q�Y�6�5��v�F-0�,������3͵����gOh�uKs����ث��b=�b^��[p�v-k�U��^��l���X5ĩfx7;�X[�6�=�Ʉzs�$[p\1�뮞\����tӣscC=Rk���%���+���������s{��z�nU3��<Ⴛ8�M�,�����l�Gln��M]��ip������3��mї��@ub���r�E�b�<��btW<��F��q�kWGnu�c�q��q�|~<]��st�7�ވ{:�=C�G&��d�7;��7g�M��O�݋�m���A�/���������z���߼l9���l�e���HwY;��N�ʑR�;���X)-�Kl8D�@v��:�RWn}��ʝ��*8i��l�w���i٥��r.��蠡ny�ė��gö�z:LL��LD�r�m��)�����b���N�D�O�$�#��5�.kK�0���\��T��Ha���M��G6^�K�Jg{�f{����Y�L�*h(4�|DLp�aY(�3/ގ�]z��Ҭ�%q�=^�mĩ��"�g�x���5Q���%�I�Q��]�$��~��Yų�"a莛ؕw +
�L�iu�-�2L���(>�ሮ��=c{`6�a&��SW�ֹ�U{ �
��^�|�	��@Ӆ9��M` x�0�}�RwK�1Q=�E�S�׼��|@�/ت2�w��ލ$g@E�Q��j�w5Wb��i����\M��m����`؝Z-��͊p��m��	�Rfi�e�̀7���m�1����:(��\?jn �#����X�A���Gk9y��⫷����Hd���ܼ��,�ap�s�;�e캻���PN1�H�{�3uz�=��&(��$N+�!�\�����9�j��2!#헑`x�Ǒm?�s�v �b�;~�>����X\*Zd�ǳTgeL�p#�6�ۖ�y���$�G��W�7ɷ9�a�[aX\�M�8�����)C^ �ޡGf�M�Sf�0�����C�֌r����G.��J]�ޛ��*[	'���N�����V���.s�~�V/M9���j�����
���E��,"�>ǫe3���[k��B"��j����ѳ
!0�5�M�����J�x.yTV�̼=��ͯ2�-2JJ���/��f�x�Z�t;��ixq������O�,Φg��P8w��#:W�U�!L��磨��#3��F��\�m��i@a�N����Vm�}f�P̹ٞ+����e�;��@_���ِI�4���M��;�P�p��f����E�P1ꑂ sV�Ɲf{�V�O��;؍6�����-��Ӿ�l��=�ں/���I!e��X�$xQ_3w�5[����I#7�L�`�N�{�=���*�ת 2q�*ĩ��6���Řo�ӄ�`o�&��X��lq~q�vzkӞ*������2:LdWT�U�\�=Ej�����
p�2���^���N*���nq�am����F��}����TM��b��K��E_�����M\���
�@���$�Wy�k��FuCq1�s=�U4\�4��@��I�Kp8�̗N{@�؍ֈ�� �	��܀��l����J��41��9Oi���T���ݾv�剕
h$��K��4��|��ϲ����hh�m�z��Eb�o���m�	~��{V���c�{�	6�$�F���!&Fb�ϻ<�����l#
�:��l�^u�8,�r `���ܝ�
��P�if�5I/�;�P����C��N�R�ge�hfUX��E�=�Tr���q��]��V1z��z�aG�ԁA���Iv�rn�=P�/�0�F�HfnM�zP~p�	6�m��%��mt@�~«� *� ���t��~��7<���y�1q��ٺ�㳷��a��s�H3���c� e�oJ�]���ri����\mͮ�v�]�v/���5�]�y8�ƎԽn�'x�窭u�z��m���d���1�h|���^w����c�
+�|2MAH��y��S��4�b���H0�����u��.����mݡ���{�T�Q�8�9~���8���7��u�0K���b������R<"}ʣ'�r��ZX�ˡ�%.&�� ���Q���¦�mӟ`ttn�m8_�!��=.�2�e�Nz9�����ݴ�Gb��:�r�䤈.���0D�Ϧ�ͺ���������3nMH����	c�W O�����U2ix�����G����֡th�Lč�v����R,�>�ewT��@C��Z7�p*��W����/'\qW�F���Nצ��(�i����f+Z@Tr�Ŕ{}1<Y%w��F�Ǒ�Zϻ����I��h>�u*���L���9��HJ�9}~εO'Ɣ��S9�~�;JM�}�I��I�TgbJy9��|�2_̗��	�ɣ�y'o�ڧ��� 8՛�d�$`�;bx5܎A���ªR�<�0�]ӥv�7�ڻ�� �*�4]�PΓ����,������]�u]�|:q5�zaOJ�f'�Ps�������@!�a��:���k6�1$���A����H�D*�SE�ݮ
z�t�a�R��Q"��L���;{��G5xxyP�����;'��bz,��p�x�@����P�Us3ؽ�@��P��IWfVˣ�ŠL	]��l��/��9�P�-F��y�)[�$X�	�X����L�j5â�ǑU�����	��o��j3݆�_��"�D��=ߴz�s��G�n^o��&r�ǆ��3�w��}�QY��4�طkܧ/�БM��Ğ,B�'=�R4�s���˯�DFH��΅��H;u�w�?���%�Rc�@�|w��K����d����j2(M�*_��N�g�=�h��X�g�\
�ȅ=q7�h�w ��{���~MV�ͦ�%iλ��~��%Ap�h�s~V�y���{$`�)�Z�����*�����'$�M'�,B	6��� J%��_��*gmhA;��n�S:K��Y�����p`��z@����>e�3�W���A��"e+S-���)�G[�h����X�V��%�g9K��,l-R��=��=�u8?&p#���g������Ō��g�I�:�n����!��p��/ր���^w	���uQ8��<}�E_�t���M��}�u���\���u�M���ä����=KBw�K�i"����$ȀtRk|뻡�`}�T���X����4�n3hC�Yut#�7=�9��:χ;��	�d�ڵ/%(��
.+����m]:>�!Y�.6{�f�6�h4�'h��+Y��q�P��d�`�>�s�ڔxR����#�W��7�~��o=$p�<A=}|k4<�f
m"�-Of���{"lTO���}��������_�U���w�[����kSt��yp���
M d��%�T�d�QS#��T�~ڕd@�2���(`�>��r���؝���[-�A̳*q�p>��H����B�r���;|�I��Y��'z��ժ	����>N���M<sE��j_�c6{AE����L�^�	ޫ���B��6`VW�̫��9-���/�1sj�F(��[��u��Y믟������y�zeAܒ�X��7�cG��y+ ���|�J>�x;v|B��W�{Bn�-�T(E�D�`�$�]_�N�rj ��ֽaՁ1s.�N�_�J�ɫ��LB�Ywy1o|���Y����˭u���qlm/f���νŃ[�$	�* �6���׏�ޑ&y .׷<}� p�#cò�S�W\1��=��ٍ�Igd�/n`	�KH�BY�L��ݫ���Hē�$�����^�0�`UT��Y:zv�Ξ����$�?��l	�Re�
3��ݩ"�w�##3�r�V]���%E,FQN0��[�����0�v{�t���F�NM��N���=	ܝ�,�y(';g������l �O���V Z5<����[cx�C,۷%߰� �Ne%g����i�gT�e��F�S­�yL���k�ݛn{�2Mp�0����s��^��"���ȳ�<��l��JF��Rj�Ӭ��ʇ��r�;n�����7�S"�
�ا`C����C���eo Z����f�8���ڑ}Mn@��S:+ѽֺa���ߗ�ֺ o`\�y�  �|m�� ��Z����b��\���W)�c��g�Qy\S7c���G�3�6�u �o�n��ذ���3���W�h�:݆���]��{M�#w%�:�l뗺��f\%ny癊��^Ngۗ)�8δݶ��7-�u�{��������d��>�}%�$���8�����{ҝ1��ZI�
f6�OU{���8�3���O	��}��f�D�+M��tMp�~�*-�J>>��=nàN������v�u</�It&�8-w�����^��DG�J4���%�m�ڒ�*/�L�]��lQuڊe�
	I �,3^��Ή�9ʅ��ao��*�q�*�Ɯ�Cj��/������_�8J��A09�}�� �rr��2�
&go)����v��06��>�~� v�OQ.�b(��]�c�,#6bch�Or���tl9�Bïs���6;�̄��}x�:��ɡl��jH�����UTB��/�׬��^��5��i� � �b��'B"�<���m5�4�x��[t���e���kn߄1�B<_w3WP�n<���ٹ�렠w��I4�N{�f�7v���\�_�$�'M��X=�޿c�YAثL.]S��Gk�td�*�f��^��.�S��Mni!X��U|o{�a�Gr6n/�~Zg�gM����p����m���ۡL���R�!|��M�Q�6�f��up�]��j�j�ёbݸ��E����,�vɰ����罨1b�&<=����gZ�<wf�nȎ�ͨL�Ur�,ɓ�67o��o۽	8e�N"xn��)]�>�S��
X�9{'ѻv�$#o�ww���.v�W�a��uZ!EZ�3������<4��&�X�2*:�}�QSgc(TrKm��z�DB�Q�{�h�֟i:d!p���S]T���9������N�̺��;��A)_���a��Ϫ���Ж�c�@��M�Y[<<d��H~,#������>��[���J�������0�=�}=��)be�H9�dt��x�`\����O��W!UC�ʧ2r��WU�d���ߗnv����M�6eg?x�h��o�N˻�#XA6�N&͠>�h��/z�!�5���6/��^R�D��H��x.3���m:�k��p~NZl�0>Qr=�3r�8(���隑pc|G.�'���87
'���ܚ���}��&J6j��W����\�)i�,�ζ�7�Y�rΔF��.oSv�w����EC`: z��5u�'�����u�	��.��u]�>2����3���KCn_�Zq����y<��ʽ��@�h20w�}:c4��ހwL1���T�]i���[RMu����;iV��i�.�I���E�	w7.��f�m�� '`*�a�^+�3������Uu9��{�)�޼$P��kuk;VҖ�e�FdL��1��<E�{�1���\mW�� �`�^g����r����r\ow��I�i��N.���8���z�ޱ����K�(��s���i��9	��1<���ji�u0sMZZ7o�
P������8l��F۱�']��m��h�c�?>$��T(����]
��2��=��HIa_����&s�;R+2��j�Ϫ�W�=�n ���
γ3~�s��z<o['�Ϣ_$�޹	����ko�������	�J��+ƨ�
����՗�F Y�3�&��K ���(}���K�y
�
�)5)�lϮibO��r�-�da�O'T���5
U��O%LCq�+��P��}�kw1�ck��\|+<h�:�l���{;��{���b8��t+:���s]��}:�	
G��L�{n�d��wH�A☊�~{���1�������qqlc����K�屔'rd�v����1b��.�[JQGJ���M�p�5[W�(�]���2��W�=lq����SF-��gR#0;75;�CNi:9֪��)���E���s�S���*�a���}��Ԭ|7��{w�HԢ�_A�>���Ԯ�{�G�Y[��f����i�Ŝ�W(�"��^wm��� �:��շrӤ�+��)����meq���
���wJ�U�2��f^���MĬ�(�ٗ�'ly1Wt���镻0�^[�i�!`�v��s$o�T�mv�)v�XD�8u�yy�l�R��I��t����"ar"��4iFCP�ڿT$���=��k[gA3k��{W'�l�����~�%QO��bL3�6Mm����3>�r���	o�����-��	��D�إ3��Û�9}��FN��ɋ#�.q]�Rze�a�>�HW�#h�';����6J utL��5d���0��Sɖ4�.W�u��j~ni�ׯ�ji��<z|��+��@�J=7O	*���A�Yd���e���CИ@�G<��c���n�w3��������7��J�[>��,�X3�g������)�+�.a{~+;���\Pg����v���@���pݛ���6B:�O���rug{֤t{�H��,�AAS�i�Vj{˿\e�o4e-�"���$K���R�������c�=�荶[f�uuAu`(׽nb�;x�-��ʍ��f|2�3�wm�s�b0�H=/zk�]#�J�Y����:���S�@b js1,�v�{��@�+�)\�5��6�	Ğ>&��PZk\w)�n��GW���Br���k�R}�SN�d��Ǆ��֙�4SVs�ׂ���̫�h�Ϟ��������� ��mƖ��@���   ;�U����wg��u�μ(�E�n�K۱��(G�W��o\�2�x5G��(�y��t�v,]����I���3�m������9oml����q����}�zf�ڢzZ����>k��xҶ=v�v�ʝsp����ߡmeUk����N��R&��Lǿ$�����|{�������H,�1q������/$�*G�|%|;�˞;>\u�+�i֝�\��pGfц�(Q�R�x��zל޿M��h
� Ҁ�ċ����y��̕^n���������yjX�B��ّn2^q��洦�{q�q��+s<g�h��̱+ʵ�L��˅x�BܙP���S3X]�X9 �P`�����)�'>�L)"�r� ����ū�={{~�D��z$Qo��o���'��r�_tv�"� ���_k��r��y>�v1�3��w�~T��+ו���1Ʌ3�>��9��>Qz�ٽsip��ni�����ra��S�Jv-�����n���<
t�"*	v`-cUzv�^�<Ҁ|�s��y7����ψgՒ�5cjX���X���z�b�f�h�Aaju��v���Fcn7�ٻi
�!A�Zoz�9�#'d�ʏ�s�~S<<�����;w�/-7k�r�=pgY����xV����n��v!�unl
�*�O�x��3� i~-��D�ӥ�`�À	L"�{��M���/������߿{?���b�x{c��^Ô��k�[cmʹi���J��A��}�ΤW�\�aB|��y$&�.�Q�C�����Q&q�=��|�	�d�^g�~�f�A��R�(�U�m��
	3����*��U�s@c��X����D�ͽ��\"��H1���Uv��*�*;O��mf��a4���p��t�z�W7M9���D�^Sǽ�6�n|(Py�i���l{�{�����k۸�'H��{K��o*ja�r��(�,���0Dr�;~��U�8�Y(6D���qs
Ԛ�.l��<j���>  �D����D�Yd�;]N��x��0Z��}����̂M�>�ߝ\'��~[�޿M�=�Q�׳ՖP;W�͍Jq�ҫ��>��`�gk���7A� 2�T�:���.���k�b%���W��
�ݗ�7�l�ի%�n;bƝ�F��J�V�s��f)�)׳:��h@/"�w39�~U]�H�c��I[���YQj��L�ʝ�����f7f�|��wf��k0��.Vβ<�	�_��O�@6�E�/dh�޻����-��5�)���e��y����2�=�R=T�����A0A�j�����Bp�t����%�~L�$��ŹZ�"�IZ�)�:�\�n��2�.o���4G?gW^��g���b�)�%�}�A�a6�fE�{T`�NeEe	:Z���l�5�o�JQ ���0c6<̡��Ԉ��('_�i�8�D��p< p����SH�%nnxQ����+A�5���}sӎ��s9�xj�I�J���oeo���{ڦnBG
���3��oz�^�l`�lT�"K��0ta��ݮ]?'�GϏ*����י�ۮ�ü��.w�w���÷�^�e�����~���?�J,ߍ�q95���� �#��s[;T'Ozlom�����w�:�N*i���Rcg�=�+7����2K��صw ��B���b�̂X���kF$����]l*�$�V����[�&�
#��(ӿXb�q��(�Rܟ��c���e���]�hئ"C ���M�zl�c߼32��-����O�Z8��kzg� f{�P�5�s�1ƟO�p@�bhU�R���w%̔���ӳ�vʽO6W�U�LI�].d��P'�5>��1�����x���ͺ�oan��%
������L�j�i����|�49�߻� z��tJ[�Y���m�>>3ӷmQ�A�9�%uU�:8����D�{.���r@6M�r{LH��~�&��#c����O���ɯ#��m��#<%�����B	�-��"��� 8p��{��(nҋç�b��Vy���v7���}� ('�c��v������ �M4A��,���Þ��g�5/D����Eϗi���۽o4�Ɵc3���C���A��×�-�_9�zsK��&���2|Mͷ��zE�p�t�<K��]҇��?qڦ���fE��*oWC���һލ3��a���nOp�j��YQg��2iQ�r�1.iY4!4�?��*�fez�t��y���7_��+�}{z!���2�.�}�1�k.<H�]֘iwP m�++f���n ���� *���n��(<��5FF�!��=�gnz��� �-�s�ۜ����n6��9�F�<prE�;iة�9��i<S���*���OO�6�w.�8Ĝ���v��yA1���
�8�F��L�.כp��^�'���������k��M�aCrS���zk%4�N�䇽sӛcR[&d���74uP�31և�#��^ե\�G'�ꠈ�Y��k�*Iw�uu�{.}V&�E#�G}��;�h�9��~��Q+��(���\Ʉ�tQ�F�pa{)N�bB�3w��>i��M���D��O)�>]�|�c�9"���89�o���AVj��#���^�C��Wt�>���
��%�;-���scw:�e����T���%�R��Ȁ��Q��6�Rِ�j�`M�������I�{d����j�	�P:����3 i��N=#}�r`�[D�A �3Ukή�@��2��f@)!&6��cݖ�hM+ZQ��//��b?a9�R���C�0��Tэ��m�L0HN�+o�ʉN��Pe_�3������~�D���\��pX��#�b�b�zfG֏�Afь$�^�vcp^?:���P`��|�V�H�ގ�Ip��wa���⃤���g��4�� �#5ӏ#��j� @L��6G��UH�Uk��s^��u��.�Wv'���rϳB���Xܣ=z2uQ+D��)���f���`R����Jܕ�����E�[�f*n&z�v�X	�i'5$�b<`#~�RDq�d�5tω���i4�.��g��[u؛V�ūj��=�Y{�y�=����w����w?={�J>K�EZk}�F�L~�A�Q���\�4���bY��n+ˇ���n�;�H4�!C���G̟�J~�]�01��l=�m|~������Ǽ�1�Ν˃�"j�q��-��H�)�t��W���Z��(H���T(pe�� }J~���2��.���{Y|�B�B> ���������U�s��۩c�%�H�q!y}���$���f3��DJ�G��"�j��do���r&mLׁIE����n�1�E[Q }B=���3��U!x���1q�b$B|��$g��9��󃩺#�W΂�7��og&$P�0�@�qD�fӇ4��~}�4@P���/�L��&cn`��>"$���eMJ��A���PY��"Q��v��~��! F��ď�!(�.�	*��K�&�&)�*g�lU����|Exb3�DF#	�)�"����q	�\ui?2~�m1�����3)L��~��u�q�jT$�%��P��_4cql��u�^ìm<�CTA2�}8���U�	�q�W��P�p��0(���Z	�a	p��~~�u0������;3��w5�;��ۺ�Ʀ+'y�W��j��M�	�<��9k/@��`vb�뉱W|�՞5x�R.�Y�8o�<�{ꯤ_�u(!6!��H}��8b�<���۞�c��1yE��#�ي¬�c��x|��D`��r/0�����bb%���b`F#����e#�(��"Ǆ���������H2��?oS/B vaщ��R�\��܀0 	�,BG$�S}�nG�"�q1�@�-�"f�g���#�&4��#DA�P����D���\;?`'TxD1#�(A��n�{8�l��d�1�bG��Rp��c�}�+f(L�A�>eկz��Xb�:@��{;�����!�l�/�����OvP��e� }�~�0Z8o�L���:cQ�x%C��a��nD1��*�e�a�b� ��"�eG�޴�0g^c��Z���j��IKVe,�|��H������#�>�DD���`
�_C�=�v�b#tǚ��ڳ]9�>�d�Iq�2�@�뮹��j@�I�w��Dm��~����B$+̩rc�� ���R.�Pb�g+g��BP̲����>|��L���k����e!�`8&��$z?D���f�^!#BV��!$�1&=C��������>~K�D�\�n�0�t�E��"t!o�q��E_�<&���j%�p�uh��U����*>�~��)}xxc�#�Y	G�'��f�G��]�~���t}G#sQ '=٨�#ȑE��F ��|�V�M�9*|D��4#�yŒ��3 �
�p่�D@�o|�1xlGL�����FD�a��Y�\�2I����u͜��]�����D���.kC�8{CʿW��MV��	����f�e�����9��ڠf����my^e}c����
CD�0DH�Q�"&w�g�$p���,G�M��� �~���`H�6[flA�1��8�2��� ��Z? |�q�GЄ���X�O��W��>���"��D!	����S,D|T����1�����"G���>?��-@��S�/����v��驓�v�����x�͈��Q���F�C�|�]Z�!i��E�&�_}��u~t$��B),���tb.��F>��[�H���i{�B$A ��͉u��� ��و�G�A |G�v��/���!�>���{z�6�m&%�#&S�t��Wl����	���@�������Rv�Qc�|����##Rf�
���G�FA1B%r�I�GRݩ���&6	�	�!���H�Z(��޺�F}}���Js	*TҊLjB2"�2B�*<9�^	A�Q�����	����i)���4>!���Af"��o�:�{���8~�:��g�|A� ��8�F8����!c��y6b��B"��t'34�h(p���"�0�(�B��U?��˨�d6�����b��1}�"�ɟ�b?| p ߗ�q@;o�-DƏ����vc�)Ԙ�}n��w_�>��A+D�_D�,*�:��oГ-��>�!�Qa9�MT#���6i�+ ����F ����ފ�*^^� 8+�.T�ɘf,�`�5�>S=v@��b�_������]\S�� Uw�f�͔���@pU [  ���Gk�����[[�V���\��v����*]�'�gr]�Y�͞�۱Uӹ���e�h��l�Փ>�:�{�{/Q��^��گ9�D��V�c���:��r�m�=u�K#�fݥ$ǵ�m�<�ݱ�p�i|��$(-C0�0	�ڨ}+�8��3�Q!���� ����j ��}w�w�phB(≪Q!�ZBF��'�x�A2�-�F�·�9�z4E���Ǎ����LCm|�P�N%��\�:�� �x�a?-F�G�g���DE�4r��>�I0F�7���bx�i|DCH���sI����0�)�3G��$�>�1,��r�]T�i������H���������~�����JW/K�6��ۂ�m��q��-\y�AP=F/w]>i�$�pAne�q�S��*+K�D�2�/�1f�۾S#���D�ێ�}7�������(ᄛ3(ް��҅��9Y�fD@����K��$�]ݑ������HD�w�D;�tr�?0|Dy�wkCFQ�tj��" �0�͗�s�S���b���
l0n�/�C�*n�f�0�<ji	q�����2��G� �Z��0N��8��_�6��=��}C���(�UA[ƹ�!�a�������7��	�=*��l?�L���dÒ(�C��TØ�s{5�K���w�A��d��&��La�ڗ� ������t��"��j�_{ޗOoǣ�j�@N=a"]xZ����A佾�����ip�H^�oY��T~aA[�#Wv����#c�糂=��E�[�Q��>��SCT&������޴��F�s�v�����8��2���eer8�\�p���՜���vM��)8P��(e�R!����vu3�CC�nL�����d�r��R܌����wvΎ��p���]��/w+t�)�#/�
��$�&^B�B@󀸆6*Y
I�]��w3XѴ������	�t��A���;.�
@eր����ԷY��Υ��s�˴:�d�_^'�FQ+��.�B̎���v���wu�ɖ��&Cʰl�!�������Tus؟�5Z�K��:�����N�a�d�ٞՏQ#l.8M�~Y�[�f�;Y?`�2���z3{���h9}�m�²{/j:ӕ����ӕc@�u�C��CC޼�:Ы���Y��@��r�j���uQ��gf*�·�|���t�r���J�����9[�)�l�={���e�7�V�+\�ŴE�[�#)X��R�)��7��=9_3j��:ͽ�.�:h���VOZ�{`U�)��  �m��ٹ�      P J��w@    �R�'`p{���;�w:@      6���      �]�j��B�    
� ��    *�    �����qN�Xz�.r��W��m���C���sv�k�ܡ�쎬�#������wep�!��X�(7�X���:�K��w]���/�k��In8;p��t�ui�:��$.y.�<r�iv��[s��V���Æ����nNLqǪ�u�(4�m蹚�TE���b�ʦ��tK�l0��nu8,�h�]�x�c�p�����+��ηdyH-���9�[3�����{���c��@R�]>3d�h71"tgbs�{]��"�1u�d�i��盓�JWO;'���L<Jr�]v�uq랈�vw�|�˃W��z
pv�q۞Y��\��Q�6;v�k[����0Y뮫Z�7[<��lg��-��a:�ě�(n��Q�:�۷a��;n����'u�u׍i�����S�cX`�Ӳ�ؼ���ɹ���v8�|IN2�7d֥���m�A���K�z���f�XS��Fn]��<On"\��Ķ���k����ŎW��͙k��JNd:��������Ν�܈�%���gfË�����۶�\sڼ!��N��:�V�y�8����׷m���N����lWE/	Qc3���/��s	qXz�͸:'vn�_m��6��2���Y�\����_/�(n	��C2{�~���D�C�ŝ��?��>��9%0���T�����#�LOC%(�'��s���N�m���I&�P �AW�q�t�N/E�5�	%��2�D��U��C2jIY!r�]�#�! Dx�<ꚯ���}ѩAFL�ي���u����t"�(4��"�����({smm\Gh$O���)�'�"�b3�ގ	��.��1��C'	��Q�6��M/1��EIU����M
�r�l�ÁY^@��buݳ�a{ѱXr�~;ci��+�c�PA�%zԉ ��Ⰷ���V;��]	^��ys�,̻��~�9������߇<<��w�dWN��$S�Cq_5��wN"B�L	�JD��׹T�QV=��4���9�hs�uZ��;0�~��ПUȓ�/
r��7;�w`�e���Aco��p�xw��2���ۢ��aP��Dom)jc_i�6f;I�qn��2�'f䟼8��:���+�/Lj1�N����P�Z��w"��P��5Suqf�I���5��׬{� 
-&�]��n����c��ub�2!�Hp��� �����T��%���g���s��*�����N���:*(�PBZk�=�~�X��6h��ϔ�;r���-n]�.a}��4Yw�Wy�,}�]V�Q�y����-�$'p�GA�^�$W%��?Y�Ǫ�T�8H�]&m��)�癒^��s[�}��1Ux�Q�B �Od&��%Mvv�Xe�!��5	�t�~��aS��M�~���zꉈA4l����x38�%nˇ2��C���%���w�3��-�2+�#�WQxD�x�QQӠ(#�z{}^������T"�ȜEy�hP�.#wjh�0i��ڙ����׾��

�
��`B������{$î��.��x4vXB:Q�}�NC�>2P18 >4f�×��Fb�_H�%��h:�X�ia�l��wIpp��'=ߧ��￷����u�o�
��v�~���l�g��r��|A� �>L$\�G��ޗ���0�(���]���&�Q�J{S?&|hH��ڷZ�����<�AmA��#M8�t8[��Ӛ@l��iJ9$�]{Um:�29�����n �ʧ�/� a6O�+\�#���!�6}��S|�,���G�K0�R��2�Wg�b��Q'E�� �+a��٧���-�\Uv�	:��N�ف��1�#�[��)R(�3sz�����l���q�7>S&�k���ngd,���a{ue줸�Wz�$d^v����%8�*%ロI7+�B�J$�Ѡ��q�@|"bNG��%L�/�LH5֦d���z��D�|0" �3�7�^�	0M:h������z�&~Wj����Q�+z�U^�``�t�~���<��#·�՗�N�>|"������-����|t�2�.6���$ΰn�/��7_�(��ƨ�-��\�+J�K��W��ӷ+�X��'>x]�Xu�D����~�>����!��"YK��K7��Xj0H*�9���5���R��{��a��[{�뷨�j�Y�O��7L([|�i�??Y*e7�=�c��U񉽘ȭQ�ߡ��]����3~m(�_U[�B�h�Su�� ���]2�3�"t��>��
 K�wL̗[|�#�rK�ΙGf�P�X"��YسAno�n�f��A�M@n'����L���]�G�K�'}�ç�&���S��Ks�D.��	�j���(��xc�&�Lc֟Һw4�w3��f��7��� v :��U�^�]@  ?���u���z�u���a��ƃm�]�Mc
���9F��ۚ�ۉz��C�U�sMC٥u��:I���\v�rOj���n۳\�[v��ݤ��s�uz�^,�v���Ǵ�]���3�0.��M�!�uu!�c�gœ����G����U�*rP�P]�vh�L9�
���^��v � �d��{x�Fsu�ުuL���ʚ�2�����.�0�Hʠl[�ŧ;�̫�$0� <���,��%�L"��1�C��G�i�z={s��iT�@�A>����L���)[/l��==x�6�\>z��_��l�ĠP�<��sO���?$bI��wUԴ���+�w���ٓ7����Z	��z�G�=X�U4��#��.hu���&g�>���K�6@a�w4���mu�>�"��B�ET�[�&�_f�I�i��6=ڐ��]ɧ�Y��� 7�Ё�@g��z�_,�,䣋��	�S�zW�F,
�mz�Dr��l����I�^uD���oĤ�)��F3l]q���y<�u�oQ
�.�^�H�<>53�?N(����_r���5k����{7��B0�p#��٫�a�Ez����4j<P�\�kꞪ=O������ �6��Y�}��Z�*T%ZĉY����LK��e��n�95I+(��yD�ج�㆔{�,xz���-�N�u^O}�f�Йm&Ǐ�q����8�U���#��z�sc��OƔ�ZW(�v��8�S�v��Sq��[>�ju��q����|j��U�8|;�-��(�q�[Fe�"����^}��J�޾�+�m��h�r"QMy����5�:�p�UP�:�p�*I.�o�܃��@����ǋ�XlС�;��s��
Ap�u#���e����{�$w{	�$P4M�q��@#�#UqV�����d�qk�>�$��k��`���137/tnp)���Tv�C3k��ڛ����m<gUwHm��34�$�}ۗ�����uNJQ8����^���?m�A�[P��#����}�p\����}��1�_C��+�u��>'����e�zĬ�zd:GЍ���S�3vH0ۢ�l���m;���tL?�J�ߟ�������mZ�znͭ��l�����1���v9Z��Sz��c8��t�5���E�]n���%G��@�b�$�5�;���pm���D��&�j����r�7��͐�<��¯	n�8��n�b���6&L4Ap�3�խ+��~���ky40i����Y�����
#Պ�Yr�pX-�Q1Ɍ��Xpc�� ;4�[y��$��U�8��G�v�� C��wb�zw�p���K�Q�Cg�\R�;�*��_&�+����K�q�Dz��^(7{qL���L��E<�°��&O��DH�erx�dv�Y���z��G�U���|+��]'�f$�M,��}�n������p�#"}6��u���V �;}��P��Gk��d�;C�}��xP��\)�'�����$�v� �a�SՈ9��dz����r!_D��I�^) �)A��e�i��t�.7��OJt�m����cw�d�&Lz�����#����k��kCs<�������0*t�a�����ӝ7!��Ux��;����7V�ʙ3�=��?C�՞�`3sK�_�,����T��Y�n�+K(�.nEq��b߮u�>f��9�*u꘦k�OoVY�����x�*f���Iχ_jS�YRd;s�c��{��-A�]T���R�F�w�&ܬ2�RG6�|�����7����d�-���t��{!�@�,�bz�&gV]�=�WV*���@�nz��5p��%wL7���2�`���Vl�Jz�@AN����ã�ǳ.���	�0Q#;e?n����:�����(�v�1<f��z�W�n���-&P0��6fH����ߑ���}ܐJ�m��L��ZI®��cx㞻��<�*	�(��=���Q�g2����L��LE���lW��=�4���7"�I�g��ah߲*+�����W	�Z<��fʮ2����HW*���B7zEm�!�g��E�b�,�L�1�l\���N��z��2I�M�u4Q>���}]x�;�ӷ��z����X���׼�7��a��&K��K
���:fL]	��/�zEA���L�n��Nr���� �,L��f�`���t�TT�z�r���n£�rl��8V��(_�9�X���`6�`��ݵ@[@� P ;���1r��J�>��#o+�
[���6��}f���{�۱�{{��d��fW�v���-�y����ݻs�N9��n�<mZ� ���(6�N�qc��e2l��z9)χ�P`�vM3��9��M�Rp�g��"�����*�l�p�W�w�e��ͨ�oۍe����uA���{XF�Du�\�xxl���
<��#+��x��U�ˡб�F��e��O��������E���9)��`ل�
e+!E�D��UϬ	�*;���������*m�j�F5����o�7Fwk���f�04\f3������;<�
`����	�^+���ʔs[�0}{�Z{�и�X$6!u�v8��Kw�1����-�|��ł��hɼ>C�C�W����/���(��&����"=���Խ�q�[�	��r�w7f�Ъ��5�!�,��N��(�hK��)��fܭ������)"���۫����	���M�u.u��I��`�i�T?c�,�8P�Tܢ��C���φIH��T�v��Kö׹Tζc�Ld�-���!R��YN��Θ����$MׯT�p$M�A���!N��kvl^˒��ݱ�dV�+��K|ʇ�����w�};�3�����v�Ƞ�K|�ʌ3�TM�m���f�{` SA�,��#:�@��'�6]�����j�1-W9��m:�8�Οb�;n:J�{ ���/����}ԃ��X`E�h��r�8�#����S4����y�S
NAʀ�B��w�>o%F����>�v��3��/�O����0V,�/O��Y��YP#ٖ7o��RP�i_Q���![;u���7����+DN���%d��՛۽7�8p>�kئ=W:F���B���}��ɄQ	�tp�ţޭ�<#�?Fu�N�%r�a�2H>�훜TJ�n�mem*�(�W�z�fq	�h&�q<
���Wݵ�
�xgw�.�n���P�f��Kx�xL״�,��5�U�Ǩ�7<��d[-��Ơ���1mn��pU�޾����������LP��߭�����i㋧���܁�A"�'Vf���.�齭O{��Xa�5���И���U�F+V6S����m���mk"gL���wPJ��j1��"j��/e-�X��ȉnm��}����Aj�enL��+��}r�qy���T���~�k�S\� ��o�ث�Aܭ��x��,���H`�4��vZ^�E��>FF2�ɒ��!�^�8���*�4DȫXD?Kd-J�H:lh���kwN�[j�N���C�}e���¬o������`x�\���1� �x[�Q9*/��Uln�GE�-��4�7�t���d��o`�������4�91���=�h
ٸ;~�j����i�Áwn��]�����I�t[C����^z��k��#=^-H��I&�d�>)�;�����[s���×A���gn���X��bsL�Z}X�*��{.7���^9�{�:�W�̖�ބ-)��H����eV������=��+�J�[HGѷD��]��\-V�ّg.T�<
�y3N|�� /�Ug8i��45!�����dI�I�	8�ffffe*P����J��U����;�>;���n[��(�r�����CG畩ͣ%��SIQZ`Q=DLB��i�QJ��4����-�h~��T.�W|����������sbm�Ծ��=\}e���j�|�a�W�"���)b��ѩ���*�/��߯��K�r�]*P�2a:�R��e����w��ޟI���V������n��нu^��J�.�5|�_�2X-�F�<���^emV�|_	Z/�m틏;���-3�;7z틋3�f��[�������5,���J�	��DD��
�n���c9q�x�wͻ��:�U*P�<�-y9{^7��|��:�b�s�����c�?�L����oe�=FJ�9靋�|8�4|}���^m����ௗ��S�)�_Ľ%�|=ݯw��.�:T�wy"�/���/���.����r��_Y{)R���W�+ӧ�=�5�Rк>F�NR�O�}���
�o��X�-��>*v䢨Zܰ�w.67+{����}�aeÖ����ĪP�8<�W2��R?�
IOo�>�O���U��/������~?UZ���u��/G���}��u}���J�C�����J��[�G��ϣ�'r�λU�p[Ua=�ф�^^x/�OW����ܗ��j߱��5J�/wF�>�w�f�޿az��az��nqU��-�s����B��	��~�m�U�/G�ZT�zI�s[�ע�霋S��<o/Nf3
�$�����ܑN$'|<�@