BZh91AY&SY�Um��߀`p����� ����bH���$P�}>je�����(Vd�$`�R�UE d6�� ��� �0P
�5�� �� �@Y@�  ��@ST
 k@@Ph!J4SJ��
�� �Ѡ>>         k�S��(�S�����
�V�   � P@  h P`@  �������]�k��&il�U�:we�4mv�n�K��-kn�`��۵܍�u�d�pW-r[m���3���q����m�5ۻV�T;��uݷn]��ۛs��wwht;����� �$ �� f��*B�*+�Ѣ5V
KX���JUI�1��MR#`kD�JM4ƅ��m�j�*V̓�Z25M���M�RkI06i�5�E�-l�a���"� �+ @
X��D�kF56��"m�CeZ[-3L�k`��t�Zm)lm��X��[kDif�iU��,JI���d����M����X�fhm�4�)@2����h��jI6�l�J6�,�d�0�I�iK[V�b$ -)M�[d`�CV��(�UQ,*l�m��`Ym�jY���(ֆ��kE�Pn�:�%m�ղ*�X��j�3h6�K2���6֥+Z�Y5�U��2kL�U�3[Lm�X��U��kjM�-h��j.����m�v� t �h��m� ̛j-���ZmMm��`F�fBP)��Z�3Z��4�C����kJ���jֶbf�Mm�*m�&V��Ǝ�3l�*q�����3j�6�i`YB�6�YF�SKU`��-���+4-�Km�a�2�F��b�m��%$�1�����-�ʪ�D5М�PV�9P�Bi����B�"�2�P01Yjj��H�����R��m�Za`YD�3f�@�[$��k06d�fZ,��M�m�b�V���mM�4Р4h�C�͵��bȥ�����cCZSj[d�Skhae&��Fե���5@�mX�@�6�XX���F$  �4 
 )AR5-�����kZ�d(m Z�����
�Vͣ[Mm��l��m��hZ���B�ժ���P�k<�C��
��  ��z=��h�T�`d1#�10B)�IIR�      Pҟ��i�1�zh��L�i�B)� J�P� h`0��6H��y��� A� I�@�D�L	� LɀV��"\vb�c��gxY�P��B��xw���3����Ww�k��HBI�����o�]PL� T�DW�AQ�>��ǲ�~¢��>U$�X����H-D킂���u�apn��	?<BS!�Y-�CRJ`S
���Jd�Hc �))�R���S!HZ@��Z�h��@ � RB@X�[	PD* ���B�"��Z� E��@U���� [ ��	L�$�@c [!� )$�l!
I!L!!�$���Il�5*
�Q�*��,d���J@���L��B� ��@$� ����HHHHR���-���%�J`@��R�L�I B��F��V�5�*a��Кa4�L$Ē�I%%0*�&&01Z�B�@ā-�$%2[)�����R��1��?�ǚ����O�a�E�T4�a3��&1��Ċ��,R
�X�PE��F
ʪ����>����<�,���҇#�HV�)ҍVb�w�w�Nv�)&����( �M�3�ov��y��a�Bݻ6�7hcs0�&ZM!y1U�R��>�f1H��*�MqTJ�zэ�J�m[z�髗KRYom��Pt��?Xӷ5�Ө��M���T��;ń�h���p���Fu���d����4ɦE@��Y���r��:��[�Q���/&\�8pe6-��Qf&J�on��	r�vfㆶ�
�#gf�vlIi^80˨�q3yi3Q)%.��YvV!ܨk	׆�wx� Lآ�v ��y����+n� E�l��W�9��^�������B�
�%07U ��(�H)5z��{��}�P�v�����i;mn�p]���34J�.&��Qm^F!2�6d��އv2�e��*��+i����.�Њ�8�ay�YZn�u4�dZ���/U�������sH���9d��aД���DLViQBE�)5a��#̼����ٷe�����l�&�s�Ǩ-pG�j��ŽK-<�1A-��]}B�|��5��d0t�7̠]��Y��:�K(]�x7lT]Bn4��GA����@�R�\ܖn�VX��3e^:�o^d�6+��Ow}{W���Ի9�����Hbq��d4�o,��Uj�6�m��Nǭ*�Am
�����Qi���9��U�]���Z�hٺ�P���`�ݴoI;%FFY�h%5m�b��[�wJ��������/{}��ɝ�������mV��ڭ�����6ֱp��MZy 4�*9Y�T�f��Dݬ��
�M� /��N^;E�/-
�}���-�jF��Qh{Z�e�:V���l�.͌/b��y�Q��;­;�����1%��&2�-Ah	U��X.a6\�X*�E��ոʉF+�q�HNe[VYuN�:���a䧘+e��ႳFTq�r��E�r��J�jS8V3+0��Hm�S13{��pm�яn̷�or6P��F$[F��v���,⬸a̵F`���o+
�d,VJQS
j�ۥPPj��h������8*f,����i����2��Im�Xs*�\�kz��6�D��aM��Uu&�ɖ���j����ح��3@�a{CA���T%��P2!�mڸ�1e�)��=e��)՛ٌ�Ī\l�R�tc�Y�QwS)��Vf�Q��T����V��;xu��M�b��f�,3V�薷4i����ݏZÒI��[�� ᔵ��ɚ��i6=���c�B���u�V慕�J����a��XD���Snf-M}i�"�3o^M-�r[B�-��&�X�9U�*.'��*��NZ�H,?�@i9���VV9��W4�Uq`u��6��!��N<CL�{�n��{�q��s���Mhư�[��=-k��խ�{4�{wPȚn�U��f�Ѻ����ZWit�����f�}m���޻ԁ����7��'P�`c!l�@Q@�LQ�M$�5V��LB�N����IHi�v�.�)(o�L$��D�e!���e�k��Lij�1<S햚"\Z�����r�E����X��/p�ڽڅ%f��)�cff�a�X@�X�7���N�[v����%k�2�g�ҽ��ic�b�P�V��\�RB��׎ᴯ"�c�a�/�XM��O/KF�����e�a4��v�<�R��ѦK��)�63[.����vҳ����Mb�r���衵�X��w5�����KJr�%� *�Sol���F�n�Gn�XC.üz�f�Ŏ0�ׁe,ɧ`	�En��R��ёN٨�+q��d��R��)�Yy<���C-�B|X2����wY�>1c���9/1A6���]i��a�ԡ���vc��w�M
w�,��m���.�VAqV��v����]Se]ū+(�� ;�������w�/�1�GI���)w�wo��&���4�*a^f�J��1˚�7hQ6ȨRMeA�E�9F	r�M�P�܍P�X2�dpн��E]^̼,I(ZЮ��U��:$*��U�DE�aV)O7Um�m����A:6�v�P�l�����ݎnB麽���n����D�͡w[O�Ɉ�En]�y�W*L�FM̸1����Q;x�]�@��Z�[4�f.^m<qa�,��:�[���fε� �DTTp�͈��5�U�׵R�)jY�*B�UAʀ���4�Y�Dٺ�I`F���K֚%o���J`�,��YH�b$��X�5SB�)�Ȳ*�b 10H*�� ���)@ZB���$�IJ�M �h�m���y��֓Z��gkVP���e ���Q�`����ƪ�����E	 0�2�2����� �*.Nc³j�藱b��M���h�C5�,R��Q�+ZOvRyo1��q�Լ-��+{�C5�MA���V˚�ݠqÑ:#"�@�(a���;mF�	�nh�%�+	�rڹ��Ù��.e]=Y��sy�{��{)�=�-ؽ�F�iل�!�mݭǢ���@ �*�d5�W$�T�i����M� �/K�ZxE�䬻R���kkg�ܛ0ںF���U���j��b��i�v���[CD"��l:��j���S ��-^���$�"����l%��Vj-Y��͸*��Q��.��.�꧵��N%�<�n��JÙy�\���"���Cׂƥ�e�,(VG+>�gI�qo+^e���"�n�8XX�M�f�E�¢�D��w{�}���A&�v���t.&�R��̺1�%
3MX*@�^�%f���u���.�x��70��.��)����1�Y$�8ٺL`�VU�׺��udw��ϑh��c��*D��N�8dK�B�Q�!����/0[8�̱�0-�
����!	"��Y�75@�bW�SS]�r�D[*be�W��-�7p��m�V�Da.�Vaȸ�3B�ث��K�J�d�Efe�[��o~[�
��,ki�u���h�)��xpU�S�Iv��5?m�4�'�'B��w�Rߔ [���z��\�xh˫�z���T�J%S�
�w[�+V���ub�ݹ%�&�� �w��%���Ve:����xU���I�[��
�٣E�f��T����ͽяn�K�\M�Z�Iҵm츖l�sq-�U�u)�@���v�_9�=�y�֫}9fӐ��!���o���;|:��I���A6E��v�E�⧛���v�&U�6��}�!�mT���mm̨Y�W��	��k���C�W���UvL�;
h�	����é+p�tZT٘y�۲�'w���]�[QK͡�v�s3��qް�.��U����^\(i��"�˔�{�{��ԉ�2��4�HLlh1��k�GZ5�rB�L:0:���/U
D�C�Hc�
��Q)
�XǬ�X�R�ƕ��(D�&�h��) �LN������*��S8>D�����e}�b��(MX�wA�n�v��ʬ;&�TZ��	J`��Z��oE5 ��b�M;�:szk�ΐ�,B�J4��T�J� L�.9VUQJ^'rl��Ԛe^�X`Q*l�4�Vjɰ�w��V=F��[a��#[zC)F���J] �H�	\#خ<g#���]%��#(J�tʬ��H�q�r����>� p���Ҁ�6E�+2T�$�܏���It��/7kh�=��	F�s���<!F0��m���j8l4��#��2���i�Ҩ����a��aټ@�+"�nT��B�~���o�oe�-;@�Xh\@!kX�F]�mm�2��0�����IU��)Ju�b�M��B�T �сӅf�`Jɉy�q,�4r�Y����bMc!v,�6n��5��yJ�cy��Z��J����*���z��v=P�p���jⵙm�el��*V����cQ�9�lqN�S�suM�z`��e��.��R�T� �m�R�ڕ��Vc�@]���g!���U#G�fV#��:�a���2����l�#F�R3�ī�DF)*U&�,#"� ��1���	b��dKq�`�,�@�M�ܔ�42�.��a�B�BB2�,�PN�e�E��7�}��^d����ܕ��|ŝ�2��A}u%J �x]=�^�5�us3��� owQ&�ջ�w��'z�;%� ���	łK��r��;Tŷ��Ym�Y���4ۺ)a4��q�v�u�,��-"IQ�4�5��v+�w�M)c`�EI�b��ݽ̕�c{ce�L�pS7��٭�n�Ŵ\��Ǘ�xD�PL�b���t0��K
U6�ڡV`�U����ڻ(%�#�U���B�?+&��A�g��7$,��P��r�+.�#��oH;�̖�����xÒM5e=�+)8�t$��Q� /v�Y5z��yVi�
(��JH�EFJ[ �X%�A�K�.���4��r�\Yn�݂NR!dq�*���TȫLi[�,� :���+i�bׯ)�ůk%�~H�@�4��wJ��0�N:�6A�d���-7�I�]cyv���d��ٗrT*�Y�NB!THet`�J�LN�5aV�h�4��cF蠓ʟ-��T@�2#�$jU�gn0q�8�,����TM����p��2�Ԋy-�I�h�t(,�0cPS�̍�Lv�mw�6��B�A��c���s*�v�^��yAzʭ�Y�L��Ί*3ZԬ�Yܗ�y�=:�ݽw{e�]�k�M�
�{"ǵ�L��a��4�ix�B�� M�X"�DbGIK1`��Ŗo>x��]ѷt��k�N��7*m̈���tm]
��a�2hQ���״*���)֡o&�Rܵl&�7���*�v4[[����Q����a#�,�ŉ8���9ck6�T��.�%w�T6��+U��"� ��B<�̩�G���t)�pk�1��X���u�=�ia�������$ī����EHn[W�i �-F�	���Z��n9X,��:��^8�䖝���-�:@h;.�6wpK���\��H�v�)���[�a�r��ʍ��sY��.��X����)��p�FR��CU'> ��#�-�^LҖ)���]�ȧ�&�Уn;q�D�mn��(B�e1��7"8*ŪǪ�G�.r&�K���]Ŗ�($�r��pvb�8"D(xR��	b�NZ9I�����4j�&��&���zƤ�h�OoY{y�^�+2Qܼ�de�#���K6������Uw��و}h�:�6�f�m���d��GuM��cT�[j��ڕ�m��n�J�pm�Yr3�3>���Y�s[m̆�`6M�n��8���G/w(���R��e�۵[���8�����̮�We�U�f �����#z�F�X��kr�/w/��"��[�4��$�<�#�2:�Gv;&�Cb�8蓴�IvM՚�:��������U/5�۱Z���z0�N�l�+��]l�u����j�p++jȻu R�Ră�3tq3m ⁫��|.�m$�dR=�7W��껗��k&0��Hn7|�sf�����q���/��ٖ�wO�)����Ia,�(m�:9Dd�cSE�*�Qe����xV%�Kx�xC��y�cq�guK����`�W �Њ�Õ(VRzP���YƂ�!LS����G4�2��td{�Y�=ӎ�� �D��l��N���)4^���f�݆��A�f,���F�RҬj��@�i�E�!�i��soC��l�`ޛ�uO`�3I� 1�&Ȍb�c�R�Ť7r�ˉ��{N�@��8��&ح@&֯���`��ˮ��e_�1K�wV��zu�))����pZ�Lf�;j�
h�ltjm�JѬ�n,M���.��Ji;nʡ�.��S]M�oPH.a5J7s
���eɫ��Ol�A�r�]Ɓ�En�
��Jw�If��.cS�ALĲ# �f2Z�fe�]37��m�MW�#"&��e,UaMWEU�6�;��zN<��+(�`�BD����GALJ��t��]�7,9���84�F��"��yU�qk'A�D��ԫ�-�
�B�7Y�D�ܩ/hV����{����w�^fn���fp)Q&��\��0"~��AA�^��~n����*h�x�����f&�FЕ��S��$��+.]�G�Q�JQ<w��s~�M^�dzl��\Cw^KűQ��o-J���������M��"�ɋ!�A�/\8n�Z6��dn�e���D��t�n7²��e�5�������� ��`�}囯9�a�����.�k'WMV��κ���n�d5І�I�R�U�(���責��i*$���Nl�s��*;*tr��4�L���d��?��_��$΂�3MU�&�R���� R���3�L�3o��������(ޭ���R�������;)�)�n�-.�]ѕ'=n���ow������j��so���u��.��X�vJx�1��b�{�^���{{���.���L��M]v�_b��gS[I�ޓ�:X��᠎p:6�;��npYOZe�v��Q�;�*kYۼ}[�m� 3kz
�8eu]L�g�Lj����Z�̼5
�B�t�h�l�}8���Ucz���3�S��	f!ۂ�+jDŨhm�;��I�q�s3*=ڳ:��Z²r���Vԝt�J��VocCbŤ6�K���[P�a��:0i��2�f��Vk6�©d�ח��v:S!�Ĭ��Ѡ�S�[��o���]5�v��s�l�=wGOs����z���(ְ��m�S1���h�)Yw����1�#>��nV��e�$VA U+�`��eL�ż�G]���2Cm�/d�B'f�v��[{�tme�,��D�F��ke`�Ǎg	wM�f@��ˮ��ݳ��4�cZ�ȉ��l��y�h��R6�ɑ�MB[1j٩���C�rDe�p�6!�+,��-84�l��
�t�f�N[ٕr՛0=��ugo%9o���}�6��}�K7�|�7��������<��)}���bt�Z�.�eX�֔�f���P��fЅi�3�[�W �h��8��=�.v����{��C؝�	XN�5���\U�)�fp��X����ѷ($z���ҐX+�f��h\��d;cC4�m�NT�VS.�ngK��0����܉N�v��h��,#-X���ȣk��"a�nɼ�GD�WԵTb]�38TY`�s_ƪ�+#c0��'
r�*I��.���x"o�I���Ԋ����2����M�or�}��Y�����G%u|Q[�bxj�g��\N��VWgAy�.s�����ؔ���&T[B+Ϡ�/��sz.Ƭy�:��%�Z��p:q)�q�n�g��hw[�s�U�3b��5Qט�,�)}�l;״���F1zxS�Y$�]��u��"F+q�P����{]�p��u}\�^��W+�2���IJ
<�c&r�֡�M��2��E�y,�Y�����ܺ��D[����)���2-��η)��'-j%#�����4�ɗ}]��uM�u5NӪ��]�x�e�D��d����:0����}+�n��йX�f*ʽ�u�60�h\Ո����n�ݺe(�l�3 tiQJn�f�m�j�t'���:W	�r�9�������^3�}z<��@��E)ѯl�M��L�j�P�n�;X7S��8r���eNy�a�� �@�¹ǋ�"h�^�mA���.7����j߷y^�Jhq��<�7�y� ح�Vn�u��-n�Tټ�c�i�k�n4 �a��F�U�0Z�NFb:ӳ�թ�N�e�*�7����f�L��x
��bʝ���"m[�.n��E�K9uF��]-�ޛ(�R���TR��XO��BK�M��l�˰�t��oZ��5�����XT)�԰�%�BiJl���Z���!�lV��g�di&	�0.+bI��rl\��c�2m����%�v^�B�.���Ԧ4�ٜ���Cu��;�_4j�� g$)��Gb��|5�1{��>��y��g���Ni\�Z7\7�ŉW9�hD�knh���P�������n�N��~�Sh��"��;�c����yqз�<�ٔu�/���&Ra��QX~c�0��oN�Ԕlm�(��g����e�[� .aк�q���/6�P�ز� ����cⶲ�慨R���䯪�v�u����[~!�;��r���	6���ZE8���n��b�1{�2����_E�Ն��6�0u�N���޾�{{Pu��frtiʠ\��9Z��e��S���^��5�z����j��ڇwtǨ|�iO,�/2��<ø����i|�90����Wf�u];m��g��WYCj��'V��{���v���$U9t)��b�׵�2����n���J�᜜&]^t� c,JŇ�Nr��SzEZ���:��Gg�b�[�P����
�����йE{��c�p��`U�b��f�9ٝ�NZ�Ӕ^|a�6�8ٜS�L���"��,�vSX���KY�L��2����L�Ӊ<��O4̷�w�`�u��up�(�6�O1>��m�!��`��ںt]�Y�t^�uW�v��r����`�$�Sڼ�R��'�EV���*���S�A�$�s5�p�M�.�,{���I6��oN뗴6�����TV�v���^^�D�����;�����e��u��Lĭa;���8f�h��K�V�O��(�tfU�L�.�N�N��A���̳�6vI��ve��9�
`"��u�n���y����x��};��|u]��D���}յ%%K^�+�BL2������++iRy}�V+���V:[Ser�f���"+AG�W" ��Y���!cJy�3X�m��7���p�9�0'��=�J�����F�Z���8�W��R�:L7����۳s�7���Ðr&��'n�5yQ��56�����1Gz�p�"Z��[5�36�ܫ�a�`��8�Ě!��HU�~q'م)'�o+%X�u�#CE(��[�[[��n�����o"����\����%^!�EGC�؂����w���4�p�҄���f���ʖ��ʐ���K] N^`�4�*�=���v���[�0M�`��w�]|�F��t0��nf����2Վ�*6�̼�]�YS��� �a[��˽Yv��8mYn������S����_se3�;d;j˭8;�0q&nVL]l ���k�wδ����5"�vwn�T��N�~���)�� ��R5G4���-]]�eo��4pnm[p�ٸ��C�ϻ
�yw�S5�Ж�D^F%v�Pj�I&���f�0#./�m���<)�0�9�.���H|��m�Q���\��sW]]�׃YJ�y(SD�n]��ԳQ(��
��� �Z(G���]汜�tu>��Z�g)���V˨ث�ۇ�[R�s�]�^�be�n�fBs/�������\3ssw�w�T�����l���,�R,�ؒ�ys��VDZ2n��� �HDV2BˋK$���.�&9��z�>�� VEB�)w �ve�vBtei���/�-"�go<�������S���;�0�0�T~�ٍyh	2�y��yr3�TM"����r��װ�� ���2�㐶�K�V�i�Y���(c5�6�j^5�� Ty��Զ]�0�$5w�1�.�j��u�54I9=�V�ܷ����#t�.;���R��{�-Z�O��҆`k���.�I�T�ս%�S�*��KR��<u��0���2�hb�g9x`�GB��[�"��}J�w�3z����[Y�/m>Z����Ħ����#�)�mf�ɷ�]��H���[�﷯�����	��3q��+�̹]��띳��Dkw�ϸ[�*��/w����؊�nJL�8������Vj�*�+���r��SA��;V�
9KK��eh�#'����x]t9�pb�SR��ݒ��â�@m��v�9-�BO�]���3����u����]�*�2���&l����-��b�r��VB�s��蝫��U6��R�M|Pi���w��~n����lz��ͨ�Q�����ٮ�66b �l� 
ln��m��[:_�t]�����_��[��h����5Z�;�o���͗�n�v����(GH*�6�r�]�2����ǒI.���ĨQR��!Ubn �	p[�W��)�d���Y/.��X�J����Pֲ�գ*y�n9L>�T3�d=o4(mum��G�
ܨ�=�%u+�8z�b}ռ�b�wX�l��w@q���ھC��%wcհZ.�&uq��d�W!Y�u,��[u42d�v�ZXU�)��ug`�m>}M�2K�I,Gj#N	xKMΙE�WA�fb���[��E��:��
�I�K����u��]ot�&J,'��H�v��8�/�Jw��I5u8��6�"��{1��Vy���;@Vg+#1	Gh_	.��Fg�љt��)�M	6�C��F�Sۇ��ᗆ.0�:��2���Hv��Wz��5ۏ�f�u��[�259Gn�m$V�Nr�̼bsJ�	8��o=�nqv㗛��}��U�\�>�㼹�9�XGB�Y�LM7}jD=�c��y��L����㗥�Jx��,��CQ�.��:E�Z����>k�y�h�ԷxW:軴iVo�[Wgb������k5)�I��F����jR*ܬb�����YEU�E� ��DnLn��2���3�P}Xܜ���OI*��w�|-ـ�7��1]AI7��h������/���{� 5A�w�a<ͫ�-�I�#TUpP�ꛚ1�Z9��ዧ4���t@H��ʂ�����l���Ox_Rĩ!3�
�Oη��Gs�Q�s]�i�WC��o$��.L�kk�X-�f�FX�)c�uA��6a�g��k��c�]ڲ��ֳ���3)���x,T�o&i�Hp�IvFb\�vA��{1�f�b�Z7p�Y�����JQ>�3>4������q�kZ=����;A�N�k{�҂CT�z���jwAuw����t���ٯFfr⤗7:�ި�����u�
MI�[����5�g,��� ���x�wZ��h�޼.�ެ�WPT��5 k6�N�j	�Mv��J�r;Ot��:��`L{�嬼����Rg�Օ��p��.�e��s����T���%�϶V�զ@j`�N��:�R�bGG�^_�JGE�,a���GY��u4��56nR�ogVt�K�ٳM텎NgL5���7]
��r����ܛ��qj�W���J��qA����'sܔ]��k��NJ��(Gwvn'"�I��f�tqebvv2�ɽ��M)b�<x�Ԋ����<�o}+��^�3�U/�W;t�RI�;�U����e�Oʿj��̋dq��y���;�2���#��ac]Lù�;��Sl�]urT7�mŗ� q,���6��"��^�-�a�vi��i���LoK�����W�n�W�@��VY�L=C�����':��W=�3����2�9d�-ܳ�Ub��e��r�-���N=+,��܄X��1�J���/sIË+E��T��c���yf#�x�6�0df<�b����-�Rͷˇ&�1�ƻ8�Hb�����y$��`�e����A]���RaJρ���e��������hef����L����b�6a�ax��9g<�j.��d&U�[�+&��7Tn\yTJ���$9ʅ�f�e�_Hc/���O����V�
������M,��]��F#p���-ذrL�ʥs	b�[�tnt�X���mSicW �c�ktv#��/��+.a0'�z �d��5Z� ����;n��ib�(+�,^�
ҹ�u�$�>�:ٶs���)��>8ё�˻��ך=�&m�zl��1�ynX��w�nϺ<ء��׮;\��K�-�������o��K��.7��5f�����\��q�0ۦ(���S������ա^�W�ٳ3�`�-�]ܛ<s9��VªVɀ��)��\q���W6(�	�ϱo}Q杕���DT�k�$\�4w�f��R�t�F�8�E��C�˫8m�v��N����ѳ�\O�P�b�iV��}�i9�dn���n�J���'C�.�r�<7ؕ��8��n�n�U'MD�J����.+OvM�fI�ۻ��l�|��S�ف�v'��ls�O�����zr�Ie�W���wcU����7f-�ӟl"�5��p��p
��.TХ@���;��ȥ�s�]��'#�;�	���stG7No6�IT�Mj��ܒ�*t�)��gV�t�m��"ڭ�˛;��B�rH<��6��@N����`�2mMv���+ox����ZI��|p�h�Ũ���Lt�fK���Q񽗹������,]X�.��!�Ǚle��4fZ�J ��y����f	d�gs&�HO�<�g���i8C"�9D*(��@���BlL��-A��0�cY�c��3��� � -�]�Ӏ�3����"f��"]��1 ��)mA�}� �Y����2]۳,pxt6�J�zt��q��KW�ޭ�ME(���:�	%��`VV��p����j���9JL�"��`ɥ
�Z��+r��+#����ZRg�R��ʹ��kF�[P�udS0m�0�u���Q��mA���*+*_U�9����s�ob �fV�\���ݑ�3����4�L�X`���ᴺ�g8�E}Y��8�1*��a�k6�F�p��S@��}|4p�\��S�v�k5*Izfp�0ݼv�8������@hՆ�f�ֻ��9e�L��Ԇr�Ī�y�rk��m �!�K;��V��st��7D������U�:�KU���	6t�ج��3�P۷�\���{J1���-�7��ݷ�vLT����^���ywmY�eF.����K���6�m"��t�[7Y��C�c��],7:�m!G'Z�f� ���D�>_u�aT���9$�/��_�]'s0�"~;�cS�`�F#cݶ2�еpR�ǝ<���\{7�y(3�.���ڽ�����ۋ*S
nn\�;q�����Ju��T%��!r�-�+>l�YR&&���	�9Rm�P�8��Y���m�Uש��s����;��.���7y�V�i�'v��c���so85�n6kj�&���f�)l�V���z��� Rt6	�K�X���n�Y��[��N��X!<ݜ�ږ��޴���%A�i�e��Mep�y]�hT?<B��i\[����� �꿞�Q����!r�
���^:�UD5D@5�v�}�[M15E[�"N�����I M0 )�(1d�*�HB�')���q � ĐY, ��i��B����y CH���'�$��)!!�-��$-2C�8��@�6��!�!����-�!L+U I6���Bi�)	0!l�	& ,)��a�T��	�RS$�0�z�8��!�dĖ���H!��	�
d+����Ρ��R�D6�� O2w�r������y�-�-�]��7�$ר�RBRL��b��a!L
Z0XO$�I�1$���ì��L@�
�'�@�	�C�6�M�$-$v�v��[	[�$�HI��ca�C'Ԅ�`RB�$�% m$�i�XHi ��d��!l�RACI)�t@��KB,))��RHy� c�$� �@�����)���L�L�BCL�b Sy �O!�ܒЁ��k( �A4�sT i$)���i�2���@������2�YD)��H��s�TS$:�i&0�l�^�d��2
il��q2/[!-$)�KB�$�B(d0�I�i$���L��4�ld0������ q	��@��!'U!��HI�B*����l�I'w�R�6��d&$�HBy�<�0����)���І�I�)"�:�ת3*���8��F��Kd��P9Tu3�!���	^�q�:�1 ē ���))��I$&$��Ĥ�!���	���ԑBRLf3�0d��\B[l��%�tR@)�bHy��8��VPM��!*�$�4��$6�Će@�q aII
�\�i���� �1	)��,�q�-�$�Ԥ��A��W���;�f����4�Bq��RE��)'�m��7ue!)$7�	-!�.�=�:���`K���%�6β��4�Nw�&���T�2r���^����i�α���-��1��f0���bM�'�AaHā�m ��ɂ�@Y!B��<��.J�I�8��`SIT)�2s.�Ci��ˠ4�m�^Pi-&�m�qĀ�M!�*C�ͤ�-�жm��M0�Hm-����NoV��M��E!M���7�Y6���CBE-%3���,hs}�1���W��Yid��j����Z��¤���I�7�-�*ɤ�9��P.SRS�[an:T!1&&в��}��0�ظ��\��b,'�m8�NQF4eq1���i�6�`q�]�I�
��1���g.���;o�y�É���+�Z�]!I:�s�Zm��_G��u6��9]���R��/(���7��8��|�+��P/R���c���L�y4�
=R�8�|�0v�Ku��<��5fY[���˚|���҇��S|���J|�}vq�]�Uv�6�!Hj�W��=���s7������c��*��J5�%��s.���8�C|�ӽi�k�ft��oE�풰�Mт"��" �c��3�ɯ��1Y�������i� &ւ�0Ѐ�D�b+]��J��RLQ�,�����1��B�\���J9�C뒬��u�-�Ҩ���"�1
	8`�0��!X��&�Hk�l["�L�L�e`���X���_k�۫3s,��h[�,v��)�ZN9���X�:\��<˼��&����Y����J�:B=5r���I�d���/�xB�*�v�J�JM�m�mNૃU�]D�BVH��6��L"B�3b�-��!ǎ���<����'ꓘm�8���f�;3+-	b~����-9@ki��R����@a�*���a_ "�*C� +ʬ�2�Gi����Z�`�� �ê�1��ř	]k�O�G�eu��X\|(�:��#�i��PT��>J�X.(��g��R�.p�k��}-�s.��U��摙�3c`ԼIX��n`nʇ�y*���u�v�w ��wG>��R�wwtY�ɼ82�8n�&ª��)Pf�l̀�ę���Rbv�pjGM�XM�c)���j�qm��$�n;+U�cp��b'	���&b������L�*�bB|��Kz�WO"�VPǸp՝�h�*b����)L̚���*O�j��QU�7%��[r�-7����Y����$ۏn��*Ӱv��3%�T-�[��8�w7ʳ�9�}�]��!���+H�N���u�����j�جB*�;��E�Q������+Eٱ���^-���kLeXa&��I+��T���ӛ[.Xkjnh�F9z�xK.j)EJ���Q�()&�C�h�X۸ �{�J���C�c���hk�P�r���kt^�R�X	dca]��O$pƊȌ�|8�k� �"+�l
�2h���dX�X��jP�ȥE��2�_�������+X4���iʘ�2'ғ���OR�M�B��"��V�@��O�Xv9d��w��r��Y���hE���
�Ec���8�W�:}av\�֓Vh���ޮyX��9r���۹c+o�5m6�ܻGy�yB@N�l㶳�*�Ћ*V��W�4��αLsɴlwE�6�&�w0yV�cTCW�� "cj3!d����j3s���<;xA�P�fU�Bլ{:��|li[M��f�*x���q��*�`㋶N��FQU&&����صJ4�.8w5�4l��=�L�o�H��w���Kuݛyz�y]�aF#�/n1E}�뻶K��Gpt��Vu��$+����.l����Y��a���S�¡��F.^�t�k��A�votdɨ;K�m�A������;�ޑJ�z����l���1С��񵕭Ω�*ʗ�$�P�5zo�&,�/��J�mvK��ܕwL�w:�t�3\xJ��6/�X�a�׼Ϙ2�>�-��[^�����|��{<����	Pfk]ڙg8NkYNH%Y�nm��5��a��]$W��8�!|�l����뤶£w�^Š�@bw�W7���i�,L��.vk5�5�Ȃu�v�&��o���P:\�D{��YﴸŎ´Ly�K\��ź����:�H���M�-&Sq@)hS�{
s/;�GTǑ��]�	�M��H]m[Ӌre֋ujn����oi�Ɲn8s5ӟDDD}DG��>�D��O:e�����r��.�V��Sn�>/&^��yyd��!��4�b��*�	��ì��
:w��fԎ����u�]Pi�S��su��$	<��� �$0$:��e�I����j�N�Bu���Bd�B��d!:�$Ё4��i"�9�$�$�a$�oy �Hm �Cl���w-��>ֵ���^���ǅ�{�ATb�D��QT�����`���EQaIH���V��"E"����hEEUQDT�"�0F)�)T
���r�X*,=EEDU(��EQ���O��b���JF
"�X�E*�D`���"+�`�����ʸ���X�Ax�Q�b"��0DZe**"��X�T��p�QUEU�Ĉ�`��Eb� �y�E*��EE"
F*Ȫ$DEeU*E��"���TE.��X��Q�������c��"��
ݝɃ��*q)�G�b(���QU�+q���(1ICB��QU;E1`(*�AS�P( �}��	�H�lk�Ns7��1+>��DTED���TD�R�*�V"3*R��`R0UQDb����E1oeAUE"��ԡTQ� �3�DΞ�E�� ����b ����T��%(��]Ŋ���*�TX��P�Q(��@aw,EQH�X

�b���r䴈*�|��TX��W+�%j�Q����.�������(�m(��#+��D]UN�������ʡV0�y��7rѹʐsfݛ���:PUUDSteТ�gs&(��1�������(�"�z��V"
 �`��De�j¢�i��X�
���U���$ҰE�SE:7�2""�z�6�2��:j*(�8�=ۘ�ȝ�(�Y�'��������uAm��J�" �J��"�G찵Q4��Q�R����Tb��DMV�]��
��0�oZ~���2
$y�]��ր����U;Tĭ��ɨ(���PD��!���'n�*��DA��0X[K�Yu��,y��`"���ʥ��6�S�H �����Ǝ���Je�*R��"��-T_��UUQ�9��4
""u)m���SmD��c�)T5���z�U�֪������7�)/���H0UU���QuT�jj�(�1�Y����$���a�sX\c�M�
��Ҟ����TPU^��SU�(������uH5��b���DE�j��s����PD��k9�O�������/��Ş��)X�	@�v:�s�W�t�k�������|"�ʱTUQ�JR5F�S*���P��OYCmr��A�f(*��EEQC�|f.�QV�g�?4AyUb�(���W�V�C�S415���*�Q�F*���1��!ƅ��7���]*�� �7�a-���	ɼY�/���$ǵ����̺X�z����iHj�b��8�+3��R���TASK���"��q+uWti��S]��)����]c��
QG�<]�H*,U�嘢J�fz�l��Z�������ݮ��\���>��ϊD�(TG̤k>��R�Ƅb�����{�E���,X�?2����5����Qz���������H�DU�(��z4/r��5@�Z�\)�b0v�iB��JGۻܼ��Q �`� Mn��I�MlV��ʳ��u�ƕ�����xvҝ��v�u�,UU�ϮS���M�2�(���뼠�Q�u�r�r�-�1�^��ˑT̠�W��Z�J4%�)^��S�*|���<sZb1����1n��33��.ff��j�6m��!e�	[�5�Z���q��P��i푣 ���/��eO-�ؐ���&+��{%:��t��z"���7�9��?���X�u�+^�w>�3	���3,ۨ��o�1��혭��Wc���5����z�;���i)�ڶv�`u4u)�Q��j�(��z��ڔ��)��^�uH/j�D�er�4Ц�)�����
�>�ۡT�(�[F��4u���P�T��3Z��V�AX��g���?k��kZ�c�{����(S�>�0�䧭"(:�^H�H��P��)_�d{T����ᅲ��O�E�}���e��J"��p���V�G�U����U>�����9g�H��S��G�ib�k�9{��v���r��5�����JE���Z�Z�J*:��}�j���dƓ�(!z{�u��J�Ǖ��*�TO4v���(q�Pz���{US�cBq�o�l~���_&����6�̟�@�Lێ<��^�M��d׵�G�s(>I�<�;T*v�F���C�q�߬��%�����&#q���V��*�(�ϵ�4
�C�r����UQQ�ږv��(�E�$|���?AH�@2�uG��7H���WϞ����
F��/��Q4�,�
�}\������PR���aת�U1�7Z֢("���>�^q��Z^�w�ތ~���b��3�m�)�I:�[��6MA�JZ*�b,Ԭ��vf��s�o3���9�ۜ�����Lo��{]�X���)�K�IWG�T&о�5�L�%�W��,��ǽ��"�c�
���P`����^�I�k�hTq��S�L����^]�Y�E���u��bO���3(o�>��H�(�$�D����O}�aC�s�u�%��U�u��� �����U5��h���gF��ES^�Ͱ�Չ�
Gl��V�?���W¨^�)�񥝩��k�V�}<�A����,T��S;�^JOV���]�u���юe�_�c��s{2�FG����i,X��^^�[4}T��:�t`��&u�ژ��f&X�C����oN6�vl�����UU)�)>eu)�貑i�����C�Y�wZ*��b���Z��W�s���բ��*�}�0S���Z�����AAT��{y�v���SA�;c)d�`73+4���J��^#�B���֙�-X��Tr����:�|�5��B��P���ڬ��L����^��־�j3�ZK+�d3�����q���ە[;yGwE�+R.�p}C`E��OE��EͯH�_b��c��X�xVM���Ҹv�����i�f��\U���NYm�
k�TV(�p����v�ݛή�uҕuc���k]�tv���o`�T�oU��5��H�N�W8�'�=��7��>G|��\�QH�`��e6�:��Z�EO��)h�U2�_o�iK֋󈋿�-OUW;Uu�:�Z�^��{�Ե�""�S�}��6��h��-�y�U�w�k�U���R��7��f�TQ!|&<�#�3J�/i��Af
_fv��,�*y'y����0F�٪���qU��Ֆ���n�.Qˢ�]�i��d�C�hqYt��	$}?D��}����<�B	te�Y_	Q�w���":�/��՘�Wm+�������Yw���dE^{0�ꦐ�
��`d��J*)�.�gͺ�r�ٮѝ�p��\��e�Ԯ�Mn����[�|��h���(�]��UR�_��ѩ�^���*�|I�}�dwT#|혢�w��4�WMY�ɮT6"�c�Vq���뗝�6��N� �hF��
e���Y�~��M(�QO��y�Z�FڊfU�ޫQ���z����ڜ�����p��>���X\�����G��N��g�{���M�{��Bi��l�,�*��};U�x\���QA[�KA�5H�ݬN!O����ATj��i�58�U��O7�ڊz[�w)��es��9Y}��H��i�i��\��P��ϾѤK�G2�,sW{����_4��}�Y9��"[���p�5*[B΋7)�Rf:��X �".DL���B��Kc�8��݁��J�@�"bѽ&�G��;_]j���]4�+��ո!��g�9��I���T0rq3�	�}b86MΕ��'�h̚/#יޜ�����3H�U�J�)�D�B�nj �ى���D ����|���8�D[��Ds5�6�UB�4�Mb��ݷ�Sq�9Y�u�S+-�-����MBɘ!�X[Ph��D�#��St�U>f�[MТ�t �0˓���d(��D +C���on����u�X�m���7tq]�9�u�L:�݈wj`���ܥ!u)dn-��x�J��VU��mp��0�b����k+�%i�f�]g+��y}ڐgX��f]�e�w5��k�ҳ`ʳe%n@�i
yn�@�VM�c�Ng�q��˿��CL��#`��$)?;��j�@|
�j��@���>7�k����֡�����"';v&k+z4�8���{z�Qf��_�֌��IWV�1�VlP>ˡf�ր�GJ�P|ٙ\I�����u���]�A�]�e,�ժ�\��w;Tv��u-�����b�~]ή�Y�7(/���j�&D,4�`���1@	${5a�
jy��=U��{
�.���E�u5E"�~�=Jn���m�O�� HE�I�Tomw��O�,W0���Mލa�q���}�tҬk��U���W�g�����2"D�Q�߻�٨�l�,�ic_+��k�w���D���͝�b����2���)��s�4���Z��P�5�y��WK#P�� 9��E!7DlDg@JD����[\�55�:�]�2v@�(h!&4�I��20Lcx��q��9˗ƞ�i�e���r痙ߨӺ�͙�����q+�,VQk���`:��?n2�ۊ�x��zX��߬�-�r�a�sW��6{~�;w�~^Q�X���K��+'���G�o�*��������p�B$�:i;�Ū�H0�0�}�4C���tD��-(���f��]�׉i��ݗ*���`Ъ��_{G���ްݒ��mtQ�j�3r-�~q��@I�>��)V��&h*`}.w$`2E��
��(9|��.�gL�Q��cA���G�Բ�qHD	�Q�1^�WUg]w
�p���Ǿu�Ō�i�F��ssh�T/�\3y�7��j�߫����s�Ҫ��̓^r�7�ޛ:��vE7[�Y��32���16�T"���ֳXg�<��=uڮvd�[b��%Nx�x��.e�(v��]��&�ݣ]ͬ���Ů�Y�[�/�\�6�@Ruz3jcY�9�UV�G�I7qz��f��74�*ea:mv���5�-;}f�"R3��d(.�P.+7��}v&tmX�.��1�eny/�<��x9t�ʶ�|�ך�Teg30���Le��GP����A"�P�d��%W��̭n��v�YSi��z��&咓S�ӭ?V�0 @�0�G9 ������
�>����8�1I��|�}�6j�c�]�O�վ{�W'�ڄ!����@�,���#��Z�mI(�����f|y��z�^h7��N/�~ы�������*�z�k�6""���D�+n����W~H�u���kM�U�Є̒]R��>�����R�����4]_s2g�����2e�Z(��{&'��=��Ϛ�͎�� D��*�H�H͚�<�ݖ��m���{�_�|���w�^�����3�bZ�I�z�[���s4�˼}�w��`Ę�WQ@ ���z#�����X6�b�k�Dq$n�ScKDW
�W;�'bL�LV�a��t��8�+��+2���Q�
Z��ϵeaJV�y>h"�G�kU�S�k.�m����Ku�Y�T�N�F��bZ�����������`��V���ތ���e4�Zk>>�m�k��;u�Qh.c��<�P(uN��mY�o���ڽ������sq1: )��v%?*~Z�Q��g7}9�}���d��:� i*��y�l��;/_j�b�~ߴ_q���A���qU>xt~��g�㉢ �J����d�8��%ZVØ�>�5+M������w�׺��ҥ�W�S/.����"���n���a��1������C�u��
#�^��ި���W &�q� �-�\��bbb�u��11�{�@b�cC�0#	*wf��(����~y�L�;�{��5�� ��S$��_����N�Ci1q���IL'Xy�tB�)��$� y�����^�[W��+ꄷhE ��+��X��ovI-�&Є��5rq��g���'yP������3�HN|}Up���'��;��Cl$�5 |�- �!�R�L�2C�|�m i'P�>�!�׺`��8q�]s����r!��{R���}�u�Q�X���7�wG���W�;tb�wo�%]�����r�]���dtf�����B��j���y������ZT�\�������X�f� f�W!�����EFE
�.�������Iq_�K{��ܫ���a���yE������UE����L�ö?�S51%9�'PQF@VQ���>����y�*=�۸x���@��`Q#�*���|cG֨��'I���.p#����,�$͓��͸u*�e��T*����bu�{�:>�}̧]��[�~�~�P��������u��W&a����"%��,E1��{�1�A[���3A���˦@��q�<�
�a�X��@|g�ΔrO�0����q�>��?�k�U���T �'Ig��Q�Ukxa�Q�/,��R{�a@��4i�11Z����x◛�	F�A"�������xw�n�T�M3�fS���Z]��T�}�L������2I�¨��Iy� _ۂ�j[���픬cp;N=�Ϻw1(���|�x���d��щ�eО���lX�(��dT�$E�1A��U��6v��^��
M�w����0�,2�fuݿv�=r�٫��+�������CS�� �T�n�-9!�0�8D	s�0�@���8��xӒ�:h�e�`��w�<���m�T'~�8.�7-�(ߪ�-��_/I`���xn�m���]?�X�f2�C��b5[�-D���>͊r6| R"�Vj�dK�cHU�)o�uwX�a�:��래\�7��h,r�er�Q՟3'Y_7ͻ�ϻ�����`�{⿌!d���9�` ����p�����՚�I	��`����^����>�ڄ y����ܷ��}[��n��޾� ��RBGڰ��ʼw��}���gzk��0��1����M�L�3�^6�}�o��}�ޒy�(}�����\��`�Tn�X#sfdx��^�{���NVd�޹�B5n�e��7�5L���$�ͦ�'.�ѭ��,�ME���q�}.W������k��\-���	� a��E�H�O�-yP!֌�H���4�~������@��~r����@*+j��R�.O���抎a���w-��Mܞ�1����3�R%���}��`��t�f�)�}t���޽l�G��X��Zs8%������eOF���Eی6��㐗��O��B�8Ma�`��2�!���z��;>٩S�˙Ѫ#u������u�\2��g��^���sL;��W��B�p��Ue��kE ��9`JL����˔�nDBTĨ٩��9Ue_�N�aO5\��=�m�T7y�п|�xhsA�'փ�B�<9��F)�0LA�����S?	��%H�.ᘺ��	���FO��@lOW?
���	�F'nP����`![宔x���)�v�gp+��u�:�O{xg�Q2��̘��P��p�����`ޫ���\�����0f�`/����N�%���J�<�͕ ��[�t'5/�ݢ}UC�=�6C�bf"`;���B�Ƽ=>gd���~P��b�A�`(��P%nU�pE/��l�5�J �@6.������;��	��såW��}�3Z�C�:��w�>�i��|*뾿?L��j�n�y���W�l��דg
�u-)��{Z�|�����r�]�>�0U�~.�×q�0G���.��e���-�r$��jť D�h$b=I-��H�����"f���b��_s�Q����ȾY�uu5���;��xJ��%|>������ ,�3��}@R|�aHy���=(��������vk��e_4�D@��0��!���u�G�}�4xJu�L63��0Y����)�\Q�"��Ӓzp�X��"!v5�1��~�Os����=֏�7B�I�9?Dd��~$���_q����5�K�0[�/"�͓�s�����kd�np�YYS*���Q6U���<�kA3�B�qT��Y�����[��B�o�zw�)�[��\D�n����b����.���/ώ���ͼ��q�Y[ʛ8F�.긠�[3&�/�@�N�+'H�#�D`Tn��yR!�4�'<@篏��N{vsή���J�|�ތ�ޚ�]͒�!)�]�v�m*�Ŝ(�n���GY@��Z>ϫ��C�w�`�3��¯�"\��j�H�#T��<f��j	��M������?r�o�M���T��?tc�Pf��j*bc�G�M1�}�Z|�j����oxw���uZ�ύͨ�&��d�R�'wvk�L�'��G��kU���zm����%��p	Tu��}3R�k$D����ߑא���C�_e�r�����Y�``h� 9_��� ]�$(]c��~��p�T����ů B _[�A�f��>ӳWU��뼊��S��:�_����g>�%E�w3�qH$V�*l�V�vV�;�}f���;
��D�+:�%Fc���V�,(Ь��C!�?	`���>���
@���$���ʻ*�\���^��Y�WZ7����3�@7�Z��պ�s]˯���掉"y��m%��²bcz*�BȲ��v/h��kQ�d�b�3(R��n���~24U�]9����\"����<q0ܣR~9�#�wb��^�T��������eч��sAB̪�
Cդ��Pl���3�\� �o�l�B�M�5b�hKJ����o*e��io���q�NJ����������.����:OҌDёnP�f>&��N�粨�c8��W9ٿt�N��T��@N�t|͆Lo��^��[gr�ۜ;^~̝<��S�j�<D��eJ�WM�����G�����DcFj��J�ӀG����;u:�մ�Xݮ��	������vև�B-��]m#UԺUW#@���K����Q?K�~s���w�83g3Bv���A�����f���fnT��ޝ�%�>p��V��WU��g�o��jR`1�>�a�՗���[LYc}��^��ˤ�ߵ�LO&�4�:�D����q�o��q�V ��P�����fU��`B��nR���L!�OJ"b�k
:D��Bal�DU-�>uV��`�a }����V�Y��ۍ���R������S��Gk��}�X �KV�� ������p(|0��+�<�����h��4��b�ӯ!qF:B7�K���:;LU���?o=���(�ňO޹ E'T�ň���S�14:��������q�G�R]]ӻ�m��]�f�p�������7�w�D9/&����ڊ��"v��"���fh t��&��|�IĠ�nR�Q{H����J{ܟ�PQ��,^'�x>�>���q D��r�(�T�J�&qG��ʂ�.��U�l9��*��W��(��|"1�Pq���;�# ���u8��s�B��-�^Z�+��S��1F�[0I�)
`�f�	<���n�D7����������T;�E�^+=�Q��p�>�c���e����k,g��c^O�˲g&ۭ�)�T(���*<>��S���
��)���1oO:���¦r3�8瑩�����~��ڷS?^�BI�,�)a6��eUJn��I�_Ut^]���L��Q����R��b��M(".PL�f�_m��G�������ڼ�A����g<:%��k������zsa"lҳ.�l�8�nR�2��qWIL�n�d�5����N�\�
���E[*�M2_N�����rˡ�wi��R�i���ͼ�M�����Ʒ�Gojj�nJX`E8F!` ��c��@:��Ȼsp1��@ $�*ڱAt5��^X�]��۷�ƚr�k3��b��s�D��+@�D�XɊ��a��{�y��}�p��]>|�Lf:~�<!��^�W�q.�ߔ��.��vQ:�w���۾~��WUwW�s��9�L8F_)J^=Jw`�C10�s�?
���D{M7D
��0D^ڵN���{uӳ�f��
 �%�B�@��EO��7�r� .vL�LGT+J�Z
�cDT�Aq/;
�S�Me��<x��ͫx�R���|�V��U����4�i7�dѮ��CZ���	��y��OъW8�$�܃��J��j�V���:������)�]*~v�FI�P��@�Ҿ�fY���8&f��a��/N�\ȑ ��F<H��S{ԌB�U�8TG�9�ԩ��c�۴A��S������Q�`_��	ŚkF�JZ���V{t��"{��ѽ_�NU |m�^*�h�����~�6~B��S��47�v�}��l�-����Ƶ'��	��L���mlI{f
���Oӓ�n��fw;Te�ENȼ����q$c<�]�B�D��	���}z\����s ��vb+�QS��E�~���:�댳��wH�{�m팆�Lv���LÑc�$I�w�L+�6�/�yJb/mdl-�p��r��B^��>��y�{6��ֳ�so�?$�Q����(AUD�k_������1�B�� eӗ��.��k�������fA����1��h6-W�Vu�2��BS�Ֆ/m��OB�W�!����7˳�ǒ�$e%(�/�vv|\���,J���j�%\}W4���fau��+T�M�Qt���hG�U��@��T���s��Spa~*�=���)b���\I�A��_<�a��3T�n�̊�ZK�ȇZv��_C�1Y�h"w)���Y��x%mV�:�C��X읉���3grf�������b�GoP���SݵU���ެ�OcU��<�5�q��Q��z.��nѼg�f<<�wm��c�Ql;m\؉&Y��ήAh���N�
� �	�E*�M�jQT�_F�=��WW[�m�8�R�U�Hh֠�'u&�ec������sj�-���a�]���D�P���n�Yr��ڈ����J�N��{]�-:����7�7X(YO
S�˕)k�nR�@<U���B�sd5/���Iu�Q�7�J�W^�����T I�!�財�b��()Y3�&)5�+��ᷯ��0G�84�a��i�(���*B#�V7˹U���k���+�U�������a�Y���6�V�Q<���k]��t�O�����fizk�����j�6x���M�c9]���J���{t�`�\ʾ�8��ȍZ���,c��55C�Z�lk[�Z��v���,μ֫n��c��KG�g*�Swe��y��f� �7RL(�A#b�a��a��
\͕��^;�½��
2�)��K3�Wuv:��8���w	�C�h�))(l���-vp����^R�oh������7�a� �t�/�BYh��$`�3��t�V��`�z�Vÿe��sx9� �l �!��k���޹��}D٣�-�E#ͱ*����=m�����ʒi�=��o&�`Ee�.�����2���޾{M���eH�����aS@����o<:�f�c�]+(Պ�!�Z�?2�d:�V��Q-�����&6�Nd(���ĳ:'3���%�&u��*�$��C2lc�>g�X���Bj�1764:�!3� �{�ia�/e�wn�]L���Wj�Qvv}���&_��T�u��y+�۴4Y�ےݬ��d�h�q|l�'�&���vC���ϵ���V۳��n���E�ILY����T�d�h���Xq��޻�][ٙž�vqU�GI�r��s�V���j�N�;��3�U˾y�I�ޥ�����w$�=�髷SiP<6���d�k-�,feǝ����:���!�~�諭��U����M3^�]�'��--񽩝Ŕn�3�컫1�q-�Z�&s
��իW�*)>��c6�V�:Y}P�u�X:���~�����]�O�~G�աYu�D0�p��u���w����U��tg����#ۓN�{:�)`�=?;}j�z�H�B̼�o�;o(\��>��x�*}�a[��?�>�ʁ�.a�Q21��L��1���rQ���e�Pel��Q_3Z��oW��=^���?]-N���33!�'�����	��Z?`:��L�?(�1��,�0�ș�s��4��H�W�G�,�=�]����;����=�g'f�݃�|�Qg*h�X�{�f��<S���
8�0�q�Qս��ͣj\Y0yʄ\T���oz�
=�Q��{����{�S
Y�օ��՘�+`���i^U+.�҆>��TET��r�� ���m���}q��b�j ��s�v���	^�6j���[G��9��E���.�.A���\[��B�`��D���-U(\�-��y�~�q�eC��Z
&�.���!�}i
��:װ8�m`��13�(#�(�IdD�����*]�R�L���B6��z��K�m�rdƀ<�gOMo	��H��`�z%OD���ZQ`ӱ5�U�U�e��tơ�NN�P��b��_#��t�ܧs�[�C�٫�B_K�d�b��;a׋���0O]c����T�0��T�K�=���tT-�FGx烇51û��ămpb�	mX���X���ML����5Շ�U�P�wu��V6�Md���G����1��UU ��׮ˇ������<��(I�>��&,g0gON*`I��U�@*d�(�9����f�DA��;�����b�3��#�De��Tf���#�sI�8`Fؘ�}Cg8w�[���R�WE�xaZ��,m��e� ��Z��A,4��n���v�`������-@F�"�w�C;P��bV�ST2�9����3+���]T�O��P�\p|7��0�G��>��q��s1��mQ�WwB��I��(��f3p��D��DG�Ϸ��E;�=v���(��ȃC��ȓB��H�$ɱ
`��HPx��D�׳%��e]t��@�)�^��M.����U�p�dg�����L�J��O�d��+nF�V1-:�� 	��b'>Pa����9��1p�K�s�.A:��>�yq^Ȟ66�G&g��y�B�"YJ��R�YNL���]w��Q�����"�ME8R��R�&��a�Kݣ*!�����]�y��m"6eJ#Tc�]��񅼚۵^r�Z�k���/e*`��0P�W��r0���_��<�Jk=��������:��B�y������ҿ_���_�ݐEg3| ���?�g7��X��|ٺ���7�v�F�ՁJѺj���]]��$RĄn��i`W�)U�\�*x�R%_�R׷O�Xݧǵ�m~;��
��m0=�c���L2�x­"�J�o�]Epn�T�t�W\���.Gӧ>;y��Tq~]���VL��4`�ו
(
#�eA���B&P�1C��+u3"s��Y�,�tS9G��dҖB�`[�޶�H~|�@����ߕ_��i?��l�uw�A�/� Ta��)�;�%mُ=Z�D
�ߢRR|��0��f4��90Kc����]m�C7�-�CE;���);��g�[ɶ��?�a�*oc������ �vL	�(D�� ��J�̓�h
D}�T���,3pe�d�^�,f�]U/�{Nk��*�o�b��ԱI_)[����oy��Ů���sv��]���u4^t�Q*��+#�nr�5ԉ�n��go�����dڰ��0�=�"����0#PXkCiȣ��`(��jԆ/d'�oh�La�`��-��DS�.�u�TR%ϸ�·����}�7I�0Ƴ���','��i"�F�dx)V����ӭI��}�bԉ E؋@���@���z�sÖz�.�����x�"�;�6f�f��ꄡڜC���b����9W��䝏%� C�f�}[:Ħ����0zE�̋iI�e3^�9�P��/s ���P-j��������d"��s9K�Ly�S�1�5�\���œ�.w�/�2>-�.��"5|��^��Xi��;��I���(�R;�����&b�+���=�8�����{+r��B%n���G{ݬX�O��D�_m�0���|%S7|`��"�Q��P��d(���"&`�9��z�(|�}�t������Q���B�o}�ش��jꠉ5ӿY�HA�Q11"�S��O��n��ćK|�ؽ���!0|kY��Bپ�����g�?��	#pf#6���b+(%��em��*w�������Sa|��iF����g^z;f$EK��뜨SW�=Y
~���B7AP��n@\�N	��e���'^������|\��yb�k���P����_�W�)���j���@��<����	C���K��9�T+����P�O.uw鹩�ʼs"Ϋ�)GU�<;��"����d��S���*��g������=QT #P�4(F��}�Nc��6����5�8�֝޴=p�����ٍ��xA��s3�nhA���[p	ZP�d������Ҫ ��\��"}�1�jr������+��a[(�׻d�Lۘ�@z~�uxS��z���ά-� ����M�X-/�p�����[�֭��o\g�TY�6S���h&�'~�Q8~S����S[ݠYJF����t�.{����{����m�PǤ�X��r�y�iw>PB���������Fb��U�l��K�6�9w[�[��=�]ߐs�R/M��]ڂ@����q��۩�16�s��Ń۾��4ywW�:f�E?`Sy���0"V)�.u��Ӂ	���77<�g��׊KS	y0#өG�uT��m��'2�}�}�\�fMP�Ggi���8[����=2ߧ�� {)�j+���j�>����H�+_ej��S�s��m.�K������)�£g�(�]���eT=��J.'� ��T��wM�*O�W2�Ae
�{#]D���<Q��L&>� ��4��;�2���,��^4:�w��OB!,&�ԦC%��R�1'�u=F|� 0C1�i�1�M#Q@��_! ������2�F��^�	g�,�^�z~�!����`���ϬY^����R�Rچ���s����j)������
bE>��� %�6>���?p���-�Fs���(��x�@���銒�GBH��IɅlO�{*��r��EC��B�\�s�5p�RNE�v\;���i�ȷUR����z��ё>m�t�TTH�g�R'ԥ����I�5!�R��5[X���*+�ª�m��H��r�ހ! ϝUÏV7�gzpZ^y�v��H"Y����#% ��=���2�T/gw0�U������������+��7"�C5Mr��^^V��^�c/���N�t$!p�5�f�LTy��E}�V�TR@������Iw�N혰��H�w��d╣
�?0<����������I0!��PbXh���©Qݵy�w�Kw?r��N	N�o�m���U�ފ3��-ٵ2�_C�v��d����b>��c��{fŖuۇ]����1��yxZ�%{.Û¯�-���I�Χ+zN�H�\���y��m��.�8��V>� ��By���TQ#�T�Qb�MՂ<!+E)�/�qF���d����E�D�>������J]�]���ޤ�^LUז5��:G�y����Fz�-����q5��zAv���
��11lǾV�PE޺� �=e���q���1����KsC�p��_e��!&��nR�����P��2��B?."�o-�L'� �B@EA)B�jr�v3�cճ���[��@�Z��K�9]�rm����a԰|(�v�{n�S*)��gG��D�m6 O�1s��2F@G�O�~�o<���5f�HA�zn�D�A��R.�v	��_wDYmB�;wb��v1��#*&*ʫ#�S�U  ��0�j���h���"l��)���6��TE�p���:�h��F�����(��+��BٙbU^R}q��w�2Q�Q(�p��4@�>��J:I�&�g�^gWu�nEz6�	�n���c�O�:�1h#��͵f#=I\t�@�J{7���"c�p�X��n!��S{q~�%
5-ع���gz�9�+]l��#��W�dm��
Jb�0}�/nb���Y������a:K���ۦ��:=�����9����q/@2XW�-���zv��?��ߪ���g��Y	}S�w-g�qr�$|�|��K��������#�i0jc/��{��Hy���}0[��O�B~V�T�=r��9�����HLwF8O�*
zQ�
��w1�r$U���X��ft���vy''��ȏ\d�B�9A����v'���:�99���k5aw&
�̀v�`�3�_u�@�*�X�V��Mܪ�w���{{�ŕ���;;��[��!��Rn�>L��5�|�ַi<�ɂ�.����sq���J��{1�=�=�
z�b�Q\�UIG]��oLP��5���%��f(c��Ƃ R��O�C�6|@nzd���㶌`#W%	�l�K�����~H��c/z�_W�D	9�����>��x��qD�;A��A(�[��6Ջ�*���v�^�n���6�"s��I�"W_�A��0`B'r��sH�#B����H��?+�G�1t<��(�8�U�>�D��Iɭƞ.�ѻ�͠*`[��?G}�����_8:��?"w#
�I'S���`̒М�S�v��$ �?�3kjS��&⻻lx�~$d �ۆʹY�f3���p����\�
��V+<6�^���DG1�|�Q�M{8c�B�����?0�ѪQ3H�����rMɎ�A�6�%V��Z�}���������u�l>��  �H�O\2�i�0g	غ�	`}�T5v�U~9�R�	�~f&�6X3�/;����%䓞��?]����bEO���0�ϯ���F��b��bq@�P��U�m�̻�0L)������E
��mT_8ޘF=V�ن�~��D�<�N@���5R`�B"a�U@����*�h}RbT��#K�2�E"c{+��~���b��J����l�1]��,ue��~���@�`�7mG��M�+�W�R��y�o|�NL񺻡p^S1�h�-�9FBZ������~��F�z�]�g��㍅���O6�̹�����@3r�Ǘ���w+�Z�cz~Ԡ�� �7؛��D��0a^{5��B�靘�ʎ#~= ����p�����
�7p�۟%e*PZ���o�K�lҾ
��v5��]*q���<Y
ͨ�i��K�m��oP[n&��:+�/5A�Г�*,��:��F������}�t��R��"h]����vv��6�촋���^�{��-���r�<�� Y�I�	]|���[T�*��g`���U�a�I^�P���P��{]��~�yz�_��|a>~g���[<�� �F�̚<a{�ۧgb��������{D���% �o�Ec|z�]-�j}��Z{~Yӳ��ǵA�%H��1uiEkǳF����r^��08{���|f,ć�
��jH���"w}���q��/ۈ��G=�?Px�{ʝ�n����3�,�w�Ut ���U�ϯ�G��#jG�?Kub�BQ��DR�J'�9D�>���A�@ylO��O=8&��軫��G���+Q�#،S�@A�K5T �^*���gT勶�E}��=�����~��x��W4~?���NÃs�B�i��թ�P�����H#F��Wp�zi�i26�;�s/B���}":OJ����x&��f�;�0�(�J�����!Dϒ��n;o�& ~ޓq�@����5�h�5�����X�� C�5[�`����i
�f�js� s�G+�낹Ӄ˹^d�]�=IA��@�w�R�)�'ڢ6j,�-����tT�ɿJ�-� ~�m�S��~Ź���R �'=U޻�k���[p�~[�jn�ipq"gʻ�\{v<���^yT��b�q6͝�5��w�l�I��;`r�sJȼ�t�����/ո�r���=Q1jm4	����]���ok�!ް�1=a�z��y����#V���j�Wos4AM�C���U6�R��J�,�Ҫ2��FTn/�ͷ;{�F���ټj�Ӗ�<MR������u�����8��8�s��e��\\��F��6o��#�{b�E+wP��w�36P����v��(3C{7���,�k5���/�u���4Ɨ��n��o���~8;�/�@��n^W��M����ɫw�L�������{�����׾��3,~a*����/����F	�O����T�\e'���
�8�zָ�`O�(�*	��z�5��$ɉ���W�i
G:���뭷�&����Xȕ�vd���й(V�%�)����^�>��8_mՉ��p� ���m�	��9���W��i�l>7
i�y�-uJ��:�b�}��k��;cC������[-�[2&��P��Ph����'^�L�w�瓷U}�	R�@dx��,�>�UJy��n,����?)Ѿ��y�	̗����wq{@Q_z�kۣ�\�g>4*Fӌ1^꽃#��{<�l�f�Vz�A��s���I�ʇƐ��B�XVno9��>j'#��ԣH�@�˵pgn��q�tJcf���
����/5Ǣ��M<�n��n�LI=8�@9ҧAT���"�\o��ΰ�Ѓ K���1�g�U$�t�x@�Q�����Y.�M���������W��}p���|Y�[W^�q=�#�Z�f�Y ����sҢND�)�̏��H��݂��ϕ.�/1>Y��5�m,+��_L�(��x��cj�le�l���m\�(t�GQf�����Ƣ�b���-�e=��͂�-���ñS7K�u}k�vU�6�6h����*�
����ZƮ`�=�C�<o�KqPj>@�����=B�����JV˴�B���ѥ�Uy����Y�w׫,Y���M7�6���kT�2�ܿ�N,��v��=[(�09b��"��w�TU���Cܻ�K��SiI����R����;[K��ռ[�8ñea��W^�ʶ�6��CP�f�'j��]�9�a�\��к8z%@�Ps��qqrA1�f����Q��^UL�<��"�ђv����d;_��}}�.f��%��Q�5�z��8n����!�Nj��ayb,w�Zf`��1PÙf9�*�����v}���w]^���H�|�S	�ɪ7'�د�(ϥB*&��!uWX���3��h�� �<�FY�*�YTk�^�@��#��}Q�;�^�AV(u��+8����1eM�?yR�31DG�.��HQ�vx��jx���-��f�{�7��>�u���LUߢ�(>��FE�f)���"T�^n(a��'��ߕ!V������#7�j����*ݹ/��\���s�'m騦8{*�ma��;=��1�R���:�~�>�I�L��ٗ��{���!�x�@S��؎��]��9�qC\wkK���A��m�S׉���W��/�h��#�l�L�=ތJ�X�z����%��^(
��q����9X��ކ-O!�����v'����2�(Y��oDqh+"�(��ؔ-"��4aeb��{�����-F"��E�k��{�0gy�K"����=��z/�j�S k�?T�U����m-l*�X��>��yitV��qb�N9��>S��=SgQ�Gjxt2{���X$V�� ���{L.t���M�Ӡ���Y��~�._�!v�ژ��Cd��ݨ�e�`�>	�m��}��"4i����U�UԼ����]�;я;,`�+hΥ[,%Z��Q#9��N�Nw6>�㠮֭��\��֝���Jڵ����^nНy�Y�쨩iF�}ԵV���a\���A|76�N�"���^�Q�!�!}]���[Yu��'��F��q��L�j�
��U�Qn45%}�Q�`���EEF_+����y��U�d�����B�Rݹ��A�=��O,u��D[p+3�_I�͛�R�A��Q�K�5�<fz���T4�gI�W����~�J_�˴=0e_e����ꚫ����dt8� �_:vEuzj��}��&ip�5[l�u��h�(M ��L��<�[��NH�0�10�;�[��!��.�\�v/�������u�b�L�O![�G���b��Hɺ¶d��z.Z�\���ь��8y�s_���2��>�� J2*1Nh��_�.�$rL���ē�_Ε��tt�ú���q����E�#����h�{)`X��lNr� �B��?����zC����yߡ�-�4���7��M��HY��A�=���O��a;�#Cz���Cv�E�*�]�b��c��`��b�5�t��J�n;����8��9cB�����I7\=�mg���ޥ��:UBU9��j�Ľ��_���c����Eʺ-��I��P��j�dR��cqǾ=k����˩�H��Jꪼ"����P(��q���WR:�=y=��gJxlנ�ۼ'k�	����B�]gf} *�I@�mz�	M���0�dK�2乿ùz�v�"=���Q����f�nE�p�;�q�+3we����,*�V�}2���خ�nf�㫥�+}�=��ҽ�49�n#%���|����'�&���^Ԗ�X$&�P����OК�׍��na88����1̂�wS{��� �^��]w���>���c+>��}_W�~��X�P�ɂnd)�-Å��a���ٱ�{�9N+&ټHb����ة
���b��e�[�z�л�SzAJb�n
�BoX\���6��׵1)ݭ����\��r����*�w�D��J���g#f����'��[�­q�z��X��,c�/�Z{�\EnU4�~�Ԩ����\G<WLQ[y3�iE�z�9�1z����KEŵ5
��a=(�,�N�,y(�nYW[����Z��n4ګ؀ؒ�B��;@ˠ���Z쬹|�6���!鲚6M��]��{�� ^4�j�	�2@]x	��tR;!�z/�Y:[��+�-�6�Cjf�%����)�����{�nh·&R��CSv��#��%������स�u�8�.�Y�9��oWpnf�1]���Z��-�e���6�d�Dm�Ťs?M	A2�q��&f�.��vc�N��MUXHi�]�m[
t��@���h-/;��{����a��P��0�*���#P�v!u�4]���:mɵ�91���MH�l�Pu_V+7B7���ĺ'>�9�J��q��;t���BED[[Ȝ�wM"�%Pc���� (T�;;��\����e�U刯�pZ���8��P	5v	�k�Ld+�wF���;Q���x⺽S�Q3r�E�/[�9xl�7z��9ND�Fu-Fل w�*E�q� �*y�J�p0��=�(��]O�����SF!�i�gS�'���.\���´�i�D˃bΡ�������8��Y
�F���ī1�`e�f����tc+�eXzƙ5i��l9z��βD�"&S*r[�ͫ��&���S���wR���<'.���F/&���֦�K����[w�5Ž�BL֎e3$�f�RUZ�7T�_��x��V_���9K3��Q�\�F�[!���_���ճ���n��p�ȮiZ�3�}ټ䥽��WO/CYX�NQ����yM,�T��ᶯ%X�K�f]Յ:�Dx����ݮ��M�����!p�W=ݞn�(��{`��O�Wm��;��݇	<�#eBe6+I[���)��
t��p���d�ކ��]�G]��v�쫠EEW-s�
��;Ugf��[̕L؄ʋp�R�V)oMxt�*��9�4�۾�+u]�ݽ|U;�W���vɬ����a��r�yj9v�p��3\��:�![6S��6�zj:��u�J��}�	C�Z[u���j{�cg��eœ��bX�^"���V#�YGq��.��%�;��nu�Ņ��q9-3��xg0O���oKo�#��#����_apz^�Uer�2�|A�d��u�^ѷֲ����QUUU}�������1v�\��	��i�HI���a���ӷe%��Z/����,���aW^ޭ9g9������wx�q�x��jќ}�+�'�ݔ�0|��(��$����5�{Q�Z��O�4�[�Ux�&Ί���`p��o�^{yl�ٺ���1��m
�/�&Ԍ�+�$�Ȟw�V'���2=9�Qs�Z��0��tҘ�b��R��b]�^�7���M/�P�LM(�LShI��gM۳�"�+��x*Σ2��.f�d�.��@��G�c�I1K*�ݘ�����΅4U�4�BjWK��З/�Єϲ��Ո�Mr�M�1W~�v��b�?,�=�Q��ӫ�^߮��7���Zكp��վ�9�Ps�"��_n,8b��Z�v�=�RX��~�&
	�E߮����E����c�������;�5I��0@q�מ�.��Y����>��!U	�D;P�Ɨ�t�����^�c��s�7-�j;�r*9����3�U��v]&E�H"�P!��t'!F-�D,������p=>N^���k�q���@]c�W��Q&VG�ޭ��+ޖd�Uۡ�=)�M�,t1�	M�!��^��[a�0�dL)\=uH���Sb)A��2as��}u]I9����yȽ�z�!Ha�Qq�z�zvjZkٕ�Q  ��L��[^�fP(U�~��ʧ�A9�\�+t�.7L��K*�}�J�8�:��'�h�Uّ0Di�6R%�b��{7��_�a��~0s��\,@���I������j[�ȱJb�Ìs�ȸ�B2� �K��tiQC�ٱ&�N�#u�n��X���l�3hԑĎ��CDВ�GW���G{t<]*Y"�w/Ms�+ ���F8���yI\3�����x\.�B��;x�%aڨ;�η7���E��p��CW�sʎ��@�����o��A��EP
��L`�/��C��=�ә�˥��Y���+�B�ۀ�R�`����w�@T�M�`m�Ne�]%&&j�3����s��c$��wW��W{��F�M1�!�y2f3��!1S"t����c�;�^2U@�ܫ��SL)�1~��~�:���.�n�ox�ʍ��>�&�`�c�WAZx�VƂ��&�uEؼ�1Eco��lj�/�80:2+�ϒ�M�î�w������I���~;�B�t��P��2�[�X�8��Pzu`h2�K��B�z��!��<G�b��q�E��^ɬR��`���r�����S��H9���w��q�v��p�1�ރ7厩���tN@ЧP�]h3�O����?(͜^��dM(ay�����5����Z��s��X0/�&l�Q�K���)Q�nl���1��Td+n�X��^��|aWeH򋫨���'�Qn�,({�#"���<������˺v�N��6=�7�ҋ���-s3PMFf1�NA��W��*�G���G]�������V��F�Ê�4��>f�c��:��]m�Z�H�A^�|�N�wMݷ�Ӏ�neg�9��{�ǔ"��o}���;&���\��:���2	^Q�Eg�J�a\ney��Mi��k^a<�wM��,TRl1�0�ȩ��tUa���������g�۱��h�2wQn��	XJ�cH��r�n�),f�j�F�Gp��R��q��w��5���E��ν^X����Ռ�rPI�&�D�1�n�J,W��R�q���n~�}�׮ﵟ#m������J͞~��Y���J��ڙ#4)����4������5$xɎ�˧{��{-�g�:<��KͰ���+�����9�NX�P������`mr�86o�~y�Ƭ����2�S�D��0v3�6:A��T���>:���I�����y���H�"�s�����Q����1R�+�8q�*u���r�Q�֯*p_z]�6�܄=��z&l�7�M�˒�}�1~�|��U��G\�Eq����c�z���B*q����	q��H�i����cIY���z�B��r�jө�yBx"��I�ku?-7�r�|�>�+þJ��t���F!b��*!D�C����k1m��lؿе���۴�~�� ী��_
WM�G��.�Q1��>����QUТ�^su�_�`m�&L߳�".w�%�����̲���_a�@;<�-lu�m����)$�GD������(���sj=Gf1��z<�ؘ>Rz�F�H��F����k���~b���Mc�����E�/D��U��&k�,�ǘ&�Ѓ�L�\L ��P}d��3&��{*��x\9��c���H�>�=��(�l�'���c�5T�#�r���2�K�89�L��:�ҋ�a3h��I7(��)���!���ݧ�8��ܤ_.t�{�ݎ���[/n�@F��u$�ʛR-�c2m��]lP::�aP1υn)JgX�e�Q��*�C�\M��7���c��C[���ٜgf���7?c�>��+����� �6b����^]���bW���������<r/B��f[��z�b&�U�b}u�W�)�>7�iO�K����R��c�s9�K:����������^��ut�z�^��P]O���tc�����q'���oA�y�U�4On�8��vO�:bԒv��^'��GxL���4��݌�̓%1	�Y�E����a��[u�ʤF/M�ˬ��B|(�?~�P��s�u�)��S�����V+�g�.M�b��w�F�O��-ڭbb���-H9"�A�N5�Ķ��z3�f�5ֺƏ-��z,��gAѷF�+�_S����oR��\�HbM���3
6@�+�x3]+eo�S���^�4
�p�}���L���5�62m8�{:&#�z%�eL��[w7�$� ��7U{���{"(&���}S�M�ۂ�yɹ���W~�u�*���g�&9T�qK�m:�EF;����|U�ɚ���E���*�����19�[�B_�����$����ݟ^��Gt�_��xT��(^>�D���� �^ɍG�[-�>���7�.)/H��)-h�UOED�^ΪL��3��B0���9���R�k����2��q3s^���H�N�7+)��x^w3;�WQ�8�yq'�$���u\�[��U�q��A�6q���d�6-���e���wVֱ���
��t׶��m�����(����C�Xyx�w�V$w,0N�2�0��Q����0���$���nh�w��Y67x�&�%�T��&����P�3���D�����.c<w7/�g*Wc#�k�W�B^P�	��0;}�I�U	�I#wW�뉯/�6���c�����q��N~W��<eqFn}������%]�b��^���9��;��S���n�=�2y���u���M���[��E+;I�y��y0ZX�v�o��MR(�c�ʎ"��>CE@yH�\\�`�)��nn9�$���Z�!*\�N��꣭��YRW��s�`�/ٛ�N��K-�� ��v-��X��,`�)���"�#��)G�� >�V�i_><��W��Sy�Uz���j���,Q�Ez����|�]uᵊ�le�@��Od� ��|�u�؞�j�7YV��3�k<nx��|�E�{��P��0�;`u*��z;�2�Ϥ�o(V�aK_NE�q��p�>o7����y==�����Z7Hm��"Oi�eb����{;u	=�M^��otT�%�J|T,z6����U��WI�-`����o��M\7OM������+1���Þ�u�V��(d�����^�LnVxi���͋P�"����x+'u�F�̋�Q��P$r��box$�nn��F篪8���+����PF����!�(;{D-2��f�V�EܩMN�'�xR�a��k�U�t�Ө~����A����y���s-�]f-j%�3wZ�X�*�s��d�Sz@�d)g�i�Go㑱O��ڸ�z����ռС�c�uŒ].�V�j?ff�s����n}�|�=�:�x_���vU�Q�T�ܴPr���ع�U���Ü>^Z>u�;��q��/������]ԷЊ���A{j�{����"�GEMF��ΥG����~�����^��f�*f��CHw��c��d��iLg��k˵yX���8&)hOn���#fA��7����H��du�����Eo�_�ƛ�q�3 ΀�DJ>����!��z�J$���J���=�8-�Q;aL�����Fҵ��M�#�]P���`y������V�oF��?���t6y�P��v�Hؘ��b&��{�jt���[��o�y�^��������U
�7}(�@~̫��b�ǯ�#,�g�w�wvIJ�2w0��}����MQ�zfT��y�#4�p�fY����M��)����-�U��{�����qfw+C�R/�f�L��g��̻.�3��nX��o��'(���N7��k���k�����?%��^�e���W<�$����Y	��ʗ��.�;��d���=w�V�=ܰ�iq��l��4��>�&q�y�[�aι�䄢P�����[&�pە1�&0/�:��z����h��(�'��%ѕg���3fq�ʇ��U
��p���Tu���vSp�ݤ���C�h�jC��]�Ɏ+�d=O8^�p)PX����ΩȗL���X�4��̤�P��O6팫����C�yWJ'״�]{U��پ���e'��$���yXX��9��DV�{
��&uݭ�̈́D��{�1�/�A&��Y����ǲ,�]i��j'�M��"�X�Ķ|�;#yN^�֘�ݷ���֜Qg��xV7�h�}H��(��Hev�p������rs>�rJ\��T�e4M�@�/vaצ�M����//�r&�9�E����l��FCӕ:+�h5����+�M�R�~�к���Nm��+��^�v����p����y��X!{�������z�
#'���c��iE}�q���3ʯ/i�b6�0�Y�1>��� 6{�����˾��>�4>ޝ�9@��9�D����E�䡎����W@�ᚵ�_��}�H��e@��"?mN�+���l^f֛�6�Q�ۋpz���K;����j��=�)�M��Z��6e橉�]_{��>���騵��3�+M�P�D^k�;U}쌨0�h���qpFr���]�v�O��9�K~�%�{�L�x�CͅS�D�@j'�Ly�U�l�|a��A����
�}i�(N�ò�M�2�b��|zr&�P]1��� �6��a�V{�-�:!�~4�3�f.���R����#�\��� X����ɜ76���55���x��	ف�w5�
�9F�4Y�����gȈ�*bk�m�H[i�G�@6L\�z5�Vb]g���9��� \KH��cv�m�3e�92Z#���`Z ��&Yr�k{�иP��Y9�]a
�a���=��L��Ϣi�Vt/<�tU}�r|�|���c�X�2A�l)Ӷ�7���Z��}�)�2=�0��b�*.�`����<���=rUE{s ��B`����v+�k��7�o<�_]�Gec��F�>��G��[b���z��X�I�;
==cӻav��c��D�6�\xA��q�Z~)�i��m1��qϥ�Q�����	F�6��wo~À�pZYiyԣ����H�����zE��1�65"��=�͑�ҡl��#�bq�sY�6��!�����-e��9�Z�x.Y�:􉯏zҨ��G�?f;Ϥ�l�
o����j<	�ZmC;��]Gd3�ن��]��ǝ�����#����@��U���,����pb"���ިh��xex�r��Nϫ���ϼ}���븨�c���K�Y]��f�Gu������ga����Lg��XS�/VE~3�:�*�����c�Q?���mk}uVm����Q�e<U%�K�٢���Y+�F��.���%��=¡��Q[�̸�t�����P<�Ωp��P��S��c�Yg�I�K2%�{��_�ħsE�����Rr�߭m_mȥ-3�g�����N�guz�k����x#��	�l�%�Ѕ�udng�}"j�ʘC���zn)��X̐R!��ُ���q3gV��R��,kl�Ew]�ƧB���Tݴ댃�8j�G�)g�7.����ND:�큘�WI�{����d2�48��c�6��sp���˳/��'p1˕;���~N��7�d����t�}�p�iF�F�ZLc��.2�n�OS��vt�j'���W}�/v��э-|�R�k�a 5臙Пj�o>�U����2]z��q��{樠�p7WX�٨6�	��'<��S���5Ҕu 񠟥D��:���}2���qa�َ��S���3��6��,�ۂ7��e��Ƌ~�sl���b]��`��<�蔋��
�������zf�י�3��e���u�~p�g�rW�i��ƨ���p��u�2�iZ�˞�żG�ة��)���rv+k^Ej���u�_q��%)'��������&��ވ/Z�A�Hn���S6�E�]�e�F�����Et�q���%��mu��rT#��p�L��Ǌ��f�)���+���_�>� ���Q��5׺;�:Q�Tx���	��z�+��͋V�bf;�ُ�Uپ.aE+�1��
I��5h���w���TM8eX��|�p�uȰ콦�~4
���~Ӣ�e�[�H��^���i}�>�}ѐ���n-KP^�'�g��]��]<�y�9�|����+��|�N��K�>�������7�̗_ �_.�p��6T�9�1՗IZ;M�ﲐqm!a�֙��&�����ζ�o3Sa��ev٦�ڷ��]���.f'Y�3��Rכpux�W+=�*��oL�u�.�C���>Mx<���^T��i;��l�H!X���n��G%eɃ��Xv)��[�ʷ\u/t�
��NV!|֟n&�f�z�*�\�k�WQ��um]��sx<��<�2eƒ��Tpdu�iQzzm�p�.�y�0�..8���5��\�,we bg��se0��|�P{��~u�z6���W����Y�x���\~�����v�ӻEut
�ϋ��{&`�#6{�#�ޫzz�6uo�݉N@#ɿ�	��������/)4c0����5�7)d�"��w�	��� 9n�q9��5=W�<�3~u9w襴=iM�p5ug3@�<#�u�@VL�YP��D ��������L�Z{c�'��y�y�y΅�]��>�4��>�Sro�V�§Q]�Y���4GT0��P��ʽ���;�\j[�����,��{rګj)�{۷2��m<"�w����/�/Roa	�+��c���1�߆��T���Y�����z��R�%�r�������EU߅Gj��w�-���&3�gS��~�h۬��9��9R�[Ƣ�W�L ����CH8&ӝ���>F�FJ��ڍ0���u�s�F��Qx߽y�߲}�!�4'��8N�"��L���v2�$��7�pPħw��n�u��5}hk��@22pWO-��F]/�ܙW�3xL�rwA�#W�gl( If�^\�BJ�r,�
�����f�+��3�����ݘ�P�y�9��1n���lЎt�:J�{���q�s;&8�d�fkѬ�nJ�͜�v�P����1�(�u��'*,���oi;WF�������#��՞�_�9�f3	�0ewfy3��!��3���@"���$.�5�XM�8^��x�æ�ܢ--V.������XBN�M�i�E��ʺ���D�F�ܸ��_fa��f�XЌ�$�
��'n��f��]�K��a׵��g�.�5j﯐�K�em{�]]��V��m^�l����.'��ʃs�ejo/�/u3z���U��˹�^p�����5�R���+)H�a�#�{�1�B�3�"|����ju��2��O����1�ƹ9�l�������Z���s~��s�q���w��b��D�O/,�w����uj�b���}�>wWѺ�R���j���6�`Z]?������wB88�J�ȧ�k
7)u�}�8�<�U�
��f���FՎV+��P�V���N�^ĥ �#^��$+kM�F��(��oR��)Е�0����NtW��f���K�����)��cOhU��Ad$�wF�M��� \2�gy5�i�j�|���Ts��:�w�հ=6�+;A�����)޶�2gK����EM�9����!PnL�̹Lr��t��� q�ʺdF�q�e蛐��[R����=�u����0�K�>�*h��N�ӆ�<}}{�Hi��j�T&�ܦ�N,�8@�v��Jn5#�T�MѮ܋��m����!/(V�����Z����,��Q2V��@K��������NR�:ի2����ɓv��"u�κ�j���W��Ў��r��i��Ϝ;/��\�i���ͱ(U�ՐX*�l���C,{��yw�N�,�����1�{�yZ�D�jVU���_h|53v0�۽]�/��l�)}/�]"�.Q�f�-W���A��	H���0�I�ҏ����&S]�S��[���4iٕ��x�EgR�@�D%>�e�B��,}S0o%Aۭ2�k���5S��Ɍ �a��V��T�&�B.��:)���6��](�����%Z��^��]�V��t��|h�1������j:�6R�s�]�H­۫f��(��8LI�s�mU��9��"�դ%���ffL��Aqsc�*����'X�y�N��R8خ4�O_iY�gt����M� ,�b��g³>DY�sY2��yån�+�TG]!oM51�o1�o�;��M]ۋQ�A÷ؕ�x�0�R��7MgF���'H�is�NsvS@ȻE3��yRs��K�%�!��+���������d������&E^�\�GtV.Fު�v��RLl�hw]�>�,vegeus�6��h�Av�v�gB�@���������R�-Q�g4��}DGۇ�J��\��g�ž�kM�&E�ssU;���"�de*��+Vnܜ�A�Xf�^6�fQ2
*�2�n[�Y~/��/ב�� ���d�+�!�>Ne�_J�ܺ��e�Q��˒�G3�|X�pf�>S����Wh�/I�u< a���9�����~�]cfN�����|c��IKv7���r E�����i=��`�����V�{zfg�1�4����<�\z�^�:�w�2*�3o�C�����w�_�l�W�z9+U���M+��������+��n.�F�7F����dz���L�g`q�ˣd�$V����a^<h�O����(z6�FQ��O�*��x_ȳ]�����c9�A�3��N)d�cS��Ѯ�1����ߏ��f���_�cv���m:�X�pW��aޯ;��XmWJ�#㣙�{�H���i��T��\c��Xň�T3<�Wz�:/^�3���p*���� t\QR}\�_�OW��ؐZ�w��y*?~��Þ��C�.6}�z���M����U��~���%&�A���>k�/q�~�{_�{���tcs��Fy���!F������5��oH�:TO�����ڄH��W�
H�Z�z�}�ؾ�W�6�4O;���Rk=ocX|�q,��̈́nes���_����|��{b熮��ұX�{f�`mG��r������]7�0D/j-Tl��`�7���J��}�m���Y�Y�Ndk�8��0o"�%]E��szmq��%t��23�C�A�5��|B����!�8�e������8�,ޯ߷=���ͳ����~}D��>�, �ajz��3�:�ј�BP;&���^�F�4Vn�����G3���6Dz�����P��d���wDi��X��1Oʢ��b~�.*2���7���띛Wү|{`NMI��ahx�8�	k�C*�T�2�d���>~�W�����aۂVD��#�}*؀9G�ڿu�N�EW��aˮ=t,�ybJ2��B͉�E57��w� r#�E�zG�]R�)����g�a?1'4��'2~�7V35����mxx�h_�����L����
)v�g��)��q/M�_��b�h��!�4$׌��+�*۞�Tz�u���s|(���m�q7g�mD�ϼ�X�/WtV���iU��b~�6��ӸE'�@)�����e3���� ױ��}]��,�:mG_��ۅ�pW쀣ң��=繞��Z9�P�,z	K#nhI��Vj���{mc����(&�tD�+�8M^w���~�WY EP�	��i�^�Q6\9.���9=����c�ޖ0S�6'>;J�Y}��uz�a�~��c��U�5b���ӭ.2�z�� �)���WF]*"_cRwl�{�g�P�]k�]��t��@�����)�m�����O��8� ��[u��\��e�i�V�Rc��&��%���I���u�z�K=v#�N*���8��l����X�u悺�y�J�;������z�QQs4�ՏjT�$d��8��ݥ�
���ڧ��4�ȾpR�<��u*�����h+�i��'
�$/���	�;��鱕Q�=y���j&��]O��B^����<��#�v`�'�n�Tz;���wo�����^^0��;�V����VC�s��������{�2���@��O]ӻ����h�-��x��q޺��I��D���&D�wpS�&iK�X/ۃ�.�m�L�`n{�RXv�#j׈���}G�����#�^Q1D�
0�����9U�����%_�u����6����4r��{^o
Ѿ�^�}��x��ǳa�B�Sl�N,t���yn��/�������/���.a
A!+���3�k�q�Hp0l�͘FLu��1%
�Hw}g�T�h��T��19��������V���%�Ĵ�W������a����rD�^��zJ����zo5X���V���<��4'�q����Ck���"��|�庫�ݩ�窺[g�slI��n��!��kTVL@���e͓��'5���Ȏ�y�r6�p��b�4z��\}����	3��7b����?}F]��v�ͮ�(��v��]�j��Q�eo�W*�îk<uJLW-�;뻘�;/��Y�d]R���}Ͷlr���*��ͷ��vN˗�Ok���f�*�-r�m��k����S�E���c����lTfñb���qDq���5�@/\����(Y�����OlA����2I�Х��'��m��]ޗ"��$�g�
�o���6
�3��&=�>�j@��:}q����7�3�3{P��~M[]�8�U��T/��X�ȅ�N1�܅�M�"�rz�B����Ͼ��ώQ��5-�N�F/K�Wsha�
ν�ap����L�u>������;��72��7(�ر�v*my$wG���g��]�1DQ�c1ٕsz���<7�ׇ���:�@�*��H�
!��]k���w^s�;��o��ވ���kj�v;ײ`�t<��k�\N�A�T������/<qZX"�[�]����v<�7�B�t������c��\:�w�'MЗ����"Ƨp�����T�5n�ܞ�h�Ӽ�r�T	�4�"D�}�F�n9����!������҉�ӝ�BH1��`�زA�*���>��J�!y��x��N�}�G�6�[����\�`2L�)^�b����W����A�heMm3Y�g�^�8I����1iV�'�9=��P@Ke̹��"V�e\�0ј7}r�>m�<�&äs<\�!����c�kMd<^a1S�����Ǔ��pԽK�M��n�"�Y�}|_[�B�nfov:Gb�1���OQ��2�+��#;�Vm*Y�ts��L��G׺ws��ͪ2\�m����췏o~��rZN��.ə��ې�;��(���C�	�=�b#�5�dj\��z��~�����.}86l�/'��^Z��ӫ�+B�jÊW�V�?�J-	=s/Ʃ��:0�p�_S��x��ѫ�zs�z'���Oz�Z�S��ΐZ�{>����@��z��꞉I�HM��p����Z�ёt{P5�?��5m��'��{����V�nЛlBs��+v����`�V�Y��
��ӕ�O(+�H\vo�n�P��y���;�;r�M�WM���OXHF��y�^ik
����y11�q�� �uG�T�.}1u��������Fϕ7W�x��i<��'>�lj5!S*�;Gz}b2�ڊP8���
�-9�W|�S�*|W�p�vP� t�&���n��R"�����t`�#'��NME��%�����cyC|:l@�%)N���2Q����ˊ�9�H�n��{��=���ۑԤ��2m{r���>P|��
��ߦ_3��^8|҆�{����n~Y�P�o�B/=��y/�=v�8�����ק���9�uq;�WP����{�t���98�|Jt�U1@�|Фb�k�������B�!y�~�'�
�~�U��,��߸����A��?M}Q8'u��mڰ,�k�}�����;)��M�K�N���Ú�u�"�<,w?�.��]�|-��m��{�3��;ږ���E�/.W�L�43����
*u���s����]���M��{�w^���^L�nv�����BY�,h�����9�M�1�b�z�+���a��W+<��1^�N�v��]��:mϳASZG��v4�C���TV���(׫=����W��#v��ߪs�E���d�|$��_�G���x	�W٘� ��a��`%pi�~`�<�������Py�Oq�@��۝YQ�xO��>/��uHsѥF���Qש��17�;�(8*+_��^�Wcg|n�����F���MX#��������n���j���؃�Y0�]�G��J[����Eg�բ���]'�Uw��U�췺}N��A�tX��NϤ/{�Q�{U=n�/��~��y�Q���������9�3�Lc���uXb�Yx�����w||�N�Q���A�P=��
�F������,jGDﵷ|₼��U�7v��;� L�]�
'-[3.�'#��&���'�<��[��+���Y�Cz����gcμ[� ��~�,Nz�s�Dv<����.luӖ�g�J�-`bh�w���G�t;�=BgY�\� U��.�gWz3�+���0�p���O���o��@�Li�r��`K��wl�p�G>�RWW�©=n�R��n�Щ��3	FT��ɉ��on�F�		 i���d�������^�Í���d��]�J�J�i�博��=C��#�S|���aH_I+`^�H�o�ᙏ��b ���F�>=¦��pl֗��x�õ\Â�LM�,~kިx~h�!�鯜oj�O+آ)�ۯwO�K�0Ni����w+{2p�U���k����3�]���ut1%ou��&hE�.�Q��	G��e�@����s�>�ڳ~�{s&���0������a��
 ����R�+�7�3�9ch��h��)�x}z��bVc�S�{���]ث���mu9�#�9�O�PQ|�v�<m���-��r��h��P�W��f~��b���[X�6�H����4�TӸ,S{mya�k����\z\^��^��۲����xx�$��(K�)zVș�g����g����:��h�:�{�����;�h�Q3�tg�3�(��a����W�!��:��py���݀**2��5�u�ˤTQy����Hx�G�-��v	�B�7J�@�L�11���To��{�=��JV|�j~�{O�별˭��N����{����u٩o�Q@�=�Q����	*���T�f����d骊S��N}���A���=��=�vD\�{p'b�`n���[�F��g�=堓	;�_l�lk
������O�B���w�g��0��*l�Ⱥr���|�]�׮��Y�!��h�������U.����N��+��|>y��	��E��*TM�P$�N��1O\��Gێi�wR�X���;�!O��JI���_M�_.������)xA		��sV���ԹvW+�>���]Q�G#!Z��Dߢ��2,�¦�_b�n1�����u�F��e�|�䍪��~����O�@�#y�&3:�����c#��/\õ�o"���3���Fb��)T8�k�a�ӣT����0w�&�o
�V��[��,�~��ؖ�P3j��~��/b�3P&�>pS�3ꎋU�@��<j�t����9r��Y�i1*<:R>S8r�Lc�V��1j*���p!PjF{���X��NFl*2|]�A�Dߟz7�y����:��Z�p��w�Nq�ⶻ֩L
�M�ó��|�� ��zF�Q�x�T �������:S�rɏ/�K3F��J�80ߨr���j�[�Rv!���Lm�C��d��V&=�tu%�~�91z���j��LcJ}�z~�&Q��'��7�p�:S��LP|^ܻ�B����9��{54�Hܖ��|��U0�"�*�[8������$cv����P���[�䐲�V��xeR�M��]�#oAu"/l��XmNkͪ�b��BI��PlJ�wgL
���O��JS��v����+���2<�}�T��S�j�:���k7����q)�P�1N!�&A>�#u���λ��t&师[���tu�u&w���y�^]�x1��j��'Co 
����J������J�vSN3ǀ��<벞�C{��E����2���9ˮ�|Ne� �����m�E�S���cY��{	��
�yT$T&���D�#�y0���r7�v�F{|�0d��[L�>�E�f��;��GEff�1��L��x�φ�š��K��VN�ɤ�W��8�p�įOd��bW"�&m)���Y0H�]�i{5�F��'?�&M�qG:��p[7Ҷ�£��
��P�O��Ե��G�2�_g����u�`���R#dy���ة��į�|����6}��vѥ)�GTK�����}�N�1��O.�1jE�3�f��}�И�E�9��xWg�0f +��2	��*�;vl(;2?r71yZ[��%�$Y���WkV_�ۥ7хn��mfpnc��;�a�r�rq��\yH�d�F^n-��y	�`�C���.�����.OS����Y�T��/�驚�ɊE������^rP A��'l�O:��Sklo%�zc� �r�v4+��n���R��ydw��[{��&D�M��]Nʦ+K0R[X�%�!G��=��3 8&-l�����#��ﴡ���t�c���:��]��~r[<�MG����j�
Ϸ�VF��z�F7tP���+ g`,�w>62����f��Z4E�
�J��n��F�f�6�=8#hTz��;�癨�ϵƗ��������*����E�V�/��	�L�y~5�	f��
=�ʉ|yeN`�B��+$H�Bsqf{(N�5���%��֜l�:�Ҳ�Z�.��_O�˼��g�yr��ײ�,�U)�bvdw0+M`�����o��Y>���/�>��aV�8d�`X�`؞�2�8j��wW�H9�p�O�<�{&cuR�$���*/߽r��ߝ*
�_����w�ӽwq�ݍhw��n��U�0,%nnI�
����4��|�=c����x,՟ae��[�̋�G�� �jF��F@���8�iF�qQuYqU���s��H���	���2.���\�6:��������0��^b[k�n΢9��o�
d˷�4����tZ�AS��� TV�/M��-Xɏ���l֏�Vx�I��B�ۺ����$�.��EZ�2Vã޿B��cC�L��{��� EՉ���au�K�p�`���S~`�֣N��t���Ȏ��ӧV��}QJ�&�S��l.1qP8oCP {«��i��A�X��S��z� yo�O1*�[g�=A��t����k�;��:$";���5��{��q��&���B
*g��T1��.y� z]�s�Q�y.j�?.� ��Rdw-��ߌk,iP�HYϝ��������D��T7
��"m��z~��˸����	��aɌ�+��}N
��2�sӝzȒ��.��	�kB���7�ݬ�v��s1Z�+�*�k�;6����W�Q�4��|J[�+8�.���*&&���T^�K��p�q� �3���!���P�K}Y��Q5�鎶re�ʊ���Df*1	�6.b�7(���j�8�ȴ�0�;��jn��l&M��^��a���r�Ϝ4M��w��1|�F%|��(�(K���-��YI�������G��w�W��Ah��Gk�1S��ct��|��vSŠ=ɶ%@,ƪ�fQ��!��jr]�X��L��ז*a��la\�g �1!���j��g�Z��l������R�[�³6�\�M��k����b���k/ل\�&S�o��:����?�Y[��N�\�gs�Z���u	-�]D]���r�f}%��5��X�f�(+�6��e�K-��)��G]�
�ܴ�$W9�N���(��n�ћۿY���熦�U��6mk{"�d8��uˏh��ҹ���o����ե�x�cٍ������'Ӗ"��<�I��q��f���=��N� u*w̔gF��v�w�2\V�wui�&��mdd�[y�}$[���]ԭ�"�&�(�>�ߖS˗i:;[QYl�7�n�.��P*�4s�z�wʞ:	��&�,�U	�1�{�u�
Й��۳��R�t�A���޻"�N����u�LN}/	�xc֫/*@�&��|!���x��s5
/%��U8�I��u��.��L�}�B+8��\3UZ��M������6ü&���VKqj[w�����.V,��f��vk�+�W�2:�4�o1;7+��F��}%��Bp[%9=�)�Bl�&�8Y���]=��M�V���ͳٽd���2vdt�ZG��N=u
�vj��zZ�W����]6�K��w�lfE�:֫�B�Ծ4�V�uJ,;�J�	�.w,-sxY�D�� U���9��q�zZq.�6I���Pf�����#�����۳�[�+��m/K�f�ݩ�+{j̎nN��ku��L���T��I?�U걵�+iS�:0��V�_X�Ѱ�Й#7g]�Qm���V���XV��U}6�E�5�I�R��k9D�.x�������4>��D�rS%[Y��5�Jv�z-<`.G������̥��W[���,-$ч;���x�6�-h��*cv�,��CAR7�f�;]��� y�����y� ]{�+j��B�+%�0d�}y��Xm�k��D��/Z�4���
ŕՋ��0[;�z������ai��n;�6ӛ$T���(7�=;�N�{jCٹy��^���&�u)��ˤ�6-���8^�\�S'���սۅW��@{��ӷﲬ��n�b[^�Hhp�x�
��`9|�Ԭ˽X�sn��w��l̛���H,���s��\������[��s���Y&��J�������7��#���vՀ�ϹA�Y�~�L@��o���W��SeQ����ML!|Mq;���Ш(�iX-#cMƉ��6:�H�Lr+�����9�D����jгY;(w{&ɯ�;��cu_�%�c��0���a-�u^Qry-�s�&Ei]�<T׹p!m��t�F��)$�0}�"�} z)X~��/k,;��b<��LQ���FkӞ�B��ɵ���jp��Wi@5(����NLXf�ؼ�aPv��2���y2�x`�ٟ#!�
���\`5j2[2�J Z��{L̚/�_��y��xU���LE).=R���k�r�c�e�Q�`�NvqDȪ�E|���c�2~J�h�˟*O/�*V��Q�!�g�`��2�=Iz�ו}���������Ǭð«������ʡ������{�Q|:���w���HfZFo��=S7F�QqZ8�����u՝`��<��y�p��C��n�����s�s(�Or*c�����Q$NNQU>���(1�	SU�#�m6������c�����������_d�Z���Q'���+˦���F�ځ^�a�A]�boU�B���&� r���)Y�n��_I,Vb�7�V[���z�=�}�๚��]�k{dq�W�g�+z�QE�/fr8�CI�h]l��8�)+���6WN�N[9m�!0�9|;���t�y|[Z��?G�l��s��ך�7��&$@J{�v_�w-c�뷉�V�d^�2|�N5%|�B��W�MYД;��jz纣+z�@~�#����N���(�7t8_�2��`�D�&���tV���9>�aKVI�Q<��ǉ�����my�y_�Y'�i��)����=VdC0�����>'�.2��Aհ_�� E{"D�2��A�e*Tf���9����t������F��:*�6��QQ�*���Sy��o�)-�zq�q,�S��	�^��wx�FK�1Pj� �-��N�J+Jf<*H�� /KΡO��X��6�kw�O��k�ɘ��(���8��?��)L�4�bo��r�l�ټ][S���0z�B�(��n��ѱu�.9���^z3mn�,1��Ա�5n��˥G�v?"��G��S7^�������+�1^6����� <�7�Û���2��[��������+��B蛟,�mD�lQ���ڦ�Kރ$(��zI�jyNȾ��]�GT@+�n܈{S�u���7*)up�2F��Sf{�C��s�ČwWV]��{ʠ�ť���T��l�So�s��Q,eg�A{�jt�{��xZ�[]jXj�7;���rtD�
r��h�BP��yfP���;]ԾH�B��3�b�÷b���8�4q��3NX�Ã���n����b�t�&�vR����н';�ױ������7u{	�S{�B��w��>�MU�Uk�V}�*�.EH�tH����F6��+f�30�����4��ݤH�hA�����6�U17{�]z�@1��N��魫w>q�/�h�g�j���V��8˂�
�ħёy��ËX���uT��"�U�>p<�Q��Le]A�md��di棨�9yXef-sQYjc��.8��ֽp
�y������o��<;�M�C}�ri��b�"�=D�5�@���b�}U(��z=��\87A�#/�Y�go=�Ә��y���N�~5��1[|y��N�8i�v��\���R�'�{4+^I�r���	ߏ-�C�����Y��+W&�&6������Ύ���l�1���/ZbB�]Z��kC���c�N���a̾��A{/�e^W��g
*4����x�:��dѬ����E��T��}�*m�3��eW՝��X�]�*�tl��.���T*Fd�� �G��
�O!�����D����uŸӖ�L5 K�S�k/@��2>��'�������y���7]��Z'�{.�sѭ�I{���B�7oKal�~�1:E��q�c�(�m��P1�'`04)�]�Z�0\��5[�]����d��7SD��]u��k��fa�T��e�޻�؜��0�ٓq3�{�/Y@K��A��4�̭}�)�p��0� ZX��Z�\8�f�rwYI)����r4L�g����~��a����u*�o����\,ũ�	��'�LT��gǭ�wyn�9�'��)�s~�=tD81c*�BK7�*�9O�a�f��,�0����S�|��*���p��J���#b�MC�˧*��}�a�1(�}�luŨ���R.]z�q^�0�s`�����p�����H���z�	˷����*.�a|��fF�Z:��^��J�)"Ѫ�E��wm������ĴL-�t� ��[u�bS̲�ʱY}7�֏ؘ�XZ���X�]h7�~�-��E��fh�;����5_���������CuG�����)Xi��q��c@�&x/�*�S�!�,^>��+n�$ת~����gX���p�{ٟ���t�x�,/��n��Kn{0�3�y��ǜ[�&f��]���<���	K^��!ੂ5l�}�j��~�����!E0��k��Ď���_��<����v���r�}�\z	��"�V�ܡ�d��mzP�bz�pzMd/���tW�tlON�!.��_E(�\0D丮���Ȕ�l�TJ�1C�=S$�!�ۿ	�9��	ܖ�6T�ɀ�'�J.��uLk:ݷ��F,@�}(�yS[���s�BK��c섺�=;��>O�����q�E�pn�����=xb������n� �[l%&���)���ȯO��M	���X�Q�:�e�u6p�|.WvY�������S�:v%/D�{e����OGE��¡.�5Tg;M�O�^�
q�����U.	�aq$
�����;!E*�uѺ�kGUbֲ��"��(��6J���Bg��Gj/��/U�K�1���i���c6�����U�2��ў���a�l�Ӛ)����	sî���4�|���3y�*� �m˅}w~ϕ�1�d�E��N��װfv\z���'N�"~�U�#���%+����KV/�����t6���ʧ�P�
y堆�Rt)��J��L36l�_&A�!1���D��u���7��x�����N�J0x���k�<�بQcZ����]�Q.�Od�#��k���X������ӵt������&t^:$A�.l�l/{sR&�=O�S��U��+9�ؒG����ʣC]z�@ɇ&�[�	����ƶb�����<�)@iA��Q��/(�G�f�fU�͛U*�]�N�@���i���:�M��ʤ���ӝ3v�F(jC�}]Խ�n��>�a˨fW�c�z��/�8H�R���kћb�M�����YC���}*���'/�Z�&������sЏy���X�}�qץ�����V7\�鷺J�2�G��+f��(���6��Zr�5��K�*�]�2::�a'Wq�c�W۰ۮW���o�{��HC۵.����g+Iܐjk(���z�_C��H]7Ō3;��WK��*[�6�K@
��{�w�m�t�:�2��{kE��ɫ/�7�OD��s�/�;G�c7��XY?�G?�n�����b��B��,/�_vn���=�\n0���t���﬘{�,=⒛����#9\�wzГo_��Y��kuQD{0���׋�Q�HT�1Og�����Lv�����G����ST˭�H�W��5��è`o�0��K���Y�7�MW�����; �W^���;�⭷����:*��Ҭ�`wW�ED�u(裏�~�#�I�f�{����7�ޅ�1v~�gU�mqEF������`��x����Qy��	)S;����˳�N�����.�>#%���=��'�a���M{����9M'w�uvaN<��o:$Ƕ6�m+F'P�*h������ekh���~��WZ�%��5�<���J���p&����#�M�[�N�.�>��;T4�]�6}B���Ǵ�,6WvO����
��F�>�����c�5a��D]�~Nc>
�q��'ћF�0�	�-��2���##�����N�6m���l�v7�����+
�'�:Bs�q��pLr���"N.�̔9�X-B}ᨕ[����Vr)�������Y�kQ��1��A��85�[���:�t��
vOc��j 2��!��ݺ�^�`O��<�i7c��{�ܢ�eb�}H���-�<2�Bi]��<���n�\%��gJ���E��wO�Ne���\�]�Q�2Q�7������ڑ�ӊ��@�k`�>�˃�Z��1j#p��s�ߝ,	�k�C52qt�3��	c��I�˽q�|Q�'�	tjtyj�^ۚj�2O�<2�O�,s��`��g��9-����W\���}��*:~�!��ՔtW�=�1<��p�;���>����9���� T���=!!�q������Pz����8��])vx߅N����}�h�����;w
�0��IbU�ZJp��S����2:Wzw1�<�H�Y#I�
�E\�k8��"�X���_�������p{B��:�#�j�:�ի��`�N{�΃�=v�E�D���"x��?UTh�H��x'<��c�Aұ
��5,��D&jΓ�~a\h��HC���U����E�pL"��fOO�1_��\�5��������`�I.d�%�kϢ]>���&7�mq^���*ǎ�{�X\�M~V}������v=�B՘��@�҄6��NC��=��&���`ӑv��&�&+��	��ȧp_�D�y,\k��e�K-c�)��?I���Y>�[�Q�~������7ڔ����X�ȫ&vG�7P9�sL\
ꃐnMzya�b�u����,
�<r2�Z�[`�J��Ԯ���t�����.�Eă��W]�*Z�D�U�	Ľ;��7Ҋ�U�r�ySt�w�2�p�ЮѴ>õ|HIի1ۡK%�ikWTh�2���t���:�^�ܫ�Y4q�s�@�ܻ� ���ƻ�����Trȭ� M7,vg��{suO��(Qo�=��Q�S�g-��a{4��x:#���I����<y#�����m�u�O��La��r�bn�1��K� ��dytC���o�_�S�ڇ�u+�{�
B��VI~���>�œ�7:�只zM�+�)\S�� �gF\>.�#/���f�CJ֜~)��{ҕ�qp�� Ek�B;��k}q$��=��sLM�3z��������P�1�_x�����U��ލ\�z.Ũ��/:�U�3bH�wS�=ϼ�[�2��އ+���I(�Mڊ�Zl�ʣA��חDҵ|/J75��r�>�>'$nϢE�,}�ݯ/|���)��ߴ����^�@|�j�펚��q˯{�F��O<3
��z��D�O0�ж�b��T�p�����yוә������
]5f�����1W���u��v����������t1_�P���w��5��(��%l�����0�eG���^����UT�VEG*�=�I:=�{G،�)�K�}ۋ�*�T5�5}�*����~��jwn�H�
T�M�M1=*��̥W�.��"m�[�K�15u��*�CT�p�`������!ާͺ��P�tH3UK����>�����h�����l����������u���Û	�x�{��nd�JU�rpN%���t�K8��\ʹ�����U�A�^�@�6��g0]{����u�(��U����v7��bs��|+<ct$	/�nb�)b_0v�������ɝ�����4_H�6�z��������R'���!28[�r�EĭO�=UJx��z���٣�,�S+L����M���"f�M��
��w�=�TǨ�w��{�a�+���x�9��1=�
��5J��T���9����&���p����4%(�NH�fN�+��|=vZ9����IdY$��l�*�h���65l�`���sP�5��]���b�(�����O� o��r�h���ھ��b}�nE��B�g!P�>Ԝ���A��!��hF�jdںKW�O&�}�o6��[��N������{�Ā/Ҙ}�f�+����H^Q#�:=�=َ[�r�eZ̚���B���=-�tܸ�x��"��1Ԅ�y[�]�ݻ���-�j��)�ܲr2���H�J̳�GoW>��������νr:����y⋃5հ�{��^>8��UC���H�ݑL��ڊ%3	ӉNgo؜��T�/�<|k¸���}w����dP�jz'N���N�$�q��d�µ�b-ȟd5@:�7g ǭL4Ӛ�+��-f��ޚ���<N�5Q|�q����7J׺o��-Q���e���WS/������T�+���>�\�]J���l��Wј�êP��%]�.-̔,`�R@��5}���)}Hj�`�RYW�Y/G�[@8%.�7P���2ׄy��$�X���3��nܙ����j��=�V�e4oI�N�	BY6�d)�����ι~Q����q��^��� j��]��zM���Cl�ŏF�����2�ړF��s���� ii{�΍
�?i��(5�Qv`��W���5ޜ1u�-�t�vz�J�}w���X_&�t���Q(�<�*��=�
~Pf�w�v�w������ޢ�(Y��N�߫�點֨��Z���Ќ�]n|�n�������rT^�~�"��K�Q�l�/���(���M��k�,z�9�Q��"g��:�s�a����"����(Y�h��1Xu��F]B>7��
�-��g_r�F��Yd���t7��,�Jb�����t�i?F:䝵��C�A�b�S�
^��d>Jc=��#�K�ǧՒJ�0�(A�-ێ}���������,m73l�
ܩ�}��Ek ��@0*�\7��L{%���X��Z��zQV�͏G.2Ɯ�����Z��EO$�-�	�m`����a�����Sn_�)
u<j^�ڃ:�q���y�6Lwm�׎@���XTK��)���o�P�6�⁧C'q��s�*�ۏj�'@c�������ؘ��ᕚ���5v��x�;�x����2XM1I�	���@J�9F�J�Y�2/��$5vw��37���t���'���sT2��z������\��}���Tv�K�N�57זy^�Σ�UU�7{+��v�[��>�v� �:h�wz) �i;�}鬬�w~�*�	8��a=�}�3{;�{1dDE��K�&�&�F���Lfm�J	qq�z��ƈ�A�%��z^\���4g*��^6�a��Vo/�<M�����V���/�M1d��_���8���ہ��M0!2���N{Y]҃��V�KF
DNAs K�K��ŉ�-��W��k~Ձ�#eզ/������Jt��ǉǦ�N!V�8��ҿ����B�Z��u_U:1���8�C��&��δſ��U���e]
a�4ȭɛ$"I5t������f+ ,���5Ԡ�l�@ ��V	m
s7��o\�N��w��Z����=��O r� ����o�λN���_�����<�0�`jC�$�$�a���j�\���%27Dկ�������M�U���Ԇ��JP��1*�n��E�F5��+�7�Ɲ�r0to�w�_O��K[xkg^�-�ZS+�����v����7vZ�{<��;�}��k���ӂ@��{]�r��0�f=qݙN�[�R]�kp����/�[���&�6%�n7	�N��L}v�^��SL=;��[��[�YD�e}��֭��qd��L����/���uǓl��D�L	�h�SVYEA�$-s�w}���ÝjI;��@<k\x�w��f��zy����5͗�TyW�}SH$H�1P��7�+ň��)0�aB���4I�ĭ�˻wSs���M�v�*y�����n��;�+t>������?}j�������8DDa��}H��[:�TsY����܌���ԭ��l��t�	/�Q���
���u�u�&9��ZKKa@t^%�n)��(���W�]ie��e��v��mAx�(��u�%���S��
�՜d��YR4r`���e=c ���N�.+�h����8�*�u
�K)�������ݠ�gJM]Y6p����;K�Y��;Q��m�����1�r���
�f�j�ݡ�;�oV�q�p�.�j9���{���-��$y1��Ŧ*@Vn	#o�dFz����s����p�2�1��z�[�:�]6K�}��s���&���%����&��ժnSK���_{ރ��:�u*p��(V �m�z6A�Zy����r������-��*�l�E�u��Ȋ'R+**�
Y��]�ɯ��{,�) E�&Ȉ��:�c�l]]s�C+q��@�\&�K��v3ـ�O��1��'oi��mYھý�l�Pv,wu.���;R�ݕ��7��iV�' ��9��ͪ9P���T�oY�wg)@r���vN��1�),Ffhk��A�9��a�3;�Q&K8�.����][c�}�\�Y��P+�����J����ݹf�K�`�~FZ'k;1:9k(u����Z��BkxM���"5x��r���e:����zv�"�M'���8��sbƨ����<�=K&ء����,����H33+7,=��G�7�՞�aE�&\�	��@ �M��Lt�̾a,Yy��+��­nڮ��q}0+�no=��ލѮ>y)����z�eɀ���p�V�t<�{7;
�K*�o®�N�tk���^�/�.N�VՋ�;�>Z�y����m�=���	����օ�����UH��_g�%xR�q�	��M���wa�cÖMz/��V�n���E�o�`�Fd��ax�ޕD�/�M��k��PUő�m�<�4�ULϼ��ע�r���f������4��^��#M�q6��ٛ8�s<;�T)�YD��=y���"�,	�$����FΪ������Ѷs�7�����ɉܛHa�M����5�T(��?5㕕)��M�y�P�Kwֆ0�]yޑ}6�8k���ҏM�9�#wB_r{sv�JP#RC�����.S��޾�KҸdI���\.���p�I�!�ia�Dv�>���u�E�(J�*��\��{�<�1..(8Rwk#J�]�*8���:�w��	�xTp�J"�R܎"��+o���ۛV��cU���©OϦ�����a���0^!�~N���W��Og*Eһ��mn
T��08�3t���L�廗7�ŗQ��*aՋ��o�k���K ��a��^(a�ZP�H7= c�ʋ}+��9�щ�w�=rl8���'�]>�d����]�r�wu�6�(0-g����Iq�*��. �]���[δQv��>��rf�=��_Nl��V�=���,�J���ժoק�-���w��u.��Ͷ,[9Xgn󔤄�C�иg7�(��U0����#�Ny7k��3>co��=�>5�zajpr=��]6t�İ��/�O�ϔ]yn��x�b�Cײ����ƉgU�Lza���W;�ou�8�*sa�&U�ECH\�9Y+fn7�=���R���>Sԥ�Iq88PZ�8��Z=�@׶��]Ѱ(�N�G��֑��ϲ8��y=w0&�,W' �����(L`J8�I�H�Н�05����T�u�'ܣ�b�O�(۩F���sG�R�d���Fư�>��[��#�]z������l1-�
��ڼ'�Q���v���"N��4*��*�f�*�,N����,o���yl�n�>�	gn�.�N�X��l�9�ht�.�>��}�=��t�ol�x�P�B�;�|@þ�����^��KN#�hG�6� f8�0'���eA�"NwQ�S�&\�gH�}�l�2��Z>��(s*,�(V��Y}��;ͭ��Bsz2�ؕ-תf�F�����]�2�Э91� (���t�oB��:���Mt]���r���K?P�u}�x;&w{*4����=բe�3�d��E�7a�J�UM��ɗ������4ozuj��x^�m�+M�0/����������tN�u�5;�ۃze\�U��b�Ԩ������E��TS�g ?"��A͞{$��u��Y��Z6���k�p��ɡ՛`�ڶ� �^�{Z�� ��>
6f4��,�%�:����D��M193�!�Q_��5�w����K����;pe�3����X�M(�jd���0�]ǻc.�l��+�n��R�Z�d���w�Ln�b��Aft�	vZ�X��6���E�T�'�/a��#��M
�d2�����y>���G�\�mL�]�ݾ2vv�߻g�1�_'�y�Tl�KrD����#�sYu';��4��[C[2!_�,y���Y2󔭞ޅL��B{�@B�V�}�N1_��콭I�Wg���m�Y��/�5�ǋ����]��1�x_O�qd�#�}��8�\o� ����tgE������i�b���ٶ�'�+t��T���톡h�x㌟���;�Z")\-���~`����qmM�+T#�v��/�d��/�3k�Fq�-z:�w�F�㌸��UM�Eq�2�e�z�@��1w�"ť��Mo���i.F�)�T?lcr4�0#S��k�8����Ž��Ýڃ��ZR��ڻ�����6��*Qkm�\���-��yJ'(���j��L�7B����`M���*݋ӝ��AEQ�3��tf�3mfWe�{z�R����57�mos�f�K7��p�/n⫰�,u��[�����s�3:�Iq���ͽ��gz���hŇQٮ6��l%��ic%ѹ��qn޽po+l��ya_i`L^�Ru�*�Fb10+1�r�N�O�.�y�"-G��')>�Ⱦ����<�ȝr�j�
�+�0|<�ޠ-N�������w
'C,n�+0"�����s�-Z�6j��~)�p��ڍ�z�<���_y-��PlrR�����!���!Y�o)��s�ɛ��uT��Gv܅�ҳ��>�)���i:50�}
F�R`{%f���߯���7~28m8pj�uKٱ���d�@������B�^�h���t�����S��z'�y8܊��[b�jv�=�� ��Vv�ғ^���\z����Y?q5x쮫�}޺��1s�]�Ip��>qu��

���^"�?S��t�����"l_|)@\fY]]�0ch�'E�&�Քv7g�쪋4��+|:���cˤ>���H|L8=�~���I�]ʂ����zk�*��́FL�(�e-��}���&��|<�L��r�9O���M��أ>�r�M��r�7����SDA���~ȅ���f�u�m�:PH�)u�~��ih���;���s�o�[��n�������aǵ�Do4��;��,{CL�]��^��V:y��wNӖԬ��c7�%���T��-
C~RM�F��Mm����k^'Y�]�H\qJ�K5�W��N|r%M�ZN�K�����c��]�gl�%V���� qA7���D;06����^sW
N��P���]������M�����6�F5������N�鐘�	/=�y.�������;Q��&�*zr;'�K�S��E�Wsy�8u�fH�nҎV��ݘe�8���o�o_]|'��B�g`��o�&k�'=����g�_Of����\�
�z�C��ݹ��W�S��Z��2f��F�Uuz�x�UkS���cq~����)L��OM�]uq;f�;S�^��xv���+%����Fy%�S��Hz�Q��c`&�4�{�K����D�S���W�3G�v�lnj/��bLhKj%�\���bI=�Fm^'�,�lܕX��Y���Y��kn%�'v����m���+tWDϲTfk{��FA�V���MH���� �-Q�ޞ�%���8|����쭓l�+���@>�L�����]b��eI�Y�a��3٨\��5��d M�ʢX^��ڃx�X�fX.�U���Zhq(둖/$���4@���]>��y�E�K���S�1U:
����t���ɬy۔̇��w)u�٦�*E���hot/b��٢�.�N���&,�儺�Yk�����j,� ��T�1�úe$���t�kU2�7;4�q �̵����>�'���q�
=]���t�[P�u��ԁ�:�y �wjxe+o
 �V/��uc&����ଅ���}I9�-@W���z��3qwJ��ܡc�<��`�R3;,�(R��������U�d�Ե��"S����k�ű?Gy�1y�g4��ۊ{�c�Dv��~]�(mg�r��]�	�Y�W�X��nI��zI{�T��y���qu�x �B_�	�?e<���v��m(��+�=�L��m{���|�'��>����o�w�,ij;�G}��u��zh�n�[�hs�8`;�n��L�C��5�Ӂ����Z�\q�*����T�������������0|��l}���Ϧ|t���(Iȳ�n-k�+�-���]�P�]ڑ�ȵ��ؔ��po6[C�A�޵���3蝻�,2f��p�[x|}��:\��4����^�ɯ%_��s�_���l�ى3D��b�Q��9�p#}G���C�0U�.p�<�ڮ4iw[�����q�jA[�Rہa���һE���m�>�;�e`�f���Ks΢�Ռ�iK|��b�۠T'�6�%&��ǧ��k�\]*}�
���Q�j���eCŤ�z%T��]�j.'�!�5=��jr�Ҋ�\�5��0H����d���0[u�����´�%��
VK���͵W�\�3q���'��,{ư�xA:�fk] ��`����qd]v���Y���ȴ������+
)d8yW�.�^X��6q�����0�x�1��`�*ςک�56}��3=��%B��{�U�{���T[�����VB���p�E�9��^|����;�bHq�:�C��!�0@n��W��1Vh^��	��Oݣ^qQU
od�Y��gT���G&��%(�\�e�k5��]Z�	˼? ]�'�|�޾!Oƻ���x����2�xV=���k�ܧO����0~�**�^��c#���ը�{��6}�7�W�qZ��Dr!�%�Z��@��%�/�s��
'�5Z�p�3���0̼�yj�]�2l�Q�h�lMF�Յ��iPV�~gT��b��U�~e9Ӳθ[C<�-��Yȱ@ncJ/�Џq�r� ���{�6��^��w����n���˘����;������Y����/� �kW���B�c��8����kȕ>B����������gy~��V�N��/�/�nǫ�/�e�o�sU�[TA�s����k���+���c���I>�F
�f+D���<滯��e�˩���:79r7E�W�^�ռ���b朑`�݁�aoc�s~�4�^?,XOeJ�ٻ�!(�m*�ju���y�;p+��7�NЉ�t����c6�g`$��M�a�0���-��&ۼ�,iQd�\�陧r\�
��0�L\L��w/JV�jn$��-�P�˕����m����G��c��͔s�cJ���h�߸Jl���:��[]Sp"O���ٸ�kH^%�|�+$��[c���ꨯ�f�N@˩�n�ԇA-�w���w�=��Y[vCy�k����M���U�oA��¼�G2��S;�הo�}�Z^
�V:7yǲNg�E��/&��aI�/��y��,[��UL���ߟ�s�L�^q��R|#�X�ƭ�Z�,��b,ZX����M�3Vƣ��o�1�*�ו͡=8��/\�8�L�VgK���'��(JQ�wK���m�[��}�ضBr谄;诚��x��f=A��_�w�y�r�I���]al����T([�u��˽q=5L$b�v�޳u�̫@x���!�8S5�#|s�6�PѐaH�q�wy1a��:���Y�����<�c*���s�bm�{L�1�A�w��Bn�WQ���B�5�4�E�&��{C'���;}t�V"�3c�a͆x�ŭ��[G��jTb���v���ԗhA����G�h�:�ۿW*�KaA���*�2��rW}3^����cL���v�n:d_�ڑ�����tw*��w����0��-=���/4��F��!�r�%_B�Y�]����}a�����|.�
�@� ��u
��ֆb�34%õ3R��Q�:�|8�aݕ�*����]e*�n�n���&B4ع4A����/'-�mw1����T���6�]څnrH�.����g��vr���ʗ_r�*^s�t�ծ~��F��t�l��y\��#��jD ��'b��q�o^߽�{w���<���Tx��o.�+��혪Ŝ�-C�	=t��>�.b�Ui��w��N�yۮH��fR��n�����R��3����y�ݦ�O�U�|�@�N�A�J��C�a�qV�T� en��Mz��2B�<����bn,G�D[��T����W�f����J�?b�,E�"���vO9�����e�u�hiʵ�j����0�f<!]C�և7�����(b�����q�mI�6qf�z�'˞FyTb����:�����2��;mO=#�E ZZ�=�}FJ7�bQ�ƺ�z��{<n�(�t0�X�X#]�S��1g�M�����4��Fm�מhp��i|{�[n��T0@�f��q:+/�W1��'Lr�.���xw��(+Y-G��fd!��FF���=X�v�'���~��h[kT2x'_�А����6!���N2i�������v�}��*�K=��cfG��u�}7�'=��+�c`�>��r%�a�,��<]��7X����ݺ��wvPF8�ǻ�XAQ6W�^2ҖeDK{�*�Ɯ��ڶ��V
�w�Rv��]M4:�Nh���^b咲�-�|`�wz�� �j�v�iX�@��X�^�],�Y���8H�����8���_��vC��dN9��\�+�Ep�����v�ex14?0��:A�Z*��w*v�ڽ������-k�ԈQ��b��3�{�n�^̜|�� ����� �縃�T{(��8*L��n�F��.�(7p��u��tL��e&�N�h��r�)��'�Oj�-�Uv�u��"h�s+7�1�U� C0n:����)@�D{١B˘=�-�>۰e6�WWx�xOg#)�.�~~�7�1�|'�E�#�){�x�~h$����
��x�>�6U��?�P�L�t;<~~]
��f�5h����l�W3�\&	�����[}zr�J.ɻzMw��v�|��/�ƻ����U�� @<k�x��2G/�1���8�怍ӴF>w!C�|��j���o�������%^��w��3gfZ���s\��!Vc��[������%C6՟b��3UğD� �Ma�bv	��iK��Pg-I��u�nӢ_-0h5sd\��M���|S��;�q��a�y���<1��3�=�O=E��p.�fiU�:��]�hT �o�:�.��O	�X��T�P�YUy-�\y#<�8�V�����M��k���^�:�1�����'�J��:�Y|@Zl��[!!-�ͅU��\r���+{w���@��06-�y	�7:�D�f����	��J�u+pgV"vv�p���ѦW
��tZ؏)��K��͜���&K�3�8Kbq}��\2�IY�|ԯ��8�9d� ���to��oW]+�p08 ���C$��2`?Qm���w���2I5��������Ww�ʹ��V��gkA���z&g�UY� M0�����x1bg��:�����5B/��
�{&X6�C��]gTk��;�*�T�1I.t��O%Z��S*^��d%�7�y�|g����W��IIz�<��pֻY�w��l��w�j���G�X[�n��3�s�:h�v,;�ʾԁ��諒 �nw|��jLrb��6��^@�f�bhx0�H*T f�;�=x��*�#ڷn�G���w�x+�)�h��}N��T(u�����Q�����ʶ��UiA���0Jp"M�e�U�Jm��h�	��e�V�S��6�9ʛ����J�N��1���{L�����od�XQ�5��,X�H���'�".P�{t�Zy4>����@�X_n����[������������Λ�o!��;�ڭ��f=V�>�V�W�)�7�g/��/1VI���92�+TgWwt��h��\$��m�}�z�a����u�I���O��m)1+TS�4�sT"���k^9����/R�˖����_���
m�*\�v`&��Z�Р;��t0D�=��B���v,7xj��qpv�Qh�ԕ�ܺߚ�Dn�����b��
��WKʗw4���/�vH0�}uOl��T�}O�D.^���7Hu�{|C�W�X��r('GՇ��Ư�%�e�i �.��lK�"�f���������!a���z=�����Z��~�^ت�4���睹� �[�Ѩ����zV r�M$]-�J�d��B:�0Xr���G�N�͉�rh�+r��!i��%�NDg1�ڰ�컡��.9�I��+Mc7�r��F�{�W!/�v��|�n':�V+i.A�hp��9��$ג�L��]�>�5�]	L(LC����ʲl�ɍ�A9�
�lL��s�r�����W��Y��1km�껎U�wW���G�G]�n�-<�Ưy�E�iSy��s�0s��s��℘mZ!�ѳQ���*V�Y�XBu��Ҡn�1��Ò[�VjbƥO`i�	YWh��ѐn��)�(Q�h���B̳î�s9���m��>���$'�:Y�
�0������'��N�F]������:��KZEbs�:q=����r:�9��1N�n���J�{��fccC/;�f��%��g�#�R�ZZVU�Z�+�HK"�&g=�*�$
c�~�|���ts��u�t3M�t4/����u��*;[A���W�!4�ـL����E����V4
��;����]�|��WuGOO�s�{��p�S�V��L]	��&p���GHY�x�C��왈�m>��x7�;Vw@���K�yg:���7+����x�(�s��*�P��돆eL���ri�V�]ֳRJ/�:YyՄ^�.=ж�Kբ�11o���k���}��`�I��V�`�E����i�bc9���8r��`�����K8� w������[�+u3HT@�/z�mr������7��*��Sf0�dC!�sv]���v�Q!=p���4�8U�vR��ܨ��:�G+w���r��Qb@�,Q� ���U�+1���V]I�0�7��w����9�5��ֽ�x��_VZ�0G��h�e8���x�=[���*Gz㑙=�yI�����(��5Lz{1�[Z|Lm�]t ��.���%���U/X��]�~ ͆x����]F>�^��NX��uߐ��_��y>ȳ��Xv/7���1~�=�G�+��]�;��Q�&c9�@�L�7w���������o�1Y�	�Y�f�>�2���2`�Y�BU�,CB�[>��W�zAP����?ښ���	0�ꗣ#а���t�obV�0��#3���<O�����Gr��<3g�c��<E�𘢪KH���D�{�|e��y_Hwt�>Krnf�Dr5�����GlcqQJX��Cϛ^�$�U��������6N߽��P~nh��ì�*~��{C�NJ3��b �q��}��G}q�}��>+'�t�kxz���Z��f9�ٷJ�����ߛ��PR�f�V.k��Ù�V��'U�R�6v�f�owN��v�+�3�.\�(\��W�V(I�|5����]�S�?[�9�\\�p��TN^��*L۵�����i�݋�_�3\�^[�I���N�����0�Z�s��I�W�T�:fk#��j�,����J3�������&N���VC����1Jo�6���2�0kLJK6�	�kK�vؿQ7u1��XέO�.��u�ڷn��񶎏z�ޒ_#�ϭܮ�.�(>WB|d�נ+Q�e���~�vsԱjJev#J��*ЊW$Opn�O�������M�u�3�w'G��;^ׂ�[��y�P��gi/ų@��c�Eg��.�yֲ��}u�>큓eh5�}Z��#[�W�]��~?�p�����T�nު�.]/{.v��瀍0':�L3��p��z_��������p<�w�c,֮�HX���.��wN���ػe;3P&@�~]��f�ɡ�V#"�\+����ǌ�W��]��a�����'�<����r��j��0b0͈,�[9=�)��.�[¾�@b���ku��{B~��X&)���^�t�Z��0�2{$��oђ��^+ I��l��מ	s��]�w/E9c���T�C��UK��t��
1�3�x9��vG�t�zj�;O_��{,SQ�`�{DR�v�t,��DܮF�g_rC��u��Nz�l��6j�>z)�4vjЖ�h�=���]68k{.`��E�v�s�,�uķ�T�&���Zn��Y΅[e�R�{����J�R� �Z.�Zz8�(r\�ؽ��y��Պ�$MBW[]��3�Q����'oަ<7ҬT����֋=�8�<���立����-(xVo%>O��w�"й5^�3U,�Z����qQ9ln���,vﯯ�s�٦)R�=8+�Z'�
���!�3���W_9�UP�=$h���;������S�r�������&��X=B
�ڱRa��S�cf���+Ē�+��ZU~���&�������<�QIN�8^�R�����N���t.U�*t�;܍;��#�{�
��x��/��~�8#w�79��.�Ǣץ-C�Sⴞܞ4�ǵ��\UT������Z�3Cp�<�=^����š	�n����A��p7���\��q11�n�����~'{k�ȣZ�z3R�G�g��s�޸3A�X���fݵb������\���\��h)��^W��*��\n�W�P#���d��d?(ݸ��MV���Z�_gz{"�!-,cY���5�.ۊ��c�$,��H��-���fg��brZ7;#�H�<���M�.a�m�*�Ը�>�2l�~��\f�`��)t��U�l)�]w��*�?e��YR�5����Y�� !��چ�mK��]�| �����1�\�Շ�_C�C�8Ŵ��R���Ok���M���0�.��"�����D$А���R2I��7V�e��%�ŷ�Q-��+2{o����s��y�����Z�)�S1ܮ��d�a4�v�a:�Kָ��X�V�/x�R�R��>�s1Y:m�b��67h�� �X� b�t��&(I>&3�޸������켹0:�/e��N
�q��"N�}��xVY��AW`Qjh�����B����o�-�93�5(�����v�m�����P�RU�J�)	����A�w觷�����4O���B�T[O��N�I�w��Ӟ^���!�߻O߰�Y���@�ƺ���*�u�;�����ś>�<ߕ�����6�if�6���;��W:��:@c1�6s�Õ��qr`�5T�^{��F�o槗����'?6��W6��R;<`F�.pm��{qt�uB!dxB�ytӘ>�'`��*`��k��FJK��j�x�Vo#�"��N���J��)��QZM�d$&�ik'%��ܷT_>�	`�ț9ę8ݳ�S`E҅��TyvwU��U�S�Z"Á�X�ђը�bO�nvZ�6�<2�:'Α�/���8�pY���F�Y�%Z��3�5d���27�Ϭ�#Y3��}Ύe3G���)��Rk5��������+���ⱺ[I���f���s��шf;K�0�����Tk�=�=�t�J��7x�q�
�O^Eʦ`
�:�6�Wuƾ���������K+&+�'�,L�tk�V�T�q�7��(1��5�3�*!��g��.���ƛˉ�>��Y7r�B��Fz�t��Jt��46�/N��U�a���{[�45��&Ks��G�g� �`�~��	9�O�=&d<'���;�C��i yZG�켖�,�xg2<������ɓ��vż��ۛL�υ9Z�{�m��𧻌ʨ�EU���feI�|(\Ѕ�c](��P���l��	�t��BW�5N� �Hb�G��m�(�dC�b����=�gr��n���ޏI�v:�8J�v&��yA M�����_�팸�t��qL��&+q��t]��⇇{PӰ|�6��|�H� =� [Qtߓ�㢤��G�]������L{�I��|���pf�W�b�����̮10a�(4� z����wQA�u"MB$�g�q����t�����t�÷$�8\n�}�+�ʚ�Ys\w�.�_8+�:����gc����G�l�'|�VL���:i׆�)���;t"f:	�cg�+��pܵ�h]p>i�39leio�	O�8����-sx&Þ�I�������	�Ru�s�ǝ&a�ʱ���3p���кAû��J#q3��&~�>[y\%��k9U��c���f�&m�,���ۀ�qt��K%�v2zM��=yk"�FU���o* RSvvd�걔��ZfQ|7n��|۹Y��S�|2ht��I,�Z�ڲ�3v��-7.rI=�;�9�����;�ߩ��&����j�p�{a]N�"�����t��e���L��h����h�iXՅכ�t�X`'����!��t�p�=�<��9&VJ1������q1n�&���s&�x.a�����3Ml^�6��?b��{&}�c<�iџ�[ߕy/ڛ�;��r~�ݵ���.����)��*�x�T'����{��(�~F�oM�������r:ބ9�׷��X*0z�~��`F���V�0!����q��_dRcרj�/��l�[��Փ���3��,�y�Qx_�$����-�Lr�\���G&Gc���o�]��L��0۝��h�T���G�gv�����2j';_�g[�-7^k�%7����ʙ��(�>�.y�]�U͊�D��#��x���=0"c�M�A��ӹ��^	�ṗ��cU��xȺgtڡ�=�m9|�N�	�k�]>��~-�g���3dL(B���S&Ϸ�݇DjoN]�]�uV�*DW�>��=Q޺FC�r�ދ˫�ݱ��Q�}~8�㼋;s�'.�G�qc�U���d�|53+h������L���"m$��Pm��m���4�aS�/+q�Ws�s&��z�[Y`��Ӡ�M�/��e^.�R�H�
"��v��؈�fQ��aj��r��ʩs�FWv_ff^4����8lGk����ײ�������)mm�!�2]��g���1��:p\�t������B&VRNiG<��jGO('9�p��L!�@�>n���o�k�\�����sJ{�%��)���@8WP�S�W�6.DV�HdT2s{��t��h��v��=��q(����٬�/�'P��7*T}��O>���H��d9�<u��B����ʙ�~��г/����z�g�M� �R�T*�ƽ��vl��=�+�d��'1���X`CQiWd_5c/+)��he�'M�NXXi�����۩�lB���xW�^�����;o<� f뇡6)�}Y��TI����N㱐����*�E��R�c��`��(���؊��c���c��Y[>���89n�$��>ߺ����b�OW:j��`�ы�ҥ���=[��T^��*��$K�����W���կ���]��-��bS�o$��Y�+X2���o�_L�1"rM�6a�'9,=5�j|�zM��#�vd����yY��������߽�Sy��gj��8j.K���=ټӇR��i-5��8u�Pʚu.��*��թ��m��]��wв�v����.��|��a�����ϫ�!G�����utH�!���Y8�����F��s�(H�H��39�E�d���d(����Y�U8
i�x�.��z'+�.�������䐉٫c9��k
�Y8iw��ɵ����Y��� ��Ӝ�gg��a�0Ou��V���5���%c�ܱwL@�_�o}�)}��]XW-��ߡ�%=�++�p��z�g)�A�A��J�Z؞�u�R{��j�POż����;��**:����=�3ڤ95����N	�����(b,�g5����ݐm�憐��S��������1쿚Z�k=cЫ<Ɂ+��{�����E"PT#���HKS��95��N>)
���G׻}v�_ٕȨ�1q�wP��q�չ:J����3�^���r�^���"z�ۀ�G�i��ﯽ�[��8�]���d-d��H�m�/2�V��x2��R�/6�.��m�K9e�s�����$G�A�����{�.��27o��WJ;���7�T�uZ� �7���x}�r�U�Ьa]{)LR�;6d5=�'��9h�H�l��%����B�78d�7���*�K^��6���nb����=$�p�
�!�9���T�ԯ`�6�P8���X=hG<j����&.6"�}o�9�-��q:QU5�~�ʄ7�c�1���C��B�nn媖\�:2�1��O.�`��r�@�v.�R,��ݤV�b1زYZ)-�H���{�9��cw�q��k��[�έwrý���g;2ԾeM�����ή�����j��d�	���p�e݆y���Y�fI˼�2`�袁��3�n�+WJ�yQ�8��DMR-�� �t�e*�E�X~!�-�2�C�Hy�c�:h	�;g�G^쾺��p����ڱ�~���8�ޡF+��`|�U�����r��d���</��7ے!/G5k����^������g����>��"�b�C�����F:����"�.C��$��5/4��X���wb�xI����v�ō�t{o�'��8_z������"���io^|���9�*�!Y�]�s]M���T�n� d��g/(N ;�,�<2�]�%z��՞�X�uF.�M	���
�;g<���Y�h�b�s��ݰ�_<�#�=>x@^�
lEt���z*�l�]��PAr���d����3��#��Q��8�3g���x�ɽ�_�R�7�K�E�R։��H\��;G�u�����~,nӮ��ŝ��/�T�v��L�Y�0��KP�m�ڋ�S|_WL>��'v�Ϗ_-n�>��p�B�\8f�LÉ�x���o�M)r\�Nm�%3s81|�hT4dʆŧk�_;^����fN��OF8�Nջ����j�j^S�,f)��`ؘ'���t��;)�ӊ�O:�V�f�ݠ�n�����D�]��5m7�Z�N����Q�8Z��6�x3)#|P:�yYa�_>ï�w������4K����`u`-^W��bS�W�7��/֟�����{�ᙾ�s���^1���eD�����rz�)�\�z�7o/],f�W�r�k�h��J���;�)[��wX�*�$[c��7�Q��yk����ޒ7J��޾n�^
���
b��$����l�aEz.8��״�jGV��^��|o*E�s�ص�
 )�s�i�⒜�:q�X� �/kEd�iLv�P4�'�.@&H��N(�.9�����Q���:�Oun�{uL�uP�S�K��Ӛ�Wڍю���qH��[5�fR����Ow��~���V����	�Ze9,�K�ɝ�rj8>:�\�{����U��x����س5�����ǭ���6� Tդ����f���V��A�c���o@[���
i���ػ�����mSl`Ĥ:2�y��bA w8�����r-�f�M�fs�c��s<Sh����ʝC�֐p�\D�nF��sS4�m,����X�X��a�*l�F�ȝ��;�#.�j���,y���6� �޻]�/��(p�:��ޱӦ�rp�I�ĝ,�2,�0�!�����JR��v��t�o9��+uu�*�t��˧����dW&�L�!i��b[鎃J���}W7OHŻћ������Es�cZ��*ާ�+8:�����t¹V��W�W�o1��w~��( z�Ǯ�f��0��V�ݜ�e�]Q��e�U���A����r���T핾V������ƵV��V��S9�u�i�f]M���
���󗗆<����M�}�B�g+��̊�r�������(J6���][��u��,\��yֺ�IYD9�̈́6�o�Ňh�m�ϰf]Q��\�g�������uوA��l`D���/��V;�6!�	�ި���C����l��ZVî��x�;69�70CA�"��v��3.��1 ����
���k2�ɦ��o��B�5��m�PeC���A;[�*��b��kUt��Lè�dĲ5q	5�7B���zC((�PHafȊŗ��,K��ea��>��mXF�yY	���i���`ich�Fs"L��}c̩B"�evv���!&X���� �+4�9�´�54��^�d�	�=մ�+%�͔g`n�\��p�r�b/tPY�3w�S�Z�p^�Ӷ�ovAN�{Z�M�l�k����z���n�VR��	c,[�����J(�\ m\�����ٺ�x'\ڗN��I�sQ����iN��{�_\;8�'9��RL��WQ]� �%̺Ve�C�;�Wh�k�{S���;���|�
�xΣ�'�7H� o��w����{��b�Pv��ruYT�-9J0�
g3�`�W�8��d5���1zs·��z��Z���|B��I혛���_*S6�{�m�_Wn�Ho�oC�X�b��Iotʵ�.��7|j�iT�t�	h�v�>��o
���X@�-�Y+;�y2ck.����C����Z,��r�����7{03�(��bo���q�t�+$��.��m!��ݦ�t(��0լ�.~ �K���q��Z]ݦ�V�Ƌ�/t��ެ1�m��2f�Q�G	*��@��e�gmڶ�7{�S'>����t������L�׭^�\H��\��h��a}k��7�D�a׎�O	l��ק���ݘ�D���>Y]yI��˱%�A� 
j�IF�G��n��| ��X{kz.��9���v�}z%�$�_t�ެ�.o.����Ei� s�uf:a�����ww��+zV��0��Ӵj�뛮^��a
9�X��R癲�k!s;W[Qr@]����úX�s9@���.n���
�z�k.�kf��Yy���Ww]vdF�b��<(��`�Lrӵ^���ѧƚ1fXv/�.'�Jc�)fk1F��/hj��h����Lˤ�9{����0�h=�e�)e�K�G(ūgmoW;�Vh�)�إ��5f��Yö�8F�w.���o��p��y���w'�'Ƚ�q#$���p�����רÊ���cen쇨�;P��R��Jp]�m���D�;p@R�vC+��<�2�w�)�b�V��]_>��pp"%+���Ra
�șXQ�	���}�}M��{&����8�[<��wA+S 8���Ӟ���<AlDp���]�f���Od4���m�t=3�L��׳�ڊ�P�Ķ���S G%=�g�=V����k4�_<�k�M_r�1^rq6g���ٲ�΃�^ks����Mgcp��l������W�ޗ��U�|����{^?_����!�bk�ײK�������}HV����	6avs�k;R�hQ9�Ms��h�-t�42�
������i���K�tٴ��Wzܱ���/��0aȡ��j6{�]�:�ki�40� �H{�QN�M���ݮ���୫� #ԏ�c�ѫU�gӵk�;dO�H�}�ڀ��w���$+��ix���L8�9�+5V٘z4�`�*:;&<,G=�m�
�)�+�y�|�
����b�y�':&K�V+aڇ�T��9�Z���q
&��l�dfV��OO\���ѯ��������rW��á��>�cxGp�y~���^Yf�cP�z��8N��4Q�u��:R���N�&ŋ�xe_!�X��L��Ȱp�]I�X�j�{�	:P;�#�z��C����X�>8_�����\B�
j3Yf�G����§͚ؔ�8پQ"z�Oe�
4b����̓�_��1ǅT������zhe��k��ssu��{	X]ɐ�����=�&�����f^�Vv�����X��`�z�n�8�p�&�ǑI�X��N�_<q\��1�I�����H{�P�o¯XE+���4���z��~ۯ��s*̛���$�Z4t�{2l�����>u=�ËZclLp����s"/�_�f�?nj�nd�)�x�*k��ߚ>>=O5L��{U���Lg'��,�p�G�B\#P�|k����u_Lp��0�;�4��'"|#��O��..�U����+6�=��\M%[ӯ�����ϑ��2y}1�+&䂭�X�gWM�ѭ�����s-bȶ�=�@n�~���`Gt9��+;d��M1B:�R�C�=�뾶��j/���+#�rq���`�Ȭ�woB��Ӣ�m��:?4Ӟt�����<9Ut��MQ�m���mx�6e��d��t#ѩz��R1���^WE��D_���t������=W� ��2m�V]g�y���q��`�$!9��=+��uJc�4!��s;�!1��/�p����j~zg!�E-U���
2J�-�#���	�
�g��_�`����b}��:�P E�頛���a��,��Z�����V�ԉ嚑ˤ��hǩE�%`���f?R�D�@��
�-�uu1�z78��y����͋���s�я���Du:�8z�ЫXcU:p��ww]�W��n�$:�e��=C]h��*p9�i�*om��e0E���x+�2Lа�6����P�Ɣ����N9�b���#tE�Z�cjE���wy%%��ƆB��{��k|�ň��W��ƪzk�:��f����iY1B�L��r�{�����u�Y��W�J�A/����Ջ h�s覽*��?�f��q��Xe>]�0��5������tuXV;�|�[隭��]��;ٓ~�Q�},7�g�r�F��33+��ϫ�Z�M<�.�����b�][�ہ�ۤsn�Գ�wQ�!Q; ��;�9G�3p�������Kd�hW�+��V�����x
oN�G/ߴ��O34yw��}N��7�WZ���D��}-x�q��0_���b�Vg��ׂ��R�eb�pxp���cݿ�R��M���p�bg�p]h�Md���m\O
��Cv�}��/Uqt�b~Mh�r�����{*�3��]�T�����D����n�|cp���ʣ�#l�ZU���y��F�*I�ۇ[��M�C����h�ϙ*dg��ybӊ�U�o��hޕO�6�8Iz<rv]�$\)[�����W���'��+����3�eHQq��v�����kHL)�j����O��*�.���}moO}z�H���lS9��m�*]I��WG2��KY�X�uk`�����4�q�Dw����)���5��L�XH�mV���}�:�^�l�I^s
���u��+-�����F �7}X����M�5��Bgb��P%U"�(��j �S�)V��^(]~j}
�v���z;�b�O��}lz�w����I�f�Z�1��U>����T�@���Ҽ���o�9�JΆR�<�)N�Q�[э��^Y�p�|0鈞V�eOu���F�B�U{r���ItMԐ��f�����Ge�?�yJ^]w� @�k����ǲ�M4�}�r:Bb��BJK\͕|Z�&n�����HF��Z�vr��}�#��ywV+9��������&c�/��K`gϏ���8��j�{���T]�R!m��,K�p��L�|���S=�70���=�e�s���
�\�q��l��d-	gg�c�-}� ����ǚ��Kr��\�q���<)�L�61Dw>�P�������o���,��UuG/7���0��c�eEl�ȣ�m��@��v���S��#ׯ��q���[�e��-��w4}%0�_+U��}��>3U��E����8K�$��Y��U���$2F�t�f���ih2cH��/`V�N>Q���:�*/Oۻ��{,˸��/x庻�,�ch|v��ީ� Q�+x��p�0���)2��eM��'JK�~�e���jY�\�8mS�n�^V@�s�fŽN#;���PaY��mF(P�y�A����~`�%ݔ�
�e�n����Y:\�&�\C�RM�r����i�_�4u�4m
������`\�7��u���D���Q���ws�[��Y��}��=�K�#j�!,���zFl'�9�8�vm���v�%�ң6�&���q�Ue)�͗�mN13tcO��t?A���֑����~Y���f���g�G����@�3ND�w�DN�cPK�ٛ3��^�����r��[�CqV3,��-K����e��qr���~�2���ާ��[W+��[[���N:Ak����2 \�]xҨmҖ*�]�oʅ��(���W@[��jH�i����d��h��������s��x�'�'t{!ejN�ڋ�S�z.�ع5���.��(g�a`ߏ>���Fl.EY��2Vd���J�f)T�qi��?Q���sgT{0$E��fs�u��{3��Tu洚�t�cSt�!�F��o9m���J4@Jb_!C������(Í�~��0�5gwu�fD����5���yVw�x-M��Zc ��Щ�۰�×�{=����K����<.���� r�{r"��(A�Y��/�f��q���+�����*&ʢ\a=��E��kpe��!V��z�w��z:�cGU�����#�2E��q�hbӽ�r�6������(MtЫ���|і��`��Xb�Zgf
r�0�b_4�`&�����*���"z�w�5)�X���Oze]_.F(*�L��\��e�v�j��A���FT������w����.�!������z�Ě��Nr���t�ƥr��r�:�^y`�Ʈ��{�� �I��#~�Z�<:G�1�j#��$��)�ߙ��93,FM���I�ѝ�Q73O5��w�s3+��H̜�Yq�]�����T ��{s�|�a!B����d&d�\�[�pa��t�N�k"����Y�(C���&Ş�X��JP��C�to��+O~<_�������$��u"��s
G�z�Ʉ��J:|�̸�N���M�(I���fGP"�=�2v7�p��9e��.̛=��NU(	o/�C뎓��s|o�_������^m3�Z��4���k�V��y����+�Z}�|����˻k4v�	qX���=�o	�\3i|��B#��nid�:�_^�(�W>SS(,�źgT{ �0M�%��<�0�0������}�Ww����<�[���Ǻ��t�<�!<�;��#C�k�vZ3�՗Ԩ�|<�t&
�W�sQ�`���%�yp'#���:y��H
7�4x��T��k�����e�1K�|�̓2��a;IWZ�����;z��:	ou�w��p���1��mLIVj$-�s�o7r��o��{o��١8%�M�چ�T�X��!Y��N$��Tn�� �r�)���&�j�՛���F,�8�	v+%����2�����[�×�`Q��'.��]ҥ�~���X4k�8<���J6�-�����kY��ԁ�����<��kC��ͫ��32]~��X��"n<�9�l%	�a����3�Q��m�=��]�J�wS�ꦈ���ȫY@����/"��a�"Ew�B�2�P���3ݨS�Y�5�K�zX���7��c�Yѳ�q��K�x�a���nD�D���{��q���{�z��E���W�<�;t2�<s���:��Y�tW�)�>��Xk�k8�d�F{8�P�`��TH���r��ԭQyj�iSz�EtV�j�Q9�'kqlpx!f5�U�L8&-E�t��\jV_D�����{u.�z�V����euLY��tϊWj222V�����,��
+�S׭TUIY�O�ł��\b���x�@l�[.?z��ϡTԌ+��Bp����]ޮ�:�@��P8d�[�ϥ����2�v;�������e�H!��΄����gŬ��m̱7�pSd�Z'|�� ���ɰ��ܞwO�*��o~��6���]<-�W�.S�����;j	Ci�β���4�OvR�d�U����3i����$�7B,�O �^��*v�-�i�^����}��	�U��Tz���9J=WI�xn��9Ұn��T�6�I����ths\�R��uu=��/²h���2$�n$+�	v��ќ���<-���,��
dz��ו��C{:as,i��N����_]���(�Vǫ��� Yo��c�HkW�|�_�*;ԭ�*�G �AFOD������('
��^� D���Μ.��q�x_]as�|\��=e��}J�����~���B˙�����m�u��>��U</�k�Y�"u@�D5�if��mwK�%(3��^�5h9�N�>�MKj�RُU㮆`q�39NML�cDv���u*�ƘY�`oE�ZቔI�"UĤ��Ɵ-^��~��ޙ�R�t�\J^�^G���8t�[�/��Aم�B�����%��� 39�.`f��b�z2ԡ ���p��y�ϞԔ�U��B���ŋ��B���_`�u;}zDh^VO~��YY����e�Ӯ�x��N��bt�{xj+��Q�,�Z� ͸\�Jf/���"gʦ�{��)U���&�����7<X����I��{^�PF�(����4��S ���r����%���v�]�����˙���y8�<��g�����jt�E]�NYZ^AE�����m%��]ֺ��-:H�G�I��{	sfj]�����3���c+b��_Mi�.'�ַ��H��W8�>�wGxa�lb�ƃ��ܧ��5���J���Y}݃�bQ��ğ�B�`>K�o� �-y�쩵9��g���q�	�A�L�\]��n��pk(�b�@�;�Q�����B5r�'��=M��{�i��~Qy1g�4=���Of�3B��1Na��x���=�S�Q���&Wܖ�X�L��<�Ȫ����yK����u�ȏ�����v��D�".�%��=F�|T��/}�m�����>�S��X�X����^�4ev�!}͑�7]z�f1ٛ��]7��z�*tY�w���w"~�������9���B��n�����6�b�\��d���S#�*��vJ�51��|3�w�3%Ee�.���x�c�,;Nu�p\`c�oG�ڌ��D�~6��\ �&sao�2H��9�ב[2�Lޅ�X���/r.���Vg��Ȩ�7{��^[���!�<#�c�����&DL�i�9��݄�gT9���Ϲ�'��W����j������Cq�HW���<�J�����v�~��Q�8.��9��{�3��� �)����Y��COu���<+sy4�%l�[�V[����g0)e�#��u;��%�xj�elz�+U�!�uBs+1e0(�;�n��Y۵L��2�i�&[A����LM9��f�c��E�����q}���賴�B�;�H��|�Ī`vX�]M�K:��a�6���x�PT7ϱ/I���K��련�V���Fwr�z(�a��{,����e���R�.�7a���Cq�;�#[2�b`]��ݵ��C
�.r��}_��9��U�Р�bZ>�}HM� ���4,.��k��������Py`��pg���U*��ՐEG���$m��Z����И�#�\���d�..:��"2��HF��+����H?(gLdb���=� ��
OM	�K�G��R��-�Q|ԓTw���5��s�uu�G�G��h�;�칵-����X�gA�x+Z���W�1t'ү�c��FG�+׏^`�WCg�.�v�n��/�mg�0��+������^1q>�y^�=lL��/���=iy��d]��:e_z�O�x��O6������d�G�3�xc%]9�T?"�l+�t��}	ג��Gm�«���e�3��R޺{w)���q-%~{����P���`+	�r�l��'1`�g�Q��\j�p�bh�V�t��P3���Y��f�Mx��_�ݩ��gW'_�|fF(���!���YW�l@u]���p�H����¹g�m'�0O��tӹ#��V&F���O���{%��������+V���T

r);��䜽pi�l�2bk���#wpM��ݏf���{m��&���V��ϓ�%ob �w���Ǜ3�J�}g+L�#Uuv_�WKe�t����']䷜�݊:oR�Net
vsS���;9�|N�6�Usj�VfL3`��R��U8��[�THj,��f�b ��RD*0�8 �Y��P���h�/�V�R/j����G0Aq��F����*���J�a������Vo"]\Q�- ����%:w��Z�%����]Kb�ju0��E��W��@����hu�w�J�vl�d*ל[���P>�e�G����W:�.��N�1�vV��Tb���bn�uhǔLs�K�0-�Ku(1�S��,bT��I�56&(IyW��d��Q�|A��s��Y�v�VҬQ�x�uٺ��P�X܆�[1���r�i㙝�j((ʽ�ұ2s��!Zvv�z*��`9 �̻#kj_E9)�Ql햢�l�2��F�R�E������@2�-�]����^n�ທ+g'F},zE�5�*P�׹�z�"Ƚt�,�:�j��t�J���l��H�ԃ٦�+N䜞�Wf�{��v�s�br�y����U�2����E�Y�.���LK���^f�+��;B����sE�#z�0�Ss��9�j��V���;��SyV�����!����O�M)���SX��t�Ӗ9�s%!�YiM!�z	��seӭ]go��iWPQ^쏫rt�w��\ܡxy�Im�л^%h>:�Z�;?�I���(�r��TM�6�J�UFʺ�w'-�K�7�.�E�V�J��o������Vp�L1n���T�c�IX��D��� mK����egG�����윉w(K�0`���!9&=+�C�t:�$�u��Ŧ���瓹i��b���i3l�-ܱ]����[7��f�;Uo98<޸�������)�f�����`��X�E�knc�}�r
}�*c���c����˥���t�h�x���۠ޚP�kHi�f3��렧g1��H��'~\N�RI�Tn6uL<�X��Gj
Y���Y��m�\�X+;i	��H	��K���\לVቼ���H�ꗺ�@z��
j�^Jy��&D/�����xǘ��g�u��9�d�3����.�-f��v�uI��T%Ү�W}⫶�є����՜�#���|����C#�;Gg�ifp��aΎ�h7�&�
	��k���ֶ��b�	�-�4W}�'����	����K��m������$4u�:!|��bCWA�(�R�z��k��]�M?Y�u� ¹S�����`������Oe:5�λ�tK{.NcN���F<[���$��m�L��ͼ�ӈ�"���̤0�b��I+�r�ҷu;iX�-��Uݖ7+u��M�;:쓋S��1��F�*������ĥ��c�9o�~@�Md��$D��o
�Q@t��9G��Kl�v��)圜Q-[X�Y������u:;��ɱ��AQ|����r�zduĴ�c���������j���'O�/E��|3Gx����v��V`��1w��� ��8(��\�/p9�γ���H);뎣�{0���m������u��WE���b�/wR>��Q���2��}t�����_��j�Nt9�Q5fE���ֵy�f�c+�W�G���,`��Ɇ��ﴤ�U�2��e�	Jn�n�N����d�DǙ��}\b�����"�`K�lf�z��ij� ŹWd�_LZ!�]N����z@�T��/�ލ�>EMd0m/U�����L�c �Q���u0a��|,�bo�*V6o�Ӿ�n�u���[��r�Ke��ׯ�cu2UB��~�I����;�.��X�YW�AQgyl�Ň�sY�����p����ٻ����zX��{�w�b�<[=Z`i����\��]#{)\\��j�H^�պ@��*�d1ʧ��j�;ko�w%��q7W��*P���AEe$y�
ԍ������2��-�������ܖ�hJμf���`��	i!�����|��b�&����PH���rCb !�-AA_m�]{O喥�9MvL\�
�{��.�9	���I҃}���\�I8����F��5y��$`����e��ŉ�̥T�X��1|[Lt]�p����Z )D���1�\D�o��sr�w��գ������L(��ٵ�6�D�W�W�+��"VZI�Ԏ��bcf��X�@[t�dl��񍍨]��)c��6fa�!k�m]�i�*��X&�]
�}v�V��"���(���������I���7֧aƎ�����p��1�
|&DLPA�~�rf����n �{wl�nԪŜ��G[ះ�E�������/U�$X8	AVm��ʔ=l��"�[xo�t�_�+���{<���'l
0�}�qS\3�Ay���	 ����"�&������3Q�"���>%r�5��W.�s0dQ�$$��kk��B�ʫ�m��Ʒ;�Q�;�o=�OQ�hdUZ��z_4�8^I�{>1険r�X�\�q�z��sJ��v��
̆52[:�l�8DAV&�Z�
�6ˁ�u��0����,��
,�-�����;��LR��㽺0�>����}���J�	fdK�]��t��m"K�\�ǯ��ss9����o`'�|�Y�(�&W�/l�:��*ۘ��W�Wv�%g�*~/�{t��g��(���|�6���wx��]M��u��Bp��s��X��h�'7E�xg��i��7�U��{�x����&�
�v�G���׵˞L"K��{"_T���X5'�A������q����S�;x߳6=�o�ϑ�+7ߟ�ӛ�1jµd�˧[}o��Բ�-
�Va>ns3�g������{e�8[K�wa<�P��]19�@uRީ�!m��q�[]^��	�z/pHmb�q��;H��rDlWEk�4gF5֧;�_vq��1�M,�m�ko�
�Mi���Y�����9���>ؖk�Nb����r��bo�b
�i����/EQ�=�W�z'���oC���8�?a��F�Ll^l��ط%٥��-��Gb�
��T5���M������|��#y�#]���m���L�u�7�����R�,Km��7�n�R͖��qu.U�_k#+)���BoU�7slq��c���I����L�m��C���z �)Y�;��ˮS�*u��vZ{�EW�P"x�ѽ�e_+�Ya�-��"�d�.�e>�������x�â�S�&w#��g
�2�Y6��}��\��������J�#��J3c�������W��5��oQ�&u�]��Au�ݕ��j�J.fp\�����2|1�~���fӼwp`0�ͤ1��]���Vb�sV�����}�ٽx�-�"�����q��3Po/�
&�Bz��k�����[?'$Io�=��OK�W(���ZAVz�.���uh.�ڟS�!6�u\�˥y��K��v�V�q���6�,�f!�z��ߪ=����j���m����Q��.�2Vm���l6��+�_.�H������.���#6r}��'�tg��f�4��Ž�CE}A���sd��z�1<�1v;���L��6��Sˮ���ڨ:i�34��ۜ�pu3�J�w��8� ��k:2�B{�� ��{����p+r�v�9m�9�%_LL�@�ݸnԞe�BcX�Gԅ��{B�U�
X������!ʠ[�K8
���Z���g�cMޭ�{����2�,�o^β��@��}׵�B����e��Lb��-��ݒ��7s)�퇵H]ؗ�k�[�6�wm;�݇�m�/U��R��Ӊ'uf>Uy�����^(�ٌW���G��}������d���U���3����O؁�]�f?!��Pm������
���q[���2�	tp㮎���C�;�H��{15B,Q��ʹb]���x�T!�5�B�x���f,4�Ƿ��uիY*+��{H�(��X�zFm���o)|G�ea��!�Oy,f4C�B=��O]��h��8̅�c֕���M�RJ�JS��<ԕ������E<U�|��
�l�~o֒ԗ^��[��w�w�w�=�0o��v\ʋW��"���[ ����?߯7�1��q��
:j���ʷ�
�㞱����tŔ=O��|şv=�����R4��� ���Y8>建j�*35�z�d�N��!EģG��N�����YCoú��?EK�b�̬�U0�� 7)Z�����޵�sn�]���皿{$3��ɧ����_V���@���9󣰞X.���q�����yF���}��q�-|6+HN�zM娬�m@�R�Ż9ȶR�..�mۗl�8�+R�W���ۆ��6]�a9�D����/a�{O�M���k����g;U3�R�n��WZ%+m�N���s_yt��3fF�Ǌ@1p��8DH[�7&�if]��A��}N�6S�M���8UBb(O�>&{��ys�j�{�b�⽝2�]���[͇�1/\�1�'���L�zU��'bX���C�A�el��v�<O���`G�'�#�����0z�V�}�#�ٙ�6�+��(�7~�=.i{���!Nc���rb�z�!]ەz42�����t�ɷ��n���{���NL&�1/D�ʬ��u�*)T˯�Bd^v�M<��_Y�Q��_�ج��s�,�Mɉ�:�P��(�Ä{=R��_�����ǠY�j\>�6�Yv�Q���5��)v�������J2�x���c������8����z^�N� �"�:[fͫ3���׀�Nη��4z����q�g�s7��>[r��`ƨ���v��^�%���vw���E<r�&o4��C�q�]�d�Q1u��'w�y��(���N�s�7���P�ߡT����&�����MŪ)a�j�3wt:u|������Zsc�V���7�����@H�Zgz ㅎ��(jg.v�J�<� 5���I狔���5hxG�"�
c���W��*RO=�CKk���-6�h��X�ڝz�w�|�b��YX5;0f;�M�<�,ݮ��l�!e�it[F}��jq��ת����Z�q��ڤ��%�^EP��V�z+�y^��׽]�}P��1�L�U��*q|o�j���ɫMl�?�uǽ�Y8~ �B0^ܨq�+T�r�c���]��q�����ț8Ӭ9zey�눕:����y�8N�Q�)��
ݞ�!�<��\9�9({,��㒄���9I�*�ᩱ�G�ت��J�05�s�&�{���lK[^IL�f�l�EByў�����_b�71�����:;I�ח ċU��X��l�M��~�w�-�%�74\�zgՙ��2ƌ�C��i��A��4���b��u���4T����y������������;0?4���O-͔��t�GQ�&v�'���]��O�&2F�N�o�5g�6a�k�j��-�D�y�x�-��Z����c�Q۱;:��{j�z��\�hk~�Sc@��n\j��S4�ܼQn���,ůC�D��@�����J�(��בu-
�ճ~Y��K�I%�N�xc��ﶶ���Fq�Ļ������ j��*ޝ���ed�5R��U�m�d\�����#�Iu����2�45h7�5s����UyM�H΅�lD�|Utz{��T�⴯����Q�A~��n5@Ł�X��m�>��T�=����?r��gh���c���
Q���/8�"�N���=y6�\�������rʵ�td�gҴ�wdV�z��f�O��<�_+����ݼ�L�I3�ݧ��y�tO�~����:��߁�X���t�f�L�`NM�V��/��^��<���Ⱦ�h�l�=�3ċ���)U��Qy�,{�Ԭς�����pe�[9~��a��Y̶��l�ۖi��$��Zzg�[r� �;��_R��:<�>��+��U�̼���A^�iklC�j6ܪ�kp��:��.\��y1n��k�����G���Ǉ{2�e�=n��3V���ߒ�հT��F<4,�S=yhT(z�
�,"I����O�]=�۷� ���G��~���?������T�E�~���
����u[,q�����r�$g]�U��U���5�+o[��M�7/���uK��Ǵ�N�� �
lE��<ū�pc{��Cuil��Z�ێ�[j�0�"*,�CPE^���z���]���fe:d��eb',�d���t�}��'�bn����`M������f����3:Z:�n���-��/�I����D���׷�3^�f�1��H�&w�Q#���� ��0��_]n������(>�[W>�B����Os�G�\��Y[�*7��C��� x]ke�ͮ���ݞ�:RDj�uݮK72K��g�Dg��[�y[J��W5��S7�H٭,t�(���BG`xi-q�2~�n_�܈������AF�f����*���LP�Jie�fī� �8�'��uFE�Kj�$F�9��\�����%y�/������\l/�O���{��y ���R�Vuo�H|�����v�{����=�1M��OJT���(���}=6��@���:��m5T*iSX�Jx�u'eaA�
LC���v��\[H�P�4}ceiR���.���h�£w���$k�7���?v�>�E�(>�'����r��qo�X@/bY��v媐'[�hIk/1��n�0G�|�g�:c���vFir\��+�<��P;7.���`���W�Rqr/t19m��n���=��mJ�X�C&���Z�휲]ZbK��>%����ۇ]����y�\ڶ���r���<�F�9јZ�N�2=����X76�������s2�Gg��w��.B,pDMrR\*S���� ��x0�z�X��bC�u�`�K���t��/ �!�2�t�ey��x޶5�ZI�G/����GL�����j��7���G�g���zN7L�,V��x`�W�����q]���ܮ�Wf'LOyv���K�M�i���M���*��c�ͨ���qL�ї�!�r���O���G�/���tבU��x������H�	��"�[�DX��%��hY��J7�]n�ؚ���P/����Y�&-	���؁��2E���f�NnȠ���vWr��w7�Ų�A��LB�~�&���BW��B^��b��)t18��F�קg�ʦc	�y�n�(�d^�{z��b�G��
�����=yt��g��Z�{H�u�U~[�]�N�c�%[Ƀ�ݬ-魵�M��"���Y�@H�gacA;�8��-��2��N�A��m6���*e���V�@r�+��C~A���@v��X�y{t��ڋcZr��wL��*sA��d1�v�s���,�r #O�RWz�j��SE?}���ښ��^��+�����]Y���ȝ�ӼB���ei}u�E�V1��$��r��n�.A�mR��5�3C��kGv�ؔ�Ӎ�{;���2��\ŭ�R��I�`Mʻ	�+K�&�q��m����^pcGh/n���59/�r���R���}H�	���,ܥ��ep�z��X�&G��p���!"��^7\	�2�
�|v&�}� �Z�%
����r3le]��w9ݏ7U�0��
nE��R#��Y��^�Vk	|42lhy����k�y�>P�B�s���l�d�W��ӞG�GWǞ*�F�{�2b��v��؊�݀��&BX�L5�E;B�ΐƽg +Y�4�wi�����ٓ���n;�Q���]θ���V*�/�j�ܾ'E:�t(]�!]��rn�c���wv3���Q�;o�D�K)b�Ҕ�w�>��Y�qn��U��a��Y�#�&�����tv:��7>N6\��s�X�۶��tn�R�;�9�Ϻo`��J�Z/�z��`��0^�3��n֋@H/�4U���&�ʙ�5�c⬾�J��k�`$�H���V���Û�[Z �꽣MU᥮����f)un��+���S^�;w�W���W&p�,���>hJT��:x.�lޮ�U��{�)��5����snQ��U�s/z.Ԣ�V[�Ws�Q�tg5e�̅�gx�m3����5�i�Ëpګ�I��w��ڬ�O[��ˇ�x4�lU�6:t��s�	)EcV��3)�t�e���U(E4b�����n��grKy7�k�V0�9�gn�L�0�ꓘe	ɐ��q?P�0d��)�IYv#B$�3j�l+�L��w>�9 6j6�]*���f]�/]e��L��z��w��+�]-�wZ:���p8:�<r��0�V9ځc��Rf5	U���t����Y�$ʚ��X���ِ6�����z�^$Nv�w5CVyK�|y���V��/jŨ�Mgd4��9�6�_Ȩ	s��+a ��N)G@��%\n�Һ9���yI2�󱕳v�	е�)٘%�n�t�_uk�F���q�
Ϋ�2+)]���w��T�1j�l��3�g7[ջIn�����uL����T5i�E>Jq�����d ��v�,%����}jY&�!gF7��m�7���i���=� 7��7o^�6�`�
����qo�Ë�F�m���^�j:I���xu�[ϫ2���㕪��j�������oV���dJ����w.	��w����q�ƍ�㈪�z��iw3�%ķ�xޫn�w���˚�r��q&T�k
k���V8I�Yk�@6b5��f��w̺����fI��14Q��cݵ2]�s��DD}j�n��ʓa���v�*�ܶ8j�Y8�T+M�s7u�U��f�e��搧��������;rN��Y��ٮ��gY�f�"��v�\W�[������ô�����3��A�0��q����΁����=�ݚ��1��Tj2#�d�IK��z�fa� ��"�f�q�J��LVF�1����ⅼ��o�}e�O��|q��ڻ�L����o���"У�0��z���< ެ�~Q�uM�55��}���V9{�Y��]m�ޮ,���ƿ0|��< Q�{ �󎞋�g~�@mv���O��/U�j�p���:�/���������T˟�
ऩ���Ri ��D��D����CV�2F\On���۩w����-���wR���r�U1�; T�*��
t�w�㚰H�&	]4��k�y�yxH��&Ǐ�j��{��mؒ�U��[w�������^OH��ΨK�.�9Բ���W��o٘�0LT4��Q`zrba��n�S��uʸK�qləDt��sB�5�%�a�5n��A����mṃ�Z�xs0pd�0bC�Gw6b[ER��B�Yj�K��b�:M�ΜҲWAs����k�����G2]'������.�{����u�ԓ�'JO"��eq�YA�.uvح[��Z�WN�i;U�0uf���G��]bi��
���t��n|���O��.�J��P��M\>���`�s�� g|i�х����6LK��?ע�����	���N����u��>��<����\�~���|ײ�^����Si
�C'�m�O��;��~�f5z�+��녶�f"ӯ�g�Y�n�n��ˢ���.7�wE;�{:�B2p%ZinA���I�b�ǹ2���ڃ�4�����ͺ�s4L<�O��X�� ��v�73�#�ym��Q�A�()��i�ӧ��ۭ��96��l�Wv:jt���̔�I�(_��h�E�P����\!P�]�w?��ׄ{�O�3ձ���r7o�|[�x.6?v���Õ�ꖎ�5�n��z��o��}�,#2�X[���RS]�Y�{��n+��H��)Ek�ꌜ��.Msrr=���>L|V�{n*�fU����l�^Ф^��%��t��6r�
����Բ�ñoS!ܠ�l�=`K���GV�~�_�r�V����biỘ*;�,�Xz�Ck���'�Pm$ o1�'o力���.�h���Ppw�2��U͖�2�Z��װ"X`ӊ�o0�o]�w߸�p�	�4����Fp�������R��3�`$2M:vyܮ�OW�YS�E��s:}X�~o�]eb�<�B������s�B����Sÿ
H!�}�y=�E�����Փ�l��ދ���y3�e��ʴ�.��U���s�F�lž�V����f*��hu��ߦ��P�L�Yq`��,+u&=.
�c����ٯ/gyB]�
\n������2aa@+����1%J5ѳ����j��A��E]�c��fޟ���m��������D��k�	�K��NG��t`�����:%�]C���a�̎���\�<�W�Ȝ��۹ZE��^w��/�b*uo{; �:��~�wp�)�t����,6j:?��&*k;G�g����[�eEϚ���Fz=|3��M��m�X��רּ�vL����/Ŗ�h��
�׹~�x�ߪ�N'��*�hrq.�o�U�8��8��]�Z��y#�w�x��W%�Nwg��P������y������3Y}��d��˝6	b��\�#f���V�3�]�Uu�q ^�]��Tܩ��-m���N��r.��mC|�w�]A+r��������=�n?�1dZ���ϲ��'���:�ͽʋS�H�0��C�7G��ޫ"�������$-Cc�;�he��s�o�^'����Xre������;�~}s��@P�e����)�])�.Em��Շ�J0�~O�jf��c��5������v�?bʋ�ɏ6��6.�W˥��w�'�޺�}2���]A�:��Տ{8_��ֈQKÇn5���Y{��N�Z�?ͺ>��vW��r��>r]����&ϗ-?����Z5UǙ(�ҜX��ftw�e�5�!
5=�Ǣ�����)��JKJGo��;W�Z��sf/k��o>��������[�/=΄�S�5ŏ,��1��xL�;��;\x�������-.�.��/4@Ѡe��6\鄱ƃ~n�A���O��jԺ�3Sfla��Lk�f��_,��3%4&r�J��s�9��K�|�ڊX{7�u�9��曢�K��v��1�Ś�֮��4���-��p�ש��o	��%0_�����ݭ�u�oTёh�ŁWu�[�ձp�+Чt�v�
=
�h���-h�������c{%��Z��-o&�jΝ������p2��O�;7�!���j�d�I��%(�еpG�̌�+�
�=6��i[��U���ɽ�c�p8������C-"��U���]AO���}�	h#��zV]d:p��vT;�NB��!³\j��=ֺ��˗�{9q�0BqҜ��Ͷ���³�*�C�8{��C����L�,����5:�vwn��os���ط�I�N�@���g�u0>Q��*�u���j�7�O����N+���y��^}fm3>=�ie�=�Z�k
�ו>�d%BB�p�Ձ	���nf��S��@�/~�R�ܰhկ�bm�w�t��Ā0��ݳG���{b�����|��k��/��eT���{�Wޛ,j�7({7[�>���F�0����k�_��P7o=�qsޟ�j,��ꨣ�#q�W�~�L�!7w!8T�n���s�L�oh�Wr��hY��f�q��N��ib[4��UC��ywݔì%�c�{oK�������
/���*G�u-W\r�I�.(f����@�n�fm��f<�&S�p�SȬ�Đ�~.�+��lR���{)��o�u�e}����&�Z+��L���l	Y�r�F0r�F��9���C�sw�@�7�J�M�&��*��#��s�� j.�*TgG^��
x>^��G�+UT{��~o�7��eaD�H���V��	K\��x~X��c� �jkŋ�5v���Ӟ��{�SwAk���9��
��o i*7�0!�ӗS/��$@��l���V�=J�-]O[u�VZ�`'�`�����d(���JQ
o�i-��ճ�Z1�]������8�'c���7FSQ*�)/v%�hp�ב���R|��~ǂzu�ǋ��s�$/��W�����|���?��z��ׅ��*�G�q}e��A��e�`|Y$�n�/�T���~,���y��o��Ѿ�.���?ex���/Ȝ�-�oہ�y7[�"r`^Έ\6Ep6ᮚ���u���C'[K�$�Z�Ic.җ:�,��진K�\�ڻ-�����m��@�����������9�6��5�SL���N��P�U���ن��톮sPg[|p�uMd��:�v�As�'�|�7�������Lp�H2�Y_c=��fW^��㖐�K�gƻ#%�gho8߳���ͮ��b�uL�o�SEa1�P�M��³��{q�\2����r�e.��U��1eU�6��8��1����S��,�V�o��Z�j��LO����7B$iڡ��]�@���%�&=]�:7C�ӌ��D5O_g��w���+w�[m����̡�׬&������@a7��\lF�>S��˕��(�7�4����Z,�h�)n<G���<XkS}is�^�o����=����wMV&-�g��Q�4i!0�������:�Qs�yE�G�#���Lm����U�	����Wj글�}�~fyg�_���He�pU ��Z���T^�RP�3g��J��[�E��w����������h01�qWZOOnP:r/$�� �d���޵��0Y�ܽ1���V�
{�u�=^��'~$6<^2�6൚g��l�������&	*XOT��0�v����맰�U/n0e���t�S�*T(��+�]��f�&[�czi�W�
7���w^���S��jdN�o��L�S�꾛��]��ir��-�2��r�x�4��E�j�%�I �"p��3�0z�ݿ��C{��᩼� ��W�ߦ-HcR�:mm+켓�<�;�2��,��� �mfb��u;�̵���a;����A�{�F���Kʍ<No�G*Nx	�X��~&P��U�����:n�~�D�P�����F�A���;��c�&��_��|�+���rzpK}� ߵ{��[%���Тf��e\�5��lR�:�h�1;	py�t\{��\+)\1���D�z�ԣ��+#f��S/���?<�![��Ѡ��w�l�7�^+V=4@��ˠ:��"���#[������H@tY]\y�J=z�
����,����;w�큼G�;=����E�A���tr4���\�e�s������V����ߖn�<K�ۥ�Q�K'֓��g���ތ_�_������zl�z�dh�pfTMϣ�y=9��3n��'7�r|����Ev٦,ۂ�ۧ��+/�v2���oHN�P����;b'k�6�U�¦qե�`H�CH}ڸ��)�W̲��4ٻ%�|�׊���˵�2ܰM��b�c˩u��a�^�ٸk�V����9��6�m�wS0������nu����r���WT}w��Aw��:ꆸ>�j�e�Ӯ<�ć@�\&+,YgW�x��dw�}�0��������MSӮ�2c�`�瓣�$݅�u��Ŀ\/�(l��jz�Yi���/U��ˢO�3�4�{��\�x��4��~o�|�-�¼h�(۫��<���g��*��/�����ڇ��.*"���{��r�sʚ�%�1{�h+���n�Um"��ώ�����O�+���[��)�b�u����a@!�L��u�"��vf�X�bnӪ0I�^�qTɳs&��Ū�$B�y�ؼ"p3fA��SX�]<�&�����v�)rf�8�{~0s!e)ܬUO'��.�W�"��z�����~�K���\��9�ޏԸ���/���?���g�	�>D,�.�\�
����禋��:e���Յ��O�d�ߧ�RY�� �=�/oϣ���v
ab���:0���8y$�0C�=2�d�[�B<�v����+R��]#��u�J&����w�T#�;SW��Z��d}��G2aςT�GnԸ�\�ǇU�u�����-Ê;J���T3���<5sԥ���v9��6�kV95s6j�^l��@�|��A����Eܯ^܂��Uo�W=�5��[��:X�����C�*��z��fֿS�3k���:�Q8&�X�b��7i��-��n�c��3ٱ�'}�=d-��
��oKmc(3��'eao�����~U��+D#����9cEC����b�������9�g�r�n�酷]��� z���Z���ݗ�\�G=�Wʯ޼�Ɣ<v����7' �����������B��K�Q"�jX��_�q��#q��1m��l�h�ʙ�ڜ�8�pAո�Tq����тE�n�ڞ�����ӽ�~�R �k,)�D�ʭ���n��o�ݤr��&)G���X�����z�t�������T[�3��̮�[ٷJ�Z~��2�,���!�0��Z��^v-�.��5�J��U����X���	�G)�Yr_�$�]*�˪�C7qj�=5���B�39���W�s�ӧ���>�ҵ,d�G��[Z��
�mA�UK��F�Ze=��,Cj^�^&��m-19�Q��Q�ؾ��@,��[�����,0�^t�dl>_w6��Ԗ���,W\궳&�4 �6��fC�I�����T��(��p�(+o�������,., @nQ���a~��H@ڈH&H�H2H� C*�B��)���=�T���K�[����ݧ�((�晟������o=^�3���o�����%�\r�A�F[���0�ӝ���1�����I��� *"�[��f���4
���\TQ�~�u���,��aN|�'�~�߇��z8��"�t�6Σf���`V���t����p;9�t�(�}ܹ{�]��d����Vc}���7���J�\;z�Ͳ(A1^E{(���3�4��m�ޔ�=.��*��fT�k1n�T+7^H1����E��ڗ��1m�.)�nfա��J���Rl�4\��B�8J$��Y�E�6�j�<�%�*p챘oB��#���<j�-l��٫�4kv�n^�wZ�ɮaC�[ڡf�j�Y̸�έJ��%(�	R��Y)h���f«j
�m�'/K��M�� �c���M䫭�J�W!��r�:hc�W���c��� I�R������;�ZuY��^"ibW�wWAL_*�)] ��#�������U��Rq�RfE���g&ḄQ�9��^��Lqd8�@͂;Nf\j��"���P����k�ݙ��F�%�vj眺�ܾT�P\7p1{���S_1��{��;�&��p
84�4�f���֛"��zwX��T�ǘ�#B�r�^Cx*Z-ȶ�il�O\�p-A6�T�i�R�"�j���N8R�IvLL�DM:��q�*p�*a���2m�"��6p<,k�h�m�l=��n�B�i(&G�u��[�1K��/[˗�쬈Ѵ)U�f��q*�cP�n�aEl՘���ψ2Јc�z���'1f!b�[wS1Ӣ�1�R�`x�L9ua˅?,'���pd�rP�F��Zʻ�ũ]L��ste�5������Ӕlv�kg*��,'�D�7K,��B��n�D^;V��eXÐ�^a�eSjŦD�:���w�LSR��&�uf�Tb�LM�4���k0*t��
���U��FuVɵ�I�q�
j�h�L�l�*ԫ!N���r�����>
�^Y��ٗ{����(�֞����!�,���{�ZaҸ¸䵦��,G�v~ i��\�)m5a +�F��Q�̼�f�ePEV`@�(�L��ϲۂY�-[;RIl:`����В��NBhMʬ�u(x]��dvf�������@�aZP���ɕv]��n��6�蕐�͐��P�El���(^�.K���5�t�'&�2l�N��x-9��g���߁��t�4jøp����"˔��و���?i�TK�r��P��]d�D+�L�V���F�9�aͭ� ݸ+l�ʼ�{ZaiL�`���;��~����ޠ�!.P�+t-��wr	��9KJ&e&�T�d\��RL��܆Ԕ��#n��[��P ��w>T2��8�U2���$e��)��P���R�Vc�]XbH�M��	YIm�U����˗�j�;C8h \��l�bk���ô�6�Q���+̄��78��GY��UA�� EU��A�  E H
���)Q  �U�  Ab ��,@�VyJ���7S�PPEdd� �+}zܿւ#>6v�K�3�q�!����ʢ��0`��,�盛R�0)uv��[��@ta/�݂����$��|�rϛ1���
��G@��+�������
���9�M���
���e6m�h���y`��(O�*~n����#G,/E��EX�n�9lOWg��QDWY�i=�f1�x_a�`�H�7��U�Efmۆ��8tx�EZ{�2:u��n�BB��%h�3-�5%��/����H�Cj�PUR6�Rl��8��"�����F��e��Yo5���5�Si�59�QAY�F����g/Ej�'5���������(+$�k5�(��}�K�
 ��  ���IW}�GL������ƑMM eR�)@*��Q)�Ơ
EUB���:��f�hiR�ٵ�BP���%\���R��5(�)R� ��P�]2�j��`@�����   �          	�QEJ�>          @^�  ;�
^�n��� z  ��QO#kT;E:ͫ&�u�:(8 h���v��`���:A�tU �U�����s�_>�` P���Z�҅�t]��x�=��h �Wn�ڍ��z��7x&�Z���@�芈*�C�V=  ��P$$=��Ӡ�9��ֆ��@
����
'�K�
Zɣ���]	U)x���J�ٙik7�Wt��TZ����{]0�G	ã m�kBe[�:[g�:����ж
,�(@�2���D-�w�J��R�-���*v�#�㔫��;l��4ր�x.�j͵z�u�#B�ٸ����ݺ�@�����ȥP�))J�U�JP�  D�Q!j�
4���ZQ��b�p+GAց��5���5J�laZ�P�J�ug�X��[fh��M��L�J��Ĭ�,�k^��B�$TT=nԥ�����J��Yӽ�H.*Su�1��&0���Q���ݺ���5f�bؚ�hOLH���6�64Q4T'M$TkE]ے�mWP  -]1�+i�M,�U �J��5����k�vu@VeJj�kd��V�؂(׽��R��k����t�j	�m*.�u�U��RD���a�(Q�:�U��٘lݝɌ�a�Ҳ�2Z����݌�[m��]uf�+F(ݺ��e�հ�gp�UjRK� 	k�Ӏ�  �]� 44�ak����l�ڻ,��5ֆ�R�rHQ����n�u��6�3��u�ݮ�X�(7��Z� �W�S����%0K,�cBg�3��(�F��r-;�u�5D��"ڌi�M,1���5��{\0Q�[�T�#(��b�8�ōP���U%�ʢ���  u)��Ui�mQB��$�
�[S��&LkM�MB�c@�ʰU*��]��"���k�h�V�mS�4ר; dia|΂Q�)\ *{
�H � EO�0�R�   MR�HК�觠�y1��O��%*�   ��F�$�@   	OB�RT �4��=|n��6��o��;z�<\��Y�\��W=k��z�[X��������g�uO�'���?��C�Y�^���B���_�D��HD��HHy�"C�i�����i����\�tސJ~�
c?���VI�����H������:��P��`����v��;0�t�:���D��?�Dʐ)W[*�˹X.;�$nK2���]�E��jKTK.�$�ĩ���g^�������V�cF�*�f��Y�tM���V������� ��YFp0�ܻ"�nv/)��$����(���fֺ8K�K�U�tޖ�+#�d~C�ާ'��3=9���DRrZ�@E���f��rnX�hb��� y�K�:��J���.X�+/�R��c?S�\%�Ԧ����j�w�m�x]t
-�K�l��B<E�i-���cn\�2�h��̱.�7Ч��6�K��Y�&��t�,j]�1R����@���,�Q�Oi���.��fV��8��dK�o��a����ͷt�Õ���J�E�=��:��
�2�8���=nn��r�GyF���O'u=-�0���� %��M���:mU�>@���̪u��ús8>�BIU��B��c�"�������3��-b�=��z4���j�{�=�~C��D�̇
�8��>����aaqv�۽�[$�����u�:ݚ6���\��|Zl)e��k�zJ���U;����u���e�q6�̕�0��;`�-�#�+U��m,v��?��H�rѽ݈��2u�����kiVbcIG�/���X[tQ�t��)�|th7H����ڻ�+B���c٭>Χy�ɾ�ݩ1��\�uǆ�iسY�]�X�*4FM�p�Nٽ�xn�4�L�rS���70�y�d��E�&ʢid�\UH����{��chc���D���[�fRsn-����2VK%�ğ��~�w߿}o�O4�����^�������d�_R��|����������6���/ENE���Zp����<B�`�/��GV����D���<�?e����<e�M
M9,ga�PSȕ�9�N3h^�F�]Or�:�jr?�]B��^�������)���YHvv���d�.�Pͷ�$�S�y���~�8������*q��x��I:<��p����z�@����p�
q�8^(��'DQ�����O���Q�'"? S��=8G��d��zw[�64>�]u&�a��j��H��e�z�y�wki���JZn^E���s�B? u]���b)���Kڳ%�N7?G�M�?#�i�1�WU�:�܎��v�7t���c��4�X_�=���)`������S�y��u�ΰ�U�$u���V#�d�'��``��PM�V���pRǑL�.���,���m"N�"������ۺ��P,���m!�]��%�+n�	.*)8�]�Hm��,J���q�RL^\�x>���i�¼/� )�����~=,��e*�~ͬ��.��IV#.:h�����g�@�8�W���	)��T#��r'xOgC�D�/�)���Z���Rt�)LDC�$�=��C��W��T�)ʚq�~N��w����(��:)��W�y<J�8��<{�O�����q�8S�8���8S���Ӣw�D������SC���܉�t�S�'N>�S��8�8������d�9<{���=gt��'�
q�> x�T��p�Rp�Ā}@"��^���x�x�~N?'����#�O�����S��N����<>$��P�'=�_�8�����q����8�ǉǩ�N2p�=ǩ���N=N"q����!�ӆ����&7Y�\�A+z�9�&[]2� q�Ֆ�]�Z���ucج�J\�'�'�P�Y*Uͬذ̲:��Rv�V��sڱ>�Zδ鑖2����-�1��|�lX�2U�.+�(Yy��m־���z�.w�BξW03?$��k�rw>ͽ�P��_\�pu��Jj�r2�t̋
̹ �T6��9d��E�pE����S���$�ثy-�ml��v�l8u4s+-��	Ŋ��w����d�I/5���2�&,�uLuͩ�@~�'n@� h�H�\ �<��I�*���k3C�F�ʘ�����)޶^��jm�;��r�ugF ���یc��0�rr4�mh�����n����(Xɺ��b��2<�cj�u���*�mҽz�p�����*�m�4�`w�J��n�pk��I�C!)��T^�t�F����Ty�![�0��{�b�&�sqe~FS2��f���م�l�6ىA��u��^�D��*Х�C��쪥�+�cj�����r:oR�����fnԃo�GV1��k���̒*��;�f�7x*�73K�у1�/!��2����oe
��Ѻ?�aԭ���9G�҉����[�X�q�&�⮊�lV����ԁU�՞���� �)���$~��� ��]Y�&�r���;��_�fՍ�Rk$c*��g0�\ǖ�5�`�q�tk@2�Q�kT�SX��m77l#�"�sh0���!��%";0��Ih�y�ҍ�*�
M�ʷB� wV^8�L�*I{D�Q�F)��6�̓F��a���Ż,�Vc�X�cN:e`��i�i�)-�xN�m���&���������:�$���7���Qt^�Xo"��Y�6�J]��%mfM�Z��`��U���E�Â���5���5(���@ �l�G6��?#��,��V���-E�<�e��,�AƩV��N��[yq<7-�qȖѷD8*͖e�&1�n��y�ڰ-���5��d�S�^��xq�	���P�jdt1�ᙗ�C6�H(��HU��e::��AY�� �BT�ܭ���n���U�7{5[�e�O�f�9�j��Zә���BD�zI����e���L;b��ɼ�Ӂ
:�&�L�sd�`��fMn�7J��gM��jU�� �
w������P�*u�Ojn�b�D
J�f���5�܈��1}�����.���+a,��r��o3��ciӽѺ�`e٨2d�]�8���t���$i!<v�lق��^D#
��65e��Wq+E�bjE7��y	0ӽ�j��G�&��bhi��0R�v�Mw�匐�5����4/5މTT�ɠ��[ L�z�BQ������#���s�y@Κ��&k9��ͼ���T����M�E^EJ�X'�D�$t�U���ۈb�v.-��$H=u��FA�Q�EY[t�L����+N\���9	{i��^�V�6i���Q�5�x8d��E��r��(?ߐ�o�ۻ�q�8S���ǖ}{>��l��mSt\�tI\��h`V����ܦ��i�V^+�(�y���m�M�	�{���Ο/��o���Zsqd�RS[�����j�uŶ1)j4q�XY-]���QC5����G��J��ǵ��5N�v���KF�õ��7M�w�$��̅�V��1ݭ.c��[�y��`$n�	BVb��,c('��N@�����V�w�t¿a$50U� KR˫�4�lA=t�n9y��p1�,�� ,:JaV�R�uy�$���u���%Zr����ɕ�j��ݘ$�Ԛ�*{{\$e��Ы������ 1eF�BDY%~-Ė�r�4��t5W+@�̺+wuA�:X��A0l�7+a�����gr��0����f��錣���'.��vl;%<�9��6�t�W��YV�w`�{cZ֡Nʏj8n-̱p����B��t��xԪ�TکZo1���ER�J�M�`��D3v�l��6&�~X��yn]�m���q��aw�0i�
(7��1]��'e̢�1�cWm빒��:�3
1�uFб�z��v5���*S.�!�)�e�����ZHL�6\ܲAb�EQT���+�rS����x�S�)����!�+ �ē��'h�6ClA�F�iʡF��`/����p��6n����h�b��y�plʗ)��/��CQb�)n�!�U/L+h[���ST/@&�Ӥ�qIb� =[��d���Ĭh�7Z�ִ�ꥊ�Nc{q�c�씱���5W��� ^��)��>�8:�v�N,�v�-���m5;�<���h]o
���'8�q}�x��{�X>y{�I*s��}*i,�����Nb�Q���|���s�����O�u�4lY���w2fMގ-޹�N�vB��>�E�fģq�����*�
�)��e>��ڪ��÷����bVӁ�:��I;�T��M�ٽ�p�� X�Xj)���OC�̢'M�S�wf-K^�q��
�j2��R�m��gPͺ��tҽ
S��*x]%�6m��ݔ�R��x����o�e���oY���Wr�>W&knl�h�r�<�_��z�i��������񿧎��;`��T�[XmJ�X�x��nu9��}L�9�c�t��j;K+0�\���y�'7�Z�c��Ԛ���rn�P]�Ngma�618ˉ]�l�h���c�"��uU�	,j��L�����z[M��j!�N�<��F�J��:)t��6�@̲�n\'�3)d��T�њtk҆ǱL�+��`�Uk���5��B�^;�l~@�B�V�D[�Rn�!PY�ɓ�y���ûѕ
�,UX�#1�DJX��8�p�V�ӡ����m6����aս�02��u��FXܘ���7nMͶ�ͻvpY��*�nm�z�Ӛ�X��RTV)b�����:���ƥT��9��B�#�w��R$�'!G�E�@F0P��'�=�~�{��`����r��U��5&�� �L��Wg��S�[\�D^<x���9����?�	V�,���[.^��Sx�ͥj��e�O�V���H�����i4fY۪*M�t~��? ?R�Jn<�x�Ǻ-x����~���Ͼ}���S��U
Ԧa��,�0j�l�q�m�̷��͸�������?�d+f�����x�:P�g ݸ����C K2�Ry6daw��%����V��z;[�)�G%M��-�fQ���ei)���+�41�Fh�	�X�
���)�(�	y�7v��0l�;"��.����,?�]�ƶY�:�C��!��$$��6�:˫D���M�I�AE3(�6����9��??��,�;٢a�;���Úa85mM�s���kF�dtD̽��s����Zͼ�Su�6�j~�Z���3fT���p\R��԰�št}�2� �];�e�w��`(�+;���b��XHԓ��;�W�-�4�Ոzvi����t,']VcK01r��#�B���oi�6�e2�^8�P/��6*�,��fŲ�h�T�,��%�-opm�Q���-8�*L�����	D� R�SRbqeu�t.�ri�,-d)V�ҫ�,�V
�"�R��u���Sc�/L8��&K�5���4��#�8��fT!�(��# P�%�;g���5z�&]7;�st޼��,�mYљ��	�(�H�Y�p��R�����
ҩ0n`������L�ܥ���b�-����pP�9�"0)S�t��Q.͗�K*� #��N�C�]�K`˩ѰmQM=���@���ɒݔ�`ҊG6�� 3�ן�O�����T}23vU���nl�s �I�u��r�a�t������kxF���Q�\I��%��������5[j�F��f,��ȭ���Q/MG��5dT7�{j��yS���6�ݵwĴ�[�4�˼x�bG���7^ʙS�b�"Mv7NY#�%�}9^>kV������^6�9�D��z@ڴ�=9U6�j���HZ.�N���BUW�D�7)Fj�*�r�"3e�`��͖,��o�qӷ�u2��v�e$��2���A&쫕[�r�w��	M:%A��lf��2�h�ר�G$���e[�H�k��#/w���NTѧl&�)�&�d��jT��X�5nJ��Q���2����7B� ��$�$+�X�z��d�г�P7�2ʃ��)2���x�qq�@��u%Vr�[­ʷD�OCN�/#���.�i�X��z,��ьh�UחF��S:"LSM��;Tf�A�6aUq�%�W����B�ZT��y[x�%��2C�z��̷��R,�b{V)���i���9� ��*c2V4r��4���f]k�0e�d�Ճ�0ɤr+ʘ��7ѻc�gln�S.����N��bC�	A8�'��Y�U]�/�Q:W�B	ʆ�r�u�\�s���N
`�e?��0#�v��Y;�a>ie/ȸ�����v��	���[��1rm�j)���ߩ9�o�w�̧j��,�����M�G��kv*P	�i���J�:ҫy�3Z�kT'E������ܼ�T�N�O7��!p�Ꮀ��;V�
�)!a���r�lUM�3�ю4-�2F���skm��]��Gk��md�mm�l�U��m6�l��۶�m�v�m��Qy�7�H�I�#}$o����>�I'wt�H�I�$}$�����7�H�I�#}$o����>�F�H�I>�I�$}$�����7�F�II#}$o����>�F�H��F�OUm��T��@��I$ I$�E ��m�4����.�m$�m��m��]��mKl�1��[i��m��m��m��m��m��f;n�[n�m��ll[n��5�m��m��m��m6�cm��i%]��md�m�m���v�m�]��mm�l��km�e��m�ͷ[n�M.�f��m��V�v�m�$�H�rIJN��8���Yur8�:u��)l[�>&.m��*�Kp���<<�y�Zq�E��w �:�)V��٫pY�)[��DJ�=�LoS��.s+WA�N�jY�eL�er6���ʴy
=b���X�2���'U�=��^�ʘ_5�fV�.����&�q��c{���Q���;;�.]q�V���o=CJ[�0
s�h���6�Z{��v�5��FK�b<�ռ�7�,�W�:��SA3�n�,Q��kIݥ�w�f�����)bN�b���c�&R�2����5λ۬ڼZ��6�3Gr���0���vv��;:������l:�i��O�̔.ؚV�i��@�A�&�dcnz���,���B�d��ޚ�h�?p+�����wG0���?�&��d�*�خցj�s���g*B%�wǸڤI��m[*��aٗٚ{Xi�{�ѡ��cUr=}Yy��8����r,˭opQ2�;Ӓ������,7\X�����{�s�M�,���z��N�78=�P��"�����.��+����y9�ss{�^~��_��} ��ݏ�A+��аAS��s�NLk��6�������	�:�yAr���=N%���j��*0�h�K6�!J��ww�k�7�pF������=��V�-ִt�]q�c9ف���5ԩ�s{����mE����m��p��L�m�Vw���"z�)�����@v�����hgA������"�#|�a�g��{3�mr��d��T���N�q3{kE^��"2I�w��ό��2$�n�����V��[ٔ�q�΀�h<�8����0%��n�����݌\P����.���k��j��>Z���&)Eh�@����"�o��4�;`+g>�z��l��,�頖WVo��<9�<�n����֢ٻ.�c�f`:�`k�������Gn��O	ë����]{;�ׄᱶ�է���o8�w��]S��bØ�qd;	\t�S�u�	u��1��e=���+���Q9:����q�s޽9a��[b�a�yo*���1	�S]G�����C!nJ��q���]件��*]8X]�	s.���5p�!�i�vǖ�G�4-�nC�w�P����N��`�Ν;d��6N7H��ژ���9Gy�F�6k�R��Y��7��1���Kn�cn9
1�x�S&�������n����;m�b-K���yȠY|�.��	���k�e*=�Dr�u���0�ջ@>s�t}(vC\5��5������(V32[Z�Me�+o2��ɇ\�ѳ��;n̝\h�1�徵&v�
��3k���LnX.�q.�����ݧ��Ym��M���:r�������4���@���Ts�C&����.=�����+1��L��#��z�%���՝γ��-W�8mTEv=l���n���Y��%�B�\�^�Yg/-Y�$�Jş��Շ�v���*u�ʺ�0Y�����;�aq<�8�')��[25��Y���^���)&���Z���w�:�o{A�")��l�D��ч�u|V�γ�j�w��x������6��$����$Du��o��G4����gFlɌnۻ��u�X/�^sp�|�֍�hq}�$�Ev�/��O\d��i��rY�g(�Y�N)R�Ż���'MYPT��o�[�3*Ն�;�hs�S�e>�;�o��x䏻Aï����3����+�����]�K9���G-��4�����x��骹��ra٘I�U�b��)="%˩T�������=�<�d.��B{���O��΢7�0Ex˒Z}�T�!.͔UkX	���3�떢���w����R�ᇙD��u2��t�ھ��Wd�ӝ�ǚim�Z�)�wBV�Q�hqsh�=N<��Ho�L��tf�W�͇p�ev��
�����U��ޘU�ߒ���Ɠy��V�|&� �-���"CIX�՛�yYI��"���V�d�����\tʊ�̄������+0�s��j�5N�W���f۰��au���}*&�-��c��$�:�w�\�Y�0�����$2xu1U�eoG"�:��9��6l��p�����b݀��E-���t��uAR�[��r�1a����.%;�ޢ�.[�;�GY��TT�3�Y��K�1ٿ�5�3�aC�']]��Sewqׂ6b�Tᗐ�d����
;���i���s",m����X��m�=����ٺ��ě�FȦ_�n��2\��X�)�yח���c�ft&�Y�VaTH�ܛ'e�r��+��Q=��W+��])ul�,��H���hDs8����v�o!qO���ꌿδ��z�J�Vk����Ms^;�f��S��"1���7�o�,��3�
RA�zU`��4���7��'L��Ƿ�
ۻ!Є��sX<����xٛO��0��k:F�6���ۭ�[��2���x�|�`�6��V��0�e�z��V*�f�t�to�u��qڅHT��>=hꀍ������im��]��c�Ok�)���g�b��;� �s�Po롎nE�xXg�ʾ����\�8n��ُ�8�SK'��^.�:�I�o/h�J�o��:3t!I�͘4Em���TsVK��������������zj1V1���ՆZ��6�+����&���1/�5ˮxa8F��<[n�f�6bԡ���_�F��:����)Z�qh�f�Z9i��i�"*��P�rlq�V��`�B���Y`��k�y�Co��
s��F��,V	�iҠ2eZve7݂3!	�æ��!X�W�q��wv�b�D/�iS�.
��J&�dn �%	���CT��4a)!T����mAA��	�����9�G揮�h��l�6���̶@��C�<Űj���V��!*�\�	�-��
�'�b~��3M0S�p>BHڦKS��	���YY��0�~�.j��H�qq�+�U�#&ݺAJ�M�8�d/��Ի+a$v��*��2"�U(""B��b
$�BB����3eM��<|g���˥"�1�п|���I_-�&����auĭ+t�id���h��-�O:�]e6G��|�Ʃ���$��\��xxy�%�[��U������!�i�d�g�|�^s퍦k��Jg)�F�+e�dٻ$눺ɤ���o�����G�o%��f�u��t4ړl�ԱE�̐���@��%���c�+X��ݴ���ʏ�<,]�O���Ǽ4ٛ%�m�0��fy
U�X}���3�Q-��_mw�}�O%��a����W�盲yw���*���� ��6�%������E�F�9٘�Xk�{���E݇Fn�?�$��em�cI�[!n��6���m��:H�_m��$��Ķ̥Ѳ5���ı���J��u]k��t��3��F�p�g�W]m
l�Y3�h�y��fA�K�By��?Ϟ�_3�7]����F�c�4��L>�wg�ڒ�H�&�a]�Xm�u�4�7b��Y����2]r]3�+�t��ơ�.��p��ġe���Hb����|L���X9�ٙ��{'���Or^�JR�t�6�?�d���[[�tt�Yq�l��N.�o!�Ә�|�Xxj�9ut�md��WV�l���,�*V�I9�4%�$��fѤڷd�:F������\��5%����n���?xK�:�Ś��M.YT�u�ns��Yd���k&�cX��y$|���/=7kS}��ꍊ�N������y�D�����k�݋���4�xX�ϛi���l�a����]t4�wnl��16�-�NƺG`�˝vٛ,�\��Ik=e>�_'�$7VG���O!����u`�73;Y��O)��ZX�y�������YJZ]���e+���ʛ����S�[�%��bc>xyb:K�V�vE��X�&e�&؝knw%��0�t��Y��#d�t�S&c�������,��7��yhG��w�󩽷E��1�3L�l��He]�ǎ<�԰�ӕ�?|'�xQ�#(�<bm&�D�u��W-���9�[��]f�ˢ=M��0��������Ǽ ̕�m��&MZᚰ��L|��3�:�g	�e|��DY�/�����BI���l��^���q��G�A��[��Y5����T�T�ڗV�I�Jݝkm�Lyv"y!m��o��>>��J�0���E�k�,����4�LW���/�x�d�V�>��o�eU��x`�0��#"�ř͚c�3�V;N�9��m���d��Y�5fH����R٪��0��%7k�a1{�/��?=6�����(�!:����lx���,XVv�,v%jJYJ2��њ�6�oN��um�7n�j%�Um�Q�i�2I5In��El̪Y��HO\�u�i+qs-��+-����/�u|�o��]/Dnͣ����Itkf�wf8�`G`�_���e��7�#Ϟ�et&�#&�3��E|�-��>�W��m���D��'mmh$Тɲi9�j���kn4����6�[�t�9��Җ��65��:ݤ�al/[O<��|�m�q���6nu�S\i�f�v1J������H놚M ��&F��͍��Ԍ�j�zV���cJ���є[��۝$�#dI�ߩ��I<[/�;C*�k	��J�7cQ[Y��������u�?)���G[�	v�IKm�C3}�i��ih�.�Ѕ���c��}o��6X��ĕl�-�-�E���j����e���̺�[0�4YV]�jm-S,�Vɵ��15���2B��i�-2,4�ii��흡T���R��֭�d�*��[��-,)R�nVY`k%��r��.��Ft�:mte�̓���И�릚[�͢MnQu/0��.��2���UڙJ�.�dͅ���h�JM��IQ�M��6����]�6�ok�6YHhɵCA�պ:KY#1l��h�
Ɛ�p�YG&��ֽ���)t���j�E�#�͚��1�\fi�ePp�u�*E�Y����:�]�k�e�&����[���kGK�h��jm�'!�n�[v�$�[5v7ll��mR��2�q�h�z����k+0�J�!�Sh[��Isu�K��&�M�Q�XK�Ε��Ų�v��J;l=+k%3����Sm�ӫ�M�,�e͉mن�N֊Rٳv��^Y�bv��l)wLC#l�(����e�+r�뙤��L6�H]!F�W���k�ɳHW�fF��uD7�UM!��iK/���(��t���n�(�!���Y��e܊WY]��w\;ZSI_WX?�AQ�D%��M�ahW��J�F�Qv�5�Q���W��*�eZc�\�Nu�5˰1��pe�%��Ộ�]���ꈕ*q��o��[��_\�<:����tܻ��q�6��Z�^s���B�wTnVlK�-��o��緈�4�F��%S*��L�ŀ�� F����Xi�ͻ�5���1h0�z�9�Vgt"�ĺJC8��V:�u��A�k2ܴ���V��rci�$�%��Ȗ�Doj
9c+LU�Ve�/
��]9�s����i�{���B��}t1�uN��k�|"�,�#}�9��Zx�Q+r�OX
�"�vG+��j�a秭m��Nݬ5u�P�-+"Ƶ���Wpes�.�_'&��K�Ñ�s�Go{^Cc��Ҕ2	����v���v�=����-�-%H�'M����b��8�7��,��䬀�$��ޒ�*�E�$��N�a���O�4��9��I_q��32
��s	� �î�I�so��1/L�z!�e�+Mf��f�f�5^����Q�=D�r+ǔB[}�N�]Qq}{��}��rSk+6��k��Aj���g� �u�Hy}J�t6ԭz�B�C����.���.�!v��:���ᬡ55�Uk����|�U����O6���v�5��nH-���x����mfb�`�ٺMT�]�0��0�FKctM%^qZ�ǽT�֭5��֐�j��h�o����<�%t��ҭ�ޣ�lv�N���:�X�c%�Ť��[�*�T�}[��M�24U�#v�U�N�9�X6m�kkO]\BR�)]��c����"U��f�k��Y����ۭ6!]��-r��������spN�ќ� � �x,����7�-��..:��{}�q�q�T$;�P���K�"��4�.�H�rx���Mr�|	i�K|�H�[��o�Ux�Mp8��+2�|B��q��>'�q� P8�q#�����8�P��8>&x�wwG��P
�(|C�x��|���#���w�S��;'q���
wz�uC}���8�q^���8���ߓ��4���ǻ!��������~x������ԯO��tx�^�wx�������;�'������q���;���;����^=���pW��g�L�� �z����
��ë�
������p��x��	')�'G�5#�w����<y{���;�W��?U��{�=�t��?<�T�x2q�����[��;�'qߓ���T���z���vNʜ�	��E�S��ǻ������/)���k���o`�N��u�*��G�Yǟ=��'|�R��@R<�Bs�^�d����^�~ӻׂ'�a+��M�w���'o�=�I;�^>�T��=o�߉��3�5�N>=��y�yJ�C��;�ާ�>?����}{׌�����z���+��|��gה�&{Ǣw�Ǹ���^����������)�P���^�G�N�s�:��W=����N�y� }ǅD+ǉ�����?Zd��~N+�^#؟
H�R<���{�o���g���~<���'z��;�Ǩ���Dﯔ�(}O^��T�^��|�={�!ߞ�װ�W�?N�>C��=N�{��py�I�@��~���*���ND��`_�<C'(��I�J�#��� �Ǹ�W�v@"[ o��<���wT�@��'D�	��w?5��������^�?=���ߚ�2w���'��d>=��^��N�>*���~Cǻ��>y{�O�8>!��\<^�P�w|{��w�
���T��<x<~'�����w��>?=�><�!l}��p�����������*��S��"q�#����#������N�g�q�N�^����N�w�'$C��q��ݞ��^9{�I����|���'��}��${=� /P���臒p�S�'q��!�?Y�ݞ?'G�^���C�C���8���'W���D$�����`��q���z��z��Ǐ���C��ԏ}���~�q��q��&N�u���w����{����Ax����2z�9H��9yz�|�z��=g4��~N^����S�$�@�}�^<���{���P�����,��=N
�L�rw{'�tO�}@+ܧעr�糃�#�w��}�E�"wǻב�C����@^�iS�Sǌ�Ӻ<��D�����Z�z����������w����q�N��p~J�ϵ�"w�����,��v{�<�P��� z�T>}�q�3�x(��w�^�x�N������z�C��;�{�
g�#�����N�����<z�T��O���7�<N��P�#�{ |{�z�D=J��t_����~��|@��N*/|{���QbyB<|N�@���,��w�<��wǴ��'|~���g�׌�G�^��8�x2yӹ�&�F'�!�������OZ�~J���|�X�{�!�����1�C�?18R=^<'뒏�J�����+��~x>+��C���'x����:"���jY#������"r����~�w<O�}ӿh������d�N~\�I�
�8����_��X�"
tI'A"���Io�w���=L����R �@���>��|����{�_��=}W�R���w�_��>}�x��/��ߧ. m�kg19"�#��F!dnB����}N����_~~��3����5������O��}�<z�/�#�/����>!^<{�1�+����ʞXUx�vH������.�́l8�ּ�/��x��Y;���~H��;�����O���
z�yN��r�F�=���|ϓ�T�oa�!��S�'����>?�;�q<�+��~��/��C�W�~K����x�B����(�x_�|C��w�~����+�⡴=��,��/������Ǘ{3���޽�S�=S�<U~Y��	������z��@�3���(���`?�u��9G��/|����|�{֥{ľH�8C�5se�'�rT5�FH��5rI��T��_���>|�bC�n��C�a׿'ǿ>�ї҄k����߱�߯�����<����g}zY����B��o�)Qp�(�w q)��q�s�q��}x>!���?=��Ogv���Љ�{ +�}J)��z=^��N>��y�$O_�;ϐ
�������ߡ�׏��|x���q��~@S�{�>�t{1�Ϗx�d�w�O8���;��d9��  |N�����!�G�x����ux>'D��d����q�����S�ǈ<[><w�8B'����q��zo��d�S�'? ϴ8�����gw}x����S�'}}C�bwW������� ��82x��G�8�}`�w׿'W�`q��ޡ��
q���)�^+���<wz�S�� r�C�8����G�t�d�w��^�Ǹ��W���P���^�~Ï\�(S�^*w���k�����^��DHw��4T����}���Ϳ���eޙ+'u��/n6��M�G���y5��4�x�O$�Ʊ͑,���L���cE�=Ŏq�G
ۭT�1)��/����u#�	�9�ZD6��hh�2�d�WdF�((��(�{�݃�ҳF4�����*p���A�&��
K�Q�j��՛��=ţ��6rRQf�k3�w5�n�
�u��머�(�t�7:�̀�܏-5��H$n����Z�L���TV�!@�!���,�-K���W݇\]Uf��/7;^�$�+�[/�;���p�3`
f'�{t-㑬���̮	��eͰ�-�斗ȳ}��6�d�^���Bj����G�s����I<N���2�T�莰��N���gz�NVZ��#U�ǧN�9�	|2f)I��y��m�����_}�^���X��Q=����9��l��a֏�7kL�_g��5�9��Q�;���,8; v{��ߐ���m���s�����	�-���x~�>�w�NP��?��w��<p~�8
�z�9@���8#ǯN��~���W���_��W�uUW�ɗxhy+C">����"$|����"��W={�$�"��iȈ"i9�U�T"wD�PS�D�ZU�E�=b"ua��^T9T+Uy�7������|��G���B�E{�QA�-"����0eUQU�S��/+�(F>�D^�'�_�G�U_dy�Q��ofyT���@�Z"
����yܼ*����Dx^TS׊������;삪�<���#ȋ܈�	�/"�o'PU����0E��8EUS��TQ0Q;�PG��*Y�x_^�XA7ȓ���U��*q��V�|$�?(?!Q�^T�l��B���#��>�ʀ���"����E�|�{�~�,�*�/t��n�Dy�=>�#��:i������@��qDFN&�I��ЅO��2���y쨊*���x�"��lEyt��aV�}�k�G��UF3��PD_��g�>�(�5�YG���������y��OgP�Q$�
�����{���������/�}���x�����G�UG�8��[��EQE
�O!�G������U�NDUT^�NQQ���Ɂ���uEs^E�(����Q�^�k�����;OlQ=�v)�^���� ����֧���`H�PA�c�>N�{y=j�^�U�Q���瓒O�y�E,+f�� (�AR��Y��W���?ȼ�����A�D+ӑ������g������f��(�O|�
�1��T����H��TP��D�'}H�DG�}z}cܼo�>��ͤ�'�U��=xEOҶo�3��o�$��H��j2@^	:��UDy�t �/<��D���������#�(�I3�,y~���5u��g,�ڿq)Kt���L��m����|����+�yz+��~��Ф�����-�:�|�<��~��QQ�O�/��?1��P����֢���&b��ǵ"����t����{�����xX���g��6�U_Y��@�v{�I���P��[G�!�{��,*�%���ٷ���D"y~'�{��Ǹ��!�{��VB+a[�2Q?0�^��*��_�!���!E��<�+hO������՞K�g�gCN~P�Ϟ�?<�����T�?�ϟ�{��D��I~~��	d�QU�7�&{}X�^]f﻽�����}֩�����*�O��+��!����M%Q�$�����ó��NW[�6�A����+�~{6x��r`bD{[$��^�G�����{֌�$�7���w�I�X�S9U����Zx>??��
���s6�p�+8(�	$!/!q,2"R��b��\��Wx�2g�}y8��,��i�E�
43�2PA��g��5J����.W���ԕ��:{*�}�z"K���7k� �t��ITh������zq�7q���!
�w2�p��P�8=OR7�6���X9�}MHWk?���B?�{�>��j�o��y��&&֎��Oł5#
k@��IDL�Y'�P�ډ����O�D�w.����;4�ӆ���=�F>[�?G[os�m�{�Xf���F�s��te!����K�!�j�ޔ�nu`gy>�R�2A$��2��\�+7Yl�w9V9K��p������'����\}�<��=��ggNî�Gͅ��:65t�7ҥ�b��8k.��ӵ�&�גj�v���d��������T�a<�4.��)n�I�ծ휶��5����ټ���V�̼��d�K�SO���(���������:~`���W�ӫ��Z���m$d�N���~�#�}��_�Qc��DO�%|�۬L�#�	�����={�z=�A�����T�7G�!~ R�϶��`WY����甆�B1�e���۞D���듖y����)��x��Ջ�?j�
Ә�n����]'<�)����-����I򗿿�>~�w||g��� K�$tO�c�;���ͥ~����A�l?���:�S��E_�oT��qJ��T�tH�9���|�}��f��*�B6�DP�����B�(j;�F?.���iBKN��Ǧ��y�6��������rd�J��������*$ڐ��.�'�'�ǘ�m�h
�fE�'�}��O,Z�U�`A�0>Ͼy}����r����Đ[��vy垡����(�"��*�&6y
(&��-���<-���e�W�/7�0"���ۯ�c2�'ğ4��� �1^�A��B�h��g#XWk�H?~߻Ǽ��痼O}�x~��{o�v�l���mTX�<4��"������Ұ���-�HfE't>���>��OZx�_���}O_$�eV{:��QF�Gڡ���@��JA"�byg���=�ґ����&E�'��WW�gĈ��'�-�}�4���O��4��#���4��T�����h�@K���0U#͖�Z���qw�� B�3}��߭�v`���$���N�Aa<@�~�D�EA��24�R2iӴ,~θK��<�*�2벻����3�@��m�A��O��1y�a�~E݈��I7?iE0�:����܅R��_F
�jd@���=)J�H#BY��L7���o��3(%�6W4�{U�B�����G�+B?��Ȥ=� n�������4�❖W� �l�$!l�D(�p�׎�2h�����i��ix����e� �_�)�>��\r�kd�h Her����%�=g����A��Hy,����|��i*	����ľ?�F(��l��y�~�4�!%���Z�d�Y����w�^��(h�4��ؽO�{��.�r����M*ƶ�=-6ejޖ �:��0��N�w9���7��r�;_��A��[����VR��K��(��*[ѵ!�7f�ؑ��#�.γۜ���Mr\*�^M��J�k\�^�?v�TEy�n�d�돺�y�qC�#� 1��!��^5X��~����N^�X ������;�O�K5A	E)�G�T��x�g�=|��������*���<�y颂���h�T��N�!h.��M��'}l4Q�w�^?��y^_^>oo��ߘ��{-^��R�L��أg�6P�"B=�R�����ʱp6�p�eS�����݄�İ�w��d�0��D���{��x��O$'��4�,����G���N�hU!��<��Q�d$��P6�&���x�ԥ�Vu�еw���F}���Ǐ�X���b��hž�)<�tD��2(eQt�?��Er�S^�(@*\�H�rk�i���N��l䨉Kd�İ�Q��m�KY�����w~��#ύ���h�
]d$s��X$ W��\�'�Oѥ�s�s&� R�g2ͫC<���`$�H���a��K�pBUY�7��:Ld}������c�P��tA߬pO�W��׊?�TZ�׹a�,�T��6;����_�O��bV���?������#��ĉ���heIݫ������0�BU3I?�x���C����$RA��F�/�!3m����.��|��$�
O[��1�
�W[:�)=kh�o��{��n�uW��QGq�=yS�0偂[���:��	?����f�@�_u@��\�=����+����
VP��[��e���h�y5��wX��^۫���:�M�}LQ �� ��)��(b]��4�Q:���Q��e�I�\~��wvn܄��%q�������j�.چ4��a)����M)S��?6��v$�~.?E���Pd�~'��S������Z>i�y�rԈr�Ui�������L��J����i���݌�^dZ�ںwD�(��>�{u���p�3;4�E�;�A֑;���k@�^f�#p_	Ch�`���n��{��Euo��ɥY;S����X�Fҕ�d*5����ޱ�k&�e�5���3l\��6Lnmvx��7�`$�������O�����Ŷ���������o���D�����b[C+Y?��\fD�����Z[�[�:�@�(I�$���[�-(R/5�|E��<@�j�D�H�x�����aL���j�R"+�}�0�@�U�,JK2��q�Kgj_�����{׿�qD%�C��t�A��@E��c��q!�H�J�L2�BEfG	8�� f�=�/ɷ�Rf&(��v�M����aĚ�X�S=��{�5���?-/�5��O*�Nw�gdEJ�c�yk�9�����횔��_|�0�xM�-ߝR�l�=�\s��Q>�a\Nzz_g��Q���@y/[v��7�Ŋ��#�I�!��
?�=�D,�ސ��{��B��GL���$Q����O����ȵ��S����yܻ^�҅V�1;+b�uj��r�x�#�
VI�)��#N1wۑU,������G���L�ǲ�l�8Q)�Uy��}��n����@w��e�E]*��f1�L4vUvx�x�i���K���]U~'�⛿�S/�4	��2��4�O�t7���/���90�M#a��s�+[���|���;����d��VDÎ�Y�����1X��4kmj
[d3��:��3H�D��Z�a<��<��r=밗��LY�W7r7�+h����ғrϗ���8� ��~�B'B�e�J#
8���8 �#��K��I~��IK�j��ͥb�*����ˊ�=����pOOV�^���Oɚ���L��҅,�d�	��4��N/�2�f/��$r��#N~E^�wS1�XU�[w��H��x�����Ը�s��w�Mօ�C+F�yjӉA�u����_]ƃ� ��r�^2�񊝚yM�v�`��N���,���=��L_i�W��<�>��
����!�Aɭ^�;iU �4�L�"Y!�N���K4�؆*�H"C����eԫ�nvu�u$����K̀�$$�g���BX�i�L޸��8�%3n{��W�<D �h&6̜�QL)g��F�#D������~�RK���ݚ�.{���v��$ɛ\���v�]l����6�&�e*,=r/��xEۢΝ�QV3��wWF�§g�HJ��5����9��2�4X2��,˄���g��^ ��eP��햅[U��U=�q�ɤ��Wg��rW]w^fE�b!�ܩV��r�n�J�㒐���Iy5��;�"��A{��HЏ|��~Uu��YTyt��䎪��|K/Zα�k��!Ti
p��I:�!q~���#��Q�XA��y^I�%W�m�� ȫ���\A(�L��&����Ni<��J(������D:����+��ۙ�ͩ�NA���-�h�����q����%�q��8��Q���Je�u�~]��|C�)k�=@�ř�~q�-��/r�Yq���m�B^�2Pș>kR�tj�r͐�<S�<g*>�H�5~�`��[�c(�ŌB��*�$�	�ˀ�L���$j��׽�ٻ��ēɵ��]��G!����2�;o�;*� ��t��j�Z�T�-Tf1w��lƦ���NjF�!6��9�����=W��[�K��]��!"��%:����:���Ӣ���^b����\�ɇ����`������B�g��6�?����u�=�~��������ϟ�߳���o�=��������xo���g����v�m\�^&�5avmvM�K�-����+���*��sE.t�{qh�l�y��[���ߨ��|u�oKaH�b��$�(>�D�)Cb�)mdd��]��N�6Q��5?�������J����e
�!'F&.�#&�a�I���yG͡:U��m5M!��b6K�Y���S&��ЛgR۴�\�\�v�ٹ��"���� qIy����{�.�^w{��b��]F~QI4v�[ɛ��UB�,�D�D�95A��I:�n#l
���(%��0.�>��'J���)��K�t�%N��ݧJ��$��g\˿c����N��a��O���t�޶R�~b��jD+qmD��RWO��ڨ��{wB<�2���<*j��������KBJ�46_�x6���-G����rY�͜��a��Ϊ����]~1�D�y�94�2$�@�ěQ�"��f2����C����X�'e���ò H�u�%����"��h�M�p��
*ESm��/ �y]������� �\��h��Ā9˷�{x}T֢ӊ�������H����s�@x�M�5�:&��Q�^����a��{�zuv���_�g��mV'�aty+�:9���Ƅ%a�.�{���ůr�BO=��m%O��
��\�"��Y�B|�_u��ե9H�(cn&<��žK���������r���S{YB�^:�6Б�&d�����m��TqO˷�n����%"�� ��sx��}Y=Ф���	�S�%�r�B���"�֨$A�k_��7v,T��I��Y�H۸.ֆ�.��1�Q�\D�JR���|-�ͺqq���.�S��2��B	I
[���"���Z�;G�wxu�OfW�vd'�r�3�����p�	R��Z1�I�23��u����Vڮ�@uLv=>�"#����Z���Ap�MQͻ�{�������e{sw� �m��Â]xgy�-��Ԋ��C6 |�~�k`�~�2o=��^ĺ�&I.�0���Ω�g}�s��Q��~��=�_K����:Eu�S��{D�'�G������Rk����1v�ї�����P�]�n���	����҉��-�F��ǜ���̕��@��~����%�{s�� m�֫��L��:�T���F�*�x�䊨I a'�	.#���kƐO�FB�S+�-�Zn�I�0��g��`����h 	iMQ���A�\vV��ǣeLi��&F��w�lߓ��G'�02X6�6��׎�[4�D��X���5�Vtb{N��3Fi;���T(�]�'�oT�aȥר���W��m�$�����Gf���6���\�`��x��ˬ�^{�`�TN��&z��9W����/��4�o*���$=VVk#ɛ��t����i`^Hzt۳�YE�V<�0ݰ[m�b��l�HO7��<��Ӣ��sv,~�	Vώ����
>���>z^�;W�#hk�?n�L�d��W�^ƫ�%f�^֥�.���ѱ���͖F��i�Z�
NKS��w�O��w�7��$~%(�8)�gf=��9�H�8��Muݏn��cW������'vw��g�loE��b��~�,d���g����=���5� ��#Q n�m�T�����D�,�1 %1�*F�Zlm7X�0J�k����=szt�1
���U��1��y��a��T�*�E�đU6�}O�[�$Ą��Eۻ����-�����C0P��Xe;�3~���u�2���_�(��h�$��f�U��-Yk�>*w9h�lx�Y�	nU�R$�/$�.��͎b{��<T��� �����,̻�]�"d�ù�G��1�DVx�̜��>�7pp�����?�vx���w���?}���ϛ���wX�צ@��1(-n���Ef*܌su����G��Y�cω����2:k�Hŕ�E���N��d��{r��;�����ѫ���n�:��PR'1�w/�L���|;R�^������.,�%Nk���d��Ө�ɫ��E�MV�'�D�����zן]Ӽ�ʫl5�N���-dh��#�"0��?��;��R1��;^�z/�;�
ㆍta�� �H1����=R��lJ�����S�"��Eg ��%| ��T���&-��<kruL�AYlZ��B��H�������(����7���ֶ��
�����*��8	^9�GVЕ^�M5�V�i�Ԣ�5�Q���ƥ� ��α��yW��w�^�f7��-��j��U*���f����-��s�]�%���+s���H��4.�`�	��x�ȀK�Bv�߬d��`�s�I��YEJ9C���6��n����mJD���^9g��3:�*@G �;�s\�k��N4cn
({]���9Е(4(��u=aإ�N�'B�����ܶ��D_x�u���ڲI��ف�mR5!0Ѕ�Z�8��#�:�/�x�I�o��>������
<��z���uL�g"�|[}}B�Bn���9��oK�n��Z\[�xY���q�G���ꄿ:�m�DW�M�q?q�T�˨���ء��Uv �]N�zf�V��y�WX�>(#ŲX��^��Tݒh�Rg��(o2D5��ܭ%ߦb�)���ѭ�E��	�Ð���.��g��7�%Cƞ*����q�]��S
�p��k�phF����Y�k��N�Ɔ>=��%b������=|f����)V������J���%�B�gG�>�>��O5�1~KWd;պP�,�V��\Za�oBk����s����R:����NHھ^����Ԇ��Z�yNǼw`ȃ�4��=�ĘT�g",�׍��'y�6	��"���zG4��̝=�`�����Wd��ҳ̅���]�|<�.6=4���H	��b�	@�Y]ԩ�,گx;��1�O&�Cg��awGn]V�/{�蔼����<l�۷̓�nD��̈�����-G����b�`�<Iƈ�`��m�c��č�*����냍گ'j�7�!� �y��0�(ه�A}G�y��˩oU��
�5�)Me��C��p��9��rw�O�z�z�.!�����_<i<�;�7;��vs7r��V��=�t&�)V��!�zkk/�m$r2�FqNF�W�n;�y�f]m1:���)??sV}^>#��[�6��X���Xe�;��Ƶm�iB�Qƿe��Pf!��+�pӡ�؍(|��z�Q��.���S�X��FQH�@�5����/�Q�5T:��l�8}���ߴ% G��5�^0D��T�H��L�'n��Vfs;}�j˓}�	���S#ʦ���Z6l�{	T[�Y��I#OzC�b��=�M�����^�gK1߱�쪫h����W�^)��D�����!B�%�wnX��fM�-wIl
$�Fid���U���P n�P5�2oA�1B	�>Se�/�&��N;�/eG6ws��`f�n�+N��ăPj�uij��vۜ��;�=�=��6�$̜���o ��m-ޕWz����
g����̈̖R�*����u���kQ#v�����o�C��x�7��_GZY��k�D���XD��X��	5�ճnMSI�UE���Yf%u��޻.��M�R���������z��҅^f_wX}��S�� K���E�!MQ���-xǭ��r?�S�yZBY2���J25Zʉ���`�o���s�y��Gj2�Q�1�YA
�ڪ�^�	��ֈ&��fGl�mPQM91�����%*��遲�jy�'Ց�*��]`�4eS��؂��e�_�Ė�6�Sux��.�9�}4����ezL�.�0ҽ����J������[�%��i{T֖v�JGfU�à����b�C��:[Ha`�������T���W%��;���d�qa�8.�+p3�W�����i��o��rey!���l��r�֥�*�WG[�tz��iZB��'���h�ED�[z��1~��������+sU+�nܕ����W�iu�L���x�IĲQZz禾dri0�����ɪs*w�n�`�B�����W2[҇7�3�3|62��>����{U`O�-ѩj�{sO�/ɻ6�k���O��#��[����X���n�����C.�e���E�l��=�`i�̨Pikq�U��5����a���7;�{,M�D���^e3;�����8}{yB��C�I	d����n��CKQ�=
laF�m]W��C�[/s���%���gR�!B��pC���;bE�c8�$��y�!�;�}��d���i�)�#��n0X�Wv���mfn�,�8���os��"���n�ňytU'�)���uf!"�"b�{������rBQ��zA��v�K,>΀G�lh-GZ�nEp۴FX�/_Ley�m�׫s�=Y���N�Dxٱ����¯U�28��1G{.��Û5�lt������-��tKi�A���WW.���{�ߣ��#xAL����N����h���r�G��2���c6a83u���&s�eO��J	���}�
�YS$[�z�.R�v���sX�HX�ý�~XW�Z:{��r�M接8ή�-�#s����u�Wt*쇜1V��n�4���*H]��o��ѻ}�
���}l�|�5�|Z]�;�׻��!��R�j.�Γ�L�o&���"�k4��p/��7����k1Nt�4V�B��Y[��LU���2q�f[t�20���d�ɹ3��K0+9�Ӛ�^�+�J�umH{P���ۥ\z3�v~r�Wo=�I�Y<q�� *⥝.�¶���O�Ǽ���eYOAE�*��Z@�y��LF�Ӊ�c�nՈL̲��%B��k)ܵ���պl�쳮�5�a��7���F�V���T`�k$���M����̵�®J�����hJ�Z.nv�3.��UV;��u�6�JI$�HYI�$�nE�m���Wm��k6�m	�]'��6w�ا�)�m΃f�WcuWQu�McZ7��{�G���t�&:����	UEiU��Vs���>���n��'����V�wT�H>Qt�i�F{���Xz:�鈭�'s@��Ĉ��wv��7�3I�W<���ԍ�WC��̴�"�~��+���]|�=�l����ա���[ma;&����bb��.���O��N������
�7��q�=���!����KQ8�d�bm$���v{�D�X5<�b���;�
���W5��l�P���1�n������`tSʹ]�F�e�����nde�H}���Y��7y�#-z���,���Oɫ��au�g�l#l����珓w�ry�O3'Yu��S
P
H1���(�C�(&H+k36.�2Y2H��}�'��[l�%��bݿ;�u��I3�6w#�0ٝq��Y��m��Ynb�<ћfc5�5�s��J�ˉ���<�Y�M�32�����,���K���-yZ���m4f��Ea��f�c���Y�(�hb��5q�,��a������s�6�ԗ2�J�%��z���$�[�(��.5�b.m11���ɓi��k&������5�i���oX�,6�֌&�\:�v0Ԛ��5Ė"��I5�Զ����[%�K�]wKm�k��K�"��X�˳	I�1m��,5�m�Y��kf�3$��Mt�fŖ˚mRM.��kH�6b�$�-�&�)wdiI5��MLźae�Vej:�$��l�-b��������~~���yhͪ�i�����װ��40��헮N��m��ˏ9��G߭o%������%��X:ɔ�U�vKN�)X��H�^� �\B��[�������w�x�o,�F���]q��+L�3��C9���xn$gW-�Wy���d@���gH���#C���C�~����4C+�B<���)���:�����G���^��S������t������C�Og��=������:������z=��I��"V?�#O������~Ŀq X��|}{3���}��;G�u�N�g;ese�?����w���?�߷~^#���������5<B#����N<x��/���>'�?)��x���W���߈//�T�]�CǻĈG�|�#��j�>��E=������O�ݒY�����xl�I������\s�y��e���_+��{���3����7�B;�ah���s�7�x�9A|��3>���x����﯍���y�����}f�P+ш�F#�
�?�?���q�u{�;��o�x����=�^���(�l����e8] |3��>6������2����	��؅Z�!��d~�����K���7��|�N�臍x�/�|r���P������;Ǎ�O�?�)�����>��K~�x��,�O����>���Ў{��/y���4���&�2>Ư'�ٙ�^k�j��z��z���_���<OǍ���'��B�j���t�{���Ӿ=��w����������������g��d����^���NX���}�"xǏ�a����\_�?��pm��h�}����-"���(���#�jp
��q�4��S��w��%�R��O�}?��3�cMv�<�>�����;��:��G���/��������?^�|M�q�~=R��rw�6���������ȁ�6~|�:q$�[_�}d}�$m�c&g���(�#��(��Ty8B$z'��O�|��/��:2��������W�$_�i����uH��?��Ο���4�	���k�,C�{Ooy�z�����N��{���@�s����?6���3ޠ��<G�����~g��zh�F���wo��W��Rr��?�?{;����{�����`~�/�E��<��}|�ȧG�_��
�#���/T�|����>}�}�^�ZV!+���Q�D�����O����'G�-���|s�������������z�7�#�f�(���I���}��uC�g�?>!��b6��D�Ԭz>�N�x�L�<�l�����_����=%���� |{�F�B6@��+�X׏v�����~��������?��gg�nT��vCԮM������>���ޜ�A�KL)�����i�BBш�Y�0���~����*�����>!~N�$Ak޼W���������Ǿ��=��x��{���ϯ��ק��1t��D�C�=�}��:I�^�y�=߯{��=��w�+�*t{!�*���ާ����7�~o}?�;��=�9x{��M9-����wv�n]�}t�]1}	�u�r�	�Gl��L�����3�b�h8�i�hz!��������i�wot뛡r\�l�����U�O#t�$���pY�m�/,����u�,�w�G��=������'u��
�Ǉ�;��}r(}�:��y�>���Oh��D<L���{��q�?�~�x��̆J��s�?��}M�q��G�G�N;�_>��������u{�����jwF')�������~����_u�A%�S���O���׼N}������8�[o�$f;�瑌���(�����u���`���y�צa��@\
k�D�����tr)G[�)�r��0�>'��������_����́S����C�!��|�o|�>������ϰ�Og����W��^����J���S���?���~OY��{�߼1�e_�~�����`��9�`~��tW�'����i��B?4�W�}@�WG��43PA���u{ￖ������}��}?���~!�������x��|X_ T�1��{���k#���:�/�}�P��_>4����@���e$,��/��x�a���������~��g�N�J���t�C׺X{��z������{������]gO�'�C�'OЉ�s��7�;������P�������(�<�1�0��~�6��׸}�����1�%��o������������{��7��懏|JעF��'�L��%CB��a���S<d"}O?9�Ʉ��F6�H?'��"s����z��r�@���rp��p�����g�[[�����㿓����+���g�?����9?<~����@�~H�����bT�?�����_Ӎ�x����!��|���|{!^﫥C׏�ǼK�w�_����"y��g�QK��ᴇ�H}�Wm���~�!�p/ȿ�f�f���Y���T�?ݓ%��O����~=䀵���?n���������ѺtC=��C��������׌��+��EO�y�T�?���g������ﻪo��<�x�C:�y{�x׸S���Ε�|�xk�}�f��ߠ����J��>Ô������j�O����XϷ���_P��׌�X���Ŭ���=�{z'z�bx���y�x�UOɑL�c���ힿ?ӷ�y{�������'z�𠿀��J#����Z��s�ʼ��~�q�8_���]2�ףo���x�~�����ﷳ�߄"<~��������;y;��vE��䂆ӏ��{�O�%������;���{8����'x�:'�����y�f����;��#����dh�H"zX*b��i�Y�v�;�wz���a�l���Srr�80��xU��Wnv�F�������mwU�@�Ov�
�r�K���j��L�
��53 �Q��b����{�w\��G>Q�p��}q�ϖ������}�u�����of���w|��^��^�x�����B'uxzt��c� x����"�������oӼG��w��/�3⻼���@s���(� ��}�[y�Ծ�3���/��<x�b��x���x���<C��'���|��O���;���׌Ǒ=������'�w��*}M���?�?�Z�@�k�?O?ۋ�����+^���>��͞�����?_=����R ����_�37�]�ߑ�����~���j��0瞧_��:�W���y�n�C��T���������i�3����/��<rp���$��欁�� Q�;���m~�/��Dpnj��(�d3���7s)ω5�j�o}z|q�P���2�b���3�|3;�޹��A�Q�I�2h��J�Q%�Mr@E��M`�'�����u�3�d�N�eM{e ��x�������*��j!��oL�B
��=(��� v�L﹡M_�,�sf`�O7���^p��#�<���Ǭ( Q�1�BH�dJ8[��x$}��ޗ���_��fU���$�U6�� )�ǆ�E���d+v��ܛ{��6�������!ֳ���Gƥ{,^�4�IW:�Q}1�����S�)]˂F�������|7��L��+��zeD���W
�գ�o��+`r����{��H�bA��`G-^�m]�A�~��=w+�h�3�	o�������wݡ�����U=:���s�էX��>Ȅs]Ot�oh51�r}(uK���Bt�`CI���~���GH�,�"��%�ݞ��%��<Jz߱�K*��u��W��V����⒕�w�Z��S��4f��¯�5�k�q���僣aOW3�NP:�-������6M�p(d�gL�{}��G�pM^8J�'��u��{�U9������$+�������Mk�=)�T��[����;xj�B�X�F��ۆ��f�2U$HQP�=נ�w;��u�-��!$l�t���PL<f!tn�r��ݪ4`�bd0�aݵ�ƍl��k�VY�Śa�f�6������oDЖ�ԗ7�e�Ѻ�MF�4%��M���8�3v�ؕ�)�{��d���o����������k��J�T-�8ޭ�ߚ�)`,ڃ��a�t�	��Bp��,��^'��,x���ND��������.�����~i�N#\��R+�4q�ةY�!�˿'��I���z�3�VL�ȫ�����w4�^S���gu�r�q	��yM��{�y�Tks��Z�)Y,Z;�J.	��c5�MИu�狔3��������і*�Ϻ툖]Y�n�-ٲ;.ĸٝ��ů�N�ӥn�q�V���H!{ΛG�����R}��X������I�e��G��]73W[���Ư��CИf!�d{(�$����"3]�fMo�lypq���7"����χ�*#�nt�F��iO�B<�9�_ 7I:e�^���s��̪��uu�%��X|�h��hFKV�#]�,&���˅�z�����+
�^����WA
c^�e��9��?�׻rO��o��jg��6�����`E�C��&x���6������FӴO0�g�7��]�.�϶<�M>�ݞ���#���N�{�1!��}��}�U��ˢ�5�O Ǯ��Y���M��ķ���(jR�N��Y�r��^K���:���TH���n!��Ѥ+bUyl��R��/a���Z�H���T�.�b]{s�׎��an
9��誊���̌�כ2�mC͸q_�E�d��,��A�b��
�[_]�5}+uE����f>�æ�hq��	��,������aV�n���TpѶ�9�_2�uѭR:
�_0��=��ceR��o;V��\Q}��h��L����k//
U,s��3���%�*��e ���yۢ��f��(k�]$뱱�Gӗ1｣%ej��ٳe�^����KC���\r���v V�̧Bơ�n�h�^p�e�|���0���2ꊃ=�eA����\Qa&�i�5k�i4�l��y�y_+�ɴ4z�rJ�V�5�8���і�m�jߙ`�7gQ��T��v2W��ṋ�T}u%�o�}Z��Vli(�F�ѭS�*m$�߲�#Ҩ���φ�؆�~��R��gII�����fٷ]A�GH�s�Bnv嗺��I�hQ>�Hw�*�v�S7���o�<�d_%�*V�ǣI��V�h���V�2��i�oç���zn�N�>�^[��jNҏ@o���L���350ۅj1Ɨ�:MY�=8MY��c(�� x6���`Ƽ��\w}e�G~TSӟ�ՠo>�:���z}^߇і�,����6U�
Fc�s۪���~�F�'$a�'��F�i�˿b]\J��ʟR��P�qOx��Шn�)��u��Mes�{)�]q6����kړ/�$w�yY�m����0��!Prc�5'���`�����$}V��n��:{��T&\��v2(���n�oˋ,�{�Ei�RrX��X'T��"Ǎ��{������&�I���u1��s$ɞ�30�kd��h���.�����D6�wƨQG��zT��x���x'���)Kԛ_x!w�'n��)SA4��6���!m !,���`Ж��k�@�;`��3	��Ɨ�:��	`"$�A�i%�6��������������ca~�OSW�nd?n�}"J]�ǵ,�兀v�E�ĵ�j��vǻ�����>��Y��H�UL�Z����8wb[�5��w%��N��Je�V�i�j�xgF2�1]W��@�v�!�铪�u�����V��}C�&�
�0�M9+� �����-�\�d�z�%ٳ���3믩3��R��&5'��&#�{O�1�+��p�q�/;6���"`�W;�'A1,��K��c]S�b;�� ���%��3A���zi�`����7ק�I�ɪ�7�)O2�{.N׌��b[��	�F��:����!���y3�S�ɝ�
��|c�:e�WG�ɽ�����Hؾ�y� ĝ]#9ُE`�a���>��˵����N7�1�C�Y�;l�Ew%��hy��.��(��V-�=������M�a��j~���AY�qXk��v�~��[�~a��5,}S���fސ�O%������t���C�����r�����+p��т���5^�����x�ǰt&� e�z�l�1�=�����U]%��}�3��~�^����_�Cf�]QK6�J?�u���:]�|V��%h ��WF�Tea�
Ǵ�e�=������
Y�l�q9d��H�����,�$#e�=%��_J�u9�l��?4ZZ�.��wR?UtV!{�R6КK���$X7͖<C;<�$x����&O?��G�:����(�0��q��L/۞y�a�ZŁ��|���Y�ἠ���/m�YX(�S"�*�#���ʏ]���xo�.ɑmT+���?'��_�k���=B=�g������(�<M�ۅVt���2��dߟ��,X����}G�q��8O�򕷜g\@��In ���]qm�?׋-_)8n*ɞ��N�*�cy���|d{�Cǈ"��Sr�@��W' �9���8y�*u�ܚ��� W�-c��:�B���Iq~.g)ϫ�vϪ=x|r	\��q�W�;�\���Tk��x�ं؅�^��<����ı�{!�������|aQ�o��1��-�S���/z>8��;��W�>�&���D|;j�yt��p9*ڑ芮j�y�8��yF�k󩤑���5�r��g�+��7NT(2�<M��\�/���u썅
��sW4#c@7¦o&Փ�1e����B1a�P=X-�j�<[��Lf�)Hu�}��m�����Y�ѥ��`���_-��T��S�\~^!���U���O����$oMb�F8AA:� #��B>���8�\�=ʍ�Y�}�n��e߆���[�v���%צεe���6�31l�����2����c"W5�l����rߦ3I�:��L�x��R 鶍�8�B���پ�UNz�f#"�4�p�7uia�x��&Ѿ����]�Pʯ]�)���騙�c�`cR���OU�`߽�Y�SZ�w^�?n�$����µH�"(Yԗ���7W,�a�Y6+)�%�vL���o,�׬�˥
��C^���8��voO]�I{+sy�ˊ�)sH����͊�O̕@+[NP����R�D�.�U�6!wt�a�vS�NF6k�ETb'���ɞ%c'b:��fO�A��s�'j+�c:p�IX�~;{�Upn	&�:����RI���������N�'Moc�#nV�d	�˓3m*�~[����H���=}�HoՑa��wyah�f]풤�@e�O&[ξ��=s�֭M��ڑ#BF�A%��f�#A�L��bv�w3����8�QU���#�Jj�p�[lYt���y)e�5�%��1��b��$����%�6ę��Z�-�jY�A�KΛ�h�,�d�d��:i3,�u�[�'�a�"3�)��8��O������}۸��L��J�eB6=�&��IkFO{<Ssѯ��1��H<�#	[}�#����
 )Ҍ{��;�6+���� �V1�o�J;Z�5f�n���2� lV�SP�	�x�M8*j��{���z�'w�h�@����'9���ܙ�G�*�_L5��)�#o�N�B�"���H�jv7ܠ���5t��j.�&S7�"v&��GV�U���8gwB4��ސ�R��)#BFan(e��k�����)5��r���� ����P��2��(��pL{uW���,�e-�����R9��P����{��A+��M D�&��%b�-1�axT�2��b���_�ë#�@�X�Pf�h�ݰ��W���#�<����+����:<IW3L���[�lpg+�l��>�,Z�1�]^����N&O��ޟ,��ʁ4��h%�{�>��	*H��Wb2g��Ҡ��F��)jT�ez^a��{)ul#��>(������M��� �����{�Ƨ�/1�.Y;�~1O�z*:�{Y�K0&�Yx�U��(:��I��2ި�A�P�T��B�9�<�4��s�y����*�VSJ}����'�^�O,jdtDDH�F�'�o'�d��hB���i�yޯ�/M����B��B����EnĲ�k�;�u�"�n�2ҟNӽ��`�(�bh ���O#�u��.�>�����˓��N �q!pz��a����cl?�bC���Ũ�k���f#ݠ�In��x�9�U!/�ՎŽ/�AH��@��_�]�e<�#�av4/�n�ؚ���mw�ʕ��O{Fİ���|F�|��gwg
��K�m�g_z�^^��yk;�j�IǏ|NѐI/q����@��ܿ|�o����5q�X%��{oۂ�ʣ�ΟJߏ��t��ղ�Vm봂���cwu������; �1q������ą.+=~��[e��S�Y6� �}�c���5倥aժ�#I�X��eVa=���L��f�<�@�]�ϱ�
٘�5W��j7ބ�渊���r��t+�R �,��&��[y1�Zi�^f��L:	j��R^���&�f��fP�Ma�چO J7G��~m>q��ڭ�*b��$
�V���d��͜�Z"��L�˼<����]������✰1�
	���<���鹣hF㤝P26�7rE����J�ϧ�`��<�y�mⱶ=�(�ƹ�tf��<k��{{hl�u���l���	?yo�@�����B�	�G�vh�n����;�T���f�u����&�~��T�Q�̙(y�#����p�ݙ��r䶮��SWb�uaҠ��yo]����6����~���g��Z��M�>�Jh�x�Aӭ�vԫ�(F���GI}���#�"Q�{Bܬt	�F'F�LwD�b���Vg��$69P��]�\o��`�(S���l������0o���N��P�K��F1#�١��0��gӜ;�y�ˆ�23Z��22Y.0�º��$���E��f������p�`����N�����4D(�r���t�y����SW����!�Xj5J���/���.�3���$���Nɉ�v��٘f��q�tY��rk��oIR���亮��xE��Ӑ<�v�{9��L�R��N�Xz�/�N}�s�0�e����MȈ�WukT&V�����v�|/�=�p��E˯�tF�:� '�o�I��;ҏ�e!2�{k�����S6֙n�x�d\�>َû�7٘����lQ��(��!���߶o&���QWOP���@W�&ٸ�RiK�Ǭ}P�g�f|�=*�\=����v��h���%��Ax��m���(��V��5'y�z.�_�����j��:� -����h���:qN��<�y;N��>�^�3�՗�$+}��0C�����tID�V�A��/3��J�����I��h��Sf�Z*#f63GLy#w9O���A�-I��ޏ�S�x����>�=���e(�.�y�E�o��aV�(b,6.6t�os/�+�D��*2f%,��U���=�3���<�>�mh��--f��[�-�H�r]�6׬��k#��TC��3��w�l��D����$#ѝ!	ܺ�s+�	l�����«���ᐗ���Z�v�~^}nD���07��U��j+T}� g6a��c;�8wHg���WZ`6\����FZ��B>�%(=#�UV�]}��.;��@��@]�/cӁZ髻�dVr�F>�$ƹ�Í�W�c�*�*A:�����6���(H+o�g�7�J�j-[��Lf�8ע�+��{�/5#�<�,Nд|�� ���/ J�u<���a@�*�uN�C���y^�u5�L{����^Y�3��%Vq�*X�s�R_�*�%
�B	V͑Q9�o���t$2����^��񒾘��)0q�o�wuњNzF�9K�sCx�h�L҆��������2��9
���=+��V��C:95���Q�q�4�
a����������g
�K2;�64�q�x~��n���a���8�=֔��s�p�t�V=�%�G�>PY�2w"y�Q�ts{{�Q��b��Õ�%w2�SX��H��C��3p��r]Dv�q�z*«(u�7*j�!O%d�f�Y��..�7�Y�V�T���X%���g�c�I�Z�w�:���v��&9��9�;��-��-�e��:�;����R� ��<�����sYy��V��[X��)�9"�+�f��f��M��ݼ�0��v^�=3�;��\(rz;׶��D������eNt&s��}%�sf'2�t�Z����]wn�Б�Fޙ7Z�5��rb�<#�s�mb�=��[���t�����pڻ�KE�;�#�X"\�9�L�+m�9�FO��N��;c����>�&�J��2��4t��=�s�k�T�o�P����9��RN��}ݻM�"�y/*q�X%���v㵎�>�oL����q�\	��#=QQ�{�e[v^$�oe�:���wL��l��̘�!|&�ʰ�x�3�t�,�!��,Pͭ�L�=�9݇[��s�T���E˾[��ج2\"�|�u������w��%&t��6N����gt����c����u�&��&I�'��aY��k�o�9�ӛo�I��H؇������y7���}.��TTq�ؕ���u�m��{`Mo�o�&���!����l>ԡ�9�C�Ѡ�EӔ.�F�Px�9�mj}M�����g."�x����^�%�p���պ��˭%���̈:�9�=;s+�{��]�38�N�c�7���^�Qzw����5E�ٹ��=d����]�wr
,�-C���*�Pl��=��^==�.�Q웰�}�wmiz^dpL��IeKWX:נ������ջ FPu����YZf>��>Bb�Z�`��)�Ф�K��gN5aJ
�9��qX�rQC�W>݉�[\���i���=nuZWvn��l���5{��ۈu*:f4�WA3߿~�����I�Y��ٽ��igޭ�je35���j�wt�:�!sgf�u��M/��y�t`��U��0�]O�R?��i����T�'���>d:}7H�kۓ��L�����Q=5o���O�&$���]u�\��j���s��[�k���W��Se��"�.�?d��|&����dc懫�v0�(@��l��MO��2��ⲩ�
c��y�t^ߠ�~j&ԶQ�����1'��e,�he7L cv0�]V�����Ӗ�.�[��A�1,q��OS^F�2���kе��fS#Hы���K����"������Տ-���q��Z��3�dA���l�uvKq\�/�2"k���XJ-]F���F�*�=�[|���dxF#��Ch�1`�f3�77��=UҮ*��1�Tm����5!eC!��}M����ւ�H�J���2�n5�e� �\�� ���ګQɗ0���'T���w�[�c��4�UP;�Y�`�)u�����&,D3�v��ιF_�Huc��l�vU�5�j:��ޘ��O>��s�hDz0�
s��[�Q�
+�M�p�n �|��D��2��I��Ė�JNY*�)~����7�y��"Q{w�s�
4A���E�]��Y������Y̺���D��t%�vJ���ˍ��:>G��l��ݮY𛗳�H�F�6�Fz;B�T�=)콭o�e僾�(��@��>�G��\�|��8heu_��$cqGknUV��T:��;2NG��)�~̬>�d%����r���ɣB�Bu;�(�[v�w�\�q�:���^>�82L8̎~�;c��Tv#
̈́�����j��=�%{�7P^��({��Qgb����GRrO|��7���5X�ٰ&$�e-q���ƚ�lm̑QRS4�iKm�^֑1�y3�����d��&������΁��b�
U�#��f�����'��w��r�=䛝�?�?�V�|O�c�uS�o�c�5��^|���;^M@�$g+��Xms��k�N�����۷G�ΤL���� �jf��w'��k�m��������`�����[$	5�Dy���M]����Ȳ)���y^q��o��yo]:8ob�g�뽴񷺙��˩py_S�]E���v3�ǹ��{��ʏL|pΓ$�Uܿ�I�e�Pi��B�d2V��#W(���_��t��`R��I�C��ӓF����e���!���>�ۗV2[Z����n��U=�5�:ϕ�v�+L�Mn*��l(XvI�R�i��EWmJ�7Z^^�b��
�ݗS�G���}���k����3��^��;S�T�Z�&sḏ�N&=�R�� �5���Wjm}I>������./V�	�>Jlg4⤑ъ#���^L�c͓e���
ƃ��g��J�!Ǒ�_�2���C�q����2G��+E�n+�ų�F�i�w���Uٹ�bҞtϐ�zjN+싏�>S�k�c��Q?�}Tu��w�F�`'�x�� N��C��g;3����pM��3<n�D��A���}N"��ecVuO~*f�: �i��"rs02u
�����;N�]|W�����X��+�\	��c�b9�l�w;5�T�>��õ\Q�����nșj�7� V]Q�D����y,=��~��Ys\�Y�U����)�6��l�;+*@��Oc.�F�r&bWuem�gJ�g����[�-�R&�tŢ>}ց=K:�f�)�1�FYo[��ʽ�.����;����ۜ��>Q�s L��yC�伄�KӥK�G!�v�@����j�vK�hw�ߙm'	���^�)E	���=]&":�;��~�g�GT��n�<ҷH�����W��i��}TL��1�z��f��2�����-t��+�3��� �u��T}O�}>����T�W\�����iB�ǑI�I~ޫ:l7Won���H�Z!L���i���\~(�7�O�=m�[�E���^����w5��Ǐ�U�H�yt��="����0I&Ǣq+m+�V�-��"�����D��Τ�.@��Z�3���m�L
ޣ�4���ҢcP~ ��j��@���`�I4�!��M���B������D��z��s:ɚ�ӹ8꫸Έ�X*�s����-�]+�l�~؂^�U"#��X�S�Rr̫��6�M��	!�h�r��n|�M��MN(/}�����o(�������H_7��u�I�G��>8�����'�:�fZ�h뛧ދ,��u�S�N;��k�̘0��G}����ʾwF)�L���7�^�2����O�7a��ɓ[N�P$]mOS/z�;l�B�3�ٕ's�x쬺��Z�Y�:�p�$�2\�9SUƶs�g8����J��J'B�T]��q9S;/��<��i�{������W7���A�@q ��D�9-���ǹ/����W�KNˆdگ}W!�q��4��%�%׫(W��S��vcB����@���^�˧�g����̗��w+$bB�q�-�����T�@��X��Y��U�]�u��]j�b���\XypWW�$���c�(Udͼ�g�5��;��a���d��oT�����/�z�Y��+�_�zq��b2�yu�c����i|C�^^���&&����$逩��}Vg�֦?�>�`�|�puFea<R(p�ca�y�.(��5%:��^�����,���m��G%-^ïᔼ�%<�鯛��ީ�M+�O!'���{籕M�"�"�Ut��˫kc&n�s��3�G5�9#��=w�J��w{�[�h0~V}'�2`�T�{A�*�|�$��̷x�V-Ϩ�����"S�q}��CcH��f{F|�z�=wFZ٪����ձ���oӄ�e�i��L�ϰg;����%�[)X��[��)�1���Ԑ��9v�E��O"V�s��ޣJO���n�P7�7�4 �g�X��^�<����C���.�>���j����Bn��8إ7;����/�>I# �~����W@��dꅮ��A]g����3��3��Gݥ����AO����j�r~d��܂.���K���C�B+!y�pt����䢓ˢ�j�����6(=�u}��Lͻ�EOW}ˠ��� *W���h|f�=�z�A�Cȡ�*J� ���f�"5>d:�[�j+�X®R.������zD�I��9�Vm�/`�]a';P�DuT����$g:���Z��$�(����������Isюl ���S�U՛��y͛k�;��?p�6
�S�\j��rж��9 аCX�<�"��[W-.�7��MZ�-��o{J�u�H�|G���&3|�P�_Z�suW�?Y�=��T�+�^ynk<BȌ�V�k0���9�:�=ؗ ���̺��u�|���f\�ʉ±ɬ{uZI����ߑ�}Jz�=��z{F�(��E�r��F���״<(������m�!����޸��PT�F��<�f��]0!�p�5nh/^j�A�ѮK��3��9U틿oBUdo�G��i�DDk��T��vT��c���Hu��z~ytb�+}��j��@���b{�6,�G%%��בֿ��c�x��N�P�LԽE���N��^�u�{�z�u��t.+��׹�s=�\�b0o��ʗw�x#K��Zv���!X۩��E80&�E����%|������+��A�$jg���_fZ2���+}�&?T����[�0���1�8��e�K�������ǻw�f߻��!
��oK��ưeo��ҸZ2a��φ���J\����������>��6z��$�Ѽ��q}^5�(�FF䔚%V����o�ܞ�O_y�U�U=,���'� �j��;��Q�7'ս���I BZ�\^ō��W�p�,���(ƥ+ݫ�o%ɦ�G�zu�C#Vzuq>�*���G)�%�ϯ��۱g�#� ��Z��>��(8pT�Úe�&��\��]�Z���pcM�	�׶$�"��`����_�قՙ-џJe��}�qidw�R
|oM\��N��:�����/L7qL�¡���35�����;;c�*�d�B�Y�������g.2a�/�9R�f�swH�b.��Z}~-���W5�*��]hؗiZ��7b�k)-&�X�b:�\$�1S7k2Ζ�U��%�U�c:ݣ%���fy6.ي�ql,�Rer��%��k��v��N�J=�H������_�Q�gi&�w�4M;oj���e���;1`�j:L����`�^�����a\+���l8�'PsnV9�}./�Wzq�Z������5���"m�^�-���~�T^���ꜙ9>iI
6Ǉ���������W��>�g�Hz����/Ν���60n��zo�}[\�3Gj|�ֱb��TSA����.�C�V�{*Ņea	��Q*A��q�~��ح2-��{����x��-�y9C�>;�w>dv�<&�9BDlG��6ӧ[#��������6[ѡϾ�۟=�#��j���&0�'Y���r'��p���u�	J"���l�[�s�Y�����(Z���@�LE�����u��%�10�^žv,:�*�o}�b�m��+E���9��e'��E��kw��+���K��W���u+�{� a�r���p�5[*��d��I�|�b9��$��R��;k���z�� �Uڐ<�G�#XG�|>�9�ւ���C��sԲ��쏭�k㬩Q͵;b/E�½>Uw��Ck�rm�{�^�[y���w )��z%#��%e���t�K��Hs��qu��}49�C�I;�>1�@�S�G{i^�'�m�1R� ��a�Х�(��V���{�5������٥�h���gx��=r��e)�B}t�x�.�v�upr��%!��/^�R�"�egl̒vv�1����k0�k|�+�����/���hui1�u��fA���N:=qJ�y�$/D��s[[�����O+j�(ȳ�!�����~�g�L�5\�7X��
�Tf�S��\h6��}#�o�@���f<6Ҳ�!q��jKJ�^$�ZÝ&��z�'x�U���������k�~��H�ʯTF��{?kU��-r���O�Myb�D#P�V �q7��1�WQ�И��X¸R�\-���2</-c�O����e��@��t��r=�}*T�O����z��j�h"亚�b~?���W��c�oH*�Ы3�d@���g�33C=�<T�&��s?o�^x�����He#�Qݺ7�����}>6&{�;�V��d*5�"E-��z�z�i�|����a��g!=>�X��9Ы.:��/>�D�g9�T$�q�*�Gh��k��o)4f{�>{�7�+�����g��MfV���C8]y�m:���F��䨋��<�}U��5���lo��Y���~�7���0��O���'����C�jv�+{ѣ��M�b���JW���;�����wև:m8�p��u�ʗ�d^mb���9$Æ7H�mt�Қ���onI�TYxA]�)��F|t����8(N���f�{n�RC���y�_��1��<w�^�}�	O��=�5��R���ִ��[u^�˱�����{_��q"�M�ى�Oq���q� �?@��]���Ƽ[䱵#d8�@��K}4�d���:<�Z����]Z8�.ݦ��;k�3'�e�f^�)6eg%�̭�b�r ��g,�RCq�,���귶s��R׆�ޥ���fd�?�)O�]z�D�)����}=�z�g-�E
����$gj���
a!q�,��D+��+t��m'�+"-E8�<�w�٩���,�<�RN�Q�!���Oj}�c��i��s3{�[Q'��Uz��ƾ������yNY���u�]ނ�G���Y���,��H��9�G�`�d�2Θ�:v��5y1|�ʔ{��~}~��`���s���Z�g��C��4��uq�#U$	�U�q1iJoR���]�s���0�٪�h��;�g������B���ow��T�Y�^
@Z�U(�n�<��aK���
���塚)}�J����B6��~0��HdVÑl���u�����"��L�)~=R���N��Y�%F��x��?Rz'��\#��[�Υ=����9��T:n����K ��-�;��!�`�zV&������5�\��|�栛��\���HgΕa�0��~z����U��K��3�j�imq��k�JD��`jz�wj����_���g����фK��ݨ�����c�wfc#z��7U���P
�M�A�Y�����bR�+Um'{��I��~��ip�g�b<�ХNq>�����Ǆ��:�[�g#�ɈW0p����E��U���}���^�?-v�8�c��W���{��{B�8(�[���:wMWv�*�����n��4���r�cw"F��|�*�������%"����y݆J����-�����]uV��q}P:�+�{j�os`��cR܀%K�߮I�P�H�]�B�o �_�x�x�f�/Cf=u���)<��������,L�W��&f�6ɹ���g���}̩�|�[f��̡�����n��"���X�4�h!��Eؕ��W6괡�'w��>��#�yN*J/uA^
m?_O��äk�nUj$�������%���oBq������:#�T3}���r�r�{m�16>99c��奟��7��`��}}�Q��n�W�խ�	�cG��<�ǞW���=67���p�������`��6r�.��L��\�;����,�f�7�.uN
�O���@��9l4D���lȜ�)S|�Q�Z�;���{7Na�w62���ު� �%ND��v���V�?��;�p��Ƈu>�Y]y����@�{U�t/f��aٙ���؞KJ3Soɀ�-����d6M��b@�3=β�t���)�.� �^���3�Yo|��:�,�C��ف�AV$%I���������q�vx߫1e̬�r�ѻ=s/��YiR�u��Y��/���Ό��z�kd$�5�4�Q��>���=j�#DN�/�s|X�׈x��"nV.F�tDs�}$���Ā�=Nc�=�⨁�a����w�U{A�.�϶͝�ĺ�x4��
�
8�WV>�dٕ�dea�����oj)h9١���#J���=��75��5Wje˒@�B@�<y�g+Dif��#]X�f�p���,5���Gu��JY��F?��Q4AL���J����̒�jm��%��L�G#̙��M�i6)-���m��Z�2bj�˱e��3�ؚ�2�d,�&.�&b�`�"f/�㯶�4�r�ɼ��{�}彃WUM�D+��s����AQ�㲉�~XQE�7�>=Ա�a�VN�/D"���]Xű�m>��_Z#�����&���x�[ץm3>��-�t�+�D�:�������o�;o�m37�#�;Mx��,�����p'��$��L�nfڼ1�늨T���Y�	xR�7��;o�F�O����e��L�,n�;���GdRk(nQ���b���E2SPBr
�;���kϝa��>�4I�6�����İI�X ��PDe�-�X�v���w_Mx�e�6��W�3��4���Q�0��mژ�s��^ͨ�`��Ւ�ψYg�g\~�IK@'hNf��%tz�$��f�^�'��#cy�hg�O�Y���yBDjN'�ϲ���Ғl�_H�����YU��ۦd5���������"��>�ɳ�F��g�����%l��U���t�3!�}�+�z%�M���DSr1�T�4������`����)rzc��]z��P����K*�_ys��a������1��͉|1)h!lmj�o/�2t���Ȋ�f��C��r��&He���<���զr��,󞪈S~Ι��K�\������%��b����z��?>����w7��u�ҦI>,���]�BH��#�U�}��;_U�^ߔ���5!��{c|zC<k_���7m�T�Vpv*+�Gk0N3SuĪ����l+���S��։���Y�9�ޮ�y4�䖶��nU�t���q[�|�^�6��2���3G!��[~^om�q#��{~�X�&��-�ρxu���۔ҟ�A��=[�n�S���x-�3��u�t"8�'���ꔶ�ON�0�ޜZ�p9�+�34+-��xӘ��BT�1�m�$n�+zh�y��n_�N�B�i��IW���,�K�v�T��sB�q�ʗ���]�.�4N^3���7̝�zQ��;HL0V�X)!$�}���s۹!��G��u8���-�k-n��ĉ)Uq�b����ers�SŴ$�H��Pv�y)�妳d�6VoWm�6t�"v�{�l�S1�CV�7�T��,��`��:z\�m7��
C&_q|��2L8��>m����ܪ���ѷ�6rf�޻�w63���8�M����E�ճ���F_}�6e���k!>�A�N�wF�s�k��X�K����L��:�X��E��Kk�������9�7�:��6���+e˘4gRkG>���j�a�Y�b6�m��2�p�c�,h�)�R�i����1��9���(ч��sM�fv^՘��gj�&*V�����9v*�ݕ�W5����s�����[��s7���]�
omL��aRO.,60�L�^7�tc��0\)�Y�^��0܎�L//��,�黚�[0�ᦵF�h�ÒQ�7�3۹۹������I$�[5�m�i&�ݶ�ݭ��md�h[q��RH�mȣJ8��c9.fn�oC�U��%�o::ʼ�{�g纡��'����o1#:���nf^��Y�N𗧕r7������j����L�7+��xj�Y�CӒ�r�ݵ&�m�{��0M��P^�E����WaB5��>kM���^��V�����3QZ��7ٗ�`��M�˾�&�]F*9l�y�]Ά���{�ui.Q�P��B�sM�f�T]�eu����L�5 =�9�����g:�*�6� V4
����]v��lk��S��Sܴ3,7�uӲ����x����h�}?u��Yyf`tu*O��m�5�h������	�jW��L�	j�=����>>O-{�K�.u���B[fB�#�'J�%U�H��:o^�e�H���Ҳ�H���i�.��V��bRko�T�w��O�.�B���嚷w�Zy[�n��a�&��Ƕ�a!7aU��2j�v�3��b�t�[�\�R��	tt�e��9n�zYh���@��qY�W4���HmR6�����l,�W�.#�iF:0_6R���Iಚ�����<��Jo/k
R�Y��֣�j��/e�#�k+M(�Y�KfqZ��}���Śl/f1�2�k�e�&�3&�e�W�t��e[�|����І��7X���j��mְ��#,b��c	��i�R2��h���a4W����[%�4)�ڔ�̺�e��a�k�3�ǌ�fT���%,�$��W[�&#����2f[�FH%Ē��$�q",^��dٙ��	�ַ�T]�'��ւ�����fv8i�K2��v2���~&�P��u�0h�mkF�JQn��/E0;�-38���m��_��?~����{۫H�}�Ʊ	y�������.���0:Ἣ�}�$'�s���g��>��p�(9��F�I�j>��6{�	~����N~hk��ݡ8�h�Ō���3��O�x3���Pnh"cf$�PQQ��_dT]v�]u)����U��PnL��>EmD�K�y[{:�T��[f�er8'sH/�Qں��J�s5
���a��Ơhtfx+3uZ���F��;A(��3:m�^����s��NSʼ*�S=��
�n���֝ύ��0)��v��u/'�ǆp��E�V$Q���^M��J��{��`�����{�J����9��򄽅���:	�I-R>�|7'��mU�At+о���m��ӊ��.�h⓾�kc�Vw֚M8�}1��F�>*�^�\�LPU�����gQ{�G����o^L�4]�w=�'OMY������{�}�m8�#_��,�P�&��UvZ�Y��l7�:��L�����:��_�*�d�K{Ŷ�xt�.�����'ԉ投I�e>F]х��0"�N5C;�>�kx��v������c��ձ�5B����ݠd�Ꙁ�ea�Z�ñi�7ofe�x�l�n�+*3蓩��������^RK[���3~�6�����eP�L`�a�p�ġ��($�Z؎���U�=+
��J�M�$Lo)��t��^��a;����C�O"b7����͸���}ږ��#�N�쳧��~��:4z��.-��s�ا}:sp"�N��sVy� �7�=�X���n�:�CB�^s\[�����j��{zu������)��=���Q
�D���Eպ$��a�[}�1g	Lx�BBǊi^���+���*]KȽX^bU�?�X2��z_�)'d���O���g0�k&Lȣ��<w�f%<%S���I��xV��%[���G`���[ފ�t{��`Σ�F��2)U��nQ�褀�*�  `H���m�#���~+�_m㒶"�H���\��a���nŃ}\G/F�{)Or��CoJ�<��� z�q���&u�j}P|����oɾ٫�ƻ�"�/Odn��W+~sB���ͩʨtU��U�z�|ӻAϟ-Rv"�eP�3�-��Bt�Z��~[��G���-x~Q�.�=��.�b_t
���m4���&��Ƿ�]^����_�N��u>̼،��x�M�,�br�:J��Pg��vx#���a�28��ga�׉u�[�����/z�9=c������{|���W�Y.�6wc]���>_��R��6VDX�`�_{6_K�YL{�{�$��J_?�m��Ay��a?dz}�|��vW,�I�8���e����P��zt�x�ŝ6�i���\v��\G�=���1bYP�P�������v���n(��\�5�=*�n�/OS5�j6�s.z��������
9�9���ҵ��/�h��.p����#!�4���?eY� !W_�X�ibߑ���cx�t�ڒb���oX�5	�'�j}ڕ�ז�L7O�WL��'&ˉW&�x�w5���ZU��%Q�#�rE;�Uei�R�{�O����L�L���욂إ�t�$�Y5҇�8�1W^S ֥�m`�'u:ɻ2Wc��x����vEE&iuĎ���J�'o�ｂ�Ubx�>��<�v��~+�Ͷd��o���;=O��.�呑Y;�.�՟[�8��?.i��%}YWi,*}�p-mvϮ�J%T[�S���1�=y���{���Ci��6M�L�Y��~�Ɛ�2kc�n����=0��?�\�ݟ2B>��]��]V��[�+����i�P��[.{#Ty1Z�;���2�.T�O�� ^L�G�'���xg�7�b��|�7�7H"-6�P��M��E�j#��O��
��ӳ5)w������>�×5��It���'�bv��s3�kuT��:0���$�ʳm�.����>���[sgܱ��K�8���j�H{Y74X��#��E},	Q���m���Q�ܟ�3xC���Ԁ����.����*`i����
Յ�����>%��;FL`y���'��˵o:;h�<���W���`_�|�ۘ����^�.��ҡAlpv�.s�ݚY�W�ve^79�έۯK0Ӌ/~/�P��Q��'ѹE��e(4hWe��t��&MD�r�!���������Y*��?oׄ�@h�R�̄X��;���#��g쎝���g
�Χ�-�)3%&QM�d��Ѓu�թ�HwWPZ����ܽ���\�1ą��{y�l�jM�rr�3*�X�C��:�4n�_���[��f�7��*a�>j4�#�[4�Qk.�R����%sJ�ڰ�j�HX�n��K��1vnm��չ��M�J��( ���ʊ���ː���tk�W�o/-����a�wK�=��L.S�Ǘ�xs6���U鍗�,h�H�̨�1�S��m!u]�1\��ƻ��}wqU�ϖ)6o8�k���>����=�޺h2O�ϡ��Aٽ�3��5�:Ec�=�<6��NdwD��	D����F' ѳ��o"�&��b������2t�)�}��bY~��U�˻[֯}��<��ȍ��l�I��a.@C��%8~�K!�W��Z�l�ݙ��eC[�H0h_
9x&�r����>Gu���S7�;�^�:��%�j��g�:��Ϫ���e, j����^fs�5�pb�oy��S]OjbnN�j줟[��̮"���b~�ր��T��J�r�w� y�X��$�󄚾~y��GNF��}w{�h|P�/�	�6��iah]vK
-��:� �;	����}������aA�M���eL�n}�+�Z���j+�q�b�{�7)t�y�B�,��T\�0(]�܎]]j�0����RΊ5S�[�
��MDxy?c?F��'���F���13���_�E���ˏ�w�z�!�
�e�V|�����Q�����#
�U��|S�Ư4��	q��j���DȢOshᬤ��Y9��I��ݡ��_y�9>����x;/�U��u��]�!�9�0�8p��q�`�#q�I�YZ��ѓ���+0��՝��Pea�f.�Q9%����҃R�\k	�B}Qv���m�u~��o32��޺��ɼ]�Y�^q󢡭*��_gȕ��y<����1�DKx�	e��l'�W�=	}�}�US6f�.&V6�-7GH�"O�D�`����C�0���˄ۥo���Y�e���׏�iK�e;�{C��9�<)q�pnO�%�o�O4ʹ���~�;<���&�he[�NrX�a�}��~v5u�9�/��|&�c�>�m?����R��4��Qb]�2�ݚ윎V���F������0�9�y����軗u�pe������kn:��n����م����ɈY|ӏ��:K�㭝�c��l�ꉑu���ݯ\����_��P��~��u�_1͟���ۨ�OӼjh�݃'�TK�j�v,��s���B�r����>�^}~BlR{�)�5ǉ0%D_�N�� ��������ӻ��^��Q�����J�j��3a+�3Ȝ���YE�=���}w�8�E*�K��a�eОT�hŉ���F=��NDQ��H��05��c%c��C������G�Ӯ�EF
� ^��35#v!z\oD��1�4�<����|Ŧч����� ��&h���Hs��L�T�@�M)NI"�l�/��OQM.v=,�^u��hgقe��Y|/�350�AB�3�V���E�N�>u�7`����K$����ձ]2�M��4%H��\�]R�A�ndwnRށ��҈=��C������7��5��,�Aj�ID��D����p+V���+��퐞�����l0���g�(���kK�7r�V�~�S�2���oeǷt��B�t�+�N�?��"���pgL��o��� ��@�ʕ�"��sdM{��h���v�E�VurN�5�l|Nd�!Z?�,$11s��$�3�uM�b��sg��|�x����9��؄A��s読�
kv��F|��+S��V��������@��fY��>�1�X��tݟ��$]`�f��q��*δ��eNʮ{	#��e��g�	.|���_��|�'?����r��#��;1Qq��l��ޖs���7<��	�b���.nf� z�|��R����~<=�j]��*{g�L�(5�$֬�ft�iKcx��wY�ݕ�5Fא��s׏}�!b� Q����
�+\;�����Ĭ��2ID��1k
|Ԡ{�twEN�ء������[�O�.�V���2F9��2�;������}e�9t.��,x=��NO��-U�樄���{7��0U���JYog�o��on���>���Q/�]�ld�n]t���b!Lɠv;���,�y�2����~�R˵��Ԧ�F��1��A�42b��C`���$`|y���4>d�_��8yTz�����y5Ed�{_�6{ �m�n�4�}�Gk����C���
g��'R3	�3+-ˉ�N��,`EV9��wA����� (�Z�'wi�E���|��V(4�FG�	6t�Z:uD������M�b��X߲K��N��Q�Xۢ6-=��x��t�21Q���8�G�{�xA;A����&��"xv�4���(��Rc�^��0���������Z�gȈ#Z���z=�@ӹ �Kg��E�q Ҿ�\<";����d,�>>�����P�F�b*�@�Ϳ
�/_d[�u�7'!y�����c]C������&�<������-)J\��=Xf������1yf�U������P0f�?�Gg�����i1�	\/�� e���Q�}��GO)��L��F{�Ϫ�GK~}�D�˝�j�ٳ�Y��~O~�������l] �>��������Y�ތزu��~̟�?����y��_��԰�4f鑎�%�����%;t�1O�W	�֧�B��9zz^�v�iMd�9v����Ik�be|~�S�ܬ�-+N�5�'�b.W�ekYM�^�~I��|7�M��Ǿ^�N�l�.�*2z�������nZ�h�ږ��!g!���Ί�^�����_Pܟ8���S�^�i)�lO�q{��3�]�+��eOv��/����p�p�
�v4���JǑ�"%��-�jMns��ڣLlU�92ԕ>U»����'yq��:��^o)r/1�wvo�-�*\,B6���M�F�������������n�nc.��B�u�"�]��u�[zBע֍	7��#����2�}P]],,ӿ�BQ���c�f�g���c[�k�.�i�9IsW�Y��&�t��I��+<o��j1�=��c[�f�km.oiI.�q43��Q�$(�E�`:��j�NX�T�9VW/�Z�vc%V>Y�>�����z����NCD�q�=�׃�+�\
�k�c�U�j5#���\��4�+�j��3�e'��&��k|^�oʅ��-y���í|���E���/o����;9T��x���y�*�$4�x�^0k�;kV*�?R�m��{IV7B7���.��v��Vbb���&�"&�i&��� R)9�z�Suh@�[#��^���(U̡��U;�rv[��t��=�"ڬ�un�1�8�	C߮4�oKĹ!L��}O�����b{��́`�'��2F�S~=��Ok��C��n.�>t׎{�g���}g}�k�G�Ѕ|jyȺ�v�_���N���XP��פ8�U�/2���������z�9��(�ߖx,%���{�i,����%i��?�7X����+��1[� �C�5{v��M�ퟡ�r�VFJ��O|�=����Ǔx(z�	m|W�g�-��z�l����Ի`*LA�w�l#s'�����>����b���V9�q�G��$�H�MAZ�)�^0~�}�U�wI�{��%���Z٧T��%��o���z�q����nt���'DQ灜��Nf��Sr���c'��?�̙�jE5��fl`�u�]�1!\�t2�fi�:Ogt]Ӳ��
[&u�5|��9��i���Cp,�}θ{�f���"�.�r���Ng��l��W��.�-��d�!4�@�	�ĨF`��++ڻ�Jm�;�K.Xݐ�f+�j����1�9�rW�)��T̺�=w��]�L%ܸ��J�����c��DD��B>�pԾ'ɜ=�}����>�L����6Î�c�C�3����W�;s	َ���w����؛ݽ�B��6Lf�]Y�5t^�u�_V�D���덾������+99Bf/��0��������u��{�9�\z�5=��p%�-P���rj���Z��ꏧm0`¥�������6/G|�����IV�7����W}���.]˗�m�p1u�\nLOo������e�+L$v��tu�?8�bq�G�x�;(�H����$���uZ���R��N�2��,u�*�;^��<ǳY�oV]UD��^s m����VZ�Y��'*�9�����Uw��\z�T
,7���&�\E���b6"��ܽ��y�����6����2:2&cF������J���:d�{�����VR��õ)¥w\.t���;3p�8'��-+��H {;��{���Z�e�e�;�8�d���[��0��0���85�k���Yн�Oe�]�:�<)�]��,<��s~2�V�# ,����랯�8�n]h/y�����}D�=~?1�W����I|��q���z#$��ض������f��eh�=��/2��ުhv��t�T�p�k/2|Ȝ�%�~IE(Q���� 񪾎(��A�%���3��F�eེ��o_xe媣�z�iM��I$^��t�������m����	+�V}���������Zu���[A��S�g�-�F�ͭ��2|)�/��3'_O�F� %��)��t�{�	ʩ���o�0�ߩe�	r�_}
��2��6W��*��)m��;������eV��[�?�;);��Z��9��1w��t�o�P��9����تlu�Z��=�{Έ��ni����egۂ��@Pm8SQHZQ�)�"a��r3x���0G<����З9�#B��0�in)�W!����4��z��T��)�����D&3O�t��M{H�M;��6��	Rԓ���p�ScWo;�I�O���b��Ve���a)[�&qlu�@A��Y���h"�l���i�6��a:5��y�>3�Kb�Z�,=�J���uJ���*߻�K?<���%���]���t��7B9��e]����Wy
<��8��pJ�kD����ȸ�՜�J��7T��Զ�U�W&�,0��N���Ҭm�h��f���;��L)*��h�k�U�ߟn:���3J�P_$F.������*�Q�����f�����)ߞ�.�A��RY%TvT�P�b�C8d��J�S
�f9mH�N	����Q1��m����e�5�c���U�>gAL���Z���1��P�nm�'J7�`���첨�(�)�5/�������W���f"���n����rxB�Ui��p��F���zΕX�0�e�.;J9���T�w ��U����ʾ}u��qnC}��>�*Ɔ9���/��?���c����L�g_��.N���G`��̔5ݸ�6��n�3����[�YFV�K��q���a]�V�ڱ�dd���j��r�߅qǦ;�t���]CE��G���f���ml��`%Z�n�W��9��N��SSyH]j	�״��lA�Ⱦ�홝�����us���&���l���p��B��RTfٜ�Ȇ;�1�\�ٌ+*C�{f��%�1W$y����j������28]���W�s�nN1����7��u�m)�����'i'6�ݎ�7uj�%!�v��u�CϺs��>�4eHs2���]:�x�l�V�oPO/����:��n�J�i�1S���@qd�z�5j�A�$9{�KW���l̫]Zd�yٹ}���$�/�*��{��:���7N�8��%�[�_�5K�c��,H����v��s�p)��+��,w�P՜_\��ј+j��n�r����D�w����lf�l�U*j�1���eb�.���gU�����Y�2�m��d�2N�Vt��@��2�����0;f2lgV-���sZ��SG`�i<zp{�j�esF讝���m֩c�,��B�i�7{�W^B�wԺ�AC��3f1U���NƮm�f���+.�]FSr�$�zz���}�R����j�`�x+.��C�~S������~��q���G!�-V��ͮ��f�u�n���9:��^>�b�Rs����E��ڣ�*b��j`}$j���W�|>��X�׿�sI��.}�5����di�ߟ&�����o(�{br|q
�#B�$_NC���2üa-������|2�ݼ���>��!�^�����r������Z<���t܀^�f�M�j����ߤ��7�Q���u��"fϯ��M�d{ZO�-o.���V�~��SIw|Οu�We�C�9��9���R��1�I?c��:ϲ�N��q5��S?v�
;b�����|����{u�ɴq�k��|���8]r�컾��u�#2.�s�mWވϔNf-�i}����4��}�FJO8A<=�t?��^�F[�A ��\��3*~{��ۣ1�=r���{_�G�޾a�wLٺ/�l���ėV0�����}�M�A*����N����2a����Q �3�M*�����{���1������`�+��������YY�$�@N8r�̺>;�	k^x�٧֢�g֎���-(�X�	z�!N;%Jcۧ�����껷(q�����A���U@���~;��]��h��tV`{���b��[I�$]L�R=����/���z�C��H*��5��֑�Q4�]Һ��D��	�*�ռr�dEK1χ��$4�kq=�d�gk����F]I1k�ɭQ�V�غ��Y�|��,�i�Mt�/ace6���)���J�X��"�&B:�1�f�Kq5WY&.���y:��Ӥ��'d��72��s�����\�K��V���b<���_�yj�����d�%mh�5�][�Z�B��K��z�#�ძx??8~��Sj���x񏤅1&gg*^���V�D����\ق�@�W>z����b8��{���p�Ɲ`sC��(���&@�
��$� ����[,����X��߼]e��E7���T7F__F��a�G��T���g��P��������G{�^s�T<~�@m�1T�ϟO����F��G��%'I��D�iN��q�\�>RzqE~���(2�5x��aK��M�hn�Zi�(ӑxL��'j�}K�]fw�cbL�WY`�܂w/��vo����ͥk�g�=F�j��γn���Q�%�G'ъ�11v����M�d��^�W+���Ė�O���B�ꤪ�c���l�c��c��_�_
K�I��1�.3�Ș�T��58�Ҿ�=rw��������e؁���(�V�ɰ|B!�º<q.��콟�H%{'�.��A�E�uڧs��:�﮳�e�x�kL��E4�5uqFtIEM[7.
�e��D8��1��݉5� ��^F�܁��N�*�s��q���Q�f�s1�;�\�M�ϽC|��kӦ�W��5�����u���.�t�L��Fw�;��/��/U��}�<f�Hk3v�u3�����?1�yU�K��oU�&�՚��ۗA���};����v%��Q��W��S�����՛/�W�h���e5�d�{��
���_�ò��u8�W������~��j����0T)V�ԼT�u{J���{�=[�6����F6�Z+-V��(���'T��A^�MEdB|�\�r-ْlc�l����e����k=c����kM����k�N��6�g����""����`�𮟔A�iH2OB雉F��k�6�n�Un��}qN)�O���ge	�ؚ{cb6M,�WN�;�M�	,�IZݸ���f�Zo:�������1k*��E�-J�f�.�ᑓ]���1vm۲~��6o�����=���|�Y�������h�mX��߈�O�w��(:�hO��|������w~TN���r�A��F�!�-�˵SX�辙�V���e2��h���hC�tu=H�~V3�����r*�W��ֱ(�����Z2<W��hnw�	u���뽳[}Pi ՙ�`��TU�kZ3;̈́�V������im���9];P��;�@�����;��s���0d�ËF��۹2��ޜ�wq��w0��)z=���+a�S���*I�1(/	^�ݹ��k��V�zN��U��������{��8vsў�"�\u�����4H��ז�W;�߱�=��DW����s�C�V�k>.��#�͢$>�7��tpWG7���>�Yq�����^�����0�z<����WP��p^�=�5(u����<�h �y���;Ԥ�<��b�ꈛ�M�aý�>�()txFӭ�^]	�pv�9�[��|+�1x�^��r��9X<�=��2jհUײ};�;�=a�[�.�k�L&�Rm1�/�S��]}�z+�.���k�.���>��X����_�̫w��\�y��q�K�'bZ긪���**jv�]~�MI�66�m���N	
PE8Ra�̅ȓ1�W�f��.�:x�f�K��B�O͇�
���֠K£+c6�=B\o4�5s׎�[��UA'�Vڻ�5un��	�4zӰ8o�p�N��5f-(��ogK��\��Ԛ�\�/+�V�H�k	���#�B�}�?l�!���~�7��d.d��ޫ~��	zR̙� ��ͅ���Tts	�ɗ�.D��<�V�]������3!>��J�mp���=}D
�4a�l=��6�gY�t�`��n�	7��&�;�c�/���3��;u'��:����������K��#���s��~�����y\v��o!�Q���<U��n�r�QJ�O�d���E���T���磏UV]�����} k��<�D1U���l���a���t���TTj:��^z�2� �!6C����+���~�baP|Q���D�]���"溣k �����#E�ذr� �ٹ��]���L�����4��M� �jŠөO��Mx��\��^P���}.����5"1�`�")@Tj8����W?�l���k�ѳ��yѨ��.!�ҡ
#}S�]��I�>�:}�(s�3S4�D?u�ܕ�ð�z������{�?�f*:/9S!u�[ڼ�#�/���%3<L�d�q�|kO�b��7ȯ���O���>7,��}h���Ƣm�����2OA�X%� ���,;^�!��Ǖët���p�]U���j6�z=r�'\խ;�ф�팖}o:yE6���&7�˯r���+�����ym�s����(e擉꫇���)z��o��q�U����sD|�r�;�G8q]U��}�"�f����8���F�2�םŶQ<�,)�c���k-����[5J�ӟ���������*�_�ʝp2�I[�?!�6� �
E��&�f��JHA�V�{$���i��n�]-�#1R����f �kd�-��Kuԣ&��潮5�gK��FYy��ُm��r_n�rV�������*]~�aF�;gzv��ˎOs�N��J�C�f-�^,���<�l��d�
'���m��r�~�*��Jy�ntmw5�W�ʭ%�� K���_�(�X�z[���~I@6�~��l�`/�6���^�v�k�l2	��*��"����[�6��4͌��X�����/Lz�|���̨WÝ`�1'��>S�pnz���'���TV}4:3� �D�����>�/�l��gxWv���}���|/�vN���p�m�|0A�C2@���¢=5�5�b�zΈEel�\����O̅&�U�z ������w�G��G�<%�*fѺ孊E�i����w�i��m:�f�ɭ�k��N����EP�epf��^����r��g����U.Q�M^Bl{O�2㤞���O0[|{6p��g�H^s���^\�+�g�7-���$V��E��1�NL��xq̣���f�WJ�f&+z���#�c��!� �uS�*�gE�vV�|&t�bY�
�18�t�=�Xz���zua�ޭ��,��i:��:���H�+ D0�$�ŽZ2�j�}��إ�2������B':`���4�� �l�����^�W P@+�����[uT�/K��4|��3�yH	����:i�7
�H\m��B�q�[�Г\i�C����*#s�\*g��t#�wR�:js�:��xP�h��7T>v_V]��u�/0�i�E�]>[�*�nd�J��=�]jj�`�t��l��e'�n�jb�g����.NV
��J7�8�7�� xt� �'�d�	��g��({oo)�v���FDЬ�*&�V��r�3���]#`Jr�G��_j+K[�dn{3��_!Z�ߴ��L�G��>�9���b�9��39%�D[�����1}5]���k�#x��.�.��uw����z�q=u��f}T�T��\gOT�m<��I�v�J�_D8����TFߩmj�:�K��_Ǐ�(xz���gw�w]�X�)�ʓ�H*εwau�����xF?����v���yٺ�������U�l�Gzvu��蠐�)�	?�jC5;�Ƴ��~�VG�C��ݗ��ē��v;�Y;��^�?z��vm!�6��"m��i�J*a2�Rc%��S��ǂ�I	i]5�e�Nҭ��iFɔD��ʟ2��F��f�m>�)T+l3z�:Uc��wS2^�Mb-e`ٵ9S"mc�8&Õ)�nЎ7���nu;ը����N��6����
bw�[/}~NϽ7���v����֔��Y�=��EՋ͆7ζG���ig�|�0��\���h\4��2
�W9w���o�?|���Y�p�C�갏p��u�'8/���~�[��߇3s㵄��ʽ�����R�ү��~����v�{t�w�-.��C�L�{���*�\V��]L.	��Ő*.�1��W����E��E��^��ַ:������BW�YYU~q�<W��t��S��%�e��^D�7����
��n�ּ�a2��<�-��(���ݼڣ(���v����	����̑"�_�=�m�Z�S����Ԫ���~!��	��;
%���i�	JCٰ-M�FW�5��;箫���J|v�^S�n��dw�����u�	���{<�[���k*��vN�WYo`|nN�oD�	k�t�Ǐ������1�㦮��d�.R��rD$�
�b�G[����t�m�5B�k}��b�.=p�=�}���~���br���p��-�݉-��q�'���Y�m�@B�i [��C����W`^C���x�q�-X(WC%�Q��9��ܻ�}���=�&05�IY�Q��۳%.|:d���m��_5��t���>șP�!�7�������:[�ȉ�.0���4T7p�kr���8r9�TUa�"��(�@<���(���*��#�N�9�����LЭ���g#���h+$�w"�����j˂���nYg����a��\��`O�&���O�ᬵz�W���SW�ܛr����p���o,m�^v;�}_;d}�~���ʈ�Y�z�"�-�%y"��cT� A��%�=1@�=,�U�HS׽��ƕ�x��,�Q�R ��[ ������2�yd��:�/1�g�e��#��՚R�c�9f��&�/Vv����G�������}
	�"D
G�hYV{��zd��������
�hDl٭W����7��G��R�zu�U�MӟMk�~~ZT�ܣ���g�-����$����;7Oeuq��SX7w=O�n�ݪ֟�:�C�3<��|~Í�u3{�6r�r��*���1�Ջ7UgӞ�'nj�G�ߥ�"��f<I�E��{,c�L"Nꋎ +V椟l�//�%7���U�1Y�i�l��V��dP���W�hH-B�+��^l��gU�恝[j�$ѹ$�&�fv5���y5�qO��_��st�f�s��Р�����zm\��;b]wl�aũ��g,�~�����^�eΓF��,��)r�&�e-M�s$+ �rXfl���l�Fa1]r�I�!aB��"�0����@�3��\�]d���W3s�}�br��x���I�}j�CȻ���<E��"����_�o�P3�0���c�o�{�/ҧ��̧�R?�U7�Z�K6W�$K׀%�fsC�c������_{+ۉ8HP��Sk��0�=f=ct�gO\?�1���^���f�e���
4����' N@�P�v��;�aV|�r��&*��W��}�0J$���Jd�
FɅ3[ȉo��eׁ P��8� ��[>X�D��6���R�Qv�'�M�c��ځ^D�R�b�Ϧ^�΢�����{%�})�Ȼ�g����k}�$�WG!{���fO8������Q��fw�ƻvg��w�_�
u���P��y_�������1��4�E!O�9��>�Y�|��^	����>���h���Awj݈��V�\�ZAb��<��ަDd�>�4����5����<B}�"��{���J=��P�
��8�d=��C�{ڦ���{�������}�da��, ����ߧ�:��xw���C\�z�W4�wtj����*��.�"pyK�f軕u�1�$�Es��M
�K���n����6���*W,C ����Ph,����B��k����n���7y
Fm��D�I��C����:,[d�lh��	�kX/z��������Us����>���R��F=�f�L�T��>|.�<�ԿY�b����vl3Ý�*;��L��y�VNљFk���P7���ߩ��l�@��׍^��~�d�*�`~�� �-
�&wL?�mT��E�ҭy{~<�q��C�#��ﰩ�^;��p�2�@�(��{�WM�FYa��w�x�Ɋ�re���6eMa~ܣ}P&C��T����2�7�xҖp�]Ot��SԫֿN=���|{�E#����H����'8:��FU���Y�Qv�\�}��������re��h��gr�u>Η���c8�=���p�)-=Vp�ѵr�-����dF^��x��l�|�XO=���1N*Qa`3�.���P8����#yk��)�<a:�p���]d�D�\�꺕����=����J<��bh�;�{(m+��î>��a����5�k4��K��X����:���:���ڳ1��v[gS	��`o��ߕ�O�����wۀ����g���rfF�'�(i�.p���m�r�QoS�8)�%������e�r�{�Vf��vz�ְ�я�3A����5]4+�KR���˅\/��Z�%���\C�$�����{��=�#�Br�L�Iq��:�`�fVMU2���U�h�$����ڮ�����-�:�.�^3��'BO��#&�&�9#ICI1J������˺˺��� II$I;m��mI��m���n�ݶ�ĸ�n#pa��_f\����_-�$��j�IU7'��N�^�N�=���d��Q&�!�la�0v
�s{\��y7GNh��(R�8���뺺Wgi������E��L�1��zo�ESRѠ;�@zk�nr�|(\{v8խ��	LsN��"��aL�:[7}���E�r��u��݇@���PvX6�e�h\��jK��
#�+��m��^�������g�Ⱂ�h��ӊ�ރn�-hPco5R��2Z[bt0]�Z4x�X��P��1���n�J�oj=��s]q���:��8Xh�I"�[mr�ˏ*LYd� �n}I��I��6h�FDJ�
���i�b��dT�F<��Z�2���l�/�������R�IZ��5wKl���<�B�y���l����Lնrbt�t��ntԺݴ����Sm&\2�6V�zj�X�F�ng5��7V�Z�e�<��3�c��&ʷ,���eD�u7�&�Ŧ�GB��������OWI���}�/�I�!�f�7n�]��Q�g��];l�d�k��].�H�:��ٺ%m��ͮuv��A�jBŗHkl՗cCGR�.���ݼm�:bΩm�4��iy�$��<�xX�+n�Y���b��g=*������r�:B��0נ�j=[H73E��L˝��srA���)Z��sD��a��M�ɋ&��.R�U�R�]�5����Rs�&+�0�П���gm�&����1�]�bY�V�J22J��%�H������ێ��~墿X�[�҇Zt��(n�r�C��v-+V,�.]�4�'�Wxw���+kD��'�]��˅AJ�^6��\M�{z[}���":J��Ü�r#|ñ��/G�J��n4�T�U��K-X�{,�S^p��}̻x�����������Q����/�z��м��'�
�/��k+	}Ï���̏�Kayuk2����h�P6pH2�p&���";&Q��D?��~���x���x����]���f�ԏ#c�ڝ3B�9{o3�I=\s8�4^����vr�\p���2��n0{�z�8Q٘�u.t�#�D�f�k.�����G-9x�]���}ly'�]��W���8����]�D�̃������/���mه�=!QӹI��}���A�_<^�~N�=�Wxmj�����u}t���x�3u`��朾⛝�E��}D���_�5~��Kw�-7:��Uc�L+�>���TNE�Z���>���G�u΅�󅚮7��{w��Y�í�&��5b�s�w��{�Kuz��,q�wū�:q����ղo�,��(Д�~�}��}F��x��=bB�v|6�/A5����`m�o�}Qv�>̢Y�j�Y��3���?͗!m&�rB��FB�*'��&�=��Y����>�;���Z��k�Hfvݟ-�P�>S4�"1z�s}���kE\����1uf�6-�<]�����m�ܢ���A�m>��8��9�eqq
�R<�����I^I�yP���8��b��
���ާ�v}'?z��}�:;շ�4F��`=$�Yʕn���������TH�Z��GpU��UV�Vh�&z�^���3!>�\_H�<�����
Ev�.�5��鼿�	]�N��NC���qѝ��{�wd�n]��mr��_PѾެ�����`�w��2���]rD�ݾKu�=�qv��8�����3'}�\&�=�U����}Ȕ����+�7M�	�+�����U���s�#�؎��,CӾS�.\��o_ћ����Y��M@{>n�D,R/uu�����{q-GL��"VVzPB�,�:�բ�̎u�z���6�^�YwyE^N�jti�W�5?wnɲB>��n=R5��e?z�G��E#��D]����¯��a-�ڑ��d�M(.~�$ޝ��p��
�^�2t��C�K�1A��g�'6�	��=������pe�����r^��ӫy��3��9��}ˋ�����E8������~�u��m����m�|^c��˼ɓu:�vW��dq��7^}jEx��{����Z>���JW�{Yx��g���ن��շ�^��`�SM_Z�i�4�yT��+�k��g\����l�����{}�"���E�!�0e�R��q�w]
����7r�.Q������̗�-����T@ޒ()��:pn�z�W\�Ͻ�.7�7�oJ<�h/�ez�o%�L>�����7S7���NI���1��0@ W,�gEu�K>Ş��b�^t,��q�8ٓƴXJ��i������X��s䪼���������p�Cq�>W�91�#.�[���u{�U��w/;�h�S9����	�spR[��w��f���ʍ��5.�������MڭB��}62�bs=C?}:�����O�褯O����>f��K��,�1�R��)2��I�U
��;Ǆk�b��$^f���c��-.���q>utcl$Nx��P}0{�]y�̘5f�B8�[�~�K�n������.*�Y�N���u�|�4�}7��p7+q@]���i��@k�9~.tL�tM>����"�:���.w��ܰ��ϽYob�k����l/i��,H�B��@��cQ�V�.�����UЂ���p��5�c��Zz/�=�*k�J�z5v�q]xW�^�]�|A�G���v��&�������^�ŖvKH�`�Q��]���d��oe�ᅩs�1�H:7jȜ�wB��j�ѱb긲H�RU����p���eU]#$��{]��v����T0N�D�\�ި*��݂�;���D5P�&�3��6&�+T��K}��<�X����<��O���l��mEu�f&�ecԒ]iv��V��i"�j�v��ŖH�"Jq3�e!���yb��]ם�Lһ>U��nw�4�̄�^�%��G�|4������}*6���ff�ݾ��n�^n+`�!_=��)2������g��WEG'wa�C�V��u����{��̚!>ݵc��e �>W�0^����g�Bu��(�r��*T������k�W	\iI2��sNJ�7���r����㷯2�{=�i�s�������\�I���؜-U����}Ej�����U��/ܺ�'|�$��˃��5q9ww�����������Ƀ�4�d���s3��_�#� `�rrϯ�L�U��`��rUf/_��`�bڗs��� rxND��\)��S���MQS���շ����l�̟����!v�� �T��n�Qѩ�Y�}̸�����wNs�&�s�J=��.�G��n{o�8T�g�1[�+f�]�tN5;��a!�Ѿ[P#�ݭ�7�ӊ�c��Ft��\���_vh���nt���Eԛ��\x5�ъw֥Κ.켝���}���ڳ���V~��.��V�?VE����tr��뻯�,�r��7y�A��w�vmen�&�gS���&�^E�$3t1έ�7u<�}�p����Y~#���g�q1��_�N	<����S�X��<�����1��1� L%�Hgm�����V`����EpEϺܦ}*u���3���z�y,���~����U��ݭ}7���uTX^�J��%^�w��ھ��K�뵵Cv!*��eG.@[�.���"�UX�8�)G���->��>B��>�D���I;���)��.wV=fL���{�Z�˫k�D�v؝����9����ͥ���� [Z'�59_Ռ����[��ƻ��I9]K���>��VG�����]���]s�s�K�@𯋢U���u�S��Ծǔon���*��5>�T�723���ºy �����:�"�eDMq�y3Ɠː�ć���E�`sx�9x^]=_��+������R7���W�{�CK�t)���|ἓ�}��q;ϼ�z&��|�G	�H��F���V_tT�O��4��چ~2�
$b��#��JH���[w�O�{�u-��h��T��s3!�^����
��bW�KEu��'}s��PlӷF�;�[ҧ71-9'rM�1e��N�A�WD볢�V�����VA�vE���bN�6�-���� ���p��,�t�w�c���l��o��Qn\�d��ݿsӟ|�^���%G�O�Z��ۼv����\�y��X�.��P���<������;��ᵛ<]-_Zvv��u�M橾x��6�c�a��{�_1�vQ̾�B��6���K����wns+Ӄ�1�#z��7d�㧐_FS;��3Ɛd���G��jf�rUf]�f_����;���l�������VC
���H>T�aO�OT��a���z��!���I4�溹�,�[�"-��{Z8$�[�u�x��F��օWun���}f�FM�'�����J�m�eø�5i�t&��7���g�{��0����Ͻ�k�/~�R�'��ـ��#�uw_�3٦kiuY�9� ����L^.��S��4'�4�A	�n@#�f�u���u�����n'�5�~x<�ó�y!����!"��ϱcL|��zX������X��M|�gY�����'�W��}����@T{=�eC=UZn�7��S�k����ϙ�v3�إ�8R#P8]T\o�ekť��\�b(7���)^t/A	:9C�}J�f�V�R�N��ZY�.]��"ú������F�!~�m7��ܩgW�#�"�{i$�U�K�wu	�9G��x%m�gJ�g��rY"�Ϳ#�!q��ꘑ��AqwT�����v:/c��ɨu�(�Z��'<Ļ�;���r��՞��[[�
�Q�j������t����c3=\�\��\������v�9
���j.�ܨ�B*K=հ�(���KА\/̭\*|Em-M�����㶩�!5�þ�=H����=��f(�?���_,@}��As����5f�9>�Zf�'��̇[����|<z����=�}*�XĴ}���[��G�}i[4Y6�&���2o����Q�_?�y�N�'8Ts�:_�c<�H��7�=_��]���ئ`n�E+$������C�}��g���G�R.���&�<\T�p}G��uX�[�c5��WKp�8�"�P�B�Fx���MC�s9=�;�+F��F�k�2����	�g.ُj��l��!�ϧ���W�lh���Ĩk3��?�W�N^�z���'���
K B́�Qn��?(J�]F��O�	��(��5�Uuлާ�ѝq#�������z���Ջ�Uf�u�eN�;N뻤d0�<n�\r��jɝU	ݓRw��Ђ>4H��W�5X�w�
�]A �q&9gQ=����'�k��s�|:�/t֥g�:�pT;ɠ�cD]-�&q�ҏ�Һ.�&��e)vm"Kd�å5-Yv4�b���]��Z�h[�%�֖[��T�K�Է&��\hp��dƧ�bG�uא㔌�a�J�#+m�c�/ٌퟬC�e|��W�tɡ2���1��\>���w�T�qL�{̫ V8��;�n�������5u��fLtF��D�cчY�1��w�P���L@K>��E�`���2����ʹP��w�c���ʪ&�;.�-�<��3!�)��I���PD��?}+�����z<Jn�o����t��3ƀ�����/%%��t4��=�*E�ca�#TTwpډ!?}�%`��Nz�	䑯<�L}F�o�iT�HE=���*���f���9𪥇��z�Wou�|�~{�!h\�=~�$���Wb��X�(���� ���
|.='��w�//o����|ɛ�w��*^���c�7<�%���Oנf`�I�)��|0qh�����5��2�29��c,b�*ʞ̺��}��Ԧ�����7`�1뽸�..%NV#e�̆9L�y������n�!,�wz�X;Ӗ���2�<�FR�h��J�~<M���w��k�R�&O
�~v9d�,�H<�!W�mb�ov��M����gN�S�F�=���gkZ5�u��VzMxH\�,��$я��Z[�jej�ɒ��㇏�$�W_Nحz���%H5�@��D�T}�����	�C�.��fly|�g�Ai]{iY�Å�l���4��m��׋۽���B9�N��E�:ȗ�f�N�Y��&�i):�������:����EfUlO�Fuz�m��z�"���H��
e�i��A�9��s��*w��}V׏���wjf�?�R/��s�iJ�@��ޅ�Ui�^����j�W�����s�;\����{ш��IO6���yJn<�Rw_V4! �����Z%�Q�͘Ǝuƺ(�l�u6���i��Z�N����|��}/�y���Ϯ&��ʹ�8;<�[�A��ZX��wr?��$�+���!��(ovu�ǹ&{��`��:	��ak�{7;[��:.��f�A7��5^���W.�G�uR�{�z,�8�nQ��uOm��#��sԧy$�~B�X 
% I�	i����[���udCPA8<��
��l����Z�}�N(�S{=1����n]���3�0��J�w9�]No�1@�{-�6�E�j��7���b�+9�.�;.`��ge�d��(�з�����ZM��/o;d��*4�����3�Yk�AoR�W������b* �s��+'VԜQ�O-z����̺�oj���Q��T�݂�}Hl�5-�=2��.o���p���m��g4v��'��O��7k��2{�j����û�l+��5�){���%-׊�c�Ls��᯾�7Ϟ���0N\u���39��{oם�7`�~⺳i�^Q�I���[��[��}�}�t��$5�>q`_��^��4iA;?U��|����ΒwMT<��k��]��3��������m��u�?%�װ}W�6��g٣,rR�(2��p�?&�	�dj�����z˺��ṀVNG�P-��lTDj�:���efUI~}���>���]n�g�Sd�mVs�	9�X��ݾ�}����g?��Hg�=�ݤ���Rމ�Ab_��(d�{uz�۪(DB��0to3�Ê�����s]EE�c��;�>���=�����{s݊?����{U��Q���b�}u>7�v#s��1}���,P"`'Z򘼛3fT�v�~V����e&�ue������Ic��f��d�ċl�s-��1�Ϡ��B:j���N��93p�j[ ��`�p]8;+�	�U�f��L�8�*�3��̎D�/`��r��3}^TMp�o�xL����:�f;{nڙb�԰ �[����h�R���s�}�I�s��z�9;t�۪������b���ʰ��IX�&���v+k���ld`V�wʊ$K�v�w�O<��������w�|��J�����~�Ҵ�]��)>6�v����� �_�[��8���:���������ww)��<{�S��?4�&<�_>m�W[��v���p:Z��U}�b��7��-��fX�`�zF6�l��4���<]M�.�qgUxhڦ�S���%:��+�]���}�����ea ;N��NN[X�>�2���Δ�YKO�{;��amu8z�[��Ȣ՚n��vR��^��b���"�t�M�l�a��V�$I�+���r�f�4&U��j3�:�?Q87�]�y7�����7�d��'7��W��h��%f]�=���g钧���@�t�mR�p6�fv��F�A�ֵ9^�'E��n� �����;gA� /�8��,���N{Q�Vk�.�Z��T*���܋+5i!�d�������[�Y�W+�E	'WP�痦^NK��J s7x�ٽ���E�y��&�
��B��u�f햋��x	6�V��#y}�$u��o�!��ۤ���Y��V\Š��J�<x��鱸e�W��$������].Z��1�m�[E=��v���S�&�ή���7�!Ȟ�-;��C�M�N��x<��K�1d��#Wz�"Ǉ��c��+��<�,16�q
�4��e��C��[r��oK� �8��pǂ�kW��bt��YR /AN�]h���쫲�X^;��gl\{��w��fK%�؀˵q�`�z+8a�ȫ�@\1�+ASQ�ɦ
���#_.�V\V��-ڏqģ�n�i��P)�.hN���.V�/:�j�L1I��E�����>���ԹLR�������p��9vq�Ξ�G��tyyux[!&4��,Y��ԥ��$�����Y�]qC�����ꭾ�� �"�K�ˊ�(���o|�߀��9��R�XTew�qF�*S�|:�d�wr�]�;{�E&�};����oAX�l\��^�6#|��W5Uv�{08ߨ��yN7�@ȕ�ײ��n��)lw,�`eA&�!R�=.;�=���f�e�?s.�O��C?GE4,���垚�o[�G_�W�=��lq�+��a��g �St�O(E�헹���L�]���;�/62������}&c!�}�}SVu���G|I<s81*��W�,��]�^rDe�^O��dOM2:���kV5Vى��൉�^jm���=7r�6�����u!d�#e&��j�.Q��&0��o]����6�.����l�*�p��a�_U�޼���N	�K��[�|ޫ�ګ��'v~
�����Tq:�6����>3B�?n�� ��=�j�+e�<�������,s�Vd�w�rQg����t�l�"=#��O�������!@���ϰ]���?�|}~��{[�15+�����}�Q�_U���r�Wr]���zi�{U;��:�$�ηw��
�Lx���f����/]����;a8YY��}0k/2fi̮���6�$���[Vi�I�m�<yB�gw񈽧�O݄�7{���L�{g`�/��z*�F�nh�yg%>ףN�iC��b��&*��&�qi�%u���[9�M���|���K�d�`tԍ+�䇆�V[k��K;jI���Z:��#��]n,`�]� ��B4�D���Y�u}[�wu��\�]�a��N-W�=ءG!9H��"��X���`�&�4��I{7����\��ÿ|��E��Uۏ=7�Y�:�`#�dA2xvoў���N}����Y^����.�#d����|/�|�Â��]O	8$�e����|Q�}��{�y�^Wj�D���	�?5�4��~R#�N��J���R�����J�~V9���U�0�����n)'ݏ�Q,�Dȥ��Ԙګ��l�!���Ky9��#HW��:�����/��1��T:j�|�n?R�����~��/AN;��D%|.N�9\�+iU����4����b=ьwsۊ���l*���ٙ����t_�*�,>(d���G�V�ɍ/��YI;��IU�BYu�~͚�ÿ\��-�)��O-e�H��Q�������걏����w��u�}��ȶ��jq�ޢ��~h�һ�1U|rq�@/A��3Ngz�)�x�n�ᯡ,24�&�+�D����J"���l�����J�GK���\�{��Q�&�vm��4�T1~�Օ����o��d�q�ۚ�m[�����t�]�U=W�6!����,�9�V�)uÁ��X	�D�e:���W��o����f$�P�WR���hR���Bu��v��2�P��
��KF�H&ٍH�<����s�>�uڱ��*�rDo~��+��s5���.�]_�t�1�����o6�4n���������Q;��S�<�`�y��f�T��~2NO��{I�C���FNǦ�ε�^QTpA���u�Ә5�W�G|��n�@Q�}�3g�}�=��!�uĭ$%��J07Ҏx\v��D��3Y�9l{w]=2|��:��6"/`l��7���ԛ�~Y=�ӷ<�J����d밃��ٴ�;����K\�T=1�����,C��EX���1x_m��zf�!�Z'���؇��>�|�F7����g�oG]Md���4�:*h��e<�N��j����W8*M{�&o� �~lz���Jӳ`{2��;���4�j:���k���z����~y�oi��5ё��~����M��fg���^髬�M�j8��1��F3{���p�ˣ�Tz�+(y(%��n5*���:Ƕ	��$�;�u��h�or]��aT�I��u;��pG���TP��Y�j�7f-�����{&2k��=�A��L���2.��ᛖl���ǅ��������7*p@�'��Wzmϋ��Uy\"����wǈ̼k���Q[�D��ξ�U�Y]#�"M|�FE:�=:���<�YPxM����� }�2Xg��W������Bs녨P~�����w���q9ծ�L9s����@�	[V��̱� /c�m��j�ٸ��O��7�q����Xڈ���O+.s�a3�G�l�����-�Xm}�#׮���ww�=8�ǺxK�;�����Q��Gٓr�C� �G��æ���r��E��Mg��U`�\�籡�L2W;b�".s��6�E�����Q�浄��]���IJ2y�G]��ĺ沎���|^�/����N�w1z�ۨ8o
�J�u��8��ܴ�d�n��M4�����t	���ݧ&��{��N�����/Xz�����驹&�0V�+1�"6:���p��u��{���8������W�������}�pRVe~�]��V�ɸ�+�7���+���;��´!Sl�v�[�y�&�A�T���p���u�9w���N�J�g����N��'�/�J4��멺��:s\4k�GX�NE���]�D߾?{�}�����D�z�������7Q�4��̳k-����Vu	��w�SCs�G�Γ�ƌH�[�<\���{��j�oĥgu7��oH��fY���ScO�S[�0U��ӱ�L�p�`U�kk�{/N.,~˴;:�|��(t���38����t������J�$�ef/er"&�qcݗO��2;���,�W8�m����8���j\Z�����{��[%]ċ�!h��0#Q>@���$�٬��q��hI��FօT�>����=�v�!n�e�u~�7��@�r"�������Yy=<������������W��;���K�c�=�q�"%���"�۳�����]x����yK��[������	!x�%3C�����Ŕ~C�#�c}��d:�Gk�$ji�}�vPkI���>��y��=|�ofx�U��+y���y$ǲ��"ח��w�U�<n}`dEkNL��P�� �g����M%6���5��x�J�mf�ק3���U"�B���֛��KZ�ej��М�����>�o%�'�����}z��×
I��)�&�鎯$_���2|ɿ_�����������|�Z۸���U�i&�0f�t���2��F�Ŷ�If����I��-�<ƺb���1�&��˜fi���SZS�[�͈%�$��ý��=�}�����>j�#a��y�{~/�P`_=��$��[���܄!x,0��:�
/�kH'��e��k��Tt
�����\�{�ZS��;��΃�z"�W_d����*�tol�q�kDr ������9��o�S��R��?��Q��9�TM�o)t�,kSulii5M2K���wy蘻���ɩ����M>�*+��X�Q�/c�ۭ+�Lj�����Vo��o�H	�0�׫2��8̓�����C�����=�1��[����c�����?��.R�/����ztrI}�_����ӝ��徂��D��a&����g���,W����ֲ����TJ�X�k&��T�����_wp�)!�+'+�l�G�[��k׭fo�������}������v���y�8d�f^.[U���ln����L��;~g�+��u�]���HO!h,��ז���{O�и��=�1�����/��]~�&���H(;��n�z^�6�x঻�c82M.{{J\ƺ<��eq�KBCY�	e��h]+*�gi�Y�gݝ� [6����N����L��u6'i��c�gˡ��HN����s۟�.����~i�H
�9\y���+�KQx���i�tT��R
�/���!��-e�����d�B
�2�;Nǅ���N=Y�o���{��#����ѥ�m������큢���j'���tZ���; J���g���Ox}A?��e������N���ޜ���E��m�xlѺ�3-��_�n�y�
�ύ����=g�ƣ��$z{$���]5)���*�߯���w�.j�>�C��:欖��xe<�[�7�!��H�KӿV��!:9�{ʾ����</���������\�>�G\�D���}��(�ҥ���8R���Q��ͫWb(���M��L1v{{b�5I�V.�O��=sXz���2���߭�K���2�Ư�n��i��pu矻� T��ō�g�;Ɣ{c}�S�M�/�̫�۴�lB"���q2L����q�["0�4u��~�eq���A�0����3a���s�]��}�Q������a��t/^���VZ�
f��O@?��w7d��+�5nI���sr�P`,R�h%�.�uЏv�ԭ�ӣ��v����6�f�"�!m^fW
c3A�X�vӒ0w�B^�-.ju���x@Ι�n�n��2��������?�r��<��o>��em�]�W��b7I�V��Qޝ�.��Cs='6"�Q��?Y���ѵ�cNkQ!���Y�R#�"_`���9��g�J�7�ݷ�c�b�O�F
sǙ�Ϡ߻o6�/��Yѕ�5~yu9�JtiwZ�e��2��z�U0?+p�^Z� J��k�v���i�>��y1h��~���s��nakT��o���y^���zɂ��U�j�5B$7�@��pQ�Y���n\fí?�GN2��V����޷�β (�b��b�_��o$s!o>����[v`e)툯f�Pҵ�� �Hx�|cn]�\ߩ~����ݢ�=��;!�Ff�+���t���jc~����iɹ��B̠�$B���n�'���ּ�+w��&e�@��_N�oomu��E�c8}c�]yPA[�FNgNo�幐a�p���jW�l���U��ݾ�k�mlmF�K�=�}����������PU���̮�m�B��j
����ǬewEw)��Ař7{�K��U�v<�?��5Yym(�!��jRr��$�w�,���n�> V9�-Qc��]N!�Ć��{�#Vl��/mJ\Ե�C�ZS+
78��l��	=Ӡ��{���w�ԉ�!�tV��uбUy��P���� �(���s��F�Q��ڞ6V����Ѩ�ڻ�}�N^^�}4�g���NT|OU���jGwK��FO��_�N�:^�W���qK���С�Iפ���M���m�ዘ񓎏�g��P��R��=^[��{�^�9NRq����>FG��U�L��W���/�k�7sk&���Ud��H���߮��?H�ޮ/
u�����W@��r@�n�BB&b�u'"�#�]aT���C꺐N,���/�,�[�C���㿩v����!�y�yI���"�@H*$L��li��^[9F�K����A�C�^�b&az��򵏤��Ċc���Yjk��	��}�c��J���*�h�D%׻����������i�J[��̘d�9y���p+�m�X��>Ӑ�����ɮ��o#�c^�f��l��/$������4�K�3��,^�Ͻ���սyb��>�N���=�lG�y��!�kc5����c���*A:���eSN�Gm��t���^��ܗm3R�����(iU�4��$	)��zN˓�#�e�E��WVh�&�����C��+�iX�[<�c.ŷ�m��6[�d�$r���U�?��L�)%ei	�ΖV����-r����ض-�_����J�uVe#�hILCM�1iv1�]Ma���M6Tଝ�{���U7�6�����bo>����A�	d�wV���,�Y��,��7w#�y��T�^2�����'6�Y��d���{�`f���z�&@kM�,��d본�m<<T�����{����@�H����n�L�[�ֺ��V�����a̍	2$*6��
$7)8#s�����g�O����WpDo���HBcX�}�c�G��ٵ����{;
j�x�ZʃQ�ë�R>\,��� ﺩ���gGLLg2=U;�f�Ԟ	�Dg�p�^��x��0uzB7���X� ����V�v��r�6¯���>����Ff���W\:�'zgc�[^��;rv���=�ƥV�9�~���»�x�:X���k�xS˝��c��֔�_�|�Mc�1�#Pb�����A�8J�/�{��xzy�*Ƈ>�08��p%��j�+=�ϳ���s���<+(Cc�+�����Z�z{j��w$7~7���_��xa��v���&�C���չ�X�1�'8��ծ�s;���ݻ�ѼT��t̷��s<,ə�JךN����G�^U�di��p��<�.=�Z�����|n��܆tEq]����
��K���#�y�A;'�:���$�l�*9mB ���4�.�Żx�Z���{�-�r��ڕ��Ⰶ݉t��+�9d]q�*2qJ��Qf�ܡ!����f����+�p��k.W&�\�j�N],�_�U~�2�-D��ʼ���R#5<7W��+��d[���4� ;4l�F:ΒS�օu�C\�n��Moz�HQ�:��9c����VU�={����5��i뻐謝�&��I������f~yۂ���:�bw�<A��wo]�!w6e�Du��J�Tn��uj��a����6����ҳ2�β��2�R�c5�q̰5��tYD�41:u����e�bU���%p�*b��.)|��z:�~�s_vWn�F�Jq9t�&v�	�MFw���0ۣ�[c�4��Z�3?+�M�c�� r�[���kX�n�{}��5��uŤN��άv��|� w�u�T�J���^!dV;�
*�zs�&L��16�I���6����vgH0f3��W(�}o�j�����ܽ������i����Y]�JC�Z��GW���w2�s��믓����r�ns�t�5�G�-۩�{������w*	۷2�qȿgm���e-i7�.hͩJn ����,�nZ��P]f�"�Q܊g����hW9ճRv�h
3�s�F�]kpN�F�S���Lgj�������[<k:�!�Ida1��Q@�t}��(�R)$R�I#f�r������>��&$�JF�-I$���a(�\۝���n�۶�ںm���Y�\ojaE�D���z�=��u�	ȱm���˝��wQ�'����{�+Z�p_l)��#Ne��Uʚ�^�F��S*1��1����d����O�>FU��b�&�h<uvs(�8�u�v�I�6Gt��U�.!B�^ތεټړ0�욜�����YmǨ�E-W��g���$�׍Rۡ�6�-�ƒ�;r���i��x�ncJӐ�y��ޞ�w���o���K�$r1~ƿ4��$P�n��C�=Z�w���eN #�CN���L���Pn~U���Rv힬�)�+2�6B�Ir��pAO�4�с��v-� ��I�A  �P���MȻEw�����?���η�F�j������[�4�Y�ىl�6̒,�MZ;�HlyuԛZ�.�.�8���E6ٗs��ۛ�i�βi��\o���Z�%{j-�5�s%��'�����5f6!R2�*fT��7a314�%��c��ٵd�6�-�:i#u)r]h�d�6i�X����uᔒ���ޒy��md��[���V��ĺ��n�aby ���&����ud��)<s*��&SI.d�h�[s��LU��R�<��Ւ�QzFHnַd��]u���m��6��V�v��2MX� �٥ֺR)SG^�V?<-ԝ�{YE���t����$Ό�f��,��&m���	k��c%ش��&�s,�R[���%�gk�J�[�Ib�eԝ.Ý��tծ5˺ˏ�'�H��%�:��a����+;n����������y�4ه�:q�',�Ȋv���g�:6^����i!.Vs#Tw��ۮ
�6۵��<<s��u�i�f-Y7ec�[V�O�b�˷�\������ ��/��:^���D{\UeC�z�1A[ԦA\��ܭ\�(���8�g�p�:���*��n�����O����ZD���>:٩���hN�Rƫ_�������lK`�]1?o�?�n��^�O.�}nZ��@�xh�k�n}^���舆]	�ך2�O!�{�	@ɰ�|��f�i��hE���z³q�O�����#����o��:37F����ѭ�lAL{����Z��C�*�DZ��P21Gj����w��;q�%x�篽[ʾ��!�W�ju霹�v�(�s���N��6�$��ʖ2��8�ҷ��bf�=;�=�,�U.�,�����9c{@��t�Y��{�b������XQ�>�'x��M��>G���X�-f�/6��NήҶ!���KsSy��W|GUf��ըu9N�ȿE�ך"p6��I[	%�U<G7�����)���c�/�w������#��ӫ���.�+��a�;��B7��}�5����v�l�W�^S���d��x��}yɺ�g�`f��x]���]�F�:�"�[ESAD�2�f��H�ܗ��X]�����,�<j���t�oA�w�Ϲq2�4:f�(N������X���,�d�ʦ	y�+�Uf�]�q�~6z�*A� '7�(ǓXt�1y5���o*n"ꪽ��Y�w�v�C�ʧ	è/:4R�6& ��^�cA���/��"��:����h��|���Fc�[�P��F��,�����J�VqK�[*�����5p��b�hϯ���hvNm\w�v��kp���f����X�
��y�f�o�e�t��r�(A�J��o��z/ѻ�Uٸ�35U�vav>��Vl˓�vDf�/���w1C/;�\a�à|P��5�6��0}�ţ��=0�gs�8Qꎺ���y�5���_Lq��RYS����@��9UMuCP��I�q�s���锻�Ck��Z���g��O�ǻ+���]�5	{�V{!w͔�>�yz�~�5e_�Zb��9	�vΪ����]�1�::��o��7K��y�s�ZʝBQS��w~�w���*u�;�� �ل
�S����U���G�����m�Ѭ��t��դ���1}�i�����E1�1�r���dMw+�)-�,F��7�ۏ0٪����˂�X�˩W߶R�yդi���j<o8�)O�FWgwt�5_�
7(Rݖ��}>�_l8����bմ�=�K�K=��oo�{��e��i�B/�*����7��1W@fj���Pżn磎�&E��L�2�6T����E�}Z��+Ȑ
Z�|����W�VM�MV|k���o�R'�*7^-�&��Ұ�NUuW�[�����L�U��J��2���uS���}�\����Rs�~I@.=jwx�}���ݥ����vVOEV�#z�����v�'4����Ɇg�
��k���RGK#���{I�\hˏ�___��L����`�q�w�\�;��~�E�2�[/�ݛJg��e��B��7O�|����~[ae�^oQ�GGmH�nH�����R_.~�I�s<�)M���o���e;8=�ϯ������;R�ME��~��>7Ux�2}��W�����q����Ⲹm�\�*�*�;���	a!�5����b��ؼ�����\�o�^��:e�[G%ܿQ��ʫ�7���Q_%w<�h/K�.��B1���N��W\0K��Ƭv�qq���VF�]N`��a��S�l�mǮ��9��u���l8ۍ����ͨ���fj�{,u�d�Qu��t�_���A�HR-7��)�0�zx��,��e�H[�K�+6ƎI/[����'_�I�,۴�,��5!��5&��A�!L�]1�n$+#�k�&���]��"��!�Ӝ�v��.�9���5��Rp�l\���.��9&��m������2��x��gq�O'ooN�)�Ⱦ���S����WV6�Ѩ�}gu����H \����A��F�ع��>�q����9�����R������m�h�w�t��3�E1���1�P��+���bwU';+6*UМRܕ~b�o����Ud<��E�р�뚱�&�uL����Zg��j��^�vJ�pHz}��p�WĽXyǣ�����LÚ�*����'����r����nO���Mh�QDjK,��qz]�4� q+#"���Ovp��1��v+\#�BY��[({��wEL��aW&`��8bQ��{G�zn3�8�ǖ����+yS�YNO
Ws�<����v��6�{��b3]�}�+�2�j��=~�{W��������d�=hFN�ʅq��P��Y�'Îmh����4����~g=>=X��t�9�1�հ�YJ��n�O:<F������E����v(�&]�X≛�^�IŽ��6���xC��,�uh��+
��|�j9�V;j�/���o�C�0qk�K�� �^��}�נʹ��ȍ���ߋq�@�w�6�H�Wf���Ǔϟ5�'�7�fɺ��秳ﺞ�^�LlM�j�Y��!DY7O�ӔC���Y9Jr�rP���q��tR���ﱮ��r�W�0�*zc�X�s˒v�Й���{ᗱ*�r}�ۥ�0�A��9f ������uTM9p��;��F����K�ƳӢ����ܟ���m8���{=���f�39<�֚Cη:���ku1�ĝÉ�%�69�V���t�Ո��	hYt�N�mُU��Qu�(}*7n]�n�(1/��n�a�}qu��m��1[(FS�o�r�������촂F�}]���\�u�����ok=��>|����vԺ�lJ�I����C�uNEY��������5Ef�u�p�|��\�s!��H���d�T�y&|��ޗ����������Рԅ�KIl�O�
 �Q �Z��c)�s5� �a�^��}5�� ���E���ro6fV�I�k�PUȰ�J'0h�M�*��]�H��gTڕ�i~��ҹ!�L�����m
�ٺ�6���I���66�]ꗸ�ow������G]�'�yWͧ�Z�T��T�\p���@���R�`�4|x�=���l�e���qD���˼��mrs��n5�^�Q�7�}1�dy�H�%��ν�*
�u���V�F�7~Q9�
r�������V�]�2g�](O���g�-a�թ�$�ELow`�t��ȏ�� V�_���@?�؆�]�����}1�	������Ԩ1�&ou9�:�������953g�W�v���@!e�>ظ�+q�V�[3Yk�*�C>U2"7��8��T{�d莾���w���+��������������h����v��}H�@��T��\':3�.���v���/�%��<�z3�!��6-��jm&�g���i�Y�8��(�,W��`����5N������6z\�x�U�b�gHt1���PAxpڧ�3$�YX}�&$�r�>�Ӯ���F*�ݗ{Y����Gp��t���;���׻��C��ï��a(I�9f����*󰜎��dث��x<�� �E��Wm���\�ǘ�ǭtJd�aKW��uY?��Q)�D�1���@JK&�3��پ{���$Ka���j
�;r��λ����M�wʒ���ܸ�:o)9�;9��'9�3�����Ň�%%V(���鿗u�ߔ��Q�Z<��U^~�WR�w�b�b�D��&#�>_�S���Tg ��NS�gu$�o_��nF�݈�P��c�*w5���WS�k��|;0�^���`Y��A��鋙� ��;��?.JG׵�tu���}q�x�X�k!d��s2��-��yW��w��
�"�K8��.776�}��/��̀ ;�UJi%zcʆ��h��kڲ��l�BRl���
	��D	2H�H7ԧѝ��ĝ�����Cj��<>�7�� #��[n���G��+^j9<!>���Dd!��@\]�W	_IYQ����ή��n��:��;����\!>_;�����X�Wu<�6,����&��Ye��~�����{E�!g�>�%N�W�D��y�	��a���/�*�������SY7՘�`�1���{;��CX Cq����1N���3��hSc[�e_�הR�K��V%�v�6������
p{���uvJ�J@���{ �.K�M!`�.���sskhM��'����N�20��ڮ���R8�U,�4qŖ�p)�@ϬHj�z �r���X/�$$,�
��	�X�s��3HJSu�)#�4��[dem��륭����v���m.�����Ji��i��I�t�[	c��;E/R��V��{�Z{ϡ{urJ������a"���ͮ���0����=��6����&��d��L��u[��P�� o�RW�]e�|��b����G�p���-��>�#���˾	^����Oh��Խ�}��/�i����<�{���kt\�QT��,Rh\q!�0�f�m�IRN���\2�}� ^��"�΄� �T�k脲o�G��R0O���ٛ�6�<cCRBEi8��{8�ی��+�ڙ����^x�lE����d��g2��h�ig��L��N�TW��5q1��� �f�/G�Sm`��Ӎ�U�&D9�=�r�7v�0P��S�+r�lD��WMܨ�r�|�j}�@4齻�jl��.&��oX����$ұ:�p=�������?E"�T����I���3�\;3'�o)�Fa������GKU�ߣR�Ĝ��_&ߛ�[��]G��Q+����z�ۮO.�z��W}��B�s��)ǯ�5�_�s���wp�J!tE����C����;�P�����\Ό������P�}�7#�db�P��r��q]��LGF�Wo�G�<긣���}
_�a�R��y�οm�dF�?��?\4U|7�g$4W��!�`���#��5���%0Yj�Ԅ���{Ț�uX�8O{3��y��ٗMP��v�;q[���� κً��Oˆ�Կ,�w}ٙ�C����M����� g������d��Z+ў���3V�pFd���3u[z�H
ß��V�hs��$FVV�tO�2<�v8���
ONR��XXl�TF�u�
T�!���ɪ|�	/*L�;�Uz����7Y����}��Uƪ�!�t	5>�ui�۪�՝gŢy��0�uz�z�ck�+�s*�v��v ߣ���wL@8��ڔ�Lo-ۙ�Ίk�6&�^G5��ؗ��-�y~�������u_���%'Фޕ.�oA&	R'o��7(���/��<2��4�ӤP�V<Ve�U��u�v�����U[�k�3��d��� �r{����^����fz��ҝ�d8-��蓋e�dsH�X�x�4�cۦ�^�SE��E��W4V�|�]J�f>zA�F��
��4��\u����{�S�q7]������4���N^�S�r�����S������[�ˏT�>�3���M�_�(�@�ζ�G�WWr�l��f�v�1>��cC��������np��k)�o��챭�R꠶���CXF��r�|Ύ[��?�o����k)묳re�܎�BT�}��_l��Ⱦ�0��|�[��[��0z��wiKލ~�ux���u�hu�	V�I��k���ᔧ�{��ѱ��}Y��eL�-�t�R�ӗ�i�6��t��慫�a����-�L ��N�A���Z��׭5>��K�`�G�������w�"���~�^�n'_衢k&N232]-^�ݫ���l7���T�A���G/3��=Ә*A�.S�J24�jC!x�9-�r��W�uS�Q���,zbL��N���f4�Gy�r��������;[[��'�y�A�����(�n��W�]���>�6��N	�g8\9ͤ��B��y	�L�����ѵ��w��
��1�;z�O�T�����U�r���Tx����A�����c��]��~���S'�M�_jY
��u���������5�d�gn�u ��բ0�t�LI�(Z��H�v�g2fe��v�j�)�}����@v7�۫��Ɩ;�m~�6�.���Y�9^9��g
��ʅ��s�#Cw:N�����\��oaDV��-tA��6���@�ſ����=�^r#m��" �{���v��P�m�����L=���M�c�I��Z�3�m�� ���^
X˙-һʴ�C���XJ#����5G+5=S��<�8$�/&s-��F$��R��\w�9�5C����4n y��H��̻���\����+��k`�g\�O�R�w�?q�j���t;٘��i5�K-�"�h7U�ܺ6�B���2pu�G�D?!�Է7�*g�2]q���WN��3�5}��m���lt�+�f���#��&�ڷvQ3`MBNƇ/L�aߥ�^6��� ������Wv�`[���G�6RrXۓ���7��i�{N;|�[��fL���������H�y�3��&
����Tj��ݴf�VR���.�^6ʺ+5t��6�N���Ƃv�<`�U�hUuSqa3]*f���vY�5���w2���k�����2����)=X��Ac�Mr�r1U���H�Ƕ/�9��x(�/xu=�^V��d�7J˼�5f�ޔ�O��{�:#�sw/V��kt6�C�7�y�Ʀb�ZxTy��:�Oa�X�	�X]Y�*V�8�ZɻЬ�X&�@����zG��;���I;�@�Ot:	J�rV<x;$��7K<�	�-�s&e"�i�{���G��b�(ECL��������[��t�D�B�l��ǀ���޿��=�=�7�v�bX�Hs�mAל�-+��Vۡ0�J���%�n�ʳĻ]���g��j�\�0��pꌫ�L�Z�<���z�0�D�ܷ�C�!�[g�6��ZH��=�xѻQ�ў�$l�llj�yW��a�7���r��;�t�ZI��ev����r���ߍ>�s�H�w�����@�f����KUȻN�t�W[amv9i:֍��p�,�].��H��#�jh���I�L��K.ܼظ��d*�Ov��c�\٣��w����'N"=����  	�.z(�
ޏԭ�9�*�L�y�$���q=�ػ0!��3ռɖ�/6�F!�A��U͜{d)��P1F��3wދ�iD�id8��T�(�L�m=�'R�v�w{q;<���Go�Ԯ��us;��W#&F>��&��(2�1{7�A<����D¢^����i�Jߏ�?Z;}>��F3ӫt�ec�C3>��־�C��_��>o���v���]�do\�vG�#	�cK��8�	�$�rЭ���	����y�?n���o����qE��O�S+�P��.8pT�:,����di�J�ׇ����	/��9���LEF��Br�Fp�[H��q1����g�k�#���}�~qo��p+A���3-t4��)���9l�+`#��G��q^ڍd�^����0��aq,謜V�}L�x�-��0H}>���s>����G���ʢ�N��E��Hr2(iu�|��ן��Ǡ�j�y׺�:t���z\]t(��T1��Ǟpw5wu�D�[Ȼ���b������q?_1w[�M8Q�[/J�x���Ȍ����w{s�}��$��� ���m2k)���I|�ҟu�ZⰑ�tH�O�<Nv��\��ˤ�#�L�^�*N��cr2����\��'+��DN��9B��f��4oX�.T��+SbIܒ�C*�+��'zRY����t�E�g4)�r�h�`��U�^�c˳<G6��3����/��U�:6�e������Oo1�b��j�����:��K�[-&�V]JZ�֕#SW7A*,�˺ۜ�&������=Jou{�������{��[��3�򬯰C���co"���Ź��G��y��|�~ω~����{�ᇍI�]�ӯۈ'�U�Ag]'��������^�N�r�#Ҷt�Q�u�{Ӛ��&\e�]<��GnV�����`�ʋL\f�N=ܓ`,���V�홝Z�����("�FX���j8b&"���3�ؾ5�"�kJ�g�$�_�z���n���mu[��<8f��
�B����֨�sH��#ۓa�@�9��V�Q���[����=��f$v&&|�u�,v\��Wz��ER$�c��L�ғJ�G�g�
{U�ֲ�e���(Y���>��W,)� m\a��Y��d8~����9��/�^_p�7l�p�n�-��"5�=��Gn"�<��io�Ne�t�H�Y���p�:`י�{xnc��vZ�oR^�q�2(@*Q��o�on��g&��S<<v�Փ ��b�.�O�π�~Cu/��n�P��Tۘ��N=�)�����	Mzk���yR���d�_I����}]2P��U��qz����H��j�u�=��ER�T���ã+�<-�J��sJ�Y��Yˀ�4�+��U�(%����2�ݝ�q��GaF��{���H"Kl�5lT�H=���ؐ�w�{+��l4t����Ӭ������rX���?5o��}f�,~�F*#q��O9�	4�iMOً�-k>"{!\�3����eYm5��k*�>��4 �瀌���D��n5Hĝ�ɞU����-��A�RZS��*��W۝(��WP>���WB�n\`&ؼ�;!�!k��'��������`��_9uΗw�|��䧰��ǋ�����P��a2}xv�+��d�!펥�WFF�^Rޱ�!�^���|"�uέ�R�{(�$��r����U�:�i6�����Fo��:��n_ffm�=��Jƾ�;��|�2)�Mxz�X�BP���<����xy�����7 ��|hh/9y"%+��"1$�{:�e�D�/i9��s��bֈ�d]��(�C��8-e	>��CE�Ɍ\OQ@��E6G�����VǑ�nd�ON���۲�^�0��}+5���J��-Ƞ�˫V�n�c�/��?	�&�q��A�fB��)��&k>�R�W�q�s�_������F͓jBWMnw\B>�9�*6Rϡ�xޱ9���f�^�;��.j�F�Svj���4�\ίT�8�l��@+	u��E}�b�;Z��1MwE�W��j��I�9b�sj�1�t�y�L!6f�#�f�҄�ye	qn��]�!�	�����kz�_ک|9ͬ0�Wz�����Λ����B��y]��hB�lr;�b ��7��i�Vܷ���N�{dJ4z��=hBlުڙkDQ�Uv�b�r�o�r"6E�a$:]��"�}����q�Cu�f�sR{7���*�vYS�e"r!�,��I��|���G�/.<tFWs{�2��W����m.آ5M��.�e�"'�Mr�*�F1
ޖ�'!/,�cSs�S�Q}��OG��ձ;��+�Ϙ��z��s�e#����r��$%�l��6l�*,��s�����E�_Ok�����"��=ke�A&#b9�5��p�,_���Nkl�r�"��6�:x���� �/o���������Z��i�+u&7�1/u�S�3��^h�kj����_�с�A���-��I�2�o�=�n)�\IG���X��@�!��\�dISK�����m�S���0`��"iC=ט�V�����3�J��̑���T��D�cn�{I	��۝N �ᮊ�!ﳜ�w�{�f���3J�]=�ys4e�cG���Bv骩���ވ�;��F�Z���V.uyV��N���T����u^2<i�;w�n]���;��0�.1q���GK�y���K�6�D���Lvھs��b+yv��ĳ��%6^T��rþñKS��ld�q��J�����}�ґ ^X�=�$��oRF��!�sgGWd����^1Pz��$dnoo�yn����n�l���b3����_�&&�%�WyW���*�>��3z7L� ��̞q�Yϥ�f3��{�hQYX�T��o�^�{���.��0P);�}�,:� �y���v�2����ś�lLtJs�Y&�{��G�=7� �����ھ8�E�f�Ծ��)-WP�Δp�x��_1����%5��bFZ��h�}�a��?`��o��d�D=�Q��nA�� F�DS���Ϯ.i��6�i��{DЭ��F��6=��	^�T4��//L���I�SWWW�k��f�6P�iױ��7I�6�ڧ]�([��� ���r�� �
�{�����Y.^��/}����ϗ:�7��u�����C.{����r(���x@B�b���\:k�"�83��߶5���S�9������or�◶�{o�p��]%�^�W�`�V��2o��1oϵ)�:��g�����A�P��>�`�^�V�`�_(�#鎲��^�tJ;�-ص��;ª$Ѕ\��-3ٸ�͆�gh[���VUm�����FeY"Ygک՝���vѣ̣//�Z�M�2�U@u�p��n�	̫��{ab��9*͎��kH���Q�uΤʺ����B��׶�u-��������x\%#?揞w�8��qf�	q���m1���Iv���ɦ4��Q���]M�ԑ.Q'I��b�Ô�h���o�����(h� a�v�/����CP�z�D�;GlWjL����I�=c�������m��x�q�:�d��C�5U�Yߠ6S��?�czw9V~�f&�0������ �C��>+��{rv����ú��Ӫ�hq37�F7�(�h?p�p`p��.�1�JgY������I���jg����f��ں����D���R&ц6�r0��F��8�}��VyR��eD"�ǳv�,�꯼��Ny����c��U�e�$7��^(� ��qC+�دʍ���=j�R��S��WUO�%O'�	�0�
���/��*G�v�����1��j'���k(q�W�qU�\7&pD�a�>�s���t�7ǯÀ�����O�o⭽�:�9�{��b�+�U���*��d�'��oN���5���|�f�]SW�h�w�fw��ڔ�Mo���z:�^��S��;�~�6�-�{�A�bH��Q>��޿��@ö[���:\��2ݕ4 X��<����������O`Y�Vߖ=�&��q�_y`��L_:cc�cpY�(��4(`fS�7>�M�Ә|��@��|�	�=�����onG�x- `ѯ�<]z�>�S0��佖��*�d3�`V�CR��Gb�Z�;�I'�����9e��u�����~���ff�O�R�/6�Z3Epth_��6��^[�ٲ�j�xt!r���¤C�*7�F/אMS��&��53�}hi�s{�O��͏m`�(�@zY-'
�.jHb��g��>��U5�G�L,��l�B��#��R�wyA�_����Y����Y�I���u���z}2������S���6=�w)�+�|��zM螕��Ǚ�@�����޸�!��2����s�����}���ZK�f���4ifqx�n:��^�� HO �W��ꉎ�$�/��B�R����8O��0h�Fkht=TzT���>�Q�dWm�-�8�fZ�}{큱�#������y�Rxm#�W�@���u������&M�Cc&��n��L�8��w��2����lT{�5Ez���%y��^����Ds.{: �k��D8����Ą\�W�HF�t�N)���r��T�(A甩��z�f|��͝>�i[s�������4]��p���K}[����wF����m�'�86V�5P�o^C"���Q���z'����|���VJCЭ�5�D��1���v��ñ�_Y�Y�{����Y�w��f�1��u����v�������q���x��{�%���ʔ����_ ��j�ŲM}�z�W��u�,�y�����8��̴&�N� w�u����H+MRl�oM�o\�M#��u�C�ZBa:�����裔���(��3�؂z��h�E���k�ɸ����᥎��Ӣ�&�K-F�����&����g~�#�9gr�*k�t�N�H�Df4��/���O�ag5 >//
��y�U�ĝ�"0I�Y[�H{��_��z�y���9��;��,Sć�G��Wy�{�N�UfU���ٳF�[�`�%	?�쒄Du,}���
�#Ѝfmߧ�եAz�`ɼ���rRT>���#j��
r���R?h3�u74��F��j� �}r��v��ɹ�����5DU��4aTme�U�^��q�;Φ���8x�*�^�Xå�ݣ�d�?]*�ʝ�a8'J�{6��%Aљ*߸�m����'�}3ǐZ���AA�E�����~Yd��I6[�fVK\Q�f����D��R�N6�[�QN4�$�����Y�N9?/��=������t��_}{���ƽ^�ff����#I��O�Q�$.+�Ny�ȍNĤ�������7���|}%�m��b��wR�O�Թ��ȼw�zp�]�kt���sB3��n�a3Օ����= WP��c��߫G��p^h�i1��5Cą�6��ei�Jr���1�xzW45���k���s�{LQb+��V�(������ڹ��'b��M����-���.�}v�a���Y,��X�|�����y��!�z���t%�����5���2�_�bS�߸�����Yۓ�{�?j����_�1���(V��}}���|�v8W��I�ǋb+==h�<��Ǭ�U�Q~��1�U�y6�ghy�6�%ذ;�t�]�����B���z`mI�����͕��|���G�.�FD�
��j���/&���\�7��x��-Wj�y�mPo��^Q�����iL#�_h��+���P�^�CL��	�,{k��JFШ��	z�
�MJ%]匬I�I��R[�X%�a
2��Ί�h�/���'�if7�"o�����=�(�j������Wif} ����ې�s�jQ;Ȳ)��N郞U�0��LO��ν���^�5n��VO�N�;�P=3wٝ;g�^�]F�dw���藘��Q��)�.�F�ʤ��͕5ꄣ�u��M}�C��7�A֮�NQ��R�3X�����#)(�B��`��'+��7���7���]��ʞ'Uytʺ������.ō�]{*%AҲ�#���V^��u����;�P�M��qҜ#�AR�O��r�ɶB���l���Q�j[l�w��{�j��ݠ"NҚܖe&U˥u"L��	Y���P'H;��Gwkwt�ދ9o������Z#� .��ws�U�6����8y�[b�O�Ѷm�ƍ�R��=�f��Wlef�Qq�.nt���$zKi#1�.<X��E(���6K��MX״�M[	sA�m�j�v�́�	m"#a(aM-�x�]y��Lν��_j4U�G�PΜjׂ�!��ti�#MU|�*��Q������ �'M����0����sY>���>�}(���X�^���1?4�QWMߕwh5؝�}D9���һ��}�E�8&���	CD�'�]�"��Q@����B��}��m8��MEX0$~�3M�83ț	e����\"\&K`��O�Fu��R'�ί��I������=��^#�Vc�Qv<��+�#�1�k�]H(�L���a�S���&����s������(� �ka��o��1�F�^Fi�F�9εlK���왁�裧�2s\(�z��1m�V
��]<}���gf���lu|�}93�t^{Lyv������f=�qT�	����8���a��x��[�/Q�}����#���:�ꇮ#�H����.��y���f<W���O�8���B	�3k9��!�X�j�}�"��N����a�W7wz�z�%Sz�c�f�WM5y��dN�K�"����R�]���5�<$c�Ӫ�IoL��3�>�f-1�Z�䲷���
��Z����א��:7��!��DII>}ƻ;y6:\�����$��	^��l�9y&���d�\)5t��k(�!��w����*o�^\����%�e���Q���6-h�g��i�3z�{<z�c3�WP�7�E$bat�;]ע���PY�͐�e��p'�\���-u��t� �Vfe�[W�P��3o��F�A��x�])���v�ӨMJƎWb6e����Ю��v_tV�,h��,��0M��bW�o2`{b.�DW�i�ll!�9����x�:�Us�w�#F��3����\9���v>�f��H��w�֑i�N�Ӣ��f�}��{��nr�8l=ffl��eb��	�b[�+a̮}�t����3���5z:E�kN��6����p��ݗ���8�K�wTG���Ƅ�/�w�H���a{|ucf��8ŗO�X����pRދ/,��C�)U��$��Pڡ��T6��w;�鶆�9���V������r�i��eh��"t��V;Bft�1�IĹ�V��ஊ�����ի�[Z�`�=���7�m..�T¾��/��d��Z��q�ה��],����-S�B�kw�x-*_vIM]�%���b���77��.��;�1�fZ�r����,v���u���
�#\��������J)̔��ѹ��	*�l���� �����Ab�2����k�]`3�LA�tv�*_�^eZ�]&J�!�8��R������j�xw���I�������h�zJ��e�ij�gw�\��j!SYaӮ�
ea��u
������Y���ι$�t��m��X�� L�!m5�I?I#E�$�I#hB[�H�r%a��5�U�V�Z3��;ˡˡ����7`�*;3Z	p�1d9�ǀ�^b�.0��گ{t~��b��e��qǲC�` Z3C��U��2w1l���}ۃ6�t4��V]�j隹�1ur�EL�ӝ4Х��У������L~7L˶�d��I���!���T�����6H�ʌ�箠�v�E��h=�c@���{�a��A�y8�?'��U������:��0��T��u�(0��v�ɘ��M�
�pg�+U:�I+��5���,���M���MwO��j
�L��(ԪL�Oc	��U*�B�2���B	7���.�S�EI��d�a!ҡe8H�iU& (��&�n���uo��{ �:���>bs��;E��.k}����Zel���>D�n���$��
.Yi��5ѝ2���M�K�{6>ۧ�E�H�!��������"�ɝ/G&O�gK.��G&��k���%,�6J�K&ƌv�is���k�cMm'9ܭ��K�!�����\��HfZޮ֨��-���������a�W���[�m����B$��n�`z٧�g�f<�d�Ռߖi��mFv%�Vg��|�񤸻-��,K�jF3J�1nZ�l2�5�(��m�IsU͸�͑s:�,\�	Kum�CCM��������=/I��i LX�%F[s�4,��$�i��L��˩S9�8nlA����*�ƺֱ�͗Y�c�v�1�4wiMYRM�ݝ]m�jLC&��QT��z]���%C��h#�`�ȫ��z��Ǹ��x��-���x�s�	�٤r����6Z�!��F�k�2��KH��F��q��Xpf."[��.-�{9�F�l�ݔ�Z�3��i�x#���_�T|���Q�q�,[Q�5k��(���(2��ʟ�*��r�(��zG���ru:��K��צzݷ<�<jO��� iB��;���u˘��e�eq�̎��݇�*O�:�wE�ʍ%���%�FDR;���w���Vk���8��2F��y(�4\=��w$]���x�'͖b� ����fb)A�\�g3���g�Pϻ�\9���&���� J׼�T��û���N)~|r\�*���1�lԼލ��
��T��A���Z���u�Q�5�{�C��G���`��ָ׾]M��A�+r�3�������Vڻ�+��!�R�5^Q�?>�MJo�9n�8��!슧N��P�s��b�9]��d@V㺰x�.c�}/v�/�&tՒ�H}�<�Ǽt���VW��^�n�DV��P�ިT�-Ѵ@]C�j��=��LB��;܊$b��<)F�
�s��U�r:�D���R�w���Ҏ�>�;��溛�#Y\  �W�R��܀�����.*�j�z�I����x��ߎmX�Ѻ���m'�����"{�/W�0�87�\��rb5�W�H�Ԑ��\�E�/�+t6<�΢T6��R8Y17"!�FH�e��f�����J�f��ڙu���]��
��M�wW�|��و�^S����ې�m�,X�饁䦎H&p�*��ҍ��W��� ����YHc�2���R==���sm[��{C����,�-���<JXT�4Z�+��-�f�ٶ�����%��׾$�D�+y��*W���{�ܣ�cI��
��)��7""�l/
�`Fþ��g���>���""�g'�"yD��d*�ǌa;A1�&����'��F%������Y՞�6��>*j%����������̦u��U�g"A�5���p��Ɍ P���
Ʋ�gfo����A��6c�I�h^0^������=�٤�^��^\W���a>}s� jYO�3��+�M�������S��yt<�+r�᛾��L�c���6���J#�-�n=J���1{����0�^DmӍ��b_Ds���\a����,�L�TKq'�\i�3uj"����������X�Y�.
*�߽�*���?}O2���1	��B`>�����V��SW�q���G��6UI��g�+���T�J��>�q�,�?43ZIU�UIRBa,�"FLE�`	Hi�/���e��7�ϥW�k�F���������Z3T=�-�ɚ�5��}�Y��'j@�۹���v�6�g���N�/�H�.�Vt�n��ݡ�\�ٟ(=eo�A�Pz�|���r�nvNE��󨺗�*䏺P�i��ъ��f����8�ˏ\rQIC�^Ph^u߂�&�~��_x("Z�`$��Z��]�)�T�fm�7Ӯ�kY������\����V�*cyv���iR�q�������B7����oi�&oS;�I�b4{[�r�p@h	���{nI�0Ĝ�/�噚�yE�#�����%�������_?zE���fvP���#{=>�E�Y9ўu]���υ�WLv�	 vazCee��P���j<}^��Cq7�v����蹗�s�{��YC�T1�I���c�؞��"�[v�꬯�>���y^�����w�φҎ�ǳ��s�';����G������%r�]���=vC�8B��ry�df���x�cq:���.��E����}��@O�Ș:G�|����TSN�wx����'�m:W�ɹ~�w$�.8�*�|0������1˾��B���A��0�E�)�#�D��3p����B ��d�r����b?+��i���ˌ��x;�E"��jr���l���C<HY������7>6�8��ˈ&�f��E]�P��.��Wbs��4OV(�c������u�We˽�3�3GMvqX�Yd�_P���yȟ�e����jGi��|��n��zf�[��爿�������
_�㚱�j�Ϡ�SFz
o�'�����|�>���l�³V���m�!Е*�}�.�V��}���Xl���l�GlY�Tl|����"?��=��zǤ��#�n�ÓC���dg�h�4a���*��ڤ���vY�j�k��Eh���v��m�-����#7t�f��K7���C �wU��N��F��$	���´�Խf
�Հ���DUF۱9��MM��yv�����3�y���Mm���5�CgZ�fz̴Iu�nK�칛�VR]-)��R�h1�ĕ��~����o.����VY5*D�	�1*̙�(�r�`�g^W>Gmv�v�Q�����P� ��_j|�Ô$]z�|ǻP{v2Gb�:t��޸>�@@ʏEFo�Fr-������J	�S�=�-�܌K�a���v(SL�"����xo�ص���� �8w�_�y����'����&-P���I�_	.����Ď�y)��m<Y��B�R��Vud�O�3�ř�-0�&�M'!H�,�,��&�`��gȊ�U3��Q��KΜ�&{�ǤqҸ�ڌ��Kږ���ӝ�+��3f�� \�I��|ØoXsf$��H__���������7��6�D��r���mxp�nr�'u�yDz��o!DwxR�]������+���K��p���?��DD\���6=R(#��ޚ��[�ă����1�§ڴ�(���`��<������m���ٵw�G�V,@ԙ���\�.�����:T��"���I�����9�fsL�4S�oB�C�|z��p?m��#����.�~��Ǟ�#>UA]�"�q�8��=�� �R=$�N/u{��A3�Q��p[� ��*#�
e�^�\��G����v��?;�>Rf�&t��0N�P���9(��yW���m�K����Ǵ��!n�:B7M�bc�ٳqhY�ޑ���ď}�!_`}u������^�7vYje� �u�u�٠	2���Y�-PQ�fV�1��Nd���B�,�vRYC1��۾��χ}e�_��rY�˱J�d7���V�ٮ��J������@9x��Ւi~�و���{�a�2�~�-�"� �a�XA�M&��Я͢��j�_G%�)UO�i��UH
{�>ZS�=�zz�kLͬK��a*����}��5��{|J�դq��ܡ$��������cۦ8J���y{,����v>-�����$�w5=}��5t��y�]\-C��ol�T���pQ8�{�������r�2��%˓�g�	/�ݻ�'��b;��ﴤ�����ψ�.�m>#ם����SV��~�ۈ�sww�$r��S�8�l\��#v��Gdr�X������v�g��@�JQ���V�s�y��1�x�ny/1]�P�p�a���9P䞌�
�baļ��ѐj�K��:����ĺ�$^��ЂK�h!� ���y�㰃���X�藍�x������#G�~>ލ��B�Y�j�B1]�O�=x��V�9���![�.�@�E��/�Ǫ��l	�\�Q���}�
2�	�֒���>��)g�)E�{�#zgɷ���dU�h�\M�����@IB@�����w^1�:^�}�?d�|(��[�PPޯ7B�I�o0�Q:�Wi �61;w*{�����ݵ���!\�[��\�ӊ��t��,)�C�W�؉��!�U��ov ���aXf�M�̽K��ۛv;'s-�k�]g_��g/2����u\�
rQ;Αљwq�2����N}�p���u6��ںǦ�m4���'���g�a-�[~���W�EN�l�.j�-�Md%5KJF h�k��eֵ��m���y=�eT/F}>��{���1	T�ƶL-���!�m(�/���^���Õy7[����Z����x P>��`z/�ifޜ��7G���������9�����^.0��hs��Η�yy�C�}�.S'�~�������m��)з;z��v�dF\N���Ʊ��}U޴�WTS��ϤPM�emJ|W^Q+�u�w��^�|=3��5hNx]����ǞB�G4��):��иwN�U�jy���T_d��O{)
��a<F&[�w,�7ϞY�k�ᴃ�^2�ؕ��b��!oa�6��T��ڶ�Q_a���D]G�^�A=
� ��L���2���+r����Ͱ�_�m`Vs�}$�.���YL�٤?}���C�pb<�. �{�^�c�P�@���.�g�Mf?�����[�|4���{�7=�K/��8^Fk���[Y�i��0K	{,����r�@븮�+IW�NKٵ��3T��]����q{G}�Z��f���D��Z�ՋMuI�I0��A���oG��^���h__0���K�v$���򲀳!��{H�e�`�屡&.̳��}t�i�3���)ݫ��ιL�YRRT&�$�T`P0+ޮ�1�h����]C������E��df�ܣ�s'U9k�:T���2nsw$��:����^���y�V&MBg�����'�yC��=���_p5��Si#�u=nJ�<�#u�����jv�R��AD��L����P`��Y�;�ىs�����;��n�d�S�u]\NG���Y�.&�,��x9��f�#��Q��#	ނ��fm��x'�z|o���U��w�C�nT�Fy ���R���
��I-�Bx�qz'ҧ�h���=��<��Su;}/m�uT{ޮ�R��ߑާ�/
9��"���F���\l>�&��B�#^ࣆMl{��>hJ�������"�"����	����E�1�{��#6c;��,;mq���Զ=*���ۤ�<=&s�,�Ԇ���{�mb%�NΈ�*Uh��������xL,7
,�ysdG�rWC���)�X�}�Y=��eI��%�q��>e<����tv�M8~��4:�B�L��u�~�T̅e���N�{Б빢����<[�/	��(���/�{+0��y:�� �:�}���7��=O�]�[p�[�_����0�.֫c�vnj�w�[�6ܶ�K�;3u��������ߵ��ܜdt�$j�%}��lm#l�����&2��T��W7u� �e�����!�K����<s���&��6�#�q���bbƽw��ν'so�=�ff��8�n&�[��f�k��L*X�ʝUP����m� ˾r���y�:���꟱�������!\4�9ҕ��l�&��2�F�[*�]�	5�����XCk��Xel�[i����.��/���V���v�X�$�9��J�&��.k�#���Q56�����0�6+.Qr�^^=�V����v���EE*֚��Jaݫ������*~xH^�oIU�M�����/��}u�����c(,��yd��b��7uy5;��|5B��m(���� U�6���]�|w�!ϱ*�iq1]�S$<^H!��kۍ��$e�M|�3;��{3g� [.�Dgw�����-Fɦ'��ͬ�����Mln�~8�xy�yZ�:{�;F������\�h~K��b�E��jX�[:��r�<�w��1<9��˻���x1y��>�~>����tD7N��r�F" l����O������QǵK��z�&e�U�q##2$r��r��F���d�B��+��P��Z;�Ӂ�{��8�vS���7�R|�K7���ݔa�C�Y�_](��֕?��W[*7w�5h/K��|Q�<k>/�ޥ�U�r�o�lbyy�
bS�z�ek�Ng�>��lK��q�,\G�{�eK3XsԼB螭T[�˫�sR�U_wʘ;�:��\�Y<r��
5s>������z��G���"�NE���Vȁ��{;3�u���z#�J���_V��-e.c��嫼?��|�WxL:�&�{Яr4�T�`�ވ��~�Ő�hF�4ܕ�j�:h*�@4�6:w���o9�|��\O5��Q��0���3�q�+6mXUM��.��:�M�	���ovI���x���d2dVA��-Ν^�Pv71����v�LO�wdٷ�qb}�]n��$�{��pNX�֝�r���{ò)ů��U�n�����/ɵ��R�ZAy(/twB�Û(�4�mL�`��0�����f�����5��]�������9����lD�����0�^���f�+��D�$���z�u��5X_��?���ݘ��Hc#v\��	�-�FN�:����O ��b>�9[�Apn]j.�#����o�����ΣӃ��"2���'��7���&�OT��.=,@LnI���>�:,ǂ��*,�K����Y�}&�KT2�l���5=��
P��K��X��o��ߔ=�h��o�����J\���wNv���&���q<�V�nfs4�Eu{�J�om������ �HY�n	ʲ(�0~yޤiA�w�������j����l���r�7�%�:�Ŏ��|�B�z_�>�k����C�Bt���E�:�3Yg��<˱��J���6�3Ŭ�_l�~����14�`l��ak�$n���K�d��7�srRx%��r$�'�4Q�\?%^�k�bNo�Sl��6j�̙��W�EL֨��i�}{ǪM�}�/G��x��7/��ʴ\���pq�lbr�y��{�N⺬��.�V �����Cu��k���fU��,����gn��ך��Y��\�cu<{P��M�LQ�\^"��� u��G�;2�E�+����
;��^k�3*M��9R��D������c[�~�tK���,M�|i��=�~eK� ~�G$���ez2�L�3��Y�\��MU%�XL!r� ��NF���ͥ���)�Y����q}
�g��tΏ��gա<�ȁU�'�j�_L/JF���j�QS'8N�Ȥz�qS{aW	<h�UU�Q��F��E�|�Dp����O����lw���nbn�ty�Ӛ������ϪM0P��|��h��(�[�{�횑�}>R��|t�&(n������ϻ5,���yq�9AH���׵�Okz� �]+�7]�S|�"�g��n㓋��N,��Uu�xh;��[X���H��m۰����I䒼�dX��;��Ԓ�G!�V���N�eз�;8>T^G��fi�Q]�߆��oj�ͱ�@�w�LE���F�
��>|���+�О��Q��B�� �r:\i	�{fQ� ^��ߖ՟fg�������n�����Bi,ʴ��	f��&�xg�����������
���P$�f�����S;-Et¡wWMnʯ-� a�[Ir<���fTqM�gP���oa����U@�~�L��٧]��8�X�ٹo�(�.�}~1�qb}[�dSC�O-���]�^��X����t�PPhL8���ᱢ��N��U�_�k	\;��3:j�؊�����~�%*/�J��ވ������漣����T�X*��}tDi�U�QY�$BKኪJ۟����"C$D���ڻ���D�_�������y_/���k��|�_No�si��������^w�\�4k��sp|�>WT:�1%7���4C�JH��!VEO̻ݢ�S!jMS���7F� �p-���I؞�-*��N�b�Y֐��FB�Z	�M�?�Sgh�Q�K�o�R�̷�-`"mn��b����u���Z6<�N�F�;����
�Yu�m�x��J��
bYvf�ƍ�H�^�;gU\�����T�P�e�Mʴ�<�o�j�U�}����l�[{�f2��O:r`tos2��T�r2�*��Ɍ^��*<o0\�6��9�J2�����y��N���W.`kee���)�)�J1����㗗��֞^�Ж��sm����l�A�e�D���e��nFM3 ��]D5�m��j�e��Y�Р�dB��a8P�d�S�Yֆ:�2�hR�1��Դ#��h[�$� \Z��
k$،�%�2��eۖV=M�e��k-m;�IKm:j��Y�;����%'1L��կn��ڥ1ɗ.-_���'P�كC4企Qz
U�Y�el���ݢEشkw�g	�u�YF��)X/�,������%�c.wc���t�!]{V��X��#��6Gj�eڻݧ;�c���RØ�hb�4�޹�Uf�Tu�*����%[�Iڔm��� �Y�Ջ��!�mM5�D���g$9��U�'lU��*6��4��7�MP Ք����t�]�-��H��*�X�D�(�b�B�Ь��WG3m�n�bYgMչ[x��:�;tp`D�����é�"�l�x)QM�(�led�j�е,��sq�6���TN�$��4�����^���3M��!���ɱ�~�
ôb�mּNXw�.��{��Ԇ��h��M����a�l��e��Rk-mby6�p�X���9.��v�nz�3�mz׮5�=��D&
�L��H*�A�E0��/�UU���(VH�J��V*�$YRd����|?(�����>�B$?|�z���o�!�k�"C�D���!Ϻ�XD�{O������nu���!ߴ"C�W��m��$>Љ+ϫ_��/n5�Hko���Ow�^�;M1!Ǘ��1AY&SY�Qd�ـpP��3'� bA>��� T� �(4    4@P A� @    � @
 �@P� H>  � ��                        @     2�W/=�Ҙ�x �s^�=I�A^wr��lt�;�z �y��A�+ݼ�齴���wo6��Jh������ڏ=���V��A�B����@��a��v��{6�   *�   t  B��:� P݃q�h� ���U�<�Оüt�x��z�=�����6�8���5����@i�Ӟwu�vP� �%���m���
�gg^�P�^]� ��  颼�͊�p��׷���/j�y=:��y�
I"�s����޻����޼׽`�I��q��v@�����+���^oz�����o.G@� �$� :     �ޔ5�W;�U�{]������ �f������������z=��I+zΗ�eM���Np ��m�5/lUV6{��*=�Z�eRJ�{�
�@ mR����
�� 81�Ҋ��g!�(�w7\��)sNZ@o{�J%�2�T��޷EP�y��h����
���LF^ .!��*NT  � =  �  ��s��%�s�=m<��b5Ar��G� ;�wwU�N{�)z`^gJP#����E*q�u;nl�#��m�;��^���z4�28 (  6���㇠;Ԧf�@��{t){dO{�сJ�t��T�i%q�:/v�*��`����3k��fW6T�V����Ѡǀ�s:P)xh   �� (   G���@'u��5D�� ��iJ�����R�k��(Y�� P\�W�B���J� vB��WFanY]h��G[KNN� � �uJq�tW�tP
y��gE(+��y���7����m��tH�xC�DͯCA%�݀�%-r�&����[a$�ZJu�8��E��g����  � � � ']��m=�������wZ4�^lD/6$$���Ȫ���� .ὺ����l퉯 3���j��w�+�$�wP=V�"�&��� ����R�b��t��8j������ T� )P  "���IJU�  a�`L4d�'�U �P  � MU"4 h i�P�IT�  f��?�������n�~�Zw0�˟��*�C�%����:�ns���/���vm��C�rY��1fc]��Y��1fdKbX�f/�K31f,��D�3b���K31f,�1b�K������8���3�DzC,��!���C4�c�9��6�36œx�3-Vd������j�����5�c�g2I2I�2��q+��ߦY�)����y���PI��r�7�eǻc-6uT'L��uu�R]9���G�&�iC&m�j�C�*��HwB[�M��lnc�Xl y(KSVb;6 `̊�$5��7k�P̈7H�m�M�n��= ���V�26.��[�Av��We�uw������Aހ�Ȑ���	�h2-N佭�eF�ٍ�"�h����X$XLB�F�LpV��ô�����v(n'{1Y����ɬ+RmAGK���	u�-0{�zAM;KVA�]<wzcr�#��$4�,�ଵ�K���j�Շlѻ/(l�R�go(j����^:� 5�0�K/��I�- ��y�&�ų�[�ݐƅ7Y�X�i��`S�{j�m㡪�؂���4��n�+�p�Y��7t@aw�E���CQ�W�hb"�!�%�n鼕B]
�S'3/!�3-T�wbX��_D�w�`�ڻ�x�>��6�V �#t��r����hS�+*:6
ּtD�MBq=��V���� 5K*:Ѣ�VV��"����;�J��/6!zs@��Ӈ2TT	J�ۃ.��.(\YbD��dU�1�2�p�B�i
�3) ����3o��B�Z���r���$��jd�ܷZͼ��t%��`�`S%&F��7v@����qCb�Ī��L�1�ob��XS�ε�a�ہ���(�F��.h��շtg���:���yll��b�wZ���]��0Иq��v����~�N��$�������0�њm�̛�Fő	e-�nc��ރ�t�� �e'jA�&'��[�iZ��i��P�6�0ĭZkf�g��JT�X�����b�N��2�Em�@�d
�&���O�R�Z��,��Q�EdzQ�lfA��$B�3��(l6"!�Q��ōG��{��{Smj��{;�թ�g6�X�E�q�c��\*��4�?#��|�W�d13�r<Z���4+���]�2��/�+{T�{�m��RT�ຸ�Q�c��"��r���N�Rl�m��ّ��C+]���l;��X���@SūV<4�ݽ���E0Z�)hO2'.]�{ע�L������6t��3{���"l�k!��w���F*KA��44�]��h��}�J5p�iv�j���n#���[#
�SVک��!j[������O)lv&\��ǫ��u3V_�*)���%8����7z5<B���.=B�B�b�JS�+�����b	
�5S��S��6�)�zތl[xp��D�>�:��6�z(��[��K["���l�뿓�UU	CĮ�F��8^b3t>Ƙ�slVC33lVIG.�n��2�K�f���؅��q����Wynm�/	-�{��щ��X�����e���h9@�)�Aj�թ^���X�e�EJμ�^�ĖB�}{Ib�
�����!$sZ��s\ĸ,љ�b��kT���|Y���*f��޶P�$��l= e��q2%�l�ř���H՚ܚ��Y�.�Jj((�A�VИj�R��	{��7�j̲s4R��kld{���bKU]�1��Y7���b˼�H��R�}XB���#�����a� D#U��W@�,)V���/a5>����S/w2�p��Osp�a׏a.�b�|�@��֝��^1-%���,��T��t�U.�&�	�V1
6�ۡJ��7x3L�� Ϥ�Y��³�/P�e�I*�P٬��׏�j:�v��:�U5g�����"�}pf;��u���A��j�c�^M;cd�t�T� �U�ɷCDv��e੍fmU�k�#B˵z����<��,7WyL\�N�V�a?��Z����
ݢc{.�f�܃*9.:�J���@���Iܨ�x�n[��� 扒�m�wGw��E&r�GZ�j�̷B���e�h�i�Š�� ��ti	���eh��.�_�|A�Xa��6�cw����j�o �l����&:�w��r ���X�����4����#ќ)n&VY���M�i+P���͖ ڏ�RR���;��jB*�"E	l�S@�[iiv��:V�����z�Q�<���ݕ��[n�0��;�H� L�sd8�kwS#�ZD�Bx���wNĄ��Ʃ��2��llr�W���tE%&�elh���,-�LR�5��ט�7�r��Ԗ�&Ĺ�Ŷ� ��Mm�/���f�ͭ�4ٚN�C˄"^#)�M1s.P/�[����Sr�4n�B�[�ۘb̗&C���IXyHVj{���1� Ä�.�ٰ��5q�́����'�mb�YV���+>$ �E=QM���`^���2jP�hY��t
[��5�JH�{X�5G`	D�mEw��8v]-��A�/^�(<�b�1� �GM�����l�Xs ֭{V��7�[��0Mz/0���B�6ޗ,�w���Ẽ���eK�X,Ґ�G,L�6����h�ecݣp��-ԗ��*HV��ͺn�7X��h��t��$����S5�y�o�71�{6��ݔћC4]�aE��i��4#�NKy�U��Fj�KIP�f����b��Ukj�5����BK���U����3]���1�J�Ňu�����#�懐R/8�W3�X�i76��-J͔E���"(˔�V�Z�����&@�ܫ��w6�4�Q �� (  ����H�v>���[�������J����SDM��R�4m�)	��7���s.��^�ҧ,�v�ˮ�k�q<��uu��5"��Rc�ks��G���#͐��z& 9���r>r6E49恖	�[��p� �ܕ�6���[*�XV7s)s��F�R�{��DяC��$m�v�g/�T"('6���ځ��x�Aa�M�V�0ړ)Fl��"E$b*%�R0��Ov�qԒ���&n�n�ט6<7v����E��2�O�!vj�l�9D�;���[H���PVՍ�zM��D��%u6��4��
+�4:�Dm�%#mj�#��+=ۘ�@�i]qb�oZﮠ�x���WyV+ ���OV,��T�Q:򔔶��%5� �yD�bfm�G���c�t��8��ͦF�n�4�E�F�.�S�&��gUt�v�30zə�rG6	�2�={�%��#��3yGT�U���RW�wl��?eX��;;���*�Y{[�6���	�{5mԻ�YwB�1��㺗�!��i�΃�С�$,��rɸ�^�L�n�2�K�n��ԀR�-F]]�S���*uwpE���^<EY��-Pf=�u�[��x�r�ј��g#��ZŢ��ƪ�h*N���%���v�&X��+�]+92�]g���	V5�jÕ��"�{,j���jΗF���xt	/~9�-��fK�ݢ���
Z)��7��(+R���"nR��+(f�鬄`��)I, n��%��p4){*�qR��T�%�1[7��Y1$ipS�{�Mb��&vh,��+,�J�\�5��:�NS�z�b:$`qᎁ���kv�U�.ѻ6,�l0�-�h�9Q#��a9R+�r�o,j�Z�9wV�c���`S&܌��J5u[{u��Q�Ӹ�"�M\�/e�z�fbʄ�u3rM��nV]f�ߧ��ꭏ0R��cU�),�N�\7PeX�#�P4u�ʩE][v/-*����Y��ۺ���1$ܭ$�wj݉f -��ʵQ��4����%⹍�+/ .֩+S�I?�(��a�B��aJb�t��V�˨���uz��5H�.}�^:M�[��r-���P���e�l"���$�
����sAxu�c�Ʌ����"�Zt��w��?��H���+� .���%f�z�d�R����p��l:ݦ�cJ�x%Z �rd#F�Y+P��Ԓ���W�iX�'	N͖�k�9SuN�L�u���0h�\����V%����a�S6��أ��u]�KȎ��A'�k��Z� �G��"Yx��b�cmL���km۫��b�nʏa�r�Q��Q[R�F��E�F�j��v)--'��h�b��ja^]�,l�Le�4sFR�B�N�X�wZj�Ġ;�e5�lQ+kq��CR�ۚ/F�&û�B���Tܭqnc��T���۬tV��b^�#Z��r��5kq��e���QQ���� �mf�-A��X��/
��^���1���-��3q��^�ܖE֓w.ȩS�e`���㙁��q[�`<�����{7^l�n�FP��ͷe��E�ʂ����޻��ձl,�g�Q��YrmЭţ)��M�O�5x��#M�ֳne˛v$n��ͬ��D�͊����L4K�����M�%K3Uk�Yl�/2Z��3��^lf�V���	�;����DG�!{.�ъ��E���[6]d�f��_��+�F^ .�d5aF}&^�k�{��xs֮�a��Nk�i^Bi����c*�ٺ_7a͵Jd3+mk4m��X���T��Re�;�P���]���죶&e؆XW41���;Ze�(����5�ڈ��D	MՔ�W`Y�R�:�h(ɧp�V�Y�3.�\KXs�ڼNV�!�$b�&l���K�$�汚f�[u��7^��67+�j��F��A�3߱<[�����nJɰn��7�*X����Hd�[5@ D-4
He̻��]��I���^��n'weTo$[ں��I�xnŤAT�EZ�@�!v܆˭������X(	,��ݠu�ٮ�o7PƳ2�̢�պ&A��Y�ySg���	"^Z-���tm��,�P:���3W&ĶD9y����-�Jܨ��80e`Y*�R�=>�(�u.�5fbۑ���W�Q[�b
ɖ�h6N�X���pL8Sïh��,2X��Z�>�Lh�h��d�M �b�nd�j���/�ګ��u���yyXEq���N5��h[ge��U���b�o7�13;Q62�I�esh�/o36�쫘jʱ�d(f�&��݅ �i���Z�\�(ܨ�Pb]��E͕�Z��÷��YR�f��L��r
��/��'�k0LtFfS����\{F�F���FPh.�1�)�ٗa5գ��:F�f(�	x*�L-K�i�U�k��2�/,���/t"�o���#�wFu�V���f�wy�eg�=w�bLW�V�&)WPn$`%�R�e�"���P�,,���r^6�3#�x�nl�[)�r�S� �pW��2��b@�`7����J�*�0$[�)˃2&~�p$Y���]i�_U��	���_k�y
���ЖfD�f�G�t�.�Tri�ı��L�6�WO}肸����
w��!@?��yK�A��u�71K�N`ͤ��ɶ]� M[d/Œ��ݢe�	�n[�F��4����<��<��R�c�[���{38����r�+����F���0��p�������Ί4ܭ;�]��1�z�Vk��ouQ�R��F��M���c^M���
���RR�ܚ�0`����X�8�V����K["�"Ɋ����U����̣P�L�Ee���cu�r�W�L{i�R���/^7WY�Fk-P/U�Nn��6i�Rf^j.�MY��P,���y�.�C�`%U��*�y��ⶽ&�{�>ԝ`W�g�
yMSt\������2�AVe��&�[���r�摬D�����u�to��f���f)�T���չ�겞�PAv�
�0%އiJ��۩{/qQ��+Řh��$œ\��͛X�]��AJ�ܔv���.E�LYC17��>�H��nml��F<7�y��n�PZ����Ɲ˶
Xʩz셥�ŜX&nU��t�t�D�$�sxۚ�N&�M��%�\5P�w0u�Az*VB�m�ɇ�8�F�˳Nvc̼B�AX����y5Ɏ^:�u���H�h��f�Wi�A�m'�ƍT�l����Ӣu��=����Zeئ��x8~́!�B[�쬚��y�.c�r���(f�^nm�5`�?Y�I�>�h�l��F�Ŷ^S�;�H����:����Օ�r���h�(Gw\�׎�nΰ��F��$�km�;_I �\�4l5�p��7v$^�	�]jF�5L�o+���t��Rk��%Ae^li,����cenӕ�֜����� �jnV���Zj`��.��0A.�1n�Z�%��2����P�>n�n���J���p6���u]�����ܸ�N���q^*�yXo㈚ѯ�`B���AD��u���jQ�p L:kn��]��
�5���/V��5GM1r١6܅*,r�"C����;��o^�x!��@LT#t�Ҧ���0bב�㣐�"�3ncP�+R8ԧ�eI��t���iE�So�,VVJ��2�kZy`ۼa"�5t7��7VT�����^;XU�	�
�d�R�Ԙ��=`֫�&�b[0��a�r�m��;��^0���t�/2��EZ�3���T��
y�bX`��N]m��U����Ge�����a�� m��ַk)��n����d"p�kW-�*�n��Y�ŷ����X��lo���t�jZ��O@v+2�X���2�Ztl:�3S�oV�[mb�7��i��ښ[�k��3nZDc�����擶C�ݵ%�S�#��2����M5ɱl7QrN]�lUbr��m�kHH�����2�XcO�f�D[��ք�wO���� KeH轋���h��tw	�Y�*��q�H�r�%)[F%�4U�ۇ6��Q`P�'
˵X�����ʔ��`s5UU@UUUUmI�	U�UUR�UUUUUZ�h��U�����n��e[(�pR��UUUUUUU]UUUPUUT�J�*�U Y25UUUUUUJ�][J�*�*��UUv���%V��6������j���`�mR��sc�����v��V��[�����V�]�]�7N�9�R����r���hqv*q��	P�;�3�۞�qg�n����v�r�5�'���ӎ���4Xŕ53&� Jt��Wf7<bH�s��鱉5�]�h���L��P
�D8&��*�D�z��um����;:�'=-,M�F���C��5(�s�r�)q�c^^؋���ג;���f� �T�������h�s�Ny�c^��֭��r���uU��n0V�9�lvz�som�fC;��u�۫�<psƞ;�9�p%Ɍ���yK8�]�۝i�����9��6��R������,v�����NĆk��nOR��M+�Y��aB��mەˎ`��zz������� �6֬�Y�;�bn��<-��[ݎ;vݵ��i����n�ݕ��ø��b��Lr����u���tE������nZՠ�xc���3�����)cp�������/b���w�[a�Z��%� ��ss46Ũ���;��v�����)P��r(A1�7b"�řý.�;���NN���r�b}q�k��-���7n�;E����ݓ�����m�F̷2��[�O[U�ѓp��ܾ�xy��ٛVz�ς���Ʊ�f��K�n��Fw=j�F�p\�-��ڳEr�{�ی���mwi���`�U�\����;�a�rd\�-tc�!F:2��=6�i.ΉМ��bᗌqŻV�9��d9k�"j���n;yw<ۥ�yr6�u��Q��ڵoV�š�	��vx�x�gs*sۀ;�V�;[�4:G��&.ݸ�.�=��9��[���;��g���Ř;s�SI�K�V��8����L0t۰�iҩ�݉w�����-�2l�<6n�$c�%���c�C��\�2��m�=������wcI�ŻY�z��[��ۮF�e�^q��k�ۋ���h5�kr\=�N0r�������:۸�����ֺݫ�l�5fJ�o]�n�9�'t���N`�r�k��{�c۝�Q�q�Ѭv��y��C�m]��:�7"��t�&cO��֝�͹uئM3r�ǵp����-�,f�wI���m�٭���l�mf���̲+���/8�^qj��ϙ#n��Gv���q۪�燎ܾ�� w;S�Ƥ�Ӹιѫ���\�q�pI�8�{qn<�l�rq�\Z�q]��a����4[y�[ū�ݮL�9��YW�gys�rۇ�F�	7hk��R6�ݽ��zk��۩Π�bM)�:��q��&�sz��<��xo��β�;K̻����p�ˮu�vwV�r{9�7c���Z�nl����;ڻ�1]��G�sp�Ն���6A���M��6o^�^��x6����f�k��ς-�jY6��kv
����)���e�i3�rsc�|��������#o.R���n�'X��t��q�7[��B�����۶����܍����vڤ�ۅ^�pp����ۍ��g����,vq�y��6����q˻�8��Ժ�/[���v�7b�rs��c��AƳ�ݭ֍�:�&��"�㍜��m�]� ui��:Pul����;��֌gDsy5����Y˱r��URg��X��l�����I��q�9F:�*f���vܬ�hB"S�te��[�x.ہ7��&W���1��6��^��mf�q�fw`諎|UӔ2���u�QQۦGtn�N�uv^� �m��Es�{[������N^vԨ3�\q���ɝ�tjvE�p���ك��惯\=�b�FV�q���v�1V�pr�zݛ����m�R��YxfW���U�9�v6���<=����C�8t��LGN��\K�J;nM"e����R�-��S����U�=
P�8�������`1�j�Y�;eGؼ{���Qֽ�`#z�Ʒh�N�8!NFw\s49.�D6w,b�ޣO�c!��z۱9�p��m�}6�;ol�M8�9��GL��uɅ���h�/l���\������3Wn�]�`�����;m�Ӱ�.�zq�y�[5����WXѷ��뵷;�r\�<���x�'g5�ݽ��:��nn�s��[d�ʂ��
E�]i��6s ���㷫F,;�z��� +@���*�m��\�qØt�k�۝���ͶշM�v�����ۣv��E��X���["k�v��n^{�Sl*7Aҡ��C a��x}=9��޸����m�G ��T�c��n����x���#N^^N�e�Ƥ�9;�&�L�r�ѪyW���.�+u��n�m���r5�*��/=N�nd�K/`b��dyc6��z��5ќ"ri����A�����݇;�'n�{���J7z'7�d�ݑ�ط�m�@'�nZ��cX�_:�N�3�EF9�]��Y��n{��Mc�� ��]��2��$�G�,��i����r�=q��۠,��	��ɺ7�ڰPl�*8����N�7f�bU�܁[�mۮ�Gl�H�ɹ�N�y���l�S��lgL]���v�׭v��ObZ��b���ܪ�;`ȁ���m��ȯ<]����N��Z�l��s�6x��ґ�:��9��<�c����v����<A���1�Q����q���9湽GqvO[�7L��p�0:��ڳU'A�ݷ�]��z'e���m�q5ŕ��a|��7����v��{.�񳈮�����w����Y�ۍ=�qǝ�7��Yکwh�nNvSG<հ�jH,&kF3���2����\�����@q��e���y ��%�ok����� |`g��S���i��l[WdGr����Ɏ��ݶ�n��M�kk��6^�Uv1Ƕ.Ե������*n�tg�8��q��F��׭�V�qt�7g�s������9-�Yv�v�|Iʹ��f=��ћ�'�2���m���y-s�2��cV}As��B,��@t ٻ�����T�:M�<學��\�ݎ��-=�ã���v`�:۷Gj�q���Cr&󐃋��ۍ����6��s[�������[^�n���N�U���-�n^[pn�Ǟk��=�;�7kl9x�
Vz��`��fA$�9���i���s�������;�s'��jݳ��3>�nU6,�a�aj�un�=&�hHv�<��{�{aK�<��ή5f��l������Cn�.��Lܻ@�d������%�8��=�ۍu��sř�ÖG�Jm��[��N$l�ut �l�].�tq�!�������ڏ=��n��+`z��e�w�n�[�2�q��v�-e��ɺ,��"�Ź�M>���}�::wn�xM���1�xà�ڗ�WZ�71h�G�d*Hk+ϫy33���C7� g�q�wg��>�׍�+�g�	-]���wXp��ݒ�Cۃ��Q����;v��K�9��`��ÆC<��u��E�� 3k��X�ʖ������.y��<��w��[�M��񬇅Nrtvv�WW=qm�a�"S���٩�r�����M�
���:�i�s8���Ɇ�pέėi�t*��ov7E��Lj�zc"v��HEt�]ټ]��m����v�urA�v"xs��.�<��\@�<��{p��gG\<��h��GK�`ۖݮ��������3���7ۀh� d��[=pܱ�s����	� ��r��p��v�E�uw;�}Jz�e`�7Y9х�x��s.��O<	d͸�z�)}��ON���m�� �nv�m�ێ3�E��8��tۡ�ʼ\;8��j�qӮ��.����.68��m�u���[p�ڹxj:xu���l�48۠��	>�3�7��v��=���cn@gt�k�A�=g���^�x�Ǵ���ٲ��pvyy3����3�፜4��f�Cw^8d6y�cE玵�<@s�<g��KhUB��P25j��!Q���Y�[3vs�c^M�ks����kZ�t�\)�I۶0�N�U�93�n��	�ɹ��wq�YzF���'��py��5�4���n���[m��N�ڱq��͡더���ڶw8�;T�k��/^�$x��|���f�.޲�9E5��`3%�ծG�:۞V;^B�9A�ɭ�n:��e8|.���Q�Ǯ\��[g�h�yW�ۓusx�#��]r�N�e|���mlu�^ثg��8.=�M�=�n�/7F�Eam�֢��GnG��z�8Xv]gg���y�9��ư=�O;���;u�vv�ϮD���m�-���vۭ����Jrx�L�\ܣ��u�G-��6�z�g'���a�wWv��j���Q�r�
�Y�j�ɼ��m�]۹-�B�t��o�<$=m��A��ql9,rcgq\hͺ8AD��ǟ�#�`������V'x�tݺ���F�9����UĜh�d7V�=g��W�pr�ecm��g�b|��b�q��[X�5�+e�v�Ձ Ɠpn�	�O���utvK�N�V������5���My�h�Fq���w��ϴ�u��&���kruL/s�)9ڸ�퇹:�u�v�zS�2�tH�;�u�yT��[���1[J;OC��.;��@���3�r�X��w���`�mE�8gȻ���n��Y�uq����M�y;n���-�p-�a<��9Gj\\����\��z����6.�<��i�����b��.(�H7����i��f�Bݻq�q�;\ۜ<�&�03�/Y�<�.펋d�Y�	e3��H����PU!"�<�H�.5knn��#@��8E�{���=o �B�;�x�wn�Eϔ\���ڍ����ݻJE��c��g����nۜi��m��x���yأ8U=u�N3��+��Urd�&�_�Y�1,K3���ŋ331f�Y��1f`���Y���"Ėff`bŘ�3K0bA�$�bı��ăI`f,�1`ff$�@�%��bİ1%��$��Q��_������s�����C@?����j���MCh�Gq/����x�^��G��L�u[;\��P�V�HUh�~��W1�s��������q9�0�-�qQ����3v�=m��d3�-�@��QT��ݴ4ׄF6��c��*M��%�ʉ��U�J��vK�n^�?V�Y ��3�#!R�`�Y�<o�{~�޶���C�GO ��N�y�"`,V�������"*.�HZ�>h�a�(�,�Y�� Ր��M����VOM�uuHp8B�W��=\[��g�k���c��H\���/��4k篠��m�sK��nH�^m�q�L��'���B�He1'v��,O��"lƍou͇�¥)��Q�W��K'�l��@��|4��g��1WZv*5w|��"3�T'�H/M݊t�������14�BW�Ηgs+°߽�X��3E!G�7r�gN�6��p���W$ܣ�R��Y����
┍���qv;��>��t.l!�[�t/$�gȶMRհ���]l��F�=y\n�ɹBQ�i�tf�~ǉ��P�3����i����S�j�E�ThF��.6ԬA����d�u72�uH ˘�M�X�:np�i�ú��7�;�,h��I�b	)����y��8���u�!�0�8�sӸQw�m��ػu�	sC�z9�W6�M��^��)q�m�g���}�����T����3���m��8��෰x��ۍ��r#�n�`v��^qֶ�r��ػ<[Sve*��-�9Lp��x�l�VM�'�3d�:�S��z��6�p÷gz�9թ**F������w�{����-|�&��=X4��j�%�������t�;�[(^�rJ���񬡃|����(k�����N��=���B;�߅�ڬe�j],�"Y[���S�^i�羚=�kN�w����K𺰎�4&W]���ʱu9�a��ؤ��xB��a?7�|�)�W�I�һ��0\��]v'��`�7n{5��ڷ�)�rd�
�{D!�0���-���(@p�x��Q��+��ixjP�&�fzgu��F����E�oa�M���X=�{G���׀�!�aީ�b%�%ka؋J:!��&��A�L;.eK&�� 5Âلb{#�#(d���4���M��<���^üB1�>X�>�Y����J����=�@{R�������]N�m��m�η��F��ڡDZB��Q�,�ml�˲����J�7[���Û�NP��$F����G�yCU�_�Yc_��8���r]�ސ���F�h��W��cg"�����5Mi�R��0p��̺�1W�F�fǁ
�����R�Yw�\k��M'5ֵJm>�t=�O/fj����W*�#H�z9і�%��U�Y�q�)�ٶ/�lK�Q�
û��±e+�T��6������m��	���[q0Mb��Z�@�fd��;�����+>Z�cM�H:*�Y����F�G�v9��tx��&چ�M���\޲u;�fIFѱ-�Ytg�֬M��V�v�!��"�oun,s���Z�u�T�Y��aRk�8z;�W�yJ� 4��[�#�j�y�>A!��^���^���Y�2�V1�m�79�G��T�O��y��S��(ڒ[On�j/��������&p�$�������p�Ș4�"�G6[��܅�:=Kq��~���FxQ:f���p�+��i0qRU�f���F6�����&e'��F�VZ�H��v�H�ub��\�v���`�p����I5l�׊JF�
� E�.���B���y��tH ���Ԩ�rw%C�+���ӻ�j�4�
����<�Y(���\{��Um�Yz�,m��2�Z���>�O#p�ȇ�ny^o	&֣XJ��u�Ѭ�����{�7���vb2Ꙕ�:3�a0���`��ٌ'-�RIU@��܏�z��M�����_;��17,��j��!���zu\�Y�xn�e���n�fS(Q:[*�U�z�sv'N�^�T�*�:�]X+�s���M�6d�|�6���#������G��}��޳�VR"�4��Dkk���w��yy2N����s�ҝ�H"�[w���s�?k�e�p�S���M��������F�Ѯ�Pٕ Dr�A +�{F��"�1�ݶ��銖���i�iY�iv'W��1��A���S��Y�n��tyYT3�3.�w�ZM&������� ��T��(XQ*�2�N�}e�֭m�]�Y�>{���7�gvh+s���Tw��2��� ���+��Tj��qb��@9=������e�+QoC���5Hú�^lܻ�E�G�Y�#�R'N�U�Ļթ��*�j�����m3Li��N�W���*P��;�mڸ[0y��I��aAza,�.)cqA�hv)0����]�v"h�C�����K��	0]�N�wbَ6��%�;,�Z༰EN�<���}����x��[�^�Qza9uug>XV�T�u=!�|h��`��;[��k Kk��߶�.@h2�n�;�d���;�.��Za܆�"����"�DC�3�X0I�4���ժ^�����`��S6��L@�;{^�KO�f�M��E���/�cK�T�Ϩ�M����:<�k���Wo-u������}�yH���qǠ��swU��hh;�6�N��շm��P�5q�7*���:�qG���^���V2t+&�h��e�!�Q���A{u@@��x��}b9�=p�:��r��2��^�5`�
WI�'1W��I�UL�,�>Q-�i\��X�Ƌa�� �a i���mv��}�.S�e]
*υ�Q�GwvD��_ͨ@|u�%e�LI�c�X���P��8�X���$O�)g_���,߇�Hj�c��X��7*T���){S��E�k��<�7!Sl���&��]�$�m��ۢ+���q\�k�m �)�ݱ�ݝέѱ���Tg��2�c[>�p�@�6���;�^û����d<�6ּ��(Hs\��U��^ܬ�7I�4`�ϪM,�L��@�a�"����j��2�-HOj�x��qN=��K��zv�,��zg��<�а���_��*�a���)��w:,S���⮯���:����{Pgm�ʗ�'k�=�Vf��ٙF��"��F��
 �8�B4X��7�$�K� ��p���5��tu���Jm�E���@�4��QV��l�Y-�TaCl��įJ��ݣ������uz�RJ���,W��պ9G<So��j�4��̔�����ep�h"w`�,�e�1b�{L[����o����B��7#rI'[y@�VJ�TKP��i��"�2��;���M��xC9x�4�{�N{ �ϥ��v[e���G$]>�4KF�?�������f��rC� z���;��$�\6:ݻv�r�dh��2b�SOK�nǧ���ٸMYy���l:��sϮ �mn�nv�JG;x׉�f۵p u�U�݉wg��6��0����rW����N���z�!��Cz�:���F����>��S��U0�8����p��M�����Ѡ�}v�"��uj�?1�9��[��o�[�Sƶ�s�����Zl���f��(���A����lz�<8P�.Ǔ��P3˶p}�e�`$�H���L\���'jb4�k��ٖ��P*9� 4c�9��N��x�np;2��i�;a-����9m@��52��nڙU���X�NԷp�q���a�vw["]b�#Ob�a�X�f$��U�	l$F�@���+ch���F:4����Z���!�)�k��;�c����f���i��W�Yw\]B,�}�ٹ~C_�m�)\eV&�:'w;Yy9l|w�hA/$�wg�DP�o'K�OkI���{��f��\�ip��n�'uF�d�*��r_]�W��L�g�U�>��q�Em)���F�g�w\��9B�|k����ݩ��+4{({�Ļ0�k�_w��ie��x��u�F�ضt��m��G����[X�-�_���z�{a/m���k��N�`���G6G�n�����<;T/��[�d�EE7Law �T�z��:=.��5��
��e���v>��&��>"�t!���eԝ}���l�+l��[�ѮW)����ZS�5:��̟���f`��
bfnj�<�,݉�Mo�!]f����o�}����Z[��Waݨ�ce"|��\G.��=�]H<��I��\6e��,Ct��948Uv���o$�{�Y�q�޽���2��L�=�sˑ��u�����dz��QUAQ��}��\����;0EV���r���em-F|�5Ƚ�^��>�|P��f�6T���s�M/$
;g5�%)w�Zs��b�������0����BY'��6���8��̅��$��JTt������aC�L.I ��4��Q��R�T���D��Oo�z���B�Bɴ�X������$ 2�O�J߯9���C�h��Er�/��vAմ]�z�,CU?E<rωJ]dHڀɍ#!{O��%�y�`�	�%��d�V�]cTi���1�h�oՔ{ܷ����x㊖�����np^h�`&��29������^����8*ӛ�c�L���`���(X��,��xɎ�*��g{�co��{�1�������vO6M��е���ʲ��v�h�LmgcV�P�V)�Ak��~���]�HBG�]�+��N�\'��|���{�C-���*�(��:��ϻx�٬���zE4@Zk��
a���0)]�57p��p:�����0�*E�xx<�]�9��yя2�J�ۺ���_#�*���^[J4���6�k��F�����+T&��6��Nd�U%Fk{t5j�M"�-m	X�	<��K̝MN�2��.�]_��4�텫���h=]��]*�қ�DEX���7[���2�E]1e�	�|4bԨ,Wg��>�\���|c��u���_�VH�H5k`޺�8T�6��El{�;������\k��(
O_�����IxY�:��B�2�U��Bov��)|�C���N�Y�8]j6�;�o�}W�}�7�M��m�׻KC:���]�l�_����%�Xu4�	>59�� 
����>:2��V��tS��o�sV��&h��!�V�����ybi0W�����'���'c�N�"%�����{�*�â�ɦ�l�Ƭv��*ݸ�Y-',s���mǞ�h-��)S��RZ���?w���5;V������骖2��f�ɡ�#6 �E^�O�GK���o'-�;%��P4I���̶
�yrѧ��,��r��,N�9��2�'��)3j�n�a�M�rH��Y�d/.��+��{��@��tA�40���Wt�4��6�]Z�/SJ�ۣG^GJ�������+�m�9/�dȲi�V���ו5v#�ȗQw똫�)���O{WE9pHHl�4Ka�W���ܬ��%�v��:Ҽ*�7�Ҩ��y-�>��N�� ���In�2����q�g�<.�@Z�F��\� ����jZ��C�����F?v��+�<���퐷��y��\��W\P��{��'F��ي��u틂F����(��+3��فu�/A��J'=kwS�v�GE6�:7�bB�,R�M0�h�Fv��J���:�mq�k�����|j{3k=]����S*~tt=����t�'ǒWqq�w#		���8��HG�NǢ�<+���ͫ��
tF���h�����%>n��Qd��#Эf�\#۲�i��wJ9��N՜%�u
�ݼyY�ᠱ��n�F�n�3����BYzk�~�W�SKbyz��0������9W�2�
i�Cݞ�eHT���u�4�;c`ڥ��BR��P�w��{�^�H��c�_��B�ߟ}�^}�<������B<��+~��>�&bܢ	���Q���A�*��Y��J*QU5���7�V�����N�iT��>6��uv.����{!()ђB��'�5����@ڭ��AX��I�t�t��	�q]�N�s��p�xd�׌m��xky��#��Z��=sKL����O�w�oP���h�ٖ�d�w�I�j�ݰv������p�P@��k�����u�]ؘn���'^����n�
h���[���N�Y�\���� �캆ض9r`󬼐5m�3�1Ѽu�&��Ƽ���j�g���˵i$Չ��,�ǶC�������'\��;���j6@zz7Fu�[��❴\�Ԫ��&��2sm��������7mU��րVL��&D1�iX�PD�1��F�L�E��k�ֽ/�x�����M1���-m&�D��4D�]�;�VUf�뱚g�C�K(�j����uc��v�Af*gY^Z&&i�"��n�� s阺r\H�"��^�.��.,`���$�8�z#]� �U��,5�M�,7�h�.P�2RP�G���߳���{��Zv�x<�׉�=�E���:�����v�s4�x0zu/n��8`��!�4Ch�|� �q���u�J��(	my���\Zk�h���6y��>6�:kZ����MQ����+X'�|X��@i�h]�k\�#h����ȱ8"�)@%@ޙ�� z'}[T5��WuQ��B:~X��.q�k8����XT�]\���`{���h�"�6������x�fg#�u�#njݙ:<��@-t���i1u�S�mC�O�%�o���0gZ[��eڠ<�L0�C¦2\M��5g^���pJ�a#�Xf�q��t@:z���o<P���,��y�g��`i㪱��e`'�uTn��])˷2� � �#�U?7z����ID��C�7�:׶��^FY��齶(�n�x���I��;\޼}�i�4-pP���c�x�s�'oOv�懆��g'R[ٳ,FcjZ�?wR������?Y�]�ַ4�f�����I���J���}��	��Q��C�K�U����9ud�ysM�v[ˮ�{.o�U���j|���@��:�ѥ�N}�!��Q"�x��!�d�I� J�ͬ����È��/�'��p�����ӵVFi�<�t�C��{�mf�"!Ꜣ|����̽O�K�_B��t���+��x�蕒�㵝�����k�N�Vev��� s��Õ�ֹ�6)��[k�=vz͊�W��<�iP��y%�㹦:��n�lҵ�����p,�ޕ�[�Ӣ��[���tV7�V�����30k:���>�*�Ƿ�;h��nb�Ow�G#�Gi�����#c�M�'�xf�Xk�i��F,�YMC��ܿ��ѸP��+�����nr�"__+���b�
�$]�A7�+ę�cL�A&�a�����QTA��'�fC6�ky�vn�;p�'KPe�QV3r�b]Q��삺�@[�$��tLX��Y�L�'F4�/�VG�kЊ�t���c*fF~�ݱ賚��q�W�K�����_��Tۼ�{�
t\���"�v+����68�`����̴2�-I7w3�u��黣٦��x�M���<�7�Bz��f=�cWp�P�۽ӧo9�B����=�t&��GW"��b�u��Uj'Wb��Ik��[$�]/��wq�)LN�ׁi�GT����Fwo���o�V
�����d��*�m�VbZ2�]<�0�P�H��$�t�������@2������9y��Z#|<m�7m8^�����R�����x�򬱛Sq��gk;�9�h���q{;9�y�t�8�����˻]��y���'����y�6�g&�ٍ�k�c�an�0v�K;q�8�]�b�v��b�����s�ַa�W�d��ٳ�E�9�nl���n]ąì����î��V�b�˫Z�"�;g�����ʝ��6-��z׳���{v\�x�6�]��6aw�q�Ub�'u{Y�x�k�"L]�j��{n��p����<c#�V���v�=�u�����Z��Gq�c�Gi�����sv�r��W���s��ۑ3����{.�p3Mţ��^wfݍ�-�������Qq�vv͔��غ�����$f���koAl˻"�N:��N��w!^.v��v��q���z�������E�ۥ�@���xNt�o`3k'l����͠�D�0((�#�ؔV���2A�u�۶g;��\\�mu���'Z��6�e�uj���rvWrd��.+�rf{�qŔ�L$pl�O`�̽%��n��o\'�jzXcv����Rnф�Ecő��pW�-�e����mm��p�"�
Q㶶�4��n��gU�ێ�h���V�Nl��;I"Z�qѷΞN��η^VCt`�Ƿ��(����'%1�x��u8��������sd�ٶ�v������<�k\�k+���v�Ź{G@h�{];��F��M��Ɓա�9�c�yݫ�[#Ʋ��i�����Y6�;n���7��duC�[q�c����Hg����u�7]u�g�z�v�4�4Y�-�N��ܫу;���s��i�\���R8�$���u��^6ϋ���:�q�{�S��P��X�����@ƶc���j�$AJ�� �8'b5k'gm���;����bϲnNq�у[0�%��XN���\�p��G �V����gm��.Ϋ�+�����؊��R��/�鋧�ޜ^k��4-̇� ��y��ެK��k-�Q]~����=��|r�R���ftTH;^Q'��bOm~�^2�ޟkX��5����V��ؒf/ѫ�\��������TnɭT2b˽�9�����I���5\�i�n��[X傏����2	}�߿iy��[��@��J	}Sf(b4�01Q38��/�V���hTI1/��Е1l�(-r���j��Hm|(�gu������%�:҆.�S���̂��$Ej�Ȳ�]�}>��K��`�f*���m�JӤ�Vig�k5���2�bfC0��{���IpPLX
G�G�xT_B_�����Qo���/鳂ًBZ:��M|�|C%�ӏ�L_����}}����o�޺bщ���ļ~홟�b�$���kJ���ZP��XĿG�c@d1C�/�|Mp1�ި���n�J$�)BE�6if�E�K�ݡ����3� �vg�V��Jz��1�u�*�����Z1�־{��f��	X�i��tZ1{�{_3�/�3F``N�E��J���&b�EE`ק�k�J~k��%�F����a�bP�`-��/����|%x��gt�%��}V��������*b�Ǚ�|C3�^v�=���F/�{�v��ܑ�*-��|pKF((%c�	��T�S&������� �s����`����#�	l�kbJ	~4|%Jsw\�(`&-?W��}��n��i7��|&͐�ϯ��^*fp�.�Oļ��%�k���-�~�*b鉙���l�y���޳BfhI��Z]1Qf���s�y��zE�4%�o��Z�����K[�Kjo�3�{ڟ}�m}�5���Y𡋦&.�k�ţbВ����OB��SePи&/�S6$7�i}��TZ�X��b@�1p��[��,\o3��~�1h�d-�1Q/��O�7߸y�LV��6k�������p}�S���K�2���3����&%�"<\11~w��0�����"-2�g�8� �~T�bit��6�~�;��f����Ɵ��Mxφ%ؓf:G8�4�vg��)M���8E|�`4x�Vmwɇ�#����"��Z؀NPbtv���رF�;�{ZPe��1|g+TK�|QoM%�v5�P�d�ÿkf-���X�x	[�Z�I��7�**/_�֓2��̆1p��1S�B">�����g�)q]�l�n; ��1��e��B��|��#lMu0Pj7���2�/x�
+�A;w,!�t�c��ٸK�S]�����U���.���*j[M��� � PK�~1S2��7�b�N�7�ݩ}�τ��(���D�t�ė�J�����~�Z133��>�ĭx��O&�d�����R���5��6��߻q$ă��d(-
NL]�洲	-��҆%��ŉ��fw����>����VR�m%��:�b�q�Lh[#6�&>k�;aO��G��]�~����#�������;�YD�����w�T�%�-���k�f�L��T�ň�ߴ��_6�i(bщ�8 �s1�i<�G�sS1a(DB�K�+�_�P1hPI�xY�V����o�f��"y(���іY����f���%���GZ�[�>�f&bb�_sIA{�lY�iU�3��ץ�	��2���������{���$
�賦l������D!��J����}�����x�i]�ZZ��1��t��ļ����b��~ ������b�(g#I��M�T5�1|A(+����P�F���O&��,(54���%��}��5�G��/�$�f��1-K��wK���^�i-	�L��q��/Ն%MG�K\��r͊�XK��9�ք�Au�kB�m3�v�'�"#|����#�-�����uwkN�o�.��f.���]$.��!�]�T͘�bb_���2�}�{�X����t�"i�WE,�i`(~1lTJ�P͙���P���𾇽�f�ēg�1C3F1b�k�?j=����;��"RUnRc�r(�uFd6�9f�`4�������MI"��br�%�C3����>k�R�*Ab��@��-���J5�{��-�Jo��<f1h�`bщ� �rhKZ��v���X�pI111�f|c37٭'�.k��ܼx����Z�-k]�����X���Ή?��-�D|��$�M�uT�.9�Ԟ�6	��jX���7��Z�-�'c%V���+^ks;QA =j{EX��҇��-{w��&��d�u�<��(���29i��A���{)��o���I�|O`�W6���f�78fӬ��w��ۙ��*L�m�˶��슸�ׇŻ��VS
��;@��ڮ�gp8�ٞ�\����=OLU����	l�H�ޜ�'p�k*�;�7�}w+V	�����'�.��b���@�OZ�ɦ���0ɜ��ۭP��i
��6���x#��$R<��=��Ӵ�������JT@�I;�ntH�u�Г^q�}�`B��(�L����Tn̡���O_n�^��[�� �׾n���r��T+eGx��/��:���f�[Ω�ZP���D?^�&�{h�b��~`Sw�ӓ��?]�&�EXU��#\ OW�w���
��[�w��u�g�W�5}}m�.���c7��õ.��8�n����ݹ���ޞ_�C0�A�Xf�uD�Ӟ:T�~��a{P�B��<HqGV��^�Sڿ�������\z�hs}�;ռ/Z�D6O�)�1�ՅX�(3GA'd�g4�'&{|iח-��A�*�b]�>��z`����\�
Ѫ��}M������B=e+��!U�n7�\���a����� a.�j�<A��]���.9���.�����'e�ת�+�%�[.X�L�m�O����޻��~�����	l����ƗZ�/O�Cb��3�l�ژw�=�`U��
�ܱ�v4+8�]�u��lV��e޵:wm#�<�������фc� G�[ ug[��]v�oL��Ţ&b�ՓF/rdMj�nl4�AÅ��[2���E�0m����6c�=�[qkX�7:yyyS�GrV�r�9��l����mT2�:��iPp������p���X����8:�s![����-�6�[m��w�1�ٰ	kv����,eq��קS�/<�*X��F.7I���3՟ggvi=p#�q�guVGv*ۮ��N-�Z���	�ET�j(̹&6g��B��
���O=k?2b�+�B�Qa�B�����~Ky����G�Cl�h4�p�VQˠo��h�C/�JJ�z&+#��&[Yp��GA�	�����FI���g�d���2V�ת��F1��vu�v̖�͜�u^����)��!��璁�ه>(�F$]���riy��=�q]�v·�|�\��B\W�,��^�trmGU˭��y\����p	���;�4`t�XKl�wp=�FCWE��H�X�*�dgj����|�M��MT4z��>�,���9FS{�M �ؙ�R�5ի/8K9�e����|4�;���MN���<��g/VxU��[H�����űH�����~9V
�YF�  �����%���r����|s�v�d�5��77���=P�y�E{�s��Ȁ,WP������g
�=3�/+<<P�Q�۬W�I�{ڑi�	����X���؋��ڽ�낊�����ww���iv󞣵��G�f4��ק��{.�u{nq�.�˰0>�Ă�{ػ��ʇ+i��YN��Ժڇ���g�݁ā��C�u�P_�{c�.�o��^����C��i�������O_�����Y}A��2nv^p�Zv�mm��,B�3Ml���;���y�;����+���`��*��2čIǰB�N�T�kk�v��TA���^����n�;޵�MW�8�����B�_9�׵�I�ZGè��3��RG�2��0�(Rq7O�s��+7@���CG��((�.�3f����� �q���;���|޲-�h��9����Z���VH}����	�g:��\�*Ѵ�(ǡ��)+1m*�y)J[��a+P?,��Fa�^@n�3�p�7���g*R	��-]���������C���/q�[�:��� �YW�C�*���`�fe#����y�ÅQ�GQ�o&ń0u��7�r�y��uo�����CMb5��2�B�x�����s�������� Ѡ{����I���oD�B�[�0�aU/Q����Xc*��ya�Hg�,E۴��?d�?�r\�0
0u5��-8�R<N�P*��@� �㵗�$}F羞%�ɝఊ��*@X�h�U�$zH~�B�Һ|o|X����+ZJ�l}��T��r*�u��c��[�ݚ<�
�<���}��ҫ
�i��5r�)�ղ����C,�y䣒uSrQ��&�v6�o#��,٪��q��C���f��;�&�(Ry�����APru]u~9^G6�<ܱ�;d|<NkK}�����1SR�7����RΈ�$�`��Ɯ8��ȭ���!�G����W��}���v�]��@qe`�h�b;ٮ�4+r�#��~��sz�x+�|�
�"����hp]�{n�`[�,����(Q<|yy�3R���:��<�/x��������
�F��{����'�#��Ir�~�Z��7�>p�W�� �^���TO����8�r�Ç�@>��k�SR��^�nuNBA	�|�]bK=�b�wɼ�#O�I����m^ Ǡ�-��¢v�.RY�:=�b��dOr��O�8��;��,��8���U魪 ��b��8"��k��~��	+��"+"�K�cA-h��m�n
P|#=Y�3���=��'3����M�U*���T)�Lu�@��7�.�|�Ҝ�� ��̓���!�nٽ}K�ߑ`�����e#幺��I���k�Zo�%Zmȱ^ron���i=R�%N��h�b��tu�6�&�ۖ㧆��j�j撷=��En���������?_�W�4t�#v1h��XU��(c�!�c�a{[�;��c_�� �y[B���@J�uI �4B�3L(�ݙ�Z��j�� )�{��B*���{.s��-��,�X)s;���90 �3��C�b��=���5��O��׊�n�vE����>�I���@���uo/)@���N�ڋ�Tq��ѳ����!����a6�آ-%]�/!Y�u՚�8o4c��|�ݲ�Tz��j�����"�u�<�C��1L�T���6�Jf��mq�S����4��|����oYD�g'��ux��_���VF�W��\���Փ����y!� �b�M�4���.wcmeo���3����p����
�)�CJ�͉���n��+�G�ы�y藺��*�*�H"��E�~�cLx!`���]8�C�_�/�H�׶��e&����"��vr(���<N�U4.�8�gb}ն�8o֚"�'�<���Ѡ'$�C3��`����Ǐu��D�^L��{�,\lB$�%�ӁƯg��	�s�\7��3O;l��f��z�:7�9�۷G#T��b<� �OD�n��t]�����������_v��V���0�S�FЁ����p���*�<頮 +�L��+i
�ViC����B���g�(#`�-T6EB͇�"�V'�����ܶ�^�� �qr�=�~���N7H�촌�ۀ#�g-K
$�;z�2VK��s�띺v}���V@�[.���m�Y�Th@�Hu�^�|q��9jg&���i_\R�^\�㨯2Jl�ڄ����{�I�p���O��O2�$W`T���[��b��v���AJ�G:�i��o��Wm��x��)�������x��D�����h�m+�D��#��u��ҝ����y���n�����et�x <r3�w3:x��^N/%�o��]��c�>�u���r!�,�n
�u �!�m��]��;,�'����2��~t���Wn^wQ����F�����]����\���uz@m���n��u����b�vX�Z˃�|+s�rS�42�[;�u�s�Gb�`^v�*���A�(�틥�+=�6�swc�,B]�Ң#5H��0��F�p7�I�G/T�d�[�|����VR5���A6^p���Po<�D�W ݣ7�x%��3M���tϼ�LT%�+'�xF�^e1�N�em��e�[dF���m ~%j>e|���I'�_u��㯾1 �Eڮ�H����}w�>��J�NE�qI�r�Ǟ�/]�����v-۷\�DI!%�Ur�w��.�zz���l�Q�dk�U(9�s*gb����.#i0��KjbY�g}8�!�-g�^����6k��	�����9i�51\��LW�'�����z����Y�s��o�}1���T�OeZ���5��c���5�ԏb�q�Ŭ�� Y� ��XH���P5<ϡ�Za�n��[�7�1K�����k����:��[�aqm�ױ�JpY�9^٨%k��޻g����V�8��F\Ӻ�z�A���'���d�����,��fd�kA�B�9F���fv�ح]��4�����u��>��F:i�f�0_��wy��@�9	�o��K�7x5 �|_�$�0D�ձ0b��d�hN$R�ױ9襅�$�IZ]a*��Ɂ���^�D���Q���\���f�h�5u�Κؖ�޼�C���u�����򒮦.�w�AlY��eo1V��L�r�����](XH���Jy�=�nά�o�AʘΨ�Sc���~[g��Ǎ����FY���VU�l�J�9^�oA�(e��td�.ǐ���#��⓺�	to@�T�Y�)��t>�8��C��1�j0���������()hXI�.W�׽��X&+���"�*5��ڻc��TGƼ����@�A�C�N��:�g7��^�i���X�ҫ	]�!l����Кy�1g�_���~�����0˱S�
���*^kf����nf=�J*���jQ���r���
:B*�F��������??m�iݭT*���t��Lvl�[�gh�Yւ��S-!Zrf�3k�V�B��o�[�cؼ�j���w��J�3��X%U����B%w)�g���\ ����X�1����N6���=%�u��鹍^H�H�0P��+��G隨�f��+=�c_�-x�C��Q�:2@�Y6lmz+q��C��0���u?zV�d\���[uۺ��{o΍J�[�O�yݾ����#u�0�\�;F'0�B�$I^tE��"bڶ~��k�����?y������0�O;,#u��ytcpQ]�<����ۄK�t>ݡ� r!��Cv��V����}����/�,�=;"�+�A�:�L��y?\����}�o�^H4�y	�n�/eW���mM�!�#T]I�EM�]&�DL�D`��X8˻���θ���L�sr�۽
���Q�N��47a=I� &����QcbT�C��V0x]b��������y��Z��M���1{6�s����Q��l�0a�ۢ/,��^��!$�BE����=��x����m�����A%��1"�۴���xv�ˣ){_�����N�W�gV��cإ���ʴ���Hp��I ��B�{*�9�mH�q7���R��i���׹����G;�9ؖV�;5f���ynߞ}^f-��n���9��u����`x� 7�w�����q�nF. �p���g�7����Q����?y��X��+G����C��F�K�TW5e.��	m���UWޔ(��t�0��
'5��[��F��7�i����(���"��@Փ>�x��W<&�pq�Y��{.�۞������C~�;t��)DC��q�!�]i3<�l:	{p<�=�v��7�qc�_��v(	�\~�k�����w��k�3Ը�u�����o�N��X��W�>�1����c�G/fؑ:�&0�P��F�o��7���"Y?LC��'!iֺ��W���<���C��%��&(���5��-9�>����=�g�����r�]��m�.+�jQH�/y���Q �FGaйmb����:���L��:��Hx�v��v�I��]\=t�g50�;3Z&��[k�e��+�4��t��p���)�yZM�}���:us�+gL��lR�������\��ʣJ��+�f;���w͠����P�?[�o>۩���ܦY7w���JȄ\[���#�&�̫ێnb���],9����0��M�幘B&��	?L{#.=���x�bYN��r%,�n����=���"�y�lb��G�Z�Fs4�͘��L=��1���*ٽ�/�is)�ηYᙠui� �7�K('�%�(�ƞq;�Ր��$�1;�}�r�Ri�7���X{���[�wdW]��l6����t۰�m��؎@��>��>���D�[��59h����6�̛B�0����v��=��A�݅�}|n���~%�l�����/pU�@�g�����Y�Q�5�㜘z��&\eô,��(gX�u���ьn�{��9[C�YE�V�v�{)�+&�e·�኎n.��9�v���L�RY�w�(�8}o���*]C�0 ��*�3���|��hru���i��̸�X�.�RU��z�^��j�3x����8��8���9��xz��`���@��%wSsf�c���y�#��M�y��^�y
[��������c��r��aX�[��R��呮���.�Hu50���Τ��@+�����k�ek�]����x����{/�#�\�z�y��`ݳܵ�ӣ�9��vw��Ղ���!wL���v��&�R�PA�����K�����2v����7��WI\6�[>V��t�`�$�~���٘�u/"K�����| r�#[LYԥ�������^���3K��Q��[�>�ϱ�ٹ���^���.�q�%����Jܑ�j,�h4�.+����z�ѩ���� ���ϵ����(v��H��^�t�W!�{�3E��f73m�wZw^M����>#�����u��u>
��^}�y�V<��({H��/�y�uޑ��}���&��F��*$�.Dr���P��kNR���Xئ��.�^ບ�(׭�Ǎb4kG�y����;N�����mÕ�wu{EP)h�(�H�f�(f�s�46B��5�xgQ�Cw]�{qyu3��*B����[k�CWڈ���%�^�rkѐ]�y�%z�{)&zo����ԉ�PT�L$�J&�A�� }&-^\Ƀ��]�^�$��پ��z����E��{j���/�t}��<���OGZ	�u�8 ���{��y��ov%p�0��5rL��k	��"�w��m�����t�s�b���S����n�����1�gU��v��-�|�8ۧ���m�s����v!
�Mi�"��3�wDT��)��`��5m�DX�ga�{���K#j�v��I70upv!��\�ll��Q�st���o[Oo(�5�+s�����Ev���ю�g�k�N$I�n�qp��liwl���Ex�[O������ڟ���}����l�񵹇�;aTAt�+�����P��o�:b���؉Q�+^�z��kt�.g��*����q���w@�?�l�#~ȨS㗉�F�\ۛZ�w��5׎���_�s�<���*���qJ��=z�C}rI��J͐~�w.���p�mWO���#`��v�O����:<�,�<�&�d��e����םzG�v�,un�1zkƈ�[�����EK2;�:�g+C�sf.��Y�� �#Vn�6/�v�Q\TX�.:�7Ϲd�)i4w�̏O�>�|Z���M��gu��ឫ���I]Ѝ��U�ְw�̨�7�������jrA8�S�f����9S�i�9ޱ��-���QӁ#Z*�s�{�P���S7f{�E���|2��J���{��n��ыv���iZ�7f�+37Zi�6ߛ@2�*�i����n�v���L$��h�?{t-��V�+�{	j�h����/j��_�V66���3_�I���Zͺ��ֵC!� -��N䟙�&��go"�3AN��^�ϟ���<����ԕ��<1xl�y'��FUV���1��tT�9qUݛ�Ν�m�=[tM��Y�V�Sܦ
ݽ�ڮB����^��(�-�Ҏ����'Cv9d���n������zY�ŹV�č
\hҔ�ޛYfH;ʑB�$�l��o("T�������ʪ�Id����`@+��Ļ�݆j�� ��u>���Q�ڝ�I��m��'������\�'��k|o�0�\9e��ŀF��xWUWp�CJ���]o_h^�dVK\qU�â��ȕҙ?Vv]�]�i���z���T�p�" ړ�q���'���]�?n�[Dl���sQ��>�<��I,4]���77?J__w���I���/^Np��.����vn՝�����c���im���30����,���;~P���~_���Z쩡�)	�7����r��{u�]� �nL�k��6{`��_ui�W�y^�����ϲ�� �	�3}2�����v<��>%�FM��p*{�G���5�^�~PFxOt��L�d��&$s{�gP�ڱ>�kǈޭ�:�,���CA{\��{:���Nyw�ޒ�
�b�?z��e(�\^����e����`%�Ӯ-Z7S���Z\��W\j!ѸI�g6d8^HcŖʭ���@����V��)��<"t�>���x���z��ͼ�K����|�Z��}[
�s	��wxu�ӎ����Ѵ�F{1�y])��/�.�� wH��cokf��6�^./Aqqm��4�5���kţ.�X�Ԕ��tСA��ƷWziF������|�_�_����������ծ�c�4��{Q��6����䴢Z ���=�R7��6��gڶ�=tu���ݧ�E~�̡��Z��YGNz&��Q��N�/�wu�.<2C	r����xe�l\2w3P�M�<_��*s~�+��Ӌ�}��,��Dc�gs�m��/��?G�N�z�%-����G�n�R��X}����2�hz�T~����x��H�VR4��1>�(��Y���֗y�# ^��ځ�F[�2�T#HBvL ��������3Z�/����G׾1U���l�Tk2Vf�>��[�w��0��[f�9�ss2�1��z�l�G�_\��u�r��q���N��\�d�붂�KkR��ܵ�p���־}�=�)򫺾�Ӟ�q�|�jI�\�9c���=��ڼb+ɜM�Ǜ>U��ړU8�`lB�x���k�5��)���wZ�cƌކ�N��^z�
Jf�ԯej۰V���tG*x���+V9�M�㾒)�_��1[�w0�:�j�sq �֙�*`@$�9[�]К��,TdC]P�{�6;�+5"�R�WU�k��5̹E�n輻|������>e������ᾯT��8Ԛ�������/���*rV��QT��[6"����Tɬ�	!'�Bn�-�	�#^�s^S�>1Q���x��fj�B�e�^�oރfJ��tT�(�T����2�36t�o�&�#�1��h{i���p^M6�����qOA�{2W�_��bwM�(�罙9�����ٛ~-�0;#��֕y��|~���{����L��o<�.���� ���+nЧ���I&��mXk�Û�˗��*^50֏�n�j�W��sT�H+m���W	-bŒ�q��a�i-��26�$$���Uc�_s��ք��q��$V�Ꚉi����%���-����>}뛏j��CF��(?��WAJ�����L��斓�ZMoe^{�f�lI]�ddS�X!@�nG�z]���k4��y�[׷�V(x��Tk�˂���� �HW�5f�$'�e[�#��M�y��{�G�κ�}g��u���}ʥ���m!MGn��U�(�f��o����FF:ܪ{i�UNݮ{�?RcR����&��w����g�.�)�b6�c�C�C|ȏU��g�[
�`�Ȅ��Ջ*vՂ].�����ƛ�w�&n+��9!d�ԟ#��,^�褾�{{�Jmg,��R��J�1��L�F�ymc���\��
���"������yP�W�im����8뮽x�wF��K�z��-[��W�jWӶ.8Iق���s�z�w�9+u���;ĥ<u�.�%#v]�k�����p�g�Y��bz§A�K���N�=m���$<����k{7<��;.}��ǈ(�.ݵz�*�<N��5ٺ�kX�yx� o�{�oӯ�߳�hM��� ֛ױx��K��=��ڄ/v4��T'� �F���)FaA�宬&�G�ᅯ$J�ߒz���F�e�a �ηǹ��D�?x�Y�!���i���a#��Fl��]g�X47g�.����4=���ey��wmxU�������[po���o���l���)*���,/nq�[fȼ�h�7k�%�\dei�F�~Z'{�������zυN�v�\�oB����Ѽ��sʧW���b�}������<���_]n��M�Vz�lH�U� 
��,}��'��.�<��2�t~�<�Cu��*��i"��W�<�����vX�z�X��j's�j)���C�;O�mk�.�x��~�V�0Q6�
�y�f*�iR�����iH7�b�ix=��͎�{�eyT[w����̬��}K�2>c���H�	$���%z�K9�[��r=#�����m[^3x���t�O����)z%z�j�p/��k��&6��
�_�5���y#F�l$Q�~R�3�9�&|=c�h��ӟ ��`]׏��=�t�/:?��Z�󒐦������>����B�*�{7r�ƒ�<��꺵Ok��w��P����l�C��ћ\;����=N�����;�WZ�6ld���]���:e������h�NxUFk��J�c�'+O�?1�̩ʣZTW��8�w���ƻ��5��+Ԯ��5� �a]����'��]�v�dz�y�erN�m�8�V6[bWg������r�_Ϗ�]΀�ļ����P�����i��/�w{ŉ���^=[���P)+
�#�蒅w�ܼNb<1��Z#Z�;�����u��J�����n�&�ma��VB}]ӽ�hϮ�_�/ً�[7��-�<i�������DK�J�*5�9&��H�ݶ�XY�^���?V���Eyv��:P6��#wuV�W^&�w��xm��;�ro�޺g}�׎�(Ք��O���B`;2nX�|~�� ��v&7�T>Aw��l�ˢ�W��rc64NNJ˺r��>�O=�B.�Q*�-�����uk����o�}bAͥ1���#Q�����/��x׽�.�*�(�!Y;^����S�1cB�{�;+��M]�M�]�n�%tl��/5�:Wx�ޜ�e.���ݞ�*�O;;��}ﺛ�WYy1�vW�xv���T��x���T	�S%jZ�#v���~�����3~�u�缎�L�]�c�7��}O���k�«��+�����h�����Et2��JӣqQ/�v_s�rWS��y�˩q>�k�]l��V^�ܸv����]�=��Y:�����U�,��0w�"�t�=��嗵w\`�b��9�z_��/�U�q����B��2M�y=��]{w}���
yk�DhU�{!{ަ:	C��QIn��b�	AJ�rX���tr��/g�5�no�^�{�|�d$��x3~:�K>y�2�s�.�t �>�&U� k���,����dy�\&�-�Pp����(��f�ن��wTtO{y��&��oiy�Y ������V�8i<D,�"ǽ�t\/�a�~����g�ԫ��RD�W��@Ճ殮������×ڊY������U;^�8�e:i�>�bhejW�I���~;�W
N�(P�]�N�譪�=��O�S��'Q��]e֦�ğ#62Ly��ь.rA~�R���;x�T_?��֥N!�Q��DW�ĽmlO5qƓ����%N���\��`%߾��=w�i$)o?d]�Nt����A�*���}gT�q]xfJ��S-��Z=�^G�{7W�蟪���[UZ��E�r=2s�2�q��X��`��^ǻ�Amx*-}?Z�*��\�E/��ݹ��N�6���vRU��Y��C�g�
+�[�N���!Q�7h�ds�O��
\&�uw�_��]�w�H��;�bNIn��bp7�-;�e�ؗ&r�ۙ�8�kq}�%�����v�6�q�D
�kX���.� �5Ր;�Hmo�Yc��b� �YL;8W���ĝ��%31
��^w��k�VLl6����V�Q�����g#� j�zώ���	X�� I�'|���ܯ>�T�z�nU1�^{�з��8��I���g�^ح���}%�,='=�n��%AO��S#vg�ZcQ�M$��^M��e���6*�o�v��r�V�ʿJYƣ.��+��CpW/K��#@u}���4�Gh﷏���{�<�����xN������8^nϡ�7��"��g��B�c`S�^�lB"�����L�]`�ٕ��-g��m����L���F���Лm���X�Ip�W�J��-�#���j���/5uw���-�f��2+�O~f��Fb5��1���eO�
�ݼ����Aj������wB�m�D��Z�-��+}o����sY]�~�>��{Ff�[��o]w޵K)9߬e{�ҁ��רX��ha�L��Ru�ڣw4��ot���#U���=�-G~���4Ƴ�1Ƚ�U�aho�}g�Q6����n����������{�;�B�B�R>#}jdz��}�3�sk����}�{�9;l����5ALg"�.�y�rޱ1�����xxp�re��o�A1�(՜�E���i�çe��c&���Z��8pS'b@!v�9��<Qq��5�]�`�f}�ݸ����5O8�{;��J��yl]E�]�R��p���v��.8Q�ͳ�5l��cq>���6�0s��.����v�x{ZZ��/r���#�G%�E�-6�lc�s���^���+xϹ۱��b �K�V����x�8�턞�zE�ke�#�JЊ�1
2��b��cI�"k�Ѫ�1�`
I��}硥���L�%�y!��US'�E���~8�_=f�qy��<��K�Sk[xw�{�4a�Ƭű�>��Unpz��,{�\�TY�[u�fg�⬙|'�k?W�V��t]K��f\z���=R���mz/r��]��՞�qT[x	k����Ϭ���Mp��w�+��x���v=�@�Z���t�`ܗ�հ7F��V�;�\�怓yh���D�^�[���i�G�hse{}���N���{(�����q�ކ%n�Oх����ÙwFME�>:7�[$�mc��.L=�k�ݞ\�䂮���Ϥ����N� ~:T����H�
�������K���w�$5�=�mHA�B������o�ޢ���9K���K�zd�vMo����x�-۹k��޻�]CE`��5Ss{�0�3맺EQ�Tٯ	V�i߶�r��+�M�������������[R�xR�~�������!�Έw�d����{�xQ�캈�{�����FǱl�4�̥�����[�[dU�(�K���qߙ=Á=�̉��:p���Uq"�y;�֊�f��s��,{tŎuT��ϳ��b�J_������zN�T��XSb���E�,>ʰ䤀�3'Wmu��r�N����yRn?�
aѵغ4�
���c�b���0� 󺩝�ΠX�!.�wB��Uu]rh��׮�ұ}���v'X6�;N�ƾ�1���[���˩�a��owe���N���W��;��E���5�KG_�wN�����%;F�(�R��Ʒ3����8>{g&@��dGc����븮����1n܍�*m�:!å����x"��"�c�4��;.�V��aİ>2�έ�S0og4&i��ј3�Wo�r�K�F�z��	�O�,wWW�H٪<�f�^ΙԨ�{��WIF������w�!�À�oS`�aDw(hJ�c���C��.����H��v�4��/\l�ge�C�������U���f�'F�Hа��T؈F����`c�#bKٔU��;P|�KK ���5/kM���t���R΍�]�2�5.d��k�μ�[ۼƴis�;Yk4J<��Ü-2�ūN�cS�N��s��N�U��JZ��,�r�:���'io1ҷxີ�3��}e�i�X2�)#;#g
�,D�CV��Vu��}��]ll+2�#Ԝ9C7k�n8u�B�^�)��ts�t��,w�n_L�5��T]�W^,�T��FN��ϻٔ�]N�4¶�h�����=�4�/��}�}�
U॰SK����}���.�(�m���;�j�/P��{�w���r���j�f����z��|,�q�{3��ҥɩ���VUWUP]!5F�6�H@m��x��ks懍��6Nۊ��)�v8�:�'d�T�S��+Ev�眽��]��7ncM���5�6�nn!+Wmͫ��^�W��;0�m�N�1s��R�*��m�t�[��5��\q�;ݺ*-!�,�)뭊;����[Q�<�K��T�O\=��á}��/$a��wg�+��;�;�O,��]8^�/�׆wOF�e�nw&�	�7���;n:]�]j�g�[A�	�v۠�sm[�N����X�j7(�v��9D*q�ݻV�v\=�z��8,�����:���<�+��c��U�W�7��d�O;�v5�;z�N������b�M�T���n�7n�疱�m����v���;A@�L觇�Z���I�������r�C��a�Q��q��K�7 rݟn+]�fxz�KuGA�r��%���ϸ�^��7m�9���w�mێ5v�����d��1��<u���Dc��;n{s�q� �&P��xq�>1���]��;&y�N��ѷ/����u�p�ם�Gkz�룮m^�������=
���2�k<i�x��rq�r����+kJr:؍��]��b�L��^/oZv�s�u֐�[�6ܜ�9r�Oc���Ք�nz��;ZM�.�z����F�d��f{�۞۰rb�,az�v�K�'j8��;k�HH<n3���Nŭ�:*�y������q�i r���n)7�N�/��{���Kp��P<O3Od |ˇ����ۜ�N�۝>���b�*�z�e.���S���Dlk�n��3l�%���3^&�m�7 ۟U��ywd����=5HE͜<=v�q�j��j.�k:����,M��ռw x����m�+�n;1q���Ϸn:��pl�_^��oh��<9T܆fx�ks��t7�i�C=�Z����m�+�x�gpsT��=�淰�n݀ut�t�d�w�[\k���1S��[$��ヱ=�Ok<��>�
���N��uK6枣y�IjեW���mgy�0#��a�\'z�C�H]Z ?�>j>�k�~|O_�5�2ǆ�����
YF�I$�)���dN�t�;;<�pEĝ-u�T)Ļ�t[�����ٹ:�����*��=�ڈ��nq�9�뛻c�˗^���(?J^���k������{��	0Ia�1Q�qt�n,^(���[ݓ���A\7�5+���m�
��[��6�W�!K�|8���,��W���E�E����z�bfǕ�-'�q�ix-cV$ �F��ͽ^s�~�z��x47j���qs�؂+p��ʋ���\�@,]����x�JX��E]�=@�VL�͋�)��l7>�c�텺p��S����{�H��<ʞ�Gd�C�\��>��ްg�� f����~̔���\{���-&TE�./�~[^�+�w�^�L^�{.���r��<{�D�WRׯ}���șʚ/V�<�c�c�6=�1���85���,�N2��}�?IK���p/a�^1�/?
BI�won]}��j4���U��XE��v�ĥ�'���v��^�.	�8����B��h������q�e���&��5P���(A����{����3,���a����bٲ�ٛt�U����y4ڭ������yzB�����ٔ�
�U�7x
�=���ED�^s+&�L<w�b��C�|RH|����1��LS�)�k�_xk�<��[�[�~dx]���x?o��s��|+b�d�:�y���!0�3�/���L�{Y��>��i�K�����Ə���]W�F�{v�Cg�>�~��v�}{E����^)��xU�娐0K9�rK�֞z�n[�2ȿL�MOr�V��]�4�(��4Fi� /�EL�d�ik�9��~2:��<{�i�(��׉"�e��٩k7ݤf��U�P���90�l�����%�퍺H��O⇋l�B~��\�W��Ea��I����䫮�89��:i������,:UW��='�؇a��'}V�����h�G�~���G�'�ߡ����1�^��]e1\=Z`O��XR̯.`�0DuH�0�ATD<�Hn+��Q�#��3�s$�Am�;�
먾�氙垟)[�s�v���EZ��n��Ɛ+�k7Nk;���o�&{��
�uS/���(�ۧ�MS�[�J���=��㈳�g��-��YX��^�@��l�Օ�G��]����iu�x���uS��G��;�Ћi������_Lђ��o�G�W`clZ{�*^�����Ԝ�����7>f�`�n�uaMg�7:�v �Q��u֭�o��&j�ͣS>��[jt&"�U�Z���{5O��q�i׺7�]���7�3�j�F=Sp׎�QRݏ8˦��4��B)��q�<4FH�Wt���GG�y�N�AU��iS%9��[dw�|*q��������}t�'I���\b���c33s�(���OȰM�5gJ�n�!�I��LT�g�φ�2�X�o���ع׎Tz�t%���'=��QG&f`Y绳��ea�7,T�b��M�>u^׽����%��k�
DX��ʕ��j�]sݨ����A荜�uJ��#R0��^�Wg*�m�>�]�r8l� �IC��b �
$���#�{��2�No��'��0ͫn==���0z�����>��&,f[r�ճ���,g����ymP^;=�K�P6}~�4�о��2���}��Kg�lۼ��0cF�	א�n=���I��*"j'^�[����z��5� T�o�kݕޠhX��f���m����P׸=o��eV���х#��D��~sP����z�)W�{TNŉ�e�KY�z.�u//�K��_��"�kۖ�L\h7ŵ��-��J�Y3bF��{Y$�8�׎�>~�i�N8�1?{��Zڷm L�k3�ɒb=OoC�5w���u�-��ZNӖՔҽΏT�]���~ŹS���i�ݩH��³����}~��Cᾧ����\ ^�I��;�Z��CW4g�v��Z��1X�m�x��g���'F:���sqכ\Tg���\���n(���ڲ�r�qn.�M���|�Xć+�8�9��Z��s�q��U�N-��D��:�H�����rgt�v��rk���p��l��ӝ��I\Y�U�p<!�r�뎞S�gq΃�y-\���'i,��0>c��O�ޫ�J����bY��졦 �l93,B��c}y��$Ä�	�~b_�{}i-���ɱ�د>:�
j�K�L+׸Z@����6�B�V+�Te�W�<{���׻{8�������:=/�����3X:�JBi�	C	z@eyÜ��~Ȇ��-/��tO�k�Tu���n'��T8�	��(�,,A)��sh��q���9�c����ݞ���)`�@pu:6�
R��GKe�o چ��x2bԔv����llT�m�D8w�T]E��lM��>��~�k�f�+ê�k�W��W��;�wLA��/��=�t���0$k��r����"�z��	�V@�������ͦ��W �岚�]��^��k�=y���9���㏰QW	�^ǝ�Y¸�
̧�]�杚��?t��ȼ<��I�|S:zm��4�9����%?�J�T���l^�˳�\�#ۺH5"�>Wzꈷ��(���D캤h�_!!�f���I��܁��a�[�BO`,��70��{{!����G��`W]�ݭ��<+�1��a�7�JC���B�f�������MC�yZ4S��#RJ�)�cy�ϪV�d`	%�t���vt����;x�]8ko9��J�v��un�Q��ե��ߛ�r����a�K�h��]���"Ք��[�^z��i~܎7a�d�(}�>ظw��4������L���> �������a �Fج�[��RCPpV�x�fk܋�"�',^�d�=s�BU2��Y��9^��P��wu.�j���}��e��m�p��b�d{+^�[�������ی腻^��>	�W>����k[R��ә�έ�#�"���z��F��BV^5�~I6��p�@C�`RqO}�s00����s����5�����Qj�t�fm������t��G/��?��ƽ�~SB�|�g��(q�ti)+���.��v�υ���z�?�V�f�PVz�$E<w
U!�\9��l'=��ll hE�:��l]'kw(O�	��[�t�#�7�^�m?^���u���RǕbX���hz%�f`�%WJ҅D���Y��,�u��7��پ�6{8�Hǡ�a���Bۍbi�y9n'�\����w�������J�EQUX��]��նn#��Va*�7��:���Q�q�,<�7��������z%�o�`�˟���z&.�mͩ�se��l1@��Ӏ�_��t#�G�n���΍;훌�Iu����ŧ$����w����d�/tl�!�v����%��;�2v ��un?��=~��*9�x��D�pRp��
��:��㟁ܜ17����U�`V�_ԫna�6�7�7����"�ڌ��g�l���8��������qy��E
ؚ�y��`𫂴��¢��T�/=���naO>�Ȧ�s[��t^��՟�s�2`ɩqZ	����~�"�ǥ&oq���F�Y7�fm�����G�կ$��k�����r��U恗��[b��=<̐���u�u26�{�s��l��k�p�n`8�ّ��m
���Z�@�đ��ד$NdL���"{�.<C{ݘ���r��F%��k��;1Q+n�,{=R��J����4zࡗ틇1�a��o�����N���I&�>��ڗow� ��CM߯�}�W�f���Y�B!�Y�Q�D�X5��4ۊ�V��n�E
�j����s�w���dK�"*����阔f���Lf{�Dj�^��fJ���*�ø��;[�γnίft2Oȕ�����c۬���-�����t��ު�e�X>̆�Z�kC��]�:����䅕Ni����ܬӆ�CN�=��o��J��`B�'�Z�x��=)]7J�����f^n6�ڛp��!�rf,j뽇������8��u}�\g��c^i�b���/yc�ɛ7��Mr��Z����Nu���;���L0`
��zn�p-:��J^�����3�O%;��;3�uQ��PE �ay��qO�����ixk�Im{u\�eK�}W;텺a�5�%�z�`�{=����D�:pNۚ���Ԕx4Jm�i�1�Of�=�?Z5��r�Ѭ��* �����}(�\�R��VP�Mu ��6�����������&�k]}�'c�C-��P���b��8
��S��������#��>�Fŀq��ۢ{�+7[E��W�Ku�.�l���L�F�<���8�ѡ���>>����`f�>Y�/��N�X�y.���d��Os7�_���&CMlPw�U������|C	��Z{ާ�W^:��
�:�^/5^�Z`n-̯*>^P�����k�d~��WQ�6Uƻ~s"C��ۙ�ѡ��J>.��3k�b)�n{(d�빉_��O9�n�8:u��8&��㗘�62�
�w���n�N��6�e�W��hI��*���hO
�� �s3ڱw���h�P9'T�bWi{G��S�!�Ȫ���9���'KNe��fM�.&$�ݍ�0��M���Q`�-S�l�ݨh��}�[}��U���fr���^L���:ڍ��G�*`���m��Y�Ip��nէ���1{gͨ��99�<q�����Z[�T�n��Jn-B���tu��[��U�^�&�72`}K��6�S>�rZ�\Ι�'u����*�b�y��g{5r&v�;;�okk��6;�����k�k��#���q��ܛ��ݹ̧;���EGX��^xD�D��kݷ�8+u����y��?I�K}4_��y�XVwc)M^5�M2_�li�u�SMF��&Y�=��,���Э�/��:���\{Sn�bu�Դo<��ث��@�yb˕�^N��=��碌�7Ͻ�?�JE%�U:(\��"'T��F螮��u�=��B��j�m��=Y�N�ݙa�-%8ͩ�X�O5�)(P�%�tg��]���a�2�Hj��Rb���b�5Ϫ�WV8���Q[q�=�@˔EV����|D*�ҴC��`��N�zMV*�\n}9����p:����𹸌��ê2a ��r����V�<��粏zO���*�on)� �1[�U���י7`�����h����1J$ˑ��t�����,�r���(�Y��p�oaK�=y|ߵd�Vxn�n�8�;
�k��9�� t)�U#q�^��#tx�� �p��	�u�P/̜s]n�����63ݱ�����h�铞j�\B��lO�G��u2j<yb�с��{,����W[�\��4��v�I��M �(	ÆTʎ�}Z��G�y.�?+�y�[SD��ꖨ喝q�u�+��%*Ԕp�J�Λۺ�#���1b2��o@�2g5�~/y���^��]��}�09� ښMIt�M���ͤ8^	\(�/�K�{S:��j�!��5ޥ�W�g�7�״`d#9�^fⅽz^$�!4!od�P�R����Ӽ!�wvK�c��%X��`	�_;����6�y�A�Q
�R�����:^�e�I�we[#��U�ɼ�$�2�d� �����u׽��n���#�/E�w���14Pg�#��s-���z8���z�2eO�	�;���`ȼ���xpD �p�QQ��B�W^i��W��Y=�V.f{bH����)���wa�P�c�!��7���g�W�qN�f�1;K�d�I���S��3����#zW�<�w��zu��{p0�&lL��T�:+ˡ�B�Ɗ���3�!֋5�.���?W�T�RE��t#;@� �pp��-\z/5�ͅS3;���9O�l��ĥ ��ם�:�!A��F���'{,Y6�����o�R%�E@�a���*gnE��JQ��W+s7�&�@�U�T���T{����a�A���yjv���
�\�G�"G"��38�V����d��9ղ��e�'9��i̯Qpʌ�[��ڜ��(>pRI��S�8Ǖ0ב1P�*�~�SFG��@�u�R�K����� 5�ny:��1����s���Ƿm�$L�����p��uf���1�bYI�k�8��<���3͇Dڭ� O��OL�N^��Q�'�XY_BP8'�V�ҋ{�Ӄ@���^�t\Զ�f�kܷ���B�:�����-Wh}�q}�vٹx�3�F{V�⼏0<�1�lN��:��"�N`أQ��8��߉�u�3D�������o.ו̗&\U�{�-5q��ʉ�l�O�UͲtȉ��Ū��q���HYl�P�N`ݴ���V�\*&���dҶe��EV��.T.���v&�����5^S�%c�Q��;a\������df�Ǒ䏚%6+�R|c��@����\wn�z��[�7�WT����&#��>����э�o��j\2f^Wg9���
��%y���u�F�^�id0c����e�H�Ϗ��(?���T�QS걡F�Ǝh���<�7�B^/2M�u�#�w�Q���t�8�&�gEK�(��Ƣ��Y8)�u:䞘2�����a�f9�K��=^�P��=�e������0�E�P/O���D�U�kS@�=�OT��f�2C�޲)@�N6	�'&ZU\�\rV�i\�׮9�nZ)0#(�A���¯�Vܸ�o��N��H�,,�~�ۑU�ӨB�O�Be�>dU�ȥ�qJ��+]~4q��� 0l��XǵS�aHו�/Ƕw%��B�k���O`�b�:�o*7��]���@-L���uJ�ɘ�J̅�q������;�=b='�$-~�US�U�DoX���ĐS,����'��4S���U?}���Y�z%Tɼ��x��;�����
�(���6��d�y��CϞ<�B���{���&G 2���T��6b�\(�#�o����(����.Ʈ����ڲU�][I؅�\R���Iv��q4��V<ݩut��7��2��}ò���)�onIu���B�F�����]`X�AML��)���	*֕YZ*M�.�}�u�zw��,72d�# ��&$���QQ�7�ui��)���R��9�E��u!�bŉ�9zw*�@��\;*s�u�Bh<�ӕ�X��0�+�Y���n�
�P=(�xVf��oSG-y�N��yn^�8�[���C���ḵ���'[��|j���mJ�R�i1U鋩*�՗y�qz�/��ŋ峵��s�xRƶ��M�m�' �w�r��������6`9A����F�P�l��k�z�'b�<��x2�-U7r�=��6�����J��ܬ��K��@T��yW1��ҬrkAP$��V��P�c4w_A����K]�<��Ycu��ԭn�E�_I�&+�[;2
ڸ{����4�}�f+ֻ�����v�z� 01�9oӲ5n��=���C��'\ǝC+M�Tk���Z���B��ʹ�����1>�k��}���n�ul���xt�@b9D����Y���x�wmM62jxL�Ʊ��aԡ+�Y[5�����3�Z.RS�t�d�8�>�o�f�L����A�mِ7&W�:�Y�1P`xN;��jp�����<�������u1�]���7b�9���P���VTl��,Ը`SV2�/B�p#�#%s��B��؍�w5�ft���_z�(�{<<Zi�Ȃ�h�UКi|9��Q�#�꽓��-v�扡�	X(Kg�ĩ�3��+�_��ˣ�l���G�Q�l�1ƚ[X�D�uk
o4��h@	2I�s��<h�,M�����h����Mi�ϐ�\��0�&�v��q��B�W����vT�vw�-�f�f�}2�:����M�t,5O���k��]�. )�X^f����ҶYY���PT;�l{�]�7b3�	�.�R��A;�s�4�dK#飷�y��Sm[SbtD�c���,֬�����ߤ��B�W�z6v��Km ��\����;[��Q���T���+O��cw��$���T���my%���_�>=;H��x,,ɮ��;$����,[��=��E/����\Nz*����VV�ONϺ�ڒ�ln���]�!�e\��W��K7��"C�J��J��Y-��S.A��g�٧J��<����5<��l��X�V	6V��B��O�Nwn=s�gI���-]4n�Q�6�1����{q�z\�p��N��b�|�]�8�7��A�ģ,��:�U_SY����Eu�:b�Y�
q(^�\���ev=P���[|�ޡ}Q�V�;%�_-1���9�7n�3WR��j�$�-���%m8��-�e���s�(u�=�k��i��:� <�p���'���kVz�vx�;=g�'�=�^{q��Zq��%�1�'�]��s�znt���ݣ��Dz��<�EBL*x��f����IJ�NS4[G\���tq�)�p�8��q8��Rg��W������s�K�X����sr�8ݞ�����x㸋i��vڶN�go-Ǯ���r�7S�!ve%t$��h����75 �^�Q-7���j�U�&����%��Ƞ�A���%�`��G^�T�`r����)�����n��X�R������Y�m�1��k��W΃{[��Ȥ�ӳ�H�!��RLVK��D�s�\��ނx� �* �mݮ~��L k7nբ�Hr9�Z�i>�b�m\@	����z����xgSZ���:�.���h�4lOl�p���|�{lb�릈c8���wy���U�]��غ�v�ץ�w�Б�'Ϡ��o�w��|wp��i�w���*#���w$�i&�� j�^�M(X��\ɺ[��}�����=�6�=^
,�:�ni�JXu���-g�*N�ѓ� 8M��JG>̹̎�RK�mCP�c�Ea�s��z��2��8��FC�����l|���=;;F��oo�.�O�˚��_<���*2�F��9:��0[ݺ���Ó!�	�m���[��ף�^�7�w��^��$�3�����2�8�����y]3n�+2ص����Μ���deYl5,'��^츜�� �qd@LY$Uh۽���P�fq��緺�:T�I�M,�Ι��<HQpV��E�w�×m�&U^�AJ���C	�{6�U���8�.U��t��ɺ3T*��/��;������v��l�W�xrWhB��5$��YO�~�i���wǆC�p;{�fW��;�� �(��'�g'��;��S9t�qS�}7R�N�E��<`~�0.�ʄ�Gn��z,{[��i�ӣ�����z�v������}�~=���L#��� "l�`�����C��ۊ.'s�նulvH��
���l�H�t���fH���L��Υ�f�ޭb��l�g}��8`[u\��˞I����LW���X���Os��e���#�S�� ���u�&���i����CE&`��j/��Y��ߤ��5U�K�U�k!��r���Ω�k]��#\�m�o�2J&t��s7�iϣѸ�L�Me�fC��z�5��e�y������'�F�)�KK�̩�ƹ���Yk�����^������{T^����B��a�q� Dz9+,]�݆@�<6�RGy\�鷰29Gr �I&�i�d׽�6���;�]li��>��8*�Ysx�v�"���4cN#۫���1���l�|HH.R5}8곞�'r%uѓ9�_�t��k��>�j���8,�����	�����n�#�?t�|�nz��;W��bv��g���U�hʙ�Y�gc�nNx��l�N{^K��cLP��Ħ_Lիm���T�G����Y%�}4��_��^��x�z:0���)�u�+���S|���*ԛ�}\ee�����|)K���8���+;w�;'V����e��{�M36mXZ��Ӻb���ž�䬄����v�W'��X�SXk��1#�F)�5.8���^�@Ǝ�wX�Ygovsz_�z��3}'sn,MJ�/l�ע(C�5�%���Rg}�s�h���ezWe����]�+��~m:i����l�U3k��O�x�/1tk�E%���eF���bs�F���7�W�4��!�͡�}5��Q+�{�����7M�5�g(MO��@^z�e>}X�����g{���wq�-��9��]�G]��ͦ�]=Q��Ux��Z=��w}�����paAP�h��No��c� ��П�c��s����:��&O*��TO*����B������F�%ne�UA�D�ĉ�Ml
���A]��[�y���i�*���ζ\��(�@��pT4گ}��vNx�x���S��L��d��|9X�Q~�/o�'�2�1���l��k�s�� g[5���ܓ��"�>!���z�����ی�ixy{Lܷ+�K,�6{RH��Ș��D\g(�
ĉ�nm6��ȏr�Ÿ�������C`�R�9J���=Eo�������w�s}z�wZ:�S�ǣ��ڠt��5��3�\qT�T��cc�:��9�3�T��y�6�{�9�HE��V�8���9���|�p}��]����+�ۡ�{�U�9w4ɦ�ͺepː������2�Kd{��x�Ro4���B~�%��A�7C�d�6L{�Ȼ��w/]R�:�$Kέ�rgY�c�l��k��b�캩���!
e.�$o��lӺ����˗[�����μa�{��^M��Q��5u�%�.3���i����!ل_l�_ ���»�Ə�d��^	�0;�Ђ7�I�����)���QAR�7�|�k�1M\�[�3j=��Ȧ�Ձ�Amֶ��c~������^;��}f��'��j"/ћ�<
)��Ǐ�Î���{7=j#�G��$�Q.�v����~��')P�6Yk�����q�������=�۴�� 4ϊ`��>G���5�ߧ��@�5�7c;5�}��O�x�Qs�z4U_A���^ʉ� �̸��>}���!�2�8HX}
��'�*��ϲtG��9���Ѣ@�#N˻��:�6�>��j:62�R�7�=,���3G����蹭�w;���K@�@;����XP'���Xv|-�Y0j�o�\���ɝ�s^�WG��.܉2l��'<r�4u׳��v����Uåb��%�N����ӧ�2D%�`lp�P$�tNm�V���騡j�J{;q�(��X��5]�@h������;F(��O>Îl}k@0[��#���Ѷ^�Z�fl�:<R�,6����d��̽��b;���y��>�V�vy7:`:����˻o��u����v�^��-9�lrR<�j��s�H�&q��ش�Ի�I�4A�m�v:1�놎�-��P�t>���oX�Ɨ#�vXHA�֜�!��v�;V���Q�v�#λ���=[nvˍ�.+��8᪂�fU60f<�M��re�ٕ����7B�Ν�#�q�jCr��v����p�6l��;=(��[��r���{FK���.������&���cB���������$&�,�:��7G��j�%��"v2�j֘���N��&zmtז�Dj��T��;�D��h�g�ŉ� �Vo6�u���ܥ27JB�ϰ��vc;��������	�j1q������8�'�}�Xe`&R��,�h���po,��(-���h�ׁ�X8�e��vRN2�<r���I;�ˡ	�����8��_+��)<X��I3�vWqs]����Ru𸚍��Ҳ=�Ot�P	�j��o������͟/��Oa�P�=�7x�����ԣ�e�eb�vw��7��=R��m������ v)�P8j�O��7~>

h&�{I�3r���*�/)��y9��]ָ[���fHT�Ro����A���&�-��B^S]B�������*k�<��Mzh���<R%��>WV���Y��co+iɈ�=���e+�yyKu�;U*��˶l؇�s�Pҋ��˙�e4�rq����L�|��*٘�g9+��qH^�`�b��<��1�ϕ���Q���[O�4�fڎ��\=9���1��]�p��Q�I���Q'�cc�����1�%���6U���}��Pn4}{,i�A[��q����Q�W.�nnc�yvȷ9�'�4�g��8��#�꽓��m�Q���i��}*��	E�C���*�t{7�	���z�=�p2�F�:��=���B����[����w[)"v�2F��Y,���L�ٶ{v��P��l�m���b���D+�{|��~�g.��v)�܉鴪ⷔF�XMO�oU^܌���"�3]q"8���,���N�����( $a��?q�^�=W6�n�d�^7ą���7�ݣ�O�Ǒ�ZV��t�Gb" ��v6��{ �˰ϫ_'xdR�G�������b���"����G��B�[�pq��y*�^�uz�f�g�t$��Uחc1�ǜΨ��g��uޑ�p:"�-K{K�ݹ��y��m�ߘ��~�5,�Z��i6\�S��$	���)F��2��k��6"�ߠ�5�	\^�u;g��������{1�Y����I��>
��g��h��� î!�v�jɽ��s��.u�lWӌ�RvL����崵�4M��_�s�)Wu�<xK2rZл}��j���}�����h� J�]L͋3�wLҋ*����>��Nǻ����9�K�lx�	&J&�-9�,�	7j���D�Ϗ�i?�E5��n�oL�]4�R���<o�$����8W�_7���gx�D������;�Be)Q���r��Aú�6����YU��s�EN����7�x�7
[�����]���]3�t�Wi̐˫�EV���ݜ�j- ���6oƵ��w�ˉ���B,��2'{�dB<h��8��y��SxL_���K"NڲI���[6����Q��V'�Z�v�ِ#c��D�)�\v�*͏Sy.ae�/��FD��D������`�$Q�ٌ���^)Zx!��vv�$� NKW�֓57��8OL܏3�{ԑD6jE�-r�8ț�;���u%ȃS	��+���ȩ�'8k�q1w���fME4��lS�׊�|��9���ky�%�K4����v_w��6�,�Ɇ�͑-��ySb�*v�/f�,�z�n��Ѣn�3�z�(��VTm���"y���./��鱦�P}��^�V���ڳ�+ ׋Fv[p9ۻ�&g���G�npI�w;&ωUW��������"U�Zq��+v�Ѹ�>�<]e�,�۶��q��9��P'�Z�y�G�c0�8pJ�`\��~.��M��|C9{%�z����r�]�⭋���:6	��{'A ��dl=]f�i�t5�]Eӥ�#��
�^u��u�*eT0ꂖ��7�Y�FqS]}�l��92�5�d��Y�.xo���� ��#/̧9���=w�G�M?cU�Ԥ�ۿ�a��l�^�r��.51l=��Y&�Z-�o!J�j�2�}�{��t�ݝ}�&b��R}�P��+�C�g�/����2�Qڢ�&��=Փ#b@�h�~Dlֺ[9s̮u���b�XX�L	7�q3���E����z��Q���eB���.�@�n{9L���B�혆�F���=����������o��w�C��"*�B��9�ʼU�~��x�O���5H��Bڦ73,+:�j5�n���z�����]U�b�k����$�^�fb��2^խ�ԓ���s�-�
%!�]�i����TD4�2��걄�1��BvɪEH�޴fZ�:��s�V|��j�Xێ���1:N�i��ݰ+D�[���4�D8��Ӣ�9����?��߿�uˍm �_�Wzk�U�f��t���l����ܮ����]��ķr9�M��u�� ÆB,�P5���z�K�_M�t���RKB�g�յ"�!��F7�����_�G=�!�s"ϼ��>���Gj˪ z����ۇ=��%���l1�@u�C��m��s{R7�jj����@b�y�0��W\��#�=��徽��'���W��ZS�
+f9Pվ�Y1�`����SY[k�+z���B��J*dR�2���$�B�pu��<M�mU[������/��0�cW�+�k�X�U蛹wX7n$+m��9�n��f��J�J�Z��)�l=��u�9Q�4ĘA���[i$ঁe�y8��Jtv�{Y6�����������9��F��;k R;��/\r ��4��5�t�Z���f2�,byB8�����cd��g��ݸ{�^
��6{C��.z��g�]m�KX�s����ڴ��uF�[�v9�!�)�����n^w7:�I�Uݑ=����,�����gf�vܽ��(�i�[0`��PQd�My���[�˜�<�]�Ϊ�ۊQ}�w�7=3֘�WWWywV������y�>E�IbŞ�ֳ���'sy�3һU� �e��/&<�M8Y��F3HZ��EC�\�'���0׬�&��������b�^XZ+�������G0a��d0�@�}��@*sv�����;5AuNğv)���;�5<��3�X�A��[gӻ��K��WV�7��6I)����)a�z.���6L���nP�Pӑz���s�T�G�0�аX�\9t0s�+������]}wBi!0,��g�Zk%[_=��t�Q��B�K ��q�f��΃�ŨW-�s�L#�j�古�-`^�S�c��P荸�}<g;��r��[i�s#jw���ѝ790Y�Ñ�3$h�9)�ne�~g�d�\O��P��=�a�5]��Y�+�hߪ!�/�Ҝ�9~�<	�A7�\a.��3W��^��c�H�@tR�&q��|^n_e�K��5�z���ioD��=N
���\�-�Lʃ�P�Nz����[)"[�����u���'�,���=��Xsg9G����	<����)M۬��k=��%�J��B�\�w_�a8�K��t7j�MV�}����ٯ$�nM��=��Y���>9�,ށH
(���E�};M��׮�qb|]�s����+�ݡ{��-��0~�k��1;��Ƈ���1�E���\F�7@�DpK���t�*&���V$'@��C�t&�h_o���(��Xv�ٔ.�+D���T�KHQ��*�<�2����ݳZZ�ڷ5n�Edyvy��u
OFe�ov��j�_5N�k�-Y����A�kE5��U��a1�}N��������Bu�سq�ٛ����|y��v.3f�-�d�2�x��R.a�p�����B��)��AU�e��35��D2�ƳH#7T�7uq
r[s/�mf-ןKqRP��ϷYF8᫵��Αwe����NP��&��WvPZ����ؚ�����>ˮ�u�.�5f��{IV����i��fF��+�rg����zEK�{�pq����'d�U�+&���Sv�����61��O��b�wp|77E�gL�f:,Y=]��of������9���)�`�#i:�M�}�p��r����,�l*�J��RT���.L�ł��M�M�feF��t��f�wG��lW4��X�}���3�9�]n�iU1#�U��*�3E;�H�n�2Y%e�i�'nwtx!\m-N�RɻǢl���h�v���;�*M�\��Ø��#T��'�gCqv��{iۦ�`��;�j�Ȯd������Xu�"��j�Uh��X���]@T�m����� ���#�R��R;/�7(��[vP�,�ݺ�u��ݦ;c�p�o8�oCk̈́�콯mp n����v�=q�<�ζ�:�ȡ:���%���'�l�.�;'b�ǵ�ǫt��+]�F+�rmO����wnv��0�v�W�Qm�x=�z88��R�9v{�6�.���,��'�ٞ��̱�m���ܵ���4۷�	b��ɓ�v�, �]��ckp�/S8z�.�� TA�RWhԹ�n��2J�� �l7XS�=o.���:�{]�s��pG�����|7_7�Qp�S�g�-�����n�j` {n��=�i �:�s����m�s��Z6��#��t��g"�=7��Ȋ&��ɲiC��ڸ�k���u���T�ͦܞѫ�X�]l	�..^r�d�]����;t�qc���2>�����!y+��s����m�Rr��Q�7r^��4��5ہϵr�x9�T۳ss�Λ�׻W>�om���Vy�<��nv/:�Z�u�H8wS��u��d�޽�N�� ���݅I�FB*����g�v\�l�t��OA�D�<�ml@e�����c�v��>j��d<r���7q��g�\�vM���Hvh"6"貚��E��<��/�v�v1g\z��n��Y`�����9H�S�X�z7,��r��cc<ZH;�O(v^�����=��t���P���O+�꺩��6�����\(&�����Ռl����lIq��<���Wj�{ynV��r�t/]�Ì^Ս�nZ�7C��q,� �x��خ���^�\6�͎�^�Ξ�q��*�!ܻ�^���;��<a�s'��s-*�n�W�cZ_klfx%9����n����n"�c�\;b�u�՛n��8��5;f+���/ ��.ʠ��vlkv�����q����ۉ�խ)��k��]m��<Rg��n�u<v�ӋuoI��v���,	�� �y۞i|�ܚHݺ�3b:�����I4[�.l�0��{c�N��\��YQ����2�i�Pv���<Ia�Hi'<�U�'MX���8�v\��Vq�D�	����$�H��H���G2���'��۲��vu��G�YR�"(X�Q���>�x�Tt�o�>1K��C �h��Y����æ�*x��G�����gݣ�Et L#�+�sqP��n�`ϩAЬ2%�D�ku"�sX���FvC=S+���.�L����弳U��m��ٵYD�Vڮ5;/�t����֟��J6蝧��ek�R[���o�u��;��w�����U��D�l�	��i�Mr�ǯ��`k���B� ���F��{��y�}1;�}!�Ǝ�%�$@h6�_��Ļ
�zEx^Ƙ�2l*��S�C&oEG�`<�2�z�빊+�S�`b�ʋ*��@�7Tƪs���7�4"[����T��6���A��\���^�/ç��L-����2�mnT�f�͈���ryzU�����>��S��g�$N;/gq�el��5������!�3r�E�1[��]��iP;���!]��O@�a�i�s�r��}�9ޗ�m��v �f����y���i��t�oOS��l�&���b�{���>�u�z����e<��f0���޺�L�r<.�����g�S�s��':�G�n�Ѣ��6�5wf�y���v5ز�ڋ>�_hJ�£�#���l�y�B����������K!�\���醜hܘ-
����vmL��f`^[]�8��"0V�}�ri+�i�$���G]G}\s�	�h ʘgp��S����B��>	M��r����M���:��H�Q���3��Y����z+��r(�T={�x���������~A��l�4�^+���y7k�Dd�RR��u����Q}��d-���F��b��#�@���'�ټ�'�*��2Ś�v�hb�z%\\�G��uJ-V��	��[�=3'b�|,������+���`7���I׽��χ��y9R���i�H��R7���}i�I�vO����D�-���C;x����a�����9ִ;/%魶���3 �a︩���T��BS��v�/cgtH�
��՝�v�(7V{������[y�ܞ�9����ju��N����p����������~_�꒺��L:�s/w�3Y� ���ݺ���z�t�`�<�M�ӽ�r�1���a�6FD����2�b���#�s��]����(a]7]u8g3}|�>6h*s�k\�[o�*������]�k�3lܱy�tN6��*L������5\��EړƚȒ�6�po
�"c�Z�.�Q�K�PT�mVf�)gk�1�����v����{!PfwUz50���C�~쫶�DA�������Gv��]��=�8F\&���^����2�XNH�Xtף�Qθ]o���*���nz$��uι�#�<���n^�ƶ����0����2;`�3��F��Z�!�ĩ��`�Z��i��~aL$mc���j[j�f ���+�*E�����<�6UN$N\'���Nџ],�	��~���؎���8�.�*�d{:gf6i��$��7��^U�T*3E'�5�D�/s|��7�Շ�bh'�Rj ^f�6qng��`2�`����(J�M4�0��0
��vM��J����Dg;��^/c�j�utM��o��/9?{�`̞~֤�I92:�g/L_v
<C`2�A���"=�E�~�3c�>6'Na�ܮ���H��Χܮ�/�!���9ʹ7- wU(�Qg<����Q�Ȏ}��sA�!_��d�o�@�����>��c�f��z������V�*��Lj�X%��\f��O�xt���1:�Ҁ��[�����&�pxO�~$4������ɘ;�|�r`*�hdnw�X��e{�G�Զ��+���m��`J��� �*݉k�ߖ:V'�)�T_L�Ğ=b���m��K�6XN����Nm[�o��9��Y���p�Z�U����\���"*=t�5��9��vꮛV�;����k�ӻu�b9ͷ<k�K�n#+�	����ې{jq�[���[��XF�39��0���nkԡ�^Q���5Z�vި`:h���Q3\r�ݺ�[b��v��NJ�iۮqm�A{^�n1�L� �q��ݞspgF�{t�����lg��W@�F䍞`F��:�������>_W��g� eb�y-���A�l���ؚ���Y��.�ӌ�>�$0\7 h��F�)�61�F]w�qh���#����`�xN��l��sq�����7F5��t��B��	��y������r���{gN.�M��;��W1}�B���I���jU�ʳQ�nw
'<�_�������mX��Q�2��f���;:Fl͜�n�va6�l�`��,�>F{�M�o�s��R�]�'%C\o��"|m:�WNk�mA�c*mZ�RX��W�5�Q)�G�o��|�J��湜ڃ�A�7�nߚ��92�<5\�*q�LQ�w3~�Ԩ5�ifKmn����?)ٻ�ok���D�pL�k1�O8�˲���_y��Wڔx`�z6����60:�pv��4mR�n�fT����a�{�TM��@ �\�ٿz#�2l@&��۔M-㾽�zj,�JZ1���	�'�d�ӊ�Iog2k���tB�F��bц�L��;	_!�{���%$5x&I~M�R��Iء�~��Y�ћ<����.	&uLR]��Ej���;3�y޴�����2���O���}H*�SR���^�9�(���ϺC�X�����*\��Fq;n���+v��w7�u��J,�f�T���M�Q{���1�s���]7�g����	(e�
\7�+K�͹�ܞ�7כ�9Vh܌//���� V���3:Y�\���u-;��u���T�V�M�E
ٓ�ߏ���rt�k���z�&74Ù��`3�{Z}�@A�ʼ�I�����u�H���K�D�j��4ѣ�I���ӛt�S�܈��F�#$u��~ZD�c�܃�t(�o
@f��f�r�M�rQr&�N�W��=�p��O$z$�8-�}'��C����5��Czo2�-ROz��R07���s���_1F�(/۫�&ڃ��]o�+:U�0�&o��x#[�X�}�z��j���tp��ՙ�uA�=��k��阩8�7������"��W��G���ڛ'��UǴ�y�A7��U��2�Ws3�~��o�����(�Ң��\m��f/#Ul�i께�j�=y����9[՞ڗ�KqS�{W�j��9� Lt�+�2o/;b��۞��yj-K�V�B=�d����/? 2y'�`Ƴ��3[�~�§���^}�Y��܋1����&bM�څ�Z�����è��e�O�����c��kho���`��4xe��T�Mz����`E9�Ct4'_}ި���C˽�1�9�Ah�
8d�O5���?��%��)���c�Մa�Ozg>B1ǖ�Z:�Vf��\")���L���F�)x��C!��Ϫi�:�c�֩�Eւ- W����W���&��89>�A�F��r��,3i���r:S#
�|5>�ȸu�#7������$���Fi�V�w�*��^�u7��L��Uq�r����HD9ђ��T��sZ���>""����أ��D��
�^�U]���O5�I0�L(N!�I�x]��'�����&�z)C9��f��]B����d$�����\j��0�0&�Eں����q�g���D�Y�$���<�h�6�l
(�O�V����C���m's �2u�#��Ҧ/ 84�Ѻ%F��X�欉]�������M��Xq�;���ħȳ�5�sq���@��	Fz	p�\�9�.�̕����+׷1Sq%�b a��\�i7�h��͖�N�l�՛��na��K��3>i]��ݑgJ��tǰ�Uu�To��ʊ�����&�W(c�A������^��v^n�>�� � 6W�K���cMEɓ|�9��Ex��R��'W��d�Z�-�lK��O�6#E5�ǲ�b|&�� �+�α9����7$��Ҝ{#G�� �H��b���N)7q9�[^EӅ/p��窡�Ɔ�z�Y�z��B��\(9�|�M�"&�әA�+Y���dx��1Y�@<��6��ZH��j�o{��:�Y���ww�v8��f{Ժ��z2,[ l���{�vcMy�n�M�xi��t��<Ձց��ϣ�� �e�qHV����Ur����xu�gc��8Q��uh%h����f�kX2<p-��*Y2kT�*ᘭ7F��OLM+�x���L�VL�܃W�u黰sa��Y�1WV#�"���.-U>��=�j2�9�"]���lV����z��mM����m��ˬ�����~�D6~F@ͯ���O1DE�Lᱱ�����{�>��{])��4��֧�Ű���r�ˑ's==srlx?4���#bV��2�i좎��U�)��F����;6w4�c���u����;�Yda:�`��l��U&�͖�'5��u3�/f}o��Y�͉��V)���e�l��܊�]&g�΄��-'�cZ�Kg����\�&=ೊ!��Y~,"L���V&v��Ɏ͙5��_r�x}RY1��u�Y#��;�Yq-�}nǠ�q4M��*�eo>���q����+Y9|��|��O(`Bp�,g)�F'�-�ʝ�%a�; �^&{r�n���;�*�v$���F�&R��b�p�``X�d�1�ι�Uk]t�+���v������مr������VL��~�v�ߟ�UqtR�G>����#�i=�v�]4h.1��0�I�O`�ݻ^��Cݭ�C�A�n�F�zx��'��*t�۶Ln�[���ђy����d)ǜ��<1�vճ��v��(e�b�ܽ��uI����z��A�m�z�@�v���cy5j�E�ۗ��ʭ�-@[{9�v��u��]gs�q��z˻9�ʵ����mm�u��TdB/�Z�q�>資�A�ELLhn���ܤPn��1���q�2He��J��	��]��-[���ّ�N]�U�2��5~4٨��Ǫ,���5F���j�~�C+חv�L~��]�؞f��UQRؼ�~���}-ߠ	>� 	�UB��Uf��ܼ�l�ڑ�œ0k�� o2J�~߽����	!<.\;���=��{n1��2�	��PX$�=ѽ�c�/l���v|*�֦�u7� �&Y�l��M���]���gA�q�fj��:�'#?���M}���㫪�<.��t�=W��H^j�<���KSaFsI�[i�qR0X�y���sL9�!
�R{&�o����B`�M�ݒG	Cyܻk��^]�m�%�zn����(�'��:/iA�Ǎ��<�c�� {p��ݎ��b�u�ܯ��.CVwIʬ{gb�O����'�1ɦ�e&`��9�t��7GU#��^�oj�c�t�VA[+eFy{��P���~���C�j�5Ɏ����车�U�2��Es���6��e��0���5	����1���f�O#þ�]�4c:��1Ppw��c��oط�+�pv��`��g�J���C2��/Z�[�u���J�["��Wo�/�sӝw-��P]���ST��a����fRkw3���Ӻ3��许z�w#�`'U���!�ӆ�� ��M���/.�n<�Uｮ����
��W��Сe��(i�g,���X�cs�[v�[�nd�m�A[Zs�����}h��R���Z,d����=m�C�8,���и�SZ�ی��D"�</+_:yjY�����a��$���x�a�7E"��G���Bn_	Q�q�|�$fA�bs��{`C��~@�W=�6|ݲ=�:��n0ox��`%��.��d��"�ዅ]���:���V�s,(w.H��B�z}y������� �;}Z`VF蘞�S�`_�qj�����/��2��ne����i�H���E-��[��K��ݕ����eS��g� ݦ���N�L���*�E!�omW�I�䨞���P�@!�б	����w{Iܭ�����ܵbM�	��>�\H���{�C�v��f�"������H��9�&a�s�*�^$��1��)u�������~B���$�X[�"oW�n���D�&6a�{�v����QB))c��U���TL�z��d)�6��܇X5kN����I�W����n��eݗ�Z��ڀ0	-�"vt�e@�5j�(����3{_,ߥ�&m-�7{[�90vţ��V>=Y��.��:Tm�/�g}����=�>�r���V��\�>v9!�g_59�&�y�������m��
nr=�]�
L��8@�|�'�B�Q{U�:�P|�v�4���d��yұ=75�6�ڭ�\d��GGBF�%�P�6�X,��%�kD���6n٭͹/UT;��q�{"����]0��㓪��py�ע����n&wd��`�y�p�Փ��J���QI~�9�Я53Z6�+1�+��5o��LF�[?u]3��՗{I�,d�Z )Ƚ��a}�'���\)��D�|3~#����G}x%�:�*1�FL��y��Y�:���qT�^�a�ϲ^=��x��2����O�����d-��h~	�c�aXd� �-R�h�;٩�Qh�dau�[���d��2��Ɔ�����sAo���E���������a������TU0q�aތ"i��mͮ8A@B��_a1����z]r��TvT���p��>>�;ؗAc�ʥ����>^ �ÿNa�͟J�wS  QM H�&�%'-����S81p�f��pozo��V���b��v�eG
i�J�
�C�gh���p]��]�L��q{U���P��D�\8�����m�Սw�L类q�df�l�m~<rWT�{l��"v���7�2�%ɜ:찀�M����H��Qnt���L�{zI��v��/���T2��9�#��)I�����ү��`�-��on�l;��^`�`�;B#{�ӈ�e�S�u�J�ۘ^m����aT���%ڗ��aъ��W:�����V���sj�;r�U�Ѯ�yu�eo.��Gk �bֺ5�K1�,��<����w+�%>	l��tEGصR6�S�R��F���rS%<�k���]w^M��6iѝ9R��M�3N��5���v�j첤$f�Č[���flkp![���{/�3��ۭ��,*�iW�|�V������2�d��0Gv��_�sγ����&�sʙX�Rd����5��:�]_6��U�ÝeL��Yr�U$�v؀�'e}0o4�5G�7 ��mf2!�����"���x��G�W˫��N�%=.��w��Nͫ�^����vβ�5>B��ꕁ���n��h�yQR���Ϸ��o2t�v
C�NN���L�n�9�iT��C���IX7�m�X���7It��Z.
�{�5-]C}�r�/kl]�G���ŕݖ\p� O+����-$��Vr�t�
3��s�1�kE��O {X1���t��,�Q���/�@P��ݕ�����u�ia�^���Z�wcK+8)jCYC.�*2��B���v�FT�ȝ���B�	ʹ��� ��*�=�Eq=OE�Y������˄�W��E�;v�]>ݰ�j�-�oH��7֪VT����g��g�:t)}Yʳ|s�"To��Kw�X�q�rvjvy��z�:�.�8C����`z���q��	��'�#�  �N1B�H+�V(Q+��8)�wxώ��-
�U���ckm]+]���}*�ɞ�S�="�U5��n���������)y�㾈��u�����b���k�:_����F�nuDe!���
9��ʕe�{6g��P$�]v�)�ȴ���ɷG�1�Gxߋ������!�	�9�Vg|�ǏU��W�	��Gg��~�0�'I�\���<a!��cɍ����O�=c��3Ao>n$���kjwݙ�4u�y����z�uY�Gа,�g�&_�L���_^��5�#k�V;��D��G|J)�[C�6���'sR��ê׊��\����*m�ŖW{#s^�O��n��S3Rw�OQ]��# 3����Ru,�Őz�c����HÀ���VGbbK��&�|���m���s��������{{*�Ӹn7��i�o�nk�3�Ʒ)F[}Ωŭ��t �}�ͳ�ĳW��g������C, '<�m:�ۓR�m	V_T�cW�lt�R/��t�!�%��h�8P�·n���GyESU�b��k�V)>Y[���]J4p���ެ��2��N�WͶ�5W�}Y`P���~���
��km�l� +�Ѷ�֫Wf�Ҝ�S�b^{b�wJ��n2�vP����Q�xڭ�D�Pm�����,�"�e�m���Q��U�������i5՜�s�Ը�Cn�7��F"�ۮq�c(��ŭ�[�Iᝍ��[�Ե������GJ�L.���u�k��'��[w���x����v�t�؍t�n^g�96�"n�'�|χ�cǐqk2���l��G^~7�]^�9J=�&6�aܝ������@��~a�3�c�y6D�l�(�n��e^sC�z�7�[b�2r�\(ׁ���l�U�NZ���DtOH�Pΰhf�х1���Ȧ!j���C=�G6���i	�2�q��q���z{{�A�j/sgX���l�h�#��L��8ѻ�o��М<���,�]W;�����#��_����)��l�/L=��O��	� �l�u˂w��X�����3��2�2���:RPPhCpUO�NJ7:�ݪ��g�ؠ�5荌�r3�ŋ�J�<ph��F�@��G
��YP/�Q��i�v^:�.z;x���|���6���d���"D��|yU��9�~��]���+�>CT7Y5{����MڄhWj���&�?E����b��]h#y%�e�H(}~�����n�u:t1�|+}>���쮟"���S���Ū���y�������'`��g����{�f�V����8�f��!��l�ܛ�o5��7�F=�����T�͉ؽ�YRGj(�Zs�ޏw�b�j��SG"���l^IBģ.MX.ヂuy�u����}@L�ܜt�ԧډj�y�du�)ϵ���{�VИs*���z K>�ދ����Г&���|�i����
ǚ��pkN���+iJ<],�?�`5GcӺaގnv��0���F�hVXR5Bm*�[l������C�a�Q���U�!�J{%H�\��_}�9�3ϣ�����Q���^���<d�����Cn=�`�ʨQ,���� ;2���a�u���b��}����� 
���ջ�81��٥UX|d����v�'}3��!�<X,��R9�홹᱘*���m�;�����WY1*GQ���ڸ�/sD	��N��E-k(�����+���n���S��U�Uʎ����J�7�t�^�3j�ْ<�(��6�{ϻ���~���(��f���pȋ����&���`�2n�$��4��2z���Y���I��;K�tq��r_���>�R����S����5�2T��vLu��K��L!�n`�>^��>�w����{G\i4�t`��i����nv$�懓`�@T���j��WV}�^Y��%{v���⁆�E�H$2!���y.Gq�Ց2����!X	��j'��V����߽��bύ[�ǳw�u]@����*�~]^�b�NǱ���V�BS=p���cTk�2Z������S��r]�:������a�	����59�8GQ��Cv2�l`����m��s�6�aBI��1j�����C��}�"��ul��}�|��i�'^�,i�q�Y�;mR.F�=-�Hiעy[�U��1�8�uº�+�^��(� r�F0��yu*f\瑪sՄk��v��i�������1�U���3V�y�.�p8yLWK��p�}��,���q���y�`w�?z3A��Q	�	�TF�'Op/otw
�������s|&��U������� �ղ�(��rԷ1������
���i�)s���a�J �����j�u� ������X�lk�>κN�����=}K����v9��D�8:�W��(��32+v� ����{���b���Ρ�W��E0�	$�2�ڵ�oFs1���ȘX�y����;��6uMژ1�r֞1�&�""��({F�\�ٌ�(m�$�0�Paxv���В���q��xm�^	r{M��s���1|f�>T�}�zeB2E�jojz��}#�3	 ؄\.����Uw9h�<m`~����A�d_��ʊ����.=�&��&D�uC�E�xY魖�wB����`� �"铇��q̝���-S�P��=��#n�+у���;��Y�si���#y�n�M�X�\ڼ0��R�ܻ����z��5��4e�i����#Y���J�j��T�P�fL��{��¤�kYd�/OoR��r�9��Pt><��w"���{6�ּ
�2 l4j���7��^z���u��uV�A;��ɥ���jFgv���nE��a������ǟh���T�O7L9�Ժ����	1�j@�#u�S>��޹�nwa���i��u�MG����3a�9��_K���/��ھ�t|5@>ە��:1tNǢ���j��+�gd���FB0��[m*��JOz��78�q�b���u��*���p���2T7�L��]��c 7j�3�[��!�-���M��������+(O��eg�vўL�ν��ј�;ɪ�L��ש\�W��GG}�^��,��gD��%Ap��#c�:kdNb� �J ���;��9�:������hˀ!K�)�6D���qS��y±��j�Ov^� �4��Dpg�tTx{����	��7�Ҫ�ћ=�ؗ���$��Ό���9V�H����j���f�*�¿��p0Z[���!G'�Kp!�3D`�B=��b����,��![���w�M����G{7~%37�7�7�V� ��!�幖=�r�ٲ�����A�9M�&�= 32����.�C���~o�P����y��K+�m�q�7Ϝq��0���z�"�/[=�nN��/U�M���vc;t��n���]���|qVG�G7��kX�%t�6�o; i�j��j}�η1m�wcCӻr0fB��J�0@�#��s�H����ˍvҧ.�.ۮ�tхvb-Ī�4�W��*�s������t�&�\��;rg�uZ�v��~/ķ�_��GF��&��~��VE9��~�^B,��z��b�(��w&��U�r�|���#:'��V�#5���d�33^w� �gǷ�L��(��ނ��n���c��\�o���1����5��E���Q�
ho��7�6�A8�{����+��x��$k���O;�{A���K��C�r.Fs�<]�k�9�s�r���L�P�(��E ��;7|T��qГ��vb��I~�����;'�$�<wn����xq=
(6!0Ru٭*�܈j\(�]�a�1�;S����jU��݃�rͭ��Pb͹J�X)^�b�S�Z���[g��NdP����	)@piC̑���o{��P�
���r{;�Fs.���q6|��$�v��6�c ���T� �<ٯ��
@����4�� �a�7K��
Fߎ�Ln�K���[�]C2%�[rj}�>�w�_�/���Z+���9�n�c$ja����_��7�L��7U5 w�)�h���-����zd�*r4ߢw��t��`�u��M����R�}�3'�)�Ϣ3r�~�f�ݛ���;E:}&V�V�+oʬ�����	�> j�%�
��w�B�gk��[��}R�ҥ�=^�&l�X�h���b���HH���5w��������gg����5�����o�|�- �D�F&^���-۩�3�G�'�n-"�n l4��"��z����[fR�>��e<��W=�|Fb\{�T�>��"�9�r;Fj�3�01l�Q��Tt%p�r&��S{�2��Zk�N��j���Z3�-Y��<�2=�j�g.j8E<^�0�.S����Ѫ̀���s�|KҊ���P��c�ݐ}n�n=1���(��ʃ���{�Fe��9�̕l����	"8Ȟ6/�;���{�W3:e�ʮ�;37WPy��왪������� ?�*�Fdl!���ꉮ�`TQ��]��&3>������4e�A�y���)�4��F��b��W�&Q��ڧ���u�- ���K�/�?�����yE�Pg��h��;�ϋm�R����;j��D��Y<���ʥQW{���/|�Lo�Go�xPT�P�j3��h���~a��5 �qM��5�˖�C/(�@q�ϗWg],[X�O3�l`爅ݚ���`��ŀ�v�*[M|`�-�0�cѻ�����w���]g�b��X�G��ì���c_����O?Ek�ZNZ<U�W�U��Zq_e7���!AJY}�&v9gVr��O���ɐV��L�ň0^�*Wcu�|{�'�W�-����Ca��$�8Y0/���&�1r����JOWq�r�gzCu����}
�T�:z6���T�w_���A/"�H<�X���%�~!���~h��sJ�9�8��v��t#O}q�6F��y�iL��ЀrQ3�׭PKȃ�D^��4��S��<_���tI�Z!���U��|˄�P�p[���O���v�tD#�������'2���s�uY�����������x}$v�;+�k��{�68�sr'X�l�m2!���8&��͒=K5��Ȧ���}gz�^�X7��xgul�5���7�w%=B��B]=��/g'3	T�H�Ӿe�a��d$@�#-vR*�L�T.�k{�����o�~v�v}D4�p�#ү)d�nn�7k�;mut���Y76���7��YY�ظ�R�uY�xf�q!w�����v��ɫ0�U?S�Z��0�`��~��c��ͥ�#�#�o��v���1s�Ƚ��g�zƤ"
�3Oڶk��Or��B�G�¶�o�H������㓏���]�$��{{�3��<Ia��d�Xf�G��������X�lԽ����m�Y�db�Q+v�H�Vc���Q��ھ�/����7����)�N0n�Vq&�����6Gb4o���{۸Bw�QQ�5W\��v�_��)��Dt���cb�1�	<��v+��R�x��V�e����YaXfP���J9uѫ�je��u�.bgI~s��N�T���T�>:�PZy<�G
e�y�U�V����H��`A�N]׃��4�B���rQ�7�N,�l�;a�/�1�����ޟ9�m���bډi��������B����߉��=��H�=�"
��,�l�F+]Ӫ{���\yd�s��~~�5�Mոj�(L��͞m��]��v��%�2�iȁѫ]�[��l��&=�l���M>�W�;�o����r�)�W�/[��?X�6�T}7�w�1����C�IU�ER
F}�T����'[�~KI���EN�����v;e"�я�=+|��q�o��y6ne�e�5�7t�'د0����������㏌�[.4�T�mN��>V�,�8.��l���oPʹAz���t�3e�m=}t�DD�q7����
�u�I���uF����ѵChJ�lNT�w����E6<ٞF:��D�z���Q3~RJ���OW���(�sUF�γ��#w��1��b�����e�a�W�m�4j[���f�^��	�#��֙���Ɗ�� C�R��?���G�i9�ĺ����6��V���n�����כ��q���ǋ�'�3\[(�P�<lm�t���t���P/&8��qn�sKm��<����=�$�n۩gk������ힽq�'�|�<l�m��j�N��Xm�v9z�[��g�R�89�s� �����񎋮�Lx�n:�n������ۀ��[��:��{޳�e��'�����t����M�t�;�Y]�9r:_*��`b��]{�/��"���\d���\:��׋h����L�2J��j�vGV��XwIݞ�n#l�R��;kG����ݫا'N�G{��\�y�c'kΝ]��@���� �7�J(
X���F
yF�T_�:���M:"�qVݱ[P�u�D{cg��&ܽ�0��
�]E�U���E��������/�x�[>J�*����-��6վ��nRxV���'1h�Vc�Q;��/�$�A%����.��f�f��fT�j�h��7/�i��A�m���dU�ލ�(��8r���߂�豾�%�*\W����pہ
(u,ŝ86�m��˾`Nb���쫁�|zy��}}�E�A��Sg��f9B��'�����T3�*�nz>���Ш����L��f�ɢ�� �;���wG�l�ٺ�D�"������G{	���ݙ�Hk���2yZ���v��.��9g+��[w�)�㷫oO�x�p�hBi�قb"�[Y�Ly���k#mD���wM2�Z��u��2vrpW��< ���W#8�q�u��y��غ˕?�fvݛ��Fury���g;MEύ�F�Tr���oD;B諢:���8z�Ktk��Me,�pX�M�ώ���p�|�B�o̑�ҹ��2]�7��=��}�:�U�~��H�Փ)ж��8h��y�r����wc�c��ew������}Q�w�5A��;8���70�x��^�¸��7�Y|��bc��Yc�mw����T�뚮�>��ed7ԫ�gU�;�V\o7v�WYٔoB���a���`����뽙e�6�Bv�_k��48�}m*2�,�ga�J�=�X&�U�NgO�~L��Y�bc3;�VS�u���e<�uv��s���d��)mr/�8��@VJɕx%�&�J�>��z���˭U2��sM��s�9��Z[v��!����ݖ>f�!��oq*�������m�K���l|����]L�w�j4/"V�ol���H]E[���d����!���O]A��^�HMq��@�wW��*�͠I'�gss�$�;o�8�Egw��kO-sy�"&w���%V)x�W=�;'C�Wu�M0e���+��R4�:\���\��]t���SSYm�,̲F�,�����m<s�b�Z�oK��35F��^,�?�&ً.�#�;�q���b�O(�AC^2�Ր<�U�.�;C�#w�<:�oM�����L���]=չ�ndß�����ۢ���8�5,����uV��Έq��� C�m_-%��7�XB�/	�"�V1{�DI&6�i6�$����R�L�D�URr������6=�vz�X�;�:�&���)%i̤vD?kZ���D1
c�RB$�t�O*j
�%�¬nN��mc�v�S��qa��=���Ɲ�On���@�q�At�>����������t=�c{N��y�z������c9�e�B;q�ǘ�e����8�g�.+�����wi�N7[�R�q�r�K��N�Ϡ�8 ����A�b��N��/
�V�s��cݧ7]�{u�1��gP��n�1Z�i='�z��EU�DA�E�;�F`-����}��n�����;�pȜt�.o*���Ӯ�$cv���Q�2�t�f���ۍd�׀;�����=ƫ���`���`�v�h�]��h��*s�1WK8��w-փ�g�ά</��X؄"´�*!�U�Km�c8u�V��㨈7��6�N9�q��4g�2Xnw#������Rݖ�ۧrv����Nm˃����1K��۟F@q�u�NzA�op����W��Ttf��r�サ��㇂�*m�u��۸����[m<Ѳnl����5r��yc�,���o\v�:�Z�eE�'��#ۚ6�jT���n �����[7Tp�6� �:G�H�d�6��wj�y��t�^{��i�}M���xb�$q��̀�
�B[cvL%�����9.+�v�WG(�i.ׂaQC�u�p��Ӌ�1�v�ƷU�cam��q�'[�WGn��Muѵ�*��]�ۗ��������n`w)�n|�N�&.(t�f;uq���t��8��Y�1���㴺{bwF���[��93��53Ǵ������l�6ǎз7<�u��M���!��VJ�f۰1����w���u��kCݻmg�&v������ '')�̽Rs��q�m��qq��m��6y��r�`�8�wl�[�z�ѠTV��k�B�-Mnh�����>�3b�Nm�nt��-ț��^k9yM[���M��k�s��q�g�����m~��]�==�B-����j���?/*" ��֏=}7�ϛ��#���l�X�+ڎx#���$?�����n-�kGe�*gq��v�n��`¦S�n����A]l��{������#�&�H���T�!�ث�	u��B,ƕ��>�}Fr{��w�R�G�.2v#�]�H�yU�.ֽ�*�E���U�s86pȠi�A$A�&�r��Ln�<5�� �o�	w�wKq�XH'~Z���d�,��!v����j���\�&!����1S\gBN}�*B�
�ǉ�z�U�H��;�`LC�ax���du��p;*v�ќ/��/<�d��;��ʾk����e����qJ#�L�R<�l�W�j'S!�~��%Q��P��f�_mż��D��-de���N����T>i���a\ ��U�ӎ�lI�����ڳ�M �=츹�lv.k(�����xVA�3��*�c�r�]�58�q*��8���f(���>,�"f�"/���/u�ғæ2^�ƣc¶�v�����������%h2a�m�b{o㶷ch��0���nƤ�8B�[NT��yog�����T�]'@���8Oa���n:�����f��S�����|sk!��5ԱC�w���cS)7�}zsw2)Wy�+��ˎ-���u$���u��s���Xmm��:�gw������^�"�G�̢U�.��N�{q3G�>x�I-���J�F�>��a�dӻ���1�z�b|�S]�j�힪���ln��f�p��m���]g8����� �"�u N)�3�j�|d�h>������3֯mD�ӕ<��L������GQ�����$��0��q�~�H�g���]�eA��^'`
l�ڊbpu5W���HF�b��u��'c1�-���7+/m��H��v�b���k޼�(ɅRa�j�e���K���%G�
,�(���\�&ٵd�3g���jS��	�S.{���co�p�4�+�d�"�u{���j��jEu8���o=z�L+���!�"�PS��u!ك�^u��X!�[< ѻ�^���]�TQTi�|�<CS=tn�t�ms��e��a�n�ݻ�c��'Ju�7��۔,b9L�=wu��[=����������>�cD�59��,�\n��ʙ{��%�pZ%���,��t��#:ѳ6��@��w���v�>.���8������c�T��Ze�\_J��}~��0Ō���jn�1�IBp�Ͳ�:��&�����g\��9��uJ4֭��u��b����iҰ:vVk��I�/��m��RgC�wY��>d�A;ʑ��r���z�y��[��+#3-z<I�Lɖ�U��aZ<w+�U1Ӟ.!w+�Z&AO�y]��
l�=.����ut<~�v�����Vj�w./z7��&�0�b+��`�>���ʽ��t(���{'���&o�n�F*�J�^pd[ۺ2F�ֆ��@�*M��K�<���US��ܜ@/�Yga�݂ �W�m!���N�J��)��0lG;�SÉtr�v�����F-�ì�.+I����m*�v$���p��y�W� �P���w5<jK[�c.k0����C���s=��U��
���c�C��{�V��˹�^η��:�����r%%��)���ocai9*�5гEo���� ���|s-8���y��d���y�,TT�;����v��ǉA��4B�C< Xʼ��������m���T��2c���[���>��:|�tN*gL�~���WM>�~z�2��9л���! ���L�'���ުځ/�����^]D��5�'f�ײ�隊�ZP���[���/�)g&�e�Lj�+�`Q��}�I����ue�-�~�=]Tmt{��A��H�%��ĺ�qVs�8�Z @�jA}1�L��5{�� W,�b㺡|�ћ��U�Y}����z`�O3z�m�'� )c�;S�13����t�ۚ����Bi��ꥳv1����:C��{zͦ 	N�ͮ q3��E���c �vv�pl�+��v�{r���m�^.�c�H�\@#��7n��g��2H�q��j6�*�#�����1��^�\��t�k6p�s/%8��G\�.�7��Cl']c�t�Ϝ��v�0b�L�;<��'� Dc���ONZK9�O<���c�����<ql�6�4�3�y��,o m�h̄��0a��t��Ch�6s��s�N����^&G�M��r�Q�TϨM����{S���xr�����=p�)"T���[3=�Ɓ��a��[|��ᑣ5��uk�	a����RWT	B5���E�m�� ;-ɍPt�Vy��M�Y���v��h����OI��v#_2�wbUx�j�f ߻gGluN?���!��}~|�Q�m���nX"�i�ny^q�[�tE%(*(�G�v�{9���n�+�h��� ⬨�X���>�����2�N����uDI^��0#�,��A�:,a�Ca������x|]�I%�3ン�e�����u�R�\i�̆��t�t�2�)o��X�^�f�˜��	g0غ��"������/ ��V��UR�MS݁��V�~'(���m��J�7��X�^����aH�{���H;��k���[."<:5\l�W��֑�'�|��e��<���q�7O*���fWFմ,z������X���f�14c�U�s�R�)惺c=Q��"�V{�^�gw!�z�j��w(� Ji"�&�r37��r���1>9�Q<�s�#�����=�E������5�.:4E�{WX�p/��H{gb���I�+1����ע�ТaW�u.�w:�z��1eژ-��|:V�o63��h�hs��q %f/teht�%g1�kT�b��.e��؞M��lzoʌ�K�*q�&�gk�c�Ȗ`��teIܙcF���譪&�1�^����qI�R�<�p�D1�ɳ����sxq���>y��Իy�x�$s;���nF����o��+DOzd>��j�ԉ�4�7c-
}��6aS>ɺ���h�.�&�*\G���x��=�E��E^DI=�3<6"�`Jox]��Vy��T\dI� �M^����u|�9Nk�ҍ����Ɛ;�;���vg�:�0P 4�P3����8��VntNg>ȇfV��e��ӵ3}�qpR�2E�m�#��0��3.�We#,�!މ1��J��=ZG)����ͩ�rs���!h'�[�L8b'��P"wȼ9�1�v,����3r&\d�{Cӣ����m=V��ߣ��ET���"��Uޏe�j|^�SS׵����
�CL��q�=���W9���}��nu�3�η<Hi�ۭu|/f^am�����O��<�Z��������+y9Il>0q��9�yR�}�F�����,#P't,�^�"�솵k�]Ԇ\�w��`:j&�yL�vB{x�za�tm������Q��ۡ���z�[��3e���5�wT���˭>�B������\ꢍ�*K]q����=�?�(��Y�񼋃�NT�X�`�F�`��5o\��ڰ�n��Z�}]�`��C�gVX=��ͻ؎�x�.��ރ9��h&�0�3yP޾�[Ks���x�u�r�=ٻ=>��)�pǗ��F{��(߯�&'c��=koҡf���"�OXz�����7�6�����A��0�@��5�њ�i\�E��ĥ�PY����Nz�p�c:W�U�����5|��y�Q�	�'tB I��l:�In�D*G�k*"a���p�Za6<$��"�VfVPq�q���4Wj�=wݚ�����;�8�s(\y��L;���	[ƧT�����\�Z����t�m��&� �D�Fm(	�䘾����~��~.��flW9�픲��ϮoGkގ���|/�i�����:]�b��Y�(p�	�
x�)��/:9-b���+0�J1��brD;Ô�y�A��M��/�Wl ^ɺ~�ýך�/�p�9�M���� �P8g�;��t���^���m���Ƈ��泫N�FHH����w�u�D�ut3�Ϲ/+�����>�j�+�D��O�_9�;f�\1���߫0O�?���&��E8M�K$���5�{;S5T�Kڻ�W��x�����!��Q�}�0L��m��떨��r��=��h�"epG}��v^�,��-p��pT}a4��v[���kU-�P�|2�[1d?����;z(����&+sEa6��ol��J5��#�M�V%;��}\%n��Ω�x
eU���т��{���~�����"V�n1;��Ӫ�!����l�^�#�oc4��C�زq��Q��ZUR�OM���C�G�9��2p�Ia�i�.�g޸��^�vT�P���ێ��s"V�����j��������
�V�WN^Ӄqڶ,=�&;;{Ofk��X�"p`�`��D�_?Eh��?{�*�:�J��h�Om�yd�S�:���[T�(n'��y��i^[u��-�e�+V�^+�[6��ι�3{�����?&�~>�ᛊ��ޅ��ۙe�C˵�Unny�6���=r"��\0[V��N�*en�H���Ve�s��]g��ԩ=�َ6ǿ?�?Vf�e�TR��6{�G��5�ő�GDN*C��/B��lX]W�{מ��C�m�_&���Fz�ȵk��N[S�:9b#���s7��7ڠZ��Ii���%����1�>3�H�a.�����6��w3�5�7�g�2��{���L�S	/�T��<(�yY��Ҧ�wM��qmڞ���q�I6�|�<z�V��k-�����7ۗ�z�s/WAV���^��{�g�mVwt���%$��ϡz8��ߜWמUD=����s�g���ޔTx�<�+�p��X;��&N[]-2]�O
�4v�釡�o7k�N
�c-7J��kb�{����Qܱ��e5ӆq��1R;o&�^P�h��a�l5���Wn.�gWk��uƷ1Y��<v�����t��D�V��n0]n�+ك�v\�+7O]h��c�N�v����m�j9u�)݉]�=�t���N��9�`M�/j��h.�ٍ�zb�W�;֖xiN�����g��2q���uL�	v�A�#�6�ss�:i���qa���8���6]խ�+�n��]�X��ny#�o��O��Ɲ]h9����#U�S=�NH�B~�x�	��ν�y*pS��/.������w�/��s��e�!�U��<;.yzu�T��P��tԸւ��2u�$"��\:�N���";����p��k�����=|9��m�S>n\����:��FΕ�J2"g�A�.�Ys]R�]��B�_ 
I��i(%�E7��7m�Hn��\��-��-6p	,��fO^o����*�J��z��0ס%�����g�̙�
L�\Ll�p<���:�mqS{%X�ի_Ĕ[&��=�F�e�;;���!e�� \M�J�J!V�F��:s��������ͅD�@]�T�0N��]�[��u�����]��*�[�>A��x��6���ɪ��4i]5�C�ݨ�= �ϕQ�~�˦�o%`Xk�we��^���ttl[:��������S���\��n��#~)��T`�̚f͛�{����G�E+��8 ˌ����4cf���2s_J��Wun���W�V�����+n���!����|�L�Mvm������;�5W��C�ݼ�U7C2��K1��2#޷\q�K�t�K�$w>�R�G��c��j_�։����ӽX%qL�\��zki��7��^j��zy:�-�+%d��*4�<�o�E�/�˃�a�͛5�]�^�79Г��o�2��뵖��N�<Y��M�a�71Eq�=�g�|{Qӵ�G+]_��׉ %���{��q��6Hr>K�o>k�s�p=^�v���A6���n���wy^4O��ީ��� ��~y�,�ᷙ�>} ��B:�kF{c�r��]l����2C"8e�q2o��E��Bct�����fMDj`,$U\J�DDn�b
۝|Uj��*��1�������	�ͭ���:�{4.��r��j�0�]g��f=�J� ��Mf����1F	҇��;�����g��pX�Ӕ��[�ř5s�J�U>���S7�U�r�$U�ӭsm���^)��y�u=ɕuO�^/<x��*�n���I�P�X�z���C�涳ޯ^�1��;q�d��xl��2�k��^�H0�0�GNn��#�v=��Bm7�E�R.�u���ۜ���Do�*(�R2s���X�fy	�Mٽ��Ě�b%ҿ[�T+����x��j�[����fb��ޏ(����,(�O�o)�g.�gw���sO�,ڃ��R�`���6V�Qj����������艫�a��<���BZGB����3�O��M���5�vjU�T�7����8O5^NyW8�{b�/��~���c�^���Ɏ�����d��u*�/5�Htu�����Y�o���%X�]m`�w��j�i� �R���37�p_Om��d�K���� $M�����2O�û��d�ܓœ/ϳm@��8�&+�n�jBo�!s�v�;%؍��5+�.�gz��=�eʭ4��R������*�ŘT�f2�^��?W�=�YY��̬߳���]C5�3.��5��-���JR��zk(I7�t_�zԡ0x^#�ǻe���t��燉k��D�<͈�z����f�p��Jt���ߥr�wI<ͦ=�����O50{}�Y5S����EuϷ��D�9:�L���T��oC1�Z�	e�BM�]�0.zN�&���k����Ѫ�ݒ-�N�\+z�������h�MITs ��������l�S���W����h���AHW��oK�L8��!i��3�و�;�$8M�A>%y"ǟ�{]�����旾N7A�Y]�FC���:�\%���+���;��}����O��ޥ6�:��S��Ȫ<a�6\�m��$�*�|��γ�<b�7���ɝ���d#�/�M�2��qE_T���4Ţ �DZ.��c=[��1p{��WPh��sc=u���bKظ��o��S�۝{2��4grmCd��/*K5vbp��qp��}V?{=����>y��1�C�:�cw����[
w��S� �̭��Xz��[��^�d��k.�Y�i��DOn��+�*�	g6,��ȘΒ��xZ�Ps�宝�ۓy_�*�[�SYAc������罴e=����R&ډK��/[��[��sz
)кmg;��ǉ[Z�6<�}�֢�:{ٴƩ��:��=(ܷ*�DIe���Q��w�u5mԻX�.�р��;1J��1�.��Cgb�쪘5��h��Z�n�"�Ň�8��(�$��X2�?M�J�����\G
ȹP�4;��ͳX2*͙��u��.�칹���y9�z��S7�`^��k�4n���η��y�ᝆcG��W��Ȩ���f��h�d#s��u�}B�"�[��cR3k��Yͬ�L�����X^����Wch*�qY��e���yhG��_fn-e+�gwT�κ;�W[%�˹��V�Qn�3�M��@)9�Y�A�����uv�q��4��7.�6�j���z�<����w<��`+6o�n�i�2��x�W���;�Zkp|�ӧ}û��y0��Y�L�7��`�ꔶ�H�X��X0U�؂Ɇ�y�+hە��wF (��,�ۣ�i���-�g��/w����(�;+h����}'gomP�i��ރ��&2��͋�k(���=:�ssGV���N]ݣF�<�l��!7���|K�7��m�l�	�J�Y��,�X.�u[��种� #�I��gƛ�N�&� 8�b�G�D�����nocN�[jjad����{*Wd�)�V �F�*g�����aV��!t
��V�����ɒlkh�"�wzx��B�ʹC�K��"��y}�}�̇&&�zf��&y��H�w�S��灺S��sZ{�#=W�o�m��-�\�2��|����ء~���0��S�f#��)}�{��H�� `<5�ճ/\E��g�
4=&v��k׹d�D�a�
&_jH���������� _�M�h
�^���퍙ɛ�|r(�v=������/Չz�;��p��=9N��u�@]s�7���YxŴ�C��D"őי��GtZ��&mW��,s٫���[�9��+~ɇ�*%�j �!!��?و�աtU>�ܛ�WgJ��|�d �<ΞT.J��;�f�Y�=,���ł��-��`Ǩ8�����a�2�JVר��H{��ݝ�Y��٠\g���ުn罜:�!�m ������7iwtꚞ��ўj�����XZ�p3��"�pM;��]1�Ѩw��(7aU����{��ĳ��B�zL�!�+b��7�.E�K-��U��4�6_mv�d���&��iw���*�h�q�����S&�#�]l�cl�������αP�iaJ�܇��7�&V��C��Ym\�3���;.Mz08XRD��$���2\In<�v���W<�N�m��2m��w=���
�9��]��<�^�g��~|Z�9���{.��C2t���FK�K�k�]��ǰs۲����7;�ogP��ϋ�V]����b���|��ۛv3���px��;9�F^H.�\k/���ͻl�s��#�S���;cLsݻg ;�X;;�'^����U���_M�����#�n���2�K�YmV���u�4oo<�� a�Z����R�#�TlU�ʅ�����ʞ�V�Ez�����X�,�jɍ�Y*O?#[SX�y�c�3�3�iLq����%��a��~޹BE�g%�B�p���K��)q<�L���/���c:�}���S^{���n1�RU%�DPvnr��؁]���\���n�y6	i�-��|��<��'[��Q�����RÎ�co�+Qٝw$EځaΏ-��<���1O}�g�[��f�n-%	 6��eْhguw�{k�ԞU�������/��������Ưz�,7:f*����zj�W]
	U8�}���k5p�O��M���
Y��=ܑ�zzV���Ҍ_�I�+�;n��j�v��n��<d@�^'�Y.��&�vA��2:���/������)f��#W|�e0	�Ww�a�W��y5(��
dny��6s��<��W��^.*7a_�͆(�њ�װ1�h��ʉ���W��]��j�t�D��Y��$��BL�#�#	
��c�L�3���,�ٛqcuU�i�-C)�Fau!�,���k���f"��6*i�ӓC��O�2�Փ5c���w���VՇ�(9J�Mf��e�B���6:T�n"��:;���D�:!"Mjr�l�����PϹu�?1Qk�7C����?tq��`�%"lę�L:�i���'?�^D�/��Էɴn�G�v�5��@g��w̖u���=s$��a���J�z;~	���G:0GMs��r�vx��Lq��<{J��1=��tL=	��x�����jVx�<�8-[Mg�,󼬕D���L�hlt��c�DdG<�l��y�]&4T^8dO�#�j�&Փ]���gvn6[��w"�@	y��pwd��4 ��ͷ��3܁��L�˓53��q0�T_��������ʁ�q���]�e�H�Dn��ǻ���í��М�B p#p|�&֐i�c��䙅Z��u�ҬS㻼��z4nr^��2E��=�����z��C3i=��Rb���7��E�L��6o��.�XD��0�tmOe�4��:�Gj��3T)Q�-ޚ���ޠ=ۤ\x�5vyD�j輟�>Y5������_ZW�n���!�	t���]��d����ώB��.��\��b���tm[Zu� ى�0����un��p�%��I`!��m[ 6��͞��h�h�7Y�(�'��V�Ġ.�?2����RV������V��t�ZJ��4��NF����@�F�WE9��e���Z�����Gt��T�4ImV� W��z{^oe�ғެWh�pS!�����6!M]�H��W�A�	�LЊ��Ĉ�Q�����d�+Ѽ#|�̡?5�7'��q{x�{7#�E*��������&K�~-��t�8��r��5��e���U0�Ҝ\��#�z�~�aV�ѩ�yt�������HA�.�����	�������+o�$��)��'ˢ��]��ֹ؝�1�;y�DK�9��]���U��ﻕ��fƓ��a��Ki!������"�r+�[��Na﯇/̔����JU��s��ж�6�&���3��m��h��5W{���^����G��r���R���s;̻�}k0Y!d�H���=�b#bk�U��0RM�&�-�Dug���:��%�eđ�#�ޱ��m��� NHF���J�*����ؖ�Nx���bv{a�1�,y�?1��e�o?ut��?���N�E�U�G زm��ξx��:��v#�+�6fg�뤽9�w�ͷ�^`�}Du�C7�NVV�Ӣ�-7]En��V&�>���cMW/q�w
#.������pp�2���F���;����O0���m%�\O��ijwoMn�u�зֶqm�S��p'�i�}�Y��Ѣ�
����n�C��V�֢�0X��V���;�"\�Y�IG7O]`�v�����4��<|E .��?~'<h<o:}���k�_���Y�]LAz�X���Y������ߔL���;�o��D�/z9�������g�,7jfI�t���{�iv��i)f���Y��ߧ/m7��9�c�c.��Q�������b�i�Ot#��|t2$Cd����dq���E�5U�[}3�ױ���3�U�z��z��+&�U%.���=�F�v��w���0D��i޵�S=[.;�	'�����fj�Njs'n��E����3P�LgP��'e����%����OOY��i�dm�B�����S�d8�5H����7yT���ӂ/��tӆ2��Ѻ�R��!��]F���Ļ�AFhم�;���ܪ�@�G�, Qm5��cM�I�����F�O9���[��r�'6�������T�S���;�8}��Yy��ds���(�	���B���8�'~��o�&�6Ջ<s�3�����畃tyC�����zA�˻D��Ep��L�����F�r|J+��=���:�G��� ��`��Y�.dg-~�;ٛ-Mgq�x��%�T��&3a�������k!�^��;��N��3WxOB�-��ʆ�w�M�		�wRVf�K^0��U�Su֗r��%��y���r�4���L�z1qLG�2�R	J�a.%v��K6O\74T��>v�ϙ��'�=�*�v��ri���y�v8��7��ZF�p�n�uc�.��r u�r��N�:Yw��f��H9���NC�s5��#T�p>�f��6JYΥz9x-aG*�d�1Z�����6�Ӽ �t�W.u��]p^��^��@�Cۙ�����z��K3�W7\:��H��8��smO^8��-�?���
{߿��_��b�\���>޻�b���<L�,E���k�v�@ �l�l�m����q����[u�ȂI�N�����$n8��C�甁��㶱�7��g�ocf%�Ú-��&��&͢�yX�&�������� /�1�tjBD�[���#��[tzdu����r5��&�5	�A80�g����H�eaŤ�N)����7/f�=��s�w^�����_�R���~�F�M?=y�lE�CD#%߯�
97I�|�7W�Ҡ);;~�';	=��i+*��|瞝zp�젍lס��~����"6םv���5�#�Ν�\�q;��9U��z�"�$�3�E���|�"a�9�2�F_�'�*$�N:�V�4�)�4���j�OTM��&4���_T�7�ф6���L��3�t0���(G���I�鯻V�Cz�7��?o=�'�I�`ѝ�"=8�F7bj�_$o�����+�<�΅f�캭�;�3�U�=1^=�9~�nM�r��#r���
��Bʺ�ӹ��=gӑm�;���B��@#܌"a00])��.�E�Ex�����|p𚮑�_oz"9�7�1���M�H��B9���/=��G%�8wd��J�Jn���Ƿ;[�e^��4��4E��ÓR��v�Y�4El���e^t�}F��3IO����z��e��q�.w�yڷnV�<�Sg�w�N���N�]%W-��� ��j-0K6�}bN�:G���F�웅���C�W�H����Ls�S����0ɄRj&ါ��l�Q1���M|H4���"�(��>OuM���fd.ŭ�"w҇�1��~إǅ�ˋ:�0�Ms3Wk`����'�Y:V�z4��ɖ���-���m�,��Pcf��+�u�4��l�U��2�_Ep�6%��]#����/.�z�1�n��\��B��Q�s�sj�:|Z�q�n�K��̳㇇��P. 3tM��gB����g�{#��=��F��\v�i������i9*^�_S�*'L�Ja!�v_T�+*�s�mΪ2�A�	���;q�
��8&Tp�=��0��$�lĉo}�h���cI��t��������c{y�W>V����^�a}��\n~;��T��ٟE�A�qw�b}z|{P��P�R$-�]�S�;9^��-\^�+T�����@����d֘8�<���}U��Toy�J[�5��s
�7^�=���'�'��zlL��9����>�-�`6�O43������7��P�۹o9H ��F4'�������= ���0�˃��sAU�X�(�������Sd�����"sgm�>S���o?'+d/A�ɡ�	�Eم����f�y3'�R��bDJ,lu��y`��ZPb򭊂��:���ov�<RhvubE����}�s���]
#��)n�LTkX��Ê�8�V�7/c���]\�n{OYM��h]A��Yї1/�8@Zu�D#�ˎ�g)ו����敎:O��P8�Ug�I�!�XI�W���pPWP����S��;;��~\bD�Y��3'�����Z��/G��Y6ƻW��~����SYBb�*����8��ԗ���.P�h��3i>t�]+�,L8��<:�@Bzg/O#����Y�� y4
��T��U���=
"f�Ӿw%���1�4� g�gvb�6F���C.�S�JO��D}�G1'Qط�>�\͓��u��T\��`X��w�|�W"�a������O=�^�����0���p ��~~�a��G�q��=~��ا�b��Z~��:#U��ܡִ�Vq�����qRw't7��>I�@_#hQ��p�G�k������h\S� ~?(^~������y:+���\��z��{lԲ��|i�`{u�P��������~��c�.=ҏ��(�i�����n��
�����M/{ַ1�>��*	�9�+M-�"+g{�r���#��˂a���������(㬙o�%��� ��eB����/����ܱXQ:Ԟ�>���v`j�:G"Q����D]tͮ�����$M+i�vY�Y8�q�� M�hE�Bv9򪬽ڃ��:R|-�_�����.ʃ� ���-ճ������������A;�W11g,��UB���z�
�qS�q�7Hɫf�B�{i[�k/8�뷖��k_ƹW�Lz9(PO�X�D���g��|M�%-��X��z<�Bp��p�[@�)�Q��*��Ê�����njx���z���l���eo��I��<6�^@��x��D��k�0#	�]�]�{��h�*���kG�ץW���g|���+2o�]�����Y
�k�M_��g��'&U�����;���~��cj=�cz-U����Fn{�/+[H��U��15Ӝ�B��p�p�:�zhs���n�����=�~��ֲ$YHR�FgӢ�>c/f�p���v;ps�2b��]�㐷�{������6;��Aet�7�_A7b�lh���O��Uڧjh���
�F�81�7��{st�¼٭��.g~��A$I &�X�9S�N�t���-��YY���حWFb�qV�1�5����;�wC��G�:�}jə�!�G����_+��@5/�F��t�u5~ٍ�ʀ���KH>�8������ݵ}���(.&{ޔV��N�'��ѩ�Өi М�Y�^�sn��炘9^	1{]e���;���
�ٽ�F$�=5u>��;�p�i��k��;�1zW��u�/|��|m@&$v�Z�W������m�螳:�
7�xrj�D�Ϫ���ۄ&%����枝7D�4�)s&����;��\�ɕԫp�N��351��LS�n޽�Ƣ2�F��
�ph�2v�K��
 �;��6��<=��dLn�^�j�c-�뭉��ܢ�9 _����V*J��,�v�q ��CÝm��n�<ܣ��&(=������7Z�����aۅ0uE�.3���Ϫ��x�6��bg)'���l�:�/�kgv��x1���(�%�;C�V;$�ަz����';m�\���9Piɔ����=�}ߟߏƺ���M�l���0sw{5�N��D��Ui�ͳ9Y�H����>��P4�H��u֖�39�j��`���àcP;�Ղ#�(�zsue���%��`x�zݮ��=BdbK���{��1!uHw��,���ț8:��9I����U[vxW|y6<C3�1Ċd>�s�㻗O��6����;mv<HH�(|�X�6�Omd��7��g�6x�GP�P-�E������{��؜�f�\�8XC�<��]��D�N-��s��j#Dv#����~]�1�sQ.;;6�wi/qiS0�_^�M�3��2.�b�p��L|�'�;R�>���9�#��	}�82UJ���U��*������s��!�aB���rb�	|�>g��=n�{à'��i������1�d+��@{�73� gw}���\���V=Y�u��A���tQ	~MSMP����g��1���6ݙ�uen�xo?�OK��0���qBhO��sP[�h�J8��4�Y��*�~���w:�V\�+>|>a�"�BEEl�ƣ���M�fW�/oTW+���'���RN��u�̨`��7��W/�1G�c������v��
xC�^eãY��Pz!��L�a1|s���k�{��"l�b�o�u�_�!c�f-�<��"ģ��;vb��V'��m�y��O�d���J�3�O�$�+��?���s:�����mu,>���h��V��\�x5:�ip�۱��瓆�˫(P�Z��������1z�*�n��z%�В���T�h��^���+u|_^fjon��-J��޺�2f�du��Җ�jq�;���^��=i�.�]�+1�1���ū�]���Q��4��5-s2�r�7�#���-7�t�F^m��t����m�u��l�5�)6Wa��}ċ��]c�-�o]�n���|gj�%C�V�;���g5�[:N�r�;4.�[��V�^��n��S<Q[[��H�)���sY�#�Vॽ�Iae����`殦v��*�X���;�-r�+ �aѠ���պ��ed���ù�o͋�5�h�o�ї��6��}Իl[��M@U�>�e]]��W�����wL�PMh�d�z&	��j��W�5X�%3;:���u�DI-˗�&]�s%� ��2���ϲ̶p�RT��Fv*�7��dT~Ցۮ�y�����\V�:V�:��;/Qä�u(����w\�[��vu`5�l�X��p���=�k4��S�6�u�!Z���wq^ԧx�ը��r�9�L����U��V�yo+e�ޫ޻�F�\��o%.�.��m�uw�#P�4�QN�On>��E��e`%-�8;�p��VPm�쨣/w�6�uK�֩�R^2�bV7mз��m+|(�b�Y��Ě��wnK5��uǓ��hv's�Vľ��[�Zɼ�JP��,�#\��+6�tT�$5.櫀�Bb�j�Ш�j��ګk�����{��Q�z�����N2\�3<�7�w2�Nu[Wfd�ې�B��qɮn9|���˵lWb��>1����쎮ˬ�����b2<m\�I5��p;����O�v���wW2�-�X`j7B�V��PT�����ew���=9�k�{:%��|�E@��N�obxޞ�"��d�vI ����v�q�3��k��9�cō����vQ8��3���xIx�n�k�ʍ�q�]�9�Cj��$PC�%ȄՀ�$Pei�ܐ>4��չ��N�60�栍�.����u�&�:��c�${��H;�87n��"p��ڣ6�9�-ASًzsv0�`0=��]���=�OA��3Ч.����ɑ����E�<�V��lv+wL�3D�ݹ�X�Lv���]��B�O�^�c��1�$�˶;W$k������T��qm�Wk�˫T:������H�F�c�::ȕE�.6��R���1�a�4�{zS]k�u�K��=x�5���V��^�J��o0rϷn�q�=�	ڑ�ĸ�;L\��{(\�8��Tx�t�c]�`����w�w��q:8�����[v��mV��0��z棊ɵˮ���GN��Nۋ&���dɻ<��ln��Rr$V˸��w`��^��F�汶��.�5�����J����ks9�<�.�Z�Y�� ��5��������v�f��6����ݝ�Ü�,n�ȇ=�1��L�PN�cB�B6Л�vG�&v��fV㝱]��{6ܶ���d��k��*:P̶�P
��TBE#px3����GF:,��gq��W5����、/8�.�+s�7�m<I��0��޷/O�j6�d�)��#��Y8�KOv��6u�SrNNv��Ee۰7l���n̜A����������wH�=��te��3��(��e����=�Ns�їh81��'g�ni��:�á�s������v.�m�s��`�;`��nȁ�q��k��v���]as���j��:f��~�.6�gˎ�&.���~m}�^�Q>��R0�m a����B�b��x��S��{\��F��AHWç�OOlvϓ7�j4��ERVI��۫�ma�ra�XϨ����玒k�#ֶ�cگ/￟M����~��k���D1&{�F}�E��߾�IN~��yJ$�َ5��SB�~�glţ�����0��X�V�$D��nu������w̢C��s�L��^��i|/�ftI3�o��KM��?6��P�F�&���W}}Q������օ��b�1A-ƻ:������z�k�g�j�.�5����w����P�� J����Vk�c��_��s�mtќ�.���6�#�a\�>z�E�1���o{�(o|=�Oo�w�uhŤ���4D}X`�Sf(!
�=:.͒�`�o޻��A*/Ѡמ�u{���Z詋��H/�̾�4f3�ҟ���e���ϤOw����婢�.���PQc>!��?H�ys���PSI�����&-��O���!��^)��{[4f'y����/�ٸ��,�����}�Ο�gߗ��ǻ�u&~<bG��J�|%�;�?oX�b�vD�����12 ��U�+��]�͵�\���?1�p�(hΞ-x���{K������?(�2�j�uPW��0�V*���/�<��G
�~���"�ܪ�ò���1���c{`��*���
!�?lV�����\3�E���$�__{���_8/���s~��'�#D`��b}��٘��\��B�E����F8@�LAffdŏ���b;�.�MS�P��&k��Q|SF~12����L���4�S(��ٞ*���w��im2�e��m��+`�:I�q;qv-u�<@��S<�{;Z��z�f�񢘧���֚��1$�_�<�xٝ:%���f�|*"ow�H�#�~�>`��_}r�#�Zؿyo����PK��C�$7�3�O<I�T^i��0��y�ycLC�Cno^��9�Fb��]"w8Y%įI��i�]W��V����ד�[�\e�U�׌����+g}eWH����~������G?���SX��3:(io�U����
7٪��I���8}3��ф"8]�H����^{��͵��Ι��.�JS	Mk�.���x��@����t�}#��Ӫ��b}��wy6��Z����o��jţ����e�]/�w�Wm_{����j�"����hL���e2��mf�l���f|w=�bf��}����DD�Y����b�{o;���}�׏��/9^oB�d��Vb���J˯sY�q��C0!�b���:��ι��Q�5��B��oz��ҙ���ST^���<���ټ����-���n�6L�G���6*$�mb���3���d�!��'����D���2b����*a��<�?���?��B���_<�%�1+��~һy�1~1�1�?	1b����������`���#�������x���7{1Y�hK|�y��JG���7�f�P�	o����^ֿ3�|�^綰3d�W}��I�V}���i~�5E�&.�}�����w��ipW�~�ܺ1t�ś�Ku����y���ϻ���&.s�D��k|]�o��=z�zb��2W����pT���hL�g���&~��h��[>񘫟{�_sp��@%��Vc��T��55���s����RP_���F��[�t�ǔ�L �`��p�.�F�X�[t^�.�8����ڀ3G������_���w*�_�O�-ǉ��+�t�IEǞ�*��]�:0XC�@�� L\��9;?myf��҈�1��2�H�D��Փϟ�,���z$DpO޿mN4����
[Wy�L�3�(-�������>�[��g�o�<`At�3����(%����}�ߞ^�KD���~�h8��!��]Q�=�O�&%�E�_��r~���0�@A�Q"8|�G�7'*bM��:1��Q|c�X�8r~�~Ǘs'��� ��I:��Z1�ǽb_6�_H����Nm-vB���esĽ��.��/����9wZ�W*}���V&0�N_t�S����̲��\7dM�"feؽ��ݍN&8�͹���b�y��3�iQ.�k����[�y�_�NW:b����Z��C�����E6�1��	3W� �g1/{��7s�c�]gQP3�dxG�x`�f����qCuU�r����"�0QB��	S�٘1�fw�w�fh�|1~�gL}z�?EZ�&]��׷�o����b��\����a�-	7��\Kc�_�;��p�(}�҉u�%�5�E�q�&�:�&~�>�.͈�1��#�����4P���S@��	����n%	�	
q)�H������߭��t���L�E����c��Z���Js���Q�3���FgY�{�f(,�rc�!U����DU��Y�'ƽ�����LZ�׋�1v�U�οNg�#����}����I����Z^nF��Gx�G���d��]��@K��%�8�!��MpJ�	�i��*qJ!��EM"_e�Ǣ~�P�Ȓ�m�CY��p���3�7mDϜ;��oW8�i���8X�V���?�{�{���2�C</�1|3�b���߿wJ�fgϑc�������o;�f>�(G��G:�h�(!�9y6	˺���*�t{�H�n��U��L���!���+{�y��e3�Z\-i3�&(c�5��}Mo�=[�g���Pζ���k��������Uc�~�$D!#��gy���S����ō����ŭɉ^g�؏;���o=!�!�P��D������E���w{�OZ��m_k{�~�[>���G����b(k6vvX��G�ª��������sj�<���K��>����_,6�A} 1`��n�������Ь���pG�Cy�����b�!�rn���G�:����N<�}2�!�����}5���AxX���d�u]t�ѐA�8q�B�d�L�%��n��K�8��5 �S����I٬��|����b7{��b�[NVn���ִs�v6K���{�vr.i���m�\##H��;��e""	\BLQ��b�����G�F^����컧���#�E�u�.���n�����\[$����9�t�:��m�'jy�k�]����'>�ŭ^�k�կ]����j�t�����N��m[r�xG3n�����j��x{	��n�����Z�ݥq�m�$wX�<��k�o"�k�A�v��k[��V+T�-����h���]ߺ�/d5��{�d����Ͼ��CD ����ٓP�?@�R�1�~�Aa�>�u}ޞL6���&���#B��Q^k�쓰�OH�L*(
���Q�A��F����ae�M��"0r�r"2Oǵ2bם߹��T�kg��j5�}w�׫x\C�W�Le�*�>#A4zL��҇ф��M�^����\��C�B�Z�=ҴQX��>�*�+�{{c��}�$x0��L��=��>jd�?+�=����u=9prF'��1n�7z��������Z��n�|%҉>���ޅ�g�wyZ���g��~8p�At׹�i�B׶L�̡����g���ABe�"�r?G"&p��od�A݅��.�ꚓ��k=:x��`$qr!.9��W�uWJ�Yw����O��I֯hc�%3�F�k#�'��U�":�B�3U����/g��	C�;/^pP��X�3\�6���%%�0G��յ(d���(��"�E8w@0B�����c�fՊS���o�D�"0�N��$��V����4%5U�X�_LWgezL Gf(���\~ �j�{t�}�u�;�mQ��V��L�]�����x�{ѯ~DU8�ey��l���2�>��Ǜ����Q!�"���:�{)��H��1иC��n�>�w��"�o��.�V��7P�Y�?H��F�3<��4cj$7�{KPr�o�:!KQ��s^j6'c��i0�I�r�����Nt�����Z���m%U�`�f��k�Y�ķ�}��LT�����&k����[8�xb�ёP �P�S��T�~�~"�ŭ������I���]�r����wu,�:�V��i��^�wB4v����n���0e\Ge�R�t]����D��v}���&;�=~w*��"e�H�cov6��9�1!��E��O���%�r�v5� ��ȑ�����O��xޮ�q1��,4,1[7m{zy��&�@�g��Vuv:�-�^9���;e�nユ�up"Yǔ���#���(!�o����q���p�2>�����FG����mE��}�*��2~}r;����q1L��ڎ+���ޜ�<糪�̀=�󄑆�*��F��DyL��J}Y�/�\=h!������zU�><CK�Ԣ��b8DZ5�7o`�x���N�!�-iik���3��n���ۢء����C?W�L[�wT6)�o��f���?D�(�U"������8T'��SV湝�8~<�b�w#Y� ��F��}"4}�]�n��}��CY���[>^QS��ۆ(Ej_h�p|DaacEz����!c謞1�%S����Ƒ���Ƀ�=�/���&�7���rT���:�2������ַvϲ��T��$�j�$�=]V�n�Q�_�7bk:���+P�Ȉ�!o���߈�l�g��3ܼ�����bh�B,��cR�ݷj�Dw�  �2ٌ���	��3���ވ�~A!��_]X�c9;�G�E�Ty>������a���
2-�Z�T���;�㗞����}�����wb��Lk�U��pv�f$v
^!���^�O2�J(pDd��O�)�W��M�@��g��>�*:�e�l?a�����ɵ�u�j�m�`�{�G�v��	^{/g�hBA�Dx�ߠ��{�r�Ϣ{�*P�ta�rC?s���Z'ϴ�c������94��|��83{�����/��P��Gc昵Ⱥ5>-�ʝ�#nq�+�N�	Bn�p���&ih�ˮ�R�ݦ�tNo�ySgs*�v���Yc}��!AlAjn��:U���j}^������z͆!��#G\v�ɨp!��} �Ԥ?ڱZ�jo:f���#5& ى��Ks�?
�~M1g*I���DN���Q,�nq��ܛ�& I���J{�I�)�#�،��~d�%D�w��Z޵���&�g��!'y��t�!��6 �����#\�);�n6���B�Q[�?p�j8�as��R���ޯg�_�l���r^('�����n�6؝�b#�n]�f(}쐴.�ꔈR����u",���,��p(Da?]D��x�㡏�@���|)���)
�
��:�3��N���}E�H� ם̍�/�\�变��J����о<z�\`�".���<���E���ɘ�G�O�s�<�;ܷ�(9*�cF�v��;���Ƹ�w1}0�b��M�2$z�Q��ZPc�V�����3�E�\#qTOt@��L^��K��0��DĮ�\��Ξ�"hbNP�pQd�t�>�M�z,>�Ԛ?���ݻX�z�8'!����N���'��~��/�'�r�w��zp|��x���Ӗ:��ԉ�� �1����`����?*�xm k�YY����}lm�=��E�\�f�Ymp��
?m��lD����C�Z���X�MoW3"��)}�j����a����ɻs���"I�gD0��8�ܙ��<	~D�'{c��^ ��6�t0i$V)G�Ц���'��M#*x>�s+P�wq�X�69ϕ����}Q�̄2�q3B��N&@�z���؝Ϊ�Nm����i�^��,
������O�^��ac.��~�1��^��+i� Gd��r� L���tL�o�ē
yt����ˇ��tR�^�����d�VK�Q����O��9��	8@,�n�P%�3��{�oB�NE2�ΉF;/|��ޮ����ћ�!B_
0υ���qI>q�'A�_.>A�J��2�'�| ��{�f"��}QN�~�E�a�n%s�M.)��=�=P�)�f�d�ET=И�%N�� 7�snꡯ�b8A��$�����2��D��^�fUz���,�T��t�鉓6��]�g�LP�G��;SW��L�2��E���M� ��b_��Uo������A�v��[&�f����n�rۗ���nTv�e-Ӫ9z�e���ڻ�-�-�� "tA;�>��LK���E˛���>`��Y"�V�NG+62���^@F
.&
6��=�{�^��3�Ǚ���l(���H<�D���eL�|T�D�=`��;�$�I�p6l{��\vkH�-�?r��k�x�vW%� <��b|�$Q��g)�b��z6�;~��̂"¿�V���X�Ww[繑)�o<���*������,}�%O��ڧ{�
6���0G�F1Gv��������=�z�
����M�O�M�d���q�k�L�i��J�z`U.�p\0�L�Sb��w:�?B�

s��8w�����,�{}�ӝ��V���ʊQ�X�b��%ĭn~��kz"f���\�}1����ij�3b����K*��FM�:�2��Vw�S�k�W���դy����]L�70�<�� o\c����5������t�
t[�c����Gf�6���N5�����Ė�Y��h)���>�#�Z;���,�8\�ͼ۳�ƹ�y��m�v��{'Q���r�{7�{p�<nr����h5�½��'T��Y��d�5��R��C>̻���}����a�k˻V�nx0�<8�8�I�+�P���񲖪^��D�y�s|̝�P=P�5�P�:�=]��0pQi��tX�B��ǐf���\$Y�-���({��i\ȧ��ג>#z�tD�r3�d�u��Tn���g�9x �yhޑ#s�r�Up�{�Y9bD��8�$>}7���H��d7$]�_^BP&`�����ou`���W����r�~ڏ_1Ul0�Hl����r��ݍ�u�OZ��.h��K����c�})v��9>���@%��GK\�#񼂰ʏ# _Oj���f��$_�t�F�r��|^�}Y��צ�����?�@E�,�pn��?Zq��&t&U�L%�Jt_L�ѤO*�L���&�j�{��hF���<W[c�&T�N'�B����eb����`Q
��Y�{��)wC'�!ŗ�����z��jjj�ft���t��'�y�^�E�<��oq��G�'ET��4ן��g�����(a����U�QU�anopA+��㉝��x�������(0-���1޵ZЁ�B	��*k�{��M��Kw�/bs1ɍ�C��� x�DI,<��ye�s��Oϝ^�;����j0f������_\k��蚊�������l��J_�_��z
�^S�4>��*%I;R$���C�3��K�%��d��\�SS���Ldxθ|��[p��32�)�ĝ�NĜ^�ٌ̽K�̽���r�v�����L���`�Z�4�d���&����*+�� g+�t�x8�Q�/�C�짶�*$P�=�����5�Yn�<�|���{w{|��k��0Mi������'3�ޑ�:�dus�r��L��`n۩N�r^1�q��=�R7e� �Ї���G������|E�2�s�����U�D���).ޜ�R;��{/�8��׾��ˬ�[]�^��ޤ���4�2�<��3�my���]LY��*e��Tl��F���d�{��`�t���Ӝ�w}�&�t��:#�����zI�G���&:�U������̒�l��<�<7uH`���v�fX�t1�}���;�I��W�ٶޘ��QXNV,�>��k"{Dس(����r�Y����>��r��>Y:Wb�S��֪)��n�<�my$�,M<Fv��T���a�3~��PuzUi����Ҏ۲�;hfόߋ����n�����Q������dq�K��^�5��z6<y��M�*>��1^[=�O������z��Sۏ>�ީS0BSI��:�tfL����̨h�� ���Cc�el��/��o�u��E]�\D�
�g;lGmڜ{㺻��D��s�}���&vl�I�\Y�<�u$4�l&.&�0��Ti�u��Dnv�"�[�Q�sk{J���R�	���P������]��,�yH4��Rų��3G���N�?!�zU��H�c�	��.v*�7�^�ڃ����ya7@t��\�k�9�7B�3�(�*���1�v��9����b�V���Y.��d�P���:Bg����}o{��V��4�C�2�)4n���}E<�4e�dT�64�ݱ3�MHs\pV��qK����z,�h����+1�Y>ڛ���0����_��N�aD��%	&���Ʈ�-��7snr�U�M�˜-��u����<,V��;[�|�笻D���aǨ5��<6�F�b4����lÞ7���8A%�,σ��qYY�6��+	�YX�%��JFd���B��c=*F���N���s�qj9�!��a��:<�\�B���`x�-0~`s���1��{�Nqy7�Ѽ�D���4±dv�@tšz�i�-��� �͏I�;`�S��T���^ð�y�y�J���Ea���C,{�S}����h��q�E�{j��|���WL0t؃�=8u<��1��g��v��nE�e�	4�hd��������d�K��Z���\�
tn]��&��>6[w+K����w�0�f�'� a6��r.�y�4뻥��!"T��x��/i=9Ma2G��ؚ���{x�t=�D����V��r��h��S�A
_@�Ȓ�ً�U�ً1fg����Y�3?�ff,ř��K31f,�iff,ř��fb�Y��ر,�ş�fbř����fb�Y��1ff,ř��ř��f�,�Ř�3��ff,ř��fb�Y��,�Ř�1����fmb��Y�3?�,�Ř�3�%���f�Y��1fg�%���f��3b���ř��fsfb�Y����e5�q�Yp*�� �r 	 r}���y�H�YJ*HT�
�&�dV� ��)M)*� �*�Z��h4�F!U��&RRL�iY�h�QP 
T#�  d �D�R���	
V�RZ�P@��D�QTQJ!$)*�UR�
�R��AEH���R�M%"�LkMe*V������i�k��;e:�j����Ylf���e�j�6���Һ0�A7ZU �ow�������kgz�Z��=� {������Ν��o]��x���w�ۧ[�'���֡�����3ۜz:燯:��k�ޮ7���wv:�p1���NۻO#�-fV�)F2*��Q+�zw��Zu��7��Z�wj��mz�=gb��;{+ݻw\p<g��î���^�j��9�o{{6�f�9z��{��^[�b��͸w����n���L�R(�*	(�o{���Iw�[��)�s/O�wnGx����w�{�=Ǻt��y��J�[�r���꫷v��W�m������m+�������o{���w��Q 
�JD��ӯm��s��6��t�����w��Qַ{ыwg��t͹���RK�y��rʷt,ݳ����ȶ�zsތ̷���5�L�J)`i%P�J$��ѝ�Y{Ǹo:�j޼����Qs����mZ޵�����ݺ��k����k�z�=���ҵ����wkIV�]9��rJ7�8��V{u��T��G�*T��y��.��xk�Fv�6;�z�KC۴;�׻��׌����v�<��]��N[�=��ۻ���;g��ק��^a'h������W�͚�B�"�!EQ]�]v��{���5%�ul����޺z����^w��ܬ�t��Sݲ��{u^��n��]�3]ۣ���� �4)�-D�J��J���vjx,�O]�{޶�z��o.�=z:��u��4�l^#�����h5e3L�����;���ᨊ��JB��%Q�s5e�r�Wn�w�;�I\4�����8w%WX�]S�mu��[Z�v�mm� �{ e)U M  �{FR���b2d41�L��C ��0j��	JU 	����� �T`   I������=OP=OQ�S�����?������g��fM�3���=��������=�o���H�M��� !	$Ԑ��C� !	$��$I%��$�	$��H�LB!$��	 BI?�/�?����]���p^��y�;�[�w��zr��o`����ԫ�F�|"������"�cB`���-G(T{�%�e��	�����2T!Ojޠ��ɍ*-��Hw&0����u�=��2���;�Y��	�l��(ռ9�]����o1��j�#�$N����h��&��Rҵ�a0��*"�whdYP%��4�q���F<��`f:�j��][���G��˸M Q��F)L8��d��ۭ�AƮG��:��R��sK�d.�WW��x-�4�n�J���6��J� -Ɔ�3�Q��ya���o.������N���ò�v�/ugMѵ�-�#lۭ���YGM[��%�*3\���`�v���leS��P��-�nXx�!�4U��EE�!�$�r�8r�G0�ZveV�XVژ��*B�ƎU�V�~���{;O_O�f��;�)�i�}���R���>�a�-��g��W�d�Zv�v`�Y�
�g�V��xF�8�a�͔�����7G��d|�Hc!X�*Ad��R$4�x��Cl�0:��C�y�H4� KT�1�Q�̴.^�Ck�v10X(�7oL��gl�v"5:�Oh�j#���v���0ГvYM]���k�)���#vY�a�(�f	eqEr���=ǵr�� �:�L�!ZmԠ�˰ⶢ���8ULS\�P�W�ބ^L�U��YU����Xs�u���H-�f�Xc�ѻ�R3RN�4V��Z.�`�̢)�0ѫ�����nʆef�
ͷ*[��i �{��\X�IW�EF7vlv^���=QVT��Y{���	���A��53y��z�"�)ۻB�Pt~a�a�n���l�Q(/��!��)��
�\��3TWv�Ј�m
��艭R�����%�/".o�
��82^͔^�`�ь���PK�&�G=�ɶ�L�;�C�Y�HfQ��d_BdM�KT��f�����&�a��S@�#w!t�,=�w����,��ظ�f�6�K-�d7I�+te4��Gܕ� Eq�1�yZ��{TA7��&T��jAlFA[�#8�BI�dܕ�T*3YZ����t�[�H����82�^%5 �qP�7Y�ɷ���!-!ZM������'��1�Y��q�U:��`�Q`6��qe$E�h�q�ۑLI�f�����G�Vҷ�����t��v#v��Vz�;�Q�6���B�Aui�aW�А�D���onl��5m��v�4H�u�v�v��x��k��fäQЌW��()��x�L�yBi��l�%!lj��nSG2���6w1٨��[.��F��Ɗ5�껻5�N��m�ôF��Ў�Z�4���sOl`Uc]e�)]Y�Mv�7S&i�����ϭ����J#Y��I��1軐:͆�kQ�	ݭ���8
2�%%�w��Ɉ��D���t7[����AEGm��5��[�F���DA�D ���tbB�r�YZ���)�0`��:b��)v�ɚF�Y����}%�U(�{z�:R�ܗT�Et��g~v��J�i�컈���YM�d�O̓$1$oI��6�(Xif�EZI��X�����fgR��4�!a�m��dd���Yq��N��/�gRñ�CϚ�����C��X�'%��&��#����n$kJ*�XV��Ͱb�4��vvCF��$�-�A�w�nU�K�֧T����KE̊�e�5-)��-�yfɺR�����a�g�gH�,�)=��������Q�;�W���
˚R�B��I�{���޸������HP�������w4�zY��.�!t�tj���6��x�M�Ե��xDeGe��:�N��˩V ��4��R�]�O62����B�k��ux�P��&7&�Vқ1�c�7V�ZEƾ":k1�ڊ@��TU;o�(躛K6�k�BM�����wQ��>3b/���4�d�`������H���wY��;z���1�T��Sf:�����������ʘ�[*��(��_6�b��vU���dʠS�7e�M,͡��]7�z��( m$�����-�N�*�N����Q��U��Y�/p�J*����hq�W��b�ڌώ+�NB�h|��LƄC0�B���9B74\�k5����n��>�4��$"a��yM����t���(-�EdY�����t�]`TZн[PY�(�eK�PzĔP��{V1a\h�I�Z?s*J�*7�,=>ݡ�!�d
�K���"�@�ww�.��y��5���R���G�nB̪�;��[��uB&�m}n����41�cT%��� �V�8N%y��y
�ư�ta4��,�2���q�(����Ҏn[�Њ�H�fa$c��D���uB��	8�����~pm�d`�s%�]Y�cW$:k뫲>�Y;�3�5�M�3r�\w)�`�ŊTC �(�� ��b(�mkKr��nA ԐӰ[B�ݬ?\ի�K,�4�.䪱>cRܼ͹h�BnF(�3j:[`�˕w);"�D@�2�N�a��(c���*�8S.m�A:1a"V���Z	�����a�z Y�$:"'�9��{���y1�eԣ�ɵGj�����	�qS�{�R�Ls-
����j�SR�W�/j����p�d�f�b��A�1�&���H���oMv1У�5莃S7^��ڌ��7,#*�VZ	�V����chV̂m#H�	6��.Tϋ��a9�z020J��5ǡ����ݶr��Շi�ˉ;n�J���ذ��h��<jDhm�H=�f����$�U���̈́�ӱt.:�&P/j\^���#�����-T��2�N�-�m�)���t �o�4�A�% Nё���������9���f��)k,�e�-^#F ��0b�����]%�t�Ċ�1�d�ӈ[x��&՜?^��4/avwf�м�����z�
 ����RC˻��_�+
 ��0����C7%�)` K-�&U���9�T�!�k �l���b��+m@�-�l\��,�Q�*�`ne��5m��{O�1�+1Jqi
�j��Zq��F�`�n/@h�3^(e0p^T�]��t�i
�Q���u�ї2�`��%%Լ��0A ��Ȣ��DX�/(�ۮ�]��d����$Je��ͻ�i���%�ڶA�x��
�?�� �)M!�	;Y {��T4!yO3�F�[;U�w�q�M�V�c!�#���&u�E�[g/I�h�P���KC�FE���
�x	e��t2��$3�M	���W,Z�0�hf�F��xi���[�ۘk	d9�����;h;Q�%�)Up�	df7��!j�B4cWMRi���M��
"�X�.�,�)2�|
B�BK�n�P�^�Ȍ�����f\d�À�h�ót���i���e�lY�ZEc ���T����4ےS+l.ͤa�B��Z��]�V�a�����r�m�r(%b�UP�>
��A�.�cE¤M�����zm=�)wM�KmTta��CWY�N�>��i&݄I�L,��.�z4ަo-4��$�AOv�L�:ʳ{�a����V�����VPk�戶���Hb(^�7%�72ӧ>�f �o]7*�")�%�t��ޤZ��ܤEkt�[�_#���!>_V)��fZb$ˬ�N`#	�ړ�ݙZ�-�r��T����!�s�X
)r�Y1w`���R�x�ދ�VO��OlR���c�ZUnc�� ����mR���E��V�l\�սkPn�skI��v��9��dP�RS��:s,���a�`�h<4 U�V�e㽸�
���Ջ�CZB�h�[�|���V�/.Li�Z�u�ZKvZe�1��2c3nc-]��`n(mm
7��ϰEyb�F
�r2����S����E%շ�j�Y�A5PE6ӏݘYɔd�sr��i:3!�*M�&Ң�V������]غ�d35:�DK�b����W�KY���XWo~n��W)��Qa��woߛە�
+XZ��y������9���ׅX��4�ef!���G�ӌ�P���*��:b7�cR��oM̼82"��-4�J�8�@m"�!��<���S���_hҭ�墊:�-Q��2�����IYv�h����t��(�w�v���2Uֶ=�w�y�Rݖ�s	$YH@��K,��|�����i��[���,.�i��!�ޛ�-���@�o.�is"% A*�V��lmDCl�:-dy�3F��U��TH&����VJ!1��;dbT!�r��0YyXh�p�
���5[jֶFm�K_ē������ �n�%YWl�bk7����ꕇ�huֳ*j2(���&���-)��\�!��k���썂���VY�d�aD �j�r�	�,�4���ᦫZ�8�+幔!"��J�� ��ͽ0^�A

?1x��yYp��ѫ�[zH�{X���N��6�G0" ��LU�^��V��Xs>"`�^(��L5l���u�(�P$�)*�
\�Uw��n�S��+��U���	�0��ֶG⪪�u�Iڏ4m�H$F�mŅ�E��*��y�F�@�b���̶6���u ��%��tI�`˴�e�9p8s�G�5*G���j�3�6:����˾f��0ċ<et�f\֤�ɳ�Gf��z5����L�����r����1��ݙc�X�˳T\�,�+kq��X�*aђ�V]�ǋUre/�$#�Ru�q�%˫J���n�߈o������5Q��+Z_#�.�#E�b�/n֙�P���P�,^��+X�iԼ��L�F�JĴ�C���f�չt�[������ޠ��ُ �� ܄�Wk��1du�+Ff8�Tn��������� ��5������#�(�4��.�.��b7�Zku݆�A��+I��V�Q�UѰ��Ú�M�7M��R��S4r�,B�\�*��]�p:�@"�\�.�$ШA1Z��Wk�[[�Xc��X� S�%^<ʑb�Q�mY� $5��&�{�yp��Y����J�GK�h��V8�EZT&�%��QE<�b"*��m*(�j
,Y֢�n�E�j(�AgZ�)����h(�A����1�A|��9��86Zţ�~�*��E�D����y���:�U&vV����kE��j2����bQ�y������./�T%F1�
:��&� �;J�ר��`�����켕V��q@M+@�{�f��S����	��䲝=�UU{�Cz�7�s��R��3~]�_��ĺ�Q��)�3=��:sPh���1��Ac`��Ut����C��ؘ�A��*|.�Ჶ�M��:1|j�s*>U�WeR�5��ҕ�[Y$��(�K
'lɲ�\ٵ�����,��/�_21�gO9{˵E�<�)7��r��v�V��٪�͚�3h�\l��"��*�w�TW��(� � �	N2��3K��71��p�ֵ{����w3����2x0�����A��T4������-[��)iL�p������۽���%��K�ݿ��^�-\��|�M[�P�l�VG7Y��"6��k7�4�(����lJ�&��X�k/��pXP�KE^��3bwMՔ�%�P҆`H��Xy佼�{���+��"bQ� &YD:�0be���DDpt�\y���O� ]�!�+E�;r�����M�R�¦}����/e�oN�F�7�<ɬ`sv;��?^�^:�Û/)%-9Z�r!J�f�B�������f]�V�,�j��N!LG��Z֏Ȅ��jʟ3l5u��� ����dj^��h:U�	�0�L�0?�����������Z	ϵa��[7����t��?3g죶�
�D�
KԂP��4��f,r�-4���DT|��()���׮��/j躎kj��,3Y���07.�"�N0�Xܷ��U�G��dK"]�P��cF��S[h�����p#	�HY��$�(�ب�WT���|�$u�[7Y�q�tͻ�&e��N��xh��wV�����k5u��<d�*��bҝ�Z$QJ	3Ml6��lX�vN�fN��gO<v��XaYf���%�����I[i^S�ӎ��N^����(Қ�Q,sc��u]A��7�
1�0��Bm��#��|lX
dD4��)zwO���*$^M�8t�Iũn��54�@�j�E�͊��,�Yd��Q�Y&�wJ����p�ʧ�hR��4oMfKwl�*��P;�b�Z@N�e�?Y]@��ˀ�ѧk,�4D?"s6}XI������f����m�_ؖ��u�(ⷆ�.�F��qP����B%��oQ��f�U��oE�S�hĴ�RT.
vl��La��be������ܩ�2a
�e���0�_F�]1+2X��72�Z;�wQbԅ�P�0�+i˶�U"t���O>/�x�!h2XB�ʼګ����W�V�θ�F�`ǡ*)B^��l$v&��hC��W�G2T�
���?"
Œ͒o3M�Q�7^h,�!'^-<����/h?Q}�_��ySay�y�.#�˻n`�/0c�����݄�$�	�!Ǚ�gD���-q3��C��L�#"�L-.3��0��FE��I�K,�-�l�d��{�%�M�=����\�TI8�\�%��}"I%#}S���݇Y;Z嗠��<R�9;��Ƕ�(���1���Y'#�ޘ�or�޴:�v�d��޵ט��x��K=il0$�D����6�1.nBzI����(j��6Ѥ{j_;��x�k�$�����K�s�.���lL����T)X��&���o�R���<̕zbF���\�E�]��fV�HȦVqۂNp��Y&s&r�{�$�y1�����OI���GwYh��w���#m�vxn�Vf�sn�gi� R  �%Z��ٺ��"b�$�)9fg@���yyws�`����9�c�wĢw:�&wI�#}$o�V��G�1O�'�=��in=l��[�2���'<̴�Y�qR��)��z�;�ԉ�N-�}7x�"IE�:7:\4��o���&6�����J�we���ݾ:���t���eJ�U�sN'O�5}�μ}���ܗ�¥&����j��rva�bJ6щs�>r��9Yw����D^�+I����nkҏVEk
��Z1 ؉bۛ��S%���5/�U�\t�^�*��2�4�a�eX��v�����b�����vǽ��o4�=���NcWue�7��+����н�a�n��5����C�%�0��[����.KU1�ۊ���'h�JW��[������f<g\�j��%u��9.�l�^V��u�c��W����X]�wB�h��9��OȈ���K`wZ��(�p�t�y���j���ytaR�f��;0���p�;��k����N����w�e�9�a��Ѻ2!#rm�r�=��u\s��|,�lV�k9�����VZ�f��*f���2�	B^u���y-M�y�(������;��=\y[��`�\��BY����>U����xJ�[�[X^2A#[��ȮHiT'<�{oGj�U�	P�/.I��X�#�:��h�P�ɒj%�`6�����1f5�m��&q���U�:��l�T�O(�	�RY}��v�o���'��� ��U����30A.]� ��>��(���wJWvr\��-��N�h�,7yϰ=�I�ût�W"v����%w.�v]�2{�of,���9�w	�3vAdD����:E�#[����N: 6���ظ�6�=xz�ws��A���|N��Z��hs�mA7&�r7��8:�`)QW�W7L�ը����(Q�ɓ���-%�(Nd�8��H���ǠT;�Τ���s�V�������zWZrI�$�,��-7x���V�q��fn��3���k6w�=�wD��} �>��+;K��Qub�Z(�;�䜣��~K�q>���k.�b;)ׄm �p�����]n��ָ��Mgw1���X��D��%=�wwy.���ܩ���V��́�əۮ��G��j��p�S�.s[=�I��ۧq��;�#�����I�p����R0������v �4���w�a<F�6��vuK�wڹ!��oy�2� Xm�r��}�O�xM�Y��,��ֱk�m�j���a�Li��Q��<K���2E��ݷ����o�G��S%�ޫF2a�����$٫!�I�ѭATr��s��شd�%`���'<K�f��v�&�";���~f��U�*S�Mμ�u��.3���m�3$��Q���]v�p�]���6��E��U�K�R�������]�i[x�"KQo���l�H����SY՛���{K�ӯ(��4:`S���f>�	m!�e��y��++�c�ԴZ���y�U��uVL4*0U�o�����Pթ=D5.mU�ԑvp�(�l�
�l�(9/6������\�S�◜�-�r���q2z�n��;ś�	�V�-���9lv[Z�*�Ml뷹��(�i3��*�wm�O7*�/��q5�;&�4_hHe��6I�j�(���V¸�Ц�}JJ�4@�y���S�����-2	������K��'��;o3l��i����d%L�v�����Svc��mM���loKm�Π��JY���Ӄ��������A�f�H1�r�⫔�*�$�ќ�'.��3m�X��ێ����
��|	�N���f�ڰ�\�9A��C���=���kx,wM�xU�&j�;�FX�腝:���z�W�;/���`�4���̦a�l��=\gN� ���'+�\�d���m����H������BF­�NqIT��U�Xo���(�2F96]��!Mյj�e*�;.�UN�.�n��m�g,�f:�:�]�$z�{�s����`���3o�z�"�K[O���+�L��q��Ve=E����]׍��9����p�/��%"�=���e���< Oy��(īg��4�4�/5f�{�3mÝK ��,��B#��j�ŝ�\�v�839&���B�e]��ڷIM�ɏ8u��dݍ��L
R��8�7Q}���(@�I�;��ݙ2�{|v�����H�b�[P���GYWG�e�k������]�T�GfI� \�޽]�ЉRHKȉ�"��gs�����$�'��m�C��:��9�i��1o�n�u�e�a|4�F�G� 9DvwgD��Qw+�1��h ���7]22�&�u���`�DF���<�>��w��y�E�_*�L�.U����v�<z�A�x�%D��2���Ŵ6圐[r�Hǎ���b�͒u��nY"����Dt+�fvMRV�+���T�7�߸A2��7�+͖�9x*���S�����]�ɠ�,��%��g*�Uq�eB� &j��D��&�s�{���t)o�����{�ȡB���Ȱ��x�m�[Z�պ�S	T"�u����J�x��q0���m;d(��G+�=) �d��p�;�� .E.�Anr�"����-�����9ˡ���g-�b=��l]mE���&�����Jed�*G���ɳe��HVd�fM��õc��w%;|.�͜�����o,I�\C��L;�iq�����5�T�:й#��;�㋸v�3p��Q}�O�ҩ�g�����c�鶎֚"�o�:T5��|)�W��\=�����@�L��#��a�t�d�����hL7]��}�K�Nؙ��ԗ�n�E5����Z� �qc�u����v��V6�5��OgZ���=B:��+�75���6�\���%;ޱA���K�ִL֭�;���˭κP��:��3{�%c��C�35:��B��C`)���p�ܽ��K�0E9ԏ-�V$Ӽ�Z�&whM������]�>5ԥ�E����uD�%�fA�{�����)WIދA��$mo<�yhIu1HJT�,��aSL��w��j���c��A��Xө�2뭗x�8�@�
t��h�);�y�Ѳ�r��R:���;v6!��t�s.b�]Owv1qy�qF^uN���U��������.t-u�VMo:�wG�'&�z�Wr7�uff�\q�i�^����N�=�
�F��Gf^�f�S�k0�I�I�xΘ��'$X;7]9/ya5Ǥ���t�I�*QEut��#�,j�q��ꙙO���ܒ4�k���nu=*�)���9N�紷{�y7��[{,W@�WǍ`��(�,�ϊ�X�q_r�̽K-���<�(kv�R�{b�R7��;vd���۲����$x�·�h�ww[�1�g���>�ȶ
�k��w8��K�	sߋvIWn���o}�r��f�@_b��=eLq��v�8ѕĩ�^FnӼ��w|�pC�Ə-t���\^�n���M#�O~�C3p�N��=�%�y1�FXc/��;��3��Ժ���ڛg��PK��AU�h�|�ɖ1i���bc��d�����K�����h��oz�7�fc�ѱhKx���
tFL�sW,wuXッ*�2�贷b�m���J��wfj��q�w8��n>�JR)F��J��&tPуT[�1{������a*�\���HG8O���6I���`2&6Q���X�m��fj֭oS�(�	7�n�L�㩒UWr�A�7KSXj�Cr��W5�NK̙��3��[�C���t�:(��^�@려gr�ݱ265S$�1��僘ŅL潨Ս�{}���0g�T��M$�T��wx)����h�x�7k�+,���I�[՟G���r�Żu1<�b�>:U	�F;A�4���M���y�36�R��>����q�8�� ���cm�(�;5�\�T;Ϸ&���q�#�I�����B�=Y�O��U*���ѽ����ۣ�92gj��:�Π5�v�杷H�F^托��N�U�%҂xz�Lbn�|����9�wJ	���x�ƺ�M��\�e�F$���uQa9��ns��Ӷo|g�S���m��.+�^�^�'I��3;���̈́u���%[�nwfi���I�2Ӑ�B�х��զ�n;�(��5��|S�q��5F*_dK�6`2ɩ����qq��Q�a��Z���)��K\t�"���'�P��rz�Q]��Ŷf�C��Ïq��2t�� ғyZp�/�X2�,���G��
��v��s�X9a܎�ߚgv�1ńXډ<w�3,��AK��c��^�yG�{�4��cV��AM�t��s��ܣw���
=h��5�P�d'���Ӑ���u�4醼�^e�N�Z�o��Y��^��|�?t��#|��'{P��ǹ\wl�>k��~��x�` ���'��_5m�da�ɻH�?(���,����/��|�x>��YF��x5��+^Ŭ!���ݕ�;9��$�
���#�\V�N�ם+�"I��h�ɻ}�n-5��J� �dc�
��n��|�v�08���� �F��	�M�u3j���kX�Ν}&�����\j�eqs�.o+��)E�j�3��ם��}ݵwa���X̷�`��Fm<�O�B�]��e�ڳ:u^Ǣ�t��̲����
M����i��d�;x(�&��6��ٜ�@�*J���T+�q� C�����\��O#�/�:�D�嚮��/�k���'$J�bc�}|�#Ϻ�N�3�wT��N���9�E�tYZgvo7Q�Y��,�R��v-v��\�d���k����{ӝ��.�,����Ak���h��K�{���Y]w�e�t�����;V" h�VZ���v�,ur��=[.S��MwF�4U��h;/mi��6e����W8��N�h(�yw�2ت��S��9V�t2���m�/`�(�f>�:�g_%R?��.�͟&ø��c�br+6m��eI��>�2;���S=B^^�g)T��X�Z�7g�����`�u�Z:�.@�e�u�0\�ys��86��ֽ�i.A�im!r�JI�]:m�r멫l���X6�2Inf�8�l]��LpɆ�-Rf]o��ޡ[��*�u�l:[�{GE�d�f�6�Ҿ	��ۭ�r�e�iWʭ�\���&a���أ1˥};Mb�y�G���c9�sZ�4��r���Q_3��rj?fs�S�䬛:�Y�b:G�f�7�qBy��۱H_�Eۿ���__f����S����lL���0��Nf�w��n^ ;:]��|.�,���+Q�m�V�
37�ʎ�v�<�t�X���n�Lܚ=f7z�.6-eH.@���VKj�z=[B��U�/��A�uY�c�q�<��Y�U֞�6p�H��ʦޫk.�[4&�/��T励T������냗]�ĺS|�nm�����ň��(ʱ�d�*����=��u{�N3�����S�s̴ƈ'��>F-sY>y��m��n9�����D�3{.�	�UM���c.�c�}i����_b��l�sg��:2�m��a�U�,��/��LPZ�V��ϔ��/�<#���7��vQP�U�t�7	��<��&k$�:�Z�ޮ(��
�%n+�j�)�K�d�Z&�f�uϖc�>��C}��n҄���󵽝ч����w ��	罣�r)�8i̽�17�H��@���f�Ӿ"����@z�D�0"�j�3���[�5P̧�#nAA�u_j4i+ChW3\(���r�U�۪  }5���(��q+�wP���/PGmQ�`��:��2����u;r�ҳh��,w����h����tq��FP�W��w>���Cm��/����G����{ul6D��kj�����i�����"�UVY�yǗ�����ΰ��`1aKmL�*��4I������F_�V T��сz�,��O�Cmv�':j�Ԯ�`�֔`����E��e7�*��N�f�����z�L;M�Z6�&�
ˎμo��W��#�<��.��V9���|�;vf5'0��	�Ղ���Õj����g"��7�M�wԍrwa#&[in��b����6��
�͑�`lXu��ț?;B��\Wӭ2��]V�^zjv�o)���7��#am�8�v�wb�_���v�ZmFn�<�/��y9��WO�����S��I��V�q����5ۀ�ti�n��4������i
����N�o4*f&�S9�oorv.���U��8�`�mb��X���k�s��k��Xܷ>��<*2%��q��G{ChcU,r9u����u�����c��>��$8���D�������Ɇ�gח;&i!j�n`W�i�"��t���:��^�]�o_h'���S)���/4t��j���$Di�1oGZ\,;/p6�v��-����b���v٦�>䋭���A��{k�uKM�xߑ�ܺ��I{�'��,캻B��yɮ�;�
�x���҅�k����y�n����in�MU��S�;ol��oPą���}z{%�5��++x��D���8��U|��Ը�K��,2n�me]T�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I5�kZֵ�kZֵ�kZֵ���H�O�!$���HO�@��k��,�}����z~-M��m�؇ƞC�&�ow:��Ô�C��j�6�����ٹ�ّQ��X�엻M�*x���Yb��D-|��&�v��+�k��֎����A���n�j���I�Ǫ�e���v��X��
ѷ�o���j7��r��u�1�/���KRYjI�]��� 8l��܇35�����[�q�93�V�뼛\;@�JP�<*�f�)�4��]l`S��H��sK����¬O�����c鰪�7�5:�I�݋9[��b�6б]ו�-W=��,������0�Q�%z:�-��o�R��ݽ�s2�-��ZeX�.ꋷe*�n��Ev^�Ï���S_�X�ʔb&�u͍�f_t[���]g���G�]���}�u��.��F6	П�U`���'u�%gl��*�R��롥Vt����&*��4�ّZ�Jq{Yj�J��Æ�N/%HTP)4��ݴ��ͧ�.�w]̘�v�T�Bc�C�Y+:�,�[�%�	wJ�gU�r�\r�ҠE��%G���Ȑ�ς��I�f]��i�ۚ&�5�JSE���N�K��hҒ�+2�Y�K��O��wt� U�N�;�����YK�v�n+�2�@d�S�I����W;�٣Zh���I;zw>"]D5m�v��.��)d\]%R8
f�;c]�4������������w��]o�]�������]\��>��OH�mj�Os1��վ�6o��B�)4hޟu�56�����X ��cn�� s�G_9�:���2'.���	���TS,cknk!m����^!�м9U2�����n�o�`��;�����ƈ��נ�nȮU*d7$'$wY��ئi�rWh�\]�Q`�Oc�_Qk&�ëc�Y�]]w�so4�8��l�'D�C�����c�/p�h��D��΅5hڹ.7�7z�.N�`kKSΩ�T���	���
���\#���S��yEo�L��T{s;+�D}����j<�B��ŮJ�P�B�#W���n�ܽ��Uu.Z	w�h��Q�e�s���Y��LY��8����
�e�a�_vn��|�R�u�����q��bH) (H����A�����/z법B)�]�����n���%��&u'��y.���u��G���v�C��oT\�
7+f�N���,Kה�D�Q��I%]ͤ���"�9N�M��A7D�b�[���*��'q[��IÜ5�])�6k��o��s�\���������9�΢�^]�Ü�� |/`r�wz�䗭�r����2���
�J�r�.M�+����]YJ�:�gwv��D���v*���4v���/��ٓl/w���:Z�찁�x�s$��]^�Z*v�8^�Z)/Z�GҮ�n��~٘�:�iY�Rm�y�w�A_E]�\9yI��'l��}�Y�zV���=~�6s�,��r��2�r�Oy�#w�qLK���O{�z�Zp�U�A��梁����^�<'i����8aີ������������kSh����2j�0�L�ĐăKҤ� "#�@F��,�P��5R��e��rK��n�M#��Ù[P(&r{�\�����ܮ�2^fFM�`�\G��n��c1,�hN�3���Tp��t<+�+��$+xV�)o|vy�&���@!���o��^uvz}��w�(f��Ff-\�N�E�U]�%ѷԸf޳ճ���[������S��-Z��1Y���"�d$v�����T���9��S����)�����O{�ᴐ����ݹ���>;����f�9n����oi���:X�%t�!�-��V�B�T�"ާ���M��O�p�o�9c��mbCGS�K�[�:�m� :;èw&o꥚��34>��QR������>�����ly��;�J����v�_Puqn�o�pz�
��;����u��}V/�"��4��ݫ��M���E&yzq�:�jo <i�[���,P���wuq�q:@㗼x��}��؟\z��Q�ꯁ����=��y�Gss����Op��(w[J�=o�F����{��4�5x{�׏��灈BOy���zy���uۤ����\��yw.�:JwZW6K�5���R��Ew����o�B���		�s���$�$��o��O�ߺ��9�`���h�Y#�Y��9���K��!�.����i������Y�{oZ�+�󘣨DXb��*+F=�z���Yr�|H�%.����c2��w�3��=�c�D�d�Ϟ����Py���sҸ\����������	�W��s��ܫt��b��A�������r����B���m���:0VTD�LE,����4@�Bf�D?�����J�j�Z\Wpj}Cv��(���ѱ��1�r*��Yv�R\r^m��ۊ��C]MK�� �%����t�M��\��<�F�&����|)+��U���^��^~;<�z*P����w��bњ�� ���\WY����9ܷ�r����@y�����9��4�^j��@^�}˨p��	Jۋ��C����R����G������N��n��}_}8������\��J�Cg��엻��Ofj	Z�E�Y����WUWfC�e�^�x�f���X�4����UV�wT�w�l#+��#7���Z�U�6`�
�g[8P����֪�F�!��Fm�n��Ğ��$�י�{�;�����7�%�p>�sh�igm�*��d�kt>K,&7�|��>��\�x��=�O����R5�����>��le�������湙"�E1c��� ���VʈUE�H�V�Y
�°Tkcm��"2\Dw���5�����1f�{�1��},�G��X�;�ݘ���{��0�u�*O����r�t�	�s�I���
f�(E���Uiɻ��s��딹F�������U�s�ǒ���_l�J��%�J˗��U������ ?@�w��D��}�}h%��3hp��[��_.�I������Q�'�[�]Kȅ��wդ������uP[8�OR[{����+h�bcӻ���:�}f�v�x3�EN�!(����ƛ��_UW���k�׭~�?u��Yk�1�N��w�A����Gl��Z�ri�+�q:ڞ�~��˻�W��}�9J/I���i����;r�g:��j�wv2weq`>�/w:��9=��n�$�Đ7�y�<�j�x��i�n�U��[��Q��p؋o51�Æ���٬���(~�}B���g��g��Ԙ�,���=���D�Y�L6Ⱥ�*L����Q��!xzg�w��X\�:�I�����$��Z+���C�`���9�(`��m�>~��u�$5y�~����띿s�OWGI��/yY�y�6iy�n^Noq�Y����ѯzw�� xr���|�ӿB
��L�����$u{9+�+�=�v�����=F�7�X�&�w|ӈ�����]�߽c�� �d�u���{�\�{��Y��o
�7,m��vՍ�V��dD[�6�v[�{1u���!��0>�{� 
��ڗ�}m/f<p�a���k3��{��vFc��W�^V�G�70�fM�d�ܫ��W ��y��[/������/`E�����jܟ9�۝�a_�q� /sr�8�g=�s]�7� C�ԇ�{�u������C���o��7竚��|�Q�n5�jG&�R`�H,X�­��{�i����a�9�e
!+�*�tվ�ر+[�vJؔ�����W7�{2�8��<wo��7���2Ԭ�$MS��K5j@{'u�h�ml+0���+��r�l��;1p��&���|�߾�| �{���Mc��NɶaIқ��h�J<U�I�����x����)�
�3�K�_�}�3;�9��g���|�g7��t%�ϟX�Z��6��h�cu�_]��g{�u�I$�I��z�ߎw�� 8��
���ޗ�h�7ls
�!��&�M�B���>�;+��j̽��ւ�_/|>�|Vm�r4�V���R<�vt����롼���T}�(͚��z/��XmY[U}�WaG��̙`��Ǟ_�I&@
������ϵ�����]{�M{����Ԋ�Z���v]-N�M%�<�<��Ώ�y���5�{��~�32e�#$*R�*�J�:5�|��=�`��恔t.7;s{��Z��hhKuf�������"�Bިn�+����0�dr���]���2�a���hBɶ�=7��f��1�wsF���7������mS�bf�F}:�u�N>�����ZZ��9���:nU\��WuP�DO9��K����V ����Ϸ��uu�8����9��ߕ��I�@���%Z�#������*�Y�bs��T����a�ַ0#6�Ìޙ��=�cO.��}ߚ�g�=��xc����}�){Ͼ�H�^g�L˧�˙s$��V�0�T��^���۷@}@�o_L�W��s���M�eK�]`'��0A*�������^���f_d)â�o�ڛ�ˮ>>_<���O:>�:C߅U�v��ޜE9�t}�ۗf����oU��N���w��˯��wK��D@$��/��i��B��W۫�N�'�-t8��30ؙS~c�.��9����*u���9AkD�$6Z̥�݈L0˹��8.d�EKR5򆃍�$�&��ϥc��s8��;fw;��O m��x|u�>BBO�����ݘ����$����Z�wk�����4��оP��P����W�W�:�<-�_�W�w�:�t낪]YBo�����8�r�>
zĩ|}~"��e�=-	Ww���[ގ��7�| ��u{bf��-�M�甍��:������^�%C�{8ضd�Y�W��М����� s��'�܇�{�����_�g�2^��os���e����6�
�u[|�:e��������k/���<��I$�Cώ���������o���zƫ�������{ķ���Ս�'Hf�h��j�O��!�\R{�\渘�wYd��ˠ�E�+�����:�7-�L�b`�U�U�|�q[f��*�)�97����i˳�:k|m��nW�S���$��@���k^���(��zl�z���g�]H���E`���ڬ�.ؾne��ۈ0x��F�h�[�8�K�.j�|Dc�E�m�b,UqWT��+1t�;�����5�;��Ҿ���l�g�}����@X�b��Ӥer��;�|�f����,)O�-wB�����?�ʋ좾.���S��1-:;�\�&V������eZ��":��E���n�b&8��7��)P�Jx�o)��e��)��w]�5�cv'��hk��tӞ[�6o]�����0�yfQ2��W������6��F*�T1��Eu3�6.1���2�M�6�nw.�vݚ&�Ű�NF�W�}��AQex���J**�Ӄ�UĘ���Zm��  ��F��H:T(�/���Sj���7���t�(��ժ��W�i�Vx`H�nĦ��t�0���\��V�����)i�e��!H8�h�D��RsAďĄ�l)���P�-����'-�\�<0���|��c�'Q��"Dw����Q���ٰ�Q�Q;)��ɚ�醴y��{��z�!'RIXJ���X@=̙e�<�PeHQ��p�����|ٱv����:KK|���KJ�]��N��˖������h挚BjӍŦ�8��R�|���o*���D|�7}r�����3�++0]i��3*jշq�]|!ԵV����>��r]�uݬΛ�V]ډ�I�2Jj��/d�������vv���q_5�fH�q�b��:v]P�ypצb�w����L_z�����ِۙk� �O�Xr9e��[ܝ5`��Yrvz�I�]��mLO�
]wE��3H췹�֣���4�7�#Rq]�S���5wm-3wV��k��	��L/�����ᇞ+M�^L��:��9���װ�j=����#{���&5�PO�7׮��]�7ܥ]}���Fq2D�,�v���g�9S;]�2'�׌��3��=݈�'�
_@�F���)�������%V��{��IO�'o�s¦�7:��<�d���w-'
���>�;�4ݫ�$���l�\��"/���j���ݪ�oGN�>��qT�Ϙ�N%%g����n��3n��[�̓�y���@c��c��.��0�!j��]��gX�C���Gu��͹�M�l�S'o�m-�"*�]�nN-WZ�)9|�3��Uu������}x���AMZ*o"{T=fJ�Xz�p������4˻�-q�w_:��f��a���:�[/�Mn;�4gP��0�l��&�������gM�d�kV�j�u�m6������y��_O��u]�K:Ζ�PX�,��vGe�B��܏h4u�ь��\LKj)g�˫oB����y���Â��_����f�s
��9&����Hd��N��䒤�I$�I$�I$�I$�I$�I�C���s�4�_=���ԣ�O�lv�v�ݴ_=�=˝���Gk��db�r�����ϸ�@���78�T�r\�Et���,��@�cV!̯���T3	��kp6�؎~L��Z��Ӹ�J�2�d8�1���|��y���� H>��o�S^��=S�. -1;ŮO�s`S��y���"�O|�#�Æwn%�zSu1"U��1)�5�횼}�� t=D.�!Zsژ���~�6��J�SI�����o�VE�nuI`Xt�S >���o#�{���ӿ?a��Ǌ�I")"((�!cI �,�d�YDP��mȻD,�Ӵ2D���}5�'5�ڗA����YCMj��E���C6+�;\
ki8����C!'�9%�� �����,w@���]�௜u¥c��ڊ��\3�L'G2zU���e��7�hĎd��� �������Q��C4I��N��Rl�,����|����|< WX1���qŉ1+
�ź�6AP�VhF-46�;p��b�
����`7�Y�>���9+��6��>��ɹ��$�u{�FbH�`-�f�#.���Bȧ�RA@��n7���2����p�4�s�]��1Pn�Ɏ��Bܽ�"�c�Wt��d���<;�А�Wv�;��|�_���y���\I�TN�B�����Ӱ�\�8}`�4�'��j�Pͦ�~�����0zq8أ������)OUmx�*mR@ݨ�Y񌪼�M��+1�d�Lt��r*;F �-�hi9/���Eb~��p���U����}�h�|�G���v�vJ�{1}��`oj���M*s��S8M���}�a���Y�����g�i����I/d��o�\M�U���6^�L�cݾ��H�_�iP��u9\s�*��-x�\a`7"TY�3����b�RY�}������ �J�R�9�t�Ų�d%\�e��k���"�m���-�5�,w�nY��z�<E�ߙ'���_[�>f�T�T��u��Rc�L�j!s���ù���@�g�@��u����LXi1�a�O���<�c*i%gRq���:"�<�����M�PyC�N�?'�d�~q&$���O7��]��fι!y�T���B�(�����-�X(@��s}���{�{o.��{y�]Q�PL��!�����5�ix*�0��zOoK���v�D��7ޤ'���x$İ���Y�>�us��]_����q>a=V߰�5���'��OP;�ԕ���<O៞�<�AC�1��l���cY��ߜ������Z޷��==d���I�Ī�z��U�]�u����|�y�~Ѥ�B���i�'�|3���eGVHc�~O����z������a�q i'�z�<M�d�O��$�q��d�7���HA��0����x��+'����g��d�,&�8��f�����}�<�>��6=�=�j@���@�ޓ)3�����JU�\š�| d��
�yR7��pL�h��|>�z!>L���Mi�݃���*��Y�u�uS��۪�F^�r{Ւ����j��#D�v�n>7W�j�u�gM����;p=;����I���Є��s�2��k���oQ%�Ka��N�*X!���cup׎���;�m�8�M}�摙��}�5~R(-xw�>����D�� ��}C��X�ʈv��Gꫤ%MA
�5K��4�:�O�Շ���kc���z�T�#�{:{x�6�f�K:����
������U�.T�'��ԗ����-��!Y���^�����Z�m���{s_`�@ɢ��}���:ƿ��X��(����+;�C1�q*bٴ�T�,���0�URI.���eo�y��82j]S��ca�ݝ���#�<����˜Hi��sb7mnjS.Z�=��		������C�|��C�{�����pv�
����:s_wk���Tϡ�xr��5E1�}�`dAp��[�UI�}����iÁe���uD�N_ ������ƶ�Ma[����pT���tk����sT����_v8c7��[���'�	��i� �x�����{ޜ��=[E����`�B^�a
`��߷;-y�[�;ېy̐ժ�x�$�)&4��ٖ!J��Dʱ!���_zg��:��Oy>@�}��k=5\l}u^�qe���w!�*8�?c��T����$�<��Xqd�����}�~�k�rv��1}��i�{�/�ߧ�!5��ѧ=�������} }����Fp���
l.�Tdq��)�f�.?m�������,�x3u�n}�@���ƶб�	P�k�;�~�s^��G	�7·ctFT=�f�2YPi�}0s�E�;m�7W'NFsy�zV���!�wзns��
ke��U�![]%��>����Y��2���!&��̻��}�����ᦰ��s݉�9Wm�㮟�Dd!4���*�$�KǕ�QT�^���H�o�̫�����9_$��Fg�9����������K�*��Fc-Mǜ���ђ���1�o}�Z��a��� ��C��L��k�o�Ad#�럈������M�$�ֽ���ϯ�ǻ���2�O6p���s�mTS����J�k���d|F�A�{ެK��
ڔ�����y���tu��q����_��~��o����:gՕ�>l�I�TϨ���:x������v�nWuumz�`·g�.�fQ��˸0�:[!
~��<�7����}0�9�j���ٔdU#������ռ�f����]�kT�9����]���&٪����Mc?!q�Dρ��["�̼]dյ���� $A0X)���D��XDE yl�<A�iv�W�x�Ky��F�������~}�����e�5��]T�XPTXL�R1�kEt�1dPF�(�X�e~$o|M�k�֟p6VзE�s45�֞���ye�.�ӷ���<���5"n�������Z��=R�:9��7<;��JX�b*�Y~�����e����W�ܐfwګ%a���1���HB��kO}��=㭾��?��97����綸�a�����p9���LE�'���9�N�<��n���K�I/Zx[��0'1��]�߾ ���z&{����J�J^o�/jZ�N;��.s1�!��HtZA�wg_��d�u@ʳ+C�%��}���N3���m0ĩ�J��{tՕQ�����l[+VX�>H@�b���#p�|�KZ�/���ZFͺ��ۏ�~��?/j�y�_�
���~�?��y�}^"9��퉎HċuR7л*�{A��I��~��"%]o�o�۰6�m{��x8D�K~<$鸟��p��B�ӳ�!��������<|�/�]����V�|��C{N�I�7�-�6<�gpW���C�e�ۓ�8E���5[���ݕĒo��~���{��^oZ�8�J	!*�Q��~��}�����q�~k���ЙV�ӎR0��י2������1^Upv>�,�특�wԹ���2�a��n�OU�ժ��~���ӡ���ya'<|���ٿ�'���9�CC���$^��ٝ̕�<�#�ṑ�ֈ���[�7�$�E ��fDo�yN�7g���P6z��Ǹ̬��lɖ����>h�'��Q���g�	>�=3}wI:�A0Ra}��x���94}F�íR}$�9�}���0��.���
e�^]M�V[��N���k,��� mh7��jsQ��ͷ�)s��>�>���W���v�А��1�`���0�p{���LO]%����',��lH�%����9-j���g��L��޼�d	����n�ǂC��c!�"{�>��B��ZŔK;5�7�0���M�4B��Ǯ��JS�3�#��<D>��22]��K8� 9���KO.>�#¹�a�����P�U:��7��L���E�D
"}���=��	�S����>#��L�C��?D#��sx�3�푨������y��&#z�m>��ۮ��n��wG�Rv�o43�47�ov�Q���EX��wzA�guƜj�KP���[}{
{���-��{���7t<�f��@'�!/�ݵ�˿<��[��v������Ꮸ_��m5c</��7R�}�!��s����
1p*���Z�.��2W�L!�{ޠ< ��\S�4##��TJ�v�oaZ�Ǿs�SIj� �Ӫn�L�WK��jR'�sD	��&�T��c�>��[�<]\�{�[5�����{��,��TZ�Sܸ���KCp�M�.���d�n���{�2�5$i��� K!NN�N��lTc�~s缀�g�$�s��w�'�&}���uM��Pw7?u.���U&����%ゐb(�~a<�8���B�립���RC���Ў8��n�f�;8����O��#�+߽��YY^��3�#g|�+�%w,��O��6eSf-��?����s�����ӯ<�����^����
T�W���,��mDU�H(��{���kZ��3Z(���W����{V�;��|Se�
��D(�_�6k~{��Ξ}}�/�Yj�5���FP;��\�,��^�q�c��G,�G ��&�����04�ټ4[��6LK5O�M0����*���uUyV��F���^���:�o;��S���5�<��������
y�s�� ���LJ:U�M� b�G#�;���_�>o���d���"�����
�%o�z�Q�fck~$%�0!���x���?�^���Ow3*�YL*y�y�"����O{������$��;(~���/6����a�k�+�N�*f�-3�u���Թ��7-~o3���I<O�	��ل
*; H4G���y��`�t���U��8x��b�ٲ� S���o�'4+!1�A��L��M������Q8K�>��o��럥���p���5�}���� ��uDY^�`�-9������iXm~�Y�x�_L+]'�o�
GG�
(o�'<U��rMQw�`�G�73 �:�~�ޅڷ.4�����Y%�r��>���׋�G�����S��D�+DF� ���y��h"w�[�g-�M�M�9�9���wY���Pj'Ζ<���k%m���
�{�3~D�|��;Q��X��(�C�4j�s.�WXbR���
aRT��L˄�X�d*$ċVE��ehىZBAb0�Hb�"��莩��3$"��-Ǝ��P"��Aakb�9��|���k2���.TY��C�ۻFĠ�!�[��z��-�2���MWgb5�I����7��_^�m*���21C�>c�V��Uڙ�����/Ӝ���A�Mޔ���V�v��On���Y�o9�#�%����'�{s,s�uu�Bw9��>�y���~���n����#H�=�L̫�>[TݚI��*6��� �4�u�`������������R�Wǒ=��m�yfP6��vh�䳆+@���J9�
�G���=��+7.�8��RZ'd>�ۺ����#��H�`�誛�U��/菣��uh��
�&�W�y��T�/��|��������s�[$0L���W�4��X�P��dRx��F\q�����ך��$��nEw��}�;(�ᩍ��Eg7���ҧ�����W���~K�� f��fw)rߍ���R�,������'4 ��:^1n�N\�XȽ"���g��'����Ap���86deɢU[#����&�}vk����v��4*�����W��qL��O�I8D��.�?t²b�@��^����-�c�7g�1}�Ӣ�;�{/���0?j�/%��j��C}3���
��$�y��ΰ�*��{:��i�{��d���V�'���N1`�nV�6�n���|0h�UHƁ;I�a% �0%ؕ��㤛a���ѭ��r�[�W��u���bg6������e��	ru:�M�T�-�=����ao<���2�,n�$��I�5#���Ss�*�Ɲu��a���I�/_w'a�BB���1��H�����H"fJ`[W�J.�N�Z*@]��d�	!�AH���8��X�b��7P�X*�ph�&����k{�yӷ��}Ʈ���s$��4���^
*8�2�U/4of���F�ʥ(P� O��)��h�W�ެ\�3g��w@ַ:���su�κ8�U��Щ��������)�u	��7E�;�1��&�X%�Cf�D�Ba�k�j.����W|>���O�L���#�*Hu��b1���v�[{�2E�VC��O<��l�l��yoa�2����@</0��2{i�����`:�}n�c�R�U��0\���1Q���8�-h�i�1%��k��&zӏ^�CJ<lTY	7e���3��m��O�$�Ӣ�8��Y���ae]W!�^`T�̻{�����Lrڥ�sWs����Y`bRԹ���=�7�P�]xp�ӷ/:�l��6Ҷ��=c�-ܸ!$?5ğn<Z��֯d��n��G��Hd�9#��� �fiMe�x�t�(�uo���u"5���o�v�1�݂ᕛݗ��,c6���l�PK2d�\�'Hq(s/ 0uL��.b浱t��fέTOi�ƹoWY�{��[�����-���"�>��]��*3󊫻i���W�{F�̚��!�3��"y�n���n֛z�h̋��]k	|�#�~1#F<B�v�X�;����x�� L�q�&ɯ1�Š݇����D��&�T��)�;�hr�#�y��ۨK���Ue8��t1rٟ%)�a���zwc�ηd��Kri��M�Q��jII]����^��rY�[�}Qev��G���9�:���Zw� jk��œQ���73H}�wj�˥�yM���z-ow<؊�����R�c��h��~]��F/�ya,/Ϩ	�;D��Rl�����s����/�:cl<)"�N�u1.�N�w���s�����8�����g�͗�x: ?�G�6�����}����h�!sk�FKϨE3�j�H��IgH^Gf����f��.��_t�vԲq��'xNxma��bzy_^��b<��	<K�"��;og2�|�em��'
�ws������z�O��T��w�e���Rъ�5w�q��)�㊸n��P�9*v:	�9�Z��2�ZB��eby
oN�'�^��W!�������[�ָz�&�;�2���l[��c-�����[���;��R~�C���i��9/@�KQiޔQD��q���m��y��x�.g��r2��M�2��AA���\e<�,4��_����%���_UT���L�o��@|)p�~�]���'T)��V 쉔��z�7�Is�!�������s}�"y����y��N�Vz�\Xu?�☢u2F&�ry~.z&�T�5a�9�>i��1�?�$�5y����=��o�n����&8
�y��w"�%��]��i�b�O�#_U��q;nj��x�Hk��L�s?���H��f+�5bj����ʋ��g�/��9"�G�T�&��设�����9Z��V���
9��	�R�*���U9���C�z�N0���.~���N���95�3w3���_���}��Z�d���� �9�� �;��A~�4�}�	ʤx�CVc�ّ3���(��++��]�3\�6�ǥ�J�§KN��a�h���g��ϯ٭�ߌ�Zկc~�E�r����{dϹ���!ALY.+ؖK����7��f(f\�"4E��F�6f�m��U��DDDq�+��1QH8ZȰ�Y(�QF�m�F�b3��C"0QV�%��4[�u�=�/|bd��Wsf7�(�_Ho#��N�ԋ�� ��b7דUn����b=����[4&!Z�&,7T���W$�a�r����0uF�U3����<�H�r�%&�,�|W��'�C� `#{�TI��m.�8:�هʢd�z7~�o7��~!/��������9�~J4�w%B��m�1՝�t+�8q{	JMЃ!A���*`}!)ڳ���9�#�&VI��p�g,3@p�^��]a������}�s����5��?���'��d*��(�(v��.��ʱ�K8'���cGTZ�i熹wү���.娮��)"�xo��ۗ9���[H��I�j����r��$t��dg=`�E�(�~a�J�Bv����!zθ8����?ZV-Ǟ������{c�#lΒgs�Q4<�y5��V�������K��$��"�2E$��!�S���)W�O�wH���s�ߪ�|F,��ω��f��W��]C��Be��j۪���#����-�E�\H}W�<�$*�0s9�J�s����P�s��Lt��B�s��PJ��w��ѩ�خ��4�;"wA56�*E(&ʲ��t���$�<BI���F���Y�'���6lQQ9b0*6�ϟ9t}�;5V�:C	�Iu�Zz؏�r��>3q��,��#�J�OEz2gd�z��Kb�sgc��y
�ץ��!G7$<��H7z�5��w���5�ǎwW\yһ �AP(Q@��:5U���.{�F�>�gZ��@�)e�<�U��ޫҞ' L��S��M
�0�=�}RC;�}��lǿ~��޶w��e޽�h�h�".C�[yWVM(&AevA,*��ܕ��ܺ*},�iҺ�xB^����V��^m��T�N vT�J�>�VAؐW&~WoU�"� 7iH�&�U��2�1��Ť��S���	~&9Y��A� r-�v�^����)
R���Y�iMد�*��fl��>���(HCW�־�����̻�R�02����}�Ҥ������V�9�d$�P�ѽ+���x�q�Fha�O���>����{=78\�5%�Ր��5��'ߵ��|fu�ݦi�{��}��Ю!Us��"�U�s��;��o\��k�V:��e�q����r�ia_�9�<B�����x7p�w�����ֽ׹o�޷��;]o�$��.g�9�g������K(:�����	3zC⁉�۴����r_�9L�-��!(� �)���èVJ���m7�V+-�x�p��h��S��<.L��1����@���3[�Iup��h�9���J9j��^v�+*�VP-�ic�S�,��w~���<сP=�6~@ot��{������{����w���H~�B�7$"�Г���y/�ל�MB�"�s����)@�ǵ'�����';pp��i������X���˼ � [x�G�v�g{!�{Ͻ[b6m�BF��d6nk`<�5f�3)x����kU�u�]��a������O�Nq=h�]���:���Ù�L���0ԇ�-�����)������G뛸.r�_�5�|w�l�/���0/.Ǭ�ac��R�H󇿷����������ҽ�}$$�߂C�J�X��K���g���P+�O�����듘�7�X��e�o:�Rh{R6ε�Z]�2��G�
4^2������Et�um��z��+���,5:9,'P��,��2��죣��G1X�pGD6n1-�w؂�u�m9�;so�|'~ߟ]cu�3}>]P���3����!�1�p��Y�šX,�db�V��E�@�(�Ց��R�#�JFX���ʑb�+��Iah��TR(��e�p����"p�an��M�m�H�i�ۗةm'���[c�e�F�p�b��:�\Y��i��[��Ų�K;W����n�̜�E����(R]HL�pTʨsiu��L+���vppj"�����k��#�St�/�b�V��W�}Y4�k�O��u��]a�UD߁��q��1C�:3��̹޳Ӄ.��1a�bk�dތB��ϒ�d�m��p�k��X���C��K����o��5���3��;8BVn��y9pNpw]3�)!��ۖ��DAh����������$N��|m�:��/\ｺ;�5q��E�7YֹTxا������a���Cp�ի7���T��Փ�P����,�"�>�{ݧ|d=��Ec1?D}���{Sh��lO<'!q�|��'��f�&rMq�D![���O�Wp�b[3�L��ƭ q�i�*�!x#U�����_�����?2A��Î_��D}�����<��o�8�� k��T�k��Xu��H5���gBnH^>��~�g_�J��eF1���W�<D��.�K�p+��7�[ώ����b���7���{���LY]��f#Vw��B�&W+����W��m�"�D��ś-�3���6���ZQ��}�f�׈u[��/��?�U|�h�J���@��jӪ�����>�:X�&vqL�jBb6p[Bb`�
��ڴy�'�}���sk�W�7�F��f��>�g Ղ���?P�[j�:��@uz ��gk�m�/��	ܔ�	�$(�h	i�Bf�V)��^�w�K����|~X�F)�-׏�2<l*�h��2�ޜ�PA��@F�}1Z�s�iO[p�c��y�Ț�v�}9�.J��Ѩ{���o	���׎��O���{}r��~�����c���S��yZ��P�Ɔ��E�^1~���suZ��	�h݆��Y{;u�7�{Kp��\>� Z�dd�A0�q~\n#菅�޻����}[A���Q�wR�G*<#0�Ŷqí�����,�m�3�=�OA��a�3[qw��F%�,$��Ų
6M��Rǈ��~�Q�`8D�)�?GĀ&7�97A�ݭ���u�N5$�=����0d�� #�@KMYr�㖬E������n\7�����B��r(�6V֧�3��q����|=�vS�eI�<Ѻm�xэC'��9u ���;iw����nq}��d� �XQ��� D�C�M�?r��~2ǿu�3e�a�宙���I=��}H�f�ӛqr�*Sh�U�0vEjqL���� ���uGk[v��Ւ�8�4�����D�,8�k��7����ҜYE�n�a��j2���$̾�z���a��w�w_=�8v����ܓ�K�{�׃�@�}�~�W�+�W����/�R�^s0�9��Ѿ8�!�k�FO2N����\����j��ةQ2������_y���1���pϽ����Ry���T��{���˽�D�����O�gk�Q>�WH:p�1{�1�y� �������y���}{��<ܓ�'��kSA0��y�m��\��h�V7}G�!Z�s��E���*�8HA���際�a�$��X6��"#��6_4��¢~c ���^w�|�t����]�{a�U�afLb�������7��q��q�G�h���Q�9YC���1�t켉g1�~���k��Hb�7F2카�\ҪCP�z�)�~4����7DWu�ӹ�|,ߡ�P�@���ɿ~���'�۸�3�Y|ْ\������<�-��j���KƁ=��D�����������h�8��Å���DFM�����������/����^��h��!�ݨ��$uMf�B��=��H�G�}���߇�5����:����!�u�b���l�3/fs��@oO��?��-�fev�m�d�����֍I�F��.�PS)wgn���m��ʂ��!����ʺ'}S2|�H{�3^�f����~'�q>h�G��BҰ|�=��f����X�=��k�(��`12��};|��m���:ڜX|w@�m\@����!	����X��k���w��/o�{�`�If���ܾ�;$i{���C��e����}
L�ٙ30(�1PG�I#�Nܔ�hm?,]W��1��(s����;]�a�+�\��[j�iL�b��\��c�Qއ����F��z��j�,��r��b��z_��ѡ#����H�}����}s��c�k�ޥ͌����&��&��N��"�3���L�'v��z�7��,���(~֙ϋ���k���P6Ő$��@߿]fVL)h.�B�@[eƵ�{k��*��e��w^�wCA6V`���M��\��p�-�Lvm��j�(�
O���H�E$"��>}�s<��~����3A�̓����s��-�y��SsLc���9�P���==�(�e�'G�}�"�<>��Д�D}}M̧�=p��E�I���kScf��%3�;���k�ݟiޗ��'�5��1�]	�:56��+�^��YΝ��D0����5�~�;7��~�3[���nm];���ȿF/�:��b��J�D�J���Of^�*Js���>��uP����w�|WJ�c��	�ȩ��54;o��]8fo���1ա@dB�fۘS"�A�[,d��-l�5H�T�Q
�1��B�,�ZX1��"#�%.w��u�����FAN����Į�>�݌q�l���3S)9ô)\��Cg���ʬ�Js��4�q涥Kຯ�O-\;�E�rI*�eR���~��OM������sl��P{��E�1�0��ڟ|�<��)��a���}@������ DU�R0U�u>�p���o���gs��UZG�7��c^wi���Қ��*3N� v��9�'Q��W���tr�y�|��p��ys�t����\JL��x$����Ǒq�&��ee�3����,}C��έ���aʐ��MU̵1$�Q�m�u���1�kynEpI����>�J⯫�(ôV�l)˛eW�>�Ɯ�;j��Y�v�K�Ǭ�c�	Z���P��Dp���������y�@���o��w��_��/y�����5�Î��T�N��QY���S��;�"3�m'�x��o5� ��CIm�����ux�U%����H$�@>$�=��H�cH*y�ij�<����r��Z0�AN:f&��&83�d>3r�$�/��⨭�A�uW�"3����]U���ֶ�j�w�ν�	�q鬳���/1�{NF3��w�
x��;�B��}��gE[sOWe��\b`�iF���~�8�-���P�����}�7����s�糢1o(rk��pJuӳ��q�M�e�Z\M��1��b���\Օv#$bPSkF��j?�s1��-g�нq�7c����ھ�&K�#c>i��7hђeK31s5/�F}����;�s}�ـ�!F/�d�痞^]m�`�dN����1���#��+�H �Cj1)�Љ@�(�h3ff�mИ�@XL�hԻ���ƌ�湳PSb�w�[��i��(�E��y@�~�� +fI$wF&�!�w���SoV�`!�S���a��b2Y@�(��w�s�gi%��Z��рQ4���_��D23������5�>�n`��@baG�H��'�FY.��S~,�4��+�$1����K2ͺ�Zv��OP���ᤊ g&kM��V��3���P�^Sv�)���w}�9y�L�sC�|�4�
F����č��"��Zu�������^���\]ʴ́n
DTG��4�A��Tvf���\��ɹƉ;�}3M�x�+)[��í�S��b|��:�V�[B��Ǯq��6�L"Q�m����_J�A�6}u�d^���&a<�B㗾���Q��܂�4PY�.ˀ5l�)<U�,��)c���A����7Ȝ�S��qC�{8��Mi^%�m�b��%���
����+��gk�p�ʺu��)�J-U�%���嚲�^;��9�J��l���퓔s.����wC��u	9O!��
V�Wd��f1�9e�[����+[x�׆=;����݉k�3N��į��-��颛uZ��5��l��L8U\�wW	b�.Am�Etk|՗ןp��n����=@q�r��h�6AG�P:��3,\�nboY�oVC;KȢ=$��I�.���ޢ~�c��uܤ�'�H��m�X���V��Noq�K� ���Ә]�+;{Y��U��ٳC&>�C�u�XTn�wʒ���颻���N����-iq�W-^�"��jh�D��-�F�ܗy�f�GD,������=���&c�=J�↬ �~_\���f�nv���#̹�>��6�Go
�LcejOh��k2�n9�I��$�[K0���p��芾ȡ��V�;G��LmFF����f�	���[�dNQ�7R�����#�2Ve(�U�$��w���2���E���Բ�:\,DUu$�I$�I$�I$�I$�I$�f��]X{�F�0������U�ӵg�]�o�LF�h��V�f2��D�D�+�1;� ��e��w]A�*��e֗��3�9��h�_s�׍�*+ƈ����jO� ]��Ō��,*R�?z���v>9_�s��a�r�,�Si��<P�\�~�aLi�� �I CL!�}��|��������E@�<�J>�\}��z�<�c�5b%�"e�*��=.e�%�7	hRbi�!L��8lI�g�-߽�w���).gyܞ;�����U[��@�!�:}v���MH�Y�_G�7�� �[��ۈ2l��ѢY�wI���l�Tb�Ͼ�y��W(��5}sԐp9CݿG,����|9�'j��r�^���+�%�0v3�P��}�]�>�vj1x��i>Gh *��Fs�g�jʀ5�
��z����/���np�jwQ�5�fQިy��δ|��naڜ�ʤ�Z�DWO`y��e���m� _xx{�Ht6&�$�M����6C]N�Ǵ�_{�T\����\���6b&4��堀��`�5���?4_�M�\��*���P���E����f�A5T��=�*��J�8�����:��S7us����K���J�x���Ziզ}2����7ǾA�N��N�γ�uF�B@~�0s9<>�׺�]������ѸΑ&q����#]�1@Ee�>&��r����0��C~)@S�� l���QoB����4оU�H/��ĥ�V�]Ú��c��(��~4��C��݋���*m7��ʻ=}Ϲ������z]\ֻ��5�������]W��>�ޞ�{>�7���Љ�+����h�0�_e�z]���c?'��x�<���R6����'������7��0d��Sӕ����"�gf�����+Y�;�:��K��n�h9��i�g�b�[G� ���oi��H��%ex�S�+����4�}}L|���cN8�R�Hޢ�1�D)31Q �Ї���f[��^n�;��_����'狨J�u �:�^,נ~ @A�@F�y����d��0~-�_��)������� |(���^��~e.�u�U��yȽ�{S���0�<fi;���,�9K�Z��³���M������l�K��4��*��ꂄ������7w\ӓ�����/����m��N%���<w��G�| {��ɛG4y+�I�6��Mg=�y�h��{ T =��u��kn�Y�.��*�2���0mh̬g�/����A�
L�:�D�GR[������g�k7"��z" wG�1���E�F�%G`B����WaN��F\�+q������B�U�S@M8t�C�ru��b`	:b��)�S#��?C�Աՙ#}�3d߽�
��͢�U�{�[��UJ�1�B�Qv�j���#��a5�N�����Y=5��駙^��.x�{�>�����/��]�@=���9~Rǹ.��3ra`�ȯ�#[�Wn�y�1o.��ͳwF�|�ިl��}�8�[m�����ٮ��?(1 cB1G�f��T�� �X��6�_gR��D*�t�N��qK�����5��Ac���w)�O��>��λ�>�}�L`�X�54����&��\� XDCVZfb�2�J�C�OK�ӽ���^r|�j!Ɲ^%+�Bu�%.�I�|��n����n.�%���HQV��61M*��驀����zf�V����>Cp["y�o���$,��o Wj��7C�jT�P��HM�G.E���.�K-��YB_|=�.���P,�Y�x8�֑(p"�a��ko�%g�Ƞ���">�}-�o� �V��j񆼢�2<5��C�L�tW�x�N��'�.�s��'�kҊ*F��]��l�+V�V�4�����}����w�K��o�r˭ɵ0�C9Qmt�����η�oWʥ���/��gQY�+�����
��#���� �A����-�.��Sl�_g�L�o�=�Z���F́|�P�ĸ�*({�e��0=My��x���������o��m�<֛|����������
QI X��i~�y�y��k�`H	U��s�v~O�\h��J<ի��?z�78�/�;6�[U�*��N׼����G�.����}�x8Pco{��!�*�a�vpTU'�\��Z��䰖��ɩ��L�d�T4d"�&2��E�K �˗d&2�T`�j"��
O1�<+�ОV�F�n�|�d�Xu���kO���Si��g-�뱟E�ED{s1�M9,��q��)����F%�fS����V`\�-	��1n�[�^����t��t�� c!���w�]��Gnwk�?I?u�r��������v>����.x��jH����}]!(c����z��A5!�p�g��y��=y�����g��f��m��Ly��[yNt^Ez�pMh��H¯4���!8�2D���y��[���$(�����OTAE����A��s(\֢|ԕ?}V�PmxS�zD!�%#�ꑈS=��>DC��cmN���;BN8��2�rH�N��x=�y��� ������J�
8�Oh��͂�)M��/8P��I�zy#Tob6�9J�:;��S.8���ځiY��}Sxd13}��6x�[p���՞�fV�*��lN��
��hs��7{��:�<Ў:lf��2B`%R~�g���c�`S�uֻ�L�ߵ���BI��	K�a�_��_3�����p�
\EqJ��R��"����=���M��*Ĩ�oT��{��e�q�����zvu<��:�d�J1��wTfazQ{.%"�v���Kn�UK��ʏq�2����?|�n��
	ЯNd���;2�\F_�z092��u�e��/�p���F�=�|+�i�����h��,,ު5��xD�6�-~��j@ݬ!(�tɺ;������n=�Ry�( ϧ��:@��鏾���]E���8Ҫ�Y��|���}�D�ﾳv�p`��O��d�y۳f���][�E]L���='�.�F �"��������g�~T%K���xHv⛏o;�G�*HĒ����=�~���M��8�>7��,I!	�ힵ����55�w��]tչ�����#��@�^�^���"���	��V����F/3{��w�Y�M+H�MzY%'��8�zc3X��Q�\�<�(��&v���.k����͆��}���_��^L���N{�đg¾������l�~Xb�״'E��9
j��:{�Θy��-o ͆^W�E�%���X����t��\ǡ��_�ѥ���9���)]Hc�gq�K����{��%�]w�r<i�2LAý��x��rϽ��~̿�nƆ4Ԉ��L9�]w��H����=��q��(1�3�E�H[�2��$Ntǆ�o-��+� ��z�BI�?��$�}�|?i�;����G���_��y�)���ɮ	� 2g@�zz���V�Z�i�b�Ʋ�v�7j��z=ε����K�:>�,V���2�����Ľ}E�p��D��*�&ܨ�[��Ȯ�
��{3�kf��*��霔��)ط�/J1vE���{�	6sq��3�jHW�в���}�S��f��R3����}�x��k+1K�H��0-��۴�6��CTT��Q!��7 m��\��g�/�y��s�������CŐ$��������~�٥�">��U��G��oHn�}7��Q�tj ��m�M��25#��-͎:���J3����S�6ˌٔ�C��������,�`HO�IVk�U����BaT<,nK��"��ּuq.��e��P9�R���2·�:��r�u_X�k/w)�`��Ҹr�V�nX/wF#S�:��C֨6r��#�o��$�Oۻ��#�/����oo�<�UX#li`Y�ࢄ�}�N'��K���o��z`��z#��R��Dϼ�	�Kˮ	��d�b�W�` ���O�����bY��__��~�牿�9�lȪ+ ��@���������_��m���')�/��B�F����s���zp	�O���Ϫ�,��xw�9o�Ւ�0r;3ȅ��I�}f�}��zݩk�����r�Z�.q��a��LZPE�b��� i�2-:E�r`3�K�7_�A)�B�x��+����f�{�)����f�N���:�XY� ��/�o_��I�3YBPȚ6�x��أNᕉ��N����C�Ͼbn��J���Ko[R}���r��i�D���_~[J={=�O���m"�2������HEz�'l+'m�sgx�CKH_W��O3N}���հS��)J+"e�r�b���b%�b�e@�_u���Eu{x�N������*1�����n�ۭ^���jo���3��ĉ�dX��
�9�)a�<�heLv���p��}0��/����>��׮�MP��>s�|��@<��c{k�.��.g_�T�.U�<���ȳ���un����\E�G9�Y���I��ӿO:1��^ش�L����84b�TC�A��_�D��j���DU�^�]�h�փ&IwF���K8��b��~�kCWlzr%��U����+M3o�'bWOu�ӴA��8��Ԩ5,aF�5���vvH��F��7:zn��}=��s�+@���}w�B���r~��7$�=Fl-9{�N3@�]wv� �.<(��&SG��l܊v���C���>q���=�{�����p�*q���7���)��s��V���v������@��0�SNR�<�hls;۵�Ƈ,1�!q�π]�9]��F���g�gk�]� d�g2	��m��d��@*.E،���c��{����ӣ!�əG.Z\���+�"��TL�{��Ͻ�5�h� ��|oH��W�m���{.��f�3x�<.�d,��7��=Q�*q�.����7�����&��BPs*��JML3g<��pl���?�>�d����"2�"2'�<�����d�Q�}R�u/��ޗX�l�8l ��à���^�Y��3�UE2�w�]ey
��{V�4У|����g��J=�h��~k��7�W{�fv�k�֭�S���9�F3�r�����f�1w���D}�vܼɾ��~�7\���ˍ������k��k�UE苬�2'�ٱV�ڮ�5]�6β\�˫!�T �17F�]�ΠD ؅�g��\�'�͖xxvU��Y{�$�V�z���W��̛�ޟW�L�vg��q��G�&T������qyab������h���'�.�Bo�7�~Ϸ����s5�~}�����r��mE9�Yb@�g�gh����p��wjr/��h䮺��c�^�(��9#އѻ�ipr�)I���Ʉ��O�~�)\��)Rjj�b���Aw+�2I����I��Aw�y�C_)G*��ޡ�V	?km`�fQBB:��\/v ��7f���>U����[�O�T�W���j�E��� �P x݊�)��X�k�Y�S��ys�\�p���r,\x�`WE��[9�n\H��o-���_b�c�^�AQ�T��fP��`�Ὥ�tH|-H�ʳX6��8L��+e�^Qv�W=�Q9J�1��0��q՞0�nf/l��<be�]����q1�?c�Y8��ԉ�B*t�gK���{D`�(��@AF�3-i��E��Z�LL=�&�����[ۇ7��fx�:�̕�]9�C}ޠ�+YV�,:���b�GE��w�$=���{�-���q$���:�[)�^SZ�Oz��tʯ��]�ۡ�}Zsvub�F��y=�}�u�ˍgX4��@EM=��黛f&k~o{c�4y�d!�:��!ADб�S{���EV{l���m�qib��
Vr�Gr�D���S�4��,m%ך΍7��!��͆�7�桭��J�f��Ϸ��9]�r�ȧb���=��?`���9:4�.��0�\�wzJ*n;�*�`R�����F���Hy����Ѷ͵��N��g@N��kaY��e���:k�Ъ&CX��.�쥅�l��Ո�)_(��z:o@7D�u�O#q+�R��f���tw��G�%w1,���C����Ф�u�i�6�on<���7Ş� ̛�tb�f��1U�c[Ά߼*.���3h���.,ܴ�e��Cj*5ۃ\�Af��V��K{���Sb
�����q{�v���2�n���:��rN�TJ�)�Ҟ���ҼґS��JK�Ty�=�<\	ɹ�Pt�[�N�^`���a��-�)�[޼�n��i��U��#3�v_�U<vuX��r���0뭆O���;�jQ݄�p���"�Uv`{']���a0���W�+&[z���F��n,�	ZA�BWsd�ٵ�R1�A��#O����F;%=|�3���oz&�g���.:B��_CH�z��r�nL*5n��h-�w�˶*�+%	Kh��w�Lil��踯���*Wį��9!uD��P`�V��6XBK�k2M�C*v�m��ym4�2&ڧ�m�]JĀo
�n��/���xu`㽣9�=����u�D���m�]�9��wa��+võnN�Ru4��JnW��.�O�cwR�f�s\���\�]����IWm]㯔;�ض[J�����j��yFD�(��e�4R)�)$��N������Y���*Ϣ�=��Ա�&�)t�`WFˑI��.q�1�s�?lT/�j�w�R�g�%�WOML>pg�=3�t��2Y�&�Ʀ�Ou���U�eù>����7�-�p,w������P>w#��#ʊ흘M����6`���3�.A"���6ˆ'����:�]i�o�1#�<��0@��~�[���f_[���̭��bz˛�^�]��]eyC��W4��-�:�;阆\�)�I/H�S�@gs|�3��|O���I;��s��fkz�v�}�����8D�S4#P�Ǵ9���d�ā��k;����y�A��~߉���Đv��${���/T}�\DDGf�_s��O%�ԗep]��ra�]k��vz���ꦢu�=5��1I�%��"`�n��:�p�|
�I����]���ӿ�{殬<�zv��pj\�e���5|�*l�ftpRk�'��	'�Ģ�ET\�f�=��ta�YJ���+�]��p�Sp�$a�^ν�WK�r��f�µdb�3Ӆ��L��	G�u���n>��l����E�G5r��L��K�-ɷ��uM�IS�$���fwW��f�Ñ��}陘��v�Ί��Ӷ͊F!�Tr(���+�]����s�;)W�i;��y���!�����(qd�)��Vz	�T��Y��>����(���i�f�K],�t�t��6T��ª0�7n�;����Y���ɋ�%��Ձ!*a���">P�*=*�ϱ�4�P�	�9?����ϖ�}PjP�˘Lo�bY�<�CV�������0>]DM�dM�'�c�����i��vD�Mfǻ���¤��<t�D�Ɵ��7�^��O��[o��v���7|�9�R�y�d;�ͪ͙;Bc/���s�j���A�C����n�|\��u~�5B�0�J���4���:��;%�[�q��P#�m��&g���F�Z�,��=�$�S菂-���3��������3��~�{��w.�[~��W?n�<�	��u��Y��f�*J�D��! M�W�U�TFV+�i0�'4���E]r��`��f�a�����ٜF9Y�D�,9G�,J�QQ�9��Kn}"��["ǻ+���W�&��yh2�2�n+���F,!$}�m7��=W͙H����˘]L�=�V��˨�T�,���Edd�,���ߢ����Ps��U~}�cG�	�:��"Os�7li��O�0\���ݴV�e�-
Z����v��1��FI�����W+=7.�5�.=息�������q�/�BS�0�
�w"lFf>���vp�
�#N1���o����8G���u�5l�qi��-�b:{��3s٦�u5�/v���~�����p�s���v��5�g��DQ�(AB9����}��ו��7\:M�����b߶3��sC�	V<�F�Z�l�	���2˚�����wj{J�hč��2_8�Dx7����.l�3��UE9&���[�N���5�P�9�n�r�rr�sx�C�>��c~U�u���'�n2�������ߟ~Λ�����X��*�Ҳ�@`�d��R�dA�Ad$Q*��o�����,�Oz�;��c���]�ܿ�X=��>=(5�3V��Ʈ��t�{�5�d��)��g��F;e�ZTE��oMB��.���mC��%���]lU�hA���j`��gה|��֓�e�{H�B�\�C�X��L���)��7Z�.G9;0�g��}
ߠ����c��@��A"看jK���-˚��T}b�7��q�}C�7Ukv��h��W�����^  ��ڕ{�6ʝ���+�Pvrjz�<�ud�fhNjn`~�c�"��B,߹b�t���
�VD��Pݛ�����6���;�D�|ePk�I�y�]e�������y[<��s���%p�?��Zϣ��27#�&I�BU�*���+y���À��.�7S.&
�;���N�4:bxʚ�6�R�y��N��(}�m�L��߄̑~M���=Wm>��l6){{F�^�XG�{&��~����w��o=��'������ߏ	:t����50:�T�0˟�^�����9�}y����{�iD���F�iL˭3VI�Y TbH(�-�$�1���5��}~�F[�sX�z�P��V+U��&jH%�w9/�̽E�6"�c=�f&��_K�V���䣯vp$_f�~�ŢE�3]ߙ��������TP������5�-`��.� )��0+N�e�`��#Kޣ,���9x���is�K$�6��@��o�siuu1�N'5���m��{ia�M����s�}�J~�y\�!�>��9R�ԭ���e"��
�,`�r2{�&��8!?(���C�w����~�|�F@'��^ײ�R��4�o	��#��K�Mab�<o�����|�Ů ������x@*iI�{��@�9>�t�����ѧȨ��u½�5��Ϲ9'a�+y]�>iL��5���$�-�"���ܤ ���Յ�b�0�T�P(L� �G�=yBw�>�-���O3+=�	/+D7��/y���+9&�I��;x��O����Fj�)�E����v�݀\p����e�F�G2/M4�\����������y��[�sFf@�i�XA������ѭ�_Y��$���{�f��0�+as ����� UlTY�;�Kw����x�)h��
��&�����yv�-8�D�*j���e�Ɦ�^b�`B�-݂���K޼��94���3�����=]��s˭T6=L3�{�u	���������>s.�X�$Cu{3�sU���7��Vzi���A^�����1�� +��K������m.4�H��璖0���[q�O����=�q�3��ĭ�ۇ._���N+��{mާ`�4^4yq{��o|�+���s�{2�m�\��t�98^�KNc���,�g��F �ph�񽝐'��j�VͰ��PL/H��j">�=}�ސ�E�ϭz�C&�_R�����a��I�O�Lr2�H}{G�͒��0j]!3�"���~����WB����]D[� Tx"��Ϡ�(Z;rJ�w�᮵�������*�c��RG~�AX�5N]�b��5����O�y���{�l�Z6��@RJ��)>�W�����[ݝ�������:�mZ�4�d�9ٜx��̻��գ�U-�8�;�6Z��2�� va�2���g����n����14p=���FDR��h���t>^=�A=�iJYX=@����0�j���3!�����HV\�/}���O�!�{��z�ns�V���䮝MY�]U����<.D�:�|=��<��.B����#(���3�J�T��U�a1I��>��}�B6`*�x4��5�0S����f�a����C�<�m��Q��Xɜ�N�u·��c�2Λ�7%+���`��T#�:�����t��'a�Eku�W.� �W/S�[���º�Ot���l�v	>'�i�uپc+/�R�g�������cےsZن}������j1��7t���xd�l+8;�Đ{`$4(1[���TfJ�]����љ��DB��˹2X�vn}b<<�=,�|6�Hz���v�ہ�Ҕ�i�t��W$'P�x���i9�+���P�tX3N�f(�H	~�|G����g��K>r����((�Dkάْ��Ҁʾ�V�j��:!�c��x��G��W_i��OvU�4��K��yQ�/r�4�Q+�nT?���d<�ݯ�y�4�OP�}����V&ʶ��vt��y�w)WE=�̽7:�C���m��=3B·�4�uoJ�#�z�#���+�Y.�W"�q�u�� d&5K�y�v��!�5�Yf&�l��_�|JWx�ny�f]q!���OU��J8�OY��l60�Q���vQz�nDHpr���3��{�-����|�r�7.-�Fv�X��#+�am�ޛ�u�i�t�G۳�\�<<�o�Y��kNk`��㸇~�� d���'f���T���<,])��ȧO];�?!z������V�H
/(�^�[^�W1��C���:i��1^�8�Ԛ��q���i�b�v�k`�^��!�62/Ԙ˽G��XZ�1�oX�klT7�g'����(��BҎ޳W���(fh<����9x���³�����`�bDT`�Pa �c�a�d �VB��T�(# �`b1@PdFA	#�"�;���{�1�s{Ç9�y����yzV�<&`�q���W|�+ڝ_f���pR��}�;�Hw<�RJ�V�옃=�u`�l�r�(x�g*1?[P~N���J�4��"z%h&��~��e�o������/�g�o���6�vK�>��U�b �0�
���e	��(�V\l���WqS}�X�]�������?-7�}����ʛ�D)��n{�Y^�9Z��.�1�u ͼw3Q�*�ot�H�E3sM^����ڹ&hv!8޶�Qw�&�pVzA�����z�[�'GV�ks� �}�`P�ʇa�`Z��@=H������2��{Î���R��U��ʉtH�?x6��l�����}}����u9{�	��ts��s��jf���X��JJ�9z��y^+��ixڮF2U��Σ�nj�⨙"�W�-�;^������_���J	rC�����os�Y�r���3��6�{=b�ۯ��D;+h�5]�>8��(Ӷ���k*���j�V�4SW)��U����nH�l�E�!�w-ZO�#�QqN���e��y�bo�)s��q����Hh%m�.�ie<
)Uw�{t�4��;�.]�	�Y���rx���I{OsOH��[���]?�����tG����ΎJ��m�J�B�.F�CtE`c�k�r,��Mf�7l�e�_@َ��t+�2��G��{�:��j96�=�p'�Sq��ɱ�>4�!�n�T߶�-C�ؿ^����C��i�	~F�o���c�U�������1�'C�i�WW�\���2�^��j�xnT���9�2p�7�nk��9�^���WBq��Id+l�C]�������ä?B���?VS��x{�N�լ[WQ+@��1�ؗYP�39B��~��:6������a�	'����7'x���g���y��{�r�߾��?BE$���5z�1�:��}�z^�%��=}�믖H�1gK�#Vw{��M�����{���Y�Y!'��5�|��泞R&�_I����~΃o��8���3Z�2�1H������a���??M�
�0NPiuv%���$N�������I z=֎�gyuN&b�nw���;��e&�h���6�}1M�Q�g�+[�ں���(dB:��u�PB/v�r�"����y�M���&�l��ɐ�� N�R�h�6��U¬wowe����{�<�J�9�e��+6�2�������:�B�F���rڐ�{�Y�����%�WIܷ��.������g�S9"jsy��S`,�2�-2�H��=w�S]y0b�h�B���2�@�|I6�b�Z)Y�A�#͙�sN��`��ܸ)��J[YK	YQq�5�a��!���S��Bbxi�l]R���"7'n�m�����Kx�5tSt�{ҙg\T��u91g�A	��`��ه�f���h��Pl�T��؟fˠX�w���D�BQ2�m�2j�w���U�6V�k 4��F�R�4jۄt&��x*wr|��1@��FF&��ȢIܫ�	2BF@�k*��)����1%�)Wl �Q�_ �'Q����$E���@/�r%�(22��m91��,J�i����������)ܷ)�v��v����N�;u��0��ɷ�۝�����=C �Hm[�q+_Ʒt�<F�z�iMp����v_g!
�S����[rs�o�2�W֟0w-��lԫ͜��{���o-4y�=�=@w�1�Ka�`�7^9��R��Qy�J9Ob�1��3Q.��Y��X��k���F����֣]�b�]�{=�����=yo��H:�:�\�7R���Vi䎱���KZ�`R�s�!xՓ��ɔgЭ�+���\+��-��F2��+`2�U��¸(`��y�-c:MVV��.�Ά�ו�i��V�Q�5�[���H�e;JM��g|��fP,�ms�!�SGmut�IP=B�H���V)\�5z0.����m,#,�]���34A��Ӝ�45�q��<���Ӂݩ��p���[�t����S�W��ծ�w3$���2+���F�+��&_tɍ�L����E�\/!a��wڥ���J�(Ha�e�o�QU�� f������E������j<��4Ag:�F=����T�p��Aک:ɣ�W��Bf٘`�X��)I�7��BSV.���w˓���G���a�M�'�k�o3�BM&|6���]mc�A�1|�5ܻ3v]e�y����M��@�}�уP�FZ*z:��C9C�qZ�u�l�˂�]�:��r�BT/5�8RpR�;{J�-仅3h1����q�cf�c鷗a�f���4�BY����1{:�+)!����-Q1슪I$�I$�I$�I$�I$�I$2�oWY�uI�u�L\�6� Sud��5�-��g��F��gd��Bs�o/(Qr��O�5�l���d,"�n�e�p3�<s��'߼��`?^#�]��,߰z�6#��#V���� �k�p.�U^�>�p�U��N��7!���نɊ�����v~S��1Y��z��W�t���1�T8c�����_�}N�]j�|C0<Z�!`'|�v�NQ���i�aKcfx*8䚇t�f3��{yd����5N��t&�z-�.MzT�6�D�6>�
�fg��M"���8����f�4���E�����]�ǌ��j�=�5�lv[�b�ȍw�wU =�tO���}��y����!����ξ���� ��!����Wn��Y@��%��!�]�^�ǢF��$������>��l��~��OkG8�D�#�OԄ�[���P�+k�4ҙ��	���o)n����/��ќ�x����e��
z��휊e��}��r^a�A�cצ���R���i�Ƭ-���
����|3??C�Z��	w	�Q,�7��hB�������AF���Y]ۍt䤮�c$w��mŝ]�M"�-r*F[�voN�%�H�su=G)`��ZZ�h.FL7s<M�14��ɢ�cH�ɜ5'1�4��4F��<Kw ��6{f=�$�T�z�Gj�d���{��[_]��,`�s97�C8�g�i��\��HW9զ�<�$)��/ښ�dڣ&��D@����e��IQ�h_�A|rT�'@� 	{��tp��s�N8w��}�-/z�K9Kc��2��l27�;��?}�j����~����E GϻϞ'�/3���_�ǔ����Cɳ��C_jk��Q�&�����f��%�[��F
cb��g��}��~�(}��ӛ�Q�3���&�������yݰ[Oc�j,�6~������1<yrM��R�چ�zy�:'����g�ŵ=����=`
vaO�$�j���	>~��ι]��o͙M���z?Bް��9�2��s�d3+��!�l�wM���V�D��.�E �~����Y���(�+�}Eq�&��ǥt��_q{e��:Sը�Z��gk�j]u�1}n��oܻ:�Mb��b�˅���8c���6C�Wb-F\q�RY&p2�1���GG�]	O�X;w�n�w�J�j�4k��I3��������E2�_�x+�nv�K�kf�h症��׿���?D�46���i�[Ő��&�GtkA�P�>t.BC�
���\���GJ��\�6�̺̽�w�5O=�����I���S�k^�z-��q�}Օ�r����
��d�ۏF�
������Ҩ�s]��1�V�ɓ�]�ó�[���x�ܱ�G�>�.#菘����nUar�������GN7�i&��i�7f�l�Ƃ�Yr����be7��C�����Ґ�G��e��}E*؉G�x+�t
A�Cm�K6mhBP�BQA��:C��cҶ�ҟ;#�,�D6t8��z�8�޳�7(z��Ν3w����|=y�i�Κ���<�5�غq�.ee�����@��?33(a��`�+��+1���E-Ii\�p���9A1&&1W,P�)H��V�e(ʔ��y�������xV[���௪F3b<.��aEL^r���j�v���p�\ȣ��J�k�Ie��I�Ӣ����k8��$�畉C�Ո�t��_��]�vްG^�^�{k*5��
�v�4\���3:��6q\ H�v''}�mr�x��yϏ�x2��S�D�"OX�ykÅ�Bj�פ|�K��`z~��VJU�$a]pO��,{���F�VpZ3o�;�=���;�*ZiTN#��61^[��g<�/d@z���MnV�e�(�7�JI�:[+���4��Q�� ߀�j ���fAx�߅���(Ϻ�f��sc�0���DV��x[7�)�L�l�h�0���}��`*e��sE�j�aT���Y����׶����AnM�P��C6U�������iw�1Z�=��H�����͏�X������=��� w�{���>�z�DG�*�4o��ݻ� ��,a5�~��f�]���#K��p�ze����u&^Gf)�$��5���|�z3�����t�0�̩��E$*�Y@�-~�ܬ�QmƵX5`~K�v�E��O�l��dIR�Ἑ���7��C �1�]`w]����;v��ڭ�����ē�J�ȐJa��bg�y���SX#E1��ˇX��A y�7�2�b��c��RaČ�����~�G&<w�[o�ꩧ�a�c3%�r��n%��K����.Ǯ�c�^%�G
��:�f��w�F��ށ� Ϗ��r���ّ��(��|k��1�	��^gv?�5CЭ&��]�<�����ߔu�,4~'yUVG�����o��Ǜ���dB�YG]}�G�������0W)�SL(�`LiR�w~px:���5/t���p����s����j�2
��?YOє҆�ls���8=p����A�Ŕ�H�|5�i�b��1^/G��m�7Ao+�R��k��L- ǻ�	�z�-�����k�!f \�}�^z��{�WtOw����1�]1jʒ�C�ͽF�-��>�[��߀����{w�����fQWwf|I��*�p��\��]]mJ���4j��U�| �(5�簱z���K1`�`g�%ec�s;�.�̮G�u`���yj2�s�&Y]M>���Z�����\s��~#`
'���>�1�A�?��R�\w��x1�/��)����1>�9���O{ƹ�5��/��gKۢG���ϴ��K��s�]t|w�3��HB1�y��W���"j@�4Ğ��gV,����s70�[ߕ02��U�����1���zй|S��*g���ǧ`<h����ñ�p�_=�68�CRֿh�阼6�#�=�p{�Vt-��峄��D:v<�s��"n��pA@�A3� k���yiw
�c4n�g���^�{�8��r�V��� ��C��z��De�cס�q�FM��83B���W,��C�\|������r��	��k�y�N��6�r���*{�m#
�:��J�z��]ג�>QW=_��ۀ���X�n�6�id�`��9�
edy�/5�y��w��uoO#8��3e�L��o�n���dj�RD � 	"��-�1�40����}�0�d��)a�zу���g����W���x���ړ`:;LX6�c��pv+'4训' �h��&Qس�}o�8s.#�v2=FQނ2���_�6��g6	؃�+���7r2�xz��s2�!A�&�v����zp�)ݞ�4�mdc��I���=����o+�_\�zFJ���)秧1�&=�.�zu���y�z̻�-�\�8��  2��v�#PX�,�ځ� =�:�,���Q'����X���pC_�M��@�b�w6:e}�_f�|�6ψ}�����HC���:*�m�x��</�C3���60��d���4�[Iȗ؊�/Z1[u�K-���y�L���踔#�E�G�����}w~,�D��N��}B�����˜b�ok��V��'��UĆ�G
��Ɂ����J��3ֈl{$�\�I�U�yܹƆ~�$G�r���]x�s~�~����Dz��S�]0�U2\uw��o�@ސ��]4�j���%&D"=�s���_}��=�2K�!G�2�[RH�2\H4rVdf	q�P�B�,�
�dJ�(���i��"�W�볳��"�x�ξ]����9K��J��� _�8'.^�#�s]mp7�ɕG���YڹᲰ-�n	c/��"j;�I�f�Gd��Y�?G�"~����sI���3����E��7����Q3}{�r��8	�n����/�������v�bچpC�� <'��MgV�˚m��3ʭ3n'V{}V�#o����Ո/W\�:�qP�b�i(}��	.�#h\7f���@AuS��~�w��㵖p�S����5ށ�{�.8��;Ȟ�ω(j�R;kۡR��Tv��>Եì��K�`�a��zϜL��F��=���Ϻ&�J,�uU���5'�T���H�c���k&�6��G^!�'��u�j�[į�|h@>��
#ޞ��*(���c}#���s�V��ʻ�2b��q�M>>����۱z,z�+&��Z��ǌ:�@���TJ�2�8~�4	b�f�i��{�m�":jq���#�O���dp(�#��
��U�	?M���JrH�0޵���ї%FV�)KK(QDZ+�D�
���UxIwa\��L}ZYg �iy�5N���e�������R"�Op�M�A5�N�<r�j͋{bSB̼�aꃬ�LK3"�]�5;��g�w5���3֫���dz�����Q��CP_�K���\ x<�;�~� )5���Դө<�j[�B:htb�X̋�]�8�d)Q1�x�Fx�����KS��:*'Y5&�
��;d�u���)��`��X�3߯���{����?D�����]uYy�6)#s��(�_]=�J�i�/��������� �Z�lb�,�^�}�݉�`%	��~�s�4#��^s����Zi��
��x}�����ti�1��ԤrMs	�� {ޖs�7]�������� �)�a���O�\�<w�Ұe{�:u�7��wk+��r�SG6����)��Nh��Z�c_#h_)��Mwx1�=C�*�4Mxŵ�qL�n�w�̛Mҷ2Eպt�H�.~w�&
1��o���y/��K��,����tӊjC�l��I �~����}�6lP7���v	�=qK�!Y�Y�-fC7�3����6���==I�70�s��{xxeCf#w����K盅����z8+Ss��R`Nٵ�{4i�3�a�`ސ^�V���2���E,�8�;L�牑rě��9ŷP�ʌ<"Ɔ�Y�x�[§XLEs=."��}e`��6�~�/8v|L���� r����!�x����V:23Ț|����~w9� �,�g����j2e��2_H�h[w��xf�R7�0�>�ig.�ݬ��a��:#�y�[
�ȭj�b��t��=e�(���X3r�zp��J��&c����#;�h�^��Ը]��Xn�S�9A�qٛy/�[�qyv	«�53!i�sQl﨟�麇ǧ�2Q������)���[��c����#�m�{�]p�
?�yh7�����s>���C��.���~o�m1K��1���y�����1��w�s>ޏ�	��g��i�mΤ��L�_uN�i�o��g1Zӡ�*&��)��f��r>�X������+�	��<b�\��RA���9�6Pz8�7:A[�E�����H�57��uad,p
�s���϶i���$Z�vs5��f�ӘC�9��1��<vT0��	��@]���wh
�n;��И���_�__VU�B���f��9�99j^m�N�E��e�S�SwN��l]�9���7��[z���̧�e�o]{�g��է��
���s3Bq�/S�����ͽ�:���5����m9�a�%�r���L*Ƥ(�J[h�v��)�ҧ����l���}M����`�C2񊎊�;��]n�b$�B��wF�E��m��f�Z�`�Vk�7����T�9�uq҂[-��$�~) �Le�K3ec��+�&(Ͷy����}�&Q- UPwc'yO��Q:�-�P��Ӗɝ]:֭�L_0���;m��Z$��YAQ�Ⱥ��&��w�Mo6�d�1abWyqw�����5�Y�)�ٕ�D5}E�-IDQV?|5��Ȓj�'��<*Qx^jۓ-�f�"��Z{�d�{��	M`���4�qн�����h�ar��1^ �]�0$�!vz�;ם9�q���ws[��R�9�5�y�'�QI�V���M%��v�x�Ωu�r���I��՘;���)%\�1_>+Y��\��S�rvP�r��\�緰k���"�a�aۓ�;���絽��k�ڤB��·b��i�)d��w�]�W�]x�2�<�1�O΢���ː���V�ͮ�u�RR�d\�(��a<@s1��'Y�1r�&PW+D���ˊ�p+j���ϯ��!��:5O��n�F-�|zݷ�1#��/F��	������D��m�֕7J��K��i�⯀R�:�pvc�xقޑxnL��]*3����Hv��&�K���9#J��9�Z ����y7]d_v��f@VixU�J�=+]����Zw��Bq�{�l�I�Nj�F�;��N�m�j����K���5��)�KPZ&gZƷV�V^���2e�RtsNO
��o�62G�;2��5+
Q�j�����x�3jT����^��M��-��Lʻ�B[��:��/�ǌ��B:���ž1eh�hǬk=S+�Wu5�w:��,�p�4�$p�˸�DU�Ne��0�ok36�u����;�֫ȸ
�n�mwc��`�H7�P]]/���w�R���˻)1>nQ��;/ ���՝ٜs����OD�u�QͼG��Ń'E:�7��I�W���KT��]%�\��sV͗��+�]�2�<݂�����{4U���U�2��8�)�ζƙ]C۽�����v���-.[�����C��8mΣ�WsJ�Xѧ�-��o��`M:)���ۻ��]f^b���b����!�_��Q�
��G@�HƑs>�@^o���y�٘�QP	hp���2�B�%L7IښU����bfߤ�!.�f��c[�"���ɍ	Р/7�|t%�݋�z�5?�O&<b������l�w���������;�s�ea�i}z�}�������z�0�W�Z=�{Ó�G#�Ë���8�K�}Cb����!ߧA{���X!����ۢ�BU7����J�$O&zz�d�٤��&�J8z��8�eCE�����p��\kѨ�LA뷎���֩�8l��M0�x֣O�\�7��Sԭ,�lp9�,٤#'�� �@źi�׃��5փ�,~2f�=��,K�:��V`�r�t䐩;��ضr���yިQQ�<�s�-��S��`��DE2	jX_!���	N�GK�v��9�a�>���_}kB�ʈhS1�0��~$�A���,�]��9�$��ֿ��-���x=�]���p��Nш#�dےJ�AMS�9�_*U��;�FiL!Z�j�h�u$��@�f��~��4�L_0g#�5���_��8s��ggG~���n��0dl�Du*��XBb�{(�������?�P�-U����{�x�.�W4r����c6@�}yėy��	��n<;ᷛ�<y��?,U�2�Q���k1�q�zuW��s�?�U��^3�3r�M�N)��N�S�r�XǍ��@w�Хa�c�{�1�|@x�z��0�3�WZ��=���ϟ7&FBs91oNȼ�����djfeS�x�����M}��ٍ�գ�:]��i�˹	7�����a�g�6_3YG�sb���r.mVr4�>�l �N:ś��EJ�mk�ك1�"��r.��K>��:o;��_{�\�I}�����o�2��1��.Vu+7Z��jx�j9�H�y�X�q��p���A�k�O+�Tp�7DT�p}k�e�,Y"��Eh��@d�S�����+[E�T�afιu��e�KJ,��й���Kk���[�YLk�5,Wu�U�����X9Hٕ��+\��o+�o���pNc5[�uv�\rq�K���\���u�2����&8�%F�i�3�:���5[Ja�s��g�����-��[b��v�Tn%�Bc����
�#�<�b	�`�^�-dG{��|^M�/��(�ir^\B�DG:W��͟t��D��@>w%���W�r]7NR�Eӏz�G�������ke�([���]�kJ�&�����0�W	�b�Y'e�^~AY'��W�j��
��{)>������]�̓5������(~s��u�cYt�?!7�������wx4 �8"��7���m���q��:1��k911�A���z�*f�753�Y����+a�Ơ��m��'0t���QFm;F�a�����/�rBN3�>s#^� EL����슘���)������=��}~�A {��n�{��Zf�@�ƾ��c�z\�Z�St�y��o*��`�sT�O� �~���PȒT�ċ7�����۩HL�y�oh�Q�+F��aB�KEG���鐅�1�ܱ�M�Lʤ�Ǉwg
}�����zYXl��7Iu���cO8�:n��a�O���	�y������!9g;��� �k��d�F�A�okNB�"�=S)����(���{�
���0n߶�nf7~�B��Z�����������Yچ�����O�&Gs_�7�A"^E����
�a�|Gß�U�q�:�+�����u{ϻ�����?2��#��r��������L�y�&Na�~�3����x0�^����G����z��!����J��k�A�Vg{�?�;]~�zb"�'�K-}1S*V�iᴌH�X�:kJ���U	�X�-�݈�7�lK���|ӯk��a˛�lG	���~ }��R�B�W��Dչ��g3�ת�9����ɞ��|��u��g�D���^���*���=lA�3�yu��<��?�i��I"N�����L.�[���̏
��깽���[�D�YJae�"ė�����5���̾9�2.�ruh�(J����Rf\�?�0ԛ�t�f�������]������=����ۮ���:�b�3���:���G�5�$ۭ��g��������C�"�����Į�9*����G�O��q}b:��u���g�ٕ��V��md_���3f�u�6=n�Ec�aK�Tj6�Ia��J�=�o���E�|�����=��/�bC򭂳��T
��M�����ݍ�w2ϫ%W"����~_����H�|�����y�������DF��{�{-Ϣ�`H�y_��-�-���y˯��<�̓F����}33!��}�:��/���ݞ��?�����u� �c��$��J��1�4zi}��}�	����99Kbl2�C���Z��W~���+y��̓M���Y q��
�)�zV���E� ����/������!6����p�Cq}|�oS[�UnC�2$mlc{��o��W"�>={�k�
�u�B��`Di ��6�[1�b�*DED+(���m��Q���T-/�4+k����Q6��г8�d8��ս���W'*�n�<��.C�b��nA��Ft<��υLuKv��c�<-�$�eЦ
��e�MI$�A0n�fR�\���;u�&헧v�FV�ҝu���G\�����֟?��F�EB�xg=��#�J]�٬��SeIʥ�}Ne���I<�V���>�l��~��sK��s��+	���P!��E������4ud��.7�2��!��S�!�*�:?1�m3#�p}ο}�;瞨~��B����Ic��uZ���	�28�A�cN�
U�"YP#�'ګs�C�[HT>�O��=��^���@9�+����<��#��b6�ʠ4r�Ύ1��D�F�S�:�1�.����O��\sϲ_��  �������/���G� �	�|�f���n���|�긌�"댱�ή�L��o)���fsӹ$�a�4.�����µj�_�V:�i�K��>�:_�tT�0�$�X�,o/���V��d�U�5�8�34�k����<*�� ���~�
[ HbI"(�2��ϵs[_��C����3̫��A+�ʸ���8���]u�oGdˬp�In����������n�]����v�-��cG��C�n�_Vĭ�F;��3��N�c�:���f���)}��{�E	��lg�Vz��=3�ࣛ3�[6�D����uj�N�>��ձC�	�:1�yZ'�����чk�ڑ@;&��E�0��&�KW�Dq|+�Xɷ��G��0�H��NZ�mj�m��f�f�|5�xğ�R�Us(F�;s9�v�Q����	���B��Y��~��xnO�|Po6�)��ʞ��]b�b.�e���>��=AEƷ%e���w�ۍ�%�"Ы�fP�솦�*s������~v��������â�?]�#iH�V��_���BE��.��͑ϩve��\��Y�.�`;j��f�����&8D�ЀGSN˭����>��7�|�h�ha�d13�������|;pſvb�q0�YoK���ǻ]�����}���� e�68y1�a�DG��5e	���K�`���(!RKj҅�	c��a̕F1�R�	dL ĀZLI�$��r���&];���m��^#e�T|ں������O�7(�<�o;l�=b����o�ܬ�([��g2����y���gn�v{$y��/Ή/4�D�[���8�
��_��쯔�ζQ+'{�oIXW��ۉ�s1�qz�-BX||H���]�P�L.0���������gU0�\�;5ց�)�aP�&r\�G+(��u'��Z���۪�p2e�P����y�|;�Ƿ��ݴҎ���*��q6�eF d�����{��+�BT�J�C�,)��ܸ�͸.w�?6z#�0�!݄�;�u����?{���^x��t�b��޿�L�h;�*�.�J���Ή�e>Ѵ}Co�6�l/q.޿'P!��"K{� ����y��C���W�}��R���1}4*鳮A�]KRf9�Hj�i+����yV4#ʯ�P]�J�s+|�,ؚ)����g��:cYt�#�<.˶=��s��r�כ���+d�� ci��2��ƈ���xҡ�+|n�>ҠC0�vbP�ڀ���QH�i.��u�ti�"�U���P"¡�9���{��s^�<�z��]̪�5��%wW ��.���Hw3�N��%��y=�p|.�0[�2�8��N)#]�i�g�Vy]ea͒�Bq�"*�I��A�� �Z�$O����7�S����z�v�y�l�aqV3��'��"�n��{�/�xL�q���
Y���B;9���y]0f�e��.J�����Ǵe��&)T;9=C(F�h��&�z0�`�]Y2S�9�}��x�#�[�v�g���]�}��e�K�=�`�u��].���-*�"˖1�m���E���taT��z�Q��PwZ�Fpl,!G(����}No�!0�w���v-=`Td׊�u>��/FS<�'���1��)l�ᑓد��l�d:�^�!
8��*�;��b(�>��[y��x��pae��h���Ab�lI�����UF{{LޟYPc[C>�B�S&�no���ڳ�󩿑���9A��ț�A4�Kw@J%��j��ػ�2���`���SY��J�rY�챦�h=��6R���Jw\ƾ��-Ƴq��q��Ưi�8���V�b�]�u�&0�,���5t��.I&�2���I�)s*�e��Bm����(d�ROT}P�}o7	$�����b����x���<u�����<�t���NFL5�K��y�A]��W7��U2�i�]r�a N��s��:����צz�y����1�fп&��t�D��?nT��R�犭�EMruTa:į��L���癷������)P�x+����p|��(����.��z�y�牛�Q�l�c���[K����n	��z9v=����ơ�*�\\�V�X_{��H�S"����#�28E�ܨ))9q�LMK�J�Cs#���}��I�����p�-h��7���!x���3�4;��h�-�B+���SK\�_���0n�J����G5�V��5�.���Dd�Dc���@/I��ާ\Xqv{�6VS��S�,[]0��MM����G2�y��:�����w�jٽ`�'�>�{]�Z�O;%�'V���AV
�:K���gwf�9F�?u�&��F��˳K�it�����"!M�i�3v�ね$��a���ќ���ט��$Qh�(���ˍ��Ս
�Qp��8�\)����J�t$����Y�����El���F�|��8:˃�<���������F'��,���1�M5t`3�z��Ufo(�\�[��,5�o�d(\���}�����.�����_e��DB�	1D�[r�7�i�"ZQE[�%J
�Bc���!R�Pj�F�O��j�I��͒ݫ�H �ߺL]\�b�$�8�ٽW7��0H���� �G g-�BՕ"&���	�j��|,�)��@g���%nBˮ�wx��w9��1i�t��Z�0��a��h�	^R�(2�F��,��e����44��q!�
)�Y��E�0�P�L˜w���$�f�ո�5�f�YmH�n7"*,�kܝ��4�<ޡq)YR�̏��\�z�v���(�匰�v2�wN�H�-�w��}�ǋG^�����"��ϱTΏ�H�fݢ�c�\��7y���j����z$�/$��<#o�-�;��FNU`�)��c0�F������ܙ�we�b���h��q����Q�E���=���M�#�
!�w�T�##.�dF�Sq:�&h}7�dM�7t�-��@vV	�r��A��S��S{٨2fw^eZ��F�
�:LC�F��v1��/2d�D�e�#�<3E֬sR��]n�3���KJ�n�yi����m��p��QQXG�\�fʻ������4K��#s��y@��tDeKW7w��H2.�@��j�aR������o�΁�u��g$eR��[챛�3N0�SY	p�����P�@VN�8�)l7iԈ�G�]��X`�'��)^�& [�B���"�+�s������n3B��:��?U(�-텽۽p���cX����n�ս� s�&6�`���]��r��rn\�,m(�e��@��1fP�&�u	|�fQu�&c�Ģ���3�;<�}�����L��˧�*v� ]Z8�"�\���ȉ�W�Gw�𧒂�{X���:����d:�����ޕ�]�͓;��Y1�]}�WF��xՊ��d��E�t�!Ҁ�(
T`?M��qe�.�S��:+\zqV��E�P�V�{Je��U�[�5H�fL���b&�๏HM��tf�eA��[Y{s4��,�z��q��SyWz���$�I$�I$�I$�I$�I���i��C&X��r�����*ݬq˂�@Eg����:J_#e�S.��b"�L�4u�V˜
{��ʥ��r��gz�I�/�� ��yx_�������3���y��m<�"~�7[]-Y��zr{��abO�uk��茟��z#S�9���9k�̇��*������L��
�v���=J�n��9��,qrC17/RU-Зr���Cx[i����G����`��k(�&b��X�]=���&ʉ�Xrz$�1�!j�-�y��Y��1g�������&��_]��}�}N���\e������Π���R�u���Y+6�'t����fu�~*�^b�q��1���?K�y���z��u�>�_�=�rI�s�?/sw0o�=S�xR���RI��Z �j��m�Q�N�A)�Oi���u��tq��¤pj
�,G����R�^��V��3���2{��`U��p�@*���[�h������9ףCSZ�:��^l��__3t���}ϳ�2�F��P��)��ݑ6)�,����Ά�ŭ���:��i�U	L�����q,k7�f�v�=;ʵ��^�1�Yƶ�n����ں)k�|��/̌S�����~�#�h�7��3k�9�Y-���ү:�S��t�-�z�O��f' W��Qd}>��BT�r\	��]唠&��z������ %��V�v�'�պ�OˋK]��1�W"���TR]&���^��`�=��g4��S^�4���5���~2�`g�~����s�����}��6��WK?&Rʪσ�3�G���j���
d�M�{u5�J��2�0������ا�e�#s��?-������� �vZx�t9f�xrlRV�^�}�a����9TD<��f��V���k����S\ͦwܕu!4J&�������;Þ�����9��}����}�8�w~�n��|��Z��ĩ��qJc������kg��}��__=��}�� ��u�D�rKL=:3�v�W@?~�����Tf�o21}����!�d�fC!�BH#�-jVaF���°B�T��"ȶ�
(1�hH�
EP$A�*PU�l�Y��VK�R $���c �D��DHT�o�׻�(�� ꭧ����V�kސ��$N��ڌ<�z&_]]�U��	���u��A���>���h33�zx��do%��ɮ�+4� ÌՑ2M��lZ�֫��+��Fmd�*�nˎ#]U�i�:k]r�J�,ON�#hUՃb#<Kr[�ոN͵�Ԟ�d�z��!�9po�\}�S�Hnl �����7{�o���{�w�r��AT�Y����|]��nyİ��&��8KI��E݋x�vJ�XAAC���?|�������#��Ȍ��2������Td����.D&Z��U����x�Wz�Ͻ@�����m��n�_N�D�r\�'d+
mfϾ��zش�Wr�DËe����n>���v���%I���j$J���W������WP7��q���æ&Dnq�⏱(!	�_߼׍���6�~�浧��0)@��J�9����5_\�����u.�<��؎�8��u�DN�3������X)�Z�$P�K浞o����2X�˞��'#����u�q*	g>9�������[k�ð�@�\S8g*�P�n����<30����|�*+%^�ԒH��{����}�������1v���ī������3�ǯ�WV:�6�3#\�\8�P�GwޤL����U�iZw��h S6�i����3�d��� 2%#�x��(�.�u.����<
�#}}[�;�2b�I�O.m�E{o+����{��OxM�L��s���@���=��pL]�hs�+����eՋ����y^��#�o�չ1����>dc��b����p퉚�~������Wx׼rJ��T1���Q�dU����W{ϕ�e*?2%����
s�WL�?6"ge��Uʵ݅+�@���N��^l��se6&�	����R�^�)߹e��hgVhsCR��"gBS���3�h��}����`T�ɸ9;)]�*�4��#n(�qB�E{��/�ؿ�T��1l��-Q�� ��
&b5DqU���
e�|}�y��{s�s)t���Л�|��L�W�(�F��i���+WUヷo`�U٧I�S�AoWl�2P��� W#�LR��t_e���m U�`�!�]=���,��?�I$�o�۔�~����!�]��w�wT��l�@�ס�ZC�<��d��T"�R���}��>�t��,5����f�bփ�ڥp��{��֨¶���Z:D�rN7r�um���s@6P�؉C���_+3w=�\HV~�n��4U�L�C�y��1V����*���ul�Q��B�Θ�rV���¤����1]�d�r|����d����A� E��wu�Z���g��x�>m�g�=y�nv�X�q��];�a9y~9Ũ�t���S��g���sS�v�/�{ǿ�����ܼ��e[��Zê��	[`���e���.�v��9��xe��"����u`#o�h�;TY�T��(�h�����yL�`~���_8���U:���ߚ�3V�]�(�"H�X�Je����:�bo��+�ܹ�rһwT5ݠ����t�}����N��m�=Q�crN�8>�x���͹ػQ���z�H��3��Z�p�ߟ�)#(hv*iNۀOb����f�L�E�qqc�s/��*�Ũ��l:;�쓁��x�LkG��!��m��y[�����?z�+�hV<m]@r�x}�v4rR�'�3aL�D+y�c�-,7�V�����)��_��:���V����[g��u�"�1�L��sza.rV�Ыg�ݻ��g|8A����|�տ��xF��b C{�/}��
��LX�t�Mh�-�Ó;�0p�*-Y��}�E^^�Rka/ ��Z[��K����*�+�9v4=�c�YaSS����p�z5=>��2퇉�ז��R��|"��#7|f����gpJ�f��yt���[�m�<�.9�$>�_��������N{�������f�bs[ǳ�WM�J�M��l���F�#����{�B�����]}�٣ �kh҉l�A`�(���������_��w˵Q�S���u��5V�����r#��)����7JsR���|����<r��S��@��%��k�s�^ֻ�cg:���[��g�t�kM��s��Z�0]�H�Y;������(��5�]��g]��f/D�8t�r������R��=uVɈO�U�f�,��o�7era�ך�dT��v����:Q2��-x�!#5W|d!�g_z{�� X,�|��+ԩ�������\�\�ᇫ�踟���q{y̒>����LZ�NLT��3n���6��Zn���+]��h��W���~�5��ƼGD�+�3�*���O��gP���_RU��f��<�{燰� B����"���]\����<�X�)E�Jt�ȹ�X��`��P�S��"&�����N��o����?mz��)�#'�N6}�:��՝A��x�s�N(�}���ßhp瞜y��	$�w�^���.hQ��*�C���i���׊��WiR�w����<�h!Rq���sQֳX+�P�,H,�)�*�Z�im���"E�$QMP�f��y���g��o�,O���ɀ;����U���� ��W�4��w=����yem�R%F)`q�g�����=�9v��^@ܻW����I�5����C�+���W�<�vא�%v�/"p�#9{���i���G�{����ݭ������]T7�}�f��w�0/1Z�����Pk�q��ln���ZS|{���-��Z�^"A����*k���A��L�[;,��������Ҷ�8͕V�3dĳ�"#�8/�v��S�붔����Ǻ��9����и7>���sPR���qJ�+7[�t�	���X���Z(��f#�d���Ky��o��4�ww-����O~�;䧸8N)cҎn�y�EJ�b�x��A0۳0�<�zyR�m�X�����g�-N���pͣ��n��:=;�qr��{O��B�o��r��/3h�F�̉�[p$���VDC��~�G��馭她�so$b��"#&�y�s/y�㔻��N��O��t�:��L���ж���jM�|��8(7�(�;��Z1�����'���ql�`4�5�\r�ȭ�⣦u�Zr|�F0{�{~������}\� 9�}�=u���s��o܈���d�7,�1LFG$���_��6��P�g�ݍ��~u�=ӇI޽��L��{�˻Z'��4���U]�a�rg�6���j���s���Ab�{��c��:��9���������ܝ͇���PkFȆ��m*��;ڧ��߯����4������
�<��㽖
7�շ��������a����z���l��,�!��WF4l+�\�ƹ�y�V.�gH���Ypyu҂�̧��P��CKT�aq��v����TJ�-gs\�1�,�3"��ղ.1�[�.����+��ȁ�Dʥ��{Y�/�����v�))vn���ƕk��I:%�'�9����3i�*�c���[t-�F���=�}HPȯ(���em)���s<�{�F�_T�M]������]�o����hJ���@L[(���(��DM�4.��I`��Q�%;�P�\�G9�nL�cS���$1�-�X� {�n���u&����o|�8�`o����{��mu�HwdD�W'��8��p����DA���d`wf��׆nvߗQ)z�i�݅�(�6��NJ����N��ͺ9tJ�b�s�9Py_�G�ǫk�����~��V��W5}�)vH���$s��K�Ț�S��C�5=�Y�y��xv7'0}7��|��އ�T3nX}�N�#���{|��Aۮ�~�b�%>�S.������C��#��s��ϢmB�vTǠ�4`#_�Du�:r���X6x�EX�aP5�K��}0R�I��7x���u���~ԲCU�"@d#(�x�*��J]�tS�!;�NΘP�J!���Xe�I��Fp�ѹ��0�BHA�J�|���CxLI=�a�z;Ż�·�d�����5�\h
��O;������X`�,f���^3Nf��ww*���	�؈��������*���Zf��d�A5��A���3�8*"��W+j	�M$�*�r�����w�r�|BCU��*"��J��a�������q�Ou%�-����
�6Ȏ h�ȹ-ɸ�vd9����,|�`������C$�nל*�V=��IM.����s|z�Gy����1!�O|�e<I�<Oy`s�e��=��.�L3�ow{0�D~�~ RI}w�M�N��e:���p�y�kv�xjV�u�R�bk��56w�zf�u|��;�:��_7�q��E����D�k^�9|���r:� ��9�� ^4�}k�D��PC�p�R
�	Sv�<��`�fw�;.K�8��E��]�rK0�����;��5���}�9�kp��up;7fp)bjn�gwT��^���T��@��mή���^��Ȧ���)c��9���a��}'�Ͳ���pg3~��7�J�)|�@j��oE�AWSޏT�z�g�of�Mg���P��愪z��2��"p��@�:EC����M�rv�I�5������oӏ����8oZ9�Eo8��F��9�T�d�6�zZ,G|��e,(ݠo$��b]��vν$�v�:��֓�)%��4��#�t�f7������/������{K�#	�oS����Ey���m����)V\���	�w�9Q50S.��6?�V�]�z�ܟff��Q����|�Մ�7W�&�CQ�;h���wF�<{���+&m�ݔ���f^CFm�2������Ud՞�+�u��B�x�s����i���ٹ�2�bw��Oy�uSp"*��P���<wfJ�h�6�=��Awm7�o6�0�/p=��8GL�$1�MQǃ#�Ī�1�{�[�৮�9yc-t��nQ�����c_H�//f}g�e:�tW;�s�i\�$;���g`�2ʰ�.�Xy�0>n��r�mZ���� C���3�թ|��{�h�YՖ-3Z����Uv���X[��U�%��y��.��O���w7��]��Jɯ(v��������q�	�A%�g��ή��X�r�������]V���$�K�������_[�]:�'4�r���ٯ��1��[m�[0^օi�ʾ/��oSt:7���Lq_D}�����M]G蟾�����"��}*.�sg����m!m5�X2�fT깖"sz����N� ���ѝ�z�f<"#�҉w]��_�͞��F�z��M/C��J�7v���<�O����N�n,��� h�	��[�b�ߖC�Jò�g��O\�`�IrϢ)��� ;S�T�M1��v���R�z��kʥ�k��o���j��~��@}Z˯=9�=q4l)kjf����{/6ϧ�K�Kg�]UJ'�z9[q�.�/�p��'��x
w+9퀲�����Qƴ�<��2o�{�QÔ���� �D�1EPG�V���Esn����`��X(��Q���֩kTA3+�ժ%�-U�b��()
"ۅ�TTZ�,�X�g�]�]9���^���o�u��#l��;:���Y�aݐ1;)��Zj�����#!��p���P�(�Yz�Мh�����Y�ݷWڳzp��$�M���E��>�>�}��+t��8���ȁP��7׎�,s��j�I�2��O,��W�_9���fwk���lf(B���f�䥋Ɵ����^�z��V��3pUu5�͚yG* �}��7��6%.��.�/*$@��M֗��BQ�'5�}rC�u0���%��-4��/s�g�  �+�:1m�Ulxed#;T��ģ,������9��̺��Yw2��i4-�S9ˀ8����{�vJ7O*l��lcs8�%r�lL�s{|AطcfҪ���ZA�1�k�%�|4R��b�|�Xb]��&ۆ���j�^��]P`OD�!.ۘfF$PD���֍��y�[v-�ǁ�&��۴�R���T���S$�\%̛�(��9���5
��j-
��^Ś�=����u�y��s�>�������j��}������ �����kVU��
����/2�VT�P��!�T��Ε��h���r��|���[>=�*��G�o*B(.�c�E�u(�g�=.{N���q*���  N��j����.� ��x|��L��d�.��j]�w��b�Fls��7��wu>(��^���g\� �����v�5�Ď�0�J��k�)Oc�����W���v�������@�잼��7�M�`Q��I�5�[B3Uزe�,�t��T[�C
��Η�����N��V+3��uz�����]^X�{��y_p�l�6�7�%��]y�at��5������3�����L!|*xէV:�E�bW���V�P��z�-+���w��$���3���r�S��QvV�\K�3sqD�`��[v�қ���c�g�����v|��#�Ŏd���*<��v*�����A�`�}1C�S���)RB�=DϮ�w{Om������U��T2ob&�F�;�%Xb�º���36����Zt�K>PRТ��I�5����=߾��x�I�@�٭��~NI��¾��gǖn[���&�W�5Owr��V�#�i�� �Q?��;r���w����<��hE=�>��{2��ŗ��	�{D���n�LYh[�2;B���:/�Wo��J���L�< :%��k"��~��LCy�f�8f�-�޴er��)fB��5�p�w�g�O�\�{`�_9���y�W"�\�n0cJ�E+U�(�q���8{]�[�@����ڂ���^�p�F�l����]�|k�
�7�r�L^d�G��UǺps:�@&�57StcY�jo&��P�b�;��ϵD��:�V��%#W�ǁ������{EZ��ܹ`	������c۷� >�|�a�����7�8�&]<	P��}�
m�
���w3'��
R�H{��$��F2��8z{+���ŧ[\p�X꜏�U��A��^����\������ẓw��^��=�Y'b�.k���iU��9�St���f�`��͜ߙ��雹�s	�F���aS��ٗ��<Wf�����/�E���	N틉zȥQ.3�pX���������ח���֏��>����z��Y��a��,Y�L(!�N�=7z��*�h��M���(��rD�I�$ ���zmo�q�fzک.�m	C�2��}%Z��rl�ki\=�w;���ȴ�+�|UUޡ��uͮ],'h��ؔz�n������g��$���5Cv��ї���T�68?p�����q��Ď}�����Ln@=��;n�*�W\�f�q@��gs�ke�մc�_y���̌��VF7�e�ȏ�>=�J�%�0�O�G�%�����Y���=Z��W�m�1���<�����;:���^ޖ=�w��{+M�g�H�f(v��b����א�u�c���:��W\N'���6i����87�����H�mEM�M�y��W;�L萃���y��7�}�O^�j\/Uݸ�C������51�<i�޾ǯ���<�ؠ�a�����Y&�M}���`�n$K��]���(KN��s��=j���3�љ�|@D�
5�\өT�k�J�\�F1�,`��F�$H�
E�E�.`U�lBق*�c+%[jR�BO��d�$o8pf����Veh����NG�}I>��w�Fhn��U�#/�4���NQ�e�-�u��d_m4��R������6�7�L�c�#^�׌����G���ph�TsH�>�1Vz�3ٝ�l�����x��������4��`"������0h��M�7ѯ;��j$�0�wP��W9N����/aK�u�ҭ�U��{��u�1��^O�n���ޤ�|�O޺������ܳ�ȵ�����$�^\ڌ�:s��=���yA�'�Or�Y���K��������)tfb~����&��u�+�v�=f�v����{�{ړ���̓�Ld(q��$�Wu���w;(fqg{;�'�*R�1W���eT&�����)x�`kt�\�z��~�Hu���t�������IGEr)Xa4�22 Ud3U֒��K�:�>�W���.�ʷA+1y�ݥ�^'�j󬍑�+y��*j�j^��N��s�����X���ۃ�ΚE�
V�N�����E�'M���:W�;#�WW�e�.�m:�[��g=�ץ`.��ە]��p�k�v௫��Ih���rx��;#{>�t�r��)ʸ�.3)�6flT	w��j����)0�,����#ʕ�i�H�x-;��e��+��r1���+n�n3ѫ6Ff�̋���b�Gb�\1��+�n$�a�������DK]ŷ:�䯅4�fʔpe�yY~�ti]���0n�t�p4�rJy?G�Ҧ&���о�p�]�P/�l�=������N�b�&��~κl+������\�m�mj�r~j������5����ܽ��m���9{�:��ӥ��0�$�Xa����s��Y6����f�գ3�ة����t�k8���GP<�#��J=V6(޺I�G^�\!���n��
�bza�3�^�]C�M�����_� >��E�:��M}���d7�TW0��gZ&uL��Z��΄�H�KF�Y�k��@���Cid}��pBm�^��ꎋw$>���%�`y�x]tBc����Q͙Kc���@�+�	�>��$}hF�N�q�n����Х��/to����%)�0�X4o���e�Gz�V�ݰ�>r��Vn����t7jF��Yr�p��>�3ڪS� ]mGpA~!g�A�w�r)�T=�E�s�u��%��p�钿U��}�L1dU�f�Z]R�Nr�#{v��'���H;�����T����ݼ����G��E�k�%��c~՝����|�B"[�`]kCHi�Bb��"�mc"�)�K��u�u���3}���o���b��:�˭��Il�ò	�M�U9Q��ڧ/��6�t5���X���kv���Y���ۢݬ�wݫ���Q�t�I}{9kͭr���Z�O��\�O5T��f�M2�X��7�0RO��ԝ�Y~�V���;Z���M���3qF]����]��5z��W3��u� O'��!H�S���}1ₑ�Շ�S��w���y��a��E��i���C����>����tU|�j�K��H>�������";�+�~7�� mJ��L��v��5��w�De�g`�� ��4m��^mY�?pz�v��1{`��K�n���L�Ý+�;�:*�Y�О:+��)R��C^��]�Ρ\�d}-��k�D�[�ͮ�I����EZ���#��q\Mx�O���$�9��a���F�a�U��bzN�b�o�z���99�^��%u�]�3*�
�φ��
�վ3���4.mϲ�;'Sy
�3V)�WVU�	a2�a��Ύ��A"-�I��ʬ���i�Z�v�ή�m�ʸ݁�Tԍނ��������8~#�V�P����������%E_;�Dr���:�ޚ 9�QNt����z� j�쯺3)to��o��;����Y.�c<d* ��4Sh��WR���f�s7�\A)J�Z-��c+Q�W2��7P�XB]@L%�k��7a~$��2N8�S�7�(FG$Dho��|�h"���elS:��p(�40BeQ[����7�I� ��)"�/�%ꎱ�����y]v*e(����||޷�zٵI�ٔ�z�3��z�vCATW�5�Eб�C��S���BA�[����� �����鮊�F�	�!i7�5��I�ڻjE������|ky	 Z.*��? ��T� ���}2h�(�í�f���&�}�v�$Q啴��"��`�4M&��K�P�B�X�)��TU����[,Bm�`���1@��3=�;��Wi�a�3p��~+&��k��=����7}�Ή[��b�-�{R}ݢQݹqEFt[��oz�^�Cy<�ɽ�*�gj��9�'��t=�A[BSu��U�:�\�����w��t�,t�\��:+N�Qv���ۇc=T�e����ANp�e�-/�	�.���O"�;�۵���,�}�-��+pI��wCo0[����s��ov�95�7bm�uf�_L����m-,*X�� aY�P����V'�kw�O�1��Ƈ=�������#z&��7{�0��6�#i8x`@�z�r��	��Y�,Z.��Xy�����qbrcC��0�ݼ��E�U���׌�H=Y4��!w�S��+�)�b�*7�,{rӱp:�2�=rv���\.����2�v�Z��V�G]���F�v��d�p5�R�Т����J�e��]t��t�ܻ��>ŏgE��F�Z6T��1U��}ݥ���R`X��9��w}�WW$t��	�w.Ö��L�BF��[��u�8d=�]r]����=�r¦�ݣ\�;R�p'GͬɚW2�WSIq��b`���W�:�Fw(��C�-&mA]`n;�a�	�(;���@���dT2����Q���vA�B=`�À :mIǩԗGh rZ��3x�8A�rvp]�IGX�oBB��{�m���o�a�0g�Q�؎mĲ����rHl�B. �k�����[��Eg�@�a�iR��tB:+�o�Z��.4�IV;��^��X�r�QܒI$�I$�I$�I$�I����@�Q>.�B��$�7ǷG��u���p�`йYXz��{2*��f�eۃJ�g�#S�,�ǳ��(���Ǟ^����5b��갈�g���fv����y��>���e�
�Hfc�B%֍��[��U��{K�hh�Dq8�=��۶돔��Jnw����? �Q�!��\y�̝�.�����_v�V�߹=�s%��[ߢ^�HpDA�*��q����]Zu��ޯR�t�bXO�lْ3w���S}��c2I�G�?1��}��u� �s�=Z[��qT�Wެ�&���EyN)���{n@�t�-�����pu����r��|{�`ff���l[�q���c"hnEk��M�3/T�=�P����>���e����\�t��E#�t�g�U��˨��������{���M�[}���7<K	�)k�T��Xfjjn3d$*BEPX��, c\��C�L�Dce�Z�Ԕ[
���TĪK`��9�}����j޻Gd/3Yr���ֺs�a}�6��JS�`�]�����CBiͱ�w�{��3JH5����gG;%������X�s���I���J�굑���P3`g���\R\:�V��zt8���J��~����~v8�%��Ў�i�p"�}}�;�)�ڇݢ<4֮�J��]8I�g���_y�&{����oo�����2�A��o0�]��g�����߳�߾�ǝ��w��������!�xtr���Kl��~��*3RK5����i��,�
�
�r�_�1V���C5��p[� ����Ռϟ����q��o����u�&�����6��3��r<e�c��B6X��S3���I�W�U`<�A=�׿l���}�k���N����^������U��v*�R8�M�u�T��uL�崾��$^��ão;b��Z�C�򣇷Gr�!wC8��LvJGG#(�C\���Qb�#v�����r7Ʃ3��֘=qR�1��Q;��]�\^�[|�e������ӍOw'b�K��hP��o�M���U�bK�Ks����κ���S�ȇ���m!�ԗ��Ku/1�sީ�c<>�}���f�ˀ�4�)&�Z:g�X4"����_f���Ř����`̞�Tu.����"vz᯾��W\�1Jbu��: ���ĭ�n��(W��N��¾>�R������OL߻�~q�{����t�)��o�x�[��Jb��O2q�ڵz�j�I�u�����H�JW��*�{n����UZ��7%I6T��rX�7=L>��e]z�����ҼFl�|��XXfd�R�������q>=<�u��(X�;�U�A��H�֭���L�:���R���᮱F�2T�v�෸w�a�ɮL;����ܡC�#W� ���wu��E�A�=}B��>����v%Ͼ����'�_�SS�w��+.��m�S)9�I�:��:��2���>G��ﲅ{Pk`r�RYM��f��~�aX��͋\�O����h.�;�ile�FL�ᶚ��F���ל71��,h����X��yꗋE=Ԅ��uV@�r��\�Q�9hƬ�fv��}u��=�(@p�J9GJ�b>�����l^��}8���T���o�!խ!��^Sy�&��u(=R��SԺ@�O�w����s g�.k��7��5�F�T���7 �!u�e��R��H�D�T�e� �����9�\(������\ּ�Ɍ�.����%G1��XY��W]ˮ�W�6����Z��|p���
;y'\z�f�b�8�ײX�'%8�jg�v_�hĻ���Ba��[�[7�א�}��jn�y[�N��Z����h_]�m�sm<�vz���U�;!�.��p���O�̃�l��VGj��_&�R�U�-[v��3 �z�������Ͻ��߼�vq���}�5l��M�m�c�R�s���P'9�@i�1گR=1�F��#Z�[{`�Pvv������Ɍ�M8�H���Ga���:0��}���c����u{��G�r�x�ѯ�;�xeiJ�6�@�¦=��A����KT��j�D�Kk��}Y{��f���m̕�[u�|wuHPbu���SC�}^����/�+���O`#$�M+H|�'�N�DX����b*��$R2�'���g�o�����s"�n��s����P�)����b4{��)6�݇5Pf����ب��鱫*�Srmk�􎆴�M��*����J¾�����[��GC.U]�V�%e��m2W�GOI"+;��~���zs����xS�)��}��ێ�]����[��R� P'<��b]9�^go��5�}G�^�OdT��÷@���%��咍���̄����W,5��訌YS��|��}-����yg� <�~R�_�1QfR�!_���[� ���.�wa46W�Xq��DD'ͪ����p� HǠ&�B��z���]mC��{��֖CglC�#j;6�+{�j���YFP"Z��9�DGO�N�+����B���^oe/��ϟ��O|Ý>����g�=�Y�N ��w�m1�Y��DYJ���#�CD%`
Đ�R��\ߝ/��y�yr� ̔Fi��]��&�{׼��2ҷ͜;�r���:9w�*�����Z:�����#3�emL�����|��=�Oyޓ��^�>��U_��Fw�j��#h�&q�6g���4+����3��wS��t��.�2���N
��}C��wJ���Q��{�޻�;����������zQU��e�єY}���Lv��3����4��v�sxx�q=)�F�E�K&����O���>�ƳO/��| ��I�������[��ؗ}��j(h�{.mGn�z�37�S7�
fz�`��������α
�ۯWL���.�Ͼ:b&O�S:y+����4��b�����F)�u6'�T��T8�Q�=9�C��&�`�}����S'�漸�aB�������M)snOK#9��f��։NDfB;�Q��732��GS䄡}����51�2�.�,��?#�̓j!|룴K�uI:��mwl��X	��êt�:z����=�ÕM�\���]����,�{�Q���m���T� ˟����2�CP�\N�gQqǢy��x�@��O����#B�|�݅Y9�m{�G^����w���A���%�}�n��q5픙��}w]�"e���m�Q�/B}>��H)���F3@�mL��z���͜d>�L�}�&���+�9#(�өP���
9�F���ƴk�a$��C�3�����}w��TyP�J�i�(W|��.6�s-�u4/֤�����>�%�r����3�W��n�����^�w��Ih�����A��}1м0j����������XY�֊(���)!� `��ko	v���=������gWӞk<V8]k6���{޴z-t�ˎ�w�^T�T��o��ܤO!A��w�v_xb�Y;�����U���]w�]5����w ظZ"�O�NKh����X�m�qv�Ĉ����T�K�p���Fs|>T�s�����{�| �<sM�=F��4o�Sr�j�BK�X�A�=��ՕwV�]9c��sE�K��oݤ��..~��|(�Nzt.E�J������۵�%��}��{wN.�n�WK���8p�XS�q��&}	St���:�<ۅ�L���a�|e{5?-�G�2�H�}����c�z�	���XMA�@�\�*z�w�ܻ�֋¢����涾���zoRqjK����O���h}��Y~��K%@B���'F=�B���Ƴ� r�K��m-�Gq�F�e�:�_a�����i{���vړ��;X[�=M�RP����7��]�,l����k��^��1xW��>�o�J���uWb����.>���m�Y}2���v`��ބ賈���V"��6�L��]<[�鍷T�k��>�?J�§��u@xN�G��q��j�Q�0>���0Q�fE.�-㝼��� >��R���:٪zz�	��ߪ;J#>��z�b�{x��x7u���C�{}���XOg^ʺ]���)-j͇z�?KYC *5F(�'�1����^4�t6}oK�]��:-m>��UW�[��վe]��zL�u��÷��;�/�[�:b�39x�0Ei7{Қ���}۾k=������$���H�O���O��B$��-��$?� Bh`@��t��	(HHE��� 5��߰�$��?�$�	$����!$��ס�O�?����!$��o���������O��$�	$d� )$ $�����$�	$�g����II��������$I&�7�Ē$��II��II��k	$I'�_�o��滛4j@���H�O�?_���	 BI?�@��}��׆��w4?�	 BI3i�p?�����$�	$��XII������d�Mf���`��~�A@���@ ܟ}������{V���h	��Jٵ���H�,-E�,�HT�EL��,�B[�9�@m,#V֚�P��Imbf�PT�`�6+l @�%A%(J�� lj(" �UB��!���������"��T����K`5C�9)V�)T�[VVZ�+Ki��M����SU6�Z����
V�}: �s6�V�d�f�lfZի[6kws���"��$i���T�;�k6t�Ti�Ctr��� �E�Ҙ�G      �     " _U���S��C�9��n�Z&��m���4]�r�f�63�����Ƶ���w%���{=أ�v׻s͑f���f�n�����n�h�6ڌ�Z�Y��UKZQJT�N��t껻��۶wn��fֳ\��u��b�u��Ӣ�r����أ-u7gD�&���m�̡Ѻ�h�[j���]�-�[k[���ܳf�5�ۛ�KZ�[KUHV�B���YYC�vn7mt�t��WCNm�unk@�WWӮ۶׮��Uqι7w��UΓ��͵S:�46���ղ�m]Y�m�ݛ�;%hأP0�U)���k]�a��ASʩr��wXrMm��S����軻vn��#�6���@���[h;�:������,m��(F�QJ�Á�N��:��V��:]���wv�m;8�;��v8)#���wkZ[#��Z�pյ�n͡��ֺ�t��IʢY���EU)I�u���ê#�Xa���aպln[n��]NqlWvS�\��;���N�4��uWu)�t9Ѻ۷j��}�RM�R�l�QS�ҍm�d�$�J0�:5�ږ���;�u�۷l�`5�;vqr��u'4��K��]�]��Ύv�#�1#wn��7(T���B�Q�쀧ݺ`ކ˴\�캫��4���ݥ3�gw6\wwe�GI��{z�n�f��륰�۬���\٣t������\�n�WZR�_[��R�Xԥ�[B�^�ʌ�K��.]��X�v3�kgtݕ@u�sN�}z��SN�Y6e�g�c�M��/rvU��a;n;�h�m&���m�-5� 6�eJ� @ "��I)R�   UO���1U�A�14b*�	)U � E=�	�T   ����"mSjdi�L�)����G��o5xxcE]?9�s�ī�d��r8UAk�l�;Lq'�9�� " DD?H�"DD�� @�� D@���Q �
� ���� "!��D " DD�_~�� ����!�\�6?�_�Io�%	����fn��n��Ҹ6b���I���BkH��ͼ���%�?����0j9�td���ؚ����^����\1������z�z��9K�&��wS^�H�[�@�*�r����ma1K,�ڎ�t��
8�c�wh��g+������8_�h��h�a�wg����wEQ�H��V/@k2� ���DfQ��R�]�o�
�r!�v���Hn�;�F-D�e<9�)ъ�V.�]��%�]ۚ{��� �}
¢��MC�*J:����Xk'f��BH ��D"$ #F	 ���B�Ջ���/6��^��Ι]/�\Fm��cw5�C5b�B���e$]Av�x��t�.����"�r	tr�+6�[Ql���۽��;k�x�D����L�"�b�� d�Eǚ��D����De#�!7�\P������ʎ��wOv$�����v+�U�r���ǽ�w���6)d�O���[j��rʃ��J�%��ܪ7W�ݠg�.�m�*k��Y0cr[.$,E�V�1��t�)A^4�&��p�S���+=.:2�j�.���p�y�E5�V���r=- �t��ҁ����H�q��\ ��ۄP����%�`ɹ\!����h\Y���&�v+��W7�]���������#sS�l��o~�X�>��+��*w��[W��ct*V��v�g(qE���rū���>�0[+uDm�=ҵ�S�M׭K�k{���U=��րy�[��mkгhԻ��zє��I����
�
#��3]� ���v)��{���r�,�mF�!h��V{0ET�2*�]7F	іVMl���T+��A��*�cB�� ǰ�E��P�M�Ң�.Q��a{f�j�ā�X��AR,�hL�	�r�ܗ�Dvd�i�I ����C��Մ�ܦ������t'Bft�Zp�n�������0b(jۛ�ܷ�]�kp�!�uj���#Y�9	p�Ae���ʴ�2p��3:��:A��a�D���b�Q�֓6�Է��!��w��ө�칐�{���7f��x˺��j�	�X�
�R��X��<��܎��Q�ek�gU�l�i�Sc.�Rw\�O1E�n�SU!z y�Ǎ��u�F�_q�`�XM��4�R�ˉ���@f���J��ݰM<����r������s2:Ef�hU��Q���VAul�i~��J�t%��q���{V�5�2u��!v��%l�
�x�T���z/q͌��d���8IMoL�4��x2Z/1�	n(�p8Fdj[�6@��@�Dʚ"O*AzZ;�Ҡ́��[�F/AGhC��fU�z3�n�C ��� �N�˼t��;)��Ko6sd]e�w:�t/1�I�CO6�K�u-cw�4879;Q��2$��D��V�$�:�n�� X1@āGj��d��9 ֻ3�+'���PT��v�VAq�b���0JQ]�D�F�6۵��5�Nuq˃�5���v�QDB���k�P��&Yr؆�+Mn�Ԋx���Q���ޝ:J�^���Sm@񚟵XE�su0�wKw*(U�j0��-Lˣ}ͽ�|E���f�\h:�$S̕s��EbF�"���/�fS�2;.��d��wjv�J/3vĪSyHf6�F�wI[�JT˱w�s
u�����4�l���4��Ar���r��&5�6����g)�5��X ���Z����Zw�l�	�ղ�X]���cU2�s�C�2ń�k؆�����HYZ����(�?�v_[�˺y@A���L��	V��Yp�$`%!�S�3�����gHs�h��%]�J�ҩ�IK#�%RR��Up�MIe�F��� 3z�N��+�at1_��2QLmܼ.ƽ2Z�GRa�V��2��J�{/&J
n�������_'z���a<��]�A�T��J'��F�`e��du�
�;�؏I�uad*w����a]�̼;�,�b1�F 2  a��@�`
""0��� �,�8�"�@� q	�����Y�]�<�r��b7@�KQ�+=[��)�]8 �DTm��y��� ��.b�V����zH6��1߰	�`����;o�+�y2�N�[�F�Z�uB�^�K��������˄>ra�]�c�K�m�WR�aY�'ZݮƂ�MSS�1�����s�t{j$2+�B�Kmu�P�8"�A��Y��J"�u�d����ٺ�It��f�j����UՌ�0����#I'
��Y��q���q�Q��L
7J��y�U�onS�	�U(*�����6fNU���iu��4�9vv��p���Q�qm$�0� X�r���h��&�VVfS
�	���U-�����Y?���)^��M��rM�/
�3�:��rQj����"3p ��B��U�Oj��*b�3I.޵Q&6��YՐ�����:�T&c4��`�C(Y�z(-.��v3Q�T����)W	wyL��U���th
 !�@Uo�ܖ�O+P1�nm'��kc$��1:��y;w�P��)���l/ � 4~)f*Õ1��1m��E���X���Dn*nVY�7R[!Z�,�b.�ƴٸݣOhŖ��V�:e�K�5ee�@�(��M�c�iZk^8V��U8�)�{��jNr� ��X�� ]e^e��U'pUg:.d*(��I�x�E7B*F�X���(�9K�[�֯�]&�yi�XV?%�v^�B��9����n=�J�B���,f� ��4��Ml�Y����eCK�7 �ve�N�hG��m����/6�7c	�Z��8I�����n�oC�P��
�mm��w�L��d�v�%���*�\�R�N���QX�w���hT�
�v(�F��b�Yu��E�C)7b����&����<=�ڕ��8P�oUeL,��\�J͘DmVK���B�{f+�*�hQ��Q�Au5[	Շ2�H�ǅ�^� �ne���w+u{B��2���	�X�1zԼ�k,]����ެxw*�ن�q�/��C[u�J�����M���4l�M�4nd��R�&Am[w���N��L��.S,\�T-[��^;�71���vz� ��Ԧ�+ep��	�v�ͺ�t޷h�Å�ݨ���ΊAn��Ú7+%��p��t�Z��*�oL��3ndyoj�
�2@ZF�t�d��,4�g:So9f��:�jޑF��$��,U�4+n��+c�-4*��#Z��h�k:�z�Â�5v�/u�	�[&�kjh�oqܭd?қo5�jz.'��Sh8әj��b�rY�bҬ�xc9�V�V�8ݽ�C
�V�2�X2�,�XP��d�3r��uHt ʀ0�v�QV�-G�NV}�q��t�q��۪j6�e��V��]eZ�*��-���w(%M�x%�r�P�4H�2�kh�2핀&1m*�KIA���",V*�
�35y4�F �;5����[e��gX��&5�q$ ,�S�@� a(�0.�X�:t)���«`���N�i��u��+^��(�k^��c-��A`�ݹ��p�O�R�l��T��Da�0Eڞ��٢�ȞU���cbe������Գ��K+K�d(���d�@�
��IV�V��r�ј�Fݱy��n;��i�����C,]7��+(���yb��7e,��".Ccj9���uʌ�M�������]�%[&�4~X�Av�je7���^K�4�[�4�r�kt��J�
Ȼɴk����DեbVŚ��C����Ғ�P�KV��v��h�.�Tˍ�J1[���@�ٿوCY�cWy�!.ș���,Lyi����&್6�oI�ҝ�P����[ub��I�ȉ�l���K`�m�3�+��(KGE
�H���6�gsh��d��d���"CܻA�Ơ�G�.�b�����q�A.����l"�8��Y��Mٳ��Mט�L�9��Y�S7N�B��qCgl�J�:{��@��q�RY��H���=d���4E@�Z��+HCV�k��/:�;.�͖���b�X��d5�yJSŘ%,��ܵve0��{v����U��z[GWL��D�ݚ$[���b�Y��=qm3��Հ%E��A�Ա7375�`j��ʈ8�tTd:�pm9�"IъWx�Ӈt	K������e���h���])ViM��'W2��3*���J�9B�ࡈ��Ȥksr�����Z���=�^�AT��%��LH�ۚqҹ��?������d�f�&�Kq�N���R�FH<�T�z.���(�,��u����/)��:�
Vn����`}p���׮��бV�:�eƳ�ׁ�ä.��JX��G�Q0��3�1w1-&��֤�9=�f�u\��h�]ƬD�201٭F�R��m݊��R�,�΍�OE=��7�u����p�9�3�eB�DBs�E5�*��Gk��3-V[�7���Ĳ {y-�y��u��A�dv��,;����.�_>M[{�N���tn�i=�U�i	2b��Qe��@Q�I���E�O
�����"�Q�1�(��j��w`�����ObB){B�5�w��ʻ�gxv���!��*d��B��<)W�6w��uew�VʸJ,�4.M�T���%�v �u���t��UhՖ�H&�
P�+��A
�gJE�d�$� X�а [��,+bf���ޮ'��ܚ�GL�S��d �i���Iv�76�I-ɪ��&tj����+8�����c�l�X8�i�M�J�PT�C-�F�r�Y��DU�U�A���(Z��j���53wy��,�����|	�HibκX���â���R"����X����*_��j̣H7�7#r�-���c	AA��e(f����9 �SvA�Pʻn����*P�DfU��۝��[�a��)T�1m6���'pV&&�Q�[jR�u���4� �e�)"qĆ�(�6��՜z�X���n	�y��l�ۑ��@m�u���:�hu��� ǪZ-F݆*7rD�d��v]�xʱCuQ� �ʺE��@ԅi��	���h���M�XD��v?j@m�f���ȗcZf�W�D!�
�u<�ǲ~�V��pdW� 䬫d�����7���]�wGD��&v�I�P�ͼ���k�
6��F�V#n�����SMO�fR9�0�E�� ����l���,L�_�a�Yc&R��A��b-����y-1r�\�@M�Ǹ��XbF��mn:{qf�WM�8֫�Cmf����&��̦*����`��ъ����E��J��<�f�i����%7D��c�i�z�S�[���������ʡ+u#2Km滪�~'�v0"�5���hEbM�W��Xu㟳,�:+,0��b�	��Ym`�ݺ(���h�N����Ѻۚ+�!&Xm�
��މѥC	ǹu+�4Ӳao]#uu�&����$�����1� ���fe���F��Kp�W�=8i��jeè�5b:X�1��o�¯3;te@�o� ]�y��i�ǥ�`�����JM �2�m1 P�ҟ^A-�J�
vk:�:{�C�Z�<��kP�Z;b[��`*�ݰj��h�@@�]�v�犱��3+�ɗ5n��"M�����q�K�Ո�L6����C�}2����\r�+1@�AU��S�-h�˂��tw&f2ӊ(�5�5�*i��իuX&��72��%VZ�͹f޶��R�1�� A�J��@�h2- �ui��f�ע��S] A&F@�bRX(ˬ5����SQ틗���t����7�i� *�>�K�䮋W�ƀ��"�v�p%d]	�A ����i�p�f<����� ��͌-M������w��7n��D��i�H����n"���Y�ҙʑt�n�Sr�ѹt�+ۭxۈ�՘
�sD�I���Vh�M���&;�vƮȵ��B��Z�+bw��8���Hg�٘6�µEW/!զj�����DP�Q�͒�p#�i�(��9h�� ����{�T�8��8�������(d�V;�����JI,e���jִ28m�i�f�2\{`��7"BLw�9:�f�8�M&T��Jm��^��y	+C_�W{�0�ɥU�3*�"���F`����N��&�3������73� �ׅpm��Xq1��X�ӳ!�v����ޠ��3*IoF��&��!e7��K4�nk*�5c����.P5�IN
�zJcS&�75�4��&�-{��i�v�r��R0P��A��D�?:��\��[�A=��?b���K��P)��ux��hbjS%Z�x���w+7��7W3����F�C��TFX�q�/CG�u�f;�<�(Գ*+�!"s�%D�[6̫m�1p���mc7��MZը]i36ئ0�(�P_�&r��K�5�B
(���H�se:3�4;5��:{Yu.��XY���hC�phwiң����Ƶm�{�����(5b��38�����	R�����u���]c���fH@����ͭwM8��6���T�H
�����gs��.I�e
۫��h����܅����E�e�e#0�7��wD3GAs9�,,4�E��WN�mӠ6w WRt��T-vE�,f�7��A��9���凂�zh�Yab��v�9��\V�-<V�U��*i��u�Ţ����Y��B׸n�U��;�I�Ĩ�-�=��R\D`e]3�,�l��*,�l
���A��w2^���;��8EF��f:�{���Ў��鸤�%8��H�ϝs*�wZJn���/�8]ww~�Ǭ
=x�6�/T��7�H�I�#}$o����>�I'wt�H�I�$}$�����7�H�I�#}$o����>�F�H�I}$�����7�F�H�I�$}$�����7�H�I�#I�<ߤ��w��.=H&D�%�I%�'Z{c����|�Ki�c�(���MK�uѹQ��Z�Rm5�P)��5rg����N�o��i�G+�����i�`�"F�����6is���^�0�y)���L����z�67F됶m�̈�΍��j$���us��}N�s�}ʹo;u�������"I��b��YŠ ��~��u��$����L��|��DY��j��\l�@��yX$GGĴ��*I��q���'p��No:�W[�WA�Eu�N�ʲ/i�%�
�V�>w}�k�:�$�^(Ak �೻�2ـ�%��/iq}��$����i�J����<�_%b�%���tK]���^����]p�Wsfw��6�ZoT](��n]��wj
]�%�g1��[4�Ž;8��7w��w�} �$�l�f匡D�)b;oG'�JU�\��u�Yh�b�����qIܕb��=D��P�B�x��zt����x�= Y�ؑ0��%7�7˴���v&Z�@;����Ů�C��e�rq��л�H�n�n<�Pܡ�y��Y�[��poCQ�����T׼Y�����ˍ��6�3�Nٽ������s:Nn>�N�ư[�/���zwI.sm���\b̌��s��P��K�V�oU�㚛�(�rv9��i]˓d�gm���5����D�$Rc�}{ET�U�h�tr���V0�O�zr��{1]���^�d��6TX����fD�oR��w�;�#� P�ά�|�L�dq���7Pڻ�u�Tl` ]�G��MO*]�̉Q�X���ś	~̰eQpdL���.��NM��9h{��#b�����&:]˻[g����U��u�%Fur3M��h;t�Ʒ��C�xh=ڸ.��H>��ղ���|��x��+��a�f!W�孫�������q��_ou���|zeou�7֒���y�z�+��s0������0�׉�:����k��׸��y���9ͣ���q#^qRhS��5�^^�=5�h��z1j� �m�wv��I%hk]0�Y[�$�t�">�Χfms��V�'W�C�0Y�[�z��A�z�z�q�C�}���"��:#h���t�T�!�F(��O�C�y�Ktΰ� P��bz{^�<lFve�)�0�:w��ݣ��������5q�ބq��«�uwyLl%�6�Šhg{
]h;|N���r�f�8˷vЊ�tI^������ֳ5f��]����&x��P;6[�-wrY��7���۽�P6j{�?����Y�u-�nH�`E��.�F=̈́��>į��oq�\(dv��wF��d��l�y�g8�v�t�k	ԣҸ�Ɛy9�)����6C'�gMҕ^�S��8n�яk��y����J	�o)n��ky�V��A(�Abۀu�m��٤Z�����]�)uԅ�z(���tpk3޾��R��i}����u��Ǻ��^
�TKwt�i&��bv0�Ǩq�3I�B����S�������t�v�"O:l�r�:K�=6P]o�wc[�|����f��j��9慄��&&�1�B�_s��Ye5���6�Z;�l�[;�Y+��U1f�RVW9��i�*%���3G�!'�	�|"є��+�˽&���\�u��+{EZ�u�t��UJ�Ø�p!�z�.�MR�;���򦊏�5nv��.n!.B���7j)�[XywS	�O.��m�N�2*�
�F,��A� ���z��wk]��7�pt�۫1umY�v��g�ac&�O�<�}���V�����q�q�̧��lST���i��έ�D�ŻRii6��J�u�IÖj�ԛ"�!t(��Rw}�D��5%�`d�ܜov��7�'ϖ�"�9���t��v�Ј���]d����,1�d9�&���;kk�oZ�wx4����� ��ʮCz�ʽ۩j��r�j�z1�+�Wl'�tĒY�3:�ܽi�(��8�a�X�z��'�iKES��w�87n��M>�nL���M�:��R��Ҡ�wyn�(e��J�y�m�⛮�� �YD��$g^����I�����=���*��;7�1$���C�h�p�w��f[j�jT����ڶw���B<��9���lܕ/}�=kF��G]a�{��2�ݡ��gI�,,���ц�Q����ˑqٳ^Iӊٱ2�dB�qЧtؾ=Ќ�õù]Zٖ���8�?9>@�-�X^�ə�0�*����3{���Q%G��7��8�1�����R�<��3�4�N��j����V�n��>
�� p���3M��m�
C8h2�ZL�Ug��7-,A1ٴ�nK��w+k���y4�g�,ÝK:�,��K����EC��wV)`P�����dt`\& �����Ten%�r��O�V��;\�����e=�Th��mg	��nt�%��ݷ}D0y�v*��bDeM����n��Rr�:V�Y���8�VX�f殡]A�����^@�,o%��$/�i��\ox;��TqNB�pL�[��oi8�8 כ���]�1�j�é㊹a� =o(���D���UCy���DJ��d���Id���8������!�aKZ=cs]
́�Kw���Ij��,�t��]��6�4��g�N�F��w,veNjb���pu�����|�u\AV��)��<�:�r�{*�P�j��r�ܽ��Z��%�p��.�oA�K���ǣ[�O m��&�%K��D�9}G������VI�ƛ��["{��.F��t�[G�f�r�,����y�&���W|v�/��qK�խ������:�V�`��c�Za�lPV��g�;�X�Z���c�3���z��`��'��X���ݠ1b���E�n����[!�h kct�V9Vo�E�\��Ļ��O2����F����+\�3���H+�N��/-դ�Vt�]�y�ޤ�P�ׇ���O�e�.�%��H`�R��p|�^Td� �'8r���X�w���N���:���9`�����K�9л�ͫ�1��Ȝ�ٓ[9��m�ss�[��W9�Ԛ!z�����S���f��Ⱥ��K�2]��X�ᗷ&7�B|k��5Ǎu�@�Æ�@��:
����U���6�\j��͎��ԘB;��y�ށ�J�y�8j!ݮ�g�r����Z@���ѝW�:���#�iJT7Hn�'M�u\�=�}-˻�!�U �i���|o�ɹ8F��-<��ZnQ�Lݾ6 �&͈�r4�����Rm=��l�ڳF�;�O_	V�ڣ���Fl�����W��V�6I":f����o�ٛ���jgI�?qUE���1����f�|7�к�T�����}B�u��n[�ۦ������`�T��oD��l�5wt�Vp�o�<���ٕp��߭5m�c�t��
�2��[���ek��$䥔P�m��y��)�DF6���*WN9H�c�;Y����&D�6�ټ�F���!��V��N�h��Y�)S����<�lWe��80�}����f���!����^�Xy͂��i��Bn��Q��X}������x�=KL�}�q�\H��qM�`��[�[Ԭ�N��u�j�n̴�����N���f��m���f�����\������#��\ͦ�r�.�4����ፔ�lX�"浸��e�	�Avv>=i��MC�)��v��'"���s��Aq��^Ю�m��
��t�a�l+��<pShV=�;-qSYm��7��ݣ�.|P�E����|�L�z���A��=����]4^�鵲S�l��-kE0�o=WWQd�t���͞{����O��:�ݮ��g,�+X�,�B�o�(��{���3,���U�e������&�L��Y5�����֣��<I�ɒ�[[)�f��t���Z;Q�I��8s�f��鏶�hua������<)�pWeڒ횏���c"{�@�(uF�gL���v��{Ig�Wk+S��G�oh�hέa�⣃,�l�¯�j��O��[��G���,m՘�=Ȏغ �	�/v��^��(+M�\o]��� )�����|�ė�:^0�uͥ�vr�s�p<%�-����x��$0�]�y��ź�<�ə]IV��Π :.��2��xv��Ś���,ӓ=��*(����\�3Zȱg9��w�N ���.[�D{('$�s��A��:�r��X�h�������������b.V; ���${A���)go%֧�y�̂k�Ё� v�9]�A�&eh��g�PG�\5�M���׶9Wsڐu�%��]!�j��u�0�Ջ[B�fi�ͅ����p�T�<�����Qn�W�&5ܷ�Ϝ";��_n3@V�L��{�.~�'�fXŧ�_\�9\VTq��P�!G�s$<ga�Mٓ��f7D�u��}��q�7�qF�5�g+� їn���lվ\�n���9dlp�:)�\�Q�:ܼ
'Yk���������9�{����o8��q<	�[�ش��z���: ��wvWC�5�~�(��j���;��JD�#Bgs�9ࣸ3j�t�O����`�,f�k;���N*�G^��]�ywrH���ePl��S��R�:�&�v�2]����@�9�QBd��x��v����ΝX�&#��+�²r��wu��&+2e��m4�Ыͼ��,�d��J�̺;��Be�L�f9�5)�~Sr�4kt�'-��],dt���[���`��I��/k�V�ؗ��J�;K3b�ݫd��պ[�ﺻ/�#�	�Z`b������u�D��0^�@��i��J���V�#��>k9�Z"h3�1���y&�Ъ#q�$���G^�n�Jeus��{|qMZI�dڼKw��k9I���y�\�"��({�h,R�����4��j\�F����%)9��Mͫ��ՙ/3���,���F�ы���8c	��+!Ĺ4�l;r$_!��D�R�r��TukK�K]R]q}v��\�Ƹ>`7���a�] or��M9�Ue��*p����ŷ����N�&��j�*�	(�� ����2�6; ݍ~���Ǹ2�_ss&��oJ!L�7��
\b�]���X�r�C���g�Y�Ҧ�Mb��
�וۓ��c}��AX퀯qSSLF�7�65V��@L)�U����P�\u�.�u�\�hT�-����̡vQ��6+�a��y[���/A�z��������TWv��TE���(+�[<�(��+M�ě���ݭ����Z������;Ph�𫸺�Tm���**�ZL��L�PZ�Ӈ#}����)�A�!E�e�G3��^��.���s�<U7{z	L���JԷx>۾���!{ι'����:�c@K\QD�J�㾢X;���L;%�:�\�GbG�t��$A�K��8���j�a�y�]�����AfaH���X*��E��7�����g�TG�7IKNJ��.h)�T뼊.���EX�0�d:&������.�͛���e�L�YY��uS�2��.k���]��4��A�^Wر��`�l�c}�}c?M=AC+v��抾�t&�u�oVu9��L��ĴO�g������$6�6| q�r�aZ ���H���NV�{y���
y*q]m_#*�bD+mn��y��խj��Z�`�ϝF�}z�u5�hL�adID��jeu����T�)e\�I��8�ڕ����*��Y$�K!�w+���7LѮ��X��+�B���镠=!r��|+:��_�~z>ɓz�ג8>�M��3�m雮���j�[	]���Q)��������u������n�+��ò+����enb�@�|$�8��z6V���N�+�W��I�z�����26u���Q��K��ܠH
VK��MOtþ�B�i&�^���k��S�W[}t��m�|�D���j�⺧u��Cz���s^sy�@;���-����q^���V�0p�r��]6�)�pX;���<��y�g��
݊�HgfU�Oj�5$�]�7[E�60�Ѯ9:6h���W^�ܻ=���V�Ken],��IV[�E�J����΅�b��E\O#��F轡�3�&�,@9���k�(��g�v���A��MVlY�WG5U����,h۔)�����a��YS�c�mrݾ�`Y�m%G�t!���\`v�w��%�A_mNI�^X/WQ�+Bs+���Ց�[���eV𻵭�u��o��}������µ�r�.W�
c�ǂ�/VKvN=�2������ܾ����BaWA#7N���֖���!��sz�	�2~�Ք� c���U��&��W={���U�W���6�oVڱ݇5�p�RD�{�qr�N�Z��s��E�ם��jN`SS�\N�Вc��-�Oq|�=�Z�������y�����Wn�Ql��Ѕ�.i��\��4��n;Y[�e#�ĸ3�u�/��|n��x�m.[|�k� �t;�Gw-�+�[+�\aU�"���qnRW2�쇦�N��lQ��DD�9�u�pP�Gll�8�e��W�M;1ba���6za���������&�+݂r�ܕ�0��Et|�Wo%CS����u�Z�!l��]�Q�^N7�r ���tR�5 5Jv���B�L�����u�L��p������κ&��Y��mJ�;��z)�:�\[2Y�����HҔp2uE�DF^�皵h�(v: ���/T�[�_�g>B�`]��dS��s'c�H���].�p���|��^�����8���E˻��
�yT�[a��ע� �Y%fH8��.���,U��^��s'A�AV�Z=7"�H�(�:T�g)����	�f�涯9��&EHb��m\��q��e(���j��q�;�P��1l����$[�7�Toѻ���Ԉ�ۈմvSU��e7>����������mx'����D���D��#` "" D! ��X��  B_��'{�i_Ϳ�#�6�Iq��;�>�K��G��q�'^s.��kyS-$��P�a֞�g�L|���6���J�>�aӷ�(�/�$����C^���Om'��W݁�:�ƿ���U���e�4��ܫK�y�9�@��dg:�l�S%'�2�*��, ����	ӆ���Z6�f>��m�]l���:�c,8.�Jޡ"����:S��\���b��>�;��J-q�MMV��(bF,���!�U�T���$\�V�*�wT6N�""K�]Y9� �L������4��SS��2g�u���I��98*ޢ9�.�?'0Vl]��@[�q�iU�޳�*�;����0���Ղ��a�D�ŧ��yCe�,�v&�7$���!s��7tQ���H��`���Ob���f'����������!��k:2Iw&��C�["�WM)�sw2�n�C��u�vx{��\io:s�Ö�J��\�ū����D+�g&��z*�jn���8>���V���sX�s�}�^�X�V��_Z����/�|I�5,�Vޡ��m����j�=�,4ȭ�r�r�����rѕ��Z����].ᘫ���m����|���Y.e=k6��8�̳z�v^o
V��Љ���	 "gu.F@;=�ow�5�كE�ҡV�}�.!vndB���uJ^Y;��Z�ō�� DD����n� �ؽ�\�G2�=�s�����
T|	y��Sa�ó���3���U����n>��JNd$�Q��q߷���\c� y��ۃ��]	��y�Y��L��/��ʛ+�g(�uC�+k�����PG2���ɁN�m������)��5c��\����7��cp�yu/K��Pt=^�>	«ZC\O�1�<w����o�-�z`֕,j��!��`�=<�����	M׀g�euѰ<q93}�"� ѡ-��H��a8 ��lfD0��h� h�'t� ��3���E�o'3��:�ٍ�

�1�4�3�m�j�OQy�Bf&��m���
5u�j���|M�B�^����X�����`�H�m����y��q�Z3eή�Λ��;��~O��I[�4�����rl{C�os�{�i����Q�z}�򇳨�^exx��;]̙�
H��ȓ�B5�t��,�~[���5�7{ӵ��x|z�";�r
x_�H��T���zt~�k*yW��ǵ�0	 ��E� ���;��.���:V�2E�6�˚�Av9y���� *B a �DBH��0��w�hL��9V#�OTl����Ԯ���oQ�R�!Y΂t��J��:v�_���f]#;��1ԵoZ��aC�s�ӕ���'����}�'�v��
o��'�]���S<���B����/3ǻ��bQ��~�,M$�ݺ�~����0P�zrG��٭@ 9-ՠ ���{���N��L0(s��o�nV!N�y� D��/#�C�������+Ľ4��[���7����Ex�ٮ���h����sȽE�X�/��Rv��WܥK��Fe�|Q��K��GTɯ	����)nȴ7m6�~J���FL�˄��o���`�9�K~9�tA3���8f7*.�s{_�[#�?C��6�~�6�G3���c�������w!M�����y�˺v��;t���L���<9,��P;j�Qx���c"��`Y��n�<w�7"�l9��{.v*B��9E6f�K5wm�
��V�-��D�����R��'�	6������Trb �$ᵉɍJq�o�׎� ��i�$X�
#�LD ,�#jX��
�i'&	�R3�:Tx �ܷ�s'��5t���q*&	�/11W9:a�r1(p9ժ[5�������u���y�4����c�m��K'���7�y���;3p��Uśm��x����iK%���l�Gu���Xt�T@�׼��x�_��x��ؕ�$������f�;��I�]{LW�c-��4�p箦i	�i���:�cܾ�,��RQ6s�v9K�����dm�u�ؼ{z��y� �5����[���Y����꥛�~�=��rmn�Ly[${WawU3ޚ��6H��vS�F��w���hq�y�����cX>L՜b�S�"�W��mԓ{����~�lD��p� u�s���Y�����@�k��k�$̕��+�{�iCPK�C{�N�5ñ#{��;3�ݔ���.Jz��r�:8�:��E��Gw�
Zn�0�{�Ƈ����2����K���Pu4F�ZH8s�.rBSh{ʽ~���H^c%j1��@�^̾�B�<+`�b��ѡ�`�,�
a��z��H�6�n�%���n���D�V���Ef9� �!E>pG2�-21������� ���\���5h��u�:Z��Z]A�����+P	��>�v��}�S��sG�Y��I4�n��q�԰-Q��Y	V��3��
�]@��a�&eШW�PwJ��T��t�}����b�����Y=�2�"j�)�	�/r�O��b�.@�by٧"���~1����g܊1��'��$iW��� {&�������mڪ�K @. E���;�Tn��;`��1/|����9Ue�#<5���	΄.cHW�[E�׻r_��������<��©��	���^� ���Y@_L� D@�����#�R��;|h�]���"�\>Y�����F�/�I��Q$RW�-�ZSE�d���r��~kv�I���*�V��ms�y>/m�TDz�<�F�Vnac+��;:h6��#��`��,EoyV�Kj��L���q۵�o* �1^���ܚ)I�.�" �1./9�ˏJՎ��ʛ]��7�_0�Ǭӫ��r��ݒ����e,�X+�ٞ���"xa��L��K�8��C^�V�ܫ��3�v e �$�2u�k��Nb�y�2|ё��\�d�)��Mi�Y� 6�z���m"�orU��v��C�0Qb�Y!�P�D���n�y��,��9�t��m���M#+"C�&�e�I.Z=�LY8�]�۲S���T앸���~�Sl�-��vZB��5��_sy�c�F����Y.���o����U���YT; b����cpf�}�{úǭ-��i�5�,��u�D�MY^�tlze6-��3��֗��pK+�ܹ�צ�;8|��ƢDDw�D^�|j��`�޵U�O
���w{�u��`�PgN=q0
_�Mx��Z�a�Ϧ�z�j�B�L	%��_���en�����#B���W��+,:�I���v�������α}�gKɆ�Q7�fs���p�,I�t4�Ǌ��i)��9P���|�r�� [�C�沧�	X� �#k���b��U��o��͵\,G��v�
�T��Tg�]����t�*z���2���k�
�&��ۋ��PG}{����Sܶ�ny���P�	� ,���""<`n�_���t��Gg0�����oYkh<��<�{yV�WD��=�.g{��Cx�
���=�v)�!´=��o��S�:�.F �oHdf�l�AH0`�� e(���|��aZ>��,��Z��s+��Hj������ 8A( ��0�!�P
 �bp��\��+�p���%���v�\��O/A���buA;�ٺ�,P��dR�]�n${WokJ��o��*$��Yz�x��=(��h������i�a'�J�z�s�p�â�������0��t�;S�K�1��s�z׈�����D@�U{&v�oC�N�G,DF'��4 �n�����f��S �q�b���x[����{ν���;�
��:��m�jr��;�-=�jP�$@����í�-<I����
ݸ��ݺ���c�q�c}��q�ު2�;�����gzzS�ua�6(�ޚ��J��r|���ew� -��TD�'�����'�����|bԔ��I��l~�v�7qh,I}q�K奎s�]��{�0+0�V3�i-�=��(x8�������$m$��n�o<�[���� �E���P^k�Q�d	�0~�ו��IN�8����z��t	�*iC3��-ԗ<?fj�"!���� ���ɳۋ�����xj'��X���p8+��V��R�H�/�¥ę]��P�vc�F��8�ǒi��cɗ��}�r�y]����k2�Kf��=L\"C(�H�I�(�+u�	�N�8���"V=l�kS�ل$�#�F�f��ɐ�����ۛ�.v���V�Dǧ�,vkCo��n1���3�qG��ѹ�MU\�`Ǫ0��u�� \D�#9��-Z�'׋� SjJ���9��r�������W_ca5� ��:ۖ7����w4X���HI�^B"k��T k��V�G;�v8j� 5@���I�w��̴�]��ք:�5�����=�]id�ç�k9׈�^�(^�b���uAx7��O��ed\0W��f��c��"�� �{^�qʽ��zA��Ҳ����	1(*#��yآ�`TB`E��@n��m��^i�����I�b_!�q�Î���ќ�� Dq� V�@�zU/Eu*����k?H����J�uƅF����"<khVi�5���0��xj�X�/��Eu���o~&��;�U��c��}�1#��$�<���g�HS���3�Ӡ�� �n~�w�Q�*�7��/;q�C��9�$�ff��Ub���!d>�Z��3:���0#�`º�ìYD�J�1��d��N�Ls@3C0�C� /��U^� �G��*dm#��\n��6��7rq�!�$ h Rā u��͛����4\�z���˹u�EVҙJN��A/`��n
[����|����6w'K0Rs���V�Ŭ��8�����i �V�ef'J�P4`��'�R�)YN8�. P��M���]Ҩ@� 1H��w�g8Dn�{�)]�hۏg|����|nr���~i��&߼�p0eo�3�d�L{s���g�������",��^1b��U��S�-1O�L�_���k�^,kgI�tY@\*���%�*\�F�x���DS�;�sG������\L�t�J�7,x��B�Y7  ��b�X����g��*��=V�ߚҎ��yy��:������\=��u�������yoH&�	�F/B�N�A�߮��ds~���W��X @����.V+����{�ANZ�f+�ɤ�����m�Oi��VV˂���h���8�6grg�Q��^�R$�b� l�����S
� "r E҈o��NTe�b���s��a9��A��Iؽ��S 5�\$+�euꝛ�[D{�D:ٙ��?y��Z=|����")W��PJm���b���橍Z���R�Pl�w�ޡZ�u����]`���1`VռI\���+sq�Q���9B��������U�[�T�hqČ�.�C��YѱyY���S��t�c�F*JKr�b���F_�o:P�h�G^o0.��X���4�O����?n���8ۦt�Z���4�-Vg,��+y�}5�D[Y�,�I�\��'yMӊ�������/�{�̨v���zD�h��7��S(��?�$~�A������xe\�S�@�.��V\��� ""�GU����ּd�7�C������׫�5�Mڊ!��1��2��ѹ������>�_���$���J��rGE('%��w+x��M>�;�?DD�҅y�G��8/q�]�/\�	���%�@m������S��Gth�-��b7V�&���m�u��V	Ϊ��QՕ\��}u���� 6XTǈxy�U^�8��)��$^s�&�7���/+v�Rb�̏i�Ǐ��R����?xy
6]q!�q�k
����H�-���� s��D��P�d�u]uW�>AmqG$9�t�Fd:f�Յ��=H�d�ia��cax�&-�NYB��.��<5�k�Z�+�=�:��[s��ӊv��a�W����3b��$h!f�۫�p��C�� f��Y�zӱ]	XhL�쥖�]��Ãy�nf��O��(�%����"���$��/�ʒ6,���Tr} @.^ԉ#��$��.�;qL��l߯{����P��:��W��ix���̥҃��MbѲ�F|y�s��̸��f�^x1VuH��r%.������������J5��!Kƫ1�~�{��8)(ebh��6�8��F�cQ��Ƭ�B���զ���A�O�J<��mq�2��V����q�i.�8z�N�s��f�Q���]h�̤2_Gٸ�HX���F���P� ߭�C<\ ��B��O�ݻ;\�� a�0�sw��"�P]ot��`�����|cr�d�(�Y���&���G�#n�w}^��ϗp��-�#�G{��\�G�
-[-�g�}���4�q�́ i	Gd��" S��:�ozS[j���1�W��	�_Uiަd-"���9�N�)B�p��k�{"Ƿ�g��j0�<u�$yoh��@C��t�A��PB��4���Ɗ���7r̞r�Tt*�\'k�d�<f���u������#Ug�솥Q�h-��5@���j����]�eւ���M܆A"h�EZ�����0L����We�
T�A ���K*Gh���N[��#������ZS�R,�T�n���������6��c`Y�&Ƙ0AeT�e����;R�@t�@�A"�t˹� �%s���(�J9�A�K&P �P1�$�5&IN\�PdCz]1��j��P�H$�f��D��GOwj�% �R�C�P;Y����_C�D&R���o��%�����nmРX۴sm�!�{[�`��z�j����Z�n��N`l�.ȤAgz�f�Mњ���m�;�Qɵ�f�Ԡ�^VWY$����β]�Һ ,ʰ�0Y�^Cj��}�^[������s�*
�%+5�a�8cņ���(7s%	�I0�72��h�t�/�G�dT&hr�[��@��Y/cC3I�P,��4#�/�.x��]�>Bj�p)[W�l�	�9j���y�����#
�6�J@�*�M4C�ȨJ�"���uP.�$�H��� A$B�W���'��9�+4j3N��u4>�!�w���C�	����h4y� &��&�6�>��M6�(i�d��$��'B0jh]�1g��{�:�"�eH���p�q���$�G��ۡ`�e�L������nc�l�N�����Ӽw��^�Y��(�!ΤIE"T���S���1Ojh��}EX��`�9z�G����~،5���*��Z<�_�7�������Lm�3���un�Y�Ik)�!뉜��Y���y���!C|�e�54k�
��Ыyl�z$Ԥ}�h/���h=@[���]f����z���)�!u�[J�e`2���8�eۀΑus�����l<!���:ܴcW�ogdT ٤�P�u5*(r��Wu׈�ռ#{�6�}p��̊�i�:�ͷ3�m&UXɼd��_b+��Iٳ=�}'U�坒�<���&'ò�X6�;��LV�dU�-��이{`�.lQ7眨��e�ë�T6�2F �!-��-�L�\����@gSO�on]IY���j��z�F�2WwWX��UҜ�0�YĘ����mZL5d�ɧ���o�]n�	c�F܏4(0U�6�J��҃9���νZĝ� �*�냱d�E5��\;����i��mw��֫;��)�Rp}Ȯ��r��z��U#��EI,��"�N3��j;�ge������g���[��ZW̼��i�-�]fC�*o��vkVW<Y�Ǹ�=!lʳp�26�"�Z5�b�y�{�1P	�U��
�[*t�AW]��R��2Wۅ��U��: �96Ħ���5�,�{�ѫw�bҨ�kV��x�q���3�|*�7{�Vb/���\ %a��)鬴(IwHZ����Z�oi��)r:M�*XʍE����v�^����]�c�E���<Lp�9�䧲��;�����*��]o�z� o���N�с;����ΫJ�gi[�;Qwu��捱���m��v'Ү\݉,��nq[w�9��SU����فD�#H)�@�!"�,�q�#�`2ՠ�H1e����@D�@b|� D���,��B ��3�Ƙ�yŃd �Z@/���7�����H+��0���0DD{D@�#�!&�`I@��rDp� Q��\�@Q�DIf�D}h``�r` ��Q��@�QG��0�Y�1`og�x�}[W�_>�|�5D�0�mDP0�(�I�ޘ���>0c�qh�1�(�`H?�b�� �!��`�1k�Ȏ1DC=���,ƃ�7�Da� "��@��ܰ#r�Y��r��C��G�@ @$G�3��3ɛ1�e��F �bM`#$a��5�T x���"4��&�|C"�ey��ȀH��!&K0��d�5�~���ovs�����r�@�2`h��B Y�ڈ8�Di�0�(�<5@)`q�1{y"(
"7��	0�g�!�d@$| I b $�`��@ � �$� � 	" ���Q�`i����"M F�,��Aw�^�\�P��� � I��c�& $<�] ,�&��Q�1�	d@&�N{��#��	qF�0�D]\����|�HdB1c-E��,�� a�5rk�iZV���Gϩ��A$�b(�0$�F0	H� " ~P$�4b�E���@�&8��+|�"� �>� �@�C �@����B#��@��������d`k�k�Z���7�k��@��fL�t�+P04�1fHG�q�oԈ�-@Q�@3 �>�̘���?�!��#��FH`"���0$��t��@dY�h� M�}�\���w'�o�$Q�F>KL	>r���D��Ř �� Z��f�" F!���"��4X� I�1j����j��i�c�ɘ�i�x�y�d LE�%�$I'+=���ʭNװ��<t�E���`�Ȃ@$
0���H�H*4�	 i�3��Y�b-� /&`��& F"Hv��*@
 ��(�@�D�M�PB<� 1��P���<���K�Q[�RU�*d�2i�c��Dd@�(!�<\��˟g�[�3���@��2���BҒk-":���49���ؕ���������r�U�;���k�6�L���*#9H^����P"�!���׷b4���R�/�f"L#�
0,��Y��ԀO��"���,���$��##EJ� �0�#�{;n�M=��04��DI@@�0�@v�cD,Q� �. d"(�%"};0#�x�D@���p�F,��׬�������	o�aDQ�&�L#�M`��� 0c�D�@fL@D@$q��$@&0я@���- q�!F!�����J"#�8��� �"9�}�6h�gbsB���f�d�1��0Ȋ # (y" -�#�
 I�!�n��!�,�H�BH�LQ חR@�H�> " 2#��p$��hC��/	�g{M6:�Ux2 (�!�H
0�dG� 'Ƙ�ס�YY����
 ]�t`@���x�I���6U$I�	� fߦ,�2 I@�d#��E�`(��9�y�~~�J M� �P�����Z�2F" !"��Q�DF�,����B�b0�fX��c�H �6D��f.���o�6�^z�x�� �\�Q�����#B0�#�2$��Վ"��2#�����C1�&T�<`qd00�@dB���b ���d� �8� ����р"}>�>ׯmta`Y��(�@$bC����" ��$2<A�F(8�ȁ��h� 0�& &ǔ ɤ#ڢLp��@F4�>ً1B1DA?0�x�1 ��ˈfL
 [6'+�]���@& $E�(���( :y� ��G�@�L@�f#" `n!<�QLe�D|`d�ޫ�`Q�Ŝ#�i� F�_�� 4������5���e����"1�6d���>j	�� a���� ��'L ���I��P(��@f1HY���,���F&~�P���0�|cLI��"=�> �B����@���*�w�4e�⌍r��g��!�=�s�-�1J�0��0  ��#�	$P����TԼ�]e�tަ
]��+���Z�K��ŬnA�[���cW��2��\C�@�R��@��`�1�����^ӆb	��m�wg�! ���� 4D~#�#Hh�">��,�0F���� �HD �$"4��2`Z@aDA  �!�GLz ��7x��(�A1d`2!*M\�u��>��_M�ݿ |�dQ��Q�v@���H #=���C�8�g�� H1���@v'$��w�#�$��2����@�8(�dQ��� I	
ks�x�J~���NE �@G�
�;0>#�LAx�#�b������	���� #Z� z� � Lr���H�O�Y�#AC t� z���Dx�c�ȹ�Ɛ��`Q���r�Dy�'Y��&|5⍡{�o�Ɛ��M�n�IH~���~�SIm4�kr�4�ܗ#�64@�o���F�J����[��jiþ�����!N{��6vOL����S�T��y:��hQp40�*e��mƩ�SGwp��ޡL�Mռ���#~_>��~o�]�;���n!k3/%N�U�*��8Ĵ��N1|�h���7Rfo3X�&W˫�� �+��i?f\��^�j�g�S<���Fc�/d�B��N]E����s����e��� �V<IϜr:=��2sPF��!�K�� �;����O��]t���nߺ�s	�b��U��_��p�b0��m�b��������۷y�-��5S�r�Ԯwq��l�%�����;zE� 䡴+T�%����Q��������MtK�^���mH&w+"qC4d��󱎥?L��I��{� �u�<4M�36X������� F8�@�8$C$��]���uņt4�֢n��2�Rgyv#Z�1r���:��*WG�}muH�(E�8V�8������uM��trsf�Hf�n)Nu�5�z��?JA�C�Ih��&߷l�΄���~筎��\�>��C�4c��r춻��%B�J��e<�zx���恙����秕z�7^�Y��z��� ��4r���ѹ͙1Eop��Dq��tEy��-������Dr�P���c�D澬�r^�1�Q�Y�e�ud笯���>ɺ�H�ƻ���4}��!���)e�ߦ�aR��tl���aj���W���5��Z<����T,>��Ƭ�7�~���f�<����MP �_��ȕUUO~;��{�[Ur�J0��W[\Y�}��-�3��ڢe� <�:�W]���4!�tc�\�_H���٬D���oV?����W3�B��v2�o���[cۗ'��K�e��S�� �D@�r�8̲Dߐ>����_�稏{jf�u3�1���FUC��L�wNN�B�gr�՞n�`/䇊�3<<�^������I�&\9��
_k'!�@gk�K/(��ʧ�^f�5TV)�eK��*�C	~��z�@�8f.�Dy*����u�Y5���x�R��=��Q�T���U��h;*UWl' ɓYZ���X:	T�y��0 ��%|�W.�b����������_a���n��ߨty[U[q�p�*�A
�ħ՛��Jk�w;��m�S������.�V� �U��^"�
���b�k,ʶjF�$��A�1��Y�ܵU�[�Ǜ��{�V��t���X��l�b""����X�#�_4�32�YR�,t���HI���i
���ޝyW�ڪ_�).2Oؗ`ױ�H\��P&��d��KV�sj�?*+n���OΧ��'�}5��C�K��d�/�_�L��lq��U��-kmj<�T�l�!ە�[�����WO����ܧ���l�.ň�{1n�3��8X-
d�Q)}�T��]��@ z~q^�� ���"�|$�1�M|��ݮ�#��{�"����5)�~.S���Ԣz�w-�wFC���06�ݜ�wL��s�w$�H�Z*��[��c񜧐�z���J=��s=� y�uG��d��)�pn܊Y����n84%�|ޟ$���9";�#m	�M��y��a�f������/���OQ���$����l*����S�R^F�߻�Ut�J�[аve� ^�r>��-{�%(��x�>M�f�]>�]�N�r�ƭ�V\�S�P���E��w�_z�H�g����I�O-+�'�
��؆.dA�5��i����Z�wު´;l�����1�@�LA�$ mD"��LA�$�U�l��%��$���|$�T���?k�<�������S�Z4�Ya� |`A1�`�����M)Z�e�ۡ�qS��.�Τ�WT���LΈ�P�&��33J���F'C�Sq*9ә]�^?�I/gE�I�.#��_e����ǨU�b�/45��]�AH�����6GSSr�jW�'�GD�1�v-�����@w����n���5�ֈ �H�1e�4�HX��y��zR�3Q�)��Ѫ�Ǐ��T�21C=`fҌ��ķ͛0VD��X��q����s��8��F�X�2�e4֮��%Ȧ����McQ�5�����/3���&�-�UB��؈ 6��A��ɹ P]��{�ޖ�G2�|�#b�l�3���Ҡy}�@O�=��{{�����ѺyW}A�H�y��o,�@����[�����u��$I@���_�3��@D@��y��
��i�O��9�	��rG?jo�HV3���W8�������#'Q�K�����u�<F���<jz�'�Ø�i����U;HM�bc�d��N[c���S�l5��D�4 ͷ��Y� ���������vB�{��_fʐ�*P��hy;ʶԣj��ҵW�i��s��F�>���?y�ҽE��Z�᧕J�"�:�K+�_L�ˣxx��L�fn/��p�tj`5�D�$l(`R�QS�^Ii�n�2�5�/ۙ~����Q���Cw.����%�=��T�9�O!� Mq(|�˹�֦��X&��oy�����,lx�l��A0˻�z^L鯴R˻��3�f���3;�A9Z��`"��Y 2!�f�*ܵ�\�Nk]��:y�飕�H�_oVMܪ9|:,k=�o#�����������D�.�j��}I�������k���#��Jw�8��ٕb���^?#�I���s��7��n��a)E;�{ޕ=����(:���_�ށ*�۵��{�%@7����< �abﲲ�5��X���R����[���3���3�
Q�hT�J�'�SRј��{��T ��kVM�L<ATЭ�e�i�~ff���Q�oP������o��[Y[c��Y��Y����ş�� 0����'�t�����������>�zjD��S��2�F�]��w�X�w鱬O淊cnߓ�n�I"w���d �hE>�$ܻ?X�ð���#/���kC��%���i�������B�0=����x�Չ�	�9��Z�\�0�~5B5Nb�8ijg^0�;�-~F�!G���T�ϋ�@v��{�!�FU<�z���<  
� 
�ˋo7�\D��<e�D���#/n�f7\�V�|�dB��ϗ�YD�ޱvAv��,h3��|&��0'��{�������ߍs\8����4=x2����K�ɛ��_=��_<n~>�s"�����<�!��ӡrQ�j��|��ۗe�o%�d�m9��h�,f�0�<��H��3u�o�G�@���Wr|�CX�^!Y>D%���gh 8�,�b�* H=6e����[��j�N�8�cb�N�w��K�A��*�Zz_o,���i�%���l�N��jL��`�.^�F4Kr�S��q �j��o�K[B"	���^g�D\�?y���/�u�ğ�G�WB�!}`z��;�-ke���0_ˉ�̈�8��'uԺJ���� ��.H>���/4�4��>V�V��:�����ţ���" � @���j�7� �z|��o镙�e��è�� ;�3B4fv���a�Bw��|<���U&�ԑ<��l=�����j��l��t��G�g��g�ϫ1���o�Φ��>7�DD,ڨ��cΨ��u����8��IQ/x4]/%��t�M�{��/w$�3�����9�n�;�$Cy�Moc��n�1��}1j��bw�ѹ�l��ř��
�'D׵>�f����)���'}�G��\�xßn����h}��עJ�Y�W�
,Gy߮� =�+��?�T	��~�OKͯM[�n5��s2r&Vv-�i�����0(����q��s�\" ����Έm����g�k��9s���4��e�]��.�^�:q�c_t��$ ,������e��ϫ��i�<��`��A/���[����/6dF���?��K|���I)����� i� �G��S-�O�	��N��@1�|a�ݩ(�ȴ�&�Gz��ƅf������cf�6��Wb��!Z4�۞�Yڞ��N�aL!=]:̬�r��Ern��5�/�Ocoy:G��\�Nw�}f�]�uu�#b�A�gV5�=���b��Q�$��$��Ia��J��~�=�%��8K��s�欸�}�Od��S�[��Vh�,���ؽ;�s�����ԃ�1 ��9DN1궼��S2^L���#��fv,D\�sPbc�v��5ѥn�����!���^%}�_j��GQ0����mP>s�WM̵�7T���DS [B�@Fw�7���h�|A�{����5�uC�1�o�O���>���"�|�P�k�>Ք��!��i���o;�n��BE��w>�V|h�V�oN��M�a�z����T�O  mՈ)���[�01�Fe��I���W[n���v$d62
+r�h�N�Ufb ��,�'���`]b�M��?(ڞj�/��D��g�a�g��LEܪq��*����~|D� �9GWe]ٚ7"��;`x�Mil7����M\���<b��s�j�s|�zt�`pS���z(��u!{�2�F�?ZM@���1�\|C�4�g��������p�?]�-u-׀@���ߛ��g�}��O��*�V5�ϝ�2���GSsT�-��tV;�yW�wZ6}�F���!ﰿ�[��=g	�?�w3�2��յ��̾!��ь`����Aa��(� �!A����]g�I��ρ�Y�����M��UN��v�,! _b0F� ��$�hAD
Ch!���!����	���&'�n��u%<��U�4q���S��n���}�Ї�_��2*/W6�s~ЫHz;�>n����ͮ�^zn����oX\�Z�0� 
�$���}wx�{����yDl�Tn5J����f�ى�c��]>�X7A����w�J��?����#u�t��]�g�y�9[�ז.P@�F�\� {��"6�ܩ�w�y�B�V��WT�DE�gԑ�1�D_������􊾍O�R�����/�xK��;�m߅Ľ�����W_�ו�4��݋�ΗS�b������3�\�I��v%���Y�}2~GɜA5U�S��Ue�KĹK3��� ��f}�J��u�bJ��&�>}So��D�ߓc>��>;�W�բ��循���]~k�y�'�6G�s
SG�d0g��MQ� z��+r��7>�i1�t�.��s����<�����G��hT�_�2�{M����)P�
�����t��e<��gƢ"�\k��H�gֺ<=WB����ҷ�9�w��� ����7�SV8|��TP��qV���(�8uSo��w�٨��~Bk{��ai������u�g��
��S8��Y�4����u���?
��T;3�fo6����>�}5AU��ݦ7M\��M����^�x�w����ܟ�O1�=���������I/>怟�S���xR���X1A1�dI	��ž~λEK�7O���*�<�4�pI�u б�3���l�D����9�C��U�8��|Q�T��}�t��+壛�j(��XBh��]N�pU$���A��	�n�85X���cMN��r��l^�-1��b��ӆ�E `y�+�J�i�l��;Tx�'�;Q
�_1%�5�u�0�(��4@�iS&H�FK5��tS�DEJ AH�a	Z�A��N�$��A
�޽�72�E0e�����wY������.�b�ޜ�A�ig�.烔<q���z��g�y�gr��vq�,h�q�ݺ����6�^C[��7+[���MV*��]ѹn�-2٧��ճF����*�j;�s�A�v�dҭ��x+7Í��
F��i�o�5/�rm���v�����ڹ��H������)	���7���j��\4���G�	6�̰�K�T&��Ws���G<�8���8Եs'>Z��m�d�G#F��Cp�K&�j����B����:�wPP�uE�%�Wl���h��ha�g�E;/.����$��&S���%n�@EQ?�Q����<�˨ 2�H�.�n݅
琖j8�x��ڼ34���*��� \�0�1�0�+ ��6��4���\O
�n'�cUp7P��Q����C0��i0獣�0�,O8+�&ݳ�9�0u"�ß9��
=y�j��~e`w י!�sѧ��w��y��ڌ�P�MX��Pr��6W)���r����f�:�*�%�׳�}%[\�ӹ�m��N�l�v=�Rs�inD&v��ā�XN��;U=�nZXC�7'T����+�U�Ӵ�f��\5�C"��-N�J����P�z�vr��h���Ñ�+?Mo���ή���F�am^�A�#��YhD�m6�_>e���[s�X���)Pf�V`�	�I�/�Ku����6+�;׮��Ʉ��w�{D�`Z�nX�m��M���]�@�W�W-����Sh�9��j��ܻ!N�����}�
G����t�s�Ր�R���������lˊVǑ;��molsy߯8�M0�� �f2T�s��6�z�|�Wd����&�6ܡJo-\�We�ӀG��w��Y\F%�MB���6j~W�`Y;pw*q�����rDf����P������iɻ;�z���]R��
5B��@~��ۼ�x�ٕf_G�Ne�3VÁ�W�����1��[��\,4G&H���h]��t�;q���}���ډe�0qz�#ue�:S��û4� �=��z��]��;ml�j�(�݈"��V��]��,&�݂���8���{�m�F��Km~<�ܻ�w1v,��J_N��'(�lZ,�k9D�MD�s��%�9��t�,B�f�bO��?�źN�Ҫ��_
��Sv�Y	�fv�[D5���Í� �&�� �ę�X7�+/;��+k�j���BS<��4��V *�l@E�R9��k�m�����;�eu��ed�}�:�*�Z��Uµv��H��M�$AɊlzD�p�f��j0;q{���g[=�}�SU�3@��kz��6�|����׭&����g�M�ue^iR��}�k�틯�\�7Om��j�Q7�� �>��5�
pݓq:��v � 9fo�cf��;=x��$.���ww�|rj���q_V������X" Q̌�<UW%8�Ir����M��x�^����_��m�rڠ7>M�9\�d�Y���*e�������f,��&f	��9'�&���;/����D6�w�V���R3`�/$���юK��M���a��?
����r���#������%^���1<�ƽmYk����>Izy��y�$/y���d��Sw�@=��uO�����	���T�y��-�u�֒
i4���'��������%>X�d�MV@j�*b25mKUD3��J�ٝ����To�T��x���ǔ�ծ��tdzh��Q������~q @�?Q8����4D��������U`8��q�٩҈�P��;'�^�E�S�(n��h���D^��8)JZ���0�ic����}1��]=V����� j�4&��� ���~�g���U�'� @�g�K��W~�o+�г~�½�0ҡ�t@�AP�C "	p��$ 0I$`�AC=���f���س�j+j���RU6[����8%�0$��N�E(CR$�A$	%�H$H��B �sL�ò��IV�Rq�����䗓��vk6���aȇ9:��ޮ}&͹��0rZy[W�o���e�CNJ���5,R�u�v7ǚ�s+0��n}7_�P9��d��;�0�q�v4�z!ۮ��AS�K6W&s�L����o�I�;{��[�h̯y�  �zn�Λ�$�y=9�Fz�9���ܞ/*��GaW�{[N���¥r�ϙo䲼�D��ba����)�hV��?}o��m�K�Y�^z�I�F�����9�W'� sNG�T��]-L�Ks�(�A����u�kՋ�G	�����~i�����nz��ʽ�C���6ׇn��D7>� V�^@,����!ʴ��m*�A%�eU��ܽ���<bX�=�}���A3�xb��5&���u\m�a������< a1�@�!tB���i�����rCO�u��D^ȗ�����s�j�5�T���4�cI�(�7��+�--��I ��C�HI0H@캺i'�K<��kr����6�iͥQp,��-Uk/k� ��|���W�he��
�~I��
�Hm}�BV˴�01=�����1d�E�˓y341��V ��Jϳ�wX ���Ab)o�H����!����*�w��n�a��m�r���w�Ϸ����b�t��P�' ��iK#��7���k�k�c�#>J�Ix�U�R@�?+�������o�#�i�%���"���$�L~�G��gA��K?l}��:�=�}w� O�^��j*����٣/�]�]�`�'KE���.i�`����n�D�Bqm�dxo�o�xv���꡴�}��q�r}��6���kfrg�+�Ź��{u A7HPs[�.\���}�k_Jlpzk��쨘^[#��.�v>GOž�Q�5����qu'�Sw�ؐ�7��ϛ�#�y�Ͼ��>E�D�� ݡ����F�}���H�&��Gy-��J�k�z���Pu5�^��Mqx��F��e_`��^GD@"7���JK�}w���C�zw�V������b��aA"	#�]�$���4�,��5������<5�}|�(Ҵ�Ξ�]�K%Q&׏�;˃���?W�jZϹ��V�4�w�4ۤ#F��Ҕ+��7{p{4�:���u���X�T|��" l��#���9nf��Wάu._�=�}��e�D֜Kr�H8 �;1 ���� ���{��"O��@ �ݷ}�}��{`�\����oXH��EE��)��3/���UeI4Q������fZ��ɑ�|�="j�<�mg�Fi�d}u���&���h�?-�Σ�;����|�sg��w�=/���q|S���_P���,�M_}�UnAx�h=�� E���Ɉ W�g��l��:;�%��l��0ό�����L�2=(��U$q/�h��Қ�2�z>�$���U��y�e@�	̴
 |@��r��>�����f�Maj_Wk��|�;�O*�D�-L�4���I	��0��:Xf�4?�S����Өm���{EvZ8��'p�p&Q�.��J|��ӹ��(��wr�)/VE��>��pû\x��u��VU������옙��ǅj'yѭ��A���RU�@�E�0��zr��ǒ�\77w��?��
B��Z��?%kX/����Ѫ"Xhڨt �]��w6>��z��_=����g;O]Irv�$=
&�y枭�N+�O/5i@�L�{lȿ�����y�$=��Ū%+K�d�� 3�B�2��eˋ�U*O�;"�)C��Q�r�Zq��FDm�����O����:���Vߥ��ΰ���=vl;��4+85�;ab�[�_����A�j��x�3`Ƕ������xyT����P�z8AY�+���f˘s��jg����׮q�̆�E�Wz��g4&kvL������׮zw5s�v����g�בV�)|]	֬s�^����.�<(_�x��2���T?L�:WN��Pb2������< DU�S�P��}7��W�F�g舏���Aיa����~d}Y<��'uoƽ�3_�V�@s����vsX�N�->�[��m��=3S���'ӟ?�� #`�f���5�}N���1� H) �A�� � ��� �H&"L)P14�*�����|o�8F��r��L��n�\���$�Apa@� 
(�$(��
�9�ԉ��:��\���B��hN�]���c���N���mK�G�8+��qS��G�ܕ8>K��������J{L=@�q��mC���XT���T��)dF��AUh���.�C��U�Ѧm�Ԗyw5�.�Og؛��yee|���k�Ρ�7�>��#��	u}�f;>}�a=�4.}�!�_��0Jv�ȣʨ]�n��g�c�e��0�ܔ�[#I�!�LA��{HV�ww̲�-	^&��uX������eB�@�5�����9^�m��
�T��|�8���Цo����h�U����LwvKѕ�ˁڮ��hW�O6��;�^&[x-��og#�\#����E��}%U~DK�����o:T[WBnt�]9�c����7n���.-6>�Z���������Ѯ�}k�2�J�S�XWtK�OZ�>{�9�I�u3�G�@���;���(��f\�Ғ�9�p�P:n2fDDV�*iɅ=�e�Z��~�4+��Iz�����[]�^j���{�)�(���$q�yr$Z�g�&"��`�̠.��2����Js�K}�ޗoK��F�Q�f������V���`!;�%������^�o�.�<K ow:��w3�zv�~'��@Q���M�&_��}�i�	�}o�)3��k��1�{��p4��B�`H3�w$T�o�!�Ѡ�n`1�ct����;�����ώV�@�����b|��N�m�N�5�]�;v	�7�}��]O����4 ��R4�8;�� }x�-��k����Y�p�T�B�H�#1
꾄�сo�4������a�Գ�%��jhha	��m�kJ�5[S���Fr�v�Ҭ�}�|2/V�͞5�h�i�����ٌ�%����|Gu��o��4���q_}^%���W�j*!���4�w~��)�(���fofH`N�g�	1�U!��M���H&,Ӆ� ���z��������v�B��p�3�I����fM�0~lS`,n�����۩�z#���.ᶀ���#����}�g� ��Χ��{L�˚X���
IvN��>�Uҽ��q���D@4	�ʟ �����uLH|T��@d@��L��bʗ�i|5T�D��O�E��ֲ֗�,�mi�w�oP�)����A?n���C�J��U�_��`�Ȉ�[�dY�7we�ӏ���"߸#��q �6�y����K�}���[9�=H��O��,��T�/�a�]g��^���r��U2j�I�4Ս�	*Q�cV��jB�U���Q.yXq�z�`���;�v�W�$�n ay���VV^S!N�����1��T��� c�0�]V�\��ז6������Z����8ɬmR���yO�>gg'���������\VOr�R�9�����#���=�1<һp7Æ_8�t�S}�>�|� V��-_U��~-^�c�^x�14�+�UDƨ��7;Z�z/l܂ȼ�նg������A �	0`Db$L A @&k�=?1�.�)>^Ŧ_�����\x� d+�c��w?�PWIU�����J-�`�GlҸ��i��U,!�d�L��}��C�nI �!=\(��j���ō�|َ�W�x摟�/��5>{���Ua�%��3����5�����~����&�����37>ߦXG\=�����4mK�o�?}�
�34L޴uR����Ðb��Q7�y��s]��|f�lڀ�+�(�KS@潮�O�kN|����^�ޙ��$�{����]�Ou�����+����2��=�8W���_����f��8cB�c�/Y�/�C&&q��ɗ��B��S�
n�5P�iG�m��n�w�"��GJά�������:|��+I�XϮ��A���[�!��z��-�S�{�%��u�=���,1�iؖ}'�x����@DcXk}׶�!H���J���E`����eG��d��(z�����]�#;E�"m�kN��&>U_����j�%��Ok���{�G6�t�\"�/"��w�d���m�\�a�I�T1��1���7�3�A�;خ�i7[�����Q��j	��Z�)u�E�vT�JL���JՎ�h����wsWJZ�.��x������ݹ��>���Z� /���M�+��X�@�?]��`�� �y� ^��*Ӽ�Wn����rϪf�
� e��ov�[:�Sj��~�ZL����x�DiL�k^9-��v���c�y��Di%�7
���^�����9�w��ݔaG���>M؇Z.����f��^�N4���"����ӆ+�`�Hi���P���� ���IWW�������)<P��h�VM�RB}qn�rt�F�t+�%������2�m�q`Xo�Tɼ�f]���z��S� U.�3z�ť����;�ge{Xs��M*� n����~x�1=m�����x���������a��{79�q��,�G>~�co�vt��ϩ�G=�&V��᮵⦔�DO[;�/GR�u�:Q��fƗ�w9Q�1�)45�-�F�F)`v**�;�׌Gh>X��zc��jt����������7����z{uNk��{�sWA���UF+�If Y������>�|3�c;6r��^0��_�Ƈ�y��r�În&2�Tq�Ս�@6=�)����2|�H��&�� e���>zfC����*N��e��p�F�� �P�noz�S�x�
��w��A.]��rW�	�mt�)�Ž��"j��̜T�O�m�;� �ݠ-��s��4΂��.���ZU��-�6��D?��C2�o�)�Wղ���B�ߦ��ODo37[�zh8��$>��È�o\3��5p�4"�¥lٙ��]�����/�Q/��;�X���]�[����W��]���Y�t/;R_:��B����D
��\�?|�B�ow��'�2�*�w�О�
�����Z��a�$�uFB�W�e��׳���7;�v(/G>C>d�|H�7��&�����4r��~��l �g��4+7�f>Һ�.y�Hy�w`��o�����G�4sf4�d`�\0}�FldQ&a��b�L3gf����ȯsE�����[�� EMKi��b����UF�r�5Fh,����fb���w��u5n���{�ؖ�Kηs��c�zO�}���d5�y����c��:T�^�V�!T��yç�`C�?W���vv�C�j{�dD�Y��{=��vh�93z3$�;�_P�=R�Rv��Y&�ܻ��1o�1�����M�T���E耣.�^�i׎5�\ Yw���S���;��zܜj�s.��������P�`�HA@,P�@"���_iψ�=y�T�ڽǣYͳ�4ղ�)����A�b�LJۈI��(p(�B ��P808J��6s��kbH�Ks�Cjۭ\�lޗ�c�H���p���Y��F��ڲ w�ʮ� ���m���]�vQKC�$�$o�����c�D��w�x}������z�>�7խ�_��b����U�s#0ʳv�4[Z�Ұ\�z�Wٻ�/��Pڹ�^�v��� �$�$	
��)-zw�PFs.e����)������	5�I�W�1�:͗�쿟݅Ͼ�X��
|T��ָ�t�wʉɓ�/�L��
�㋪b�O��֑�uo�s��L���߸��L�ת�.��l��N��Yz\1x�,�Hq�B&*X<*���D؞������wS��c���)<��%}h/{�A�� �u�Y���G~� )���{rT�D� �+\�흽��o*���Z�WN}jO|�It>�Uc�]�'Fġ�k�bP���$I�Ug��t]5��,�B�}]OSN#��FM�=��Hk�@�3K{^B_/�]��{���̙�h���z�I��i�vy��KR�v�7�%\�u{���5~W~w��u2�V�|ڔ̛u��K�(\ ��H�u�-�ٟUJV�Z� �I���c����γ�%���K �|rɾϑE�����K���Y���i���T�Q��vh͸ߋ�|m�����������_�E:��A^��~	�d��H7���ѷyA2�,�U�,��]Բؖ��$F��0wo2����A���"뵝E��7��;�Z�5������c�0+�ԙ�V�pڠ(
�$z��8�K�jwE���J]��X$�9W�(�8+a�A��2*�l@0"�)�I�'y��(�*�TP&�C�I�&ab��a0�gj�������׫5�J�zC�7�����gz���-c�rٙ� �!�K	�ЪW�d9��1v]^��d�;}i�sK�\��);닭��{1��e#��N�ē�%�5�-��h�d��c�sD�KY�Kr�X��������1�a�60n9�F�Q�8�hy;�E�R�޴��^о�*��Adӝ�h�a�9a��@ؒ +9ʕ�{��ŲV� �,r!J��ܻ*�zQ�j��T�^k���]"��2v���{ll��L50x�yb�b��.�'4:3���C��1�k�6�(��&/�l�=./M�6b[dZT��`�$��V�i����F�;+u3����C����if^�	��~�����񹣫�v36�MU� 7�@4ٳx�TZ��[�e�[�.�˽P�:�5N�u:q(F-4�uNu�m�y��}��M��N�A��yw!lSV�A�����bn-U�}�;���X��R#��Zb��7$}#m��p\��3T��8���g���^�
������P���^At4}F/Y��og@�hZ��N�H�\Lv�3*l�h�]����i#�rKΛe(�w�w��XS�.��X����3@x����Ɍ�������`VP�oqprwl����T\#N�v�uwz�aƧc��FT�1��z���ܓ��I�X�P7W�$�`�/��Ć=��X<;C�|��՜�Aە&�<�9A|�#��|�mH�s�=vTO��k+T΍n�K��q�m�����Q���ͧ9k]
�`�F!D�g�F�Sj���=�p��s+t��m���;�ݧ�u�t��)G(�HG�Y۠iڬt3��H�vSt$Qu�����A�.U�İбa[�8Ðu5�BLv�O"Wi+��@c����5�^�4ĳM���73Y�- ����:YwX����Z��D���q>��=BP?�8w��F:�9���H�����N���]����t�w�;b��V�]ugo
��NG_���n^��f�J��j���D�X&�^@�Xz�玈�k�x�(�)���E�V;C��\��	�n�,�Hjƍ#R�qt�����ͬ�1�ӷ��	.��ѻQ0K0���M�?�+���V����x�
�kd%�R��t݃V֍&��J7�k��Xޥ�m��s{���a�60�]��y�f�������g�E�y݄�{f�7Y�]-�ݘ�gf>�6j����}��O�T 8�¸���;w�T���啒Z}�r;����;N���f���w�;;����S_�͓�a�����W/�i��nɁ�膈�0�z�=���7uct߻�9��k�s�^����+���]���N�}���2�>F_\�g�2i��TPb2\D�`'�� `��B��#1R=J�zpz9�<ܝ�Rm�n��n�4$��C��8�;��qb6h�mW37�j�+2&u�R��o�v0�(�k�W�߇�z���T���yxY���vj��llyݓ�<�m��k�9��dV���F+�g�^�=��鏬v� ���"�y�w�����ժ�s���/����4q�9X���19zP��%�_2��V��lnٙ��2T �ḅgeS�5TrdݔjhT��Ύކ�����w�Ӊ�}���X���Ol���fy��t���l�}��6D)W��2d\֔Vf>�75)i.$vً/m��XB���y����
;��F���բ�)��U\D�!Xg#(e�<�H��Ojˊ���j�Z�)N�
�e"&/
�3 8.�����}T�?5�0�N�F;�C#4B��b�W�ߪ���Ҵ�_���L��  $�@x��ۦ}Nr~ś)1�i�m���ܜ2e ��$��4Sh �����E��\�H��6��k�YEF����ZW�C
��]������62Χ!JJTk"$uF��vV��/� m����}k�i��;�#�9�>Q8�����{�+i->y ^ܑ8z���@�f�}b���#��Z��N�*;:�!>�'�sD<^�I�T�����[,+�m�{�WJl4�)<�p���+������Lu{��g���f��%�S'�i�λtθ�Z�5�����t:ɼ�%�>�R*��ջ�?���.]�ʝ���|��#cSuɳ$(�y|�S�Z$����#|��I�
_��g��|�n��{���d
�V8n����wަ��j؁� ��D��.C��й�f��nWX�h����%������}�>�bn���>:���v<g8g�s�qt�;�����`H�+��Bg~����bn����׹4D?��ٗ�:��V6���U2~]Dn
zk����lU�@�����ɵk�D�I�8 c4�b�w��x�$&�Z��� �l�4�P(m�o�fB[�|umSov��w�����7�v��3�SR(Y�e�:���pc����}�2�ˣY��
��llVc�J������yKh�3O�\�~���/�9�;���x 8�Cw|�י��n�Ղ�)@�D�"�	5�f{�ύִh��#�-S��	���[�" @!�tol�u�έ�*�Xm���v�6&
�Ip�ͽ�+(�\����7��h<b9�ڔB�x������KX��&�ާ٢5��EB���}��h��DjT��9e!�i���>�=�9yR��5{V @c������V����0<���w�j�Nr{�Q��T�
��J�xwh����S���]�6��'��KS�J��L2�Ꞣ����7;�8n=Q<��nI�E5E�s�0�WX�Ϊd��'�pU]��KR�N���Y���ׇᥱ�
��Uf��Mz�5���w���A[r8���h�;�|5����Y���������F�M��hs~�W�J_i�&�OG(���&.��z���1�ً�z|*�w*"����T�.�`��4ܓ��rq)��{P�s�-�u̙���9�p5��>�# ��a�r7��b�[�C�ߙ�21Z����Ш�E�C#JSڸ����o��it}�4aX�+������w�m�ю�?��o`�+�C��A>-C�.�UH$��A��Y�>P�*�7/�<8���Z�͗��/J���o��:��ܝ�k����A�|ތ�F�l�yZ�������`
Ϲ��aB0� �@G@� 
e��w*�d�i²v��e��S��bfia���Da"���4h���S�MQ���ꑾGCG.=[�qs{�e#W�;�����5�����4v�B�7�fZ�Z�kf�!e��O���\��C���3�~'��3y���1�g$���zjH�ʝ})��i��ƻ�γg��{��P�'t�����+GrS�N�Y)������˫ 0���YE�9��C����4V�66��j���*Цf��:'���P�E�������OC���Wc��'�L�K3SN���٪������P|�5��/�剿��<:F�I����މb�}���Q�X&;o�4f\;��G��l�O�����E�DO��J�&���\�M�"e[�BM8m���cJ�ˉ�6�����21n�Q@o��ME<�NU��z��SUQ:sf֧����y;nܐ�Y�vn(��R-���we������t�0�&��&���
rz�=N�d}�9tUl>�;�(s�DlmoL	��Y�jT��m%[u��yM� 9RM���;��BF�`YW:j"�)��asüs��(���2�M�r�T*�˾�0�ю!���R܊���#�M�>ӥ=#�F�D>T u�{����Y�*i�Q (�1�f� IU܊���y�D2h�0���a���U�_h��x�|1G�򯹭���ԑ�5g_ I"�v�C�)*�Bb�u�
�X�qp��§&ݏ]��+�U�
V���@J�uڰ��f ��iT��B�+]�������]�b��ͷ�/���|%waT�����=�e��ƒm��``��CW4 \� ~�5ﻯ���O��o1��2h8�U^�V��9�f@K�у�_(3��3�-]o�]�st�&Rj�ǜO�}K^��^����2�{�F/I�9Xc���c����f�k�$�q��@��OW�ܢž�yh�~[���Anj�G�2!���-o������	z�dMr»y��r�H[���&1p��^�Z�UR��
���2["����1`p4"��p���u�:�n�<ڥ��vȍr9�[F�/һyq�#A�ɛ,i�,�}���cU䩫Xե	2��m���iwJU7���Zb�y�=���.��:J�U�EC�z��̻���=v2���!SuQsx�t{;�4�${.Y�=�]�h�|���g��}��y @�G+�g������zJ������%?ۈ��A
;U�gΦ�ݓ2i��wc�n������e�`�<)|~�P��������]W�G��  k*|���(P	�� "{&�6��#��mD�ƛ{�^�z�1��u��] �� ��V(E���l>���/�NVʝ@tv���>�EK��ب����e5Zp�m�G7�ՍK�ɧ��[ͬ�xy���s��<1k�i��yt�Ӄ�}V}_=eO`&{�߮~���/"��>�GX�c���x���$�ɱLN�x�\KDt��r� ��:����YKF2���O�U�eK&kﲪ��U9p�A?�K��*^�Vz��ܜ����Ga�m
/{���������K���`��U�ҥ���ԋ;����x���f �"D���>�7�����2���t�j�y�F9\o��べ�:��:�QR+x�x״�]�㞹�aZ�\ۚ�tS�|��˺ҵ߼��������nw��*LԱ��+��ܺŕn���V������*�����ϱ�/��.@&���q��e�ފ�}*e��Mhɷe\�D���]�yQUŨ�i��NG/(:����qD�`p�y\���pdɺ�؉k�v�k�����Y���%�뗽���Ǎ�����O#�gM/7@i�!�B���nw}�`ݗ,/�~�`�����^.{�ʇ���b�b'�T!^A>9�}pL�w��1f1&�Gj[��������G�4�T��kNP_b�V�����w:�Z�x��{�k&ɮ��#ٸ��?��7�>S�1���׃��x�=v��h�V�Ֆ�kՊ�;dW�����6ԡY��&��Osapst`CMmvѰ��==�;*�1ٔ`}K5��]b�l�M��B���*��I����LQ3|�Λ4�W΅�S^7�f�1��hݾ(�Xyv��۴O��jud�#��޸�T����3\o=�aP�(����j�	^uBΘ
�"'�w|�:֕�Lh�8� ��F @Ƨiք�K��������E@���K\V	��(g~g�F�w[��G7"C�VA�81)x��{8 B׽6.]��D��x�����|���)�=�kG��o�t	�:��=���+$�����e3�{���f�����O�s��i<�`4�jFn#�S�TS�j��Rb��B`�4���m
�b�����\� ;b�5Sy�3��)�^�(��ϸ.���H
3.b%�\��o�3�w�E#��u��:q���Y&��|O�W�$Ҳ�;��{T�����5���vtm��uwi#1��/t�3�����Tߝ�܇�7� G��L+߫�U�۶#OvS��۴6�/�m.�t��}�h:()��X�KH��_N��L{i��[W�<YWw&.�z��ם<r��7&�������j 2PU�"13��ʝI"����Y�5��gP� #	"jd��0-���ȏ9>��N 'A����|�hp��)D�i#$�h�v#rv���ۜ��D������iA��c�'��gLsj�'�/����3纘�;k�uvf�D�c.z�m����=p�u;*��A�i�ɟ7�;�8yqte{�L�[�k~���c��z��WW��cs)���t�aE�V�(v�뜾����� ���I�_�k����7����w��K��-��o�K�ߞ�G�M�	�u"[����Cke��둽:׳��q�-������ � Q%�_�~�1�;tq��Ε=2l9�El�eɓx�!�/�VK^<��M�o��U}e�v�ѯ���|�6�!hx�}��7SI�h� �����{���Hޛ���q���o8��A�c+W&�����~��=v+h�F���:p���*j�/�����.��(b���q3�~f� ^f'��rǞ|a�ҩsg��U>T�lN��nؒ�ťO�5��ҹk��޶��̈�vD�=�ͳ�`�(�8a����?4A�PGk�t��O�'-�ݦ��ZR�O3�$XD�	%$I"�$H� F�u⪝sݏ^ICۇ!�j(L�-+�<&C�$=VaT��{N������ޠC����H��a�{o�T}k�l���t�Ztռ��k+�2<�[��M�\~� f{�������lsr��r�j�o������)�;r/��T��:c�6��R�U�z�6�A�}�'��ܿ��7/K��Y�.W��9����2�V�Ӯ��w+K�ڴK�7{a
wit������[�W2��&z���[����cT�
��9��;-���f���z���:]Y������Fp]A2d�v��1���ӭ�9���}���޴�)����_�C�߸?o8�K9|���6V�O�X`D?n���3�ؓ٫�U�#Ŧm���yy�En���Ż����6OJ{�zn�z+I��4�O�>� w�Dx������vz���pL��tF�>��L���A�K�[�r�\s������pu���yހ��-�v�vul�lm�S#������U�\��pY�`i���v���� a���x�k����ؾ,Msd�6m�k���_�нlD���A Y �a	������r�\�U�g�eҗ<RAV"��x��}A�� �m�!P^�cv.����a�zݦ��FVi�֫�I��e�0��q�U�gD�M7��;��
�5ί�gVu�å&NS݅�Y~��ὢ�B����S3H����ٟ��kǫDͺ�`���۹���n���Ӌ");��3A<��E����^���T�Ab���K�I��k�1�����a�v�������f�*�q���DQʜ�W�F8S�lt�S��B�ā���ƀ�����g,�H��]oD�J�=9cS'�}\{Vk
�{��P�ғ��z�N��107����k�vc*�����6݂�T�)[:�����u�����z�Qx��C<BML�$�!����:۪�z7XB���۞}�g�jVf�����5���S'�=��lFd�$��sP����|�2l`�U4S<���&�+ܪfo`�t�٬]*�YK���_5ǯ���t@�yq�Rw��M7~M��=,�M��.�'M�3<L�P{�1�f���rZK�m�x{�s[�"gw\KQ�f�!��n4�+��y[�n�eMnS+Q�mIb�?ߠ]���5E�^X9II�Xeޙ<hH!�y��
x*#4m��Ս��82�\�l�B�+����´@�oZJ���]���I�)�jP�s2�!����bv���IA��]�f��r6I���8I�L����P¥L"i��� �`�ϋ$�M��ȼD=�j�4�z_c�;|7*Ԩ~txut$��ˤ՞����L=���o`�T��go���<�wL{6��n�l�l]_,Q�
fv���b��0����/��KY�{ �y3�%��ȕw�8�����H�b4VS�j&�32<�ѧ�VR�{8KkD9w��it�R��X����nT�N����G)�Lj4�f)�s0R<�S�i^m�B�MK@��c�q�/@����1k�,���2��г{��5YrR�+��y�l�^6�x9ыY��X��0 ƀ7��E��-��93nD��$��,�zB�n0��C �d��6��t�)J��U�d'��ҝ�miD���R��}t�R��#c
 �5P��Qܺv��V\���7�x�u�7!W`�IM�E����0*� �mZ��Q�ʵ9c3�U��Œ��K�DteL���J1��VKB�u����܎��}���hȽ����]u�]k��u��g�+��Ҷ`f�Y�Q��suZ��nu(�:�g?��'���o�}2k�9V!�����xʕͥC�Yoz� ]kp"�-� ��Ơ�]��(��iAn�Ҟ�E�p��^�͙��VѬΣGج�f<����F��}����g�p.�F[�ن� s�]��;u&�u����ƼY��
���,&���Z�i���Y���Y��,�+(&�RT�j,O/�p�G �GZ��m���!
�d�͛��ɠs\��{8�\��b��V 8�V��Z�+������ЃHFZ��44��Њ0�b�-'c[V�����כ�J��R��K�L_���#i��:�U�&ӣ>�s\��to�镼�D��s���mqw[:~	�%�܄-�+XEV�d6�!�c�� r�o&�[��|��^lwMvַ���v�NM����/g)B��o5ta��6����X�m;n.���S����QU��	���^�& ;7�EQ�-�؍�v��
�Xw��r(�D����hM8;!v�����U�zkC�qt܎���w�-��`؄l;�{F�'��y�'V��d��W��{���
�қT#�𭟹�c��'��kn�ko�qۖ��|�V���h�a��E��6�]�Ǻ��pC�=Vl�ׂQcr�t�D�r�n�A�-=i��^�
��5h�����j��uw��}�<[+^M\�!9;F���7d�.�A�}�BT�]�G�Ԕ�5-��`ww�u+���(T�hy�bRʰ�i�:����\��݇��sC�B������D�;�ݼJ��}��W�i:ԝ]�O��u�����,�W5�ח_+��I��3�A-��f(�aT:�FWN����P�5c�l���Zuѝx�eU�-�ñEF0:u��ҿji�W׬���7u�0�u�����م�8���&��sӾ�U~��<�"�{J9��e�8���4ld�m��v6,5e���K^;���R���5Է��sk�'|�����j�{|��t| 
���)���,�|]=w���FeQ�c���w��u�|���-��l��Z�S�p�Eb�}¶\.�}����oi��b^
�b����'�@��{�sr/5�nfV�e�~LR���:���F�ג��J1 ����zAh};w.����i�;��������y��o�I��|��>;]-~����i��.盘E7Z���&CC�Dj�^���K��폃0(�U}mI~�4�)�q9jq��:��!�nsU���`DX(*_���79a�V�j@��2���h�j���ɣRI�3����T����[��>���Ox.я��:_~�M���|�+k+�滀n�/J�g�N}��	�z���'��'\���3�)u+���L�4����&Z	�^]���|�_Yw��|ݠ����,r�O���e�s�M9��������6R7�aUR2%��S�^^a�:�"�O�����6�z��靶���y��&�5J��������m~��u�M=_5w�ψ�W�ez}���}�,f����'߳E��k��q����(9
3�sot?_=w{2oi����g�{��^8���fs����Ι�������:g������Nsl���[�:	;�ڥ�	��%P��>������!�ֻާ���ءzVb4F�YWP�J4�:���`�gdn����]l�v-������ȃ^er˨ '�.�u?gMo��5�s�[�L�eԧ6.�銛	͗E7�����3�@�;�j�CRs�W��s-;���K��-�c��S�[p�C"	��iP �;���M�w2-8/z����C�5{S{����[�P;i�uoc��[:�7v��ל���Z/*�Η�f�)��+�x�N�����Q��w�Gl�Ƒs�:�y��ƄXgU-�z^��9��d�؍q�f�$u%�#��~����}��ܡ>�s#+/|w���ulJOM8�y��u�֛��DQN�L���+������<ߧ�h�'���?�O����3\Fn���L���{�8b\��Ѥ�>~��ΩO��M;�*�~;�'����rZ����һ��q7Q�`��)6�.�2-��Í����.�Ѽ �7�`��MvP��|��l����$ @0{��9�~��=�H_.�O�SJC��
F�Y���^��ܞ���{�E�'�V+����
��a��2����4i����Ŗf��7�eb|RH��Rz}*�i���J�
�k@�lR1��%�k::7�n�*���s���x���c�P����EU��&SL��y��1�K��Ie���l�ܡ����u;ی_.b��|\#� h�
#qro�vf:�v����q�&.��wC�ʆB�+�x
C��	�õ����C��h�]1q�� �����Ju�޼y@ü�����-����ɚ���+���tچںÛ���������"�ukp5\׍�5�d&�>�8u��yJE�k�2��۵�t��{��l/�{ӈpO�uJӎ���W��xX#�n" Ue�C�K�c���i��R�lg���'��%��_v�'lUp����M��#��56_4�Q/[go�9]ML.#w��-[3q��%�й�Ic^7CF����ۼ#v��sN2}_�)�zF���m�����7e�u�L�k;���ھ#<a_��9�����r�T�3��Ά�Хkx딌=�,o��K�V�ݬم��D�;c�w {㵔��{�8��Ld��Yu����o��i�a�_��c��.׳�W�Y��F��1�D@�"b�ӇM^W�3�8UVU��H�y�l��� ����v���@)��1�i��T陵��
P���3 T��}DP��Xkp�pY<6�"d�F��Bv~����Pa�
��iM%s8;4V_mvO3�`��I��r���?�^�܌X!nt޾��G����x�Ph�s8F\s���4��ײ�meNY���NP�ww���:T�,O���7)���� 
3C��{��k�}�h�r�W<��avck�,�r���[!��/�w+%��q�HLS�ɛLvyi��g�תĩ��׽�MF��9��xW��;X.��i�\t��¯��m�YJ^��햭u������L���Ι;��μ )���d��3���}!D`AA������[����7�P�^�-'�4=+�]��sU��2�v(}ǘ�ԃmt�?%s݌t������� �LS���	˴w��	��rO:h���t�L�{��6q�s�]^{��ET�>���Ւ���^�Ga�n(�)��B�*���A�3�ӵ\K�l/��[��;�R�GT��A���:q����s�k�^
l�Ǉ@��/Nn2�႓{.�=j����S˵�'G�Fu�5���"��6���W�@Ů>1�� � :O��/�7���\�fv�a@�̹[��R�Nq��1$�"3D���Rۥ�\���̽Y!�'�lEd��}��3�9���}d�6��f�����%+`�Uq�Wy[�p�q�`�fc|��C��IET�e�$	-zlOT*���N�)��G�f���)F��=���G����d��ƈx�<���#l�xe����SKK�V�X�h�l��
���~_UG�G���b�x��tO����g�`'D {�����s;˃�~ΩY��/k��q|���l�K��V��U��ߤ����j�/��E���1_1x@����x�{������p��v0mM���l�O�=G=Jj��ۧ���y��C��I��}F�[��C�	�se�=�32hdp4:k��$s��	a"������ݛ���W0N`�+伕'���q�͆�fwR*Ǽ����\��MLt�ᱛf��k��"���%��H<��q*��o��gD-I�w���1[��*��8�h�-��?�m�3���B �)���A�0���%:a�q˩ǵ]*{���p�ݙ����ͪ�1�(�F�)Y���A_�d�M_JJU���U���6���g��ܹݺmL]1nN-Z��3;ki	��k�(o[[aH�X��dqa�(��%◟�u��E];��f�:��� k �C��RM��ͨ��h�+VV'�2jlZu��C���8�v��X�i>�1��z�wfwf��1:޿��>�&>ꓯ�{��v手k���	��=��I��^��(�����=$���5�_=����*e?����o���t��Dԗ��ͼ�o��q_�'���K
^�of���_�V���QR+�MN�m���!������{y;FhvZ̞g՜�#�S�/���]�js~�xn)%c"y�Cٹ}��#���}�{7&UMD-�AGRW���[Ӕ�f�43.� m�s���i�=���}B������W*w�2�ul���򗳅ž�����;M�\ö�ݙձeZn�L橝S'��j����q~o2���?̈́�7<�}l�dv?����x��g����?��߇/]�4W�cHf	���<��R��SC'J~[2�)�m��O]n��9��X;Ǻ �(%�ӳ9�AO��<.��d�ۣ�oC��/�+zleg���,gi�<3Ms�������w�v4ee�Jv�F��wW�i���l��n��0�;G���L��>��*�g=q3��2�.�iU!����4��ojW�.n���s��U����N)�R��,/LEI�X ��Z��y�ۮ�~�_��f'&9��ݰöγ��*ҥ�د]�@�Ԟ;l�X*�O
�F��yB��/N��ru�~��l�>��E�z����z�]V�3��df����ݲ�Ѵ�^��o07���3%rL�u��\�M�m�����x��	�ONN�g�!��0�����>���^�%`1�be��S�*.V��6ŉ�6}��<݀�l�fڸ�ghnu���\���c�+7e�<�ƶ�5���W_K����|��eH�L�s�nڳ���5��L�p�V�U+�G�H���7I<g�P4~��m�SV�F�*���:_h��d��U̬W�R6�+n�gGfGѸ�]��*�4 ��z��'��_�t��. `�%L �  ����2��DU��HF�b���7���8j��~��&�@I�pCRokx�5�'[ s��"Eg�N�`���t��u#.h;@��A,NZ�%�~5wk.�{��ΐvkm��[ˌ�Fs�A1L���.��ac���8?o�F�B�GW���t��oezC�& �L��z����yi��Sq�I��v�����lSR�w4B���[t��p`�Ot�"��s�P���!k$�{)||/�50��~��ǣvS��"Wv�˦�&7�!���/24�x.y�C�Y�ݺw\�V$�z���]����X�M�O�����"�NI�?y�,�w`|�ވ]{"4�������[���g����lT�:״�5���@~am;So'b�m�t��lϽ�U(�4�k{I����m�h��{� 2��`�Q}��n����[O���FvB���Ym䬎�{�E2}�ko���݇�`ٓw� 9�lF.�O�4���١��=L��Y���	�#0�w��1�_Eb�u�y��|eߔ*4m�m��yWw�Ϭ�Z�0:B��8���x:�#�KVW@��E)�1!�yl7��H������bQ�[�G5��Z�U�&����uv����t�����q9�C���u�g.�]����[���`��\������ɗ�in������E�YM�t�H�9�9om����A�:�ϔ�;�����ev�6ۊ{�R���b그���0���Ć��*�4��.����(�+� ��o�����rS����~m\˹�ӝea����wgT�9M{���3�����o�/��Xw�b'��ߣ�eh��
X��U8��c��0ǁR��x��X��DϬ �)�1�T�p��T>N���5��63^s�ϐ�����m&@wf_��Ua�K����o��Ɗ�DD|���{�_v��{��(��j9��Ꞅƛ���O ^��9~l3�ئg����[�GT?!�ZoB34�6	I;7�kSŁz�O�����`��G�����3M�/��*�!��W;]�<e���H'y�0]������ff����{zM�G7�6<�Y\i���Z�^��p{�8X-�d��֊{D�Pܫ|Љ6˫�:o9�b�X����M���F��b���]4��U���U��c(de�	�c��U��Ɂ��l�����!@a K5ÂD�,��T���*D�ݭ2��o��p��8/+ɰ�H
�/FY"���'zwy�WC�ِ��<0� �7;���Y*�1�|,�Ȓ�K%JI&¤�@0H�+R� kN�,��5��.�"�n�� X)�a����n� od��g��Sy6�a:5�hrCY�ͱQ�F���E]�8G����2���z��k0=Zw�U�B줚�w�G�ss�+|+m՗#��m�^��M+N�$x���T����#���[�v�rv��FR�Эpikd�������:���jl+�X9�.�����E��1��8�5%^R���q��F�]���!su����L��
q��܀ㄘnr�����+��:R��S۾T��Vl	j��%��q�@Z�Db)�,ڼ<�7ք2=�ĕ�X���y�gz	�O{�鐔���#P�Dt��pD���RC��A�` N�j����"�EF������Z3���]�.���j�r���cZ<�aU:Ѣ�wWuj�_p�ЪݪXf�E:ݔ���f-+u�Y��X�S�;�+�Z��F����$�I20�^v�a�8�GP�w׫Cݶ_p��i�:�0��s���	c!��޹`j��N�i#C�c��A[�7���E���*����I���ο�oUw�4���Сk�N�F��H�H{��XsѝǸ�K/��|M��V�0�IΦy�npwr���kef��\�΂�`���do;Op���\�e��X6%��"ط(�n��b���f���ԍ�~j��@17�ѳ�d��Ι|�JǼ��G����g{k��J� ���]�<d}Le��v˗\�=.�rsL�X�������yk��V�&^#�;N��2�[�RN���3����������2���+*p���J�E&;�����m������u ���^G��O4� I,u61*Q��w}�NP���6,�݇�Z��a*N�n�\y6�AU�_.����s�n������W�D����!Fr��>GNSǆ�ت��f���v�ׇ����Y|��/��3b�Oor�j�ʝ"�E�}x�n"�]�*���4��]`=��ܧZ������]v3G�����yԈ�]�ܺ]���w�p@����/�XKcuµ��o3�1c�B	� �����1)�	���	�n$��qVq�7�N���s��Y\�mjPCD~}��M�4U��kr_�z�fnz�}�xw���Vwo?��s�mGH�W��K:�q�c�F�\i��g���%�s����n���Y�vղ�D�$�q�b÷�&�Kz���ܫ�{6�T��ZH�	��� Ѹ�noPv��<ѻ���gK��E���L�NV]l�g�ɻf7�����f��i��tt�6����"��cZ�	Bh7l��R3�E��Z�h�1 ���Z���gM��+�(ܨ~��;?M���]X�3�n�o�I�	�y�΅I�3��{� EsS��:���"huJ�*�u�,ޕiZ/c����x���h�k5{($�1=^�ƺW��,���/t�7޹l�q��oLc������rыjcu�v�	�j��ݓ����Z����Ji��.��_��� ��]ӏ�`؛\z[����hKW;�=��}�-�P����@����7�����r������6��c�[�Z��&8
����ݛ�+�0@�lq��h�l�)ڬ���D)�u��j;y�� ���z�ˎvϯ��g�|~�!��b��^�n�d�LG9��/Y�+�QV򲞭̜���2�ｻ��B���[ĵ7��,ûj��n{jw�-���Or~Hr�Q@�>� z�g��@�@��z���b�g�u��$��O1=E`Z��V��WuY�����o
0��r8-��������滌��[t����"w/*���}.�.,:���l�d�᫲1�R�w����u��	mQ�9�*h *��hw������ÿJ���x��'ã*�o��n�szS�F]Uʖ����Lf:����6q}0LD)�����]ڭ�}k8����LNܹ����B�ݬ�~�N��m���lݽ�m��ǜ��ws����5{͔��)��M�)Իբk��@v'��V�-V,�>h7帏�' u��s�S�e��g	�3�������mwo /���oy����\e�p�~��kD;Mf�l��J�������;6F]�jn��}�q�K-�{�m��	�4�͕�����TO.�\��w>�z�0(�Xbf�rV���`s�ת�s��C�����u �U �z��7��\F��c��'+k6^%;Ե���LgV�.k27U��*Cp�D���dn׻Wf�_\��N`Z�_9g&8u��Z��t��? �$L��Q{>�u����Yn�O��ݥIMկFU�Dp"�wh(xg	� �Q��X��$�	mR�1d��n�`롭`z�R�;{W��m��|k�ZX��pb�}]ӸM�hC|H;�C�y��4f �	.Q��I�qZ97{Ks�u:<���L��z��u%��+p��R��Xk��=�R:�͍Q��[p�\B������:���z[^��]���9��[1�x��f06Cs�������=s�B~���)�����]��Y=�@=��]۶fc�L:��p"D�g3�۫��N�!ײGr,�W��Û���0g��8�7t�yw�������x�2�N/�F���].���_� }�-y�vS�w�d�^U��b�oy����l:�܀Pҫˡ`B��ˈ�W������^��Բ��HP��+@��D�\��r�%m��ޜ�G�gw/}��z��� �b �r�~�(:�'�K�m}�'Jtf����P�Q���u�e|3�{Zwy+w��	D4z%�a���g>O6U��5��fh���L����}*zS쩥<�q$Š	@� ��3� Д`"	$��J����x�չ ս�7�N�,��ո���fwl����`�D"��Q��A)�&PE@H��i)��=��<[{\�D8e쥸X��+@�}�!�[Xx�5:;ד���:څ�/o�o��Ӷ�DrW\�������O:bz��;�^��<~K����s̟#�������j�5o
vf�. u�em��35^������Qs�\��R�>�ݦc�b���绅7��u%	�4]_mb����&%F�`���Tƿ�꺺�|ε~v���%��^����u�͝}ө�\.��˧iT�Ќ����;�rh�>*�/��ҙ��+�}0�/xw��x��U���u
ګ؝׆�Qfи�u4�{2����G��Sk>���Nl���һc`�m)1�S�3�����#���N����T1��Gt[of�e��Z��$�������Zk!��w�U���͞�7a���5�1V0>t���DY�u�_�x�z��I���U�ǂ��ɞªx�
q���ƈ�
�������{�|���(R��a5��hUl�`�&*C8g`��vfpP���H�������ضx��q4����)��,V
8�]1�A0҈(�D�� ĤL�]n�T��mV��ӻQs��}���FK��q�}�K˘�����w5�18�qF�K���{74�U2�\�.*��-ߚS��yڮ�cU9u7��-����L�
����N~J$T���PȾf�fF�a�S;m���СM@J���duy��l��m j�[�k�����ݡ�6o)ҥ���|y;�[��Uâ��W*�j����~���QY�5j�t7c����j�W
�óv���J�v����@Ve��̔9��w���L.�;�� i��_xUd��Ů�}#5����7������'ѩ�ve+��]�\�-����&
����C�d��j=�}�
C"�֖�!�X�MS�/ol⬪�x<�u���O�l�����'2;�Q�PB��]�CP0����k=���μw�I������p�'�0���N���k+g�;�����]=��U�s���"�V�\ �pj���
޾��P�-�������ك�����ֺu�ͳ�f�8Y���]H�),���L�� D2�qd�BU;�:]�x]���3��[�ӭ�9��Xw�j���t����Hj�=�?�ڷ�y�β�Ӗǐ�y�_�C(F�*�����s������'��TQy��܎��.�{�;�E��[D�6L36۝�`�do�N��VO> ���9�qa�-�2:T�J�R]d�\��yu1���1Q��d�tC��Sy���>ot��wv���%�p��v��l��D�ua���.u�W_v	�~М�g,�>n�:Wz�B�#�g��e�g.ʩiތ�(�I[|�y���2���S����S䟧m~ܖgmϹӔwp,��?]y*�~��֩�5=�Z��MТ���W>�i�J�����K=���c �%le�p6i]�֟���R�r��hB��ӫt��U7���S(/�q�by�]j�{�X�""FX����@�tb �:g����<�v����P�!i`�%��5�m��F�&K^�����P����h��ϕt/O�Om��}U��Gǭ���?}\'���b\�"	��H# ��J ������]e�3&�o_
9I���vx��ђ�MIz�f""R``��� �nX�'u����F`{l]s7������Ԟ���&\�нx�Ms�-gv:����BT�'�ۗ��g4^��I��|��<��5�dI�;�!����ߟ%�ж���{D�Kr\��0~OL����t�]�`�{����W	CC�3���>��/��[7�a�Prg��N<��G�����p��4K�F���Q��L��t� �R��?h�ϴv>������������ ��(ڨ[0Q�/��s�D�r�S�`_#�g_[��n��&��U^��+�����ҥs���v��~�; u��E W������<L�U�y��a�)u**)�ݕ8G�l���/���Oؤ_xu;ȥ����^�jAwK�'�|���-K�o�<��[��i������~hj�*q�7)e�O��.�x�^�q}�����(�$�������*F��G�00%��ﾮ��c�ZSP���t7;)��hԲ%Wt�4�vs��[0ne~�Tm���k>�w�Uo>ܻ?	 �A$�1DD|`+�U��;Y�:��:Eʒ�����x����* i����`V&�>�(%����Z$�LnN��ٻ}�ˈͳ�ptc��ȮV7Ф�Mv������>�����,3�}NᲪ���;{�Yx�����
��/=�B̸�W�oǘ�]N:Jz�����K�Ǜ�"�V=*9op�->���e̷Q�P���7�w�2 " }G;�a��Qr���E�ʮ�g�6�c��9Y��#M�B�}*n�D<�
��B�nf���iR��#�T�i4k��1�ﶶͲ���s'}Խ�n.�[�]�3S�ׁB�^"I�tS�T�t��t��� _�T<D�]�L���z�|�$a3�����G[c>�?��?�ݍ$�r4�#a�g�`��2;սh�K��?���'�s����x	��r��D�x�'h��o{'�3��ՙ1��o0c�S��4b[�Yh�֕�A2j��~��-]��4-��Dnc���^�kW&���"1�)βvjs_v��Cm�f�}w�n��:�ʊ��w�x�&�����|�{��8C�ȢJ
�`LA�,��u�U���l�+Ưx�p����Iۉs����Gc�و��D �eFh| "M4�7b����ۖ	�!�T�Wf~�]ὛbR���!޹;�8k���a�s�Hi���t��;�'�2Zm>=�ݼzgw2GY8�1�]Jb0w�ńic�K�-=��fӀ#����;�'2�gg{��fl���=�)wf�u��MmU���ch�-�߄����Ǯ����z�����j	�H˾�[Ks�a�f����jt�C�_KO+�;�Q7ٴ�Amc��74�#��'W���KC�}�on��d�|�o;���~C��_vU��]�1w	.�z��͢�%��O��^�Q�1��n�^s�W""33�:�� Mz���3�/�WKW9?�E�Tu�DD�0�]&�Y�3�y��v_2^x����\���$�<����K��5��ԧL����m�6�3G>�[m��(�eA�=�^L�|��*�փ�yͶ�Ca_����p�Fz���ه\�y�~��n����y��Ŕ��F�>.���4]�ϳ/~��"�1� ޜ�~��3*M�8�t:'�w�Wr�J+�ݽC8��{:`�)\��摲�y^�\h�2�:������A���ja
��v��������W7tv��#����u������(8��6*�f���-q8T<J9�d���ѯm&ER��x�93���0@/]�6������:��>�2����Fmi���P2n��GNM�ͫkg�J��|�	�U���k	�"S��D���u������*��T��ڙ�!=�ěY��O>�`�nn.w��{{֧���j�������Nq��^G��L���w����]]��klv�}]��ߎ_7���y��y�}��G�M�:�}�`���M�#���ܭIʷ��7�.���&�Q ����8>���-NT���eJ2xZ�������h��-���˽��������~�3[h��z�W
�����cDD3 F_R�Z�����G�2��9м�;����{�8�u��F�*�Ν�.��7ۘ�ӓ"U7�<ͧ7���}�� eCȤF�;�Pt���ӳD(^�[l3r1�7h���f8 �Nm�.�k(�C)G��"��	�E>:�����g���1�P:r�� ��{V��]���WiS��qw�:�`��uu�U�Uŋl$�d��
LPֆbFSa��?�� �X�U��T�{ش� �����GV�]��;���j����w�Z�"����t��%g�\�ʶ�c���Lُ��(�5�=�-�i���њ���뤝��ĎӱvN�d���-��fr�ր�k��?رU�Z����]�՚2���N��o����S��=S{'5�.����Έۡe�ӱ(��n�Q���I,��&4u�)κ>F���t� eI߯3xw�k�r�7Ud�J|i��!�e:z��F,�ᆬd�jh4��p�P<4k��[gEV�B�L��P��S�*7�VFZ�`[�xj؉��$���p�a����g[�`OJ$��R�09	M�2ŗ	��իJ�d�ڹn��K!U��t�Y��4��!�L�m�+_<�u��Nؚ8v,��j{2d�p���I	��-?���"�Xm����<-"F���@�U���S#�I�2�B�d�n<(%Uv*M��`�9'ę���1
g+�ڷW��x����&���߯�����etS�}$��$��0)�aT��f��G-!����1�.�j/�`�I]=E��,+ۮ���`��Y��&�L�CAg=���[���x��++��q��f�CQ�i�)��s�"�tdd~���p���PC4]�\�R;[�X�V뤒�<<8�c(ŁJōG+�Z�{��>�aԞ��/*��Y�c��[���;�8a�]S�{�Z�ڴv~��&�#ZS�J�5{Q����`f)F�1�N���	���P�D�8�[�F�Vn��U���J}�n[�*�?K��2=�9ll}�Ir��]ڵ e�*KQ_ABm!���w�6�����绤�Vsy�#F�X'������n�k����W3�c.r�X{TOok7�I# ��vQ#�s& �C����C}-ECa@=��5�7S�8�W��z�S�5;(���߷eu��D:�%/��Qn��9�K����+{�WmW�c|��aEoVМ�l�I[����g4���7�)�2�Z3��\�-\���6����������{�r�d�H�M}��������=�#��۵HY;w��Q=��&��L��X�H��l�T�\x���������p �ԑ���#B�l���!��˹Q�mep�w1[��N�����+�4��N�HR�y�,�oz�I��q�V�b�/�@y&��C�2�·�_��r
�e�#w]\;RR�Z�HK�o��с�͋ꔃ�5f�CVo�9�^sIQƪ�X6���
�uu�/k@�� #۲����I՚��f���29g>�������a����oC�*��qۋ%0^!�� ���y��FuM͘��e�:"ɘN�x5�me¥�
i�d���?v�{D�ל�R�������H)r�����@�'F�;�X��M��~;^ܜ˘��{���@`��lMsr�Z�p+q5�Z�O� {sd$@o��}�D��+/����ׯSڶ3���d�;�*p3�.��>�������󓛵u_�:������t�sg�����2��9�Lˠ��s�����#6����Ӳ�t\��)��	Y���C���_/�^^�]�iZ�e>g�9�C��'�M��_�*�-�j��.�Q7�9�֝��^��0$g(FO����.�_��[�S$p��\o�׷{{%���ʶ'g�1x0�;�;��;�O��{�6��B�P�&��P�(Ժǿμ�*,�����$Ȼ�q]*��z�$�t� I�$ H�N���W˧dms���'7�pZ��q�H�턾�z��z�̘�SJ5j]`k#���ʋj7�B'gf�I�zZ�%�5�������R�i�����aL�iK��9��|��hi
�4v��=�y�foȻ6�=L�xQfN�ۃ�{>ئt�r�|X���o�{���޴E����s#��h��(+�1����������^F̸�V���յ�,��[��^���t#Kq�9������s4�l���ڞ����.._���е2kS��ي�Q�3_t�5�'r3}���391���}�[e�2ҡj@�������Q�4MKQ���.�zf^�� � !�����ֽ7B�g�SK����^�@������a�o-�[x�q�;t�M��,����T��[�T��/��Q�$�y��3y�ܛ#� ܗ%�h�c/����ұ{Z���
�}i�U��:��n�������ѿk��4�i�"P@�/�� D�"D�9yNf���L�����rS{9:�d�=҆ցF	`�H�0� ƃ�ah`�qC0�6
!\\�]3�v,.�ݽ���a� �J=�7L�!FݾY��R��(D�]�Pvu��}�Q����Ubt��z9����F���Q�ѮhO�*�����uF���B޻���3�&7'yUD	�I+��l5���O����џ.�4�����3�}FZ��n�^�\s��[_u��,G���ݽݦ�V��>�ښۈ���@���|��unQ��6W�_�Tn�w��C�L�f��c��gžn-��*����xvC踌Iƞ�Z�.I(q	R��6|.����ɞ�}�E"�h|���H�r|nACrBJ��?��lcB�v�0����w]�b�Vy��]A�z��5b\��3����Vٷ;a����3�VQ�8��p��Y�ճzڱ#�:x��0���,\���<��۱��g��ߪ�K}����_|�W>c�ϼ(�,|��y�(�
ff�"�_��3�=�q	�v�偛9r�xGۏw�M9=�|���֜�7��GddB��1�|�ޱ�Qe�Nf�{;r+Y���WR4�����&�8�a��A� �3��K7k�r�3�ʽ��-֌!J�or�Q�9�X�Sd�*Lvy��J�[�"�6�H��r{ս}Es\g��٭w]@<]����^t�ld�Ԇ[b�9�l*T+�q}w[�|�^��U�X��;��
 Dv�(�8��Quٻx��V��k\��V]�\y��
����/-oj�{PJ��[Ϲ��3�*���^�������o
~.���v͏��=2{�W\�'�����.>��n�Yc�o)�9Cnֳ�k��7|{{E�> Do�F��M_��;�Z�#�阇�O�4&2�n��B�M���w���>�D���짡�C'�U|@v��q�H����M�a��du��ھ�x�u�C�Fݪ����.���A�S+ys˹<V��(��8Ov���ص�h�Ӕ}���@�W���\�*��S`��;n�c]�T�ޗ�3J*I'j����dS���[�d��]���GC�x�.����_�nF�N^��f �IT+,>�݋q�����r�Cvs�ʰ�������ݚ�T�ά��T� c���pÒ�0)�N媕�ܨn�)r>J�h>p�=���04r���	�Vܞk�3C͊5����y>|�.����-�徫.������Y�C���kQ�oM�	g���G�g��D��|׹�n��f�L34���n�n�QJ���*Oq�]j�j�g�uެ����s�Y9Oj���t�W�*v+�\��U���U�����40���F�Z��<��lU��bZj�����h�
�f�_nxm@�w��B3C�Ba+�4op�!�(۫C���.{hf��ߡ!��׳}�J�}�ڴ��͑�:�%G5�Խ��;��Qݡ=DΚ}�z��W�kr��}�z�# o)�� �״�����7�|�{w�@��upl�Sa��<�ԛ��M�{x����A=lcؿ(a�nq���4�cD����Ÿ��Y�K?}o�,�қ�<����َ�y���\y�n����ܮ��m1U�t�a�»���iQ	�5�N����A�A,,H1Cd��`� ��P>�����mZF^M�v^��tl�R֛y�\N\���F���&#R���C$�	 �7A�TJD~�AH-ud���n�һoU���,�G
��j���OL���Jdv�[�y`T�3ktI8�`�_.r�s�3��P���ٚ�}T��}p�׺���Y�
��(�Z�]�[�I�n�nu1���4ZsN�ќq���g�������-�k¿W��)�ڗO;dK�MR���O�O�ޛ�x��X���:<u���*n�m�e2<B<*`��u�MB����6܃fQ�f]V�4�J�SQb��"J.8Fr�{Ʃpri�3o�g[ӛc��.����y�>�o
&��ʑ�Ɩ��N,��C1g���i�;���Y�DĵsS�4�uQuM����u2L�ʦ�4/"�x9�f{s3�>����^��-� Da��L@Y�ڬ���3����@���o��Z���k�䷉�_�������ޯn�gĶ��*�j�5�*s�	��r�qPY~�����T˹�sRpp�z�N��v]�qe�����_v|#�f ���1id�!�k3�uݔ��ʼ�n�D� a�	�4��8��d^fFo.�%���=8t����o`�ε���':к㿻c���]�8�9�Owm�+]�gonx^SF�M���:�\�i�(bϋ����k�;�X��Y<]���U�6�ם�M{�-�>�U5z�����n8;�_>�MSCv�c�3Ų�[QC���\P��uu�Z�dS�������n�����gN`"��@��zF�����7��Cz��4|N���1t��E)Y����;��>��:�9�_�s�e�ݼ�7�����Ʊ���n���ɺs�k	l�kM<��[&'s{^���{`fct��!(�5�4��E�.���9�Z�_��`-p������|�t)d;���M.�>\]�Q�?��iF}&�qD��x��H��Y����­b����T�v�l���G63ozI���R�uArǙ�z��i�L(��9;i�[�L���S�D��E>"��ls��oy�;7�s�EV?	��P떊�NB!��ndn�`�Af" @1�|�[�n9+^*{^�=Ӌ�n�BXHЙ-M-�"e�������$<Ch� �TI�@�e��"�g��ͬjA����۩DF�g[��	����XRM�׸��x��D�%D�z���dkf��)VU�2�<�Yk<�젇���{�]�����=�]��m8㏲&J�ަ�xJr��ri�mz��e[�U�X-� ����{��1�)����OpQ�%��X�VL^���G�uN���2>/�뗃��a�A`�bD�:�nj3|�":q�f[�ry R�������1���n$���c�]:����ouXk]oJyv�U;�j��y���W�M��H�uO@��Y�`sl�x���s.)�C)�Ա"�� ��<�Ռ*���{����AJ֓��2�Й�=L�@���#�}�u����4��Of�p���T�󴧃�.��	`�������MR'�k%�Ѹ�y��-)��S��}��'��QC�k��^�Gf(zH����s�k�\:2�@!S�}�<���tZ�'�?��x���(Bi\T@�&2`~B�Q�'5�.�V�5�����LKL�n1 � a�aDA���1N�dS͂2�Tf�DD/v��(,�ۇkS�Y������w45�Z'7��[{��3�%�:���Ù:�ƚ�j������͝??Y��SW*U�n������D��";8�_۝�<���k������e��iڝ���H��5�3�������<�v�[-�o'fg,m-٪7��us�k�s�/�W�B?�G7�t[�u��?)�6�o����R������bZw	�lU]>�{VO*�L
��0�l���K%��*�D�mg#�]����pg�j���U���s�X̪�����(d����S�j1�=�ut�l�:oK��b����Zm�)G(�2�T��T�aunc8����^��
���{Ƽ���� ���=�!R�5�.��g�&栺0���7}�;������[��#�1��i���zމ&�{Q�ٙ�y���d����x�bc���k�g��M�їL�;�k>�-��s����u�+ ��+e�fiP��j雷'݂r[�I�c�� ̢�=*���t�	x��\�]���m�-�-k/�Sr�T�^\%��w@�V�����<�������Cꃹr;;q�5*�9FFwk��̰�xV�N��Ml"��h��Jo�u�}�,\����f;��q5?V}��ϸ�gO[�+�ϗZޗ,󾾹3:��Xǌ�ȫ��۽�Ϥ]{+�^.�{�>T�yЕ�/��~`�W�n���1�cԼ@=���l��V����~kf���ɯ/o]|�?�;�v�Z��e���?�(E���[��%x3,�u3*+��w�ٜG��+��h++XցϷ��/T$���{iY�'?o._{�,��ժ:c*��������������B$��Tc~�Mj�V��w��kz��WW�E�K[8XP��Y [=�QM|��1Sxv&�O�����5��^��&D?�Vu�ܼ�,�w�+iqݔ��T��ˎ9+����&8���8�*=���w|��;�X�ϻ�7�;�`y|���:�W�~s߼��M��M���Z��,vh��6eN��aL��ֈd�ѱb�SBw;�p�7@p��pr�5v�r���P���QTg$��W�;"@Lͱ�����_Q���)@���Z$q/�ڲ--�y�!6Z�r��cVI�t�
}]��0��eV�l��6i�D�$���hBع��KQ@��@"���12�@��L���-&µ"s/��uvZ;I')K�C�}�k���V;:ؾ��K'��b�(���p�9M]�і�k\�M���<|ou��x�h�qG�p����+��9z��Z��,$8L��:�ov~59�8&f+�9�z�Lt��O^ܾ�ZI�[#o35\��tK^^i�x#�\t;$�c�YC
��j��/��]]G1%���Y����[�/��E5����I���u����疳���\{h�b`�i�,5&���-�gp�.��`�xH�D��@�A9F�H�:MSwX�0Ѐ���ê��]�&$+P#
}�q�<� QU))0�j�� �l���[�	��F��͚/M�*ٽ�����6l*;#'[4Mp���.�3N��	fp���Q����[�U($� ƤA�
�����9�%u��b���fK�2���$BcZg
g��v��V�����\��ы�*��P)9uM�hvn�P�oWZ��t���s��L��ьG�U�Y7�>���rJx����	�Gw ����=-��'~�+8&�i�zͨu�;�\��zp]q ��x��{�|�2�7�3i�+5�o��������ĸ1}����Q�&'� ���3�����e��qR���B��3�WNhji 
�1���Q�8�N]m
�j�6Z]���c���۱Y:�=O��v�0ԗH1��dr�
wK�T��J��:��y]�C��YKѫ�����Z�z;@(�3���3��ntu^��s��o-��i1FYwn���E�9W&��e�
���w.�P��x��坛]R���S�[��L�\�;�N��Ȉ�Ix@`���`���NW�*�DT��9��C�y�n�85E�\��6�h�Ƞ�ޭ|�{�M���a�%V렯�N��/x�䕎�͊�>U�s%*� @"�;H`���K�ۻ�E���1#:�eH�i� 
�>&d���u�FCJ]Etj�U�0�()�_0����8�؛T�~cz�m�V��.7���{v�u�v���#J����Y��Q����n�fښY�i#�����b�L_�H��}@�AJv�}֝��B���n�աk/6�؁���<��͍3(7�򴆗r�@t��AM�V1�Ք�����Pz�c�t�i�z/���;����.8�'�_I.ya��R�ns��V���;m>�N$��\���X�KI��Eg6N�|��[-Y����t&sV���-Z�-d��>�:j�q���;�T�ǲ�^�ǤE���@�KF8�Ø��L���	��P��*�ї����[fSܡ�]/3ؓ|�*����ϫP�ng��s�jd=)����Ԟֳ�6t�C���Y�:��>��o�:��I�Q��b]���	XX�kIj7��v78U���{Lp��=�{r)D �DG���W�m��~���d�mڗ��޶̞�z�����水�:ɉ�h�0�����όE�a�b ��0�{�s�;�o'2�q��<��33)����V�64��iS�J�;�a60݈���[�v��l��sE�q�a���o*�cTN�S��������6/�U�4�J�u{�����p�P;	��,�h�o%��oN�*\
:���T�6N1����5"�k��\�}%A���Q�|��{��}���2k����v��}��բ���3�]I���o��$ i@��94v�ͮ�5k��;MD~��b�Cڍ��0�~˧t��UAUo��G��ح{�N|�=�2�%YT��o���q��I�P�Jĥv8��Jr_��z2���U��&w���v�H�Fॼ�X��>��%����[G���3����S���gh��l����������4�yY=���|��������a�k��>��@�<M��B�\�V_�{�5ݧ�GlJ�ӻͧF�_�։��b6*�Ϧކ��Jjĝ��Ly�M�ӊ��_>s��҇Nݿyß���������z*���ڮ��6N;����4ы�����lW����BuzX�Uf�ҩk-�)Ĩ�֌�}X%ڝ��}�����`'�(�x�����J��x G�@��j~���J3O��,��dy�B�������b~�*1�r����S��6��㱦���3�����͎�b�a:�e���TȦxZ�'Q���n��)�t�E����}_�͝�R$]����@�� ��������>:�'��\����z,��#w0qF]l�,����wg�;�D!�H$�P|�����v��V�Ӓ������n���p�(�`2	`K8�N�%�J�ӑ/(��q%ͺ�[�����5S��`�#wY�:��m��A��F��bR�fͫC��ݚ�	�Օ㛱��i��$]Y���7#o�q}��\�����V�*IdM��0S����L��7�3ف�|��"���W�v��ŨX9'k9'��o]��a�����{q���WH쉩I��!�O�]�F����w����@
��� @>�̙1�@�ۚ�vӈ�zqe/XoZ����uB�?-�W0)p�չS�� �#n�4s<2��;��}��'U5����N���.�G����x�jTL��w<�a<�+�-�q��Gsn�v��i�������͂;��A_g�&��*������S�Ǿ���9�ߨl����:�Yg�C=���j��L�T��.��q�H61��o`��;��:��i�*L����������S���c`�&B�N��Ȍ��=�	����t���p�y�]M����0�9�y�����m� ��q��K[�L�z�]A�o���ꥊ*��>�(G�k����0��گ�
�v��������q-冦�٫"����Ƶe�֖T�n%��vӻ�h�q��yVslw2v�&^��s����Zj����ߪ�>��x}���>����^��,Ƶ]�$�~|������:��uxSN*�e<�Wh6�ǩ�1
i���-�T!��CC���^@�v�0�u���=E�\��1�۫U�]J��t�`��ܽOw�����Tb�բVJ���f��us����AbB��sU]��CΗSe1��gd��7esmY,�+��CT�mO���a��TT���O�/Z�]��3����f#F�Q�(�QB�f�����qxH�3�X�K�T��]�_u�_����4��P�h[��*r2�^Q�6�ᬶ0�K�����˩�{�>��|~׫���\{�s�\�4H��-��QS����2�1������:���5|ܩ�e�^$K_�K"i[�K���0j��8\�h����������_��~��\� ����V9x6�}�L͕��z�;��dӷ�FҒRDq������T3*�u_d���Cr��NJ�=���3�}�m�h���mo-Wݚ����- 0�1���-��-�8�Z�|��9�;,\@�o�L�箠�&��uT]]m��ɖ����q��� NS�Ģ%��
��Y;U��Cj+vXSQ�;��_�������� >LOfjv�;35f�]��
��Sn��٧���m_��ö���#���Y�6�v��_MQ��<���[[խ=�����~^���ξI�]�f������y�/}�d�ºY��٩�v��N*�E�b��fK�N��ټä^���4�pN��s��X"�J�eS�M8�W3���voq�b�E���{�ײ�H�w�O��S�U�f��k�Rϴ<���i)e�!I3wK��c���>(�R�z-�L���#`#��d�}���1 �_oov�?uĵ0��e�J[pf�q:�+�*����zw:��~被����C���û֓ܞ׿EЀ%�Cr�Ǿ��?X��H4a���Y� o�h��G����{��7.�`29D9l�y�� ��PSf�*��˓5��EX�K4i�p�Ү�ڎ%�qks�ʐ���%�g�}B.�N�/�����6¾\(�]:1���奾㜾�'����<��(,��3�B�+Wi�G�[��k��i��ܞj�]Y�]6��f�9�8fr����z��D�z��I��b��F�ι�T.TD�8���@����l;����[wTw3w����h�^$惥eX�ECL@�;[VEJdR&/Cv���WoN	�}��(���B)�j�j~��Z᭵4_Ik���A2=��^�5S^�#�d���p���V1ڢ"��Y�9�x��i���A�����3s����[�/��
�_<��s���Jr����+,�z�D���n'����в�t�'�����>�>�3�ٝ?C��^ʭ���_>��G9�ͳ��N�`D\���Y%W}�X���Z"�2��<��k7�)�c[,���~�h��ۗ��.��)�1��caAk�}wCԈ���ݶ�b����qU��Q���#D�֋M:"�����2ʡ���`��q7{-7x�&��o0��U��nt�ngX��-��g���{+�l��Daj�+Q7���(����V>�雎;K������g�;al��u�*�*�L�*v�� ��������V�l�ʝ�C�F��,툑w|�k^��<� �T�0 �"	s[�޾=u<��ێ�p��&mt�/sP
k..��`m$�.;���;�_����l�vnz���G��wa���~]$�D@>��5G'/Z����W��� o~��މг���pe��2Ӑ��Ҟ/usb�C&@87��������5��u���:��5�&�;�'�ч�H~ܮ`���OoMC���f��;oz�xľT���mx�;���s�᧰I�QSR��zy��|�����	6����٦I����;z�w��&&˞�MJ\'[����k����;�:�5P)����u�5�b��������7���ѱ�Z�� 2d8D ��JHJ쯸�DS�B�u'}�:�L-y���AC�����mUP�� ��H(� �`� 2 �b@�4�{�%Ov��Y<��3'�ͷ�<pZ�ts�
�gr�|˔gsG]�	�*�q2����Kgl+o��F�v�]�q�[�>�1^��2+.�ѩ����c�U5�S{Y�?���e��e]�yy��ܠ��x=�7>��^'�-�#{2}�/p~~�)-�Y��&�uZ���NZ�]Y�yq���_B�Q�Y�iG�����?c�=W{��mW���>�F�zP
����f�5�����U2ё�:;�T�/�A6dD�DX��7;l`[��׻-���[���ݓo8Q˧�o���
4�b��cvi���~٩=���q�=e� H�B����t�����}=�߯U�|���V`� 
1��N��=��==� 8Dɐ
��i���SD�,�FVc���NMg�����>�~1P�ǐ�(��\�ͮ�6��gG=�KZk�/&o�'(ΧcH���'h��5�r��=1��o�<����p���y�罢��cx�����`�k�ܭ�Wf�*hù��Dk���
;�������[�� x 6>B�D w�e���X~X��j=�1m=�Y��N�`�#� 	<b��MR��ə�r�˷��);D�~�V����t�p��-�	Δu{�ƵvZ�z۫�@����/����4�B[�ۮj��Յ�V�,i^�Υn�q_}�6�z��#�<J��<����4�jн�W��"1hzN�UU�`��wV<B�Y{��i�q;Y��37���F��*���_U̸��ς��1O\�rþsEH�
��v�L{^m[8-�[#����"�5�9��h�tnB��\��[����O V�v��K�a���k뢲k��#؀O�^�f�ͥ���u��Y�ax+�Ug�|���C�欯�{�)}G`nF��-��Z���L�v\gJ7�5�l�M���{t��9�%ʅ0�Տ@K>�3����-p�/��՗5\?HL�{�]V�k���+j�b��D晶Jؙ������޺�_�x2��TK�pvr5�XivH>Ȼ�)ܐ~�-�,�s������?v��6*h��q����n��aw��f�aϱ���m�3��3i����oyu��37��z�8���9��R��0j�\`�	�H�|�Ma�z�,�a�|P�jm�#��]�h��J[oo4�r0�E���W�vT�*�_R�N�T��N�"�T�3�tV�łN-��U*�t��d�uW~�)e�q�2�����m��{�;���X����x���
Fg�����ʌu�:���N> 0�"7�4��1�7j���p��͗ՖM��/靯c��=��b�F��3+�[�uL�S��j!��w�H���#2)�>����7�Ena��n���l�qRy���W�r���G����n����v���IW*A��`tH:��MC�úw�'�̠�]�w}"�������o'�,�� ��O�]���{��� C�g��G�_�:%rMs��r�M�y
��|ߺ�p�������[	�M��?���[�{�{�x�hxi�F��{�3���Go�M����4|!��s���)n��a���󽸚��`���Pu|6��xf�K�d�㣿�-��I1����#4n����;κ��F�-q�:�RhM�o-�B�����8�ȳ��d����;�|S�/Y� VX��7Gu�f<tK�t����{���)l���d罝v����X�ca�ww._S+�es!�����;����צ�T��C*�^�� ��7^=�.��箎��}�X�`Q~�����Vy�=N�Kk�r��@�Fʭ�H��V.C$���}t�+H=Ի���C:U�;X;"��*��_�SZ�CNͮy+�w6��4H&"�Z(S�w\�U�ݗ,hNg��;"YSVL��@'V��$�q,�M�)�	L�Tԓs�P̜5h�#f��Xj�E��	|�e(S�0�kFPX%�LZd8�̨RE!Gi�y��@�, �E�E]n֊��R�dU ޫ±����%��ִJŌhoKބq{�6vN�}:��er�/3��D+4�u;{Z���Kn=�yXA �w
Vֵ�NP��ɩL�tݼ�{��ܩWJ��*����Q�&�1�'9�\�������	b�^�.z�n�35Y{Gt�V�[�3m����s�"6�:�7��E�U��-�j�:}��5]WoIR�f-q�p�:He�E��W#��ʦ��ڢ*��Lط���ө[���i�U�u!���8;)��`vt
)&c���}�m�αJ��\��nZ$�%�f�B�'x�QS��E䒵�H\�zR"f�٫m,-��r`�*D��$V̣��p�f�I�e��W����
�QJjʪ�/!)�q�OH�J:�l��j�f@�d%͑W�n� ��%
���<Y��j�N��p����-���<u�q�A�&��ټ�d�\�\ʺi&��JhQ��L�����[&�~+yu�2d(��`�e�Kd�H�}$��%���L$�
n��;Z&��И�!U�e2mea;^_v���N�C�Rmh�=f��XL77��@Hټ����6���泼�jr������Bgg�'ڄ��ӗ��N-Y�	w�r㋭�Gfv2�H ��.���2d�\���J���.�����9Wj[�
��.�z�:�aJK����%u��[��RT���`h�ջ�e��z�#��/Wuǂ(��Z~2\栎dgLZ���\R�챨���t����}F|��:y�f��`�T�_�6TN���v�ڛܹZ�zg=�����ֽ��h�6ѡ��I�9�/�J��u��]�`���o�)�>V����9݆��l׭�-���`����<l��YC�P��0�K�Ⱦ۬<�]oZ�l��3�y��� r�LPp/�������t$��_Q"�.Z�	��!�É�������[�V�M���κwv
4h[CYW�ƻ)ѵ��}��լ���t����9��v;�3un�(�VX72P�d�� �64�ӎ7��#ï3���oN�4L���+����ݪwү�o�oI���k�:qiȲa7�Jq�޶f�J�oS��!y����9�U�7�\�le�Lt�u��Wt�t�z���Ոrnd�X��Ru]n���CY�+2�]�ԣ�)��Vj;�/Q���9���!�]�쾤n��Vr�\�Q��Ή�F.C/f���(���vз��r��Dꇦ۳��I�\��D�6�V�P��.eI��&u*�G�E/G5������r�����~�f�T�t$�/�8 ���ȩ�8{���Rm�3]4�g�V�w����xz?i�����M3�2�E�e�Kg�{S��H7ܽ!Љ���Z�;�JZ(pp�7]t��e�Xv�{v�|x�I�&��LuҬ3�4���C�CeV�޷�)�-�pk�_4��T������	�;ľC�T��]����-����[���^e�Q1hJ����b��݈��v���K��|��T������zK!���	Pƀr���6}Z�l��)��w�83wü�y�N~w��I��>jffP\.)�۷!ލ<F	<�<md�8;<@i`b�a��64	iޒ1��+���`mD6s/���w�o����@~�b|�_'��B+z!L0e#`�GC�;,��\1i~���>�2��X@�|x�
p�����yLئ�B��Ϧ]���g��	�h�+���%�oi��Q��5I�ؖ�t�Dh-�ȄP I�		�$AA	#�-��)RX��ro��y������ԯ����s�B� �0L@0b)@�A$5�XD"�D I�A�.�j���ξЩVKz�ZOC�A���+a�H>�jv!mP)��sz��v�\$�o:�����+�����pǶ��c�5#D�f�A��K��a�au!�}ݓ���>�Ph}Ī�(�_�>�u��<��D_y��ƛ�c0�Myx}���}a�q�vwLJ����5��\��Ѫ�D0y�.�%l�.[�>�Q��pG2&�ƃ��"�&�E9�������r������o>����&/j�N\X�4���9o]�U�2�`!L���t:,�\k���L����nW׻��r��73�֬f�����K�OF,�O 4��d���H����c��[�L@l�/lOu�A�@<L�ЦzN��3#8Qe���f��K\��і)i3�B/��W3���L��'�<�&��WjO�z���xrJ��Qg��#�8ʿD*p����%*�ڴ��?398U~�Uᅱ���"YC��8�J�t\)�:��{ ��B6m�+�2���}z��7�0��a�:qv��V�E�O/4��Z�	UV�p�Hdt��x��ow)���5�1��hܮe�o�ڦS�I��l��a˴$��iS�xw��m@�#M��f$z�d�R���Ȼ:��e4^MT%5X�$(���&Sh��	�2�b�Pe ���Uo��$(̍���!M�����:�m^�e�Xp�ur�7��{'Y�_wq�1��VLG�����<�� ��_s+K{�꬚��gf��gys?~�C~�=���>�&������R-k5TAo���
����f�x�W�M��C����r`��vR̾-�L���pK����1���aVcH4d��#ny���z����}����)��X��pf���2���Q8�������:7o��jr���w�Ha*���ls]�����C7�������i�l�M�"�f�v��{w��|����������тI�O�DhEw�4n�)[��&ٷ>ȈC.Y�]{"�!���۞�b��Sai�)�f����|���U-����}�-�� �<�D�*��v=
e�t1�wʰ=�\~���䀽�+����^\.�|{7[��@+���k�lٵ_D�r\}�H�ʏO�hk�@�+�U|z�����KXB����9�a��;;d'�Q�n	z�Vw9�;n8V��-y�{���U	��v�m*S�N���.�kfox�L�������W�_����2D� � ~۰f��.�i�3�Zf��'����f��W"�0+� Z�ɷ�2��UC?9P�^�؞>V-��VKP]�[�*M���\z�gS����_9�(�o����`�M:�F��K]�<؍Ν��叮�I�3��	׾��j��;Q#���wu��=q7�@-C6������; �C/�����L4-S��ڴ�5��q"��a���v���_gPQN�Nw����#P��s��T�zܓZ���=p�#����)E�/}7��Q�әS-8'��б���0#�;�J�	AXay[�O�����Ĭ��s�d�<{�~�L����U~���D�因������#� ,��37��7l��$U�F�����PAG��u�?2���y����間J}�˴7l�[�����Qc¶�ut�#'�9v���&�1O�+[�/��b�hԼ�8>��G�Cʳݥ�GFV|��%��Ο�"�3Z|���d��fT�������}�^Tx\@g�����B�p)��I"�e��'O}�s�-�j�im]���}g���K�������C�K����Q�`������{@G����!Вn^�>���t�b�?fz�H��|�4��n�)7ڲ�*�[���nM9����(�D@$!�]]�+����у;)e�R�D�h�wb"X��Ս3��+�i�]��9�ǵӭW+��c�#Yw�����:d���8k�z�1g����֌�Xa��.����"��or�k4PO�׋Tw�݇\�:a]N.s}]M�f^h�)��5%�=Ż��*c�R�y��i���8{WA�L�ߝ���p�=q��T6oưc�������j���.�vh�gd�y��s�)�3�s�R���X���!����\&t�64�kG{�zx�I�Z/�߫в��������jy��	n�u;<���>^�__T��lS�J�eIЩ�0��MD;*����K��=@�|1v�_t��s�w���wY�E�p̾^ǏU3�����m����פ��l����R�V��d�"Iߚ�F�=�ӭ^SE�W3��A�{���޳�⧲by�'����o5s�H.ͷED,p�Q/8i;�<�;̵E���lP�ٔV�m��t�S�i�5+���\7H�����\���k=r���SlC�;���£����֯�M�������Ktt|>n��xw=�� ��*p�Kv��a�+�_3�����Q�6h*�b��c9�ڼ�q�O4<��L�
1Qv�]rvA�R����{;��U�KD5�s�4aX�Ψ��������;V���s�芣��ѭ��A�+��a1��
s��H��L�,�Q`���'}PMr�	�Q�v�M1��Ѯ[���6���v�t�;�����5���Ԣ�|��F벴wD0U��Ս7UW���dp|�LC[��i�s��<A�tD@q�G���)U�L���^���s�0�|WwX��k�9R���R\��t���Ag��T��]T5y�]�>�6����&�������Y��:��k$��W�&��Gby��v|��-�;�&od����.,.�O�ȳw�v5��:��`�I��Jn:?S^8}cz�q�YE	w�4�v0�v��7k�kB��{���y��*��ÖY�8=�r��s*S�0}��p��,7�m�uN��wU�pκڣ5�"pE��Hd��q���u�����Ӿg�H�O��8�~���Uu
^pu�ۼ��Ad�e��G����S��mw>�rx;�l�G�'�)�f�z�&
�hEA���݋�QQ��U�di6���'��~$�� s����t��e�I3	4� ���"����G؇ E������ը#��J���RA�lш�$J%�C�(�	�d��$QPH0fx���.М�-��х��޽�Am��[��yk*�KE��y�-N������5M�5�q��+��]]#Á[��g��۴Y��Vo.�:k^��g,���e�K�U�U:1�6c���u��v��m����Qz,���1��sE���U&=J�׺��0��u/v��M������ީ�:9�¬���[��R�Ꮹ�&{���U�������������cu+U)./>\7n9�-�8-cSR��lC$m(���8�??��2���Z�{��]��k�YV(o�#����/+�ݠR��CV��6wܝ��h|���� <����n��u�����T����h��c@j�Zo82i�1�'(�75[!+����+f��T�q1�1��9�D�C!��hnz�mwl���̟f�G��
�?��/n)��r���vE,�."�%~�:�oH=��h�Ln'�T�5�:m���_4��Q.��[�g[͑����ͺ��&���ب5�qT?**�����1}9;Q���k�%�j�l}<�fi��������*��ܜ|�T{�$���b",�D;~�t!O�������a�q	7�*J�R�C*�r,���00e �q��u�'�P������U�Y��hb�Ekk�9� �=Ǣ�:���K�;����K����κ1a�V9�ãʒ�]��n:Q��N�Η�w���eNG_��@V)>�W��k�1���Q�hj�/�ٖt\������-Wf�]q�R�O ��ŕ��7����t@�``�O���.q�ppN�)~ىu.����������L;j6��m}�Ffm� �ѩV�J��5�!��ez���7[�����]�8�c%�?MWVû����wQ=�U?c����$}n�jD@�J`�Q� =�y������u8�S�_�|�ԟM{�R�͵�Xv��w��]�W�s)��7��\��':�K`Oձga:d#"�0�T܋޸�,M��U���U��ϸu�ϖ�o�D7��z��H?0@���l�;c�w�0�IЦ����z:�NLܨ���a�6���e���)U��Wên�f]���i�RϨ���<&��w'���7��V�	R.'�$;w�����/>f�抷���<U���:�B�����M�S���?	�� )�hx�+�ԋ�\3QدcȮ��4X��W�/'��u�G�J�U�Q�N\e���]"h��-���K�ƐC� +��$xo��I�i�2t���A涻�����;L�^� J� ğ����:�g_WL�Mu���M�/pnwNE�ʑ�곅��$�J{9}Y���cޙ���,�N{�W�3���Ҳ��ϐ���iA�t։�ffna�q)m��k�U��դ5&8��6z���y��E��k�F���S��Nx��=[��Ɠ�z��E_�s�Wr�5��ɾ�v���5��uP�z~�3�m��GnN}}>�2�;e�QV�f�o,�k��%Cm�ɷɉ�
��m�x}�����"b���ӛ�\��+��*�v��mr�t�̴3��i�i�"�@$#̫���@g���P]�e\�r��O���ë�����d�P���`%�\�̫��lՄ��_ ;`눞�{�U�[;Z�9d�ĉ��#�V�_
��A���KU'D;����]K�FP`^�����%��$	��x�
�M6��֌��.���;�7���#��v��6�oz�bn�S�ވ4� �M�䲔��p��烷�[5�W�]�U��C�W#����̹Ǳ�}{�w�g�ˊ���0�	�א��Q����t?��5 >H�-0>0ɚW #� P�2��+��/s��T��S.+rslvi��)
�E��`�I� � �`2�Y�KR�೙d�$�9�)�)��2��]c�6��3�!�Z�]�"�g}�$m�a�;@Q����g%����F��w]ήk��#�;�����.U���$Ǹ����[�.֦n���V�»����j��b�Ge����u�����*r�&?�ߗ�j� �#vI��N�+����8�q�D����K������\�������3��P;�����dUA SL�:1A�V#��y�ה��_��j�f�nŞ��;,}��[^�����E4���-�!�b�pc�,���-�tf�SM�Wy��NF���F�z@
����T�s���XP/6  Lk=�-q��)�k�b��۽T�\HC��2�+��,�����Kƣ61�,4HF�猛�`���u����XJ��o�Pt��*]�]k�7�+Ӑd?t^�1ژ5�"�g�kҮsO0:�#7���J�ݢ��4�ʧ���6?G��{k�^ER�z�@�X�2�k����y�Ld�l�ʒ��5�	��F*�\�"������S��iN���u����)~xw96]i�]ù�|��?�S~���B���n�N@
7��Ϗڗz�4��i��ϫ���\��ʾ�����Y%V���3��֚�tH�M�P�'N*��DC��$AޥR6E�j�rH�4��3��63j�a�x���\PR�1u+66x��@�֘�q�QS�ji�#N�O�fI6��J˂�F&[`��8�Z\,��Qa%HqS5!B��e$["X��&�=fq��SV�K�8̪�c+rW�����ǁ��-�k�� ĭ9۲��#*l	b�.��ra�F�e���u�8M�B�ݺ��I�ƫ�
�=Uv(�ƞ��l3.�y
S�%��dl	mQ!�X��_��?��D!K��u�����>�q9�Z/ainN(t���č�1:2֤4� n˖����d'g�[�s)���,/�VU#{G�3u�-�����Gu��鬕3�BW]%Jҕgf�����K���m�ިA�Ŧn��%�S����kD�T���^�;a�J�L5y�\�Jp���q�y��KX�nj����R��8#x���DN��#*y>,�8� L��&�2�B�M+m!ҍ�̄mb�]!)����wx�T�;����&Z��e�x�$�` ӄA�fr�ks]N\�k˧:;{f,vL�
I�aq6i�@ '�M�5%��B����B�ѳ=�$��K�I�*�[���� ��+��a7;9�fʩ���FF��M�L�ה TT)���ܡU@V.�����U9J!��ٻ�]�ۺ�I$�H�|H`c�!]f.�z�5p���b�f��F��� y0��r~�;	�{��ف>'E��j���gq����qjZ�h���k��ؕ7�7����v�����CIw 2�gR`� Y;�v�	�S)�}���o�7jWu��֢{|6�������d�8�"��f.J�kzzN���Z��{w�����|��e	-��(�ŏ��xҮDn���|U,�2�0�ie��������c�+�%�����'Men2܉ھ	�������-��v�̢�Ô�]ŕܪԱN��������9P,�4*���뉚'M�|{^�QF��Pxd��i@�ݦͮ��Jj�[�ǹ�[ۺ��6	�F�5�8g<�:]��'��î)�k�M���,yy����LN���282��~O�q�o�WK��2%����H�F����N�ĨB\�a�r�'�|u�Re*��up�&���2�I�}Qn֞
~&�r�x�X�.?���p"�uf��I�}�-\�٨l���+����c��: �_�ݞ��6�;f�	v�d!��Cۡ�,��8��'9�2e�L15��Z1R��k.	{
o��qs�w5�^���epzs^��K[H�u1x�|�t����+���,r��싅���[�]���]��A����A�{{u�.M<�P�Q��@���7��t���b�ӊ��3�d�v7�iO;�k�"m%o�l]�#;%k	�Ͷ�Q/@�ά�6���o�ZW}�!��V��.�����;�������/~~p�5�ޭZ0	���U�����(�P��J�@$h����D��P��"_t�Sَ^^�ٰ�O�5^-{�[b��mQ��Pg���+�`�|�0z����
����	��W=*i�lL�'����}1�ly��}g��1��ÕVpi����u�D�z��i��<���9�&��v�4��LD�!��j����w�͆K�eH����f�7��W۫�J�.���Plvz�>��] Mey��~*}�������OG�~��Ƿ��XkwS���{u�¿QK�ö}K;��� �79����4T ǳ�V.��f}�Wջ�S[��5-�{'.���j�L��̭*ٚʙ��_�p�3�V���}�H9��۶��Lq�����\%����2Ys/�5ydX6uC'�je���<̣UCv�!�~�z���8���N��Q���o��)q7��������5��Yt�]��kMW�5�$$(�4MM�Wh��u��>�ه�S� ����IA���7L�_|�r{�gu]�np�K1��Z+�7o��ػ�Cj��""	;���8�j$@L��n�I��{���2���F��D��4_<]¥���sq�s�h��X�:c��Z��U�F+��a&�gG��V���J�Ҷ����qj�m�/Z��O1�W������j��q�~�~�=�
n�{��ڍ|��#��'J{v־�W��V�9�(�n653�QO4��'@D���b�;G
�jy�3P��I�Kс�,��p�������U,�}t.�ʧ����o\fЁ�^{|'7��q�?y���+| ��"R.V�w�7sl��Ws��[/��}~�
���\��eu��\�i5�ʆ���f��R�,9�]ߧ"}~��%��o3��o{&篍����#�:7
��y��.�(�ӳX'��)U���s�#��Ⱦ�.���(Rܺ7b-��]\���5��w��Fr�w�L��U��1�0�L�t	e�5�~9�g��߽����T�[ܛ=��L`���":_�U8~�(>i�Vm�J����g�9��rj��!�=���8�@���^q���c��+^���$���ـe��<��<�Skw�S׳����g9��? ���r������u�cے}tv�F�� Yš(��o}{MO��rI���e�p��X5P/YDDH��d��k�%I+�.'�*½��e��f_��7��|�^\�X���pZ��ji��ۄ���������p�|���q�c��ku�3�j��<S�`��ʎ�_`=��!�Zr��M�B";g�6�<$�_u��lV�V��v���5(�o��]�t�a�1�t���R��}�{��[�{
$�hWI���&����{hW8%��������u�s��	�IY��_�Ϩ*h�}�j� d�R��Owa��oy�P�U}��˺�.�iM�Y��TsFk���<��p����|���H��˦�����w!��"*��l��K��q-�،ηӉ��){��:lJ�6���T���4�1TԱ��FXQL�"�CK���mgpVs>���NrR�M�[����������v�;ü֤s�ǎs�|2���F�H����cWCcr�.�ٍ-)S�37�� ���1���]ٮ�B2#w�:mlHjjt�����2{���/bI9-۟z�WJ>���"��+����/��;�)ߐ���+����� �so�Fͳ���zm׷�y���no#��_Y�W�i�>�AK�Y_R�;Z���&G�H���Ԝ0��r�(���������j�$ټ<�J	�����`��; �l����s���;[#��o2�v:P���4�~_�j8��U���圏���"�&b�|9�z6'�/�Wk��vۘ�wr�|8���"]ɨ�87���[Ck�xBVYF"�W����7��_\vKOL�3]N��.T�^ ��on�%�r��{4�3ϫ*_)*hwk)QA���U��/�l�>�o;������܊�Ⱦe
W�^-Z�6	����Cj,)8=����~��V��^o.�uK��tM[�����s�q��.�s%7-A��a$�d-M�Z�p��x��8�C0�������ʚ�\��6'��S:%���&`�r��/��ǎ�H;C��2V[{�^�.�޺+�xu.�,aܴB���̕i�'��n�-��<���`X�y���O��L�tȎ�~V�Y���":nN"���ȀX@�e�ŧ�y̙�9����e	[ἧPy�[[����%C�&z^��ْ_��شݗ�J*�NTt��h�B)���)��)b��hl����
�k�6Rv݆���a>z��z���������vbhLk��"aI��ܙ�;b"���S9Ʊ��x�13�N�~]��)��L�_c~8����a#Ph@�h������ܭ9<�+9�&g�̻r�%��w�EL牱E	M��� � a'��
%�'*��Ul���s�F���F��ms�Л;�mSB�B�IT��� (�R���!�ǵ:�r�;U�Zd�)����5�8��W���}��5���a.�i��޵��v��y�F�I_S�ֲ�g<�*����v�#�N��qOm�y���#Tu�����`ٕ�9W�%�4�h��>'�mOa|�o.!'p�yi��/�þ�w.�����S"�j�hw��@����Oy:1���n�)��e٧*_��ݶX��¡�g��+�N�5��=ϫe0*��n�C�[�_2��*i��6,��3U��r��5Jvy%W'���0��tt��i�D�`��.�<Rh�����X��ќ���<��p��0Z����ʹ����"(T7��E�t�����G�h��Ek�?^d�Pֳ��Jרm�Q.�:L6�SI����7�Ջ�6�bu��]K��{s����Wׅ7cth/������ku`��v��W�/�E��r�m	$8���j��̈́��N����ؽ�+$[�(~�o��k^�D��s/E�aɂVՍM���uxԬ�1���'X��Bt��}��H+�ח2um��O1�||�>�����Hs`)P��x�W��JNfl6IM�`�:��:�	�ϰh���f��  j\QL�F^�]��ɒ['*q4�M�$�,3�6�~��-�Gl�[��ݲ9�}P�u������(��0� 惹����2�f���7��������c��}r������iX8ׄ�_q��E��֖Y�y�i����B:L�O[�M�mܱ�utt_�Ɇ�e{y�]�#�߀����l�s��j�Z�Ͻ�y�}朥�#6s� �	��memBvh�=�1-�2�'�{�j�U�n޾h��z��*���I��L(uT1�8V=�W�C�R������O�rH���x��_���n�+���&a�ۻT�CӐ��*�T�O.��:��u:D�M����3�Y��o�+�۪�7�=R-��U'�7mt�0#�ًk4;�I�n�u��ǆ���+>�-w��=|���|�B�4E�DUy�n}��U���>@�u;���й�]nB{�&�-����<.��P�a��gC3:J����5>��(����ǃO�9`AY����ɘ�%�>_x:�u�������r� Qg��ﵫ�}��E���h$�H�W�׻�l>2������0�Ye]�=�d�(��o5��U{ؤ+�7`�f�3dY��Z� }<2����Su�������031�/�L^�Z��>�B$��D�����G��+0j�!���7��X>���/oT ���$	 �0,� 2P�.WL����GԻy���W�	�m;��}���7��][g�����2-/����P�_ɧ�dK�3=���ר��B
u/���'�����}qz��G
c̶��� V���W�=��|9�ћwL�O[r�^��?3�Ew>s^�ɔ�wN�ۧ'^,���Sʪ�mJ�f3����
c'k)H���4�#yQ��V�T�R�tM D�(�P҇�[j�4��R9)c�Z�ў>�>9�R2�����8+M8j3Suք�;�FE��CC
�L=�j��+�jdfn�])g+�,����j�n(�f�M<���"�a1��m��ZQ%�Q�o VXa���M�f�H���gt|�u�w:SD(Y��f�sYR���T����0����^�nT��>u�甌��z���;�fg�3��6�	���v[�Ĕ��S0e*�TL�U\גB^�_��d��]n����Jտ�����J�����f�m����.e��t�Iڥ��L{��k<���umA.��[R3/�Fi��k�k�䶹��Z�"���χus��̪"�a낟�w��
�N�S�=�
�:W3!�B�t�j�o�C�c�[�Cc�[��Og����̮�9���jd�2��r1G-r��)J;�唎;�_y�U�L}���:��B)$~�>փ��1��C{�go-�:�Եte�=Z�<�y�>B�h+�0Lέ�5����|������u����F�Wc,7�WK��c��OV̛��]�,<�vrf�:T�#"��}�2q��߳�I.�n�Ř��q;x�%�#g�C�rsb��T�������˼\N�UU�^�&��tȑk��7e�m���Y9ŀ"mD����/˺R�;�6��p �����������{8��*|ݚh}_}�w�N���fϬ?�wy9�������*�|��ޕfn�xhޒΖ�S��W�m�y[�,���fhM_�`]���mHϡ`Vz>Q[�\����p�M��Oi��C��D��PzL���E�n�����:��X���<�v�U�V�&~/UX�����G�뻺�)�ӵ��:�n��n&!�C D�d4橷d�-�G1��FZ���]\G-E�:���X^���d=��Lfs�4{h��+�q���G�δ��?�)]X�������_J5�J�K��Σ�w֨������s���΋��E-���@�*�)�1="Li���،<����@L�qCT=y��=�l�U#������)Ϥ�8�T��\^��C%�٘��{��G����pYB�b.<� �&���F����c��q�vW�׽�.V&�Y���#dw��� D��4�f8��@�XE�=�����*me��p{3ʷf�w6sCc���>���	XT@�Q�$�e�X)�����������*�l���;��+������u�|���#[�x�;Hq��"PH,�2��Z=����]Y�oa��2߸�K`�>b�m��#w��96�侪J�J��+U���to쓷�Qv�������̔��D�jw�W��ۢK��K�;�lӕ���t4�XO;-!�	�{�Ť����咫��:�|7��W-��N�r'@|J�ѽ������|�si��}O�˟j�|��ȶ΋QH�'��)�\%�5O1m�r����R��d˞!ޝ�V+�Ȏq&	�{ꯊ+ u3�(@������m{��*�u]�#�]�O��J�x���U�^:�>?��O��q7�OT~`��{�ߖ)4;o��qy_,&���B#O@wA�{}��;V��U�p���"dY�.C�6��$�}�'�"�=)n�T۲*gM�ex�)��[�x�V7��t`HS�X�!]��mfk�v�~��������1�w��v�r�K��ZUk뺵+\X��ל�K��E��}�����)��5+���)^�X|��D���䗞�Y�zP˛��}�����P~��#������}y�����=����� Ke���'պ�EU���`�]V�G\'�v~=b� ��;�h�\���Ip#���k��{}]��.��r��&	���1k5�cK8h�-+���R��h`�]�/��x�yL��z�Nξ{fG1�v7�U�l��:{5�g�X�V����g���O�|��³�A[��Q>"�Ǔ,���z�LBJ]knEw�t�����x�æ��oQe���4�g�S�놀"�����C49؏@/��F)c¤����j��{�{j�?�O����=�dm��Ǌ�ɉ ��"Ͼ�2"�Wv0�"�3���8�u3��J�d@�""���_�|�g��㹚��,)".�F�@F/&��=W�
Bi�����s�5���#nd�����`��0ݯr�5��Ս��	@��[_�C�6z���J�@�J�!UF���k�X ���y�d�ΪX˶8��O�X3:j�z���9y��[u
Ԫ�m�3R����>����P'��R��<1	U���`e(|�t�� |memOK\�;MG�Q�[���y;����'��&���gUP_DH��b���:��ɛ�����#&�4�]w����f,�y��Wd��(=膇e��d:��l�Ƈ�0�WΏ�Xu^f��6��5����Ѝ�>�{#�視��ihbo����٭�c�ڸ��4���Fb��X�`"�^h�K_܋��ll��w�L�f���"�����AĩU�a<�:�]�����5�.#�Mt��95�P���� ��@"DG���   �� "	����� DD  @ �L @�"  3 @� @g�D@ |D �@"DG�x ��� " DD}�������" ""?�:���?���~����"" ����!DD �� @ D���?��D����^�� �̏h��q �¿� "#D " DD~���D���BX�D���������BD� D@���� �8�޿ " DD ""=����J���l@"DC,��~�� ��H� D@�������(+$�k92�2 ���0
 ?��d��D����Tm�d*�BAXڈP�#
�&��(�)��JR�m��+0��̶���	
$�R�mf�*�*�� ��J�V� �EQ(J5�lU#F���JH�J @�Q�*����AU)*��*%J�A@����
*�UT�i����YjUT�B֍j��H�MJ��W6*E%N����6٢�R��
�5k��R��f�BkmP	�*k�UhiJ��U[���j$D�5����	SCU�0    °    eAc:kmv4��X�m�R*��UUf��V�)	B��6�H:ԓ��l��E*���V�Im��J�**�$5�$	QWmR�`��ںЪ�+��r�]P�n��uMV��v˲�]�����;5M�Y4v�]�p�*���n�4����w:ݴ$�ںM��cP$Rle%e%�ER�S�h��T�̧L�EL�j��t�cP띛X뜙Jۙ���E��Z��k2N��n�N������ �-5@YN�X��	Ze���l.�ۡ$�-��(ڕ�:]P��9�j�S�:� �M$�X�  ���F�"� ��L4P	i��PD����T�U!.�
H���� h�3J��� (6�N��MQ���Rꔖ��;���( &K�i�lt�TУi��u\5�ZY�l���B@��UR�;�[�RRΜ�h�]��4h��@R��Vh*�c�.
m4m��UV���j�L:j��J�M�B�7UP�)Gm�*P�* �9D�5����E����Ml�7�h,VCZ4�5`J�����A)J�u9�������m�,Q�:th�d�Ċ�PIF��U)�Z�r�Z[
���t�  ��u�mA�X�;�Slu�MnЋ
d�d�:j��:�]n�t�ɝ������v�n�NS�+���Z����-�؄�(��"�IRG4i���-l��&�mUwP�ۻt���ZgnK5��v��Ѵ��b�m���\һ�T�ts)���f�hW:�t(�rp� 
Ct�       =�A�J�1A���a%%T�cLF�  ��$�R�A�S�2CL��bJD� )�6ĎC$�����Tr�L��Ȫ@Pb8	����d|���_|�<���� D���� DDL " ~� @��D"#�@��0   �����p!������x�D�]2*]Z�ЎX�4E�&K��ԫ����mfA�d[i���1�X e���٫�7��Qw?R�m3Q�y���+���vs���oR�R*=T�3"�1P:Qml��t<��tN��d�D�����l��)"̿��^���~[�'r���|� hB��� ��d&3��A6�E���UЖF�nV���M�R��<X9UÒ� <;6�*��Yk� X��!~J+2��Vu, $�K�$���Yl�5�"�.`�e��%iQ�Cw0%��P54"!�bF��)�b���	�E�T��M�z���G��ѯԦ_��͛Q X�Rk�e6ۚ	(GO㛏 �Q�7ٯE�ФV�z
�����}J���[.7�[�Y�Xи�R�@Qٜ�L�a4it2��wSmcy��z�ݭ�j�Z���bYhVVąbǪ�����@��9�K��1m�fÐ��r"K�r���F�{@0�����/J@@5A�䵟�֋���i��L҄e°�
�=�{q*6ԉ�z��}g�NB�����2�թ�iZ��V�m�.��v��
�����3X��T�ѡ4X�C�H�FU�N���~˴���,�sX��ab1'B�b�Xt"�Є4�ʼ�n�b�-çJ˦,�U4�3ǖ�U,I��Y����[�~%0���ՙ[�Sj��"�0U�:����M[�u����9hc4h��R�噀��a��)=�ҙF�r�-�t�ܥ��aw PkF���bW�f��-���L[cs.P:�����I�
�ǡ*��dQ+�84�.P�k1�zr����F���7:���&h�-.w:��\x.~����r��5��
t�ɪ�$T��+7(T�Mc��3��tɷ�����e��i+��Rƭx0\�I^ܰ����
ٔ�JX�&�V��t�nVI!*Q(!wy�Ԩ]d6�3Xe@��MÖ�W�:љeV��n���1L@��ɭT��e(U�
�ޒi�i�k��:̡5ה�0 �$��s����o�Di�fIV�"����'��J�J�J�c��w�--��5�\1�ݱ��4���H�p�W"ƀ�En̓pb�Xh$���^k̬4�m#x����w&���HBN�	�7����D]OůJ��Wi�y\Z�+y��l���-V�Dn��E{�]:,�u�PT�Se�W�L�hӲBsQTpj36����lQy6e&�V��V�W�O-( ���Z�S�S�m��''/���冧U���*B��#��6�WO][��]Q8��(icώO��Uz�B��V�q�0�9�h�@���F���%l�n��s��'9p����k��+J�����s@��O2�l�!7~�r���z���*eJ�j��}jR�&0���1�,�7Eł���cs,�:C{t��C��Ս�XJu�"���f�M1�h�ãR�)�/@2��t�Yk�F��퉵3=T���,�z�HX�+h�f͚�氦����FV$��j��H�n[Ѳ!��c�Y�X�!Ӻ�5Q��Co-b���K51�e���j�!�����{[�.�)-���f̫蜱Ӕ,��q��M�D�1���3i��*���@:�V� Ȍ1D=��h��}�#�3�kR�쒞t�wi	X?YT�e'7�0K�yYt|��%�q�-:8eFj��ֹe�[yA;�)�R�H0XO^(1n�'"��=D: Zj�v�*�,���	��k��*��ie(L���H�1+M-�n���Z�e�Pn�%���6�kt^]ֺ�	P'1��xw
86t��4\0�ͩ���a���4�XNcХʷv�V�j-���I�r������4A�M<l��L�i�Ȥ��ŵ��v�퉸�B��˻k �p�%ԉ��l�j�'�Pb(�i�(�W�t�Yh^��]`Su�6�]X(�����J���83J�w��:,P�:h��3ݡ��V�d��Mn���J�V�1��+���nn}q�f�z��$�l�����c,;y�k^c*�����̉�������0���a������Ď��d1Іe洚�&��ȳi�7Sh�D((RR^7m�.�(��L��̆��;�%�ksMn̊Q��lËK���b��1�xHO�n��L�R۪Xb��B�L��t�\A^j�F��0V2�F�n�����N��˼¬*ܺin��0!1(��a��hX�@u�'F�]��1��V���Y�%�%�� oa�,-;�FOҦ ����P����� ܳ�b��RI=@h����JfŽ[���Y�x�ӁԲsT�d5u��m�����ڒ�bCXB�М��f��\쵐�w���T�e�u.��si�t�t�È(�{hm����j7v��e<�x�.�ؓO2��a�ӚkK��%@rR�#2�a�v�-K\R�aWQ�j����;�T�w<���8����e�oF�*%�4pA�����.%�-ZqҌ^f4�t-��4�FQ�`I�]�Z3�"�jS���D�,ViH�j#���ѬB��ܛ��*TKr܄Q�����#�g ;*d|�r�3xZNT�0��]v9V<%[4�f^Zb��>���Z�#���W���#��$ݰs`HlA�'o)Yi$�]l�5�9	:p�.�*A~�oX�h�^��  ��l����v�L@݃^p���`�kr�FxC³SH-�k4�wuUL�p����8{��2ԣ!�e�2�1㼵:4q�QTi��QmEۺ���\;'+te�Ӣ0��L�ݯΠ������b�7A8�V��
0�k)l�GCcVrb�Щi#���-�Ǐo7�<"���X�]O2ջ�D���FK1�PbɆ�,�ݤŭiض�����Y,�d^J*ј�$#r^������8D��H��2�1U�^������a�dU!��t�{���(m�@\/�D��hĔ�x�uh�÷5�2�I���1\:�-�VfnQ� ���Q:���6-K�fm��86�"qB>�C��e��)�:q����=E� ��R&���j �/%ڶԙ&��4��*��^�(�����bZ�t�;�3U^��8�#3P��J�
Z-�m������V��e�����C����t�تk�@��P	����l��-ŗ��Y�2U���r�դ��Xå��7��Ø�X�.9�)	Rn���Or�ŝ�1N��ɰ�t�j�/%��2�B�Y0����M�H����HSBa�Bɫ��@Y��,���X��J��bP�E��ۋ�K�nی�I�t�p��nlSj7m )<�)�*ËLS/����q�,'fGV�W,U��Ca%�A��/�V�ji]͔�ǚ�n�FRun��-�A�ӮM�K��������ۼc�FثZ�����ƶ�G��AZy��Q5i�1h�x�k�1|+F��:C��P7@���ʴ��4KږEi4,A������{���^J)JY�(M%�7B	t7Y�ȭ�`�ksv�	�*��RQ�QJ��;i&G����*��d㺙�iMܡ�f����l�te�U�æ��5�qF�A��UX�Գ��N�T
A�c̦��썝$�x��ɣ�T� J:@�.s0����]9�u�OX��#�g/,�UN�p���ut�n�ҭR;C����N
�S��֬˭�k%�0(Uf�L��5y�D�/[ٛ{�N�l��������(�ҥ�U,Ѫ����zc��,d
e�f+5�]A� �EW�ɶ�TM ����3A�LrᲷF��2����/r̀HP'(���je�Z�eĆ=j��԰��݇�vRj���B)Q��W��B\S���LB���2��^d)( ��՚'�ŗ�#e�F�0�'�PT�ܹZ���l�t�IKa�5ޣ��4�a���8�9���W!�꥜�b6��˄�Zb1���#D��Ia^
358]�3ACnU�+���I�mԣ�f�L^����P40��7��A����j,��T��Xi�U�M�<�r�N٫�r��uH=�X��\�!J�CEe��.*�س,#���1�ճo
%�� ��� +7���t�WZ�<5�ֵuz�hթFė���ڕ�C�Eٛ��kv�`pJ�YwOǕe��I&b߈��V��M��mf������ 7z5;�Ԇ$)n6�gf��J�,���=q���1"���l�D��3E��9U:ΆI�z��{34m# ����m�F�f�+d���:�pٷ`�Z�:l���\��r$��Rh֝�Ǖ��!n����(�D���e�!�
���R��+kU]�r(�Cj�ۊ:�=E,[-SV���=�sMjo��݃w�æ �D�ni�Ǚ��Նvb��n,w6�:��`EMBN�H��Л1(N��Z���]�f�HX�$��bT�xT�TͲ˳v��15��*J+K���iͭ�^in�.J�H���:�5b�٠j����T�B�`�Ø�:i�e�[��,�3)����u�j�H�,�[����ݰ12=�[�]f"�OL�Hdt����[oieb��jd�T��%,+�zA���,q�v0�h%1�%��A�,����lʸ
�0L�i"�T�d�؛�i���L4�'X��.�ک�~ؖ�սF�-m��Fld��&ebH�7���Ui�4�X�M��еwz)m`��z�Gu�t8���"��Yv������E\s&��Y�d�PD��j�C2h�Z�bAK7>
e̹4�(�Kk$U�[H��T֬W�\ʖU�MՀp�q����e���TA/�Y�`�����D��ԭ�B;tt��=�M�Wt��]IF�(e�N�;dJZ\F��oj�v�?iX��t��	�f`-�ı���
E���R����-՜�3ha��)ᳵ>T���ˡY��7�h�Sqb� bx��s{����ޗ�Wt��	�/]��Xr��4�3m�wZ�@�=`�\�~6�� �r�@�}�Vj���]B��v5�[�[oY�Bؖ,��"�CZ��ě��**5�������h�IY���+6��,����a���	[iM �a��cBɹSNP�!0�$�1Jڙ6��š9�էS��s-�:�V�T��sDux2��	B�X��-]&�p�&T�`���n�4a�&���ĽW��詬�p����x��^��Siބ����?[�
���TQ˖y�,:Jks6�n;�5���u�I��~2�9EhS��8t�Td��Չ[W6�j�e%�V�b֚t�䠅a�F!U53�-� Ȅyx��{Kѕ� ];d����s1ܹ�Q,�w�ZY��/u봂׵8+0#C6/ΞZZe�JYɓ-�Y��&�iU��"�����-7)�#�#�(+Զ�Q��L�%+�=��c��'p(�nt #�h���cv0h�`��Sk�h�9rq��7:�F�G�&Eb��h���Ѵ4bx�����Jo��欧��v���X���X�����j���[m&�8
�˷,�g���r��6s��y��ml$lYS���.�8R*D�2��(S�u�lX�;���ݫ���[��6�y���&_��o嗳6�<�"�O��T�mzP�#��6�MV5RJ�f���4ٳ.h�%	B�,(*gke�C)���F��$T�đ��%76e H�ob�k�x�fe޺X�<��m�`]Րa���̻N�{YZ�/ ��dU��ִ�[�N(��H��ݩn	�{@Sek۰�~���kTY.\:ŧBE�
&5��=+p�����cr�̅���t�u4�mL*��0'�q�zm})�-�,ܺ8��1�w�Z0\�k�m�d�n��,6�+��r��Z̭���Dԉ�Ҷ�k+[�~{�)%���K׈���i��/4iF^�u*�z�"�`YV+���Zr�YQ`��E���`�[>����q��ǘְ����l����t�u �2��kTO)�kKWnR@cPVܖLܩo5e�4.�
��:�,pnjj��@�^
YIeHS�Zec��4;"ت���8�e��f���4Y��B���'R��f����L�,^S�U�X���B�J�.��x��'1�F�˸�[�Ɩ���r�Z7V �?12ӈ��,�?e6�?G��ʅ-� m��Q��*�J��i�o�R�d\�V�H�9Ann,Ot˧h��0ιY�(��x���e<8��_׶Rw�0��h�-�w�-:
�n,��A4Խ�)���u nإA�r�J�]�t�W �Ф1�5f+��:�o��H����S��@Md�T暳�%Ѯu%��C��,�B��b+\�3��&���KZ���|\�i�9vnm��˧gj�2ZX_�a݄���n\�Z-�aa�Y��͡n�#��e�Qv��z�/�5�4��I�,(���:�w.K�����F��Vanʃ��f�RY���S�?(*�[;�o�dͷ��J��.�e�6��+������%E�R�h��FZʰ�V�3-��m�:wPd��6���l��\$\
AB�%��U���3r�t�X���sQV���1h�颡�R�Nb
�n\b&5�p�&ČM�M����u���"�̈т�P6M�o$67ulCh���կ�1P���&v�
A�ͻ��-�r�;F�&�z��2j��ʀ��a� -���m5B�M�&��kb8Ա.�LǪ>��J��'�!.��h���a�z� ;����v��4���ސk	�Ͷ��yQ:�=�?5Oqf˘��M���9'�M͂��w����b�[ȯt��0v��vǔa��[k ��I�i�w������aT��+�ufG����^��l&
�űCb�"��M��l��54��S�l���W�j�Gd&>}$o��m�{t24�p �e�˺���sm��#}$o�����Cm������rH�6y.Y�H�I)���W�f፮�%��#}$o����r,̜����N�Ϻ������}���{����*7�Kx�+��\�\��s�������t��Di.UͧV��\\����Ѿ�7�F�IF����)�A��J>�������1v��_>[�Im�ϥ��ǹ�$o�KrBy�w$��'�w6��wf��,���faye�:�ģ56���M�r�^M��k�[�Q���o,8�y�>�x���W��e��v��>LJ���ub`��\�gM+W�u.�p�{�\����%n�rм�6)��r��ֹ�7��1�-�7U�D��@�[b�N\�CA[;0��A�i��8DJ��CMg퓳8)�C��{�T���q������5��[�>8�7n_Ɩ�%d̟�\h|����C�|�	U��1��;�\���`������%��t����ξ��)���I��+�4L�C��V7�_c|��w�m�s�.���i�����2�VS����ڜo7�Pٺ]�.�5��l	=t��kd�������%q��
xZI������v��2���泴��+��.�>&�Z�yD�'�2f�[o1D^T��� u3�r#�Iۣo[w�r����_>����R)��,ʦ�k)�}#��xe�u�h��{Z�Õ6�^Yݔ&�Fwz�
P�=��`l�����ƚ}���݋�S�Cr]Z��6T�ír-t��n�V��fi@2�ycE�T�l� �^XT�8D�]֎�M�ɣu-�;�l�9�v_tAbc�b�ff^Mv��-�ܵ��ͮ���Ca��7ظ�R��8�ն�g�����e��:-H5��vK@��a+Q�p��	:�LѸ�gP�"��j����E�S��9�u
:l�]�-#�'�]�8k7D��@�v}�Yɬ�v�Q��;�b�DS��
Eu�S� �L�C���:���Kv^���%�g�c��A�(]dЫyݫ�b�(�f���v��tRЇ+����t��Z�����7�y&*Nr���E_+Z�V��;��7e�@Bշ�����F��M6��܊#n�v����L��m���Ͷ��+��Cn�j���v2dAnW{�+Gn�]�Gt<�RWa��6"�w�u�7�Aںww��!:]��[݈S�f��rƅ
;ӑ#��WJ��A�q�ޮ$5҈YMfT�}�K�<o>����m��&l9+�L��U���Pk)mua��I�ۍ���k�D�0a��wmѬ�$w����"Id�4��;��b$�=[��F�ZKFe�X��m��wdM�V��mps�t>p���)�x��˽�	���`�L�̽�x�ǹ4*�F���@:�g�˔�Z�m;U�q�J(fk]��\�Q���$���j�5Z7T��f��� j�����-�:��*Ү�TH�\�F���ˎ����X8k9��5ܓ�sܐ�/փӲ�fV�.(�iIv�՛�J��ݍ�Λ f%:W_w�삱5�u�7oIK9:�%�w�[�k�j�F�DQl�`��jH������d㙉4.�h�˖֝�G�"n�"Έ@��{K�v�OJq�V-X���)��j�����uX^��cס�K��,Vq�q�r�yt�Ӽ�

Y���k����|1��Bw9aZޮ��SNPCK�»Y�ڏZ���R�S�aABV�u t^vᚱ���qF��>�y�S�~��ऽ{\�n�tQr
bK{.# {,�Ʃ�e��"Q�y�r݇���:�+Hܥ��2����7�	W��F,87�;qNUqޡ�S-79d�ڶ�bVn���o~�{�B�D�:���z�3}0�b�h*�2,�C�&�,��O�İ�OF&5��97�'�<�"�=��霺�3��V�i�t�hT�J�˭.����(���� `[ê��m�3"��8�(���u��+��\ȏ;8Yڳ5v�����{�R�&)�+��\�L�Q���W���5��SaS��ƀ�9�鮵Q�z8�G�4���pb�#�9s*$52��5ve�Җ.�l�/-Վ�[��rk�8�Pt��jK�"x�{w7� U�1�+�`=��EAܰ��Jt%�eh�6���:�}�
��[�\.��W����U�
��4Ss%�\�d�1 f��!Ja�E��u���t@�����:5^�W[���6t%��<Z0��W�^�iؔ�e#Ȝ��u�2eʖ�&n��>���:Q�Oz��A�O+EK�p[������ar�>��+!j��fW�'B��6�q����mZ{΄5��R�]1�+�����n�:��W49<7rK�/{�ż���PT��ݲ�r��*l"���OR\{azi�����{31ed�V�=��9#�ʓ�ХO��۸��:"Z��ә9�YGv�C�h��l��\]�;�I�>+�vΣz/e�Wx��4;�:���s2���f<e�)�n��u��+�7���Vx#N�fɊN���ۭW�ʹ�WJ�ӇΑv�:���J��ޒM�٩p�ח����vJ���*����� � ��]8��hx`x}]�T��`΋Yr��.S�;�f��st �xe�]ggdT/���%4.�/_-
\�LM�t�o�/_;ސV�\A�%I6\"�U�c@�\�w��A��4������3 ���M�m4���E8�ޚ��otm�R����@+�C���.�\�\qg^wGX�L�{����pK��m�f�v�n�S#�\�����{V6�����Fb���.�(y�]��	)����m�ۥ��
e�.����V+���eN=1ҙ˦�qki:�P�&�bb!C�����Ct�efh���/:.�]g4��=��A��"(��N���P�,�t���ü'�;J�L:t*](�R�f�������}{���/<i�(�82xJx�L�Q0��Ǘ����Ar�nj��D��A~��e'�OwI��*�ʐ�k����5�D����4�|B�H:v/�j���	}j7�K;
�C]�"�jC�2�(�eH��U�Ѵgw)��7"#U'�D�����m�}3��u3y�6�]$CB{W}I�X�񶨫�+M�Qä�m��� r^�%�6Z�ő����4���o$�m)��u��_<�sQ#���ګ���0JB�(��R��Ӥ��ah7n�E�H��jZd� ݉
$��`b�8�����=��j�멝R�e	��Y��:dř6�d��f����Y��Z�Y-���Z��F:��s
Aә�ok43�k�eaE���	��`��7s�Y:W]2���-���\MV���JvQ�|춧B�n1��Z�f
�E��v��D�*�0'A���FV�]��i����/���WZ'g�V��8�5���d�������_�_�i�)�����O��έ1�9'GQ�wveZ,S[ȇ��szj=�Xq%{��콐S\�BOW �d1R�L�N�wD��Q��[u*�s"S�����*��]�ʍ<հ�;�p�p6XW�_ahz±���ǥ%v��H�]Grݧu����F����,�g�`9�i��bJnf��+���x�k2��í�d��SA��ʕ��&]�=�Yj�-t�EP�ifaq�wnл��qE�+�_��_�f�U:E7	� ���[�����7�`�'Re��.�f��(�(6�VWY�"P�L7ܸ���יJ�˲��w�(h�Fd���kn:��)}�N7s&LZΗYI���W
Q=�1і�.�a�y�o0�T.Ү;���&ˋ��u'��]r���x4���Wp���X�C�o�>����ݦYW�3��W�LS8%�z�>|t�m:� Ͳo_\��4_3�scp��g^ތx �R������5M�_^U�ܶ	�3��m`�GP�L�ST��x].���jg3 ,�N#ٷ�KL�0�]ti��x��K���T�Ԥ�xGM♀�7���7�n��W���¯�����z�u��LZ�n�n�@엩p�4��h�Ǽ�.� X�	��Vi�f�nN}S9j��QO�S��hD䱛)	��sb��Eb�vZ��	.�;W�w�
�nb�p��a�+�pf��ͥ(t��z����X�YHN<7>6z���O�%�J9Xz�>X'c�_w=g$(�����4��<-�*��ۣJe<�f^kp�ýLN6�7�����/0�U,@K7V_�љ*�v��	�Fn�2]�����;�T�t�ٙ%�t�'�	5-+��^:�u8����f�T�Hޢ9�B�^!G`�i�x�6��]���!��cz�_U�f���4�h��&d����{X&���L%�}z(.au��*���-���ݼ��k�o!9�uv������÷���{2˷B��c��5��;��1R��S:�H�C�x��nk�:��>t1K|V��0�A�7�M��Yx1�wY�9��:$����v8�텮�Ŷ�պɶ�Z��Y�����'[�:����R�3y�i��hm��n����{S	Bj�a8a���)N�A�P�z���_Vn`��G\��̓a��Y\��������+6#���۱�u=Ra�y.V{�b]˞�-�����;��b�l�7$V�<m+�̮x��JN�AH�]n��0��C�Xں�@E�M.�욚ڄ�u���q�����u�J��N�a��q���`�(7Y��4h���&>S*�����a��+.΋Z露��*���0��	r��X=ΰN�r[}Om��x�l��ko 4*#��q�Y"���e���Ӎ��EY�����8�Xݛo���WGQ�t�����FIt �Id��F���Gx��v�)��,f���́��*0x���"��uq��f����M����ЍX�ޚQ +��M�Vк�Ԭr�%#�T�sݥw|�U��b�T$�k��J��Ff�����w�j��.�gn7y�܌��JЕ�'�U�xsr�3��k��3���˺ht��媸�j.�&���+e�3��4�.	x��dy�m�m\�l�J֑���#�B�ڎ1ou,rk]hLٴȬ'(u j���/�.�})��Y�v$�ˌv�@ޱo��<�f��v2V�Wԉk3����k�oP�)��r��m��:o&T��Ρnd�����s��w����s�Y�3o_YO���5Wu��/_p�nM��A�4os9`T6A>�5kش.ĸC�R����<G��ٝ�N��wq��k�KN;?=�gu�;�Ŋ-=i�r��v���;�[��-��2��`l�2���e�Gr�ƛ�57�$X4w�єrI"���<�I$r�"�Q2�803]F�^�@�I�tK),�b�<�+�̚�t/�޽]N`�$���Tp�^���{��"ZSV`�~��jʲ��{���o:�`�3GW%ڷ���j	�[C�k��ܭЫ�U�D�<v�B�&�ILR�X{�@`6���
��Ņ��6'�+�JMt�.eu�x �)k4I�t����+��hX[z/��#R�[D��9�90��&���5|��:7�x�:�$٥��W�305����7f\5_S�t�+.���S�A��GZ�^���wH��C��b.V?b��=���![��%�3YA_n��:V3q]�#Оn�j�>��d��A8L6D��~�}G8^
TW=�X޾�)
ul�	����5��h�o(�)!.���JVZ�VQ`�Z̸�s1KSE*�Yv�����O��Z��`�q"�^��Pڴ�e�5P긮���Hv��B_V���3�[M��J3��2�h�Z����h�q��8T�3]5r����˃⠬����.��6����}q�ĨL�s�j�[��o(*s\Vf�����[W�V�ܩ���Wg��.���j��|�l����֮���J{]Y+�8�X̛eJ�[��������ki�IZ�x�����_�����+|(ea��\��u�#֐��Jɝ@�u�)��B(���,q���f�`�5w��Jɬ�jT�����>Z�V��.p�z�}1'Ӱ���Y2jb�2���+j��'2֥y�����o"k���p�3.s�γ�:�3�2_j�!�-U��#km���?#��]s��w�q���V��������Ԩc1�d���8��=@�!���v�hu����Y����L`��v�*ۻk4A�WM9�0��<�]$o�ҷWc����n��NC�p�P���+zV����	�o�z��z�`{�ìU��A�K3��n�}�GJ:E�,�6�7ƺ5�C�*�ʻ9�V�MNy�s�o2�-����++;��8��J���H쵂�2�Zj�S"�.�yee��1jG ��͠7DD�\���3j-�O}�9`_gQ�����B�!�U�R;�ǔJ�	�����
}w��KG���mbp����D�����F4$�:�9g'��1oG�ƀmVӢ+�5GM�m:՛�b<ԥ�5f;�JQB�]*����UhP�����! 0�M�šx��m�� ��t2�b�x�Va��t�k(uueb)<Ŋ&����1�55Ħb..3�nP@1f��yD�u��h87��|U��m��v	-==��zKۓ˫;�i^�}�cE �������a�W��sy�RX�rؑ�E*�b�ݔ2�G����3M,*�og~��GɃ�3������.��Q�@`Rc5�WU��UZ(���2:Q<	��Y���3Ӳb���<�l��s �^s�Mi���I�M�m�k�����0��:�%4�<�K�*�1y�/-���,��7:�^ugۮw2��y� eg*�U,�g2��},[��
ۦ]�za��h�4��V.e��;9���.,��M������G�.L������=Kc�Ԭܶ���=[Z�ͺ�-I=X�1���]e�5�Y�9��n�6��(�����̌��*`�3J�ܦ�g�mp��D�
�+vX��g'p6��N=+l�ּ�U�|bÖB��6S�����'Q�:�Hvp�dq�r�[N�d�;�^Y�6d��H D@�@�� DG�@��1�"  +��x_���͙y�*��sD�J�h���ݬ<�_V��}�o)�U�J�oa�"���k�ǳA軬�2�e�u"�v���.�˷�(G5S�p��]�E���W�v�U�ur�wk%;��.f�- ZC�]n��� \�Ԯc�A�V:�M��>K�
cH���9ٽ]�ՂTy:��Z�m���գ�IbR��Yb(�i��-e,��O�F���Y������qV�Z�J��;�ºsp�!���B
�V���`蝭��ei��{ľ�q�x5,BW]�j[�hb�ڍ�/��^b�_T�9���>�Un��j�|ݙԟ靋�nGp�I�$���r��@躔�7�����P��3�����X�����;���h4��P��u��	V�~�c����L��̺��!���:��]��͋B'`�{Ceo�v/�jY��꧛a�'v�wC��K\-n�v���n�����Ø�1,��ZTR��l�U�f�L�DCΏ�[�kz�XV��V	db��A��e��v�vp�Z�ۧ,>Ԧ�[�"�`�;G�B1]�Z��nE��vֱ}\�ӌiK��2?��w�o�(ﻋ��;�2u��ٗ�QU�N�E�V�ZJX��_6�zl��z[�|xQ5z��N%5d�e�,Ά�wg	:��(�|u���N�#z��w>{*1�>����.���C/7>�)wT�Uq��)��7z1�C��uƕ{�S�}" @�nܩ�>��^uˡ��ff�r�r��k�(��Yc��΍e�҆G{�8-����l����uko�
ek1&s{K�T9AʆZ�����ٵb��gpݴ}���֌�z�T���6�{`屧�:p�u���ˋ��ٮG��y�fꕺO���������:�}][.��7�V��>`�W����h�2�]�z������DP�=�%�Y���Wwq⦟0=Έ�����e�ƣ<=�m����]�$ko���{7L��	o��}��*a\=���m{k|;��j���lA�=\�ӽ��֍���i��GW��ɦ�;9x�>u�6�C.�y]bg�pwԬc��t�!�����k �p:�k��y�׊�	ؽ�lD�~��,h�y�خ�Uwl>g�s~�V3��"u�f�Nc�uwY|�%���Ӹ�P���F���#���F�}�Z*�hݳY2�xX�x���C�x�K��Ǹ%�=�Y��u�:�>��V�"�� C������W&�B���wM���K���9�*;�q�"1|mX����ˤ�>�Fw,��[�nCʧ���4�r��^�k�B_;�J����Pl�z&�yq�k���rm�<�OVպ�v6<
v�����eD�����{F���9W���ŝj�<��f0��{��A��Ք���Pu�t�4p���yh�W�[d�.n=5ڛ,�����F"���✖�.u3�����	���/��*b�U��t�f�N�~�-��b���5�,�/pmg ojkO-������t�~�ˉ��Q��FL��2ĭ������GD�Q��jjFXy���L��u��`��¼��D=��p����B�MZ�3Ҁ�<�+'�ٶ_�'��)-XVR���fW�C���~x��EW��i�)!�ec>��@S5��Rƪ�cռ��Ú��8������~�薋�~-�7� ���U~�I�G��Mv��ÖL��%�t�	�i��x��U��(0R�v��{:�N8m�Q�mI����7X�������鯒�c||8yDJ|�21�Ck�ָ�q����'}[r:S��7ֺAτ�xio3��2czh��zD��*�mӱx%�+ZS-g�G�vƧ��l�p�k��x}S�<i��]�^��X ���`����VU9^�M+V�K�A�I�w��گ����hW�ܱi�TB��׷��U���s┻�:�"Z{ڭ���h���~y��si̋G��bS�xi
7�j6E7�"��6{��yݺ$�(��O�T|���m�sV(�.�����$�@��O{�iEH���T�>�G�	��Xj坚�&��2k�Am�v��u����K�Z ��Z̮\���O��Lؽ�E2w�#I�G`�Э�W
[:��L��ü׌}�d��Dئ���辶w��L$ײ��^_Z�'������=���?%���]
��y��G�	��6o���ۛ�u�<�c�8i^��]�z�������?,</=�Px�+M��V{�b9�ffǴ�h�KF�ѫ	.�6���+��r���3�`�鳦�%3��
���e�l��n��Elk�kzҿ�x�XQ*i��F��wܐ�f�(T�Ek��s���=cv�I3M3�[�;'�p�[wt���Ȝ�%'8VŘ�#o�N�1pQ���n���[�R"��PU�~�p2���fv� t���}��~�L5�ÍHN�V��U�1ݜ_�f��\��Gݕ~|55�������sd��LS1�+*��e_�����^�����.6ɮ��N��s��v��4(�¸��*�y���ԉ��*�Q� �T!�R�'���I�옞e ��Ө�����[�h�&&j9��o+l�5;ǰ�>�V<wG��t-�uɂ�2�D1��ʐa��Y�K�uudK�B��Hsvu�����s+{ga"�A��e� ��q�wY,w��*t�o��kͱ���
�g��zߟlj�������]\w�"٩+�Zk�X�gk	�sU�ă���,�����L<�-S�Yy��>��	����7�xU�:`��B�(`��wxw�q�zz�
Z<�gP�<Ÿ�9��ۜ��v:W�˻�\�Α�vw�zC�/'(�B�Y.������6����3y�r�p��:��R�u�B�h)�^3��#ܽ}�
�Wr���%�����)���[��*���ꅿL�H�Ι�c��qh��c�#F����;W}��P�� �tH��S<�;����:l2��7~�甘��l��+9�Z�^WL��}ܶ��}�4�zSUv:���ʊ/	��=,��y�<Yɟ/ݝi��D�%�Й�����w\�u朥�`�,j3S��d��q�8�>0
��s�}+}�Dp�E�'�(ڬߜ�*b���:�Mjh������˔O���z,�=�˳�g�m4r�����^����f��M�^u|���v?=����0��{MIc�u��fX@sz�I]?,��Yk7#n�,Yj�2^��X7Sl�N�;�����·��va֖uC�A1'-QQ�fZS�/�/-��j�Că���P�J�_hY-E�x���ص�Uss����P�������r
��,nF����G�[���O�x]��T��z�竀W���dn������
����<<g[����u�B��ow,fi8�����zu/��Lq:F��y����m���:��p��ٖ.��{Np�CGu�j#M:������^�OT���r�W�rc���Ϗ?o��Wڴj/���n�uo�3��&�{��K�k��xxy]�ϑ�I����b�����VtԾJ�<B/��C��EyG�׏�+w������ۺ+����N���۝��$�yF!�%{�7�ؤ�f�zt�;�[���ˇ���X`��݂�^�zЬ����J��5iD��=Z�on�^�[�g���/\9^lW��G�_�'"�ۍ��T����۱v�쳯�n���O��4n�����kp������}�p��+F���s_e�,ޕ}�z�ޤ kP(o,�0)j�G��~=��Ib5�P�)�I]������mNQ��);�j�"��:��ݫ�e.յM���������a��,p��݂��e��sxt�%̾�	[͗���,@0���,CY���=r�i#/�\v��+������fkfk�.�m�:�j��Q��9�^1�xb�t�Rb�Y{��Eȡ�Z�0D�����=3��:�{
=�K�̉P���m��8���=�~ޜO�y��L˺ɳi���� �13�f�x�]��#u��F6�+�s޺�Q6�0t�]`���7��
ة6��g�w���w��_g'k�p�׹�h���³0/v޹bY�7�\5�b��
���gU���KD[ơ�C�l�]p���=��vp�mW��=��_�b�S��+�w�^�]*��Na=�w����9D��d:��.�|=\��� /}�{;�V������v���q����]�`�&�L�՞�J,�r�i��b7W���P���VP�0,��#[4J��L���^Y^��b�ypv�eE^&��N+�by輩"��C��~ݴ�]�&��}��{cB��:�85���a���L��k5*��/E�}����nD�\Q�v���/<2�mOk7O�VZ�ֻ�%�����`�sR�).�'���� �̹�gf����%M[\�\x�ާ�d�o�]��u>V���C���IԽj�˔�� �� E�ĝI)���5�̌So��-��C�#mcS��)C�6;�=_d���{�ݎ�c��^#�N͏r�#
���4i�j���6��zlX����?yt)����瓖�Z9R��]@۵�b����w�n�K���?vf�g�s����3�ZiJ����}�Ό���v��Y�4�ړM߈�c#joq��x|���+���(���p�o5.��Vpn���2w^Լ�5ZB����͑g��;P��e�s�e�����b�6t���;���TI�%Y���vzSo�hָ��&u��WC���;V����w����$�u�N�s_~�c���z�:��s`���e�����[�C"�0o���U�?7o���s�D{��n�z�G���6�G]�� y�y�&�����".�c-���oNg��:WnH��%�g���q�h��+���;�uIo.J+U��lm.�(�k}��Q�רYe_���Ų�zΕ�������R�(�a]	��=~�S�xJ�*7a�i���ة�����y���+�c�k�@[��Ηȷ��^ˣ�>6N][3��KaJ�҈wq����t6��3k	����,̼�cA��!��a�5�NhSmR�*�n��c����}�[��$����Z��՘^��+)q������J�xgE�A�tdw�[��6�.��LN��s�<�:Wo��5^���?qe���K� ��0(\B��}O�8��$���=Z��U������¸�ܾ��S��'L�AG4+�r/��pp�*����\�U�0dB�3u�3CH��V�s�ௗ��̞�z��S�MXPYF�=��>78>���9ϕ��c:v滨��k�}jW��5�P=^/ss�.c�u�����&g1���ijKB�	�vl�:����.�h{�.Gi��5Y
G�gV_6���S�@���X�1�P�+yٮ�Ms]AKH�o��H��s�k�k�C���Y���nkyN����Zʙ��x��O]Z<< �w��
��\:ʄ���VS�X��PwN�n����{�ɦ�����}��7nq��Nz?`�D�����m>�{�2-/v�6{����7ތ>�!ǻko�g�&`��<�t;�4NuV�>J�]W�����θ���w;��e�*��_��/x�Ŏ��穜�(�;�9��X�X��Hsʂ��n��/��D1)s8�-Ng�-SwW�>Y�0%�RY)��q������:��fL�k���d�9Q��n��Z�h\�]ť�������7��Ug���ok�A�}�,T�`�5���/���q��g3%[d�;�a<��z5˴NK��`���j�\�V`0p�9f��{V�H�b"oݞ�$�>���#����3�b�c4e�!H+���;�΀�t6�{ڳ9OK� ت�X�oe�J�vm7:vM筫\�T�����x:�y�5p��6`�c��֞����7����]#���}}I�b�߆q���v�֝~3���\"KwF;���*Eu�u���+���z�Z<�_���#��WY��z��\��Z��5ؙ�E���Ǡ����M������<|-��3���eap�WJlG��S��<34^�n��I�qns�y*�]��&���&���co���P
kM�T/�w�
y-=�p7�ޥG|��u�J��iC�2h�75`�vΎ��9��+[E�U�`�T~0u�CΆs���g�e4�|s��M�]QL��gez�eob7�R~+�Qr*�=����up;�u�5�K/wf�v_�F�*ǡQ~M�3Ƙ�I\�o=����h}S�Vdyt�i�:�Z�����&c�#��܂��ǵ�|l!LrV���K����X^�-�_Xu�GIv��9�/o�nϢ�����Y�4�!J�|%�kյé�uh�f�H�rԺ��K��@﷩�h`9�gl�t���U�
��'C^mq}��caP��X��묜��]��5;����7ZĞ��Y/W���T���ؚ�{�)w1k����b?r��~��
V`]K(	7��=<vS��;�Q���M��w���]e^��{ݏ��t�����GO�]��_\�z����{^̗�����q�1i��{;�N1���Ӡ. �<X�	�����������t����90r������Y:*���b����.��{�n�K�U��??o��ۉ�_��u�y�]�7�v���G�ږ�
�uL�x�5�^��n����vі�e�&mc�a���s�v�b� �o���o+���}��rQ�r�9����3s��������v�{KW��qx.���M�����~y^]ǻc�a���6*�5�x�|v��wy3O��L�ib
�U#���u�z�������4������}vr�Ѐ'��{s^u/a�u��'��_�J7sȊP*�~����;U�2�gg��xJ�Q6ޒj�o��t���Ïkش�������[3�`iQ}�bٺn��b�����"5#�g�����!��kh���<�u����Hhu��</KoMuᶱ�3q�-���Ψ/;�h�H��[��4\����U%uw�a�������N���������w�� ��/ �M��9�Lv�.Xw6�E���<�Z�70��ݜ�95�+R�Ȯ���ͱ��8�F��XP�%�+5��ki�t��Z[[��؀����u���\��Psk���y��n�M�����F��Z��o���ѫ-��:Ћ�k���1��;u(��2�I>����+f!@];��op[�-�Dl�;㥍Q:c���k3o�8L�P���0fጆ!�����t����J��Ѭ�]֡�TbҐY}��f�8벬R���e�!��kzrѺ5m���U�I��\�A´�z���:%3r"�a�A��;N9پS $S�*h	�	Ǝ!)d����Z{$�s0^�0�n����W��GM���
�������#%�9�
���kW^R6�w�K�V���[�a�&�zW"1B�+��S�dwm�a��/k3^m��/(��]p�$é�M��8��a��1�[�jv�,�v�'1Sh���F\w��	hS��&�Hȵ}�5��Hp�|4��� (���q6ng�kO
��cpk�p�Y�]jڲ��T�Q<y+H��UӀ1FĂ��v�]��ٖ냏k��9���Fm�Wd���ݶ���n��gp��%ל*7ǳt���^��+I(�+�{rT�I%F�k�)����v�j��pݵ�IȴA�G&�e�Jͳ}/��X�ʜ� �yq݊�ʳ�r��9k�*]��jGSyf�'E/�9�
�tf���V�[Y�4
wGq87mNSr�1,�Us�9��]B�@�`���-�N�&&��H2��1��9��6]+��r ��Y@wdbZ�56=��{�)#ۊm���k�Ѝ�0�E�OW&�U�bV�=���+\�Lr�m[�Ƌ�x.�&�sW]�����A��i
:׏"��s&	���B��11���Ö�FG��^���B3֠���:7� ��g����CnJ�gt�;5����4�i;1VP��.1�yv�U	x�F�:�x;-J(��=3��A�K=۶h
�=�٢j�i<s��z��Q| %�䧉>;ռ�쏩k��{�[יa��+G(�b���S�&��Ĳ�F���|�:JaRO8�g�4����v�y+z�7��wn`��,���J�_�:A4�Z�Heـ�{�>�k��1�r�c����^����zt�X��N�0�e��u���U�M�̾Wݩ՞��e^��!�P
m*��e��DDXX�֞q]�

���E!��y�};uk��)yIջy._VΑ�B�=�^p�f<ǽÕ�sC{��-�l�ɽ*�ɓ�$��6�8n�偖�ӧݭ�\�s\}��"5���5ܻX�޺�ۏ;�;Ȩ�N2�}ܓw�[�k��snV_-�J[������u���)���2d��1���.�7�|�|���e�N�</��'�vX9�s�'��0���i�Z񈯔���� =��� 3e�E�͘r�� "�������Q���p0�
#�
�>!�$�`�,��J��@&����槵)~��^nm_�FHLN��"�w��(���L}H2 o��2J�I�cDILF�j�0�a�քI-��2�A"<a2κ Q �8�s#ϙ����p�C�������WV��	��$o(�b���$�dJ8b<|/�">!���gؽj"(Ɏ1�U(a$�/�z��#�	2c�4b>=(I&>=��j����|��q�H��<Q�"Hd|cLU]�C?�1�C">"�0g�C `�\I�0�>"%��L�6O��I�G�3G��$��"�#bH���[��zG�3=��ۡ�<@�� 2�"��dxę o�`h��{G�E��$A0Ny�$G�q�D~����0-��u� |`#t���(&,�G�@2�D"0����Q�dl�O�ŨI��{{,z$��� 2<c��Q��P�I1F$�!&W�	(�H���GJ�	Db�P����(�|�I�0<Y��A0���'d3� (�Y��,�����~��|_��Uvv���gL!���D����> 208�4>	0�C1_ e��1��X�D"@����B,���h�����r@IE�I�	t�g�����봷��/v� ��"k�GZ��`e��(�c�@�1Q@�F�@�dA0H%jH�@I���1������8�'9�0(�D6�}��� �0� ˞#﬽�'�g���~Df���� �> I��ȅJ &8��L~ " w�X�&!�B5� ͑�0N�� "#��I0�3�zۊ"B4��[�&�� Z^#���p[~��Ԩ]��s�LG�
"'�����0;�ш���d�`G��L�@2��jc�=�IHY�L���|D"$�H��G� ��7��e� �@$"	h���M �e\�u_���&���D���T��{@�"��l��]zȁށ�J�Q �9t`=���Z��N��S���Տup���X|�:�T29��=�=�O��5�i-n�:�&uY\��s���;��Lכ��1�Y9��aI�fӊ	t��or�c��9ײv��i�.��D2�cB��%`3$w�F$ H�J���?x�"��`D4��04�w�0(�2@��|`&�1d|D#������|���znoۻ3�z�"hGR� �@$30��űf",�T�$#Hfs�1F���� p�Dq V�;#Y��m�Ӝ,�,����|G�P���~1f�!�
!� �1�=�`|�3�#-Ɛ�a��Ƙl�	���]!����@�j�DI�!Nt���>"a�y�}2�m�V��.�F�7��(�֪��� ��G5f���v`a%gLa���q�dE�$�"����@���c���� @w)�1F> ie����I�x��oWvj���>� x��H�h y@&��cH� %�Ę��D�1� �(�Z�� 1B3�x�f� H�Z�"���4� ����戉 J�M��y�Խ�}�ݓ��0LG�Fܸ��|c��, �1ő��&$�H��0(��B,���(���G�0�"O׎"HG5�B(�<p(�D�nO��B*� d�y{�u�S�s^}�o�'�!�<pы��`Q IDi~lU( �4�r���Ś I��ߦ�QD3���I���0�s�Da��H����1񀍑ib(�� ��:`F�嫞���Y�ϵ��f0��f 'f�"�B!�L� $���� '�x��I�,�f#��qFd��"yC"���5S��3�:�2#��y)I��1g}�I��}�k����7z�҈�!��"�1��R@cđf�`cB;�$��B0��"#�,��m�,��@���I�?��(�Z��6`W+ `|~�!RT���Oշ��;'4ߣ�4�0>O�k���,���q�#�O�ɜ=���{�+_z��U��a���VW��5U�:�F|EZ
��ـ}���.����\�Ⱦ����@�]�oLfa8jnS�|���GV���P��:�۬Ў��Í�3�k	��'(�VӒ���\����9WL*F�X�:n2oF]�qN��z�d�.�jD����5=ݮi��?p�������4(*�Ԩ/o�� �CIS�z6��^*��������其�Y[��|vO�ӌ?{njS<�^>��c��XuUv�ίr:/-	k/�oVi��V�·�\����
�I�͌>����Y�i�)'��ஓ�n�8�ۻ��n�YC��G"���j*�e4��pHs�;��u̺�z���.��{��㰋�۳�4�,�[��j��u�wu~�Cټim��:��ezY=]:,(K��zEeb���N�Z�SG�&r�b�Y�S>O!�o9�CZ�1K�6Ňֶ�-�nǄ�<�η( ����ݼ��{�7�.�$c:�����.~"j�$B��/�ZՂ��A�æ��+o�>J���>��Cբ�pˍP������+1u̮���]�i��Cw�7{
� 7��;o� �2b�5�Mޞ@*Q��%q��G!E靋*x�gf��;s���@+zg���,D9k�^1�2��{��)����]���^��N�M�G�� �uw��}0Ve��jε�ʽ�(,jϜ�O�:þ�u���k�������#���h�k�+OV�"����a�c�-b-E��w�f���d4�ֺ�m��#t�Y˻5�;����"� :̭
��/:�����u�Z��_<aƗ,�\�h��ز��TY���?,m��H��}�f��ñ��]�_����6瘶�û����δ���c|u�״���q�P�kĕ
����W��R����%^J���c|����Dǿr�q^w�$�y�!6�3m���m/ 5[��+ֽ^"u_��_r�:%T*�^wa����t��Hq��۱������ 2�,U/c����U���6+^�I����o1���]$u�qR�G�8��ǔ���M����z��R��<��Y��Wٱ��~� �<����U�>�p�;��x�,�*[���Ё��y��ؐQ���>o|���%��a����)FR$ky���tvSċ>;���n��=L�h�G9}������c�Qx]s��^��Ҵ�OڊΞu�������k�Q�(x�z�WTZs{����[���yx�U`�q������{����];�3^��ұF�7iIZ<���.�YMmپ�k�;�qc�|^����������ٛ9&���M$:�O�7���&0��}Aq�t�O]�f8�Ib��*/n�̰(ZН]�x4qN���.Y�����|9zȳ�N�c�K2��.�ǆ�m��L�u��V�����c��.��{Yv(��x�������F!1��$^cH��kʪ�R�5yY� ��[b������Sۛj9�qX՗�@��V(��{���Oi�*~o�	�~M��׻�z=�͎�,�w�K�<-촾פ�዗E�8�P�i��B�e��c�f�oH�r�����<�W+	z A�g�t��=���"�}�}#�\��q����)�!q.�t�k��xe���W��f��W�~bL��[w=�2�5�=��e����ݽ�+^X��uX$y�ReVGޕ�6��I�c� �V��ܽb�'�x���yS�Uݩa�͹B�=,!��|!e�޷���S;B�կZ�	8xp�7�R�>�05ߔ�/�s�[���"�k��7��B?7o7�{6�",��B�>B���'�Y�u8�ǳ�<-�4{� 1eX������E6�K7^�
�rq�;W���f�iۋ�����?"�q�Ǘ�J#��y�T��R�죉�U��༏�V��q�P�1���zP��9t���������{�y��0��ch���`E�aw��z���y��-S���T&�/���v�s�waϷ�����4�qe�=Y+	d5;k��9�VU�߯��n��r�
ڋ�-S���j[��P�'\��ͼ��؄�r�k�9ۨ'o�4h��ƫ+_t�gTϜ�w�mh��zq|����!�ʠU�a�r����<!#�0=L���F�y�/\�R���{���Ƞ�K�H��{��W�ޖ��?;L���α����le�����he�뱾ü��zy��
��ʯ��ᵩ-@�ޑ
�+�y�S���0����%���_� ƣ�t�m������I����
�ZC����
�~��̶��^NM�$�ۺ��,������~��<�^���z�zy�¯b�;���]���T���p�q��*CW��wj�f�⑻)�
����0T{���b�u����>GX��y_��~�˵���Ye����|r�m�!�]��~������k��&%��XO3ӭ2�=��xzx�~7c�$�����<�oW<����v�ڴ c�QA�{�ܢ�'Ƥ���^AÎA1�!R��#�J��u�M��iq�^Fu r�ZYu�}�8�{�;:���C��X�´[��{���8�<i}[�iκ6��S,��v<"ơx
��M2ߙOcLu�ǯ��Ox�s��>#`���*��ж�X[��f��at�R�u��:��v�Ը����$�V<A���XUc:�P���Fo�i^�ݵ���v[z�Lo���J�ný�rɏ{K�Y��u`9�:lnvb�+�{�=~�Y\+��aڬHz���8�`�o����7���K�[���ABzh��Z�Ҵ��joߏg�O
�ZD��_���6�o�mLT��{[��h`��+�ч�<�76���_-	���oo���#֘�P<��1�	��:��&��{U�{۹��s|%gW�־�"�Ǘ,�V�,��O5޿0=�{�����D��}4�5�QyB}�c���'�6�.�����u�*Xo�J�zBO��9XM%O�<�gI����`���I�n�0��nJ�8b{}9C��x�h�ںW��V��e?Xv�k�y�zM5����1Av`���.���N�|h\��hǴsOk��J�q,^mD���-��(�۞di�X7����~k��<(���/�y��t7ү�P�e�\y��W
`�;0p�z��R��x��]�>�p�}���.ؐ���wx�JT曺���y\��K����������um1��9�4�
h���S���w\���ma����`��۾W����B`̞��_hhJ��}oC.�}6�����V�y�l��������o��]1]YWC�jMT9������2Q��w��N&�Z����g4Mv,ץr���}��}��xݜT�G��]�PGH1($Vk�xeZ��!���wê�Uٶ��Q�A�mN���n��t�-WY���|��ݩ�=}t��s��Vu��ȏ+K�Ճ�2�V��D���C���ݼ�|�^|������w����n����n��^�������+}�䎼�2�3�Utޗ�k��^���WaV��{P-��|0D��g�5L�C�/'����$o��e-�ʶ��s^�ܣ5�I�r7��5���p�\(�A����#��oֱ,ʼ�v��Xg^WN���.�hm�֐��Һ1%�_�V���F�8;���8�yϩH��|�[S>g:غ�'b�L��~M?N�]�;Oyfy���ح����܃)�Rw.r%0�����6=Z�9����W{�48f����N���Ż���{?^r��o����΋��P�߻���b�z��D��P���bv���g+R��z*=7��[Iߏ<��|��dz/��+|vMx���	�V���I=�Y��38&Y'�7����Q�H���rF��_V�o��^2�����{pC��@�Sj�NA~��8vgu{�b
�j��P�;=���TP��ڏO�'�g�H/�P|<���o��������2�P�t�x�O2��{��F�N�&�D.)�A����0�Q�'-�W�[K:��,ٱK�w�dq��r��+;���i-S�_Ǜ]�z��ږ6��֛f�\s�]*r�l�[�DK��/�*�k:� ;�j�A�o%���ݵͭq�{o�/*l�&z��@�^�딴�C5j�ίQ��s�]�y�U��[�N̞M��b�C��5�f�$��u�_�sV�g�01��C/��s\����*���*^��R{{�/k������Q@	���sL<�@c�/��D�0}��*��}jG�������{~V�&����z��$_�X�u���oU�����岝�[�[}�͠w�ދ���{�����W��T�R��zK4"�<�o
`�7�5 ޯm�[5<g&�6[�E��w~�0��'�s�z�b��~���$��YѶq�A�ي��!�^�Z�&��E������b�~�޺�i
Bt�>��/8"�)�[�{wWh<����@�E�x�4}icLxL���z�%@P�+�|i��b�p&c��=�Ż����w�����4˖�#��Tk(�}���>�`t�Nԇ�͐nF���
뭯S˃ӡ��{7��?7G}ֳ̲E�H^���L�]��x�Z]�Ǐ���Y��T�v0�ȿ_��/s/F�#t�^yF�o�W �B��]o����2�eE� �s��%S#&o^pŝQW2�G»���:�=A��]�v�%� j�;�%.3d��#sY(���o*<��W\��\u.2�]5Qy͗�5�'�Q�9�os�L�{yY�{��<,w�������g���{��!�J�V�'g+�
���q�y�S���UCv|V�zz�����7��g�~�>���w'8��e��9s�Nz�k�~���l�
�O�g˦�`�Z}������O:�rKw���+����_�6�k��;�e������u~�U��O��Wx��uu-w��z�l�!������ܿU��=��Ki�P'�ҍ����z��v�Q�"K���s��ӻ���Juދ���"�x���7���-l��Y���z�������ˬ��q\9�q���K��~=�AN���{}�|GZ>[�*:_6uy��J�#������O��E�ю
΃�%nt���о���<;���z�T�}�.��\���6���	V_���uk�;O�l����@���f|�X��˒q�j���t�x�g�B�Ή���.�s&xr>^����[�o��NԶ
{`р"z�GAR�U@po�[�D}#��qW��9K�GBt7ll��65���[���\������hޜ��Ӱ�Kp�FU��]D]�5��)� w�,�v���B�bQ�7��^o.�!CE:Mn�"&iӭ�� �/�1��*�s� r����%�[���S�e������\�����ˌ;���m	Kk��Շ�,7�U�u�P��`:�w ;-G�S��X}Bmvi�~�;|����,�&�J�MN�m\�6w�B9O��[ʞ�.g��ʱ�qJ<3��S���_66��a=�"��I�}V]N�L��"�^��]�Lż��,��'�ϰN-L���G����l�c�8Fꅹ;���-��hJ.�4�,;��j��k	\��t��Wm�x��*�+A��;4�}4jP�Z��՞�*���1��N�̺�`涋�خO��wr�tz��R�� FHum�!���C�����n�b%���i,q؝�\�G<�����쭠��n��^�ռg��]�Z��$u�p�j��V8��`�դ&���MK��s1�2ɫ[��������t3)�R�SlE^Z�t��4h6��՚�h�|�A����P�N�`� �P+��d�Y�OT����./:a��wf�7U��H��d�o���,����U��"���w:֤�2­���W׹]5K���U�f`[1wK�vj�\����4�q ]�By0unf�ỏ�>I�����k���iX�x.�9�bgtf�MjF�"Js��{���,��ܼu�BU�o�MaٗL%G���ܺ�|-k\"���i�DD�KCΒ������R4��3��B{���k��|�q�:#��8{a�S�|,hʅ����e0�G�Eq��ت�V�,9u��.�=��?q���)}��ɇwQuڦr�����=�v��X�q,+n�9�:�v]'>aafE�t�`��k�7[t�s���C|B���N׭�pN������	[r�]�6� �۴�1�ړ��{ڐ�A�;��L�e�/������V퍥s�fN������������8�l��f=�3��'�&��n�4��&i�����q�8_^��v����ћ;��CJ���B��nwL��ݮ����Kw��iA�E��wT/O�ҙ5+n�����jf�gT��V�Z�N]�3B`Q꺙*���Ⱥɼ�m<E�5ʲ��0�$쁗�*����x`e�/[���J�&�dYyE�B���Y�բ佴�\���c�s5gu,���{7U=�X@���&��j�]�N��}w�ކ�����T2�M�s<�x������-����5��C9L�S]���8(uc�y `f�w<7"������Ǖr�[E�xx%����t��ҍm��5�^h�巙.ʡ
�u$e����h�rw���@ެM���E[ճ�=��x�����(����9�n�^��Xx���5NR��(���*Y4��Ӻ�t�0�뼽��de��o*��]s梥��_J	_n\�R'�t�Ƕ�bS+Rj�7����]�z�n/�<E?j����jz,�@EV���=������ʿVWo�e�S~~ǉ����fb��@�t�ޱ���p �V<����w��C^:�V�w�9����>�~G�h.�92���׮�3�N��7��X��2��ݦ����:��f�-��}e��V�j$ժY�r��ģ�㖺86���ި��ۗ��^Z���n{�Zip�l�3�|����<'%<������}wҽ�d?:�ܸ#=�2���J>U�筎�wIUcFY�wՖ|Q��=��K�gس��n�%,��~�)DT���[���)3H=�I�r�.�n�ԯ2!^$�i�]~��c�ž�n��������ជ��I�Qn��~lW���|B�#eO�b�Q0��箕w��#�q{�\���d���{%��&[>=�&���u�j����?*�G��n����oI�ڸ=@_������i��^�A��g��=�Ï��=wo������
v�F4-�o������� |EMh�u&��D��E�;n�'1mub5c/���I���?���]`�� ��p�Ď�7*�-O�*�/]v��'#�45L�OL�/��2;��nM�h2�˞�[WHaT8�/{��*��Y�(N��R>��;���Ņ��y�نv)s��:W�O]�Ur�U���*��-T��<=/P�|4�D�=�����^���o������йk�mڷ:���5��}$���׏%��{�H��]%�ײe�;θ+���kǾ�}�������\|3Q��O<��b5�S�Mm�<畓D"��F{��Uv{s�{���}�V�ļ�הK�;���J�U�T�����8v���!M��(�ظ�:{��ns[[��%����Z�����/��z���p���	����N�]/E_/�4'ޕ�����ʂ�T4�ʐu�۔y�|���c]�C�D��>
1^�ѳ��U73n�
z�C�����ｘ�1m��QK>Oyt�*e���mKk�<��Y�$]�?h���q���@W���΍u��Ug-�=)�ݳ�bUй���L��#�<-X6:��J�~.�~*��,����$V5���O5��VxM߸ ��eq�ܿ'`�&.ژn`"z{j���_yF��Tb�Γo�ku�c����^�	���Θ���c��gK�н�f�W��q\�f��ť���.�:-�dJΔ(�V�ѝh�6f˰Qu�|ݹoOj�Oh�ΥY��{dT�8��|HO7+n��G35���u�G��%k���_�E���Ϧ�뻟gY�c�X(�2{9H�@����s��٫�3���sݪ��s�ϡ�n�q��eŶK��嵯��أ�<�=���٬�����d�����	:%vV
�ct�%Y&�: <=r�����>�a��ǵ���G�]�Nz���8)\���W^<,ڮ`�������m����7m�J��|��_�o����z1�ѱw����?zb��>�U^-�T"�*���S�Z�6{��7�|�Q��V|v�Z��B,�L�t]ா^܇��[,*�����u߼�h���/��׮����={H��5^����;�9���䤞ͩ�7���}T����<��������ɰ�/
����SAٞ�����3�&��q����o���DH�GQ�z��^�β��^���u���#�m��<;�q���C��{�n���;�|�s���Zo, ��lQǕ<a0(��ݙ��;���鑼~VV����^�F��Ə��ε�u��K=cZWC/BKz�y�l�J���t��nݰ�qÛ]�e+ �&��aU���w]zW7Qښy�4�Z��c�9h���w������t�]u�yC8得�r�j�c��o��0ejcj���X{��^؈�>\:�W����5�7�3iV�|x���Y�Cw{e5:�_l�&��Ӌԫt�²��`!����++�<��u���w�UC�����K:T��^�9�U��Ѣ��A+|�.�?��<��a��;���'��|7��o��M~��^x�ms;듵���J�K�(��%w��;|=OWR����s}�{^j�K�oʟ��/	Uם/ΐ�z?x�U]���h��V(_�=�(����:��3ԁ�8S��z��5�V���lt;���.�w=N�n���G�5��d1;3��k��<�i
�{e��԰8��4�w��L�W�]u���R���ST{5M/��{woj�>嫼��|$�]"�C��S#����)������\��n+�vtv��`Q��`���,�#`�U�}[����0��9����k�,�9X��x9L��.���Y�*�:�߹Ǡwo�s�~��F*���]}g�,P��7^�%Ͷo`�`\��v'}�r��k�tx�;�g��^� s�կc)Ykë}v6���q�3��Qu��a�+`vsI����}:��2�b��ֺl�4�8rt�,a��(����غy&fp��|�L@fayPv��2/�U*o�V_9�Yӏ;�[7-��N[%�g�qwΘv�6)�w���ώ���>H�l��g��[ۅ��{����v��$�,�������_�*�b�z��t��&9��o��u֚Sb��^�W�T�z�k*��J�P��xb|on���N�}��C��;��Ʈ���[o��7�1s�*Wev@1W�o�=�`1?aOOoo�)9sz��w�����8u{߬C���^��/{6~Z���\������Pͷ#N!�3طo��V��y��]o�j|)�������잋�5���
�ٗ�X�&����CL�׉w���2F��rp�P�t��>��e�/{3^�|�/_�ax�*�x��et�k��������{5x<P�8B��X�$6������3P�LyÕ�+��\ ��o�r^��vz�`��/B��߳��ܴ߯,�z��A�"�`�f�b���%o��?xu�cu�����Q}찅�B|��ۼ�].�1
BRZdG#u�|��}�z���=�W^�����)��Ԗ'ں�z�ٚ�AT�Q��;b��x#��Dg���¬��B/���xz�`��ҧzb����43ɼx]nC�J��{nr�zP��n������ެ���ه��fR:E�����C��,�A����#vo9��q�YOYܢd�霤�V����e�T��1���rs�.���oR3C����Ď>�/�N՗L����n�4ܬ]�{6�e�.�pZI׺tz_%'M��i��#���uʮ3wwY���~�u�<���;B�z��9�t�J=8�t�;�<�����O������`^��r��g* �kυ�1�6yW�E;r���"A��η����wyf^^�Ӿ7�U.��\��(���Փ�����Tix�.���>��s.����Ǔ֧�!�Q���E�洱k��Et��,����}x����`��ToW��2kp�k4߫8�b���%�<ptP��c�R�Uvz����ؿt�5R�e�yu ��ߕN�ǥp�@�:�`�]�+"��(w���U�(���泳���q�\�ԛ�:���ŋ���ќ�#sx����X�A}��Q^T ˧|��g��~��A����^Cs��r����Ql�����>���z�x� �o�he��p�␦�^��^_����1�M����:}�0��I���UV:g���ԅ��2�� ~�D3��[�N����y}����}�[}^ǽ��LTF?%J%�z��Y~����7]^Yw�f	�KPR��!cgF�B��`��Hu�.g�mh�]�J�WmRjwa���}j�
��y�A暺�]g��������R�+��z;2�OMɣC[�8E���wo�NqlQ	j%�x[2wI�"���8��[̢U�,�t*)�V�a��Wt�}9�F��y��i�Vk�y�q�#��D���������wy���>)`	���)<��{��~����/Ͻ�k~S-q��,��������D��q��^U�s1���o�Mp����5_��p5��J�י8p�ɟK��B9�L��1��CӮN�t1�.߆�.���ؾ�i���w����ӜWo�p*l{ ����T��ӣ�ʯ5�ʠ������θh������y����h3�O�*�O,w�E�c��X�-�s�ul+�}M���OO:���Ʈ��'��늽�x�������</ߟ37l *���Ԡk��K����xi�����=�
��f��S��{G]O�����Fz,4M�0�u���V�:��RdQ�����yW�.��:���=Z.����_Q����f��@����W��v�4��m"`���}~#o��R�|���^(�����>��z�h���r��qc}���'�=��C���B�_my#��9Z�����úF ˴���e>���`�o��]i 8{�]��e�t(���^r�*��6F5;*!�u�[P��V�wh���[�%Fp˼��Z�+�(KO{����5|��y��KK�3�tp�7 g�9��[��x]�:�B���P�����ښ@�=��m�G<�{�;®���m=�N�>~�++}=�Z������2�U�s�V�^�̴�S�^T=��!g�x4Azk����v��yr>�03Ij��v���w�A�ړ�ħ�r|'aG_��yO���Zߎˣs���~�~k�ݹ�ȍ��^�^��Vnl ���wAw=���A�{+�&����%�=/�(j0�|�������W�	)���zJ�H2]ң����8��8t���/+��UMìWv�s:GrS�:�l簗�����xU�����ڒ�<5c]��fr4�=bg�8�r���8֎z���{:�2��=���ϻ�����B�Fd�)��PX�;=7�F�m9^�\F㜖U�^��|�%3T'�:�������r=���<���/-����T_OZ��w�e�[�f[��
v�Mq�~��	�=~��y�zy���o����Z>#�����ᇥz������m�]��p.�Ev�u,�W<:�o�-��ح�Z��"Y��o�Q��/ʏ����+�3�����1rڹ����K�K.mc[AtH����
�\���i�ݕ/p��J3X
la�xN�z��ҡ�g���~uw�l"7���u����xtJ��@;���N��=�s��U�u}g��PQُ8�g}��<8Z
���+0�e}PfE���^�Z�Փo눃v���U�µY]u��[�=��ps^���g�#��Lq�f ��&��8��=KO�iӫ�ׅj๎2B#m��O�&=��h�x��nke�����]�8�ɼeJ��M}z��xn���������3y���)Y�SL7#Ɲ�<��
��RCY� ���/R�W�BºN�%�B�Y*v����"GW5�){$��qp�Z��{\�܀�_V2i�ig?{T*̫��������}��C���o̯=�OyKO�rjY�7�_6�G՝j�w�V�LFI���~X��JsY��5^]��Y�1m�T��E罛8�=�d������X���ʾ��1�@�m��ٞ���}F����Y�7�a��Ů�������ow��{)m,F��[�䠷+��l���?K���G�>��_g{n��&򒧮/�������WZ�
�����/@��/ݝ힫�݉6X/�b�����#�:�Dy��7��.��S8�k�_X6��B����2����fg�����M�;��9o��+�"ƭ
&i�TFԘŊsEu�K���MoּdL�Vm@	t��5nIj��\���WAh�X��w,"�:��F!�e\z���A��]� �E���mowC}Y{q{�)9j�ҍ,FW����1�jCFy�}K�(�gm�=�K�3Ɵ��Z�xMWj�p�L�����='���^f�B~~+�x	,}�oootg��U�g�{�]���<7�:jEW�?
[v��	�Ol��~�x��VMH�`��H��R�Gc�$e�*{ҏt�C�qF�$�2�F�S!����(���{��]Wx]��輯���;�����s�nn n�X��{�s��q�孤�<�=|�ʆv�7�(��뺿qi�5�b������]`�>/��z3��o_����2�����g����Vb����
'�Of�!��<��U���	�<��d��M\��O@ >S�
�ڂ�w�v�J�[~�p�]>�}��
�^�_p�s~GOv�}~Z*��+�0�.��i��Ut����N�����9Ϸļ���[���'��S6�߸�{��H�Gg��R��������I����ь�{�XӾP̅]�U&3��N��ww��`{ՖC���^����:��Z��p�c���[/53����_�w�2a��q�,���[�(r=�^fF�r�i�:[kY(���X���K�]�7���8��nd(dzE��G���̓:K]�o.5��������6��S��cN��}F��}�'�c�q[��ڪ4�^�p18��Q�!Df�cc&&l�O���`M��ۺ5�-����a�Gh$,2��jrh�'JY�A[R�ڶ�V-YW�V�hu��j�٤8�M�sK�U��e��l/��͊�̢�;mf6�����w��I�����i`����s�q*�]Fn�����l.A��w�/�����t��QH�:��Z㲋����}��6�7B�v�[�$7V�8���]d��G\�mb1�\�C���v�#�YX��ZأNb�|ݍm��n;9ٶ�����j�r��7eHƱ�{����<���`��`�7���]7~�䷅�z��&�_ �١�_l�:���&�R��]�YQ-��-�0N⬗��,��5qa��K���^�K�����3Xo���Kz4�&��Q�p��`���h�����F�c]i9��Dm�gKߊ�w$K���J���NG:=h���,Ńy�s�u�`|u
���b6k.�:V�kٻc��ľ���E�����6�>�"[ڦ�VĮ��h8FŔ��f�;�)Y]��.r�;��V�S���eb�oS��ľ�mm�f�"���R�c{LJ]鮸�[yL�钌 7�k�]����ɳ	��p�=�t@��`��X]Z�ȫ����2�s�m�u��rL6z�W.��<��,Ŵ�nZ7Cz���*���tSa�+����'j����oBvwq<qv�I];i�a�����4NX#r's�5���݇(�Vу[�ҵ�n[��`N�t�w9�_����_v���E�cwUL��ۻN��"<�.o7Ɖ3J��|��X�fvYJ��܈)�}k�۸6����`P	;��,#��ʾ`�uce�z7�u���Vs�Dn�R����}�fm��9V/�k`B�s��t��ƌn�Rҷ��4�V���kG;�E�Nb�u���]�;�=O"�BU�@��긱����D�
e,]���]2���@�P�pE��Q���ؗ�N�u�z��z�q_	������=�;�d肷�'��W�;�5��g�q=�NX8��o�Gq���uw�a�ĩ"C�ݮ��:�ۤu�e������o�ڱj�![Mg���\p9b��6$���c�^Ѹ���eW��� ۬�qͩ�����I%���c��V��]s)�͌_b6������:����B��W.@��@�饃�r�P�5�@v���a�n���6�]!VN#�K��:��6iX��+�1-wY��%k�
mغw�N�g5��N�{����*l��q<���� �Ǉ3�!N�ȠD��t��ŹB�\�`xң)��]S컮A�;;[�]3{�9�:3�;�y�w��o��Nv��6�|��૴�c�.��eM�kF���}��DV���֮֯���z���5�p�w�bJ���ow2gs��bT�Ǔ�_y����B+�]��F'����Z��I��ڈ��1t&#�Y>��ơ�<Қ�/{�����|�yע=����ϧw���%S|���^>��*! �\T��&�7�g����ȉ������9m>~��֝�w+J��>�Q��C�����g����! ⷴc��T<��T���w ���;�G�T�gy	�:>��:;�&�o�0_I�f�Խڏ�Y�W�PBR��׶��&��¬���S��_��X<��n�^�y����z}�s6�{xW_�zs�A�U/��G({
�V�w������F�u�߫s��%����+"���}�vt�C2Z��y���a�8�蟚��}Lǜ�f��}vؠ0=�l�WY�r+�W��V�3��^���Hh�x�S�����r��`�������5\���f[w�D��<����2��get9�}B��HN��?Wv�.�x`��_S>�jv:�nɞ��̿��g�=�V�T����#��sz�����L�~�i���o�5���(����U;�$��@KkV
!r�p�;��B!��
q�f֎�wn�l8«:9���ׁ������k�EZG.ql<��koEa��1b��,a��ft�(3�ta{�����qԗٛ��u\NNi�p\�'�(�4��0H,t��h�r��eP�3�V��9�>V��}3�-�J׺�n;�W���ǮY���׫ۓ����wf�ߤȵ[���E�G[1�j�>�F����aq�������+}�*��F�V�9�����o܃;Q����}+޾�����u�����9��m��;H�P���g�nXnV��b���B∺��=}��4&��!^�|`��W�<;���]�@�B�o�Ծ�T� ��*��6G�$�s���е�\9�,|5��^�==&�{nmއ=X�wwJ�j�;R�9�ݺ8�i��"[��hr��ۣ$�!����֮���~���}7��坴�}X�Ӭ~o�%ݛ��J���<u�����-X�:�*�V���t�@3޴����������ϧ���}\�}�C/=���ȅk�>^7V�&6��[��Mz�ޫ�!\=�O�{���=7���o�c��N�{�%{.�#�p~0�n}Ϯݑ�<���V���k|G.t��|yN]��=!u�stVN�*����p��,��Q�����n	�K��d[�Mv�h06[ZYub0,����$�-��`�:�-�!4��g�l!96����z�mҙԑ���9�e��=@�GWB+{2�;{}0L{w�cvG=��SJ��$?V���8)�&:�RK�ih�Y����j�����Ǜ��VN�5�`��%8_�hW���tP�5+��W�W5�~��#x��M� {X�~r�Y��]�w}c�x�m��r����A_�z'���5�B���߽P�9�������P7��Q6�|��龭S-�o�,Uᝥ�c���8�]I��e�����w������fr�H�.ޞ�;�i6x���*���¥�(ͭu��R
�0�+̢W��4>�z�0<����sE�z�L��sWW��V���V󏠉]Y�`�q�d��������~�KzN����K�s��P��L�f����}�ѧ�/����\�A�H�}�@E�̭�ݯ>��Zǖ�P�J�\�.)_��˄'ك�*Â&���=��J�,ս��ή��s�I�4=�?:c�]z�c/Q+!qrï�}Q��!����#����W�;����ļ�#��['T��5y:�l过������{�^p4���er��q{^��xM�=԰�G��ɛ�37{�b��U-3�N��L���iV�*��W�`��S��;�_�[�޾P����sX���R��l��t�%Z�c+,�C)��ZMo7����=粜T��48M9��*.�J�:��<����Z�΀_Up�5[��ع���>��ڏ�x��;�ݯWHo�{z�z�-z�������������	;۔�.~{�!��Ǩ�������h�����	�}����G�f׈�IoT�v���^���^�fh��%�g�b��z}ow���Z(o{.8Ȧ�N.�D�� ��Ҵ��C6$�̉�^�蒊~�;�nsu1����.Oy�	>7�5u���W0q%�m�"=�s_����Ms�|�MIM�6��^G����e��*�Z|e>#��D�q��s�jU��u;�=:6\J�~��o˷բ( �J�����Ξ�2}y��ҷݥx������*�ZVY�Y����b�$A?hG��f)������M�8틆�^f{�QTpw�zo�ީg�Σ�-Hm����@I���{!W�eu�S�7D��^�� N�Tu%X���7�:���2�_���go���C�����,o{�A��k��c��HU�&�5��U�0�n�M��Mvs6=2��pzS���A�\<�[���B�����A*j��чX��]x`��bj���R���ʥ�S�M��fHjn���\�5kӨ�t{o9u�j鴵+r�gW)&��uQ�p=J�l=���{��v���b��lv�N|�K]�I�Q��$��s� + J��9�0::����=i�گYo���Ľk)�7��j�{�c"�Ԯ3�z���j�5^ޞ���O�����n�ۑ�)D���Y����E��/P 8=�| l}�\�5���!v�{Պ���x{�� 9dq�Y"��kKI�A;Ƃ���5�nǑӼ�c���Ɨg#��
��P`_��:dJ��[� j����H�wX���AWM�ϥt׊U�3��'I�/s��a;{o_�fץ�M�?\s�˗>�)|Ϻ��	u	8���S����*W�#x���ieK�;����gn�/0޵K�����!37v�z������g�X:��y�2>^Uer {�~ՃoG�:¬w��Dľ���r�+�1T��O�nbdu��S�A<��oBN��f�)������ثZ�V�Aoi^t��WtB��|-[�B���!�:����]l��-�ij���Ѻ��)��U"צN�N<J�y{�&x�4��K��o����ę���ז�U���C��n�>�t֖�����c�^	^|����~�H���St�c�<hb�E����z�ؖX�R��3Vާ*�w�/��ir9Ԕ#d  7l�;���Н���Y�Y9��Vjbw�ǟ,w %v	\k��}φ�$�뒩f��6�+�lV�7oVc�%���)�X�����N��ܯ{����W2���w����r�bߐ�����KG�}�eԽ�xivk��w���<#�N���A����z�� ^Uu�2y���CG�x��o��m"���Ď9'�x򠧶�4��ޥ�)��a�>;x�.�Z�����r��[����}�j��k;zg���::��kg�v��o��;�ؗ��|c�D�[�ލ߰��"�#�0�ں�-_���a����=��U���Qdt%���\S>a����>����՛�;�f~=à�;�>�����{Ƴ�*m���u� #L��ʕӅr�3�ϵ�;�ŜQ��j�l�3���u��Z#��'Qw4�إg�u-�Y|:]6������������n������z�_�0�x�M���׷�,աl�^�Q��K_����׾/(���gZ��Ə+��u�h��W% �O5�xǦȓk�{��'�R2@ty�8}�x�{bX����x�������H;�4R��'��>ɾ�-^�RnΝ 8f-��nIeև=�qt8�맘Ö���u�l�E����W2�}�Bu��۴���,sl>}�Xn=j�d�����:��MAY�<�]�T8̽�7L;wP�$78!\Uk��{q�5�mvb�(�N��!o���n�Es���-ܛ�
}��.Y轋�˞qֶ{�R4C�(O��5'�lR���h��D��\��<�MT2T=睋��\�s`��W޼�\�=�9��W���ۜ���[.�R�h;� ��õw�N�W�uefi9Ιe/��� ��b��5~��.�<���`��Jć}}iU��/+5T>��C�չ&߻�&���-MDڥqh�l,���	R�������y�"��_DƷ��}�u��y_^b�8d�k��f�W���UףC�={��i���WxV�@�ː��ms��m�*�����{ �/`~�p{�+��]n�������j��㡉�w���y��O�An�W1«��U|6�Q�2�*t�8�<K�:%�*^���0�}���짲V{�{)d�s�u��t:P��g=]͋!�b�����:�&����u�|���A������oV,��ᚶ����n�'R���U/���Rjr�H�g����P�=0�W���Jq�X�hs���ј�#w�cd�c9i�%�Z/v��p�����:�t�w����r�y$xCֻ�B�\�63i��ʽ�9F'y�]����r�V��v�8tk�B˳٣:�v)����,u� e����*��K�:g�FkV�>)��'3��ճ�P����w׳��O_xZS/[���]�Uu7���Xpl���uLU.I�tO��gg6A��u���f{�c�,�r��@r,�	�s?Dw_����y1T�p�U���;��s�ja�y��2��_wbn�U�=sB���r��f�j.�?WS#:ep������hml��u\Zw��p��7�^�K���4zVX��F߈����s.q��M�t�½�Of�{�.$MA�S�Wv���خ�1�ɲ�Y[��O�D u��o)����o�Q�r��ȩ�mr�d_~A{uĶK���K���m��3���P}q�>��6��{�S�S����v�]���7�+�zr������T�D�N���+���ڳ�`��n�qj�,����W�	�1'7 �[>�t)�����B��׫vs�U�Z��7�sC������a�j*�#���%}��El�A�68{FΓo�4���~W)W����;}�Īo�V^�C�;,��.}��뻢uI���.�n��1A��U����������r�'\�(�����[Z��e�W���[]S�vMd_
��Њg���SȈ��z�X4챿��S������H�%�`]yge��p��n�!.�Lݝ����ڍ^g;�u4�T�c+,+5J���-�G��N�9g����һ��"J#�٠t��#�ˊ�%��EY�K2\"�����;�� �zʫ�OUP�5�H�H����=ac��\�0��)"#[�=�0�3"�F{�&�/$��7T�m�,�^�x�\xxi��q�Z�����fm��3�1���Ye��\1�=4=m�6j�K̪�Y[39�٘o��d���5��a���rܹ�>14�Iœ�zܼ�f�Q��o��B����J4��J0Nߎœ��T�x��U�mSa�gq��@r�u9�a�� ���ly�\6A�So�gЕr��/U`z��qF��_𸉊Y�Nn�bNo��Ϣ�7cj#���O���H/���~"�:mzݓ�����v�����T�n����w�c�E�o�b%@x�����N�yx��U�3z|{�獍~��h|�����j���n���t�o�bDZ*w�9�^��#�vGv}H�2���;G�����2������ѷ�"3ͨ��Z���F2818�:�ǝ���~z�=q7�:�������L��}��L!96���0hj�n�;��'��*��f�<[Tö�a�/�1/C�J�3�܄ڃ羨�5�dQo&wr;C|�O�x�yR�<$�3>���0���{�22#��H<�g\<G>3/Nw����&����[5�e�"���\Y���1����p���t�[����W˫��30\S�����U��M��q8�����KH��-�n�u���nݦ.
�Xm��*�.�3�v9�����R�2�:ͦ�E��ວ	֨��;�WT���c����3Q���g�Җ74��*L�EsY�3Ġ��7*��J��ٙ۵{��xi��T8#l�����=F�C�/�f�E����q������S����4�L��ˈ���.u<�{���{L�<�*Ȁ]�wU~��P4ELs��g�2Ċ�lN��� T��/3�r�5Y�\�w*��-DB1I�bCg��[��L�-� #�;���X���.6�H�Oo�;}"��W�L��b)����:gW�z��}��b���}��wn���LvK�a2�677'��A̘�V#�|��a�Yb#3w1��s��v�]]73[K����Ņ��
�������n�琽��'j�������&���o.dW7ƽ�
�����f)�^����uޅ��^���ud��lZE?p6m9�P\S��t+*,/�VV�rg,�Ӑ��[��I����$G��"����c!�`7�|f%β�8��۪/XooF�r����"��s�o����^�&��讞�w���^S�7���%�i��*�N?)��^~؈��P��z�?&vx�˿e
���S{�D_��$�ٟE����QĹ���z���&��s�C���j�Jem#����:Ľ�S�lX�y�t�u�%q�M��^V�v+����;�-A�����!�E$�TCiЧ�ӹ�U���,rʏHp�qXNui�q�Y&WM�8ċ1!��P��±޷s��d�VtX���s
z��LnϢ�N��tݮ'��V�i+1(*fYYLi�"�y��X�SUN��k���Q;��fK�e�ܤł«QP]X�j�L7�n����řu���o8�����Ϭ��mM���lLm--m˴�n���=ӱ�;q��v��;��o7d���w������cA�m'���L�7n嗣�� }l�������SǛSA�#�M�[��y���ࡣ��Ӻ�z�=ᵜ�����6ڬ�gbR���O���+	����e�\%Ԧ���b���-��.�]9ҧ�؅L�Ϛݔs��]��3a�WKEH��{twr�сr]H-�CQ��o��M���f�w�$�c�7�С�gn��Ď�B�c�$��],ès��K�O��RhP�!JP����m�-��7��s$�9u����^�Y�M�9���1Q4��n�h�ӻkA��yu��4��Lh+�pY�p;�4���f�T㘡�̅���pN�/�פ�����.-&����nN	q9Q����Z�[�aUʥ=�T��W�.����Q�����N��ч1`�掎k ��Iݗotl���܊ 7v�B�;��#�%n����L
��.��+�3�ZuG�c��n�VU��9P4�u�
Tl�C�e<��U�tu
�pΰyu[۝(-��!�5�k��e3��I���c[�a�6�{[L��j�fb�R���.3��d�Q�O�A������*T(s��܂�������� l���UX#y�ҜU8m���9I*=��;V�gN���VZD���,5�"�[5	��^�s��*��NB�����g8t>=A[�vSQ62��x�yͥC�0�`�Em���VVS�`�]\ͣ �v��ͱ�v˺yu4�r �oV,*�ˢ��E��̰C�oo9_�T��Q�����$��6Z�;"A���VJ�̎gI;a�/�W��5�L�5�GI�w�;����)t�n�q��]�J�N|�jﮂ��v#C���ԯ��X4objG���]�+��@��k��3��V'f��i(M1�ó��`Ǡln��������G�g�b��N�Ŧ����\��k��[�r��_�{]���}�t�����Fjs�P-d?���J�\٫��!SgF�XP_Y1d����s�=���7�� �k���fթ3�B��_`Y6�7��e,�ns�U֜���Ζ�=�AR�M�+�yi��v!�<�`glw���@o���Kt��� :����>y�p���<����Lz���#w3��+{[YJ]n붩���>�c�N:8��+͕����Чxm�6��qG��Z�����fl�]P�e�U��W[�3W�E>72���}{��{�һ�_%�f}�ö�����g��&ׄUJ���ET��{�� ��=�j��ޭ�c�4��Ѫ�<k~��I�x#�^x{�ّ�)z��0gPQ���.��{�(#=d���j�̈�s��ci�L>
�yU=�qu���Ե#�8����W�íK��ʠ�{k&�?��<jz$9�����9����謬���M}-n
��\�ہ������Grg4��YB��h�.���3��Н�J�x!�^]D��/*�ywU��o��z�i:�껹��ѻH1��㘐��e0{}ns��+Ŗ[�Ǿ�c��^�����t��N�C�������y;���6�&'���S�+���f�%dM`�P���EӰN��+�bߣ����q��5���B2�rwM]�;w�7�@�����z�son�����L�ÿ�#
T9#Ԭ���c�b[�'t�A� u���'��o�gz��/��c�g�@?�V(w~o'F���\�G���o;�|?_C�K]뱛>ע��V�ݶ�z�ė¬ޘB��^F�]��J0~��X�b!8�q!�=?s,�he���ç��(��96��\�Â,G.�փ\��/6Vf<SA��
�"�Aqa�vA̛͑k�RV�ݮ��!��ie���z,8��J�hDf��k�\r�8���v�Ww��J\zn,���鹴]���x��L�Q �:��@�t��{{[A��-1�vd]�5B��o!�F�w�)��߁���"Y�@����S5���hC���g�+�����1�����\�u7Y�n;z�z5ts�w��0�����Q�E^���˜5#fw��E` �E�D|_��;�t��ҡr{�J�wѯ�xEzG4">-3=>��B����&��߬�u�e܁�v�D�1��=w~K1�ٵ���7�ېD�A��:���k�1p� �fK��U��G:����}bw9�1�n��GV5�@^Q��m�c=�MtB�f���B�T��)h�|2�<]�;t�[��n���s^���]O�_�@q~�L�en@��/;֩�{T'��9ʶ��B�Xm���y�*ۼb��[/t�����[��{@d͉;�d{�vν}��`�*�`V�ߒ��=-�~�� ��J�\����Vk4�������;2zv��K���_���r���X��j�����D�Wm^`n��O�Rۚ���x�"<x
.�k�3w7������p�`�;�Q�N[}������t���Hu�[�E���z#|;Ģ�4�n�FKqR�,R�ڪ�2i@J�`s�����TuML�D�Vճ9�,����2���Ғ�YX(d��&�
��6jVY�YӑxqO�aՂڜu�߆6�^�q�ʌn ���<N�2��q҇&�@�ޥI�>F�7�6�fT�J�k�.-���5��)��q{������
$9��ovA��Vs�Su�Ny}��/��8=��UN��[OF�T���9y��p�g�b|���;'\�6&�C��
�1�]�����[��>ᣤX{�(�Z��t���FU�}�uӾ�0B�¹:� �=�Gʃ��QwnF�ɼpg�Ӱ�$�FÓH��6Qr� /C�p�p���B�&�%�;��{t\nen�"�s
��vA�n����f�Lk[��B[�aߊ��r2\��KǴ�5�Ռ�uK�,�G���/~뚚��#R�k���,K�f����&�	�;�"���dg�.�	�xLf���](���o�ƶ3l����؇y��㚖�[�S�*�y��na���ۅ�xY�(a�� .xf�}}G�d�:3K�D�Kܲ�~ި{�>jz�i
�}���#~�Z�8�!o��
�����L�gr:�*�G��@���������7(M���+�z�hwD�w�m:�}�,x��o:�����׀mvp彑��C����Z�9}۷5џ|$Wΰ�T� ��~ax
�+���<'HgPg!/:�z< ˮܕ���sQg&����w
\�����˩�6��鐦^D�r��v4r9D�>2��{��ٞ��G�k-Q�j�)�ʼ��
�@��Л�~/sZ�k8�͸T��t�D�T��+9�� �[U���*Iq�P��I���Xn�u����������Y�k4ǡl=��1�u�}6o^���A	�Wq`=�L�} ���u�qV��sGNn�vHvK��"����o���7R�D�=s:pw�đ�Jf�/t�T�Y�7a`�S(���^�f�R�oj.�'wu?p��<3���@b�1M�C ��fW�'De��a�C|m�خ��3�t���.�}:a���@Y��k�X!��3QEwm��q;⧟5���Fئ�]_��dj�vI�yt�����0cz7V��#\\��z����\Kp};�&�u�������IU�:�ι�J��kZ����s��\H�͸��	Όg=P����^���N+�v*�}�}.��
���(�Y�Ř�Dl\g����f�x�~������C ��S7y�e�nm�����xAy��Z��|��t8���o�>n_������������'��Fa�
ݣ�Dxϩ_uZ�u
 [���5AV�|j���ݗ��w�����.k�gK��0G5OfP�}��t癙�!Զ6N���7۳����n�O �G�7?��������+�n�q�q2�̾d�����+���z6T�K��b����x&�@/e�ʹ>�uw.OKyrN��7¶آC�T,�A��K�>�:���"|�w�dx.
nh� }W��O֏��}A��PR��<JC;
�����#��1+;���N�D�̱��t\�38d��|�Y�+�Ã%�ۤ;L�M���k���,��2�5���!���XH7�T{&�]�)vQ������*������L���\�G��.;��/D�>=|�}�EX����:SC$럺��tvڷU=��d���	��������mI�w�_+���o�mJZ�����R'�N1�se�=xI�<�}�g�2��Z�Sw+�����n/�|✯�[Ep��������]6}j�������0����ޜF���'e�T'&�c�/O�D����y?q�W�-ULxVI�y_}ً����W�O���F��ߣ����/zAT�?cY�.�¾�/-爈A٭᧳Ǭ�d�ϵl���<���馡��_y������v~媳,8�%X��"Qa�)��|O�Z݊����rx�UA�����Oc�B�̣�L��hF�fG?di��Iھ3 �g�g���O<�G1Oܢ��K��s�"��]�������䛻�Y%	񀮤�<F��e�u
���確W���{/8\k�|.�LUx}��K�:o9w-᾿�G��f���I
C��I/��ŭ�>��V��o��ިEzc޾��z=阥��m�g�j��U����ibb=ј����6�[;��	[����JQ���fE4V>�}�M�|����R����Ը:�:�U�����m�3��s���|��L�8H)6�C7�n����U���+v����N�T����؊���1y���U
H!�X����*��+���]8����D��F�S��.lv�������c���M�.L:�Yvǝmv]V��ƨ�q7������s0}�[�T�ٝ�̌K(0�Є��n2y�U���{9w����wT@w�f�����&��J�Õ��fo5�g�M(ͅl�LW]�bz#荀��5���]frضrH����#�Ή�к�O���L{Eyos�@Т�9��K7��n�Ij����}�F�ðX3�<K�Î�V���u�ˡh�~�B1�5�����@�O�W�v�=v����p�I��d��=�N��۬��`w3��m�kVt�
�y9C��K�9&~o��E_��	�����to��ӱ�J殽
�1,�U�qe{�t{����L�l��Z��`��@t5�/ ���/ߚs���D�t;�Wn�� �����I�0����s�����3.e���!�VE�&V��oڸ�;y������/�v��6>����i;�u�H�\?M�G�]vl��W���W:�p��� ���X��������};�����m^������j):�������}�yY�_�d{&`�������HtQ+^ kG���3BaV���W%����>�~�Q��=��:��?k�`K�g/9�q�a]�;�i��.zz���:�rYD0��-]���â����J���cb��]n�>݂��Ŵ��dgs�7�v�j���̱oL��+��q;j����7�`���
2�v��uh��޾���F�#��{���܋�>����I�����*�Q���$揮��˩��=V�:��X�,�HW��j*)���������x��*ۘn�5*�����y�����ٟ�T9��{q�p��ɟ����C�|�f-;���u�ts�ٯ�%s|�E6��TRI�<�؁��LE���M5D�Ҳp�ݘ�c��ݢ5�x޲�[�N��M�N�d�y�]3Kb��O��+ʸ,tK�^��T|�UL�ڞ#k8�~��J�����	�H�	���Q3��MF)�9�������5��b� �t���z	��24wvT%�3u�:L����F��W;�	�no`sr��6�@�΢�}��̺�޾�=;���y���:1\I���@Њli�8��˹�aDS�C3(w�z��:�b4�_�=���{U�\mlB��5�pf�fS��پrVN��X�/j(�{G��0�wѷB]���^���W��\<��=�уQ��&墠t���3����wS���ҭ��� �Oz;�ֻ��,D�f��8 Y�\���C��y����Ϋ��-��D���t�թvF��i�h��!�yeNGHH>��BRM��u�"�V�$ֻ7 ����4�X��t}�_p*��PX2)Z5�0e�[o��B���sռn�E���{�M��:��}�ăb�Y93��kA�J+���ۃmk7Y�MG�����s��(>�)߽�e��S�b�=�,��m����q1�&-v�"��,�S{Xx���xw�����7::��Rg��"l��=�+���l�M=�&HU(���B�Xf�b�hky��w���l�c�s�cT������5���ʚ��0��$-��t��^����{�e4<�-o�l��n~Ds[�1�[��ʔ9��R��TH���SЮ�ɀ�V�"�L=���}�w�˱֭|%8���Vy<T��F��������읎;����%[�1*�Rwj�ݺ��� L��//s3��&w%�6�ь*%.�}�p�et��~��TS����P�%"���Q���ҥ��6<�'�q��+zk������h�ɺ����e���9�Yi���d�5<������vb@P؍���|
�����/��Y���j���<'���aΞ�:wO�8����&�{_Sw2T�V��Mr��{5ly�ݭ��E�ܩ��g�d���pm�j��8K�g���ῧ&���0_vf���$���V��)y���d��LY�^I�M���¤T�݆Zȸj�@��zr���<foa[3��=ᆝ��5���t��h���C��G����MJ��;��ه�m}�
��;64�Nu:�dI��B��{tau�]o�m����X�1���;}�T��3�.�u�{}7����@��!e$���AZ��l�H��g" }�d
X��6st�H�j{X�V�T�b٤½�Ӹ���" ���_w�u�=�D6ZU<'nr�O�wa���q�Q1=:�FL�rQ��foNp Y��\���צ�'�~��3Emg��Z��/�W[VUH���S��|���H����rwj#*��x"��9ض��z�2�냭XX��i�~*�ʢ灸��3or��������;�K�S.�s��78�؅����g�)26̠2+
f�)ɚ�L�dU'7�������;��R�n�K������������"�Q����ʩ ���q$)�>���z+�U1�}Lh�Ļ�����*��>w*��ջG�^<:=+�X� �U��U��&)���y�F�|DA�/���|'�:���]�oX��a�t�o����&P�n<jeK�+]���׊'�f�,c7�=���nhC�����^׹��ݗ�
A�${�c S�zV����d��<�ܜ���v\���3F�7=;
�'״D.����3�h���w�բe���A}-�R���ZgTt��q#U<yXЄȭg�9WL��k�������26�H��nZʽz ��*�hյׁ�)6��{'<`LH�;F�l�b��H��N�a1�:�M�7wl�?o6Ὕ&a�$C<�� ��ܶ�M�D�����8�� ��)�g�2	�ݓo����W�W�Y52�r��٪������oj#�cb����|]��e-����¦�F��W�ͱ��os��%UM)U�s.���r#�[�(�Y-��Լq݃����/Vǲޭ�>��_W�[�dg�ǵ�Y�f1B�ə�`>1g�����M�m��y>���Bf^չ�۝��ݑ�(���]�:����u+FƼ����|傟��u�y%��������+��!�(ڎ���S&|��)�q:��]�6��=¡�s�e�'�K���j����;p��ϺŪ���eP}�Դ	:"l��#��nf��8�}����&lHU9r��/��v�u�o�Ư95ջ=}��~U��=�9�HuL8_��*/²�L��8^˨�*9;��d�T؎�40�n�F»g�wֺGn���e��]a�C��+0'����H��}=Aq���h8�V�Χ׭x������;�X�3�P����X�qJ�ݗp �~��7T��t�F�'��7�P�}�����;�s�>�˷^jMDzq
p���}2���� �,_��t�:%�Y�;X7�|N���F��c*gY64��pW=��[I֚T�ۣ�6@�)�,��8k*`���ܰM����CU�?1��t-��T�r�����u���s��av��۫y�`����W1H�}��P�ld3�Ⱥ����;�7��d�Tɒ�:�z�tھ�\D[<:��R�K5+��6��r����N�����@����$3j�¦�:�������<�̺ZVV��{Z�{ڪ�]��Z����U-��U��K�V>V7��ضgi�*q������B��R�DX�QS]��i&��I�r]G�V-t�;�5EHXR�����KONW��[�(�����`��4�i���Ƭ
@�ބ^�T�q��ubΑ�kp�Z�*���Y�܁ڷ�u �X[�4y��c��p\7����h:�tl]]���#`:�,���۵Y���0�����i�WA�Խ�w����mەDw.�����.��܉�{j��)S��+�Y�N��5ns�.�Q��h�3%ĥ7ٝ�a�q�d�m�m�Ht��I�:���f���N�p�'�v�[}$�����3N�!;��_�Q:_@������P��ړ5����W��NMl���3��	-\�Ý�� �f,�]Ѥ�U�e���t�}8.�p[x��[g�e9V�f�>4�O^G�S���`�5;�_
��[hv_ۻυn��.�.="���_+r�Q~u�[u������tX7η5'ZΧ��Bu��*���#<&c�H�%ʹ�uq�8L�Et�jt��E�{}4�XN���J���՗��������ȳ�Zw����ޜ]
��>��F����U��꛳�t�tx�hJ�00u:�ض�k_Z��˒���b�ݗ!]�����s���:�j�5�ݱ��v��w%�25�]H��:;M�N�k�V����v�\Rjj�A����v����E��ᒞ,q�B�6�*���
��A�V�}/&��1��4��"��%���9�]��)t�t�ZV^[f��H<��ՃS+mǜ%!��������Nbv���V��ot�"TI�X�7�<����� n��=�B\�j���"l���2��P��'��M(�@kv]\T�Ec�����������~��U66v�Q<�c���vj�z�5P
�� =ۍ�b�3n�=]�'�+6��	&s.+�Ew׭v�#��<�D!.�ge�yZ�����kR�t��t�J�6r�7��!��Dء��r�l*R:���;y[ewKUi{yսNA�]�YR�%���hwͫRӵ �䘋�2U���ĕ�`Cɣ�h�����O:=�zu���<��]r���[F�Jܾ�u�JPf9F&��x�g6-�k��~�Εzm�4������hfc�<7)��m�yH���xs�5zܻl[}�j:8(�x˵J^�n^H��I%7\�٢^�y�I�q>�2�H�la����_GR��Z5n�E��gj���X,s�.B���c�*�f�3h��rg%wB�y�BZ�b��1ܝ�����髫���YݏwW4oc�'E ��fb�~~H���n�J:����盙�^���;�;%��w�_V3�k�yճO�%sƼ�c5}�ױ�9 5~��z3�"�Or�Y��B�qâ�d��f\n����ج����ع�K��Fw�S�Xrˮ�7zeפC�r���t��]���+��_�=�e��<�V�^���W��vl�k�<����B�Mb�]ML���k���SЍ�;w�2���|E� ћ�u�y������	�1��F��wgU���U�ޙt���G9�Q{�zb�oý'�̾@�JS]B5Mw��f*PnV.���6�Wrw�.ћϵ���h���`v8M}o{�������;�9����>mq����sF3�wFm����b�~��χ�L1�i诒cĐo֣����Ȣv6PLT����c.i'ί4s�IȞ�M%���@ȋs|���ju�A/Fk�ϴoo}~���R\8�>�R۽����^��r��g7�WY�3]Uk>��[����������PI��\�S�N��O�;i�8��{s���ז7�ӑ:�%�M�+�&W��*���A��d�y����T��{y�&����L����z���\d�I����ht(�n���q�uՏG˳�+C�4y������y��P��)���%R��Յw�+x��G3F��X�*B��e����@t'j)���ێ�Zr��e'��{|�����>5�+,GTK��T���D@T+++"q��~�)e��I9V�Ԁ�Q�|w;/i[�&!���p�(�-���gQ]��;�3�>˖2��Z���d�;����߱Ү����t�'�:K����c���<����J�!��c5����,
��ZW&�6���t�1���H�i=X`�i�D5����t8L���t2ўʝ!p�]Qك2)��xe�v���T�1���Ŕ}n#*��Ɠ5�n[&��%%;���	uj^�R�������r��mM;J���R�x �z�~��T�<	�L*S<V�ҝ��!��8���䳣���r�}�;�^�n6l�exH��&߲&���b#�*\)@z�&�6__�oB��wK4V��D]]b���x�tW�\�1���u���&J��^���{yK�D��ٶ=G"7�*��]p��Y���%��f������N?#1�G��YU
D�r��z:�1\Vǡ�wY�7x���0�ɍ�)R����=ǰ��/��uAt��'��X=���ɹ�ī�f����ԯ/���6r@�#�d��x9T��`PBŉטx�e���,ɷ���$�h]�ق� �&A�sc���t�XN��fV1G��՞5cs��"�Ӕ��+{�8Z�mX���t!��_.�]+a�yB���^i�8�Qr{nǞU�5�^	��[�u�����>�ޱ����ݕ�9�s��x�u���i�*y�D^n��e��ah�c���+,�R�1�E��$˯GOB����� :�]�^&n�Ǣ�F ��9B&����=	<w�oP�s/��8{�P�i���Wp
k�g"z�K�Z�ˎۭ�=^;�+�U��<�n��%r��mm��b{���|l�;Q">��q!����b���=��X�Ɯ�=�+�f-�̝j�����g��νV��GV͐Vm=<�,I(^|3�N����S��ޜ���8��@T�3����N���*VQ�Zg^�j�����]N�R���yLz�YF�H������T���'2�O\G|�# KQ��r�xS��r�Q��J��Z��r����i�F$3<$O�#�J���t��É�ʡ���)ꑛ��S�����Ȟ���D���T�;17�}�>��Pq�A�y�R2ˉ�C�n��G�����7�nߺrorW�\�r�vO4�ڡ�*��g#k��e䮳 ��&Ў�>�Nr͂��"%�u�X==���pp�E�gs[�eE�������:��s�S���W�y���Ga�%������kg���왵R��$2��
]��w�|�/���i�ՓH�Eg����a�n*;��#k��R�v~H�I���dd���M�f;}3W��k:)TX\�9 �}��7<���G�w����+Ű��w��@{tJ��U��k�� ���\�@�*{ y)�/�y(�o�tczϦf����lz��ѹ�z�G��c�B���+ն��zro�{���'�ۓ��v0�]z�^ˌ�+քz��Mp��;�}�(�w���=E୉�Zz�,[@��OF[o��Ǫv�7æL��#��蚴�z�fBF�ek�=/�i�C�֋�|/W2M��w&,t{5V��8_UF�ݗ�,�f7��}��9m]���h����53�l�$�JғQ��5�j�-3^]�١���>��ݕ�0�C�r40�g�aԦH>�jf�{q�^���D_M �\�J��x=��y{H&s��Ȭ�����>Ę���}�@��FOMM���H���1�TB�}�wyq�a���B�1��պ�κ��i�q�����c[S溶?O�ϳP��y�k�����:,��K�YB�z������2(��^<e��j����8׮�BRm�`tn�q�r���K����l�Q��Y}��p���3n�!6�N�Ѩc�
��H���o3�G:��f���]F^�!k7�S2��GľK�k�H: �wm�mE�@:e�ӽ���|,���ue`�*��}��:����5����{\fboz�b���o;2���D_G��3��M�Еt1�ʮ��xfD'���r���P���QAzW�K
G��u|���T���c��)�iݡwS�.��g=�m��4f�W��K�S^e��EY��w����=}��/U�����'������7�[`��y�UL�t�C�D�o����tŸyy�{ݜ���*��65)Y�:���|��3*T`�-i�鼎�&�z�聽/^���
�=�%��*˼S3/;ɠAʡ��g�M�.0l�Wj�C3�t^�A���MKD���B�>�ً��)*~F��^��N�=�'>ιu��K;�S�̟<��]]�#����+�ݻhݪV���雧8|�65a��T��5٤z�Ψ��zV��P�N��Vu�'��sa��S�7�c�+�\�^��w�;3�_>T��~��iKXd��LD''���P��@���s:OZ�$�=�-���[�]ݖy�>~�H.�p��JT����WX�BuO���2|t��1�K�\Cr��QX������O�*Iy��mF�d���Q�
.������뉛����ׯ�P��+�D��;�B]x,������������c���ӂ���4At ��hnM�%����l�"�0���v<��&��Rj����.>'6b�+�')�_�i�A+�:�Z&IX����uЉ�
x�<����\��������czr�շ-�ǽ][��7>��a.���7z/�?r��nO��Ϊ+;�������M��^)wQ @I�k�y����7	휆װ-ҡ9�>�t���qfÉ;����O���_�w�����+�}��]�X��#�=7������>!�Ǟ����޲��W�v�s�f�3�\̜�]~��X������U���}R]%�*�k���:����?�=�~}�˵���ޛ%{��":�ZZ��}�#6_9w��L�melf��=��.�i<��$I�ӌã�\��5����q�%5��\���t<�gݐd����\��2�m�jPݵI'�sZsVr��V?=��=�=�����k-�:��􉖬��{���rPG;�A}彽�x9��5ѱ��_��:�b��epUt��T�n������J{��K	+���w�k`[�D<�C:�vfE�~V׷:g��f�����Q.��EF��Ύ��|��#=9y�j��]��̄ͨ��Mapn]�6n<z��K�;b�{s��	�9�j�bG�tP��6^�^�x(���׳6Nĕ몑�U<���J�<��N��]m�"�����T8���dV?k���#��ran��i�L�1^4�>X�
!��̒2˜�������6e�f����r\�+���w�EY5b�3]����:���kۛ�zT�ϨQ���M�V.h}�͔�ڝ����"��+�k�(h�E��me�eڙ��������~Шe�<]VO�m�y����˨�RX��d�>�>;)�F*='l�U�Jm�p���,)�\�^�U	�@W*gG� ��>���|��rL�W�7Zs ?wឦ=8��[�j�P��_7��R̹Y���8���1#_�f�iJ!���F�&�垘�!'�N��4檡ֵ2�ޒ�v��5kC����:ȍ=�7�_m� 6��]+���.� ��Mi۠_w�J��Z<�3��
ٵ��X|�����ʴ��E��]V�;�#1%a�9�&z�t�!��I���UN�nr��H�\�UԷ{�5/^�z]~ieD��[�&���9����ڧH�s1�gfk��|�i����꾗[���v�zfW�����9{�<�Aŷ��(��d"�����꙼�vC�ƙ+�p��N����L>��>/*/x^mMҍ�����*�J�RИܪ�ؿ@����.\�2�m���ed��~��S�D*��Շ����΄\t/S����]a�n:�"ĭ��+��}�L^��Y�o�]�,�����K����lf������\�K��e�;ݧ��*m�}���Ȧ4r��$��e�>U5vwI�X*o\)7�×\z��&�e枥��	Y���r�c{m����)f@ ����mK���j;��G�c0<˫
ʥ]�"�j6B�w�HM|�-���-S���b�GCs~����r��+0?TGx�{b�Gzʓ��:��Wq�{��տ<���IW�e�[sT$���1B7�fE%OI�OUz����X<�c�ՏԼ��;V�V߄��;�5?c&��[�l�����/չ�%`��`ָ����ڑO~�I������Z�9\�L��R,n8���m�w�4�4ˊ8^�����U����'ҩ!�ܾ��s��F�f�eGw�׹N����i�I�F1�����ץ���3���?��V*>�7�t,��=f��9G����U)��qE<�#�˺c�쌈Z﹪7�};r=�Z#�>??�.���b�ucFV��<Zyj�zQ=	Bb�#Ua���c{�q3&����\ϢN��ͯ~��e���M�a��\��AK{�H>w��Wk�|��hD��g�ᱜ�>�/(�z^�t�	g$�.��1�Rٛq��@RsxU��w�U94�c��y�VQ�g��\��%=�{C�r����ْ.G ��[��v�O�::בӅ�a�� ��\!v���W�1I������uIp^<^�|}�w�v���īe[�@9Օ���v�R�%��;�t0�M�{H�*z(���*L�X����6������K�`�w	.l�[�W�gw.��vQR�WNa����F�f�ǯt-�����Ӷ�<��&�I���2_Vqw;��	d�8"������4f�疇R���"`{5�۷3b��U��D|���'\"�G7v���:r���:Lv)�ټ����ּ������抟b�c��a���Xà:o-�bº����Q�Pz]振U�<Ďf��/f^�[�i��\ٛ,_�UG97�F5��M]�������;e)���InZ��E����A�.]w_��5ʭE	�P�.(K']�k��/�o��G�&��_a�Ꞿ=�f�;�����Y�ׇ�"��	w���E��l���U�����)CK#a���}�I��t�{,MY�����\���j�0�eݸ�3��S��eَ{��"=G�rϦ�V���E�/3S��&=��K���X(�QqˬF�NW�=�R��vc?�L��&&v��.��p�tl�$����>���کa�8a}﯇].z������>��/e���|�'j1�^�|�s͇�4�/D,����hmT��q7���5��<����ܿX�S�u+VD���'农ս�Ձfp��s^��㴽�1v$g�b�X��_���J+BZb2��>B�)Oan�k��z�{|���:�I6�4lps�歘���Oo<z0�*������%�'���Z���&^�����4R)��X�(�,�J�T�c�ڳz�A/9왘H_�۠:o$l�W%��Q��Ѕ��qK� Of�.��ʷV�y6n��7Ezxl=�R=j���\��>>�Q�fr��Ja/��cqɵ�; ��ta�Z�F�vŉۜZ�tLޗZ�9=�
�.G�K�N=��2��2�)r�쭄�<��B��|��q�8۩�+�U��y�:��S7A��q7`s�D�3�+����i�F]=᏾j��{���q�ъ��(��Cx���<�nEG�gQ�����	�ޑ�I؆�^-�<or=ּ�vҴvrjK��b��YG/ۖ���x��{������W�:���f���e|��������{��X��r'��XxM��s+�����b��&���<
��V�����Y]
��SǳL��6+C����	A<r3+�I/B�\[�w�ϕ�D�SEB�����ɨ�3M�c+f�i,YX}��w.��U�j}`s~G��l�@맡t&2@��x�d�u���j`�zLg��A��k�N�7�>i2w�w�l����lTS�V!!�v=��]neo*�?�D'�~ wԥK���+z�Cu5L{�hQO9�P#w�=|��s�۰^���u��}�t'�����H4��S�B;�6�H�{���8�u��{�Gr�r8��7W_%�2��v�.e>��w#Tww���b�WQ�
ìR�nk��N�j:E�B�<g�͚嗸lt�g��m7VkG����iz
��y��𱻹uDŀH�*����P�le���[�}Nƶ�A��m�P9�j"��yr�s����ތ��7�lh�KA��	{��5;hldAm:�W ��7���HW����i���5�����N����Sw�
G7��D��ʙ;q�b�c�2��D>� a':ޢ{��sQ�D��蚲�]��|�=:��Z�Lk��7�6󀔖>o����������w�t�6�%lQn�Àl���uuA����[��0��PMdLR����v+�O6�v�.ΜB5����e��ޢph�wN榑�W+Y)�i�ýrA*�zŜ��Mv]���[L]�����N�e�ɖu���Bk ��+]w4��t_N�r��A��C��2��:�]j[]G��ъtAk�#F��W6�"ŗR��ebX4��n��R�&!�3n���찪��M&����Q9�.D��`�`�j�u&��1A��9+����eH�D��:s:]���˥]v7��q�����ʣ�j9gsh͝[!B=�v��*k��� �,Y��c�Y8M6���*�Ÿ������=��vKmK뎲`�dg;h�X��0HQ����een�oa �Ф�Z�����D����;w�|R�f�@p��ۙ�S�2�V)NQ|�c�³q��/8ؒ	@��3�����B���V�Q�����GZb�k�Ng?6vpPCs`�S9��:����3����{MF�Rwc��m��z��ͬ��K�U
�/;���R��o�ۧ��-�U�:��P┝ϫ�v��۸�oZ����:u������W�8����6T΍bU��c�Tt%y�c��\R\^Q�	w����9�s��cΡ�y���m����Sh�qɒ���7Sx4��|���Uk-=��:b�gi��o8R��nnL �Ǜ��)�W�����"�w8XO��(�f�擛-�뷍+g��eɥ1j�1zOs��٭�v:�ܣ,t;,r�{�kw�2�=i^wR���p�_���L�@#R�G�j�b�cvx�YC2^�V7r>��K�\��@�XR�\&���&��i����̛5]n��VW(�Y�
��Lar�1!Y>�!(���7uء5��"�����sJ\6Ѳ����Q��%n%m5�!�����8$Qt3��z���[�y���g��s���%H�-�|�KZ	������w.�9�U�f��滀�1��v���/��f��v��N��fn��/2��n{��g.�`�db%8B-Nz�r��Ǜ�3:����;E�%�H&�8���5�;�1��Ǒ�&UNc��+��������=�����o0�h7߯v[���k�:��u}Åv7i�W����(���8Ю: ����U1�O�ʵ��L%��Q��ve=�^��B�Hg�ݶ<���($x����fZ߬��"u��[�im>������Cc/�}ɻ�? <���;�Twޣ�R=&�)��rc+asx}�͝�'ٻEP�R�A���%�\奙bb��F0���?c|jn�{�/�rW��	���O��UN��_%�"��X){m�~��YȏZ�=º�t�0!�72t٬\w�w5(3~�g�w9p����2;�1�Ĩ.��ن�����݉���~��~u��ɇ|xW3�	Ն]'jq��7A�05��=�e��/�]��/����y�R�i���̽��y��Mm����(�kݭY��=���ܗ�cT"Ȏ=���
����91 8o���"cs2u{�NC[�1�O+�Y�[�{�q ���O�~���;���.36�	�3�:j�:YE��^��R3�'����ܮ��姂[�I�4�4Y'��7��/���?qv�4?-��g���a��*�Z��S^��o�f&��r�kV>|)�lGp��T���[wn�/�67|�+�����r'�4d��$��GZ��Q����hLwZ�����.�.���
IK�#�Ja�9"6s]�"���z�)M���n����f���뽬���X��9���Sydq
���2��f;)�5#U�-�]>Yv�g��͖��Ǣ�������,�-8{<cف��s.��VoH+J�;���lJ=��S>bqOmMz5�G�s9ޑ8����spa�G�@UE�+:zS0��n�/=�u݇]]0��k�|�p��;�aeG�˒+k�0�z[���;�t��E��3�vp�s��Ƶ�Wd#��P�3#��o�lW
���ȁMy2��ϵ�}��������\����KѺr�Ft���TCe��3�\D�5�Ѿ�{Pp��[�N���$u�U^���#�5tc������O�H헬��������4(}����n������M#������G�Kpp��k,�*�fgؒj ��,�s-��G�0�����d�L�2ﶄ���O�*��)�ஸ������Ν�u���Jg�Vj{�4�W~q��(�k^xi�����\Y���Fi�4��t1R��ЫS��^��({�Tb��]c�^+������Ex '�.Wwǳ|�=	��Ҵgl��p�6LjO�'a�Mט���~ҕ�7F���7]n."D�i�yJq���,{.�$Ff�ޭ �=�<Oe�',�u�M^��޺[э�������Uv�0�]J�k�ۑ��FӦ�tc�ټ�AD������s��ڿ�uY�RƔ�w��%�E w���1|�-��t-���{)��KS횈~�x�zu=y+�>�V���U��<���K�?C�k<�VA�}=Y�m�,��zGD���S����j�
a5(P|q��+�3�|b�%�kJ�����^^޾�qpNO�k��W�F�e,3
�mu�{�9Gx�z�]��C��^>J��.�|N�}R�z=[Mұ~��j�Z����w��n�����I��[ݟ�o*���4w8h���R˾W�tq�\W�p���DD�EP	ު0U���u��f]���_m;�< 9�&Nv��װ*p^G�B>�^b�b��x���Of��P�yL��A�[�{����g�|�x�]�>0�u�Y�}2c߬.:O1�ڲ�ɭ���/v-���*|����(�1�tn��|�TЈ>x������k�~2b���Tl�}]Bs2�iM.�Dϕ����b'Y�v�@p"���xwr��L���g��wQ]޻]�	��6�EFZ��SC����z��zp��Ƿ��3��w�~�Ƙ����S�wYJo���O���א�+�����o�mI����!�n�;ɴ=�������;�)[d�.�
�cӝmi��Gn�5�b.�}��3}�*��m�6�{����Ħ�Ø�孺
�ㄲn���Z��O4mpzxj1�p��Z4�)F�;�I�٪��}Y�d���*
��r�o�kY��a<��LΣr�8&�Q����{Us2��s{�Kُ1P�^�(y�
��o����㻕���<Qz��H��"||�f,��ጠ�sj��I�gt��*�EL���P��\or��&�7+�Į�z'����X'�!�h>Qtmk����ѳ�UU�h�#�� ui.��gX:���<���{
�
p�r��ΜE@
����H輝u��*��+�K����E��jf�s��%x���ȱ"�{�U!oњuq;��ot�׎�����_��;��ߪ�=ޏ�p��Q�C��/C~^>��cs��y`z�G
�+���=�o��js��rt]�dXw3��i�M��	ޮ���l��P��l�㒠U1}�%�m���6���~�C���R)҂Ӭ�"��\���uC�E�
��砺o��әw&��8&�P��R�ׯ����ˎ��qI���Z[3贸��u�.�#֤� q�Q^��|�ݞݗY�;�;9X|U���b�s1&!W-U�I��ǳ�V�BQʄ���z �wd�(��M�Y�6"k��S��0���<ǭ��'v�磴�Ic��Ec���hW�ffl6տ�e�ٳ4�P8gJ����W�����ϰa�M�`bN"�P�d$��fV�&�N$Or��~)	�����f��<
�-r����M	c�us�AS�w=[���m��B��wP��x�A�d���j�l��r�� �4v��E�s��x�CM#1!Л�ɘ��L���#=�~�N�t�eγ;׼u�d=��s���U��ٌy}UDb^t�v����B���!�#يO�m��|g���;
��f����t�1v(��s�c�6����ہ����j®�>�l�lիEJ=4�z�Y5��V��wVR�y�m^tG�ȋ~��z:_@f.e��>���s�}��k��#A�b��l@�o�ː������3鄹�Aq�.	D9�THS7)�EJ��"V轱A��~��uѺ�5�܁���g������2���u6�X��E0�q����}?E���W�]M����}�������4;�L3+��7;f����8&��7ۂ�!�W���^��i�Wu�Te�/a�C�U\���bP��3l�4�b��ň��e�W�F�x'�u�+�1_�Ĥ��DU��כ��<CTi����1�e{�;��QN�g�˼��Ы���6��y�w�(M��AQ��"��;��W���LM�j��u��"�%pN��U}[t�컕����=���^2X@2o�=Y����ފ�UA�kΚ/w�\�@]em!����
N4�X��*T�+F]pJ������_t=/M��E�%d�E0��k,�gbvm�(y�r�Z&RW)Ҥ��ڨf�Na�E��I��#nnf޷��NEb%����f��gT��1�c�����zL��t8��5,��.}�v�yU���o[�7��Uy������QJ����|�� j&|p�l��t�]������=NN��.9�}��|=�t݋�^���6�Ó�WNE�ٙ�!κ�
�ׯ���<q�;v����w�D��������|\R8�f��Q7i��q�17���ܛ*Ň7�g�_n ~���[����q�}ǫ���r]��'(��N"����[��7R�k)���s�������_
���!7.��K�p�8J��N��n:�<%2�z�ҧރ5c{)�h9 ��Rz~�\^�W�4�	�a����po�H׭q�pU���N^�u��=sx�_ʗw^���Y��b]�>(tO�Dv^xf��#�_D���^�bt�b}Mq.H�lN_��}E�y{�QyVT��.����l�U_^/����F��!�2��]W�-�sG�:C�򸯑�����_?��Y{~����:�Q��BAc�7ZN����V�eUE�OCޜ���*���,E�/@lD�E#ƨf�߭{�Bqt{}�AX��C�{���Z2�u�T��YYhVg<ۙ�$L/��+��t�>�r'�����bU�n��r��N��M�������p�K�ht�.l�єq�وm�.is��3�ʸ�t%i���_Z���.ٙY��%�-.؂��d���ZK��_Vc�v���*Y�hy��jjT�F�]��8��q��j�̋=��:�7��x�s����q�S�������v�R͠�-��c+��*���|&��k�4�4~Ma�{��yS}��s��ި{]�ա	��D,
E���)�x�uøc�����r�2�µZ��^�l��F��)]8�^����j1ȗnfGR(?1WB���Ƣ�®�҅>� �|���n/��E�л|o�W��y�N{$� J�R�_4-�y?�+�Q�W7�����_�Q�vGS�0gYُ��(���bܚs�Zp��'�%@�N��>6��}��^���dzYW4�7',魨^�/%>Մ�6��Q{9zhpys����)Z"'�'���|~,��Z�;�	���{Ϲ_�Jf�p�������C��:���S���D�M�R��"'f"yz?AJ��W,o�q����~n8�UFU��$����u�{�����2����+�-1�׬�&��(�ܲ�_�*����GdB��������r�g�g��wx�y�����*�qL�P���ߪ��腆!���Bew�O��"���U���&b���Pá����HAT�ঢ়�ɮ�H9^�D�܋�Iyuh]��)a�П>��8B}�����V�Z�/+J�#��H�4��*:�t�q�ʖ�g�O¢�[�}�tS��^�駹��T�K��x��'r�<��V�Wse�{����֩i����.�F�O(����ۃ�dd� ���?m�h;�o������b��&b�G�����;�Fa�=�d��X��:�Ftm}���7&��j���J�����_�|7�����+�G��^�]'���I�~뎘�Qಕ#;��#�j��;~�1�����B��׹���eٻyb^ս�e	BTĺ<���W�15��&�s��J*���H��j1u�2%E(���ms���K����z2srd�1�닖D)���c����oK���2e�~�OL�
���L9��|*�jb��L�H<�e��V����MW�F�m�?R	�Ƽ�*E�d�*�&�LЫ�-����0�1�/έ�ڼ+ܹ֭�T"����=+7�e7e�d�v���T۱P��.#�&�jH�x"��#K��zj��Dz�ϩ�a�z��w�w)�������b.���n�PDc�P�J���g����t������C���#�0����+��߻�S�ǣ��'�������X����{���z*"3'�YDCΰ�:��=i��I����u��$�/���%bUr��k+�SwR�Ӱ�3Un�Ffϱ�u+��$���u�k_|ޘ�p
t�C���]ꮜ :��^8����{�M�����0h�O_wC��.�w)�|Z�[�]pDd<�P賗�ݑ��u�a �;�<!�����*9��w6�Hy
�'==T�s�<����_��MM�͎�;)�V�;p:U�U�.3�RB��F�Z�(�c{�~Z�ϭz�ٖF��9^6��h�̅�Oa-�� ^��
}�(�s�f�>XMm܄�����(]N'�~"Gvc?���S���A�^Οi��=m�5�:��5G�@��S[��̧'2.��]��i��G��׹S�w^#��3�o��;oD
uc��؝|w%�b��
��@�빶�]�<��VY�l��O���
���8_��ܰk��y�aЇU�Fp'�*�PeA�>�ѣ����z�[�菌}9MM��TӾ��r��e����T"�'�k��Ӭo�#+�c�8��2����B�T��Z���uѽ�uzb�P� U��?ua�0�U���m:P�C;�t�/�b��U�{�+�6��{��ܟ�_r+Xm���9�q%�Q��P��0��a�w&��s��8�*={^�5ܣg�������t��>�����/�T]ot�|�]a&g��!������&*�}bpF+|�:&�/'ڷ��:E�&����U�o�O�Y��5�˭i!F��"�f[)Tnl����WJ�T]f�.�M����ӫ'���L��{���$:^�M��|��U��
W��tl��� uzf�(G�{��٫)��஋[ߖA�gu���Q�ʸ����|�ۂ�E�y`�\������^3���yb�\>�X�D��q��V8z�c���8��tc۸�M��5YOjd-�Mɢn+<���2BSU����!�،���e2�PˏU˷�z`Ľo�#)^�ٹ�ٷ�)�~^��*��Ά�i�>��K�Qi#��Ї������Ѡ����zsșx��`���q�ʻ�λ~��^mֱ��([7�	݌U�9�1��ƞߗ=���w������JT�g��z^��<�\8���������`������S���hF��{���mK��-l��R��"���9X�]j�߳���U^���Q�v�(����N���3UPaު�?w+���}=��,[?��h�]�!.��غu7�v.��Gba_����[S-�ʈ�ԝG��9�Mzd�pӏ��ƨ��k��������ۛ]*�>���ٟR1�����T���St3�r�C��^�v%��T����|c�H7:7l��99�{#���uz2G ��7o}�tW*���٧���jϢ�X�_�y�#e{�|���`�|�v:]+z�{��ڗ�6t�t\��M��K�;���DZ��lY�cH��q�!���G�V��͒W^#�����r�����n��nmD�,9�QɈ��&�څk*4Ջ�Xl�<L.�G���������Y�6���n�0�+���s��RZ5�n�q��r�EC��+����|d)��̲̕�{�!]f�gm���⸡y�K���R���a�o��$���S��n<�gug&��|2�����n%���h�vQ���3�����y�X���Z{%�uv��AX!R��xkNd9J�=$��U�9��6v�X�M�J����S�a��r��3U�]�����t����l�Jj����	����F���p��|�*;�w�:���|j�N}y��08��=�X��.෰�="���mc�0�Қ�����N�nL��殽�hf���đL��\����CK�ڥ�1'��.��廷�QI�A��+��٧�PVNN���_���ևA��1�����Bw-v��o�V�]�r:56�kYx�(̬.':KӶ��0r�flm�zЩ�KVI]��B�e��*'��i���Ѧ��ƯȵŒ�eӵo���fsa'cy
�\�
l+���h�rȾ�`�0�it��B�f�`VWR��z�>Dc�:��Ց[c�봥���gb��[y��K�ŧ:���4�YW������D�S��kn�:Ws��
2��+k1�������_-��f�ӣ��]c\�J�fcw�W:�x54D�S,^I���8�<̉n^��I9"zwHa�m�m\���+�eq����N�]��d�;\2�l��#Qn؂��n�]t�R�(еzK����[!��jWhZ��n�z��NQY��"a��gj�Q>��1��Y�ҔQJ�ɰ}R�)�]]3\����s���ݖP��@a���͆u*��.D���lQ�\�:X����e�E�o���NB��5�̾�k�4��0*�"�m�F��ݱ��1�����^*ƫ�9�5������PM|�#�ޱ��{#\ ��«��H�hMcUm�J�t#�Vچ�<���^�;b3Yn�j�]�n����M���u)�������N���'�bO�$q�\�$�aᲝ:z��c*�Yr�xa���AZ�Y{rgd}ht�2�1��z�5�5��ǓP'CW
b�:�[��/�r�c�����p���h�w97�wO!���Pu:�t���q�:��=YD7�EyY9��rb`�T�+D5Y�ݧM����!�/�������_����mJ@5t�>m
<%I���R�d�j%hލ�g���Uh�öU���)R�_oE�BiA+�NEԮ��/��O������!;��f�����*�G�Y�+�t�
^�SRo�fĨxj�� wkW3m2��P���~���_$8QɆ0����ҍ=��K��N�g��9P��5�{%I�\k�-�
�/��ü�k3��t�@k-ŷ�u�2C}[�>�&�(m�w&�0]���N�e"K�5�;��;\�T�`�	oeG]���no%�����w���]l>(#���=����Ӓ.��O�+a+�2=���Zg�ez�=���-Ȫ�u�󻮾�?z�EC9-G/Hi��\U�9���d��Gq Q�,;�9,��	�e����u�]Ԫ�V<7}�`4�p^?H7n8�j�q^ٻ���f�| }�u�Y��ݓ��ǜ��޿Y&gۙ�V�R��Aj:���T\�t��p�h3�Bc���>	d�Ԛ���C{zR�]�r�>~8���s�Os����+���]���!	�u���Q�;Z�U���97�_c�7�n[������LC�uQ*���W���{7ק��yf�o�{TP����~U:��l��uN�C��]	�m���DӚ�vZ�u4a�}a_ �2�Ξ�=�z��U�n�Z��~�D���M7��΀�,�ג�gD�����Ĵ��5M�|���v��Ec�.2���mǗ��{����}�I;�nlM`������r�M�z ](l�~Ep&�{�#��{�U|��L؏]�<�@��L�W�K~ݽ�p�X�l#~��%��0����hp���Mǣ<��p"9+!�~aw���o�@yTDD+>Ow�L6�-��t��1e����C���e&�[����؊Թ�\���<pjZ8_q�WWas/��q�8b��Z��Ҷ.|^�u�E
×[	W�k&_&�ϑ�7�[�}9�X��O���P�j�ǎ>�em%:��r �VɊ�fp )�}_�T�N���O�i-�:Uv⊿1�f��{3���a'���w�4��_�cN��V�.<O��X��w�p翿+>k�ݪ������(ku��:gzj'��XU���5�\����W=�2Aq��w^Oz z�ܫUc�
���ݨ���t�5Ϛ�0S�D��闆�tϣBd�s�f"�h�ʮ�s�L��n�&_-�ee!:{׵����-���T�]�P����:�f�n��vj�c�t¼��=��-���}Y��.�&)	�(J:�X��	�Z��B���ᱴ��xZ�ǅ�� �?`k���]��9�ڱ��cJg�s���XG��-�V����͂��~� S�vN)}Q/����zj��Slg���ɡ�7t񈙒���V��w�c!��ڪ�����W�H����g���� Կ�����d�ϗW(p�pz�U�	�1	�H�Vל]>Rw��z'4ok��؎���\-#����f^6�%^�n"���?4��B=S~��MT{\����qXU:�RW�V�@�|2B�z��v����� ��ׯ\���UWSԦ$scf��)N8��FQU�Oj����ޞ�t���R���ؚ����#R�V
�ةCćǍi=x�7�4���MFP��7�T��v\��;�Ҁˌ�;+�B���p��;i�q$�[.��.|��M��+:y�)A3qJ�#6�w�4����#/�Gx5�߰��¨��������9٣ow�'G{�:�6&��K�ںC��Өغ`)v�3;�^0��x�أ`�gnX+��g��H�#��w�o���:)�Giݸ���`2r6�}b�W�� *ٚ}��J%�q�D����xz����.ƕ�3����ߐ!G�,,�g�W�+3�X���h�f*#tB�Q07�X�c���`h�<�jy;�	Hm�{�ۣ<��7��<�Xo��2\u p���x�]�[������E^�;>Q��>���;��a�*�0R�d�Y�g('�8�P	�2;���jG7���Nv�+4%�n�/���2���^�5��U�ͺ��;K���������2�|�K ��ٛų�f{O.$��w��#�>�bE��#��rt��1s���~�9[���$�� �ǣ��|��?�bE�=\⟞��o}W�wWY�uR
R�Y��g>׵[2�|�U^���W��^7o�6}�*/�5n��[Z-��ы�Ø�'���\M�$�JR;��)��n��sT��;��P$���RUC�ݼ�)98�j��]�ÍߘWL]�&!�ڤ1���33�\WG����8�����C�%�8p�9J��9����Fg5n�}��r�uu#�{B��l�uz�3L����X'1jdɵ�w<��*�íB�:�:3'�0aX3ծ�<��-Zݕg*$D#�S���^^��N��# �W6���y��8R��#`��Y؇,�V*q�14z��Οq{PY�I�G}�ٽJ��NF��lڼ� x�f�'���UoU����t�70d��Y�q��R��Փc(�^��h����V�:.{��������|�||<��}k��|��EAT�eg<w�Y��$�&'�z�q�"�"^��*��7S�fJw�B� l2�)�x�}T��������Hລ5r)�%Hx�O"���*/:6��2 ��T&f]�2b��%�4�؎	��b$ױ���Ut�-Bk�����ꛅ�N`���Us������ϖ��sQ��n���w���݉��7��Sz%׭�ٞʂ�s["����I`�����B�~��6�jِ�����>��Q���n"����e(�wz樍�+��o�����jPl5s�{�pm���@�7�g�����w����:��X���_]�K��S��5�!��T7[/�fU$���v�s��n|#�!P;\<�/;�o���7@��Ɏ��X!���i{1�U�U�1z�o�d>�n���C�7Å�
�Зw�����}��f
��R��=�S���ܻ�b'�}�|���S��NFq���{QQR*���~�/@w��ۈ�V��x����Fɨ˗nm"�D�n���8ʱh��2Z�kU>�]x�A�]s��,�٭�6N@	%o�;ќ�v����̷�p�Z�ď�N�:o0�.-�0���f�I9r'�B��V}��Ɨx�2nH��E���x������w��>����t�.�����,��
q��\x:��ϲ\p�T���<�u����D�Hn+u��9��9��\lE��'��,�&�C��k���5�SJR�}xFwr��/-ߐ�_�\���W�Y"�ڪ�RUl��gɵ�*C�e���h�]��_���x�E(k�ߕ�/q���y�&��n��:�7)ך�YqU��r�=��÷�%vz��Q����m����雅�8]T��΅���G	����N.K��H����	68�����}�19��U��:V����oO�}�;&}U�n�ľE푕��B�v�Q�菊��c0��z�P�f�w�K�ds�O1pۘ����z~xN�O6�{%X�j^�N�-�q�[�dsGMژ���WF<��|e��(k�u�h���o3�ٌ޺Rf���>�i��w��]��y���5@�|]���.Mvu8Wޘ3*�{���W�/ K�N�yVT)�S�ö���@\8�|����O�}�65:����/7�ՙ�z�����P�=����k��ߕM_:��N��L��j��o���=�[����Su�}��e�;���Z��^Z���L�{$�y]���c�F�.l�I����X9�;@�ꎳ/q������sr=�z�7QYMwwF�9���K��
��U`���hV'�����tek��p�9s�(����>�˯;�)w4��6��h��gI�I���9�8"-T��e?m!,�g�������ql��w�킣H��b�a���}0��W��s���Wf���{�'-��/�c�0�fv�Ak�d?d�M3���}vv�5;T���O<��v��HU�6�z:�{x��zqʒ{4����Mlx?T�r�::�d��ј�����ʤ@��V�$��'{�4�E�u��V�-�e�gpt�`?/B�R��)�ļ�<C�%��a�4���;?5�I����w�z��]�U�<�C�uj���^���т�xD�K�%�<������̿�ӧ��¼(fW���Y��'��P��s��.�)�3��������u��/,�S�HT~��Lh j.�����º
��DV,��^�q���1�7�n�eo�'f*i볂b���t�X�+�oI@Wr��v��=K�}�J���,o�`��;��k�}X��&|��ѷ����}9d�;��¾T�.�5lY�6Ͱ�5���7������{:ޭ�^#�v�E^\��uc��B{�����/J�*|*&_v��{���#w�n��J�D/\�-~ǉ%ϧ	������'^�Axf�������]p���q����^VI��d��u/�����(�+�o��Wf�=��"U���)�k�U6�!ze۔��ZH��Y'fS�A-�oP�!
�S��'4�՗L�	�����d��H��$Xz,�r�&�-����IV)�`�T%���j��#�s1.1�:W �w.��+v8h�;w�Nwt{��\=ޢ�mÜp+��7�|g�m��Fɖ��.��+��!�@���gk�����]���d۳bc�R��VPs�37|����yM�ú]sÕ<�Fp�}/�ƺ��Z>)�a��w7aM��k�DOA��$�s�L]/LM�鯦y��W�u�k0�9�y/��#^oz��^����������VXu����}s���+B�]S50w/j��j�c-��K�y�>C�c����	�;k9������u���f�[�����?������;Nߒt����E�r�2Z���^D�=��#e��k$��xE���׸kg�����wY����y�7�)�(��k�(��ޚ]뜤Fw�"Y��^�~9��%�eĿvPm3�#d�{�ۏ���l(�s���@��	�i|��+{����uw��Ӿ��]��y�p�<U�x�Y���f�{������D��gͿ�/��p^y� WkC �Ǜ���c"=Ǎ��S�<��w���u�t���W����ϗ�����^��~�y;������a��'d� \�t�hlNc��p�j����ٱ����W������4�y��uџ4 ��E��X����/!ՉR`0Ġ����K<����M�h��+��(;k[�����bM˖m��񼲨gEϚ�ӷ�dW��q.�C����o59�d_>3+�ؤ��C�
b�Y�E'����%`�Ej�����4�{M[^�W�]'�+F��U�}�9��˵9�m�ZS�Ϩ�X�^�s�
�f������~��}������z;�w�h���lPj��u-\O0I�՞N_��=�M��쯽_lNz��~��%>SI]���ݩ�µ�MЌS��>�3%҈���ȕ6�'m������f9�@�k�i����i�@D*<���o�Ls�޻6�Vx��t& �hM��eґ^�{�1j��ϯP�&�/�927�T�_s�o�Q�Iİ�k֏�#)��E�l�s�7
�`��6={>uj��U��u��̌���6�e!="�93��3cF�pv|	e�
�=kcEF.�<D{�x����r�R�ko��.r�"C����*�3<��g��֯���_e�"��k��8��!N����D3���[ˢ��bv�̕�2���b���b	�}�>�I�q_���^?.�=3v����������}�S��[�U����5�u��n]J��
����Y����=t�F��e�%��#�J�Q�|�Bk��9�>Sj��S�џV#�+6ߚ!�!���K�Yg4�r�;�ub���lۀ�
���CD!�'�/V�s-rs��9wr�tz[W��H'�U�k#�/X�����jNݍe�݂�ač9IN׼V�)S�/r�嘤�&,�jIs�㈻�׶�nm81,,�츯J����yԓ�J�rөݚ�����#�k��C2~�=��B�"��>��OAnF��=;l�w�jb��W;�%W}=/)�F���q��e��ͷPs M��#���b��5�虭![}��ՙ97a��H˒�c��5v����}i�^T��"0Xh��D@�b�{GUh��m�ʊϔyI���i����<�̫�C-��퓝�OK�ڬ���}|:Q����4
���#N�EͲRs�gc�g.�j�S�_1�ɪ��
9���i��n���C�}=f����ўҎG{@S��s�3q�s�;�4:��V�_�
��<~��}�����o��S^{��=�#��!�J:fTKka�N,��dء���l�a�����l^��ܥ��f}�Ӓ�9A����_,U|��#���~Y"��ZwUs(��vH�{���"o�*�VB��95�}���=ġ�G�ҽf�~r�7��1�w�����|���y2`{���;<W�eG[��w��y��-	pԠ�Nת=���z7ߘ?�E�&`w�����We�qN���Z�F�q�o��f��}Q))�
�O�1�
UZ,e����>W��I��[�	����<�W�k�vA�W�;�n� �t@�T��fF_�fZ^��w�I�5�M��`��t�X�v�Op
b~��`Q���)����zK�-��*e�+Hw�{�jgw�cu��-ʊ`*��[I�%���{�D�>���;�M�Z��+�Z�vm&�G�417NンU˶�Gvpض��[Z_2�ح�^s��q󃷻^m����-ն�����>s�cGu��e���݈���/�g���.n}�v����R�cx(�6g1��w��us�-Ƕ:��Qm+�E�B�5-9�K8kق�{P�f�������3T�<�����?�nuԫ�����u�y�+�rc�r��^�wv�u�&`<E���Y��v��7"v��v�V��ìg��
�(��<�ߥ����,��%h^��ʱ)dCy�i&k-�B��J��c��.�.����G���p#�7>������L����}R9>y�Qa��5霶z=6���3_8rl9���έr� �	b����s�5�d�wL�����q�N|�@�}���MF�>��&��5Q7ީ�ne,�pC�n)V�&��}�u����^��n��Y����&�K��uw��j��֊�κ�=���^z��Z��S�/��-��|=I^=BߐS�[�Ͻ︀k)dѰg�2��f���;WB�ث��K��%��@��8vW�7~�Z���ʍ�hd�*⺶���tb�d��@{���mq�r��p�/��4�|��p���V� 7�hIw�,Q��1�̻���>E��B궅����{.33TH�9�r�����qUI�Op����������U:ū}%4��;I�+Uo<=�a̫�X��r��_<��*��s�ֲNw���i1��6�z�a��$��!�;
���7+72tړ�������bȨ��rW3;YR���,�죆;��
,���\���̽�vo�U�MK��4�o�w{�7^��Ѯm3ϭ��2vݠ�Iz�����CD�C��R��6epp�E��_�f�h��X2�dgi����pt��''��`��Nb��m(2�E/��꜇Q�W����
���9ӕ�uq��I�)3�9(8��N�p1�q�Ǫ�i=|��9]b@�E�Ҵ ��.;�[�V7����c�y��<����V�@�,��� *ǀ�8�!���ғ�JVI�z�E���P�c%�Q�'U9[e�mS�*
�Y�^�`��6���������gYre��Y�q��JM]e4��,$U�a�p}�\��	�oy������.��\�0Wsskk���̨���ou��9�6�_Z��a$�<��}rA�߱�B���7I��k�E���˙����\��]W�At�LѶ���R�z�N��{�������Ku��p{C���S9y��M�o(���,�ff�uZpi@Vt�9����,���b���� R;���y%ӷ���\�x��9g-�{u�ܘ��e+3C�`vb�(��Z���Ep�\���!E��?�W6�6�Kʺd��)׵b�_*��w��n4xi q�n<n霫Am�څ�G;���p4È�/�(:uc�;s�X��y�{�}1Y7�J}�[���1"Osf��I�8v���e[9�q �^��4c�K dҍZ�Y��Ę�����@L��8V�ZQ��.�2�Yo�p]����F.����_^Ih�_Y[�V����8�$��<����SB�ޠSnc7iJۤ���Z�՛��* ��]�gs��cw���(R��]����S݇�$��PHkxQ�5m�X�	���K�o����L�q�wu��ܭp�Sϯ�xj�(�D>'Բb���,�����k�j�V�.����5�{��ih,�cO�@>��ld2����b���+}u��*{Ċӽ�c�#X�<�+��xŉa�P��tc�i�ꝫ�����@M�
�R[�gb��+�6w&l�U�U��m#+�6�����rbe�bȀx;2�-�xJ�p*2�}=[�*�[�7]�"���\y������VݴV.�Ƹ��{Br�so/�P)<��y�)�{��W���,΢�5���r���@:a㼶\�a����} X�et�k�<�A�u�+Q5��Xa64N-�R�O*�}�|2����.����e���u�ḽD2��F�v^�sCE˼�[�N��M��m�7H{�a�Y������Vs{�r����[P��.��%Z̹b��y�u��o��9�x���k�����X%e���Kݾ��L��y�	����e�1�Y<yR����o�,�Jsm�_��Z�|2�ܤGZ�pSy�\�.�<*�u"'_QK ��oo#(;gl*]��B��o
�#-He���Zźk�JoN/�m���Iuj �������9���ɒ��V��7�˘Ժ�������Nׯ����������G<6<��u$��q7Q���vX]8��� u�������)2~���y���F��篷,o>O��&c&Б�WI����]B�e��� !I�����ٔ{�-�ɴ���C?F�/+���T��(�t7���9B�ǩ��\�1Q���;�y�x�t@��.��B������c���fpڤ�![`eZ3�+:񞌚��)�e���緶�Y��U�8�O�}�1UՁ�\�����k��C)z�������	�cj����H�1��Yz��R�F�$ס�(>���>�=�sG������ݰGFM!!��Xv��U�L��榇�U��<�F_7ր�ɮ�Y�Y�ӷ�Ɏ�����K��g�����	�\��9��^'�Z�U�,� �ɿ+$�c\߳0��x�eSc*�+|g��Ay��eۨ���9����f��÷��b�E��G��SQ.�=�*ԏ�c=i��'�.%���=}����̎�7K�D�����1�<-�C�����p��u$��v��0 ~�q=0��{� �7tdf��^8�n[є���ƲO�yФ�jYR3o�6�g��p6�z�GnK!�L��;&�F9�9��քb�����ظC��}Wz��:���������%N��ܨ`ᕓs�{��2Y�tjr!ݙ�֩kba����w\kB��+/��ZKRD��ͣ���S�������]�Y��&��g}�[��l�X�Tf�C.�ku��S�����M3���~�3iadu�U,��ܤ��D�t�ES�Oj瞌ާ�1"��^��x��� M�/x�jB-k���2>ع�LǸB�L*�Pǣ��y�}y��#w�c��\��Eg���Kܮ���i��v�N֤�+�;U̊L���T<T(B�h���!�3���sݢgk�r5x,�>�J��c͓ەe��e�=�)��Bd)NhW�S���a��sP׹2*rʌ�wqK�m��,��[Hh/|���tc�?g&G��Th�)�Vb�B�w�;��J�ߥ��ͫ�hi�����@���.�u-o�,�� �С��cq�wd�."�u��*�>_zn�8��ɣ�}/{��`�2�����q�wO�iIZ2�l��oɯl��L�zg�Q��205|����y{BuE��z�z�J;4�a���3}:aI��S�9�iK�4�JciYk��=r��z"Ϲ)R�*"��z�c�N��H�w�;�^3Ҫ��n�'�}FT{dh嘷�܉��)���6u�Pu�{�����Xg���vkL�OD��P��u�v
 ��4�-=U\M�b��uےs��u}Wy�1�u�3�j�{�F�m5��]F���F�<S�����n�`]��*r�J/l�:����=7�v ��wZ���:��9�0�|t�&w���ɫ.����ݮ��W�_o��$Wcj�`h̨�,\���v���d�*ٍ��F�s�Y�e��޳������]��ٶ�UF�r=<|�]��,�r8�LH����5ɯ|��߯Z���]���v��U��ر#���wyNy
k�X�n���_�e���ۢ�O��x|򧬾�d�(�!�����s�ٺD8T��]��hJ�&<y�[�6T�n���9Y��v���:	L��fpH�s�|ƿ��q���s+����R� �I4��ہwp����"+�v'/_���BWE��[ޮ{J+x��6��9�m�����F�l�|��z����G�8���b��Y��j=��in�ʩ��׮�3�����Z�Ơn��WWy�S. "���|S�#jkg���ř|��g�Q㒶U"���9��M{&ի�7�&������;����"��5�7g-J�K�J'�����r受=|��-��
x�َ|ܡ��N���QNa6�O��#������/�+���u*~9+����A������O��������{��t�|�fV���é�*_�j�k�Y!9!��,gJnn����闺��b��*<h���l�z�q�Ua�n����|�-c^wD�M^��{�Jg���4��ŧ�6�T�tt�s5�ݺ����V��T.L��!�oe-;@J`[7���Pt��Y]�����V�nna�p��� �MM�i��z�X��B�N�qC���$����c6z�e���g'��D�6Jٷ���iX7�s��d﷍0}�X�ڴ��7�f�{x��c�?v���1�+���Q�MJ.o2 T�"L]���fG��y�8�^�~5�=qw~�����n��q�t�4 �L���)��3�R(o�Y����>�<j��C6��Dbrd��6��i�oK^s�f�;�:>�w���G���%G�Iݙ߿R�~՚�v��=�1[�X�WÙ������k4:�~��=��+�m�z�y�'2&nk�.�}u�%��ӽٜ��8�s�[��jz*���n�jB2;6�c�b�'f*�Y������ �����d�޼پ�/[n��z#޴b:}����:�����'��(��.��z�yO�/{��9��P�W�O�ݯ;2f�=�(����d�BQ�CJ*9�d�����ے�]�^=�"t�b�0k�Y{l��]X|��.�U�}Rz�Sӣ=��CWL���x2��U�t��5V�Z�aѝ�AI��%��(��IB�fo�p8;tOs�Q���}<��;5dw���S�����/�NN-�R� יCޫ)�/=���������,6�)c������u��������6�s��a��B��G����S2t6rj���R�P�|q�֤j��yf�%���k�h.�����_n.�����+)��d��s�!�!S]La�}���o���Q����5�Ҝ��VN�lY�m�j��U��ړ�����u�����Y�*S{R��}��;n���4��v��/�3�^ZZ
���=������lk������Z3:�������@�g�|i�"��g���S�io��,}������~�$��;�v3ҹ��j��w��+
<*|�����1�v����d�ո?_�4�f�Їg���B��ٝ��=� }��n�t+�6~b3��Fo�ETm$�g�~�]�L�2ݵ川*�aі:��[%/ث�N�/dNW&��`t�5��dm�7�㗋�[�k�dA�~�����)N�*��l��w�W�,���ը_����.N���U���T��%�]G��Z-�[���"�Xi�a}xf�uU cc�'�ه�L�ȣK(oa��F�w;�@T��7]��}F��5*��o��Z�b��&z1k�ΈJ��}=;��l�+�1�l;ǵ�gg�[��$y=/G.�%T��sq/�����I`��YW:��V̫u�^>���e�����щS��h����p��)�z�Z	UM���1{&ɇP�	{[�#tn��'{����+�� L&�+��l�y�@���Ι].Z"� 立��(���
���~y��?v0}��v|�nv�S���*�[-�L�sRF��uV���"ϸ�.D��E��CO&�̰�9��}5k��d_���fk%��[��V胠=s��\\�F�dE����R���{E�HU�uڍBM\�{��9�#n� g3��:e]^�2�v�4��N���¯�B�y�3�\�+�e�1��Ԫ�_lH���V���\�R�y}E��^�jw���l�nrxx�t� �z�i߱�!<#=�%<���r�&�2�}��Q�XĖ��T�v��<��SPEa1�J���_����:�dg_��#���&פ����*����j�U�N.�=�5�����B��oNh�k�SǱ�+÷���Rks��@�,4��~������:�陮����`	�kj�����f7�8Lƴ&S���S`�{��N�go��zY����]ۓ��; ���I����{�.�����8o�:s���s�*�(aUt�ǟ�У��[���w�,��}�,v]���!?7��<�������� ��ş`w�[C��F�xeZ�'�zC+$��p�
�?�z�����}�Z������ ��q���<}���ї����zEJY�3m�g|�A�޻�Ѳ�<߳"�ѵM�^�j���ʧ"��N�;����M�١k��T?z���fB�&V�3�V}�[H�B�|��.kὖtW�kЈ͸G���@���U>�ϳ�����rUc���:��j߭M��SMM��#7�5]��t]v'�4��F��9�T������E]V��2���
�"��e�������_@��[�/"?/KK!��Vu߫h)�FE���uZ����L��ڴ�����U�����u�IR�9g�f:;j���A}wwu��������j�AS��u��ǥK�n^���QXVHo��V�y�`�҃�]=������m�mw
�Y\�sЭ���L%v�O�5��-��^N�G�$�����,���<Gpu{���h�>�wv�w�
��o��}�V�g�}�#���W
?�v	����v�C�J���@��Y[�O=}^a�V���>�De۝������"f-�d����@��܋?Y���qs����H�׾۪���>m޸�R��>�꾮����������H?W��h��<A_OV��ۛ??�t����uT���v�϶s�'wؿ=����Ps���K����t�3O ;w#��HR���b+Z���������k�~�<��w��x��ҿ�_;P�����;�W�H�W|���wsE�o��bݯ�E��y��A[sp���s�R�O�jX��0��s�p�M��~���K~�L,C:����Fc��+|2��u؁��vg.w7uK�c	��)�6Fh�����_Pxr�}κ�bf�7��_?}���Q3(ws�1n�����츻ɬЎ�_ׂ} �ۥz^�Wz�'�瓯�v����o����@�=^
��%�n��ּ>�=yzZ�E�,u"�]���̞޻v u����Ꜽ�"��ʞ��~BL�N(��e��b����^aκ}M�������ױs�F�c�����NL�c���0�����; �=t��S��zo�[�b�4:�d^梩��wC��*^V�W��h���,���d�T�ܱ#k{��.�uчn�0�h�M79RV�9f^��b�&�>�JnXM^��ɿ��:�b�b��j7,��t���f�.�{���Õ����s�ZľC����-��Ѡ�z�r���S����Oߥ��~O�AjM|v�W����ѣ�Z�T�ǜ�9�_���a�<���ˢ��D^k���mF��u^�1����ĩ}mUϽ! Ǚk���ܴ���r�|v�������E�ݬS����s���{/wH�l��Ǽ]�#������q���06���fM���@�b`������C�ήS�},Շ}�d��F]�q�-�����g#Ez�q�f�m�g�!A~~d�hnkBTc���TD:�/]�B�U�{���e�V�Ň�g
�r��6��Ի�g�G7��V�y^|�6����y��z�ɐL뇿X�����oa��=Ob��5"��}��s��闞��NE��ȶKaG��fE1B~[ݕ��7#�{��V�b�#���6�x,�ڽ�k��o��N{(Ӊ�����=7����tۦ��vv�l���pʟ_�3]�$1D�����������R�J:���~r!)p�^z�-�쪞�Uq��9�����:鐫����}٬�����Q���=�xP��Uզ�?����
s�~-¿������%Ĵu�ZXhb�����c��O_�od�촒�M����?��f9��©�y�}�%���ܿ��V}y��D6��g �9��kzi�w͝���g{�}��F=����{lu|����R��"�y�-Tφ�����8o��h��F��b�ę�Eԉ����7���S�m(�etC���e��b��k���)�aCM����J���Ѓ�z�?�����JXj��3��Kz�vX�뜎��ۣ�E>���E�H�,���:^�2T���sv�P��L��
W�	�<ݺ�g�׸57s�� y�������j�	�fe�ڮ8!��(P��7nf���Y+�q���e�2�\�vD�����r�Ԁ�,�[�ϡ�\�qWX*�}Z��c�ɮ���t�.��z�l�Yݪ�x��],�@���{=e��_���ϭ�g�O*���|]g�û�����@����d�ow������uW��O�q%yzokە�;�S�˙;}S֣oky����N�h�����CT�?Vg����xWRwՕu��k*|��0=�k��2��_�g�27OЖrJ>�DO/��fP��t}IN�{��ßn����~]���4!��ӸWĿ���,�O5e�^�^tΟecڼ���]�����|N�����>��k�K�����o���Z��gO��z�R�9>���{�'qN*�y1O��I/�<��rN����x�������b͹�8�Mh�����M��%�p��u�u_�#�R�y���S��o&Z�Jm�}}0�� 	�@�L�T��W��)z���>K�GA��:^��}����>�^��κ�{hd4Q��5Uv1E��� \�(�Sڤ���̀����e3̵�^�AjOׂ���U�y]N�O*���W[��9yʍ�������3�сdP�hκ�<ӡ{J�8����ԁKD��,~�G��Ժ(��Io����o[�����Щxwu�pJ�I۩['_t�֣I�]�Ν+H]{`|s��\��:���ַ���,Q��X �;X��]o��߯g�<ŝ�g�eeD��0C��+g>�����ο����4����1��CD��;�n}��<G��(«
/�GA��s�VSq�*��	ѭh�En�ḭf�dŝ���� ������Sq�@�k%�ܭ���=�,߯'���N��1�1��'��	����+!�=tzv�}���i����<+�#goٯw+,��[��� ԭ�?+�3�2ԉ�jXs�:~���ٟuy�6z�P�şW\D���cƴ���1�Ηf��r��i���)�uRɛ���v��	��T���y�\0ߓװ]�a�b�zz���sq�S��l+�v��A���_b�~��К�m��_3�31K��nrC�Wyp.�k�>�k�����)�G�3��͘��K�C��f�#�J�����ƍےiL��z��DIa��	4�cS�
=Dze��܈˺�ױ���]��ܙڈ��9�]};��+�.{�o<�\����PD{�X�����ш�A2$ὐ�p<`�~��L��?+�[c�~���}�ǭ�j�@�������|���gm{�X�>F�t��@�Ԁ��}f�����sa��:�uO��eJ�_����ɺ�=�꾳>7>w�y�M��������;2}�edN��� T޻��K�_��[�o�7��7�gKV�;��J�w87�m�A4	gi�F�6y"���5R������x����߽?��V�l-��H(ʙ�� ����w0�u,�t��e헜��R�5@�4��㖺��X�@��nr%n���N��+1��:�k�R��Zy��j̾�*�ϱ��U�k�sVaDb���a���\�Wq����:����;�b�tݗiN��Y��c���Wr���QsJ�J8��\�Iu�#����;��2愜NqPhԬ�/�<���{�.l)��c��u�傦�V M��^���L��;l��T�u�)���d�[�T��{Z�]�HZ���O�sh۸��9�ban	���Ge�.�([le�1�=@e.��+-Ŕ�#����1+�̥���nn-Y5��:�뺦u�N����lsE�wL����ֱ�n�N७��h99���Xe;�7 �Ӊ�T��6+��wJ���E�['XU{��V���biJ�X.Jz���I��{{��� ����vNҗLi�`Uyo��Q�f�D��@=�N��M��4. ��
OC%9���݊G�5�m�3&:y�z^?�f��3�W�xEq]�p[���qm�����{�Ԓ]��v�B�+��Ԯ���k��^m��K�z�wP�k�X��ڋA)f|�WQ��t��{'t[+[n�:F�R|�����Yk5�dN��d���*�U�����R�T����]�J��%s��e����݋c.ü�ս.GZ�9f���K��ힻ����%v��+��d�7��N��NwI|'Lw���z��,�C�1<��CVli���t���F�W����Χ&��ou!4u�R73�����ռ�D͢5��6��˳����),b���6�<s��].���,u@�%1fС�6Sk*�M *�f�[�ӡ>_�:����hd��]Ik�/A�!+��.g
����S-��*՗����=�y�5A��ĳ%=2Q�{�	Js��2��dCrޕ	�n>0�7ýY���>�A�8d�f���'Q�Р��"U3�{b�9��W%s�c�d<2�t�h��Y𥋧N�sP�[M��rރ.�8�"^�|'&�Rb�p�5U�U�ۮ�LJr�m�xYV�c|:�W��Q�J�L��=Fέ�W:����^
�q�:��%'!�s�]�~g�ڥ�S�%Ź������E�uZ�)���^Nc2��NF�K����l��)�ݕ0_+䷲-��Î����X$��[3M��Ǚ�Ft�%-�Ǫ��#r>��wX�ar�Z��'���8�@�B�r�c/QIf�\�첫Ln.�Wx
��v	=@n�Dx����-*ߊ޹�!3�纐�q�q�05�Ny��ws6���ӫ�υH��\@�VӖ�[��*��3�v=�񝤝��*'��uڌ��q�aU��2�冂�4�5�O́&��r9FfmU��!�+h�u�ۥ��z�Ű��i۴��憴�+��λ3��D1��(a�Gi5v��9:P���s����,7���nS�6��1ӣ��J�T*�O�	8{q��Mq��1?���߳w����y�=���u,�<�;B|��{��s2^�����7s���9��7��ч<�e���g%�Ө��\�`@󯃃u���C�>�v�G���3��ho_{&�z$�R!�T�y��5	��{��<��ۼr�9١�&���`x�d��S��eT�ȷw�y�N+�6jp�cٙ�lSΧ��ީ�m+�������w�t��|n�ؙ���8W3=쒉����6\�1�c.���>#���7�X-k�s�_G��w�鷑�tU�����<d�?6�n�ؙ y�M+�T�疪�2$����s�ߪ߲棩��~�ޅ�bcK�黰�%K:A�L���� ӷ|k�=Ogs��E�9~�5ww�B�h�_ �>���ӱ1w�ςή�Y��9Pc�W�t����=��#����(g�\����R�G��w�^�ɬc�4`Ҍ�î;��pW��K_Gܷ=9@�'�t��.�E�+u=W�**�#R���j5M�}�1����r.}�с��	�|��>8}9y����G�_��ê%���'���30��n�nTR��&ɬ��pJ��%_���_Z���kc\M�0�����$���tr�-�����n���6-��*���`p����:��KjE�x�"���ţ0�]�⩲h��D����G��fl�k�7��b��[���/N %��V�oųV��ݳ�[ v��o+S�{[R�onD���{Z�륭p�K)�c5����9}�+�4ɛY�4�ywܮ����W!Ns�:����/H�]��ul��gV��Jo��w��D[�����u���"��O_#L����!
Ԧ{&t>�=���Ǘ1E�j��쎭_|���7����)��`w�����S�vr��߄���8�?4�6��D�Ԡ}��0�7=5<�wz	n�����S��������N���dX����x,Fem8��=韂�Y��^"�W�ydX�R�#����Z3�C1�O�y.SG�홗��rܰO��B�&�DvP��{y"܉�'���5~~ܓ�u+��>>ބ>J��<�of��Zq��d�%�?�g�#Ҥ_�Xp��ݪL�?)؃��})�ſ?Z��WO�ȩz���B�d�p�r��ZLz�-<Dd���G�:�o��>rL������_�'�ocb��ӝ������<a���Ǿ����v��*��9E�9ǁ�9;�C@j)��jo���(��?��D�C��Z�RuL�4b��!��z���t����~أ_�zjc��I���c% Lz�����ɬ�����DJN䗂����ɒ�@�yZ U�%|��*n;�|z�*�3�'_lV%��$x��"�K�s����A��US��T/������W>���"'[�xL}۷c�OG:�uv�:�{�8��zϨ݈fLT�<m} ��װ��U�བྷ����<;=�z$������mN��e0��֟�J��/�u=/+Ty��j���5�0,>��1Vx���ϬO��J�����I���׈M�V&j�n��'��6r�Q�ZqP׼�^���9ox�2���6s�h���;����%�#HrҲ�5wi�q�,�t�z�/��羏y���q�\���^�c��b��^a�1*�yQ{~��3�ݏS�c3��v!��&<}0#�A�������V�1^��c�Qz��>��>�yv�y�x�UפOYZxm���W}]z9<΋�n�� (�
�0u�ݾ���Q�?�sR��+����z�Ոci;�1��!i�QΞ�^�8ƾ˨v���{1���!�rjj�x�/�p�o��O��HZ&#�a$t}�2�q�ˑ��F�5�-{b,۾	��&6�D{�
��9�����G�E�cfb�\�b�mƙ���@��+�^��C�����2������es�G�E�ȡmKY��zF�C���UR�����_h��m�v�8���ǌ���\T�����G�'��Y�uZ���r��Ԑc�u�Kԡ����ˮ�����V��~�~φm>�}��Dr��wΫ{�t��~y�͞��ܬ�'�UG��ٚ{v(3=�2�x��?��M4>)�/�X.�YZ�S�;}����`j��6s�
���^̀3�$'#��YN�J灊�?
-=���)�y�뇺�z�Fk&�Yӯ����oFe��y��1�u�w�{����z�h֦#��=����e�����X��g���ͺ�W�Үv�TO\�nr`@S��=,u�v��x�rN�o���n����B�[������֢�����H��p8z��}m� s� \,Ze��6���ٵ�3���-��%Ϸ��c���v�-.��G(�ص�V����x�W<�P��}��։Pإ�����I��U}uۉ���%	�E�"��5	O���Ғ;5�|��Ǒ;sZ���d�}[�6�q�E��e����,��1rf���qb5�"i�{���L�)痟
��x7���^)s���v!��&˛��{c� Ӟ�Z��>�P�����nN|7"�Լ�8�B�t|*(R2;���I�%:�#�Tj�^���S������7c�/�zW�XǏ�q�[�� W
=Ӫ*�c�,��v���2z7F�g�H�G�#릯ү��lZ����F�f� �&O����{����q�>etfKR��Xf��~�+�J�4��e���׵�߽��݈|H��Ctz������ρQ3$�O6-�=[�Qs
�o�c^W��:�|6�C�W(���W�P����fp#N|��y)!G�T�ѕ�n�6���CW'�7Ztf�j&u��ޥ��S��t�a�W@��n�ˉ}�V�X6�̰ۙ&yg���	��Mc�iU���a�ijr�<|(����	�B�:��m��`D�9K��1Ώ}��םQ�7���)�u
���_Ud��{�e��¦~Vʈ�m����
�������C����ߒn��w�2����E�;g԰�~��� =�d^��3����M����?-��NUխe�=9��Ap���v�H�c܅���r��=�rD8�}�J�ǫș�.�gL�~6�~��:S��=y�U3o�gj{� gَ���bT���q)}1|�1��i���4߽�T���P��%g�[ض�ֲ���fޟ���Vϲ��K���7/��`�ѭ�uY�:�},V���|$��&cYrQPU�����f�T�Q���u*'�	o�$��a+֩P��r��\ڎ�kܹ��ۖݿ��;b<�̑Y�&
�l�C��k���T���ѝTrg�v�U��Tpp͇\�Խ����ن�[R<Eu}*�8^���.�VW�V�Vv�Đ���e��{�3}?|vK�ۺ"����/��d?:cU������D��=\~�>v��R#�⏒��np�U3��vH��d;w���g��Ck�)�L��z�,��p���{o,}/՟f���yH�w�_C�"������f��QӸ!$w��7�Y�����L��L|0�xR��׀�RC�gč�{���~�6�C�R��������N�gҙ4�o�Q�W�bo���U;�C���E8��a}$<�F��*VD}��*\�Φz8ٞ�Y|*���q)�:����:�{�0��z�Զ<~�?J����߇U���J�Ϩ<��j�̕�I��)���n.^٘��̗Tz#f�dj����-��ǆ��.��w��>���|��Ϥ��>���^y,}q.G�b����w��cٜ��#�\�^�Μ��E��ؠ�8�C�/՞Z^�m�4�h1RGɈ������T�z��ݘ�▓t��@���i5a�!{�Z�?>�4���K��
�sG��ɽ��%�K���r�	���dFi�y�G�D���SF�w}��1c�(�����+�z����p�_��ဏ�5���P�������������.�^]=u��êX�%E�_�E+z(�#�۷�h��]}����e�	_�����ǀ~9�� җp�YA��V`Χډ<�Ͻ�X���"����HǕ5��v%�s�Em��֮��V�s]}gS���A_��H�zB�7�o�<��H�+z�Ae��X~����l
.������kYz��W���!o��su��V�}�r{z�O]W�C��	��.,�S�|�U0}܏fG�9��>m[���9���`����t1�~�k�E"��0� ����w{wi���_���.Ǿ꟫NAg��{FI�����3�Tm�Yi+�;<���y_���C�V+�9�eaϜ��c/��s����9C�E��c�o�Z4�Oس2_�� CN۩ƴS��d!Z��.�F��:���
����ӝCd�I����}5ٹ|1��I���Y"�I+��܄u�}�>W_yd�+��ﱏ�~��6F{�hW�l7Y)�.�)>��5�*��q�v��"��n�f;����W���9;~�$�3�ț~q�P�l�_�ù%Ԑ+޳��!��3�/NM��`-��Pt�U~	z~��3}��d��srW:�2ܶ������#�#Ϊ�^('s�_#�X	��HLΪ� ��2"�{��64���a7y�V����Ez:�ۗn'�ݻ�?S
|.ʡ�m��V�f�^���D�!�.�00� �=~4cº<^|I>����2T���W���.����������o�V����P��٨%r�7��^ Y ��;�oZ�89YS�6��H�L�bzX��	�b�&�|Et�}����7`}-�ϖ
Ooec<��ԅCT�f(f����G�ݏm���4z�1�7u���@}�0屎=�����鯊��2���F�� ������\��T����]K�����j����k7��B�MH ���㘻@U�� j1Y�N`��E��_�U�-V	rB8a,�JQ���
�j�Ķ��X��f2�Л?H�b^[��+����cm�K��L[���o��G�n�c��6-dI��;;�Lkp��xn�\`؏ ���0�m��9\bGU�����]��a
w��@^,�w+�!��-����l�)qQ��ݴt��o#S
{��V����
���P�^�+ �M9懶�H?{�<}k4;�|�jG���@�y���6�F>~�Ʒ.����r�o��՜�؛�^�-N���-F�� ���M+�?L�]G��=���vR�����f�� f,s�q�'i����!=3��w��zp�0�=k���|�\�Y-�!qa|��r�D{�ds���7\�{�t|F0^���A���zE��+w돡��Bj��D��p�=
��1��ʰ��h;.��v�V���	7�.�'pQz����ڧ2B=L�~t"��ǝI�"O�k�)o3F�Gʥ��c���/f���c_���y'nN�W%��
�_g{/9���L�(���D1MB8%}�0)!X�|�ˏ|�H`��S���0~V	G�T�2�>����׸\��
.�ގ���s��ߥ�!������"��b�8r�V?������J�"b�ԅ��'����1�ME�X$	D����M@����c��Q���J�o�*`�`E�L���|�Pv��|^s���YAk��z�|Y����ϵ���ğ���m��w ���i:�]Ʊ�j��L@�zY��*8Ǿ}�urk�i��'g3㚐�~T���z���ә�D�,R�/�w<&�*a�w��R��~7�1��}�p1��<iT�!���gOޟ�t]��scۙ�vP�>QEX��{s�|��)wu��6�t� �s$ě;3؃,�?LC���}d�����������,��*�(�R����nz�c�}�J�nl��ޜ0s�0!��<l�/`�� K�/�!g�^ر���l�0��ѡꉏ�D�FY�_*���H
Dm���hgF�Ϥu�}*E�f�r�i�n(:f�;�H�`�!��r��ݽI gtV3����u��� Fn�.��h�,�o��8a�r�Q��x�IY[|{���O���e*U{��<ݧ� �ܤ����)�Ζ���w��Nȫl��n�����g4���"��s;w�ql�|�ar��@_�����:b���NZҪ�d�y��X���BLar;6cOȩ�=3ִ��y]]�˗e!�,k׵���6�ƺ��k}[�q��}shE�?y͑�\��#�~�~\G� (�kf>Y4F%�`�n�YW�$�B39�B*��1��ʛw#O�|�O9���z�Ĕ�?Rj(��r�}HX�B�#,�@���*���C�GTQE� Ue�j*����s xS"_��ݼ4$q���Jy�^cܙ�ÈY��t�0DO� �#��&��yY��ɏxL�8�����r���k�1�[�;D�:�}� G�0"�%�����R�.�b��<��"`<aʇ��3�ܮ-����t�P��^k� ,�`Pg�"G���N�ǹ�t��y\j3��'����_�?V��	��y�<�����g�⎐߄^PE+�����*�����	�ut(���@�'n��!����&�@�������+~��T",�,�w�F
�[��X�9F���K�k*{�cX��^<Y�G�ꏌ��43�<�t2fH�ɳ���PR��FL^v�q$YR@F���ƚF�"0��Ϧ�.c<$g�+��y��n�����&��A�DP�}����s�W����v"b�������ζd���:vd���.�g��Q�i	�����ݽ�}D\��	@�=<��\x��9��z�>�9�����v�##��9�_:h{�2ߔQ�mu� vzm���Wb�����f+g$�0�h���4�2@疩���lީ�A
��V|aǦ>�GԕGݷ��$d�����A��DcH���L48����:�#g��t,�J��^D����U����q��'��T�n,TP�+�m���]��T�u
־�L���U���+���tt��]��������efC�\hVc"�6rk�Ð����Jn�;3��񫶎[=���-]mm�Ӎ�
�*G��Zw�6���=�P�c�+�b��콧��G�KZ�y�F�dMn�Q����.1ց>6"k�؀� �TC*8�%j�M,������F�`�P�!�d��X��eՎV�/$��OU�}��vvu����W�H"�2�ciD����ц&f�Gͱ��,�cJ1�\~7���@��sD2L	���� TG���4�!���?w�􏾖���fm�|>7�:T8LD�����V�Qr�a�G݃d{T>�,�	���I���2$��1����7*���b�;�`��*G��{z#�;&�ݚ�}~�8W�PLm�A��**)R�[�S?0�z��y��v��vо�� 2F�όag�VG��y����� Ջ,�/U��=U���F8�j}����H�-��Wgoh��)�"�G՝c��ƈ+O�Q�F������">,�7\a�_L�C�F!?(��T��k@�w�����ӤǕ8��G F&�)u�^�.�f�>0k��J�r@�P����3��p+\Y |�X�X0�"�q}j�ք�,����z�0=�d��62�<}N�Dw�k��,E�+ta���s�]��v����2-�����P�f�f�@&*D+�X�@�!U��΍��X�P�
aʁ��~��c� �#�V&�bQ$�&}��x�|�=����9\�V�=���J�{f��w�1Dt�$Q�P����aF6�LI����3e'�(����ci tAI �|a�T>ں��� /WTq��N}vE�BmMg�]��M]^����V,f~ݝ�@և��HC�0�M���d@d"/�7��0�;��ޱ$��A,��H���b�!-$���������c�0'Q���Fy�*��E���֤�x������� ��q�C��T$�>A�
>� IG�l��@��� ��j*�O�Pȣ��w BmD_�f/yl�!bz��<Y�0}�D��/	��^���ᵝ�C!�w��f�����e��bW������|m;	,E;�8�7է���{"�tNK/�]�뽖whP
���挾��C!��Avvgs%ŭ9��y3{q����6v�z�vrՋ�4���������֭���>��W��ȼ
p��f��Ԗ�{���[p<G�����V�����P9�g���4�p8z��2<�p�da��W��?}�0>m�l���
a����(�B6P���b�${��C�����%�v�\���>0=��u��j$�uf���(�� ��w��2��iV�@4�*w�����x�1$ W�G�{�ɍ1�C 2�(�Z��MS��ѓ�[�{{-�_\���#����@��.� ��x��Ԋ!���X�^��#HG	�grE|��=(���  4�@#��$� �p���I��/�	0�kTv�(����D���y�*ZG�;5��*~�W:�x�`��;�Fҋ0	�/|��2@����x��f<��](
���T�p�F$�
�Di��ƥ0�m��y�Q�+
�_1c�P����e�����]z��חѽ��>0�
0,�'�؈����`|b�f"�"ԁ�w�E���f~A��DG܀� ��
��DV��Ta�?0=hG�j�'�َHyC.v�	1��Ҁ���;V+��6�ys���}Ӽ;5t��4��FԱF0��#{쩈-2>���q��Hв(���sTV (��S i �@*?T�?(��DN�(�@��n4����@�Z�L��� Yy	:�r�<��g~�ύ
�o`{���E� ������ 0��bUl�/�$@���|D~1��Da��!�8�IƐ4ၩQ� F��H�4� /�@f8�32P������ �b76�)o���:g�����O]n�C�I�#yF��bʏ�D" !HQ I�D|@�c���|�Y���*~���DC"��ؠQ�8�F �Q��0�G�� �0؀��` C�"H@�Ę�"�c��t$���9?/���c�w��(�# ~&(��H"�|@��d��D�!� �b>�N���ڢ��" ���f/�qdDY�D > l� E����>����d�Q�c6�$G��0���>":~ }W����a2}�n�����b>�#Lt�ʀ$��@��I0� d��>T%d
"���	ܙ�4G�"����6��7+o<���"DG�D@�""?�D@�""?�"�� @��D"#��� DD�D"#��� DD�D"#�" @��"��� DDz"�� @�" @�Ȉ"DG�"���� DD@D  D@�  b @��D"#b @��b��L��.O���V� � ���@  nO���F=��J�� : t w�o{v�  M ����
(��ҚP����� �@( �w� : � �<L҂@ 
    
     @ )E�@ �  P � 
   ���(  @�� =��[[��/Jw��=�]m7\��U�4����< q�m���w:�w���l=oҞ�n[�T��-Oo.V�{ޅ쭴����p v�� -����١��^0�:�w�� =_*�Zv�hz<l4(����r�l��{ъ
 �W� p�B���wV��(o;��Ay��h<CB���rTTzy]���  �   �    y�����7�3���yۤ v���z�*�����ё�� ���[j�庄֕W;�W�*vם����w[�-t�1���]��G���h�o8�׭�(( hf��;���绔��we�� ���m�z^w�h�n��h�x�gc�{�ۻ4ᶼGEؠG �E�E=����<�������@�Y�=νtRF  P z�   @  ���Y�^&��wy�tzqtQ�w;��:b:�b�S����=��l��z�E��˔S�����=z������+�[�� ]����m4y�\M-���z @ mow��ڣ�����طo ��y)�oOӢ���s����o]��ǎݳ��w����v��;�;��Ξ�6(���{F����
[!@
 =��   Ҁ@ �KomT��{�u�iwkG�9�:�m�����ON��4� ��m�m;��ks���E�Ǽ�<��g���*�\���k��g^��^{�k� �  ���o=�JW��7�@S���
oy�a��ٶ�k�������{{{L�7E� n��z��y��5��7f��{t����Ӹ��tu�S@@ �x   @   $��{�s��xn����wm!z�<��o[F=6G�m��PWv��x�����+��n���Z�Gy�ݽ.�w�r�z�x�{�m۳�򽷸
  ��Y��ma���={�ҵ wF�r��ha���ް���t�eaӞ�]�v۷W< ={����׶�+�w���wyoCAWL��[o� �?FD�J�   "����I�   &��#"OI��2d���5 JU   � MUA4L ����JF�U   ��w�����ﾑ�~j*�Fp����{6U-�KK�f���:��yP���zP�h���%=
�b�������� �Q�}��>�����L���)�����[r�"���Y���8���gX������|7�j-������0���
��b�)e����u���;��*p&�q	�0����� �'�n��ɴ�L7X] ��g��{�a�L��?	P	�@ ˑ$����y�Uҋ��,�o�э��hQ�Ӑ��2��V:�@��$+X���-��%┸ұ����V��;J�Ȱ_���m��ŝ�+G�����V0�I���p	�"��cENxO�g	�KO��uZ�/���:+FP���@fG�0.�-���(�0�4��S��{��)\���AS5	�Ȭt6j���k4�}ab����%��#µOϩ_C��+��y1�+�@����l�}�ҍ)��A��g~
�c9w=�o�)0��\��/(��la�*�~�rҧSmf��Xyk<�=�uK�+4l�8X��x���z�ݐ�L9����ɮ��s��w�Wi�J��3���;%#u)_��0z�t��ml�SKS�L,�5sYYu���Ȉ�{xBi�)ѤcQwK����Ї0_^G��7��f�Eڻ4�һVJb=�ˆ��p]�"Hu2��7�N��zB�9�Z��K������'��Z/���y.�+ΧE�Ճ�[W�5��gur�L\���+�v�8��W���ـ�I�Y�ٱ�ݵ���.p�}W��Y�3�=9��	A�;U],�N)��w[�u�7wySVO\�)�.����ˋ	޷˝��l]|�����\7o���d�]�)H�	vQ�;�Mk���c6��9��z[T\Vn��V�G�CSP�YHQu�w�W�8%K��mq1��ҹu�m�r���Nņ�h�ܶ���ov��ch�Ë�ؿ`T��]��9T]'\�=l��شp%�-8�:&�ʸ�nRNS�T\4�qn���ܘ{%�rƅӬ��RAA��WWeW�3�������m%Ƒ��-�Ac[��Y/.&n�Q��f�Q&�7{KEf�I�!~9�Z�F�kFՇ�ֶ��]e$]�^���Yɷk&�D��'e��%S�^.���L��̌?2	�|'�x���'Ӿ��Ԕ���$�8'ӿ	�N�O�b~�c�c���~�H���q�~���'xN>=�S����"wÿ@����~��$�;�Q;���N�@��N���u;��؞8:���,����G�O����<���x�r5��cÝ�n�m+���2?b��-�b��0��B�g**b�]���S�:��bR���3w�jf��r�8ܣ�So(�)o:�7m��;ӷ�K�C�9i����piI�0i�4�ދM�*�w�F�kK;�^ڑp�bx�p��)k&�ٮ�r3��6n\'�,�)�����R3B�飫C�S�:�Vܵ]}!�ͦ��9u(�D�ڴJ��ޱǭLο�lD�+���8�/�I͖���*s���y��9-kx�"�*u�����i)�!]l�5z�����	��f� ;5���a\�i$h�7�B&1����{8�;n��]hu�q)��[�[)w:<�''!+�����=�w�����]�f-��s��Rh4]��r-��5[�[�%�>/v��n��Et��ٺ�+z�R�"�D�6�e�̤��U�L���uz�5-��9���Vʚ4�%��
���Že��]���of���L�(X�;�8�{iP)I]��*�Ҁ�6��VL��
�y���k�b��;,���W5���+�kjm�Cg`ذq��pBgf^����&�S�Usnm�y�[b�t ,)F��墎��U�=;�E�OUe��
�T�vԩշ�h�m����T�]���5�:�ˋ4�E��b�h�6��c��Û��x>鯭֫꘡�'tQB�`7E0����Y��C�lљ�����5���U�A���P�/�'�X0r�/�����-I�A��닾��2n���"pu3+�����t7��{	�ń���f�Ic�s{Q���*��$ޞ�w�����;++\8�e��)��q[(bj$���d�6�m̺���)~n�8�U�n�P,+(\�bQn�N���ꄅs�f�Q{E�g���uyHB��Ot��P���pH��]x�}�&��nB�Ά�-]�v��˙~��k)�ʻ*��.����l=��s�S!�̽W�r���.��C�N�#5Ld��T�r
3;�w9����MޞeQu�t�6�<@/��F����㻣�N�Z�f�}cT:�7�YM�	�xE/���"��k���P�B;��j+.�r~XQ��ٻ�������5��bZ�w//#�⻵�EY�DM�Y����C5*V��kuv�n��]9FU��nZ��(���anb:a�bN�q-��L��*bc��4��{�TRn�v���3CTTF�#kk^f}�(�M�2���e5�Z�(,0�ݎ^�y7�u�:���](�u�rJ[�]e4o	���ܷKtK�B�癝�bc���W^vagV��K⬿˷w,vc��*�]�Ε�\'�ຨ����%��F�u?c�#"Ȣ_���&MJ� �q?�P0�\ʘ~W
�PJ���gۊ[�G.[���7N��嶎�6-�+7y��&�&~��ҵ�ĕ|��2�o%�QY8 
LZ �0p:H�r��+�#q+^�h�f�{fo�d�fdʜ�B�@�L�˪�
�2�1<��+m�*ީto�B�f,�Om^�J,��rƫ�H�r�²e4Xt��X��X�w��1�n�
+bh��f�S^Z�A���[#2Ԭ�M���:��WmUn���0��4[4?��c��\k+ �V��V�b/>bL�8�e����ݹ$�Jm�:�fbI/u-�y���^���?~�nժԳ�UӨ�Y�RbZ[�)���K�y`��Ҍ�	��t�"��N�%��'R��׍�[�����`ܺIۃ5��4F���"e���,7oa�)`,*;�0�YH���Y	ۣ��!�t�����zA�u�a�R]����K�;h^l�q2Ma�~��_�Y�n��LЫ72��$X
�l��1tN�Rd�R�
�SP*eȀk�J�LѤ��p�mc�{ł�ٱ��-_¨��Y��*L�51�Œ�f�D�1�
�5���-5�PW�m�Zvɥ����f�y���&���[���
<��P]�m�%�d�7�]�n�n�ܴ�*�h��+.D�M�b��7y�=�)nY�r;X!�ˑ�b�����6�A�B����%�Y����-t�n�!	� aw�yUeڴfh/-Y�I{(����V�g��-��*��݄�2��ƎC����g/C.��e�ǽ�d9�Ȝ��P.�8k8�s��9�^�k>�۰Wb��}��f��jU�Њ�+"A�8Fan��,���Z��)YV>f�$[沜\�M-�"���!��u����,ٶi�`��+6� �e�1P�t�cNk�!���2#�njŬ���'�{H�
B�(���j:��5OIc�5�su3t��fͼ��W��N�ſۨЦ�)2pb�m1�邬n�v��h����C!I7�,�-���-�Ja�y��6�m޹W!y����r��-agf�j4v���;��f]5��ZRT��*d�S-d�ʦ]�Y�D&�J���uM��!�c��v�D�"�)�QI'F�i�:l�Y9p���;�U�W`��Uۛ[ɞ�$_�Vf*J��f��3�6�nJ�1�y�~4b&��@B����)������L���?S떡��tAQ�rfݧ������V{[�����n��Hr<Jِ��A��nKt�G�DF\��Q��)�(/�@������:Uc���t�9�̬���#Y'.�m6$��!xwr�J�r�ե�u��6�Z����&D�fѫ� �6`�ԠY�H��#�W�-8��5��M��6�a���,��!<�4Q/C�r�����7N��j�\�$��d%F(�rE�Ɋ�ba4%���cw�b(��7eT8�D�������D�ZS�oD�5hH*��H�j9�]��s[��8�l\�bg��B&d�X�����	u�0�%E��!KP���,.-�S�5�ɜW�͚��Х�B=���4�a�.ލ���:tf����#,LF�f�©RdY[ �FR��Fʀl��e�,Eê�XR������k�)�lݖk(�ɷ@������o��
�Am���x��nn����l���;a3�+��*TZi`��c��]���K��K�7�(f.�l9v^+���f�m�Ta�#�)C��&��\��(�G��y�����#cX��.���J���Y�v7s�rƊ���7�1���9NU�-�ۼڜ���8$�P����ޕ�u�4��Tͬ�r�b弸,^m��+hq���R�Nf���&�%nS-f8w-�Ũ�,ܫ��J݂�-R�r�r�v��	�$(\6jjxTT&l6+���n��8QQ�SFgp�I.2mL�-��!�E-�ę�~�2��w{��.�=�k�sx�P���R,4yѻ:!˼��췗��(V����x���,�朠�Xp�qn�Cn�b��*��*��?av�+("rҨ� �W�l���Q�׼;��?@0�Xw7[�\,�]��ev꼻;3��23XBц
���*ˋ��#aei��G!,ke-禲�u@�)mc��ևY�X󷭐)rL�Fo��YV�:������<��ugQG��UH�B��+���M5��GZ�l�c�����v%���O0�껬�@ط��"�ϴ���	�Q�� �r�D4 :͹tf��s. �gQ�u��f�f�N�k	���d�/[��%�����I����qR����̳�'�X����ζ���܂,ڵ9����Р�m�u\�8%f��H����\��u]�Wq�Z��{Wb��em,u�X쾢�N=ͮ������U޻*�F�)�yi���O�rQ���1��,� �+��D���t�7n�v�$%�mbĕr����m�'���
v�!��t��o�5C�M>���X��]�]\멾�k�]�����K�a-�����Y�ю����nN;W,��2���tyD�����f%mށ���b����y����ek����RW�#�L�zL'Y�ؘn<ǰ�-�����u�^feiv��_�=W;ol�Hy;\�ٶ���0U�҂V��
ɏD��7zʋ�8���B���s��D��b4P׬��kWY�u@%dU����ҥc��^il������SPT��g>��ijC����-��v�@����e,��$fI�+����7�*\wy�X�����J�f�.2�#i�:��;�#�ٗ�*+���{���3��W'^�4G�Q&Г�ğ�w.�K��,n���I�oun��u�aɄ�-�p�"���hR��+�K4`�N����iީr�x��ӫD�%ې�b5Y��Y])J8��Y�/"h��5���$E5��A�N�jw�l�5~P��y[du.xS/�1�[�_A]��[] Quu- )�v�y&6fRO��W��u+�J�7�i�����쮳DWK)IB-��g����j���V2��]���i�K�:��Y�&��A�K(
0�����Z�~�LS"�췣b��W_�r�۫����p�1�����3��VR��z�}gM��������I<��%}u1�g�}sD8��W�����P?$����u�eR������*PʮoF���ŕ:\g.��w����V�~���K`� �6��y�`ܵ�-*��%�T�FlL]_'��R�x2���cma�ɍֻƟu�eƃ�e`�|���;�3�to���
�v��e:��k	�ީv��T���]��.3gP�V��V�,VG�S<o[���iaoU���P��ܹ�9ݲy��o+7��j�Xd&��%��1�#b42����	�=gT���kf���<@����ۉ�j���u^�pAUx`�QsBr	A�D	��R��w����2�0_��ǔ0��[��H,�c���$#�w!������w7��ꗪ6+���1���B��-<͏:M�\91Ǳ`�9[�{�ΡW[-oW��U�Yg��\��*/a���X9`)C`6��P.����!ڒeD	Qȡ80i��u2 ��)�&�����F�'m^Q��W۷,e�xq�,w8{�`�Z��k�E�QRUт�
��f��wA��L]]'��q�2������]$�!n�{��Zh��)㔄OsU*-�;�[�ˢ��ͫ��w�v� ���&�J���#A��3v�{���b�FnĶi��<�h�у�z����E ��H�[���o��6�ڋ�oUV	�8I8V�f�p�=Fq�����O�mAb��E6�����J]J{6��i�YV'�ؖV͏X-E 	Z`�gٲ�����z+3\�On9�N�#Cv�`R?�e!���l�h�www�t��8�=���?6,�g9��D��ͺ��ȉO�z�?���%*�b��+{���^-��7���VC8{����(���J��l��)e�W�� %ɷ:\�޽� �zv�]�HR��cͽ8(�U�a5
���MiS5���H�2a�t%�Yχ����<$tǹ8��.�[�Q˽�I����5Q�MA&�ZE�ͬ\������*�e�2�Z�ق�<Wx��7R�cL�j'{u4�$9S��Uj��Z_Z�����*�'5~��.6�Hw!!��w^���G�ɷ7�[k/0'La�+S�Su�G6h@
ͣ!��J�f^V��h�[�]�����y_Y�9^jq����o���jV�և�WNx�A;	��I����K�Œ�.2\W
30�n�v
UآY�i^m>[��@��A�e�%^oZ��y�7K?t[�5�	r*w���s4�C���c�r�ɻ�\ڢ	�f���q�YO�x﨤�u��[��t�N���Fp���	��1iP�V�>�|��]5WmB�L�:�.}w�b5iR/�ܙ6�Ζk�������ُFhYXN�LH��P�-]h��qGu�C(��1���,����Ą��d�?��G5+;���6w����P�P�����Z��-��kt��h�-�(:�P�*��rS˭��V���Z� ����\.�khZet���4���m� � B�BI+ (Z ��l��ڀ@@Y!]!0n�n��|�}$�����7�F�II#}$o:H�I�$}$��I�#}$�����7�F�H�I#�$o������7�L�����7�F�H�I#�$o�����$}$�����#}>��II#u&e=X�V7B�l�Ժ��mm]q��B�[�i*�.�VۖZ��۱4e�Yl�
J�p	W�����5`[���iscU/6띭���۱j�m���d-� ,�-c��@ �����qn؊+\�`ڶ
ݕʩ�V�nu4m��7]�K`+n�����e��s�z�m��+m�+Mnn�Ͷݲ�.��5�V�j�6�(;i�V��K#��!@���0h m��fV�ªӖ�VT��%��K���YkF�U-5u���}i)f��#��u�ƅ�f���&���3r�ꢘ�5+q���X�gU����Z�:b���x��m1�]�ɥ��Bm-�b���ۋ��Ih�	���ԛ��(�����Y��CM��ԃ=̾��v��Ld��KWT8�32�ljj�1�Iˊ��Z��(�aqڂ�@Im�O��؛�	�ԅ��v��LƔ��iq\4��m��g��Mc[V/F��=HM_͉�Xz��CRȁC3([�4X�n�XB�t��1֙�j��,�^�)R�+l��]������ᙏ"t��'$��vk�ѳ7R˅V���y�f��ѓ���5���K���=��i�Kx ���5�w����|nB��[y�c~�|���if�<�Ϩݥ4e0�������C2ߒ╮�]\�َC>&�7���KZ6Wbi���`���Ф�Z������I䲲�q'��/�k|������}�f#oieX8O{��	=��-�ͤm��`��>T�B���:���]|��M����ٞ/�2	��S��v�[	JYD+`5vƕ�Y4v���x�����e�viB�*��J2՚k.�Z[/��y���s_����HY�L���f�e-��b9����j��~���g���;�%��\����l�ЅJ��(����&�����F
��[��d��J�E�)f��]��I�#�p��@�Mh;E.��MeX��¼���*ĬYnBV�Yc���6u���Gg�1�m��@����As�G�o�ԕ�>/�zY,o~� ��͵���Ҷ�m�ޮ��@�&���ĬhhV�a1H&��B�@�}�`�!1�#5��}���䑸2����-�#��DGm�Ԋ�in�Ĳ�2�p�]3�q[ĸj��be4���C
-��,
�0�b����Ofi��\����9�dͥڙ���ea�Mc�����.�V����1K[��|�`}�A��c�x��씸�?	j&�Gѷ]��0�P� ���'�� �0����s>g&�lM����n����if�V��nPM4��jb���c�?�R&'�^ԅ�����i��鰛l�4у-qi[�͎�L7f'm�q�9*׮�
��.���g�����m��F4��mDl[�i���hC��4�.�ζ3\�6f�R7;0Md�b9r鄗�5P#�����Q5�G"m��V�	w�����mb:k-R޶��>�׍M+�Ys�1?���/�h9�
ł�����Xm`	�,Bʸ�-�_�鑞1��ث���q5���kgj6X�����Bѭ 14ִ�7a�3Fe��iAHT�307F���J*��=Ͻ-�wf~����|��*���$
Y��[�А�k��l�:\�Y���7��=�X�������x��s,�kl��-��F��5Ы6���w�Lm���&���m��y7�@7f�ri�����,�Z�Z��	��n�Ё�صCu����T�ci�49	�B��Z�AW�[f��q�4������+6��¶kRWa4�L:_.ތh�m�p��S����{����5��}��h�F�K�Z踋���t��	nb�j�����`�˟�)ۼ��ۮ��l��ZMi[T>�P4P=���(ۅ������SJ�f�mP�h3
�\��K-��?KNOu�v�clu����3-�5��W���6k�l���v!`x�-��FlT�;st���m�v%����Eľ�&�eRPt���_��ϖ�˗<>�{1�,7R;GZ�&��:ke�n�S;������a���W:�1eAs6f�;��i�]��1t.����]�0?7{���%D+�#��1���g��z�6�Y-%�u���mfM������ZV�f��S@.R�H��y�ix�w�h���\єV8�$b�|z��|���>`��ۙ�g�jJ9�'�aS7�@IZ���]�m;Z�:Rۭ�@��+�)�%��J�n�����%$��`�6ǿ�}~g'LQ��mB��J����5�؆:&�D�i�������T�_��@h�1])1qn�^�Ņ�F�8=�.���K �!?��v�\�7Kt��<��2X�)%�e����dk�<I����3f�w�/�Ҷ�ݲnщ�[�ձ�Ĭ��z�!�<f�q1�}w��k�֣��GB�Mb`,0�oc��Y���V(��ɑ䧥fK&���Tm����+P��e����6�ke&��9�uV�H���6�{A�a���%�%�ؘ��\�ՙU���ޟ4} ����X?+�e�4�a�`ˊ͝Y��3jM,v���
�t�n���C\�Rl��-�Td}E��:Syc�����ިf>���Eq�ЯB��T�c��R�����D�:�4Զ���޸ü�n�J!I�ZF�1.��}4��չ��ښY�#�d�$��`��m��}5o��p��,�Klmр�.�vt�����&���Su
�%�qn���S�-���CR=��5DMX+Oі�vk=��&�[V�����F�t�vЛ7HFƆm���a�w4����=مv�nAd�B,6f2�t�D�	�oe�X��?w�����^������dk��m��-)4� k{:���	U��B���O�c�Iۍ��y�`N�����Q��d�*���?L�W�fĥ��ĳR��w�����7����x�3�S1�v����3���;�.eݮ�%Op�%�f��ˠ>�,2٥
e�2��� ��j���Z�`1-��)zş�,7MA����7ߚz��/�;ac���ie���4!B|}���:�<�%�:Va�f�kZS���;)����.�7�a��˸�%LfcU;e�Q%M�UA��Y5�"Be6$%Y��KR~6��%�G��[�^�isw��OyѨ���֌�eն�ms�h�R|S'ߛ#3i�j5f7�>�k�z�a�Df�s�[\T4�F[��딎��]=��hln1G�]�i�u]�^��ЋSY6n��Z��Eg��LB�Ã��,�@�l>��̡oaߛ���S�,e0P�ŭ���;�I[��3��vں��j�l9v��7�L�#ƺ���m����%�먡x���e���~��Ȟ]3y���B\��B�F�²�T�ԋ3�ѫy�	����.��g�4=�PU[���.ؖ8̮�\����vJi�2�A���f���h0ml�*_��ٖYo�دWd����3t����oXa$b� ��������͌7F��-�0֛	�If*��/І�}�����'�#�|Y6Ʒ_�z����/�U�6Zf��he�CR�\n�ā�j� �����b��}��6��f��&�7#�W.6R�����5�j�O��h��ŗe����������o�J����ϱ���:���u�Y�>�@N��J��[�w�O���(F�@S����A�_L��Z�6٫�.nA����y�\f)����P��5�#Ulf���޳2���ջY�^��~V�,�/��i���"{�0����5]�ϛ_%}hQJ�v����]�c�뮭m���1��WRz����@����q���*~����Ua��a̯�|&�e�m�~y+�=lK�i�@r�P�B�cD�WRJK&��%&�_���8le��B"8+,6�-�o�,��/�?D�5��[e%\��M�K�l�p�O�e���e�O˾fz�D�����bb�%�(-�h��=L�'�ֺ/���-ڠ�ﻩ�[}��v�i����H��l�`�6����cts�����<��oa�rn�	�աI�j�Mjb����й�͛���ԙՉ.�t�
���,��Ç^6h\4�˶���Յ�}�!�2�hyf[�����hi�����.`�4�!��&	�>�M��:m�h���͉Zز�hK�����ѹ����\3S���o_CY�wM�eu���]�v���j�!��j왌W:n��$����=�L]6�b���Bmq�*m�k���䰛lԫ�����i�5��Lf��5�ƀ!7Ň����x8��hA�ʺ�ڿ�_6k�u�c5ڐ�X�+��l�[�ݾm}(_w����k���~`F�lLu:��o?��;ɔ��NIz�5
KB0-�� E�5͚��4؟6�7�L�V����՞W��3�,sHv����c?��^T��m��P�k�h�cQ�?��0�|�➖�{JL����v�a4ф�UHS.�f�u]e,u��e�ڛ��5�=<��U���g�w�͙��h6e������-�Q����m�r��E�,��m�
w�K��mCc1��am&��B�)�a�X�*�4�DΛ��-l��{6�ZX�*�K�.��94cUҎ���n15�-mv���@�����u���UW.�k�]u�)l�8,՛�eءSZ�1�	m�#c�R��6~�@�_^S���)k
����Ϗ_z4Uº$[6��Ѳ� %����}>@����F��՗EB�R�����d6�K6&4B�a�[���T�|4B���ic(�1Rj���M2v��+��P]����"�)=f��c���Svi)b�t��@�m�1���Z٦I�h�iuְ���
5�0`����`�yg�	�h���`�i�m��W�60Lm��C-���$֓C��#(�u��b�ОJX�fZ�2��˶��
�f&5�s6���ƭ�f\Ѕn�ƎtfͶ���wS����l�JT�m�m��@]n�,3���$f�f�����F�v�]��e��cp$��J�#VV"��� �a"�jЙ��cZBV�=z�e��s�]��4�,5��R��s��GZ���Wk/&5�t��e�����3ZCm�2��C.��7-n���ռ�������V@8qB��ɍ(Yv�D̚`���jWGZ���B�j����I��o(X3]Is#oc�g��6u$�[��)����m�GKl�%�B�.*�͕��#6����j��\HZ
�-�d6����jk�qM��v��J�+f��@i"����±m��Ѵ���x9�g���$=��i.V.�,��f�3����m�L��4��^cK��SB%��d�X8�hY����]c6.J�Zm��uͺ�K�������N����%8ř�T��D��5�h��
�Nlu��skmg;g[gkX��i��-.��[lU]W?��+�_�6����F��j��f^46�v��fcKnrk��$@�l�������$��-F�-�)[��jHn1�O��=@_K(ݗd��f	��.�v���,��ĬƵ�Q��a�b<K]�pl^5se]5(�[XR�p��vԶ�]�Mt։,[���8nҺ��)WS3KZt�=5�W�*��H���.k��:\U��J�l¤%�i�U��-J��Xj�u
9e  ��)TV�ݚBSM�[�.k��R�*�ke1)���l����j�SM��Y,��.&�CF�[���նT~�এ�f�3[����va(ƙ�KP,�Pl[0����lD�1tV?Oc�C�	�n�&1�u�Q�h".(bjb��+4E(@Yp[����n�e)�4��k��$ݷ�t=�u������0k��l�-������7%i�J&���$�W���i�)�4��M���j�������-�-E��6\�U&�[,��`Mo �j�L���?K<y-�pYl��E�󽯊�M��r:ݡP!�tԤf�ѯZ�l�i3+i���yx�,r\��gSE��R�1���7�F�3�?.�䤾��m�0���@�6��etqag�n��j��Kx�Wm����Ev�Ѱc��i��\��[r�)J���5�Y�-�T�ѭ\Ӕ�#��T[��)�n�|z�����l԰��cw �Rv�$��I!�n�K4�]�8�e��M-�0�lty�Lf9���Q63�2}���i����E��(��ۧ�O��HT��Zhk.���z�F�z$��g6�q{�3g]����K�#b�EE�V�Sr������*���,�����A(0����OāZ���f�8��R����J:Q��[5qb���dsXqt�t3�{M'�| �Pq��5��1�Ϟ�����,an6�E�XG:SYJ�r[[>{o���f�K�V�nfkDm�Ի#+A����T�٭٢��c��J7[P%st�-4��9�]r�N��3lMPv��(�Z�[�c��l�B��+����L�J��՗�\mY����P�c1�EV1�:N���:�N���-��֮ѵ��\T.��a��[��l�v��$ �ԡZX�[��&1],F�'L��J� ���,ΥI��@q�i��Z��&�$f�7�]���pwX�te��+I�=C��M��&>��paI�G�m�{Vf\RĹ9d���2�u�f������]���,��ٷˢ���`�
����LGJ�t�V����E�iVB6����RQ,���kx�K�D���@! /��c�����-�H��]�3y��tN�y�w���egAOޗ��Ϟ������_=Z3�eH�bc�g����Z·���H���������A���y���)�#�,�.�ݒ��բ��E��[�J�x��|���!���f������YS6s01j+�d��GPmټJ'����>�2#�5u��k�a\ �{���}�����ե;�s��*���[�V�M�_,�tVYh	:�Ĉ��(n��JEԤ�\���槽�=+j;_�h���b���#�ݩ�*Ccw�i:���N�a���#ў�^�~�y�H�M�=,g����_���~ze�+Q4Z@���+l�q.p��Y�j�/��0���64�Lh��J�Fcm4m �'vlY��~�u��ؽ9�oZ��iU6�3��^U�檳n`^[��|�o��nd��*#M�E��aC|��`'i,%y��Y�Uzm�ki��x)Ɗ8L��<��>��B.�X�Y�>��yVe�{w��8S��Z���&7yh��HT�D̴�5q�����]�����:^��'��WoL�M��y �~�������
���ܞІ���N�������9z��n<���@��x�����y�(��5�4DP���)�`"2a�n-�PZ3B��t��zi�W���~���M>�@�8�mP���f�GΊ�$�ʸ)�KD����J�w(���rܕ=<k������V�G���,�1Iy����R\U�,��B�2�G�^P+H>�]4�@���"m0��*n���7a2�1,�.���B�-�.1��m�� "�Er�7��h��qe�=7�/����Y��P�<��:1n����^+7��s��^�=���u=H�<�u^9#U@��_^Ń�Eﺽ�RCw�86aj�=�V�ٞ���f�f�b��o�����C78��"C+�Q���5��=c��R=��Ķ��$Ǧ�N��"MN�^����L�u���6��3�H矋h��������`��m��3u�m�=u��#V�˩t!ޠg�p}N��:�'|[)�3ee�W�yh[{h3Z��F�j��7ɬ���֪�謒���-��WA�Lɤi���~�z������?CФ&Ĵ$��8P�W�=�s̋���j&���y�%@���L�:�D�D�<s�eߦܹL�^[;<�^��˳<A#�`��#pw��9Nh��U�Ի~���٧�O^��}���=蟳/�Բ�d�i��0^��8� �j�e	XS8�S\�t+
J#��ج���R�nE=��]�k]򟠜�|���g��]�a�" dϾ�Q��sI��L�Ku��\]���������ڏ��t{E�[�6���������Ⱥ�N��m]��:
^�ɰU�p�	��V�X�����{�]:��B�Z@�����"�m�-���\`��ST���R�{shVI~��\����
�{4�q��J���t>Q��d"bpNZ{OG}���wʁ���\����'L���n�E����[�V��d,>�wɓނ���pоh�����y�:l���j�[�'	ۣ��7��"���X*���e�.�x=W"ڏU��8P�l7s����V9K:v�վ�����ze�Y��g{\�
�=�0�QMw�=\{�>ٜ7�ܾg<x��Y��Ů��/�����K���T�J���B0�zh4�u&�[4TЋ��K���-&��b�]H�ڲ�VY�&&�{������eQs���6�&b2�-2��Ш,���*�z5��E��=��ٮ�;}������ᑾ{n�
ԣ3��qd��3
ެ�}>�cb�2��YRln�����W��?yӚ[��[�lpEpU��ɴ�Dխ����#���vȵ9��ֽ�W�I�1p��MT �.�Fl���TBpɮ��H�<���h��ZQc���;�����TE.BO��e�:&�гg��fvow|RA���;�\ףվ�ӻ���g�gv����;��['��L�+�z��&S&0٣	�!�8�������=PԺ�U�c풷v�^���x�
��Y-BBG��6��s�s�,sF��8"Ԭ�uǴK�H+��8Z���w�8��h�ю�l�>��x�=O91��{�}a�:-fe��j���!t�V�g\��Y],�?_{Ş��YhVGV�U(hh�t���7if5���mm��4�!�̈́9��(��WE�l�=c4œX����0u��ةr�C�����6n��u�u��#�m��v8�3��c��ղ��a��hWk�0�mn��sqɄ�����7�暚�*�:QZRiN�r�,8��ۮv��X�q��6�7`íƷ]ոr;������}�ô���u٦�[��
`!H�3�S;?
�2��j{��y��}ݳ{�[�#cu{,N�q[i���:ظp^�{��_%1��E۔gI�3����Q���I�I]����nM���y��^^��V�ޠ=u���6RCW��I좟��z�]�mw���J�<�e�̏Vj�����`��YFh�m��7�����F��.�;��.�p�!��8M�pE|��^)3S�����h�9�����u�bu��(�t�
��'��/�;��m��-G7W�ݾ�*�u�u��imZ��FU�w�72�#vM;�wǘ��N�)dd�ov�=�^��s�������M1�-��R�a����~�$���~��T����]Ed�FfE\��;�N�a�'���Z��ZM֘���.Q�����דk5�78��ˊ̅�0.������Kz�z�<7�/T@�l{qqӤk����_��v	}�,au0����_���߰f�)��%7�B9n������d�&z������{����o�v�r�ȮWi��ͰwY�{Y�.U��z�5;�X�Φ-%�xK�����J�>ѯ7�Eg�H����ݮ��т� K^�R�榎�������Ǎ��H�6�)o/v�۳�ּ����
���m�504�us�6e�b�Tc����k����y�Cd�:$P�N��F��Y`����M;��Ϧ=;DW��~�}���z�wBofcM��kN曩���.W2K?s�z�����Bn���t{l�����l�4�_r�b�L��=���߉�E#�ܽ,���̵��z�;V	�v^T�f1\��W��I?�������f�B����	�͏�����E)낔��@X�ޛ^�k�/9�������`�~�r�� 'y����*ߪ3N�1I��I=���`�V7S��j�r��}S:�_g��\�z{�B�gc���!��ތpZ,�/2[]WY��5OA$my�d�-�%��ױG�%����,�MО礻ܹ�w�j湿F/�@��N���t)X��M�g�h�2�$�n,�<7�s��{q*��݃TQoEһ���\�w�9X|�wVX��DAZ��g{D��liP7�1�u�~xr�U�����x�!�&�B�n��� m�f�c旪'����CW��_
"�ۉ
�c��V�Xk㗚U�I�9S���y��Å�=[�Z͡>�� �[��I�I�є�p�T�@���Y�xnԢ�5}���Y"=�4�4��׵cAݯ�پ'�=�����/gZy�v�-,�t��/[.���ꡥ�d�A�����m��R]\��a����m؞^Y�OP�I���l��n@矖zc�0�6�ǒ��ĺ�]M�Z��w���Wm`������CO=�;�rU,���O��X�ϯԯ~\6�xj����`�H2+�o��KEw�����w��X�I�������Q���딮���R�\�4�����{|o��j�Τ�_�5o���:���3�/zw�nǏ�O�51�H�J.3���&SO3��T����7h���֏\@8J�DIh�W��%�kf���|0 �'���/0� {"T�k�P-��<G�J��-hmvZ�R)���i��yGy�u�bݗ� �ٝ� ]�BSC����N�O	��j����sn����Īu�����(]�{����E]��<F���!���{͞G�z����+�mg7c�a�#����  j��Zk�;7JK���,���a�J4u�k+�ފ]K�@n�ѕY 2�P\"�I�,ۼ��G�~b�fћ{��v����]G�j��2�j/3A�)P	���80K%�A�<:���[x��x�w5;�)��;��xu�4�u�ۿ����y��g}����� -d�מ:\��:�-%v�ܡ�?o��.i�3��+qT]�0ꣂ� ��^o�G�lw~�=�3O��9�N�+��R�Imh�{6��rm��ݾ�n!rBi�fm_��v�-�Dy� ��Pw��w�
���?yC��+��%	^#��\0�*(PY�&�^���s��O/jw.�4���q2�j*qn)���wӵT�V�ݟ��,,�kjgK7G��f�-mdp�|�����N�FL������U��}��Vf>���8�lS�mu���BZ�=�"ov=m�\^[m������Ɏ��y�B���Jie�\�h^�רBcE�l��1�َ�ZG0�kK	u�t4vٵ����a����GH���yFf*5SSkcj�#
�.��&,���E��ؠaG�l6��h!�΅�Z�뒝v#3Vium���O��:�4}�],,e��mwe�Z�v��T����K:˕#6֎����Չk����~�}����B�	���A����5��u"�W��Ԁ�c����T��h5k��J�:��D-�������s��qN�֍��qŴ=�-���E:���v��5�:�3�C�]w�P����/�XѢ�c���=�`��_�WN��,y�JN}L`��ŦŁB��g�?�$H�=���I��z��[;�}���y�v&+'bU5iL=�>s����=�U5����!J�U��w9���e����j��zkdܯ=�Y���&2*^�ߕ�������.���:�~�k��{���!{:W�իųӘ�����Y�������ZC���m����Mj�8��%P��ug�	��B�@#�����.��^��j���xB��. ����V^�N}|��Ւ/^T�K2cź�o�ߖ���Q�=]�[-b,TVa�k
�f6޻kK�5�2͠ۦv�]m�bݣ��Z(��I,��%W��E9%xɞ�:��{�x�8|�����O��b�N,���'b��!*$L�����Q��çt�a0h�����k�=Vv���O�{e$p�9��j�N�x���*����1n\Kd��&�m�IbΚ2��������~���\�ׯ�oޙ�{6~��^b��;fPQ��&�������wP�W��˺Y$�Jʄ�
��&�Z:ߦ˰��w{���ɒ�<�]�YI]I�!��`����}R�mh4nkw5�=,�c��P,��{�W�5��%K�y���&)��	��H��a��p�8�=rܚ���B
�m��0,ʹ��8�}�q��J0p�;���/:E�6j��������{�;ص��0j�g����oYoD�L�[�(�n��ޱ�],�|�h��#�U:Fڮ��ݙ����nJb�l��Y�[�M���^��k�GZԊ�ڊ��!�g���<�3�������)�B�}�cq���T	�k}H���Q�2M��?q�O̮�bl���=&�l ��?X�o=�.�z�q-(Ux��e�� �L��m/_і�Ub�cu����]f jد�� "I�:����b�W��}{ߨ6��].^빓#?D�I���C�y��$G��v9opy�L��r]��36�K6�,�2����DŚw�&ԋ3QmP<ƍa�U;7{v�>��q�p�ue��#y2�u�F?b�a�c��lJ�2�guo�mt�؎����o2�w2�� ���\���q������(v;5�*8��/gk�E�a�����^�|լ��N��V<�N�V��V�>L�z�S�WՑA�#+zLQ�{�RѰ�Au��}�&L|�C0z���p��Whv��o7reg.��:��lf�{�s��Y�:�����3p��n��է��;�����K[7��Ǭ���͑@���Q�4�:��n����d�U�7IȀd]�MYe�jedU�td@*��cs���&J�I=ĵS��ZXwOt�9g��[��5���!ѧ�	���s��;7z��̡Y��%�r�(r�a�0o@�*�H���mW�
K�7�_�Pn�Zײ�&�
��k�o�*+�6"0�����$M��f�en���w;*����oS���@$�4AߺEu4c�ٝ�����oo��ۺx�KZ� +�d�vD���E]3o�V�%u���=�]�:>���oz�FkD��O�.�W}�4�9�3��㛽[�:n����(��%�����v��J��sOp�M�/�^�JL����η�Jӽ1�� /��w�I���&���)�����	{�����&i�0Ky�r)�+��@��wn�����⟛��m���c��4��n�n-u�}��=��ɡ��Z�����_��@��W�У��Q 2���~�4�����ޛG���ٌ`h�o<c��&M��T���D28���#�j��|Lz ɬ�:�_tT���ﰏ6g�N۵��}g����g�5�4~뜶��4G��#�����uK�}Ə=u��<�_D%4}G�bDPB	>0>�G�M[aa��%�9?o��K�%���]}�?p�BQ�	G�F(�!�E��*.H�p/�� {���G��$T���dϼ�~�M~H�dI��B`G��l���:$��q�#����?���)��llƹ��+5\�7lV��u�l:�u�J�F��M1FK����z�����'#�� id]-�?Qڇ5���>��7��#��L������2(�<d�$�r~�����ݏY��H�}��9qq�Jث[�Z�����wh��d�e*Y�i�:2^R`z�<:�}u�D��@��t������4�G�d3��?V\��|�,����Q����"�fפ8��+�#Ƣ>��B�������|8���-����(Q�����{i|�Z�b�BT"C0��~n����'��?��)�wU/�ޏ�(�@c�V�Ox?#�dg@3�w���~���,��i��|��DicC���R�X���"���䣮F���K�?Y�����q�:�ߠ+��?C�l�O�����')�$ꑇ�W6�������X�z��'���Ҥ��`������>��f�^P��׹�E��GM�V�mc�ބ�u�-�?q�����)gfum^�Ǳn��386��E�B�P�i@��rjn��EN��&����� ����DV�JM�D�O䛸#�
�g�j@F�����?��� ��@��|>��q]rz��v�n~�H7u>c���
~_?|(�R���3.���i~����ɡ(F]k��Jz�����MBjf6R�ٻY�A��a`�U�c�}�VԳݡ��)�j��[^m��hc(����>�R���ё5����wi
,��t|$�W
 ]�u�/���P�~˙���M��^R�X��a��	�E�9y���t�F�//��$`2���Ͼ��dE
�[CIy�����6�~���m�j�5�f��t`B��u�� Q ���M�I�G�?Q�f��@����ռ��?"(���}Q��y�to*~�	��rtš-CF}���2E(�6���Q��'.>x~(w�t}����4~��	�ϟ=��8�ǖy|�����fz��d^G�@�L߆��g��3ر�YG{]{��.0�$A��y��M��s�I>���26`G��~�����u�������J��7�V�k��|���[��Ni�ȂLסI��x�8@���"��|h�R`��'�aI$3G�o�"Hå�G�?Y��6s������k��PO��'�Q
����z+���ݔ4���I�>k�/`3�<a�ժ B�l���茏��ȡ���o"���7�K��NI?	:E�>��d��'t�g�W���	�S�~&"����g��q Y�>���d�$|�d���l��<~]i���	E��>g�����ҡ�4[v/g=YD�	,�Ad<�n�$H�RY8!e?��3�Y̰1dI{�S* d��Q����3�32��U�#�r�s�W�n�p�/�[i�+ˍ�Z�H�m��b�66d��qdS�i0�*�`��p�0�%�R�3�ZJ=�h��I5)�v�E��o$İ��A������i��1���M�Sh�7�i]+���M4���0���B�K��:8��0ۺ��u&.�u
��Oj_f�%�,ь��l�iIN��K�]5IĦe����y��f�,YeZ�iH�L�F*�svͻ�g��� ��Ui�8����ژ�љ�mƁ	������SK�55��[�]��~����'~�ϙ>�;����,��#���	 L�����P>�~�@j	������?�����l��d��� �$� ����L��S#�kZ߷Z���	���՘��zt��۶çtcv�6�뫮�a�.4��WL!x�Q܉��?$J()jZ ?Yq�s�q7�,q�lV�La]5��^\�s��%�u���x��� ���#�>�����[�����@�� �HO�@P�e&́'�,��g���@� "8������,�\����G�B#ﶧ�#'�tca'度q���JҪK�O��?Z��M�B?}�d�H^ɟl�1��#� ����:#��	�6�=^jvkʍ�DB�">#ֵ�p), �LF��"���֯K�>�����}��w7�4�H	�
��������V��?���F�?�f7�H�<@���*�il�.�I�x�!9����"�G(GO�F�}��ת^LQ�������G�V{�}�0P�p1��h�?Vn��`G�~�Gݵ~����K5�Z_T���X�}�{�"?m�C 2+�����~���6�@o]��H�sLl>�r�4�� Aꁵ��<G^���?x����@;�Ϗ� ;�I��5��Ģ��2v��{駚�q�ͻ��&���"�Q������4a�a�%��4�Fa�ٔ�����)L��O�>��P�@���:��G�?q���mH!�����c�ş�`�$}DG����"{�<?mݿVC
��Ͼ��@�L��+�57hE�(��H} �'��4���xD)A	&e��d����+�HG�Q���y�dY�U�]l7oE�<��o�1��0�wx�wi���Y����;�U{�i0۱�c���l�B0���)
�]1�q�1��|H]u0i�|�<�����og��@A���?|	�0�J@F��SdA�Y��(����۲�?}$W>�X���Ӥi�'3����q88i�
�CI���O��Q�>���|H��3t��~�~�Q�L"�o|�ˏ��l�#�~�n����]�4�=��"���z�0 �W�a���b>���ݦ,��p��&?s������5���6U
�S(s;���j��"��H�k��bpϸ���/ܾ'�"&y������T?��@G�"��ŇPn�bH�Ӈ�1�>�n�:�r�^����}��v��V���iQ��[j�i���o�[�N�R�j��#��(�0Y� g\l�z�E�h���G�)�8��3�u�<�>�7yC������?"���<~��(�Q,��m/�1�?	#��Q�:�G�x~�ϸ?��v�)u�8�8,�7]�)�ŭ��٭[cv`�8���-�7f�,���6ֲ��m(��Zkr-5�cI��'����\��<T�_J"�g��{ |\a��ǈ$nT�&ա�nԾ�������S2�l "H�j8��yP�E� yL�G��`i 2��F	%[]�����:���㩉1����|�k��́b���	�0���D���]��+�3��Fـ��qE��K|t�"��|O��^� Q�Տ�<F�Ydxοi��j_������!,�"T���-�n��>�>�>=������jv�@ȿ�,���($�S r����Eq"g�?A�c�4���ގg�O�,8q�0���d*B�	ws6��!��x�9|v��+p,�Rg~��/uVsX1��ݙ�\�U���Y���\{��P?��������Ӱ���6��V�?���>ߵ�>��_���8U�SC�?r�g���5jđ��^J��4��G����O�k��sc��}dPf�>g̆d�ky?��֗�&�b.�;rU��zo��"r?N��0���>"$D1Q�ސ�E �,�T4~��G׻ 2 b[�}Dg���8h��G�3�=�����Z���8� Ǽc� ����?�1"���E�Qu�e�5?}�81I����Ujj.?���8�̾�~�C�@'��f��6q"�k��e*:T�k1��H�Z�����TX[���.><k{�5�<5�aUA�m?��ọVF�?���c�//�*n~����#��p�Z�����B�&����G<~����#+'�T�p��0G��0fV��-L0�,�ڡC�y�mm���_�ҍ{�� �4D�p3�*�>� Z��~^���6��e��� ]�e08�|~� +��Q���,�ޤ�V�4��J#��W�e��:�d�(�	?Uv�(��$���A�����:AY A����>����(�~�Tir�H�[�ޏH~j�צ�(x2$��4��֘�*�~D^Dt 8�G���_ADi�\k\�_�b����>*tj��V�R���}���'�#�-ys����d�P.ycQ~�R��/ф1�|���dDAHG}B@�ג5�ȏ� A��aӕNV�^/f�+�a�b��^�isD�+7:wH�F��۲�kn�PhN�F���mgAb�n�r#-f��س�ji"�|k��%+z�!)>�~��Oeɲ>'H��?A�9}ҐB"�F1)�L�"�X�$}��c��vG�������DD���~��C� x�dm�B�>��uLLׯe����-�裼�N�($�������~���I~3��L4W�q�.vJ&B"Rm"�H������3a�gT�6�����㱍6�[x,���.a+n��hMB[����:~����N�zm����?{���N�����E����H������~���N9[��YpK^��A�(���5�u؞>��(N�'�ߥO-�g��42$����S_i�<B/#�� �D}��n�x��O�lǐ{6��廓2DM�ç�Ez>�yk�DA8�U�C?���R����(���$�d�w�|�6p��Yu��[�������(E�\�ػU����~�3�oߚO���y�d7�O��|~'�/Z^"g���@E��ϳ=E��ch�`|~����Ԃ?Hr�Օ}* �	y>R�hv�_
 3��x�㗎�)�%"R!(1)W�G!���Mp�oj�LD�TQH�ߖR�<�C$���Ó�"	u���W���?|��F�{>i�$�@E\:`�I4���C��=G��X��Y�=�� �E����ck��sdEmAS� ��
4~D�5P(d����8�:D�2���ݬ�{��{���J��93����}�lH���G��#�-�?]���ѥ�<"�S�-�~J��\ig�E��)��ƚ�xyL#ŏ=��Ab^J��am���z�.�;}9ջ���k�������l����v��{
{����w�*�ȗ�ج���3����٣ �7?OϞ���"�� W�́%�k]�&�JY-�,C5 �B�aٚ�](�4��"MCg�m�e����Fg�K���au%���f-�q�:��)l%�MD�)�n�p����r͉Qh��V�n�����9�V�;	���fSF�!a���t}n����⿷}~|�x�7C�Ve�V�6� \iq��h��V�Q�mJ[�3]/k�z>�s<F�iXm���Zn�`�
�����onMl*����M5K�f��q�C$�*��?G���>����}G������"H����� Q�Z�����������8Ԋ?2 OS܏�S�;j���ɠv�ƶ�G��4~�k�q�����zb��[v��q�4Oj+��i��)��KG��.=q��|~��ݫq���/�	�>�Y� �VO�O��� ����"� �AP�kk��#�d>���,��������� �#�G�źb}��x���{�����il,p3�k����O�0s.�}���i��s��D�(�2 �f��8�͖G�"�emmV��V	p� a��'Gnd1$L9OȁD�O�7f�>�^�?�NB+#�D|�>��ퟎ��z�:�L�ՒR��[͇���<��-8Gy��awEl����a�Q~�Di1b(`� "0r��*"�@�Y� ��2D	�!��s�,�� ��H�	�BT��*婂~�H�08�d��S�Q�����'�������I���JIO�'����/��a�����a�&>b&cݤ��TkQϽ����@���(��]H��P��7
@��D��Fz>���������hƪ�O�-���/b�ނ��"�E��s��P���~��5)�ؔ�m���]I�Q��B�8G��V6Q�!����c��K��F(DR�R鏻d���e`���W��|~���q�d�0�=����괓9ۂD}�� ���_E
���'�-�Pg�x���b$vHb�.�����}R�K�m,��R��a�l�t�.	#4��"_��:��[V-T۳���w��}m�V?f�_����[Y����ޥ��o�bx˻S3zgq:���>���<�>���A����]���F?}��)cǉ����*�3��,������D�>?��*��} �z���'� ��}�5�VT9]pC�
=�K4�����/���d��sҐ��:�#�?y��!A?a��u˒>��8���:��$or��;ݡ�����@G�~ef�����쿿G^�,���i�+h�!K���<D�8{#�?Y�(��
�>�p�,/�~Ç�#H'�}J���ޡ�TQ *��,����H��� �O�@F.��P���7��LZ��������a�,��$QC��>����qg�b���"��L�Ql���?|gu|O� �߽�C�(���A��h��5�����ޝ�����g�WZ~�D~�#�>�����Ǡ��G���O	��nߜ[���'���	�")�2Zᰳex�eaՔnnJ��!4��ew�Y`�]D6�d��'U!O-ȗ������Q��a�~�d|����<E�N���ӓ���`��*F��m�0t'�Ϫ{�c"F��a�1"Dj�z~�?I1��F;��l�;�����\�V͆�v��~L���~��0���>�GU�J���^G��Q�!�b�[�SN/��,�����6D�]��W�M�"�TZ" �����wRc��Q������j��o(��C?I��7�q �ILL��Qb]� "�>��&�����6~v~g�4Yn���o���<��d+�rNN��d��D�1h��Q�iNM,-�Χ\���;nv�Y8g�:�lCP�w�is�:eZ���<ӓuQ�eI�ɪ���� �~�^�`\//�����0ɢ(�l�H�<~�	��}���v�X�B�K�~��ǍQ�������:w�aG��k� �=Nl� a��S׊�L
����w����Fv8�g�d�
:>�=Q�yd�4�k~�	3��� ��ן�׫5��������-�R�n���	��O8�0��_��弘|B;1�T<Y�G�t�,��9���Dy��vT�y���#��,��
 m��a�N�4�dNE����G�(�q7�ܡ
"`#��4� 3������3�PJBc�)JcYu5�Cka[lۆh͘��R���B�KuwK�v��5,fлo���2�I�@���#�|��,�]0[_x�<��k�Xg�}&��Hw�q�Mﺾ�4d��}U�ަ�g8�ş����1�W�F�j�����k�:l� a�Vт���NY�˂����c�Ɩ>�����\0�8�k���1<���|��I�+|"~3>����?
"HC8Y$m@]]/��#�Qn�x�<�q�G�~��_A�F��,�̪�ǫ�~��������8w��iA5m+2�Im��o��}�|0Qހ"*@ہ%;6폳�(�������d9�o�_o@�&>��2E�8.���8 �'��ƾh�t�F8D>#�_ր�	^���}�=��?}�����<O�����n{`��6-ߝ?�ÂLH0��4Tǹ��"��}�~��x|��y"20����	J��.>�?x���~�۩b�G�װ���[��[��KO��3��L˔%�������B���@��*i����Ƿ���K]���7���[�,-gM�>v_]����[[���wE����p��L�>��_���K����otI�)&:��?},�?
G���O���J ��E��F�7;~�zB��1�H*'h�$�~&\�9����/7_�ϖQ$+��'���$�o�ߛ���4�nD�j���\Q� �"d��%�D_w�O��ߝ��笿��ԅM�Y�XLCUѠl�-��M@6.��*�ΞV���Ђ��L|Ȃ	>��ˁ�IGyGϗ�ĉ�,��R|>���0��?�A6E(�O�>����i���?�X�������@��vD���B~F��}�J��I��T$^��~ ?[��6&�б;C_��kw�Q'{+D�	FL�A#N�����9�ǩ,�F�`���C��Ę z#�3\�tD@��|>?��Q�@:`x�Y���xco���"�;,&b|d|I"!	@�J�_@��$Q7Z0mq�~'�2���މ���$ ��@����&|S�Ϥ��'����8�'&����� pE��0Fޏ���{K�q��R.�2@$ײ6߷��/:���jz#�p� y{�,��/pO�1E��ydb�Ce]��Ȉ�	�H)(+7�w�?kw�]�rs��:��]U�d���`A��u7 ������^���_n�lس�����]J��:i��^ڢ�1
"�,�8#j���>�!�D�m��Qb#����K0h�F�R�_b9��6b��^Sq�����@y�����l���6��y���@��70=�|��xFU���;�X��q۴���	۽Sz�V�q��W`��m�n���u��L˼����z��"�lg"��S��꽳��ՙ�8U0��ff�'Z�t���
��f0M�/DKp�����)�l�h�51��rn���Wk;>5�toZi�l�3��/�[ܷ�t�����M�O{��8v�A�7]�__��#Q��݋��$t�Lw��[�z3O\�jv��ml�.����Q��wj�\��Z����qk5����u�jޝ��lV��ohn.�IL�bv�4�;mT���xoo��%G�j��.}1)���*����m��v��H�|��L����dL����p��q|�<²��{g:�\YCR�ɑ�t����#�ί�F���r[����
N��9�Sg8�d̾�%�q��@y�7�	�ت�0խ/������ZX�S}�ާf��}W��*pȝ�'fU��N�l�w��i�����O�a��8�P^IK;�؃���$T�w.�뺕��-�#��;z��F2�%	�6�[K0�Dp����x'��heܳv�cP_^d��$1M��.K�`܌%���n���@��/n��7��gl=tʊ�ڵI�qQ��W�oEʱ��f�����,�R�� �g�q%e��::��b�	���O�iCV9�ӣ�}&9;wJ�B�o[��l����q�c3)�˦��2�J�����o�Eْ,�rmX��f�)�z�����YW8^e�Z&��&��n�٨[�0��q����$���>����w^��mn�`-�V�%c�u˭�������Ս��«us�T6�����k���,�1��7E!�-K@[^c��,q��w9�e�JE��e�;l�v��4��uI��J�݃:��Қ͔S�5�#��]E�&�����u���\�eX��m��;)���}.�\��kc��F�d�1m�W����]7;l\C<U�- ��ғc�a*RS�4��amѡic����kR�k)1\�2خ���e�`��v,)��0�v��P�\��Š]��q��X�]��(EhR��5aoQ����o{D�܂AD�ːu�,Ytm��5��.a��45��6�З�h�[��_�oy���k�&��c�h��s�hT0-�Җg;`�7�
bju�$�5Z�Qٵ-���Kn�ft����N��vf,e��tv�)�u��vv�V�]m-����T�[{b��$.��3֬�	G46�5٪�z�)�kHRj��բ`|���q�Mm,%��R=i-�jL�{v�UsA��ݪ2��Vmt-�K,i���-�8uw��g�۞��i���Z.Sr	@��D�L������W^�sc��]5�Z���D�������e�*�M
+i.&�ҧ��K���2�V��4ЍFll6�Rc"pm���ԍىy�f3d6v��j���v������EԴ�{�I�n�ī���<}��y�O#�h}}�[Om�M��|�GJ�h�RҰ�k���� tt�%"�v�4ֺ���i��K*������{�g6!����7ˈ4|B��lnl���3�k.���95l�a���ɛo�M�J�m�X/��W2h�u�v�҈7\l&i=����%$�����=޶y�����y�%f�����&�[�X\	nZ���Ck�%e�Z��g�jj\�[�F����B��֚]2�%��.���Y�ɮ���MMrSh�ųo���.�X�X#cc�,��aĩ�Ka��c7j1�j̒�dt�fڦ�K`�Y`ˍu٘����m6���r�sM-�I���vB��*�Eh�bl��
�}Y!&IOl1���+#�i*��z����	C�QNx�fe%�1�y��������le}(9��3�#��K�\k-!���-�n�$�me�8��WvABmHۦŸ�"�H���,������[4���-��l:��)���6�՚��X[����f����� k���8.��嘤���HSSBq3&�t���8��n�1�L�3^m�`KJ�.5�J(�3�-1��e]���	��U���.�f]ֶ��me��ȍ2{�#�tH]N�i����0�f����F�9x��~G}��/o�9b�<�M/)�ϻ3���]�þ��!�y���;/u���E�W�tQ�9B�{�~���))nkX3֮b�"�0ϧ�q�2�j��](�^�z�]�x���.��D����q"]Ĝ7~�̣m��^�����_���7�)F���><MW�gei���\[��eOp���"NTYD�>'eȤ���W�:yc��k�9XؿGͦ�wj��QF����^ѨB�,�0Vf[�o�䜱n�O���7��^���>-�NF�溢k�Z�sEE>`����:������Ң`9�����j��'T�����鸮�co�")�)�������rD[�3p;�[G4��@���M$=� /B\> ��+���c���si_�o��=H��{W���f�*4���F�	��Ej!V� hkuu�30�V��au�j6�-��pkn����@��o���lH��ło�lln$#n�L,�[S!���J;�dT0��bW��
�H'f��vڑwR�����mj���V�����ǻ?}g�����7RWݹby��jU{X��4tW�#va�X)����f���ٽ��M��ҳJ�s;,�v͹:��N_3܂ǃ5�ܭ�/�vk�(l�,���绡�g�b��ز}ff�}1�tm��=��di����_w��i�#�8yk$�#==���	�F̶�@d��q�yM�P��-������<��H�w��v|�G>��R���R�ہ/%Je*���7�YW�Q�[~׫�8"Q�Q��;��q޿r.<����*Ws�-�P�Uu���u�:[�baRH-�u��<�X�5{\�j>3B��>�.�D���;v)G�ۇ���
�es��P� 	m�����L]���^���V�D{^��̑��^򯑹����o�[S�� �U;Ë�3�:���2�ƫ�^���sF�Q�Ä����o�91A�K)2�(��&,�im�.�b�J�X�1bh�1v�S[.+�毀�P*��i��c�����3ƨc��8�������`Y�bs)ӵ��{/*�2����ݶFмu@�U �y��s�6�Zk�3l,��0q����)9u�w�����p��%�Q:e�z! �� �����<�Jù��I�l�Hl��E�."�J�x���ݳ��ˎ�xp��ޜ͂�J��R��Jp�E�B�
�B�̯F�Jt��!�;tW,A�雹��<�PJ֪�6l��wK�����+!��êZ{��t��^P�8�F:�}emfk�8���]m�YQ�U��es�S{zwe��UfU�����y��Y���j~gV͚���+g{}f2���H�)I����~ �R)�a����5ʥWT����l�EĢ��������r�ZtI�wN��]!A\1���r�<ؾ���e��6������|��e^"`�$Wc��	�L��6�k�^Ԏ���~�E/vm�!��pl}��6x���B�q�`�I8����W]�y?*r	�o�:;��UF2d���A�G�~����_��O����(.�(�B�jZu����u���<�jsl2.�j��0\2������ζ�yƍKP�m����GU�^Q5u7�$\�F��h�O�Q*>�Κ�K�g��Ԛ�j�U�5aU���sk�O�׶��Ƽ����=�ٹp�I�BM�~Ō�j���U���r�T���� x��@����ef �o���z���/_(zD�}��4��kH˥�>���b�M�"D*7�w@�0�$B0�J���8i2(��ZE���.>��SW��p�p�W�/6�t���\��H����"��?U�Ǻ������y��[��>�<?��1���r���w�xE$$����1
*��Ⱥ$䂕��`٩g���bϬ�E�֯�M9�^��H����:16)[�WW�=��S�����׈��)�7���j������y�����,r̬Ő��'�]��۬]Q��aw������`sn��c����c�"Q�`!�Ϗ}�ϗnTɡ{��s����l�o�^�b�3�{3��BԺy�E�*(����=���cգ~�Ի)y�yr�~��~D��2P!Z��K��X�e*cT���]�2�;f ���%-­�\����O�]Bw���/��װj��;��Adju��es�%OZ���'=�j�k�}Y������Vw˾�K�)F�BV !�<G��;k�|�gMl���yy��u׳}����6��f�o�ߗ�	_���<{m-\���cB�Oգ�ȠN�)��\4۳�
��̼��{T�fK�E-�qNg����o��w~�O�6����tV��|&�*�V���Y�u��{� ����P���ڡ�J���M�6Vz�6�I��\Gw���1��jz돬�ˣ�s��b}��c�W��l�$R�$�Y��E@E�6Ϸ�+�������Ū!�_}��̍�v��_��{��"��7�����{3��:��(��6�B�_v�`�;\&��*��X�#�<*'�+(0�3,$&��i��\b�p���n2.�ls��KFC�;%m;ǿ��4�a<1����r��Q%cq"T� � �u��29�tqt��#{����V����K.���[xv�ܔ6$w_�x,���A�������Z��Aժ�l�ٍ��I]�f���,q�4���V�lvDU^�[n�}��� z�Qy0��X͵�cvx�;vGZ��mu"B\�6��4�h4$�6��h�V���j�@�M�F�n���e�9�:�Ё��13f`L��h,�1�m[���my<�Y{7Wv�ڽ��Ҳ�,vnm�(�V�&a��\���+srhl�RP`BI~�;�����j�.�_*��[��w���+���9/����u�Y���ތ>�QM�"P��՗mb�Jar�HJmP%�SY�sq�r�.���q"����O�k�F;��j��_j��Λf���"�)��L^�ZD����_fn��I�TiSQ��J)��H��tw@��/D�{Ê����Fwsxk55�����平�xtNnzund�w<�����flL�)��-�,Y���*AI��Mj����m֍�47�3����%��vT&c�;w3��1�;��l��n{����a����~bGS�sG!�����P�"P��oُ/���j�?�����M�ܭ2^'�u��zM�}���ǩȷ��X��˫��E�i߳����>�,��Z�vqul]��Dȅk�n��I�Q�1�aie��4f՛]5�����4�q�
++p��@;���4λ���l�s�3��Q�f�Nd���w]�z�tj�{�r7�:Z��/�ٔj}��	��RcQki��D�G�%�`J��m�+%e����:y��W�=﷧|��a?o�s?s�b�u�����n�݀����L1�+n�U�r'�ʖ-�7��}�����Jn�1*��;z��)f��R�<խ��u���>�(<��6�G��Z����{����xQ�$�T��K�{#���9�\QxRђZ�Dp+�g�;3:���}Y�l{����0g.Uoy=39�|(<��dl<-._w�N��R���ݝ/��������Y�7s$�LA�2�/G�<I%����W����Il�[�U���PI�@{P�n$����]�w�׻7{{}�Gދ���|7����n���` �D�Yv+��pp�:4�����ǡ�D��!��̛�w����T\/�}�d{Cۿo�_�>�vH�	��~�M�ܸ�\��4�0SFnH]�Q5�RKb�)����	[���2*�*Tܷ,O�o�/Ӕ��׳���rz�����ɲD�	�W��򠆥J�?c�z�dǣ`�w�G�AD=��F�/sFfX��/LJ�Z���ֿS�>Lu�ã���^)�d�|�?nc�N�0`1׻W����^����.�L�.��o<��,�xg���CL3�pQO)a��4�κՄ�7�R�R��1���G1���R)+����Vv֛"m���
��x��4l��/xð�D���Γe2[궟;Wr~76]��W���l��>K���1��+�w��ur�Z_�ύo�.��蝄|s*%o{0)�!@�$!�X4R�笧�ۤ�s�X<V��wb"�Y��ӝu�<��n.�͝��WeV�F{=}F<�ͺ�:�n������n��}ًO��7��ҧU�ϐ������9u֨Ŗ��D�9�˴����M��ZlEƉ�g�]��}n��{�S�h�}�)��{/ݻխ6�1��F����b�M�1T�pFl������5h]��\�pY�bDb�J�Һ�n�����YP����=ʼ����{VW$��&zT���t��V�,�6Yݭ��U���{��G��o��(&��
v�u�4"����������<�->��Lie!��>Y������Hύ���pQ�<v8�{{f�녈�=;�yN�1Q�0�m�%m���8<j�L���~N��U�Z��Q^�c�X�TJ8DOq��+�Zo���ܚ��/=i�D�!ٍgJ[�l��_�:���i@� ;��+6���{��W%�an���I�o?�0~���#�
�}x�&��+�j��jau;肩ܣ�x*��B��R���78�r����ʃ��LX^���w�]Gsjiw$(>�؃�3L�B1&�|5�I��2�7a�`=�7���=mxQd/;�iݒ��[AB�4r`��~g9�b*�Y�	ot�Z�V��$iFo�{�ꯧ��6��g�}�ν���ss�o�l���Z��5��������$�J�R�s���k��/l�a��fG��f��Q5%Պ��7M6-�F�a�����"� ��˝��5Q�PI��WS�$�o��	�!�x�[�{����*�3��J*�"�\��}�=!!汗�]6��R%��3o�
|�w}�7��]ߣ#Î#�!�0�m�0̻]J��[ub�c��E�YąD�,��?C���!:������!@��G�dJ��(0bG�T��)��Q�"0��S��aɷ�\�L�pg_����
�#/�ccu'�u|��>鵦�ي�,~ͯC+�ܽ����^�;���9NJ�"��H�@�vx��\��՛�+o�nO�}�쌕��z����D_�����=Y3j���]�1�o��s��,����oob�m�� ���__sF��0p�K
�
Ԑ���]�{�w�-�����L�-od�Ddfo;T��/Cp���|��N9�t9��^����8����5��F׏;g�A��;+%m�p qpW[{�]=�qI'뢦����;iƫ6#9݃Jz��籁վ�É�[��l�����冶ݓR��+���X���k��j��5�1��]��΍�-"m7pɒ�I3>��ޙBj�*g9e��e�he���"�F�V��U���!R���-���u�ڤ�����y[�����%l��@F"���R�X������z��B��SՔ��d�����la�aek����,[�#P��h�g\�^a*X-�u��VTSR�p�e���݋�
�CM0MS��3&�����lЈTc���Mش�JWMM���E��(f���YWmY�{��Kns��������T�HX��8�5����K��`AV82��E���w�vX�G�����D�T�4�[�a�Je���zz(c����	�/���X����Ў�
z��Qٓ���㧶G����55�WZ���u����N�����0R`>rt���V���R
��r`�a�o�lvg���ڭG齔\w�,y7y�F0��wPѨ�`Zi��/)�ܻ3���m��?o4�>�_2�Gk��*vB�Z�<�5%/�Ρ��>d���7~�9'�T���ȰPְ��+�j�.3.*��kueNuf�������^��o��5�wj#�Q�RA�i��&��3�h������p/r���Gp�����߇k�V�h��^d�X7kyS􋕕ْs3���BQ����l�������5���fJ�2�g���R�e,J�d��̯鯥}�v�*Lܬ�R�����,�s���m������Q@�䮌J<~>����"z�zo��J�R�uQh�	��w�x�c��}4�"��Jl֜y���P'̹�%r�V0�� 0׳&Og�Kx������z}����u��I�+C-�)t������Ō]�b�����0p���&���˶(�t�@�a�bZ�Й���F[�@�!�����(��;������ٔ��]����J'"ZǼ�X��1~���p�'�6w�H��'�Ke�J	�߮7�{*eae�vs���mor�w�L� 
�y��C�xϣ��3�}۸������V��^B��my�����2҈_r�"��SD��2��A%��oLa/��L���UDI����H\��{$#����`}�٬�I���Q� ��F=0:�C5�3�ax��Qg�LN0�7ᘥ�Mb�Zj�SB�ogn��d���ouu��Ω[�s��(ו{8��V���z恂�+X�)çz�Z��Ds�ٓj$�sDތ�g�{�K*�I�+�I�H�! 
���k�]�VK���6���iq�틇��]��1�e��O���S���"+w@_���6�e�dE�,�³���}�x�����ު
n���f�bjf��g}�n3�YSf*�Ud�w�������v�>G7�-���Bs=���s��
��Ů-�{���^˟c���_|5OCc�p����X˓�Q纬���u�Y�L�
�L�)�5�QRf�~"�.�y�0sd��Ɲ5�o�o2�c�'e����7�H5Ӯ"v^��, ��v�2��_͛;�{���FHK�-W+3�y��SU�˭�0��J<	�Q֮;ܞ̵����iPA�'�pV$7`Χ6~�ٺ5ov�*��}3l�-��`���$�M�Y�Tu�7�2�˾�	mN2�4(wY��.�C3���t����c+d�ܽB�s�7x_<�-�4�Iۛ���,�9������[,YW���ד^�wGwu,�ңb.ի�H�!��BQYQ��}�_�G�g�+L[t�N���R��[�gL�Ұ��.6�I���;k�Ckr��u�&:�b#-V�j�9wcgv��o*y�I�[団��b�`�,�˓+�#�k� ���v-Z=]�qv=���;��B���ƟoBr����k�x���ZІ����K��,.��\��εϨ�{Vneղ�Vec��9qIĤ��kɹ�Y��rסk�"ke �M����]/y��]&��F�ݙ]�v��a4��Y�F��+*0
uq+�������R�D��9��1�ƌӷ��ux�R�6����/�X�挳���˹6T��EZ�+r�os:���w���,�dYG;���բs��b`��n(�x���v3�U�S3X�*RpTS�H��]̧O��ԨY���kW�
�|"����zD���X���\�S���݋ʂm�(3��Z��9�zy�r�\y�sF�wkVv���abͮ�C7�/�����H�=��o׵��cS�m��wt�:�����9oy�v��h����O&�@QG���.�?��=�}��]�F]���Q,A��<���nV�b��R"l��w'�{�|���fОduπ���>H�R�K�}s\�'*�~x�~DM�h���z�Փ/�ݧ[�"�/[I��j��	��3̄�7�����
���Wff��d���8~ri�A}����0��W����9��$i�5�~S9�Y m_�0�6}���t�\��)��%�XHV�c�՘rm��!i]�*���]QИH�`Iz�%�p@��FAI$������h6��?��֧Ҏ�����컋�u�:E���)9�j�{M��~^��sb��=�"%b��)i	��)�y�ٙ{��|����t꽠��M�L��z����N�}�[}���V�J>>�{ ��g]Ds�5�z��7|��x��P�������<�hy���h�����Tע"%�sPP&��'[��㗥� gn�e��T�0zf�7������0�Ð��un�� {l���m�ݫ�'�[�j�Dӂ��iN{\~�]��ݘ��35�D�l*�{^^x#���罊�w��gyo��C�*�ԟ����+{���xM�#�4�*�*s)��tr�>���To
�ʶL7[e\�xȲw;њ�{��6�nD��=X�ez]�o��_���d`ɣ��Ђ���J13���XfU$� ���1g#-י�o����H0���ͬ��ԅȹ�o���%��Z�����u�/zmN��h#�����7_D@X-�n�|���3�*1	�Q�0-�wVW:`tp��͙�me
�����I`�+
�#NﵿI��u~/��=�Gq!��e�\�o��d�Լ��D���.����)vA��ڏ.�4�WZ���uT�֮t�(؃�����`>�g��5�s���#�/A>�1љ#�	�����^�ng�hA�&܊g�����q��^nK O{�hns�ΣV�	���7���Z��I��n�k0��B^�>PT��y��=��ER,�{ʪДh{���WEg�w@��})��{6��(�vG�*�<=�{�I��Q��u&�Bd2D4��,�G���VC=K:/wg�R��"��ʽ��f��х3�Gܷf��1�ߡO����b�K
��g�ohk�폛S..z�no�UpC��YCs��&��b��s`��2{H�W����w�:��릘;�$l��QDV�v��a
�ja.��W��F��q���۶Ƙ�Y���3ZLz��R�t�p�yxLhܠt�F+7�W��6�0+�𿋶�9������9k�P�\_��ϛ��k�)W6Z��.׵��F Z�M ش��䫶.T���n�vt�hX�ۮ�A��m��T��S\H�[F�d��>g�V�l��q��.�� �[���R���f�RPҦ�qi5X��f�3hBl�r?o�<[mHw�%��8��FU�.pd���	H�pĺ4fS:��oc�H1j˓B{Z_��1�u��v�k���]	��mf[�WWSd���u��ZJ��̴�ۄ�F�l�]U[2�6�;��LmO�3���S0���{6d�0�ڳ�ϗ�\[�3��t�}�I+պ���Z�����̞5yޱ�%J����څ}�^��
'd�Z�]��tWP�vɨ���d����]wL�-g��������Y;��F��Q��TX�����\��s-����O~N���y�_��(�����j�>�1N�b����P`�m�S��y�Bj?�)�hko|8j�qc����J�˶���%�	����a�K��`�2aj�����ȬB��Q�]��s�;~V�#��$�������l�Hɦ"2�㾥V�y�T�	}m0}qW�tEZ���N��N$P:V@���߇"��;����p6.���oQ�\a��Q�ᢰ��Y{������T,�����3rC��.g<+L��Q!��Q*(����?�����F��<��&+ �`���>�WC��g��)�Pq�f�u5q�SJ���i��9�����$κ�ن��TI��!Z6����3�\y�<���=u�CU&g�Yz�
�~A�����?J�|��%-XT���N�}&�\|�����S��D�n�>[,o�&gD�,Q��wko>�3<�~ҘZ|?�� �w3�)�}�ވ^� �����IF�q�Mo`'�c<]���ǻ����tĭ���mKJ��_wVv٤oj&��D�{]���|-�hq���|��	��ƻ��n�l{��\�j���H�E%5\����1���V�5Z���ƫ�=�ڟG%~�Qm����������9�}�������G�J�|h'R�i��q�ٝY#�e��׊�粏��Uzӵ)��m�?g�����(�`�3.^}�5�elDWw��a+z����wm��b�t�7�}/�P0~�F���,Y�T	5H���3ޱ�ڴ�Zjl��4.G�ɿ>Yo����Q���RY�?R?��|�Ю�:��|�G�������j��c&���{�^�1`g�F�)�}�}��Q6�f�w�uR�Wb-+�U����pB�Dn��M����w�-�]�a�#�v���w]��fk���~j��r�G��ڊ?{�6��O��/L���*ʰ�s�>}=��}�aM˞�b��d���0ϊ8B4�E��S�PR��3��mi����>��b����O�}}��j�w�z<&������_k�i�?Qgm�k�|�$nJ�<�=�(,�͋��w�<r�wG���S���8)%eL��͵=�!�LZ닪��5J�a�=�J�I��{����L&l����R6	6�i�K�����\�-U��	3C"�N�on�rò
<��J*Gb�]F�i}�W��:+ˍ3m~%�}��J���~�j�ξ{��מ��L!W;��tDꜯX���Ո,qB�%��������dl�*&�۸L���,T�W*nך��n�]E��<��.��/WNޣ�~X?{ԙ�Y�Lms�c��e��='�C�^�@��?7	��s��8TX��v:�9y�,��$kI_Z��'S�f{�gu(�~���J):�lnK)����{��1do�Dǔӻ�5O2sY���0L]'��ĳޥ=1uƷb)iSr�ڦ�Z�2ke���m
�� �ӄRP������wE�w1��S�5�������6<|C���w0g-�C���N���UU�>�O����HD����I�3"#0��.Y����#�#ݝ�>
�5t�q~���>~�̯�©��xj�%��ӱ}
5*,���qPz"j�zp�sK��oR�3\���A�Dݣ(+�>���H�&A\�/�#����I;ݽ���{;<�<���O��m��S�SN���7b��(�G�u�����(������Ю�;շ;�~���\���6 w��ϕxÏ�GЮ��r6<Rn���*���~y.����K|<�W�ô��Y���{j�N�苊�h;b��^��e�ffh�u7Ok9�u蒚ۧh��k���K��B�[�\�ե��{������٤դ6�^ۯ|1�~�\jb��g6���>9�r>�M��o��6�~؄�4v����j�����mͥPϣ�|.p���(���p$��yG��Y�r)@ꆫ��o���gʘ`Vf�5���n���$��6Z��M�����h���C`��6��oo��0��� ��_Tž^F�XE�̚�/z���?>�Dmu�~ǔ�C^X�ά�^��ǚnUv��D9ٿ*�e(���q}��c-�0(�������3x�=�+�v=�5�!�+�N�:W(2YB7-HV���h�K�<t�EeOۍ!}X��2 �z�!!���
:"�y�e��G��
wK9��R�����;���>�_
�X(~G��F+a�����8��e�)T@���4,�z��:h�u[�ǁAL��!@�����8����5U���>�s@�K�s��.�}��&����@^B�yR�w6�<~~���g�fa�Y��j~\�)�4&V�w��@����?KI�^>�ʈ�V�+w�3�����$쾕�9�\�z��Y.�G�����f�F:��oUWF��|x"���W(�C����
8�Q�kW>��&Y����yy�m���8b��Ҵ�[WI��m�F�v�<�t]��NJg��ޜ�:{��[��s&��Vm��hn�mg徇��mrL��c��2Y�C�hK�e1z��޷L�`����%6[�V�n�ۉ��HP�fJ�K��������&̮�6e�M*~>���ĸs(TMMc�3v
Ji�3�v���(f��[�O8�1uk��pS�+oha�6�:5����If��*;Ck��h[M9h^���^��f3,�i���-��J�u�L�f�a�c�aA�.��%��n�l��۳�3x�s�^rN��`��Yf�u��\G���JUi����m	<�}�������}8����z�Q_	*c���Oۦ2.��g����=�4q�S�޷�w�i=no��)?U�q6YD8���R��wiO�� j��7EWg(Cg�������4*����}�Xo=�
�˚�f�a���ߠE����c��lK��s��;;	��ב�0Q�R�e����aČ��%k�f��#�4��d0��˂�������5�S�ך��7e�C+��:��N��U+c�+=��n�6��{��$��L��R��2��I�m�u�|�>5QD�Hh^����{��흟��ܝ�O3|'zx��f`��L0��MoS��D]�Ę6N�0��VPo4b�~Ju�}９n���s˳�ydk3?um1�|�y&�����1J>��02�֩��,���&�q`�-[��;��̫�Ox�:ћh��Y�uv�Hbs`��j������;c�X̬��-�Y ����%�s��'�a�g��U9�Lr���j���g��2�wu��J=�0�F8eQ��0D�Q�2�)?o�|@��(�\2�b�A ��f	M�u�jKqYK���0�{�p-�1�#��D��8 O���w.N����gM��|֐�*�c�"@��Qcۜ�P�z/K8�;�3p�)�N�Q��܀��GH�_?����v�Z2��1Y�-ԋh	���iz��f}γu|�����x6ŧ�}�1=~��!w�����T�"�uu�Ƣ>$/H���k���ʏ�ސ�)׳ѹ�#Mf���dT�L>�^"�q&tL�ڻ	��#^w�q��Y�{�������`~�--?:�?���q�>�����U���x��"_O��qgO��|�.�`T�ڋu3]�$���=ܧ}R{u�zZ��D��DA��or ��%)�S%%�p�?Ml�Eu'\�	��f�Ǐ{X����֧�� ɛɻ��F����;�lf��naa^,?x�����D����匂"&T׬M�*M-J:S+�i��͛Z:CpBi�]5-m�6�J;+)-��5�����!7��9xwM$���NfOea]�ܕ�c��]^���sǟ�K&&��� �����.��&�rp�ݱʯ�A&p�$��3�*����xu�5��q5|7���<�ݚ�WvNf*�7#v�[���#!G���Yw�v�)���簾�U1N��p���B-�[.��U�H�$����g�˔@�P|�ȫ�j�k�_23�<{c:N
��ȕ쁍�9��y��f��ܳh�ʙw!h<��a��`�F���f�Em��J�.m�\��O�_�v��/��R��>"0{/�d�g���Hơ��ȑD���"�3*V{έ�?�n�����"-Of�i���=y2~f$ܢǼ����k�3��ֈȼ�K"|T�ri�lP�O<:+_W� ˟����^��HL�A��@���R!��_1חJ��G'Ѷ�n�|T)�J�W�s�=��s�M��Wme@�s���%>�΢��
7�>{qܯg{*z�fL���Z����O�&�k4��j��[6^��1��A�������s&ZQЙs1p�뀍��Q���_�6W����j�4�U�[���F�cv�Tz`y]�����7�&|+m�����+:�1�@���!c����,�!h����_��{��K1�~���I���S�Wצ��:�yy��2}��J~���x�VY�u�� ��������z#���˴�Ƿ�J�u����`o]v���UMt.���^���Xb�ڌ�b�$u�z���G�p/���&Ԩ��c������x��(I�s�]�3=1	(!JI;?_�y͊������~��2�{����Hd|�ک�c&3IM>�D�Jk����l�{�?,,Ѵ������y%�_�-P#���k7�V�og��f��ⱀը��
O:��w�a���1];e`��H�5I�Ӈ��G��難w�`n���}��������gb��%�9�3-���Vmx��!K�:��/U��d�z�~�'7�S����n�}]tdlW�1Xk1��TG'O�א�7��M�
����3g9Ǟ h�����4�77M-�Pԛ7�;��\M��	.-u�~y��씭��Øm���O�h��>U��~�m.f��+Q��WP���2~�rզ3��E�̎��1+`�UY4(qr��"L�d��|�~@��@�hތ�0�e9�;5w�߹:y��ѥ�Ы4�l	�}����nw�,=�L��(���[�>�k�!�W���ۦf��.�QO�;}< I��_�ڟ��D�\	��$�ly��w��Tl�Tz$�6�m
p���)����Y�oz(nw��7O���n���@T%L	�>�}bqV��AR�}΍OE�3\���{/̎�/jz��&ō�D ~�&6/{Պ0���?~���s�Yzd2�N��c�[Φ�3/;}�4}xe�(��3�K8���HՀjr*�$g5t������Bo�}Hsbj=�TW���9:g�v���}�����E��\�u1��>D{>G�1��j�Ù�tT�����]0�����Ĝ�y��� ���;�/s`�={�A)��c����y�S�k,���<#y��]}�Q�=37��Vl �2os�6)��q<WZuԘ+��N��j3S�"y�� �P0\%��jQ]S�����^�0,P�wu��D��H3	@���H�ZUpk^7\��lf��<������Hm��w=ް@o������_'jdKD������G��1Wuػw���牥Y���ݻm��=��`Ld�5����<�(�#T�A}ܷ�}�2P;i�+n�Z��'=TU_1R�sCdJdG/.�����'���c��6���3��r��°D����(ؕ����pf���7�.,����Uwٽ��e�..Q�80���0��H�u.��Α���i�V�Zș��2*���cQE
�O� ��I.Nf�Ex�N[a����M�����0�d�e{h��ͤ�17��ߙ�5���Ѳ�l�
�Au��d��t�m��='��Ρ ��]{]��:,8PӼ,)R�gB�������+��{��ۗ�iX��J�b�3S���p�F&[\�;v��5�!� ���{A=�Usͳ�Ac��Ɩ.�fq��h+$��t5�VL2fm�-�Z��p��X}c���G�.�wۂ`mQ�V�:�_N�]��[;�Ҩ ۺ�����}]�����ʃ�%2d]1�е�b��N��\r>ͽ5�q���z]l\�&�Z[�u&�W{~�c폤m��dQi�ѷ�y��]Xڻ3*���U�ٝn3+�1�l/� B�Q�m�V���c�Ε4u����j�H�Qn����{�٭��E���fF�qe.4��.��"L#2Ү%n�	`J`��@V±a��Yɰ:m��V���n+��B�fnʌ�-[@c����[@�5��cWf\ �Xi�UXf�ik��>�x=V���Bf��٥�K���Z��h7#��C��1���S\Y����T�9�>��>���ǣo���>�C�iCR��V˂�e\�!@�.�m��7Dq���[EΠ��k�w[l�
i�Y��[�`�je69�mY��4�Ks��M|7!t�e���U��`SP��� ^�vi��e�b�p�[3���T��a}p6���{�x�/;6CM�} �x��٘U�A���Yn�lM0�����oS\���:Q�X���G'm+M�H���V�b�.p�˫d�y�fj�$��ƺ�ne�Cج�'mm
愄�ִƌ!�5��)�8����س]p6ݑ�Q�3�gX5�܂̤
�[a.�~딺�Iq��ɫ*YMY�[�=Ynq��!�lM��]j�d�mX�����D�S[l�l�5�oo��V���\u�e�/�c�d�ف�Ɖu�7ZF���A��e�5)`͔�ʅ3��s�KB�a���P���RV��z�ctrWԷf�M�x��R���/��k*�H]�v�-��� n:��QP@��[͗[*Ke>�Ꚕ���:[�kp�Y���5O�{L�#������a �Ѧߍ�]*�Bӆ��j���%�-�R�ѿ��������E,U!���ˋ+�M[]�s��E	�"rk��wR�⢆~���XA���6],���5n[(4�2�v���i-�f��n��'﷉�\pC�ʻ�m��k(���f��E�e����e[n*��E�c+���5-&ÛM#�����s�W/8�6�L��f�D.�K�5��µ!�8��]�Ɩ�XL��h)v+.ȣ�h�vA�l\��Ttq�H~���TZ�CX-��k1�`� ;m-�[�
Sqn%���kZ�M��,m��ٰ�B�[Me�*�G�^�9����\�5�J��V8���Kq��A��sH9��tҲ���sQ(b�%ƕ��%�[�Y��Q��a�5b�����v�]3@��Ƭ������ZP�����@���G��	c�[�#����K�E�����R�j3[k*���m��)�Y�ߗz��7�t�n�1�����U�D$ ��R�JX�R����0jJ{�E�ߦ?��c
��f�O�;�}P�/=?L��y}I��!�B�r��H���{�\�3��8�gԐ{/<��G�p�sɵD}��~N�*2�P��{u���Ǜ��o+��&��_X=���tx��*�q����Kq]ъ�X�L�1��W S�����B���z9{P�C�n(`��I u9�{��Ḑ����̡�����̍Y����2�`�g������q�W��3��}d]��f��=԰U�^����ܺ��#�f`��*Lʘh�6�'����h�����9�˽�{�e��?~��m�&0�W�]�N�l[��O|�ó��K1�g8���xy׼e�sχΌ�ޱ�W��?�b�	K��~� g�E{;f���I��A%5���n��0ǣ�Ea���lm)�g�h2�s!������'��I)�w�D��k�����"�O��-�M*����SS�ڕ�im�iu]�Ǯ�]H�Y�Jg�ڬv���EY)�>�����v.>�R���+�L㏄�26&�=>o�Q�)n�}�=�>�V�� X�wf��Da��>UY������ʼ�X��ȱ;B��f��{��A��>�������fb��pTQ{f�$�^��sYR0] �xU�`�����)gD@m��ݣ�|��eolK�8�!��3��g�4�3՗�[<9��w��)s��g��N&�*�;aȀ�+��l�*����tyȑ�p�\���_ݎ�W��=~�u9P���y���Zy�vwk����E���͟k9�W~"z���= �(�������Nt�bȳ�r�eD3�^�� h�p̃�]	б�J<i4�d)A)+��!�x�v�[�6Q����w������
��O�p��X�kD_�/�����{M�Q��$��ȳ�UhN����B��[J5^�d y4� ���y�{�r���X�G�Y��1���zتP���ozb������x��g�o|�)˓���(Q���c��3�F,ZÚ2�}�{܇���eNj��V*�K�Ibn�ԙ�{Gb�sf���M)z�^��V9,A�($�Kmw�#"s�����{��飢�5�T�͵J�Z���Ä��s�oh�+����cκ'�=���;\����U�\�����o7g�jw���i>���pP�Tʔj�c_B��iګ�T�]�^��&e�}��z6Y����+>�2jW��0>���uC���l�T���os(z6Q�\��z}CO\���$����a�Y�ǌ��O���/^��]�0�ֽ��C��]uډ�Y�R��	�	�q��nU�x%�����F��_��phCn��뵷}h��Z��.f�7�N�ܯ���́��,�k���v&�_K��qt��Y�a��)W{޿2���xS�Y�ªY
���mf�����*T_I#����f=�^�\0��I<�MS3�{���yu7H���}��#�L9���d�����Z�r��QU��1ͮH��]����q� ��Iq���L�X��H�nir����`���D>���E�����~̄RaK�W��B�:��>?*���,6��Ct@��^�{�#�e=S���-I B���7�-���K�b�v�[t֗MkF��K�ٺ�Ю�2+H������~��5����޶lD��X���wm}�t��=���]�t���&�DX�Y�����m�@3+�T��2��$F ��uo2f,��fށ�C���4�A����))K�Wj�_�+�9;�Wڝ�	��j�����12p��ƔD�>Qf�˶���������}Ͼ�=�߮��?J�(�ZJ]��~�UTN=�UK`e/��ʹ��|]�{�؆*w{�#��>nv��5�z|�3[�X�l�Q��I��p}�GF Q"b"6�f���*���f髜��s5�e�)�}������!-��\�t?vJ?v)�=��n�T^���~�u�/gT��lT�ww)r擧��c�w��]^*H�2xts�e�"��&���l�`�d����y�����y6z�F}r�� "RPeJB������_a~i=�_��?��1�t�"`�)�~?v�W½���\�g�*�5C6���ϳ�>Ywmg�U�_��Z�g<��l��S"Q3]�Y�Օ1\���҄����n�3Q�R��VkGe�l���R��({ե��3w�P(���)��~�GU�h=�����f�Dn/�n+�9vô��E�Di���V���z�K4+�#���e�;CK��Ǐ�gh(��yu��Ƴg���F}Gj1dKYZ�͟``'�n���ǯ}�\�� ������T\n�!��%��%��{��P&��գt,��Y��鿧�Uȑ�Z������f�N&�a��<�\;�f���ch9��ؑ���
��is�î�O��Ʒ��4<�7���ETn�]�[������F�����u}'޾B��Y	@dJ�WV~��w*��1��>9a��=�ڗt���w�~�i�w�@0�ϑ�P�C⑴� �I�O3�gaȐ�/���-���ڈ��^���\�<�����{�L�fI�(V�:��c�N�TC���*Mu]5z��"�Z�<_�U|f�갱���Uh3�m�^e�n���r��;�Қݒӄ�2�1�st�������K�B��g`��XD���K� ����B���;�.f���t����(kΆ"���v�5�3\\�j��k��ñh���Z!, D�kk5BX�m�.T�k{0�Ɖ�\Ks���ݥ����g�Kt]M�v%V�
ٴn�&RfŃ�5tlvU��:��5+J�-]�`����e�]IX�Ed 0�l�0�ds�kMf�``��ųT���p�7gIj�`�7g��Й[����J�m,2��gMYm��Pc�*��b��HmdΛZS�	бД�}��30A�}�ͼ̞KF�>����t���[�͋i���V;�����U�=1�]�j7��Y�;�w��MG_�խk�����JZW{p���09������O<�N��u�����=ҽQ��Ǟt4��8Tj1\�I�i�Q^ ۴�D�%:��^�k�޷P�.�z(��BV���Z���D����Y��0�^vP�"��W� S�.;y1<}?{*D|��w�	T���-MF��'�Q]A�Q��Mz��`L"~3L��·6�(|��~��^7>ÉC�O�C�L�ww+3uc�E�(�~��
4�1Vt�C�>�h'��)9��A�ۯ'M��V�Do��)P$��ߋ<B?J�(��ʿl��jD�ʆ)�Ukʬ]�-(���"'id�w�W�N��Rؒ��'Uޠ�@���O�6��y\3�8��E��e�"&�P�U�(#�m��Ǝ{hf�i����0j�������<{Y�QMBk�!�d�?Q�(�Few�ȫ�"3��Ir��~�'8(%Y���\Z���Ϋ��iUm/}9�|�}�[1�ز�s���3П�N�H�PY�DVU!mG��kv�lxe��4��=�]�2A_�]7��t���mwwX�)�_)y��.�Y;Ǻ�Mvs޹}[s��uȇ7���}��oq�V ީ��>���M�דT��*�}���N&�rcn��.�F]�)~�>��wd,��Ξ�:��?p\F5cq�{��gv�k4��D
?b��F��lQ#��������/7�/nA�/|!��ձ��*	�A��@�ޟ]>��E��ځ{�,��n�K	Q��*�-�gs7��uY2|��,ۮ^D˲�n�9��ј��U�_L��H�">�GI~���`�~ձo�_vo�z�C��w��
�T�p�|ɀ&���=�u��3P�]
�/n�ۙ��ϻ�C�__]LW���Y,^���!�C�]k�o�ʙ�6_�浟��N&?ڟ.}a�k���x@L��6�!f�#q.����&k�A�:�D����:5.ʹVR�J'��`M��7�k��H�_)D��CZ�!�d�6��e��z�m=Y'!��Va�G�}�������3ђ�[Q(�֗��c���Ȳ�~G�U���@<t�(��|�/o}Q�>�at#eP�7��US���s.\�{��*�`e��G�7>Iʡ�M�}��2�!d�`Gu[�����}��ϓ�,�B�y��O��7�D�G��g]M�7B�+�@�r�fT��ڷZ����R���{�fXD�lD��`���RE/R�+a�F|*Y�Z��W_���Kn������+�CZu��/;浔%9@��a�-X�G�"p
�1�<o�}��V�
*"���r��:�}k$*R�K�}i�gH�(,�T��ܳ�ۜ���G���fS�M\���'ݽq(��%(.eIBgwv�n��H"X��9̷N~�W=�+�ϼ�����Wg�a�<E'��$����3��
S�W4��3_�۔Q���E*eU��ӣq�;\�[.�����0�L���v�(jSUœ
fWv�{EPUS�)����?	ڨL��.���.���釪�cs
/�s����w99�G��L�?z��}\^Уy+�5�5�[,����)�����~��B�����E�^.4����dl�4jx�MR���]���tmZ��L�݅@Q~�6'_rŚW�#���k�Qb�v����T[o�&�������};��{�����*�,����t����������y0��'�	��Վ	��i�v��F{ �w�a�SM���+r�e2�,���~�`�{���E�z�WƩ�ސ\�O�%疟,��c�E{7ڻl����r���x�k����ј�����,�Vŏn�KoGP��l�8;6�,e�����l+�ս|���z����V��s��M9w�n��D��`w���~�^L��v'����eHQ֒cr̟i����i7��γ��4|%]K��&\µw],�8�V$���+�@�8�c�.B]).��A��6d�m�K��C3jWQ���]Juգ��l��a�����^ƶh��:��&+�\�I��y-DO��D�(�;�������,)�;Xό���[��ج��]y������*z�P��Zj��jE��}�#�.�QbT_F�&Dz+�:�pe�@5�^��Pxp����S�]�K�������<;$s�Z�n*�&8�
}S�39�7�.t�@�'�FeI�JQ�̩H3۽�^��x}����TT���fx�Ļ�گ�5f�`�Sy�����]n�;�1J�ΥXk�G�-��
+����W��}��	��ߕ�:������Z���	e��i��!�|��*��?Ug`x�~�׃唏�S�a�ٗ_7��+.�D;6�-f��?�����?pÙ��� 	�w����|�ϯw��1����<�4���N �ݚ51���]��Zj2�C���G����������L��F���Ӭ�s�]�vୃ%fYYV�À]�E˄���L��f�����"����J��OW.�W=�\G{R��3X�zdI+fTI�	D��{ky��Rl�91��ծ�,��C\�y���Rjb+f���3����ڕu���M`�i���^���U�I,(YqcVۈ�&�eˮ�e��]6
��ǗK���1�W[Y��]g�)�4]�[`)_Y�z���h�%m
7 �XB��0\�
�9�Ԍ~��3ɖ�u�vt&�D��J4�uK�n�鱍-ŗm�e,],��tu9u�[�3H��TZL���]wm�6�E�Ե@hk��6���G"���+��ٙ]��B�\��U��*����َ�~C���z��S5�]TrhY~��e]�X��a_�N����j��mp/��K��H��M��}�����t�ѥ��5�еg^�̎$h���$��MuZ}���?T��:\����D�_5��p;�6�������`(*� �����v"eL����΀��K'mt�'ơ��4s�ڠ��#nv�����J$WYAÙ�(������)fv���{��>KR��Pn�K�9w��{�t/Wu����V�/>�o�_�u�������]G����+��r�Fߖ��_�Gz�$t��<+-�����&f]�F)����h��,�*!�w��f�W����2��{8�{Ϣ��$lY
���َ�7O��^Ի���bt�2s���=Cg6>����'}�ޛ�=R�̗��9r�z�z�f	��l&J�f�����[aT��v�É�i��˓V+,V)K�+)m��	�����h)��Sl@�4��Ƒ�N-tE=��&)A�P$�Nb@S�������*�6"�$s�/Q�=uv���S�ʝ!��׶}"r�"!-��;�Ƹ��u����5�z��t�j��Y�F�?�p�X�!�ފV⃗m��5���˪�]���/�s׎�'q��1�x�z9��%`A�n�,�Y@nH�y�������!����:�\��o�
��E��Cx�˘����]Q�%������̈Y�}�OE�j���l�����K�+�Sܼ�0�ƺ=q���m����f�glˉ눐�#w��|�j;=5(h�*� �-��]mV��ۭq����_@��#� �-3�'z���l����.�ҝwOt|E粟�ھ���ȉNT��x�x��F/�rGG���+��|=�f�e8���
YH�*y�J�0���_��P�'M9^y���3�<�!H��LwlkT;���=9*Jc�CƼ{Yή_}�؉%uq(����:����u�h1��SS$��$���ZD"UP��HHP���w:�9�5��\��<�."�}�\��Zk�l�Q�2)}ޮ�a��S�����n#�h� 3��/\�c�b�͹��a�) X0"T�b%&^L�G�jy���/]U����w<����r}Jk4���//���d=��uuЫ��F~�w��K�3����!�����3���@̑�"%)�[M/FD��	�����芴9y/[�;}�����#�89k7�cw	��u����%���ْ�V_I-nWZy���h<%�-��gU�oD�jM�-��57^>�*�b]+��j��"�ĩ(fś�өY��G�����=G9�@�)�ut��S�~[�3�M���3���}�/z�'��m$u6�8F��Y���h��*d@W���@ַ]�0�o,w�-62�޾wq���'VD.��;�E�ls={a'�B��Ʌ�h���m��ۃ�Mi�%�{@�(�J#j>�]ŭ��a�2m���Šh�$��]X����V!���1l����x ˄I�q����ˏjԙue�ɂ��z�Y�:�X
u��)K)��wa���GkF��y�AzH���ڗ�xR���c෹�]��C�^�O���Vo^��ЫN_��&��e)�P6�_RB�T����K,��U�03��o k�X-""���6���e��h�S{�k)_̨���[�:�n�V�"�&���p��F&�?jS`�2���/�Ҁ��6�Sƭ;�i��x����9��|E��g2R�aK���$�h�z���s5ց�:�1l:یc�E�-�*Y��C�e��W����\F:�J��h%�,��u�*K7X�Q�I-YH�y1<�9jk��6�e3��I�ݤhV�3ޱlԩm��c/UH���Uݺ;��)�u�,�����{�Y�Y����S}x��9��6�����Asy��f�]͑l�ӫ.Aɸ��%
K�خ�5�\�ӣ�o�}$tN�u� �ˬ��~сq4�Ǻ�,���<�����s�<@Gֻ���u�����;�?��DO�ݒa�L�Yۅw�'
qC��{���#a��o++O����+:\;������蝗!��j1Ji����4���{�zlYF��R�O�#;Aȉ���*�{㫞���}�kO�f�S�}MGW��^�]O���[�$n�滷�����Y{`����g��Q����Y=�U����Fqu��}D��@�L�2�Q6s)n��6�
f�kq�Jo��ѭ��]`�K�Z���e��[�_kI��5��������3����k���yl���=c�z������r�!��S��b�����P��/H��g�H��Z�b1540��Z�FȢǪrr������� �$.I���
�P//0U���R�[��&}`K�W�wZ|*���n�|��Ϸ�a�4����[�Q�	�9*�	}r��3�;(EǊ�	@�&5�}�^���<D�WX]&j8�d���K=�/�짻����1�z���v��Qw�z������-��ŘS�����W7����-�q_�*`�7��t��s�7�qe|v�l{��F�U��Ѫ�G+Y�A�ѝn�6���W�Vd��m�ӕ�iB�V��$xn������ȟWxI�����qe��+�$�$M�bȦ�3W��.�\�f���;�E��v�����	�W���f�w8F��lF����StE�e�@��=�)����H��<fL������Vѽ��^�U�α5�����8_5���rs��Ʀ��B�Ũ��x�P1���nf�~FV~������䂫ƕ��?F)zHW~m��u,��7�>#�7�����9gY�Wf�.�����FU{�Y��F_�8�L �H�k��4�WW�.܌�ľ?��oA~����}�'ΦUn��A�@��ʸ�d���Gۯ��c�u��]�\�o�s�A����}Q@��1�;�ȕ�ۯot�^���b�y�Nvg-����I9n�^��/ss;t��[����A�h����0	;}Sm��~���?b��}����J���P�8�J)�{'���qq��v�^׭��]?=�LL�O���G�銇Q�[ދ���/��ؾ�d��v"\������~���wm��A������ƻq�ۿ�D�Vk���SQ ���/�tڹ�䈎ns�� ��U蚸��{�ׅ�LL�ض�'DL�ƴZ��=����7!���}o%&�cV֓�er>�G�sF�a���^�Y�+�w�w�����X�B��C��j�˔�)��pI(��� ��A?TԶ������k`���Z��n�"65	]5��K�ͮ%�R�t\�J���S]l�gB�$��kB���������ۃ����ĳu�la��}�n�f{ZT:�]���mM4���m�;�������U��1	��V���������i���rD�d�X��X�s�u�--�ce���ݛd��&��-K�zj]�;QLB�J��a]1Y��u���LC@0��F�jL�ꕨ�fB�A�*d�C��Ys��א�,���[�5���v��,*y�u�+.:�R��r�n{�t�öz-<U�}=��D��@��]�~q���D��m<oّl�٭�~//ݚ�7S5:�v�b���m�PM�g�F56}=�wL划��4�����^�X͝�u:��u���o�9��	�"!)"���J=w��*��u��Ǐ�|�eI��׆�:�p����+���������x΢�u��~��A��U����d'̙�yɄbT��K^��g�A�ۺ;f\A�z�4Xs�Ҷ��W_[��G�$�ϳ�E˙�J�����K�Py��7��6sZ�����۷ECښ��(#"S&T��a�t�d�����{2FM���}ٜ�o��_:����8���p{1�N锔w�n��CG�;���`��:��gU��=Cݙ��o�0h���Huc�gM��Lݥ4�ź�nՔ*�0D6�B5`Ԯ�s�l�q8F"H���C�r�\j�s5\���jGg>�^���q��ԙxE�p}V��A��zS���Ct���A���eZ���;Mǡ�!^RU�ɕ&J�S"`J�R�s�n|i��x�eϾ�a�|譳�e}��:g�[��9{� 2�,�6WL�yEi���z-)C񇅎��M�W�T����U`N&6}�B���+���.^�-���7T4��qo�+��H�7�w�&�֏����)�9��a�nṽ�ʷ����0q�����@Ê��V9�	�fe�زa�"r' e�����˟(�lD�Ş��TJ��ųf� ����Uu��;�DF�ρ�BP�$�$S��&,�#&mAlL.�q;��\�fx?xh��l{�޴{���bm���T#��6��>f�~���9�y7�F�b�zX��]㡸zY�_/6`���-��k,<���']:VV�����!����=P�k�њj�,�T���{Lސ�	�Ѝ����]��X���.c�d'Z�3h�6��]z�4V]s�R��JJn������	lR�jj�T˭����JK�_*\O�y��]E�к���Zg؈��ׯ	us��~�`��B�S(�)�k�ߤ5�\W���ڈ(I8H_������X��kX\��S�B뜐�ݞ�����O�|�ř"f%,�s�CNB���Nuon��}��eNBX�����{߹��������y���ͨ��^΋�~_����x�l������p���9լ�����ųc>t�\�!PmY��Na�>"*d���Yfnu�ט��6�
�d�X�fQ��� =��ײ����S��n�*�����8f���Ip8��Η�����
B��ʕ10���{G+j�7�G�/]A��OR��
���bʵ�����oy�K6Gʮ���M��a~�0w��Lh��5�yb�&_��������v6�}R���`�'ٽ뮴�ѳ����=T	�dn��'ʕ�p�ڸʌ����N��]�P�$.�(�s��Y`Y�x�>�K���pF��g�&�2����Q,BĖY[SK��Է=���Msmˡ����:��B"��[U�6�%!�z�¯O��j#�T����3	�)�3�f\yC���~|��F[=�o��!O;Z���W�3�D���)k�a�[�cgK�w�&���]��ڶ�4����3ܮ|��4Cȅ�t�}��䛉�c���f���5��>�罐v "�+�F�nh���6�n o@�ST�}�J�ifۙ!%�|��nh�Ӱ6&�̓�tee�}}�᥽�F��6�����?m����?1���s"f!ȕ����wIw���:�;>��7|���y���N�Lj�]��c v�AW����� �Ң����7ݓ0V��& �"�����
�^��QR��ߖu���Ki%��m(tu��|���"k�8���Ѩ�u���M�o�|�Wߩ*�`�[�O��Ӻ��Hz��5�]�q쟰��ojEexVe�q���3�}��ZK�d]Kh�l��|�{.."H��+z��=r�U^�ݫ�5�(� �?~Rξ��&�	a ���@u�80�L�&�Z�u��\˨g6����k��w���S��Y1����N�K8;�^Zχ{����C� �v�NMwt��i��m(�VZ|��q�׵�I�O�-�EA�i��;�h��~��_tA� ��Q�a7k�\��k��W���w��u����0����L}}��wu3�|��5*3�����cp�X�#����"�S�dKu+C�f�9�=J�&��k�ߚ)I��t��ʋ�}���|��7[m`�°6�Fw������n|�A�Q�SϧZ��EG�m�8�� �'�;Ƣ�Q>X��E���G���Dsf7f��R���#����E!qq�c�U#�\^���d3���`��2��Ҥ f%Vku�.� ��5��p}3�(��슬U�U�p\��m.�*
אn�\����]Zo���y �\�6Q]��+��U恱D��o�ۥSo�j��T�KqJ�������=K^���!���l+����y:ދ+�sPʁ`�*/'@̄���-���Ϯ�Vkt�*��XKW\2ʱ
R��a����<��
,ض՚1�B��%q0V��qud`����y�}w]B���3F��Unڹ�4s�����h�^L�au���\Y��v���gE-�k^�K �G�3e��w]h[^Bم�7-�"�ˤ�Yf��������ǌ�kGu[k�	��5�F�[Ɩ�6�1)K�ȥ��-Ռs���s6&ƻu*��l��`�(bR[S���h���KB��QV����K }犞t�)�s�Y�=(r��N�s�Rfy����׿i����5Ԣ�L�8���س��x䦵���|�R0bQ�*DĤ�����7+���R��_(��.M?�Do��Ʋ��������2��}��N׹�q~"8�.��&�q/w�#���zNfᘕ��H��J���5�آ'�}�=p��i�]ۋ��p���'�uqG*�����޺Y��^��E�Z쳇�,�M�����"!��%,V�gH�DU�,��7����}��rd�v�+އ���-/z}��I�?}��:��z�����DdU��o�=�s��q�û�u��p������}�	|�<~�̝�L��gI1s���V�>����g��ܭch�ͣu,���Pċ���,v
ңA0�ܢJ�M��J��t�X�K4�q���an�nm[�i�J�v�����ª&�U��� �}����j�B��^��tj�j%Q
���Qqv]M)�����z6�����N�)�~ݓ\
Q5�ڸ�j��8GO,�pP����������?m���01N�u:�����HzZ]���g40Bfct��ܵ�B֞�_u��s��K��
\�_N]�9��[-�/Xs�o=�8Y+�ޕŮ�S_Q��>�~�~S��dz�}j�ʰW�{��QО�-o���T�o�`�޳|��[����������R���}�_w�3w��أ��LC��U@P�r�6{˶��L���v[K|��[�>p(�ȗ-mW�]��H�������5Tt���������˳	��#è��z ��i��G{�[
��Ⱅ��ǈ��]X'���W��0�ysa���]Ӗ3+�8#��Q6"YRa"Tɕ	%wX�
���̇�f��˼0V$�$Ҽ���g�N}��S�T�*���A��x�Ǜ���|g�[�u�F���}���|�O�?X3Q\ˣ��c�5&��iE��&ɮ�lK�]ɮ-\��s֟�=6V�`]�d����w&Ko}�=���UU)�㷫#uMdW��>E��{��fb$�R�nr^�����0�G�Rʪ������V�,�|�ﰗ����}�o���0FxD�['e�VE��y"�#T.���w�SWu[��@껾#,�{�n���1���� �	�)R��w����W_;�;ǫ7;!f���j��t@���&�׮H}�rR���Y`��������.�y���8�om;�+{��f�y�4��)]�.�^򫥷�[���s�H�x����.k��.��K�b��7��e�IϾ���ލⲕ
�����s��a?�4�eJ@��:(�/N�)M��;ܯuW��Z!�%z���������ze������]3�ܹ/2�j,��\/�BQ���������i���ڼ>껳�.�7����&|�i���'m�Md�����B�El	r�1uޠ�v � �s�����>Eݓe�$O�'�_Ga������ߞ�]K�-�؅���M�$�5�SMD�eu��k�k��*\"ݝ]��q]Z���fs�;=J���gQ��%�#��WD#�O������uS��1����f��Dܼ~�H*��{>�c��P���NV w\��oOqp���}�7�~j�_���5��U�hT��;���MH[��4���E�ULH���z�|qc�zR��p�ޓUr1��%6�XQrN��]Ϸ~3˞��7b[O�<���L�3��L�~�#��T^vh���(�{4gW��c���� �.�H��H�2�/�'2�@�%F}��k��s��\_&�Jw�Ϝ���^�R�+��:�+v\Wq�r�WN���UD�ɃX�T������=wi��8�Z�[3M����>Cx�*$��U�O4��ƀ@��:ݨ5���t �fM���;`.��u������Ռ����.�����&��Z�|�jwt�	��,����s�ie�r��ܘ�se_�dm�.*z�7tR���3ݓQ�߻gϹ��uѺR��XYZ� �e�0�M-͖U�'h�q٣t��w'8\h��t#s�$̮�̟�z)�vw�'۾��&n:m�!C(��ܩ'�� W���+���{����ݣy���~���jIݳ~<�h߹gӱv���B���4���Ķ���x����y/{���=��iӫ��qY!jU>ޜ�2�\n�ܯ@�������-���{��v; w���L����'�&���z�`*�]�^�+�k����=���vQ�b������]xstry�7V��.���s���¬��}�g������K�\�lמ��}�����Gހr���䶮^Տ}��..��������Y������O�L�w!κ�ou��D�'w�����
*��ҁ�'��ї�N�2��N݉�EJ>��m��f�Uj�-����|'�㼦}�LVo�<��Kηy��|�sC,�����H�s7�ۑϺM�uc��������}�]�F�L�Y;}���B�y�1ga��'�\�,�W#W�����f�ڜ,�;9M�"IT�;'M�P!P(e��<�p[q8�Y-K�4`��n���Z�[ɔN!O��A�"�*��gWV�^+z',՗v�^�����gf��a�t�̱�v�=�Zu�{P5�#��j�4��뒞拎u�B�k*T�u��Vs�PIcbl��f���ݖ�����\�\��ɡ��Ȇ� }���\ι�뫶L���l֛�����z���|�)p)M�n��Lh��j�m�3&^Y���=�1KFY�f��##(1�Yc��"�R-bӳ&�Bq.��3d��1ZpW��l�+"��S�6w�7qe��7��nS�o�v@6��;n�kV�XM.���������:63��r�)궋,�闌��m��Vn$��4����nV����9�U��w�e,.�\�v���&���G[��!�:܌M���o��H���Q�,���7WViAh�g(VYXphf�c�-J��f��i2(ão���d쎍4,��*K�%˗�8H8����c+��pX�(b3/qK�2����>YW�Μ�;�e����ͧ�9P\rwb��r|dò�Gc��S�bH�V��[���y�D��h=�n�1�7;�8����.���O�.˧YBݓehȺ�R���;pk��&l&\��K�]ܳ*=��ɽ_cT6t�;&�AKl�j̳��1P"���6h"������JEX��9�-D�/���r�}#�yg�0���@�ڔ�WCQ5�[m���X�v�WB�Z�m���Z�v����u�6.��*�H�������,)���n�m�GWSm.��s�hYM.lt����[!tm%��v�;n�Q���Ƿ�r`G����C��b�뵕�~yޞ�I�1Q��
�s.nÛt���3	e���\qk��\74�&���K 9���(�8^��,�g)�u�Ya��R�ك^/;?��>��$
Ֆ[���1WI^��Fkm�����҅C2�87������4�i�ik���0Q�4a����s�ɶim�-ں.k�"�
�]��H\k�9��֘.`�ұ�r��ږR��r�)s����,*�Mu�MHK�d��iy�b@���3I��Ա��������=��	1t�  �՛4s۴ͭ��1�1�u)�����΂�;���.�Ջ��顦����C�5���T��n,�cF֬7m`Gl\;��{׬'��XA�֮��q�"�Kn�Yf�0�6
k0�hmkL[LFY��&t��XJ�
�
��+%-��*F⾺{Z���[��Z�Ier��e������ͳ]��^Qm��_��KY(UQJ�i/�ش�����\c7��Ҩ�jM�������+}�M��I�f���<[4=�m�U5��)��&1��ۭ�Ms1n�4(:^�t��y��]'��!,��5Ĳ�7XBg`���s3��e�ڍе���uOgP�9���%��]pb��5�mr����W�<oz;[`ܘ�ݎ@����8\��K٬���(��i���<Chk\kv5"�0;SF �}2��4}�n&��sU��Io`�/6f��)`�ی�h�B�!���3�}3T-�]i	WPpny�<37*eI�Ɠ����Q�Ѕk�F\�� �"����\�[�@o86�c%v��@�[�X;���<�ԗ�֔w�V�1�R�n�E*�!�s�`�bk��34�R̭v����64]qWl[t��X�,!�h�A�ҡʥGGu����V�~��x�𪯓9ma-1����F��e�u)�o5����^K	v�d����X�e�����LJ776-��T틖�Vh1,5�n�j��Z�&�+m4�t�Ŗ���[0A��ѵ5�CMtձ�ekv�]
.ݫ.tb�s��/&r�m���Ѭ�&��fnΕW���P��6��5��qa���.�`꣋KSf��A�L�z�iM�G�g\�ln�33l��MRWM��@Фn՘��8KI���uqS[�cmm�2��0�h]w ʪr��{��^K�w���f���]+y6#k�<��wR��>�����(WfG{jÝ�~,X|�����W�t������XY.<D$L�2�d�3��N/�Ȏ�L���)��<�a�U�������hOh~��ߪ����]�/��S�&�ۺ�P��5y� ;����~0X�k�������Ƶ��onlZ=��5����Uԍ��kiX�B^�F<�8�']�ɔuB^��~�I
��ǭg۽}���[��џ?��(��M��JeA0�u�<��?w{��[��^��V*N�{f��e�{Mt�1k��t�9c3��N�
T��-�܃�aje@����9],����oJ/<����.ME{#�Ӌ�fO����[�3Cb���p5����Uˈc���BC{qWM�Y��><����5����("hi\�S6��,�\%�\�͗
��k��*v�h9$����DB���0��}kF��4�k3��lI�'�*��>a��������{Nʱ��TX�����Uj�Z�Q�ī3�(�����IJ)J��ʅh�*�tzu�߾�s�����X1i��!�[�M��W�H�:uA�+/���V��JzQ��7u3E+y�r6X�j�ht|%�%	�5�l�ײ=|�6h���G�������h�0�˘U���S�^��L���9��u��-HuL��߼�k�活� �0�e-=>��6]U-����ΰ��u&\����zvM�u{�:�h�q+��띕�w�����E{�����]g�'s����wwN��s������%������\�\G���+���u鯬�g���I�(��W���0��e��L�mr�󺅶��{���ɣAz=J�I�_A�ZB��1��{(�̚�&s�U�}??���_��?v4魯���i�U����_%���0�/�'���@��pE�c�������_j��'���b�h�$)�5m۪W]��x������.��W[�����"� �;*�?J�/��N!���I{ޯ�J����Tu��5蝂f��k���Y��OH쵱�^^��{��DA�>�f��g�ϔ��{���I*IB&e0����]��weGnGq̸�N"�H�r�G]��~�J���El�q_�^-���~kW���~�n-�ʦ�ַž�+�?E�:)YHRPR��g�^|s��O|Ai�6�ﯷ���>�ʃ��zݮ�؄}>�(59v��k���ۤfe�+v��U�Tۙ��rɘ���{˰_�c7˺tE�|ܬ��G�����_g�{���ڇL'W�澑�y۱���=�����-��m4�2f�Yβz+e�J'=�祥�&��&������Ѿ�|��*�0����1{�j/++{���{�Ғ���.9pT����U��*bRQ2"�%(���f�[���Y��C�V3; ���ʝ�#�<��*�x��Λ��p����^j�S������.A��n;�Ui
QD� �"��̯1a#)siR9���b��\��r%u;D�S��C�)���M�s���bV�R��p����C�DD���:�W�pL�����H�J�}�w�o������<Ip��S)8�+*g�,ܬ]�zS�~W$vYy��mh&�/o�|�֎M���*[ۋ~��^�@���g�C�%_*���l7۩|^���o~��>7��$�B[�eHs/>�v�UX	���ݟU�$V32B;%c{��,�=��U��>�b@3k�ʲ����j8Twfhm�sMy�}�e��ޝ�%�	2�����.u)�_���C�?t�W�t^���s�&m�A���BG��EMJ�[����IU�.E�g5o���@���/?C��-=�����C��ewVb�.�j��[�H����u|j��z��/U�\�WhB�e��~@9���n�,�P�|���7BD9-;Ι��d����!j��6�G�����鵉թtH�.t(�MH�x�L85F��GwU_g��wv����{[�O����Q����(���ƚF̲������34,z�t�!Hۥ�t�.��ô���-ֶ(H�����\8GI+�{˒ۼ�HUV5��. ���.���o �)�E�1@��w��e�ಛs2��ʉ���I�#O��U(�G���/i�MnEvfaD�8RԤ9�ƭ���X��ITe9��M[S���ua5{�o�	|�����)X��!P���k�f��o���+��÷k��5�|n309��S9���p�Ӻ�^k[C�黔���z���C���f�M�p��}w�n���Y,��z������#��9��-��L���nX���N�u5����?��>��:=�a��s���5:��рs�k�w�������ֶ��>Y
�������9"�d��8���E�?o���y�~.�x�n���U��N:B
'��%6��I_,Vwm�Y�ʫ_�*$OB�R�HV���(�L�j-��+�u�ν&����'N[ؚ�m��j�.�7���7NA��0�ݮF�2o�i�x&h%L��C!�I�+���96���\Z��Ԇ��8�Ֆ��c�J��k�|K�..�-��4)c�q�i���l��FB��x�	��]�Z�e��XVg[]4ؖ�f�v�$�<�i�/l�5�8�I�92��Z�Bm�k����|{ݳo$3f�"Q.G4�O��yն[�j.�ZGT-�)#6w�8fд3n[my���]K{��%�mk7�������-��\�r���L�� k�Ǝ���
M*�jmXՅ�%�ʬX��-��km���Uӹ�suo]wF]��2���n�{�w�Ȅ�^��yWoȏ�5Ad�ǌ#N>��ڱ�Rd�tE#^�OsTB�r�;܅��~�æ�}�wǶҋ���H}��򝒦O��ޔ����772߷R~#1zB��j��d���a[�>��Xc�y"UL�6� Ӻ�5y}9P��yP��usr���j�1�i�h��lS��o��6-S^ݗ겲<�d����UE��e�e�f;�E"��"IBNY��*d��B�ܽ�y?m{�7��wϚ��k�w䲙��z_�;�U3//#G�j�k�vO�[7��>Q��q��I4`♗׃ו����K9yڒ9G����:�n��y��.�D_�;<�w}���O���c�Gy�qq�n���y�w�"�T,�	n��qS.c��LYsMu�Ζ^�U��͒[-���B
JQ�Be~�%��{3:n�Af{'�y�OY܍��v)�l�lWgjy�W�h��KƑ�=j���R�Ҧv~��B� �BB"%+�����zy�ء[���+_�ڶ���o��-�J��|�]��+ݺ�műu���:��h�M>93B��Zk|eJ�x�Y�7�]'}�.�{�Kޘ��Ϧ���g��o���Ŭ�>�/���/ye�앳��=��z� ��̅��4�WJ/2�m*��q�I~u�cf��r(٫����l=�{9���$�{5��l�	b�������OJd#�C���i�����p�,��3}RN6=}}�wӻ؂��S�3ޯ:��ȓ�&{_1��`Hʔj�6��=*���]�=W����#1S�G��� �DL�B�D�]�C�
炢:׻(T��W�g<�����A������S(K�*�rzM{�E��׺��e!/�Z�]ύ�Mo{�s�n��ף��۸]֝��%c\K����e�	����]���&Pa���	��g��37+;:�2� ʆ)�������c���e)�A���XS<y��^�P�i �ul�d�� ��ə�kϠ��'���y{L�t�U7�+E�_4^C>« үG�{�.p@���K�·���W�LTwmҎ��3�.��7�$$&L���H珑����3w��߬����	�쬟D|+��Ǜ�F>�Uܶc��Ҧ��Z�[��m�V^e쩧y��癙L��[Y���g�k��V�}����2˭�Ac�Vy��R���ΰ�t�;�zc�=�V�^�.�=VC����(��)"�6�f}>S�=/��-7t��_��9[�%��N��Z����F����^|~!c|ܠ*o=�\}��F7��=.o�l�&㕛�c���Ty�%@�Wr꩝����4ù�����ê�7J�'}�i���f�R���]�t�A�Ծ{o������w"�s,�KC\y���sojP
�MJ+-,���f��y�����V�F]�H���E�'i���1�4�0\�K|2�]4���.Ô�{=%+�I���!U��������~K�)7��g��'���t�׌T[��f)?}�z��
�R��fE뽬ݱ��[��t���C����ռ;��v��uv���^ՒiW�t/ ۰ϴd�a�|�������s�[�~{s�i�P�,����u*��mÞ�d˳��~��~�/镞������fT������t&	5�BwӴ�-hv��GDzDt�BT$�D%��|�Cq�>y�lb{0�7�{*��^v>�Ř=1��|�{�j��f%Nc�ot� �ِ��#�V�)��J��P+�.�:k��D�۬��+-��צ�ʺ84��`��f�;�{�_ޓdϺ�ME��p
S�$	��Wk�Ff+]K�j����Zk�j5�ܵ�=\��Uz�M�q����#ҁ�Ε^��뚻����˒�l��h_����a��]3�·m���cV-���]Y.��[n�,.��
�z���٦J��GX���κ���cf�N�B�ޑj�4�����"���O�cHw4ڎ��?n�W;QQ�]�@S��\>���@�GI��&%��
����2�}�~��������{��=�ʚ�ѢOx�|�?y^s�k!S{�*���w�~������g��*���Cy��n����l֞����X��S܍\�p6a��Kz��е�1Ӻ���ʑ�)^{Ӣ=n��GM//Q�k=U��ё�m��^���f��55���~�i�O�i����s��f��Wℙ%�C�2�\�#�=�xbB��}Ȭ��g��`}ўϺ���s��m�3H�@�jZ���S�`���m�c-*�+�+{3|W�um��wr��tp��Q���<�{�Y�Nx�t�<>���ydImp�o�x�����gE����y���� ��������7r��O^Ջ{'6S�C��;BU���^���a��&�]s\5ikK���d��c�d�ղ:�l�	Y��63�-�*�2m�-�Z�{��XgWKL����z�<��J	�n��a[�1�fѺ��6�`1���5�ɩ��ݭ�١���z׬v�)�biZ�n��f:h,��l��F,t+`8)�f�Kz��A�6Mٻ�Vj�������)a4,���V��ݳb��Va�f:^�KeY��d"2�t���Aί���OuȊʈ�Z������(�
+w�Ǎ=[��[6�։�
��Z�����8���N�����z�NÉ�����aeל�1�oT1���3���q��6��t[<�Y�ˉ��kC���׬Ec
X� Jzo�Մ�.u������M�!\�U�Ӆ�e7I�[�&Y�o�^Ţ���^=�}��Dc6��3��}�#4��Q�D�\�e�8A)A�g�<$"&���GZ�B�xܛ���_LՇ{�t��Y:�-ϔ�O�	��������S�'9d�X�A�A��j��)�~�wt�s���/�����i[Y�7�6����t�����~��*ݕ���ɨX�e�b,��i�6n�z7�������F���B�m@o�����5���ܛ,��xE�=��k9��L��q��z���q,��@�Rp/��3�kqj�T�VL��*����%����]y�b���[���`�z�B<��0�0��� ����KuJ]w7��َ5=��^O,]��tFLYfx��xp�2��qt�^�nddE
�#׾�{���j���E���}n����[���ra�/2]�b��4�ܪ����L�m{�K~5�l4B�U,�w�͙��{��K��U��(5��N�V���K� �E��	�n�U��%�e�5ۥtK����*v�Wd�:H���&}/�wiw��Y��kt(�F������o����u���8a�s����
8҃�������tOm���}����=Yu}Dq��(��ǽź0�-�T�ڼ�6��E�B��ڑB	S����q�ԫ�{��'��%���{7���tU�{��W�hH���.Ȟ��"uu��s�n��5�$3rd\��ڹ�(�	�yq�U�59��Ovt|�·�!�s<6(5ãI�vm�ۭ��-�K3�u_-����~2;�:���g]>�W��P��E@+3���]���s��oSV�-�4�l h��hK���G�#?JYE�|�̴�7��yk^�����e�Ֆ��z��%m{�嶾z�⼲V�0+��{�@D����W';��a��.䶧�e�p-�j�j��!��MQ���3��^jͩ\Ǡ�+soP����GG��]z'�5VQ���I=����˸��C1:bd���T8i�vr�]7����f<�FY��^s�T�󏐄*8�;]�MEr��R�jT([�C]�]�y���$G3�íRg���q3��qlڙ:;�]��Y/�i���nb��� ��L��J��.#��$�C�c[�h+�u�j.WU���*ض��E��t���B�y�.����r��6uq�Vݩ+�{[�gii����,�*j�)��V���k_U�%�K�gqc���o{6�g$,1��l�Ed�N'�Fo���N�ݗv��]W;��M�2�d���b��!�J_1V辎���=ډ]<�����]i}�e�0R�"���өB�WV?C�L�h�֍��<��w�ܽUۈ����&7�t+4]z�G�7�9��I�ZQS��`K{W_Z�YR�5�+&��n�3%��[z3u����kV�k�\�Wf�m�o�����vN�g��lۗVMԭ^9�~oqX�yu<TclZ4P��e�g�[��]}�G��
ڲ��s�]9�$�s�^o~P��x~��v�2a2�����[X��=7y�J��0��r�X��NM�P���h\�O������ǵrU���u�	����K��*	��4ӭ���c3dZ6�p��������yu��.�W�x�(s@�ͼ����T=}�
,����c�O�˼5_u7���ܗҷ���C��`�4m]'Q�v&���o��9�l�T/�oVT��i�L��-y�փž����3'D���n���4�w-��nt��I'wI#m�t����(�X�og;�0��]�RL=6����{Q�������}L_�G��ͬ�����OK���W���(��!%DD�]����l�lh�o�r�xd��� %���I
�tǺ�/��ǈj;�V�g����dQʛ��4���MDoH0$�B&TB�,�鹑N��;�F�Y�b�u(յ��+�fv��`l�{@\���5��4l�|�Z��5�Evd�ӛF��v�C�J�aB�;*�jM�3.�1�,F� Wk�:�+u��e�Ɨ�Sݬ�JI�jZR����O�yd[b�����o���L7�g�,�C�k�7��dv��k{ַ+�M���.?#��7�`�ߴi��:� -�R��]�蓑�o��?i�о/-���G��Ϩ7Q;19��V�
~n�ȁ��ۅ?w۞�5�.¡���M> ��\Ai��]to���j�y_�uƮ�H�5;�1xM��}w;���Y,qr��G]+���y]M�X�i<?R�"`�%%(t�W����u��ww���u���]���I��>�<��S�×�6~i\�*7
&#
~��n�#ھ��\��Mb�ܲqVL�(_-i��"Y�7�}\�z���:�/L�������w���f9N��:LA���D%m���<�va�zUz$TD�z߫D8��b�>�o�=���{T+&l�CY���Z�Q�g���|��K�"@�샯kg���Ѱ����r��GN�2Z�M�٪���5 ^�p���ٚK����ݫ0
,���g��N�e{6��Y+��Z��C��w]�5�
	��-ˈ�{�cæ{������f��"��%�͠������"�
�$�����k�}�P�w�������s�ђ=�,�h;�������Ʃ���LZ���~����띾�o^��_k���8�v
���d�(�����J��^��ʅ
�x���-JX1⫣��VǤ.�����:k|���T�������e�^��6dR�P�ar��ή徿�I�u���N��h��Wz��|�up���w�Wx-�y�C�����h�����t�-"��a��b�~b	fs�h�Gz��Fy6�W���8dHjz�P<����J��}�}yK�~8��L*��+/�ȹg��{��.=����x�Km�PH���3;/w�������"�DU���j�*��'N;����Y�217��.-�XRS%��,��m���bhѸ�Դ�[�[=7V6��l ���v�[�aqiA%�j�Y[��;�,�T�%+J O�m�"�5�
����Y��������� h�u��6��_���:��>�v�G�[b�}e�v�lYMM�Y�
K��pQv�23q�W0�-�KQ`ku�뛒�æ��%m�o9MĦ)�A�K�D��@������F�P�����50�]oj���7L!�\�3�t.q,�Eu�v�5�]h�����桘���u��tPJ&����u��Th�
^�^�ҫG� ���>���6��N\�����[��jSǧ�c� r��ah,ӍG�{>��v�{,}Zg����z���ʽUh�H`��
��b�.����	.aK��g�[�vvm��,]h0�_d<`
"pAOJ�u�eF8��2m6��(��v��g��#����t1:�Np۷a��˗��NJ��Ok�}%�W[��׾.�J�*e!*eJRY����:G��D�#Օ��l�ç����l������آ�w�������D��o_�g��O`V�+c^X�כȖ��rx����eB����7~h����aٞ��Y�!ЁNDΑy��˻ҦF�*<�l5~ܽ�j����Oy>���'�_�Sܫ`�A��������kˉ��f�[�;XX��٨�F�R��9V1��\r�&e�ѩH2Q�����R��o^����<��X�n��uy��N`��h-��ڼX_�1�����O�^uY{��m�ܼ9�nU�V��i��z=/V�`�0��x�i�/�6��]˯;!̢(�]���F�N�u�/�n.�k���i�����)�	�{]Vw/�6���o+±���r�OOK�Y�k�{�2�j�<��*G����;����Uz���ILv_�I(��b�}��=y1{w;j�)�a �L��9=����y����Q��'�UA�m���P�\Fl���m��*���8�\����m�M�{���%�A��6w��<��ߴ��
���I:��Y]�K��f%jn�ꃕ�f��W\���o
]힝b�߽,ޜ��B��S��1��J �#-�������ω��u�G��u�1s��C?N>znY7Y_W�v{.:.�� ������\�����n�{@�~���+J��6u����&��������*]*��5�u�\i����ܺ١ll�K�4�V�mNz"MF�#GXB�
S%�!|�ߜ������g�>�?�̽0de�ս��=Ϯri5ܺ��w����`�=�%%���;�檦�O�߻��9L^���a���4��v��h�
�\�����J��{���(#�ڜқy�y��U�ܚ�u�~��8ʮ�$@�h7������I_s/˜�����^z.��s���c��1�gr燣[w�^���*�%M��s[��v7�dۗR��Xi��<�A_=��@uJȾK7�`ۡ��Ǖ���s��^9��Ͼu�i��ᑏw=��cGu�v�"�k��JT���S0��Tz_?o����n�{7wZ�
���n�޻x�Uk{w�Bʓ���4g�y}��U���zn}�.X~�h(r@*��RZ�y�o/�M65�8�Qu��b���~��>������X�,�n �'��k5��+�������|W���D��Yeh�* �� ԶA�ᣣ6�G��3J��˕ؗR�I�fQ"�T���T�N=��O���'���1�R��3��I�v�x��bU{M��dgf���83(���Y��ݥ���' U?�ޖ�}9�,{�I���7�uZB���+��v��K}/׆�Vz=���3t�.�EKݛ�v�=�̜_x���Do��̬���D,�J" HR�P�֥�\�o��c��6�+O���U�$���5՞��m�26��s���W�;Q����Z �=�XF�͠%˘uw����S����<v�c������"/6��7�+#$}�a׸��'�\W�o޸B��$��m�C��H�䳒bw`�=�Mޕ���a��ʘ �j�]���0U�����+�[�û2M�7.���,����xf�U�Sw�{�L,$h��z�ǋNa�k���sX__P�}r��=0{��"�|]�j��dy�Φf��e����<�6硯l���D"5�� ����qٺ,�)v]l��u�ًP���hmPfَ�6i��u�k ��������G�~�v����bD�k��w���������V��p���f���{�h?��;�j�Ir�^��'΅b,��D�&����~����a��.��T�s���Fp1�����79�CR|��WR��^��OP5=�L��F@�bD$e&�{�󉔴�IQ�T��ٝ��l�o��{��}��_���:?8x5|cIe���f�M�,�ε `i-B?&���:_�=�}�G"2��w@|��y���
��ԫ&�L�W����X�nz���VJ��g�B��e�5Q����~Z��lX�*��=�W��13�t{��-�l�Q[ϴ�tYu��(�n:�34�WW�j̕WUQ�.��Ti~�Y)@Js�Wz�M@�V����?TӸ)�!�}�M��sq���qO�.5P*s�k@��@Y�u�7�E�kuEN��T�����Էݷ�Ϟ	�~kE��[W�L�dścT�9L�K�Lr���K1c���6��_,�ZAԲښ�F��P����pP����R�Z��4�P����[�+�]�{vm���,GY�.n��v�.5��iS4	u���»����>�1�i4�R7�v!��(�髨�T	r�3m�nM��XBbd�kc1l�2�m��WX���mr5X���;�bɥЍ-G�h!�i6]M��%�D4�͌ݩe&�k^�J�ZF���t[s���]�%������~���FPL������y9�����;.-p%���ՙy��z T\wC-��VW��񜺝/FL����l��j���~(P��I�㇞���
���BrUw��Of��]Y���y=����ZaߦM^'R��Ωz���[k/!aǷ;飽$��M�Ӂ���T�+1�K��|yԋǅM�=�����ewbT�5]q+7q�N�'}���[�?u���7���5�=��P��-tv9N�c"������+/�FO�vX�Ciʦ	f�_#�e����*s},�1_��V��m��:���=�Q����4"����8���p��3T^��������g���/������z���fkI�䘟��P���quYg�DN�����?<�9%��]
JZܮ�\�����*i����4Ҹ���R3ϋ3_��[���@p�����UܲP����>���Yڦ��_a�66,F�~�U������]`��.]�|�7���?e�ȀT2�+�Q�{K�����[��O+J�Ec$h���|ۛ�|���!��֬"�ʷ7edGY�:��4
��ι*N\�f⬾�l �M魍QYj8��tת�z*o�m콝��������	Y8e-�*>����K�㧫���>�7ٿ~�Q�G"�(s�]�">�����w��t֌��>�j����&&��lk�O���.Y� 6a���l���D���uP�
�6QrTy�Y����=qr{a��U��-~7U��}����zt�|�2�r�T�G�X3o������U�ͦ�2�z��I'�!�,�jC����k�/�OÍWyn�����}����6��f�w��D2��gvX[~���uU�:�g׃��留�^����j��"p��
 ��e$	p�����mK4�f�A�Z�k�J�]inSL�F�SA�]O�h R��}D�}��P<l�u��l玳y��d=��:^Ww�iѓ�|�B�V�����`=���������fekD��ՐM�=���g�����<=Oy!LГ�|]����0�辄��_�"���*PW�s.�X���ݺ!
21B�����W�����d���ˌ{��\�b��۾���tDf|E�����n3L���oi��N,�F�5�.����Aۈ�MJ� ��1n�N��hZ�r|;z�+��w��x��̫��m�����qW�᳊{ХW�U�2�,&	Rҗ}��I��}=ԥs�w���Ǵb�F��v���l�7aӛ��j��y��Ѩ�Fm��I����Ȝ�s��]1ZE��I�%	D��=>�.��_���k]6�o�B��v��
Ѩx�'WT�{�F����dD���L��'c7��ޤ���F˵�ts �����qn�xl����M���n��)cp˛m�d�5jS]��������V�S񌩘��%z3!N�$�7y������1����t�L][JIC�~�k�AP�XX���u���ߎ�^����I��B#d:=]�a����|߯>��g>oA��S�����~��վ��]ޱ��|�\��H՝��w9��c�A1�@�2x��n��}��̊_>��$6�H+^KΎu꽕�Nb�{���e<���2�͋/������;�{����S��{5�>���	cT�Q�����S��|�����E��8S���J����<q�5�`���nߢ
����Yrc�XX�w�m.�G��y�Y��n\�6�uX������	�L��傎NCDc��~a廜���`�_^<�;�V����1��϶ZJ���R��k���pdLTT��S���5��߻�g��V�U������v��y�>W�A�%�e��&(�:����(��K�Q7���;s1�}q��;bv��CM��ڳhB�RjGQ[-�x��M�M�4�kK����I �����N�~��wԲ;"����f�*�J�[۾��٦	�f���k�2ku��p��?x/�7�w�]�R�DÔ��{�vW�e\^�V�p�w�w�����|n�/}��U�W��:����c����t۞~��쪪̞��:�ϧ|�d�-q6�m��=ݛ����_�ݾܯzf:�]�a�9^�����p�U��n����đ��7S����Э��`Zsg W�������[���Ύ�݀m��Ԉ��"6���]I/�;7c¡j�T����3�Loj����[s|�׬�}��#�-N��AU���o��;���UeX��݂S8�bW_G��*ךS/g��l�����24��YW�-�������z��J"M*�uرs��bP�莙�7E�μf�;\�v�3���w���F�ݗOp��-�p�s)^V��t8��zeGf�'��ul����]�j�t�Nrbڕ>���3�QlՍ��v�A�]V����.��kk c�e�(�BWu�V�[[�T|�a�{(I�����a�,ђ��Q�K�����b����#�����Mq�[�Ʈ�1aB���d�UjK���l���-�;�z�2N_n�5Ŷ^���Ón��>SiJ����e���8��ԓ4�����f���E��T��'��娢@P/WV�%��w�����[���������k��!;� w��6�7q/#�[/�N�GW�M� /y)����s[�&I[�U�7��xd<��j�ovv��_�%Pf�lͼ˥�0l�.�-�gC(����Hk�f����QY�|sjЙ��t�ʁd�,�ȶN{�*Ʌ_��X{�|��)W��XsA�S M��Mi�+��u2��'��;OZ�ネM'oz��L<��.��J�SNgfXVޙ-�MV���é^X�Lǝ�|�5�i=�{�V��Jb�@4�Q�W3��OŁw��<�Y���r�[=��.�5��Ռm��Q�:�8k;/��{�����;��@��c��y'isgn�?nK��Ӵ�sjQQ�v0P�b�I��B����)�ͭ�w=W��Y�)�3���o}�iM����y��Н���ε��վ�v���Y��O�YeZd6���(Z�m��ݶ�������x�Gm�ڒE�t˫�����//,e��]�-���`���k	XS #���m\%�F6l��ͣnř�R�����v�uMu��6m`C���k`�%�c��=n����{hkYt�itKe��n)`��v���.����u��`������%=KdS�Թ�b��]�+J�m��lѰ�a�(��V�jb!4�]P�����ǽ��g���*�w��==��	&�p�ZBQ�%�[F�u�Pa�)��]6n��%����.T�Z%e�*�\�K��륥��Pڲ���y�,�_K����3J �gZԕ�q�iUfa`�gXG\am�Jl��*Q��J,���7���`���Z�{2�e��h�5�K)�Du��i��7[0�#�j.�(E��"SUݮ3��"Ɣ�Q��]l����!����\�iWY��Uj\D��6�W].�桮���o��z�h��0;)��`弗b��mH̚��Ĥ#������#��7�f�)�K'���1cam.����kn���v�	f�Y�ƶ�]u%-�(��I�K�6F��1����0�3}C�3�>f�[mm�55�:j�:�D����k/�Z��5c���*�p���
܈v�j��ślֲ-���>5�iF~�W�i)4ŖiFV�.�f�*s3���nvi��l���� �-�큈50b\˞k(��ls=�M1Օ�w~��OYhS��>�(�%Y�k����+�MV�e���x���_A��6�t��/��дZ�oZ�l�b�h�X�LQ-å����XW�łY���g:���%�(�Wf�pL�#���L�vigˬ=m��5�ű�MHűF��l��
B�e�uc1z�dW��J�mMa���]D4�h�Y�i4�3���fr��,���SLZ�%:�H�FSP�)���tfH�Z���{��Ɖ�]���B��aԔ�˶�f�[�G����Wx3���>���e�02�ݪ���R��j�ґ����Z���.�K�j�ƚ�&��Bl�{+*FRi��SXY�(]a�ݐ�͡�M�5q.&��+�Z�ۥ߻��M�ij�ñ�Y�\��X&B�ݙ����5-K���;Ǳ����L2��f��1.��,3�P�"0iv���V�2�m�n�0.�EX��~:���B��NE4����-�5�V]�����J����aF~�����t����KB���3&+�j�ӣEn��X�����jU��H�.���λl4&�B�!�����l3�O%��;j3lMc����6��
��0��1��לu �t0 �Y[�����F}�o����B�?""���g=>�L�Y�G{�5]d��!�U�:;���8��Is��x�6���x�aL)TLʑqbH��>��3[&��8�f�\�o���>n^p�]r���7�!inK�̫� ��6��KD�^H�|a�Vx/e��d/@e�dR	=�ۢ���
��i�)r��x{�U�S>]����>>O�eќ�m�LFb��*��_}˭������D�]b?	D�
�~������x������a.��̏(�s-�)��?�ˏ�э}Q����w��b�3�=*>��R#B0�@"�7!�ro��|ܻ�����u���kvW���}|�bv�;�z���}��S�U�3�K�Kf<�:��,؟��1"~Lzc�c��Q��˰��c�sV�� �љW[Ke�R�G\DH�Qd6}��/��K�μ���O@�(�1u��pP2���r#w�z8����i3������8��#���H���	O;�]s{�k�����A��i��_��}clo
�QeA�X�U��ݟ���+쾽�JnU�t�����Q'�gs8b��/�c1.�0��v{�
�m�;�f?�����>e�7;ȻǺ�F��>ɯ�����]��zw��x����1�"��0P-���h�X�mG��fdxz��ɪ������g���V��5�oDE��9��F�SW�'۷���fǾ)�����"����H�����{O��9�������k���o{¢�.�||ڈ�==�^>� f��m�9r� �8��{~p��w�w2�ѕ0�)"�]�p'Cmlwf`��<Uà��9��`�����9�EVZ�ݨ���wS�xPj��t=�ǃ5��?=?$OQ�9ٲnۊ�EB��]��iIa��we�F4�]�)#�it��v�m�T���9kV� ��VW�H}�h[�K�@�}�<��c�-���]�[��a��b��8R9��o݇(�p�0$�B��$����؏��S��6��k���
���֌�F�?%��x���.����q��W�q�d�C8]D�t�|P*aĦ��'$&[�[5�L����y�w�^��]BM/ힼ�^Y��y��Y����`J�x�Dt�̮�%�s%ZJ�yg��k{��6�$-�,�+9��'s��AP����2�=�	�,׫C��w��d�>gw��O�Ԍ��E�~7շ����Z�1��Y�uǧ2����V�1M������
،$J3ހ�՛��gۢ�V9qS��Qq�ô��օ��6~JA�JBJ��R{�J�͕�}��"9WcMK�m�5c��䘽;t�Q����S��|]-���������=n�׻��"��}���m�Msh�Σ.��XA�'[Q��R���j���)��Į���0)J"�������|� �Ծ�������W�������κ>�[}�|�nи�����w���!8� ��{�Ýv�;�n������b]q�u6���ӹ��f���(YX~3契�_vJ��)\T~�|>��){��75A�r��@G  ��5�-?���Z�(�����<!���:�_��xl{
���ɗ���ٺ��v���u��u���n]����˃��b!@���l�=9^�ps��Vq+$I�}i�,yz߫�!aE���T�=�0�p��E\K�k��c̤��A�KZR�U�5�k�V `<t?t.IնLćr�{��]�ݵ�_[�Ѵ���"'��ܽ�����JX�a���_����--��n�߉o���~'�|=*UtI�*N��1���>]�7�����`��幮�>��9ݵ۵���B������J���)DD���A�[��P�gb̀��.�[�6!0R�%m�W��J[43��d�nIPB�e��{r�}Yz�&��7ARwf{�D�uO��w�e_mf'J��U��5'5C�DM�޾U�S~�Y7��__f�ɽ�?�S+��0 �|s'&1�����O�}��عy�Z��t�ƎW;���ʦub���m:���ys2�<�� �06�O����r3=�K� ə�D�_+�{���_M(�5�0�*Ÿ��>�I��-�f#�1��\�\�`��z]3Z~��?F�׳*ӵ���sW��*���?i�v�-��ᗂޜ����w�S���w�Fݤ.�U��ٜv�=��·g}���xd��Ʀ�O���>�@���3r_��^�7�I�r*ժ{eWXݨi����՞�3�HU�V�C��Ԧ�:�U�	@��{����L���=,ŷw��ٛ͞��a����ԝv�L�]����q�n�N튼�]f] Z���f9�t�;�b{��)�ܵ�SV�)Hb:١@�v�k��/[kE��@�î�k�\3�R��X��[��ؚY�Q�$v�Z��.!A6��Էl$��eU�DX�
�;Gk"��|��(F,��l�7�l{v�̫�p�Z�l-C���R:(���ں܅avq������D*5[D���t,�2�M"�b�۵q��&cm���G��l�*�]�Y��A˳-�f��I��X�Z�AZ�P��LfE���D�d�lu*�I������aJ��)��9��韫ߨ���q�������
��q�R�-���;ް^a�GfV�n]��S���H������"P0����ʯUfM�xP������X�]���w(���Jј���N�"�]y��T�X���媇�ݏ1~U��v�>ϻ6K ;�n�Z毟�֚=�l)�ʺ^�~K�[������o�~��m�Q��c��b+��:��F#��T�pY��_ȩ	�8���>���FzF��&�-҅�e~s���WsO��s��-U��!��u�4��9����g�m�P����ͭ�`h QZc������z�2�޷U�=�Nv
Giz]�������d��>Y��y=8t�g_1rB��gKu�g��V18�_z�ɿ4�8��?s_xi5�ku���c6�*iv�Y{R�4F����Ό�Y�tn�����><q��o�����!�u��]��u�b�U_���`�ƙ5�$�=c�c����@��u�д�s!�=uRĎ�
�R��AX���]�k���.N��G��F��ء������Wg�׹4L�`�CVzp����3}8��y�6�zݢ��z�V;l�}�c�\�YoP����-�]���d^�y�#hf��:��n&7�f�vx�YJ��}Aɳf<�������7�_j����j�30��6��ǔ�a�U�T�y��g<.��_M{��A[J����n�X���B�\K�Q�I��8����^<��&fT2a$'=E��s��x�����Hy=���J?���l������[5�8:_ئɇ<=��>���jH�������iV�Y����AN�N}�f�a>���z:�_�7��Y�����px���Ѣp4�F:"��ٙ��E�e�N��Y�Nϭ���S��빡� �H0�Rm��gK��A��5�z��QR��ip���6�J�k��Kd���y|׽ˏmkس�2�����/�ˬ��}����}o�g�{*�p���qVO�l����º�WX���_cU��P�c�r�ល��Pb��K��IQ�ٛ5A��8�n.���{��U��<�+��q����k���I��;P�!��՝zբȭ Q��������Ի��'�z�=��י�{��%z�c0wD���������}712��ra"�rhWv��թ�feܜ��l[�8��S��$�
���%e(/n٫���Sgʽ�%�6,KV]:ʺ��˧�Ѧ�4��B��f����޻M��B���r�GTV���s~�L�T]9��}���f�[%���K�s#���|�L臨{���,fW����r3m߈��L���O-5,�oz��v!��O�W�ε�:	�O��R��[.{���߸��	����mH���{r�WO,I�?[y�o~��J�O��v��5;�̫�z�U�o�\���*�en;N�v�t.blYG]]0ĻM]I`[D@A-N��HF�X&/pf�$y�g��Y��	Qg5'���z	T�vd�3n�u���Y�Ȉt�-�a�}����}��%oÅ��T���� ���e �j+��]Ϋo�˺��'�o�p�9&��ގ�d�u������JLҒ���J��	 ʥIc���+}�r\fx{�A��p�7�	j�[��M(�/������]Rq\�Q9����Iڨӥ!g���>8%�����>�&F�ٹ)��b��G�7h
��Ӄ�f���q�sǏ`��}�|�i��^�hP�Щ�􊁳7?v�L����~冽2&h&q�/o&r۬�s$�,k��5���y��C�d���:�pT�^l��`V4���E��ZHI��}��g�!��*�;ַ�AƘe����fE�.�����_�eN8��5�b u���}jfb'^�
鉓�����#����(2�̻��K�«SycV��Ƞ�m "����]5[��ZFT���vƅ�g)v��M��AvYR�g��lTK����v����O1��l����ܵT�{@�"!VM��v ��om�sn�v�E��N��p%����Fbez��Xf.:�lp���6T�CI>�ۊ�u{*M�kP�ݬuY��&Tȕ�w^iݍ(�]�8k���h���ƪ�: qs|�L9�� �W�t�>��Sl�5HP���~�]	�v�Ig����C�O������NT_��z�j���' ���REL�m��}3X����k�Y[Vgte�ɉñ��L�UXT*��|v��+ܔ�K�{=��8��)��#	�E�{+���Ʉ�(�C*Q���Q��L2Cު��K`[�ﳬA��1�vF:�WI.�Z�q���/W��[x��YQ&kv��ʁ��I�ӻ��Ɯ�Wղ��n;s5:���i*�v3S��C���FR�ϻ&,�tkJ'�*n���-װ,l�)ۣW/�TͷVǱ5��,I	���Mh)J�X���a-)æ��]R$.���3�CfM.`��V	��l�M]C[�q��I��[c��V����s6�0E@4q������i���avpKԈ�&�w~�o_v��f녕&
ذ#�*�؍���r-���mKZf�hU�E��4���kc�o5C2�5�ʩm�d��h�ێ�T������ֺ��r�Ks����m�l�gmT���`%�s��u��
q����Tt#p?�⛿`��o�|[�kO ܞ�(u0%]3^���o�qQg>ܮ\���_Na�۞��m����-,��ҋ7�e�/j�<Z>��n"�7U�1Or*}�f�7:#������隺xo���������I��\{��>@^BH�%-�jX�Fx^�ᑓw��A$�o�'�Ky���T���w{#��=�;G�(��߼ް��usC�vi�lRE��m8�I�� �hiu6�I/�7>��W���E���扵���X���<��v�՜��f�UGu�@��L�o�(pV�~����(U�� o������3F��a˽����ڋ��Wkj�g������^֘�?(�;�sU��H�&�(��	7�cq����[5�6[��M�.��t\�az�]d��4æM%��RB�+m\�Us��Z�?��?~v�-\\���wn��V"Tp�f�,N�|b?}y�'�����d=>��ނϹ���R�K9�ZsWO�罊]�R���aJ6�'(�?utʥ�.&�4�����<�C��vu�+�8�gxWr��SQ�6�^n�:D��=����Ͼ�ܳЎ?��Qt��_	(��w�^��	F�`��gw>���x�  � ����4{˜բw�~��ɘ���a��''pF����P�����{���o���>�B��P��#)�kJ����Zv������^'���1w�*�1��]5��i���N�4�
ۋ��$b�H:���{����j��މLU,�8+j�R���3��!��?p#ob�eEI��[���2�d�y��ŋ�L�An{ݑ~�}lA^B��Y��>ܹAqa��X����|�bW.�1�d�9��V����s);h����T�0V�C	=���=���-�ϋӶ����7�Y�m���<�~z��9Raov�L{5����뱃��8��ZTV��0����g����������y�v��ܷ��n�M�sK���ɰ2�~�QWι^��r��]�_}�9���iY,#`B��N����trU�f�^�ј��w����+����"1O���X��	r��hpqō�-TGT�i>{u�*��Q��u3������﫲��4g�G��_�k
55S�����ƴ�	�O���pc�xS�+"��#K�]���[{�r�@
�4ndI#�-u���l�ne�F�� oa��1eܺܓb<��t�]��㎈��R� �n�B�]pot=kv��������v��5ֶ�w���4��H��sd�͛,��xX0JpKa[�0^������.�3i�o9�E��V�Л��E����G�š�-+ɷ���5����A�&RV�U�c7�,n����>���Gܐ���H��5.�����H3�j"��[�K���o |�k�k��%i���3���nN�E��$Q�9_�pi�q�
� n!)h�{.:��Er�k�o9k�E�I�}W�z�V�!b�U�g	;ɬ��JQ{ۛO^H��6��`&��\�8	8��l�\Z��Lk�Qq]p��hv�pB��{��u�l��j�3�S�T+\�C��q[��'{ ���y��-�s��Ş�Nϩ.��Zf(+_�U�5oO��Y�viXy�k��w5��+��ո���L���ǝ���:�ɼҍ#��u+�_L4y	�e�%�l����m1�] /�m��Mf!u%�����*���t���ջZ�����jS�w��o.m:�U�w���iU��s��+�A5�xwc�
܇?�ފ�y�[[����_	�)�'�Io�����u�h���"M�TQ��c�7��ZWǗ���{<�_vJ[�;� ��E�x/�ђ�����2�E��3(���#^��>�ރg��;�0tLML���;���]W���:��ٲ�gv�W+���˧�`YEx�+�L�b�~ܰ*�r@�&��N�b�c��KSU��u/z2x���m�����Gʕ���w�b����U+��_JҾ�K����>|¿�6��t��e�R�)5EL���!�~�+1�sfs+uLL5Zl�[�h�z =�~�j��\��)����~P����o�2�^��bϨ��O�5�{s~����f]��<<��m���l���'S��w�ڛ7�u��g�7��ծۭ�4��mOg��/2�y3ķ�񉕷t��\�oD}��e�8�x��W�J�%��E��$D��W���U�{�S�+s/��}��ν���nv��m�|}K����]k�������
�$�.��2}����3�)��Z��J1�׾���� u����w����ۼϼ9}�
�B�-�Hݴ�#�������[��i�<Fi�����f�%��L���퓣��!St�f�|^X2�a�{uK������F�r��i�O�2�D2-7�R|̙��eM�织"H��osFs���~�ʫ<>��O�<*U��W|�l���^�P���@QŐ�㶸L"Q���+(Y�BX:^���4��[%����ͮ�ے���l8�� ��=��|;�_���͠>k�np+�:X�r�v�S�g(?m�V]�}�`w��[��p���g�d#�J��p[ �uΪq9Q~���y*�U��7�����Κ5�:t��GNg��/g��υ�Z��}��hjܙ��k�J�, �����p�s����5yK-/�̾�w�����q���v+�=���|$�u��]��{'Щw��ֺOj�1zkҀYaPXJ�&��u�V�٫A�����]�6<���oE�{7(6�w�H���Cûr�oElE�4Wo|��n�]>���<	�VB�֑9On{�kuL�6�P�^y������֦a^�y���8��&u���V&�_T��/C�R;�]:#	41q�&)e��L��y�^���Z���mDn<c��������]I���u���Ua8H�!�$����t�t8���ɍ-U��֚����9�pK�v��M�i�,v�ے9�%)a��U�6�K��[jɍ6e�#�Yc͙�5��"�"P���^Qn�-��T��	������e�\h�]�t&[���{KkE��v��j�S@��?��y=�ѕ��nڬЭ������&�\�K�Yi*I�L��v����f�%ņۨԖ<�R�;k�b]-�YV����6����]�e����5�����iK�T9�.���;M�"�ec��-�\t���{w?�v�?�|��%Ut�s�2B���,�~�ՙ��^A"z������>�����j�݋H(O����^ɓ<��<��]�����K٢�m��h�����������ps]������������~��/w�^���}��U,��� /L#1�>K�o�J����[�*�]���t��^���y:��@Ǻ��D��Y���Y�<W�10௉��0�)���\�P����1[��6�5���$ѱk�D�.G:���W��[�5�W�K��Mob�O��h_�&!�	&1X��k7ҾGv��'Ie�}����U�}��=G��9�b����u���}��_ Z�y���ĭ+��k��q1��f������w�5hݍWCW]�4��%uԑ���l����u:�Dj@����s�~�۩�$�C=U<���}y۷��u��:�	�����򂌔���T����x��.C�";����d�1VYcҎb�{�t�y����gW��e�Y�m��(������'-����5۷j��r+��n�Xwt����WM�gS�i*�La�H�.��m3�o��'�mB�Yu��+jkJ]�ݗ&*�	�}uQBc��ª5��[J��}�?2AȈ �"a,ZtwX�]ڃ��u�CGq�w�/L����M��Y�5q��CcwK�/�i{�x��7��yc���g�A)�R0�����[D��+��C�=�7=Y���*�-~�u[�vO�븾��m�e_�&rlJ���2��Y���6���5AS��LD�g-Ϧ�7�c�(�x��������?���Sy�AM9�Ρ���עN���LQگV_R�\�x����-�`�ua`%N�뭁m�3c�6�B�=1�)�jMi+mԭʁ��+v\��n5���s�CWk���<��-͍�é�4MEl�kv���p|h�ϊLr&ѿwow���2m	ss��8�i(0� �%����G��;	g��0;U���3&�=�����>S���cn/E��]�����ƾ:�����<o�U𬎲�Q(�T�yGj�S-K��ꭕ���rb���jӹ����(uvw!��ܤ��ȳ�S7j�fa-�LI����9����9�wg%yg�'����+y|�p�t�@S{�S��oG���Nb��V�|���D��x����L*&5��DĖp�S2"���:c0����Ns���r���4�]��l7B�R{��w�}��y�e�鳘Y��Cޣ�lrJ�d&�$��٩����q�Mܿ�o�-:���`���*VzmN��c�W>���"{�EBH\>�弛�qo����O��B��di��m�u!��m���SgM���ԗ�&�X�cs�.�;k����N�l'���3Z���Sq6�T�	�����;H�F�_E�/o���O����= �N�*���˂�R�rbe˼��}�}�\�8�e&�d}l.����d�J�������2�y.��|ݗ���X��Q��L�t���Q���v\!�����2�������ت+L�pۍȍ�DL��{[�+'�8���I���_Qօ:I\�V��S,��׭�����2�|�k0_5�F���5�N�o��}���/q��)׏խ-K�_�Q�HxQ���׻�6�nQ��q���i���ы4�YCki�/\+	����f�5�◸i�h��=�^�����B!����d8$��0�m��6.v�=����xO�0��˩s/mf���p���Zi5���s���sw��o�z9/QO���>�\�D2J�~
��*HfR�4�T�� �F�WZi�,�5�.F˴%�K�~��p^��fy^���;�pƊo�|�vY�=����z��
Um2�:�9+�;��p������ɱW(�e	����${6*�6:�V�'�VD�!W
X����o2�KC-i�5x��\��������P��학�Qޜ�'&��\8d�^����x0�xK�97�5�x~��u��=����`�6������Lz�{[�٣2�<��|�@��ЍH���<|��s> �����/����q�S�>�O��4�
�	FZ>嫓�^B�7���.����7e�����YE�����~�����j����i��#�v�{�"�Ѕк����L��"��Xʽ���5m�|��{qf�̢e�ʹ������o$��h6)O=.f�%���R���Z��*�g%������o\4���Δ�7�\�t�� ���&:��G#�+Yh�+i-`6���G��jLR2組��ψ$�%&.�j��h:�R�9���<���w���%������Tv&�,x-a����|�\.Z���&��+4�2���/k�33�v�8M�$�KsLD6
�ɬn��5�I�b�hic�0�l [K57m��X8���3��%��V��5�6��B� fi��
�k����v��7�[�[�oGG���p���.t���G��k\w�@x���̔>���˜�n.��4��g�2��oF��q�����,/ca��1�׻|V���g�:!��d$e3a�Rs���0u��g݊�������P�{Ю���b�pޭƗ��]
!�ʍ�3�r�Z��bs:T��o�^k��[�X�%lN����Ϸ�|��n���Ѷ�i�B����ޓ�����,����^�?#���z���СH��Z>�;:iq�-�Z��ݲ��<�8����W��%O��=;�k-g�p��2��0���V�~����I���L�����03_5��˩��o��QQ������V�d�B��ط{��ڵ����U^ϧ�^ͯ��D@u�T�,���vt&)�a#r
rA�p���s�u^\娎nY@� 
M��À���w=�9x�V��Y�n����YܟE�u�boۉ�Kbs�����uz���վ�r��_�IP"IH�1*�_T|�n�����f�7��mә��y�+��ՌF����u�v9��]��;�
re<x"Z��J ��d�TN
P��s��0�B��ĺ�U+�5� vyn�3��i�mw9�Q��۪��o�C�o٩�򪢫T������r>�/�랣,�e�9>���UH�����=�n.HX0(1��ғ��ѵ�5��dBa��3g�}���7���uL�i����Z�j�=9�99 ���
�YY���@j/aL����Yf�i��ݬ�Z��Μ�Z������C����J����w�յ M;�������^�i@���L&T �Ʉ�-����4ø��(��p��e����퉱Хv[��H	uv묫Wzw�6������'�G�h����Ϸ8ynlѶ5+]�{����{@��}����UA���$�~�<�ޞ^�0�E�!yeÜ�f����&��%��Ae߀�DY��Q��Ψ����Y�ky�K�,�\^�ŷ8|�ݦ��zr�4S����(ӽ�����$��]H���{)��YC��T�s���]���A��ȅv���V�N̕��s�)���R�e�Μ��h���[�ɳ�	�Dq�l\��=U�:�ҁ�s�Ńrm빾�wQ�3����R�׺��6q)�2��9�$��3�ӇN���L��Kb 0��[���1>{���Se�:�^瀿c�[�#����$h����7���B����|~z�6㉭�@���Y���dq�al���u�l�n��-�7Q{6.���%�ӁX�>�9�=�ץ��;��ا�'.���l�^�R�ԫٝ�WOc���{5��9��z�a�� ArZ��ʆ~�����J���e娺&�p��_�jGe`��ڙ���k�&��׼2�U�mX��8Tj0���(��G�=gO�������׎����S�5;���ͷ;�iQ��ȏ�%3����Z3WN�4��O���ٷ���>yb�}@�8ܞ�u2�=�x�����]fUd�Oq�쒈ʝf�7�ӿ�K�rb�in[��,�u�֨�X��Ux<�`�c�3e��I�|�'��u���K%D�ЮP��w��}�y��g����7��m9ַ���E�Y�ns��&E�Z{���&9��v���@�ٖ�u#q7mU��Y�ز@dTj�D�j�Ҹ�H vX5'Gd�S<�(�ۘ������%�cϏ�2�n��3
�>���5�spEQ1�s��$Ovǵ�G���cn�F�?@�y�����g.����ߜ���%��Q?C�b�C�p�[x�m��R���_�������2�P�@����nٻy��|f)����C��Y�,��f�ضzB����]�(/%��ܖm{ޞ-eE�Y${�׽x��B����
��ަ�Ow����R�������^M �^d\��=_'K�l��e��{5s�9�W�&dJ?�a���e�Z_
�hHux�ZƳ�~w�|�ϫ�AOv$���T ���|�� ��(��2�c ���[�U(����*o��~eB��T ��T ��s^o���T ����/���������P
0��A+�?//��A�k���P��n���B���:ʄ=��=m�Jy��֭��ۦ���*y�T ���?�ʄ�n�����۶��q������zz�u�*x��J�w������)��������l�8(���1O�r�E)T�\�ݕvַ�� u�
y�C�Z �Ǡd�����u�����r�v�a�B] =
�{kY5@ת���I�l�U�+��{�    
          @                    �       � }�%>�AJ�m����^��ʢ��v�Q�� wM)C�*\�z=��s�"�q����� /xE�\����p
�iJMJ�^���HZ��z�wRD� ���������y�{X�{�y�z+a�/-]yt� e�=�Ť�]-��ؑ��q��q��]|�և�*=��e�     �  O��*����Pq�d�d����Τ
Q�񆄂��� � :kA��l�h^1����eA��(U=�<A�� �� <�����9�S�^1���ʪ��AE��:�RE�j����Jj�w� ���v�nc��,�C���O��)q� U�>-�UTJT�� �R*��]�H*<@h+�%u��OF���6Om4@� ���}�         m}z튧�H���7��D���Ԏ�ӈ:�B0 A*�8��0�k�=�v��A�J�^��� `�f�
2j{0QT�P �=�{p��^1��%�8 �{�OΥB������W�IQ���ֺ!x ����۶+��ɠ�M+�g��۵ky�ک[�݌��@v         �zŶ���Iw�/1�y��<����mG��
r�p �����aA�.�^ض�y�
��=����� s���rn��n����Rz4�@(��� ޚ��w�ރMV.  ��E{�==IG��=$\Y%'��x ���=�^��㷶�նE�����zw������P         ��n2s��{;��o����hB��=��om�| �=�����E�Z<^Gy�U�&�hD�pK�c� tu���oG�ůM�����yg �M����)U���@�	S�c�3S�5_o�����RQ��GҊ�g���CF�7\x x*�t�qz*�@�1ݾ�}Hy�N���1[�4
S���~�R�   O2bJR�  )�6�5T�F� =��A�*   �����@  OH5J	� ����?O���G�ү���%
kqMb�W��I�O8���'tԡs��,��P�Qԧ2�P�Q�BJD/�P�Q�$�$�"?�IBIDD�D$�DB�O��U��TeL�����J?$�al����,�V��V,G*��dT�&�pi��Gv�h䤅�î�)$@�Aѩ%ȶį��Hy)�j\ME2s�;*�$V�`���
�1E=��z����_=�U�S-�u��mۤ���٨/R�����!\�csWu�	B�[���x9����u.�J�]I4U� ���J�
A-ڀCwn�ۡb�Zv�=yM����NUB�xr�J*[����No?`�{�zj٦7�o �E��|E"��܃&P-�f[���X�V��{�Qv�kK�G(�-EM��n��Π躘��5�N��L�.��њ½�0JE�dL�h�TAX�F7$�N<˷� ;/oFT�nV�ɮ^,x��ˋ�t׻��˦�����Mu���l@��Y��v��۵Vq�tBqr'f��V���n�9�� ��ֱJ��91M�V2�<ܸ[��WF������ �L�0*�NV��[�M��˾g��l��ѥ4җV԰åw����q1��$��<�*^���-���ŏvܸ��m�1:V�6�Cp�y�K����ޖP����Q[��Q/,����#��//!"a�6D�V]m�i"�FQ��S� U�A�mj�S���%컭Cw3CQY�����coY�,�"^M�P��E��XI��Qէ�V֜/��:5�JQ�FD�	��i����B�qMh&�\��(�4"�4kvɗf,��Ixd5f|�$㒊�·Rwj��jݜk�7��C2<�g&n:�ض���r:M 4�t��U�e^3���U�$�d�ۃ54/#v)&e�����t]�Qn�qa�(�REYr��D�3v�J��	��$�;���[��:e�3����]6a��TS%5�"b�8)B��-��FiTu�I+n'�o!�ej��L4� �������{e&�[�@�M�����vX��[�j�LțB�JI��`�*��lU��KҋŸ	�aSj�'���^�������6,)e��rRv�m���s�/H�+RX(
!M�[y��lCK�֫�l��8u��*�Ҷ�>��Czb��\(ב���a�L��b�N��t���s B����A�w�+y�nS\������hm���n!����������mKYI����ײ�%d� �M�<�n�f[�e�P�+��Z�f�p; �H�^�Ķ����ސL	)�r���փS@nm:�r��������F�Zs�-�%��UxJ��{�g �� �Y�lU���ʉ��2��cq,:ej��eJ{�f !",��A�9Zbi=y+p<�� U��^
��oe����@J˶�Ge�f�ᬸ0l�Yg>қo�^���j��<�@�ɁۥE2���.�Dݴ��Hz��ӻ"��3
y+"��7
9Sc�2Ŭv�t��������c\�f��w�B��=�Le��7^!)b�y����P�ͨ�Le��e�rp�K�q�e��/�܍�v�4W"���V�
bU�sP�MpK�s�S��o ��Ku���mB�MHc�ϙj��K*DC[Na����5�w,[��}�S1U5�ԡ�sR����y�� �Y�h����v/"��]�!�\Ԕ%a�{dVf�15S/b7�-�	��H��X���S	'Y1�{���W���y�n��m�{2�
�ohZ�*-������.J�3�\M4������&G���.�Z N^[�V���b�=�uyp���j�Y0
�vr��� �S3Ng�ړ�Z5���:����Q<��.�0ņ�������fM.�f,S��^n�
�r��4
w��q�"9o~Ԅ�-5�p�[�m�$ژ��,SF�h'u�ƳwE3!U��؁�j54k��_9eƚ�y��ZHPF��rGiNZ�Va�%��KmlVʦ�`*J�1��UyWDbߎ2t�
�B�׆�����cVC)���ʋ7#5�D�nN%6������t�)��LdIjV�E\E���b�Q�����n������0�ۋ]�K(Ս��k5����%�
x�y��F��)�Ϣ���R2�*Ɨ3����w]�Y�?� ÷�Ǒ��G���*��v����z��.c}lk;}�r���\��|���T�C!*7����V�9x+e���6fB-O쬽L��s���:̦��u�bY��c^;p�ڹ�,�-ަl�*S��+�c**[w̒�Wz�i�2��㭿�ѷ��'���YCe�i�®��"��N��K29sn��~ۂdz]ۗ�	zkׁ]���܂dv�7��%���DMTD ��J��pË*e��HD�N���6��n�b=�EÛ�5�kt�Ǯx!�Wm�b�:[&�i�-���#i��@�Sn�m����R��:�z����&�A��rTg]_M��o���㏥*.c���ӫ:��Q:5]�����Z�/4�f��9h�dv@AD�k����R�I� �K�gjLk^jC�,�ucq԰I�u��C�oR26�������&��B14��{r��)�i<�A�w42&<�5���B�1,r�<�7r"NF��:Ev��(^@�0��r<x�lĠ�e�a���W�qPՆ-�oe\V(U���!&��Xx�(����iգ��$�Jb*�f���l�k��:@}���׮�y�;���+r �f���;�9��.�:]�fc\c*;Z^]���r8�,Z5Y�u�@����s`�mi�X�0�ˁ�D�ڏ�u���L����3%Î��խ�j�]�jQ��H� s�E�]f�)LA��^5T�r�����0X7�Х�^*���2�s����(+�Fj*�C��r�WW,P[���u��.[�ۺ�^����B$j=SjL�w��'P�ҕ��4y������G�W�y\#�w��K�#��_��h���\�!��g��)��X�)݉u�VD'-:q
H@��"�J�$Uٝ�����$z��1�����h��������-|x��V��n����4�Î:��Go#4�O�nJ�U�<�F���������5��OF���w6��Y��)
�;Ku�����28ayW��Q��Yd�E8�����9m�N]^�	BIH �$�)ޘّ�mh���v	ң 讵�e�*_>�<��*�-��xB��Z�F�'����Q���nT��&���N�II�K�j:*���pkH�*�s4�q»��A�v}�7i�oU'��if����:k*�Dm���j���a�b���)���)2i?1}�s�4m{�ڕ��
dZJ�d�hQ#�Ӟ����ɂ��%�=%)%����9	�b"U̴��3�OW���邜w���3ׯ�.�[�/yI�|niM���ZI �N�b,Y���ʒ�F��yj���sT����W�֪lD��y��� HKB�"�&�i�ز�5w���c�9u�&l�Maͬ�glP��Nm��Z[��Ч�O���\�pD)kT�ar�)X�ܚi>n��1vEAC&R�br�752�����b�:��-3PQ{�u�&�q����Dɪm3X�D�hhu�H[��y(<׷�(��n�2�T*Ś
2�!U��#�=	��o$Ƿ4)[\�6K%�ɒx�\fnUP�U�P�5�\�P�l�Y�J��չ���[EbV���ӗ�^�1ښV�Lj�Ī�x��>�kY����-N`�/�ͶI�J�B�nVV]�t��� �Fϴ
�*��ȩ�-%%�%��j�1{�z��5�/>K�^c��o(Ŷh0�'y�$;��
�%b5u팡�T-H��y.�[��F��L�ǗL�؞m$MIt�~��c.����66�E�	Zԭ�Jb�3�0;���-ߚ�����j��6���5��������e�Xr�J�E�AXr�H��c�D7u�B=Y~X�&��M�J����]9�D�	��gN�Bl��k����zۭ����f��Ξ�h'dR�9�\e�b���˵ot�-�8��ְ�ܔ���aʰ9d��Y_/2:��8ոj8v��Z1d6�r^�'aOv�*͉f�G1S�-b�Ҭ��*���%`D5�qL�cX��yZ$��6�-�۷��޶o��ii�hTrI�����D��ӧD�.$�M�Y�v��ˇ����Y`׌�LөڗA�	S-�x+n���ej$�� ��Rk�7�����1�p�P@��H�.���L�F�W�m`ERf�&�͌]��U�k���� ѵ1Z�Z�ek�cnӦFIji�*�ۤ�*�D��V�ͬJ�l�d����0�(6ܕ��8Ea�Z�h�� �Q��ɲa�(��J���雥��2ܴ�2vl���b�tE�Q�4]̪���ըoA75ZQ['(^	ta9���U!���Ghɓ-r�Ê��ja�m��*��O
�뚴��3\�HI��'+1��h�D�V�^V*R�_%�Ų�X9t�j����g��.�x�NXж��{����e�bY�ښ�؜ �y�R@%�^;(�}q"�l�u���Rt�Aу
Վ�܆ecܐh���I�Zji���IZ/i8F�z��n�o��G
��UG˥e�J�������׽�商���Y[e:\�H�-h�Ό���;�@�X-��m;��Fμ;t�麼w�k�jb���jͧ��F�be�Z��McK�t��	GNP�4bn�֜о;y�d�iշ���x�W���5�Fm�������.����eJE0�ɢ������,�}�XƉK���	D_�8p��FA����a�h�ݥ��lbXT^S�
����S7cS	�vm�LKH]�r���:(lR�S�LJ�P����D<y�s�i�m���U3�3Rɗ�s�֊���(��Cb����EN���1��8Ҵ�v�$D�$����p�ء"�j���{�T�9��So/1���.�@��h^��w��`Z�a]�Ϋ�st	�H����&�n��!m��T�Mȵ�!�&T�E�5{)��"��͙nac����;�b�q�y�iw-ӎj,�r�]���[y�XT�l*��tM��!��In�:�[Xn]�+l֌ӗH�w���܁AM-�srS:��m�ñ��-:�[��N[��bT�*����ۄ�m;X���-��VFԛ��J�&0�!�Mf�L�2����,�Z-d֨Ż�6�-"��XC*Q�ʒLY�J�̔��7&�*�5�9����ͭ��b6~�2���,6��oa��{�9��9hf�e*�Ʀ���P%\Wn���e^��r�\�v��#'{sG�12������Ŵ��fōl���֠�ȕ��P
���+%f��h:��dx�����֫;�.��D���<:��YT���:�`��|��xڑfM�����zr7ɔ2��Iz���ۙ�hAȒ�Ga��R��"adŒ��Z��V۳���ͺ����J��y�Y2]�[��%4-�AOMśu-<�@�L|�;�����
�d'�p�Q�B�����6�%����wSrV��]hтV]��4�
�g�ͽ@){8�"噆{���G׆���Оb�Pn�NśZ܊�6�[2�JJ.�'��-�ݱ��?fLj�f�����3jo;qF"m{k�?q��� ��{Aw#�{Pk���s2]��Ad�eIY6���l�(UY�F^�T�v ��AL6Dp���ֹ4�!g8㪻�kk);jMw�̪ý%�)�l4�n�&����5bdk>�8�v̡A����|��բ�S��2Xq�Z���n.+%��	�+a(� мxn�KB+3�7�ӕ�y"�=��O���w�!Kt48��׽WV��v5j�CN��b���*v*�v�/�Vm��]2�1-�M�wr�Z�!t�!T��bKN�.#�+!s�>��bq
��]s$�G�ӹ�-��]���o4�^[�����kKobp:����A�OT���LcoX���K&o��9��<�����+��4�#�E�p����Ԃk�)gn�2�m��.W�K��|=�B��
�^�B��k�mr�E1��}������~���DoV���Z@N<X�:$�d�Ƹ`�M�\w�k�1,�{�ݎ�
���^n�&q����n+��
��,YSo	q)z�'.NG��+��+z�
�oB�.�Z����L+�i��A]���:��:E�2�V����v��˶b���FZT�(��ڪ����Rp�ne�F�lSl7N�	ԤuX�{x,
�kf���3@�P\�6��v��l'zi1K@Ìô>ܳ��z2ޱE]л�3i	*ls�v�՗C��T��2��Y6�/F�P]�j����{h@ʳs7�E=Ų=Ph�`�m�Im�(e��<�Ov�d�k�/>X�s;8D�հ�����4lA4('m�	����I˴*���V�*�/S�TJu��YMc�fŭ�Z�ʚ��,F2��󆻼8��v\1����8�G#N8���L���d��I0�Ŏ����҆b�}�(���k5s�����t��~�6����Yz���b���V�۫��'L�L����3�"��ҽ޾:� ��>N�����C�s��i�8�Z6��1G�{�NU�w���o�)���* ^^�ŵ���P(��.f^`L
%�n�i�R��Ĳ-���{�D<U�FS2H���y����*�̒��_�F����__.pnCvG�]�^�7gY0e;�H�T��)��.wG��o62�0^ܽ�r���[p26b̊��QD3*�.��#�xNy_�Ń�����
BYK[���2�����nx'�Q�����#d�3+n�"U㻼��ͭV�c���Y&�2n�&;7v��akV�����Q�ΓY-}���'N�K9�S�aȻ�*�M�P��\���F�j�M�]9t �[H�8   �R�J��U@�UR����!�ݱ�R�Se%��v  *]�@` (1�ƹ0~|�}�M��iVVV�-RT�ҭU*ʦ�Ya啬�[�K�]��SR��UUUT����T� �mUUP/-�@UUJ�U+l��-�3+�@��M�� �����w�s���÷�����-��k'i����w�w����t�t��C��Y�tv�8ml����2����Km�v���m�`��;v�<;�pnc�nȶ:��"�=�R cn�^��(�I�v�궮�W�ۮ�;l< Wni��w�:�k���kvwZ���u�h�.���a���n�]�i�u�.��m�����d::�6�ܽ�e�|0Ͷ��w���'AV^���p�(���a٢�P��[�,�wc�d�<]�b�;u�M�zz�#ӽ�4#n�㰶�t�.�����n����n�2%"�pu������n݉L��w-��tv���i�ٲ�"=����Nr��2��B�)9=�y�x��}�
��<���x
�H�8j�E;��SN�Qv��˄��X�"�9N��)많�Z�:#�w��sq�lAq�<gW�z��{N���������\c3�D���>�7�}qg+��ۑ��3ۗ�*n�H��b#�ǌ�c&$��u��n���;q�m�UM]�����с����N���,9�'b�*�6�+�� �M����t��uݣG�\�;\b^�5>�Aݤ8:j��p�d�\r��z.9����S��Z��0�ˋ�+v�h4`3�\gv���̛{Bt~�]��I��A�F:v]�Ó��6��S���+�_���%��m�^|��''[X;\�����^�5��������w��u��7��]���n�4�ꃨH��;ds��S���[nhcS����5c��c�p<I��Y����<��F�/F�n��۝�npt���$ܝl�"�a�tZ��R8���f��k���=��wd=��
�'V{4�&�v*�{zL�ܽ�^��a�T�j6�s��9w03��@*X(a������,�
,V��w.�[��������g��j�j7	�x�m��s�q����;r�.Ľc�-ۋ��Ёc;��Żv�<�Ks�o.����ٹ--͇�����^���&�;u�,�!
��X��]l�If0�i�u��\���n�zۥ��v��瑻<Rn��㉱�5�y�`���=���C�s�M���u������&y�ף*ݞ-��Pݢצ�q�r$I]����c�X���pv�[����S�v��y�nɧ���)����=�a��	�y;u勭�v����pR��f��aM��Ӈ�N�/J���đ��v2�
hy�%s˶X'�eyx�'g�p܎�{-T���轇�C\h+\m9g7F{F5Ʃ^�:�u��cÍܸ��}e���Jnf�G��Ӯwm��:8]r���lF�!���axi�;v���u��d�Ds��U�e����5t��q�yؼA���Rې��lgom0��3����8�1���I�/�=�V��:%�g/Non�.'e�w��=�q����.-�۸\z{<O���8��m��}��p��^�=hֵ�w}n�v�Ӱ�������c��&�L6�}q��r�^�:����h.&��:�����Yݺ�k����i4���iM�=�v���N���J�R�d��:'�Vt�s�u�۸1Ϟ�UA�c��4[XzoR����Sgkm	�T�tq�b-C��m��6��|q�/{vN2=�tby���������zAD�8:����:6G�n���7#b�6L���G��N'�l��+�����^@�@gn��.���f��,f�������hj��v��j�n�v�ϓ��B�@T��U�Aܛ���n���A�zd�Iح�ݪw�[��]g >��΃v�n���'ۄ۪�}]n�0�W=^+��}�_}l��S��z9n�^.���L3z�[�m۷V�Z#\�:�\a훆�kV��{62NGc�Q�فF�g˵tvC�8'd}�jzF������:Z��/;���d��Xy����}m��cF�nm��F#]�<蘰d&"�#h�LLh#��cw��93��Mn��g��7,�o(R'6(�.��T닠ζ�n�v��(=�q��Wi�����GW9�ł]=�rt)��x���n�@$��a;������-���9���c�vs�y穑�h;��@�x����;� fȇ�H��ͳ�fuof�sb�.=���V�tI�;tp+gչv�8Ru7j��q� ��ˋ�l
gduk[{�g�m���6���ș��"�<����0sn5��v�w���v$C�����Z�;hnRYv�6,c>M6��G�8�'k$s��Ov�^�q¦Z��&S����[7S�GF�Î��c��,��xޑ����c]�!��GK�ɶ����C@m��P�KV��7'm�[�8��xk�	r��V{=%��z���xu�ۣ��s�ϴ���A��v���<syI[�8��������[v=�NK��bp��=s�d���u˷;�v�v��ټ�q�ė����ٮޮ��f4�u��G^���#��"����n|z��8���U�v9�1�K&�jݕ����vn�8��f!��Xةb�V��~ݶ���pV֘�=��ǆW'key�� �/h���֋c��ǪM�m���j{s���e�Ē����}Ԧ�=T�<9�q6�d�vv��]�ڸS\𬛑�\�zNxN��M�VݻZ�� �cy��c�F����}p�M�vǶ�^����m<�-��ݻ|w��Wҽb� {8
z7���=��O%�i-�o`���D���]�Wm�¾v9����U��iw�!���n�#uֲ�:<��ѻm�㍡���]��ާ�>������ͻϟ>��q�q�9��.���z�όg'�sF�I�l����h�2�n�q��"y�v盱
<8ܛ�*�ָT�l�ϷY}���[%uͱv�Y�N$â��A�];����VΫ�uv���=�6דnL
rtX{s��[��H��tk��,�����=�O�gE�c��K��rfNCn�M�׷�jM%��{Z���9��	��vཬXvNw��,{�{+<�&�ls�iK�;%�z7\�Ohqٞ;�j:�x���g����sw<�޹z��vu���z�f�};�l���H�oT��<��z����V��%+nN8G*���\��,=��tgWb8�]��Em�/�9�r���d�f����\��]n3&��΍�e�V�{��	i`�kӸ����:�2V9̛���^mצ���W=�>�.��r���Y������/F�GG'S��p�`^�I��$k���0���fn3��w��Ŏɸ��a��;
��=��r�`�mm�m�)�N��뚃�8�r��[.p�t�;��§e�˻)��v�oFی^�&��n���Q��m��\�KӸ���u����۬�d2��s��IOX;���gɞ�1����[v��tŶ��@��t��ӫ���;;�&��Ǔ�q���kz�m��*d��]"u����!&��o@�������I��oR��rg��ۤ']����F]{��<��u=�+v2r�g�Q����3츌�U�v�pxŪ�ۭ���y���5nf���۬��{aε�v}|ј.I���/;s����V�]�Ql9M��0�s'��#Ά����v�6J�g�ݪ�x��D��v��;��;Lm�iǭLb.���㭕�qɃ�p۷l퇤�xd����<�;�q��c�[�6W<ѭ�n��.i�ӛ'f�{p������l<�ܧ'n�7;�ι��r�r�yG��읞��\F��m�T;�η[oN�g�>�˭�n
�s緥�q����x��n��~��)�`48���>I("<u��;��Wc�Gl�}����>�ͣd�ڝʵ��=O�4IĎ3�b��Ί�6�u��.����[�1�O6��Eg66�������m״�^F8Gq����J��C��Ş�Kָz=�8�n7O]v)^L<uzș^���>�9��H�/2��H�zt0�����<@A�(���gy�J�����x�d�k�/4]pmnƷ')Z�Thݝ�\��R�\��]�;��=n���tD�}N��^����n::@���A�,��C2m�ѻv�ͷv�]+ϸH��h��u�v�� \G\Ok�v��S��ǵ���]���k�r���s����W���q89]��n����&�v����d���-���<�k��$9��i��^K����*�����/1뇺����:�����0S�������)����f9�f�F�<����s����Hm�a�d��nr�8�k�u��ܡѷ�ۉҰ��v�83S;�{Cc�c��ky���	v�b����#�
�������`ۍٸ ��:oU���;�}�@��CU�6���1���S�vr�q��pI�]u�7m��Z���P��:��j���m�i:<THi�4�ݱs;����<l���z����k�Ä�z�<;�vCps�
�e��g+�v�[Qlr9�5 nz|��m뮺�l�<��u͝�v���ck;=�ru�џ4�;^��Z�z5/��Lm�mm�.�n�s�n�v��홛n�j۲�]�;s�^�������X鳸:���U��U�� ���WY��b�]��{Wc�"s���Hc���ێ�\��Ԟ:t���u�ԊK����ud���v�7K�p�:��jy�7mZh+�{�����P�]����=�n��O�R�a��g\h@��Ĝ)n���F��v2b��s�˻S�{F�&��u�&�79�v���{FVľ����RlWX�mͷk	1p�1�n��:���E���z�u�6��w��y�q��m�Mm�G�Lk\��v�=���X�Ϟ}�y��;y���M��9�L��+��5�����.w�[۪�c�H4p�Ƹ��f�6S���R��!%	%�d$�$�"?k��%
#���$�D@�C��J�O%T�:*R^U,�\���ZR&	�\�+U[:��V��F�m�8}!�A��z��{��Ɗ���KZ;���lsvq���뇮�H�<�g<rk��W��	��I['.iF�ڧ���휶�{k�Լov�S��Ygۀ;oBs�g����q��q��+�۶ݝ��y۷I��u��\�x�7)q���o:��ܘ�Ӷ��$��,q����K
v�n#:玴�:.\r��a�c��8:ln�'��Zcs���)�u�v}��sӬD�z�L,i3\�K���|rhx�R�d�������{a�u��y�tnv�5��mƻ��ۀN`l[�ݍ�sթe�g�j�KC���z�rudW<��8�Ĕ�92 ����;�(@�	�u�sݞ�5v��2s�=B��O�;NpF6��c�̍V�y�9�1Y��X�3�������h�Gh;nݴ��.ún��]�vu����b7�͕6�4a��a���+�x��:.+�=�^su�n:6���mfՂ'�ٶ7�e�;�,�¼u���Gv���ٷ��7iD�^�����٪�.R��gv������X��Ǯ��x\sFɞxGz��3�0�tr[nS���f����=]v27%��)��-(�=\�ַi������\9}�s{uS�b�mp�F��&Pݑ�H} �$� �a�t��F|���&Vυtbl��ý�gה�H�^t�ORl��Yw�ym��ήk�z���ڳǇ��8�]�vc�pA�\�[]� Q�w/������Gv�X���p�Ǚ_a��"6�[���Oml��<b���7\���;,�kl�`�{��!�a9(p�T�vSt3���z+n璹��^W;I���u(�n��=��'n1���9��S�g�ۏ.�u��R�K�s<t=Gu�mۗNu�=�����'���m�[[;�����J�7��蝮��;{���,:wY�}��`�7`9I��uѶ ��d�n{96K!�u���y�w����@�0�P�B�Q�dB�	$�~������Vgej��	Ojmu��;��Y5�����v�F��aF�&��Gd�x�����b�,S���z�q%�ܩ�퍌���v���y���6ss����;c��g��ԝa-���흽�X�<��c�睰m��Kw=��O�ت�����Sۛ{-�9qW��ݮ�H!�V�8�C]x�@]9�6Ηcc�����z��@�\�Tt��{˜n���;����܈�/���d��˹DS��vM�SJ��D���?�aqJ���f��t*֘�͜/s*�����
���H��Ѣ�!^��`�%p�R|�?�m�T�K��"2��ݒ��)�v�7꯰�ˈ�X�����wB��N�{�{{��G�������4jD�r6�1�3��{Ȫ�-����%N��7��]��D�z<UI�ޝʷ�;5R��:<�`���.D����NAx�'��,/����o�3�E=��$y�`F<|T̫l,\G��v�V�[I�zQu,��Ӎ��Q}#J=�U�b�)Xv{0*]�J��v2�C����h��F�%���*|���9n���fŎ�s��Q����G]L���<�mUx݇���q]�˺�z�l=�>�re�zID�nO}<c��U�Ul+�Wm�(ҧ~���w\���G�M�wfm�>��d�	��-a\��O���{��	[�e�}E�g��u0��#�[���޵���;YS�aVEmJ8/pe��u����6����<T�dX�f�vK=�5ݠ�v���n{�ڼ��}���C��U�8���V͐�g;�/۾�\k�rs
7Ĩ�1YA���XL�:ǽ����x�Qs�XH`���P玭�삱��##��e�&����N(=l)bZED�6�SλS4�11����],�^��링���$��&g�e�J;T{�ԴSZi#/�.v�V����fZT�T��Th�FKOo�oL�^q���]V���j؇�;��n�N�l�_{��XJ���zYE�ѿ�L]e�H���*����2J7��kc�*v��f���{l6����=;���G&ۑH�rv�+�C+�z����o:�l�Z��.��*Z ����Jݻ��^I��'���G��ps�[.4�1�2A*����{�fft=)%(C�8� �M��R�ұ%ލ���-z�Q��'��A�s��i�h�c	H=~��y7_�i�ΫӲy�.T�<���{�*���2���i��NX ��m�85l�Z�ɛFx2{a��n\j��'��p/R���&��K|����˻|��.]C�;Hw�-p8�f/�a�#-���p�ڮ���e��C϶�F���G:X�W:�������t�m+�=�/7j�&ie�}r�n�1���k͐I�@�NI=�a!g^��t:�;Ֆ�a�b��b?im�y�V�/���}��������}��i"|�������v��㹪�O�@C/�X�����'9^�����(�]����{^t��zMD�h$�6S�m�+��b��5�$�*�(��w����؋���/n.7tF�,J�<�B4���%��N7`E�c�]��M�9]G�Z��ޖ��=V�V����V٥t����du��T�x�;z��D��w�(�
�����7ݯsf����A�x���\�"��y�Λc(�������1�|�b��	�I
����'$��r�W���K��)��V�����w��_e�!8���s�&��_X����Y�$�X1��f[�墨B��U�M�;�gt1����T�P]��+hޯB�O�5VË,��ܢ���Xj��r{g����V
|�1�$d����򨰃��S�*Rf�h�ib�ٕ�� �!��{�ռ��Lɰi�FbF�ӝ��̂4��t�M�56y��;9���\ud�z3\۶:#]���Y�ӵ�ۗ��7Qî\7`����9���� ��^y��o��}�M������U��Uv;�mS��&����J܇Wz��DD�\�.D�)cgM)G�x�u��2�܅��D����떓����#r�Au��i�bt=5�ܹ�oy�ǃ<��P�!.!	$��r#u�X���m�K�ymkS1g���2������Il������1�~�v.�(m�X�H����Ѻeze��a��!e>+Π� �HQ8�t��@��q<�a�V,M��]��؆�z��O��Ɛ�831ݩm���֨�Q~���B�Ae�Ԡ�J����ޔ��^\���}m�Pov����/	2��]��k8Ҭ���� �[�桡�^jZ�;mVZ^e�6�1�t)&�du���n����ٖ>m�������J�[���عN���	�on/6%q��^у<F\��u��n��H<=W��k�����S]uZ�Dy�>\����`4ur;r��դ��Ͷx�����݇��d��qWn�(��9C���{`�oX���"N5�Ӟs�O���lUrv�t�c��ds�Y�P�]�pvn��\nק<���k[�1�������c�s�c�n;-(aa���9.3s��iۤ�F箺�0��[#q-q�����[Gvk�#�I�k����8�i��w��E<����&d�ۻ��u�3�6u����s[��q�j�sB�������o�+dr�-����yR��JGkh�t��{�7�ت;�tu�ž���j�����ӏ\1��)�:8O{M�����r8�$�^�V���mz�����w?�G[��YyEZ$��C�.��$?s��[p秷�W�O�c�%$9eH2��L���]�N�1��i�X�����4��U٫=��V��t�um�f�#TM�TJ#�8���cnI�G�*�q����s=�!��\T�j�A5�չ���Ľ��b�<���3vQZ���*��g�x���ee��И$m1�^qu��N{F���P�����brmË=��
q7a�%>j�NN��I�z����d��}��ZF5~��WeD��5OZ�Sj0`�W���{+aW�v���Mt%3$�'�
H*�G5���wx�JE�҂�Gg`U�����Rн*vEy'S*f�dTB9m�7�on�K�\�yq��=��]��FۛR�w����ۊ�,d붬X��z<��7��{�MT���̞Sz��Ϊ�<\��Ňg7�9� ��q�#A)*�S}ڎW�gz���`�P��+΃��p���PP���VXV�?A�҇{��B][�>9JEB9���ܹ��R��u���yo=����=Wk��[�D�Ρ��4�7mo�8��ݽ���e�"�篥����a}�)��I&X�cF�3�?��&��EZ��)�$�UrP�p����3���g��S�&���sՔ~����hAc-�ްZ�޷T�^psr�YVn��{fn���ݛ��o6h���jVKF5QU`	�Uy�q�1d��사B�I���bH*��{&Qbs��r���2Wf�e�A7��MA�E
	�G��O��}����;x%Ϗ_��j���/�N�D�"){���\��=�.�N�8S��Ӵ8O�ƣ
��ڍ�.��[���K���#,g>;U�G4�<4�x�z*yk�%�Aژ{V�������1ov�6�w.�O/�X)kb��Bz2Ъ�g{�S��w�7]��K{s{:9\
��p�����R2z3j׷%��W�z
�n�HTbۓ�gA%w/@�B���O�e�L���v�َ�د�tN���IhI>���8��gol�J�_�y���m����	H��w�%���C��q<�_�U�C���B�u���W���9�����^���G�6+���ɓ�a�hJ��lj���y4<�m��]��۰tW�w���p��qe"��f��&�]uA�{�}��)�;f���U���~?,_es������n�<��ľ�H��#��p�Y�]h��_��xr<x��DͱkWH���#��pz���KT��_�������P�ʁ2ى)$�2�=�ӧ�Y]�MX���RJ���c�,�\bN9��
���U�7]�i���0@�*$ہ���=3`+�)!w7����jw!�=4���L���;ƂL�6R�=B���^��T�N�-��o^+�٦M��oVL����{�Pjx+��o��x�f��щG��$��CrF���e�-��C��`���F��`��"$(LJB�jb��ƴ[��z(fO@�8�VD�Q�F�U��u�^��^�V$�w�c�ev+"�3�U��k�m�n;�����H��=j���p>^x�'���.����n�Mrׅ���q�$ R�͊.byUy��-�$��<r��e2�m���;�P�5��{ǹբg�N���Η����~6V�i��e�ܚZ(��\R0���~Yp�pϽ�qp��Rn�e�RЕ�=���4���`��T7ږ��W�vs�-&�\@�Z%�`�����W�~ru��~	ה/&}9��fgJ�麑��\\�C]cԱ��Q��{i���L��e�,�t�9DN�͝�c��c`k+��V��	A�ِ$x{�6�R����N�W^G6�<苄 ��	�@o�Y�&�]�s<�+,xn�}Ɏ鞪{�q�O.u��������`;�T�b�(�'�o^{�PΟY���Օ�w���܍��+7�6��g^o�n��l*����֭�xqRM�ʕ�ܽ���W��\3o�����d��j]u�j�ͣD,��6�S��{/\�n�ql�����.>;B��i"�����������%�p�CKϕ���kz��n�n	�O4�jr�8�����倁���)9��]�{�tX lF��m;"=��λN2��黭�`��v\�T�zq��m�����pvg\� �n����l��]&vy���`g3bA�-�]����n>�4�u���s��m͊�%�.v�n�I��d�L1�;��=��
[�?������+7��j�P#;iN��"���P�ߵo�QW׍	B�^�Ƕ��/��̀��͠˼r�:����Ӡ��n���CK\�pm�ޫ����z�c�l������.��P�-�fϖ��TG�����\rS�f!Č��d;Kɳ�y`m-��J:x�U�*�U�lp�%���5��]������4A�EF�nIpt�A��B��N(�oЙ.`�a���7ɘ]J'��,�QF^�M���ڽد	.,�U��N�6�`�h��KG!���j��q��=���6s���j�S��<Iv*�$I�k������=x��ճ�$�_e�ݶ�v��'/Z�sp�r7.)86ζ�-����v�-[�D����k������dw�.K� ����5�L��]UQ����wӥ,�i`9�������2�:K��;u�z`�&�)C$+0W��4[kk�`R_.������>o�6�d��(��kskl˖B���ے��P�mZ�)�ֽ��{�4v0?�͍��Wr��{,y���{z=�(ά��9ΤH˙�{k��b6�������IT��r��q�$�
��Қd�_uO8�z�Gio��PӄVj�iKԡ���nwxo�ݟ^Cr�)��8͙��C���D��,�xigbǛ��9�����xU J?W����L�[-�7��#1�REoo�I	���ݨ�x�Da��VH�_�#1�P���ߡ��l�(��@��3�:�u|�/H;pO͙;ǫ;sA�J���֮������G~��_H��ai,�X�D�Ykqn�N]8��gNԸ�K�k*,[\:֒�;k��H���|�4}�^N��Ļ�K6�V��I�p���;�.�q��x˄�����;j%��OL2�r$ԑ�$"W��X��U)�h3��43=`�{L��u^1�mz�����+�C��4ѹ.����@�nБ�&b��z�݂��Do��]7P	_{>
cL�ܯ��t��c�Zԑ#v4@z�Wa���v�i��: ░�/kR�÷;b�n���G�L��+:�=U����	%��f�%����IIU��K��U��w<�@���B'kuډL���\~;�}��f��m�'|ȿz<&��ճ�`'��B'�s�����K6��/�1�fW�-p&����7���*ޜ3O3s{e��G5�c��u����ʄ��F�d%�ux+C�K���Wא:�NV��2�9���mv�^�Os�n�8g,`��]0�J�ؘV^�Ȧ�����MZ�Q���'JpQd���I꾒��ˬ���4��ޝȂ�{]W9��KB��mEx�d��K)��U�ߦY�2ɧ[i�ṯ��]պ"���jJ��wd ��J�.��F�n\ƭA�*a��F
<m3}��:��`���q��WA��K/@�^���:�b���{N�W���=ݢˠϦ�MM���S�J��ᴾ9�'�Ef���"L_*�ۭ��ɕb&T�ĬM L���T�����֤�3j?*T+&��z�Q���d�{���4�_'�FI�i����	�\f�N�>�vw
Is������9@�;4ݚ��?c0?xyh}�u/#eQ�I-M���݋)m_`���.g� �1��j���V٨�=�B��Qm's`��H�*�V�{���1�q�J`���V1j-�EP�o�c9|�����:��6�C���i&hg7,��]�m�(����{�[�B;�m0
�,�����E����}�tS `�)jgw&"Nfgp��)G�ت���y�X8qQh��L����qX[�;�[)��N�"v�V�sg&��ٞ�}:�O6�rc���kzA���UdE��h�H��� ����yb��x���Yܠz�П�Rmy	��E/+L��.l���`��fS&�u�}ֺ���Z��	�g�ut��ґ�5v����۴���&�	wuu׆IQT��Tr[8fTt��r߹�e�fOK�7J��C�1���ؼ"�d[�5�I���Tad��|M��c�Cw�3�(Dj2K1��5$fw������kV�`��axx����W�yℊ$wΫ׌��m�|�Ul�T��ιZ�ߗ�Z���_�ڶr'%�u���ͭ��l��:��b��Q�Fx�텷j��yG6tU���H\�;�t.j��$�!"��/�^�C����W��O�� �מ~��Gۻ�T��8��t�d��=oL���,qx��Flr���'9�<��Ő�,�P|�?=ڡ��I��f�n2=�,M��Xڙ�J��0R\Z�¯o��el�s~�%
���D�N�(B��R�n�]��xjͽ�sv��$C�~X���d�r50�&�L����)r�U�Z�*�!魨�����fU�I%aTT쮎(Pew���7%˶�X��Y���G;VĦ�Hɴ�sq�g\'�"�V�'�n?BF�K�˂{
��kyl;�K��k���y՜jgR�wCoU�y��mK�*(��a
M�A��c�j�y��N�;���^q�<��k6�if�5�0�^��mp�4~�ɛd||gQ)T�����873����!����'���E�Ӫ�j-�4O�����=���۬��kp���=}Tq��VB�! q�=��!j7�6ܙ���]��o�m.=}kQ)Jkr����ƃϱX��F�@��X0��wJw8բ���ә}�,]�C#��"dG����У�)��}�6������9uۺ7�6^�{���$�)[r{r�֮��Vu���W3���x�P�YW��9;Y�G�Z���u��T�����w.ef��[�͊�s�b�zP��spQ?qe��M������/5�;u�efr��� ��UeJ��7l�<���ۤ����Kﻦ� ts�l��ήRȐm�qG��L�����N���v̻d�Y�K���P�m'!W�[�D{``�]�"��ûX������ttё���62L���t����V��lf@��؎x��v����9�#��ðe8n���s�]"U7�6��Ǝ^K�:�F�=���mnΗ�Az
� +v�*Gc�k�-xX��ξ'�}m��E���Y?�˾';��Y�ј�d0��ۢ`�P-(�ϥ��H�7�S2�V]�3�]�z��]��ܠV���nU�QS�^<�A��PZsX�_�S�ly5ކ`�3���ݣ�$iVhE�����Y�kK�zi��<��!
@��2IP1�ݫ����w��no^6���������3�y��X��mvC���J���@�@mV[[�����_s2ֵ���%���^�alu�c��da�nجt�I6��4�ڼf��nظ��>��=��M�L�q}�~�BT4e�������!�cǃN|{(b��{;Q�����6-�Ku�i�]�u����8���)y���F�sC'�bݳ��l�#`a�Ftl��ۛ��盙yc�q��6���OVnޫ �ʉw������(��rT����^�pL�e����?u��R��]u1����I���S'l��&�9$�a�rG~-.�\K�u;������_W�ʄ� ��[�F�F�hnL�N,uwL���]����|f��ԍv|ˇ4�9�)�c1Ц���ɜ;�aI��{�4�����`-�5��捽��-�s�Ƨ�����Z��E[���J��crI��KF�[b]t=�3���O5��j��mw�Z��ʕ��'e��]=�ܧZ�����O���u�(y���#�Y�O�:"��u�um)��_D�T�5�Ӿ�;�7���|�^<�&N��%����,�|(1X$�@�����`�>��}w�᫨�Y�h�E���F(����E�#|�׵r�v���Ŵ��.d�1K]'\��e#WK�n�`:�p�e�Y�n�˘N��[\����F
0�i�u���Z8��b���Y�rE��=�m�O�](V��Q�^�;��"�un��zQ��f��`�H␢ɑB�r,�1��$�ln��]�#���݃��t�Y�{��ot".83)��8����sP\��Y0�T�C�}y�`^��)�)��xͿ�;��/vu�ҽ��c��ܫ�SHZ���aԟ֌Й��kzT��M[�t/�-����|�D��]�~(��Y��ց�7 n��pG}/e5H@^�;��옂晦�e{�����oJ�^���״2�>pFM��n��̲�e>�X���f����U��0��e5��c��Z��k�[�wP�iǲǗ���k^��E�9�]u�}���ڠ�Kn�
�T���}w��RZRv��R�����_A�;�n�1��]��Gn���m7z���f�z���֫��5#
���o� �j���]��x�c�'%�T��7��F������e�����t�a
3]�����[ J���J|^k��[s��sr�X�`5���q��"&�)�I4���Ї�k}��}*��@T�v�q��ӥ������f�K��e�*��2Y,�m�{�$�V0�����5 ��ٯ5�����i*�ň��}���h�Y�i�5o��y�P�}�*巓^gUP�ͼb�����	���nv�����X�j�Q%���3�Y�����������kJw�+ݻ+y��_fY���)�0B�e�:�_���l��g3�+ٴ���O8���l�����eτ�/N)�0#����nt�㺲qr��ټ�ݮeL������blQ���e��,�C����*��z(���N|��;7�F���&M'���^_����˾l_�>��5�י���'H�#T�L�n�k{8�s�v.ڴG7i��Pͥ.��qS�[sT��&Bʧ�Q�_O�����wAT�@n�a[�$����W#�2�u{��f��}��:(PV8��
�nRٻ���h7F�4r�*�0�khn�������;e��mL�,���</!��U�����E,ʦۦs��,�q5��n�Ϥ����m����$Z���ffHod^GTUNB�3��^t��گ7���(��d��[��	�޸I�8�k��o�F�$�����=��Z���5{ӂ��6j#�)נ�99�'\3�&0Hp�D) �c��_^��.?C}cw��A�(vlʺlM����s�/=�9�: ��U���)'�(��0�^�+�n7=�X����+�%�J��h�|F���,b�t�im�Of��h��\�Yj�˼
��3f
����fZ�x����Gd�ջ4݅�c=W&Jv,n��n;<r�/nx�������&۶����e5a�i��r�����6�O}����絭�&e�rE��N[��:q�U�t.�T�m��;C��3��e6ޓ�3^[����4�qv:�&,[���^�%׀�u�(�$x�Wϱw]��ݜ�V��q���sKn���`�WK�I�۷bM�+�p�Nf+$�7[��kqk����Ϸ*�
�vP���p�[j��W8�iN��YB�N�P�y9 [�M��D�9���g����1Z��Zޤw85�;�g� Z+��O�h���܎�,~�&5ސϯ��֥xSf��!wڪ<�^8jȿn�=�.K��jj{\>�~VEm(�^va�
�gV��{)ĄL��d{%R��ٝ�-
�-Qs��vG<�������z\z�����ee\��u��)�������ב�i�$"ۍ��/�����ݭ�V��Gfu�ݛ��w�U�1͠ﺦf�l��WD��l4f�e����̩		�����FP�41Kj�����D�����n�^�L�b;7T� ���G�Y̼���h���6���y,�]CMXw-Z| �~����v���zP�S6�tb��u*���{k�j7]��힞6�`۝��L&�m�t��YK}�/{�j�w�n�7�Z#ѪG��mg� T���3�����/=w�Wy*6Ůș�D�iə��U
E�l�_�,e`�w��+ٌ��,32�Rj�
��"S�Ҹ-��MW=ƞL����\�(0��!B6�m;� `���YDaN5;o��c�v��;o����^W�2%
�8�:��-
�k���`�f��դ�E@�q�#�����F���(c>k{��J硎�d\��j���� u[���������Ъ�ⅎʍ⌞���3��:{��N��B�[۶v\��K˞��)#�� �:`�:��W^�y�N//M%�����hE��[?s���f]�p��J���]�=�����s	��kz�Y��U�����.o���akU�w��w�|�{
6��E�R8~�� ܭ��t]�tum�"�k�����6����+v{p�Z�$��W%�fT�m;���D񫱖�%jmt;��גU쨜oRu/g9�kO���d��u�I[27�a.���=����*�Ūr�:Ӫ�_N�ɶ�^3�-�5_H׎�J�P��e-MS�o^�ۢ�0�4"����$$#�O�6{zK����I�Ys��U�_i�o�Ү1�S�ɣ�+Mі%f��^��N��Nq̹f��'B��PA��xcT�X�W��ڕ���ޡ���R�r�A�^����sh�!)�i�Cq4Zd�$���h����Z��Q��k&�_�7�@��1?]6���,S��zׅHy�t`a��˒Hn����Xݕ#,��H0�m�d��p�7��΍X�S��˃�K�{ W��m�V
8A��<s���\^�z��e$�r8�@H�Q���,��+��vU���Cv�:��|�\�I��g.�#,�	�)�Bn�fy׹�ڨ]u
�z `G��ݽU�E�v�'���ܟT}�~N���N��C�e�M�2����IJ8"�ʾ�t���d��s��w�~����4X�]�3�!��O��_;�2^FoX���6v�f��rٿ('F�'S T���N5����w6{�sH�QwU��n5�A�J�k��l�xs�x�V��T"�/-��$�2�q�"���R�n��V�H����.������#{]8��̼��:�j�)�
�_v46.u_`x�gx�.��֠�{�G��B�ۮ��0B��n��은p�[�O�^��3r�\�M�D7����yg���<�;ޞ�-̿�������C����Kn�A�B�
��+�{��gK��Y%�lJ;uy�㛝z8(V���<f��������l �&H1WU�%hQ�b�؍qչ�磕��W<`.+ۭ;��"֩�N�["��3�7�[�쮊��.�%P׷��{�h����4�A��.l�#j�n��f��,�QD��*ʅ0�i��rKB(�i�۲���<�v�����U>ٽ	�ȼ�)�ɝ��b�� �����r��i��C�Z*:��R�n��gz�G���*��ޯe�l�q;��)4���W*������~�#Ed��H�d��w=V��B�t%�q�.K"�?.�������t�J������Cf��F
��f���Z.������t覽6)��Σ�=adO>ߪ���²KbRr���ٟ���w���/�(��<�ٽ��QϪq_��\��}!]��+"�`0���`�-!#D���_����!ۄĬ���եG��
K!z�aP�����o�k/�r��ZB�)
H�Q�i?{t�ZBd���H_}��_FF���洨ൊ�V5���gS>S:���_������t�K�p�&�P
���(�y��n��(>��~2�٥E@{��Z�Y�X8�XY��0���X
w��۩���T�� � �HIFK?]ehrޡ(����3�n֎��_��[�XÜ�ނ�t��I�no0ws��5���ϻ�ݭ7*��c�A���	�VG0%�ilY��G�%�w��[N�@.{�C��oxw�ۜ�����s^�Z��Ӏ�K0��4�0�le���k�ft	��`$�y�~�MJ�!�ֶse���sYg�#�wPIc��(��QےK�y=H�k3�R ��­��xr̡�9wk�b����N���"Ezqi�齲k��
��w�:�+j�W,<PVkx��7u��ܯ�C�t'�;^��3kw�+8nj崅+Zyۓ5�c���G��'N�z���K����(��!����o7�T�xT������}W���Q�&���-����7gI��U��[�b&[ʸ]��+j��ZvO^1�'���FBb0��y5�K�QT$��ם��cf��-�������^f���;����<��ҝn`Ցjoq\���ə��dGhA\���3ws��h��R���[�\���!�pJ�s_9\��)R\��v�5�t��ɱ0�ɂb|��ǵ�̮��,�M�60���e���S��װ3����&3������R��uZے�ǻ�r�mG��嘁���["崩Ŕ4P�N�K)���B�4>�͙���ݹ�/L/�fP8P-�̍HJ�Sݣ����n,�)1S��+��lj�F	�bђLᒔ�m��X���u�c�6݃��{D]�o�rXk]��\���^���v�v��m�����m�N�BeKX��'~
G���)*7��gLM�n�[�y^j����-���GA�ݶ�۹�7��8;Mf�gu\�����ݻ_F��|x������#nsob�'����^���@��M����nx�L��ZT�2���/j��N�iI������]g��Eѝ��s۳��5;�ۭ۱�m����ݽ���`-d;[������u�-�ǎۀ�M���o6ۯ�>8�w�Gb;&sД�;��r*���l���	:��_ecr]8p�d{q��J�.zm��=g�ӷg���t��^ĝZ2��7�{��h�{�8��G����<��zȝp�v9r�`:v�<k�/i�eŹ�+vzg�ּj��{mݰ8������;v�������8��f�ll���nx����'3�lۆۂܛZ�v��;��=xl�6�5<�`�Mouy;��}����7g�׻���=�r]<`�`�W���K�F���Rs�vv�����ݸ�l�����n�m�r��ŻݞwoOq����0]���vf<��֭�1n�0� �(s�fv:���Ƕ����wn����`�n�9靻�-{q��)6�m6m���.�ܮ*\�u��w���ݾ�!�j��}RX�ˏnz��snƳ��*u�t��g�ݹ��ˋE��=q=�y�Sp�s\��]�onr�ཀྵ^��.�O�EpCf�Ӷnɺ�]����m^��ЎH:��v7�k �
k�N�-�ֻ\�y���&�Hg� ���ȈjS�2�	N�E&
s�iX{c
Lq�R�p�W�N���gG�\t�V�<c��˷�۵`�n܂h�Ӷ^]n]�6�pu�n�n�pB��n8|t;��l:#�&�.܂���Y�V��j�n`��NwhE��g��
�^%�>�Z�� 놉+=rlup&rl�������Bd-[0��z�9g]�A�P�������r�m)�%�CWa�E��=;F�K�˝�[W��ʫvO-��q��SzgU�[�c۱��A�U�#z��+O\1ϛc��幞 ����^:�=�!�]�.M�^3z]iN��mv�ڹ7V�m��h�V�p�Nm�ì+�E�x�ų��������֬�;Z�t��G^y{m�����m�\s�>J�#[�nڻ\Z�9��/6帰��R�̎�ú��������\-��J�Gअ%�lՖ���j����n��(�/���_Kz�͕uܼn�٧�[�X�]�����Z�����J��!�L�L�>)u��n�ja�US���$�d����m*��U_���4 SG����/4�Ƈ�5�`��(�۸*�8�9�6|5�<pX$�!�k�ʸ��B��H?]��\��H��ͧY��w�yU��?�S��"�4ܽx��;`��5%-Qp�Z��fLg���ԉ�{��L���YX�ucI�/+qW[>��-d�ϳ����9�2���V��}U�&����Wm,',��]�LpJ�D	��do{H�0P��Zr
�Y���?5(���»��xO?5����(�s]
�^�7�4.o}�+!v��W�9p�/i�y�Z���STP�%���W[�~�A0;�U���2>�C��QY �;�%~<$O�-'�	ָ�#�������<F�b�?gt�0�n(bS3)i�|8�\|�Iq}��x�ܟ
?�I�~��{'~��7��!Q�p�r��.�^�z�=ָB�p�dCF�����W!�U��~�!��o[�뗝����ʶ���Ccq\��1�<.��) p��Z����[��M���5dxVV\���E8�ܮ+I�+ߔذTA��P�>����.q�@����E��% �m\���J��j�ǧ��I�*e��z/;��՟\�Y�����;��������t�YV���<)mT�TD�#�A�y}��@�%+��"�IJ�u`ɤ�����b�!�Y�vt+fMޫ�Mk乇��4��*�МN��� ,M9���o�=0]��\"y�x���uE��Z8�w�D�FC�s���|"EDcj���x�h�__ެ��&;ztTC)F�G��z�y��7�<)���>����:��n��Ţ|��[]^��ULm0�i��o�~q~�(�a�l�U��Z_1��)MƳ�3\"��v�f?���v�k�6|4�m(�eP��N��GJ�T,�9��/M{U�@\j��Un@Ub<�J��@�L�D�U�#Hε`GM���l�f��O��+�ͫ��&Bɝt�)��ۊ����F��[ND���j��\��(XGȲīڻ���G��$��{�d��E���t%D)<%�_��*r�L�R&�T�U��3Sj��,�"���7���HRB��]� �*���Օ�C�o���ڡX�.�ݱ��x�T���K�HRBg R|q_{}W��ΐ��4|FKT�(�B0������+`���8�M��o�7Kf��^9�j�ۡg��ݵ��v�OpحS�)����?A����சbc�w�,J�q��gm����՟z��)����2������}��2�}fϛ�7~q8�M�Ǎ��Ԓ%>�j�XB���D^�D*��K�'CR��*sT�:."NxA%
�0s{��%�{ڍA�SϤ���|D��b�V����ӏ}2���L���+H���=��m-�ɑtў����#��>w$�-��׿�-G~��v0�&�i9/�q]i�J��Vm�/}뫅�&q���Ⱥ'M_�{8�p�`�M;DF�QV��9����1�jsL�e���r ��u!k��&�Q�S{sK�s]�ճMnǼ.���f�]c�wX�E�B?[�nX�n����k�����,^8�\�:ԋ�Y	�I�������bӸ�V��a�Xj~&y(7�NP��<~�(ѣ�n�y��|������iN�n�c�h�#�7ą򶬂��=��W'��RE�����������(��SL���L*">��;��0v�������p�k���)|�Ƥy�$�v~*��ZZ�.�X�����N&]�g~��çH�:C4~e~��w~
~�������m}�wZ��4����/q+��%f�U5��hȟ}X�N�Z���0��a���4a�s0\�_�k�|�	d�&Xy9'B$�@���5s\�i�n��<���1]����� ������WW�5�Zƾ��J��e���ΊE�|���#I#^L+����>{����K���eǖ���#Bח�ް���>�aQ�0_kL��:�.#�p�M�9aR?��/�?��RQ�NJ�@x�w�TÅ���#ɰ(��ou�H�m��b��KG�gqT��WU��{ٍ,щQBT}\�����qZViڣ�D�鯴xBϽ̫XpM��/r��U���z���LXP-��$]S�m�,��p�oH9\�֐�]�kx!��{]W��Hⶖ�+ ���Y�Z m �W���O���t���se)ZoE�,���KE��h�>�{����
��v��	k�<�6f�t���Q�`a���/�kD�|���⨆R������C:.�	t�*!T��ժ#W����Q�;���Ł�*���2�tJJ9�,���+������Oo[�j�1]�!��g#�K�ŝ�������ŽhηA�j��r�D�t����i_�pi�`n�[m�=�c�D�[�4Vo�B���/��L�����0�Xĵifz�53C�KL�+K����f8S�b�9,V<ͺ�S���ɇ����C/�XϟG<nw��{��Kȷ��6�-�P���!M�k^���k�)�rP��JH�2���خ��%ľ-E���}�jxC��C��2�7���lV���ka��6<���o)��y������GF·����}���Q
�֕�g���/�׳Ǫ4�������_U�˜.0ZB����XX���n����������28Y�aDkY,�n�Q�����Tf�d�;�V10�S�@g���4��)�8�U����%Ji�֕u���K��ֶ����a��]��[F��u��i�>�j��4�PG��8+0Jύ(W?_����X.��]��ΜR�,緵r!�%�����<@�Do��?	�����#�(�%H�n�v���r?'����}�u\.���4�5]����?����m\,�-ض~��o����m�­��ZS�H�{ެ��ӡ,Y�ݢ����0��¥m|}�`x�xu�,T���IM4����iVؖ�_�����Ԙ�(�$�J�=�p�W���`���%/,"k���á��H�'_Z�a�s�\}�v˒o�|r�sZ�`���~���5�#����]ƴ� �9+�l��������P�u5Y.1�+၎H��9��ެ]��!�	�J�/�Y����ܟ9���y?i����zW��DB����}�җ>��JK>�l؄`��bRN��� �x�)¢�<je�չՋ�O��}��|�����1��W'���mu�t³ˤ�u��r�n�wz��WYHt�.�{`��o�;�N���$�{�%��Z�L#�-���d�4�
%���ek��xo:�	�C�	�+@�{a�������r�H�i�e�6uN�֎�����9���u�qV���M˸N:!�I�n$��n��c�u�Y�b��eܸٞ:a�͙���<tzM]v��F�Y��q����E7�zz�Ի;\':��wm[s͹�N��95�K89��ۮ�q.T���G� ە����b�9�v��nl�u/��Ƭ�xs��G2ܪ�W:,�^�5�96�j������/�?�B��f+��ԋW�����`F�׈ ��B��L������DC��0��%��"q���\�=�5�u��@���}��h�
s��Z��:.!20�"\��4�H�b�o�&hTL�M$�R��k��H��g)T�	`}���5��D2�o����Ŭ:�W���������z��Ovc�L'�}�r�kbTC�}�x$kL酔FFX�����+g-�k�Y��zk���X��s������v�E�)�ӑ�:�T�<-���+��01�BA7���p���U�RB߷��A��_~��?-$�	"���=��­~�qz�,���+r�-�C����8�{�+��±o�V4ǩ��Y��k&G��I-�k�������c�o����>�=W�Z&D������-c��D�o��XE8,��Ⱨ�?D�l0ED��t�N��Q�����o��^#E��ݝ�XFs�VG���\�$�L��E�����uƤ1��̑E�g�{U^�--��O�X����T�!�����r��/�މ�����L+#�I)��q��s�q��ऋ9M �4��l�����!t�칲�d)e��s�ٽ�sӍ*�Ä�3NBi��'s����6�n����'�N��\�B�������cv�.��%'nHLr��D.��`��
��[�Q�ݴ���Ǔ��V%�E~�1b�9�V�L���<�Z^>㎔X�5LDlTl�c?ێ���?�=�G��8]&�)���E�{�[0��@��*��D
�\���MT���d�,\#���� ,�ᴰ	!���Ͻڸ�p���{�N����ϯ*�VMZc�>�k�Ԣ�co������OQ?G���hh6��*�=��.T�w7U۰����I�%�Q�NTu�O�`��g~!������j[��{j�a�OK,�C;֑�T괲�"�E�V�{���v}�W���B�'¼��w�F�wҴ�4�Ӡo:��SR�J���+9ƙ2���ȕ�W�Wτύn�C`�mQ%�ݽY�Ĉ([�SW��Og1��]~$� J߹�,Ti�l�6��*焋80�#��-�"��/_�k�q�k���y#��j��sUp��w�~�,��W��3Ǫs>��Լg�����װ���5;�e4���P�\z�֮����*(Le$Y眯]^[�������=�H9&Z�׶Q�V�ܫ��)
��jL,Ѻ@{X7��
&����RG�,&ΊQ6Ր�ڲ�	y7?}�Ր����S�B����ko:�f����rFc��
��]��s�R~��V���?�a�iX�������b��m�	�M(L_/�C�T�R�ě�D�̙L`xC�}T�b�>7c��C]s�j�쫭 f�Ϸ����H1�+�=�����i�gJ5�-H�RjM��KM���i�ے�����z�ҷ�Qb�7Z��c:�$X����X�/n����mT:H��i�B
VYU!Ԅ/�_��>Z�D���}�8%D����{N6��z�J�㄄��^s��b����0K~��v�WN��������=��΀7�,ɘTY|�w��p�=STpF�ia ��.��#��8���˚#������[ǆ���;뫏��<H���u߲��wޟ����b�=�l����qK 䤷R~����cƫU�WQL,�}���F������T-x�FI[�7��s(�ْz�l������j�*яE���u�Ot��Y��-K��kW��n^_k�on�ۦ��Q@�u�d���!�@�[�R�+�����5��X`��QB`�ʼ7�e
H�8�VX*$M]Z�L���G�I���D�}�-w��좾��b]��e���U����kL�.��:��[�����k@q�e)(�
�[OHù�wՋ~h�f��X�� $2��3�mʫɏ�'�����ho��_Z��A�\ؗq��E���m�be�"%H(i���E�I5YP*��{�kDc�m5E[�(�p���r~�������z����*�
�N�SD�S��n�$� �
���gu�H6��V��|��F4�.�7>�ZB��d���S��Ͷ �F��A2E�ڦcN����4%�r�&�m�ָ�G^���L��&jܛ����e��B��Ѥ�T)K_q�9�Z/�>�bd+$�(h�r+���-�����)ؤ8Ӷ�B��8���W'E���U�߈�?j0��DTP?TB�?t�vVP|���	��$��}���)P�dҧS5Y.qĊ�(�{{1V��^3'�n���Α_p8D[��(��,Z}!:l�/�{�֐q��Y
���"k�}��#�0�G\�f4��Z��
K�o�����.��k�����4J�ƺ׭�,Y�[�3�%�c�̐�_�"���X���}v�ӝ�V�8ٓ3&�׷7l����~�v�_�d Y�%��;"SO�-�8Ґ��"��}���i�&Q����J���ٜ-s�L|a�\r*����8�.{� �KV�ם#_5d*=��Ώ��q/��g3g�s�U�}����%I9I2E4��ެ�/{�����m2(��j���jش�{Ɠ0��l� �ܿ����W�E���.�������n�[ףnM�3�dR˦o���p�8P�{	c�+�f�H��}s�%�0pK�~W�������d�ҥ���T��pi�@�~`<���$���?5ƍ�ֿ�4�n���c��o�W�I�!Õg�Y��Bϲ�>"�/�G�{Á��p�����8�i�����Ǭ��q¥���@��V6B���U�&`�d`���*�\���8�s=�����R��)�f��C"������9�����Qq�����OM�+p[��߭ߛ��L�b�q��׽�X�`�ֱ��WI����0��|��kA
���,"Q�������~�b]�,������_�D�5�*�%
E��{�ź�d�q[�΋[Um�#���K�RJ�J�I+��o��0�և�_^���]��)]߳�<G{ߺ�����g�����~D�=��f�e��f��g|���Hg5�W>�E��$��?��[Ǡ),��wp�X%��Z����;�o,K�<�?�~E����~U (��-]�F�]��%p�i�)���9�g�# ��M8b�d�0X�CW����W�/����ZA��sj+O2|����RGFYb���Z_:%G>q�,.�%{�u\,֙M5��RT:q�Ԑ�<�jp�	��:ISUV�,oF#=�ZZi��z�~�����>���B�כ���F��׆�Y{�vԷ$�T*=�nH��u�dk��qѢXBk����/)κ(��Ⱦ������}�{��c�>�{���q�x]0dw1�Nz�L��_�-qAh��G%�0���7��ߐ>���`��~����k�^,�"�
����{�����W;�+K�zr���q�N8T5{)ms}�Ĭ�х�%�id{�?r����(��XP��0�#���5:{~�=vZn�����7��i�ڗ�x��ՀpV5,(֥ee;�v��ĳq���Mǵ����uq�_Ǐ8LQ�FԐBn��6�u@�=��0��^��-��Ղ�ۄ�4:y{Y9�c���`���㧴�g#�v�]�k�ۍ���8:��S�"z�ڶϯp��rЧmv�l�^i�we�qr܇:�;����;mn_����y6�ٔ�(;j���Z���3ī�줤����]�!+]Tx)��8�c���d��oFЩ"��ף�K�j�uNϢ�ֵ�U�/����4�=npk���5`y�n�PkV냙ힸ�\y�x�j���������{����k��`�[w���x%�p�B�af7
�O����o���F�J�|~�]��Yu�0�Cw�˽[�p0�)5"�/�(B���w��p�t��Ds�M��$�^�1t�c�'I�����VG���f��R�����T9�+�-�?�)�ox�^�DP�|M{�eb]/�8�U��S�H�޽.0�h��,J��*<#��+�6�p���������T?����
�$.���LK�lc�73Uqzе�p���`�+!T�ޫ�u���qb�x/r�W-L�j#�wt����E�Y��/���K�����q_�>W���+g��������+�!Y��P��jV��x�#!l5�|ۊIY�����׾*���ݨJ�����Ĵ���.��iZ�4����z(��s�@2��D�ؖ${/�kE>u�� �$t�1���~+��Ӯ��9�Bv���o� C��j��t�ưn�Q��	ln9N83�#�H��"�$P�W�}�^+���](薿l�A�C�����Q����#]{e}dޥGEX��тL��U��U��z.���'@]�b�3��UMv���ՉM�b�>,_H,ܙ#���9Y���8�Ų��̘�[$�e��v�c&��VK'RI�nn��v�W����y�17=ߢ;�Q-�T�[_KCf�U��#G����5���z��N+΂Zg³��VVmb�#�G~Z��Y���b_k�E���*�i���i�Q�Ӳ$/V_���E1�UHꪳ��$�[�0OU����V%�{���Hv�{�,n!a�T=��Y�Wx�U��\ܸ���������J��ż�	7Fm_��6!C5U�/^�׺�����<��1�n��1�}�!��3�Ȕ��_{�R��U�Udj��|Y��#}����M���B�>j�hK��p�%�ـ���A�k�Y��F^��Ö����E �+��|�)2�I�����8&o�����jH�$]����&ʿ}1��� ��j�VG��x��RDML�t�7�����^�y!}���=WD7S�p��%	�@��~���w�)��ԖGm��U�\�����*��Yj����?\�{�,�{�oL�q����a�|�g�*�s���GD��Θ ߳�߾��e�q<�e\/�vR����!n6�+�w�x-(��,�5�-а6�s��k�9�i~��׈�8TH�I	Z&����L�rST��3T�.|�E��(��RYgB{.��U�#�0$����@P������W�m��J�*��ἲxx����2�\�{��PDX@񢳘-�$�	�߳�Z��8����}N:"�R_������\'}M��2(�i&��J)V���x浑�݋��q��v����Hppv�s�5������ݹ�����u(��� |c�2��Q�ts�Y�9B�/s���F����O}�+��8UMq��vE�禩���+�+~�N��l\�u�u��—�"����F��t��%�!~Bc��dQ���Y�	~��i?4��:��j�H�]"i�ܙ,x�r��Z�ٞ�j�uR�e*w�r�1c���i��u��W�J�f�-���#
0�����#5�$YR�At�焉e��r�v����U};����M�_G�����øo]&�QC�
�
����y2 �TD�I(����^Ǟ�Z�ܕ>{-a�مE�}�\^��}Y�8R�5��{9���R�E�%0^L�Kglf�ޅ��p�jӘE�W�|��e��]&���*L[��F̎NʍN�P��N��mL���E��9��B^C�>�ܟz�1�~V?�n��5���Tw��8��_%�d��]��f�g��'!�`�� ���2���Q�ьR\�Mj!o]\Z���������M����!;�mR���z�c�c���A�yf�M�V޴���ۛ�
R�Gy����Cvf.�r��;<�[vN�[�S1�����-�-;SM���ݢȲ��ٶ�!b�>կ%��֕�������0�A�y��������b��j9JQ��.vm��U���e��W���4��n��������Np����[��7+���z��̙�:R{��IR�,!PPn&��z����K4u∏�C���wpI��7~u67��J�N����퓮�{9�#�ʬ4�G��]TeIP���E����,�y74"/)�Ԅ6��m���k^+G�2�imu^ٸ���3��yu�QX�)Vf`@�T�L��h�)ǫ��]4��ҫi�u��b�GJ������	Fhp�礑�6�]$rR~��ɱ)H�sJ �x���<$�x���#����YZ���o��B�M��O!�,����l��{E�X �y�
�r��.�LZ3j�6+�h�p��v:���Tv%����3+R�e���RK�c�Q�Z6f	��l�ފm�y41C��a;�?*Z�Z�!Iܼ��5�M�e]����m�TU�Q"_	��+���i�	B�QIB_X��ޝV�6c�09�՗T�h"�<��jZm8	���q�G4�iy ��D�f�z}��Έ��K7�.��/*/��ГƇݜ���p��JGo��{+HZpX/{��`��eؔ��*+_���%��_-g,��纭V8�]���L�b���ϦIH�
�R�5V�Y�9)��D ���:@�L��s}S�-B|`�F`4QBĸ�$Y��ù�Ǽm�|�׺�0���&��])y�[L�W���*kv�h��)�
HS_}�CZf�̥dܿԪ"E�~�N���1~��ڐ��"ၗ>o�%���<��������i�sX�������([~�������ZR��]��=�N���I����\h�_|�Ù��]��i��� Z��-~Y�I>�.�'��u�ߗAx��Bf7'ۦ/7��� 8ன�H$�H������'�'���!9s.���/Lve`Ĭ�V��w���:�����C�x��#i�"�8C5Yޔ�+'��D�&G��%�]N)��z�Ó�tXiZՇ	^�X�����������#��UC���@Ii�� p���8�-�>F7 ����? �
�`z�ox�k�.|��J��Z�z�4B{��xI���
?&��~�s�&Ô%a�d��4T�~���g�J��(d��z`��wU�Bѐ��4�X����Rg�o�h|��ЊT��T��G�"&1��$�[c�tS�:�<x�+=��_��|dL�t���E��XB �aGn������R Dy�@Qb�T)�	��qZ��'�EK�|MV��\�nW����M�y}6�rZ�٬��,sWI���e����S܆n���9�)�fR���1j@Ey�x��&V	R���S��'�u�-M���i q���-�[]�ZT��gV!ߋ�e	i8�a��N�i�b��+~ۭ�dڰKNʕe�e[�h��z�_���t\~u�
�(�h���7��|�$p��K�έ��v�W�#��!J�jiQH^�iн�����ƛ�� Uvz�D�C0�~�%r�س�x�
og�
�LM���3�h�*Xܒ�������Ց���\u�]5MPL�.�ΑϘ�"�K�f�֝�{��h�[dp��m,�k�Pc�ݫ\#�}�\i�d)�	��:!����?c���K�s����E��ȑs��W����4c`Gw/��D8�Y^��;��Z��$*��V~]���jB"�ΖY��l����F�=�\�����*k��w�F� ��2��"�܀W�߫���l���:;xD�O��k A�Py̤]ʔ�炣D~���+�F7���տ�ૃ���x�:ޏZL=��'ԝILc�i75[��2�֤��V�+m����zsDx��L��hk�4�h����P<����a�P����Šd^g�Z�^�Y�V�S��^�c{�<0����Z�>���X��ҒȾԆ��#wߵp.4܈F"n(�v�t���A92nfy����G�*�߹[�0R-"�"J#���+)�婏����R �:�D)4�%�W��W��kF*"ǶJ�aX��/?�������#-�h���������"�J���:�5B�FA�V�}���dQa� 
����z�p���]ƛ^-�~�i���DÇ��{?;}�N��P�?)R�6Z�r� �7"`�~��E�ߋ?B,�gi
"⍻�#�Q�����ʣ�i3��BVC���'�����`���f�<�]�������E�
�:�仴�I�{����u+�b�^��Ͷ�5�f��s�>>�M7���j�m�BX(Ia�r���@q&�@�]�������{v�N�[����6ѷ;��7��_q���֥�Jku�cl	�1�ɑ�S:�g����x�`�9���Ǝ��m]7�v�x}�sU�c�s�۬��4����q���[��E�t�툻���W=]�%�^�`�<�m���نԬY�*\��nBm��Ξ�ഘ�,]�n3� v��FFw"vW��vtL���V5�
��;��шͮ���mط]��g8�Y��t�45�����7�Gld馅%4�I���HU{�k�3?+ E���'�2��K#\��|#���`��TD�Q��}�O�,=�<���g=���%7%�ۆ+w0�߷�+YmQ:ؕ�JE�{�&E!�����̰�RE sU��BR�Eg�Wޜ�^��+��o3����Ɛ�ϳm�`��͝Gϝ綖�H�,�D�Ih�,���.���WH`h��(K��6�7�s���>�����gm�p��>�/pw��/��b�4pt��	��R��asZ��U�%b�)(`-�����gEȐ7�f&/�{Ԯ2��|p�rn)�����R�w���ד��;��,�ʲ/��|F���vE���s��ZY������ی8WG?m�0���� a��8�M��W���^ʒ����<�&<�ֽ��!�������Y���EG³���½|(�{��b�ŏf�,��Cl@�ణ������7�Y"��;qE�^�{{��g������v{��4G�r�(�%�!�Ʊƿ�Ͽ�����e�3J���&��ݴ�R����f�~��<Y�O�޿�F:�-�c�r+�����'}0��g�p��#�zlP�u�LA�D�q��z�w_־����ۑ.�)JwӼ�]1���%5� �MO6Ec��	���8Jx�vv�V� �����tmv�N��ÛRrS��eUUy/#DR���!X��)z�{�ʸY�I��--j���[�+�)�4�#6V
�o�izg�T׮��U�y�Z�Ejn��A���tAooޗFw��ja|6u
�X�sK<��M2���j� �w�K�M���>s��Mˮ?}�~�=�>�W�O�ֵ؇A�I�#��*z=�`Ę�4���娬����f�7fT�e��z�7l!vtQ8kZA���pL��6.��v3T��ϕѵ���\�0aϧ3�8�H��\�I&��m�v��=���i�(��֠ �#@��aG9��(k��q����{�;G�՞��вߺ��eH��V!u��I�:��j��	ߥX����3�Ѓ���{ά�Ѣ�r��M��/��ՠ#ED���=Y
o�������������e�����hH���"󽺸�%�1I��ҡ2W�Y`����9ɘ�Y�H�|A��9����795T����������Y��DGS\�s��m+�`�>�s}Q�pfZkHK��+�y�Eg��\h �'.:�R�[e6D,�eO����I4B�D�<�ힻ��}iv��U������IAM4��ށ��JE�MsU��ѝi͹&ڔG)�UJE�W�g��b �w�][�c�y�N:~�,���{��k>���8�����}��RA���k�P� �Y6Ӷ�Z�(�+��k����.�p�|��������ߦK˽m&ݢ��2�æB���y\�n���B�z{p���u^pn�,�&�QD��W� ��j@TP�P����}�����M���������O�=�w�����J��d��	�a���o����p}����I�tK���b�=�Go�\uK`+2��2N&Jv�e�sI�)���9")7+��,;0�Xp���҅���no9|V�G���6���|�"Ζ�Re������V${*A>�B�ёd&<��hUY�vq'��he4�/B~���7�-���O{�k�r띏��1x�Cf�p\П]2�4���-��h�\�駅�8��$a����gE��t�,#���Xp�ڢ�W7ܬè@>̈��~��p�O6�����)����g+�Y(�.�FG|��,��U�z���:��j�����%����ie������;H��^|�m�yр��s���#� n�m\=yI��
ImQ"	�}���x霻�^���2>ưbӅT����]c&�p�ܗ�KO���E�xb��]�f�:2kwf�ލ@I�9��J�_��}W��	i
E'�tؕ7S���g�9�I���O��/����}j��: E^n�+���i:q��V	�[�y_�-�
i�H�����4c��w�KL$�$J��j���������͑��M-�>�$��)ʡZI�B!��+&l���]��*�^��P����m�$r�^���k2� ��ن"�]d�-|%��}����q{G�Ai/�F2��l�5ը]�ݨ�y�Ɩۭ�[X�{���\ۡ��+����ߟ��7Y�c�ވb���H�޾+�4�2F���~�Ƌ��Η[��kܬ�(k����J��@t�����_����m��8;�~��K[n0�q���=�!}ެU=���تrUmi�(�W��Z�*f�8�����ã�����U�$��Y��o��i񬿫9��V�%�<�f{�Dﷳh\H��'�V4�*��z��0����f���͢0d1��{>��@
$c+��<��p�r�� �"u�Yb���=<)��L�sUkы�(�[LG��$޿s���:\��
|�@E��(���xU��0(4Ъ�����o��[��!�=�s� �:)Q]��qV� �~~��3"���Gk��j��	�ۿ�E�k�jX��Y�	#�'���j�����Ac��A��L��;����ӧ�����;�IB�u�߽�U���|��<#�R�K&�R��H�� r�i�	QD?t;߿m����D�׹W���e^��2t\{%�-�[�t=���c�)s�Yˍ����z�}���5��������>���HE	B�8+*Sd�TP�M��d�L)H�F7}d�~�2}�DE���=�u^ 8�v*4�P�8`�yO�z]����o�}��82�TB�l)rb��z��1����n�{J���!�)��V�Lb��ތ�!�_�?�G�`�Y�'~%�n���vݵ`�6$�����M����f]������g�vZ�;=]�+����z+"DS���Y)���굄i��|�S�
D�/���b�<��ڴ����iYC0Rf��׻����
O7���_��%s~q(��v��@��z����"HhW���V,9ƤN�"c�}��⦩��L�����8G����X��e�.�+�W>��N�Q�G�g��xH� �JϠ��*��r����\<a�W*���8@P߽��~#A����Nhy�� ݾ�Ջ/Ҵ�^KI�[�qMׯp��H��Q�e��t�1�0��WQ�}���YRX���ޫL��O���q��iM �s`����p���^��㙞�>qt�.D���V��6ኆC$�3���f�8�@Rf	X���P���'2֐�Q��	I�<F���.tN,?Y�E�����?��AĘ_��;e
���_²��..�L�9��%����C?>D�A���R����Z�w7Y�Gkg���Y�@R�ݤu~��/�Q�>�V�!p���.ڲ$!r�����&d)>)I$5y2�� �-��,LY�͠�=Y�`�u�i�-	{�6�!�3���V�����ݾ��0���*U�,'3�U���H罿b�p��ȪY�e�BbeE��qZ�h��%D�ҕ ��2��*�tJ_��I���~�nd������h^
�QH��lJ
��^��*�%oǠ��ʴu�=�w��!�Ga�Yڲ�
\��ˍs"��Gk��l�n ?Q2���a�rJ��@\��Nb�Fs�m�ke����ۏGV6mr�YK�0�j,�j���k��l���c���8#��:���s��$#�)�e�2)��f���9��sسa�݃7B���(wTl�;G���O��˸�S�Sɥ��V璳��&�p\X�-t��X�i�ݝhvl�q�v�x��Y�j8�L�BN���uPL]�;';�v�G\�m ���k>�l�\5��R	�Y��@��sӍ�nw��{�o�o�)�KL��2G��{3�'#��uج�#�1"�M���N,�$�'"D5�9K������j���L��˞㏉��!Q	�>ڵ�ڥ �����$�� QD�����.E�Ln��T�u��2� "H�`��o޾+X��>�U��=�h��A���M����1�rN4߫��|q�짎�7bb[&��ЦoޫH4f�>GC�$�T28Q}��ӊ�kC�,������#rg�B_�R�dx�w�n1��
H�Q��x����+rou��ٟ��rcZ-m߻�q�l�qBL�h�.��T�0�e]� ���s��9���s3���>+��l�/7щ��c�u� ���^,-�9\V�`�q¸�H(�w�?�����D�@Ä.����]c{VE�3��đT��:�~�%x��U�KkL_ܘ�M`��9V����?G�aÑ
 �!���2~��B�$x� !�n�)+ f^���=�I�	�f�]�ƙ�x�����ǂ������rziN����K!�"f��-�E	Hs�V�� R*!5�Dh������[������߭1	#�5e�F
H��qZ��À%����&Z`��[�$���~� ���:.	�}ۑ+�ĨLA�������a��9��!�+$��7SN~����08�p�7��F�ݳ�Z���wBu�i�.7-�jjf��||0	h!I�pT/�'e���LX��?nz�nJi8���`�_{y�k�����Y"��&[baO�q�e$�=͕��V�7?�Υ���x��+�ֈn4I��9��G�	f^RW-�x`�[�^�6?pj�
�u5J�@�qYzR�̬$ָSM,�O����a�K?���j��%����{�F��i��KCr"�+��S���vg+�;���� [�w %���s�Y��k�K�v�W}��v��?>������U6�%�[TiQuJW���V%���
�S*I>K*�@-���έV���ȋ�������2?N�Y�
*�_����=���"��G ���"����`��e_���`�4�+,_�=�ϛZ'�/2�V��O�����>��g�Q���+��߼��h,{�z�~�"�,B���᦭u.(�}^���#H���ݫ��������өQCu5X����J��a��3��^��^V���u�<n��U^��(Zx�uȆ�ƮS �����zԐ����g�{��-�n�U�FV?�y�(u��DkC�Y������<~�M�����#�4B���y4?@��FSR$ܞ�#�\�-	a$�,_s��in�R�PI��(��P�D4q�y9���]��D>���,��K�G�j�dY߮���_9��<|x�6�o�0KL4��fr���ι���7��X�/��SC鿡w�����5�ڷ��C��5�o]m�������ÓWk�(�۶�xn�:�c]E�L��<��� ��RQ����[�!���e�����KG��zZ�'��F��vʮ�X��U����򜅌��e{�U��۞9�*��i�vl�
��a�b�����W��f+��妈ӢSN����$�,�T�
�[�u�������0�ز?�+�$����or��!Ӱ�@�Wp�-{�ֶe����1�Y
HL�R�˞��J�ݖ2����ㄆ�΋��u^�p�k���r�}�KYr��ig
E�4wt��K�U#�:USU�-8o�у���D���{���p� ������,�CѱFW�~�����,J[�g|ڟr�O*�w��v�^���j����8�\����F�Wj4(�u��:RKi$��ޜ�y:��Zؾ3�k�#��W�__�׍�ں^�'J��򎴙�b	>#�����ݫ��>- vc�b��'�����u����HI#��f!օ��ᴴ-��<;=��L,g��:���V1[a�h�M	���M^�U���U���P/
q��z (���ݲ��7��@�E�X1�^�%\�QZ��~�Z�3�.U�q�C�7�g���p���vvuܓ�B�>G 
��u\.�E��dn�&'�A��~��~ŷ����9^<1��0��$��<��ݺ�Ӈ:t��"Jm��r�Wmp{�0�d�5������N<$b\����?���j�1�����?�`���-E���X!�^��3p��en��r���Q�*ƨ:�4���tM�>!�ޟM�k\��gr�0�+#�l�@X���j��z�g;+	������(	��E�;�����^�
̾�Ko�j�}Sd{y)rSf��+;�+RF�i�p��U-T�>~���**��A#C���h��䢄���-��x�{kc ��W~�v��� �R�%�$� Ͽv�@�B���å�C�f�G$���+��� o�����0�{~�Z�]8[}���պyb͎
Z�a�j�o9F���"����@�.�ڣH�x�V$�{��!i�Bd�3��H��D/��qd-\p��j�*ww؇���kLAg����6X-��YM�A��JZ~d���.��#��D��)&_vaY�֍���R ���$��1-8&W\��"F{|��Ϳ�o�Y�ޯ���!|���X'<�mr�d{��Z@h��⮽��B�����֙�Y'Abj�e�ڴ��n��i|%E�~�|��Σ��2�f>o5^�͚Me��`�@m�!����b�%L_a�c4|1�����v��6q"�Y�s)Q{�0=[�����<�P��B��j�[(L�o쵦��i׃篴*d�Re6��[�_	���$ RP�'-��ެK�s�UG��g�{��Ah'��ҷB#>��t�4��I-")� ���VȓD��;�Ԋį��5�p�����ã㏺Ꟶ��q�r�a�ǽ��/&��Maj�v���ګ'�9�S�GN�;<�q�#�^��;�E�G=�uD� �C_�~n��}��! C�I���(a$��SB}յ"�a�H=�⾈g�1b�.z`�S�T�?r�0��{�}ߕ�2�o��}�+z@A9�/��E�nd�����$z[��(�Bȉ֧��C�����;m���Z:#�:$U��f(�l�g_��|�|�Fz��ix��Ķ���"P��߰T`����:a�'��U�	��IB�4}��S�Q-�W^�b�֢D�xk�k����Ҿ��/�cM�r=�)T����[V�8.�ѷ_m�	ֳ@�@f.��Ea�$�M �?�O����{��W�=L����"���{�ú6J.I�L}uq����X*#O��TE������|\�u���zNh1��"��?B��>"��~��c��$���1|��-i��^���-\s��B�K��S�}�}�I�d#n鋍�2^z�i|c繳�����P��Q�`�L'� };�X�Z�3�=k
\��(�UVuw�Օ�����U�z�p�����y�+��U[h���nuL��M)$*���f�$��f��F��߻�U�ΊL$���D��q�F����s�n�l'FM��e�Y"���>��\t�x�XY&��b����~�Vl��!���?&�y��w� �Z���I��Z/��k��7����w��Vv�ɱo����T4��{�WYB�e����3�J��a�^�(�p]�Ρx�l�2n��U��Q+ZUd�L�reL�O3rE{R�o6��NM������mЅ�*�!h���.�Բe��bΒV5���4��@	�o#�-�e�k&,[��W�����������[ݽawS��ur�FY.�d3�1gl-��o���.�`5�aI�RN�E����nF�0o.�Lnnb��*�8���%�k4vT��\T��O5�Mvc�׺��%eM��9s˘:1�t���n�{̳�+Jj���sr�U���j�gK-�ݼ=�|;"'�;a_{N�C��6���}=���RZH��,�s����Vt�9>���a��_N%I|F$��+8��A+����{���S�5�+%^f���de�ë�T�c2V`Y��٨r�b+ןm蔗�fT��w#F��R�4o1>���=��bM���v��=[�ע���Wp孒lZ���ea���j��ZV�xJ�GvK��$�b�n0U��zaM�r��kU �"`[�?n"~��������^#|�V:9	�!����`5�e��%�.�U�7���FfQ�WQ#���0(��x�ZlO���	�qnP���"�/H�WU�iY>%�؃Z�._������LS��
n�vZ�T%z�#�MՄ�q�zX�ME!����^�Z������C����|��0��@T]qR��� +T�h�h�R�*��ĩ��n�n�{m�8�ᳵ��;Ś����y
�ltq۷l.�э���f���X��ŵ�^��^<	�&�y:��%���i�m��r�P�P�bm��\����ն�9��N���V��J-ǩ�݌w6��uk������'5;���ݧi}9�%ϟ&�����ͻ]��uۓ��y;!�g<w�x흮d�v���j8�ص��q�%��p�n6krj�ph��[N�a�ۋnݳ�����Sp[[,�絢��;�o۰��<������q�u�\Xmך+�í�H�h+���E�6�	���y�g<�WFn�Ӎ�v�m�7H���ɜ�8��H��܅!q[����F�Z�NyGc���];AuNL�R˽���[�������6�88z��-�!�.1î`w5٫r�^1�k�Q��Н�.�Sgn��N3�غ�;��wF��灈�����;8;zB�]t�7�Jr�^c���iv��s�K���n�{p�#��*qۇb��/�R��H�ݞ���d�z�mv�m�p�ܼ֏1�9�4��h^8.����n�]�;��g=�$ַ+' �ڀ�g+�u��^����q���c*q�m�n�W�'a���s�\/(��
��%1ȑۏQ;�ǳ�A��󵪰���Ӄ�ppp��N�u�DWn��h�v�O:�N��}�ɮ{l9J�8�򚃈ݨrs�%֝3q�D�m\ru�"�vF���<v8�">7=�k�k��x�FW<��1��īm��.u�f{N�2�۝�k��:gV�lN�_n�8.\�r�d3=s˻=v5���zگJ�1��WU�6�/X�t��F�����N��y�m�qsZ��s��kV��r���ܸ�/O<�:z�n�ۮ�!�z8���HtK͝�"�<Y��۵��Mu�6$���f1M���CsEK��;�;ڱ��6	�s��h7���'*����x�!�An��$��V��d�H��ѭ�o �q�8�nwv�b�u+�0N� �k��`�qo<����[��]�����֮n]�<�V�[�X,k�45ی������[��Iq�w�=q�,{s��[�ώ��S��g`��i�"��Gr�iX�K�c ��j뉥jűO��-���L���gW�F��K��u�kqb����\V�	��ۮ�9�^�D��n{��E�p�EV#y[l�z���b��l�٣�\��l[��E���^�JP�m5F�[�M��v�ΎK����J�F���3�C<8�ȶ���b}}q����=M�c��]�ǽ��?�ug��{+�͐�h#��[�RS�J�[V�?J�1�>�Vp}�^�'���z����A|��_J���uA@Yɓ��B�����t6oOfu�FқlT@Q$g���,I�@��4
pdb��M<��a�'��\W�\maݵ�&<�:��W[�9h;���er����ف�,���뽂�|��jkv}*�"���HD�e�.b;C��vo�L�͞Ί�_�ɩi��f��u�
���o̷G�6�~{��>���#�5�6�IT�$�!�IJ��c3�y+ng��`��hQ䧌�E*�}~�n�:A	��g\��(�)�e��K�����@�mWS����9:��D����u��n��<�
�˴���:�Qx�J�1�,c��ճer���I��i]�+��~eS�D~�v��X8���@�����$��^���`��es׌g�l1z�q����o#2"���Å� �0�����f��.�Ġ�>�sr��L{g^v�{fL�Go������ww��Q�Ƅ���ϗm�z(����
�r.%z��њ��mf[+=Il>���kyè�A���U^7���Ux�]P��[�9[-l�����w��4$��&�\� bՕ8+��U^#=o�V�6�Vߤ����~�oI����H`�hUSDw��>񄙆�i2\-��Cؒ,���Tw4��^���F�U�{J�b��3��h�q|�Hg���3��4k]��<r��$.�ܭӦ.�S<{��L�E
����K*��]H�v۫����m^%�T��z������$B�-|U�R p�&��o���o��6�ݽ�^�Tl�� �Hٱ՝Vg�o ��hRUOÀ��IP�b4�`�77Yb��!ۡ�řo>�]��V���nI����a�qD���:<�1�):F��{K���7l��e�����)|��{<���_3W����ǂa~��6J\�E���(#rC��������v���_��ݫ�|�,9w΁�m�ɖ@��*ytݖؽ�q�5��^�sl��K�s���(����F8�rX�e0����3�꿺��Y�l�J���x;��z�h�}aw�%�?����i�j2�Ү�r�����3�2�̇x�"�l<�:t�
��͒-��lo�:к\3{v���3.�w�U\��1��w�9�8�����a;��ՙ�r�}T��ICN`)7��I��'s��dܼt˚:{;}v� ��>��KR�v�N�M�o�zn,�M.��w�(�誶׫Fn	;�}bǝ�P�|q����9D��V+�u)5)��C�n���o= F�K��+^�_�_nC^�.�V�K|�/��'T������JW�tj'o��X�>?m�sϴ8���G]��۞�ɴӘ3k��wH�mú���.�.�6О��١�`�@%��ޙ�e&ӣ��9ɂ����4� �.�����=�"�<u���O{��A'f�wq�;�)j�0(��#re�l���tK��y�Q��pd�<�t,��P��wu�]ʇ�D�I�x������/�k<	=(.�剫��;]�$�[�̐\�颃{{\<�EK���4FR�\��r��{���ޮ��!rq˰��}�>	PGw�
ܳ)#_g3���b0�-��^#+���2\������j���̷�WfTf�:UR�͖z�%Źe��y짠���^�S�6z(�[��Šv��^����e���o�2�V5Y�ur��̵}������i�	��t@��j������lG8���=Y�O?.T[��%x�hڈ1�^U��B���d[�o��#j2#�便Q�;�
 �Ϊg���`Yl�<�,����6�ҝ���r�r����v�JŴD�����(i⛒���;��Dv�^�a%鍹[��lא�3}�����e��d>V���~����8,��c����Ay�����=��~��f��݌��IWD�"�P@�i�4-��)��;���@�e�"+墈S.�ˤ�"�l��{y�ƏD�E�K2��]�yz�̛��&-�$`�F$|2&S$�"�g)���z|U%��|�ڏh��Ҷ�n���9�eȤ7��������~
��Z��$5�3;�Y��I��4B6�a��~h$�|�,�xm݅�*�x������Ƒ�����R�Y�\s�]K�k�H*oB�H��uVd�b�~6�/,��hY	nO��֯������.6�9~��؝�b��B=����+8s�{2��+�[ʅv����+#M:?#:���';W��&����|w9�S�8x)W����+��_:��ֹ:��+�yuoJy��h&n�Mg"G��wձB�d\���9� �Xp�Rg��vL\��۳uQ���\uv��3�^&ǀ۞S[��n;n��;vd8zxy�a:���J�4�t��WWKڳź��8��;�6�6��=���Zv�e���/MH�ѳ�\�=��ֶ�&����6�wmjxI��c��s����n�@ʺ���]<���v;q�\�y�m��H��qn��mv͵��.��f�x��0 �S�p���=�����1�ivi�hWv&�l��W �q֖8{v)vn80���צ�H*�ˣ��b�]ޔ#DX��b���p�=0CZf�F8+(ptR�]'�cs�2���޸�N6�p]\��5\�~�:<�5FwL��J�����}y3�ǜp��}�d	X�EkV���z�ǽ���R�H�'��cX��Ƀ�H�k�餥��[g<�T���Qg~�>toM��n�����E���ҎSx�q�����i6�y����a�k¬��(�d<��Z�Gn���������c���j�U���^�]���������v�_��[��(f?��Zdu�	5�[t1�����֛�{Ke�U޶�;-M��n�4۪v�P���rd@-���m�]5`e
~�j\	�c�{�[`?2��:3�E�ca�XAݼ�l'��L�n{;�nU��tOs���.�E ���C��&M�B�8�!���;���z�|���H!B�K���؂F�M��y��zKe_I�L * �rJ�FE��˶�3{�]���8�3ٯM�زr,�Gװ�R���GJ q75�Kt�0ܠe�p��"E�^�]p��(��$g���M�rmmb��7h��J#ݺ���c{1�p�r,]\�:�Jaab	E�RnJ�K'�D���gUY����[�U�r���~�K$ҕ���M�v��׻�na��H�ç9�1�HN}M��ܗ	��K��t7Y훮P��]o��'\e�[>4�u�ǘ�¤���=���i������vƥr�N�O�g]ٞ�5�FbD�R���JA�v�Ώ��(���ڨ�vM��ە,�����w;�n=N�N��d���̖�{���	;�ġ)#,4Dd��pi]��%���\q���=Y�og�.uF싈n!�~m7'<�m
����J��&U1y=ݺ!�<b\=�BEӺ�����ܯ��ub�o�aC5��V�W_W�dP2��I.��p}���̸*˕��������J.;}����e��u\��_-�w��c[k��}4tG��1����M��:�!��էӊ�s���p�cV��)m8}��Q?p�<����r�6Vt+
�V�t��sX��p`��U�%fI�;:K��*F��T��u'��R�৺Tw\�N�s7��1��gl92c���[��0�C�P� VKWx���fgk���v:^��h����x��'�{�I�.�g���!T���~'����p�����mT���l
l[p�P
rv-���q���}�yK�-�<��>i�K���h`�{|�TN��n�d>���ו!�b��r}I{����~����=�}|m�ڍ<�F:���u��m���r��1j�-���\q�qWl�4�ۑn�_ꆁ/�L�0�f����+��Y>}�ĦR���I���!��į۳N'D�5m�F
�Q��NI�
H�i�]��y���2�wߣ�"v�`㢥v���V�u�p�:|��챮��TyW�u�9;1#���(�ޞ���3���UT����ن�c���]���o5%v�B�	�ݽ`��z�%I�R䘍���#-�~�G���J��V�Ѿ�+}��	"�(E��؛����һ�R���0V\�E�nd'x��c2��b�#��3s�K��HB�3��B�nG�!Dr]��Sj&��e�&�[�py���Vf�t��MUy/T]"��>'�pV�ۻ n�wȓãa�cQ����9#]΅{�A���X����W�z�{T����a8�vfs�W_g<-Ǝ$[Jd�<zk�;����>;��\�5�+���S�g�l��y���u�͍�Z�=�;�8���H��%���{0xd_=^Co�1�����|��Rܮ�s���Q{����`�l�On�ų�𮝌݃(� �JJ��jص���`��wкI�H,��U�#F_B�'\��*�Nf�{��8���F�hM�x$��^
�U���`޾���U����B[���8����� ��B'+_L6Md���%R��8�<v�4=��y{z�d��T������	uT㠓R{�Ek����Z0�%�{�7�Һh��v{.�G���Y����x�����O����FqL����IݐW���ۗ�V���v:��8I��ԄE��ȫ�����g9�{k���(�؋�F�Ķ�`��ey:�	��wt�eo�T5�<�6���ܬ�0p
��Y6`Z��g:���tEL�f�X���N�l�qt��gfP��m��7^��g����%������������8��u��mlϣ��j��dE�,Ʊb�#���r ��=!*<��&�r�h�^��[���X 	yj�q,n���W[� ہ�M�t��ޯ.���%�ti��^^�<��n�Ս�vm�i�`39zpom��="�/mc��erl��s���ɯO��麖�cs;<unx�rt���p>Z]���YI
��Yv�9��Y��;S!�;XM�9��9����.�i��U�G�{xi�0�P�T�3�a���~ߜ�G�#F`���($����:���[����h�G�v
�u���K�xy���*��P佰}�͹��<���QB���gb!����{`�2�V���:�D*ʵy.X�k�Q�t�q�?X�ј!Wur���#�<�̕N
�q���ăbF���rG��Kv~����лfI������a]�b��2��ئQ��{��ə"ڽ�9����:a5��܅��lDZA� �-��y�P�eb������z��7s"�<�>�D'4�R�=��hr�u�N���������^�n�3Y��Ϣ���B���yS'����r�L�~��K��fY��gSQ����o�W� ���@����u�|Ȑ�%?p�5�5M����N|g���&z8m�l�جv��9n��71�.��0DJ"|ۈ��h�$���~�ӭ�v�I���x(3�����v;*�Q�����p�	�zݦ7����p>��{׈�XP�P�#r:ÞH���p��؉@�^��fV��gvm.�:��'5�N}�Ѝfq�&�m��؀X�ބ$f0C��At(�I�X�N}}��{�hVQ�=I���!�����2���q�e2zws�6�+��{���_�';�r[E���c-�ۂ�`��W��{=�s���x2|��k �ů^!��y�*˷�[�B�4���dxs��ӧ��'�(H�P��D�l��ڠc��=��c�v%��ޝ�٧�sj�N��.,��ɇ��/(�%�H7����&	�����M�'�Ά�	Bߐ�H�/�wZ1;n{«/�u�AV�e�I������!Qaԕ]�������,��ղKc{r{�m���
|�!8!�3(��f.���Ѷ3v�q`�7gW�v�s�4A��$(�jG\�ю��3y��m���QI3��o�34�M�o�֝�c��q�j�_j��ܒ
w�U����<� �"E2��3mЯe_����³�~��68�U�/� ���2�*��N^$su��-6��j���i�I%>�Ř#�7��W�_��(ὯF�)����O	Lbڶ�-��:��窥����f|�K�!l����q`�-}��s��k���],�Ux���[TxNoJ^ѡ�1����p�o}�2^R�wI\�z��^D�!� ������ɖD"��ԧr��p䈬rؚ�O��xL�ͯ`!u
��t�!���Nep���M���M�vt�4�4����NN"�E�\f�R�f6c�h{�Ű�0.	�iӜ��&{��Y�$YIWh�5Qֲ��X�z�ml[Z���4޲`��[��˓���8�����]�l��7�m�hb�"��x*�nև�J��St%+�6�Vw���:1di�ӯ-i�\z�%��#�6�e�a���%n�Ys�zܬ2S���Z�{��t����)�[�i�=l��w;�t�ҮF���\QL�;�%i��l�Qn��l��y�kׂQ�_�[!�w�pҰ?����s6�@�h�84w_K��[)_�a�z.v�H�~�S���iW�!�YE�LjK�s�<����^Tgj�u�xV\�8���^��^��pO�YF����8r�K:��Ӌ��Am��h4�瓤b�٩�[p�&3�w���W��m�uR�ѣu��>k��,�u��MX�R�J�[�/��L���?��Ūq[��kzu�u�ج�U�죻)����.�m��g��VV������m�]|N��o�n7�ܬ�fL�1��Z�j�ٻ۞���f��c��Ҧ���{��tp(OV7
dV�χ^ԙ��k�jv/���<:!������ ��WZI�Et�s��o���s��2���f�����Ze��v�ֿi�L�D�$-8� E[�q�F[�:#t��Uo�N�nU���{3LȊ*#���Pb�@�>,x�<���r����Gz�I"j(�E�QǶfʕ#Zw��@�<BV[�o�J��s1��y���kb�V��u�c���mW`��|��߈>�;x�XU��q�9�7�����.Q�%�m73��=�Mb�8Wmn����)d�||]�֯'���z}�������vG�B,]&U�����b��}��&���u;�f�Sq�1�G�E��M��������z�D��d�]/���V�-��f�6̣d��΅"Վ����ξ���7��ѧ!�	�jG�_!`#��wt��#�QaumXԳ�sEu.�9Ӈ������+kn̩s����6vVr�6f��-�D�E	=����j!���Nz���Z��R'��
���p��+:���)�zo��"���N=F9���H��NQ�2�E��G���Aa~��Ye\dw�{��15J�Qxq#oevn�}R�1����ҊH��0�o-��Y�|�)��rA����OyԢ�({�ѣ���dň��A'��̡p�����);^�1�{0���O��_^_j�Wa������+����n�.�z�-I�O=m��v�A�7
�O]9ݎɗxcu���v�w)��I�xw ��ep 3P��\����'D�W�����r�VoU��V���ބY�}����/AGoHSiG����d�"#n<����QD���o�?W[[�ܩKr.;���+�l)ڼ!��A��\MN��gS��9���^Uw2wjϓ�j3i@o%3B�T��!X�{�{c�Eu��xw��n�y%�k7�v���%�/��;�p2![��M@�&H
��lnTZv��P]�����3�
�>�����{1m�2��Cc�)Ҭ�L�vӹ��<TӖ�݂hr(�l��^Bħ�;��S�;��.��N�#v����_���;w >�!&R��x�g$NҎ������m�Ȼh�!�6�eba@o�L��Ǫ�g�;en�c��썊����wL�Y�:�˘F��)�1԰˫jI�:��yX���
���
�e2��t��!�H�n���p��D]��:(��\�[�gt���Żm�DJ�zZ�%q�#f ��tn�^�*��»nKD�pX�[�Y)�l[==�Lmݹ���n+����۰WI��y��v��m����ݨ�q۞5�n�<�r�P.�mU���3؜1��p�]�OvڷB�wÝn�j3������'��q���f�!�����{7��67�n6�)MMv16�[���u�M%�'Q.�vv�/�[��f��1u�qg�w��9ԃ��`��T2�l�݃{P��Z��U�������͚�?8��A�>�D*��_��x��k}�/�qO؛ݲ{!��f;�r]\ã�Au� �EW.�/g��svW�⺽)��囁+�0ā�����'(��-p�^���h�z����{���6W��Q��Mgd&�S�#���BvT*hGu�}���j�	H���kSow��^M˿O���P~�AG{���4j����*�&͔���y0f��>�n�~�I".�EfB�+���$�����^3���+�!����ylJ�2���o�Ia��,��+uQ��Tn<��՛���$\u���f����
&Ѫ�φ����Zь����\���)�����x�W(v6��۱\�9j�I�X)������+b��s�v`Goz���G�w[ҥ�����/�Kk�HLW��|1��^U"��۵�$�HD��Vlyb�ϻ�t鵞��E؈�qa鹩c/�ZY�IU��R��Z��o���A�U�V��Ԃǈu�6kz!÷b�k���+�\����/L�]l������9F��}�.�k=���~x��,���fo��v%�����{��ڤ��I�AY���t�&n��i�E�uOw�B˼0o�k�۪5Բ�;+�����nP�[)�|���	I!_Dܛ3Z����im� �]�X�>��F�`�������T��k��N��U{2�Y͔="x��)LGb�wv�9����HȤ�ǎ�2�M�n7 O�/�����N �s�U'�3ۼF�^���ۖ�ž�}�Z�����MD����u���ѧ"�s]���skM��a��ണDi(RNI�݇����c,Ʃ�$"��:�MDV��g<�ǜ-��I�-F��c/;�%#f����u8	��-E$�c�>N��nuK��dD�t�G���u�z��~�۝Q����I[��=�������VG�|oA0��h�юOc��@里'��Y#����L�t���Uܕ��b�:��̣Zio��.���U�����V6!���K�?C0����[G3)_T�׈+n��i>����1S޼�
͞�V��9��mn��y��>��[�8"0�i��>���������5��Y<0�S0�n��O)�(oe��K`Q�,��=�
��(�)��Y��α�@���M���9$8�=U��Tgz�UZ�f��C_�>����-ʾ�;]�C@�y{���3�]+B�G-�=f�ޗx�l>ڴ��^�<l���\�v�Ihp��t�wZ���\vz1�m.�ۘ�ۍ�4�{=����tK�Xpi�d�{���(1U�pV��<�s�)]�Z7�i`���;�ղ�Y"��藅>-�cA��I}�/�Y�r~�)0��߼�f�壗;�iY�����:��8R"w�����iX<S��OE�0��m�}�X��!'/yhhEFƜ$�
��z1�Ju�r��L�h>;��Z���xG���#}��w��>�Gk�^��U�e�t�}nH�"%��}G��v��O{�`��l֊vQ{�4�e�h��}����H/����AY�4��%�5��z�ndi
Q��w��,��O����'^o<��XXk�D��Z�1�iKzݹ]�}��3��O�l��B����7�*i�%4"* d�^ �9O���d�~������s��ӭ��?�t�;�۽Usޔ;۾1Ldh���w_鍶�?YC��:z�M����Y��h�y�����c��؃]j�읦Y��p+}��h&Xc��^wW���jnk�}ϼ*\����q�r�O��0�>��~W¤�����O{(f�+M�P�\ eYÀ�p�o�n=U11�2.o�uN.�H}N|^�V�銷��RՕ��mM�}�5���gn�"�:���Ţ�#$�BF�Mv�w�~�;���62�ox�4x��{��+�����j��=�徏�)X)\�yLv����ߓ��Kf}�H6����I�F�����H *Bܲ�!٦��M��/c�;L?uڻ��[�	�����������w�.��$�J���K��q�$NIV��Q�ʳK��<�?��t{��֑ϑ�йp*���W�T��w�x.a$x�Z巚�Ow�7qqݠ|;I�! �Qb�W$9��[v�M���z�{���Z\����(]��|��D�KvG!2&d��5<l��pN��z�uƶ�r=��̜�BS���r�x����a�#�6���quF��U���l����$-��]Ԑ�q�]�<�Z鸺��L�X���1�X�-�s��y��Wx���!�-q�M�ē�z�p��cZ;uk��m�% \s�l�ZO玻�[����ə[]O��8aյgk��m��se�ۃ�.)��К�k���	\r�:��0�Нasv�^z��W;F�q�3]\gO��Wu�n}o���;H�'}�x+s�2��x�
�~��������)J[��=޽��=�����e�q°M���e�a��yթ;�:���ISU�o����>�������M�߶X��]�t�������$�I���~A*\�EƊ1��7�7U�cl��*Pꭻy����{�`מ��������f��^	Ȟ�z{�1�tA����s�˘QJj[pc�C%*ҹ�ܗ+^����iڶ3�n�u����.��}�oý���W��ȴNu��o�������˱!I�Q�a!�"i�.�㙃��ga��qt5��c�{=�4�>p����l�x�#A������ks�IU#���g�>�X��.�n��<��ɩ���òۈ˭����𛈝V�^�V{9|�N77h%.���+'7�mu�:_ZT��{ëދ��>��Ф@&y�ت�*��XWA�B[��
A'n'��MR4vW>��m%��K�r͙�ʻ�թ�յ�4D�_�[q�m��9,)i�̙u�o�uǮ`1np�6�t�u�p��yhF8�+62�P6%�s�V���aR��+=G�\vݑdҷ6���A�*���״��v4����q�����6�@�T�[M���5�ݱ74��tSrv�*w�����~�o�Z���o�bDt��ۏ���	����Ia��p�\RJ��A�����z�HL���ޢ����7�U��݃��F����HK^�E��ËRl��+����k�UhE���e��I|��_y�",�{����9P�d���{���W�h.�Vz{�:	�����d9�\u���k���]˭Z=h0r��)!1��pa:	8;;c��v�+=���a#�g����ە}�B�%2\���rH7�)>X��&e�,̩�O�OTy�D�;{��}�w��GQr�A�~L�n��;>=��
	�Ԓ�e�Bc�K:�+�y����a�!HO��n�Z[�F�~�h��w��ܰ�^M���Ӫ��r�V��/r���B�|PƘ{$.B�Hӓ;t����*��2�_o.�N���V�f���І�����2�m�J��Z�ž�E�ۚ����;��E�J��.D��z���pu$y�H�ݸ�3�AP<�o�G^��I�:�[���˚�P��P�DA�I�����:�m�6��G�X���1Po_`���WoטE��<>y��X�)��4��r�Y�������,�o���n&Pi$��o�T2��w�H��c8Sq[��L����"���[�q���k�A���=��t�(.�*Ĵ�������BQT�N��S�p��9���V��SkA���s�XƉ�[�g��H~k�ۓ�Zz��k��~�DPu��c��x(De)ݝC��Æd�������o��jd���Cٵu}�z�ʐ��*7���CR$�:Y���;����C��M���Hp��x����8��1��.�f�ѸD����خ�>w̭[X&Kh%��-GڍΞu=o��V�
���׈�)S���bWȷëV��㎼�g��%��d��Rj1>�$�IW�m#�������~�j���C���á9�*���n��g^������N�J�sr�Bf�ǋv]��Si�8�mBq'X��d�
����w_^V"�ͨ���)t�ɅtƱ��L|�gj���7�h�&��(�am'j���|`U�>�.�+�����Y9b��xv?F]��Gy��V��v��֕ԏyI�g�Xn+����ߟ7҂��`fJZ	J�uIX;+��v�-�1���+�;\�ckm��]v�]���Ԏi��K��+��d��g�2Ws�vTVÓV��
����oʃ5��G[��X�2���Ꮁ؄B�*��WV�@mK�*G��p�Z�<��ʳ�&�oz+%
F��iY�����9B��~u����Pv���I�de=�9r��83��c/N���7l��&X�黍h�.VկT;�-��sn��^�oX�恲W��}� �!%���(~-�ʿV<t�+� 8�օRe���	6zs��M�@Bo��om�d����Sz�\������g~��pU]�os<��O��A�I	ax�^�D]N�|vk*R匇����ΠaY��i����&7%���.C�_5��Qg�����O������ư໋'.q6�d���×}���sF#Ћ�B����M��|oW,�/
ԯF�*��7�����eJ���<���
�e^�B6������	$�*GW��q{����"�<���'�~�:7������s�J�#-nB�v�~y��%�?b̩��z��˔�9��8�r����r�+���f��Z/S�|������V5�0|*V����\�2%����܅,Zp^EF�U�,������[����s�RG��D_����f��vo\m��]W���]�Q�=�&�wr��X�w����Ro��7v'X���(����Q�M����*��ͲE�q�	�}�ef�F,���p6�?�����c��<{oUxS�[=1��ˬ�C�F;sjĆ�d�5���c��Lv�����*�Wk�GJw`.7wۏwU�!�p]����_n�\(������o���h��^r݌�Ӧ��m��^��,��c I�צ_;�Ǌ[�����1d�Ī�n�$T];:�Vt:����X���7�STU���X$���z�[�$mi/ha�wv��cw�{ښwy�]�8M�����L�Y;s������|�9��p��2,5wK�j���*[Io4�a΋[�tQ��^�H��Pc��Va�Xùp�i��}*m</�pb���3f}��
j�_`�/��l�3kQ���[�3x\��v��������MJ���8��i�r	2���9��كi�\��ov�;vD��ln5��e��g�ݲa���*+\��ghx��K�ܾ����� �pr�	˳�zM���s��9�n��z;LX�x9V�v��B�;Jn��Nً���&Χ`��&��v�a�#�����̈́9Sn���)'�\�uܤ�d���\O��Ӌ>`��S/`���{f��ѭ.�M����nޣ�+$��kpe���m4k�m��$b͂��A��$�@��y�y�sq� ��c)#�[�#�+9.�7[��ns��7<�쉥]��|�^[�-:�4�v[Ӷ�ż������K�&�A9��v�X��!��t��N
�9�#N�ǆ�v�Z��M��-۹Z��nȷm��΂�xy1��v��k���pn�9�{q�M�n҃u=�u��9�Lq��]v5=n�]<��ӻ��p=��p�frxWq���6�=��`;u���%�u���rv��n�������LU���۟6��ۭ�r��M%5��NܝG&�����::���ݖ���/�]7YKV����{%�lv�2�S{�V.�L�3���۶3٘�rvy������ާn�v朜�C���˂�Tl�ͥ=�w�x�b�m�ӫg����yܝy��왎Ex4Q�'am�ig�d�����<q�{m���
�lR� ��rlg�pN�:}Ү��Ǻ8��c�]��zNI;oH��±k�n����n(
�/k�呦��;v�ƜgY�mR�6�m�Y=(�v^�����ݻ'm�b|r=j���.�����v�`أ��n��,M���FNwbۢط��[g<����J�ݸ�j�o!��ݣ��e;1o�;2ݹ�kō1v��8���/ms��m����ۊ�ϳ�v��-�v@8���4X}���si���9th=���X����86��{Sm���l�o%[�Q�nw��t�6^�o(n�`���qCJi�[�l�g��c��labI�NL9U����Bە��l񝻎�lcfrN��ݟ]\s����N�8����h�2�%t9���h��t�j���^n�LpO]�}�0i5�5�����)n�y���mص�O;-6�\��݋q�p^�ػ�{�ִ�>Z%��Oj.��֧�\l����c�Ɲk18���g�N�3��5W����,�mW��5����t�A��NZz����V���1�ev�,M�S/Q�K/Y���	,7�������L��aP4�R��٩dR�O������јq��Y����G��~�w�A�z���]���Ưfp���ʼ&�4�WvD�_)$�h�7;ſ�U<%@��['m������3O�V���ަ߻P{�ԩ��󏹗|�A��6Ⓜ���Im����~64xj�^�y+�fy�:�RQ�5
=�޺jI�g��w���e��%s�t/�U��5+��3#���r6�tp.�=�<S@�	����/?of0/{�S�y���w��8�G�y����z��h���Vs�f��E[]�j�h��؄(d2��{�Lɢ�C��g:v��ѣ�|���|�8�YS�#���}�ѩަ]FN��q�
��}p&��<5�S#,i��(�QOg�r�}��z�u�v��me�u���UGlm���	&َH�f&�_D�sɃ���W�"9H����.��!y,��⨚N��^�|�Q�A��6��G��Zy=)sY��P"LJHt؟s�]S}��+�a�����`�����ɟ`�ͼ��;{J�L-�=^2����!�K��N�rÎr���/��Z�K.��LEƲ�N���>�7��n.�kY�����w?U��	���όC�Ab�,�}�d��m��ƓQ4͚����D �Ѵ7���x�-˼�|�IF��j�sw�a[{�G{W3ݨ2-cQJ)m�?Z�����@��ޜc�N�:��4z�>ĬPO25��R(%�3;X��kݶ���Z��z(�۶:��-bmDX���
�st�nJ�߭�<x�����=�|�N}�&Wr��p��݁ʅ�I��[�qy:���%�;���u�&�#�rv9�֭��a�]�eн��;��9�#v�6���"܏No3J�Sr��K"�/j�{:���y�[}`����}�b�q>��%f_)ٱq�V;�&܎Dڎ(�-���A
SڍOq�FۺY;6$e�����T�	�}6�)����[J�
�o��w�sj_�1�}*W���!D%ș-�����<0y�`��Mr	�{Ϙ����e},]u�A�F�����uy);=Y��[ޮAr�N�Z3g6�$,,:4_n\tj-�N���5J����j��+�|����F�1}�R�v1|}qy�o���g��DZ�O�%B*
XJ�q��u�5{�C�wG�y�Ss<|�X^`M�2gS��� Lo4�ޮ")�y��֌�z��7�{w_��S}/m�e��P8"5���]2�.�v,��x�W�\o�w�5J룖,ޝ�cW�����K�cW�c4�{}���,
2���l��c�i��b����4s>y�����ZݛS��FJ!�`K`�O�%�|��~�͟u�����M���rރ��9�t���g��+ʭ\ɕ���膃�tQ��
�tr���M��ș$�����Q[��[�j�}F�Џ��P�$�n�v�k���l���!����	v%�30�t��N��H^Y����܂]������t&�7��bD�-�h�+47�i�l���p�ׇ��a��>ս��މ��q�%b#��g޵*`w�1`����α`�!"1�t[������|���G5�U���~�-�wWK�ݯ��榨�у�_k��Y݋�ov�k�j
�o��]U��rޚQ��jX=�ЏكE�їcM��H���zX�� ����_�<��!���&��G-����Š�u^~fdp�&��ݯthd�9��̊��ؔ���Ĥ�	�bS�R{��ڒ槡�^=��Q���kU\�
w#���G}��Q�"��QRHo}���̿���CO	R��a��/WCL��1s����Q��;C����C(C�������=��b.l�"�0����i���?.�
��>�|��"�u���ܓ�=z�d�t���\P1�A�k��O]�}��ζ�d�������˘T�[%:�tM�4r���Jꟼ3�[ėy���|bx��歊Ցsfj�N��LBM2;�R��' @���<G2%�秬z�BM��7{�OƩ&ޮ�ȷ1��� !
���dEÆhʯtQ�yröz���x8���*a���v�6bI���a�C>:3{w�i;4��x���d�/{�ryZ�iiݎ�G������]�<z:��cZ�5#q8n}�(�ј��&!���*\�Ȩ���a>*oF��R7*i�kڌ�!�w�A���ѶPo��C!�ݛ6��a�V�x���w$mFq�l㝸�{Aӛ�8�3\se�C��2�9��-��w������rm��g��VumL܇`wm��myK�a�3֩�1�[P���� U��[Y�]��\�l@��N3����_6�t���c׭ﾾ�E�0�' �<ֻvXVv���T�WJ�m�WCC��v�g��#�x!�9,M�J!˫d�GΎT[�Iq[��V�#�X���i�s�x����Ӷ�g���D-�f�Ƙ`=��<i��:�+�F6�MGd��E���.����_�M����ן#�pos��p�i�Ԃ��9\6�<۽�A��	��	�"Z.J�,���Үy�����np�B�Ѩ�}�b���3R��mV�`7��F�:��\q�܁�o�gyb�z���&���rc�8aQaʭ����6PE�/[���¯K���U����W5�A��i�`�\��k֗*[^3��� @� e�c��ݣ~�eТb{j_N���J�7Q�}�3�+��G�dG��!���>N�V��;a�hzE'��#��
�;%\[��;ƍ�/������o`��^>�'Ľ�I���<��+�E|�g���[}�Y ���:�)�}��j��b b�jҝHݸ�*VYp��!.@
2��
����e��rG�!	aI6�`����f��D���_�ۅ_`�a�Z]��p��B���vZ!z5%Ō��$\q���ͯ#zmUs�n�eX�ܹ�q�Y|Q����\�����4t���=:�sib��ѫ[��e�>�2�_wM���W�jof�3��l�Û,#[F�����x�L�$�-Ȃ�s� �j�LX`���Z>��~#��=�8��|gS��P%��W��Ē�I�I�O�WK��}g'�������K�)���^�	�ܔ�'%�[Ǵ%���� ˪���O:�}�{�y�8�MD~2G�����3NmIht�r�t��L�!!*;��3��~-�ܪ��CP�k}2��x�^��#�ug�%c�I�0�rc*�F{�.����T<UswG_�u�k ����ژ}]א�TJ�wM�IxV�IYi�{�����������x��mq�H��!S�r�H�
�s���m�V�������Q�]6��"4!��JVzx�%<���ٝ<�
�V��ɼY��͕�ۿ��_g��2AG����P�4�P�4��kk^|�?zV1��$M��
�ԃ�d��[��LB�����-�����)�9�,��	zm�>��\[U��7�6)+��9*��sZ��S=�)*N̺%�wJ�]+�r�pwYA��M{f���a����Vu��57�Z�C_7��7U��T�r�`Y;M2���w3D�9[��G��T���݉��/\�W��h���+�I�G+����ρ�n#��<~²���(���^�3[�W��+��.���o���L���p8M�c7 ����ei0M9hE
rIZJ&l��Ws�i6�󠼻::��f�Yp��$=��j��=.�J�V�ECݰϾ�����|�~�F1�[Q�@X���lxt�qc����m�56n*�UGV����J�p��z�+�ט/5��$m��i�^���Ž�K>�Ϡ���gf�5n�"�]�=z4TA���=�)�ʮ_��}]o�Ϊ�~���E��Gw�Q]���+ck,w��t���ef*/�G�3�F�Dω,9%\�ya5���u;�����q�0�4?W�����F�t����Uw�]a�Y���n�$	1�>r6���ԩ)���`=�4c=^�nؽ�~^�^2n�c���q�R��;�Cwӈ�X�r�Vh6�w4ڥr�� ˽;܊=-f��������j6e��`Q#>v۵\6*ʏx��W������edH�-�ɊFYL�q�C��:��Q�k�6)�o�'^�٣�S-6����D��]�t����gs����q� ��(�mN��8��exH�n�����h̦v�hS��m��qF:l:��R���!L���}G���:+}���Jjs������h�����O�i�m�$�|��<�bQ�@p�������K�[h����]��2�L=���<��S�(v��b��R�؋�7��yx���C[* dA9$��-ﮪ�*��>���X�j���.�y/=�*�!����<o��o+��7S�*¢�,j�@�A�Ab�o�~�z�-����]��)'��ނ��HK	�t���r�I���n݃H�\�7}��\`�4�$�
9�?���U��G�lg��Ln���ݖ�5pNݲ�A+D[��#Ֆ3;ԮŊ&7�_�3I�х;(�=ћx��J�ĭ�əR��bq�g�|�]��q[�N����kFPOH��sMܝ��� �Z^�q�1�n��Y,t�@[v�h�H�^˪���-1�]��B�k���e�����NoN�Q�Ƥ(ːp�Ş��}���ȉ(��_[�]����r;v�� �un�.1�n���͉7�:�!g��0�<u9.v���F�swUP�=���v�`�Uї��l8��o:�U�{Zt�������0��F�dѝ;�8ˌF�oh��{�PYm��j���]�w�ĳӎ]̚s��Q�ٝ���{Q'>�k��e� RF�%C?˓!}?uҰJ��_����#�g��YR�\�S���e�C`Cz��gb�g>.�ת���4rl�%&�Qa7%R�8�;�u`�q`��3����Pr���!BN��b?"\���|�zj�)�1�����N��k��Q��$h�U����ߟ_`�QˏA��ҍw��b�K����{ޝ��e$�wAv�۔�|�n�Ɉb$)@��9`nb�onr�ﴏ;�*�A!���wAV8�官K<�U��D#_/:���J�{��Sm��*w�2�.2�4T�W7��-����I5��>1�8k�'�4�����:��0vW�X&�(���\�ꕳr�ꪀ�4�˳p+e1�5ݛ����z�������ڳۍ�U�3Gf�P�B	B�Q�Q0J�I|ǎwf�a��I�A�	�eu3ϣVގO�^��И�?k>o��-BoH��=�����	�-���BZ������N隊_C]Xn��K75`h%��e�u�D6�T96�}�oo.{ڨ�5��|ZU�%����]{2�6���m��6^�U���_ij �{�V�"���r�^�Esy�QiU��.9�0�O2$ �v�QmT�݇G��E�#�I�!� ����ܖ!�G�;$��Z��k�5��_����Ϧ/m�p�{wʟ������sv���,��Q�$v�����9�0T;}����OTu���/]<�t�R���N���[=A)�i�z����iٵ[(d{f�Ҳ1@O�d�ni)�}1}��Lc�T�AP;�ٛG�<�y��C/۴=Ҝ{���C�!�/yp^{��|�g�]~��ۖ2y�s�O���71Ã�t������ڛv�\���;�Z�h�wB�Ã��+L��k��M/z�z�IwO��]���Ք�T�}Ľ=�D�+�������ٴ|�/�,�VNK�'������E���Ň,v�L6c]='x�eA��v�ɐn����{[��KЃ@{p=�[�v��J"b0Rn)1����f����Ѵ�^}�	�����p���=��4$��Z�$�nu�ag:W���Ic���93ם+��uo<�k�7��R����^�䭐`x��J��n�el{ݲc9���}�J(��]mv�gN��\c�S���eV�v�u�2��zm���.�9:�ewR�;s.}����A��z�)�l{+v�YL�����ѫC�ݢM���9�4����j�8��F���nX6y��sLU=�&J��z�F��x����0މx]Z��.�<���Γj����\S���r=|����Lx{��s��ʴ�PJd�L�ʔ� 7@�(��m�nV�V;`�/f\�9�;��m�o)g���OƬ]�*��k�&4�'b�X3��"bCx����\y�L,�����R�9���b�A�7M�T��\�=�:�T���wX/ �DK��.`ȸ���6U��ô{q�/mH��f�ɭV���*��bӳ�(�^Ջ�-�!E-�1��ܫl��̿`�g������i�U�oZgmVM� Vݧ\��J��2��{��{Z�k�S�fQ�:}=�X�jɻ��0ѵ�5����BW��:����u�^�(p&s۠{FJ����7[���]Z�H22�hh��ǅ�������i�4��i�.� ��PnMf��ѻ�aT���Y��1��5m�k��Ub�(9v+�D��̀�����5��
[w$�eWV̾ξ�m]�'Vh�=k�.�; ��i���mLm��*Ν����,�YJ�.��ڲ"�*�XP���T_��
]��K t�_��j�m�����-���I�@��F�������n9�Ǆ��O�m�W���q�ίp�-Z��힔�������	G��D:ÚW��ĝ�rxn��&�까�
�.��m!d$���2������<Iп,�����qOgV��|�|���Ҭ�|�=]pz^F�l�>�]�Q�J�_F�� ����\Z���i4593kˎ���沓��$��h�l�		�'s��O�/zJzkB�.U��c�p�wzX�n�s�%��uT��=ͱr�|Z��(l�	]�Y�1+��{���'{Ҭl��}�l�s؆�'W�%2bҤ��b8�S<�ur��8�g�;�\^���E��Ɂ�+K!X�n��ˑ��<�-]�ee*�a����o�����Xo���!�򅁗,;Ƅ!��Y���RD�c&8[�H�8��Ϋ��iqDf�7�n[�W��z!
����{�!�	�h-��~��{6a�P��&f�)=h{t�)I��=���e���Cx��GI��a���sZYzf���GS��7;��b.��q�U	X5���o��!��g5���R�F�� �Ebw=B�d�}l�Ե(�Ϯh�T��s�{bM!�
;|�x���4�+_f���/W4_d��Ʒdn�[$mU0����3�GAl�Om�rqmZ̝�l%�-mr���퇞������@8��w��.o���yn頥�*�*� �׷�`��lsҬ�����=��>��T)��~���ǠQ��7$���W{s>�y��Po��Ude̾�<�͙F
PIܙ��1i���m��V���]���LNCY�l��BLQBNAd[O6��l�.�ʙ]y%�\Wr����F�x��4�1:÷PE|��c-���\-�P"I 46ߩЇt�B��Uu]�VM�op{�!�\��V<�&;��*��yW;�p��[���O��2vy���#�
%(�����+���E�uEG��#[N빻$��zC����;)܏E��O�ݛ=�j�Z#F_=#���搕����b��⵹��c�7�;�+;0iR�trˬҞ�#aa0xQ�M�u'A)��N2<i;N�Vʎ��	u���f�f���;��wܧd�J�ܗ�\pJ�
��t^�sk�m�L��������7u=��	���S��L�x6���\�����rpT��G	�;���rg��yx0c*o��O֭�B�ћ�k���ۇֶ�m���v#s���:�� �nm8�l���aŬ69ls���c��m���h��xP��Ӟu�`��0x�ٴK7�kk���[�{�L�Inި88�u���*;[g�\m�׶�㒺$�b��v��5�Rm93��]������i��*�%�����%*�9]����۾�m@���.y�{�(5oz�g(���281W��f��Wxf
0��f�}��an�5ʼ������)K�n]wS�Q�KVn�f�^W�|�;�g��2�G̻��5��O<�5a�QrM	�r�bMr���`�Ϟ���8I4E���u��"�[�z(Ҳ�\[��%�rD�]S0ή��M^�P�����S���m܌���_C��	�r�˫(���r�^L@c��Vhg|�	d)�	��m�<Uo�����=#�s��GnF�R�#{��EmW�y�f*.�]��u��3Hgg�HjdX��Y�S����C�o]0n]n�=\�R\�Z�;!ٳ�Y7^�^qt'nA�g��F�+]���㐭�u��'(�\{�D�ۜ��M��e�)�K_�,���	YOk`�Ĺ�"�%H'$�Y�w����1�d��t߫
҉i:y�6��D+�uⷥwm�:�iF!p+�-������� 4�L+*��$�ᴧ���7H�O�)�7W��pW]Y9g��:��$0���.na}��2}n�����xAvx@ߦT�wdմ�J(���^����*�.O[�YD���*�z^��K{�����t/��JtX6Ŝ�p�0�/��Å7����1X�}(��}����l�M3=}0Xv��]_k���PKN�L��	����f�nE�;)�
���,�M	N0�F'_�$��fof�ލ!�B{��w��yᠶmѧY�619��{���T�N���_ m�|�7���M��r��+Q����C���%[��q��2���M�c�[d:4��Z�=B�d�%)�/�2��r�ίt�^��󸈭]F��e��A-����
�V�nHO�;���
��ۦ5��Z���BC&�s�"���W^���Q���O2�׳�#�5�?hq=X}s�<�?��I�ià7��Ԋ�����(��I~��H�n�ߺ]IM�*���=�8����Dm|q��sM`�c�B��o	�u֋�P�w��8k���ạCt�-��oݻֶ�p,VT<㻇n�R�Vg����2�dg�$�U���bF�.H){�O}��64b����:ޮ���i9��S<+q7N�椨��1�7gNRd)	D8��#�QV��^�],��d5X5��7K�$��8�!��K�C�6����P�
<�6}�3�©�?�*�D�MES�RNu��(��vw-�3���b���S�����4k�ͤAƤ��������Q��^�'{K���W�./M�]��#L�7��T�����6��<���(c�C"�Ie�m!Yr�8����nI�����b�ȑ�Cݻ�G9��[~�^+t�F+9�UPݭ���\x�!RDdD���od��,�Vl��.w֪��$OR3�̺�VJŵ'�]������!s���7F?�R h�����I<�*:�,B�CH�o���r���\���h5��
E+w��g�s���4�*���ʨ��4|E�`�Z:f��5�nV�攦kr��rܫ�ϠCV���T�.V@o��^�)U��m^�^�U�+�K�R�a� RIv�\ں���ݵ#~2m��̙��w�R
�� (V	���:���� �ه| 1#�������N;f����ln�՗W�p��K�גq�;p�k�6���ǎN�<�#D���X}�_e[5��Ws7y'�u��X�6��4���?H$E8D�.����<�J��+�>��ϑ-������_/,C���mS��>�x\��v�k�,cg�<��C�^�^n�若Y�M��Y�8�zq�_���2T
8A_$��)	�c�p�)�N"�#��R���#u����<'�6�����ǵ��]�luz��uW�U�tX�$ف��L8��ԡ�����x�u�ݎx��)z\�~iQ��4|+/��EIX�/~��G�x��ӷB+loGo���}�K���}2��T-������A�[|u�-��Lm]�}IpY4��5��{]{� z��T�;C����:�<�.o_K�r�n�YX�i���<?{�ޚ�����3	/tK1~�9Μ��-�v����4ooeK�Y1[��Eh��1��K� �FR۶����.@ݒ�h�û3n{q�n�Y�"���Ի�v��^͎+��gṅ#]n|f9˟X��ᄸ;��[���Obܾ0Y��Gi�۶���[u�Ӎ�q�iݻ��թ�;tk����(�,a<��8�v�ڥ��&�Ur�n�/����伃;cqPe�qh�3�[t9�7P9��9iώ^�)�\k����۷�O}�sα�Ľ��q��TTܺ籬8;s�V�m���y��:�p\ ������ԏX�cq�Yu[����p^�3h}�t�T��l׷���H5��	Ñ�E��
�i��z��o�zz)�F�Q���uG�30^�Т;�c]B{>�`g���L� �y�
�Tz�z�ߔ�S���ؓN^��F�9䞶#1&�@ܗ�iַ:�V���YaO!~wݾ�Ы��EG�O.����U����YEa�It��'����%8~i�%�\�a�-B���߷:��7d�lwW�9�҃���}1ݎ��E۞���v�9u��fס�Bu�Kls�q�I�"G �q쁳��P4�w�/My,��N���ld�'��Wtڝ,Z��Cy���)�T�MP9W{�P7�����v�EC�q�b��B�W��I����t����<Y�\�8۵+v5m�������׎Fs��k,+�xU���}�Ap�!��{��oe^�=����5
�]4��?*�\q�Iн��p0�a�`$$�^��0��"�_W%X߈!ۺ����A�גf]��T�o�
���4�,����z�fF�d䙱��F�'3~E�{-[�f<�r��)}[3��}�J�P�ǩO���/�s����צZxV�,��S��z�τΜ+rڏĶ��ݤ��_ЀT3��S�����]�}U�rz�{�ۙ�i��gC��P쩔00U�-���c:�C9�jS\H�|TJ�I���'Ƴ?
7�U��\7�7��D��%��b�M�&�oGi,�F:���ν������������엌)>��Q��$vnL��z]�Lvt����s�K����O��'B��ڞ�'�
��[a�9�;�̋���V(�4	ΦZ�\f�p=�u���#��va�ga�� ����kvDi4p[f��~������1��k�H�7�yY�&���MI�J�������[ނ�B�������,u�Z}{!!I
�l��9y�Y����dt6�Y8a�3��q��s�L���D��!۷Z<���A�gW$�nU������U��)Ym��X��AW���gZ�fmP�����w�&�J�V9���U�Y]\9P.��b:u����%�^���yZ��v�N@�ͺ��e��i�Z�&_!���t�yb�a�go��'v��]T7�P���nò�}�Xj!�����J���7�v��]$t�~�!R2�j >{�|q��4a�{M9<r�L_#^	
>=ػ�^��V���1�J8���RS�t�q�U�R�J��勫����t8ҾʩY��#�}j������%�g{\��]�y�m>��D��-H���&�i>�k�%�b:f �*\�Ѵs81�J��F�Ҷ�J<*��y�Y����P�f6�O&j�N�+����gH4nOW�lu~R���{̓n�R�b&�q�9�f�sȵ���˽fr�(r����=�9uۤ�d�/5$Y����Vm�3�b�d��ia{<��~08��\0z�C���0�L>F��V��-ǉc.�5�}���>��l�\�����H]E% rJ�Jq֫4��~'y����&d�D�g�Y�ͪ��z��dRx����lB��Y��[��ƚ�O�(�i휱ob^��=�x?�'`�f���a|G�R�0r�=�f��@��x�d,���=���;/5�#}�}�ϛ�g�&�����	��η�v��.�j����.y���Lp;Vp��W^��[�"�-���<�|l]�����hHÀ����x�f�r�Ŕ�����6�lv��t��eON�%����w��dX<]�R�@6X�L���>���N�dzK�����Ņ�-��J^<�#��I���d��qÙ}*[����kq녻ۿe�9GFk�HݠaP�'*�4A�y�8��qoz	ceo_z�jmlMqy�L�6\*D� ��9��'L�����F���U�yhg=��^а�U��׮�Y�^���c
���Og�浱�����mN�����h���C9^�]����)W��j�a:�[KnN]�u��h&]����>��5Agt��;��n�����ʩ	�7�Q�1��b(�!�୪�^�2Mw,X���)t���W��9Kٽ�1v@��}�}l�_:]��k���˜=U��ݝ��j��1owf���8dm[���2��K�ue-:�����w�i��y�ּ�J�p,p�<�fT`n��M��=���k���ל��d٠Q���Z���pl�]N�\f������svN�rF7d�Vz\2v�k��bKw���ɵ��٣���{����z��^!�A�%h(8�!b�y���k�)W{�^S�� z�Vg�����p6�k�3+����_�'eMN�:�w^�vy,��2H,~�?u��c��)�U���/uu�(�j���K�
=I郯��ɪ�k(��Nf-���cEH2Sx����������;D���3kk*����+�����+k���o��{��l��%�z67��*G�#�Y��l�e*����^��R>�QJ�1XNr��p�{NS�\��Zy5W˪�{�>:pj�,vGݮޣ\��"�:�k��fx��_4�ռ���r)�Y][�mmAgwy|�|���ol
t9�o6η�"���H�k�}u$��Q�������#U�f[��{�3d(m��fg^� ^B��+?��{�qC��)]sUmc����6L\^ͱ�ֽ�������t]R+Ek�3��aMt�O�ï|f���'�;�yZJF�ƶX[}���&&�8��4�]CCM[Qf����GFo&^�G�k
�krV�mn>��:uh�&�ۀvB�i��Y�>��[�6�4F�(�e6������s{V������A��m��%��W�3mꪩV�CjN�U6�ے�j��|��t��M'^�Ǵ�d��=��=qöWy�t���b���b�V'D4�SV���i���j�����}=��]��L�mk� �]���O<\Ar�W<�ûJ���r��� ԭ�6�me2��֍�i��1b�\�[I�������xm�x���]va�u�6ۜrU�u˩�y�۟e��G��P�/�-�n���ՇF�6�Hsl��3���������ltxR��Ƿn�:N�lb9W6!��5�ۮs��B]v��KV�;hw��F��M������];��\�l�q�u�[K6ツB�OI�Kӯfn���n<��j7�6dC
홮��x�箥	�N[=��]ƁÚp9���D��k�7-�0j�r��m@��vrueN�ss�sN7>`��=��q�c���se��ҮQ҃���=ϷI�q�8�7��n8��V����w��W����v� h��}�]�s����v��@gnu�n��m٠�Uۖ8���B^�ۜ����OT�E�z���^r�]����p��p��ַ1mu�[qL�wj^�պGv��=71��"�i5����3�������I��u��̣��l��C�a^'��N�e��6�tsF&��v��sΩWe}�6��u&��m���av����Վ7(�Qn��ظ'���u��Zd�xK	�g�=�a��/[M"N�(On��8�޾�}���8��{Z�w:�؅�ѫiĶ�6�;�zz�f���O���[�\<�;�S	>i�R٨zݛ�X�շSyۓ[���ﮍ�|�<[^��r���Ŧv5��+fVv��m�,l��'��hS�΁!��v�ﾻ#��v�%,ۨ�������ι�1��qې���C�A4�nTSjK���ɺ�s���7�9�su�u��5��ǡ�^ښ����[t�P�Z�`6�`9���c�yЃ��m٧nܒ��;3�Ӱ�͎���$�UEwc��ۤ�ݭs�nSc
&;=G���r\7;{Ӗ!�ʾ�tqu��[ǧ��-��eMU���v�^�<I78[�����04Ga�ڛb�]�-ۋ�c��͢�wQ�g��ط`d�1�-�[(��nx�]�d�%7j�0�u�s��KN�mV�cK� �n哈S�u��y<�{<�u���M�l]c��e���O�ų[��[�1�a��-є�|�����%�ͧ��R�ӯS��^�Vw�}�:e7]�kF���҉i�1�1��
�����߫���'T��d��R�"�훚�!��t<~��d���U�����;���9c���[������6"e�~M�1�gѲ�spBt)'�z�,��ޝ�9p{*�&��>-e����W�,��~�u����`�5X�+�B�G�m�F�g<�L�R�S�^'�V���|΍����	����cn�[W�e��(�����(I�� ����a����Q��;��*��Z���k����7>�T�G�5׻�f�sc��
r�������q<�F�G����\��yzC����b�����+��e�n�Eqq��}.�0����Ed�)j��>��p���^��o
'��q�˫�e�k�jLO)�<�k��Y�ӝ���xے��ŵ�o�<���M�33\N%=��q]�4�G�v�c!���dn���i�S5��2q��:iÌ�}��]�pz[���L�G�p�Lm�M)����:X>�캖xƁ���벗��9�3=�|_h�k��d���N���RF��l{qT5���HzY��72�a^��&�����RQo%�{��c�b����j�M,I�vf�̵Uo�`BUڴh4���W�n¸�-��V�i�9w�[���׎��U(L��9lS�M���]�~cD{t���"ǈB	bFJ���á�(��y�Ə���>
ӎ�c��Pp�ՙ䵷��|I���֙;%�˧��xEnH;��W2��j�t�tWX0��VOW������r$%�Q� �j-v��/�"e�V{>՞��u{�&�3\L���!VQ�P!3�g��&4�ך��M犱�6�֢nܳ���ԣ��z.4�m�<��� GEe�ݺM��#�&��~[�c�������a%z�[�^L^�&�)���_�3c�4�}^���І�����l�b
7(���-u��#7���i��L��2�A�E15�_T}�r�w�h+�:뱛����#�0P*1�8��]�$iȑH56n�X��b��=��G���U���.v,�ᆼ��t�K��G=ǂh5��.��{�f$o�9S/%�CaY�hM�$\�I"͵^�n�*��ĳw�;}]�Ͻ���/�Ꙋ�w�N���М�K/h� �"�S%Q�ٴ�s�� �;ו��zఆ�^tZ��'�P{x�kc�R��H�v��ڬ��[��m�^�K�/��u}�[��QwϮ���eX8�Z_jf�{<�䕻ܝ�ux�r���%�ˮ���/��ܽ�_Cg@���ڙ��I��[6,!�v��-d��ZW�yk���{�z��ś[�$�B�NR�-���.�A�Ml����v�t�����h�ߓ��[�ۓ%˭c��"�,F[$�e�¶���>�y��~�Oh�
���*�������+��}�����}&�v��8���zڞ��9+��9���l.�
�G�޳�`�~1�ay�v���R�������x=⯔y����ՇWAM���EF]$�P��>�4�����[���*X�rCN�]�z��{�*��vG��x�lT��ٹ�{�g�FT��}�3���ºg�Y�$E4�� ���>�;CZ:�N.�p�^@�/��*���A�V)?w��y��v�~}ߡ@��r��
�qF�-)�)I��h^N��Gm��X�s�tv�����WEoh�`�y-2���+ˈ��R���ޟrl���ql���G(W
J��6I�`��'����n�f[�s���ۇ]E]Eb%3�iEsy'rv-j	J��ǻk;ޥ/�'��&^�D�g�w�����isf�!J��aڦem8����2H���2s�B�W�0ec.�����,X53�B,����ʮ�d������pņ��h��Hhg�H��A#MB�rL�-D��Ur��Ϩ�L�Ʊ�xQ�Շ�O
�b�^�w59��4N�E��^ȷwЎ3�
@g�OM�>;"�E��8J��싻a�L��8�4�ZQz���x�h��g)W��ݽ���-/F��}����j�/_ggVM!�O_��l�l�; Ee��{g��&;���+�]��|�%�����E$`ǫ�^b}��gK�t6��j����Y{5Y�l�n��ݻ�6���C9��66<�]Bs���-��Ùyg�"����}�6�N��sf�m�H�0}� �܀����8خ��ۧ�3�vloV-p�'y1a�q�A9m�lFn�6k�hm�|��8ۦ���K�;d!:b���s��8� g��	BJ.�]�lĞ*��L�n��ƫ]Зu�q�ã8l��r�p�=���a)��lc=����������:�v��^��e�q�Rm&�:㞚s�p���c����y<Y�G�u����\�\{��.��l����'k�6���ؕ�g�[p���]zZ�������G�O��ut��<�H����Y�ӇJMQ>�����DRGC���b2���R�P�}z�X�V������ZIj�������k�UN�虤�S��+�ά��KU=��T�-^�4��e*�Z��C�]���[�ȸ��tl�����Y��W%	bVgJ�<�����g���f\b��1��mB��)�C�޺a�ćSu��M��ݛ��}�3w����U�+����i6F�K�Շ�޷2?UĹ���B�	�B(�ynEf�OY���k�}.:��y0w���{�_*${fZur�*��nW�3��x���B�7���x��)?���FQ�FԒJ��CD)�F�ծ���nm=���7a.}]�-n����WG�~or�L*�WЂ��f��cT5��z�2V[�����O'�m�)���r��YnH�Jہʸ�dq�W�;P���/�벍0YZfV��\��T�s1�䧔��F�˱Q4�T����tѣ뭇�n�+8���Ҵ٢��+}�V5�)���5F5��]^&z?g�3g-i\s�&�_#D�_�g�VFq:�S�OԠ%L����y�y ��5��8k�B*u�'B��x��DE�Ҩ6�;��ˏ�/.��}���îCu�,MӴ fzxS޷�\��=�>���.�GGn�ν�N�r�\�:�U�پn�eŤ��t�N�HMy[ـ��f�t�B+������3���Ǟ\����{�u��5��!ؘQ\W��0K����wI&\�h�Ⱥ^�V]]��T��'l�eZ��x��^������^��f)p��r�c���Md
^ۀ�zF��k-��h�2Dd��(8��;j��vP�k�dH�S�t�ݎ��Z�i����$@r&$�0��$�v�e&Z��W���^�vG���r�#���+���]��luJ�����Ɛ��u��⢕J(�eg{��uה�<ߤŭŖ�X�w��;��f�&�x������w���r�s�@/��U���Vm��C�4� �0$��F�Y�B� �o�x�(;������i��C���2*�E�#���T=Ԫ�֍��-ۗ5����#I����e;Vn��ӯ��X
��?��e�4+�&�M6ǒ�'�ap7Vײ�;�REE�!Y��l�=�H��}m����0���Eq'&��X��|�
ڣήݘ)
W�w��{�`����_`9�j8
���(�X��n�,\Ȩ�/����e��m�3��Ҿ��]��+%9e  �v�em�׫�v��"��u����f�i�]�b\�l¬Y��7#��o���nŷ|��j"^�)��/�,�ݻp�v���[����A���۱uv��ɞ�S������U֙>��z,�0��Ay}��[uG������=��yB�yZi�%�2�Ga8��Ы����b����/>I�z��_@*��3����O,���:�m`ŝ���Y���-Dן_+�l��R�*��r\������?@KH�NI�>��|o�@ߵI�x�����b���̔q�a�5*B�-{��5{�-��R7�D�e�Z"�����A�)���槡����O�]�M�~~u�{��P�n�;�{2�&�:�ԽV�b3�T����N�w+S��'Y�ےDs~���ק=`�rlts�cs)��4,4��y�K�u}��d9�,:�*�Ǯ��JW��,O$&��J�a�;�v�{��ف�ʒA����3����z(@��U��ۏ���.��w����P�\�2w�^� ��wD`+Gq�o����+(���D	�$��\C]#t8����F:8J��\\�nK�(ѳ��5)b�e�1�,�M5�9_���/��8�y�[�A�aRDuy�����s�)�e�����et9��/c|6�Gn�#���#���q���Hro��
��!wX�lp����Wp��R����װ`���2�*��K�V�[��o5LP��yaD�
�j��FT22KI�ie�h�Ӿ�J�u�2���dnF�����l��rW��JB7�ɵ;�J�"D��݋�ц	�6������MM8͇>�C"�������<�OR���͙�]sݮ����9�w�^���7���Ǜ�¶�Z^HK�s�#F�(F\qKƙa�F����y��$9Ԭ��]���_�|)a����E)s�Ӫ>�.�p�"��4ZGj��b'=�M`��׭w[^Ŕ�#s]´a�A�8�]�7f<�ُ3�1��<ۡ�*.��Mo-[I����=8���;�,E ��S���vl�����3�fͰ+�Ӄ=�jk�M�l(�ӽ���X�ӹ�)�n�qn��E�]̀Wn��#��,��БGZ�m\��v�j����}8�^�T��n��Um�댓�{[���s�.�ٶ�����l���ɚ�a����^��x����=vn�j���q�"��IIN�z��I�S�]��gD@�ח�[��\.��x�3��uڞ�uو1[t�3h}KtZrs�6�V;s���"�@��q%$�����,�w���2/�"c8��Ïh��16Nr�5���rټu�d��?��w��G^R�Ɉ�I���' ϗ��CLo�[�E�V򫗓�Oz����^$�]ʁ�U<������u�v%��U/8��zoe���O�PT�;e{ƺ���]Q��R�Y&ZU!{��^'ٛ~�P]܏|��X�(5S[�����l��(��K)�m�;0�(�}���<_�-��I^�x�A��U�����?V;8P�d͞���O����:Ä�W|�u�ÌC#1\*d��������qV���Y���nk>8��B�voI���2�Rb�V�`y�I�E0���uR��G����?�ݾ߳�t<���Z}�o6�D�;ewn�z������]����Z�8��"9|��Xg��Y%������<c�J���Wr5����[�D���l��+b���Q�S~΂��XAK�~�˾��-_�B`2�4Nu�Vf�@�Ujq]���f���6=�XѶ=Z����ʺ�}A��yT��ESF�9��z��WF����:�4�F*fb@�RZ��U���u޽�l�]D�qNFGs.��[5����^g"[B/B����;۾�sܩ'��;�<\>����&R���aI�8/��zU��>2�L���f֍�~���+��bS����o�cohc����@��Ӫ��������ڷF�yߢ#�:�*�G�@ț�I0�z)J��x`���J̯�QKg}�H�D}���~P6b˾μ.�����_Qs��?3)`Dg��Y8�y���aUl�-�U�(HA8ADF�w{���D�U�����5b��d�WE�n�S�]���j��K�s�ާ����&Z��e�=�	�B?�VƄ��c?a���౎-v�y	��I���y�zլpխ�E��ke�U��n/'j݅��txѲy]�,��{r~^8���ӫ��Hv�\��vP(U~��uFʞ�����"Z~M/��{�=��Q���J�g(۲�$B�R��q���{B��z�yҾ�A��u���?QR#ޞ�8x�ϕ���j|\iz���+�v|<�KVT>������s�s�A�of�En��Ɗ�&
$H�rg�Ú������X���Y�*�����;��+"�}f�ܷVU����^����n����S�c��%Q4�kk�k�b�4�W|�IW���90>g:�Fw[t2�RuYU�t~Ռ���z�|�K�.����X��V-���� }���P���=$Lv�ݭH�H���) F����hm�˷��v�	�T#n��6S�@褳��:�� �GǷu�b@sUf��1�a:����G>����/����A���µ����v[xFGlV�����SֵZ����me�<�&�ݬ&V�b����r�j���g\~�"�{��ܩ)f��Wp�1e_<�m�q;���U�X�Z�s�D�e����:ʙ��R��Bcu[��h��"�/�z�!MjC6eHn��dZk(��ƹ�{<n4�)��4�q���^�:����C���e�2ܰFL��%+I���f�*�Y/�8#u�ݼ�$����]��p�e����ma��[kQ+!�#T�Tc2��.��=Sw/qcg3�|uvgowp���¯`���b���o�����|����sPɝ��qnC��J�R-��R��v
��Ն�(����h`�T[��{�X�Vl5�ˍ������Zo�� mM�X�٥(-��i�E!�7���W+yy�������8�$ڧ/­	�ŰĴ�n�'ďU�2YpP0�9��_��L��oW=�s*P���JWi�\�P��<��=O2U�2��3�V�ݪ	aҖ����}�����:�խ������C�^�탅�A>9�)WR!�GI�+h�Y��}Q���9'���-މX�e��s��U�4�I"t�4��b����1�����|�L�����><g��~�$���_O�!h�>�y�����6kS���Ĉ���_{���F�B�DW ��b�P���C��#�"�dv1�S��v�rD b%��c��� a�����^�iPf�S��^CA�M�~��fo�U`�H{�}2P1�ȏ����~5Qd@��B(��\�C�������PY�N#�?���LO�za#��&�۟�NQT!�Ndv;b/4 �v�o\�t��[�\�X�k�\rm(���U`�)<������7�}+�q�?���{^q��c�Scg�Q1�7/�W�3}����A��t�R:{5L܊���XՉr+us�le�̦T�)˪��8�	����WƬOg�_/_��<>�@:��/��i7��@3g�~���K_@�w����֊,�1}�Į�B��~e��/P����}�Z�G�Pkz�(��"3�q�_;��
"��|��Z���7{>W�ґh�"�r��9�$�X�wu����;��G��K/�g�_ÁDD��LIO�N�*k����SMC6	ffw1P)
M��	��̳�j�h�z2���fN�������f�q�.�KJ,UW��iO;=��1/�IT@fe|\,�Ĉ!�Z�[գ�K�̞����X�����̒�7�֔��˖��8�;�w��|�=ҍ5{������geK���+�Pz숎���n�y�y���m�>,��D� 9�{�,!�A�2D�}�|�H|�� /v��fθ�aA릝��3Wۙ�k��!Dv\�V4���ZK褎c�E�\��9Ŋ��0�(��5.·[c;̜u{��$獭CϮF,�S�V}P�3]����(�PVB�h�©[\����A3�Mc1t�3��S��A4#�|-�R�^4�ڔOۼ�lvs���_]�21�d®��Ϝ�w�����	����0�%WzP�b�N��Ϻ��F�_���@�-IN��Օ	��3�}D��>���`󳺉�?
xX�>�~��t ٌ��D?|!@{�Uq�dm��\��˯�θL���K\95�G��#���^��f9B8�
9�Id ;P����mq�B��k�E�G*�+�Eg�W6��@Bۃ6�3H:��Cm}��F���T�R%�N�ƕ�~�iQ������1}�@2(���OY7��G��(���9	`�C!�y�_=�S$��>%Dt�����V���P��eܥb��ܴ���դ�$��GJ>��?��� ��s��dq��y;r��}�R���c 1P�Eϯ�����!�*f��"�#�j4M	P�HN���Z�� N�] ~N�ê����`��6~D�#���:��:�-C� ���I�>�w�}d8����A#��o>�WM-�X5ndpPV���k�1��3+��;qY�J�6�Z�2Qؕ�:�JC~�y{}� ��u�՝�T�IM60�W�";����Z�uj[cN���
Pb:z�r��-�_g���m�|���sl���i��k�S���1'/
��O�C��w !q�l��X	�n
�'�,����U*��9+v"�R4����]v�2��l.�ax�n�Of�<�.����:�5�]//J�M4���rgu�3�p�m�	`���u�m�n{Go8��<�_f�u��{</p�ۮ�n3��۷��t)�s#�2#v�g�g�uv+�q��]	خ�d2e�h��r̆H�L7�D��@�� (���u�"0U�;~�D|��L�"i���kz�χ�?/&@<��[ ���c�c�y�������a��qF	�9�ZT.�k����~!��LY����M��d��P�j��%*+P~��yW��ȍ.��U�S���M}�(�#LIkYS}r� ��>�!5�8��7gh��tU�B�4TA���~欎+ipP?.�x^���o;�!2/�}��9���NdTUQ7
��� "�ԑҫ��ZX��K�MʹiP�A���������o]PU�6��x�����݂��!" ��:VP��ϡ�N̡�h\㌧b�(K1�K�p���L�ML8�JI@Y��!�:��|�������x셗�3V$��p�%�fvcD��B�o�W�>��m-,J�q_M�אJzD����qv_V�>���|ϣc'�����O�?߼��;lV��G(�lK_l�P�s�`c�	;�����p�ɆQWN"��7��j2��_;JN��*�
�+��긎�F�o�x����!d43:gha�~������ N��Z3��~�Ø�e��g�v)x�.=t�t���=��y�n�՛�ًd��iN�!)ֻ5�;߭�̗KPЖ	}w��7	i�v.BbX*!P��*����h�Ɉ��	�%^��:�_�Ǎw�6��ڒJE|�Bϝ �QU��q^+��8SѨ	#��,����x�@ϣ8cqP�YGC*D��d.�zP�G	v�tM3�~�qa�X����];�z��}ً1^37jH���;o�`ʻ�T{��ԢF��g+�[4EG��Y�
�M(֬�{�_o��7�J�
�̜V�%�-��p��O*U��iih�D��*]F�!Dr̶�">Y?{�_	T����DQX+#��Qw����l%���S����(p��7�,=�>dYW���q$k��.4�p����;��gp�g:��ߚ��#I� ��#�F��Z� vz� Y��bs�<�
�_2'*)�O��ᝃ�B��hռk���JDH��\�[��ZE��J�;�ن�iQ�!H�������e���B�Y�y��zoK �6S_}�z*O2�	��#�wE|1 �5Ə�3{\P��4�����I�0��Y������n�l��H)K���>��}{ȥ}�U��5�EW&!����r��Պ��XaQ��D2��*,\�o��	2�N"H���R%�Mϳ�Uaś�~%R°i�Kk���	��;Oe�����\�:����QO ݓ��	���F�*Zp֐��ݖ ���|��ʞV�IEG)���v�,��F����&s�x�66�?zȫ�0�����d+���;o-:Ԇ8��R�#�d�8-;���_H�h�LT�R_�E�c����Ϋ ������-¢�'�J�{z�oH�jR8�u�>rZ��V$#x��I�Of~��<�<G����
Ӻ���#�C�����,���!��!��a��ċMΧu�>�Z	`����$ި��7[���`����ݹ��]v�F��.�u嵆-$��6L1���+on��_A��ب+�[~b�Ř�Ų?Fo�͓�������^$��ύ�Wq��C繵(l^�cN�`��o���b�FB%�~�(�yS��2X"�d�$ ���ա-;�zY
�w�7�څm�T@�Eg�U����4ȳC��F�<l��>�U�Dh�a����#hݥ�F�`���U��~��j��	�C����dd�L���sψZ(�U8��Ő>�W��ե��g�
�����[�ඝ����? �%9���ƾP,0����Q]��7b����&��G��E�α����c��hʒ�W����;j-�CnU.�h�*@�\�S]aƛ�v�8�y������ %���t|Y�}� �!d2O��{�ƽc͑13tW��n�R���a��ԦB�d
"W������?o���#�2��i�II&b\�+�8N\ՆT,v϶���7�xKqT�|�ͦE���L�<.��>@~��b�:�_�@�u�
���8�����!v�:�gzv$��y��(�m��1��Q��,�8���d~��}�N�~�C��f�������%|ǀ� JÙ�^��~񳣚>��}�R�� !���3���{_s��C���0 #�|�#-U�!��a[�8�|,���l��P���>�@>�oe���7֕���|Ⱥ_}�+��=��:�1n��	"=t/.���N���LD��;�s"[�k�B��S��e���As1��cq����2�ꃳ	}��lN���cZQ�p����Q�ˁ��K�!�or��X}�b����zᮿYF�n�B�s���O���)��j��K(�Rت���}�a���g.#1��Q��De*�5����~6�?~�)
Fm��l��{�4���}9C�\Q[U'��K#�	�F�R�Ɉ(dT-�C�oY�@���sq��^9��s�3��<�߰,��]ޟ
��"V`�G$GG���@;N����#1Xď��E��\s �97�&�a��@�X�E(�nՊIkCMz����A!�r��J�US1D�+���!\�,�O��X���+������g�^ί�]z�)|�Q�RP����� V~��!�|a_]��i�{w{�͜}鶻�B���y
���D�:G�a�[Z������t�� m ���P�J}7�W�"�=a�?qk8����B\;;|-[.p��Y�qBb}j� %:�1�g�#1Y��Cg� �����4�E9%6x�<I��]�d��1~_Y{��2�{�}�7��u�<�ULo/%ޫ_[����U�1�L�Ǫ�ۦ�7PeVܿ���G�����]������wpQ�y� �Cݘ��6dp0bQ�/ﰌ?=]K�" ��S����$'����V�iU��6��Q*k��q�¢Www��We�*���S~�e��D>�}	��kO7�<���o y4`U��a]�_k�y��vi��'�C�@�A׷�.t��e�{VN9���˲&n�lQ|��e���~�_�xm"�"�p[��g/JMۧ��p��l"��u/�s�ֻ�G^M�8����,f���;tg��E�;Y�%��r��z-�	g�]���݁�}��x��ɣ��΃��9��p�X�'k.��u����ɹ�n��vC��u�B��$������ݲ�p��v9�N|�8�3�3�ut5�� ]��A��l.6�L]�i�vp�Nط[�[y��\eݴ	�e��Y�7]��cq��ίrv�t��R1c7S�ûQ]��;�m����'����w�<{���ٕd�V��Vڂ�}U˼��Xh����v�}O�c�J��',���T��6�О�������B$���D++�1�m�$w�نc��Q�N�WeRJ��X^����,�:��;� K��j��AH��Gw�)W�n��
iƊ��(K�݁�{���V�>��޻����dI���p<���'LIB�uU�,ְ�G���0�;�!��G��i�Yl��L�[e�*ۓ6��){���65H��$x��m�@��
�!�>D4�h=��b��2sz��g-21�I�����u��Y)���l�{��������������1�==\kᘅ�!H}
#y��V~��|���v�W�)����P@z�����*�}�{{!��?�t� :��Z=x�"Jq��̷f!�����'��D�����^P�ę}�����k��ץ�g�j��!ݕ
3,����if4��T��j�F��2�|��`�3�7����lύB^1	"���v8��t�m�L�ʽ�b�m5�l=���ꕎǵ��x�?���߽���|{�"ZHV��3=G��`}1U���jgԒ%[�`߭��������s��qV���=�:"����_�T�>��3��
p �=�&Jm�jI`^/��/����#M��ʆ���I��2��s��-�@��Y���o�K�73 8�dY����Knx�꼒�������to���8i�*�{ V+�����XQW��=WE�Ĺ�c�$ @w���w�@�ޟ*TG�*Л~�_9R|��@2��O*�4��]A�D<@�+��7ն�Y�40�Nj��.���sl��}�32S!m�}.�b{�d�W���0�;��x+���ME�� �p�=Ѝ�&��W�0����O��|������i�l|K ��}�0���D[B8�!�B�+g��*�ȷ�a��0$oR�H�$i�d�ib-ن��vLu o��J�,
���(��ӯxe,:-���&��!����G匄T��2@��t:FP���{�w���a#���ejQ�%��	�l���]��~�/����'d��]UaQ���?f?�$/�l]���SZ���7�l2,m�+#��ۍ�\��	��\g�E��c��W�[���.�-á$�ԓ~�_3�aa���~�f^�E5��xF��9��{M}·g�~^�*!f�i�v_�wn�Ǥ؍JB���D$~��Mh�_>��Dn��W]X��LQ���|�Sr�]%�"�lĻ���7��_'�WL47�}yg�{����� �9'�Fv�p��w{�%��D@�}N�%���Ԕ�8�A�D�*�#��d�@V����ĺ[�4Y����_��τR&�h��b\�i���ϋ��+����
�~�[a�� ���^���M�*wO�����S5�-?��M��ip��W�_�,;�W[�/��JF�UrB�׳ٔf��Ί	=��-;����	aa�[(q�o&�G��e��W�*���mz/X��p�A�]0��h?E}�2�#�y}�[�3[�A� �kI&LJ2#8�E������Ŭn-�C*�N����Y�>�˧ @�I��0����ʸh|�|$@i�}"��s�#�Bx�F��y��c�XT�,�ٌiD��x/��P��0���b��D
��	�C��v�=������e�fU�<��ӑX[GXW^�L��1QH����:�
���!�?*_D�m+�xY*��v��@�zF�~�����=�Qu�{$*�~�X�G�Gm��ɹ�1��:�N��1�:ͭs��^9l��٠��H��G�<��> U/��w��P���uB�&�|��{�W�� ST(�R�b*��[�kw�����H��T��{��~�����!���SD1�H�&R1Ã<�`6_O�4�7K�z(o�����ھ�)\���䆪f1�"�d'�E���S�z���dD�X��49���ܬ[:߉AJ���_B?����@�d
܀�j�������ހfhc;}���Kt�&�j�7^�NyU|�OϺG�S^��$0�Wb��0Z���V� ��_Q^uR�7�y�PȂ$�8�8��SR`�p�H%�o{�T���FNh�����G�e�C��@��"�Ŝ�(������F|v�,o��{�Ưo(+2P�z%;.�5�N�����٥�ˣ���	��4j9v���mz����ÚJ���a�J|�׳�_��k���R�2�Ͼ��8�j$����~��U�,�~�����5��@I���u7A��f���&�d]��o�U&մ/�~��}7�҂�� �i��r赳7snN�pf]�N�v��q����ť�>.N�ò�͹
��a�ϵqg���vz�wl��u�kR��v�������/�)�h��k��|�`"O?�@��(`���T���wk�IW|�����ĖWr��;���	��^�Fb�.Ъ�+P�/k�-��1�HYw �B���*]�K���@deיּ�A�\_z�
���#d`�RH���7�����-D����^����!�k���۩�/�F�|p/d*�&H��Q�3�mL�.�_t~��!7�钒oFZ��"�k�j��\���#c��ސ��
#k�}2%��<������g��d�V�yCJ�=�F��E�;F�h��싽ԤQ2�ޒUϊ޺�͌���P2g�O�c�U;���B\mD�E��;!>~_78�Y��
��,��[�]�S.�gv=(LMw{Ůٵ���(I(���	(I(����IBIDD�$�$�"��$�"?�	BIDD�IBIDD҄�$�"?�	BIDD�$�$�"?�BP�Q�	(I(���	(I(���%	%�%	%�	(I(���P�Q�$�$�"?�IBIDD�IBIDDP������T%	%��������e5�]H��?uU� ?�s2}p#A�'JZc�J����5*��4c�� �Wwr��
ڀ�j��8T��ڰ�$B��ʺ9��h��Fځ%�EڊJ���T *�E@P(��!RQ*�@�)D�%B� 	 �@��T�@UP�P�H ���
J���(� �JR���a��Q�t�[+7�:�[M��x�4�\�������N:$������qv�O\����{w��p�޷{}ڽ����EWwL�s"���(r�@�H/=��m�{��P�J&� � �v;2��Aɪ��;7Kea���m��UR.�(��J�s�$�ns�HEWu��*�>�"Q S�(*�Q�� U�Un�
4��ve����Wa�E�a�ͺ
bΐ	�0�;�A�@�--b77@�N� &�m�cq�ن�� J�z�t�����W�`�E�%e�MEJ�u΢U�ۜ9P���8�E�D�������� V��5��{�碂�8��֋ѐ/� ���*�� 
�O���N����P;��,�y��4<Z�p��
����@ 
y@� S�e 8��(���hz���%�A@�u���� �<�)�F� H���R�� >���@�hhk�w}UJU�hP�z�t(P^` �� <@
3�Q��]  ���)JU�B� ͅ�t ���=���j�� �${��  ���T� (�H�JT�U�t��e�T�biD�g��Q�1��]�JR�-����B��K�b���J#[;t��p�kl�v:�5��� IB��Tq)���r�4nDPs�������n��]o0����`�M�	9P�u��\�	U's8�\��LJP�� z�H�P��)RQER7))�&�%u��6ѝ�*T�9�A�w��&�
st�X <��k/�绮�i���>��lRY�"�������ty=7w��"$�v��� Q�ۭ� 㺩N
 ���aл {��k4:���G!��۔|����y�*�]j�[jyZ����w-��R�O6��{a��^��Д�T�!2�J@ h"�dĔ�(�  E?&&�T�e!�F@jy�A5)P  �*U4eC�  ��JT�h`x��������%�����U7�����	��7���_33j{����Dd�r�H��Q�#z�ڹ_�""D(��Q�BQ��""D(�����Q�#����
"�!(��!��I���Cc�h�彍~��Y1e��;-wJcB��&�*cx�)�eÚj�!�Z�sw"��zV�h�VHѴŪ�H���f��݅�Ձ�|��8��f�.g\�f!���m$�f�4�����Z(�dԼ�k��bd3�]�
'UJ�X�l���ܺ�3X��R�r�˗^<�]���\W{j��Ez^�{�w/0�� F䌪C,jz�-o��c7n��
�C��WV���cxq	(?�-nhّ�ěT��P�L�j��$'$�[��%��΍\���В���C>��r�b�;�u3�+6��-����J�z�P@*0�)s�x�74-�7
��&إ��~�c
K�RRYj���+�i��O�Jj���IZ��v s5t�re<^F����n��\X�^4u�1S�V�C.�S�К�/%�pG��3�v��Ҍm��D�L9*��0"64������W��s�^;�Q]��ԛ�����������;
��칯� ����� ��p����&�q��{
��p�@�u���nL���SEѬ��]St�'(�FC�*+5�"���P����oU�V�nv:��6�+��I�E���t�m�}pQ,�mJA���¥�TTZ�{�-��"��7�k G�å`��Ǭ^�J��hb6�
WM�:@ʆ4eD�#���&nV<��Pt����9��D�^�ͧ�� - ���*CoU��:�T��M�r�r�bf�����KP�x7�M��EDb!�J�	�ܶK�ՉG#���t:�,�mG'�؇���ã��-��5��.�d�(r���E�I�G��I�%�M��.��A��ݘ�k���rh��ngS�m(86h�dYD�*�R�9��c�."�RX�4�
��5��E]���儞a�G^�9�(���&��f=�-̚��]'�f�7gxiwv�w\+����j.ur���!�T��,��r�i�� K�`$��Fm���aY h�Mz��	�*,(r,��J��8Ӭe&V��o^[�e�x(6�1�	���[��:����k֡td�(m��q��@sTŮ�i0lw��[[@���*��ޑ�g��7wZ���B��$�+A�:Z��܅�ƹ�'V%IR��e�U0�R�U�
i��N�v=�����S��$W:HǏ:��(d�H�6DW�d��r��<Z��ur�����뭹����[͘����Y�'%Q�G�[RI=B��s�����߸N��ìm���Ar�fjSs��Աt'aa��zY��5z�jުp�%��c�&�جF�VNZ<D<���	nP�y��^�)2#E�O�xܣ^������ޕ��+F֨��֐�7{c�f�"�kpVL�73u�@����r-�߲�j�����8���2e�x�O����F�q��a��U[��w����%�b�Ղ�̹j�Y�ʗ%�ҵ�{d��+ EEP.�v�aa��&˅��)(�؝wbQP���
�Z{2�Ȱ�ʰ����lY��{�(�Tf�O@�\�W���G��BeH�*ɦ�ɱ�시Qq��O�����<n���ȿ��wh!4,;g���f�3��n�`��V�K���ͼ��Q	��XՒj���NT���|�_�u�U[VFe;�L���a�/w�.���tY¤8i$�G1�h��I=�n1���7ʶ���:N�{��m=��u?����V9��T㳵�^ꚫC��� ���� s̺���<�Ȉ���,�� ���h�U[�����}Mí�����͎��n%O� w �f��w�c�;��M�ء	��6a�݅��%�Zr؇*e�Q��t-�
w1<1��EmШ�fp�x2�X����jF�w��Xg�4���݁7ic�e"ή��F�[��Y���,_ֶ%{�,<�mX�çD'��Ⱥ���F^�*�In9{���B-��6�a�yZ)��5�[uwm�YS �	*}���Ѡ4�V�v�i����k,! X�+����/	Ȓr�N8�+J���d����[���Zk\V����n�-9f#�pe!ѯ+yN�F��2���Y���=j	ҥc^y�s�F^-��+¢�1Z)*��L�F�aUk=s��Pk@�A�Z͛�wmI���n9����-�SnaB��5*9x��Һ���-���&�-\�Zb�3�	Uh����)����!֩�.1�'KA�:�QaGMȈ�޽݇FE�J��4����t�~%ש=Q�J�&�p�t�MP� 3���9�k.��Sr�qY�g0��(��
�m�[����fR:�M�]���SҴ�˾G�:��r�ҳ��]&NG��*,H�d.��9f�T�����(rl�gMފc]I3s]{��-|S���pG6�P���5"��^�[E���m^	�J�����jn-.a�, ���6��r��ۏ*�<��ٶ!�/Fb��5s$X0�I��E�A�/�;��V���6�SV�`�������S�5C�1�� L����y5ۗ�7LR�0^�љ-j�B�W@�R4�^j���ܙs'��̋��p�D�A����^�5j)�T��+/ ʚh�Z)�N��-ɐn���q�:V��aې�T˂��y�3��.�5�ve)v�e���r�h���ΚV��fӷ�^�iN��Kh���fs�Vf�����&geJ+u�r�K�C� �䅕���aC�J�oW�QYz��/=w/u�m�%����n����F��������l�4�	7*׎�Y.�]㷲���yŜ�N�4��xϜԛ�6�t�\�X�VP�a�:����\��19��|���Omlp�k�b='3)i�r��������K�-���.�+m��bs�Y�<w���(ll�kM$��W��F|.Ǆ��������f6f�2�uf�ѡ�[���f���v�t�FI�k-�ڞ���Q��ta�;�\��p�9���`H+�iݝcMٳ+u9���9¥��x���}�J�{h��j�d��e5t�:#�J�%��r[H�`��وa� ����S�ɛ��LFX��wMk`�aU��ժ4���Ż�<���qʞ�SnL3I���ZJ�)e�u4A��l\&�cy2���<N��l��@����+ܫ5�1�qթ�g%ٺӸ�m��*޷�����ӌ_��js���r���Ϋv�B���v�w�����w��8�ۼ�ުp�.CX�c?�gՆ�A��-��A��"]�+�Kb 1�%�#�ݧ��d Yե3���`�\�/�aZ�c�r���]!.9s,�p�5ڳ�C�V�}]8�R��{*��)w��x��MP�^�,1B�֘Ek\2�I�K3j���
P����U�&)J�֕u
���c��]*\H�n���<��gh������-:ϸf�JO�v�������V�|Z(�X�WF�wR���.�!.��=}(��M9�֧�Q#j�h:�V�����3KC�*�|j�uS�E����+��*��p�zIKyJ��(/���6�>Q�.�|�d���.M0�彬ܚ=b�}�*�ܨO۰c�`ײHț�������1鵮����C&��i��f�*�+�y�	�:5e���w:�5|`����/0���ֹU��"zm*��>��j0����r�|�I��}��$����e㮢��n3b�WґB�4��,���H"o��pZ6�t���Q��w
T������"���	�&�Gq���GYN/c��å�BXFĬ�H�@���\���׍l���l�id�zɺ�YY�&��fQ��9s�~.�o<�Jn(@%��ڤ!���em!t��O@�X��f���b�^��,�j�� ��R`k�Z�嬳F��`����-�4�'ُM��I4�h�A�"�س�],ZM]4A��wh'Q�	&{��αG6[]ǖ���@�j��1�Am9Zyv�#�e\��!�9 aY��t�@�Zf��N\B:������J�O�Np�66D\'n�LM�n�t�5�����R����BACu�vIk�6�3k�n���0�?I�%\�Yc7�I��3�u�oD���ς�+,4�)�~���"�ԌZQ̕'ڮ=��B��&�-fr�$�݄,��K���I���i�3��H8��-�;�ܜ&�}��^��t%c90v����T@2�a�Y�8n��Ů�������Q�S��ڻ��m�&`T�elc�)f 5�{`��s*�Nm�kj�9��-�4�0U�q� $�dr�a�v=y6C�8��@a�wi�MT��&H��^�t��Z�� �D��W�|4k�DŇ�)# ���:����*�0=Z:[%)���YD3*�LB*�L�<iSDr�M|(�Ǜ�$&)��BH��-���^�C,F���cNV�Jnhg�"���s2�t��Hҥ,�tl[�fS�	��&dm��#B�*��cwzq���H-�S#�Gcd�:Jʵ`�a�y7��4��s��ZG����j������	V�QRi��m]?��WeEҜB�)��j�C � ���[2 PD�a�d�̄\b�sA̩56���G8�f�6IF��T�u���QײM�_*ywj�H���V9@�e8�[i�MK&5����C49L<��2Q9��ɶ��%	%]�P=���1��RͣsE�0 ���
Fr�T慰ջ�2f��c�B�����)R�[�-���#C�M	<�x�CXe3%�5n���&��M�n�����M�m�2mh��ܯ/=�Z���i�\=$�r@=1i�dlH�HCĠrC�M�$N��z؆���S�,����N��m�2ù�No�ͥ���$��bko��Do#�tt7%� W���h#�Km��fH��]���dܺ���R�b�!�4ōї��2]7�Y-ŨL��\��L�r�V��ܸ�7��ޖ0��­���%��&��]h�����W#����h�љ-|
��hմ>M��[ �#�zT��H�Z�䳹b����Yp�-9e�SNc��(O�{�I�6�����%�![7����
͇�G i|��WR۽�l;�J��\�� �D���.i��slj�R3y-^��T6 ���|���]Ymwa2z�O)��X:�2�0��H WN�E��{ݡ�m������v>V���c#�x�ˆ0kk4(�W��5ޣ �WRa�hh��	����V!^]�J�����V�V����Ml�1X8H$&��F�9��q9�ݐӓp�;{��0p�H6��º���U{\�-�c�s�,O�����I�:��{�j�e]�:l�sB�гK!�vI�Q��:n�(�Vw��t�+Q�͍�2	�K���ӽ9�v��;����9,����h��z���9.�$�4x��{,u��ܺ�R����	�ODJ�1V��31�*UZH�}IQy�r �������j;fn�����58s5��P2i��2r�"�@��xoL�M�j�JC,!�ybŻ�[� 
�R��ѵ;���xkv6)O�D��ֽ�^'�,?1�e��CE�RY,"K>b-]Z�E�w�J�Ms+jԚ�lC�
��v��v�P'��,a²V)r��P	ψ�/�RU�J���K����8~En�E�3y���w^��ɛ�d��Ѝ0�t_��4魞�@a0Y��L�LARp�TZ7��VF �vs���B��w#�l����3J�]�	wv�*�&���$��Z����:�q�ӏ&�p�p��}��FFd��"�7��9����;X��m\��S�U�sg�*��a6���Mc��Ƥ|�m��v�6.ڔnh���J�l�"��U]դJ���lfS2�w]�ˀG[Κ4�h��1#K����!VJ�?�]=��Ք��VS��/
��ţ!8�P�E-��bS���r��oIYGo�F�����R6~;X�05�֤�ڷV+e2n��%h��}B��F��ZQ�aq)��R������[c˦��6SG1<�7��KCV=h���� l8�Y�(5�]w�=��Ov˸8C��7h�_8�*�E;��2nj�yt�����lL�e���*r��Mۈ-���\��d�ĵ���AV����[����{��=V�I!o)���71J���6���Z1W�<vBM�m�+�`��c+���L�[43u�{i��� 46��c-�Hjşl�Ri�CU�4*<���(�V�f��r�B�I[�{�a~���#<Yͫ�1E��Vk"C�@�ώ�4J��!�,���KJA�1��� �9��B�Zݻ���tS��`�k*�Ĕ }��$�Q���6P�D&��6�k ����C�.#Hv����f��&Ωf�ʸ��p憨Ck�B�H�xG��niؕ�!oS.��A��T�be�t,l�FU�ȓVX�F?Z9�2ń�mͮ���M���t�n]V�x�9V�8�c��3vu���0���3P��^��~63�6�1�&�
orm[7UvUu����5ۀ���2��`8Z�\�B��cv�[Bh��dC�0(�m�%�/^+�M�!c��I��pt�K�� xƼ��K�PLyW{���[�!v��2�,�ƌMؙ�dS�L��	��K�D�	5�ܣQ���.)�v��5BF{gѨ;^A�:��r�c}8�`v�]��c��?yv׸�L{[�-u�e	�@s.��1�A�y��a�_�mW�ʣ�=w�un�	�]K==z��[��d3���L��ܮTj�6ҵm�˖X��bꣵ� �����AP�m�-(0S�����겪�h�g��l\����d���Wi��Anp�Ի�wV�u��\�ng��hY�KX�f.mb�X�Q۫��:�5qKѼ��=]���E��%��=�s-��3��R{un^a��������ЁN�6�Fmlu�^[t���a�p��w���q�i�{W�������c�6;,X秨����d�·�o��ɲ�D1�����og���C{ue8��>㍝\��pm=��s��ݑ��M�`�W�^3��Z'\}�5y���!*�M�z9��F5����8�2Ss����nܽ�]d�C(9[Y-%��٬1��T��,#���ci���,`�3����[r7VKk�2�v��&�Gg�n��]m±�Ψw�.�[]�,?�u��J��0aTm dV���m�z�g�\��ݲV�=���eyOj֍���Uĸ<ϫCڌ#!t�����A���"�i9�붓v��\�`�7Dv�C;O���6��N����J�[���Ⱥώ]ӷn��n�e9�Ť��7V���wd�[��.�����}[׭q��4���h�oM���N����8�4h��52��5e�Ł��SNq�Dl��L3p���F�e�G[p�޳u�:�����`�uIaL�b�ٲ�!�n���Y77IkH���hKlYŮΕհv�+�� ��cv�ݕ���)��������:�!���]5���4
*�g��Ϭ˕�5v��q�Ewa�x�cpL�K��)�ǋ��/9���dG��̴��u�k�;nd�%��gK��x�t��I�;tg�P���W�I�r�����^�Ep]�hn�睼m.�l�X1��պ/-#	�\h�j��}%�p���;<�j�tqo��+������m'OUӔ�z�$�Ӡ��z�)$����v{l���cB�%�^�:t�M�F����1�<.L�s�����C��@�]����V�α���!�Pp�iv�B\ZR<�x����8m+��)�ִ�{f��6��lu���ke�av�eہX�.l�(��n��gM�%�xu�n�k:!�E��&�����l���Ş��J��{��/�'nrN��&�r����[&L��s�;����P�]+H�4I,!q�i��h-�*�g��]�1V����@n�tq׋q��z��ns.Px,���ֶ���W%�&Pf���5��g+���]�#N��n���Qwvt�����%�ak���ka��f��1u۾�z뮞�[�>� n�s��s=�ے,Eeѐ�m�ܲ���P���{q�U��ªp�s��//g�u{t$[\�p����E(�4�ux �w��2��ڸ��t%��˦�,�x���a�t�m����ٍ�u�Yl6�fգ�%��ff���mE�P�J���4���mm�(�^h"�f1�u����۝-���Rs�ShR�Lm�NK���2�Ы2���M�l9�>3{]�2\���WmF�v0�̤�$�6�t�@���Rr�9wu���ێ����x�7N���b���v�ԕ[�Z�Ce��qm���S�:ۇ�'.v]`����\�!�r)��j�Љ��v��O �t�����u�Q{3-�*2�cz�ӭ/���wWj��{[^ў�6y2g�
'n��J�"㰧e�U����捓�|@�%�3�=@�6e�S*R		��6�+�fع��S�f��tM��B��	M�4hl�HM�	D���,Ճ3��8-�����+���C�r�I���(���<�j�fH�����3u�pl��R��=����͚�nq��u�
Q���<����4�h�]̻b2�u�t�z���1�t�p��� �-&�;`�p%ٶ�!���B�r����jL�Ԯ�c��71�V�r��E3uV6�\�ye�h�6P��`9�]�볹^א�K`��c�A��[m�κ6��m�IfX[`�K,��]P�	fl).�(З7���=�n1��7��h��i��݊��
���L�:� ���WX��2಑#++�3�K(ѦV7l��.c�V���ͷ�Ge$���z��.�0cX[WA5�t�e�V-�S�"a�:3si��1��ۇ�'����\q�m<�<���s�']}��	�y�Clu�Ujqg�<^3�&�e�s����8b�����ɘ���j��k.�m�4Z��sK��b+q�c�r�<{=��ɢ�����kb�M�F��:w�Cz�j�g�g<�<��.�=.�rg��380Y�lsr9�m���l��<��u�t���m�D\��/-��>=\3&�E׫P!��3"�F��7ny{"r�|;d����=��-�V�󝺽k�Z�/�a˚�5x�J�g��Dn{t��_KE8Wb�t�Cv�cN��{f�a�]��6.�w\��U�G�W�B�5�z16�ZyE���c�a� sȲ��9lE��f���t�Ө��)wKv��w�V�up����w��a�5Og�r����U�����]4X�ĺu�iq�#gR{Ko\��'{��[�v���Gm:.�%�ݟk���丹-�vݭS��,�PAy�m��� S���.;a��]^�-��[a�eL2饉���M�kǘc.�%5�������p���K�����V��p�9��c6 ��]���s�������:%{�][v�q������84��.�,9��Cs�x�-�k�4#�v:�6�����8�)��=�&�\c��:|�G��؄��12�\�b��4
���%�l\;�<���B�2f��\g^ֳ�U�筎b��s�u�=��D�e�;p�=��e�F;;�F,vқ!pcD�v$. ��Uں�[!۟<l96z�y��cy$�y�����l��[N�g�6���R6��p��V�O[Y�;I��պU:E��97'Y�;q�:�qu��çy�ޘf!2�˝�0�M©6�F�p@����t�V:V<cZ�t�T�#�\�׋(��Q�nxL������\��pn�u����ٸ�W�/8ʘ��\����Oe�suۧ��V�7kcT��m��2dS�����M�5��5���dԾUx�n.�f���ZF�1��:]�c6İZH��XMb��o�쾬�ϴ������1+��c���v��3��S�oe�lv���nF���\cn|��Ɇ��ѻ5	�� ��s�����Nà�)�n^o˂���`r�%k13�1�T���9Ґ��-VŚ�	�&��Ш�bqq�k����J��pu�{:Dcq�l=��vڗ��� A:f��S�6����gKh�Ӭ�]��9���g�.2�,��6θ��g����Gq�5�<�y�ģj&�&�`f�JۀE��FT=�h�q=��[���+*7Q�$-���T�;XKH��-�Gi.!�2b�q�΀gv7n6��x �L�46��Ί�u�*]�.%[�+��z�R�չY�ョr/6���o=�No����n��-��\,�"�귀�8���7m���Қ��N.#���q3<������7��;ng��ȻDY��I�ㇷra�u�@-���v������>����-�Vl]�7)\����N����Y��b�CGj×Y����ی�I�D�tc[W���a��<c����9�9�v^���>�s��c����m$Ʌہ�⸸��ι�-�f��F�{ջ3Y�y�1�oG���'���l�o۞�mu��7X�Ez� c>��m������u��V<4�K6�-�q�{a�`)�nݰF
+����YrA���3f��8��t�c铇A'6�K��Hm�bҴ.DXTgVlյS�Kf�K{u; �=�r�6��N�2G]�;ո졓z���N�����e�W��l��љ�
̣Zq�`��=T�q�_\�׾`8��%�[wgq�E�p��"��꒮v���3%�����Ʈgb�#����G��EW�`;�ѹ::q��s�yn���<cV[0�)�ٍ�t&�B�����:�u=<�^C:wa������=v�t��Vհ�\��v|RG��F�8Iu��Z��F�F����ԏJ�Un�4�9H�g3i1fme��
�r��/4����[�<�gS.����t��N܌d��P�t$��-x���CV:}�㱛�ù�9��k���bT�A.�2R�����#SV�(Jkp�6 ��>� 0�)�=�z�$����ʯ=��]�x�LR{!��8�Y��!��%][s�W�Cq�NWfx�w��.�P����.��sm���<Y���:�no0/�<4���ݗ�N�\�F	w�wI�����-�ܝm������&�4(Ǳ���<�!����n.�<Y�"��CQ�NU+j\��*��.FBJ�V��u�k�͢?�1�ۅ>��K�t�N�8cF�y+z!����N]�	cr����d1Z6��̈́�yEsp��]���v�0uN�+�܁��܅��]�� ��૎��nr���V!mJ�-�����O3i�׷K�F�rt
��҆Aj-[e�2̂nnֳ&�u�Xf7���9�36�g�\��n޴!u	��P;I\��mڼ3�m�-�\�����Fy^���77�ݼe3���OW�pG�]�G��GY]�I��W�������C��]�$.��:絿i�P��_]���8
5q5&�t1�fhA�o]t��4�]y�s�
$څK;9��pc��1N�;ƇPolF������C����ɼ�V�k�N�F�bG��݋�kk��,c��1s�4	ue`����w[d���31=T ��YNrŸ�$������ƪ�\����0��.�v�y�Od�
E��Bkm�e��3n�ldbF���-ti7F�ˮ��D���42�;��k�,�K�R2��}�rv��[xn���D�ÚU�![����[��b:-�[t�T�")P��(�J!(�_��S
#�Q
"!(��1�!DA
"b%������r9t<�8vZ�"���	YYm-n��\KÃ�E���6�����JE�\�����s�0�AM��A�U�\���,c���9=�͔U�@j�Z��Ps���VVe���,jJ�
�FӲ�ϝŴ�c�I+�Nع_��eM\Ş�<z��^9�ػm2ɕ����ͣL�� ���[��Jr��'f�m�rk��4���-�]�/N�X�E�n�a��RN���q�؇;��4XG����.��.!�K�B�i��'�V��z:Lлm��%���CG.]Uz��7\��D�O�Q	�;�Wc[��	�C��ҴI��q��ۚv]s�\��� p���n\�֣�Z�n8��9�4j���{�v�6��9�=�����E\��:$�{L�X�XpM�b�"v7��U\����W7h�xA�d��#�n�w3�)�/'u���X-�C@�%se0��)� u��.�����!u>Nj}�>u��;R�n�G<�V�Z3��cstܲ-�I��4�+���P��1�rsKFFA�cl�=k�V�:$j�:�Ђ L��İ#��Lhdn��̖���2.�/hܜ>N���E�]9�����=RM�u;5X�Cce!�#EY���wn�r��>�xܡ��78�����]��r"[p;78v����Gj�ԅ�T�0 �#�׎�,�nS���%�� ���5���fi�9�K4AF�P44&%��)x��s�eOcN���)ͺź,��q�R]2�m2ޛ�a����{q�uB����6�B�,�6�ƙ�6U�u�xnC]��7�@���	�A���5�&tK��KS	�v�fz��u�fN���L��h(jB�A��5�-����VGen�Ÿ�QO�ݝ�s���)��n$M<@�8w�����^;v;O���s��4\�s�+�sr�۩"�0a�������%�Yy�l����='1L]���3�<�M�[��u�oz���#���툯���w{���� � ��P�@(P�(P�P�$�P	B���$��A�$��P	B�������Q
"!B	B�m���P���V'-�ˬ�15���m'm�Ӽ<\s�`nC�v.�8��V�Z�l�(BkrR餭��l�0�X�8q�����vy,�;�� G�1���7E��װ�����5bѲgEt'����V�-�R��$m��:͗ld-�0�c��W;i#�{o&�KT�6���E�-�CZsEyіg6�k������W%/M@�<=�u�'7G7'>��d�r���*=��?6���X��w��"Q1a�%���?���@T�
�����;�&����w��U�c���u�����<m�%;���8o9j��Ӽ����ô�
굮��x0&Np]Y���Z�F�oF���&����T�x�vf����5P_b��r�L��n���+��-v��M�h/.r^��Y4��D񷊤b6����0��e.����A"pv�I*9��V�}���~���k���ë3r����)�dt���@Vo6����,�V6 	m�.�%�Z�$��~���:���}��G,��7�b�fjS{rWm��ew C0���]���<���ڨw]�*��6 zQx�suO-2$,�!�	eh8�uY��쭚P��#+vHvf�&N.C���%�WX��j)�F��~��6϶��t7�]�aP>LV�,����y�I�ŁX&�4Hj���'x�z�0��]x��?\�\Q\y��37'��֫���(��L�t֑�:�A��ç�<��u�=����tG
m��M�/��R�����������i��ͫ�x�t���d��:Åԫ`%E�c��R��k��&6�X1�e�0q{�e(k�2g�}盠,��dZ����gs�����G�{���_�OVUW���-�=LȠ�r�iꝁ��6���wpF����9�	���aH��f)�7��=����:�W��G,T�l��)�U�2}u�^�!�԰GE4s�ر�L����W��c*'ܻ﹑:��֗�ܭ�cv���v�m�yK<�$�z�ք[ݧ�ћá��C໕�J���7���g�ځ�1
�<���^�;h� ����62���3�w=���x��z�;�<m��os��C�)�u��^޼�t~V�z�T��	q�1)VNP�;Y}ո�Oir���m7���0�b%��a$��IrC�ե|j���~ڼ���Sx`^���˃8m+�C�~^��dA��ڲ��A�J�����X�3S��[Öѽ�oib`�q� 2(�K3��w��Ĝ��Գ�Қ��o0��ŉB�X�&��*u�VT���CC�QE�3�׈��R�l���e�{j�����u��0V��P�"ך�e]���]������]�h��Ӂ|U��NpfS�H���V���$y~���e)"���q�JFs�M���o(Ϭ���w[1<�֙��N� ��O��d�<�b뮌�Z��o�V�y��kÖ1N�8r�8ʅI#y���B����fK��c���I-ּ ��9�qv��)��=�z�ѷ7�	Q��X�ZiJ7�tUS����K������lr-Р�czY�g[v��mq�(]��ٕR�Xe^2��s��H ��T*=�m���>x���n���˥�
M�zAt��E��+�=��O�z�yg���{%)rDP	��!k����Yw-�,�0{=��^�K2��}��ezՀ*7y�Y��I�Z�]W�x����Iޞ��H�-�G��U�;�\�����+�u����R�j�kV^h�]�5�{+�W����t��L��H�,�$���.X���QG�Bx;�b�5v`�F-�N�]B�+�_Y~�R�v�1�:���Y�!Ί`��*F�:`;�!��娇�_7>�{m��������i.�xo=3:b�h X�K������84Rt�^e@$�D�I!��eS������Е�+�V;�	�_W��IȞkŚ[��+��6����>߲F�Sb�J��<1�Z>!���Ɉ�q���v�z��4]����Ǭ[�m�&����%5�&D��"Z%n!a�gǺ}�y�~v<�<L�z.�����8�%�.��7k�5����G����_g�C�s�}��u�5s3v1gK,O57���WvQ�o���!����QF=;�|�nڭʙ��tÙ*��Y�M��B|ː�7�i�%�58�;V�i�$��ﵿS���#��T��>*ِB�9oe�g=�,�E�mK�@`p����Js�6�^�D�y���:F���C��r�J������9RA��%V�pO�����+t��n?hp�?)�z��e�n(�l(܎6�e����ٛ���}�������ys��Y����1s7�y�wH�mou��&خNLfM5޴��.������Y�'�-e��M�Y�Ω�m��o�]�u��[�'5�r���ɕu�yCQ��uYF�c9��	8��3a�XK��5��v���Z�	�����p�۝<fwns��v�����ximޔ�L�w�ðaۍ�#��f2���IE��5�Y���ԄX�Yn��e�
�.��Ү�i�b�ù�0�]�d��h����n9ے{%�x�r��7�l����n3ಪ�rU�_k�/1́p��lFT���V��Jd1�63h�!��Q���'��o���!l�	��c��j��M�厁b��A���]�`[���V֚�e0�a7�$�����?�ʲ���@�]�+�1Gz{��C����כ��G�C��G���C����+��؍�Ć{J5��(]W.U�6���>y�R�r:�Z���j���~�ʒ�=զ�êp�P9�0"/v�I�D������@�M=Iz{`t3lӔ��QE�A��O+��q6�y��.��lٛ�׷����Ұ��#�]�q�E6�4�,I��%+Wyʼ��x<�I�+{�Ƌ��P��,��SX̗V��u�$y�f�P<��[M�κ�~밢͘L00ϻ�i"S�����E(fmx������C�U�}&KY�[�q�`�ӡ{U	f�7��6V֝�)� �U�`�6	ŏ88x)��ܔ���:��6�W�W��������QB�-DG28�n�=ۛ��`줍��|�6��^h3�c�I� ��W��ƺ���)z�j�M�шAJzl�i�Ppf[��_1���矟Xz��L�����]�����
�h���u�R����4�e��X	�8k���ӬJt����3�W4a"u�_K+_%Vc7��l=�
iY����J�����ʇ��Ʀ]��*
(G�PW�	�UV�)rGs�
�1��X�Ű:�M^�j^VI8D)'�:�O*�ikįP�f�֣��sz�����:�ߪ�Yp=��}�d>�xM��.�����Mq1[���P�� �܂�"2o���N���ӻ�;��k̣p�N�q�`T>9����T�k)tJ�nW��fWz"B	�u�}��x��:�����z���m���Қ;	i`�i5�	0�ԩXT�];A���w12�f���I����5@Y���jw�u����A�w>+#�Q�Ƒ��{�1�M�ߛ�9}2]YW,�"kK�4O3&[R�b3�M��t?~�ӹ~�ϴ�^	�P�����ls��y�����-��!˜.�����1![m����gz�^�˷S��]������u���Y2Ȃ�����˷Du+��ט�{�,j�����My�NWq`�Dܶ0�y)*�/w�'����J����*��q��}�� ����Q�&�J�Њ�6[����X�{�M� �c�7)��A��=��_z�08I���J$���Em�|_Rm��bV�zחQ�^hR�V$��,U���k�1E{*���Q�W��vg]�fE��
D��,�[F����7��{���k�v���zإd'��tk�����
<EF�=]�
��!�O˺�8,�����}�s���P����yZ��ہ;V%[M��l�HM�(�!c�]�M�q;lT-����>�d?'R����X#Pa����U;9Ee$Ⱥ�V臔���+�CS�|E�g/ٜ@�	��}�S�.T�DE(�I8�Ks�E�z�pκ}��ΰЂZs	����Z�@u*^�h6�+��p�T+���"�ߚ}�`:/Mϧ�"���u0�������*��+��Zh5��nZ�y�ͺͲ�%t��{����zg��<�!>�u����՗�Ii�"���_��w��U���`Z�|���qK6;��(hf� 7�-;� W�wN�%��,2+x���7�e詳�K�k��꯮��ӻ� �l��V��}2��╣k���y��]!�d�[��Y�핚���v���R���-�
 �xz��ᐶ�1p�y��|F�dV�T�Z�A��w�]��b��Mq���L��l�1&����6-o�Hh�Oi�*�O:z7����uq�KFgk������5ru�v�\�l��^�z���3Xbj�5DKYdF�i�"�/��[k�1��N�;~^u��[[tk/&N��=�o4�+���q�9��H�4�V��L�E&�PT�4��%%X�!�
�ZR���4^��3LkV�����q����#fM�A� $���C�ٺ-�H��0�>M���=u�&��(��{�/]bK���F��ٚ��kY�M��{4T"G$}�k'�*��jC,�~|v���d�w�~�j̢Tޱ*�wp�p[�}��Da[As7,�4����@��b�iR�5Uj��[&F.���#P��Q)$���"�=]������v��ݺ�G�ʪCHw�p]g|�I}�:~ܱ&���;������<ڿ��C���p�T��g��4^��:�l�d�r��s,�e�u�f֢�T��zv!qul�J��n����VY��d�΍�bn5�\�	@��j$Y��YtR[�2������2&7��5����r�9���ėY��H�˓\Xݧ�Vi��#A�Y�:�RU��������غg�M�1��`�ch�p�6��L��F�E74�Q�h�n�u��(��c�l�W��q�{a�.�:�fILcSbQ���!�r����!�m��\ �㛧�;�Ί%�����K�����h:�7���ۍ*^$Vb0��E�9���p��b-�ݢ�n�rp����)%��tɂ�2�Z����+�i�9Ǉ���H͹�>��w;������n�81�#v(���7>��G�mO�!0���.�7V�,�ӵ\���{Q���wp�����μjr�a�����pr�1#mE9ϰ��M�S!������V-杰����*7�D�a���kh�P�j�vOD����@} �Vb� �Mӿ"	=���v�r��w�����Sj���I���i�2;<���<�X�EU����Q#H<W��/☟I"̱�*�A�\ٷ�M��HO%�ٻ��=��/a�t�?Q3-1X���ힳ��_#K'zw"�s���Q����ȚA$b�2��۰	u��Í�^��=w�51�%�tt��2ͦn��(���2�IX�i<���:�1|?{�_%��0���L�,��h_���1���U>�M	Vdmg
��5�qe]B�����/ai��DHB����Y�2��ޞ�gc�W��w�qH�opB�Szf�ϘqH���ujAD0�eڴ���꣇�\��a<ꙝ�Ct.eL��W̓.�NN��I������)Ò�*��E���+�H�Z�&m��3og�ܶC�uj%�����w�e����&�,4�?��>�ڍ���R��*P��<3
�X�ފ>���F�d�f�k�[T
-
�;^�0ܻ�yz���<8�7^SN�_.����e��4��W%-J�0������Y��WT�G	YY��VF���k?t����m�*Ξ,�u�z��E[��M�%�㥥҆m/tH�滑O5Zj��a�h'G���.+gM���=���x�4����E1��Eh��+쬽>Ʋ�1�¼����m�1��*5
�y?m���۫��rǟ�u��9N���v��u6��>��a�P����^f�k���z��ű����H%u�C+z�]:|#)u��yU�-E/U�u!�5�����P��=U{�SUv��<`i�ȴY�¨�Jr��RF�6��8�
J���^���A��=u�P���� �]�����zQ�]��2�Ӝ!�Vh����x\��K��VG+��<� �lR�ޝ��~�2$�>eӯ&R��1\�m����������GA���D�2�G�<�;�Ψ���%].��>�P�V
io";m����s�[wr�
w���8����Q;��t��׌�X_%��q궫_���J��������fe[.8;kS]�x#)t��<�!+s:E]��=ReK7f��6�8+3SVX�K��k��H�5���:��67r�-��4��q��N�ɏA�{o��;��wk�z�0j���e������K���<6��*��i<xVRU`��ϗU��Or骲�5��]9c̷�,ܛW�ູ7�F�Ę�����!�Uҵ[ �Wy�n��I�$ήs7h3�� �-�st�Z��E�OO�THQ �z�r�Ƚe�K��k�	�n �%w\����ʸ�EӶ!�V��{U�N]�zʀX��F7��\�C�cx��Q�s����'�얠����*�E2��õ�|��M�����h�&�@	/�a�{�1[W+�u��y������f�Fɧ�]%����R��)��׷���d�f�JY�}D�C��FM�
��;�U>Վ���]d�MJ�ZFӭ�ӫj�ݴRۯ
�zx@\Xl��-�mR�zY�^U��YYD�ʑk�J���o(I&f�I��Vt<��g���{�ӱ�yw!>6��E�C��ꕼ�6���8�/^]޺��"�᲍�5"x�C��+�N����t��ڽHO��'�rx�Ua�ySo/��X{
�.�P�*�8yfeٟ��V떯�e4df�@�.�<�f]詇�[��vx��cʕ!�ܔU�������I�
�@�nԗ�f^a;,[lM!�W#~&́�!F�/	ɼI��r*R��(�qG�^ء�aL���[\{(�~�[��M��IR�C,�7�k����|������?�?����9�N曵ck\��+uR	��M��X���Ҕ��+�aUe�~���cJ+��]򼡂4*a^�OU�s"@�Rgqu�U~�f��J�a�˨����j&wC�0"�*F��q���f��nar�!�7E���lDU#6��;�n�z�uC��g�����n��w|�����ZR��h��� �zS�o��y�n�ʕ�ܮ:�Z��y]௡oe{�!t�(����vY��[�g�'�~����f�-H�{�X]E���Rm����#7kA��j]��3�޷xZn?8�ٳ���wgR�!�&���r'�XK�Y�~Ș�s[#`�h��x����n뫂�u��_[����m�qD�V��ed[ՄwXTYߙ5�]g��nf����m�b{�$�wݸ�v�d��a�do�ziX�;)��W���1���f��mE,	LJ�[���Ԏ�_�-Z���Ќ{t��-�-a
��\�,�V#5�fPM5�5k��a�l����<�߉5�t���ݟ��Ȫ��:���ǩ�00�}R
63%�G��H2�9v����y����e1��3�����V�ϕi���	
�����-��dl�rZ��l�Q��>�1PYӊ��d���]�|��˯<����B�f}�E2���Z'��Ȭmr�o;��98�m��#П=��Z�S#Jeu<�o��Py+�{��¡4s�D� ��YN���@�t�����,�֚�Э�*�4Ы��ɫ(+��"J�����F(K��j5(mD��ѡV %+z唪�'�mu�������L�KH�{��mU��Z#��}��3`�(���+�����8�k�L̢�\!^�n�{P3�-�KF�^D��[�D2�Fm<�=��1�t�X�ofN-Чy��NVL�2ե�����!�I��1�]����nCgW(گk={p���ugr �83�!��{e��u�x
�')�;x0��Ɲg���P�S�\m���*�h��Io,�ZX[���Ƒ��X�2UyU1�N�6�f͵��${pu���7�뎹t���Ӕ����n�}� O9��t�s�4,�Nɸ �۱
n6���i�G�{]�"L0����(�^nLˡQ��[���/���s�����:�+�����n4CR�,��b2� Žܼ0��ܤ"��k��#d��.�f�=V�I��a㚥;OoЇI�������d&$,D$�(3�\קϋ����ޗ�-��*�%3u��1���X�x��o��"D��V=��v���B^�Z�.*ӔmY)I-@�	G'S9�O���]���!��L]�K���_�����^��f�q��@]q*ϣx�� �����Ĥ�-@�E��n>��u�SVf����[��{t��T+��W`����F;�f���j�����Rep��M�S��gaɿ=沍�XfV��.��
=�y������Ss\�aE2������:����Xʻ�/�Di}�ԯ?�G�S��{7Bܳ�P�Y!B�n�.ɍg�d�<T���7a���YsK�AaxՑNP�5TK�W}<�m�C}�c��`�目��y�)c�L[}���ʽL,�װ_��u�E$�{Z!U���l6#TK��q���o���u}R�YE`X��=�=U�MtU�[�3M[�t޼�wU 6iv+q�f7�!�y��}����D���͡I�;�*[��֩�j�;�u�¶�eu���E���#W�i�lL*��_LkH����.�儷g�2r�M�⌦�!4��$t���$�yUS���=�ܝ�<���Q���v����Dwd��5u�6���W�}|3.�MFL��)��}dB��B�V7_Y�	0�	�Mf�VPwZv�Nb,�dк[���7���-���h]Eep|c�Sf!r9����g��G�U������LͰ�+�|�%)&:�W��dP�a/m3��k�:�V�L��'	�U�5<1s�T}��X�`H��0�iO�;�Ց��S�y��`�K�j�^��n����bw����&D�q�WJ�'_�^rC���\�-�q�P�dzJ���C��|��3�u�B���Z-��0�.מ�M�a3!	8��_d>�+�34��OM�p�i�������<�ֳ�ϴ�w�!c�U>)K�zo	2Q'/�g���{�����ߍ
j�#tÁi�\�JASZ�z�X�{�k�C�!HSW{�%w[���E�g�,W�X��-��{WQ��QVg �w%-�4qL�o]��5Sܠ�S7urX��-�������]���}�S��k�ML�(o��͸��Sε�ѠDb$L���e�k���mIOm�BV���⃈#��h�x�chF��j�d@�
�c����ͯqO&2Jz��Ci����W�n��U���ۄ�ힾw�����6��e*(��a�Ȭ�b�"5�qޥJ'� u��?Q��+�}uu�Q`ؽw')�&[�[�Af�n\�whq��8cS"����-�h�ѺҳV�]`Vb���k��;�{���tD#��1<�)�7Oݳ���8~H�v���{9!�	�8��nڰ�@���^��)3.$���G4ͦjƒpE0��Ԟ;*F)q����WSw�D�X#�,��}cO.�U0!��Zx%��4EK�w����C&�\������j����h����Y(��o��-:���Y�}�zGe�3�v�w��}���O#�Z4M���i�<�r���B�z��9g��:���;	�خ��5^�|1�$�n�}^Q<�ƂR�2���Yû����j�8ɛV��O:��]jݢҿ�6�-;C��h;!�I^v��h����zȻ�:rw���CDm�Q��N��>���xl�̴��A~���t�%U��Su��}�7C�}�[���o#�Сy�*�K#�����ҭ�W]A�ZXl����0�d�	r0�C����-�1�6:v��bÎ��h�T� �g�9����v	\����H�1pd���E�s��e�n���o�ҭL������䦴���p�h�����M�����~�P7��0PuV�����8�,��LNG�_Q�/�[��Lx�{Z�쎦ݕ�s�PL͕7jm�Qd�#�E$6n�d-ػ�*�{7I�o�R�pջ�:����H�ղ,1S%��0�^ƺ����.p��)'J4��u�<����}F嵓h�6n�q�2P>.N���>8p�[CK:��*�Z
V�OV��G��#t>���B%#�N�}����j�D�v����ub�ռl�Mt��yT!������2O�:zQ�,߃4��W��W�)�<}��lnXo<N��ȶ��m����zn
��=vV2��c�!~ީZV{��+%t�Gզ��T.��׳bRf+�x�j�՗�Vړj�6	��+;L����c�:ɼ��s]���v�A��Z+ ˲����j�n��Ի�-�7�3B�6RBGs��d�W���.8	ۇ�0��i��+��V�������c�n��{�^V��f�#%�v`�h�l��`]�ם�nB�c��Jv��q��%�euK�W[3��q��@���`hݒ3���y�5ƹ��m���l�ю;!��Oƪ�8��Ѷ�����1�n�+��T6Lɸi��x*K2�9Cй�ߪ*�_�◣6~�c�U:����R̦OWnP%��I���v�l[ݘ���:
�SM�02���R>�VU��@���v��xb�Ug�U��J.�.T�QO>!;��5�s
]BzU��ѿ���/*6���6v��!�i$�*H��{Y���Yï2q�.N����ng��j��>%qq��N,>.�U��(TA�<�)ƛsF���Y�:_/�}�~��y��u�k���}]t�t�Qԝr�x��1��y����\ok�z.������L����G�ݰ�ڋ7{~^3��UTȢO����۔�֓b�R�\�`+�w���2��������9�+��kb�����:�=m*م�e#$dH)�8�HCó�HB��=��^K�m�#\�F;X�s&s�HO����F�k.�Sλ�89m�W���)��'0��)i훌жݍ� ��~��D��4K
 �O$���m6�暑س�#�wU~YZ�w�9YPB���&�jl�QY��]Xr��^����Jd�ڪ�F��Uw��E
8������yG^e�����${ZVo�Ǻ(�tճX�` X�@��G[����ܮ%���ߴ]�)߶���](f��z�*����m�������H�dA��RQm�Q�A�%��px�m�ۧVYGA}�pe�CLB�eJ��'b�E"I�P�� uqM��{���n�;��.C��,�NE|'f�~�)$�oQ���fUxT ���Z�ۡ�uG!��)s*;�"�a�c�;�_�o���˘�+�y�N5�[m��=�gl
�Spw{�X{gV��7(��"�]�*�ٚ.�^��?!!���ɽ���{\n�ٌ��llNs�Y\Jn���]gx���2�9���O;���>^δ�a2��Kb��r2f�E,�]�Ƴ:z]����Y-c�����l���Q�vI��Rm�w~��x?w���Q�4�-���U��e�`���Gk)c����:��/\��U��~�|F�R��f��h4�hC&8׆Z|��|~�i�辣�ҥHt��Y1������;ɢ��[��&�B�v����'^HJњo��Ĩl:���� s�R+˨5��fP6j ��É#�ͮb��31f��/ԹGa�j�e�m"x3�_��̌�!�H�k����uJgK�#�d��AE��ݜ�x������^�]��W�o���y&��=�w`;^����,菓�,�2�������G�����=�}=vMn�v&���,�|4�uҲ���m�zA�cgJ��������ߺ�u���鉬�ޑ�&��6mx�J"6ڶ�y�6���O�܂0�sKep\�^r�17�w!�
�Zu��O���fԪ[o�2�ۆp�wk�"�y[��8�14-/����1��zS�#M��h2���1Q����>����+:̾j�j�U��*��9\3}ਐ�Sk�ɞ�1mZ�X���[�~��5��q�X(G�5��2%�UZ8-B�G�����t���ݻ�vg��8�^�a�h�+�cD��Gu�J���aIƣ����{�pU����>Ï�V�;)J�X���;���2ҿm�5�L�^0A��Uc&�:_�|C~/J��ַ�W�M+o}�X�W�[v��W�EH���ɺL�6jh9�ɼ{\�Ϋ����O+i�ݛ6d��ϳ�ט���*���D.Z��U(UW7�Q�18�X�~��̡����B��A�v�Iz�;��M�b�lw&�D�B���"��1�Y���R���<ݡt�1$��W�n0�[�#"H�b�<`�u���0퓇ni��i���b�W:����5�����>o�<xj�t��BV�9�n[��� �u!W�6_;�Z�{�g{�u��=8}�n�ֱ�q����kb�۩��uA��6�>��^��cpem׏�f���G.p6�����pt�S\����YF��������!D@��n8�ŵOPjS��"������O�>=�6W��춁{���H2΅$�ڶ�^vsLQ�랪ɜN8H�pF�Dm����SڞV��Py����8NM�u����
4��]o1u����f{ �#��M�b��t�[�(���2�`��2�p*�� ��^���z=C��.O<��t�Z�W&�6�'^�l#�P�6og��\R(�O_=��,�"�nyĐ�w�Ͻ�~��5��}J\Qӗ�I���s�L*�S�{u� ؆��|����Xu�M��b�7g#kj�]֎y��o�l�:���zqyOt�A�O��R�N#�~�RKA��Y�d!hb�ҫ�'�ܱ������񺗃nu�+���"��۹KqZ	�v�u+�	��Gz��<Rc:���dǃ	��g8\|��^���P�6��lv�n�rPw�Mԍ��x)��Dbh��RU$Zrê�Q��+
n����˶��f�
֗l��w�
�����!et̖��U���������zȱ)����c�p�V���O3yRR)�x��|�
�.�(�+�0͚wV�!{m��m�!<;ג�y��ֳ-��"�آ��/,@��o%:È˛�Eډ��Z�w�#��{y����hne��<-�+�t�|/��p��t��Ȫ�ٳ��x{�}Q��&��<��V�+��������Y��5,㰝n��µ�Of�܌G^K[�Ø��v��P�פ�gF������
n�z=�͆qD�U50j�����:krbҲ%H��aT�[>Zѻ%&���N����g������s��¦�o�暍q����*�f.��Vc���|ȨS�]�
�Xj�)��*l��ѫA�g�l�n�':^�'������vج�no��Y�vF>�kv�{BL����.�ݮlWx�"�s!��^P��];Xwj��Yx4=_,P��n7ֳo�n�7�Xۛ2;�N�U��*��#[�Ԟ�]����k>�
��n��{�w��g��" ��[@/.�kgc�WOH�mr���8�Ƌ���x����	�#\a�	�����nb��P�PGx�����7\��<e�%a�zt�e��*��vk8��e8.��׭���q��^�ruz�l�;q��n8\�(�{Dy�˚�+e�ȕ-�8�*�ږ��p;�ۜ�����s��͊\��x��������Uݲ�n6w�Y�VS���7��_�n8�v�nݑ\{��ܽe������W�?-���호��=�9�B��l�Ek����ԉ�Ԧ�������m���̤.h0	H�b�l�5;@�e��H걓%���Q�<�@�V"�8�R�7Yk��
����.1 ����n�����[[э��'FV��.;[�9{^Va����^y[�m�s�l�+��ݴ��]�Ӯ��Ӎ��u�@o�|�h��"<�/,l�<�����d�qI����b<8s`��ɋ���뭧JRe&�e�4x��rA��[�5Ye��k�z�xF�Q��6 ��0�g\K���ݐc\ŲO����Tu���e��GmV����^1HpoY���|�m�����lULi���m&b����og�C�:�f��f�ג!Q�>�8e�rW�����+ט%�J�2��%�ڹ�.t�3S�.�+n���Q�Nk|�|�G�]bNy�#����#̫kr�7opC�d��S�:�t��ю���b���&.��l����0�ج�4�[.Y�ٛ�6q�J�⺣#=%����Tt4(ф����P�8T�f�G5��Z�j#.Ńe`��v��۲�9�p��Օ���f��.
K���G7d�ttr\G.]���k�v�1�5�pWg ��] ����u.L���{vMà�;	"�vq����j����ZƆ�f�-e��s�䒭���f�h�p�+�"�),5����@�848ɘ�!��>�֣n��
g��i�,�'
�<��2Y��\<\g��]�p�M��]4r�h�XF�CM�^krL�����SV��;�{zݎ��s΍�7�8���E�.6�-q�2D��rGK3���!`�H:�hzf��nM��@�N�6M>w�acM�gtF�WP���	R�;5��.3uw��3-���Ĕ3 L�dX�\��4�}t��p�)�q8ɵ�뀮��e1Z�.Ԗ]g�"Wo\gv{�%Y�����4ٻY"+SD��ѭ�8�Gnmr�iu�,f2�WB�����5��m�c9�r��y>�|9o��]K���cl1�PI����]�tW�����ŏ`�����,U����][,��N1�<��#����1�Ɨu�'�uم&`�:�u;/_�8{��'�
(R�jk��ٔ�0�8ʃ���8s>��������{K���B���m���i���u~��1�܄d!��c���֖Uyڍ�fK���OG.�F�s垖A�Kr���8q���6%��x:D��w4�\b�B��I�\}积g{��Y�Y-�}'Ov����M������l�;_U�E�^��λ��]�w�W̊�1L4�hE����~����}<�	�/ύ�Dj���˩�X-�<��6j�se���ֺ��,Xj�J�����[�k��=�ղ��*��L7Y��������N�'mĝ�MЛ�g;xjݞ�sG�~� "�+�\���ǂ>SrmE�n��ȭ�����K�Z�,���˳Zy�&�XhcT>`�j�+)�(O[�Mn��&�����=������z���a�^���X�r������XK�^�[�(n�=`��XTu�n�=�M�j������T�d��G�u��QJ�uٵ��;����?m�c����C��.맭�ƪ���7��=t�����_||�sh�8L	��;.��r�R�:C�I���*�:ʆ��|�(��*r��6C�K�Ty�co³}mn���q��M$7$�Ocg�0�mj�t��3m�cm �]wI�c����U잂�9a���U]���8H+3��cTW����t-���u�_1�&,E#��}¬�T�fX�`ߔ�2*��v�:ᄚ�oE�A�>��2�F{%��W�]>��w٥�&��1y�z������w-�H\cD�fB$J��D����`�w:���NN�n�%�5��2ɍ6ཻ�v~Œ1�Uu�.PɃ|o�y�@�i=�����C.��[�Y�|�̿#k����*3����MCp(\$�����d���`�>�x���p��Y��ڑi�V;��,��A~�])���(��%3�Z^'�1�w���1��Ǜ��]�⯉R A�)
X`���x�}U<��ܢM!Y4n���X�W��W#X�v�s�����n�d0c��L�A�����m�SǽYN�S��;k����*�����{=���^������H��L�k���"���w�8��%$������J&��3O�W��g�ʑ�꫼x����k��C"��;�u4< /t�3շ!����Z��:�a���~��w���ʸQz�������JQ�Y�:m=�^^����8��aG#�p@����~�}�b�#�����l]."+ӝӲ��xA5�3�-V�1-��� �&(B�`݌�m��9���N���Sqؙ�nF#��Ʌ/�y}1��U�uT��]�_��:�O��� o��?K7�խ����uY-�<7=��4h��8�1��lB܎�g��ƱA{~�~�zy��>�Vk�����$
�]���&q~Ͻ'՝]�*����P��!-�T�(��-��F�G�ꆢ|8�sW�{�uT|W�{ݱ,3��vu��c���}�����Ս�d��|�,�12�����γ�z�+�N
�Vڪb���;��^3˥��͒�UԘnX�n�w��� ���S;��J�r�s<������n�i�Y���p�c��,ξL��3�j�F��n�ݷ��U��o�Ogn����o�蟂�y�^�"�kp�p���ò���z
)۬��4���W'�ըXy��{��f��l��gk2gҕ�tV���č
'�J�'�c���[��v�m����A��Ωy2nnS�-��j�t�S�ٛ�=u������=&����9�rw��-��9��"��Vl�n렡9�S�rg���+��x��q1M#�ק����lpS�FfY6'��9��ڕ�l���{ө6���V��^��̹}��ن�X�4z���l�v=�
�FHQ��1Ô;P������|�����n�h��Am�\Ip�����K���7o��*�|�: �i���)?xȟ��Uǧ�]VZ̵=�bXQ�T���W㍖��6����>H��n�ޗ�y%���i�4�CƢ�f$�Tfĸ������c������\9�7��]�/</������N�C���򉟣��ܽ�%M6n�*��f�y\�/�nŲ�ց����A&�ǃ�k��|P����9f<ܻ}.ӵ��"�<tm��2�|�*U��&��U�w�6�*�T�=Gc��D	H�����t�R1�B��T�4 �f�v �[Hp�l75SP�]I�s��㍨���LԦ-�lU�Q�+3L�� L�e��X��ey�{6f�g�+;�� �ܝ�'j���,�]n���:�Go���i��>Hp�pfγÞ�Q�:n���v6)7�-��OgV7j7S��������<
�z� �n���z�Ս��z��qv�mg	�&��g �nC11v�c�k]f�t�.%M2�م�����^�7�^���z�,�r@}M���s[�{G����	+#�պ���"?�u�{-��_]���R8�0� Q�c��Cm�n�CY��x���vݪ:����g�+��U٣@�K���A��V��lR�Q��.�%>Ln,�K�ւ����F3{�ޜ:~����ǭ����5�ȏ�4<!��N��<=m�u5�s�ҳ��o�ѻ}������s�+d2��$ф��W�C{������:nlg%eR�R{S���GM.��o�8a���g:���A&Ϥp��-��wĂ�ₑ�o��T�A�Ս�O��Q�Eg��1Ӭɺu�2��tI�1S�EŒz��˭�[���� 7U��-���*$���M�a�O��#&|n^!�ݳ��-��F\G��ct雞IH�]G)�^����u�A;����vz�맟���q-Vr�O�.Cg�M����Q^Sʲ�GN�'C0i���H�D��ãa�O�R�YM>��)�̳�P����ޮ�),�����j5�ӹ1[]�a�5��w�p;}{gut�$���<}��X'������;Q����
/+m�{��s���)�9�l��h'z��<>4t�A<�t���ب��u����l%F�>�zo�?_�1nO&�`͖Xl:������Y[����e�!
Ht�]�&��'�z�Z�S��Y��f��:=�B+yL�X8FWŸAD8���x�om+��,R{|�vw?f�8�j��r
�>�W�u��M5���g�<���z�hq��]��3�e�d����S��D���=��L�,�y���h.��t<x���o�j�C�u��~�\����m?Y�=�@�/z���.�kl@î�WM`LB�0�3-�[1��c�![x͒Z�E��D[.�
�m@�R*���$�?n�E_K���P'���g�F����Ł� T�	#[>�>�O����xa�dl󈂜1�e�"<mÎ:��/�˯Ԝ�ɾm����Up��qwDy��!&��w��so�����|��A7t�q0�3!��{�#���}Te�i�E�Q��q�<܍��BejUu2h���'��j�S�\��nq��[�B���z���[��v4�6K%�=��!�"�Bs����>yH���t��׍��k�a�[���
6ԐƓq"�Z|!��{�;zD��od7�;rI���U�4@����3[�^�!B�03:��o���΋3E���Aӡ�h�Ss��m�Y�	ŻޱJ몪�_7ca�m�����ڭu����yIn*U\��X�)�)����~s�_+L�W��7n3���
�/�%�%ɮ+^1�H�v�qYTҢau�J�c��8Yj�X�6��Q�&��$���_���/C����=#�[�_{�zB��=2�����,=hݝ���L�F&�E+�����E��ʒ�QO�qny��Ž���<���Y��j��IҐ�
�����Z�.{1����@��ů��0�ߝ�T�eb��Oz����n�}~�=lN��͡x�[�������FI%P���<(Q�J�&�����������/|;�Iʁ`P�!�͎�ëV˖ov�v�����(���=M�D�omf�~�#v����ڌzb�ƈ�2/#׺��:�fP����p��Fe����J�j݄I�a4JEl�n3CD�//4$͝9uǊ�sx�ɵ'�
��N͕�s�܂�i� ���P�k��hmw��`��us����L\��<�e-wo��)�w��Y��3~rvs��ޡ�gO��G���h���J�^���e��	�72�93[�i���ޤNw�y���g%������@X�rnG��<��Yi���(�e��v������/E1�x:�k��ӔŁOT�ʪ)�]�yƳ�	�����=��R�*4����u��.!��N��4�d�hK�5W�Xs��.x�I&k��y�kך�ĤR�.v��suSf�i�ŽxN�28��9 n9�*��mR��F��!�E���GU\�w�-x]\���^��vޫ��*n��ep������Ӿ�d6��4S����An�՚o��Zo ������s)���c"�=���̍Z�Q�x�E�7�:���Y�����i��CSZ<P�n��N�S��8y�T]�A郡� ����ಏ0���,��JtY���}Zv�����8�r�����b�^l��T��V>� 1m�(E�d&�|o����2{h��j5ݑ�*��[�����ʹ�ițA�MN۬��:���O((�R˳�-��6!1����e�E�Jq�9���Z�l����M�6V���� ��l��^ 1%[6���-a̮�cQ�v��ʈ�6ȍ�R�	�&�	ϭȲ���m�/�M%�⢺�����;���"k����<kgtp�*Cg������������,g��S��Z���ة=AVʇBtgm	�Nl':����0<q&bُln��nQs��$A�Auɡ�B9H"�a׍5T*������m��U*�~���;����zze��L\gb������5o�mo��򶳴6k�J��=��-ܪ��P�h�����^�ei�������N�e���	�tK���w��p%]r�ݼ&���@#�8��K*V�T�k���:;��61�p�C�wΟ���n�ۯ@�0s-^�֥�/{�)�a�����B>t�|�7��E[\gkW#�2�M��������+��G �^X�����1�*�v�zk���\{yо�FL�'o?DH� B/OrL��1��c�s>��S��=�
����L�&㛔�2P�B��U��-������\����-ߥ����ߎ��Gf4������T�i�����sTަT��I��umb��x�i�M�����ǫԳ��ֱ+&��K�q���[�P'�sn��P�9
�G��A:_�{���x���g�~�^o�ߜ�b"bz�O���+dͫ�f��6:X������+���IDX�p�{�1-�4�|����{g����;~�l%<��ʜTYo��/�K"bm1j�]��3��Ҭ�*)���i
�/+Z��Dd�5�{�������&wb�#G~���y�u*��˄!ή�ux�_;W�g�z�]�o���b�U���R6�FB����W�~�9�a�){̪��/���;6j����}ZP�t���ݔv��Ӌ�*_xb��wG����󿱜��6�ɷ�#ׂ!�����c<��W:��b���R'���ϵ�fh�6�{6�'���59|�+2c��I���iIr"ԅG�����^���o��(Ըec�7ie�=JX�X��ا��ꔗN�Cؚ�$�QN�Y��}w���X�-�&�Q�؞S��/r��7n��n�iq��H�lA�əC
�q6�o/J���н��1����g�����S(N�����I��nyE~1W^S�{�O.�N�K�9BD�$Zq��n.����)y�ާ>�%�����3T|A���Iy�~���
w#3�����m��V��;���ʥ&}�Ey�<�н{޽�Yr��&M�<���_���c�ސjU��W��yMR�)��t&R�V�s�[�F�ʺx��em��~�0�����V�$���ZmDl5�/K퓹Mk
��ga�*�"R��.��wh������s1�%�f�Rw+�Â��q���Y�m��V����:w4�Su�m�ź�N��v�r�]{�x0��+@�ׁBzP��#
{��B��IW�}6v����cVj�F��Y�wx�����A��ő�2��:�3�3���w9}/uQ����oZ�Ml7d�4f�U�ӡd�a���bS��6wr����-�����V���h2��z�Vޫ4���ƴ��YA�=3��h[����Q��P��mҷ_��w#����%��){h�ym��蓸&S��t��L���Z�H�ѻ/�d%V:��=�����f�r�҅���]DL|�1�#Y���:�on�u݃7��Ү��;Y��WN��Mz��&�74�מ��G�w-P���N��e��}׺�d��/���M��\�J[sKϤ�wF3�`\{�{���'i�*֠���2�&+���N)��Ew��C_j�v�3��4)��EEk�y�\�,/kM$���Vˠ���Ν��U4����{,j��mkɫՋ=x���O��7=��2�K�3+��EX!a'��y7zʔǢc�(�R�|�i���1�6�Y������;D�w�����x�a�瞑��;���hywۼ�<�T̽��)�]�3M}׺�!ۙOL*A���v��zń3|�PU��;�"��5�}�y����M�W�+L,9��5c�)��9/�Qh���*��6�~w_'wG��	��V��+���r�7��y5�"���;]yV���OIss�yp:��hoϧ<�O�y�@��n��;�G\�;���wA���j�qB@��DҘH5R 2%�/??
����������rN���yH�$�A����^�-��ǳ�$�9AH�eÄ%��	��U˚�pV�*:�~�Ϻ�O"�s���\����l�k|T��A���m���HVr/�� ���f����B	Mm���B܁8�E��3)�W3���/�xqù��o�1څW�D�u��y��������[%�3��2�%��=}�����2�q������_������aؘc4�Y������� Fk�}J�+(w������`�W�n��l5�=�Z���'�;G����^�t.���]m�&*;�h��\�DJ���;��u��v�z`�MO]*���w�{�9ܖEusR�$#HDL��AK7.�?�cܢo1����9c��S�s�yr�Y�E��j��e��>e�h�%�{PA�Vjx�Ǟ�K�7+ŷ��1�qe�ܴ�u�R���	uVL�X�+)�D�jE���紨๦�� ��⳹g��ѥ�ׯƱ�7D�z��+Բ�0
h$7׼f�H��m`���{��R8�
c'��#�)�f������A&biV��ֆ`"��kY�t%Xa�U���h��1�����D@Q��(����/׸\��X�7����|}����N��n���Z઱�{A.X_�� j$q��e�Q�Qn���c�����{w�=�@�TD��O�v<8,�tЋ�{�-f���<�-[��	���{���5!BB��JA�杺>��ϳ��4�5�/U�o��˭ң��	��ffΘ���MꤽT׳��[�䪱o{����#F [�&�ѧ�su= �hX"��{ee�ɧ �7�w��l���h�y*X6+���S*��x�{3ʯ3%J�Q����$�(Ҡj�#�K��B�6s����"n����i.��w�r��O9ƪ���Ǟyu Boc�EK[�z����HOyÞ�LP�mf]��,P�Ƶ�i�GoC9�G��4U-���&x��R%\���3MvJ��C�ol�`tNE��������[-��n�e�a�c!#]���.�v����X��b�Un���nTA*VZ��D+��(K�V�A����i֡7[Q#\�Ce��T�$P�ȅ[���#��d��ps�/\6,d��'A�$�9�X��5l�52�ׇ,[�ر���A��qB�<�㰽I��gNܯ\Nl��MuN�GWY��^N��Ǳ���j�'�W<[d��.kU�ό����j+b:�i3R��K�ۚj�$)7�B;JU�]�C�^$5j��ʻ�o��c�N�UC�����:G��^4/RR{�M�{5�뤍O=M�j�އ]�m�t��z>g�d�W�YrH0YZdGMCe��X�<72�m��]y�f�ɋ�zy�x�jjp�*���(��+k���E�ؽ_G�k;��e"�rH�e��Yw��;Us:k����7�̐J��fc�� W�r�!�)Whk����!G�����kuaJ^j"�>��I�X�F�LxP���L;ϱ��UT���c���Y7�'^�U����[�74�}�՜������D����'>�Q��[�[�)Q6ِ�#����Y��Ey��GnJ�Nq���s��]o3L�%�+�A[��o��uo��n��zG��T~��ۇ��x��f0R�����\'�ph���<���7ݮZ-vA/f���~�n�AȊ1D�]�b�R�#nj���uDf,�!?�y��ɟ$���_N��oޥ��z{e��jP�W�8���W��n��.��e�!e8�jCo0�6V�6���H����$C�Z�w6����
��yօY���Qṻ4�ۡ8���[k.����h-Wc�:��[�o�42�����[�Q�q�J�^�����ymj'5x���졗u�@!��{��hܩ��]'�)��4Z�HP��rGx�*��G{�&�^��w�mV�Us&�w�}F���5=�"����)u+�R�������B����(T-B��8\�<�Q����͋��=\�D�<�e8�]K�z�Io�Q\�G
���Y���{�=O:��-�y��w���?|�� ��.Q��|<˞^xܔT�=W��[�pB
M6'��V�x�u��TZ`�+&�V�s�1��bb�T�D�d$�`s4h���di4�u)�[v�d1�ł���&b��U�%e˿~���a�]v/?�f�T]� �����}6�Ɵ����2
��D�+:�ӡx�v�^j���%1�i����Q�>��!Q��+��a�
��,��w<T��.����Iq�0?]޹޺^�{|�d�*M�wd�g+��r�Y ��۬�_������RI7=��Jb���Ų6��%R��<5���]��7�E����i���δ�v����Im[�v[,�y~�SQb̧A-[�/�/F�κ�� �U�-��Լh�)A��'[t�f�7�E��[��9Dv+�}��x+��h����f=��:zk��#Ѿ��=2��u����p����v�}B�ޛ@�j�]*�*�Z�P�u�J`^6�y�����e��d�W�eC��U�S��d"G��4��2�WzPz�j;�f{��������(b����xrc�0�^&��Y���:�	�
k*�gCMI�Ƶ���v�L�8��nܘ�n�i��R�l�kn�l��"q�{R�%C�w�՟���WW�I.��TK>O7o�`��Q�˙�_o!Z��u�vZ�]�WDi�*ۮ�1Љ�)QF䒧d0kz�s�]���&T��T�JӰ�1��hB �}�;G^빝�|�Dqe�����q8�
�#J�nH�k�U=7���W��e<-x*[I��{0����Ӻ:�����3҆��_P"O�&R����6��$���~��7Dn�{}��?'ޞr��T���.j�	��3D)d]y�1��Ľ��9d�ޥ⥨������HW��Xg��!��8!�����GK��~O~���.�i\�u瓻���w��A�53h)�[z�/�9�ұ���M�R�L��	�!R8��VZ�u<h<�Ҁ�	�uMÞZ]��&r碧���z}�*��/���7G�k��":�����]��]�@��=g���p�؋�F"��L[(�Y[a�����kʮ>��ݕv��=2X�`�F���9=b��cj:��2:���������_]}�}����ޕ>�AXL��K�G�d��ں�>J��{k����7:+�#� oں���Qm��w�n�B�Z�my��X�9�cE�A_F}w�@-Q�6S�߆�c�����Y1��t�C�z�l����KI��ʏ���䭷tlx/0u�2���W�0V���s�C.��j��_�|_�F��]Kxy��b��J�}aE��Lb��OFIQm*��S��~�R��{<��>�V*�ݎ�Jq#-�܍e�k�̞��LV�P��2@p.\���h��W�]�����A����_�}�	�zX�=�[��öכ�&ҡB���
�-l�)*t����=�*f]�j���^��!`���ǭ��8aK`�ըҧK7���K+��﷐J�Es���%it�	F��$�i�ȉ��f�!hֻJ�,
��r�rbі�U�nw<C�	�86����D���n����u�z֍��M��<LUȻr���ͬ�������&ı�c��MJ��̋FP��W7Eb��h�na㶳G:�*�X�VS�>�ar��s��(�P�Ʋ��)n}w#�� ���̈́fx��@�5F��z�=]]�m<�2t o$u��9䍮ׂ���1�Om��/P��rWP�)��#7�uןϞK���د������,���N��zuUwR�t�,�iK����������T�=���m@���,��%����u�����p[{x���g��sgVLi^Bˊ{�XE�_��ޮ��P�-��?ĉN�Zꂸڷ���0uH"a%�,�z�[.W��?Og,��#�HE(h�~�3x���u]}���y�\�t���>�lkU`��y�X�F��������,��T��������3�n�"�it����U�H��q�z0�1�\U�q��FZϳ랻f�����]
�I$*8�RD��VmM���~�r�{�{�8�/�?^��o��v꠪��/J��!�s~u�h̨x���ߘ1��|U�[�|�rc�Ӻ6�p�P��a4�#53���ر�\�����E����ތ�}x )����"��^����Nj{��e��G��-� n����C8M/?~ӿ|T�u��ό�4�U*��}��t�S$wI>.m[�ڕ��A]A�e^����ub�y/�N��$�>��C�m�	�++w
�q㭕�U�-��7W.����
{*��4�B?]�=��E��r���3k+s�߂���d	��Tƿ'�:+��W[�5��p&�"GrOaJ&����K���6ǙeE<{���/V�7Y��U��6���x��'*z���s��l.���,�ƴplD-T��l�<��̿vxR�t�n�>�5���n��p�o{z]w��`E3���"��p�9���!kF%4APC�"�>�MDu��'.�R1_�c���^�}�l*E�{���[�b}�Vo/rk����K�gl�o�����A�Abf�%�V1a@����>.�rz๝���A�F�L2�9p���_���Y�/3�Եm�!�n����㦰#�������q>�ڕs�$}�Eu���q�?w�%�es��=~�Ņ>�x�
��Df׻��yu6�V���1ud
��+��(h�e�ןz����<�5 6�[���	����c#���w��y3фT^A=Ôi<��s;ru�'w�t��D뙏z���]_]�q,clGT��oK�
=r�[5�3*f}�뱒-h��Iȵf;/��)���V`���l�����d��J��פ;�B���P�f�����,D!Վ�����YU�͒�7<�.Ěƃ`��<��Լ�n�L���.�^��}8�""��GZ�7E�ޗ�e�v������7Y����'
?yW�M��װޅ����:vz��H�]��9��o+x���Lc	%�Ԃk��ʶ�s�焢�=���̱+	!�݌�2�QIǾ^]ԫ�,�%��ݣU�y���zr�o[�Qy�\�\P6vVU�E��7HD�_as� MJ�DX1�>�8[��Pjˤ쪪4~��������W�][���&@`��.�b�9�Q�U�ϻ����F��߀^l���R�7D�VAw��d�q�{�"�&}n��Y}uU�J��Os�hOb]�T��h�u*�X]ۤ�Oy�O䚚�D4vu"�$�r:��!�y�hK5d�X���{�6�O��\�ȼس�]�ET��縵�o���(z�7������Oϫ�՛E)��UVߞ$(����^g����ۄ��˭�|C�������ŭ3�z��[�N��0Њ�]��t�L�{�3����Dtz���$�L�j�Y 9	q9{��S����X���΢��K�X�7�m��ܞ&�.�����H��N�Ϭa
M�Ht�欟��8�������#���x�Kr%�=�����9݀�t�cv�z��[qWIXi���!$�Hbέ�
�t�r���眵*�u�I�r��o�'��U��=�+9b߭�^�M�K�]Q���Y���Y�An��~z�"�v���wWK8v�c�]�Z�s%��
���]�@���R�U�<�<U��=��<���w?{0(ґ�$Fa�GvP�k̯nt���ph�v-;P����C����CNo�߽/R���{Oh��ſ||i�<f8�D�y1�+���v�I�e�h�]5֙Λ���
	lE=�L܄�[����yF�G��̛� ^���w^��(�Dx]�"��"�XV.&]:�{�\��5G^�j��������`�R��on��<u_�X���N�"�l���:�ufՐ&�t��Is��ǢsU���'u�x�5�E:^[�V��{�t#͜���e�8��������0k�͵w3���v8'qlt�
�J7�N�^ܴt��r��s|�%�/ ��{��'*U`;��VB��J��e-�9��{R���I�ݮ]R��v��L[Wum�Թ���ĠAk��*u!8k��{*��O�,����wQ�����+]u�;���V��z�Ĵ���Ru��H�{`�;9�[j��-೚��T�\"��w/^���U�T�~�w�L>)g��n#��O�G�S����I�i����$ik�H����vc](�����wd�];n�����-��&L�C,N-�MK��R����X���xk�[����꼅�-�P
T)u+�i�b�뾛dmt������	f�w� -M�8��e]qe�Zطn�[):�X4$ᆵ��ʘ��).��o3{��ٔ�53/�	�껤�)ŉ�+�]�J��ȉ�h���3��nW��j��[ ��w���lk�&����+�'v�O�^Y��O�}8�z�'�$�A�ł�}��/uP�z��]y��>�P��W)�
��sn��Pz-S"6��6���;�7ۮ���]G�ejδX��&�;H���wj1��2���)VᲡ���u�k�s�����Ky����������NX�8�����=��!�{�����;����q�1G�q]�^�r�nvҽd��eͫ�#אm��/@��P:~K�ӌoI��A�wi�o�)X#���6�t4)���<�0�I �c���ZwO�9��0�N�@Ev�YŲ\O����Wnƴ"\ށp��x�Î
2��u�rVRfV�d[z�2���@��H\��Wc0bKrU�J�1��;[�6���Kp�iV�����W�5�c���&7^v��n*lu���t�
�z��ٹD���ɻ�pW��E��aۗ��@�sM�Q��cf'�����<<��7��x��n�}n�2�L�QJ&��sL˳��������6���#��C(��:�3%Q��k
���Z͝��9��b3+)���˗�pі�t
�pݷ-Մ�[�]Q�gX�hH�
j�W�B@c������j1�\�9�6����@�.�;r<{c��m�,.j_X�p�-�o['eo`��M�n�t��9����#a�z��x�监gM�Vf�''Q[Z��;����z�������FF �U��o#���<��p�=����E�8�mՋ� ��v=��+.�֚`��ځc�l.U��I��gm��&����ޜ�y��q�����gF�##6K�M�\�S�ES���㍵�سmƱ�P�.%��
fU+t�i�ūI�x%yn/�,��2ch�!�x�3�8w=\�]-���֎� ��6��m��U�+���Kv�mZ�
X��q��Sk�z��m�.���� nX;��[��Y����h�f�\ԭ��w`�Y���\���m�Z�}��	e��fjۀ�q[\���mE���`U�:-�� ����4�i,̳RV�Q�E�-�˖��`��̍#���[hN��9��v���3On���vEb�^Ǉ���P����n�)�s���&q���qk�P"%�B3J�����dۗ���Md��9�� l%�$��0�f�q�ݜgқ��m��l�)�;"�
z�:ɜI��N����h�����v�Ӷz�0��z×/kwP�ܡM���,7r�����z����ܻ�m�l�"�z:�\۷7f���SU6Oa�=�Gt��wCց�,[�`�W.�Zz�{q[q �^=�[�wo��9�e�ѣlwmN؃B�^�[��J�/�����t�C6��],�����L˥�\�A!�^�i���%�H��:$�r�PIE\Z�`�3Esk[C9��̦��IV]�ʒ�fbv�*n��.Ѻ�0a�\n��=�`���:k<'�7w#ħ\o88�6;g;�i�6��s5mncɰ���Ӣ�=e���E�6�E]n�u�E��p�f�+�'o�I��z�Vg�R�Q�5W�ͫ#DȒ�-P������SU�
���}K��O��s��X��߾������i���
�-�
�Y7�M�~ʠ�\���屑B�,J���^��D�F��5Oas�.ڱiB�Hʹ�߷��x����},��ן{�)^�Y����1ݟl�/�xT|*$\�2���[H]��'!i��.��1Q%A_{�:�y0�k�����:u���*ې��=����e���1\���/��,HY�u�d�_}��ր������	�\��߾���RE����]�up��Q˻dZy����X�cx/a�Ob��ro��W�(JU� N�<Ֆiߏ��e���r����x���_��N��9��&J��A��"%�{7y��zZTB��
��ٓW�پ	g�"�N[��iW����[Â��	^߮�����{��j��D���tE��7����6f�-�x��������2�.� ��g���]8#P��r���מ�3�5yn�b�����w�J���ma�A
K"����,K���W�'��]Į�e�q��s�<S�1����?E�ٛ���Hi�@Xv�,�� �~�v��N7�{A<e���Gv�QΠT'�Vq�{s�qq�b�Q]t]�O�u���y���^D�T%\mg��â�(VB�|�׿Vq\H��${�]�Vp����������!3�X�n$���`�w;�銋HSL��&F�J��A>�OΦ]*�t虢�.���-�cXa���(
sQY��N�p_N<ʟ�\�����(�o7h��sk^���^+��@.U�z,N�ߡ�Iiu]�M���+g	sA���2�T���lj��F�m�}��W�&z����.�I�0h�/�_�xXi���ZI�9T���oV%<|B],�N�!P�"������[Q�}&{���������ȩ|�!O��߃��qăR6�r�L#�9E2���X��rpAD2{.}���ƈ�U�v�"e�!P������uZ�Y�*�K�s��{�K���0� ~��S���V���֓B�E�j��oܲ�q�,K-� VEy���ߗz�eLˢS
T�fjr4��4{�+HW����+ҽ�W��>W��B�N�߻�j�<tY98�ĬW�ڊϹ�VB�;��q��.Z���SJ���-��Z��vi,X�x?m~��/�d35Ь˜EF�{�A"�6݌\����{T�UL̢��T���):EG�ZX Y\���鸳�N�n���L�Uڻ���������i)$�Ƭ�G!�~�m3��	��*Z�K��}�qBം��;݅�I�Ջ��sU�k:��߹|�T��{�S]J�B�GB�m���Mv`b�Yn��[�v�5-�i˫�E�]�#�W�,!2%��&*���c�ZB�i�.�|+>'���7�B�<
����ps����}�O�kl��g/�Xp���0K�U��g���ӂ`-��_e���^N����U	���-uN�#�Q
����H���w8t\{����-��Z���a�"��
�s3-���K�X�)#�'Ә�Ц�{���._\��^͒,���i�7=�ͭ<.�}�Yɺ����}�� <CY3%��u��Ú��+h;�?�����u�(��盕�<F3t��u���S�X#�)��U����kH���j_���?n����eYdỤK�*�ٴ함N��ze9B���YΦ(z�)d)�As# �5��k"�iKc7Vk�8�V�6�Ӡ����0S,Ľ�ǂW�ߝ��0����V"0b���RBu럇E*U*��:��XFSTqs�i3"�{����xMZ�x����a��\�,���(V/>}Q�s��8*�+"�5f	YB�';��cND�lj�^ %/����GVMZ��D,��Ū�Ɛ�	i$h�����w��JFd�-�*�;���XO;�셇� �{랺�0�\P��!o�M	׳�sz�Jt��sO>w�zR��Ţ��E[����~�V���̐����H�X���@��}��^#z�@�?cJ��h��/o��S�.��K�.��&�
��ϓ��pϱƮ�6;�.+����X=U�u�׳7c	��d*�ebF��}e��ow�7ZN�W�ΌgO��|�:p�$V%e�(T ����Y�ɍ�gc�c������z~����Zy%�PU��|@�^�Q�,_{�昼G�xx^=��Y��$6@���_�E7Q��)8��_p��!Q��X-�
���\,���*�<wN��o��I�4��|D��ެXG�{*Jۉ��K�w~��S��iia���������y��pbb���\�z�q��� �?��|7��3�$�h&�(�$y�cm�
N�@��;�b���ڸ෎����UD���
hn���'�H�Q{<�ZG��M�\�Ĺs�D1IB[mt\�N��}�+VpB֤,o%7;��'VO)�އ�m��RY�Sp���ҬT!"��~O�yW�K�i�����qa��.F8�j��,m���%�>}�ZX�x)����ѥ�s�;K>3k�1aR�D[R���vԣ���u�^��U��4ÒZ��.�wxs�K�}/:w5|6G�{öK3 �l*bohϮ�ZLk���]M�[˼�tJo;ٵ�i
�ܨ�p��N��ݐvQ��ep������g�V��U�/��,O��{�w�5�S�Ad)"E"���_�f�̭����}�,��vV�4��p��{7w<pW>�{V��V5g����	`��s�6�\�O��p�'����E��~��w�b�8�X�Q�D���t�qe\��[-a���8�w�����2�a,#�Wdmˊ����_�����V�fDH�	�'�sU��Z>j��WL�V+��"��{W
}�L��lLdӑL
�;u }�N*�^V.�5g�?��1x��i}��D����/?tr7����=�����fV$E���]��:)7�-ǥ0�I�����}Y��跺����>�3��c���>���wUƋEdP��E�2��}�|daްR )�vRb],��۪��ޮ��:�W?W�,� �\C�����|y��sMAj/r{/_nu���פI�	"�O>�uZ_,"��6��\������|\b(�׻p������D�+�\��xTy�=�[���|2��WEDa���
�߾���E�I��J�1����y��￪;��Z��yW�&z��o��:u}���X��Kq9{�3�\\jw�B�4��o�bo�rn8.���!:p�&�W���}(��ܕ�X����'��/8S�ޖ�.�#���Y:�e����������p�kp�K�d��e�n��|Y7�������?�k�i��d���w��z����Ͻ���K�}�\<-��֐c5��ߧ�-,��*!2(��dĊk��ˎ
H�ܞ�7f�!
��E;6{~��	�4��A�?�K��f ����td���v��=���|GQ4��$�J�U�N�M\*��#}d�"�|V���Y�*U����r��(E�qJ�@��m�FMuڵq��>�u�.�ե�Џoύ<�h�T�k�[w'n���w������=���j��i���{q���p76�yBd"�,�\Q
�.�ft�x�r�km]c����Y�פ8�m���p5�콶�������a�GHGe�d6������og��>XE���l�vLtv��{���Ɩf�mm�;vt��[oEb9�tgU��C�y�	���q�VJ9�k�-�.�iO�N�<���/:��(�YﾻZ/!L��R ��گ����p��#�0�G����M�ƀ�~�z���*����#ㆭQ�f
Ky�&��C��)�Qc
i}��Ow>�sRԧNfUP�u\XF�"	I�T&A��t�.��{�/�~���q�|��L��V5e��ʉ�������\:kH1�dP��w��I��b��T.S��}�����-|!jh�}+k�ܿl|-#�j����˞�Ӛ�m��4�ib^4VU���V}ObX�������\�����F��a	�g������D8I>d}���_�
��6��dVO��j(RCZ�faq�YI̬�IR)#��&�5*P�����SkD
ƥ���,�Ϸ镊x���H>��-� �k�v+�$9s	����ku���}N��d뾴����p�B�|�ҬX��9�s��_�³��iT߻6�F�_)M]RF���߇x�b��oS�����o>�M*����{��pRt��!P����K��>��sӻE������'ݕe�����ۛ��4ȑϥ&GK߯>1p[o�.c�$)��?��ݯZ��>����Pi���-���T�����%��em�5�G԰�j`i��Lʯ���/�ڙV%$��%h���*�ZXkh�S�ۅ���Z-4W��<�|'�LYm\�N��O�{����d��勧�8�"�
N�M��7��1ol�R��W�<gN��?n���1A��,��:��<��1�&1�\�
�"������:/w�_ܮ�7Yy�i�����]ɐb�����]�Vs�j��	-���˱@p�4Ů�༥�s�]�uNq�i�VL�/��-�KJc���v��kbSN9�yK������	��ӉV���Yb`VdȘ��s�[�yƐ�>w/�Q!�g!t���o{��&f�GT��-y��l<�Գ^^���ƶN��?|�k���ßm���U�{��K�i2���t0��F�Ƨx��>��Tx�=^W�&^��g�p���l��c��S.��|+��p���c��:T���<J���)ada�su�6�r�{��6~��M���#�_m+�bf�km�jH�Ӛ�4^ㅊ�|���Q�[����%������գx��?39s�|W���j���Y��5D`������B�U2�&L��Ťpb�6S��X5�R�[dW��Y�X���hSb_i�������~b���iY��R���I������T.��ىk-L�b^n�,��s�ӂ�
��TI�x�;Ɣ�{߽��Ǽ�cg���qv&0��=����9c�L�V[����Q(�1,,���&��ӷ]M�kXV:�B�������J=m~6�LO隫��ǰ�Z����n��U�,B�t+y�*�޾�E���@H�.��f�7���~[�w���+��%��1=s�b�;�ޫR �p
���8�[�����Kr��aN[�34�ipS֬T �x%b�h����Y��]���r�9��df���`�]�����G�
�RD�G>S�LK��
N���D�����ڡp�.���������3�MSV*�x�g����4��}����V�l�"w2���g����g�U�G�˗2)[S�۶�c�i;l�T�]=�Mno~��J��fv������P�m�fI%�� �rj��lRd���]��e�*�Q��o����(ɾ�R�-�#̫짪����J�{��J�zB�yr�Sn0X1/���2s����J�#�B�[�b2���rJ�y?e�+"�W�~����}''徯�јEs�w�8%�I	�b�I�~��-֬�!��M�
Γ.պ#�_k�������.&��z>���+g�#���\����Ŷ�X�ܩ9�J�4S����r扡�
����-#<��\#��b�;���`�p�&Aa,Ɣ�"�~��?^=��KX1o_��3{�f��������6�'�����X,"ϊ�R�u���gjH�E�	a��LRAG{��ֲo��vw�:���C�A)�xݣ�5��/6�"D[�(T�J�BD�,�9��l#v6�@��`h���*��s
m�Z4T����ѝ���E�"^�P��n&v��aW)4V�S�
��ϼ������9~�>�|B��EE��E��|���[�<BY�E߸����uSg6]L���31��g�����K�K%�I�����M��sr�c��ۜ_VI�}����,(ww��w���ƨ�)�ٿ<��*+�+��+�����<q�8���O{R����{��,#{���/o}%4�PT��uUk��}�������C��"�l���4��\���ZdP���E��<K��)x�=[��D�f�PB��i{~�|�Mq�QB�i<tB�����,������X��j�$�����ڹ��T&Pԟ���5��X]�������H����{˛K��{N,J���S"��rbn�]��8Ԑ"�S��U���8�7�QZ�)��fW����o땕Xv�UNQ���*�<Y�W�y��%M;�"�Ιh\Z΂,͖
�׫�/F�Mn��-œJ�l���=��2d��přS��TO//A��~������} ��ЃA^Bθ%�_#=�2<5o8��\|�ɅD�k�N�53���EM]�q+4AG���OO �>�RO>��E����Jm)�'��w�&�0Z-�mt�0W5�f�y�w���c�>���P�[g��;n'��׎�"Y��.�x+q���n�ʪvD��b��^m�����?�瀑*(��ä{.gk�M���u����aYa�}��y;^!QzeQ
���r~�qѯ��Y�}|�WpJK>�JĪiL��8+��Z�<�'mI�3�֝��|k��D'�^_l��a
�V�VD�>��;�������̽�cL���EB9W��Bk\)!��J��!�|]��epS��K��|�4�7~�ݬ]�OvԖ.d�|k�qZ�ϧ����G�������[0B����zA-�D��\s\-�t��]�� q��8]����`��*�9�@D�Dyf�=Y��|VB�^<ff�6�[C��p\� �q���ߝ�#u��,�6�Y#�Y$p��w�u�I,�Mʪ�*�q.K��?f��`������x_u�U��L��1iI¡o�=W�k��AP��vZ�&�������1��lֳ��!�^e�:=����Z���}Y��V��!Q	��ym��n@*��uE�s[*�VO��\#��t9�7N"��\��~�t��b2�aq?4�����!Hī�����ζE3'e+#��B�}y�@Zn5���bXE!r��0���}s�}�Xv'���㗨�u��i|f%����Z��]�7�i�"3(����/�6y��n�5S*U��KںD���g��*�3�؏,���� vx��V� �񣶥v��{-�cPn����WnwfF�;�F����x'��y;�O���ݩ�xw�]��d��x��&�M��О]E����%�$�;QǮ�l�Z#�a{]I�VoO`��A�mS]Þ��z��M�,�_9�ws���J�R�@�nYv���T���1 ����.$\�n�n�/O;�=$�1����x5����an����r�GM.��Z�-M���S�>�ƯC0�J�����"f��6�H��0�] ���O�+�X����,:�Z�8s��v�9��ӳ�����m�!I"RG��:X�����~q�)ru��&�N�7�/[�O����U ˁn�T��p��A𕐾����KE>�~_\��͹�NO|�7b_d;+=� ���v%�|+��Q	��>�G�_����>�o�J����#�W5b�#��P{1�����o!tVr{T��I�����}�,���j�.��'�ɍ>��8�db=[5S_;V.7�L�q�L"����\�����	ӋϏ��?�}�����
��s��WD���ir�R��#��'~1e���7�+�p
�[�_}�*�U#uJf������/��p��ޣ��K�}k�����2{ʸX+"M4��s	��<��.$O�K�Yh)�H�B{ﳦG����e��z�KJ��;��yEf�T�s=�u�-!3��)�EG�t߿~��P"@T�$���$x��	��K)�JY�<y,��\!1y�9ab���}�N��b{�z��h{��YV۪�
��͵�<�E�O��Q
��egܛ]�!P��S�
�C�Y����:r���}H&)ʚ�N���F4� F�T�9aN�`ܮ�W+�W]�9s���n%0�#>�����IՑ�]ן�B��W��'�R�''��Tp����@n}�z_yw֖g ����l�_��ણN�[�wM
o�}.��qe��f��ي��SE�\��X����S���=K���p��Aw�<���s-"�dQE������r�dV,�\�%��{{��a�r��es�'���,�K��Y2���Ϲnf���w���/D�W��!�ū�w	:�{pEϣH\�9�鯈�^��Ŧ��tQ�o%IuUJ��3윶�\��Ү�>_VpJN��Ǆ�V-|���zp��]��n�]X�X�c�O��z��3��c�\L��6�PQ3N�ń1I
�->5%�e���h�%��! �g\O���Ĥ��څg�����b�p�Ku�;з\tV�`��i�"�1�|����P��5V�U���]K�LU
jj��H��Kŗ�~w������4��gx\-><�෢[�Y@Y%Y�_|�j#�nW���L��B���>��b�-�X`�-/��է���p��x@�}�Z�>�u�E��M8^�9C�����2�2ԎE!n�;i�%G-�b��N���.�����(�{�6����g��s���1\*#-�S�Dˍ{��
�	x��.���_}��kw���V|@p�*��W��Ր��[H%�o��\�[mI�����b՟!��R��XN��:݂��=λk�j��:UM6S�O/=��?v��)X��s+4�k�\���.{fD�W���ݬ��:t�'jza����+K9�M�~�T�3�۟I��_����\��NB��aN��EJ��C,��������i�à���y?^��Ѽ�/��X���(u�ծ����i���Oן}B6����}��o��8�z\y
� (Ϛ�;�}6��D����K���*kH$�{�şxڡt]#��^��~R�_3�����cy=�|����2���ef��|Gŏ�J�6�J�}�-Z�'Z��Ő���V�ew�s�.��1��� ]w�O��A�f{�U*Cɦ<��ז�b�rl�K���HE��҆���ϩ@7��J��Xq��������'M���r3.�%$\����WKsY�e���8��qF ]&��3u��A���W.da����D��F�
�m.*C���
�\q�Ip�%Lm�癃��Wa�i�Q5WQ�Gu����ʝ
C�kT��.M��8��X��^�tp�j�̉��h�V������v!�.�^H��,9\�d��u��cyG0��*#��j��厬l�bm�Fe]�OzU������l�$��y��۽�[�A�s���fH6mX�����wU~�R�V}�g�ĥ=oV����j�D5Z�Z4�FI(%V�Qk���e����Q��ɳ���ҧs�kr�Ë;WW��/Ȥ�E�<�:�7�u]�O�}sZ���=�K���$u�/�"\��mN�b}�[�0V���%pܮ5�E	L���C������CUAA�=�]�t8�}���͝u�����hĞU��J�JR��͎�O��"�ZI^WA�R����!J�VAf_TM	�L�&���`^L��j�t���d���B�U�D՝���n�䡕��N`w�e��H�-ޚ����z)�H�u.z;B�yE]��5j{)V���3پ�����l5��UNl���گ����)uW��A��ңW�V���`�iC��S�Y�GR�{���72n;�F���S]!%/	^V��v���Nf>��>��^e�L�c���j�U��n!���+����Қ�+���p��zT��������}�@�Kz�VX�����ik헗	��Ľm/}�u���?�:��j�-)8.��J��F��W˼�ޯ�y�#�z���ͥX�Ƙ
��J�,�*�k�#���`/E"��On��6�WNE��߫�v�-ƕ�o���ԓӟ|�Վ��{V.���/k�t��Ր��]�,6Ñ� )$6���$.�
�#E�M}�<Z��u��ia՜;ߟ�������|)��G���eq�+p��iw�T��g���HX{��X�Ort������:B�S��q��
��՘������H~e6T��(Tiz:x�Ѹ�����Ǝ�sv5spm�<�}����]`*��R%ASG�V8RBfۏ�!_�ߪ�Zܒ,��ő�]{iY)"�~�@�aQ	��Z�3����"nup;�MS�ɯ�����6��i�j��d|-�����m�6�aYrQNu}���UI����rI_�����2�6Ydn�O۝Α���t��?eeg���ǥ�b��kg}��=R�`�M�E�s�/�ϋK�p���	Q>k�����\-�#��'�������^!H�x[�/�]�E*eQNf�jjx��</|����Fx�0VE_��ڢ4B"F�S꞉X�sｊ��s�/D�vUD>+��ߎ]����'�4��Ng9Y�^=!Yn�z��/�"��f|Z&��Tʙ�ʩ���-�����sU,%QN�rD�&>R��#���2�5��	n����"\4�qV�H��Yq�
�K��Ϫ���*!e8R}�LiU��i=_�|%, (����}���OZe�IԳ�V��-f����S1�}�Z��,��`9���%,��6dbp����8���VH��!�K�}�/��%��=�(�\(K��M8�j��r��y�v�4U0��z������ym��]V]����\<*�Yd1U5��_��p>����
L��w�)}3_;������p�K~tF�����p��SL9������XF���*�z}�˿�����75q�钢��e,&��W�����-4�˄�R����U]_y��G����e���F
��ӽ��p�\:*!}74%����Ӝ�NBo��RD��p�RE?_��	����r�U����hhXY�\�ޫ����6*u�	�JB_��f�s�Jd����K��� ϟ�BL�� ��R}>�]|!�Ǜ9�ݿ�h�� !�A��ث�ʇۯ�ȓ{0�$9h!I�S�{괼p��Y��Q�nq����حO�1�|,Χ��=��G8%��*�[�ޓ�����Z�����g������?!�/�������5��n�+!1|t�����Oe2(L˾��-w�y����.�{U�����,�+���*(^����5�i%	�Ji�"�!_��O�&��cr5	N����(�.�V��E.����.*��/��Ϯ��4R �T.�%���-�9ͫ�K	�i��bd��>��J\��mQ��:@�K6����n�_�w�����^:�aQ^�l�����鎎WZ�������2�!1IG�*R�Ʉ���;�� �R�?3�Օ��A�)��R�������ӊ��]8VQ_��;K�͞��ta6vR�,������ͦ���'������{�x��;�=��Y����\ڽ���z�gv��J��魱(�iA��ȡY��.Y�����r�C/ҡ�+}Cj����E*��`��m��J�53\%RheYj��n$yI�z�'��8D
�"b���.MP�a�u����v}�^ɱm�䭍�Zф:Ԛұ�J.�{y���j{s�� ��l��+�f�eļv�|�����ǂ
�E�AnN��cF�p��[4��&��J8H$��H��-6�͈�t����nQ#N��h���O�uc]�'R�����eAG4����Kͬ�綹��Mh =���2�١c3M��~��yb��$�&nsvꎞ8Z,O]��p�׃]t+!R!1Z��;��|�TG���;�,F^ܾ?�xo�y��򎒥��_Y�[� �0�zP���{Ő�F��S	��4�E/3��̡��:�1hH�QBT<�JĨ�������k�Y��־-���8/S��&��RE�߽7�9�R�,�)!I�1Z��"�B\>̔�W�?��)��\!^�A���z�����:uw۫���z�6mV4�������P�cU:m.���U��p�����ФV.��}��M!���+0[fF��6?_��%�Ƒ�mu�H��HVgs
K��8D��f�r�E���_l����md�������j�"������"�2����{�o�ڹ�@�[-l�_���>+��+!vZVQ�
���Ϟ%��~�ȨVD��$�p�w>/�>b�ㅒ�X+#
��qS\��-�}�k��#��r.y�xG�R�R)>�쓔ƛ��2JR�T��	�j"�
�B���ѕN�<i4/U��k��׎��^�Ҡ��_[�V����_��Չ|��L��}m'�6j��+C|�H�	�p��mY����~���n+�-�j*Ĕݥ�O�՗qc ]7� �rq63���V9	��-�b5O��␽n,VB�|z�.:{��,��� {�ĵ��?�{;1�¸��²8*�F��>��U�i��~���Z��B������ݞp��p]"��iQB�IBVo��{���)sL�N��9�R��|�*�WM�ךjE W�������{�5q����n�Y�X>�jJR�C
�m�+myy��%m%6�����"�h�҇,NvXA�3�l'�e�uI�q���o�9�K�>�WMg�,_O��p�Bdp[N����jg����)���3���ָ%�	{���15G�v��n��7�.���|Y����=������uϯ��f��,��˞x�\�������2���W+�E��s{�q8��p��z�*�Ǚ�|��8\'2W��}���p�
�ֺ,4�''|����Ĝ�uԱ* �������$�	�S��%��,'ٷ'>�8颓|�{�]�@]��]B����w�q�w79p�L��
#�1�w��k羛����2>��ұ)k�z��eqVgs����;��w�R:E�i>��,��O;���Ș���uk�3D�dpt���&�.����Hi�}p&P�fW�3˝���uJ/{ߦ�����(T}��/U�|WWU����k�!뙷�o�m��G�م��Wn=�p��S'�>�h{���43��%�y�.�5ѧ�P�a�����*�m��y0�&˲�Tg,��6;BG\J��t`�Xq�(E�.���~�^[�xZ.�+����K�q¡QxՉIg���zb_tEߨ���'�{d&m6 �0�<cq�z�-z�p���)|ɱ��>_OɕA3D̪N��UZ\4](@������_y���^#���;T�?Yz�2���0�ڢ3���"��Q�y�Ң�Kr�����v��y){]!X[�+��ST�7[��Y�r����h=�	!{ӯY�S�L���*i�\��]�_5b�5��Y2'&{���lK���}�.z�O�4�W͋�{��}��x^���^�\���e�L�t�>�c&��+}[T�ۣ��h�u/�Ta��GhRCԼ6�R���$�͕��*����	r�����yc�8��t�8��z�ㄜ4�X:F%lj�j���L�&���0��j$�|�{ҨN�
�47EMQ~��Do3�=�[��z�%a�w]#OY+�腺�K-�&�\���𳫳�`�>��).�s^��ξ꾑�?�q�h}�b�4Rn)�M��Hz�d�y��V,��{����I)�����E)�US�Nhnh�����*eB��(�H��o��ݑ��LH�֬�#��{{χ�>�mWމ�w��£�z��)��ZB���K��}ߍKO�(�[)2(��p�8h�B�xE��8�X�m��s��{����޶�Y6X���t5	a[U�����e�����fĻf��K,��Z&�Y�/��tY�&�x��k�ќ4�o�O<���/5�/ZZh��rK���
�~�,���ұh�f4���]�������yՕ>&��]4��~!�z/{wӋ�E�N#z�	�.׫��jhR����,���#�0�G���-�AW��t�������a�*{BX$��ږ���p���T*8++!;ﾫ\ɞ�I'E�"��ϖ:��[�}"���/�$sO{�������f��o{��\�.a�Y�'v'EB��a�4�s�E�ED1v�K��XD���o�kZpX`���E?t�:�.rؖo��rGմ�����xՋJ����}J��XI��"�t��~��δ��To|�Fk\���aܞ������s�gL#�9�n�xF?���Ra�q')�����Z\=Ɨ�ƙ�ԫp�榑���ivr}�İ޴��2\��g��)�4���S=�����&=���h�g*��i�n�]M�-Py�]h�ʒ�s�*���­�D�UlUסw�n��3�ڲX�?�z�������N�]0�f4����Ϫ�B˒6����;Wم�����3��Z�W�<(dXS�/�*��;B��gĹ�WD�w���u���;�W߈��D
Ȓ�RԑF	^{~/�Q�}#�5�w����8GEy���N83���,#��f�_z-���5߭��@ʊ�%B	�^�n�W�Y�"3u��{d;h��Ӌď%�v��t�d��uxW��E�r�[\$Z9���`�/w$��^�]#�&���,\#5£x�߳�q����ҕc�׿c��,�{3�_eA�G���|�j�M8WϽ�KM!q���}ƬTg��^8w������:�Y<����i��T���Y����������w�&_�����,� ����[�WP��G��_BV?���K�5Z%�B�
���J�[��#5�Kw>L�)92�JH�_�!r�����KR��氀�0(Q$�k�:G�Y>ɸ�!�a6�Q/"��T+0@��~{M}�w/�RB谎w��ie�Ukb��K�l�n���|�H\��֕��5�	z��p�@2�Jmʙ��� #��QR{e�����Z�k��"̦s�ܵ�q��ྷS�2�T�"{�s�!Vl�T+!����|F?���B�z�MSJ����]��~�_s��M&o�)a�mԫ!s��}��	�@:��j������V�5êJ��XCz��;K��L)�y��+BPg��ߍ�趞Q��r��_µhL���$��O���Ց�-����JJh����,\�8L������(EG�{W���^_��n�]Eާ�����î�P]3hQG9_�6�k��.8,���Ge���Q�Mc����?T�ta�(�0ęD��fhTy���X�Zh1�]���n/:��\bK�(��Ȑ�K;��m����*Й+a������]�`熦v�(.�^ʹg;��4�kQѮh���������9.%�K2�S�Hm�1/=��`:�q��]���v��Q.����lf�e�.���c��V��PiV%���`�\nJ+g@g�M�t=�{E�uWk��a6j�]�2+���	��^��ڄj�{	���@fu�f�L�ی5IL��tA�rZL��>�V-��^_�Y�\2�TE�N��.}?UƋ�9 (��%h�#HO�r{�$�����Y����>�	2�=ʛ��p	!I	��)��0ّ��b-���޶���"B��M�f�d�����{�D|-!�"߮c9~�im75٨���d�ִ�{�K,�s�;�Vv�$�'�+�"σ���DiB�}�������|�Ƌ��gW�����y�"erUrdT��'�n��\1i����>���q�WO��H^Ʒ\���O׿�G���Ƶ�ϰ�b�0Ra��}���Ϯd�F+�\KK�������k��my[����#	}�_3�Rܩ�QEQ3J�h��]��I,�d��y}����V��/�|�lX-�p����P�G޼��Z���:Ր�߸����7�p��8ҭ���q�]{�B�3�V�om�KS�s�ZG�Ց𾿾�yJ�L�t9�S34dH���8�����	|��+����q¡6�Lv��M�y���֨�'9jc�2����lt��G[�-�%�"��{��mtO���H��s���|/������>�/1m�"�Z	��R������9�����2k����,T���P�qNd�Q�\��?H߬ƾi��k��AI���a�i�Yt�������s�V� �T���Vݣ*!{����k�]��l�<%�2$�cT&h����,�� �c�Df���nl��jkm�DM�;�����������d/K�=�wT���j�߼��HVyӤ
��s99goP�J]�U!YQ�ͮ���ә���i<Y"u�Vڰ͂}=�]M�H�+��m5�:&]���^�B�u9_c3}�9���T+0R/7��Dw�W(��T��gy�Ԗ	4`��]�fо���L_��y�����^W��G�dy�vO�|��?m�͹e
����,��d�͸N���h����,�	h�D�Ξ#��޵�p���s�����i��U��.�s�r�R����'U{�Αm�p��)�T�D
��O���K�+������|����N��L�)L��㤞�\kH�Y�..|�L��s����XGǇX��|<GE��p_mZ�p�@���ٻ���U����RO��R���>�=ƕ�WRߵ�������7��0�|p�'��� ,��Dx��Փ����#�Uw���w�wW�'u�6}W�yE}�|����dbƺE��.���g|S��G{|�XC/�cVB���G~���K�6x-#��CܘSn,_}y����3E�.[���n8W�<�]s���9R�8\܎K�:�ֶ�:�On�xƇeX{c<W7	=ja؅l�ʨa&�\��4�4���V?�y�ξ}��jH���ȱn8��3�����Ր�y1�r2Eb�ip���|Z_}��-y4ңH�Wm/[[]��}�1�	Q��/���,v��St*�5-:*ibVp�Ց�q_�OAP���G��5�U��]��=�XE�+*��s�.8*�RE��>q6��3>�괾:/(}��{�Z)�j�_�mP���)~���_F�/��O�����OJ��l;ns5u:p�!Y��)��	����Dh�����V'�(	�zm`�p�4�ڿ������&��F��.�n�Z���<�}��hk
�.��Z�Ja۱ʴ�ɿu�}�LΠ�Rh�(�{B�2{S^���1aw9�1Q#@���E�u%�~��ޜ#�*��}񞵲�}�Fs��j��,�	�1/4T{���-߾�bó��X�����7�i�&�M0K�l�>�o����U
��T%����߽�Uǌ:GV�)�����w�9���ͯaze����f,RG5
?a���eȌ!�����xY�^��$���,:h��x�Z/�'�ȯ���dN������履�U�dWS��Sɢ���O��isHD���4ŢW׆�C��ټ=��-ճ
�&��lSKω���4e�sfWKn��=�m[��{k�&�#n����Ļ����W:̦QI�*���!i/S�D&H
�����jH�O��e�6��0�V�̿���q#3\`�ڐ}ʻ��iI�'�ﾜ�����瘟����v_�B�bRG���Z/�������u��6hX,�eMa�K�zW��\��J�	�J)����I�D*>��&D��t�ZX�����O�]yw/+�M*�_B�b��Z�3faQ��(��g�����*9i�b��_kx@�7&w������h{m�����/[f7�|���J����S�6
Njl�IV�1	X���_��^#D�Ș�7	�T/[b;O&ԡx�x������}�)��f�7B����w���#��nR�{kHb�Ϲ�q�:!F����k�}y��	��ڑG$v8F���2�d��6����Gއ
�if6����--L�bZ�£����U{>��'�
J���;KH�gz�?Lt>���\l���v%���_U�W0�窯�h��I��ɳ{gYOo�G>YpnQ��බѽ��~��|�~A��?M��[�"5f���,i���t?F�h��]Ǐ�~���������8�E����}���~��y<���L	x����g�BT"�����[�Zt�5#!e\��,O�Wu^�_|ר]{�+_
�~�������*ĸX	]_ݛJL!m>�f,�,D��3K]�f�'^[��iM�+��Y���7�+�}˗���Q��ck��i�\�F���l�����nt�{�kJ�bѫ����i�iG�B�Ҳ������Ɍ��ͨ�Ya�����ɴ�pbRD❥B�;Ɩz�Ϟ%sKT����8b�Y敔GŐ���;�ӳ"b�����j@TBﭟ`P��t�I�c�.^ϸ�i/qАt\=��5ʿ��,��.��cs���@S^��4��{�.0Z%E��Y��όKٮy�X�n�u�e��wU���D U̷���Ux��SJ��dX������T��jj���$JI�T+"M>�ݲ�f��3n�ҭ�kmt�]��7���g�}�c4\��g��?g���	s%��&��g��KM!�B�������L8B�Nx��fH谅X|��"�jjeʥ3S.jq'�|ppj�	�����k�������ߧL�<��L�	�\�l��ֈ��/�W��Id6�ۃ��^�����ǎ��g9[Ia"�z����|$٧	��S�B�໎�V���27R�5N�³H�Z�p��)�������$L�8%4ٲ��/��Y=����;���,}���HV}�F��-�Jp����|t�E󒕋D�q�ϯۦtv֝�R�#�	��\��UNTz��y�T$l�ء{ҏ/N3&����=*�c��굦�nj���۶Ε��5WOk���oɁR�Ү�Nڛ��Pnۮ6Q�;#���5�8��|W�"��vT�9�U�jy��w��p�r��km;�:��wurl������%�M��;.��/�]�h0�b��&n�z�Z{65��ˎ�j��-�|�X�cѺ��$�)P���{V�ko�֞��U1��; ���̥
b�t�c �\V�{���ҹڂq�6�!�B�R�"�٣�}���+�ę�R}z2'H�̹���������}u1��͚��� Y�^�tf�{k�p�T=J���9A{XVk�մͳ��X��֦=e�Q��F�3����a)��k�g�:���B��Q�3�M�7�Թ�uEO���у�ꗎ_�(V!�GFD��ԅ�� E�&�$��|Kէ(2���-���q�	���x�g�e���IW�3���s��R\���&䥜须f�|� g���;��-���CT�IX��U��L��,����r���m丯��\�õ�d;4�Q�e�5W��%*�0��-����y���j愨W{6-TR�7Y��Ņ�*����Jmnޓj��嶸9]�%�	�v!G#m5�"fu�K7��֘�_��GG��P{NG�cj�j鸇3EHGlJ*��u�3V�c��h�����{���BS�_7�r^+��U%}�]��:e��^��)Iн�2��Z[�,�'A���*+���u9M�;���3�h{����b���.���h�5�sR�,thE�U�v�(3�N��˷��q��4K�oW����I�s�ka%s��']��|��Y=nؕ��m��<h�.B�}��ɶ�9�k�ZD��2�-f��=G)�6���.�Q��eX|XݹǱ��̈́���9�aylZ�ۓ�$x�*W��8�OK��	��q��ƞ-��v����"ae�|��K��T%�7S؂��cãa[�5]�Բ�T-�9s�Mmu�؆欄�R+ W|7k�҃���;��t�.ǭN��5E���㘱�x�j8箬��� p��s("l�gqvW�n3��d�.��1��oAs�pNx�
kU[��c#�a�.�Ns�q��L<�s�C$!-��T��0�Q�6�����y7��A)�Jn^�$=DBn�L�{#��1�ɝv��m�p	�l5����l��̭�`���r�����]�:���C����r��vj���nN ���;��{m��wAXGB=�ۛ!x�s���%5m�nCx��;���]�G�]�V;lh�`�c �R�İW]m�2�−�Z��hYk�[N(1z7��[<Gmcv�Vz��]s���\�7S�n����Iw����-�{1�Yc6sM4΋���B/�۲]�9-��#H鞎FǴ�E����'��ƒ� �vu����ük<��6�<re��HJ��hv�z�ԼJ�[�']q��\�o$ p@�\(�����Tf�
P�c�$Ѯ�-�A�:V*�H�J�5�l�&3*����C���k���u�E%�&J Z�&�1��5!,����5+����o9
G�4��Vz��3�T����x2�u�i�����m��rH$��$�3h5��w mO8O�N��9-��s-Y�h�O�6�n�m�ہ��\�=iGb�Ҟ�7k��dpi����¬���a�bMFKّ��`�f;��ans��ގ����<xxBܮ���ZP���,�t.�vL����.����E��>c�;��طFd�@vw�׮"놓�۶��M�d�˭J�x�j�ӻq��p�M*ɕ6^�/�3jE7�]��mǵ1��2�E
�\�� �ː�\�l��l%��'�j�5g5�1���^���15�n�X�fP�D��ݲ���]��C��Ql�p�&�f�r�����xle{�-������>��%ж-`C
r킗:�"p
g\1�MXy�JwF���Wvm�f�8`�T͢��Ͽh�݋+�)s\X7ͯzm+0]�,���D�\��ϳU��\p��Dh��fc�}�,�#��}t����{;�O��)�Ӥ/oۥ��a1�³�-iY�>��6��o|Auʔ��/|�y`�ʡt\0�5$�.����5Z�>��z���ܽ�B�'
EDl���6�f+GF�N?�S5=L�=�_��e�Nߩ�[��,2�F��W�D�'��*��˩���^t���n������,�:W�� J�zle�!=�U���������_�����E�����^�49no+og�>�f|=��;LҒ=��>_*�ЙG���$�����S~)_�8-��,�*TŃ/ou+�w�VE��EM�%��շ8M"���N{���|�m��cN�����_�e�q|N�bϱ��y6��lu����0�4DLEDҘ�x�f�Ռͦ�����b�`�d.�u���:����T��.Т3���t����bZ��Fj&�_r�go�>����۷����O��`8�tu���]�l�ʭ��Ҳ�6D�N�Ey�I��s���>W鯰��[]��:��W���hEbZ���Naꚶm�0K��f�IR�wkx����U8�׍Z���	��ǲT?ǟ9[�ݶs�w���6_j=zv��A��
R<�,�{n�O���"G_G�2:�k�%���~h�}��3�׼lL�6ʉ�&�0�`�̮A5��-�{crUc�Ms�
��#���F�uNx����of̴DW�Ӻ��T�5�$�1I*����Dw^���Viͪ9�2wu���;�O�CO�����"���+��s�U}�f�,���'�����Q�ҏ8Ye	k�V ��XJ�Yv�jp�*�5���эb�e$���Ϻ��<Ǫ��Q̪�{VevQcX���]E�^�4,W��Y�aC���z�-7^lk��]Xh��j	ྃ���6�r���'d�p4=�}�WY�������%gwT<}�6֟-o�\Ǒ��ABOwtk8O���"�h$�r'/Ө]����0�:�-�Y�yh�HG�  ��m=��U�d���1�Qaf�Z���bb��E-�!T@�zuowۖ��K�0���h��+^Zv�Ǫ��p�<�q]]D	�Z��vw�F�<��0�Y��9:�oz�'��q�I��V��pɺ�~�/�~U��@�]�!f����N�����^�7H��w|��g�{�`M�����ձ�mW\���\i�ӥ��l�}r��M�b�r�����2F���nL%����{�|O&�rw'��&Qy��n)��9|�غ�M������Ղ���]6m	���	[��̭�fxE�����>��^W]B�ք�w.{D.y�݀�i��y�=[�ߨRW]���Nw*ҝg��V�o��;��6#s���Wvn���m��]����2�:��o��v��Q�rK��u�Xrt��ˇ��vZ��YTy�߳rS�\"e̑B\G�"GiX���Z�/fbG��߶*����'����Cٯp�`ב�7�������]
�xz�h�\j6�p�j�t�ں+�=��}����wkL�k+ڞ��#���>mٛ�V#>�/�U3$�٢,w�MԢʕ��X�ue�%��쫺m1��f�jޑ�H�h��dZۺk��X�)`J$2۽��>�f6
��d4��.�&+�D�}Q�^�_r�^"<�E�L�z2����
����:��OS"��u�N��^55�=���Ë�Y%k�E����kh�KclI-�&m��lR(�c�56.�.q�Ļ`2�0�r�8t��������p��]fQ"�g�ס՝��޸Џj��q���x���/��|�f�Z�fw`"�01F���ْ�_g����8�߯������,�G>+4��˼<�4����r���7�.����wV�HI	���i�h����^����.ו)5N��(�sE�"�*{����ӫ��gX�4��/<N��a���=|��i��k������6�����������X���\�}�-yYI�tc�u	�����*�Ⴝ⽞��^���}0�ט,� MA��H-���9�m�S��%D��z�<��[���h�칻�9S�W�m#L1;�Nk4h�c�z�C���2(K�
X������ft*�s%�v@��d��:��#�c�I1�Y��Q��^���Ok�-���~og"�E��%�e�d��"�q۱�E�[�ڭ��,&u�p�F������cɺ�x��Al>���cN4��dݹ-x��G���#a��������y�HB1�+�B`�������i�#Z%�ظWoJn���\�P锥�;ZY��fhb���=���q���[�p��t�!�;nnBM�C��r���u�Ķ��H��C,&
aѵ5�p�ΐ��0[�*�]m�r!���r�1�ŵ��[M�9�r��\�a;�{�?����n����7W	;���S��n��߇{Q�KC����9�ؤw='o��R=�����-ģ02�U;���*L�=ycr.�7��Ǚ��n�y���N{�h�Tb��z�k�Q�N��U�|���^�w�^�x�4��m�����.)˯�K���I�t�x̪Tc���q����+x��'��F��5-v�˳�>u{����W2�N��������Y�aZ�}��yk��k�M��k6e>}�"E�c����5u�k�:���W�p���O:��x�Gt��)�P.ȑ�yMneT����ó�鞢�dʛ��z��u�}㽉��.��z�]�������^���Օj���/��n�#�"��nipU�M��ó=. ����0:�BЖk����06l�����g���?5tR�-z>���=�����hľ�~��|�,��T!,E<��-WG�2o_���rfae�,��	���a�^�=��U���i�~ש��JQ�-ѻPU�k��L�		v�[��Hp#yQ:GQ��1n�s����E�y���c0-���3��ri���?Ntn�Qn5�����ʃ�{ЛY�u����>�{z��1ƵD~�.�/UY��|�v��f����t���m�k&j�p���>˄R�z�o������}�����y��e�M&�%δ��0�{|�Y�0�~� ������Oy��A���n��Uv�e������́���%��~�1����`�bX{ȫP����m��P螐-�������?!�%�w	����~
KKn��jou�K)�y�@޼��bR�����GX��4�:����ˣ�Z�ٵ��^i���1�f�,��d��+�<��W?{�����f�!�}�;3Yx0�ԯ��{7��{��yH6�N�Y�.��q�(?w��US�VfO)::�k�/c��$��jrR�4���ݛ73�x���k�[��]5�{���#2&SBR:����a��sC=�RO7/���C�?R����5�N,oC�*�(fm���[�˧-i�X�v*�C1�͜��u��j�W�Y����ʹ5��q���S�PWT���ʣ��'�#���x&&]b��]m������Z��;�Yu���X�������_Y�+|�;�{-�2�.(Y�{O���Ư�FT�5𶚐��&�N+�[��T�G+k]+���ֆ�s���7<k���:CJCUf��/<yg���4�����?u��y-1��Q6Υ6�l�[g1� g[o2��d2���صJ�Gb�-�$Q{����(X�]nUv����-�k�^%�!��ʍq�`[�,٩o;��Uj#w���6�S�]���(���1I�ͩ�R¼D2ͷ�X��qSݳ�����QFf���N�m�QӋ�շ�;���$���SJA�������{]�؉c$�`Y�ۣ 1�
��>ǜ�������nf��UβA%UU�w���2���<#�,C���NX��_;��Ǵ�q����U{�_;�C����R���R�--X���y�4E��MN-�ke]&��{ӹ�@�d�5�]��}h������x�ٛ� �՝���&��4ؗ
=|�����s��r|���|+e>�lA�b�<ʺ�[��ym|q���.��,�A�zQ#����,�|�:h6b��3�괝V�[6x�,��YSX;jF!�ݱ=�gq������)��Z6DU���,��[��̵�X�y��,B�o���:8iE���X�y�:�s��'*A������*I�lD�����,���齖d�=~˖��	��_��D�����8�����̫������H�[@�*�Que;�I� Z.Df)�Lc)���*ӘT�ވ'gq�]�V| �S�۪ɦF����u'n͂��_yﾟ��`Zʌ��'T�}�:�|a��z�!��$�ݝ�qx)�{K-r��3�����Bw��`ǔ3tTʐ�:�|�q�N8�)����ݭ9����hPy������qP��z	�9��,�W�<x��jXۦn�7���Udc�^����Ә߷si!4��բ�j-_	�^��}��f����y���G� ���ނ0٤����t�,8r)L�@M����s��*N;wk��]ot�vp����ƭi=[�98�<�[��n��Iz9��u���r�D`w��=�j�l��&�խv�"�f����;U�:.�}��N۞�r#��ڴ��u�;qN�5u�C[3��n�yQ�J����U���B0;������T	�@'��;cmm�i�:�^@�=�t�L�:��ͮ��2��X�n��]�gK�'	�ܽ��1�["=F���:7��y�l!Ha�]j�\(}�7���:��ea��C�z+��<����[��(z���d]i���bXS��y�Q����)�J"N��}����y{�b�`,A4�^��_l'�������\�A��A�o�]\��ę����{�}ւD�U;�Y�)	^\�sϰ�ͭ�y��������0��Ƴ/ӸR��,��JQ��]^RG\[�v`�&8�qH�|���C]�dI+����y�o�:!b$��~���_^��l���_���ܑ1��?}��%�K��<���������Tڼ������0�R��º�����ed`��&� (}ުv��-M�sS�uj`e�M>��SƉStL�]v^q��rΖ�'Rx݄Pሷ]��s�3�!f'���K��EH%<��>~ꪥ�!Wힲ��v���}9���} E4��������s���A�Tp�!��Zr�e��}Y��ֱ����uB��!�����Ճ+H@�M߰�����{���kK2+y�7��Ek��h�|�;r�PB�ۡgV��y�<�x%�]rhY\�>Ǫ��R�'F���خ�wgi[C��;�Ӊ1�B�QI���j�R�f��EH���g�y^,W��g�>�Jض�;<_mé���Վ��ƞ��Vd�+!QSw�_c���m��O�y����l|^�V�T�J⓭��l�W�&��F�y6^v�;�
��e�������&)
��*�1ow���l��X��Ze����<>t�t���t��eH��?X�K�A�efk�,�k�C���������d�Y���a���k�ۦ��{q�}�44@�RQ�x[���qͳ���mJ�k����m����;�ƀ��K�-�z�F�=���t�-W��w�<fV�JF�p0�0�ӏ0��|Ws��B�M����{xW��z���#Q�F���@��v�{K���]�|6�:j{�:�}�ˇ�3�0܄2�d�^p��Y����5����Җ�BJ�����jy�woJ٩g��,��Jזzڈ�DӔ�e�ҥxa5�@�ifk*³
դ�m[֭�cn������Z��Є	�ʏVh�k�v���e����\I��n��o�x��»��vv�T�;�t|�*͊Y�����}��8
q�ϱO7`��jWm��s:�p9��2��6�N]�jv�ܮ:�Ӕi���y���'�{N$|��m"���d�?5y��7п	ni�-b���I�-z�����9]�Z�����ӥ�����c��n� �g]���貪@t7g��v��/z�#e�QY˽aj(-l�S�,���Wz��(�oMn��K�N�@Ep �)����\�s��X729]/��y�X삝�펜쀅��&���-
����|�v[��2�N�v=g�T؏���ikj��iAJ$e�31	���l�vq蝷ms;H<�[�'���[�U��o�X��'�wN#��	Ӧ	���	Q��c����,��{1*f^���{}F%��n�#���S��.��u�#j�س��E���_�&˗���A�C~A�6���"V9+��������7Nf��ٕ�ς�F��T,{�,#��գnbd;b���٩���s�G|wYۍK�Z�*z�6��J�݂��h�{�s������=�&$3fhs��Pz�o��,��Cw���tŮ���q��IAn�W��w}��Q��/�D�S���;8Zi,eH��l�-���TbW�����X�r+���5�	V8��q��&�s��9{���'ㆎ���Ƿ8yH�l�Kp�����&fSiٞ�ʿI��<H����s�@�y][�Ƿ�(�96�l�!z����k�Z�[=�a�.W5��̫ ��
����>�O!j��#zr�4�T������;��Ѫ����$�n�\�����[g������>;+mPQ ����ZJ�W�:-,�1�WWX��̍LC`sA���0kXĕ�飃l��=|)��tuW-W*��.�j���<���_�A�9uЦ�ͦ%�����?O:kZ����x!�'"LHX�ȝ�jfN�wz�w�^y:v�jR���H�ŁUTR�<��>[�]FV���)�e��!,F�;���a�\NDcRI	A�!�k_";<�nٖ��̢�{�7�;TR�䒮���V(����{v|�mw�6���EN�۵�!���,��%D��J0+��l����<�S}^ԂoA������X��o���F�� Hj���w���G߹�_5�N����s�W�o�����U���k,$!.v�ls����MѼ���u2���Z����)�7�M��]�N�Y��ci4�%I
�GWy:��xu���&'�C�wm��2UX��Ř�����;N�ln&����G�*Z����ћh^���+v�V%���O�]��g[�����Ј�����W�,ˬ3H�TU�~=q3���R�k��ȫ�(�>��|�w�ԟ��#���E�K^��s}W����S���k,p�������r�����AV�N�߫uC9s�l��n��yo7g5��ݿ-�	�v�Ubʮ>���u��䁗-�-�v���o�=��ΙY�N�<Au����.ʨ�K���b6����m2-){��o�w�M������ͅ1tʣ`�L�n��Oލ�����3�{b!�ܕ�n��{��[�g�(�+S���&�߈P����uo=Ƕº���W� �5�q0���#n?7+��C���וֹ�D��h��%��n������33��;TS�9ċ��f�$ʛ���C"�&��$
�Y��2�coZ"��@�ܟ �v����
w�Eέ��T|K]"�z�Z�YJu��]w�o������l�,h0�l&t^��Y�^��B]�Q�P�����'m��QX�rŪ4��)3�i�5�t�l3ZJъ�-j��Hi��#4�\��F��]6�n�.6�`ܯ&9@7v��s�+�w�6ϐ�xힹ��л��a~�'d���N���#�pW����aJ�`[cJͥ�[�1g�a��D�մ;Gg=ƞ0���3�oBr�h�z��Q:p�:�����=���'.�̠W��k�Vظ�=�9���n^�4�%e&(�)��P���Uu�}��@�Ǟ�U|$؉�6s��ͷ�W���8V%�<���~�<��� M�5vq ��ȕ���+%߻+�9�spP��\j�_��T�^܈xK▒��>��LV���g+�<y3�V��w�.�w� �0�`;6�=�������ϣ�X�|�lr��(�{d�+o
����Y�_6��ӫY��l���MO��궵nT��A?~;�a�z{a�Z��w|&.u�J��\T.�׷X�Y��ݏ3�I.2�g{cy�j�Z���*]ٴ�����m]~~��Q)n�duYW�Z>[�l�{�u��{d/��{7y�^(��5�:�U]�R{��k1��Z�.���^b��K��m))vj�+\���}���-�mp��X�J}�mpwE��/���"�A6;����skS��c�_t�����,�c���3�����CM�b��th��ˋsr��`��H�����R̠D�a��4w!��zsQ�J���ˊ�{ï�Q&���������P����VC/s��f�aCU�s�{�v ��t}7��~Ai����5�z�1e���|��b0`��,mD1A��M���w�{qLnaF��U�u��O��}�ҍ��,׽_�f}�v%�V�a��{�G��W>�Ore��:����p���k��f�7��_zv�I��׆�=B�4��B�Ӻ�$��/��S�r�Z��$e2d�+�L�Rv1G��?b~�[���_C[[�ޗ���S�Aƻk�\����qru�S�Jp��Ympˈ��˛.0�Z��xq�|�a�ϲ�]��j�WG8��R.�i��_;O�Uڬά���;��uc����8�.��V�K|��7Y鹛yu]�Lu��%�f7q$T��b��6�n󕂪�F곗���wW�7�g��9���5�p���X�_�4�/�b�L�9�@�Y��b*E�,O]M��+���Ƈ�Q�rb��X6��i'f���t"����)��6T�h��W�1�+�����HR����v&��8oL)�[�'u�{��9���܉5�p�M�����^4�,_�=�ӊF�P4�r��Aխ����}f�L�ϩo�{����ݧ�n�q��tNuv�Myya�u7�Ew����b&�8Qͩ���^e��r��8ԑ�T���[�uݾY��*��)��>:�R�i�S,WN=�|g\�}�S��j��_�]=�y������Х47 �7#*�Ԧ���͙H,�g��9�m7�<]��^U])xEd��ݣs��ӧ�
�8��e��ooM�}ޒI����v�n��u�%�э(=(�4
p��P�JR�cw�{0���LvrJ����K��DٿzW���N�]F\]j3趆�%tU7�ʌmw���m-��lE"F8nŧEq3�e�j���Eq��6�b��=|YK�.�,~�锵������)�[�}�(�B��5#�i5�N��{�qO�i�Όi̮�p��=�Ÿ(�MOz0�1zΝ�M�o�U�I�чs>Ԃ��z1ݽ�W��ש�ȥ�ؙqi�WI��SW�Ci��M����
r�����$=�{�/�z�f3�Al������|VS�:0���d
��)?u'37��Ȫ����fq��z� ]���Y�[��9����C�S]lUv���pX8cCh[1+t�%�����X�4u�Itm�7��g�����\U�|c��ZG;�D�<�]}���M���B�`E�*6Q���s������-��G.A!~��m%��ݫ�m���t��b��G���o%]Kb^̶l#��^����׃���Ȋ��s(M�;�׽Ǯ����R(�M� ���:�˩Wrs�.�����wz����pw]^��9�C�y��r�=��W�� ��1% �"�^�U��PCվ�{}K"9Vh���+ș�T�[�nq�Ɗ����7�;��>߱c���s��uN�����.�EK�1�r������h�^7+�� �en�O&�w�_��>B����%byx�|P�{R�+ˊbr���5�+M�+6%T{ƃ��Ss�֙������8�Fz��X
�j�u��w6���c�D�9�L���=�y�������EK�.�]>�bюA�G��qvn�`�jֵk1���C,ɵ������c�%�e�n�lm�c$�B�ʶ���p@!�cD��Au\�I��]7�[��kT��N10��.[*��"��EYI��1�3i�A6�k��[�3+t�Y[e,�^�<��h(�c�>��ŝ�;{B ޻-��c�[l����&�!1��5���;1M��`A�sa�ɦs�H⮚LF$*��	m���F

9	����O��ʻ���j���6����]}7��j�ۆ��$<��F�p�f׎Vx�u�r�S�q���8�0?���
��*uWD��_�d�M������� ez�f篽ۚz�7f�s�Q���+��w��dq�i����ǲ/��[ x��#�ZY�z�Kaʲ����OHk����4�z���b��T����`j5q\)����K�+w�MY�Ǎy�U=��h�F	'��g?�[m�*�gq�<��1]�0'SO����Ũ��Js �\HC���^V�j�����Z�����Wm;�z�oU�x��mq�^�=B�)��S����3G�<x���u?@��гMAQ���U�if��L컗g���f�.��F�X����.3@S`�%��$i���oI2�R�ޯX�׌�O���	#�ޱO;SҶ�
%�Veܡ�n�pSw��b!�؊.�q��|V�+�m���W��O.|6�S�j��[z��7Q%y��[�8��A���ە;2'g0��3I^byڮ���a��nTW���p�4׷,�+M��g���a���w9��g��VsRlls�U
b' $Y�A0�K�N�}�m��3Ι y�e
���xśLً��.LY�6=�>��c��)v���J1���38>޳^�!�]^p����%�����|�Na��]����D}m���J��l�˥n��6��1e!#��ނ&]uJ�m�92V��0V涢7Ti�y�/kb�^5�"�M��B�k�*�[�y���z�ǿ�'�;B�́�rA6u^�������/��`֒�n�W�[K1abF���Q�>����y�L��a�����1's�+c}��=�U��>
÷O){�g�{i:�W�(�ǃ��z����U��)K>�N���^���;u*��_�3=X�|dU6��%һ�jL��q>�E�u>(�&IRC�}R�^���T����f{�5T�ӧ�w^�7U��3r���jq����Xق��4Ҭs(,#1��{FVi��(�5�K�iS����$e%�@���j�"��#kw�;_z���vy�bU��{Q�{_Z^�!4��޼ �22����}��Ϻ�Pc	z��k���K�r����������Dti�Q����ן�fK��S�U��%Á �8�jѻ��
��.Y���,�16V�l�[[h��g�} ��^.^�}Ŋ��܅[���B���WC�{4�kq-�U���Q&����L�(��Mv�an��e��yֱݱ��c���>�u�y;�>=W-�u�s���.�{��l�=� 7��f_`�^����Y�Ø�,��lHjG�^}�޻���Ղ�|�J:)!�E���Y�*�ˊ�8��������á�nuU�礻�Qi��%��E8�,�u������}ޠ{���e����ϐݓ(x{���/_�2���J�y�U':�TIƔ�M�Z��W���ɯ�;�/��
}�&k�N����η`�R�	4���>����:Q������W��lv�'a}@�ɣ��쵑Q��m4�V@;����^KVN9��a�\�3C���&��̡tę�t����Y�Lf�w���jȒ�R'�i�>=���;��F�z��%��>�O���@3;}l�����z8�Z����}<2�xg����H���%���9�����v�6]6s�N��wm����S�5�6ؖ�b-�-����:���Kץ"t�/N<�/{��.G_��V_n��S)���d[RF��G�q�e�,�$d�چI��O�bݺ�i�*�����8��uc+��nȩ�+�w��dTW���m����Ekd����=��I��w�����w���%86�}����YW\%/q�Ib�ɋL��X$�ʗ�;�7f��݈����J�y:��)(�Ѥw���
�Ju��F�皮ԓZ��{(�>4��!�}�GM��AA�m.��ް�;�����}>�4���fFӆEg�8���S�]aMz�]8�.3��N��w~7R���1�K5F�c�Suү�/|fY}�� E4~�r���c�{�e�����:�q��®�*���E�K�⌳u�)Xx5Q�z�Tu�:����"Ng�y�̔�p��ﻔXn�в��!���y�t���KO5N|v��&���Uz ����9�[���������8�Ip���KC)�z=�ƥ�(��*�V��\q�]ht�OT�j@`�#?����Z�(���Y��+��u�p�w[���[ǩO�q.-"�;l��2CV����\�`�X��P�v%q�l��|*�E����5Rː�QI�:n��t������� �Z���Ij })̺��].P�e����x�AN�U��l溥hNkronj��Y8�ȋ�r�Ս�Tc��!��t��n`�)i0�:cMl�s_6�Z�������
���q>Xd.���g����6���QQ)���y�؛��ާ��^�I�S�2�f�t"�
��v!�5��#4�$G�wރ����VW8Êō6X5Rl����m�~2�c�P�1fm�X}�]Yq���ñ�n�v�'X��G@Y[�*"�"�i�}��ll+2f��n�ީ�%wt���{�Pi��Y��%�T3f���[��I��K*�`���>VN���KZ:��C-��k7X7(�bEkLz�.wk8��B�X;�C��a�`8�]51�����Ѡ:9.��:1�/d��L\�ν�M����;]��������W�&�������w�,Ǖ/I��3�B�	����6�h1������v�ԇ�?w���펓eJ�j�Ѱ�נٱ`ڙ;s�1���G4�(�*KZ@2�9;!ŧ�����rXM�����όt�\ݵ�5�ق(���\���-7������܀�^ѸZK�[/m����t���3�Wn�=��=���I;Klu�`斃p8��I̤<k=ܺ���y��uJDz����rkS!v�b@�w,l˗i�<�'��:�9��xiu��w���ڐYwgmCpz���	��UOK���f��<U�c���Q��ێ��\Bf:�+Uyl֐sp�I�qM�ci����<^'��g�F��d9�>�j�w���S��+@6��M�ȑ�.��6���y4��I�>�y�޹��c�]�.w��4���$�:��nV<ق�m̢(t\gL�V緌����Yc+�b��u�8w7[���ZY[��v\v��㶝�`D0nŬ�ĸL�IE fM�[Y������[!�9��##��v�%�3��÷�>՞�bm�C��W�÷V�gF���-��ωm�g��%�v��`йh����oK�T�V2�\f�����^,�n83ܭ�mV�"m�9��^W����V@,���j啕�8�h;C��R/�)լZ��#�`}�g�(yƞ9"�:Ml\g��J��t����Kfiv8�b"FK���!�Ea���B㣬��H�H	���2V:�P0�P�cP^=]�囦X٦]u%����2s�=j�!���R�U�%���eU�]�V�/4d���
��볣��7mu���C�xaC�n��[q��zt*g���BK+�1��&.�p��3�:�e�/c5U/8!s���lqA��lY_u�
�����WL��Nvչn4L��x'd�^���3I۱�ۇ���^N�z�ٷq��s�Nz\Q�k�`L�YG����.#j�6ա4�u���+��g<�#�ǺV8�س��n�3a��Z��Ʒf�.�����9�a��, ��f�mL��j�m�#˥��^WD˩�XJ+�B���3��a99�v�z<Ti�vZvɢf�N���+)����'"s��5����wm'pA��t�l���ܼ6����:f%ᐗ.����4�&��9I��յ��i&\c��fv��s�e��cla�80��9cc�j�p�)�,V61)*�ι�)����Z�1�ں�Ηa���9���[s�^��Y�1�t&��(��-�UGl�T�٢��v��r���p�� p��ޘ������H}	�A>������lw��㛔�(	�G}~ڌ�#/�y+�X�:�4��I��08`q�=�.�~=����{e�~���%��Y�#�W�-�G\�{������oʔ�瀦������j��C�=�V��h�")��-�<���EJ��:�J=�����w��,uI�v��ΝJ*5y��*��×F���b�Ya�e
HnՒ�ݭ�4��������JSG���~�z�R���~�{f��u�z�94P���~�P5Ys2�T�w}>G���䶖�ڏ2��"<�����~񪺺�;`���8��+�N�mz�s>�p�U�CN��~�����L���	,�n��l�n��^L�U�t[[�K(�]bR���.��f	l�\�RQ�i^Rok�C��G����^;�U^�ɼ��!s��1L>[۾��NƋ;���0����Qת9���(��>�mm��Q�Fް#��ʽ�Vc�67w�:C�;�����󃢺Б�FS��Uv��Q�[��N���+�ث1^�FG
'i�ˣ\��7NK�����j�e������<<�M����۠��c~=��e{S��7D�$�#� �n8%S��2����;��������}gȆ|ӵ�]�X��տx�{�Z��O��1k�[~�~�¢L���#��W鲰T�jj]^��j��Y�eyN����f:ΔMk�T#��}TJ#k4�K�ʗ���E�:�hv�m���N+��,-�x{
Dnp�@���Q��b���~{��Ɛ������<��Z�{�U.�E	�}��.�R+�`�6�	������4ܩ���lBC��=+n�$�b�\��2��H ߽:ӫ}Z9�=�b���}�+]yS{k����[q�|Ͳ�I�;9�y�l��uB�'�F�h�(�}��c� ��ћ;:��a�P"���{�fk5�6����N����^ܿQ��^-���W���(��$�O���ǹ�k���\�'?v�:;��� 弖Gz�y,�a"��~6"���e����/m1�6@E��C̸�LEI�\=Ef���l�VGY�ꭶmW( ��B_QܫYإ�9�@�����i{�oW3qx��f�$����<6��F�7��Q�>u��A6gu�i`=':���e�x�����z��y���&<wXB}��6Uc���R�vpah�1��d
8r�����A��UR�ʛNm�W\�޷��5Rޭ�n>�{�ڵ|�ݾ�L�ͯ���?m�ϧ�$�+��ڼ,b�0�s2�d����`����W�A�ۘQ��JH;B�N�*�e�%�����=��O�x��_!sSw%1��9��2�ʨ�ci�BB�0�FG$}������{)����N��4��/RC�MOM��o)w�=���+Q&�w�f�-m5�%g7۾Ӿ)��J��XXqĢ�'>EH����+|s3�U��(�e=�m�.zQ�rjMY��ڼ�v=[��l;&86� ��N�±X���}���(�qp�cj��kr�w����{(�"+w�^)��b���v�Xݞ]�i�4T��u^���.�GL����Ò���ͬhf���oos���	v�*�ҧ4j����w}�%��A�ﭝ�9�x��3���ܷ"K�\���t�~:î����G��,�{����A���j�.�=��/q+���|�at��I��fmOW�]~�E��B�*G��2n��B5�J][Mg���@,[��w;k/bl�mv3��e�˄�\}�_��t��+��{V|�v%{�=�T�I�ژ��5]�{'1�/Ӷy�N@�+�Y�,��6��"�h�Qr&�JG��}uvm��g؍q޺3�Q�t�HC�-{_�G�u���R��I�5�gU%������C{*�V�b�wL�8�q&ĔqP���r��|�죓6��sS���4�l���ע���1)w����:x�VfC:� ���HrD]�����tD�iѩ�)��5�εuǎ��r�|�<��ΔkԹ�3ܪvSZ����n�{�8 �7$�$�nI����rRWOs�L���U�{ٻ��۾�K�.�uBt�{{���A��t����b���(�r�.x����'��͎)9���MS�{�{<vU�F�[�C
Kw��5^�������xu��}ܫ�����7I��������]�{?.�n&�0cėc��2�v�j;LR�A��΀y��,Xی=wy����Oj��ㄍ^�
��c;th�Q�w;r��1��E�*v�����d��3��ۗ���U�l1հ#��L����7=�n�2H`�,LT�&���s�[������:w\�#o^����;zDڻ�^��7=-j���դc�;��72���?m�@}��*��0���f��k���r�k%�v�$��[�)���ff�3(�"�3	�U��A������^�w�����w��ϹV,e���ً*2:�gLӻz���qN�tB���0���M$MK5W��Zՠ��������{XSE���K��#������Xqߖ��X�7�GaP��)���*�r=�?<,���t�yC����ԭKb:�7y��V8��f�a`Hv��g|�n�^�c{�u�=*E$�9,�'$���=ΧP��I�<s�/&��X&M�o�V��3��*Utj�����GIЌ[�x�se�����"t9ww�/���(�l���-�׷7 ۾�\Oxh��שW�uY�7{lś�ba�'oI�e�W;o�W_��������
��/B<D �A���.��e�m��9�&.�{:���^	ch�����0�U����.�;�N����=^��>��9-�ηF>����1�d5�9,�e�CKag�
#�fǧ�m&^�6�R7D[2�&9!���+}V��w|��j��H�f���z�=�Q�yd;����!hS#�C��k�G���$�q�GXtn�Qr�޴.���#�,��񯘓�O]	�E<��X���:��؝�{hz�k�i�o5����>��/X���}b��}��|��U�{�(���$%��e5"2I_x��]b����J���!,$}�|z򷺅c���P�K;��� ��K�o�����Yhߘ�n�����4h�p�8�a�>�9�E�k�2eW<�*�����yy�mg~ɩѢ���C��<E(X��X躽�^!s~�=�6��h�Vo��w�j�j@��6LLF�9�����tD�6a�+W債a�� Ӑ8C�sSm9�j�k�F�$���B��WJ�+����	]ء�u���iBA§c��u�+�߅e	w�7���ñ�brݞ� �ѷ���%̧[s�k���Q�f��ö���k���j��oOӝ}iYv�kyPö��u(��7�Rw���U�q�uZt}�y����M��(��y�^�dM9L�)�׼о�>��B�����O���C^�}�x�(lu�~4ƹ	��r���}潕~�E�K7�[�`��hKɽ��'�/pf"�1�7��w뼲U�۵�t�$^�I��f
6���\+5�R�׬V���^�X����'Wv�3/jD��E�$G���2�nP
�ûHj4��Y��ݳϛ���Rb,kn��B�Z�����Ȑ��՞x'�[�g�w��Z��� ��.�Ń�%�IH�p�O�{�{H$9&S��������sf	'��*�u�pN�w�
��8��.@����Z��G�,�����GP�$E�n9&h��20�Uʇ~Y���2o�S�T!yML���M�TfueJa�M�����_v-�l��ЩT~�sw�+��w�;�k�eص�4m�e�8���Y�^k2bkn&��8�s`�����5��v�3h�G	$z�υ�8����6pԫ�f���}�$<�Ρd_{�j�Ŏ=:x�lX���i��l*�p�37F�ۺW�>���}�a��/�w��w������Y��Jb�-~%@���;<���#��Ɖ�	=�*���Y��!Z��V6�g�"�bvz���y�H�g�T0���Б�$9�.Q�m���_,|k�<�U]���<�5����e���n��Z6C�u��_s�� ��û:��~�)M]LM��E���2�-����x?��N�Xl��G���Sq/
�qU�>�]�,�΅]�|�O�(+�h�^'�m;�/^���oƖO������vX
��֙�n)�q���r�]ݎ.xV�!\������R[����?r�-|�H��%}{3ړ�����	*D��A��5#����f����Y�*�|#���ߧoVJ��~�x��>�I$%��UW5@[A9'�<�в]i�'������-Њ��V3^,��S���a����7)�8�:�X�Sl�9�`&��d��aQ.����^�b�/�˱�]XUYN�J�ԌMwc8��O9���x���]���&��Ww�(}C�q]�W�EF9��n���{�,����]7+�z�Z���?S�s��N���I�M��f���u�U�v%�/ӵЧ�<���-3��xNϒG��`R�i4���Y=��V�-�r8O?<ڙ���^��53^ܝ�+�*ܣ]�7U��A�K2���ǽ Zk��4�m33QG�ݔ�w���N����8�)����Fס i�����DVk���]�R�M��c�����G��:�)���y�Ru7}���Z5��� ��T�' ��:���Yힼ�cS�#���ֺ}rJ�c����[��E����F���RB�Օ�3��4^�Q�N��̽Ἡ��[��Y4�)�恈�oA���]�"ଈl)�x3 C��m����ś�.��/lUKD�,�x&;�F����tb��{�V��R1&m6��i^0��n:X�m�*�f:�{gl�v�Z�j�н����츱* �ݳ]�����lq<sSּ�x�/������!H�%&�¸V���Ƣb�WYKh�c"���3l�qo�ه�kz��L�D׃�㇒C��Ý묪w'/7p�&&�H�1�dS��Ypn�.f�8�a���D-�R̰�'^�۳^�ɹ/W"�G:�FX�#6]ͬ�΀����0����M�q�v�.1�[N|�����E�`���g�����{Vվ�#+2U�=~i�fp�����Π�V��S���M�Ls.�mK�
uFh���v����V����D�}��
�U��ڧ/[G�b�>F��,VR�4:��^�Oz��9MLaN�v��E���.���ʐgzU�4}��3��y�$�m�u��p7EZ��v�-���r������y203>�,���R23S�r3d���~�<�c"�g^�w�x�v�J��d ��W�K�l��Qk��r�]f���[&]N��.�wOui/��?}<~I��X�1�U�����",�w"��[���H�	q[��7�yu���ܓ��N���Op�5�"�+�3��;1蔑�r��Ds���>���."�maV�5���s.��Q5�XMI��GB��/^��(����$�����3#�~V�G�Q
S/�zk�!i@3v��W�Nyi��ws4bD������*��]���`��f{�) .}
2�q���u�������X�⺽)"��3�z��\�9�}<���2����oS��w�ԥM�1A���E�\�|��>\Τ����t��*=�@M�����/�w/������ 3���A>]�%���>�muq����-]^���!�B%�����yHgj��N�5�S�1轛>�h��#��諈�GU�n��+�x�
4ׯ���l]�> B��zk�zde�t�F�G^U�����{C�,�ߝ���s���y�6[v2�(���b��o&�Og���s�V�"R%DsS1�e�싻�.e�"�e�V/��_C��.�d�úvT����*���js�W]K�/���w�λQښ�$c�y�ד�[��+��TP�^�p��p�4�-L��gbOc�-�篴�\z�$�)zo5��}��۱s��\/�����MKي*�"V��i����g�ҡRY��ĳ8k�vΤb˕ŋ��b�e4k]Kp��lfm8���,a*���{���iN�$����^�&�I��P�@I�9��+ZC9ǂ��dȂ����qq�f��_��Ŏ�>iP��"�nn�wQY���b#�Z}[���^����lq�:�#H���Un�^�K�[�p�����2߯({9�IYB�!NN�X(fB�l�UY�,��|��JD���|ɴ�ZZp+��S�U�K�He����z����tꂓuE�Ed*���OSR��V����ZQ0�b]��U���$.�%�g�]�wysA�^^�gs��U	���;mm嫣��i ��N�ay����Y�+k�u;{r�:[��e�����u�5� ��o*kv�N	�������y��3jR�8N8��I\��9֮�����rɝc�>OJ[�<3��v��<	�-Vy��R#��X�Х�Z2^�'i�����W�����z�yZ�������^���
(�Ju��(i-2�7�V\�g#:�r��-8�]�痬�2!@����:�.�ܷO�qf��鎻8Ωs�tc�*�V�6�-a`51$}��	�Wtr�Oް��+/m͒RA�r=�G2�;�~���BK5�#Q`�r]X���"��n�����L�Z�Z�v
��"R��\�Ы�7Z��>�NY��}�d�;�u菔L[����V�n泲�7�;Q����G�IMްMe�Ú%�V���[,��6��X~;)��[LI�3�3��>�0��˫�_G��żB��3�� &����g.4�n#���˹��rm�/$3�y��}n�w�:�Gke{`ٕKѓ��0��h*�zH4�Z�z����b��UG�I��ЧlzX4jh��f��1�wS��G�!W�)񛸗��^��d���:���9�=��人��yt����W��&.f�j��c���b��E沷���q[�t3��`�C;ޘ�)p�W$�@�̲�E��M�`���R�WU��oz��|�X�mӾ�ͷ�k�f�e�����n[�]}Y�����=�;�?	���x޵�ʋ�>H��X��}UdV4�����<�;ي��2&��\��������7T���6��i��^S>��q�Y�����Y��?}+)�|[��.�g�DԅGUH�Y֢���w���י�wk�Q�"��w��qW\*#גȊژ�{��J�<kbZұ`���tZ.�ߋJ�㢎�-��-zO4�ki_�pInn�8�4��-$P��$�'�����9��U7.iZKd*�U��S���4/m{f�5�u±%Z�$�;��\��{9�}��I��I�"�I{;�W�皘'�d���dcW!$�f+r�0��j����Rp�S9�K�^����o���������B2���/U^y��;�����7Fʑ����ƴ�"�h���O�����,�J�%�]��|"9�.	^5DH���{Ԯ!-!'ƶ�Y
ûE`�&G՚Z��s��rv1_��G
I��
˦��=6�KPĒ�qP��l��F��9�L�I K�Q3T��#�&(T*�Jȅ�*~�WH�=^�c�%�[�L��{�VDQ#�.����FF�/��0�P���IG={u��r��S-.����^��WUɅ�s�<�^ƧOV�E�K�v�KK�ۜ;�$����˚���R�D�X�
	+���Efx����E+�YDX�/;���(�jH@��3�v�cN�Tǧr˄��m� �q��{٪�ä1%}��B�����O����,F�4�3���x�+^j,������RW��Os�N�tP��D��%$B�_�Zd%�LR%�"�f0�X�4Iw��+�3pQ$*ڿ����e=������k]�����W�w�n��J{�fjDJ�\Iq�ͨ{�\����J�;ӣ{%�+f���Iv
��/1b����J�[�ND}��|.l�B词%d$��
�|{�A#�s���9��>�����Jn�iE	-#��y�D���S)C!x�T�, 
�=|���u������t�
#H袥���M����kUr��!h��
$�RG��םƢ,Q���%�� Q~��o�ڙ��i-��-QBMM��ݶ���S���5�bh�qJ��Gk3���!0ܮ�k�U��n����ܞ�N�p�rmN����-�ME�O��X1%��"E�4�Jk��H!+"#HJ[��o|���w=>=؉F�{�,F����o�B�N��DI+}<���y�ӿM�^\̄�TT�^NȎ�Dm��XB�.���q\A��Z���5�Iԣ�(�E
H
��̪�ٜ��zT���-%�Rb�-���:��(਄��b�%���Mi�Z$�缝GD��I��l�u[9|��o"�]V�j� ι:��TiX�J@�%bTBZG���K�e&�T+��c�H0��}����봢Ί<B�Aӫ=��w5�A���%�"3�%��ٸ�fV�Bd{L�V(V(��{��%�J�Չ*����	t�����|�)��i����ȅ�Dۏ7
ĕ�|��{��v#Hҥ����K�X(
��
{���{.mG�T���	I-�Ĥ��^緅�I!){����XB�d������a�dGf��}��+� I1i	I �o{�r���RU*r�Dh���*!I �������q8A��It��\�!uc�G.lǞ�??�U��de���=Y|.8,�S��%"�%=p��^;Q{1D���IP�J�4��Y���O��pQ�]4����0������W���2}�)9�u>���gff�+��Ou��Lm�艱X�_uj9M�y��R�w�^�~ךY��>�n�~�����e���.���M�9ݺn��i�뱴m6�Ff`���g�!E����v۠�e�=��c,ط7���1��27:�dLh�Y���8x��XQ��&X�����3cDm	s����B`�tW���U/im��:7ŷ\09�tVܠ:�j�>ҡ�W>2#��1��a8�b���=C�]vi-�+	�-#+�U�����4
mȝV�W
\j�D5�l�F1�9B�6N�^�{�}��s4=n���vܔ���� �N-���*J�J����BdC,m�](�������ظ%�1B�*]"[YCI�w��kP��<�D�J,�%^ǜ-H�����eO���^��%d1D�'	�{��`�Dd�r�^"
��"��N�MB�3P�nFw9מ�\��{xYΆ��H����mk�E�\ɖ��_��v�Ud���V.�Np�L���qy�"�Ge�K�H��vmQ����y��B�J+��.'��Q�G��t�g}|;��u�����s���
jh���Qw����ת�#g�࢈��z�\�j$�������丿O+�x�+y7��i	m�Rs�~�dޫ͈��p�8�;e�XD&G���ip�B�%�f�K��+(d%"�R�{g:��<���c#s]���/���J�T"������y��a/��u����צ�H�.
��
�sF	H������
��fRE�N�aG}�nҪ�j"EH�k�w�1_U09 ���^�0��!Z�J[mP�GD�.2�WU0UB��S�USFD��p��EkQ"���⸍"�u� ���s6+Yؙ������2�n��E�9�
0��Ԋm�
o���O�u�K�����=6��к�� S�#4:�Z_7^��[�q����tm�z.,���uh���L ������i�U��3�&�iԋ���O�=��ag�5���c��w	x�yҵc��D]8�1+���P��2DP�/�I
+�+۞/���ڝ�;�i�+��d*=���Y�Lp���7�Zi
�P�%$���tyuP�eT�榦�%�L��A��E�s�v>���������:��F� Ѝ�X!���x֤�'�d;��r*y���lW�]cn�ǴpF����h�ۏ�����.n����а�6�|k*�F�ޘ����Y �K�T�h�>�M�d^��+*�0�B�B�(w~���!i�{����S�l{��8��x�!Y?��!��ʎb��s� �N�ܒ�$%#�Z]�m���r��p�%b^"H�/3������Ĺ~�sU���~�H�/�RW�o��\#��)�b�M8K�k��׭5oDICR&u{�����efB�3os��5��i��E��\�hbu\����H�UnJ��qH\BV%$ �~��^X�}=�Z) b��m�b��y�T�h	p���q(^�����"j��,��bH�&Ȏێ
�dC���U*fYI��*�j�Q���H�SmPm�+�x��i��]��'���\�vv�m{:\.	1.��SR(^�_�Ve�LJ�ZՖAׄ_��� �#HY�,t��"R�$���Ы��߸�R��U1M:��<��Ύ5��n�	���¥,��8`g�]�<К�n�p����ϩ�l��ۓ���ъ����Ś(�+�K�k�٩JȺj4���E���p�O�[8��]�Ko�"贇�K!x�!�g��!I�Ve�w���NE	HbI�0�J���v�����gKNM>�;���Co�%�#��.
��;�p]ޫY�L%B[֨QX���ee��G�-8��`B�D�.߹����$!���u��9�q"�o�I�$*)�fj�U	iF�'�sd+�>��ju��Div�P���ܬ�w	�%�*��oǵf�e�h�ܶ�ܳ^����Grn�Ci9F�/�q�B�����']aK6mB��5��S���L��KYW���_qK�n�9�����0A��R�g|\�j9�Y
Żsc#3���ܙI�����F����@�����Q�!M�$(���B����zn���T��x�%�荹�sz�`pj��6�S�B�E��x��=1D&)(U9t�뾹��|��N;-`����}��y��7�!s�%�iMo]N�:�Oo9�?C��J�sT�*+Ė���DP�&.�+��,dn*4F�Ӯ5�r����/·�~�=֐E�I�`s���5Ɩ�>�DI#ښ�FW�XCZҭ��B�'�1<qG�h�Y�ފ���JH�q��J�e3U�گK�p��M��k,ae��p�b��GT:�QSE:��^"	>���z�6�-:(�j;�TE�*����q�����Vՙd�JJ���O�C�Q�������[�~1s�v���
��<�M�<�n&��٦DoR~��Y5K��±sEfx�
���y2���$�щOdQgm�|�x�G���E�MI%�-���9ӓ�ΑK��(-� ��u�?x�����'����)��߻�#M"�dVh��L("lr���%���ۉ9�p�����.8���*ZW֫�� �.(��-�)��!Q������J�GE'HR(�.R��t��M��q����J�ާv.J�
8g\�Y<���d����u~�9&�Iw#���%�!O����ƒǗ��}���Q��T]���O��b��C�m/��;C\fw�U��W��ӷ5�p��0�Eqy��{ˇ^�ѐCv�%)�D� ��.��\�ce� �Mպ��P��㠅{�]!�ɘTp���ܒ[dМ�!�Rꌍ!T�(���	X��ɵ�i��!�?@@U.�sW_����OH�d�<G;7���'F��b�TDs�w��M̐���beDI�}9���p��=���M*�C��K\�ݛ��Ȕ����ˍ���F��du�n$E��Q�N{�܇z��M�ߺ��:#�RP��E�9�p�|���*#I�u�|�l��l?r��Y��	�����[��u*:Q$G��c��&d��I��4>���k��}N�R�=���7�k�vc�#������������A�m�#��C�4��^�^���i�d)!W}x{sSW���T�5�g4�$-�".6��)Ni3!SNh����i�f4�Uʊƽ��.1��`��Ƣy��j0�S��}���p�D�B\��*�u�D�АEd_}��s�,蕠d1.��-ީ��uU-Ӛ.#^'�*�{�&*ݩ��W���a6{��g�2�*(X��a$A�bȽ���G8�R�owڮ�|<ڴo3���=��ܝ��%U�c����w�d�'�'̬��߄s4fA��	��#��{�{}�7��u�Y #e_DQmQ�)z�܋��=]�{�fm�<��5m�!���,��ϵ��ԞO��i�_t��6��o_�Z+��*�o��s�����g���f[�q�!�:֍����V���f�(������_u�����n��4.9�[8П<fU�໋�OW�G���":y�)w1<�OJ����5{��s����f'��D��� �j@i��R(h��X�M�xv)Rā�sי����Rm�ux���i.s�o��6�uY�F�[�*;��k^�m�7:�k�1�}k�riv�N]�Z�FXYe"rʶ��t26+)��sM�[�����p�0��=����{	�CwiVw�]�-#>�|�v�����.��Vl]6&��ffx1s�lD"#�m��R�va�Y�R.�,aIP���}{���I��ZU�}6����	_9�~���6c�U/��W�̜��1�k|�->�mimH��h�_s�N��$�2��?�~��N�Twj�4��ҋ,�Eb~��)֧��wjU�����DY�+����v~'h�hW�DH�����ih�H����놄	x��e��m+�W�"��{׭u�v�L���1�|�S�g�ga`������p^�_mF�w{��x�)�w�'Y<��|XG�Z37}Σ�^�8�8TG�Q7���;JE���m�c�����6ʮ���)ԝ��˟B4F����8�]�x�-��Ӆ�#d�VE	vދK���\.{yP��>v�-�S
���iWy*J#DZ�{����yՆ���%d-(WxJ�=���dy��Y��ɀ�Y�[�<�rݬ��R.�P��w�oMٚژ�jȱ{��;=��r�wŨ���"Tڂ�J��L,ƫվ�����E6�߄���׳KVi�YJ������z����#@ct&��\®��UۛX�`�MXl�ؑe��	��-^�`ÂZ��U�~�?[��H�_=��/&�EÜ��#u�H��ʯ�}��Ä">iL�����t�Z}F���m�ZgI[\�!Wf�*�^�kHE;�:��t~���
� p�$)�`aV��[��F�+��Y�C;*���!k=^�C�谤��2�jPWt#�"Ɗ�A�q���b;]�{,���z��wbE
˖B�Y�x�|���Z&jn`��W]QT}�J�m�F�"��_|�-B��	n��	s}^�̮C�q�۬{϶ú��`}��m�㖳Te�
�9=��/�ߝI��y���$�7��[�{_i�[�'�-=��3�VjU�{�ǩww��m����vo�Uq�M8�#i�{=�WLx(��U�n��u���\1�MB����#)U/�n��K�2�7_���ދD�����2ܥ���Z�^��M5^���ޫ��8�>�V&����w���'K�kJȆ*"E��'}��D�Tꉗ3EMU���͚Ÿ��oű	h����o��w��Es��%OiWZ�J��b�R,�K�*���׷Tڙ�SN��\���<�P��+hG{s=w����������0����h-��TvNKw%�[u�q].Fitq+��P����WJ��1H;�db!>A�#r�`��.u(�aX"/}���iI)&��o�OJ�#�x^��N�~�qغۡ|��jn~7W��f�{�T���U�/,�=�qs�5D��{���5Ļ�w@��=�ݧq�n�#��9I߽\S���{}J�q8�$��9�ӓ��z�������3������}���tڵ ���=��Y��u[:�G��Z|����(���̥%�����V&}=uɾ+�P��Wԥf؅ۥ��K�D8��#�a꾳+��EF�Xs7k���)��o:m6��$��g��ձ��My�"��Iʽ�ωݯX�j��!�����۶���+K�Q��Ⱥ�x#)5!�cp,��y���|��C���F-���c��j0LST�@�3�|{���諸iG�j:s���#)E�i�M���ճ�5`U�F�r�x;]:.�b ���^#�K��/x��IU�\!�����;�7����r�_}���K����+"��B�^�v�=�-��~�/¾��.0�B��F����SJQک�z��yM�H�#��t��v��	©� zjT����e�a�9n��=�����M�=!��2@wg�.��4b�Re�!׫ܨ�Դ�5
���{d�*=�ب����o��Wm56֖~��i����f{�TG;�!�2���ݟr����=��͇^yܔ�YH�Kn��B���ݛ�V�7�X���>T��?Y���9�8�g"�H��p�Mb��N̪O�-��#ۺ.�wE޴����9�9\�@{�W�ߖ����Q��N	��u�og��5�D�ݬ�O|�xɞ���W���p��v�{��B������V_�a�)2�;ܫ!T=���t���2��W�NI B3N$�ϟ��ZS�c�k��Qf���oĔC|��:�7N���~J:�|U�:@����ͺb��;h-�w�{��V]��y))��g����N�U��:����SϘ�'��C���oɗ�V��Ŀ����޽֝aD�y~��F��f������r�����}�6�|-6��!�{�[Xԡ��x�E�hWw1>=��)�ڋr��;y������W�X)-�����<�}�o���I�X2ͩ�v#�P�z��n%�/;�gh,�Y�B2��l��.B���C;Ҟ�G<5��ޯc�1~�4��z�%W�I q�(`�i.]ٳ<OUI�ʥ�KpQ��F�S7l�%t�$ ����!�	>�\�Y���4�7��Q捯����w�Q�\~��/�,|�v����y�ͦ�=t��3[C�G4CܤV%�EHJ��	�}<�*�j�������X�R�'�}U�{}�׶A����	���ǝ��*������Ш��7�["�	�p�S	ȗ�)ԅnƱz+��.UB�'�z��_��cݬ�֎��7�5�c{�Kp���Ӿ}Q�y��xl~¥���X��ո�(H�&�7d��A8�qoA]C5�}�Tq��f��ǖ�J�%��Y��:N7@ޕ|�+w�US+興Q�"ʈ�Q�#����Q�#�DDB��DD(�Q��DB���DD(�Q�DB���DD(�Q���!DG�Q
"DX��Q�#����
"<�"D(�j"!DB��Q�!DG�
"D~��!DG�
"D~��!DG�
"D~��!DF�DB���b��L��0����� � ���fO� �Uw�E���   (  (�T �PH*���� �  i@�@()@
U  �)_|  �        �      AT    R�   T    �h      0G��}��c��0vo`���tu'��y����UE� #��i�<vrѢVܺ�5{^O!�zt�0�� wov�.�/J�^wv���Hi��%j�;�tQ�6��OI�u� ==�q�n�A��ѡ����V�:�p7��i��@�=�{Ğ�c�=��j�y���a�wF�=����Z�X��     @   ��5��r�{�������os�o\����� :�/�-�4iŧ��F�齷��d;��j����{��=
�{�X�)q��6�m6vxΎ�
;��owKz� ��[�N��w�r��#��d�r��omٛw�PГ�ݯu�@���X��nZS���ܼ��l[[i-��-���     z   8=z<@�y�ZS�`�N/C�h�� {�ݣy�
�v�y�{9���F��K������ dK�݃{tu�Ω�S%f��aml[m\cA�-���TP� Z:ST�+h��7��5ŧZ�w��󫢭� `u�מ��ԫ���!=���={es�砬��$�SkIX��      �|�4\���c��ho;��-�Ѽc"�m�ۡ�cС$��� ���֔�Mv�C���m�3�v�ixã�$}�x�ݶ����� 8{�أl��uW��=��u�$���mm�f�M��=
z��J˸^0营�����i�(Z��u�9�:cyc�l�g]5����l����1�Ɗ'��G��4(P�}�=�F��;�u��r��|f��o_w��0�v�lho���$��Y�{�     (   /��j�}_w��Xm�˻i��k�gR�ٷ����JY�������t�:�u �jr=��M�s׶QK3���A�É������7cLz���Pٛj�l46 (�}ށ� 
 >�x =x4 !��w �讷�Ѽ`�T������.��P}o����OCC��ZN���h�������­��.^K����~%*�OP� S�LI*T4# 	�"��#)U&�d ��ʥA�*   �� ��  4	���A��M?���W�c��m}�U}_����E���yK�M
��s�5��l��� I!%]	˟�@	$$� �$��HID �BK�@	$$��B@�?^�~���~�����F�C�+ŕޜE�
=ۚl�nK9����ȟ	n0�B�M��֥x�p��f��n(�żX)77C9aaR��G\)��p,H�{S���7�o~yN�q9�{�4dI<��^���S[���i��8SU�6������z�Ӛ���7�����F\g�'n[���v��@z�@��D7���3.��3n�{bK���QH���P�3fD��MMԛ��^1M�ު�k����FN��ޗ��\��:������:�٭���pƹ��,H{�x�,�=�x�x�1��b�WX7���Q�z�����������s͝[��e=Z6�eP{p�܋X�����?���=����������
��ͩJ���j�X5Ǵ�]t��5�����F�];�Tr��OeL-�3�%\�޸]h�:ݕ�L_K�o���cK�}N�A�\%pPNr���'��|z�Hv��k�����:¶f���^��j���Z�7kXy�Y�;���>�A�>��x���@-�B G��e]�j+4�]:��k��Ѯ�]X�l�Evh���wuG�w>3y��f���bW9<j���i�Zh��Κ��>��a�t�G�z�s�{�g���[fKQԊg���^��R��,~s9҃<�c�_A��5�^��;9�n�s�/$�͵G_1Թ���2�6q&�sA�9��Bd�b�T�\�c���"�/��\�A#�$�ט�{YO�3�ĳ�Q5i�8�H䳛lLC9�c�;��G��z9C#7�8�9���d���)��,���2��-+e����z8"8Vf̱`Qy�8�T�J,j�4"�R�����#�7&��� �2"�u���J�0�,E^&&΋6$�,<u��xVk��Y���m;�M�nȱ����;:�f1ݼ��	E����QH'6�G���(�+igGt�X�r�2Ҭw�ٷ:Y�&<�؎A�����W�n�l����,C�+�����W�k˝�s�v�:`��42ic{�k�Rι�C�����|4 ��z�I{�9�5��N�=F���t[�.�c���p���Lӄlۀ�r��XK���E�'2��	=I����ܭ$s��2�
訳�e9�w��	�+��-A��m�9sgvwY�83�sx�W�-�M�(cA`��%��;m�X�<SU����3^��&���oz�s׳p��Q;�r=����pl�joJomZ���}�u��0UH@�4]%��9-Pm��˔���ә)ckG�҇�U�v[M�p�f0��&2��.�+w���]浩H�X��p���XD�;��	��4��m��\�I�:Gö��%��X;���Y��|eg{���u��>�M������-t�ʹ	��n��󣱌Tn�quۉt��l[�p4(^���s�2��=Ɇ.�Z5��rv��AС0�;�.Gz	Gs<�	y'��ӀӒ�X+���X� �`�l���t"���C�˃��C$�9�B7��h�a�Lgu�剳�T]-k��q�^�ȡ�&HK	���B�z�-�sI���rv��N+��\��R�#�3� �V������w�珁q�cx��NLޔ�+rm�0L�Ore��p�S�yh	�g l�7�=̫S+��q���H�U��L5%���@w�Hd�B��ё�$���T%=÷���P^���&Jɂ�/������7�!����\�-�5�8��!�o8��pE*Rʖn�EP�z�r-8{7�Kn'���C���p��KN�6�˰G���Ow�ł�V��Zt�
���6�.�o;vr�E �"ܫx�3����=�)I�k)��`v�����.�����v��Ru~�O���Ӭv���U�{�o\đ����3�3�lC��鹠�iu�N�n � 98Ö<�4<���ŧ�����X�ީ����������`j��v�rG�����d�b/O wqг�:k억�l�7GP���X��U�&�ٴ>�f�)K"�8��B�Y�Y�压z��rS�.�<�=U���y�A�b�V�k��o_'�	�v�u�ҩz^9v�ԋ��D�أ�Lz���K��]�f�/ѭ*샣��B�cñ�v~��+�����t��.�df���n�r�X����X0��Ef�0����j1��=ݪ�\9^��*�O��c���ظ�cd�ķ{��.#z� ��`��M���@���^�'��F��61�k1`y�U�E�@kKFg,�nGD)<���au��7����{Jq]��8�TF���GMX 뽚�u�&@7wF�S��뵃k���y�8!Cw���Я%�&	0g:2
���6:n�k��df�A�YhNzx�l�^=Igc��YLPW[�P�MLDxM#���Ɛ|1s���:�괡ѵd[�nl�r	 ����hN>Q��P�騜��EB�(�FF��lWc��rL�hЃ�/^ᅺ��+G��h��[܁(K��t����! b�����./�C�'�F+�f�ư��H���\m=f�L]9,�oQ�3wY�-E�{�)I� �9!�!�kYG�U���	�r���/r��	��{�%:fu�=���ٻ���T�`��^_��uD8��D�8=�[!��y^/7����6��b�������� ]��M~��λ��z.¯I.�XD�*W��`�]]ۚ�}�(�r�@G�[�ch 7`��`'��?Q���=��e�v��E�i�7�!mcc
�?.��!���#�!Ǥ�TJ2��V������)�{� ��*��s���p���(�3
-vG�Ԍ1�@[�(�Y��,���������f��_AQ����nnĊ8��Gį%Mg}��#N-�@��M=J�g*�s���6�S�Z��k�½T2�2=M&ǂ��4�Ԧ@��wM����r��0޼ԃ�M��}9�
3�L��0�5M۰� ��k=;R�s�F����:�"a*>ʷQk	a����Ć�(B����*�lAϻq`��3pC
cS:���p��˜1��V��x#ʭ��e���"�OG�u	�B�M�m�4=�A1+��ȷ�I�b쭻�v�6o��d�w{p�5�ÐXI2ep-�Bje7{����������6��J���Ѻ4%.m7�<���L����m}z\k��'�]{
0�[BۤJ��TO��5�bU�Ynd�`�tR\�k�ew.��8v�+����|9��}��8���w�VMݲm}Z�hHag�\1�'�h�	j!ӧc��9�u7gs+��WNŠ���Zjj�QѮ������y��Q���ܢhwVۃt\�sF��U������dLec����趮�Bd^syy[�u҂�9��`(�b��Z�YKښ�ƾx{����-�.ҡ�,;P=�����Ԙ�څ���bz��J�T��?��Mݫ����ķ��[���<+=r���M�C�{ӿx��Y}�I�.�ӑ��v��0����Wb[���k����K�nF�a-5BA,;Yrd��h�{5҂��XS9��)�a:b:�Ĕ-�7��d�����v\`��)�e=�P��B�cjR�͆*z性9�۶Է����wl�6�\�n�ܛ/f��ta�9Ӹ���;�i�+Y��#rbkV�hQ��?iT���8�4.��swk��x�v/ۺ�c�≹�DQ�v�V��ZY&�'�uz��dYx�y#mm�EH�Q63X�w.�{���{�=�sv!���M�w�$1%��=�����5ݳ7w�7�çle�1N0S����WA( q��^�.귦�ψ׵e�[r�+_�޲Ju\O��s�\��<J��0I�Ni�E֧op��͙Ƕ���zu�숞�{*=�"�$�\�$Š�$��,\:ފX6)3��h:�^I]�Uĭ�I�$�n�ILy�����.�yf9ׁC.�{e�3���g$^����q�;^�K`!����Ԡ�Y�C$wp��n-W�e"x�G��BDQ��̇ĳsJ͙^(�7;����'e맲KN����K@����j-[�-�L/�����;�,����Ʒ7dsK���������sD�F.��.�+�M��[l���O�ci���E�C����I᳕��� Hm%A٭n0�]�!*p��MPp<�ߵ��u��r��{�n5\9d�p�ۥ�񳳑�f�� |�s��o&ŀ�T��+�u��^�n�ݡ�Y�*�kIݛ���B��-;A��L�Nt}C�],�ă�u3�` �wiGsI�*�<�{���|���2	���AJ��1�7�6��iDM5�8im.OU9�7 #S��Z?t�q�/���y�^kGv9��u��K�Zx�o�$E::��F�}�С�XLM����@����a�  ��p��:oj���u�Xi�i`GB\5p����hb	���E���-��.�e��g0g�Df�*J3�&�V������?�X�e>���|�"R� ������<if
�;/r�CFsr�� �tl뿋J�;Bޚl�\a�͖#ϧ�_9��!W�k�Zt�w)6�s���ʋ�G�Ὤ��V:�4v7�ңF�]�Vh��d��w]��J���q��������lf콤�� ᣏ��8�m�R����h���N��܃y�M7�b�Rv��hs��]vGs_��M�^����ʜVj�7����z�0I���^åbа�Xy��Ӎ�ѷY2Y���k��t�m6^R�wv�F�)�@` �^�q㢭��G$j�j�.�od��(��A@	�}�~7�y���َAj᧌�P*�8�Gr:'m%��C9rܛ������]�y�3���N�N]n���:x��V�ŵ)��wXn�uZ���ua|��2��
i�{%���41�'N�;l�S���0�+��x�&�g��}���C5i�-�[�S���O�2�+�����c�94�ݱʕ֔�f!��{F%�N��ܺ�yZ�v
3�ߊ]�-Ko]QЌ=��V>�{�R�V���L��!񻭧����,�rQ�R�H:	#e��z�3z�{g�7��x�R��p��I�C�,�n���v�N�a��8T�Lc;q,�����wkn�����!"�j�5�8�-zc��s�����}�&�;T�=�ot�U]��N2��:�=�	�T��w��0��D�u��i]GO�s�l��P�P� �%���:�k�s���IV<Q_��k�j����f\wzL쯖,���n�ϧsK5hLo�d|;�w���Cݜ�&��)G�X�m-���f�y�v-���bn�	�#�U�I��	')�J79}���������i����.Nh��Z��/BfI�U17 
s�p�\ {�i�8�0�1	�i��fJy�K�6ĕD��y�����5b�l��Wk摁�v�N����+.]uc�$؇2QѺ�Wc#�u�y�v���iLܚ;]Ǘ+go��_���_M�]��n�u��l��㸲�s9��͛͝�w_o�Uv���P�Э���\���
aG���r���k�%��10����,[ҽ���Nn�s8�QKr�a ]Pm��L2ۭ��"�ǳ�L�v����Bdl�4��Q2 �	�NtB��aܘ�����aZ6��7�F����f���Wgc�%y]�r��%Ջtm��$�S���@vB���N_�d�N�n���W,��sU��6*�x*�	ڮ�V�a�ۥ9����D��fj1�ܱ�{P6E�P,�����z���x�I���9R����%6u�5���ێj�!.�!q�q�����L������=X�C������;�:�ZW���nt{/Zm�G)w6����H�}f�͆����k�h���?k�LpA6=T���e�ҽ�2gvl�U�LU��Z3��r��I���%����n͏b۶ŧ[�<��-E:��G��"]��+��H��@SI�x�1��N�*q��1;����fa"H��{����U	�Dj��e�^u�Yz!�V�E�s#�{�I5�qJ�G�s.&�]�3����&	�F�y�4vP��Z��Ks��֬�ڝ<�O9�@�mj׌��xt/� �x�x��=�p��E�UOǟJ(�v�Zu���X��g-�U�{&�5`��xTp]��$'l<�B��=�u�NT$cX��NU��ن��	B�dE��vQ�D1��85-��e���,Y��W�{��g�����&�r��D�z��+��	,������Ž/e�t�A����������&}z�.�/��g���,)V>���U�f��ۢ� �<󨘧���`~D�b"�oP�L���i��@u��z(��-�]� !1:�vk�vƮ�|9W�r�Z��E
%(���u��p�+��f��2J�GtSS������X\i!BhI�r][V��u��s\ɽ8�Z��K�\�I�9���LntoG.7���d�ޒ��[���	(�.����LѼ7{7��N��BХ��Z�ܽ�Fo$4���H݊��.�Z�XS���Cӹ(xd�G&++��G_X�4� K�>��j�B�6�c�&��V��������o4k�����8�{�����ɠ���.��߰Pԍ��ʜ�2���*��m���ӫ�L�%[��m���;�m��V�gf��"�uJ�J����)�
�����F��quة݉�V�����T�C�vͼ�S���-X��۲L�C�
]�.x��ƋV�g$vT���<:��H4��r�W�n���Dnrz�۶�n�ESu&ݶZ�8;Y����֚��$k������x��V��ζ��ٹD�f7n��������羚u�usqk�p���/��Ƌ\FɎ�#�C���wn�O��\I�G:c�t7���p�s������YܧR�3��O]qvtm��t�+��V}7U�/n�x�]�mf����n�v������r��g�m۱f8��6�ك�=lm�Ѹ�q;�q��L��Oh����� j��U֝o2%�i���ZԬ��Q����� ,�bl��'W.^�kY)���n���d��c;�^�v�������K���U�:��}�q��v7`R^J��5uՍv�w�p!�탳t��vƅt=�ƻ&�M��(v}4�¹�t����qݛWe\ݢ�jy!�KXfMv�ɘ�<��Z:���C�gJ�!���g�g�7#r�횷E�Ѱn��v����4Ϯ��weG���U۷�-�Nܨ=N��tN�
o��Ō;�yM�D�a��@��]�nSu獶�X^��0q%k�/H2��.<�떜�%�,�5�n���ݚ2.���q���H]����n�"N�z�i�[�=cq^�s��-s���>;tr�շ�s�V�W��r�u�~{��[@%l�5%��}����.��v�Fl6��Ncs������C��n�/��N,�=�=�L�>4݃�M�ݶ7&��'�c7�M�p���r(nI�<�K�M���1���=mq�ݔ�WAk;]sȷg������{X�g\�a�ؗ��/X�y�9뉺�N⩸*e۶�y���W��^�۰��y^�rC�؜�C�tq�e�v��4kkv��Z���&�	�q L��n6�ۡ�;[��՜(V�=�R���=����j�u�W@�9�;��`��L�ps����#���"GWJ���ͧqPb��`^�Wb�x���c<��78�#=��u��<��\��ݜ��-�ې�71s!��U�\tv�wk�f7T=��l �ۍ��vԘ��'�gŁ��t����c�n��V4v8�u�[S�@s;>)Z��n����Nȋ��� I��9����^-.�[�MC���n��;����0�������	�<q�m�]�v���mn�J��Y�p��#������[�ݳ��2�����Nu�����`cn�b7:㫦�2;b-fu�c��u�;&��c�3����sJ��<hs<�;3�m�Z쥄�[1X�%/�5cZ��p�=��O�9�u�"y��F΍������wt�텯@���sq�����q�Yq�k]����[�j�q��7<�7 ��.�m��:��ɛk\b��=��Nw!sm<����[s�ׁ�]�ʇQwe5���D�:\���ø�Dz�F'�pg����3\��$m;]2�m�K�I��v�+Z5���^3��L99�\���u�].���MUbc�.�q(p���lU��c�s�{l�m']�\�ۋ��6�s�g#m\1����k�^�C���!bĐM�k��$OCE�����SS�9�v�%�{�N�g������;��[re��=sa���r�۠���v��T���x�6b;��w��𛮟3l,o#�vxM�<<kN}fyf!K��ɳ�wn{`��Wo4�Ɖ�U�9��ϥ�.:��1ڗi�:��AF�z�w=�t\�&�m�v�-��X{��rs�r�{[��gc�h<(s�c��n�Ӱ'n��m��wbݸ��:.[q�9�+	��w-j캗vm�g�l)�U]�[ru��=��q&�y�w�)�Ǭ���݁��ðZYG]��sN�-��Ӄnv���Z#s�b�$��I�ѹ���<�%�� C����$�����kM8���x�s�ZN]��OgOb�P�f�oc�N��pQ�:^���ٟ��&�ۧ��H/f�x���V[��\l!�����G[s۞U������p��nD#���J�q%�&mY�S��;F�ڦ΋�X�=�탮3s��ru�W\˞�ݭ�tӊ}���q���wX�Ӟx�oc�V7[�oB�X�'���6���J��!\������w��=<l-J�n���k�=�����5'G:ʃ[�L�{^I��v�]�g���m6����M�m��M�_�����#������v[n"1�.�*e�u�;�燵�"�6{]v�gGmϻ8�mH��3�fc�5Ƨom��lNݮ|��qc��r<�+n�g��vƽ[��0�k<t�G6�3�^l+Y��6�9䶬�nn��M��8�˟h�n��z�����w��m�;=�q۩�����jN�7n��6�d8-�n�z�j���3�J׆��m����Gq��G �I�;F��d��{�Z�nu#���}Jq�Y���MA�As�ﯸ��m��[�@�[��|�Ũ�v�Ob�н�|V���lo��oq[����� ����ێ; bd�3vf2�v�v��g��ʶ�=h��n3p�9նf���>���&c�oE�����ׂMʾwB<dzۣ�ۋiCu���v.�+�Uέ˓v������m��H�붱�������Z�ؘ��A�����duc�v����-����k�B�^�zò���꬙���ljW��nJ�m�]��������p�q�W9�:��u<�km���\�.���j��d� �	ƳL���
��_Yz���˳˓4�T�N�K�f+R�EPZV�v۱�-s�Qw�/�m�۴s%ĐlpD�+u]>��gj��9���*;f�7cn��m��]���:����B�=��,s��;ۓ�j�K�>�{�2�z�l�x�n���^���/�f���<9n�6�v.n��A�N60�(�x=�<�M��n0�y��ןV��3��m�)���� 7�V+c^��zx�vu�"�������#���t��n��Ƃ$Nc[��4o[���\��.���m̓7ݎ��ū�tlny��´�e��a+Ƣ����n�tkձ��Q
�/\���Ԗ�7Ff���Q��#�xtMokF�G[�"���I�<\Y����ֳ�����V;{��wv���-m���{>��O,,�Ǥ�s�uj��<�kqc�7Um��ɀ#J�qu�57;G y�U��\2��'��=1y�F5��s�Lm�.��Ì1n�w[Q�]�t#P��i���iv�7@Om�l�U�jϐ�M�����ٻ ���xۑ�E�a;�c��͌��Jc��6R=qq�C�GGiPű��#eю�`�V���//&�)v=\u�b2KN�gW�NR'��)��u��ɀnw&L�y��<�z�mŸ�Xn��7k\k=xӆ��n�S�
�Ϝ�]�m�b���}wn6�l�J��NQ[���m׷�iؤ�}�8�N�3�ޛd�#������B�C�X
�B)�Z��rcV���lt���j�[��6'ƺ��u��RA�ؕun�'�̅@O볒x����m�e���qv��;�W8�Ѱ�x���p��u�..���M�ۦ�:�;��%vȪ0�t��+g���=�lg��V����y�"�"zlG�Gg�ϓ5*&��^Tp�B��X:w��]�Nؒ��x��a����ڻn�[u���
m�]��ceW�&=�I�s������l枅�/lAt��W@;Xq��7ێA��Nz�su�{\�r��Pe��)����5�v"�@d67�Uǫ�u�xv6�u,��E)u���.5���qՇ<nwv�2�af��\��/�ly�y��!�흉{����o%����g�x��ݼ]pnx7'�8��n$�OP;��s��GX��c�����Ӣ�tKɝ�ӱ�ݮ�[byⷧ\��@g�G'S�K�;9$^��8W;M�t����}��Ѹ�ó��z�m7������<t������해o9�]�
@-��9�h��M����cR09m�����ۖ,�����`�ύۙ�_mg��m�h��x��	�t67-��u�8͇�b�k��s�!�l��s��9m>��6�;E���3a���..�8��ݷ���-��Ş���vC�vΈ:�݆���h;=��PC�ig^U���� ����N� (���G%�� ;z��B;�ͱ����
Ș�Pb�:( �|�ې�����"
;vg;�S[�g����c��e���N�k��\��=E�P��qg��	Z\�hz*Cq�]P������+�rE'���5�L��'#���]��5�nc�ֆ�����7<&����֖�wg���y��만i�m�έ0�oCG��nV���n�m�yθ�Ma�ƻ;scg�s��ֶݎG�ě�|#/}J�WӴ��pn�m�ı�y6W�p��9�	K���֭Lu�ns�t���6�Y�;ګ���mщ:���3�;��A� ���c�1؍�����}�d)q���1��S��i���ϷK��p�8�/݅�O���z�yC�'kz3��l�M��p�]ۇ��C��#�:"�m����Ƙ���]>�'�nu+�����j�۝o=�v)zn���d�Ŕ�fŰ'����#�+��^�}�ڽ��8�:��ȇ�v�
�T��m���crt9�ki��K����.���4����t�cۓl���W���O,p�YQؓ��;V����>����ݤ7�s�l��g��c����-=���u���/j�x[O���V3��O/e�s������X����B󻞹��d�����QH�̱V�8d���R;�m�����*�8Gl�-�v�mF����緍e�#��om����]�k8��?����'����z�gu����zT]��ŗ���Ϝ�`�=��6���>�7uګl�n�k;�f��FD�g��$	#��b^i	/�HI1
D�F��b%�T�̵N�ӊ�n�n�0Zz��nx�s[���݊����z��iA�
��3l�^;:7%E�౎ٚ@F��AZ�5dV&��O`A렩��q�+B��_F���s�v���n��2�N=l���'`[����un��#R�n)z�@��Cv+���7!����:�5���8�\�v#ai�aw`��N��Y{{gt˄Yp�+J]qs���K��+�^�{��.e�p&b���Ch��N�x��u�a�ڡ��g�92''oGk���+�+� K�ʔvͤ.{�K�Bٌ7�H�ٛ�]����<t�vg%��%�AM� ��x�uZ��:=�v���vk�N��O�os^�[�{�#N�=�ˠ�[^s��\�ӆv.�l'nsv���r`�v.�jWqk����YS��\�T�k[�<�n�W�v��6|8������xC�s=�G��Lr8�oh�M[��Þl;���^�y5.��2�&������݀�4qc[�t�!��Z�V�'��+�]�w��aޱ{<�M�9kq�u����˫'[��c���<�h,plg��1�,��wa7kwix�Oaz�e��91;WM,��&ٮ���`滷���M�P���y�x x��c�q��oO8���I�vB�K�q��р�qĪ�wt]l��/n�&�}�[{n�h�Cm�в�7>���i9��;;:;�	��3u8���@y�9V�0��k�=��@�s����M۶�n8ڌ���x��hrWnv9zlpc]�݉ELpoYv�^��c=���tr�Gdy}�g���kv�q�����/�zaF���p��Y�յ��1���$�-�;����i�lv;&@:�M:�^ݗ����TmRe�M�v�ǭk�j{��c�E��Yϫ\��S���Z^��0�[m���F�<Q��Gwτ��w��$\K���Z�;�5�7c���{l��كv:On݌���+eA7�������*s9�����ň$٤��@� ��	i!`� m	  $ &� 	� 
D,���/ӂ�ўe��n�܀gr��x�꺺+u�L'���[I�۞g�����M3����[�&�n&l{p����'G3�-�;�'Q�m���X�`�6{>��/giбvR�Ek�^���6#Q�gg����k=�/v}`����D��x���xci�5n������]�Q�M
�J)BA
�QA�t[$�[5Z}��z�w獱��C��rs�����;9G�]��gp�ɔ����Q�?�Կ�������j��Jf�vh�o�.ڹ^C�B��f�]飭��I���r��Ъ�%�-�&���ƕ:W��C������P���i)wd��s"��
g�nS�2�Cƙ�j��D���d�|�by���7��.�B��3Szz�ncHh�!J첪�W��u�N�=m��.�$PV]�AQM��F�-�#)�����+�J\�t����C.�Y���,.n\u4bu2�+o�ʪ�bd%w�X/�nBd��V V���B){vO�y}%�7�=�%=Pں�6���c-h���J��D.�=��4��6ڃn�#(�=c�tu��p5��M�v=z�Gn��ݗsX����)[�𻌬�7�3����_�Z�c!~Ti�����2y�۔R�7��i�2o�A"؇L�M0�t�:N�jG
@�1�vltsK���w)�\/������k�ui�`��z�z_�y�ê*��#�B�=�jX}�q�5���̙��_Y�ǎ3���x�D�!�<ǥ���󞔋7�c�����vm�F�+cp)�.��OEۨ@ Ec�e�.��N
aIzx��㔽z(�԰C�|�|$��/u�Pe��l}�(`���DD���g��D��/��/�����I.�J��'w�/N�ukl���z/�ow��g
k����uH�&�XBѾ���b�~�Rl���X2�b3D�R;@�d7������1uB��ݤ�i1ݐw;��7Q���Z�Ҫ}�w	^�"O9��;ò��q
%4�0�Lޠn����gp�<������aǨ ^0�� "��2*��8��c&�{\ߺ�=x:Q�yQ1a%b����n��;l��<��_s�-Q]�c#�ֿ�1]{bw��<��7o��"4~6���E��� d�N^s�5Y�s{��+����ėDEO���M���S���ch�$�6IJIH6e ���o�5{"1Ӓ���<��;���g��=�ʝ�_۳��2oJ(�s����v��4�2Z���b���R��]&9
�(�����8�~���0�&��k����1��ݮ����|ڪ[ *�%��sej���:MU���t�z�#��س�*�ث#��a���P���}�tӰn^�$
%-k��U݅�r	e8@�T����+�[R�]�����
�V���d�yh�Eͷ��"��6������(�9����M����������6�\Awey�=MR
`��n���m��OS�qn�'c�����t9�Ҿ����!�9�GW��8d�FD:��?gv����������r�6�nӉ4*)�)�#bCk���U�R%Q�L�#U-]T��_������5�}�Uz`޷W��������hY�~:�ߌ����o��Ȁ�����r;����~�C��3Dq?��E���ِ��[xK���z�n�(O���~��^?è�NK%%�r�܎���~9=WT�#�ϭ��L�BT9 4mz b��Vh)��])��#	�z�~s��h��O{v���8,�L!pl�ek�{�w>�o:-&q4>H��'Q:Cjv�Nn��x�����v��s�� �]�AI��fs̺�zxg?\4���U��A�}e�w#�#M��F�u�=Ǳ���9;�m��ٯ�m��a�mn6>�R�[��<����7w��������u�Ǘ�ephjD�-Q�CCD�aIDEJ�n�9�mk&�8�˥�A��6죶�������.�]$Jػ�n��"ȆM����#����]g��s0ԗ�.�V���yzw��2������������D-�AZ󜔎G����f�)��*<�Ϲ-������c�.!���6��m+��-\է�2~�?�$�~��yt���ͅ�p��6u��Ig�.�<���}�o�xuD:����9���bmȪ��:�(����.��r
����m�U��0�E�w}T}U����.��>�4.����:��)/�;x��U�v�G���I�]��2;�L��Т�>wʍ�d�B�%��
1N)w��{��)"���j�������A�ߺ�S��&V��==U����_�Z��b��G�{�i�*k����������M��-�<�0e�����9��3��"q���{��=��6g;�=�}�:�`u_�:�t�NN��.�vfK7�1O��E�cY�x��wu�-�q�GlQqp��~~�1ź�yy��6��l6xr��8f0���pێ{�H^�Ն�9Gǂ�X]�{U.�uɶ�FQ���/&�v��%��H�2m�^]�vr�{��'3�Vx|2�kێ�b�7]�a�s��=�Z�ѝ3�������aKEیn�\ [>vλqr�ؖy�6�۴j����ˊy��r�6��Lܝ)�S��[&W�Kt��|��ۚ�]�b�9��Ȩr0���I	��zP*��Gv� I��o28�Od�N��fB�7�27��b�Ci9nȢ1F�Y�<R;A5-��n� +@�L�"��S�0tף���^�����8��(����BG-/ۻ�3��`�u��DY�=1�$���M�A�#R8	i��g��j�]Z�|�B��]ə>�&��3]��ڦ8>����#G�V�n�ֱ�\���g^��&�2���O�2��C3�3��'����F�1Ή�����E��^2�j��}(l�S翃#GAl�S��vz��z��"�<4`�
��)�~��҆g����2{\� �qy�Я �ͧ�:���_U8~mC�^E�C�SKkX������H�Ӗo_i���`�\���̄�J
�m���o:ޙ��	�]c����sY�?�����R$����[+6o�=�j;3�앦y�Wj�y!�W;�[��[b b�_X���}$c�D�)���1�����e���û������=~�2��n����{����ޒ&���ٱ�����%ӫ���7��'4oh!@�fF˓+C�N�6�'�Ύ�H�Z�,Z�i�"0�Ӕ:Iu}�켭N��D�/�C�{˦�~�V�x7�υ�h����H�1�����J��������?o�l�Bp������1e�L�T�h@�?i�;���r�;�c[�p@C�D�-�h��P�^����֕����W(Y}����H�!6W�*���L~y?a�����5��� �e�^�u�K�7@ǜ,�y����.Icߚ�@���Ɔ�H�Y��XLs��<���{��u�`�s3����^0(���)��nN�PUvn�|Y��
4J)	&C��Bc]��|ݷ\����N��km�;�R�%LH�q@�����T��C"�V��?�>�M�=�ݯ�)ztf;��25���E���^�f,��J<�@�OS�ϣ!7�Q�-y��Q�ꆧS{$ Q�*Ɩɪ�e*����&f}k�W�/��(�ZB�Ə���}��z�^Uw26��ā(���~�L�[d?���ΓA��Ԛ����`O7�L8�׫¹���4��ֺO�����z��۔�:ӡ�{�<˘x)��{Ӕ��ί`T���X,�@���R�|=��Q�8��lYex�Mo��� Xb|�h�&"�?7K�Zx"R��H�Kʬ^�?.u��c�^�o�t�e�R�������q�`�(���-�U�a�'�H��[�
^,=D�}�c�qB7mü���[�EVd{�D#�:PRp٬���uyJ��"�[��h��86��K8s�<��&BTm�J1A�u���v�me��P<��܎���B��u0�*F�1��Zk��!;�u���,���;��%�yNȷ�����tք7=*��]=�Cofg�s6D!�DoО;�OI�y��7�����<���c�b�����v�%d�ոA�WN�Uh2�?gN��5hWe�-�����`D,�ǅW�rH����m�o��`�:�%�� �:3�}�t���v���'�{�\�J�3�
M�ι�h�����JF��@�>�4��RH\m�QŸ�����9W�]�g�ӯ��!
ݜ�Di|���/��ޒ�G5lvwyo�r�$1�Y�q�4�w{RDc�e��%�v/yo{��e&<Eh�uƅ��lD�R���Ǆ2p�)م�8ak��j��^�>]8��7�]�u��f�j�L��t���(I�!�ǆ��fR��2P�l$Q)�6�s銢z��6��^՘�C��F�,+���+�{C�x��=��m�^�973��+=6�2C�Q���;k��dl��[���˻��e�vt�<C#�6���;a������0��p��E��F<y.�wot���h61��m5i)%!~Dpk��^h<r+F��K�eH���o��U��>�-W��D>����|������ug�v��
1�>I`nB����8��[������uގ��fƻ����Z~�5�IfΡj��^��~����8��&�REVB!O;!�Yw���}G�z2,��g�"j�ge�
qV/�$y5O�{�=6Fȍ�Ze�?	�|X=m��b��mO��su�����BI,�j!{��E��C���oN��V+g�c���K�#� 㼠;޼7��*�Wz0r׆Ӈdz����p����WA��W=��������u�����6�_%������Ĳ2�����3r�I3�e,qe�x��4a7���g����`0nKlT�p��9���q�������v7f�:׈��#.�Xn���T��sl�T�p��F��lՓ�.B������uO
/�蜱��8�^�k�����v�f�����va:�`���Y�X���鱲��ck��g��D �Bm��۝h��c�"6B���]غ��F�y�{uͭn������d��VRm�,=���χA�:���+���V�W�+p��K�S��W'Xv�N��-�č�<�[��!�v�t��K�S���web��W�gx�H/�G��5�gD��;���d�e�ú[`�w�7�AV�+�Z�{��Q:�����e�ulVҋ����6���%���}�Q��U����ŧ���J|7=�*�k���$b9#��i$"���H2��Y$֪/���r�,cj.˾;7%����\WZ^!-C�M�udQ�*�b�'�F&�l&d��o�����ʺ^�5Z_Ѡ�w���
"�E�G]�N�����o	�#f(o����-_VMwB�m	5���|�G@�J!N0�N����=�|�*c�q��~�/���h�n��~u�qxmۑF���W�F5�C�Es	���}[4���H=�6�l�����:���ɺ띹�)�U�q��u�u��kH��Kہ-ǯ�cy�3D�h�/��q�G-B!]d�aN��Uf^+��`-��m�Pg=hQQ�"�cxx0��\i��mHk��3>�=+�9t��Ы�:�D����hD=�唵�ۍ����e���;�E���z8�WQ�x]����=dǠ���;{��B��:��L3��e�����ј���� ����_�B���a�L��R7����y>N�eն���\uCS��[��qϴ�_2Y�Ǔ�y	٭wN�c1#��ΰ��	����^v������?n-�GG�%Cc
����m���Уk�V.��o͆Dw�{�ǽ��V���$iWdth�`���r�d_H.�l���|'$���Sr2�-��Q�ϢF⧉��o��aå�#�}�J�b�b�:�afLG�!R���AY�/08!��n��J|�^�ש��"ٞl�&���@���V�b�ΰ,Cڧ�k�ǃ�s��8�e���-�	�FW!+Q�)���Gj���B�4��3��+��A�hݨDa��v��j���-ںB	�Ɛ���k��t�پ��P��vY��a/�Y9y�hxj��^
̓i��= ����Ȉ�ݪ⠦{� �|�!��Ш'_D~�����u�KZ�ž���n����1D$�d�(�M�M5�N�|Z����`����rZ�;���2���=�nH��ۀ�px9��g�uqbY|��Wb��ʝ�) �x8�zż^Mu��͛UORṯ�@�;)]&��]Ѓb*u��t�u;��n�3�\���1��K�!�Y:ʞ�C�;N����ޔ�
�Li���0q�$�Ə,4`x{�[������1��D����k{��5�P������m`������;W��	�cD��ޮ3>�̸�@���f��᮱�xd8�/	u�ͲΟL�|es�{����u�z\��zr�p୦.�)z��Ozp��79��@�8�~[*}1	���Ok� 5P�{�z3��bB��x�嫌��FU}�o��9�U�j�$\��Ro}å�&�����ח��J9�t��Htn��n�ԳaHS�1Λ�&<��@�[4�A��IQ���󻼍�'L���7ƹP�$�Ud�L��ܜ��6��چjI�9[6/J��k�:�{�M�Ї��7W�H���C�p��ҟcVq$�<w\;����h��+��`T�N���gV7V�V����r�h�\*0�n����P�4W=��Wc��u�gl���Di��]�0�������;���x�4���Ӻ�]��y�D���5丽9����cȌ�5���}Ay�ܼ�.FMgᦦ�cnv'����Gg��]瑌j:��4٨��vA7�d�r����Mۆ[�A�R��d8�M����Y[P=�Nq����L��F�6��;������gA:�f��0��ݧSXh�N����B~���w� Yܬ��{����r(@�S�:i&�I��E�8o�~i#J���r�iO�Z+T�Ah�"�4~dq����m����sy�R�?����;�t�oj����\R/a�{^D65vڜt����Q��x�}B4�@�9(5�5�m�Wκk���ޒ�ZS)����,�Zn�ۓ�����&[�g�%*5h��?|4������D�ۍG/#���q��uv�a{.+�θ�ڹ^ޮ1r:�.���9H�L����]�׽�lH׽�l��G�yz��0.葻��/��͹^D�C:����ym�e�1r
�H�lD n���/�}u�hq���֚��(�yL�����;���8�a��#{�pL��U�[�V���dD�u$vV�К12;�s�|/t=E��O;j��dޫ�,�����G�������+z������T�q!g�3a���c��7Ϳ9vi�r��j�M�]Na�?A}�N�7��Ӟ��@���p8`�2����Oi_j��cx�l���|f�Dk���K� �_�I��ddᠧ$-�z�@c�`9Q��]�^Fh:����x'Q{Q� ��VhA �s�܊����9um%��4�^�z�}z�?TB������l���A6'"����zr��46�hy�hi#�43v�k�Z���U�i��	he�չ�t���X�F=n�0<wʙn�?�$�X��V�ȥK�<E��N����߄w'������]-޾9o[
h�TLo�_Wj̙N�@a
����(D�ݔ���v~�Z��2�|
�8J2P�FE�)�"�Gs�4*銼�YB�M�Ǵ����~K��p��PUc��^�Cue%3�_K�����6�����`5���R����p��NC�hE�?	E�Ŏ��d�Ϣ���|E�;��C���?���z�{������V��>����m���[ \i���=����j_��������X���OB�H1{Ӄ� �7x��l�����ah=#x�VC~ձ
� Q�Z�-�(�����'�/p�����Rr�
��h>�R�U�~ܻ�����n�g��{��W�e��W�
�r!�i�eV�~�q�����P|&�,����|:����i~��o���+ꀉ��>�|�0:�p������Ϟ���:��q�Tv��j�ځ����]Wm�mA�q��W��%dܮ�����sU��Uڷ`����QV-��G���L����,�|�bW�j�F.I�6mpsN�xw��<&x��98s�6�n8����[3�Ӎs��v/m��.#�3u��1��g�u[��ѻe�\]C�\�z��Al�f�k�v�\�k<Cy�>mFlu�V���f��R��b�#����]�ܸ������<�s�s ��v�j;iI	���?E<ޱY���"�u��6�	��R����%M�	_U�����\��:��i��C��!z8��%�N$�60�B��.�Y�-�6���o���� �5ڲ���{v��Fp:ux>?X����~z�>�Gբ�1 K��Rp���9p�f0Br(\����Ⱦ���8<GVT>����)�R�Q�1�F�lV�hg!]y��ZTBiގ(��bs���9>�(�.4 &H���F�t�ȝ���Fz�m/�����~4�ɔ�k�Fg�z��,���h,���r�g��N�J��2E<F�@}�l��'e�D����E�Oݳ\��N��	�WSs:�Q*�M�_dVcȅ6�z����Z�5,V�dO#��YF�������N���<u���L�Lvx��wlGY���w�,�Zy���C�d�����Z��d^Yj�8~�i���ޱq�
�������yh���Z�l�WU�;��^�0�|es1��y�-Z��������?ѓ*��3���c��Dݪy�6#���{�>�Z��l��.��Do�{��^Ȉ�p2��B�|dN�(Q莌{�_qvͳ��;�!�(p�)!>�z��~��`��V]��i
?m/�{:��2�7�A@{i�W!����s��1��ANJfl�Md
��V:q�u�pcP�nZ&n�����cۄu�N*tE!���۴Բ2s�����g;����g�1Pn0CLB�q1dU�!�`�:�s�?]�o�z��ȗ���<"��&4~f��<��o���j\�.v�ZïoZVn��G�)}7}(�w��`�߾D$I�hY��3��L^k�Qu���B�w��KUgP�s�^�c�~�P�h����eI�J�Wav�QZ����uNe�E�Z��BE
��1i�;f{m�`ט����Z��A��p�-p=j�(Ge���V �����n4L���twi"�cy]W:6�]�*����]2������
�I�<���f�%�Z���A�����*0Di)�xB!@G�2��4R�U��ٳ$z�?��.�YZd|�z�$�6x��#��k֩[vu����U�굳� i���$`��,Bc���uR|HG�Ԩ{$)�1�vw���Ĉ��U��杧�v�^S��;r��4����|-�ͮ�˼�h��<�o!q2�Jwg'r�p�
�luJ���X��e칸���r�	UeW��Κ�/y�����:F寜�58,�V�s�)YK�T�Z8'c)C�+?-����;Z(��ʤX�P�l-��fh�H\���7��g���JBD�`�cn*���?#o_��b�ag��~���Գ�{Ӵ5�e^����1�,����n�4��u�*[1w98R�R�pR�C�DƭUg�ckq����q�q��\�d����t� f�^ϸ��ؾ�W⾢M��,���*��E��6"�a����R��*L�B�B�|��݄m�=O��>E�����DJp:"��.A��w��|���c��,�2�1��
(������}�x7�"?Td��\Ǆ%՚*c:*M�OιU�}`�CȲB�Y�Ʒ�4��
<g`v��~U/��{ ����ci^���q�i�U �Q"�g C�!�2����^?31
���~L��	 ��8�)Pd;��d]C�'����;��U�=ݸ��h��H��"�U��Ўخ�"�Σ>e�oWv�v+S���y#�rU����Ś-�F�0\NU�j�������ATV�+�%��#���5p�c/Ǖ��%�t�;qU<�C޴�6g�@}���"م�N5�\�8@e�Τ��W�Q$6/�ͻl��lھ�zl[�rz�՗s��~��a�e�W����žp�+۾?qS���z��HԷۡ�n3D����-ūL�_��)"0��F]((�]7��M�ti�R���]��x���6}�e���6Èq�j���{[�����x�#�l���jÆ��Z���V�P�DG@x-x�B�.8�f&~�!�nݵ�,�`6j��!�;+�S���~���(�5�La$&�zc�^\%�#�M=��י�]��jo��
���Z����M�y���
ښMc�;0_�aS��:�r������/��ʓfI'tn���F�Ҿ��ױRK-��F6���cUkg۲��9��nZe=�`
y�~���W���h:H�*r꩙����ȈGN������
�)/:(G �K)%1��B�O���-�u�5����n�q�B��?$�Z�����dޕ�a��߽��<�>0b�!!�b���>>��ţ_t�*�񙻽�t�P�if�#Y;�ď�GC]M�^'.^��"��g�
LW|��g�9������2"n�K?H�d�U�g���ڝ�G3�&�t�uݖ2�y��Y��y�uD�9��%^��-ΈN�sY�H4v:3�ng`�ݸ�l��s<eP�qQ�'oh�,�dN	v۶�:cv��0����䛱�²
�����N@�A�(WZY	�%�<fu�"�O�c9Η5���=�5oXKş�ݢ�lc�m�݉C�� ��b�h��nܦ������h4�Ds���&@,��.\m=4R͗f��]�Dn22��"#L���~rrF��_�O��ƾ�A���,��ΙM������������{30���M|���<�L�X���l�$|�51<��/=��3��5��LIÍ�d-;�]rU����T�PZ��#'#n��w��:���$삈�ތ͎)I���W�����]ʦ')^+��Wb��D����Z�����CG��S��/eev!�>W�n9��(�
�Tc|al6�,@ ���kK3D�w���[����n_�>��X�OU��� �k�V+F0!Yp�Uؒ�
.f$��0�ݰQD��\a��@����6�=��Q���a^Q6�"�D�ҏK��lťc�O F8�	��n+5>g睵�Jw�L�lgu���'j����ꮸ�B�,V�Z�fO�W]L�k#�3b��u������\k����G/�h֍W�Q�
�!�+�k!?�8�Y�|�A풆�<�~�=���8~T����B���|a�ﱔx4<څ�&91#o��ת���{b&�`������z���(�Zf��ĨC��ў�'�K�dX˖3T�{�Y/��-����몰����;5�Ր�l�G�����D���w�Vy9�e�_���!Y(d^�f�^s&�=q����l묣��YSC,�Yj}G�_N�X���<{�1D"FR¦.���Ȇ��>�4y�)C���s[z�57&�\Fہ�d����ܙk�a�����+M{vw��"~k���a���O�Y�2V���������\/���幷v�Q�.��ȇ���ۍ�>F��6�:E��͗U}��ڰ��80E��HWk��s��C�Y�}��U��q
�GN
ݿ���dӃ�g�r��]��4�Q�iϣ�z����85aH�t���;���,m了��9��V���ui��q�Go�"�I��:�zrWoN#+*Bu{��T,�fGgz�-��roq�jB�'7[%%^:�<�֬`��S�˻�@�A��>�ۄ��=b2z��m��8��qw���
,�W+��F:D0���� p�@��y�~t�>"�s)�g];)vS��L���B��5�� ��u�3��r_���q]�����������;�����Z[Poc�	[;�@�j��\�t���Y�Q�bhr������������`�u����8S�������2P�4q���̿y�o�[k�ټ'��3��N���U�3���?e{V
#̶�*��^Y���Nk[�1��K�Pڛ�w��G=Ikm�Kj�ڼ�d���.��G�@@ĳ�6�{㽁������ (�����Co��.X~�#��l�=(n�}�ݘ\P�����1t�9�3���s�Ӟ���v9u���{T@E���*�?{�,ɖ*����!$7�k�Ȳ�E4o_s4��:R�.�����ec����Ő��细��d:B�YhTYS�u�z��߻���X�|2��o���:1��*�=4B�޲��:Ȝ�y@��w^X����㯹�d��a;M \n�Q:�(�rX-�5��ث����c�����n�$��A̓+qR_-�����ok�J�ʵf����ξdq8m�>qI����³A���J�}�{gUpTC�u��,x�֨���,���걯-}rB��U�%�Z��Y���g�#+A�ַ���5y����Od������3cp�]୩��k�'��wIr�ps��$�+W��ct�XX�k��
(n��ݷʶ�dk�C����J��^=d�(ז�"����*�h">G��P��F!������#E�ܒ&5x�I�fۭ�r��lV;K���f�U ��Ӣ���	h(\a�ц!���0��Ez�(��z����b[d�w�t�w�z�2P��CM���7a��z;LN/(�nZ<i�5��[v+r��Fu��*`��ľ��o�6n�͑nz��Bh��|l5z*uz�VR�v��џ`�tc0G#���U����(�k��)5���F�z�9��EO���zz|���k�>X����x��������ޢ�Á�"�F��\��K)T�pp��.�r*̒4t˦UtWm�19>��W�B#��7�Ұ5��7.�\@EaWƊe�����u����]
�Z,2bq����+W�O�{�>���#�I�Af�|��y��۾�����1�E�#>�<I�ol^�U��:��FX>�7�>�I,'�U��]�L=x%F3q�{�7�++JE>�|pH�~��{��Ru�o���U$�Ҥ���G,��s{�]�0�R�.�,�'�3UL%�"4⏩�lWs��H�{�BK
���z�̖l��\p#cܯ��:)��<��Vj�ޏ�&W�lg}��A�}�ٱg&�(N1��$��Uٸ�`�'���T�A8.�w�o�l��1��M���^νy,������w}γ�M�Xw�R�e��bi����>y�ٗ���`��@F#�4ڈ{���Ud��S��{�'hfK4�x�Af�u�ʂ{1h�n%�j7�U�&�I���b1xk���_0(16Q��|X�K�CΘ�]+��E��e�7�˖R���I�����z���_y
��'fe��Z�q�H���iZ�7�@�|�s�k}H���7۽v�7�l�[D9��͵�yk�t�����g;�lnP�XF�\÷b�C���7����s��uG�h��S�a]��n�Y����-���*T�je17F�%�ANz�Oz5��î�3æv�u��g;����Y]���ʸ�tKt�|�lV�������Z�P:��0:�Yu���1�&6��l��jܷ}m�u7<Fܐh�?�U�f�]���t�i]�ӽ���A��m���tڎ��.��0����Y	0���q+�G��C��y0�yAQ�'���o�;��M��K�J#��1B����Ѝ�Z���\��U�2���R����8�	Y����8����H0�z����}�on0�vf���j"v�\�xt�:N�ϣr���\�s��\q��ى�]���7&�.HU.�-�zxӚ��;\s]k�ӲN�[�Mg\���`7i9Cn^���q���ռ�L�v :鞊�As��3ϷI��� �	эp��{�{e۶4H���ǒ�v�^�����qk<�Y�Zw��ڳF=Ip��\v:l��3g��m0I�|7����k���v̻\�p��,��s׈��p��l���.M��D�^���P�����wY�F'���mŹՇ��q���v^�L�:��tzk��ry4����v�;7)��Z�+n��m���,^��YӲ�r���nu痵�n�8��ƈ���C��e��f��S׃o�7�N�oq���mʾ; �e����;{;ڏ1uv �NN9�aCqA�錙�����`^1V39���NO[����	vv�׭��0�'�1g��;Y�D����[v3�c#Z��ܯ��l�<2Z�uv.�ۡ�v��bmݹ���g6�ɴ�|nsN��m��n:Sv`�x�Πvn��عz��'g��cV��e�U��qZ�ڻp�{���]A�Cδ����ri�k�0<�d�����H�B�O\�`x6�ncslޞ��1�ɧ%�U��"n�Y;4��+�q֮.%�2a�����NnLY��h�d�qpuƯ
xJG��ۚ�Þ�����i7���<i��6�+ "�c�-�R7^.&��m=q\kF�u��;;��'�(�s�Z���Tۥ��l)�c��8!{��ѻ\���s�����Q�9��ܕ�[�=�R5��t<Em��ͭnʱ��kg�m������N���q��X!���9��q��{lG���@�M�J>yw<�nb���#l�������Îx�]�VnL2���x�k�xWc�4h���ܶ�nc��O�E��nj�:���9���w�l�,m��t�;x,�u��-�g4��u	�v���m6�b�[��!�S�ܕ˸��l��y;A��h6��WfNִ���o'Y�T�g��#v2G=�՗e	z�RO����6FR�6��ٞV��@s�'���.����<�����X�b�i�棕�]��%���7��N�n6-�ճ��m��p�k=����Ț�sɹq���p�m$�ͥ�k�rv+[�^8�ر���]ۭrk����{E̼��3XE'8:]�j���%>��z��;�}3������'��B�jO�kK;�����6���y���\��Xq|P����ȜT��j��[������C{��!OT�;;��n]�۽5FbqWڎ��0i̥�T1�罒����f��ιv?�;]�#�����e�y��\�D|���:�Y�#)�����e閅vi�����+�4,�~�>1�d�5�K2��/��0=�"%���q�f{wNWA�]]�7�w��=���kԪ�><��Ӿn��ѣ�
į}AScVs���F��/�Af�y<��ƪ*��-[��P��Q��Wg.;��M{@��S�\Y<�g���hː8��:=�A��LUrˍFo��C���x[a����P��t�yI_m�K�㧭�ծ�Z|p=�`�N�v�k�΁EB����-���J�U��_�`�[��D&�j�ym�Vʎ�󞏫���՘��4̎m�u������s��bb5	�!vu�p	�w���a}���^w^��9؞�}V���e��b|C�vCa�'�_Y�Q�9��TL=��ųGY��Sxm��_<]�8,C8~檛�m�f�L�>y;5��BSj�xja�̥�q�w�3
�Í�W�6�t��΄C�B��D��~^�c+T�Ah�Ϸ�f���"+�=�wԄ�H<,Wī�D�n�r@5�o��t{�qFA��Ϣ�$�����N4����X4#vj�U��&�/-��̧y��j6-ؘ{O@TfI0�K�B$݂nʯ{F�3���`���N�F�}�}��j�^�[r��>�mO�=�#�yj���u'������_�ͷ�1�	WL��-L�E�D�4�N�n�P;=���۝!tzf���&8/i���#]��*��0��UՈX�{HgI�×@��i{��i'�/�6t�5{BAG��G�!������D���ݯ ���v��WZ�5xO�5|�ګ�����l�d����!��ח��U)�ݜ;��Ea�:�a��8��XZ9&)$6��H���*{���+�O��mt�G>C�b:W!=WT9E���D��:�3q8�<��L]�I'+��3䆆���cޘ�\�1�'TUD^kλ׺&��[X�V���J�=ҡ���/:<~�׍�?d��ce�4�1�S�k��2�o�bssM::Є����~��_('�rIpm��#��|U��\�N�Q�^�Y��Ѥ�v��^�� �2�-SK92�[	G�8գC=c�[���|V9N]28�84�~��X���jN��c��2�1egg۬я��ǥ��l��Ǜg��&�x:d�Pr���W72����gyNV��kd��0�v֞��������}�m
1�۵�.�'/#ڃ7w�`Xryp�4Cq'6���Z�i�zׇ�}�����1"	�;O��0�����?o�t吾�\Imw�>�>�%M���W��O_і3W/$^���eY�R�b��~��҈ʾ,o@CpI
�p����u2j�b��Y�O�*��>>s�f1�
��n�ҧ�ƍz���xx�+rU_�0?�fI� h�r�Ȯ�Fn�=���x��l2�E����azo���i�	)aD�^�⩩��n��!ۋ��ŽLL+�����R�t
_:Uǉ�%�����/��l!��1��f�_�6��pBk��ܡ�z����m�>�(���$�rZ�>FCQ��g���@�̫��8΃�{�ś�CV���z�Z�h����#�3�#��:�ۜ|�~�-������B��U�791><Uq����qv�	��'��#v*��q�#��ΪR��ogLUpk�G�<A��x��5^�*�,��г.d�\<B�N�:3[0�3�t24ҍ�Rr�����M�J�W,tͮ�+䐼x��`d^Ӣ+��iȹYw���ؿW�f{Fg�b�9_e��g+q�@�H�)"�.�$&F�W+=��������~�y�	%�
��k�ۣY�0���g�k�c��w�Z���ZM6O�O���E��.�]5{��G\��8́r�e��"��D��Z\7�������{_v�?AnqQ<^�D-�Wp����T���ޔ*����h�U&mQ�+�3=�bJ��A�%H�=�l<�A���v8�E�N]�ߗ�a������I�M�ʰn��c����4U�:dՏy�M+/&+^+�Z��:�{UYz���]�D��-0�,7��4X���YѺ�.��"�.�ܗ&=��^�z���3��M�J�[�g ���vb�eʦ2��c�+��\��L���1�C���I�g��9���(�ݴ��cO�J�j�GaW�>�R����ؙy�ۥ/B-��u>�`�t��������ۦ8�����ظ*�4I�t�Cm�� �j�8��9�O]���dz��^�+�(%0��x�M�U��X�#�����.#�Q��UP�hRJg���Nh�ѿؘ����V��Ud.�'�Z�F�[���]0q�6�;���²�YY�_g8�f'!F�%Ȟ�Ė�;������>0[ϸ�=�k�+R�e�<��hv*���2����w�>�J���l���23ͷ
i�#D!$X3�tNWz��r�Q8ʹ�}ޱUi��J¯آ��zu�͵��Z����>�M�ex�>etR��,����?�J��T��ØEW��ɇ8��I�n�cr�e[`3���+�`��JB��Eի�U��%�g�oC/��|�P��MV$W��I�!�)�)ш��ǯA��g�\ܕYRu��O����eR(~�_`y�F���!&�J���r��!@���o]�<�2d|ݣ���Þ�Y�x�v���K<�.�W�u�m�mO���3i�2���ѺX.�5�8���U�ڪ�[��ܞ�U���ZY^Q����=�j��G(�_[���K�8�e�a����
'���ߋ��ҷoɚ�-ֻ�|%�;�� ��w�z�m(博��|r_\�Q4i�
�cӜ/��Ve}2�I�����Gd?N��f��l��=����x6La���*;�����2��*JŖY�8�Ed��j9�Q¨��jwT�9#q4�]���fU��	E����L�7 ͦ���T��f��Hׄ���h�d�K:�}:h\�?v���=\�/D���EB�3��<o۳S|��]):<�]|��7w,u)�(�=�]�����O��^.8Bq($PE#�몀Q�5w㣼�6wٔs��z	5�+{H>��=�K����tl U��B%�~��fL�~���8�[ܸ:���&��7ɰ{1gi���mT"�	�����)Q5�
�-�����Z��4s��]��b�N�n�!����6���+�쯍)�l��}��Ԓo�K�t��q�5U���U#��	mw>ȸfm�9���n��	�;�6|�1D2K�x��L�9j��H�h#�>�E]Տ{.�'��{,��L�&D�rA$�ƛ�u_6���k��6���ڡ^��Y|ll����!;�\5��Y�2�1�3�\������u�Zj�Z-q>�ѝ����W�N�;���sѹF��D����t�vg�s�5�%��l �;�_(\M��G2D��:M��l�<K�'�{����V�ç9��0S�׽>@(����J���;|���6D�7-��A ��O�%��8�f�]�)���*�{=0�Y2��_������ǧ�SBz�G����z^GLD=W�ὶ;�.�"�{��,�˃���T� �Y V��]��b��K��]�Ӛ����dc��4T�mD�2�M�8�#.P�Uf�}oB��X	�,��iU4t'Sq[*Ȩm=݂�%O1�U(6~���rl�Ϸ��Q�%�бB�ӻ�!��y���%�Y_w��ѕ&��ֵ�K�hW�&�Ր�)�hT������P��&zgU]ۙ2�kYi[��	�@JR7f�.�ʻ����^_xɽ�TCW���=��ɹ�̪�U�e�I6[>=1�z؟.�����$���l��R�����������{�+���U�ZdF����lN�'��֐z�) �ۇӗ��+l�$���;V�6x�eY=��C,0k�7Jf�#q�gCKdZǜ�����HR��j[����/:<�j�fz:8��6�9 ��"�H+-�Y-�~*H�u�6A��=��q/�T�����k�<�)�T���O�/˭��]�,���"�~��G�Tt�9�8e�s\cz�6:[��vz��g̹z���҉��8IZ���,���v�74�us-����3Ϗ�V�{�'A���|��Zk�[�^�l�����l�֐|��on�f���a�!A��qƤc9W��������i����a�[@ ����[���(�)^|���hN)�5V�3}@��,�5�v�P�����D�)�*3$2��W�XC�2����7�Xr	�,��
��Y����� �g>�J���v�f�&V�%2�I�)ѧݿ1g/2�<�]��w�M�.�,���>�c1��+TU�諏;ێ�{�$�W��p����C�뗽P�D"ڌ� �����(�#�ϒ�b~G�����4������8F
�nJ_�W��!�X�w�'+��3�:~ƅ��9Ǉ78[ ��u��8o�����=ؕ��=v���,w�er������nL����\��Xa+us�=���ΓO3/�O}���Lh�E%�Q�V6��;�JN�\���ɻnvpGkp��]������,�n�6�9i�����O��d�y��s�M�\K�.�U"�����y����Tn.��7ex���K��hCss�vܦ�tv�C7���N��I���5��������n����8�Ћuͱ\���X,�<�NT�*4���A/XXi��n�.�p��[Y�n:2�����)5F�ӂ��
PNH�b�X��,.��lv��[��#�l�޴���e��f"P�D�cL��M�^p�Y�,��dheM��a.�{�^�wޥ�D�`ꡔ��Z=�&*!�8y*��r�#)7�/�=Ц�H7"�C!�,ﴼA�
矼�_�ͽޗudjA�>��`��&5��+�<�C�R8�"�r����?v��݃(v�'�q:ݥW(�$� ��Q7�}E��كY�q���r��[~~�"�oM]iv���C����
�WT*G<�=x<ٍ�$FnE����U�L�r/y׍���b�<7��4�[�}���âŊ�2��S�=�z�זO�d��>T!m7�&R��b�nLUٜ��o��$�˺?*�Cyˇ<e�s��KТz�\缝�i۬&`�ѯ޵�q@`ۀ�	n����.� De3�n"۱�n��.}gx������{\u�_��;�Q!˹J��%�y�UJ4�-��cc���˃�~q����\�	���s��І�}�͡=������fش��׷��6�����}5��Vl���:�vCX���G��Y"�ڎ�'��.�����MI����V���p{z�{�r�}�b)�'�Q��]���QR���qn�yl��[xUAo�e�Ƨ��8$Si��x��W/���7�oWq"�{�_��͈r*Dgv�J�D$x��xiy��mW{p'ٽ|}�wi/'�6R��d�Ґ�z�Q{f!I*��ϣ��9M���uH��x�yo���|���Ifs<��)�Gm��玭Q��o���b�i��	B�M�D����g�ë��bq�1��d��=R+}��ϭ7�
������hҎ]r	�^.�A������N��i/;�6n��y;�y#M�qeN��zx���f����Q���4��ܟs�O�=<�Naƙ��Ɋ*��'�C��J�3u0kq�ȁ����߉L��ُ��j �^_@�?E#��y'�f��}~-�1��nvd8�6��m�M�c�]y.�ݽ�8�~���|��2��y\A�cL�$l)�
�o���,Þ�]_#��鈿r��%,��xR�nn0k��\� ��yu��*�3֪O�вn݈_�Z������rc�
��j�\;�2U���8�t����eX��;|=i3FF�+�Ozg������=����Z�"�k��^��ql�ζR���z�i�·;.Ky�/��L^2�a�`��46f,���b?��S��.��WZD�Sw}������u���qs�`��{L���HU���z�(�����l����)t%XsU�ؽ��,-�KL����m�}����.B�zw������S�NV7�G@�oc��P��TLq��˱����j��֞��H��:t'���O�m�*�H�]�{ ���(��1��ˣ8_�c�tW^]}�j|����C(��o���=hn�ˎ���C*-�*U]���-�ҫm�b�G3݊`ĵ{��_f�S��ٺ��3��� �WC
���ghd��V�x[N���$�v��m��9GK��]QQG�т�l!�\��X���N�2�zg]fg��Wύ-aݪ�ƒ�{3��Ggh�a��\�y��*V�]F<���,�=�Q�ow�>a���=��;Z��u�Y6�Ux�� ���Ͷ��mJ��W���0'O^M_��T�����d���*Ԉ���"����T�*��F@f;bu|坏b�ji�j �R�k�\�V��F���H�X�5򁢫��$��[�U������s�Ϳ�lۯ��=�]����n�x�)u�zN.�;�W+��X��;X��b�u"z}��d��U)�|�Z^�d㎶�zH��S1G�>�x�_MR�I��n��j���m��6�����a���k�2ѷ^v�/.��5_z<��"X nFJ]�t���
c#�+������u���|�é��bi����^�v�OIRu�%׋���.�UH7>;k����3Sa�����+��y]���6����{g�Sd;Y�<b7l�f�1��7/=�Ʈ��7���;i�n�B�
z=�M�0o�>��%�m���$���;�V�ѭs�|:N.�H��ç���%�;$-q}���vw|�w������]��(�wo�m��n�s<;wѧ׭����.�ط֊������3�tQF�/;�	,��y����j�J�>q���ˉգ�c6�?J���7��ļ�y��dc��p:�^���u��*�3&}p]o��B拽��/���F���a�z�y�x�����VA�8Q	��p]yV�K�J�����׊����K�n�n��!!��C�s��)�5��*�L�&�<��>{4���]<���z�� �ܘ�9��b6w��S}�o��XeIs��>xC#$���˷j�6M���R�͗p,�(v�5���Y]#�zĳ�������^�>Y�J��C��/P�����9:��tw:��tQp[6N7[�!�ܗn!28�ݶY۰���.��z����<�4�b���[�ze��I��ߔp����*1�����0�Ɔ�k�~p�䢰�J/gA������7�$g�-����G���.�z������{��]�"!x5�}O�(�&��
����ѫ�g���`�Ν}��u�� h��q��ȥ;v�8�xuz-�����ܨF���T꫃|��[����6W�[�	X��Sљ༩3m�J4�yڴK5^�}��b�=�zϟU�rYܐ����<�1��G~��}˞V�v�A�Y_z��_`��^-�{�+W�`�>c���#r�-�71XK�#�*��U���s�r�.����p��ȩC	gx��h���3�	7tH)j�y~�Uw�hE��u���ф�P��d*����Z�8���y����o��>�į��3��q�Oz��´��X����J�U��'�� ��΍��ts���vxb�j�c��V�VSR�1@�H.�[Nr#��>��&�  g+m���<ix�a����7Z�F�2��+�{{��;��i�`շ
p��	�vv[n:���ڱ�C훦u��L��lk�^,v�n�Sz���r�r>N��ৢl�[;�L��n�ry�w��||��g�w^E7eq�3�/��������l�.�v�7��������c��gSۦM�n}.�Ǚ�)0M��WH#��X������,ǔ����`������{��ьI�=���L?e��[	��W��ʓ�߅#I��Ar&�RGU�E2���^+�yof!��D?	t���X�^����̗��b�^;��R�'�:�Z�vGz*�%>�%E$�>�\�)>�<�B(S���hfyx�A�Fzt{�V��F*����.)"���dhH�-H\�80�nR�}g�����v�P�9b���؛]��P��q�z�f#����k~/<�P|d�+����:����9����Q����N=FN�Uz�W�2��0s�ӯ��[���h�t)[O}ƽiؼ1'q��V�Aj��ܟo�ߺ�d(�m�.�m�<��W#��l' nW����,�!>��ݞ�iEn�R9G��y����Z��	��<�a��Eys#z~�T�J�ػ��5�٠G��zO8��Vh���f��P	E!��:��r8r�
��k��xo��Ha�P�t=�
�{�|{oCF�9fN���Q!7a�5�I�]w�G��#�-�w��cNگ����Ϸ/p�'7���yӗeyP�"}��zr���Y��i�/#�ݞ9��X���-~ó�|RN�},z,��RJ�耕܇��K6O4�	����h��S�.w�7i��_�(.�3�����n�+�h��$�m�	1ȯ}��\��⏤�a���
!k����e5�����L���,Y��*!���	���(V��"� ����,��1�/��D�|߫��/��y#LQM��=�S(��ޱ^�Ͻ��nCMel�E��+o�T��>-?�����n Ж�-�k.SFnն�H����� �;����i�j?������CB��OXT)2��;��߰�-��������jϕuz2�;��V\��w����⠖+P-F�Ǐ/>1��ggt>�(��4f���Tvo�G��b��U�u���8-w�8�zQ�&;�zSa��^e�P ��BX�ے`Ǒ��0�/X��{���:�k�#��_9��Y�>;�]xe˜Kz�]�ok"����9�Eu%d�9gm��ln�����vN}�i�܎7�^Vt
GqI�%��a�L�)��=��NyyO��5������-�#*�}~L��Pia|6������p�P���o����a���H�X�]���[��S���^��UJ���� d�QMFD$��GD�u\ُ���:���ʵ�u�^IZ�U��H��'5��OϝmN�-�²�w&[�`;����N�Q^�c]Q1��ܔ�;�38�)�z��uP���Gf��,h�.':�D�g���o녤M�<�J򕛪(�� T��ٔjRh/x�שW*��'0��?IgX7^�N%�W��6��.I�^EV?��n�e�&���g����9M�qX��B���ǲ;�o׷{��*�nA�Wd��?8{1�Ѩ�22�&�
�T�?iM��f�4��5{�h��{e۱d;��[��:�8�Rk�Ŋ����p{�K>��-��,��V�����pRػ&Ug�bȣ����{��J�|�p��U� *��:��ʱ��JY�ΐp�+rḻ�;Z�p�7�(�p�����˹&���5��K�%Sv��D� ���Me����Vޛ���b �����!u�W�2���O�����, Z��i�ݲ���(��{�=+W�LWh�~���Sf����G��r�+)��s]����ޙ~�Σ������^��Y&����4�b0C��B|�rD������=�01�k�ݑ����5�qk�cnq$Zq�1�^��o������-��@��ó��ܪ ��&Ե����F�s�#��Ԋ��ɚ�='/i��XJ"(q�=��Zn���{`��w��Fr��|��]%tE'�B��V�|�:X�k=g�7�D�O�L��f����p܄��)	E��f���UFg����D&��=w�|�4����ssz 6������M�J�'��쳅��c����FG]$nZ��<"gd�	���S�q�f�x/H�ʎ��bB�nf�2J�����6�_�V|�]�m���X���_��O~Hi �c��z){:�=�Ja]�Aڡ�}R��zS�/<6!HQ��mw��L����T;�K�SM�Y�J�d���m_�{���jVj���aݾ��O��2z��� f�h�6um5;=�O!�tEY��R��W��]&U�q&0�쬽�X�zv��UR��G,ccm����]ۣ��cu�\\��GF��#�;E�����Yw=��l��;fۻp�ѕ��m�&A���]=`�y�[i%��Jԅ/���0i[1xb�����v��ѸN�9#�D�	oU�Z"hP�0��4��Q�`�ku���t�xm��7<s˷[����ۙ�y����vx�a��������]�3��zE6�!������sW�R��z6�F-m�:��{��q���IЋ�2Xq��j����x�,��`�m�fZ�<f��
�k���0*x
��Y�x�1yΖ�ٶe���1���$F%pWv�A�����U<��|�!��X������=W���\���T��v+	��fwJB�h�p��a�H�N�0�4�FW��wa��E����L}Y<W��.
m��E}d;�U�1\�������������Ě��`���=߫,�<��ܫ��fBߍWI����|}���#��oם ���R��˷��=�Y�M��+�/���BP-#���6����<}jϤ���6�O'��^��ډW&�!��jo�Ď(��O,�w���fG6�q�ιu���rmd���� �f���f:�ڎI#ZQ��[D"D֤$JZ7���5�a'<8�ې?}���Ǌ���T�?��Y����9�pY�ϋ�KW~7�Jj�B!{�C9��}{cv$p�'���W�u�qGs�.$]AM�P)r��Am�,�L�'k�k���[��{�&�}���t���)�A��ְ��'%gP응�&�����|�ĥMe1MJ�c�x�c7�	��� [�Sa�V���S9�/c�uS��~�r���N��3���*�f9�{��k��Ҩ����?P���sޛ=��	����w�n�H������'�A�Hk���􅠆*�᳽j=;�5��î����}4n"�R�:pU�=�Jr�����oz�0� �9V��-`ʞ~����`��T��RT��%�<�4NL�3yw�p�N�;�fC$1��QQ�;�m�Ok�ei�鳾+���x�a�ʴ��t��G.5��g��mt/��T�r��:dwa��ѫ�z��\m�y�˰s�L�d1`0�6���f��y��Πhziݬ����~O=���̜/������UNL�{��7t�B�v�V�0uaH���f#)�tc�<iWO/�[�ɚ;�9=�Է ^��y����O�M���\��G�4��~v'�MT}�ރI�	Mx5c��jU�Z�!-�'âD9�W.�`����>�<}�Ss���l�k��HEn)d�2�.vw=�z��t���	�y{�f�&���@���3�Y�G8H:G�5�l���yz��}�pu�/��x��>ӿ]نh������B(�>P�R�J����><��г�|�{�iW��kE�%�*�������I�l�2���~z�6-�ޑݟ+L����&�7�C��~^��_o�&X$|D�c'/pYY=�:��!�a�����&�W�6�u9����#���(!Ѵ�	`�Q�+[ts�Z��;cg�tmƼ��<�h��M	l\W�r؇�p�܉��^J��Ͻ�t��ƩP��������0�)����Vg����^g]���������D�V���Gwv��ɳ���#���,��^?
)�G��P�R�.�%ԧ^V�����N5��0��H� �����<�0r��e	�u��j��$%�c��U܅3껰K���z²%��}�K���|����1�r�L6����S���`Y���Z�x�m� 1����Q#��mY��{^�����%e�_RI���^=�'�{���#>�����޵���|*SFy{������.Uvk�����*cJ�E Cǖq�S��.�ܤv��)�ܾ:��ƴ��X/�6M��wT�~_%ho3�H���(ح���'�أ;�뼤�� �0r��)�}=����Q��,�����Mt����DǬ�޾L����9gZb��4���Uq�J7l�-�sڷ:�l��&f\��nroQkM��(KREB"������uw����n=���!��xq���U�G�r_C���'���$��߆�'&�D��U�HH4 E�"�֫j��A�p�h�h}�Nr}O<�Þ����8�sZ�����$��k�~_|/w�{�X4����%�����Oc���W�����U�J�w�V���T�c�X�=��:g�W��q�[\}�1�I")�uf�+�]�P��Eɯ��}�׷�?d�^��\,A����W�r#�Z��Q�z�f�ǯ3)>�< ��c��Z�9�IW�R�|�x���j��w
�3Q+����3�u����P.�g�˗T�o��]�d�V�N���=�K=��	�=�/�������v
܏�P�>l� guʽ��ؓ*�T{c�}����ŕ�<��l9=1�c������d�����q+n�nL�/�aQ�3�JoLi��`��t�ϗY�6�:��so-w,��~c-t����;%4�R�`�V'ov�p	(��"�<��n/{N��Q�֋Ny�\���͚ˮe(U:	��X���Xtu\޼�k3�
��%��}A��\�8��ᔔ�t)�m�h���<�h��	�h#���t%I�[�bw�΅�p̜���=җc�Q�7��[�xCIu�X�\�t����<�=ҝ,��^h�O�J�sA��3�U쮻���-������{��:�OY-�w&]̾B�9zs�6�&��Y�@�B����[������P��ͱ�c���t���˒���u�����P6��z*ϻ�Ր��M�s*ؕ�チ��^��L�|��XA%�Y����G�v�v���Ŝ
֚�:昶��S��/v����4m�{�J��r!R�ہrq���~��OM���r�
a���4�>͛j=��9���
Ĩ G�y��఺nh�Cg!ṡ��e����"�Gq��(G_y/1;ϭ�h`��t1����9��`x��s;rG��u:U�%�wѾ{�1�����q���Yҧ|N����S˷|���v�3OˏK�]q����7�b�nɇ�T�����}=�^�����cz˛�G�z�/j��8X��+���Tuj}�����̉�?�a<;�@O<}�r����Ś�Իu��M+9۲�<u�id�{n{��=�4���r!��ԍ��q�oj6�1���ݬ������u��eӴh(�똥���������'<�@�V�7=�pl� a�e�y.g�%���a��q�0v޺��8H���9�����k���C�j�]��֬FX�Dv�]�s�B�r=c�U�<�a�䝷��&�� U\h����a��n���\�a���V�l��5ڞ��6<]�s\d�!��n�+<6y�]�(�Ű�����h,KZ��u�Sb�W\9��.\3^�[�|3v���r��rjq�{q�8��v�K��N���v�}`C��e���n��=��]����'�uk��b�����Pީ�-qrn���Svv�qfp�H���n��s׎�s��vyw�P��^�z��H�<�GH;�4X8n:�6%1��ݻp��N�Bm���|GE��4:
=�lq9�ܔ��^�p�oM��� ���n���@�t*�c�쭹��t�"�8k:���ö���ׇsՅ�!�:D��v����p��I��I"�y���gctu�5�q��O�ͳ��rWp뷏c^�q�dokk��^�.N��d�x�������;��<;��\t�{n^���ȫ�����W\���c���&�u�ڃz�mL�[�5:��f�g�t��P�ӎŝ�'�۬�\�̌۞R#v;����נ��<r�n1>��ˈL�d�d�m��mq�y�8�.��*mm۴kf�e��ۢw!��{�q���WZ͖�ڸX�kH���bhD�V�R�B�S����n��Ni�v��.w����*��t��˷I������u9�hM���y��ݔ���u���3�=G+W<k�+���g,n0��3v��q�k`t�t%C�T��^:�z]���]�l1
�f˞MǴ�{�]��]K�cv��	p��j��5g3&�,T9@v�n������l<���t��y�pӺs���睃�֡��2;Ϟ�H�]r0�6䣞��m��m]���w�㮻��/M��S�x�6���{q�'n0�V��޵n�l���=��l�ln�iE{!��'s���&���֌�w#śm������]���l܎�r=���y�Uq�!4�E�'kq�n6������Y��pq�ˮB{��u����q�t�<8k����cZ:3���DA{X��/Ta5�@�'i6x���\�d�8�7X�筙�.�ٓ�<q�[��b�;٧�(�	4���'�S}�^6�S����M��=3�&���1L���Nۥe���6�m�U�O��DC���l�cpb�M��\=�J�j+�[���q眴��~~~W��:�!���W�]��fWmM�,�?(H^S�P��O3s=5��{�[�ˡ�^���㽏y�.a����vy/_��)�����_��x�-I��w���	B%(��q��%�u��p	����xu����aħ�u�^H̓���<���+���<��9�.?Y9�W�,k7����������Q:��{�V:�8Ֆ���&7LU_'Aw�ʾ�����F���T�|vcš�l!�M`�Vh�
q�6���:���7����:�Ev�0]=;1����/��u�Y����m��6���v~�|��:��P�z^����	����\�{�޺�'�خگY�f�'��= �E .$[��N҆��ީu��D�g3uOڻ">&[�pt��f�vkO���U]-�x�n�3n�MNT����\��ٝ�+�z�sk����Xh]7���{����*E���0��69d������-\$��	
��#B$w��5B�5�w�LD$F�/u��S�%����~ ��ܳR��x�^�po{b9�J��tA��FP�HБ�qU�I�k]��������>�:��nP�~�Jɓ�TL��q^t5��Y���������[<��a@>�`���"�+�Ke2v!���1O���9n���2G������{*s�ۦ�W�:;�����/o�������m�h��4�}������6�8����nF(���۳լT�Ջm����sۭ;q�C�u��3n�]��=�5,�x����������v��I�]��H��,�'V)�Ƙ��j��y;��{d��n�����s3!DA���{ScVr�����M����Wl2n�<Au�O#����2�<�*�ݻA�y���aވ�B�H8���kNu*���y9�T�ϵ����k�.-s�`�lw�U�I+&��i;5Kw�o�&��#������`��z:ɰ�3��5��
�|ʹ�e�+_��/�SC��-s|��x�X4��2��l������N�v�S��
७��{��^`�y��"%�x��M�u1�#ٳ�?#t=��[&�C�������$�\&4r�F�Y0��{��,<}���5�����ϓ���^mQ}nA��\=��*X�Y#�76wQ�Q��e9�Ƒ�ɰ�����%�<[S�8�f�h=G5�!�c
�"�+�Y��v� w�f�ٸ��Cy{�Yr�g�L7!]3��M�����=�ڻ[�������(2�NH�^L��A�^��P�y�`o�%�9(���ב�27�z���;~c��=���;���׽��x�ND1[J�e(�N.��Mܬ�g+����|6�����۷G��s�v�W'����q�=2�װ[�z��	]��� ��B��� lL��.�&�n� ����v
����gz�ԱU�*əu^���3����U�Z�,�������odǐ��be�q�ޙ�D���Z5��$��̠�ǐǃ���)���6�t�NԺ���ڡ�1��K,ɪ��e��cW9,�����p��<���W/碳���w�����N�õޔ����D=-?�Xs�G~_ߧ��k�2�s��ع������8㵃'�,���F�,��-�n�r��i�j#<6tr6,w{(��}��U޼w؎T=x����wν�n^b���$6o��~Y�1&�A~���ÌG#i�`���\��VU�N+2�%��ߝ�q��>k��~_?8��c��,ez�{_+�^�d-ϔQ�N�X�����h܄�<�q��DD3����U�m���3wj���V�^չ��l��P�0q� `bE0�c��2�;�\X���z�4껾�k\+�^��[J(�*����|K�A�<1Jəb]B<��O�!�9�7�3��{Fb����SY��6�]�����&�L�����D��xo���j�6�����4��kUlR���a���c���Z�x��dH2�r=w���O����YXk�6������,=��	�x<������&�E��-�3\i��n1����V-�'��ic��;n[�I���0��-���f<�;�{W�xg��p�d���,h"
z{:��ǝC���s�\q���e���e{s�+��עK�ak��G�Xr�y]�b̥�N�<����k���l��O4�^�x���[X�p��D��6��OL�rv�mn(�WL��ݶ9�g��k��٬�9Ў�q���w4Y'�rY���7\��a!z�8���v ��"��B��d$V�m9Ⱦ���^�S�W����(��Z��F�)���z�g��w����Uor�Wm�ɑ�3�f�0�_t�D�|��W�Яg��r��^�^U;q�Ğ��r^t7�X�t�=]�����/L��6�]�HX�&L�ʑ�A�xg�{�׹�鐀�<��nҟW�F��'��|���p��s�K�{�l�OS��h���##���_����9bǆe���S�2Z~'��G�{�o�d�������~P|���G��,Ŏ?d`�#bBԇ��iw��lfe��w�!����L�D�Vi�h6�}�W�t�t�0Z�����齞�nW+��Qu�+GU�`jT"��$D�E�{L�=.�{�Q�!�/������m�hI+}r?�-�8j\ʞ=��*�܄�YG�ͭ�7�p�դ�G��TRo���;f
�����=ּZA�q�9r9�)C\��<��������I�������\�����Kц^):���(L�I+4gZ	*+.uVj�j��zlֲ\��[�ϓ
a�n�d;:��Go��Mꛪ�RD.�՝p_���M	�퇽�ta��{{^�zH/f��<��3�ƛ�{�U�T����Kn�5<[X�W��d�'v�
��:��������<��!E�7���[��IEk��Q����/)�ח�4�_N�(��œp��f���E��'��x%�N�]��<*���%�}|�`4���n!�<��»;�a>^��Z�w�\X��g�yö4�א�o�ռ�^�}��O��y�ᐕ{&<�ޱ�wڝ��&�q8���]���s�s������q��7&˵��*l/�)gv�ݹ�a�9*�EvI��V�A���8�q�>N�?bX���ū������[�d���ݛb�G�')��d6&�1�W�Ly������:�c�\\׽S2��]�AK��~a?����U򒄳���g��č1\�5��"Y!��Vc~���PXe��������,R&��ծ�[Q�Q0�pC2�G��O��W�wDu?���0Q��MX�㩞g�j��wڻ+"H��[�{��3�τ><R��e/X^g2���;,y'��p�����2�n�y��W��1K�tAnz��yJ�%)�^�����/s_{/������g�saU����a���!�R,Ij��a�����vH�H��|g�t��NIy��x&>U�]R_��Ň������������H�,F���3x�5u�ggt��)��KK�WsF��u����Ei�r�Pi��{y�~̞��q���Ւu_�CIto�}un;T����ʕu�b�����,�>=�hm���� N�Vw�(��g��f"�ޛ��(a�P�I5L]��X,�f-W�tɝ�+�]�sJ�,f�|�ޚ��fM"�>h���9�1�t�J�T�7d�\�M���^������N?=S۩���~���8���Zd1���=B�fV����woe�����C���5)N�3��5��z{%�=@ja�=k5f!*�7�oD�/7���o��J��/qĺKq�������u�I{���"��i�6���}�/���=X��`(�&"�������������U~��F��p��t0�\m;<��;n�gJ~�G���hY}�L$��(�܆)�ܐxg�T�	���p-p�=���,1[�9C�Q����6p7�bY9�~>xp:��Gꕞ�/貈MW���}��b���]Yq���O�����c��jt�p�8[�II�s��7�Ϧ��#e�^�C�aV;x��(1�s�P��v-Ra�� к�y=��u���5'�qWoU��+K�"0BbH��蒛�~��w�Ux�d����r�NYh�����;��6u�L=�h׼����ka�ϳ�#hA���r�ͮ���f˱�]+x�Zs-��G�.�FT��5%zA�S<�ɚ/i�z��]�݋ m�u^���Q*�"�"	�72+�=��_b���Z��3��*�W�睭鍗��-��C��z�C{�5�t������S�Ix.}l>:�Ҏ���uj8=k�K/Bޛ-u�	�n���{׆�߅���B8Y��@��ۣ�t={إ0i�+�8&�ط��K�(�;��Y��jP�d]#���\c7������Jhx8[����u�������Sc+�̏u�s��c��t�{lP��-�a䇠w���N�(:�v��۝��=]�,M�|5lۈA��N1�7g���gs�E���m\۠�bՎ�/c���EW�*6�^M3����)-��dq͞��K�r��Lx佬>��d�ڵq�ϋ<=����C`�&ϊ���;nAl��m�cl����{<չK���H �ܰc�����r�t6������:��M۲!d#�~����N��O���0�u�Ƴ����#n=���a8�nH�p��y{�%�t���|=�D��G�ϰ�V�Z��L�D�h��_i��t-���P����C&������'���)uuUUtw�b���S��!^l{0C��kݮ�j�OM����G~�UqO�5r��X�t�z�JAl@�����wc�r��������uh���,� �7e�u8�����Z�?bB7W3�a֬�����:�?9	(`Pȓ1��C�0�����n7
��6���|��v/{/��^ƹy��E߰Rc�JO��7�TԭW��ꏢ!�IQ�{O��O�$�,��&-�fݟ��;$�g�:��^n
�O͸�jI��D���#�x�j����ofzu;39�1te���-�"��Wҫ�L؈�-cš	��������.�͕���~���j�6�˸ З,b�i�zn�[��ׄ>K��=�����ܹ��i�&�y�{S%Y�EW�:�s9�Ѻ]O�/�be�Co�^�wK�Xo�����s������R�*P��{�yOg���R�-{j-Y���X␍B\��
��UWU���g�(a}�mn����l�*ڞ5oky�n�3���1�����o� k��ؤv��G[�&Q�ÒJ�p�_���o[���a�t�9D��������۸����^����?�{�C�+���Łc-��1kŕ��[��[�K�z����Dk�c+��8��������	?/EiN�Q^��[X��Km�������}�"���!�y��SH2f�q��l�5YP**�5PZ�2jU��=o�}D�pѷ86n���A"L��G�߳�	m�w�׃*��+=~�b��M��w*��y����jD�驪�/q?H��>=n)��v,�&�-��$�����I��{}��v�l�9�k'a�3�.KI�+qg����S��{=�1_-�bG�`����
�Z�}�*�q��
	%��~���ʷ_E'��w
S�Z9y�?~��w��B��[�]Y��u��hҰ�&덌����\�!^���`��q&!��)�wǁ�續H�k=2E��U-6�Ud��w�dq�}����Uq������̞��Pk��k�3{<=�pB� 6��1����>3�����!��蹳�%)������'NN�z�H����C�m�1�X�[��J�NL�d'5���3�Kr��=�\|#�l�
�k=Sn]����n��i���(��v-�V�����3)� w���W˼M�s�4)��ot|���iu��U��Y��9:���ɯC��[6;�ܝ?���Z��K��L����C����&��`n��eʲ]KY�gˡ���s��d�������q��{�F�@ɧ��g�m��D�f����W�v��X�@U�j.X���CX�ag|�
����
�d��9Î]��E��b�-�ZM�u�������R�;�[�W6s�./�:����̽y�0�d��Q�IsWb���,�ww�u�'�zN���k=��\"��3g���Y������>�t��_Nl���3�\��7�x�rRc#��Sܙ�7�M�p��iB{�,{�n�{�U��{��m��b}�]'UQ|�$-Ⱥ�ןe�*�@�β������ �e�����Y��u���1� ���1w���,큪�Ês�~�g�Y���ںx� ��e<��ɮ�NHև1f�5AM��,K����m�Q`��C��t~����$�<9������[�๻	�'th9.�E��/�a*&�� �?�|��s=��Y]���I�m�"P4�gG�����;�o�vZ �J��O��h��R����T�{"�;�
�b̚�����s�tG�p��F��K�M�I#�z��J�9g�*��K�$ ����xT�<��o����r��ڳ-zu8����{�5�#���g+}=]__t�nu���^F��"2b�^��#n�n�!�1q�6W����[\�'-x=�7}{=IT�����\�� ��Ua�*��e��<��׫=�\�7�I��e�� ��'(��nGY����F�����èŗz�hݿ�#���0c������c����g�R��涳3N�*��7�����qI�M�!��d�b��+�+ν��Cn3w�����]	����hǪ����lu���ѥ��7�3�YlYBIRIl5!�/s{|�ھ�;-v������柨�S�t����+�7����둸��o�o^'�X{ݣ�ʍ��n�oF���n��58S�[J�ֱ���b畋hp���H��Qyӽe{��7�˸w���#{�y�J��}�8���ҁ��o���>�R�tG^���_nm�ץy{'���sߧ҉T�͹5�8���KR���.�����v�ju��U�0�mTK�DN*(�Ө�z�r PuRBon�]��WCgDl"Z�-k�N̩�n^w��\�Q��{
�����m�Ӗ}^Xx���f�z$���U��/d�0{0���
8�n=�4r���ِN��,W����ܵ��[u;:�Ha[���>�"]8�09��Z8�D��Py�Ky���=q��Q$�vko��vz���.��^v�fΓM�G�3Fn3,ك����w��&�B �l��>ڕ%_����?&��v����fg�ٽt���y���@���6-�6�ݿ]Y����� A!�HA&�:���#n�='���@G�ﱋ-��V��������^��#���W�^:�����H�T��)�:ax&^�c�ݕyu�GKMr��`�Ae��j�Qca��.�&A�����lT��풄��l�\����s��շ�6f���� �B!"J0�/bn�dJ;kus��K���4��Ӫ\s�UǝK&��Ln �냝��\�El��`rZ��[���6:����*n����A8�{�]@;<u�Q���/<lu��u��l]ۈ�s�1��;=z�I���1.��c��g���u-̝'e�����-�]��;nP͙7lC�捻v������l��c��s���5؞��u��뚅��gf:�O�����:��yⱶ�ٜȻ�҄���ܒdW�i	�C��%y,�;���&�=��t��o����t�DW�kD�+����Cy���5���&4PQ�$/"1 ��޼;}�$���C���UrR�.j����{bCo= ��V��Ϯn����bg���)�8�S�C3�b��a�BV+�>���{�:|�a�y����"�
@��זp�Y��g�h�ź�~�����Oj�7��GT��Zf�&(�Ư�d��9T���7������]
�Ȭ�P�ö_:qy�o��|�fw�x�o��������ޢ�ng���mC�H����_����9���p�v5���ܔ[�-��q�f���A6��b���{1�}[����ͣ|�r^�B�FTM тe�84�.����y.pj����qqu�����ݛ(����H*���nl��[b�wSn�S�2�r��jĳ��]�G�Ry�tw��M���`*�r���@�+t�NB��e �T��}��|E=6�|7���}�ݝO����7��w'�I&��npQ'_q𪋛{�y�ן�9�/xܫݛ�-�V3�5cV�.���<�S�;��	���=91�s{V��}�cu9Mj�M$�+���Kٻ=dr!�>H4�(4���vFZk�-�����T�<��c���\���V�Yٜ_�N�CgG�z�����}��Z�l�`M����f����v\�}z����Y��b�P{�p��W��������x��鶭��}��T�y��^�TǾ%A�M�)�M��+޼g�kʚ���=�<CW�u={~U�uq>C�l���D�����n�Ut|�셳w�f��YD�W	!P�NŘ1pM�q�,�k8��6.��������{}T��%
H6���U�w?W緮�U$�.���|i|�g����~4�I�ը5kɛd����P��yyuvp�J%�╙��Ϯ�*#ב`��J8U��0��h�h��T!�κ�Tf\�.�2к�P")40M]�������"�8�P�w��[R�N�Ftw{�:��֯�`K�ne���,�b�V�ݛz��6��w�&�i�_+�&e��t�9��׭و�p���|����i�O,����၃]E\�J���vgV���c/GA[�偖�H�����7T�:�u�8ɂ�i�m���>��}�K�<cB��Uk��~m��{Ea��3{g�ظ�����H+��W�Z��m�����z�*EV�l��剗���2ӏw�c5�����8)�W䖪K�_��;������m�[�f�y.YP�4�v9�q��ɡݲ��ء4��؊����H�k;�\7+���p<�iuuޱ�ͨ�h����u�Gv����D/}Y�ݜ��̔*��ns>,����%�#�u��{o`󳽱U���6��7�_gӽU���"G���?v>�����{FNQhH�L�f�8kɳv7����t�O���`�����uީJR���c�ǽW�/c�N����M�D�F�I�!�,?<�	{��u}
����m����M��7t�0����9���I���,���t��������Z@�d.��AMכ��zD}�H��7�'�za�ȳ��!�JԭC0���a35Ú�'-c��og���*>��&� �	fp���K�s��{V��t�Ѓ�ή���R/XZ3�+�w���U]&]:匈(@~���~~w�v2���"�:�\���3џ�l�az�c�;O��z���Y{.����)U��_�G�<����vA�5��yX}��ؠ[�:�Rc��͜�uYdB�E��GN��-�i�����FAb���������t�'�|��%��F���mw���/^Lh��P"�M�KO��m
r]����sP{���aR��w�N�봣۞�{�n�f[H+�SƭٙK0r�'�Q(�	��[zO��\<�*�;MA�����G���[����m�.Ԩ(�Q�vv���������c�uW��PD�й���O_������J��N����ד׵�R/�:�Fw�n���g]���k46�կ7o,�mǙ�-�,0�Ww%�oow%{;V��������;�5ݭ���Rt��������W��������0�+���s�<���ɹ�*5Y�l�u�$���{������3�;�.;nl�VNJ��yݮ'��o7L
l�U����[��'��E�n��A��rq]�khOmټJr*�wZ��]�˞ݺ��v9�Z26��Ƹa�b����}���Fu�lŎ������5�m�7f����v}H.���]�����M��DkF7@v�Q�l��]M�Y]�8U�x+�aj�Ak�[`u���mnή..�샃��R�8�j�e�y�6�Em���[��c���x�w��1���0�ј���r�'��>���_Wge��8H�lI�$��{<dc;�x�z��ˮYk�8$+&���<\�DL��������Lb���_�c:�	2d(�E���@����V:�koy�L�@U��"���=JJy7N=oz����(�/F�`"��(`��웵��k��5^�Ϲ�ӊy[fy}p�hl���Aڼ~h�Ǹ��J�!֩~Z3�=�r5���!.A�YpC�rڕC�������Ի��}��U�u�I� ���������e��\�o�D�lS¤��L�<n\�}�/ڋ��v֎�jΥx��p��[����7>Iv�/�w��c� �5�KeF�㞈���op{*�{���M����G%�+�o)�۾��^�x"�sen�vj�$�8�-�e9!�z�R�@�v+��H0]jy�n��G�ci�nq�x�ȶ�yT��n-�7�D�E�^�C���M˽�O^�yI�����}X���.��O�Y�Zr�
ү'�f�wf�U���;4����{%H�6c���Z�=��љ��B��.�޸Ȋ(�D�E�u��~�T�.��Gw�Dw�(��>��={� ��f�F.cX���6};}[��\�M��'J$Q��5mC�g�`���v�7�ٞ����[uwך�-o^�P��x&�<��\���e����)����
D�ʪl���r#ȋgy*B���i;��ִq�u�7��1���{�0]�;�:�+�^����z2$=�N���t��Q�Z����n�Rn�-�C��0�h�\�I�j?]�%��V'�s����>[f��Ϸ�3Ч{��}��m�yGB�5�v�}�ˁ��p%��׹-����;��0V��Ory=~�O�x�;��#g��~�J�������v/{��q%0�fˌ[�b��x=�ǅ��o�����zp�j�_����ߗl#�Iv�w�z��
��y�1����5�V�;������G"��:��TԂ���>M��##=}'����t�����n�b���׻�^JZ�:L-o�!%�Y�SA6�R��6y���q�C'^��t�m���Ѹ-�Y�9�|{bE��/p`[n����v
~&d�H����p�X@�Rp���5��˨�v�	"�-���R�􈹤�O��v{9��~̓$�=櫮��C���I�r�8Z�
�ݖ����)�,�bgQl��s��@��g^Z����䓋�x�����0삪I��z��C�gvd�X�zU�X�^2o��y)hs�M�*�uYY%���R��0�̎8/��Ԋ�����o�������4傩6>����/��0j�����n��k[�{�e��B�	����vt�֪x�bddL����b?Z�E��+���{�]F�ޡ+�FW����"F6�.8��/�.�w������p9i��c�#5I�p<����Et9��P0�{���X��=�ebL��t�*��L\oe�F!j�\}��rn������{�&�e����Ə;z�t�=:�מ��C��)Q��7"��Hw}垃�%���yT��ׂ��a	�{b��M�,��=�������n�т��>�.�������#��Sqz���9wUuŭ�ű���fEK-�۷k,[���d4Q�׹'�����y���{gF{��z�(�vד��.�<�5�b9*���{��Y9w�}��#䁅8�F୍׶y����R�1�8�������Yp6j�o�"{��=!m�4��#^�T�襁����۱��@Dl��N[���,vg�T�{Ʋ�ZL]x)i��׳�6�)�)���3F���o}��-���Rq��p�]D[����<���4W�nƌL��u�t�ۭ�����lN_Y�����>�nM�^�G}���+�ePE#i@�RH٥A�^H=�$�ʈ�{��yh��gm{����3X�Tl����+��C�c�W
�w}�4W����]��Y����,Յ���Nn���/fp��ʞ:{�ܠ�_��\�����n���cBn[�۬��Wa��f���${��!<�n����K��{�Xξ�r�n�.�:zOMG�}I8
6�O���eton����BI��}����"W��m��7�����W�^J>�h^��N��ܳ�g�S�H���}kuu�w�Q+5�:8�
x�oe�H���@o��]�g�� S�����W��&�x����ŷITya�Z�����9����M!ٷxSp�|o.�M������a����*��_�g���I��S��d��Z�3~�g��w�BC���묑$�)�����57wsK�y�s�0ee�DՈs����rv ����xz�ȗR2Y���5�<�j%�s��ީ���ИT����A:z\(Zp�������z'ӑ{Fr�m�aG�L`���<p�~n3��S��zqH�n�JK�u·&��qAY����R���s�j�V�]*H�[�!7�Z�R�l&d�E�T�JGq}��8�"R�p7�<�9�����ط]���Y��k���Y��:2ZfWlQ��i�YW+�

�bI��u�S�r!���nk���d�s�·�c�u*h����[̭�<\����f��9֕��Js��u�I=�R��e�ԏ��=9��-�2��P�[�$J�y�軭�*�|���ނ]aQܴ戮�s�v!A�f_Z�!�����=E���d���8��Y6Dc4�n�Q��[i���V�v�7���g�F��n{xRn�q���84]�X�����-��d�v�r��{T��n8��%b�p'n��ܫ��y�^I�Ξ�6n���;Vۍ��U��#	1�m�g�6۔7�nu�Z�����:Zv�u��<=�z��E�/{'�����ۚy�e�P�u��q�9C:*z���EJ�Z(��L��F�I�&2+۞��W�zŭ��n�q�1^N{�T�3���G�\7`��!un���q��Q�=3��Q��p���]�\ݮzi�[/����[���޺��yo7<�7�.�gu*����n��3����kJ�cX�U�W�l�TL��bDMZ�Ҁ�^�C����i�S6z�-�;lt�{�m�Ʈ��Y���N�^϶�H����A55n�6���l�ɽ\�8����P��]�ںYYw1۸)�{�z+{K<彰���.�k�ю��7�!ss��){h:���v�����k�=sӨm�ۄ�s�jw<���Umz���Rd�\`W�*Gѧ��r&�޸�x<�ZF���Kwms�M��׎��or�
(SH m�Ehe�-�#\g+m۴�#�:Q�L�]=�9팜��ǵ�v��@0t�t�[]�X}��W=��mv�scv*���^9��ۍ�`$�m�X��r��������;���{\��D�.,�^����ͷI���v��Һ��i��-�w[u(۞|��v6ɤUʶ�gmZ���űx��� ��c�v+��zSe��]�.y���^Z7y�@S����秄ۨU���9�[k`ƭGl�	�B6��B&���uz��s�e�}�;���:�9�}���A��m�^�.�Q�,q�K�6ױw;�h���<���w���9K�M��nLGVb\'g��ݣN}��Y_/���p����˺cz���c>v�W�k���\��)vh�P��%%ۉ�;m	�:�:�����3�ٸ�.*e-�a�c��;��:��9�Lu�j��j6����G�哶��,��s�x8�������1�6��m1�'�6:��t��ع��F���ޯm�ӛn��N[��1u�Z���;�F�O^b}�}n-�s���xz`��oX�N���p[n������,k��k�����5����A�;�mc�s�t��x�Mv�q\k�s���Iq0^m�+��9�,�b�7�חCp����Klc&��v��/�^��\�u�sʞ:W8�ND�@#pH�d��g/���	^ąc4~]=���r�+�kg�i��(G��>����g�X2�����	�.H��G���f��b����M������u��� ���@�~��B�_����R�Ǐ��a�Ƶ�ۯ���r������<��ǑmQ�)�m|Gj,��R�Y+��'�U5^�vÕ���-�)�h�A�S9p�}�DN�0�L�;��TN��B>���r��S�	h�N����]�j6�.��,x��W����|~�����[^���P��Jv����?A|4�@f꥛F3l����V�f\'��;F�@���N�s��;]�m�%S-�1�d[O.;ؒ����
x�3��[_L|�8����!P�j��T�f����#�?|vU�����f��SD0�,�V���Ts��^ϻ�h�A�̶�h��d}�LδC�}!mK-�����酯K�k�Uꂔ����d������G]���f :�ev�]����6�LK�g�dɑ�.�p䤈BhձE[WU6�����?���{3�8Ի�
h�=�k�k9�Tï�l�;p��9�xZ#��%����kF_�i`����9�UV{�\.3�=rx�o�|��W�Ѭ��u��h����q���i�ÎA_6D��1g�e3�>�a���_��8�D��G��.��o|=� T�쓷�qv��{b��Lڟ��)L�t��ko�lX���k��9C����QI���x[���鳤�:ˍ畴9�C&�Vw��hﷳH���協탯s���D���k�����,؅�!繿OZ�}󩇾�MSX�h�y�}U�5TvA;Kjޗ�Q�}M(��ｔZ1�:h���z��|��N2��
?R�*��C�w~�f�;F�׮��[�o2y�-�{���'�Њta���4�:�a͌�ˀ��08$�_�Oؐ�|U��x�dߨ���9���3��ݴSD3�
�����z�n��G��F=as8�S5�_y��v�q��=��w��gY��cV���+�X�����O�-,��
�%�Ǭ�D��]����¯<���d#���l�_�ϧ���}����~�3��QM}��OXU߾�:ɷsơ������M�}����=|j����-��*�L�A���16C<�A�'ѧ�-��½�;'I�ڑ�k[s]����n�eܗ]4��P���%=���J=(�ZW���_6��y��e��E��>���fs���~f2�K��y��g��o�9��D�ߺ���-�S�cG39�gZ֥��]�^�K���I>b�PwV��V��ֲZ%���Vy�|��y�Ϧ95�l�U>)j��eʎJ����b5�3�ST�~�$/���h�D:�	���0�/<��B�Eozf=.����:��d�io�i��F�d�%��zR���-��Fn{&ѯ�x�[>�.g%�~��� ������ݯ~|nߺ;�K"ӆe��S[�s �=A���vw{����`��ܞ�v5C�ᗔ_;����D�IﲌA�/7ۦ�"E���:��4� u�?�ދ.yu���7�c-ö�h��=�@Ԋ���e�oK�4�F�g1���;�{���C���~���fw%[���f5^��ӈ���Y׍{�kX��yy�E��e3��XU�>�s�qL��>���޾�Y�7��ʅ�����C��$�"H����ax�~�(ޠ(���}μG��w��d�}��Evx�{��G��ۧoY̓Y�����a�B.aÜ���s��,-��K5�"�t�Ǐ�Q�k�S���?ߧ�*nh�@�<7Z��nwo/\&;O�Iwm�vt�UX�Qɜ��-�v�=u�(R����;�{���D3.}��Xc�w�+kYm�j�شTNR%�f�1�U�!��,6j��0��}=��,��[u��vM}+:im�ҏJ1�w�����8����m(�Ǧ��!�	V�燳��k7�/���{�_ow%S-�=[�h��E4C>j_~��/���`�!��"�M_��,����oϼ+��&�y�SX�:���u}�6GtPv�m~c^z��S)����Gӟr-��7JZ�<������7�ʹ!�A5�~4�~�����s�yvo�??�d~���A����(��!mp<�W"ֳ_X{;��5�>��z�_����hKam���vk�0�g�|����ڪ�F=J�N��u�x���%����F4C]ْ�!�c���N_-7�D5�ĵ���=8}~y�&��V����lJ��sO��)o.��/��t�'z�Z'^m�q5����*js/��p�ڄ���Y������hƏm9�2c6�a��-���	�-���Z��ׯ�> 止Y��~���G�>t�˄K9Rχ�T�q{~����J!�3��Y���"�|����7)�5�o�/����������V�̦��k���ӟa3n�ˊ�n��5��0�V� ��dH�`�8�VUXE(ԯ����.a�
as-߿N���%������F3�P�M��r���g�h�9(����mu��k����v�ӿe�޾^��x�_�SF^}��>�0��t�C���$&IO�"QRT���U:��h�|��n�m�#�O9�b8�S�̝����5�^uK㶸l/��Ư����[�]e5�S޸���W>�K�!Cl<�>Ͼ�j̈́qE��C���l���D��~%z"YK_A0T�UF#Z��'�A�Q;;�l4{��)�5�jZ=�Wk�]2Z�s���h��o�{�R���q��ߢ�����
x�,72m�Ӝ�Y�kDmH���B)�,C=��@Z,c0��X������Qy���ӞMu1�"��!����(c�:ϙN.5����d��R���Xu�]e5�u��c=���н��Q�'j���.��a������E�j� �a����R��o�d0�Q��
8/u�Z�K���<�nk��l<��e4Gq��ֳY�yGܮ�>8�7�v�͔[�c;p�������rl;��v������6��uٽ�ƎM�c�!}P[�f:�ߥ���nmX��� ��͐��.���'{���15��%�}Z!�e�Z.,��\ǰ�^��o�K�.�*��L~��F1��e'�:w`ݫ�Z".W!��n�՗r����7�e�p<g`�������{m����x�⤮��7�F�dӴ6n�;���j�!�>��D7;q���^vwVS�b�u��[��}Ӟ^wN��E��9On)�lv��<n����	ӹ5���Վlr)y늵�nx�m�&�v�������y�k9͌lq���v�ۛ[���q��t.G���fd�ۄ��ޗ��jg
p���kR;��.t��h�%��-����vW�����[�}kOA7��`�e�X�g��\���dJʝ���*甋h�L�:��W��,'���{38v�s�יO뀶�߹���Ǜ�h�y���-��-� ��i���?hjV�D�W�[z�*�E��ĸ�@�������8fkĽ5�ɚ5S�k�r��L�y�K:ִK��.�s�g��>4S���\woӬ|�<�}�h�q�Ͻ��s��S�SDq`�8;jq�[l���I���Q�{a,'~��{�k����1�5����n?ߕ|;y�!�nvT���O%N]]t���>0�_{>4K��n٬׮�{����\�������ŵ,�SY���?6����a�dp_�O��?x���lل��y������|�Z���ܔ[�G/�k�ѕ�W��h���RGb� j��8�����3?~��_�e�݋F3��� ����8a�;���
d�1�aH�|7U��гd6@�����Z1���KD3�̕�Q}�_}^�&o=��C�25ķl���%��z���S��T���֛���6C\�.dؗ�cV}c�+�ܯA�b�Ș�lo�Z���;�Z핺'�d�v;pv� Z���i��ݳ�8x�5�K���is	5��Q�q�>��@[	}���h�CM�f8ϙl���]��شgb�SYSD>?<a����'.,�{S��<F��_��2�ؿ�,�Z�˖�մUB;�ψ�
)AR)e{^z��5^�iW[]����a�~'��;��iz�d�Z��FW���P��W�R���dNN��5����^툻14Cd^ȳX�}�j:7̌L\����.U��(:���ng�P�ֈef��r�7�7y(���î�d�����^��B)���9�ε�u��\}S]�{Íu���hٽ�|�GRX�5,�4��O��.���xu���oZ!�!��\��ih�[R��U��ESgzu����mf{|�|�����rrg�B9���f���.�W��~�oJg�sR�K��^Kk�)�.�o��=8��=�~~0�y��h���C�1�f���ܷh��L[E1��\ŴO�o܌�%����\=����@��<�nw���-k�v�G�����;����4�t�=:�>4�%�E4CV����P�3�
��3 <���}��rz$|_G;�q��,���;uٰ�D4K�����Z#�_]�����-fF;jq>�{�{�9�o"t���&�l��3sڦ��c%ǘ�=e9������W��)��V�-���尕�iy�u��~u��|~���8ןY�p�����=pu�|�}ɾ�δQ���hBȆ� k��ƀ1��׋���G;O�S�����d���:�C�ץ�k`��q�X ����-�v!
 Cڀ���K��_�H���#�g7�5�T�ˋaL�!vw:�L��%�cu~���s���֩��÷���}P�4ol�3�g3Q\���KU~���ߢ�`�*���K�Hz���QmC%�q���-h����-d��w��g�!��NPk�o��;�Ϟ�=�LP���>��AB��uoE�}�cȫ2�hP�P�0t�M��S����M��o|���'K���֘��7F��n!�G����^�A�D��C�)��ﾛ.!c���KD>�vO>��[:7hU$���N�q���="����j�9������WȌ!ֿ�z�H�h����4�D�f��F�#Z;;��g�ن�m�5��������[��F�}�g��p�j=u��4�˛����K.d���k��E��0�-Wnc����j��Ї���,ٕ�ޒ��?oߦf��k��r�Y�Mre�1��v,&#XO��N�c:�v��۹d��ڔ}k���<~�#�Z��ߑ�+�fv��Ѹ�c� u.&{5R=Q��x��|�s���;n��^�Ǐ�붦h:iY�ߞ����5�M�ì����}����Ƹ��"�!�ϭF^}�ɮJ-�d���μ����XL�y��n~����)��Km��,�����˶kǭ}Y�!�͟s4�[�YX�[N$>5��!c��J�_��r0���M�~ߢ����eCk�ۃ>�R36Q�>5��aa��{d5�d��4eV��׌֊��=����IX;�mw������·a�	��p%"����~KmDS���4�	��8G�q�0��Z� �D�2�u~������5�r��a�F�r��S^|v�;����E�2|������~�}���^��8K�N8��ߺ�~�b?�Ww.#&�h�NT��>��aK-��k��,>s�Hu�U�{f�k��)����q�{�`Q�~���ۿ�O~;W�2��gz�u�T�J��2֮g���5�Q}YZi����E���05X��o%�|�N�lʱ���::�f�η��|�B�����>g��r/q��-X�j�=;�BKL�7Nj"h��ƭ��U�_a�ɴk�ږ@�p�t�|oO��;Ogӹ�h�D?���-��;꿢��k��W���k5������g�
?��w�Rm[$���`>{��W����sE��c�"9عW�2t5�	q�q�7m�h�����h�����ߗ=��|k�����ۋ�2=R�8�\"�{/�E�8>��HKͅ�A���-N��XL��nO�yߢm�|�Ć0�Ƶ��s�g�8ԕ�f33�m�5��ڏ�N��T���\|ko�~���G߲Q���6�?%η�YFr�q�C�����h��2&'��kn����X��֐�*�S��O~UFj��L��S��4u�_���V��+.����őWJR�[-{����ⶋ~�>e����sK��.�P�{�g~�ƾ�Ađe��'�k9��ڭ�Kf�.�'Zs�u�C�R��<凞�՚a���4z͔S1��í�=���P���I���3�x��~޻���]G����B�݈��]�B���������:ɔS8�ۋ�[���U�?ھ�Eh�nZ����X�DC:�}܋6�N:g�nl��1� ���_��Z���m{K��q��q�c���[G����3d¦������ѝ���7�e��-c.�(��=��[G>��1��e���Ǝ������c5�<>��3Y��A/����*f~K�����;{�埝1�[i��837�3�,lW�ֳ��������:�|v��{���m��L.lpu��{���6�/��=�I��艻s�u��u���ى�{qsWcl�۟<<X�5�Z�tpo&��u���?������M]7j�=��="��l��Ub��7+q`�D�>|v㱃.����W�\�pvH�[��.@���N��k���q��(x
C����������6����۹��۬�f��ko%e���؋�p۷�5��lv�4�X�N�KR!�.��U5�p��Z.X��l!�������wHKc��1v+��
wj���{1e"����������4S���L91����xÌ���j�$f���g��eq����S�}!��}�׾#���n����v�5��5�w�,��ֲ�Ɇ�e�dDGt����c�����K�_&�K��5vm��o?���a�)z���nz���Đyq����s��<E��-ԲZ�)�<��9Ȱ���0�����羲ɨ-�GdU�+�)b�a<���Q���{��KeG�7X�J��5箵^�Tƕ|zo۟}S}m���O�9��Z�g��lwm�7HD�7y�����Mt��ϰ��F�v�}l8�}����6jYȪD=���E�s�8�Dh����[f���Ao[u|����s�"N�Y�:��{qh�]I�N���[]�s�k����[_<v�j���9�vQ�-���:���_�Ə_8���u��ln/�#�ҏFz[�����"X��m6��e:aO-�*�0��{�v�h�r���*v>���{���;�D�O�@&��P���(Yh��Q־����2�O���t�jnܖ���jn/�����CH�m85\lN5g��s�j�*��f�������;�\�A�l�`�|/��@�H��_~�!���d�.�2�QM}�;G��(���`E������߈��kpǽ��g�t�f>�5�/��el-0������]"�__k���`J3	��|4�.�$�[�K�������/�5�~���������AWk�w�nt[�v�滗��hv3��5Y��ƺ9���G�-�L����|t7��n=N$��s¯���.��y�VB�e�Z;|�S\U��c�w�0<>4KD0��َ�?����O�>~�:u��<�#�6�K�pGP�$q_�5}ޙ��e:e0��o݋F�&�hȢ��^2�3�#�����:a�����K�:�Ӈ|���Q|�ͮ?kY�0t�}qp��Ϲ�FִD9��Z{D��F��[?~U
�-��;-[��K(�P�Ĳ���1M���b��(
:GO�2�\q�{����3Ƹ��oXK-�xþ϶,�ƎTd�����w�fs�y��ƎmJ�-�e5L��pn�.
&���Q4Z5��Im��ڄg�f��fq�T��1�%�d��{9��n��=�.]v��\~h��PSE?t��f���|��p�8p��������c:ǥh�u�~(�ı��}����d؀�g���8�jJ27�:�+�q6�� �|n7mEh۝ ܵv�m�;#n�����Z�q08q3O���\O�m[-�r��_eֳ͚�
��x�e����p�?_)��f��ߣ�mr�7X��w�l���>5���c��rϯ/�gZ�EEJ!�.�~���jZ4!�c��4��[��Ag��h��4@Zwa��T=�mr�}��WY�[��2���=ߦ���%����x��T������D�CFLCm������lQ�?��?��yl�;���z���{�+��)"�2\����C��A�k׭՛ɰ��3�n�4i0�h���v��ݤ[M:�:G;=�tk����`W����l�%h[(ؓ�P��1�b,��=���ZS�T�$y�"4��d{ᥦ7ϰr�.iSj�(�'V��3,S���V��z���ͣ�W�K��W!��k	�������Q�Y�j�]9��D���g.�j���]�VW5�n�.̦�WgQU)lͶѨ:6xMk��qVNHzd>��q��=���c>�Z��s�SR��0�7˄Ƚh��úW�2��;td3��o�=H��\d�Ym��7oRk��9�2��ݝ9[�&�U�W]�vX߱�.�A��6���`��\NI����%�Sշs�u:7���CG�N����=.ץ��R+V��z����7ԅRL�;�ٲ�E�J��kr��}�7��Fp,�ν�J�Z�U�L�q�<7Uz�}�ud�&�!G:�P[n�����H�T�;��7�,��f��'++t����L�ф_5�s��E��w:���\s�co�-����ݽ(�x�QIշ��v.-Oe�(<��st��৴���
��8��l{F��";�����<�^ABa�a�
Yl��(�Х�s.�ػft�3r
�@^�ݭM��ڽSm�Wn��N��N���ҟ%#"�Q�Ŷ�S���+=�;�Bw{�5�t��Β�
<�Y��[X�]�Sw�c�g�e��]ka:�X������\�.�MlW �.����n�B<��#�CϡDrH���Pcܗl�0*�vm�������h;�k=s��Vrl=Ƹ�u�ϙ�F�s�s�ϲ��g�M{6$�>V�ƠCV�\�W�c\}u�����=ϫ05��ˇ�y���Mܮd#��R-�l(��شw�e��E�o�����a3�O>��C�~�Ֆr2ߣ���;�E�u=f���)��~�EW��φ�QU)c%�sK�Q����Y�����a��s%c)�>�<f��v��~��_W���,���ޚan��׬֏�^ڠ+<@���D#k9_:�ʁ�8ᢾ�׏Y����n>��-�j�ۆ��r�Ev3j����;i�pܤ^��+�>��`z�g���o�;�a�*�턴w��;F2reSF�/�N����-h����.��w�,*�1�/���e��=�a>�[>k���Y�С�3�d�<3Z��h��}6c�DC�Tq�p����E��G���g��ᡜ�%���J�6�>g�E�v�õ|7y��,9��h��K�@{=�T^3���,��Oh h���9����yȈ=�w��U�Z��0�D��üH�҈���0I15kZ�s!�1��x�9aC��F�Y�M�!M��B��_E�6%�m��w��s�T��5�>|?_�q���*����uϲp�`��E\6ڮ�`*��zg뭈�ji�Z��d��Ƹ�h����FE��8�lrg��ь�Bˀ���)����}�h��QM:�Y֩�޼�,'���D�g���}y�W��P���g�<�+�M�n��}��٫iA��Q��|�w�\�+���d5��&��D���xv�f{�ϣ�j�
V$t朏^l�gᕹZ���o[���<=+Ͻ�� (�:"*�Nj��k�����?{���q�}�X�W�s�f��U.�}��;Gv3�2Y�c�E�w�C2�YƱ��f�j-�׿}����O��z�I�m���]���	�ۊ5b}d�Z�dŜ�z�P�L:��B�۶�m���p L�����3w��Or'r}��~kLF���ш��F�g}��~�_�̨];���)��v�rA��k��p�"v~q1fg������\�ճ��-�{m�6�wvLh߾�⟛�M6Z��ے�a�;󽡄8@�B|�_E�X���A4��+� ��Z)�~dw>�י��SD4C}�!g��a�/�O��5�>��ŝ���G�O޳�S7�w�O�8�~�fxFQF�p�p`�H�E�"�g�> O���<��c�}�],h��%�9�/}7�e�y�T2ڋ�Q�$�����3歟L.�=ȼj{~z�<�k�ހ��06�߾�e}Z��n�S���4����tM6��d�T������g�/-�������͚�{��{/=kZ3aq���/}����u�Z�{�笖7��>�Y~k?Gܾ�ߘ@U��g궟�`?���4�0���G�2cj<[=��L��KeL�U<F�^�-��?l����_>z�>;�T�MǗ��s��u}S],8������L���Xlo�,>�֊|a,�_�q�+��v�hҮO��!SE�O�^�����
���ϡ�7��p�/:(Q�7��y��C9kv��m��UnUVF��X�b>�"���1��L���)9s�f��[ `��`'E�d����6�ˢ���#{�5ڶƻc��%s�ܹz*W��ɍ�x!�c(�$;x��t�9k�y��s�`��f��]�և\��mE�x����Erb[8K���:�q����mɥ��v�1����:{s[�v;'-��l���x�j�u����nYk�K��ۀ�j��ڭ�!Q�Yn� �
�����nN�v���`���&Jt���-Z�R�.��7T.���u���.��kr-G���u�鍟dca���уם�m�m"�?6��N-gb
j��SD�Spu����ßO�r��Ù9-u�h��:�"��ck>ܺE�<=%�Uyc��+teBe7�ǭ�*�	V���}��g|diono�O|ƻ���h��(u�߉1�6��E��Z��r�@`���Oμp�	+"�U��ޗ�+��x��.�d~=?V"i ��>��qS4j5�gb-0��~��2��F4[G��ߡn}\�5�5�N������UW�-��Ɗh�V�Z1��"B�r��"~�[X���%5mg�F����Ф����⌔�Y����o1��f�����<�ę�oC�����W�+=vn޿5�CSݬ����t�e4K�䇾��Z8�%������E�UB��޻)�4K��/Z�������J0ƣ&(�2GtF�=����mcV�k�G�s�]�C�V������+]M���s��x^����|1�}4S��w���Z��J;�;=��C�h�}�M������-�d��>�wf2aܿ���p��	S�e�=���rU��n`bz�z��ly�����$a�I�9v�P���޿5��N�`���k�>����af[
}�J-�>�&��N��?hi����^��`e�sy���;&�l<���}A�������ز�5����f��5�=vb��O+��Y*t��F#�Aۂ�o������h�W|R4j�˃._�|�B���d��5�W�ſg�M9y<;��p���R�`�H�c�b��Wo]��v�(V�بZ,41Wei�����?I� |���E�d�	��a[%��{쿣��KG=���b���C̽���އ��</O��p�f�di�����6mF�eT$���b5�d�K� )���~���O�㶌+$���a'>�-K+��E���on�ξ�k�u�c槼�|��6�SG&��_�E�ϛ���7a^��Z�m~[�|m��Dm��5�kY���`��n�ʂ>�{늞�Ǜ����B��j�,�����ָ�N��\"mz���ގ�Sۙ
e�8�oV���ߟ���{���h�ծ����D?��ƈ���A@Y�Ł����5^��i6�����Y����3�:+h��)�e�׹%�ޚ��e\�u�t���g�9k��ذ�c����Tof�>�}���ʆ�ܺE��pSX2�o�~��y���Kf���`F��"UP�\�y^�Mn0=s��^�2!�9�=z�(�%� �
m��>�a�3��#����Ʊ���U��q��Q�}P����k܄S�a�<aZ"����Mfr˯E>CF4CGf�~�/������.���Ҟw�A��ѹkN�\gmS�zβڶ?������F˿Uϧ"uKD�2�l��io>�۴u��3�0�oO�}z`}������W���a�g�#����p�	��������\z�װ�38��֥��QR�I��ֈh�cR�Ͼ��_�5�Z>�������۴c�7CN/�g��qVg����3N���F��4,������4�42�{Ӝ�Wk�1_٣��U�vٚsVts�I���
��a�̯���_��6�gZ)���%�������M�֏�-6CG~��jb�U�ڄ[M�q��"��Hپ��z�KxK8�n{�S�c;���Ͼ�8�Y�d÷d���$�,�Q��?t�b�����ƈ0���4}�\���������w�_ӈ�G���^5m]�q��m?ߛ�ҒY[�QR�4����K��s�P٬�F����6�g�2�ư�d
4|�܌q��]�
�{}����q�	|羞g��q��5L�|���#�B%�2Z�`���)�����?�~��c�3��`FͥŦzx6oXc�wkpX���08�{[�ݹ��jUF��[k�zpҏ�U����vgq�d�ck�D3ޅ�[�Fg%[-�����a��~v��w'����s{�4{ <��;r��z,�p���Am�^pS/����JQZ�[[Lך�W0MB!�-�ϙ��r~�G~����ݳrܕQ��y6�z-U��f�F�C\ݒ��1��T����f3�q�7��r�Pᢲ��Y-cCי��[Du�ߵ��_�b-�qB[)�.���J��!� ����
7���@��"�~i��݋C�D5QU���uіt��sÓ�~��1��!��d���t�в>�Ջ�5箵�K�U�������@?Ie��t-[U�O>�����߼��w�ObѬ����j�Y�N;��&�%�󂚟Al��^ϝ�Z�l@����e뢑.��<Ϳ|BY�m�����U�/a3k9�B'f�+�l�^5	e��坓L��z��ج!��>�Kh�6�Ԝ�Z����֏d"��k-���r�9�eC���Yfim��Ϣ�[j�ՎD��_���;u�q~�?E�@��������~�L�E0mq�P�)�@ssދ�ބ]ƌ)�Z>��ݜF�aU�F��B���?N_��R��EA��țy���ma���٬�;kA���r��7�`��6>�x��-�����6���ÿ��<��c��)���{�ɴk99���
��[G��m|�k����e��h��>��s�1/�3i��YMy���泿n���_q~�,�F�(�:_�=����Z3L�sK�q��(��{�������G7�溧B�����g��d���gخ�_͵�oJ]f�l�S�W2~�F��AN@{  v�s违��#,�7�=���wa�9���D�%N��l�/��N��u�x�������^��kl��t���!q�����M�Z!�>�y��u��h�le㵮޴S�MS�����F�\hq1���ggb�X���˿���ږ�m��Yֽ��-�N����^�k��d�1���B��μe|����cRr
ko���n}��L����aI��$O�����~�G}[�NkY�۷H����C��%�w��"H��Qq�%n0�U�;��j�-������"�*aQn8�/w���/�k"�d���|�k����t�����ذ׭���KCο~t�5����",�t��a����?G��/8�|�8�py��'F�8����y��;��t��weȧ�.
{���n��*��k��1^�B��;����sf{Ʊ�br4LBq��� vi큸��8x:�v��]h�oQV�����u��/V��s���vm��q��z�n.r�u�B�p��$��l9��vyϵ6��N���=����.x�B�m��l7E�܆q��j�� �۸뗳��H�}��]/�� �݌�sz�`�N���-��ٳY�#��8D����wt�'`θJC!yv�a!1�ڄ*��M!�P�]p�F�)�E�����s��;7l9����nG'l��]�Pn5uV�v�n��Le6[����۩��Ƹ
ae{�k9{�h}������3���Z'�H�ؚ��/��k׿���C77�~C���S�z���D�@�g��7{��Yϡu���K\e4s|�0 ��&��Ur۽.=y��4���BY��u�oܩ�q�X��c�G�~��}��-۫�3�[�h�D5�KC�%�<��Vy�^����m���fd(e���,�������*`���)T�fb[��޴KD?��}���a�q�Y-z�y��4��ɵ,Ɖk>��9���k�|p��f�C��-���pq�/���\�1���;�aM?AM	���.�Lăf�)����q���տ�Fd��}'B7��ͣ.=8a��%4����6��	�t���ݰ�����MG�}����m����uW7�F�{�t�czיn�]�@����~?����n}!JC�����Kx�E���,h���;Z:z��+�F����~/�mGW��s��SS��ߞ4�a��2l)�>ct�5�k��,'�}���h�MR!�DC���{�rbo����wб������.'���;����M�/gwN��h�&�{4�+5��MOQ�����uߤ1��ϲ-��l��Ql�������U���ոf_����`�����nnO~�~̙q{r�?��k�n7��ц};�d�	k]k�����	#*��f������aL>ȯe�>1���O}�V;��V�;�g*wR�Zv�0��n]��C��7r<ꆂf���W��a��8��DA�<
����y6�kK�<�����\"�]�D��}Q�\]r�C?g��iäʇ��hY���s^:�d3��E9�٭d��yW���ر�o�oO',��KX�ٚy
����-S
~��l��`���̹G.!�7�^�{�h�a�u��^g�\�*��}-�3�Xm��M��g��2�Mw�o�9�~���h��Q˅w�����<��l��d����浪��Q�㳧OVn~O0.\Q�(�_��0���Ǟ�ry(�w��l�>�͘�}�պgYm��!�����=�Ϛ-�	cff�-�S���>k���b8�5�A�Up��$Ɨ>����=
��^im�4�㼀�[=�}ʯ��ǎ���f�#����}�#�k1�^��e��!�?��ǘk����n�����5�2�m[r3>��ѭ�]N�l���|o���n��d��N�v���2�V�e���:㮸�ФKnN�;�Q�9ӱ���(��S*|X-���?�AG�� T_Q���}WNѬʅM־:e5������'�f5�"���l<�s��A�u��k�"���n2�X�g*v�i�"=�v��h�;����5RC�:qO�mc��O}H�A��|�q�ϝ����F\/���Qx�T�;�0�D�ݩE<a�������֊{�
k8�Dg�~�F�g�bI�s�p��TεL��c���ŗU����/�U�z�Q�6:��s�h�)�h�M�l�/�}]ͯ�q}�C����
��UO߲w�8���@!�*q�/R-��4�6���^~�XV�[��hS6�0Ģ�S�;8Vmv�31�W����a�Y�@.��@s�ƭ������ ��%��6��_и����CY�cE|��
l��SQ"rE_?v��ĞJ�_����ܑ��C�e��}��;�T��}����[XZ�M��#��)�q��9��aag#������r�fTO\�4N��E��_�*�Qn�KE��y�?�aQ
P-7���5��>Tޖ?�(Ҹ��ag��mBm��E������)ߧ6��/��}��Œְ�M�����赎^�ao�c-��h�}{�a��.�S<�dKA�77������:lʾE6��.�q�K�ȓ�ݨ����ώ���Y�:6w8���g�;Oo�1�qۦ����Ovan_�S���4�k<Gg����D������v�وm�vKh��^��|j����q��~}Đ?~@"�a���y����=��<d?�M��;�ڨu��)g��¯�zU�J4�|����5�\�V��_y�r/�{�-�nlچ{6W�ƫ���!�>��ϝ��=h�S\�;s��=W�9����}xvc��>k�_H-�=�C؈���u�9"bjuz�n�YƎ?�K��}��b5���Xяޅn��,�����gt�!������ѿ�<@�ø����Yp��Z)�	k���~~p������\z[��4��n������� ��K"e��5S���5g�&4fF�3��|�#4<ïy7ȵ�F��h�B%��O.>�mε-�D�a��>���ɝk�C}�}p�'ݻMy��^�u�p!����U2�NXs;��E�Yǩ�k�ޞl���/���re돎V�l�u]��8�ƕ�g�,��a��h��g��k׵���n�5�t�z�l-d}����ƫ�����KϽ5Ʊ�G>ˈj��}�M��15-�ߞ״�m�ٛ�mn}=�c�r��=��c�4C��!����֧��~xpi�;�Cb���,�ګ0N�]�7�m��6�tgI@^.��ݞ.ں��%ٷ���c[qZy�/홠���nu?�ӻ�{��-�h���8-�f�����S]e�z�>��^���k�{Ɇ��]��xռp��֜���g��>�sϚ<�0��vv' !���f���K~h��0���[������n�$@�nCx�#��������~����eؿ��{s�.�Gљ}�0�C]���a��![9����;k�������_��kƩ��d[���ˉ��i{��)t<�t���ߗ"�H|��p�p��cr�$�z�P̨:�-�v����8��:��гa"��c@ҳ�~4n�W
�^/�j��M�>�eg}��3���}�v>�K����gN^�}h��|����%�j/Y�o6km~��!�S`�KD�4�~�C?B!�߈�r��^������Α��֩��Ss>��7賍w�(e5�SD�T��ذoZ!�՛a,(��O����g{�K>}�7�k��<�[D=/��O�$�:�Y%�5��:���m�Ym��FF�ɶ�[��ȆcE��A,³�<�s��/�;���v��K����[o��[h���ܾ�������h��G����Pv|�����fE���lD3)5_x�k&�4fU�#s$	�D���K|(��2nu]����
�c�3}����z�=�{�k�8�L5`��6Њ��V���J�1��K���r:mv;�j	�{#f�=҇fJN��-���<���oI8�Z?���#dL/ɽ=�N��ݮ�Oj��wyu7$%\,�������鳎`�p��ۦ�1]�ɦ�q-��|2���%��]	W�d,��C��e+�)?�h)�=��]��h힎���х+��Y�I�=��v�:�r/
�Y��ɚ*���jȓ(�a���[�-���[}+^t��[��2�P�nQEڟ��7p.�����K#}�~�fgl�ɽ����f�G}��м�r8���g��"o�7l�wm������zo3)k��ԃ<=%��k�/e��:vX�9m:���&-��.VA"�]/e˓�3?O�r; ɉ�;�=�O�ޭp&��v:��eQ��
J�em�(��#�d�S�U29�޾V���>�b��nq�Җ���Yr'��#�S���WR�2���������K��DtE�4Z*��I�)g���N�Z}�c���:�I�y�Z~��۝��)Ƌ�ϭ�=�WP�����6��jvN�'��NI���C7�D���i��/��������>@7�[ݗY���0�g�^�H�'n�E���������N�傺��c�{'K�K��6���X�)J7�(��cj)��G7�<�ww�KM�69IKKjsu`1�=��'m]9w]��a����	�
+���68<0j�Ui��#�! �c�@8���d���Fe�������)�n�:�v���}�_)��T}d�`Ѭs=�'3��G�ܢ��c8���l�=C�����ns������s�9���2�Wn%�(;vom�w2ӻR��N6������89:�����oC�C��Ӻ|<%]�^�7g����fT�nۈ.K]��<�v���H��B0���z��n�^Dgl=�]c�MP��u��g�m�g��;=W���R�]��*�s�@o���u�muWM��<��D��i��WmƷn�]lqt�6����=�;eq�F77�n�[��`׍�DMn=n�\�u�9\����ݶz��]�l{ݸsk(N�/y��ѻ6W�t���>�ۧ�x��R�.g
��X��Շ�8B�l����컎���#���9km��v�pqNͮht>���X<�'*�z܌�f���m� ��!7�7Z�(E�s�fw\轱�Khj[����F�s۳�B��N�a�[n{v�>u|�a�g'�c�(����`��a�l�{`·Q�q��Ls�uˍ��F�F������=ϸ���iúޒ�8�x7���g>z؉��nɰ�ȯc����^��=np�s'8b�9�j⻂s�U�a,�5[t�㫆���.�t؊��k���m�f^�{gp��S��ϣq�A�j�gU�
�G4{u�P�Yڤ�n;Ҝ[4�R�"$�tysQ�d�,ˉ�S�z$�sK�yw ��ڎk�v}�x7v�s�{6����e�C��L�n&I�-y��rT��n��5	�%���q�4�kr����ٴp
議��piګ�ŵ��b�rj�t�S���\�۠6��w;�n�v��N���7={wW"��Ӥ����7�<�垳���s�k4D�W㛒�J\�v���:�ی���S�k<��t[k���2ǱxԼ�n\k78�����
.cnD�N�%�D�8���(��;�^�X{�f�%x�m�#�n�N����8��ܺ;L�;	��nݗq���=[��B�9c��ܮ�s��8z�I�����N���kS�v_}s�6��]]�L�����k����#8����?��7z�v����.�c���qr�]���٫(����8
�v7��*�;�8Ťܼh����b�ͳ껝֫�s0�t�8��"i�g�����=�u�ػcv{�^�"���(��)�!!l��ǯ�8)�e�0��{���a�q�r�j�E��>�w��0�[�\�ьmO���8O�Nfz�_C��CF4CD4v���쁄~!�������4~����$�Y]VP-��=�����J��K0CU���}�γ۵��g2��5c=�E3�Ǐ�߮mK9���K1���%�r��Z���jYO}�z��,�{Њ�~�^����}x��Ǧs�=��a9>2�/|1~���Q������	M;ئ��V���hׯ{
�#ӯl8��A��W�_YfV��~�/_���Õq��D����>������a�{��{�y��j}{W�.�9.�Jު��5ָ����J�_?����r,��V�����?O�Ԗ�_���$w���݊#%m�s²��Os̡��%^��L�C�$�:���:�;��k��9����Ah�3���sYIv��j�m�$��߁��s���������$\��Ԕ��0(:�@d�kŝ��m�E�� +3���-����]�
��qW��t�����z���z߯����:���ښT�I���z�*ЛLb7�����!"��0���<v��ݭθ��o�T��~T��m��?&��ĺ1i͞���՟t�m���C"��Y��dw���� ����za/���^"-;{�2p�s���Ɩ�uR{2�{Ϡǽ,���z&9�Ū��uƷz���"�o��kb?T�u���!LPm4��Β��L���NW,1Z��|}�=�ύ��YU����f��:��b����)W2|`��R�{U��xb�]�he=��kU��v���M���J��r�`�<ݡ����w�V��uK=�F�`�$rHAn��J��Χ����I��W��wK�.:�M�)-{̏޼�l�ݺo�8��zC�e8c%DRl�x��zxiخ���ە�:{��={py�A.�2a��&'Hr@s��3x����v��\�/˺�58O�}�n�J��>W�K\��*h�=�NYg}G�5���)Ǚq8�ng�<pa�usF��ZG�A!�
mY��c�F�1�]�x�k��fT�e�o������6�uf6����'P@q_�PSު���+ٕmN���V�ы���s�=����<U�۾V����1��@���:�3��\�7�����)elR;�@�Ѽy�����+�m�Oi��ܗ��S�U[��
�M���Y����F��^_V�_cl��c�F�A �8\�'&�G5��2�-�̿<7��Q��t�*��K����|��mu�(n��q�٫Gc���_�[�O�e��CO!�P�V��u�_�x��*@z�-�#k&ׄ�6�gi�j9�,�,`��Y�ny}�}x�x�b_ZB���XQ::�J8�����0������6ヘN;�m�7�n����l�}�ͫ�����u+֤�+��s�hZj�]�_�]���rlK�tcQ���V���|ӣ��`_¢l`P��R+����]���1�r�p���-ނ�#��c|���5�UE�ux�I>�|/��W�F�fa�L*�W{�8&�ߛ��,��쏢g9�{<i{�k��qۉ�X�}'|l�>m����Jz��'�~vdb1�>i�6�ލR�k�_���XR�Pd*N�լڄ4�WB�U�����I_��U[�d"b�3�+r!Xg��I�m~�;�z_E�)��=�A׋!�:`g_Zt��%�3�7q,�	Ճ(EiS§�fM���c��5{��K�5[(��qZ���E�q��6OL�C���c�Hڝ����ش[������B�g���Nߵ��R��+�����~~�8kI����+썶c�Q̀�Sn���s���E���	�󐛇�����#<&�>�����a��f�ex�i$�֊����_5~�</��<��n��� �0Gx�D2\�2�
H�[IVJ�W�3Nǘ�e��`/�xw��Df]7΁��:���~W\�ֻ���*��M�������������ILH��(�{�:���x����U�Wc�V����[*�Ǝ/�^�h�1 y��Wއ̼% �1"�n>�.�n�g���DP�^�n?�����S�祻�Y�@�I�
��r�i�}��Ŝ�מ\�ߤ���WǓ���i8��3�=�f�Q�2�z��(/�%d�C�K�E5u����x<�����̗*����Z���K�Aʚ<�Y�/F�M��ڈE5:�
u�V�ˉO�[�ˑU&�\��_i�Mӓ[�L&��Wvm�o��'��Bv�)e�=E�&����8څv閽<⇵�����<���*�9J��=�Ѝ�ɓ�������q�o��63��s��n�^$8���v��
9�n��0��vYtݵ���n��<�]�y��l˂�c��g����+� *	D �n:�(:��l	�Ys���8���6�ש�V���P�z�����vp�&@B6�-`��B�ӷu�H,�`cq�Ǝ�v�˞��t�=qꈨ���kլ"�%?v?��~����7����7|ՋNv����~d��ި&_������g���}��	#M�$'$E�ͅ;��gM���g�92f��25$����������lr̙*a����x�����|	"D�aFI���͝^x0��2\���X����G�?W^X��NN��y�;�e�{�+�����/���t�|a�>�s��oѨ���G�f�k!v&_Q}�Xp'OMX������3��v�>{�2��\Ys��l#$a��a@�Z��c}����a�s��cjOv�]���]�e�����݉�68>k�Y�@<5}�})�<ѿ'l����OWb�O&��X�f���-�)��sX�<=�G��A������.n�=;Pu�q�9;�p���8�FW���0��{�u?[��[�>~:l��O��|����S%�\�z�#���Z�`������^��x���^3�xkdmB��彞���x���V�g	�wP�S(��f-\�9¹m8�[R��)�4f�̿���wN`t.����h3�C:K��[��W_�QȦX�����Ϛ���]�o�|�s��e�tUO��f�aT�%������2��ީ�^t�ׂ��˯Y]k��2���]Xt�b��Ke��S_o��0u�{��,Ǉ���2����X�M%�Z�"�vs����=f�}gꆻ�U�?�q������"_-`+�RO�4eJW}&�yN���g��hX�*�c��]��j8�hD���#K��B/�zU�I��F��5ᇷ��/��G؃�#���/�O�wė�6�@�z���[?/{\�	�7��v�����]''ݥ���>�y�kP�����l;6[��۳)B��n�7-�݉gn�گ���d��I[՞7��h�t��)��A4y�Z�j� �;�kw�U��f��h}dQ�������[,F\
4�Q³^j_!������Ďe{�G(��QZ�A
;�^�"��d(��^
���ǽ��o���WK�a;N��&H��ȬA�C�\��Y�uZ��{��ڒ�����i�lIv%�:�w��R+.]�p������˒����q|__41)��#ZX�z���q���~6I�R�j�d��W�%D�ӹD�4|�xDUuf{ih�b�EG	�b����6a�9$���ܬ�{FrCG����w�%3���n�g�)F��u~�>�=E�m��u��D��6p���/2�=ƈ��|��n����I���a[!�Z���A��A�]�8��-�󱗹�����[�la����C�j��h��<8���cʼF����L���A�Ncqr�=h�56��s�)��3�*듷�ν�'l\����0���8D��� W��]dH�qO|����M�u}�i��/��*e���{/'����cc��n��0��|��߾X8�Q�6EP�L;ץ�)p��7޽��C}�.�f�4�Of���,F��/���c���{�s�2Ͼ$�w����ZCv��퍸I(B�s�ԋ��Dm�]����蟽.խxf9r�W��qow���1���@u����M�̫�N�X�/#����"~p�!6r^^[�^���jDZ�R�;��P?T���i���ϯ��{�?V�%"ń�L2ߐ�p���`�}7(�iZH�1G�`W|r�Wט~���c���唯{�j�Y��ܨr��K/R

��4%�2ϖ߽��}��`ܫn�i6⑆�*H�[�J���WyWe9�>���Jf����{ᗗ�ഌl|,j6o�٤������!�L&缏�6=��/��0�#HL
u^�8�(uĝu��ҕ��ڷl�������\�v�� �"DS"4Q�E�s�������f���e���*ְ�d1}~����Yv���{�]�VT�Eb�<~���{\�
��a@�i��nFo$A���]ٔbȌr��7鱞��*�V�FNb�N�M��6:��/������I��������lr����BDd@�RK���N�:�n���/�ǺyT��г��w��=z�/c>���+}�i'4t��z��=`�!a�?FD-��ww�]�5�
���5�5� k�tϮ�=��������!�W~�����՞��CYo3��o}<����Z͔��{*�y��m_Hl��p����4u%+�&A�=����I��;��B���[��c���)M\�Z�C>���W2j���4�]s������*��G�9X��q�:nl�o����Və��(Vki7A�0f��O��x�j&�W���R@P.�-�n[rs=75���n������Y9N�����֦c��p�xZzW�#�nwGk�Ϸk�%Y�z��͝�F�9a������ӌl��w��&�ۣ�$��nr�;V4[��Ɓܙ7��്z����ۨsei��v���^�p��{>{<�n۫<�;ŲThL���J����c*S���s��n'��6���F��F�j7P����hU0W�{?r�5�:ݻT[��+�i'��]Y&ݵ��w��k�?�^�V�����zکp�
��O��;K���=~{�/Z�t,n���z�^�Jź������%4�i�c�\���|�ƽw��J��n��S�P���Y岸wq�5NN/�{wԍ���Y��Jp՞����Hϯ�_;�*��i��2�)��d0���A�� �p�My�5��g���)ncy3t[��T�CO�o}*L���GX�~�,�ДS�5�g�<Nr��UҲ[+��rARt�=�Ln��{������*(!V*��x�[W����_¸�M�&�gi>���^�{h�>��~0י��D�RH�8D0�ò��J�ʅ��U�a�v%g�Œ\�A��B�^{.�?v��_>N?U|�W��D]��o��C�
�޶�x���g�/#�c7k��1�8��+���%/0sѶ����a�ۖ�r�wm��!�Ux'����f!�o�q�n˲$��QwU�}�w��|n�^��U��x׊ʥ��ڭ>�[q�9�Q��V���1��Q8�}��MYt
�0|����J{�*�;�p�μri�qou�AJNx��RW�MM�C���iwu�!��.	�[�WIIK��d{���3_F,E��2���x�@2�ގ��b	�E����J����+���f=3�/£/��7��#�'��pA�'ڝ��E���N�%�+=G�� �
z��S�>��J���6�垊����q����������l�K���O'm��B%��TѾ��|%ʢ�:' �sK�Q�8��y�8��CE��{6p��r2���-u���_"5[�ؿr-۔K�*hܝ��'���;��ʟmX�9
����q��|MK����ͮ�������m�'�;���G�KUP�tg:A�ȷת�r�`c'7����M����XW��V��b��Ҝ����Z=p��5mKP���g}ݩ��c��	d9�l�L̀_=/]��n�i�J��=���U�g0�ݴ�=k2�wU�#�3��������h�ED*�.n�Ťnǻ�XьY0[���Y�.��[G y��i��֑ٯia������rPy�KJX5���Z��1�5Ma�8(��%P��X�^���f�(���� �|�{��}�;������Է/����h������l��
���%��H]��m]���22�F:h���1gw܋KX��g"�1������L�����t-p��U���p5�
lֳ}��lJk��X�`��|t��{҃v�sb�쎵�,b�[��+k�3p㏱˽�ns}�����w�-=��Y��s\���e>��\z/GE�ݓv�'}Db(��5Ǧ�|E�w}x✥��Ӂ����*��\�;����_.�vc�4�l�Bmf��������ו�f{�I���ˍ��$�8��W{@0x�{Z�f�<[��i͓�A��# ��g����?9��W�<S�t�wh��h]��B{5yЧ��p����H�Ј��׳�Q&y�*{ �y8��/5��/�8S����M�� [����=	;6�7�D�=:y<Kj+g� ŝO��6�L�<�D'[P�9�A����4c6�`����ةL�:�^.�[�q�ʝ����I;̱��b�B����h;b�è����'F�m�!q���On&�9Ԥ����
�܌��3C�dv��h�1ɺ�5�E��ϸO?p�bAoL���tE�ns�6\��9ᓮ�e�ϨnѤ�t�o�R�&Nk��Y̩�(k��М�	�}U2��v=p�Q#�2����c��it��t�ed���P�r(��E���D�Ѹ%�/:[��6t�O�%�1�\c�ކ�w^���AM��ݣ��B�~�Z���Q��4m��BR7��"j�&�%t�[��U�4ќ�&p��g�3���+�ʖ&wIwq�CU��B�ùF�<[!�!�ƆZh�LxHt(؎3�FU�i��f��'��=��S��e���>�3��L� �A�$���v�s[�����!�˽{4�-��W���(sN�e}��?�x�=���E���1���:]f�b���F��޴����!��Q�"{X}d�Юب���?#�#�@�ɽ�\{i;H��{{�`ͨH��a��X�h��Os��Hǝ��b�	`cG���nŝb̂��@�k_��h�_."���hcH�{��G�it�5؄[���ǭ%���c��Ӫ���ޖ�Z�<�M,A�G�3��ik`���%���陃�E�sb��s�*h։hƩ�s!F��V%�K,���cBl^��v����H�"Y-,a.��]>�4���T6ET�3��w�F�a�[nyh�/js�{3]O#���l]�NUaA�YKT"�RZ�����肘u�[5���h������#�&D[���P�\5ф0��mve0X�j����a���؈μ�D>�4Rĭ�gF����m��ȴ\�,`�4���%mp�ץ%w%�l�.eMK p�*��hX�-��b%����KZ��]>MϽ�̚2��IcB-��,V�{wذf�"X�m"�ﴖ�>�y�U.�i��LA��T�;��Ţ�aL�Q���{����c:҉�\�7��zֻ�p]���e��e�bи�mvD[ �kH�ʾ�l֐k�T�q��i%M(�m=~ȰX�>��hF00�����C���F�b�/��
iK���L6�m�VЩ��~��<�8м�h%�X�hF6V{�SR�9P�pDMN!CF���%��zy���_Ƒl������i(b`Ҿ��zlM�h�� SK�D��_m�l��ݥ|�kB)��b�]k�֒�t�FxgfOJ���o��[:wR��tD ��x6��7z���C� �UȽ���jz�οi���?�^�d} �#ޣa^=���<��\w��4�ZK����>�kU�Z���ⴡm�B�R�ik�
kE3F�lK�Xv�|�k]`�!��LJ�R��䒽ʙ�f��;�r�L�@u�hV�)������I/nw�hX�tэ�c�{�Ɩ�kXh���mp���y�,<��C�����w��:�|���G����80$Ƭ5V�Xi�=ns�(��,��p�56�ټn�����9N���Q�\h=��"����i���U����a���vdrV�)pҶ$eW����l�f�&�L���;�K|�^��}����?Epф����U@3�T���]����(`KI��O�l�$]5瞚��U13.b
���5�U�m��p
�hT�^���W/G�z��&�u�,JX^��޻o!�	i�K0E?D���l4�:ĉ`��B9��� �u�/����{�Q�֖���������IhIT
q158�k�X�LU Դ-i�}�hָ���+j����w`1��=˛@K4(r�fU��\9���C�Ӫ���;H��-bU�֍j؆�g��%���mn@�iT$�zK�(����ӄ X��IU
W%,/4�%���l�����q%-"{߻�Z�{ ���L�4(k9 ��o]��d�S}��\�\@*��;�#Y�46�i*iD͗����N���-�s���H&`-CF�(e8h2<ZtT�N\�sQb���怦-�%��wީ��q�7�1T�hM�hP�%��������:X��D�b:���M�	HQ^�&�����]e�کD0�[\���lP�kK4�`�� �ߏ������JϞ�]�C4��*[Õ�Ms�aܶ��og&qf�:I���C18�n��A�t���uY�8�8��f��+%*撦^�h9�h3vۆ=��m�C9(��C����@%Øz톭�e�wPS�ݵ�<�:���U�QW�d�N.,0��:��ޱp�a���ݡ��z�k��V�M9�<�)<��A��7.��^�m�D�v�VO�u��n]�Z��I�����tؖ*9-�)nѓ=q��X��ڳ��t����a��[6�����n����=�y�xr��R�f�k��m\�n���h�+�O1�3$�N�n�]Bi[��Mɴ�u1ˉ����>t�~\i�P�{���&��͐V�kF8h�^�z,l���*chR�v{�!�9�3��>����b^a�\����������p�|�k8�x�cM)��6�b7��n(6�U�K+���{z^�bT�bR�W^�͂�?7��>����8#���Kw�͋B��S	�4C��1�\T�2D��6���K=~ػBƔz�Sb6�}���FBp���9�!��M+sP+i+��e����#vWKLZ��k�(֐�zZ�4��"�s9Sb8��SA7�e.��v�bG[h�-no������u,i^�K��V��� ǌ<�w�]ߦ�s��b�.<h��D��<r�#�AN5Qh1����+hVͦ����fy�z#K�����%�`V�����{�hX�[�"Z���rG��;5�4����(`ToxGw��/��c{=ص2,`%��	[����̺��P�jjl8��ey�إ�L	`>ƿ^nM�H��5lQ�������Gȼ�_��ڽ�@�8ĥ�|�Ql-�#o���{!vҶOb�KP�4X�1����L%�E��1�[A�K��ad��H}u�ڏ9���� u�{m �v��k��e��;�f'�dҒق�m���3S��u���J�-�T�r��[��z,KZD1c%�j�:�?_�-їҦ���1����E�bcwo���X��H�2�;*�Gs/fˈA��1*b���]���$�%�8�ѧ ���8��@[���A~��ء������G���>�޾�P���)��n��[����\K�ڨ�Ѯ&��ثl,�p�.��^n�JS3�vf���<?���4�λA�D0��˂ֱ�A�o���vN5�U�y�R8��p���"ձc��������Ɠ)��H_`P�U�s��t8��A�a����s�F\$����c�^�[�K��y�j�sa���
�sxe��y�|���O�g�׹B'��]��8�Nr:�l�p����d_&m�� K	܉7�i-��� :+���J������=��Iw�nm���X��cd�9��-j� ��*�ANXz��M�Y0b��q��l%����q�,֔�jt�L�<^r2 u��b1�3���V�{M(�����A�X:�F���SKZT鍔��p"�������b���1�H�n��9�5�1\����a̞��k�	kv]��c���X�eu����=�Ɠ�ɶ�'�[Lh�����e"�֗�y�㬾�����������0��uƽ)pv�g�9'�n���-�vX�nG�1�l��-5��ᚨ�c�d*a.�KI���d�0�iSDp�K<�~��b��ܸ�MM�c3;������'��9]<�d����{\����C�M�iM�$~�</c+j&��R;�0���95�o!��Ս�k�S��2�q�̛��)��ryܨ�=��"�֊j6񎽻6�x�m~�C��B?�� Z���Dw!�����pF����Zҧ�:Ҧ�8��C,"�������\z]��ZX��ҟf�M�2En�g ��i�[%��߽8����?y� j�neJwW���k����C⩑���O,��a� �~Ds7���}d�(É7���*�nū�8*�R�mS7�9}t󌿼��U�ɴT�CZ:�ۦ�eT{}��5��p�K]h�*��q�&���r�7*����L��^�}����s�ZW0Gf��}|j�7�,Us2��M�����c�SE�l������-��Ծ5,��j9Y���FN��.�\���n����*j��ݼ�C
)�F�M9�Q֊�5�u��cǪ��z�Y6���)h��RҶ�=�h���~�δ6N�MA5�2�@�׽��$
�Ҷ7l̄��o]�%�F!D~��x�n;��3�"�MO8�q�}z��;O=��9,�^��b�aj�wK�/�:���,���L}�����!�B)�5]��V��eKa�q֌�	����4p|}h�ƛ)���:Ż�뾻���]���x�5����z!��M��f����iSw�L��{�IP�n��A����\�K�%��	���A���/{<Uv�.�qG�}��8��;C�:
`C���wBȞ�/���vԳ�<dz��3�b�טj��Շ|ta�?P"�m�	>M��d�$6,��Y�X@���	f�7��fv��q�<���ۋ
f�5�U�]���C����$x�>Y�1}�{�b���!�1s�SA=��Y܋f�b���%�����:n�|�*J���M�{5/���?G��sx/Knu�uг������E�0��r�r��޲���;iK"�)��R�K����5,�W>k��TbK��Z=�v�n��4mg���l��k;�Aa�dR6�r�c�_e[��ڳ�:9"�l�w:q+�Ǵ����re�{�OB���x��5u�V��5���l�����pD�F������CQ�_��0b��Ə�o�Y�J�h����y�h[8mKd�C�C��5�pҗ^�v>�W��y?p��#��.����Г�(w��rY"�\����T�樅os��9��vp�"�!n+�9N������m��*%;�ִ��Ǯ��}���kZ�l�w�>�ǹ��Ǜ$��6���ن���N�V�Z�F�!e��������Z�ZѬ��7D����u��ҶUE+(�%^�\iG��oX�Oe0l�<Z��+�黵o�w}�N$���<�q�#��@O�v� {+4�m����4D?g��PA+0��0�j%n|5����d0p8��7"�P����W���"˜�z���g�
�D}D�XF����p b/�3Y�"�P��U�ݡG�A����y�f|x!D3�D�ϸ��zq�ݚe,�w� (!i�ۜ���������:bD�S@=
�w�n��X��{��)�u��8���/�^��r�'\��^D��ڏ6�zM��e�ɝ>S�Bt���)�0�bj����z�MD,�e�@g��M�a����w�b&~f4>���z�O�j��E�qY�%��J���8�yt�4Y3u�{�5o�~��rx,]`2��#y�$H*���q��M�"d�I���u�s_.*�'�E�3f��J&Jq�..Fbİ';�[~�cʜ�4�U��bs��m�Ͷ�[&�b�����9{s�0:����z:�K�$�:��]p�+�y�2m��ƞ�y��9�m�:N���;e�wd�T[������}ә,�sU{/)�5NR�~��xeD%M��Wm&��Y��<�:��;	�H%�ֺ6p��˞ڻL��͕ڸ�{C�]����m���g�D�#c;a����\<[�+rNŤŝ*�9[;=���#�X���r���L�6�e-P���T�B���oJ4��j�{ﷅ���-�5符��͝,�|�����3�}���ݳ<�i�$��Wv�h�O�:ѧ���'ŏ�e��$�7"r�RGc2�U�J`���}yƆ糇��0�;�<��ny�d^F�:�� -���V��V:�3��jn?��B�����n��0�"�E}�[�u��>M��z�>Y|�Q�Z:[i�XQe%�vāWqp��|j��Ķ��T��	�8���z��b�;�z�vvv�S��f>�G�ӌ+7q�f1F�NՂ!��\����A�$pU�d3�!�p��/;.�D�%�5�$�7

O� �:��5|���-!��Ѫ�^���3�oN��1�wq]����ks����{�}0`�ʘ���-���6l�?<�����6ZFmh��[�����T���f��q?��03|�b�8d@v�`y����J�����A<au�o+X��XƲZ�H$%��BEs�j�����vΛ�p&ׄ����=���n�q�0���nH��N���b�k<m���^�4��XL��:>����{��Q��EV�ѫ'�ym��~�Q���0������#�_BF�n+��̋��t�qͦڢ�Q�!7-�:j�M�T A���?��wH��29l��9CR/���f�ɯ��|�W�`N�U�ŧV���	HE��V���}'%�t�^����u/��o�YFDƃ��� aɶ��nlR����<�Y�Bj���L�=�X��j�h�惫=��Z)��q�������Oc����B|w����Ƃ~yک�Z��u�����򑤜�	��m��}���������7n�G������F�I����[���^f����^���*���8��J��W���M
8w�;��􆑞Bj�t+��oty��J�<��ڤ�",���d��1qݏ2�v�"��݆��NԠ���S�w}/�ʿk��G/F�bN_�ޭ�E͟��}肙�u^���؅Q4шen��z�|[�����+q�ʧ �V�ɝu]k.��8:퇇�;%���=oXƐ�'����l�H}�W�4����<�#�a�Y�Oe��E���Cn���NU4���1����E����r{��sYB�d�ﾄ��%��R�.A�F��h����{cf>�����)��n�Q�k��ʫ�ުa^�ν���	,��_{EU��O�B��'���O&����V9��MF`��[���n�~B��k�̓�`�����o�6/����,�l�\��z�yxCÔ\��;b����r5�.�Ž]0�QJ=������t�o4�uIۂq�a�_v��6v1��������[���d]>�5�����e��#�ib�S �Hn@�)�ô\�)"EU�<���z�YV��^G��ㅚ�ݞ�?qjxe��������uQz��/J�D�:������.�	�j����H��WSr���}&<�!�s��ډ"ma��w~�՛�wϷ`��E�Y��oy�8���u�w�샵n���E�n����i&q��
rg��ΰ���m�Z��qZ�՜�8���7j�w"<����V����9�/~�����J��|79�>��3�G��4�?��D���a�wF�{�H���\- �{%o,g�8D� �#.DN?v�h�{ݟ!}%����.)��d���s��O�E��$�2|.z�xc��T�wq��8����z����5���q8d��#�>~,H�W�⫱x蘫k�C�@0��rێ��n�P.�۵)V+U&�STKFW{%�T��.��~��1�DaA�$-���� �]H�R�7�ͮ[�fM�upڗ�*7^������#���F[�r[��]&WF�	>�g
�&�Q��;��,��3��;�ɹ�n��yx�d9��DT��	�AO���6q��^�/S����z^g�����b�0��S�x�^�(1B��ܴ��x?�r�6���Pb�y�R�}BW8�4Ү�г�x7$��^�����y��^A��T_���ǳ,۫������03�� �������s96z�-�c����b��p��n<&FH�,��D0L�vظX0?qU�UKov=�f�)H���j=����<v���e��7ǾQ�:����%d�����bI��Q�Wں��F��������R��t��>�x���[����~JB�������N���41�}�x~��%��h��%�,��g/��E��$US�?��'k�nJ���H)5�G�o������Z[�m��.<���ϧ���@wL�9xnzlԟ3�W�S�m7O�i{�x�f��E��ٺ�}u�J�*�xɮ�H��4��!n7���g?M��w16�ז8��sӋ�ȑ�3]Y�ڊHl��2���ۘ� $���� �BK��$���HI~�HI I	( HId �BK� HI� �BK���_� I!%�I	/ �P�HI` $����I	/� $����I	/��HI$��� I!%�I	/�b��L��̀�(ϰ� � ���fO� �y����V��UDUR�Ҫ��\�.�R�R�ʐ��Y5�j���C(� ����"������J�2(�!UU/�           @    (        @    �P     } h      � �::=�����/;9^3�G��������n^^��&ڙ����{��[�w�촻o:��w��5[�-��<���]� ;���j�;�ص�����ҩU%Hvo�������ꭷe�u]�)�� ��*{�y��m5���mU�W�ã���o-�o]�:�� �y[Ӌ��ᴷ�w��#Ms�\�{��x���s�V#F�m�J�      � �.�{ly�mG�vYϻ����{[m���/j�.����g]o89�j����r�ovn���m����w����6� �{j=4�'=��u�/w�Nt��IZԕM�v����cz�ݼ�{XZ�ϯ�� ���V:��o|w���=�ww6�ǳ�,ĝ������Z�۽��nsex �^v�z��n[�z�u���o>{��V�A���l<k�;��{��Q�sVqMi;J��       {�{>�ۭ��o]�Wv�޴����Ƿ{�ض�;y��)�8�� q�轟v|���o�w7�����[��ƻZבռ��{]ww< ��z://)��v��{����R�"5S���v�j��X�ҺS�[� v{���ם�=�Z�[yn����l��3�q��4�m�Q� ��h��{��U�ݹ�{��y�����7�ӥ�m��NWhJ��H���      � /v���kk^=����<�����kL���ڝӖ�^w�᭛�\}� >�*��E�oe���ׯ\wN]�ot�)5�omݣ;N� >��*���n��W��w�: �	)6ʕU���z��۰x�^�m�7��=�v�p��{m�<^���v��.��u^��[�ݽnΛm�� p�mKms��Q��dy����U�k�o^mMa/閙�.�I*P6�M�   z     <oe��ׯw��@� n�>�G�w
�w��:>�w�� �ڨ ;�ۚ���AA���r��aA�Q���y��!DA�^ � ���k� tt�o���TT����s�+�> h:���� 
�[� ���{c�c�����(d(�Y�SG�����{�u��-�0y�� z�>�^��a/}���`���y��^0� q�t(�� ����*� O�&D�J2 h)��4�TD ��ʥ@J�  ��D�J��@OH&�T�z����O��P�����0~*��_�����>����2�$j�w+*���2Tu\�u~��%
"%&(P����(J"��D(��aBJ"D~�BJ"D�%
"B��D(��?������ɖ���`5���w%f���!�9i`A�z�e�B-���h;eǖ��b���l.�l�pJ+-�.u�,�	Rx��J1*��3��5�xq3͘t+����e]�Njπ����CxI'�*\��L��16��5��䏆^�Q+�9�����H [��V��J�b��)ųK���6���IN۹	��vND*��+�c��zqQ1�[3�a������d��=W%7��U-t�S��(̖�ql�n�8��s/Z1�+-��r�4�c�p�9��X�*hi����-nSn�V�:6��.���a�N��YhYV�Ѧ�-��x)�h�7^|��t �jJ��AwPHF�n�JeŇw5�Ѧ�թu�^6��T�7z��A����ST�:��!l�u�y1���|�ԙF*ʕ�fc�C*ˈ�������{������, �N��Ytj%`�7�a3%�aң�kS�ced���T�٦`K.Uq�Iu�Σ@*f](���F�r�ɳE�1���`&����&�DH�7��]�{�i��a��GR��f��y�C�?��!F���Ȝ����.�m��4�-��� �{�`(�7��r��F�\,C
�1>�	R�^Ř��C�ԻXS��w�ol�eVE��Ե\�y�]�m�Mv�Sp"+
���E�Ŗ4au7�(�)z{����J��T����@���7{o���تe�x"`k��di����G1٘niQǋU[��[y�śELx��F:�\$޴�<FQ�"��icĕ�`7pl�ٺ�a�6Yss[�/f���f���E3C{g�N����6���<r�*�kCq7�21�%P��A�0$T'*��w�%�T7���l�����b�5��?���s�A���Ё�'�����⨶2������6���5|��/�l�co�atK�A���}
��[ڦ�gH�Xu9��0�N��e��eӲyבmAwj�u���u7���Z����+e�ӛ/i�P�j��YRW��%�&��c'^Ѭʅ�k�0[�T��{*D�E�	x��d��YSS��U��II-�Ejj��K,hk�e�w�2��k�+����̧�R�]��V3mfYT�F�M�cV�%����[��\���3n��F�j9�,�$�n�خ�:4Ƹ�ᷚ��c"�("��c�w1)!�V��;۳�`c�]h��ڇ^#k/N4Lz��t�]WM]�L��qu�[n��w�nY�	AM�/�%�;E�ћM�z�^G��{[�2�6�i�z4��#c.F��j� ����S meJZ�l��"-�L1'����)��V�Ţk&��g�K H�5�ҬV�ܡu��YB�J��lJ���a��]��[�ى×"ʗ��AM��Hm�66�9%�I�](�)�
�U\!�����z!��G�����73���ln���� v�H�6fK&Z���X�@�(�\h�1�f<k*mc�(�4���g4��b��0�yr�ݫF2�e۟fl�M�b�O�)�%5��F@W4��O��54S����_a�b�ܘ.���.�����!eåUԀ�Ԋi6�[�����}�3�l��ʠ��S0S�/3\��b"�°K��(�LzM7�Ǩ����#h��9
+;Tk�y.M����ɀވ��Y�Μc�ѬWw>�\��p���5�2�CW��֩̽�n�nm�Lі�[lR�K)^�(Qp����3(+�|�2wBy�+&�8 d[�]�S�r*�"P�"�9��w�w]4�K���ӫjٙzeʼܩ6U�	L���`��S�eiU�t���.bJ;0�R�`d�b���id5��a��p����\���ԺM�f���Z��N����5Ki�Y���PBn`���RR�H�N��Sʼ�@
ͦƆM�N���FN�ytYu,�8ԄKw n��0��n+5�Mr�Y�vX�3�)j/[��V�gE^	&U�@�Oq�ws ��Z;���'��м�P����؅-.�3{��J���cj�Y#Z��*��0(8qZ�z��:U	�y��*Iͅ��zf&�PQiܠ�މ�E�V��ӆ�+�1��������g%�ĉ�:ֈ��u7^#t��/%ғVVP*Gd�EG6�2�v�Fp�D�
51㙖�3/m�Zʗ�D�5iA91	��;��R�{q]VFn�]C��R�2k��l�[m�2��`�<�(4低�2�^U��Zҁ���!P���O]*��%;�j�j���
m�F ��CdܱYnc��U�Ę�u�࠲���LZ!��OgF���K�4C{x`��νE�����Ż��[;V>��u����������n�n^Y�5X��^��ren�Bk\:�4�K�V/!�1{j]Nͥi��Y�d�0�7//�Gkh��p\"��Un�jA�bi���^;�O\��U���̼�ʆ ���ڀˉFV=8f'y��#�A��-�)Xr��[k��W�
 ���S��-�{������ Rf�Ymbf�Յ3%n>�,Hn����c$�@�Z��uj�q]�I����H��������mU�AR�L۹up��6sʐSee�mT zĔ���	�v�n�C�wɵMǮMoה�-F9r��j�aн��R���J���)�
2�����ַ6��
�r��q�u�̧�Ry�b�BVAi�2dLTR0i�I�d�$���]ȋ�4xt9c��Gn�#m^�V��%�ܱ�%m�27���7eث_�$�߮Km��]b.E{��?A�!�lm�d	:�L�:��h.!M@7�F=�ī2�{�#p�jS\�l�BH���%l�e) �eh?
֚��ٟ�C(<�Z�(�� -e�/R�6�f�ƣGc4�J��&$˹�֩@�&˙��'E����0,�	���ҳIZ_��XC ��Z���+y{Y���H�u�e��.'�ޝݴ�R�AZ��N�i+�,|�X���]1Q�4�[�N_�7Q�A�+_ѩ���B�c�a�5���M�$t�7�3 !�Fd�2�ov`?Z�&ܕ�
ժЦ��m\�U)t�.egƴ��g<1f4�����}�ޗE�vgMmX�C�w ��e�Y��T]X��V�'.���,\�x����sIs\4�(��if��+d�td���u�+G<��i���a�%)M�K�ݸ�r��J��B2$W�0�7o�%PW%3Ml)I���D@�HM9��^f����%T9�^�,�ڭm\�8-^�� ��U��A������")��w�]�p����ױ��:� ��n�.*��0��[�zJ�atu��X(迖��D]E5�V�m�1�YBlK.Ƭ�e���{�V<V4�`��U-wp��f�7��\�k��[":s��B�̫�M�z�ي�nz�m2���w������ʲ�$�T�V�:*�p�0g3Z�0l��0�Z��E�\�Q�Y��M��h1�͔�����θ�Y�d�Uӥ�|��ĨEu1��r,9*�4%2�U�RM{�(	6��U��JFB:.k�%��̭;nt�uR{r�fn��dy���7���niKJń�{l���N�\5d�j=�je�F#��ɐNʰ^�+wb���jc� ���A�aٷ��8^*���:T+�"�v2��������4��CcD����(*f8v���gt�6�R�B��X�,<e7u��ɛ6�*�����bn5�6��\��P�oa�N��b�����슽���㗃Gh�t6L7�˷v7R�Y����dKl�v�͉#.��ܡ5<%�S6�&1#�eެ�hnSS�
�h�m�����z+kZt)J4��4�k��2f��n�`$�R��^�je�ڗ�cjC>��IL��`[æ��"-�[����l&))�̣Z�ֵ�.�˦=L���3�tL�ᷔ7�D�丐�,ś`�o���X�4��΀��E�mi�R��(e+�D֪82�۱X$TK��
d�vmbW�t:IC���׎&>E�G;�:�ɱP8]<���j�%���Tvi�7 &C��l���7e1��4�H]B:4M*�}�W�Qgd4h�5#X�ڑ�H�4��@��i\T�!{��[bM�V"� 3%ѓ~�Z�����.�cׂ�kNʁ��U�n`RͰ��;W#�2���6�09k-���,L
��KDwe=Iݖ�>�[�q�&[�*'@����ہ�9L��pca�RDN"���͵�Á�1�k�+��3�Ht�,T�ɀn5c%*õ��u�6ӻ�{u���0��/Jn�9x^� }�lXђ�/�%�����G�$q;xҔ�܏^�_[��I͔�Bͽ0n�w�~�U2kf����4�SL����0if�������[�]�gN*������0����n�n�-a��6M��~MTs�mѽ)��6Nְ�%q��k0Zm��P�Eȥ�7��.���ve�ؖ���uO�[�T����k1ݨ���8v�1�,*|���h)��O��:�E᭺Oaݰtn�8���^�ڰՓI�%^�܄ӉŲ�%*�a�:.�mE��U**n'wR����e�ou��ϳ�[�:*ȧL{��KQw���B��w��(2��nV��[��N(�Q6��ɷF[����h��QK�D���Cj�y�T*J�Xu<zt^�G[���I4	�w �w�w�!o632��hV�҃�sd��X����0o2�;e�*�ͫ�,�@�l��h�KD}�̡�V��pe%��n�F�ڊ�rX�4�%��E ���(���3�7fȦƴF���gŪ�n�k�Kh2&���%n�?h�)��r�ћ񩹚B����.���j��l闭`�V�3�/7���S�-�b՛���a��%�:q�#o0���QVl�6�VȁA�B���jeooQ�fY����������J�&� �x@Z�a�z���%�J/6�x������퓦��.�!�{�ՑZ(I��-2��n�V�U���G�Tٲ�� 6�HDHѐi��̔�;��̧r��R��t��H�[u�9�mo8�ՄK���*)3]��C����%W{�՗�w1�Ҳ"){���Z��5�d[/���R�,��q�9���8�6��n�Θ��PJtUar�6�T*��EyR�ś5�jcWX�MD�#iW[���ѓs.n���k^kY�77�yq]����i��-�6Ju�e�u��yLR��%ne70&�Yin�齳���td��졦��L���ۘZ���w�n��t#�
O�M'�t&s�rL� }`Q� ���M���Q��7�&�-%J`�-�m5�m��%3�l�#a���R�=��2Z���HΩ��3y���'���(	,���(��B�,Ç>�CYYSi�+*#[��[�qކ�]�!���:�J{��}�6U;ʄfOz\e]7jβ��B�����#9f:܊�j�:+��>5f���kˮ�Q�G9r�]�T�r�m��U��[#(�����NR�)7g*��T�T���aۛ6���pa�F���-#���u��2�i�IJ�j;@��n�����`*�ר#�Bzoa�/cW(h�i,XJ!�{7okoPT�Hm�4��:JIbm���X�`)��9e�R��ܭ��fؗA���V��"�y[�f�6j��n����jƲ�:I�Na!�7-L�����b��0`����jzԄS�(�)�h6Sz�C	6he]�1I�i˳�
0umJϋ�$��0;���l[�6�L�K$E��s.ɱXP��flܦ��� u�'�iF&X� C~��Ջ+,D�IJ�Q�ݙX��1^�Ƿ�)���DQ�`5/f�Y��3�|�7.R�u۶v[7P;aJr^T�3�h^%�lݼ�;t���-��J`���[�k����E�F��F�sp��o]![�᷉X��W��&B���w6�Ը��5֥[3rH�2Kb�9��e��;%Ŕ� `ӯ,��*!B8�,��a�gm��\�Γh

��1��}�a���P"��n�BN��,-�[
�&�v�V*�n*���j����EV�5f5OKK4��X �,�4M�L��i�%�/����L�dZ�PX��H;�3^�x}v���)�f�P3G3NYʹp���o	���,��2Q�h�P1ٻ3�oE0�Ř�n��o����v�1TU0�T�v��Y��[��t�Xa�$�hyJm]�f�V�q�5|��,� r)��d;�SI�I��x-���S/!�E��������KN3-��@YUp�oc
n=�]dvM�,[�K[ò-L��J�Dsr�P��Gr�N�md��dݥ���lPPY��"��	F�˕l���(TJ[�HQUJ�r��)�rebe�fcW&���U�����ՠ�J"X���&]�W5s)�Z�1xg=S5����D0�i���'
��H�r�hڔn"6j0�oLñ���9fe\��U7$)!��p�x��dG(fB�,����r���?<�	� �Քv1A�`����(��U�l���[�d{kJݣ[Q�/J8�C��!�T��B�Đ��4қ�-��������k;8jD�.iٹ0���2m���Y$�͢v���j:Ë��G��ULD�PQ�Mn��^��Qj�M�V���5f���O+#-�p�n�,K�ۦY��Tq�0���ʒ:�Zw!�kp*XM��в���E��9��u���Vb���v�[W5�� f��v왛��7E
�!�����[�˚���Xv�I���:��ڀ|�=@���N�â��Z�b��l�'��^htK�]�re�+������c��:n���/L��%	��R�	*����:��a���)�ٵ��^^C�����,�룜�An��M����ն�[����;��n��r�F�O�Y;�Ɔ�nF�sWcu��nZ�s�<�ӱ����S�[��'�1�7e���{\`���;[&P�:�ɯ�x����.{F��s�6����7�ً�����+��{=vǈ��α/�nJK�]��GM�u��b��m�۷w8���ˌ��R�gs{r�'q�kx�S0i�4�kbm��[˪bg����u��W��I�s��BwS������=����l�8�5�Dx�ӻs���ő��v�ڊ�\}GŶT{�7n�˺쁢7�/i���tٱ��p�=dCp�r�t�N�ˣ�9�܁��������v]��A:��9}����6���i�KcNn+N4�;��{ �n�)=�v�Ի�ݳk�5m��;דu��Z�)[ێƍ͚���/���y��K�qӷq�^'�J��/m���x�-�p���x�AѺ1s�F�v�4�O��N�We��m��'���s7;[2�**�݄�\�u�є㍎Q�m7d��f���Z7)T�e����l�u���}��!�_��s�B��Ln���Í�{-́��!�<��p�w-�<�$���F�UKe�Wm�����<�x�]���������J��,v\�u���Y�Dd���׉�v9� ˽P�D�<m��}l6'Þ�rO�z��N۩��:m��{��]��<��a6�M�<u��]KӸ�x�xlG  ��9܅f�i��������q�Z�ݸ��[���oX��oO���f�\�m�Z:�������Բn�o73��I1̒Zݍ]N��*gd��@�f6�k.�v��7����aSDg/d�z�88㫨��1�pI�Yݗu�1�ݳ��T�m{9��g��z/)�n|��q=�S��m�8�Ɩ�������xM�ayՓ[h���;���.b�<<.��m�헵�Sr]�FK��X�z۰�L�rv3�"��f����qZ�d�mr�N���c���]w��z��M�cg�1�q�\j�Zp�X�`�8M�m�٫�of;u��[&�s�gF��-ӍT��θ��s�G�`8��:�lަ8z݄��1�lݞ��M�ݤ����Mm��/d{=n{`;	&�M�b�(�Xl;A�N{8�89dnk��xΊ�7n=���r�vȚ�]�'��f<u�"|�I�f[m�'n��p��K��n�3���J�<;�g����'	^�b�?
OŋIN�����7��i��� ��vC��bt��.�Ҹ����1�g[�c���7Xt���5�'gF�v�ݻ<A�6 =�f�Ǌ����^22r V�S<.��{�pqq�������q�N헇��N��۰����,0��]�۫v2�ۥ���gt� �hڎi)���1�wlY�vV�x%��6:g{�Fz��nfގ��u�c��N���OO�i��r�cg��rx��,�Ϭ��3��R���J��O ��(�]���m۶�;M�=F���:�xl�j�m�[mW����p����@^��{!�mY�㶑���4�N[�FFc	��3�B��ksN������؜\>;]v��P�`W�1�7�b�0A �������b�ы�����v��;p��d��E�s�����vE�c�-��-���8m�:9u�p\��q�'c�(��\W;����]ɋ���䢕,�\��V��}��gc�&h����k�/7Z]�ݫ݂�p�|�=��v�G�Nmt"�B��i��=�����2�ӻN:�Χ�5�^��۞y�7�`��&�:�*�'2���۪��Iɻ��W����:ؤ���Վ:.Cf��أƻ8Iϝ��.�{n� �N+)�d�ÍړJu���|����M���˭�^\��p>4������v3NK��-:��h��vf���v�k�ܺ7oY�<P�m�nc���]u��<6����S��sdld��Kqs��@|�ǵ�m�/;�F��6,��f��ܚ�wkm��Ɂ���9�"�g���yd�������C�%��N3ێ�ji�Hw:�6���^�����n8��t:��^5�v�oG�]�f�{����Z����t��3\6۫9Ytg`��v8�+��wv���C�̇1Z�l��E���v[WK�Ⱦ���F�m�+pƓiʗ<&5�q+�ջ��ǝ�F������nEV�:e.���Q�}�t�;½u��nWL�xy����X�͋y��\���Z��NX��MJ��mN�5�W<���Pt6g�x�;��nxn�4p�y������jM[��"c����w�x/���ۜ���k��lv�j�NѷE�tvӭ]��#����3g;��Ǟ������+�ݲ�l���G[nܛ�ym����)�S����𻫱�/�j��*bؤ�p��uv����EC����9��&G��Ė�X�n����㊮���3�=A�8읺5jM�3�Vc��nwW
`B��8��6�gW3�s���<u1n�} fq�.E�_�ﲻq�˧�sn�[7g��ޫ�]�ۓv765�'[s�#Z�ۦ�ܝu����qn7#�6�w[y�ە���v��Y܁��,��ga��-s���mv�=�uoh��c���;���8휸�xs�unq����⁜�-����n1��6��綸y�Y���PǬ��u�@��<㫝Ot��1;��"c�O�k��U�n޺�s�94{Ru�]�Sn�v�ݓ���ci�5�P�]���B0�[l�;p�tZZ��V ˻�ۑ��ܗ�cl���`䃔�Ē�>��-����/;����8f���-�ޣ�� g%��_n�xN���:�9����;r��2��g\>��V���O<�`N2u`�5�Nӳ��Ɨݲs�������
Vk]u��'[��1�=7;]�؟e�<��."szĠ[�q��	��c��M��5`�{RͶ�Z���X�.���<�ə���.�R�g>�Q:ST�����E��vݱ��]��f`x�����gq�^^6]V�=RT��t�ײ���T<o�؏v{kZ��Wg���[;��"rv��6COcj��i��/'�֌蝸�@��|����_+���ro���gs�!Z4��&����۷^��9����Z�y5�A4C��I������K�{Q�.�M��]F5��{h�t�I�y��۞��a�ja���c�mu������zS���m��g]sv]Vf.7[��z+c�W^��ۍ��]���;Y���w��	��-˙�t��^�Q�j.���2Z����퀕��k�:�.�rqoC�n�p��Q'nw�5�0�.����;����/�M��/�:��c���������jx��f�Ƶ�X�B�q�\�����]�πԑ	�0n9{���kn{nCV�m�8� �,�u��s��y�'m��c��t���iL"���3��!>�d�$������aN��/Oa�<о1�Yq�.��m�us��ø��m��dZ�nވweQ�8آg<Nl�S9���m��rm7gv�N�[�Y�ۯ'VYsci�6�O�躻p����Ӄ6�nݙ�6��r2�%p��6sp&�hx�Z���n�}���ch�d��6�rJ��m�R����=��m9�qY̘�����O9�t��=\�k���*X�\@fMs�g<[u�+A��7\���[Pq�[K����{��jzzg�6�ɺA���@�9��������ࣈ�����R�+/�sb.j�)����ط�������n<% \ܛ�gͶ�����s�;nLn]X\�gMu���qb��n�dQ�]�s�J�X����m�%��X���s�'UjJ9�=h�+��c��x�V��.�| q����H�Ͷ�и��W@�G%���X1��q������$���4���܏n�����۰"��l��r�U�KXmZ9�[�xmkV��n�g�]����6�B�l>E�c�lgi댎���Om&b"�/j���>�����<t�%�o=&5���ݳ���{{ܴ�vhɗO+�ӧfy�#������A�V��nV'u;&Qae�dLU	�h�BPL�P�z���Uu�>]퓴Jٷ@8z�x7W%��Mlu�ZMd�l<�{7g΂�;n��xv1�앨�bM�*�>"8��H]Au�<I˼X�9�%=ɹ��_9,���"�A�V	����[%����z��Į�=tz���=f�n���{qt��m�8$��f'{=c�l�, �����p�K���qh,�;f���:��s��6�c�ݷ6��E�ݶ���{wW��&wd
��f�r�&y	6`�nu�|:(�#�]�=��Ns��l�f�sWm�wvnJrr��ks�:��r�U��+�W�8G�q��s/�۵)�ƾ��!���q�ݻ�s;&r���ۓ�0�oG���k���<��`/���0c����Gl�m�������C{�v*��Of������]�+��)�{m�\<C�wj�5�r�u���ݻm�g6�v�ӏ]c����r�R�������<���K��gţқ#�[wh[t���8��t����ǿٹ����x3r&|8�VxCeS���N���y8{쾭cV��a�Q�q�*���.6z�w�݇��l�7\�g�9�b���^B3�mm���w@+�eڦY�V�J��{��Wr)6�1���Á��k��s��^�c�������;���y8��m�ۃs㮅��N�ڻlv]{j9�@�.�;��jgѭ��y�a�W	�wm�{*')Ru��n���o Gng�;<[QC����:�Y�;<���t�v�'c���v�;ORg�hh��^[�9q؅ES�Ӳ3W0&���i:i��8�Gs��B=�s57���m����\�<��e;&䭙zWE^���v8��ńw�.v��'!�hx}���{�B��!~�D����Q��%
"I'�{�����1N�,꓄� �m�����\v��u`��L��'3�6z�am69|vޞ�ݻbr���Eӗv�A۷],l웣��7n&� ���p��҈T�)��S���u����G��{j9�<�v�焰���Hz#��{xϗ`�5u�u�!��+@㎊
�UAE�����(�üm����L^٭�=wg /\�ku�D��ggu�UŐ��gs��5�d�mom]��!m�k���7�[�۳�3�i���d���J���oK[����|�ǝnf̑��n7o;�cJ�v�Z�3b�W�j�u��]UqY�8��2">۰��M�<ۇ;�a�k�[6���Mn�m�q���wc�՝���n�<jv�\����! ��Zvb�cnAm#���Š�$�݌��s�Q%��'b�ouٴ/���t��n؋V��+(I��mu�P��g��w�uL;Iũ�W��JXN��t����|b��[�1v��p*�qE���.�S�g���]v�W�竭��v�u�98�n7M�(ٞzPYl�V��۞���ڱ��j܇L�Y��vN��q2nm˙�����ٮN��ge�G,J��M7&qY����P� �tu�ۇ�qqYȞx�k��,`��
8��a����v۷m�j��jl@kGb'���pqsͪ�͉5ݸ�.�����������������u�	gwl[��8����c�Ơ���.�.�{uǜ���e��rOTq��6θ��oS73vGL:�q�cz�\]+G:�%7 k��<5�{v�X���4��gsԷ4���E՘����f���n��7/)X����pz�@v�E.6;e�$�u)���O�;���͞ūom�8푌�Z��b�q�.���� ��sڈsf<�C�j7pGBb�z�X�c��c�X��rļ�7nɫ��U�E��3�A��p{I�����n�.�s`�d۱xv��u�X��=���<ö8\�L��Uj���$�DBJD(� �D(@�B����� �!DQ
""���(P
!$�W	%"�� ����!�`�s�c�����<t	�e�F8��狎���෋l�	t�^v����j=�즺ӫ���ɫ�l���i0n5�]#����.:x�+�=8���R#=���:�	�8;k�:���.5��S
��X��'!�${>]�t����k�g�P�/�ۻGnGv&w��ng�p���N���'=^�	���wu�+�!�cs����Sl�8x�粋� ;��z0b��ڒ

6���K�?��_���?VJmF�Zfd�#R� 9lY<ڱ,�)��.
M��B�GY��8�l�kJĘ�����Z��I�0q�b����l���ȹ�Mvx\f����rw~������ʕDX�m��f���������R�h�X��1����Q*
<��H��f�,�!�JK#�i�yS���]j�4�3���wV:{Q"z�,��s�l%�$�-y[M� ��j)>w�HK��� ���τ*��W6����:t�)����ۆ*o�U�Q�T�X�e�,�D*���j�8]e;����������^.�ZxBn<�q����m���r�6�W<Ke�;�\,+$dp�
dp�٪ip�raX��$�ow4��C�I��"�(�'4\5�4*��J�U�>W�'�]ЖxZk|>�ŷ8�;b
�r�V)#��B��P��������i�4����!K��3���[1�k�3��xK�ƫ���J{��g���;���擩��h�e<z�b�q<r��*26�ޚ�Ӊ�SE����%��u�d�ۙ4��ܤr%s�����tt��!4��sټ�%!��ڟx1�IڳYY���L�^8��}���Qm϶���V~)�V���W�ͫ	bu2�
�^�}�!�'O@	�;V3�xԨ;�s�1G�,��h����p�o'EyԺ�����y�b*9%���p�+&��b�yÁ&Y�����p��*j�'[�<�+���n`�C��1vF���u�ӺC)��"��*�%T�V�(���[tN�vߥ�U��V��٦�C��Z&\uc�d��::*tٙ��}�>��g��	V摔��J��o;��0m�j���3����ՃYWGm7]�Ԃ��J$Nwr�J�%I�fvfP�NJ*U]�H�H�w}*(+�^s�^�%h#��}�+���p��%�F.��Skp.�Nũ��Fk��b���s:I��Y�XT����]���t�85��y9�8^���lch燬�3�v)�uڸ�sc����~?#1%�����C�f��M�b�:�"p���iy2�T E���#,���*��QRT��B����{&mU�������;��Z}53|�}�P^{X=�ҏ���Q]�(����H%U�� H�Z� �\��7Gv�P��tz�s�����<��UAMyسQ�R�Ϩ�Z�=�U��n�*>2Hwi7���2�K�MBF��躎�>�h�0�c\���)l��|&Tf�pa&�Sz�(9	�k(�����UޤR)�B�M�[rm�� �,��sԚ[�T�,e�l>������F��v��ep��9��{S�����1X'��x�n�):@&�,6�������B��U���n��)ُ[ܨ���N��M%;A�C��pYz�F��Ky��{�������X�� ���9vI6X't%������F����hKa�Q7��T����*ޤ���z�����hhr��Y,�2��C���ݮF�4�㼀��{��rR�[���Q褝%�I']�G�R�^u�xV��b�����/��K�Z��1p�ӻ֖�#�R����#�nc�է��o7y�1�7"�v���-��Y���T��mV���(Z�V�d��1�:)]]��C��u|����ʲA*��AQ(��ݵ�j8�yiFVw��4+b:�[�t���E"���+Y�[��{�ʎWK�%=�K�9���ޓ�r1�^*l
Ooڵ���σ4Ҿ��V�op�[V�j�cYau��%Hnk�֋V�o������c	(Ӎ�^viUS]^ױgy�j�z���QU*�)n�*�Ӈ�&0��t��@�N�.��~�5|o;�+�Ǌ��n9�X�j�q���mY�4�b.���]�W�<=8����^a*��YQmA�RZ��W!�k����F�5/s޹� -b�3��Oq}�ie�5����vn&�mv=V��K+�s3#��ʸ����|n���f�HP]Sk78I�$�o����6ڬ��D��a����^�ᒘd�0�U��h��P�J�
J���rk9��T�U[#�6�_q~�~�m���R�^���w���]�r��X�����j:l�R�_ R����x����ջq���Gϕa}�=��D;���b���u����$��O+�Lھ9 i�]���zw�M�f�%:^��W����-�XY�㵂���6�7�(�ú>��O�M]t�&�j�l���D��}����S���˯Z���SA�(����Y�\�2���X�9���5-�+&�*���v���wu���ó�ޞ!N�Q��n����3]F��^K;��n�qn۝ͦ8z�^}��3��=<d䀻��K�S�z�Y����F�����X�9�T�LgGN}T7mչ�O��N�v��N]���3�v��gv�$�r`T畣'��l`��#���Gtt���;���u7n�\I�{/��k��rk�M���`}�4�j��}v��DɊ�:�����I0����s]m�h��F�8�bM)H�
�V��} J"3���Zݘ'k{uɺ�]8�u�N��%Ϯ�r�����V�&�<����tn��]�Jbh-W��-P�9��y�@����������G�����~�%r��g��;�=bќ����2�.��zx�4�Vl����YD'u�F���&Ѯ������X�n�	�	V���<�=�˫�ɰr��+���B���Z���I<X��J	:�J�t6����@��D���6�צ�E�ML�5s�ڬ4�p%�\�G�hɈW�$�/^�}��Ѽ&m:]Y�	 Մ��e�G%�6�)-�J׭-s�l@�3r�U�[��j��մ�	��ju����Z��E	��޽��� �T	�WE�����{qW�Ʌ9݃�x�B�7\ŌlE��y�
�f[`�-�Gl�sJ49m\�v���TJ���W��dʺ�^�yT�NX|[�g|T+�
�h��J�C;�h/�n�tŎ>�+��eylS�ܶ�$;�u�M��ؒ�{ұ��Kx�m_�e�B+����ЖIoT��r��;�owW�\���mp1Rj�VB�X+EX���+O��^Z�xH�ɝ;��v�s������H��L2ؠAI�w�F�C��\{��l�5.�~�lQtӍ�͈X�i�v�6{���g��-1أ�F�ʽ����(���+�h�st�[>OѿkǞ��n����t�=�vkR�o��䔯]u3��1čZR��8/뎅ˈ>���T��5�y��)F�X�ۥ�k�y��z���n���'�́�m�C5��J$�/x䜞�]L��#\��]h�s�����@�B�%�??�Uut��J��uvd�vڳ�a�wBm۰{2�鎆��퓶{g��5B�����(2U���-;���ki�Z�1��ξx0��d�A��:���ݽ+m5��$�^zW����m�}!!T𢐣VR���Q�>��<�Oj̶|��p��nI������m�|6A�weMU��ܒ�8Z�O�H����^��S^���f�4	ڍ�h0��fnd�z(�l��s6��i�R�gO�܊��\����ݛ���%2��C��q�t�F�D�}t��̭�Gn/]�[$�ޕ���t\�YoeAb��e+1R���s��^ut�u���K�?e+~z���]�X�T�%���"�z�N�`![k����h�_��]g� tpl��P������8w��G͍��A!e���8x�����t~L*t��o��T�^bi�(]�|�����~ʸ��׎�ep������`^��@�T�}��/fc}t�,9����^�3��H�@�W*$����3�T˫]�v-��~�h�H�SN�	a[��:��*�*p�T�Q��r���߷=Q���]~��������@��-
��:^yv�J�]���9?��o؟�{UbzCOv������{�Y3�*��82�E������=��A��e��]"P�P���n�T��s C}����q�}�ׇ�j���Y	#eQ%��:u�MU����]��*���v�Z��J��.㛁˷�ˆ��7�2 n�����ۦ3U�}�n�����TA+rIV��[|zo�|�wz˔1vv����ws��p�]���O*��2�𧹎�R��ЛVZ�&���mY��rx�.7�s�K(�f�H�s�vWk�Y{+_`5�eJ�h"�k>�&ƣ��V�Zd�F�Wi��I^�ogd��kIkɛ�e$R�mO�ߤ�
K��?e��m�C�:ka��(?e��\�&!���w` ��wK�U��7���v�S�Eפќg�S��4I����mx}6㎝\=��4�]t���C��.f��q[J�T�5J���c�2Ku��Wnʥ�߅k�3S��P�x�lB�̡E��z���I��j$i�=V:6� ��a���l�B��N�Joqץh��p�<T�&e,m�'��7�z�C!jn�;�ul�j8�ށG�����t�T�u�WY��ף`�$�4^�y<2g�ش9�q�m`66�~RCXL[VY�W�[h����`Q��D�$����Ǚ��\y�]�"bWe�����]Zj����(��%�mz�z-u�}���㱼��6|$N6���Z�e�E;�T�O[�Jޱ��T��{�ﱵ���d!۸�'\���3.�پ�d�䡰'Yk��á��]���(u��`l��Ł��J��/J�����{R\I��Dr�6�_�w��� ���t�ґZ]<�t���O~�����k:w��0Y�㖮�v5��Sw�v��6�&�SN�'5�V�0��u<Ǟ������sn+Zz��v�ی�7,��0(�����������qŔ�ɲ��Y�g5��=�����׮�u۟H9�&,q�Y�3����q\���jr����MC{n�����ۯ��x�:��"C	9˶��n�	��;rn4�&���铎,�����m/'t�G9[��m��N����3n���@��ę�4n	�T�2�����,��n��bC�4K\je�"�m_(f=
���AI Ŷ�<Ǉ73C�$�B���ґ��*��cӪȆ���L��ѯc���_O{��u��U��bw4�\2J���멝j����v�ɩ0�b��O�C-��b�)��;�1}?��-~�3±Y�|^m
�X�m`j�;@��ŅL���=��;XD��R�6B�MՁ���1X��	g'�a8b�����5Pw�G�������F��J��9zM^���u��$�Q_�I-��1���w�������q�[�� �{�sY��1�yU�sű�q=f�{|�s�m�H���GP�>���K��v���
�����m������� f�Xڜ�l Wɔ벏�7]k������c��P8p��Ns��^�`�S�t�u�A+'[�B�4�=�Mih���H1r��U�_{���q��ۀ�B�;P��\��>a%�@v�d��_�_ ^-�^�1܆���g[��%3X���P�h������x��
r���Rs��>�ؤ����k��dW��谊̋���J�.���-2
!��d�m3�c�%����8��W	��P��jЌf���;�������v`�N�&�(�Vn�2���P	�H�`\��|R�i�^��fR�-���_#�o4�~��j�C��y�У.��݀*�U��f�����eX�hY�t�6��\G���ߙXOE����X�췤�q)��p`\��;u�������w��}���1Л�T7���Nbƺn�4D�e�u!#q�6K�n7�:�3\��+آ6�!��U�r�,�rzݢ!�#O�ϕ:k@7毎U�[vѹ�@kiQ�<�N���J��"�	���m��%V���;��1��I���;s(*�2��π��aV��m'�� �i�K�kAȴ�����l�歟](�}(M�+�Z����C>�;WJK�%����1��L�g����s�����iVe͒� P�Jp�Ч5�k�>�&��Q�]\pl�v�]p�.����Ӱ��i�]βqӽa
<��8�|,W�|֞gZuu4��#��-��c��pG/V��3n�^��tќ���fe�D+j�d0���W/*�ycH>���[[�fWI/c7�j�P���o�.�+�n.�o�g�m�Za���;��ݷ�����I�Q�46#Ʒ���1�|k/�&J;a
<����CY����L��@�ӻ���t\7�ګl�"X�%;F��GH���+6��gl�Q�Յf�e1��DŪz��szX��7[<KN�؂��6�[ݜ��NA�㢕�y��}@ւ��H����w��O Q���Θ�^�
:�i̻x�1u;!�k%]mA�q��R��L�Sn:iʂ6,�;�cӜ��iTx�4����ʋ��z^�If��yRh�)=a�]d����W2�&�9܄�݄��P��҉�I+胏�󵊸��g�<V�H�η.�h؋��ʹ�̥�hmC_e�a����l�a�O��ր���Yv�8nС� ��8�A��7������g;�r�v��<�围��2h�VU�su�Bݶ�s$`����/�
#Β�S��Ǉ"F�c�2�u��{��f`�/:v;���7%%��9+�[е��~�wSF�Y��M�!A�a�/�^X6�,gt�È�8�96[�(��Y��*V�ѴB�x��sr���3�j���u�����.y?9>N��W�%(J$�K�I�M|�$����DY%@�x�D$��""D�%� ��"ZDf}��ZIv�K
:%���	P�HB�(�"ܾyr_�Eg��[�*J��_���9����^~Z3�Q;�B���4+��إrN�q5�iV��1��, ��]�dd�=4�GR���"��3��4���=�{�멖����2��婓csќ�����27�;��<͊�h��kޚ\��K�,'ͽ�q	��B�T+e��]t�A�����^+Sb"�8���S0��BF���@2�I��)�M5�Uv@�y���㝒�ch]_I��t��>ƥ�D��k��&d�d��+�}�y��KX��m݂ ��i�eaGK*�۩��䷚�㫡�PC���>˯q�,HyB͈q'7�ٗ�Iܯ^X�A���T��h$�$:�t�͔�Gw�c�[���C��;��M^"��v���q��|�~�k_][$X"�w!P�ZuERU`���B��{�+s��_�P�-��>���4�ˊ{U筤>$v�P�Ԭ2�y��u�I�-"�W��%i[Xzi�3ZA�]��sRt"�(F���옠��H��f�U���ì�eL���Tj�3HO�[הfr;�V�M�}��Q2�Bmqv�e,�D��V&���T���h�y�WU�Zm����ƪHzSr��Z:ה�"�w=�1S�\P���rƶ�r���<�q�람kv����Ŭ�r.�Oc�Ozduu���F�	� �of*!|d�vU��%�H�[�W���&W���{Xj��ni��}�G<D���V�62��i�W�$����uj�^�eL�OzM/2�q���f�qr�5馮�Dƶ���P�����p� ͒$��r�]{ٞ���n2RHZ�a]�i��.��*��=|�ܱ���]��Y^*�NS�k��Q_���מ��t�[�:�|
�T~!RD��W��}K��qy;�L5y��J./�$��t�y��w��mq��kU��y8�����T��
Ut.�Rs]oH�m���)��L�/*�*ܗ:e\f�<��w7��V�<u����y�V�W|�*�Mv��*ֹ���S˱����g~NN����z�bٺ�%��4����P�V��3NN� ��Aowq��A3�gdq¦�ʹj�MC` BHZ5j��ȫ@4�!�;��A�q��K��G;�V<�'n���8;�y��5:v��|tAL)�X��Wrj�)�a�a��X#§95������PX�������8���N�w�1���U�q���FN �i=n}u�=t���gb6��L���D�l]	��嫬vGj��kI'��3��vωsϲ�n���yL�<K�ďJG����v)�U�dm�8vxI�;z#�/N�^�kN=�Sn���8z[�_�?�Y���Jw�]�uz�Z�o����T�9���r��م�Y��[�Ϗy�	e>+��bp�XT�a�A�z��7��LE%zN���ݸp���u���}���t�s�I�����0��Wo���jg
�G]_[H��I��H(�I�DR�V��oQp#˙�?��K�S��o!��.J�՞*����߶��=WL		�Y$kά���I�ZK\�ݫ���T�=�Z�4oz�q��oF��������0p�Q��w~�~�<;=8����S�PPMYPAW%Z��3ؗ����0��[���Z��GW]A�g V�qb�nr��Τ��}��4t^����<���b1,q�ZJ7d��T(2�t�w�=��I.	�p�[��g��΋*�J*�!7]���oG�q�5��}��3Ԩ��t7����^o�[��-�s��ʽx肻�A�@a)$��)>�r��K"c]�w�w j�1�ݲ�=���Mc�Y��m�ԙ{�]�7>*�[̥�ͽ�q�CW"0�ЀhsN��-	�d$�zv�LGOPǊ�L�.�j�+;2艊뻃ο������F��APo�n�p�ˢ4q����Sβ�4�O��q�)�(Q�MX�B�Nϡ*5miۨ	�4ٛf\�Y�&����wæ�&�{���E�{��p����n� �4h�)��m�t���עI��oNf�ښ���ۣ5��1㽒�<�o;�C��W�E�>M^�j
cj[�������I ��$�~AXJ�/U��٩�
��6��(QcX�@�/&^��/ew�<��S��@o�f�ܧyy�z�6���K��${+/Y�r�7�V܃�V���/\=q׵���9��I/n�A�Ռ�߽�u��澜w��w�Έg皏q{˶�0��=��6��\�v��/��q��V�~GN���!�yH�&Z,'A��4�b�u=�y�1�y��G���r�5h�爱��;�"�!��N���?n_z��e��/M'���/*ɇn�Uv��E�݉�ӓiV��e��gW*y�s���x�p6��6�Cw�ew1����7k�wĞ�o���hw��mԕ��	��݋v����ui��{ˌ`������`�PV{�(;�]�G�k2��.̱�������]�"0�Uh�H�
J����K��>�qc��s���fIj~ԟ+��֫�>o�Hpr��t���y�]Y����g%z�D1I��
ESI��� �y��?8�L/ ��ā�}��V�����Hz7.o������77uCvqS��\�׻]�g�i��@�!��Y��Ȋ�y���Z����q�q�m�v��^�6���8���un�@e�{}�s1Mn��>�#W��,���������=�gh���r�I�����R��_�ٺ���EP 6�P���+ݹ�m@����&h�1?IC��#��n�����s�5�f'��ҝ�J�i����ne?�m2�d2XM�5�g'4�8`����^�\mq�(إV&x�{�i��0edYݾMk��Ni�O*�j%�X�n��ZvaG,�8�L�$W��^�$�}Z�p~t�u_���+ru�g#�N����zg�z��4x*(�4��/8e1�RV�5�.���lwtS�p�QRDv�z�U���� ��V�
�����w�Ⱥ��<nᖕ2)�M$)"�VP��W勽�v�U�ٯ��NN{�PqXkE=�M�>�R�m�W����ף�:����ʷ�9�(��Sd�p��S�Gg���n�6�Vɑ��yx��ݝ�<�i�s��S!��6�S����z�G��'ed'�+�s���F̽j����s���Ϛ�����ҁx���8�d�\Y\�EQ��M�Ň��^��-$�"le(��G��nT���o�߻ҡ�Wa����tK\���o���5ì�Uڝ��Ed�{��q��)3��u6_��5�~��t0Y��D�Ԥ��NH�
�aL��i�];
�y�s�b���Ӌ֒�Dةl����z,��mqu.��^���s�%��1-�w�L8,�t$g&�q8g�_Z;��&�1_��Wƚ)$XTi�φ#����<�n>5)�u�
�P�Rov(A�.U���4/sC�Ҽi;;/�Y�|UdLTB�kG�n*�s*С!kr����d�T�HP��,3\�[U�v�B����{�VD�����I.N�}��2�)P�ik�����Q�mr덷�D�Jc��K�Lq�<��I�sa�*;[�
/9�W�\����v�y[�������`��;qjq��h���{oC8�C\63S]�9���q�۲�]�C�ͻ�4��[��A���e!،�!q���o3�]	��k&m���]��!sg�����F���c���B�:��|�vz۶݄�q��E�<lE��u���Sok�h���v�]����4��ݱ��l\r^W�����pM�+�L�qfxծ���8�~��E?a����tm���d�t��+.�P9Q��qW��=|<�|�D����o̶�-��t�I�=�e!ǚ�+�p*K7h����y��|y.
���z��H^��ǞI��z�������ڡ~�B%��h�i����i&c�|&XX˽[떧�v���M�A�B��]I3�`x�z�Ie<�f�+f�t�4�P�$��KY�Xs>:p��vw�8�9��&�:�)�[�OL��9�b�B����=����+��I�}N�b^�|��z�|r�a���m1�{ �a����+��g��ӭ]�ȠȎ6:1�����KE>nf�}����Eҷج4�C伍���4Oʋ .X�U��L��vے
�s����`�W�]�c�M�[��*�H}��i�����g�����,hq�&Z�Q'��J�Ŷw��,���v�;㐡�ֻp��r/9j�m
��k���n��g��`R!�`u�M���[�v����\�L�L�/m�F��Y����;�St&�K��e:i�3�KX�󺷙���E�v̈́7w����q�>��|��N�}���|�y�9j����7|ܼ]�U�T�<��.E�ծ��肉�X
��jK��ǔ����O 8vo�z��VU�%����{��}0s�_R���:ݿ;�{�X5m�J������ج��$���w_W�����ʰtBc�2�ҳw-e�~�J�"��SnЦ��A�n�x���@���mf��̏Q�9�Pr˔��t)�BT<'���AD���\�qNι�W�f���Nt�^ì���
��3�[�rD��[Z�r'(-�պ
�vN.kM�7k�
�.TSE��sOj�"�4]0�S�6E{���./��}O�5�-#a(���_�<���q@�t��)����Z�h���������fv�9�ň��=��9U���9g�t�
 �&�.�HrM�3vG�[|���x[8�~��g���E�����d��ͦB$��$��u�<��y6�w�f��5VY�`��w0v���Qc��P��7Q
�I��ȳ5[���vvyJ=�&�k���[�F�qGO�D��(êu����ξ[QK鈨��[���O�*��p��X.�^ �s�Q�PL�:�M�v��e��lȬ|\>@���k��|Č>�|&W�W�c�=�~��������J�p��i���E@���l���e-P�0Ss������#ޮ���n�?-��"���=X��nt6_K><���J,U���}��K�O4)��}S������C>���M�j˽K��g綱����7>x�ûv\K��YX���P��n�
�^����rU��Sݽ�1f���(�c�3�9tV罥�䉵Z{]��ޒ�=^�U������"�E�OZ~"t�cn�V�כA
�����>�~u��Y��{u�L�gvL�K��$��fܨ�^�)�Vװ/��Ϧ蹶4*CA����"�'E�I�m�OWz.�y�.����1Y�0O�����x{�T��oM+]�t��*�t��@7u��1�f�A�Uv�����\�0ٵ��n��V��G9���Z^�:g�t��o��Da�=x�v����Uēb� �(��v�"unˤo
��pָ4�%:���jM.!qV�]���	3x�T�Ȧe�nCWR���뜾f����{kl��".��P�!Y�Eh�&�J�1���+�|����s��F���/m	�/y:E3�32�6v�ϼ�i�=Tu] �%$hn�·�ŗr�%͙�l��-����'L�lj��(`���5ś,��v�lp���KW~@?����:�݌H�{�n�Wa�2n	^�p�Υ]^У�S���r�)g�m�ߏm1�R���NY!j5=��	����~a�W�$�n������$�r�*�f���5J���ڨSw�`!-ps��%ө�ꞧ�O_ʅ�� Z���wrlz�c��ݔe�l��K�����ux}ҽ#��x�W�Y�/�ݜEQ����lب���y���q��&�N�Y����l)dn�,G�׫���_k�J�8R�b�U��
�{���S��n���X���O$iS�.��Ok�VPiQ��H�C)�x�Y��;���]"h����_<V0���b.ܮ�<u�x�猔�9����Ǯ�
�c%Ɇ��i��[+Un\�����A���wƺ�WE���V5θwn��B��/�O�\���P��U�!�au|-����r�1�le���3�F�o����5.�5�js�I=ڹeg*Z~=���l���7i���>��l�(���.�13��6D]�5}Wb���s����	6���Y:�:�d�k�Z��l%�+o$5��_X��q1����_X׀����&��c�E��K#�_�29F�z��N��`e�|���X��2.x��/DDA����%p,��F���]1����7�qc"G��h�SI�EÀ���X�o$�Sm��$��Dh���ے�ݼܖՑˁ�%�_r��<�O6H�e�� �z��1m��kj�3a���m�-�j�!��o������ӫ6��5���?f+k��]�@L�8i�z�Y5н��}�9wڞt�����{i[К"��y��Î��项�~�$W��O���4ָ�"۱]�[v�1�uc��jtO+j�N��3���Ջ�Q���]��/���ް�a�)����N������qQ��n����4���jnG�Z����X�C&�;2;;��-��*��v��P�)ӵ}J(끩�f7t�ˀ�ksW�� �3��HTK�/�����V���2�J�[Js�0.�Ʌ�6�y�3J�w]�YF�Q��[��
�K�,�s���W.˅\��n�Y=����Տ��cPYZ."���ࣶ���;�K�8�c�����.�a�hc��;9/����6Q���*�6�x�w�cy��c���v�`3���{�7�-U:�ϋ�D縓�u��p�r��q����v������gA�3��q��,��·����]��7Zp�Ղ��/Qۣ��3�Gm�[w;�}�oQ�s����8��� �{ tr������au"v���C㚘�l��y���/m�R.ے`��l�lv.ݯV��\��7n!�;[�H�ݵ{%��u>=s���Ǟ�2G�]�<�^�wg"����NEy�S�c�t�ݙv�W�7�bܻ�uu�uvY�=�3����=�GI]�yK����y�y�2cJ��1�a�8��j�Sp�fҎq�x�A�9�ŷ<�2gpWn����}���s��<,y�ywC�-v����poJ���n:;���Cӎ{<���]sZ�cG�؇�N9�zۗ��[��w���[����i�87Zz=�gSv�rl���Q��LKj��#м<q©<�������
���'8�`P��c���g[eǮع�#q���v���v��<��cu�g�j�d���ṡ������gv�GQ�z���V޷K��5��;v�pX���-�ѹ�T��x�s����-�8g�#�`:6`�X#v�snt"��3ݞ��6�<�hx��l��>M�hH�ιl\��;�oޛcf��a����kZ �v���7J=��^�7kJ�k���we�m;�,Fn��c(��
ㅳ��=��.���kFE0��C�n���N�ln. �	���7v�r1�c�u����|�x�x8n#��ڳ���\g(�^z:Sv,�nj��.�t��mK��4��q�u��(�Ӫ����L�:��l�����5��p Y��k�����G�/�=d㝻�3�%p�i�άds�	=���7�'n.7�di��x�,ģd4��э2��3��� �n�Ҳp���Ս�p��n�������0��e!�����b<�q����[��0\Gl���n7F�����-�9��ڭ
�CRkQ˗A�\��j���I�n1��x/#�L<8�D$l%��Q�˹g�7&HM=�T+�f!�z3�r�l�W�/9�\n��vH�)��K�����g��)��ŀ6��"l۴���b�`�E��q]����q�lq��n^�9���7�b���rK���租�S���	|��v�u�ʽc��$Z5\���;s<��ӻ\�p��:�[<jV�y͕qx3���
v�ycn�rkZ]ӻ�F���Y&�{�G�U�"����y�ğeA:NnsɅ׻�׈�Q�r�]�k����������,���c*2r�P�鰨�i�_�.���eϣއ�hyB�
��]N��2�w�N<�>x�{gl�M��z�=�z�<��nq�zPr2����z��M��鵶�>`*�>�m��y���F��M�{�q��+I�:�vԒ��-��9kJF���]�{]s�[1���%�u�+b�
W�a~w�J���~u�����3;<}AyǙ�S*Z�3�ũ˥�+A�~��j���wW�bz����r����&}z�����'�)��}�7|F�)�}Խ�|��I�d�[���~��yync0�6�� ��mn�u��u�6�ds�M��8P���N
B���8������E��m5�PT�k}ޕrK�W�+������>5R����Y��@��'�yj�P�h'Ղd%Zؙ�Jm���BDy��y[�B^['�i�cI�:L<n6T�O�wD�wZ���x3�jKS�I��p�*vs�7wYsM�"uЙ�:564��c<L��5����2aS�s�J��s�=V�%�eJ�j��?��d��E:��n�x��P�>����˼<T�/VNZ�5��c��i��G���g��k�{��۾�d�]��e�|�i�E6S��QDv���S�t�{E���aFa��9r�=���뼷Ҏ��a#>���E*<��T�d��h��b��x�b��[�'�o5@�E�#�&[-;��wWwrw^�V,*��ي��L��w;;r�]w���,�t�ӯ:��/#�JA�b:�^M��9�Y�I*Rr՞t�0p^�J����]���;qC�Av]���kr��wZ��ͭ[XԪ�K	H)I*�x���˓u���t}�ȥ�}Z�n��U�b� ��;�V.�2O'w�����T�^��%�sz�u'nɒ��r��bqQ�e%����E_�8�겾���DxW׽��D�n�)��Ϛ�ހ�ƻ����=2��u�g��,�{+�⧻'�^��L�H �@�Y��Q|��@�_��+��X��J� ��|�k�I��B5�xg�7b`v����`涒˧M�tLstK@�g]�X�D�sC�*� 4c���z@�i݄����+.:}�!3{k���-�`���d�/^!q���-h/Җ�|�ƽՊ�Z���y�s���v�F��^��I���6p6���H3���+}��eF^Q��Zݒ�"eH"��Fwsp��++�Ҏ�j���s=2��*=sؕ�!ѽx@9���G
�ơ;�Q�6�d�~�1g�&k����R���O���;84GHb�筷u�m�t� ����z���)��AR"]m��s�}{r��՝|%�(�d��z������ƾ�Y�]E#�vOua�/t��;L��Yo�C.�YB,,_���@�A�`����F����4��s�]mXF]�W{)��ǣQ���m?Ap�[��~we:][�y���-�<����~��4�`�f���"ԛS�gz���1�~ܱo��,�IS=Wrv����ܘ�Ty{�~M��U��va������uA[as1A��I��fM�$T�xJ~���ص�9)h��;�|��:�J���)O0ǚcm��&����7��4��o+.�5b�b
z��e�M��ݫ���'3�2�B�Ui/�`�7�K�����>���;���h7�����T��D�]�oc('{ɛ��S'�qr<5�Or��މ����6����i��a#	����9��^��΋wҎ����M��ƛ�)����&���z����x� *q��e#U�k]�s�����I��]���~��+�/!��ߒ��Y±j���={+p��,\���9���0��5�����ɯ�.ل�ZE��{����&� �������%L�����}yW��*���@�:Z���*a�?"��'��T���j�ԩ�:�wC="�um�"���>n�U���^�ګKo�n3-j��)'����T�Vz�-ח�@��D|[�~w-�9�;�׮�uys?s�a��]ũ6�$�),���ki��'m(���.JȂ��S
o�޳Y�G�6r�O2���{9�K��Kȹ�n�:�_{���%<>�^`���+��>L �iց����NC��e�Kk���Q���:�fD����YZc/r�5��g�m;�.M�k`]ޒ��f�����o�.ҵ��s2�qZ�ci��;��{��jީB�3*e�.�ƻ�LKQU���2��6ﰈve FB�h}*�L��˜���VQZ�
��h��r.<�{k�7N���QW��f���N�<qʧ'C`���8ș	S��:&� H#��L�V���:<g:��؜�)G�sq�䎻M��1���T\p1�����v�-����.�q�����G9f�&Y�.Y.�,U��篶�e�lMko=������L���	s��mv��k	���j�p��a�-�L0�<�e�`��\� WV6�5N\��q�p��2Zdfⵔ�Ϣ�F㕵V�-?~]q��9���������:�:T�=wsz.B���1*��U=��YNw\%�2y��'�ύ r�X����K�w����.�v�v���h{p���}�09byJ�x�|wjO���=z=��G����s��k9ud��Rg+xO
P��E�@e$۬�g�Og���$��NP�t�zɠ(/�:|ճO_m��4^�s�t�!�����$h�)V��|���Q�"���Kb�4���0g��p�}:uu���4{�B�;�	 �4���U��{;9��綏 r6��Kc�_R.J���ǰ��y:�倯���J�.�O[���{|�ԡg�Q !l\�=��w����﫭i`U�������/��ݍ�ߓR|��as!��M�d�g�jk,�щ�	�HFvC��Cu�lvݸ�g��/;��/k��M��Z��n�v�4C` �N�X�ٖ���#�������s5�qiNI�Gmd�����u��%I9�u8`%p/�&g����Q�,"��� �z�����˄�ܯ���7YO�/��r���a�~ݮy�֓#/4�l��\:`cߦ��}f�.'���5�PշM���c�1v�1!ނ�ح�����0��U�+�˩��s�"���o�uϯkx ���t��w�v����V��BE_ƈ"��/ \j��{G�{K�����F��묥�{u'n�m�Uy�g��k;�%>z�!V�M�TR�wV}۳�ew��٫��c(D�5��R�J��5!v,��U���{;�SC_��Ԏ��g��H��+=mᦍ?g��\�8gJ&7ޕbzճ7��b�.�:���Gns�� ���]%@	!"�|{8��[�M�G��Y7M*R�\����װ9�^^O�]�RYY�9������߳67C����݁_{&x"�&I�Y�0]].`=�OK`�\y�ܮ�u2Z�Ӳ�)J�a�f$2K@S�n�[W��wb�-�H�M��z�b>֛�G���v�av[Y�#�TRv}�gX�dSkͣ�U���P{�VÏXu�>&1Ya#@:B�o�:ʤ+�����O	��X�3�����1hܽ��[�#
7@�{�M�tu]�5>���S�yɶ��u��Ϗ������z{"����J�,��M��&���uէB�Il�컞����zd��;7����PU�/{{�i�ڶ�j-�MGb�lN�9�U�/��B�Qy�(p�I*�ˇb��AL.����+o�f8}.^��z�ޕyn0!����{�����n[R�w]�	"�ɒhXET�۽/ ��\���ek��^�~�OwR�R˲��!E��D��{=�ݛ���1$���=7:�;�jq2
�>���9�r�	��l��[�l0��9j�z�����h,X��Q����ۡ�����+�
��.�}y�r!R,���U����pb���h�N��_���P��r;�\��8�̅<�78N����񑽊퓈��r�n�g;��'K�-0p"�Մ6NÃ�R�)i�>u�+��U����(ڭ��^��砬�ꃅ����5��m���DV�c�0� �I h6������ah�=wo��'%�g�j@Ff��*�v��k�dT��$����(_�t]'�yz׈��8ͯy��c2=��t���\��e�i�M��^.�f��ڒ�LA
�r����N��z7zfK�C��ry���Bs�� ��u��z����ď��M ���N���Tv
�༧Ǯ>����ʻhr��vEP05:y�m\~n�����SV;H�������Z@�Y<��W��SُBզ�lCX`VIY�=�v�֧��s�n�����S�E;ZvH���gU^���9���z�~���uy��}�|>�{�	q�^��������X*�W�to�R��޾�����Ũ+��H\�����:�a@b�l��^�\נ(�w�i_W����Bs�7e�5M'/�A^nݟsG�G[��=�Sm\�h��kq;ٯn�XGGe��%WW��m�wGk��U��S/Y��T��{�>�*�b06:�!��e��&,OS�̙����sѝ��K�#^s�=���G�Kb��Ӷ��=G��D i.�u&Y �]��e!�=�g���W�)��d��]ۦ��!bw>;	U��hݭ�S֬}���Z�h����-Y�����h���_�3�'S����*{���<���oK���85�k˚�L
��X�K`���U���U;���a@�v$�) �5���uU�w9O6��)��k�С��z����>�Z�@:~V���T�������}�f��v��fZ�A��Ak�ek	Q��M���LKǡ�	��xS��>uu�[�B�<���4�F���ה�KT�zKv�w����3H�W��>���[���w�{���_w_��[��ٺE�ń�{9:�M�y��;�=۫�����xݽx�U�ܜ#y���b2��xU$d�AO{�г6���h��&����1ڋ��:˫spF��<�v�Xv�;rZΞ�������-�u��/m�n���hM`Gx��\i��g���N�{W&��V�c9��v���t���ˉ�=��g\�c��O��!�;{�ҹ{&:�vr����=�7s{YK����'�;	ǁ�ɣpf=����ژL�6���s�n�(�Yiٞ�sэ�ݰ����]-�����vϮ��<�:'n�B�i��7[��{<ᔫ�ܼ��:x��e��9F*Z���ʄ�h���w�V�DPv�7Z/ه���>"Q��;��=]m����.���D����V��y��\.밆2�$t�u����! �=����x�^�O���H��\�M@����{k�E��Q7����;������ ��}�Y�x���8�=
��"��f���w\�qf.D�%�T��j?vuԪٍ�sk3&���xzmͣ|4�7O�*U����]/|=���!b�,FB�ϩ(RB�*�PuL:���WWB*���@���y�,V��o���D���9[<�>8�>�/��}����/�R0��l�|o�y�V��c#�IV-3�f𞣼��$ką���xYl�vݿE��?9Rdu(n�T�ղN��p4�<
��s�:o���_36:y�c��^�@^{�����{�Uפ���=Gj1����J*�LV�7Uk��Iڮ�n���m���!J���LGq�©ǧ_{��t�AZ���#u���^:}r۰v�^O8,kx%0KYw��[��l�g^e����c��[i�L�7��ѓ~n�rͫ��e{λ!�����U�N.�G-��#_Z�8�:.�j�ݻ���Y��bn�kҬ֔8����4�ct�ԅx���N�^�xW
;tCQt�[������7��</_��dlr������Y�8���H�	a�i�Yy�<61V=�Sq���Z+��	����(��AWo؍W�Zs���}pS��	鞲����c�=��i��Ə#|N����al���T-g���{��|w�˒���!V�*M*�/z����<Ӽ��7�]ƍ��.��.��mO�Nj1�u����0�'A�KN�d^��oo��	X�,R�tJ=�Oxc�ג8�m? ;��$}v,�]Ӳ�C��-,X�*
�zW��Ab��q1LV��w7&e��)��s���xw8�s����/lv���m�.��t����#ں�]ֵ�v��l��#X���ʚ*���@Bj.���
ny�Ҋ�EJ��u�F<Ǖp�Vj�D&���X5�>���Nw�^A�O�k�9j�l�2	���LZ�S��O �,C늓5�����	p����d��ۦH���ɕ�뇇S�գ�՘F�5>3;�숖��"�����xSti����o)"9��zg*a�O�Gǩy���j��,>u�l}3fő[p��˙)l��og0:�:,ά�8ǖH�Z�7������ĲE|���J�����t��%ui�v��n������gK�L')��vnق�!�����M7�.j>z6�#Y{��n����Pb�t¼��Z��J����o5?/�d�b��>�O;rm����ފ㕆U���^�5��6j;[��q6��r�rm�>4�����5YҟwC���N<Ԛ����O��j���l�����R����$o��8���N��(��]`��9����v�z��!n�_t��YQ����c����]I�̦+�1�0�޲G!c�c�&�=��g�7������[{�S��갢�M8�@KhnV���ۓ�ȹ��ܦ{��Q�~9�F�Z�ġ�Fev�(EG��,X�j-Z�2��s�I���*ܨ����s'��������j�gN��'�eu��W��@�%,x��L�F4$%챮�<�{�MJ7�Na�m �b�a� 60:�QЬ?C�>�b�����G�nVG#D.;vuqh/�7[/�+F����ۗ�>�&���Z]��mG8�}���x�.(n;�%&�G���m/�!}�b4����]mjnpa����W���=C���6#������GzF�ӪW+Mj9��U���܋'�K&��]"ό�˰`E�d���l�;c�����kc62���u*���S���s�>5vGm��r�֋R�Z e��ݭvzܭ8���<�/���Mx��R����F?a253�q��*�C޽��#��j-s��3�5c�B�-�Mٿn��]��N�W$��{��J�z���b���z۫����.W=�u�VX�gǯ�U���\���V-�c�I�"�L��dV*��	���k�:�λt#Z)�[Dq �o�i�6�ӟ\�%��ה�������?Y������b�~X��yU�"���Y��d�bE�(�=�q�]�j�v��vJ��3�{e�q�{On��1� f� յI$�"�+���'g�z��{ٴUӆ���@PT��lw��OqB�;�c ��<r����U�(�pmP`�aK,銴[��{H���JɲU��>th�2%���I��p<c�ۘ����Aԁ�d3���z� �Mbd�޺1ٯF�h�f9���B��A��DJƶ������X�x`�����D��7��)���s��>"cA�>{����ζ�X���V�bv
��we`�]r4��c�~�Tݾ3�Һ�94y�<�-��䤠M�(R�*�s^��$�룖6*�Ԡ����Ƕ���3�֖����jy�OY��B�K{n�k�6��>�껩�Nĺ��˚(�Y�`�(wL�6�#���V���(�ה:7��+��Lp�e��݌^�(
�� �{�)\�wXodחcHh��a����P�����X)�ľ��{��o���
b��Kܬ���L��i�NU�HG�^��r0�C|����ʨ�f�bTYq��Iŝ^s����!t1|�@ߓ����kGY�����1r&�ruՍ8Ns۴ݮ�flD%dN֥#�n�U學�G%Uk�e_ل�Ώ��+����9;pl��D~�r�*��gT�fz�x�Y����f��O�W�wc�h��`�7<�+S,
�e�>ӽ�n�_��ý�󓷷-$}R�Q,�ˢ+~��g��B�$��!�;{*�F��x�p�*S�D���<�������yj(�i����hu�״*�9(��fp�1��1v�Awܻ~���Gw���q
�V�_�<�Y���*������<=�\��s¦�^m��6�##	+�;��)}s�^9�����{7ݕ>���}H*��o^T���:_9B��K�����U�5��7�N��l*���;)�5Əo*��h�yqh僪Ғ�H�)���E<��O��`�G��T�;�2nߨt���6e�ƽ�]o*�6�P�_o��{UB&�}���(X��]J'\�u�c�ҳU	YjEO+u�JT���{[��[�v�eV�լN|e�3�aʊ_f�!�S/w�[�&�l[D���)$Y�0��mum҄V��h�v�8��f��3;nn���^ں���lr�z���m�m�Dެ��8��ݳ��K�v��H��2"�W[kG�RZ�3/e͹���O`���۰���P���kh�{���׷##��n�;ݺ���K��;u�mu��۾��!�m�]�GϦ�u�nri�b'`��E ����cW6x�Op�8���o/=�ֹzV�4�غ�s<U�}���x��X
�ۉ�T�-PVI��i絽ǥ��<�G��S߷ɽh}c�aL�󧂦�UL5�jL]��̡I�u9���*�� ^��%I�i�*?nRF���v��d�������P�.��	%I��:��ﳻ�"|�3/�X�601����7㏼��f�>��)�g���S��p}AOu(u���֫U!W8=��Z) Yl )�z�B�=�_�~B)�S�g�vM����y@�_U�����Ǿx�t������/��ީ�h `o�/�]���>ړ� '\��_m��r]��s&�js�ՋۢU������<��&��_g�.�㯳@�Zr��n��[���A���x��Z8_��	9(���k��o��TVK�o�c�U�]�t^�H�S��G-a_l���q\,!�e�B�{Ϧ�O�dICaVkE:�euҭ؟�P���C�.��'J+��M��Wg�����M�==�.�C9�'��`�\��G�}�f<D,��e�iu�tLUI��>gRt���dr�{2��;O�X��z�ᴵ	���y�L�+�(U���8"��5��TM�j�k�q�L�1N�t��aIUolDa&;b�s�M����@�S�
9��\�9�TW�Be�G_Z�$1^т#\k3O��Xӹz}U+�-����VwRDA�tĂ�%9B�NsoϧB�fٳ��<�l�N�;�k��*,��R��[��Z?ck�'	���ĳ[���$�7�;��נ�`���.�"���W:pK��0w�c���n��E`6H���$4��$��[o�]�)ͨ���w�*|3�L�v�+��C2J"���}V>��V0�}��i|�c�����α�����X��B�P������ܶV�	[�%4��BZ����~=.�b�[1�/�6�3�r�\w��IU^Ā��P.�9�.�X�.��I�]���^Ej�2$���; �������{��\�;.���a�j������
�Gc���m�1�>5S�<5^�b��S�^AV+��nx0y,J>Ő��&U^�����.d��7�� Q� r�Բ���W��{��48N8'K)�6��L.Ifs��P�OwU�/���)3�"���۩-J��h�^�����ʞ�J�zj��^��]r�*@%f�y�B
v�ع�n���Mº�В�9X��=f�4��g��X,$�D�]<���>�� ���5����읚*�8�fy7<���n��:9�җ3�N����V6"o�`�8�s��R��md�&j�U���Mqq��w.��=ݩ^Z�f��1so��KS����'�/Gx���i�M����@�T�`}D镶�,�7�n����/h�UhyL�X3�J�+��7I�p����k,�tj�"�k��]0�.��m�����W3���\Z��h]ZI*�1�
�L'ޟc8j��
>a�'���'~�[�_	��܏�G�/K�\}G�=?XX~a�����Z�l�7�Q,R<����V��������*����Ntf�86/l歍Yyٛ��`6���W?�?�<�����l�T5�/��>�u��i�7qP�*��eA���q�Ď��k��<�z��5��U��hR�����]�+`*B�i�u��K���7V��G��(ѧ�0�t5�N7Vq֊#9\o�o�ѥ��p�B�X�G�p�m���~��t]���n��*��c�u����"t)f��}4�&s*��q�Ʈ���E�vC��X��t0���]�S�L|����h�<�R.�ᗗ�f#^��јET@m�tR�����L�	��A��������Djes<�-�`�C-�۫'՚�����g�ڞ�a�{�U�NNX�|�g���T�=��y�|�By<��.�ژ�ߍ�4	�A
Yw�7)����6�$��*���8ٶ�Rݥ ��[���y3#nY$�mց�I�K����(RX��:����b�"���@�|��rZ���D�;6�AD�]澘��z��]����wK�(��LWCc�F���`�|}k�5$�Խ}9�p�J�O<E�+�ɎܲVp=t�t�Lvz��u���b�%�t�vy�n7Σ2��\�?���*�E@�m>��׺zV}��N��rҪ���J���{�+1�['ʯ=*yG*.�a۩U?;�����]`�dk�ƽ������eb�f���rڳ���5�ή�9����+���o�S��0U�;u+ 
�F�P���X 
&N��~��.��~�
u�:-����_�'����a+Kj��r!�Zm�:��~N�*U�CW�eM`�¯�.�#ԟcգU����W���+�ب�\�*R�wJ`�����\,��i֎��tr3������%�L��/L���}O<d�^���n�i��==�ڞg�cQ�1���X>�Ɩ������9S`��.���^=XH�٤�-��^�~�d��]*���I\qU�;���S��?WU�> �4�:ܠ�!YʃU���f��S�0uր*�T�&��h���Q]���v�ݣJ�e�&��ɦ�����R��t���q�����!��;�%V�ֺf��;��Qa�x22�F>}M��k�0�A�/V�qr��x.s�IPni�	o���t�����s]����nu��>[;z�&���6r�C�۳���O�k#�U�Cc��cny��;�Xn97v�u�}�ݹ�P�Cg��C��u��4k�r��9��g ���v�p��9��.����X�fyP��M������ۓ�8�*6�:^��@UF�O���\ɉƛhn2v�.�gc]c�2�ǵ��{U�7fcx����<�F̒�6������z5�Q��]����F�.+{�w�0K&�n���!���t^?�����چ�����a��'���&���O��v�5�?X�B���N��V�L}[��Z��nw�������H��Jϸ�ӽ�[j�K��U��
�{�X�p�>�J����*Y��% �R$�Hk��ʕb��C�����b7�suE\b���,h+.����Ό5[61���~NCBX���]�;|��{�n��YP�V$&��O�ܖ��2�2����J/M��]g
L:tK�>�K9�᭱+��Ȱ� �eE���Մy�D5�ڷ`����jQh�r��ѩgD��^����H�v�h�i��:��u��q@h�������Թ=��0��D>e�:��qW �Y߻�_�����WY�?z��05n~ᨐ���t���\�S�w���v�˞�zn��N�$v����]eF��9�z��y�os���W,M�aG�}n����Xuh��O�؃�C
v�<U��WZ91ۋcD�����O���.\���Y�ޕ1������������V�v}��%�yG�񋓨���ӳR�|DyW|���MRÌ�`�h�)���m�_ˍ1Z����S4p�z�i�%Ŷ�n�f;9�y�j��T����) �y%�A��^Q�Tz��	��]5[z*f�*�肺p��21��
���Ɇ��V��9ma�v6����γ4E�YG׆��9N����7"�ֶ+���{��';e�q#J�+������|*�"����s�]a4l�G#T��Q��&��,��Fڣ}[��S�]:�0��_1+-��W��h�ۡ*�H��}�"vf��
 �)����轥�/��rOP V�ɽKpI��xSh�c�MR��!
W�ZXTi�s�P��k�C��uk{���^c4����J�CY�\���ܕ�Z�����K{�T�#�Q+�}ɥq�A&X�I&��ʜ��Ͷ��mk
����֍
�v:�]Vk�?���0o\����d�ӯ`4G���_'v(�7�POr�&�%R?#F���e��	]/2Vx�۳����b�3p�n|�{��,�jT5*mY*���י��+�-Y��)���Ɣ��7W���^>^4k��!�[����_qhk}r�oj!�����D-}vT���5�&�bb��mmE�FV�K$�1�湌�ωOgV�pG�{إ۴�������L=�K��J�/R��4�ٛ���mE��>t���w���o�>F�W�|G۵��U��A��6�����Y��(���R�S�0�5����돕E�̷���|r5϶�${j!��^��)HF��"�ǝ/Mܔ�s�ˋ���I�1gn�1�C�vX��B_j���%�j����Z^��x�^㢯�G�2>����o)V+5d�����/6E�X�J5%��i?�Ͳu��G�Bq�J��Z�TG�!^)
������aJb�k���l�V���e�^��t=��s/U��]b���nj~8��Cw��I�)|KM?��t�5��M}s���	6t�U���g�&|��
�ͨ�َ��3��� ���{�4U��|h�鳾� c�
h2����mI;׭�jymD��#����<�w5z27���f��&+��ʦ�g�c�{.*�lP�U]#��-?}��5��e�E���ԫ�Yо">����c�F7w�9�"��R�f��+\&�4�x�Sۻ��y��}Z�)�ؤ*�V+�*�߹z	2X�@GV�nM^V�~����֝f��˺ez=�(��,R 7.�ADеDn4̚�]�WY���^���s���+���}���
ܵL}�v4�a�J���
��krpr�
B��&˃`:2���x��T�D,�z��BFp�up�N+�h'o�V*4���{)��1�8g�?LGʅ�65~�,��m�p�w�a�D��6�g���uS`3�7�pUШ��s(
���+�"�`���g�N�A��T��/�F�).D#��ٲ�Gk- '��KO;���gH�{�}wS���J�{3.�ry2��nν��w�qjk�N�>B�h���'˽jȯfΥ}ӭW���-��q�d޽�K��X���;RO�Ԩ����ˑ�5F���P�3�p��W\+sYO3GL�L�7�+MIb�)P�ʊ�.�&[u(�dʴ^���Cg3��:�ٗ����z{gsuoB��AJ
�
�dRϟ����7�e[��q��g�#npF��N��q<�ҥ�k�1�v�6:]`@�Y弫���
��]M���i��
��k3W�~5�g�ۮ��[N@���U��x/�*wZ�
�ɫ�����qE��k�+A,�s��S���v��`��D���Q�Mp�哳��D|񅞿C>��ކ����Z�=�h��k5�{$�sB�T��7�(�
����Y�,�`�i
!��b�?Z0�v,[$P��sh��Eޔ�&���|%C��4���e����҇��U��U���J�r�u����I��@@qV{.����Z(^Ֆ�L�(������y�{�m]D����ƫ��{��B{=邓c_�,�*�T���ԝ|���T^�GⶳÂ��2���3��oIY�����d	����°��妇��f�n܇9�p�{�#i�1'Q�3�t�ۿ[�^�ѭ��,J��[{�y{�f �5��@CCe��>�ѻS�Xd�QK��� ���
�t�E�s(��_t`�C�7.p�,�*�v��S��؄�"fn;��P�7��JDl�Yۑ	զ�5�9H�A�G���nUK7X��/خ۷��_�yy��MC�J��ʮ��٭x�*��r�4� �u��}�5I�Bǈ�+U����ՈM����P���͛L�fړ���s�S�5�7&���J�04NGf��\Ē�K�'&Yn�OeIB�;r�R9���\W%��b���Yc��ӻN����$�M-�e�1��RZ��t�$��b���F�u���m�u�I+��K����������܉M�q�y��z��F��L�=GN�Ɨt���lT�Nu{+^�:�'B�- ��J��W��BB�D޹׳C}J�X�f�%v�#s;!��3]�w�,u�VI�i�t�+��,֊G4���i�r�,��T'e�9O�w&G�IF�ԛu��qغYn�I���>���ث�Å��\Z�������:�����D}�Hv��j؆ܼ9�Ý�ËvH&��|eB�!ul%v��]�9���&�u�,K5Ч9�K���3���s
c��8q��\�]!���ۖ�@<!�4帮M襾�y+^f�t��r��{�:��1�|;�RW[�G�Bt��������Z��U�r��I�!����l��bKj��Ǖr�q�]ckn�x�>v.^0�}|p�G�m��WU��XD-��r{{Y��Z�V꾠��#��C6����F�N.w�ۀ�@'D[��>��+�Wn� p!���}�s�ר��I�XI݆k9���P�<G��pA�TN9e�Lfs���f�Ƒ�3��Z�/R[lN����m[�6�-�r^{<�W)���v�q�;g��`�y��;6����k�x4wZ��N�@+�W7H]�q�\�3�g�GZ"�Љd	F}Tbd�P���^C[��#���E=N8���׎�>v����ӻa���۱�ے�]�Pm�͹6�:M۹��y�ݸ�m�Kۺ7G=7t>�,���2s�˳������4gb^�����.N��{d�[s
c�ɼ����������6-s )�v�0v��:�q콷�۞]��p��r*CJ덞"� m��ۍ��Idq��]k��{/Z��I�ٟ�^L-��l�d7:8C��˺�p �ݱk�a8;������n��7��%����/'
�s�X��kX�]u�7=�ݩ�[��+�L�;\��s�:�M��#mi�W;���W���\Fs٧pk�ki.D�D83O'���qu��OS<n73�s�֠�=��.t�ݻ]��M�'<�	p�Vy�{u�yz�S���8'#�����k��W1���y�gst.ː!��8��9G�d��v6�wk:ڹ�h���c;�Ş�����2s���ҳDp���ݵ�c
�Y���ݧ������\�
�n+y�ms��.����r�G�
�]6v.nKcS�<kn�G<�qu�)�3��q[�����7]�{r��%�Gd3�������q��p����63���xL�ts��1�vm�r9�[���C;ϵ���:��zJ�,4-�N��^�v��N��]��񞫱�:��1��Ne孶|e]����5�q��ͯY�]�wN���<C�ݷjy�]��8��zE���nG	v�v=S�Jѝ��=��/nm�|v͹��b]��Xo@�6T:Z�[XX���@@Ь�j�"Ұ�	H�'æa�l��N;&Yt��7t�;�O���Z�v�#�"��i�K6�v_�q�Cۘ5u�ݝ�YJN�s�w:���Aa�Q�:�,ca������[����,�l�O
�AZ�wnuշ�&yhO#<���v��S��]�z�Z㇇�����lv���(���rC��!pԖ;pV�z����i��Ì�m�^��Y���qpgg=o�ȴhx9��x���;;��6�;w��m�6�y��v�szX�綖�rk�m̓���\�v�M��I���]q�F�p�d�3*?�z�J@���S��U��q�n�b�f�R�)��3�ִφ�{c>�DSe/�5c���yN��_e�ƛW^֬c���F��-z[M&�U�/����<�+A�h�����/E����iC��/]AXץ?(�,m�7
k�x:X���F�Ō!󃧃!P5E�I2���{-AT�A�]1H���E�^1S�P�P�*��{k0ZYɁ���<�%��S�����bz��`m����̫�jߓ	�����14�e*���myZ��[�7�<W�}�4�O�焫�x��;�1V{��ݱ�/�4�ǔ�j񕞋�ˡ����x�^�v��y�W@}�P[Z�=#���V��յ��R�[�L���FW�m�~o�銒'՗���ڝ-[�n��
q~[�X��(
���u��~´| ��5�{�c�a�ˎ{�������,���pY�e ���ֳ��o٪C������\��l��k�a�:e�{`b�0}L}7���ove����%H �������Xj�,����c}���~�X��AD`�0q�U.��fl�ĂmKMMk����"q�K)�91g���<��'��;�}Qi�L^�v��$����-�͡E]�sV��͊�w6�ӏ�%��U�k6N���%���Hɒ�vXL��M�n��RN*�3���v�>�EB��=u�5�V|q�.u��©�Ymj���yf�Jp�W��'��j��%6���yQ�4*�������{,�q�ml^��Ub�1^��'H����8pڵ<_^p4'6Y�J�x���TG��P9��֫��*�D��vե����vH,ܭ�;��g?Q>�7=���C���J�J���l{����s(q��w�����V��<k]F\��8����L��M�<���*� Je  �ٟU�TE@���{>/��{*[��m��н���CO�y%�rv��g\��=z�S�dXn�"��nr܏���յ���s[�hF���TJ��W�A@�=�u�Bq	�/:��]i�.�Mע�u���e��%t_V��ns4�O��o��˙��N�Z�Z��R���Ay]�Տ��Zj��A�η��S�ל��{X}c����E���M�ĳѾ
��q�d���ˡ�يiț��\',u�bz���dp�ź8@�:�a���/=�(�^���z^Efi
S�+UA�������,���qD��(
_*H�YL@D{/&�s�[�<*hܬeS��3�-�����jޮ���g����+�]Ecn��Yt�u7��hm�:�an�f��̊_B��ݭ��	\��fbx��>u!��=�'��7et�o�tfb�C+u����N��g_����[eE��كӃ���ǖA7�m��u�
�)�c�n۾�O�|D��J�B����E�9f
^��T��ݝRH]}+>���ՖTӪ�Zio��WbXڃ�N���5�����<�ᖇ3%+��J����25�ms��uCA���>����.�x���m���g�h��ݔ
_u��[�x)��SŜk6흖��u�;3��B��TNz����o<�YZ����w�������3�/��>j]B�=5ԹirU�e�Nd�/{���n�:�00_�[���;�-֎c���}>{��(E+q��W���R1-S�v� �WXuG�[;�s�_}Z�g�h��C˥�D-4��ҥ^��8�<�(��E�a@��6��d��'�}d�[i�6Uq�Og��i�AY\�E�>5���_y�N=��S��pOo^����S��|*^?N=XX,޲s�J�<�c�a�DI��і��G����έ���p�W��T��x����Tq�V�%�Ox޶(�\+J�M���4�֘��7�'���D���(�i���]�*���t�z�$���D���ګ�u�sn�Dy���w��I���ܦ����xzJ2��jـ˶:[U'�nU1���B�f��%M>��KT-	l�=��x\�rGUb��'���n=�i_���a�w{Ӫ�*e_y������N�!�}�R�>��(6�s7����뻹�r��tC��0F��;tݷK<���[����6W��S�ɽz�ۄ}*n�l�r�A�KLZ����:��r�wDTF�:�>��,3�Lp�b�����V���j.��u7�ā�s���E@��vYr�07��(��UKlޚ�(���x7�W��M}�u��8��¦��z>A��yg�X���������)�ma���2_��~�5�7��y���ih5�`��I����#�Ro��M���S;<���AU�lHM����J��u+e�N'	���Hk,}��ׅT��S�u����S����E�Z��*Y-O�}��x�E�!����S2{{�S�nj�Q<L�8�Mxk�[��e�,�.�Uj�lH�2_R�����=��s���冗(!Z��!LJ�xh֘+I�Kw�c�v�!XeӪC�9�l[���|��1������[����"��棛���V.���}�<�?a��B�?Ui�����v��^���Y5v�VQ��R���.��@�N�aӖp��qP�lHͷ�w1n��]2���̫���emI(�s���A��sn��u��-/n����r���-��;@���cǍtc��<�5�DS5���[���xg�*ewn7F-˓�ݏF������2��{k6��=Xq�.wwG��vٸ�6�E*;�/�6�6:2�]n�hܔY�Ot[��ۆ�Zݭ�p;���۝�^v�9�·[�YNͱ����s1-�m�f��jMm�;s�nl�Ǜ8I���S����� ���I�b;v��.9v�[v�3n{1.օf�ҵ�ۛ���SfgPY�Ҫ�g���;�WT�8Y����"#J������Z�@(��Y����PU��"�dpQ%
z�^�R��I���M}��C?V��T*n�f�士��"�9�u�d�@����k�S���*�����;'\mf��[�c�i�Y�C�n�j�i6B	�uxi�Yh�*�R��ҥ�%^�G�Z�YO�Պ諾MU�P�$0v���Ij!Z�,\����RBv���"Q	3�;�O�544z�{�gβBu����z�ܥ�>�1��/��ݧE?{�S޻޺�Wk,|�n][����;A�$!U�I :U3T]��ھ9C7>ϋ�M!H�\�X�#S�%{�Ym��#���}�S	��0 �>���ϚQr�@���7�����f���D��!�����秞�/��V}!̼/]�q���������ٻLBQ�2V1HIl����Y�ܫW{?rj�߯���#���%�[�P��M��O�6(ui��R$hq?{�Dz�q+��}I��F(�VYK������b���z��|z{�.4��GD������ك|*RV�%��8�&�.��%�K���gq��O�b�X��Fi�����ǫ�Y�}�n>|1r��4�
�R?,��ܙ���3ڶ����u�W�W���({K�T�Q�E"�6�$���t�M^sU�<33�9`�e���c��Ǜ��	�]uh��<M�}���zF>@�*����_�w*��LljK�v�u�S��tP ��Q�����"��,-�J��ޝ�2YL���G[�]k�z��5wQl^]9?B�J�����3!W�s�a�Ӡ�}�~���AK+,�kl蛓���Y�un�;��	`������f���3��!^ X�� %��m=�Š�<��NG�S�w�P
J��׸c=�mo��meת�,U�85U��F)}uk��k��ڄ��vg��k-��0�ݦ �"�8^d���!5M����c�~*���/�����M1r������	>�� gu����4M���i+���TD��4���Es�	l$)Re�0O{{,�h�`�Q�q�6	�)n�����얻\�Xy�YB�͙�`�+�V�U�B��AM�@'���֊��nT)�|�����>*���G�>����l�{E:��<d���^l�va��\���ue�hTe�U�Ȍͩ��<�.uJ�n'o�UfԹY�]?�Й+���j���"b��V���m��.�ٍVży�7\,
���w�cS����7��b=�>-�1B��2�ݷ7��VH��X�&׈+�ې�С�</R�h*N%��AX:<�Ϊ��v�,hQՎ�S�9�c���6ӭ�Y#�<��U���dRڵ����q켩!�%;�tU�,R�W뭦ree|�u]na
���qb2J����v���{p���jbT(�i������ֳF�Ʉ�l��c�����R˩!�L��!�]���9; d�I�Sl�Q۞� ��-����~����Rɞt}��H;uN���c�z�c��)���������:�m�<u�巕��j[��[PGţhC�Ti-e�\�=�wc���嘉>W�U�~Ý�iQ%��YS"c'A��GY��]{T���f�M_5ܭ4ߎi�)J�(����z�9Z����m������,3s�w���+<i����Y��=�*.�E�cC7��A�^Cw}�UQg7���j�R�SQ�9�BWeo����ժ��ܲ�K�٭��J`*҆��E�c�9������R�c����o�[� F
z����[e���4m�[�<���>�O���W������;8)ؠ���6�NAWW&Y��*vwʶ7l�ђ���iv�^���֏����̡G�[w��M���=���|��iwW��җ!S�B�j�go;�=o�۲AI�g��w;�ÒtG�c߳��o��.��P�����v�X i݉9���lu�h]������J�C�������|��J��BU�\"����"_��֭,Ք�@������8dj��۝�I��sz�ˢ����X`̮��e:a��i7MA%$[}y&�f]g�:�ʻ��D\=(�;R}k��}9^�l2%�uIR�7ƪU�v�{��������,�&�֏q��7�̳L�E�)0����A�+טm�́��B��[��J�ʡF^����-3.�e��r*���~0g[n����myV�PM���r�9[��HIM���3�R=:!7���v����}���������>�W�k4�u��3�g��4G
 gWq&�R�)B�t�-����>/:��n�u���c�=�>�4i�{3�P��Y��t�7}ð�������]�<��Vc��$`�]���Ԇ�\}�/��(\r3=�c8�췯��죰3�ԧ��b�]�f�է�N�e������ұʺYΨ��u�)&!�ӡ]��4i��V����x!���a*}Wݡ%X�^	{� *ʰQK�V;u�����ˍ`��h�&��=����-��3\@�8�޷[��/.�N^8|��Nx�;�ѱ����=�#n0=��m���|��'[�t�2�oJ�n^#b�n���xrD�]�ì�ɻ���*� s: ۩M�����{+�\v5�aq�����=��,kn�W��%F*�O��:Lq�8���q�v��k�}Eg͜�V�Y���F6KcM�Lspּ�x˝חs�=A�iPm�M����$���n�����TDn�[+_	������M
���e�^�Bޗ9��_v&nFnӄ���zt��(m��j�8J�)-�"]����x���O+�����O�� ��)�л�ķ�I��)V��]j�1^d"����^־�w��q�Ʀ�E�Ӽ�|�O�Q@$��� �j�O�+lW��ϕ�n�w��κ
z�q7gS *;���c��ڂ�'[�B�_���6��F �`��'��$�l��D��x�kӳ����X�YB��wcz�V&�\?H���e#���_q����3�XZ�.�J��<�#�G��&��,V8XKZ����*�]�d��]϶��Mo�*d�&�|�au��,���ʭ�f�n��.�a��-t�N`�����Y���-Z+���k��{�L��5�5�D�Xǎ6� ��ͮq׳�p�5�4s��=1��7Þ_�{eV[�E�����fc?g�J�#~�a���1b��*;a���Q�u��dF{��-o�%�K�3���n��>�S�*�X�?[@"lq�V��8C/�z����ق���b�Q�d>f�V�eOյt�v=:Ң�-�o b3L�׺*��,tvqy�����ڷF�:�c�I�l��+".g���a�ʵw�O�I "	?o1�_
`r�z@�x���ִ���e\�F�bm:)5�4� [ǅ笌���v&;��e{,�5l�{��`�Z�9�y,�#���r�sjf�LTew���-���KU,t�z^�z[$a��:K�Yq�q=��Z4{�z�nS���r�}��"���.H>��"�u��O��i�����|��Ө׫���IӪ����r6ѽ-kZ��F��/>�8n`��s���Mz7��}U����ߗ��3���~��{�qʱP{bY�K��%��oz���.Q�J�2Ȫ>0u�:�f4Q�Ѷ�;]���S�b�=I[�;7�S����%m���]�\����o}=���{�k38F)��)+���*P��^��b��
�Zf�n�T��eۨ6��q����T�f>9��q(鷺t���i��j��%5}јg_:��@a�!��7ϧ��^���@R{�[����]O�,��^V�+�S-�A0���r�Jcmݬ��hg�{�1e>7�&�گ�Хo�aܨ�x��2r҅�������ėà�Ajy23][S����.�n�ϫ⢐l6��=�$��G��\5A���g�x�r�t����]�sL��E��D����V�N�D��X�!)sԆGug�c}L��y9�7�����z�li�(]�j�Ж�,��65��Ǉ»A2�-&~1�W;N�a_7V�ubı�Q��d��3�g��j���z�4��h�o&B�42��e�.X��yo��,^�y�Aa�[HS�`%��v�<�D�Ev~�
^��P�Q��> �L�u�y��3�	��45�r��*(�M��_f�i�B�ܩ²VC��l��R���y��g$�U�ykQ��pk�#
IS��}̬&E����kW�u6%��{�(*^��:��2r�u�9�쾆�Z�IY�vTȉɵ��@}����*9��ҧ4��@���ol���P8�"�*�C����q]����*�#��+1Znfj���94���G�].�$Q,�"����=���v��r>p�b=�hlf��Q��*���kG�k���ڜ��I�1�!�gg]c�N��X{8^hg=ȵs[�Py����v�ӱ0T�}�ζ�w�s�Z��X�#�mQ�4��t4V�&K��R�w^|y��[Ϣ���˛P�z/�tvRӍg�������e���|T:&#xU.�uX�l�J=�j�u�B��a����KG�txֻ[d�X6��T���j4���U��M�^��F��D_���ޕ��Zŝny��J$���K�Wh��lK7�����}�ժ����zk8�P��ja��=�^o�}��o���n�V�D/���z����-�c�?l�>�1R��B4@U��n��`H�:%=�s��r�g(׽=��ԣ�#�����>ʳXj�U�~<�ႼjCZ��������Zmvz2�F��uZ7*r�Iz�.8�lgX�xv��3v��v.Ïka��"� 6�똃��J��>�y��n�ζ�T�u��I�9�BJs��Jүr���{G\˭x�*K�.dл��ŉ���\^�D�rA��8/�V���~u*��oN�>�ƈ=��\��3v�z�?>�r�M�t�W�������~=���g_�+�^֋�7׻;�Ae+(���+�W�v�Sף�n�.��2�<jN?[5�H]\�N�ݣ�`iV��췩�[�`�&�+�ݴ�e!��MR!%�&��L�r�9�,�����9�ޚ���,y�����z��]ka�}/|����tn�rt�����P�^/R��r�W��+[�j��-v�jޮ���� �n���c}���]�h��N�u:X�K��;����w��z��1�y+�{�F����Z�5i̬
�|XDN�a�sڹ��,�"�����%�M�L˰rub׏s�w�5��7R_�^}w���%�=�-�XKn(G� lS��:�N.�Z9H�R�Uh@�6�U��;!��S���q<[����+C�φFT�T1@���?�y���+�_�+�}�ޓ.�	"�&b�}��-ԡKn�\iB�';^�M����n�,<��Nx�t�^v%�d�v�A4�T7��[$�"x%���ڷw�%�[�&x�9GҰ��hx,�u!@o���+���RD�@�]羳�f����~ � ��)&S��[�֎��rf��'`�X�z�X�u��:�S�c�Q�R��W��K�2ɘ��i��}G�G��`���i޴6��2OUޮ��Z����<n�gk쫢�&(���7��)x�p��P���9b�U�����)�	�~c�u5-y�\��*��q�����HYJ���ciz̆���|����r�A���3[F��H�|b5���Y���*�8\�.���2���a�0l��9�#��0���
�,ot6��=���=6 8�}%��WF��յ�k��1\�yLt)V�#M����2X!"U"�]	N�b���v��pn�kcrX6�Իr�r�퐍r�[ksύ���쫶G9zݫu��<[]t;M� ���w$Wn��ʭڹ�K��-m����F۞˳L�G8y�[����Yݺ�ܣ�d+��ǃRE���jۖ�F4u��8-η;g�\l]J�7> �i���i�ub�t��F����@��i�܆�b�n.\�5�f�)�ָ�t�'\�n�35�"ݹ��u�x5����G8v�Cf�\SI����8Pl]��=V��:�Lgyym�+�Ga��
��7�R����Qߞ*U�5���L)�e�Y�˔�-�k���i��T(�,)e��9�Uc�*������Ekמ�|W;�m{��[�3%����wR���Lp�j���<�F��`�}Č�ˤo�@�vs���a�G7+�p�2VZf�P��t^��[�u�x�Fj��N�{P�f�Q�-��Q��%��+�+��D���b�q0
ǯ�gӗ���e1@X��&�q e���$�m��6�2�1�Qmhrӧ�����B�Uu=��rg0i)���q]fN���0�u=��(��,��A�^��{D�j:z��QZJ�,�����&�2��mF��w!����ǢVU�]W��i�CQ-+�	k�Ϯ�:8׽�:���V:�ƚ�	~�X�{8�XS-2����F�L\�te�8��o&L\c���=��S	�h>�"��UH�m���̺b�/6�~=��/q�&��S.B�/Rp�Bm/�U��[��H|�̾��I�MP 6�y�PRԮ��Jb�	�~����7�&�k�E�Q����,���U��Q�ӏr���A+pJ#.;��G�xlo�)J�	���� Vw2�`Mv��W�������RF2(�@%r��o}�;��^��0�;��;�yeGt�?�T �M�-����u߻�e{e�͜J���^�������v.U7���5��l/8kFp��#Y�� ��U�m��t�oX-�2�g|������[��w�y�l�ھ��=�S ��#�ث��۰����ُ|cwՑ�WtɌ�<ؽK�cJ�EP	Y@�m&w$��`�\�ʸ��fM2}�t��S�s��=��Qf{����4gP;۲����E�����������w�g�x�*p�H*AL�qחfy\�6ݑێ��:��X��r�D�5�]CB�t��L6�������O���p]�[�]�6}0�o�r�.�9�i�T��v��7��U�D0�>�+D�^l�v&m��jm�L�� ��m{�p�û�N��mmw�'d�Kޭu�⃺�~����<�ff���O$֞��&����~�N�!���-��H;��H��"�6U+G�.CE}{��yP@��ڻ0-�M��X׷��6P�su1�yc9uҮ�cՁ4�s�5\��y�5�	�Y��;z�M��%����i��q��1�kSp[=K+.;A@|o���L�g�x��6z�Ѿsk��Z�c���b]���$�Y(��.ʈ�է	Q�g<�Z�i��"*��o�u���|fk��r{.�(eʻF:���ݽ!rE{�mL9�0�>����h����wZ梚i��7����s`�Œ����U���7�9����'�D�e�����D��4�{ �¾����[�[�K �a#���u���:�k��tv�NӞ!V�1��|�;�+�B�* ʉ[�[V�o�-]�����t�#�eJ*/���p�H%���0��Z9e#~��\��{��{:���آ����}�1�tv��D�04�<�F�n��qYpN��f�F�p��$a�ؐ�+q��K�r�n g�V�5w����/�׫�%\�ee��g��(�t"Wł&�7.x�F�>w.ܻ
�]0iSD���冤U�͚��^�g��o�s�מӵ�����'���^:�]2�������r��L��^�=#p��ڭ��2��G�F�j��6E3���������\��8���﫹Ū� L�R/�n�Բ��/��b���	N+�7��1Z�w�F˸�������nϢ�먽si�϶���wn�'mJ3����d�����r��DD��l���T-��@rs�mY��w~7$�	�����'|������:{7��).֜��$&^?��1]@����Q4y���g�������;p�ݺ���q]�y�=[E�.��z���t������~���kf��q�.�l�O�V3�{�3���X��oxy8��	������o�ʸ���&y��uX�!G㒛�Ծ��]��ٷ8��Uf�g�8��)�i�]��G&�5gI��H�HR��ظ�d��p{�/X ��Ȟ<�@�	P�D�6&��۴�Dmʻӛ��U��i�f���T.H8���u�{ʂK7f�sN���V��6pot��,�^Y�X|�r�EX���*�6 E[dļ�t�!�~�8"^��t��w��(L����8��&�^�ۖ2V2���J�x�w���[3f�b��-��9�̎�,���m[\v�<[;�ߩ�Ӥ?�;.�.�:���Et��U��w.y/��g�פ����P������6���U ���
zG
]Ji�bZ�zI�B��eֈ�*V����s5f[r)����J�$vJrM�i��x��Rn�T� �Y]ԏ3����V�H��AZԱnCY,�6k���������]s��݋��s�5M;����ŦuH��uno[l�����d�=l����YN�"�7�7 ���5�m�=�wK�W	��ûUc�Du�� �Վ�"=]����㋌V�=��p����x����c���X}��j�9ӫ�������]fOm�N�Ig1�{v�s2�V n��睻�Tya{e�:v��Wm��ټa��χr�,��9�4��n��]�xW��E�����1I��P1��Sj��n�Ij��.t���Ke�9���n�,��o?�P�]y��!������Rƈ�-��[��
gϪ{EE��#}Hn$��t�p�ۢg�&P��^��$��;^����=�w��M�����}Az6t�����+�~<6�:N��L�LŲ:`)~�����R %�ku��ׯl{��r��t3Z\�M�.��\��y��l���<|Fz>�.�K��aM��t�-|[T���[���~�f�|�|�y�͕([�9�(�Ȗ�W>���fYG��^D["��J/(,ѝ�c�QS��X��XU���%�A&ͼJ����g��-�����
�u3f����D�ɦ�T�>&��{>�ʁ�1�}�/�rɭ�lO��b���͂1YKqj�5����Z���-���}�x��ç�Ą�Ԧ�UjU��Y>Z��)�nTY�ӣL�_�v䕫2�(�t��k%�qm��gj�J|�gz\ޝ�U��l)7��߸�4^/f����F��&]
)�����Cڷ�R��[�7�l����_��~���H +�z'���:�(`���R�&a�c����^��죟A����o7)M:������y�=��f4O<h��0Z���Cճ§���1�O��Q�Wj}F��i�H�uu�|Q���Y/�j��M��i����OT�6�~��x��)O��׵X����oL�Ib�������m9ah��u�#eӖ����Q"�Ö�]N��)���B*�e�T�4�m�i��9^�FOkɡ�t9~�g�?�T��䪟�(9�K9���7ޤ����j�#f�g-����(��b�n�w�f�����/Y�+{xORV��7�Y��8VQN�6�Z�u�fôT8��Au�ۮ�#%���jv�ְ;(JY$i�X�$�������+hR@�ߥ{dӃ�E]�y�Cb��?�
��)ZF�F=X�)��X�o��Frt�����05$@�6~V��\�DV��+t�1�!M���a%��Vx�7�N�[^�!�;UZ�կ[�����xӫ�{������J�1����Yd�Eli����t���շ˛����,�{tq�˕.�?�)�5Ӌ%ev���`
���n�XǾ���˩��f����| ��\���v�s�PN�����֑�|�T�v	�a�����V؛�=��']]����{)C ngIT��u��3E��`E2�$\�<����j)l�[t@��z�	�n��uؘ~r�n������G��x�[٦��W61!���g}�+f�f���g��2��P(Y]e�X�i���{�Y�rȱ��zY�/y�|W��
����;@Mi}�W��պ+�"�.��&����]�����.�j���_[,�g��8����-٦��q��tձ�T偗Lpή�w�R	ǎ����Y�'f
�eʽQӀ�K�ZY�~�s�����-�O�gk���8y���!�1�N����W/g��P`�I����˻;��$�*���nOm{� f�ȩ��W3{v��j��?�_"��]�`�����fd��.��]6[)��)����d�Χd7|���y6`<P�J�w<�G�8%K��=$�.Gn�9�}kx��5j�tz��e�Wdp�"�N3�Xt}�!��Be]���X6���Z�E�w/�bT=��Z�݋z�e)~���f��s.���!�L2:Ƌ��qL�ʋ��Yc(��� Y��i�IKs�"����ͷ�oir��]����,f�l�T���)����Ԛj�tT�N��ΗS�T��і�Q����٣F�ȕn���m���3���V���Z�3Xs���^�^��[���!mo�!�	�n勫ls�����<v9���	���˃cC�bN;�
�9SAA���os��O{Yk��/��|b�>A㛫�OެgV� ~��nՊ�¼{�͘���}��q{Qx�>�D��-�mk�z<]�K�L�f�����oj�&��]xn�۬�s'���XƖ�K�/{��w	�}��i�6}vwG[�oi����E�Zb�i��c�O��Z�]r��h#n�*Y�Z��ZԚ܄_��@�v�ȃ}u�P��*�Q����/ou�	�D}�M�t4����BIj�ŮH�jo�g?�)�=����J���]�xs��Fr�\�L���:|����=��b5�������Tqgے���Je>
��Hi�E�I��g��C^r8�$�U��$a~݋���o�̞�ۑ�P�C1?ef0��4��x����Ѣ.���S�⮏��p���]�=oTmm��n�����5�bJ��%�V(�X�K�{$X�b��N�t���9�8��m�<� ��k�M�.��p�9u���m�[�1�}L�*��_�[n��lZ�[wz���	tC	\��+�:��31�E#XwsS�����u��]偟%CE�ݧ��c�q�bq�u��j>O���@�^=]�q���uΟkɈ�Y	u�����D��������pmf���0���Zzvgl�a$%e��1J��eg;Mʾ�[�(j�R�JT��e��FZ}L�';�2�+aK���Ս�]%:Z�"a��h;����]�ԙf�l5,k~�SFT��n��W�}
r|i��(	G���ח���a�w�ЧSC)WR���3�MR����UKX�Y�y�뙤@/u9*N�9�K��ws(�)6�&"���u��i�&3�ڌ&.�y�զ��z��DY��XUy�i,%mqo���QR�G�#����@l=�9�L�hc�IU�xUq�͛ޏ��Ok��i-Q�Ɉ��МZ9�]_u�^�8�ᦓnT#��_\�6��Q�c*�eIM�ݵ� ��*ˌw+�W�b(��'��z+�/F2�t�ё����M���`k�x��p`�u���3�����&鎸��/DK5�|!Zm-d�z��^�/��c�&����%��y�!'(I$��h���E�ɇ��O"k�J�곰�y۶�BQ��bMל�^.�n�����a����5��U�����aDb�wx����s<\�p�M%6=&��"�P�I6�Ӥ�\l��x�x���v�]�7��6L�M/Y�\��q�:�pq&Ӹ���U����6kN^���q�y�0k'/F�v�5�+������%���ɒ�m&�^��n�c"�AӠ�JD��H��av��1Θ�rx�V��Z'(�N.����uo+��z�f��ÈN�7��w�gv�8ݎu�x�[��x�{f�-�t� aw;aw&�g:v�C�#ל��+b�vu{n�E�1ѭ˽�H/y�V��;qӚ.Y�{^L>�Aɺ7NGdr�n�I�#ә ���mG��.��iK���띞"�u�7W���J
���`R.wg�S��ʂu�6�K�rpqǺ���[Z���q�������G9}�^I�ٶqsp����n9���ܗf�����/W"�ݳɶG4' �u�[m���xZ�q�1���Y�]��fD3���e���$����^ �9xk����<Ŕ�]p�5�8����-�X��lX�5^�ɻ]N�[u��%�g���n��`��	z|�n���.�u���8�w%�r���{=v���41nOu���M�n���kn����H��X��;˪�oB��X��e��v�j{�zpv�ev{LQѶ��l<���q�=(vqy���\2�2�z�n1�oY*��띱��{xm�(y��u���������OY��v���8����X���!��x#j��[��.|G���4�����D�t�Zy�lqq�h#�,�Ύ;n��8��w�2<�����#���\G;x��=��������y��ε��ݻ^��`��tv����'B����O�W1>n��,�{���όb��G[u;�wFl�r�h���� �Cpu�0��]	��wE������<���u��Əf�b�W��{:�5����q'=��Sk�#l�8z���:]�IF��tny]��2�n����[3y��� -r���RY��Nx7i��m���2<f1�g�[��y�#=�i7`4x��AƔ٫�%A)~�ڨ �0�A-�(Qn{=7$]O^;%�ny#�3��%nŸ��&�']���vr�Y�bp�"O[g�u��kOM�7d����,q�4	�n}n�X뛰ۭ�[d��:|W6��;�ݍ�q�I7��Ŷ��5�ݫ<v��Mgv���׮:|=q4�u���uWKT���]ns�l�����,d�Gd��v�(8�4����N�W������Ԇ���e��]�l���^϶�=<s���]�b�����ZX�e�,����9̝ȍN���'����u����f=g=�u��c�;��j��e�6�=EW�<46�ft��fuW�Z��P�CQJ���ؖO�3�fc��߯}�$n�l���^z4��]@��y@5��I�(U�j�L÷�S�ۃ-���Y�WIՇkH�JL��<�h�BI�%�ukh
Dh���4���C*��ýr�5.�Q��;����oO:h�a��ι/2N�z��]������z�@l�Q�����5PN�����Lڕ���G/M��;��f�S}�cl�� K�6�}鵏R҇V�NWz�&'�[s�5^8��X�{��4z��V��@+J�����,G��=sbD>���Jw]��I]��h�3Ӂ�YWV����9G��eJ}{癞��үH��ؐ/]v�^�&���qz0d��K6���q��%s����,����u�m0qQ�u:�������+;z:ؗ�D"I�޽����'7�b��m�^��E�~��e��<nǼӣ^�m�U���i&�2�Gz4q�g�>x�a�-z-ݹWWeu�3+ҖL��ׯ�ި���tC�gkJכ��}�*��I��T���#[1]�2r�`띓5Ly���{�/Q�C��֟q���!o�����m��fL�A����qg/�y���M�c\M;��zZ{�'H�%B+����ۘ�b�8؎���Ɍ�1M2S�ɓ���z}y��wpr���_����'��k7��rjc΀�O�Z�S(&��I�~̹E3��
���E����/'2���h����dݭKDe0q���ݴ���6���*�2uE�/.��u��j{F�P�dTLt��X.$Ǌt��=J��/vso��©}���1��Jp�� :�M|�NU���.�Vc�7�P_CB�u�E�0l�l�DW:6Y�S��8咳��|D�Mt� Z�������m��x�zg�_Mԇ=n
�V�{#�dTDK.�&ol�k�ys�0�:�����-�ײ���4�Ț"t+��Y��2�p.g<���7�;=�7��l��gd�~OxV3�%u�=+ �w�[e/f߳jOv�{\6M��
����HGv�m�Q����kf�������O/�e�15ܩ]�����J�G�Z�7qRe�WY��\��$2ӹ�]֬f&�*�������kw��2cc* 
��;����#}�L�^�%�{��سh��2�O<,�XE�$�{�~�n�,��N�i�{��{ך�C��ף�x%J�Vv�2���n�۫�C����}1������NY�^v�=d��EE��	1@�n���� [�=�E�x���o&���K\���~[ii�,]���(�k{{+��Y������mk�.x*��Pm��%�@�g1�0u�Iez��!#v�׭�7Ek�΀�G�qYb�(W�ZZ{\�s��+��`�����	̑���Ti���O*o+z:\����(�w-�n
l���oQKFJ����i�#в��@6��\pY���T��w�{)M����Ʈo/k�|��A-"���˽��պ$�ste�."�.�l�L���˙%J=�J{�ٞ�n^��K��h��0�U��znOm��W>�]�%�t9���s������:h���M�z��B��Ie^��/�2
��Zܻ�Ԝ���9M��f�1K�k�f�O�n����1=��^�[��[�9"�zѣ��}j�}���d��s�&*ET-K�}R�����rL���	� /+�B*(�=F�;�W���E����kֲ漷�8��E�
z(�[m�*�I5ϳ�٪�yJ�Ŝ�s���0/e�|��Z�����C(\h*<��_�m�v#���%{/�꺙S>���V(�w��T
��>4H) Rt\�Ɖ�Ȧ��³��۪zC���c/#\�s��ۧ���(2�,��^�Z�*��W�o\�m�es�ɬVSD���¬��ۺh������L�9���V�8�^��)͐ۢ�ʱ@bQ�I���*V��#��7B��m{�����/Fȁ�K�7�ĭ
k�	��|J�x�)��ޗ凹����� �~i �a�I*�����$�V�
k�@��^��+�W�Z�)s�K�|��gL\h��Z1����m����$��JEX��(P��O�=i^�Z��s9�<w=��M"׏��v3���rWX����Q��/���ѿ-=]�^�k�xr��fg��S�&ݪ��d(�;l�ր���Ӿ��ʝ����]IKӹk�V�z���e�b ���Ȼ˔��]��)��m����ztͮ����:�����D����:���`+On	!B�5L�p#g��m���S�'XE�gV��]���4�|b�\M�2Ӗ�#���d[�4��D��y]g��ks�=�t9���oˌ��4tJu�[sˣg��jF�c;qO8��X�f���F"�y-�{�s�֫���7@ۉۧ�2LMu�p���n���)�v;t N�K�ۄFL=���&L��&_]�v�'7k���1�Ʈ�ǧ�Wmm�|�ۜ��<�s�ۖ?����Ӝ�.��D�眵�#]L�8����EtkPZ���Sn�<#��wI����1�r����j㭲��lbT�IC�޹]n� ��g�ߕh��k)�So�u��2q�'�����)r��g�6��.�z�ݍuA���-,�{H�;`+J�("KN��fF|h4{�6���:���Od�f��C��)�yx[��Aդ�~�>кS�u�.��U'�������M�������Y�}���WuaJ�N�'�� $�Y6w�j�X^��]4��Q���Č�������8��&� ��g�(G��Y�wW���!�Q=�԰�6F�X�Jp�Q>��ro#�Z�z{=�{�A�KM�>�%�E�i?J�ie�#�B�Ż9.�;Ҥ9Z�gY���b�WtX��W�My w�|xz�a���=���Ku����ڒ�L��V�#�{�����߫�<s%no�� �3���q 뒵��X��\v]�y�0t�l4�fU�����iȼM�̞���o�(ye���R�k[���sy�غ��ة��Z���ە�tTݺ���H'B�e��}Kx��	l�9��oa]G�gJ��}�*V���a�`�6^C�/�YL`S�̻jnh�Ro^�ŉ�:�VN`�;�]
��{(�W`������\�F�O__��+�_��Z����	6zK�t{�7h�`�72k��%w{s��{8/F����,(�֗}ϫ
���W`�ټ���O��wG]k�!�^R�*<���=yo�q���**46����ǳ�9͟Muz�c��,�IC9�m�.	;�ۻ[���}e��o��k�t�<}��D��r~:�ykhQ�g��6��=���
��H��j�J�1&��;>R
f�On)Yj����řSިu�xT#S�o��RS:��t�%�mtz�\�3����!�W����|,%U�V40����S�WO����=���N.]��'��n�W����l�$���#��Yb�(�����!����X��v���T��v<�ox�.�
�0���I�g��ǧw;��
�VKEP&�)�}��Qu��^e�����{B�=t��^����v�2˓�簓ƕ��{;�L���9�2���2�����9=��`k��;$����2}�o_Jʰ�Vok�x�����54��7�fЕ{!�ڞ��gR}2ol�ʸ[�뻡�,����{+@e8a�s�ɗ��/㦥�@􄟻�w!�3$sl�MҾ�z��>V�N��X��wP�QJ�_�R'mFR-��I�e=���5�1ȗ�lz� Iߞz�̹�D��̽W�вx�us>���O{6�1mt����<;�@��	�j��ߔ��2���Վ+�Nϻ�x����k�}�l���ޘo��j�õj�m���I����:�"��ۃ8�Y㮽#��-mL�����`M����y9��TȘ�l�����G��ٗ�x�W��J��m�i��ٻ^m�Q�a/<!.����N���BF�4�a������;�Mg�\�����������c��MC{%)��\k���䥊���T��a��nUm;��Ⱥ����~����/��fו"H��I��c�'�A�#����12ǈ��;N\����\�[�����I2���2M�LF���%�+��? M�Պ4X?$���c��Jۮ�r�t�7�h=�y���#f��/f��z_��/a�.ا����_�R��G*C�&�9�H��+lS>���H	ųEJ�9
�R���չ`k���y��]���ޕ���cx�6��*w�u�.β�1�{$��$
h4ZI i����9��~FU��N���]Kǲ�>�z�k�a����y3�I��s����<�2"��b!��ஸ��S�M:Dѕa������:�nCv������[��ֹ�KQ#��P���hv���;qnw^�̬����l�ҨV�as� ��oۻ�u�G�,U٪F�.�֏>��J}��=��E���a%�s��2�
�g�4�yʁ0:���Ǟ�����/�F�K��Kb�DF�y�kw��N�@�/v�{��.p����B'e���)�� �Ͻ��.4������C�WՏ�	%�7+�ν�l����͝5�w���n�^ݜ�t\K����㎈懇'��H z=̇}�[�(z��8㩥�R�������8ٯV]�~�TH�g�����.��Jv.6�u�RA�,��l�Ͻx��O�;���+p��7*/Z�ɘg�du���b_~��M��{E�u/�zD�H�Ȥ��͡X5}�0�HN��u珅���P
q�5�\�����#��z�J��3�<C�E�����ɤ��3�oIzF�W@7$�q(�˅hov$�t-K��e���a��l�=r�э��v���tWAX��^�>�M��î'����w�\Q�Ӄ���;���Z�!�qnwO=��җ� ^���km��Ҽ�k]^ܴ�k�گ	�\d;��K�U)��zl*���=`���L�$��p���8�[���lv����5ŝ4Bn='�t�t��\����.w�l0�B!L��p5��n+��n4Y�<�n��|t��p��WIPS�P����^�yb���O��3�@k��n��횛�j�=0��`:���˂�&�(�vaFք=�R��vE+��%unM�6T�^qu��짡��X�S�����^���(�����4N�����g,Q����ъ���N[�^�+�M�C^��F��Q�V0(���m���I��,���r�٥ew���{l﫵��^�pmOyN�zv�=qg��z����Om9�Q�"`� �RIb�l�WS�����)�B��~�˩E[k�n����t�s��-;�W�u���^�wV��!�� smA0�׼_�J�(���6S���j�4=����o�D?s�h�L��t�ou>�𓄉m�C��J[�2�sx�������D�G"lbv�"�Y����zN��.��n㚌����un��;Q��UD��*4�mS�����/�,奁����zK��������v���r:��mY��d�����l˭��D�Pn���	�Yy�2թ�;������;ZC���-��gj�P�o	��|��ڎu�f__2E1��0���^��)�%�-���F��+���)Q�@Sq�]����g�j�$�=O�q��˺=�u�%on�MvP��I�B;^wRY\�b�:9y�N�a�hSm�}zVnv�=�ڱس���:���<q�I��=�#0vs�\��KyL�L�ʹ�T6�����2��禢#�!KS����o�J���nS
�M>�qK�w���ܮ�m��(�ݦ+xzo}rOF�߱�Q�8a���S�`�������R�ծ��=Y�ʺ۷�Jt�W�:+]����^4X喪�J�r�lN���Z��-��b�Y�g��c�V<�$���f�tb��9]P�`����5v79�4˝��Nh�p���麎��{ �]��nu^�*Wp���n������f��~�A�hes�h���w������k�������9yY�6sj�� [%�@m0[lg����פΕ�}S|.'E!��� ����U�T������ʹ:$x�oY�<��{5�փ������¯�I`����I���`,㾗�����wJ����ns�9�5�M[^F�׃M%)�^�N�Њ�m���jN��Ўg۬ ��f:N_R#�
H�ن�����1�U�^�����$�k|�mO��\qʸ9�T
��w6��w"Yb�JJxؼ���{���	Rr�rX^ӹ3(��-֬�ۍ:���XU�m�ﺄ�PJ֧>�����n�^�F�ޔ�N����٨"h�LN]���Y��S�'N�9"���lNWR�v����jݚ�qn-�����P� ��;���Ԁ�R�8��ݺ�q�(o y}����i���ؙ�q����-B��bY(*=3�{�M��2�T�Tl0�r�����Ko�xW	�-���m�7y������2r����'У���o/U]u�'�.\��9��k��suL#^#�l�]�"ה�ۼ%�����k�K��-Z�tm\W�i9U���˵}Dw�P��r^���9��4�ѣR���,G��6�o��on�vKn�^ņ����2�����f�����Ca��C��x�s�՚X'�3�eS4��Dф�Pn�5S-57y��+���Q�^S����/,D;�]*��^X�ą���ԨңQ�ö)���ҥε�oOH�YOs.<ABG�ځ�۹�w�tW��s-�L��d,=8��\%��3/����-�Ʊ��Ӹ�[�ѹ5f�zF���Y�f�ױ\��	i�ݕ��y.�f!Xb���Vݳx�6�,WMX5��K�M�)U�>�7�O��ai��p�pXU�X����O���#�����;�P��Y@�j�|����u�"'P��-���_E�P��=���\��W�R<���ww;��^�E��� ��l	�Ď	���y��} =M:dP_'��fm�pLYfTv_��"o.|���;����Q����x��)9��k\i�y)Z�-�U5j��ԙ������c�ύv�:7S��9;p[n.۝��k����}p^��E��]�U2�;��U�t�wwx��g�M��o,�g��&
����X��`��v�V@U����T.)�K� (��\�>��wcǛ&�R�@�(C��H�{V�o��K�MKR�q���Xm��u�:���`��9�w�����J�rχ$��'��s޽[�s�N������+5�a5���u�����zPƼ�q�����95�w�!n��W-5�35���^��Q�d�-؞3��+���b�{<�����%�6S�9Ęr��i���6��n�ľ|����/N��P��2sQb�����4�#\K�]8U��d��v&��N5��f���c�������Ĕ�u�{I���%k�b'�%�J�Aj�
^�Әz�^��-c�U�{�a�e�}�����_��mR��X�9���V�m�d�qÓu���I����6y���oC����^��7Y���yNq����i�#Ǻ묘"!B��}�7ឝy�H�1�ބE �&����o�OW����� wv�|[M���u��:[�~�镍���a��M��4��� ���j��!?8"����S=����hx�
�b)Z�w��x��$���������Ngs��\���AViNX����ԧ`�mЮ��v+��>sKuh^8�Sŋ�2�k�w-����&��=B�������G|0wl�ݾ`L�f�'n��-�
dٟOu�'&7��[Vh^�������u웠�*T�M��I�e�erA6A��f��dђ���ަ%�������by ��j�uR㻍�^ґź�nϹy����/��}ęt��Y����nh�"%��'31�ŗ�s���¨u�ћ"�H}��$ن���b�096�DL��KF����\/1[��cB�H�j��B�P�b#�I�	a%�з[/C�u9��p�;*!2K]�rv�䰽>�Y�nݞ�L0��]H�V�k�n�i��n�V9�;R�N�rs�{�X��9�S�:����r��v8�2k���vvA�6�����ۢ�T�.�u��7>�9]�<����F7/c\g��ͻv�[���睶حU��@"��9�ۘ��Kr�q�,tn�Bݷhq�zzg�=��+�b���t�Nz ם�Qݪ��^�+:|�e�?{}Ν$��C��k`��V�a����ܔ��]�t�n+Ɩ{�.����T�Y��"�)t73r�6 ���r���ֺ��{#��e����6�m����J�M#yӿ�Iu�er���-n�E��MRE22��H,����X��׋4E�h���}4	pV���^�m�Q
`��=}���v���0U�	#u��ܮ4p6�t���e�����*m{�S���3�dX���c\>ʞ��R�{�S;�,;�l�?S{�V�Y׺�}�H�i�xEi�����N[k�έX����4���t/��{�ۗ	1��=�[�V��\�Qٔ��xk��o�l��kO1{�K�*�h������X�m��h��6iΓcqz�W�Su��:�$���( �U�Pj ujf��p���O���}��Y|�\gYohd���ߦEǷoӽ�{��e*;]f!IqS@�E�%�#ˆ�ܜ��~VV�M��W|ǘw�d�b�˶�����+ή��[4h[���J	wu�+F��i>$�G�)1ӹz|:px�Ս:gUx�O+��:S�����$ިl���7~^s�*�xOF7&��mP��J���5��[a�--�nJI^�H�w˾s�7�6[��4����9	H/L�I/�_bبzf�fViL�M�v���S�ا�����[-$����-k�}5ܷtK������]*�H��^��j���X�Dy��5wjorP&Q�Qy�6��kK-w'�^�P������8��8>Wn��\�{i�'�m�7A�ﳊ-�J]��,9�v<�K��tG/��M�(��V�Ԯ�Ir.�գHk��v���琫С�<t�Z�v+�R��#X�<\�����S����M�s��M��o�m��8P��5݇5h��L�j���ɞ2h,<��)���S�6���n�z�֪����`�+�]�H,��MbT܈g[At7='C"yFf-�O.�o<C��=x�{}~>�Nd��z���|��F����6	�%�%�	�mz]�/k�:}�4׌h{X�=��K�9��*��W�zp���e��2���>y����U����� ��0ϦJZ���j��n�b� �[����[�v��������f 7u����rڢ����xG�E7�Pܖ{|�[�\}�&��������_G8��];�[}R�kUj�|䩵�l�'ᵇ�Mc����̝�o!v0�������stR(�,*6���Y�/������ܞ=�pK���qn�=o(yf�N�'��E�hM<����̽�{�4VV�s����G�:Ԓ5�V�*�bZt��nr��qp3GH
0P��<FX�V�?�Y)���{9~����x��	d���v�-�w"���q�j��%?��]�>%Ȇ.��̏~��ITvȜ��-�4Jz*�F��sy;ƈ��ٛ�ׁ�l?��54/?cR$
����	Q�L�g컪c�&B��4��\�!��w��\+A�D�č�/���T���h�s��OU�d}�1���������$ѩ��B2���]Ƞ
>t覕�;�X�P��W��`�Ǳ����'WmФ�ߚf�ީ���Y�/r[3��:�뼹�Y��t^"�HU��y7��zx������]��N��������Cc.����Κ.0��H)��3Ku^s�7���ۼ3w�[�Mʚ�%[w����-�E���~u����O�殴/��0�l�{\��-�����y�Qw����|os�Զ2I�x��E9x;Z��\�����|�bbl�*�7�'a|`��v�籧��7�ǒ�8�WKg�c{=e�@6���gx�y����-��~���2M��Ďf���v�C����|˹��kop�m3/��G�%@ϡY�b�Ri3['fL�m����G�c'e_x@Nb��%����~G0&V�c����_��_%�!�bZr�W�t8�L�e$�97�w�3�x��+����yV�������wꅷ{7)ۖ�ݵH"s�q��{n�{<�x8��,�C�[M�Wf�ܘ���2I��v>���1;�<״��
#
�8i=�e��VOf�\��������$�/�/l^JÜ $�XdP%&�M�:��Q�����:�Kͭ��'������߼wml���jC�t���2����!����ݧ|+��-�ok� ��OS�5��.�E����#��=ݫ��&�)obԒ��[��T���#� �Y�d�q�i����q̈L8��Fɔ,+BҫR$��7&!��g��ۄ�k�k�t���絇�X|������!�\;�gq;�H�7e=���]��K�xӵ��7mm���v؉���lt�����!]VZ����}��`�:��\����ӓ]��gn�	#G\����pt�@��:�` �mv�n�[���kOA����y���Pq�2tQ���w���͎H�=9�ɷ<]��۱��d.�駶�<uѢ��T�Ay]�7�c��s�n`�N{s+=�7n�NA�~�|K����Bg�]�ܥ\��K�J�쵴)'��Y�|��W2�k�����Rwy���e�`�MM������;	���me3Ə�i��V�ζ��jhyP�W�+����*yU��n��w�F˩�8wi���S��S|�/:2Q�E"��q��G�+�ʷ�@��@�KVy!�&�m������E���	폯�}�d�$R�	w/o_;��-4ۢHhU�Z����4`�ymn#��4旗����}ƒ�aXh�ֲ��K��қW;<��;6S4�Iȍr�B2���;#f��=՞CP��T(3�e{�=KǭQ
��s?br�{q��*�4y��}Z�9�ԗ��B��͚����]y���n7ɅI�EZ)�ɹ�����6�H�<�v�m��Q6���QȜ�Rf$/=G�hLh�}eB��%��x�����ڟ��WXN�e�d&���ny��c�gk�%���d���)����uf{笍~�o-�i_"�j�+@���"C�*^dZ�z�gբ�>B��e�"r�Y�����t�`z�]\\1W^�#×˩�]T��nw5Y�f�ԧ��D�:��+����X�l5o]�EX��L�tVZC:s�ٌ���~}�Gd=��h�9��/6�L�>��p7���}����ׯ"���� �o��2����x?J�'������O��,ɸn7�;٭�~�y��"Tqh��Ζ̼����l�an���`�(w
���N��;��d�H�F��׳��]N�k��ϵyV	�oJ��aJ��uz�*^l�&W���QV7an�H1)��3|�6S��Ѱ��w���խ��.�k����*��u�>�	�s��������F��y��0���'@&��h0������Ś�����i{	��-Yֵ��y뒠Z$�]���8��mͯuS����w�o�/ǲ��W�n��KUhh ���
��#��&XH
��N��?(���(f�I��(��\�V����B7F�c�w��ّKwK������8�cGv/n+�����y��~*Rޫ��\s��ע���w�>�@�n� 0��א���SV&��;��iR���C����x����&�o���}�h�\�/�s� U�����wt8���6��y��䠌���G�ͻ�{��ɬVωn�9�_R��0���	D�q\�|/EG�d��zF� ���%+�;t�R��GY���+"�g>�!݁��%���j˭�_w�}�PD����XG��qnl�%�E�#'q��B4] �2�I�1�誢��ܳ��JӶ��Ϭ���;͛Pje��M���XA�]��<v��~G�;03b��	�)���T��ܷq%���9K��9�8��n{]�n���dŇ�m�X��Q�O�~q;-��gp+<��'����8�q�t�q]��
�/f׮�{\u}Y��)sJ�X��i� �`��=.��
�A@0�9B���3�w��ў���������{ä���}�|_��{�����L��{����6���}��*�ޣf�x�	U��A�h�A6\���d�[�{�n�f�-N�H=���N������t��,�=ѫ���f�#^�q�����V��R!��ͮ˹N���/�ѾS�+da�5����n����xIv�[����ס⠜��K�)Cp/hw�9z��Va2`|]^�ߵ����>������u���J��7Vd��l�u��S�©Ã��m��}t��y�!@���� �EӠ�m��&�ˬk�f�8o.d��ې�0�!i�^&��gd���}����%�'�a9���I�ܴ~w魌ub�m��:۔9�r8�t��m�3&;vF�z1F�@^�C��ؓE�d�ҷ]X��j�rd��S=��F	o����8�z�Wr���Ł��3�[�S��m���S��J��&�������L��N�)�x%km���~�50��l,�㗴8N�o�����+v*F���\k|�Ҟ�������tAg,tЦ�:m{�~�!��|t�M�6�i������}�p�,c6Q�h��ь9F�=��n�o5��׺g��n�*�8�^�B�@e4J:4�II�D������Sz�t�h��gwX=vsՌ}������r:YŽI�����<#��l�P�1���`�}���-|w*�Ǧ��)�*�m���g��-���^<�x:-.1���Tm%އo�w�|�Oc�&�g�]w�_.�x��bTј� �[^dg�-YRJ��[��	���Ѥj�{������t�6�"��U�^.��@5�vMLv���`�#����3e�]�� 5��$�ǂV�� R�Y�Yh<�W�	�}�5���=<�M .-X�Qsh��sn�G4�f:
��&���o���ܣZm�y��В���к�6[��v��w���^#DW�2����	3���tV��m�ɡ�FeM��9�!�TO7�v��l�1J�ka��i��h�S]g��g!R�6�X� x�
I>绗���.�sj_	��d e,}}���>]�F��',�*��ŞξC�T��A�����7WK�Q�0�e�l̗sM79��Ɂ>�Nw{-�
�ǆ��5��Uݸ-o>w�Z�R�uo1u�f���&'q�wxU�==������n��"��P� �ha�f*Y�R���C��]�M�=�}�r�z���nq2fQ�
tX�ʁՉ�6{�IV�q����-䣾I^�˭��j������X�)ku��^�ދ���ۮ%M�[Rxᾣv�Kp�f+}>-Ĺ^�2pKTq��2�5�Ƭ�J�TI�E5*��dk��Ef����0��CU��htޮ���ܮ�^%�V�|�3U^��C�Zw6�*W�tb�reM��]x��-�t@�N������xsu:Ϋ����q˚��s*+w�z����4_t̠������;Ԩg#��o�L}�����{G�.�L�bc�kx�nLw�,�{�Q�]���쿤2���s�Zp+ur��I��JK�%��ݕw���f:l�e�������,b���.^�,�2{K��E�ݧ�2�p�i�ĕ�9��؟[p��7c[v�l�v�Z�:�,�..T�G�u��Y��o`tvy�jw�y���<�F�Nӆ�3�e-=N��t+�\V(6孵��`����cq�[s�5�{�g ��-�����t;b+��>5�x<;y�F� ���� e�8X��ҹ�+���л���n�[�|�n[��(.Y��/UC�e��`s���r����ƞ8y�x�X놢q\�7K��<p<t�%�G��B�W:8^�SZबE{st;�2qx��Ha�&�6�)�5�ׇ����nxœ�{yvz�={<����|�8ݮzv�ڵw/�vu��n�t�,q�+�	a�c��S��䡝׋�ѩ�{��n���gCV��{z,o�����^uZ�n��q�մ�/Z˭�n6�u��Pb;<�]�ڀ�M��]B���ݳ�֑�W"�.�<5��$�kvݬg	c��\ۇ;r\���	�VUbk"�,t#�>��P��uvݸ�:�j.g�ù�p<6�Y5�-�ݐ��ݵ=L�ڱ\N�3��۷Q�^�Gk�k��^;v2]Q���9b��q]ג�[7a�=�d;/;��1��u�M��k.�v5���l���͓��n���O6\�ُ�W(nx;[Z��m������n���+��Zg�K���Ёϱ8Ga�슷V���W��6盰��j|^�U3�V�t<�u���F������Xl�L�]���	]�箷l�-բ��x����q�]�v5h���ՙ9�WXv7UǞ�F�.e�U�s��x��yCq��pVmt�3�s��nw�OY��V��rl�t���h�qa��g;�c�MX��z��^�2�\"z����vS���y�l���5�"a3�@�Uu<�/ [3�����f�<������Ҷ�8��[wR3��;V�2]�7j�w���eї�k��m�mn��7+��i�vt���%��I��7'm�b�^c�Ʊ���h7>���ݺ5Eۧ��;0h�w_=��c�f:����_[��7�bv�瓎�h�Í����n#���l���顼�nA�����K����]F\�˂�w\���c����`Nr���f���gӷ[Ciz���X���ě9����$:�#�pv�y{l�����ܱ���'/8�z�ʇ<����;uf䃸y-���8�i���e�\76��'\�q��ڶ��85ou����Fx�{�g=l��3�`!m�����2�w������u�L�����b�����,����o��kmh��eq�!q�V9^��!�(rG�
e��Q+_�C�mA�w*]ޮ���*�CV}p����x؛��7��㋑���Ƽ��L�����2��ͭ��'�+D�-�Z@LG�����j5�fg�1�{��l�ѭ�ֽW��$%��y��Ⱥ,��r���#p����N[����4�b� ��6v��r���Sh�ʺ����w���3
�:&2H~��Ř%�p�ZD�b�������a��)�K�rR����ߗY�i�5����m�VH���"�(��&/R&�jBi��T�����,u:��pK�c���q4Z�Z`���ﻑ�٢�uu�˝X�3}����/�>�.Vӄc�.����Z��ψTxJE��&E��q��L��54�2+�+<,����dE���nwOF�*i�b.�^�ힵ�h��^�l���p�)�դ5d�t3õ���<�U��\�$�&�	<��z��E�I����V8]ϯm�{�f}�\/���U�?R�M���bG��M�yU����{S^��CBA��7�\���t��'n��o�z>���Q�k�  G�k��E-�����x_c���1$����ީ�xQ�ڛ*S
o�ݡY��C{F��~�U]f�#��7s�ڎ������6C�Vu^vJ�&F|]�:�o2b�l	*�D��nb�d5�Y����J\j� ��f��'��Ĭ��R5HL©�=�1+x����\a����v+���U���:�#؋�㯪��8���]8�D���҇UU
Z�M�,�iV�,��0��R��s��w��}�La
ł��1���c���{j,��ۢ���g�lq�p��<)�p�J���x׸��.�JK!g�����sK�>�>Ǎk�������a<�R�Kh�O�+�*�,3y�bf��K����s��z%�q5f�n�H�����q"�y0��O�d*:�0�s���}�S=�O�$ı��#)w^��+�D�Eʹ�d���.ds2��̪�T�UJ�i�����9�.|�^�I�.�n��$�T�ʾ~���ފ���p��,�gEe��J���x�}�4Tp�*�g�~�Id.]��k�*8@Y�⟪
�{�����Q��x���Ғ�N�;�7e�V�s�h�k��� �=g]�kM<�	�q\��pe79`xN���￀��gD*"_s�'��qB��#L�.#��������XƬ��^���8}擩�+��~�����6Z�\�w��+�z�4P	�K��������k��	�9'�i\��2��=��a-U)�&��)#H1�ۅ�~�c�X%�r^O��,^g�KS�������fc'�~ϵbXi5й��xp�����מ%�HRn>�c�,>|��*n�n�+�׿Wv��?-4�r���>���t|�j��jg��7��iϖ���:"�VI�6����iB;ً!KۨRY�=�n㢮>��xFs�w���#r��E�SyA�no+�eo�5uuh�Π�+Vb2�B�I����}S #�V�kê�ٮ�'�]���B��X������~Zp��	?}���K�]�SK�-Q���&�r����M [���d�1tX��{�����S4	̎����"E$)�o�����xD�������p�m2$�R,̜|k����VB�\)"��<�Vܘe�)c�oLK�D���~tAm.Z���}G��s��H\�~�iی8a�燈��7f�#�߿QB��Z�dNJ�孟�E��~�)�f����X���	�Ci\M+(W������2�v>̮��h�=)t��U�ae�&9�{�괨�*^��/�.f;�k�1��`���W��F^*�Z����o����F�b�4��}���7���Y9m�������;;Ynp�]����X��-I�&��w���5_��R�-�����}��#d.i���[_>�{���Z �����}0X&����{��iVߥ{ܺ�b��]��Ke�/�����{�ߘ%~.�VNv|pKO�}�ve+�+���m�Z�>\�	U6D���خq�������
�������魥�Q	�bR\�����k� K��JD��6�LA���-f&�� ��x]}�_q|+�*�XeOii���~�=��-c�կ���}Va��-���t_sٳp�GE�OI!�RE
ۉ���x�.���.cVU֙钊�O�z�x]3������>����I�N�������8-4U̘XE�J1��|��%z�J�H�q��f�^ylU�玮Q�_�Zi?s���p��(dI�Ʌ��ژ����_��ZESCz SNĽ^�J��:j��}�5O��K�~���Q��5�+.�Q���5�3�6h�_S�ip�+�;����n�a<�f��rހ&SJ�m7��-YOD���Et�}m�GZ>b�=����K#E�s"�O��������q ��c-D�J������+-�,XaS��ť�>��t+Ɩ�ݔ�`�v���a>��vO���V��R��R-936YB���g<�X��j7d*-��W��[c�"�\��;)�
���Vw���u�п�(�89�cs`	��s�g����7�i�ݞ��n�K�k���qf3̗>��֨�����oE��V/�l��]9~�薋�*!z���{.�.z��p����D��5=����%�|!aBR+�#�`�\�|^��2�n��%DRB�����K5�uK!w\oSVxX#�"��d8�~3��5��GH_�{�ƫ��TP����?�|ZO������8F�Xb�~�>����p��q[�
��H��ߟ���:�`�À��gvU'��\�S�7_�¯M,Y��룴�et�G2�ÄI#�����V�E~��p�iB�ӏ��ɏ_Ms��g��,G�Ќ��>X����,��j�E�������A�Wڿf!�g鳋ᒻ�u���1"�x��0#��|�4�D�4�M��#\W��t�N�/s}��/���S�(���>��*�;���X�[��W�LGvz's��_ �$],Ro�.������=siM��]�O	"���ը�9���� ����G)��_��mW���)?(?ϖRJW	e����\�$)�PS\�{���:#����A�,�$Uͩb�~��pdk��b���^%��ꨡY|U��g1��{|\.���e%53|;p�y��S��4�	Y L��~�qM��a��������YW�@�j�I��'�i��`�l�3��MԆ��u4d���W�V-ە�Fl�WiwKNu%S�Y��r�-�x.̎2P�D�U
I�s�;��C��n��9��i����`Ӹ�&�Z{mA�I��l�mk�r���ǉϭ�mg�;�c�i��};�}q�yˍ��l-xfƍ[ry݊�G/GMs<!�����i5�J�o0vA�v;�C�$$�tVI��\v�y���d��Xu��n��qC�v�
�>�5Sd����Sz�e��Ⱦ}41���[���W=���g�s��:6�����s��G�B�ֺ�P���ɑL;��m��w���=������+������w�5��B�/rz)0��c�O�E�q���d1�^�V/�H���㴧=՞�G~��/<�R���y8.�������t��4�Q)��^տvK,�L,�K��t��+oA�r��V*�p]��p���	��NZ��s|�P��%�%~���8R}�����a��eN��j"��؆F�X��d�龕ݪ2Ԁ��k�ٽ<r�
�,UL!�e_� ׼�2�3UU,��&fS#���6��q��|��/�����T?{��`�}���
F�}�O}�\��'h�����3���_G�F��[Iӱ,>緅Ƈ[��+*�I�jH^�'��:uS#�L�ʙ���D�A*7�WV��s����j��Ցg ]V�Š.bqhE�>#����9��_@f㆚B��Ay~/HB�lV"�b�S\�9��϶|/�Os��H�p��0��_�M�Y�ki.��SP9i�R�	i�J�8.q��&��uu괙��=!zڣ±w�M��m4�9B�c���iY�
H�}���.��{@t�
H2��%� _}�j�����(�h�m�z���z�yH���Z�OԜ�.�%� �f:]pB�������{Zq>ۮh
�S����C0��n�)%���.��d��O���̦�+�����.0]bqgD��&ֽy�M�KH�Q�����?�q�VsVg��3�����䐾ǧH�&�h�|p���~��w�2\H��*"�*�"�{��9
�LEEe�_-�5�Z>[è����{g~3��'A�~Ao;��_�������\P:[/n��3����>��������թQ ��wI�u1���~��qf�1Mf����I"��zk}39഑�ȯ����Y͙*"���Q�* N�ޜ�*o�\�J���!p����˝{i\�yei{��}諙��/�"�:��IHL��V	`��[��һZ"��RW�5����T�	t/	�D�����Ϛz��51���)Qc@��T?zm,	��Zd��߼�䟻wt??,��n��qbYo��Qfc����;{7��3�����,�9|�����
�T�,���ϤD��Ջ�o�Ƈ8G��0�Q�2��W{���K9ͫ��L���T�X����.�
@��t֬�e��o��8t�G�_Tp�1{F�KA�gU���ƮX+�4����XF�{�@�TE42��i��{���ۘH��S������ z���a���c��R��s[�+~���h�\k���D (��L~�V�s�@R8�AO�TG-���Sq����N'�� ��)�
���Ր���G����w�Y�;$:���b�qWmofx����L�����fW4�BλR�n�˵�UTEJ(t�2�M�y�!I���b_e�d��ǉY�eICH8`P��WJ_W�V`��������H��ޛ�%ʮ�i�2���[��b�=��K�:������i$�
��@�x�����&�g�S��~�� ��%�B�}9+<��W:�N]��9�����}8H�UzhJ�y��r��1���`��Q!�L��Ȏ;�w��Ou�[,bC��-���y�N/����ԇ��x�.������y�X�bt�~޽:��W+jH�jͶ��N�b�9��6gBg|�{��{+��ÀG�W΢�B5�6���`�5¢=�w�G&f�Ug\���ߕq����+p�Z���O��st�b�v[[t�db.�!@/�fcwy��!����x�<�:V�\��e-�u��vbz֋�{�V��6����6�&RωX,�&��s��U�_��oZ�q��*��ۍ'D������D��,rPb�d�ҏ:.�z�U���m�m����w�����慍"�N_;���z_�׵�k����n<,�ۛ��ؕP�ˎcb��i��wU�Ư��̹i2������9����M��h�������������qo' �G������Jb�Q��-רN�t�·�����eNw2mY
"�O�ܸX.����>��}HWz�߬Y&��Ӄ��*X�h����TF�J���U�G��>�˯���pTo��.�xq�p���	����U���nd�ʂ��ti��&��|�n�n]�5�gy��f�ׇe⸣�y�\�ۗ�	,q�J������G�������|u+:Q|E���-_b����c�6 `�H����q�[�qɩ��L�5b�>�D������:�x��uU����E[dX�
LƩ����{^�e�z=�Ӄ�����>�]+T�T�Y.� T}mi`�c���sݬ�.������k탰�r�P�K�ϋ��������z�12����E���c�GE�`���@[�Vpb�~�+S�y�����r~}��,x�=h�#�lmU]�k"{3F��"�#q�������R)�W]>#8���KV�>z��`�ϳ2�C���/�,@�j��+8%לⴻ�Pg>~"�.}�Z�s�����e�0&���X���8�$}Y�IU	Z-M��Ɩ��j��z����w9�t����mZL�p�;ږFVL,zC���q�}y�TF�[\֙�+%X�Ͻ�k�GjtJ�x����u8<O<�X��D�ʡ�h-h�]f��$�ml�x'KɌ�s��T���*b�4�)C)���J���.�<��|y��-D�Rr%\h��w���Q�+m�AId�_/5�~]iH�B��5G������|D�b��R����~~^̫��g��� �1)#�a��VG��;��j��gE'�&}*�0�Q:�3�ھ�.)7��&(F8��*��F���աY�b-�*�Lwc�z9>�e⋝��j+�q{\�����7_��>�F���R��9e`�KWsb_���nWSn�‮_��^	k�(���ɱ�&f{4� 8F����&%
��'��'�;��f����ZL�&���tMr��V):.�n��%+��q�a��4#��b����A�2۵����je�F�!B�I߽�ipM��c�mW6|�-�K>����	��>y8�d��m.�Ɩ�~���|k�1P�,V%~N�«��՜3fWFB�Q^��y��mQ�����~��Z�]��Z�Ɠ�ƌ<iW�����{����p���>xp�%]�*�S��V����ݜ�F��mh�[]/�>��}\3;��RY|�O͂;��'!t[�[�����e���7�6�'���x>m--����N1�ooq�ʎ�d�WQf�i�8����g�ś2��r��Nu]	s�{�	K�9i3���鴾6��P�����̮	���J�Os���\|k��[�����k̕��,�^�Olp��f��ώiV�9%�M~�,���_È݁h�,��[l�ߥN4��1�b������u��$��Q<�T*�ݷ�"�ȯ�֭/Z�Q�`��"�精"꽮Ҽzv�N�m���������W�q���s�R&xe	x����y������K̙���fa��徖R#DZ�������]>�T���߳��Аw�l=��������-�K�</�m2aϟ�u����<F��\i�����FC���\=TM��{Y7wO:��uS���m6{��͝�ع��ۻ��%�'E<[X��{X�˛��'
\�7k��ڑ����{0�����Y��g���L>��\];�,�m��WW�۶d:���k�$my�Hl���m�v6�ЯLvq��{��9�펙�X�+un'��p�W��ٱ�vr���P�nݟ[F�=^;vx!�e���K[E��n^tkC�&�)�A�\�'ai��ׯߢ��i�^����Eeo�. ��]����/o�f�朘o���h�ϻP��lX+ǂXX�ɕ.}�k>1o޼}�.�g��/c�ȑ}��;Gg�x_.6Ue��Dkh��~�Ѿ����SB�տ�����[����ˎp_msUw�}�G��#���ڒ0ZG0��V��t����.[���P��I^�7���E�5��r��ߦ�H�o=�.S�^֏�[�W�<x�B��\����h%TIN�4H�D�O�$r�b�U}����ϗ:| ���\�*nP ��[�`�Z%��I���$�}ު�[A�g�e�+LFi��P���/{��з[4�;�$K
J	i��~%��X�	�V-?����j揖���)�/��s��^�0�����ӊȭu�c��Y1�.�.{ۥ��SY�#��$��r)�>�����ۅ�>�ΉJ���/�n�մͮ��A���Z�>4ܒ�<��Am�-���?���v�b�2�!:����	i�Ր��Z跜��h�q��/8��^or,�K�
�QXE,��矻k�\�m�TBhK���{VFOH�Ype	P�y���7��q@\�s�xF�����R�]����?�_���ptl�AP��aW�3pѵeN��G:����F��͔/3��,�Y�J�IkR��e��m��4���i��Y���pBƨ�GN�Ti�Q�i\���^����n���)�U��,�ۻJ���v�-<<zh�,i�����-3E��s6�lKL�BL���Ѳ��,����l6���X�J�|�,,�R���_U�"��/����
�P���D��7sle+��}�
��6*�]mb��ї.+쏱2�<����jg�}��c�Vfm˺]չݍ}�ʭ_<h��#�x�_��}{�d//��"��Ҡ�6���x��8@)*J��Jk�VSI�����U߻�u�=�O�����x:�
�xtz�;�sD������:EϥI"Tz����y��=��D�[yu�p�H��S,XI�9G����k�V���,���z��j��_S��}�K��,�ᦒm��I�8C��䳎>{�XӍ�n�S5�gw���{���4�T�*d)2j����19kH�k��o��)�Ԥ߸X?��ӛ����L]ꄔj�}]m+�V�*�sũƤz�I���޸���,X�g�e6��B�x�|U$����L���kf%k]���������|h~]���:*�T�-jڣ��Ɗɖȣm�brғ���kEm����Dq�&� �|�6�'���y.qk�̻�65������E_�׉�3��?�[��^�4*�ͅ�����S'�g�Ӵԣ�O��%�D^vl0ͽ�^|��� k���6�J��-R2����N6�v���ő�`�#�Ș�&�(?��~��t�jw.$�Q����ϕ#��.R��7��άT`#�κSM	�SU�)�gվ�\#�it�$A@D��>W������+?/\�E�����ID�E�߹���!rD���/��׌,�8hX��#�T�Nj��
�ԇZ�N�_c��	����N�\pZ-ϱ V��[���#�8���J�w��.9�u�,�密a
q�;=#���_@U�z؀n�wԯ��0�_MӅw��k��i[�/}��B���{���$Α�ʐ�|Go����U9dMC ������Pm�뿊�{��<�7�Bζv�9r,���!X�fV��qb�+���z܆8�K9Ͻa�S�{�>w:دeN&k7��˪����7{/E�1�)��7R��A�f^��I�\yX�sn:[d�F����匃Z���a�Π�y[�κIPn���(L̒��j�pD����آR��7q�oq�eZ̬�5GS��|'R��4�7������|�N�C��;��w���9b��;4T��tI�Uȋ�.����\��p�w���M2����-�����A$��H�(s44�U�O.,���-��i�}�H��j̃�����hĬ1�-�w�w�v-���T�-��j�=lr�-�GNG����1�#��t���V�$%
��6���]=�s�u�n�Z�`�Lo3�W{Ӻ��Mqr&�L�.�nd��ӫc]@����M�γN�t5o��V�C���B��"���Op��R�sj,�Sjn��e66Ew�{6�w������;�J;(���l�Ym�x\�;NRyJ[}ܟu�X[.[��
��͏iFc�i�T	�����}*ݛ{�"��&�=XL��v��T�����E����}7�7-z��^W��c$�8<E.2�-9��\gJ�cr���u���]�G�27�r�W4�� �&�}b�N�e�#,U��z�'�{�'Q!,����Wu��O�h�Z�M�J���6�:��y�ꖷ�ͥ�n�q	K��N�VJ<�wU�)�d㝺;�mj��-���VJ��p��cN*=e�{���;ٝ �Ⱦr�.n�Em�\3j��m:#���걎�A7H�Q]���}_�ւ(+��*�(��S$]�h����`�÷�:�*���^�z���RUL���_�T*1t��L9�������K%�أ���i���ਤ Tv����S���|B�f��� 7Ð-�fn$m̂���o.�)X�}ʤcL�i�U�sj�
��0 ���2�F�^��گ��R�偫\7���/H5�֙����SO�>z`����m7E@�����,o���:����q�}��yf	k	,�h�rhUF�z-��
g��+��6��@<"o`�~�EV�5���{�y�ά\L�H�AM�H�.��{�����GM�ˁS�����Y^���J�����p��<6���\���[�Zv��7��X}���\����g���TAT�M�_O
L�(���G��4�f��s��}�Έ4�M���b�<�2��;2#���İ�}1@��T�&�m�8�%)��j�#3-���VT��F��"`8�^�ʝ8 +�gU�1�_*U�eB��+��r�����L�KeE��%�ם��W�Bx��{�.�s4� 1�c����2{�wz/��zeU*�.�}P���/�8l~C �j��)��ƅ��j�caorgi����=ˋmD��!_۾���rl+�}S�O�u�cǺGL� "ڡMY�� M��MH����P�?@��,���$�����#�'"��b
���؂�����`w��,s�BAC�{z���_l��v���y3�6�<=G/��ŀW	�@��� ٚ:P��O����9-s�0���TB{�=J�L�b�uB�����k�ɳ{��y�g�۽�Dy�,����Z�8a҅bzؾ��1 �ƕ�k7�� "kj(M���u��)�3�M��ׯ�`�E!����UB�2���ej�]�LG�����ڒ��ETx�=z��mwth���k�[���u�̂_(�˽�o"wݭ�."��s@��M���y� ż����a�{=ܛ��8�'�2$��:�.���l��%]K��zF��̔�^d� E���؃Zy��|�.��e�a#
ar�%�B	l7�j�����c=��$���O�}�i��i�D0@��GN�?{U�#7�W����j��ު�8�Z{�z�O,�j�N E!�AF���a
��{�j��?t�����Y)c�7%N�SN��l����8E�v]�-�N6yuЎ1�����'�T�SS35?/	�D��z��h���X�2�H�o��.8.�8�(Wc�4v�tԙ��굈,x7�� ���'�U��E�(B�=��#o�ݞWb���_}o�!��]�0`o&��#���s��֘ f�0F��l��ݻ�pͽ~�:u�R���AYk��M��R�l)�@"�
@��J�.�<f  7��=yίK����B�ZҠX�x�^����x�rj���$�BE� �{����:0�
J��!0�S_g�_o��B�/;�v�4B0�P*p��}�*u2�*Q4��Qi�h���礤 X�mӯ{u^ Z�˙>l�0��&)�t���[=���lL�P�=�v}�V�W�st���I�?k�B�������BN��Ze����ŬU�T��PtGT���)��J����,�\��,�Ko�~�o�m��]8}|�k�����������Q���$X��qe6��j�-Ϝ؏]�tł�Q"E7�k�vd�
�}�=�ލ��H,h�r��R�ʲ��=����޶�����Y�_�8�P��R0>��4z���� 8����o�.��M0@��J{Sms��`|ؑ-� G)�rܣ\n�����N5�t���f��Dw�L*i��M4�L� �}�V� q�iD쩱 *�<�M\�G�������B�\Cm:(���������O:~k6�xn�����1P}�T���V�'�w�����K����3�����P9em��F,��VqC�Im0
�=���Q��劸�#)~n(�)��L�u�:7����Ӻ�]7&��==��l����>�6��"�l�ۗ�3�݌��7_}�#�[���9x]b��&X�˅��c��y<1��N.���<�
��j��[���k��<�;��c��%8�N����px0˺�Fў��ۋBX�G�|��Av���G���J�Y��cw6�>�s���Ͳٓ9�]۶_]�i0�{=\lW4m�'g]�ۍ��ڼ�y�Z���7UT���G��0tD��,�m^5`)��~j���!���C'��V؎5$�������ሖ�v可%?�(A��$X?�?����|��A��u�����܉�FH �{5ќl ���1|�����]�m|f6�Y�UN�6ګ�����+$��k���vU�X��<j�cG������#�3��S�sEѐ[|lG�,a�`o7p��,ゝ!���tH��� ���3�pTv]�n�OzZ����߮���~=��z�'��Q�M@M.o}�{$s"$
@Jd�.+5��
FP���LX�|��{��v�b� �ɠB
w)���縳��>�;p�𾙡p����0��t��K6���2�i�6�n�\/{��"�1R�n��"�����~���Ac��QJ6���mq����d��q�nk��;ߤ���:����Y���Oκ�������L�f!3>緦h�oe�"�\�S.@ۘ�H-��E�}�[��P�F����M!W[+h/I]��ų��_�8A�V�)
�P�a�@v�ק��Z��'�Ts�A���Zyɐ�2�	ӲA[����� O2��|�q�sZ�2!�I�K �+�z��rB{��o����>ⵐ޵�r��\�����@N9E��߹�y� ^�N��>5r9�2�_<"�+�V`{v������r$ZxI_9$`��V_g_�Vqj�7�d�~?Fr�$(�HHW:�vlfwX���[H��۬<���D�9-I��^��QaT�Wc�B�{����g?w�.4���85br�Ӌ��V��e����1�mY t_?s���u�XF ��:p��~�e+���Z�|7��Wk�F�dh��R��x` �}�i���p��>R�z����ߚ9�s�v8Oͨ�����㠼غ�eMd� X���X+l���gs�3�4h����l��=�vQ"^�%�������)�	zp��X��X//�̥�'V�i:]P��L�EqjU�ׁ�TS�_������V.�ʴU�Y� 8�&�S/=?1��S�������2�ƨE��{7����j}��^h��6��7�͛����N�л�υ�\��� ;�$�T��J&�ff��I���E��q�lH�R�J=;�W�#�>��T0_��|`-����b��:��id���iL��}��7�x^%	}��V��Z& �~mP"�g5��XSf}{�X��"��dJ��+�!7��o{�:�C���W���{d�(�U+�޵��x���>��+������i�,R"!8�̧"���W�&=�"�2�����"]��P���o���
G�|�o�^N~z?z�k���&�v�ύ�th�
�&�����iM���9�m�ȥ���4q.G	(\�y[@�RN�>�+XAƃl�������|�����_����7j�g�Ϯ奄��ʤ��Pc�:�f��uZ����@�[�Ԋ�/��� M{:^A��L/[�^J1��������Qx
�W�-����^���k��x�O+6����j�Gn�Xݸ^�jn������n�~����e�Y/�'h�sY>�w�ňZ��B-�j�0��������t�ƺG1����$��V%گ���QN�J��KŞ���a�1}녔suZ�����4ǔ�"]�Y���g?#�b�����7$��}:���x��%��\T����[�K�+�ｵw�_�+��1���/��_w~3�� "X'�*m� V��}���8u���K�����0RP��n�Y�ﶩH^w��mov;B��~>"x�!�3G��r��C��fk^���Jf�pXI��	7�T�����:�;-I`2>ﲕ���0���>�V���HkNړ��߶���t<�B�=݁�׺��8��H�*f�͉��	��E8Kr��P%�2��%����P�� ��գ�+G�\���<��*gE�aHK�Ԅ
i� G|{�-z����2�"�cm6���0����c"��^%�i�2P�@�r���f��+��އ��K�g��Y�,���A�o��ISr�u�����@��Q�Ő�J�e49���g0ώgf��i�y�C/�.��M�#~߸g�3�.8�hnd�"}ctqo����)�̕3T�pA�4�$���\p8ᕤȾ��Y�OI<4.�Y��X*�߷���߶ft�#���4�9iI(�
i��.ϻ���t�R(��@�J~�	��N�b�k��RJ��x�(�,^^|8��6EԠuMld;h�E�
����6���4]���::�H�n�Qm�Ac��-oǻ�߭�rc�GO�S��Ɩ��Vs��k�Fw�:��дZD���E��x��}��*V��u���R ^�������ۧ7�dl���}����K�H>�_'u��"i�DY��1�m�ّ����Jn�I�&�h�f�g�x
�.����>��'�ت��o��v/�����to^ ���Үv�Ց�}]ҡ`���N�ƞ>g�Xq���\p��h�bR��Y���{�-n��@�fٛٺ���*�]�m}?LtV+@/O-k�;]��#*R����f�?�a��X}�sU����-h��*Ё�D<������ڇn�7=����zW�Rx�+`�oۦF��^OIm�Ⱥx���q�����G�bT�n�TĘ1z��>֮�a�lހ�2�5Hc����>5�Y%,��k��f��o�xU!y=��AMO4�
xҒ�_{٥�=�aB�e8�[�}�V��SK�L�g���E}�i���^x\O^*�x�����/�:U@U[�R�7}j���V^-m���]�*p�F;�1ҝ����&5n>��b��n��C~�^3�YV��	�z�**&`�;9�\���>N��)#��f����ًZ/�~8E�����%�n��Z4H��i3��lj�Tr�罠^��ϵ��$G�d¢%��ǅ4�������V.-!M?��	?�%�9�l�Xi� )�r���#�)���P�����#O�[��O��������$͵��u�������ǜC�,�	kpND�J��������bwa�i{?o6��#	>߽�YEW���8�M~��4�AB���o����Mo5Ҡ��FH�x�H��Y��\�s}����R��8kr�e���	=�gLZpщ�y�*����Ӆ��vsᄠ!��qI*ϖ���.���g����"�=��U��@ŝ7���>]\�4�|���:ab����_j<s���@vN��<)V�,V�����W��8�;���b�Д�J�>�"�C=3�#����/���Z\9���ưCS��c�Bz�?2[��J4;j��wZ�ͬ#�Y��C��:짻�$i�Be
��B������bG=��*��^�,�:�| 6ߎ�z����V��b­�w%�b��zԀ���U��:G�\���+"�խ�I�{6ϸ��AQ�N�w�ߜ�?Pw�ow40�X�,�� ��񐹭{��V,%	�bxՋ�����KSְ�΀V`��C<Q\ϸ�H~�sVa�[g�*�W1��*�9.��Ǿ�M�����[�/��
��}����Z:
4Z��kDm�H��=��o�N��;*�K+�ˏ����H����"|�$����u�u��N��I��Z+9��=��{�b����K>����-@%%�v�*
�V���U�ZpJNK���j���P�'��x�E��80�{&$TP���LV5�߽��_�����~ɣ&���u,��H���-Ǌ�k�g5�k&F��n$�cN�gc]���y�ݒ�,�2n�߉�����԰�$��f�d��c��w�W�6���L��l�/����ڋ��nW���>�g��\�Ž��{l�=�(�N�-=O��r;����o�>�KFG��B�'ͺ띺�Ϯ��z|�P�rn^���-�\�Na�<)�u�"�u�c�bi�r�6J��T�����q��դ6�yҏv��N��s�h.z�r�:9��I�n:�E��]�{u�8���ŧ�ݻ$�t��dX�Hg�lPP�zÝ��kuΡb 8Ӫ19$�,F%hIF���rhrC��x������o��爲����P,p�ӿ���,Z�����
�|�(�I����U����ȱs�)��a�}���XO<�2���� ��N8v�����U�.�.��m�.[X]5b�>'�F�<��*{)j\��.���L�m>#.�;����|G
��y�=��._��;���
HS-p�o9�ғ���8'n w=�+XԽ��e|�e��*�ck�-���]��4\�w��^�^{�5���n-�>}���A�
%�����obӍ6��̉6�k
�{p�Y�Ul�B�˥�`�c��Jt�ب>�GY4+&��fL�<\�Wͳ�3ON|[��\`�����X	s{7�
}��|���w0��s)�Y�H'�Y�P�QT2��hsKx$"��c�o���v��Q�}��κ���\pZ+"����I��|�x������ Q	��H���;�4�r!�f<"���G��7�#����_����*�
�'C>"Cs����! �R�4�+4Vu�b�evB�-`�����֯�LY
m�X�����yS��+�ed*־"����X)#�����~s�
��JRX�KGU��^Z׎�R+�FTifq��<i��n�륿+�������� uF��θ��bض�{<��k*�ݮ��d˴>��nw̕�]�Y9j�˯�5�?]Oϣ�����=7�������v���Ҝ}���ī�O�XEKT/�;vA<{V%����sy>}3��~���}�x�p� ]�s�j��[H{��n��Ct1�~縱~�m�&(Q�R[u���E�}4�Q�p�����z��S���Z.��{��j���j}Q���k���m-v�p]�����QԼh�����7X�_p��=�S�j2��oX��3p��,�s����R����O�P�X>G;r���Ku}��$��P�E���qZM�����D�I���w��%�2�宾��غ�V��������P�a]���^�\|j�,�P��@w���K��~k���3u�׍�Z�u\,�ݨVG��wJ�>�f;�ꮸ\!_+�w/��Q	�"�!����<\.�9֤�W)`��o����[��K
tUߏ�������"Ol6�n������(�p{9�ߪp��'�J#{�U��5���o�v�T>a{q%�05�d*3�"y��xX��z�a�4���u�n��2���y�!g=����\��s���
�Y?|��̊_��jSm�+�5�ɛ0����R^ưY�����W���PU�*��b����~�/������|Zdw������W}�0�x_��ⴹ�.�n��W��������V*#�Y	���X,"�K>��:��9����W�EU�'%��^-�ݢ�{q�k��7&$�Z��1gF�a㛺N[���xX?8TH'��"�K����q"�9s�f^d�>����yy²�}�p�ƈ$��g��W�\s/����[�^����+�-"�~����Q�iQ�NT+!��Ybds���96�IM�4:���,4�,K���Z�p\8��}j�V��{=מ���L����#�|(�{*���Y�5�
:.uzWX)#�=ٻM����rZ�\�pg���zZ�mt��|��O��{�\<'�W���=�}m�� ���|�����飄.�,2���`��-�TYqOZ����\-!L�ü�w@�*7�x��Y�
:%=)�;n�.���,�G�7t���WsF�m6�E�\C=GU�*-�$���AlskLf�K���>TB���?gKXPc���%�3e��I��{����C����]!���G=��L&)��B�-D��=�w�����S�bG~��p�A���҅�����½{P�����2(XN����s�~��i�
N{��L\
v�s��{�>�%ew3��}[}���Z���|�?k��eM
�F�$�>Z~:Q�-X׈�|/[�mt�Z'�N��V%�$�����'�|i�f�9����0E���Bv�S�O���X���)'딭�,^#2~�md̯)"�L�t����7�{�}��������qP���gK�lI�\q:끲�>�g��/n�\$^�񝺺��d��8�?���<[�{����<P��-��ν���_�M�Ȯ�c�`�_�u��"��* !3�j�����$wnQ]<%F�_	�M0�{��_7-��p��c����SDc���}\�k嶆4=pM5^�h0R,����_+K��W��.��O�]^>���c,���v�b��L*8+�J��.�g*S��zZ_|�3��;ǒ��LTB��'���{,�����5�#�g�i*!��x��U*�4��9�����T%��%$wZy�=���f��8�1�H�*ی�K��KI"{q��*�{t]AD���r������*���/�w�X�4H��]#1௭1+*w˔��� �N��(uO��B�p��.|w�?W��ł�ə�w��a����/&aY�����֧�
Ĭ�/|%�\�r��iQ�p�J���'_M�~�M�F80�8�5�'�m15�e���Z�ҥ:έ2�ё�D�1�J��2[X���8��݀�����Tǽv�!I	��H���?l���JU*nhuF%���5b�{ψTP�^0�ޗ
����p��r���5O=��V����ۗ�t�'n�QB�;��"�뺴�τ*1ԥB_qغ +>��_6���E|��\!բ/=��1�O9����CC
6����8&�rg�`ی*ǅ�s��2�r`u	�oE�����G��H�MH�X��c�+�r�$I{쯄��9�r�!�{T�E���Wj��
���Y;|���e��]���u����\#��z+#���Z�cq�.��T.�3@��m׷G?��#��#-�ˏ�4����-�K̿��������@%��2abA���d,$�Hľn�uUD}_U����J��D/{ٖ��!:���>�����%��VBj��S�u*���S��Ϻ�5��~�,���=���t_K��$!�S��b�W�>!Yʫ�ݿ�j*5p����w-)]|!Q�iQdd��X�;K�pSM}��j���g:y[���UPZ�����E	I��w�n�����Ր�.�"L��Qu��.�r��������Yzw��Ѻ����EQ��5��}d`��:�.�!b��T�	Q*ݮ��㱥~Q�%[�q�kμ��ONd/��v�`��4	}YP�D%W]h�C��]�ʖq��_	�B`-��֔�K "��&�����ҵ.�)��&B��	(�Q�aBJ"Du
Q�#�B��D(�p�%
"?�P����P����$�!DG�
Q�#��BJ"D�(IDB���$�!DG�
Q�#�P���$�!DFDD$�I$
DB�Q�(IDB���$�!DG�
Q�#�JQ�#��	(�Q�B��D(��(IDB���1AY&SYS?��Q�ـpP��3'� b8���T�
�4���� UR���PP$PU(U�㥲&����i�
����.�QI"�AB��  �              
Q@�@                   }��i��y��;m�lk�y��/,�i�X����x���Zu�r� =�Y 2����h�^X��{��^g]
(�n��@S���� �tt[
nX�y�b�o;��^��
)�   y�      ް {        P 7 �Mas����o8==14na��ڣ�f��h��Wf�x =�lkM��@��w)�z:�y��ҽjs+w�u�[��P�@*��  Q�    C�4(���B�sJ�LA��e��t�l7 �*�ri��s:Nڠ�˻E�nn�0%� �:KZ��蓣�;9E   �.[�f�+b�7`�l�p ;���nV�v�5�ss�YZ9��Z٥���oY�m��(��vmg���6m�r�֛�+�y�餘��w

f�ER�P�        ��i���KcV��v�LZQr�v�Xm���UZMi[��#��\��`ٶ,q�E:��[���k�9�mm�J� �;a�n6v04�)BP�$�8���6e�nnR�� wY���wq�(�;�"�sc�mA4��R(�V vS[nY"�fܸu�61�ƹ��&���-eR$*T+@�'         ��Y�۶��Zknc���u�-�v���\ ��nnB��Us����k9۶��$77;+m�K� ���9��!ɣ���HH��W[fE�r�V��p ;�-m�52�۶�UM.csR��r�T� NZq��kn\;fZ��d����nd�сT�R���    P
P
 \��kn]�Unn��B�q����7-a� �u���Õ�Ͳ�t��J�v����iER\ 7m����H�69�m�A!@ �5N,����g=� �� z�Řm��]��T�ⶰ�q��c(���Tp j�ۤE��V�F�8��T\N�&��O�*U@ "�0IJSP 4`S��B����  j��H�@  Ob�RzME  &�ԩORh	���0s7s�<E���X�T�I�U�%g#���)�[�83�O��VVa/I�H�c��:�?�	$	&�O� $�$�			� �@��II��$�$��}������_�l���^��Xfkw���sͥ{{"�X^Øn�g�{��/�Es*�i�`e�.+��ٴ�[h,��:��Ţ�` ��B|g�J�.Q>q�r�٫pQ͙mE��I㻅��	v[����B���a¯�z�����@	��<}f�ZxȤe6e�:�P��>wj��sF,�2M�-^��_%���V�*�%˛�*S)m��3^]��-��7Tb�wa�ܨle8�ɴ�CU����ؒ䬔��:[��{Bd��L�,1X��Z��(�
7Yh4��F�/�1��$��a���]�q4T��H�]Ա�ո��jĈ������ǫ�6d�7f���dσ���!���j�;Y���j��Z�Z��7��I��zko6��V��.��D6��޲�c.`�7�	+���Q�*V	b�QZ�$�g.�;b5X7�#e 2����u��V9����DO��횫Â�Ǻ+nm2fD��bϱ�4�V[8��Tp��*�r%������n}6�s0L׀�x� l,��hL��4oÂc)��6������Q���Y�fMk`�8�f��FFe�R��EcM�sW\���z�N��({f�J�2o��K� <�+�,�U·ʫx����W�l;��)h�W�u�-���i4����+�fn=Dn� �����LwSެI���E^��)U�&Ʉ�"��ꢱ�>�F�* L���"�PI<��vPe�W����xh�3a�@('y [�f���S�E���a�»O���F�CX��^�X=B�d����/&;F�V�6�̲m�`˵փ���� ����9��Jx�Kk'�g���טJ}eD=@�0zX��h�y2�Kson�_M����cM�&-6ܽ�Z1Tuܧ��B"Z�c-���1X�Z�1e���YT%fW�~����GenR[x6�r���ŸHܺ ��S�Nֈ&��z�љ���7�e*�sV(�	1b�4��N���vmd�+1
�Ga����z�0��Z�4V���Fc{V�L�b�����ǐ߇��
�"�y`�IfG
H�52�3�,��
V�qz�A��,��q�V*y��e]���Ē�*ʁ՚k@��CH���q"�A�=S�/{�W�`��h�1�Y
�Z�ƅfTYvl|
f�F�ݛ1	J��ay^�&[��2�u���0�v��1i�B�ˋҩ�kZ�]eɏn�ڶ����5��7�TY��1�V�љ��X��ժ�qt��Lͦ����M"�ᵧov���H�[��L *\Ȯҭ;�cݻ�e���<�"º� S۵l-�*�;�kP��S֘��������Z���o�Yv	�L�9W����@�i��� V�J^2��Z ����t��\{�ԋ@�ps��Z����7����M�1��2+%m�E�wc�Cn^��\�	̽��@��²��B9/̚
N��ə�)楊H�C���^,��Y�@�HM*9!��*�R9[�kjd���\�˫�~�Q7������	�-"0��\�v��74:�HVv���Va_8��������X����J�"l`�;+F���y6�֔(��QBs��ɬ�5�^�M�U�.�I�a;�"3]m��r3���j�Elxc�5�d5,�qM��4�pi�{n]��MS.f�[)��V��=��v7�Őq 2��kL�Y��yJ�ښN�! �3G)!L3l<8�&~����n��J�z�Qm�:P5~�Ux�6���Ҽ�dm6^iٙNݏ]55'3#�/u��Y���@9@�Y�BT�H/��*3P*�)����S���(Յ�E�y����׎3ɀ���bZ�"��j-P<Vm��zЇ��X�J���4g�2��u����aՕ�n������/��]�eMЮ7��n���y�i4�&;�
u���e��Z�ꑊ�V�a�=uON�
���jM��K��z�7��$�{�{!Jαo.��e�(�:`��0�Y��޾���ͭ�أ��3WB#�������׼0J��hbt�:���ӻ���Ż��#Pˬsv�c"x��l�}Wr�9m27OLn�j�R�p�}XoF�LVlcNK��r���0k�{֛�����Z^Ʉ�F�SrK���wEzGa�^���S(�����E�.COv��7� ramC/KŖؕ� @-i��n����Ղ�"��Toj�ʗP)j܅��J�a���6ފ�ْ<��Βހ�-B���l��{I�T�b�%�Cʡ?+l�>�=k��l/`iU�e)(0��*Z�,uP:�*�v+�f��Sy%栈fE/n��gmAW�2�֡��S��ի�Ѹ��1
���k��(�e�Q�/-��Qҵ^U��g�x���iP�y~f} �Kq�>��d��F��~��"��v	4���$��*4⼇ J�c�ȊU�)�)���{��ݸ���E4��bL�XbY675[6��5u�x͋.�W�2��I���z��,�<
�o�H�V8�d�3D�&�����Ŷ�
��i�i��{���$`�a�ZW6�D���6s2��-f��$.��Ki��3,��%`�H�˺GS4M]�sE�
�In�șN��j�!�����N�+ez�5s�:�|��	+r��K�YEު
�ҽ;�k�2/(-���"h�v�4����x�������lz9S�V2z�4F������y�^�R��WtԠN��5�+k�7qre]�ϡ�)��%ф�K͆�r�^f�̗N��%Zvλnj�e�`�JJS�9X��	ڦ�K��w��U�t+/ �/ln˼�K[I:�hR6&� ��PX����Cp��6%س&���
�����6��D�X�ts'�"P���g�t�CJ啄�^�Z�3m��z�ܛysR���s%2@����9�ٙ���a�r+������:�Ŷ~����.b���C�2�mF�9K�"U	�sb�2�	��
6v�R���`���7t��NCD��#��)���σ�hZ��I�Z�9���雯*T�1��i9R�f��	�x����f��&�8.�l����=�=ճ$�1�:m�Os�֐��Wd�J��P���57vQR����fe�WG	^�b��U�W���V�K�݁T��0����Sɥ2�bf^�kfL�;�)8�(�n��vf!�^��@�+�X2��j*יF������iKZ����Uդ.�̀�w��Fj�\�c笐M�h���7�w!?Eh���S��h�|<.�3�Em���0I���Ax+EջL;��5�v���C�CW�~��8�f�3>���cp]{&J�U��i7/D�cϘ'��WWt�
f�T�S]�ܙWNn�Pn��l��K=Ye�F����%V�n�� X2M5t���A�y��'(Y1`�Q{�f|��t�˃5�!X�����m���R
���ԇYbz�h��#��d�9�."�V�� V//+k]dYSV3~eˋ1�2m����fPH�'�ϯ��-}jL̎/!�,b������} ���7X�)��ʓ7rA���yw���1Q���ST�ѥ�����Z�l�ԩ�ݠ2.�+slj�ۗ�*,cq��ԃ��(�Yh������ף$�#��y�Ze�`�'L��9��z�82�+���Eh�Y�yv�?W�X����|,�B�G>�r}u>I8؆V�[�lC_Tr����2W���|�lB�����ڜ�wb����2޴�9�2w-�����r��S�p,U/ໞj;���SO2ug9P^f�ݝy�C�L��]n_Hk+.����e�������{픚%�{�x����Rt�-5,	�c���>�ᯫwUoݲՓT��9���U�R���ެD�Uiϫ^Ug�#�U!T��醪a���t�g�j&�7tɧ�L�;�Ú1Z���hWE��
���㢹;�W�R�4�1�{]�PeV�ߦ��}�\+�%��/"Ҽ�hi���;�����ȴ��^p֚|��.�qK�U�ge]*����L��o4}�jՁtob�v%�o`�y�oXƴʔE*f��w�)+r����A*X���F��ʎ�#hl�ҫ)f��2��WXմ&�0�d�ڹ��b6�d�*����W.�=L�)r���.�[�G�*Ȼ��vs�2�N���B��D��P$A��w.�k+v]��)�a�ՃS
�*�c��%e�w�o�ZW&=�7�
62�4X�F�9N5f��O��57,�)��xI"�-z�t�(�S�T�0A��S�Y��$�*�&Ƅ��5*P�֪4��ݡkn�ʸ�I��LG�7�;X"R���e��]ɹR���1�,.�S���e�7���Rb���ܴۆ
�ʆ�իGYL���:�TB�^Q�2����x����!bT
��5��n5!�<.�K���Y��ꕌ߭��#en 5���C7U7B�b���l�V���Rʖ�EW��!g������(aw���]�,�����0@��ǎ�T�a�L.!�y+�;E��Pf81Yc��J[�A�7N�ŖԹ�(�~�^Y7C�2����$z�7=�)��[�]�+5e<�СY
�Ye��f���ڙ%�7�P�E�Vl&�\�E�Q�R����5t��jd-�\�(�7��F��QKRѵ!�����M�!�e�w�d��nc�el�LώB��n�B��&�,�H�j!u��!,��*�ey��0��d"�	��]]$2)����
�����/�U5�&�h�b��WjV�A҆�:����Y�0�E+NCZ,�J�r���6HѬ3J�.�dy�EG��,��H�uZ¼���ӊiYv�ٽ%ꕰ���J̧X.�J<F|�"�tl�@��J� �!E|�@YNG�WG�j�����_�mhY[C�Z�b��]JM��{��6l2��f��Lw�����9M4e.�D]�9��%�s[]��M�2��d@"�E�ޚEM�B�W�)pS��%��"��JCB���>�J
�&�M�X��QQU.��@U�ѽ[��3�R��XׇP�r��b�o��Z�X<� H�R"�ɕ%X(�Z���Jm��F`͸.��V[`c�n\"�"�F�^���j�Z�y�"̡�X�ԭsMdwOk�s���kغ��>�����mC7w��XwJ��c/��,��׋J��T��F���N�5��5�%����,
�EJ�ӷn��!�mD���4'gi7*V'�mYl�qFhn�QV`��N�""��*�P���t� I�u��J�d�T���֢�&��?f�8���	[���];S�4����u��c�!T�Hٕ��*��C~5,�0#c���P9��g=����;G����tV}Ӻ�����D�����c���T��峽��9-Z�\����g�8�}�����JW�����o�F��۫ţ|<&�:맕�׹}�( �Ȱ���
�CfݡV R�ù0�N�TP'�򥅏Ve�E�����&
F�:�A�`;���[��Ө�N�h)2@��Z��rc̏6ֻ���Q�ٽ�;d��r��Z��mQ��V���nV��^�v"G*R���(�������ӥ�¾�qY��t��ů��$;h���ନ�],"Ťr���6e(�{Ef�&�B��)�K�\�*H�g��z�I��EKm��]�8�/6�����6]?:@]E[d���^��]�bŜb6;sWj:�&ޛw�`���FZf�'n�G��F�F	Y�rД��z3d����7(��:�����n�b~�dx�@g��j���uMs(�6���QE���ỳr�����L��N�Z4�H�U�mj��B?*�Ek�p^���н��b�^bi*.d��rT������y{0���t�/@��e�z��D!�k kh\�d��������F-�Rk9݅f�.�ʚ��6V;-�N��M��2Ħ]�t.g��4b~�M<���b�����7tM��]�<�*,�2T&�;f�G��\�L���.j�I�ޟ�d �}՗ْj��iU�͉��jN��&)r�Xf]�~YQ�`6�5��Z�Gz��u(jۭ�.ACQ�f�׮��[���0$C�8�:��ѴU�DU�Ewn��J+�M�-��*�z��KR3t�2�(�	5C�!�� H��tX�H�jFn����Z�J�p��jM��v�B�h�t�P�O�%����J���&�F:�k�)S�v-�h�K]�*�k1���ڬ�oKK/,K�(Q�c�oװ\��h�p��L�j�r*�8(�}��֦[;tu��%߭:�L��h��ިZ��d�[6�;ǩf4� n*&�Yj��v�h��5t��F,ѥ��%�4S;t��om=��cu�y#l
�B��Oi��{�'�1�|b���#C�b�&�;f�d���m��V��6�3rZm<tB��EÌ��[���F�q����p��7][&����ٲ�h�0utN�=�VȭF#
4٬5d`���Sյ��B��2n�j�mY��n�97i�f���>���3EΛ�u��k�ާC2m����2�TjRʴ]+^f�V�x^��5��Q��ɖ_Gx��6��Z:����֍�8�xN�A��WQ���Ւ��6N������j[R��
���bbbn-Ɓ�wD�e�̈q*+V-�V���b���VRUjf��fԐ�g�*6ʚ/*�t	P	u�n��1����n����3A"�Yр'�R��[Woz��Ը��ykl^��-�͌|����.Ƥ�r�ʫ� ãk ] ��t#����M$�R�J���UU:,� r�UJ�*�^-*��įb�vQ��Z�(8�]� 'F�S5*�ASwT7Q*�PW�A�u�jz�vtU���@�U�0T�ETUV�һ*�UY��a���rxz�i��v�'6x�:�c��L��\�ۋ��Ee�ú��Z=�nބܺ�mn��I����q��9�\���:�4Z�3��׆��`
��Z��Kڶ{cDJ-���<A�n-�󰸲����Ch���l���h��AѪ���ܛ���������Y{(�����<83� )�+ɵ����]98�Abw<9��?&)2U"�5H"J�7���7[۶�7]�d�qQ�"*^� ���ӌ�xmɭ:������N-�N�v5ƅ��jM�ˊ�#�e�7�v�gg����Xv�B���!W.��<���d;ۢxh�������,4wm���M��j�����]�t�cx.��ٓ�'1�&�ln��ݎ�.���ݹ��ݵq���e�^�Wi�:�d݃F^�!����c�8�C���a�)�tP��7+�"��L"n�ٻ�� $�TJx�k�j��mҼ��v��y ֽ���g��E��*��9혲������c��Սʈ��=0�햰�<�XN�5�面w$�L�y^�]=���;ힼ�ݍ���<5��c֥�YyW��v�G`cҹ�S,A�� ����F:G�gjH��Ըz����VNU��b�m]=Ypn��{u��fca���<��v�7s�z�]�4�KAm#�]��{l-�ms��d�E��G;���3��\��M�X�8�N]���3�-�5���t9ح=6<���D�Gl{U�;b�;����tj��v9g��q�������8ɮ㌽ո^6Φ.9p[y��ax���
$vݩvn^�8��&��n��\cX��Q���f� ����� T'/n�':k�����,���}�y�8�5#a�w;�5��P��w�5�le�X<���۝m��͸ktvku�[��GH��=��y̼4vB;jw��<u�w����)u��V�\�7���m"�鵸޺�.�ts��g*�f�q���&�&�q��d�6��x;=�Lv�4P�Vzi��4�[mْ|���=ӻ]pF[!���c�ȅ��H]���m�MSa��+���=��a+S��� ɷ/��������ŭv�O(�\c����<�\�.9�����6�<cy��<�==�S� �0�쓍<h\��o��/1>�� hv�<p���Qͫv�]7�����
:�wan�r���Ɲ��j�];��{)���n�;�����s���j���ZC/�9�Fǐ����Hrm6��u�ٍ����7eSg�6۴�0�f�ڸ7I��Y,[���pY��퉛��5����]�<�E9��O�&�&f�v����EQ�KH;��/�V���%�1�1�8����G9ݧk�� �g@�sn��!9�)�����mW\�m���(�r��b��d`�������ݰ���!�q�|nPs�xs\󞇞ݷ��[u����9�u�r[��5��m㱺ܸ�nwX܎Wn����u�������uŃGg��i�aX��\Q�m�O@)��l�nL9Ű'a�,�b��ўs�a��=�9��x�L�d��{p��f�#���n��ŷ1e���F�7����ۣ3�OD���Y�#v���]��W\v���f���#��۶�h�j��Q����n�8�1Ӆݞχ�/j6��u�r�'��;���1�{�3����+شk<���^=��Nv�l�k�;Z�)8x�t�+h�xz�9:���M���\s������ESMZ������7`\���ڦ�v�)��;T��-��;m�q�'����;WMv�"n7[��9����}�]Z��ݜ��y�}=�����v{	�s���mG[^���:z�Cۈ�� j\��Vc�(�=ϓ6�q��������:�9w/�',�;C��9��@-�n�oZ�Aŧl��Gd����*�Z�9���ct��Az�<03��O<Bt[��;(�۩�|5�=F��nݫn�]Л��5��C�mm����nSc:��!۰<\M�,�ݰP��׬Kn�vWn:�g1�i�z8*��>�m���h��x�d�p9��RqF-��st˭�K���s��lv-ػUntGn���1Ψ�����f|�úc�u���*�WgvM�Qۯtu�F����p����i\#������p����(W\��wI�=�����Xv�{C�ܚ1t+�^�<��l�]q�-նNi��7��z��uU#�ϧ��0���F���#��ع��N��g1=��:�l3�ocr�I	[�[��c�ۯGc�ٸNz��cm���\f0��I���$sׯm<P�朽׷^N�6+n���9��v�ّ��t[���1��"�7E]�r���h��ds�v�z�z:a��vO��*<�>����n͢q��ݧ����o0�({]�C��kB��۬��׷1q�@v�mln��	���rt�o������d��u2\��.�8��vX�ۡ�<>�co(��5�]n��a緇����v��/F
��<�v�ET]�����R=m����nҥ�[]:�ճ�ۛ��ݽ�m!�F�@�g��'ۙ��qnP�y:���y<m8��Slv�;;ͭ�����Ի��)m�8�����-��C!Y� �\�Z��غz��#�����pvp�=ǃ�9ێ���5P���[�4ՓFD�
�W�.��r@oA �R;������7���7[8���peс�W��u�\��Ŏ�9�l�L��j׶@$uV+i`�&ېD���f}�[6�ڛ}]�7AӞ �b���t.�9�h7k����R���F�ǘ��%1��$|�a�&�㾾v��];u;��N�ݐ{ggn����=�X��m�[r��Q�A�	�z��9~l�%x�"�e*d-V0(�+Z�"v�v���\m��᝞nմ��cj�95q�g��]=�=�����&6Ƴ�n<�'�����m�m��.Wn�R�׎�����Sn�����g!���֮�h4��ܻ��묜�tk����GY���rɻdڜ��� �I���L�lZ�̍�r�t[�7l���r�=�����\�6��>kѫ~�sۮ3��$��c�d/k�m��T@�mD�
�U��6�ӓ��hڶŷ�	c^=);�#���mYn{Qc>9,��8�c�e,>�Ԧ�Oj���k=nFc�3�s���M�O$�9#�8}A��y�^��쵣W.
}8��O�
�X]�˯B�nl�*vݝ�t��ٟft�õ�즪�[Ӻ�]H"�}8��q�\:4`��ł禝ʍ��1u-s\;����Z�Js�Z���N�*�#N�s�oe^�al�-�u6��Tc�U7Gv�|�#���*idS���C��*p����$-�h[p �;n��]��E�[�5�^�=�N9k�����;c��D��N�-� ��{i��X�3׮�S=�B6ckD�2[f<�d����.뭣���c�ӝ��:9�u�\�b�;l.%�7i�.ϭ̙D���u������,.��<������;#>���{�ݮv��8�6�:5ә��!S�T�ֹ�lwI�����6v�wn}�ǂ^8뵃�!m�˶Ğm���LZV��9�
���j��Z���۬M7>x�Q�W�5'=�ݲ�u�ׯ0����yw@Øո䝹���y�:�9��͜��g���^����^8J)�F\������苮ҷI+����]��:�����sZ�M�8렇��g�9�'2���Ӡ;:y��K�m�L�txƵ�Y������d�7Y��9�U��Ni������볺*F�s"Ca쉖g�sH�'vZC�f{wg��Ɏ��"�v�ף� Pv��p��OcU��c�b�]�[ǃu�:��(9��x�=ur��m�7]�vs�<�Nw[K����ڗێ��<��v{'q�)�	C����� �\��ڗ]3X��\��y��s��^'st��]��9,]�[/)6���7[��Wgn�$s�2k�R#����)'u99#j���[�zmv�6�<%ft��ls�����$r=U+��]�Q�m��Q�ݭف5�
nD�[�V3��E�m�ݰ�xw:�^/���aOP���)����$�.6u��s�pq˶�x�O���>�A�q��n�4�y]n��Ú�UZ��x,u��bɌÛz�^ݲ6�o-�[����{���,\ul�vN���:_r��!��������9�G�c7`�'���t.i�C�N^b��Z�`ݜ/��1�],�c��=rF;=/U�=���Wj���g=;���8�ݎ 8��������nc-�����Ӵs�Q]��;���tKؘ������X3��ԛs���8γ݀�v�ԗl�0�Anu�@�۠�l#��\��Y��o��IׯoC���n�g/n,X�磢}�]�ق	���&z蹏��npݽ�և"Uv���8ji�W��7FםP�b�/;�Z��S���y���v3�	�>z�<bў[��&�:7��2q�;(�ۂ���G\�<;�ێ�Wk�V��7d�SWm�ޟjv�6�F����f�m�]���yK��Ѷ紙S�P����}��ǭH�7�`H,+���9�m;_��|N1��8W�A���ٻ;&�f^�v�����������g�Ճ,�k�n]�V����7�m���r�wY�\�]H*���4��wQ�\��؛�Og���?;��t��=`��{f�f�V3��m۶�Hu��tf��nЈr������:9��[��\npr��� �Gh�șϵ�,���]�Q�scv���듢��m�M�q��r qe_��z�֑�v�s����q,����rv�.xӒ]����˴�ƌ-����$���!!O� �@�0��@;��?���K�╶�㖺�7[���u�sUJ��x=�9묙Q�]�1Ύ.װ��npc�Y^�v{l�Ѹ-�����s��Q�����M���͜�ݚ8�z��w\�v�����fq�.�ur�`�۴�a�6ZW&bƮ���[����[7$�[�y�s�Gp�6����v/n���q}v8۵�3�Ѱ�Nx8�k�;S;�i)l\�|oAZ��"�d9�����t��]=A�m���2��{t1�ۗh{l��덫�Z�t��1�s��.�A�%c�����ugru�=\q��j���\�ڶ�v8̮v�16'l;'&Ɏ.���v��;k����vO]�na��I�<����4oe #���i'��);;�)�vvwqj.]�NY*������۲3�#�M�zx�h��v���ci��Ѱ��-�'��n���;'C��K�r���Ls;^����[��x�Zn��x�"h6�[q����YN�m����Z�:(�/m��k:%���'1�F�kc��8��Qۜ:Sus��}x���Y�Ӻ&l������
b�pYۃ�ezR�����φ��B!뭲�;s������}�!��v۬��Nv��P�o��ti�n�չ���n��p[�[/n�5�/=:�5�rv�>��i��\mv�t�{뎳�X�c��4q۷�6)���m�]�h�0t�:�uĬ������ȧ9�a�^18����]�Ξ��;�;�u���۶�s\�&�/Y�;���tC��lrm>y$G�#^�vq����\N�ͨK�W��(n�v�;r<>8ֳ<�uۇ�;{��A����t��3h�{�ѻh�{v�gˁSp�/� ,�G�����ͻ/Um��5��D��69��a8]�v6����-�w��].�Y���ryWS�;<�=<v6�/7m��!���s�i�Z
��ܽ��saͺ<s�#�c�n*���N�U��T��nΔ�N��]t�hrl�لA�Og��H �	@���)( I E�)������}���3�G���y4�	�Fw`��mՏ>��:����s\g����L��a��N7\u����o6�{Y�]6�l�tc7n�n�$ˍ�1���T>w5��XGj�{{C��As�V��í���]vJ�.���	���5��ck�9�X�n�8�#�\hw���P��-��S��R�˸��sq��3SC��ow����y��n�m�����\��r��{r�ʼ�����ҚH���5�6�F3��"Io٬ON� ��.e�a��}�a'����=��{x*zq�X2d�cv��!v�������|+���i�G� �òd[����`>!ɷ\���&�=�/=���۵�8O]m�\��E�B���'�3�L[ר�I�[��ȏO�=O���x_ 9fs�`�o#Ţuf�����5���zr�5�{\���<*o��х6�"��y�ᶨ�m,G���V{T}��P�Y��N�]��m/�v'/O��X��]��ߢeK�	�����=�X��8�4��c(���DlG��bٔ*����Y�Aor}�',˖��.��4?�v�߀���i������X�j뮫f���@Dk<�J9��!��g�d9�nV��<�3	��u�Ӷ���5)��LH���!���L��%w�C�n�!Ĵ��jU0J�KkT����}��w�U4)��5��a4�3wDi��ˆ���7����S��E��y{�ĦO{�
�
{�Ί�����g��d�p��f�����2�&�8}l�K�Q�	�Uԭ��.�ޘ�h��A��A�Ƀ���Ykɾ"sOKZOD��֐��?�j����J�/�1]n���۸q��i������UKN
yN��ꈯ��,xn�N,�gmi��]m�?���Y��X;s
�k+3�t�q4��i�m���7^�٪d�jc�Y11��	������q�f�?�bG/�g8g�i(��ʘ_�ڠ�5����ε�
Kq;~�pq��:�L,Cu:��CI7�4,lPg��{��+|F���k�f��	����m�{���e׷�h-�&'��뮡���6�c�Ɋ����^;Syڮn�E���oS�]O�Q�)�m��vm�?~ǙU���"�"\k���S?0�M殿k�A��b,�WD��g�V���a��t�ٚ��㕞g�~���L�Dm�}_}S�n���Uݴץ��W��4	 |m2��F�����\u��9.ۍ�c�=�Zw<�pv�;$V�%T�R�8ZP6��nϕk�����9���u:�0ݘ���,\��>�����>�LU1_9
�~�޵�뻫Ww��+�M�n�P���z���סd��{ʹ�MU�T�m�Y�m��Xm6�[�L|�ɮ�����p9���R%�dU��<+CV�/��I��ڸq�W6��&!�(z��^�νE8�a��ޝ��r����'�ͳ�v��Y������V9�'V+�ܱ}I]]�M���j��՘Ρ̢�����ɤ�꓉�՘��e���z�������<&���{�k+Ԡ��~�jW�`	=��̫7ԷUY+p'���3�K:s�k��(\[���"��,L��u�q��G�T�X/
T~���5�>Wک+=�^��3̵z���?D��rƨ2��ɶx��Ls4AA�#��UW�X|su_�h����R�xo^̇o�LЇ>���n����v��`x�������:;ҥtW�*
����\�T� ���/�)������UU������GwGXiʘ�����Zi̢�-_���d���	op�&��{��P�Jx�0�c�[_}s�m�I��T]��sF����y
�Yl0r�g���X�-�T-`�$���>`��Vg����)ü�:��6�ǧk`ݻu���ؑФ_>D��u$:ӑ}���/N�\I�����D��m�uϮq�UC��Z-$�h2���'����uk[��I��)%�y6�ﵟT�[�N�۬�i�q�qy�l'Β"FP��\k�����˚��GdU@����團��k�p�t���a�P9}zw�Lg�P�1���	����V��ii��ciu�k4s(�g����ZF�܏�:��x��C�O5��LFdam�	B������CH/��Hx�kw�4�-�oɉI�e}�p��PS
3F�?�O0>��ٚ<�2[i)<���n�y{�����L�k����9��
80RWSm�T�~�4��X/a�PWEƼ6�>�;��6�.��:9�6��{Z�O�)��ɉ���9ۇ�Soۣi�5V�*����F�<�˴��)�K(ŴoG��bǽ@�U�[P���l��9� Fk�t�j������Me{݋mSY�'<3,�p�{{�0�������C��_WZ���v�p��wR��]& 7ﾽ �{�PӚ���ɧ;�K~��J�_$��D�:��}�����e=��ʴ����v�j��:èy-�`w�p�9Y��Sel(�	��%LOX'ez��=v�&^w"Y�Z琟h��Fۊm)"r���v�_����m�'�Ry��|�n�d�W�I�q��!z�ݭj�
�"�>CL�Ӧi����z���ż�/6ɈS)���7�5���䏷u��F0��WB��ZL2�2�!�Vӣ�)����(�2!uęY�Ɋ�(`���.4����ٻ�����ߨ�M3J߽�f��6���wjbe�޴�?_�Rm�>f�{�e���i���+��˻[�$��i�)۷�﹭T��{���SbS���i��Rw_{ש��9dU;�m�+�5k��ӳu�NȐR��ٳ$�
C��w�;++�>ʗ��WP:�Wq6��:*@j�e)~C�����CO+���u�q�����l��!�<�:JO#��'��9�H[1{,���R�G���L|G�z�呫p����ܣl֫}�[�ʠ�a��۶M=���R@���0T�&wS�����?��Z}x�Ï��8��d�6���'���YZ����[L�뵩����i<Ic���������ꤝB�4����］�X����h���5�Rp��$^�J�[�iP����VvV�c^ �]]���o0,w���[�Ӯ6�%�/R�N��,ۼ�3�I,D�Ԛ��-'�ݶ�@�3g�%v�6��;�90���{<V�Wu�Ǯ'v��ݽn�ۧP+l���q�F�J]Ѭ�W���t��v�V���7L�u�k m�Cu���)u�vv�����q�.v㮓�)��v�Z:�裂��}�mv�y�e�ÈW�����]5��۶G-s�3���(�va.�H�=�x��G6����.h7:��xLW/D�� <w�\�x�*�.�h�U�����j���;�k�1IP��_������!��ǉ��9��W�f���c_Qi�ݘ�#�^Ӌ�^%!�/���UX�˻��ks��k��m�ª���Zg&��d1�}D̩���O��ٜS�C,�UX
�����kR(���V�����ic^�Lk�t��3|��k�{4E"��uE���;�g=g��>q�ej�޽`W���X��o�@zW[e>k�)��_Қ�W���c��=y�N��7�뷾���8�N�����ь���3U�����b�6ȫ>�}}�@�S��u�����n�ϙ�m8�yS{�p���4{�woZ�i�)��_'�-�B�y��k����f���:�yU�{�Ȧ�8�.�-;�>r3{����I�ڪ������`����/���R���+�����S&V1���!T_��`�N&�
���d�ĞLa��.�u��9uS2�	�i8�n��CL�3^�32n�/PY)9�j���y�m����d��F�m�B���f���éF�-%������Q�����U��S���.���w�lճRX�b�t�f�#;(<�v����'��lt��l��=����q��?�ʡ@SJ�%�Kw�6�w��M�)��_��o�(u-�>��}S��=�p�*c֍Y�9���o'���0�<�Y��Ͻ���{�\>N'�:�>�}��!�P�����=�߼탊��!�k^�{���Zk��w���Z
�z�g���̷�����Ȭ�Y�ދ>*�͕�[�l]"K����h>sd�o�ۣ�v���\E&_�Èm���n%eCwS���;z6�8�W*�oU�kצq:���W����y���V[6������݈n��>�_G74N4���RcJ'=�a6�w��LJ�IZ�v�W�^���X��ji�|��L�U� � >B��z�>�}��w]יY@Z6�W�^�̹l�,8�S2��~���׽^�j����H�����	N{{QC^k���|�����<�x��b�'\L�����r��h�ste,�3ڽN��I��',��6&o�w\�Z|�N��ȧ^�w�4�o._�*J��b~R)_,��e����Xv�;U�T㶳�
k������ɘ%E�k���a��'45��j���Ri'r���6�r��X(�S�y֬3T���g��f�Ki���M�j?�Q�eyբy�+��*�H�nYga�G%Ƈ��mc�b.�G�R:��A��cQ��"����l�B��_m����}k᢯�z�m';SZ����Rs}�Kkܳh�oZ��6���sty�P�}�ާ��g;F���\�́�l>�k�m�}t��k�RV�w'�N�:'�r�-�U��m"��HZsUϾ��~~Mnך�͟�Z�܁wR�,�^�Z�'j�8��m�(�p���mu��]d�ɧ{Č�ݹ��+�����Kp֕uƆ�ݛ�ĕY�~��3I�i-++��u�g���u�꩷YGɕD���ײ��i��5�ӝ����1��~2�ۅ4�Դ�`���.��2�o�V�!˪Y)�JŖ�I.�{9ܽF��{8]ΰz�/j�և{fצ�D�U=�U�U~���W��&<f!�Pp�������v��e��6�>�����_~�Y������U��m��6��ϷZ�99�^�
CO����O�0��z�⢆%�������3����)���Cl������4�s��~��wL?p���U�4���V�����8�MՊ�+v�~k����C�#_)�!�7�������OW��M�^�;��U�r���4���q�C�=�kW���Rc젶
u��k��Jf�S9tO0�i2���%���K[��ZW(���=�:.y��ۜGwU����ⷷn7<ǃԧ
�/*�/���UѤ�y�޲q֪�$��v�g��޽b|��lY�ت��8��E��x�V��s����Y�.��)cY��4ZM
�o.�m}�ȫ��=�Ԣ�+V �n������u^����k{�j�����c�In�n���T�8���sg^2��t�w]��)����m�������%��P�՛���K�[3�;���⣩XE %��*��5��U��ןsVM���P�4ΰS��^����pI�o��v�Y�}��Y����rv���{�]Z3���E2m-�B���e�ksI�mLU8�c�{��
S��g���eka�S.�z�=��)���}M���AI��c��r���}�{<x�M�Q�{^��A�jo�)�������<�襑Î&]�Z��vC//�Cକw���.4F��Ng=U-l]ӗ�Z�vŎ:��94�o)-�tVS��Tû��Ůn�cU�O�߯�S�+R��A������ɦ��bCI����:2��^�?o5�^Oky�����O�����H{����;κޭ�*�C�i;�ϯEv��>��4�}Mݺ�K4⛗溦��ZhB�c	�O`]{/��۳e�u����ؓ]�э��g;���(K�k�۟������[)��=׽����0d�4#�{u-<����M��bC/��{�o>o��V���j��8�|�C��o_\�ް�Hk�7�v}�2�1JX|T������/�����c��{����D4�Wu\1��-M�{�<� wG͖2q��n�Mv�>L�nu�����=���gx_;�����ZN���2�*��q��/*y)�ԦJi+�@G�^u>`��I�!i-8����i�|���?S�ֵ�Z>N���w6jC�_]W�b��thf�Z�{&3����4��+i�L���-��l�NEY��m�������9W����>��r�a��v��gP�y��P��Y�4�~���n���6�n�M�LW����~����M@|�zI1�S�ìO�A����/����
�Z� 1�	Qd�_���&��(�h��'�~{a�-�����z4u'U��B�ùv����W7��(�a���M�n$�~t��17[�&�W���X ���o�Uz����u�1��u��Ǣ�!�XC�5���������7V;6�;�s]�`��vM��CڪK�Oi�t>��=�7ś�Yy��$��*�(D��[k�� �^/n���:4v�ͺܻct�b��!�)�{�=��bx��;	xai���z�9��\�x|\���ϯE��i{t��o/��=o3�-�������n�>��]���9�|n��<�^��]1�lc��6�ۓ6�N�g��>�O:]��1�U���0ݣ�Z-�/E�[L.��v�ml����5uH�!ȯK�,�#c�y&�j��<^��)���9����h�ϯ��n�׮�V[�����-?s��!��ZՓ���:�Z�ɤ�=���P�
L����s@wU[^�m���ɽ�6_;]{̩�m�M&}�pѾP���i�|�*�a�9����יt�*�'�ki�����3���@n�g��Z�u��5ThM'��Vo�R�fXu6��Rq��k�
�H�S!L;ܿ��Ӵ9u�7^n�.����K���
�-ը�
Ϻ��t�\k�8���=�)�1�)���	��j��6�'3yU�i��{3�1f޿3�\ɤ�Q���*�bVT�l����@ySw\EWZE=��-��
7T� ��6������
�>�^e�]U ����UD�fV�0-7�����ƙ�T�ɴ;�w�ѧ��ƕ�|���s���,��q�i��a��/�w��n�~���hw�/�%��.���i'P�PZ��KI�9�hB�I~uT��*�)�{&�L/
�Ӂ�s�^�'R[!ڢ���ޮ�L2�y�]���z�3�� RN�_�O���Q[S^�"�
�#rD�GP'q���v�a1�[F��qX��v�n�& ��/��u���1m�ү����9~��ף�
vϙ��i5��Ʈ��s�C���_0�l�yQL��٠�y�o>�һ�Ϙ[!��ZgQ�[�*f�V�\k����'�k�^�`��_�6��l--M&�;��N>~��������:�e���?M��U��V��q�5�Ӊ,N����ޕ�t�s�#��p�CY[�}Z��즩Vx�����M6���쬅&;�����ny-��g�í��1��m�Y;u:�*q��3�R����;{;~%l�'���n>�$z���3"���Щ~j�����44)�X,�����ՠ��}��e%3���No���;�9���a��Pg9�u�y�.��N3YS�}�4�R_*�iV�B���帚��iX�B�sm%�1��5�z�~el9\��n�����w�q���Tޫ�{��d��:'ܢ[�Le�a����;m����EEj���k��9Y���6Ȧ��C�Q�;���v�2��o��ˋ6�`r��޳_z�ChfT>Gmy���y�v�\��z�Y���y�O&�YR��gw�f���-�j䴻�C��w��e�6��VC���p�z�/{��v����V ��6�X4���ͽzln=ػs���=,�L�k<;"�5E@��'�,�s乭�?���6��ϳm^�>N3������z�h�u��v��C��{�z��/�vj��q��&&�z�3W�ލ;a��P�?}@}]z��K��D���U��N�w+��Ė��V�&��}__ק�ZCN!ϪRq�c5���:�N�)-<����z�j�4»^�L̳��>���wg_���~#EAH}��:F�O��,n��il�B��^��|�q'=�C���ĕK۞>�>tq����ꯨ�4�~���Kد��]n�c�ݶ�0I���a�\R]�*�3Ί�B��4CYWn�SPQ��B�
ʻ�>�܈wʢy�A�ے�v&�Rb��"�r	es�æ_;��7+6jCH����5X�޾���
1����PB��V��>09�bRVڲ�e�o56�b���4�n���:���Sy�K�sf{L$�o���C	N�7��ٿ
�0�d����z���tBo�����H�^�8R�A�y9����?jʲ��x��W�V�9
��4s�Y)-�swQ�ʃ�o����$�䞪	�R�����mBO-ɥv�u+&����&F	���^g6���t��2띝o��H�i4E�Ϛ!�J;���7�Nl�2Н͡��M9v@���d;We��o&�c\��݄^�q��1��#M>'�U��x���6�I6:��-/!���;��#�͏oΤ!��LOb�#` �^C����N����u6-��=�fJy[Bm�kb�@�u�qk�F]���1�����b��t�����f*�ɺ<fa�v:vN͠���ޜ�wm��-DU˗���W�;`p�5�Me9�
̝u��s6�=쩟%�����ewr1�{�%Btt�x�9����7�¨\���M}(�qI�e�VZ��vbŔ��r��XrL�>�����H��u����V�r�S���@��q
��(t]a��N̫�_N{�
jU�/���F)	��[�_ԯ�y6�u�ׁi����i���7@���~t{�M��Ӫ4ɽ���R
AH6'<���+3
�o.�h��P�J@�RC�D���n� �!uD��Z`eԉF�o^���Ă��k0�B��R'�S��-����w�8��R
AH"Af2RAH)�>@���RL

AH)!uD��R
AHo߹�D����ZCܻ���=�AH) � �^�RAHeQ ����(C�) ������s{ ����lH#0���R
CuD2���R
A
AH(��Wz����h��B��) ��W���R{(- ��*�) ��$��R
B��)=���!Ĕ�R
AHo�Wj֑�2��k//{䤂���i�L�e����~*�
C�D��R
A)8�I!uAĔ�R0����hJH(y%$�j�,�T��R
A
AH)��yD��R
M�BA`^��۟���q ��s>���?%$��R�R
%$��P1) � S�	 �
JI��$���R
C߯7F�)"�����*�)��I �w3) �5TAH)�RA�Jm�H)!�k}�삓�8��
A;u%���j��R
AH)H)6�I!uA�%0<�AH)���/[.�Y�?�s�֑:��#q��h���{�eؓ��T;z�RGl���w,ѡ:���]�^ ���Y8��R�$�$��R
B�)8��-!UD ����$=�����) ��
H"Ag�Ԗ�R
CUG) ����@� ��������)���i����׬�h���RIIUI�v肐] u���D�P�X_j�R� ���R�;�&08�AH)w��o`bRAH)��{_}�F�q � �4�AC䜺 ���R�Xc
H(��ʢ
AH)!�{�4%$��R� �L
H(u%	 ���ʢ
AMv� ��%���Rm��+fe7m��a��R
AH)H) ��UR
AH)d��H)�@i)!����B���?&�)-
H)!ڢ*��.�W�v[�4��I�)�d� ���^��d�U'YI ��$UL�2�
C���\�JH) �^]�H) �=�&��(Ja��XhH) �����J`|�AH)h��R
n�y�$>��m$=P- �!��
AH)
����i!�Q � ������]삐P���
A
AH)Y[�~�n�J�R
AH)H,8)䤆��) ���֩_�Y��̖e5��l��P�JM򀴇j�)����AH"q�
AH)��[�i ���(��R��!��{��[�&!I � ��v�Ă�R� ���]����3�� ���P))!ڢ��f�
AHg���䔐X�Ad�;tAH)&!IH)���sY|�k_vH)UR
i�
A���R
C�9���AH) � ����RB�j�|�R<�IH)U@�%$2��~@���R����RN��H)���D��R
IBC�D>���RAi���
ANn����D��j� �|ɬ_�щ��r�j������) ��$����g�)!��u�+(� ���}�����׳�i ���/�
H,/*���!{�
AHeQ�R
AI�) ��
H,?0�����ˢ
Ad�) �$���R
B�߻{� ��2~e	 ���ʢ
Aa�T- �T

AH(JH{wa��ZAM RAH^�gSD��R���~� R� ��[i �!�� �����
AH(UW��~�w�t�:\��W�%�ڨ��l�R���*$߮h$	Y�����:X9�חN�l�����9����7z���o���}��
Ai�I �5ｼ��%$��!䔐Y<�H,�%$��eYD��Y���I ����UO̔�R
AHk��;������fVg) �O��� ��H) �q) ���IL���@� �6��
Aa��-!��~����R
AH,�KH):�$�Q � R�z��X|
CUD7TIOP(������8ɟ�x$<�!!l�? iޭ�m�C��$�$�^�z ����BZ@�H,���v�!������|�C~�B� Đ�����jtn�Q���ڦ�nn�vn�s;1����
�h��(��1����h�[	m��V�p���6��J4�����
AH,R
CuD��L) �8�'�]ņ0��
H)��) �����w�4AH)-�%�9U�Se�i��Ĕ�R
AH.�� ��
H,�%$:���ZAH)����d���RAd�楤����AC�9tAH,6
AH) �y)!�A��
Aa���k{��)'�);���gwn��P;tAH) ����) �.���R
~��
AH) �/;��삓PZ�RAH) �9ui:�!�ݒ��)�����R
AH)��]����
AHww�X�v��e�e�f ���R� ��I ���R
B�X���R
AH,�e0��$9�߿W8AH) �i����w��d��R
C�D%$q��@�i ����Q��R
AHs��/{�I �K��� �����P�JH)�P�
g�J`[��?2�
AH) �?4�R
Cf��d��S5ܲ
AH) �5TAH) �`RAH)�I<����) ��
H)o��h��}�������ʢ
At������t�|a���AH) �=TAH(�) ���R
C�{��RYF�ʫo//� ���R
Ag�R[H)
� �aI �eTR
AH)� �����\1!}潽�Rm
H)�
d�v��2R~@���S�$[%$������S'I �i)��.�)�2}�s�́����R
AH)��
C*�)���|�����m��X�AH) ��'�A�����
AH}�٧@ZRN�HU�-4��}TAH) ���D��RTAH)�
@�(���$���R
B��~�삓�on�?%$=��<�H) ���D��R&�I�XRm�))!��hm ����R��d��32��̼� ��
Hr���X�ZAH) �u����I��^���_�7�l�~�H) ���
Aa��$>�o�R
AH,�2�:�N��R� �|��IF�R
B�)�IL4�R
C~�ۭ ��Xi��I�R
AH(hII ����R� ���- �i) �I) �������od��R� �����
B�) �4Ɍ���P+G����=�V�4��Q ��}�II39a�bJH)UY�JH)��i�D�) ���KV*��) ��
H) ���^5������\�-��ݤ��k�H)
� �����
CUD��R� ���P1)!�D���*[�>�c-�Ͽ}ޛ ��PZAH)UY��ɉ&Ф��R
AH-�.�) ���X��U�~�Y��w������{w�
O�Ai-�
AH/��P��� ���� ���R
CUAI)�2S) �7��ֈ)�)6�L���R
AH(u%$;�d��RTAH)��@��- ���R>d�{��6AI�����R
AH) ���dr�) �L��R
AH)!uD��R
C��<����4�����՜��y�7Jϰ������xȳgp�l�u�
��@z��x-Ʋ�潐��r�mO�X�vX���uK���e�nv�c��q��5	���f7cj�S@��X�np�����n��X;��s�ƌ��:�׳�N!�����3�j0�s⪍�@�V���;=���ۂ�\4��le!��W.����vq[�k���[&8յ�[`�nr������(um��n���U��������ו�-���r=uv�?�;_o<���m��뮹�. �k6燕5�ֈ���P���u\c&{`9ݰ��W1��M�fe�) ��)!�>d���R�R
AH/��I�]� � RAH"A`q�O�L�S�?k>w�1) ��ɶP�X�/�i�-%$7Tb��) ��� ��O2�u�$2��I��,ߪ�8�H,���}͚ ��B�>A�J���'+�D�����6���~�ͺ�(w�<�\��Ls�ۥ�����Կ����Y�W>'�^�bJ��|�QYUe���G0���ą6�|���!�l�v������6�*B�{Zӯ�3���z���zɏ>�����s���2wol��=�<�$W��_y_U쬪1);�9�_R\l��̪��q4؇��o{@|���5)��r�N��h�If�9�����������RN�Z�N��|�~�|��}�>a���L~�����UM��q�oTm��r�߅�v�{��l�5��w8���E���}���Tq{�!���d����U���=w�^��O_����}���N=��+\��[a�E1�Z�9�}g�Xӻ�*�|m��U��b�\~�øտ���k�vU�7F� J4��j.3(X[���k��)�������/B�X��Nd�ꓕ�oP�g�HS<��k;�z�R�I��.�̦}��<���Ϲqa��}��:���z��[���+j���*EFϙl���F����bMn�n�m�4cq�,���k���f��{&�۬�̭��r���I��׼&��߽��u=��=_}�P�(+��I�.�v�]{TOWݬ��}���x����!�+��WD,g�0^}Z`�y��vk*��)(|����T���u����潝��V�T����8F�V�w'��ȃӷ{��Gd2����j�c�Y��9�bG_^�}��qP��\�szܚp���J�O�*�=ܾ�COO�q=4�N��*i��h)4������g/E#��#��;�]&����.�m�f�o����r�����It��*��h��B�W'P����N$�mS�;���u;�ґN]��o=�^���������z}�oW�}��g~�5v��>M��n�2{{�E꺓I��o(_2�_n�iokCWEb�Y�/նi��_V��~���Ň�S�ﻞtm�����<��4�j����l�.�j���Ϩ��s|tbA|���O���W�W0�����.����)�(�>>�c9�&5��F��6�Tյ	�G�}���ܢmB���2x��w)��;U����*�AR�n��c^�>�>���Dh��|}㸳7��񐺮�}P<k٫����z�4U,�\�՟z�¼�øk}O�U��M�V���c�h�D<��6�������I�;]j��Żty���I�D]�d���u1�<�'L���v�']�T�0d�˩�V�QN��0�fTʩ6��w�����\�y�G7�)��4��V��-�/uI����ƻ�c_%�.�r�J��y$����q4���g/�w�p��)&�R�wU��Ƶ�ͳ+�]��ꔮ�b�O����0Y���w�7<��{����y'̯��f���v�� p�!�/��>E[)4�n�Wu�g�d��G̏�o��Z;gU��(�M��}�y
u��d��_��u�RY@]�5�+[�/	�FV��+F����i�wn�s�V�9����{����}{�r�OvR��3+�st~ʐ�7��nq�Hc�OSh��{{����=a�)�=�ʦ˥��%�4jV
�
�>�g��fp�+:�y�^}��/t������,��P�5̙�gMq�t��aL/+W~��y���'_&��;�gy�s�����ޥ��ޮCuP_?P��U-�YUuny���1�%r��ԩ�Nk~��ޯɤ;|x
���|&g�2O��N|���UWd��>�u���+���D��(1�g)W�p�M��ز�F0��|����o�a��(�YI� ��4�׭ו;5�Bq��I����ݚ@k�G��8�=En���±�y��7���L<�뮲���j���Hꏓ>�a��3�>g����cƝ�&�I�Y[�*�}�X{����&�=�����o�<I��>m�9�h�5��2GZ�>\kX�}q�IkĊȁ��������B��l����}���v���=T���Y�����S���<�|�)4�֫n�b{��il�s0���� V�g�g�>���
��zTnV���(ج�B��˻��^��
�E�L�v4����j9��)��k�b]=Gڥ��f����{9�H���R!���2�ܪ�(q�Ə//��C�6�ᩎ!�U3��r�sF�y��Pn�}1��nxT,�2C�H,�q�CZ=j��6�ڶڭ�����4,6��v��ZMj��\׳=SO�v�9��I�}��իf1B�������e� �E�]�Ï�8/4�qq�ut�M�fx��;m�D��7W��+�u7~޿�#�5�<a��/�ХoqyhI"Zr��<��]T�|+�|��|�>v�ʛ@���[MYk]r��o/3ahq�ю �l��ɾ��o۸X�KyMJ�@�����zJX}O��O�V���o��WP�Oɉ�߲�0�'Xik_z�m�l�[j'�|�̵���-gy:���%��S�+�<�v�б��On��@�n[2tr��#�n���pQ��(E��ފ$�_.���j���T��,<�(�k�ߴJ�O2y�o�ϲ�?9j�yy΍?j�O��YSl�aM��)Y^�I�5tc�5%;��W�8��SPNX���K��MwS�8y�8�7���J��{��i��a�,��߻{��S�ķHR�{��T�i�"��[7��<�{}�h{P����x��}�ͩI�>U,���v���X�U`F ���Q�����X����z޽z<ͳ��8��c6�ׯ��BT��]}������ԳuIVS��fO_'v���^v��y>�}���ٓ�Ӵ�/�Q�Z�����媿Ykn]�̼��ѾV���l��=�/���Z��C�����y'R�`n���Nk=�h1�蘞s��i�S�����mk���Q=��P^�.l�?}�nԬ񯚩^˻�����0��;�]�T�i������~���4������*׷>U�������E�f�y���i}A�J`i���٣�ʩ-�KG�c�o6��]Ͱ��ǵ&:�>��N7���s���7L�]�^������s���S5	�4Wu�tj��h��;�w@ٜ7]�J��S�6��5�l4�u�v�HX���O�k������'v�Ӵ��7\��yc53nd۔��τ�7εrm),j3c&�xܪ�W�����N1�^���i���Jo;�l�47���xP'�=X�+�d;?��}����;�j�S��R{c�nq�nju;�Ų�������n��>�mph�\Y�=����uJ�`q�<��qӬ��V�e$6x��dL�8����ȷ������ۗ��e|�#۩�3N�q�3���x�(�����w��{Hg��ɧ_5��6�������5a����-���wvLg/U�l����|d?Pr'����L�_����V#1�9�^�/�����y'{���<��S7^��E�Ueݖ5W�,GI1>i���T�C��7���R
���K�{M�ǹzw+�m4'���/��C���Ϲ��S�}ۿ2���|���i?:a�߲w*m=�l��+�\L�7������b���7��%,�Y����*���G�擝��u��*��}^��9�Xc{/i��{5��O�D�꓾��ۮ�U�7�&?=m�;�f0�'�e��^�i�=��l�0���fRn��EDHQ��/��ƺ���@W���s���r�V��2��q��_p<��n3[՚�?8����2��Y�N%�n�LϾߝ].<\���-o�����wZ���/�f�YID���ı���t��
�)\���B��Ki!Hm=߽��:��߫���C=�^��}PUr<���4h��-�Y��j����f�N0�2��kFe�m���:�9to�S���w��C�&�Md�R�((ϡh+'��vx�mƻWnU�zD��u�p���v��x8c�n�;If�i�����,�)�s�߻�V���Զ�����v��t�u۶L����O����4�i]����&�i�I�r��~O^�|ͥ����K;�ݗe�^)��f^�i)��F�?��+��ģ�;L�FVs��Y�襏ʘV�jJ8+T2I�+q|�o�nؗ�۹�E�k��]�$���*�xE�Sz�9X�d�ݴ~�uO�tŅ�w��������U�[|�7��
F���
�M�E��Lyړ��Z�sw_km�n�ϹF���)\k..J[ʼ�q8͉3*�N0�|�{[�:�ޣo;Jm�v�ӏX}�o�}�C�h��I1�n��>b�C��
Ow�\`|�>t��T�g7Z�D�,�l-1LN��l��NP��+1��S��:��_{�f���}��硧Ⱥk��oD�{(��QHz�`y�34��]y�m��=���u2˳��7���[��c�w����I{up�m��C�K�Y��H��)�Q��L�-�m��&�����__��D�8�x���ۚ���*�m�o1��!��>A���S���)�۰�g�c6�Nj�����^P6	\���p/�V�1)�o<�۳������;A��6����׉�����%J-�-&�K�G��\{bZSZ���fٛ�|������>f�����"��_$Ӧbf>�B��JN��H|Ї�(9�o��eE:�:i&��4?����I+t�����o�i�b�b����.o��������m��;���Q�Vٴ�)��_{�h��SiM��O{�ө�ֽ[a��wA��i-�ww��U�Y�ɤ�}�g~Q�g_�'��������{gSq��X6��u�)�)��q4��G�y��|���m
�Ş�����Ԃ�O��q;�[�.,���71�ڒ������f�+����Gy�(�*���qDtr�����{����䀵��I+%�m�� *��f�޻�������˨ZO}�l���>Lt3ϽP�Q�^��ևV|^�:L����AD}T '�3{e}���׹��5��c!uP��~g���UN�I�<{{٠�f��IķY��TX^��t���|�׹��gp�LT�11����y����Z�-�Ė��Zƍ�S1r�w��Sڣ�\N�|�W���?�N|��н�;�0|�ڷHW��X{�b�׬�푪--�~d�k=Z8ϓ��Gr��E/:s���OePH*�D���6�|��z� ���܊���g�ܸ]��8��gۮvݭ [�(�y����*�&�ǏY�����S:�ri%$���{s	�v�g���d=���A���=�8���ѧM�!I�}{a[�ru�8��j���=�J��lk)�V�2�E�����Y��}킾7[��}	ڕ���ӓE�������ג��-2�|�2�u�_�ݠ��}̶JB��u%}��֝�e��=�ju�L�����Q�_AF��P�f�KT�ꮖQNf\�y9��4�>z�������Ka�u�I�Q�c�߮pUPm�]J�)
�?Q�4�n�8ܹHZO�w���Ϲ�g�;�%7����}�c���@��Pvd�=D�n���������z��h��? r䕘h���㳷���Y�YYE���7�o!��ͥw.�4��&(�[�Z��N2�B�J�5�W�f��3��P:+�&S��mO^�w7��Ռ1�q�K��]�h*d��J�Z�o�K�\��Z3�U._�o�WX�w�4�]�r��T�k�-���̡f�9Ti���=�U{��n�5��4�ʯ��r�{�u+��)>�k�}��;���&'�4����h��)-���_$��p�����Eh�>�����_U2jӺ׎���&&�EKu܁�4y�6t�9{\���U싣��8<8�z�*�@.|�k��֐�Hz�}�e�Jg�E�5��Cl�=Y�V�ɦ|�v�gGՠ�«�����<lqV��D��gwA�Z��ޡ�UN���y��n�:����1��!}��2�V*g�+�����UU�GW^h�����I��f'7��;���N�!��%j�<�u��@�� ���.iX?W�>We��������M�@�l��h�>?��'�8����V"H�l��|i.v-꽔�N!�mo�:�3�|�I�kU1T:���s��o�Lc���L�ƫ9AĴ����v�<B��}{f���]��~�>�/�}ˁyP:�|�^��E
����L��8�)�+]�dƽ��U�Z�
_o>��֯����í���J߹�����!m��=�߫F�VZ��B���ר�~�1�����/�}��c
�VS�֙>�3�������ٴ8�>v͠��t������"󵧈�[�D���4W��;�~�k^t��Q����[���u�4����A���L�N5�ׯ]]�p��}�<���L}K�|��Ó�.�z/Ҭ�0���9�ۛ)>�kF�Ki\�����^uY�K�z
��V֕��gqv��d��EZ�HIQ�1�{P�ػT�u�o�DϽx79H^��~у�$�=M��˺q'2�gn�H3�"�2�<̬��n�>��,��-vE̝�h���HH7���u*R�[9��ﯲ�S;-�`\BL�x.P]���nbcwt� �Am�x<�ު*����-)(yV����ޱ�7`�lVx��]e4a��[rb�E�nʝ�2����r��x��!�]cg_S�ܶ�{�wm!Ѣ���;Cm����U�٫�i����Km춅 '���"Ӿ{V��;:D�|�]L�͚r�.��;��۶n�>��IP�)Nٶ�\-1t��L�����v�<�uԼo\W�Ipc���J����#[lky��ց %mՉ���L`T��%|�u<���Y˫7SY��M���]r���fm4�jt{���Q�R�E�*�]`��Ef�D�WQ#���uxwX������9�E�����M�'�.��:��V�N���F��-����B���@����))��m����|x���/CLj�-��#�*3�Q��	{�vAUNkz�e����1�<��\���dt��i;�w�9�k���,C♷�����[��)�Ypq��ô`ٷFP1K��;����g]�QVf��vgr��v�¤�O�J�}�+mA��Į;y����Vt��!VE$���hd,ul���)mv;m���0*�Uw�ۧ�+��x}�v6z�Fs��z�5ۥ���7�q�O�Ys��'��	�1:��<5q�Wl=�]Yn^Y^Lzc��|{�}j�[�yh`�h��q,g+I����Qε��a�u�7W[p�nf᧊}P]XQ���	�a�}���#E�\fW��8��2�0s���W<�4z֓�l�5��-��cf6��q�prm��S�m������Ϋŗ��nU��烷��ul��ո�Z���w����j�˳�C����i���s\�F���n�݌R����5�l���MK�˱�m�e[v}6q��^X���;�+tvڻ
;Qշjz���mk'n�wk��F4�^GX�7g.i�;��ͭ�n�t��'�aC���*ۡSF�x��D۔�4�Tr�l��d��yR2�����nŵ7k���u���U��KnM���y�v��
%Q�	WB�Z4]֪�����[W[�nݻ��ʻ����p���#ֳ�l�v�e�
�Cq�n^�fM��i`t{7B�6��tz\^�����<���86�.묜�Ӄ��ۦv�m�<(�8Q�p�7%v�7v96ޖK�xy|H���G<��8�������x�7={m[c���F�^�n�������ܖ�:��`��\��N��; i�v�\�=����q�����\c������
�7]�MgA�=5�΀��w�'��c�Q�H���8�c�=h�N�7r��m�V9�{;�S��)����}q] lp�7'湸sd��z�o�ƚ9��'kW��I�J3��h繱�:Ɲ>�lq<�g���p��ڵ��&�v.��yd�ۑ�n�H����wf$�g���!��d1n��N�N/BgW^��jw8شCA̻�0Η&/o<�[��p�p���;����n(,˄�r�wU��y��d���m�o$:n6��M�#�':=��n5���5�;r�c8��D��g��Gu�Xkd�Й,�/�[�������3˄룑�Ts�7X�[���hb�;�n��jl:d�n,n�2��^*)�N��|`�7��%ڛ�c�Nێ��Bn5OJ텟1n�a;ϬkU��9׈�`��Wr��������.͞�y��6����v	��5���k�U
�6�uƦ8�m�e�������ў��g3۴�^��2:r[��7;F:�μ�磮u��D �-g��j�W;�}�]��n��ꋘ5W�?3�}�X�����XkT��6�'��
��ܮ���w��W���u⥦���.��>�C�����V����'���;w��)��6�Kw�|�.O��5�ȱ�u�9�',�В:P�Z'�<.�y�������[imI��Ѭ�b�{ے�̺�ly-5L�>U��fj�8�{���[6�۲m-S]���KE>���IN�S-yA��[>��E��kyo�ϯf�ϒlm�O���;�m��]R����Z���[�l;�����kS�m���:ݓ�C���g��q6���^��_.��ۣ����hc�s��n�lC�4�+��J���{t4통E��i3޳i5�=�����
��
0��}����?��=�}�^�Z>�3�2��}�6���ou��)�m���>����>w�Շ��Rm�����*5��B�l�����t�9L1{\�ٞ�o���M]�Iܨ�.��p�W�VV�+(���u����kU�y�_���ѦL����R|Ŕ�ts��+��z�������%������t.�<{��[�+iw���.9�Y���9Ƿ�`Yv�N��+�Q�p'[�=ЊM��'�6��r%w$���%����z�iТ�fu��F����i]�̳�,��'�Y�����^�i� nM��l�niz��y����~>[9iŢw��8����V��8�h,�33|ޢ��xJO�ח�=�u�Z��&x��2���uM�cT"��S;�屌��u��9~V\��d̤ �P�� -y�x%�!kfˬ��	�1f%������S���oexg�Vn^�m��$����E����-�+V�ᾢ0�IB>!��ctj��4zҬ^�	m��9�O��q���������{[|3�� ���b�'-��@�Ib���!aȠ�tM����~�Ղ�eM±]�o��&��w��st�Җ�ᏉQ�ӎP��	(.��N����7�r��'A�%B����?DN1h;�mD��c��J�p=��z=c��Y����T���/f?R��WwN>�]�4��c�F����P_�j�|P9/7��Id+�ac9oY;k�r��8�k�L��o�"�[[Z�L���񥽸ż�P�SO��]?yq���[���û|h;=���E�R��h�Dī;�]���%��ZG�x�>����cA=�G_����r�q9�jy9��^<�܈q��y���*I���=�z�� V�&� �I�������w��wr0���`���ϭ�6��z�z�)9Ժ�u\I:����&V�p����e���Ƨ�j;6�h��ӣ_��k����{����~��tV1��{a�����v�G�;�6� !D���F��� �m�U�ve{!תQ�˩|Ƽ/v�{kK�ǣ̼��r�٧Nm}��Yϯ�-j�b�v�g�:���Ѧ-+ =��W ��棊�6
De�Z��)�6��>X1>*>#����*�lU94�\�^>e�Z��El��X�v�v��ҷF�jwO�-��Ǟc�����t]���ʶy�'�|�0�Z߿���ňYw7��~����4yښz]��{�5��������t��`s *�;�	���6��,� k=�� ����I� �wW��V�}���GNd"����X| ˮ�}����z[ݏ�P�L]`=�N��}��:wǛV){e����\���k�b!@Ve(��|�����_nR����,Vs.��b�۳�n'��)��;��WA���~)Y�L �c7����.�%���3��u
\�] �ѳ�8u�Cs�7���SW �Rm�+��7�&]������rh͞(��=j�ܽ9r
�s��=XV+�z.�;Br������44Ƥz%Z�����W����H�eX�jc�{3�gM�r۰ʫ `)��F�#�}�[��wYĉY��]�5}�
�9�5e�\\WZ�u$Xkp_����{�&��%�eِ]�������W#i��GTv�PI*��8X�g^�
]����<%�=���ǝ?�sv_�O1i6}ˣ���^��{��Y�ЫT�O����\�|B�v�;\t=�P0�3>��^ݝי�F���P��(�@6�A&�Z�pϭ�SP׫��tM�b���4�jj��b���LU���o{+a�����1���+5�
���ǎ�)9�(�$���Rgg�q��y�;�z�ܹ�&�췝���9�N)�&��r�M�j��\�r�����/��4��-����	lN�۲��nuB��u��5�|;^?"<�n��gB31��vޅ��{wa������Ņ:H�<��rv�;ϽRUy�h�S��'%�}�2�\���4���kH��G՚����^�!���ifi׹��K�T�~RL�ۨ�=u�~�����dSa�y�Z�8��cx�)f�W2�$z�v:XbCl���n'8r����Ĭ��i�v�о'��_�����t��j��l�H8��m��ses�k�l�y�l�գ�U��A![�9�#��hr�nQ�S��.�nm��ץ�}m�ۻ7q��l��mf;N��6�y�c.&Nu�=��E������ٸ��-�lp����u��a;����i�ns�x��u��C�)�;oe�;9\��@t64���j�ݎP�\�]d��9i:ڸJ�7]�&s�۳�Û��A����R��!`ɶ���oW6ݎ8�rn���غ��5����;�<����y���q�T��$K\K�)�ڦLٔK�Q�����|	�o@��2�O��׼�_�m!��~�}a�t�M"�	׼vϢ������J·܍�=��^�z�S���Y��Æy�]��\
�C2��F�}�V�����uc��i�.��݀9cp��<����S����G0��lJU�&�K�Jz������/��HYu3���W�gF������^1:4�N���鞛�o۳�}Ő3��W�^Ԝ�(59K��2�:�΅^��9b�JOb���4�&Oݹ�� ^\ᵾ�;Q�KJ�D@J=o��o���[FoW.ʭ�T<ayq���{=ʽs=�¼��gv5 ���_D��=닮�Q�2K7O���z�]*h�8B�� �Gv|�(�5��28uf��9�]I��Bx=�{<c<)��%��"lwQ�Ѣ�^G�ۢg�օ����9�$h�|�}�_�z���L��4�I�ԯ��d:�u��k���h�h �bU�OP����e�2��ذ`&ǎ̻�k1	���PYʍe��vV��˱>q�=C�\�]3^䵗`WfV�_��ݨK�1u<��T差���W�ֆ�Z��MU��+|nl��J���,�79��D�1�v�yS�Y�}�[$`��#��ً<�y���(�J�I���6��g	ۯ}��:�Ri�T�.��ϗ�ف��|�@`NEh�P��A7��ޫ��E?6 �nW�x_��v�
J��7:�� v���o;��c{���Y3 ������n+|�+5K�;�;���t=h���v�Ζ�,ի������M�X(��=���`�q:��p��^tb��uP��+������������c�W����'��b�����"��<)�۽Cpᜇ]����znO�I$�#��N;<v����\�gρg�AF,E�l�흮7qBz�W��$�i:���5����u���щE����FK��k�Þm�W��1��U/v]��H:D�*�����r�#�y�ܨW�� d����f	*'�������R������D&zs�z�Ԧ��=��CF^���
[g�07B@&�1����l�zm��E��˖�Y('�+��憳w5n����ܲQ�.��w�����g[ul�yO{�WӪ I{���C)q�;�VP�lm�}�5J��V��
���زN�=Ok���u`}�q|���ۏF���vwY��ڢ�u�3f�H�(+�](�f��(4M[f������qgXV%�F,o&��}/�������N��u����,:�8�x?1IJ`'�b{=�Y�(a?/e0:�.D�����X�ei���|�+��F�E���9lظ��S{�o�����$�7���5��o����GK^BZ"�-ŝa�	n7��Շ��F���
�\�㥫����-p�q�a>��K�>�IK�o���Ѻ�OV���Һ.�����"I�3o´��c�/��ih������=��׈�^���q{�ը}[E�[�Z.q�2\�\���}��M�=gt�|������պ��+�j]�^g���Wg5��5�#3��z}NV��/O��)�9�k�[�ܕТ)C5�(fDo����[��}������E�z���T�en����v��������j����C�����d:l�`Uҧu�3���(w��,.{�_����YX��/onv,�ߜ�P0\~���lW���Z�;�x�"�n�	e�9���v�-㚩nN�]�I�y�=��p��5����J�Q���M�=�3�'����[���f����"��?�S�c�M��i��B_�;�˳��I|�ְO2�[	��/Gu{�R2R���*�(���m�8���Ѣ��7�e^먅Q�N�i���V�X�s�rف�N�e�l�ck��
��n�v9���]Ԑ��L��C~�K9�w�2�+����v��������՚����ܞ�'0=�5�۪p�ɫ�����б]GKK���\��j�T��\�^�!��U����؞�@�x��-�g��%�[OT��j����JŞ~��],+M͵���}y\��v�\Z<�݈a�@�Ch��:6n���m��2����Y���#О���/g]�&Y��uw_{,������yYX*��wE�V�r�;�~�3$U��A��4�U�wFϤUx��ΝJ��Z�}�Ӈ��aܰ�����5���%bSݚ�6��y�P�==�ǂ[�{+X�����~���@�Ab�N�2�^���е�~}1���+&�h���T��������.�ܐ��5P�v���4�J����d'�f�6�b��P@��f��5�u��Fw|�ݬ<4�ʚZ�y��Ʀ��X�}+��c�5�s9��2�"�+.�q����D������p�ju���ȣ�=�ZF<��Mc�nKu���57[��wOpn,܇�����
۶9�w<�������ۨWzۦ�n��۳�;�;v�mn�Έ8�m��ѭv��I�s�<R�4l��'q���s{73ۯ9�������Ÿ����4"���s�.����;J]U�V�s����Ş]f�b�)9pZN��[Fn�\k��k�M;��=��x�)������Ym���/ul��n2��u9Z/ߚ�u���͏m�y�'�j�p�r6���������f�����M��|�u=\#�j�wo,��k>��6(��?LdPt��%�e:wV&w<��^]M�_k����ʜ��yY=೽��rK�o��~M�wMvT�𭘾ai"���+7<8]���m���Q�xկߥ" kO΍y��?1���ߤ�r�<����[��uE*}H��l��{�f��8wV�M5J���*�w�{�ĕ/\�������0��\{f�:�sKmY��X�uO�{��W�e%�v�;����(7��$Ҕ�Y5���������kκp�hh$B(�3�!z{�����3.M�wNx'6��Cz���q{؇�,��{B^�+�Ph�t>���w�x�B��uc}��9>��^��ڒş0+n��ߢ�l�;FlR�� D{RNs	�>ƼnV�1V����12k��:KS
�u�>Vk�ʳ{ުg8]�J�m�ެ��`�X,�v�yvH�m�γ�*�v�&M�w/{�r��i�����h�b���)5uq����n���jzք�����>+�Gu�&g���x1�V+q�յ�;��!�]�W�/�y
͛�*�*��7��n�f�}�>yG�����q�N�[={�/�?+�����6�U姽���F+�s�Fɵt�׷ަJ�[��K�w����w�[ͧ��S	~�D�V!{ӻ��%n{I<wբ��<��Q���1�ݝu�מo�BK�<�Dy� ��v�F���*����>ܖh�j��җ�oЬ����b(^����7.��L�ŝ�r�� �r��A�=8��/���ۑ�
�mm�[W\���j�,�f����_��&��|&]����+�SZ�Έ�����*,���o�/j�F�]�8�96�k7���܅�Z��R���(Z�V���~7f�cn�9�7r��H�PM&�u��O�̊Z�� �+f����Z�j����4��:w���ux,�3�trx�����W����'���)ٵjz�{^������ ���	%D��	�[��`aג�ȹe]<�v}�{{Ү!��������+6����}��x2͵]F������ɓ�:9֙�ɰU�%z7Rh:O��	/�F�N�{	ƨkUb0=��������9/I����UQ�Gn�Lf�v��5.%y^x:�Z��k��h�1Yv��V�x˃�e�j݋Kw�$�e��.͔������;W��*�րE^��0�4hʀӄ,'E�,�BގgBgU���K���u+ G�ɣ�:隳�qK�
;ۄ���r_Z]4;�,�N�.��KW[�G6���������lI�@�gr1�(w>8dw
�Y����&{wz���z,t�ͮ�b�m>�,Igz�����S��$Y\g=�{y���{}�3��&�nN	��4�����u3U�#���c:��iU��ЗV�Y}Y�y7��sT ��\{�Ӽ�H��4r)uf�f�¬���\�b.��@��n�{n�di�s���W^J����:��>)�Z�fP��ak}��͊�uvxY�ܶo`���1<�!�y��¼@�?�{�Oo,Bև9G��8�6L鶀�ߓ��9}ذ�gs��cZ]�y7&��,J)����+����ܡnc�fљ]��fM-n^�J-㮾������8n�9��o�Ӡ�$��N�Y�/O�Zai�{HyZ2����V���i�Cyh㩁FqץJ��okH'���f�^�"�Χd	�5X��j�F�w�I{WwB��Uf�����4g;}�"{�+#7�I�˽����ha)$2j
X��Nz���
�@w0��bt�N�<"��*��x���z�y}�6�3b��Ҭ�ϱ�B����'���[]�g>'7͑�7��z^�߆�PM)�H����^��r�R���~���wXV�[�V�됊S}n���\��ߦ+�uMp(x5X={᪝f��	Y��0K�ux,�a�V�r���8F(ۼ�o�׶��D_�Y,ҹ�����ԟ�OJ�Z�/֣Y�ܿ�PѾ��WzQ
�]j�so6���Y����b�V�x��2�k��[u�ݺ�s��7�6�]��B�d�<��q)\��BB��ܷ��y��fz�|�\�vދ�t�1���^x��~�F^�;n�'"��Ҿ��@��zJ�R��ٕ*�[��r��S(Q����c��
wqг[��S�0g��͢�W;�=:�TȺ�U��T�{����)��R�;]m�W\�����)�=�z�=:r�Ny��P����n��*}����u�S���j�c�rwq�<�Jҭ�=6�+6�d�_��{�7˫ˋ���)g��h��s~.�M�c��V�mOϕ���O���E��
%�<����ʕ�����nZכgz�B�j���U�N;�ҺXǦ&��B"%��ͫ	=�!�q�ܝK��6^�g�[2�'����`T�｢��T�g3u��sr�ՄqN���<';8v�:�����=�f�Z���ꇭ��jG:8Ӓ����-e<1����(F���5o՜�wH�n���'��v��>��ԫ9��#�->YVU�u�����N���М�o�`�+��Z8��nS��x��Y��V�ٻs��vK;,'2Lz�q{�3nO+L��b�m>�]ԫG��Ա����|��p^�{���s��hҮ�{�Ȳ���N��v��1]�MOB�@^�j.��2��aE��^#2������p�t��<�p��}�ɜ�c�ߟ����4VN~sĻG�/,�H�<7��,�k u经�{���=����D6�A$��4ج^Zav�eL�:"gS3�O�y�M�D�o|/ݘh�:��ޛ�*�5l4�������m������3Oz���>�����]\�5�7��3~�Ex���1v��k>VU��`G���; ������i-����5�����P���s|�d��BUm>h �����\��wx�g=R�>)�)��3&�iXW����h��ؘb���_]N�)��-�䮩#�ș��1�v{SVgG�b��WEp��/l�vq�+e���6�
t�j^���{w���33mEҒgVW���X�=</oWؽx5��@�J�QY[N.öNg�����(��ֶ�1f�ў�P�q�kq[�]�7n�������鋴'lm�����l�NM��k�;�;yЛ�A�bպ��ilq�wTv�ۛ)�,$0v`�h���wW�Y�W��s���m�7��۞;\m�<ňR����7/mV���/�9��;s�v���L����wC�\�<��A�n�W�9`�i��F��=u�.���m�sϫ�=����hz��(��-u����^���?z{8�Ú��9IB�˯�_;�Nk�Y/�{�T��>y2�l�:&o�(��®�nn��#"�,S���B�CE�0o����1�~���cq��t�ß��E�z�����Z�,��n��O*f�qf[W��LW+���ph������8��Y�-mw�r+��LN�>�N6��XbV��y������'�?cw�y:��A*������"b�{�����?yWe�9�鮰e����r�"��ns��w�ɾ1g��hN>�=՞�:�g��_`�� �u��}�^��_1�������M�f��G����>�^��2�'��P�h�K ���}ph�Y���� �=�Vͥ��]N�h�Z���^fJ)��F���J=���{_X�\���W�<;2�>f�&�OnQ�H�����p�ƚ����\9�/7l�<۩�vl�����[��B�X|"Z\������h����g�׵�>�,�ew��MMj����9mr��J�P��S��m���A.��͗r!��9~�����!F��H=��� �,E��t���j����L���i�2ꑸ���ʕ�0��]^��z�n�ʿWe�k�e,�z�MTĕ����>��ƪ�8�XJǰ�R��{t����<�L���f�b@Nv�o����:��y
w�Q���Ty�)gI탅v`�~E}��EP�&�A��xDAh��[�4z�h����瞥Iv�9����fr�{7:�CT���=�m�Zj�׳��u�:�lU�l���팊����C7����b��0@���VŲ�>Cr�T�DP�t7s ���y������:����W�+1X!���6��%��������)��+�ut�*�L]F0�����7G�d3�b����3�N{���׬�Q<#�����+4�6��)�q�K���y
��_ 
�>��ua�㉳u��5î�����8���N�uΗ� N���H@^Zzv��=�'5�<S��B݌���c����N�h]Pu���o��41K-�.K�9{ޗ��߈��U|���X��Y���I�hФ�Ѡgs�s����Ƨ���}`�����u� D��w1^K��v��}��h��t��V~�0=��ݲ�U�]������w煮)z�b�>F���%$��kYϗ^�Ǽ�^'�H^�>�ѳ�u�ʰ�W&��2��3��iM��s7M�V7YZ�%����x�V������ܠ�b[^K�D�ǅ盍-.%��|���9h�y�n�{sWX�4�۬��;h�f��>�g�� ���=|�5<:��D��0E
��{�m~鏶_'^	?}/�.������*=wn^kzh���x�f2h<�$�w=�ѩ�
M�W�X������=��>�U^z����S8�A�9h7U�������]{���҉��t�V>�c(��K1n�����K�W	(�I�C��uxX�<P��[��2�*�����Ѓ�Oi�_���� ���$� �s�@�=.v�F�l�9�ӭyxx&�.�*=tO��>qGHF
_����E��*�[�E����[j�şTGW�_�?0o?]I���%T�P\�V���U��g	;֙�T��6�sX"��`B�Bn���T�_y�T����h��`���W�ia�����T���V ��T�u�ۣ~�D��(,}��T�}��o_)=�51�O�R����T5 ?m��O�kˣ�ʞ��6�w:_;�n��5�.��{G*���w�?c�)���U�+;/L�}��z�����k]���Fꭕ�[�h���\Ϳs�ή��o��M�����5ߟ���9yE.��W�{���oo=�k[�粃��e��iz���(��6����U爘R�V���ym=ɽ��.�`�MT&�g���M���k��]=MI��eL�|6�TR{&�����K����:�]�v��Ș	ϙA�o�.4�Y�OV���O��gM{+�
xo9��)U��x�)�����X*
^!Za��3�l�������:�V��P��۩�:�+��ut;���d��9�v;V&y�sS�����0�,��'
��������M���2o5��H��j'ނq�JFT��=2Z2��%�y`��t �x+#�IS��z��}�j�'h{(�N���v�5-.����լY��ֻre9=*M#��'��U��^�J��w���Ϊ̮�v]�񯂝�wY\Fh��?S^�:�����Nio�9wY*�2�J�`�Y]I'��{�^�֊����ݒW�0+5O}�٨�s��}��޺�>�eo�r�M�P�u�ϝOw;���<yg��>ʻU�
ѶXIm�]"�]-�T���@^�m�rzRV^��8����/|�V
��=u�f���y�~K�c/�n�im�)V*�.80'�k��z��㨒�XKo#��i{��*�[��_������{j9�ZE��sV{�����R�o=�8wv���E1Q�Y��z�^{N�eh�W4s��ݭu+Jm!�*eC3(<�Z2��U׊rrd�{�:�劵Vh�;����Q�~@fR����ڨY滭빭-Nf����m�� `�(��8s̡nb�[���6�-V�ܼuΓ�N4;jӎ�낶:z{qWXlvY�pS�
D��WF�l�W��2)3��t����<�XHM�=e��ɺ�v�W
�vx��A�u�9�4�i���X�m��ju�8U۳�/>�ܢ��F�v���v8�^�V���"�祦��[����ua�'����E�3fö�{6]���x˜��w\16��W��4'Qv�<���3�s�۵�ñ�\4�
%���\?P�.�	���
��z���7)(�����*��5�Mw/eG.�^��Ѽk���f����sK'�ĭ�|9*d�+�y��L�ɢ�i�V
 2�{fa� 2��%x{� +T[35!6eM�z��u�:��n���&�-�9�	����@ʱ���9����ڛ�����ۡvA�N��L"Sذ�,`�j�/|.�z��>\�l����b��n+ey�9�y�����?��mz����Y���?Z�R�	�gZ�Ӽc�z�6����#RJ,�Lo����h�Ԧ��}�P�k4�D%B����/��)��?T/��S�~20�ۙS�W��9��n�j{W�Խɯ&E#�0�.��j�*��mc�j���V�Te�s7�iq2�1}�	������[��p��2�grʲ+ �����a;9��Hx�Оq�uy^���ij�
U.����m�n�˶��dx��vy����t��f�h�v6dYJ����>�m�CO�Mg}ٽ���m��3w��?R�RrP��)�S�p,�;k����Y��{x�ǔ��Y��X�!h���A&%��U�72�A�����h��u�
ڴ��6�l�xj$��ƨ]�=dx:����U��lnu	�6=�.�w���y`�5����C��Bε�E�0�:3�G���hH/�R��Vn}ZD����`�W�d����Q�B���N�I�Qt�i��W��%KLz�L���y�����N�l��ˢ��W��T'���c�[Ss]�6�%�K��_Z��1�LOqG[��_�ߝc��[�� 5)��[�Ͻ�S����j�Ëp�K��_Z����|��J�o8{d��������ι�߈X2�����`ѽz���V�������~=u�g��)yyP��"9N�m��]/ɿ`�]�g��'�Y�9V,�����hN�7�L�w��'������k(��g4��לޝ��g�J�&���˚�=��Ξ��v�:⵶MtN-��<v�����js*�(���oZ���k�3���b�}(s�V[82����0S꾻���^87j,T�ѐ�b���3v���V&�����`�	&���ԫ<X�Cc} �������x�~��5��{�sʊZ��ׯ�֘[=*u�_1U��u9e�ɻ�7�D��w����)��M���7U�.m�فz*�><�7ϭ�K�}�»lU6�ܸHLc�P�(��yE�t�������$�k��W���Cr�؃����C��4oJq���;��w��,*���`����.�T�V��R��sp��ѿ��E��s��P�~���@e��iRe���
pOv䧢�<�^�X��k���>�EbʇL������x�������n�&{,^{9����n�C�1����a��]R��ZE$�kn�q�H3m���yüҥ]���l7"��j�`nxb�
Y����_�᠏��/�;6�p.��U�G��aҟ�Q�=��&i�5�P^��'Tnx��;r�ݒq6��m��d��;������J6��/<�v�1k:�T%N~r���F�V���ʀ!b�<5�rOM�_{��S��	|�AG_�g��9q�V
��:�=���+��5{�(�g]o{�]���)���J�zz����Q�������?,K|�o���Nw�gWJpՋe����A��9y=�{�EC龪��F�(�&��0�4M_�B�yGا(G��B�D|���b��Lg6���O}�i�On9c��!����Ů�G>�P2����[HP���(�������gf�w�+|P��3N��+��<ʍ�6���X����AZ��Wwz����t��5^�+�/X(����e(z��+OgEkn��1��$��k�
J��l6������ű���Ϝ/}s̬���=6L��Q��	ҡA���ʩj��\��c+5eԱڼ�B7د��G�һ��3�Ѳ�xֽ���Q07�(�l~��'Rݛ�y�)��;s�ʵ\�@�B,rA�@���yeB��[b�sc.���\�z;p7vw7l�9����eB�0LhD�z�E��h�\��Fk�*�x�g�q��s�|f�ۤ��:�9e��ܥk.�� 4�~j�r��2��8��w~��E&BT��	4��UxN���{�b}����<e硠�V�-䃧Z��e	��
d�:m+�ÿl��vFK%Q�>^ui}]F����疬�z�W��ʵ��J���m�������/���+ �'PB��̟4��ݶ���U��Mq��R�a���޺��AH,�I��W�0	B�,VA �yC��J�m:{2�����n�z��N	]�z�c��V{s_�ޠ~�LU+K/��WW��h갫xK�*��6PMˎ>�{j��R����?�T��Mg����������5��̃������koH��F�~ҕ��,]�ً�;�B!+���:>�paz�PG9[�b�(���>�l_��UW%�.����f��[���(u1a�O���c퓭36�s}�B����Y��]�Nݒ��C��<k�tܺ���W�9���^�C��T��qΡ|�mV�:Tn���b@R��{!
b��Zr ��έ�R+��ҧWe�c�җ�t$��O8�o$,G2U���4��+1ekRi�,3��p�����dx���S�DsWf=4ͯ����J�dS��A�}����D�ᐫ ��+�Ӥ��a��q��n�m�c�v�oR��\�)��*�J�EN�6�p�XN�q������	�¯F�[��lV�_}>'�J��:�j���7��@�3�3^�8�[�T�:*�{rr���-ȆY+
���+r��9A��P�s5q̵�K���F�j�ϼ3B��:��b�ƞk�Y�e�\3���ز��gV"��N��7f)Ρ吊����_}Grxl�jr��Xȋ�]����֎{݃���G��7
��𤢡��yG�c^�g��׋�2�kE0 ����J3<ʃn�\��{mԖ,B���TCo0e��*��&���6�u����:pV���<�V8���U��47�5eR
CB�9w�EH@�!�Zj詩�����X�mFk/������Ю�M9�6v�H��a؝wY�g3�9Y�f�E�2���8;=:.�@�R����{i�=�y�`E��s��5���yJ�%�J�GH��J�4�f�n�k»����2֞�Zr�v�}�ۦ��g2��SkRI$�v!�JI 	%b�6�r�@���LS��C�hN^�dΣ�ޞ)�'h9U�a�o)���.�E�մ��H����[�㗷Y�]���D�6���G�ocI��k�gS�v�c�v:N�.�]{��[ODs��t�8��a���O��7np���R�`��m��=���֞D�� ���<��<�@h�ۍ��u�T�n�.wZy�n7��r���u�[���ا��K;s�x$uq�SZ�x��θ+^q���/�6f�X眶z�T���`�A�Ж��Lnu�N�p��y:�9��ܙ�e;]�N|�C�6���qk�Tt��\e�gk:�+�ݛxی�]�6��9�y�vݷz��==g;��[M��1=��<����xw;��u�(�����[�ۓ���\�ֆ�����x���4,aۛ�^4�;�y�Fs؝�*�;�p�;!�k���z���Tu�	U93�����=��q�f���r{�H�t�cse`�;s���=�Uml9��m�{\�a�Y��"M�Ω;<S1bθ�uj@�}�v9	 �[�u����c�m��۰b�e�W��>5����\;<��k���g���W�l���u;n˹����z��mJ�ָ���1�];�`:]쎳�+��I����q��v�[���aE��tnP�&M��9.Hږ������nnNݮ�6�ڸ�up�sgdv�۰v�8:�;�5�$��ֺ	ɗ]q���5���::#v�ݺ�4W/([u�<I�Տe-���L���]������n��n8����6�F��7d�:hq�2\�ql�j�tD�sW�f��pi8ڰtn��u�{���w]�=�ΙY��Վ�qkٷ=��p���U�e<��vYd�A�d�v��{rUC��m7�.+��/@ֺ�ٛ��j3up1��Z�C��{98۳v�cc�Yŗ{v������ٞH ��cW[)��q��L��.�HL�q�[a9�p�Ƴ�*��Ql�S0v��Mh��0��lO�o \�������"�366a��r�G�1���*m��>]m�>�GX]Y�]����ƕnݓq��{R\����#.v�ζU��F��	�XËr�l�Ǵ�]���f���\Kf���7�=m�M�v�75�����S�
�rN�mʡ��n���f;(tkiݖ�S�ey_h�\�#�+���]&��۬�E�7&���u뫵���&�q�Sȟ�_��[�e���P��uS֮�#Q��WN�������3��Ayj��y[��毲��I��U{��ow��^/2�J�+=|/QR߈����r�25J�oޝ�ײ�ׅ�>�<��u���p�\;�R�.��׊���M�Q�]{|'�}zM����Z�N����bp� e@����J��7%;�,�ZxM)�ڠ��eQ���K��1���Ox�R#qU��o5�<!�ȱN���u��a1�z���ҵ2%�L�9��Lx4����9�5��ڦ+��,ʟ{M�P��:�vR:ޚ�ك���<�Һc;خ���!��!�݄�:��=�]���!ݣ[�~�Km��V����Mw8Ug��������.]w-ĬD�P����y6U�����o�|/`�O2��ד*AV<�%�M�8+���Ɗں����+]]t�@]n�8��C�#�����
�і�{s�xL����6������Jȸ��MW:�)�x�7�+�	�{r�����/�P����ڎs
m"��S���h{����Ք3�$y
�D�Qw��ȵ���"���O�+fʹ���o-�1�
�>W�(<�U���{�EAV�=�.��w���w`�x">t��7Ń�/+�ݺ�b{��zT�yz��D�ޡ\b���Y��/���VB��rP�&�?C��td�-Dk~n���v�+��V�7o_��*:�H�q���Z���o����X�1J��ܳ�T�UL)���݉{��3U�(��<*�:>a�*��� I�G�M�m���W� �+��ey���7،��`��k2���4hb��.�SV���?\?r���-�xͷ�;_��C��{'W���>7;-���Qh���7��B��l���N����ͪF��t�����7�<}�9���Y�%�k�W����|�$U�'Y�YWG*����I�߾y��A�IZ�N�� '~�`�ur��#] �+���9-�.w�f�7q��[�ک8%e	�s�̓�O��[����������}�b�����Nw�1�ZF��v9.�U����bH����{��:Ng�֛W[횋���D6�W-�.�s+�]�gΓu�������/j�ޙƗg���ԃ���*�dPf�y%�9�V7 }�������4�ǖ:���Q2�_ւ�s���Z �x���X9%�6�Np�{�S^G����T`t0�ey�����@��S�Ig|�������]�KT��e'̊{n�W�XR/z�'v�++t)��ǈ���~�(���Z�h�tB͗+�wmB��]ʓD~~�	��4��R�I�i�/��zZ�s�q���u|����*���g��9�ZED}�_$�]cY�"_n�z�e�WݓkKoYŇ����z����䥚�`�F��Wgꂯڣ��x^@0�Nwh�+��̩U�jb����s)�Z��\�����/��ِ^%���L���i�U�6�n��I����|yY�9|���}�pg��U�{;=�)����{�jP?/������7�U�3���Y^�N��}�����x�����d�OײN^���#�V��zߜ�G���9��j���DT�
Qk��*�N�44�\�>�\�A[��K���=���G�(v{*q������c)o{���.��[��T��RR5�s(����M�������E��V�	��o巾N<���w.��zT�$N���ɚ0Գ�ѷ���Ww�f2zf�
�U�<�]z��
����?c]���N��|����m�'#�q�;�Q{���wł��޵��y�`���0!�i���	�6���*��n��W����OY��f��/1��"Ȼ�I����3�]�vm������i �2�W�G<Zr��أ'�
��5�赟f�fuxRo�R��P"����3�ЩkU�_��m׆����K(Y�Oӷ���	����>7��w�=�N����|���n��8�Qc�N��O��U�zƛ��J��Q�Tv	��a�9H�=�fx9�uU���f��=h=�eW;��v���ڽE5um����oy����5���V�Q=;%JT.�b���2�����H���]ޑ�W���eZ�����F�z�ub�'	K��7�k�3;Η��

�nmKc \a�t��۾U7�'L�c0�Ð[9�=�b��i��+lj�}k=�����ū�9��>�~����i_}%��Qs�V����yϝ�J��.k�{�u�S ��Ӵ�9�M���//L>�]pLoHP�{2����ď� ���Q�*��(�����Y�Ƨ'����g(I��up�qi8����v�y�
�2���h��>6�ҽ:���O0z�>Tc�������[YUR
��_�w�
�CG��a���ƣ�p�>
��w�.~�Y!S���Ui���f�Q'��_��tUvV]֝�g5�N72��GJ���&�tngJ�q�Cy`�r�UdY0A��|���w3��d ��%[��{f���Fޜ����>��l��o�QG%Lk�˱�ն7�M�d@8:Q8�� ���=�ŋ�Y랮{t�I��lI�%��88x�7N�����Ыn˻�^��&{���9${,��gnn�'\yܻ��\SzKu՚�Ou��m��O���{��]]�1ѳ��<�;gN޲�Zs�ۥ�:۳ݝpf���.����x�f���:c���W����vzx�c��ۛ��b��w3�7�L�un����e#p�* ��ŋ����ڗ�mP��+��t���F-n�+m� 7�<<XtvW���z�O��
�S��u�3��~_����Ȣ ;��^9�[�7��L5�;gM;�����X����[�O9(�
�u�u��G�zQ�YMNlW���3Y��$%N���u^@�.��>�&�Z�V�
����iu����x{�N'�����w˙��m����UUwʆ��{Q�Nd����ma�c*m�f^!)w��Kjj�D]*�H%������G���@C��{��7�;~V+k��Mt}6�����4��f���XUi����JwT���5Lh����g՗R^C�$���`�Y� Hճ���A���1����ؿ\��R]��ɵ����?I^����۔j�̷X�����{�Xp<�@Q��]����dSwEN��u���"����t&u�1�'`+��d�9��]k��>�Wova�v��j��s>���)+�d���ghT�B��S�����&k��;Z��S\��o/���Z����X��>�"�+U@l�~���OT9^̾fxQ�?z,������:3/��S����V�-��[��^\��p`�1�YarE��R�����|��!ׁvTS(��=d3=�4j����Yb�Fx�{Iy��+A�W�t����)��eyI����\�߈�؆ƨ���{��}K��ƈ�w��U�����M���6��+�w;X(�'�ix�[��&�mz"�mj��L
�L�[ �|�T�Vqo�B!(��ũ9ϰ֖�]}���g�g���-[P|�(�J�/��`4�^Y_A�DU�"
�ܺ�V���=��9����j�L�����E���P���^�|�[C�V��[ ϶�<A05�OMk�|��,��2�o��>R�y�=G��hOe�S:���f��b�Cڋ{#���.��~�~��uמ��7�����~~���;>�xܧ�93��n=v6��!���!��mʖlb�;��9Avv�B���W!^�+۟7�������Ƙ��Hz�2��2_/��"���]�)N�����ݕk�)ù�E�w�/��e��b���i�UJ��5��B����y�Q���^!*���C��u��bAO�(Pc����g�s\f�<����Ծ�J���(�<��OO�g.���aH�ݒ�k�j���r��x���%d5�
F�wo��ʙ1/%s@�-�)V5�ƴEj�ˡ��V���ub3�p��ْ���Gd)�9�^|�J8h˨Y5���%d�tK����g�B�v>�����웜�����s*Y[�S�q�f���r*&@ ,�X!i�B�����y�n�e�8�]��Ȓ<"����g��j�6.�斓zs,ҝJ�!%h��C�sc����.t�I�_�P�>E7�Q�4fdb���+�=���f�Uz��ʱAT�é^�\�{�{֩o{�5^�=�0�o�%r%j���LR��r�V7J����8��ع�bsv!RƬc��6Ϭ?��ַVŦ5�>x��B�K���y���Y���\��݇�)��*��2R���W,«�{1]oO�f�5��\�s�*���ٮ㝦�\�P6��>ۣY�[}�9ƴX�-59�Bu�[� �mY�ǂ�k˟��K�'g8�}iz���^��hy����I�B�w[��>�t\�x�����ۃ�՝�xB��g�N�u�r��}����h��~�����ݻ�@�j��::j��������v���F>����Z�Qi�P
+8���fyx�
�H`������I�ɊP�-
�_9=����{�����}�����	v�&�V�FC�S�:��']7y[w���{cB�M�zJ-M��5H���f\�|�-�3x���Z@��&�'F��}Z�.�昮�x宻�iH,��_](K�r�F!��)=�%r萴VQ����j�$i��=�}f�Vz/Y>S�^���̱�/x��Z�XMA���c}����(��ׇ�N�fx�J�b�oA��9S���WH�ƌ�p��޺�ɑ�d4�GZ�9ѳ��#cݬ���1��G\��M�7�q���eG��];v�����I�����,���vn�R�#��z�h.{\����5���ڕ��o.�p�,�`�x���0����6>{Z|�5��_�ܥ�<:�=B���d衸N���u�^�AR�{�	Y�H}rTO�e/��!�B��F�uR�U{������ʳ�!ɓp�\Zx�Ѭ]ŵ����h�7���6���{g���5w^>����]�	��QͥV �N�=�to厖��d}��ӎ���M֓E��3���w����@8���f��p�)��IW�
�˽�>6*e�+_-ad:y����[�v��PBj�n�'�&�_4����Ӽ��ªnz�\S����V��=]/<-z��t3��+��V��5��o{�+�h����S��"`�׍���X��u������'���)OI����ƈK[O��,`���$���ҷ�u��A������&z׀,��~x�]ʌ����8^������,-  ���q���;pn:���7�0�v��m�����i�<u�[ 2�z㰏��s����g0un�v;����uì].���z�gڎ��3�4���`��:��s�n|Vix�%n�v�q΃����z5�)���g�F�65�`��5�l6�rJ�S�c��x��v8���>a� tr݁�ƕ:�{y7���y��N�<�����y9�d���Y*"��q��g���9�\m���7�%�tҟ�Z`��k��5ONTRj��̭�.d��oK�ukCQ���R4ǽ{��}��}t��
$�Ri���}�'e�{l`>�?���w/V}�M�����c}��:XT�4D&A��/U`��e�Tw3L��A*=�K>�n��#��n���' ���&�i��d0��Oˣ|Y�z�`��g��ɩWЯ	nV}����h���V�&�JB�y}8����y]����'������� ��BA�ER1,5��b�-Ǩ��PV�K=��޼��jʽ�{��j�]2T56�wG\,	�q�(Y\u'���ՀԦg=�ƘG�v������O��ٹ��1�����8���H����f��^�mb�ycy������`A������o�H��O��3)n��ߟ�����+�ɮ�tڶ����G ��v�Rs&��ڲ�u��lk�#_='��~!Gr/~�3:C����w�^މ���"���Y�+�z��.ngQG�W��]t��;�4�NZ\mQT�%x��z�|_h�,�Z<���`�ml<��a��wK����]���O��:����Ʀ�{Z7�&ʻ��q;���b��;�wyQ���dH��,^V�a��+Ώ�xg�]O�����ww;�ߝ�����W2����i�z-]�^ѾU�R��WR��i�,�SW�5����̩W��4�S}ݛ�*��NP^�R�̢Ͼ|o�r�تĨ�b�_r��/Sɿ��W�hm�Q:��X���Q�L�XU��]���}�����A�Ե��'��T�Bm�=]����Ѡhx�ڃ:i�Օ����_(�� �
T�M�yY���>��>#f����m��dA��uY�ҭ�;���#�&�����_+H����P^��(�sJس5#G"]����BU+��vZ�ޡΈw[Ct �:ݺ��:Gn _b狤�wnR醜D "���\|泛��˓W5�����$Ɛ�»�����55�r(�ڝ�o��w��z�E#yB
c��US����;�兗�������E�I:m�H���{Mh��6U�Lʘ�gWOpB o4U,k�ù{��66��t��t:g�;��Ⱦ����{-nE�=�S�<a����� �������>�h6�%��xT��M��Sxv8�"��OR�yރ.�o}_o1M�J�eO�)(�FW,9���h��&����nG�Z�&���bj�3;;)!�..��onE�r1+���GI�V_<��`�x��T��	a�l��v�j�O4��Z��o��w�����r��I	���4�W~ODgnK���G����y
��mk��G
V�{��#�����H_k<�2����Ǩ�Oi�ֳd�ղ�TŰ��v�+�����`]�Wj�zn[I�Y�/U�9�t>���:q8i��÷J�g��sι|5+��i����7e��-��ヺ���r�m\���C�n���DڹN�+���fͣ(к[L�x�m�����,��b�׸���z���]�n۩����.�L�e:���O7�)�j��0;4hVؔ�C*��wr����tͅj�e{�#T��>���2b�e�� ��(#ց�6�s������sk#
��72�{G�� �H۱�F��j�Tε�m����՝��jY|�V	f�i�{�.I��M��ݜG;k�@o�V���Җ6�^]�f*�_jD�Zn��������f3|��Q�Ǯ�-:�^���nS�<���7#�l���ڧq_]3{�2��Z�9��&���hbZ���*g*��һ�m�/v�>�]���]�9j�$�쾧W8:����BPu�R�u5U�k���c+<�)���Vsh�A�sۅf���x��y`�H�4�\y*d]{R�K��%y�Č�L�{+b,G��G>�h.��f��9�X�\�P[53u˷u�0�J�����'�jЯWp�M�+n�`����Y];�[zjv��^��B��Q�4�I��[�K��b?�[������'�#ɂ�nW|38W%�QG<�de�M�^���/�$�ٜ��s���f澙֟�*�ʂZ�啇��3�x�]�Y}2@������.��]m�"���wWy@��ME���ϕ�Ȧ�X��q�+nz"O�������KN�u�k�g�v�nS�hA�\�7WV{a�g�^��ܹ�ȯa�,'g.|��]���~�~�f���ڌ	�'���N�ӻ�}���e���5����MyyKl���h5���K��{�ю�����͔\���9��ԾL�As�Y@�ɕ�=��C����^ܽ�������זpӜ~��R��0����}3oK��������=�i��=$SPq(�m������b�û(���j[�2�mxF�a�U�;�F9)��w�ϛ}�r��%Uuw�w.5H�Bt�*ʿ7�%�v�׍塃~h��Y��M��k���}	�X��z���=���SA��/���:�J{���)^�SF�Գ�2
�#�Mݻ��.����>%��k6yܰ�yfXd�������l뫜���Z�®�����
y��	�嚎��Jf��MY�A�B@���k|�"3��7��D�ޣ�4��E,W[�7l�SA�I���x*LS�S�^�z-4�V�}w����3��Q�0:��Th��5����4;c>#��'Len))�r&��䎶ˎ^�F�v���y�����v�m�(��i�Kn��}��Y��݆���Ԕ9�Wim���q�_ѳ&F�m���o���*5�\�V�h̦�"�Һ��{WU�v�\=��t�I!�h��ݳ]��#+�>��T��Ă�[��;�u�d�}˪P[��ݤ��zΧ�Q�*x�@��嗀jܺ`*�U�`�1sOnG}[V r�JLՕ��Ck���W*��7i{�O�<Ѕ�[�ܿu�ԯw���SaY?O{��Z��u�)ƪ�e�T���W`�ro݄Q&�d
�4PN�"'�u�tDav��Ne��u��?&�X�,{o��)㗘��f�_~>�\M}=�t'��������U�����>��@��R��%�=��r#�*�A
����Y����V��8�̋Ʈ��u��Pe��LB�vgeN�}���T@�=o����~�`�s�`=G]�ֻ����c�� �u�e��k�]�%WXa�yҋ.me[�.��ܘ�,F�r˄���걷9�¸B;Zj�8��H��w��M�����s�h6�%��ol���۞g��oQ�vh�q�&뗓��x����ε����n���1�eojg�ɲr���3���l`�9��ݶȻ��N��\�n1��a��q����R���gG0�
� wf�]��b���v6�λRcx�*��:n��u�e�ܳc4�v��\ݚ�#��]D���Z�e��ݛ����b1��Evn8�^�nr>��wMG�����b��1��}5���9�2��O�]Ԫ5e
h��J�5���⼭r/!�W�=½/+F<XHe�R�]{^�fzye��m��֚�a�k��+��wS���WPW37�L���Qwu'[���D�_Eo���0��wf�Ń�y4u�ʾ��[�>A���ە��eU���kv%^�hY�{�[O1��>Y�~G�^�.���q�0!t{��uEZY��Pܾ7��
�#�5����]���8�y��ˋ�vM��Q�X���x%y�+��rЉ�1)F��KG�1mJ%ATl��{M=���F�Ώx��hH�cӷ�+�x���z��X�)�k���|~"�ϋb�7���LX�$�ٺUʋ|֓��fc��3����xI��&3s �;�S�`��T����YX>'A��LH���9��G��(��~�-�f��r��<���77n�c�tɸ����#%v�jG��vW,v���������R���\ee�����7�|�!~���:~�
���ߞ�c:GޮU�]���V;Ol�Gy�;~$*HyS�>D�'ֱ4X�d~D��t"��{-�/����߰��*��˵Ԕ���Y�b3��m�N�U��,'�� ��W��r㛛�u��)J���~T�Mtʹ���ǽ���������<�֬���/5a� ��U��r �
a����R��X��f/x;���E���4�_��E=\+X������r��q/\ޟu�,�3<����I4:�9u�K-�+�PI�>�8Hf��f����_CG���Fgڥ��.
vL���u׺ܫ�(Rv}�S�T:�n���˭cS����f!y�>���e�xTh�	|t)�ڳ��"� �4�ϲ������H�A�s9oS�<;�)Mu2��&����%�a�aw'��J}x)���:ӽ0��Q��K�4|7�[���ϛS�u�G�NwF#�M�y�;cn �n�t��/,u��۰-׳����s��F#f��%D������~��F��<?^[��H}�V`��Ɗ�٘%�y���g'$
���)�(��>��GS.܁%��s����osp�4�ݙa�
-4�k�q�L�>�`ܕVR�N�y[��F/6�՛u����.��t�ЦM��>S��_���挕�A	�J�Ĝ��l�_k�N�4�Y^V�[��Ҳ�6�M�z�ɗ����ׯP�YG����b�ڔg۫ up�>vVwX�(��I^�����3�⼩	6VZ�r�S�-�r��\۸�t��ɶ��
�"���%�Y��>�kմ�x�hl��^���S���^vU�
��ܧ˼��M�ЅE]Dzܡ�Ǜ�w�5\s�߼��MYJ��B.��n6>u��l���RF���i�ާ��ok�u:��I��L�V�*��?�X$��<�e
Xʦ�C[��_
M�B�Þz=u�q�Ykd�89iW��]�s������@�`�ܮ�'�t+�Zލk]m�ɾ�{����M����k2�����k���=cN_M'2����)���no�|�,۰�5�W�񨰦���uv��/o��gHh\�4�C���I�pU/z��e���?>���	T��]��vZߍѷ�#�;ݠp?mzf������8�ْ���(�-"�u{���}��$~�E[�묝�kӌ.�X��<5����_[��Q�����ˬ�=`z��C6�+��
�E�	s �)ɟQ����E�ն=B�ԏ��}[�z-�̐���Q�ֳ��4��lϫ�m�a�ʮ �_G/���׋R�^e*����oUS9,�2�]_�]C�X%�(Iw�:�w�u8�F%���g�ި���-�S���v��o���"�bc�w��+�!I$���^���_D�r��/5��λW�7���^�[�r��[���}���Qnל��!���^�Έ�C�Mһ�Ʋ<u=��bn<���0w�����r�pO�Lg`�Ѐl@��Ҝ��t�1�����?[Y�o�4�?q�tް������ryz�jO�^�TlX����BbҲݶ���Uf�%[�f	Mg��b��л�\��*�w?���L'n�n�� �m\�JYP���0�
[�����#�^kǩ��Uሯ:4���nt�R�?A��+���4FX#�W����;z��K�o�>�K���HeQ �A�ԳW�"���������~G��;v�*�<���7���$O�O��1f��l�<]��G�  �4*�l�V#��r��	&lڽ�~� ��k�q�f��c��+�M7��+����w��춹Y�a�K�c�C+Js�������x�,	
e��%6�g��!\#�K̂���%���M�"�V7�+|g�Z)��_&8�ʋ��}.�����%��$k���]� �σ��Sq�VZ��`�d��kԯU����H�{��d~�6oԑM
��ڜ氨6���g�.���%|����hPN���g]۞�mp�m�y�x0Y��]�=:���snw\����R�u��l���r��;vۚ3û7�sWC��ۇWm��=,���3ٸc�ՠƸ��wu�۷��l{Y����r<lp�M}�үl
�s`�yx��4箮��]]UGmm�F�onQ9,mb��p�q��&ζ+hn��j��*^����#(mh��avSAu۸d�(\=��m�ǤЪ�2�d^��s�ʞq��%.SMN�����>���n�1��Wrj�w�*U����$QO�_cm�,������)o���m��P0�XU�>(:�Bl&����ygOY�oo�wheo/i�eZ�P&�rW}�ʀ`���ݫ���S�N:[{9X�ݟH���ړC���Y�^]{��F�c���>u����t������"�����{�bWF���/->ʛ��N�v�
�Uz���I��띆ݢ���w�#�V���h�ց�6J���?�q#w�W??9W}����jY}�!�zԠ�v#מ6����й��<=�5$��h٣R�y�#�u��I�L�U*	5��5н�}���" E�����K�rH�<W��C!}����r��VΆ��<g�efC⣔��`��~�:e��X`��4���;vv�lݽ/;v���;�'i)�X̊Fۯkv�,���L��a���"2��Z���m�k�m��^��x�a)zVN�	�}�{��U��맞����7����Α-z��%-�-���a�~����'_k�g��y�]�����.�o��C��k5�ҳ�uɋX�u*�=sv�#{�/vpS�+�{���R�t�
2�������$9�PW�>2��[֦^�l����yW&�u�e?0���wY�S���K�7G�o'i���ʖ�d�Kt�%����D�jx�j��A>��ּF;�ٴFY���k�<�T���'����&I�*��"�އO~*�M��><|>�4��T�����r�9��W}̔�����W��!= ��:�|PPY���}bf!<��x�yݝ=˜[��%���zM�'�V��h���AË�7�S<�N�V;�S^v&bo�_�����~U�_)}�F�<)���{Z�]�:�Y�9F�Y������������V�Z�Q�w8N+ud�9���w�x��N�׫r��7Q�ո��- ��v;J/6,jp�}�ܬ�^E��|�[����o r����b��{.���A�R�U��;(u~�T2���~�~˒W%韝�\9�c���gr�PVK������eg��K�����6��hޚ�sr��=^�h���+��k\��}m��p�
�hs�����_Ox֍*�2�K�]���T��"X���7�-Q���'S�/|�ߎ�gʐj��N��CA�{�h4k��}F�쏲��Bx&uL�����0�l��b]��Ա��k�P�JX��s`��yܫ|\��B�؀&�������mv���~�̿V�7�k..�ee80ivzj�o<<>a�هݬ�/����RO1�*��E�Swz��i4�eS$����B�z@���*�	����8E�b�A~V�׼�SMK[<">�hc~+�y,�υ����m�n�����[g�����\�^|\�r��0��|ZR��f��j�N\hz�n�ōV۫gC=���{5��(6(��՛�Ħd�/9u����Fb�{{���t�c���y<� T���~ɬU��@l;;;!</<k���G�OܫVKS�A�R���fq͡س��W��WC0뎟z
�`�8�Ezw����)��׊����e�:R���t>��h��o�ee���}ֺ��H��,�.�6��6DǷ,�.e��Q�B ����j�e�n~2TF�6j�9�9(r�m���Eo�W3ٹ�����,t-�ۗ[C��~S�XC�7u�x�ρ��^��3���2�O>�(·�jئ�t?9�GiS������k�Nz�^�hK>C��W�I��0�X� ����i4R�����N��}�	���_9��@��/K�$p������=D�Z�b&�\���_�䨇�ǅC��/�b�n�ݣ�~c|��QPKz����E�m�L����+�N[]�"
W�i�V�x�*�[�ѣg6���g�9
��ٴb��nr���Z��7/��Ƕ�B��LC���E,� ���߽��[���cGn�{Av�����E�S�ɦVct�Wv���&V�*Ͼ���:�wQb��^ɌQ}�/3�5�8��C%&sG���K����۫��sWX��g����bfE)e�.�/�[qL�De��]����3�:�>(4<z�}�-�9~�ZFԴ\�j�m{�7����Q��JĢZ�������\[S�{�ca����"ޙ�+����1��e��4� $K��ۘ}|Z�[+^.���;ܴJ��I\YY\lu	�1�"�]X�����L������nr�<}��:�g���{&���~�>�Kɚ&��4RL����D�ۇݺwFS��q�`�{p�ы"��Q�R�i�"�N��^�iXc�,�����l�(^���K��qAJګ����/}����U�e�_�r�xJ�z�C�d#�2��������lOP�`��f`U���,`�G�+W�7qN+S�h�<E�����tR�w��jr���C\�y
�r�Z���Y�.@�Ηf-j����َ�%7tV�N���L�9}��{�/�̜�g(�6��� t���[��Ϯn���uhu�u�T%[5�^<�2R<ԸWI0���H�xEӫEV�m��m7f����\C7g|��"�����T��qi𱬚[�|&�=�gz�,k�r+'�r��7k.n�`�]�f������pXfEg��v�a�l��+p�]�N��E,�A��;q�g�0���7���x�9��2��<��hgm-�[E��uU����[b��'>��o��'OX/5JÏ<ձY��UX�z�H��I�1'�i&���&��y5̴�&��!Q�
��j=��.ǽ:�Cpf c�E#�`���`ڲ;e`ܾ�&�Y:]�Z��l��U�;�m)u��qt��s@���;�9&7�f-'U��]�0*������L��J�oX��������)M�Y�q}ԭ4��d���[3��"#�٥;6�b�.����]��[cM
����-����)��<��Z��L:�Bnz���&�K�QhFǂ����-��*΍ɓ����=۹��q����KQ�T1V^3�����7�����J[��g��K/<&b4�
yHO�F*������4���q��������H�F�r�m]+iVd%� �R�[��ֶ�;��{)38g>�s�b��68�J�ll)�>;#���6P9�v��6��9�a�l��l���ٮ�\)X�nh��ɡ;���[qcFw]���Gu�=vq�٧/��ǉ��v�[j{eѺ�hr��[�%秝ֻ$�^U���n;k��.@*��W;����0d8:�+���G ���\���v��<��x���t����m�]n�=�q������6�k���Kn�g���G�����<kq��q�]g��cʽ�yN�g@�Xx��ۈlGc<�r��� ޲ܝ�g�;��-�G��E<;��A��������}>�x�dC���]��������[ta��L�4hyˬS�k�s���eKs�O��!-cb�J3���G/gi��˺^4Y^*��۬u�ڵ�G��6�J���<��k�{�\�������cc>ڕ�`��k��up:�7)1�{r��W�:6������Kë�E-�vA�q�;�׮����1��=z�����a�ք�3��v2�V�"��H���\vݮ9�e;��64{n7���퇋].M�ћ]Tvz۔��3��n�cg��PwVWm�;�^]��v�C�p�L���5�W:�N;n3E؉�����y�.����!�d<�lK�Z:��vp���e�8�ÏWn����=C��2�xo]v�i;t�ۅݢޓ���';n[�����vΌ��v6��;���PT���#�v�Ňr���n���=��L�p/l�@�(��v�q��ӌ���n�gv�о���!���8z.�k�J�Ɣöֽ{/N��Ŵb�1�Mh{�N&�r��ݷj�v�z�f�W8z�+]�8���0�{s��;���;+sX󍹫�	j��yL۸�ܭ��e���p�x�q�N.�ԜH���n7��l;��ۈ�Y�-��6��{-�A���cgO�1pg�:���Iؖ����R�ۗ�6vz۳��\7=y������Gs�f�cbu�!�n�ֲg����p���tu�wi�q���O�S�<&7'q���t����E�q펤CN�9b��9̷'k�;�u�/4�i��!�z���������a�Ϣ���l;�t�9�7y���Z�����95�6��9�u��J�5�k�^�݄x���[�
y=Ɨf��3wn��"͑z`�k��.�]��s������#K���>���뵫θ�If�\�}�a�r���i�"��0v�-�����O�j5i!��;�Z�P��t���֥�^�X+0���+��5�lf�`W�x�����z�3sH}�/y%���@BX|��=}�؞9���|eEZH����e��\xceo��5{�~&C_3Zy��[cё{������VY����ṨRG�zw*q�TZ��F/���D�]����[��Y&E���D|{y�q�,��h�ۣc�nEl9}�uN�G�� X���o�x������+���:�S���2��������1r��ID{�ZxկG=�iN-=qIG�#�V��]�d{hms��enw���� �U�4�*4��!�.S�b�>�Y*�O{��iRPY��t��̓s�`�4`u
Bwk;�����2㫹��l��A7S�dA!h����j�U:s��	��o����!].W���R�̐�0;�p�/���ҟ؎�⚙��ȱȡ� [�����7���N�/-
�φ�����!�ݳ�8̈́��]^��Q��������٤��Z�j�+��,V֩��/�fgu]vc%J����o�,�{8 M�,�^���gԲ=ڿ��1k�\s���Χ�s{�&&I%�jIZ��U����o����&67�)�WW�����M�n��:��VP��O{�o��h�X��6�~�R�� l%�x_*B���*�����m�*�۔�'c�%b��M�gIW��z�f�y�'uo��S��j:�R+נM��,���T�I%e�s�ZGrTi|�-���No������Eݻ�	��C�,�/Kjb[x�nYx\w�C�t����Yt/㾍��λ�L�;��mu��>�f#T5d��WB�[�+Yl���|r5���<g�wOn��ۧ�V=�n{t+��c瘳�Y���?xEQ�����Fg��ia����}3|�ૡ�l��6`����f:^�ڂ�{��*��em�F�%�,QXSEi����O�G��Ð�]��$�4���ˡ� �}�)�O^�����N���ev�������.�7�^)HF}�Z���5��n����z��g�3C���/_fGس��GN^�������͍{�q��R�y{VG��z�K�<m�^��p��W�M�4�讽�km�#�N`�f�#�;�B����̩����>yiŘ�et5�.!�b�[$ª�*�r���{4��ɢi�e:�������*�|���*m�=�x�l�!��'��(:�F�ovT��!��g��U��7���� 6�]v�	bH|6�/�M���&����w�Ԣ�I�'���ŗU��/Gӳ��1J!��u���ō��켥��J��	�)8��me r�����`;��y�΍Ґ.�;j�hݎ,�ϛ����w�t%=��5	ʱ��v���p����{{rf���z5i�h��܇���?{�[��2�����A��w�閝>/�;�(a��@
3��_���|�]X�v�KU�j�=:��ue���o'�{��7i�EO��%n6�\��B�٥��{޼��ݽ���t(&@i:�
�Ձ )陙����̛6Ũ��x�ֵ�k�^�z�9DA 76�Ŝ�|NV߆R�����e���{S�����,p�Z^��w?8��9߅[S6���NW�G<\�J��4d�ϯ0w�]�z��,^��(�	?'\�{�㩐����2��p��hf��0R��O`"+ՙ�n��0!�+7B���Ӗ4!�
9x\'R���lr�p����8R$��AR�Rc*i�+��T]��'� =��A���7q�,{��Cَj`-ͧ����zCw1R�z��ޞ�39)]zy��s���)�=�)oҎ��'B(̪n�[/k��s�ԛ=�z�u�۫�»��8Oe�Z���u,����·|o�Z�>�Չ{E�h�>�{��8�d��+uҝWr��g^�_0���~՞��n��7�]�~ם�NXDX�����ej*���o�˯�o���2v3(;}�r��*$��V�[Q����Q[}� �z�'1Zg��7��G���7�WS�
j����6o'�<�w��.+�Q$���2�-���B�����9��e�}��`��4�sc��Yn�c����<�
 �KA��ԫ����午���M��{9<���_Z����I��l�]������K���ro*^.`����.��>|�e/���M��+�T���4�Jp�Is��x�&���o�G�8K�f_���3j�x�٦F$'���(�ڒ�cY��Ռj�g;|����J��8LK�,�ù)�U�GY�����Ԧ[��7��|4���)j(�~*V,�;7S䛘#���yw_N��m �7��]��[��w*���vLnEu��ݳ��q���-��ܝ��P��ۿ��h�R�vA�cll��ҙ#p�ϓ��pOm���[��Btf�qѩ9;b�3��V��9�.n�K�mvW���qع��<�����ݨ��vM����:���K)�Gb�S#��!)�#>�3�J4]����x���枱�E�'gv`��x0�;�[6=�Z�7`�G�sӘ{&�3�ls��f�n�m�\{�E���z96�+?�q��������W�.����!����.��Ɗsrݧ׾��H����+�g��ł
��9�n�>�W7���J� y��H�)$�qD��?	����QgK�Ws�+�T/賲��Ɲ�-�o�1lZ}�H�1�[�!>y��^~��ÿ:	�Ra�A6���{<��vǹЙ�PF!Ӂ�`��:U�=�A�6 �9Wl��{�=QT�8w��5��ŭ,?Imd��-m� �QH���j���v�s��ϴ(��Ր�/���?��)�X��x)�;w���^W�=��VL&�e:	�|�b���@uZ���x�G~�PVxm���~
�����������±�w�]?{�
2�U�w�Ko�@���wy&��r-�-[X:��䍸��b��s�m�S.�N-�h�vu���)�׋�xa9���ĵO�So���Gn���nx"H��"_����ſ��vh������ځ��z�I��alnU���pOc�MPw:v�u&�!R��g'a�f�c��j�_خPZ���*�o͐�u�!Jt��
�M�=�か����I^�NV�N���0�7=6��;A���"�r�����E�{���Z�ӿa����F�#AR>�J�zz
������pׇM`��Zz�����5�l2Z��
D��lC#�:Q�{��H���v���ٿs��V��7M�b����(�1+pK(b�wk��'�u��IӢ��Aq�1
�Q��f��ӕ�;���}��N\1[�ST�SA�
��ڷ?i��g�m��z�����Nx�57M�Ԗ�!��/�b�$����0o<2��&��~����}�0Z���/"���S��%�[�Au���NF�Ø�:xe;��"/\0c<��E����ӡ�<�j��pI�������	�Nx웝[�r���*�t�U
�Q�"�_s�s�׾ȯɍZ�jDVy�N�����X~I�ٽ�D����W��M﫦%��jy�����կ\7��/�!KP4O�����.��+.v}���Z��W-wb�b�񠴡uŞ�Ӌ/,���rK�_	�yz�X�����ګ����Z�+�'�t�Ӿ!˚=��u2 ��(z��B���/vS 	�ѩ��~A���2	�`�s��iOc���Kj�!��Ɇ������ws30�ĵ���$�<2SkN=��k��
	�2�!����?;�Q�OՎ�q���)|Sm�#<��whй~'��i8�-sgvV����R&���u�m;����w���q����#6�4W�}�[��"�"
�Q�}W �̰�%q�~�����v�ڧYa�{_�H�1�����Ŭ�H�V�f?f
�a{<�t�!ܖ�>���������E��1�k��lk��i2��i��{Du�s�V�iT`�+�p�z�۬כ;3�W��٪"K�o;T���	�x���;=�fZ/�'��{��M�q�R�Dg����[��� lB,��5��z�O6�{�7� �y�Q��E�Ռ�Gy�3�[m�ѡ�R�,,�%�~�ײQaM�MPe�����T �h�f�����F=_������=�5�����!�"<i7Y����h��ݩ��w�縿+�nV{������H (TD2����S\�eH��{��ھ���v���=�Qwj��º+ݼ��)'Z���m����U��ؑ��J����wC���w��=6��/\��F�-\�Hu��+1β-]���=�OtP�Ь�"�\��R�tD��wM�}{�[X��@_�iVM*-����h�ۻ.��3�gvg�y�-R��}��7��}gJ)Ӯq�t�Y�z@��N�W�rz$=^�x��Ϟ<<�.�SM�*��j;Z�n�n�3����[`鍬�����B���%ݮ\ h
�G�[x���˻�<� ʍr|(�J'��q�����{�;"{�[~�-?��������\ӌ_���Ӫ�ejJֆ5wϷ�w�WP���Nr�-��3u0����b�e�
x��A-$��0���s�s��y��7����o��rk����MB�*�/��m��滌�#�j�wK��O���[U.^z�.��`K�|����v�-c��r���,�sO���������	�6�u��>=��Z����� ѡ�����ǵ�=䬎fR2hBᎷ���<�����gϞ�eiW��M�K�iӤSi1y���|4G��wVaKİ��6w���J?l�?G���^��Q���������z]�W��,��:�b�������]Z@����GA��r3L&u�:.h��	T.N��^�KQ:�	��G��)/��Ѯ)p�u�D�����{Y���1u���k����;�*�7��$�<+�\l�Q�w'E��^;<,�Ldѭ.xig�D�h��t]�K�/�|���(ٚ܀�ny8'��ڹS��i�M��f^i!N�'k���{y�+����8㑮9��m�r�z�Zy���LX�gWA�e�=� ��9a9�3�ڻ��;,{)W<\=�b:�����&�͞s���]k�u�s��ur[�R3���]<���lmw�]����Z���ٌ�?������V۔au���o}��w%�<����ney�v�q��tt�r�o�5�[��qz��R^EbC��W:~��ξ���}Ⲓ'Û����v��r�Vu��1&�卺�N�u��/{m'���!f��䔇��2U��
�M6B�3غI\���o�e�zݜtspWzAv\V�a�N�ͱ�Zz��H�r�p^X;A�Ŧs�{u��iem�ғ��X��k=}�;+�B����R��J[��7��k�u�W��^/���z����鹚5��7�N�vk�֦s�o��� Q�@��E�bW��_7�j����v���ɶ�K:[�L����E
C�j�y��K��Ó�wVn����H��D&<����]��[�&�݆�v�SW^�ѹ۷e݌;�%��lv��R������:����;ً�i�:�^�8�(�m���o�pR8,�6�e���{�x�i0A��9�Z��s��+F��s���5��vp��9��uǞ�֡УR)R�{�!�s2�)ѳ�L�2�%b�쏵E���YK*+��RdJ�x,8�]k��#h���vl��ɗ�c^����=��<�Y�]ǯ�y|������BK3��B�*o��*���.�h�,�DwI���{~G�<�tNx��U �P���;��jn+�U��لz���b1�l��yմ����@��%���#�_���x�t<������h�7����玕�T3yO	E,�(wPR�|���rv�ߗ"!�]���tE.����D6M2ټ��I�[�c}y�e����U�Ɩ��&��e�������Vq�ܵ�Y¼<��)Y��pW�g���Q�F�	ݾ���ż����v�b���="jڔWv�\�;;�ӹ)$tBT�L�g�}[�u�LX]�v���Osvc�7�}s�\{F�3����w�X���#�{}H	/1y��%��@4��n���ɩލ��9z��Z�F=7���<���q��;�B���hm����I�]�����k���{��Ƨ�z=q"ޥYD�@ ��1��X��*d
���s���p
���n[��M}A�7�C����J(�ݩsh��i���v����ޑ��د.�	�[���(�T�.��[5-�t���-�ჸ��E�誆=�N��� &��|��?��#��^��U�]o+�K᫩ckn����ڸ�op��~����6��[}p����M�|i�,�sQZ�.����u�_]�;�Џ$���f�t-�*��.�Un���R�v���azY�^���?f,�p4%�EE5.@���d�J���V���z�]Zzq��o����^M?���-fAWu�o4��v�IH��wCMn����nO8��Pn�W��udpQ�NU�VF�κP9,��l��IW>�`���A5����C	�gg=㗶yX�\���0v�GqC3��q�WvN|[N]&�8h��Q���3�;�3!<�v'�����n��敒���e�㜹0��
�2�4�ހ�2���;C���@�l�e\�y-�/E�%�WX�d�z�_%/a�PWNMk�*�l9uj�rޘ��L�����u��k�fYt�x�逾zY��;���J�Tr8rO���L y���K��
2�R�=5H^�g��z%YY��-��%n})���q�ꑖn��^����&�����>��Ay�	c��"��4�p���uhG.������ݼ:mr����j�u�B`���l)'q��\�Jw��q8��ۣy��PڮF�(�]��_v�J�LY�5'��c&�zVZ��	�("dE&v��=\X��GKC�YL8Qb��7}[��"�8���`������ir�=�(VX+������D}5@�r�EEv2Ki�[7��Q�-Ѯ�_��b�Qy�|�Wx��\������!�[�{�q�q���v9��rB_�<���]6���O�H*�b�i�-�ꪱ����8z9�ɤz
VW�L=��v�Ϧдpظx�.z�w�!��1��h�!��=Z���k ��ש���eN��^K��<QW{|6����?X!e����p����a���^��	��~�y�ⴻ�R�(Ղ3<=�-4��6f�_��!��n�y�Ar:7�z��h9x���S�ο^k�z �,j!�|ᬼ���Z��:�Pc���Q�ه��y99����͸���V֎����4=�-MS߯�#�����@;��n����s9밻'p�P��I/7�V��˱�C��L��w�M�w�����<�؊We+<t=�`n�/���vP���ɰ�G��V+�evhq�y��t�~�A�X�4U���ݘ����=������)ʠ&�TB�LA�y[��m��w�����c���L)}�zߜ�8*OD��u�$4P7�ߵ��Ξ�^��F�h�LUG ��q�@И�Y��Gqv�����N�;��h��� �:��|���r����ӯwc��I9nh�����nbVv���i�\)竜�Q���c��u�s˜��Ãm�V"�ǹ�����N+��Uc9+����iyv�VX{U) �����Ķ*mx&8��6��K��d��W��[;�j{�l�P(W%E$��
gӵ���ˮ�]�����p[> [x�{Tҍ��m�B7��Me��ͭU�3�=�j�r1�]��=��h*�MHKonM���g�R��3ud�*쨓.� ��W��c�|��N�Vz�t@��y���%X��ߌ/���"����M�͠�^ؿ~e�o�]���][�ѫ=���N�Wy�=�+SN�w������.Z��6X�����rQ�v$��.��o�H��idY�{(�a<]/���N��z�^�X��a��vk�CR�(�W������7�& +�!�6���&��>��,��s�]����6\9
#O/Z�%vM�[lt�&�;s����B����:�2�[^s/G���`��Y���Y�<��
��^��A���jA��\�ԃo���z��76��n�op���kv�7m<��$��3�g����㞲lL��ix5��k����;m�� �6�)x�Pݼn�k5n9�OE���0��s]:�`�k.h�D��NprFu��Ղ{%�nʴ$�qX�K�~?`f�C)��G���.L�;=���N�1���q�)���>�ن����5�X��/|�=[�H��m�M���fm�	�P�λ�X�C�z�3w[�3q�ţ��w�to�K+qh�P
���~�2HfjLc���2�P��D���qPXz���Ѣ�4�2|�bQ��W�eL4ɿev��U�}ez�I��X�kF*����{Q���h{���� �7�v5���/�Huk%���(��'v<�2�)T�h����E��xӤs~#�9�Qm���l���7cG͏�=:�%J�g�P�P�[�"���{'�u��)�6�P�w�J�i{M͒��#�.��wM�	�z�XŻ�yL4��r�ƹ�W*�:��s�H
�Y+��u��v�����f����$8{ ���F�Qm;��Sg��o0nZVs�9�T�l�I���>��в0�
��j?g�B����_lv3g��],��ǖf��4 ����@�p��zf�U��s����S�v6x�tn�{�%�Mx⼧3����\O-v*;�\�Ql����{��t̑M5ņ�7��W�f'���kM��3r�Oj��p{Hķ�oz/+7K"p���&�恞t&��^�w��k|"�Q��+O��T(�<�U�Q�	� ��eDG
��ak������ztw�(������W�r[��վ�$F���|��O'�׵ÉSW�:����![��t}�[�ӻ߳R���3zz��E��[�sGAF�n1=�nORS;�+��Aww��+��)��^e�+��^�Q����$S@�KlՏpl5�{��\ѳ��⻝+���,���{f�ǻ��g�Ϡ�]��M�V6;��@���ϳ
ݭRJ�U����Ж���6O��vq�N +.L۷8���o�%M���Ե�bbj@^߹@�G5�̯M��npg�x�ʲ4�|̀�l��1���m�^�S:x�=֜lǚ�s3;}��Y���i�#���YIDK۾y�����R�Dy�;�Er�gQ����~�Adf��u�=�����k��<6ٯ|ϑ�	��Sj�	��g�4����r�գ��W�~7����~I=>�F����EY�mnq�CũJ��wV1p�7{g)�y/v��Iyr��/^6��E�@�hX;�w�\�/B����L��p�"#��,�D1��9k���� ��F�Ah�r�Z�6�]V�G�Yk����\���߃Q8�������nͨ\���CI��K�9A���C����MEd�������ӱ��'�ၭ��s��]P�<���/|�_;3�ܼ��~U�)פ#Y�¥z�0���۵I �+j��qQ7$��K��IYɥu�#ηf�A���{n�Æf�^?�|��*?��p���X��	DZn�[��}�T��q7K���)Nu���� ��'|��Ŏ����b��r�i!���D���mY:���k���y�p��Y��R�it�pC�rfv��
W���~$/�:�a�e��F˫���M7A�n�{�<����!��"v����0FGF��\��h��^�S5>��H���=n��v���m��w�H�M� %DS�칸 ���9��po�azm���g���C��oj�֒l����7JVW���h;u����Ꙕw^v~YX���3�é�gYE�O�iw\�ɘ�ϥG]����w7a'Y&羗�Dj3Ag��6.<�(ʷ{�%���te���9(k[��s�"�כּW����ߵ;������g�V��,_�g� �_P�^'��nz���MU}h]er��4��z�3��n�q��X{\t�\��i�^M[�k6�����m��R2�!�E2�m΢��l싯�:Of�r�����lq��p�D�V��Q��@����x�U����T]M2 ����E����K>�aT�\�ۧxC\tH�.^!��m*��۩2Y+��y�p��>��Ϻ95���uw�Nɧ�_�(����aS���	tK��q��A��{����I�'��<t�Ċ�y9g��3����;M�ﱶ��B�M��m1^�@A`_�F
���?~���Ws3J�O�����Fo�9b�����\ys{|�Ǜ5�VX�b��`�o<��q��w��DV�&��34���q۩�#�3x;�{�OT��<!s�]����򺝗*tq���
q˛���*�݅�%^���\k}�>4�gt��S�
�`υz���yW��6��q�Z���MYMj��؂~�e^��vHx�4��w~��l��d��yk��v�Y�by�Kf��w:����۪���۳���mnyz�t�^nR�m�Im���R����z<m��N���W��ٕ��^�=�NĒ�Ʊub5:̮qm��Y)x�ܜ���Bq:+��7Syr�swW�:y��{�����<��pw]����k���0�ܹqmgp�7v;�p>�ast���&����X��x�T�פz@Q3ۃ�gg����g��g��������o�X�ՉfwW��8s6���rߍr��9���9�>����J��w�<x��(N� �μC<�A:����(����T)^r�����k��Z�X�!0�hoI�p�nxNӵ��bV,h3{��"�z�e*�m<$��<����x�8�ﵽ������՞���)ӄ���}�\Av�NFd�4�
�.m5,k�r��k�}K��w����)�R Ԅˠ"垺��v���[�����j$�B�q�w�����e�[TD��B�[u�3�ݐ�,TdoO��;ȉq�ۻ�$/��o��5w��vV>S��b����S4��tt�*�����Lڻ翼9����zb�Q�=X�4�e�=��s�׏�Ix�r�f��.�fvv(��jək�}ɷ�ج��1�'U�)��>�qm�Ľڸ�~�B�ۻ��u�~�������+~�T��#c[�ե�#�R�ꗭ���P�"�%42��x ,�G�\�Y�/*L����H�^�-(h�\�t�X(�z���z�uޡ�v%��ޢ9�,ɏR��&=۝�O�3�Yz�?Az0�-��|;��)�BR�ZQ��C�Wb�þǕ		�*���Np��nh������N�ֶ
���xyr|J�-훷^y���4(�[b*�$���뻚Q�x��t�^���=��m��d��	XOOu_��t[}Grw&��s۩��ssظ�|"?�d(XI�s뼼�j]d5�wՊ�+�S]�o���v�_g��.�	�J�k4=	�ƦTMn��Z�$�ZV;���F������ꝝ�K��:���Y6�u۶g����al��.�*�����o�{�%N��[\�g9}'�$W�E\�	�qf�I�]�%z�%��j;V�raT �CT�$�4Ale�KDm؛�����g�2ΚEr�k#��?'}��`��{�������򔏲;�I�]v6��Mzߞ�]���L+�>i����<q���\�']��@&lq��wf�M���(�g�G���D�6�y��a�3gs�;�f���
i�dE��V��o)J�s�Cf��ݫ^Z���_��x�oK��E	�Yi֮��٭kZ�a(��"��)<t[�7ҷ�<r�^�|���o�>��������{[�r��ߎ�#8
�^�tL���]�VkV�9
�?*i�S( SX?{_~�����>�����|fR��0�+��!�#X��쥒���q]��Javg37~%��W_��>9g�����yz�;�����{nk�t���k��շ&Oܧ6aǝ�J�μ�����[�7K*���z�,2�d��g��{T7�%�L��I��!���g<�Y��p�C~rq�!XE{\�f��Cʸ�ī����F�L���d�7ry���y���T�唋�r�z�
]=��������o���G�l�B�����j�#�ŻV�?_��V�h�M���k��WX��g�kw���knӆH=��d��=�Z����iH����v�8O-h�A,;�W�n�� ��|��b4j]��֯{��F�y&k����ԛVQ��H�v�,e��� �z*M⛷^��f�Mx�X>��N�s�
Uo�*bj<���:�u���ʐ-�vz�Μ�y9<��Cge̺sI��U:������g=��Ŧ	)�| ' y��m/W{��.q�R� w��[�j�����WՀ��l��?56�>����������r<!�WI��k�Gx��&�ݣok�VFݶ�)���>؞��fz!�JH�(�VB*m����2Q�y���̍��y�j^{�5�ʡ�Z�߽�Tp+�W�cΜ �޷�f�������*�q2��r���I�G���|�+������g����/`~¢��~�)�"��=�W��.LY_��ګܘ�ѝS�:���3u��0��ݛ�x���� Z��A{��'����_}�W�z�?��c�Ї<����P�]��v�;'"
~iJ�8��}�{�ehmR��k���v�i�tD��/B�=�ѻ���gW"������r"(��>���2魇��4�T�Ӕ�ԉ�}~2��T��|گ1�s���>ki��0��v��p>����=K���Եz�+��P��J�*M�D"9u˭�&����]@r��^���u���j��:"�ÓVD�ū
�ܻ�.�v�c�d��;t�v^Q�8mtP��G�%�8Q�5��v��d�Ev��
n�Ǘ�+�6�Xv��lJ�f�fӽ;��y�{sC��Ȓ�U����67jL��S)�Y��0C�!�5|8�m,�R��̠4��v�AnMj���o�R�Hc�a��Uv���P'�^Qu�:�\6q��mS.��)�6�z`��q�cg���	�D�H��Vd�}��Cmu���v�F7{OY�h=�әA�Ι"ܲ���l�VL���^V�k�kS#���!�6�q����wB@���KXi>�_VG�kp�XB�����Y1���i��Gm#ȋ��m+��<اA��tᮗo��a��ǧf9�n��D�x�Rm)���z�+k���Y���+<�57z�f宬�x�C-rE,n��\)�Dᩊɣ��"�K4�̰�[�е�AV�^��]2v��wy�֦� �vO���پ)���YQ�F������O�[yw(ơHo�CNV_V�n^�}�d��nl��@rJ��֢�3t����h�b�!���](��]y��cj�f��2����;��}��ʥ�ҭWu�����wJ��ux;t�03\�j�!6������/E�jA��,��y6�Hm�^����9֒��x_Yە�VL��/��V��~�x��M��B��c����r��N��1&���x������h��۝�bus�v���[�i��A�-ֱ@`��]�my*;D�m�*!�=�qb�d#"�ʌu�h|#'��wq۶1�s�.�m��	3�ɺ�x��b��X+�����ݴ���[�;�����q�g1l	�Ϭn�
m�n$ܶ�.ֺr,��Ol�n�|JC9��֭�#�N�4����X��.�.��7:#�v7:6y�×��9+z�vɐ����!��r6�������;Htm�F�g<q[�>]���<
�m�
�yR:��8c�e����O���-p����wWmy� ���۔�fǧx��۱��b&a8�m�����㭰��ۮn+��7�=�p�.M��y�q��gV�-J�N �eݗ�`�m�_[�t�>;V!,m�k�0����wV��m�nb�M��u�KS�vWvz,v4��ӓTix��{\��n���g�
V�Ϯ���n����k>/
+�N[������n��m�sshl;H67N�э��I��u�s�f�z#�ȋ��ێV��m�n��[8wjIWH{n�G���9��F�b�5�cu�.�8�l=�Llk���	��+�]�V.��p�bx�H�=��\�Ra�wCu�by�_<c�YS��p�w>xr��s��:U;eܽVd��;y4���ot::�]���9�g���Qbi��nT�bA�T�z<v����S͝��:�p�/!]D[k�z2x�s�;��%�m�hqn���Ϩv�ں���OQ�묺y��:�D�\g����3�-YÓ���ti;;"':���;]��-u;��Lv�y�fSn=��"1u��ơVN:�!:Պ��2�,�K,Q��M�s�>F����onNm%�GR�ݗ��"^����h�byah�	#�@v[B�J3��$�O7n��vv4�3�ƃ�[>�M��%9ݕ�d�vN�Z�[r��;����΋����m�e�Wg����ھ�U`��X5���&�cv�\��ɍː�A�/O��G@�6����ݎ�����a�ǢX7^�������E�<v�OkAM���<��ry�v�]�v-W9w\�Y2e�ۉg�N7U�ϝ[>*N�������G�SOO+�s1��ϩ|C�[0p��,k��{���n	��p��ۮ{$2c��Cc���Ggc�;iα����v���������'�Τ�zj,�b�<TW��4#������r���-u�s�h��t��?1Z="�븯���.c����E�
Gg��QQ�];�0D)Q]l ��/'�˯���o�^�l�t����y�����cy)f^_�Gon�	R"�\2�-��3��t��ÀxÈ��a�
t�lvfM��B��ڝ5fM�
��Z�Mc���2�o��������WNH��3}+��m�M���I����������+U���<�.��*�5��^M�&o���`�X��n�Z6�(`~�)!��·pe�un���q����h)5��z��|�ys�Im�p�ǩ�vg �Y���w���|Z�����y��a���=j]�̷�my,�	LMY%���R9Gb�H��	n���t[a��]�c��?���a1+@���4C/���L�:v�b�?zG���*�۲�c�Ι��	L��}6�N>;w̺�+Gۣ�� k�~�FW��!�&.+�ߦrD���ƣ�:����k��_�v���u
)L᷽R�e�f]�/v��#D�,��nJ'���]�y
�@�=��Ѹ��c���s��8�se� I�w��k(��y^�5�jF�{z�f�Ԁ߉M�$4o8��{7���xo��d-� ��{<37�q>��4&F�MY�~��/�zYW��_è�)�~��_�5�*y/y���/o.�<�1I�fs>�1�&C�kڷ|ֱ�'~����W�B| ��yɲ��[e4�t� M����j�e����Ã��ZV{�Yܭ\����2�#����-��km��ĤLV���\0᳭���LN�nA;X���i�e!�C����<����d+\��n���&���N��Eؘi7T�ctJGWm�w�ZZ����;/��&�����>^���ۭ�Ǽ'y��22ɇ2��ϗ�G�H"]0.����;@��j#�}��T.#,�_�nt�B:׶s�[�C�M��'X�˽![ޣ	n0dr��s!)�5��|��$��#�Xs~^�7��`�l�]�}��갓��.�\�hw�h��y�+�'�G�F�P
�
r�Q�g>��o��.��;#��n�4��s���h��bb|CsR��^-V�i��=u�w|�LO���'N����޾��~ԅ0'̳�-������_�x��QI�����,f�-)�~|�#��)@�+��������!����{:g�����m`Ґr���nӁ|���z�3��V��%2{�@m؏����!�g��V�u.\��� �2]�u��*��׵��߽��s��;h�zmZ���l�ʚ���rC&��w]b:9�g��v���[[��ݒr�&�{���OŌ'�5�j	+�xJ>�m6�xS����H����w��pHT���Be麛�g���]�B�뱀lr֯-P���jK^�="ŋN�>~wc���A�Q��y�Y,�:�^2��+é�<t�tEQS�����8�0�u�u}�kޮ5��mZ����Z}��o'�OTGa�<'����w3ܬ)��=j"�l�Z��0�Tz��~yG������f��d �����˺,��y�`0���ɗ��ks:���ƺ+�y�J�1��E�b�/U�b=B���[�]bw!Ͳt��'EEt+]������1�Q_V�/b����:	`HVy�ZZ�E�)eeqߜ(^�Ż�y�c<o�iZ�J�9��Q�C��������w�p�tM��/%�a~������᣺
�~�u!0A橠An�Ů0ϲ��ttf;=�x��95�"���Wsp$g�)t�h�S����q�wk�s�|0�)��Hg�3� �Ce�V�H�
��>���'�׹��� I�U*#D����C_�� �%��f�IB.��Wj����u�xu�����Xe�!��	�u���_�h�쩴7��Tn_�v�P�=�wR�W�{k�n�,���%��^/�e�����C��E{�;D�̨ɸ�����&�z�dT4����&C!6q�gt�v���|��zۊ��1ܛ���>�U��7�݊��w�Ko��(�����*�r$���!��-���Y�X�L<Q�l�njI7�ǃ��Y�4
���C;���Dr��o�c��.�R��сNX�����(�JgxT��R�WLX�U��T",JW�3�yyf%N�Dy�|×���a`,Y*���q>$�̥����WV���);f�����r�jչ��1��g�	���msv
�9Ŏ0���;)�Yў�v���r�6�^r�nN3���f9�l�Db%������7�h�Yݨ�7GI�a��5�����-D]v����pv�z9M�����|#��]�Y錉�nI�q)z����r�n:�۹8�U�i���v�y��y������mI���d������źM�]�qq�ۦ�$�������0S��n���FȆ����-�/^9�ѓ�~�`O6��!�ͺP&�){c/��K�Y��-4X�}��IzM��]j֧���m�N�B43=�U7�Y��YM��s�iI�O�g�����bE�/L8�Fۋ���Ovsլ?v���qϼ�w7�V�7(lg�t{o���Sr�	����Kͽgy�5E�m��k�n�r��Jf, ��>�~ �B�ЏU�����UΓg.��ۿf���ۼ����p��b`�}v�}{ʲw<�^5h�>���(!3јS3�P=�܎��ż��҉��g��vn��
4���cv����7Y����?�E�����sDP��z�TϮۻ�r����}|��3�Y>�{cAI%.o}:��u2׍i���<H�Яz�?���m7�8V�r6���Z����s/,��)��)��b�-P����/`�P��{^��Q��ӟo)k�
�{���3�]&��k��Cw��*S�N>涓WL2��M2�m��sˑ�G���S�F�ĳ@�H&0<���ؽ��p*��u��+\ܫ�c���|��	�E�Oj-�ca��)�s*�WW�U3�D�R�-�1���_�Vjyޑ}�އ_X���P��?wF�v�ZIs�\3g��
�\񪲕;���n',�]�%�k�{�vvL�T���d^2ڭ/����k�w=����X=sP����K)d
j�調��D�V����ʭrM��m�y�<��j?9��ʁ$:���O�U���~��[{v|��k\�NB�����g3�`=���w��ŽZ�l��P�����+���0�Ї4� ���"P�h{�^_��3�����z�<�'��;�/2g'W^ߕW��Ϝi�Vܵ�H����쓞�pݸ�	��6ts��V��ë$	��s�pAr����;��y�Ř��yJ23NP=��K�ei�	�M�^sEb�G��>��j���V���̴-�A��YmQ�����|E�B�;��h��>|m��J3_����o.`8.��9d�����%]d�MY�K6�O|�R�p�eDP�Tw��y{��b*�X��R�z�r�7�#�m�+��wi���Q�wrM�F��"6�r��ʍ(��e��y�rzj�PU�� �7�LāǢ�-&�m���GFqlD�Yx.,~���=(g���GZ|���{�w�0!l���p�6��^[2�c��+�����9������<�{kmX>��u,V=tk��_u<؜Uu8��w��v���8�=SNy�Gj>�1S8�frK,$<��˛�F��CY�rO{�|s��`������"��}�n}�b��ϴm՞=��֋h�[p����nýB�A�>�#.ќb���e�\	ۋ�;k�7[�� ��:��}�浐�">f�^T�+��,�?q�{ܭR�Z�Q_��B������^�՞�ÛDQ��0ID�����M�0޷"��t.��2b
e�w�o:�qګC�����xR�'b\��[�6!��z{��=�ı~�g�I�^��xw�03M����&�=���ko�V�?	a���}�vr�g��bv�;�b`����y���5.Xp��TM��aJ�m5����#�G��s�jŜ1Z� ��L	~���>`fH�?t����;Γʻ� 7��������Ѝe��2Eh��ҕw�;G�9o���IOO<X-�n���z���v�ɇ��������CaZe���~"�>P�����Ѷx���Dw����V����Y���S�I��S�-����޹j���bTz�j�	������
��V�X�m1�c���q��������v���N¿��Kk���\��h��~3�z��+�k���y&t���en�.���L�t󹡪{fuw���;|�{�����]���v{�O��׬�
т�-7�{l��]��j�����Zto��H{N����5�7��^��G�b��c3lK��ݕᯩ�N����+E7�!ʵ�IRlJ��\;���s���iS#"��w����<$�v��i��9ս�o+��`u���������q{4}���|�$P�SW��I���֪�k��㻱�ܢ�V7���c ��㛓����G:����_Wzr�<��G���3@�g��,6>!���5�.L�j͔Qy��\|v����Ogg�e��������D�z�K�y{�OhʟUD�W�8��E�sɨl�w�6<+:�e�VW�̴u�y[�����K�i�=f���]��0X�k����[��$�k�	P�F ���\����:�F�y(��=�e���<��xáݝpVuf�6�뮠��c��\��q���{��U��n���lk��8�N�k�<�mnΞM�q�=u��'b���yIyƄ���by����mcnն��w#W�����a�[W]am�p뎍�Zw(�n�]��\���7a����F��6xq�I��NXw[�������]�Qy1s\�
<�8D�9�'�c�:�]	[�ۖ��`	�,�[�����GK���e�QU��b�V_+�2�Iv�u���4��^�m	8��8�ٞ7p�s��I��k���d�m6���|U�l�%v��W�kr���}�ﹹF!�Yw�6�L�rB[>h�|�OHs�V�g�����b�U�>�/`|�Yܖ��l�[=���н){��u���ٺ������ʏ�������l��O��g�{;��_�z5��U�ȕ_���z��}��b�2�pV�����&��Z{���i�U�yq�#��Ur�T�;j����ݚ����XW[@��X�%q���f�\��j��j�̰1���&oh�]�9)95��B�6���/]�l��Gs�.�%^$�:U�K���a�:�$���e;K�э�:���q��ݛ�{s�64�pv���՞�i:)����~� <��	�"�h�W����9ǳ��؞*{�$w���%^Z�k9�CΦE>�ej���*�@Q%��g�i�A�\�p:�{�P��w�ٷ*���z��� 35f�vL��Gj���
�(��u5a�w�AWE/H�{5L�d�o���O7�|�T�y����Ӽ(�[��)��G.z��'�_�7��(���~#~�D����3D���n_�vQ�'�NZ�xt{���E�Y;��U���T�v�'Ƽ�U�v��@�G-�vP���R����'y�V���t~ڲ�Q�4�S�xD�w�HY��,��}�JT�����'��>f�|g�W��M��v�	�J!6R���y'EpoQ\�ֱ�H�Ӽ�#Q�n�\���l�qUɧ���sOO@0w���$��ݬ�]Aud�2~T)��2H]i;�cpu�5-�qp�ݦ���p���^\9��P$����['q�#�]�_��@����s�Y:�Y�>�Ӌ��ó:��5k>�������m���Z�W��R(��5oáw�Lj��~�꛽W��\������ֲy֋��@��w�{a#�-x��R�����=#G7���EzUܦ������fV�X�a��6�0�n�t�1���>Of�r���fW���Y�{�핾뀘�=��*ܛ����J�~/h��%�9�f	KK«�W` X̹݇z��sLy��܉����7r��u��8�׶8*���!��],�����f��{�0Ь�_}���]8N�#Ds��R�r�Z$A^���HT�v�Q/5*��ž���Rw�'����uI���b�n�+�XM�z���	�.�Q�q.��jU�K&H�]��]��<�����Zck1	��0�%Z�v�QGz�Z���ܱ��뾖�-��tީ��n�'w`t�%a��Ɛ�y��lcED�8��z����#foZ��YΙ��>��P�jV��i[��G*����J[�����;=�
�������{�.M���Y�Y�v9�u��x�V��%��.�<�g3�1�>�O9=1���m�Sz�V�G�K�h�w7��2�sW\
��֧wCL� B�dιg�^uG�l��G�&�DCEZ����
���F�Vu��J�6�e�����HY�{&.�I��뽨I}��2�F�d��(h����o�uf�kV7fs�|����6�M�X�T�9����S[U�m��T���-)�zT��Nc�[��)�W9��_l[�(]�Wt��J��)o>G�����HmQS��
�ۛf��{ٔ
(��H��sm5�+8�.�%��mBr�ej�g�,���`'��+�ף�f��[��&m��6����t��\�KNdeM��������Ȭ��X��Y��<M`���,��Ý��s��� ��ҳ���� �������{i���;��c[�B�l�T!P��==#м$g���r���_���`e��`��3y�b��c��{�|��x4�ߺ��Y*�^��!r�e>����>�Qv��mS����W^X�qjP*N����yoE��;[�z���o�{ёx���;�h�_5I�cr�~ꉉG����L˶� }�1ڡ3�6�Od���c��ZX���{��f�[��4��͍��j���i��������j���^=ή�4fՌ
�q^b�-u�O/黻͘��$���Vx_��R�v��@�W��8ׁj���yw��#u��]�[+λ�V<�]ۭ&�-H�� ��@�mw��gg"�0��^��@�/x�%GBJ�%gΖ���8k��eZ�Y��Ǳh�Ѩ*�i�r�:9W�_>?y&W��lH�	O�6�4�J���p���3�v��m9xƍ柙�Gc���TqHh�������?R��&��Ӽ������A�9rPX1����oڻ<�=�%��ʼY�W����Lfs�>�f�ݵ��T�
��4��NT��ꊻ�K��u;�8܆��J��zn��
�����.�S3%��*���d����[�P.�5:_��*���~��hYt��jay.Ϝ�]��m�U{��w�|==^�R5�����Ͻ�v,�]���n�тt�K��&ի^�l������G"/u����=Nu�.���Jj+���]-fD��3>)8��yq����+�T�Q�t��<�;o|�An�bн��}N�Es��['��Ub�S	�q�t<�ܿ�����`�f����F��s_7*���|}IO<�����y�ב��!��3M�����^(�.��$�]o��P�B��������
m��M_��*����@�yK�ά]qY�㼆}�D)� �s-z��U盂�x45|��C���5k�Z�F��{:9�y��I��HPn�m��F;��.�� � ��6�e�\���^��v^��C��s��=�{�������Dy�|��k.KuxN��$�M�_$�^u)�����ؽ�{��Ku�y�*��|���q�A��y�_���6���)X3�P�~��8�T}6w5P
B��ʴ����f����0u�Wb ��rwJ�n�p�% ��b���9�b��`��6ԫF���2_�EWh.�Ab�z���V�n�u�7��ie�\��^vp�R���'U&v��[��Քg���G��/���a��^Rz7j��R�HMM[c���Q��۶�]`��+��9콶B�D�Qv�Zy�^���9WV�>��n|%���X�m꺴�q6��`�����H�U�p�\ȳ�����'@��4�ֺ���6֡��F�N�j9������QǶuh��]p���0d6���Z�ݰa{E���u�hY�g�r��l���+�r%bŃe������^~�r���ynR��0�#���^�E���)]�K(,�o��
�8�����ۼ��N��U��`�F�97�����s�;���y1`�*��Ǌ}d��I�k9|4�����_/m�6��X�	���\[��+	�G���XHVՀio�Ly9���r��w�W83�#מ���mF�U��.�Q�+���/��h��Gϫh��4��뤃��R�6ج�:�����d���.��uy]y��c�=aSDy�=�W͊"�>�p�a���V��Z��Vq�寮�Os>�qU!�{�<^>"+��A�o�����|����p�m�x#/��u̍�h{�=���**��t�b�,S�j�!�nU�\O�T��K{�F���#�Y�T��\�{Q�ր��#���ν�޻m���u�/l��h�h:5\Q�8��O��R2�Yޏ������b�褳����w}���s��8��{	���LzE^�:Çq_)ludh��DP�\��]���W.�bRs�	]��q;��8r�4������]��>�z@v1��8̣��eu�K�W�XͮA%/V��E�ӦH�۩ۢ����:���� ��L��j�1��Y�-�GjD� :e�D���A`�����/u؇-$���V�wMgq��ߛ�i\�\F�F�k�Ě���ؠ7*#�����@��nW�k-,��e�w�A�:&�i�@M�� �6���T"���ң�w~E���,*L�텊�Ωɑ��+�: ����=(VrΫ���X�a��t�)���w�9�"�A��P��K�����f�HkT�>���o��� ^ι�P�Wء�͊���v9�)p��Al�������W�����smFꎞ�y��a�t�ۯ�`�y�����2�%V�u�"l����I�z��1�_��9���Oi�㪇�bs����!<��p`��ߦgIR�-��Q�:��m-�|-#W��2-6�z�xJ��J1:��S�9u]�\�+W�U�c�O*dT;7�c�v���dߣC������w<��fb������}[��[����rҠ��4KT������
�'�=�ñp�}y�|��V�F�׌�e���x��Px?X�d�Dz���x�E���L�5z2��Ztf���ez��j
��y������&2�׏Y�F��z��e� �ɻ�p0��N�."��.�s�s��z0�3O_�˔�v�3T�7�z�y�|��,<ЎU�cz��o����92�%��-�-w�e�D����He�Qo���Չ��B{���ge���f�6����\(�ʰ`����@`J�c~71���x㚕��zɽxx�gkp��ƺE��=m����vzF�U��VU*gօj@�����x'�/o��b����a������}��^�K����:��ks������Vv�v!}Z� ��,��� q�i�n.�f�&!�����Y���sf�}��s~4z�*% ��[���W8#����&R�{�QqH]���m�h���GT,����.���gy팯&��
o��!w/=8.YB�׻�Z���M��}y5�9��[{�Mg�'�Q{�[Z�r~o Mm�L��Qי��6�����]�W��E\F���i�絬�����@y0����7i�T�Q�}�y[:g�S��E*(̽�{��VS���	��m�sj�.��n��h͡t�5��$�Q������{Zލe�Й��� �IP� ��%j�q'.+�u.yaN�L=��;��k�w�Y���wbQ��n��Q�����í�C��{k�/~�Z�U$
��ei��~���Ɓd�/g7;W7����:ǵ�����{9�۫gt�c@gL��������f6ފ,R��&���zI�#�P&���E}/{�����H�M��8���f>�d�I2��a��Ϲ�)��;Uț�$������ff����w�oG��S�$m��/���ǅu�a�H)$�;({u�Ub{�t�z��"��zv�Mޓ��v�RK³ٳ=2??!ǳ|��-�v�[b�����e���Z�Gh�m	H�=�&Ӱq�Fd��p*w�q���s��ru�lKۘ�oxy�!��e/e
O��{۠��}n�K�{�6�I���M�IQ�{6rW������㡫�r�#O���2tV��-�hے��}��q��vS��L�uu��e'�-\u4c;�b�!Y7+r���l�ɓ{�W6PۦS�JxH�s�����%݊T:�s�t��&Y��f�йX+{��B:繻��d{:��l��k\�y�W'\	�G��O�y-�u9��j��i:L3�y���Y�G�>"7m�`Nݛ����]>ȩGSr�v�Z'��v��`{k�����ɸw�w6���m�ڍG`랆����݌\x���k��Sp�{�c�`(O2;��]�����8��qǮq�.;rq�qX���una2����s��6��F���6�7q� �����;��;p�A���8ލ@p�M�3�i���~�B)�g�p`��g\�0g��g��G)�[���y���p�f��C�rn���)S�"6?f�Z�Jvq�d-b��VإqZͱ�C�qm[�b�Yy=���$�x�=�P�R��-ew(�N��%a	P(4�e�ڵ�(W�X�M��b�B)VN>oͤz�GY�6b�3'd���zq�M��X���Z�셕IBM�JM��T7Q���f�ѯ/ڗ�D�(�v51s�{�����+�Q6�/�f�dW�7^p0{��y˦׷U�+ݵ+��
D��%�۾�� ��癞�R��������k�F�/���;L׆�M�b(���p��VV�a��H �TWm�]�ׇ��2ͮێ�& ]�;�M���ۑ.^�WI+���MKA>������׼lzC�;�R�Q�񣍩��	����l8��d�}n�=h��7/�m�����dPa6�v�z��f>ǚ����^�حaU�Ԍ����%n}v��WB��:6�os���g^�������ȅK���qI���JD�V�[N����`�o�Z��<�_\���[ƥ�y��>Ǡ1`�¢�h�|Տd�﬎�����M&Zt���l��)��A�u���:^;�ם���G' ��/���F�ю���L���{d�5��fh�%��U%FQ)�H$���݆IOپ�u�I����#b��}�J��i�^4xy�{�e(ֈvxY���QRLj��i����ډ$m�гS�CU.�~H��?,��b/Wz���E����L��ʞ��,�w^�$���{�s0餽�
��;gu��N��U�Z����W���88��pxi�h*�al�"�B��_w4z6����a��Ư��%��&	uepU�����6�oL�9׶W|���	���u�i]�>�(CMBm��i�s����y�-�f�2�jex��b�y;��3�h�=揝�S�i�'&�(�x�k_T�"$���s�����w��f�-�^�o���ۣ�ذ���V��:�M���d6��GΧ}�YΦ��}�!��v�)���H����+4�p�wջ/�^����,5���\P�I����G���^���I'̔���X�r�F��a�)0s��܏>vG�G������(�["�>~V��!<Pb���Ҏs��m���UqP���(����͗y�&���hVoX�#�2���h@�S��8��:?vo�Q͞j�������[}\z���}�����p�(���n�ݖ����n�GQ/&w<��v����e� ��m�7U5i����k���w��YSȗ�G1S�ɰ�D��Мun����Nbq��z۠��T���v G(�ӳ�!����G�ʷ;9�q!Z#���Կ>�QTU���p�����FWY����<:���P�C���U"@2������WȖ�%R߄F�a��h��=1.�jiGb�f[��j����j�ͽo�ܰ�@?�	�� ip�V܃s'm�Pnvŧ���f��HE�jӣw�7��Z�����+V��NY��^\5H,P�;�q��bɖ�I�$�0�������Z��,\y�:����Z��ΓV�K���L��QQ��ҵ�B�^� r����H*�K`� �n`���asש[��P��d�8����z�'�u�a7A��	��%��E]M&�ؖ�`��~Wc{^8{E��M�����̢t&�v�*�6�{qs�9L�w�A��t�Y�����f���9m��,a'�w
B��=�ٴ�[c\07767��R)2�V��� ����w��su�y�KbvީcG`Xx������kk5FCQtK=4��vh��w��l��؋o�Ti4ټ�@-��1DW�����o	ߞbB+�bZ�V�F�k�oL�ՊO0����B�d�+��m�����xV�[�;[��(;G(�v"�e�µ��Fi����oEmK��+�Z+�A_wL+mVe�2�t��Фv��ٹelL�M�*����U�oeKZM��Cf�P��լ#SL�������������`����HJ �@�P	$	'��I I?�II� I I?�$�$������II��$�$� �@�P������ I I?�	$	'� �@�x��� �@� HN@$�$��b��L��1My� � ���{ϻ ����f>� �  > w+�U]��;�;��φ:�@\8�@
(ڇ���>�^m&Z�0�]�.��A[iU�)0rs�f�7gT;Vm)`��I�t� 
�:��   �{iJT�      *~�	R���  � "���R!Tz@ h     jy�I�S� ��@i�  Jz������&�C&�� )I��<�z&&I?Jm�z��&�)�jN����몐Vl�'�H���; ���������VVCk�2,�1fX���X~�e*+LQ�1���]�Lϳ�W�ۮ;K5���
����c�;��͋y��O���#8����ҪO���'���0[���XI��Oa�$�,<�V�U�W���*Q�Ǝ=}AR��uu�t;v�0��OF+�����n��ͺ;����%^��L��Qˬ��0.�,oNd��͕�bZ�.��4�8IG9�6�	M��F�t⎟u�ӶH��h�.�,ExE�óGJ�Xh7����N�Yk.�Y�.�n���/��;	�����F���b�:--5x)���6u"�j_�OmuE�ن���m@��u;C�qJQH�yٗ���Gs{�R�%1�9�>��ge"���L'�$XLkt� R�W%� ��v4��y�T���G+��ozt�@:_m[B�U8��fq�e���S��uM�`  2��3>�0ٳbc��.�~��N�r>�>,��:�=��y6n6�f�                                                  m��                �A�                                                          7E&b����"n���C����$��B0�hS6��]��.θ!q�l4����
YM0 �Vq�v9����*�h#���LYUme������v�m�w4nˊ�&ҐQ%��h iKqay]Ԏ��ndٶ�&�`ݩDmNl��K��Kv��m
�-릒���[v\BtJAܲ�V����]�0;U���n�jZ���[�@�Z5�\cdf�/RSV#��R	�b��j�ierT6e��;i�Z7i�Z�)p�Me,��ǯk�٦���I
�N6ؠ����|�w����c�N�*`�Y��f?�����A�)��n������       �  �@          �[�rU�f�q��V�Jĺ�i]i;Z3:�Ѧ8j%-�]�RL2�!�f���������:�=  � [���Z�����D	C����>:��8~�����O��I��8��>N	����+É%(JFB{$����}r6(����ط�!3}���e`8�RF�@�b\G:24F�=����C�v��A�4�1!%a��N��Ԙ�pM��p)G���2��Wxw��ޭǚ�Ŕݺiwl��2�����I$�I$�H i>m�N[�6-��cd)$e�w{���,ie&�]�B\�'tL� ά���H"I<�Uz/j�>�!���j��x��бK�]fѴ� % !��g*�Q; 2��eξ۹�իaU}]u�đ����d��;|�'�L�C7yۋʑ[�mA֯�FV�`��jC[�l4���	oS��VU�i��5�3َ����V'L��&��q�}7�w�w� �  �P�`ki�l��]��GNz`��(j�������J�n��s�����a���2�v���������eU�%
B�]�,%��]�8�ј)&���t�P��P�0q&�AS��B�2���=�ݕmYWaC/X9ۨ�g�/t�
r|'��|������SJh���7���5�7�n��%u�f����*��|�縳�y<�i�{�^��`�W�뻡�����B��i3�U�,rQ�nh����5�����>y�^���z�����V��G�׻'w՝Y=x|3��˴��+)<��nX-���b�;����n����O=���    ]�wQM����k%[wo����S0�E�)م�E�"�fu�l؋0�2��XE�E�"�"�E�m"��)s�\��1P�E$=��ˤ��=p��nfcIW1�2���w�]��M\a)�s������kٯw�����������Ŀ�7���{�ܔő���}ߕT����2��8�g�0��w#�{8�
p	��+��s��~uAlFd�S���g)��~]��sVUHe8ƕ�Ǳ6Wfݤ�NvC��T�VۭTJ,�d�����ھfg?O�|���A����5�g�˻�����G,S�wڀô�j��`Sn�H���r骘�a�׬ߓ�w��    Iub����K�Q�T�R�M|�<���>5�]�R��Wh1�%fm�Z��xs���U3��l�N�u�8�E�c}�swwM�Yx��4!l�B��핻�Ĕ�M{�Da��넞�'���l�τ�<�|�U$��D_#&���G*W��j�-�x�OOiow>|���+ҡnݤ�m���kwm�L��ci�=��Zc����EX�e��q*GT߉-s6�p��}�Wn���%��*�F�i�i�\��z������cl��<��P���@�����u�|��ƭ�wX�IG�8���ꏛ�+��/c*q��t@��                        f٤e�U�T��I�e�[u����+u�-��������p�d2�J�[/6�M���/\�    6��I�0\T�c"���y3䒯��L��C\����bs{��F`�����H�H�	H3��U3Fn���(m���H�Hu4��% D�H�ԑLKu$
u�L��F T�\��13)���Ӎ�&b(i"X0�)$J�)�)�,�űi�"@�bX�`)��HL�
@��Yd
RX	H��I�)�)$�IL���wu3UeUYH�H�H�BRC	�i�b RX��;� R Rs R@��,A�� X�b%�`�� F2�J@�fJH�
�vxɔ�H�b%�`��� R1�
�f&bf&bf&bf8�.��y�-LDFR PR��H;^��ݕmYV`�H�H���)�e��H�H��V�o��L��Z�̦��f&bf)���A�j�H R X�c#,H�b"P�
�(�H R R R X����K2�5li1����vԷkZ#;삜Ip�؊B�sPK�_d��q%*��U�T�s=�'3���y��   �,͑5��h�	EUvD�=��m�I��{����2����v�92Ja�;�D[�i�o&�ww��ʥQú�-��]rE��kY�^CNR^���9��Si�#�+�r�ڐ���i�{wmSVT�u�gS���V��0�{4�x�g:��}�}��9z��a�x���jL:��#SI$���L���j=���*<���"��I��%���-՛ޱl�Y��w���N�8�}wwV���<�I�q�gd�.�nN+��}�!B��Xg{����	�6w�ʅ��g���I$�I  Kv_&���Q-�*�l�=���kM�y�ά����%<�L0N��� ���0�	�Է�Ϟ�V�k<�'}�۬�}�&��w}�Ӯ�<�s;c��͆Rܢ��	�]@�C)[�cwwW5VT�Lbu*,�Ж"w��6�x�{�wiwOV���r*NݳB��kW@͜�w���Y+�&J�=}ߔ,b�ug~b��g4��EP)���؝��C�����\b�+.�I$ "P��E��Ŀ+�����Oi���t�V�E^�    	p��e�k$������y�=�<���4=��P���2�7^9�-$����ͷ{��.�z��dt�A�e��u`��-$L�*w=}��5K/krq���e��py�4�R�D��i���37˚�����*���6�[�"�-Y,o���C$̝teo�:�_~�������9뾻��r�   ��wcR��v�F�@7W�e�(�#q�+T�W��q��f�<�R�%!u�6Ȭ����gp9��r�U����XT7�P��%�h�4�% �K;���%PƪG��`�o�M>���&�$`$���U;.�&���.�	�eY�R��>I!aR(K�����2V�S�a�{}y�ڵ��A/��E��ȩXzN�i�X�p�kt^j'����O@�6Wb�(M�	�$�I$�                       RVͻ���#���m(m�hUc��m�\��	�Ԓ�A�T��6k������i}���y�~;U@   ,���W3����U+}>��}�b��2Ō�P�p67�Wt%�ԒD��A;��Vd��C��
9j�#��Ô�O��I	ID����Ln�
��@��{Bd�m���kK�$�D�MC�𙲜8��l9��aKõuď��{��u��JJA^���U㥕�n���$:(;�_��-$�I$�I  �eL�&m���nݤ��(�Q7�'���8�x�&;ss2m[�Ӝ��o,II%$��YEw��5״n�6��ؽ�ew^vV) :Y&N��I2�]�αö�l�9�܁n]x�31*�}�+jc�\���)&Z�/C��מ��=|
�}&����_�~I+	Z�V�c�@�x�Tg�̕g�'6o��*{�U%وD�#I$�@  �][�6�Eɩ�HI$e����6���Rr64�u�t�{f�.���+%��?$�($E�����cq+6�6^P��e�3�R��^&�9䒤-%a;����EҼ�'���׻)e�on<2�&E��b#i�-����EZ7PSnJm������������6�:�3^��)$Hu����m��.�����Lw{%tɗr�y$D���y1a��\s�r�l'�]e��Wh��S�եZ,^ԒI   m��&����d��I"��.0�e��.����yǗ�9p�%ڨw��6�T�v(��"lNW�5��p'u�y@*�}�$��s�)WM���%�x	pLW�	�h��,hἒEQJ�Sc<��O/r��eq��N�i�3Զ���ʯN��$j�VS����/�.1���UtE��V�*��!]o��F�H�I$�   �Y��"jn�"�D��FH �p�f���;�j��ݣf�̿��?O?��>IJ6P��;��+�]qq���E,f�B��J��D(E	�v4��B���k \:	7���ֱO)�"�*���.�gtb5��S��oJ1��A��v����ʎ����$`��K��1TV��m�D�0)���ؓ���e@nL���U;����օJ�����d�� 7z�;����<��9w7��o                         Q�]��1-&��&�бZKF�L�k�ir���Ҩ�v�Uk�m�,b��f�/8    ��ͺ�e�غؙT�R�
^���*��+�YO�Y���կ2�M[I�
�aFh�|oS{9
߁{��sg�ͩ�M�X@�K֒����Bɸ&\����p\����uB�V{{�$�	
�vG�����?{9osUMʴ��I���cΚ�2�@��r�4"�P��iGC�y���=��z�ߗ���}�P    &�b�[tʛE$��e<��n�-���W��qg��Ҝ.�a�=I)H�$���gu*ۑ9JL���g�ǲ��zT���V
�mϘ��{�0�Q�z6��'�n���V�����4�đ��^1��I7�YH2�]b�ڋ�[�!��@%E�d��an��u��ۻ78�r^giέם��{�   �p�fx�a�`���ǋow�Gf�;�k;3gb���>�Ƶi#% +��
��;
�r7�RB��k���p۪�K}��F�V��w��-�Rc��ʍ^H�F� ]%P���ŝk�u��D�_j��;�Jm�Y���"��z�Nٔ;ک�p�i)$�$�S��>��D�����B¡��.������ �B������tt�m�̬��ᘮ.�ȓoxw$�I$�   K�u�|1arB����DY.��e��}�e�~��@�1�F/���[��3�%h ������]�4o�^֍�e��+�X�]4Z��M�i_bH��h�Yg�a�g�v<�6��u$V���T��\p4���fu/	R���w���4|E���Xx���;x�I%!����+��l��K��&{��2��r2Sg�����    ە���Mn�+Jl,N���� %��Y�2�J�ӻ}=��ԑ�	]��:�Vr�+j�>��U� }ZU����\��$�JR����k�9a�|i]�eъ@��U�Rmr��q��*�V-��w��	?Z��!t&�|4v��G�Ӎ�b����H�%	���疬عe�Ҷj�%�)@战0�'�CjP�N�/7r���f|����zz�=n���\u��"I��                        ejK�u�nf�Q�K�+���4Ä�[��u�2q9���W��YE�+|B.2���!�    ��r�\�H�-�eI$�$jڇ�1L�*}�md���ܳ�{�� �$����'|�r���i;Y�/+ty��"U�Hw_3�ݏYY5ڪ�*q=�]�2�m9�V6��u�$��oC�ӡ\m�ƪ�Sp?J5>n(�r<�㋟$����fo{+5�l;Ŷ�S��������sf���@    ��1Q(��
�*�a�����L���%�ـ����o��.�후���2MB�=��B^�*g��5�r�~�a��ǯ~/l�$�%h�[��
�i���ŉQ���]�m���8�����=oj�Y��/qm隫r�,ɶB}p�ï�T��m��H�`��Q�� ���R�ͽM���   �|U�&m%OP3Uv��n{�Ͼ����7�ńxy�xz�X��ߵ$n�Uhn݁���B�һ�3'<׮Ḻ81��Y��7`���cC�S�����&���|b�����q�vi���wm㣷���
gt<�`ƒ�r�nf[��F�dwS��1ތ��RJ�6���UE�Y��\&�u�I�-0�!��ư�H�	Z�֭}�#�ؕ�/�u;n�$0Dj��KI$�@  ed�A�D�(�%RH�I�j��l��Rq=q�\��f��]�IM�.T/5͆dm�l���s�^�m<(|�|�4��j)�k��cT���r�GH�ry�vcԒIIX)��=p=ź�h��3.e�GG�/NB[�������t��,�35�����=o��ݗu��@   $�m�f���U-����Qwy.�1�d����2����RH�
�#�r���s%��^�˦�w#�x���i?i%`��q��Έii�yK�;Rms��IY
�����ãT\kU4�μǬ�o��Zgԑ � J;�Z�X�7LM֝\�`��[
�aEU� �W��+���a{�U���K�ܷd���_��{6���*h&�L�T}�)$�"��G���[�r����+�Yן�9u��u~��؛xv�\m���9ao��|�8ɷ[��l�w�������[�+������|Iy_�O:�8d:�
���K��w���_Խ��3��?G��^E���P��ͅ�����o5��xW��_4����}��_�m틎�t/g�ZrӲ��6.&e��/��垬�8��UR�*f� +E夜�j�E�gh]�m������{]w����j8������z>��/��.���C�����&����b�~Y�����/1�z1�L�/y����=��v|OC~e�h�K���'����OļK����/_��.��]/ϗ�f�����\����1�r�l^r�+��}�K�W���V��h]W�j�䬪v���ƩT?,�'��B٫��'NE"��ܱ-����np[��0���^�K�q WS���sK����W���?N�h}?ۙ�<�R�.��S��ֳ�]ߓ�K���]�+����mS��<�
�<w���r�u?�:�=�p���b̧��e��^��S��]\��T��M[�.9�&�
����s�Womf�_oQw)��/7��
���z\���e_��=���[w�_�wxu�+�1nkb��u�Yȵ<s���c1/(�l1���H�
��@