BZh91AY&SYE#��8߀`p����� ����b8��  m�����j��j���P룥)� �J ��@�T���:�SMV���� h���X lm�T�E%� �A@$�%%A"��RJ��ID�)UDI)JP���*�$�U%UD%$UP(�EUT	����}��ﳻ|@\��=�W�l�ײٽ�ﻼϛ�-o�׶�����%^�{�
�wt��h�{�}Q�ﻃ�������=n˯nP��'������m3(� 7���BP�$"�>{0׾��e�Y�uwZ��|�����Ͷ/}�����H���ݾ�ɦ�kj�=�xUU�w_}�>Ƶ��E{�^��I-��S�aϨ#w��.���A�M��@S͞����miu���:N�� iVZ��w٨O�>IS��ۧ�{޴}s��7<���9h2��ן2�4o]�ٻ���o�����P=��{��i�]�;nu��s�(Q�nn�X=6e�׳^��%5﷥"'�Qxz���u�Xr�J( ���P��R� T� ����U��L��z���}��ŋm�a�v��:�w��U�3��ǡ�۶<�uU5���z�ͭ]�Ӿ��y��[������Q^^���O��T���7����E_cG{ṣ�ֲם�e殧Z� ��v�/G�Q�|�I/�Q�7Uv������A�=��3�{�*��N�ӻh�޷�k{Z=�'���}�^�=aq�;�+Ż�S�we�5��
�]�p^>�@����}�y�5�� ��B�H	H�*�/������}��!���p�zw4{�u=����*����N�}i����ztZ�F��ﭑ!�f�������<v{fy�^�}k��0�2�G�b1s{U�(��oR�Ψ)@45NP=���*��@Sީ����۹�U�{�{��+���}�g9����z���$�}�O[cg�UJ�����}��P��Wg�o�����г��rz�Cڵ��uA>y䢼td��@}��@ 7����AH��T�*&}�p}���/x�y6�澞����z��Ӿ%W��}l�M���p��nm�l���w)��v�����k�ϥ)w��{죽���Ͼ��ҩ��g=��j�}��m��P*�C'y�N��>K�Ww>�ִύ�ƽ����Os۶jvn�7m���;w����|UE��7ݷ���<�+֊}�{��
my�9��}�>�����+��{�zx��P۴
�2� w�ʤ�
	QRB%*|�� 2g�>�)�}�{���� �u�@�||���seK���1k͏C[lޜy7U*"��{�.+]���ol�q洞|�%C������ѽ��w�p����=�^��PE?LT�PFM     S��2IT�z�      E=�!5T��0    Ob�PȪ� 4`��0�?�iUI�   �@ OM*�!	�Ojd�4iO��A���H�����~W��]~Cw)�i��ï�L�
�+6."T\ޞ~=`ƞ��;��I���z���wI�������$��/wI�'ww��I�'wu�?��o��;�>��:N��:�d�wI���OHN�t�N�;�ww������I�;�t��úRt�$�:LwRu$��'R�v$��ĒRv;��))���L'u;�$I�S�rt�rN���"t���'N��'t�:N�"I:t���Rt��'wN�);�t���;�:I$�wN��:wJI��I'wv;����I�$�t��N��pt�	�I;'N�t�'t��$�$����'t�)$�N�;�:wS�D���I'Rt�:�t����N�����1;�tN���;�;���ӥ;����Jwt�I'N�t��'N�S�tI�N�)��N�ӺRN�N��u'N�ӻ���9;�RI�u;���:JIҝ:N���t�:���wwRwS�I:�Iߤ��:N�;��N�N��ҝ)Ӄ��t�JI(���$蝎��I:c����$�w'RrN���蒒o���?�$t��#��W��ɔ˷�a��,����Dꏮb
��?}���}�v�f����G� S� �daeQ��@�ut�k{�h�3�o����=G؅�Ǖ��T�>�����&#8��q����O<���jQeS]mY=t�4����ʠ�Z@6k(!���;�ܝ5CYSo�P�n�@m�p2�ֵ�F�ʚ�d���#������:w�;t�E�͕�`���*6ir��Wx�D�ʖNC�]�=���q��Ƿ�н��LNN���)�y9����1
FD�ASo%�<1A�r��ǚ��P1�����]Ũ�N��*��b��MQ0Ṫ[b�h�N��}�z[��o�˫oy��Z%�����I�k%�����Y{k�O��/,�Sv-.<n�]ͼ۱$2�fc��c̓���,͸�c%��y8�Dڨ�:�kor��N�h��<�^-{�ua�̽�	�­#3h�[�kg�u.��e=X%b\��uڦ(*��)9^e&B�#�α	�s�����f��S�X��Ճe�L��ø�v.Y}�MZ"��ah[T$/��*�����}�م����+uD�cu�����Ķ��c4td��<��5x���ywxv\�T�e�%3H�@�ɶj��Z! SwT�U��Zx��!9	��j.�2�(����E{Y֩ d���ے�)���y��L�Ʃ���f�ɔm��O{m�w#b٬�XUʆ�BX�0�GV�ڸ�4�� w#��)�X�Yn�rLJ��DB���jރi6�9�U^�
�c7z�0���y��7{B�
���g�ѠM�2!Y��R���� b1^V�iW��В�p2:�Y��l��)b���� UG�j�qd �; �LS�T~��U��e9��
Z���`�J�^��_�ͩ��,
v��U�n���[�����E8�u���V��[.�&w"nԛDDр9�tFȍ!��@�{I]�I �3�풮�V�+	?Zwp����yp0����P�l����TǊhN*�.�.�n[!��vp����R7�TYQV��̖���1Ym�Kn�F��lY~_��jī����dV!ZSw.��un
��%��

��$���y���@�X�H朕��2�D
�5��pY/�pE�B�U)n���Ār-�ʸ:��a<u��fΝ"���ҚŸ�.b|7-�x�K�0e�
�e�iH��ZpZ��$7J~��u��y�ݬkp�[�;ܤ��������`�j�Ѵ�C��5 �4)��X��:�QԀ)�y5[���2�k6�݊�6��%C���-P�{"z��:Վ������vm����d�PG��|�Ӂ
8�&�N[<�(X#6�$� �Z�`��-졔���eaR`�5t�0&щ<���5S01.����ݩ��V���+��+̎�M�-�x/x�1`	q��n�tV�ӻ7�)7��*�� Q����qd_���fvƺQK!��sLgD�ʏF;t	��uw��ɱ^,��p�%UPӼ�j��G�M9b`i��0R��i�z�ᵴ�j^I�=Z�쥙Vŭ�Z�e��P�xCN�V�YB�w�T�F�'����	��ታ�`�5�hnbYcU�:��ð� �Q�BQ-�V\��Sx�p�D�2䛥�I���
r���)����a�˥�$u"�����e����A�Qab�v*��멤�e��kV��(?�@�	����#��>�������ƀ�32��w(����L�Gn�]_$�]7�1�����.h�+-bv���IbUP"���|����>'�? �~�E�ؖY� o�p��5-��Df�%iVC�1����6K��NY�e5Q���UY�yX��T�a�l�"Y-b�����w]۹��%&�R�1�N�n˴��V����@J�(�@c6u�n��)�X�d�K����"$J$X�f$ҋ��a�\YM���j��^2Ẃ"�#i�+A�q��(Z� �b��!��kW(k��������Z�IK2J{"u6�
e	�l:����wuúM��g2�2n<����Y�;{�ON�q�%Y�\�f����(b�AD�,���nR�w����x�����-�����dO Vwt��ӦЊ!�hը�n�S)'[��������=Ofk���`���TV�O�ŷN��Z��)��n�)��H�@�K)�b�y���B�Rdt.�,TF�_�7+-˴;	�,�������(��z�Qɠe��PK��܎�ހ�b\�S�S��܉�E�,C�Y�9jq�U���E<���Zj�(bi@�f�`Z�Tz�-Gu`�KX�c��Y�.�OKxS�Od�B������*\�&*1)Hd�P�[t/���s�TH��2���Bvݡ�T��S-���5���d	�:�vL��5Qn���l[1�s�fӛ !%�Z��y���W���!x):���0��ͧw5\Ti�{��U�g5��L�Ɣ7����j>��x嗮m����R�yS����ɝظ�K�a���d|�����f�(�vP�?�@�!R}��| .�;�}˕��W����,~���v�{�nqd@���IyY���hq
.�2D$��J�n�K���Qj^n�,�Ď�Y�<;\bKK[����Ni���l
Ŋ����8vI�.��%�ܳ���u0-�8����-��X��"
��N3�eh�o�Y��-�����Ćf�z2�n���3�5"t!����j���]F��K��]�~�p����R,][Z��Uyow!@,�ȿ/��۴��7K49���ֱ���aU�l��c$�m�'fJ!6�l�9��T*�v�)`Ǘ5�%��]�)��$�h�3z��d$*�P�&��f�1�b�Z��ζ�'c:���a����0���(A��sB���Iiݸ�yCn��{S{!�%����  ,��N5CY�H�ٷ7M�|)��weN�Oh�gun0�w6!g.�,����`f��ʯ�k.�0/�eh)�'�8R�y�s&Ae�X���i�t�H/*h��n&����*o"@2O��dbPs>�	��L0�F8�v,�7��<�3X����e	F��Ud�pQ��d^��a�̦N&bR�?1���� ��%X%,t�D�h�Jv�emd��g���a�?IMbpn�a7�e�zskl��!�*R{CO�x^�QS:~�nZ�ч,Q�DFx]�Y�s��F���yb�A���VB0fK$QX{2v�<���CRyI��6t���*�e�4�<hܨ���FD\Sɼ)��y#1jF�L��V�m���t�E	�`v&�,<+T�Ҧ�HI.����#`=�em�����{��p�QU��k0���dn۲���4��o�#嘖[�F�]�_�+���3�<�\�V��T�\�rf-*(�d�r��J?�+I�Zt��h-�e	U��*1[M�[���SG�e!Cq��S��0̇"��{HV��{8,w��.�wzn�(;�|�#\C(�7 ̝����&V**���c,_�X����]�*��j=�w�B��Ũak8X6R�Y#�M�voa܈�Srj��a��iqU)���`:�v6629tM���'�׸ �SkpX��K�E�7�2PPN��e�˴����eb6�Y�* d��i��TF�g^�6�7K"Tn� �t�Mi
$�E&L���{�eP��n����[`�jD�fmM�)G3�;�3	�:��0�Up��5����#��>�����h/��}�n��U-��@ovP�2U��8�_��!6�A�ko(F�0]�V��u]R�AZ��E1�Y��eҫ��/G$5.��;�3fM7,V�"��Ȫǰ~+ou���j�ɘG�AܹwJ�$�R]�-d�� &�]��g�1֕��ʵ�&!	[����fȩaJܔ��v̼y�	��.3����se�8�(�q M�������h� ��@b�A���ni�7N�J�VF�5 ��]�/`�%�XY
S�	W�*�2��W[^��\���Xz�;��V2�˾U���eɯ�&���s0qK��S�x��^6f�/^�T��ȭ�!�Qˌ��J�SCh��m�b5L�%����5�s6Tuj���̫��s�麮��U܆�D�21�UӒAW��D�h�h�いGCv�"��`�"�ʫ�������rax��\��,p&����'��M]�YO1��ǚ�D�nP2��07%z��b%�Ȱv�8�y�)&�L�D�-�ڃ0AN�Y/2��
u���	_�Q�����H��=KpD���9.:bV�,�)���#-e�g�f�|*],�,%�1q=J~ʃ5h��uZHVs�7�V��ϪLe@�պ�6̭��`����L���2���_3�C��f��kDq֐�cxM)F���M��u`�qH�L�6�­L5�T��m͚J�t���f�0�f���--�j�%�	YE�I%!��/X����hڒ�����ņL6o0��{{)���:Í੍8�T�`BU��d2�Y>�n�2��`�+{,W�����%t�rn^�X%��;2jCV
v�j�@��
b�Ճ(Ej��_N��.m�r�Ǐ��-��+���5��8R�ʜ�2��t°��j��͠��wP�ٓrij(��^S�p�D�L[
m�ٹS++|3�����!�6��3,���X;A�ȶ82�tj`�ش�D��Җ�$P���}�6���
ݮ�h���(,�J`r�����Xn�=�CY���*��6)-'ǻu3`8��5s+vZ��ꂪ���}G�!�e�)�D|0�=0w��F�RXZ��(
 BD�ໃ��v��)�:X���0c�#C��}҅��q%q𬬺{��ed��.�-��0�:p���'?Ij��V �ӓ�x�dV4���:\��WoE���3�E���f��f�w5]�Ok:o);dtY�����e^Vf=�B-��-�_e��](�i�l��2����%�]Z��%-�*��E!�7�:i/+{��j���D�On]�f�ls����t�:�u]��国m+)����q�
�a�Yu����n\���P!�����;��ՠm�R��D��s.��+h ]Fx�h�b]��U���b�j6���XX�O�PA���j��[F��#Q9ݪ@�=�A�_b���f�)�ӻ��T^�oxf��w��v桪 l+Vna�(����i�{�a<i�&�84��J�U��(65�ɛQ���k0K�+sh�W��ub ���A�+%;R.���E,F���M��2�M�O��l��W�0剶�"�GEM!
��6� B*T�k�.��3p�SR������� ��+�f$��SaVӭ�b�ͱG$�x�K�h(��qT��#�(F�5���� �Wc5�Y�3ei�WR��y�;.AE;w��!+�����b���Qs�A'3-�.e1fం�fQ����
�H�d�r\\aM92v���h��l��6�S+�����o�VV!v#����J�Zǹ�9w9B�A��gm��6�"��u�(]\�oF��)5�Y8d���o ㈲��.A8��J���nR�`�fɳ8h0�<�1j��Pմ�H�aZ�`	*�f2
`�9q)�������S��s52ҒS�F����,�J�I�˗t����p�; *^�c�ᱧ�iƔ�
�"Y���\d]G��B�e���xѓe�FYyE4ku���fv.��!�S�̤�%��H
H�1A�VdH�qv`��c�d��wE�
��Y�{���n7v�_i�2���8@&\:�T�E�Z��:oN.r��uej�vW+��e�:�(�8[�ub�TB�ZUfW� �jK�!GG�?cډ�ZӺ/sWm�N�)�HgX7a�c���t-#u�2����i\�1�oM��*�C\6F����g]\%n+36P$Xn'Pu���M�1�6��`��7*\#�ү��ܢz�;�f�Ym�b�m���iP V7Y)"�d�`�$&e�
���y�1L���|�*n���,[ձ;,Q#n�ɎM�a�J�P�F:1���&�9�&VY{ݫtQ�L�걃6��Ɔ)��=�6\�cvQ�0Y{A�Xɘָo A��!jb[��i�9CC�?�3x��O1�����भR��-�xR�V
��"�ĳY�P��4�Q�L��4���Ah	h�6Lt�ˏP�c]��ǔvR��L�\�H�3h����Iv�Pc���J0�C�{9$ҫ��NЩD�" �\�A�D�>Y	>Pƙ�o4+�P�'(��󒍪ڊ��`�-����<�*�na"�bר��kwM������.X�1ޘ����8s�<aPϋ;�"́V���*--�G1��]J�f��bBpA�uD:�9lW�hROr�$y�;��,�f[�s
ǚ4`#D��.�^�9LH�7�ڸ^Ch�x&�2r5k�Q,��BѬͅX?�� %��u��SԐ��*1�iK(�ou�A����[Pp�Hej*j�d�b�2S�X�I���u������+ץ�73�q�2��0!��X�r$(��ed9e�I�:�"�(���M�(�c
p����E)��5R��l�̧`^b��� eCH�deT7�#��Nb���-�JX@����J�wcL�h�H���ȒG1!�N�²��ȰB�blΫB�e��8m2��!q��M��i�Ls�34�Kh��o��\�^m����F�S�
��[n< l�M���ϩ�����@x�z��������ěQ�Xx`�(S��-d�k��f�V��;9˝b����p�/נ�7L�,��K5�1��.��\Y|�;�b�(9��NZ)��f
Ќn�D51	&K��I�&&
eA��d�Dw�r�?���?�2򿒇�����w��� &��ߎ���%R��J��5U�V�&�|�3��(��TҭUTڪ��(������`������25U[UP UUU�UUO*UR�UUUUUUUUUUT�\��*�UWW*ґ-UUUUUTQU]UH@;UUH!WUTUU@UUUR�*ԫUU��j��j��Q��dj�������j���jU�UA
����U*Ԅ�I�UPUUUT�l�UUT�P]-UYYV���^j�'5mUU]UR�U�V�`r9������,(Y��!�Ɣ�A���L]���b��7K�n��Z���^qֈ�͝5�t(R�s�ơ]N4�\f�)��]��$1��,!l�������gK�a�d�z�N8�qцeW=�<��#N!�=���긻�j�uv�;O`�^Ż]���]�cl[O=;��@$�	�Miq�F��{s���DK�����qK��[&���L�Ʋ�q��r���m�����k�py��R���uL�x���g+']jF���ll9����qK���Zޚ���d���;��K��>�=o	��ճl°�R6d��-�uk�Y-���7,�od0L)3�m��Mf}�uB�pf�hq�T�:��r]r�xЗ-��u�R�1�z�+�l�0\ dɺ��Tc9���l�Wvq\X,'k.;;�:���J}�5�p�u�+\��(h+��l�CZg1�7XS+�@cM6�#@���04�m�·Q�aON�:�(:::_
-�Sg�rr]@�h9��95!����a�Mb���F@��B�j�kq��ۭir�,<�&�t��i�=�=vtMÇ]�])��t����Kl�3[�r���f��קA��OL6��6!m[�,&�цh��Rǖ�2�l�̨����9֣���	WiW�����	���O!��C��ӹ�s�l���n6�[gqm8y3@�)��-�6ԁ*��M.p�fY](B 릲/!.��d4�pK�mf��1����g��bc���Ӑ��h[)��26�744�L��P��b�s:ڸ�K��5.���1v1]8����q[;��\\��GG����!ۛ��gX6�8[<Z�v
9Z�c��;�]�9wNku����n�S�� E]�s�����D"���LGG��ͬ�-,G\#e�i�3,T�ܭnfݙ��˷ZyPø&Q��V�p[=��uv�5v���I���a�m��c��H=���#���=E�	d�ۥ�@v^�\�D������I�Rۃ%�]��J;+6@��;2f��\�gMwhB������0��!s�Hn�q\g�M��q�8���=�7`[�"p�ԁ#Tl.l���	��l�]i���v�!AwU�Y��YT���RQ.	*/N�n�@�<��	�]�!�SM��(B�y�rh����O;\j臍\q�V\�o��6����mb�Z9�q�����8�"���m�6ۏ[Lt�vw����+K�m�[2�2�,,��&�ɣ��ͭ)ؽ{X���Y�]M*"�X�ul&�k9�z2��F��)���aHDsIq]*Ps�S�H
�Hfw>6q���z�f�.Cm�Z�2��q��<h4\�-����^�)�q�Y���LVJf�c�(W�k�b�5�-��&58�'5٪�0�y{K�ř����Y(k�ȇZ9����f�]]�Ԣ)������&ݩ����]i��;0�K�&�8#��`.=�Q�԰�`mnݣx��8.�I��K^�&ı�N<�v1uc�Fm��;;�K	����v�2J�º7&�f�2��u�R�mu-�$9 R	������)�/��J�sV7�����U1��l!'�r��ڝ�PuWV�͸�8څ����*V�n���z��n	kTM�9(斆Z��8Z�%�Ѹ�`8�µc؊�\��׃��:�cl6�W�6zd���a-�6�ǜ	`ݗ�K�<���� �{MV7btG��im�JJ6m֝�ՋrTj�Z�2�Mu�ec&�k	�KȽBmك�sܲ��v��nP�����kB�4�ƍ�\���M�:�V���!{gqʋ�.̗��:�V���2��1n�y�v�z�ι�:7m��*MpMu�#-J��*�ͨ��(zN��A���k�X �&���R]ٚ�CF墭�P����R������$]ة,M\���_\Wq���\�
7�U�
�mR�(�bR�)j�X4*Ӗf�R�+�!Ou{�ͩ�7td�wf�Dz�$�LR��M(��:\U�h0�lz3���h�x�L�\�e�(�J��4�6M�sF���uu��q��W*#L�@�A�ط�����ý�t\h�R�n�u�;��\r�,^����n�1U�����9�`e��ny�u E��ZŖQ��]Dx�ɦ�V.�I��i�x%&��e,jc:cde�iL��Ȟ<��|����up%��p]�p^69:�*�Z�rB�P�9��VP4&�L�P�53]��ƺ;]�������kI������U�\u�%�Ꮃ��P���S��GV�Zd���2	�t1)֪WW:�N�hKu��['-�y� �mv�Kl%N׆�n2nz�#g�˃{�V#��N�����b��{�W*C`��l�˶��Kc�!.81̝d��[ y{��2p�[��v,WU�< ��P�k�t	��T���Y�I
��'>ܶ�:]d�ݐA�D;��m����1�l�w0�i�׭�I�q�z����;zl�i{f��l�����*'C��6�H�qq�����-U#�ԅ������(Bvۇu�uqϊ3-����ް��a�l�fL�lhW$�g2�ի�<\ÍG9:�b#��z�-���	).��f�l%B5�1�4�lWf�M(^ڨhCB�!n��7�t���tF�į-!B ;1�N����Y�u��u��Xe 졺g�c\јM�;juBc\F�w�nrmֱ�(Liw$mls�`�\rG1���#�w�usۦ}j�7U���l�.̳P�e(�Jfg���'��<)q��c�lC]]�!5�Z��"�P�v9�<�wG�Y5;-�D�V�����9rV[ʄ�#S�q�����w����V0cs�����P�a�M�v�%�X��e	㫠M��%��qŝ��Ws��nOd4��b�����\[�������b���}����ݟL��8���$`q�CWW��K�5��k�2Bl�P���d{Ao!ۊ�3��ڍ�����V^Y�7e5Ӻ�4����"��1rAa�������6��n��K#n�� ̹�L[(v����''nC]��q#��۰�Ύ3���Zlg��v�pn��.R�m��;`�YK=��R>,�0����1���9:;;pQ��wPEB���n�N��:\
n76=X�y��0�LT �l5��&�f\fR٫X5�;��-��&.8cr'm���+��.�G�۷mEu'��H8��]qg���]��V�	�g��:�Sƻe��°�㐊䣥���mu)p%��k=�c5���5�s��u}���� 9[�t]��Hz��&ث2.ś�� "i����,f[4��$�iP
m�tے+G-�av��K0�$�<��u��m��8�@�� K)��[��\M*D�eƭˁ�m�UӋ�G��j$6��L�ơ�)��ⵋm���M�+a�M��m�5%	���D��3��r̮мdŠ���l�j	���:�={GTõ!��Ve�-�X�l,�[,`J�����R��:-��R�������{!� K������؅M�\���Nz�#�b"���8�A�X]2;�]qۜh�i:�!�I۶0������ƌ8ņL]t�h�Fu޷�&i�3��.!�'k����oh��5�'�d��kv=cc���g�t�(�0uA��H��ݮ�L���J9�a6�0cm�H[B	��+ˣ���Zh[���v��6�e947�6t\�X1�wfKnvV\�n�ʋgq� ��s�}�فk��Y���tiMj��U�GnM��t�N#�B�CC�N`:��ǆ��XEۄ�]f�q5�e�X-�aXL��jL��t�����Jcb��gnE�����Df�k;��npv����Ű��/s�}���\�w^����#Ce]-�f�B��Ռ����m�C�qͽQ1�ٛ@�&+tx����|��q�!�
��kl�,Vܰe��1ns���.�nvq����C����tr�ٱ\m�*�Vu�B��xM�Ʈ2Gn����\��y�h�;i�����	<7n��x�T�s��*���ǻ56.�@��	���)��#����by4˲T��Y�K�jX X٩\��pZ�&��CF}��$e��]Te�@�LK*0n����tj܄GF^�Sv�@�rk��쎀x�jC%����s�׉�ni,V�6�`4۬fy�2�u�
�%,B1��f�Y�;���R�r۶�ƺ��J�W!]>^Z�{ułvő�Ѷ�Ԣ�׹�W���X����6�C�l���b=�f��n�-+"2�&��Acl����K�a@��!ua��vA�V@ڢ�y9 ���l�n-uƎ�&/;Tm�`�*q���z�q��⭗��4�J+�и
���90�\�����[�.t�@a��Qڬ����ath,!������^x�܀��6SI�]v��Q��ڷ��d���i��XU�fYH�B�ত�-�E�^w���Q�X�102\�Ģ�gk�J�Rɯ�P{Vl��d!�ck+P�]tu"B�l�WP ��B%�d륻���J ]��ZLr�T��+m�T �������Z]@��p&��E�x��qb-�uv{\ԙ��bһ��GE[:
�X.��:�hh_��I�I'ww�����t�;������t�s����O��çN��N��������Ӥ�����O�����?t����'N_��N����{N�ӺwOĝ�'N��pN���I8$���N�Ӥ�t� t�8:wwwI�:wt�:X�B�1���!t~���k�z?��j�lٸ�����U�i+��<]�2�:O�;sS��}:���	E�77�9�L���A�(_`�q�s��.9[�ޭx���p��:jN����I���j�Q���P�*��	��7�U��'Ԫ���#��peJj�[g�5RV�h�˙W��7j��%;j�J�d�׎r�P�ܷW��a-n2){@��>Gtn��5V�@��������Q`����rv�,���ƙ���,B��+s�v�F2�m��ɨ�����@�[�p�߰c��N�p��{����Ay���}^u�@?W��/��y��p�w��@�"�a����w��:���վ��0y2�}���i���S�2��U|��Y&5��w���dH�V���m���,���[�Fm? ��
7�g����ϣ�}�_�X�} �/�^�~~
�<V�d��ڭ���������̓q�ק��H���"�6�f�x/�=���Ec�^nJ�Y6ߓq����S�����X�Ժ����J��z��-c��0e���ڔ��7\i`r�yYf���
�3T.$��ڏ1mgT�(nq��o�l�jݪ�]��q/�⧫%[F�T�&��6n�P�c{K��QV0��4"F�5&�+�gJ�2�z�n���D�#M�"�us�u�������9���9�����n�YC�0׌4[�ې��*�g�������v��-�:�dś��Dַ/[A��G�=b�
/��\�E��`�z��� ��[���LR0�� �T��Hg7̬�.���5sᚢv ���z����
G���b�$��d��p_���:�{ ����u�ď���x�o�f��j1P�@�~8�ϑ���2ؾ�����p4tL�e]4$�F��*s�=�U֮��{�:m,E��֓�JX�� і�`��x$�����f�:x+0ZB"F����7�{ӽy�=�x�C��Q^oB�j���}WA܅�(�)+4ڛDݡ���>ZD�h�7{��ﴶ,�������Ep��s��J)�w�����; ��,q���zX*PnC �y(��FQŗj��A ��o#���s}�ShZ�_j�׾*+��<�
h�P3hifVIT��WZݾ�]�q*���+�{ׁ�n���ĪO^O<��w���vI�����mZo���sv�����P3��~掍L"B���e��dW�'�U8�/|��3�~�RQ�	G���}���u��Qs���_T�x�+�s�ȇ�/k���e��.�ӜV�rm=��N�z�I�^:�Rml� �ޔiJ���F��l���@�6/�3압Ξ
��o���e�</ćrBۘ�wP2)c�Yt����y̶'���,DDH&�`�%��!���=�;I��������M@�0�M�ڬ�v�eý��lh��\���ت����z�K��<����t~��6�]�r�w�Ja���%JM��;�����s��zf����$v�(��lR5��td�V�p�.,���͏�6~Y�me��� �A$�G��+�̈s��c׎�vj��_��R�]��J��������F-��<2���z�ӻ�$��r2�g7����'	JH�.�]��;JfgEΡ�f��`�*�z�'�^�NCi3�ts�}v�29������Q_����~@$�!"�eE,A@�~�T���Y�*��Qm*�廾kf���({�3C��h+�{֝��fc���}J��٘e����[f
m7	�w6�ʕ$��W}�������W�{m�@�vh�&.�%Y�:�x^������Ś�8,(�.,�݈�Xv�Ù�6F�,B���Q�������n��T�-��{��Vu�Y6��c�K��7f�Q@crM*��ݧ����. gr��J��eLl�L�j$��1R�,J�^���u��ݢ`��;��D��׳��yf;�^�h��jf�I��9%�1�׻��@�5ѻ��Ķh�����Y����%�Pnj*P5�Faxi�s���b6��;H��������<>�7�:��r�;� ��C�c�����[�Qأ��`�BS��3��7��:rfHYכ�Tw��VO_��-�}��'�ׯz��70P8���w����ep����C+xOܨ��ZJk��{ݚ�ٱ�o.�tǸ�pukn�NC�+�n҂ǥ��N-Bѣ,�Ƨ�s�b/��z�|�1��b�J'V�[ih���_q�ػ	L��-_�F(���n.%q�A���nQ���MtX�/E�����Cw�4�ޝ��Q*���Y�^�Q��W������?`�}N�Vz��X�P�b��4+7�t9��׶K�_踨&���:6L\���ﶈP��ut�N��X�R�r��0M/�8��H�f�A�4���gQ�	槦�[���U�����%t�,�n��d�D��*t[�L��I�,�8;/�k?#���y�6��d�U>�������G�$�/���rޭ����d�zW��ب�W&�Y�VA�о�[��m�K�͜�jv��g8���y�.������h-B*n�r����oV�W��U��>{�5�^_�]��� �
�
��Y�k/<�e��x��W�˛��蜱2e��J�J���{^JS�⩌�,9��'ٹ�k;u3GN
v�t́��I�\ �I��--(W��gwD�w�N�N�w��̡K�?}k�a�:�x K���r�]���X����\Q�Wwt��'K��]\���>�p��x��=�LCU���sxT�Ԟ�[Yv��`Z��`q����t�s{�k�zy�g3gy���7~�"-wl�e׬���\��f�j����[�&7^�ƫ��H�	����gP1ƑMR�#��]0���қ�ɳ��@�ܻ���J���K�6��ޱ�ԭ�Mt�y�Z��Thkp�q�̽[�y�A	G��:/j�8~z�|{�f����l�~岯��J׬k�M肷�y@�Z���%����α��;2U���<�F�p�WE�
�LG�3N�쵐����^r���f6�b9#h�ꣳ�n��\L��#|�C��oQ��a+k �l�z���'7v9zJ�Jqv�\���&�Ŭr��\6,�n�OL�0�;�v5=n�`�X�I��<�v��Y��� f��-L�ng�l�p�vn	�ż�掳�[�v��=�ӌ��Ku�rR=����������Y��.;i�b�3˭nָ�b)^8�,&r���N��7�����Y��jV%��#�ϯ�n��t���_�N��Sq�a�H�D�;��V=f�ڽy�~��=��� �.�zQ[�����fL,�o���)_,<��0�ήy��g1u����\AS�%�I+$�����=���G�~����oX%cr9�����	�X:e�ֱ.�3��H���Ki�vhڑ0�" �G���F�v�;Y���Z�׶ǃG��-�>��jC�=�/OJ[�ț2R��p[3�ggm�b�٠�=��v+o�4�fa²�sL���{��x3��?��íɻyL�iR	�E&���k��->��ĞB������yd�[S��I�z�����"���i�Z{�٣��ÿ��K�S���;��;�N��jϨ(F. ���a]Z��žg�8[w�ݞ�f
vF���N�\������ܪ8yŨ[����-n0�@���\�
v٥P1b����ݹ����íq���<Ȱi��s/(=O}Z��>vjX�ں����x�M� ܇¤�W���D�&�\�Ve�z�0gf��oz���V��1����')%�Ъ�i��.Wr���*�^�[7�n|�BCWDW��k��fUw9��Qt���6�n�I��a��v�p��Cs\t�qڮ1)�i�-z��Y�Q�X,�	�g�fM��&����z�u�wע��S�Aŵ"��2kv����\B!��U�d(T$�f-�.P��T��������Z�o�'�����|��VZ�6_�Vu?w^z��:����DWd�`����;�͚�7ڡ'��S�n*[\mȃ�V=��ke:�.+Ҡ��c؆*>΋n��������6���T��4&�U�����é�_�˖�J~��&�����"��Y~�|�NG�˥�Vǣy^^s�����O*�*�D�) i�Q���@㫭FXN�i�7F��k��j��E���y���~������V#�oNY�kĮ�"t�/;�׏F�&$Zi��m�|�h=z7�9�j�9V�'�(�=��_1z�5]��cRЎ"���d��J
.wI�4�f�A6�[9���jԍ�ͪb�P9�q���Qw��̾=���L~9=�������v��]���U�Cf_g#V�y
x�b��.�4PSOg,���� ��ܭ��v�x�.���ԳyZ��EӔsSH���h!��Jј��(ơW�v"/}XN*���~�⩗���=���b�KgI��R{;�j�ه�cdlHe��m�.q_�gu���
L |u
��w�Z�ᙤpsWe��w�Å1@Sa��^��7�CW(��Ę/�%vc�y���a��j}����[�����J*6{�⌁�j�ջ๛U������p�-2�6|qe|��HD�������u&$LF�h@�G9|����}kͮ�y�^x\��lP��-��G|�x�F wcL�s��so�ף.��u�z�0��һ����M��>��V�h���i�]np& is
l�)��ܡQ[]r�9�Yp�g�Ƴ�>{q�T��RaH�A�����ai�4��+���+ O�Tٳ�j����GfI�ٸÉ�\�p-U�J���T^'*L��Ø�L"��b���z���?m�\�e�8d~�{2�n��rޥK�-ҡ�v����k���,��TH$.�#�lY��$z�9�-C��:gil&�=���L���|�˙�f�v��n���]��d��ih�N..�C�Q���D�&����u뛮�dk]$k�ox����pZ���9YV��=�]� �N�$�xG��9]ᾦq�Bq�a������^�p��}��i�^���� �i��Z�8J���+ �;u {��G��-y�ɺY0bL� �
��E٨��r�T���|l�ߵ�Պ��}Ǡެ/=�\���.��W��Z�6ƚ.��*-��)c,�XR2��E"�W5�ʘ��LC��K6])�pr%���(��a�@J���>��j8Eɮ�9r�AQ�D2K�fw3.���vT{⧛V?[��Vs{}ƅ�ڽ�6= ��wقun�4��$�HZ�` PF���='voot��ܫC<��T�� ��2?g�^���ܹy�0KS?[$K�#�s���P�$#�w������ѿ�W�Q�=�1�Z�cE��Qm��>��oou;ݲލ�d�6�Ž�0^���;���U9�V�4��v�wf���u���@�ۆz�u�s;�7u��9�����%z�����cή޺�(Q{�̖�w&IO)jZM,MP��U8n2r�e�/�o���Ļ1�Q��)5Z����A�i������~����Ͱ�����ʽ�g�}c�F���]��ļ�ڨ�:r�ZƉҜ뵷�.�K7o{�4%<F�]��X�%� ��I�F�%�2���+MZKk{h���&fq���g��ܤs�������f���qlz��Gl����Cd�s9�˻h-��UN��l�ތ��1��qj�8��.�4A���-јð��kj#�(���D���Nn�ٞ����%���(���`�Dw����w5����!����d��(���p�Y^IH�� �5hp��������ʧ�
��l䗻�_e�
��U!]X���߫k�0e���{䱦e9��J�
H�t��s���1���gb�������m;�]qY���T�p]M�,om�0I����i��a�n��M�E��k*I���N�����79��h�g�(vXhb�ld孚ǜ��mI@�u*
��J�4��ӗ}�s�K(f�Q����&b�,h��kdf��<n]=y�6�Zn�{Q�Μ[1��%$
�[��P[��5Il��̵g+�xA��fJ������~��(y[��E�~���oy�Ľ���`ݢ7gXR�I��#k�N�����;Pf祆#q��uj|�jj��;n=ݏ��ޏ_i��|�bv���wj"������p�jjq���y�kV(��� `ɸ���:��_!Y�wL�w��>�Ͽ	� �I�A |	$�G�Wj��FS^�:�!~1\܃�|��*�r�=�r�]]v2p�嚏�ˍ�e�W2�ʽ�h�K:��N�Σ{��o�ȋ�z
v�ٜ봌�fm`2z:����`ڗ�f�|;Kr��y���� }^3�3�Q̖
i�k�[(��r��Z��A-И��~9�m=ŝۊ����G�gd����]�ɸ�j�Ss�WWt��7��n���v�@RB�\g��2`�w�аP���ŝ�c��y��2��I��OfViG�-
L�
����О:*5�7)��=8�Y�C�f\�|�`Z�v�"6˩��&br<�M"�dȟ<W�.a\�쾓`��uk����(O[��<�0���R���)�ajYtu��I��D��B�nw���Xy"�B���+!��b�k�nk]�R�8���K.�o*��H�o�7ӆ�D�U�o]��i{˶U�o�ھ��t4f`z]�3/�2��;�tu�ݙ�U[h�����6��m	�q�����{dp�a��*4e�U�mÙkT_����k��s.΍=���p��fggZ��wh�/']�X��ű�a�r��i�P�@������lH�!��q=Nd1��)�봱�9�&x��I���Q�1�c.���u���M��`�+���Nu�re	:hd�_���Yv��V�ޒ+kv�-��K?����^Ƹw����Kw�p�%�-���)�^�[��:V�;Co�T�@j+ڻ\(�<L������L���&S�7��䍨UuY��Um*��T��UP@UJ�R��
vUv�TQŧA[X�"
�T�:=�SS,77k�^f՛�quڲ����Hp�=�F��vX�I�p`{;�k�A���yr�n��5����;\�&8�qVںc��N���.3	�S�l�hTR���<s�gN�&�s��#vc�%hj&f�[����V�W6|݅Jꗀ�Q���+��&�6M��Wu�w1�����GV��;�y�b�9�컰,k[�6���B�6cB�B��a8�V�ٵ�[a��'P��fϸ@Gu���\�b1^�2	�k����c!��*��0уVK����+t��F1����)��:��l�Vu",#W1t�*^�Hm)��0&�%�m�v��z���$ N���X��ŻM���p�Zw:73$�l�1v�X�w�s���{I<�D�A\jo<�v��=!�HNф��I��Ƒ��v�T<nR�q���'n�����i�q�IC5�]��D��6��1��C0�����qƻmq���W�m�Zݲc���v#�����Zŭ��Ѷ�z��Ň|dawl��e�u�n�AN۳Ր��6����=���H����l�I���d1�'���7	���D�\s�q���`��$n1�]/:Śd�9�iz��K�le!F]��kL���,<'.��6�x���On�)v(�]�#��a�h�iN��WA[n:�m�d�s���v2�����c�ܘ��[q��KJS�N�@�3ٺ9�v��pX�R�ݰ�������kq��+�NL�6Έ��i�<�Ջ�͝s��ɨ:�,�˘���F�1�$ԭ�m���Y��W"<���j�Ў��CL��N �vc�(͘��[��X���y�KA�۝	`��d���N�J�Ѝ��:Y�XiBu��	ia�@vj��bR�P���S�1tk:�-����\��St��m���e9��:g�vG�u�]���T�u�EMJ}&I7��P��6a@��R���Ia�8�Ca�^y���2�%���
H�m[��oTd[��]z�ֱW;Z���v4��MՀ����:}Ԧ3i�%Ui�3�uf�H�8���k�;_�j��'����]�,}�\�ۗ/+"�9�Zp.=���$Y.A6��F�r��(U�1$���Of;�V���B1Sf�<s��kXҗ�23r�o�L��-_4��C�_̟s3Un�[�����GOʷ��%	�y����C��많�#$2����e�K��Q��n�E���&�-��0��}�m��^�F�	>���Y:�X�7j}��yÂ�,��6��3�&��~��㏮�"�y���04�՜���HY��w���i��ͽ���ضt�{>r�ER�M�zSkVm���f�](�6���C�QIJ���}XD^��v\�8[e^YNHf����t��wJd+��O37�ә`G�dU��ˈ�����>pNe.������$�0W��m*�������aV^r��&9!=�;o�g�#�u[��	N4ژ�npP�4M��3%�\�.��i �!p�mc��A9��u��܍�fN����|���UBc��0p�$h���ǻf躱�8|%7JFFJY��DS�����t>���V�+ECr ��<��#ژ(
@�w�t��Sy��$�o'p�k�r��ڼu�;��
�HJt��[���R�XU�=U�G.C�x�ۗ>Q�zīG�{����:̸�Ծ0"�v�m�%ɖ��z�����'� IRI+$���s����9��$#o��S����XQ�~�`V�L��(�8���s�le��u�$P>����b�V�o��k���j�2�ynT���:�s�,�Z��UՍJ�2d�wq��F���<W讬��^�)�)l�%N�հ��P����3Һ��a0�}����ߩB��K{;�T��PJHHA�	�&��6�)���yb|������$>��/�V��`36��LZ��럟��bUE�57�#6$��?:�Yn�FQ��_q�s������Oܜ1	�$�Vj5����T 6T�s�h%V������8ۀh �rk=��g$vy:#m����{�CrꮍA�XA��ݪ��Q٭J�k{yI���=�XӒ3�����2�D�V;�ܵG׃u0�p���3A4p̐�:��\����lE>V�h�M�?P� �p�ogW`�	�����OQ������Vg���n�9��ҺG{�P�7@��*�4��t�m�K�c��(Yҫ�ԦgD�8��ע�-D����G�o ޥ���B8c�xv��d�J��S%܏m]\RoS��k2�p��KA6C��`V���k�����4��\�<��\�(��ۚ�u[����+jdf-I7og�y��Ǻ;�� ��ԉ��i��:��fV+�o�D�@O��j�C�,J��dĉ;��iy�)�.�*�������1�t !��m>3�����ȡZ��슩�� F�ґ�cQ�W>��y��nq�;�yq�zY��+�/HZ k2��b�<z���=yo�Ǎ��䷡��`�oݶSy�'�p�@�<�(��Q.�J��:4��!��&z<N$�d^���δ���Q�W};}P��ȅ*	��n�k����ω �G�%��Ұ:����L�LK��T�v.3w��Z2{̍�]������b�dM�I8R�;%"�L,�.S����oW���,���R&$&@-�FcG�^�r=�׎��-�~Q(����/��)M;'�|�w|��_�x=�9��uΛ���9�0�:����$U9n6/3T(-�i����ۭ2�.�+2��=S+�P �nf�?w_L�*�_���Ζ<C*<zﭹ���4���t��]�s���%���f9��3Ww1_U��ngj�v��F�	���V #�=�DU���D6M������G��w)�{5�jXji��wvx�@ۥ,�#�;�=+�
ڼ��=7:wJ�{i=8K�����[n^�Mf���i�9h��Z�}Ŏ8:�Zڮ����a����;�lf�۴Xinmf�z�V,
�ձ��]E�;�n�����P`<s7<���k�i�%�ת��Y|Q�5MMq��ise1�eq�&@$��C9���u��.���ݕ�r�e�F�N��ǭda�Z<���'��sc85v�ː���i�o\q��QgU��2�cS3:�u��ю��L8����0��(�j	q����'p`����nY��b����̬.���ѼV��-�	�f���&c-niSE�R��遹��n���GؽKς������H�H�@����7���o!ԩ'�k�8�.���P8׋�,�V�z��g$u�nFQ��]	m��tz��Ow���-�\���>�`,�]�(2�-�˄!�p�rƚh<�� �V�OG'9��"Y���寿��{v^�"�"���snL�,IcIXF;���68�������=��j�����؜����B���=� RZB�f{0洐IN�X�k�[�&���?xϰ
@�c��M{)=8�Uރ�% bBV�eB�%������y���l"�$�i�(0q*���n��W��>"繮�KGZ���j�	�C\ƴ]�|���9W��դ�G��ﷶ�{��]����c�p<bܪ�:�B�J7�`*�c��9���ش'�zk{3��l$�J��uֲ>��ٶ9 �}����1>�K_M��^AP��O{n��Q�6a�aK
��>����0n�Fu�P����Bk�=��c@��s���؞�7Y�'��&9������ɿ]]*"�s	6���{�)+Z��S��"E9P�9a+f�ܧ��^=��6��r6���1r٘Y7�l�ם/({�x$��0"_T��g�p�Yp�����8�����^�(���(��Fn Żڏ_�ussh��nY�}��W�s���c�#O��tIF���A9:��.�w[6�>���s�nG�V;C{�(/�$
[Wc+��@�l�o�q��t���o�>� �e��P\�⮄ؒH�(5v���G��i�>�U�X�9�EȨ���> �}��P���㏹����d�#���zDN��:�]���y�����iC(�T���,��y����Ӟ�!N�֪t�0����$�e	�C�=g��
v�{�'�]E�W&|-q�ղ���%�7��Sfv����Eg�H��d@�sФ�K�ƄX��HR4{l�v�+2R�v�p�L����;4lt7~S9:��U�0��He�Z��RP��Z"-�BI�м��kFޏ �#2=��6᱈���c�D�]��ZUh/�*+���Bk�b[JP��1Ҏ��P˪](���4M��O����f�^�"�A�\P]�E��rs�qs�Z��rF�
<�n+�?lCFs�fYyuZ���#	���h+�(u6�D��ӈ%���!�����j%ct8s�sNvݹ3�0��ڀ��Qgw�]�c4*�$��w}�yzY�y�����K�t�|R��9�-�ۣQrH&��_JH�f�פR�G�l��7-Z�ߦwY�lj���0�W�5�Әf���5�-��0UG��l^�tl�����N�3���Uc���<(��խ;��$a�p���u��R�Rx�J��,�F�d���P��3S%����H1L��B�b�y��܂�[�� f_{&п��`�9�{3�3Y�4�9Pg&5��u�NȒ���1s[rɜ�أ�X��[�j:̹;�����p��ɞ�A�;�i�����b8�ͥ�i��6].�{O�J�&0���[Wx\��3Ծ���G������B�cS6���娖�H��a�p2���p-�wO�ԍ^ph�tE,59'8k���`V�u�����@o`�Z謓��7[w�j����f>dL�&��[�a��
QיȶM	0�phe�"���;1���w�R�"ѵǙ�y:3������6�u���a�v	�@imIA6�Q�b4����H���D�$ Q��On�4 ��*y=26����Yqs�@m���֮cDx8������� �S��ut�����w�tCa�@FU$7W���܂ӛu�x��L�2tdP�c=�*��J-y�Uhz����]p,�岱^ɤ�"$n��:*`��ڿ8����wo8z�kC1Ba�5~��df.�_Nw�h���W����v6�GB?��Ǝ�8��~��`}!����a��f�4Y����WgJ����m>/i��J����
j��bǕ�|.�Q���W���B�_��� ��O̷z�w�gX*a�$�[�����[+L��P-�x�h�՗^��	�R�2{�lq��s���U�nC��;��ȟ4�:��2�ßo;	��TL;��Z<�̹�����= �A��a�M���յ����q��������E��G���b�+�@D���؟Kr<�t��0�ues�д6�j�ܘ��J�O\W�����#sy�Bab��CP�)�ɱ�舅E�w:������|�w���k=kt��m+e�S��I2K��/ -�D�-H[*8R���W�#��ܖ��s�\E�|�����LH�Gq��e�y��_���1�q���{ (�<��������J��u@�60^fSjn4�Bg^_Z{j��1�;G>�hb=t,Qf{b��\��w�دmN�c�0�f�����O��4κ;�p��H=�X�Q(���Y����+j��:�;�p�ܫ��AYk�`^<鴴��4���Q��������n+>�{mN���jW��݀C%7թ:��>�'G���PG�-x����|������X6^�ߊCX��6�I����a�y����@J�]#����xWm�jھOK���ktV��^���Yt�K��ud��F��*�$]%v@d�!�{q��4��w s��Y�_:�>	��wQ͹��IY�i�;�.+u���sĊHݔ�ńv# �`���l��q�+	i.���4e[�!u��b�v�*
m G���LCM,˳f݂����.�ղ�v�.�G	d1!����"��j�c�0d.5�f����	�:��rv*�� �� :RN�r���c<���b��~������~��W#�k��Ņ1+�>���Zq���Mo�W�:�^3�4�̦�K�m(��洑�0rrƮb��w5o�/xn�B���e�XQ��U1�Kw�Kt2���.&_a�U>g�c�E�x��`2�ʮ@��H,�����H�k�U�?�������(��(Ͷn��Ub"�Ѵ\p=�u�<�r�U\=��x���	F��4$-ؤ�{:tzF��fr��L옎_���Ok*�G�塶��I�爵Ѵ�;����N	e�@PQ��Ұe2�݅�2�mT��
�����S���:���B�0�d�P����`|���"�S<?^\�&���Ѥ/��hb{��F�^p��i�Vn:k���'� �Vy2'����]��j�Ӳo�\
S�L�L��qb��y}�M�|/4i*Ҝz�.3��b����<�η=�P/��#�-�-*T���/�%��-��KD��z���'����v}=	米p	^�U��}���0��Z�F4Q�칳W�qDW�A2������p��%��i���]��6*Pbs2�چ����:�77}A�$ߕ���>�h}�a~���1*��8x�V��n����#��$�z%�ZL5rQĀ�i�ݽ^TzܥS/���p-\�nT�����0M���Dr8W��4cO�����Z�Y.y�+#�!g�}xe�ϸ�m-&�Istߪ�E�{#�޹�����m�ݧ͋����LJB�HTqI!I�	�,��Ӟ�fu����6��!ಃH�Ld��g��r����u=� ?g��&���L����=��|"X������}�)=�f�`�@.l�I6�aMI#��m�b��x�&:&F;�wu�x��]Lc3WΣw.kwJ�����4]��S<PL�A�;�ީ�wf��e�A�0��2��w$[^��Lᓷ�f��S�^$뛪		<u���8�#�$
��|W�nY��!���h_{=qpQ�U�s5ݮ�Xk��}���s�n�"� ���%U[��2��f,�� �ޤe!�QT���gdyח�h��I��%�w�����b=*0F���LS?/'��܄K�,�^s����T z.��
�i�Bjy�0�,�}��-���%�刀��=�2ȗ7�=�,�\W�>��[{���f޽�O�o��^2��Q9G�V�v�b�[#/ʺ���A�ȰT?�M�_�b����޾��̚�G�I���s���Ҵ�	Dg�2"-$�R��݉hK59��j�h���[Usut��>�a�;�E8��{�@8�nl�TJvz�ϸ����Y�G4���y�ѻ��i)׷���d���·E�y2)Hq���Ơo;2�ۘ���Gq�+rI1���p��1��4��r5^�
o"Ӝ��jn2��X����JY��+�Nd�D%�Q��]�rxS���Ds���ި�y�#5�`��	 c
U�VJw�>�H��>}f�t�q�o�=�,�ː���<�yhQG�T��;�_�P�c��9�{;OY��!)
	7^�f�b[j��S	w���X�=%�_�
1{<�+S�]�䦜nܵ�)�q�F����+�Ѳ~%d ��H�L0�*ֳ]'��1M��䘿g�z3-�r��;�|ٰz2O��M�������T�b�wU���K�ɡ�a��oo�YM �6��M��Y�t�ji�;zdYվ�\9������<�;�yY4���
-{ڣ�?nNyZ����F
���*�߶��>�+��p�hmC�S{�^v���
��I��/2(/٫٧�1���h�rSWQ��c���r��S���F�A�L�6ȟ?�hуuh�i��ۮ�@���%��Ȩm�PvQ����}>�c��(9\.k�f����7a3c9�O���wp]����8&�__���w��GO@p���?\23�F6΋��x�lfscbH�Z
����E�U��ioNc�k�^s����H�����9�E�m��@��z��`^�[Z�NL��={-�o��4HdN1ps�w��%�gt ~�S�L9e�C�z �VվU�!]�2=�p��g&�ԭ?	�&.�
8�X�V�Gt ��c��f��(����陦pي�X�cF��uIf�2�]]��6ْM<��3VͲ�"V�˓lk�ڑ�Z��{qJ���]��	��X]��sY;���s�+�`�{.i� ���r�TP�W:2��Ĳ�Hg8����=�Qy�W6;� c���H�ެ�Kk538�\�Uz�w�ehKڝ�9W$����ǋ0�=D0K���ș��U�~��;����w3-���+��uR��	��F���(J��"�<�Ś�nر�P.:������L�ٕ��s*ݶ�uܬ�%�ݮS;�����ʙ2�/e���Dz���aGx<')�Y�b�����և�*:����𡊍ge����;�m.wܟM�з�A�A�{N@�^z�W6M9��f�l���s5�8�Q���dȷ�3{v���WX��B���T:a:,��(������[U� k���fF��9P��H��.�����(��ZFޢ��zZ��poF��ۺ��P��-!�׌+���;����J�eoN���n�ُ�l����Ɩ.�<2�zT+&0��O6��h^�kR��_�.���y�6�[����R���)uX_����C/�n��P=ś:�-i�Ӧ�3�]N$b;j�f�U���	�2�˩z��S����
�Kll�ѳ�G����UƟT��� ��Qb�Wm��*V��t���H������Je{d\8�-�
�02o{r�)�����znf4�5�p+�1�s��5�8yN�I'%/��R��<�H�d��>�y�I�˪��no�pz�c�]�N���|�����8O�O��z���U����Ȍ�-ĭ	�q�#I�f�[�n/�8A�MEQ�d����!�ږ(w�f�M�f3�X�񌩓�g�	�#����]�7�5D�ƌm�+���oۍX�Γ[�h�/�PN��To.����!��^�Qz����y�|�y֡�.���4#C��T��߿����N�Ź�x�t�0��)�!R;5jBۆ� �6�&	������vncu*��ePќ�&��ƹ�>	�����|�ɑ,�F=7�l���ħ!v�����;=R3F��X1�	q:��{�V��0�/|D)��r����ߟi�[��l_�Wټ���7�S܆��c6�09�emgR�ht���=X���=���%��i�Eg���{k�^߻n�ws�Ξ���G�@f,�^��ߙ�h��q�j-F�* ������& ���8����J��.�w��
�+���j�G$��Ž�$��Q���L��6#
�\Ժ���%��S�K~�����#-���d�V���J���t{�r��P��i�s�Wp@%��^���/�㸳`}���J�v����Q��U<�nBv[@J;Ǖ�]:��{sHF�Վ� c���k����h�Ff�E�r�@�K&	�m
u�����x۶-���V�u��n)�l��k�i�j�i��T&�:�� T��Em&�ΎL5��gL��5ʰ���]rj�iK�BQ��t��b�j܁ێ������u)�����x�u"6>�iO��]Kj����|�u:k�M���ͱ/^R�~c��s��>o�q7a*E�+3g��C4G<*_���;s^�#GR̩�7)	���o�%�~��Me�K����Cs�O1gM���m]նoO�ϛp]$��;�T����O��>�B��������v���W\O[�띆�w|%C)�ȡ1�@�D�-*�iK�Mr9�K��v�E>�y3Tΰ�=?B{��0@�*��t�׳j�	��z�,�xg��w�{Mí�i�����nk�a8!HN_pU�m���^eg�d�jDy>8�UDN��7jo���Z� h���*m�^r�ۥLe�t.�����(jP��K<��:Q���v����B��f�C'�g<�����WFa����/%gM��d���| �<���<W�Y̟"��߀�� �����y(�}=��Vl������#��^US�Ի���h��-
�Iנ*l�<�w#{��:��ٖ�ҽ��Z����6$*���rvFr�q��h=�8}F��O
���O�s������C&H�m�bXbi�u�)�U��%� k{��LXs@\l��ǽיwxk�k7���N@�6���e=1�m��B��j�� �*v���2!;*.+uY�� �����YZ�R)�԰�V/MŚ/o�6]��>��[��=qf簓k{�J�0���xW<�ۍT�GGqE��^J
q��V�賛Y�v*.띧U�H���U���8�����\\9�Ff�nsf���d��ݮ�l����#��P��
H�W��ڋ�GT0M���Y���⢹��/H3a:o�PA�7�'EDG)���B��=�f���#&0��6c����L���S0����W�<��=��3K(��,�BSI���Mn�Op�D��k]wd�؎�+�ty�u;�㣔"[p%X��b�]p�f��	Y��Ɯ�9��bՊX�q��2�������D��Ň=��5��#�3�
�-�f�s�R:��Q��V�8W��y����LD� ��%_!pdc�O����Ay���a�S>��c�>��%CgN��B�����W�pJp@�8 �>0�3�3�"�p(�ub]o�$��� �P�D&�=��?h��8�79V��X�Y��m�M�12<<k��w�G����V2wzv�zZ
W ��𼃛����P��ny��J��)_x��kOp&j(�Bh
2s1���<ܺ��׵���ޘC�X�8:�Y��P��f�&.3�Ԭ�P�h�7��C� ���M�A��0
��v���d��ƨY�x��T��W��`,",Jg;Wn���HQ�?mGi����t�Ո"���<ȣĳr���{.���I8c�!�S�$y��ԙ�ۯEf�<��;���8���(4Rwr������f㑶�{9[�Ƥb��;{����(��O�Xj��إ�3������G���f���/p)+z`B0;�����|�.�s��~�*����Ѝ��)�S��b� ;_5N�
}kA�_��e�4r���L���*����'�� /��Sd��ކ���ket[�C/�+b�k�܋�k.F<s{� ]7�7f�/)��0�H�O���BO�_��D8���)P�;�*�\}�L8��������:�z�r�8&M-��f1h�s�zvb���>�~ʸ�2�
�JC�F{絹uc��'�SqY<����Y#1�jɟ�nmM	��W�{6���@��"���?"Q��	��fn�Bi��f��7dׯ�}^��z��>u���w YQ����0Q�|6�?e�;�~��<�1�[�H�q �"|�B-��Ik�ڳ���]T]��ۘ�¢	@���AlB��i���񯕌`]�^F���b^�d�LL��} ���C:-Ӹ�]97r.�����uk��x��.�@�
D����D�'���N��^nZ>���V����i/��^�1�PmBuX��1��S[]�!Q�xs��|�������5~�Y�b���(cݧ����{�ʻr��^�̆��p�&YL�i��@�vwͧS�\V��J�#9Nѣs48Ө�wܮaǴ��69c�K�ddV�x�I����}{��+�5��1k)�誇Vh��E`v��7:�5��>��X�\!��Ɲ�]��OuZVZ��[��xT^����D&�m��}(=Sw���U;�0ˋT ]sId�_w-��N9���TBe�}�<��ES�+;�l�����7�����v���f����+-�u�$��e�Q[G�
��W�}c�Wdp>�	����<}��C���3w��4�� �b�ɀ��v뙄5r���;��%<�پa?�A'p��������=�S��^�֧���AI�	|J�a�Y���]��e y�lϷ#'�|�AD\˘���=��8���b��.��-J���VǪ���]I&��Q��F��~�������W�캕��g��3�ف��d+=s��$���@5�s�5ݔ����y�=��� ����.M��ޫt/6w�qJ�}���"�e�o��S�2�^23�*Lu?�
�!s'^?�ғ��ޜ�ivK}f6���8|�`M;~���D~�X��4��E组�O��=o*���0�u{b�4�=�o2�$����YG=��A�i��>�����#g�G�o�؜���转�3�W��`-C��0�h�=�5�+���o���5e�	�j|g�f☪T��h1�տt&&�x}؂�>������:Mu`��(�wW
K3f��@�I��Ui��q�S۰�]������L��L���?5�TT�]H�.�s.�P���0���!�ݮb�0VӍ�μ���,�q.ی�q�i�G��5�U热���*�C���iĹ��E�c���c,�靿�?0�n�k�l����LC'iN��ˋn����v.�a���I�Pz�8���]h=�#�M��v�cv*��x��^��h�����i�����4 S�H�R��������S�7��]>ڸ�����d8�^�'9����W�I��P �l���6�q�n�����8�zr�Ydu�U0�g�o%!s�b�p�N|	/�c�^����N���O�`ƍMN!7B����1�8��g`M�)��v�XY���%��*����H�Nd��s�˳�'��~��Nm�n(�֧W.Ͱ��M���B3B(k�� ����0��C��=ݳA`5�=�����aw������ ���K̦WJc)::="{�Ej�'}w1��d�"Rb&��I嚎/Qv_����f�I� ����#�ޡ�.y����U���O�9x���(�y���=��WǦΜ�L��v�����3{뻪0���x0b�M:�:em
l�x�7w)O���M����?������Ӟ԰eR�����?O|������I5�}I{uf+=����7٢�ƣ�R�t�s/�W��pp�0�R�����RpYօjn��4A��iuj�^��^������m�t��޴�9{x�Q;{�-���+�=�E�>O�h���t��{=zZW��^`��Ww�O�q#�N�k�ާzz;貰mb�d8��y�ej>���ޘ{�췰 ���J��b��1�v�/i�\Tf�y��PMG
�7H`Źzf��a���Em�'b��w��T���v��L���8#	�1��Û�F�n���MZ�nHq~��Y�Z�bk-9�	G�Q]��wL�vA'����%
*d��.f�2n��t���P�<�g�:Ϝ9�{�?H�#����Ǯ0��`�h��GF�b�V�H(��d��M���T�~��.w�pZ-\pjM-==�8��eY�z�Lg�r��#c"�y˒}���� ��h�e0!Xdy�� fVeM�Td�E��ъ���Z���u1�]3�%@o���(��Z�R���1�Ϡ@����f�f?Z��j�F�>]yY6z8�Ja �pa��L�x��R���}���x����=��/Ѝ5q)]Wf\`�0d��`Q��,�x<�Je I��f�q�����ΣY��ݖ:�azO�9}c{��0�Im��y�F`�Pӹ����a��o�rz�z�� �g^�|���{�|,����!���9��O�|�XҤ�:�{��P������"�A�����$�R:������LI���[n�J"��ТE<쬮���� ��Z�� ��A�'�$�
�(m��<�|�K�U6�(m���;�k{��2@�]u
�vζ�ra'�C�+&�� ���k�yZ�t
���O�N��N����w� �>�T�+�1��-cj�5�.�"h��G4t������{��A�Yg /�<����Ƶ��D|�]�pOV{���.-�, ��.���J�i�����{���|�X�]�)b����&t3�Je��D�]v.�TJ�|�y�k���{���j����6�O����L�T;��+A��8�wg[�9^��s�ϫ>Y����q�s�rˬ��]��#[��y���{��j�\�P�v|��1�ܔ=���^�,~j����T}�7��)2!�*�b���_�^������\��ܰr��J�M�C7����m\ʠ�\�ːdNB���t��S��I�q{�VE�{5�=:믠xzF>�ЈS.p�;{WY�&��Gu�E �(8mR/��oʄZ��kUp��T�W2�FS��4z��fv-n�x��Wf�ޠ�5��y8�[�ɹ&��p��o9a��w]�����Xͥ�<���\!#М"T0�,�}�	�����
*�nq�������5��#���7��c�:+x�ӆ��{o8]��C����H����4�r��j�lmu�{#/��'�~�D�����%�`0Ȧ<"��J��R:WL�j�;�v� �j*^�8P��
(�֤�!.N^�8��p��d�~@��?�H'�QJ�;�e�aS�pHi'���;십��g���;���}{�Yy�sʍ�ryG噺3=�3�z���5F��;����E��G�
��S��PZݷ5�q�D�3J�3�q/�{��gH�e -�&|�9��&�~�u�����)�a�0���tX�w=+,��z�����@.{xwAI�؀�����ID�o�;y�A�w�c��<�wx *���W!]�D�+{4��Z3FfvS����˾�Xr09�A8�)5�!��d�-V�;R!�/h�����&7�ez����%���>���W���R6&=��%��w[Y2�w�FF
^��%�ho��hQ�S��9�ݼ����m�r�mܟA-��w��	O�qq�+��y�㏹t�����O����c���8���� f�޻���n�)S�c$��ܳ��E���Lh\L�L�7��X�g�e���Q�~;��.Z����F�}{�4�S���QkB�t'ˊ�oA�y>�Z6Z�t�,��z:��NeҶ���t/��[\�ժ�9�c��f�E�"��{�^����ַLU���Y��A��g�m��4ZA�M=������� �jd��B��(�L�m�}�������Z>�~O�P�M���?KS5�u5H��WO����>4�Ƙ����3kb���۹S.���Z%��<K�Wd��^,�d���n��������b�2R3���I;f����,4L���o�A#	7��c��ۘ�<dk�yYl��:A0Z�2�ϕ���㌘���f;cL�����bg ���k,��ܵ���(b=0�ae�/�wQ��)7C�`�9+<�2�X"â�`=�&߼�}O�!���<����cx&`�؂��y"�]TT�U�R�2�Yl�6��g�w�`��.�� �,���`�X���(�[��n���Q��s7/TG\��v��v��0�3��&k�Q�:6֗j
ߓ���j��I�y�>"z\�O����/�]��Dp�;/ ���qv�}ہl��U�q�p8�kn-�ֱ��h`�Q�녓\����6әv�.4�|�#�qv&e9�Rf��2ە��	��1�J�\u=i�[�(B�d�i����n��Anoe��qM(�n�+(AtTqqCX��C-��>`^�w#�9 z{=3�Ɉ�S%��t�N�_���`�(_$�!f҇�컷ip@x�p5KŮ^�������R�p�i�z,�Bp���7}x�)ŏ�;s;��f��˕"M�Vk���R.��0���v.�b��O:��-c�f����J�*~��-��t�r���y�w�����Anh��EñFj�af*si�{J���9���vH����B1'�oh�Cs��%4^�O�M��ƨ$�����̋r1����&�<f\��A[��H��z�](]V��|>z��Q�	^^�6����姢��;.���U�gq�����2�l��Nb����"5Z��:�q^���s�@�=�.W���cc=����9;���Q.��wL�z��+�� �훾�b�z7�Ds%�$A�S#�Ec6��r����{i���P��>7^�����g[B	?We�v(���+�)Pj��e�V&�;��
1���/W�G�@���������X5x"��fr7��!�R�%�d�O/Y�����tǟ<�d!�A�lB�Q��M���܏�3t���ո����`6D�#�3Ⱦ~]�3g�l�=�6"�/�f�x�o�������1n��fgӣ��-��������a��)\)Ka�f�l�1C��Ow�����Ժ-���/{|�l�~�'W;[:���6��L.���k9�^-���ku!�=v;FoB�;��ft���1�e�4���2J���ļ(	&+��˿u9��5��=2U��Y V,9��f~*�&;2Wk�f��'�'��y-w+H����Rw�g
�k��suZ�#$���v~�3�½F���h��ae�[���P&�4w��[���ZnX�׺̀v�u�F3�n�R��&�aM�k5ڂ��f�E'��L�7*)�D�$�.���c�x���QK���En�xy+����h��x��������l���̊v(�qDluw�ٷ�p�ǽYU���5�Ddͅ5�Ē��p�Z��蔵V9;�wnT[7U����𶯡��t��gN���o�6W:���6�H"T�3���������V�%�{��ё����4-�5`!�=[�t�oP��T)=d8�nvi�IΝ���'��u�p	Ej8�SVs{�cW^|)�ǀ��@O
Z.\�� �ʽl��X�u�`�"�5+�U��8�,��u�|����ʹ��b���%DC��qG3��.E�x��VHb�����[��WO8����YC�s(��t�oV�Ew�V,��2k�L�'�f����C#����쫲)�^�{�'f�7;,�I2,X{���i�(d5y.^l�TѢ�I�A�m�9��
���t��R̳shO��I��{�6�K1����+���9QZ�Vg
�֗V�J=�3;\`�oDLj(���V�'N�(Q4I��UUUWJKUm@J�J����&����*��-Q���HJ�FY�h�s�f����+�"vIH�F��n�re�z�@�#H5�GA���h��B�rQU[���\E�W�-��F���f:#U׀����
�Ѩ^׉ʶų^c�� s�h�8�"�P5��5,A�k�G Ĭ�6�V��A��Gi�vۇ�]���s�pc8:�����Tm�#����,�y�FZ�b	1az�I���m*��[OR�r	��d��8^�bh/]d�8��5��a1 �5��r�R��lH�{2���k,rs��.��P�s�:���v*5�A��n�磈�`^Fk��y�Q،�f򆆮ٝ�Z�q<©F�n��qk�v�`�u��18�.���b`������M���j"Ů.��μb��M�45��V�v��F�5ĹG�]k{"p�v����g�W�DN#�wl+�8���s����빘w�WHp;Zm҇ :{d��5u��U���>�l�Bs�4�q��f�C%���hͻm31PKf�����\�,R�vQ`Kbl�t:4-!�1�� \=�n�a�.T��wMrfS\��۷a9�x�=T��4��ex�n�aM�����wUp�Fd�|U��N�!l)㱵��p`�\��Z�'\��՗[�R]��7�/,RAvw�6�z3t,]��u��wB� Dؚ�l86	v��c6�Q�])�s]n��k�6�o[ƭ�GI �!�1���Ⱥ�>��u.��q�����j:�]x��� ��`К7W,���T��c�	
	�@]�XCa��6$��ŽaHMe���UXmu�i]��L��!
6ʩ.�Y�n��m�k��\u�	Vnm�:Iɶ�긫]���殓\�m���um�Rul�.)w���l���%�=s�%�����c���3;Z<�V,۬vr=��k5�ͭ�z��WY^�o!��nӲ�7ԑ����z�oz� 5V���9.�W�<#{�:)�H6 wu+�_a.dnmx�>�<��**Y�̾�JM����I�#l��H薋nl���v�+��X7T)K��6Å�H��a1�\#�'tl3O���GW_��E8�q�����5 ɍ&!�V��s�:8%�O�{8�ޱo�퀗6\IA�J��u�	>��m���l�0������Q�^�:�D"~��t����o^�!"��'\Okחb(y0�.$*�f��u��Y�O6a2M�*� �Ɋ���6�oֵb��`��U��a�A�Fvy�QU�4#B�W��ʛ�B+!rc��kJ�]^9e^��j�`��ڥ�O�J��s!xx��6M	<��<�Hc9yv�zn�e9��q�ކX�r8g�to��1�ɖ4A]��pbȀ�Դp���]x�@�8+s�\I��e�^+T�ݳ�SiAm�!;�zw���ed{����p��ӫO2�D�rUj2]]0���mcV"K~Ŗ+��V1�̸�&_@9=7s��掘S�nة����g��q���ʱ+p�.�KI���ya!����\�o w��$n<�g��]���r�>�|f2
E-|���!��_hw��Ĉ�C��m��2`@��Ĥ[G����	���fK��5��n�CWD�e���PU�{5Q��f�Q|@{~Y�X�*Ig�Q�"FI:g���̳W��e�5wk!<��w��U�*U: $`^LU`�
&���0��/�g�3A=�@�b����mȅ���s����6svDw+�T�R�;3i]^�p�G_ޒ4�.�
tk{=����|w+33d�}�U��Y�嗫xZ�c��u^�R�׎��|�8�j(�r�^6y���Y�sxm�ފμ�{ٮn����U{�p��(��	i�����z�vC�ۑ�<W<P�+՝�v0v{�K�;��6��꣎
�n[��^��y�	6�ފ�/�ǁ�ܝ�	���^đ���tN�xe��e���_��$s��
v����w��Gu^e\�yR_[PE8�X|�0�OԽwU�j�cO��m�&�X��w��u�he�$m��f�K�.���#��n] =��e/RL���{~���B�R�e�m����������n+�7mz�]-\������-�n����p[�߭>5��ͽ���P�0'G7ƶ�ᩮ���I F�k�&N"��1av,�Pz8�ut:�Z���t�т��L�ψ���l�0j����[������L9W��"��	.6�f6;Txx��}�^�}�w��Xkb���+�p{n�8Z�c�+��7F�M��&<���I�;��t��^�Y��Gno�!U�N�f��vyr���Oy�!hmȰ�Wpㅱ��Tu_���N��&���D����S%��/{(� ��/ɞDݖ��f�nā:�.9V���v���z��Q���/�E���0\�����۽���(@n �SS��N��Ⰸ�z���%
4 ����+�<M�1Sq`y~�}���=L�]'`���h��-=�7���U^Ӯ�ƛ�WQ����"�7KoH���w�,b��$�����G�V����}\���R |ϲ����خb_ɾ�n����\u���.E2GL�G¹oG&�0�F�X���V�����9��Ɣ.}�n.��<ـR�'�y;�R�ٌ}��K�uT�V�گS|��B�:V!�s����>|�{��ӳf6���g��K��t��c9���P�'�(��6,X�ySIsxx���Z�{���w������Z.8������pss�	s��Ã-�^�����h4�1�B����������p��9��(�5��>�-O�Xˤ=�
�Y^�y�e`����l/,좛�	�u�=�>��� e���������^��3H!W�\/��~�Dw��� �s�qW$�¹k��su�b�U�~�,�,�3i�alv�狀n��u�B2p>n=+�&N*��El�	L:*%���T�L�2��{۟���.�n3ګm�����*�J��ԧ��2���ۛ43�,��>'<R٬t+����0	)2��"�}/f����`b���O]S��z`v�H��3�A��yu,FF/��XFVP(��\o#��5�����V�G;k6�Κ+��N�-T�^ѩ�P�A&�Y�w��K7|�������a�n�WV�^�)�BCxBL�aFH��w����nn�]��c��lt]u�T��y:��i�tsn���l((0nB�L�Օ�Ͳ���{hfQ��cn��1�۞{=���jg��+�A}�ǍV4�cp]axu4�BVvÍl5%lq1^�D�68C�uf��`��lbi�����̱f[S:��<9��F�-Hkx��r�Ў�;�ے�{��-���L�M�t��� �M�1%F������%MBA;�o�RK��';{N�P�����s��(7�Tග��jdvu��F��;PMT�Y$(���,z2ri�Q�A\q���<O����q+�W�^�6�Y��T3��{;�I�'Bp�.�&!0�	G$����&#�莟
�;���K@���{te{O��k��6�t;���';)�K�4�a�$�f�4�f9���y�����XU�����}���vZ �� tXW=w:9������jB�%������4���3*|GC'ﺶ��ف��a�N\�:N�f�ׄLV�>	F�к����#E��h�����bR,��7:��f�=�+7xn7��[�w���|)F��|k5��|iܝ.�e\��V���|�1�]�0��tv��.�`����������{�+s���Rh0`Ä�	���э�Ɋ��i�����z��f�� .�kr��D���$$T�����㟎0�υM�G��\g��4H����������8���m������X n��s�'gfn�J�������hSd�ه=,�!-!����V+w��?*[������ިa�b���2<n���3��z�������x�I!�yS�-%��Xe�7���V	޻�ˎƾ t�s�"�z�8rԥ��|g�;P��{L��i�z:m��I72��t�ʌM_�Ө9P�j)�w|~��D����b�k�vDU��˺�\��nv��g\�)��8d,�L-G�<���c��Gr���ި��c~�o�OeA;̯Alp�F�5{�a>0Ȫ郦S�܂�X������L�[`Tt��S�s����wZTs�3�S��71$��z�NG��(s�4=�����=��v��)�b��/��nG�딿�U9=2�F.�q�;�S	��M��.��ao�oƆ�O޼�}x/xRWd�z�g�J��5�#/���H��G��s���p�������c�^[��f�V��z^㘥<�=ڪ&�}wl�ǡ1�
'j&ك�=8s|2��^�j������s��>�PAf	PR��=�lՠM�{���/��s*yQ��}5�*
 !����#��%�A�Y@]�!�)���NF�K��U��&�}�
��g��w�V���G��_95B0��/�5�1�P��n�þ��Z��(��Z)����w��pP�6�$�������R��M띘�������d�h|���������탁)-�Omq=N5z���֛��Q�%&����aȳە�j��\m�Ѧ`�m�Jwܷ���2D�k����M*�Y�l���m��J�$`g��>ŗ�����4�w<�d�F��R�l,��
�j�Tѫ�!�������f�v�m���}_
7�&���=�'� ����R^��<���#o8֏w���G�]9>���*}��tRY����[��G�O�Wg�Eڭ�$3���M��w�#k��Ɔc!"�ęʠ}ط��P�%�V]k#2:�:�����)vڷtUm�ͻ���E�T:Η��ə�s�VI���8bU@By	��i'�a�灥5-
d��W��5�-؁A\=7NYK"���5�o�l�IZunv����Ɋ�B�/Uk������;�F�߈��k��3x��ٽ�V0�}K����ث=ཡ��H(ʅ�@��qd��`�v'!MϲWD��F�ڶ �1�J�Z�6<�(�"�]���L_�4�Gv���JI:3���+���츛��Ȗ�2
�y5���<�fnf��n`��"m>���װ����55+e�E5�	�&g�!�d_n�[c��][\�,p��!4���͞���ۧ�/\�4�i��D��c�ǡ�P���o�y������+K��ֽwc�����qݙ�ew�I8h��iì��ڽpT-�V�67ǚ����͌m�^άIB:�i;�3v΍S���^sK=>���	.g��z�P\V��mC�P����oB<���a�	�:~����+)܏���W:��W�A�d0k�K��)c�5�z�f�֛A�ͥ��R���.�)�_����{�k����C�d`UG u��2�%w���a٨6l~����.0c|K�{%�:��/ٙ!��,�a9X�hS����w�w�9٭ BZ�0�ƻ7P� �S�[�+ܦz2��:��zJ��o{(&��Q<�E5�R��@葧^l�Q�����Ӟ3�l��Oo��K(�d���[Mv��=F�����y��bp�q3u���l�>���e��{I�K��Ƚ��<U}s�57��"����S=�y�����ﷸ�:��V����ʻ�	x�h�@'����.�m�;j�^�`��Q��x$��&S!�r@D��!m9)�cŜ\2�-��8 �*L���?IJB`p�s��0�֑CW�Ĝ;�K�Y����)�U��˦��s��3z�V��ۯ/5U����Ff2�.�Z�ȷtc58�j�e���hdo�wb϶�vY��D��ϖ�@y_Kk�AW�B���D)��{S��a������?j���WC0�,��&�<<n�k)+<���m�>���q�,���j���C(�c��"7�ׅ�`{��~�\'����\K�'=J��	�+��f��f=�tqL6�L�p'�֛2ק޷��R�~�/��A�ۻ���J�K�0*'�����"�N�*I.���h~]�U����a���b�l��D��6(��cv���f�*�B��~�_U��J�V�8��J�e���0�hB��&�B���,�w3v��tp�8�˚���EͰE��C�X�6&�*��fARmf�҈�l�N)��h��&k��l�Jmw�1�3�rz��͚�xY���1���..��P%bm�Qm��[n�C�q�͗:���,L[x��l�3(Q�^2k�Cri�s��c���j��:��v؀@I�q�	����uq5s���nÊ+����)�[�S�&�4�#�|�pCju��C��������N��ںZ�������,���JO)Xhwޟ�o:Gf�rqG����I󮥷^K�����y�ٶ*�z69���1��j��w�1����^t�Z��0{_��C!B�
4ɋ��A�����!�*��E��$�6�H8I$��Q���ڮ�p>���$8(�e!�h�Xx{w�kh��C���sR%���	ٝ�!�ٛ�j��ˆI$�5'�����������)�]C*�"��sm��>���ۅ�h=}��P��߲3�|�ي������4Ԣ �%��Z.����]�ǒ�h�H�Tnc%��6�v5�O�����Km���2�Ч35<��?y;�<�4��zjxe�/��|M-�<�ڙ�}{�\�!޽��&=8�`/���+�}lHӱ�t��g4�	��h�L���QQ�H�0L%7N~^��x\i28mb���.��/^��<���=y�5v\��A�������+/�r�����Gf���Vj�vT���rw<z� �Y�sܶ�eϰ;����Y����Ϭ����]M�ۘ�v�>*� E���	{��RbSrXͷ��'�ztlN�@��5"�{���,<��Cr=$W�{/�{ٺS�1޻ׅ�V=�]]�+|�'��6�EԸ��oz�dg���mu��7^C`�������}6Y��%D�h2dn)�h��!GМ*6N��n���`���L`�^��ޞ�\��Z�,�H�MEV������:��/U�7!�=݆�'@~���7�%�tҌV�t�Lv_�A}�H��6 �Qzŏo�<2�;�ܕ��8�j�;,��=s02�E|.T�r�љ=�X�u��9��R�A��ۉ���w'����N���P��.M��t��#��ML���-s��1���v^ʀ��:�Ӊ�3wz�Sa��.XiUѾ�Td���§{�75pe��>Q���F큓͈�3�W"�w8r���nv�'����v:��{�X���${s�;�](�8v�x{�ŷъ�G�=��O�z}�Q��2𬶺��*�w��C3�(�St(�x�v�pEӂ�Y�SD]3V.q-�[#W/]gLXђJ�:�<����Y�Kx��R��|&�6�y��h���2�����L@4���=�5�����ow.PQ@�A�`7֭oC�2*^fU�gص#j�-���|矗��ʑ-%�!�&]8�9�nMOn�)$P�pa��E�1�g����������C�ٱ&�`f{�4�'����,�Ȯ��
{����T�-�+-�~�uUi'>�t�6v�>�qgZ����B��n7�u��X�E�GW`�y�T�&M�Y�y��v�=��/��\"ʆ�u�R #/3+�����hN�;Ղf��vx]7F�*��ټ�G�_%��&�\�+��@�o����#��Ր�����o�*o`OW|�,�O�� �)��n���X/P�!����;�%�C�61���&���rY�5���@X&�i@���Ճ{�ك_�5�M:f:�����s��'�m��P_W���b���L��g��MC��P�1;q��(�5�1�ِ�}�5����y)�榹B���ԏN��\��`��>�7#��aște�"Q@-�j�_��f�+MO3�����k7<;�11�v&�E����L�R�!�x� ׷|:d�Ș�v�E�ͫd�+��ss��*�R�������6ې�>�1wܢ&��ܬ�oݎ�*}ǭs3����%s����<6��RrqWc�æ�v�E�.�Уtd�Q��=�0���>->^
�����c�x�����d*��֡.b��3���%.KQk*�5Ǝn��8Y���)�Ѻ����yN\�T(R�(1��Mi�_kR�N`Y/�܌O������"��A^�#��=c;3��e,� _"�5�f��k��&�2D���֫���g'"������,?�¬��Dg��mۏ�Hy��'+%X��*ۍׇ$-Ut�1��6�ʷ;�rPY�c	v��v�o���[䲨�
`�8eSԂ� Y�B5	z�ve���R�����"^��ê�����2�)�"qV��岂^�b�&aq���7Q ,�]>��]��gnհa���P�9�c��`����T�ڷ���:�!ui~�lm�o���t(yjoΒ�
+�s�;wYR�m\7w�M�=0�_�h��P�2Jk �ӗJ�\=P�9l��ff�ʁ�n*��&��a�sx�Lp�d�L��90�%�2qv��	)Xb����A'��sL���:N�S$4��k`�@��W���k�X�iuem���
�/1��c;G2�>�:±i��\ �������⬂�nH�9[1�s0�tS�Xrr����mq�^�^�+-�c�SA�MV3q��
Hn-��l����#�!��?I���j����4�=T�S��s���Rf_U���,���yc42S���U�4�ͼs�xX�܇�^m�
�@+u�E�p�)��L���乫靋�4XF��+�W�Mq�ts�Hk�K�f
��mC��R�f2�@m����kv\�ȷ'7;�jj�j�=1�Sٸ0��=Z
EPwwkX��8�����;�A֢��V�g�{�X����V�	n�a�t��e��s�v
4��?��R�W~�Ne��Syەͱ����s�Q�,lι��&��«_�P�]p���N����˧&���{��w�D��-v��^��g|j1V\�&6Nj�������C�O�Fh8�ʥ��t(�ޗ�����B�S�uz�+0tPm��)��y�u�Υ�YUHŨ�#2ܮ�����z6�h�Ͻ�pj)V?)cI��y�mZ����C�9+�j�8zs��߳7��H^�8�30l�F�<h�\ଝ�DZ�%硁�呧��\p�#�G��!�.��v�g��-���t|T�-'�زѯ_3�c>���{��֯t�F����c&�p�t�ە����6�'�;�͘�#�8'�ϔ�g0F�^�SmX)36�%��k]�gZK�!���~"eN�g�o~��Â�s��t�c��Y����8��\�yva]_-Oq�g�b�z=J��z6;`��5	�]_=�g�Z��շOڈ�>���t�{�}F:��Six�j|"�VPk�sX��[��_�Wџ_��@��28�f^��}��� �J`���4�F޻�b����c�����L�1�n�ۍu�X�W8��֮ �x��s��E5���8���Ǥߘ���߮��f�|��1��װ�D�5r�]�oM�l��x,�4�Z{��,m���<�H��*;���R�ܠ6��|E�yR�Gb�QQ9M�e�ۡ�m��ݮ(f�W0C]�K}AuM�r_dΥ�ݖ ̡�ă��6(u�yY6-]���p6�;u���N�f��l˃l�Ti�l��"V�!n�Hc$�C$ ڠ�@��Z�[��!2��fp{B�g8{,�s��$&C���\��LD�Gr݃f���5��0��6.[c���J�J/:�=�cc��V���Cd�5�;e!�&��M�3�HM�`�΍ƚ� hq��v�4�^��5�c�����NQ6(ݲw������78=�=l�{^`O8 �{${��r�{���pJ������1LV�˞� ����-`�Y~5��{;l���t�"k�y�p��ʄmE�fn�������	x��z:�Nl�&J���Y���ن���FT��3��'۹Lx��H�л�X+ץy��	L7�P�v:���P#7��!a�qU�$��;s�k][z��~;�����̡�x#�O����h�YѼ��nmƪ���-L×�����K�H����uL���#~��e��_P*tӟ���V���D<3�L���Vg��xH'�=�Lz�nsOa��_�wo�m�x(�n�ً�t:B�:|��ZÈ�^Nd�1.s�|r`��~�n��3�j�|n��4z��G����W'�6B��Q���8�=9o�"�/G���OEظ݆u�`����'�G�4�	U��5�*�˝�!�a)��2M�����O8��V�{}��x5:�Y�&�����̂iQ�!������ݬ4�;e|��c�;���q)��x�F��h�)S�kp�k��3*^���,{}�����N{~F3�O%�U�ۗwCN7-D�v�E�S�ۅy�]�^·BvZ��df��n���'�b[e��vLLT�G{�MC1��#uٕ�ys��
��,JTǙ�N'P詤b���i.�ĩ*���穜l.g�oDl���=�)+|q��F��v���zq���{��V�����ߎ�7l�#�8�#��mI���\��f�a��)$�m%2 ����j���s��c�^�~�Ni_�.��OVMJ��}�N+<�	�'G�;g5���y<���ډn�(8RF{:/�	bRݽ������oO{���]Ise:>�
1l�]N�s��LN��ݔ{�f�-�&���q�2T��a��ý%�,��sW�=��}�M���r�c?dH�G���������Mp>��"*E��8����&,d�^�&�k�Fӯ����a�A�ؾ�j��e������K��$�����L�{7Ç���ţ�qw/�.y�g[O�  ��^�b����	�]t��Q�j������JS)4qm����w|;R�YD4-4�in\��+���dc�
J�]���1ix�![yʮ8	��xV�IwV'�=�m�#��g:@�{]��Jm�U���&��&�{:��΂�!��@��G>�a�����}�h��s<��hM0E�a1�\D�#��AxBd^�9N�[$ֶz��Ξ�g�����q�+��U� A���㊜owm�j2F���c{-z�|�gzx{s�{��(�}��A�u��O82�8��XNPȦ��>�8s.���q�\eb-_"2�7�\JoWu>zq�7���L<2uLR�uW�3pW5����Ԑ���1D�Ɓ|��Em�:�/0A*\�=��\W�)`%��Q�����|�okb�݂teq��[�Q��E.�L��^�J���F(h6`����k�4)��zwsn��g�{L��>m=#�'c5�7uR>>z/&��8�;��������:E��/Q�g��U$�/��"1xػ;s���Q��Ls �b	e�(�'���۬x�=���*&;�=�%{}*�F���r�%/n�R){Ω�;�(j"eix��*�Y��#��j�.��>1*�-2�a�ia7�T>��,w)����8	'Wnf���;3��3<����6j��C7]�LM�\���sߥ�%�{��!��اy���{�x�R�W�gw�`0i����p�a�-����ɕ-�ce�v4Ü���U���o����~�������늳����Ʈq=�=5���M�D"� ���|�I�6����.q��I<�����Q��Xo��������V�ʸ�\;�yP\+|�t�frW�Z���p�N1�5��g3��q��j��BB�g]C�kTr��}]z|����S��^��oH�i{��Z�Y��Ի��6ٓ�cݙ�>� {�H�&2�qaqQ��4���2��Þ���}�.�&���/餠剁$�"Ӗ������#F^�]��5��\�n'�7Q��K����B�fq��v#Y�t-��3|��P Z����g��/�*����e�Z����!����ϟ
�9六��*w:��H�P��>�;>�'ٺ��w���ݓ�FOwj�݌Q~v�r1�7��#��
����lܝ.�{T��:WwWia1n�0)�'�q�0���E�`�Gf<�rЂP�aޤ��ss�j��&ۨ�E�v�� |=���<�2�`}ヿ~���'x*̀6|�:�kW���.V"�}X�4f���R@��6v^�W�ng�;�
��A�T�y�ƨ)�6Hp��)����
�����4�㐗)��d�1�Fs=�;G�O��5����꞉<r��kv���D��稑թG���vg�ݽ�Q�0i�����*x�RUlՓ��,�M=;�������ٮ̺���A�ľ��֍�5L�����n��k�tda1K���v�|�����
S�ך�w�id�8Uv�<�u�(�rB���3�m��*ƚ}�;
��/�p-�.���rj1,�j.|����a]Ae��^�Þs�A�߯8uݱ7��6�9C�FmV�-�s)�yݹ&�sy��&�L�����R�{!�[��X�3De�b$=����޸��ҽ���F�^��$1�9����6���ps;��2���Ok����n�g7�4��tV�8���=��bWMˋx�8���·�LګT��<�E솨=Q36�B��w2���8��J�u�ġ�A�M-���,��q�=�,�od6����gU��kù"e;`+���{��L:,���r�k0n%a��i�؆-݂h��0
P��t�l�@�-���f<�!�ۮ�usd�A�G�mc��͈PY����-eM�-ݰ���J��K��fٗ�,zFGr���Ԭ��;
N��7��Ƨ���Q��*k�do�r�SI�I.3A�Mca�~��
|/!o>Ύm{�=v�)���+����6Y��5�����Ǯ�|�{��>�vC,13��-INd�D��TZ��n�-_��-w��e8M'��Q�;���#w�A�8�)��_��^c��a��S�<FD����D��I�aH�ɸ��������@H�`����
H�	�:�8��<q Y�^���_c��.�*�k*�Yھ�´_�s,l�z�y��-�}���2�B�E���
�l�Y��_Q�&���O�:��k85�|;��K]�q%��gH� �A�۬ϥc9��g�3��'J�!$A�Ai�-7
����^z�ί���{,Mta�]��eM0�����O��3s��-��A�-�O�K�ǎ-��o��`�q��A�g~��Y�M���ݪ��*�/@9<n�IbU>fw^I��y�OG��\�mNKy!����UO?�{�o#�j�K�yeE����HÄJa�,W���>W�޽a�^⬧�g�x�~����0z��>A�:1��$�<�G���gL<�g���Ƞq.�]}�&�kM��:�髩u-���h��8!�:�����:�f��}˛��+���c���Ď�[8;d�1����:A�y�2�xF�?�D�P��JC0v�F
m��(�ț<-�pRw��u�uAP#��W8V���f�	ɀq�����Y��76���n��Ӹ��Nj��n-"�n6n���>˞�Կ�l=9��z,���˴e�up���4%�1c�ŏ+0yZ!$�cX.�^Ttg{�Ĥ$��,U�G�n�'=<n�=GI;���J�a�Z:&7��>JҔ�1J���,�Xэ,;����d �����潧�\�)�)�c��w���v8r��BwcFHX���wҺIg��+m��ܓV��dRw�"��T���v��^�<US���ҏG}�.z�75���i.) "=�E6Y�m��9����U�����W������t�iȑ�H֦x�E�;�I���y�-��ڍ	�dM<S�SkϪ�OoD�Pd��&O���`|+I����7�c�yر�͵���*��J�B`gn��ǌ�F����d5�؛ӟdgK+�>�#k�g<�۪:�T�J��+{�d��i�TF� �M�i(�:1vmn:���>P8Wg���ￗ��߱;Z�B;�z�����\�l�v����t�pj�.k���߽�_g�����bwTO���vw1-���%|����I��A��X����N�C���i���D]e2���?Y��,�W'm�S���Cd?�7H�*Lxn���a%�S�#k�n��]�^�.��^8Gt'�i��-��� �T��_>��}�z{B�:TG[�+jf�+No@U��ڃ��wׯ2����]G��ZO�m��gEm�B�5�`{�.�1gQ�q4�
����s+2�^���\�r�As�|���^WMZ�D�>�����L!��G��wQ��7�es��1�����������ٓ7bCф#���sdޞɍ��*�u��1��v�>;�����t9w�ڸz`�~����gD��o�x��6��he[�`xx��F]�Qǽ�f߻`j`��l�a��d(��8Ce}>U�%/7�e�r?0+G���=�����OA���Ff:B�4z@��ǳ���{�ˉ��D}��qP�k�bD�v�tO�A!�{�y��;����v�$:˖R�д��[h:�������A���e��l�%�y
�{՘�L�I�����C]k�ͪ��ߏ(˳*�����1���+��>Zg;���zxL�Z����{}�sc�,�����#�\��@�*^�o��bU�r�p�V�ۃ���x�?W8�L�{��a����ؗj�����R�yq�M�%u�g���9��7���!�A4�L���3�;<�n�4 ���Ӎ�Bf+ܢ�wHhj�.Ӥ��P,hZ5Ö]�I�ZA-t��]II�s��0��$8�}����z���������R���I�R�mt��{G@�������J�P�Y\�:�ȱ��K�6�l.^��b�c�S^��SMY�t/��'��]�'�ٲ�߄�;��-���M�KSX�xk5��򚉸_��e���3�xm��f���2� �Foը�얍nk��׸��0:�U��lPŮj���8�<�;L��2�bM��2�6EN9�Y���*��0�#n�q�J���t���L"�iڶ�:����9��z���D���;v4�H�f����6S��D�Q��h,�i��m�P5f���&!1"_FJ`�N;�����J,\H;Jp�7�vy]��16��q��d�i�����ӵ��u̎�m���`��e�X6��QKChT����#훷�7��LyW��`"7�];9I�g�؝>[�d�*`-�}OR��u$ч�wT�j_g�PI�-d>V�G]����KARꝲBc7b�#����wޜ=Ұv�60c蕗�и*����pGg:�ͩ���5��Z�הv���w�Y�H�lG9c��r���ɋ2����H,k_}9y��[2
3�ʬ�@��ym�,��X��ί��#��딘�+��ږ����*��g-\�7y����n+�7K�f�������I$�H��T�!���c��ÝF]���U��%1(;]�R�L3qk�t�*�Z�4n3����g�D��O5:�6�t��p)6��,���\���b�u���XZ��K�l��d�y�i`;.Ʀ�"#���66����%�&�HX�૫��s��,7#�8jҪ�k�'`T�鳢�D%e�1v���@�lLm;t][��M�N6BF�ɸ|5y�|b�=�yO�u�63���nc��K�W����_k9׳��Ҍ�p�-K��˝�+;f���#�ֵ	�t�zȻ�.y�wd#Z�k���R޳u�,�~j��z��rግ�9���W+��Y<��wm���1����Xp��c���B����o��:�VPɔ��n��˲�`lP�^�q� gͻ.�%�l��ZR�v �b ���5�-��r"��G�'��j�|H�c*��}��ڀ�2���x��\S�!g�sSC/�$��"H6�h���wI�*�L�߽�����D+g_v|�'��'��e�9@�M�c�f}V1�X���r�׻��d$q�]��4��]���\�i4D2_��~�C�g���ӷV��J҇Foy�X<ډ2Fo��{�
�g�m�n��Z���@w����x8�ˬ]��#��mp����1s�h~%�$2A��߷�e���k{Z���1+��r���-�+���|m.O��E������Oi�{P�t*��aS|�SnT-T����HM��t��ջ�ڣ.أh򓜠`$!�{�zr}1�F�So�q���}k�Zw4�/罏��SfUy��etٻ��ɪ�B��W$�˴�0��X����g�tI�6��!�b�G�x7�x_j�f�Y��	���2�,�v\�-LY���Õ���7�:=B���UWε�+C��5ա�jU��
�(���uM�˕�@:퇺�v�A�b%�s�ъ�N���#�gr�汤kx��	��C%Lշ�u7iVՄ��v�V.�l����[���C+�X).��{D��Uh���j����g5ջg]M�GA4��0ν�ٸ�CA����HHخ@G]a�DZ����v�QT�R���b�S�\�b*\5X�,7f�+i��9� C��J�q�����T`�;l^.e�v:�v�mk�n�vi����R^�9�/�M�ᙫ�B�nT�|��y��#yuy�e���nT�l:����na.����i�g.��8y�$�	�rj`�P�iC);R���H�1\��ׅcz�&$��s&9R�-�ټ(�|rĮ�:���;\*ˮ�4���H�c��tzsnecr���x(fܺS{���Ԩ:R��sx�7�5t��U�M����6�k���{+������;�FA�/��YI5p�O*�v�g�ŗ����xos�V�� v��t&Wp��.7Y�^vK4>i��])�s��07��+{p�;�g:��Y����s:(>������g��cw�o��V�$�����dDuXZ�j����ej�t*�Ç6G�f����u�A�[�/����5 Z몥Z�V�U���
x����e��T
��
U�m�yM��mU�`�ւ�O���۬�r�I��G\.搹z��%4��E��s��k�e
%�Bs����a�쥻z�:&�@Y����͵;+/6�H�.3�����كq�롋��\vݮ�v�'%�:pA��Z�>�j��9�-sҔ�7lvtU�{]qk�yӦY�jҥ��c�D�����D����vMI�V%ؼa��hU�0J[�X��ͦ�/A�PBSڳ/93�u*9��^��f���c�	]J�͚���'U�st� ��=s�wb�!-��a�#KY��Д ����6f0a���5����m�A���ڢ�ccD��g��cy�Fz��B���sS��&J�F�<{�
��x���.1��7%q��&2�7mo�W|�G:.;�L��f9C�+q�C���e����d��A5�lQpn�6Ɓ	�Jغ�p�(˓ �ۭ�#+Aȝ�Iitθ�-����u�3Nv1��m��j���Y����l3��9�ٵ�;+'%�M���ՙ����q�s�c����^�vt���v`��f(��5��-p0�@�hNlA�.ޤ���:[�����WA������У���r�(��unZ�ρ��70��$0�ݻ[��t��aHZY	vq��Ka��[w2��c�2�lojF��Q%�ˉn��,].�6.a8ݭ�:�� �:�ƍ�T��V*�.��b��h�t"�#k-�-v7Ey������ytv0W�+l�q.����f�e����aUP�XL]&�-��@�j���u�b�����pu�bjR%���.�i���v�����펕v��3����IY\�Yc3M��Iu\Ȫ��܃�8�&q���:�u�\T�"���|�_�ɏ�v� �k�v�Ѹ��u)�O�޶E����c��v֒d���Zgi��y9;������Z����ێ��u��pskY�x5pE�ڱ�[ssI��#ZlJJ�Vi�l�CB
N����7+�Yzng�EO*V ��룔��tBG����JM��ؚJK�~�B�]E6V������.$o���_����B�;'c��kk��ݜ9�k��D��1��fnD&�4چ� t�G=��T{��� ��3Ǖ�7�M)����`�#�q�R31੆y�]_D�n�2�iB0؁��M�TVh����	��Ҹߏ����]iB����`b!��C�Xr��q�C�J{�Ҧ�o�)@����C��Vn��ލ;	��p�E��F��f�!�;�G�}&�Ё���=�<�å�AF���?��L������bz�js�A���(�d����9&Ϧ]���׬"�m�A_P3��xna�5��gis�Ǖ�5b2n�F{.T�=��Չ��__���do��T�.U��De���
���!����Ci��tH���W\e�~��{Ƨ�"}ܻ�ļn����G�.X�9�e1g�*|	S����87ݪ^��72����w}���Ġ�� 6D���\p>8����Η1+��F�� �O\.o[R��-T��0űh:��n�ņ9�k;��O18
EO�{���}&�'%�7<������[��H��.ro�'I�6��}}����3�6������b���Ķ�l�<܈S*���sl{fV�U���R���z���1D@7wI���'8�2�pF�7��3I��L�O�T��a��@�p�RCP-P�9����FD j��Z~U��s{���M������K�ڋ?L�{�8M���G=Ⱥ�M�� ��9��ѼY-�h�D]�x��g�2�}��O�3M�D=�z=TO� Ta�f���๚���d��B|�4I������V���8*';��p�_����vn�pp`��N�`��|���y�.��f��V?J��f?g+�;��΁��#�e��D
v�B�Vm�x�>]f��F�N����/�Ϸ������Gf@�iÂ���!L�%��@Z�^=:m��v����:Z7�;�C�`3 ��n^nq���L�ֶQ��xߺ�Um�A�%ǈ^��o���{���Q�����7�R�w[hNݷ�笨py�t��n�nw~�}[���MLp[�-�G\�b�*�R%5�V�-ۻTo0H!�p��� �4��n���:>�3��=b]�H޴-���Ye��vX�f�6+�!Bt��p��Y��6�e��
m�ÄAN�7о2tA�fk�{��xU����5�(�ƾ��9�+�3���{kEb#����K�Ωf�������g��u�8m��L J�� Ƕ�$k^}�iЃYҞ��A���eh�m>�w� )'����%g`�/+1ډ>�hṸ���wpcI�|?u�z?
wB���8i7��޳��/���>��Y��3z��|�]��\�Y��|}f/#l��p��������T�M̻��C�����e�#�cF�ϐ�y�KE��{���h͈�G%t/n�{2�|X��gNV�s�={=�jha�|] ��0~�%�g��_��$���8�E���A�r�O���ʭ��r���}��t�	���4�+����D˞�9ܸ�H�50֚Otz�>{XF�f۱��5!T��컧�e�s0��� O�������s��Z���rpGn��v�XvP<� 0�! �,.^�s�8�<��r֚�[�E��fu�R�{eғ��o��{�%۝t����������Ռ�~ûqjI�$|'n������ˍ/gÕ�r�V]x�z����D��$���ЬA��r��S�ext�Aѭ�7vG���]����������o�	б7�4�달����,+�L�N��Gʀ�Mb��g0qz�.8�W��ͷ��o/��=�81(���U\�R�|���]���Et��i9\�hpc�<^^}�����ˋ�˴=��@���3A(�VZ�+����2��4:�o��}�n����5O���1����W�ɵ�N���3E.�ɹ�o�y� h��ۋ+�f�Ӆ~�+�-Lb��W_����}i%����N���vU��5T����͝ø���v�xw��kOcpk���V�X�ہcs��m�8먔Ɩm��e�G�[.��CDM�m�� ��;Ec�p�물R�����v�`��Z�ۓc2ҩ�3:�vn��H�n�kLK�v�iE�4��]b�n��v����/R��	� b:Z&r�m��lƫ:�o^��^��� �Ku,pR]�"��Ǝ,D���^��tY}�d����=�>���^0����7LN�X��W6[B	�c7g���=�G�7O��ny�<fn��U�9u����l���d��N�׀��a�=����ޘh��=�"ƒh�[����Į�5.$a2���U���G�o-�Ή����x�� �\~w+��c'WD<�5u�|�Ȁ�V:�[p������_1��3��wwz��-r�}�齰�]�+�KOٸ����e�8׏�Mfжh<�;�MR�h�{B(8LhF��l�;���2���TWR�}���|�z��z�/F;f����^7�m�ʸ�yh��c�ל�$��7�v:�U>��%u���Re��������E]���5�~c9��8gX��("�}2|�yW������M�Þ~1�%`�y�jz�Y�^�iO���(rj��By�*ow�q`��i�[V@��U�WO	���мF�$���zmx�>�����	ئ�;�.�u����#��|�g$���[FN�#ٵ˽Ingp��mQ-���d,�(���_�I�hW1��'=�8W�q��wF�I�LƟ$2���W)h�uLǡ��%y��k�˫���^[tN1�_
Pw�b��}u��3-��ˮrZikR����ತ`�nryW�y�K�+�9[Æ���e�LT�ؐsG�K�����ŋ�[�Im\��"� �f��r����5����G�]vt�ˢ���@� v�%�.e��B�W��:�z0���:�)�v��"/x��h^|�s,��f ���F�1N)���k4)����Ԓ`�%�e����Hh�;bF��;������*����i�h�pi�5Η\t
��F�JM��q�ؠ�rx�g��g����Utk�ϼ0Ҩ��������~<�p�l܌��o�p��y�{Dx�
}[���gx�ob��f���c�pj�[((��7��}�<m�
�B8���Mؓ٪�xB:=�`p��MKٿ[z��R3��P�Wʤ(��S=>��Î4>�*�(9���=O(��_ċ*�VoW�-.Mo�C/q�����k�HV�]/,Wo��׷��o�tܰv�_���{N6����kmS�{%0weՃ\<#%����_ۗj��묥�j���oB�,�<�A����
Z0��1D����[o�v(�W��ً�޿��_���n�p!����p�����=u��W��.�WQ�KLת;h�`���ն{==}�LWi�h�c�o�b��g��7�w{�n���j�t}�}֝Û�%+a�]�.� �7��@�څa\yJ-[��f\	s�	y��q+�nK�Ǳ�aέ�*o>��q�c�u���M��&��ё�ɖp�	��+��R���v&9�x��y�Q'a���t㘨� !���L����=�o3�vl�3~.s;N�N�-�ܔ!Y�w���C{#b0� ��\*����9Yy3]���<􆤇T�����M��Mr�s���{���a�p��j���o�ԌM�{N�U�g[�X���M�x ��h�эiI�p��"��J�sr�p�l�"d%�ޚ�䗍(?{P���Y�8l{)F���40-��P*��H��Q�RXj��ܺ=;x��(�Qv��w��G��{�\��{���q=�M���o���!w��*v�ln��$,��#7Ʋɮ�]{�ښ�zA�~�s�4{Gr~�扭KT�����5O��袯5��f��n����zo��o���K�kQ�
1A"�K,� �XM�gh$A����qL<�A�c��n;��~�{���-���U7��Ƙ�z��s���M��ZfA�P��[�A�����y��'F���H�1��/�b�^xꗤ6�[Z<����a��v�q/gY�r��|���*ΪT ]K���3�UE���\�`����P�`Alau�Yk|�Qo"f�*mt��6U�POZP�+jf^WN�ɏv��ϻS���gB�h+/O�cj
�2��ta�CB(a����{��4p��c���g�H�b��U��ƺ+���P?1�2.f�[��sܢ�㺦�r��]�y���먾 n膐���2�BE˻��9���y}�C˽�%_q�mO����;2��Pt�U6%�n�\���>^B��/;r��5j��h%�A�e.���{M�e7�ʷ��=diR���kM��4򖱌�|������U��&}C�-�_��ަn��kNzx�\5��ͮ���d��L��`P��1�f�#'SG��os�>��/�-���+{zͭ	�h��n���<w3��t\vٌ;!"���GR${��:��R/*���,Ö�,vNg�]�ȶ�T	�^(4y8����>�i�a6�d�i�nV�2�-N��\{�+hq��z�����	�:�#c3[���&���_hN7$��#�;���'��q"��č'�z��//6�(�eK�İ��	 �/+���;�c��wf�B.x�D�Ϧ	�H�Z�ئzr�����Ez�q���}Ϲ� }}��y����a��S˛�Y;�m4����,8aPLݦ��!ɣ�u����2��˲�|y<��ޅ3�Gc;D䪜�mP�+JL�N���a	�BU^�8`�x�9`��d�3AY�#��T����㽴���*Ü�|��������G5ҫ���*x�p�z]�\D����a5�q����ap1����hݘ#��Ǩ!%I��[��[c��0�QX�K�p���Bn�h�s�	�5��n�Ĳ͌i�X��u�^�]6�m)(��B*�M�q2�b6�m�k���:ؗX�e�`Y��P�{Z��8ذ�-n�b�(�bV���e�JĄ��6��ma�Kqs��'<pb!C��ّ-E�>�7E/c�|�`y'C�2x����</Ǉ'���ˬu/�7�x��M(�%&%��	���th����I0h���T/w2��|���L��4���)���=p�뙳#��n���i�١��Aw�Ⱦ�i���zէ���α\�{O�c�Fp9%��V�}v��6wo=��^J�Nn�B����w�o>Oї ������Yxu�)X;�qK+���	 �(I6!39y�w�=2���Xϊ�}{p�]�5+�@����-/�Co{��P@���*��ϲL���c�ɚ�SM�	?�!+�W]vr%��w�c.f1�Lo7�휆oz��"m½�fv�LW�J�pƓ����+�n|����[m���ސ�1�9R�}����$�nENכ�*/�P�{/w��ՙD.Q��<�~��;�G�\Y��W�����X�Υ&�u{���c���־���7S�\�Ԯ��.}�����s��\�M�K�p�*�_{yt�C�wV�xn��$^)�ŽR1�^�D��i�1��y���
��e���pB]y�2�F�I��:ޜ��cu�0�$%�Z��޺#�Ny8�{��s�23:�D�Y�G:�ͨ��~1|v���Z�p���إצ�����г'�mάyf�t��Ţ��8%�-= �QK|ܵ��ţ�����0T	;#(U��a��)���=�`H�&�._Sn�|��D���'�&SF=�~�R��(yoT����*��h�kX�x+LD�dPp��A|�f�ة�:s��ֶ�\:�X��i&B�������m�ΗæNʺ�h�����C21�S�W�W�!�-xН�i�[��橳��$F�9��"})�`�}_P:W30�Y�ʧfǝBf�{6��G9a�]>�w}����Qʼ7[#71��_@$G�5�p��h��پ5�'5!��1�B��� �Q=���D����W]nb�R+��3^ڧ���S�#6=�޺��T��4�l\�ݺ��%K�,p�-ܮ���)�`lE"I�۽v���B�R��kV�J�c�j�����ݮp�늇RWvV���{�fx�2,P�lQX]��w���c��D�#&�D53SN��z��TeN�_���R\���rm}�c��{ܫ��YԶ��OW{Wn�W�`��vj�9�}�B5�^f�\�X���j�F��Q]]r���<@i�p�pE#q��sn��0�ڂ&=lM��w�}����=�$[2��5rV;\�Ǳn*�8]:�G�d"_$�$-�&��Ɠu!���&�;]_tn��We�����K����~������SYϐ���1�����o�	���a�a��ë_��P�W��*n�и�w�ܣ|��/y��\��8����v���%vn��.HHp&�j9M�Ԃ�8��Q!�X������;a�,M�2�$�^���~�щ��4�oX�{�[J�}KA]ǽ�ϫ��d����^�
Wglm:C�v+]/;����ڼ�
ؿ������h�ޢ���cƸ&�|�s8:���#�27m{7��HM����'Յh�����2}3OC��JŃ.��3��n��eM�ǡ�2ߖ^嚅Tv{Iٞ��7f�O�>�������\�*	�F�wn��^,%��+�������J�0_1�jfV�Ṭ�I�e���P;�Z^�L�D��l�6a��n��gVŅ���}�U~�B�A"�l�n�ϠE�dj���U�:/
�v�g:����c���%�����1���m������%�45Q-�At,e��z�7�͹����ٙղd��<;�Ϊ�;a{����yz�G�'rg��//)�G�j+�`��@%���:�[��^W��)h� �)�p9��z�G���)�Ox]Ù�u=�O,�����z�l�%�fjMW�#t����D<U}�����4���(HxڼǇR?o�sS��[�c4�T���ó�*uvz�J�W�$�v�+YІ�wP�I��v\Lń��I�^�vEn)boF"�2���a��c��?��;@G{���'3U���*��c@f3b�XI����][��T���W�K�t��Uo���u׎�}xRKA0usws#�m����w)�T��v��є�E��[�m5f�d��X
t�R��p��a���4�$����xeMԁy�-�67[*�ᢨ�Б�oj����u�Kv�(U�ͻ���,n��&v��t�s��'�o��*y�)�����+B��!\JZ��-�V�ru]��YfrT�y�]Q�\���^	F�u�-��)T�zbo����q�n]'�ܲ7}��e���`)fhcuf�ڃ���E����Yz�7����5�_s�h�X�%�SL�0����N^�]l֩�G߲Ѻ�f��]c)�;��x����ѻ y�A����g�v�E�x[�{�wݕ"ȇ\��竆ۛ����ۺ�U���A�\W��.Bo�<�r�-��F�c���f��%fi�3�'�(@7i��Y42��K���q%ؒ���/:�Q�ܬV5Z�����J���n����zŔ[�]ա��7	��Pi��3WT3�R#��6:-H��C"��ޕ�ʽt�"��7p�3"��ڳ��S�]�ǹˆ�ԕ�h�X�Ǥm�j�]�N�A:h%���Bcz��Gf���+u;��z���Y'\5�Ppի��nXDy&��Y�?:2/����D�C����#N@����-��\N�Dz����js�ת���72�� f��Wp|�hi�%���l�Gp�i�`��q3�iq�
�gZ#^�xGp���
Փ1��	���G(�!d�Ty�}���X���׬�p8��VD� �>v�,��@�
h��A}�W|}�dX�o�{�1��<d�ުp摁�K�����x�4��W�<
�'��V-w��� �YR���OD���wT�}w÷�`[����})��{./�p�j��	��ܚ�� ����A-)n�x
�J	n�1���F������D#lBDk��۞]�w(&0oOWb��;{���'���'�|n�x��j�v��ko=�uZ�ܡ**��	� 9[?��2n��Y�m������^�Q�'��Xb�.��s�^�v���e�>�57��=	�w�泜�	�}K(C��ڥ��D8!���v}��N̵�Q#�V�[�����6US󛤣@�U�X�%�׺���QZ7 n��z8+T�(�@��A��\h禸D�w|O40a&	:+�o%G�1�ZGa	엞��8E<Ve��=�W�{&m����S�o�d��u�:������i�!!VQ�l�ܩ��	��c�Ы}yRu�K�R����](����#���0�~o����5�j����@��1�X���.��` ��ζ"�97m�`dxL\]C��pu�Tɕ���'�m��qV��Ou�7g��p���T��v'���f�TH���J3���W'hӮ���6��P���<�lc7��R�����fx��%i�H��Z�׶]��G\�'�/f���Ϫ���2�^g�^���Bm7$"��d�QB	c�����~W6Ǹ�`�U
^Ԫ��&V���+�k�<'=����� 
pꍁ�f��������}\]�������k��R&n����L�D؀�@ʇ^EǺ�Fu��hPo���'����c6�p� >�R���&�cY,�k.l?r�\9��܊�)���#�d����\��f1���[D"�
H�d�n=W^�e�سgFx !�����d�0�n���K��]=���y�~��Z�̺���Nݘ����ț�Ɣ�_-V!\=H=�<��K����8§���!�;�/c�����v�)g}Xo�<��G)����Cc�����'�}f�G��AaC��Z�C�U�{_W,�v��<kF���QC�����f��2_�d�
�U�7�tf�p!d	������={��d��f����Ug�O4��d�ล^S	`�~��W,�~�>��s=��[�8��b�2#љ�Bh�ews��|"���o��P�הΈBA��Ϲ�Z0�$
��a���j~��5���_���t~�Yn���办��wϲa��v�������ز=�4|�l��`�f��Hh���9 `hw=��;�x��pJ:ձVky78!��u
3�N4�W
j�I��;ݦ3��_����=�.��y&�� a�	e����������g��9<2�ӌ�z�b���Nu<v7g�'���p�B�.M�3a���tn��L�g��{$���W�Ď��S�����{U������=�@��7�QR�o��w�l��=�	p��"�"O����V���ô�̿u}�i�ms�/$�xx�7`,���j,{��WyzTO�w��B��ζ�b��d��쿶���Ó�{>���ű�tZ�
�
"y�5�z�c޷�V�4<��OIr�pI|�� �����3ϒ�a�\N�9�����j_�苸�.n0� q�l�z�T}�/
��G雘�ݽ4��{���ͬ#E��v�p�C�;W�(������Ȼ��:*��,c�]{�B���Y�9t���e�}!��~o��!���}�V4�8&����B�j=9�H�.:�@�ڌ5n7Vv�	�j�"�W��������6{4�Ӟu|�T��q��/c1�'W]��YS�ju�Md|�;����oN;/�_P��Q�I�vE2"����?0�&�rD�;�7GF7�U�����*��g�o�r�ns|j�۫؟}�2y�Y%num�o��1,>����"0�2v1^&.L��\�W9/��&���Y�.k��'�>��o�ʏ�ITh-@tS�%{wt5m����(p���s�4�K*U4̮�#SO�h�	q71�Y���]���U=�0_�{���3���l�I�p^:d$D��b��*�=-���t�k�>��e9����3>�7��R��'��W���yW�A�X%��<=�xbu���N%�%���V�[�G�� ��%�L@��r2s��Ӄ����q2a���+ޭ�U�}˝�_�$�i1��5�E^���+Ff���$
껄T��=D� E�F�sh��rV?&���b�?M��[�����XS{�IX<&��	��5�/����������d���ا^y�e����w�|i��N��-�9�s�W9�����>�gH�|;HK��Յ4옠$�I�],K
�ŽZ�!)���A��=W\J�Wn�-�����������J��yB�z_a�#��;��B�?rRh��OON��**
0�-ff8K�sy��8E�zEBG�ns�t��=��!��b�g] gG���jg�����ױv��6�}N���]H�?>{u-���Є�#.2�!K�<8�i�	���[��K 
+��R{���(騆B���يe��mKƵ����e�n�r�X��e�Q�Xel�����7�Xm���TF��zY>c�<8n��i��,-�W��u���ɩ����_N.WCn
^͕Y�{��A�m;���{�Ԉ8A1A�	���y8�U(�s��k{z��+�Hi�y�н#�
�ž��l��K饄�=ݦNr�b��U��=<gph�+[0Cn 4
S��N�~�1����;�VzoF���0 �^�釗���2���|$nTl 7 �����=�1"d�t���K��\!�����v�`2�p;��q��EV�H*[2�~�r�e]�P��+���q�9��uSUƛ;�Ma���1p�d$�p�#%����&�q�1Ch�����գ�&��.vZ̾g	��@��Ż�oO��{oS:�4��@��L\��t��z�	��L��:N1JL�s��U�9�I�en'U�c|��teM*��|���tO�/�,���Y2{ݸ����4�a�pA�͋R`�������2��lpTg.c��(�v��~Ϥ`M�k�.p��SD+��5ix:�֗dlʠ��N`S���� ����f,i�
�`�}���F�-�}�z���W鑁����툹�*�D�W���!%�
�ɼxA,;@��Y�۝)䭗.2ƃ�f!���εO�]CB��#�Ƕ�����Il[O'(\E��E�g��4~��i�>$�D���j��`P���,�͊��K�P:�.LY��\]��f.��.p(U#�yޣF��n��0k4��f��..45J�˯n���벼���!V5�S�^�nف��l�)MT���qס�xA"-ĹH(z�ף\����O[n�I[u�V�k�h�ktѸ�Z;s���r����
.;���v�Pg�L��#wY�=t�U�
q}��]�����8��bC��W����@�w{�nߐ[ ��Q��������ز��h�4�@ڢ�}�KzA�I�>+�9��g��½�i,&	NI���I�,��n)�n��LF�ʦ�{}��s`'ж����9�m�^t�*ʤ݋���<Kr���
�N4������ۘ�g��v��z�t6����f��Zk3��>L h�.������ܭ�dw�$
I�^�s8����"g;
�����Qb�d?��g�C��h\�	�^6f�͍��<���D���ʢzk��dnE.p��C,�YdX����e��h6��6���?x��k3�lp���u�;}ν������.eĉ�sdk�w7�=�ߧv��[�_@I4�0�Qr�t�h�׷Q�vO����7y
_͎x�;2���ߍh�������T��j�¼����4���xG�m��Y�䍍��?*)�)*5�A��4*��=��>��Ew�~7�Ԯ�w�4Q�c8�����x"����~�)��]���[1���8:�=�wO��z��5c��m1;j-��Ev��Y)�È�8f�:�@([ћ.�1�<c��>y��
���2;׭�^����萄WFA�)l2-�&/I�1\h~̵j�_+�@t����9w��u�%�E`�|�n� �sI�^{:��>[��;=]����:s�\W�/����������M3�33ݗ�1��Y�4#�`=��G�V5���	��T�;�{�)�n�\�l�SZ���x��N���3�7�g��n�ᆆ�O[�gQ�ßZ���=�͚�>�}/�_5�j���^ Q=z�Z�Ɋ�#���M�a��.=Ͻ��>�{������f�N�
��D{D���7��,�qS�'�=���c���=�X׃{=؇��ପ��]kw��z�hD�!]�/_��sx�3t^^rHP���Ӕ�rlo��+X�brd,,{���C�6�mdTV��4@ʖ�]����Vߖ�p�&��mRM��f��{ �N3b��lHW�3 �����[�����E�oUV#/��d]y�C��n	Oط}�ozQ���D�=�4�� �*��6j��CE���Q]]�R��}H`3�b�F,X�+t�B),�����&U�岻�EgL�qnD�n	'{s�/*3�b�1=^���j��h��:|u��	\��<#�MJ�+۬��՞��LV���n�)�j�
TxDa7��b��xN#�6���s��8�)�O;(vL؋��WB��.#E�,S�ԓ����y��DsE�m�l�L�;`옻k%������ك���z(��Ùҧ�s>���^�9���I����c����,����Og���s��nS즧/�O%�&L�^c�x@��/s7� oJ5���9�ܝa_WD��Q̇e��+'z�Kq���wt��`��xfzW�G��'o��3	һgs�j�{�\�	AP�P�DK;����MAP��%gW{��ֽ����m��_A�ȹU���{� Ôy�˂<���·�_�e���~��@�Ad$	����́߻��ޥ&g�*;������j���2}�(j8���c/ٙ��%�k�w���a��&(gq�y�sh�v��/���S��0A	�e�6}�+��t�W>�OR����e��C8Ѕ�ܺ.Łmm�F4єM��i4�9�Ҷ�_̔�*�F�~�~�C��x2�@�/:O�)t)�/ty�ɉ��<��c�n������܅G�S��q���>p���Y�-O=^�3`�����������$X�'�Y�gA��_��A�<�&_�9�i�W�i�4*����+-v���a�(�'�\n��]���b_�p���i��P跶J1�B�u�:�%..2�]�� (�=Q���ś����#+.�Y����ܔ��$.�!��U11៿G���io2mˮ�e�ŗ+��>�Nɚjs�����?,�>�u�V$G�ل}��H���9��((	��lG�I����V{.j8�7�KWN<D��^v�Z��_��R�&b߷R��Z�)�|0J�Uȩ�Da���[�Jx=һ����$�ͤ������1����j�m���AN��{�仴���Ώ,;�m�z�Q����\�'F���wef_;�l��V��+����]��Rh|WȰO�r�|�Oe�S�R�3\���ΗUfW�$��K�D��ɠ6ۍ�IU���X�3@+[H���`\L�h���Jޢ�zs�l��!F���L�uF�7Ϥ�����OǄ������5�TPN�8��ϨNOh�4�|SD�U;����Ź��C�uHwv���5l���c}�w��՟N�4�1��7�J�¡u�+�w�zg~�4k����x࿌4o��A��u��yod��+J���_+��B�j����K�o��ɏ�l~)�w��Coe��/Z�w8z<���;0c��4%	�l2�r)�f��\��z�d�����@��mS�Ն\����fF`�Ej�8�rM��Z��,"���1�"�(8پ6d}�Vٮ�T���qw��77��B\z㸀�"ͥI$��R�J�M\u��.�H�.����6[#.�u��8��b�gK-uF(�Y�<[ǋ�2ԩ�i�&y�9�Z[t㲶R9�-4����[k��O����i\3M�������Z��BF|c��.�\۞4"����#v�l�u�AÌq��k��Ƀ��LG;�65�4�й�����,5�%���-�a�[[p-���}���#����K<$z6J�3���劤y���s驞��&�8I�Â�u<j}<x��b��իO,umj�@t�cR�my<dx�Po�	��{�o�2������-{�x�W�m�_s��}��J��p��i�nF�Ci� -�a��@j,[�]T�q�;��}1�M8|����p�i��|O��ŕ���ck]��y����ϗ�r�6y� A"7h��.�1E�7�j�.xGz�����}�`��y��{�U�?��&����	W`���G�=��Q�25�d:-7�\>��ڳ��q}����������������`��g��b���;��዁������Tvdh�Kq�P���Tw��w
'2���u��y젎�ސ��1s�k8ρ����з|h��)���\�Um|'����K��x��L�}U�KՖ�t%��M����\�0F{2����Oaw��u�3�,jO�ؾ���=�9��V�0l��W���P]D�^zY��oו���`T'Ci�i�x6{�˱��dw�h��{���=˱lᐥ4���I�ZO�?�U�ϛd10������r٩�V�}�}��PްCM���1q�S'a��K,)��f�h\�Wܺ�fR��N�Ԅ�k�j~I%��K��u:��[��hnb]��m�j�p����v��
B�D����z��sk����j��s1]��*��I�a���T���[�	Oe�X�s/2��\��ZT�\7H3����A�E�e>ը����v��kT��%��F���B�i>��M�bv��wWw���u�����Zqa��e)�7
���nM��~��Ce�����4Z{�c�ǻ��\�@�=v�g��ui�1C��/v�c�5�y&���|c�7�0�J�O�s��4L҅]Z::�]�@lbf!#�y-�J�U�����WU�c�Y���+TӹO+��(́
���]�=�%vZ66�f�b�هU[Qv�r�Z�����pt��ų�.�I��`�S5�F<��-�|I�?����pХ�c���[R-��y���v)qt8�D��^I٪���ڕ/�/��VL�4ZD
2LV=�M+Ո��Qd�BT�v�N��->�wݵ����oJ#u��,�ov!�o��חt�V+y���v8���u�G�@n���;S2�Z�K �P`�e0��:0�\�`O��s��K��nB
���O*����v#�[���w�uq���Z�=(E�
�/��"d��t��KE�ݘ���(���V-"[9ץ�l��qe�:ڭ�3��R4��0b�W�^�v�Vj�m[�����N�j=oL�׊'�	�M �ɩ���&�>��p��j��5�T��B��UT观k���d�;R�QUT��*�٥j��ET�K�n�y��n#�օKCu��v��u��Ӹ6MY�T!�|��;����������GN��0:��m�����c+��C���ز��^���1�c��A�Fb���n��2���nڃh�l]l��"��]���pT]��g��f'�]�t�.�@L�8�U��1�om۲v�7S���W�I�Ƚ�v��&�8�*�ģ�WpݱKn
��QЙɴݥ�(��v���J[omT;F�����GLJ�����j�ɗ�:�@����ˉӓBF�n�YĜ͍L��a�.�15*�"Ks��;���h�34��:���\p���z�c���������|v^���m�v�m��iӹ:B�n���r��u��V;bs�͎#uBo!j�U:��,��+.�R�O�NY��|c�ޅ]�T�u��f��z�/n'#uڎ��r��ku�2�^5�k���nѼ���,�R]	�1�Z�YL��e�B�X/	��e����u��YɬkL@��oh3F�{U���9u�Qn�#�Q3o\'S[�-�ι�h���t:�DGE��{%�u�ު� �2abYd943��;]�KÝ̐>7d���wn���*�ݓ	e��R2ڶ�\s�z�U��s��K��� (p%�C"<a�,c��װ8��t[1���D�tn�]�[�5�BP�9��r�:��Z��J�	ri�+�6r	xuN�����^�>*X�:��lm{D�A�,0�0�70֚�F��D.�V6��K\W��s��l�mrJǭ�m�W��YT�`���m��ݪ�%��D�f70������Z�,7U�hR�`�Ym�ܐ���6*��Y� �(�[Kp�pt�X�.��û���%ե�����*�Lަ6f�篑���6��4e
�S�۳�B���vd#s�0�Q�ĉk����Zt��3pAv�BgCQ��sv��`Zk5,$Æ�.$"�:mIrƈ\G?ߢO�17�hJɾ��6{�.8!�3�>���Xy�`�٘ֈPr��c�`]��ZW���Ӎ��p�#g�$�c��ir򝵷�3�ťs+��!BԻ`b����}��^�-m��ˑz�a�V�d���z]�3��>8��/w�w=���ΐ��{�,2\p�j��r�|�����~����vx�5u��"W,b�Y9����b{�Խ�"���Z/7:��Q<P�ɮ�7�+J#t�M �l��	�hL��Y#�5x�o�h�Opف�<��k/Kq��0L�e�$����m� �\���*�}Z���[�{�IR��u����>�5!�� � ��oZ�JS�=sx�������ߕ�%���'�{��h>���Kd��Y�mFT@�~�H���g ��)���E������[!4a��l�=&�*��*�#cjuZί=[�nL�^�0{�Y�����{���ťڙ��z*��-�c�����v�m����2�Tb	aH�j���Z����嬨\%@��u_vJ�AJL YF���m��:�2^t�*�D$�h���h���)+��S^k n�ʮ�R=�f�ȡeg����o^��4k��Ÿy����14r�`9f��]]X:����9�w�ł�ya��r��\Q�;6U��]E�ހ�������ɽգ2VmX\m��n�]�����a��A�X�}$��c��=KM�;�҆O��������T�}U�o���X/�؝��FyB�x"Fw����o�V��xt<T�����K�1��C�g���ꫛ7)��Й\��w:���Mx}w^��W����L�P�Ylp�|�dWT2�=��ә�"j��u˛�Ez6u�SMH ћ�F��y{�NF��1���{��SY��wZt�f�`��ɯԄ[�m�[�4���q7-{Ƅ�U��;��	f��L�H�9|{����{��y	��D>�~[������o��8��3aV�C����d�3R�gHg���󙳧���b+�\�2�g6�$1N=Jb��ˬ�%}�:��ޮ���=k{�U�?��C�D%��r(��f��b.��IiA'���ق�%�	 wI���zu���K&b�+����F����r���ٞ��ip���0�7},�@Ql&�}�O�#`���
J��A��Y�s�:{*�F �}�=Gb��w�Y�}��KV�'�ڧ|a���k��}���%A���y �=>��c��q�'O;yP���t�r:2�ȳ��ma�V�re=3��]�B�4v�,\�p��sF)"���`��F$��\`O�.�Օ�2浝��5���W�Ǎ|��̶���΍� ߾9	`���}}>��q1ܘ+��×n{CXrљ@�,�Fx��y0#x{E��l���YgzO������Rھ�ȝ�l�[F��7���`�EX�M��WO{@�0��K�Al�z�IX"��d�1������)'V��.�ln������|ׄ���+^��������cng}�sq�,ߠV����kw2{f�����8-�!d�q�B�p]���rB�y]�+B��	����jʔt�(��(��X.�Ne&�3�����IVSh&�*���F����ӂ��n�8����=,qs���vl��������T�%1�}��+�����&IC��s_z[�6ҭR9t���)�s3���uJ7�\�� \`��/Zm`���	lGxL��U�V�Lu��W�v�(��Irh �Yp'�=c�=;��27����豝Kw�i��a��P�^n��C��["붶��5{-v��:�w�"�B=6S�ە�9��g<����{�Q�&�22�w��,�Y�%R���^|>���P/�{���߻�kk������;����rY��F���!�@f��1��PO�u���tk������ʜ����1�ԯ���Z�<�C��ϲ2 ��78��ͣiBi&�'�ӎ����G<�n�51ɒA�#g�}d�kyOg�؍�Z�mn��%ti���?¾���ؓ�Nup��kJˊ��A���I`�)l#��2�\SJ]K�V��֣�9�j�/&z�خ.y��@��ӫ�*���c������,�虡Q k��'�)�n�ܛ�n�2��V���I�ě^m#y��Ã8�ng��_���k>���/�.�����iO`��}1zwe\���s`��)6Jd�����5h<��hP�<�Mj1'���>ҖVM��V��Y�[����Ȯ��P�k���{�o�tI����E'��w���Hhg�Ul/f)���N���۔��o��n���2�r�u��%�p.^jT�6��t�į7Mee��l�Q-y�Zm������Sk,_b'
��';b �<F-*r�1s彦v�ň��rس/������e�D�3`�0i
/U��-
}�����~��P[K�yfll��s�}cϬ�D\��VV�y�Ώ�y��[vF��V���Z
3~�X���f���K��	
|`�/���y;��d�9�d��_���f���T(8x��#b��ިʗ�=�h�M�uR���!ۛ���Il�҆���I�b['�֞��`3�V꾲�䴝���[����ps�g/pU�ޟ�^l��w�5O��oz*��&�4���3V=���M�#�8�u�K#[~�/#�R���p6�yw��]�i�*��9��8��[�\����z&�,�\}�Z�׸�v�3Rm�k�z�X�ʰ;�5.�+�����k9t���Y�9���f�yw9Ll�V� J�8o�5�ΰ�d�����}�%��}�HM\�{��{&7��	�KP�9 sX�1��5�/Ì:~/�=����e	��OY�{�n�t�4�S���G��2�d� ��RZ�o<�Ŗ!�&�N�7�"pm�L�gdmڢ���b{6/:f�C���5���7�j{њ����V�5���A&����ڮ���Sg&�(ݭ����)Hk���<�O�`X����aH�>�+oa zt�\��gu]��S�a��~�1�s��{ލ�7�l@6U���; ｾ��ج��;~ 散�U�&�ଵ�"#�/��i��gFi�������1���ϻH��{��>���}��6�j	L��3��H]�oWuOeG��Zyz�%j���L`k�y_���	�(Õ��=p�=^����β���,h�?<^׻yk��W��^�{���@�p��y��YPn��FxH���rW��_W���Ӧt��ۭ�3����J:�o�B@��z}X�n|�5
Ux�Th�|�4S�#N���ǻǣXP� �a�^��
`�x@���&��s�x>V����5�z�-d6��.ζ���m%oA���m�(PL2 h��✷If��C�W9o�j�Y��.��O(E��X����b�U��uݽ�Q3�����wfNV
Q�
�+�!��̦30ѱ�@��c�ԗ�$���6�L�}�l�z�������T������a �Ah)�&�X�j��9�W���vkq���龛aPs�#/&�N���;��1��0W�ً�}�7܍�����Aޝw7��yCm-��p �Xder7��49e��WnI�dP�=��[�j�_�b=�/O�[ޕ~��ɞ�ZmJE� {��{z�t��{�����nl��!�G��89�1]=�(���W�e_�=���y:�����D<�z$����O�Le�H��%�J돡����Q�"�fu�ˋ��#`���A8y�AGm�ݠc�-YeU�&�>���d�F�9�v�K��b����s�����3��ul�;P8�&$|�ow����=Њ@8�)zn��6@ˬ��H��mL�|�ͼ���~S�S�:v�ܱ�N�jCn�ō<��]u�٬��L����T�o��p� ~7���eg2�^������5顔�}fzo����e�'�ۥ�����O���fl��I8A8M���=ı1�U�ޯ�]p�E<�ݯ;��1`�8<�#�
����S��(��Ȥ};�9��
 ��V������w+���"��f;e=~��o ���[�E:-w��n��7��y.M2�%?*9��۰Q/��۟�L���p����(�y�eۭ��#����]N��`�Ȼ֒��MTy�E(��4�R���ba��d_��ǥ���-���t����}Rg�.�$?i�q����+T���[K$�X��t�=ꚿ��!G��'�w+b��#{,�#q���\燐I���H$H�뫙�7����{{+�����85��0YQ�	cP�˒:򣹷�7�s��X���|+�w%}~F��^�e�2�:���tT!|�j2��`�x{=�J�7�?c}JN{��Əi�O��&�A�8�^uE����U��<о��6�� �o˭�!@,6!�Xd����`6 <�Ѻ��ю/E��ல� �d�6ЈĂQ��@�_��I��\��P��ǖ���������I�ө�h�=ۘv���˘�����- �v���d^N���>(��)Zή�f���'�x]�Y�Ωc^�H!�R�w�g��q�f='�r�ﻏ6S�n@W5�hC��s'�Z�Q�j����}������(3zOl�O���8��u�ڸ�~jz~�������A-��!������&�kƊ��G�����a��U�uu}2�Ɖz��5��k:�G��h'Q<�;UlȖ]�>4oq.��]��Լ�8�ɚv�i!f���W�*7�����X.�ِ�sy����Փ�qq�v�ZNH���a��Ʃ����2�\�6�nF�4���0|��Eȹ{vmq���S#���s�J��f�ӻ7 Rj�-�j=cE�i��vyc�������y3�n-nu��ix{�!�����#B��l�uݠ������ i���4�Y�n�/O�qO��j����ŶP�`�,c�؅M����f��Ft��^�E�V<�C1\ iu���d���[��n�� LP�h]�-��M��T�C���z��.e ���}�s�1 ���5�~Y�3~WW� z�s��:����ܦ�o����Dq��ȿW��]�H�y�&M���ĳ��p��x�j�7h��l��b�3�.맦P���T"�LC.����"v��\���C�!a Ԑ�S�!�	�=�ݔ��#��J��D�h�8V���I��{��q;��!Oftp��e�u�^���($��b�k�8W������/�->�W�*=�"I��1�rJO���R��%���K��v9��<J���j��j[ �d	:�$�G^��Y���k,�&<H`˙��c��>�I��+�{�B�W>S��Xk����{y�	���j6��*�85������:���8ۏ�$j�Pk'-��E��-��p`2����U���}��~�:�ՃG��t���1���(�uk���t�;8��ɸ%(d6�w�K���ᯤ��η��YJ6D��U@_9�u<c̚�*r��b�;a��%[��ܮ�������<Q���R�ĺ�$Md�u.]�V%qL�vb��i��l��w��3״�n Ee�o':�Uѭm;���66/Ͻ���'%P�s���Y�O>!���0[��W[�f5;�bDw�+GM�B3�bd�0 ���ī�E�4t���u�3Y�|�8�ۮ����TL"zx��.��;\!^40A!ue/T0�瞻�nv�{�I�4�|Q��Z����ܕWX���/A�CL�����w�*[~��;���Tڬ�w�g%�5,*P��3~]���?{&�|�v.��2Cx{�׳q���z���T�0UOb�j MU��L8wF	:L�H���@��������1� fa����=���\�fZ�W�v�����b�c[�8�<<M�X��eb3ccY	��h�.���%Y��׍�ml��N���_8�F�r���Z�t@��=�>�oK�+pߺ޸�8y��(�WL��D�J�J���R&��=nЎ������B�dzu΃�G7�_�b/"����?��ۃ�.����x�>�O�Fj�Njъo��l�6�&�v�p�-��-��1B�4��Xt���Os3WP�.� ��M�o2iջi�o��ϧ�U�X�[P'�<�pty	��շ��X�V��d����W�!�c���u�z��#���^�ڦV���!{b"�ec�<�Wf9��|Wi���V,m�)��g��&+3
���uM��aۅ1�2���z�T���ז%��W|,����@��v;�����p��ئ}���jn��g�n]|��x/jt�g�q��|��O��[z�N#s˸�s�1�����(pXjD�R��<��x�ݽt)C�lW����/Tt���峷y�^p��[=�=.GަHRep³yևﱩ�E�fz�Ҽ3l�L�5��!���6CN I��)�(U�DF��&��j������wČ�:\׊�Gd�9ᛇ(�[�����KhIׂ�w����{�=h5���Ӑ�C/�λ�=�x��!�a'�%���ƕÎٔ/�1��U|%��o�Ϧػ����傭}���B��d��/@��<jMv�N���6U�w�w�b��4���0�v��R+�f�r~ᾛwƱJ��� �2
�0�e�LUK�D�J�x��|X5p��Fe�n��ǫ���+ؑ��ں��^��#�Q�1�Q���8���r3B�bW/:wܪ*�c�F��0�y3���~�j�9�-	h��R���ɔ�ñ>��|�$�4�g��oV�y|�2�U���3��0R��3����}��^����wg>B:6����ա�"䍴��{���D�/��O���Z]D�c�k> �c�*��@��9F��w&�T��̆��n�ob�v�ٝD�}�0��Ns��l����xC�U�+�v?;�{VP��nĵ�u�6����gRc��{f��?�lъ
�q)Ʌ,�+�ŸNhu}YӦ��Wu� 
��5����T����l'߬�>#&�p)w\���K#V��W"�%����	d?��^-jL�(i��.�  ��j�e1�p� 6k$;��&��o7\��'JàG���Ü��|��J���������t��	U�Ėk���t�n\;�q'
�ۭS��St��c�lVC��ڜ�]�w᭭��by{���`�6���ۗ+�A�W.�W�BNu�����W��jA�Ů��M��T��K]p�$�go,�������η[6���#�Ju�K��l�Sfë[�s]ב��/Ɋ<�u�[��u��gl���_�7�b8�I����ଞ��G6��	�`}X�,6i3 E����9B��ۜ����:��5�aA݇���Pi�p�E��%i�@;�7�:�3��v�δe�1j�O�l#ϼw���^Z��'
��ʺ�yʋn�>�puH`m��ܽ�9t!�w.o	�l����;f�wV@uoR/_A����5���M%\rb#��'K2�%g�Y�{_5q�[�����4���@ؼծ��p)W�3��c�z�#.(WS�75w�}��&NV;f-�ɗBu��2�;��Y�cP�ұs�R�j\�.�?��?�v`X��eU:hқ�ਏ�;�Zt<��qn.x�J��A��T�m�wrg���=�ƙپ�)p��|� �d���q���M9%+����4eU>����1.�ΐ�f�n�0�3�������݃��9Ϭ��j=��O���ۚ�=�KE�XI�!��̘����E;�(_�.�3��J�e��@�����zk�gx��4V��_&D��ضa4OL�;~bĩ���^[���R�w�v���Р�&��	:$�#]YnY��6�.���t��h	찗� ��u���[m�\׫e+Y�F�ss�Z�����rw'Y�"h���jQ>�C��r��fo�� '%^��.�*_U#�m_��o�Y���s4��l/;�S۸u�A!A�D6�b��U�|�VV�J8
j�W�c�xu61:jb6��	�b�n��9&�9�g9e�t	\�@~ʋڜ�~JqðQ��p �_�ԍ�W"��)uz����a���ҍB������V`�b��k�˽/�kK��� tS7s�%<���}��zcqck��O�"���i�M4�n�:��׮bv|���e�]$j���Nŭ"���yѦ�P��:ǻm�5�;���9�\��aa�l����r�UvΗ���g�]Z�o�!Y�X(\_ӂ�;*#��b�� ���jJ��=r[7\k���A-�ۄ�p��%�%hAڨB�9t�][����|�h@�Q�64p�:��,L�Ά��2lPky�`���u�Q��P`��^W�6�|�ۙ[ļgq�څ�ن��nNMp���e�#�<n��:�HZ�
^F-�4��Qu�CZ�"�W0���ڂ�����i���@�g���\W�go��8�A�U�U\�}�3��)푙чXl�	' �M��h�AM�K����{��-���t3�����zJ�Ǵ�4�w)\�\=�W����{�\�/��� ӂSDn51G�sSG�]���'b܊�|Ӭ�6�)XqM�[n�p��/G�����@���8D���3y��v%�2W�7�_������^�s�_E�A�![7>�22�/R����&$�#z���|��ə�q�"N{���>�q6�l?�c$*�P��G�-�]F+����C�̉����;	�l��˽�l
��,��Fx�����w�^1릎��w���];����i���~0���ϻ���]�n7xt-�a0@�ev�]������9=]w��{6'ͯud0"K�x���1�-]]�R��zdN��������G���!?�f$M�^�ᘨ��Uq4����-��{3 �հ6P�>#y:�8�of�=���N)˱Jv��Ϋ6ν&�Y�k�f8�-�;�S�7���k!�ű�`x�*��zjĲ�Y"�>���GJ���J�"S�k}
~�5	�}��0nk��-8m@i{[5�WOڎZ��il�j/��j
������mغ7/;
��	�<����	�1p�I�f3ə,w~��D�>�7��VQ]�|9kwʽfyWX_x*M�s�l�fte�IM�t�HĻ:�5��v�[�:���mu�h{�b���yHߴ�Psp2�z}�i�nr�8N��NJ�q��-"$ۄ��գ�6�_
=�XaY�R�UEtm�qv�4zo�c�K�^�-��f(�^�F���e�W���O�*�gp�&��\4%̈w/s�����<�#���[۲�/�
t�^�oz���ni�<|	�T�H����(�_K�������
�YlR���u�r��u���o/oe�s=P<����磮8�+X�K4Vg�/W,��v�,?;�C�u��h�������?\Ǉ��{i	Cio����]���nn��>������4h�b��u�&���>8u�b1�=g��4P+J���� �d��lv{���s��sO�os6oG��&;1�G�A�
.2�8�{Kʹ�r�i���#"76�@�@gX�,�W�7�������s�)J���L�XӇ��v5����]V`e����L�ա��.#��{���ߔ��~ ��ߞWY����u["�aUX��ԓ>ï�rE�[��tzC���h���>�B	lIE�/8��j��4�r��˩�0�E�O�'��ޓ��Ry��Y<.D�R�=S/�D��J�!���]{�'[�8Z˾�ۀQm�D��B's�Ð/+3Wݎs2;��8_;άMe;�7���.}��{@��\p�����{�ݡ�My�ל0���hS�c჆���y�_N���J��˕t����23��V�=X,g�c�����X��prGr�f+5>�]zdp4�4 ��A^OvffX���*��5*��_!� @(��0�H���e&�c�s
�ĵ�$8N�1�!of�ã��z{jg���57�"��;�Y��m��܄< ���k�w�H_:�D��;��U�w���Ķ�i`x���`��N�L�<��^�m�{�dq�S�'�Eno��,�N>��B�b4�s����饭���ף����,3�V1h�$웋f�t���F� !������S:et���S���+�y��8%�IN.�J"Аr��{���+z�z���n�J�4�NI�w�����}���}Ӆ��{�Z�ڷ]���|�	CHv�Ս�*>�w��Y���zf��3Z1p��:Xuzƾ�L`W3r�t
=v_U{9J����fd�C`��>�=�>�Ӕ6�}�m�U�{�J�T^�R�{�{d��9����=1�m���2�ڗ�kFZ�K��f=���,H�)q���e��Qw=��=f����jr�@�h�KD���α��$���K�ˋ�&�&ńuԌˡ��01q��z��>C�������d������7�+��"�vƼ�0������+٩l�ɐ�����|��c�M���]��6ּ��8s���!�J��J��~���*��47������EM����)�i��nHª2@�u�||���%����}T��b
�����*n��_��ڛhH|} ����ϡ�Y���:�u�#�ěoYS��̼��������zF�i��U�監;,	mV<ɻչpKE7�-t��3����kZPvV�ʥrMdN�dV��̸���V��Ūv�򀪭���-��]����^�;���/h+�l-[Ab� af&eKLZQ��t�������O9�h��6�2�mn�Zf)/7���9y%�*n��`@ nsڐ3X�0�͆ۦNf^�aYz�Mێ�Y�W�k�&nx�*��
VT4ٶ��dyr����u��>����({r9�Uݶ�0�Ź�i���U�Wn�/5tm�,�+f.�H��'��~�(�7�߿�]��5"�_Th�bl�^5�����Tim&bD�W��"D��U�z�ex�&{�N�	»����]��tl<5�3���ïi�ٶ�aֻdM���5��x�w���Ǳ������Qb�̌piZ�k�ӎ�k�,��΢H���`�㍦��-(���kmC9l���F�q�u�c��^9���
�Ç�\����[D|ʎq�yϜw�_-��~�l���wm�-�*����Q��L?����vCW�iGL�^��~���>x�G�}�##M����Gζ#ϕ�%�-���[�7R��މ��u�q�N_^"�DH�(�k�� �Ē��H�+NVŭ���0�P�l]�jo"�dyc�ڕ�!��D��)�^_s���.-��y%xH��%KG쾯uׂ��v|Jj
�cPz_���u����,O���w�>�Wy�\L^'�{����j�v��xV��F�tEzofb��$i`�`�9�tD4�}�ş�U���}hl��=��i�
��?��mLW7�5�q����$�uqJ���P&� ��a�k^��Ʌ��p�uvE������F%�"n��-ʇ�"�& ����:�;s��;�{86�c��ռ�Ϊ.�`�")��645�N��2��9�rī��n�~?{�9ˠx��p2ӫ�k'Gn����î����pT	B	��,1 ��fk$�e�%�7��^��__!�᷇�ҩoH���;�w6Dz�)f��l��*m�5Ya�}u/�/����+�wUCTӎ�V1��ޣ�E��ԳQ���Ee�/u��]�U����H`��<�����2j�r�a��|�,�<�XU6gn��Gz�F;�>���S���nn]�m-��J�{��чaq��a�Im��C�x'~�@�l��B��w�7�w�u����}�����.�Ʌ{���:綼c��W��5�` �m��V�#æl�&�}��G�m�����K���s�2u��������α��UҢ�g�5yuX�n=���ъo33^9�L7
dY������ER�u�� �Z>���.���د��{g��&�� rZ�6p���-�v +3�ݷ,�u6\%�n��Oe�<��'�y���2#�[/�5��3�A�o_WW�&���2��:=�&�"~����t��p[R�w��a�64,���T���j�Ŷ-II��0,�՗gt�� ջ�K)�t��Fy�Gy<�J�3c� �l6]�ȫs!�e�n�Z�t��de��3,
T�?R����b�LR�½��|{B��NT���	t�S�or\	�S%�� H�i4���V􃕾����+	���pTߩ�ha'G��ޫ+{�Z�O�������:z���SX���8Ɇل�!8(�V����Ve���%��ok��Y�N�S>�-`�������˾�82=k�{��K�l����a~��]W��!�������26Q^���;k��䏯��|~Xb�1W�s��C凅<���
9W��X���˘��~eC�[g�9���k�{�jg%]Q���B�i1f���.�䚽��;��Ļ����Q���bq�5Ӟx+f�kLl��Vݝ�2�y�']��w��IWԋ�f陼j��m�'Ay��80�\���4g��*5xGv�B����36I��S��U=$��Ӄh����jc�+}i9;U�e��$c�o�V#��c�8e�F����-���pu&k̾ �};@ffӚ��N���H�	6�n�� ���{�����}[*CeJY$��ř�w����y�\��x[����.P��s���&]�렮V��gVwD��e�^Ab~�w�'����ec�W�_?��w���\��EA��1/�y'���`�s7_O�Ώ�e����6|��4���A�1�]�:�N�{�{��{ה��U�\G�«�/�JK%��������v/�X�����)��=>�#��� ـ� N����UO��B���b��?j0#�E�i�s=q"/{/�]/�_9�:=�^kj�)�zmg�OdN��#*|�g�5��:�[��j`7��n�̘�I��Y�Y���'+�s�3��ߢjC�a��p�6�����U�pSn,%�(�K���;��)�Mڻ
�㦷V�Gҍs���cof��?[�M�^��Ǝ�3��j3k^T��lf�j�mC~��*' ��+|�����ʻ�0��
c���Y�Z{�1��u\��7�U0t�u����J��0޾=�m���%j(�&�� [�����dٜ���U|�1����c �V�8�1N9Ej�QKLڡ���`��-����sЛ3������F6~ ���Or���^�*���w��uU�2���<^4��39��\���9�r��)�fa��ŉJ!Ȥ�����[ȯN+�������ؔ�Վ��d��B7N��'"6��fWU��.f��1�#I%I++�-�틉��ͭ�8�n��g#)3L�9-��c؎x��7
6�M� ڳь�7:.�4�/�A���nW��O)㛣f�#��!l��ؗ,�H�c��F1ܼ�8kR1H�����,k�<���e��Yi5�q ܹ���vp=L��3��&�Ѓ,� ���/348�w]�)�gV�1fYL2�Y�t'�-��0[q���	��ץ15���D���?�ާ����|� ���&m��t�cp��&\0L)R��g"ruu_�'i����|cdr���J��z���؋u�O�=j��x�;m�Z�I=�ro��!Z��ز�&�^�� �H��%�
U��}�u2Oe��~���U����,��K.�ru����	JWq8s.� �+�)N�WM$	$�!�֏,��}������:ab���}w8���1����-Z
��3?p�(�"z�mc���ym��t&�Q�~�#r�f̥�������I��/�����T}TX�� �����e{;��kVy1�Q�E����?Dp
��$AF]'vyp���)���p�H$���Ճ�`��
ƛ�+���%p>��!ݪ ���4�#����4|�k���W��(�Ɏ��"~�j9����ޣ񌈊���p�/3n؆���D́(䑥�H�o��zk�.�޸���g�Y?*}s�����y��Ȅ�H����D��gN{�	Y��u��<�^�q}��݇��YxE��|��D�i����}�Ydvk<3j���t#F�̮�;� �0�8FZ��Ɂ?c��&~�C�� �F��s�U1#��C���A��ׯ.�nPŗ$h���w�f
�d��(%e��S��N�[���Y��l�%9�"��.����im���7�|�"y)���#�k,�zM��4E��	eNe�;�(�v哇�:�����:��Wc��8����B���7�.�n���wZ//��`>utj�3�z�� ��,9��jR������L�('�	ݛ�*���y��^P �AJ3�ܐ�ZQ+D
�ޚM򫷗]�m�N�iC���GD\u�5j��14_kٶ��-�-��P�A���t�}���k�l�G^�h���;��$)�iWoC�5tJro�Mz�8f���8�j����w��O���mΓ�6Wga�CQ���Զj`Xu"�a��Dd�*�`Uh�!|u�������@�&U0�ۓG	B������Ťf����F���D=&�)��"oa�ǖR�������V��&�ܤ���=(� �.��(,7������\v'"���Q�Id�[��d=��Os�J6�`;�Ǒ;k�Q=
��.ؕ�� M����*Ι\��vY݊V�����[IL�97gq�%t_�e%E�dd���^ȕ�ƍn� �YSSV�tY;vܸ0<7���i�,�כP'�ۙVp�
���ڔaͭ f���ѕ�:ժ��9�]����e'���Y{��E��Ofuֲ�5O�ۺ�O`���WB�}�ӈ���ή��Xk2��U�Lf���fL.egP�:�\Q�
XD<���z�i&�I(M���Up�(��W��#UUJt��T����YP *��k��杶�	۫ѶN��e�X&Ka��B�mt���ij��y��hRR����.�\��J�'L^-�`#�A&�,�i��RXk[Mu�0gա�Cq�+%5Ϯ�/m�.��b�]�oRC�3�h�]��]]�BSE9�N:�d�ȕ+ѱu�;'m��u��ey���4n��f�8r�k�:E����qpg�qǁ��m�J�fbP�eƯSA�u�9:nW]�t�H��kg�]�[���J�F9 �� �f7\���D[�`-���n<��R
��jS˸�Fl�3 �\UBcT��%�vb�c(�fu�KW�d��\n#��nnŐ��ɻ,<]�cy;%���#�v1�ɗ��v������ŉ
g�3�.��ɚK�<]�t�76:X넌`�Z�h�*Ѧ���j�0�D�t���W:����v�c����6���Q2��qW�]p=,�;��Ez�ѵ��8#�I{a�J�����Vŗ�n����1��n���tt��X̺Xhu�׮��\\mP#"�q5�B�f���k���=;����mu(5 L9��0i�Cvh+f�8��n��M�0��cEc�\���䁠^M�q97�Jm���A�K-($�,f�A��@:���E�p��p'B])�d�f]���sf�%kl�Ibe�l!DKm,��[���CF�J5۷;k��{������l��Yzx���:�
v�-�& �H��+��XT�v]��)R�ؤ�K�������i��цy�{�!Gq�Vٚ����<�����Ʊ(�H8�A����������}�h�1=�-<��]X�(�����ِ�n�LVӓXL[����et��դ̛U��6��N�Q��ĮЙ\� ��k�♷mسF�
6%�p��[%�[0I�;%;�����T�$f�p 9&����L�C��Ar�ֺi@��@e�6�s]�#�����~��[߬~6esٔ ����e�'�x��y�7ܩ�)` �ݑ�\���2����@#� (Gn������ �#���u՗�����������n��������`�ƴ��q� k��CO�`2�H$�g��{�����s�~�
�b�(�窀D#�� ���F�(�8~�[C�-� <@x�@����,����g(}T���i25A�T��h?x����9���H���0��Uq�����#�_Y���bO�B�_8�)P���?p����@��� �]�XDp���?x�}B��?}d<w�C��ŝ?:;�ʉ�.��#����0\�ezrb$r�j0�uP�}�>�1�a���E�nM�c��D�t���}Z� e�UG�{���G�u <@�>���g.v�������r�� ��o�`���C�8a��&W�EE�F��{*	m�c�|:@�~&�� )t�,Q|G�#��C�K�k�B��=5{G���|]�����G�@ܙt#�����>��Ä}6�ڦ~��V����_xF��9ͯ�G�s�o�I��2"������ ;�My������Y���nP����@t�E�����`��5����~�p��@��? ��-綀e��<���?s3�����@D�����v N��!�p}�G�.Lhb8|�]�@����]�J6�n"o��@:~�q"G������P�@gᤑ�H�x����<=��O�}p��È�{b��v�X�����+��n��i�(��eC"w�g�~�{��Ϭ�I!j�ƀ�~h�"Rw��<~g�?|��o������S�<>7��D0��F��?���+6W.��)_��W�������x��]����31gc��՝��X��]�J�=Q�u��]�� 2rxTx�f��*��ן�Q�"�p��	_��ǳ�,�ib�fWҤ��~��?r�����ԗ]����G��&i=�.�Z��߄?Q�+_�B����A���Z�s�2�Q��3H���!��G���������}��pc�ϑ�_�#�Fs~���x�?q͑������>���}��� lC�;۵kﴎҢ>����&{�,����g���kﳉЈC��|g��+BÊ��|8}{�퟼F��`h er����=���	1Hd.�?�(������� rr��� 3���0���#�����G�#{�efT��}��̀9�d��D!����}� ,�H��aC�ٔ<B�~�C�~���~G�����;��k�@��?��x��Fv�Q��L��~�c�x�;D�}Z@g<-�����:~<)q�������U��G=>���|+P
~�1�{���Yn!K��@J���Z���9�.�(���/�K���W�P��� ����> Y� q��{�b��"0�}G�,p��6l`�����=}�5������:q�|}[Hv���1I�k��N{E85h��FK+�ţ�؅��Z]B� ��}�{{zb�#�Gi���(|;Q���}�m}D|/��G�~���A!�0�]C��ր�>����1��`�(�hD�EOѽ����z����]��;��{�S���;؁�v���^[Q?�<,��x�#�;u9ܾc�B���Gx�~?B7(gfV�Ю�+��e�@�O�;V�ȏ��?z{�_
��� �DIa��W�0p��f�pL�h�K��G�}�b,GӼ�����!;���D�Z�Lt����uu�ǍmҳK���6�W�u������f3����տ�8�]�w��LF�r��$t���?g��>k�~G��^P����|�q��Fxq���������A��G�@5L,�þ�����F\�5�\X�������L����7x!�f�5I����|�/���9���@G����?3���_}�_
G{�Yx���X����v���1� �9�@x�H�O������=����Т f� ������?C�OW=�pu���^�DlFa��#�tV����3�?3�ͯ�?i �v}�>���:~��wʕ�g�C���8@ѣ������AF�l��C襳y�D�b�D@�*˨Y
�`?���T}��/LS��T����(M��l$���h�(h�;�9x��|���&�q^U�8:�C-BcF"ˈF8t,tte͸�I���^0&���n"E�l�ς g}�@#���B �}a��>�����Q���"l���GhU5R>�G���h���s;u�w6��
;�Ԇ����c�+�g�=��#�$4�;�}�����F��d`6��C�Q_h_c����4����F"8F��\���Z��#�=?F��F�.�2��2]�>�לY��}Ϗ�H�\ʢ�~��u2��@�bȢ9HcP�x��7{���~���ġ}��^o�2!�i�H�W��Hʮ�{Ϭ��Ei��σ?,�t�>���,���>�B||��G̥����� ���,�����!��s���BL�H�Z w�"�/�(���!G��y��V��C�U����p��	64]s�+���xQX(>�Wp�n1�oZʼ"���K�E�jI��Xb$x��f�aۢQ���T��Ћr��s�k�h�-��A��m�H��Gb������L���K�^�9sWnV��à�^�E���i����whll����M��)����d�� �:��,�Xx�,F�핤�\����S ��Vܶͭn4��H�L2�3ZZ�	�ia��"�+3����%�b�}����{V��@�����!����e�e�Ĳҝi��Ϡ�@�N4���!�@g|�l�DR1��IN���'�bn���#������!��~�a�/h�kI4E�]�>�͉��Ǹ! va(#�V���O�bB�}�H���`�!��-?t� 'L}�����(" 0�x��V���_�=��o�vg5Z i&�ŝ@���"6g�}9s84��b4��������Y�� G�Q{P��8ңIv�B�e��-�˒Hِ�r����{J��q���N�t���)ͭ\v�{�����`}��BDxE���X�����������U��_vu��r�@�,��	o6��$��yo�&����c�~�	4!^��_!aɎ~˹��_Q�/�a+�՗�uB�,�����#+�8�3�KSy��l�H��8}���n�a���`�p�<"==����qq��7"Jp]��
:A�u�qS�/ž�v��W�v8�)�~9���E�6|==�Ẃ��t�,�`��" ��~�����ޔ��+�w�+���* �Y����w��8��2�������~\ZU�;^?i�/P�H(���rQ�#O�N��8�a���I =�G���U��% }������B(���U!8F�]�X~����	���N�B>�������^�+-D��v�yHqt�i�𲇗O�&[�k���?}���,�_7Ҿ�^�����3���(��pSng�7s�G�xtu�te>������`�-�g�t��4l��0{U�vit[t3����2��߉�i���uC�?y��.^�>:a��Փa�S���W��E���N�������mHW�?Qh��g���]�?s��secP�]��գ�=�{]��!��D��Im&�$|����>��ͽ����>���?�Cրd�\��G��kcǄ|��*���P���<@�Dm Ǿ��:7�eMԭ��p氆� BG�.�?c�X��lo]DI�����h����%��P���ç4!���h`�ӝ2�\���;�-W#��Q"��wlC�%����~�0��g)�����} �@�	��4zA"�?a2�Ca�8����&�Z�|'������x�}�`��5���^P&8��|4�?T_p�ʘP���S����/AjV�sT�R;T�O���b ��~c�p�~mG�N]����p 4�%��O��{%�`GK���#���f�"r����9N�Eh�?}s1��e����.��҉&�G
��g���9C���fE1J���{��3�AS{Ԩ
�o{�xb��4"0�"!�]���"�a���~���މ�_Wf�#ę7X� s��Cu�ʻ>�2��� s���U�~&ёHb2;���A�+��b�P~�l�]Yu�+D��X�p���5\ド�F����W�|/g�h����J'|Oמ��"��C�G��a��w�k��i�+HX��ˠ*�x��j��G�V�9e��&�Р��Ň;���0f�;d���Y<�������d"���_�R)���q�ݣP����4��X)I���n�t'��M��w�to6ol*�Ύ�H18�=�?(���J��:���ٰt��7_�7p3�5T�}���f(f�2=��T��=�P���H����럟�$p�׳�U֓TA���q"�����B,0x��^J��n7���U�F�����C��0r���p�8}�#0�Ι��Y��+�������O �Ƿ�Ɩ��8F�T~�@y�2/t�Ga8�p��B������C�i�{�p����1�A3+=�q���zxs�!Ļ�w�^\����/��t������{Z3=2Djţ�я �׽�^i:B�
i6u��{#پ�5��=�h�a���u=�p�-E���kFo*�?x�����xc�y��UN��JTLS���Ι�3���)�o=R�b���1 &��=����t��{�EpGC��zB6t�L�U/i�	�Y�$8�oe%6I�H�7@�-�0��֟5Q��g��-���u�%��v���}{��x��"&/E���(�#�o+�z.$:�G�"Q�� j��}BY�1?��������	�W�*3�7�@'�p
h������_�_x}齩���`���:>�]�]�u�U��(Fٍ����d���4�j���#��V�ɞ�,p��qzI�^���z�5xPa�d"�at���1��ܗ�yt
1�O�G�U�	�澛Y����X�����J�nc�G	��jr�ZhL�z�:!UJ����Փ�u�:��ge�.pB�@/UR'�wo��O�� ����ǹ�b��O��QB��;�@�#�mN��&�����Ѕx��|?g��������~ ��.�\�!�L�I��r��5�����N���f��E����������?d__��2m�����>@i>V�K�xp�neSJ��Z+o�Unoz��<��C�C�@�����uZ\�fV|�;`�u�y����M��;����~�Ԑ�=�=h�[�{v(���q��۳Ia�<���L��ʸ[��A�>���.���Fp�b		�P�50]�\i<X��0t� z��B�A�
w�L}Ś��i��q�#��X\W��g��;�+���^�y����uѸ�i�߯o����h~�0=)�>q��d�w�R��b����c�u�<8���/>~��댩>�ZI��`�U��V��ə������c��b<8��1��0�]{�c=km���ԏdͮ��
xD�����νh��:���NY�D��tiVϲ���e�o�vs ���=�����~�M5��HQ���s�c�� r�׽k�,̓>ޅ�\���#2Y��v��ͭEׯ�'rO� >���ד"��T,�D�!��ץЏ� Ļ�1"�$.[���ޗ%���`"���|�ۛ���C���kyw���b��	\�L��z���)�f��E����o wn�n�[��眊ڄ�]�IRJ�D*6I�,���J�����5N�ᩚ:ًXԥ�#�hK�q/6M�Y�v^��b	��Vn�iCGh@�4%�u%��.̤%qڭ��82�#f-q3�]�.v�aB�N�q�d���q<{7�{qύ�)6�Sq{�@i�e�HX�]�`�C� �v��A�ޞ�v��\��ٹIeq6�K]�HT�pZ�4!g��e���ݾ�!��c�Ѿ���]@$��x���\���}�3��u������m�&@ОE�_w�M�1��e�{ֵ�r��ዽx�|~���f̏�D:�z"C�O��ǖ��l�ûC�u%�s+v�$}�$}bGr�`-���8D(i����]�%���?c8�.%�E��W��_���=o��ߟ9֮�`���'�5�ζt�OA[bpF����%���Lf�v�i��N@�[���hj����?:?`��f{����"�Z'�ñV��];���S�n�s�G(	�%G*P'�0�f�=��^19e��{DÇƚ�=U\$�X�������2KY�E/sb>�0�Dy0n�*�����>�AG�+�[ӛ��.Cj��J��	W~�=C��0�gP�������)k���չ�",DpU����yú�Ց�l��m���R���� ��0�(�c����Fkݘy���C��/L�S� }����Z�z�;���@�¬���?{�O�`�B��O��QtJ}�����ꆊp�?��\7o�G扸y�ej���V>�ك������һ8ſuj�V��g���4�v�+(��Ԡr��VW�-��n
K���9�r��˺��
���8���.b�|7^"�KV��ɵO���v2�}�-1�g˚���<���5����2߈���9yt!Df�/AeO�fE6{<q��9jfe֚��=i0��i^�6:���.�M�"�
 ȥ[/U̚�ˈ�qaPI�sl�")�>PόE@�)}�}Gwk�{��1��q��=��b�I���k:fD�ދ��yP9��r�{�\!{&7��aH�&L��<F틒wާ����M(�"=r�o:�t�t�����@#js�v[����Z~�w_����y���n>�8�M-�];a(�(�P{»o���?f��B�);�f�O���K{ڦ<��#�X�U�[dx�5����>�O�����������\��UUGor:0&�2�@f�c�5��(p����![�/n�|/���x�������&:]9���й�1~6�����{j�'�l��Cq!�8L+���yz��3�r���ف����ا׎TL������G�=��^�+����bM�W["*.ۧ�Ⴗ�gr39�%��P�I�ٌr-��t�����
�=3�Y-`��*�<�LA����څ�t,��<W���7+q�o`qg=uTn����}}�k�[Ȋ���M%��a�'�O��'�3��ĸ�T<S��B�`����^��La*���qXg�@0�;U	�D��ӲH��uoiTfue����r������T��+%<�7�R��ňГ��}�tK�����W~Ԋ)4Zh���D�P�d?�^d�Vf�\R1������B� ��B. ���1���[�!��4�H���5��[�(�/8��/j���v �8	4-3 ���ʰ�)��V`NT��}+��7�s�n���d��ҿ_�)qh�+`���;({����J2������x�!�l�g��Y�AlL�@Zzg՘k�"�j:~�һ��C��=���Un��O޹��
oz�
��ND��=�s��s]^n�E�M��v^��0�w'��Gw�Vlt/W�N�k�;�e��S�Ta��ۨ���4R�ۤB�Xh����m�[;��y�lw��&��W�F�}}żɘ�C�{Y�	JE�*'����N�ܻ�7<�#���q��v���-|�(&gr�1o?I;C��6�Ϋ�Y��kW�H�KeWo{3ي.A�DaO�bFT,�����޾]E�N=�Y�N���ہ����(�,�1 g{0����EL��,�An����$��<�IO7����~o��;�3��t������'wN����|����t�<:_��$�wt���8�1<����t�y����N���&�wwwI%�����@��wN���'I�6wt�����Y�'I�ӻ�N��;��$[;�t��:w|���z����|��;�wN��I:I?q�=��/??��}�/O���~��W�������_�~?м������y��W�����y#���?!����?��{��t���w韆=����z��w}߫���:N�����)����^��������?)���?�~��w������ww}�{|T�����.����9�~3�w��~s�}_wée���I:pI�$�Ӹ���N��OI'N�A�e<3�����ϧwN����_�������Y��~��|�{w�_���}{��Ӥ���K>�����������zOi���w����������a�������Ӥ����H��B�'��/w���g��I't��޳���Ӥ������x����:wI�ӻ�����>:I;����#y�?oY�� X`�x!?�/�:�� m��8�t,�$zwt�;���/�?�ǧ��>~s���wt�;����O��?�}����O&|~3�zC��򟇺I|�ӻ�I��{|�Ry�?��O��t���ww^�>�i�}?���=�?_ߨ�
!#�0&����?v������xO>�{O��{{O���ӻ�I�ݧ��������t�޾�t�~>S�ǯ�_o������n��wt����|��=>��<O9�Ot���'wN��_�>��o��Fw��g����
�2��>�+��������9 ��>�p���IJ�JU!Tt0	* J��fXfZ�J��@�R�[3�*P((XCeV1%�D*�
��UI)���jJR�!)T�D

�Q*�>د�� �P@��   �     �9"���P��         (B��UT 
�9(K���� h��URHP
�j��Ph i�4� : ����hr ������������ {�]T�݅)�@dP
�tZ��=�z�f�+��B ��@  }�W%�ϩ5�9bɻa�Yf��޽���=w$����A�ʳ��٤�olz���Y5����{��u�6�ǽ��;Mm�aۉۮ��=S�F$u�.���Η���uݵ{v�9	��P5� ;E�eu�2�(�ڔ���@ק\�cml<�Ti�R�zv3US����Ekauv�N��:���X��x:s����� 㭯^��Gvd����1Փ�"�;�vQ�1m��wG��4U��J;2�J�"  ��ﯬ�,����N�N�]�t4)s��*�jUv����^�^׻� y���G$�96��f�wu�g����3U�٩ډ����k
�S��@�.m�N�]$�.�]âE

�I)PK]�ev���s����j���垽^�An��ov�P.�W1��:���ۆ�ݙ�4:',ׯ8ƅ�7t:V�T�����US��) Q%��U�b�   ��/=�9+�s���+���Ӈ-��vTü�N�+�[K���Qk7:�8t��j��[����#�+���ύ�hM9�kN��ַu.�]��U��
���mE*UTUO{ZW1�k��z��Җר�OUrƼ�4g]jf����S�v���W�u��rd�u7z�6�\�vs[�MRiM�.�Gv5�v�x/wz��1l��*D�z�  q��}�(M��g��vg�w��\��w���׽�����5�뷸v�=��Y�ͬӮ�9պB�h8w���[JV��k��-��]J�^��� DB�
T,5��::���3�k���c�\���U��Rzz�=��B�֌w�����zᲇEk^��M�{��觠:<�2��<�	E*A">�DG�  g*��t�ͧ�����p�e�ދ�Z��#u^�����E[�;�@�Tw�4Pk%s��uc]�u�x7�����aͶ h�o,kͥ��w�>�T"�P({j��S���J�   ?�bIJ� @ Og����P��T� JJ�   S��UI	�2i���*!%(��7�cF���#�����7g�����f�fN7�n�S����k�\���q$�KX���Zo�4����;�8��x}����8㻽8 ;����8�?�w �xwq��y�A��ww��;����www��qݜg�{d���o�w��	z������j�Γb@B7p�SP����y6%U���UTr��o^��Vѿ���V��[e#�a�Y�T���ySGvI��fҊKWw��X�E���N��3��m�A��o*���}Sj�CQݪ�5&�W�P������J�s���-D7l��d�CۭL&��GQ�P��%q$���V�� ;��Bm��,3\�7e�`4Э���R��t�ȊE�&�&׉U }�K'Jֹ�T�5x?V�%������&�"���$��{H��UN�@��M��pCo�%BXLG b��Ju�aI��8��F��E��AGuڷ��Z��0�0�5�y�X�z����/0P���ͼ&%�4D���hm�Wv,[�*��6�	T\�f�w31��;��t�+S]\���u�۷��W&TGnj
:zvR��Zc!�x7� u��i��*�SĨ���wE�iVJ�(Tj���0���w	�×Ym�X�_��'��{F]S$��~��pf�[���U���BrcN��O$25�V�YFT��p8��9��{� �X�K��6:�Ĭ����,�ɣoMh`)q�������j�j�v��A�a7��G����3N4���y��:̱�-^��&]�ݫ���N�Z���Ϧ�2���N����������L�ⷴ$X�P�ڊ� R�ݝ�/`��eX��d�צ�f�1S�J��z��a)�;ܐ*�q^�)�6E3�Fh٘Ee6��+ P��x��u�Ҭ3�����)��]-K��$eVք��TuKe��V#�4kcr��x�)p^l"�=��viz��{�cf���ASbJ���ͫK��̽��;E�z�5� Yw�QT�-�������b���
c�u�X(#$J�s~�0��.����ˎj�4�s��*�_�OX����M�C�c�gW��gN�53*��X��4��
3$X�T�	��6��.X �G3.��#i�;�����n�5R�m����%0ĩj�����i�l�ui���N�􂵊4��A:�V/Li�&2�P��V�푏Y�YR�33(�i1�b
Jׅ�@�FC�)��h��Ҟ�g�)��)��x�Ǐq_>=q޷OzQm仧WAUd\��钅����ȍ#���!�a��zs�F��D?�RG�D%[�">��C�Z��I��m���cb<�;9wW�i��kP��G�LZ�L��Kۂ���X�׭�V�6/i�
:��`��  @��q��ѳiㄽ�X�&Gkq�d-�t��/
�7#x+d�Q^�m�0�x��i՝���n�÷S2��Тvj��հ�cr���љJ�)����12աIVGy�n�o[�u�	T��
�F֩��U����qԂ�6^6M������b�x�Sj��;��n��LbZ�JQ:��Y�E��Ć�2��s2�'cv�+6��Hfe��l�ô�2��]C!�ƚ���B��QG��{��7P��!��l#J��[�cE�t��V<2��D<��	u�pE�gI�K�>�>��'� ��f�7�W[�u�LئYv�B 9�+a�7^ �f�EfE��t�m�ٔ�/t�r���h�����ɁIzIT�����VY7��`���vVZ)�6��@��m
[�kF�E^])hK��K�e����1mcćL<p�[������,6�i�Y@��i���؋{�l�Q�غl37��%N�.�.�L�[��f��R�����ˌ�� ��BGs'Q�oN�):[����n�n?��{)�� Wg]��5Uy����l��B�T?��f ����$���*�&le�%EǀԪDۻ�ܹ�;�LL��yG(��(�jӦ��w�r��Ov���ܧb��V��W�(�i<0[n�GkI.��N�Q�9�֝�T��VE-X/�+h�����mO��~�}�uu�}>�m�n_U�.S ��O�o�ܰ�3i��5-�����Y�6�jT0a���nE�l��F�}���*�6�e�P��7����QH|)8��8�}{��|N>�����q���8��d�����w|O�n��{�B
X���=O1M
[����[[��'9S�9�W�l�.S�/�7�G���/ͺ?g��O��w�|I M��t�b��*�P�W�<�k�Zk4�%=z��R�Ï �	q��B�{U�\��͡�n�T؎(��5�լՀ�Aj���S�d�թ2�+*ɛ�Sj�qފ�lM�2�(�B�0�f�.�=�M&�
$�Ѵ�Ɩ��y��|���U��{'p�
W�d��/���o�{����14�h��n�h�u�
�*�͗�dd�@��J��S4lD��2�zr,%3F»�BH]^��(@y�X
��b�m�X�dA�D����{s ���`dw���:��R�	�dvC�����Z2[&�h���Kkm�a`����,�G����k�)�F�9�/-�𷈬pǗ�t��d<J�w?3E,��G���|��R{Z�j�.��}�j����֢���һa7���tF��Z�;&�ޓt�Z.���T�l�^tf7���ih(�~˯�}�i��}����2|{���ǁ��/|Ud�<z��=�y��W�;�'
��}�Q �~ wFL���n��ʹ��mѺ4@G��+�R�*�n��L�V�@�Sl�ˋ?6)U����S'�'u�Uc���@����p	����vp,dMn�v�w	�M�����uIcD�w�&¾K@�ASyd��i�ض�z�#XGDk+p�����E��LͲ�J�An)�
E��)�M�B-Ժy�auf�kA"K���6VFƊZ�@�$e��N��N���[�S(m�ba���T�fT+.��K��L��F6��[vYu�8���"��f���tf�v)�Yc)��)��}+t�09R�=4h�,�m��o �Xyq��@\fB�kFhl-�0���;[M��5o�8�Ĭ��Z&�nAdCyY�rÊ��{Q���v
���l�3�ʐe�&��5��.���`�wV�ǚ-���#���TʼQj�Ra/Y�� ӥ�P�<�yASn��f%�j�Vj�m��B*�V�6�̈x���ӡ�%�
Ҩ#{�Ar'�i
�5�hRXn�����wW�U�&%c������ �R���e�7��ц��4,�@L��ےLch2�	S�2b���˘�ݫSrL�P<��1�4G��iC`�f��:��f�r}Z��$d7��uH��1�X��\��F��G��I��Α�%2*tv/��.��ѩ�E5��?XU���ZZgn=��d��[���q���g�����,G��:���0e���W�e�/5�r���&���V�
�%��`�e�0�%�k��^�h�M�D�v������4:�7_|#��m�^ﾝ��޼�+���E�<��w��^���{����^�'^��x������:-�~�>��h�>�� K�T`��T��ywa�iڟ�֘"�4nFU� jֱ%�Q۶P��c1Բ 2��43�c*ʚ܁԰�&�k��ͺ,�u�Ca �:Ouc/
��t�	x3c�Sf��ê�O2Č�Dh��lM
��{[�<�I]\(�M�Tm}`�̬�\˰�;�;Ψ*(�'0c.�d*)[�:1�)����"YzN]��K_f�j[;�l��4�Qʄj�(B�U�Y�UZjC��q9-%y��2���9�3[�Q���X��SЍ�q��;*�]�܄��j,:�r��+�V�45]kB<$��tʫ�v��x�8�#a�F~�NK�n6���lVń�9�چ`�M�I��k/Su6ln��v�^d��=&�l��c&mc%�[�6�7��u:⬥l��.��jd�"�uu�ͭ�%�N3�V�[ �/L�z����"�]�n`��Y�0���"f��nIo�F��9�[yMX��EV���r���х�(� H֭F�Y����͢2=x�
,^�$�)b��0�ͽ�!R�x[GJ�2-##*�Jw��p5C�QN�2�U��Ѧ�f��nds.k��d��`u�6��ip"D�"��l���u��tn��72�CnfEѠ1#�(�X�+h�6nk��Н��E�#U�\uV�6�:�n5{p�TZj*�:�ɑxŖ��cʆ)R�
��85$t@��`��;ǂ7�/%ɪ;X��:{���txU�G���z"��'IyH����G�{�y^D�y�8UA��S�@X�B<D"t��Q#A���˺�f�٪��Z��M�nĠ�Jq�ĞY3�^Լ��sV�q$K\Kp�̉� ���W�ˊc�%^!�t[�Rԑ�p��sV��9;�����Ւl�1-we[i��f-o6��m�j
	�ڵe��Q���(n��1-յ�Y���9���t�Z�����)$*ޫG��ww����ɂBB䧀8,�x�[OM�)J)����WY�M�:����5�R���M�WRP
����J�j#M�y0�7��gρ���q��T{��9�<�ܢ򈪢 �wk����{��P�ӂ�6�l�`������������U�`T�Ǹ^d����W�t�%�=����l�t2�1U^�D�{��}��P��g�^��~Bc05���Q�UTw2dr�gM���[r���^ۺ������Q+�[�O�J���Cl���z����f �8�5+�f�2��[hk���b6�ښ�5B�䂢��٩��V�Њ���:)n:��v��Ct�m+��B��{)}ph4uRss�<���G�Q�בl�ej����%ֶ�ꗺ���2����)Z�·�rk�c%�1�ٺ{L�aC\vu�/,[Djl��l�!�f0m�7V�Rz�ښr���e-���	1����
�1��+oE��BS� ���r����d�=��-���0?ud���ɠ��P��;��t�6U����,�asE�Z+��^�_)��ڨ՚䧶��ĩ��S��ֲ0,�On�d��)�R҄���Y�en�r�
4��"�n�u�Xue�Bf���ED���1+�H0��"-#ZE'7��"��uN����J��t��׭Ѹ]5�$���V=��{Hm��x�U��m���
q�j)F�v��ʓ4f�*��W�ll��eJ�[����햠�`�LQ�H�z�V��y���n����)U�`$e��]�{�Gz�7yslYqAN�B�;��[xZ�
�#P�vC�f���R��:�j��2ع�ҕ��;���~p�r�ͬA�ݓj�8��f]X�C`)�u�˹�"�6��-��Uw�{�u`6�b�f��Uy�.c�%aUiϲ�,E�ױ��&���Kh�c�Ḿ�U2J��0�!*�R���U2�2��ZΫY1����ٱ���a��^���	�VY��]K��IŚ��ʻv�ʕK6Ez�1�!*��eb̚������f]��*;�{�H�"����-�ڱ�`�E�y��UljMS+U;-&1�eev�L�Q��x%A����;����p�%�6��Z&O��Z�e�����¡��V��d�Y��V��KEŮ�������Ƚ����ګ��?�-@��M�e�i���Kҳt�T�*YwV\6����s�E@ܰ6�ը�Ù{�֤��-�-��EF��a)3	�ǋ����)b��ȾPۧ���$!jF'l����LöMm�M�[�r��t�N���ǳtt%f�e�<�"#�gUo��J`��@�pf�e��.=�e�nI�DEs^յ����t�c6H�*،Q<թͫ�f�[��#q"LرP%a���U�ܭZ5����ySd�^��q�i�����1X�I�B]�a�)��9h��A�;k�Ӹ)�U�4-��0�-�t�ơ���.��S�w�;��s
fԔ]:/f�oXH��RV�}��7xw�y�����Kڀ�� Źe��!�f$�����"��6cɪ�M��z�Vlq	jv�C�T�wV��Y��fj-�@ʧj�[ܺ*�Y��kp,�駙Zr�	����0��J��+Pm�nY��@"�S�e�̬U!�j���:/�Sy���nm���,�ܙ"���S��`��M`Vꂕ��ɲ��S�E�kw��`ҡ����c2��vv@[�Y&�7���E��h�cj�T��ʺ)e�*cZT� �"�V� �A�j�b-1)*�+[2��s���!<�㡘g�kBV,`Ј�k\��E
�t�an+�*`P�k���7#�5��
f���U9a�+��T�:9ͻ!0�؂ZZw���Y��tK��ffU*w.��qo�t��o�:i�zLm���@n�O1PVȻ$�ʎ�7��X ����y0�Uوȭ�C2�ኮ�5$nT���/A�F�(�iF�˶틷v)�w�#h��͛tQ7y(Q�oAf��Z�
�o�K*<��v�b��42�h�*��}�^w˽+^( I  7K2Y,E� ��  ۚ�vP-� Ż�m[km�k$-�w@   n�yL��][w&����9��E�!�	����ݜMr.��ϬL�GӇ��Yµ��6�4�ұ�u�	Ŏzb�3v^!�/�"�[�_�����s�J/CT�Gy�ܕ�� !�}�D���孑�дi���X���
/k����28n�N�G������o=�7����Q��f�7,�cS����8���}�"{�^	�� ����}@�Zn��"Cw�����Pv!��c=V���Vp���j�\�|j���w�s��^�/��o�SkC��Z�ٺ�U��EՆ��y����]h�"Q���5�;VO�x�+�_Z-�ǡ��2�M��M�X�H#:�4]+y�R��ڝ�K�p3k8JKo�9��J�T�6�0�0��6D���%�8Gŉ����V+6�+#���1�س�0���9��p�Ю���n��;R��֫���\��v[1��1v��Έ��v]�� �of2�B��aa�4��*���F��5�XX��C5U���U�Y�r��T꽸�UuCQ�u8\�ĽG_s7.�B�9�M�S�T�>u,U�C(]���aଛ4�tV�'�g�'� <���1H�l����yۗƭ\��)��51��;V�t���.wZӇ��IwRG�I���F���d��I�N�.n�=t/%	�v	�H���r��9(�2r�j,4���×Dm���5�^69���MWE��׼0��TF�0V>�`�4�5��;����]MĪ�u>��
��ް�ӯFUVR3��e��d�$kzQ�Yn�^Ǜ)�b2!�â��(�ܢF�\�$���6�;tF���-��sz�]tT\L]]�w�18N�9׿���)�헇s���1f�R��"U0�ńWJ�js-WV���#�Ӧ�W8�<+��0J�[��)�;1{C��z�n����sp�60�tX�V4����sL�H�5�Hsz����v�7%�E�����z���NK�T��6�/�s&*�My����ʈ�):r�/#G�go��YӔuj����\�9�Y�h8��R�;��B��8��)ý�6TӇ�-/8N�s�O�RsFf�d{/2K���̛�;�62
p��R�:w���5Ǆ�)7|�-�q]�f��J�
�^W�Why@=�Wrj<6V?��FGד;fλg^f��<wM���S^�z�9u�t�<��,�\�5�)ER�z���P�*&��u�����qچ�BC�NT�u�|��x�+EU*Z��Nہ�Kwx�K�95��v���{U��r���W)'�Z�Q�*�t�g���Kp̧ϯZuztN�N��I��=����P�&2�n��u����I��W]�t��[{߹Ts��}S��JhQ�ߗW%J�n7=s7#�c"���T�]�1���nk��������E�I�/
ް�]	�Y�
�q}��l�q�œ}�|�e��,`j��R�����mЙ�����(��ŴCuYז�t���;wf�&S�2�֮��V/�뾸���rvP�+	Uj�u.m/>��\j���!��n��F�[�&Ca	7l܀ж���pjn�M^Ku��b�ر;���K���p�>�uO�*(���؍�9o�����S��y'ĳ�7$�4����6�7@�%�.V�TC[22�V�(��ɖX�ƄoYa9����(��u���,���b�!��t�JU�Q5c9���`���KH<�¨�j�MVN���a�y3}^c�b�cA�?m�k*e�U�&I |�	x�UY�=,�2�2k/�w�\�B�]���ɼcE9��T�3��LΗ%�������]ʻ;.Ys`������oOU��u� ����F˛"5�m�~��%E�f'�z����~w&#$1��\Li"�:JJ޻ڵZzQ�L��
W0�Oe�yu��52�9��,�\�E�bI�^D��%3��e�뚩ue�#��f�B*�i��Q���Eyd�"=��7�^'��y�˝�}�]�n��40P���6	�8q6|���FW(��7R�c�1Y^>��5�u��K��v���H5*9,�5tB�אn;��Ǫ��l��v�Jd���[Xz�S,��N�**��K�/�VJ�V�H��S�n� [�|A�H���˖yb��Z��[�F�2�TP�6k�/�s�Y�`�����;r����۫ǐKhSJ؇�m�M���U���6Z�{X��A�ޛ�o��ъ�x�d�	�6�a5�S�vx,�$_1���ʱw��W��TR����n���k;b
�2�x�z�w�V���"ѻ˫V���)� yz��B�L�B�@��}:�_�Z�g9S�Ŧi��n`��*����2��B�۟�R��*7���$8ot˛x(�ܖ�P����H��Em�	*II����AkrJZ�y�m�D-��*be�)]��Vyi�l<�u^��髤ktz̃��*�4���oym��T�k9��Ȣ3�$t��O��}�k!4~�������p�s@�E6��?XWڦ�a?nT�e �l+ڐ]�+36
����*a�ƛu�P�3p^�%hZ��M �6Mۺ��!Q!��W5��O:%�Y]tU&O�I�8J����.����s[�/����-!���'�Td��ݲ�(�:�P�P+�D�e*(G���WƙJ��/�c�	n��f����--ƫ���d�~�	h��U���4�)�Ηԝ�d���]�t�1 ā��G92	��gک�C% cv��j�R�dɡT�������&�T!+4����څ(&�2����Q�l���L���oU��M3����7��2����@Q��a�����@�0>��4�v�-$�qEr4��
���t��Qp:3ۻ�V�[�!EJ���j����dq�6�1D�A��A�����*�0ӆab$e`���yW�=��b�m�ٻ2��x�ª	��m����D��:"����c��K�$BD��`:��*����"rE���.��l�G�)
I�(��NX��y��h�(*@���T�⮪B\��Є0QƲ3|	Oq�����7��$��Fs�sTa�[$������<��z���>��<n,�\�R�gW�M ��q$a2]m�&���h[z�l�+w���A��_�l�4iko�2�\I��>/�l�����'��Ť��ItM���[[5uX�R��f�)%�a�����3;%��ڦn������?dCF���F�$RI�WUBL4R����T���m:ХҺM���Gő�-%�ɨ�fԵ(C2B�íU�޷��e�Ra��B��2���MK`�Hf�+b��)�";YaZȷ�8h1e�R�蒤��I��ec!>��k�߾D=�;mD4��v��#�u���Z�K�2�i�mz@�s��]�M=|q<��E�� R)�l֤�R�$�6ڶ�	eE���_G�t�Yv���՚^b�L���t�v�U�Ֆb�[k�T��XR��mڦ��r�TˊkJ�Mqh�3u�J٘�uw��3�fM��T�IҗMp�١e"[ٶ�HMyn��F�9e�+���݈���F�f�2�fM։��5�t,!m�79�y��$�M��5ԭ�7����������R�c�c�bd�$�f��d6Փ��y�O:����m���7��KۢuF�1���<-�i-�-������%�����&�ĵ\B�%�+�O���捜�p����Lb��,֚��;E�6�e��V��l˰\,$�I4�պͶ�bc;72n���f.�Y�����D��5eХ��,f�f�YQ�]%��T�Q�Y-�4n�-ý��Z޾$��[���m#)������'��|���f�bk~�� �� �$ce�\|��|#)�K&�u!]���ceu.&���Ke�q�BhbY	�-����';�Su�D�:�*��I+m[�6MaK*��ksJmt�(^��\�KkI	�X�V%�e#3�6	�5�&���|���t|�I�գ��	�X�I����i�d�A�d���%�ŗ�ce�&%uƛd�n-��jQ�8�cR�)46������չ$%й��ڷR�e5��%�!B�3"�#y#TED��D�Us־ȴ٣3bB+̆�XK��<"7��ջ�͊�f!"�8��7BKua�l$�T���&1�.����䏝�4!{3�<���ݝ�Ӟ�tʤ��YE'+5�Q�I45��vr�.5����2�J[��|��R72͵�%2Hmk�l+2lfjk�.�ݒ�:$�G\F�cmn�\�!v(Iu�ڲ�[R$6�� �3K���>�[كZYd�o2
R�5�K���Z1Wj���Վ��Y̺�,.^��FE�����H��&��z��MDY!m�4�`�f��,+V�N`�k$��cnl-d��>s�x�Յ��9˙�;F�t�"�b�l���[3�	sk�`�.�^����+<��d�Z�ͻ8UФ(��R��U��:�K�Jd��K�,%�J����Mi]uͨ����Ɩ1el[uGFK:��h�s�]�5�CDKm���,���jś:Z���h�	6��"HM��[�����LJ����3Kͮɚ0�H���]$���Ǯ�Zb�L�n�[[�I%���Xʍ�[��m�tƷ1��@�3�H�餬��][R�[�����������.�.j����WVh��IlHSj��Ŷ�e�Z�)ir��ݴ�厗h:	[uu�F��U���LBZI]6VԝF��Y�&Y�#e�c%%\L��r�lس:0uf%׶�n%-�6l�=���2�R�*C8vc�޶9t�%�H9�Ch�T��ƃk��m3+������8�]�,�Q#u���7lݱ���Vy�&/L������jY"Yt�VY0A�ń�0e�ua�ι���A�)5���m�K+]L��cl4ٖlɌi)���]��[n1,�k�6	�1-�Y�Y� ��R�-q]�HI.�-������,�h��(���c7+�m*����m6�l���ɵ�.*���*p6��!�6��i��V����K��;X��utΒͺgM(���£�GC[��Ľ]&f�nZܣ5R�h��W,]�[cj:f�ԗ$,�D�-Σ�$�,�gf�9Mdm�̢\Nd�u���:����ƶɰms�d�sld���������i��m�. ���%��4��)�q6�Y#e���\l[���іc/Xk2%��KGiu���[p��&ѣ�-��mFP                              I$�d��:�h�d�2�<VgA���f��;_5�_c�-���e/�wIgV`�Q�#�,�Xb-�u쨷�H{tN�vr���S�\�X���X]ݫm#���.���Ap�NCnN.�MK��/���I����/3528��m��5��o�Ū�0R4�S�q3�PBoR�I-mJ�˼�:�^�<��:u�}+�)����N�{)���в�)z(ic�N�#W/(����h笸!;���g3��G��n�:���hXYu��p����.�2�j�<�ew1�ʾCF����ե�S�5j�]x�.u�X�R�ȼ�ê<�w�Z�Q�i�.�*(�w`5y���R�p85�GT�K1�Kkv������l%b=�ՠ"��>}Y{�E'V��z �Ŀt�ڵ{:����D�j�3Ķ�oVۼ�k�W�5K�U0s���v�3m��:ا��з1�[D����6b�S�f�L�e9Zh�ʾ�������W3����*R���ts�p���Sr�j�.�]s���%J![ۊf�����r�(�]_D���0�\a�c<�ؙ��۔1s�5��uZ�̾
��ᷴ��0.���N3L����F��V+`)�B�0lX��7oy�S6�/�n��u���JfJpEN5x3�z�a�C� ����,��Tַ;9�����_)�GlC�j����V�;��R�[Z�gQ�YD�/(����	��ɵw&Ȅ1��8gi�飴=�8-�t�+feQN�u7���)XL�z����޸0T��p1�%[�y�f�t?�Z;�낒�-�]v���r������,"�����omߢ��?&�HuV�� �yrV�P^�ٗ&�pv��Lgj��h���tI�7�D2���pI�A�� iݷd(����w�9vWB�`�0h�X�W{&�
��;̉!��E�=S����'����C�?V����ۀ;�;�����ww��^�8��q�w�;������ߧw����q�����N;��^��wǸ�88���S�%������wW�:��q�$���q����8��w�z��D� P�����|B���_�@�{��x�A{���C��w��<��T��<x^���1�����)S�,��~C��T���<}{����EϿ`}{�S�l*uL�EAT�z�wW���z�<�P�ߓ���8�|N>��|ӏ�8<x��^<OS������{ǃ<��x�/w�� #�"w/H����T�q�N�!�;�}yx���q����N���?'m��^�'G�+�x�'.N��'����^螢�@OIǯ��=�wd	�ꂜ����=C�{;�;����><�|x�L������x�{�'��z��=�;��p�޽�G��z���|x���^><Xz�S�����N><T�{�� ~�� ����2w~?y����wq*g���C�^��?��U���l8#'tC<w��w�2p'G��w�'z�Oӏ��礇u{�juN�!�蜡��=����w����/����<y�
����ǈ���?t��t{��8;<_�S�y������G�di mf�,�k�|��S_|���{ϓ��ܽ���!�{��^�����x��;!�yN~�;׼x��~C�w���x��x=yx�6�@>'x�w�
�;=�\�^�{���OS��:�T�}{��px�2�S�x�;�x��8���C��+�wǣ���\��=�{����W���^�� �q��"w-�/D�w�'�ow�zyi��z�ǏG���E;�I����'d�������}C=�� a���T9C�����/ ~H�z�vT���|O�������^<�;�(~B=�����gwD��vxS�����wx�G��Q ����'�ww�w)���N����'׻�c��><~@�����^�w��S��|{�w��>�^�N���w�;���D<{��^����|N;�y}B�;�������C�����=x?<z�������'~O�
}y�8��� ��z�P����aǯ~x: �������~Ӹ��ﳃ�����;��C������ޡ�w��x�w�<{~��
��w�����P>��;!ߒ!�<N��+ݐ������g��{��vC��^;׾!��|N��w���~@��r���9x�=k�ߐ�^�z�O>�>"�W������8��y!�.{��:�27� ~@��~C��xS����^<x^S�'d��/��w�iǶ(��P�y�;�v@#�x��N+ǖz�z�y'wx��|C��C�r���C�����
�x���Pd
��y>�W��w_��=���)��W�7���>�Q{��p|��t�|N�}H�||N��M�q_-ی��纡��p}�������^����޼w���=x���~�8�'z�x�G����?{;� ��G��w�����������}T�w��<�|x��Q{���p}x��z��C��ߥ>N��W�x*��g�=�þ'�[8�&x���S�'�@��Sעw��gǻ׃��ǽ�w>�/��ҟP��x����=������0 mC�Z�,���4����4�����?X��wǻǺ<G=����N��N<���^�>!�5gǷ�N��ԏq������d"!񈮞y�9�˩��7�����}п�w�u�9|z�(QN����^S���}|C�����^�u�u{�<T6���̑�x�Cϰ���O�~z��{���޿�y���ݓ�>=������!��>�����|x���]�����g����@����l��gH�������G�F�:<~��6E�e�>!G��^��o/w�~hx�@���g�/Ӿ����~N���D�rǼN����~���P�>C����c�{�����`�,�X���;��ē��K�*@�����+��D���^��q�x#�|$���OI~��ڱ{=Ǩx�k���}�dGǏ�d���2z?�+ܡ��>*];Ƽw�x�xC�ꞿ=�{�=ާ���|k�=^���o���g��|���w����ȿ�O�!�|��but�}�y����`�� x}�����g��@�q��Y�g=�|,�d
�f4G�z���q��P�#�q?@��S�#[${�*O'����}�"D�x��q�����'?OSHx��J��D?'���� �^��c�^�x��i��Z�?s\i���}��h�	H;'�y��P��������D���;%E�r�Bax�d�����ǭ`��ߢ�'i�<�����]<4@��<F��+��|�9�+����z�{��ǆ�R<��@�x�G��@U��.�Ď}�*}�~8��8���]x����?<|����_��?=�,�Q�>��ޓ��߾�>Oϓ�pM�|���W�I��>|'>��Ht|x�ʆC{ �<O��������{ǎ}�w��'���d �W��^��|@�����
w��;��;�=�T��jø���"�^�D�����ߟ��֕����8��|{�������={�^��||��=N3��|H��<{��`x��=ݕ�8�<�
�׊���N���^��~{�hu��|x���P7�iߓ��i��z �>1�a=�	��(8~���h3�L,>X_-j�1��O����>�����w�ww��������o��G���`�̕C�7>�O�o*��e�n���u���J��+�0��nD3��;2��ml��ǁЬ�8�%ihf�}��5�����"
��lN�����p�rf���姡���gU��\�n����]��yg.Ā��'t\"0�.׵:ސ�U|6<]���J}�u��Ի��Վ���ؔ��x���r�:�v:z�!up���/��s׭M=g�����7��\ha����GCrZ/֢��Y"��j!�.��Ц��7;n��H�o�������u����=8�qff[�(`&jm��;닂�}���N�s,Q��6�\��:
Z�n����}��˼?����;����@8���Ā>�`_�n:���~��{OrV�����{v5a�%���vT=]�p�.���w*�X��G�}�'��~N:�� �wt��㈟��!�}@:'q����?S��׸���q� �P��㈝����w��{��x����{�^��^�w��'dS��'o!�^��A�ں�or��
w=��H �~ ~%����"�������?Ӻ
�|g�	��ޱ�EUUU�UPD_'Nl(�(���A{Bp"}���{1~R�y�������>�AE��ATUQ^H�/�Q�Z�=�FΜ�<䜨�9�TQ�# ��DD������U�y�W�$�EDA���"��<{�!�/<��z"�����"�sX*������DUy��^���쨪&�*��������w��UR"3�TyΜ(��?͇�%,��3GL"w��qz|'�ʫ����N�z�������U��qQ�QsG�bG�}���6T�M#�DN���q∈�/<���AU��x�EWI¾1EU��d�J���^�{��:�>C���������A�W�ЩDT_��.O!������U�݇�W�w�<?���?�����$S+���A�����ڌ�lI�QG�Z�'�T�	񜨨��~��"��-�s<��*�,��`Ш���Q�U�hE�@���W�����S��!"5����N�+�緩O���؏��!(�DZ�D�����ygz��4� D�Q�??��I����]nX�V>�_ʕ�W�%��'UA��U�O��D�U�#�?��u���yAy��0" :~j�;�g7�}��֚�=	�$"�Dy�|��<�g����T+8F3疪&��L�DG�� ��<��ƚ@E+r���Fm/��1�	H��m1-�c-$4e�f&-��	^�M��~D{��(�����K��u����Bȯ�^�w�I%�T�d&��I"���@�@}���'��:AO�P�dW��u�Co���������'�#>�={$�� ���^��9(� �WZdI��C�:4�s|A a�9R+i��sR����O|���zeT2}j~g����+����O u��E����#"���(�IB%*c��H��&��w�ћ���Hlo��zy����A�B
��TI6~/�����9T��`�~zu��,��uHe��̟=m���ћ�IX�p�����������W��cp�X|�J�>B-��߳�����HM�����`���%����\+zs�I&*h��������0��˫$�m y <���d�E%�*������dG�br3�םf�96��5�	�&��$Cs��U/Wd̫*�mI$4<�v��P&,�B�ŕ���F�NƠW�F���اĒ�8�,�B	�HK�,�j	g��6(�-�[�$$:M K"���w˒�^/\�T��}�v����C�+\{�/�M�$���Dce�Ïk��ҝ�Wq�5w>W�w�4��5N7&��s*�B-ʬXv�F9��㸚�t��}���}'��}3$o7��d`���JI;,\9fM�j2S]�Ʒ_�mF�����Yz��Kf5�(�Ys��ᛣtlڗ:���'��_�F6�X�����5܎њ�4�q�F��w?{�1�P+e@�ޕA����S@�;�w����'FE!}��H�?�����c�Z�U!`
&F���J�X��ϔ*ֿ���ӆ	�E�G��5H�⹥�I2+~H.K���l��uy��KZA,�e��`�ְ_d�}���������O�~H�O��s�����W��$�-t�Jʢ�V�������/���^*�WDOȌ}�����|3��
��'�'�Vz�O�A�l/��*2|�A"l�J����F�CKlb�9" �!6W�)4
��&U��D!EIR��,�I{�f7<[��k�szۥ�#d+,�Ɨm���a�I�G���*���h��R$A����/�/�m_U��QH�z�_�l�u&���� +�r+_S2�����	&���OZ��2�g�{U������X8Hܡg䭣�e$}�L"$���W�A�"/RB~�A�Y��f���^�G�M7�� )"HO�f�7��VȳZ�p_R����F/��>��5�J����e��?&Z�?F��
F��m<�bB?"Ƚ�s�39�=X���,ԋ@���� �i5�p"8�7ˍ�6r�1��Y�X{	����/��q��n�١ܵ�B��ӵ�k��~'�6Q�@�#��O��4���j"����RX��1}kY,��V~�0QC<c�?Umܤ�I��W�� �����Ϗ���.�ï��r�h�N�>"��t��l����w�R���唃u��A�!g�~E �^.ʮ����D �`3�K'c�B'�����m�FO��@�[V� �%��>]Ȳ�B~���O{�_f�3Mx���g�?+v�r�"�2;�Zg��HHYd�R�r�`�{<������������z�^�����p�Nop��qfo���4����:��^ۦeܣ���,=����io僩�e̯H���E����4���-u#}�aθ����/iΡ3+{b�Z���M���R��{ɭ��f+����I�kR��NeC���$����I�D����Gv����Ԣ��vD"� �
�C�����Ӑ��*�ؚ��� Z��l�?2�9f�a�[=b�5�Ti����s��Wm&idn2��Aߩ�_�7M���eN�2�HU4�
ػU��QӾ�,`��V��A
<XС(@��	ۙÂ�V�3����ƿ"�ϖ!d�����޶!�E���@z� A.�(�E��ģc���e|��oR�[@�W[�!e!��]�3�*��z���"7q�\P�|�e�0g@���:��j�$����è�,���V���Dl=u���c��?6y��N�=�&��Q,�~T��"5as�����uKm�4��ϼNd�����&�\��XR�Νm
�#��ZH洧� Ȫ��B���m�5�b;�r	�l�s���B���@�=z<�-O�V�Vz�N�c�����dqy!��@��V���y�9=�*{׺1P#�� � n�V��/��.�13gř�U�d4��71))��Kv?�R�f�R6yy�B�sBMbUa��U�:�m?*z������g��=/~M"M����mϮ�He�ŕ�rw��.�|U���eS��o$�Ž�:�#�W�����Ax�8!J2|���I��I���>B���=􄜣l0�
8j�4<�,�C*��|�A�����k�m>��AP�l��Y�F�q�(1�5,�ˌ�e!�w+?yY���K&��1�@�VݐG��t��:�5��J�!��j��S!��@(�Hm��PY��ׁ�*p,�],�9�[����K*;�,;7�E;%�%�ռ`�R�JڐkO��׸�Kz��=��u�r��*�i�9J5��'T�3��hm�p�l,.�P^y�Q������H0�[�:B-�ͧ.��6/���8�T��$��_i�<��ۻ?QX)`3�V��]|�ie{ϯ���.¤��D&F<�{uJ	�2ȉ&vϛ��Op�5���3��7Lɧ�(�VK;wdPE����Bm���-�b۱���<�`�B��1�F�O����l���0�<t�<���*@�����jK]+�v�7~tE�I�Al^��ũ�n]��Zv�%࿝M�9����9d�f��1����V�W���?|τ-W�70������4�n�T�߳Nq���&Ѭ�Q5��p�I�U�j�.F=~�~�	��<�|�Z�Fp�W�ܞE��XI|��P/L��ݼ�M�S�=�L���E���jE���%UO�g���4]D��%T�H�i �&Uk�XFe(.x-��t�E��e�fC�g.L�A���lZv�s)*F��U3
#�j ,�vw�&14��тa�P�L���2T����\J�*[�Y��9� ��_�z� �|ٴҌ�X�f]:Te&&e���/�b��*���A ��ו���Q�E�B^I�t��{��>�H,����[U�Q}qGw������W�N�ƚ����'[>O�`R�Wȋ@��sp��oы���S�u�L�#�$Ge�j��1�.�!%����J�2wf��A�OU��@䁔m�3��Ц�FD-i�Dg2�Z�J�u���P���5��/�7+��uA=R����>㍛����[����a'&���c�	q��������[����Z-�+�aޣٽ�u�9�ָ�C�K������=�����]���뒻]M�.� �N��0^�V\�]j���IWx_�� ����c��e� �VXE�AX�.
��+qa��^���^��1�O� �"u�9h����W����R���\���,�m��yۑ���e�W]j��O�K��B�>>�7���!9h9�xS��@��� �4([�Ɉ�4�h��<����$�.�_B7�(��V��dʐ��M^m?�[���=�㱒k[�U�t��������	,�J����n��Q?,�Q'�V?�)"�]�F���Tq�����znZ�u�	�e�n",Sc)���Oˈ㔯>f��7��k~�}V��ܞ��"|��@WSL�wVS�Ź=t�C-�Ah��j�2l[��K|��_����e~>A)�L��Ѿh��9�F��9�5r��`T�cb�]��$4������ۂV{\L9�S�HR���;!�=S��"�j	�-w���#G�e�Ԋ(c�p����r2HG4��ڻG@U9t,]m{wt�����P���QM��)�F�:C�,l��oxƴHUـ�dΕJ�ȧ]g^��	�z���=V��;{'�t#C�9���#�&�d*4������V#?��vAI��?]�
��c��E�(&Y���z�$�ҏ�X��y��7�i�A+�{]�[|/޵�Q��jB�3�4
:FM��N$D�>VK��=��ڧ����^ŝV��3���?��ȑ�z����,�����&���t�CP��G���v��[�T�)_p }X��������������1���<w׏���q����� ?<
ww�}]I��z//����@�;E� }�����~�ٶ�{�2��_�� 'u�2�{ӧ�7݊�ǹ��)�͊h5�05�ɤ0�A�	��A�df�&���F[�M"Jy/��Qy�g\�I#�K*��百6x$im!m�i	cZ�[���c��#<�����[4��I)k+�Iu��l����9�ui
�kUl�$�3����d�`�s��l_ņ�2�I�ե9��N���vĘ��0ԣb@ (cyy�3En���j�̕$�&����<B�&&�
�S�p�a�u�a͆0bI @����<r����k������u��.��I]:�1��{+��r���t�� �J��T�RfT���9��z�����^���"��Ȱ�greO�2	C7&�ovJ���|�W	C]$]%�ؤƔd�5�j�W-2�����~�u���3B���#CJ�K\�\G+��"c�PY���{�Pd�����^G��Bx�9Q�MP�����Φ~�l��Yt;F�va�B��f�4"Ǽԭ�~���ˤ��A	�k{��I�t ���I.�0Đ�(C
A�(<�.e�R���ݛv�B�	K��N��4�Թ���b͈ɶ�E�)]Ig�uJ֚Q�'m��j,z*�`��H��%
��*���q�U�S0PS�T::|E��N����fm�
)��r�x�dg�hl�5�a�(�n�t����m�'s��yq~2VIR�&��Žԝ�T��,�9����4ϗ���5��~��E�8erE�-M9fq<�"cm�h>���n�4L�5"�?��G�z�R�P�A	�j��Wue�	��5fmP2�C,����E
$%��o:ϳ�.�=Jh���h�����}�� B�w=��S�bS���x�S��M���dO��Q�x�XT�"�;h}�E���;���'����S����}� p~ �^�^{�o�%�����&����#+ڏ�,��y̗&���$F�K2�Y�Ga��N��]�]���ͽ�^��{�g4�3i��������]�߄^С�����c4U�[$bQ�O��O����>{k�<�̞H�+�^.�#ж`�O�n/u�{1JUS�����g���u�͂�nnӤlY�v������H���V���_+D�~��5����>b/�_X�R�)���_[�����n�䋻��+�7&m��2�oE5�^�<�x#	����-<lK�����!���V��1��*,g��V�+� 8��c�˕�6�=7b�����c�^B�N���||س6@&�P��;��ʪ䩧J�nJі{��'Ʊ�TNuߴ-�|��g�z�%pCFqgo�5��O�zCջ��E*$�U��㮉����#t���J遉�RL���͞~�=��ԩ�Byg/R�x��pv������'�(0Ea�?�i�ww9œ�+��5�&*5I��v% }���o̎�{^!�
���r�$�:d�M�G���N���e�QݢSD����ns*�p��Ɋ1����r�B� W�X��K�vK
�^4鍧>����e��U;(��o.]���Jy��oK��I[|:�d�/�O1�M+o޻�1/O�)Q'����à� ��H�5��V|Р��;�mm��Y���ku�Gk�tb��,����,ͻ&^ƻ9I��||��)��>��(��D=w��Zн'��e��3WQ:��PhH̭r2���Ry����]�0*7�O��� Y��"K�٣��)��N��#)�p��wkj�%U>���?}v��"��<Y��i��>�m��lW���p����:�b��U;��� | �#�Ԑ� ����h�,�Wh]��D�Q{O�i�f���	�,y��	dݾ�AC�^���Oxb�yfa�&�N�*C�:��u�+ʺ�c�����u�_×��Q��k��U����e)�՚�8.?.ˈٵ�F�0V�i���@�b�N���5(�c�rG�L�_��f���͵�X� �;|c�6��T5���!��j�=X�;]�T�:���ZEWѰ�坺V$//�n���A���zh{�雲ȵm%���K@զ�-�o���Q�P����ul��4h� ��i�P����<(���C<iȚ��;�\�48$�����.wE\���ȟZ��4:�e6�P�mq��j�Ѱ�=�޶+��S��<X���1���ߕb���AQ>\Yݻ����	�E�9� u�C�ޠ��\jFN���lXl�Z�zV���{L�N��i9׆QR%=��bGϺ�[���`�]s봨#J�20I
�M�<�b�N2���l�ד��	�����R�ӠM�;�@{T�g��A��;�QKL�}B}yH3[��?V,�G�UT��2�J��ШR�hƌ%l��e��i7e����=����8���&������!_������j���{��$Q��/DQ3���J����I{�$s�=EA.P)z�{��E��im��[!,a�e��1���}я��w��挩F��ybi�m�*uJa����P�1�K��cE��\^3��.���S�)�:�S f��g{��d�_��U:T�7�%�a�5�������������i�X�W��4��d�~�C�A��o���fΟ�2���>-�T�g6{�Y�wZ��Ý�NWx�nw��ʞh�o��krN���0��u�	�Iۻ�����F�Hy�ŷ�C,��ސj���g�2�5�&y}�B,��ؤ�s�EP��݄Wy�q�Vl���V���������K�p+i�U�S)ף�2W��>��Xj���:�6z�)���=�1RA�лیRF�@X��GoԷ,{αغ�d�G��xѷB�8�z���]{�k��6֋v�"�G�z�+2�4�V�*���%A}(,ܤd�ҍ��d��q�<�,"��܇���X�
�hOU�UT��_��f�B1iU&`J�Fg��U��0Ђ�h"�N4[�2�-�YH��lҖ�T�o�ǅ�d�1K��D��B%A���Y�S.ݢ�I�����N��AE�;Su��(ã�m�K�I;)���{������v�!�Գ�5x��CE�25���g���F�ŏ{fjQRSk�?a����I�t�n�N��&��`w��z�
�y�W1�,`�G^^)��W9�w;�RMlդq!yr�c
ܩ�,�eL�kv����¥s���7�n�!qlX�87��)�m�ˑU�/������A���.[���k�v�6��
��ԟ�r�=<�����-�vϐ��p	G�t�*�)����I94wk.���U�9��hþ����0�O9g���^R�_R�U�/q#�S}��kN�c�Zw�)ɐ|�m��Z 0[.���t[�ǿLSLnn_9'fi�e���>&h������[�(9w�X��W�h�(��)��[��\b[��W�y-@���ӟ7�ڟH
�(Q*�m��S#mY�`��ҷM+m�Y
A/]f��,K
i�]�U*Z��#�+��1�fo8�[
�]�\�q�`�i΂m!��y<)4�nI$�..����ꎎo��?�I�n޸���UUmG̺g�!���s��}��]Y�z�C�$wT���ba�3��ݭ��$�NjV��Q@�~�J<o4��o����Q��4���S&+2઺�ݛ��Ѽ���l�1YXN&<�b����^F;&=\�D���4����j�
��tT���C-�f|�^��B�z�YW����g�8��0���r:��	�]O'ޕS=�E�(�hg�V�r�\�7�M��TXDO�w���rS8[��<��{b��{�q����,����4UʌZش�E��EQڵ�Ӡn�$�|�5ޯYږs��%=�^�9�yR���Iks!B���!�']Cλ]�3~�=�极�1x�w��j(�N��u��t*÷몳'��7zK̗YGj���sF.q?�"?�Q��� ��}U]^�Tя��V�[�R�Q$;F%��*[/.��$�
��J���n?��f�;}!�i�E�m�=b�V�Yʸ�D���>\��XT׬U��g4I��8ꂺ�`ّ�T�N2(�-ۚv� W��?f������$��nR=s��h�.��.$)l��s�L��CO�6ݣ$�%O����>W�:N��:bI?\�$�4�X ]1Os�R��#����� �H��K&-�j�Ҩ���T��spDbW2�O����I^�}Y'�V�W:췬�Þ~�׮�p�YF�;�ƻI
.�����
3��o��,�ڝ}[:�����M^Q�U��8�Z;�]k����_,u�]�p���Z�ߵo��0Z�Ǻ��٢���IG�qӝf�svݷ���ie��ӷ�9���a`n��p���Ϟ�����|{��p)����I�Sü��i��1Z�f�8l��G�ݱ��a�L;!���f�v,MFS�;�00/S©��Q��u��˯�mܠ��IJ$�Ժ��k�,��H2�v�X��B>�3e��.�]d:��	7�A��bQ���TM��%�w��Q��搾�}1u��?�X;�5����Jח]��݉l�QZ���ds���כ1J��r\@t�7X���E���w;i��UJe���kc��P:���:�.���K�8�B���jI{S]˃��*��pqv�)����&��%%��x�\m���h�K8Y�iŸ������+0��������SP�ed��J��lb���t����q�8������m����a�X�]������\�i,�Ɍ�٘7���쯷��UEΜg�r[Zz�G��۵���|#��=�d�� SU7.�F_�#�^���j7D�$���rI�������a!XmWǗMt���*fY	wNY�dͺ;w{����igZXM��t#[���V�}�6ŭ��X�k���Fɥ�^P��5I%�Z�۾�t
]����%�z��"��Kdҹu:�?�̕��Q�gpRp���ɷ�&�yu�]�R�*���Nɛ��1�ޘ��od�N�"�sܠ��7}X5Ϫoׅ@��aDl�R�2�fkr��+w��yA��c�`Z�$@�<��(�\.��������9��_Y���WH�J5U:IVZ�	J�=����� ������Ö��`lإ/Y��|�o�y�_)<M���J��A	L"�f6(�abM-��e���wC2v,��Rb��	T��&��f�DP��fHYflИ�$�,�����Dݶv�F����Jk�Kfb�cr�e�E���U5,bȳ=6�4�>������X��c����%��6��5v�=:�I��sK(�J,�Ie��2�[��h�����O<�ʋ&iu������o�<�fA(���1�JG�aB�lA[6�[�'W�7\�1i[R˥�-1pi�D˞wH�s$I�! ���ɠ-�)�Hc0����)�[��[3uoIu������4�2El��Q�J�є��U-�t��R�`�r�I��l����3V$�g-Jٜe���m,k�K-���"��%���V��͜4��a�ͤ�t�:&l$���4�Eq+5!s��Z�-�L�8�d1"�E��Mf6�m(D�MJ�]��붻��#5�Ksv1����	��W68���kd"̲�    I*>�Dμ��]9��t�J�U�*�r�˻Θn3ͻ
��c\��t����62��U�}�2(�m�x��r�l�nF�V]�I��؞��}�����	�ƻ����/i��2�ͧ�Y��%���=Nk�7�y[������G��;�x��
/}T��9b+��/d�'����<&�?'���_��'�(y{����3��#�#�x���@q�'�Ȍ�_��_x�q}�� E������~[;������
������M���R�ͽV�#DB�#��#g�`��a&�d��H ����ƈ�b��"DU�n�2���u|i���M{��~J��0�A{�#�N�y�S�~��
�������x�DDW��O���:~��6�Șd}�O�a"tA>{��?���d��l�f�5Ѓ]��b�}g�4���Q~C���J���$��#��H��̀܇��B$�?y�S�?�w���O��6��T��!^��{�^��G��9�	]��.����
,�yD_u������(
Y}��ș�^6.�lHЭ��"�V@�Qc�"�j?1!�x�����2g�x"�?�{=��q^^PP����������������#�E�?��ЈG�w�K"��8�?6G̍#��J(����]P����}������޳�TuE��V,�H����0��K�@����-�`��,�2��ZE�����������$7�={�x�x䭶��������=BC��q��
�)����L"����"(�&r�H20�E�,��V��q�=s�=�O�( �}��C��fH@��h��~G��u*�H���;B�$}9
�F���I� �LZ��4���x@�*�1��g�@D'�3��<�O�vx���^��j��/���(Tc��FԞ��.߽ءε�Ǔ�|l�4����c�h��$=�-|���'�N �T���ާ���}C=����W�v�&���O�y��S��'ײw���5��!�̟P-��;���lx��z#��;���HXH�|I?}DuԠ�����1S���@$"�>� ���*ؼ��/�9@�¥N�>���=�"�����x\���:[AB�~��d2Om�*M{��������'}���N���!����
�G�1��#�$�H�<o�(��xI��@g�q��߳��𨅟�xy�"rF�������~��|i�LZI�}�����H%޵�Q30l2�x�)��?��������OSI��ǟ�<缾P�N���>B�ߏ+��NU@��H5]���lM߮�]���1&7]
ZX�k\;�\͉���������DrW=������R :�2}�{�=x�{����O�����0������qR<T��Ҳ��V��$	#��������G�J�O?����P���D�|C��#�?DDwN��<)K�̰���r�7i��tjK�m�2+�}�ǃ{���F��:�ϳVl�8v�ا�}a����O�{�3�)ܣ-��2��Ǌ ���HQۡ	��F_{�����^��^�g�T��z�E*M����z?$��}4�y�w��>=^^��P����px�2{?_�<�@S<d?�H�D��z�=����#�?[_Q'�> �{�M_[���p}��{�����m���^D��|N��R�a>�N<H��ֱ8�~N�����d��ϟ���<���|{��=�}����w_I���U�D�>[�Z��u���2,�"�2/��~�|�t{��T��0��O�׌���c!�`��x�'��G��{�D����W���7��)���T�˧ 	4~~�Z~�G�I `�ZvG�U�dID����{�O+�g�6���D`����x�Dh"a 0�����9��C _�p����@ "��������P�k�O�a��~@|���#��|�;�O���~��Ǆ���_�T����?|������0��"���ݹ�ύU%i��\������,��/�%OS�T�Oi����޽���_^��h�AH�������ޱ�2>C׋V��<��E
�C�z��ņ�!�QyJ��|T�]:��{���� F������̰���~��D�!d��t��l�5��S�(_��4��Pm �"���ڣ$"/P�^�8�(��?`T������䩄P"�?a'�>}���O���L��1��עg��行�m]����X�@d{�0��5t�A"�e ����GϿ[��d^����J�{�a�>K������O�Z���?���<��:'��G�HC?"9!�i@��4(�/?p~�%q�?u ������#ֿ����>F��~4�����ȳC�t��O�~�7���Qx�	f����J�4�	�ě�Hğ!q!�UL�������?����~L�����&�����׃�'tN��D�$Ӿ=���z����(��z��C����6�W�j=��G�)⽯��H����a^�@�O�t���v(�D ��{���3zTIU�Sui���i��G��1����(�,��!�a��>�#� ��{�������>o�ǉ�;������?i����O�U��N��?�����|NS5�Tc޵2���46�g� 2����?T�^u.��6k����08��(�9Cdb@#dD�L�[�����O��q�9*)���g�~��g�L8���DY�c�]}�)�d��3��Ǽ���C�����9b�È��PD� Qt�?x��ʺ�GȍN�dVT^WT�u?bLI�0-
�LP�r�^*��k2;5�#�̧���
";��l�E=�ـ���u�pP�AKkp�����!�O�qu���x�u�]�uj��X�ӸiB��b[S�.c�G�h]�"Ȩ��﬌�$��,��<����~�OSH
t{��Ax�z�'����^"T�<O��q�O�|�	�3����,�Y���R��?9 <FB#�ȋ"���=8G�C#���
�`�\�p�4�F���4�$i���*}L�S��:X���EG�u���(�V`�C���@E�Ä��"��z��DY��� :\	�2x�a�ZG�ݼ�����~'��y�X�}�������2G�x��楱XH�4gl��c�ō~��~�?}�ɞ>���,������O��1J��w�pi�D�"��S�}�����)���������?	��9�2��A�L|f?�K�'�) I��#<��!w�zC�!�5�Ad�1n#�Nd�����mڲ�3[,	�8I:�ua�����s�wr���sHzR=W�bGB��rE����	G���C��ix)o:��o՘����
&*�m]�����!d��B�w�/(�=�^�b�>�pt�U�ߣw�Ax�����*��yD�Godȑ%4��5�l�җ�J���2�b^�7��=]��LM����5���1G
�P:��P���9EOo�ڭlmD��B���ê:�v��mq0���w��z�+�W��F�?pM3�	3�-�)��	X�kE&�/�)���5~&ޜ���N]E0�S�)_(�u�dG:����]8ʺ��5 �T�ˊHH�	�D�:f�|2���^�y��F�^wŵݿuZ�'�H�/���hV)v�J���;�|���Wg�LH@���*~���!1���-�����W2�F�6VQș`0����E���r�c�����tZ�j��7U��Ä�8�r=�W�ŝv�8��j͔Y?��U�'�t���Ns�߮� �Z��e������U^��P)��<�!X����ؑ�Nb�@��(E���2eY	~����Y�$b�&�ݧ!d^�C;hQ�歌�p����vܡp��shn�h딙�6�_^4�jﲡ��2;7��K2ifm�I,�0�Դ�=���Nev%������F������W̏�Y1.%Y&�vm���R[]�IGK��s�M�A�gc\f)!�Jh���A��H�x�]vx��w��4� �i��lȰ���E,s7i��a��q9�,&0n�]�5H�j#ӇRh�$,x&NM���[��Y^��-߇<�f�}w�j�q┲��M�,�
�=����R�bV'L���sPK��EW���\����\u�{�����uAQD�S�ܙ˴��GS6�f��_}� 5��A���ש=��MNs-v�N�VVK�S>�T*Z�W;��
7�D�d i�L����$a!!����!�ڪ�S_j�-�s���s\����:m��[~RS��9�0ߺ���j��@�͘p�]VJ����q�41�A�o+]���}-�9�ю�p��R�0�g��p%�8���P���T�Sh"
���]4�j$?�x^�͘`F�z�(ڴ�o���g�qJ�4�)�������w��T����.�
�H��鬀lȖգQZ/v~�9��AϪ��:��� �
�'"zrˠpЫ6A���Z�xx~aB��b��~�)� �l1�\�=QV3��1Xy��O����� �d�E�E��l��9��Rm���k���x����W��5\� a���鍚�m=m�x�����!��Hh�x��q�y�1��):E����$\32�G��HTߒ����v!	���:��ևl{�w���v��ZHj�.6��`�����띵]Gw���0��1�H�O��4zi U0{R�%���}��'���(���=F{��3~�W���踿=�sr��'���S�Y٣��aW5�]QUֆ�/���R�'v�U3�SjŊ��u��wNBc#T�0��Q��mq3^�hu|�W1%εk��ۤ�OE�kr�_����QPi����P�N��\�ݙQ ��������0�Orl�m�l���!�]�=��5�4�#���1^�N�dLJ���dQ՛�ǔ�IB��j2I��t���iK��.mF����ڵU����+��E!��,���)U�K綜�9#���N\ϗ���&KB�?���j}�GRKݥQ�b="4�k"Z� ql�2i^�}�$
�����<�Z�5=M�&<�w��K7������eZ������k����W�H���35�ʍKjr����W�32��!�p�T9�Ֆ���v�p��"v������/W\yl�m���qg¤��М����0p�Ϯ�l���	�Е3O���H��(ʐ����Ñ�?h��z|�Y�S5��O�!�4���0aOf��^N&Ź�K��W��뽞��Q&kw2��Aj�5�}UV"�D����
4�� 3PP�'�R`���L� ��Mq�\7���T�$��hI���{�TN�Nf6'z�����7T!��("�z��bzsT���.��'U���@a����.4j�6l���'*��
�uX^�zl#�~Pֆ�D�M�W�"���8�L�*�yST����5��)�D%����f��9쪞�ﬨ�U��|f�W
gp4ηc�~~H,�&|�ܾ��)몚1�[�UH�9��M�R&��\Wp�{Q��<@�l�őO��Mr��TF�A�TJ(�m6YNqY�ξ�s�
RWU������Ȫ����&�GR����7�\�����q���V�_	�^�m�����������{�ԧ�aۂko��2j���<�t��ȝ���x*r3�c7�cڝ6�pA�Up��`E�S�X��p�z�;��Gs�ƛ�;���Cf`ջ&F��R;��Xiܧe匌��yGl����v�7D���og'tvꣳ�H�M�{u�V[K}0�f�z��!S NM��;&�<�HAeB�+�y�lv�z ���X+��r&f~�M��E@�TI2I�-Ƨ�j�י�{T|���\mGIƞx�,�_\y��d�R�C�F�	�LQ��'���:e������/�oV���j�r{�Bo�Ѽ��������D�y��x�D*����B�_cXa�q��Q�wBh�Bo6��ԣ',- #f�NfuS�NZY���*���m<�sU鹫�;QT��j��4T�h{.}/�&s��c��ms{�SW�u�Ojn��u� ��6�'f$�j&�&��S�}�ۋi�,ϱj�j�VP:�?rT�.��*"1���|�a+�bD݊}T��K1�,�lI���>t�vo�bb��T���t+�ڢ����`�V�ɏ�E]�n�u&|{3-�����	��%;��>7��æٚ����Kj����I��8��C���%����ɧێH>/���ʤ4��nJ1u6�T���Y1�q;R[��v*T2�	�÷|��=3b�x�WIXu�K�H�~ںV������`/�0V��z�Q�<Ӹ��.�w��>Ǜ�!8���#�mE��[;��!2	cT�V��Mw�Ľ{��h0$��ʅ4h }��veg�+���\VOmG� #Iw��ɑQ���{�(9����J�$����Y�UB*�Cx��{��عU��৴y
B���1̤���%t7���s�D�VG��;�Ź�p*ǩ��N��K뵒%��I���L��JtA��#Xv��y��UA��]F��͓C%�R����k h:�}�J��f�^7���3Y��*c;$�TY���ȳ�Z��;CK�[����*]V�Kf]ʎM��s=i���Uo�fH�f��e�n�l�L��L�,B���w�M���)�����d>,ȐwXb�^P�����c��
�߽��+�&���
;����y�#N��h��W߫\��C^�EeZ�#3�� К���x���bA%B�X��>��`�F@���;%:����T_�|�)��01q(S����o�!�9p�lU�����<�cv�Ȁ/$�.c��g۾�<�ʡ���P>�^i&}��n�x�p��GI�yb�uN�X��ں�sU讵;��N�����������n1��7�0dZ0˄MLM����Bi�u��������^s���z���&���ʚ�UK{��1��e�����"�!>n`e( ��pZ$�jW��J[���nf�4�h�TZ���J4�j���}�C��k�9Yt���v��\l�P�UQ�z�"��9��m��t�V�����~��pMMUP1F��X����{'��6m����J��ل��]�c�j~e@Q�OJ��}�j�S�{���Ƞ��Y�x�oPrx,V�V���zg��2�QW��
b3����N�ir��0g�se8L�X�$vS�ƺ��4X��&_������ YN2��)׼�K�w��z�T�u�y�bjW�sR7�蟪1�Z_�Y��/���'�еP"r�X��j� �3��	D���Vl(Aob�{��uӒ�ፚ�y��Z�A�fw�_W�T7�}]=�>��会̅R�B�ͭNM�ɮ�oM�e�ûӦ���(5�V�e8���Kю*��eeK����[�Tg@`��l���Z�ޖ�꽖i� �mۢ�X� NX�d��n�`���f3LE�(�p8�k9�Ő���x��5����6X�%��,��GV*�$#n���,��Yw64��ittI��6ޓ�X��<��k�����L�#�(@A�J�I%�mWӱ�̩����)k�&�%}�K��[^Ț���s�on]��Β~�b�so���Zs��L2��^�������������/�(AT���S�`�>|$9&at'@'y@pe���&�IS��]�u6#�=QAx�S��}��dZ�cf�N�VsoאW�'��j��|N�'��of�+m6��\���F2߶Dٜ���3�v�@��Q�ʳ���.��X]i8��(�h�b�iֲP�,�Bbm�������Kbe\����l/�ר�wS�B�n�"Z\	�~�������$>(o��d�@���O:��vB5�5���}�_ 	������O�nd�q�a3�낼���*G���u�S���ת~�pfcK�|5ooeMxߓ��N1,�=��CX�F��SK;>s^��
�x��;HQ�E��#(����38F�����D����J��dտ�gdZ4���T��}P$�wo&'�9I\ysr_�JO�nr��KV�@�V�NQY;��EG�dˡf��BΗ�I�#Ɏ�h{^D�0 Ezk�՘UE��k4�e��{rױT�
���>�-<&�D��m�s�S�Q������ٿ\�p��V�XYxk'����,İS×N��N~I����%P�i����x�D���X���%�M-3�%�x��û���f�����׵ d��l�=�T���P멉n�}_8E��OSxW��;���]����T��"]d��spۧ;�mU��kȢ�5���#G֫���A@�ѽЃ�F����Ѥ&\�kzP�c��<�\�a�銅ݤ��wA����Dn��Ӏ����]�]LSB���X뤾}�f-{�Ju�<��¶��wJ��EF[��')+��?�:�_*��Z)X�}MyM��&2;��T�'��[S)������Ε3vW4��G����2�	fyݖ}�҄�D8&�ne|�)"6!����F6��Q]�]2>n�hR�pW������Lښ:�]��J^B{2�O�%Y5@�9�.�tz2t���\��xN���V����ᔄ�͎�������W�6�����T*�]0�I��� �LiN�&�W��:5����ų8�Z*{ާ4�����<�Kz�N��`�p*d�ͷ'�A�^�Č�����3)�%�����:��V����	M�T�U�%7����#��Y��OA�R�����6��Ϭy�4;r]E.nzuU��7�EQ��(p��s���뺙N��M[�޽��L/�/�O�u+��sh����"TBdt�'�A�T��W0'Y�дl��&��"�f�sj�w �Q��}V5C���]ȩ7�~���U/��gr�K���ſ��x��S �BN+����פz��hX���(c�6n�^��4�{��김Tf9��ДӁ��>���\�)(��%T(�s7%\O���I��E@=���D��0�����=뫚9�S񙙞�)|3�|��S��29�p$�÷�p��)�&d�A���/�^�r.��@����&��Q�F<�i�ڞL'+��&�(R��e�|�#�n2Ც=�0�r���`��2uy�9���6�p���H�������)�.WVbJ�zC3��i�ۋU���m�I:�$��q��p8V^�G�e7jgVA��W&C�(Y㏫�!�:�ӇN�Ѓ;n�4��'��z��՗��-���.�����k�LX����j�w³U#�w���|�y����L�O��U��K�`��(�UyĞ�W�n�K�Z���tdM�����N�=6_��A��m�ƽR\U�3S�۱a���
%�����ڴO�"��.I!c���˙�i�W���.4�R9F���q:81,��ӷ���{�#»�ǦUKb�MJ❞5�~���xU���М���f߳ԛ�x9����.�"�^|=�s�-�n����"��KeX���m���VɂwV?8(��T�!3ڠUa7�'|���$������r␡��Bj9{ĉ�"G]Mz}� ��Y�[�Y��G9@Υ14���Vz��C��	��� r�t��\j�:܋VpƏq��I�~ˠ鷮bɠ���4�Y�.AQ��mQ��-0F�&9��[����HA���	��ˏ_��i�|�u'���91{c��*���=�w�ㅷ��.��\,$HM�禮~�h����Y0��0m�xM�V��^��q*���IT;������.8�D��LNFa-� Q�$O�cn���T��s����W�ˋ9&gJ_�_ᐚ[Ò��sp�9~��6���OmuK�8ܻы�$B���1�4O���yi�1]V���,��eCϩ�Ў/�g��o�鷔U��G=�F�	U�S����a*�����F%��5�~�I�^�.e�N\�QU(�T9�X}��m�pG�7E�YpTH#Ք!�bhn{;[Y��.�^y6�9I��@�T�6
�����u�����*i�|w�N���k�c䉃*>�dg�WI��W.ԃ�uu&_<��a�v�W3���2%�	Tc>#��1�)�ɇ��fu_#�ݕ����������hQ��x���[;��E�;���t���\�Yq$J��.�hD�;�6��q��$؈�,_[��um!E���ťv�����^�'ΨŔ$��� �W~
�f���PF����k��A�O/�uoz�� ��T�~���f=�)m2q�]���uή��2��\�O,]j#]S^%yde��:����7���G0�̮�l���`����Ⱇ6��K�ff]u�q�v_)ڮ`�iQ���/��AG��cklfXg4G�ȯ��7�u)h�$�n�er�N��>Rҝ����������~�`ګ��j#�m�Sr]�Ѵ��^v�n7Y�Ƃ���EV���m΃�yv�ˡ��Iy_r�b���:�R�s.��٤�A�WC(�l{])�2��U�T6&5�JU�h]�'���Y^U�W�0��et,��UG3��Y����EV	F���=i���I������_=��of�=\X�!����U��붣����2²��b��m�r��׺�H*KЗ}fVpVAj�k
X��!�Rm*}>�����O��g��P��x@�]�M��N�g��βq����϶�G7i�L��*ޞ�&3����6���f��r��ʴܘ�b9sO_f�d�C"��Ӻ�S������m����=�鯯�&�/)kL_-/ad	B��ZNZ݇m���bk�z%��Z��v!�өyo�L��i�S��*�����̪�de��uJ�6H���.�%�v;�Mc�,"S�V+:��/�SjI�o\��%ooV�:�����їl�y\ʗ[��9�;�ޮ�%�_l���0�U�NX앦v�f� ��^���{�՜��V6�vri7�!k
"�#u>��k+d�0�g9`WdJ���������Yz�e\k�.��J����;Ox���ӬRU2:���7g4Ȑ�ʳ�m-4�\�v�ێ]�eG6�.��,nt̑X7�&����`�°I�O��>}�VFkE��7����w{sy�N��j��J��huDċӐ��!��a�m6��Ǧ����F�bu���x��+�xY��X�[�ܲ���J���zm]�Ϲ_9��p��c�rdB��*��rT��a�[ �n�(_D�	[�z��4�܈����`��k*z�jq����ja�vq��P�Y��*�t�W�o�^|W�O͛�k�W��V>��쏦�ۉ���R
~���4��VT$1=���W2#27���Gȃ|�a���{Ʃ�ZU���o��T8DV�Dł�S�]�b樥��*v�/�W���):"�'�Qs
Y�Q�2\��>���U�åUWo��4�G!!eF����<q;��2�	��#Q
�\���2�U!��]+F�8}���9q�tddr�d� �	��ՒZ,i1�I�!�4���rW���N�y�5Qv�O)��ff�.pe�S�j$U�k�����J,���}SIt��SO�x'魕���5_��x	 ���	��6&R�IL05�W�[&j[�V�C8�T�+� '�s�b ��<d�N�zi�w5�z\���;�xS�o�|�6� H!�i�LQ�dC�mۭ����~gvW��)�xOC~05��ʡ)�~K�r�j�^�_>�yj/�g��d�PN���&����t-��0�B��Pb�}���U��s�v�]{h8��EŜ�vl�}�-m������`Q1��꒬(��1�ݔ���Uq�3���;�$���u�8i����.;�m:���/Fn��l�ʄ���Em���u]m6;������;o��gJ���ǡ/�:��7��01Ch����Q��T�e3���3]�IS�x�!9���r����S���m<���Z�y�H� to���(!�H�c�B�$B_!G:�I���Y#u�&�Y2��%si�Z��f[&۵�uH[qۼ�������[��UX��k33��e��3Z��:�VI
GRXf�M+$aV�I��b�����r*iY#��AYJY�Q��m2s��� ���^�R��WZ�1˫��$���ZUu_إN�n����Ba�� ^�z���hT<�f�D��饋�V����tr��	�#+=���價ӳ�`X6�nO����+�"ұ8j�T'�y���j��3ԇam��Bp:62��̀R�:P�s�ߺ(b�%���}2��0�/D�Myt\�,X�Z��s�[�/fB���[
��IX�cS%�a.��K�$1S!\���٠�6�#��j=�����Y�B1]��@�B9>��b}4^͢�@* mQ���B���6f궵�Q��.I���[���`�L�
��7�@�]5��ʸ���0Fԩu5.NMx��t�˙A~ݨ��喾NV�	��7����Φ1��+��O$9�{���S�A33<m]�	��UK��z|&�\=�w3,��:=��T�1���Dj�Ml��JbK��4��Ϩ�hD��	��uOS���*U��X�)q	��P�b��͂��5�hRJ^�����W2��cS1�G\���g;*��6�stjM����U˾<������2�3��/s�p ���f�W5�0�f62a�N��_�(kz� �N��Ҝ�
���&�R� =��)�b|A=]�2���ة鵰
;�T��X��<�]�ڼ�Ϋ��n�U���w��Yoَ��gi��&9Tl:�M{�@eI�j��wy��4��:�p�IŎ�=}.wt6�B�	��\�YIΏQ���l�D�p*�;ϟ��fyö�U�c�}�w�8w�	��Ɏ�*��+��M�WT��'Z��������B+}����m=G��e�I��7E�j�nW_k�=�C�k:r$2���KY-������3�&�L%�21ɲܒ�2�{z�F_�C=W�!��$KS�=��	��n0U{�R�U�/�^�v&�3�>�L�ۂGħ�܌�O�H#NY2)7ߠ��t'�A[�u�ߛ=�`˨f��e��(�AKVKD7��ZrMr� �_O^����Դ6Ҝ����Uʕ/��;X~[ߑb
�;"���������5u��fE]7f�V"YRD��䣗�{�7��Ǌ6�%/M�RW�]�)��eXw�;Q��*��'F1��į1�.����'[v��^��6�D7�+��W��X=�6G�wA8p}.�S�>S�S��O0����rkf*z�`ģ(��j����䱀�<&�G]Mi��n�X3Od6"X��3_{Fi�ڂL���pS0O��W�s:�+<
�HA�:����=ʻ����B�Ac2��:\`�.�T�׺G9N�WU]V�z�H ����᷒m�9�īM��k�%�@�=�Yb���r��7Ǽ�#؁շ5�*�Fa�y�	�NEU�/��#D.�j������1�+O�|ht�SG/a�Q�������+�W_'��VR�ӧh+�jx�r�U�Z�~��U4Kc�WG�WS7�ގ8�5�Jc��UL��Ԛ奐,�m���s��dg��aZ����6�a-��m6�Ep�Y̈/�Eo���~��/H2��:�Ѽ�ȡ��ĕ��9 ,b���r��w��`���)�QS^6I�;;��v�y�'f�����0E��Ӷ/�$m�͇k;���QwKݙ[(�,��Vg���48c�,�շ���n���!jb�xi������vu��e2f=���雷��S����4����t��I�q��
l-�B��#��&8���6�Vf`G:�I�vF�wԣܩ��٫[sa��{/x�;�df$=��e]�z���h�����,�\0�G�FD�1������4�N���H��)�5�w���.4[��3*�v�is�aVE�S	�-�.�.z���WB�eTK��j��vTy����ֱ��V�T��d����x!Ș�����U������Q�rͥx��Pfh��u�w� ��㵳�] �	߰��i���5��L���z~����T�=w�	Nz����y��2��[Vj���͹�%t+����E�!>tj�Ĩ̀ȿc���È���`�q�*�U�]�1O����ږ> �?O�̮�S6wz���PX�׏?/K�3���7d���]EX?��%����Wub/���}X2�B_�IQ����w�e�r�U�L���z_Lpߙ���B�%ĂQBj�%���(
����=�&��I�\���j�a<R-�ힺz`�=��r���֛aAvbj*$������5�c��Nh&h;�=Q�]�-��n�D�$�(/A��u�6�M�!^�h���@�^��J�KdR�F�L>4z��-��3��U��EI����+}-�6�:Yq��2*2��B1h��>��ŐHU��<͞�ݹ�]+��ģ�@�օ���E>(a 5�c��M���w��wd���;I%�ܹ�3r��#�m��l�1� 7S��&�<àm1q�	f^t�.-+GfP��oC\�S�����1ɇ��b7��T�`�巔���n�&����C�?]P}��D���e�n�P���bFN�\a(q~gF3Y�x�P��A�^�X\�D�mz��t��W�Η��_\ؚO��VO��·�@��j�Y��U����u�b%�W�-�䓛�e|6�vab�75O[���:����� �M裆�ì�C�6�ݍ�\*�H��E�V��*���ݗ�=���"&/nvA1��{^��*�ʧ4��X�� N�Š��.j���/\�5W�<!��	�����5d]W#3]y�Q� ���Z�朒�8P.B�m�RxA�_4`��v[��g_O�-��A�(`��n&�2D���j�}�rP�R �)_e%A���HU!&<���A�[bvX��Y��j>"�/)����&C��׬K�9�w�ȩ4W����(b��)�5��[a�ʻR��Bt��sֲK�{��
,z�OLCgY��y�s%GUsae�1�%�bE���&&�*BFn�u5�3~s��ں�M��<]�[���)����>��,�C�ޣ���H�j���ON��c�Ď�v�J"��r�a�����S`J�!ѺM�Q�Ca��0FI�K<�Op��vi�!��[�
�ȡ��!A�����3i+�+*h��n���{T�jԒ�bΞ���R��/�TJ::�7!pu�+�0�6ښ���1��kl�0f���J5#c:C�.L�J�:�l�Ιg+���o�_Uf)�%����enGH	]��t��.������%e������\bZn��x�"�,�]6ηm�(���Ė���[��V���SK�/F�b����K�.)vL��h�8m�4��]6��J�-�+3M6�y�"P�y�yF�.�O�a��Ox����	��b�x�t�T��k[W��u�n�k���s�a��L���ߨ��<9�3哽]�19�Kh��Y��贺�����Xn���]�֡s�}�K��)�)�)��u������'���C��]=�׹J3�e	%����j	���!޿P���B�qv�.e ,"+̼�T"]Ӱ�G�_�¯(/�������6�+��b%��$͈�!*z=�E���fN��0��i4�J�PT��T�PMb�z���"Q'�5�;1�V��1U�.	�=��0�8"׮�om|�Ďkh���ew��,&�� �vS�ř�%�����pB���hGS�U�of�#%Gzջ�K��0����M��)_����{�'0�s�Z�t��`���s>c��+(xb���v�/��Cʔ�,CW�Ы����A��P��^�;��+G�JV����yR&����o/j��I�Y�%�r�衝.eR̃�^,}ׇ�G�	 s벹A;�Eޣ���T��,��zc=�������	̽�C�|o,v�ѻY��,{[�������ɩ��8��u�&��1�Z�b�(�~�|$|`o�:���m�V�yy��,5��oQ}�[�&���w������?�	\Z�sY�T���Ѵ��x��x�F��D6b��2n�Mor���^Vp5��G��7N����x��e�e�ӂX����w�M�8pl�e����j�=�9t3�cvP�آ8��L��W6n�V�B�7��D�;:�[\I��nVG�OEs�^c�J&���za#%s�=��Ȩ"���Vp��3�7�3	�>{�UR&e��;����f�|���FG�Fh8�j�e3 08KѾP|�̉���ԥ��yR�c��A/X���W��$�a�E�<W+}a��,mjP�C���w�ߪ�'���^G��G��:e���R{�륂7	[w���1�y�J��������Ww�`~�VE�BU־��=�C�j-B�tǃųEJ�Y^��:̓����(8]U���k;��}ͅ���S���f���c�YP�"i$�+�+=�~�0�t�QC���v̈�t�q�ܽ�Ң�ǽ^��*��whBL�D�����!�(��V��zP��rg�����PR�
`L���/5� ]�Y݂{����y�]}��B�}F~1���*Y1}���t0z��9\`I"�Be��/�%Ǐ�f ����ưG����B��ktTD�9 ܅r-���MOruH��yt�b���/�-��5����V�ˤ	��{���Ԉ�B���������J�Z
*1t'��}}{|���� �^i	�H��a6�����R�R*�\#ٽc$�%�]X�� ���R�a2KF4�i"P`U�{v*	�ٚ$l[�j�r���30��cD\vfT�>U�qG`�t���]v�}]F�z< �]�`v�Ru�����3T���FӐ.�K�(v�1�w�u��7�HlK��x�U7\���v���x��B�;f�_83l����"w>�v�:L��O�Z�q��r#l9�'� ���F�*��W`�:L��,��d��s���N�
�L�gaî�J71����B�B�U�0�Q�}k��]oONm_g�����X";�P�:BT���^T:'/q>����d!7b�ނ�P���[T����@V�a	�Ջ�,��ӈ�w;�4P�>E`�ą�q��=��5�x�{3��;���h�r�+�t���R|
��nH�����Omi�S���z����/5Mō��:6���G�QDW�"�\I�B
=UX3���Q���{l��0g�h���t����I�R�_ܘ�����z�z���&�'z���d�um�~�0��A�ZS�6�UL��3�+�a�Tt\`J����fw~��5D�{�=<��D��>He_�Bs6��Rg��N� ��&�ނ��i��~w���I��y��9��s���b��KN�i�*�
!���$O�������U[r��,���V���(�_]Z^����3�ϵg���Tј�k��i�.�;��x8-SP���;�N�Ϲ#~�ڿq�ہd�4vn�Z��(v�	�»5f����g=l���'�>^��>����3��/� H�e�2}B�r��]���[
re�r:]#3v4���Ͼ��y!DlP5�a#mxD=�G^`��*��%co�$�U��y�wf�)&�ќm��q��DS���CKJ�k����6��N�0S�O��zs�_v_����s�k���h���;��QO����~���7%t�⏻���!\9��t}WG-��*w1;U��!#�u{o���|�y9��8c�!���ג=�D͟8����qM���tA�5b�y��d��N(�{��{]m����?���Y�������,�	bX�ph���l^����a�:������֯�@Hy; ���:�KT�k�$��-u�8���v��ڛ(xD��E�1�8Y�ڶ�&2�ҝ���;Ui���$�`���ֶ�:�jQ��(d8wځ��񥝐:�B�8���џtf�� RN�7���	�D FY�s#������yT�$�.Q�[�:b8f�f����ĉ&�|��2�D�Xee$Uz��p�����=�l4zX��NDH���u^l*��s%cqS�Ư'og�6��9������}�ݳ�L-������\�dtz{��wW9Y^��N�1�7%�w�:o�b�DZl"ɮ0~c���s��˛/�湠Q"���*ڪ���;�N�ǡ�1c�"**�'`�Xz�O�D����^0�=30��:q�-���V1��Ih��W�ܶZ��e���������:���jذpan�t+z8ϋQ�}킔�C�{Ü�4ɡk�ބ�Z����>ۦ+.7^���)������%���έݻc瀇���WB橴��Z%4;Er�f<�Vf_w�\YH��cL��u��-�'�Iۖ�v&MGf]5�Ӣ�.XĨN���u	]O'f]�y��<˘�����HAP��n���t���$���l]$�n���6��;B��L:S�ad�ʗ237V�n��՝<'�1��bI����.���m3�.����6��7�W�ВD���$�_Y���mz��k�w�?_���:��A�1<�}T��8F���M��h�/z��@?,�C{_2Vߪ6}]$��h�F=�b�l�ZU5}b�|�,gH�&^4SM@�A��R&xs�.*���2�
���e�s�����'�	��}3��$����;[tG�ӂ�v�\z��t�^tl�lb�]�������=la@���<��^`�������)�^CT\�Z�� 0���!}#�Pq���&�_���WJ�gO�W	�`w�]���馔!��P�	����d�1�����S\�+�U�����ݹ�x�<:O=�B�5��5�9��a[�S�N&.�nF��b*27'�/X���_�����g�	=@ҫ��| {R�W�6�{n!3���&ێr�,�U�����A[�U��)XI>9Bal���#:H�c��뷵*JI�0HG�ʽ���2�Cs�7`�k̑�O M@�~>��1Y�HL�(5�b\n��2v���j2*���\H4��c�)��9��� x>s]q�S��g]T�x0�Ʌ�c��o���eH�|���o�����]{�8�
d�-,!��Ķ�_��0���u��$/�?�����Cu�J`���:r!�x����!@��yI�|����8 �Nn�Ep8D��j��ӂ��;4�
��|ȋUB���N)�S6�R��dd���H��;�������ڦm�,���aI^m��j��e�rK��DS���u%�e�8�c5�
��ݹ����3Ap!��-��acv8�\�ZO�N�Z�teZ5�j�p����^K����s��7��Bj���n��wZ�N�ngkU���`w�W���ot6M3U:��b��(]�ճ�<ڑ��P���]�Р���P�]��ڽSpR�u�@!]�Z���VF"�l��z���>��RJi�}u�78����U����.t�+��j7�K)d��ܨ���s���B�5��ӢV�/���9���m���(	]͡�c۞+H�C��r�d�fr�))H(�wq��Y��r�;�K\�H���j�u&��sx<�w�ÇWu��J���/;�����FN�L&ׂ�С2�Ȗ�zrVX�b��u�B�f�M����K6����,W*bd�w��	O%�<��}��D-Kh 8r&����V�}�åU�n�p�ޣf!糪�"w6��r�U�&�u��OF(�s�m���zE�[[�/j̥��V��+�Xhn��wxh��HFe����gQأ
�.�K�֔��p�	�`�'y�]�z&�e����.�8�38W1vN��UK9�:�C\���uÞ:Z�
�ƛJ���Ofb����'����gW:�#�q�FE|�[I���+�:0oH�1��l I(;<X��kU����s�N��G�ȔCͤ,���-b��ꝗt���^�w�g���*[�[<L��{�w�(j��'��Z�-�ӝ|bW6ծ������FG$�Im��N$��Q��6��sPWn�9�� ��/S�4�}�K����^�q��p;X���A���{|��x��Z賹#1��kr�^�}/wr^�6r�����O/��s�83�	����*e
7�ծ�rݵ@��U+&oT�`�|�ص^io�}T�2r��
T�mI�{�u�!�+m��я%���U�u�=�M��q��A��v�����Yީ:c�ª�rW�t��a�xS:��u�����8�
��C�騙mHE���mP�j_��La�6e�`�\k�V~�e�v�v	6m��F@�RR�ۮĝ�ZF�m��Đ��|�U�B2Ҭ��d�ԲF�N!�Yn�^n���6YKO����vY��L�J:���k�����\�D#�|�����++Q�����XT�WHT�ݳf��̶F���%�Ǭ�	�b��4�.�I��e��6<dT�A��"�&�ln���16�t�V�\1�F�-���$2�HMe-�(��ZBKn�F]�er����Ul��i�Ynq#�GDΩLK���FY���n�{R�&���ǵfu�����[U�fo�>y3n���݅����0��Fc�;E,�Q���RV�^�i1#p�H�ܕ��Gd�#J;M"4�kB�=zI]e���I���ˑ-��l�0٤�K���:.�(��zeC8�ėTA��5�!���ЖR$���Tv�u��Z6���f�]Y&SX��.�[�ܰ�q,�Mn�h�&�id�biD\��1�Z֣u��YոMf����̶�X2v��[l���3K�     ��g[:�۞����;�����G%�b�omޥN���=՘X�X:<"t�5��.�h�p��qsa��W�W�M;��3y�,t�4�|��W����j]}��| �<;,{Չٞͧ��#$5]��Ա��o��!������zbp�r�%f���C娞؅X4� D��D�N!z�ˍw��W�%W fY8	��۪ԯWHQ�\�&+L�IrgHk���U����$���UƳ����Cs��2�"F÷�����7�UG�H�s��?W����M��v!St��rv'��q�d�J��Q!�L��S�8jw�k<���׸��.-�%�<��B�o��7æB����U�CgF�o]_�|�#%�O���J�1.�mͿw�u����}TAw�}� C-�֭�F�b�����֦Lj��������t ����i�牍2���PkClJ�h�7���q���p���e�iq�;�DjR�O�b$܆�ћU.q��?Ut���Gȟ+��TN�K,�	���σ�Lc�!��?v�*���o��H��s� ���] �B��x�T�u�o��aW�D��ۜ���p��B)���vx�!�ۄ��F �΢nh|g!�-�?�l_�d#��>A@��N�����l�!�.�HP�>2��k�cf�ƻ��w�)O�U$;0�Ͻ��z�\P@�赣��<��}��=�޿�ߢ��Kp���>����H�Pn(�Ba�B0ZI����R�����ިw�إ�HןV�Uq�s Î\$�~J��D����Ei{�401O[d�ʮ��6�nh9��Fj}�	�cp;R�+�̜����NYS�c�̂�ZPK�nV��ɬ��K0s��UR����{7�h}������2�N}���LՌ�f�����g:BF�HakB��%�H{�����͔���=c�H��Z�����'n��EnD~f$���i`[x�U��qi@�
xU>! n���(�b��﫿pK�
�k[��|(.i	���&Ƅ�g`�'4��t��s��s׵ס׾�B&�Ln����m�J�y�nl%�u�UixS���[�p��be	�>���J��swq"�oKڐUX�7���٘g��s�#����m��6QFuڋ���E%+�i{}�V�\VjB�ѽ1eD8����`X�N5�n�9��jרX��ڿ��*���b��hM���V���U���>�
�����L]����u%�א�pa�9}+Zj�T���8�� Z��ͳ"5�����v�*LoU���;����IR)�V�""�n���-zq�KޠTX��]m�-%��՚��K�8��7P5�{E����I���W	A,��(8
����'��)�A�{�Z�\�2pޮ�4x�x����g붏g�MT� ���=9[�S�������n}�NL��k#YW=R�ۨjd��;�T,f��x׎�Vm���WD^<V
�Ā�����O�b\d`����N���.�(�\%0��C^7ӌʫ�I[v�/E`#�В�����1w��b��"��oZ>�^��O��X�Y��U�����b�RYH�M�c�|�R��Uu�#O�6T�d���^�"}�T�7��1~u�1���KKմ@�+��*���ܑğo�Yۜ��nƮK���U�c�ȅn�(��Grv�m�F�[����g`B�2|�(�K�i���u���9=��Nj�GN],C`@fg�.�=O�mĹ�S3~�0�`���^!ލ�;Z��5/�7ry ������ʥ�b#��Z��GKF�'.�fl5�e�ky��Hs�s�ȓӖ+�e�֭��؅]�(~q� �-b�>h�3��2F5zO�qSq�,��T֟?OSTH���rk=�z�ů��+�����\�����F�i�>r���2�Iw\f0Y�ڦy��^�䫬���5���]T$g�v��fQlX*+ #2{�n��3+Ւfo����[p<A�|'�ɋ�%&���7f<��2�sռ�G����33&�e_>u;�	��dD�g	���{��}��
�u���;������s�s��$`���aP�(`<�:��U�ц�r�*���ﯢ�z#E���S��B�#=��Z>f!�y{ۜ�R�F����A�UQ�-o�h>��LyG�)M7�N,�k�JS݆o�o���f�ŞFA Ͷs��Ⱦ��@w�.�}�)��}N$J����;WA�wC�֌)�΍ k���yi_Z��i������5�n��g�=})��y;�U�ͫ"M��!L�ߢe��Ч�0g����&Ѩ'�p�Ʃ\�<O��3]��u�Sԋ����?|%/G�����&5���l�6�Rx���+r�k���j��Au���]HF���Z�,�b�Y����Ah�ë��Y�쨬��ۢ�C*7΅������V�(�!� i��b˜L�4�&s3��պi��[&�+.U�O��Y��"D��R�b9��(�]Wz�ƍ��Q��0��ij��$�8d��[,�e�6��ͦ�r!ȋ)�ڒI!�T%�f�ݫU�?�!���ț��|��^�&��K�ӻ���R�}��^�i��=�u�{��
I�C)o��Ɗ(�r5���R��]q�|PZͽ����,h~�a�"�W[�����
�Sΐʍِ��x����ؼ��/��=ݹ�PZȞ�".�mW����;w}�$N�dg�IH�t#�l�����V.�p�H͸g��_�_��w۽�Yd䘍�L	�D
N`��p�>��!!��j9+`3�?�����(���GV��<�;��M�f��C��KD��	�H{�Q�����L/�ȑ��l�hw1gכFn�U��Q'�C��ԍ���7C����SXj�p�pf���Ä����#�nc��C�k��������y���/K�\w٢VZKv��L[�s��/e{�m��Xq��[<=g,��8�W�]��feM �޻�K6��5���7Ĥ�-��/��#�����m.�;P=�an&�>�.~Ն<y��:2���Ge)Ug���hÞ9ڮ������wI:U�١�v���F�������AK'�].�=�S�a���n�m�K`�x2:(g=��;y��u���h�vC��)����>n^��_t��f��µ1U럜��_]�(��2�baG�h���C}qBq�y2��כE�B�'��Z�UF{�]�	Wo Y�sx�zp��S���io�-
���kp8_r2�p0K��	�m�)m�	���׹j�}j����Iop齩���w����=��~�M���6z�E~~�;�����9��kBۡ�)�u���q黔ceA��D�	��-�<�S&6)��Ip`��N�����t�ozsm�4�vf����k���/�1)�w���*S���@n�������aG��j}쉓�;نHp��ZIϵ9�K:��)���v2�[�}|{s˶䞋�۵w�W�r=��c���\��0�'P����E�乣i_�����x�dWB�S1N�}5R��@i_���e�J3-��~z���X�S�Co�����O�&a��D�^��
�w��,6 ���������ݾZ�ׁ���iHq���Vڍ���h'ψ�=�CN��q_ہZO���;��),��,g�Jm=W�����8�V*Գ0��Kzr�\٨}�V}�(�=Rͻ��"��A�w��e�-Oԣs�p���DX
�W�;mu�l�������p�l��y����C�]k����A�#-������ד���������W�>�l�z��>�8�tľ��v1��Xd-��Ԓ�v�)T��b�P1nUmH��tP�>YZž���/�{��[�Ą$�m�~��h4\�(L�0R�r��<:��ay��0��T@�[x���3��e\45�ʵ�����[D��'Љ��.܋����������5�'�]�U>��n��m�u����cbf�'mY!�>#���z�En`�b
^��a�/��C�/p�bk��X,c�w^"���l\�]�p���+�@��ݙ;7�\zb��T�ޡܦ]�aؤG`�
�e�ob�"��uy���������5֨�5��y�{4�^��wH]Sݾ�)�1����U&�������t�a��k�UL�SQ�GB��	ѡ͕��wVf��+{��kA�m`Ğs�M_ɥ1~���	��
��� ��W3wz	V�1� X��|�
�x���������s� ������:��G�0ةZ�7�fH����Ӷ;}��M�7[ܭ�UC�'�J��3�����GQ�X�ԇTÖ��t�Uǔ�%[��ݿf�m}�5�I*淡O�Ǯ���;{zX'r��s����{ZY1�C�=���?���<]o��B+'���4��p
O��?������n����#�ݛ ��_��}�j��~/����i]c�iI�
��8p1P}��ɗ�~���Y�O˺��.�Z�ޟ�iqǩ��Url���º�$��nn�t]�rM��6�����r�	���"=/3r/�=*o�UK�S�,�6�9�0f��#E ث�]{6C6b���;�V�G���C,ٞs\�����^)��WS�E]�Z��W�I��kfF�gCB���dಂ��t���A�����^3G� W�[��ֲ��'P�0),���אo�#����?A��b��[��L�މ͔�yݨ/�-�-����Է9q����ێvoU=��Vu��)���"X'�Uvd��=>8�0]^Q�&&%��l��Z�u��N�����,SN��Y8�w�y�w�:�����JD��;����CT�ʽ�Ea	p����]nF�Ȫ_n�'�eWZ�t���0�L^�I�߳kV��O�e.Oۯ�E�>����r��.���!���I/!�����@�B�;�
a�8���w<�:t�jJ-y[.B_Q��I+4��QXOR�|=��l�v�%��
��9Z��ݙ]��$ׄP}���v����2����~^��#z��pa/S�0�ኬ����zr`=�I}z�X�o������J��;(_�di&q���:��K(l۪�l`��T/#`�=�rwZ<1S��$Eਔ�>]�Mye�y��țT����&;��t��o���k{��)����K���ձ5�)c܂qnu3^}�Ǜ�ȥZ#�2�8ttd�̃�č���P}��'Y���1���AA�b
f2yN�eP�b_��R�+g~�e�O���5{�ء��ZQ��A�}5��(�99N�Uj}n�����r*����x3�f#BQ�9S�����7s������럇�1���6��z����wH]����Vz�����Hv\�d
�峠�i��������q�{�U�ǔ�xj ��D�[3m^�����q���L�����;�����O���R�퐖���z��N�\�\�t{R}h���^�cr�}}���cM�b�u�3z��DN
����p�N;�2(���Yqa�i%�u��.��z�;@0ۧ7�sD¯+�g���� CqY�H�f�%u��v���m��`�I��X�9���c�ԆF$H�ٶΊHXH]t�a!����]v.靤��Z�ΐ���[f�k�Z�	^�n6�X[�$�A�H����uu�U�PV��^�F�)��_Qa�y��̢|���(����s���+wp��=�Ю��:7� ��,S�����-��)^5Ć�$>tt�5��>���:��X3xׯ9�&.����5��1�뮍�$��H��F'�S��� ���^�'��E��+�S	L�yPٹ��H�D��B7� 	X�Ӊq���a!�H�H-%>Y�{���3*;��*7�1;bw�,U�ܭ�1��t'�▧=ޙ�G��kFıXb�	N+�Ao����E���w�=�Շ/���<�R�[3<HJ�g��	�G�Q�ze�@�!_�Z>�{���Ԟ�x4^�I=�<EY�Ez]/;�'yt�+D����ؑ����"EF�XH�ϒ ��i���ч�2|�¯�ܴ암i�Ct�-;+k6&��Y�:�&�*��n8N���LD*��<��٣*	��6�sAzf�D�j�)���<3�Ϲ��>�,�KY�d�L�<w$Y]����ו!I�ж�ѦhJ O�W��s}v��F3Z�F��Uӹ���+�n�ʥ֟�H����s� d���`g�l̔؏j���mˏ;�����[��<�}Il˒�8�,�:9"n5>Ro�)Wy���f=B��W8�b�cغ�`�P�V�L��7��R�[S''�1�sOL��6�oh�;{��jٓW9]��s6�Y�Hk���5�w�ӻ#H�UЉ�k$�8�ǬL�Ӂ*GG5T�����S��W��ofh��=�;Ҝl�9�Ǡ��4�[?<���=N�^e/�#��A�6�;94(�I%�󇉽%&j2$s�! �HP�Yp�I�PW���~��h� ��_\}�%���R�����zA�yJ�:ZI���=�_�W�Cr�)��v�(�ʯ < ,n4Ѳ�Tb�g�u�1im�up��g��g0�<9�@�P!��|�D9�VC���VK�6�*�����!?Y*7���Vy:����F�E���PN����p"kv�=ڗEiy����v��,$5>���F������b['Wo�3S�1!�q ��T�=^���f�9��O6��P�L�_��aVo�~x������1t��uӿOU��{�trx5��}/��`�}̳9&
�)����Օi�r�z����~�mC���T�NP�	�dQ���W���8�}}IWl�	$���)c8�D����3+|�m@<�m�?EYHL�#��$qkD���(�T�;;�c%�ۜ)C����Pp0��B!QF ���e�sb�˺ut����[��C�p �[^sЃ�ضZ������$�/���d��y���{���3��j��e �^MO*6ˡw��N/�>�ӕ�Vˮ Ҷ��]�C��Շl��h���ݛ%=qEN�5�s��U;z��C���ZL��U}�V#UVvQ��>�i�N�u�%ޮ'�z��k� �K"�@CCk�'�,�c�Xkv���~�o>���ب��>F��Twӷ8�u�Ͼ/}+е��Kg0`	�4Y��cl�(���������Z���7��7��\�ϥ�TT7kW\����jʲ�&/9����Z
{E���/V����֯��+b��7������Py���_�����;|���\T�Vz��X4��v��r����<5���c0�\� �,��F�x�G����#�d������"��rjE�	Y|���M_���ڒV����(T4���CD�z�aɇ�*=϶�H�,�T�(wv����/޳� Rw�۲k���J�ӯ�θ�.�ZW��~R;�!��Ex0�'M��B6؀�l���$[�3ނ��9�ҁ<�앑j��g�V�_:�/8>�l/���į�^p%!�D����i߉�;�N��-h�:�e�=˭T�D��"ǣ����i��M��v%*�!m()�9~|�Yo�k����3UW8���QQ��8HC�mR� ���V&��&(W�_.SH�UFvv'��`��Ƭ�5�Dm�-Y�qX
f���!K��M3�&�͹ou���/�t⩅��y���+e��S��oy�.U��m����o��X��˫� �܉�-��\)�bҕ���qT��ԕj�v�0&X9t�l���Yp���jP���i���V�� �gu)�JMͼ��FȊ�Υ1�nQh�q�*���7U���JBt#z��v"��5[��Ngr���G��n���)-}G@ѹZ��|G�3p��'�L�t�.�z2	R.��? �� ���i�抳G4fj.7F��I�`���s������lƨ�zo��C&�Ϟ#	��]�z�k��x=�b��A�I�[-V�e��s4�QעV�a+�z{M]+�8r�Fx�-�ap���$�X���<�I�$�A�fЪ6���{q��>��c:��5�orΥ&E�]\}�"w9ݵ�c�#c�'BМ��cZ��Df��I?uӵ����ʄ��T��]֒0Uͽ��q�k��m�[��S=�B�wink���XZv�Amp��5oP���ޙ�(G.Ӽ�����v�[ a��q^�o�9��m�S�oT�ZP���#`��$0Hً:V�|�wt�g�kE_M0��7�V ��J`!���e��j��������p]iP�����ԗ�mf����l�:�I�}�8��K����#K�m*��x�:Z���\�h;3�}f�\�cj��G+Pg0aGI@]Hh��ŃK��f���k�xn�5�bà^lT9��b����Mg���G�^~�eW��pj��<qCs��Zz�֢�l2��S��:1u9�!�ӫ�][�γY�G%+x�������q�)�+�C"�]�0�D��wt��]�HM�_ ��z�V�˭:�g�Ow㕝���^���z�[�vB"���hв]�0���=Z�m��z�T@�m���5�>�K:��1�	��d
��Go^��,g[��*���P@x�U�v+U-�"Y՞��`�q������ �G,_MA��+������c.\|���Mԥ���K�m:�K�AcJ�wQ��Ӈ��`���oi3��]��}�X��_�u��c#*���{;Nl�r�aی�Wk㜝	��l���X��7��d4'֞_D���6�քI�:;��Uꝑ�"��i�#�ۥ+Оu5�4^��6I-��ԥ6G�ͧD�\��ϏU�z���O���{�!uj���U�[A�7K�yق��2O�d뼛�B��Ĳ�g4a����tp�v����[-�5�r�=hz��DOWB�є�T,&���4s�0��"H��|e����r��YZhD꒕V`��J��,��	a���t��_q%�f��1��}[��Q��a�1&M�B$C ��\�0�M�*5;^e�����T}�v\�b^C4G^=�R\]���f���z����z�p��}A�q���U�4Oh����n�+RyX�g9�w3R�%�E���k�/9y|�W�!��uEYWY�ʑ�U��^�r��{f�3���'Տڻ����{��,@�`�����M�/�1�ڂ�J;��ǽ"�ب��F\��e��U#7�=��E���/w����E"�=��f�Ξ����wҮ�,b��0�F��(c�>1WBL(�8�#Bn6ŌJGrȸ�[V2��ɍ$�9����_��G,>����ḽ7�����&�����>:���vQ����<��rnm��Uy��j�TdHP��J9:"�Z�\�5����۫�f3�vvH���ƔԥԷ�=�d4[5���b��mp�B�W0J�M�2a�	d-�����ҋ�F�훖�
p�\�I �[Wo�H�::���g��QgX���~�p� ����^ʍdk�#�����Ts^������?��?{'Ϫ�JW�^��� �}9Џ_~�]�z����Wp��m���e�����W6Vڜ���0�
Fs1ᛉ�F8GGF�vT�!���x<w�K:���\-�Є6!��,��
8l8�!��E�#�������ti��R�S�QĴn�:��yalmX�{��9��$��jgs�CT';�M�1^��D!����L���!܊kb���]\+@��G:��[�Z3��R��n	Χ���y�:�D���TQU>'J�GyQ'V|�f��z�O�v�+o�~��im|#��4�ū�ScO�D�����'ЧC�q��~�}7�pnw<I#}�Efp<�EF�>����z6�u�r�R�* ��ԴɌFM]�I���׫�~��#�I(-�%�*�x�C����ɾ3+�싚Ňs��^�Z<ظ.k_u�w^[|�;�\7�c��é_�H�}>�UWv��/�b4,�����B��4��9�h�W���ZR�u!F�ÿT�֋�YEh�Y$�	��N��
��\t�Zm�v���Q�4�մ	�!#���9/&��S9���t��'G�lb��B����ȃT�x�x�1��>Q>������:�t���X�B��L/�i�S�V��(�C>�S7{��E��l�ݚ�0o�=g��7/��η�7�$Ưff0�Ƌ�P���b�����$ѫk�钪��ǔ����'��1��S��U�C=w�.Qי�rj=w�̸Iʒ�<����E̩y�j:z��EH��y�^�{��,TϩDw��w�T��#e�y3iv�te.�4?-�v���K^�b�W�x(2"<��3���m��G�i�uwS-��=�Kۚ�hɅY؄� �}:��f������S�C�o�xH��{�E���l�4��Q��A���f�Ó^S�~z�<]�q�|f�z����#�y{
��
��	�[�S���R��}˫��:pzM9͞�C*�#Q�?ng*'���HU|�����ɷjUv��O�z/�E���
����jJ��fA���o��+�xq���G�|��{�Ji߳�+�1�.ݳ�r��^7� c��M��2�����,f�4$�i���S��a����Y�Kv��ƴ"� ��V���Y#G�_��7w��ƭ����<ėq9`u��.v��rF�^�|xRc�W���[�V	�v����=�D(6��lb�y��*��Nb���V��Trj�rDL�H�m}t��+y�b�x 
���܆QYN��k*���'�Q���S���Ʃ]c���U�ʕ"��zԝ��l}7�«)GVVf��1��A���=Bs��5�?uNز�(У�F�dt������m��!�W>:O�:R��{E���W�wK0W�ӗ�eȪ�2E���{"ō����.��v#�el�ˤ�E����]D I��H]���YW�{=F���1z�-p��hEs�,�d�~��
,�{[�:6�1x�pǞuZ�xs����F��c^�?f���)�F��2�i��D�����ܐ�f��A��Z=�x�`��������M�a��4�ϓ1�"iL{_y�������
*mi�S�}و`�U�����Q���o�TueೀN���h
��$��5W� ��A�պ���fG���!���b�DUʷ�+���W����[��!&�	i�b�lz�z`���UU���Lm2�m�bLm�p����Q]���WG�pq�
W�0�O�Dkm<�Y�)c�gtG�c*�P����6�Kޅ|�� C�ٳ����[\�����ZQ�:'v�y[[K]����yTׁwaOzEت^�q��/���w���_�vު�z��Gcզ�Ik�[\��v�R���F#0��`91�:�0���8����<d�>�oEn^)Rm���z���C���N���$�9���>�O.�8 ʒjH��W�o�H��5ʯU�U�M'����B�߲��hl���^�Є�̎�ݬ��!�?>�m'����~ɸ��Q����J�m�h�r	����X
a<^�Y1���U⇈�+�g�Ͼ��wM@QM� �Bl2T(�L�4*�n�F��A^�	�F��/��w+�v��W�<���%��K���e}�|�or={���c�ͅ����!��˕d���dmgT�.=Oc��9+��)|q���W"D����٩(ڳ�d��+�8���'��O�u�Q�lu����-��1}/�%Jc����نpv�J�1�'�kt\'t=�n�T8I=���ݓ,Dk�e���\f.ԩ&����!_�/�A63�y���ȩ��0�q��n��zddfeFFy���y�Mo;�-e7)X�w+�L�ݫ�}Mn���\J��G{M��B��I'���D��ZE].�[3�8e�ݢ�����f�I��m*4��:���R�j��[�"B�i����D�=<��>-3&�\�gB�_$r�h�G12�]bkk�؅lU4���Ļ2Z�MY���rIvd��l�d�G�Y.��֬v4��Y�D�T&9�I3B,�u��<��+�o*��{�Y!�Oy)G6���<��;YT2%��"�<9*Jn��n���+D��o���7]������i)Iڜɍ���
۴^s�z�~=f wYv���#\����{z\!w=�	?/��{�P����鞜�.��>C,K���J��~Ӱb�BF'	jC�5��"	�[��=ޠxy�F�n0v�<ӫ�?/:��pL��ޭ��%˩�.�N�-+��I�V���{tI(T�Yy
�t�bI�E30Ѓ�h��כ���f�p��$jY�WrR�c yp��R�i7pA�/n'7�j.�6-q�7���Dv�����}Pb�"�"��������ܛ'�x��QQ�j���ǯ"𠵾���)�ziw5��{����01��^�1���S02v��k@�ͳ�*b�鉞���5��y��l�����F�l��Y��v{�urjP��'h�髿�l���>ނ�`�~�Gr���������z��{>"	O�,�t<�u��t7���ÞV�ם5A�>��xl�ļ�Ԋ��v�&�+�Vͥ��M���k�?5ظop�aY��:��%��r퓊�����d�z�\�Qd̠�*��a`�Y��s�vL]���/.�(�=9��.�������تw&@Z��:�״��D�͂�D��a��
HS�a]�/:��\��	��R���_�Aʊ6C�(a�_͒ 	p�]:��:��&�X���a5���a��/V(���=;>�6
�Q����p
���Iφw����ʸ�Q�f�]���qJ�����n!z�,NuM�+`��N����W�`�T_���s?6�EMG2ЇLn|c��׵�����P�uǃ�FE��^��e������v�տ�fy�!�`�߳a�(�k����	P�F���D�*�cܶ�����5B�!�i��6�{V`aT4�:���͢m6�^��z�w��}�����۟o�}���߲ni�ñ�1|�"aխ�S}{Q��ɤn�_�f-(�ף)U�o��=� �WjFv�"�sq�j��#9�0��&���c�Y<�i�[}�**N��P�{-��m7n�7a��� 	z$񬎹��;#w�/��R�.�ͦ����m�hK�\rv�ڗH�|}f�x������>HB]�p�>�?Pzr��;�vDYa���y����f	�ֶn���z�\V��uޜ��\P�X�՗J�0͇�6�U�D��L�ۃL��XÚr�uq���c'1ZP�ȣj��QLrLT�������z�TE�V&e`B�1|�W��K����
3 R�ۥ���.�^���s�=�n^�8��W�WUSh�a#����%PT��uBE�rU;3S���u.7{���<��-h,�w�"Þq��q/MR��f�������_�O��1�}f�|>L�WwLnAԼ롹p��0W�k�^�b_ �fsC7�^�}�^C���_��v�+�A��f���{_�$V>�>_ۅ�}sdd(Y�J�p���8�|�|�=��&u����r�:Y'�e�TF��`�?e/8�z]q^���C�^%ܳ���z��,F?p=o9�Ȣ��ռ=w����-�Xu�G<g`������n^�s4�R�P*�BYA�M$
M�  ��
l*�`Ɏ�f&x�ՠ�ޤ$��c]HH�ꄺ������,�<'sk*�/6)����LhР�Hʺ��we��r5�`җ�^6�\�X��L�e���;��g�wb��v���J8�4F	�V��_V��w!h[$%V��*��^<3��}Q�9%���B޸�ot+��Cl�9DUK�I�&�q&K��(M��&ޚ�Se.�����YG\�)������}t5�v���˺��}zmu���%p�@�����dc+/DQ�OpB���h�V � Wnnѥ?�Yʇ��v���V��[�?)�#�3���]�p�.��M?[Ϫ�T�P�tŰѝIɒ���bS���yt|����(����nc�i���8��>��ŷ�z�S��%���g����a��'s���U�E6�n�����58#uSh�n1Q���s�TQn�����<E��k��g�U�/a��:�<m�n�J$��%B�����dV�a4G������N���r`��X��K�{3�\}��[�i&�lb$8�0�A�����`�G�ǝ�\q&�e���uN7ָU؇O���m?�~���K�+�Cz��s�?v�݆�d�����"�f���虫���C��D=JA#��Y׸�DY�áK*_x_�����{Дz�|t�l�{جe[��x����Gu5���'��-I�O�z�p�)j���9�'�}�إe*���x�Q��XϒH�;w*J��T�����q�[��O��2pq�b���ޚ�󚛻�o��R*�BOtR��t��]#a!iL�v9�Gk��Z��ǵ���B{Eսח�w
]��������t�wN�o6��t��jU�a��OU9q��<�D�Yٽz9S�̫��UB�AYn"�itCgy棛	�r��|�d��]1
�E���S2I��4���B-���c��ͦ�ͨ�-\�R�8c3.k%��<��L-�$���Hݵ���Y7a�u��W2Ԓ�BRI$�k;Jڥ�xr��Q�沇�7<Lc�~��>6�o"Ng����O����V�lPH�C�����o���=p�7.Zz��F��=z��`��l
�z�����66*��wn�Ӿ~N��{J��bB��&(��dq�~U��3�R/�;Ͷ;#P���*��A�"�D�0"\ Cǂ?Eߵ���m��g��y�d��i����֍M�����⚔dVȷY�&OfgG�&%&���g剳Pb����W�6�M���秈���&&���J��M��_oq�*w&��xh����8����+P��3�F� ���DZ�	�_Q���st�f<��+%mc<�ݼ�3��mFK��9r1��!l�Qgx,J����21���[C�N���G_ [�YaߜA��w%\H��� �<e׎�j��;�����t\�L����C)����n�V�G���M�=ͦEC��>��w����7���1���g�e��Ȫ�^���ٹ2�͊{��6O�wP���{�a��[K��fP��È����J	m��������.���mu�Mͼ[w&�v1@��ӫiw�Z�A�*B�K�M�G��R��L�k2湻G� ��r��ѣ���3�0�_dp���= &��7��Ν{�5�i9#�������(�멇`�l�g{���s9Q�Mf=���CW�x�h�E\=�;�Z���6~}�N����z�k�*�<g`�Y��'����S��>@��@S!D��}�6v�(�� O-�8
&���4���r}`�fˈ#\����g��f[����L�W��
�Шi���%6u�HZ��"�oS�c���i��#=�Z�#ZMٗ�_}��� �ӽU6�&�X�C_V���h��k@s����.�rտ|	�/m�D 2Q��EE:m���@���q�}�@>�ck:l� ƾ�.KGm�pU�1���u�\d�M9��kM�,��ڳ��N�Ĉӧ#OÌrR�x��SviQ������� �>�{~Ä��_�q�#�����hΨ�T>�3]����9�I��.�+��j��Zi5����~�e�ӐPL������`�h�aÄa�J� &R0��,�{Ւ���4@�j'���]J#�p�')������}e�͋��$�ZO��㧟�g�'����j@�ޠ�j<�H�x���"$����#B�!r���+����8�l���{+�I[A,��5�K��q��P�۝|f��5H�Y��+�1�r+dEl�z&� ��IS6#۬,��Ӵgp�ܮ�B���w@�C�G.�t�j]��s51�q�)�k;��Ԙ#��;9�p�U����RYM��ڸ�3Ζ*A3��9�G��1N��I�_+_V�5�}��e}g��ɓ'(�@[i�u����e�x\�j��P��I\��AK�]p��������3���9��|Z5�����I�H,�������j������3��3Wc
:��'uTJ��A�!��A�l=po7��&� 2�ҚQ�ǆ�NK3��Vl�`�h�*�f��&Y�;S8�/�t=J�u����:��H9��_%�&�8��6����Ǽ���8��L�����'��x�t�<��>X�1�G�S��
���B�����m>�E�0c��7*�� k����ttIC%��m\����h��U�0��Eqtz�&�'��H�7,�W`�p�����1ЕE8���<�3�\�idΘ4�]sd%�$O!�������55��cG+�G`HmoK&-�Յ���mm-�x~O/>�=��l;C]V���W���g�y�u�G�V:E�IKM�o�Q���M�.XV��4��c��n�B�GK���t.������X]V�M�k����kX�f6�&���+��5c��[�#<��X�Í3�(?�'��O"Ʌ0iV�:ٍ�V�J��Wֹ΋	5�u�	Y�I&�3!-�)[
�H�G_�1�e�1h��MQ��]�:���H�K��M��kc����*N�u���M��g"3:�`�ҵYl�a�B��Q�;V�8Z+k�	�8���E׬ݬ�ц�	d��:�%����5�m�]��,�65��K����H�wk$d��fh�tW�ɩ�d��F�jg7���jQ4�k62�0��[ё������u�VěRF�A���i:�i&��3�k"J�Y��     �G=s�/q�Ք9ѕ�(Eм/�����.�Y�mq<x'qMX���j�k2�@�c�T���ݳ�Y�V;�(��էw�%y�D�`4si��60�
]�6�W�� ��v+���wp$Mw+���-eu`%�8ɝBLOW�]Ĳqף?��gu�u�U���q����Cr���.	�6��o�����i%/;��,͐!|�"2� �U��t��!�y�k��������W2EI�R��2�,Nc}�T,VX�a^gu����vE?7�uX0?u�- �0Yp����S~#�Ļ��ytlʚ`�z����j���'T�Tf����q��f�.��|��y�C�|�^?���t$�,��#h}�[\����(�j�<H;�����BJ����߲�5q}�(��������[�Ƹ��{����pӘ����AA�`���8�+}�Vl��B�R�.��}�Ҏ�tFL��gQ����s~O��׼|��0��ه��-��#io�4eC~��c'Z262�2ck7c>"�4��Bt���㽤-Uڅxe�o�'��uˠ���.���g�cP-�6\c���T�ύ�����@�A�?3_�^�ñ]B<&������VM�#h�M:��dL(��Q�BRF�	�Fs�SP.�s˪��>�	8����@���٘�B��KQ�lTzu���ft������U2Vb6�-:s����]�k&�s�<rd�Xڤ�_~�`�Ԅp��H����Tw�s�ё���S��7��ü�N�뷉)���T�f��
\��
>�<p�8_���"�0��Z��ڣ���i��S"���u�F�ɱMl]q2��9�v�<[�̘[���DSO�K����R9>[:e��ϗ�z;׌�cj���0�#�xB�܈M�X�C�������v���	
�����r.?�o��#|[�Tƌ��D�۳���y��Ȅ��'3�wD^u��tZL\>���a�f�֯5�Jk��du�fZ2'��{UӠ�L+fh���|�S'dF/;;JZ/o׺d��z2:�yؖ�F�$`	߷��1r�7}j'H�?v���v��:5 愣z��-�lm�U�!*��m�=��ͷݲ�N���@��e���96�c-�6��j�ކO��|���}��%�}���1�P!���G~�t��t�k�[Z��[u��;;#�Q��G0���_�>��3�o�LJ�W������M�@�O���"�t��-_�wx6;:�8j*�GZ�7�y��h�"��u/���z������ս-��cÓ���h5°h��Z�s&��}7��Ɵu�d\˩��M঺PKyT�7[���;1�z�&>6�'�z��pbu#6�ef�P��H��U����-e�6��Qf�H]�Y�i�ڪ��(ɔ~Z��ס�oԶ.���ΰ��q�,߲������J���ݝ���	��謗�\/MA#4��>��Ug׸*��Rs�^���&���ð�ك�g�üvc�c�%�_�9ܞ�c����{B��7qH[s�I_�kja��}��\8?��~���� ������	Va[Pƕ���ws�hJ�O������.��򊨹Q����e���&O��z�����6.FV�H:��g��M��&K��I)HH�0��d#�Mա����V3�<�A18\7R�T���˺36����)����72�����>�fY�˕�{kãm���LmxγYk����yw�r����Wb����+�1.MA�k+��5_{�(uI���X�a]R�UóFzw^�&``�5ѣ��\EMX��ׄ�7r����ܚ�i�s��NF��7�2�}�M��D�!RF���(ʑ[���u�C6|b����Q����Ƚtw}f�s��N��jbSf���_t�Fj={��'�f��0Fm�wj��/�d���fu"�us�{�����k65�o	��
vڥ]}�Ll !�g�-y˷���������4�E
�.�#�i���y��gd��] �;�q��b:��RX�BhZ�Ջ[���U���i��B�+��U���6]�kj���5XD���<�:�ad������b�4���z �Ӷ�W��Sld�,��8���-@�إF��g�^��F��4x�\G�f��6h��f{נùFh[��
a����
q��x����uU������ʽ,>@���p�)Tu{��ڋ]0�U[�����rwi}S�F��o]���[�5�<��{�=��\Xh0��&�LV��-�H������Eٗ�ðl���G�3!2�����L��Y�E�b��"��8=�`�<�w�e@g��єkǁ�܍w�����a���ܪ�p����/�v���^k�I������8�8R�'&x�M���/F���W�U����ݠ��ݲ~2���|���{���s^8"c�H%� �U5���棷�F��'��x>�����_���suDӾ�y�ui�J�J5,[1s��ܖ�٪�9j���3h�^=;���h�0Ѯ6�t+>�d���}��jOB���K=YO	G�_��k}�~��uzߖ�$M�-M	�EuHF�hg����xMІ�M�|�r�d��mT��yV�Z/6̑������;�[�����������Z�N���@P�{�>��n����O�C2dn�xu�c�ϼ�:>����5Is�ޜ;u��4��E Z�4��ڳnk�t���xZ��w�p�P�S�{t	G�0$9Q" �H�L8.s���>��d�N�l>֞�����P��~�F�j:Z7��"�{���J��4NeN��v��߽8}W�
W�&���N��s��X����=��z m���
�Mw�*
���T��^��!������h� �v'9>�
�-rN�pQ��i����(����)�y����_0ؼ3�֧�]Yp"�4�����ʝ�M�[�p�2:��{�������@4�t`�7xO���>��0���9����gijOhy�J�+W�k�sU��B�y��)�!�X��ww�t2���O7�+�|��Z�\�����hv,� �Om���1Iư	�#z:E�FV�by��k��Jѫ%|0I���0>���2���M]�AU�-�)�{�t<}^����W��]r�P��+J�8�q#�HbE1>"�i��&��G��ڶ�y!r�0��y�9H��=�c���
���΋V���{ey��1u�����rC��j���,����M�Qt�D����WZ����&�EJ�)�ޘ��� ���]K���s{��e�>��ͳ��Zx��#�&I��e�ʘ�:�Eq�t�+�ǣ�JQr1����/g��*�<�7w~"���-W+̈hU����J
���kW��aw���V7�8GN�s̩�Y_+^�D)�ɥ��$����m�%r�m�e�-E��y��2�x���^iG#�c"��"llUnt
�d|��)�ٹ�s?����ǂ��CGVw~�i�!�Tlプ������;Q�f�:�7�Dɽ�u	�u���7��7��ܰz��Ni�za��Y�w���������A)V֠ba���3ˣϐ�D��^��W�v����h�����P�f:�Y[Q>����~�dc�i .Z��
�~
|���c�x���បEB]6[1ă�� �	6���%�hO�W{�y*r"��f��u/���<�Tf,�WG�]畼~39*��T���B��c)�p����W_���+a}�=g�]�%��%�X^o���VI��O%���DF�-�@>�>�J�F+:�X3"�/76r�W�+H@�t�؂?^T�0���	�g��;��z&�B�4&2N�\h6e��¬Ǻ�7h�i6g-�b�[����L:���7�du�{ףWTm��s���9mg�Si_.ᚙ�����[f�6�u��L��eK�me��f��;=8�	�m����O,X_�f&�g\x����Ty�
.}pCE窊���g��D�Y>�d�df��5�ie�v����R�e݋ꉚ���	c����Լ'*����NϤ���v����������q2�|K^�ӎ�l%���`h[�rn�إ�n;�/}��[T=0ܹ��԰+CGMQ^��n//��ꮹ\*�SnK���7��u`��px~���bf�;�ceb�������\S�T�u�W��~N}�m��:-����!&l�YB�]Եw�s5�r��MJ����|�9�	S�0�����q�*��vb=�p�5j6|se!�)��b�p��^f��:���휯�ρ�����]m�]b�)!���K�<�F�+g��ul쓭�ݓ';Q�d�/��fW��׹ss8+�
��y{0���"����lt�ߛq��B�\�=z.zg�s�oM�.@�o�=܎[�F�̏{C�?�h�J�U��Zht��W<���8���H�G��w�L'����z1�C�vR��
�y��U�YJ�,N�����8X݆�`{�;�YD!���᠃�t�lMP�N�lX��խ��I�΂�V�o�{��Nh�}��O4�>4�$��������K�d{u�������J�-��M�f��2IiK,5�DVĭ���8���!,%V����	[-�ݧ.��$�M+i��g����N-�roԀ�u�oiۭ��V�ު��N����'l�{��<aX��3���o�%^�zΈ���Q���z���O� �͑�+|=109М���	Z7�U�>ݑD'4x�Ӫ���9o�C5WU�d�t����?|��K��"vON��nn���%i����e�T�������(~-Ĥn"�	�)�_����+<������>���\xG��Ky��5���n�}��dj?�C�vz��5Q��߂{Q}E��c���B��W�b�!3Ժ��5=����h*������w}����]a`M;˅��3(��{��G�����@G{h`�ɥ*	��_Y��e��\+��N�h���Q&e�{ �uP�i��uiι����é�E��/ws��ȷ�y'r4�um�H]Ϫ��:�KT�^S���F�E��2*��/��0�=3�&A��@�o�����Ye�p���x\���#�����N�Ty6���\�c�1��ܐz����n�)Ϻ�\�Ut�N�:�8���������{+4ai�Y�R<S|tcŃ[ě�$��Zfo�V�rd�ov��M[v�K�,�嫨)�_b$��_r�؋(_Lw���sPo!-���t�(X���%1�����.6��B̌m���ss��ک�+�/��UtA�I7�Ieĉdm��фX��i+����U ���R���}���[�ߖ���M��n�F������d"���6��nh��r�:�\t�d�}��q_[�]P(�z�-
pe{�{�޹2;�y#njn�!8�wA���ĴI��@	�5��xe�}1�-x��'�?jɉ=3����!Ρ��>qK�3:}���;:)��č`�-��B|s��_�FL"5`�F�R� Emء�m��e���s���4d��[���<HOW�`��RK��3s��ϻ��xXW5�6�oH�U؄�6c6צT׮�E_L[�����[��xo�V�6�r�\��/��+5��S	���c�B/9������"|,��]K��@nz;J���4q�������}%m�P�UYp��&�_����*�f�AWԼc=��1��w���l��8WAe�����+����;7�X��cg��9�.��&{.&W*j���-��0�JwZU9�J<���H�:,��
#]$ُw�Cz�TfɽB�˴�GsB����^h7���4*�}����z�硭j�`KgQ���g�߶��+�r'�HbK��T�=j�s�������{@.0+��M���u�'���o��!��F�$f*H鵶���L��.Ý�u�ei+ss�}��R�S�}}�9�I9^2���ݷ���؍�ob��,�Қ�M��^�U�������
��{U�y���ޛh	�0��%[��.+�L����]�]xn�N�_[�-��;�e�f�ը�����ʅz���(qq�4�i,,A��=VQ���W�ؙ�o?#FߨpY��ڗ%g��FNK�H��M� ��n�5��loJD& ���o*P��y72�r���ȱ����oc�Jn'#e$5	4)@�F1���e}R�{�95;k/d���ڸ�)��_I�Sy���o3x:��{���g<��d� ]'p��ֵz$M�\i���vp����)�'���ӷ��U~t66;��U)k���~gF�ن��Obn�ϰ�6��W�X��`�]Pq[�[Uf����-٭�wau��f�Z�1֝��"�P����6M0H�6�\2���<=���A�N�Db�.�#O����.\�3�v�{dh�ݹ� ͗���[3��M�����0sR����#\3x�8�#�ҋ�G����Kh�_Qɐ���"�٫�qq�B���[h�6c�	�$�#H橶u�	оv�W�F�M��ɵ��1|0��|��ZE�(�[K�ؗ���hkcAt�S6	-��NKU�jˏ�j����K�j{E;k��D�������[����nUE*��U4c��L,�<l�7Y;Fn���;�"�����n��l%,�3i�dH�{*��$�L��^���r�dg���Z�}5�x{��M�L����J�#d�Mr*"�x�Q�}�Z���|օ�lp:x���Gb"9=���w�\�k����7�9LBы�۱ē9�U��U��3��;RO��?���)�ū�iۼ��F��c�)��:�Ҫ�Yug*��Lp���	�=VH}}N��]g�6Q��WA�u��n����O>�}�����q��?{��Y}x�*wwD������q�«T�n����8-� 񳶩�s�W8rl�xV��tj*3��FK�F��rR���}�����D(������7�����e�S�xc�3矇��)$�(M5�w�0V�1t��C�V_O���n<�.U�>Yy�� ��GZ<ao���Z��w;�k@N�j �N��1Z�U5���jlW�t�A�C9��(u���3eZr��n�8�����ɨ�Hm��*�{��:���1ڎ�Z���������JgY(Rz�/-�T�j̰�t��FBwb�ͭ839��T�M��F=��╨o[��;|�]�<�&v�9���e�P �"t�f�q�Iuo{3gavZ'�9���9��ӕ-�ܓ)�F���6Mw;��3�Ct�V����{W}[�����AM���.�/P�ޓN�9w��*n�K�z���KJ��ʽ��.����E�����95]J�A���70sV���x�Z��k{���%E6�9_]�(w���/;����g"��[m���O���k�$o&��l.�v�������XwAF���U�X�Ϻ��C�ŋ��7M���|�P7[���K�ܥ/�u���{�ЮZ@��9�d�ݭv��5ϚPҶ��`�;*���j�3ڊ��\yr.���+ԓ_)j�XY�m�O2�ɫi9�F��� }���%��8�c���՛��ۇ,�=R�1"����Jp[Ι
�4�տ�?s��`��H���ö�M��:���=��kז�ر���Q��+!m�!0�p[V|��2��ʮ�M�V�<�n�kv��f�O����S(b�5����kz���ӳ��6#��"���:(o�'��
��5�[���K����xl�@F���F9&ϱ�Ϭį?8�p�<�e��d�3�qV�^��#�H��vI�я`ogҞ�z�#�sqV��1h�vã��"�(T@o�1�aD�J|�Q#E��.�+;��.':��{'�J"�d%�_�;���f_$�g��h?�*Dx����blU;�S~�Y5�bo��bQJ{]��w��4���G+�S��j��'�uÀc�e=k)\\���L�Y�$aÌ�~g�ޝ�a�SC��V�q\�E�N�s�\��༽�ƺ�{�����5V3��ܛ��#�Wٲ}�.=~������
�r\B��r�t�#�ci������]j*9U����j���OR����F��9]�Vҫڏ919�|�!<M��죳6�w�^����U���į��P�k���j��F�7����t��A�z�;-�P���<h�U�D���k7�.���;6葻�km-�1���p��c6J��]���T�rՆĆ�l̲���[�i�uIL]l�[-�ZY��Cd�ѶkI�B(�I�T�a��B@��)�$���R�e�/ǣ����f&�����ᛈ>��.o� ��G�cۂ;�0M;^���i	
*��o�k9?�T��W>Le�[3M`wbH�UW�sy_B�h� 陴�9(��ͽ�A��}ꧫ$����R�)���2(��c�t"㷦���A�GҶ���i�ͤs�[}|�5�C���=Z�>߆	�P~���ӽ�;��q#ZfPU/'�eM>ɹ�75��5��.�[��P+}eQ:��=������\M�zAXj����s�O�b�Z���Pz=<��*6%�f~��&X�ߦ��m��dT��k_��<�n�]6f��L]�Aԣ;�M_[�d���ʂ=*t��qY]$��9"������(Dޣ�J�\Lv)�\�K��:�ě~%/��gOL�Ƿ5Q1H9[��|�7�_1����gv�i����{w6�$G˿M������gRCR��9}a�A���P�ߨ����K}�����/�O��E���g;;t�Gx���Pi(�Z!��*Q�Vֽ���2떊7ù#o�|1h��]�C����
~v�����L�����\��d��*��l�qc�>��0�biwNHc#��a\�=�=���_\�FEvR��sb�d۹�?a�n��v���4zh�mqe�4�����8<�ێ�����}��}Z��7$%}9�?Y��+t��B�"y�p'���]q�e�D�;�� ��N�턓�@��~��U�Y�����C����Ѧ���7}�S·�*�L�wZ�u5�a�A^���Q�>Ӂ6�)��F>�Ο�zv�n�{�<0�뛨��[1������9��﫯��p�yφ�g����J�Gµp���U9�fbt��tך����U�1G�G���;�ޅ����6�Z��I�y�h*�F�)R�F���m��̀/!]銡�c^�&C�	J��\�o႐�{G|�-ǋmm����O��D��;�+-<��oiF�Śh�4�RF�C`���0�B"�`r>��7R&
������lrA�ո<����<�Ʈ�KU|q;�Y�6��W��j��c��+�/l��:.o.�D��*Z�����.�quU9Z7�`�]Y�q2M-wε�Ij��+7�ܩ�����T�6��gC���v��ў�w�������D�*h�;,к�uOo���gE��i��'H�y9�G� �I���S��Rꂑ��̰��p1� 7u�aI��+7{}XT;1�cw	�^���;�pnN,��%L���`�#Շ��;=MC�r����ny�ڃ�U�^=_����f��܎���@`��I%W���q�լp"8vʪP��,^Z����v;�Ml�z��x�����Q�rL6]
�׽�)X���;��B˦;��K"D��3!�XLԂ%�0s0/�V��\�?eĴ�5����z�f2�*}謻�LR���:�}
3�"aT��a�4Fܧ����ný��%��	�RรfF���t��SK4-b73���}�H��Bt�mk��]������L�%YՏ]����U��呹�e�Es�^B�m/b( o��׆R�O[�w�c�A�dɕ&A����B6�̗[]�B������X҃�̿��W��{�[�X�����3��@�}�`e��*���8���x�L�޹wSu��gC�7��qe��9��cE'<j���]V��y�S��U����Al�x gyX1w�N:vV�~Ω�y���I���Sx��˻�5au(8y�kz����ʊV�����1�]^@��s�8I���3!���ȓ#j.RLrӌ(�7sX��
�^���d���1J>��f��߆,ʺ�z*od�"�̛(�͚��u����
w�Vj��w|��'����:Y�=�0`�"wM;>��V��V����L.�F�x]ǈ}�U;_'��lUP��չUFP���څq�n2�϶���t���/p����;$_�03TM����b��E�\tZ|q���XR�=~Jb��m�\h5�a�%�p�(m����jY��(��kp7c��>��0�w�(�����B���Z(�A��6�<%ߧ�z]b�s������C~i��j�00B�{!N�$�v��!�O)"��������7��$�C������B]R�Kwʶ9u�F�݈\;3�K�46m�G�������s�_�5�:Y)��h�EշQqVH�-����C|Y��c0#����Z�/}5�]���d��fg�,��d�B�KWX_V:q.��ꜣ˧C�N��ȈX�ɣM�*b�0͘��Ikv����n�C�	���U�,����Gr���N�mVb���Z;e��j)>0�
����4�e�T������d<�iХ�i�[-�԰�b(��]�������e�C�x����њ-v�fM����mX�dJ:��+X�6���+6�Y�Z�U�m��ox�Ǻ�����c�ސu%�O�.���<6�W"6}�;8d���r�b��O�Y�:����6Ls���(���g�\t~���J2�ʍ�S��*���g1{�i�4:����C��]����\�|W�7���	4!�������zr����ֻx����P$�`�X�@X��B4ل�	A�T���(�y7���X:f㦲sMǝ�і\����������n�`Z�kٳ�<0���T�ӗێU���T/�jٞ@�!ud%U{�1z�'Z�2�N�[�w�$�CU��P�&{<�'}k���mE�f	%<̽b��Oh��MsU�s&h�8<c>�S4���6�&���Ѵ1����q�����6:���r�CBՋ�2I�(7�5��gfz9�0�\���C���u��nl @�L�)�ڡ*��Y�cW�w�W��%��\J������{w,Rдq$�"�)<�BS�QK6�����Y�6�3�i� kꁳ>k��Y��Uk%G�dW����n* �V-��}׉�UfR����ݞfʩϔ�*c� ����q|CV6U�����E'�9�w�~��L�$���9h�&ڏx��[��7��D\Ö��㺁�X��0�D�_:|<����$c�i��}��GV�}�z�x�KJ�J��IrYel/�L ��=��n�H�ܪ���u��u{���>�ơ��/�����<Mu��:��x�%ƨT~~���Ov<�V<��j���I�����́�ƋS��ďY2�􈥲VoOo@>H����
}����"q���ۻ��U�y�5yKū����q �}�3�j�c!�_���b��Vr&g|0�l.�%�W�{��*6�Z�PL�ʸ�V|����lG�Y��nL ��9-�H�M\yʫz=�T��'Dr�e$�g����|ܡ{@Z�&������jz�!G���kD��6��x�Psh�Uq�?���b�h��M��s�y.�c7����+�{�'��r`��"@�]%/3nx����W�fs)�˂�,@a�a�I(��e��F�*Hv!u�g�4���H����n���T�B��:緽=Q��ұSp�D�jk㙝!�)�_��p�����zq�{kU�Չ�j*�ou��������EF��=Wc�r����R��_$�[y��Q�]Yt�um
�XvڇE(�8b��40ć��#�g���}j	�SJ��X\O�b�0r��{	�y�s���ᒌDxP�s�C�M�e�o��r�K~ѭ-j��oxBS�����o���B1BA��!�q���D2(7�ƥ�wW���\#x�xt�^�S��-a�h��Z�!ՋY7YQ�N��&�pz�Ӎ��z�Ȉ%�;O{��ۊ�R6�2�n�dQ
��g�Z���^��D.�ܐ[>�E�mp�ME�.A��=(6w�En��M�+.�z�	���>��qY���{�Y<F���oo�켚���+��i�܎Ī� O+�%�� ���gMdͤ��j�����UN���d����a7������a����H�I*�M��ػhR���A���İy�M��V�ƽB��yQ]�7��cx^���啌�
���l��W��u�V!�@�5�S1bc�T��ң�����<�]��Q�v��Sn�J���JJfS/�\I�
���{���]�/�}��u��#`K�s`�KJJ��Z$�4(�pʉ�:�m\�z���S�w:қ�׷�)�m!%mj!�\>� �H��5P"�qs��N��w\л[�
�yu��i�
�C�kg.q�J�Y=[u�3fnH��{n&�<f��l����]{���>}���DB���j�����7�ḽz�:�9�-g�udu�}>�3O:�5"�e�ß�N�zx�i���![A�P�Ʒ�w��Y����ɇR�vV��'K���{�C�����kOj�4๥Ԓ�V���#��n |��*���Z��x�~D��z�#�ޕk��V��ϲudc�Oo�"5r&���#U�!`ԑ����$
�D`P�	S[};9��xg����8@pL��}+Ǧ��c�(����$7��gb2]tS���С�	��}�8[y��4�_��?u�S�8p�P�9+�3�<���
cBP2=B�3	��2�d+�漪!PH����վIC��O��NY2�͙�k�����Z�B[��0z���=���[���Gz`ɾ-��gL(N�iX�1�b<eq��w�T�+F�
fA�{VdL+� �{�y�w�����.�+�W��M���CqZ7���xI6��E���5Uۋ�z��y-YJ��FJo\4m\��'���V3R���n�#��.�=�ۛGc��W�U4����b2[l��5S4��7ST��]ԝ1J��6�[v�"�4��Ĳ]��4�:�Mҳ�4�La���Y�ѰY%a��Ҵ��٢B[d���d�$6��u�b�?0Y���M<W�3�{i[��yY����΢w���i��1��sb<����BA��G|�V+#��<�g�[L�ӗ�7��(��tY�鶡�J{V�������sv���
��KNt�,aov�d�W�!�\�}��d�&�.�쩌�}���S����z0��!o�?CI?ڔ��lӑ��a0��&(����w�Ćz�cF�z�Χ0�I��朋ݭ�ǩ颾��	���;��jv���?pH$�p������(S[���gH���oZ�v��76�=�6Ao`�)�n�����ŵ}���J��7/c�J�֪�x[�Ve�D�c��,��@�����sk��:���Rd���$5k��*V�NP���~�7�}�<ى�8��,]{����y���t��E�\���3dQ��f���o����*cq��a���6Ζ�{��M�����u�݅&c)ɧ��׶�4��Ft8䳽ƺ=/�ա_)�G��kǳ����%Z ��jJ<sW	����3�!����i��a� ����մލ�"�f���4�&R�6t�Zt(��n�Hh�<4u	��#!�7�}	%V�h��ꈪ�)yݘ5�u��*���:�i��2�:�>���a�81��XCw/��e���]#��,Apnh2�k`��0��%R-�aˠi�E�A
�6�$yۺ�叴Ykg_�4(VM�(Uܘ/�v7l�9vv�St���%+s4���cv���%S�HYK��v'�&���NAoj#�]�9����ϋ��m]uu�4��έ��KT�\+�����ʙތmI��i�{Z�;S��z�gA��Pۦ��><�C����$,�$�����ⳍe�y}������?-� ��Rd��DC�$L��z����3�Uè�9�b�;2�m^�S}_�T��۫c�;)�ʓ^`�>W<дQ�=����}��c��5���.�[���u�L�s���4��o�b���t=��fF����iߞ�S���ٌ���Rj꼨�l��N��+A�tS�QuG{G������sj`X0�t��nkK3Z�
�H<o�u�[d����o�tڴ ��j�a�F�����#�,�7k�NBG��B a�	y}��������?~��ƅkBI�RS׺�m�p��ݪ�okBiq�Y��#��5��빪�yjw��Vo�=f�K֬������*��	��ƨ��֋]36�+�3E�a@�a�.�;X����}P�.�-�Vf���R{���ܬ�E�.����]�-w	ƅ��W���s	���
��E�J�tua�5��xuf9�nì-[x(�Șe%܎L��k�1) �F�nII�	�7#jI!���9x�gu!��543&�8E�pE��t��n��%<��5t�V`ݖ��ך�m]t�˨X8��1�v��5�pQ$Z;��.��ȇ�:
QnYηy�
�[}q��w��>o�f�y��+>ӊ�����v�C����7Vj���'^�Ν����ڰ�r�����:�+�:X��WE7�ޫ�-�Y�S��=�Я5:._vc�k���G�$�^_ź�P<.��0��*���:Y��]l�Ʀ鑗������t��꩛�.�'@j���w��֋WG���1D�a}A`�uS��]RL5$1���!&� ���۟[l:��Va��B_!�E�=�Owy���&�%�a�������2j'E@�PU$�O���(Y�e�-nu���E�����nK�Җ�e�]x�wm�SƙE��2�(�����UE�#e�I, �l�jci6v��ZF�����:�fZ�wJ�3`f�lS�d�	dh���h��,�e�c�����F"��������g�<.*�Mٔ�myt�szl�;i*�F�]WfM&��)EI�i��xU�:��eؚk)��9!����FD�Y�J9�Ў�ZČ�&�,���#���[[#�X%c�I6p�t�������,-�"#����ጉu�d�m�K�H�"E�m�Xݤ����٭���JC$���K%K%�F�ґm�b�-��l�ՙ&���叒�d/�KԂ��4k.J�h��������X�ki]r�͸��A �`�nXV[ef$t�曦!��e��niR@�Θ�G��C�:/��t�F٦D�������ܰ     fff�s�mڷ���.fv�p�-�mK�UN,�s���Vff[wO[W�,�wr����6�ݼ��jr��c-R�V^@n�q����Es��N�!5�}��'�Ϧ��(t�*�f���K��n(6�]��N�x����J"��7f�͸�S�3�#.7�$ �jK���꥗��?��/�-�>��x}�Ҩ�`��k&�l�d�K�&��if��Ɣn��3�39 ��8]؝1�|�����r3F��!Z��.A�5T�m��f���3�ާ�}���w�ٴR�Ț�4N��[Q�����y�u��L�0ڥ>��6��3�y��;štp��J0�rh�k�j2Ӌ��d�M�W��ml��Fh����q=����ϧ��G�J�hF�R6�~���r�aoh��M�+�em=Yc]~�6�;��Y��'�}W�L�	��dsUפ�8#�J��nj��]kOQ̣E�TMo�~�N=N��d<��Պ��ESǚ;N��F����>�	i�����˨��+�3*'a��B���v���k$�h����Eo����p���iT�t���0$�{����Xz_�n���cf$�ga��d!� 2�Q����Go?y���:�q�V5<:�0��	��F�TU���{���.l[3��,�p:WY2j,$I�ŧ��ԸR���Wp�!���c���ϖ�N�Ҏ~]pє��7+f�hGC.-���&s��}p�ۋ�Z���]9͵4�����q#�rHT�Ӫ�U�EJUO��фEs4A��;�ӓ���j��W�}QT����[���U�N
�pF@�^�VT�A�@�*��&]�{X��{"yGe=�����~��'�/:ִ�F�w������iT�S9��ǣ^1Zh6
�̚�� �03̘%E�WI5 ��KzntQ���^�A	F�ۿ@��A"��t�:竖>�گ���hvꊑ֯��x�(�o�Y�'�
���{bw�����5�ϳת�)��<l5��x������<1����a�.�0�%�5yė��>(b᫲��>
�t$�6X����_�����z��2�]L��2�HP�:�)d۵�Νe-�4����ٴ�'<i4v&�O���}�S��cr9���EXٽ�ܡXFĺ^a�Mx��|{Ⱦ3��h���c-ɟ\�*���NR��> �H�hcTߦ΍���Ɏ���ӳ�9�c��J k4�gu�NQ��S٘#cfc�[c���-���/M�ˣZ#�:��:���ֶ=ܕ|�d]W��l7}��vSn���gK��L�˻��WLja��=��9[|�ީ@N�5���ŋ����R�)ou'.]�~�:��;��������F���ރsjk��p��R>��S�3=b�Nb1:s�Q�AO�L���=�?g�e��t%�Oއ�'F�������6�����>�V�9��ѓZ���o�YU�5�y��7�v��(M�N�*��^ر�\��kuZ:bu[\=��0�]�k8�r���q\�΃I�Vܚ��'�7\x�� ��OpsuڤVT� ���P�=��7_��캫��z[bcƒI�
p�_# *"Ap���y��^��:~��[��[�Q::�X��&���g��������F��^]㍄�O���I��:����rIR��3��C���ʵ�ރW��V��=��0�/��\��Ϳ���Q��,Y
�a��]��+w}��;�wKAL��|�g&SiD7�
�����z�ձ�:{�;MWM��S��4��w=���#2�<[�^�}z�.._�i���@���e�N���nwݙ�{gs�
��/�w
�yF7Vz����;DO��h/^o=�em�[�
Iر*�o#0������@�V���$��/SC��//;����k-e|� Ga�1�/�d�$(����"�,�Kmk�\хI�d)�,��,S�d���u�I�tՕ��Yn�.�Q��.��e*:K$��G�:��]t6m�.�&���mX�t�Ut�k]53[5����؉�$�i�Y��rV���]W�
�?��N�)�ޫ2��K�GO�{��y�sE��+��ߦB%#�!�|E+U��1�>8�R����ˤN��jF��E��;�BM*�w���5z�)�/�o"��:��/��^����ޤK�^=��4WG���Z�:쐎���Bxl��vں�[:�s3�iJ}�W]�d�#R0�Y{�-½:7�w�!�`���z�nT���"Blt�F�?f�\�A$5�ǫ�~�Z���\Y���N}V�K��+ɮ�r���j�W5.:�������^�TԼ(FOl�},?p��z��2�JWܘqZ[���׻H��*W����z�a�t��)B��-�ûB.&M��"�Sa�E)�G�=����%l긦�*�ߡ���q�U��"��D����Tt͝2}윔��t�Ayv,~M�mՑ�.�֜i�݋K�PǏ��t���L���5�(�fwN�|r�.�Ĥ��ʡ-�T;X�s%�_TUz��VTxcu�7^22�ggZmϩ��]A�N6�5��xa�o��9�TxN���vG�v+�Y�_��U�ʾE'��[j�<�Pme��r��-��.��������� �}(��k�k5'b�]f�㊒c�s���o�i���d���f�~�>7o'��Սn�|����+�jX�I�V����$�E�J��~]�"�ֶd�̠�*�R�xH�\JwxT�,в*���1J$�U�F��p�+��t+��l��ѽ1j_����Qϑ���s]�?$�9~Y�ix��<J��7E�:��&�ƣR�[~[�MCze";�ǎo�����F��]N�d�0U�'�lE�ƻr��FN��gC�}9q!��E����v�������S2}�Z>SV�:�ha�I� �/���e���s��q�7z�K���x.��K����H+�n'�>z}��>�����R:xY�����1�|�ޝ����Va�o �^c�WE):o�P�#\|_<ī��AL-�hM�9��Wd益D�s\|�v-�!e��7/,c[y�4��Rr	�ukPZ�_;�{��搂7F�U����Yf���%���߷ߐ}]��/�8���ky��.�;�#���9���[�$�ѐ_]´�uЀg�J��:L�T}hnu��E��O�ƘY7��Y�Jb5Eh�ϫ�mrK��p9�V��|n�g!#���	����7G��ݹ��1��uu����U5�VH���5��nԽ��y=���r��]w�2��Q��i3*��<˖c�enw����r����kF����U/{�Őd�7f|���a���d�~t�&���0�T_rͅ���Q{��q;�_����ۡ��B�!��l��S���h�}��,Dg����3}Ο-�P}�M���V�����&��{��\��Д^1��.I�9�_N���s8�GA\1:tޥ�5w��vk������m	���n�m�n�H��Z�㢆���/�~��{W��}��w�s���I�Y<��8y�5�#�v`��}dF�>��4<�;�ͦ���؄|\���D��CJH$�h/�e Ď
5 ��,���U��z��@� ��3���Q=R��arᝍ��n�	�����#;{G]��ٽ� aORԳ�<�x)�ټ�wٔ�7��Fl�9�Ι���	Wng��ea^���O�0�a�JC04d�o_Q=hQ�d��:gq�+JUʇE�a�m���Pշ�U�#/a��5m�t`^�Q[�%F�^��ص�pr�u�DZ-m�Xe�yث�]�Q�9�%:�ql��#�O�\��uvLN0+�}Ԣ!�pUL&�kՃ�䉎]��Ev�٤��º�{koWt+Ň"w��+���UU:H��6�p�����<�4�Pw��)��p�F=9�Z�����J�
�Ƀ�c��򾧻�{ٓp�g�o�Y��㡴�1�t���bv��<;����G�y]x��p3���.�3��8@U�xUu�*=(�̧��hE�~�m,���A�#��n������y�j!�@�g��9�l4�N"0�=F��$
 "m�H&����Mg��J��yz���'��#����{�hh?^�z���d���.Uw�Al���ۯ#ѕ٘vr�FT>�>Wu�Yy�׽���~0t3x#�Bx=Sj����+̌�7��w������:*ȇU&�Y/~~fe�}�tOVO!/jQ�F�]�k�z)�:����\&���NfUA�V�X2�EeM	�,{�YF\v�����_O~tM~�_�@bU3�S�$#%Ŝ��A՜b�L�[��{��㲌�u
t�^�.W��[8�vb�.���I�=�1%�s�!�o^�W5���m�['ǆBj�y}RgjW9e�"ZV3k�x=��N�mfҰ�O�-$2L)&�o�'���ƴ���rf��J6k4��n��u�Y��r���$l����$�&2m���e�m�ֳI�/]�3q�,ҥ��b�f�6[�u����f�� �ˣ$�IM�Y��m>�~�^�U��"�Y�-��V��7u���P2�Vǧ����:�z�+I�$�Čn,hl����Z�{lP�G��}��I|��ڪ��>�̭�ȲfCօW`Qw3Tu�TghB���O ��1���V}^=RQH���.3�K��Ơ<�0��v��/-���vy&�"�;�|�'e?�,�"E�*���zOE)��Lz_AdsY�_f��޺���<�9�X�MZsR:�k���c��#�n�:��j�b� ���ד�w��L�L�T9F��F5qo}�4h��u�׎c�%j��>\��pn+�P\6۱��>5�)Sxx��	C1��"��Ɠ�w����&)m¨�v)"�]8�<q��2�����5�5*q�$�Y�j��_��L��uZ�R>��| Gӕ/]�z�䍷(V�D^�����}����*�Z�F����>�5W�T���Տ[�2.��]��w�Y�bT��{A�oW�m�o��D� &﷫ٔ�S�����){�����V��v(9(�&131l�^c�y���Ns�w�D���gY���j����!\:����x!�S5�F�8���8I;�|�NYܭ�ݺ�����a��ȏ���nה�:���E_eW�^�=㝾y���#�9�H��R`7r4`(Љ"	�A��F�S�¸�uq�x-ŗ��O�}���_	��9�������Zs�.�~4��D郀+;`�ջ��!̨I]��d@i�E	
⮝������U��[�����f�����W�E�3	A2V$���{֮��-�v���Jq�6n�=�0�w�B8�/O�T:��*{جִt�[~W}+A/��͉<�/��~��2�쫞�o�M�L\�o�yq�<j�oG������1��X�E;1K=k��H^�L��[ܖeC)�ɗB*x�+̂>�f�B�4Z�pO���"��=ͱ]1�:zq1{s�b6�T!�������}2�A�R0�Y}1�¡7��J�	�^�2e���5���#��x]�+�]%C���+�?�&hT��P�!�h#m�d;8�9���ޯtΨ�=
��7GFw�m*8�g�V�/����=6N�76�S]u�Ҝ���,v���t�95bM��	�C:�e����gqnh�|T��wιK�I������9�Y�S(1$wL��0({���ٝ��z��lv��xwh���a��л�`�&�<����@����shֺ_(�s۶�|��5�a�ur� ��r��3��wݘb_���Q�Q���+����9�K`�I4�ni�XQ��&�[�oq�f����m���=�����y�#wTz�l�{�3磕ݕ����J�!�)wc6��v���e��](�����>������Ǒ]�+r��3n4�zi��ގ�$�|���rF:��Z�lp�TR�J�"���N�p�v�غb��T��Y��, ��{#z�/fCZ�6hcTqz�t(fe���U���[ƥ6O<D�X�u.�3�o,		đ#�5t���6Y�E�M2���s!����p��<Ѫ��;��N����u�3"v�.�a�;�/9�����ˉx��y�v_d�ܨ^�U����\(�n����ش.�µ	zs�j�HZ3=��t��=r<�ᚖ���yI�]�{�2�5�d���,��z��ؑm��[��y?�����g��#a�i��t9�&�<	iK5]`�|5���w9fw7چ���
��vշy��؄���ڨ;	�����V��ɝ\�x��`�яSNfY�Vh�f~�$��'L�� vۼ�ɤ5��R���p[��cݣ�CP���:��Y��zdY�i��
�j��^�1d_!�;N���M>H��{�U��(l�y�}˨�
��a�/in�{-��@Rm^^-7Pr응����k���	�^����*涡��ّ��Y���aI�t���˭����m꼻�f��a����u�w<Mʖ_j�C@��X7:�O/wp��N���#B"����W8,g��� ksF%��v�:���������:�=���vt6���O��c\D�-:�]�\���=�������R�j��5-�j�O�\��0D�����ٛ��³�<�z֡�zqŌ˹B�۔�u��oS�W?�"��KL"��a'zh�v��t�g]c,mW]�*A֧V���Ik�C�7��G��/T��ɘg"�Y���y����kmp�r���&��Gwl��7��%�N���Jƪ'Q�;z�w	6�FHtZ�*�)��`v�R�E�7{����Z�ӣ�TSbD�40  ��5�nٗ՚5�W�nڮ_�}�������:/)����V�� �����ۜg�t�c�ַx��@�9��L�9��:�dӈ)���7F�syp}�S�'7{�J�Xy�vQG7D��ԝ�R��u�z^*�5=�
�}z�F�j{E�Nֶ5�7���r�>˝:����v��v�S"YU:�s�jN����ۮ������������y�.�ƴe�x�oC1ɹ��3�Νc�,�k2�G"�4E%o��_$��To8�t�p���W�J+���@���v���"]�C�����$�@7�X�G�T���k�=�	�֗qF-#�E&%���z��Æ۝6�>D����{��O���o7��jŎ��lmng^�Fc�H>wk�W�+su�^NPs�Ւ�˫��7L��t�\lC��P���}�rsxWn�:=�����+�>U$�v��}:�)icS�P�����f���WP���8-�5��:]t�Pν�l$S��n�$Ղ$�����> ��/'x���z1��'+�L�n��a=�:�9S �:]�b��N6g�iW��ګ��Q���Q@&�ݷ6c�g��2�#��H.�.�y��R�;	�C����{�Ϟd%��Tgz��S����N�*G��=c�N���8<G���O�G8�����O���~~
1F~�|�yJ��S��V򫊘|**��U*�j~��M[�/F�ӕ^{��Qa�hb�>�T�H�w���^= r��k$����LW���������!&CA�Ӑ�!	R|C�8j.�`��Wf������ԋ]��y]uW��6#:���͡ND�J��VUм�n�gJhB{~Q���>�go�6��:ݺ��5����3"=��e^S�3>5�iR�������?{Bp8���89�v�n��c8w��ip��qr��u�om�2�Z��;St}tʠ�5t_	�[�c*p�:�1�B�Y�D+о��P����>���"q�ΰvZ�r���Q��emE�3�ewڻi}�"�򭽡wgP�GB'1�j�w������ȳ	͕	�z�)�]�b_c��c��̑���Z�E=W��p.yE�����4QX�S��!;��������$�Ǻ�y�.��Q�h3Q$c%���Ld�A��U@#��:��	��$Rʺ.m�����ڷb��^�I�����h+���1��K-ƱnV��+��\�(��$�k��~�tVr�u띢~������U8V\�P���WV�JT&���ׁ�Y8���5���q���}6��Yo~[��h�I��W�@}r⟗��Bϖ�H��ӣ(y����E��+vθ8���Q<ߝx�U����=\���5E(;��}�v�/�ߞ�^t<�ߺ�T�᭞F|�ټ6$R��)6���4\"��m�n�j5����Af9��1,';R�\�㐼�������v���@x��f���� Z�?\��i����X��{EPh��`¹�/
�%��^W��?/a�@��9i^�?k��!J�`}������&dS"�?L�.�~�^������E}�rW[��k����2(����n��G�M+�f�h������_�h�:���:�(�
�Zy=�s	h�+��a_��-in�֣�@�c�[�-�ǵ��7[~�V���X O�����4��V��q�{lT`Ƅ���g�*���9���Fҩ������P��CzG�1�DU�ҎS2C]�Iu�l�E�~^9.��h�Ӯ��7�4*r������F
�)ܾ(�Si�>�b_���~�fXLwV�֚M'Z+E�Kc�s�wўS�V�e��D��vI]y��d��z(N*�ʸW���iNa>��s�۳�l��hv����ba_9hq��WFhӕ�T�C���"O���4+��go��ik���/�m>BF��tԆIm 2$���c&H�&��5�����
��ǋ��P��&X�[s��{��]Gs����0��%(Vu�'�w���ۏn���w.��"�.�3<���h�J��1��UE~���y�~�Vgo;ܜT�Ӕ���)xl��Y�%�&(�(ڵQď^-�=QهE냢y���q�[�[���:����>A�)`'��"4L��V�]�V��>Ө(��MIk{P��O3����!dۚ�c�|�8 g�1�Y���X�-�5J�Z�иk}������h����{c
�U��z��)"�F��>3T'n�q|��Ӽ��v�¸��ݑS~ȧ�}�����f�t9TY��q§�RD���r6�w��-�������X,8���|)�KFN7b^G��A��9�u�űG�w��S�XQ��nW��ڃGC]���B3n�p���0A D�����!& �18�_��L�=�\Q��5�MV�$�Z�Tk���P��$-#� ���)�ػ5�پ&��:2�zwkC�He��wv�Һ��~�V���l��~nC��J�^n��\�6��{{�E=���D� u;8����:s4�Y��L�cS��t��G�*�?ֵm-h��Z�s4�7}ז3�nqV�։�k#�F����e!�r��c�dH���Ӭ%�G!���nF<��k��-��i�L�uJ�,G1�<�_�����z�XS%UQ�d\5m1h��=�q����y�3"��'t(�I��.{�?�c8�z�m)��hأ���%섎yK��ʼ���3���,�_d(eʫ�~ι3~�B�ˉz��^7o,{��k�4y�]�/���}���f��C|
�֞�r8��2}�"N�k����>��ß��G	zb�_��n�ρ�C��bv��R�j�"Q������a���nk���\�hҁ���ޘ���͹%؋
���^>�\(�MG���Ғ�&�0vVsA]Q�A(����Rv/jS�:��=_<�$t�H¸i�F�X�t�~H 	�0%m���P�gxs��s/��T�`?~�̝Y�+T�ٍB���.UIk�UR��ǃ�QJ����
�+�NpOM� `���q�A����.=��C�ˇ�
d48˽^ɍ^���P*
CH섩����s@A�.�w��0f�Z�q�.��R��l��9�k�_b7Z�(j���_#��ԕ̪�������Q��W&��Kp�n^�7�:\��}bs�_;����%W3���ܯ39S����L)<Q���Y�WC2+���meM�^�����vt������<L�(�J3i����$v�iYw'�\�����u�=0p��m��k'�Yz����(���!9�ӭ���(7�n�GT���{���Ѡǋ�����^�����|`�/�{���"��4̅����i�SF��]�;��1�=�d�&�����"������W3��Tw ��R��5'�Ffv�M6W���4�qy%\f�VEM̅;O�[X=����w9��ή��Gk�Ǔ���_��2
A4�$P��8	�&�!�jh�S�5R��f�L�����S�吥%�l�Y�0N��k����վ���V/�Ok���V:�����f�r�-�/i"��E)����[ҏ���Js
���d��4��p�{�5@�` ޻R�Uݷ�fWU���Q�A"��>gBwص8ս�o�~K�#�Β���0�U��[�#c����U���f�����X�@p��Y��E�2
��k�u]Dt��l�53>�U�` �q�`{�nn�����5�{�F��.�/����G�xEIrjc�	�P��S��K������%ꮾ[���A�7�"i%\q��l�hE�7����zV�ݝ�3f�t<�����:zRU/����3������K��4��A�f-�e��7F�6K�JM!a4��=+7m��H�.�l���HM�[��z۲�;�ut�5ViYB�[���2mk�9ūS9����F��l��b�"��m����e'[0f�Y����B�[� ��0�Q���!1;�)���Dh�����C�q�ǼhK���{#�!p�(�����#|j���]�K5�2��^�	{A��Ω1)��;0����Z���׀�N����m���4~��� m�b��I�	��3�1����GB����ls������}���[eZ�m�{G]DD�$���[�m�J��3))]��o��R��̰&Cl\�|G�vø�/�#�B��Z�f��J0�,�j�e���$9@�n=��[4�:T�yܯP7��T�١��~B+���_X+�$3�cO��P�������� /"IW2�ۃ���7cM��Tn�ѣ�S�\V����9��̍\�l2$u�R��T7��#�l���W]s͛t6|�t�������8w�#��ڧ35Rzx��+�0�냐��b��c#��	��S��C���f�p*���h��a�١������9��ʖ^)�{U���b�H�\zt�B���#�.��a�*?���:���{2m�3�E�0��g|�U`U͛>3��}?y�.����h:S��l
��㶯y��q5j�ӽ�5��1��Z��y��ѱC�:�8s��:҈�<(sƹg�96w���i����g�Ro�S�(�d���q�N��ٚ��}�]���������o�7�hԬ�3�wC�<s��Ӿ���G��%��IX��鑚'1�\߳!4�_�@�DpăP�i&�l��L����<���sQʲy���br|���?�$`{���!d������2jz���s��17�0��BI�;��M������na
(�S��c0_,���^�s�4����E���9[�3��͸���^�TIS�=&k�-�?M���khs.���;�{>� ��tŅpy��&�!^"{L�0k�G���33��Q�N��ǯ:�R&��]�[WT[>�a�J���n�`��A��>,�����eyM0���}����Y�O��{�8�0ÿfB���WJ`
H�G�|�[*vW��K&�1sP��pt�4I���ۙδ80��(�;�9>˹��b�Y�{��.>�5[wI���]�j�2�8o��1���K9LiÆ��₎��2Tl���]Y�5�<���[R��u7��D��#�1�|n�FP�ʸI9`1�� R�6ݡ�;]�8�U����^-�KmM^������Ҽ8p�+�a�\�`ؗ�m�}��N��B:��$D���6%�N�=�Z�i��fh��bǅ�-��{��W�)�M����ǭ��,�e�����Ҽ�͋�7ͷ�WvqNb"]mr�L++����ɕ3���o�C�
������.8鸥@V(�Ӳ�2!D�p�'�v6*ѱ��S��r��;�ܰ����1,���V��;w�9/ߘ��7R�_���i�1/6�x��#d�?��A+=���"�1�n����x�X6�+k��H�D�oh�04�tuld��j/��+����uh�ā�b��$%k�����LoKSY�������c��y�`��1�=Y�s&��pU>����d&�:C�m�
�{��<�ꉕN�bџV����S��| p{�0PP����'2�j�B�D�����f�
�}y\{��6Z�;��0�R���IؔOG�M�vwB�E	��;�ʔUbz�|���)X'������b ��:K�c�U�w+ 7.q��	�)��i?���L�
H:x��7�i��a>�zU�����V~��^h�W�sfA��(��jC��T)��3��<4�s�5�;��1����`c]����ӊ�3�y�.�p�dKE%�"+:�Fe7w�Qe�|t`-sf��*�JW��nt�0;
�M�h��J���2�x�m{Y�SWPHP���T7������.�X��K�W�N�i�̓z=Z�nN)�j��lwn��o��jFdbWC_*7�����sWdv����iQ-jl�ç	�����0�芘=���^��O������_~⇼����BO�R8�C��h�r/�)M��`���Q�.D�~�>����R0��3��w��o�q����,��������m�	�}B��ٷ��ej��$/���#���	�Q����8Cz�Dy�c�(�Ig�����g80�
s������}�2��M�5e��N�û>��]]��V�M��2c���䡺Fdr��xr���5����=K�3W�di�#�F��CH7^�����1._�׭�ٹ�܀vw���wv�(#uw�%Y��+bmzR\���xf$$��E�Yn�x��o�������ڡ�ͺ��8�u�j|I�9˓x���tG�c�G��ub6���kn
Ǒ5�/B��.~ʜ�N�����2�of��Acq� Ы�2���q9ʹK1���$^S��n�K��v������S�%�B�dm#�d�U�8��ڼk�P��CU\b���#�!Ol�ǲ�Χs�uԋNze��Z"��ґP�'�=0�%�UZ>�ϒ\$O�N�k���#iG���e���ռ���q9w5e]oC�aW�i��qH�J�)�c�),z�أ,���y'�6i�3�-�Km��PrSI�*&�;�f[�:^ê�H���ޱ�od=H��iN+�V��V{����ό�u�K����kBsp󮥣L֑噭��],fl(��LM�Ke�-���7jyt�Yf��6�Yn�Yd��Sv%v������5n�u�@�f%M�I]m��Zʶթjm�ٷ�������C-�ܟ9�A�_��s쨸�"L+5�	��3c>3o��p� {+ܾ8��������6jWs��q�R�YR@ʬǓ�΋>M�u�j�>4d	:���"�fb�yw�����]�ɫ	��f�	�QN�%gB�G0�n^a���p�P��F��P��t!%pͮu�5-uЅ�
;�����ʗݷ�"'�:���f ��Q	�-���#�ur�b�x����d��)��4%�Nî�r�_N]��wA{���x��i�:�&�	���Hy��e�B��Ets�
�/�1tjY!g�ϙ������܅�Gwx�vw�@��E���<���xi��)���NW��Q�
PD��A�o-ҒtɡS�BGr�����tG{�E�N':r(�~\6�U�핢{�<�{\��Jr٩i<�^k��H������'=�TA�:�W�М���d ���c+�P�1�߷��I�۽�ϧL%]K��TUR�5c &�\X�_n^�;�@��f(ܠ���p�<����D��-�ې�<iN���^�
y!�7�_&԰�ˑ������p������_)��ByoshE|�@�ټ�$n5��ڱS�]��Q�X�K�Rƈu�$;u�]�Ԏ~E]1M҅�aqZ|�K�p`��N���萓�}Q���f&�noꩂu��t��K�������;�������9�ou��c��������9�>8�Y��dӵ��1�f2�Pi�0콶wEB1f�z���X9�nX�We�W1��٠C���X�mCl�&l���V�+�rN���O���i�l������\ͣ�]<|S�Ɔ٬�!v�Xˈ�᛭���LRٷ����Ρ��Uq��3Fb�Ag�y.N�9Xw�y��b�;��o+�ے��h<�6h��DKm�)\��ZK:�#V`.E��R'���8�7��$o5��;��o��v<��Ww��Oh���#s��5w�U;�tO��9faP�>�0" k,g�]d"���y�^-��qV��:<.�[���ی\G��]F]�%ǒn�x��{w����-��W����K`��5���uMp��ft����u��AV��l����r����W�5�v�o��KK�|�㺼��ݕ��\��E>aӁ�ͦfj|&���,W�o����.�>�OCA)���=1o_#��;l�)w�$�m��1�+A6�48,gJxV�Xj���hr�b/������7e�Rg'`�X%�
R�CYx'���y��b�Sv�]�;��-:#6���M�9w�KgE��[��hz�v�O*��O��E`N�{�#|�ngqC$�dTC�Wl\�1���I�kA��u.n�^nCP�Ķ/R۔�����م�:�1��QT���z�J�����T=�[ټ�XŽ˺�w�i�����_5�<��E1�֟)T�,��j(<8�Wq�(P$�iup�O;U[�F���C�Plk�뽲�x�\�T�:R�!��]�o԰�Z���(Jt���{�AD��h+���4ݰ�=�)�e�+\�J�}Yu��\��&u�,M
]��xX��l�K�,NI�SL�S�[yG�:Ԡ��ԕ�vS����,���4���h<`�I��)ɸ�6�*T�D.��D�#�k����_&��|c����kI���Yn�F�Vͷ6f�����Tfњ�Yn���&ϗm���l���]�3�\4�����'������̻������m%Il2�f{�y�#e�I���J2.�����ߖ��M_$���XkJ3c#�^�[���-�2"�p7j۫��K�ύ�����a���/�W��ĳ7�͙6{f�IY�ŋucz�r�̴�M
�K!qt22]��ڵu����-Zȗm\J��O�j7F�1�X1��H��g[�Ě�G�Lݲ�*���^�X2kt��i.Y-�p��A�����A�qj�H��v�Kˈ^�Wt�BXY4c�M�!]�N��U�cMk�l�e�m��M���38ГRQ��j[JMFˡ��d�)nll����I�,�i���\��m�I�7h�n.��t����m������ks%Z�t�f+�[l���͆o:�	.�3^�+���)���J�����,�&���7d�6�Œ�  	$�I$�I$��i������
���P��U���k��o���nu':�Z�U|�mډ�[x5Q�*�ӡ�	�T٦,�t���ݱm��D^��W��Xn��۴:w\%�?���J�^��6��*߻�L�7y�̌�uw�s�^����%�[R��C�a1{�f$���t�\=�ޘd�'_�%�n;��ra!SnW_�S��{p$w>Zҵ����	單�%n�u�2�1�t0�A$��[��򎟼���¾���&�KY�}�<�s�x�����}��a������C���
p��ۧ��g�@�]m��>x�W��ڮ0d�D�^=�ݙ�:�#��q%@�.K�s�}!�R�PO8�˺�q�apq�K�$�}r��~A)�t��w1��_�*�.~�ǯT���t{����v�]�Wrc��7��k�5(���K?&{ʈW��b$W�R����=�A7G�[����(��9�/�����,�ޟV����)�%�ɨ
�Ƙ^uw�ߪ��	e�/��&#tv�.}�]��U��u��ҏ�S��n$���"��i�W�rM�.��:�Nc{��،ǞҩO��z0�6�����{7;S���΀w���6��7M{�R�eҢ��޺j׌�Wp�=�;by���y��CL3��_PyN	�݀9��w� 雷f�zt� ��8 _�O�D���L8��le�9����T&1'�=%YT2�*Y��b���\6�ZKRg�¹o��P��\&|� ��_'c�VR�6^G՛�uGjX�َ��u耺W=���՛���JY.�PJUJ�:m^t䗢���iV��+�m*��ŗc�::����{�6������v-�ѵ:m�]\2��}
�W��c+l<�P��|;O�~���(|v��z�l�T�J���2�f�(.gTr�9@-:ܩ��/�a�ɨ<�7�6QXh�.����C��x��k��^�a	��Н��q�鍊���CTi��X϶P{��s/.杨|:\K�P&�Tľ��+��g!AD��h�2�ڥf�'�ٚ�)�Q}�^��փoNu�]��8���i#[T�([#wǥ� �9A�I3,��5(eA���%%�L5X��
�+����{}�T�S>��k��|��k��
�F诸�xO�/\����[��s&>��yw��0�"�Ov?
I��2�E��<1�sGJT�i�U�a����1��gZ�7��	�B�'~͛)O��/֔w`�s���BT��յ:m/1-za}^���6�
*7�"t�z�]�"���.{����}[a�6PI;f�SF�sp�6.걨�5�Gp��L{�^��5�&H{��>��i�>��)\�\����^[���)˓���h+X�c�՛�w0��L2=2z����j��O�	3�t��ȨX�/����L=����������u�*�=���ߏ��7*\̿EQ��N;����Яfd%��1��a&�uC�z�ٴ���_����kVU��m���3���\П��r2�wd�U���u���M���ut{���{dŁ���G8_wg�,!	=�E�.G�Fa�k��q��3]e�ڮH�\n_����VΝ��g���"߁I�H�}yj'�p�)z��ꬍ����%�� _�5�	�����u��Nrj�i�>��(smg@�1k��଄�a{��D�Vs���J��g��@ȩ7��hq~1��u>�Q���Lta��)�ҙ*��Hb��j��|�xkw!�q��ma^B��]��?����)ȿ���j�r3�/R���?G�����ԕ��FE�*0;��%@'�etm�v�澍)���v��֯���V�LT =�Kfdؐ��.��R�O�).݅E\�į:�x�cQ��Bg��g�3�d^�X�Q �ᢇɦ�!@8m��%$}y�ʹ��63f9�9�ˆ�+}�JZ�)�*�b��߼�>���n�����ѫV��zR\��4���uB����<���sҰ�OZc���F����7���?�۬�n5ju�s˗'W�1�Bu{v\l�����;���>�;��hU�[#/�D��z\�M+��Xd��!��Ḓ�_��6v-.�
ܡ�|i٫�ͱ�x�
{wU�2��5f�y��6.0f+���(�Bw�+�_!��v��Vq�4]��	G#ڼt���A>,d�j�z�(�Q{�t�}�J��VU_OM��U�LÌtY��IS�|�w�L�<E��Rܜ�<���u�?MC���mf�
��X�(���ݝ�і�r�J[��s�q��.�M�n��/��ѝ�p�Byh��R�颢���-$$��.&*"%���J,��GQ�m,VZ��.4��m��n��[o�I�J^i�2m1.3$�q�ћ;���:�]�%5���#c&�E���Ib��z���"RI$�<=.�b�Ỽk���X΅]s�۩��m�1���y`>s�t釈��J=�N`7G�ݺ����֩B�Xx{i��p�$�Z�gz���7ǆ�z�#h�t��k=9��< �߱%5;7F�0��w�ye�r��ܲz�zI�8���3���!�X����	��S�P=)�d�dS�^W.w����bR���c$Ŷe�I��)IAÀ�i�!�g��0�H޲2�������ȸZX�6M�bV���-�q�� n�(w|�8�Yo�wG��)V�:;:'����+�ߕ�� g�����E|eҷ���W�5�l��H�,�n���� ��dfD�B���Ky����Bv��� ������@�U8��R����[��;�w
C�33}�()	��PG�r�3����ŧ͊�D�Y]ؠa�M�{�
��)�sxU���#�8Q1�Z#�C����!�p��{T����y��_���o�{+�y�L���:���s��e��(�������(�SF��{��\T����{,5,��k���C���y��Z�啗�7��f��2!��|mϭ���ՃS���R�J�դF�;}�Ȥj�Lo�6q1��P�{�wq��岳�,.��m�ҶO��c�9Q@Zh�ت��We�F��S��J��=���z{p��&�bްqi�7���vo���KЇ��3z�����.lz_�d�CR�N���mtGxjJa����=3�+޻�a�6��-Ny�={7������BJN6�a�k�K7`݋����x����p�\�:�"_�����Ř�,�;�l�h�u��!�H�?b�PQ�߳t).�p>^&�=٨��o��b�a����W�W0���K'�lHkUw]�;�Wte�A��F4�''��tҒ(�²H�;��;��c à(�Q������,��s���	�}ϸ�0v�iw���-��6�%����ܵ�_4��B�ӍƱp�γ�F�WZg�}�����M��/r�h�V1�p�Zg+�L{���I�4cYk��2�����J����ͤ���v ���A��扱�g���B'E�Z���0G`�yx)X;!VvnT�&��YR���3Q%f�	�O��]G�aVȫ�����h�5CE#*x��Wڤ^�j����+��b���q�x�}b�
�aO��e�r��*��x��ś��.�8�.���|;��˓�1�[��u .��$f���M&��ҹւ1'�^��������pfw˜'�Z���E#񂖻6*��5�����}ھ��&�c[�omJ��`���Dl���T�GÖr�W�I�3�,s�K�ga�f�Vv����#�o��j5g�Ot{�ݕ�Z��ֺ[ۭ�\�������9D+���~%�1ҖBp��K�d�k�U$�J�����׌ɧy�ս�ﰡY�����ݲ����\Q/T���m�BkY&�v�I%�������	3�m׆Nn���ʱi����2�E.�Sp��ӕ<N��(ܵ��9rIŖ��ø��ng�A8=$l	��^���e5����ep)4��EP�,�[��j�M"�j�' ʸ�f/`d_��_�^!)���ɚ�q�].$W��ƅå�,r�ڽX����u��r*f��3��l^��U?Z]���fɦD��Y�L�A�K�]�GJ�/W��t��N�fV������Ϋʎ��fԺ���dV�0�O�.g/cy�H�Ce��F�6��C)�Mh�w�T�s�r�=�Uk�jD�,���F��8�N����SS���GS�sk���=S��î�UmU�v
>�$�.�S��O������%��b����_�n�Nu鷫� Zܰǆ�)�ؒ,��L�|�G<��.�6�Z�ƅwS�v>�f�yV<!���>�ˀ�GaK\@K�8�r+�j�:z;�!�9nTJK�>�mv����E��M3)�]�>�k��m�(g,Ȥ(n����\=�]�c-:G`�pYh�%��˫��w�sN��p��wCT�eۚ՘8���}s��(]s���N�mIw-탹��Ύ$ϕ:U�R3�3~i�87A��.�I;w�b���}�Փkd��m�:�2&5��4�a��$�.<{�)L�{7~g']��޽�����b��R!�:w�:=|8�ȣ�5�y��@��r�෣"~���-���}q�t�'w�m�e4����mן��%OD��R�Ќ�0x�K�\�xCSg`Ҭ�&!9�3�7a�H�$�7ZȜ��x��xn��'�~Qٖ��4��������U�C[k�e�=:d�5�^W�n�!���z��Ēe!!0 d���'	$Є�/�P�*�}Q��	E�]$x`���z�Q#�yAD�R>^��ML��+]R��9�tp�p��Z��C<<������tY7�q�ԫ6"2��|x+d��g.��9g�lC�,T�ȗ'޺j��O�I9��_X��h-�Ίdep�T�'ɾp1�T��^U��y�^X�������U�ݺkD ��C�+
KѸ����h�	�v�4�22�j/W�p�;�J�Vp~���\-�����w�N�W���GIY���/s�����g�n�7�R�2k��x���G �(K̔���:�pyi��3v*VV��aww�ݕ�4F)V����u����i>W�)��Mb�/�A����;�ov�Ѯƍg)T����}�YL�n&TCL�������z��!#Hit�ŉ�`�VX�]pݷBY�5�k-&�\��r�m�t�k���t]m�-�MF��&�f�%$�\���˗beSm��4�Kcv�f=��[;s/m$J�K���+����P"�zxYW��!"t]pS
�؏_.Nۉ���DǼ,���ʤ����p��\�B�84gΧ+.pTS>s��m��?T_����=Tu�^{��B�x��ɛ3��H�@�Sɡs����Z����ޫ�OK(�9`���I�ٛ�����nΛ^!5鞙H�m�O1V�l�u���������8{lNƭ��gA��Տi&]�<���@��\I�"��4pS����&���td�Z��
��~I����� ��5u���������c�<��.�ޜ������}Sa��`�.�8���s�(E*�{��E��ڍ��\1�6b��+k~\��i{5u�	sI�XÇ]�:o�l؇��G:�U�g�ۏ��%��t�#|bע���_�@��t��ڣN4s�w���P�~����m��b�ݒu��X�pE/�v�/���ج��#���\��]C���T�98��>��*�z*�l<<.�b|��F\�6��!
��+�Y�0�$�[C(X��qm}� ��q1ҕw{�lh��{J��hw��Q��U�O�v�6���g*�d��8TԻ4[Wo!+V����}mQ�����}���Ә���R�qf�b2I��'-���������W���}vin�373���*�}��]�'G\Ю��pp�;�Az~	{;f��ִ*�W���C/����r�a�ց:���;/;��oh8�u���O/|���P���(��h6R1ċ�"Q�Y��$C]	���D�rTKB_�Um�� $a:0N�~�f�3Vt(Y���md�]o]��2��w!��-"wS�d�U:����u9�-z7mI�-ȗ����+�c���my�\�W@>�ڗγ�9�ZvGzc\=�X�ŗ�Y�s&h��`�>�;�ėo<{��#8���.C.~v Ot8X)G�^r�%GRG6k��օ37Dq�n.�<c�8ݒ���y%�&�(B�����i�G����Y�ö�w�OƼ�*ڢ�"�Xɢ�Eʷj<6� Q�k�3��ƅQ�����Y�s���\L�v�ܨ�J&�@�����ʼ��b��n�&m���I��E�P�3� ��f-���0���v����3�����ѹ��l�0f�vG��Zu��	��ף�k����%�J��If�h�	4nKd��27�����Z^��������Z�P7��bE����,�b�>Ж�}5��Mm{�f3}����<���K��r	C.�5E��Ӱ�F�4?<�,ܣ��,��+�1�w�:��+;������R^��+uq�y�mw�9M"�j�}�-w����*k#���3�5@l�4F3�"����(ze�<=Ӓ�oF�~��|z\���ט7_|N�ݣ|�&�gD��ܳ�뼪g��JkD6�/�yIom�X�"�j��=�Z�J����F�~�>KOϴ�t3���˘�f;�M�q��-F�C4.,�>5���1p�,�!%ண�4�{���U1�P�% ]���}\/��CLNP��%}�(W���=�0�T�:N�({��&�	�h�^������s�c������b��<�yU�{<�fHq[��;�>���u�ZJu.4�49���g=I/))��
��-Dy2�	u W�u\}����%c��?���òꀆ��,1-O�x�"^�s�璻S]t�ٲ0�Xb��6eN
m^��f������Vcl9vÞڛ:t:�jX��28�g��f�]��i��yj����^��KG�vw�!/�w�&���;���i�{�Q�[c��N��� ��OQ�@��Az���i+���ۙ�C�L!�r�r����ѱ����]g�\/q|�7Ԥ)��Y^�ƕ3���~�6��o4GG��W�[���[�U¶5ƴoZz�@�V�T����Z톖lN^Tc
�����%l��vger����7M��U]_��9qC���	��F�ߗ��ww�=�q���������T�8 ��I��w���ww )� w
w q�wwT�8��x;��?�{����?w�ww������;�����q��W��g��������q�q���9���_���>�����廜��P�k�Tk�Om�bE��n]:��3>�h�-�d��vV�7z)�"���o5-���Q:��l��R�Wk1ђ���w!T��alفk�1�*v�n�fӫ�Ӛ��_;#�7�B��Z����H���{�w[w�KZڋ^����ʬ�I�ͩ�7F+Z�-���Qcd�SX6���	�X̲�X�{3]Zxv�2 ����M��j\�k&��R�*U�j�,2V�cAT�EV�;�3X�����-��4\�Y�r�4�ǅ�I�F�i�?�;���
#��<���6��Kh��/K�0Y�R=�UlCJ�7zێ�І0]c`��Th�^:h�J�gZ�Z5Ԭ&7�ۤ6=�Mc�SP��-=����6��\y���Ցz�H�4��t�ɡ�УhX93�ҝ�g��J�V����۽�w�N��E�/V=��m�(��!#[���,_1zXL�ЄQ��F�?MMJ�)�6�-���ZѫabP-bB��D^���
�J���1�7
��Dĺ �6`[�h�cRGQJ�m�Qk�N[�@��'(��Ǫ�@����,�Z��ă{I�L�	&f�����ڻ*�
W�
�3�*��Q�*�2�I3r؆^��Mn\��[�)CJ�N�~-��1S�v��2hfl5�ɸ��㫫s/%�H�OX�!3��Be��#�,ћt�o�5cd�{�N����kK���h~�,����p��+?;[��u�b�H�)�"�K[�50%L��2�ݛ#"B��*�`�p�T��o��Ȓ���`�&	[Yw��UZ�4Ԓ
�L]`-�/.n�F�OVa:B:��$z��M��R@CT�v$h�ň]�2nɡIL
KC�l�\tIа�?XL)��Z�˺�n��ma�[�N,�e�om÷�IF�$ �p�]lܤ��R�6cD��QB�n��9fJ��?�q��q�rw �wp<��ww ���rwq��w��������q��<�=��q�����w!����o�����wq���|?����n�������?��۸�8㻼�y��wq�����8㻿���wq�����P��;���;O?����|1���;��~�;�8����������wq�����ww����/�?�y���������?�������q���RG��8㻽���?�����)���\"��#��0(���1'|�y���ԥ=���=jc�{wy�x��("$�w�U�mU�J�f��Wv@�B*����
(T��m�)�($�ZUQ��M aI (�̔�m[B*��kV�D��ͨ����h­`�Z��U@_l��%&��l�D�BPJ�*AT*Tڵ_       |����� H<�����b^��  �  
 ( �@P1��
����öҊ��wڶb�j��=��Yg�'tKH�(�f�����F*�A���ƒ��JV�9�Sl�4�U*}�޻wZȢ�Zj�*iZ��)	C�T�VUlj�M-���B���li=j�3F��;n�>�F�����[w��
 v�T�((�{T��Qf�72�C&Q]�U;H�,�(��R��I%V��l��lM]�J�D�1�n�a�Ɍ��f�n�l0�ݺ����mݮ�F����YT��٤���4��[�[Uۭ�J���������k�����;�D�.��:7l����t�Sn�Դ(�-u�Lm:	uwwJ7�eu�"��]��δ�*�"�RT*��kF��^�����[wi㶵c*�۷j���d��X��ne����6�l��u��˛��.�j����AMm�U$N�]e�]�s�K�Ƃ���T�"R���ETV�zg��{��uRe]���j���9���V��E(�d,Ͱ�1���F�XP���ݶ�U�����z��,��Ԅz�����+�k��������4۷"��d���M�j�v���)�i۸s��gl��i�ٜ.�\�ǯT=
�vpb�h��'U�֜L
�T9�ڥQ�A�����ً�mm!��I�T�������WmWT���]:�v9�mnf�t��[���wan�Tc,a�
iiݹ�.Z��S���t-^��@+�0����-Z2�çd�]R�ۢ���H�`TT�(VեCm�V���Wr��]�GZ�*�j��:qݧkv�C,��ݻslg��{mf���V�
ݒ�WUw(8T���N�p��1V:�Ӯ���
%*+��ڧ�P��cz�ǥ�����׋ڀ/]4z�8�e%vt�F5LR�(��c�Jk^��ҝw�wU�뻵\�7g]��mˊjΗwwQw[��[5�v��ED��� �;mn�;mk�tжt�:,Ζ�6S���ɶ*2���ۥmCV��W`���tBF�Zh(�3�a�s:�wt.��ݸѰF�Q�C�Y|����)R�D��� ����J&@ �{FRR�@@��)@��  "��	JT @��SJ� �@�H!*�@�����������U'��\z��/t�����[���_D�ή�u1O�:�q�<��304�y�����HN	!!!�I	$	'��HO�$$�$� ���|��ϗk.�j*�^K|��Ji�ǹX���q�"�rf;t(����Ձ��`c*I�0�6*���m<J��7v[�]�Ñ&�]�,��d[u��,���zXF�O	g^�Y�T�6E�VʼY�%�)K�C��!�/]��(E�ss "��0dG�+�b�Pª4j�#R��ZK1���d7N��ݵv����x��dbV�1��V/H���CVAז�X�2�4�&X�J��n��4�� �~�������$^`��q��.��Bp�KF�#c"Q*ْ-n�I�����l�Ң�H�27� ^b�@"��U*���-�Kc�f�������ejv��5J`d�[V~�:8�T�`H[V(�d��ܒ��?4Ѥ�7*�
������A�KJ��7v�z� ⤌y�g�JbPJ�46�ZiV-��� Pi�wt�P=S	�E��d�X0����!d2V��šk�{�=UY.0���1������$hVl,�ĕ˽QZ��kU��i*�ݱ���f�4��q'Yh��ǋ_�Y�	l`���ȱs���^¼�� �YOD<tl\&���T��\��-�Vպ9CRBlu�^%���x�*B�����lke�����b�U�S�yV�Ԡ��&ĥ��V�Z:.l��X�ץ�:F�m(ֆ�y��EE1���LDU�t�'�����c�a���l���h�ZkU�RCl�4�7Em���mŭ��.���^X�I{�W����ڃ�|���HM
"�X��<��Ǽ�o�j��hKxkm[�����A[�"�#yV�]b���YtV�+��v�%�X]IP���u���[vG�����[Y.B����?^���%b]��-\�h�*�饭]	W��Lͼ{�s�������b(ň�*"VT����(����DDb"��
(���_��M�)�q^[��a��b�aY�V��" [Gqʰ�;�M�^(�:-�Ͳ)����R��yj���*�!�7h͋�mɥv�6v
��J���Q��`�'h�9��4`���Mڽ�ꀢ��q㵙s�O#n��;�vH�/V���NG���6�`�̤ݚ�S�]�I��Z�Yd��( !���]��G$1�`p*P��'W��݉,PK��L���Ґ�7V9~���EU�ͯ���B?K�!�����SJ(��-�����N��5���~HV2�E�R1aK�
x�<g����Z�^R�`)�O+E1L}��VZ�� U|R0# �2"���,H��(EIR(��Y��2P������5���M�5ofh�-���jX�fX��O%'��0KG%<1��V�+sY�Qnf8[.j�8�֌�X8i
^�h�X����vf�D�G!܏3��%�tfӂ�E�o^��JQ�N������!�1�&�ö��x-��(�,V�dC5;Ԇ��i1�/K75�����i	�Ƅ㧿H1f�b�d!�a
*j�f���;A6��+����e��d��� �]I�/ I4P��y00�ssJ��$l�h`8§�!�bFEoBZ+J�@n�.��U�ݦf!���9�:��6�f�LF��n�;n扴&8�lK�YLl7x����yC0��L�����Y���ۻت״�ޝ�`B $Y6aZ.�wS@���eS�t%���7s]�D;tc����V�ܽZ��8���{r��5�(��.aD:�FҐ�7�FQ��y������Y�cZ��;��I6���gיcDb���vj8bB���A�35A�z
S]�r$E��zܫ�L�i9��w��+DFcQ�M�f�e,7�KV#��{����0��Fʧ��eؤ�<�e�A5k��J��0dw+nJ�N��/(Ҡ�YKiB���e�[W.�i�Wn$��ZA	ޔJ�SHݿ�)�WF
.����-��Z��L@C�=��2�C��,�%�A)�4pSИi1�Sgc�����uj\3���sf���|�3����/M�t�UdQ�*�sVm�\�^�E���<�ᨉ[�+b�y'v�l�9z�Gh)V��^H� �6�_�9~*Q��r�O�8�fD�r9�X[J;F�5x���^�]�4X�����u$�.�4%L���e���u��`5���&R��:7��(5������	�;��S-ԧ�A��T�]���؜�Va��w&��\��]�_:)�@;�$�d!DEbEX�PU�V$DDXP�q�"�$�h"�#@
�I2��3Pkkf��,b���5Pi� ^��K�F�*��g(i�0ll��Ȗ���wLش\hؙ�ʓC D`�t�Z�T͛�y˛�p[s6��&F����YM*l���V2h�x�Pz��ʰ�F��B�Kk7h��t��)\��Gqby-n��2<��������R H�f�ͭ��K�Qws3g�f�*MDm�L���e�����Dxv��=��!�\�6`8p�v�i�.���-�ͼ �FܭN������+)�t�%LW���Z����˵V�u��=
�����Zא�wB�FSrakQ9)*�˔]*֙�ƕ�$����M3k �^ϕi�՜19�*Pb��\. �p ��JfBk112�ܼj\`,GFci��Iq��^D��Cl2�lB^S*9;�ޤ��ڱ�X��%d!��h�|rٻX0��,�
R�ږ�*���0w�����f�P�+)RhJ9Q��! Y�˽9����(�Yj#�&���Tյ�j^|��j�|�h�mI+]�h�F;(�1��(h�B�BB��⡊˩C4��d��̿�(��R!-��}�F1V�$\�(�OA�0�ͺ���r6LmېX��w.�;�f(E���-��`�S�X �v�v%��{Ofm��'6��f&vn&����.Z fU�N�SPv
#p�Ma��k�{�4lolm*=p3{�-��j���/.c�p��Q(o�M�KS�V@�����B%hسP�yX�2cRh/*�FϬ7L���g�&�X��ʨ�"+.�,���3�`���c�$�l��eb-�2�R�݋�$��@�2��]�Q0<G�A �`��B)H�$����ZɅ�v6���V�f�����[
I��EY�=�M'��9[6�	��T��yB\���>a�������5��$��d�tw�f���ɓ �l]�a�{*��w�B���3BV`��YJڵ���
��˨̬�sr�b��do*!��DvC�*̼���XUV�[5:�ںKP��z���k�΃<&&jа۪"�L^Bܬ���>�`�ǚמsW-ѿ+��1�Q�͡,
��[tV��y{K��@,��ż	��Kt��h쿖dV��&����s�m��CQ�H�"Qu�L�b�A��b��+�*m̄�B:6��p|�4=�5�# ���>�P�J:�x)D�ޕ�*��kq�s6�f������Qg$֘���6^�S�˽I]䧶�أA�$J]*��i��Tϣ�+kA�=U��'!�I�4sn�r�#)I1�.�:�'�RZ��v�XB��x5��l�Ԓ7�0%Q�d5j�A���,G7�d&�u�b�"�m�B򙰔k��g-E-�0���*��5�u�b�ݼl�EEBc��te�h��9�q��py3J<�g+vE>��:
�v��TI�;zD�e0��AF܅�c�Ao�.�'`͙��<:m�	�-E�D��YN":��ҫ�j-[�jpz��
ۚ#�9oC��;�Y���	V'%��8c��S�+G]	�e-6ػ����^��[�c�vk6kj�*f:9�h���)I�[R��bE��f�N�2�fs�U]�K��S��6v�]:��ň<�qj]�Ck91�]���kÚ�y�iyw�o��aR7�F�M�My1�w���ha?"�X$�X��2:�Y�޺Ѱ\��jIw��P�b���OIj^����ؽ�x��sR�Jȣ�u��]��պ�
��{ԋ�M^�U�*��Y / ��`1�gݔTNiP�Tݼ�d�}�W�@��w�4�j���E�J��Mm��wN��֣�yB��c�ACn���2Q(S��
�.*ZUagp�K[�-��Y�%�7�%��L��0��@�x�V�=f���U�>��c �Uҿ��
�0��kks!L���0��5�Eݿ�m;���(��Z��٭F7Zڷk1�������n���CX¢��9��mRx5��Z����)�[�d�4(���ug���;nӶU=���"�]l���Q��k��Â��.������8�]�١�/.�7t�*یi�QnaL\b��ܧ[��݋��W�-@��wv��3�(:*x���S�	Ʉ �R��N����f���4��f����֢��/(n�rL�������Z��؉K"��� h�^\YY�����ca�O)b�����*�lr�QǤ1WRD�Y�������h�g6en�@�JM�N�3B8�ۍ��Ƥ����lA����恦ڭ��"v�,l�6�2�b��N���D�f'@Z�&�z^a��ŒS7t�=��N���:v�V�e�y�`Q��)]\���-�'��dckq�*�k�(�X�-��%V����,:�W�+7鵱Jƶ����i���e �n���ٺME�CsP_A��K7e*[blIk�mRĶ³`�����4�uL�)LJf�)��x<��oZ��SI�PPD!�EB� =�&
���[��:jCOP�c:,	ﾫ��� �"��n���y��Um�۰a���7&C��a��Z�ƥݕw��&\��TT�GG��|�dם��M*�B�s~<�w���|��
�AM�f9I��9bfZ�X�⻬���"��4��&�2���M�#!�lnC�<���&� T����DoQۖ���x�gtau8��Ѵ��.xs/d����\�
e��b�0U�nc�Qn��7v'�jI�&Eb������9�40�&� ���OwMl�2�FlHF�`���"�m�u��2��̜
�n�
ڻeI6�OC(cX��c���n��SW�ܺ�Xw��n�L-�M�h[�-��ݿ����v2���LA�M�E0���X����:�V���)BY6��8�`�AKpͼ���	���-ְ'B�"�a�i���je�JF�3�_�����ا���d����[��̎��њ �TY�d��wCA1���)P���
c�M�
��V����VC�[Uq�ŕ�� R�C�y�z����+�Ci��8�J�s1P/(%H�P�Z/�jP�.��Dm2�-g+o!�W���0K�l�٬A�n���1Њ`�+(�x ߚV6�b�{m����B7u�lj�Q���ĩ�zI
�p�˚��YW,��,at[;��A\zM,�(-�+,�y�Ѧ�e+ҕ`3IY� 3��P��o�TD�G�Fn�Oq��;V�b�鋽�m�AVf�	CeZy��pAW�o]��B����5�
��M,�f�mbn3�Ҋ�9�%_�]݈Bb���������h;j�-:E�%Y��4.ܚ{Z�kp�0�V����܀�SU��R=�-�����HV�	oV�ʺT��%L;�4(�7e�U�zJo�!hHL^��S3S�fEe��R�,���7ne$�3����n�zS��n���� *� ԅ�ǒA����
 ��H�.�Fa�̑��n�dt����s ��7)�N+)�� �j�U��n2���F����[f�6)�;gt��[�Х���� ���)2�囸�l�#]m�[	�"qX1L,@[��U�����S�/Aܬ(aV0��a�ۺ�S�FR��di��k�m�V��������X��A��K��ss-㛤����S�P�ѧ��9�`����FB�Uedd+��^�D�݂���a1^Tu���ލ�h���[�Lja)���%&PU!a�&��ae�����EKJ����Q�zm2�K(�0j�/C��+a��������~��C!XF�&P���e��̥X�+�Ś �0l+ڦjai�)��Z�P�@&����+u�j��xlm۠�8�ͽ�w(����8��1�Y$V��X%%V��V�ĉ�_�*�3��ܔRd�W�&�+�Tn�����0 ���d��Wwh�-��붌�P�9���HS���*Υ*�j5n��,��x�Z��F�֊?'I�^��10Hg�>��˜n�2��\w(u�[�tH����ͱ}M��D��w֬I�b `Z8�����0$�Z�2oϮ���8*Sc>��s^R�<U��.�O0�;�;���܈L�����;��[>��O{����,��Ex{ֆ�Nw}7I޹�;���[��yI`�oV�]os�`����=f5)l�avs�+I[��Z�ˌ4��+��C��b��Av�.rԶ���[(�iC3v���a=׏����ۓ�,蓤�8���R����銅1{�C@�	�T�1��8��ݧ�epI�*	>��6%�x�Lځ�<���yS�a��#;9��'8�ѕ0K����6�ir�[(�7d���Eo�VYΚ�n*Nd�m�NӠ�p^���t��P61eM��]���y�e$��<�$�cF񰻦S$^u�bƗ��c�59e֝����Ѷ('Y]NѢ��=+�o������ߚ�V�M����b`v��d��˫���*�T�f��q"+{aT���JJ���T�����y�kڭ�}J�<`�������kN�ӽ�BK���t����7)�꘠Ӽ���75kj�t�Y�����Ӊ�_V^e.YA�ìX��e�Y�M�i����J��L3c2�)���G�c�N��$b�BT�.�P}:v�z�����Gw:����׈v�h�um�-��)���r�N��mՁ\�:ᄭ*k{&32v:�*��ć2�\��ޘ�{�G˹-����Z��ZڟZ��krހ��NM����@�K�� 	nW'a�]���غ���^�3H���5��hpL��N��WM��Z60�܊襺1)���i�!]��pwwn��)@��T���Hg1x.�V�v�qt�������3W/|HK.�˻�e�0�J��c��b�Z����F�f�y����E[`tx�5ȶ�]�r�+��Ý���iY���_Mj�t��� �w[�5|�5Ԫn�HӠ��EN�Vb��F�t���.�һb_H��vc�R�Vq<&�HoÙ��!aÂPc�Uս��aC(��q�َ9n�e��O(���Zic�4�1
N--� F�b�����݋���9�]�zv�M�*��n�V��Yk������ӜҮ@×:�\cDq�����*�b���
數�2�і�ums�#��E���ǁl�=��8�4p(�9j�6�8��
J�$���D�A���S����Zp-}�(^r�ԫ�hŴ���FA��{0PW���tTVI9��E��+�B30���B2^k�u=颵��U��d�qV�P)�0z�)�׽�w�����~S�<��BZ��|V�����o�6�V���ؚ���q�n�J�j�ա][���������.7.�\�Ca�Y@㾔B���M��{;0c���RZ\0�3K,g i+�+�#+F��75`5M��y��C�gdڕi^��ͩ���|���)�듌��=���m�ߠ��n�e�]l\voa�(�rL8��^<�Hdl�v��{����[}�����Q]0�Ƹ�3f����Q,�|x��o�MDmEk���C���1���ȟr�vv����F�.���hu��ҏA�C�W:�ڽ���q7�5�9ؗf���b�j���vGO�]vpU;S�:�2��Y����rG�;�˹��^�|���e�UԱWe�^3)Q�J��m�^�6u���i	���:M�P�'d���	����%;'��:Ƒ'ru�v�²���.�f�7�q�]���YC��أ}�)�ϣ8K�tg:u�$ø;[�(�&KF�qY.�"��b���ʄ���QoR�98α�Sf���}gVd��LV��ę�4�I�/���#�����fo�^�N��R/����Е��.Ep�F�wOnM�1EG�:j"��;������w�L�� H�o���ZlR�L�'�s߳8L�s�����l���r���rS2������F��ԓ4rh��kpɻ�6�W�����:c���幉�mx�n����Ee6e��n��IU�(�;��,x���L=�v!J��.]�2#��s�:�����Z<G�+�OT
�H�6���<�v������v�6��]yz+���ݑ>zB;�Cόm&���b��i{���zU��x����[WJ<͂����j�[�["*�Cp%.u����+8~�����
��sv��R����XVѨ��U,����41Y�F:�I�/Ws��u���Ӎf�Q��uq{�4�L}��X�h��Oz���	��c*ɻ0)2�
k&fC�3,�jɺ0A����{��JaZ��j��k<�Q#�[���c�U�Vͣ�us�|��ҏ>����9���R��VD<ș��ǒ8]�!���,�`̢��چk���J�H��/���H���B�5�*�r�̰��/{��������>��b�'�*U�#���yHwC�q�ՠȁr�S�"2�tt�Cu��81G�i�Vo�	X��qm�[�L�}�Yop��j�Y��T[n���0�� �ú�
�>��6q�Ҽ���{�`��K}�G7k-u1Q�pN��z���?5]�X�z�r��9��F�T!�@ÂȔ�\1u� �.k�K��Y1Ԡ��Gf�ud���OV�$��z��X�s�%��-"��R�#�k����7L�b)�{�4uص��*$��5̲e����W�E{���PO+��
���`�NzR����v%d�6ޛ��nd�)ֱ)����g�1�%��i]����c�pA�<�}(=v�8L'�镪��ڒuMk�*�:�F�̻�sox�����}Z$b�yӸbT�l�)u*��� �r3h��b����`.�n��p<�����N��u�#��Ԇֺ��놐`�ٗ�2�;8�$ӾI��/�^Wַs�Ks6���f��j,��4skpB������u!I��:����_!�8Y�kkf�p��]��VM�ʹh14l2�-.�A0�;��xY#�ҝ�񵘊��M�:I��l�LFh��W[6.`_r�md��|��t����xoj��l��hm��]��LX�e�|�.#�
�+)��ܴң��hA:�F���p`6��(�t"����*�]���ы���T;F;�.��=�	J��R[�Ӎ��D���Xwy�QQ�8I[i팻Z�(V�+彧;��HţEq�/���͌��;�[^�Z�T�N���Q@vp���,���|�'����4�V�a2�`����&��	I�KN@!ܘ��hθ��d��JZ�0K�F�;Wg�1�j#}}yN��@W:㼨�9�	�T�����$-�o{��[F�E.�T��Y0^���Y����g�N���?=�C��r�!Y�"N�Dr�����Cy����26��r��7/����V���.��'AE\+6F�f��-�� �ܵ�N�8�uݗ;�$/M�[��he*i�8��!�m�e
zws��Ӗ��-��z�E�PVEBLx��	�rN��}ұ�����ƚ�f�������J��/�U�E"s��=Ee���X��%����QSwF�47�(�A�k�]�����9c|y��q�y��LKDW�a�E�a�����wV�
O��ֽ�[CF�bͤ+oz���Ќ�g,�k:�rfi ���Bh�٢�8r���2��k�W����i���c컾�)�%�18�"æ��iM!�:dVL�����	kO�ǻ��wjuU�������d�I�A�f5ݏ��]P)�YÝ:�7���5��n�	��}���)vE�����i���sWQ�x*׷�#�J��kgeX�E���%�	<��疰8��_GP�
Yz�U��r�M[(�me�Zܗu�q��)V�Nr�ɡl�yȀ��i��wѬt��:�\�qԙ(ɻyV�Gk-!\�=�_f��r��Y�>}|-����i�\h�ps<�x0s}�����NW{����N��U&]ĝb���y�yƦ� �.�j=�yM;�K�1�2��1_M�fɼ�}J`���۬p�7��dy��#���K5���õ�|3���R{�2K�t�ki��G�s3���t9U�!s�n��Fve�n�<R��ݽ\B���N���\�]r#��{�n�Z쬔���Y����&#VV�`ytH�kcڽy�&�r��T_f_ti�*5����UNU�]
��.�S6�R�K��_]f�.E�u�o]st]�<��R�_VWbJ��V]t�}s�]�w�mN�bԋ�=[���4�.����$7ݬ�͔���z���	�E��7MSDܬ���S����fZ.�(j��/��-tFs��iE�_gu>G�⛓r|��sK�6:�Ab��;�Y�K������'jơͮ����ҋa�˕��)>jT2ڂ�Vu���CM�º8�޹��:��P�u�w��v(A�t"2%�)�;k8����gה�d���>�$I楣��t�6�f:��T+{�K��V����V�v�4���Ϻ&�K�j�y1�Eg,�Z!˱y��=0n�%qϽh$
����)��=�Grr�=M'z Y,EleknR��D"�h�RPY;�xZN���O����v�*XF��Z�lb��pc[��W��6�:���wyrg�<]ʶV���;�\���RRi�o3�R���xR�]�e�U8�A�D/!cy�]���9��\� ���䣮ݜ�nmG`SQ��wǐAg~ϖ��$�S��<ܺ����!���W�]"xx��y;zK�׃+����� .;�s���lf��]�Pd��=\S]�i�3�����u`��A2Q혰=�.��Μ�¥fި��S�+2�̓�;�6��<�"�=�xE�HX{��C^:��r*���v/�s-hf��⵬�ʊ�L�k��2���ڥ�f+Q�u�B�%���i��Z��W�Y�NS�F�ca�=����Q}E��J�
[�_��o��\LoJxۗ47Q6x��[��2�������0�t��|Υ�n����{*ء���;+�t�g�����+][�]�y�/�LX�C@�Jr�\f��79|2��`t���)x���o��жe�sEe%��X\��6QG\Ѯ�]��Z8���t���4��c]t�J]��H�:��Wf�^sqP,��[%l�U}�����f�pC׍�S{0�v�E[q�4�aJl��h��8��J�5~��u�K)"W\�)؛���ok|���X�sY�/��qX"���؆Zo��Jǽ���se�����볒�VifU�Hړ�^'�8��&se�S�)���kW����˕I�b9��u��ԅ�n��צ�K�tҨ��H�ji���h_G����D�ڥ;�d��V�8pWIVYT�=I���)n���ō����Ȇv]
t	ξ���9ƷEM��EZ�t��*l7� 6���s��ӷqq
���<�t��3
��S*.�AN��+!ٕ���3{����/f�b.�sx2�Yl�[��NL��)��Û�S�,�Uظf��m+��΍?-8Q�ژ�v�T,���!|�E%�r4���.�c9��mA}��p{M�]aC����T�[ٌ�b����7�m�;+s18��X� (�)�V��ClX�v�x��i�1�L�Zh��sA���Ka[�j��+���\�".���8��OpgYܰY�}鷼�%�5�I�'Ru�U�{��}�J��oG˷5�^�SB���!F�Tu�2Ơ�.�,Ts��`�Lc�.l��뮜]݀�q����X�K�6��S�ɘ����ޒɮ��<��g��F"�ý�כ��.�o0'P;Mf��٧�i�DTA���t�^Z�Pm����ps���nA���f	
'b��V�8`��ެ��9wc�>Xb����'��c��̖���Xۘ�繛���)��AG �9c����7�T�b�r��zͥ{|�F��"����;J٘%97)��n�c3`��4�ΨdWo��9�7|C��Z�o�EY�ǹ�Y�/\�avi=V�{���R�fTZHIuDu�/
��N��[��n����4��7��Ⱎ-ɀͦ�cO��N�͠�L���lraTV�{-&�,u�@vV}�t� Z��8JX�AI�� ���Μ���rza\�g<��XY��J`\gd7*��gP���_qrīׄ9[��n!��61j-U�����
���R�:ݵք�w:Cݬ�,�˳�5�;��ᨔ���R���m�Ϙ���}R݉5�켰-P:.ي��A�;�Yk�`w����8v��'	)*�LG�r���ᨹ[s�s���:����	]76�o6.��wQ��إ�4kpJ"].�y.g �E}�h���
���T�=mkK�g���W��P���=B��
:�$��jj���8 ��v�5��V�.cqN,���#���#�G5f�Sq�1k�q�.WBwE�w܌:�ʕ:�>��<`���ξZ.-I�����q�[�y���>X3���K�?n�k؞1�,~����@���CG�\��
�]N�.Z��D�ghtJX޽��n���kR��ogZ\/�+�-��AN������/(	����$fV����q�+TQbZ�X-���2�Á:�k�me�!��4%�5ml}�����2���j��s����Nգ�H�v��m�RˁUA��I)kӛU�ol\�0W�����u���	2�G��c�V	Ñ��7y�P���rO�vPB�j��+�P��[�'���p�w�]��&P�{w�VR�����B`[�-bh�b
��ǌ�5�S��� �(����	!!!����� ��! Cl OP�!���3�`@���	����H�2@�X6�6�I8� 0��I'XBq$Y$0����@!X�!$���:�u��Yl��m$'C�M�N2Cܰ�4���`b&$�Y$��!P�5BI�	�$+x�!�����0'��Hi �Y!�$��$HM O!=I'�'M��@�2�*�T�3T�6�q��`�=IԂ��I�&�HOPI�$�	�@�a��I��$'P�$'T�hi��	a:�4���$�BO;B	���'|�
BC�$�T�I�HH���:��M!6����hE�i�8���M�:�����!�BbCI
�Ba�$'��i�R��K�a+$�`ɻd�OPY$�� �N���`q x�I�	�XO{HO<�C�
2d�'�XI�=݇Y$:�*]P��`)P�I'�a�X�'l�m 8²���<I�C�H;�Xu�.��`�	*Hi%HB��u��Bb ���N��ݒV����0�Cyd�\�hE�@���1�C�	�u!��x��Τ�!�<d%��4�1
�l�^P���"���Y	�N%`q�{� )�5�1�CL�<d�P&���b��,&�d#i"�4ԄY��&�m`LH�I�l�bCibx�&�� ��4��$�@��i��!�CH����"�:Τ3����(���a�=N2gRcx�OXx�i!�:��C��Rݬ���x°4ɦ���,��P��i"�bm&�Bi	ԓ��Ć��Rx�8�����VHu'R�u&�`{j��V%�'P�-�6�!�C<d*��@�!�a �Y(������SL�)�ԁ��.������V"�����d�3,6ɾ�޲I�V�8�>3��5�(a6�f�T�1�E&ް�x��x�VM2W����0�@둆��Jx�;a�Ci<q��$�rśA9g�=���LC���/�Om6��&�i�����'RWl�'B,_S���8�|�g����r�|��Ɏ&�q���{�s�puF��O.�)���\N��q�-d�O�DnC5���ƪ��XKL�Dx���7�!�l4ŇR���ġԞ��{Mr��峭na�+\q��'�MS8�4G��.>!�dX�l�M9�Y��4��_U�l+�E�����X5͒�	�_,�����D3�Z~��>V�&v&��|J�P�[q1�^{}f�|k:��97,&.��"L�<������2
���b�˗�Ο��U��1��D7��]庠 �R(4�խt�5��	����H���:l�1)9���~.�p.�cB��K�C-��7 �C��8���y��+d--���[�1�z㻩)�D�� �A�f����8R�:ty��]�#��M�����0��9>.m�]��U��U�Pf`��v]f�An�q4����/{��x!��dw��e�]��H��w�d%W��҄q@¬��=���n���az����$է�����5 )�p��T	�zUF����]=���K�jC��s3%fZ��0��rŴ�X�aЏJ)�p��ha���<�� �¤;���f��18��ǣo�+�ъY�
�		�-_2�R}|s$������`#*\"���0�wU��]��t��a�_lago
����B
h�ܟkᕫ�bb���g��V����g13���;|!$X�v�o��E�w�iq�2)B�m�5�^+17��
�u���t�r�W,LW*V�c��ۆ�
���fT�}pB:�g�"��2��.�#4�=Y%:�NM�qm�.��݇IZX�Tux�cȳkK���ς*ZkU�LZu>��f�j|X"X��e��*Qi �`$+��퇑Q!��=*Ǩ2x벲	���W#��C0����=S��h�+�ǒv���)e"g����l�r��U�3n�^��\���	-k�u|�{�}����iv�:㵺z��K�V3�ػFtH�o��v�WFTŶM���β�����)8%��{�S\�#�eN�5b�7���b�v宒�n�[�����h�u����)#3s��{WJsgNE5L�XWz��|�&����%��f��h�4�F�V+��u��^�k"#��:��@\���"�ArS�/���(,��t�1ޘNU��r�v�jˮ�	�kȜ���L'Yׄ��v��N�Y�QY�@�x�k!��%B�J����Z���'1�h|�M���z�m����ۣ~�X֐�����md�#�3KI������q����+�gƦfTVq�V��������
'j�J*u�n�t�E�n!a���e��:qÆ��b�h�-K��!U����=�3��ړ���Q;�y���[����0�A˩�S$�:��twq�6��u�>ԩ��)K)y+>7i@L]{����@97{Zϣ��O:M�ôn����Wn������v��4gˌ�+2Ò�ڏ�̔���A�������P���;����T�/��E��B�&�3%r)�:��̫�TZ����ly��\0��7�Q�%����F�p���d��.Y[S%;F��$���a� kb��v����q��1Wt��'G+,@2QA��L>��*�Ӥ��E�}Њ�J�o���zB��w����R|�ٝ]Fh3+��ALHB��4�j�m$�I���&0�>�J��  ��s���I�i1$&0���.��@��@$	�i�OXi$+	<ݐ�@��� �$�H_:�&$8��'�IB<{�w!	�~�{�~���y��y��\޽���E���
�E(*���(>J�VT�"�DYm9����$f�EQbE&0��QAQ"1QTPAM%d�UZ�a�٤4,E�ZE�,1�`#_ZŊ(�Kb��QE��|otQ�ȌX�(DY�cQV(
�b"2,�k�h�GZ��cDX���LH�(�("��!Z�X����b$PQc�řmQQ�(*���*	b1�e�TQb�<h�T�E��jQQF0UTf4bֈEE��d�	�l�1Ԫ���(��*"�A"e�E�q�1)���S3�4�5E��`�	|�DQb:iE��1A��Ee=�(���"��U��H��Tt��A ��X%�c���G�*�bL޸�5X!p#�H�X�*�b"1ED�����+\�Eg��PЊ���wo֊*��b�Ɗ�DE�/�U��DE���TPT��QU���~͌�P�P�Q�±AA<���C�i0b�V��I*�X�Em�g�oA�Z�U(�iDTHŌLj�E]Ҩ�}ϳH���w(�Q}lETi�cUA߳^Z��G�F
*��b�eX""}j���a������԰G�Q���
�%g2���v\j�URV�KlQQb�b@��N]$%ge<�&���w�>H�J�ADQF
9j�&�*gϛѱQX(��vγH�H��b"(�{�4A���Z
"����Т",X�/�c�2�,��QV"��+�TD�Y��s��EhUP2��"���L��Qժ�J��l�S)�(������*0`�V�QS���6��{e`�"¤�����TQ)����2�`�`�+")i�w�lcm
m*�*�ϙU��0�$�GK�ՁM5�������5�|�رAc�PA��b�X��*"�=ɦ.�D��MP*���b�6��<k�V/<��XV�)YE�AH�&��R,]}洜j�{�1�����(|�A3܅a������,��8�-���6��N5��EC�ϴ8kU�3 �X[*�����|�#���E6�?4+��4��.�EDDc1���h�����=b���yْ�|� a�B���|�*�E���1E�k�J��Q���[PGo��X�{j(g��j�5AY��`|��ѿ0�SV��l����i����O�&,UJ����VW�jdQuh�X�ʞ?jPc��o\
n�F"�������>�2*��ʪ�5��`���f_�ʩ�)���7zee	ꈼwyز{6h��$�Ҫ*(�m�F�XJ&��4�X��ĹeS���&��U��R�Os�X���R��yh}�kS�^��e��wqLg�QS�3w�&Fcb_���|C��nƔM�E���v�D����B�¢�M��j���R҃�b��&Z����Fq� � 
�GV!-wq�N��e��띞{�=�X�yhn��UW�ӧEE����3�Q��h��Ȫ��*�heR��N�X��B����̘�f?:��"�e��w��
"�9���<�A��
�/�\7i�f/�6�ǶV���������)DD�b9j��,ӥ�QO�ϩ��K��lu���'$J�=�}kk7w�	 ��~*#�R+�t�o�ǔ���#E��z�"}���,�H����w�5�0�ԛLU�y1�8`(]a�i_Y]'�sVS(�PU��` ��}��q1VU-=������~��+��5q�Qwi~}t�:��׍F"#�
��!*�����GufV�V��k�����{����Q<�ܦ+-����6�#��۠T���<�9�u�!TE�~n
/��c�>�K���TEkb0ݍ�J�thD�>ʪ�j���5�nE8yj ��s������f5���_|�E��DY�)  ��zs}��w�_��V+��Wnn_:�N�!eSy��0��{IV!kݕ�8ش%5�N�+&�%���x��NhN٢ � ݻ��e;r����H+̭�!��=�@h�;�@������e���i��o*97h/k�{��8F^�%�ݪ�D�Y�p�-�<��EY�Q1,Ew[����(Z�����UQĨ���]f��Q+�g;�=x,~�/�����7�����DOmue��LJ����a�h��x8��q��T�o^�:x��!A'�!-�;���]�˧u��_���_��h�B��U[x⹼�3i.�,U}�v]�R�R�k��*8����'���9�7��Ӕ��s\�Wn�]ATr���(��\�PG.e\�r�ܘyC�1ժV�u��Zd����(��~<� ���<b��{(�xWܮI[x;�y�3* ���#��=�>5;kcmN��ݸ�ՔǸS���8��3=�Euh��g=�lUE���b��q�5r�i��������MKM8��g��o�Q[�[.Sv���_7#4�̢H.�PK�dq��-V/X�����S����=����:�Y�q�u�o`�Y̪2��ѽ���Y,AQ��[�؆�k)ֱ�3�f:*j�
��%w|��(�ݾ\5�wh�D���7���}K����"�l��-�	�D�H#�pmֱ�]I�3}|�g�^UJ��I�ىX�B�1���m���y����G>ɤD5j}�a�s�w
�ED��_s��s)fZ��s|ѳ_\Oh`�n�8�J/���k&m��rf����)QB�`����"�@�~?8���R�<��\^�Ffd�ЫwV�i`����(K��BHճ��*-�0U��'|ю���5�����M���%h�������g���_���r�������eyj�˷b�)q�K�WWYS��<j(�왫(��a��w��ܥ��[;��l]�wk����+�_��%L���4����Lm�TK/��j��f�i*�|��}�<h�YiQ۞��t�[�W�UPr�{LbkV�Tr�⮯�w�&�r�V��E�-Dc�W���mE�Y1 ��{U�*]�*���Ʌ�ӊ|��4�&�����_8�EhH>K���Y673��y�����s.>�����h���Um
�o���I�m��J2����{Ӌ���
�����{�m/Zk�昭��)�V6��;w�5�4pBEnS�q
�F�e�m&����$�ǐD�|��3�6�T"���i�ev��h�ۖ��n�:�c`� yu�=����H����*�?�ܨ��of�b���3"������ԬX�P�[��߷��f(�4S5��߂�����}���W�1���լUo��MFw/uT��6�Llj�>�G]����&bUD�s�T�~jꢈֱOoΝ'���٬M��ѡ�*���B��Y�^��Ϲ�h�����q@���Y�����*�\�c&�cUk{eb}�~Gz������.�]��Ӿ��R����r��d�4�����Nd:+�qE�� ��m.������gtx2Ɗr�c+���Q98� E��Wk]9�v�%n��"3H�{>��(�#'�fR��;���^HG$p������	 EM�z����-j��u�U�x�'�l�T�s3&\�Ҙ[�]4�cl��}�|�T~̘���Gt�WI`�[��I���jh��H	�]�f�#�7y�j8&�}���(
��/��T�<O)Ε�"����k�Q}�������ye���\D?(�i.a�Ծd^x�_M�tSn1qƭn��hpb#�7#�2~���"|�-au�at�Хl���r<��5����~��_S__����v�-��A��7`y�ڠ���ٱ<�KKZ>��n�ט\�$�!\���$Y�̂�B�G�z��@EE�Y�7}���� ��!&�{�#�k���c�1�sM��V�)ysyy��kx�L�<�͋�I���|keSJ�3���`#�p��w�O�����.Df4[co=���S߷n��Z&٥:����4(�9g��0u/]ˣ�f��A����`�R�*ք$^e� �O �~�^Q�=k��MBs|<4� ��?$���*�*^'��$�v�����1��w�v�yL�-?ZJz��/2�$h��@@Ý�(bD�$���k}�D��@�"�H�c\t�g�$��5u���m$8���UK6M�'ZMoW�s��6�t��+LV)~��Pg��b�3-[]�Gϯ=ru$/>�`�O�{��U�W�_���,-;&r�����6	�e�P?[� ���[�pO�?(h�i�P�U  �x�Q �i������|�U�&�H��]nV化�����.K���B?"�/�&�$n֩f�����W�7��]2��jN]L�u=��4h
�a����Qwm��<����p�q��p���ն^*�Oz,X1��$���7M�cg��F�%/���F�+��y�3����v����A�s7,>���C�!���*w&��*�XVI��v������hڝ�������B{VKz>��R�!|��˺"�
(���Po��vg��)����b��e�h�w��柛�s6�i�a�4$�E�|��ܰ��Mx�M��S�����)��`�v�#j,��|�|L�n���7�/�>���z��)X���rVT�gR]7���M][��c������]�g$��V���+�ٺmj�z:�1�.�̺콽�	�#k��K�i���r��+}+�07&��=�Lɶ_����qQ��$l��6���3�kMb��aZ���{�{I�#Kq����@P!��P���G<���uH�(��'R?�Q=G��9����� �ul���eݐ�|�k�ppJʵ�K2��c��"�O�v�(��>:b�7�6n�Z��6�+��8�!?�toj��|�Hk�t�1q����� |GX#�=4P�J�K�	�827噲�W�z����\��C�h��`�ֈ�SG�J�7#���h�J+:8RD7pA�(!�����@�i��ۛ3ʐ����r$@ �M�?|�G�c���~���D^����(���������XȘ$�p�>$���[$�$x��z�}�n: �f�9�/4!l������>/�	���ֵ1�@�N�=;58�=��I��^�yW��6�/j��tq-�$(��úv�cѰHD�^&qg����H!$�L�����m�]Pd�!�}�B�+���4~���>y����+�;�'���@	+'�\��$�U�};�"u��en8	� u뀌:��������=B6~d�vH���������n��Q_"�7�v��[C�&
|5�7Q������� �ʊ�̥)��7,{+;� �D�d�D|���G�
"����&�y/ta��lA#z��y���gnǔ��Y����$�N7�@�R�����
�0��^A6�Dc�]A��L��=�b �!�FܷV���&�EmmQ;�kJv��!7�m��(v��1�׸5��Y�����8q<i���>�z��)L��"I �]>	�0�YF�'y/�c�_tL��u������J�@�T���A|G�~٧��֎Z+�k�u��gs�����j=M��C۽'+��$a��.���Ue!�a��y�}�^��4�&�a|e�� �B��ˎ1�|�Wg�8��&n̬Yg�:�P��2E�V�%�y:��r�W!9:R�͙ۣ�Ѫ�����%�����+�akɧ�
��M.��M]�]�η��/������f�e��x�V�f'Lƨbu����0�t2mG����Z�&p̮M)�$V=���4&�p������������R�	��&��@H����h6�rAy񦐍��oyō��%U;�^h������B�@�����?���y��ƍ��%__���A�Z$Z��� A�뗦��R��J(ZCg�Wf�ZE��Dzx��$���`��c��!ίxa��z�	jd��Xj��?x���=�ȹP���Q�O�55��U��  ��F��GG�E�����'�0AB�_D�^.8U*@�'�C@R������
�ޅ�i�F�h��Lu�ZK�۫�V=ꃅd�s����9CHjc�g���u�b�B7��`����W����@�^&���h��:�6�5A��@���o�E>_��E\L���&�$���[�11�_�?SJ�sk2>Y�u��J+u�L?���M�� ��QCb鴑�W��
3$^�jz�(Oȯ��1�h2�˖6O��C�!�a�˾�WQ�ur����s�����T��*^G�c��:g��D��)W;gG�K���������<�!�P䃹��*������k֐�]7�m��C�W��Y緾z.�mpփc��@��M6��8�,�����-2*�Qҳ���
'�~e��@�ߔ�u�4!��t���i�z#�I|� gk�K����FF�x��:..��*�:�2�J�c�󸎨�$~d���x�6C(���vs�$�90!24�$#K�]��a��z���x�M�b�X%([8��"ս�u����%�)n���?2�Ae ���y���(���K�T�֛"s	��?|t��k���T�D��t6ރ��V��r;/Mx/�y��Z�$rdq�|H&���=]�#����{�eftW5�ˑꌜ�c��I#(R@��+�H{yueY ���`�W��)aDE����JƩs����Qu͐��!j��ô��e������8"�@�O}�>�'s�����!�f@�m}du '���h�|�<$��'�����+�>��l�冼��}��_���6\���ͦ`۫�' �%t���o;�l01qW�X�r��b�Y����?}�6��X���f�n߯J�n�N�n�7�g!)�o+'B�K�-��	]�W�ʑn6�	�<=\Ov j$�E��c�w˝(��������Tx�]Z�4�T�u3�置	�i���ϱ���!c��G*�P�~Bٙ�f�5�m����>�e8����h�	y%��������	
��C<�Q
�x�"����2h��Y������Q��j�H𦇞*�i�*�o�4��Q��l������Y��b�3�m�˲�_gd-W� ?�ؾ�}�)�)�ΰ����h.Y�x Z�U���@�׽3b�YU�/��������X�^�}؂���ܷ��0��UU������$$��u1�{!�랈�:�1�|��S2��E4I�ť48���"�6�IZl���^2�'�]0���-��0������O����YV)�e��C�� �������yڌ�t�۾���0�+AH���y�+�Y��_!�Me���X�G�ka/�6�v�j�C�	���oˇ�K��]�U���/A�(Q����jT4B+Ŋ^�a݁��R3�T I��V1�j����u��d4�"�^'�#%�R��	����m��ĕn����^��ü��y�X ���LSa�h�)�izFx��g�����<z��d^nc&�*4�7�g�͉͐�͎�>���k�vf�w���f�����b�J�S%
�Q|��A�E�a��"�
>:����$�<$pS��e4�U��@���"61�U�
��/�B��'s�$�)f���
^'G7����	z�4����F�!"��?Y]�3h�
�uϩxch}@t���ٟD#���"au������Ɍ��;��z.n��x��A��H̗Vg�AMvs���#	�-k��Txh.{�^�� `�l��-у7�Q�Q��_�o�ڀVP�V�y���W�\&��a���33JK)�c5���`a8U� �30lC3yu�_����w ���7����'2�{w���9��n�Y_���;�̜>�eL��=�{�}������,�Vw��<�\c�����澍�R���{.}��=r��]���p.�y3E;M)����kPm倊�n�ie9��E�zU����=w�Cz$���~���>�"���'��9!q���Ӳ|A��"K(_Te/D�=Vi�$T���k�5�C�`�yF;���F1���!�C3A��4���Z���V%A�C)��0A_.`�/�q}���Z-A�DG�!�1F��1{vlPK �uP3Ct�"�(����Z*���B�O{|��E���i��1�B!�h�BE�	�-�! �o��$ʧ�=pΎ:=]�.!~As�=�$6�h�(��󔆁�P�T�;v*������Z�,p=�qQ|���S�(5F�W�D&�zz1��
�dR�L�I�g@�rP8����� Yf�j%�OJ�Ck�O����.�׎�~|�wc��Vv�����,5H¶|yC9i���J=�<[^�M�i|R���Qv�W�Ȑߤ��c�_k��W
s�G�'������T{�y�����F��#�x���,n1Z��]	�o�iwc��]��Ǻ8��N �N>u��E	6��@��Z����������x�o<�P�+�N+�Pa���dn|����\<��[T`�t��54�� G��T�p�=r<͇���$�j��`�ԑ>��S;��8�;cs<hgVZ��1g�)���n��(���];�0�l�{���j�=���u�F�yF�3uz!v�2n�8��7���* �_p������<ػ��ww�g4 ���(�Mb��g�9�H���FN��z/�$XE��o��9������[�jɃ	����>�������`4ӱ����Ou�2�dÝ���V
N���8E�r\s*$���p,Y@񻃥�񀢏��L�*�O����0x�Ly�m*۹T? �X,I>!�����T��1�S�g��W�;=��5{,L���Uι� �.늞;Ø4B�ÿ����D;'���>������K�w��n�J�ơ�Wݳ5evu�&�>�{�״�,���l�X���,�sUsn���v�y����!^��td�[:r�~Y)E5�M�d���6��Go>*^Ca���{�k� �h��w���V�a4���UDA:������K��t	ІG���,(��x��^8Z9�!�A5m5pqJ��f��mۯ��U/zT>�2�K�Q͎<� ?<��|�%� 3:*���U=�T���]�yf�:"�qQS�W3K陦��u]��um̓�V��X~��8�\�"~c����o��/��9�M��>����6�Y�{����Wۺb��V�iE�]�P����i��IY�={��_=}�!�j�|z���P�Q��gD�A#ͳp�&�erO�cT!?2� �+�<�6�І4J
�iX��V
������/�
��XA�"H<�M(�DR~%��E�Ls��d�|���Wj�">L��Q���
��d�UX�����Ѷ�g�z��gZ��Y�e�^�g����I���@%�� �|,�h�ax����C�廷���)j��]\�.��ǎ#X��nE�l�Z)M�.���A>����}-���b�C-
�ݲ���s�g='C{䘢�r/��c�w"`��׃�I*k`�Ǔ��� 0^�7�?:��U5[��R�yPU���V��c�x�����*��f����;�<s�_�N4l� %r�'�EX>�b�qc� )+q8�3*h����-W��Ĝ���i�PV�T=Xqta�!����G3M ��Q�k4��"���v9P �b\��aZ\Mx����UFM*����/)q���휜���ǋ����!�������0�)$o���Q/$AgQ(2�4��l��Y����'�����d�`�e�#\�,ZM@a���y����nAuMS�J�����ʜ�o9?����B�6�����z9���Z�3�R�c��_)���1����(e�"�z�V�國��3��q�3qgB��ha��Z��WV�G����*�v�r�
���BJT2vuK�� �Uў�Z���j�XC]�g�`����:�r��H��"f��Eh ���+�-� ?��U�9d����@�d W�� �cg���31��-�5�se_��7ﮯ>�+��&�	U����6k���e�!�:u̕>恉i�WJ6�ڪD[{̎-Ք��re��t��ʯ ���t�<���L��WqN�;�;]�J��i�2E�����RP���D�#�MK�~�z_ݟC��h�B{��W�����"]Ueym�S[F�`
��������>j�|�X��>@����d1d�����J�Q�QB�>!aS[$>c\ C	����̚��˥���~�޲��$�( "��0| �����D��۰�)
!��G���	#H�Ğ����E����r��7<�S�z���8T������[c'��,8�א�c�F�z{�	*�2x��Ac�=�>(�^�o�y�M:?��X�ޔ�Z�t�|H�Z�r{�ش��Y�ۦ�f{�>!cD���Gz��,���O��t"�tׅ�Kɇ�iMe3���4a)�e�	3�!��;�B�Ix���-���y�t�օ
�ىb�kB"�| ������`V�@a�`��#�hl���y)^�����yiB	�@ri��B�4�/�Tq�y��ك��ͫ���w�D$o`@z&(ע������c�ˑW1Xj�/@hx���P�g[*�(*�J�E���������������n�z�����c�����C=�A�Q�����.n
!x�W��xVjS-}�o��R ����m�]~��i��V9�hA��6g��C&S��NtYQ����7gEb�\F�8�_pqu6�+x��{|���B+�
�v�}r��sˋ�h1Y�|�����e��{
6Ծ�:��s.3d|-�]0˭����A�5��;Cx������,�s�vc��
h�f�x~T��^�͓7�W��dOR5Z�%���0��8w�F�[Si�[��$K%J��?$��)���Mt�x���k�M�l�<��tB���	����s�T$�k��� ����I�q|��C*�%b�D���z���F5���Ѯ��?(͗#���W	x,k�Ɵ:*�D6�}�Y]�}�*�8���������Tp�W�g�2>&���o��y��l�kV������z[����l�L�8����=�_ �C��% EC�T��#��=-�~���L����#��ł^����0�q˃[�{&{֤^��F�yw�Q�5د�.�����R4�u�L'�6���K�-��z� �]�ƹ�x��A��6@A�M�sЃ�jz�x<��3Z���%jb읿{ y����s��=�A��/}�q��5��F ��%R����>p5��.����PW�uя�?�z�O\�����^ݚ|�ڮ�őǹ!��޳I4V?,��B�d$�O%�7��;��0���R����0���}ͺr��� T�h�$ЯSd��ۇ�3�w���K�}�t��TT�*/�QgL�Y,�:�wM����O/o]�4���|+O�U�6�8D>5����K��B��p�<���}R��u{^f�%��('�d��4B�(�μ�| O�h�S�F�H��R�����}\�i��t~�:	}��$j�㾿{�V[�u��m)��<��K�`�I��a���|*,�4�W
_����}�����C�A��8�)��C(��dS=�n�諭}nW=d?u�f1o���:���?�ms��۬�b�]IӨU�#��2�m������ �u���Z�̧���
�F�N�?�)jY�f�h�6�]��/G���t@��2�(��}�R|������S��䳑[��;���7R�d�Lh��3B�wE9�kiM�˨����u{$�btά��U��<�5���x.��M�ȥ�X�a��ic������nG��c�@�}���@WSA��^���j�<n�D�'�hP���
Rj�v"y����&��:RjvS޲����sj������YN��O5	+yqa��ŗ)Mm��|	4�d�W�݂Ӯ����#}su����:�W�N��%-��V�(n�D��/���'���j���%g7Vg�EZ32e�;�͢q���%�v�/s(͋5�N�V�Ӻ�P�o7kOq@�Vo<yR���a�]ʭ��s]����\2��u-v����S��'L1yu���o7( ]����!��(�@g�!Z֯��˘�vP�ו���7�g�twХWÊ`�*ʛ�D}���<q#N r�%�.�µ�.�ݭwl�+p��Rݓ��'{��3�j;����kX��B3-�)�7j���7������e=�3�����r�>��[ϴ,nv���/`�����΅�o/P�b�u3Ɵ6�:�i�ڝ�W|]�j\)qt�cΥN�8�icy�߭��E�4e��Sr ]Q�ʻ�=�J��)9e]���T��])���%���+��G����+�5�U�����ii䞔��b{��q5�N�(Kf>��A4@�un��W�A;��X��Cw�ȈYN�׳��wUKV箮���������̺PGj����Cm6��oe@:����V:����o\���s]�լ4;����1]	�<痐(��vz�{b�>w����}D,E��b34���ǈV�D4��SHW3/�\鵠s����ƛ̝��])�,8�;��$gsS`�[S�c`���R8�Ȼ�����X��~'�����V��:�w�偽EKJ����ĭA�� |rm.t͢�Z���Z�I�i��ʴ�-s紨C���A�*���������3��"�w�y�:{W��{";���⑛6Q���e5�2��U��=��B���_=B�J������0eN)7	r��.��pa���j�q�u�3-a�����9ݕ��[�P�\t��y�ˋ�/{�]@��i^lR�`��5�\u}:��.��W'z����<��q��'���Ծs:�v;o���AT�:��^]1����k��rK��<�SQ��*�]\��ȵ$�D�X0� �R27�*�h$��0�����������k�;UO.9&��������C���㢭���@��r���L�BMXq�+9s]�f}�]4��X�s{�vV�/\b7�s6�3W�?B	��H����B,��T�����i���Vi;�4����x����MZg��M'�Y��͝��u��bm)�����ԭw��]���ar�Ͻќ��.&�Fc??g<�lĝ�.�]��_}�vc�:��L�xa�����F���Z�4/T�{٭��o����c5��֞����=C?~��u:��N{|c�r�{��q�������^h�������Ϭ<y҈��11�g�4i4�� ��ퟝ��>�]O{f2�b&�w�<�̼�z�SL?;G�aș��rͻ�6��|g��x7\q��cC��9�����O�&����p��ϲ�f��.�|���q��E����Y��~C;f�_u�-��cP6��ރI�24�_}=NE�?2�T��O�:�L�I�t�_ɤ�ݳWW�t}C����{�'ƍ�����-)��u�{/}�^ە�ă��A?$�����i�3y����6�t�֩Is�֐�)�nr��?��~�k�1/�i��Tw&��q�u}�w�Kl=O]j��B��bm<�S��x�I�4G=���x�Lb˺T3�>���~���2�foH�m�h�
�(3LU~�F>��o_�s�+�L��0���o�P�oT+.�o�����e՚�bV�����I��igl{��g9�Ne����W����p��C��?����c�;�Z���t����y��i���R�?':��ۚE������o���\5������~��ϯ�ZmEL*u3����<��%`�7���S��O^�h�LO<��Ayq�6�˦�M��Χ��,�"���1x�H� d3�:C����Њ~v���éP��x��?h��/�f2������Èp�O5TL &�{ZG;���W�������k��G�M����e���Wm�S~kE*_��E�i�Y�J�j���2Ӊ�v��Hi3+���t�M'��g���z6�<��h�sF~�b3WxM&�e������~g�㧩���4�ve����L�L�,:��t���B��wo/�Κ������?x|��>������}[���/�c�c�G>=M'-Y���_y^�T�y�k�T�.���]����D�Qea����N&�v�).�Q�~��tm��I����6�5���1�J!����)�c:�:�Ɣ_�s���I*?*C���u��tv}�6��}��G��="��}�<���] �S�4�����C�8�&��'6i1/�Dƥu����}g8{���|�>��G�}OY�Ku�]7I��5�i5s4�'��먼O̺�����o��Sl���޿0Ћ��`�ߠ}�q>���v�-����{�w36��+��m��*g����s�x�!�Os9�`�䮙����'<�Z�g�sfى*m⪉����~��hT4����f5�M�����w�0�|� y~xȂ��?�V�z㬤ި���t�4����ح`�Ŀ1�^���Mwk��.��Ii&��}C%g8vW[�/t��]�	qu�1�c��ʡ҅�^㎺�_tjV7��2�6�����RL������8��}mqq=�1=���.j�y6�m�S��;��#Eԉ�ճU�ѝ����~C������K�K����T/}�6_�z�M+�^����w����+�/y�ٴDy�u�}�3�]��(bJ��bw�"�Hm��z�S�<���|��B�& �f&{K�힧3�
�:g��:O�uv�D��]�)[�"�	���#iǨa�C��Q*g�/��o]�0�]k��is�4�T*��8��ʇ+�0��'Pg(�%<���=y�/�f6-���^1M�|�>���Ϭ��߼)��ϼ��׻�Y��b�m&|��]�µ1����ܝ���K�7�����L��t�����5C�|���3ve��5��4��l8��no��*<���5G����~gEt�-�A�h�^P�j�����t%�O������@>[�� L}��ھ!�����Q���6�o����lg�߹]���4�M{���;���<Cv��|���
��B�yJ���:8�E�C�by����u�M0��q��<��+�vg)M�Z��2��_NDC���i�����~��Z��R��3��s�s@�Wղ���riy3�����җ��B�M$�7�\Iϩr�Xs�~�|�za�������9��>h�J�{��1�sx������͡�?q��������#�2?�[c��;��~k	;uy�z7ֿ�	� � O�_�c�:�[z�Y���םo'Fu�5�sT��0GT�2��M:fa���Ӛ��?&�o[�͛��S�T���,��}����,�k�{��Ew�Hb(�x��XgbiщEQf0���Jh��"@�/A�8	��u^�����'ω��S�)l6�8�z�5����iЋ1�����r�in;N'�ķ��y�׬�f��!ns[f�S�bO|��7��I~�fR��'�i��I�����yM�_ߨi�Q��@!�G� B��"
�Ԭ�&���~����w���ݦ�}���v�����4�.�L1�����5���6������Lɷ7J�a뉓�3o���h�7�5�SH�����a�M���l���1�m
��z��>�wL��fX��'�������`)o�tK�ٶ����o��cp�z�T��-��������}�Ì0�M����j��.�k���¾%�p�!��DY :X�o߈��"OB�
��5�p �
�Vp�'��ݢ�ٽ��#c��4��s�W�yQQh�fL���d��x�{<��5�Z�eY]���K�?[�
�R��:��k�_�[8��Z��:I�\)�Š�+��\v'���]a���z)�Y�:�dz��Zf��Dq�o����VeVn��1���a�K��&�^.�b�e
6���CgG�yWKc�SA�����(Y���Jz07c�g-�<')%	'�����n�f/'�Sg��i$B�%�C���y:c ��.��{�!��񩅴�����ta �����d���^W�F.�j�ך�����AZ��]��f�ز��_k��F��q3�����,��L�#���g�|��? �A^>�Kvy�c��p�����	��N����MX<y�ʒ�R�/��6;�)�҃��_25��{cҞ�t�@��ٟ)�ܨ߻�f�����U.(/I"CRE�
��_�<��{��|�\]����g����lDw���eu'M��뮒3�)�����eo���W�(���fthD�m�-JA�����ع�r��{ۗ��K��u@��X�$�ݽ��Z<�ry������Ӕ����D����h�`:=�.W���}LA�}	E	��#�_��!��7�3�բ�����s�,c��S6���Š+d���Q��>m����t7�t@`�� �6��HO�'8ڥIf��&�]-eH�կ~����$�p{B�f�_:RAۼ�.�z��v�
2-���^{:,F!�B��'/NC���xuQ��ׅR�����0z��,[�׌�]K��Wyx�^�~��^~/�N0!@��A\�v�\]�hB�'�]��6�a�(H���@�^�)ͷb�@�p����(p��۞��VeK癰��|Y���#U
��ѳ@H.��F����<� ��LiJߜ"O/+j�Q�t�u=�`*N$���Ro�%��B�͹�7�&s�����fei����K������@r�nN����n�q֎����ͳB���hV���[5]*�Q��=R�.{�����
|$�yS6(���R�
��--�M�p����{ٻ��2�@	Q�s}�)�}*{~s{*����ZqBǕAIщ{����_?z9l�d�7G]�;�\�5jO��P�����-��Zz��?���7opgk�%�{scc�$J8�k��P��������		"<gx�Id}=�����%*���W�����/��ױo�,�d���
?���<}�nd�,�G6�nx��Y��5��+��0.;`�)�*��}C7|�N�H��<���i?j,���i�5�T����yL���{	SŢ�*����^��<�*IH�D.��$�6�\�T���~�^,���_��.���K�C\�D��7ɣ��^4����Hil�	D�(���I�v��c��l���� ��֪�dY�y^5����ۚ��:��|�b���������D�<�>9�+�$`If�39ߎ?�'��r�i�.�+�#*����X�̶`��a��MWZ�*"o�b;�O�L�0!�N�%0�_e=��H�]{'�¹�4`9���{���W���g,��CG�s@j�>�Ѡj%=#�uc�TC��M(�����O���c�#J)C<P��S9��m�����U��f��`�������-�ӭ@�9\c�P��B�x��8��6�8B��UٵjyV+w-��ν&���B��rFQ�s��f�?{�V��[W�)��a�I����^�W�B���\��p���h����Gڶ^O�Hd)A<G�o��g9�̫�|���UxYc'D�G9 9|0gD�7�k4׎�n�rP�n!��!�W�g��� r�6��iKk�Îr�h'2��C�ȟ^u���t}>B�)6�o���ѼOd3`m�񐱋�Dm��Z���vpU��r�%j�s��M�j>:r8�L��t���8|!�S�+1�Lk��[�[/�ʦ�y�3P�
���QB-�U{�y��Mm�o 0fs~����3���Hqk�vW�޹�5�X^�óa���s�6;�� ��Q�����tb}���R��Q�'���᷷���tG����� ^ԯ�n� �GGyv]n|Rx��V��Z��y����dС�9�S���hq�ք+LD҅r0I8zy��H�s�?��C��Za�C�j�cUC;]�U�u��'�h
��E3��Rq�	��a�L��A��xs������;_'�բ�H�޺+�z<����{�^23E%\xS ���tP:*�<�)���R���oTx���R�Z��Oӌ���eok��8S�>24'a�ClY�����9� �(W��8�Ϲ�C-$i�C:!Wu�Jy��������N��|W<�,V�+�VB�(��y�]��]w��<�S�y\3�l�
ws��$�,p\U�������е=�����Kcs3}��~�҉x�>��g�z��������m�͹���H�r�ci�&�b��N%�\�b�e�_m]����<�O_�8�q��3��4 ��nwf��O�C�MP�B�9C��]�`*4�C������TDY�o���G�N>ŏ�޽�_�\��n�hv@�6>�&0��$Y�M�4��]���P*�:�")�^����_��@����g�=\4/oI�W,���a�u������Ŋ�ܔ�f��!AvC�-f�+�7��h�@�m#�P�j�v�w���@�|pp�E�>�2�90�4H���ܙn�j��o3$�Mj��/��*���wL�nb�	�����0l���"���t�/��{�Ք>��x���d%D�+�0���BIӋ�AB�xHV����O9�E5�]+ᏻiy�z�U�<3�P>�����{�'ǥ?{��s񶶓�t�둄���&��0�]�9�*"�1�kDw��Z�q�!��k+ק����OfS&$�\�Ϛ\�vJ�X�/�q�'ʹ灋���iZ�����t]f��`���d��uǯ�6�ķkn!DV����VXpz�Լ)������(J^�'���Aʚ
S��r�~9
���9<����N���IF} =I��!K��Q�_K51*肬�_1U-o�ds7{���*({)xf��тn�ϼ�!���N�/^�Iy}ȋ.4]u�P�H��RLq�8�)�����F	����ν6��䙡fŀ1�q(Ay�~nΒ�^�	u ��X�ٷ�&[_��f�~�Dj�|U�!%[,��-,�PN�ۙe �l���$�
�ԧ����{���w�x{��a��/z�?rlw*�lMi����
}�hkW�w���4B6E6l��c���x��W����h^����0�ˡ��<f@��F�T4w���-.%�k/�}�g�24��2i����>��.�/�9��wdQ]�b(o9��yˌuB� ӭ��*� <�H���>�����"�!���[�Y�Jn�\�\���-~����A8�+o5�dv*����%b�.���9GA�s4����ݍDw
���rӬ{z)�MA�,�[�p������Y�����e*F�ȡw�����Wm�:�=�X9o6���:�a��������Mq]f,NM{�J�vwf�sP��I[.�[�u��S�C=��]���c�Cjݻ�=�!;Z��ֵL�\�y\��a����v&�+�b�ae�6��?"[|�y���ۡ']��f�6N��b&�v$j^U�y�{FP�V�T���z�Y����:V��!���w��V�L��D��/FݸEq0|���󃡫�Es�v)	tu�e��ZR֯��s���^��{�'4椴�4M��(J��l��f�B��8�#a��� ��ec躓�j��իٞ�8%<�Os�Y|s�]�
א�����c�������x��}�,��ƨ+yB�,N�C̱���������𡹗
�g��%�ވbǱ�ʤ)v$�krKpMi���/�[��k�H����y�"U��0��F�Ǆ)k��#P �1��'ޒ�Eo!��v��T����;.�2�/1ĉԙ�
�;k�T�׶_ι1��vi�Mf���
���l��{���JuԓJk9���V齘AV�=�QO��O:oy�(f��M����I�]2�)���,s=B{��z��Y}�f����j�ödܞ�GEf�.^ϏkW�j�*���}����WO�����q���!�`��2or���s�����t�)��E'���IW{��xVK���< 噸��ҞO�"q�����5�0U� ^��*�;o3��9��Q��d�yS�����>n��6�=FN��Wn����hr��e ]��f������﫸Ɛ��Κf�^^ٔ�P*����T}���g-�����\�Nk�Ҟ/�7`,tFm�w��(a���_]�#��om��|���|)����Z�k��hB�W]����!�P��<�c�������-|���x�Vf���zr�w��ރV<��r�O���b�cr:�Ϥ�O�)���J"�/J��dz�.�peYK��:C�k���:=Jh�ˎ���G��`~F�<yӵ�}tpT4d����A^�B����i��/N�4�nȯ��B��Z�P���]ˑx�A����a-�"�M��2uBr_�^����g-<,�+����Bjk©��;`"�5�z]{r��ҹXz�b��QC�Z*��e][QDNbx���o�7�O}5;�9��^ٳ�0Ջ*�#��o��7��'Q�.j~A��a�^�������{����z-m/B��`H��̣��$��q��[�Fη��[�}�'�Y<��)ٍ#�-U�~q$;��)�)"73��� |m��h���ZyU� ���u��m���΁ţs.
��U��I�z_�Ԗ�}��9����V�z��~���n�䅔����\��X\��ݲ�_cH%eI�lu�_�l)�a��G��;'����㛄Y��H<\��Ʃ.�y�l�7ۃ�n�1�w�q�Ւ�q�}�Cɋ�S<��}~ͱ3�w��Y�-W"� H��x{�j�zB�Q��bFM������퐭�WJ�|cI5p)�:�OW�k6զ����[E�:�*�
�B�����q�M�mS�j�匹tJ�2���[(�!�sy�W�}��(5w5|�]i�]�Z�d�5r)uM<�n���w��n]r8^	��s��޼�O_wX���%��*w\.���:��#ٖ+ynE�ˣ��_Q�>Q�j/�F���x2�SG��w�N�4���Mu��ge�D��N�T��6��lWz.̽�����R��p���| �ZB���
MdY�ԧ��OiY*#�N���+G�l��z*���l��_#�P�Ng{��s�0��3ۦ!F�$����X��ϗ���t(X�>q���$��W��<[npys��Mf�Bz���ս�\�׈�݅ߠ4�� �tӁ:p�w��(�5���b}�U'>>�tbT������ӽ���yX;}]��Ӎ��R�f&���b�u��aK�:�p;���
A��깯#`��g�uH=����~���Juf5��l��7Y".��Ւa�+�'RìU��)J�g��k�vT���R�#F1�M��\�����Z�u,�Z�KG�n���]�y(}.��C�r��
���c�>JJ���t)W��û�����(���=ep�n<�F�ʋט��+��>ۍ��)<Ӱ$H��t���P F�=���N%���cލP<h�Yk2����@�-0Djh�"����#�O{o��0�Տ�=+^���Cro/�q������.�I�yn���,�p.H_�z�n�k��(�Mf�2Ԯ=Xo��p;�؉Z72�<W���U����C�"u�{��	V��HYx��:���n>�������Z����%D�բh[Y�fg-ŭ_\�Ur�*ތU�+�X��2k��Y�%s�5��G���Y�ƺ�\��H�9��垢u�_��[O��6/�rA�q7���
�,��F2-��)����.�ڷ^����ѐ֝� �k=؊U��W�'���F�Hxo�z��.�SEV���Y����4v�t�@.yz��j�o��9	}Ҷ\:]��K:L�Bǋs�2<�A	ӛϴ��y�黑�w(Rw������Uf�����,�İ����i�>8
�I�¼N�-Մ}7X&��wz�'t.;�ۊ�҄Km�*'#���z*� ^$=�6�Y�H���~���;�R�^b��Yg;��x��z�:ܼ��b�V���gԱ�S�sn�?j#.��{��&QzF����o�5��'�ޒ�^{Ń�:(������4y8}�u*�e�C��cw���d�B=���^Nuh�J!m	�<� ��Dd~��)�=s�¦:�u�㓺��=�݋�W�{y���<��5��=C����>���z]��.f���&i����t-�y>�feB�W���(5�Q��F�`�9���\@��2n��gbKH���~���{��[w;���MC��$��Ҫ�
�?aO9��Ӷ�A�u���4���љ��5sX+3qm3��B.IxV��Mr/n�Jͫ�8�Rk�ut������T޷ue�mp��A�N֜�U�^u���vq(R�)���Ζd�3#�*��]D���4T�Ķ��l�x}�wF�]��C90o4grev�g	ܕ�/�yV�����AGE��W���Ǣ�֧wv���49hp���+�(���R$��q��.K��/��Ϋ
����ɫ\ҝ�f�GB[SL�s�ueUL8�D��y�E�b�I\��Un˹�c��eЎ�Q����w��3�I���Fɵ�SCX��՚CjP���	�Hg=�9>���t����g$b�[���0ٓ/K��B
��Z����_Q*fK2��W�
WK�m�I8���︔3S������ų%���&�d�d�8vg�(&Z� �Z$�֥А��z��5i��	"�����aN��|(W[���wOw�8-��5�
�f�E^�:$j ���.������t��t���]܆Mi�J�+a|��F%���_��3+�0�-��;}�:������9�*�E0>J��C��
�ggq:됀��C,��
��ޠ�p'f���"s�	"�y/*q�[�W�n+�a�Cze�f�;�
�NwF���7��j�Ē�� �Wŷ3�U�C3&<u�L�&���;#&���b�n�f��o�[�����w��!>��º�7hS�}|(���bހ6c�õy�=���*fw�3i,T+t���G�[Z��/;A�-c���X�̕��:_]��n�&�o�Ǒs䀽evc�&����B������6/��D���)�*���Nu`B��8�[�tr"��J��Zl{]��$)fh�ʭښ}s-<��;Q�6��3��J5��I�P�ǩ�k�:}�=����-̷���r*�ΰ�N��#�f�)�6��֜��݆�Dn;�F��l�w�r���(�\�����p㈭I|W�igv]qT���t�-I��[bͭ�I|��tXiH�)n8����ڬ|9���),�]I�������zzp��U���G0
�ޤ"�S.~��J,�1ͷ�1Fu�GYcΜ[L kk6�ǎMn�j�mL�����q�l_T�����t����GF\��Gw=�+8�<�n���Y��]�ˇ H$h��-��#���,�5�@��^��;�KYa�pt��}�V�=��k9K��B���y"�e��z"�(�x-�=}�⽀.=x�A���垡�J�E)��!��#o��S��nJy��ZM�z�Y��U�ptsy���@��[zyX��u���k�Mxō���D^m`�O�4��<�jz��޹u�=(�ú�-�k#��(�9��<��Z{�3��ڶ���S�J&��4�1�0z��@����f���A_f:¸��D�[1v�CA,���uf��N�C,�ܸv���I�D���U}����X+^��~���o��neZh�A��n
�Vl���cz	ɡݹ���1��`�ͽ�"��'{;I^.��,dq�[[�Vژy��6�����1لq��5������齹%J��5զJ��Ŗ2~��v4��,���56��쨆���K _?�z+ɚ���o����H��u)&q�<��qϊY��7`�o��>�����^�u���<�{Sڷ��.���S�75a��`\_���F#PMt/g�V�Si}���w�a�'�l�`�]Ͻ<0�"�U}���5�=R�����힞���&>C�Xa.n��iO��=�LT���o�
�/Ї�u��o��h	���.ƒ�\���U�����U�j�w���B�ʧ&��B��GY�o�~��?�d@^�����U��n#�7���݂o�^����a��{k��)��b���nuȲ:�(���Jꆿl
��P׬�c|M�=~����Q�*��Ӝ�!L#�[<G�g�~��K�ґ5�|�!V�B>&��1�Q�����$l��ne��������t&%�L����������vu��DS����oҖIxꁊn�Ù˲���/�+����l��=�a�eQҍ��meF���[R������O_�`�u�/�j0���[�s���{�To�h��Ƥn��ۋ_T�ͣRL۹���k�U�p][v5�����H��������NŶ��9.���蝭|T,hLc�XCc�w��,���[�
ެV����ؚ	�fN��+���P�O���y/z���ޓۜV�-ޑ�r���6E�w���6;ݓ�t�y!� ���^:\�����5{����t�������,�_���{�ם�Ň��q�Y�'���eV��K�l��<Is\	�ed�U����9���d7�iDl�GM�)
}:ש��r����V���ޝ�(W2�o�����mL��َ�wDs��`�ݞ�/Ƨ����:0m����B�c^^|.��� zm��0$a�Sz��Ƕ�W��=mo���t���$m��P���|��3>��2N�x�M�Nf\
�`�i�Z�[�ĉ~L-��O��>�p縶<WnܺW�8e��sɷz(ߍ��|��R���/��UZ�GhXNH�s���+�xyoS'�^�����/yw�'O��a���e��)��z�/������y�v��t��@ �sx�ץ)���(�5g:�w7k�t��ux���쩣��}�F'�gʼ�{��l}����0����}�.$z�`:�۞��5��ŕ���
��K��*�m\�o���ζ�d<C�j7՚����＃�_P�pVՙ���1��Dӭ�p(��e��q�ėܰ`��a4֐�']#Q�9$s;��<��[����u�m�Sܮɜ��*k[o������0*�r�����6R)dw�o\�1��j���m&A���f%ղr��ë����կ)\B���~�;|n	�o�N��_p�U�m�DQ�5|A�ju3������UH��q�ue��	��ݨȐ�����ݠy�=��<��RU{�����/_0��}Ƹ�z:��"�#w�d�:�����N�C��C^[��pY�wP'H�ga5^I�$���dM�u�����^��'Mǲ��ܥ�m
U>^e�iD�ò�{�~L�<�F�,'�Ԋ��N�/'���Њ�6��]�0��垜:�¶k�F���!#}��n�QTF��\ߦVp��9�=�b��!�����
��/c�|:Z�d�;���:B+7y�w(�����55?����z�����}��z�#�=C� 5F�'F��E��U¯{Y�3�?X��g3���6f5�~׾�:��:_@b����u����ҽU�%�,�0�e��_mC�C�O=횥��M�aAX^Ǚ]]� A�A�ׂo����޳�r�)���<����u��;Wl^��!ėu�=�Xi;0�kε�y���g��B�#�����-ʘ�i�.̹�H��G[�nlɊmM^U�Wor�f��MU�뺅n�ڽz�d� H3]\�Hj&wXAqa3���y��ŻYfn��i\�'��>X\,�wN�����_v��v.mn�/�����!c<"4o0�˨��a}�M���9V�IP����}$y�G�'�-�l���RJ�ӯ����K������!i�Ok�E�yػW_W�j�q� ���M>��J�U� Eo���~���5��� O��[�ݧ�����3�{R�/S�#Y*n�[���ع�RV@̷�MƋ�7�'Y|��YA���ݩ:�i��F��oR<���M����SgoU����)�f���m⥔c>����<�i�[~��z��/�����MT�UϘ���2y<���ي]�]A�TӦp���pc���|~�}^����&���͸�UeR��^�p?,���󓓅b܎us0�׳��u�v��c�E_y�{͏g_-�G�
 =@��O���%'�#]�~1����}���A�Գ�s��}�m��Id5��x*����碊7zy���*K���/����A��׈g��g���cg>��x������P�h��pY�-��3L����������s2�E�`�M��J,)�u_����oU!%o?ED���V�xּ˾�iPq��4g__5]Ch#���w᳍��S-���e��'�m�m�!�n�(M=)�WvH��'Oh��؝�Y�_F@��v�<�Oi��-���h9 Ϯ+)�/��X_1o��)ү�5�]>L��I����aY�0�ԙcPe�OޘYyn����x��F���
���h��[�l�ك}˝�y,�e��̳6?b����fhn�~��w���]4YIN�- C�Ƶ_�8C�q�Co��u�@D�4W�J\5F�쩖��
s��k<6be<򆒀&-P�n�%j�̺)f�=؉�{����ǔ��;W�������ʺ�,�G�*@*]X�e�Lzf��_�k�'��_����gJ�wް��}*�3�#��/i{;O�)? em��Yj_�-V9<�H>��B�M}^۫�����ٷ��gՊ�����EG�`��u�Z�\iT�6z�<�`�;1a�=���}��>e��i�F[!�Q=h���R��z4]���{靰�h�~��D��*�q&ݷP�����ꥤ�	�ɸ�����N�/��,m3�U��Dq��C���7�MӵQ^���c+��}�����8O��0���n��e�~yd^+���{$���muZ�΋���}S�^�b�������aMV�m.���s�ShK%_!y[)^�������A��7Ft�;J6e)[��wD��ó����h^���h��������rWH��zD%����^_ �k�g�9�nߟ,�LE�o}y3^��j�=׏P��q�ޯ��CG�����R���:�K�9����[��g�Uկj7~�{��J�n��'��̵��P`[c{m7�u�ޯ�u
���Κ�M��`���,X��4W�p5��o�ٛ�S�e;ʐ���\�����I6\W�$���0�^Pj4`�wH�vx�<pj���_eY�!/H�=S2z�սs�s���x��VV
�ܽ� �=��
c�d�=��l��D�]!�̍�g#QoU��=D+9�:�j#Z�,�ض�U���*>�J�1_K���ӆ����:��N��;�H<=��o��;u�+�/ٓ5xׁ����08p��M{���Vq����R�^�v�v|z'^vZ��>Բ��Z�X���5�MscҮ�����s
FuL4T���
�� j��,T�G����᷏�~޽3���s�~g�S4�yvA!��w;�����O��`�����}���!w�Zg�&���ۑF{�8cFh
�;�bu��o~��	�b@p����A��y�^@�S��6�x��mǃ����.<|���U�OQ��b�yPD�e�ٸ���6"�1�s���8�wF���狘Ű>��i���Rfp��/���ZtN��!iŕ�Q��=Qݡ,F��QS�����֢2�C��M�� �|�	0ok-��Xʌ�f�A�2��+��l��^u��g���]�>(����asyF��c��u��-�����D�E���8a瓟�=n�|������k-/�����}�'m��/� m��څ��m5(����K�;����zg�5;�w�~[F�O����4�=;��{ sV��vv�^R��7OJ�:t�+=�tw��;߼}�=�]�ۚ�獊יu��p�lpw�C�f�^nw�lÐN�N�νs_�b����7��F�C��0�%��5ߖ67��]�R���(خ@3���S�ݹ�GZ^zg�Z����U�|�[�XW����vH"}z:�{ܫ$�5�BMi��ש��wYY��r_������$^��Ǥ]��p�wY>xʩW�Ns �^���\�h����Mojc#C�0�����c��=��B�Wh��h��@�{�+��O],��G�ݎQ9�7s�2�T(��ǘ`�Ȇ��ϣ}�	�NΜK�μ��~�����G4/��<���
tѴr^�����hT��vƻŮc��Q1�$P=���o-�o�u�S���k�,�s����u8��;�M([eW�x{��&D���D����O�Q�A��*�Y� ���yc�I��[�Ĉ´����_KN�V�	�iu�������߲Ln[�G�{�T�u�����iT/����T��هaN]�7K����;SsOr��k�b��}��I�c��DT�W��<f	�oox��ۧF�z�D�<����;�]x�Zj�T��Ş���xsc+;�Aյ�ss���K^-N7s�q�8���En� �
��&M���J��{�۝��`���+4�FE�9�+�J��`�J��@�Tu�u�H4�#���w{�}/n�׮\�L������ؽ�{��\����9l�3ԭ�0��|{����ї~x!��M׸�Ml�R�-z�N�j�x����W�������g��m�[�/x�?`9���;*{5�G���kVE�������!U���+���Ӿ�^wj>}��&Aܰ�����Қ����/_�6j�M�ZDW{�\��͗�jZ�Ub�\�{��}ol\5<U�FZ�����]���ǘ�ǲ�.�;�N���mzR�L̞	��/r����;3l�W4�k2a���XB� ���Cư:=�B�W��$󟢫]�o�&r&�v�Q��P�5�J�(�`=�a�L�gV��R��,5� ����jt.���T�Yڍ�
�&�+i�l�j�h,�Qޗ�7^D�=;ws\�̻D�,���lu��5R�ef3_��5<ɫ�er�<�n��1�:��ejڎ���ˍVg#�yd��"�H_��|�8ӏ҈���ul�,w֋�/�2e�,�&a�J����|���2�n�?FE���ΪA��A`٭rW��cc���ˇ��Xluɽ��˯� �$6=���g�,�w"��bi�)3 �x��92��r�O���ݢ�@zfi;;u����A�:A���|��ϲ���(�r7�:ձv��~����+�4�(=����fUyɜ��r~�TOr�M� "�p:��ny�^L�����������A~�P\s觲�_?nݞ/$~�-�[��薨af]x�ף3��qA���pe�CA�U�ͳ[28��w�pO��׋��͒q�J�}zn���eR���� ���J�eN�`㮆��,Xp����r�[�(����kN�>�����.A�2y!s kH�a��/	���Q�~����������u����;-yg�y��꓎mOc�/ܕ�/*i��Ij�D����G'i/��ӿh���론�b�/�X�^н�a�ʀ��@�ڼ�e���#é�m���=Hҷ�;x�3�� M�ZE��ga��a�u�bl/�ɕ��n�}�����nS�LL��z]X�Ub�e��X˧P�U[��lζ�t�]������~UN+|oQΣ����y{Á��!�����)꣞˩�X� �[�
�]��Q�m��9�}_7p�Z�Ȥ��^���ح���&7oW�c��.�3S��܎-����J�r_>��uo�e�4:D�y��[�b%)�}�#�n�FV>B*��,���t]Y��%`�������}-#�ՃD��O5�y��[B�U[�j�P�Z�[��=9���ë��L��s,aǺ���r���!�[���U��j����.{��oWK�U����]�m��ː9軥ރ�㗗=P]̎��I��7^��M���#���\Hg�/��{�Dw:}�A]8�/����K��Ec�WL�K�ZB�Ї���SF���D/ee�AI;���JSpga�l�U �D��f�V�7�{��i���0�����������^��ʄ6�"��!XPX���%�\��[V�
�xto�]�������.��[[�^6:��K�E�m��z�SЉ>�Զ>y��>ѻj���V@�67�bG��6��ڳ�O�Y�& %:m捬M��^�z�\;d��`E�ީ��՝x�9���^���QQ�{�CIte]ޖ�vQ↣�YC :�j��U�B�IHV��̋u�r��V~��,��9q�Y8b�Ci_4,�^T6VD7F�#ϹොžT���%�c�t|�8v}f�s�薨�=i{T����!���~	�F�6�Ю��)ݥ|6t�+���ȳ��K�>H(ě��i�9��Rf-2��_}���[�-�Q�����8�����'w/��:y��w��s��j$/i�W5Cud�[�N���g-�n�_b=Uϲ��/�����व(��^�7��U}G�6z�J���(�9X���2�"�][���C��}��rČZM�2g=����Sd��Ʈ��s����+4&��{0�|��-�È���F���:v%�K T���qC�#f�{�;���Uv��j9�C˽�IY���j�<�Ij��]ھb;�wO �s!@6��ۻm���hs�0���}�,a��nB��mJ�C��8���Tzw�Y.l��-�f�q:ۼ�(���	:�F�I�oS=P]��c�\��Afu&�J�e\vf�Vo2ֱ}�F�#w���v����mNE<W+�|�x��w��8���D��M�V���c��vm�ǰ�]�Yz�A���U�Z�[ME|�[�V+�K,̬$�$��j�0^�x���z嫴���7�E ���Վ������m�X7Ê�hhsD��p�/2���}e���ƭT�꺸͞�-�y�Bʋ٧��}�c.�s���i�c˦����j�J�K����L�gWIT�z뻑�Q%&7�i4�'�8@��|��t�*f�TuJ�-]�Z�.�ZȺ�c��ص$���8_T��)l�WAp�<�Uf�?�'ޒ箳5����~�m���*�)ҭ��թe���Gi����Օ��D�ڱ����w��Ϗ1ۓ[�C2�°|��#9���hN
��a�YW��mZ��\�`������X�k�%cݦK�ɳ�����z N���k�ŝ��&�u���4!�� �U�ҭl=�9�\�y�)R�T�ͻ�q+-�S�X�*Sh�f������v�_Z�f�ڕ���P�N)X�.c�{�J�\� ΋�3qh���]gn��(�moT�u"��1�]N�C�DXb
���<����;���5*�X�\�u�ށ\r����RSvd��fϮ�8+�[��:x�ՠӃ-.�y�s{���.3Z��q;cJ�����;��}���6C�%�B[��۷;l�.�͈���Y�����iv&�ȡ�H�)`�7��#[G��3-}��ؑ��cn�����b�������U�rrظ����9�}[q8�$_�vrl���Ni8�r��{ #dDl�FB�4W ��Q��着��ޠ�ԱW�/��|m��!%cv�m��Hp�+�ϕ$�)��,�	�SM1M�L��,�Df詵��ۗ9V�:���!�d�J�'��֯�쏈�\Nq����p�xh��c�9)��57>#�����F��r��7N]��{{sK^��6�l�Aj6�wĶK�⚵�I�����Wn�+�q��R��N�^����S�]��~�34�C�� EO�wN�I^��{^�|���s�U���x[*ج�.�1f��F�s�Pp�:���{Ɨ^�� ø�` z���<Ժ-<�j�x�ׂ1y�K�s�=-�	��^ߦ��o����RU�e*�L��w����.�N嫛�^I�V��x乊{�6��^xƟAW~Џp\������i1t=bD����yA�\M�ϥǷJ�.�dpl���`�O�l3�½���i]r��sy�x���	�٭:4/h��%����[M�ۣ**��,6�N�(S]`��d����/v�K��
B��>\�{8����a{#FT]8�;�}�u�jw�0��,�P�H��X�M_�k�'�����3�W���ڐ箎ΓH�����}���K��W�[y���6�U�������ٳ�� 6o�ͼR��mK���y��d���rA�;�fma�F�S�D���uG��2����cWA�[��p�zM���V���8lK�ښ��W���6��9�d1�Jd�5��L�SWn2/��a���FKC��Q�L�^y�H�����_�%�ʀ��C̪�Ģ�mmJ�)B��G�yD v<�;[&!c�c����g�"K�eIҼf��[r�|z@�o���5�ܚ<Ȧ0�@�Y��a՟F��� 4��u���J��������w=&���xU$}����Ӎ�	WOÎsb�aq��V�߼ekw�qVwp#З��R�nz[]oK,w�w+Q��$Ň|[��묺����Ǣ�3W1�IR�ݽ���i>���]�Ʒ|;5�I��MNY\�}w�b�:�!f!��ۯy�\1eztw:���V�K�*�Rtd�7LN��o,ұ�=yҹ_&�5����p�,��
�Amw���@��/��bs�u�e�~^�\�{�s����"�~�=9����-���WO��d�������]i츕�J�x�4+�7����`);�W+���(�ӧ����i�����=B�(F�;����T6N7@̺!R�׹$��6��+
�4Z��Dkm�<��Bb�6��K�`��[���Y��Ԭ�L&��^+��}�_b{��G�:��o(�r��s6�2�tw�J�7R]��c��Hm��{�v�ȇtAYr"�>�4357��p�R�'GӞ.�ף�"�tյ��`̈́��v�:݁�,��X���f�V��9�s�#�g�Ӆ@��<�A·��
�� ;3��4כǸ�;�~��: Sy�
�ɾ8Mx�匦T9��qH3������{���퍵�q2>}���h�����;���q�D�.��~/ܸS�4sVv��]����y�
 ���Pd��c�����o�4�=P�gk9>��
�D���\}[����I-�!�C"��:�$6@������]'g^_U���ܮ��|n�k�}����_/!�i����,�ic�����q�T�țx�B���9�bT�z�m�<w9��;/��g�����q!���bK�F;�38/j��.�W4�Z�C����/�Rgx��Y����*\��!�$�
c����Qp��<�Oat�ǲm:���L5�{;;��(V�P<я;Go�z�Ƨ�	����%{��ҙ�soM��vo�{<̘�g�
�O���j�TUaۤ�Һ����K>.T�B:zU���/(�^N��0�G�{� ��o,Ʋ.��8��8�0�(��[��*7W�uje���M���mm��h�!=��vi����٩\,�1�
��Xz��c,G���N�R�f&9s��NKRM���\��������/\b?W�z���Ս�l���ӫ]�ygb=�ڮtxG-+�mk�
��SH��1)	;u�y9���k<oC���E0�W��cݵG|X�N��r(���`L��֩�ӵ�r}��:�dY�~9��U�;�lG�tW�e�Id���$]��g7��-��6�i���)�D:ȉ��T^W+c�o������e��M�l�D�N9+Zx�uJ���������Ļ�J���9��Kf��g8(-��ć��>�4NQ�x_<l����n.��x;�6�͚1%�Y���;��r.��R�q�������aC/�1�5ۀ-�s2%${[�����ݙ;+�b��)�k�qU���鏙5��ߋ��L���s�Ի��&��^�W� �bޏi��X��Գ���0q��Ӻ!=Ðд�Ѹxz���)̱�I�H�S2#@y�uM��:���A�Ӕnazz݇\�-t� �u��Y���ƻD��պ�x��I�����E�aV���f��[Y�=D]+!K���:(&�d�co����ٕ�b��0�֪mp�D����T�!��ӊ�Z��ΧVb��m��u��gp��&�5;�e�6.�v�[�oiX����!�VZ�Ӟڱ�=���#�H�b��~���(g�ܞI^�W��T;9�����R�@H=v<s+�my����aV������h��^���.,��<�z�}��w�������r���క�AI3��9���zd�ȯl���#<p���K������$��T���sZd>���	u��9`����2���}�h��\��㔯g�U̞Ѫi�c{:+����~����Y�Q8���<�[�PdW$<+���Vd�t΃c��f��G'�o�_�V��Z<�%(�0Սa�����A��jw)iZ�{F��Q��5d��Z,Ўc%Oz����/�����w�3{z��Vut���
�0�ro]Z��P�֞�ط��|�˧�:}�m�~���-$,d��YJ������=(.��I���`����i)r�Tt�u����j�ռ�T�1��}��'7:'����~1:]�'��%\2��VW'��9$��1o*�j���R��%�E땶�v��.>��;����$�S���;PV��/8���P����W���,�v�c��m��B�	\�t��Z��p������ˊ�b�z�`�����}W�s��4f �f���[y%%�@�&�T��r�`/f�����#�y�
��uL�-�:q;=s�]��EwΒ��;9oe���݄�O���L��ֶ=�a�ΩG�?����a[n��pig+<��ǲ�����.���E�K��[NDs��Ƈ�g��K�ޔ2����ƴ��\}���1#��BelMH�~-D�|����/<����b��{7��,�rq5sۙϲ��b�ӅB��Y!m,n�v�1�����|��PR(`��թ�է����2���d�&��?U�`��D���աm�K;/y�7QE�//�~�i���>k���4#!ԙ��4Mi�`��SV:�2�t��;�A�av��9���|y��{�	yf��V�Fn����
�`-�>���~!n���T&&�L�*˩'-���������?$|V_��j�}pW�z�ʹ�,Og�����+ޡ�����v����#9���V�곊�Q:Y9�xE�+�"oF�b�����L��7�[KАF��d���Q���
��T���yҡgI5�P���{C�1+{��J���GH�HnEzY�Ǝ����^�Í���d��]����l�!r��]�|�Lar�[�6�RH���I��4�x�0�d��F&��6�)�Q�#���R	U��$�*3;o��Y])!b� �&vq��O7ܗEM*�(�7B��y������3��7Sr�U���ǔ������OӨ��'t~�|y��7"[���c��v���S8Q@�ye�*�f�o�{/���BǩxZ���Ї�ޱ���|^�he��m6��wuY��N송*�>ؘq��;��{A�/�י]Uc���W���UAvH��~��袳��w����a��!�c�EN�뽪K)D�̄��i{3㳟������fi�;�+(�4�z��/�Wu��N���F�
��ގ��y��Nmx�����n(�ϒ�y��;�i.����u68�,���vw�Wݛ֍�(�~��{�k�D�M� "�S+��ŵ����g^�_���샰�k�c�gfW5��Kr�d+0�ɭ�zW�\�#El����0�ʕ�sGr�Я^`��Ƥ�R�rKֻ�t�Ǽ��1w��g��s�]1o��B����-��}�M��Ȑ=�*|��w.��,���zQ�:�X���N�8n^:pF�_m������ϱLW���9���\����]���+���y="6�l�A�O׬�o�uK�+f�ޗG����eb��K3��Ji���]��T���.r$�kJp옍�DC����)�;2t���(ԙ���z�d�=7L�7��U�\��e.�;26;MRN�E�,�rr7��yz���f�u{A_x��k�h�;�{ ˋ�i�o"GA�;��v��g�f���6���XuѪ���V�*�4t����&ƽ1�!H�_z��4}yՕܩ��{��S�1�}���d[��mo���hj��g�W�g )�K���>���hJ�F��~l,��]�>�_w22�fv���;;TD�s����kP�o=�ٛᵞ�W�瓯�T��D���P6���
"+ۺ�>֬�gu��{o�0,��[ѓ��^|z�)#�`;�JxR�0棎�E[�����Ы���\u�N�8�������`�g�O%�y�u�����`��G���v�O]d�~�[�|��Wn��ZM��}�z�$f�v�wK����{����z��.{�G���鶦����ie�z�v{i��d#� Sف��A�wK����S�C8���B`�8����������}X��flc`�f��6���Z��L�%ɏ1�@�e��-@w���u�W �$�V�>��mK4��U�Co��m��B=;��ry�;���cʝ�9��fTo��y����a��7����f�ٽ}1�oD;�q�S#��t�\R:�f�Dz���Ƕ��v�~^jZ��y���Bj��z���;P-Uc�v��o3���ܐ�Wo�X�	���+��6Y���U���YP�,)��t]�r�k�˜{f��A��:�����Ő�}Ӹ��Gcâ�f��`���W��O�).��[k����^���+!��n�B"����N�,�O��*7쎭���=V"ߋv�,vx��eO֦wFw��#Y`Vd´�O�,��(((?��mF���~��	j��\��xt.��N�)}���*�nY���H���;z_\�H!����H)�K0a>l�V��y��n9���`�FV
��{�Z��|�5�Ѭ���( ��*�vzN����W$]��؁P0�2s{*�����7��q���gg�C�*�X�$���DA����y��Y}<7�ޗ�3��o�Gꢒο״&ă��c��5)�׿�QG�`|�+��j�I�*SM��(ؖ2��5+�2M�0�����]��Yv;��gF�W�!��U���w՚Kꎅ��%vHт�o`U��h�-";%���R���L;�$�X �ߛ��o֤�)�$̚���C�Z{k���j
b��]qt�'Y���.+������rm�l�B�\��3��wޕ[�t����-Oϛ��c�󹒉�}C�-����p��dc��tP��n�T�{+E%��G���Kw'��]��'�^y{?&��uu䝺���4�Č��e�I� �Q����־�(������c
ܛ>��X6]J�ˎޅgBM�yb�>�)H�nα0��s	����=��>>�̭w1ib5��
�����]�eq�*���Ȣc ^EV(�Y��`��F�V��gZ>޳��W����*�|��o~�M.a�<�%��c@��N�V{$��xy��QL�[�Cn,���nTJ�ږv��=Iz��_$��������F~_�k�y\%�_�9xl~�Wm.Ԛ���}sBӶ�>�9y�+3�fv�/'�f0r�&9�n�i��p�u[uC��̩�t�����cO{y��v��~4��+���L�S��ڏ�W�^��B*Ǎ��<�pk�4�_��rb��/g���	�5@�����Sy*&���ǯ0dOeon)���)(�G���?.��֘�gS5dyMe�lxY�c���c�ٛ�M�.��5{}Q�/R��z�d��Hw?m�uL��vS�z��=9j}<A�����;g�!�ǯ���ۙq�]U~��h���A���Δk�P�Ӽ�����W��K�����g�^��<����eb��D�:W([7�ݍ��;1R�G[�-��p`C�v�EFr���vd�/�f��<������H�B�8�kx#E��t� z��޵T[���#�Wi�U�.�R��B�.���������J��%��4*X�ЎI"��z��n$m�Շ�B<;+�Zg�ǡ��r;&l�Eo[R^����d��kQ��l��M7�u���ݨ�����{�u�5]��CFv�I���Ae.�j�L\��G�����E��3�����x��sE��kv�G4=����ܻ��P]З�` ��=܌޴5j��_h
����/eNr=H��ԧ�.�R�{��2F��3��qTUy��_
�n.�xji50+���od]L��.�q�]�W"�����u��Y����K��:���ױ]���T�{A����rv��xNV��JKjoCPO��M��tm����sQ�@s����߷��A2�&>=̴m9�U��9�j�ӣ����3}a����]��cG9��w|�㠜�3�T4ɾ�.��t,�v��x�7�Ou�[E�
H�ɕhu2S�����^v�xº���`�.��k����N/V��J�m�ʵ�W��{C�t�V��x��oR�j���W(+��l�g�΀�5YG���X���}����}�����wWw�u8�ݎ�7uj�%!�J�uFw�&:�Gd�$ �|��ᵜƾIe����&c'i��ޝ��z��y��|�4�BD�Ck"di�n��]'�{tQlֻWXb���� E�:*�f����
9����6���sN���qd�4eq{��UyDlHܲ��e���b�	ֻ�Ƶe�G�2�o��m�/����ZF���up9�JMځ>cxj����ǚ��:ݺ���Ri�K�	l��,�̩�-�DYH7E���>/n�铘��}�j�N5�&��t���s*q��O"=HV)oK�dw8�*�=��
�N���u��f���j���*�i���Ĩp;�j@�X�E���qo9��ׂ�� 4e�94n��u�)�v�'c���/�v���F���(�q�W���}Z+m�16��5�UH�+�jި�����2�N�]�kI�#�I�3`2�[EN�ӣ���N�`�3]-E��FQ�(j��;�ގ���Ƿ��R\�5�z:D*/C����J~�a�Kw Y���n�6�X�ѭ�g{7���0�i�ǃz����U�њ�/�򣪎��"N�A���	���\lP�{Z��;%��c�����Q�]b��<��N�}Z�7�b�ܔEAͼ���Jl���{S���]N�f��6�*��K�i�;�.bme�v�VtK�iur�n�q��qo+aG�����33V;���չ�w��	���dX��&CLr뉪�&!�	�F���;��EV��6�� v��s�7b]�����a`=}M�N�C˦uK�O���U��y�*Y��S�����w'�%O�`)@�0���m�D��r��w��g�"�=Y"��+"k=>�*۞;r�_q����w���7�u�M$���5u���0~��X]&��A͏6�t�×8��G��Uw(��gYy��� o���0�z$#���EDBS#�v;6�*����L�0J="	-x�e����]KLn��m�9�[�:'���hΪ�Y��g�DMg`up��^	���]���1ěs$�V`S�#���'����i��Wœ�ez����΍��;�������ۨ5 �c��١�G���tɾK���0��n3��G�1�}��`���u}���{쩉'Y��f�ɥp�G?V����
��i
��zS8K9���8���ecL����{������!��鬘�:u���t�Y�p�dV}�I[*sj�_`�\?������ӯ֊�<`^����0z|���9���~`��7آ�GyQ���Rٜ�W�x'gPP�ӌ��Zv�}�����s1Ȳ�M zY�ݗ ��
� mi�������_�U��p�'[_��iu��$��D�0����6�t�&�X��/���Z�1W����%���xEj;L����9x�q������_U�焑��u5��W�gmh�j�8 ���,}�hS�WA�Rl�_���o�si��n�"!c$]�۔�7�X�&%����=&���v���}���EdV.�
ƽ�e4|�A[�p���2����y�VX���UU/�9^�/�aȬ�4�:�
�ח�QeC]w�:�W���	�B�V�{�@9F��4"�����}�?]NT������:zp��>�L`�@Q���~�y,�����Q8�Jk��{��u�m[�r��?�M�iwS����U4�q�g ���T���E3OE=����dfX��n�J>
R����\�[����ǅM�>~�}��Ot�Q��3��W3�"5��fK>ي�j%�l���Ψ���:'��n���S�T�نo��tg��d<��˵H3[)���Qu�Z�g�W��X�_��Y�����l�ށ1��H�|�6�r�����!�)�㷽ج��]���}m�9y�~rn����8�G!�q�
�����f5���4==��^��n��������lZ��7;�N@�1�ڼ�w:�^{ele��N�x����>�t����[�:/�'�fͯMGM��ݏ�����*�ʫ�R�oR)�g� x���bc
�12"�Ǝ�(�r�����K��*���Q��4�1��;��;j�d�/Obt�e�m�+�B�r���7%;�P>��;d�U���vC�5E��V��Se�������m�1x��_.��cb�58q�g��S�S��U�9E�KVԹe�X��!v�e,8x��у��!]a3�8>�tǇ.:Ku7�x^J�^0���8�C��Ս�����6*�t�Qt�)��W<V�����Gb�OM��/��[���4k��<�;�z��bUt�D,�Ȋ|Y�:w�g��:�h�36ZVn��t�.09�����ҷrl�b�{cz+F�Lzzx5I1�e�/���,�8��v�O]���R��F�'�'<��1r�ʞ�~�Du�V��{n�$�U����{+�%N��u{bwS�	P�XqDly7rk"��J�:����w=^J�Sә�ay�T�(��q;�;�Zu.U�fY�إd�G����v��^���.w�Z��n�����Z|j��C�ϧ;�Ls:��;��Y-�LT-���fX�J���4T�y�q+��;��i�<hϼ���#��A�̽�`bQ0��В1C�Y���7������`�Ӎ�\����qT��C8�ER}j�#C�<v�z�J�݊�[��ˣ��T�X�x`=罇�/���@�Y[D��:ዪ��'��z�K��+�ewR�m��ʎ��guMݛ�'F2i-a�`���z=L�>�#�Cw�GY��蘭�1���QЇ���;��DVR��f���N�޾U�0��1���Æ\�m�]�nSb�P��2n�Ngt�C�
���^m$����>u��1�o�����ەd졃�`��ݷ[R�Wp<쮾�'��oz�U�J�b�(�{j��9u��W-���S�r��y�N��^T��)}��u��7������j�>�Qg�Đ�\_xP�K�U
�3f(2c���;�Q>�W���|+8�w�eV��6V�}��TA�l���h,������sӐ�9����f��5y.���������E�����y;%�]����Cv���+g��K���ڥ�px}��CG�3���K�^h]� ��z���V�`*�
�¿~0s�c�����N^מ����Mo�&���;��zL����Sۜ6T�C��T�t�G7vd���뜯58H�+!Zn�:<�=���M�i���/W�^7Yʯ��z1�Ũ�AY�5$���܎�#W��nY�n���f:v�.����H�~5�Dۦ;;�'�Ow4��	�/ҿb:�K��_����qM	���"a�ˋ%�z�W+�r/�!���"��#�i��/���ZR���|���>�Ǥ�3�{2�r����-�f��v�{c�=Cw+�G�b���J�\vd�#}%5�̪�Z�	�W1畎��ۆ���p]U�T�s	%�޷^O�	�.N˳�v\�f6��ԯeXք���;�v-��=ۗ��t�zj�����/&��"g���*��*Y~��<��o����N%���-}���)�w7B�J|�Y�����ӫ��I����F^�h�>X ��f�ǭ�pd����f��I�}�EE#�'9Ϯ<�����Gt��TN�ؕ�"չ��S#+wI��sg
��M�ʽ%�����V�i�_Y�y9Aдz%�43�I� ���}~���N*Ur"	�[�\.7:������6�����/�wp��=�	�l��Bps����y�70U]�������ئ��k����я�5��A��l�6���IQ���yG���۟G|j#H}�`�Z]Q �)�����lҭɃ�$���n7wD*�T��"��nN,�\�"��цcKMLZ�{�N��L�����@����)�\g��n{��K�W�jox�$A�rD�F��@�Y��>�5�x�G�<�z��!Ȳ2h���ܻ�h�(��!Y��Mu��}j�x��sV9Zky[�+�L�Q�A�%��'���N�/0��Qbx�ph�Ih�tˬ�O�J��F!�q�{S��e��s5�.ƍ��wۙ�I y�]�9fVtD|�l\�����tThm���Ex0�(wJ+��Db�U2��]lw�k9�Py�s��_D^[򸕀7�2��5c�+�4�r�U�o���3�=�(�n����{��6�Ԟ�O=����c�w�15��;ה�ɩ����*} r���2��ҧ.c��u�����uD�r�����Q�bBS)o�g�l+��a��,��ё����	:���.�q�&1�k4f�G�"L��>��z�Y�G\ �m�v
9v�ջU&ڌ�u��.N�%	K�'��L�i���T�G��c= ��u��od�B�|s+�rkʹ���Y\����.{M��r�������:M�j\�һkO_e���IQ��'���+�	��gd��I��"�d���zrNW�{*yFq��Տ�	�uL�6���۱�j<�S���Y�?$��Ԧa�v	��V��W�93nD~��ǈ~���]TN�V����0�G7T�s��3ASҦ��'nb�K�Y�ګcb&/���Y�v�@l��ٝ�\Z��lp�1�W�Qj���K�gE���C��;=��Մ�dX�K}��%����*��;��<f��>�Y��;���l_`qzѾ�9�{��w�s����E�8p�I�/�q�3�uo�E(����j�TMz���n��׋k{TaF:F�7���6/�
ګu�f�`���/������N���Db���Uu����f�:A��U�5Wy�
�;Ĝڍ,�T���h��b ��\�=�l�q����_�t���}$��Խ���ǂr��Yr��5||�!
"���47�NGU@����ڈ;آ��,@��� �����ny݈`�._zqk%G�7��g��&�~��k��kw:�yI�E+_*ts��ד��;�|I���xmf�@�L��%��� Adn��,]NO�����*�{zz�F՝X���ĩx�N�-`�ef�K1�b)`�E��a��`c�Nt[N�]Ҷg8�vF^����-W*S&�t�!]�/��DJ�Ν9~���^;2�k�^�ۛ\f{%�Bl��Ј79N���ï�U����B' �~UyG{���Ș��q���"��F�.�_�ǻ�R�,��*�3GrM�DQy� �o��|��&�EV�o��k��
ltI�ư	QZ��()�s�ψo�<�������&fr���ʅ=�8!��~�-�_R[|*��8�隑�P8��P���13������ũ
�6B*d^ޡby<����+���_���z��W'���|�X���u�/�(vU 8ǥ��S,�k--�.�ݽ�?i�%�?#)�5����V>������/*D���Sʹ 3�����_;��L�S~��'�u?Joϫ�cݖ�
�����W̴��ӪX�2}w����Q�c����3�"�ݪ�Nyz�V.���[���9�H�!����㶷�9q�`s.Q�F��U@^{;�����ނ��;*)S̢�Z�4���r� ��Rd��wb�^�u�s�j��jW���x��ֵC�� K������H�l!+��s���32�#���]Y>}�ȁձ
�IPWz�n�H��)F���n�r�Me�ߙ��*a�f*��Y��3�:�Dm-U��-���u(wl�U�WJ��if��#г��k#}(��1ejˮ�J�@�;�9�@Ŝ��툲Ġ��)w+|itorV�:�`�`�N<����.�Y�����[����bO9s<(��;6��G{r�3muѕρa9�]��E�̓�.+؄�*���U]�ӕ��W���^��)�?�#�Ț�q� ��t�ݱ����袡g5�XF�k���:���ʾÅmՎ��M�U��{�`k��G<�i] �x+<�i���b�U��܊�k��g�𕊐7�B9j������(����s{�+|9��|&[�6j��q�p!F!~�GP��|�)�;W����'���W����L�q!��Ǆ����yq!n���x������t�Q��
��� �Ŵ�z�P���h3�n|aS��w;fc|_q����'�3�/=W��e�]4-�o.JDE4�h�4��;[d�����U���TE�`�T@�F�j`p��#��c�#s9��E�H��
�*�:#z}��Csޙ�v~��]��\����Ϻ{|��+3<È�b��H�5��ng�3��w�.{ݝy�+��ϻ�K�]�)��_�>[Yϊ:8�����X_�
jw�m��гNu�#�(UA��C�����w��0��7�]��Jk�o�A�<���ݹF�4=Y�=����􅵗�Y#�l�n�TX�˄P�zb8�<�
��Ψ��՘��P��]���^�-��p�� yw�GhzNIn����aC�>G
�v�{�٨�s��p��T�&�s.E�g#���tM֎g8���!�:�sO�<1�e7SsssQ˖��[�_+VeBKά��U�'�@	�W-f*!�C���3:�\(��W�ȫv2�����t*s
nmU��X�s��d&��)���743����X ���/�u�U�'wcv�j��N�� 9�{��9u�2���gf{)9�"��sj�:�5e��>����AG�w����qͱv���O6��k�b�4�.{��,�/y��}b!�}u�� �:��7��{q.�b�*�%W�Uk��Q�}�֬ǁ����[����-�ˣW;��q�9�s5�oE�,e����d��V�z
�5�O_3u�^� ��W�I<v���U�ϔ,/X3�9��n^�f^g�sy����PM;����8o���j�	�ɯ�D������,��B��=.;O�l��m�f>��}�E*ר�膎W�r��3b��9g=`p��	��Ϳ���پ�s� �w�4bz�ެ��wg�nؚs�<QPE+�%�Q|�Vh�pS�QD�@��9M}}f&����Cƅ���B��w���c��cw���1.�b�싲�9"=��U	O�?.REd��Y�4��)0�Jk����ba�Cc}iz�o?G��e��T�Z�د�\�8k�x�ˉ��>��u`��D�v���y�����N�{�*+�2�A��k��Ӽ	wS;+z%9�N;n�d�G4�<7�����Voo
z��c�o5'r�K��\���R��ܨ��8Jٿwǋo���\�1��*�)��;r��U��Ib������B�wd��5�}��S�r2����Ҹ��u��7�u�RYͮ�F�v�U�J$ǻ\�p�oe�)��[n�%mu�l1��a�^J;�l�O��!�����eg�h��'��L��T���ǜ�Մ����e'<i�陠�d(���H#�OZmm�+�鈏n }�(�b���I�s�����Oĥ�Voc'FgIk�U���ݎ�&�����
�ur�X&jBf޼K'Krr!�N2a�Fg��nkp�=ǫQ{K�p�{#�B��RB��pl+�k�Z��XμY>%#Vچ�������'R[�%�<�&궯���?�5��8��ͫ�Ǐo����v�;��ci��fpm_�]��&@�Uw�*���'�k�g�Kc�̱g ��]nob���o}O�s�?�_�0�wV�B�ٛ[�8���cZgT���C|�P<�/4�is5�ܞ�ffR�P�������`AZc�sr�C8:Ʉ� �~��9q��O_gSn�"ڳ�ˬ�X�ӆ�a����%��A�/'Qm�\����bDd�R���f�6/���Ҡm��m�a���d���E�x��W���mû�
�],'�En�j�a��WW�6P,jAΨ��6���v��8�u��M�p;�*_Pp_��6C�}�t���+�CWf	��~����"Cj;Ⱦ�k������,�:��`|�w�;������!����Y��#U*us��3��VmX���t�ٰ�wT�P�ku3��Y;DV�Ẉ|`I_�}B]i��z��i�y1}�k d��<En� sP&�v7j��N�[�l��?�3��+�'wLBޮf�5��g�;^�g�ɐ���Z7�\F��ċI%ym
'�r�/H�;�Pqo�f����ƽ�f;)�e<f�qJc"��ٙ��/��`�`5��*����z��Hѹ�8���5�=�0�j�	��f��8Uv�)~��F�U'T5P�6�Ԍ!#u�UVT���sK�ީ8�/��띭�4��źc�Jea��1�<��9c����1,Is�wf:U_}W��q��n�:���L���)$*[M�XӼ�1D��8��9�ɚ!�#�Lr-�x�j�6v�:�|��5�W�9��*������s] �
`B[\��{������X����r�}��"\��˨�S�r}�4�Ǭ��ȣ���;h>�s�w0�H�9Y��('6��t����%噄*�]�H�Yj�D�M�--�j	����Ͼ��|u&f�C������n��� �����uU�0��a�vȪ^�F�2��(�����>�,&�]U-�<����$�je���4_[���۠��Z�_}W�p��eS��ȔBƖ�q�8�ˣ�R�;T=�dU#�0�W�fs�vǴdk��7��o�"�c��-B�� b��Y;z���Ьn�agӷ�\��-���S�_W%Nc�}��_IuV�e9d$� _�WEc��4��
BG`Q��1�2���ƴR���&�ǒ�s�*�b�0.�[؟	.�̄p��G�\�^�'�-�[�V@��6hr�u�BV�d���{�U����LS�)h ����WQK'�;*g�	�r�ޜM��c�A���� �\j=�?	��;���eLV���ꭺ��J��� &	��)0l��M�9���J�^DQ�0���f�_!�Q�45����W�c�fS��(�+,�ŷ]_��V��FJ��<o<�P7h'S���]ħ�����5ޮj.�n�ҖX��̫�[FT�cn�Al��������Ӕ@�r�%p �R��͑8r<J�GOe���^><��k�ڕ):c���KmvsD�0�Vd��[�H�R�ۻ������t����,r3��P�a*M��u`njX:�n�˵�\��馯�u�D@{l�mv����M��C�P"^�R׫j�n$����#CZ�Hq��)�ӫ�yڢ�FĴ��`�u��@�
����d'��](*o�խ(P{ȍkcǷbjv1����:G9+VM��2�{�i�[�@��b٪pq�%orn^	V
�8K����@7�z�9�/4h���Ht�*�����������Z�F�m����O:����Eq �e��^F�W� �}�C�^�^���5�H-�w��䓭�m���^����e��r��)b��oZgB���l�S4SN*Y�8��ү�z�����ۨ�g�Ã�2=J����k7:�Iӷ�i�:2c�2��̉�\�P�̕e���{�+n�i�g�M�A��r��g^zc)�n��u�L�&7k�������m^zxV�D��9ս�/mp�e|n+���(y��A֥�u�跚NK�^��U�Ɛ�s���.�3��~���Vss�_0u̡���_�A:sЀY�Ө��DWE����1o�py��=ǫaś��F/y2~*/MhF.�!�<�@L)��n#k���)��'�M�K���]����B�B�۳�"n��J-To2OՂ�����U"2��q������)ԁz�U��:�r�4*�{����>���G��}�^�
5-E�q#2�5�.����媽^�>�ۊ1�)u֧�H(�i���9ޯRJ���Gha���ҿd�q�+ݾ�Cy�7�.�{ւ�+{�!�2���@�dy������:����f�j56z���l��=�l`�UQW��ga�Xg��iױnu�����'�l-r�V��v��T���ι�Գk��/�9��众Ԫ�$y*T���OU�aY�=y9�/`�9���'`�����>�K�ڈ�~���;Pk���'���8H�Ҍ�n���\M#��k�Q
�`�܇UaF��5�s����f.+6���x�Z��-��~��(NR7��3.'ڏ_&��E������b��+t /��9���K#yF�z}Dj����T�tz7��vڽHy,���|��!X��>���Ì�z*s}������^j4��<'5&��r����k/���ig�Eg]�/�8Щ����C�=���&�,r�C���ɯ'%d� _#�s<"��r�r�^n���X]7ڹ�5��!B��]/��Ң��h��e�S3Z��w 2�Q&�>�6j8丐��U8�Y���9ON���T��G�,2��~�����������}�B�"�E;PLVD���l���wQ��bw��z�В}���|&�^z�]�)����c܃x���F]�-�οoUm^%�҄�'���^G7�vR���}��I��caT�U[��/hv��V�=>p1B��=H,e�3R�&b�c=`�S~��We��ufGlp��_�%��xVZPvH���JV��6#.n�#��o��tdk�N��I��W�ڞ*Wn���������c#�݇��g�k+]�N���=	�:�<Ǟ������m��nE���P�Խ�v}��>��S>
_ya�n�@�	�^X��IR
'/c��Ϗt��Q�YJ�9O/�[=��!�������r�_��x�w��s��fxr�0N��lu!wa�f��)u0���i��Me8/W���.�R��W�n��r�[����O;�s�DE|���L������0ff�;��y���Z����P�k�p;}:E��0-g��*��j��}
@�0�;	���QYQ�g������:(��?L�[��ޯUQ�F,�r}���ݎAes���jx�����I��R����ʤ.5�fH=|J;�g�lg���lȉ�����fvS-_^��I���M���t���Ǧ�U�-Ĭq��� �s3V��s�r�vCҖN�t(���!��^L+=��Շ6#�QJd�����'O�{��
�\= {�oފ`J�SW����i�9{��y�>A鉷=+ںo:�r�!߅i�/���1(3���*����7U-�Q��V�{������{�0�Т;ق���U�"0������L����Kd�d�C��r�`q�טC�K��e�Y��S��۫��M�6ń������'�x'M��(ʔ��x;��맹��k��:<'*B31�ݲ Q�_������6-f�.��>m�O���̓�=���gM]�w��,ﻢ�Z��W���s��3�,��#��B?S[��Ƃ�Y1�}D����:�v�G���}�}۔�r�:�<��n��U�u���1Q��ȖەU�y��8�1�[�L��_oZ��ĕC����Y;Kn 3�T�Pr[@j2���p��f�}�k��i�"��t,��p��y������.��8�pa6z�2�d�Ru��hH���W�fN�3z�ޒ�8-Y���sg6� L���=*j��8��f]b���W�BF�<����'�8���z����D�]Rv�,�4�x�����w�گ;��P�S��u���fK��l�s�t�H�9?\xR��T�w@���P���\D�E�]Rݪ��7���ݺ��Y
�� ��=�}�{+D�,�vjκ�v��}��ïb1{yw!>���b1䩬��7�̭�q�t|9�LDV��W3�u@��G���h���yߕ�ΈBH��x�����6s�֍����{�s�ѕ�6'S�<���UOk�)�e��Zۋꚜ�BhIt"��o��/e�]�`�|Ǫ��������m�#w�x�B������c��\��[�!����'<{�r����xr��35ᾂ#F�1�S���+��NU>��D�߮�y/uqYy/���.Yv��͓��Y�kY`��2 T�Vg�X�ud���)tS�.9
��o�����r���LK<<�\�e�^�^t��뮨�>�=�H(޸�+��47�����Q?fw����G�^��j���ݧ~8}!�8%e1��n����\zx8��2|�陿C�*[S1��3{ґ6��96���6Ez��w�׳c�ћG*͚XV@�����4,��.�t��Y/I3�OM����1�iumG��I,�D���S�fց�d�B�n]O�b��%C���Ua]Д}�j�U:km!��e�;w�زV�n`vP���l͡ƶn�H�����m�p���o�8-Zw�9[+u+�`bWO�E[�EK��nR�o�v���p�)�J���㓂C�mt�fS��Mf�\��OBNx.���\&�d��uy�oJ��3�/v㌤-R�݃S���i*�c�9|�z�a��Ӵ�>%L��T��Svd�T;n��sRꖼ��t[욓�u9xpYBJ/E�X��M]�,τN�yT�4{���2�9�>��<���hV����׈�c}6�tU��#��Ԃ�|65�(xZޛ8Wbo]�ݢ�0����u=�Aށ���67�na�Ȧ�����
�j�@o2'e�H���?C��lp��j/�xa�K߭�v���#��]�ڪ��]b7QFK��*J�b�{3�l:��v��D��p%�ї0G(u=$S�U�ai �/�~���t^�<.�)S����ڟ������N�!.��j5J��� ,�8M�o��5ѧz��,x�GwB��ej׳��ïUƿg�k*�vKf����]@����`Z����`���e���p�Ĥ{�UՔ2�B/("��r z��'�9��1��*��Yk6 R�H�;�I7���p[xa9��A�%5�51��h�������oGIN��!�X�]���'u�hdZw%©8ki�ӓ�k��F�w����E/feUe���K�ͯ'S�$T�kJn۵e�$O�Z�S�&�Yv;C������9q�}{]d�&gf�]_��\�d6fv��hق�g�����ٲx���¬Q�w �:��a9��c�!�/Vּ�<�<՛z�*�Gs��=�&��K�GMd�>5�{u�s)�RR��bh��7���>�9�kݽ�;���oʌ&�f�ߢ{��3~�M^�ղ�Ҫ�0��s��Tp	�d��C7�5N�@�N���\�#u���{z�k�']���0��r�Goճ�v%��b��ƻ�|���«�ŀ�������2xu�r^�Ƽ߰�hҭ�2����W*n�9��<��\+��7����/�QB` �IVr�4���W9��)��[,j\%��΃��j�M��3���+��祠��2�٪	��A=.(��/�[t\C�W+Iw�[u���۸�D�f��^�Է4DYm��]�]N�y�y^\�w�u���{�K�oy(��묹���nn�� 7�\��B���#�x�T����`ζԞ���O�:]��'sw�O�#���_��_��Y'�k[�Z"�f�?Dk��N�oM� �����u�5PƮu����Z�D��V��K��eH���q�hY��t��Ԧ��0
�����J��X�&��aǏz��.�;'�\�6��m�$�^�g������1E��������93�<4G���RC���&=�b�B�@I�Y:"!ݍ�%ms�*�<�k/V���w�qn����#F�u��."���L�B��dW����ٟt\nh�@�
vE���9a8G\'T;��������6c�W���]u����q�桡�|8�
nM��ײ�\	�;��v(sA���@���qXA�Rq!���c[��ȉ8���M���j\Cr���a	[��g�+��9\�<l���vϧ泹�=3�aY����Οku�aT<�mM��d��M��3'�� i�9 ��$�Ap�d��B�څ1�3Sz1�Hd��r����j��bMdpե����uI�Pg�g�ݏ�ӱ�J龼~�,�
*n�U ٘��53v��6\�_���y��̚�>V��P�u���D���"��IU�iv&P~�Y���w0���|Q��δ1O� �OU�i��"��j���پs�����.��M�fJ���v�<��]�x��dO�/��@�N¥��Fo�.�x���G2������+C����ˋ�iyyE�"�����Y�w?Rch[~���Cw��[��vZa��3�=�ѕm��7*u�Eu�-�b�S;9�\�q��!�N�0Q��΅�l�J���f^��=��_5iq6+)�΀�*`ڽ��u6N���W����W+~o]�ר.�i�-����s�`��3%�Q���=qL�c_P'��卥ү�VK��5��2F{�8�Nk6�Nn`����Jyr��m�[��ߠB5 p�Bg�=��ֺ�.���K���l��������A1bd;3��ދ�˹���##����M�پ�G�/.���+`�n��W��|Ԋg�s��	cV/Y���6�ܽ^{1���P��:�s���g��F<���xm�=��/v-y�XU�1���5=���#�e���B���x��H�_�XM��Y+4���V~ֺoMMz�'x�Z�4�~Y�x碼-?[4P�t{���U�TK�(L�ژ4e�X�oT��+Un�<�p��&n-�l�����;��$""��λ�4}����"4�b�G:�
c�4UՎ��Q�.|,����|�-v�x�?�����UJ~�]�׶�=�S��F��Kͤq�5w����P�"�1[�ScQ���QY�=����eST_F��X�=v{�WX"����V�K.��Q5�&�}��=����Q {R��8k���7���:�#;��x��d�ŵ���M��pyYoC�q���	*�	b��9�� 2�	��WJ�4�2�(�S���O�����wj����(F�Ƕg����p6��S�D�V��܋�� �u��KV7�<��]C�́�[��T综���XH�}7)��z�3iK����M�A�qN"	�|=;V�/����8%{����3hpx�����q��c��Q�z���� �}�u��o���v&��������!Wрy�����{�#)mD����{WM�(Wf{×_1��O�U�K]���d�j��R��vb��&��I���%�`S� W�a_P�h���o2���ν�'6S�9��gFV��ލ}�Y{����[^��$^Sa���ޚ��5Ð;�	>��_�)5W�,��X�ƟaGP��,]F.:�Z���a���ge��&�ݝ[�e'm6tnfӵ��4Q$mU���>0�e9N�Z31
w�rV�r������&Dƺh��f����y;�V���������U-(�4mT]&>9�Ww��(�w2�=�4�\���u���#�����G��]�Y;Y�-he9z�o~ش��5k�~��u�-�)�-雔:�͙�ߪ�tk���7��KpQ��8B�O�ۯ����ͱ��Et��e]+��W���r�*��ǧ�L'G�PK�nn	���]	����f�^_�υ��&��c�+\���u���}��kb�w��%R5e#�/2��� ���ҋqG˘0����].6%_u^Cݤ��;DưkWzp����6V�7��|� ��Zj�ĕ/Z�,g[3)�u-��A�f1D=���БkiT�^R���`k�T~��y1���J��}�t������Ct��G�k��f�	�{`]�k��w��:�DH�ST�M��fl 柲l��\�f3Ȕ8�����x�O�s��r�I�]��26mӵFK�AX��Kx�Dl8f�σQ�j|���y
���0v�l=���m����{�Ԛ�B��\K����ގ���(*"����0aV���ſ�k�_�'��Hz�U�_�~ٸ��^JniS���7���T�#�����??f�
�Q��B�T�>��� ����)�˱9��lcp��^ݶ�瓨�>F�'gU@�U#�cE{����~����v�̥�=����C�fduo���*1��*p/B�3^csw/�;�+M�e�L���6�O|1�齰z?d���>���k["��q���=tq���PM^���ж �7�[������e�-���k+ �2��J](.}]�>57)�vnکzE�Q��f��-C5豽q�z�V,u�q�΂���{٫�K��hb��f�8���,�i�ø���MYʷ|X�{w�<d��1Q���P�$~l���2�E:�2�u���.7ǂhM�}P�ձru%����ujF�m�H���.��bؚ��X��[��.2΅�E�d͘��d3uN;L2�W�k������R�4�>�2r�i,꼀��U�(�&��<&NMA��X���D�����y��'6�R���s�}�I�s��z�9;t�۪��-��5V���]w`�uٺ�x-�a�&�E���U�F����?R��`c��0r_J]Q�ʵ�'.�nJ��U�e.��`�j݆f"l�wP.|뷖����S�7hu����!�����%Q��҃�����ͭ�l�I�4:����6�嵋4?�/g7������f�uRǎ�T W=	k^t�Z+I��<�8A��k����\Қ�m����OJG(s�Q٤e]�X��;����=Q����K��u9݇^-�M�ʴ⼡Jgh�r�Z�N� ��Z�V�+���Q7s����k�wM��4뵣�!3�4�����Oz*n���4\��CՊ�	r��k9��hM)t��3o�\5{cv��`6�Հ�2�wcy�N���P����9�͙Һ\��W;9t}��7�}o�f�����uER��UèZZ8�N��n�PN��IZՁ۽6ỵ́��$��c'�Ev�)t���r����K�wGn�3��@1��t=_W��~���mƷ�.�:'��@*�l�܋3Q��2s�Z��Z��,�\n!R��η�����Gug29��{��h�dN�
���o��G�ʂ��M��1�g��u;ݩX9plp�x��9��U�=I�6ô�7:��5�*;�����h:��ݗ��v[A٤p�5u>����[��ظfRl��*���*�]��#|�@R�o4��"ї��Cqǝ�9p#��;T�V����zrj�Q�h��t��n5�r�3|� �z�<�w=�k�mdN���~܆���\�Q���2���k�w�wv`s�Q�%��iŮ�S����4M�Y;�^I[Y�!�M��Emg�U�YWL��Q��h���[�y�I���T� ��>�mN���l1�$�������=�|�C�:H`Nݧ6��<��Hâ�-�.�V�,<��˘��/��=wS�|��Ki
ۃS,�־D�:��YE��/m�	���b��p5cܘ��[�]n��&�W�|��"6��@IF�7��jƁ�}���{rB�t���Wev�pk'��63L���t�'H�7�e[�ѽk���GZ��N�2�Q���u��H6:��b�g�����\�]�M�۔^��[�l���H���S�;�XѤp��퐢/p�n�[�C��%4��o�ڭwC�=����:�ޗ��d�/q%o��Vs�����)�Y-�H5��^�����Ok�n�j��]je��	�#���Vl�5Բ�',u���c3nrV����,���]n|CM�j���x�*������bҾ�fvN�d�b�aX��]�L���g�ԴR�Z9q�������ﾦ��X��%,�ׄk�z�@P��rL�'u<����+j�_qӫ-p���
�I�=x���Q5t�]�mH6�wL�l�M̒Ѿơ�G	Hg��A��2�c��u�eN��0j��֢�x�����ף5ߺ�w�]��K?I\�os5���:����T�I�Dtz����:󕊛��7�RMvE
������e���}���oҫo�ݶ�z�����2K4>�m����Lן�V�*:5�H�x����e�y������+�@~)=�����Tɻt�a��QU/��D��a����Lxr�*��s�=G*�|��4�K�+M����\�x�Mag0<'��^k��q͂�TN��0Kƙ&����j�ܓ��=^��w�!�	ús僩._4�/nB=\���_e�^�
w���.1F�h?�a�Ǐ���|����E��]OJ�v���E��ڇ�4]!�֝���v'?cS���W6���;_E�W��jU��ǃ�(*. �r@�.�2�F�+ƶ����Yrze+}Њ�v���3g�������P;�Vx���mD���w�z����F����P�6��6��&�_�\r�E+B�0�&�z��Ez�ׯ-��]������yNi��,���^��7��x��z���Rz�`������nk�i��q���'o3�3�.\�(^��J�����PVkg��7R;_jcF˳��8�Pի�[�8*Qj+��>�������s{K�����+��W�M���G��Хn��O�;ɪm}�:.�w�8I�ə��#��`��r}|����ɓ���<���e��ܟ*<ܨ:͋�:��wY�k�]b�K�>�M���U�0ܴ���7jG�f��}�ɰ��g&�ԛ�f,y���`ܼ;�>E�P���'����8����)ݛ�5z:�^��K �7eέԧ�|Qb�c��v{0q�����Xś`t<��-�Q��p��>����1��
��I�*W�/Ms㎡&`|�׵���e��!�G������Bw�t_�8M��̍��#>�n;�{�N��p��k����lgP��h�{��g]����i;��:��}u�Q�	��u�]_�����;�<s�!\�1+{��Pjͷ?3�W��/���4�^����A�i� �Y���N�K��P&Lyؘ�7��/�l&��I�=�7#��'���9���U��˳�:�
I�/ƽ�~�R"d��NV�WD���f+fDeDN�v�f3�LVɠ�=~�Έ��,K�8	����2�L�NNօQ�j�g��Dq"S���x���ǹ� n��S=�4_v)��� �����Z��y{����	n��ۚ]68kNvp�*�*q�6�u�5�q���Uo(��H����2��r��v����:�]^�Lcԡ�ē�I�tj]��>�|ONya GM��͈�?���l���>�+[��.����Ԡ��2��o}�J��r��6z�!*���)x{�硻][;�+c�\'ù�f[�S�C��t��gMGbCY萧�?��N�����.~.f<�+�^�*��}�,�M���	��\Nw�Y(�,wќ�3�Jn�o5�������np ��Gٳ�wuxO9�ӹ˰U��r�+!HrD�]PJq��ga��Y�9��;�Y�o�N��9��f����{��{D]�Nq��*�O�y�̟q��H�:vpǥ�`���F��Oi�B�r�y�o`]0{do�h[���g�u����ٴ��ޚ[���B5鬈�Bx���m�+qͫ>��X �sv�oi�L>ۡ�tc�#sb�_\��#|��3~8 Z��B��ɹ��}N�r������
��o����3� 'T�<�`�<#�Dl��Cdpg�Ꙩ�I�v���9�}�{
��}���u��^2�;20T����]�>C@������"�'x7q����=;q3u�^z�]����ve�Y+]w`w]�^����Su=��d���+#�ٲ+�Q3���z�C�r²Nϼ7�vlB�!��U�U����wf�V\P�ͩe&���HK����v������w
἗q�ƨ}�o>WVUf#S�K.Ȩ��3t�w��S�Ղ��h\�ԗ4���4䫬�^�_�q�\�Bи��Z���/\�j��T��e�B�b��f��<ίk�-�|��n�/��h^�~�Wz������"��R
Nuw;�]i�A]i6�e!@e{�`�N@�k�s������1Z}5�5���@�qN�����	{Я
A/�������g&OC�b꣍�[�/sz5�S9{Mß��U�מ��֠�(� ���Ojm��!�v�:�eS�8*��vn�:�uz����~�,h�0���C�v��4�1K�Y(��c)z ��=@d�}C�ΐ�f3b�>=����)NGX���iJj�#7�5St�x�OU'����D�Q
�uG�o|b�K�,tT%�q���Z_��s�_�Q͝o��o	b��y�2ͷ���[n�_Aa�K���>���v�~_����_�:�v�(V�~���yy�#cqX����+=1���s��Pq��S7����o��\̃���M��"��A��x��5��Et+&��Q6�ꓝ�T:!�E�C��ouW<��1�=��%/2�ʞkW����	���N�M��s�����6���n��97�z(t�s������뾞�r�>;^�{+!e`�D���;�&����B��ع�o;-ֵu9^0� (�YAwX9�^Wh裹����W
Lnar��x�.W��b�b�`O[�[�hU�v�� V�S�JY�Z�El9}u�M`�d�Ӌ�P�0���R�g`��ɩ��-���[ݣwr��� �6�ع��^�8r���G/fݩ9�а���P���q��h�^��3���+f%���R,�7�<W4.*��j.L���hk�o2�.�k��4����T��r/P��ٙ�`/Z���5�٘fw�a���x�Z���>��gk����e��[��nPkJ��5�t���e�j�~UwQy����p�O��
����˭��v1z��6��D��1 �K�~Gwpb��+R	4L1�,�uo c�m�����{�;\i�r�.S������D��V)B����q|8j�꼝�eǜ���2Z���,gDF>�� �ވP��4�OD��:�0s;p-c�|�`��r�߁C,�Ag#T�N�n	��M���$8�Q�d�v<[�?xm�J�i�[^�"��h��uUp�|�*�?#kb�T�clz���5�K�Ц�Lm����I�S�����߬��:�5�а�S�*��{�t9�>��싎��D��]苂�f�iy
��;ֹ��)̍�Ps���؀�Mk[�Xg]���T�>�]j��H"̌A?�0����V���	��wv����3�\�Cj�u���q�l��
_a�v�,��7�͠�ur�k�v����f]b͖���r��iU��5�T5����	t��91�wt:����y6ީc�g��u��˥�u��}
nh��Om��U�٫�(��§\a��:G����J�;'�L��mR�x===Z{-�]����6�豛~/�ېO]������dd6�{ߵd�)t�n�v�I��Ὅ��:c��s�6��Ev�F砺^��3��}��\�+>��E��n�֪���J������~^�q������"7�I/eF	p&w�y�K$_��\�y�H%�i@�y�J�f�:9�>����c�����~���t��vȎ�],|�~/@��o��x����~�6[�+¥û�?kB�6'�Z��OB����Dzn绍�̃��<N��EO�w12ؘ.r �uD��<7��Q.<�nD_P˅[m��Hֆ���Bӣ�������������\Q�u¶�A-K�{U	{y�]C�z��8��^��k�����,�����/e�@�gy�:/������.'�C�z�SMEՕR+���7b#����g�ڎф��9$g�>��;y�ś5�$�ŅV�{���C�J#\����#˫|{t�m�n-G��yS5�G�m�&����@�����.��Q':�����6�zV�6�h4��6i�§��Cv�E�V�b�qs��
���:�,�7m|�>N��mŀ1��ap�&�K�>���	�f�v{I�ƒ�oi9Z�R$f�h�(����v��s;l�ov�R绗��z��z�h�@��n��O��S�Nb���9n��Kw�vO��Y�l��=��⹕C�s_ợVR���8�sG�@�çv��w���Vq����i�2���=S�~��;/'��\.�pՑ�+��UV+����v������߻�8�L�V&}>ꕞx<�����W�1�M'���8>��Q�ԯ��/��w,��bU�������tzm;�lo]���说z����6f����rhYՈ!�H��kb����s���C[��VR�o]C:l�p��%�u<�[T&6�^+3��nn��N��)�_P�K�R��W[2@�%֩�X >��&U+�{�~]pd���-G8<&ęʬ$sSXX�o۴˩�"�����n��3MMnh��t#7����fxm�N�=�>�;�b�DFʻ��Q����7G�6�W�n�b����K��J=�\��B̈��z��:��MW���=g��	C�ו�b 4�����]&o��ɝ�9�YӅ��D�U��W_od�|Uulljk�<��P}MR����}�����T�f|�]��B�� �t-=#l��
n�t�v�o`�aw-���-�3����٨�������"�2�l͔����#�+��f=ދ��׶��K8�m2)o%��]Z�f^��k����9ڴ�#�����T�ʋ�p��ZL���7�7*\�Sn�]�;�k8u�ru�R9Γ�47iL^���%�q�F���Ut�#v�[9����M,�:<Ȼ
�{c#O!���޽4���k����g̪��%�M>�)�߇���U���
�Tzʈ��/���_T�g�ūj'R��L�+X��4�ұ#4o�a��/� S����]q���{���c0v�$��檅�-��J�G�ݸ��1)k��e�I���;+/o��qj�*2!��sի�ޝ^��*q��;�x��2L,$ʺY�'g��*|FTCq���
F�Uzg"�߄n��kmr�����?qs����"闣z}ֻG\vyGM}��9�w\����МJ�ȝ�Uٹ�W�u� �D���#���QV{L<p,�S'xT�	��\h��u��=1��o�	�}�R T�wv�xҮ�7k���}OkQ{}m�f�����\�?3E����ǣ�7�RxR�	��Pm�^��� �fM�9
 R�2	�0�p��x?zN0�o�����v(��=�{��|Ì��L��+Ş���
�.�������Fy�0�"����E����M^v=�O����?`�b�e;�g4Nj����.�I��Z�bƖrYS��F�Q��Y,�����hn���t9K�͂�>�����F��u���2m�!tRbD�V����W���ЏSlg^�[ǯ�Æ2`��b�l�ѧk^i�xK� l��.d��X�E+��>�~�m۽�,��v��@�C�oc�2�l��tfZ���ѥ���G����\�jF@~�z���#tqMV�������n58�j�i��]5���.ء�;)ZĬg��z��=���xs��r���v,2}��e��35]9'�Dl��୧��t�z��mv��I�CHp���:�NM�����m�"�� ���Mz��K�v*%��6moo��2��^��}�M�V|�=y��YKDs�N�nf�c��띞��A\��Ky,�4�n��s��>�Vvּ�����xv���^�w��3���C���޺�"�Ro���&f�@u�j�Ӯ���~�>��jIV&���j�-�S�u��_)��_��P�JW�&3�y�:Af"�7*ͣo��
O��
sƽ���0�z9��m,"2#���^���kw���uU���G�I����)���Ϋ���=~ku��^%�Σ���95L�=��ޮ�&�D}į�t���W�F_�8�������`R�yl=��e���G������=|3^�����.���O�p�5Ch�SS'�����{:�.�;���������ͯ'���Y��ީCQ�d���u��d3���G��{WZ:�t�*�e"�rɻ˛�"x����#��݇Q�pj{ �ql�.�wjT!E-6J���ڸ�g�J�q�n��j����N_jk*�Qm`�q-��¥���Pܫ�o��ʇA�l������C�dK f�mp�ĹH�q�4GQ�?G��b\�l������ ��]+pc����_�I�x@�G�g+NW-��
�����%C��JX٫��I�i�n�NV�l��&��T��u~����բ/f�8�A$��E�SAW�h�y-�6ixA}~=��lg������y]fg��ި��ث�:xb���EV���/�0�0I9�苬��MB����=ܼI��Cܒ���	H��Pf��t3�D+�Bq�n���w��lbx�iS�h^�Y����v\�S��23r�����b~�)�1���s�^p9&��)��*��`�c*"�L ��tے��)܁��h�bB��s��v��Q�:�mt77y����P������jorXG~�p=����jpk.�M�
<��f#QXs�ج�'���1��r�3�;���6|�kW�M�����h���q����5��d��Yeh0�n���mzg���/?O�*�}���]�ʱr\���\�J�}����LVǽ�e=~���9��A��*C�<�,����&�C���ն�ٺ��k�� u���Ϊ���l�Bv\�n�wI6ͧYGd�ݭ����Lfk�&d�+^i:�-�\pD�"������*ާ�X|
p�n��.�a�;>Ћ�:jIn�R{������ŋ��c��V��h6\��4�of�qv�-���ԽG�ݩoqj��b�r��V��)���V*�WƝ�r��q%�v��Q�ɛ���h���SY}�>��V	�q_}U�-�е_X�[�Re]�vg>��Xe��
�U���M���	Ou���DR��(�k/}]S�k�o�+DYIN����S����+CWX�"��ڼ9��+�U��Zz���ur�o�[�?p9>�M�2�ހ~�cj�Z�;~YM��Xb�W�<�"*�^Ng,@d�U���É��S�8�%��)�ù����j���se��W72rW.G2���v�����ks��G���g%ٚ�5v�+��S:������ørk�$u{i4�*S0X�H�a'��z����|�^;�r�f㿔�/�0��3N���(��M���q\���b�֣4��ׄ[G�^Zu�1����oF��9�TQEd5�0t�c�Sk)�WS�v�u�N�k�ۑ&�8��Eáf"����[Yۍ}�fE�8�c�8*�E�[�ڱ.J�ꃐѷU�Q�ntx1] �K\����w����.�W���wӗ=�n[�ns�T���	зn�=�,o8�eܨ'n��e�VvՀ ��`���SsD�P:;�A���bfo
�z7yկ���9R5'b�v.� \�GZ:��7����f:|G�`Y�+7[���֬��S��|#�XǬ&��6��m�w8�=��e-���I��8ګ���5�7�J��O�Cj���1]Gn���%�|Ñ��0e]�!��{���Us)��YI=�}{���Kl�����v̍���R�ԫ�S�Y�]%�jx���V��U��v��qs���=]v'c�lÜ;����ۇqG���{��#��P�Ő�i������Ƞ�;�ᑿ�^aݼ\D�ٓszp���3w��a�2u�N����C�c4j1��d���X�@v�0���l��������2gn��K��ٌB	u�m؛�r��t���w�wݵب�:�@k����0����p�j���uj�}��u�)ʋ��_�E��6���1"�n�F"�wU��<T� m%���X�)�	� P
�T�,B�NCo"Qứl�ź�����7�~z�o����[[����/2�eL��c!��%�P9���6���i�m#�Ŗ|1��YWك��`��X�㓥J�`�A
�v�������,/���䱕u�i�vPް\�E���4s��x�;����t�9ʗf����2���4��Y�mK�i_Wh���a'c�kN�*��1i�t�V��s6�k�XQC�Xߢ�,�V"�|N4�Cz�\��k6���W�`orU�o�<�EK�` ���b��-B}h%"������1r�������������¨Ct��{b��7�żA�;�w�RY��\n^b:$�2�`gs�Rs�4��p5)��L��;����-F콍�����dz:7O�u/{�e�H��j{��<!�W���衽s�4	��t�{��kKn�x,�Y�D���TGj�3�zn�7<�HSX�Y�a7,����ʂr�"����Gu�n�\�):�[A��6�x\�2���4e�~�=q�q�+ċ겆ʚ�~��׋*Y��,�yo��F�c�ͧ��G�i�v=Zݳ�:W���2:�I�AЭ�ܺ1��oyl���ꛣ�Jzs��v�%3�Gm͚M���\�\̊&#<�]�ղ�ƃ��J��mϫ���c����Y�]�y>C"2}[o��#CS����Pر%^���v��DVwm���/�"��mY�N�r�Bvg��a�k�ۧ��a�z��|T)F�뉬�C�Mؼ܇L{ �|���4���~Ψ�#�l�TR����NDΛ��k���f��Nm-�n���s ��/� �n�xy6sհREh���(�J��O_�G��up�i��w`�u���y�S������@�#0�<k�t���ܓhU�u��ʧ]tQ3��+1Σ�'�؋�aR�r�ۛ�KY�7��j��F�հ��p���	�l��PK_`Fk�Jϻ��<j����;���L����j�S.a���=dT�;�X:i��\������iR���8ƫ�b��`��4�2���b�֍��?���*���wJ٘Q	�(�4d��)L��Vץ8��%H����h���o��6)hFc�f\�yм,\����5��,�� V�d��ӳI��Ȩ�z"u$t�>ʋ��w'�j��ў�6l��K��$s0o̠	��DށS`����U������^ffye���y�t0y���2±��l�m%WZ�t�JT����{|�eM�P乇�{��>�ˣ0�i^�Z��_�{o��v:z6�������dB��Mܣ�������9�����R.͉�$?�~��2�2�w�wƷظu��:tdN�&�R+rh4<ɞ{2ت��:n�+6t�
�W����J:f����.C˪���x��~��4��@�Q= '�B�;��۰�/Y ����rYq��^�?��o�ܱ5�t�Ϸwv Wm��;i�.~{1�W?�K���9WO$�?���x�u���j����զ�)�^F���#���[�}k8.��4?WT�A�mU{�_-��Pz�"��*bV��8mEU�݅v�ǒ߿��W�Z�;��#��a%_���^��ī��Gg�Jv�d�a�2\���9E�#�� s� �9ͪ�#����yAU�ǯ����-��zl�Cw'��V�������+.�$��v;���V+PVmru�X+M�`i�Lu>�2��4�Չo ";|���7�A����ר�q�o�ܓ�{	�'f����*�\��}6F�=�w�b�u��{v�4�b*�>�Jl�f����	{b��т��F
:��� p�S��;�r��Pv8�w^�ȷ���}#�^y�ܴ3��W���ƽ˲��9IX�/�����.�?	�N� J�N�<+4Lxc��E-x'�[Vd����n�{���C��[j���Y������Mx�F �ԇ��a�4S�i��Qz���x́;��B=,��:to�mߪ/V��=[lo�/v���G��$Z��q���O�{]KV~ړg�PŅ.�C��#���U8���u��"�R�J��:�!�(��E}���ʯ��"'���سvg�s^
�T�̶Ә\���)�����t@��p�l��o3�9�N)����m������@�
���E�Pm껵{�K���4=���6<#�:X��U9т"ҼJ�eз#"`q�h�q�E��w b��3�+�G�.�����fҴ�j���߅>Ȉ�z�#m�1)מtb�D�n�g�dB{U�hǱ�S���#����D5��3����v�^YT���c�����u��Ds(W`%�/+ዑP�ek��fHw���mb�]q�R�"v������.H�hw�>�Dǧ&��7\�� ��^�9�ْd��5��#F��ŋ��͖����
5ŝ��YSZޛ��䔾e=��؞�3w�O�ۖon�7���.ؽܵ�=ٙ,h�O��/��.������{����Q㒟���Zz>WN��WV{z�+`ZL{U�cDe���Ĺ�4z$��.�6\g�� ؂��/�]���&-1_�n��$����9��zr��j�"��ծ�f!A���뼳(¸�O4�gd��;��1�V�J�Ï��r�Y�+�o�~�JNǋ���`:s9��{nz1�2n���9��Di�P������oNW�;����ʨ}�f�ۦ�A�J����]H/��[�ݧ=�[U��t�>$�kW���.�k����F*�zL]��2%�l)e9�8X�~��kΈ��ZS�$���pr��詹���o�iV�߁l���ȯMƎ�\�D����5D�OO��S+M�7����Ayf��#O���*{�s��sLb)-jm��E2|��m�X�h\�k1��?cV���t��=��ݎ�I�֌�yF˥���EdH7΅T@��6���� ���#����;������}�����ᾰػ���T�d�I����{�jG��z��Ʈ���x�"���q�t ӗ�)�x�ܱk$ϫs��8V'�Tc������w6�֦RW ' ��b�yE���ǉ�e�S��,��rU�N��i�LE��\��f�;��~���f��_�v�I7fX�~�ǹ!xS��`�Ŏ��	R�ī�^�ٿD>
�E&3%e����}e��� 秤�}�3�
�hBa���]w�d��O�"����m�9�c�=qi��klS�p�"0�f ��Q7�
�&� ��@��4M�4ٿ�KE�S��3��,��x��-=Z^b弪���N���W�{R�L�D�u�����u,��������X��)�:����A���X3v�O��p�ÆA~��W�͎�0��7��f��.�A�یǲ5�b�iM1�Z��uz��������y�ܔ+�-�l�H	���'lf���!�Uk�+���Ͻ3O4�ǃlݯdU�W���@z?fVD"&�����J�0M�
��.���fbS��@Q�[MɄ.Ǔ��.ٻxi\h�\�A~�]���٬/{4l��B%xP��I�VS�Y����+�ǧ���̩��R��y���V�Ò�{���ۜ$����v6���'}�Tk1���#	��S�>
<��-FѤB*�	H�#�r7Mrt��ֱ�����R��|@���;�C���.U����Q����z��Su�Ǭ�~�+Z���4D�k}[}="�����ζ;7�����>7y�:�reB�u���&�*5��e���S墰gQ=�l�������K��鯄�C���{�u����x5���uv�'��l��O�{��Xl�h�g����W>w����k�ї�j�<
�R`�{�,�N�[�	����H��*x������(<GL�y��ﵚF+�^p�<�ݖEw��-%Y��ɨw����f=S�t� �-m@^n-{;`�r��^�ٹf�W.�������3�����_�@c�ڡ���D
���%�]�
�\?V��ޝQ�8��z=���#�;�Lq�����5E��pA�R�ؠ�澡�d���5��7��+s���\�T˳Z+ݪH�Iw
�˜��Ei���1��8�����l�!�>�^9���W��FN(|#''ϯ��o���1Ke���QS�f�6���,C��d�R�U%&f�τ���h��_�Ki^N�w���|�;Y4��|�dR(�t.M�\�ܹ�9'uʒW��$ݫ�.��M��H�[fj����5OoD�����:ɱ	;S2��^�y �]��^�΋n䴶�k��V��&�h	�<,ŉC�MO+�J�.�\O��<�koL�^
�7(^��<�w�)�l�,tt^U�p[��2��a;IWZ�����:�v�
���vOU���ow���q�k��Q����$FF�8k�Wѕad�g971|l���铆5W.9@j&�7�1+	��2[�*�%�KȄ�����E��1�{������13��Q2vw���OJ�@�+� �q%�l��O֝���N�(�PK�o']]���ꓓ�f���?��N#��Ү�3�����ܡ^nk\�L����F�~���ڢ���h�0{��m�H�ξT���P�u�$̟�gv�Y=�U��ݜ���������
 WG{r���ne�?z�ICocd���/�����L��S.����c
h��.�Q�8}�N��Fr4s�$�Ct��K��s��FW���	]�2x�j��P��"y��L,��-�=!��J1������1�ːg�쬕�Un�Q�{hV�����~���\�~���H5n���畚�.���ʊ���j�W�$-�oԯ�n�{�%վ�}ѫ�Wv`jʭc����nzНց\s�����+ojX4mpC�ד]�7.����ĥ��j�u�;&vfO>M��i^���S�]�_�^�F�7�)�r��96����ET��zr���߶��z�L�1�2`�����J�#+�Y�"`x3Y��f�N�S�U�H��Ι�W����3�IxX$n=�W+/�<g��yd�q��+~^��0�^��UT�K�rkN���r; +%�u�ho�;�^-�@+4�e)&J�YOA�N���S��"�B����gf�=�s+��sd���W2Ӻh;���^�q���C�5f)�	Y��Eui$�b��
F��g.!ӗN�n����fug,qz�֖�UboVVc�h��F'֝��/�RQ����)�.o;n��w^W4��i�ׇ��ގ��I])��x&u\z/�C�gy�ý*��z2�)
b{:6����dK���D��߅WK*!��vc�;n������ڨQI���?*Vf,��v�a�n��>�����wr��cF#��^U����G��;_�\�,+�UX�o&F�S�#{�j�]�UF)S�5�G��hX���|F()���H�M��S(A�B=�Q4���=�Iw���kkO.�΋�\��Z���"��O�ꌘ�2;_��A��T���vW�GxW��J��t���^u]�`�۞�F�o�M�	ߠ������1�����[$-�W�t�^/}�Y���tfI�e�*
��թ*�c(i��+�s7��J^FގN��u��zHP`m��v�j�/�y�;ݫ������3?yjkI���w\Y��;1�~�r�)�0�>�:������3�S|�c��g��U��g�����9�U�*�N��;���~���9���1~?����FX���YWG�F`I���D�V���[]��jA����I���2�Z�&k�;/@vc�k��Ա1k�E;�J9;�׫zgL�1T�u�[u,>���NcR�=e�V�݆����U�p�&p�3M�3{�����H�p��Q���h,Kc�i؄GuK���ف�xb��y
�%��^�Ǽ���M�f<� ��G�K��b�z�sM���J5�B�ʸFYs�x7�7�,��Voe�
7�3��Pȳ�^�VN�/��D�/�B-���%-�M��bLL㮝�Π��َ��)f�;o��p�3pn�ǷƩ�{�'�HB�غQ��� ^�ʩ6	^o���
�
�}^սg�{����d�/r&�k���v18��boL�� ��N<v����J�fEK���{eF���ah2�}�����\	��A5i�(�>��0�C�<,�ܻ25�B�P�g�
�h���_�㫞��>V�0���,�֙���؝��uM����qQ{�n����}��|��cY�˞�oe�+j��I�X�����wh��Լfj�������}t����r�2ߍ�FVƌ7ЧI�5|���/�'�o#x������tyP�h�^'����=R*�c�v������b	�~�/k�cǭ'���1B���`��ܶ&c����5�f�%Z���⊚].�᳘{�dJ��XMG���LeX�;v��]4fP�<ZRŝc�= �=mMh
��<��uo4F�,�Y�-E�<z��
鳮�[�tM���
�՜7��L�wm8��n����D��s(^9C7��RGk����3�ھ�x����������W�|N�mhi��}��U<���S:���2����i�U�* O��q!��Os5,��$�BPn��^Ze�S[C��;��>�ˋ�B��f��W��ˢ�h�>o�̝��̈'����>��S1�L��ZM=��Vx~����8t��6�wD����?HP����:���P�գ�"�f���dG�C�����*��O�\ڟy�3=X���}��1�e�H���G���3�=ٓ2�E��允�:�<�Iհ�������s��w�yp4���k���U�f��@�����k���^����R�n�L�w��U��:)ױ�.�C���OԴz��t<!~�f�=���\�C�f��^\2S+��W�]�.ߙ��Q��`߫Y�S��C��a�-v��W�ysxHf7�v�秡�M��(�Hs:�A����j7P�Z
��6���(ƽ~Bt�?6�(223by�6�#so0Ba�gy����1e�����b�M�F���P�p+1H�b�ϰh���K�\�^Ïju+na���Q1�	ql�<��m�Q�d�_�w�ʹŝ8�nk�y��q���V&F�Hb��^��=�:�-��f�4��{��q��x�ZJ�B�¥��m��+v�x�c�䡄����Ҡ�c[0��l�j�^wX ��'^���;���}�5�q�sn�)���
/vb�+j�27+�q��s{�cH��D��������J����W+��*��[��DA��}+��u�w��C�4�x;qwN��Ã @�޶jEL����Ks)Q��i��o�w�z��L£%d17Q�@�<�c�]R�֊=۵�-]t��[��$�R��U���khH���r�t��Ƅ����JSo�PY�X�43��ڱ�1r�c	i�]�<s2˥F����h�q�k�t3[l�ĹY�Z9n��zVEe�v�
����W��X����=%�*�!F�}Y�2-�p����%tU�x_���d^�sI�X�NW�:p�j�|�6AU�f�A��g��rD$��M��Fu��1f��*�=I�l՛"(�rͭ�:���C�cĜ�}�5Ոh��јF1G"�i�q \��8�]]��1mf�%��Bk[�f��t���3 ei�'���"�\�]�z2ys��Ȗ��|�[%\_�UgR���c+5Q�������;���ƕ8}�e��P�s��b��iצ+}�IUl'ب��)����*Bt�|*ڭ9aʁ�	Ǐ+HHAw�qb��za�l+)���Jł<߲��3K���mJ2���E�V��*�v�w���j�Yǻ�w2���CGRg�eq!�/GՖ����X�:��c�YAHWz]�\��y�����Rj�
[C7���_�#M<��r�Q��/i����\s�U��Y����+7����5	eY�sMO{��)I<���V�ٌ�Ry�RQf:W��ȹ|�+�ո֜�Es��$u�M�f�M�.�phI(v*زZGv :p�o����NI^��U$��t{p��HI�X;'Vp�3�'ҷ�bw��v^f+���R]�`��7+i_Ph]��-|�n�Ą���*�������h�q�V�fu��ʶ�w��= �~f��|%i- 3�eڈ��=�e�w�l^��+	�z���o �X���H��=�m�ͷ"3�}���c��@쩘�Ee��Z�G����d6�*W��,dy`�T�r)�AZ�!����z�o���e���<]�fwc�}g��꽃�4�������ӈ괬�f4SN�1asq�ѻpN.D�-������ǂ�y})�)1]C�l� "��|:��;N�uw�4������|+(5�,Dm.��d��+���2�X�	e�㲬.��Y3se�U��(.�n��C�;H�g���h<�f�*o"̜ЏAn��l1�9Q9Bvtg�ɸ܇�V�<\�j�mԚFȺ��w�K���.}���ػ8n9`��'H�s���w�_m�(J���wn�sJ\�{��S�5z���v`
����=���8I��Y/�n��hG�͹���T��'5�*����iLX�����S��s��պ�t��-s�Y~�I_$M��[����
���O�����]t���ې�I<8�5N����of���H
 ���0R��Q6��ؿN�j���#P�����k���nNH�Σ�:oU����g{��f}(�L��n�/��Yu}*c"��w�K���6]NG�3ƚR9h�4���u��ً����8��q7˫0)��E��<��`_�:%BUalv�[d\��ދY�{l�90&�0��dAN�&g�A�O��b�x�J*�ooE�	�Bg�������@v�
��(�5C���U%�U�R(�Ϲ,:<���n���9�����i�6.�^�ߋ}����G]��0|{1�˩�w��V!������c~G��&���T��3��$�<ߣ�ǙFЉ�zyM\�n�r�U����a�̗jz6��k�;�P�U�����&�I�����®3+�r��+�r�u�YF4jU�}���H��F�md`�&%��\�8Q���٣�Oߠ}������ˤ���%YZrZ�b/���8���X跎J;N�m�k�^Uj���D�	B\��;�P�o��\*\�f!/�t���
ȀQ�#3�{3S���pm�}�+w>�Z{�	��4�CѺ��R�E��3	�r�7�^�GEr���ƺ�)`���ټ�-��v�!��G*{�M$��ϗTb�F]�o!���M���9��e�3	�@������/8�}۹H%w��P���^9�n�c�k[�5�����bK9R�2�f֐ϯ!�ARu�Phʧ�u����.r3�i��Ѓ0@�d��Ƨ��������1$NË��]�>�F�^̣<=�8����L����T��d��Vb�Qw���ݙ^]ڞ?e�ц�������C��o�g��F�2�v^�7�S����9\�G�z�c��TX��-��&�k�FT��:	G���|�����F,��ޏ��Ч6�@�UFȉ��p�+Զ���s"Q���/������n�w�\q�1tDp��.�����!n��Yx�H���"��:��Eo\�b�1�\��rl]rb̸�"�`D�.ђ��W7f3n�l�yV)���rT�U禵՚�f�\ek�Doo]��U]G����r��Qq�7~9J֓t
G�7kAp{*�9G�Vz�r�Y}G�z��sw8��a�of=���<}�mU��l�^g0����*�&�>�ebcfB���
�q}�]׎��8�����d��}B97���.�y�G���f�PYX�ݥ��Y����u��5F�~�5鬈+(��K޻��̱�tf��Mg�q�I"�
���`����оH��ּ	���D<��[��\9h�s��Z7��bΎ�)��+j
|�կ�����wU���ҷ6������aS���wǅ�Hd�(�8�;C���t=�k��*��_�"��p�M�:1R��W7}j�J����^����'ݔ���28���#l��pozu^�#}��u��~����+|q�I~��G%Z�E�ރ����g��l^wӺV���7aN�����<�2����Gw�=VtW�Üs�wm�!?91����H0Rv�32��jpR�zk���D<��z�	�+T<W��3��q�~����n/$u䉟�.�Z����~��,�O��ד��i��1�`<��]���B�_�B�p٘�w��M�9_�
�Ozv��e�ֺ#�z�_�J���w�'z1�s��ґ��oKWvM�[����t�O-���}�$x�j�nO�Ww���$C'�9�N�������?+�?i�ew�>Ӟ���4ؽ�w(�N;A��U�C�m�W'W^��>�'�� �L�����,M��ᢢ�q&��FRj���W���z��2�߽��҆�:~��Q6\�p�R]+F�ۼ�9���3�P�c���qeu5�yE�G�JC]��5.�F�ෳa���kJ�P�h��v��j�QWvX�#-���9Y����� �{q���|x�؂�n����7@8y�Y�K&���[���.n�vI�sO�2؞��]���Z����q^��~}��/�$�#L�G� `�#;ٹ�o���6�N��K�)�7�&� gi�0�Z��VtM��il�&&wǦ�N�1�9F��칍��J�� ��J"�jY>�ݴ%G��8��k�Ӿ�e>�Kz�x�ԭ�=g]�E������B�S�`��2�����<L��=ҋ��� J,K�a�༖ڦ�ݘk����O�N��{���L��(͊2�I������=Щ���3~'N�19G{FZC[��Fc�U��d !����ѮfFK�)�)w)E}�NZf#�FG�w�F�u�"����8�^�D�T1ϴO����W�0�yC�Ow���������}xZ�-D�Ȯp>d${VY��e_nW���z�pLw��/،��zxW�_o[���z�����=�Nڴ�g�C�k�D��Ù2��ɂc�v��=7�m�5�І:���Yg�`=�ӣ,a���盿��J��[\�y5TCѱ埓���y�}����3]x�p�;�u��U�����u��ߤ}_��pˡ��֣��@)�����wz��<�9�Y�E���jĂ�M��[C�`�y,iY���m���b���4:|���z��j�hWeh�e�*��̽����؎:�<K�傘��vq$M���{r�	�j)�Vx�F�P9�v�O3���2��L���Ev-��n�7?U�<t����K�`>�(��0,^��VO/p�Zq�QWq�f���p%gMd��Y#UC^�p�Z��D��_���E*��X�Yb<����yWW�= ���1T"S�X����OF�=YY�bҎ�`����_�mx?\@4fiq��w�-��x�Suw���n���f%��R���8/��� �Ɖ�.g~�w���p����:�SV���fL�3[�D�pd�o!*ѓ��+�w��ۂ���u���1���uw@�>ٰ{�ui���*"ӑ3�T����"�_��g/����Z=�Q�cj�u��ɰ��U�	�	ށ{�s����P7��"Yާ�5��Z#c��d_�.3Ў�U�����06:���v���;բNFn�Ċ����x�h��{��я;]g���n��x�~�J�˼�����}J={�v�H+��=�ʂ���Dul�|�@�uU<����Y4��E�����r��za�UolU:X�ŝ;C�<�vō��1F>����0l�yOe{#���zEM
O����׽�Q������5��(��u��v� \&v����ڠ���	�l��3�8us�𫈍���M<��cm�MD<b�g+�0å�k�xT8Z�C8fAJín<�-�*�º�&��P�G:И���Vš�0����%F.-�~pzL���y")�Q3��w6�U{Q��0�?11:|��fÖm�2�9�b�F*P�|���+2:��H�'�v�Np�F��E-���r��\�_J��ĺ�\�ʹ`��;�Ī�9�5%)��~�-ĥ�TL��ԫ����ו9� ��=����-���g�w}v�`����G=U���t`�W�/��3�q�xnB���7/G�zb;>��;9}�B��n����\���r���g�����t����ѨF�G�snt���6T���� uHǳ��{�@돦l �<�=�~s�_z����s_�u�v����󛓗��yA �7��䲱_e׷,[=���!'��re�Fg���tҪ
ց6�uT������{�Ƿ���CG�FLa}����Ȉ[�^�E���c�I�Ǡ;�c��5Ғ)婤:�H/����X��[�	@H��֥�T
�
�uo�Dq�j�L������u��.�u�#Vy��nyU�:cy��yZ�%��fD����1V*���O<˨&2�tflf`i���A�}�b&�<2?���Ou���iƍ|^=��F-L�;��q-�/��'���9����A`GY�p��V�+���Ts'CΤ�]��~�u��Ça��ի<t��+B�rVV��;��=���9�d0+���aC)5���+-V[��z���z����������2l煼��nP�����{���:��Cx������~{׎'� n�k�>�D";=	Sf��u��r>�vsZ��涰�,^�#��f�TYɀ(��x���o�7�2r��f���|��@G���`f��ɼ*e��,�:��I������Q~���{{g;�m�n�Z�S�}f��a���j*�h�3u��8�N�޹`��b������˺�;�wrz��\;�5��#���{�2U省]N�^S1�l�m�l\��hk��p9�Xnm%^����$y�o|�>
���������Ŵk�W����y�KW�~��Ń~,�q䯖�E"`�׷�x�dn�G+�L2�3 Fk���ͤN
���y!ܲ��4湾�oAI�z5���;ث�[=�f�^�"��Uj�+*�`�L���u2��Qw���il�Dz��M|�	3����މD�WWSs�����>���xW���+�Ƃ޿�A��Kˤ�mE �m=�t#/�]����3|)2�����b��~K�GyP�ok]�w�JK�l�N�H�55e��c�]e���f.��S:�o�(�_ZI.3�=*���܁U�v/h5�4rUb�R�\��S@�
�6�Un��a
	�����j�uվg�-7�Fs��@�b-�n֣a!dӄ\�nuD�e^x-�xu��6Sjb�f��$㏎�b�������/j��s3����,���7=��1ȵʶ+���Xv�\���J7"t��S��#H�~�?Yq���=λθߢ`�Dm��g6�N\^�޷���-O���O��s���WDR'���&&J���b��L�ޓ�6�C���o	/S�vq�C/�*��3�����k�%�a��w�Ңn�0�O�߆�rh���&H̏qK�}^�ᙡ5`v��ܯ5x��CLr&��8I�eyyr��fMg��V��+���έ��	}Hf�쨞ݘ�f4����y��ZYz.P��N �>;���W�%�P���}�]��/�;�d╛bsn�Ч��t�����9[^����^�����m�kr{s��TLi�[���el������Eȃ�܃��EG(�̛됫]y{<l����y*DK�n���=]C��e���qn+�'�NϹP>�/�!�Kgu��pˇ��%J"����x%(x]n�ۭ�x;�@�{Qz�I�T}5�%v�"WZ+B7��s��a���}�?�����^wi=WH��t]�,u�:�Մő��+w�����l.ވ�H��:	�יIZ���1�}cK���:��լ��ج�-?dS4��l4�N�ጲ���ҧ��ە-�����W�cȖ'�m��xr�}�XE������;g�y���c�^`��O�n����U�xp|�=f��^K�Pw�@n5)��d��s�&��/�<����R�o�WY��2�KM�[��S��:ZW��ts�����3���J����ݬ���g�\�@�3g�1�����~1z?#	EG
�LG{���~�XmV�t��3��7Ȩ�&�_ED��c���Ko!вu��q�"��Mh�?`�'+r#65�+H����v�I������+���ybQ.�:=	E{q����q�`>9�ŝ�"�"�����(��w,yI�>HV��WZ�=Ϡ���RT)!V�������2Y�U�a}q��Vb���i)w�Ԧ\!f}	z4���.�9F֣�&�>.��T�ň	��۩�L>Kü�3Ĳa��b����A�
\��*M+�����b"�>��W�g�<g�&~���r��R��TZ�L��5%y�pZ�Ii�M��H�Ӝ�q$�<�T\�q����v#�M���ԃԿ~�&R�]Hd��Cm�ڈ�8�z���O\@��*�� >U�=���\2�zy�C�͌��<5��m�l��w�ll�\)@��B�n�ir[��+�<�ځ�p��1fV��� ��w���q�C�t_1�C��j�w�����[��T �� ,"/]_t�����/h��0-zWw<�`���g�g%8��nD)V#w�;rⱻ�~�YQ��(�/7��;'C���PDC��&�W�L���(>h�[�	��y��[�6���DY�U���}���ޛ��̞�,��c�qi_���_����� ���TNe�W'�����[���ۓ�ob��~�����T�K���uh��rp)�H�!�����oʜ����<�IU+$]���,~~�J�x�~D����8��y���i�31\�Y>x���=����F�K��Ժr��3
ϡdD�'��;�s�=S|��߈��f�ԩ-d'��c�5E)d��ֶ�!�o�)f�U����b�cv�V*�7��uLI2�R�28�V{\�-��7��3P��}�k����n���_�Ю+���^�x��/D]u�5l��9ޅ��{�����چ��s�}���ۃN��"Wx{5���ӑ��p����pV����.�ʢv,߻I�*n���m�%� ��NP���Tq�9	,�lR�z����r�<U~�0���0敟��ͦ��ȯ�O�>Ӗ�~/`q	�>�d�Y}R;b+N���X�.U��w��%L��K��A�W���b��.��c�@&�����Xޚu!�c.m����ǠZ�#�(�� Htu��Gk�8rʂ��ꗗ%. C{�eYq�B��\��X�Ι�4�X��Id��஡ o,�H��]�|%}NPe��l�kS@�'y�/s��.���!�uCi��:�z�Mc�t���$o�Dk�յJը�9��\�	�o���yF��n�rH�Xņ-p7�	�Ӥ�m��6#�](��Q
�wj���P��NS�v�N������������L��J��r�x*�Y��'�;�2Q�(�Q�h]nwQ�L��9��ӻ#�#�<�WJ�c\[�y|Vq��;�w@��0V��p��W;���,�e��w ��%��[��>��Z&�؈��p��T� �K4\ :Fk+ n����M�#w��x�����G�L�����R�p�Jf�\��bYE����a��Y�#�&�����tve㽿9\ Q����k�#LEǻ���:P�~|�����w՝[\1��xsK��'��%]�9.�n�UjxZ�1�V_�%WJ5°a�M�q[��iS��ޠ�e�R��[�B򒙵}M�n_T��e�065,,�]]�0�,���>hJT�݆J+NS�@]�cq�qS���WM����a�����e�7,1j�J�]*��f��sX��a�:�Մf��-n)́km���{�AvW��-G�,s(0>�]B���bmVe�5�t�ʵ:L�d4Y�Z����$V0R6V�;�5M�2g.*=��}Wzc�]Snmi��usxwj#�����hS+�f[��xx*���5:�G�4��b�$}��ൡ�T������:Yg&t��p�qw�v. *O�,I���ԯ�k1Y�����
�u�F��rt�i��!�7N� bd�Y��b� !�Pi|Y��ٹ�B]� ��s�N���N�v�W�,�1݂�����[�:P�5Z�0F�zƜ�V��;QP6y���6�9ި�5�V����ʘ(MZ�V� �v��}K�6��>Y�L)��g��*��0Ą��8��;Wa�����˩I5;�u�7 ��2�b� 
'����|��y��]f��+v<�i_σ��>FM��f=�!�q���B�mzRÂS������lmb��=���E�=�y�+��#w;kb�Y��siZ:�Ag�c������4���g���b4i��ӈ�n ��5��qTs7�:�2�ټÅ�v��*mM}�ٝ���&h8�z��h/'R�1�7!f,����-T�Ё�;�(�kY��ȕ���ԀvG4_�۸+:dv8��J��]LM�b7�b�jV����b�.q��5�Em.}�"�9�,��ʊ�6X�&ëo�F5��uIz�d���\:$uq�#��z���aM��+[�$�t�-���4u3�b>q���jcd8��!nb�t"k��&�*v>�:���dc�S�G�NĤIŴ�'Jن�gL^;�+ކ�n���z��\W=³���/�{h�M�+�$1Y��+iU�v\�"|q0rw~�b�։3�Z��ml�c�ds\��"v�+L���x���w���=	���%3�%s�9唆۞�!�k�}�==���X�/?X��/4��;
y"C����ӯnb']y�$��۰�8=���b|�Jn�v��SA�������Wwb�w������*r�8��m�W�޵X#:0֦p�PY�DF���އq3(ckh��)Q��[VIv�����~i�x�w��v������ʶ�HƜǲA�����5���`�ֺ��ң�.����SrFX�o�hw�j�i�J,FE�Vv޻��n0k"6�鈻<�<<�Lgl�]O�k����GJʑb�~��d}+�=-�f�����Բ~�~&4��t��8z�u%v�V^�:���W��Q�i�>w��>�ڬ�n��z�m��k�.���:i���g4dp�������I��=����@�ѽ��ͭ��Mb��U������Ķ��˳VQ����9�h���;[E�z+b���z����*�H{��t�:����I�s�@�䰁Ʀ�bp׉��󳱵�j�����'Lj��'hQ�5��b;���2*��b��TX�X)@/-*G"[��P��8,)H�u-��i��(�r��rvbҸ���7/�K�Vvo������ƪ�@�1=�yy�1��4�>�ǎ�n�l8]��e�g�>����=wY���d3�h�U��Mg�Yײ��"*h���m�8<(]��bՔ�Lz��ۄN�ܷ�������.�5ݯ0=�-�y|��G��q��(������"3B��3��D:��#���d������V��v��^��p}�넽�Ӗ'bhW��.����l%�.�Y?e��a6�~.���h��7�%��Ө�b���VX+�%��{nt�D�6�8/ܵ��oꮘ >���H�7J�pi�F81�WyQ!!w�Nz�����!��a�8�n�z�dԺ�2s�ݸ����Gd�����+A��W��5��j����>�W�t�p���w_���d�[(��{��$�� DӋtF��VEa�����x���W�v��tN����Mku�����zؾ5���\��CR�qo�7��.��C�����V�y����:��t��Ǖ�AX�Q�BƼ�6.�:�]�t�-�ĝ��ρ�y��63�:�9�\�����΍�LRy�;��������9yۗ�>��'Yw'�t-S�n��q_M�C_G����������;�N*��b��_�_ogn�5T�ƕ(�<n�����Veu@�YɽLmŸ+b���(n;�.&	�ׁ*�y9�h�-�s�����Wv\���%�Ph�@e�1�&�ֳ	��u��k�gLa��A���"�-�r��9�1�.�%��hUEۼ���f��܁��Π�J�8@F(h'Y���չ7��X*~��i���0x�?�|�b��{�
Z�����G��;�q$�qk�O�U��|��3�᢮�L!�q�'�T�4g��C�V��xҤ��3�Sf��?I�	�Z7�;~~���<}y�j��^�[��y��AΕ�Z�T���6�U���g#mr^�f(�SHT���J��,~����` )�9w)�҂�5�̜ܥ�.T����n�)˵?Q��b�5���ͽ ��g&��ݎ�>N����7�z�署��23�e6�u�^�p�j4 ���VEW�ڈc=Q�:�)������uNT�eȳXg_o�My���V���29��ח�v�1�E��hM��{:/fv��/6�KYR9_zEtO���ǋ�V��W����g=qG�͜�F�y~�.Ɯ�k�yU�@y��gr�̲�a~=�D{�ܜ�P�:h��*���Rwҽ�d��Qı3Pv���Y����솺��YJ�#� a��*��N�Q�i*Ԯ^�۫0>�y�N��aqw.T�I4�.�\ä2�İ��,h*�C0ᛯsp�e|�+���P�ϵk����c&!6�ʖ�QJ��5�X�wt�?M�7(��+Tq��ꎭ�[H�R�s6���hq��j.@.4���َq��~���흥�u�O�Q}驰�w��zca��7�9��7EsV	=�d�yMx�]�ϊ�J�!Q֔�nԳ�mЪ�Fy{��QGgF�Ez�������!c�d�t�Sgګ �JY��cw�o�LO�I`�F_�����4j��<�*�Tȵ{:3FTH'�C�r�υ�D���<(�*� �"}�}u�v�Bϯ�r�%��c���Z�o�V���'�CwS����,���#�*y���S|Z�:�!ݬ ���(���e�6�,��w^����w-y�˙�)�&'Q�@{w.1��xq�$Y��%�ӛ`�j���Q-^���;�r��㮎S��I�bN3�
�N��.��R}̧-�*��m���讙�^q��5�Eb��ڪ�������=:�9uMu(ؗ�T��S�~p澍�WI��p���sKk���O��&� �W��(�A�Q������;b��55;�S��ˑ���C���3,��a~��f^���w��qUs��1(�0�\ K��/�Hm���O[��xi�n�q'p�u������f9��S�ВƔ�YS2��H:�Xֱ  �Z�R�y\����=ζ��x�Z(�AG�M�=�3���k�9��D�빼��wV-}֎qҏgNA����S�k3腓O\�*f�B�lrE�{���Ä�{M���*�yl!���q^������I�RF0"���S�3YN�<�u��k�v]�Rz�v�Qqb�Xҋ��sV��<MN+��5�����Q���}	V���<�*W�zw�:-g�W�K܌V���]��Dx�}x��.����X�F�UD�,�m9��5͗z+���"��B5��{�ꌾ�\�(��W����[�[��3�����f�
��<�?�5��cS<3�(��K-ɡ��j���,vs��S H�����G���<lF���f�n�-�q�,�.`���J��T��=�US�٣���EOn��(������k�x�;"�/:����EuG���뀧��C�S�Gg�O»�h���^�G����~}lS��./Wd���:DV���v�0c����U�;�x^��L�4��}�H��^Ӹ�\��r61�Zt4�ww�屻o��%#t܋=�+ue�4G�����ȋ��}��[�!�S��x���ʍȅ���E{��Uu
��E��ӧ��H2���/۝���3)d�e8�J�`sۭy���]g`�KSv-�|-�
u�xʰ�)0rȞ+���i�{{��E�.�\������L�ˋv�V7�]��X��ΒJ�,�8�qZ�k�h�%`��ժ�֋!ۭ��}ٱX���i����F�9����J6�Qv�w.uy�eq��J�l��hT���2���U�fC0�y0�ҋ���O���a,�눲�l�pt�>�S�A�u����w<Z���œ��]t7��C��~��?�|�a�����ȧ�x��e��u��ξ�sVv��]}}c7�Y��4�9E�ߺ�:�~^}(DI���VY\J5�נ��g�Щ^Wgsv>���3���s�#�gIBN�Ei���֪?x����Q��u��=���b����M�����-
z�C}Ie�Ce[�bɮ��w2B�C���p�>6���8�<���}.�U��g����Q}��*ݏ�Dx,��RJ�[�޳7L��k�Έn$F{cF�м\\egX�ɍ��j+��¡������;�f՚��*b� $)��R8��L��u�{�(C;|��xN��&X�Ju�L���5>4o�~�;�~v�<��	=s7ӓ���O�]��%��b�1���f{�RQå��{Exp3$߻�e��1'ѝ�O�ŷl[7�m�Uԝ��6*i����"nΧa���t�=�۹zz�/�(J\8s�!��F�v����N��u�ŕ%%Bff4XI��ut����ɖ �����sQ�}����;��O��߷���)c��'gic3��t�xc���S�՚n,X�k�W�&�^rt"�׽v���9ėqCƥe����iJ��[��ݏ�pn������z9�!Wܡ�㪠_>�+�6=q�*r���7��^�z�s�W=��JL�^j0���Hg:�D���ё�����	=�U�"�5��� ��Qt-/;��v�aZ��c7^nu�N�׉��R�D3	@j�T�eWV�R�*�^���xUz����K�f�s1��H*r*A�Z�����3�.�.}��S3)Ó��݂f�����8�%z�Vʸ�+�{uC����y}ºL��x���a/ؚ�n>j��fw�E��͐^٫~��&��MJ�Ӈo��p��w���A��b<����V��SP�!�=�1H�Db���8υL�o��t�ԓ[�kF�p2No�4Dj�Tˉ��x���7D3lط��_b���۞@�ۨ+�
���rb�W힕�~��/�8V�/'\4��մ#&uP�#c�Z�W��z·�_�L���Tlu���	Rx�Z����׊��{랍 1��m��O�/*�x�^lߕ`�zf���x ����CR�������;/J���(�+�]��f�&[�c/��Һ/y���t�f�jՔg2����X��������c�����X�ԗn�۴���36�{�%|1J�X�\�o��J����X�8j铲����L��}�*�}3;���{��&x_���hǠ`+�����pj�u\�?O
��
u+���udHuPE7:+9�<o;�L/�זo+��9�N�v礕��@G�6��[����y����g*ӂNlb&�K���>�ظ�[�/�.��8,χx�F�J�1^�7�<�����Y�\P5�֞yX*y��MＥ�/�]Ý��HU@?,}�P�ʸ�,���44u�a�����JzF�!�=���ѢjjX�����w8Ƿ;ga�_V���y�m����+�ܾcI�6�aޤ�F���H��i����E�eO/�s ^������~y�@�^�SΣ.k;+�3[�����jS	���N���� o���rB�p+��%h�̦��L�Mo�ƻ��J�b����7Nkѫ`9v=��{��bx67�	�F�4���o�U��z�M_����r�e������]_���btɽ�_�$8ǿ(���y�3���_��G! ���k�_���u�To�m7���2W��.��#ni�r���,_���^��!���b����9ǟ���y'�Q����dh���B��kgusxo#�j�Ea���v���]��a=@s�ޘU�����C{��o�5������wZ%ͩ���c�Q��<�{O1�fI;VW
]Pq�z�>���բ5�fuq��4%RUjv]�L�+���,��Wu�ŅȋW�ofi�r��1��c�ux���F��2m�U�՞�u�#�$uwv�Uڻ/��[�'!�g�	�Rh���%�~�_��}��:���v+�h��vv�&)���~Jg�sj�D�&�����e�ߎ�lm��Y���!t���{���k:��
G����mF6e��*̓�k{��Q�xx�3�s,f����By�����==��Y�q�"��CL�nO�bb����Lc�l�I��:ja�FX�dG�΅��������v��
�,\�E�U�i�W��GI_]�^���#�ڨD��]2�7y>8��(�n���7�ӣA�s�d�8��R}��t���z��<�w��f,�S���D�&�K�m6&Aa���6ĳ��=5�F1 l'L���èU����h+6(��b�'��-dQ�f9�xvAJ��7�ݗ��$��E��<�v��Y6�����5�.��v@���b6���p>�&u�&��s�I�8Д[�����'�1�Β�|�p�V�G���{~���zwV(ﾫ���s5�EU��� �,ŧ+�k����v.�ގZ�ݥWٕ0i�)���jj���ǝӵZSf
�&�;��:zʮ�n���.�vv9��*W7�ݎ���ò!w�N����M��V�M7�E�5H��m�t����5��t>,t����#=� 0-R{s���.^�)�Ǽ!�F1�����ہ�g7��#+�v^�!���	��]׻��y#]��d��œ�b{B���&�����h�{"������ٙ3޵�B�hu����nEy�"1*�#�����Е���;-#w�Ǉ�$��ev��ҭ$�C/��Ż^���lr���wd�s*<&ǧz���b�d2)2z���W��7}x���2�3�"�]gb��Ն�t�k���_�5?,���3�#7w����?)X��dO���z�on���Xq�W�%MJ��_��G�M��V�t8�b�_VGU��FC�^+k݊z���c�y7�/zuTxu�3����1�ƣ�
�='��3ӔQ�5W=[]!;2r�^�#7w�A�iNM�מ��V����� kꛝ�}U��1�2N����ۼ:!OEؒ(Mb�?�yH���WG3 �jV/�wۺ٭��f�=���?}�}W���9Bj��΋۸���.�s7��72����k�?)@���*ZQ:��h����]vȏ՞����5o�ɇ:{4�V=2��]JyZ�s�+R����!����j���x�>pv0�]7S�^Ҏ,�թ6{���%;�u�A���P0�B���2�R���,E��Κ��6"���$�HO���HI�$$�$��		$	'��HJHI I?�!$�$�јfff��a����}|K�����g�T�ςY1�JV��.��G�Ai6	����V)I�R�*ȩ�.�h���Z�T�ƥk�ѭ�,�s�r$��OM�LٷV<w���s �cB��h�����fGR�.����bƕ^|���l�-u�`;�Y6��.�1��+Fǟ�>#U����(�6>SY"�5*��Y��S���U��au�
uE�A
���G�1b�/L��B˛N���Wn q=7Z2��kq�ɏU���C����#��eƬ��*�J���f��ٛ8�m�O&�:
��)��c�g5�t&��̢4���3\�JTa��q6��:p$T�[�m���n��x�Z�����U��˩i^��,8v�%�AX��Dhǔ���˖����&�;Y����*<o0\�6��9�J2�81J
�뤳�4�Ytƻږ��T��dAQt�c��8� CG �gq;��5Lԣ(�ʸ��Uำ,��z� YБB�Q��W7\զ���^�@md��Yt�Vf�(!Y�*�N4�.���u�����A���p"u-7�n��$�&�gS:X(�z�s@V)�K��/j��˥x���!Ű N�TD�5ɐ�g^PpUޜ�b�YÆ;x�n_�.�Vn��m��cn�:�����%�
��R��*�m+)ku! ��ڻE ���.l&��J�x���X�jR&�j�@V��ͬ�����̪ ����ɒ���[pK0Š�ܨ۴%0u�nޅv
��Q֪����X� �c�@�5p�B	6C��uP�*(1�Չ�bTO1fSx��֨���LIVP��ۗ�-�Fk��#2C�VTu�i�G3#�>q �Ք��Vc���DQ�$wv���Na��
w�K����Ͷ2�K�{hZ�ӧM�q�֪�^�2@߬F Yb%m��mdA�[�M�r��!���ɱ�}��h�0ۭx���H�E!�H�Z�H�H����
�Z �LU\�E���%�k��4����ʫ7VW����3��333�! 2��$� �� �`$�$�H$�$ ��0$�BH� 	'�HO�$$�$��HI I?�!$�$������!$�$��BII�䄒���	$	'��HO�$$�$�̐�@�t��@���
�2��^��D�� ���9 ��>����窰4�(T�!@�E��,ih�kZ��^��*��(UB�US5U��e*�-EJ�%Y!&Lĳ+Z��͚@�EB�R� P	��%U:�H����@�5*�%B��TEAEUR�AEAIR�J�EI����    ��rR�P;`s���\��v�J��ו�5�ït�$�����{=�{�u��Z�u���ol�r��]�8s�
���(�IDRq��[6Yۺ ,gp�I�\���5�'nwhkYF���K�u#���h�۸5Շqֵ��fp\r+cE�;�t�iF�%*���WNEk,�%ۮ���gqwm�Zv��\wwp�V��P�n��@�ɻ�r�!��m˝˸��î���%a��'M��e$ʕ$�QJ"㡈�r�MV��N��
���\w@6#��]h�\�W��1[+Z��y�P\�[�j���:i�@IU!\:�iI�sGZR�a���p(H��;w�c4�����f�E�]����ven�die���iA�jJUR�q�9�蠪us�h�N�úq��t����&��@��p�QJ0�`����� ���X $�RR@�qҋ�����6��!��@knծQJ�k�:�9(����Qc��l��kKU��v��`J�a)T� v�6�]�wM�4s��ki�Ytu���譛n�nm���:tu]�u��k���43�Z�iu�Q%*��jUm�H�n	ΣA]�rJa�eA��
$;���S\8�5s��(,)Tq�;[Megf� hR�E8���l�q�l�R�7m��n�\��뚡'�V��K�;���8&g7:��Z��$8�S��J� @ "mJIU�� a�� dbL�`����J�C ` "�CM(AO(mG�z����I���(�h�%p��o�f����$����F��y�*b���:���g�"������;�@E^�@V��TI��$ ��bI ��|� BI?�Y��_��.��y\�\��֝���;��2��&޺��:Z��4�+2����4��-�#O*�X�j���F�q�A����J�{��P�5=�z�*�&5u3������l�W3��I�u��:]�,�k�ѶF�j��.��Se���͸����Qn���`�Rܚ} ږ�� �	���P��M��lP�!���$7�b>R��,|h��Rm��!��`m!�a�)9`s+��ɫ(`.�Hx��C�!P��0�C9@�i�M�4��AHc!Ă��o���X²!�T���Lg�2i�	�$�Cl�q��~���/��YHT�`m!��RHg����=Hx�m!�Hq!�}�7|��<�[��;�S���y�iSL
2��)f��7�H�N���6Ú��^M	;VL{�hI�,�������<��*i8E�B0�����y�E��W#�����l�H��	3�
�n��]����ªb���hB^[D,y2�h�<�t�+�)'yHʳme;�wjn6Ym�H�H-: �Z�yh���S�2��,�F���S5�*��+6ܩn����R�)�C�{�m�ܣ�RM����ǃw��U�1�1���:�H[å�޻�y�2���-��vj�
��!TfĤ�ش9K��6/`��IAI��X�Q]��wB")�*��&�JV$7o7���L��xP4��������*�f� ������qSфa�c���J�*�ՊXfkm��[C�CO�e%d�v��Ր��Y�qQ�(b��pUܺ�����dt��xZ�V���X��NZɌ[
�����F��Z�hn9����I�M4���P�3V� ��)V�Z���m���L 7S�h�*4&M8N�c�V����q?�������8��+E�ƛ����
'E4�X���+��XVi���`�!�֫L���Q�fVB�P� ��9)�d*��	��m���䙦��C/i���i[��F��V����{S+��鉨�JVh!u�����0��hHF�V�V��ƽs"P̌@1&wq7�M�(�2����ֻp)PVl:E�y���6�ht���OD�-
.�ժ̐����A���X%n �Ɂ�Z1�{YR�e`g	��2mMǼ�Ή-�h��Z��0n�jjB��{�(���Tu�
t�uf95ڤ�L���f^SZ7?Z1�Ci�+P���x��ۥ3X�t^��i`nͦ�tsh��Z�	�xB�E7N��St�Y��͠[yf�S�`4��a�3H�""h�T 6ΌH]n]�k+T80�6�^�XQ�[�[A�.ѹ3H�k5�T��OIx�J6�ާ��E7%�+Em�:�!��ҭ4b-�wl��M �0l�	�$��I�nbͲ�Y�ۢ�$�d�T��WE3��)z�|!a�m��dd��y����]:l�r��K��{<�e]:��40���"付��sDv»yĂ-iESK
ӻ��P&�:n��a�, 0��u��V��l	�IH]�^�KE̊�e�5-)��-�yfɺ�W$�*���O/Ԯ]R�Tkh64�����r]�"
:sj���Jނr�^��L^�h���yD��J�쳢�iR،08&qT�̃2H��@��F��yf�!��YI���������Z"g]��\�u*�zf�2�T�����U=x�Z�p��N���]f��7�f�\/^+���ÓX
���|Dt�c�8�S���v��Q�u6�m�׎����;8�$���|f�_5qi�rɩ�3:f֔��s9���˼�yM����,�F�z�K�ȳ�Z���mm,�����U��jҋ)���^�bʗ`��mJܻ�@��N�,P�CS.��y��ɻ���rIy��-�1!�] b���M*�*keL��pLr�3Z������o!Te��7�S`�Z%~_�(4i���K�n���Kc��j��b�TG՗-]z8����E�o�3^S}h�� �11�y�Yi���q�]#�X�9��Gv^��w���L�ȭi�2쵲�b�m� D~�3#rh-&�Q�<7��:j�o�o�p�-ׅ֨�h���]�z�[.k5<�ej"�L��&�	;�U,P�-M��JI:s41�cT%��� �V�8N%y����s1����c���,�N�L
f�P��Zv�hY�mQ"L� V*�&��"���⥺X"�PmYHm� ۆ��r�J-*��ƮHt׮�C��@nG�i��H�{��j�ZU���ީ��.�Ȣ3Xj�;��M;���UHmӪ�Mh�V�\�g�u�ٴ�j�*Z�źJ��T4�[��,ح��(]P=�C�B�ۗnu�(U� D7K�p�7�
��o�;�;���sBK�0POo�6����R�Y�A���#l�V�wJ��ʻ�7Z1���k9��!Ǌ�
81�Ydl��Af諵W9��U(T��1�Щ_�t�RJ;������N�L4�Ȫ����̰Ra��)ZY��頮�:|�ͦ�"�umF��=��ܺ!��1
ZL���KB�diE�I��r��x�,��w��#�8�\z�^,��g.	-Xv�+�����d��IU�x1(�X�dJ�:M-�BD6����ӫ��=��^(���2�{R�j�F^�]0D�@�l�j�2"5Var(4�r	A�f2�!��$B�Po�5�Ĥb��030R
+6��8ň�h�[w����&���	j�0a��u�(ݧ��-���%cCb�M{Wa�b�cÉ���ߔt՚SoɰV
Oc����`PGb��Oe�)�Ԗ�ˢ ^Z]����]�Wk8�;�u�ވk�g:h�w��5�քh̺��.�r���X���$Ct�*�
.Ѻ���ݧch����3)'���@<Ҭ��,V��I���gEY�bwl2EiƞQ��A�L��`ň"Ê�U�lU�x�h~�E�ѱX��=�oV��ֺ����i�r����눢��DX�/(�ۮ�]��m���@S�0#Y�sQT�y(c��6Z6,'^Q���f�5HP%�� l��nR���5yf#u�Z�S�n]��r~+v1������=y1�C/@� 
1Oj~'iPB�c?�mY�Q�� �ñJɡn�fD
��m�wVh��MRӴ��ҫְD&a�����R�!�p ��ccp^��V��v+1-"����b����-�^�����L㘘k.Bq�ܣ�!N�%�C(F�j�F\LX�@�7$��4�r�����%�T���kJ�]M1
��8�9��{�-6��D�`��luf�,��m�,b*P���.��eӘn�� �Q����K�X��p�kaej�6���+I�1��[b\̀j/���B[�*w��yk|���-A����Bj�� �[��!B���K��0ó � �f��<�{a���ՊNV�t�e�)���伆�Zt�GY�H"��MʻH�b��ʺ@m	oR-y�ܤEkt���~����5�Z�����S%�B�-v��V�S;�2d��~��/'�.�1*��2����*��EU v0E����֜��Y�CD�kn�V��-<U�m���:�9�ڥg[l�0�t�(�1Q�z֠�(�֓W��]$soّBIN7x�a̲�˙�Y�5���h�ViZ5����(/C�v3V.Mib�˺���P;t[x�������@	%�]3�,(3&1�6�2��l� ��r��Уy	���,X��[�F^��1P�Lv]1L�r�f���Q@�j�iǊ��,��2e��Ni4��mm7���0��n�
h
�k޸
֢%�	�D]m��%��K��F�o䣧r�G��r�v���d�Z`������K��
�0(X�*�4��<R�4��L���p��܃fi�e(NTWZa�1�a1�Eʷ��^Cv�r��M�4��v�i���_5�ۼF[ۻ�:E9h���D�E{�9h��f�M̻W[L�E=7*�	N�Sn�|gnpyJ�%]kcޗ{��)�M;x `�t�ڇ,h��,�����y�W�l^����i�CL��klyGbX4�˹Z�@5B�c���4Q�-���赑���O2�دED�i߽l��Lk��N�
��"���"b�*m�-*��Z�Ӌl����uu�I"M��Z*�,�`������ך�7�Vm��Z̩�Ȣ"v����j�8�������w���i���v�BT����`��XM��F�~g1V������mQ��A�w2S����WB�4�m�ʽjQ�F�ʯ&��VL�)�%�H���{X���N���-����e1V��_����E�~��Oo�)�+S��F��@4
�n�&f�v��i�Q+����� Y��fݫ�t����([��$͹� �7�����V�8V^c�����[JP�*��M��[P[��JT�q�$�0e�X��*�I��v�~eZd�H��aQך��;�2��L1"�D]2Y�5�:l�l��ٮqލx�~g�4=�{�\�y�o�i:j�fE�/2�� [�憡�{7dK�I���+k�����v�v�5�
h���s}�E:�K�V�<ݩ��Mﻛ�wn�	��������+j�����n*���b=T�G�fUk�b�Q�RN��n
���7N��cDN�VݣWjܺr-�r�K�V�oPL�v�ǐQnnBe��5�혲:ܕ�3k*7N��GUf�Jt�ke���٭T�85dr��Z�ݼj��.`�w�$ī+
P�b7(˲3Ӆ�A�.��'l<�`���.��w��2!0)S�t�2�,^˴�5�t*�˒�!JRM
����Gf�'U	V�T�T�x�#f�QYF�g\���XF�I����MI��N\#Bc`u��MB��X����(��o1QE6�]�
,�QE7h��5X���E���v�Qb�4X��YQDA�y�j��]�;X���*���t*?0EHf��y�5YjHP�6���P��:[4�&�(��-f%�o�x�L�6INQ��Ӏ��CJ�$ !B��Ң��><f�,Ơm����U���h�iZK��+0\��p����Z0���K)���P�Q�u��t�[xy�//�K����w�|j"'��0QF"��t��<��h��5�����:hC�0��`�͗|��j�<g����v�Tb&�q�!淴��n��ы�UۙP���E�lOۧA7Zvcn�,�T����V��ٵ2@�X����V l1vr� P~�h
�,G�V�a�<͚�<ٮs6��5��kB)k���h�x�uy�7�SH�(��DN2��3K��71��p�ֵ{����w3����2x0����`��rV�uB[��vmY"d��2�XE�_�P	m��9X,E��t'�s&s��j�vp��jj���`^R�8ٺ�.���kY�Y�qG�����KbV�7���[Y~�nbk
�h��p�lN麲��D�*P�	��Na����ws|��H��F��e�����voY�Ӝ5q�aw���U�"�nm]���!tP�mK�����d�t���6�.du�Mc���Di��㫬9��QRЃ��Q��"��n$*����!i��i(0����Wv��ƞj��(�vX̏�����4(P�n�Íx$��҆i4� Ƣ���_�����LԡF�!C7�;��,���1�Y�ݾr�M���ֹ奺�2�+3Y���M+�.�Q�u(�̄~�SAl�i�Fݶ���*�˷B�
�5D�ĝ�b;��v���,�vyC35��S�G���
��!��
9�m�?T5�f��<���<�$u�[7Y�q�tͰ�MU1�����Nl��
Y-Ck���]w�:��6ش�p�(�h
%�y�kl�,�WYW``��z)�6l����X��+,ߞw|Ɗ�V.�5�՛�	���
<�F&2�!�N�k�VJ���P����T�q�����Jh�bi쫹����>6,2"M�h���ciU+fW�iB�Q�Ɗ�'woP�E	@�sK�V75�*hB�A
 �bcSat��^p�n�t�y��z����
T���Y�߅��E�J�[�9n�b�� ��
+y��b��ꈗ��+�ѳ.� D��)
����` [l�N&�9��q�Q�Ye��ǽ�^:8��l˧��õT%��k�h��u����u��g��D�Vv�:a2��V,K�U`�Ѹ��m�X���S&d���qcBat�utĬz�v��6��X1n�Ն ���]�䭧.۬eT�Ҡswu<�~��+.�t
e8Ju�� ��yF`����&VV-�`%��%+]H�Q�shS�@e=��N�Ci���I~Vz��N oq�5�L̗�d���{�8G��}�o����7�F�H�I�$}$�����7�F�II#}$o����>�F�H�I�#}$�����7�F�H�I#�$o������7�H�I�#}$o����7�F��H�I�I#G����<8�������np�cQ�	��^��L��od�������峏"Z�O���ġ�d&C�l&��x�Z�#"�I$�%�yCȶE�l�=��&��|gf.{�$�m�K�����$����)�M�7�䎞h��3.N�mŽ׭�b�(���1���Y'#�ޘ�or�޴:�v�*f�ֺ��7��`d��F��I4J�I#i��'���_%݄�!L������u^'J�rKL
K�t�W9��*M�V�����eB��hP]�i����Q�*�c��W�!$o�˥ȤY1u�n�en���eg�$�oe�g2g-'�k rJ�����Q�d���Dwu���zn�Iq26�g��5fn�1��vv�@"�"U���ݛ��r&(bO��֒�7�SЂJ�����^�bK]�(��΢I��F�H�I镻���F���On�Z[�['�V�L�&�	�3-8l�T�A�7Jvvޤ��5"D�E��w_M�$Ȇ�GQwΊ|�Y�/����$x)Ȼۭ�A�7e���ݾ:���t�ƻVT���\�4�t�cPQ7������ܗ�¥&����j��rva�bJ6щs�>r��9Yw�����XV��w�J���J=Y�++��hăb%�noWuL�v�F�Ծ�V�P9q��{L�R�P�dӵ���c���;��5ޱj})������q��0�XK����-nTaun3�[���
Sr��n��5����C�%�3_:�\uGmܔ��(�ىwr׏���M�u|�c��A���=ُ�7��l	]y���K��.�ׂ�1�wX�&��z�VG��н�,��j���2";��'9d�RzJ�<�jX(lˎ]��ޔ�]A]T������Kn�u��Ե�zJs'\��r^��2�İ��h���]mv�i��ե-D�{b�D�ms��Vw֣��!���v��V�(K�n�7>ǒ��'����.�@l�s���ˁd���v���n�-��4�hu9�n��p,@GM���%�7tҨN*y�ގՔ���/^\����#�:��4V�Od�5�B�	EVR��͘��ɶ�X8ڙ�n��}7Yɝ��Χ�2=���b����I4Osm� =#\��ל2f`�\���.!�}4Q1s��73y3�8�L�0� [v�#��&�ۧb��GN�(��wk�b�Q�ݳ{1g6H%��K�Ly�s�"%.�`�I�/!���q��������鷱��#�ӻ�hu�H���Wc�t��֦CC��j	�7k���I���J��깺fv�D��.�@�L��H��i-�@Bs&�ė�D��v=��P�u$��C�����M�ͭ��Ҹ�ӒN�$�e��i�ĥ�2����I&����{��QfG�'t=ڐ��Ϥ'�v�������]X��;�b9'(�|��r�'��e��ш�_�$ �kR)M�$��;Q�qs���c��ر%��s�J${f���]ϣ�S{3�>�#˙��3�]��j��|6��1N��l�dI&�gn���t��G�^f.1&����H�W;�K�؃�Ҧ�GU߳	�Y�3��]Z8`�}rn��}�L�G��Ο�q��)Yb�h�\�-G�V�
�,Q�N�R�fq���ļ��$Y��������(�s�d�[�h�L7}0���5d9�=�5�*�]t⚮r0��Ĭ{}�v����ւ�Gu]]�dʔ���^k�����S�֙�[�(�Z]ۢ��E#�{=�^��q�T����+���S�Msi�̻�Ҷ�D���-�r��23w[F�J�ڶ�lK������הf ��0)�_[���	m!�e��y��++�c��% �5��Y�M��i��Lx%F�9��J�ZG��@Ӥ�"�엛g��E��Eڹo]�ݡ�M�m�� �"����/��-叹x�a��>�G�ݣþ,��M
���ښL��������k뵹�N-q�e��< f=O7*�/��q5�;&�4_hHe��6I�j�(���V¸�Ц�}JJ�4@�y���S��}��ۧ��m;�;�m��|�f,�|�p�Q�`�����#�^��7����58m��`-�"Y���s�K38�zpv5�A{]�� w�:��IZ�[WCk��wz�]�_H�ӥ���m>8�`�j�!�̇Fg0����)�5vՆ��Y��%Z,6���d��O�����zMv���(c��pd��)��v�f��Rk2�l��But��d�+8R�d��<�@�<�ͽ@T�0	u��t��̠c�:3�&;�5��穭e�KwY��WCzݺ��b�Z���N�7�W���r���ոW�GC��!��o`q���+U2��!����1m>�{��De3�c�r�)�/8�m��x�)��M\W��-�Q�+����̺{]G�	�9;e�l�q���Z�ɉ�u��h��c6.�Zj7�sr��a�zb��.D�{��U�O
4yP	�3f�޷�xk k:��r���b�lb|�g�_RA�t�nɽ�0w7�PȺ�(g9�$��.���u�t{�&^6��۝/+\��\eNvd�0����۝�$����!z���Z�Ѳ��un��ژu�d �2��E��L[��n�cX^v�#h���Q���,bT]��Lx��)�n���Y�u��ya�˵hd2�R's��'f�\�-B�V�`��p���^$;����(V	��ܻ2��/%9���oP��7Ab�;�M��޶�e<Ɖ�{o�Ю��5I[,�۬lS9Rl޼C}�	�H�)�X�l��i��W5Y p�Ǧ
�8�6��	H�;GI:;'T��;��{}��4âɠy�ݮu/tQ��w#-���o�B�ݻ�a�:�rۈ�0�q�uئtv��"3�6�]�
}��SQ<	�ӶB���r�Q�Ғ�Mm)��"��ȥ��-�	�+K
�̻�C��3�1Q�]uc-f�A*ky��Hãh:t^=�g����ɖT�m�5ٓf�I�����̛{��j�[r>�Jv�]՛9�G��=	�X�n��w�d�w(��)mۈ��R��B�k�X�7�.�۬��r�UE�x=7Y,N����	�v�qӕ�}-9Ҡ����Lb��m�ݺ\8ѫ\P��WȘpg(�V�-�E�f��Wf'iR�Ӂ�&e��%�[�QME�8�yV��1�X��G�*�*�)5v�mp5��OgZ���=B:��+�75���6�\���4✨м���*�%k��,�\�4t�Կ`��'�Լ�C7�bV1�;�<c3S�J��kB퀛�L])�^�K��̦_(��@K��o+�@os7��-k�;:���{nw�h�n
��˞���x��rF���ˇ��d�S��Ir�,"e3�/��]��8��Mj�7T�JG�L���e
���O��5��N�pY-{'|o;:6]��n���# ������CU�_V6��qb�Bͽɋ�{z�@ Y3A�\�Z�+����u�NM0;FJw1��I2���d��F�G��Y��	���Y���h����ܒ񼴢�y6H�43k@
��a��8;��ۼc�t�I�*QEut��#�,j�q��ꙙO���ܒ4�k���nu=*�S���r�W�in�0�o��X���]}e�-رZ�k���F]ro���^����Y��m�Z���s��@�iw.\ޭ�#i�-d˷���7:�s���nL����z�<�2-���p���޼u�RP�וc��Rv�T�'ub�ӳ�oX�%0l��sKp���&8��v�h��T�/#6/a��{��Q�8��m�x�%��=Ɗ��fneZYØ�`+�][Yt�/��iq}��6����'Y�zNI�'f�⚵�+<|���9��u	؂�wz�q�*��bk"nL�������A�&���4�pa!�V3�����⫭�VPe
�O% &�5%MK���ݙ��[�np�n.8F�`^�Y�
�1I�4`��^��-�� ��I��-l��r`ukܝNn�}:���[(��gc,c��e�6�X�ՈK���oz�R�C �P ��v�-6�E�����*�#�{���AЙu7����wj1�-�hj�[CrEv��J�� ����V�R�r��w�iE�."�i���;����У|oW~w���s�0���uI�u�$ͭ��G���r�Żu1<�b�>:P�q�tc��Jx�T�}��W�s3mE,�
S���\����r	�6ۢ�s�ZϕC�����c��N`�w�.J��ͩ�y���F0+"/e�]�iA�\P��&S��Π5�v�杷H�F^托��N�U�%҂xz�Lbn�׃f�N>���431���)gY�F���H*"���-��E?�6����ϵ�~�1X�:v�8L�mLm�G ��.��&���o'���f�$�2!	�2Ӑ�B�х��զ�n;�(��^C:��X�3*����漠��Q�.5��=�2R�U�}e5�k��$]h���r�+0-���֢���]�l͎�%*d�-=�(d�m^ �&��R_d�e�Y㗨&�+N#�5��u�k�:�u��{��{d���)૭����fe�\�}Hv-J���9{�4��cV��AM�t��s�:-��F�=诘��Fy���[!7��뷅E�KV�Õ�즛\w�M#7��v$b�e{��C�7�*�\lt���#-�y�[��n:�+y:�=Dꈛu=F���;,f+�Tmkt�~1SO˔��v�P�������X5�`]�w��=�5`�:��(ZV&��&Ԓ�+Oo���pMZ�:�^t���d���`]�v��4��/�S���Uԓt̫�{���Nո@(ݵ×A9I�.�m���ֱ��:�lǅq|��h�%��W�]\���u�]�ux������P��ڻ���{��f[װ`��f�δ�D.����Z]Ӫ�=�'Hj��(;�xp��I.��pc���{q3V%��z�*�%�+��9J��G)�
�A\t�u3������Iw|.u.�]�����ն_�3EhNH����*�0���%Jp恝����'I��Ѣ�:,�3�7���,��u�U�»�6�V5�z��(S��s���e�S[�yWr���\ܴP�%�=݃��r��!��ҫ�v�Dw'j�U����%��Y�G�e�yZI���L���W�	t�fk�%>���.^P�én.�:��On��Vf��_Pyp��4����Y����P�7w=�oyPshfV-�����6�f���	�KC�b��we�h(ƫ�y{�]���b�j�ݞz���"�u���
kk,r�4�k����n���̛u.�h�=	���m�wIfq�N�9+Qe^���r<�췋�T����ѝtث�hμ�N��.�.�V::����ֆ��W�7��u�n[��,uв��o,�R����ɹ��t2�{�8��^�z��@�e�SR��qf��ۏH���<�nf���s�q��Zz��L�v���;�0S����ۭx/z�pe�.ҏ�e9�������3B$���c��ECJ�Si��gs08�4�>1V`���A��ͬ;p�`���ը��K@��
�[7��7��t@�F�-#0�dQuLұoE7#	,�ژ��w�a�k(U�BoB��NIV*��^�Q�.�t��]L�����SeeX^n����x*͵/vF��ވ�QK��#��e�4A=��>\�CӞa�)jW�{y�}֦��1�\(���A
�gf9OBŧ������f�ևDb���]B����-��k��n�_�x���%��g\�x0o	�������7��<&Ս;�5Q���7�p���FTwK~9���7Hes��)i�Sz�Z���;A��m�����,eKe���-�C��̫�@)|���Y�սVAbV�F�F�Vl�k��IT��
�j�MB�;�[�o��((>��V�+l�d��k��:��Y�j��A���aM;���вU�T�հ�K�P�����|������Oo��jh����o�>��7��3X1�b��Ĕ�����C����ܛ[�q�f�+4
���$c���V�CFV8���Xc�G���Q\)����o��)kN���r+u�,�fqw��s��g�9X��H�)4�T��<T7o����r�眹�[�_g�WN�`XU4���2,��WA��4R���>*��w+o(zi�du�-���(�b��P1���#�ӺEX9��Z�Ǩ.�����s[��2�ὃ��q���#�7*ŕ���`���]C�ǢKC��I��Z��I�Eέޚ<�"��2�\�Z�v�N����,�vEyN�5]�w��\<z����P�g&�ݶ.Յ�w�܏�S�[gAys�n�9�73�B/�ۤ�8��h�%�:�s/���7!��3�k�x����Ƞ*ǼSʇ���cG3���T�m��瀬w��$�{n�4���wL��t�m���u2X��T$cU�EZ-c�MuqܠV��ԭ�/1uE6hζ��u]��\����|¾X�gˊ��#�Y��K�:5��ï�ܮ�L���Z��;����7�"}X��F`+(y�bFi�:Um�aaG����5���;�քw�.���k6�����$��-��i�bK�$#\�J����Z@ʹۗ�/5���o9�.3�cD�EWK����,�E��me+�in�����mfXʔ]<�nS���Ha��kc7%r3&=��k\�ե8��N�4g���h!v�E-���A4�AU�ǫJ�L"�ruj3&'8W�WMSe�V����]�R���&���	�[�8��.��r�kL���t8]���YsS[k4\����6�N�N�Q	���y� @!$�ђI'��H!ަ����k~�i ���� HE�M��R,���l�J��̒IP�oV��$�X�!�4 6�H B��@7��	.$${d���@"�I^!b@#��M�HI�	 q�I ]����	 ��HBd u� ��HC�Ci!�$��B!$��Xa!&Z&!	8j�@�R(�!{jH$!��9� d��ܤ�x�H�����q� $$4�	P����!|� z�
�.��`��� 4��Bo��I����RIY �A�I&�IRIXHVI9l	�	N�Hd�`M2�%`L��P$�	���N�!6�7�̄+
@X@�!� x�5�d c$�G�!��$(���̐�C<h��&yH@5�d��f�Bi��2BT � [I7l'�j�d�'ud��H�$sB[d
�e�!<a�RR�C�c(f�u�5�B�̒`�=߸B�6�[B� q1���1"$�Hm�c%� �	�K$�ٴ��(g2c$(��dĖ����wI���IY
ɶa�Ce�I����dr���d����5s$�VYM��<C���)�G�	��1#��hC�3)"0��P�!�L���&�I�偌k��Ią���@��!�F��1��e���Y'���ˀ�P��l�(d7��}��A`m&�OT���[��)
�g���M���C��B���mXɴ�6Y�$� b�i��&�O;��1���ueM�4��ӹI�]0�cD��("I�TP��x?KV�
�˴�M�7{[/pj8�v0 �m�Vs��9�"����ռӕ�q?� "����u ��:��������fk{�0X����Z��n�n6!���ɦ[�Σ�����lھ��/o.vnu�dT{pV#;%��aGʞ#���X�*�_4v	��]�2J��}���w5nЙkd�Nfu�/����ͼa�1�Z��m�G/�E�	��L�������R��1���о7cu-Hdme�&�tngK� ᳦�;r����8/'��,���ɝ�~�ɵ�c�T�P3¬ir�CH�K5��:�4��6�is��aV��I�}s;�ٶ
�d��&�v,�nvA��D�B�w^WL�����ZS#�݌����{���<E�}z���3���l\��*Ƹ��`V�*0L۔:�mN�,����]�k��K�R�DԮ���Y���v���x�[��z�^�Ջ��	YWNjT��iP���:L��}X���v��ya!��+.�UgJ��Rb�hN�N�ݙ���������8jT��Qp��@%�I���O���p����u�ǉgi�
�]�����6lj�%��\@�t��u^KW/5��-�*X�;Tz���ˌ�X��R}ٗl=Eg�ͧ����B���
)�3��ѥ%6Ve�1��������ӴWM:s�Ό�n��K�me.5۽��Tˢ���N]&
�vӚ�\��f�i��/�$�����uշ���ܻ7�8��qt�H�)���w`��\Ȝ=���C\C�u)*�a�u��Ø�}��y��$�$�k��=���Ϗ2��3s���_WX����V8V�n����j�5o���j��JC�����ҏ�a���vm=�癆�q�:�Ջy\�͆�`CfG���� ]�͊�e�o����\�+^1M`��t`����}�T��\�{���μ//?��,�l>��I���R���AMB��i:�i�pە�*��8���
�Qk@!�2�Tk�p+�<y(C#��0�v�^�Wwp�����Sn\饍{(�m\�[��,��X���Kj�e�{w����OG*����V0����7�<�]}�g�]{�P	y��Us��v/����D7�gup�J
�^��Ȃ8wP׳o�𵖚�U]�=Z9j��2ZI����C��UY��M���@�:�[&��$��d#����1$�$XEDD �
�sy�nw�9�߽�ޓy��&�=��0��q�ț�Ӕ�΅gv�ŗ"�7T���9�߈"�z��3-��ST\��Ϲ����J�`�q��[E�g��(��Z�z��^;�^��\9�Ȉ���5Ӳ���1�qs`v������{2���:�/��U^�8h���[��Ԕ��N33.��o!!�ܘd��r\��?l�_P���NS��'���9MB��ܧX�F��J�����z�]�[�hG��]ٓq��d���-q+�>�L+"�U����+9(��Y�˩S�r<ҳ���4��]��]��n&F]t��f����L��QX��z��_��[-@�T奄*j�f[o4bU};�aeTLj ��B�k��	��׽O�M��ĺ���x.���#�����#�)�˙my��j��ɪdt�M2C,kJ�((�@t���YB���0�p�v��n�}4D��u�lef������Ur�2㈋1���t$�$a��6⚍��97���1���m�A���M��˥�o]��=���j��ʥf����Rw��c�� �p�x�,��"��&�^L�Tr4
_E��r�ua)��ے됙]I_;��^|Et�w�^�߀�������h���Q݃��$��l��hs����s9�}�<�m�3�5�l�t]oϡ$4{���~�]�{�*�b��ic��Ѐl�.�����]�a��1+�����K��z'�Q���f͞�H��<3���>��W�]@'�q�㧙�*������R��f������]S��#^��n)J�"�J��K���E����´I�:�)��N�w9ݾ"!\"MA�k/5���h�9�y�v{��<�^j�v��Def�R�!pAc ��n�㠱C�˸������%�y�w������{;�_<���o�UG��/����W`������ղ/��px)⻢6v�	���vc����N�7@+Z�V�E��#��֣Y���2楫^���r���չ"��7�(lu^����u�;��ץ�>�W�^ئr��u��~���=��Ļ������
��ژ!���q���Am�m��XFDFu��r@�����hz�r���29a�]�z2l뾾F�����1���; {�s���/��秛rC葀,��������=3�f�w��_k|�����EL�8��h��wq\\Nb�;�W��y�\=�s����{��=�s���@� �"�|��2��3B̹G�>��{�x�}ԥ>�Bi�elt�y���P��cZڃ8ԋ��f��+1U+��^�<,rÈ;s).9/6��	���J�!�����kC�Mm4��t�5S`�,Kn��V̦�n�� �ª������N
��L��l��7EY0��S����c�7��Vf����S�^�&"Ӏ�ME��� ���m`�Jq:�f���3���sM㤴����v[a�é�/Uz�i��b�jb�v��UY�z���p�i��k ]f\���]>
K�&���Ң�o��\�Up���u��Ʒ��E���{ު���7I/k�Y�X̣-G.�W�����~��p�O�u�zռ��B��K��t��g|ߙ�{�<�]y���_9�^*�iy�o��'=�ː���#��Km�1����x���y�}���^k�} Y��y�s�N��=���$ �s�d�0rTUŎcl,JX�ʪ�[*!U%"�Z$Ud+k
�Q����Ȉ�q���}ʚmg��i�c�՗K��Gw;�֯;�ݘ���{��0�u�*O[�{:��4,;z��V-�d䛹�rɴ�ݥѫڲ��\H�1�U��u�,k�k'*��P^t��ހ�T��L~�P:T�jc{�����߾�|�fvi�F�jbz�����U����G����o�p�}�Z��!H�i9(�^���3C}���vq��x[ֳ��Ec<2.�쯷��t5=y���i!��і�{3�ٵ�:��`| ����g��Խ��`���]��ZGp�Rt�w5v�����/���'7юr�U�FP\UUA�m\g}�+f�'0,�Z6��۵"�ʃ���W�_}�2D�5�`>��\���^�^���I5�$��y���3Z�_�����c�<n�Tuެ��\fa�64D�ͮ��������O9s��I�cDd�`@$"z;kC���u�S���O+����m�u:T����h��m�������'��m)x|�b��7r���2��y;�w�٬�R���r��{�c��}��d*�\�z��q3YO^3Y�pX��ne�+��C��5Ó�L�h(����s�Rq/����t͛b����r���:WtW
��H��q�O;��q�hq��#�� �wRo���es�����]%-;N;�����5`U����֋��y��7�<}���}��]ѽ�Z��O� >|�J&6�8�����VK��U��#��wa��[�D����+�;���#M�ô�{kx-� ��]��6b)`o{�A��˯�lđ�)���wa�hP����P�Y�3���7.$d���
`��v�W�$6���.^H7r}����{]�չ�i���w�
0mæ�cMH��2
L���U��v��4iu���T��rTM�\=�O�m�ՉZߡ�+bS;�[�\�M�]"u:6;p=����]Rw���V�*�I>]��3+�ǻf��伊v] �*�̼ާ͎�z�`�8Fu�a��z�UBB�ϗe�Vg2;.�]�u�,���'��Z5|�ڕ&�'-V'�� �l��T�y]9"2��Y���9��Itֺr�J�3(͝��~n���W�g���3���_HxD�@~�`��[���3уջ�طA=�!��q���-|`d�N��B½���^W4��T�-Q>�*�yggޯz�a���lOٯ�������Z��$ndJ"k�z��T�ڴ���UpԹ���*�w8�`  ��o^�8�5�Q���N��ͼ�ٹ�VWM�,v)�	ʼ'jj�/{v�;�}���}瞒�I�H�p�ɖ̌��AJ��F�+i*��-�ڧp�y���U��y����;����'t�#{��>yٴw��On�
!\wx,A�gG.�z8��rle
�/r,�̨+^�\{ŧ�u0s=���+ï��<2�tenU*9��u:���Q��G���g�u���Ga�}զH>+^�����N����oު�6r���^�د{s=�y�ߔ}~�B2��}�����)��ɻ��Be�]�J�=֕�;�Na�6M��:��W�L�)����Aݦ�g�tű~�\�w���2ov9�ֈ��C<Wu�LիcܠfS��о:*7�DD����9��;cK >����W2�]��������J�O�kz��)$C{Ƕ���w�����9j�#  }x;�>�6m̜�Ȋ�6����7��df�UT,z�ݹ��~��9҅��1��"
�\��5�8ӯ�ri϶��n@�A���u�%��}@MJ����Ӹ�Ycp�zc ��f
��<m�ay�b�b���G�6�v��+]���� �ge�^�Q��j�4t]�s6�Ė�m"����\�`03tI*{�R�[U;�\oN�{Eb���и��W���t�������<9�o�ۍ�c9Pѵ�֌v]]��sBܯ��g#�__ƅ�^��ܦX�^nV>�F#C���_� >��K�Qux�lM.�Z��^u+Bg.���g.��p�A�2#�r��oh�2�>��UC��]�y����Ol|�_s�+���})��7���v�U���gy!�r�)���.<}�����wz�޽�3�I$�~;���ݞ���y_c���8�u�cE�]E���(s��;{�b�R1"����"�b��4;�� ���:��r"�Ӹ �q���ܢl��*4�s/8jx��P��©�!/57�\@Q��UQ�/F�/`���j�}�*���r��wd��]��I��ۆ���'�#���!R�˚����e�cWU�{����q���C��s[�p�R����#a['��q��܇kr�^WZ�VC�^����P�]r%�.<��<ã\p��D���4��c�:y�h�6=y�4e����X�w}=�+E|q|GS2�Z�gۢ��X���׷r�T�	���]�<q7��i��c�������O1��w�5�K�i�-�7��?cA��,8�S��?pR�Qt�*1Tb��+��y�q�,�a�m�鵃s�t����0�#�cnkY���Z�t�{.�k��M���,�|���[%S��E"�4�
��eT|n����h��SҨ[BA��:�.Y�Q����c�(�WN"[� ����n��'������+ ��0�DZ  [-�4�#�hVt^���CW��9�r�P`��ys\�û�-�����
����\�إ���u�6�i��O7�L��}5��W3�7��@1	:�J�T��$H�� ��d�,��2�*B���#���7��͋��}���Z[�`o
ZV��0�Jw/�\��_<(tl��G4d�V��y���m�kw[ݖ�紫F�ׅե�J�r�b�r���
�t���k2��[w��KUo�(���ﻤ���Nx�{�'n�wG�I䥗:]���I'�%�))M��w���&v�=�$O.e��(m����D&���n�y�im��/Xb�m�A�<s�T�ƈ�٘x����.V"7sD˾8c[���փ}�ަ	G�qV�/
��*�G��D�)��c]bݝ�x.!���B5'�[٪�mV���u���g�����g	���80��c)���ɜ\�V9�5�u����r��B����:��;7�ppx �� n�J���;v��d��YL�]z�br�v��ȟo^2��ξ��v#��3()}�S�f��pnA�1�r`)-ս�M��k�v)z� ެm�C�Q��;���wct�M�nՆ�q�@6T�|��{��5��6V�Z����b�����\���wML���7)�잧�H�^ͮ��b�t��q4�wwb�E8�KTB�ʱ�j�#�n�������^��/����y����ܜZ�8�JR0r�.gޮ�����)\�w99p�׳�	t79vº���X�v�2�E$4�v7ܹ�&#7�Z��'d4�u��ت\z�S6*�HLQÂf�9���u�j��׏pZ��ݹ���;4�����:]5�Wj�Wu��U�G��$�Xt4��]����t�D�ќoT<�L`���sIĚ�ge�{`��|�9�)[�����ފ�U㋪r~�!�|��Y���n�v�x���-gǲ��k9�u�V�b�r������q��{X;��.��5k�vml�Ȗ?���e��P�j�w1�H�GF�?4���s��z�����`��)w���Փ� ����n�<�R\�<
T���C�W��_�~���'R|]>2h/~p!��.�@���&�j��CU-��+�=;����>����!ttL-8�@��׌��m�reL���ׄ}5���iv)�+�q6WV�D�RX|]��8�����ߎ�$`��@����@DE�$X���1�,QdY@@>�����Ow���N6
1cGl��*_�S8��o�
�5�?g�p��_}\���k%Z���;�s]���}𣿻��{��+����^����{mj�);Ƭ���1w~�X�v�L�i���_|���O��
Ͼ��`�uU��4�-ms-�݃>��{������_;���짯�u��lA��ԕ�f�9�nw����)0�J��h��*~��iv����d�>���?�!_r�(�I`�, �*w�|x���"�6���E즏@��9'1�z�b�M���죵%�Lv���I�l�:��O��a��5�2�xw�	 ����|��x���X���'n]N'�R���M��������MP��Lp�ҝb ;T�8Y1|>���\�1�b���S��P���<󶶗aW�����bWZ����z�DƷ>�$I��ٖ$n+=	ީWZy���<� ,|>z%`T1{D�`s��ga�'�+WEnE��@[�Ÿg��	�^"ߙ��7^�k�/������s�U�� �j-^���Ͼ�$�Ɇ)����g��u�������6B�jr*���������V�;�=ҮG{�:)��π]k��a�\��{G��  +\���"�q5��aYۯ ��3]N���e�hVk_z�����}�v�ۧ�s?����p�����4���6�Y�X:�P�X&=Hi od!�u�χs5|?���8����}d�0�bJ��d��w�CS��'P�iXy퓬��P������N��B~�O�٣#���� �/١uLH��!Y"�K*�Yl����O�Doy�y�Z���٘8n+uu������;r�똍HS��ށ������툁z��z~tĹ�;�RJ��sS�W8K~�]z]{/�Y�	�߰�5���'�8�=`y��J��x��o�L�zϐ�6B@a�{��R(O�������~ַ�����OY"��L�l�O}��g�yԟ$:��I�$����I����.��I��	�"�+��e����3߼��޿����;}!Xx�`��'��M8�&04����!�i'Y>��'�$ ��-��u��O�%I�}`,�OY4��2T�O�o����ݘ< ᙡ+(g�Z[�~p�y�2{�d:� ��Nr�+� >�v�y���9��$�6/z�����GT�Ba�e��4�P�_�z,����_�-U��GW�X����>���gƈ�L9��#q`�ɺ����+Ҟ��N�� ����<���JG�._����g0����׶�;LZ��W[��W������KCY63ͧ��:��܊6%T]��HL��ͻ��|��}��������=u�s�)LJ{ES�+.>b��t�j��L�B'�彗��E�ޮ�(�V���v�q�f#("�? >|
��f|�^��e�{��^���6����3$2�"־p�gJ�h諸�w8ьܬ�5�	��-Q.i���J�s�k��kPî]��f����5�&;Vn��[Z���%y�<U������O�w�r������4���v2��<�f�̮ˌ���/���o���k��HwO5�����|�_�j�����MV�v�{��tn<!�䅽j�r�����WBe�,P����&� r�y���J� �� ���� �\���e��1��!G�V��ޮa���H\��|�ey8�2�����uO�1���A+K�"׌�|>����=n�f��H� �w�yB�"�q
��f_ne��iY�v��j�_"���q��|�EA��u��POZ���/�0E�~�����]�y���	��̾;7�~��y�}��G��4�A�Q��ķ���~�zLW��ߌ�������ME�Nړ�a�˗��ߛ`zy�	�G�9p�a���o*�Su�}��膣���UH6S'���,W�~p�uD�rm��Xn\|�joZ�v����~^��=����c[hX҄�B>��}���s^��y���m���n�ʇ�l��K*</�{��m�������o1oJؚ�9����r�"]�Ml�}G���C�I�$��W�~﷚��}�,���kK��^���s<��{�1�p���"��nt���WД���(ǁv�~���j|W^Q�˩��&��*��?z�n�G��=�]�z��1����>r�+1 _���'KF_hEF�{����[ߧD��>����G:�|��]��f����������h�H;���S�}��
�~O�ۃ��/��Z������|%�ї��x�ń6�+x��뼚'jj5����W�����ė|O�(��ջ5~J�Zz$MC�������Z�8��f&��3M�}�vV�ƴ�Zm���'"�@��ޘr���ܹ���<�-����k!$��L��E>�]�3{+�$���S�萅�Ǵ�X3�'��|~�����;��R�Ԭ��}�>F�mȷ�����۽�O�@PQ`�RQ`�`���
��y�������_��[�O�ok�S�>r�Q����5d�f\����Ҥ�� �����d���cZ+���"�0AE��c(#S.d�N�� 1}�ewP�vU������P�y�p���ܸ��˗NcR&��*.���]��`���/8Pã��Cq#ñᗨ�u%b9���՗����������}m��p���E�7��?I]��=����������;�z1�wA�y�� Ë$h���Q˔�%�#�;�Dc>��bkʆ����\LLQWBe�!�ϋǵQ�O�  ε^�*uT�B��Q��;f�b�j�7���1݋Oʗ��E���cs�9���t&�0j�OwfZ}��	ܟ��PU$rY*׽8&bo�|q��š�[�U��܎1s*D�.�_gH�Q��!.��h����o[K�ݩ{
#qI�|���7�  ��u{��k�������R2V�}�v�J�O0�D,ŀ�y���!� ��E�����"�<2zw�%��ϸtƉ�F���| ����/������0�����ؿpW��a#W��w�����cy�(�O,�jԘ���(�ŵ�@�|>��2��y�rPŪPH�	P�ʍ�߼��O��j���M}��-�9��tbp�<�޴sz'C%�0�=U��;v�'����Ժ�~=�Ԕ��� �����&
��;���w۽�p��U�U���s��ܐ3���	j�cISs^�$jgx��[�9WȒ�	��<�� �<>}��{�t͡3-ː���7Q�ͭ;��P�N���]F��JϽ,y@���_�}w����ׯ&��.�Ĳn�D�[e+��!�}��A^7"u��6|l~�	 $����XM����QY��1���I�>����	�A!����o���S�}��-�����f���`ͮ�%{�37<1rj"��=k�R��;UOZ6�7b�*��9�y��y���e�g��L��޼�$��7��9Y���`(l���.�}��%��3�i�F%����B����?���|�.����D�⯊gj`G+뻬S/r�Ͽ�o_��y������;���z�^�o��]"L�(u?c�Q��*�EsW��pIc:��*�[물�Y �Xi4���u�|7W_';�|ֲ�:_s -�����di1Ճi�.��u&�+p�Ӻ<���+��u6���5�掖i���f�F��M�jo�f����n�{�m<�m�y�>�i,�O�A��TP;��鴰Y�oweW�;O��bjDٱeKF�Y�g�*����cC�g�ґ����_{���2z�;�g��|O o������sZ�y�/��{N��]�6į��3��T	�����p��ЎXS�}�T�I�^!0��&���s�r~�]�j�C͵��ɏf������|)~���G�W
<��&*��Q�7!�u]n�z�S+޴nb}�@ָ�./{�A��Ԉ5����|b3��[�V������k�!���g��kZY=}��.�`T�ί�j}��(�{n1���P-�ӕ\V��sT�z0�������A��R�ɐ�O�/���+�*pA1��tc+.\9���D���=�{ӧ����~�>���R��F���=��׺�M������@ ��]32U���<�
� p:����9���F�[`�+B��a�x�V�zo���͗�,�l��a#(�D�q�LӯwK����H#�_#�\]�LavP��P��-�h�&%���]
�N�L�`���4��k��[��f��j��^`��e)�@�s:ݷ�HV��vR[B=��*�/@�[�;�L�l>D�ll��5�YV7y�cr�j_�R�o�q=$��[�����y�GY�_��C���ɏL{k��2��q2j\���I<�K���9\���4|5��Tsb��*cޗ(�8C�nRq�U�j�A8��R���m�5����߹�\ω'��Mӡpe���K�dw́��Qa�S��7��y�k��TD��?�9�m���+�iBhb��F�{*����#�ݳ�J �HZ�{#�⨮�� )���������s^�s�>�&)�Y`	���,F(=}w�1B].F����F���a�+)"{o����*/�3��W�J�'#O&�Ea�zt}A�+���˴ �@�$a@}r�*PY.�&�y0��вi�(C�}1ރ�,���?�R��'СBcg'��"�S�u��g��ZT>�� �:��-R�6��.U�k2�d15sF��2��u�%)�( ��U!EJ��̸H�FB�bLH�UdXVV�����!D#	�)��+(�i���K1�2@�(0�`B�h�(�L��(H�� !��|��|���k2A��\��Sz�%�v��ARCP�4#��������Fu5]���]&:w[4�wsLAV��`&n�m���x.sP�4�;�;��|qޮj��[S��sx�PAq�2�]I�ϤU�#'�n��_��&��I�Aj�N�M�r\�B9�eN��"�>�}&}y�E��?Á�i��ʠ+��܆?'��E0k�(��Eq�h?�y_���Dt��/�U��ѓ�˸c�����E�{#&{���y�T!, f|>f<*���G�0y!�~�{oy7?\���YR$=�Y>��B��Q5���^��]��
��iN�������}ۙ�\[�3\B~Bss���g*"G����_�)>lo��'�O�~"��]r&�$�)�=�KIR'E��=��+ةX!�k9����8��uu$��N;��h\G� Oo���^�_��>6�޳������h�ix�����F�=�<�����_͊�l�<O�K��c+�Y�=�1Z�Ѣ�"��+
���%�W��Y7��ު�N|������� `���G�P�8Z����~���x��Џ���7������p���S-��ơM�j*T��h�21��]p�6u�_��.�Y.:%�8���D=UO�;2���s����IՁL�
�6���)�����ɠTJ-��Ak�Z�u*��"�]�2�n�h�����<t�l0�Z�@�@dx�S3��:�բ)�o"t^q�ݳs��wD�Q��XQ�G̮;b��s�I�;�u��É@j��=״ �Ԍb2�mM�|�_Wu֮��ߜ3g�y�/_w'a�BB���1��H㵲��]n�����^�����Uw�J��5b�D}�	"	 �P�rF*N][��Ę���T���wR �":�Q�b��x� AuEQ?���ұf���tK�EGYj����Ӹ=k���u�f���R�LK"��c?�WHZ��k!�����:������_q8�
�i�۩�دʰ�Vɟ�4�Tkr�b�/��#ˠB�O[:lg��vLs�6��`�f`�)�RC��`�fS�R��)�(��ԯP�e�5Zk*�@����z�>Z��y�<q��NF�[�0(�1~C	x囵U�V�n1�E?g��j���y�=��xė/Y�WT��N={�(�Qd$ݔ oO���˯�`��+@����W���ebb�3��{�6���
�Ay�ou39�I�[T��j�p�[��"��B��Z�0����ц�
 V˩J��7�Z*u.���tl+�m7Xz��]&O�Ѷ��N�G�\��	=��jJWZ��sy�:IS�!����RЃe��5�΍�Ӱ�<w
��;�̫�0ծ�gsynM����枧��8��6��Tڏh���\�\�'Hq(s/ 0uL��.b浱v�1��2���WM�����D�o[����'x�b8����o��v
p���h'�b�mDo�����}b���*n�%����-��S��o�r)���n����� kKݖ�}���,�mU�� L�q�&ɯ1�Š݇��܉�蛥R�Ȧ\�h]����s�fd`'Ʃ�3"fu�a�:��.-�8#���˻�u�%�H�[�M>�nJ� ܫRJJ�t���z����[�3��{*�a�l��y �0&������&���nf��
��ٗK(�>*�3�}݉��W��4��o,�T?)��k�b�G���}@M��$}�Fe��38]ĵ���si<��s��Cr��v �G{���ԁ�T��J����^R@����!��yΏ�Q'?&�WF�j`�[׋�λ����0vؽ��i����7�*NsacV"К���h�ڸ�1:����.�ᕮ�
DF#k;������� I��\y����҄9�Z���^l�@[�yg�P��4p<�()�n�̕ni��:iKF*X�����짻�*�ޔ�.8Վ[IH������`��u�9�qH�k��9�J�;z�s�����MO���w����՞e�8�^;��,w�PU��0nka��GS��os���I�K���^ip�����\|[��W�S�h�
�Y��ҫ�TFg��>g���e��	�����^o�7��H����t�R�M/�"N4E}���r0�rRK��6����u*�U��:)!��3����{�;q����}9[J�c�IF�Ӿ��>�d}�s�잌Q���\Hq'��%3뗽}��	k�L�(b�� �ֽy�dM�IJ7��KR�����   8>����zl����v��8*`O���W�mT��P�k�j1�+.RxU#�k��$�_)�uOu�^����7~v��l�ԫ�E(�_do�|H���f���j��h�_��wͰ�TT�׏��+j0�Ab�ZW�sdG�%%bQ�G���	8�X^�SW���ǚ�cd�_L���eZ��>T�"��D�ݜ�P>�_���S� �g0�߫�!�������7���{����.o���e6UP�y��V��y1��6\T�h{$G��ǬC�MX��n�'��u��B4�Bz�ey}���߿R	�)���|��1%H���o��Y��J�"P�\�"4E��F�6f�m��U��DDDq�+��1QH8ZȰ�Y(�QF�m�F�b3��C"0QV�%��4P+,<��e�(�f��=�KK�����w�;��n�OA��	JJ>謚SC.�l#\������(�j�.tѣ�>3�S;K^��h����Wȶ��^����o�z���P�Ե�H����]��j��*،�y�6#���� D�C\�0�y)Qs��2��=x�"k����S�0_|H�-�_W�4���@�T�Q�]�]�TG P�3�+F�
��S����^SV{����g���Bvx>y�>��{�O���R�Δ�<H�&�opҲv�CXTG��_�����>�,��`0���5����0��7n3Ñ�4δ���^�~��r� {};�.ʯ"���T%&!%2�<[
��`�7H����īM��A�NFJ�b�KyϨ�a����zKyG��4ey(�z�M*�Y�#ԕV�~b�"��!bAb�FH���C����;�j�y�z�Ǿ���۫�Ћ���mP��CF�����L�_�O�6�M�+6,��t>p��&S�
�)�-n�3�F	���2��d�_��2���sŸ�,�9��vz��u�HP�9{P&"a�F���B�d/A&��J����|��3�l���gz�����t )2�`Tm���μ�<���k��:r�=�^"��|���*���|f�]Y[fF.=n�����d2:�z��r�VR�l�yBH��9�F^,�����Ҽ�{ީ��$-޼ֹ_w���?J^���ߺ*���P�PNp����ב���zM�Ĺ�h��>�#���O}����-%^��ٳ-����]#��	�!�{��}�혿��$�@6�F/�����6SȂ�LJ1��Q^[��G��h�n8x��f.v+%n���*'�D����f�;ȑ�ш��2�����T��^Q�}�y�Q��&����V�1U���dp�&V0������^_oLTF�`�N5�;�|��fb��R�9QϟJa~�[�گ��5��7����ko����g��M4��7�|��o�HH$m�ղ��m�F��遅�80��A.C��^�Q��#8�#B:*s�gu�s]����W7�h��B}�{$���~���n���M).~UNdNK�v��.s��n.�L�#�긫{ɢPA<4�ϳZ_�r�֜����|��i��us�7�$�v������9�?~�ˡ��W��q��_6z��+�6ܵ�%O�B7ؙ�7��+�[Jn�{����N:Kl�K�юS3D�`9HJ!H,�ai(�s Q� A��z���`�^+Ѳoic2�O���2�P��3[��3���nm%��Z��D��Q�To��|���Y@��I}y��[{� a�'��j�l	��`�k��9�4��n�po�;�7��$?@!rf~�ߏ���n�?�S��ڧ|�#
�^�v�GBǮԂ�_=�y3�3�k$ö�B��}Ac����i�}#` ��� ͩg�c��H�}>x�W^���+[���ɜN�Y׎��=ކ|j���r�n�ߤ�G�T[��Ƨǎ2z�h�7T\���Τ'�c�~�pA/k��/�x�3k���r7�Zq6�55 �7y��yD���+�"�z6V-$�����(`�W.��A��焄���CgwǺ�k�ߛi���Os�� ���$��-��`a�����֏tY�R^�ȸ���ǗIa�t�fő��
7��|^�-���F���+����s�Ō��S�����L*R�wc��,z��{���L��b�}�vߛ8�xr����W��-YS�=������]Я�XC&cr�50�1�B�Yd*�$(Ũ�!,�R�PPE�#*%���F)H���U�"�XV
��і(%��(QX/ꢍ"��2�>�Q��{�Xm�l�:�:�1.�s�/�R�O���m��M���@�Uqf;��"{�}n��t,�\1�@՗3#�J���E�mI�8���Z���+)�N�����DR�幹��Y��Sw,�z�O��ԍ�o_*}����E��	lX�v���6�����c�����
AcPϳr|ud_���~&1G�0ыO8�����ߝ����.����5�����HB�
������ɔJ���5`�_u���x-�ͬ���RC�'`�\�,R�M=�n�!gc�>�A2��7��t���5�}����6j�C�\m�>�l���#�
��=���S����+�����B;�"`�������^��P�C���_�-������N����Kkx�6 �A6bv3:n�)�r�6;d0An-d�����ВL-�]3��Mk��������_����~̀��o;󀥣�q mW��y�r�i_[�7�/
?���8� ����▗12uʏ$<�X{�sz�g_�J��eF1���.�#���d&���LK�ɿo<t_c����31l�6���`������f��COB����ƕ���.Ǘ�	�nv���S���g�Vs��C>r����]�{L�(����%��Ӧ���%��Ja_pwİ�������3�������{eo���	��|�~�����|��}�D�Ɏ�=��zV�w�8��E.ُ����s�vg�%^�~����Q���I�+� ��Rˁ��#3uOPCc��A���#�OĂT���K���	���w9
8�H�y,ݞ�9zN+{t&#���'0e�ݻ�"�CJ9(%bY[-����}�3��� �$�o��w�����_��,�,�C`I��$�ƭe^�I����]妽���MEL�P��k��Y����xnƑ�VK�Ȃt|-� +�����ũ�H-���>�I�f�c=�W^�6R��v�WqΦ��`�<�glba&�%�~��e�]�;�m���Q��ѡ�8|��ey�^E2=p/��P\�h1c�U�D�G����	\mXT�9.�?{sۙ�=}�~v	|��="�jI\{I%!�.`�٪K�v���1;7L�+i�S�p��l���b��#��f���i����u�=����?zuL���ݳ��^���/j���K�ݔ6�kN.�� ���������������AH��! �H* ,"��j=���>8�''bc�8�Z��a��VV��:�(�}Y�M���͗P̛��|sX/����B|W�|������q7�c:ɣ���b�SU���Kx�^/ȥ�i8o��K̶_���?x9�K�'�[ZD��"�mR<��x�Ǹ��|�)Tv�\���=V�Vq	+�J��V��´���\��HwB7� Arl�y�M���3�)8^���[+:�髧�}�~0�8v��|.�����o�6�G�㺘�<q�`�O�agl�G�U�Uw�=Y�b���Z���˚�o����K���۾g����w�&�I_�|?ob�,�G�����K�ZZh?*����йt]#y/[��i�ظ���C�9�1J���p����;�ս���ؖ�L`��׽��y��}:^w~�Yp~	m��.Ox�U�����wm���s�V돺8�^�V�9@(%3���:��#�K\y�v����竘��)�گy=7A�EYq{M��z�=%>�Mr���D���3Vb����L������P���Lm�]���,�����?{ �2��?g��?f_G�����?v��WX���x�{���q�Q��N���C��K��,����,��=�HOn�Iټ�̾��5���߻�=�%����l��Hئ��u0qWǌY��6pܮKˁ�j�z'�R����������ʗ�zks������> |��aR�v���?XWaVk������wc�9����E����w�v��������w�=u�3s���NzI1�4?~�9�Լ����$�G�CɄsF�?����v+0kɞ�����k�9o���-��7�&Y�9��jOL�	�����z@�ϝ_���潺�������^߼���oc���i?���5�m/�=]�zk��|�I��3&fF*�T��lY�H/՘3�W.t�.�5ϫS �v]�4��sOm�A�2A��r�ݏ�Gz�~YF���"{��ѡ�����Xٹ_i���H�@U�P�/�|������ʉ�k�t���Z��]p}6���m`��e���2ʻOR��!A��mu7��aј��|o��|�1d	;7��[���[p�8��G�H؄�/۝�G��)":�U�ږa��T)ݓ����Ri]�s�L��^�ue�\C��	��Xg������o���{�:�G��(g�#������2�s\��^�Q�����������=��Ͼ�{� >[��<��7�֘��f4NȶR�sc��j�@�j*���یv]�����K�0����0�u��ި���c�H�R�d{�Yy�3�J�J�D�V�ˊɿ�&�%W�òVj	���W�%}J���o3s���N�&
�$U��ڂ������X���h,A��<�A�^@W���`�D+Fi��2)���J����cT�UKe�c-�*2�me���ZR"1�R�]�Z�u�ξ�_�u�{��K�Zڿ��r�m�e�3��I���+�S�(`��}]U/�J�(Ǔ5uW�ùs��]�C1��Hg�=y��ڤ��Y�Ix����|4��XʤXݪ��$�u1Q����xܳ_���	?dT�y�O��>�g�\�����2%�϶c�3{��y�svU�6{�֗W���;}*{�B�`���F{bsy*,S�#��7+��g.�kg������sj�5����hE�;�=��#���7"���[m�����fn�~R�����k2\�E�}�͏8G������[9��[�SRq��%I����	z`m��kЀ�^�a�
�+���$���F�[=U�9=�צ5��v >|=���|j��'��w HP���x����WH�7}V����!�Q(`���'�R��:9ő`	��0���=�4��km;�G���H�H#�GbG�zp���1�YC k�����<��>g�<�ֱ��/���>8��]9�݋���y,Sv��7۽jfYF~�p�u���b�dɦf�s4 �=g�)/��-�u�WI*�3��ĵzv������r��U��L����ߺ���Pm�O�G�;����'�xg��gDb�P�ח����g5��ޞy�^F�뵀P����Ep�v�m-���d�J
mh֞�G���a�i�YĮ�J&�V�MASvl�r�;���ȪIvD����3*��C
�.�ɽ�f�o��0D!���,�\���˭��������ۛf#�:�Dt���(V��8���K�`��4���ɺ��	���c��V8ѕ��6j
lB���bkt��3V��3�,�?�*"��� 
�R�mcb��*�X�s�,9JY3(RH�)��5��<�5���p�g�w�s�gi%��Z��рQ4���Y㎎����9�:Jɷ}�P̹�����hv��X)��w;ͺ��5�5u�YXi��WvHc�����e�u����f��Q͝�I �L֛%H���8f;�l�`���.S��G���� r�<�r�14��i*6�K���on`�m	�P�N��A�(�{J/E�ܩj.6�H�F��!�����G�*Pf3����'W/�-k�I!ڜK
�e�״�y6<��`qq�A�>L�ۼ�D�[ɛ�����S����d���<o�M����>O
@Bj�&�;!�74?9�g(�T�nAi(,� ���c��xm�U��3x��o1l`_3�x�u]C�W_^_>)=F�W�m6݊�И��0*���Y]��;\k�&U�������� ��,�R���x��o�rT�9u߷Dy��D�vs�]�CC��u	9O!��
V�Wd��f1�9e,V���(:��3��ǧvvPW��^v䬸�a7Ι'c$sډ)4���r˺�L8U\�wW	b�.Am�Etk|՗מ�Uv���)-�z:���(�_(��l��
�uHfX��8��޳&u�i�#�Orwu��S�`~�*�v�����޶���^Wm��xV��9-���:�����i����F��ׯi �mJ�J`wFu����&���)���hs �p&��r�a��� �ji-Ԛ|���t�y�/;xc�P�kf�"��n����
���Y}��Me�C;/�S���m0�L@n^4w��K��&r�Z^
�j�3u+��1���� �3�/��p�/{ �/Y.wIE�r�;W��e�v�p�����74nta��ov����w�I;}[���=��UW����Ug�Ju4���� ��yW3N՞Qw-��1���Q[���}�K��x����/-�7�V��DA�� ��seg&�y.��>�o��6�8H��J����<�q�\�*�����q����c&vL{�@�Lx�+f�V���~N�"�x#zC�)��F2H� Xg�����N��W^Y��h� ��*tC����>�9��#А-<��L�Ex�{���F�΁qi����jD4�P&��
^��{�*V�I%=���$x<��v�G^Xj$Z����0n����_Y�q�*��Kﳲ��R�]�p�/�1!4�Gl�L��ߧ3ua�pV��_[�%48���-�;�x��ծ��ETO��<^���r���"9t)"7ؤ>���M��1{�����{�G�{��8}ބ�4@ByƄ�W����k�uN�\�2h��HfD�8�39�OFl�fa�{	À�I���]aۭ9������Jg� ��u!���I[ޙ7�}�=!��r�����z�z���34��堀��`�5��²3+���ˏ�y��i��Z��on/)N�^�]�EJ��ٓ1��{�.T���ж��y�������Dڦ���h�h���!X��Q!�[SS�{��o|����1���5�}u�����,��ɻ�\X�g��3N���P���� �s���b�&�8�vz�B���i�)S
��O�E�V#�� ې�2��p�3| _��x����e-�E�@b�LS�Je���T��۹�,���}���]>g��7��[�Ϯ�g~o?o��Ԑ���GDwz����ڕ��)m��/��ܺ�y��W�W��qˢL;�5D~���������$PR?��ʻ��)|>�� (�5��t���S96W�������'��hq��9q/���Z��bЫT�]rM�a}�%{"��N���c�~�0�@�G�����R��cJ"���Vl��X��PL�Q2� �ݏc�ߦ��b���4N�e$���5ZDb���h���a���W'�M�7��Cl|�#��$����\jHE\������3�9�6���'r��.����yé§V,��m�we��)b�kU�8Vv#A�6)���$3�'fM����J��g]Jl�ndi*�Zo��˾kuh}�*��
Y;~U�"���s���| �8�������P2����ʁSi{�ꫪ�n�C�ʼ�0�{�s�Θ��tsR�tօG�S/Wފ����\�V;��J{��}�׎(��ʼ 0|H�������Q�"���(�^��w�N
��{�wR1\[�yi���g�-�&��;pH�@&�͹�X��)i�=����Br���CO	���T���3Ĵ�XnpW�Ί=�U�n�GҖ�Ć�wA��`�R�!���~�~�;�֫�r���}�����O3��n<
��f����h�^b�>�������i����"�ݗ�yrE$�����[���� `(@P������;��N�Ʒ�~��_��m4P]ӯ�`�B3��P�s���j0��y5�V�Y��7���H��ji.7kMi̹@&0������$�Be��ʆo^�鎜��ӆB��P讳�04�v���.�I�ym�F���	%�K#�f���5��7+4^݄����y�n�ã�1����> �i�n�g�3��e!|��8TG_��j��鳻�(��:C\�A �X��zpb%�5�lr>��6�ħv��X� ��Nx��!{�$jC�8�\�z8��"F:� C�}NfMԾ�G.��+P�^�W�'����V���r0���+�R��*�Z}.1`P��{H�*$���^�M8=�8�Qִ�i}�|�Ps�5|���Ox�T��W]��k��H ��g�wQ���2� �}����|X�Z�i?/�����$<4���b��Zקa�\N�s�n�1�����׷�s�6z�� �1��`A@�) ��/ߏ3�=��^}�_D��.ڍ��ݟ��p�4hgn��W�e����8Ѿ+y���F�K��R1;]��XN�ݢ�02�����+��hO_���eFj��@3Vcㇺ� ҁ�c��[�NML�&�fK$b���!e0�1�X�*,�Y �\�c!1�b��QB���)<��r��VMzD���vvU��Xu���kO��Φ�Y�B�[��c=Q���14䳀>����Gs3b�sp������\n ^��G@�Qأ�4��ӈ�������ULgZ��r�Ǿ��Y�1C��k�8˜��աa~CS��ƴt���⯃[��	��T�ɪ]<�oC�3��sG{1H͟}��A���C�/-�`U�#^C۹�f�a��˄pn��Q��y�4�6|�=�M�p��s�2Rt���};y�o˞]R�y�'���}�*[����1��_|2mk�b)�)� �F�9Y�X�FIU�����d���fIՎ���*Y��y������}Ɉ���>���^�C~�YhV.w5W�x�Ȇ5�Fvcm����Jr>���:Ꞣ{w:w*��Y�yD�Zu<�e�M��*_���������3�yqr�^]z��&\z(E�5w^Wpz�o��62��o<�=�-�S��|÷���y�}�j��{�BR��w�a�^8�`(���H�a*EH
�"$��~w^������{���bTg7�HY��v����QA��;:�n�C�n%�u;�ҽn�i�����q+8�Q:��ק����dK)���{��dBe�N̶ve�����cсɔg�����_��iy�.�҅v��4����/�|,|"�C�
���~�f/O�UQ���J�ȕ
%�&E`J{%��h��������߿w{�GS:|u3���#e|�Q����9�����x�ȨH;���{әי�7.����j3ǅD���!�Ȉ��d����F�����i������/.�K��$bI`B~��Z5z��Hw5d�D�#�k��՗�b/QD�2��������/ހ�>����V�{��(�e##���q��+���~��eo�FE.��ԟw�RV|<���"���ca��1<Y,�o1�������y�ls�W��c蘭?@������O��ۣz=ǝ���]�͔���.��Q�DhՍ�5����c��l�N��x�Z��"G��=J���i����C�G�M��M�4�����.���m�:t�7��u�q���1��`P��g|cs��GJ���!@��dq1s?�yY�^w�lZ���|'\��O��Å���<�r<D^�F��1&�8I$�B#��;���-K�O��	���d֟��3���
9l.��t<�ƺ�yӋ}Gp��Ǻ4���������Jsƒ���_K����.S ]βa����"|�6���'�&3����5���C���2��w�~=;�N��I*�a�^fg�Qɐ�CփwXm��C�}�yO2϶��+�R�X�������?ӵ�Kd@ʥjX�]v��H��]�Db�y�^8^w��"#5��3�Y7n) ��̓�%�+����W����S�Mӟ�^�<[	�R��h�H��k2X5s��p��E�r��yr��}�K�>��:{`�	d�5�5I�F�EP�02��b(�=ߚ�Wn���zs]�_]Z5�p<;��[��u��WBan�Q*��:�I��Xc'S�8�r����+gf���)`(�ǌ�9�c�]t�y�u!t�!
��K�|7��ei��Xa7��t�~����=}�}R��Ao�h-D�( �Ι�YEk��M�����`���iZR���>������Id("��/��>}����3V���
%�g��'�&ׅ׾+���~�d�W���:z���mN�+�xM����ֳ�_}�繗~�Z������� I��>�ξ��;��I�(o�=���<*wN�aK뜔�F��_D�H�d<��t�~����{��1�K�Ӝw�����z�����k���^��T�W/_sR����z6�m����\[�9;dq�o�ﾈ���b�ץ{�S�ʋ?h)����s`��:���$��K�� ��TY�\OZ�_֮%���?�ԩ����C�RvA���s$S���a=���y�];�%����|k�h}�-�S3.R�VD(�2��s-$�K*"Ă~ �����ۧ*���AQ}(�Q�t�2�
޳������3�W�C�N�e����l��R�ڠF�n�v���L�ő�\�>���]}q���؏��z<>��Ψ�2��0/��~ь�VW��xhw?^=�����QQ��H���V��$5}˅��Y=�|��1��c��>�z�V�rD10��	U���DMe3��̨;T�3=(�ܩ�h-�+8�8��.[�+�QE�+����>}0׍��uM{�
���t�A�-{��,�ܓG �ݾL���|-r���k��}i?��oo�r4�^���X�<�g� >o��]��(�c��$�,��q��J�_Y;U��P�-:&������g�q��u�=�0)�񶳎�K�K���-l=�/Pl���x|/�"���N�(��[�1!��5Г�����>����ꐄbw�
N�68��5�O���d����` k��^�Y���@�9���S��D�k�y�4�c�e�A#��yL��0d1�3(��K�b`�Pq*����gw�}��<�]ԮWW��u�tIඵ�Ύ�W�m�o���C$`�m
8��W[�f�Օ8��o�Fw��Nٌ�o���x�Z��Ή]!c<K�\�T��s'ۻi���
@�Ȟ��w��8�������z��SυG$�}�T�.Ǵ�.V=���x�b��+/ΥwY��c�D�d��=�&
��*Ͻ����n��>�s�I�"/�|�̛ػ:ֆ��ts��`�2�r�5̚�'���Dwv�&�_(<�}�=}�7�xn�z��@{���۵�_��q�0�#��Â�W�=�q!�Ⱦ��䙠����gl�BN�í���j��D䵖���S;'����>	�G^E��῞�����Kc�����Ϛ_���<H\mT(��d������Go���7��wϻ��H]�߾o������:J�E�W����K?c�F�#)c��E�ڬ���~���˿U3b�֏}{jgg����������ǟ�%xM�u)��%}���o�HP����!ٻ�dv�I�%nՉ�X�"���tVI���^�HhX�*(��5�@\f�G(�G*M��n�����f	GQ翮�9*~s)�cQ	�,���,z�b��7]�S������Y��� ��%'R�y1��u���,�C����Q�e.ٯ�����]qY�e]	G�9��eu �hj���z�S��IPt����*�~� \��VK+e� w,��g*����*')Y�<����:��-����G�L�k���<��&9��z���y��W��]��|׺�:��h�Y�(��e�5��h�R�������޳:�{p��W��T�Zy���k�2�o��[�7��T����ʃj�t�����` �{�<�ɫ��=חg��C����f)�^SZ�Oz��tʯ��]�ۡ�}Zsvub�F��y=�}�u�ˍgX4��@EM=��黛f&k~o{c�4y�d!�:��!ADб�S{���EV{l���m�qib��
Vr�Gr�D���S�4��,m%ך΍7��!��͆�7�桭��J�f��)�}8�epK�4�z7�3j�������D�NH�}#�<�R4�.��0�\�wzJ*n;�*�`R�����F���Hy��ϣm�k�t�ݝ;[�e��g�+��V#��t׵�TL��:]��K�7y��R�QWV�tރH{)��{Z�L��.���Z�{V��X��Kq,���C����Ф�u�i�6�on<���7Ş� ̛�tb�f��1U�c[Ά��
���m�]������6��]�5�din��n��t��-56 �>�`��L}��vŌ9�t#��Jn7���XK��̦R䉼�H/��w�A���-a��:Du�*k�2��Y�����T�VF7w��|��A럲���;sWN�:D]�,�;\����Xr�a�?X\�wtlڍ�0����"�Uv`{']���a0���W�R�.�w߷���i��@'s�+��a���5A��#O����F;%=|#�7�����h���g�յEy/��-[F�sA�xF�ȝN��z�^jYEE����q��0i������duP�=v=�Up���Me[�(=wF��Bf7�� _em�}�`�;r�bT���@@��X��B+ks��;5�o�R=2�c:M�A�.�>�߻o����&WS�3���i�pX�}�7�;�9�}G����X�[�K5�
z��O�u|{Wr
Y �)<>����1�����Y�T�M�Ԥ�O�;-7�cW�����}����f���:�Z]II�e�4R)�)$��N����0/��/'^�&g�w�nu��)�Z��Ѹ,&��>���c����1lI��/��ys����a�g#����}U�GR3��$��[�I¬ٗ	��뫱����l�OLmD�D�Cp	�:���yr�8G6�Ly���w��*!W8�F�Ϗ��%�����}��}��t�@� � o�Ѕ����XC^�El-�;Q�m�䖴�������e�X�=�5�i`�y�?�� -"u�tRoV���F� �Nsy�
��V��c�[�p�8d��w��B��^=�a��U�.מNœ�p�n�I�faz65mJ4ȿ�����̹����Byn������������� �5�^�k����:��Ϻc5��dN!�H�t3��D́���ޮٺ�␥�/֞���˟o=�|��׿�,X
�H��G�ꁓw8u��]�������y�k��m��P�{��XL�,\b�ٌ�o�s��y��{�v�F��	F�K)B�`T��~���{�뽌3�׽
�yNZP��XV��S�{x��=��]|Y�*��Y�M`��\��I5��t�]^c�Y�[�n����o9tէ���L���$�G�����{��!�T��D�n'9�:׫��9��2��v�c��EM�f�\`*��ՎD�.�������W{����3j'ae�rH�B/��)A���ۈۉvm� D�T�/����fj��{��}-7ˤ��=UQ�qS��9�����ܢ�1�u��V����;-`��9��[��vs���]�m�r�!}Z��p��a�>��'��j��"z�a��hDR���F߯=;��j�e$;��}<�9�DpN�y0;/�{�Snz�eF�����De��	d�/�A+�}h|3�v���i����qiظo7���]�����Pψ�\zx�K����C�yH7���me;��<��9���.,��o�y0 ��M8^<e�J��iZ.ǜ���	�����Y��f�*J�D��
T�=�{���}��ُ�;��f`�C�h֊��t���iֺl�X��[�t+6����m��+�EGd淵-�1�.��\���3��G��6�qA��knlb{ۭgo�����mHfd�'�����U���z�ou�?wkH�AW�(4Ú�� ��dM�H����"��w|o�I$�}}��W$i�l�����.���Ǟ�������®��J;��h����0s�
9�5M�T��N���s�J@�7v�[7���<�߶����<�.?m����$�%�>������~�]�|��I~�|;����f��,��PӺ������_N:�Y�u{����G��f��J�	����� 	 � $� |bk�8煹��܏U�L��1����3�3Eo������6O(5�~՜z�_���>�7���&�=&KW`�e� <����,�R�����L�	�[zV%��v�NS�Zl6dN�"�]!�X�4v!/:	�ۘ(i���}w����ٽ����ѰՕb�IU����H$"�d�"�d�!"�1T�`�u���
i5u�'�}�r�]f�-�m�����Ϯ�e\�Ü�z�i��ʴ� b�ʵ�k]fN��L�y�c�^e�D�;\��Z���X�}��o<0n!Q�T�Z(�)u����׊���x�3r�1a�w0u����J'"�G� �Ƀ�j,������"��N��ar�HD*:�֙�(>��Rb*e9Q�r�Ŝ��|>���i�M�;9]s��rEx��o��LG�!zc�u}�]+�aw�m�q��ػ�ٓD(�u-m)x�c����9��g���9k_+���.�j/(��}н��|	�8B}QH�Y�NQ�菡L���Z�����HV�})c���WtQM"V��޴���eK�䎉���3��+a{�zZ�8��9�w�Ocu��C�k,>��(��M����%���Y�F�н��E��t��| ��+�~�fka����[�Z:<5�
<!:��#yRYj����n!����G���W��<����ER<,�k&�̺�1ud�ȕ�F$��0�قJ�C����]�v�q�t��m c��&Wumb�Z�bf��^�pÒ�/�����˗��rW��*p�����xf�G�����^�i�'�� ��3�u��s������H��.fyJ�	���!���e�S��5P=��6B�4�Ɇwe9#S<�"֘��u�V�:���ˋ��b������5�I��{��,K9�=P|T��\�g+�SI
�-���]Pz���'���	J�t�gPzU�k�c�����"A`����<y�{�>��ovY���gN 9�Ӯۥ��_�|����9i��
D)�b@t��Ԥ��b���oNyO�S
��D��=����ŝԨ��ȟ��n��eD��r�]+�`�Z���y'm!D���1�t�;C(Ux�@!�\���G����D��o�d����bM��Й��GDI�B!e���tP˜#��)�yg��:�)y��䱥bn�rJ �~_w8��y��JUi���o:d|d\�#yni��	T!�a@.�ZߞC����n�H6��C4I+���Kj��1�Qȉ�я:�rV�E��]X�]��i^iK����B�>�qʹ���8�3s4p��e�I�1���(ka/��-�=y-d�w!��}��g���M�k�5Y��A��"FC���y�Z>�7"]��$~�W����rcM�H�7���r!����|=�l<C���l��=�g�28�i��X(9��o�7/���q���5��.w�{*,�=��r�r2=����bE�/R���_��39ݾ�D:�x��&i�|����>p����V|I�vOz���]�}Bك]�:��C������\�0=��|=[}n0I���p��u������Zp��9��Hf�	�\ƭtC���F*!`���Os���%�Պ\����������},����C6c��(�Q��l`��[���0;��diI��YS�]L�!���̓8Գ��O��dRѰ%����VH,�a�K-c�\�R�"��gmD,lu��JY�"�l�z
�#����c�q eѾ�֭�l���0`��!�����r�)tD��<OG��օj��	�ԦQà�PN	���d�7�v���u�Թ�n\&-�2+U+��]B��)&����}�|���Id��f>sE��￾�J��8�{��X{���U���lpo��D{�U��r���E\�u��c�zZgz~��͙������:&������>��M8Ⰶ�mt=9��V�T��A5�ܽ��v$������QF��G�NQ�eZ�K���E�(˧�V�^���"��>���/}e�c_?,��V:�ưd���@�#3{��:hb�]]xgf��g��^@����Y� �ܹ���}��q����őV_F�u�*�b,��9�=�#�6�o��62oW���u�3b����#���}q7�{q�7br�6��%WҦ����a�[D���a�C�-���2�������(�H	�xz��y���}��5U����ŏ�
5�ĳ�6d��Ai@e_f�+q5]�2��K+�N���m���nM��C�%D2^wm��]ړշ�$勴�����(��ti����p<'�Y��z����	���c̘����~k��R��s�ұ�Zd]���w�ם5��oF�>7��]b���w��V\�z6J��ݱ�{�[�����<�.�qcT�w|JOx��*F��"-u�p��Y�A>�m.U�ɼ�]ą~��*�+�w�5���I&���N���������f���k!�T��$��.�4՟N�o8�+�b�q�U�� �ٌ���^Iw"w�wJ@�򺆾�`��/�T�-_�]�p�B�B�d���F��Z�q��W���jt�֑5#���*�5 ]������<g�@#���*���h ���Qa�]n�g_�CC
���{����0��p5:�ܡ�(Ԯ/m�*�&��v6kj!�AR-"��g��|>�~�O}�]���z���s_�P�e,�H����$�`2,!�
�bZY"
�"Ed,bF(
��!#$c�Yg�������e�D�*H�Ī�h��	[�𙃖Ƴ7y]��jt{6���C���;���C��悒T:��ݿ�d[��:&IW*�l�^��{:�����Xb�֏ajx�Ӱ��ؗ����]�&�V,��S�	?<}]���ryta��OQ��"��zPR7J^��n9C��X������3��[�ӳh���Ͼ��V��r�x�~y�~����Y؇���_>u���t�҇R��U�f�b�(p��=�����B�����ݩ��
�+�N!�n���5�<Kɝ�u9-�(�90
���KS�rI��j\DmA臽��f\�ʷ4�v���~�|�G�|׬�;��ϡ	/}<�G]���E|�������f6{�g�-�~q�e����7�ｑ�_GPn>���uT�ʒwcQ[e{�~�� !&a���=3A.HsYJ�`f����a��B�_�'��Q���]���&UuFp*�8sST>6n  ���\���j�1�j�R�u����8��1tZ�^��դ�x*!�)۱��9Q��4����:��wغ"��slJ&����Ȱ�-���]-��w�S�w����ׯH�����Ɖ�^�
��@9�$��dA=k�1gL�Eu�v�T�و�|���s���>%,/B'�fJ�n;���>��|w���w<�rI'�s{�4z�j����̧��DGL)T����2"�{b���W�^���}�eEc�&�e-��GG����G�~����ÿ�0ѕ{��kg��B��ʨ��e�_\��ɟEƑ�.{$9���Fzc��e`��yz��}~�0���d�D��k���h��u=~M~t�{���|�?}H��5gdԢ�#d���I���pMʕՉ�Q��Le���"���5��������/kw��<�n���~��HT�P����PHU�gB;��yp�0$�~�>�n�7��mb�h�պ��\�)�uˮg��Ϯ#HI8�3���m��P7��>���k/��m��'�>���5�(���C�M�V�{�62�x�u�Å�PB���5}ٳ���-� C|6�������B��TC-�~�jH����3{�ѿwݼ���b�£v�>V��
5�S���������ۛ=�ti9�n�xQY�o�PU<զ�E�.����{��sI����;eI�jN�uݽݖ�)w�Efi7\��BN�I�^L|J�ͱYK)�[��f�u˸�n�_�F��j��5A���i�;.n��T�zk��|�=|�i��59��i)�k�L��u�u�D���)���1m�M�L�7w�5��wy��|9[x�م4�fo�ӻ��(&�.
i5R��R�VTA�{MoXo2�k,���f�&�:�f��X�q�"�=�@�@�ˠ��B�7�^��Y�y�{p�<�vZ��&U��eR�waU��K�ńۭf�۞��sc���y熸�;ДL��p̚����8�.������y�e�l�_�P����"ZLW0 <GQ��I��&�4�A�Һ��5�q6��wΥKq1���iEʠ�Jn���L@�u�
W4��3��/K����f�mҊ�2�T��j�bg5Zbw{Ѭkiɍ��bVL����JV�r��r��7n�طi 8�[���Io�}#��c0>M����ݴ�d��JCj�ۈ	Z�kwN��lg����	� �[�e�r�t�R�R�-�9�7�+��}i�Crތ�J���_7��<���G������p�3ĶvWmI�6k��5$��9.ų�D�xvK��p����M��	Y:X�[�p��ۏ�sj5٠6/��M�����^!�����Dҕ�p��U��t�
�v)b,mA�/���x:.)ˎ*5d�!�J3Э�+���\+��-��F2��Sa�R�>���Iy�/�.]��[��#���'X�e$�<�q�x�޶OD[)�Ro6�;�nw���g���쮇�op ���"�F�Y�:Pe�z涠�P�:ﻱ�Ih�y�9Xhk�ㅰyˌ1����O3��Uz���]�{��D�ާ��&Xe���\w��7i^.ǭwk׋��s��˧Ϫc
�.�ߝ��T���e�]���QU�� eU�zI�0^M�7�*L����7WYO��orw.o:PZ(�Pmgml���kQs�ٻ&�&2��q%'`��/D�x��=jS[�_LQ,�wY���YMRR�oSU+V�<�r�ḫ��c�
]��j3^�{OL�0r��x�ǧ�
S�^�+pr	'+Lj�����W15���S:f��,$.��L����v�*�+kP�˔6�I-�!�<��뛽s�[�nHĦ�&��d�ޯFb�w1��7�H�r��hsЦ��x���������u����}	έ��XX�E�ׅ>X����<q���Ż��wM���l�?gK(����ƪ��b<��h�U��%ހ�Z��ސnWo�Q^���rȕu��잇j!_9(��@�NX����6o6,��c�z�(Cz�����5�M0��tZ��uO�.P����	�^]'��dg��M\pWP\V)|vD��J��
�I��U��>Yz�nFfO9�Y.q�wʽ��_U����^����	�c"�g�@ݏO� =����$�F�<ݖv�T�59>��r�p�������x�;�o�Ut��6*�:�d�>��٩�5��:L�<����;i�W+�8h���t#mX�{,�>�DE��}��R���fe���|>��5���'�Ϸt�ϼ�U� +#e�a���/����i�D��(>���C�םf�����ؕ��z=���:=[7
|��}g��.��?k��2)fa���V�ZU�
K��~�5��y���/9�&D�d�oQ�
��zkgs�]���ewn5Ӓ���-�����uw\]4�Ĵe����C6X賈u�Ws7^��F!�=�>�F��D<�d�JO��/6\��8^��pz׈'Q�r,�&�M�����e�D����<<j�圳��&gNn����C��=j	��*����Nŝ"š��b��j�}=ص��>{��u�ɰ�U�TE��T����u\��Sȣ�F%D�H����ɩ#�{W^<���b���Q�V����v`�.�oc���?|0H{�:��.:o����>$|��[5y{�})"�A�
�.EuG��S�9���!�Б��#���snK���(p��-�Oj�����?\)_=��M�7$ߘ�����,�k�Ei��mw���� S���U�3׽~o����Gm��sIC#pm}Q�ƙ�uϷ��X���*Ts^sv�a�u	'��~�׵�t����^Rl��sbFd��W-���;�~���<6�ڈ�}̙pfB)����걕�K�|OQ����Ƥ�G���I}��{gt�OV�!k�;�]�".�^r��N�
���{9����T�ݗQ76p͓Sl�f�M=��n�a+��s��F��5=FF�D�!ׄ_/R� Z����6X����,s}D��t�]�N��·��n���D\up�Z���"���gq֩( {�>��̣^0�z�����xra����y�n)ϓQ�l(olX,u��k3�y浛�o�5O=����a	'߻tG9���2���"k�q�dE��!�.��^�x9��~w>����%�!��߻�1��[q��ysbj�[)���X�S�qS�ϥG���'����Z�b>�c=����>������=�%X+^S��X�̞�;ו�tBًk�|���|>S�9POHR]�A�غ�f��z\�6%5F�u����0:�R�\T��r�t"#�;���Z2���;A�8ÇN�����T���9�C��OA������1�"
�\nB���|@�و�0��0i��e���cj"��$��U��AJ������+�(e��$YZ+
�2�eJ]	L����;�.q{���e���ޣ}Y����+�]b�P�=KV˵���%h
�E�KX��#��^�����._i,p~�o�A��P��Jx��f��W�����E�� ��l���
9��@ozDa�2��O<��_x�./S���ԧ\BS�94$Vbc��r33�ʏ��?SR{�u[�/�n���t<$���ݾ>�S�g{���ǖ+F\ WD�=�g}R/˼z�/#�P^Η�ڟyי>�bLV��PR��뙎�aҖ���� �dB�+ ��5�/~�\87��iS�R�q	a7Қ���-��]uF��o�z��i�*v��JBtY �*7��a����Z�n����U�|���I�{[�c���{7����hK�vbo�G�X]���XS���|+Ϩ��^μkA|>�N�:^՘�j�f��H"{LQ�g�ƥu��ŧ]����t,͎'��qGc�:����IF�E��;fߟ�u�t�1c�2L-s*`��I
�dDE��"Xs{��o��v�:n����ꝿ�Z�Eǵ�v���0^<���O�Ч0�rk.�R8+�aR�a���d��r��n����$���9���d�.����7�dn~�`��^T?�A��ѯ�&�[����%�keK�ˁMV�C>�f�G�E��\s���FI\zF��q�tʅ.C���UF���Ip�ѪO���Ө���C�wr��p�w�8�{��zd<y:~��6v, OC�{:�="}��@ɝ=+ٓ#�SJ�\���0�I��o�n���^�����_'K��j�.�����a�c�֏�9�l׷�~�ywWn$1���5'�F�,L�ʍ�����d_8��1	�^Ygn]e���+��ﾾT�z3��Cܸ/Z��I^����j. {}�=�qm�7+�yT�.�Y�k jBt���ԑ������{�!�J���W����㻹�S��NJ�^�a�"-�3��:1��sʅ5���;u�W5oNx+�x2��p�-fd���y�����9��gp�
��h�W5`on��U�z���!@1��=���V�ZY���8��++�K��sil�]fDvk�l�ۛ���%sٹ)�1Ho���<߇�0 �A��<�������c� O�z+3R��Ŧ��3���Zz|�wU�۹庣SH�3YzH�f��Փ�9:#{�Ӌ`ѭ豠��e�o���g�_�鷟j�+�3��:��Κ1�D4���㕳#SӑR|���m�ʍU��`5���+����W�<�E��~��Q�$�F�1��Cal/h�,f@�#,|e�֟�HU�.���#}F�-[k��/#־`����_С#�r�L�{8��0p1P2�.�_�Z�P�Z���Z\�86�@=;��u�u�d�c�I�����v��㿩��o�3����o�9��I��=�:��$b�����2�{�VB�b��P�NM"/LY����G���R1��f��\��7W#����|O���J�u}V6�j�I���	"~ �DTH�_ct\S#V*��! H�l��顆�k�(�?p�8-j\v�J���=�P�;�W>Xڽ\F;Ư�nԘ���b��R�;Z<�H�f���H�QkmG��w8q����.$4��:د0��t�5ge
gb��پ�J��F�i>ܟyC@���ҾH����5��u��,�h�3�ߕ�6p^Ƒ�&,��r8>�1���%[�I�?[kt;���Ţ���SQkY�U�����1���#��  ;2!y�)��n�pP��U���!�X[F]C�O!H"4^��Y@��0�c���\ɗ�j���~�ﾁ�U��|1Vt�(97��NVMǴ�o#"` `�T�g�^E�m/�{pkXk��R�c�ٽ���5�jP�[f���/��Ao߿I>@���"���y�J�ӆ�U������U ��t3<!m1���EX��ow�"v�rw�Uv�*��s�s�s��u��@�k��|��9�S3E�iD/94:w�M����I�6t��:��7����Xױ�}n�B!�|����q?&����8\2pLC(��$�� ăG%fF`��)��`�&D��cl-џu�ӱ�E�]��;8�dS��˷b��[')y��w=� ���`��}�G�s]mp7��*�:��on
)G�ٷ����62�~��g�z�_��>�|�~�p�ח�-���qg_���VnA���7����>���1Ѥ$�Ʀ�5I�1�k?����j�~�[�����#��c��ѹF�K�%v+At.�3<��bC0������ڨFC��\^&@�
뢜 ���bq#�`����/�q~	�k��&�D]G{����`�%lu�*�3Hc�(ӕ�K��ܽ���D�j�c�)ZU6�G��< u���l_�f�fxę��U'�;�%[��ǊsP@Y���!�D��D�Uƥn!�ô��<�c:�aXkE�x}���h��M��b�1�'K6�\]�ﲲ�d��Ր:\mK���'��X;!j���C�w���gj#��U���c<2 �29��dt���HT�upm�=^�O�#����CkZn	p�rTel����E��Q��J��K����j�ˣn/
x�hAu��+��3��+�J��d�Ⱦ��p�%�N�V��v��w����e� �G]b�T�<f �������,��t:��R,�=j��������� ��"Ұ�<�������_���u��uy������3�)���> �m��z�Dxu��"6GC�w���sV�͙1[IF�yR
���|N���������z�v�)��v�:�H᱄{�{|��I�:p��}u&.a����T ��u>N�!f0��3AB������슨8�(f9Y^{����C|��y�{�y^�l�MC:�/.`��1<���p��T�k�71�t ��۰���4��fW�����ljuY��,������)Y��~$������_�uڅLd� ��3.�����	�]�u�cﾼ^��i����>�^|b�7����A1HKs�ɅS�).2�Q�������N��}�ރ���mgֺ:.ЉH�,CҸ���V�� O���8��ُ�;�߯�1M�w���ő"�d3�y�f���w����4~����70�s��{xxeCf#w����K盅����z8+Ss��R`Nٴ�re�騅�kkvL���iX�b9�u�٫wo�X0`t2Ƥ"�
SQ�3o*G^�z�,O��M;kq]�7�����<��m���ky}�y��w����m���ٖ��"����93{0&&]��hVx�.�*�0<4K�^b���.�Q������{��5�S����iy�9UM��a����c��5�A��!B���#��)�Xh�[:������� F�N��uo��&s&u@>}�>���F���F�d�����O��+|IR�j�0'�☏*���Y�Tr)�8��}����>�^����G�� �jq�����Z�+L~Cai�X[���=q4�oԽ::*��%�G`�ġsV�HVa���|>���}r�0 �o�,�����ǻ�������=�=�&�Ť�p��+�5N��b�~�r��l�p=�Έ��e���s	�')[ �)?y����p��};��w��m��۝�m �)�@"�"�ˣ�<{T���f�6Ј����2�Gʴ,c������5�Ms'�Ot���et<��M+H���+���K�fT�V�O�q�$����y�9;E'�.��#�:�����O�Ȇ�
K���P�5)�G9�u�M�{��V���@+"B���	�\�N���76�T��7�hֳ����u����C���0����)m�]�̦J�:�c�0M��w7�\���<�CH�:�p�tV��pm�
�w3�$���42,ESl�s4�ֳ��Xt���B��[����hД-ATch
����aL~u8qU�C�Z?��Ը��A�{;t{�q|��E �u�[|�O�-�:�u�["������s��}��L�4�w����Bm��z��i�FI�%w�zn	�{�[՛�0͙Z$ASW��mʊ��x8�b���ʫ�s���y�<*Qx^jۓ-�f�"��Z{�d�{��	M`���4�qн�����h�ar��1^ �]�0$�!vz�;ם9�q���ws[��R�9�5�y�'�QI�V�˯3��ڋ��d2����c�Rv�t����������as}�RJ6�"b�|4V�ú�"3�6����J�3�o`�k7�E���÷'fw-�����#w/���ٓ9�e�	����]�/ޛ��(i+��f�`N��_'��QD����T��V�ͮ�u�RR�d\�(��a<@s1��'��+��Z�8��!G�u�s����o�n��}�ٜы�W>�b�gwW�iuM@�Qr����`�x&n��uj�X����|]��W.�^�cN�|�1��������p�`�ϸU��Rۜ���y9��H�
1li^��;�D���&묃����@��rZe�1K�����H��mu8�ʗ�gzt[�� m�4�:m���;�GlE�����K���5��)�KPZ&gZƷV�V^�����n�汏�/�ȋ�m~�a͝�kh��l�W�$�n��R�l]���Zm�	y����K���'fG��+�w�q�j=����rQomb�Z�G��N����x<:Dk��s��QwȊ��kV�Ӱ�6t���2��4EW:��^E�T�uk��mc2A�������}�������n�|�����$LuدѮ}VUɯ��Y�ۘ2V�r�6��x�s/�N�u
o5&��&�*7"��9ҺJ<7�������ێpK��1&����4�.̣5��W7��Wᕘl�ŹS J�M�Ss�q�����66������Z�U��غ��e}C�z75=1gt�M��pZ\�e5��N��x�x�`ҩR����u�;]���i�M��mv��\Kx-�V���l�.���7�^�è���1#�V}����
��JUy�w��}"B���PÁ+08�rA��\g������3!k��c�.��7Ҙ'���8��5N����[�xf9�3��^�c��p8�����%�0�m��&/��U�f<���g�4o,�h�?~0]���4��z�0��}�˸y���4��GGP�5����:��`�*9�D_8��\��	�{Tg���/�N3>�)�"uA�w.�0�Cw�^�^�M��s.���]���4忏��xh�޻�
��ً]��@o=S:�f���z��l�/���A��9����P�_fD��������)�����Nv�<Pȥ	;�]Ȓ7�E����U��t\�!8�.�r=#��/�,�n'�㓐�d��'�Q�T�a#Ƽ�5�F�{���p�|Ȃ��1���QD3;���x�����'��S���?û�v�e1�^W��:q󽮦���Xh�o�m���41��Շ/���Xd�M<�Db�u�1N���1]�M2M��hpR�v��e�I߀�|1�.8�x^F{�l����**���,��F�����4Ǫ���	r;������`d
�3��QʟD(���5e�|6��_Agg{�^\�ڭTtB����*���H���JƗ��Z�������=,7�s���� � v�\��s�U=TV��7֪�z�gv������>���	V6E�l阼2�H8[3S�Yވ'n�wƩ����|����^v'fI�铧����D|���������vFOeD���9��D��qz�x�c��1��w��M��[���k��gӞYVv���*,���'��������~���k_7L�|}�ר\e�]x��qA���{�;�����P�NZSk�xj�Y��lG���ۭ�����Z�t���q0��Yj)-b��TYEJ1V�a�Ӑ�Y��F[QT��ʬm�!���ṴĆ~�~���7�����=��01�X9Hٕ��+\��o+�o���pNc5[�uv�\rq�h���y���b�y�9j5c�4�QHȺ��}}�Py!������*7���nMmo[�M�4:�q�ЎRT�4�w�?E�^��{�=��/w���^�;�޵�Y�˟q*-/C���w��q������b$�}���z��U6�1C�����r]7�g�a�R>�IE����G�لZJW<�}��COIŪ6v��Df��Z5Q�D�dzqG�V|~'�Ű��,~�D'ڟm(�Y1���A�	3�:� �W���}Q^=��-��$f�dhڛIk:�WM�xWi�C��6¦��mt\�����ă'&ǈ �	��D����LVz�M+|S�L,A�g��H�^���vJ�\�ݱ�e��*"�3��f�/2�ܕ�{׏�o/⟀}��k�Y\֯���H]�P����0�J[��p6��:ٻj��?������\�i 8~�*�O9sU���$�%�5�k��*Q\7H�t����!���R�u��ʗ��D�F�2�]��:3=���v�H�[���s�+�zA}�Ö�z:E�y�)��~���>y�r)B��hG:\������-���n殱�w� 
b���3����f
Jy��Nl�,�';���&��Ve=�6H����celTC���1�%?/�����Z����`�m�=�w?s1�1=s��Z�Q
$N���KuZ��t.Qc���K�e��I��<~�A���������{?d��"h{�� +3����Bgt���}a��v����g|�g�$�{[T�m����o�?}o=�Lu���o<���O���'�S�P&�ftX"Z���#g��_\��E�o��aE��_ذ��ȇ[5����_p���}��}�9��s��:�١�����ɣc�C{�u|xI�G�ޥ�}J�(����~�_���g�����\�q�'�#	$�;��U�k�z�0?ou��L�:ؼ��*��˖E�.�_kܯ;��|y��:�V�:�e�%N�D˩3.n��0ԛ�t�f���v�>�Evv^��T��k�S�n��ޤ�ɉ�L�o`�J���1��΍�������Q�e*^����Gr��C��G�D0{v�q{&,��K��Z;^���Ng��@�;˒i>��kN\m����ݭpD�g���3��G >s2��4��;;��{�O��wy�Fzf�`�+�ć�l���(��+[��&���ǌ3p�u/)2�s��g�����}]a>o�1j�W���wL�R��_WO�wj:3W4��,���3H�Q�nA3����/�5�G&z��;���5{�p�����a�����67���uG��^�;�5r U���S}��q؃,��>��y�p�]D�����|8݂�:�;�[�* #�}���<�c�6��C��{�����ٴ�i)oP/rN�L�-C|����@qz�����e;w��^��[C)L����rٍ[!R"*!YD�l��ڍ4�b�i`e+w���\��P4n�qhR��|��N�V���y\��"�$�й�C]���5��ҟS�v�c��h=W]t��Y����h�����^����{��	4�w��&c.�O����dz~�V�yWm��/߅���r*$�@�~�Ŀ{a�!J��/1G�
� P>��lJ:�ǆЏ{K�1&4b�q�e(��m=���Toj��C��/��@b�d��j,e>k����Z�n�r�~���GAu�@�FP����B�W=W�a9c&'`�(a���NʼH���"�/�'nrxS�6���z.fk�{����=R}����Xм�w�ҮC����:a�u�3|��@k�^�[�NV,<�DB����������t�9x���tH�1
@���J}���O���ε׆� �A����t�jy�7�f��i�Xr�f��'2j�$c>�XV�\�nt�G!K?|'=��|�Ֆ��]]X��7�1h�Z�������NMݶ8����ߎ�OM�Q��:�
[ HbI"(�2���}Ϲ��W˳\������.�`1(ݎb^�����k:��YĶ�\���v�{V���:�_Ml��J�Ǳ��t��˝��f���-���n����n#�z(�8���\��K��\����@����N���wnB���,���އ+��=	s�ӏi�&u~��Wq`�Oy)��d@J�|v�����+G[�ӷ��M�.�ՙ��\����Ώ:�2W7���y��9�_�a=S$4����>�����4r���ĒD�9��x��j��Q�A�>\D�9<M�q��9�Fk�4*�\���P��U�����	�ڠ|2����ߕ~�:�׼�9��{���ٷ��p������Ha�t"����	�x�ϭק����y��K��nNer�+Չ2!�갶�G�ߑ��o��_�����O��<E�E=kBƳ�f��YK�#ibg�OL�",��o��f;T���T>��(w-4��3w��|��:�6m���~��>)8ASVSQ�(L�4�\�D!@�
�[V�,XH���3fd�`
1�Z�H�"a$�bL �&[������7Pxl[K�g�Z�Z��S���
vf��e0��2p#�Cy�a�}#}�"W�ݷ]��&wihK12���n�Cy�6p�9d����N�]�s~ʌW\t�,xw��}�خ`��晎��6�}�?u8V��ď��zJ����/�y�������1�.ޢ�彚�R��}K�0l��F�°B�[<���v�T���Ztk�l��n�-n�׾�<���}�w�^RR
����_U	ACQ�o�%����gЇJ�zfLE�����L�7�#�5����)@u�B}��w�n���?{���7���#ixY��_���Ҷ2E����}�A�դm�p�.�^�8�Ω�T���(���8��e��ۅ��Y��uۊ��<;ޑ���}��-�eE���^�N.Әe�6\��!����kD� �e��I��o����p�9�V�e��N�ď�>Ro#�T�*��C��[�����.{)�\K�����2P�^yG�zTl�3
�-�t�&13$�H��i.��u�ti�"�U���P?���l%{=��xyO�鱔w�!�@��T�@�Ɖ]�s{����t�2��&8S��]Yԍ�-t�Y����p!I�˸�j��yY���e�����6� ���^����	J��NʪZ�.L���&�F���%�H�F��ݜެW|BІqgTԳ��P�A;����'$;~�ዻ�ڠ_��/�).����HHrr�`^k�(nd:�7?:Md66�Z5t7R'���I��Zc7gIQ3۱~Ͼ��0��&��߽��jP�=ͦ�Q��ځ�����@�5� ���"#H�]�_]���}���1��b���KB�q�f�~����M�|Ͼ?i�$eW^�b�K�d|���Lؓa´���"yܮ+�������y�����G�۷���.�;�����@> q���KFl��	+z(�>2Y�{�r���^j��f*w���>��G���:G��i�m��]C~�B�����j�}�~�s3�c�O�����)TU��(�I�7-�ٿ���Y�1
���.�a2��V�5T�f��)��V����n�V���;�8�Va�T7P޺�+X�d���+�g)��l���2S{�O o��Z�B!�3���ڗq2���y�3#�p�y�I$ϾϷ�����x���8뷍c�kJ�O~��6�P�Nۂ��&N���E�/QŐ��yߏq=����f���X2@ ��{��{��Z��A��k"�4�3�	i҆]V%�eȊ)��^��H����[U��y.�����˩��3���W� �mx}�}�^J�G�z/�~�!#��Vo�*����%�ސ��T�m@�*7
����R�쏩�Ӣr@�ͱ�c�-f����bSJ{�� ��50���	���ݨ�B�6z+t����ˈ4^Ku:���|O��>$�lϧ��""J�A�6Dpk62;�V���K��p칉CZ��	`�Xj�Q��I�^{G���O�1p��uE����*ME�(Y��H ��VG;�n-��,5�QN6"����`�#M6s��7��Aq�lZ���> �^wf�Q�~�+�0v����P��[Qg��_��`
�8��ukXO��U���]�m;;�5I�5�[o]Vf]�_�K�.oO�f�i
l�B���h]��&�#�8f4%Zb���[f��f��:�#at-s��K�� ֬hV���4I�j�M\�g_mث� S�bf��O� �u��^�D�:�8:˃�<���������F'��,���1�M5t`3�z��Ufo(�\�[��,5�o�d(\���}�����.�����_e��DB�	1D�[r�7�i�"ZQE[�h�.�5�љ�b]�f�e�$��'Vn�)ҨVnT4h�����c�Dm ?>kޖ���Õ\��v�u^�Ǽʹ��u������CFu��V*�F����XtܭI��߻؇w�_;�s�N#Q曇J(ŭ�\��{�~yC.R�ww{i��]�NB�2ҋ�ZњCt����,���e�N&e�;��Cc�Qj�K�޳V,��tѷ�f��N�f�OoP����LK���|�[J�^�*D�W�Yt�WYx{�S��u==$��m�ےn5�/q�ݻǋG^�����"��ϱTΏ�H�fݢ�c�\��7y���j����z$�/$��<#o�-�;��FN�׵��`JT�8����P����]�}�d+��p���<�Ts��I�����+����4+.��DyL�c��Vv��țrn�&Z9�����փ�T�G
���Pd ��ʵ ;ȍ�(t�4���IcW��(%�x�3-XD6��Vm\ӕ�4��3֮��T�uj����-6�ޞ�k�\4��TV�X�e]��K��J�*���-t�Q�-#�e`�ҳ G��7N��f0����Q��?���n���lU�3Vu+Mg5N:��s�Y��x�Cw���.����Y|��8�q�R�nө�2�1���'�ի��9���twY`��̐{'^�.x��v&�$Е' 4��<H�6�!�;�rڸY�/p1x�J�����;���@e�N�>V��pˏ�f���%�X�Q8�Ŭ�(s-;2���n�	|�fQu�&c�Ģ̽�9.<��~���|�\,�y0�nP .�]`�P{z^�,{+q'Y�qҁb�n���r��:��nu�Os�RP��� ���K�J���k�Zi�ST��ĵ��7`���dS�1��L���rY��q
P��ڰ��ml;w�.�Ñs�Q�jlo2�.��9���� ��Wq�6&4�BTqz��!��N�C&X��|�u����X�n�
���A "��]���%/��੏�@w�f�uښ:�+e��;�	\rX��� �o�s����!�AA]\jN�����WОQ��/��Z��Ώ�rxP�c|�/-�Ǝ�^y����q�O�s믿L����}ퟏg�9Ku�M��1�U��f����nn���!nx����d�ytw��@7ʵ�'�Qt^�A�Y��\�}.H��/��HL�gU������m��k��}��&	޸��/���=���Y\oyx'k8͈3���ü̐	��y�_�c��g�ߤ�� uoH���0;ٚ�=�����v�m]�Ǧ
��n��λkԙ�c{$5�Zf�C󶩋�y#��:����Շ�O��������R���K�Lb)\'�.'�DP�w����[�.�Y�#����Fw�r�u��%���H^��( w�c��ߥ�t��3�\~�a>~�8��}󙎵cz�B7ગ������g�ш�W������h��f�!X2�F��P�����}͔�,�!�yg1n��hq�s��*��z�BS7�x�t�K͸sO+O��4�Ʈ�R �۵I���k��:��p7a��e�
�b�����7������9���o��rױu/�����f�i��x��C} �R�Ω���a2y.f���ڗ�Q�>��v%�v2c�	`}"t���!\V��|���h20n#~-��+�;�b\N5N���0z�Gb<��0֕���<�D�N�(�����g1�|�����K�����əϕ|�Eyne�f�q�B:��g$�f;!朷�;Q`y~p*U9t�MC���mO��uU���  o��j�s(z�9�TYѩl8A��� �N2n��k��sF�EQ���`lZ��J.���''f\B�?=(_8
���\�n��W�s���Ww��5��ʥ]�$�1���i�`㛉�ӷ��y�l�~��ªc�<�CƊ8mVKɋ�
����4xC����7�e9M�uǯ��i���G��Q�d�c ���*1H�-��eZ1��T	D`��J�`[ D!)��*T� 	 $+X�(Q%d�/���7�w���9�.�:�i�;�'����b;�X�ц��屪X���_\�LPe<<�e���ZVD�n�NZ9)��,oq΢T�(fA[}�����NЎ�����h9\(!f)Y�S��t�Vd|�	�۝�˓qtzG����:VlE�=5��>�	5<��A㵞�jjiE -��7�}�K�&�ذXȩi+}ZدC����U��(.��$��!���|��{���7{�y�����,�
����F�IF���ڏR��Ñ��s��cظL��t.�^�d��u��K﷌Y�OM����0�S��e�s�7�	�]5��>P1x+��^r,�Ώ%}nr��.��Ox"uAx�K=�WR�]x}��{��+I�?|sH֣���Yѽ�G����,U��{T�{Rd��N���ͨ!�si�Z���� 	����n2$��e�d<�3���$Ji~�^<�[��#j����dږ���ݶ{5kׇv]�����^P�\�j~.�5����hK�B�O=۾����ł�U��E�k�z��w�1�y���<��|C�EC�����f%Q�Z7)�����K����F���y[��.�
�ǄX��1F�!���X̏��&Q��f*p��~�R����ɟG\lM����b��rόT�L|�7޿E��*GiZu����*��6�E6Wc����`#�w���˴�LoQ��ތZ�2�<4���e�F�����")N�D�D�ܳ-��0}�f{������<���}���6��HL�z�9�a~9��ԃ������\�~�Wu	~�(��Z�>�u&��k��
ާ�T��q�"�J&e����cr���Ƿ�>�Y��H���s=0:A.���:�Z���Q�c�B-F۝j�q���'�>m�Q��w�R����	��ܾ���s�
ʼ����PgECDa�Y3g}�GαT�
���U�������q�\Q�Wߡ��U�>�i�U��+��:^!,?Q����#�B��lsaR����:ˏ������2��F���`�f#TG�Q+�YP�P�]��el��]�9��y�h���\��(j�-6.�"�i���+WUヷo`�U��'j&��͗���M�<�$I���kl�5�ܥ����c�uweW\�{��>?C?y$���\nS��g���Ә{U��toY����kQk-�>d�f�o�:�Z@��>���팞��Nm[@^*����?W���߷��ř�X�ť�H��cb�����RN�;��[�y[\N8gL̛,�R�w���1��Bm��+�&=�頺Wx�?\3�X�_z�{�5�����\8q��i�4���(�6����8gɚ'�A� E������{������P�c	���Ʒ4��]�ؚ�W&��U���mM�W�%k
F��LJNs����'B�þ6�y����@��[�y篙z�w�in�0���sa�����x���R`����i���\_V�L��+�%[�up����d� �3���|o�o_��W��?s�>^�����3V�]�(�"H�X�B�W9���������5�߼�aTWٹsd�,t�m��W[+��]�;}���qS��m�=Q�crN�8>�x���͹ػQ���z�H�徙�ȗ;X;��3m�g��dC�I����E-9��ꁸ� C]�t:��@�Z��+���j�!gNMC�k| �T���汫��ߵ�ƝJg)�-Q��9��WPER�k��X9Z]����O"��L�n)�NE%��@�c��X���ae�ӓ7U��Aqcby���H����ǋ�Z+�2H7�``��#5~���yY���;
 P~�z}�X�t���3��q�M��������04Y�Xb�o���^�E^^s�U�/ ��Zb1�=��_���f�>��=(d�A];r���w^�g9A�.�D�W�j�QK�-?A���G>�D��5.gT�nB�V�R�k"����:����D�xK;�bl���[uW�!�xl.�
}�ˆ�����x���u{9mg. �����.*��c>_>D�
H��eR�FHE�G�|c��@E�N���[�i[�۷�lt����L�;;�����t�5(���Ḻ��+�u;܄	|���޻ف�gwY�8��q�"\�"s�f/_�i��#mms��6c��w��u^�3�kaвT�%!g��A�n��aJZ�� A�Y��|>ۿ+'�cϳ=bB�3 2%���Y�Ĩ@�\�EN�j�T^�=A��z��'i"�'Ȫ����{�P�C��tX� C�?{��*w�{�����G5ޱ��l-$#�b��{=R9|�kOl�"��f��;���U���0v���ާ��0��Q�Vģ8��L z��vdޟ�8�3����h�cs>����,���5#�2�e̺`���ӛ+�*�mJL=���*7U��ޤ��
S)��3���*�9	�����@��'T�vS�c̽�W��n�N�ܻ����WY��y�o��hp���~&BI>x���/=����.���E	]~����=���~��'��)ik���6�E�9��kY�ʨE�$F��ŕQ-
Z���RU�"Œ(�&�T3[w��E��gi�<�>�W& �f�*W���V�&�t���,iǚ�"{'K%�����J�R���u_U�Z��*�0�(��36��Te�WV��,�S�w��n�WO���t�˗��}^��zB��s���z��!\Ⱦ|f�d�[ӧ�qb�#���r�j`e�cu/|��e*ȁe�ޅR[�Ʌ��>|�6�B9��ʱ]w�����t
]�^{'�L^��n)},��>�q�
Ѻ��:KW[�Z�m?�0a�����/�Z�|v�v��zo�}
D�g�Ժ�xz�/��V��+�)�lT\$@����>��i��(���Dn[�I>�7��w�K�3D�k1_�7,������� 	^��{4C�NM���{�v�h숱����k3L0eymލ#k�te�[�v�q��?�����ߞ��:0�y�3+n���JȈb�~���w���{�=�-�;��;y #L�5[�P3�c�������j���]�S�4�@�m3g8ԛ6�D�Y��Vw�@i��w��9�v�gv��٧2�jP��xH�t�wڞ>f<~|~? ݑ=�Π��������9W��{3�Ы��#[.+�"��s~�v{�*��1&ffzw��c�J*;`��X�蝍�f}�FpM�/�ݢr~� �E��ʌ��SQ��/�F�v�x�Z���B ������3���y`�g~��pksC�J����
n�^OM_׷��2��D	g:=��������ǣ��Qņ<ZA���El��T-�Lz�_�gO���w�w��l�����s7�B������5��������I	�o���>�SQf�΢�e�w*�˾ߚ�<�;�{�LVk��>2˓2)\�["��+Tث&������he@�s�t�ӫ�rw_M�Ф�ٺ�Ӯ7T�������n.т��__u�잽���:�̖٧3��x<;��W)W>�A�p{�����]�!�ɡ�y���y�n+6a��χ���ݾG���]$)_�'��8��~���P��'��V��5 �f3����l�e�(�!�������\T��xԘSq<Oz��G�z��N}�P�r3�{�ul��XQ��Tk�������=��F�KUIL�!O}�Rt;��g=�z�2������qzb,c��F���T��2�ȍ�C�7:<9C����	Ρ�=gf��v���+u�~g�p����c���܁�\�[x[����������x��%�jD�wc���گ-�n�q@-�a�j�T!���d�����:��V��>��}�st�|�7�s��uu�k~p�@�$������y��6o��2u����]��є&�����J�Vx����������N���PĮ��]�e Sp���YXvG��e8�.�P�J!���Xb���}L`����Ri�(r���U�약O	+Z8"1b�\]Vt�#6	 �@�s�( Tg2y�-�W�:�)c5����s5�{��V�fZ�y�Ul�T���_�`��q���� E�j#O0��q՚�
��3U�ڂn�I,J�����W���3��Χ0�hP�H���Q�ʲg����cە�޽� �7�[y��q�a5�)�h@E/�&�7��vc�%��0�s��2��$�v��T8����&2Jit���s��Ԫ;���F�{�[)�N i�{���/��1v�a��{�ً�j�cݶ�[U�J+YD��X����t���x�ԭr�� �'�4��=�jl�t��(��{�w�uV�o��	ċU6&��ֽ^r�ͻ��uH
AǾs�@�i�4��@�6�����]�����u�2�M��y��Ws��6���I��n�pC:���`;{u�t���v=Tu5�3�MI�?N�W�vgB�&��VwuI|E�<!�EI�kD+/������ku���j9�r�:>Úｌ;���sl�뀷���]�{�N6K�Z]	lb��`J3��kK�	C�o^�z�p��0�U��%���6_8�ç������}7ۓ�:H�Ѭ�ܴ��vsx�|�Y2�uoY�jo&Er���ל�F�6��ӵ��]����C�i
��gsܦ:=]7��[�\Zp��2�uJ�9knB���R�w�eJ��3�)��c;�琎�t�{�A��6����)��[�һY%�	���Sw|s�u3S2�I#c�*�˳o[;�ٙ��SO8�˓�0���
M��5��%����e��wN�4*��1/�V4\�% �T�2�
���6x�:>�P�8}�9S7�j|[B���e?�ٸ��Yk���H���)�R�0Y��x�̕�mNz&���o��n��@���� n��#�t���$@ᦠŕ�Sఙk�w^�6����[C/.�]8��[�jf��Dפl��=g���v�+��q�x�&���α��&YV%ы?���d�n]ͫU6�����c�ue�
,���G�!V��.��53J&�GS�u�L��+zr�W ��!�B.ܺw�>W;a���UwzO9�VJ�a�u��y�b�E(zsaKi�}܊���+����y��ٙ5�+?�ͷ9ڦGk�Ei댥�;GQ���;m��J�v��uj�q~����R��8�X���N0>�|���%ʰ�\Zjt�B��Yc�3>���n9*"){O_i��r�y׻�I>����Q��b��
��;�C��+z�>��Pvz�(�B�d���[>!i�K�g�6y����^ȥ��ѻԧ]�N�����������R�R�jV���h��7���t{z����>���/��V��(o�\*�v�<�����ݽ`e��;)-1z�FL�]c	̟��tt@xd;J��پ}6��oۦ|I��Z�w��*Pb��;A^�z��⿷�Z���UR����$�;�"��v�X630D�L�SX��*�%�����m���!a�=�6��[�R�TH�EPGWV���Esn����`��X(��Q���֩kTA3+�ժ%�-U�b��()
"ۅ�TTZ�,�XԪ'�|��OU����;��V��A����g
s;C�ҧ��/.�.�L9c�uԺ�qG���BoS�ξ���T駞��)P��[� gG��̦r�{��U��gU��K[;�F�$��.���g��^��3�5ﰶ�7ד4ڻ�ދ�;�MW�ޫ|�|�'Y�>�#7��VL5f]��eٟ�|27�E�����Ѿ{x,bʈ�;�>����=L����w>�
��qtn���WQEy�2���  sV�<�����ѫ�QWR1�$��m��D:k���qƶ֢{~^au�t��n�g����W�7inM��A�]��n�5�T���p�t�ޤ�ME{އ�G�_^f����Q�V^�����7�ca���̗f����|L�&T@��H��1S1Cz�S������斚Zs��Mu:7�h-�QJ���.������<{��,��\����K�V��E�[�#ױg(K�D��zTD��]���n*G���(���.�C��}�.�x,�{	�X4wkNYG���i�j�4�پR�o��+&Lש��w1\>Xբuu�|�ǇJ�A��s�w���Ӯjxw����  QB*� O6$93� K����Ǹ�WN����T�t����_T��>����}u�t߰����&g��Q9�*�؄�n��dV���w]�ݛ˝�X��#�ݵ�sj��,��A����������nة7�a���z7YG��J���;8�p��7�$��%+����c��w���ٛ��[�{B��|I�#��0�[p��DPPRf���UO���§���A����B*�y1ջ2u��hբu���,�wf+������u:=�Z�z���.��K�t#���;��j��5�}�jn�[�~By�A��e�nc�k�D'�#���G�9]!��ϝ�vV�'�Jgg�w+:���b��2�15Z)了K=�M�Yy����U�_�%^�▯�;�����4}���[lt�򂖅�}�g0�U��'�c���꺪�yixW�����`���B�,/Fƾٸ}�ո������'Xۨ祙�{����ޅGr!�X>ɯ��@��9��1�<�j����8�ǹKY�V�pi���NsM�j0]�� ��y%R�,�X�\퓞S8;�u���[8�����/xG]���g/�%ש��NgJ���y�����_���ld]���V�1���R�X2����)��p��ے�'����^.�c��5�f����t�NYS�_'��Uy��Fh�=Ӄ���R48a����cצ�*ܓ�g��]DgFc��q��٫�rY���_PN����rE�"�P+e�u��p���!�������h���yX��Ot�"}.�w�{p������L����Q4T�w�߬|�]W�3�![���g\��\_��QY���Yf*�f+�|}��S��M���jb� �Z�`��T�&��c��œ�l�9D���>�._���`Ê�k�E�/f��߷�ͩ��{��tR}�|<F�2v �}�C+ِs�_�-�J������ڹ�8,�^2F��� s}���J�=|.=>��>���
����Y3���2P}��:j�6w�M��q2�}a�W-�p�IK<��sQ���{������i��7���W7,����U�B��[�L��f>g"Ӝ���^��6�.��˶��˥Q�yz9�0�u�6ٮ�ڵ�eN��.
�M�	��o]E˃l}n�[�s��:7;��Q�Q�u��
�y(���D�=j��8�gd��/cٽ��r�T���o:ڋ�>����.!�C�ﾎGrv{ 9���'6�R�ÿw������� �}Ӳ䅕)k����IM�U�rl�&���:��-�d=)�_V�����c�}3�2�U�Z�<�kj����Qc��_>�6E�j~t�V�����uM�b����b�M�N��4��ޙ�ʡ�C����vɢ0�E5�ʶ��W=~O���^���in��[v��mٽ��T���}��=��O���U�!D �Nf~ %��Ye�a�kN�R��e*r�����h�#)���QV5�f�匬�m�KE��."An^�����kp��̨��ߊ���3����b�7,ԙXG��y(T����Ō�o��u�>�7��}��j�JNED�^�ơ`4����.��-ug�o�x�Ɣy�3�i~'���3���}>�>��8��@��&е�s�sc2������=Ӱ��1ILf�ǞkcB�{�Q1��)PK̳9�H�.]3�����/{).�n��/��O�������26�<�@}�خ�g���W�?���s��vM{ҍ(nu��fo;3:x���]g9O��[���u0>Z�8�~�{�ϲT靫|.#2�щ�ҝL�=�m��|W׈�u}L��^
����F�n������_�GV�|\��ޤZTn�q�ls���Ikݾ��/���o]���s�e!l�r㤣������d�*���Ly��Tq�����I�H�b��n�ۋ��v�B��%�X�mHmgNʂ@w� 
�֍�:�^�������Q��Yk�q)^������]P���@�/�N� �^���˷W��i_gTeQA����9Ө��Z�ofN���|J��;��I��"������%Ա<n]�ɑw,���T��w�^�i�|�!� �u1�5�j#H�����{s�2y�����)��}�g/�C��	9��N����]st���������"ЪTS�\�ay}B�f����rz�q��u�;�¾˥�2onB����(�g�~y@�ﴳ���I�u�1���$k�^f��E���4'�8���-�G�|�d�dd�d>�h}�A�,�^M8~��w��SVsg��'���� ~
�!��nQ����1���Q盃x�m���M3<�w��,���dtu˒8:���cb�뤜dpc���P?������fo�t��3Y�����2o�إ��"��| �����*�VT�yÌW�C�}&�rW��qKh�gC|;�U�ڴC�ʃ�<P"�/S����<ȫ�R�;»�ݮ��XvL����%v4{P�ᧅ׶����O,\���
]�ק�� ��M�F�c{u}X���\~�V0��Q�b4�)_����c-27�Ր�ż}����ǔxW��G�Bn�f乺:�u�z��S�o�?wysfF�Qυ�+ιڎF	���7���=���R�gG�}��b��,ElףMѵϩ�U�}�����H;1�œ����m���[�:���}<��<�Æ��h���=���kZq�]kCHi�Bb��"�mc"�)�G�>ߙ�9h�̫XXءde�*=�62�/_ &�w7ke���[�;P���}W���6���ӵ�,����K�9�ۓ@:QM���9�&B���N��o����}��9����������D���I�7Wپ!V_k�FH�i�s��f��W�z"�*��;b�7�긣�ͮ���s���KbS�x1ίz�r=��;��V4j^�]�S�/�f���}#��-�݇{�eb�Y�e�Bٜ0��_��%_�W2f�v�?}����u�v��~�UW�֨0��>���_��xl^_����S}VEY�x2'�x��Ĝ�����}���$$a����~Q����2��9��FM�X�d�;���"��: U=gy�q��E�3�U�q:���qW��^��ƞ�u;>]�Z�↹$��fT��B��L!�q*�bub7+]ks-.foY��t��YHһw~2���.WL~���׊���;�fD���ژ�0�k�u��U���,�)c�U���5�D��zk��ˆV&�Ͱ_�PK]߸c%���m��si�]*�c�q�(���s~J��6����¹d�e�
W� �	ݾ���[�� ��9�w�S����%6������z� j�쯺3)to��o��;����Y.�c<d* ��4Sh��WR���f�s7�\A)J�Z-��c+Q�W2��7R�𦹽��9f��3�+��d�q� �to�P��H��*�9�1�r����1��7��<����S)��qqy� *�ʥX?4	�Ghf���3{|ü�=:���~��)G�.�����<���ͪM�̦�ֹ�o��5����
����B.����Ҝ�Z��^��o�pz�o]�����et���/����3�&�j�*z^&����-���]��.�ΗWa��#ZO{�DH9@�Pohp�7��!6�#���"�,���Y-\�Y�i4MZ]"��P���4�LL����.Xj�bl�̦�5I����<�N���W���VF͗�i�nF��H�}v.3��	�N��l�L\��OjO��J;�.(�΋r�-�OC�+�(o'�Y7��]L�P�'�<��t=�A[BSu���7�OF��fv`iks������\�o-u���wG�;�s(�|�ݝ:
s��/iix�`O�pe��x�)�dnݧ��7��:kYw��u���G�mct�ݤ����h��Y3v&�`�ViE��{N_&��¥�yr�
Y|oh���y���èS��vk��]r�k�^���V��65M��3m�6�㇆�!�,�`�*��V����nf�҂�)����#]�F�{]���v��Wta�1�� P�A�[
���&<�Uuw����mS��vUպS�9�jo�[`�\�i����!��7mŮ�uh4u�L�K�#�N�Y�M��4�{��G//��Ei���uK��
���t[XTmţeLsY����X
�%&��#���w.[n�ssA����`�=)]�@Y���c����v��i��;���X�^{w�r¡�����ڕhT�E�k2f��Ms�x���٣*���>U�J}�6tP�G1��u��I�⦕(;��Z�+|��V��#�DѼ�fD��N�n<e���Vڻ�Rƀʻm�m���|���X"�L`/���B�c|[l-D��h_��s6���a�����q�$���Y���f)�c�q���v-𺘃�w؞����o�{�"�}��]ϡJ�$�f����!�50�xö&em6�uևb�*\�."�ͩbUﺷ�l�U��|�W1��:=}�I�4ȇ9�w6��,~_r�Gl���|g#b����f��>�#�ZeGe��s�8zk�Ӱ�uD2.Y>�v+M�W����C׽��<��3�Wu��<�n�UKVi�ɱz~�["��R<dh/sD��3�j�t_SmuTgc˹�z�<�͆�Yd������Q��ߔ�A���q��}�G���+�~>�c7B'lf����z��l]k��u����	��<.d���������Ҷ	�?���i������E��,q܊6+=��sx�	x�B7��޵�x}F�C}s=nŞ��`�G�&W�AF�6���;���7���Vn3'�a5�-r����MC-�c��HB��Xń`K�hc#�@��H�`̶KTZ��B+`�R9�  ��~'�E���'n�dݖ�Y�Y��l�j�G�.%fL�i��)հb.�k`�E��4��黉˽�oz��$��k���ڒ�7N�s�R����r��N�+���o׽�v�v>�Z���Vpެ�+�b{�LA�pR;v=G�0��݅���
���!��(n>����
��u�>��;�_������cs/3�N���f���e�۳[�;"�S�3W�٪���կPGg�1�oBs�����m��M߆��WZ�6�^�r��|w�sL(�*Dc�v\�;��%ڔ�>��~b>ڰ�}y�+>k�����^�NP�~�w�Pt���><J]��W�S�؝>�5���������x�ɑ���Ǖ��+�*�uԞ}��1s���^�ޕ�׹�k�K��|��Y �x�P$�@�g)�M7Q�Sw���3�����"��x��V��ךO�=�;����fc�R:9Eˬ��o��U��u���,gfq�e�=���p��"��q���#�w[�۸b�Weo>Ebrr�g+��J2z������/�q�Kh�ߣ�V�F�M9��}�&�K{}u��l�<��$�r��y]��}%�/2�T�n1bl}����q��;�r�9�t��=v{W��)��C�����&��À ڛ֠�p����A���>�P��=Ӆ��O��_��h4~J������=B���-ե�����M���W�88�E��n��U��u��p'���"�e�ܶ�]g���yS\�.1c�\{s�ǽs�����}����R}���C����gԊ�N�̣��~��<��Z���<��8	*��\,32J�XVVE�5�w�1:>zy���w���yRuJv���ڍ�};��]N���6�	�PN C����Ou8FV���e�r$�G��.��.�2���l����"'%�MG���[̗RO�-��	�ڧ�|4��@�W����P��ٛ�]�G�{k��2W�ՏK��՞�����Xx;֠!T�AQ0}��;W���q\����Zˋx�� O.�`\����U��p�X�D�������������* �VNȩ�v�&yc��ˍZx��*�'���eʊ�|��N,��S�^��g�w-�}Ҙ�u��N�ykZ��]�7�p���	��& }���l���Ug�	�����Z�������v��lU�^�IV.l:���6>\
�š��X�������m���L/���\��K_M��|��s���$��Y���8WN����
=Q3v�1y�K��,A���8�jg�/�Z1.憷��f�N-�l־B]�������Qxց��~�K��
�(��(�4��%�����T�uc�s�55�ϢaF��d������-cNҳ������(K�r� �O��L���:�2G����������/�e�hb΋���5Lq<u�a�-uA��^�r}���ꪐyg2��&]F�����J�`̲/fO;�	�=��xm�P��V����}�J�z
.ϟ� |�=�'/i���7����~��?<]�����N�K¯ה������f�QR:�薸�|��p��f��g	��<�nT��Xq��,�}E��:�Y�י����w�]�C�A?pJ"�h(���0D�T@Y"��P>����ﯼ�St5m�j���
ز^g�\�f�ur�&�{;�����qu[�J%ZrF*GV�_T�|��_\悁5����U�H��<����t�4�%����T�v𘽧O���Vz]�iI?~��kު�߹?1>
7SS�c��?u��Ŋ�Kj�vz`e��p���o���y�y�~V�몯V��*�;RB�z�:4����ٵL:�w%�i����Z"�v����{�� �������� ��"�eh��p�ql��[a�IZ�Q���Fr4c<�� �>�o��u#9��@rL(uR���o�e+�����k��Ev���rd���+���G+�
O�v�&���� v;�9�Բ�S�����vU�5�q:uî�-:W\y��W��i���R"�0�T��(E�@B��!+ V$���淽������v����f�txc��:�޽��s-+|�ú�)llC��y��-��壠��v��3��8�[S;��ʋB��R��ٖ�	ʺJ����t���(��ՙ>TFP�l����+(ؿ�s�c�Js_�*m��ܘ��xD���}>���{ (��5�s�n�
�����I��.����u����v��XQ�L�o.�Z�ڞ�yԪW�gɬ������l(ʣ�Mҡ)��f����/k9���\k4����
�gT����}��{��P:ѽ�\��w��`L�[d.���a�n�2���9�WX�|v���[[��c���m2�ʘ4�GT=��4�F�uE�C���Ǻ��wV.�p�Ɉ�b�9�+��Hwݴէ٩��k�y�-���b�>��v�rTK����dg06��]�"��)ȭ��O!i��'��Q�+�q4�_b�Ӳ*jc�e.V��9�ka��*t��=�a�\��K�Ĕ5êt�:w�--��
���x7ϛ[�3��ZA�Wu�du� U��^�\�����&s�9��#�a4���K��z���(�I`��QϱY82�C�H5�cz�U���g1��h]��0���ͷ</+5ebQċ��=�o�'��Z׌	Ϗm3Y����h&5f�t��W	Ŏx���+�3^ʫu|lj�u>ێ������]�ǿ�ϴ>>y�����I��z�}O��_F�N�"xpO�	Q���n�*gT:���Q÷z��H�~��yó�=�qS)k����Kp)�}���t3�쀻,���@�Ϋ쒯�{���e`a�y�0.�I�Q�1�R"CI
:5��{�ם�|�]�����U���gWӞk<V8]k6���{޴z-t�ˎ�w�B�4ܽ��}5��\�f�i�o�${��_^�h��Cؽ��y��^;�k.�{�k��'c��͡�M	�vZط9��4�㦴Uh`���tě��.�SO���:�e���z��v��+LB}wQ4w2��V��������sm,G�s<�}7�[R-u,������2^�}�N�F�ۙ[վ6h%�g���8�����]�^���O{��ۺqwdkw`�a�|�}E�w�P�����C��KIJ}�����q9#YA������n���BKqw��e�yM�ޭ�zc��ī������>���^�]��f�f��_�r��k[�}��>�]w�7˟h,�/K/��U�d� �A`� �W<�z��wқ���8_J\���#�|s�oc=ӲI
�۫�4�9��^�~u;mI�I��-�֞���T�([Tm��&+���T�2���~�o'��7~B0�c��J;���9����#^ߩ��_}�.F]�|L�dW����~�ȋ��M**��mE��ө����m^�k���}������<��Ž1�d�%���L�d�D5��:D�b��s�H��w(�v�a
Pݴ���s���$���=�3G' �R1�/Gt��4�¯`E�>u�'x7u|���r�u���$΃|�ﾽ�x�U�k���!;��W)q�\��lŔ��oִ�+�����=b�p w�����{B�T>X�c�Θ÷�8��u��M�eHZip�J_;���*������;x���+W]^ڰh����ԿƢy�GR���W��mT���ny���,�[����"����������HI��d I?��T$
��HI!�!I	�H1��	$	�$ ��� E_������@W��W���l�yx�� ���������u��p�U�Xq�8�G�lĨ���]����m�*�N��W5�y��T�P�e�MœmD�����p���\��-�#�)��B���m���9�	�;U�.���81��L{{R)c5btU���jmV�,YFDԄ�L@��Srw�l$[N.���@ł6��Z�M��M�rC��@��x	Ǜj;J�����bM`��Mh�(K6.:�OB]�	+�0�t��  ک@ԥ�l P7 �q(ҧ�Z��X��	Lwn�)�V�;�e�X��h��������m`������_�I #`I  #!$�$$����$����� !��@ �@��!K�����"�"����}�(*�X��������3�*�PU��� ���b E^���~s�Ld��@W�
 ��!�|�}� E^v;�G��\���"��]�~�(*��� E]v��1AY&SYyu��߀pP��  � 7'�`a��{��V���h	��Jٵ���H�,-E�,�HT�EL��,�B[�� m���[Zk5@J��%����AR��Tح� �P���*J�������U
� �Zb�Z2�PJ�����YR*��U-����P�Z�RImYYjH�,�m��mf[5LmU&�kcX6�4����N�H�G3m�5VI��͵%�L�͚��͑�"��$�jm�u�5��1m�F�`jH�C[!+l�U�����     �     4� �}���n���^�{���;�L�����[�w3���{�{vͲln��W{��{Ȼ�u�N^Z���ݝ�{oW���&/wn�s���{�:�۽�Z�Qj��VmdUR�R�T�^��ݴ����8����w��{w�W����3ovm=o=�z�]����lۜ��u��6t��x�������i����Y��k{������ޯ;ח���{��mn2��yV�[{�m7w���Ҫ�[K�M�����g�{h���ܛ޻�ާ�<��G�������۫�p�骳f׫�w��Owo7{W��u�y��sכa�oe'y�rm��޽���v�WV����N�ڏf���s����l�P+liU&��-��]=�.򧮂��n�-z{�[����{��k���Wp���f�܆�Vk���ޫ�ޕ�����Ͷ�U\q�-�����yRT��f)EF�E5�zon]3��x���^����or�wws�˫�F�{�v�׮�㞚{w:v��w����oyu;w�ӗ���Um�t7^�u����M���6٤���UR��<�=t���ވ�]p�[��a���1�K�p��s�go{�m<׽�Sk{�{������o=;:��׻V׍�׵��[�n���ݮ����jp-I6h)�Q^�)5��s��}�%�ޞ�OOmڕ�z4���u�l�ݽ���J鹞�����9�gl]绵�{]�{ѝ����;ڽ�ݯ^���*�l
�!U%-�zSm��pw���o�[{��]������x���W���l�r7�{ܝ��ڧ��������4���mֵMי�ݷ�ۨ����{���{���m�=K�=��ђ+�j�-��RZ5��(V���_o7I�3Ӟ�yz�jǍ=�Eڷ{ml�yz�Jy��{�{�[g�v��5z��m99�t^�W��m-ݵ�{����w���I�ޝ��gw���ꭏT��t�w:� �@2�R � S��$��Q�  *��6���a� T�T�&2���	���   1%$)?Rf��F�<S���!+��?5��¿\�+5[���o�`G
��-w-��i�$��?��D����`@""$D ���"DG� �����B ""?�D " DD2 �"#H�D�����|@��t��sp��W;�Q�J�MD��w(�&e�w��V=�7[J�ي3D&��	� #�?6�t�4�j���H�����!�S��bj^�X5z�F��-<	oyG�aǠp�j��bj�wu0e���$R�W)��iYf�S�ȭ��GOXa�����:�v�A���r��� H<�������F���7vx
�m�tU��j�aB��.�	*�A-�Fe��/Ѡ*16���7"wj__$��ӽ��b�J&Q�A�Ý���b��:+�ZQ�ݹ��j��wЬ*(k�9b���������vi�4$��B"A�4`�R
.�P/)�X������i%�	������f؉f7s^$3V+�(�RE�PWo���A���.�.R*� �G)��iյ�n��ͻ�|������)�M]\�$� �.��L\y��H[9ؔFR1^rpj5�����i������t�bM̜	���b�̵Z�,쟜{�Gq��0m�b�L��l
���~�,�;���R[9a]ʠ�uy��q|��V�Ҧ�*u�7%��B�YEi#�wKR��K2a��G�=L�aR���-֪���g7�DS[�jZ��#��@�@���(}��.g�w�u�
�=�E,n�\bX����|��aټ��ś�=�"ngb�8�qUsx�Iʘ*�)�<@�75;Vʎ���U������
��x���yp.0�wB�j8wnvr�Q���g,Z��x����Q@�����+^�=qT�z�����-�H�Q��pl�h�U��&ֽ6�K�{�ǭL�pX�ۻ��P�0k�5ݢ
���b��g�1A�}W+Ρ��or��a7�UL�"���St`�ed��;��B���(R��4-@q���{�] N��%�**r��f�n��H��(�"�F��a���(]�x$GfA�V���Hٺ?]�XN]�o�[���o0Bt&gI�
��x���H8�"������x�� ����wV�J�K�5�s��Py�̫L�'
�31��^c�VDKL��f*5�i3k-K{N��7I�:��J�˙
����vi�w������F�p���P�%(,5���cʏ��E�Pf��qqXvʦ�U62���'p����TYa6�-5R���x���Qδn���������N�-ܸ�y�t Fi��T�m-� a�����g/�kj�;73#�V`�f�X� +ʥa���V�Q;����z-d�7BPh��ț׵k�P!L�3'[�Q1�a�NVΐ�'�uI�*ۗ�����QvK��C�����H-G�%��"����ۇ�fF���d
�D�A���$�����*�J��u� Ta��v�0[ve^'�?&�2
��L���,��O0n����D��g6N��U�XGs�
WB�`��@$4�j��R�7z�A�qs���*s"H�HK0�5n�HS���Zr�Hv���I��1c�k�;��y��EHK�wle`��*JA]c���I4l�a �Z��Y4�W�;�Yxo;�l�D-��x6�%K�Qba��-�n����=H��!Y�E�p� ����U�%6���U�Y�7S	�t�r�B�X֣0Q���̺7�<�޷�QaZ��jEƃ�r@�<�W1Jz�V$n�*�B�&e=�#��K�J��v��jT���7�lJ�1w��cktiA�q�t����L�y�a�0�Q8[�ZΜ�J��;j�J�)�w)-c[ci~��X�r�:�Z,E���������xͰ��[)P5��+5S-W=T1��,XK���l��� kq뤀5���M���b����e��l����n�ȋP�a�,ŗ�FQ�e8C8h�q�,�t�8f��0?�U��ĪM*��4��9�U% N�juW	dд�P�$i�Z�7��\��fC�ʱx3%�����k�%��u&Aek:�(]D���d���ώ��_��w�����x�ڡ�%@����yx�aM�^h�@�GP�ʀ�C�݈��{�VfB�{���6ܬ�û��& #(�b"0���& � "  q��`	1��@� I0�0 ���ܝ�U�S��!�M�#tt�b�չܲ�Ӏ
�tEF�Y7��p���+�lZ����k_c� ��N����`Ҽ��-d�`|��T+%뤻[Ol@�]n̬�C�&E�)&;��Ժ���u.��A�u�m��h.��5:�q�`��}�':A���@#"��,��P;5ʳ�+��e����-g\OZ���ėI��`F�N}��]X�s?�]�4��p��U���m���p�	���t�m'��Zv��< ��R��jژcfd�]pޑYƗYm�I#�gjN'	�.5�N����w*�M�����m%efe0��@�;N_Rڌ)���.��Փ�]�r��/tј�7 �2�?��%�����!C7L�*��[��M�!�34���Uci]՝Y�țX3�EBf3H��$2��,��ђ��KQ;wc5E@`ъ�^�p�w�˫�Q�� 9�F����V�M�mQ�����y�V�2I�hc��Ǒ÷x��ҝ@KX��	G�r�b�9S���yѤY)*ŏK��F��e�3u%�����!���kM���4��Yn�l#�]�D�cVV^�t����f:F����Qh,uQs��!b���}1֤�  Nh`q�"�U�X��RwVs��B���I�����LdSt"�kqU���R�����席j��j��U�c�Q97e�4(���.V�����4 q̼R�j=�H���F�u�
)�T4�jSp�fX���p�:��ۉ����cn��v0�5�pK������jn��F�=�jL������a��q:4�٦L�7h�X��R�E�u!id�\��'pIN�/��HP�L7b��ol�,՗[$]2�pѶ*()ۂjZ8S��}�]݃���v�VT��H�p��4�لF�d�+\$!����b�N��I��*��SU��Xs.�T��xX�e�@�
��Z��r�P@���(�c)�`�ՈS�K������.j��Ǉr���j���kD5�XT���y�T݁(��*�F��t��F�Iou!J�dշ{.=�� ���or�2��%Bռ�)U�3q ��`����Jm��P�	���Wm,ۭ�M�qf��8\ڋ.<L����l9�r�Q���@�u�Z��6��9C6�G������#$�hO(vK<R�Ks��1v�i�����hY�RHj��]�B��m��;�@��Ib5�!����(���,8*�Q�hB�^@���m�6�������C�)��Zơ���xh�6�Á-9��q�,�%��-*̷�3��j�j���ݑ�0�%i#.�5�+r�U�	Jc7-�wT�B�'h��m��zT�aW�ѭ��7A�w�����n��]�nE�U�R�N���(�r�T�ǂ\')e�D��/���N�3.�XcҨD��!��"�b�n�ЯC3Pw�J�`ӳX(�[ձ]>�p���rcX�@���1D"���Q��#�B���,*��ݑD춚)GZ-R���邋ֵ�ٶ0���4��ۙY�4��+v���I<DF� P���ݚ.̉�UY�mV6&]���\�-K8)����B��a�`&N1���t�h�uh�w)M�Tm����㸱Iv����2��{
r���L7�)~vR�X�"�66��)��\����� ��,�z�RU�j3G��iV�SxIy�丳NŰ�ړJ�+V�Jɴ������F���لMZV lY���}�urܵZR]6���#Àij�ٮ�ܭe�ʙq�1�F+a��^v�[7�1k5�j�0%�4P�剂�-4�Cuq�$�q��!m�;zS�*5\yKn�]ۉ<�6�͔u:�l�-��re`�[��	h�A���f���m�t,�url���H{�h2��(���P8�x��T�K�̖�-s��
Րl4ݛ;�T�y���Ú�����3q��T+�6v�ԩ�#�W���
Y�%�� ��
�ܑS��@[.�DT�E��a�I��5k&��X�C�����o/I�*5��FCQ�ה�<Y�R�a����WfShG�nL08.�\�ǥ��ut�,DJqM٢Au��^�6-������;�X QDPy�T�Ks3s[6�K]���wEFC����Ù�$��5w��8w@��X͌�N�\Y�F�.��Ґ�f�� �us!�o	�2�9�9t��+
��L�F�7)��IU��ݱe�M�"YZtĈ���+��jS�qo:΀�o��VI6k"i��T��U*�d��uO1ע�n�Ab�"ȊW[܀@�ْ��s���f��������z��q�o�㫶\k?-x�:B�h䥏n�|e
��8ss�iLjJC��&j'U�j���j��$Nʃ#��k%+���ج�,μ��4�S�Cp��Q�+1X�W���?`�QT-tD';dS_r��q���32�e�S{`i�K"�����G�N�PH�vGk�rý�ޮB����շ����m@F�V��Q �搓&,��^����$�joL�Xd�[?��R-�c��.�v
�x����!�D�$"��-sYgxQ[����`p�p�ka�a���͢�@�kt)��qܳgj�VWq�el���ʣB�ۥJ�N�\AGb
wQx�GNM�V�Yl�$�m �a����$�&t�D^i0K�M���o¶&oY����z�ɭDt�>�Bv�h^ԗl3sn��ܚ�]2`F�����
��|v:��u��f�t�d�(UI42�l')�{tE[�Z4qi"�������#S7w��ʠ/moፗ���� �륏[�:)�%". �nՉ��R���8Ƭ�4�ѳy�r7+R�!m��0@����R�n�]<���7du���H~�5TFe[܍��i%���r�I�&�j��2wa�bn�u��+�Q��ȟ��J��&^ґQ'Hl�ҎSnp�MYǪ�-V���y@��ݹd���Z)[��
pևP�I�{�z���m�a��w$M�J�7e�෌�0Q�U�쫤^aʔHV�?��)�v�o���5�H�c���vkm<�v5�kuytAP2 �7S��{'�Em��Ezq Jʶ@9{x�{�.u�0�ttNN�gi�����˽���p�n��j�b6�i��h4��ve#��	�[b���J���������2e*�4
"�k^�*7��(e�tܬ{�q%�F$h-��q��h5t��j�6Іmm�@M�j�YL�`��mm�V
�P����_��T\ܴ�^c�Vn���_�J�StK͆=���W��8u�,
�ڻ	�l��R0c$��k����p�Wc,(�SZڸ��V$ݵ{����^9�2�3���
[V-����u��-۬(R��ن���)�_������rbe��P�H����T0 �{�R���M;&��7WYbm���bI�{\p�� .��vfQ)Y4i����	�z�Ӈ���֦\:��cV#���y��,*�7�FTF�0ݧ��6�Lz\n�,ܔ��R�.�&�uѽ)���ԬЧf���4=u���F���%����=� ֫������G`��x��C2�\�sV�9$ܬ��L~�kw��X���j���M@4<��*+lL�� mR�4\�U9Bֈ�+h�Grfc-8�B��[c^�r���Z�7U�i�Cs-~�Ua���ې�m�j�u*+1����!�	v�"�V��j�z+%5�dd�%%����Y��5Nعy��wJhx��{F���s�+t��J�}�h���-7jgVEЛ@�D	�0��즞G�cˊ����*
���������9Wxh3v�ͤK��V�ԁ����!V�/,-���)��OV�57+��O��׍���Y���4I��hef�tњ��k2a���glj�_<�+lU���'{Nc�����=��i�+TUr�-Zf�ܼ���EU��.�:��2�����0
n�KJqǸ�L�0,����n�Mp`�n��N�ec��(��0L�����YP�6�kC#�޹��0fm�%Ǳ�V�P�r$ ���}3��m�����eH����M��7���5�w��	�U\s2��)���f	i�{鎒lc;Q ���cs1�Ѣ�xP�؏���=Ō];2'i�9����	;#2���Dm�Z"m�R�S{���I�沮�V0�*Ȭ��P�4���52i��s]�L\�nR׸�떝�kw- o s�t��IC�����E�4��s�-a���U��W�H�� F�2Qš���r�1��us?Jz�D`I$?%De� w�B�4Z�n黣�c�.��K0¢���B';�TJU�lʶ܃�X�6�3x-խZ�֓3m�c`�Ҍ%��g)^d�I#Y� ��h�t��6S�1�3C�Z�ӧ��R�U��x.�f�;g�v�*?�[��kVڗ�jI�+P҃V*ۃ1���ڰP�*9kMP-<�8���Vd�]�����tӋXCi麵HĀ�Nl���pG?Z�䟖P���a�f�]\�]�P�@X�N�^f]R3 OHsy���tC4t3�A���@�$P1h�5t��:gru'MQ��A��d_��kSxn��L��Xx*����-A7oS��u�jb��m�Yᒦ���7Z�Z*�)՚�-{��5X:������J�r�3�\� ��FU�8b�fˁB�̡��h�t��s%�Q
�S����(`��QՇ�������քtw5�M�$�)�% �EN|�Uk��Sv_w�x���뻻�v=`�Q��)�Yx��ܑ��G�H�I�#}$o����I;���F�H�I#�$o������G�H�I�#}$o����7�F�H�$�$�����7�F�H�I#�$o������G�H�I�H�I��$�����q�@�2%�,RI.�:���,ws�[M��F�7:j\Ӯ�ʈ��*�ʓi�ҁMwi���<5|�u#}WN�9]��\MsOs`95��$�)�K�v�2���#�Lm�d�f����Ա��7\���ndENtmoQ%����M;��w�[�[�m��yۭ�ݍݜ�̙OV����- ������i'Ԯ�
f���x*"�m�W�Z�gB����"8:>%���RN���m^a;�
sy���j�z�+�
wU�{Oy-�P|��9��\q�	'2�BX�o��1���,�{K��w�&��O:T���Q�Z�+.�^[�Z�܏z�Muϲ��0`üp$y��z��@]tkr��+�PR��/�9��٧�-���7���+���&3f�7,e
$qK�z9=zR�B�.K�R�F��GW�c�H��^Y�%]����Ʀӧ�gV+�q�Ύĉ�6�)�Ѿ]���{�2�� 0���$��-wR]�k/��e��jE�v�p���j���͗$���z�d��zڈԭ<�l*����|��Dv\lU���Q�2v��H����ә�sq��v�5��q}��kӺIs�m��B�df��xfr�.�*X�P;z�����Ek���msHB�\�'k;oF�Ѭ�Զr&9"����*�r��@5;���ʱ�Z|����̳�i���������&.y��Ĕ�Gc2$3z��K�&aݙ���uf;���f; �l�ٺ��ܛ�r�c�>Д2jyR�VdJ��ŝ��,�0XK�e�*��"f��gavrrh���Cݐ'�F�l^1��]��=MfҮ�+���*3���o�sAۦ5�:��A���u�
A�wv���~��_nC�Չ\�+S0�
�-m\��@Ǽ�|��2�{�W7��+{�q������΋��]�{���0de��V�L��OoL^�������/�m��s��B�����i鯋F�[ыU�mû�V
H!+@�X:酂��9%��mQ�u�u;3hs���r�):������K�U+�;�+�*;������	�F�o��ꦱb1F��
}�*���[�u���x����a�b0�(�O���Ӽ}v�Ą�^�-Ǐ騻���#�>�^�����ca.a�-C;�P��A��u����7�]���W\x��HB�&�h�L�����4�쵝]Q3����2�q���؜�k��Ͷq��pԞ��ʁ��S�!��ԶR�өm�rEK(^�t�1�l d�)�%|���{���C#�Λ�7Ok&��e�����8!�k����sXN��Ǎ(�4��ϹM�/9�<�:h.���(��<��p��{\0���f�vZPH��yH�t��[��j�XՒ	G��;n���"ԾV�N���K�.�.س�G�7k��Y����ǒ�XףK�ǆ֠;�V�=�E2�V�X뻥CH�5�{���=C���H=0��h^Wl�u��OvC��k�\�y��f�Lq�j\鲂�}ӻ�ޘ��d�K6gt{W�la�4, ͤ�15��J2��|6R�)��w���*�ݛeZ��p��\^ҩ�7b����wSN�Q(o�oA�8e�	=�L�����I\�]�5�}�b廮^�[�*Э�c���Wvŀs��֩t2j�}y��엕4Tx���s�79sq	r.~��P1O
��˺�M�Byuf#o:vY�T�U�1e� ����S�X�
휹�����Y��j�˴6;<�6�|I���fZ��@v���ۍve<|{b��>'Mu^uo'v-ړKI�M�T�N�U>��i�D�z�����=� �P��,�'.��{����>|��!ȝe=k���F�@���*�%-=��`�C!�7��y�X�]{z����lh�'��^Ur�n�U��KU%���V�[С��]��a<���$��1������L)F�1��k����M�8\sHZ*��ý���v�Bi��rfWgbm9�GB������pΡC,.�U{����m��t-�0��$�� {:�_d��}�MN�I��1T�9ٽى&�:`�Fۄ�v�2�W�R�4��Nհۼ�����ϧ�#f�{��Z7^b:�s�V�N���:N��a`<�n�6
�^<F\��͚�N�P�͉��"��;����e�����̷WO�y��q�h�n����L̡��YWG/���9��n������*>n���Y��ǧN�:�|��8������w?td^�T�n�ڷ�w���W�  �t���nfkl�R�A���f«<Ł�)hb	�ͦhr]^Г�[\��ɠn�<)f�Yցd�B\�.wf"*�os��aK�w����C#��1���^R�+q.�Z}���A�j�5���v�)�Z��F�k8M�ss�A(��>��!��k�WG#*m�v �tnJ��ҵ*�|�aǲ��C0_5u
�p%�=t�Z� _U�cy,�)!}KNwj�{��'��r���e��v+{Ha�q� ����$��I�W$�OU���yG-^� 
%��Z��.VR"Wm�ȏT�$��K&�8�Y�e�vWX�{
Z�����r�Vl��[�GNKV�	`v+�&Z�e�9��m[=zt:6��c�*sS��C����eVS�o;��
���L������K�W"��U���,f��v��x�A,p���yw��zR]x���=�rxn��4�*\5*'y��8v^���MN4��"�ݕir5�k��<k4��`�ư�E��A5��r�㷩~�k�X�V�m��i׺�C�����b����<��r�b�&��Y���P�m��<�������(�r.kt�'dV��@X+��8��ʳ}*-�^%��"y��PŬ�77@͖�Z�����A^��u�yn�%r���e��n�'҇V�<X�*}k/yu�/E�<�C*��Hs��J�'M@�i9Ô����s���t秙׽ǹ�6�Wb_�΅�P�m_TY��&D�v̚��؄�o3���Zܠ]r�Y�����7w'V�b��`7�vEԭ�\���Z���1���X��)�<k�"��7->qРUvgn���A���U�&lp��F���n����V�̙�Q�wS<��0vΠo�����f����U��dP�JR���Cw�:mc����K�n]��r��L�<#�xM��7�i��b�kr�Zf���6lG{����4v�i�ރg>՚59܊z�J�N�N�3e��%�|^���:���I�44�6|��ݎ�CS:M����-����hgfS5���r��%6�G7,��ۯn�r���0.\&�����ڤ �z'�c`�a���b��3|I��]F̫��N�i�o5cs��xVٗ��ح�6�+\�1'%,��lVs��YL�"1�u�&qR�q�D�(i�*�@�/h�92%y��v��4�&y���F�wh+Fb�J���)�m#b�/%�Y��^s�}��#4�v�]�F�j����l��O�N(�w��Z��r���Wl��K��Zgl;�=#��@��s��os�:ݚ���e�v(s�CU�ve��fP]�%v'�5u+o���5��%Xu�J�d�x� ��o�m4s��tI�t�7l�Cb�a5�ǵ�,��Mb����L�Jj�OnC����8���� ����*��v�nV T���se�a_�i゛B��عk���ng��LP��Is�2��._v_s��g���G��W1�4=}�:���M����d'�kX�)�3y�:��%��t�l��7��}�(�Զ�w6�9g!Z�ae�|�E�0 �����љd�=Ҭ�-G�T4�4R`u��ɭe<w,�h��L>L����Oe�4X�3��%�И�ڍzNÝ�5L}��C��w�!�O���.ԗl�}u֣��b�C�6�8�dL竷\vK�K=��YZ�_�>c{G��3Fuk7ggf}�U�}�
��z8�Ŭ]�cn��I��Dv��(M�{������AZh<�b��z���(Oh��v�X��e$�m���;�m,���K�C��/�n��;Ǥ�!����C�OV-���^L��J���u�pe�q��3ö�6,Ԗ7Qf����qQG^>���	��E�9�Λ�%
q��1r݂#�A9%���Z^!֫�W-���GP<�ȅ�&/ݶ�gط�t�r��m�fΩ#��.�K;y.�<K��d_V�Ȑ�Y���0�(hF�`�8z�=��Y��*h�7��ʻ�ԃ�-=��;W����ެZ��3N��l(�6�+���Y�}�ְ��w����1�忝|����j�q���d�[ߕIs��>c2�-=���i�ⲣ�$�1
<�!�;Bn̟��1��%ӭ���k�@��7��9^���u�f���p,�f��#c�!�Nj�B�q���Q:�\��l�\�4����L���X���y����M���ť��׵���o=H[���!�s�1E0v�V~���O�R'A#;�����WӦ�x�&w3 �I`5�X9�MܢqV::�>��˸ӒD�>�*�e7��G�*��י5C�y��l8u4� ؝��Ψ2�&o����N��t��91$Q\����N뻬$11Y�-��i���^m�]qdc'�P�e��Ej,Rf�1�ѩO��w|`Y�[��Y9o�Z�c#���
�5��m�Me��{^��ļ�:W9�Y�f�[$�F���7}��}�pH2� ��'���S��%�Y��
֨+N�-
VB�����Y�b�A�)��ts�6�օQ�a$���:��w�S+���������j�O[&��[�U�X�L��{Ϻ�����@��A`
�(����!� �R��0��_&h�9)I���nm]X�&��y�>Qf'�r4�]n���L��X�%ɠ&�`ۑ"��%ʔK��2��Z\�Z����b�>5�����Vh���{��*i��,^�S����V�-�0����Zt�i6��WIU�ID�i e_����k���6=������4.[x�Q
dQ�&�R�$B���ǻ��G<��ޕ4rh���W>��ܝ�{��
�l{���b7������r *aN⬴��2�"�Iuk���[B� )h��\�/�Ve��͸�I�]����ܽ`�yz��n��7���].b����r�,�yA\����D�mqZln$��uv�h7��5� ����#��eAڃG��]��J�o��qQW
�gVRdP2�
�N�89��p^��N��
/�/�9�ȽJ��!ue'۝�⩻��J`��u:V������t����u�a=ǟ ����Z��$�To����ug\�a�,��2��;<S�α"t�\�����%��T#���ힾ�W�3
D�%j�V�.ɼ�h�m��=��8�A�JZrV�!sAN��]�PivwHEZ*�]���!�5����=�wFl޷m��,*fR��훪���L!s\Ե2�i�o-��5��*��ō��g�����i�
1[�l�4U���4㭈�z��ȶf�gH��%�}�=ԇ��P�a!�ѳ����8
���:G��<�r����5ht�S�S��j�Wt�![kt\�̘.n�kU%�ԋ�|�4���{���B`|�"J%��S+���r�1K*��N~X1ƞԮ,��VW
�&��Y#�]o-��f�t����!\�B�M�L����/C�Y����;��9�L�������m�A��soL�v�gcT"�J����M���5��ج���S�5l�f�Sv��]���]4-d8�+sb[�'Taą��Ѳ��N�u�i_���=XzM�Կ7��Y����&�*]���@R�\����L;�T.֒j���j�;�u��O�v�:W�DK����V��+�w\�T7�ʱ{H�5�7����or��ڝ7�i
%j� �	�)���hR�������P�̞G�Vql�@�خĆve^����RL��su�P� ccm㓣f��uຽ˳��AemĶV����D��e�$]������]f*M�U��:�)�n���9�`\���inf����Vx'i��L}pd�f����tsUY;��Rƍ�B�;��Q.�6�9�;F�-�����2T{�B�nu�l�x��rP;���t�U��u�'12�h��Y���>�Uo�Z��\���m'�ON�n��+ZG*��|�P��=�x!���d�d��s*Z�Nء�Om��@j��!d&�t3t��N��ik�lb{77�P�C'�YOP>���]l�hIesױ_Qo`���Y�x]NX�cn��m��s]g	� TK'�g,���<N�Y�y٭�d�5<���	&8hP0�rޤ�w�ە���]̬0����_n5v��a�����^`���Ε�ΣM�&㵕�&R:�K�9�X�����l������&�R
�AS��wrީ»%��%�^.`����%s+.�zjt讶��DNC�7]�$v�αË&Y���ӳ&��OSg���l
ػ]ϲn��')��^��	K4WG�v�T5:��N�^��2�Q�������y'"	޼wE-уPPԧi;��.0�$�lq���[���� ��]���Z�j>U�ضԩ����s��ų%��.��9D�)G'QP��Dae��y�V�pr�c�
��"�NU����s�(v��E9Z72v>ؔ�m�zѢ��ޫ ڷ��%�����	�T\��n@�(��H����z/ŒVd���R�/��X!��{�2ttoţ�r.��b�c�K0�r��)-@�vokj󞮢dT�*.���˷�R��Lf�m_'�����s�yO�E��z�F���X�}H��[Ge5\
�P�q��>�hݏ{��ׂy�����" DD~���" DDY #� ��?��!  �_~L��ҿ��G�$m��㣺4wz:}$��NpQǄ�y̺{5��L��6�6i��x���_Ksa}��Ԡ���kƝ��G|�'Ԝ��*��n2{i=����qՖ5�'��_v9�d�b�r�.�T�-f���뺹��L�� ʠ�v[D���N>�'N�[�hۭ����Iu�>�끌��+z��;�;��O�ur�(v�N��:(X��E(p��:�u55[ä����bΣć�WAS�����r����1K�pY)�u3��u��s���x`���LO{Hɞ���;<�S�rpT�Ds�]P~N`4�غ�9p��f�t�$���gvU�w���a�=�7�z�
�9�O60f���Yj�L1nI8�>B��]�.�t�f�cD��͇���m�����������!��k:2Iw&��C�["�WM)�sw2�n�C����u�RwGs'm[���l5��Q���ū����D+�g&��z*�jn���8>���V���sX�s�}�^�X�V��_Z����/�|I�*Yl<��C���Mͧ���<{*>Xi�[D��[O;'��+P74�����]�1WG��9ߺ�A]z�\�z��Dq}�f����8�ő��m��$ ��Թ �x������+f��J�[��ĸ�ٹ�Y�׫)xlpyd�J=j�6�� "<!�wЀ��˚(�RǼ�t��b���^l��w0���&L�#�Uc�nw[������	9�h5C���2=\c� y��-�v�ǖ�-���S�__�6Wn.�>Q��hV׸;ZKEڠ�d������`�oׂ��vYc��t�����G�M]�כ�K��i<�����:�{��U�!�'��Vў?�ލ����Ֆν0kJ�5i�����|0w�Ud�OWL���3�2���8����S��̖�6�uE+�ó~�a[g-��]4G4y��:^ ���L@� �����|�k�Ɗ\wC�Кa3�m�j�OQy�Bf&��m���
5u�j���|M�B�^����X����7�0�m�^m�|��y�i��h͗:��:o�#��>�#�@$5oM4�����rl{C�os�{�i����Q�z}�򇳨�^exx��;qL��
H��ȓ�B5�t��,�~[���5�7{ӵ��x|z�";�rx_�H��T���zt~�k*yW�롈c����|a"ȀN��;��.���:V�2E�6��Av9y���� *B a �DBH��0��w�hL��9V#�O:�3��R1C�]�1e�ޣ���B���)��m@t�@8�ٗ���Fw��c�j޵c��˧+�O{i-�L{��l�Y��%���E�.y_y�,��ɘF^g�w$/ĥY�~�,M$�ݺ�~����0P�zrG��٭@ 9-ՠ ���{���N��L0(s��o�nV!N�y( D��/#�C�������5�^�X�n��p���U���v�l�jy�Y�R�J��9�^��,~�����3v�uL�{CJ3)��9f\gyǃ��{��2k�e-<t�[�-�Y���M�a��̸N-�����`#�����D=�̮�cr��&k�+dp��p=Wfޏ÷&Ш�u�׈q4��v����)����@��w�og��o[�A��~T�]�Ò�P�ѣ���W�_�JF2/���)�v�3�q��r.V�C�ʇ��b�*�c4P�fo��Wv� ���n���K�x}��Uzd��&�t wSֽ*�L@Ĝ6�91�N"p����`"� ����@$a��0������H�:�±�IɂrT��N�)��/9Nd�ۦ���� ��"�B$�1�&�s��V� `���Z��[�ﺋ)�]��G��N�N�V=��餲{*	C{w����1�
�\Y�۽7�L��攲\]ݖ�Tq�X+�E�gM�D{�^����|w� ѽ�Aj���M�os�]Đ5״�y�X�C�d��-�9멚BpZd��'�p�i����"���EN~�^G�h�v�/�ޤ*^h�;�n�8�T���Y����꥛�~�=��rmn�Ly[${WawU3ޚ��6H��vS�F��w���hq�y�����cX>(՜b�S�"�W��mԓ{����~�lD��p� u�s���Y������d�O5�ص�fJՊi���u3��J��HR���,��w���ݔ���.Jz��r�:8�:��E��Gw�
Zn�0�{�Ƈ����2����K���Pu4F�ZH8s�.ri)�=�^�M��$/1����L�f_A!Y���o�Nz���0I
c�0��=@��$G�7^��gr�k�jt�B��@s�P�5\�
�E�C=ѢQ�_��?@�3K�{ۆ���]�KV�K�6��!�T�`�<'�����o�
r��h�<�>S	&���9�:ږ�;;��*�1Fqua]Vk��l"y�̺
�|��V�J�����YCLWt���VOk̀����w�l�}Kܻ���-"�6'��r/hȷ��\�XO"�q=����U��rɺ�5���;�G�v��R��dD%�����W~�~�lt��TGa������c��Bs������r��ܗ�*��!<{j�(>$i�d�Bm)��״ 0"��P�7C@�+�?v������v������]�Ep�|*�Ak�+���_��qP�H� �.'j[촦:i�=�P�o���K�;{�����?X{��������Q���m�9Y�����L���[X��a����Q-��Z�,5��2�2��n����4�z�3�rhd�	'h���� ĸ��.=+V;��*mv$s�|�g�OWW��:�ѻ%C��XZ�W��<21�]D�>�cl��k���q�Ɔ��$�W�W��t:g� �@�@�ZI1��;Uy����_���H�X��Ss��=�=�@m�
���E��rU��v��C�0Qb�Y!�?�S�@�i[�If�ܱ�3]��lI|Qc��dedHa���l����%�G��'K��vJw3Yʂ���O�Vӊm���;�HX�&�[�k�x��r��qz��k%ןM�1C8j�����*�`�Z:_=l`��O����;�z��X*���\����gZA�-Օ�WFǦSb��9�iz���P˚zn|���Ω�j$DGz�@��pGƯp*��U^*d�\}7w��\l�ut��� ��D׎�ae��L�n��v��*$��Xle��<NҼ��S�� �b�3N��RdDE�ԋ��Z6CQ:��ۅ���r�L7��3�����bL����u�<>�IMOl�ʀ�'/�䫗n�Z>5�=8J��Y�_��{_���}�Fm��b=^���W*�wң8=��Wf[��4A�v"�Wu\����3���^ X���;�ܯįz��[s�l�e
Б �9	b"#� ���U��x-WIn�$vs���@�h�����ȝ��W��o�UtJ:c�2�w��T7�`��߻c��b��R+Cڋ��2u�P�� ����m�< "	 ���,�"^�O�{�$/�w^_)�f�=�յ���2��~D%RF0�1
@BN�\��+�p���%���v�[[S34��]Z{��l���rj�.�dR�]�n${WokJ��o��*$��Yz�x��=(��h�����㔓��N2�5R�7�᫇E{l⥲��0��t�;S�K�1��s�s������D@�U{&v�oC�N�G,DF'��4 �n�����f��U�l���P�H�ּ-�����^�Ŭn���w���\]6��9Pu��V���5(a F�qA��a����$�G5롔,��
Dxww*�]neOOu8��UH��ZK�DwSƅ��=)�C����z�Mn�{ڹ>Y��2���F�"Z�ge�打��oi�>QjJ}���6?\�M���$����u��������&���&���id�i-�=��(x8�������$m$��n�o<�[���� �E���P^k��+��z`��+���*qͼ/u���j�.X4T҆gC [�.x~���dDC1��!�g�	��,׻��Q=������\XŢ�̬�r��_	�K�2��/�N����8�ǒi��cɗ��}�r�y;e�O^�e�:�ͱ�z��D�Q�v��QV�Fܝrp1�e D�zvS��Cw��T��M�}�l
(A�	i��{;Uܹ3�,���8��٭�:���'$�I���F�Y4M��z��7Z���@23��%Yjׅe8v�^ 	�RU��a�<�)[�ʙI���u�6[�������5���:)	7��DMwʄ~��h�}n�C� ����'���Y���8Q��Ї_F��ur��)�r�K'n>sYμD����@z�S�ƃ����p}�+"Ⴝ5k4`�OD���� ����{�U�3I���J��$Ġ���Y�4�� �.O�vW]�m�=7= �{i5K�0�"_�q��_��͟G�lD��R�WR�,�>�����T�'Q<hTj��,r#ƥ]80Q�~m�\���UA���+��;{�6p��Y�ү�=�;��I� oI'}�䄤(�=x�B�ǂi;��������Ě��hMM�?I�t��yیR@x�py�%�34���י!���P�!��g،��� ��~b� ׺Vy�v�$x�p��c����B@x/�r��il�A��l������q�ްۛ}�rq�!�$ h Rā u��͛��I]�.]=X���ܺ+iL�'PR���o
G7��wς��^���;����)9�ێ�+�b�B�\���ʹ�D�V2��|�0|qB'�R�)YN8�. P��M���]Ҩ@� 1H��w�g8Dn�{�)]�hۏg|����|nr���~jl� �o�W�2����2X�=�������`߁^�d���DG��D@��i�}Rg��/6��]B�cXk:L����U�G<a.�P��\5{� �^6��tw*�v?-KCI����2��nX�㖅d�n" $ ��\�0����=�P0��WV1�N�֔u�k�Y�͢z��äv(����/�kj]���jP��b�(�T�m���VG7�}��x��Jz�"�aR�`�Z�p׽嬖b�)ܚK�(�~�6�t���el�/ʸV�����fw&q_�hu��!Lf(�ʛʾ:U1��� 7"](�&����FY��={���8t�)h��E��m~T�y�	
�Y]z�f����4U����,���qš����"�z,%���& [�^�j�ըz�U=u�wqk����\���
h����$���x��s\V���b�W9Zr����n�D\aV]n�R��3����-�qgF��f8ntV�N�������T����ſ�<��f�t�J����`]s:�K��i��!Z/Z~�ż�q�L����i�Z��Y�C�+y�}5�D[Y�,�I�\��'yMӊ�������/�{�̨v���zD�m�7��S(��?�$~�A������xe\�S�@�.��V\��� ����Ǻ�U���y~{4�Z59�ͯWpk���CI�c'e)�s/E!m��}X�w��HI�7f��䎊?��{����6;�O�N�O� {�@��^F�>��tN�zc��/�n23	rPw�jz�:> �T����!���ϼ�-K1Iq�홎%aw�b����C�eW-��]m��~� �1�rUW�+y
n�	��I��ms��;S)1Q�G��c����r}Y��<��rFO�Q;%�Jp1O��B�c�2� �x�C�XJl�����g�-�(�3���̇C�ѡ���B0������,3w,l/$Ž��(W�����A9i��V�J�u�4��tzqN�1z 7*�����l^���ȣ�,���uvn�:Hw����)���
��-W:Ƴ�H��׷��AV�h�0$�>[�Okr+=^U�M�~FT���dO.�� �p"��I��$t�t�ۊd@sf�{�\ܮ7ZiyEj��kDQ�J�Һ�JWe5�FʰM�M����G2㶏��Iy��Y�#�mȔ�""�`k�3����kGxB��Vb9����}�:pRP���K�m�.qy���� ��ۍY�����MSV����y'���eI��W���F�]vp���j�^�J�p�O��^�R���-��y��HX���F���P� ߭�C<W���WQ���gk��>  �.n�d^j�஑xl7��ܼ�=�8�p�dI�}t�H۬N��4y���� �y��r�w2�B�V��w�� @�E,#��%gs @DQ�=鈀�Ρ��ޔ��Z�)��y����k��Zw��H�sk���c��@�OK5网c���35G�:ג<���H� !��B���!}�HY���cE^VM���fO=2�:j���2g3mq��U�[��$Ic��R,��	Gw�S�����u�9�hu��AmƱ8ASD7!�H�6QV�'�6�L�孽��q�qEA�&r��ʑ�&������5H�F�r][�q�5y�o��U�,Id�3ҜaFܻl1���,����\��x'j^��(H$Yn�w1 $�u���iC�21A�d��4Đ��)˖
�oK�;��W�C������Y��(���S�����	o%i�+G���N�;�.RWX8A���W����6�ͺ,-}��t�Ol1��\/r���6�[��ӅX/��)Y޾Y�St&���m�;�Qɵ�f�Ԡ�^VWY$����β]�Һ ,ʰ�0Y�o�!�IԾ銯-�Q��p~|�Ў���۽��R��M�jQޤ���[GP��yY��F�4��:N�#�2*49y��s x��������Ǩv�	��Ɨ<u��.П�5ww�+j�m��1�-B���o0_u.@�r0�jԡ�	�4�D1�L���"))�WU�H�`ʡP0AD)�y��"qJS���F��4��SC�7x��4:�`�=/Ƃ'��l(�̢l�j��|��Sm"��&LMBIa�Bt#��ڳqL��#�"! fT�J�JgGh�2AÒ1�����xx]Z��������XV��}-�i�P�^�w�����Z��,�S�p�R$��*u���D\�ښ48QV3��G/]�������[���]r�ܥ�}�՛������Lm�3���un�Y�Ik)�!뉜��]�6��6���(b/��榍z��!U�o-��D�����R�-�y{�ˬñ���Q\��:D.��i^��WS��u��p�.�t
�ԥ��b�!=���V���a�lኄ ;4��Φ�EU�*���跄oav�F�wϮ�ّS�7�[��������I�V2o&��؊�|�R�F�޳ۼη�E�bw�7�]�.d��`}C�^��k�E\r�l���G�.���%qNyʈ�X<:�HECos$b�٫"�4˵�Z�tu4�[�n���0�8�]%����+��t�%!Vq&3v53�V�Y&d���b7Ӯ�s^���G�"�c,aeѮ\�w0���MG�d�'u]�,wW;{���y��.��1ʠ�O6�����U���	���8>�G5�r��z��U#��EI,��"�ޛ�n�X��UG�'���ww�ޘZ���yw�Ӣ[�̇T�S���$�x<���q�zBٕf�J"dm"Pشkj��8�b�"����wd�T��h���ҥR�d6��ᚩ��� �yɶ%5��]i��g��f�[���E�Z����]���h�����Wl�Y��J�|%�r�+_)V[��С%�!k���h����nإ��7H�c*5��uۤQzr��q�uLu�����5���g"�vܔ�Bs'p7��!�5Ƅ�E�,���.s�|��������|�U�J3����ӎ���e�	�����t��y�VӻYݜ���*s��#�#�#��`Q i��
l�4�F���K1C#��uh1YdC>"*�&��:,��B3��"&ЀH� a�>1�+�q`� #� ��>M��;+};�
�� iF�4DB��,H��I��@�@e�P!��� �#b}W0��aY��Z� ��\���"'Tq�&�<�Q�v�3bLB����5_V���ϭ�f�D� �"Q#� }��,��f D�F��F�0�}J!��.��e% "�d3 �%�Z�2#�Q�b�DC0�1��0���h��c�0��w,ܧ�}}\������	�i�d`�f�Fr�B �Q�<F�F��D0B0�}Uǈ^8�B0H�0�DI��ȣ^q�  {�I��20l�n�~u�ݜ��;;�#ܡ�1�G�� �1��F�`6� c�3
0OPJE�bL^�H� �� �Lv��f	 �H�	$0 � $�&	 �0A A �� �`�`#�a���G���5��]�W��5�7�xH: �b���,ɀ	=�@0	��|G4�`G�a�Y	�b����ADQ��ƌ�W20,�}�1D�F�Qf0� a��{��\���V��|7Q��n��I(�0�	0�LD0��ߔ	#M�mCj!�<I�,���0�� $�@!<�� +P1������cP>�@f<b0�n�" ����֦�������c�,�0���9�1
� L"LY� E�@���"8�KPr��$�3&#�C"O�x�`�j��"8ђ�$B1�CL	"0&`�A!�#H}�}AW+�o�����Ib���O��">0�`qf '���2�x��(g� F(Ǎ=��b�B���@�(��C,�Z�dB1a���f �ZDq2^i� dId	I��f�yr�S��0,�"{lx�Dau2 �	�|}� � J�1Hl��(�f�a��A� ɘ��I�����8
��D H&+�!�(�'��`��4 �uq>��-��TV���e��-L�{��� Y&J@� ��Bkr��3�-��5��\u ]C�A�s�iI5��V[����w�lJ�ˉ����wWITTz���ܾb��줦�h��f���DDg )۠> �@<�#Q� # ;���F���@|E���I�b�1�F��1>��	� #D_��>1E��!���Da�c�Z@� B{��gm�)��c�� ҈�#H�HТLa���8������E�� dO�fq�/Ȉ @� s(Řޚ���?��؛�-�"(�:d��	�pɢ"L�� y(�@��ɀH��0"d��1���@��"�(�28��!�ID@$x���� �@'>ϸf����Nh],с�,�Ԇ!p��D`� /$D`"�$yD	1��#�� x�2��	�I	�#�" b����H	G�DD|�N��� (x}��>���i��Wj�D�D3)F6l�����@��8�"�"> #"<Y�D�.� H��"4�ʣ�01���Ř�B	 a�2b,�c��H���Bc�5��7����	@�	�@�4@�#z\Q��#�Q�H� D@$��""�@ 2"��
0(���ő �~0�(W�F",�"+2�a`I �ȁ�@����|�����Q� 8ݠ0+�
"<a�b7P�$a�F �@�|1D�>1��Q y�D|>@28وf"�Dʖ�,���"H�B�q�@$3� � �;�0O������#L1�� 2���Hu�@��D ��b$�G�6��<����$���4�{TI�B�Ɛg�1f#F(�'��F >�qɁD�f��{˲������=T�?��O2�����I����,�a�Db��'� � i�̴��� ��;�r�
 3��q�4`���4��`� [bw��&��^�V�>�"�@&8��̐!���A04� 1�#a� <`#��7P�1��H�F#�3�\|E�a�����Fa�i�1 ��G���!Qh@�dO�}�_6�gY@��7r��8��J���c��0�r����� � �"9���E)�.�(uMK���PKl��R�y]���ЭR\�6-cr�ܨ�ws��8�u��R���7]��sᏠ�H� �R��3X�tY���H@&0�)�H� �����0H���f�1�"�|�,� $��0"L��QH�&�D��������"#�,LY�F��W>�p5ϯ~��|7o� @d�"`AFݐ>0$����fb<���0��#Ha��!�݉�	#�`����6D3�4��& E0�
1�@��r�DB����#ҟ�7�����@�&���������A(���4�~� qDi�`")��$��ր`��$�&@� c@a� �Vt��E�+�z`:Q!�.d��#��D�& �G���^o��n�ɟ�u2��I�KC;�6�!��%!�VZ�i{��Ki��[�馆��ɱ� �;y��b7rU>g�܅SN�5ļ�
s�oy��zgv�\2�R�<;�շ|�B����(�S.f ��h&5MZ�;��n�xC .-d,#D��\Z����_`���]���|�O~٣��
�t����މ�/����L��k�"s}d#�t�'�˓�߭T���A��*z���=��`ӗD�j��]�e��� �V<IϜr:�{�d���/�C6���$w�[���s�}J�����Z��]v�w�*[Ղ�3w����a�-����� 4G�$8L{n������LG=�n�\m�C���D�;�Ag�����G����Z�SP�˨��{���{v��&6(��R6�;��8��2LDy��Si���-Rdl^��H!�r�h�͗ZPW�t]v� #D�D��!�Fj�]�{{���:QkQ7}ÙG)3��aQm��K�+�;S5��\�[]R<�tN�N$���'Siu�z�^�;�e0������2S��u��@��i I�zܖ���Wuԓ/�.:u�Բ˔'�6(|��C,vyn]��hM����U��R&��FG��f:��f�]\���B�(�x~~F�Kd�z{-]�;�Y�O}��Hg�yq\ۢ+�]7�m��>^G�m\#��Э]!ں��gfz]��s�1O��]��z���n1S웪d���k� ��O�ٖ�� ���:�+��3��h��T>7j��M�ٯ�
��Ƚƞ��a��H�5d�����d34�����.s�	+[�/�ԣ@ ��p�w���9W{�6b�7>�q�G���Q�ZZ�)D�]��G�ۼ�d�u"���2K�3��X� z�z������~:����M���@�x]Fz�ܹ<~F������NJ؀ k�A��W2�#~��z�M�<��Lt��* �]v�!���FUC��L�wNN�B�gt0��J&2Bd�9�<}W�Z���ؔ�⍆�Ջt����GѕS�pT�>��{2��Qu蝹'�Xz�@�8f.�Dy*����u�Y5�	M��O�`���\R�bD�"��+h�çUwa�˫+�nը��}Y�4LDD�� ~_���5�Q���M�q]:����L�K:{�,�Y�b��$'smuҹPh*_�g"���;�>�V�5��N�u�|�ˮ���@;�yw׈��z��q5�e[5#LA�����ec��>1yfϷ4jY'O2���^>8p��϶"",_��e�R?%�O33,U�.�C��ڪ s*)1���{�o"���<���<b]�^�!rӡ@x�}�{-Z�ͨ2���	�#�}?(��r�W��`��D}�*d#ЏKF;c���?P�k[kV��z��UnWX�T�{�2��e3�v�Q�/����U��ws�
ʆ���#���o� ]�;���ꩩ컷M�fc)����PQ E
�Ivb"���{}�]x���o"Bi1dW����T+�Y�H��c����x=T���C���髊��A�|�m w=h��-o?��q|k��o��(��'���D@�e��Ԉ��-��w<(ef�k;}�h+��}&$sKÉ0'�<�UTG�h�q����b�0��Jc��tw�✩��}�K�m�v«�o_�?�%�h��R\\��kn̲��f�r�d��PiJ#*:�u@Y�WO�Wxӻ��1��.M��(z�T���;�㯽f$z����Տ��˧���E�l���C*9o�l��fi�a1��]�����;&�Hw ��I	 I& �`� 6�`�&	 ��A�	���}�7��$���|$�T���?k�<��+�+��f���i 0��� ���b�_l��gUvXݹ\���
�Τ�WT���LΈ�P�HZ~gwx�^��B1:�MĨ�Nes$c��ԑ���t_���?�.;��_W��hp�RW]Р��Տe�9������5,ɲ:��k�R�Q=�:&׳�7��D˘dL��WD5ZDK�<�\�~m߄���_`�; D���g�����m����_*^����3iF��rB�Le�v])|OY�[���+n��e��i�]��*K�Mu^�aMcQ�5�����/3���&�-�IV�4��@��xȒ�>MȈ�ݟ^�7��̼.H؂*�6�� �8�m*��D��m�����O��g�w�����l���߮n7��t4W�ӯ6Y"J��������"�_@��*����>�4[�X<'�����3�!X���\��/Ҿ�t��G�,:�B>'�����{(��Ȟ������
��	US�����&1�6N+���;�Oq�9��]_4N�B�L�z!���� �Z�RR�2�:������$}�*C�B��u��*�R���SKJ�_I��e�ύ ,�������J���k_��TQ*t���,��}3\���j�3y����m�{Uѩ�ם����muD�C�YRY]|2�%+��D����o��[S���%`�Ag�(�%�=��T�9�O!� Mq(|�˷Z��`�65���3������3�A0˻�z^L鯴R˻��3�f���3;�A9Z��`"��Y e��m�Vn��i��9r�$�m��"Y}�Y43r���豬�A����ֽAM�񩝶:��]:�-�&�&w�7h^�ᮣ�H�/��)��W3fU�LJ�6�<��%3K�sub��C 5���i�zT�{{<0��"��t}���^�ه��Py_H�j����,]�VPF�=2K��*X4�����</3=�j{:�%ƅNY��e�����9��3d� (/���FI�P]����0/���=�<���8]}���tb+k+lu��:9+5����Y��>�p`��G��m��yi�֪0ʾ�k�˯
zN��]�cE�W�)��^$�qPm]Q$��KE`�M b�����g��vbҚ$e�Cg{Z��/��;He�G}����n��`{�˧��ū\1s���_��0�~5B5Nb�8ijg^0�;[�W�m��Ա$c
&&wؓn�!�FU<�z���<  
� 
�ˋ )�<}B�V�F�-"���yyRd畳A�:�`���Q*��]��R=��	�=���y����H���d��Qf�د�v�G�J�����ķ�̄=�L�,Q��r���e����g��t�w������T��羞ܻ-;y/+%�i��SD��c4������A��;|�?ޚ���|�@�Ǣ�
��!.�s;@�9e���Aă�fX
��5�.V�d�/3�|h� k�vK��8"\j61Vr���yew�O�($��Ge��wV��:v��`��G�/vȁ�%sW��?}-m�&" V}y�r$���EO\�9�?$�ޮ��B���'�}�Z�v�]w {���� �L(pU�AWIV�Ҥ Y?e�֐����&�|���᳛�Z��q���_{:�Ј�!ٛ�Hoy�hiA�fY���b���_FF&Y��!2XԈA�r^�5���wVˡ;���yky*��@jH�]w6�HD�pm�a��6CX:C�lTD*Z�א�#zɜ�l��_���DD,ڨ��cΨ��u����8���IQ/x4]/%��t�M�{��/w$�3�����9�n�;�$Cy�Moc��J�"���Ǚ�}��IS�TW�ř��
�'D׵>�f����)�0j��`m�M׺ub�NU�}��ٓ��Q&8Ѷd��=������^�LH��uV�U磧�\��z:RK���q�v����� ����!O���@V�ٹ���Z�����z�e��S&���,�+����+�N;lk�*�33c�iLć,u�`��l!Ѹ��O<��`��A/���[����/6wn�!Hb�|��7/yww�=5�T ��`  ��3���jS�BE������pB ��(X(N��A��sd����]}X��l�&�5q�J�U�B��A)]�����l��V�÷���W/l�W&�sY��D�6���z�:����y��vl��WP�_3p��Q��X֨��_i��)G̓���2=%�R�*O����ܔ;�{��.ֵ��ښ�_w��]�ɖ�T� �,�#w?b����S�'{R��D���epY�qxOi ��'���1�UjK��6��P��o��<��{���{�R��i�3��<m�DҊ*L��~���W?Ut��^Y�uLᬐ��@�1 �.D`G{�~̟����Xױ��3�!�۪��}r|��?V����_	����I�KN���cy��v��/���ڳ�G��;zu��n�Q7>�Q5s�:�� @۫ S���������/9'cS]m���)�D�=�8x�3^ʕ\��n��'��D��~�v�-d�|c��A�ϡ>-�6x�{@.at�]ʡ.R�����C� 
 & �)�:�{*��5�T ��<g&���zˇ�ʦ��t��/�;��~��7ȷ�N��=1�ޡU$��QT%�U�tY@;&(q2�|��]��;�P�md�}��V����G�堎����5;�z�;,�W�7\Uo�`��� �>�S�aԘ�so{��ݶv�T<@�^��E�(���-Q\W��"ÖR�΢�����s/�HdjA�c>2�$ PAh(�(0�,�@�`@@��yWY횤�*\�囻y*8���ET�;wk�w@ b�k�5 �Q$#B
 �Pp�"Am�l 	�m�H�.	�⛨��IO,��r�`�T�s��5�j_w4!��:L���Ͱ\ß�*��폛��?)sk���w���oX\�Z�0� 
�$���}wx�{����yDl�Tn5J����3�l��1�Ԯ�E���Of�8�TQ����bG	"㼡LM�wZ�Q��2��,\��&�̹Z* ��Y�Dl�Zi�1��]۱�ɳ[HK�nDL��#MbJ��W��6�uQ�H����Ny���o	q�y-�𸗼�V�����fL��z�nΨ;���?r�K��4� @�b_zO����'�|�į,W���� z��fե����
���Δx+Q�Q&&c � �[��G(��R�|��e�mv����j�[�W���ɔB��tsװ)����3�>�ȏ�F�\�-}��M�R~���*�+�m�������>.��DO=� �t��U1��̧��f�;�T3�=��#_Z�p[9���&�.��>0@:����t*�)j�+}3��{�J a= ����Վ0�U �4>�U����#�m�6.�;5�o�C-o}�a�=�l�X���[�k>GhTł������Y�4����u���?
��~B��7�zr�ok�E>�������������*G��J�kƣ����6���y�b���j|�W������K&��/��:��VPLu�Bgm�o�_�vW1R����*�ʧO+M!�z�@��J�FqQT�h�Vq�#�G5�bwJ�'ܠo�9��O�N���|�sb��E[KM+���
����؈7WA5-�C'��<�b)��7�Y��f��K��Ǜ�\u�ȂIg)!�r�U-0��U{��j�$��j!Yw��JtkL�:aQ#h�D�Kr�*�C.UHNL<���I�D�
�(���.�JI�
 �*r��.��ˀ�\�m��a*go�l27�#���Kzs���3���ﰎE˫������'����r��Aevn]6+t<����o;�r������b�y�����-��t���5|���P>�Q�[�B#�0{$�]���Ӳ_8����AE>DԾ�ɶ; [��h^��O?j斕"�w��'X�'K���JPbY��Ap��TN�4`$�2�.�P�fcx1\1΢{��8����V,�R�̜�jC5�ݓ���7q��,����Ƀ|t.�z��gu�T]r[�v�D�f���v�϶x�PC���i���U*Re:��mbV���DU�eԑ7O'2���Rt�E��[�`~y	`�����w��om��3N�@x�b�L2%�Z�sR�-�p�����v6¥ۆ��X�\��W ���5B�(aۊ�$a�G�iB�q<��v�p�,��T��|���(���r���܃^d�f��ӆ��;�ż��mFo�P��X���͕�b��#����h����Lvh��a����IV�<��}o������/v=�Rs�inD&v��ā�XN��;U=�nZXC�7'T����V�+�U�Ӵ�f��\5�C"��-N�J����P�z�vr��h���Ñ�+?Mo���ή���F�am^�W��b"v��z/�2�SD�-���us�R��ά�zP�`2_,��O*�lW�w�]q+�	+��2���Fݜܱ��uԛ9�{��^���!���+7���vs��;��vB�kr��Dr���#�]]p�:C9���p)d�����Oi�6e�+cȎ�9E6���9��לr��RR� w3�Jp��/:�*�^؋�嶀��hR��W&C��t���j��1�WB�Iu�P�(�̈́����N�Ċ<at�� \���7�*Tdt9�F���rn�o�,�v�&WT��|,�&�T._D���׌��Ve�{D���Շ0�iU�2�����n�i*Vĭ�Wɒ%e�Zbq�.��g.�f����-Ø��o�̌<
�ޭ�:�{�3QZWNy�q���L�G��N��S����}��+
[N���rn�ytm�SOW=�	��#�:���h�]Ộ�Q⌥/�Sꇰ��E��g(�	���wSĸ�<����Sl֌I���طI�zU@8c� W¡3T݁ �Bd���CV��.m� �o1	57��$κ��J�]�z����5D��!)�KܚV�+ b� "�)����6�M��|��}Բ���2�^���J�H-Y�*�[�����ɾ�91M�H� NN�+ڌ�^�D�u��ŏc_b���n�m`��-�"m��}�W��ZM��'|τ���ʼҥ��7���wq�;��äBP�iO7�Ԧ@4���R��d۝2��|�G�����n M�c�	\��<�ϕ��~�G�^�~��k�)`�D@23���U\��YUu���D�teb�~|�T�����[3�-�s��#���vJ��p|�a��`x��#^�]���Lŀ������|�H]���~�ɝ���U�"_;��F���R3`�/$���юK��kx�N�l\x3�����7F�+z(ڨU�ː��͌k��5���䗧�ʧ��B����JJ�7ql���.G�V��Su���w^�A��h���@q�L+Z*�/��j���TJ�q*@^*� I��T���8|�J*����n���L�>��F��HOW��yyM�Z��%�M ��>R>���?O� c D
�����4D��������U`8��q��}m�u�3cqj��OeL�1�F���O���>pR���I�a��ǁ�e�����jڷ�s�Ά �Q�����h�zԻ��<����Q>�k?]�^�r����y].���6﹆����
�`�H0C�! A�I � � ��f�7�v�ŝ�Q[W��������ܬD�h��/A�&$�t�)B�&"	 �I-"A �ED�-��2��g�%[-Iƞ���[�oe�`��@���=��*&�v�<7�sMH`�򶯆�#�]Oz3���Ά��'ZjX&���� �o�5�Va����n��"�sk>ɾ;�ɰ�$\�Q�=��m���<*^6�l�L��~�����ʓ�*v �����Fe{�� �c�u�t�	'��Ƌ��T�2�{ۓ��Pو�*�ckiޗ��^(���m�|�%���$N{�&�5P�����\�7�^�Dl�מ�Rgѷ��>1�m���	� �m| @EK��e��dɤ�=2���{�ֽX��p�?��;�>~�=��L����8�<�mxv�tCs�Lj�f�����U���iU
	-� �������X�C� g�o�A�"��s�cٸ� ��CDv�Y����S:g��8��,@��K�]x�EnE�N@�L�;���f�^�%�dkTT{8�侊���f��Li;�&���}wM��T	 `A�p	 �	&	��sE dۼ�=1�v&/{�Y�x�fҨ�\t����� t[�TIa�R3�1�@��N�,���&d-�5S
x1�����Xɋ'�/D�\�ɘq�Դ0@Viy�wYF.���@�=^<]R�gqn޶���_��}���Y���C���P���*�6O�9K�)-WK@��P*�@N2a�8�U�R@�?+�������o�#�i�%���"���$�L~�G���8��Y��~����t%@{���@�0��%��UB;)G�F_(���/��'KE���.i�`����l)b��	ŷ�u��}��Q�ۿߪ���ג� )�@��E*m}w2���Ͼv;������!A�l/��s����Ⱥ��exC�'r(�<}T���x+�G�	m�,a�(;j0��p�o)џ7$G
��}U�|�h���@�CYAW<���oR��MId��{�J�����1C1R��kؽq���S������$�wc�$��V��PI��{�//C�7�l-��h`<$D G޻�I=?Ni�Y��k7��/4���\�M�H�$,��ü`��b�H�d�˩ש 2|O�N=Ix��������!7���F��]%��ۇ��bu{���9n)�����wHD ��oc��dN\L��J*ۨpO
�e���l���Ӊn^� �f 0�!���UnT���YO�OX�b�}�.y99EW�q]Sj[j�a�p�ޯY�4!*�3-2j���&�6R���_,�_[B"92>����)ms�"�)� qjB�����&���h�?-�Σ�;����|�rR� o�2�Qw��*p9�u�Qŝ)�kﺪ��/M�3��>91 
�L��͚gG`��������� X���t��6�(ivy���a#����})�,g��R@���~U[�W��� �D�h2 ���b���`�`��3r����/���k�T1&Ur�&/�Z��iʒ�!%���a��t��F�����-�P����EvZ8��'p�p&Q�.��h�]�i���K�;�g����"���s�pû\x��u��VU�������X������hA���n�x���.)�(o{Ӑ$6�<�bṻ�-�V+�3n̬vt�J�&ϔ�/n����2�F�C��:�����[��j��=�����\~4��2oܹ|�>���@b�D��V��w�̋���z[�5��ax�Svލ��"'h��:Ԕ�����^B�h?	v��\x�K�5�K�dAf�QN�/�]��.~���^�
�3ga��[=v����i�Q�8e��qq|gv����=��r\��c�w�}�W�<�T\�Ĩ}= �f������f�g����܍Vd6J/z����S9��3X�ffo'->f��sӹ��us���D�<����.��t'Z��mz붟�к��t��VW���ͣ:��n�k�F�	ЎD�z����< DU�S�P��}7��W�F�g舏���Aיa����~L�ME���U3s��b�)��v���uŢ��0�N��6Z}�����s�3ßG�y���t(����n@\�}N���1� H) �A�� � ��� �H&"L)P14�*�����|o�8F��r��L��n�\���$�Apa@� 
(�$(��
�9�ԉ��:��\���B��isw.�Xp1�_j'TWJ���Ĕi6'GZ�4�>��d���*p|�=�����5咔��z�$�i��������S�ުay�#Cv�F ��c��A�w!�۪�]Ӈh�6�jK<��Ĉ�lz8�&jfI�le�;U�����_]�|�a!ί���gϹ'�f�ϺD	���%;F�Q�T.�7WT��1��2����t���S�&"{I��1X;�ww̲�-	^&��uX������eB��߿	�	Bu�^�2z��w�mz=%_B{�9ZZW�nqX����� ;���^���\�tl[B�n2y���a���2��mD#{9����oz,����U�/�`c��Qm]	��t�����Z����Yt|.U�Y���wN��C2�um��/ZOjk�ɋ�N�z����y���N멝�=� ��$'��������e�p�d,�Y�Q��˒��èX�[�)�qow&v��[�P���FB���mvy��W�y�h�t���Xh��1�ȑk)�D��g-�32��ʮ���)��-�3z]�/��U1G��dn�75[��}���P@�狳N�]z�����,���X/���q��	�?�h�(�@f	�&�ؓ/�q>⦻��ܪ�9ڞ3���Ƨt�#�hD#����gn�H�D�bC�J�g0���{zb���i����+z x��b��1>Wçj6ާd�.����>��.��yG�� 	�`;P�8;�� }x�-��k����Y�s��xOx0�c�z[�|Eα	��P�5C�����=�JD�>�W��+F%ҸMV�������]��4�6�f��E����ƶ�?��z�;1�;Ĵ=&L�u�ݴfO�-�V ��i�����Ғ�y�f��]s��L��j�Y3R7�����Bw�D�l����uL`�U�"�$�i��I��{=w���~f~g��}
�N4�9'�V0_py�6����8QM���T��;��n�莪Ct�������{C���t�:�R㯣Z���f���5_�W��_?B���h�" ��O� H���ú��|T��@d@��L��bʗ�i|5"�h��������z�Z��q��ͣ�=�o��Ku5�P�$>J&g�=Cӆ���U�_��`�Ȉ�[�dY�7we�ӏ���"߸#��q �6�y����o�}���[9�=H��O��,��T�/�a�]g��^���r��UW�9R}�5ci�J�b�Xբ�Z��Єi���|���<�8ǽ^�MX��C��)��@�$�������dHC HWֳ���qR�VLp�����
�Ί첿�{������u,�,���Hn���><����:��JV'��qY=�\iJ\x�KΚ{k38�������J���|�ӡM������d�#&�ɇ�y�o�E/u�S��I��TLj��3s��Ǣ���,���fy;n��	 �A A�$`ֻ���r�2���Ze��O�t*�s�Q!^��C����*�I7ҍ-~!Ģۖ�v�+�F���(ak'�fv�3���rH -�������{7e�f86�^��Fy	�.�O����XcIi��otn@�+�vGj���l�/u�}�|I��ڬ#���W�I֚6���֟�ۏ	ω���7�T�i�C�p��=M�^c�Kv.ۊ��\|��8�ٮ�QPF��v~�Zs�w�>Z�^�̼a ���>��`��ƭې#\�}7ᕻǭX4�[m��½�L΂�E�e�5��KQ~��O��"�J�w}�m"�j_�T�]��r�}�w��Lϵ/�p�"wgh}Y�UCe�݊t���FV���]@�GK��0Z����=7�"X���\�ڻ����F��g�y���TF5���{nR������O4V)�:a�W���d��(z�����]�#;E�"ogMN��&>U_����j�%��O<o��۩��p���D�n���K
���U�VY��@S��3�/P���e��b����nvNk�K�F٨$.�qj������R�)2�3+V;q�_U��])k9��n5���Wӛۻs�a�}�51��  _!w�#��p�˩4C�u�ofd��T�\cxչ�5��r6��z'�+�̞(YE���g]�mW��+I���oh�)�Mi}���"�X��{�xgÕ;��<�G�<=�)��
j~WKJV�!OT��v���_������xj]Qk�P�8b�6 �T�Ɛ�]$4�7��V�%]_��JSKެ���(d�4@+&۩!>���W�:[�s9uЯ����F8j���y��Ła����˰���Z{Ja� 
���P#� Cwg�.�\��a�+�q4��y�VT��v��kb���-����z����*E�3���}����|�`oK=�ϕ�����]�;z��~Q�f�@I��x|�EפҦ����f_I�Ob^R�>��RTȕ�t�&_�]C�1���q�^�N�8�&����G�G]�};c�R�\�}{~�s� f��~���COnD뮦{�sWA���UF+�If Y��XY�g�0��3�g*�ѵ�	?E�l�hz�n�.,8��c*eG�X�^aD3���O�M��;� b@|D�4�(�L��ṗ&l�#�f�K�y���^J��F�� �P�noz�S�x�
��Sپ�K�du\���z�]5�|�oe8L���bs'"���}��H7�h}8\���t�KE��eA�-m��Ɯ��ϻ�ݑ&!�M:���>ԩ����� w�[�^ϫ ����ֻdG�zᘿ�	�����+f���3�*������D�/\�]c��<Jԯ%B�����Q29�9�q7����Φ�P��y����' E�>h/�i�H��ك�ÓٙHh;��OF~��ⲅ�(y����E��3�Q����j�Ǿ���;C������ρPϩ6s�$_����Gр����9@@?t�r�:LhVo��|/�u�\4�dUx��!xm�x7>D����ٍ.l��\0}�FldQ&a��b�L3gf��M�^���� �>����n�ݡ�:��u��W*0;��I T��4'aP䌩\���a>�'�:+nF����q��sC-��w3T/Y���D�^�V�aR�rb󛧻|ލ�EU�*���P����/�j�^�eA���p�į�1җ����yKiL)���r���n]���Ø���b�&�*ANo��@Q�
m�S����. ,��f�)�e�J��H=nN5c9�r�]�}s!��� �����X���E W�K]mo'.�ʅG��[��jYYb��P�}�(Tĭ��ĘP B�d"0Y��C��Jg9[�[D
[��"V�j��f���D�S����}fb��l
�j��c*��;o�����@#�v�E-6H�#}��w��# �&�k�{���V��q>��}$o�[\�/B�2=�#�H�k����;��4� T��{��~O��_w���sҽr����0I0H �T(U
���ކQ2�F���HE*0�h7�q�eH̏	y�5����
���0º�L�ym���Wz`��%����A\�quLAy)����<.�p�{b��޼;���@#)�Z�[���wq��jX^7�OF1rPѨH�����UE��&���U7P������T�wc����&D�}�����pzO��NRϟ.z8��N׷sے�b x�`�X��@��l��߇SyT=�*�j�s�t}<q�x/�%���U��v4��6��LJ��xd�3J��U������(T_WQ�|��py7��y��." ��k�m���DE���&pZ"o���y���gA��z��ԭ]��9UC�.�^�t�_�Uߝ�4]L�z�Fz��q�@�:��&,���@{�z@�GlϪ�+n-cI$��S1�z��O�����s�%��d�gȂ"ڇ�'3Z�!���5L�u6�h�=��0��ߋ�|m�����������_�E:��A^��~	�d��H7������ˌ��V �6�UwR�bZ�*�F��0wo2����A���"뵝jfa����h��6R��2LT]�jL۫	�8mPV�=a�U�?cw�N貶c1 iK����'*��Gl!�8c� P\6�EU� dB"U�4�:d�"��Q%V*���r	 �a��,T&��T��s6Uᗺ�f�iT�Hv��T��Zl�]b*�٥�v�[37�d>)a8:J�L؝�@c�.�K�؜왇o�3�i}K�zE'}qu�yf5܌�{�I�⹙��d������J)�)��a�%ͧ�艗�h[@ �+��ݎ�:ge�m�sc�$k�c�懓�t�w1Kzӣ�xoB��ϩ�Nv\n]e��l�45�k�bH ��*U9���N-��!c�
U����T�҈v{Ugj���\�8��
��	��7��{�c`쭊a�����4�X�m���	��쨁���q�y���(����"�K��d����U82��F:	#�U�Śmi ۽��[��,ݧe�P�߭+K2�U�f�:1�[ڳS�掮]�l�4,���D@o$�i�f�Ш�wط̤6/�])�z��u�j���t�P�Zi����ۘ���$�[���'P$�c��]�[զPf'���X��`�>۝�M�s�)�M-
�ik��>���I�.�J癉*Hl�_[޳�V��/u�Yi��}mu�RS�/ ������g���g4-JҧY$r;b&;s�6m4`��zOs˴��9%�G��^�o���Үp�/5h��a�l�zʙ�<@��vL��`�������	����������[�Ҩ�F�(���������I1Rt�,V���oGrNj�$/)c�@�^\���Gl���\Hc��U�ô9��.mY�T�P!Bk��s��B:;���бFԎ����j�l�wY�&����͌�n%�P��<�pÖ�ШF�bL��{$n�6�A����G�G2�wNO��Yy�S�=�zw[wH�"�f���;�O���U=�|S�u���v������`��:Yr��%���
�}�������c�2y�I\�Zݰ떩��r��%�o$G`ٹ��9h/u�_^��˺���pn%%������������s���1չ̭��G��WLuWwX��`�Nns����#ul�(WR�҉R�����xu��ҡoZ.VQJ�*�EΥ�mu��U��Nx��ׁq�B�B�頍�[c�;?��a��6����@��w|�oL��E�5c�:Z�fӎ�:A%�\z7j&�c&zy��j�񇕠�u:��B��	i�т�fV`2�[.M2�\��6�ԲM�{�o}� 2,8������;����<�8 l�ah�/;��olЦ�?����,��ܦàM\?0�o��@��ʄژW����b��j�]�ܲ�KO�nGy�85�i֔WC����w�;;����S_�͓�a������O��r�{ˈ���&���Nk�+������)�^�_S��߾a]5���u��]�wP����癖���2����fM?r� �LFK����R ��y���c��MTԎӲ̫]�[�]r�w��.l��fm{$o���b�w���v���d;��Ǜ��rP�n0�(�k�W�߇�z���T��H7�1�号.v<�s'{������7�-��ّ��&=�PI�)�"��݋�n�c���/�Ⱥ�}]�/�{�zxi���(��[�h@��20��4(�4�DB�f���\����$���8�b7��}}��MEQ�7+�P� �i�iH_�Փ���:q:��#��� �Z�'��ll�<��m�o�sX�q>��d�"��]�2.kJ+3Y�����;lŗ�وd,![��<Ɇ�@���x#U����m��uVI}��(R�� ^��=�.+�G�y�)j����pB�H��¡����{%��_U:O�h�;S�Q��������:����j���Ҵ�_���L��  $�@x��ۦ}Nr~ś)1�i�m���ܜ2e ��$��4Sh ��%	�k"�Y�}�Kg�\v��ެ��T��oV�"X��f��3�wR\�{&�*���Y�� iC�CʍdD��ٽ��їÐ6�Noa����4������(�v�m}V�������<�/n:xz���@�f�}b���#��Z��N�u�^���\�<6	�~�)t�F���`�_KoDC�Z�Sa��9I仆���-��5��o���9�Mvc=���D��<y�b���KXf�~�7�.�VM�,����Uܮ�ߙ�-�)r���xSs��"s^-�||�mu���ĩΚq6F��U2~�b��zz]3��0�n��{���d
�V8n�����MU`ձb ���\����sH�cXܮ<�>�1q KU�?W�h��|7���Q�|uӳ��x�p���.��ߨ<|�����SG�I]�%j;�[��su�U�ɢ!��46̿9׈w��z��ʪ�:��'�*j,��@:ߍ^�띝����4Q̝ q�q�f�n,��b�
�[�`����.# �^��E���YU_���n�Tu^w��v;�}<�(>vM�ݻ����ԅ�b�~��,���9����c-,�5�;y��J�S0Z�����>�֕�pp!��'�y|Qι��У���D��V���t���J F w!PMV���)�ʈ��P��w�
�x{�$��C0�� �ѽ��փ:�(M�`�����0ؘ+M%�_6�t���r�����*����kjQ
��S_,
�L7O�-b�8��z�f��K��h����)AŒ�Tz�.�x���ZF�b�ϧO}N^T��3^Ո$������V����0<���w�j�Fq[�Q��T�
��J�xw�SS�q߾��7 �ڗ;��l_d ~�R��qt�å���ք��J׶D�ы�'����<H����z���L�7�?���FNЩ��y�#�o�b}k��1�Kc�j1+|��+]����kQg���^�+nG����|���ݔ�NY���������F�M��hs~�W�J_��}N�K4`F�L{l�%�����'�¬�p��,Q��:�O��f;�P�Q�ȟL�ck+`��36���ʹ��u���8�VJ�j�^��2Yy��m��n�~f���kg;
nW�B���s���iͻ*j-���z��{E@��n3���H�6�oiN���?L��r��=�xT��>�B�UP P$�$?Mrϱ��W!�|��®��Y�%.�xt<���6�2v��媮�bzIاX�u�L�Gm�m�:Dx���g��C0�@B #� 
����h��rJ���`8��LA-������R.	��C$ѣL�b��j�>6gT��:9q������}��j��t՗��ơ�1Z�]����\�����K]KS��lք�3��}�7"�-N�_���c�=���;�t� �~����x��P�բ1^��>d]ۧ���rl7:͞V���3�Bh��KW?S@��N�;md���ׇ{K.���bxe7��K��<\�mZl��Ù��c�B���h�3$"�B��9��*L�meu�Πw�\��&�fji���5XS�ٞy`:�� �����%�|�7㶷��H��"7�q1�<��.�;z��$�Lv�^h�|�~�7)=m1pw�q��q��`��e�'GU����\{���vp��}msG.&�s;�g��`�y�]E�w�5(:�w��j����a{��ߜヷ<�N�۷$ F9���/vT�m�w=]�lM���Ճ����@���[x旔��K��U��n����wJz� `�0H-�R��R�n;i*۬���n��RM���;��BF�`YW:j"�)�
/��3'c���@i��0����:.��w�x�A�>�)��#���W&�)��7b!���߽_Z��S_ �D ��D\a�h%T[r+�ν�4e�d��b0�����*ۿ�\�<j���yW���r��H�W3�$�y;B�����H�1@�
��V;�\\5=��ɇwc�Wi�أ�Ŏ��D�� %rκ�mX�yܳ r�4�VT�Z����Lr��cv��\������VD����`^�t�yn,{z�#���$�C���-5̴���@?Z�����Fw�������BB�U��~��� ޙ|{��A��!�yj�~��3���2�P�~�ͷ쾥�i��S�O}�w��q#���!�v�Slv0�7���v�n0����_}=__r����a�=o�#Q3]� �PR#kwh�T`{���S�0��	z�dMr»y��r�H[���&1���������T���!������f{v��8�uO}�VT���w�g,���>�H}D�Ĵx�W��\W�h=�����d͏�4�?�u�� �j�U�j��W���ԭ/גA0�DSN��[SHә"ǔ����7G��	|�'�;��˳�y׈���Yg�]*f�*���M"I�˃{�{�A|�бq�#`��*��/%����^f���PK�eM`��h�v�Ŀ��IrQڮC>u5�왓M7�Uk�sua�>o_��-;��K��`-R���o>�Vb�R8�~� X�S�^�	B�L D  {�7�_I%�L�<�Q�6�p��:��b#9����( A$aF $DeU��fg;[���t�ՃhWz��Rgb��-:�����wx�3��v�K�vgZ
�ܚy�5���ׇ�	M=';]����N������S=Y"�6�[U\�S�Y�W!�*����Ϧ4�a�K�96)��k�h���NXd���S�S���Ҭ�s�%;ɚ�C��R��*��U9p�A?�K��*^�Vz����-�e�>񒭊�7~��_��� �#�y���7ܫݥK�=�w�;i��c���D�s��$}�o�ϧ��e����u�F���7������v�wY��x�����0(.�j��y�V�5:)�>_m���Z��L�P�g�Dp����w��*LԱ��+��ܺŕn���V3{��{��w��VW���W��{  �x'c�І{,>�WDk�S(��2kFM�*�r%U�b�kȚ��-D�L�r9yGxu�r�D���!��Ћx�%�K�"Z靻��s}>v�Vff�Ijz��"L1�k��;����Y�@���E#!�[2��J�]�?�oF�o~��&b]���mn�&fΫ��<k<J�tX��s��/�	�.���,�$Ј�Ksw�=�n�Q���8U��Ӕح�,g��3�΀����,s���ɲk��H��n>�O�����h�d���u���wnXW�p���[:�\�hX׎Ս��5�"i��7�(F�u�ɤ�S��t�l�E�CGhVK�'Wq��yR{0ΫO8]���0��pN���e˭a�!�����B�3|�!�5fӂ:oj��b��ѻ|Q������h�������Gٝ�q(�_K���f��{��
���'��Q^����y��h���w��ִ�
cG��� EO�
15;N�'�BX6g�8�����* ���E�����l���ܾ�wn`�>}��V��ڒ�*o�_���-L]�*e���K+�x=��S�{F֏7�����r������#��õ��m�ﭛ��ӿ)?M�:��t�]��	����OuQN��,����Ap'=[�O�Q�����_�������T�[�n��Sr�R=�p]_�ʐf\�J/2�u6�LA���(a63�_�1Ӎo=��0���~�}1&��a��{ڦ��͗Q������o<��;�v��0Y̽�q �0 �M��}�{S}}.������oq��ݱ{���ݡ�A}�hyvۥ����A�@O�zŊZD�u�Zc���[W�<YWw&.�z��ם��nM��M��AF��@d��ꥬG���r�RH�dih�u�c6���`�$ML���F���]�q�-y���]Zq:nPG�C�'hj'�I'�G����n_p���xk��n?�#ǎm�����,K�3��1ͨ/�,��>O�|LϞ���v�3����S�B=o*.�v�cv��q�|�۴�dϛ��^�<��4�#o&W-�5���ر�S�[]���Y���S�7ۺ�4r�zP���9|P���< #m�`@W�����i��j�wN��2�|yE�z�	}����)�|_�F�N������<�_�픦����$-������ � Q%�_�~�/�}u��榵.�ܳ�u��q�Ǥ���Ւ׏-e�m�9���_Yc���tk�yj��_(���Z-_m����{!. 9�v����qr�7���{�j��=��S���;$F�8����N'Հ�ٷm`p�k�jçnn2��"�� K�I�黲�,�.�8��k��by��,y����*���W���gUL�ө�
������/Lu;Qi����+s	[0��-���:}0LE�9A��AG� �J�u�������[��]�JR%fa�C���A$��$Za�A� �Q�x��@��cגP���cڊ�t%{'��r����!��گi��rq���z��+�{�#�-��Q�4��6�-_2���yy��W6dy�v1[��M�\~� f{�������N���q
��V�^Z#n5k�S�v�_qʩӰt�nl�)�d�L�Hm� ���`O?M�7�n^�h��\�5s�sKou�ed�Q�]ݠ�V*���h>�̍�Ŋ��.[b��殌��SӅ-����v�uX�<��qs��Cmۿ&n{��7�I�åՙL�o��u�`�2i;���e�Wi�Ɇ�}����`%7�*�e㭪����7���=eg/��������"�����V����=��5]�<Z`&��aN����V����[�PY!�!�3d������nQ��~���B#�D�Wo��׽}��f�k�6Q��x"e��2x�]z�C�
૜��l�������;���1n������dx���[31g�����K��6H��Ug;l}u0��L<M5�n���|X(���Dl��V�}��8�x�؉#�@� �"08�Yu-M��� \�U�g�eҗ<RAV"��x��|h^�Q�`����x����f��zַ�ư�n�DQ�+4��Uׁ���Cgm�*X<e@����ײ�u�n��s��ŁՄ]a��I�Ӕ�a}�wɻὢ�B����S3H��a~l���#�բf�h�0`��������ڷt@���iő�����~U��\o�
��~7��X�:7��Rp���&�`�������]��{%ۡ����T2�)�����e,�;%�9"~�1�EL}L����aj�@`s���m3�w�$Ru.��v�T�L���yq�Y�+��9C�B3�z�N��107����k�v`LU+�-�j�pO&�4�h�ۆ	K4	��;x��ڋ�?
�$	/��JML�$�!����:۪�z7XB���۞}�g�jVf�����5���S'���_}3����5�,�:['���T�L�'���4�r����i�kf�m�2�_Wz�Z:6߶��J���9�m����]N�i��n���g�o]�藟Λ�fx����Rcf���䴗���$�t�fD����4�&����e����[����4%=kM˪�'�"��T]��A����U�]�Ƅ�X�-P��@�9QIU�ʨ�tҎU�x��N�JIJaZ N��%��e�o�����֥
W3+2���h v'h�Ld�me�fj-#d��/Ä�H�H*XX0e*Q�� &�i�2&	\��Iف�!���C����������V�@{�ë�%.��MY��(m$��9:���
�M��v�ki[�ʇp��ǳi*��˃[D��j�0�������ؾ��)��������~��6�L�If�r'�B���r�n�+)�5]��1j��i�Ք�����Z�]�m=��rQr�U���Np��Z70�*��w��:a��F���9c�f
G�"*{�+Ͱ�Yɩa��}�n!����;�b&-xŜ�М�T�����X�,�)G��Ɉ_<�6S/X�9ыY��X��0 ƀ7��E��-��93nD��$��,�zB�n0��C �d��6��t�)J��U�d'��jsc4ji
Ѹ�I=a��'����1�D�p��];UR��.a�cټn�����+�I$��"�]RDhA6��r��eZ����*���%��r�V��ʙX1�r�b�j�����cq�s�}|��8+Y$ё{[�X�t�]uWZ�7�]e���'
�w����uVp�A`�\�V����J<�����'��y�F��L��NU�vE@��l�2�siD��V[޼�HC��Ka�(�Fq�*WmmJ�P[�4���c-hײ3fk|��k3��{vFk�S�����}n�]S4_N�V�ͅ�]ޣ�m�u���&-ڕ���ƼY��
���,&���Z����M9�B�Č��mt����|C���'���M���z��]ڶ�wj��m�p���Jd�9�HU��S�Ngm�)Ӵ.��eEsjk�E����y�i`��V�F��}F�C��Ę�ծ�9 {����ң�������yyH��{���UwI���ϣ\��A��.�[�TJ�88qY6�L����M�-��!oqZ�*��!��\F8`xp 7+6�l�0Aտ��� C6
���k[��N�;N�&���[�_.��uf'}�ĹAh�X�ұ�����;�N7�$w)EW�'^55�^�L0 voR���[��t�oj��Y��Q�����(����۫��r�%W	�m��r:��Ӻ��nJ��VE�e�`�B�f�S�N�M��4�]&�1Q8"��6�Gx�[?s��C�"$N-Y�����Wa��8-��,��n�P쭔��E��6�]�Ǻ��pC�=VMU��(���Y�g"K�f7N Ћ�����wI�T��\�d�Ka5�溻�h>-��&�n����r�^^�r�� �J��!*M.�#�jJK����;�;ݺ���R*]4<�)eXT�ĝp�n��Hd���g9���!vf��y��"i��n�%[;�T����jN��'�RN:���T�d���k˯���$��̙�����J����ut���/R1�{���j�
�E����:�nʫ6[i�b��`t�ż)�~��g˔���������/�zg������`{�B`�*���=;�Wﮚ#Π2 D=������z�n62	۶�T;.Yfq��׎�j�}j�u-�3{3R����9}�}�ڽ��)� _��?x���^���o%��O�_x�U���N=���/��[�"�y�Z�C�p�Eb�}¶\.�}����oi,��b^
�b����'�@��{�sr/5�nfV�e�~LR���:���F������|xcr� �>����}���k�n_}����73������do�.O2Z����wE�}��4��s��"��_U�=&���'̲zj�����pL
zÕ_[R_�9J~�NF��ly�,�z[��uyz$�Ƒ
K�s��,1���H�[�����V���4jI2�`��pq���V�@��G�]����1�gK��I��=O��у�sf�я�,�R��5�Ӡ�H�,#Iǁ�����=�&��J]J���Q���q����A�9�˱�������).��ܾM�h��,o�������Η>�3���9�&�F�l*�@�D��yK�|����>��~�i�R$���Y���;m#y$��M�j�Yy	��������������N�i<M]��s���0���g(sÈX;�.�M粑s%������(��ͽ��|���ɼ1�fWWu���@x�u��S϶�è;:fV�kW_dO�X�2"ÛW�9Ͳ*���lv�$�cj��&+p�B.�
`�X:&�;��Z�z�R�#b�M�Y��ue]@r5+
����g�M���[��^Tu�eض���{�"y��.� O�]v�:&~Κߢ�k\�&����R�غ3�*lT'6]��oc������;�j�CRs�W��s-;���K��-�c��S�[p�C"	��R� �.w�o@�6�dZp^��1Ǧ��j���e��t�Πv�$���Z9p�u�n�1��9��N�^Uŝ/��pH�G�8�3�=��:���F�|�zI�W����*��� @�Rv���DD�8suP����0H�KpG<�r�����c�P�]�����;�I`�ؔ��q������73����������o!�Z��fFD�=r;w���y8�O����3\Fn���L���{��1.s�h�]�?]zgT����&��Q?��ʏyZ��-L�����i]��̸��Ձ��a���uj��laƙ�+>]ӣx@�o~�!��;�����α\��;�3�?���eQeP��T����9T��3��C�ʂ��j�SQ�g�MZu=�Ǣߓ�+��vo��Zً0�BqQpm�4�z����3\��2�>)$S�f�=>�l4�Zq�J��g5�H�6)���ӵ��7SE�H��.�796�9'�٬�|�i/��X%�)�Y(c�}t��Wg��S�C3S��w��\�b96��Gr <��F���	���tL���n��&.��wC�ʆB�+�x���mp�o�Ũ��P��(�LA�x1%j��{��}7�P0����}�M�];��	�7�c�ې���U��j��9]���훙o����'�<Y���I��<^5}���?H]X�>p)�'ݺɺ�a�	�2𣉮�1�FuHc��kYs7�#��5q�y�U�)v6�엲�f'E��q֥^��{�O�zK+־��Nت��S:�%VG[njl�i̢^�4��3�r���\F�'JZ�f㝐Kk�s�2�Ƽn��s7e�xF�e���2}_�)�zF���m�����7e�u�L�{�/�oj�mP�[W�d�l||[��}mъ��w_��gCQ�R���u�FЖ7�l%�ɫd��l��~�g��������T��wd��m���n�o�E����y���No��<�c����2���W�7����" ��V�:j򼘡�%ª����E�ϣf^?Y �@m��u�_[\��S�6cr��*��3kt3t;��"u��4�o�Q+���Ź��5�R+���Uf
:�������0!!ҚJ�pvh����fu#�+ww5n6�r��Xu� �mv��J���u_���<�&��N�p�����h^'ݯe��ʜ�7Yޜ�����K��*{'��Y������f�gv�w$׸�RѲ�:�"y�\���װY����>�C�_��V KGn㤐����[����Q����_��֬����4	������_gt�`�դj�}o��y��*v=pس��ԑ��;��d����o����@o��:򺈪��bU����AK�򾐢0 � ��{�Vg��y�K�N�b����Ǯ�[��Yr�[��g�(��b=Z�ηkw"}0#hGŮ�*��!� T��1r���TA!�[�I�MЙ��ɕ�c������rg®��t.sF��v0���0�� !�[E!���\�W6��8ft+a=�_�?_eq��V�M;��8耸E9i>t,�#;qJ��Z��+����5�S�r�L����v��yz�a�{�6������]4>>i�����[�����ǈR��@�LD�]>�ܾ\ު��s���Q��2�n�]Ki9Ʈ4�@��lhh��hSyKn�s�Gs2�@Ud�������m�cT�`�OK�a��Hڋ���j�TW,���GQUƑ\-�o���Y�����ow���J*��-� Ih�Уbz�Um7Jw��|��-��^|�g���Z� 1���\��&H�+]Gz���KF]<	��4��o��6��.F�n0�mNW��T}d|�[�.g����D�].{�y�f�U y�� `#���.���:�f(az;�ҫBӝ{�`�����L�.�Zέ�M]�nɶ�����T_���z����˷����2��
�)Ï���2�x�ͻ�_	�om��������y��C��I��}F�[��C�iB~��o{�̚��;oI���d�XH����os��f�Ct=���-J��/%I�}{y\{sa�Y�Ԋ��87}t�79i�S��lfهf���7ȃ��\�%��H<��q*��o��gD��}��yM�^?C���)-�/H3�޶�����!^��Ay����35~���L7�9u8���OrS5n��ww�3j�L@�@�(�
@�`�!��6Y��4��՜����f&��ɳ�v�\��6�.��'�Tm��+i	��k�(o[[aH�X���Xi�8�Ix����k��WN����L�GU��d�z@@��I�z�y��y�W'畎|�*V-����g��Y'>�>}��}���{��w�� �M�-���׺P�5ׁ�{�'-�݌:��	�����{=6�Ǻ��
Q�_Q��vzI]�k8�{=]��0T�/�J끼 wW�	��,UR_�6�=�,��NO��2�����꿾��<Ө��&�I6�����og`ʽ���4;-fO3��z�)����ӂ�9�g<7���<�!�ܾ�u�Y�>�=��*���㊠��+��­��N3_ 0�e�B ��w�|m9'����U:j����|�r�~�/�V��I�?){��-��Wn���l�����έ�*�u�g7��]O�z���G�@�>s�!��l'���3d�#��~��w ���(���ϭ�r��CE{�4�`��1V��Yg/YF��+�[4kj,�S���U�:��x�@E�vg8/�3��P�w�+om�o�T���@'��aT��L�m���N)�쬽��������YoR���;����ƦT�cl�F߷g�ܝ��Gl&Kqcw
��=�,��{2���s=wS�:ojW�.n���s��U����N)�R��,/LEI�X ��Z��y�۸��� ��x眜JF��Y^,��>a��a��z��m��^I�Q*�xW�+�"��h'^:g�ϖ�S�^�(���]��OY+�߆vT��ж�w��^�6�K���������d�I�Π��>)�j���$��a�otx�	�X�}��f�0�����>���^�%`1�be��S�*.V��6ŉ�6}��<݀�l�fڸ�ghnu���\���c�+7eĽg)b=r�1��.],]��RՆh�ʑ4��V�Lݵg;��6k�5����:�~�76YEQK/9(%b"븓�n1]�w�5��=lx���J�X���m\V�Ύ̎�q�-�U�z �t}�y����}��:~��0D��& F u�~�Lf"*��Z����wR�j�s�fL�RM��!�	�`wԛ��!�f���H9��"��k0\�~�]κ��4�@z��'-|�?���\��ogH;5�����P�9Ǡ��J�}�S���]dp~߼�|�䎯s���ߒ��� 	"L��3�{�}���Л�Mǎ&#���r��MJ���,.qm������=Ҹ�[qϽC�`Ѕ���M���������dJ���{��	�����Rt�|=q��7��%��ґ��m�f�v��s�iX��\�$WhF�??�3�G������~�tg%��0���Qv̙����^�{]�E�3��[+r}�w��3t��͊�gZ������^��dߔ�i��94��|��3T�%��'�bk��m����!�� ˯L	�7��U������ߪq?_Q����̵��J�釹�S'�ƶ��nj�M�~����P��?�w\��y�f�m�Ek��I~���F���ؘ��ˣsw�.�I�1W|hDZb��H��v}f���@Y���t��Րa�Z�Z�wr)M����a���r@�Ht� �s�
ݚ9�v��"��5�L ����_�^���w7ӉΪ�;��9u��h�Lhw:�����
��&��^L��Kv����0�i�5y���Y�e��_���x��>��w�������Rm��X������v������{�k���Kl���� �7�3v���3g:�m�Am\˹�ӝea����wgT�9M{ӝ��.���[�����X��>���k�c����GEu�:Y$M�u��$RR�<UŬ{w�g� zϘ���df�'K�Y��������	9���H����6� ;���z��Υ�S^k7�ׅ�$������x���2�����`}���uOBcM�Għ�/`d��6��S3���c-ᣪ��-���Q��DA N������`^���g���;��yE��}�`��g�qʅ��p�Uō��rrȫ�l9��LDD.���"!��J����Dsy�c���f���\�����k���ޖJh��N�Ʒ���l����*!ŋk��`[�!�4hF*�L��I�]l�l�ZoAf2�6F\�F:�\�����h]�t�3�q"j��Ŵ�U���1 ��%t�ݝ��Ɓ��z��c`�ӂ򰼛�D����e�.�_rw�w��t1�M����	#s�N�z���0Cw��\�(��T��a,*H�����.K���`ޓP��"�-&�~ ��VX���&��u	{�%u�=���ɵ�	�q��C��m���4����B*��71��uU�]����N;q�;Y�ܩ&��]�ű���
�
�ue��~6��/yp���[�<U�f*x��j���uԭ��o9�Pգ)t�V�6e�r�Y;�]�T�MM�a��3GMƙ�2u����{j���h�i:�!��xF�Q�� �nc=\�n�vv\�)p�ޝ�8I��)�`�z��+'E��ҕ}B���oMb�`KW��A/���� �N�f����a��V$������+��8��N�{ݨ�	J8��A�5A�AOZ'I��$8x4궪�l]b+$T`I_j�ٸ�*1e��;hi�݂�a�V��(��5��*�S�M(�tZ���:#t*�j���N�e=j��I[�j����ڜ�܉]���*4��$�I����;U��z:����z���ncOE)�q����v~�H�`t���V�4�wKI��R
|�q�.n�Y�n�⫘�>��ʼ�����W~#A��G��Сk�N�F��H�H{��XsѝǸ�K/��|M��V�0�IΦy�np`J�ɭ��G�Ys�o:
��G�ݑ��=�*��sa��9`ؗcĈSbܣ�ص&�����F���/�]c��vA
b��DU�w��������[\^��K5���+X��;�v���1���.]s�����i�2�cD
d�܄m��/��b��&+�f��P�T����uM)����4����g��//��2��	�p�4�tRc����k��&�^�	�K�wR�q*H��{�t�M0��Q�a��*Nwwڴ��5;�Ś۰���Z�%Iݍ�k�&�zj�H��(���f޷�fB�h+:�a�Ѹ$!��S�������`��ԣE�*��٨hp]�*u��0+m�_6�#��)��V0�s�J����S-}x�n"�]�*���4��]`=�R�r�j�ګ�tH\8au����+��2e�R#MtH
Kr�v�;y����ʇ���a-��
ֆ�|�XŎ�\Va[�4bS�����Im�qVq�7�N���s��Y\�mjPCD~}��M�4U��kr_���������]8��rt�woL�jˠ��֯���uR�Ǽ����m2��8dK��K�ifݙ�����aU���^,�U�$�T ��A���5C*�U�k s��:vػ�qΠ�3�y�wii�<ΗOD��̙N�k.�G���ݏ3��ف_L�j���4��:`QWv�e@�1�g�4�WW)�"�I-w4r��Wm��xL��w3��B�۔nT?~�֝���V��X.�i�ͷc����ʍ<�gB�����"���	�|�D_q�P�N��u� ��2z��~8�������NcFsY��A%Q����x�5Ҽ/�g��{�p)���d���szc�Nw�{���~�C�%1ӈ��|�%J���o�k��n�)�7�ә~
"���]ӏ�`؛\z[����hKW;���$en�����&n��~����ũ;�X�9�J�w1�u�΋<G@�Nw�����^�c�[E�g9N�e@�fr!O����P��ϧ �?��&\{-͗�nz��K�a�������l�vbb8���1x����yX/M*�����nww%�s���|�Y��E;��7j�
��f<ʥ72s���-�:�ת��." }j" �L�o�}"���	D���b�g�u��$��O1=E`Z��V��WuY�����o
0��r8����������]�ux�-�W{��ʼ��{(�B�ˋ�=*�[$� uxj�a�]��)s�{	mQ�9�*h *��hw������ÿJ���x��'ã*�o��n�szS�F]Uʖ����Lf:����6�����&"�v�r�.�V�o���_��}ۛ߻�ϩzV}�B�����^��C#%�Vӹ��v��d�N��wN���U�|�N#��:�`ʖ�y�*�ӄL�n�B�7΀��gZ7Z+A�y�2�n@��Yn��x��@�o��6Cev�;�u�]���r[�w�;�t�8_�8�3
��A��:�A�vދw�$���2�St�c�ˎJYh|��kl�@M���l���(ހ4J�yw�B�w;���i�G��7K���� 3���V[�/���C����ݹ����7'S��^M��'������tߟ��b��¸*Cp�D���dn׻Wf�_\��N`Z�_9g&8u��Z��t��?�D��&P��(��m:�O^R��2��VnҤ��ף*Ѣ8Q��<3�A�# ,@�a��$$�#[T��J�\6� n��V��5)s��oh��7ư���%��-���;�����P�}9M�)�K�pn�n���w��8�S�13��>�˚���y���Z��m�Zd�5�fͩn�ȣ�ѝ�6�+�-��?s5嗰��%j3,�2$��Ӏ�kqvsEζcZ.k!����2.�_��<��|]	���B�;��Ȭ`��n�aՐ������ǻ�_$wˌ�{6AAF����.k"(u�܄1������9L����M�;���]�c��>�^-̹S����VQ����K�����7��uN�L�Kʾ>lV��5;y���\�ې
UE|�)ެ���}��i�;����}I��qpe�i�xG�λ�����~)�Ƒ���G�gw/}��z��� �b �r�~�(:�'�K�m}�'Jtf���ԡ��q����8�g����
�V�̬��mL���}oz�W�<_���UA���H�6��Ϲ�N|��J��'"LZ ��" �ٓ1J 	@f �Jt���I�-[�[ЉSy`���˝[��Z��gv��pPP&
�B**e�$��eT��H%6Y����ok�(����|��P��]�B��]���nrz�Ӯ�� �j�������N��Y�]s�2�����^�IY��yU�+�W�w�,��M��3�>GK%�a`��j���
c߫��&ض�rz��[�o��j}�з=��Y�zw.�Լ�-;�7PV���u}����^������;�S������:����o�$��z+{�׫7c�L"�wgU�];J���n�dl=����@w��Vy}�Ɣ�V�_h���H��;��߼z�Y����ݎ:�mU�׆�Qfи�u4�{2����G��3k>���Nl���һc`�m)1��gen3o^G%}��oKw:�c������4�Yv�y�I1��׃]ܴ�Cq��p�����=�n2ç�Pkp*b�fk:Sd�",���/Ӽn�Yä��B���OK��$É/��IL������N���Ug��siD���}s��Ru��&���
��ڌ��Hg�����U� P�T�?��]/�M�g��WN�h�&�ON�b�Q�X��b	��@ UADS#�kt?2@}�j��oe+F���;�>���p��Dd��''ܤ���+����sXS�Z�aN��q�-��sL�S*U�B�,B�=��:�v�����N]M�r�+��S6¦>�tS���-���2/��ّ��FgT��i�=ŧ4(SP��ҹA��^mŨ[+E�H�������CwhwG��t�k�d_N��V�8�p詺��ɻ���w�����q�����u忀��V�l��Paي�l���w;ygz�b�E��5}����o��chCv��� i��_xUd��Ů�}#5����o{աݑ�O�SR��WC�Ĺ�[g�?)0W��?r�&�+Q���HR�֖�!�X�MS�/ol⬪�x<�u���O�l�����'2;�Q�PB��]�CP0����k=���μw�I������r��N#Da���o'h�V�xw�z�R9u7K�W��V���jߔ�F�v��P���e	��{�[�^�ᙝ�<�s�:yY^��ȁ);;�D�u�Ӎ�IeO"fg! 
!�+�$ک�9��c��ܬI�����>�mq���DGx�9蹠'J�P�Ć�c���ݫ{g� Q��!�9ly�����42�k1r�;+ܧ;����KG��7g�,]~��wV��x���l�fm�;,����^��|Ascbs�24�Ϋ��u5�3Ժ^+��ى�ˤs�E�Tj�Y8��;�T�^G?�"���!��ݼ�4x	x�)aݮA�n[8~Q1QA��1�μ����9o����g����J�\�^�q�������U-;ё���+o�O!5�fY;��{"�w�+U�{zDK�[�w���*e�~�k�=v��֩�5=�Z��MТ���W>�J�u=���&�(��G@��Z��)a�٥w 4wZ~��%K�e�~�N�ӣ�T�^w}L����dI��u�{�DDH�K��~q�� �BN�@GL��~g�����s�UJCd-,����Ͷ2��d�k޾^X|�T_�����I�?/��������#�o�W	�wؗ8ȂA � ��0` R�$E3�4pnYD�ɳ��R|�s���"�4d��R^�Y�Ȉ��� � �u$�4��:�	�j�<ј�.����V�fl��O[{y\�
�h^X�Ms�-gv:����BT�'�ۗ��g4^��I��|��<��5�dI�;�CK÷�}�>K��mM�������S�`�:������]��vn��W�Yl�Zq�p]'ו��ܠ�f��?JL������ݔ~o������D��k`�^���)2[�� ��HB7����>������#�fg{�sǲ���t�j�l�F���o|�� �\󕢝{���:��Vk&��k.eU���Z/K�*W>Gl�w죱 Y�Pz��ݭ3��e_�̠�=���{]�f�ƶ���	C�6Xy��K{��R/��:��R�um}.�jAwK�'�|���-K�o�<��[�S�6^�� ��J���G��������W���w�:?Y�R�RAK��>�>���H߻���&��}��ٝ�t�N(s�=���骃��[�����^
u��z�}������ؼm��w�Uo>ܻ?	 �A$�1DD|`R����3)�3C�V�����ro�#(���:fj�A�=XdD�\������7h�91�;@{�f��W. o6��ю�7"�X�B��e;�=iau9}r!YKi�Xgt.���v*���;{�Yx�����
��/=�B̳�����4��i���^��+�(�w$U
ǥG-�ŧ؂��l���<��^�}�}S"""�s���u*y許yUЌ���l`Z�'+23di�HUڕ7O�S|H!w�3NK�4�pg�}J&�A�-1��kl�,�K�w2w�Kۦ��(ռ5�C51��x.���$���|��"Αt�˖�q|����2J�����sWS��ܱ�����gn2'��`���cI8܍,���j���(u����oZ2���O�x8	�����2y�<��,<��%���Ť��g5fLu�������M���Z1��fÐL��63���z�����렉�";/��*+�Xu���Y;59��Nk����T��Ʒ��h��EGo;�<U
�I��<�����2(��D���`��0#�s�j~;[5J��#�)�{41Rv�\�mj���vb�5Q 8B��H�Mj�آ�����D֐�*o+�?r����ͱ)O���-;�8k���a�s�Hi���t��;�'�2Zm>=�ݼzgw2GY;Ϙݮ�1;�b�4��%�f���y�j=U�������w���[]�6wq!��;xz;�R��P���ګOS�
�Ѿ��߄����Ǯ����z���]L����}�<��6��D��S4�jt�C�_KO+�;�Q7ٴ�������b�
L����f󥡰��������6�w?;t�>�>'�s���s����K��Z9]��ט��o��^�Q�1��n�^s�W""33�:�� Mz���3�/�WKW9?��q�f�5�4WI�6i����j�]�!(XMf<U�3a�� /N�|
m�w�l8֚R�2"�{ٷ �4���mm��X�1���y0{i�c���Zy�6ۡ�~Ks�y�5�חfs��)��y������[OSǖm�������v�>̽�3��(�zs�A�z�s*M�8�t:'�w�Wr�J[�z�qF�t�J"R����#d=�}a�2�T6Uv�u�GɈer�:��ja
��v��������W7tv��#����u������(8���n�fx]t��*%ղkueh׶�"�
���rY�����M] ���ݛ��; @�F/wή���i̲F?)���֝Oq�&몴t�۬ڶ�z�·q�T�*�d����)��n�OW۟`7Z/�\���Ѱ�eH�ͩ�b��$���jy��Ksqs��K�޵=����YN{�|���+%�y���=�w,}:�WE�`o�Û��Wj��������<��Z<�>���۝y�遰F��t�f��v���s���c�ئcl�>�����H�;C+羻A����d�d�;5�)����LZ[���z'�ћ�����M4�,f��k�B��������cDD3 F_R�Z�����G�2��9м�;����{�8�u��F�*�Ν�.��7ۘ�ӓ"U7�<ͧ7���}�� eCȤF�;�Pt�����@ ��vh���Km��nF<F��f8 �Nm�.�k(�C)E��"��	�E>:�����g���b5��t�:)�6A�����ƻ?Cê�WiS��qw�:�`��uu�U�Uŋl$�d��
LPֆcfSa��?�� �X�U��T�{ش� �����GV�]��;���j��Q�}k��Jʻ�ӣȕ��s*�{Y�Z��3f?�Т���T�P�Q��k��3`u�\I�}h�	Z� &�'���[���巭��m��b��0�c&��쮓��
��\wjޡ��uӥ�=S{'5�.����Έۡe�ӱ(��n�Q���I,��&4u�)κ>F���t� eI߯3xw�k�r��X�'<��=�����w�p�X��.��i	��l�xh�mF�Ί����f��.��Q�ڲ2��ܫ�b&���C	­�F��ٜmn�=(�K���%6d�\$
%ѫV���r����2B(�3M�V�fC��k x�02����|��^�;bh�س-��ɓDQ�g�JD&8��2���]a���l��� K�Wt6ӱL��',��E
u�q��Uة4.�I�P�H�of2n��)��wj�_twQ�Ҳ�P�f�"/�����etS�}$��$��0)�a�\�3Qq�����qj��Q��w0u�����U���Y`J0�u,�r{&򡠳��v�-�nf<}a��G��p3y!������9Ցܺ22?hd�K�Ya�_(��.ˮo���,`�u�IV�Nq1�b��bƆ�#���-�=�KR���Ozr��zo�ͱ� í�TVd�ٜ0�.��=�VmZ;?Jٓr��)ۥR������V03�k�"B��	���P�D�8�[�L�A�\����9{Uy�iɴ	*��i�+Nv=��\;πk�+�d� � e�*KQ_ABm!���w�6�����绤�Vsy�#F�X'��Z����7m���^��n+�ױ�9c6V������H�H>y��H�C�Ʌ�R��_[C��������ݚ���`q��4�VjvQ��17�n��玈<u�J_md�ݛ�0sƖd;k!lV�r&�ڮ����4�
���9��Β��3���g4���f`Jm�����j�/�W'k:��p�?f���Vo~�WL�		�����7b]�x~���{�ػv�'n� ֊'�����S8��:�)n� 0�/*f3Qј2N��"��hZ����7|9w*4m�����+z\�߽�A����3}!ӬR�^r%[ު�s�k����K�I�)���CC�/��عn2�����	�)K�U$%�7������Af��JA��a��7͜�9���Uq۬W��*�uu�/k@�� #۲����I՚��f���29g>�������a�k��\�L�u{��1���L�k;ӣ�ˆm+WčWҺr_�E�r��6!��?
��)�I���L�d	���1F�ۣ"�8��v�f�_�з���*���WlYbW6:!�,�{rs.c#y�ۓ}�ڍ�5��j�����$k����@���H�߫����urV_9��ï^��lf;���ɪw�T�g�\9#U�'�t�����ݫ����Ԧ��}7Ec�L'6{M?�=� zΣ�d̺�W:��/b3o������;/WE��b��������A������,t�1�S�?L YO��h��9�I�}����
��$�5OEE����|���N�K�D�	����>5�����������.��ٟ�ޙ�m�5�8�f�o�t��pg|=a���op���x(U
 ~$�J�X����ז�E�vټ<�.�WJ�(ힽ�9]"�b	 �N���W˧dms���'7�pZ����$A��_e�R޽HfL])��.�5��f�eE�ۡ��t��=-B�����p�E��l�{������H��
��]Qh,۹�C.�+j�q�Q>@�w~��52�_��Нݲ�8��lS:^�K�,W	��7�=�}�wZ"���ٹ��I�KY���ڌ��n':��0=)�Q�.?��n�5m}K �僆z׶v{�H��E{Ne1��b������!��6����*�����e����Z�vv�Tz�y����oK���;����П�&Q�Ɍ� c��/і�Pb��o�}J����jZ�v�u��2�� =���v/��{=ꦗucYR���{9]ye��j�[|��4��C��,Ou�k�yJ�V㧒���U,&v����k	<�f��t�&��f 7'6]��f2���~��p�+���NЮ�֞�\����{V�M�O+��0������w�\��( B
�D�"`"`��3R��&F���a9)���b�N�Ck@��0F�a@cA�d��40	r
8�!�nw��L��opl�s�5��`���Q�o�zm�ԥ�
7�F�T�k��p�{)~96�X�:���nl�z$�n��}tk��J�����w�Q�(�з�� �w�I���UQu^d��J��3_���X<��]��A��}��9��aA������u틎p�Kk��%���;����J���ٛS[q��������9[f����7_��G��&h�3t�1��3��7���*����xvC踌Iƞ�Z�.I68��Y�ٛ>K���d�m>Ϣ�z�>�=���+���Pܐ�Ҭ����!X�[A��l;��1y[���y���=]��.~l�Ȏ�~y�l۝����^��+(�]��vi���ٽmX��<Vf�FA{.B�~�kr���gH�󋊫[�L��޵�&.���[�� ���7���0�j�)��x��~oC�?�{z����A�6r�������q�����&��ٿw�;#"EF�� ����؂�.�s7X��ۑZ��w�� sI;�΍2`���f�H ��(P��B�����҆����jh���*��ӛ��u6I��g���W܈�1�:E���ޭ��+��=��k�����4Up��`�'UΤ2����aP��\�������fsMz��W�b� �0(��L�|�"E�f�M��Xn��s1Ytfyq��*�"z�������@u*�o>�oTcgdU5����գ���]�qD=/)�1v4�����tr�D����Ո7z,��귔�R����kY����U��=���"7��r\��~Ӧ���=�ۑ����C���J�nr�X�fr����폫�=i��)�s��ƾ�;U���$xq`i&�_���:׾sj����IUv��vGd��b��L���.��Z��=�CC�bעM�9���-����{��	s1)���S`��;n�c]�T�ޗ�3J*I'j�����D}�[���|3���O���]w��s�
�|܍z��ߤ�@�VYއ��þ�+.��n�N����:T�������ݚ�T�ά��T�Hc���pÒ�0)�N媕�ܨn�)r>J�h>p�=���042ܭ�vBm��'����b��B-�b:^Aφ�.�d �p9o�˾���im,��S�5�޷�̄�	3��\j�#��3�[��\t�k��7qe3{��Vv5z6�4��d�ާNl�_��(m��H$�5�Yo}���زr��1�\�c���oUQ��}Ӗ��wj3��}�|��ыC=7���Z�P���9���h�
�f�_nxm@�w��B3C�Ba+�4op�!�(۫C���W=�3e�oА�`kپ�>�mZu����!�^~=��g�z��ND�J���sE-4��p3���&��=��d�F �S`#^�;���߸U����M�ǃ`���Y�6�ܧ��n��Ž�p��	�c��C[s�PxݽѦ+%g_w�⟎�gU,���h��Jo����;�Lv��<��̣wV��F�u�i�����n��gtl�J�N٨�jv�8&		�� �Ii�$A�L0U����<hJ�{�S<�c�^ʛ ���sϒ�r�W6o`0E�1��N� �$�I	����P)b#�

@X�k� -ul�u��x:��M��g�8Vn[T�.�z`����Z�ά���5wF��RY'�7g-vv��W:c9>���홫��K���{��ߢ��Qu3��C�I]0�����?`WS-�E�4��=��	xzN��-�k¿W��)�ڗO;dK�MR��],ԊҊ�H;��>�b0��T���F�0�Sp�[o�(`�����S��Qj��W�uD3�f]W��qn�*;�,W��I@e��^�x�.M;fm����zslq]���|��9����C�ѹ}�<ij�d��o�3z�����ξ����TV�N|���t���N%=�n'*U6��yx��h�3ۙ�)�����䅗��c�r�y���j�����iK"�r~w��_+C�#�_~\��P9f{=������9)%�f`�V�Z�}�}�9���e9l��,���S��g{*�����88?��z'U��;	��8��j|z�/�>舳vMb���|�5�ٺ��N��^v�S�f"L 0�ƚX�d�/3#7�j��T��:nٹ���|m�b�u�7{XS;�'�0]�Nؔ�$��:�_vZ���FSF�M���:�\�i�(bϋ����k�;�X��Y<]���U�6�ם�M{JYߟ]����lw��f��OwUA���c��$�<��45TM�4+K�ݭ	� ���_pS�zLp�7[_n��gN`"��@��zF�����7��Cz��4|N���1t��E)Y����;��>hl�uQ���Uk���q��2�vn,o;����d2n����[!Z�O'6�ɇGI��׼�w����0����HJ!Mu�-�y��q�pNCyFV���X\>�����|�t)d;���M.�>\]�Q�?��iF}&�qD��x��H����k�i��X�>bz�&����&�v�͌���� _��7�A��I)�̪�\Y��9;i�[�L���S�D��E>"}�{c��{��ٽ�j*��M�j�\�R��Fh"��(�E�Y��@ �t�?��[�J׊�פOt�w�l��P�4&KSKd���k*�~"�!���`"G�m� $
�!��$C�L���mH4=�][u(����u�1�ӗ+
I�����B�"\��u�u�oe25�f
蔫*�f�o,�5�w�vPC�V׽������=�]��m8㏲&J�ަ�x_kEz���jY����Tx����������
�lǬ�B[�w�=�Fԗ[��0�f�����ҏ*ꝃ�d|_)�/��:�>���F�8��u���f��Dt��|̷ *���_f@���n=QN-���(c�j�>I��L>�n�u���y�׺�5���<�;d*�ɵeg���v����U��$w:���Yܬ߰9�s�[~�d��L5z/i�}&F�lJ��*�3m{����AJ֓��2�Й�=L�� ��@�������}'�^8f���|�)���;�X"�?b�>��uT���qtn(�c*��Jp�����wROe⢇�ח�z����P���m-��Xע�te
�B�t�y���赲O�~���+@
P�Ҹ���Ld��u��=�����}lQ����'��i���f 1l(�424&�l�y�F]������ޙE��plÑX����n�:�F�o� b�T������Gy�5	.��\������4֘��Uǰ߾'��l��a��Ԣ��T���󡅹�4�r+nDvq��=�;�`y����/��YUz���1�;�K	G���ٝ}M��ж��	拷r�n�y;39cin�PY�OK����+^��~�~�;�u�k�l�)�.}z�s�屠�4v;7����fWO��Փ���Ȋ��ų�Vy�Q�Q#�W�w|������>�W�B��g��
ʧU���Pֹ�C��w)�>|}Kz��M�{��P�Й�+M�E(��C!�EH�5OV�3�	၈	~4k����9�^�'e���" 3�e(T��k�3��	��.�?����j��~�j�m���5H��v�`�o���AN��� <���	�}��ۅ�#/���k�g��M�їL�;�k>�-��r�W�\H��mEv-
"��hV���NKb�:�pb �P���� �%�^-��+Wpn�x�D�Kw2��7(5K����_�wtkx_�����}o�
,�4>�;�#��{�R�Ôdgv��O����j�/����^�_���)M�γ������{�Ͻ�� 3S�g��<��ft��R��u��r�;��3����x�͌���]�޻=T���,�UW`�ꯘ��H48T�� @ ��v���o[�����t��Y��� ގs�;7��^Y�<�]z/ӷ��][,%����B-���ݎq+��
�S2���7z���z���f����H�$�]��y���YrL����O_Z<�fw6�Q��U�uU7�͜�0�7���D��ʌo�I�X�ҝ�����o^�����������b�[ow���u&*o�����p�^���k�w��2!�ڳ�^��If����X�K�쥯<b�~9g{ζ}�����D��YG��sSqw�kꁌ�.=7�N�/�6��~Z��/�{��T�ɰ�I�1�kJj�;4qe2�qqQ��LEkD2vhرf��;��8r��8XZ89��Q�B��(
��飯	3�_N�᜵ &f��e�NJ䯨��ǔ�w�ޭ�F�6��Kr^d�M��܄�8;XՅ�p�=Wd1"(U��*���xQ�I0@D E��.gq��P- �� ��L�P,b��* ZM�jD�_mZ���v�NR���1�9�vv�X��b��1,��q�ܣ��êH�5w�FZ��r]7G4?���m��V����lY����T*fȯ0o��&Qj0nذ��2T8��M�����(����K�L���1��m<{r��i'l����ysxF�,uyy����Iq�����e+�Ty�o��:�uuėڕfNJ�eoP�Ւ�kI��ؒ#[���EE1�-gS]p�@VٽV/jx�5�խ{�3�T������!"%�.�U��tM# �5M�b�B����t*
�LHV�F$��y� ��RRa��	2V:�4*	;׸����Y�4^��U�{�es��l�TvFN�h�6�v/�]�f��.��!(�!]e��L$�P$I�2�H�%�ջ��vs�J��t����fK�2���$BcZg
s��v��V�����\��ы�2�6T
N]Sv����5[�֨aM6��%~�+t�c�}M�Ϥ}#m�ܒ�3��h�:Bj��-(Byu��a��k�}�νf�:ӝˮ_Z�8���P��x��>l�>o�f8ӲVk��$5-�ݳ�͉pb�_m�� ��LO&.A�>�guo��˛��!o(�/5�f-�����@�c�;g*��q���3�Ղl��E;��w]��b$�u�z��i��)����A�g#�XS�^Z�$��ky]�;�wu��+Ujc.�N�_��[oGc��wv� ���nH�;����]��M�lT���H�G*��X��PT<���*|/���k�V2S�x�w�I��&�Ӭ��"3D^8"c�`h�)�J�](���'9;hc[o?-�G��۫��fЭ��կ�Ob���|��,V�]E�)o��y��,�OWBJ�Wf�S�*��9��q U��e\��Y�wv�#��S��fGYB,@aCQ�̛���r��iK��yF�\UYb���e�
�,c���������3���4nb���[�N�X�$iAt7}�7;�7x0T����;SK9m$p^��w�]�����)�B��)Nѯ�Ӷ�h]�r�>��ނ:�-e��[7���]���e��V���^�����H)�*�<:������v
^�p".�=/E������q@�wT��yd�+�"$^X}9T�[���2U�`Ĳ��O���Ӊ*s�9�goVg�R�x%�Y͇Ӫ_'�#��Vzèpp �	�պ�rV��Y5�ϣ���\k ���E�=��P��9���}�)h��s5�i���_�;J;�_:2�Y_u�l�ƨ�E_�r���,��	�vwo��s�jd=)����Ԟֳ�6t�C��ܳ&u�6}_`�zu��\����g!�V5�Z��]��Gn�0��������׷!Ґ�@�Dz[��}V߼�0��N���Y�P�5���m�o_Yg���-�ai�u�Z�
a�S5|#��(� '���	�.s�[��{y9��D���� � O|�麏O��`����<�4�㹶c؊�[ս��m�F�8�4QJ'6���V5D�<�/Rn���͋�UtM/��^�b���.���N�id#G#y-MzuqR�Q�ݜ����q���Ty��_<W���*3�J3��U�v��]�Q��@�Ms�*9��]\��[]�'є���-��)ع]�VH& �0�,rh�]�j�9Fwo�n�m��a�wR72�
�m1�"�Z����:��E�Z�Z���{�eJ��	��]���C��
�R��J��yF�俏��e�d<�A�L�_������Ky
���}��K;;������3����S���gh��l����������4�yY=���|��������a�k��>��@�<M��B�\�V_�{���Ot�ؕ��w�N��7�X�lU��M���,�Չ;_@�󸛅�oN\��Y�:r�o6=�ǳ��|xww�/��0U�aV)�]�rl�w�=c}Ji���6����^���q	��cU��GJ���7)9	��A��LT������Ap�O�Q�����{��@��\����>�>�f���Y�S�����g��v�ꆩ���d�	�6j��N:���s�ƛ��΂��c3�6;y�Q��e�S�MS"��jȝF�w����A�7������\��e!RE���?��x�:�}�?ns�B|�%ʞ᡾�M@�b�\�r7s`�����i/�gv3�p�B!�@p	'҃�T'��ӷ�R�F���]���t/6k��G��KX	�bp&- �PyE��$��C+p�qz�q]��lR�r�dLX곚sH�p�f�[y
���u�f��d5eB���k��ku�Vs�����_n�;0|m8���w�
�Y�m����9�t{��S3��W�{
�)sGި�6辆k}S�vI��I�,�[�m8�pn�ts��c}=��;"jRh�HF�S��kѧw08��y���@
��� @>�̙1�@�ۚ�vӈ�zqe/XoZ����uB�?-�W0)p�չS�� �#n�4s<2��;��}��'U5����N���.�AS�OmJ���n�,'�er�^�?�j;�p�÷�5[H֎��v�FVl�w/_0�N�So±�M&�o5���~�̆�Cdf?1Џb�>J�g�}�֘����]$�
�6�lc1N��Ӕw��u���T�?Y�����y�ܧ%�珏N8b��kڧ��j�&�z�gGI�L�
�u���γ	���W�|�5�vm����n7`�kvi��Q��x�(����GU,QT����YB>��0�u�Q��^�~�T��ϰ<D]㼬HӉo,57�X����5�V������q-�Ӷ��cE��v[���c���α2���%�8gB�ŽP�/6�Ty� =K���|��N���Z�O��}�������y�/'>��9BW�4��SɅqփo�z�����ɚM���<��;��(
їqHǄ�Fk���~�ZF܈G2=���{N������or�=������Q��V�1X!(wl����}���w�$�
 U�U�Mv��t��)�?S;$�)�+�j�e^���=#j}�g3�R��^�|�z�:�.A���<�317҈Ͱ�DJ�k5핽6Kr/;��ifV;
}��=�S�Nzu�(�ۃNA,���<�#-��-�u��)��EV5�^l�#2�&�P\�����v�]ll���[��y�D�n�e�?/on�/3����㫯y��W��ʘ�Y��D��T�B&��4��_c�Å��ֈ����Ϗ\�A��S���7
���]��:����S�fl��`���ݸn�&��6����#�D��E�"��T3��%e_r�.�*T���������E��+����_vhO�Oh� È�c���{��$�S#I��/D�p�q���3l?���k���uT]]m��ɖ����q��� N��{�U�F.����*�n�2��;��_�������� >LO�����՛v�*L]���f�N��m_��ö���#���Y�6�v��_MQ��<���[[խ=�����~^���|�������+;b�^�����t���S@�+Ud�U�
�9��̗��e/�y�H�{��i��
�۬�]:2�E��=^ʧ�8�q�go{�����&E���{�ײ�H�w�O��S�U�f��k�Rϴ<���i)e�!I�wK��c���>(�R�z-�L�V���0��G�`>��i�}/���d������~������;�N��>�ӹ�_S�E\�o�Z���A=��{�]Z� q�7,|{�1���hD�F I�/�����N�z�d|V���4ܺM��H��=�U�G�@$2���0(�!T��\��;H��f�0��ZUѻQĴ.-nr�R �^=5ļV��O�@E݉Ý2��_r�Ü�W˅k�F6P�<���s�פ�sW�g����|�{�[�0��E��������Zw:�'��D;WVcM��Y�m�i���'h�^��"ޮ��5r�����9����'�aod�v�qOd2)��W�l�Q��ާ�����mx����b�1 3@�mY��B�q��V>{�X�	"2��F�L�U�S�ƪ�m���K\.�>����z��M{��}�ׂ�������5VR�YϤu���CM^^��'�粄V�n|Ǻbcv�>뙦v폝J�=���s�����O/�M�P�W��@�_w熳B˩����W0�p���ft��u{*�w�E|��hi���m�7�t�o6?�޹dN��K��ܱ�)E�e'�y-�:�o�Srƶ����~�h��ۗ��.��)�1��c !�t/��z���۶��S�B�\��*��j2^��c��i�DY`о�x��ù9���P��˒Q����3�
�Z�Λ���9%����z�evM���,-]%j&�e�����Y�~�����cp��f滭!V)WzgS��('57^NGƟ:�+e�T�:�5���glD����Z����p
���H˚�����T���3����[�ؿg�Z��tki%�p�ݥ������n��d��s�-[�>�s���3��&""�uY�99z��K[�{�������</j]fZr�S��lYd����۾��������S}'[=���q�r��������?nW0_��'�����C�M0v��t��},;�|�U)���v;|��O`�΢��W\�����׳�9�m{���L���/9^v������&&˞�MJ\'[����k����;�:�5P)����u�5�b��V���}՛�����؋ȭL �	� �"`�%$	%vW�l�)�o�'}�:�L-y���AC�����mUUH� ��H(� �`� 2 �b@�4�{�%Ov��Y<��3'|���䍞8-h���e3�P>gMXo�pMP^n��g W,.ufCЅ��I#s;J�ٸ�-�s��u��.�ѩ����c�U5�S{Y�?���Tw�K�-�Ē��D�6�=��=?�y�>%kV��l������ˬ�<��/�M��q0��2���<",�����.�����|��ҏ}OS��~�bz���Kj��(�a�7�ҀT��Wk1CYY=!�>�Q�-�)�J"�Ouc3	<��loD�4�q�\ǘ���{1�ۖNo��r�B}�REΙ�+�F�����w���Rz)�02����$[�u�u�i:|���uؾ}�߯U�|���V`� 
1��D�\�����x��&@*6-�wO�O��XY�����7�윚�Z%�KN|E��B�C`�2ms�6�X�����6aE��$�wW/9�3O�X2��h��5�r��=1��o�<����q���y�罢��cx�����`�+�ܭ�Wf�*hù��Dk���T;�������[�� x 6>B�D 	Uw�e���X~X��j=�1m=�Y��N�`�#� 	<b��M�:12�lj�KNe635`��K;��e_<yh�G{*�(6�S�B���V/����_M��in����\������XҽǝJ�����mj�����+7L�����u�B�e^���N0`�����ߦ]��%�,��bq��8�����K��lyX�]ȿ�}�o���\h���g�pH��R�Xw�h�!W�=b��2��kͫb��dp�q�:�]��G!��m΍�V�0��ދ}��?�I��
ޮؚ�~,�Ϫ˸+ɸ�fJ���}b�砿�uG3ch���a��$b�4f��=�깫+�^�
G�Q����|���\�Y&n�.3���6�&���=�u��g�r�L/0��c�ϻ�o��'?��\6�_�*ue�W�=��ʫa5�k��~�zʢsL�%�L����fq�]q��ȼK۪���;9Ԭ"w*���kt�]z�9�u�R�>��\?v��6*h��q����n��aw��f�aϱ���m�3��3i����oyu��37��z�8���9��R��0j�\`�	�H�|�Ma�z�,�a�ICA�� �:v����)m��Ӊ��L}�E_�R���}Ju;�S�L;�l�0LuP<�HY�Z�	8��qT���CU���]����a���vB�/�9�gc���`���c��?��S�:�(}��C2�*1����K�8� ���N�[wC�8HO�wۿ�����{�靯c��=��b�F��3+�[�uL�S��j!��w�H���#2)�>��X��i��[�z��G�/w�yn��e�eRQN"��T]���s�Ju���J�iR�`��Aחh 2V�{w���"홙�vĖ��Q9��m��e��`�|�����Os���S>^=�2���(��rk����琩>�'������m�>�~��Y�^��v�KbVOt�x O->h�ދ�I�}�2;}�l������?K��,�QKp/��}�d8�������wv�����5B^�%O��o�bI���T�f����اy�Y��ܑE�n2�X�p\n\�١FW�0�lHS����2�ma����iz�q��'��;��1���ywà��1�g�nR��%@��yu�^��O���c1���]�yܹ}L�Ͳ����	��E��W�ox��D�sM����ݒk�q.��wl��k�%M��,`�(�V�CMī<���{%���@�Fʭ�H��V.C$���}t�+H=Ի���C:U�;X;"��Uy:�R��l���\�W8�m+�J�H&"�Z(S�w\�U�ݗ,hNg��;"YSVL��@'V��$�q,�M�)�	L�Tԓs�P̜5h�#f��Xj�E��	|�e(S�0�kFPX%�LZd8�̨RE!Gi�y��@�, �E�E]n֊��R�dU ޫ#���%��ִJŌhoKބq{�6vN�}:��er�/3��D+4�u;{Z���Kn=�yXA �w
Vֵ�NP��ɩL�tݼ�{��ܩWJ��*����Q�&�1�'9�\�������	b�^�.z�n�3����ڲ���M�Lfp�'�o{�6�:�7��E�U��-�j�:}��5]WoIR�f-q�p�:He�E��W`�tŃeSE��QXn�l[�z�iԧ���i�U�u!���8;)��`vv�ں���͢g����Mo,�D5�Rh�*�UA�Q�aW�4��z�y$�aR�4�����j�K{��0L�"r��+	�Q���8�
3m�����pBiv(�5eUQ����Y��'�^�%Z6m�5k3�d��ȫ�7H�J
	y��LU�.��5J��uw8P
�@c��t�:�q�A�&��ټ�d�\�\ʰn�MIL�Т-��S/gY�N�M�����ɐ�Ou�U�\a-���}#m��wt��n�0��)�tb��h�'+Bc��MV�ɵ���=y|y��+�=;��I��h���qa0��*9#f�k����w���٩����#�	�e�ПjK�N_Wq8�EdS@K�S�]l;3���A<�vh�X%�5׳���k۳n1�n��6�Q�mz3�f��\u�l�{ԵKP�]�wn+��J�0-���X���E&��,Vc�X!Eiz��<
�^�h9��s��9��1j42Bȥ�cQ˱�X�ѕ���
�K�t�.*�-�ک*�;Zl>���[2��7�r����{o+E��z1/Zђl5�C��-`��s�_�ˌ�#p�����XS�|��a#�s�պٯ[�[�ݸ�=5�x"���Yj�D�=�aΗ��}�Xyt�޵��Nlg��y��@�蘠�_1o1oٔ$��_Q"�.Z�	��!�É��U����[�V�M���κwv
4h[���-�vS�k2�#*%K�Y�˶��K�sb�w^f�݂Q�!��f���#�WbhW.�@���7 1�י����y��f&H�tC�Vqnn�;�Wӷ��	y7��A�5�8��Y0�ŏ�8�o[3F�\���V����LWdv�Ҫ��K���Q62�s&:S:�ewSޫ��s:M�Zcv��972Ԭb�:���|�~���eJ̥��D�E�(�m;(������f�z�an"�v�p�/��.U�Tԋ�p(���D�#!��NT]�x�vз��r��Dꇦ۳��I�\��D�6�V�P��.eI��̓:�b#������j����p�|�����y�q�^�J� �{hdT�S=���)6ϙ��v���+k���P�g����l|<��L�L��k��|�������`��/Ht"q�����ĢFҖ�-�]"�xV�^ݡ� �>���tb�ބC���D��|��!�!����P�[����85�/�}B	*YW�Y����\�_!ݪ{w.���zn���ܳ�"��e��%a1��G�)�Gov ג���Y.R��QR�_'�t���,����%Cʆ�p�����Keo�M׻�L�����#�zp�4���A_EDD3��U1��3]RN	<�<md�8;<@i`b�a��64	j0�\�yv��̗��^���;;~럑4�'�N�<��fN޷Y��G�������с��ه��oF>0�L���
`� �><V�8xq����֕��,X6}�`��@��a1��
��[&��n����T�-�hwN%�Al&D"�0aHd NH H&" �0Io��J�Ŗ��x��ܽ͜5��}�t�띒���b�J �"	!�r� ��!Lb� ��tCP  �wf�u��J�Y��B�z\����[�A�KS�w@��a����ڕp��u���+ڋ����֭*Z �Y�a_G3���{�:\�{����잞6��*�C�%Vq�T���v�p�s�4_)>���
Ɠ^^d���X}�sݝ��R���^����\z5RA��� �?��Ԥ��������pu�̉��뻫ȡɣA�f0�1�{y��:��\7fB|��"��/j�N\X�4���9o]�U�k`҄�cM���[3���[o��F��i[3�vmYʏ^�v����5�S�(��T ��H^�0:td�V�v��ق^؞���؀x�9��L�&�s�fFp��#�%����2��1��,5�3�B/��W3���L��'ٞy�}~+�'�=C�WҼ9%b�(�������_�8e�}����gmZ}�?398U~�Uᅱ���"YC��X�J�t\)�:��{ ��B6m�+Y�e��צ9�y�ޫqӋ��j�]���K�u���UlW��A�O���cnnӃM�uz
+�֞�ٹ"�z�'*�(��1�����m��k��u�����@6�q���=K2r�7]�vu�� �h���Jj�HQ�5�2�G�L�[B�(/_
�}�p��27��p�6���Ǟ���{}��a�x]����Q�gA}��nƊ�VLG�����<�� ��_s+Jw�	�Y5Ob��t
���~�R��${	�7_t�o]Y#������*g���wz��	��񾸐w���垵S�:ד`iN?�L�c'rGt�*�H���n`�
�A�%&�p�������&��@l{�G��qM�}*�}��6/H&�T�c�J'�א�4§F���NU����!�^B�9�k����?hf��?����M1M����^,��ٞo`O9�ɉ�Ѯ^��O�ߛ�$����=������+p���6��e�<˱�;p�a�{W1�z�p���Г�Vs�(Q���MT��o�>a����o8&W�O�1�:��;KJF鎾��X&�W�%� /|����3���`_���>
�􁿚��6mW�,ܗG]Wi�Q���  �x�|ꯏV�E�����5�b�E�a���	�Tq�^���w�ێ���^k���Bv4ݲ�J��S��q���ٛ�<� &������W�_����2D� � ~۰f��.�i�3�Zf��'����f��W"�0+� Z.��՝m�{@��{��*޿K�f�/Q
��0-�OO5ë�>�N���_9�(�o����`�M:�F�-w�b7:w7��>�i&x�f��'ES��t~����rɆQ?��������@-C6������; �C/�����L4-S��ڴ�5��q"��a��l�������S�ӝ�<#��"���ÆnU zb޷$֡��O\(����t�O���%^��l��2���l�P,d����N�R�BPV^V��`f8�q+'����>��_��!h��I~���D�因������#�  9foa8nٽ�H�̍9SE��bt�N/!C��|h�m��q�Q���J}�˴7l�[�����Qc¶�ut�#'�9v���&�1O�+[�/��b�hԼ�8>��G�Cʳݥ�GFV(ܗ�;:~���xd�i��ϝ���g2�g����������<�]�g��p)��I"�e��'O}�s�-�j�im]���}g���K�������msR�>�x/�c C���o{���
_�I7/C�N���J1|���=d��`���Fg��駝?,�wiI�Օ�V���7x�ri̼�̱DB " iʃB�`�v��W*�%��#	� h�؈�7r�cL�J��zo@sAsq�t�U��gX���XJ����:d���8k�z�1g�����xVq�/�ə���_Wd\ڝ��Ph'�T�Ū;�nîf0��9����_),�*6xu.��f�X���S�y��i���8{WA�L�ߝ���p͞���w*7�X1����H�`{5z΀���=5�gK�E��h=�TA�#*^�=�״c�1c��{�Ξ�ƯZ���/^�)�j���w��,�����}�嚞Ce�B[��N����O��W���8�jIL�)w��N�ب��[����!OP �]���1@����������"߂��N�����vܞ��vm�ph"d����1*V��'�V��
�'~jQ���N�yM�\��
~�?��;�gE�Od��Ow)��j�R��.��@�d��s��gS��*�e(��u�;2�¸m��n��u-L����o��� x\�l�;�U�Ƴ�.�nU6�>#��ݼ*8�XNj��ћɈ���<��GG���ay�s��j��.Rݭ�b�J��鿨-B�f�q�Z
��D�X�G7��&\m��O6{6��TG��\��zT�@�7�/g`�uʹ�h��nv����+�����"wSc�;�j�Z�.y�Tp��5��V(1�qQ�&;�����eo#i�(ԹtO��c��#:t��(	��w�Ҩ�p���y��-�3�6���v�t�;�����5����B�~��K�lbX�3b}��n�I~a�8>`&!��L4�9�b ҎaO�kQ�gw�Uy�>��@���ǘsо+��S�5͜�a}^�.MԺDH{ ��E�}�.����.�y�_��wR��{�pD���z�5��C+��c��<��;>Kq��НГ7�Z���LqM'���Y��� �΃v���X7�b�қ�����׎X޺ܯ���(K��ñ���DA�]�Z�q7�O?}�^�T�r�=C�g�.]t�eJf�p����Ϳ��ޗn����,u��#8L{�����3ƺ�Ҳ���ѾC�E~Ҿ���_�/8�]B����$��Y%v��.Q�|�˩�u6��j�<׶o#Ǔ����@�^u�"��Pd�����*ŻZD�;#2I�~��+.����$#]"&YbL�M'@&!%�<��6��y(����00֔���x�iZ����H5m�1��D�q a!4��l��D�*	��U���E�Dތ/<����l-���S�YWRZ,t��ijv.�缹�o	��;�WP�neut�oP[��r�_n�-gK�YY����z�ky������/�V�U:1�6c���u��v��m����Qz,���1��sE���U&=J�׺��0��u/v��M������ީ�:�:K�.���w�GFO��Kw*6|�(��矯�l@(w ��Ջ��Κ���,��'�z6�X�GR���X0'�z�'#Wd�;:'Ô琛�NW�F�w�ͮEeX�� �W����fJ+�t5ihcg}��z���]���l۳1��RwYՕ�K~�R;ȥ�v�"�c@j�Zo82i�1�'(�75[!+�$L��9�o���eۤݔwL��A.�c^�5�24��'����ؼC>����qq���`V�w��}`v����E�SD�o��Z-����鍕�����Ti��<S~�����wLd�l:�o6F���W6�x����b���{�ѝuΜ����q�X�D���Z��vgǒR�Ng�-C<�������|�T{�$���b",�D;~�aB�M�ew�}LÊ�o�T�����t�Y�1``�A�L��N:uP������U�Y��hb�Ekk�9� �=Ǣ�:���K�;����%�����]��������I`.��w��(��'wgK�;��}2�#��� ՊO����v3uTw���K�tve�/a����Uٹ�\}Mi�~8�������n�,��ES��˜{���_�b]K���=4S�vg��y�&�T�������6��5*��R�ƹ�=��Q�~���7,���˭��g��Is��k�fZ0�WuޱUS�;�*A��G�閤DԦ��w�����GS��:%���h���w��(�_��jHgyz�ِe}��S�.�}�h,���B�jv�o�\�B0R*s�I�MȰa=뎂����]��Ō���3����50N�3;�֩ ��5c�ʀ폚�ߔî5'B���5���I93r��g���*��7��V6!\s����v��i�yK>�$�/�!�7��<�v�"��J�q?y!�s��enYy�7�4U��'��Xc���(�$�]�Б阬\�TXs?t�=��zz�{���j;�y��� W
�e���.����[j��lS�n�3WH�+�j>��q��+.�
���I끸i�n�8C(� Py��� �����9�����2����/mc�8HFu�t���_]�ˤݠ���t�[<���8Q�i2O.�:����ՙ�J�=�i�0?�ͤ�й�v�zzVT�9�R_-(8����,3370�8����۵���j�����M���#�^g|k�{����v|���'<^�����s�I½VN���9�+�`��	�d�k�d�g��A:�K4��g�ۓ��ܜ4��}�e�v���D������/�.f=v1\�)Xw�t�ࡡ�n>��q��ofG_�`�OG�م�G�������'�=2`���y�uۜ���5������[۱8߬f\�{$"���<��,	�Lʿ�f�XI_�����7��[��!���䆍�*掩�ep#����}Rij��~�S@5�w��޿#�}P<$�y�7;�aYɦ�=U@:ѓs%��yg}����r2����F�m�Sv'��U;��H� �dݮK)O˷�w��<�
ؙ�r�e2�ڮ�*�����Ve�=�����%�>�\TO�P�f����q�ud������C��9PƤ� 0����3J�`� "̶�
�{e���&�Tˊܜۮ�6s�!]ȼs��`q�0`�@@��K!C�jS�s,�d��3e4�>�x�S|�v���f{d#���]��ޒ)6p�٢F�\V���r\��Dm]�u���[�B?Ӻ�0���r��}gy&=�|vǂ��v��\G+j�0��-x�_\<W�����k�ꭻ�͍ͰkO)ڬM2ע���	��u�b�c��9�&,� �w���,��d�u�g3�l1�~77L�;TS>x���yC*�*��!V���7�)e6����D��݋=�vX����]�KC(�i���[�C����4X��H���9)�*�wx_G��>W���`�"Y���>W��	�����w���Y*�������s��6��l�ȷ�2���;v��^C�t�s�"M�(WUJ�]a1�4�oޭ��K4u��z��z�r���#��kx�z�����v�`�|Y�{�jZ���Ӱ�'=���Us���6�N֡Ф�t����xK��5b�ķ^�Ǩ/�Ͳc&Ce�6T��Q��M��1V�A���P5�'����J��D"]ׯs�ܥ�����u�w������M���Gi��U�8	9 (�zk>?j]��^ �7ͧkg>�kK�s(^�w1�|(-u�N�J��*�gUӭ5�$葅	H�*��N�U#T�(�u�0H��J�l���n�i�X�:p�ͫA�9���l:AqAK��Ԭ���cY�Z`~���uEOѩ��t8 �x�K2I�LZV\�B12�i�b��d䊋)(�C���
$�f�AHHSU}����Ԛ�P�\��eVc[���|���5f<_inC]u�%i�ݗ�S`Hs�}����z�n^�����d�B���ՠ�5�M�5]pVy꫱G.4�B��̻��)NH�G0A��%�IPu`o�9~oX`����.���<Z�'4:��^���5h����8,�ӈ���$l�і�!�pv\�����;8uZ�әN�u�ia|R���?���qm�7�\�;�ΧMd�����*�JU���_#��.ZWU�Kz�s���T�MN�S�I�qPr�S�Y#����W���h�*������F毸o>�*q�Yc�1��1M܄D�R2������R�hS(�($Ҷ�(�\�F�+����x��w��KC��ɪ�e�g6^�9�bL8DQ&g/v�5���V��s���b�d�0��V�dM  ��٣P�Y,T)��t$�֍���X	%X�\�M)V�݌����zh�M�����eT��L�##Is���t��*�����P��+`e�{r����t�l������ΒI:G�6��WY����\']�,5�3�2��8IŪJ�<<�u�O$o:FE�Zv������/���F��8�-V4WK���J�ط����v�����CIw 2�gV0V ,���[��)�Ծ���7���r:nغ�Z���~���v�@�8�"��f.J�kzzN���-Ty�����[Ӏ� �в���Δb	b����iW	�7F�vV>*�~�[La�Y{l��5�z4r�����	W,!a�|	�Y[��"v��xz��{}�cKd�]�s(�p�<�qew*�,C ��� �(�+n��T'
����f��r_ײ�Q�}��Y&�D�a���l���Ԧ���\{�]5��]��F�<h��g�GK��`%�\,:�r�ָ���=|R�7������j�H�^V�j��zX�t��\W%�fD��X�Iè�<)݀��K��8#�WD�7����L�V.� cd�]��WI:-���O��]�d ��R��fwO��8R����cRh_{�W3�j/�).
빁d���x��K�{��ӆۧc�.�l�?`z�b{t5%�^�5D�<L��	�!��ԋF*Q��e�/aM���.}�潫ڜ��,�Nk�܉ki�� ������n�`�ԕ�bU��n
m�;"�lc�V�Weds�v��s4�s�|���hK�O/;��T:{u�"�wM�G��+c��t���Y!]��ZS����I[��CWu��Z�l<�ku����]#a9������w�d3;��vჹ��0�ӳ�gb�T�y�Y��&���Ҡ��xkӄ��*�� i�{�͔[�l�%U�4BT�K"Z�(W�@���W�*��c���vl9������C��`�6���3����{>D�=]�q\���{^{��k��i�
U|����|���?	�&�E�ܘa��}��0�U�E,*�c�]k�*����9{��ᵇ>��4.�����TT����C��.l2XE�*D�a�fi�zn�}���B�����g�鞔f6�29�m0��.(���Yg/��\�lv�ۻ�0�{vK���)p�vϩgx�9 @�2��1�f���}*���ϴ���~�ka��f��q�,�w	�0�U��rv�Bw3��&�#����q��~�o�I4#�v�ۥ�yE+��B��"8�o-)�TWk@��C�RSfm�줟UP���7��~���+�>S�EC�#�f�d�
\M�&��-t��2|��V]</!n�o5��ךђG&��+�By���{���d�BI�J$��A��
���z���f�=�3��˷8i���̭�⛷��l]㡵Yρ���I�	a���&DL�R���N����'n��+=��p�kt�\�l�%c4N��v�#�uъ�(C�D�����m�������4�Z�|�-Sͺ��_a���1���~Yܷ�Q=MP��=�����ǵ�M�/w�[Q��y�t^�On���j�u*��2e��ƦzJ)�>���9X�[gh�B�*[��Է��`�,���M*����U,�}t.�ʧ����o\fЁ�^{|'7��q�?y���+|=�D,�\�d��n��2����<B�}�k���T︼Z��+��J�[I�.T6Wͣ4?"�9a����9��}�d�3ߙ�γ�Y��l���7�sG��7
��y��.�(�ӳX'��)U�����vFmՑ}X]WgP��tn�[�Ժ�'c�k�1��[��&�6�6�;\�U$c�a������Zk�s���\����<1�Z7�&Ggr��Øw�C�Ck�ʧ���9*ͳIT�_b���?<NMU�$;'��G�����{o����/Z�ޒx�Trf�l�2�~QO�O���ީ���Yt{��=��xc{��&�:ܥ��c���i]{rO����`x�"�"2��j\���$�`9���X'n0e�U��YDDH��d��k�%I+�_��a^�ㇲ�M3/�招�a�g�.`�EK�-
��}�4�@�m�zXt�x`�\�8^>_~R��1�j�Q�P�F-m&p)��C)��^H�����c,���W,w�c=`v��K���<L\�ƹ��8�b5P��>`�K��'A�����m��E.�g���Yz�6X3a��< OWV�U�]�%���`�Vk��7Lq�#�$�ِ`'�%fæ�~s>���1��M����HE��|nٴ1 T��{�\u��wL�ԍ)���9"2*�h�t�C1��r#��p���g�zG~.]7&��;��� b�v����+W�݈��}8��b������Į�mO�L�ͳM�MK̠e��b)�4�ϸ��wg1�O�8�����u���"+�,v{E+���2���o��دFS�O�w�kX���ܱ���cKF
T����@L�"�]�2���b.���;]��V�d55:vw�}O=�EWM�$�����6�s+��-�P�Q����u�K�*�KK��N��g7a]P���@@����;�6��A�^�A�w�M���=�������&}��r���8v�י�bL� ����8`!���^Qʑ�������j�$ټ<�J	�����upE ��0[(����v��5AgN���[̹���;Ʒ��3���Z���ھ����s�SD�]/�"���oF���j�cs.�s��]χ���MG<�y���׺�^���ɚ�E�S<)$o�޾ ���>���Zf&��=�\<�ȼ��ݼ(K�+��i�g�VT�RT���R���͊���/�l�>�o;������܊�Ⱦe
��y-�O\�&g֨�4�E�r��=FU�`�ˀeR���V�gewv\��B="�,�-�t{-�4v�1���B<�������"�D�
�C�ۅ��TԒ���Q�<���/^�3��cP��K8u �K�l�Ym�z�`��Cz�q�Ժ���r�
L:��2U�EkP�GZ7/�R�C?`x�϶"��^Z�3��";��Zag�o0��8�wgc	 �|�~�Z���J\�vfxE]�+|7��=�kz{;aû�~��K�&�1t�p���wӐ٫������9�����ʹ����Xr��:�Z�e'm�kA�k�jǬ�Z� �ɸ��� ;�*�>��`��m��%��X&�ђ|ѥ�Փ����Rک��Mvsܧ/!0K�|}����K�9��QA��q�#�ǃ�r���`�<��$˱�/2\�pkdT�x�P��ݐ	8DQ,!9Vf�fo�����ס�ϏBl��MM;I$!SdJ.����KS(���������V%h]�p�#�Ƕ���Hy^~.E�J���ڗ݄p���z�����c�r0o�H"�����k9�Wh�/���wӫ����sF�DOӤj������2��*�D�ƞ�3��>;j{���yq	;���N�ax&}��2��N'�sH�"�����Q(�"'��N� �B�=�/�[��c}�w�r�u���e�܌*6zK»T�CP[A�^��S1}��I`γ�Z���
�˧�z%*�dU�<�)9�]ε��އ��uL�&K7qu1�E������w^Gr�:5���HrK���W|m\!j��pB�o38�ٶe�Q����MDl�Z�N��'*�j���q�	Z���%�GI�Ӫi>�~}��������u8WR��^��pt�U��M�X������1t�X'�y���f����$�|5܀�[BI�?0���}%�b�)x]T�=U*�gN���v�
"�@.��%@.Қ���VEA@;���W�J̑Cx��.�u�ܤ'@���6*A_&����o7*x�h������]TV�C�(J� �d�����i9��l�%7���;��4'W>���H]��� �H�qD-2{�w��;&Il���ӕ6��l����9�K�8����o��#v���5�BE�g��p���R&��x�����6t�4�����y�iy�}G��o��"�[�
w��E�`�^�}�����ZYf�,P� ��50uq�6�wMAz��j;R5���~�&�=���v�v؏�~M<�ceC�֋U�֞}�{�S�4�,9���PL�k+j;�F��щn��q$/uCmWʾ-�����\��ХR�[���{�2�L�é�aU��(��v�����O�rH���x��_{y�v�
��Ck	�CGlv��.���=��ʡT��{c�v�!-{�t&��C�&�۬Cv#��۪����R�

����{��b�lŵ��$�7K:��1����Jϥ�D]��_;�*�:��b�^y۟d� Uf��O�3��V�h\î�!=��S���FОg�_�W0�e����%t��w嚟u����������XVf83�2f+	bG���2=�l����Tb��$�y���ߑ���:��ж�䈒Jʤ�H��&��)j=�K�s�5�U�.��fN�������{>���u!؛ �؞^���U�q�
n�����&f/e�ɋ��U=���@���Ȑ`C  ��8(�c�Ef@ߤ5]�F�����=�e�઀X�2b$�A$&�dUP`��g�����f.5k4�庾�M+i�]�� '�Ѽ����<慯i�i| ͍�:�&���/4��� v�^�.+})Ծb���ˈް�苋��8Se�%�h�W>����e�Lh���ۺgzzس�B��Y���+���f�L���vv�9:�g%Y	g�?��N��}�F��9~�W���Ȥz\c�M�����|�T�T�&�4�*i��a1�3k�wS�5����R�.���<}�(|s��e}����p��N���u�'�ðёxCp�¯�����-�J��ڙ��۴�JC��������l"Nq�y�y��Lpwk��ITf��� �iy�8�J�P�Pл�ܵ8��{t����������Ulv<�o)7��]W��;�Z�8��c�UsTȼ{�5��f|�>o3o@�+[We�\IN�e3-���-Q3�Us^I	{�|tF��>	u��7+V�O���}*�����u;;�\�a�
����K����Iz֔�UD��h7��w�!7�O�r����k�䶹��Z�"���χus��̪ߑ|0��O�;�V	�'W�ʞ��O�}i!+F�U.@��׿Pƌd�\�ǎ�f�����_���Wj�Bvt52|��YA��)��t�95��Ǚ�#�^�4��wc�t�1��RH�}�&��O�ot�����Q��M
��L����Ýdo3/�M(�]Ox�:����|������u����F�Wc,7�WK��c��OV̛��]�,4e�����,t�"FE� >d��}>�Q$����bPTO���㐖���!��<h�N�c��;��Z�6W���o��][6��!okS�ː�D�5�eb�6�}U�v���)u�BR� `�` ��}W����s��^��>n�h}_}�w�N���fϬ?�wx�m<,"	�Y�dU��i�*��0�ѽ%�-�����j���rY����К���f�jF}���r����}p�M��Oi��C��D��PzM7����%C+S�u�l�+oW6y��<����yJ�m�m-�Qݛېy�ݸ��jb8rףU�DƳ p^�0�T۲v	�ˣ��Lv#-N�h��#����_P^v~�9ҽU�������^o=�G�v�>��-�}��O���  ]ՋO!�_��|u��P�d�T��<�>7:�L&M����zw}��E�@�.�C@�*�)�1="Li���،<����@L�qCT=y��=�l�U#������)Ϥ�8�T��\^��C%�٘��{��G����pYB�b.<�!߉�3>ѯs=(X��\nݕ���l˕���pzé�� �@%��0� r?�q�V*��:�J��˖�R���ٴ�͜��X�j�O��y��@�0�`	8�z�
yr1���=�ji!2�sCӭ����v�b�z��6�9�/���vdkv��i#`�yDm��0�/�����]޵՘��Nq��-��T���/6ފ`ز7z��r+�4E�!L���˞�c�dkﲫ�b7so4��V��������$�%2H�_;�Wn�/�.���NVK����a<�\���'��3���C?�;��J��V�X�og��[����N�����z��~�a�9�U�?q�<^�.}�M�7��4�4��v�`Ԇ�oeUJ7�	�~��u{�^{�s�;ӾJ�}R ���$�?o}U�Ed�{��5�>u�+��QT�+��9:�}�|d�U+��(ܮqjc�J���SZ�)�����^4�d���+ݾgW�Z]�#��g �[�̞�a�xݫ�ހ��^�Ri�G��g�"�1p"���'{��?X�Җ��uM�"�6tئW���q�X����Ecp{�(@v�>����ٙ�h�0�^�0��C�=���EW��E���w��v�r�K��ZUk뺵+\Y��oo5}*�4rS�����#'ӍJ�6�JW�V/��3ǩyy%�Vi�3Yn�u�y��7���
�Y��,�^x7|'~k�������E/��%D�d�fd�f}��H���K<Vn�Ǭ@��$|@�"}MK���6����u�5�k=����^�v9F�A0L$$��X�i�Y�F�i^�qJ����vD�f��nm�3�1h
q8:��ƕ���Vղ�΢t�k��%��ڭ���0ϯ���-C�g�����|E�&Y/~�^�����܊�:>�ٝ�X����"'�MG2ޢ����S*i��x��� E���4}�>��x[�>��p�}ó7C@�ѵQ�clxNs�-����u���&A6ۚlx�옒�a��,���"+��wc"+39;�#�7S9L�f{��v���4�<�c�IEs�]Ϲ�%�$E���B���c���g��!HM:��[�YN~#沛�m̂|YԸ�P ~eAF7�j8����瑛�[#��2��l�<I�L�ʕ�B8��gdא� A" s.�\�o�T��lqo���Κ������^D�l��B�*�[qc�j\_�2��_J�Ѓ�J[^v�!*��Ԭ��ΖY$�����,�Q�rV�,i^N�b<aD�I��rgk3��/�$Ob�~��]�b�����d}�	r��G����
~(f<.���;bo���g��*a��>[(��'U��CW��9b�Lǚ�E	��LhF�y�y=����\S�4��7�N]�l��α�m\�d� 8�<a�����$����>���Ʒ�L66MK;˦x�3]Nf�EZ�
�yv �T����s�B���q������
��]#=NMy<����@"DG� "#���   �� "	��"""@� @��� D&D@ P" �� �" ��@��� ����D 
1""?� "DG�׀������ "#�+���������{� D@��1 D  ~��  "��o���D�����0 ""?r=������ D���_� ��� ""?o� "#?�,@"DG�_�b���X�H� �� "#�/�_� ""?� D��~�����Q#��ۀ ������?}��D���$` " DD_�����e5�`	��hl�� �s2}p"A�|{*6ƲQ! �mD(T���i�[MR��VR%)H��R�� �Kf[`QR��B�T��R�B�KA�@U%P�@ j"��%Ѷ*��BUP%$P�  U(�Qm�UT������U��J��IV�@�E*�Q4��M�H,�*�@�kF�HA$U��zh+�"��LUUtl�X�FՅY���@P��Da�e�5���֕5�T*�4�EE*���ҵ"R��IRD�����   aX    �����5���SY�J�ʩTP���wj�A���Gfj�jI�U6wj"�B�NثU����%R�D��

����]0EKm]hUU�k�C��R�p躦�MR�e�a��r�bd띚�Ƭ�;j��b�EZ�n�T��v��n�J�]���1�)62�����T��T�ڴE�*mfS�B��[�ei�c��u�ͬu�L�m��[L��h�[V���'Mۉ7u���G]�̌ T���
,�Y	�CL��2���Sp �im��@t��TmJ.�wr�ֵw\)�L i��F,t  wI`V��M�m PԦ(���("H��PT�T�*��h$S[tn 4 ��@�N�d�]\��ـ�w)uJK]��h� %��4�:\�hQ��n��Э
�˶JEH! U�Ъ�K����I��)gNp4�.�`4�w�)JG+4M��6�6�ډ��R@h5S&5AѥY&СE���Q��ٕ(Jk�I���X���uU�Z���6]��E�+!�R��ISavp���T���ATU�`�6�(Ɲ:�Q�v�bEk($�ZP��ͭd�v�-�]�Z�n  CL:鶠�]�)�:�&�hE�2A�V5Zm�s.�h:b����qr��t�]�S�)ѕ��D�Jm����BI
]�ґP$�
��	4փFj��V�J�f�����t�mݺSnk�3�%��K�P���Un�K����.i]т*E:9���K�E4��F:��K98 �  ��U�      
�ѠʥJ� �S�0���C1�#�  T�R��F �)�!�@@1%"P �WbG!�LDD�R�9Y�bL�U (1��p�T�>f�bே>w�i�����"DFzG��@�""& ?q D���"���@�"" " ~����~������2�$��DL��V��#�*cɒ�ou*������Y�Ac�ad���b�ǖi-wvj�FM⥔]�Ԇ<�L�r�n�b
�hê�ݜƣ20Ԥ��U#�ȵ�LT�[F"��)n]�fY��!-��n��)1�H�/�vAW��t��ܣ&�1��o2� ��Y	���M�F�c-��t%��ە���Sy��r�Up䤀Oͱ���VZ�Ń; �>g_��̹��K 	%R�I)h)B[5�f�����;Yf��ZTC,P��	}�@�M�r�����gX����@ak�*�SGj^��p��.�k�5)��5w�f�H;T��jYM��J�����6dM�k�j�4)�^���k,��R�"��ˍ��VqV4.;��Pvg*S0�MZ]�����X�}t���kfB��zEeX�Z��!X�ꤠ��021N`��+[G1��%?����ܴ�6Q��+z1|#�ҐPh�-g�u��;��n:S4�p�/��i��J��"w^���Y���b#{t��jFx�V�hլq˩*]���qB����;8� k6�E;CthM)��4�8�ѕhӬ!�_��=���-��t�X�IІ�X��n�!82�%����Kp�Ҳ�7M9�1��Kk�m�0=�柅IL;zh�ufV�Tڼ$l��t�����V�f��3NZ� :Ԡ9f`*���m<�On��Q��K:7)c�B�]��ѩ4����Y�t�a+4S��˃�-�f,|B���J��3YJ�tN�8K�(Z�E���c)�ѻ�`�MΪc��I�$KK�ή*B����=�;ܽ�Mk@�6�B�4�j�I),J��0�X�v���]2m��ᦙv�J�0���^(W�w,"�Fj�¶e+��,ɧ�A:�2��HJ�J]�n��*Y�L�P%�-p�ᎴfYU��DGu�$��D"i�kU)xA�}B����wZn��fN�(Mu�1 4� *��1E�:�`Y�RU�H��룉��R�R���������KDo"`Wycwlj��M8��7R*� �ȱ�(Q[��$��C+V	!*d���++�H�,�b'��ɥ1���BCoEF��p�S�kҢ%��mW���Gk&�/b�KU�À����^�N�!�F��T=��n��S"4쐜�U�Ϳ���u^M�I������U�v�J.���ּT���x0C����ux�a��o�DnE���.��û�M��U��V�*F�N,�
X�s��c^���-�զ�wC2�jZ,P0n�Q��cI[#�'��w��\+�nm���*�Ү=�!F��!$S̴�[=HM߱������:�ʙR�Z�`_Z��	�*|2�w�)��q`�62��.����#-��ucj��AfH�<�0a���DLChZ"�����f�� ̦v]=A���Q��{bmL��U �+0ޢR&��1�f�9�)���lGQ��'z���6�1��l�m3��Vm�#�t��TG����X���"��Lru���ڰn�i�!��鋬JKmb�Y�*�',t�,qB" �s'Le ;%��cy@��"2����ջ 2#E�Or��6��d���Z��{$��i�BV�U;YI�M�#���V]&6IDkg�N�GQ��k��Yz��PN��oFT���W�[�	�ȭ�OQ���]�jʤ/*�Bi���f�
�"CJ*(dR,�J�Kn��eh��YpŔ��gm������u��8BT	�wB�^�&�1�jo!y(�x�$�0V��)r�ݥ��Z�n��s\�%� 5�!� P`�O;�S)�y�) vqmb)��;bn7�o2���%�h�u"D���+�'����Zd�;�1�Z� C�FX�h�ͧWV
)�-ƪ�ҫn,Nǒ��0���N�2��whk,U�h�0&�[�0򒤕��{q���$⠛��\E"ټ+Fޫ�	$�[-d�*�����e�Ǘ�ʰe10;�"e�A#���#)��am9wr5q#�%�t!�y�&����2,�z���Z%�

������[hK��)�S2�s!�2�Ʃ�l��[�"�v<�0���`�X���Ln��h۶p!����fEz�S+v�+WW�����Ռ����[��Coq2����0�
�.�[���LJ)t�n:�!�t�ѻWie�yu��(�VeIzo	l;����jN��ѓ���-+&�T?=� 8�@7,�(���DT�OP�)D6�?-ҙ�oV�C>�A�m�+4�u,��(�]l&[yt�`@�6��؆�Vл��'3Ꙣk�;-d"����5�x(]K����zj]43��
&F��if+%Z�ݧ3YO4�<˱�$���̻�h������P��̽ Xv݅b@�B���XU�t���`5��4�=�N������q�ѰJ�k�M{��0�����u�V�t���8�s��5��w �0�R`WjV����ȮZ��k!5��R1Z����k���&��ʕܷ!u:g4�q���ʙ*ܲL���*�(&W]�U�	V�!Y����kyl��C0(V���*z,U�kD7�����7l��t���VZI1W[3aNBN�\*��
�_���8Z5���� " ��0����� ��`ל7���X2�܅��Q�^��Œa��.��A��US<!�/uN�̵(�tYFf�̽�x�-EN��gTUl"�[Q@����I��{t�"=S17k�na.;9�X��N5��|"�[>���՜���*ZH�a*c1�����M�O�vwVw�C��n�Q+q<Q��r��a�K+7i1kZv-�iau3vVK2����f<Iܗ�>;�)E�(;�'l̻�Um�h�r�p�qYHn���"�᢬
i��-(�Z1%&^4�Z"���p�Re1sLW��y���m�@,w�TN�����R홛i*����P����9�o�
sN�oo3��Qx�)iT��1���;l��v��&I�`M$(ʺ�W��J�h����ؖ���9N��W�uN6���+v��B��p[me�zwy�-�o�*i9P䭁��vG�](�*��+�Tx%�{���Kqe�f�c̕j�4ܰ�i-�V0�{6��u��5V4ˎl
BT���t�ܺ�gB$S�q�2l8�8Z���q��L��r�L�o~��p��7qRИv���j�5�m�K#-'�);��X�.v������[��+Rr],��#t��ڍ�@
O.Ji������&ap4�\GbK	ّժDU�{��l@��Iy�j�nK�FU�Z�Wse,q�����[���pPst�D���~j��@��Ɔ�v��)��*֤G�%awq����lPV�A��`MZt�LZ.^!��L_
ѭ#�N���,T�0��f��,kM���ZMKEmmcn�⼷���R�e
 �InЂ]��j2+s,�ݩBh
��T�fTR�b��I��3A,����t�Y8�eZSE7(h�� ���[.�y�z0�kMe\Q��f,�V.5,�ӭ���aX�)�w�#gI.�<��h��9 ��8���.�m8 WNv�j�� u��Y��)�S��>��]]=���4�T���.��S��Ed��7u�2�p��mL
Y�DG�S/q�M^c�;�K��f��S��%��m�9r�
"��n�Ktj�vCus�����jي�lWPl ,QD��2m��H)�jd��q��l�ѹ�̨�(��ܳ 	�3Fj+�y���q!�FZ�q5,9�waǸ�ݔ�Z���P�Tk3U��2З�?l�S��7�F헙�J)��f��qe��H�z��L.����7.V�im��&-RR�a�w���7�ee#0�jwu�t:�g%X�����8V��cA�xH�.�XW���NwL�Pەv��j�u�x�[u(�٤��l(�/��#Py{p+Z����f�&,�GiUn�Eh�"ܠ��j�ܫ�RhV&�&�A����Yos��6,���D*�d�l�i�%)lH
����l ]0�ֽ�f��]^�5jQ�%訶��h��vf��ݷX��]�Ǳ�Yz�RI���2���SspY��_�5�@A�ލN�!��[��iY٥eҸ��-a{OB�m��H�y0[&�51L�yv�BDN���RF_��n�^��H�! j�{[xѫ�
ƀ�41��\6m��4V��N�.�-�%�܇I5z��5�j��i��[��0:�7�-A��YqA�.���4T��
��WD&�
%�ڡ�⎢OQK�Tխ���j��Z�ı�7`���*Q;�r��i��a���=�͸Χ��SP��R&��&�J�,f�����q�Y��%I#?��1^6�3l��ݰ�ys �Mi���F�,�Zskb�[�K���9z2ΫX�6h��'�:P��:��1N�aÙn��`�8�o&d{�lZ�� K:��d��$7lGL�r��n��Y��/��+.6����YX���ڙ)�2��K J�ސi�4� �b��,�	LwIm�mK2��`�2��5�H��6�4�&�fd��-��"�˨6�c_�%��oQ�,K[l�ћ0~I�X��.��p@UZF����E�)Sf+�-]ފ[X%jE޹��D2�)n/��oE�]�*F�j�WɣtD�E��GFY1*+Z�̚%�X�R�ς�B�.FM%�.����j�V�! �5��2��cu`:�cE�q�EC��wUC��2�EGj%�k�-9u+F�Ў� ��bjU���RQ�
pӭ�����eڰ]�FO�V25�%fo�w�,y2�n�v�d-��ug1L�d��xl�O�(�2��E�f���+T�AX��@�*i��F�島���U�'wbK�@c��0M ��v�ַP<OX;W)����nH&��P)�bU��n7WP�z3]�F9V����r��%�$�ȧ֮i1&��
�J�Ee�)��,x(R@Va�q�Ǎ���?k�;�Xvv��V�S@5�ke�вnTӃT.�L,I!R��@M�D71hNh�iǔ�2\�wN�U��%�.��^�dBP� �&��WI�\7�I�$X>j�ۻ�b��{��/U�0�*k)$���2^$�EA��d��w�,�B;����B����"� �r�^G����Z�ͫ��Mw�v�EhRa`ß��Q@���0B�%:�bV�ͧZ�YIn�����5�(!XF-шUML��Gn@2!^<p���4ehN�-��w.EiTK*���})��z� ��AN
��͋󧖖�h�R�rd�nVe�ɴ�Uv2���n$��M�f�H�!�
�-�-�ok'FIJ�%�A����jA��
<� �Z*:0X݌&X2�T��v�8�\�z�M΃����ɑX�lF�9��C4m�,�mp���ၣ9�)��ݤgh�&z�(e�2�ڻ��`V�I���2�ŋ���j�g�����M����F�[	T�wK�����L���
�j["��b���j�)��V�u��nG�6�I������e�ͫ�'ȧ�sU8[E�^�%H�u���U�T��B�k!�M6l˚4�BP�K�
���D=�f��ц�d�&1$cú�M͙E�2[ؾZ�'��F7��;(��dXud�r�7s.Ӡ�V�DK�+o{r5�7���#��%&wj[�e���Z��*_�9���K��iБkÂ��F�=E��&�8��Xܼ3!i��]?�M6E�S
��A�	��o�_JCoKd�7.�-��Lh�ø��/��y:훭�K�
�0��6CV�+sF�j�5"t���������
IG�Gf;���&0�Eh��Q���J�޼ȷDXA���ah֜��TX$Cc�eF�C&�0�Ϯ�nE��caq�u�;��cl%�k?]2H1��r���lZ��۔���%�7*[��YtMEK���8N�K���Z��8d=���RYR䖙X���ȶ*���N'��t�Y�r1�m�Ц,=IԲ�٨��l�)���Ud�E�cu�R�ˤy�� ���xQ���3�ⱥ�;�/�V�Ո(��L�� j�a�!�M���� �2�KlHg*�q;ʸlR��e[�5T��%��/DP[����2��)�L3�VnJ6��):YO:(���픝��L2�Z/s��N���/t �M5/E�Jg�e�@�)Ppܷ��n`/���)F�MY��;N�����%nf��0Y"�9���	tk�FIb� ����-P��X��0L��ɼpo�֤)�_W6�u]��u����ڻ̖� �ŧ�wa6�|��.ևKE�Xuec3h[�H�E�]�m)e^��K�z�3�oK
)��3�˒�5013����[����;lY��Gb ������
�����ƨ�Y3m�tҬk�Yr����Ť�'0�Qf��75���0�U��ǋor�o N��*|���4v�*�	�P�Ij��`t:ܦ�2�%)���U�9���Z4:h�tԭӘ��[��I�n7I�#r�Fe�k�d,���s"4`��h����[����uk��T0a�I��B�e��n�n�p��ѧ��޼�L����2�(�XGA�H;���{oFm�sFMP��h���؎5,K�S1�O��R�i:Iŀ�K�yZ0EA4��Xiކ� ��C`�aݡCe.�����`sm���TN��O`��S�A���8�St�=NI�Ss`����cov��V�+�"����݄��ov��Z�.mn�yd]�u�����U"-
���Y��xd�F���W�����	��1lPؠH�C'm�:�;�M9�����7�5�������	��I��}���.\ ;�`����9�$\�k�H�I�#}�p��l�q���ܒ7͞K�c��%Jnf4U㙸ck��|�H�I�$}$��K3''$��Ӫs���*�t�F⤰��idʍ�R�$���W4�"���i�����]9tK�siո﷗&�2to������GѴ����j�s9(ҏ�m)�x�t�]�m�ϖ�[m��v����nI�ܐ�r]�'F���;��ل-<!��Y�^YkN��(�M�%�`ܮדw�������oac[�9�G+ϼ,�^+��U��Yb�]�uO����]X�%��)��J���K�\6���*n�:!I[�ܴ/'F��ckF��;@��e���LE�,�y���j�/o�,أS�%��F���=�Pu�lvD���Y�d��
p��`E��+o�\u9��>B���Mkl�V��=ۗ�	Y3'��6po,���� �Ub��tFeN�W+��0i���9Iu�] 1�2�����ji��y�9���%�0���W��9t]��x��˫�8�mst�=̫��e��6���6n�j˹�@�u�O]-���8<�u|�5I\| B��v�=��z]��L��u���$�
��dK�����^Q7�������LQ�00�L�\��v�ƃ[���ܻ�?F��Ͽ+�F�D�en�2���t�H�&_�^z�i:��V���p�M�זwe	�Q�ެ��2�n��3��#v���ayw�b���:PܗV���@A�����A\�E] ����l�P�i�X�|>�)C�>A�=�,WA5��b�h�Kp�[+Dz�]���X������]��Kyw-y-��k�'b�yu��.4����35m�Y�j�}�h�΋Rp9ݒ�!�J�l�:h��E��S4n:��/�������6��{%�ꥎoB��/WsKH���f���=Fq��.��_bCVrk*��pu�؇gQ�<��]}��:j�/Pǆ�.?F�ή��݁W���Ib����Pf�Y4*�wj��"J<c��%D�E]����!��:0�,{֬�;�&M�^I����� �W�փD~��o��M�t�m�z;��{7Q��qGSM��7"�ۥAݬ���!S'r�g�.3m�x(��Fjǐۧ��t�]��[��^�J�۸Ws���(T��zCi�����b��v����$�N�w�+�ŷb왱=E\��AB���H���Ҷ6Px�r���t�SY�1_p����ϭ,�j��y �ɛJ�4;U{����q���[]Xzuz��}/1��&�e��tk.	�/iȇRY&�+�����"�V��֒љg�$�f�Aű���c����[\���.��JG�D"7��v�c���43��s/{3��M
�2G���f��Y�r�3֣N�ax����s�2×5TF�2��:��7Z�B�V��+����w�Z�s;���%|.�늴���R8�(Q��r��h B�F�V��j�Mw$���$8dKǵ�������*�CR]��f��R��B�7cf���ىN���]�; �MwnM��R�N��b��V������[&X5���;�-�g�m�v�8�bM����嵧t��ț����""^��]�@S�R�u��V's��`uZ�ob6t�V�+���kR�v��@{��{��^]=4�7B��}�6��+o_rq���XV�w���@�Ӕ����{��ִ�=����PP���@��f�k(�\Q�/O��c��߬+�8)/G��;ۭ�\����ˈ��+��agy�H�l^a܄�a��BꎵJ�7)cü���t;M��D�Gs��,��S�\w�m��M��Y,v��ؕ���m�[߻F��аE�*N�vqޡ��L ���Z ��̋&��	�,�*��,,Sщ�z�NM��)��n��g.����U�s��a]�wZ2ҹ2�K�2���!v7�Ay��p�um�Ȼyb�'�=mr]n�켨�2#��Vv��]��2;�픲��k�� vW&�;�e���젩`+�T�.1�/F��k�Ts^�0���0}�����\ʉL��M]�q�����6�uc��V�p���=�,�ڒ��8����@y�n��u�QPw,*�ҝ	A�YZ9M��θtB����WK���0dA�gB���p�-Y)@�����BҘ|�De�]C�,��-��i�ƶ��W�����u��	a���<.�5�U嗪�v%$YH�'63�l���Yr��I��,�ρ&��Δf�ާ�PpS��R����0'g�\�ϸ�l��Z�Y���	Юyo��c&���V��e���WLG�J�{E�i[�Ǝ����F�ܒ�)��1o15�-w�7l�ܫ�J���mԗ�^�e��u����YY3U���t� �H�2��)S�ov�=����.�4�NjVQݱ���/��#��m���oϊᝳ�ދ�jU�3|��΄���̠�6�a
y��#�{�
��M�}E7�ӻY�b���y6�U�r�b�Uү���s�]��N��;��w��yvj\/�����u���!�$
�r�ywH*;sN62ZWz=��3��\�&�C����j��6^w�Y�����IM����B�:�s1�-a�������0�Pb�RM��D�iX�:�-]��r1�+&����5:�SbM0��3QN4�����f�Ա�=)P
��;�˳�:DWYם��E�� ����l��}�tٳ��[����W.%���;�^Ս��1EnF�Q��#�a!K��G{mWo,BJr;t8@[|��n�m˭'��yU���v:��S�Lt�r鷜Z�N���	�o��P�hb�.��<�Y��|5�΋��Y�*{�fsb���&��43�,�9����;j��	�ƶ�����
�@J*���p��:�,9�<F�^�� Ƴ�K�� �g�:���5S+L=-Ǳ��%2��\�[���Q.�P_��I���gr��r�*�v�u��n�+8�>C>E_�R��嚮jk�_Z���¼;�/�jȽZ�䌮J+�R,��v�m��qáMȈ�I��&�q5G3�L��]L�`���IО��Ry�_�&<m�*��kTDp�*[y�������`č��1dw}�.�+��8[�8k�Jm�b6�;��H�p���f#���
.l��C�t�$nXZۺn��$�ږ�6�7bB�=��s�+�f>���a�Z��z�gT��Be���c�Ι1fM�!�ٽ�zV`얶VKxs���V�z���<�t�j��������XQjq `Bv��*r���B�N��A����z~; �U���:ҝ�{m_{-�Ь��d�V�Y���x�]�|d/�9���	�j����կ�e��Zf���.K�G ��։��h�0�e����;��yv�t6�W�+Zu
~���wAC+�3�D�B�NI��}]ݙV���!�#�ޚ�hVI^�n{/d�,����=YT�S0Ӯ�Ƒ*�b�s�V�J�\Ȕ�.�튀��r��O5l<���+�����Z���b{��n�q�I]��R&Qܷi�e������(��K=�ûj�{��������������-�̨p0�f/2��~32�alɗoOi�VZ�]5�T9Y�F�\}�۴.�.QwJ���륗�N�M�w� B�<�V�*�n���(EIԙb�K��ه�������Օ�q��:��_��./>t��R�2췽�J5��7:�+�ێ�5�_f��É����Rd�%�OEc�te����j�u�5�����3:+I����@�I�}!\�=r�.�,��/�ǢV.P���Ϥ�c��i�U�������	n��O�)�N��3l���%�嬍�����"��׷� 4Ԡ�3�t�Sw�וvw-�vL�$[X.���7�+{K�Ĭ$����@$ӈ�m�R�<� wW]|u�^>7��jf�"�)3��x�`%M����Ƅ[����}������!`����qîS��ۼ�;%�\*�v��5��=��n�%�k���F�Y���T��Z���S���9,f�Bg)�ؠ�X�݅�ց{��K�A���k�� ¶[��11XwGJ�\���t�iJ!r^��}z�!�VR�ύ���$��	n��V��O�	����Y�
4t��u��?�c
����ҙF�!Y���*��S����6�K�=K P�՗�"�fJ�݃-īB|)�����L�`i<��e���*�1FvfI{a]=	��MKJ�;�N'{�,>Y��*�7��{�W�Q�>p"Aͅ#�c`�Hr�(�޺W�wټ��M%� �	�#��b��	��md	n_^��]Cx�
�o��{Á�G/bwo(+���N|�]���)�z�����l�̲�о����}b����T�&Υ�9m���^09�[��μ�w����R��8n �yM�6Sr�V^E���]�fNdm��+a�~ݎ6�ak�Ǳm�5n�m����Vv84��	�掠�v���z�w2�m-��=c4��P���N`f��S��tT.��u�W՛�,%Q�>.�`�v�W$&b+w��m�)
͈�-5v�uOT�n�C˕�����r�Kh�x�;���X�-����OJ�s+�;����PR0W[���;os��6��PwSE��&���;�r�0�d:a639.u���ӧ�A�Ed�oy;�4��`pM#j�ɏ�ʹ+�`e*XG>��˳�ֺg,��J�30�*)B\��GB��s��ܖ�S��A�c.[x������
��f��pVH�?�Yz�냻��`��Voj�3�#V7f��Ĳ�����b]/��/ᑒ] .��Y4�Q��h��v�]��k6��q�3 v�J�4x6����\n���E��&tSg��u7B4#V$���@
�SlU�.��+��H�+ \�i]�!�glX�	%Z�pҫ����E�c)�����K���ۍ�D&�#3�R�%r���gܨ�������r��::�j�8�ڋ�����) ��w��yC`��K�^6��r�q[W3 eҵ�d�Gt��ЩB���C��K��Z6m2+	�H��r�˷�Jl�q݉8����]�7�[�n�,�Co]���U�"Z��>q����&
utܲ�[{�N�ɕ&�3�[�)v<0<����b�n�\��aL���S��t�U�s����;[�A��PeM��X���O��Z�-�.����Eb�侶gj����y:Z�R�ӎ��p��z��qb�OZb\��ݥ�w�N��V�gL���[)�8��f��\�q��AM�I��4e�H�3��,RI�ȫ�GA̭�Q�W��?{���K7�خ�$J�+�&��7�WS�;E	/�Fs�U<ץ����Ȗ�՘%���Z������D�e[ξ�9-�����G6��yy��CgV��Z��7+t*�UvQ7�P�	�RS��������¯@�avz���ƆvJ�R�])�]e^5�Z�t�>d᷊��ƚދ�"�ԯV�0ut�L,-ɺ`���_>�i΍�7N��6if���L��b����مWW��h�2�˧@�y���G(d�֧���a�R!%��7X���أ��r�V���Ic��VPWۻ������W�ƴ'����O����"�PN�&l��_Q����{7��
B�][%�n���w�Z"��)�HK�#5R���ՔXq��.:j�R��J�F�]�+i!;�yփ�}s�&�H�׸i0�6�'�aT:�+��v���P�ղ�4��V�e����̵Z3V��>��*�u�� � ���L�M\�cA�{2����+"#&tK��j��n;�2��\u�*1�������4��

������s:����w*o`������=hZ�n_)[0+jAF�����C%��VJ�#V3&��R�+�rqy��{E���sV�^8=���W���)
�
GxyC$y�Au���3{��gP ��pJb`Њ>)�d�Y���2�]�}�k1ڕ-��"�������� ރh_LI��n>wVL��X���o�l�ڸy	̵�^h�#�%[�Ț��\6L˜�s��N��L�ڹih�Ukz����r�:�;�O��l�\�����u�f�ձ�=���u���*�{"�"pu�8zcOP=�p;lꫝ��C��t8r�l�9�53��ʶ���l�Np=f�3WI崭����sj���S���7.m�
ޕ��jt=Bp�Ŷ^�*�����a�Pc����[��_p�Ҏ�c$���`P�J�r��`U��S�^w\�[̾K&�����l�=-R�t��;-`���V���ȻK�^EYYvyLZ��;9胳h�$W;�xڋo��ǆ�nC�X��o�kf�CP�|�@�Ԏ����vqu�-�]�x��Ƒ�#E�X�:�6s�/��kiQ�	7��Y���[���[U���Q�Sb�N�f�X�5)r�Y��ҔP�F�J�����Z,p��}z�@<�b��h^�)}�n:H2@������1՘f�]&��]YX�O1b��g+7:�{�Mq)�����۔ PY�?^G5�j&�*_y=w5]�KOOwj���������W�_v��H9D~t�&��Xl��E,��aԖ-��${QJ�ص7e��.q�����K
����߇ly��`��_��Am0����y�mP��F�U�g2ƕV�2��F̎�Bc��B�m��}��옶���æ�-%����#W���ZF4u8kRySxb�z����v�L������M<O7�L^u��a���8AhMΥםY�v�̽�D��Yʻ�K)�̬��K�B��}�n3�(��"$U�˙G/c�`�1��-n�Geff0��Q��˓;�C�89��'OR���+7-�껆�Vօ2�n�DROV3Lml,�Y}�vVu�m/ۇ�ͳ{J:}mApes#+lJ����Lҫ7)��a�\0�y#���ݖ6�Y����u��E
�<�u�%B���吺���͔��h���cμR�:�Yw��Ӽ%�藖s�8�� =" @�D@�""G�� 
����3�f^f
�����4ң�:qB6�k1�շ���s��qy�[�zȴ������z.�$̾Y{�@E��3��r����T�:@yWl�fg!��p�\�/��N�w���@�P�[�c�*5+��E��Վ�A�i<O��B��+yl9�voF�G�u`�N��֣e�-�c�h�X���X�;�o+YK }v����Q��}Vi�0+��U�֫R�E�2���Ɯ;�m�Ђ��շwy�:'ki��Et��/��f�K��oZ�����n��#ט��W�7�a1 �O�U[�uڳ_7fu'�gbᛑ�5�ChC�!�&���:.�;�s;w��/���'-l��!�wp9N�ƺpC�Z$����ltU���X�2��p�$�.�u�Hx7Gc�{�Wc��b�Љ�*���[�d�]��Z�b�:���q�ݶ����E�[�]���št��j�B;���!LK=hĖ�T��:�qY�S#�����Z޼���ՂY��bpCYd�ݥ��;�֩v���)�V���#��t��Wu֨f[�mv�ݵ�_W<t�@����q���,��
;��窎���}-ve��UcS��xiU�֒�2�ͽޛ)����M^�yӉMY8�D=�3�����N���;k�Ӽ�ކ~�]Ϟʌs��1��e�P��Ï��]�2�\c��yGy�ތvÐ�fq�E^���D�Dz#۷*{��םr�l)Y��\���9k���?g�X�ns�Yg4����s���w;.>���Z��|�Z��I������E�r�����!�-6mX�?�7mk��g�u�:�^��1��M���X9li�N�8E]z���2�Ťe6k����gY��n�� �;~v�����h��m�WV˼cgv�ՠ)Ϙ?��hp���Z*�Cgޢ �f% �z��p��{ao:��x���s�%do�;�b����`�~�`u��r	��n���Ǎ�>F��F��v�e�
�F�g���^����Z�A�x-�{�Wt�j�u�mj�Zk)���竲i��N�^,ϝm���˴^WX���+�d]+Hx=�6z��0�������|��v/a2߸�+�y6+��]����ߣ��r�wY�ӃX�]�_7 �d��w{t�:)wz�������lѫq֊�kZ7l�L�%��?sP��/R����q�	q�nG���gίO�rբ��&��?�:�{ɻ�Фi���m�7�s��wJ��C�sH�_V+/<�2�)����<�xV�[���7|M=�=�W��������~*&T��^���\q��/n�\�x'Sյn� ݍ���Ǥu0'YQ;��u��^Ѡ�|NU�k1gZ�O-3��*1��n�cm�e+᧔w� �*�w^Z<U���2��Mv��!�z:�ш��=���%���L��@�<�+�nwq���
���y0,��lӸ��{9����=�A�K,�Y�ښ��w�7��5�,߻��n�)T_�|)�6фw<��+g���=�*�f`����mt��3�]j�=��p�>�Qas�3���P��B����9O/J��q�m���溆JKV���dY�����fߞ#�QU���}G�H{YXπ`�P�a0�����o �v�0���"5@y�������%��ߋu��@�$z_�wQ橓]�bp�7��Ig�:Bkkx�2��e�
���]�v�ά�F%�f�Rw���2�� ��/��{zk�x��C�"�o��5�,�u�w0I�V܎�����F��<Ğ[��̘ޚ<�ޑ'����t�^	f�֔ŋY�������[;��9�D�^_T�O�|�We��9vzX8��t��NW��Jջ��h�w��E*���?�,Z�w,Z}���+5��Õgg3\��.�ΨȖ����oF#�:?!_�a�\�Cs"��:g��B�����E�ǈ� ����wn�;��1�<��@�w�Պ����7gI7P?����ZQR3zeƸ�/����g-V�gf�	�=L��[G���y]j�F$���#���+�*����|S6/w�L��H�`�5�+{;��UΦ�9Ã�8����u�m-z�6)��uw�/���{�S	5죮W�ְI��3}xEm�{=���i�:�C½Bħ�d>��}�{͛��2���]m�>��NW�zoެ�����d)���g�+��~�A�����wٙ��0CG=�ѥtj�K����J�=�����*�l�	L��(�§k�Ys�#{[��m�[��޴���^'G
�lcQ�!�$)Y��3Z��o���*�X��RL�L�����Ŝ,V��;|��'0II��f7���S�h/L\o��/۶4<��T��cc������yY���4v��j�_�Srp�R�S��a�*ŕ~Lwg�a�Y���?x��e_�Mgw=��x��\�$�S��y�ʬ�YW�p4x��ׅn�i�>���k��ӹ{�ƫw]�Gy
=p�(y���l;��"u?
���b ;tT�'���3Rn�&'�H=�t�,{�D��V��'	����u�m���.MN��(ŏ���紝h�r`����c6��{:�m���]EY�P���ݝd��x%|������H�}&YC��/�f]�K�*ʝ<����+��lo���»��#�����=��bz�W�ȶjJ���D)Y��F��`� ��'�'���u�0KT��^c�A�O�v�q5�l�`�0�Ѕm
�>-��y�����/��3�1n(�b�5v�8:�����ǲ���5��jݝįސ���� ��VK�&c=~�:��k0<��Ep�������=ԫ]gP�Z
o����/_sB�ܽ�	g�9:>*�}�:����ʽ�c��o�6�"�}��}�Z:6��HѾ�2<���t�%;�%�*��,N�{�nN���ǹ��߭y�&(3�/$��o�����$+G_w-��z+ޔ�]��q:����b'�K�7^D�Org��gZy<�4�xt&n�=��]�W7�y�)o�-�����43�rN=ό��\��J�d�*k���6�7�3ʘ���:΃4SZ�)�y�=�6r��x���1�`�����M��h�/�;zn�<Y��s��_:��<�ݏ��Ok�i��ņ-� ���E�X�D��m�ٖƞ��WO�"�Z���[�gZ�L��;%���[7�����*���ų�]��F���P��PLC��GE�A�sY�������j��� �**҆f�KQn�#��v-A@�U\�뮮��9u@a�3ƺ�1\��°{K�Q�->�����S�.^D7G��3s^�y��U�}1Y��=f�5uk�6�Y���s;]pЩi�����N=m'y';އ�K��N���ch�烛|�+ζ�\>��e��Ǥ�Ӝ%���qڈ�N��f�6C�<׬Sĕ)#����y���\�����������ڋ�w�۵�[�t��;I���~���Z�1^Wn3�sRtj��G�E�p�U�5/��������|��^Q�o5��G
ǝ�+pE��2v������x���y���i��.�Q�dE�^���)lY�ޝ3��V�.�-���m��4��`����+011�R�#�ZQ(v�V��۰W�)�C��5�K�W��yh���IȨ��`�U9G�:����]�;,�盄�g�S��~e�y��,/}yǦDm�b�7yfJѱ�����}�7�_v�w���
�-�JZ���Å��qߏgF8�RX�zT3
k�We���;�S�x{�N� Z�H�����j�YK�mE�kEwC``��㽱�gb=�7`��2Yoe�!�s/��V�e�D���0`�K�B+s6�D���F����W�6�榢,'�򙁚ٚ�%��[c��Z���A��sr׌p���3���^�� �r(hV��:�~����L���^g��"CAT<{z[q��<���u_����^`c�S2�l�d;g��>L�٦�<�f*��o�)Q��
������M��fWA�)��M�/�*C��l���짼��E�ŗ����\;��dZ0> ���ݷ�X���M�v��4�s��e�p}���gP�00W\8,=�l���U�-�m,��T��
���,W�WJ��EӘOj����+kQ*�Y�?��_W=ok��j^���ի�b�n����tow�-��sX5	����ug�o�ҋ#ܫ�wyAE؍��9��(gf U�;L3q�����?�9<�זW�s���^\��QW��g��J�؞z/*H���P����m=g�	��`{���Ш�λ�g�-�c�=�9x��J�z��Gtv�{�f[�9@�w݇��Ao���[S����A��u��t���`.Բ
K�I�3��;�s.gYٸ$G�7�SV��A��5���������c�]O��hnP��n�u/Z���;9G�;9 xƱ'@�Js���e3#���m�d2�H�D���e�P�M��E�AW�+��'^�c�����쓳cܵ�¡�3C��|���|;���^� �2wO��]
~:�s<���֎T�$WP��oX�����[�R��3�ݙ���\�Az��<�)V�R����m�c3�820ݧaa�|6��w� ��ڛ�}y^&k'
���
<��n\<o�K�.�U��bk���DW�/"V��y1�f�dYƨ����,qF�j���i����qX�/�!�0��>7�GUE��Vj��lݞ����Z5�4�u	�vt����ը���]�,���%�g�S���߽�������b\�:�7��i7�s���PȼL��UyO�����Q�{��ީ�&���ͳ�D���C�p^mI��"���H����w����ә�dΕ��'u�fY�n�z�32J�4��R[˒��f�K�
"��pfTku�YW�lql�޳�e1t��`xG�T����WC�k7�_���^�ʍ�Dozp`�*y0c}�E�c3{�����Ʈ��4s��-��W��􏍓�V���R�R����}�61]��(����m���0�s/%X�l�Hf,XyMzlS��T����������,.�a��2�-�� V��ǵf�f
�\in'c����q��y���%��ͮ˧����\øe+Ε��>�W�c���YD�����!{�
Ы~S�N=��/���V��t�D�`�����/���"��S PQ�
�~\��i�*ʸ=��W'�{�L���`L��8�����+��Dt�'����{T�SVQ��d�O���olNs�`�΁����0zZ��Z��n�xCW�����˅X��i(+=pə�j}yZA�Хp݃�%�����˫Z���o��VB��ՇW;���=��E/V7C�zA�.��vk�S\�PR�9��-Ry��\�����P�c�Vk�:ۚ�C���}�ֲ�u�^3w��V�5��B�{1���>�zoՔ�'�TӀ��[�~ci^�ri�s���f&�Gۜ{hyS���/�!vC��-�O��挋A�ݡ���‽� �����q������	�+���-]���U�O���U�,.'Gt��+�v��Ŭ�Ye�����K�(qc��y�g�J!N�jc��/}���`�[����J\�5S��T�����e�G�rԖJD;��t�w����*��N����.���Y7NTs�gA[��ֻ�*WqifF9�D�@�(��@���F%Y�0s����u�E��2��`�1��G+9���C��%��O8 ލr����;�.���W0�՘;NY���^ՅAp�.X���[�g��&χ<����>|�ᘷ��`�RJ�0��es�+C�^���S���R��6*��4��dR���MΝ�y�j�>U&��u�.��z�Í\"�͘$X�<5��w�6��>��z�H�84�_R`@��f7�z�����CE_����W��ю�b��=
�]g]C2���J�}��?��/z��-z���}�^�,��{V�h���v&C�tz���'�=��z5�l-s�u��wL�t�X\ r�҆��)T�j��������e\[��^J��ic��ð�	������G���o��]�KOp����Q�"7s��d��P��)�X,�s����b&J��g�{�:�e���k|)Y�M?_�j�fDTS.n�^��[؍�����T\�J�hp>k��\�]wM`���ٵ����bѷʱ�T_�}�� �RW<h��ko.��T�U�D�]#Zi���;����������7 ��1�n_S�Eչ��=R�e����K}��wQ�]�;��C����[���-� ��gM</`R�	kZ�5mp�bZ�1��9\�.����P;��i�F�qY���))wb�nI��כ\_v��ØT$m�#�9����'+��l9�N�a'3�օq'��K��|�3B�76&����]�Z��࿘�ܶ��s�R�M�&O���q��Tg~�hA�]�}��E�W�%q�c���>d�tw���Wv����.^�<:?^׳%��~�u�|DZx�^�듇t|������(�.�Bq1<<��G ����#�]%��Lܤ{��/3y�VN��7��vu��}��R��i%�������x��s�G��t��ݧ�iǑ��������S1:M}����۫��$0��e��bI�X�X}�y�ݴ�F����=���w�5c�ܔv\��Gko�����=�p/#������^��3�p�~lz��W�q���E�tv7M���u�/���i���L��S$X���H�`��(�}��-z���5��M,o}p!��]��t 	�e��םK�k�j���뒍��"�
�_����N�y����$��T@��������s�$-np���-+y���#`9F���TCjX�n��9X�ae�.�H�H��m�F���*�r��ƚ�=���+]m뾾Re����]xm�EfL�sFm9|��Nī�19v��u�"�{6p�I]E]��x�//-t�S��qr���C!-�uǝ���=h�#Sj��jS��oF㋖͡�a�D�O=V���-��g:�Mu
Գ�+�{�3lj�4��8�6	o
�MCq��w� �v����!�6 .8y;�w�kpW5����l�v�b6�E�u�4:8ѥy�V����";�tj�b�fN�"���=�r2��J+3�O�p�6
وPN�b�ǜ�KyQr���cTN���`����N9�"c�F��c!��ob�v�� el쒇6E84k0�u�j���_u0��:�T����j�ajޜ�n�[|�:�v�D��<�p�5�k2ΉE�܈��z�Pk��ӻ�,Nvo��	�ʚx�@q��JY85D�6��,����'��<��U�-���|p�¶��3x x:ŉlNcB�i�Z�ה��]ã����y��Xm	���ȌP�J�2�ǫY�{��l����כ}":#��!ƶ�D,�0�|S}c#�%�j4|V�ڝ�K$����T�(�7���=�Z���ɩ�2-_nMojR._-D:� 
.��!M�����¦�X��5�r�GZ���d/OJ�&��CFt�Q� ����Wgwve�����4t�yD;sQ�wU�.�:)�m�}@v[��Y�-�	u�
����*�i�p��J�J�ܕ$�IQ�Z��o�&>ݧ��c7mwRG�-t�ɺ�hҳl�K�岧;-H)�\wb����\�n�Z�ʗA��Z���Y��	�K�NG���]������G�p����NśS��ܯ�K+\��l�P�'X)+`�xӬI��u�����m��{/�M�J�p\�=� �P���9 M�h+��JH��`$7��#u���1�E���	�y��O~!���5�S�[V��q����ɻ���b��+�f)�B���Ȳ�)�ɂk�Ƴ���Lp�u����z׺���P���3�'�F��+��.?)�ۆ����3N�l��/Z@��U�&q�z]�B^>Q�N�^�R�:��L�PgA��v�¸u�h��.�O\�$ިy_ 	}y)�O��o<��#�E��2�����X`����>ػkvsT�	�|1,���z�_"N��T��9�Y�70*}��p��ޭ��=�ۘ(�Kd�/����:��M#V�Yv`.��O���wLv\�X�pW����3�����7��L2l�]p&��w�s�/��jug��W� 9HuT�J�bb(t5��WuB�����Hup�wN�Z�í
^Run�K�ճ�k���v�2ُ1�p�{����b�i�"roJ�rd�	(���y`e�t��kAr�"��i�ȅ��l��w.��w��v���N�*.����w$�éG���'\ە��Fn���������:���l"�
i�̙2�j2�����9_�_ w~�A�ӸO�zkI�w]�g\����L3�@�Z`Gּb+�&8���@bg5 ��YDi�DC 3f\�&��&*�&h� F7�i�*��1������d	!$"蒢~P	�c�,�����J_����W��B� ��C1���
"��#� �R��#L����`��@��G��3`u�G�hA0L�H�D���@��N5����}�c�.�F��m��Uպ1DB aF	�!��B m���(��R�N��ȏ�F<~0�/Z��2c�iJ�D	1�垡f��L����JDI��x��hm�_�*9�`$�)h���WsDF���<b�{������� ���c�h���~'�y� M��qa����$�0#����0����k����r�/��x0�cH��䈣�1&H�� � #��D|9�IL�lI�\b߮l�df�b��cǈ�];��">J	�"�����"�@�!A Y/S��qjk�����0>0���`|�2 �LQ�0�F	�U�J <C#��ҠQ ��:�8� �#1c`rPL@Di���I�Y�� �7VzDx�1� ;��߸��9���]���<Y�Hf4�hQ& dB/�ψ��1M�L3�E�W�Yf#�x��,�Q�E/&g�� azZ<@��&;�@��QDGb`E�0�;��}��-�-ݺ��20���֠i~��:E��Đ$LFE�(Ѣ:DYL	Z��'P@f>0�B(��0%&(��,��c�
!��l�3�2�h�2���/s������8����C"({&@�c��G}�r!R�	�-������$ɈD#�j 3di���(�@�H�<�G�3��#�∆Ѝ0��I�$����|~߬>�*s�������1����b��tb<B i/Ø�,�<P�#ڄ��j@�`qC��� >"� "0���j %	�E |`|@�D�#G�=]W�dɺ�<�5��0e^�?����"��^� w�d��H=N]f�=օ��S��6���bouc��\:��ī�:�N���t��F�fS����vZA�[�N����]VW46������@t5��k�Lb�NC�~�R}"�ك��]8;�ܪ�w�u�ݹ��Aꋩ���ІG�B6p�ID�����I =ҫj"���"H�9� �(d � ]�L
0��"�_Ɂ��FLY���F� .65%�}^��������"���Ԡ@$F	�� d1lY��0U=" I����G�E�,��.@�N���x��r��4G�"8�k��,��"<D��Y�F(�Dq�f &�o�f5� H�q�F<D�ss1�� a?1Hx�#t>�,�ڠQc�S�6Da�x���XF��{�L�{���˳Ѥ� �1u��|@� &{���G�Y��>���@D�Y�b4���C0D��1�@���o��0>!�&$�GH�cQ��YdF�p��s�2�[�ݚ��w��#>2@�"Z P	�b���� 	F�q&<D#/�|@$
#ք3�� �E�� Y� #֣H��(��,�%(�F|y�"HҁuSbs�|�/e�d�d�z���.%( �������qd|��I� "��
#��#��
 ||a��"ȓ�㈒�E��@�DG�#�
8b dۓ�.���1�^�]w��.�ןv[����d4b��@Q@ߛJ $ \�$|@�f�@d~7�a�F��8cm@fL>���c� �!�B>0�|`#d_�X�0;�A#% Θ�)�j禧��u��w�{o��0<Y�	ÄY�����u�1�	0�(�	� rRd�"��F��Q�D� x��Pȣ y)0T���� �L��@�#�B
R`x��Y�{e:x��{6w�ޅ�4�"�F#��d���A �T�F��$Y�a�Ў��1��"�Ȉ�/��wK#�P(��3c�0=J>��M��� � ���T�.�E��m�����7���#���Z��}K/Ⳝ}H���rgb@���ޤ4~��`�h���d�UiΩQ�V�����`�_i!bK�ŧ�6*�/�d�q�:�|GC[��N���=}zՄ�cF�T9��N���4#�b�p�l����n3	��tCմ��u�.d�>NU�
���:�Λ��ї}�S�6�����ڑ-�}���Owk�Ca���)m�1q��s�
���*�騀8��C��ލ���׊��z�yv�}9am��V�����4��ۚ��*������y&�U]��܎��BB����՚Ev�U��p��W),�oB�h�c��ë��Ec�JI�ux+��[�*���<���P�i��Ƞ6�ڊ�YM?z��N��]s.�޴D�K�E��#C���"����Md�9V�!���{]�_�P�o[c%�{�^��OC�A��
�y�ޑYX��nu�������I����VoTσS�C~[Ŏ|�ּ�e�R�iͅ1a���Kw[��);��/<�zwo,�^�M�˳I�N���0y��H����I�;'�K�քu`��a��=����ϒ�.�eÏ����h� r�T7����恮G
�]s+�b��WkZi������³��������=���Mp�w��
��yE��\{���Qzgbʞ"�٨��N��%�
ޙ�g�Z��f�������j��o�Wd;�׫kӽ�cǑ�<�3�]���6Lՙv{@Z��l��v����"D��k���n+ý�r�}2��G�w q�-A��J�յ�.%w�b���X�QvwŮ٥c:�=u��|wH�8Vr��}N�m+nH���+B��KΫt���~�v���q��8�#�;.�6,�}Uo���~6�=~�zn٭���s�`Wg���/3M���-�0��Ŵw�� �xX�`5�<�?.bT6��%B�ţ�q�E�/ԧ�x��W��������;��Q1�ܻ�W���I:~�M��~4G�K�V�/
��W��W��%�ܪ��U��ם�i���1�/xDRgy��i���������K��u0xAUc6t�׼bRl�볛�A��gDIg�\T�Q��<�3��-��{�0e,^�g��9�,zf�ev��l}|߲p�d��>pg�c�;DŎ�<�0�>ʖ���4 F� �k:�${=���,:>�`{�Ck�8��Q����o�l]��"ώ���[�E��S4�>��_b$���x���^\��:�DW��t�3S�����j5�{�{.C���bTt�7ރo������+��A.�^>�X;�dz��n��sy�N�Lץ���Q�M�RV�'������S[vo��3o�X���@k�y: x�>Ek��r�f�D���sI���M��sI�-f�P\p�=��gY�(Fء�J�ۨs,
�'W`��F��9u˖sE��t���^��,�S�X���̫ǩ�1��x8S&G�B�E4����Į �����˧���]�/`�ge�"G��|�Q��Lu����+�Z�T�ń�^VoH+�q�أCz>=,���ڎy�V5e�=�Պ �����/<�}J���t_�B>����^�wsc��$�����{-/��:xb��x����-�{�Щ�t���Y���?\��~:�>��^�c����$��ow:h��g_H�.yo�j:��
y\K�B�>Z�*{^zd>ë�� ������_��&����v̯M~Og��Ymq�z�oCc�ׁ=�]V	bG��U���`�M�zRf��'U��w/X�	�^/y5�T��wjXo�nP��Kg��Yj���:|�T�в5k֡�N#�����~Lw�8�\�V᲼��Z���;Џ����;ȋ$�FP�ϐ���I��A�]N01��~C�� YE�'2�9my�M���׮§�w�����5���v��ai�{��ȯe1��R�����|(�T�;(�{�}}�/#�Յ/�l�k� ��b��r���ND]/duƨ��&~F;��^i�:r��<;t�dX]�|ް�9�~mT�f8U	��.��]�����s��167�M:\Yt�VJ�BYN��g-�h��Օm���p[���:��ƯT�#!��(��=��*r�o5u�!/�Z�v�	��q�&�q����#��3�;]��Z"*�_ ���xfr�q�m���y3H�A=�>ѯ^{��3���5^��r()���8�k����������O���$���lo%&�a�k4zZc:�o��&��ޞjqB������B�,xmjKP47�B�
�B@{��'�g��pn���IE$�:����1���-Û}j����os{=��»֐���w��B�_�z�-�.���m�,6�i�>�a}�0߽0%��o}޷�^�h0�تƎ��v�{:��=�/\u;hʐ��q�ڮY�8�n�g½bG�L����혤�v8z�ϑ�>{�+�W�����t;��Ycy*0u_�'�B,fWj�_��*��=��01	�m����L��k�A��xߍ��F	a�l��?[��+�&᝵v� ��Pg^���(���5F ��p�L}�T�6��Ҭ1�{�v��\kב�@�֖]g�y*����NΠ��4����Ƹ�����0yq�F�V�A�s���k��"����^�xL��S��z���8S�C��<�Ƙ-�n
�h�-����ٮ��C�:��`�N�b���u.;&1��3��c#��Xε�%�Q�ǸZW��ms|��ݖޣƓ������Û��D�C\�c���t7�XtΛ���J����_�VW
�{�XA6�����"�9ā[墽+��w��V����P��'>��֬��7�������¯֑%x����wM�[�[S>)���糚.�
�4a��O7ͬ���Bx55[��~"���-�#��rDBkjί/	���l^��`��	Y�뵯���H�q��)U��6��w��l^䀱yF�z�#�M4�z�^P�{��z냆+��M�K����]{
���R�^����{NVC�S�+��d��"��'&5�{�[��/r��N��NP�6�"�<6���U���O���}��Mo/h�LP]�&����i�S��$��1�����DvүK�Q<9���x�g
>��Y{��䧤�_��O
;��"Ʊ�k����6�v�Ay*�U8�=ީ<ԃ��>�WtϷ\2_t�*<K�$#�7��]�5��9��q��^W(}��ǆ�k�b�~���.�[L}�x�=��9ǃ�<������3u;Xp��A�7{6��ag���3'�Cp;W��Ż�[�P˃�M�A��c镭t�=�j�#p-f�fLWVU��Z�Ui(m�m��q���S�����(��y��]�5�Dܫ1�_d._t��7g)���Wq��J	�ŤV�i�d70�Çp귕vm�;�xPrS�<:)[�`��-�KU�cm�_4�wjx��_]!�\��U�z��#����`�̣�*Q+�#�ꩀo�7o��&�.�d�p!���&�z[��p𛫢W�x�������ky#�7̻�C��_�7�����W�97��U����c{ǟ/?��S#E���Ǡ�4�I��d�Kn�����ק�(�sRd���x�Mx�y�:�
/PF�$'�����K2�.���j �ו�S��꣋��lu��f���I{�ꕃ�Æ�*����}<6�s�R.d/V�ϙζ.�{���*{��OӃ�w�ŞY�yA��.�+`+��7 �~T�]˜�L+f��hM�V��y�1�U���o1>�S��u@qn�elG��ל�58g���||3���T5���&�X���9�44T=x������Ԩ����M���w��;�_ �uY���v���D����B|oշA���Oo�n��	�I���$�Tx�=����5�գ[żx׌���8yC��4�>TڼӐ_��N��^����Z�}T!N�`���&0v������� �*�k�Ǩ↡v<6?y̢;].�6S̩xm^�7ѼӴɭQ�n�g�>���&Tp��y���ή5 �lR���)DY@�9���<�J����x�KT�ń1��o��6���v�5�ٵ��J���(��Ļ�l����ʣ�·�H�ھm��d�kwmsk\d���Kʛ����=EP5���#��-0P�Gگ3��bq�d�u�}��S�'�w7����7�c ٪�'�]Cc����\զ��LC������42�,t|�
�?k���q������`z�6ǀ�Pl~o�%���K�l9�z�'����Z��z���>�ߕ�I�7��^�g��C:�G�`�[�i�(=�u�l�F�����n�h�w����<^��w0�U���=�Ԣ���ޒ��<��6��H7��}��OƉ�͖�Qz�/�߇�4|�Ƭ��ؼ1߽7pI8x�tm�~Px�b��G������ɫ&�~"�?e�X�������8ZB��6����F��Jw�������"f��P(QCk^7�ZX�+��ޯ	P&
�g=��\	���b�b�n�:�]��=�2�l�����`�zϷ�3��S�!�3d��4:B��k�����A�����~�M��u��,�b��z�Sw�n1�/֗y1��b��fu�;��-�/��,��Kѡ��7W�Q���v�)�����[��2�Fn���Qu >��maIT�ɛל1gTU̻��l��θ+OP}�Wwݷ�b@��j�K���$���J&&y�ʏ0)U�-<�m�K��ET^se��}��n�t[��o�<��Vp��8����h>���-��Ľ^�E�E��ҷջ����B����q}��x��Pݟ�������:����d�����y����?m�}�\�<��D���C!��8j�������(V�h�d�5ySμܒ���x���b7���������Yzx�>0y�]_��c���p�=�]]K]���9��0k�=�yv�/�hD+Fz����Z{�	�4�|l��b;ޡ�ݷ�g����������}ҝw���xȼ5=���wv�[;煪�jz�����o/.2�!r�Wjm�R��ߏp�S��q�q�֏��
��͝^fy�����i~y��ã����AQv�c�B����[�=k�t/����O��:ޯ!�dK��j�7���sU����C����6��w(����,8-���{�=,])^9����p�!$x˫ɞ�O�����$V��3ӵ-���4`��Q�T��P�Ŗ�H�U�gR�Н�[.��xlu��u|�(�)�=�Z7�"r��7ǜ.ѕf��C�v�ckJip����zqл��uĤ�,�˶�P�N�[�ȉ�t�n�A�!��cuʸ�� �������o�llA���Yl!�.�� FW!�p�xv�������BR��s�a�p���l]D��+�����Q�T�VP�]�n���)3�p)I�ң�S��CW;͝ǳ�S�h��˙�!�l�R������f͍�hXOxH�#�m_U�S�S>舺�W�kd1o+�K9>I�s��S(�3�yGj�C�-���:�nN���E.����&���rs��W7�m].7�ě@p�'�ʫD��z����(E�-V�)�g�3��t6���r�hӭ�.��X9���f6+��o���ܫ�����Q�[@�Hqs�����+9�y[��؉@m�ZKv'l�=��&pl$��{+h+�[�sװ�o���Wo�{	f\,ڡmՎc�5�i	�.�SR�����p̲j�����2����']�n����[W��� 9��35f�� _?�e9��6S�; 1�G��Y+Vt��+���8lK�ăΘr�&�٢�c2�<`���%���*�*d�=Ur8�e(�ε�,̰�p����u�WMR�;+Uw��@���ݚ�!�9'1�ƥ;\@a��L[���8n�w76;vZ���V%��|ؙ����Z��H���s���oK=/�/xP�e���Xve�	Q��77.��Z��r��f�0R��ml�tT��!6���P���Z�8\iΈ��~�2�tv>��FL/Qí�\q36*�fխK]h"�K��o*��a5�
_c�ra��]v�����:<eݬnV*�KJۢ�fΤ]�D�ϘXA��`�2/2�Z�n��V�-���r���7ӵ�u���z=}iVܻ�w��%���+�h����E���8��y� S7YD��bE+@c�ջciC������v8F(�gn�zf�A6<n�(�ُp������	�=[�M*���	�ss8���aעt��m+6tf�ľ)PҮo%Я����3�wk���v����{ZP|�b��K���t�MJۺ����-����5�ժV���uG�И�z��J��ur.�o+Oyr���(	; e�J����~���Ļ'Ĩ��I��^Q|�еv�n�h�/m"�"mt�\�Y�K-sz���Ou�*��	��ڽA�hS���]�������9����Gt\�2D�6�bKo��}`�F��NS!T�nq�N
X�B��]�Ȫ�9!5��iq�\���`�	wv:8�:8��[wD?��h����m�K��B�Ij+c�Z(\��&��d�7�F�o>:�V�l�Okt^+*�v��8�d�N|[�נ5�1x��S����+y�J�M>�`4��],(z�/gsj>ʡ��\���f���҂Wۗ:����#1����Ԛ�M��=oWrކ.��OOڽ|�zn��<�U�g�G�;�~f4�Օ��GhA�ߟ��}e�������=�8w�g���%Տ%v|�y]�6׎�U���o's�������L��5���S����8�+�̪�wi�u��έ���Ky�m�Yq���ډ5j�y�w�(�x宎M��ow�=�v��𗖅c�w���\1)��>>���	�O ���%_]��o�ΫD�.�l̥��Ҁ��v9�c���UXіl�e�qyyu����,���۷��K=�.߯�Q#�s��0��L�qfܺK�ۺ�+̈W�#Zy�CG��3���o�ۼ}/���q��g��A;�xT[��w_��G�_�H�S������L��y�]�kǸ�^�=����<:w��s�I�Ǐ�vI��|���]qڧsu�ʱQ�[�?'�}��vv�P�>~>���j�W��P`���Oy���q�]��C+:���{����D��Ɔ����,�qSGZ'�EI���:9�k�ہ>	�[]X�X���,urr���{WX:�� /�\*q#��ʇ�S�
���]�"	��S!@��4�訇�����u�����U1���D-ʵ:sJ����������1aG��^q�a��\�vN���s\��x��ʂ���U%<�K�;�=Q/c����l׽�:��n�)��!�4.Z��@��ξ�q�i�FI����q���<x��Ip��~N�
��{���_r{:�4=f��f�S�+��z��[u9�d��9��.ў�zaU]�������b�1/-������<R�Ut �g�{A��+�i@�Skr�;k�.%����[�����Iff��������2K�}^��~�+���~�.�ӧWK�W����	��z>�}�2���>��@���s�Ƹ�{��v�+0O��W��l���M�ۦ�����z��|�{�f4�[nz�Rϓ�]1J��r����R��O<wVf	~��<}�\A��A�7�� U��|��]du�Y�w�OJjwl���t.y�-;�9����V����_��_���"C�tvI�i�y���m{l�w�?�Y\mw/��X<�ɋ�����ڽ�zk��CQ���������o����׬o��s�+�kX�����/DC�نoU솩W ����h�it7wK��@lY��
8պ�gZ1M���]f�7n[�ڲ��7��Vf9Þ�Y�N.�_���۲ �Q��wx��fQ�fAIZ�"�W�'r���s鷺����|���
7��R;P6G>4{��F���j��-5��j�*�\�s�{ۧ�|"�qm��nG���mk��v(��?a��k<@�/7�� !&�{�N�]��¤��:IVI�΀\�0~������om��y;u��{�{�����j�
W)+"�׏K6��6=�o+.��[}漼��iR�>%3��[�v�4�{4l]�mtOޘ�8*O�_׋xAȨʤ�ĺT�ֺ�����_*`�U����=�Ћ8�=]C�+���!�w��
�m+�x�]w�*Z'{'���C}�뭸�8(O^�7}�W�u?r��mgg�)'�jwM���_U)=���!�"|��='nrl"�½�,/T�vg�m�v���3�s��/��+��,Q�mޤ���3����f#�~�y��[k�=���j=���^�[�G�'��@�*�=��V�� 8��q�OL
2��fgp�ǿm�:do����n���Q����ls�y�v�R�X֕��В޲���irR��r;z[�l!�p��}YJ�2I���Ud�]�^�FG���v��{�5ֻs�Z$%��w3w��B#W]eP�9o���\�Z�XĤ���)Z�ک��V��׶"8�����70-Mg�L�U��=�5�w���MN����<�ɭ����*�:�0g�p�J��#��j�p��P�$wtF��Ε�%�W��lUA*��h�~PJ�/��*O4���h�ǎ����I��_��;��b_�8�W�>[\�����u~������0:�@��ǫ��S�Ԧ=D���e�ך�����u��Uu�K�</ޏ�:�Wc�<6��Պ��r
(9�8s����� E`N�޲��xfզ �=��~K���S���'~�Ą{FMG�rN��x���2�C·��}�5,<7�7���%���]A�a�ԡz;���SK����ڢ��yj�+�	�H�P应����}�o)��<�z�=�����ݝ��}Xs�@��'{ƽ�2��>�{bV�p8�L-+Îp<����K>�V.z�^S%wˇ�xu�C�ʥη7�q������a�ф����qW_Y��#�M���sm��:�<���G݉�z�s���#��Y�dW���k��G�Z���]���<�q�w�]u=z�J���k.�8_N�.�ةv5��%M5��9�y�J0{��9�.�^I��+m�*GS�^T�g�����J��U��{j�t��ƽ��j�S��IlY��]ĳ��͊i]�5zs�qy�ϒ&+8Y�V��o�^��_���;�c��s8��}��g���ʰ���{���+b	�zgF��lu�����W��g;��ʩ>R�T-���ۮ�����y�P����o1���/��=���\�J��]�LU�[�O}�O�G����
N\޾.��8|6x��N^���{�׼�����͟���c��g�� �m�?3m�ӆ�y��-������^`.�[�Z�
F��7sys5;'��Mz�g����e�V2���~.��>��]�.�L��bܜ1�=�/wO�yYj���ׯ�>���X^?
�1�>��]:��{��ww��.���^*��g�'����>��L��Sp�n����F :������ݞ��=n�а��7���w��-*�0�+�vH�C�,���y1	[�l��|��j���T_{,!k��(����#�K��B������y�;>cއ/�{Uע�&+duJp=�%�������f�PU"Tq������^����}��Ћ�lh����F�#���ޘ��v{M�oD��P�ҧ��ۜ�ޔ/�*���Ǭjw�%ü��a�x����hh�3=:k����,�Coc�;j�Hݛ�ky�F6VS�w(�/{��zg)&U����Yf�?�Lak{�􋽡���ǔ���v�=1#��K�D�e�6���;�ۿ�7+tͯ`����u���I�_�tZa�H�y]r�����`x'_�]p�&|��Р���{�'�N �]>��E�9r������g��~��ܴ��,�ʀ"Z��k�o��G���Nܯa�Ȑx�s��C�m�]�Y���t����K�d�-o�:�{ud�x����^��˼�r�ϰ*�˯r9�������yGTekl�|��,Z���])b�-�:mz_^??x�a��3;������>��7�� ���,wICn�"���Բ]�ޯ(�k6/� �MT��|�]@*s7�S�q�\3�-�N��,W{��Ƚe��j�~�:gw�����6��gW-�&��N��qb�s���g%����>��3@�,_d��W� 2��&�YŽ<��t�}c��W����\�ƺi��[=�eu�O���ޱ�=�/��}j\58�)�W�-��xkƷ;"�ve���΅�v�.�z�;i�U������!l?��H�����V������"^G�_n(e�_w���W��v����R��c^��_��u�}M�W�G�ف�f���8fHX�ѻ�=X$n�kF���Z:�w���T�Z�]�a��_Z�B���fy���Y�h�<�m��&�+������̻��rh���Nekd��S�B�BZ�o�̝�@r���3�"���(�u�;��ʊiվXw:ŕ�g_Ng���clZ@m����y�~�p��ļ��%�?g%�`���|(�eϊXE8��JO<�^�l�l>C�K��vZߔ�\}g�'����p���-����}�nוu�k�{C���\+9=l�W�\c���5�N32g���Ўt��k6y��x}��듼n�z-˷��k�v/��Ze��AF��<����:t���
��+o+v�(*t��2��m�*����*y�)���p{�ea�~�Z�S�ʾ���jX� '�"�b���][
��Sj��S�ά>��I����c:�5Ư1>y�4ǆO����� 
���5(�+���9�.bž~;t�x����������S��t����Kk?c�o�����ԙ�c�!p�^U��K�N�謏V���~{��}�a�Y����)�2D��岝���0w�H�'����_�Û�G�(T��.���W�#��sφ��o^���<�t��o\@��x�:���d�P��z����^H��g�V�n�⩃��2�%&rO�;�jX6��9WZH�i�c��l
7���������Nʈ`�`�,c���w;���	Q�2�9i�GV�EJ�����'�:�M_11�b0����]6����{r�ᦞm��0�T+�}b�����8�E�=[{�:^��𫿳{�Ol�O���
��D�e��:�m,�l�̬~��մ��3-/Tꗕ{vY�^^��羹ݩ<�\��D�C��w�ݾ����c���v�)�ܟ	�C�����S���ַ����5:��_�ǃ>�nz�r#b2W�W��U��=�/��]�r2pP{���I�}��ID�xK�
�<�=���ꮼy���J~�oޒ�R�t���?v,~�K��USC��ݹΑܔ�N��9�%��~� �^{}���v����X�~-Y��+�X��:��o������/%�κ��{0�gi|*3��.k/|󐹑�>�x5T$��M�`��NW����%�yW���/IL�	��wr<�gG{���h�?O>�`���l))�U�֯&]�sV♃�<���Ɠ\|߯�*ǂq�_�E({��n�[��1>֏��=��xa�^�4<|�{l��[|�f�\���]�]K+���jxv+pV�}p�}��o7����y���%.>�D�ܶ�`�C�R��˛X��]�C1u>���W<�uǚq�eK�/쒌Ŗ�e�����4�zY�x3ߝ]�@[��;�<]v��<;^�1��5yӹcyOz���Ub�_Y���vc�1��j�O���4J�#�_T�Qc��ׯְ�d��� ݬ>B��rp�VW]f� V��r��ײr��Y�H�xS�E���,�ɸ��!&�R��t����Z�.c����o��S��	��l��7� v���}��r}jN>2oR��}�__ޠ�k��!j�v2*��<7��C����
Vn����~�7�»{��g�#=�KԳ��а���	i��J��*�@�ȑ��w
^�+k �\:ָ�^�1� /�Ռ�~��Y���
�*Ǯ�����/g��p����u�!�+�|�R�眚�g���WͲ�gZ�]����|��D_�+�&Ҝ�x��W�z��Cv�[n�#�Qy�f�;�|�**��~�V?�2����jG�5�F})vg�(jQ�+��Vwƍ��|�qk�og�,)�[��f���[K���yy(-��zf�+��O���'z�����۪~	�����ry�4����֫©�+�b���;�{E��g{g���bM����r}zs��΅z�v6��7˨��%���{�2�{̫�3=���,+�j-SsN��[���ǃjH�q�B���tU�&1b��]vR��sF�Ł5�5��P]/A%M[�Z��'%oU�Z9�>����N��nшdYW�z���Ps9��s=D�@o-�[���V^�C��
NZ���K�Ƕ���j%L{ڐўx�R��>��pw����ֽ�Uڸ:F�8�huu�I���}�י�P����^Kx�����gw������Wm��O�N��U�ݯ>{S�*6ߧ�/vU�R%�8��*���Q��a	~ʞ���0����Dѥ�<̠����k#�'J=o#����U�r�z/+���B��(`8)������=x�����\h9ki7�;O_/Dr�����<��z��Ze�Ge��E�zGd�Xp�ϋ�g����[�ĥ����Gk}�Y���zl������=�ٹH`��%�f�{7��i�=��7}�W�Ž�� �邹�����]�R�߽�<WO��j>B������|e\�_�ƃݹ_���m
�tL8�˹{Ś}��]<�_�1Ӭ�?C��Ns��/-?a���u���ͥ��'��.���#��{1�vE�}~�ERG4>�C���4c=��V4�3!W{I��ӣ�����+��e���}�פ/"�Φ�a��>��}(���CL� �.��������Ggd�\i�=x�u���J�f����\��G"N��@��J;kF�V#�pR�Wl��z�>�[���Qj*�����$d�$Β�p�ˆ�f�)��l���%M������ӱ�_Q��tI��VǪ�v��9W��N%�d�{�Q���ɉ�+���X�nwv�x�n�b��r���	�8n��(�҆VbPV�Ԭ���ՋVU��e�nd�n�i(�u����t�q��Cf���csb�3(�N�Y��3>�o��mh>=�3X7 �5���J��Q��$v��[�do]õ�î��k��42TE�,β����D�-.F�_u;̓:�Ю�����ձN,nb�WY7�Q�'�X�n�:i��6ݳH�VV0r�(Ә�_7c[d���vm����p����M�R��f��8 ��; ���.��(��lwWM߳�-�B�`ɽ��16h}��/N�?<	�T�om�TKf�{B���%�a��K;8M\Xk��fCe����7}�&���:6Rލ,ɵ��e�.���>r�b#��b�Q���WZNb�QF����n�禬F���w��ΏZ���K1`�w��k��B�j�؍�˲�����n��(1/��)��D�?*��'{�mM�ϻaȖ���ձ+�1�Z�e'}��N�VWq{���9N�6U�槤X�����/��[`��ȩ���vT������zk�"D�S'�d���WeEkf|2l�Bf#�;Ob�<' �!�|+1�F���*���) ���̄���t�a�ܓ���ˠ��:s1m=�[���ޫ�n��2�D]�p
��چ���9��Їݝ�O]�RWN��j�hk齴��܉��e�{�u�wa�5մ`��4�rۖ�����5�ÁNn���݁G��Dkg���S4�v�Ӧ-ȏ;����LҸw_6{�-��R�9��E�"
m_Z�����%��N�!K�3���9�X�iލ��i�՜��Q���h��a��eY�m�DNAՋ�������#]"�1������&��{4�������QoS����m%'q��SȩP�w�;xz�,i�n�� �*��E�{ru�L�{v�Pi�,\b��l,'6%�S��Ee^�9��C��s:����D��: ��ŉ�f����w�����OrӖ(�����e�;�C��EX|o1*H���k��ε��h�e�:=C��趬Z��V�Y���%�X��8͉>F�����n"i�YD��zev?H6�)��sja�b�k@If�ó���p��7W\�b�c؍�2�9p 2:θ�p�P�}��ː8q�.�i`��%�C���z<�eۼ=9ͭWHU������ι�M�E�+{
�LK]�Do��G��Ƅv.��ӽ��dlӰ��뭩
�*��Opa�m�H;�����S��("h��+D1nP�vW>�4��`nWT��.�C9���WL��Nh�����k]��[��;蓝�;eͼ_+:8*�<�싷�YSjZѽ����y�Q�é�������/�����Ml�"��X��2���̙��wX�� �����m=<wЊ�W{}Q��`s��ֽD)�``6�/=�]	���O�&>�s4������}-ws�7^u�wG�~�3���cnIT�"<�W���7ʈF ;�,qI����쵵r"j�}ý�4N[O�����}��ǒ�=���c{��~�~=��{{�;�H8����7U��U2=h��6�7GN���Q��!Y�Ba��;������L�{Y��/v��Vr������5텫�	�=0�.�r�����+�g�����^az�8��x��ͩ����^�����q�Kǳ����ջ��x;|nE�鑳]h����u�{���2JȺ:��j�>̖�/^m�bXe7:'��f�S1�-Y�/_]�(}�,U�a\��U�>����ײ���&�=��rt=���u�)�<}��y�W?`{ٖ���/>�#{���{���]NcP��R�n'���݃y˱�-y��υ{Z���[�g���/�n�OxU�U,�����ޢv�2r�.��g�}����:��ko�������UN��*�}�Ղ�\�\(��Јjt��z�����ۼ�0�΄l����y�r���xZ�V�˜[%%���Xmp��X��Khvٝ����F�ǧ�bh��u%�f��E����v�;���J9�M?<��� ����T+����'NkƏ���E��L�pR��ێ��C�0q�rzD�������x�;]٫7�E�-V�n���w�V�mZ�Ϸ�Ѷ���\uG���/7�xǽ
�jʻ5�����e&uw�'�� ��hm�_J���l����b�785�o3�t���9l+g7Y�Eۖ��zؤb����x�.�i_fzh�ɯ>W�_;9g��O�9|x�9-Ѕg���/��" #�
���͑�I#��� �-fWw�g/נOOI��ۛw�ŏV*�ҼZ�Ա~7n�5�g���uZ��/v��6Hd%�����{j#��߆�s��M��ygm3V*4���G�wf��{�R���x�~�~V?�J��y:��:���&�z�Ƭo)f>�����,W*_{�P��f`�r!Z�*���պɍ�k��8�^����Ww����((OM��s���{����^˶�����;g�[�p���dyk�5��A���0��˝+:�S�ftďHE�u�����kc��"}�+�f�3��;��h�R�����S]�Z�֖@]X�:<��|�	3c��%���B�M+0��B�A�6��^���t�u$ju9sz��CP(�Ї��̰N��L��ݑ�F?|Tҧ~�ծ�9�
x������Z"�a��F;�ڵ:|�l�����xՓ�MuAX'�	N��!�/J�����{��BǞ;w�g�8_���}�Wy���X��3�v�\�yp��W����z�zЯe�w�T/|=�㾩�T�~�M����:o�GT�t[�Kxgiz��z��=�Rj�Yp�t�s����쀾��Y����!˷����M�5}<�ʿ����}B
3k]{�T��gL7��(��,M�{��^�L'.����G}���7�������U�3��U���"WVxX'�u�o��z�F���_�ޓ�$����\����,.�)Y�=��m_d�i�K�=�C�1�sR9eg�zs+n�kϪvֱ�=R��)CˊW���2�	�`�J�p������}�p�꒷��5oy{3��<��v�wΘ�C�����J�\\���Tk��~�}���z��U�@��.��q/(��:���=�^N��:/���z=��7^�;��\���^ׅ��pu,<jh��8`�f�����X��KL�ӡ2�5�kU���9��;�f��T�+�����7��;�$���7tr���:�5[3:+�V����2�{�V�[��r��@`Oy�>�k�N~�ʋ�����O+�a�օ7���\2V�&v.DA&@�r����6��^61�N��k����޷���^��r%*<w�{|N��,K����p���7<w��u�����}(��B}f�>�FQ�Y��0�[�1ݽ�=��i����Y�=�Is��{ޟ[���{���ˎ2)�����>~�&qt�;�Ő͉>�"} W��$�����ۀ\�C�~�"���{O���]f�q��I{�w�e���5�\�>�RG�eͽᗑ��(��k/J�V�O���1os����r;��N�d�N����_�w�����h��,R�'ww83��L�^y�4��i^&�{7�gʤ���oV{�n�X�IO��=يxmw���8$Sm�;bỗ���U�ޛ�w�Y�3��Ry7���c%��U��Y]x����97ײ;k�IV4��6M�Τh|h���aiW�wpY��fq����8x����v=Z�-X���yɵ�v��`�5�ۻ�};S]�͏L�!���}P|�;!V�u�P�}�8��J��;4a� ��^3�,��������2�f����"e�lhْ���`;&�B�Z��&���]yZ�m-J�ܫ���I�|,�Tk�OR�i鯞�t��id��4����)���y�nTy��	*�� 
���bNx`���E�r�OZl���[�=�/Z�GgM�#^��Ȼ�+��^�⭚�,W���.��S��}r:+۸��j
Q.���e*�y}{K� k�o�(G�{���]���b��#�Ļ��Y�zVH�q���}PN��|�q�۱�t�;X�8�����¬z���Ι�����{�;�� �%�U�s3�]5�yL�g��{�!����{�N�����ř��@�w����Ϩ
_3�]BN1�8T�2�=�rJ��H�/1�+ZYR��vz��۽��L7�R��d<羈L�ݮ��~��1���(^uL���Y\���_��`���N���Q1/�g��
��U:�S�[���~>T��O=���Г��ٹJyu������*֦U��[�W�=0����_C���P��{�f���:z�[&y�g�Z����n�9�}�:fUEH�铫���C��I�r=�R�~��p"q&}csu��m,���~ۭ��h�5��"��urX��W�,>{xߢ�;�}DT�,�O��f�p�����v%�:ԣ��շ�ʸ]�@���j�\�u%��=��=�t'ec7ƖG#�C�|A�U����1���	]�W�+_ßs�	%:�Y�k��J�����՘��I}�;�!�j�}�$�}v�Ӿ5w+���<��̭�����o��ط�!dx9�����tYu/v�]����Gf���S���!�nx~��l�����]j�GL�k7xP���:�y��u�H�9�q�#�I��<�)�%�w�{��u�|ώ��K�ֶ���z�������u�zڠCv��ޙ�~�N�Φ����]����?�v%�a��%�w�w�'�Ȭ��L:l����W��B;Xf�~ƻo&�u>�{Y	kr�WϘ��;O�#+��f�gB��ٟ�p�9-�σ+x�f<C����ʛr�1�e@�<�2�t�\�����k���1gTG�'ڧ+���>k4ֈ�l�I�]�0v)Y��KfV_�M�8?e�07ü���>ۣ�}��E'޻'���!�.S}8{u����h[;�ע�oh��������1��ֳ������y�Z>�U�@+��z�1�$���=��T��t�{�7�ؖ>�yzE�?�7�,<{������7ϲo��KCW�ԛ��H��k��Yu��p�j\]9���0���{[.�r0A�0Ú�rP�D��wv�=��K���w�E��;�>+)���PVq:�n���/x���%	�WZ����hMD-]��5�J;���[��j۰�\�E��}�w&�n�K�z/b�*��u���ԍ�J�=�I�����Z)zQ&�8=�,�U�y�b��<W=#��/�U��0;�OfC%���v�-�z���˼Թ��$0p�]����YY�Ns�YK��dE��6����_�(K�O?-{X2���!�_ZUv=K���U���unI���ɫD�g�SQ6�\Z#�$:j�T��7�F�t���uȸ�q�1��+�q]x��Wט�`�GY{�� |Y�U�'7�u����^����}�7U��{&�)r�9�\�z{J��-sy;���5������{[���<�~+�Z�cu��bz��x�^q��S�P[��p���U_��j�J��9O��{J����,_o��-{)앞���Yq���hy�>?Y�Wsb�|ؽEk쯠��|ɣ�s���v�)�g�}��=��Ջ6��f��,��|[���T�o�UF��pf����+�0� B�L1���*=R�F�=�弇:tf;����:�Zf�{�V�ݢr�*9�F��γ])���vp���I���з�j���nw2�sQ��rWG�k{x5ܺժ1]������h΢݊hsu��*Kx�y�/"yJ�tR�Ι�Q�ծO�e<$���wul�?f������&S�������e�}�]M�{{�2�="v]SK�~�.Y�͇Po��l �sY����K>ܠ�P�5�n����1�LU<��+Ua�r������a�e:�̫=���؛�g�\Ё<)��5\�0Y�ڄ�����Ι\&�-qu��Z �C�"a�W��l�=�M�׆}C����1{ѷ�8�}��%�˜q9�h]�p�mS٪��ˉPb���Ý�'�z���+���k�l��V���� ld�C�C}���o[�Tbܳ��*`[\�Yߐ^�q-���'h�����G�� ��m�T\G:��}M�Dg����h��7�%zݣ�B&;�g�8���J�ޜ���,t��+�Q#S����f*���;�ۨ�Z��587yUķf�I��2�Ϣ
x��m�į����ݜ�v�d�������7=�3Xeڊ����l�_b��[=�PnM��ѳ���M<�5�ߕ�U箭��{1*�[�U�����o�#|�˟}.z��Rc������Pu�Dp"f�')�if��\���8�J+ f��V�`Y}�n��T�]�Y¢��"��ij��"+8Ɜ�;,o�a���{�����IqX^Y�yr�)�6ۿ�K��7gy�t�yG26�W���M.�)����
��R��An�tQ�iӻ�G�lû���Ȓ��vh�,a����Ii�QVv�̗���E|�7�=ň1����S�T:�h��*�k��XX�w3L:lr�H����A��,�Ƚ�ў�ɂ'K�9�8��1�u�'׹�'�pf�eֿovy?Y�~4Lžj��;�Y}�WoMDkƍ����*��V��zvf��Y>�y Mnk{3z�.`όM7�qd��/7�z����c�jv�ҍ0�R���d��5�;�'�U}[T�s��z}��`]Nzf�;r���aW�k����Y�4%F\���X���Q�6�Ǽ."b�f��ؓ��3��ڈ�ca�(.R�r��{.�����^�d�j����]�}��z�?[���:����d[蘉P��51�9�wS��^3uUx������c_�1�1��$��;�[�����;�������FNo���;��H�ݑ݇�R-L��t�����u���̱���4m���j6vV�>�Q��N>���sw�_��O\M�+�N�kq�&).�3�7�_gpSNM�fn�������	�~��+{Y��V�0�i��K���A�����!6���>�uT[ɝ܁���u��8�T�O	8��neL+'���̌����:�Ǐ��ӝ��,��ɼv��V�f�e��Gos�p�|�(l�E�-��w�.��0ho����4��if}��r�Sv3\N!}�%*R�(���k���a+���i���Vi�ʳK�~��ݎ}wF��g+��L���i�l=8.��u�$�N������ ��L�f����𴥍�4��ʓ��\�f�Ʊ(:�9nC�ʯ�ҧ���fv�^��u�g=U�H�#)d�rOQ��������w~3�9�gj����~����D{�7�&���0��Ë�O*�C�^�$=ʲ d]�_�pS�|��̱"���x01��Ì�܁&�Vx2�ʺ$Ǹ�QЌRhX���/V�|�9�{��N��,il���E�;S���H���S.��}��qN�����~_xzض�E��_|�۽*C�S���L�<͍��	Ǣ:PG3&6��H��)&}CVX����g��yݱ�WM��V���uu�1a~��8���d�[�9�/e��	ڪ;>�/b����˙��Ev¯ht�E��aצ-{)p�w�oA��ut]Y5;���O��N{��zGD
ʋ�����:���*����~�~�	�>ȫ���X�G����G�6������ѿ\�<.�'���z�䗧I�F��+�������W���f��o�v�
���zlyן�"8�T�l��C	��;�r��B� �:������÷���1�g�b�d,q.y�+6�g)I��\�P�}���[H��)vŢ�/E���1i"�r�\d�gi��݊�.;nE}N��Pbd�����$�yQI>�t)�4�jÕy+6������4�V�Za\w�I��A��1"�Hs<Ɣ7w0�w���Y9՝�2��\�tS��S�w7k���:ճ�J�J
���VSv��ı�q��&�S�mZ���N�䙇R��l�)1`���TV<Z���۫*)F��qf]g6���)��d|�3�<�aC�z�u�KK[G2�1ۀ�15�t�k�w5��F���}���(>@C��ᰲ,u�X�D<�I�g9�0��۹e��|n�[99���;&�����pEH�SlV�/�f,�x(h���E ��Oxmg+�c>`���;DYؔ�����<���l�n�Yj�	u)��-�����{yK�W@�t��6!S73�e\ꡗxy���F����R&q��ܺ%t`\�Rv��n���bSa`�Y�]�I;���(s�ۺ�8q#��P���Gt	+x�K0�����5Ԛ~�R�3}���oK@����FM��\�+]r�pm��h�i�b��{LTM<�2��Z;h��ŇZ�w9��]f�*c�
�\d\��$-���U8�(c�!oqv��K�u�8 f�#��I��z�e��D�NTe��:ָV�Ur�OsU5p��ˤn��u��5@geӫ1ta�X&9����-��we��8>�w"�ݽи��D�H�I[��52��|���@�����V�]Q�X�5�U�x9NT$]jB����O/aƕwB��3�]V��JjtHa�nZ��L�.�Rn�d����oM����8�ڹ���T�B)����/.�CtS�b���+����
� ��pi����:os��G��h��N[z/;v�RJ�u7��E���Y�Ӹ�?Ֆ�/���aȄ0��Bu�#ק�������S���3�g7���PCV�ݔ�M���9�&�^siP�?�6�[x�:����)WW3h�)����slc��]M7܈;�Ջ
�r譥�Qah3,���Wǀk�($�C��j%�q�3_遍��Ȑ{ospՒ��#��Nǘj����Gc�:�e�Rv������E��dJ].���y;��rR�ӟ&Z�렯������5+�t��ؚ��:�}��gP%����L��Չ٩gZJLq���>X1��0��kk�����ز�7S��i���q�*�����ܺu��tD��}h��i]:���w�Q����F@���E҄36j��D���EQ�V�LY)j�"��a��8�� 7���jL��Ь�W�M�M�3�K:[���Uu�1B��z�����l�T��Sz)��^Zs���HDl�����lP�z��� )u �pa�O�n�%���#������x�����`����R�[��b�E�O�-AX���0�
�sed�cm4)�xͶA�\Q⠖��ur�GY�2�T3�t�n������QO���8;^��^�����fٟl��b�C���h���R�z<CU12� '��G�y�/w�x��6x�j�O߮�Rx^�W���dm�^�h ���o����=��Y3~z�;s"z��rX�uS���p��O{�]d-�5-H�iN"g9�g����R�'2�)��ɷ��x����u>tr�N{��GB��++)���SF�K[���3�+���b�}æ%�Qܙ�1��VP��B�-�7���.4'y��d�Q8ì�ʦ�E�~}[����N�:��qz4n�F-����$>�L�[��n��J�e��q��X��ꗺ�s�a�<`�@ӨP��7?b��^N�~�ͼɉ�{Et��
�9���YX;T�oft���J������C-e�i�r�ow9��̼���WoN����)��3~޻+\�ۧ��!-��0���H�+?�,������w@f/I�A�/�Yޡ1K������䕊]ߛ�	Ѫ��W*Q���N���W����z�fϵ迾�a�m����%�7��kW��Wy�Ҍ�{�1��N"\H}OO��*G;Ơ�������<vM�z�+p��˭5��,�͕����k2�H�P\X|]�sds&��ԕ�7k�u�v8Yv8#�&��үZ�1� ���N#�5���3����"�6�nmy���"��(�H:βt�1]&v�^���ds�L@���gP���tѲ���yu��jⰈ�kP$7;4T�z��8��3>�ƙ���7s�6�Lo}�C�>�+]M�hێ޼��]��ư�L7>좠�hQW�872�Hٝ��QX 0Qk���9��']!���\��Һ��k�p^^��ȏ�L�O�2P��3z�F	�87�r]{Yw k��%yG�]ߒ�s6mf����v��3�lt�{���\g *���+�l���μv71�X��D��~��=�Սz�j��s��q�]���q�U.��Z*�L�z�j��=����'p\׶>�S��_�=Y[�7�����b��	�y��r���P��fg���^}J�v������=�m�|�����3bN���ݳ�_h��-J�X�7�C��OK{�j�_�u>q�ҷ�-焻1՚�670zv7�b�̞�����w���GE�A�"l�ܿ`b�<k�����y��9�;�W���S�Զ�636H��K�������tt79��>�Tg��ğdꁼe1:0�990�e���h~�ވ��(��1۽ђ�T�K��v��̚P���=77�USS%�/յl�f����&�̣�����VF�
53�	�¹2����jVt�^S�Xu`��y7፼��p�r����9{O�����\t�ɳ+��Rl������,Ҥ��K�b��MlnJa��^�}{�p����q��ݐk=���T�}Ӟ_l����j�S�;�Ѽ�&73N^G=r�;Y6�>N��>����x��Lu�fy8����<�h�V�
)֢'](��Q�b�_D��t���0�N��%�zQ��#�A�ۑ��o���#	;�����7���\����='*�P�I��{.N�4^��[���=�\ºy�s۽���Y�S�뻐��w�p��;#����0Mduc$��ER��1����߃z榤��Լ����K�ٮr�6��BsƎ��ȫ�h�˩{�����Jh~�[���"|3��!�dx楣����ʺy�ۘj���6�x^F�D�f&���__D�EQ��=N���CQ.��,����tσڞ�ZB��l�s�ߢ�N-�[�B��h�w$܎�g����,3w��}�v}��{��
ឧ�0��N��a�&u�ο=�.�5�]�\9odz��P�e�֮_v��tg���5�,�/��^�
��	���Kδ��2�%z�n\�Fɨ/:u9�-��=���z�)�d)��2�|]��Q.O��+�^�vg������Tsک
{r�(=EB���;u�&柋�ֻ"�.sn�:aQ6,��
�i���3��vu�Ċ�\m�.��m�6��lmp/)7u{��#�@t��1�[c�G�o_M�׽���BoC�XwS2_H85y]`���U��Ƒӛ����6��:��F��MԬ�/�\Μ�1$uR���$Õ5�l�X)T�;-;��W��Ժ�ڋ����O�;2O�ƻP��Sb�:�>����r�X�h6+�����0�����_N�s���`5���~�L�Q]�t��N�����kr�Q�)�W�}��ݒE�c]#,�|��ލռ}�2�޾�7�R�\N��ɪ�]C��>m�$��UF��3�`��Z֣j..\�xW6�n-��s��T<#�#�e1ӊ���_r�GK��®�4�J"kqf,��m�4�ٻ�%ߠ�=&���P�3�T��D��y[�y�r�ym^^up���_�}D]$|�������������k���G�	����|��h�3�W�V�]B���D�PU����~s7e箝��k�*�������L�Sٔ/�y?�9�fi�u-���.�E���6��1Dm0��(��M�����mo�3��d�L�3/���|뇅�kJ�%�^�����치��}n�	�8��`2�O��]˓��\�����(��5P}$��Ψt�爟<�����p�U���aS����Pr1��O��¢4�t���7�J��C�������1�,e�xj��2��#6(�x������y����7�{:.����:��*qL��c��t�D|2����ɬ�m�]�v�0�-��y�ʹ�a=x��kS$��1Q����i�<O�_1�t�V"�}sN������>]���Owz�/�{�w�"�c�-{�w�Rn]��Ǌ�w[�[R��n"��T�퓌F��s^zO/_p��EL��{�������?�j���_8�+�V�\!�﨨�*���M�Z�A�~��"�� }�p�����tU	ɮ����$����O�j��KUS��g^W�vb���F��{S�C���{7���(��y�ސU"���n��K�y�"vkxi���#�-s�[=���<�zl�i�}���r�1z0;���j��;���	V$�H�D�a�b���b��2�ܞ;o�PC"ndk7���3(�S!������n�v���>�Y�����+��S�(�jR�n��Ȇ37{��v��|��&���IB|`+�4�Q��f]B��y9讕�5��������S^{|��뎛�]�xo��i��z��e��B��x�K�aqkgϦ=ն���m��^��7����zf)}~�u�����p�yyoZ@���tf'b�gͿV��8�V�p;��z+���ّM���_z��G�_2~�uԭ��t�.���Uj!;�<�[iL�g���*�_: G{�"�
M�P��[�Ax�u��f��Jݥ%�vӬ�>4r��"���^b���B�vV#��q
�-
�a3�WN40q}Q*�����=����d���B�������Sz�� γ�]��[]�U����3�M�z������d��8�vgg�#�=�!9"|[��lc����]�ꣷ���Y��f��e"pI��ҷ��k��ٛ�C��ƙ�SJ3a[7�u��ވ�#`,�i���Y��-����R'b�.����Dl�.�����t�^[���4(��j�����uZ���on�F��70���p��fnD�m��Z"_���sc.9��+��U���]��'i�>R{�Y,/Ox��x��&c���n�`՝>��NP�|�6NI�����W���cp��0]�Ffҹ��B�K��jYE���g�l7S3[=����'{h��+�~�����<3�,���۰s /"�2@~RuL1z2�.�>8�!˙nfbHwU�jI���"}[��!N�c��"���ݨt�����yN�b�8�x���{o�]�"�U��~�e��Ψ�=z|�-�}� !}+`�=�N��/i���[W��a�tG}�ڊN�;>�k<�x�Vm��ɘ�l�0�x7J�W����糌Є�U��{�hk��Ϡ߻ETb��m`�����������q\w�Wf�a<�^��9�r���Q m�Wp�t�� �Fҧj�Xأ�W[�O�`�z�m"�������]��1ڭl�B3,[�7w�帜Nڦw6��,'�'f����:�Z*����v�4Q�H��2�x�7"�Ͻ�;Ro���|J��jf`	9��-��v�bOU�ί:�7�"R�gڊ�
b�"���f�^.��GMJ�9�cbb�k9`{~��g���e�^�x�<}�g�8���P�)��N���y��6k��\�+M�5�dO7v i�Sp4��MQ24��77f#ą�:7h�~�7������*<�y*��3�r�L��ح�S�u���W���7S:����� _��R�3��1�Cj�;�i�;TL�u�Q�f�de�(;�x�MB/*X�#�)���m�̍ݕIn��u��*7q񑳰��e���܃}���P%󨻟uqs.�7��ON�b1|�xDu�n��Wo�j�4"�y4;��l��Q��������3W�Oo2���UmW[���s��ٔ�n7vo�ܕ���9�ڊ<��8]�m�P�A���׫gyU�n�$�ut`�i�`��h�<��tv��'F23���4�D���"��ގ�ŵ���)�<��N g�<�A;�C��h+��s�|j�Q&��;uj]��g}�}Z3�F�y�YS��O�1����y��c�H��I5���)�m��=6|�w��
����V�{b���)P�{��5o�o/�^�y�����_n� ؇��NLŶ���k���r����Z��kQ�|�g.����eJ�
w�`a��昶�r�(��[y~�u�Lyfɋ]�H�9�"��"8�jD��~�0;�Ύ�����ȅ�,.O{���np�{+�O@ꉒJ*��V�u�����l������2��9����**a�'|!j8��r�(3	u5�)闫"��^�YM:[��2�[������{��:�o�ԃ�{9|"�+��`,Ն�Ȫ��n���{�r�u�C_	N>��U�O�;~��+d"�i�;'c��me�V�,LCJ�ԝڨ�n�a�H:�����csI��q��tc
�K�_z�7�]#c�����A}q�"�H���lTt �q��z2��;��\h�
ޚ�Gn?{���?�n��2?~�Ng�ZuDs>�MF�.�/9�����6#t}�_�/u�o5��e�xs�Z�����	ﱵ�s�����*�o	�����̕1է��F���6��[y�kn�Qq7*k���59:\�B����e����3�o�ɪ��Lݙ�t�I*������^d)}Y>3SCyגs�lz��67a��.�P������(o��V�ǲpxa�h6�G�2��'s�2�uPŇ1��B;='R�|N��a_f ��qƍ�<�D���u���:��]i[�ck;��6l�v��hUt�z���a^�D氳v� �YI'9gGPV��o;�1�+YȈm�.�c͜�:$ڞ�:nձ�`X�i0�dƴ�:n�e�H�.~�W��}�t���O	ۜ����D�����t�LON��=\�T@k�FY��ӜD�,W 5?5鹉꟡���[Y���t����Õ�Rd|��*�;�{��#�����ܝǚ�ʼ�<D^�<�v-�x^������A��{��g���r���n��k�ܭ��uz}h�N��˨��z��/��!v�����L��(����
rf���2�I�����-pk{��$��c��[���<�c7��pgy+q�Ȩ�w=�4r�H,Doh�I
q�*����'ULtSF�1.�.w6�
�yO��ʄ;����n��W��J�F�.�H:d:�e�Ɋf!t�{o�Ѹ�n�����s�	����c�~��-��k]<�,d��)��<��R�J�~��n���sن(��OwuABq���x��}<W��y�m�e�r{����+����<<d��'�+���'7'/��݇W"pl�Ѭ�N»����a�z��$7����h�r<4�_KT����V��)��H�OV4!2+Y��U�*(���*�~��v����&"���^�*8
�5mu�kJD�;�^��(Nѵ�.س|�'nS��Lq��Sq���/���̈́�ogI�@m	�O+�  �-��d9��<�$k (��q��̂u�d��{.����ML�ܯ4G6j�@���c�&��ڈ��ط1~v�@y���Kf'���ѣ���slh1�Ǭ�&IUSJU{%�ˠ�����0�Kca�/�w`�a��KÕ�췫}Ϫ�o���V������@x�oY�P�2fa��Y�o��yn[n�O�f'�P���nwv�}��dtJ0z1�`N��ax��Jѱ�.��'��`��|]k^Iw}j�}����8G�F�6��:�8�ɟ)�
z�N���t���p�v��C:���rƹڸ19�zN�(ys�j�>.��Th�-N��!�H�ۙ�{n� _e>s{I� �N\�g����;n]f��q��Mun�O_no_�F�*�OqNg�S忊��S?���=
�N�wY4U6#����������������۬��!g{�X{���D��	�-�>��OP\~;�1U�s���u�^=��w=��V,���(ã=�V&\R��e� ,�߳M�;|] o����6�T"p�:�z�������r�ך�Q�B�;:���L���Ee<���{] N�p�d�����l�Q��Xʙ�M�'���{:V�u��>���䍐8�{K(��ʘ/&���,p����P�r��d��r��9�b>���y����䃭X]�*v��bX'c&���R#l��1��2.�2������d���2d�έ���6��W����D�J��G������\�b�s�}��=ĦP*���p�ڹ+p��jδ��_Ľ�x�%�.�����(ֵGE�����f�V�����Kf�h�������6-��iJ�zĽ$��g�}���5TT�b�ZI� �c�ܗQ÷Ջ]&���QR�e#��6��ӕ�V�
+����6'Zz�tvq��:���m�/\e*�X��sZ�<V�ʡupVv� v��]@,V� �cm��\���gu�mZ�a�E�@�e=H���"$�v�V~�(!0 u}Za�@�Au/i�Gfe��v�Q˻�r>oK��kC7"B&^ڧ{j
T�1����{��E���[��D�TF�5�8L�q)M�gb�m�nY:[u�m�+�Ry��$9Y�)��䓳 �9C������I-)�-��ӸE�so��W�N��=k.e�{�'趤�l,����7ӓ[k�hL�{KW;op�fr�hً2�ti'G�bu�4]b�N����:-����NU�ٱ��$Sב�T�uX<MN�W¯��������Gۥ/K�K�H�����W���T_�r��fa�g>3x����Iֳ��쐅��d䊠�1H�	��3	Fsm%]\b�!�_�;��;xQn��p�*�����Ҷ���e�:����`DF�r,�V��w}7�B��O�aꑭ�2�m,Un������..��u��N�F6-���֨�2�w���we�Wv�%u:��G�.ΧZ�b�lm�{ݽ}]�C�B;̍m�R/a���~S���U�5B�m�����Z��w2�����h�8d���yP����ʠ�¬��t��Kɲ>A��#�7�����c���fWl��]+�<֕��٫=���-��`���q�	He愭����f~�������n�7H�mV2�O.��:�����d��$Z���8���/��̮n�**	�f�J<�ݗW(��X��z���2�8hߺ��M���|k�DOs�0x]��`���T¤��v�rA��Lۅ`�Wq	�
ͧ0ĂI�ˊ�]�u�]��)��1E˭��}V�md.�dZԼ�'*�:��a͜�M�m$�6(b5ܨ[
���o;��V�]���Z^�uoS�i�t�T��{�z���jԴ�@*�&"�̕w��3q%{�ǲh�>t�r��e�Ώa��e5�t0�\�z.=Vѷ��/��sҔ�Q����3�͋C�Z����s�^�u�<�h5tq�����u6[s�R6������^�.�V��sچ��N
*�2�R��[��>5�IM�(6h���e��eO�L��<�jmu��Ԣ5V�[��{��'�ڹ�k���ː�|����J�����12ܙ�]Э�oP��ؽ�w'Eo�;f��u:j��,�wc�����	�H뵙��񟟒 ��웺��c�l9��uרdtN���n��Ռ���ul���I\�2��_v��A�@_�����H��S�Cܽ�}-Яp��!;e��!.���+:>�z�.z���Q��T����벍�Ş�u�����<)��.��q;s��z�W��jYk"O8U��W�|`x���sݛ,���.�.f�ЬSX��SS+�"���6��#aN���,��|o�4f��{�b��}6�Br�c�����d;��f��]-��Q�d�D���E	�3/�?R���WP�S]�l�����8C��M��ܝ��˴f���Dj5q(�X�_[�^����<x�uy�ǺNo7��O�\{�|8\ь��т�n��wئ���7����j�z+��$���z;�{2(���4�x<�˚I���c�r'�}SIk�c�2"��=����j�Kњ�������_�a�ԀW#O�T��cd���t��\�������VG%L��UZϨ���'"��}��;�u{/�$T{S���v-���w�E�����N�~�u�S~��Aɕ�z�ʀx���E���Y'^h�h�}�&��w	���S(�cAlޣ)��9�x#���
)���v�uc�������A��$�%^e�-4��c*s�T�3�a]ƆuJ�+-��у���1ʐ��Yd���	ڊc�8�㥖��}YI����<�7�=�O�F:����e�-.�
��Ȝq�h߮�Yr��RNU��� "�m����V�I�n�z��4
5KfmDl��We�N��,�匣ᖡ��5�{�17�t��lf����>I��81�";�"�:�*�Hk���F��2�����z֕ɫ��E,��6v�'���#�OV3aQdk���B�:y��g��H\-WTv`̊cƅ:�wFݡmn� L{�}j�e[�ʩd���z�Ɇx*���IN���]Z��ԁ9���ǭ�f�r\��~�SNҭ�=��� !^�b��zU?B�
������fqcz�0j��,��8���nNļ��[��&^#�ɷ쉾j����J�
P�i	�͗��Ї�*�����=�WX��g:)��/�x�u]k�ꉒ��W�!�^��R�0&�m�Qȍ��ʢ{�\;whks�n'ٽ;�c��;S���G��Q��VUB�2ܽ3^���W��c�z��**"�-�c|�JT��ƿoEdq�.%K�!@P]>>���`����n|q*��=y-9��+��j���:/H�Y4���U>��X�bu�.�Yt:92m�鵉,s�`�1ɐh��jg].�V�zٕ�Q�Ec5g�X��䈩��0�J���NV�V �]B��˃s�J�i�P��9ךn�6�\��[��r�F뗂c���]h�4�j�O���Gr��7�87et�z����8]m��{J�k�������CqvXZ3�>�
�"��La�l��2���г�v���@��q׉��q�ш*�BǎP���7�1�BOĀ���>���a6��6kn�9����Ȟ�������mOW��
��xGm�/��	G����[f���$z�%N�H��(\Hg=��X�3zDb��V;1�8�g
����bs'Z�����<���s�U�8�ճd�OF�&�J��ӥ0�ǫ�{��;�g8���z��L���0�&����ʕ�s֙׳���yq��y�S�T��5�S�VQ�R!�=���n�0&8�̻���9����f7܄����꜇��m�R�)�e��G%� E��pщ�	����<��]!�0�z��i��Jz�f�~�a�vsr'��,�'iFfU9�M�_zp�O�j�~Pr^B9T���g��[�ha��f>����n�ܕ�#�݂�76�}
�d�Y��� Yy+��&�I�#�ϱ�S��`�~ȉy]x�Of�ƹ��A\'Qu����AYEQi�Gh�g,m��ƹ���T�.h��h�pd'G�i�F"-aŧ�wZ��=*�&mT����k��t��_0�� Zhud�9�Y�x�0s�mۊ������D��ݟ� vp`{�:v2�fY��L��ZΊU9�@!ǟk��M�*���C��}��J�l�p��������:Uy-w���;qt�W&�3J��Jk�����J���]޳险����{#��b�tnD<�޸Q�e����z�dJ�m�yޜ���������s��<W^��闲�!
�����S\6���s�5�#����CQx+bjV��K�4�k�с�����ݸa���3?�4�&�)ޣِ���YZ�K�ZG��鵢��̓t��ɋ��U�1 W��Q��e�#���u�ww[A�elCi�Z)n�D!ML�p�*����t�Mt�KLחd6hAc�O�"6wed�7��\�9���u)�ϧڙ��q׵31��@-�(��+�f5^^��	��r�+%��<.�ϱ&;�{}�kP<�����Sc>�F���DAx��w����_o]�\vX~��G��n�o�5n�s����r�vu3�z����������3��T=���g��&w~�΋%���R�ÖD�Є;���.ow�u��̊,0�~5Z����5�`P�T�c��c�;�R��8:�;i�o)V_n#\*`;۶�M�S��j�B�A�6�*�����β�0eWQ���Z��̾��/�����-��cQqP�}4�a��'p<YX4
��b�Φ=x�=čm���|���^���ޮ����t�̽`���-���v4%]z���2x��	���k\�0+T&)u�P^����]_>�d�=�X�y�o�wh]��˦Į��uEuM������י~@E.��Vm�]��om��EE�=�~hz�{꿉�l�B��gM�V�87y�S'�7P�(�3��'}~]1n^f^�g!�ʇ��JVyN�=���ʕ:KZ}:o#��	��� oK�תj����zI~5J������hr�t���Sdˆ�7ڪP��]��jC��SB�.�P���6b�G|�J���ѵ�W��gӢm�ϳ�]y��R����'�-{�W{���緱J�wn�7j��w;�f��#�Xk{�"�Mvi�"3�%d^�U�;��>�{՝s��{\�gc�������;W�q�������ϕ,<'f_�y�R�;��	��u�2|g�={;�Γֳ�&Om�f�u��Wwe�eϟ�R�ˡ�%eҕ&(o���*��S�E�m��*�u����ܡ�TV#�.���;���ʒ^w�'�Q��=`�`��˪��&=�:�f�(������ {���?7���З^ �;6�D�g�4sx9(�o9*��d,MF�.���iIB��C�v�"��a�4�c2�I�:Ԛ�?��ˏ��͘�
�I�kF���ePJ��V��V+�i){�t"yB�(�&���W=�*ŭ(�.0ޜ�5m�c1�WV�;��ϼ5XK��?�ދ�ܪ��s�����h!�6��b=W�]�Hl�^c���M�{g!��t�Nj�O��%gG,�Y��N�n;������쯢�J�_w�j)�����M����}~ψz��6��w����]�\�٬��3'2�_��V!�3~��Ug �Fk�T�I}ʾZ���ά�?tO�|_�_E��Eu��w��^�|�Ȏ�����f��͗�]���)Y[���d��O"<�p��0��)r�a�f`\~ID�c�(�6���d����1�;���zڔ7mRI��ֆ�՜�ᕏ�}��gOi���tZ�jN���"e�=~�qp����-�_yoolb��tld����4�X�9\]"��;��dg�5R��>R�J�n;��Z���?Pλ��ّu_���5�Ι뷙���=}%��K����Q�'3��ĸ�F.��N^w����A��h"s!3j!)�X\�aM������س��ŽzNz#�����#s��W�
"j����M��%z�r�O$:9ҽO*2�Ӳv[eH�>�C.��{=|����!�H䱁��[�}�wS<�E�;���<��z{s$���+#+"�oa}͙jY��4��u�*
����VFX����D��+z��Τ�����v��^�$��f�b�A����h3e;�6�v<7�����'�
%@lC*[Y{�v�`�`-ecߴ*k�U��w�~� ��!���*�&�<�DϦ��B摊�I�#Uhқ|��� n��
m��9)W��UBrCPʙ��%�ϻ;�f�(�܁�8U�֜���xg��N19���ڴ!{W�M���.Vzs;� ��H��景R�v�>�	�yg�9I�ӿh9��u�L�w����j-�)Z��d'N�#Oz����`����A���&��@)tZv��z��O{�5��mz%��(}��nB�gg�k:,U������IXaN`���]%�a�alt�S�[��"�8W)Uu-���K׷��_�YQ-�DV�I��F`}#�k.`�v��9\�m�ٚ�u�)�nvD�jz���ſv{]�������x�N^�O)�qmൊ"�����.z�o=݄���q�C��>�Ӱ4�������O�ʋ���St�j#l$+ʲ���&7*��/�"�m�˗!���G���C�Y'x�����Q
���a��y�s����wpCWXq�����+s�
��c�S����p��Wg�'�>i�R���Y�-fopuW7�����w3o�i�9Ɗ�G9��b;m9��)��;I0r}ϕM]��Rs
��
D�0������ɿy��i8�Vf���X��a黾�Y� 0+�5�R�A�"Z�����2�²�WwFH�ڍ�о���_7�{z~�T�A�b'ؽ���ߥ��v��������&�؃.������N�<U�DB��^�&uo�"�'�U��n�ŕ	.�1�P��2Y�IS�a�^��<�y�F �5c�/$��յշ�5�N��O�ɮ2���?oE�t���nzIX?rX5�%�#�m6�Sߥv"}��z*>�NW9�=�ԋ�%e+�q]��5���&�7E+Udc�*D�I���HG*�/�5��=����YQ���S���D�q�b��E�%=b��8d��p�C�L�={O�%�Շ�J��{��o;;OY��Q�"n��B
kGa�FO:�r��{#"��j���N�܏kV���O���˴�~X��Xѕ���AD��DBP���X~���Þ�\LɆ�t�/D�W3�S��sk߿(Y`.�v��~v�)9�R��������_?4�<=��lg?O��"����;EE�5��{�v�f�l�P��gz���NM;��3{�wU�k��m��p�Oyg����ܧo���d���+kV�'����Ύ��t�D4Xj�9�=3W]�C$'�n�Rj⯻��fR\���x睦rzE��*�V� �ueD�m]�����G�r�o�]+}���}ʞ�.�ʓ-F�30�䱍�.;}�ko��)�ń�K�'����ˠ�ݔT��Ә|�=%ѽ��q��{��&�E�����.���Rw3sL�՜]���BY5����5���M���԰=`H��}���؇��Umg�=du�����ݵy����r�N��s�o6r2F���3B�e%�y��ؼ��o{�GV0���wذ��7�7�{��y�+�p�1#����ٗ�VƳ�r3��f���Q�M�эpl�W_��~��*N�GJy/�/�[���Qnen�Pi�]��Mr�QBe�$�� R��q������Q������wz���OC�٢�;�u�z5��ȅ1� B]�~w�~ p�+���o��Ǣ��P���w}E��l�o.8�^�Vk?�hfWr|5�3�wnf�=D��vc��y�Q�kF�gv�}�����	�o(����V
2�\r��Ӈ��bT��]������S;�`	���싫���+�=�%�fO��axgv�Xg_{���K���|o�$eO����@o��}_ Iڌz׷_ ���a�%�;AK�Q/�j��U2�\M�r��brO?d}��/�="T�]JՁQ(���a�5o{5`A� �u�׾�8�/h�]��V7=W�7 ��Ж����Ez��
A�X[����޽D��4v����M�M��9�f+�E:���7
�).Ʈ��k��|(ֲ:%�1I���vG"���|��3
*�,��U9��v�ެK�{&f�����	2���`��aø�!w�D���ٵ��2�ղ�M���M�^�nT�Z��'�2��ϹTz���R�K����rmc���)���D|�V���bv���7�֡�NOyB�����@ӏy{ ̩�
\�;+a)�+��к�u�#���z�6�y����yvaεv���l2ÜM��3����q6{�z�OExcf�1��v4b��p�6���#=k!ۃQQ’�x�u�Bc��{c�v!�闋x�܏u�.]������>r��=�VQ���븤9��^�/ ���=�ι�:ٯ)r�_#~��+/ �^�,��1�\���};����?s3�����F;���;�Հuz0{��WB��T���DSv�͊����r7BPO���RKн��]���Q5T�P�65��72j8����w��ٹZK�Vd:%�˩oUfڟEX�ߑ�[;:��E]	��/�^�Y ]fo���9^���Pg���(Ӏ�M�O�L���s>b����ՈHg�r}W[�[Ê���	�߂��)R�z�Jާ�MS�S�s����_)C���������p��e�I�7��8��-��Ї�*���ͦ�:^��&.]g?��ܯ��2�GM����c̮.]���O�h�����'/X���h���0����:�����F�"�O��sf�e�%��bM՚��2��E���o<<,n�]Q�`8�����&�`E|���_S���Pm���tTg���^\���m`�w�%���+R�z��^�3�N�[N���2FvM�ô��(>#{f�{x3�m���;㓹�0qT��`����fQ=3��N�yCX���L�,Q���XIη����\�u;��&��Wcr_,N��V��mE���%%���*"�n����B�����6�:�[[�p��F��]GPlv�"aV�iL=��Y���݊��͵�K��Ѝo9<f}�{��:���0�ӹ��gU��JlZx0�\�J��ޱg(:�]�C��3v���z��?4���k2e�C&�6P���7���]�-��ӳ����kA��#P�gL�;�GC���Q���4b�Z�6Ѫ�uͺ�È�eԻD3�X�%�[�`���t�۽a��,*�qSI�$c��No�'��;�>ڀ��]F����Pn��J��*lR 9wN�Ηc��r�W]���|�'x��E���Z3gV�P�r�ADݽ�J����q@1�v�X�NM���~J��n&w0�v�G�q���R�㬘'���6�k��cǆ�<�YYG����@<�)9��1�iqt�8�#"����Y�9���s�����S�_.����m���6$�P#(L����P�7;���Tz�{q6��֘���S��͝���%��`��sD�����*�Q���]��w�ޟཱིk=E�;��B����l�u[�v�ç1}�e�:�8�'s��ݨ���-�ִv����j�)3��gU��N-�i�͕3�X�d�X��	^t���W��p�E�b55Ne���X�n^e=�[A`�bh�4�rd�v����^"�_=���UZ�Oz�o�����ww����*[��=���Jn��Gp,��ȷ]���F�E�#��9���u:��J��#�riLZ��CL^�����kC}���(�����ǻE���̨�F�W�ԥ5��;���6��%��Ի��چ��ػ�ݞ(VP̗���܏�fc�*$�3���	�tF�	���d�m��&�W[�)����kVu�­�S\��{��G�C��HJ )hM�v(M|�ȫ%�:��\ҁ��l�cngn��[�[MaA7F�;m'o���	E]�t^��$����gn;�z���a��R=�w5�ց�e��Ee��]˨�C�b������'d�)ݻ�����$Y�c]�����������̼�۞�y<�ˠ���Y�N�S���ܪuq��ΰGou�N�x��	v	�,59�g�Gd�1�x	�S�����}�w�f�B-���4Z���ݖ�,;�vZ펭��B�Eǰ�]���hø!�;A�6{���N4+��!�gtUL~S�r�DzrS	z5�Dq��Oj�%@P���F�m�7z�A�
	<l|$!5=ٖ��3;�k�C�o)���[E��3�>({������rn���0�f�����ԏI��g����\�o�gl	�n�T T�z��{	w�9ifX��aь$�>O��������ܕ���ga=��!UFS�w��m����^�f��r#ּf��D���:�u̝6k��Jߣ��\>�����̎�*�b1*�~va��o#@l�wbx*�~߬*_�ps�a���ua�G�چ�ee�|�x�Oe�ch�u���n���{ԣ�y���/d��@�;d�[E���l�$�kVGju{9k���%���2#�lq<&B��q���NLH��Ev�iGH��̝^����Lz��y�����@'�j�_�o*���z��ˌͺ��rL�Κ�N�Qnf׺�Ԍ���}:=w+�=�i����`�M(MI�k������D��]���n��.Fb�e�ʼ�o�ע��مI��+ܲZՏ�
y�[�4}U'�.��۾�͍�(����4C�4\���/j�.��ֹ�c�n9�֠{�z'�K�˭�űR�ĩ ��Gs�E����yȤ;w^�JSkv��ۭ���Y����k7@��'kNh����YB�loL�r1كN�zoH��`~O�]��9"se�4q��#�ƥ#��0�F���`q��˿g���
�ҵN������d�TϘ�S�S^�o��QĦ��F��N/�t���G����E�UQkJΞ��=+FE[�GK�o]A�a�WL&D��Z�)\=/���YQ�����4���e<��&{Qn*��ݜ/󻱭y�����q�"��<��½x�2 S^B̺3s�ze_p�}k���%o�;���tR�n��ѝ&�9��u1���7b�o��1rV�Ӫ'e�uW�����]��qy�:���R;e�>� ��hf�n���l�����v����y�SH��53y+Q�R�,.��0ʺ���$��9��/��c�/��5~d�C���,̻�=�;��ʾ���|�x+�6�z���i��}x.����U�������ߜf0
,�מ{�7x�d1�kEE"k�j�b�T���*����W�vJ�q��j(WX�W��%���0�^ 	�K�����5�B`�t��[<z,����F	�}Su�+��߅��nMѣ+'Í�Eۋ��#Z{�CҜfjw�˧���w�@<Oe��hI�+�l{�'���E����cl�o(���]�2�R����c��Ѵ���6o5Q�Ʀean��iv��]VyT��9]�fId@�ū�LG�5�E�����}��s�����f���>�O^J�O����UE��O)�<b�������!U�u�OVo�t3uޑ�>pp�z�t mz��B�MJA�.�������	A��Ҫ2{��o�zח���(\\���䀸鑳�K¡�]A�^�Q�9��ttP�8׏���K���T���Vœt�_�r����"&���|�g�|z臒j�0���g��ʪť0M�38tԲ��r�w�\(f�v�:�Tw��q���x3��C,C=�W�N�f	�����u�
������W��ؾ%^=�n�S�Y���;�S4;�|��@��u?5Y���*1�l�']C�VgL������b���2kG�,��݅Kf��ʟ<sv���8�w]���%4"�*��{���Z�_����$,�WDМ̫�SK��3�e���%���}��P���?^ܱ>�=����/]�Ww��j�A~�ͳQ��u���0*��垜-�q��$��Č�������"�������R��F{A�i%;5�8�
�9tp�[R}�k�{�m}��*.��N��V�9��±���[Zlt�۹��t��qrğmJ��[c�Ͳ^�ru1)���5�kn��x�,�ۦ�u��|���\��m��얍;JQ�N��lvj�h�Vv�%$`
��y\���.��wF�O8q�3�ܠ	�d~o���\̽����R�c�T(W�
|B�����i����k�7�^��>,��7��>�c(,�ڼ�{��<��
���S,7r��wWܪ�ɪ��1+��������	��h�]Z�`',�9�4l��Uq�(��G+ ZK�(���wu� �c"�®��*��b�P��㾭�:/'G�D�wJ������y5�A��t����F	^27�2,H�ĭUD�[�f�\N�[�<5�.�=�-so���ꄡw��\2uTz��ߗ������Fy^X�§��9}�n���Z���|ܝ~����Z~Sn.��w���"�;���$��nx�L_dIA}�{�͆�{d����dp��Jt���%ȷ9`W(E�#P�bB����.��}��]ɩx�	��2�Թ����*���\RF�"����-.!��g ˫��� sTW�3_;wg�e�t��N�V}5qئ\�I�U�UbRc��q���P�r�! ���>]�$�$�zo�s����Ƈ�2�-���1�|u�ݺ����>�X�{QX� ~bǚ�����o��vE�l�,TҬ#��hU�j��>A�s�x�l����>Y	%�ٕ�	��ܺeu�߅�Bl�k��9�ك#}���K\�{m�SBX凝\�T��OV�cy�}p�;]�&�^3�qY'7���$�����q�*F�g>�sG��n^(��H�F�t&��f&i�{�=H�v_���]'�s����} i}}�ꇻ�ĕEf+6cE_UQ��*]��Ą&brЫ�r��w��b�S���ep��nN½��f��!�]�(���X���c�,6�f$�������ϧ�:��5j�R�M)ޯ�Mz8��Ք�vW��"߱?^�����|:������`��cH�o�ب9�'����.�&�on��a.y�\i˂Q|���wR�;��U�/lPt�ߢ�]tn�fcM{7 w�}����&7�L�ze�8�M�V*��L!�r�0��O�b��U�r�Sjj|;@�{�.�#��S��;��ٮ����	�%��HoU��lW�� q�tUs��o��UWv�z)X�.f��9��=��x1b+|�"~��Ѻ�	�h��LW�q)9���e�����f��n�iD��N�dTS��Y�2�"�4*�:�M��w�o����~i�TF+�ȇ�������S}����v����\�|_V�+�.�gG1~}"Fg's�����Vn�o�w���Pf�����0Y[HgᩦB���<FV6s��4
ї\�)gut���K�{}�C�a�Yǻ�L=��;�؝�t��h��։�ԕ�t�2��v���S�m�z���m�ۛ������X��pAu��Y�����U$��q���,�ޓ&&�;*9MK.*K�g]��C�Dc*<����9�U^n|(�;v�|R�};1_,� ��:[4=�7�a6��0|��S��㋎|�E��v]7b��W�"{�ͼp���ӑq6f@�s��¦����/�O�gݩ�����#��$����>�m�M�e�.\F�LDMé�D�6�&ʱa���Y�Wۀ��<�{�u{�q���3\�x��I�:�ӈ�5s1�y��T��Z�~'�\��쇮��W½c|�M˨Ǿ��\<�N���뇳S�������	L�^�t����X��Dƥ�@6�ԁ^���׫U��4Bu�d6:����5�\sA�l#ӗ�|!�\�>��׆���VA�ca��z!O�����;��W�;"�1ׯX�"�SE\K�����u{�+_Qv^^�^U�+�ˠ��t[ �W׋�6�ѿ}�g�:WU�����N��<�+�i�������^�ߢ'�����o��X��օ��{ox�խUQy����-mhʧ#p��n��=H�Y���^���]�EzPV%u��^�V��h�&��VZ��6�h�S�
�]-� O����o�vtX�l������1S�do�n'�6���*���,�2�ehvba�\���r�8�	Z{9`yWֺ`��u��fE�{"��u�K� ��jY9���V�빗՘���0hJ�r�o;���?Cѽ�|��-���c=�ڄ�s"�o7ίM��t�)�1��B�m��6�>|���;]��h1KrwX���ʮ�+�	�z���<M�Xg��T�oe��z#���s5hBem��ej,
E�m^*p����%7���́+�V�uנ�[:��j��WN-W�ǫ�ڌD2%ۙ�QԊ�UУ��񨡰����O��E�+���1�{�.��hU�z��p��<�������~O��Tw�������}���k������vc��J;�#��X�&�����&=	�	P����<��8_x�W��n��U�.���:kj�K�O�a-����^�^���C����hw�V���I����(�֫N�gy�^��W�������z����/ί@A�:��f`/�q��ȃ	و�^��R���U��e�_�'���7�Q�n=I9::�w]t������m2}
��Lx��-��(�J>�,�W능>;�����al�A��}Az�������}�#�kny㼳ʠ�S;�&�zw�uz!a�4���]ƷS�F�����p�s����d��0�Gr>��U-x)�r2k�W��+w"��^]Zct�Xo�'Ϻ�cN�c#�<e�չV�mK�Œ�B����M���J��]'�q�Y�k��0���_g��׺�i�y:�5���^-��ܺ�22լ���v��nh���Zj���K�Q���=t�8�v����"@&寏�y����>��t|1X�8ɘ�����`��Ç2��f�aY" eV79���ѝ_D}��ɪ�����o��ƭ,�W���5��;�$�hJ����챗��Ië��x���iTx,�H����H욼���ENߤLD��e�d)Ь*5�}.=�vn�X��uowYBP�1.�/!/��MD��I���/3����&��'&�]~̉QJ%����\�t���c3y���ܙ;E/z��
pb1��:�����l��p_�F��3B�)=Sf��
���'�%�2�F:�ի��i:�U��ѯ[|��Ԃ}1�?
�cY%
�ɡ�4*�%Kux�����k��`v�
��w.k�U�&���J��M�o�=������C��T2�K��I����&��}��0���{Ł�3�ss������n�*�1�򘋿G�r����_���>ұ����i���'`l/r�_��e�}�5�z����w������I��o���~oV".�x��b�1^����I�Q�-΂��OC�j&�d�b��e'�3Eǹ�:��	X�\�?Z��T�Էt����[����{]J�;�I?��]n���7�,�"���1}�z����W�>e*�e���k5B,�Ĩ�f�%����cˤ��u ��V�W\<�:,��wdh��{��H;���~����
��/�gc�͸RB���OU/\é�?F�`������St�c�ǎ�qշ����mUt���T�������!��럖���^��e��F��W��j�.�!t��Kff��F;��tJ=�FY�O��[w!"���p��S�䟈�ݘ��C�x�������oW���Ez}#[i�w����Q�.�/�䣳)�̇K���h1u���u�T��׈������N��Q�X��'_�{X��B���<kz�m��{=�U��{�9�S��b�wB�iv��7,�6l�Xt!�nќ	����P~O��h�龞�V��#�NSS}wU4�}\�tY` zr�����{4����������/{�̼��@f�4йa�+����>�G]ton]^����(�x#��XA�&�3�~acN��'����-蘻�%Un�^�
���3����'���܊�{��1�}IfTg���/+�>l�q�Ɂ�-��y�:��^׸�w(���9y��2{}G]'f�O�v=�~K��U[�"_7�XI��4�a�)�n�	��X��
�>�������m��i��m`o8�r���Vy:�Dv��ZHQ�2��ق��U�7:��үY�K��s�������ha%����r�I���|{#��xq�����e�".���^��J��3vj�fž�+�����w��y��@�/��+}2�_�v��s^X6�z,��an{ ����6^X�C���=Q-?j�U�����v�=�����(f� MVSڙE8Srh���+�`����y����i�#1�b3�L�2��r���^��1/[��GCW�vnf6m�Js������9��|��y���ZH�!�>����(�h$iu�ޜ�&^;�+�&d�m����_�C��u�p��Í�3�wceNwLE��q����bx�]�>=;� #"6uҕ5��8��,O,�:��{8;�e�E%;���'{������������=�R�E�K[2�!T��H�=aV!�Z������W��}�xݨ� �s4Ӭ>��LŕTw�������1�Oa������{�2�kK��z�.�M�݋�;�؄W��%,V��q��,u'Q�N}S^�04����=����@��am�78���J���46gԌn�{�3�:"r�������\���|����i��=�3����΍�0�Nl����i�G���=�M��v�ʲ�<c�i�~g��E�>���Þz��^�%���_�'�0�]�N�J޿��z���Í�<o�]�W#�x$R���"{������{�ǒ1�B@�j��;c�Q�U��d�׈�����ܮ�vy۬%��Q8F�hTrb#C�I���Z�J�5b�V9����4��� �zrVeͼk�s���.��ï!��7��n��\c��P�w
�5t
s2�,�%u^�HWY���lm+��(^o��%���{��C��	*�0���ۏ2GY�Yɪ4_�mu0z)9��l��8ݔc>|��c%���oV-l��֞�Gd]]��VT�+әR�OI"bxv�8����#c�Ҫ�����f�\�7��l�d�t�:��.��/�<FҚ�����l.�0�k��/C&� ʎ�]����0����ӟ^moL$l�@���'j˸-�5�H����X������m.��ES�ۓ;09��yZ��9q$S7C2�4����D�P��v�jLI�e��.�n���R|�{�
��vi�T��S������ê�|5��s8La�7���P��]������U��l���M��^;gJ3+�Β���.E��Y�rĞ�*pRՒWk��P��}�ʉ�*�us3�i������-D�d�Yt�[�y�Y��I��B�=
��Z-\�/��(L:Z]2vЮ����T�%�ϑ�N�rudV����)h=���أbV�a�R��iξ*�:�U�>�j��r����p,۴���pB��d�
��fj��p���mA�ٱt��� �X�W�٘���βM)����nc�N)�3"[��5�NH���sl[W*oe���\k��8��7�q�2����-E��[� �iG[��@�,T��4-^��3v���f8/�����[�ޥf��Vk� �Afr�ڲTO���Lg;�dt�R�2l �T�
f�WWL�/�<��m���j!�e�2uEPgh�sa�G
�wˑ+nt�z�,Ζ��.j�Ym�i�ǧn<��u�i3/���(;
���eQ��wlfn|���q:�W�����r�b��>��s��F�_*@H��w�@������@3F��p��9Z�X�[u�Ҷ���U����(ẗ��،�[�Z��}[��b��p&w]Jr���:�rS���������ĉ�}W=I<�xl�N���ʳ�\��ys��PV��^ܙ�Z1L��h-ޢMfMl`q��	����Ϋ��qK�\���nb �\2:;�*]�M�j��e�}�N�-���C�l������VQ�{�^VNy}��/U*
�Vrwi�j� szK�ld@��pk��@ib6xFR�]��O�B�	Rgo��k�(��Z7�oY��uw�Z0��jD���T����cP�PJ��u+��K��S�b�|~�HN⾙�.�(�$ʻ��VF���6��ԛ�Y�*^�b@�ĕ��EL�E��,�*߄�-�&�ra��:��61��Op|R�h����A��T4y�n��@�d����u·K�0�(���r�eD�:Pǋqm�']u���V����
v�ɱB�iiӣ�H��uN�F`���.�9�[�Q�ob��G[��s�彬����hW[��/��g>8�4䋿f��z
�J�̏f��V��YA޼�c���r*�]v��믮�޴QP�KQ��|�W�z�f0)�&���Q�\@x���K>��|Y@���ƴ�`Wu*�Տ�d�)��� �ێ>Z�W�n��D����j]F��m��d��q�<F}�7��_ə��kU��������Z��g���&�%�4������9ςY;5&�uv��ޔ�~ܦDϟ�9y0������$g{��~�lr��B{/��u3��~�ֆ�Uy(~�M�������ۖ�$���q3�TJ�:����C3����CcEY�[���*poe�N�~�=;�S���0���Deb.�Q4�]����Mh�XW�<������}����~ۨV��_�Q#�!�M���2�;+�<��䡙�< �!%��-=��Se�1�r�w�X���ac(q����fb+�oN���X!�裮uܱ�~��@� ���\	�^���m���_5�/��6#�kO8'#�5�R߷ox녜>��[ߣ���r�3���$k��q��'b��G��r_�]�c;��U
ϓ���kG!�)j�Yg��}���I���h.l:v"�.q�"#����z��\����C�\|N�,֮�t���_��w�B����U�ɗɨ��wM��_Nz�=����"�ڵ�㏮�[IN�5܈1G��b�ٜ
B�_W��=Ӯ6}��Kb�]����q����^����I�z��]��,d���ө/U���o�:ƫ���9���Ϛ��j��x:}��v6Ιޚ�����lE���C�W9���U�e̐\i���דހ��*�X�B� q�j�79]5�s���87�eᥝ3�Й&���Y��Z%����7u��ɗ�}��YHN���i�F�Kn�2�(�y%�/>��ٴ۪#ݚ���0�>�Ef<�yf��D�Vo�˵I�BGm
��/d�{֦�м+9��xlm-�^���w��,����o�c�t��~Ǭ�ҙ�������k��{���c=s`���� ����F�TK�s��z)��+���v���hd��<b&d���U�x�]��ogv��5��'2�� �����'p�5/�����Y0���Ç�7ހq{Bo�Bt����O����Dމ���6#�F���G����Y�����W����uO�3C*��Tߠ�SU�4<���VN��i����!畼��+������݇5<����2�H9su��"+��U��)��٣��S�4�Q�UbSڶ���w����:�$�AԬ�f6&���pC�ԡ��v*P�!��ZO^>��F�9�t�Q�'j��2��95��z��2� �����\&n�e�Iv�˃g)˟1vg�J΃^wJPL�R�Hͻ/]�&� �g��Q�z��"�0�$w+8�$u���:wNG�h������쎵M��=�����}4�6.�
]�&��E�嗅+��-v(�<Yۖ
�Y�R"C��j)�����Ίx��wn,)�X����X��r�
�f�G��<f`�g\y-a�����;˱�vL�v�v7�Q�K7������$l��6�����TL�Ʋ�7�@�y�oO'ڞN��Rm�^���3���mO1��(�L�F@9⳾2�zV�'g{�C*�W��τkbO�m&��t����1Y*�b��	��9n̎�t����e6{�ӝ�(J�	sۺ���̺��W��MlfUu�n��a��}龠�e����5��.ovf�l� Y��ˉ5E���Ű���}9C��G.��2�L\�"�_��V�k�	"��.����+����ؑsOW8��o���U�]��Ve�T����VAt�j�ϵ�V̬�1UW�|y�-W����lD����[��֋vƮ4b�p�)���3W�~�0Ҕ��/�a����\�U5��N�xT	)"6T�P�7o7�NN&Z�a�Cv��w��zɈr��ia1�������=�.C�~�P�6	sN\;�R��r�oo�Q��[�%@�c ܠ�]H�д5�8�]^����:"�!��9�	�Z�2mt��$3
���P�N�Ό���V�k�F�+��Cֆ7eYʉ���~w���<S����#Ǘ;7�^u���xH�+pVv!�)Պ�j�M��s��B�k�B�Q�z�voR�sӑ�.[6�/�1ٸI��3[�h��w�?�5��b�p4���d���+׺��(���������p��ls�_%�'�_��m_>��PU5�A���z�� 	�랡�iH�ȗ���
�fM��Y���qа� [�JC:^8�U9����o{h��8.�M\�~�R'�H�t9ʋ΍��̀,(�	��{'̘��9�~�4�#�B#蘉5�o��]3�P���64���a�+��\���1��q�� �f���83��}>�b`�>���މu�w�g����Ȱ=���X3p��xDP���썽ڶd ���O�mTh�C雈�%���J/�޹�#o���[����+�ڔ\���C�v0�P2����}h$:���b��$4έ��"(��h��<��{bf�l�U���ٕE�+�k�����s۟�B�T�:�Ǝ�j�&�-��1s2c�6Vo� �^�x�U{o^�|���[��)����}���4%��n�-t�7vx���x���`T侬7.����m_)p|T��ӑ�}z���TT��m�_����:Cv�:)ŕ��^&�'F�у�j2�ۛH��8m[��o2�Z4�� ̖�Z�O��^7�g\��K:6k|oM����I[�!N�g.ݾ)��3-��)V�1#�G����:��G:�%f7٬RN\��Ѓ��啟uu���5L��>oDx��{^>��$�]�:��~c��+���������8⃣B�m�^�>3��2�|vxO%�xD69|�5��ns�m�m�o�Wtt���K,I���=Z�~��GA��Ҕ��^�ܢ~��w�+E���W+�:�ģ�H�����[*�Y�ms
��Yr����;~����<k�^.QJ������s�v59�m	�����N���u�k�\Uz9ܯ�y�p���]���z2�C���u����f�tU<�s�m�ųQ�g ��0S��ƽ��R"�C�/BM�N.�$���mLNt�Uh�Ε�7{����{�NɟUx[��/�{dez�м(nݱ�j�#⥁u��>���*ٷ��R���S�\6�>���^���č����V<횗�ӵKu��@�V�Y��v�03;Uр��'>�~0J�}�=*"��c7������h����Zr������o)�`�@�P=�c�]�]E��w�ʷE��z5������ӭU�
sT���k%5�;�+"���y�CM�N�~,i���ufn��}z�p�.�l?`=A��qw�SWμ��ӰoS2���s�f+�hVǿmt=��o�|��oN��o�q���o!�4�0^Wb��7X�ѭK�+�`h�aVh��6�����z�>ph�G\܏x^���VS]�]ѹ+d�wR�:��­�UX4������Ưks�EZ�s�4N\���/1�������]�0uͻ�$��Z&���tcl��uN�U19YO�HK9���fkd�[3D;.�f�`���0s�Xd�6�L8�G��� ���Uپ���	�q>����.ٝ�1Z�s��7�L�d��]���N�)Gc#�8𝦽�f�^����,���r���9:�D��[�.\����G�0#��f u��=핽I*�����)�r]b�ս�r�Dk��*X�����A���
}q/-��l�X|�'ૅN��dcyr�]�ޠ��d�h�-��Z����ez�`����=A��Iz�>`{~��%��/�t����
��"nVm}��p�=���h��c���ĳ=�7�}���"������ ����3��𮂨7��'�׷�`m��y��5���[�Iي�z�������/B�,
��Pܼ;蝻�OR�o҂*�����!�������_V6��ɟ<94m�&4�t�NY;N��p��:��[}ͳl%~#�M羦g�:�η�y׈QW�!�]X�P�� s����Ү��
���ݾ�.��c������3��Q�"�_��Is��go�}f=��װ�^�d}�s�|W\!j+�~�!fו�i��(��K�~��FlA
,
�[�1�٭B�n�ȕ{�v�u���UM�H^�v�;1V��FIٔ��CKD'��0�B���;I�85e� �l�:�6�"�R9t��2�;ɵ�{�6�t�U�m+�	o)`ھ6����K��t����˳��Jݎ)���S���e�w��p�
�5M����}���e���K��~��0@�DF3�3�f{���74u��~ck�6�ؘ������������+�C:�A�q��\��O/�$K�񮽆e��Xw����SbB!���m�I0��SK�~��k�f=�k��#�r�K�~�כ޼�%W��������𼕖q074\�j�
�к��T�L�ڧ�ځ&�w}�5^rO��X�1t��e���`����>x]B�����V���}��h/u}�|Nӷ���|��kܫ̖����@�ב!xE1�g5�"�^j%�o�5�����4]�g.���l�Jl
�oZ�J>�-w��z�)�����w6����fb�rYq/ݔL��2�@�v��+�}[
>��iwP)}BE��_$)
��t�]]����ŬWu��z�;�}��ax)�ٹ^�3�{~(��?q��o�K�u��|k ���+1������DXȏq�n&��%��2��|?/����t�F�2���2yCb�׹/|�ǟ��N�u���egy'�j�gI�5H0�;�8�Z��*�"����lF�곸o���?�e ���}+^C�{]tg�  x��om�!��,�z��ubT�1(`t�1�� .���y={J�(>������a⢘�r�j�<o,��s�t��Y�{h&\K���:v1��Noό��v)$z��m���VFu�I�tp���X2QZ�3v���$^�@V׺�E��I��Ñ�|�y_F�Nipr�Ni[yV��3�/V����º٫ǧ&/w7_�0�h�"Gs~�����DZ*�'[�l�KW�Lo�g���f�x@Sb&;+�W���a߯z	O��Wws���lwjhp�~t#��Ϫ��t�(��r%M�I�j��5�uَ}�!��v�sw�w�
�%o��[����ꩃ7�ͺU�&2	�3b�t�W�^�C����s��9ɧK�NL���5����Tm�q,)�����/H�l#�q<��k�·$>͏^ϝZ�d�lv�n�s#/�r�B��HOG�eNL����Ѧ��Yx��OC����Q�����5vq��������@˜�����~=
��� �l���嵫�0�/W�d��j��@�=�HS�~�wQ�neC���1؇�3%u���f%��n�؂C4mO��hW�.8�׏˅n�F�Čݾ���b��*b�,�<�{h��V���s����t]w��R�}½l�<�k�Dmo�"�+�O])Q���{�h}����ҁ3�q�<�鬁Nc�O��ڧC�i��4gՈ��ͷ�y�Hnzz����FY�<ܤN��]X��y>[6�*B�5<��e��Kհ��\���-]�E\�����s��	�u�����&��.�p���cYq�`��q#NRS����D���ܣ�f)+I�.��\�x�.��ۛNK*�.+ңb���u$�����wf���6������zP߽̃�b�P����ϲ1S�[���N�[0��<ژ�����U�EK�}�{y�h�Yj:3m�F���c�H�)�:anz&kHV�j��fNM�e��2䆇�X�6�]��9|(�Z~��,f��5>-����Z.��[j��Ar��i�����?�*��{j��d�fS����"1��D��l��9������ӮQsl�����ˤ�C���z2j�!��l1��k��ۦ��k��_OY�n��l4g���������\�L�B�Ü���M���U��²���y:_w�v���g��מ��6�zH�9Hh�����Z�G"�%�6(t��3b>�`��W�$�)n�ٟv���Pupw���_2������_�H��A���\�#/]�=��*k����
���y�_�|�mvuq({����Y�ߜ���G��{]�w�|����,��L��t����YG��뷝�j�KB\5(:��g>�^�������j	��xa����U�\S�࢖����o�{[�D:Y�}TJJnB�S�Lz�V�o��{#6O����b�V��s�}o�:��;��P}������ۻ�&4�/n���ٖ���C����q�q�h�p�2��0�:�������� �i~=Jm�|^��Kl�
�e�����Z���:X��k�Kr��
��{��l�d�e��Q=ϫv�j��SyV��
ǲ�ݛI�Q��MӸ���r��ݜ6-���̡֗v+q��\���|���כ}E�w�um�'��5��Ϝ����k>Ye.�wb:�$���C�4��g�챽Ԅ���
4M��y����\�q펪!�[J�f��MKN{���`����=��f6�>�g���: �y���۝u*�e5�<og^oJ�ܘ�D����ݶ ]d��fb�a:ݫ�Mȝ�>ݷ��0���+q�º��+=�3w�{�|����;IZ��2�JFY��zZBɚ�KD���d;��Ү7�{˺��d}�6�\��ϳ�wDs>��S)n&�lT��O�hTXbt�zg-��M��������j�8�F\�H0�X�f%��Mm9��9��@�%i�`ӟ/8g���A�Q������zTM��|웙K2�雊U����z �o�koׯ�۳};�p	��R�l]ƿ�Z��5��C�3���C1|*}��3֢|���}&RW�P����V�s�{� �Y4l��1Y�8/4��н�*�����w�If��*e���Mߺ(֩��2�|�,
�����1���,-��:�\o\�>�3���7�><�4�oՅeH�]�}F��z3.�;wϻ���p�����b�,(�ˇ���CU9�u�.9=�URuS�\%�3@p~y�w~���N��j�IM9���n��[�vXs*�<kc=��#W�#v��;�ƀ�u����98�EL`<��ޥXu~	%�HuNc�a������6��w����*;v\����T�9;$�(����:&7��/Cm���xSR�>�*�����ׯ��k�L��n�L��h1R^��5>7��=�3T�"͙G�)Q{���م�.�����k;s��4�/I��|�!`CS����J�QK�t��!�k��{��-��t�}\t��B�
L��J/�ӷ\d\aq�ZO_,z�WX�(�c���2�ˎ�V�}Ս�noAX�h��)���U��>�%b,�
��`�9�v:44��ҕ�p޺�fiy�9�Gs�l	�NV�Gf��T�ʂ�V`W��:>�M�i��(�mu>C0Y�\�d,�o\j咓WYFM-��	aXgn�*�FBx��|�����=K�rB�W3������#�;3*:�6�t�NC�ͧ�֤.I4O't\�y��o��'��l���QE���A"��Eƻt�y�/��U�]-�tm�)�T�����^�+e�*/�R�k:\���y���^`��D�l�20��7���V�P�'Dm<te�/�خrp9�����Ga�IAt��n�;^.�Y�c^��u�7&&*J������*J+��e�Q\-�,c�HQe���͆pM���0qJu�X�Wʬ;��腛�@rۏ�g*�[xv�q��u�0�4����G�����<}u��_LVM�r�� ��H��٫u�fN ]���řV�nC�@1��k5M�eR�4�V�Va��&,���<8�N���`�K��̆��[�zA\vC�u<���y0�v�׀RA-�V��c���<�<��16����TТ7�ۘ��R��"h9V�!�f��ʈ9�~���+=���kp����i����a��;<�i�[qV4�Bf4�.�[�>��1\pA��{�h�+\!�����������,��e#K��*�>��ڬU��� �<y�a��/���Z3���P�k����uآ�dJ�]v�ʞ�"��n��i��3�)��r�1bX}��+u���v��j����Eus�{��Ԗ�Yث8��č�ɛ Un�g��H���E���'>��yز ̾�|e���
���CV�
���qH�.�Wcb{�&�ᕷm���=�u^М�&G���
O)�mJ|^�xU��o3��w>��ܧ�`w��x�-�'XG27F����H;�G!��:�P`�e��ME��VM��m��Sʱ��m_�a'1˯h�Ŷ�},=n[3+F��3��Fݗ�����r����ӫyv �[nM���wp����8������bu�����(틅�B/�IV�.X��{��o1繎f.o#Z�B�-4	Y}'uR�o�*S&���rBf=�p��F��gOT�m����x�9Ҝ�o�#֨��w)ַ��b�K��
��H���F��!��������
�r6���[°�Ra���qn���Ӌ��`���]Z�,0�2{�|�2d�G&��)�M��5.���ED=pv�F���i�e����>����;�I!�M�w=5��N/>�c&}�����L���,p(hQ��9���ϓ�ቘɴ$k�j��w��P�Yn��@Rg�jj��e�o�t�m)�|���Q���*����sU=~�7��7�P��q�o�5TC��|��y�-.7K���Ы��?)9��{ٜ6�!�V�V��@�μg�&���hY}e��9��n���r�?��bUu`l"������f��^���?��n�ڪ���?Lz7�^�~���Ѱ��5�Ge
��{ϰm���Co�b�b7lѓHGHz'An�uu!�����us�#ї���/2k�Vyyt��rc�����3R����z2��{�7�B��ND�<׉�V�Uq�8H;ro��"��7��=/^-�T���ʫJ��=^w�@��"?<�{�8��ٳ����}خ}����K�OGyJ�#��Zq�I�K�r��_p��0�#��R��1E淹�y�mOb��c�5�5{]I3:�|o� _��OL�6���@;M�]���� ��e>:�q���t) ږT�������eq��޾�Qے�{S0n�ɮCQ�lNw{5��,�c�v.�7�C�U޻{΢(;��,<��"E�S�qE7*8ed���� ̖u]����wfwu�ZؘF�=���Ё�:
��֒ԑ;~�h駷T�~���)��j�~�ɢ��ǟm��#[*V>�Pˇ�Z�fG���6w=c�L����XYqUK��+7)+u<�$T�ڹ�7��LH������,D�dlK�4���Z��"L��.{�1���S
��T1��#a�^Dx?H������03�Y�����+��>l�]�ӵ�!J�N�@s"�7���E�
�(���m��q4��h���\�^;�O����d��YF+�p�c�x<�Й
S�ƦTå��Xt2��5�L����(��A��~h<E����.&A����ɑ��>Ju՘�д��N��R��w�jw�j�c�%}376�o���KC��K-c�&�(v�&��|]�6ˈ���z9����ޛ�;��h톁�K���X0L���6�Di�g]��RV���i���k����,��ûTC�1�_3x#��^НQk;ޮ�/Ҏ�7g`<�N�Rc+��D��R���҃��VZ�3O\�~^���JET�
�����ӥ�R5��N�W�����[�	��D���Y�9f-��"}wJy�7��Em���'������/nݚ�8��/G-T�]h]��,��4�OUWaX�2�B6��_U�wk]t隻��ѹ�F�E)tƗQ��:�c���;�q�`$
��Bҋ�=��*��OM�c]�&��֬�}΁�}Np4�9'ɝ�;7rjˡ��17k�nU������ڼ+bE3*/K*���ݵ�Y9�E��c{;��;Ѷ���v�d�w��mm�x=f��h�6m��@��\�G_=s��.��7�=�m��rk�9�����־����b�� ]��Us�6,H�y=�]�S�B����'��}����A.{�v�Ɠ��^<��/��<��<f�#-����n��!�f���ɏ}���͕#��D7��Vzǯ���>�S?u���8\��1�络q��䇜��;Ա�<�M?�v�]�*�b��H��F݉��쳳Е�f��G����҆��.��M�;���}�cf$&�Ѿ�#_/#^�m�F���+��xtX�/Vo;��D��Z[���p>�뫌�z=38����)��qATˀ��8_�ښ���4�1fF_'���mx䭕A���c�q��^ɵj��ɬnz8������H�x�~M��R�g��R��)��G�\�c��_'�Kk�B�0�c�7(i�Ӽ,���S�M�S�z���>��������}�]J��J�y���Pg|�n=���pr��zġ��>B�^�t](�3Y��<t��l�������HNHb�Kқ���6x�e�q��Cʏ,ge5�\|Xr���Fǭ?_,�Xׁ��*��W�mm^�R��#B� ��qi��<]]%���z�n��?s5����-��a[�KN�����dT'�WehyB�.ը[��r$:�H-Sy-�olޡV1�dP����P�:���I=<0D��͞�|!8����=��m��1���V�\���;��Lc�"��$��������>���ݶ���Lf
�i�}SR�˛̈4ȇ�B�7���<^t�2��ߍm�\]ߡ.�Aꯛ�=\{�2� :>7�{7��fԊ�Va1C��φyO��͸u���+�M�1�}��ל�ٶ�����)n�冦ƪ	Q��wfw�Խ��f�����}�LV�V+U��}��gr������u�gh�
��y����@�̉���cˠ]{	n����vg&�<�6��;��7�ڞ��x��Z���ͭ�阽�ي�Vc��h|�!�jv��7��6o��K���8 w�����c�3;Υ�;�~��l�#�K���^�S�lK����v�T|����k�̙�E�J�%���.��zg�Ҋ�w�"%��G"v䭗i׏u��3���V^�?m�V9����{�_T������f?���+F���Ì�.x�z)�U�ò֡�tguPRq{k�t�G�}�P��ٛ�N����n|mO70��Y�;w��a'n�����{��5�P���v�}�gp{����K��X��z��<p{g�}�s~��ͭ�\��Xez�о����?�̝����;7�;l�yu��2CY�Ig�pZ��f�� ���Wۋ�������a."���dT��S�y_b�%��!�Ɣo �3�C3��0o�Ӏ�[�w�{���8���n����Ʈk3]fe<��Vn
��Ԣ�p��Bۭ��_�%�"�������������w�u��?��<�>��/�d���Υ8��.����"���e�ȫ��=e���[��`?��:�_���6�N�݃�L��}F~�v��m��
�8��2�Loݷ����:��n��;ٸ�!��%��v�â6g}kG+� �q9/��
卟���zћ�UI5�����}�8�̷mym�J�XG�e�����K�*�ӳ��ɳs�:�C*�w�����Z�Yx�ut9�
S�ʮ�s[6�]���&���j�=�w��gxl��U?b�d�Q�{��iV�z�l�H��{�_^��]U@����a�4�(���w�Q������=/��l<��Q��J������X�����Z�����ON�E,�7���zh���b�������GK�ˇ��U68\�K��=�eRX!��Uξ��U��*�u׏�))�psww�otbT�w�;u��\;��dޯւ@USg*�^ɲa�9^����}I��j�g�
�`��.�	����s�9�Az�=a�.s�FA˖���9����3�1±1v�r<�݀�n��݁(���-��%q��V�y;�ԑ��u�EU���e��4ˑ*�Q~����ɀ��,;��h��MG����!ٚ��ss��� �\�f=��C�8�aD�T�D�u�jR|�v�P�W8� ^�z�c��[�H���{ΙWW�L�]�M3zS�!�p�萼�}L��.J��{�k|5*���8�8U�b�2T�_Q|�0��ڝ�Ga[7[��%>�3��w�{HO�p�O'|���jɩ��GpCa�z�1%�l�9�x��(�@T�XGw��y�W��<g�������<���;�	��&lo�ʦo�����|����n�p>���;Юu�Ӛ.��T��g����.}��� ��$K)������*��x��fk�dĿzD9�ځy�s��Y��DN1�	�塧��9��|C������ޖ}�G�"Wv��)N�.}xo�'������������ʺ�U]3���t(�ǖ�C�:���*�_G���C}��O���p�(�+��.�@���@<�qg�ǣ���^V���ހP��,�\*¿���&)��}ֵ�w�<q�+;/�oB#�h�lE�e��y� ��R�w��~��:�w���e�l��7�ȿtmSC3E׷��|�`�z2�Ȧ����!�/�{���vhZ멕ު�|���I���镟nV�8з�?x˚�oe���Z�"3n��"�5>�o�O�3����j�\��X�f}ή#ڷ�C�u �T�SS|����Wb���FF��I�.�Q���z�%mnxw;�WU�:��=��B�H�9~�9��t�+3�7:o���ȏ���R�{��՝w���oё����V�u���S#(v�*�/q��m;|97�p�T��A��3���ڠnA� �_]��m�<�3��k�Z�PT��]ur��R�[������V��7իu6���Oi�g�k{�3�a[]¶�W<�+h���	]���:�e��l㗓�Q�	!��"�wK=�m��^�i,i��O��ݸ��¿&��qy啣��Cn���3U�]�f�&3r�P��$�P~�V���D�W�F��r�aƏ�Qv�g�j��}����mY0oh��<+27"����{:hv\�f��`��)u�꯶s��w�:T�r϶����0"��=n"�"yb����?"�G�W�շ�����úĝ7�~e�U*�i]�3���	��v/�}�=w�>?�*��]>Ì������R�}z��֪;2������Z៾�>2��u�^%��t�����6�{3}�N��1 ��0�{����X�k��G���y軐V��>B*�\씅���.�9Cz�$9���%�if���z{R�_��Σ�;k�ј���̇���]v s�9݁�˝��R���c=�q��#���7����s�����M����G.{�L�����[���c��..�k4#�W���H2���^��W��޺���y��㝵��a���|ǡ$�W��|�u��9u��F�^��E��r�H��b*fs'��݈b)m���/3Ȩ�2��k��5��#j�`�����W�s��_S~�n�.������\�Ѿ��>�')S� @����@L45�����/O]9�v��pޛ��X�������p�����ʗ����f, �s1�`��5�"w,H����E˾�B�aۧD�!�5SM�T��mG�����I��R��W�7ro����uعX�3ڍ�)��]'��Y�����*p�j�;6\��ֱ/���v�m�v��h�ޭ����?���:������z3�ߓ�Z�_����vs�th��?1�8�s�}��y��︃n�蹼���t��[Q��]D���i�~"�*_[Us�HA@1�Z��z<�-!����=u~�'��B�p�k����\�u����0[9�q�rH�?|}<��}+�L��>���h�� pX� �0�t���s��Ǆ;K5a�e�=>�їu�u�q=�5�Y��^��`���bY��P_��3�Е��'����x��У�`^�s{w��qa�Y¬��ܺ�`M�sE�.���A���*U�W�7������s����d:���>D���=��|t�FSؼǥ�H��d��Ǿ0ze�)�q1�-��Q�癑LP���ej�M����u�Ճ�X�H�'rͫ^76�d��[�S��4�v����M��4�6鵳ݝ�[���\2����yIQ#�=�z>��:��y�T����귟��E
\-���Kj;*��U\k�NEbq~�����d*��v�vk9>�.�z{?Oh/�ui���};���_�p����}�fÉq-`V��=��9w��S��j[�6�-$�n���}��2Y�x5p�x�}�v�}{�7/�w՟^`rQ��� �e���ށz��gr�����c��e����_>0/wT�����k�U3�:c���{��.��Z.鑴>��q&y�u"cj����y��[J6�]����o{X�?Z�+
j��P�y���R�v�4 ��oO�3xGz���������޷]��5��#�C����O���QC��R%�,���L�*��ݷ�9��7���za�7n���5�M��<�^G��2�@}8��7Z��zF��y���q��+��ś���q�J��u|5�kL�E�3]�4�=�r܃}5 3�+��3�yW��\U�
��_V�1�rk�wE�+K��ޯ�2Vwj�!�WK:�.>f@��Ywý�!���wY�Sʢ)l��E�����n�����*�d�Y=���'��<#��U�)�I^^����yfCN�����N�T�����~��}y����"���%3�� �Oՙ�|�p�ԝ��e]hb�ʟ'g�A��ò5L�7�W�����%����Q��{�(+�A@��^�r��۽��l����cc����/﫻 ��Y���3��G��)o�_�`0� �D�����>j+ϳ�l��R���(b�������Y���޷�NFO�rŮ�	�S��LS�:RK�O �~\�����o�!���u{�����na� l�C�*n�xEo�y�It\���rW�H�9��g���T�v[ɖ�қg�_L7�Hg�)�3U������^�� �O����n8玗�fz+�a{��ר;+s��_��s��U]�Qy7w�@+�:fT��/��� 8>��L�-{���Z������/�~�WS�Ê�v�U����^r�t��sG*赌�4`Y9�3���4�^Ұ�&k ��u RǑ,A�l���á��.�*o�[�'eu���1w�7��*^�}\��v�E�����'Gu��g�b�J��^��-W/a�쫵���Ci$Kh�V=��.�[�f������1gcYǽYYQ2�L����Ϸ;?nb3��)}�#=�LC���P�1{N���x ���u�0����om\�Ք��h��C<�tkZ<�l[��n+Y�Y1glt=9�,��3����}8/�zw+plw�`7���+��}���Llp3	��|��)��p�]���y����y�|�h}��
�����k���<����D����7�5+@������̇�"|ږ��Ο��)6g�^x/�M��T;�g��W/}���=����s�ه`�\���~{D�B=]T�f��F�j�D��jb�=s�^@~DF�7���C��eX�����+��rT��
���f_�����ߤ�t&��l�lW����R�&������@������������j�w���}sf8�R����󙅾��ҵu7�vq�v�S5�^� QX`��M+���C���Q�tsw"2���n��AWgb�7&v�=�BoW_N��
�˞�[���W*|0���'*i#9�tb;�L�8od;�._�w�,�������_����m��~��,e�*�=9"da�^ž�:ϑ�;��3� &jY�zop����g{n�E��]S��R����7�rn��z�:��ύϝ�^A�Sf��9�};��xN̟{�Y�{0H7������5����M���M��ժ��>ҵ��N��h�MY��z�Ѷ�H��k9��T�6��*�^-�=57�FO쮕�y�
2�f-H>���]�7�K6�%vY{e�$+��P;�%Et�宵u%�.,���[�;�w�����g9κ�7֞l�ڳ/�F����o��`Z�՘Q�����z�+�W+�w�0f��z�~N�X�7e�S��6n`X��ܧ�p��\Ò�҇N!:��"�]w���v�N�7̹�'�C�5+-���9z%���K�
kp�����x�`����h#���;�+�%o�*.U3�gJ|Ft�uY.V��+4֠�i���g���C��6�:�rؘ[�b�9Q�p˴J�m�x�PK�2��qe0�ǡb�z�J��)lC ����VMi=N�:cS�Gh����c]�/�&>5�e�Ӹ)ka�ZNi��N��.��s�̈́A��ekҷ��Qh���^�uՠ�X�R�����:�Rt#@�����:�5zw������u�^B�Tyټ�3tPrӠ1�|j5��2xB���Nu�uwb��b�tɎ�Ao����Y��oL�U��\WE�\�/:\[mg�t���$�t�]��vP�
��1���+��=�����w�qR�޼]�-��V( v��JAY��.��p!��(�����ś�·Q���;j������G��n��S�5�8m6�ʁ��j�y �}�A�5v��WfR� �	\�'�u6tx7b�X˰�1uoK�֮ǎY�2ģ��r;g���:}�]����d�9��ӻ����_	��y���K'P��>�O!�Մ�v��$�ѱ�;v�ɸé[�HMb����x�45o2Q3h�ibͅ�6���b�j
K��e�ͧヺ�K�5vKP*�LY�t(x����ʼ�E@
�ټ��4�O��N�zw;� �WRZ���aHJ�)K�¢v���|�ʵe�kj�a�t�D�Pr�1,�OL�f^��R�ƾ{L��ܷ�By��>���Vy��4��wN.Y���	�E*4(6�ȕL�D�ذN`f��	\��� �(�/�V|)b�Ӣ��Ô)V�kb���˺GN4p�H���	ɵ���\��Uo�q6�S���|U�X���aTxR�:�v�Q��`���s�yt�W��}N��k�I�f�z_����w��	A1ni�wqG2�QGzV��o�b헓�̾�S�������3�JsweL��-�v|�べB�$pV	9����j���i���:@IKkq�+�܏�9]� �\���'IǠn��>�:��G܃���RY��:b;,�����U���݂OP�'�(1KJ�wⷮCE!�L�9�,�s�C%�}��fo�Í�*<���s�R,8�-��t�g��늸p��L�d�gi'fgJ��]v�-�h�Ue�̵9a���8Mv���3 I�w܎Q��Uk�vJ��+]d6�b"^�ql*�v�>�y��,��?����Ql�F���M]�n��N��=�7��G�&���.�[��ͩ�Lt��Ⓓ�
�S��N�u��\g�O�nw����s:�Ob���K6G"�П1���^�zk̗�:�8'M���/B}���a�-�|}�Y�C���*��#<����]|ä���O�ݱQ�/:���v=���ɿ�.�{��(�p7�MBj��qO �86��vhw	��C%�>�.eT��U3�-��^}S��EM��,��fg���n��{o�J�3�C�wq�7]��}v��k�&~ﱎ��{$�hes>��7�|�X˱6�O��>5��V �Z�D�����]�:m�l��k��=��� Oͫ���&HqJ��69媵�#�~'�Gw�침�jE�߸��k����zn�)�	Rΐt�S"�~��4����S���7�q�_��]��FP������H.��������L]�s೫��C�T�!U��3; �D��e�H���e6��?;3��y������2k���t�.���=�������-�NP?GI�1v��E*
�OU㊊��ԽfiZ�Se�m�`)0�܋�F�4`e��}�8� φNN^c/���Q��ǯ���`/z���!���9{�������k>`\���W��b�ָ����wL*�s6qE�&�}���y}ED2ơlۣ2<�p�ʡ����\<��;;���>��ڑs�;���<1h�(�e��l�Z7�Q!�g)��<��6Z��6������ӈ	m�GU�@��qlա�l���]��[�����ԩ[ۑ4vp��֥��kG8�t�x'�3�_k���2f�u�%�]�+�-c{��S��N�.8 ��7d;[+k�չf���������%g�]|���7��3����*�r��B�)�ɝ�oOi�"1��EQu��?;#�W�(�����|��t�X���a1T�ݜ�+��+��*O�:��y�;�u(ey�#M�MO!�ނD_۴�A����T�gl*nD/h��b��%�' ^ ��[N?dOzg๖C32����Y/��26�V���LjA�S��K�����fe��ܷ,�3����Q�/��H�"q	�:��_���$�J�����ҫw�+ٺ��}$�$�x�t��+����%?7j�;���v �9�Jtqo�֦����úr*^��}P����d�3���֓�KO*���Ϋ��cϜ��>n|-��o���G����ئwt�Et�s�G�3�}�ǵqﾮ(*ݼ�ʹy�Qq�}�N�P��JE��)����1�-����=�Q1��gֹT�S)���~�޽��]0��n_�(�����%��coc��@��!#~�k=�.wQ�ӹ%�����d���=�V�`�_%(ʛ����ʮ�����Û��v�6	�1ȿ����s��2PB����UT�z��*󷼠�Ϫr}H���v�����α]]�Ϋ��N w���7b�4�_@=�u�+;�r�/e�"�An��{���+7� ���k�S�}YL<����R������COK��y$���ګvFgMqL�pU� }:������Ң.�i���F��6�u�St�U������	�'M���l֜T5�=׫ch[ƞ-�/�M���<zfF��ji�mD�����1M]�th�j�7���K������s���v�!#6W����X�>טE��J�T^߫��7c����ı݈yz���L��Pz�oc��&3��W� ��T^���O��ϣ^]���u�7�u���V�^o?6AU�W^�O3��ۆ0�
+¡LE�F�o���/�T~���ԟ�
��z�޹�b�N��r�HZw�s��׹�1����u��^�f}�DHl\���^4���;��"�2����Iw��l��b0ѷvK^؇�6�Bf2���������hw�����,���~�٘��+ص�q�c/�@P7>�J��������說�,0a!�\���|Ĳ([R�|{ޑ��P�|UT�5'��1��c_݃=N=ez��>c�� �n��f`Q���|�`V��\��5$�]|�(yg>9ur��'ć+�U�z��߳�O��ko��e����];�}3g�~w+*���Q�#�f�݊�{ḛ�-����M�xb����@ֱT����f��;y��͜�B��W� �	���S��R��b�䮫�OEk����s�b:���޿G��ɪt�ù��<5[љqC��v�Le�|�]��>h�^�5���5�rp.y�t�(�*��V()���b3n���贫��U�;���lOG�]d����5�ܓ��7�[�vt��V��hm��:�����D<u%�����_[D�����D(5ͼ�;��vmtL�l}Ke�s���u��&@�}���K�v��%v-{��e(u9��%T5�o.5�T6)B)n�ys�{ik�_]v�{��z�Bu�`��q�BS깻k����k_'���N�ַ���3�V�M�\xeb�}��5�9�L\���8�X�C툚|$���.>0�y��¥�^��u�W�\��m��{=I�������@4�V��O�0mj�q���Ȱ�/)�-���
����s��d	N�����W���3�Ǣe�z�2������ކ�V1���kV���tꊧ��$.���'dL��ч.�R3������F%�������� ���}~��~�=�~��]�ԅ�uw��-�_�J풫��M4��Y`;��`��j{7b'�����/k�-3�ETL��)S͋tÏV�\«��ו����_�P���*��/~��ٜӟ:�^JHQ�0�ee����=qÕ��M֝����c-��xo���s�;Xp�Ð�w�r�_yջV��,��I�Y�2��bqSX��Uu�3�A�Z���
=ᾼ�gBw�N��[g��f��~�R�s��~���Tu�����
s]B���-��Y>=��C�zb0��ߕ���;�+��A�>`���|������u:;7䛧?��̥�ǣ��o���,:��y�E�OoY�d��o�Se*�-�C��y�ӕukYpN}�P\,+}ݻ�;���!o��ܡ��D����)�{��1��&j˽��2_����)�Δ����^v�L���ڞ���c�?fX�*}��J_L_9F�}c#�7�wU$f��"�IY��-�5���42���⡭������u���Ek���j�k{A�bN��K��+Ǫ�	(aɘ�\�Tn���p���/�ba��J���[�	;t�B���DT+��E��6����.c|v�o�u�؏9s$_�mɂ�[*������c�"�>�gU���Uz���3a�3�/l+��6a�Vԏ]_J�N���K����������$jv9�f���O������8����Θ�9�0���|��Q�d�W���7Ԉ�8�䦢[�5L�F{ݒ2A%E��}c���~��s�"�Gކp�(��#�yE^��K��gپ�^Rn]����ȡ���;���y�Tt�I]�|���Fc��3C=�"95^Ԯs�� ���#���������ԭ?;�3-yS����M,[�Tv�Ǫ��7�N����EE�+��GI�ѣ�ʕ�s�
�3󩞎�g��_
��x�G
fε7q�ά�^��)e���^��-����ҫ�Fn����AUc������(hڥ3%G9c�
s����f(D��%����هzY�xǮ>�l>��=~ˮ���?7(�Fs�">O���p�D�\K�����2~<��X�g ����)ץs�'-k5v(��#�<�ǐ��g����v�?T��bG.�|{m@e����wf$����?}P+��MXp�^�V�6ϭM},/�����G���u�o~��c���:���o;����q^}��;vy�ѿ�z��X���'�1���^��4������,<���`#��a��!�q6���A�$w�t?$�K�FחO]x�p�2�ƉQq��Jފ>�����>�W_Ddm�셙BW��C}�ǽq��c��4��3�Pb՘3���O1s�x)V-,}ȵ�=��1�Md6��C8���[z|���㕷��_Y��iC��W�!��=ސ�����v[�.}�;j��ކwPYe�V��|m�{������:�qZ�^�7U�k�[Ą��\�u<��Ge\�ި��{����P��;�}��(�ǯ�'Lw#ّ�G�脲ϛV�g�'�|<���4~���Ac�����H�ƽL:�&�=�����t�:�����ﺧ�ӐCY�ђn>�n�g��x�ZJ��*�l^A��4P�*Պ�}Xs���F���=;��� }c�P�Ev@�����<V�7��,̗�i�Ӷ�q�V�c˯ѣ}Π�;h���$����P� �f}�5_Mvn_}��G?4{�VH�E
��!i�pϕ��A�)
���c�h��E�͑�����C�k˅d��O�8M}
����y]�v����Y��p��h��efNN߼k�*L��&ß�o�*�7�0�Iu$
���;Ho���Kӓf��F(�T.DU_�^��6L�E�8�#�ܕζGA̷-� n��'����W�	����H�VE�bR3��Hc�C����M�>��M��yկx�^����ۉ��n�m�����g�u����jפu��)�y���"�(�_��p���O�y��|��2}�U�9?K��y��*j(e<w[�բ�3�/T<��6j	\�M���W�@?u��ևjVT��o�?)��=h�v��	�_]5�k#}�M�Ky�傓��X����!P�:Y��g����wc�bn���f��}>��{bL9lc�}>6A2F,�k⣀�L�o>@��~��5���!b�*��&-g��R��?D_�)Cڇv�{����P��SR '��x�.�}�����Vu���<Qo����xU�\��K*�B:G�+�?Z�)G�-���9�ٌ��&��"X���v��}����q��v��e[�6��۹D��绲��Yj����S�j����6#��+j�:��a�NW�F��`�9Ʈal%XB���P�-����m��C�*����\Tg��m7Ǣ������9���}��x��T;W�
�=�Ny����Z�M�C_/Z�Q����>��y�|�M�Q�����˳p�������ug=v&痾S���k�Q���鿲J�O�8��Q���{��ݔ�}�7{�4��Ǯ�w	�v@��'�@�L����ޜa�%OZ������*�Kr�\D�_'1�Q����4��;����W�/j�@�i�G#��ޑq������b���qQ1��=�DB��}sr�:��ˁ�r����ꩂM틴	�Gޭ#0��ƶ�̐�S/���lǩ��Raȓ���[�ѻQ�q������ٻ�-��X��k2�Iۓ�!��}�������y���6J>"}�S@��	D}L
HV'_52��<��)w��襦���G��7�ϲ>��u�"-B��g7���{�����k�}�9?kv�����Տ�zD��?xңH��5!}�	�:�5Lw�QG�V	Q=�+��P+j�k��n��R���ʘ tS?%�_"�y_��#�VPE�1���B0���s�p=�'�(g�xy��$u��@��q�~ڮ��<^��Vf�
�1�j]\���u�G����8� �92C ��;r��r�$�������	���Dw�𻔦Ů���ia{���f�C�"HDw9�����i�,\���oݔ>ϔQV>�����(�J]�s��>@"��1&���� � O��e3?Y +�pi�1q}f�K&�oʽ�"T��������#�wһ�[�'sw���r f�'��0�HR��j�Y㗶,}�+��-�?:4hz�c�#�|іlWʦ)(��~�� �ѧ��`�J�k�����d�Ι����R1�,�Hcu܀���oD@��ǫ�C{?]h�}���ˠF�Z9%G3[�eNjܩCo��"RVV��b���7�J�B��7i�H7�)0(�/�zs��yg�����*�$l[�y���Y� 0�H�|%�����[+��)�\�o�W��p~���N��ǣ2�����=^m��.����E�͘��*lL��#�^G�Wf2��HbK��D�6<M�񮽮��V�vǜir�\�F�O�sd|W79������#Zُ�M�q![��U��e	!�����~P��0�d�A�������S��9n���o>^�1%<ԇZ�) ���R�nP���-!�
�x�:P�Q���QG.�Ybڊ�-ǩ�#\�ȗ��a�o	d(i�d���&l0�}��C���)��ɺ��VEy��c�"!D���q�����������eV����Q'N��z�@�L��|#a{dT�˴�Fq�2<�r��}L�97+�`}�:��"���� X���ǈ�s��1�n].1^WZ��d��?}s��կ��{亞s�*}�>8��Y�����7��J���.�
��z���a�]
#�}P(�۪��Df")D�	��>�Di�>�.<
߾>U�#,�������E�>NQ�G����Zʞ�X�0u׏C���z��&$���>���<�l�)��@���1Eѓ��@���IT���񦆑���4���f���	ǠJ�/j�ۮ|��mx�F��uPf��z��F�z\���y}����(�i��?: �@s��#i3���(G<~ˁ�Y��T|ZBkf�36�oF}_Q*4�P%�O1�3W;4G�j�޹��y��r����~N`�Κ��w�`]p���h#fǘ�(�'����0�4��=�g�"��9�b�u{�7�a��B��U�q鏾�Q�%Q�m�dI�"���#s����0i5SǍ {�nΠ����] R��W�0#6��b���}���0� }�&
�r�kgtW}*�*]B����<F�~�Uu~4���>{.�l�FF�,�.��Y��W��ȳM������/.�����N��{�j���c�vKGG[[u4�iB�J�Q�qE�V���Ͷ:-��wT9��J�ضs;/i��Q��֫^vE���[�c��C1K�u�O����d� ;�3ʎ IZ��K-�|�.��Q�~X/"�q/��3g�uc����9,}��E�}����v~��U��n��Q$#g�a����lqw6�Ҍi����l3�\���g�~4��s��D�nHg>�>O��z�#掠�����y��⎕�>�x"��E��T@��a�`����$v~��dqxL�#�m��b�ʁ�������jX3��%����ɣ�f��_�k�pkoʆJ�D�T������5��^@n`�%�/��fH� ��3�Y��懵�k鿩|@5b�#��`e�Uf!&�>��k�?�R5�eo����;��cH��gXÄ"41�
��@��=�dx�|E�~���0M�dW�*�䆑��O��68��<��6>��~~��1�D<bn0Q���
]vW�˂�Y���`��\�6Ta:ņ/����
�@'@V/V(��\G�Z���$ $#�ް�bi�@�͌��S��]�����}���Xa}u���+������i8D+p'�2��ه>�	�J�
�8�=�AU`}s�t:�<�=�r�|`���������Չ��I"	�}G�8A+�| p����W>��nbw�^٣���"LQ6�g�b�D#�XDQ��SB%,� L�@I�J*6{�<G�@RH3G�����"(�����De`�]�D|ЛSY�l}�WW�~�9����g{�P5��Ē�L��c�&�� ���g�#�zd}��I �ㄐFK1��#�آHDKI����19,C�n>X�.	�dxr�gʺ{�~y�5�,�=6�t=�c��#gC{���U	(ϐr��@F����%��*�����T2(�2|dĝ��Q����A�#F�����@��|�*�_��h{_ײ���mgj��m����پb�z6�:(�om���e�)G&�N�BKN��v��i�-D8Ⱥ%]�����{��e���뵹�/���t:�]����qkNd�L��kl�z�͝�ޡ]��b�>9��ms�/�eu�kkd�����2/�9:�+u%�B�����'�z��� ��44E&�hY�F��(�\����4�`"�`O�cL�`$|�(�`Ǿb$�.���=(���B	䧐Ǣ${�����w]��=�x��b��]@�"��#]F���|G�
��>�����Dg�U�P!
���Ǳ����#I ���2cLi���J1���$�E���d��V�^��t�'��/���C2w �ˬ@hi,}5"�dl� �׬|l���A �ܑ_(��J'@g���1P��� a�(��=��RD"(��L#��
 ��h�/n�u
���N�}�ʟ��ν?&;������C��*#L��x"F�" Y�;�*WJ�D"*U$� Q�$�Qh�~1�L%�n>^q��D�@�ª�E�����/�f���?hW^�9���on��@Dq�8I�",�0#v���Y���� `�]�(f���dG�sQ� 4�$�䂥�2��#�d��Z��Z�	��c�P˂�L|Di���+���Պ�yM�^\Ŧi��t��]>�dG�1$��,Q�D x���*bL��@e�C� �,��"�Dx�E��
"'��@4
��0� kQ�F@�0(�#��0,��!#֠4�}j @^BN�#\��/�v߲��B�����D5�y� �@�����@ B!�U["���>�D3�C� F�x���d1C1�8`jTcH�"#�f1����1���> i�d��$@&��ͿJ[ﻁ2Ι���~�S�[��R`�Q�����r���R@a!����#_1b,��`
����"Ȅb����(`"�:�C"#�`F���"�Dv 8z�����>1&"H���3��]	?z��O��������� �1��I� 2��=�� a$d@󘏭@Ӧ �F v��dC0Ȉ'�"��\Yb ��)�G�D$� ��>0*�o��M� I��>��@f����U�28�L�}�����m`���� �� �1r�	 .P<@�D �DF�08���	@Y��!%w&hǍ�BȹF}�zd��/M���9�"��Q D��� D����� DD(�"DG�@���� @��@���� @��@���Ȉ"DG��@�""?� D��D@�""D""�D"#�@����@�""?� D���"��� ��@�   D���� DD��
�2�π�p@uZ� ���9 ��>����}�U   p�ݎ� ��W@�  ��
 ӠQ�(  @4:  �� :  :  �V  =th+A��	D��m�B��a��F��6�h4�R k �)Y2-�&CI h 4 
u��� �� �4ΏUy�^�mJo{�R�Q�;��
��:�Y�<�{ޖ��\��
���횪�q:zh����C/xz �R�m�.�[+m�-�� Р fR��U�H�^!�B��y�z #Ҋ$�(�6�R��{�*��*���T(��5�3�
tk���ZQljV帯A��)/;�D�-٪�;bO�K=�v(�+�P�  z�Р���AA� �@d<'E\��D�ܠ=0��ݵ����7��u��n[��ZTs�ǻ�Cl���ݷk7�]v��\w����kmS}�w��m�E� �״

 �l�� k���z;Y� ���:͊��h��wsE`�!�� ��ϰ�$!��������b������\ �<��� ��u��@Q�   k��@� 4�  �� l�Α^����</N���}�}�wwt�5�c�{a�� �N�w��׬M����y6�1���-���cj���{�������Ҡ Q@ Z{�ע������P��z�m�;�<J�G�n�_N�t^n�5B������e������������
 �����*ncvWݗh ��h}   l�  ;�[��a����G��ǣ����ly��P,i���{�l4��!�`yz�ab��;h���8:Up ;��+��y�p��h�yq� 4h �ܻ�PԵ��}�]6ڛ� �vݏg�`�M���>�4����o���n�J��_y�ޕ��m��{�V�[7��[X��Ž�o�|����  2��
    P t��=��y�xAU>�Q}n����AM���cp���ym+�ޞC6<��EUS�7��}�ץ	�>�n����^3݋[e���=��  rV������ݭ��Ӄ� ���B^{ݼ0���{���s��֦�u�t���cx �����m��k��k.Z�Ye�U�� S��LT�@ 4 *~0I)T@   EO�&��R�4`�j��ԁ)U   Ob�H�R�M0CC&�������OS@4x���}�C�'���1x���_�3��w�뜞�o�d�,�x{<���%��33Թ���ř�W����w��w��w���w���{���{��x����݉fb�����$�1ffCř�33�,Ifb����?��hq�Jf�����/�>����|���q���J���
c3�e��yna��m{��^mnw�/Q��Ƹ�ޮu���~�v��ZS��8w��ڇtr�Zs|��B2{��z�gn��=7�k�����y�:���b�)Z�Ib������ g�ن0����N.���7��84��|��{��ƙ����&��s����R�JǪ�ꏲZf��*�"������tcȭ���2��9X$a>&>F�W�0	VEEMd��x/@���g�4�	�_�
�@tV����/֝�%�2�K��� �%Sc�SN��U�R����x��j�-�X�l�R8���8�.���Eؼ>�]b�
�?>�}���G���n�n� W?+;����gJ4�����+���}��k����c�r0R����oi��������J�M���]a��L ��9�.��Ѳ��c�tS�����vB�0懪�,�&����_]ޱ]��(6���W�lH씍ԥ�W���Ҟ����M-L
�0�����ee�Jjon]Y��z49��,[�ہ�8.��{�!�ב�M�'ٹQv��:4�Ւ��o2��b�ȒE̦��Ӆ�tސ���u�֬cR�A��l(,}�廧�V��.��K����b�`�V���h���\�S ����ݾ�"fU�}�i�`1ytvlswmf;�˜8�U�:bVpL�N~��Pu��WK&���|r����m��TՓ�!�h˾� ���w���w��_!h�E��x���ꃦ�;�v
R2�]�xf���"��d�'l�>0��]	���+l��!��v��(�:�;�+���R�B�����d�\��6��\�t'b�k4a�[o��添v����^a���_�*|N��n�.��]�NZ�Z8��bte\C7)')�.y8�Jv�b�nL=��۹cB��n� ��ګ����]�����_P��6��H�y� �����,��7N���n�J(�I����k$�j��-c#T��j���[�Y�.��.�/GIm��۵�v�"XU����
{g��o����cFh�3D���p�o �3���(.��.��:-3�8/E��1�����fzp�ל3�C4L���h����4L��	xg��ZcL� ��Ƹc3���� �.�i�Z`g�i�<3��3L�����{����v!����j2Zx���z�@�A�P}�±\z�H���%�U9�-&%.J���os0�{֦o|�7.��<�6򀼒��v�]s�;o|a�qx��׳���Ӧ��c9�g.f1D�q��`�Bs6D@�HHx�p��)k&�ٮ�r3��6n\'�,�)�����R3B�飫C�S�:�Vܵ]}!�ͦ��9u(�D�ڴJ��ޱǭLο�lD�+���8�/�I͖���*s���y��9-kx�"�*u�����i)�!]l�5z�����	��f� ;5���a\�i$h�7�B&1����{8�;n��]hu�q)��[�[)w:<�''!+�����=�w�����]�f-��s��Rh4]��r-��5[�[�%�>/v��n��Et��ٺ�+z�R�"�D�6�e�̤��U�L���uz�5-��9���Vʚ4�%��
���Že��]���of���L�(X�;�8�{iP)I]��*�Ҁ�6��VL��
�y���k�b��;,���W5���+�kjm�Cg`ذq��pBgf^����&�S�Usnm�y�[b�t ,)F��墎��U�=;�E�OUe��
�T�vԩշ�h�m����T�]���5�:�ˋ4�E��b�h�6��c��Û��x>鯭֫꘡�'tQB�`7E0����Y��C�lљ�����5���U�A���P���ް`�3�+Rڸ8e��[�닾��2n���"pu3+�����t7��{	�ń���f�Ic�s{Q���*��$ޞ�w�����;++\8�e��)��q[(bj$���d�6�m̺���)~n�8�U�n�P,+(\�bQn�N���ꄅs�f�Q{E�g���uyHB��Ot��P���pH��]x�}�&��nB�Ά�-]�v��˙~��k)�ʻ*��.����l=��s�S!�̽W�r���.��C�N�#5Ld��T�r
3;�w9����MޞeQu�t�6�<@/��F����㻣�N�Z�f��Ξ�y��yo<��[��z�Q�(���k9T&P�����ˇ����q�r�n�n���@��4Mcp�������*8��hViQ�oVn��-��MJ��k�]�[���NQ�nh��V��J-�6�[���`X���Kr���6�����'+v������������}�L�������י��u�"lL�(�M`��
67c��^MŸ�iε�qJ%pܒ�ʢ ]I���*Q�I?A�r�#!��E,��Uם�A�ն�=���/������4J�Wv3�kW	��8.��f����n����O��HȲ(��S�5����8?%ʸ5E�٨�����	S��l�;qKyh��uv�f��~I%&�U�v�Λ���{���)�[�Os	���%���7�=��ȎI��P�e~dn%cK����/o�Fe��p�2�����(�^��y��e![l!V�K��+1f�x��j�GBQgf��5]�Dc���(ɢ���70b�g��S��1��w(�P[@ݗS4*����Z�غ���`�rl�4a׶��h"�u4 A���E��١�@�՛m���YY.���&QOf��?���ɻ#G��^D�nI2R�b��D��٘�K�K{�p�����O�ߣ[�j�,�Ut�,��Co�����v9eA���@X:@f�7U��d�[��A��'l�zFXd^�lJ�5u����N�����7H�Q,GEж�`ٻ{�KaQ�	��:�E]�B�N�hf����v�&���s��dt����^i�B�eˉ�h3ի���Z�ͳt�42f�Y��o"�UseGQ��tZE�LIA�
���iJz�ܗ&�9
��đ%�»vȋLR���%D�4�Ck+FT�o3Q5�U�̇6�R��������=A^�E��i�&��K�Řf��K�딚ޖ�n��x(�mAtS��tD�m���w��ݺ�q���+1�֊c6tf:�k-�nMѢ;-�7.Gk"��yr;SX�y{��5([{���k3�0������9Z��y&�o���k[����Ӎ�Z�4��Q5%����7�['ZU˻	4ee���-u% �^�]]J˥�{��s{�98�]�p�q`罂s&���}۷`��wZ�z�G�ԫ�41�2VD��p���iFY7h�]�R��|�BH��e8���[NEg!�C�Z�-���Y�l*Ӻ�otVm0�z�Db$�j�*Ɯ$�	�C-+�dGH�ՋYk2;� O������Qk��2�t?;�j���-zk<4��f�U
͛yg8���ɋ�Q�MRd��j�ci�X���!�[)���B�o4Y�[5��Z0$�Â�sVmZ۽r
�B�W��Y�Z��ͼ�h�J-��w%�̺kk ���WXTɘ�Z�u�L0���,�L&�kq^��Cj���v"�n<E�Sb��N�\Ӻtٌ�r�=�wn�t������6��=�H�8��T���)t�]�f�m~ܕ�b\�'t�h�*��@b���Ԝ寅��PP@z/lg�O�Z����F�ɛv�T
�6�o�Y�o�c=�g!��+dTΈ��N�w�)��~�k~���%����rv��b5gJ�|��UΗg7y��p��k$�ح�Ă��/�]c)^�\���֎����c�QY��ȑ��5v$����6)xDx����F��鱸��l0ӽc%���'�f�%�z�V�uQ����b�mwgw�����t��q�ξ����֨�Ж+7�-�ލ���0d�Q�P�9w�^�B�\�AEiOI�ա �~8
�"!��=v�hXM�n��@��m�r9��p�q���c��פVT%��\�4l�K$
4�-C�7����eOX֗&q_�6jǫB��	����ө�nd�z6����ћ�����茱1u��
�I�del�qL�f�f�NnL�!+�[F����ݫ[�ů��i�vY��O&� 67��b[�ݿ�4+	e�[�M��Xi��^�����K�#���Ȯ��Qi���u�ǲ0qwcڹ.o�.���������x���1���Q�0���d��Yr�P�-�b�q�l:&�� �!�b����*^�fU���j-�+PV&P@�pǋ�R��9VĶ�Gn�jpF��0����B�b[��zV�����S6�Y�I����y�S���FۭJa9��tB�����L���ܷ/�t�r��Z�+v
(�JU�Qʽ�d &��p٩��QP���@�^����Vҩ��p������P�'����!�E-�ę�~�2��w{��.�=�k�sx�P���R,4yѻ:!˼��췗��(V����x���,�朠�Xp�qn�Cn�b��*��*��?av�+("rҨ� �W�l���Q�׼;��?@0�Xw7[�\,�]��ev꼻;3��23XBц
���*ˋ��#aei��G!,ke-禲�u@�)mc��ևY�X󷭐)rL�Fo��YV�:������<��ugQG��UH�B��+���_�i2	�����24�/��7���'P6-�����29{�f�qD3�(\��@�n]���ˈ.��ogiـ�ٺӭ��h����,���	Cm�Eh�7R`n���\T��qs�,���dV/lne���(�w �K6�C��d��?t("�}�W2�	Y���+�1�W*��Wc��g�B*^�ث;�[Kr�;/���Esk�}�7�a�w�ʦу �b�Zih��휔hcp�g/K;�a�H*��9�9��#�M۹]��	i�X�%\�;9hy[|I���w�HrŹ]1����P��O�(�����oWW:�o�e�!az(V7M�hE��Iì��sFa����:{��n~]Q#Ge4D&�[w�u<��X���f�mq�pr�Z��p����H�S2ޓ	�w6&�1�D�K`��l"]e���ZCA��W�OU���$N�5���m�2��r�������c�1�޲��,����5\���Q7�؍5�=�aZ��k�P	Ym-�t�X�k�W�[9x�@��8���1{Yϫa�Z��Gy.�n���P30)��K(�'	�`J���~��
��m�&*@��n���v�+��F�v�ي�t�ɹ�ٗ�*+���{���3��W'^�4G�Q&Г�ğ�w.�K��,n���I�oun��u�aɄ�-�p�"���hR��+�K4`�N����iީr�x��ӫD�%ې�b5Y��Y])J8��Y�/"h��5���$E5��A�N�jw�l�5~P��y[du.xS/�1�[�_A]��[] Quu- )�v�y&6fRO��W��u+�J�7�i�����쮳DWK)IB-��g����j���V2��]���i�K�:��Y�'KV9�W�r*�)µ��f�N��1̋AWe�gx�r��3�X��]l�@$D�Z��LMʃXW�����(�g��0��W׋�9t}���ֈ5��y�b\��nv<@��<��Ӌ=]xʌ��K��O[K�<���:׊���fy�۞��l	��9u�H3�7���k���[��w(���h{�iU��.2�:3bb��=��-J������+kLn��F4���.4K+s�M!ܙ��}�ePV�)�&{XO^�K��"�d�8j�Oq�:�j���ڰ�ab�>ҙ�z��m�H���z�����.��!�퐳���yY��SV�� `90�Wa/0���nY��8�E0O%�:���+X�4�ש�]���`���M�T4����^ӍK��)&��O8���y�k�x���m�n[�/�f��`�-�[�w1�Fhڻ���rF�w~N���z�K��Kt���rm!nd��fǝ&����ذ_���gP��������x�ᬳ���.Iu���0��U,���Q¨J�`���I2����P�4̂Ѻ�i	�Ք��V��w���^#|��(��ƫ�ۖ2�<8�;�=Ջ0
ُ-n�ۢШ�*��Z�cq�k�����.���|8�Y���X�.�d��t^��扭4LJ ���B'�������e�@�f��n�ڻ{h�Z�E%u�	�z� �K�]��]v�B�7b[4��g�@�T�h����O^��"�x�^Y�{�2�Xc��ݸ��JYfp�p��8���z��	��鴟~ڂ�Gx�m���������mcH�b��O�e�,���Z�@�����e+�R�E1��ţ��ª��1�u�_��CI9Zٌ�p���黖q�{wk�~lY��sy��M�t:9���������JT�O�V�3%�[��8o?|��p�&-u��Q���7�8�cvR�x�� K�nt���{�A���޺/Z�����!�zpQ����jYz18�ҦkY+f��d�n�KN���˵�xH�rq�<\9հ�nF�V�̕��WE*��b��X��9Y����y��Z���WK[�0]����&�jZ�Li��mD�n��2���*bW
�U֫B��[�z!c�\%Vdয�^e����$=������h��6���me��0ej`\�n�����Y�d5�)^l������tk��6�o+��7�+�N;�۝��U�mJ����
���'ba7Y�3{���~ز^��K��Ff-�vn�J�K6�+ͧ�{^�Uh; ��!d���VۣO5F�g�zF�A.EN��f��~иL{�]�7}˛TA1՛�n:�)������]kr��Μ��7h�5�!5f-*��G�o�����W)��V�Ϯ�,F�*E�Y��&�c����p�85v:�1��"�	؉�]�E��2�(�He�f1u�e��؟�����G����gs����b���;ABBº���ol�+��f�J�qM� 6"3��%@@L�[��J�6�p lTr�v]u�k�*�8��`H[hI%d@
U�@nW��+��s�wt��g��ߣ�$o������7�H�I�#y�FzH�I#�$ozHI�$}$�����7�F�II#}$o�����Rd}$�����7�F�II#}$o�H�I#�$o���I��o�H�I�3)��0h�ڱ�W��S3$u+��he6y�m�rl� ��[+[�MJ�P���u�����K�m���v�,�Z�����89�Y�U}J��W�i�*�R.��5V�Ԥ�-����Hڑ�@@�#r�녀Hf�9{`વ��`��}�ʫ�P
����
�A[0V��PAUڪ���G�B�5T�i�j�k��m���;�I�v�G�[���{s����r��2�'��{~���_�]��쒯�t>x�]=m<G^<�n�9A�ݵ�8ǢC���=(���e}�J����m�5˘7n�[��Om*ٷgr�v5�7�u�g�7��:�j*��l��S`;e��Z(R��	6��h�qɍZt�u����?`թ���V�ݨ(7P*u��]Y;g��v���%v��9Η�m��Ô��G�n�xEp��G��X�h�M�`)R,�cj�e�\v�]=�4ܔ���Vܩٺ�?Ӿ��1��r��9{����'?w����fy�k�h��'�p�3�l 7��k�#��\wX�=e�msn��݃��UX�&\�М�4!�����n�vy��|@�����|�(�"z�Tby&+�b�������~�����͜�s̐�G�}�����m�8y+u��յދ�����7�2w|g���n���������}����p���;7�{����O!������B�^�Ȫ%8l�0lF� Q��swErH�<����M!�����R����9ʲ�̍�1��J��D�傳��>��V�}ס��6�M�q�t��OK��ۏ�|��
b�M���_N�.���������2��x����;���/����u��}q�;쑓����nݓT�@�D��Q5��t�:0N	���9pv��:[0�X*�ƚd� XWb��\��.KΞC�V��H:=rm�ܜ��#�9�#�ǀՉ���Q�q�6z�k�ۭ���u��"ӏ�}��<�䝿���{�um��5�9�g�ȵ9^��(����[m�4Q��9QFReCr���=&֢�l�(Ƭ���}�G�I��w�N?����^۶��L��؝�n�[���̶7E�d}����n�]�؃�X0*u��&7X�d?����뭋�v�x���h\ӡܺ��������~��9� ��֌@��紌���e���E�N4���	�������1�=��,�N�d�c���|q��#ď1ߑ�۾���qq�N��d�vG��r��UP�%���tѣ� �
���`�+�wsEU��UcU�����Ywc��/Xh�z��Y��dͶz왰[p\����&��U�66\p��;��<u����v��n��7K�L;���M�k�;{������X��t�Nۊ������3�F5���
^�vi@�#�R����]<�������}�}O���b-�8����3�#��N��L�d;j��Ɠ�6yvܻq�?غ1�mu���!�v���=:q��h�<����.ݱƺQ�a�]q�^�pP���*M��b�
P:����{�E��k��l\7�N��;���9����{�v�m�M��n�1s�G�5�0o������m��t�߻���x��/c��@�۸vp��]��_n��[�Ξ7N�I>�]z�
�u�}�P���[Q��BG��+\�R��Z�KE�+���ɽ�5���;xۯ]�M�����[���Wm��m��p��)��ܕ�s�[\]�~
�����+�a[(�N����دd���鵇l=w�cJ\ྞ�����;r��F�O��q�g㠏������y�N�9l��ȡ���6�X,��-�7j�6�sf�r+�l�l��Gd6Hn�&yx���.��� i���z�Ӥ���#�r{u�p�������۷kc��*j�:�n6+�s��`ۅ�����}�����Fңb��p?l�vEȆ�5+u���o������+�K����t�ʘV��~?}s�i���7�%�`�U��D�9�++�$�)*%�U����nn���>ɍ��Zø������s�Z'��g�w.�{��*tj� z��yr,��`�n�0d�n;�\�6/�]�����
��m:)X�o�y8�x���ʃ�ZD���,�r��d~��܉�OS\+�h.r����9���Ϋs����7%�_Z;�����cΫ}��|�Dou�r���np�rc�9<jʋDQ�Q��PL��ds���L���[|m����u�-d=�g�����x����V�
��*�벻d��'*����sr�zk`�ȝ����^Cp��T�}���o���~4=s�����r/��5�4 >�A�ܜ��|�n�7}��{u������|���s������؝<kl����gA�E��*�xb2<����d�BZ�ʍ��>�2&�I�8�W�0�»��t�nS��Ā�ws�}Խ���=����<g��Y�OI�5[m�ȿj�OPJL6O����]pv�=�l�D�$]`M�<WE�F�l���l>8ާ��b�C���&;����ξ/n�˿�|�GcnO<ah��=���w&���s�%�b�1���ç+�+u�k��7�;���&�nn?W�����Z�v�t�4i7tu���·q�H��7���1�<�n3Ǉ�����h����Ͼ�t��gY	�8��{,�������s�N�֍Ɠ�`�?F[a٬X�6�l ��mZ��ƻG:���*��7v�p��ca_]u��ø���Ƕhԭ�䵭�����Q��m��}�p�M����~es�ݞ��=�y�Tp����R�$�_=���d��Xߴc�Iۍ��y�`N�����Q���l��F�@�#֚�S8�l�����ۜ_ߌ���!�s�:B�_��nM<p��\R�HEW���Q����7gd#�ɾ�:�z�j��Av�����;:�n4軶��e�Z�X�b['�R��?fX *eӱ��x��f�]�}ɟ���x��<��wk�gn�>�����yNɾ۟X�:�z����n��чh��<><v����g�s}����Q~z�.��.��K�LB���
6��A������~1�z2�'���0�Ў�.�8Q�Hs"�P@R��~�jFG�qG%ߝ8C�{)�~����~���:���Rɏ��q���������ꨴ�R�&����;e��Q�p&���Cz���7ømj���!��t6D�)*m�є��1�j�G{wv$�6��P�jv�e��܏����}��$��W_�_c>�vM۞ۑ����wۚfpl�p�A�Xǰ�������]����n��/;*���{�eSptvn|=cH/r��������S� 4�lչ���x�vh�Q�����{���c�����]�u�/;rg���9�鬞J7b��硻~���Pm�"���R ��7�16����׸D����Սtnz�5T��	��E��=�i�S��kC$�$Pp��K;�~I���d:ځ��:���s�ͯr�kr��x��G_U�Y�T��ض�=b` �!�!9T�v���~�k�.�<�3������qO����*~W���p@僨D*-�u�w�}�cy��0gl��/՚o/h6	�pͅ_���P��vzQ�+�F��6=�ۯ}������v����算v� x�w?Ͼz99S����ϰ��/c���)��U�sX��q����H\msߔ�d��k��'�O��M�&�q�o\��i�i�4�tCb ���`	5�v�״�0�&��;�����8Ega���Z u�ّ�RF�`XЍKN��
�X�j=k��wonw<h�����=?�=�oa㗏�یb�9�]p?�n������x3�ɶ�Ƞ�u�EU�BUV\+:Z�Sy���y_|��n�����V�8�=�;�8������\�޻e��R���W�s^��tm�ŵt��7�^N;C����mv�17l�$<�����ǳn���Q�B,�	�Ղ���Y7`(�1x�hӺ$�ss���u�u�jŉ��ٰ�jF�4��ط�v���!÷��2��xb�k����Ԝ�%hdEN1j�
����z��.��{\\i�\�nDx90�s;mb�xixp�m8���+(ՆA����X�w��v"K`��U��f4���@�8�"����w����ǾwY���A��� �YF�n���L��EY߃��=3؜:+��W�8 �^6���~47C�r�F��>�?���]�BS�s<[d���;�!��~�m��ߙ}��p)l`����œN��[��j�	�n̙I�����+��G����p1��ය�~R}ɢ�	�Fu�o���}��x�v�x��g�q��=g�g꫰�O;OM�6ݭ8������l���R��
�G�sX�PhU\v���.���y	�lg����:��?�|k|�7����L֚��������5>�c�=\�͍[�V͎@���]������գ�Z��!����k��l�ф����q��۩�<�H��jٟ.x������#]�֐���pR��+���
�<��fp��F%�6� A;����nr�ql��YCvx��ɥ.�mʹ�<OD����}�������d�2Y�}�~�� X�n�z��N�;��nc�w/߻�︓�0�y����Nr���=ڸ��n�����ɓ�T�|4B���ic(�1]ӱ��mg]Ҏ����*'���w|��[�n�9ס��v.m���h�ܣ�X.덷�\̧nN]�AƊP��ʥ
�S[Z�*��N�u�mt��'%��m�M�6�	�r�2KA�%�]�o-F9�כ���v��g�A�a���k�3���i�#���kQm9-"�֎a۲3YxqB��������k�����m�M�U[#v�0Kc�y��cf�mn㨎��o:T�[zL��c�4� X��7#��uf:��}}�ۢ����#��>yy��4�3�zu�H�]q)�WIO>ú�iN.qAħ�O��ݭU6���kwgf�Z�:.$|#tz�B4���2�aJҥE��5q���e��r\Jh������q�ȫ���t��;�9}knz��wt�uɝy�{T�����s8�������[��çh@�ͻ��ܮN�X]��<8M<&��uRf�u�� ����F�ڊ��z}�K��IV�=����2N7o��s�W=`���:��mm�/3��nt[���<ly�Nn-g]�ʱѧb��g�+�n�
OY��v�.���x�e������{��{��ѽ��ř��5�,Ib����ŋ1g�X��{��y����������������s!\�(���`s%R� �o�+���o��>���Z��ٗ�M�ݱyY��X�7cQ��-@];-e��HP�a���0��wk��qw��w��>�4m�����Y��H\^3�mV8�֔np޽c��{sŚ�mY��v&��-/k=��/)v�jr����\n{i���ݽ��%�!::�.�O����cp�/�	v0b��S;s֣�nܻk�Ht�2�2���V���� p��*+`^�v�]V�[�O$y͠�/:��Y{V�k>��rA��������'\<幧�Ay1�w�:�:_��x��ݽ����nSl�s��=���ψǭ[���a����#@+�PT�I؂1�H�����-���a�l�-�z��wc��8!Q���G�ۢy��7+[��{��u�Gm�c��̞0�Gq��Ɛ��7;!n{[�F�Og\a݋[uז�Ņ��Z���a�[)��V,���@��_kcK��϶0�Z��Vq���|e��Kg��㒜���%�������&۵��s�鋄��ە^����w׾��n�rg��v�'\���:ߏ۵��p�4vü~4gs�PU7X,�;�����{=��﫧c�_lu�WCm�n�p�8���p����9�'
[5�Z�i5��B�Wx7Q�}�`e�;��n>�8W;�6�'�U��)��n��|�;B��.{{]t��g�8�r�����ۭGOm�&6��^�7�����๡�.vq�*�Ƹ$FT:�
��^lZ��;ۇۃ��u<���Z:㨚�{<��g��������s��:�]�T<��T�FVWDR����?V�p�M/x�9�Nd�M�[,�yzK<
v�'of���/ͪ��= vF����JRD���~���nߜ��m]������<�bL�T{���v��0�t��<��u���a8�юGa.��! n�����)Ųy�Sm��e�Y��jf6;�ͱZ��ڷI�\s���EFS�j��Ϝp����5��rc�Iϔ-]��bX��BIfb�X�31`,K1$�1bX�31d�Y��}��m��ݩ�%dٱ����/�Siz�T5��3��t�^�y�ֲ\�oj踻s�C������D��qq�b�.�dJ���7q�}	\÷�o7����\s�v��w������J��S�A�����7�v�����7��a��f��"�\�ZnŃ���g�+��/W��\6W[c�c��m�P�<]n.v�[�Nݽ��S�\�n��;��q�^��g��H#��3���d �!�r�y�n���q��#Fo=:n�կ/����3�b̬�)�[���_���^�^����Fx��LtC L�U{��XV���a���W�y�^u�C�"B(9�:�O1[�;�y���WWae�{�Bz�Z�P� h�3+t	P/Qo��83�J��U�}nE�ZVs0H�5���%⎠۳x�Ok���V}�dG�j�+�"��a��wö���n�j�B3��)�U��ƶ'��p�4�Y�謲�ݝ�vcĈ��7Yʦ��m��1Fh�F��D�) ��I;�l,rm�P�Bdn�Z*�����Nn�_�"=���췐zd�a����{�`�d������@�q��� U�ƨ���͹��O4������r����k�N�"�W\Z�N�س�������#�zsB�V^�E�א�� ��Kk�A��|�5���[�7=ʈ�dcv�P�9���	�K	^a{V{�^�o��Z}}�d���}��A�*��̡��V=�y�����9e^U�b^�������C��j{Ʉ�Z"��R&�s-4M\E�o{�E�9�u3�h��vΗ�����
��P(�C��=�^!(aICnOhC]Q�'w�G|��ɜ�gk�T�`�rx�Tj�{N���{��}r�9�����ID��dO3qn��јr^��k�N�d����\w
hi����j�NWs5�>z��9k'Y.Ԥ�H�$�k��&c��ܷ%OO�e`�r~���}F�<�E�^m�;�u{��{���8ue;Cڧ(�l��f�(�x���UI�˕hT�Z2��(����V��(�֢�^l�4L��A�h��"��g[�ŗ���d�ֆ�afs�B���P�Ż����xh���q��z,��g[����#���x�aTEK���}{����I�x�م���qZkfz^ve�����+�徺�o;���/x�d��f����O������D��]�I�+�;tl-�����wrģ�Mhɳzձ��L��D�8��c��n�
	0z�U6�Y�������nm�leԺ�P3�8��ErW�C��-�h������<��^9����^���o|�kUztVIFKH�m�'��2���-ؗ�V�w��3����!�RbZtRy^�w�ݞ�9�E�q�5rM���<��MV��PE�b�Y�9���n\�t�-��^�g��ٞ ��z^��;���4u�*��]�N��������e����y�����>��'Q�����g�E����9yۓ��ζ6,鋛�vw8Ŷ�Y9��.��נF�P��ɧDVh����քV�/SƦ�0Ԉ���ɨ�nJ�%d��J7����.��V�_�``��G�S�=��-�[	W�`yf����]v'Gq6��w/A��*�O��C+e,Z{�MLֽ�.�{�!h� YX	���B��{kfqL`���t���I���Ь��{��Oͷ���iz����/U��|���D*��������S���ռ����N�5��>$�)w�ڷ��#s.�X}�'�+;E�(�|����*�nt�'_~�&�\N�Gy o-rE�]���U�����]��z�E����p���n�����Ԭr,�t퉫}��E <�˾�������x{ba�8���vz���}�8ol%�|�x�͖�{�}]�]�5�^N��]S�mEdE���#RT&����r�wS���nquј�;�b����:��^Y�&���u��hl�LeQ����6������'7C��f��Oѳ�f��������_����b��Q�������N�ɍ٘pF��+vD���v�P�u���R6!�BR��k)�ﷱ���^m�ľqu���Q�`�x��AU��GD�F7s^�mf�Z��_�'<�Û�5P������ҵQ	�&�r)"��jѢ�Ih=E�ӾS���:Z�aQ�m?_X	��4Me�fϮRKU��b*<s���5�i-�-�l��ex)k
Ҿ( ��#�֮�_o?N�L���sQS|�{��2��T�k�:�Z��u�c�E���^���x�
��Y-BBG��6��s�s�,sF��8"Ԭ�uǴK�H+��8Z���w�8��h�ю�l�>��x�=O91��{�}a�:-fe��y�Mٺ��c�<�sɻ�}�����)˲w. 3��⛑�xk���:�jU����,=�x�v��g�.����u��v3����@��B�����2����vG��'<u��c��+c�V�{h�n�V��y�����%3��j[�=���5�Ν�_����=r8;�w�0k���n,�0��S�����</8kk�Y�x4����q}���g�b��q��� kqֶm�;��4��(��m��������v�1�us�F���XX�*b�ܝ���l\Lb"�	$~s�o�����|�|]n\XE��)6��R��Z6�𙭜؜񂑪�!A����ޑ�i�
��U��3�E?5���:#���;���x3�}����o���+�V�Yd@�=���?z�(����/���'�p����߀�Rf�g}�Kv�ZsJsyՠ�z���pQ��'X�\O��_�w�{�<�uZ�n��}�U��Z�4�F=��=ow|	VM�o�2��I#vM;�wǘ��N�)dd�ov�=�^��s�������M1�-��R�a����~�$���~��T����]K��;��qkj��}d�8��RO®v���6u�������&�6xǘ�Ƨ���kŮ4��!lL˥�E.�<x�޽������,[�\t��:��9a��݂_z�{��]L!er���w����YI%i�vsf��u}���˙k��^�_+�m�BfV����"�]�oc6��g�Q�f�V;e����}cW:��D���/��3��5+��F��}�"���v�/kF{�-z�*SS��wr�=���,M�����iye����UiB�,�&snd#J��n�z͕#$^�4�X�s�^>�����Ŭ�B�ML+�a�	Ɗ� lX����i߸�}1��"����̽�׫pD9�J4�}8+eͪ��]^'�2\�d�~�6�w��ݭ$R)�;e��h���~��o�ċ�9y����;Ȥ{ۗ��<y����o��mɩ;�5��\��8��r�������s��|��MvD{'8��c�~s�|�3�m�����-"" �6���48^s۝ϩ���&��;:���@N���ݤ&b���n�3< >BY~��\J��~�j�r��}S:�_g��\�z{�B�gc���!��ތpZ,�/2[]WY�%	US��6�7���
mz߱ǲ����,�MО礻ܹ�w�j湿F/�@��N���t)X��M�g�h�2�$�n,�<7�s��{q*��݉jn�"�^�E�2�g��򋼷���DAZ��g{D��liP7�1�u�>~�P�y�����	��jn!nf�� �� m�>iz�}{�]8�613�KTU0�/�bQ��9y�X����9:{��ެ8^�սլ��-�@dv��G5�.h��U�M"��_��&^F��^zk dG�������h;��Z;7��G�S�{��D���N�<��K������=۞�2\�њ�Wl�wF�±��Y�̑/j����۱<��r����3w�����܁�?,�Ǿafmy�%��tĺ�4����on���9FǾ��{fw��Y�s<�_>�o�_�^0��m�X��ŧ�����dWx,�J�����]��n~���Q��%yhJ9-���3��딮���R�\�4�����{|o��j�Τ�_�5o���:���3�/zw��������h���尲X*���$��gi4�=W�D7�nє��1���p�+ވ�����K��ͱ���`$O/(^a� �D�,ׂ�[X1@x6�f�]�Z���b�S1:
ӗ����Ż/� )��;� �R������
�$�k�p����u��MEP�T�qE����'*��9^����x����C=��sX��<��>�e���W���n��>��G���7�@@Ӝ��b�Cs����v���㧵��8���NH���k3����FUd���Ap��&��n�u�����Fm�k��&x4K�Au$�'LÙ��s��{W*rl�T����D �ïk�E����asS�қ�[s��w�_	�A�'Y}��*��מZ�!�w�A�]��AH�y��~��Ѳ�QWj��p�����曳8��EEݓ�8,`	�.{���$y����Ov\�������Ai�J��-�t�f�#y�M��{����.HM>z!��wq������V<�Ni>��
���j�iX��* �-5'LDC�&!��ш�F�B�N�ڱ�ڌ�c� �F�$�j)c�j��-��Tb����xvIag�[S:Y�>�,h�7�kk#�����l�w�2egf`w�j�5'���:Ȍ��=X<-��k���9��5�"��Ch;Ϋ2����J�;���?�u�og�:��7���z�8����n�k���8��[T#���K�7c2�\V!�U�`�X|I�+��+�B��Tj��=�jB���Y�Wn�����#�[���y��ܮ�/Gv�n����)���kq��C�d^�{N�o�|�G�A7=�9@�M��}�j[�fwv�=��T��`x�����I��M_���ۑ�ۻ3ۥ���}N:{sbwrYI�N�mӻc����q�MK+d$RLD&y�p҂VwS�s���qN�֍��qŴ=�-���E:�s�:��So�q���¾���4/�XѢ�c���=�`��_�WN��,y�JN}L`��ŦŁB��g�?�%F����I��xR��X=9��_z+Q�{�1Y;����Ja�pq��ס�:�ZH1y�Y=[M���e3Kٕ�ȏ*�m?N팬�d�!⌊SD^�CH8E��i�p��~�}[���M�"�^�����[z��B>AxFg���w;k�i�7'���95���l�Co�՞�&R
� ��kʨ$�[q��S�q.��ؠ����~;Y{:�z(�ĝ׈^�R�RQ�c�ѿw~Z��uF��Mw�l���PMYbz{%h�_5��=�뇦�A��[���+���j�e�q;A�V�x��پj�h�ח�$���?�K�i��X�՘oN"x�s���>�[W��	�	;��`Q�ݙ�t��&�<U�M~G��ָ#�)�Ol���6��Bz)ܯ1q�[��}f-ˉl�@Wd�ͺ�,Y�F@�9!33���O�~�k��Z�����0�f����_�Q(���q��
�݉����wP�W��˺Y$�Jʄ�
��&�Z:ߦ˰��w{���ɒ�<�]�YI]I�!��`����}R�mh4nkw5�=,�c��P,��{�W�5��%K�y���&)��	��H��a��p�8�NʙF�j3�ìb)U˙����n5iBFN'wS���H���_��U�`{]��/rg{��f
M�l�z��^b����4Eτ��>ޱ�],�|�h��#�U:Fڭ չh�{b́��u��/2\��4��V϶�}	��kR*j*�T�������LZǮoW�>2)��U/l�nH;&2�-�{�g=�\�ʏ)�o�9���~ew�d����6�`V����t�y�Dqp������I��0^\����"f0f���sj��ƫq����F*ٯ��6	PYI�6ݛ;�$K�j|�M�3�,����1���GO�W�9��ʢ~0�r���v����"�1Vf0mp�m�Y�e]��4�fM�f�ڠy�Ú�vn��}gN�����qPF�e�&�R�.~�t���k��2��el���N�遱i#u��e��eY���ع����w'3yEVP�|k�Tq�3�^�$�j���wAst�7n��YoV�g�y֝��(�H<|�f��V��"��FV��������a�뙼�DL��Ԇ
`��)j�w������(n���]��uG���7Z�x�-�2��t}{uf�8�Y��5�ϫOO�w�o5f��o;��Y�$9���Fb !�2$�"R��Uǭ��wN�_�8ko�*��Y�ٳč��W�ё �����;ǜ�+$�[�O�9ia�<!�Xx��9lWsx֮ SL�F�,'oe��Dh���/72�f�j!�r� �X^�dH��p��3�k�P�*��WO�ʉ}זr��h�k�*vY�#������؈�0f��8�6K��ݕ�6����f�O;o) �[�~��яgftRޚ�ځ����n��-jX �u�U��F�=pat;�Z���&ք�uwl����ͽ�U��m>غ�]�t�X���S��n�n�黄���Ԗ��2���ש*V�=Ö!6���x?E)3�4rw/:��
+N��Θ ��9��'�F���˯l�v�wxs,x%�OlW[�X��x�-�ȧ�b]Uݺ�M�G�~o�~���*M��(����,M����E�f����=�����yyu�]T�<1׋�j�Q%��{��ͻ��Lfi�Ϧ/�Ǟ�����?�*r��I%���t��ɢ$�?�SL�[��Ͼ&= b�Lu�tR��?G�a�+�-������L���L�K��pϻ=��X�4G�8�#������uO�}Ə=u�r5(_ �����݁$QDDF�?U(�!I��.Ը3�w��:�Ӛ���u����e@�$A���!��~ȍB���d�T� {���G��H�	�@OOy�~�,�#���wc
{ҕ����bbP��0ws�"~}:��L<=i�d�nյ�Ȋ���c��[��������h(�R�
ų\$����p��2E�ڐ	���J��x���A�;_�//�]���Ͼ�p��
$���b�Օ�;�M����� "�x�_&�JF��b�N�S��vuZ)P�,D�������ה� �Z��V�B��!�@��t���H��l�8Y�Y~��Ֆ��~R�����6�����o�9=]���Q�o��Ī����|8���.`}}91e��"PP�ۯm/��O�,XH/тb+G~����o�}<����uJ~��If���[���|4���� j]��Y���ȗi����Oj��IKEL\�ļ�z~u���O�-��[���|t濽_p�|j�3��׵]O������@��Ԇ�}2����?}d<�=Q$��l���,!���_���(~p�,k��"�#��+^�����Bn���蟈��i������:��c�طib�V��yS1�T�u02� ����b�߼���~�Di���1Qާ߼rZ��R��3: ���^g��%N��寛~�s��i虉3%k�.,���z����_}��^��8�wˋ�1p�.^9�	{�{W�/�fC?"b��Dx��\���,���""� ��8yϪzx��n�v.� ���"��k���:M!�r��d��h1BZo�w��c;�ۼ����[4��?�LpqeH�G�j����1�^���������촶�r@�w�_�x�{�Æ~��"�՜�?{u:@�V��~D`(����k�(N6���%�K�ǽkJgt�����F͛��2`C��u��@Q ���S3S�"o��'�4l�"�gѓF��x��Y��������7���	��qi�aK�e{7$�(�q�mE�!5��
��%ڲ����۾��̇?}�9k��@�2c��y��̍?-�g�iE�|�0W��b��%v<�"�� �`�+�r$1��D>q���h�4ͮa�Xx�F�H�"�߾x�2sox�el�-q[%����/�Y�>��k�z��4��dA%W��Nf���+��$n��p�}˨1 �P�#�Ih���1�"0�(���7p��zC�_D�ϰ�Nsg���S!t
 aZ�ٯE~`4�����\i?��d7�Zb��{�y�ē�N�d7��y�(z�m��ȱ~���[�}?t� |?o�$�I��3��d{�7"HcLK��&$���>���K��Θ��ِX�w�g���5���2���[�TX�
,:�~~�u��rq0Ǎ�3b�g�(��ᷖ�y��j!�d����/���$wseV5�;Wc2�����E)����-/¯�C�c�ࢿl�w���|��H=�^\n:�r@@B�K�P��nUl���q����������`��t�����ݩ��9�!mv�09w�u��8�l�q���n��;kHYm�A��p�q�����[�������ku��ٗ<}��m��C�-�J	�f�������N~�c<vz�]퇛�X�W;��(q�{	`�M�G�ύq���m�����m�W;�]�� f����Ƿ�}q��ض1�V��u��tuWZ�u���=Ð�2�ҕ�r��ߗE�ş�,��z����?�,��xbPJF��<��5�#�%��bffzfp@���M��D��,#IR��|HFH t�\��$[Hy�ԓx���Ş���5�L��1>����gy��ĿzԾE�>�Ĩ��^>w!%���,����, 0�d|4\�Lb�ׇ�TŁ�v<\��{73<_���ߗ�w4ļ=��֖�,�~�����n�t�	/|~�,�%�P�G� ��e9� #�~�i�3�/��]�x�$���.��ٙ��|,�TY��<���-��|�	1xz%�≸φ��m�%�R���I���D�b��]�>Ӥ| �'�Y�0���E� ��#k���kUy��������g��j_I��j��^��.�æ~����,fDf G����n�%#Rj�i-53w��U�E�O���q�'�J7���#����Y�$]@D�����@��c�D$�G8gO�F��M��R� ����~e�!]�|�u�#�O�6���f���}g�4}�W��n��X���@�h�lE�P��q'� 3��adIH��a?]���~�n��vlƺgۚcb{��$i�r ��j��<G^��@��O�8~��*[ִ���[�w�W�snx`Q^�`QGn>'�U9���������QC� H�yS�q��;v3�r��cl���Z�dС��7,odݹ�=3��_�$�@���M_*G�?q����m <D��;K�d�ȳ���Q��!ws�?m�Ϗ�"C�9��t�$$�8�p�+�"�bz@?#��|co�	!�U������������E�����Hj�Ӻ��_W��ϩ�WPb�Ź��0�wx�wi���Y����;�U{�i0۱�c���l�B0���)
�]1�q�1��|H]u0i��z��d ��~
�}՝v�7�>g�0F"Zlֽ-Y~~��#� c����"+����=�EVi�4�������#ĆqpZM��2>��<G�x�X�{'yw?��gk����i1Qolo|�ˏ�ج�#�w�_)}��x,�?i�v�b��s��
�(�x�x�L^���5t�F��J��kL�{37����#!�І�a4M�r�?)zX�(���~����ϸ��§��'�	��X�LY�?o��ָ%L�\1xdLy���!��D��M�Q�\���qW���Kh��n�r Ϡ}�mGÂ�_d���b��\�ڳ�|~�3H$������=�.��p�?"<�@V@�Ln��.����*�(}�Ǟ����1~D���u/��c�����g���6��R�_s�gO�ÿ��~��2���F`E%r�<ꬣ�ϡ^;�7iȦ[��9狵Cإ
�����i�ȴ�5�&�h��Nx>I��<x���8t�#������1� ����[�8��S�N(�~��D�7탤�"?[�?D�o:�n iG��`��$�N�`D�#���W]��LZd(�1s��>��t���%�5E�
׉�S_�;�qcR��#l�g︌"���@#�����3�>	p�����>��h�&ϴ�򖧏^}��~�� A��	�$�ԉ�[���8i��pP��pPK\�@���~/�dY�y�pI��|w��+�	|��~Q�tw}s���	�Ń�'T��vN]�
K�V��X�h�h�#�_����\ K4ԙ߷���U��}'wfdW2yu�Vg(�W�T/�p��ѹ��9?|� G�?���|_���Z\3<�E�{�7���D�7em���Y�>��fi=��Ҝ�����}���H�|�8���tLWL�����}Z���4����s��s>g��n �iD]Û�&����<�����`����j��Z%E��ﬃ�B������h���D�Mn���Y�{���8h��>�I+�{oEV:�h��	3����~k:p����O.H֜1>��5�w��gݽ�V�L�E�lP]���P<y��O�zV�(�a0����I�-��۪�&.MOgN�F�P�wnt:v�V;#RRIo��<4]�LL�ƕ�>�8���2���n��ҏ�\|<r`fJ���2կ��8����?V�tJ>�}�α��_�v0K�?�|�ן�4���?r�3ч��>j��ެ]ڱ2�*�jH�����t�gǦA&/�w�`�{�Y���#� ����� �F������C�Lb�c*@� ��N w����>d�oS�U�M8����tU��>�P,� ���Wo�C�I�5-������x~}�3�y=1��=� x�E��G�q���F�R���런���������hLxI�F�"�v\�"�Ẃ&r#��j>}�S�"�^D��̾����}b%�)`U6�����=2�?a!����
��� �+�H����i���>�"F�󟇶>�|E!����@I�FD}$�9�NUJ{E�Ϋ𮧇��"��-�D�+7:wH�F��۲�kn�PhN�F���mgAb�n�r#-f��س�ji"�|k��%+z�!)>�~��G��tX���LI���o�KUM�PWGh�ԂOz��������ދ��~3�pNy���y~�Y藆t_�q�Q� wR�	U��(�\|��Qޅ�����w:x-��S�ei�Ǐ�^��sp��+�c�B�Wln֭�ub�-j�OT�؁[zֺ��}��,�`�܋vc��r�]1��/5��b��ڳL�Iy/L��f~��x�����EI�����gc�9S�~���,��_������ytB3ң�q����nӇT�lt\��3LR�/�2����&���#�39}�q�#��~������OC�bu[_Z�}DYDB�0���^��^{ a�"�*���'�� \�U:�����{!%�����&�"�.���܏F,�_i`.*�#��D�nW�	/?5L�g��i������J�~x�>���?Q���B^�s�>� ������/I��� ���o+?�l3��z����^d����T;u��K�=����^M�j-��B�	��3�(�O������$�+��#�i��t ��$I'O�~�11+~���w�t��~�5�e�D�5�����wN� �D,�xb�Ά��Y��VO���?	�͑(���V1ֽ~�6DV�?QP~H�q�G�dA�U�@�\�|G���,�!� �?=��ov��x�����%��!�}��A���<G��~����@�3�e�����Ģc�K�-�=���;��M{<<�#�G�n(�d)��2������=]u������������l�f�]F��;cy��=����;ʕj��K��V�c|��|�e�рh��7x=Bm�*`GB[���'3^�=s��^6�݂��oGM]�s��\�Vݸ�;Q�uy���tx��a����gr�s��*%�T�!��e��cN5��ؠoV���m�:�&z��Kcet]��";@>جiւ��\9�g�߻��=���r�G�^�s��lO�7kr�:����l��l����\%��JA��Nr��:n}?��w^;��urv��&]���mu�����ssK��Kع���]&m����MT��,_]��3�7濞�Nk�6���}����> PK�}vb�\8�|B��ȝ)}��8�~�
 0�\�G���;n���F��#��Yij�G��d��~DN��4�?]j��Eƴ�=��r��R�-?�F�����i��4��\�����~-���Izً�o�6�%W桀��������8�A#� �E����Z�HY�6�hQ�ع���{1�Oǆ~�^��YJ�%���n�/OJ�^Ο��s3p>�q� A����HG�<G�D�����6d��E��ڭ��
`J�@���-��!�P��Au~�9Ǟ�<����K���e���?G<�~u2:�h�$��䷛8?}�y�@zp��4=�H�7���������!{jȁdQ� �L�˽�*"�`�d�gb�"�}�������M��fm�$��9㻜�̼����2B��� OQS��ot��K%M�ֽ���PJ��Z��o'�s��S�ȼk��Qn��z��{8��~g�/��e\d
<n��u�e��C���bKM��C_�<��L�x�����ګI?|���Ƚ��z
ی��9b��H6y����~;���GiU1��Ǡ'u�1�n�8��"���}Hiq��X�|���qxS�\�I���V}�^kY����~<n�\�G��>"OÈ&Ȃ�� 8��,_Gٚ���{��H�r���ĢHU\���z����B��k|G��\f!26��S�ͼ�����/��x Ku�����??m��O�`�1Թ�bh�L��+�b��M�;��7{-�����/�X�3�������X+�b�87�<���]ڙ����s{7���=@C�0D��2����n����A�o7�H��b8�8��\	?}� ��V��5a��n')W��F6Lj�n>������5���r���+
{��iE]i}�_=��,��DY�&�,���q��-	��=֥:y�c�f���V I��cH�ݡ��$}�@g�~��{�|t�{fc!�kLS}��?)%%Q�e�ݶ��x�x�쏬�g��;t��.b]<;��OL�� �Y��E���yŏ��I�uȳ�5GD*r���1w�����{��|���<f����g�A"��5���AgI�~��:��-{�4��4(��[��}0��{���!2D��cR�����__zm�?h?y~����h��b/ݫ���3�ɥE����{7�~1�Ǯ��>LW��2��u=��\G�BK���b ��X{=@{"rv�s��#�v������8��ǵ-��N
�B�[�/>5�IW�6���>>�=2R��/E� ��_#<>���3x���?2��ѧ�W=�C�L�R�|	(�|~Do��L���g��}1�P3��$�;�V���]m���r�b]I��L�p(��wf��:�i;n�*�4��F�#�z�Q�}J@����(�I�D�6B"��쯃V��@��-&�L��}��]_���|�<';��n��7�zd>)�;��h�U���r��E�Sp����gV�)F��{�O?	Z��Ě2fo��[y#�?9wekY��=��Ù�f���G�k��0���<�uˌ~S��kU��~ꓡ�F��57yv�:S�U��Σ�97UR9���|p�$���?y����.�V��/Hp\=8$�NԿ��ĘŨI��}���v�X�B�K�~��ǍQ������:w�aG��o�}���VF�0���vq��	�W�?7q�\!}xq�ϼ�p�u�3�h��<�z���Q�[��IQ٘�H1 >qB�b��kE��Ry�{0�%��,�	-�d�����0��_�[��r�Ψ�*2W��:E�9;�7��(�O�����=/�#��̟��D��A:@�fHY~�sy�@�&�_�r�8��,��	i���3���0�-Q��j\�O3���K���:��3a3��;7]l��bK�a�S%��&�D�� ��j�-k��4����U�2��(�۞�מ��R$�@������M��n>g}��#F#v謁��3&Nq����?I���ǯ�#�W���� �R:l� aQ�у/�P�q�vmY�'^������.�6i�H��5�?U�.|`{>�>���){/l
#��(�@DI�$�� Eur��TJ��s� y�䨏��S�A�F��,�̪���տq�ǈi�CÎp��$�j�V0e&�����3��4�2��i7ȗ�
z~����|k�g��^~c A��E}�l����-d�����?,��DI�$��D>#�_���	~��}�N�ޟ��")	!|�\����q�A��I/q~:`%D�/���'�/�fx.k�߽���G���##��@&폲�� �G�?I��V�)C?|�{
��?��ǽ�����s:X�̹B[��Ozˬ04+��q��������{q�l�ĵ�ݣz��*u��R��t���e��n�[���FO�~�7E�X��,������ӻ����C��p�k�q���4�OO�Q~:A?��.�.�JH�# aY���[~�zC�R1�"����`M���5w�߷OPbDx�_��K�oo�1KA j���Q��D�"�2�"����|?����y���8��ݻ=G��mݤ.�n[8�m���:$��X�X�(r��v�%�|���D��:Mk�B������I����u�.��h�K�7 A�r�L�7=y��<�yw�}�����i���G蠖�T���F/n�s�yy��0<�J�2�Z�;������Z'hk���c����$�eh�A,�� ��R�W�9�$t�ǩ�ߩ��W�������ļo!9��<>�Bo�{KF`��G���\�{߼�9[8�뤭o�6�1�C`�'�n��QhPB��уk�͸G�~E_.��oE�� ��A�y�����>k�N�g[��]!��Xw�]��ɣB��C�4 J��\��ȹS�
 k�s��}O�J��%����#~�)'�L��J�qF�w�/�l�qHl���92�%f�����n����9_>��c�ʯ!��/l*7�&��O�~ݎ��^���On�j�g������9T�!�mQ��b���=3�wZsqn�<جb�9��>S�����S�=�L+��)ę�g!=������9�g���{�&f}s�����eo�@~�+��ïr�V��>�%g[L_�x�bsY�n��ˈ'n�M�YZ��#�Ge]�DC}�q�޳9�j53.��ӭ���ٱ���(uN��3���$Vft�9T�
]����j��;�+/��@�!6p\�-Ûד#�ȩy2A�~T�#�u�yq�d��AV���V�
s:=����{gI�0^ݴ����'n�su�u��n��5n�ؼ�!�GI��}����4��֧j�F�����	m[Wv�ic�	�@�Ȫ>�r2>"L�U�K=�m��;m��ى)��N��gm��u�v����į���_w�Ϧ%3s}b�]��@Q���|��2��o�<���RcwVl����C{��/���VR�ol�^��(jR�2;�b��r���h��X�Kx[!Iց��<�l� ����Sĳ�#VQ( �>1��3�]u�ڵ��!�s���K�o�����ޡx/�j�W@%N���d�ʺ�IЭ�N�x�;�9 �]i��5��@�J�)g`\;{�]$�ʜ���wR�xE��t�oS���^R$�;Ыif���p��/₽�4-��n�A�j�̖z$�)�3#X(B8��nf	��0�z�m�]��/n��7��gl=tʊ�ڵI�qQ��W�oEʱ��f�����,�R�� �g�q%e��::��b�	���O�iCV9�ӣ�}&9;wJ�B�o[��l����q�c3)�˦��2�J�����o�Eْ,�rmX��f�)�z�����YW8^e��ƥv�.Pf^��{X�O�ϧ��Io�}Qg_^��`��ݺ�m���'Y�^5s��?u'
��@d��ڥS�⩕�pu���cT7�q�e��8�wg�]��x�//\�����To�~�든�M�C�M᭢r;�t������nˁ���;x����c��y�8nю&��o��3�4�l۝ǭ/f1�uFGY^��A�¹��Y�6��[r�.wV�V2gs�j�;\���v\�v�<�Oi26�y�d����'n�y��C� ��"!j�����S�,�f�Vm[��РQWgn�ȹ6zN���q~/�����cvgv؛���*��vc�]v��/�
PR*�,��?;w]I�eu�g��#10�b;e�Z�=V�l6M�n������	i�
`2�s7+Fz.�5��:�o (�<s��{��:�)[�*�n�$�Vw�d�J�����ٺ-�<��s�v��4 K�vu��vwI���ƶ>,���X-ٸ�q��=yq�ܯS�8��^��!�LX�^����y:�����ý������,I}�n���ǩ�t�y�� ���GP�e�LUdz�{����@�]5)��v��ƒ��l�Q�Q"�Т������ro���H7Q�H�Smî�&:�as;��ڪ��wg�=uQO�qgc�i���OW�p������J�KIE�����=���hКnXJ�f`�B���Jବ�.r���%�����m�qum���ޭ��I��u{<���?>��{;v��������n�pz"�����(��D�s+�؍#��h����.�;��^�}�;vH��W.q�ͫc�C��~�9�A(�6�n�͑kV�r���(u��x��F۞ͱ��bQ��2�N{p!��G�M9����w[�X��ev��b�\�Ƿ<��f��=]nr�g\s�3�u��/W�}�)r'�qQq4"��{F��nMٛg�{Cb��q�����m��N�5�r�;��c�L�֫��n��>�uż:�7Z��Kg���[v��U˫w�*�BL���c�	ejVGB�P���O/3۝�y��{$u���>i��ѿM���/ۨ�#js�X�v���\��i�ݽ���V�vY�7]���ŭ�B�lu;������;�I�s��m��(�=uk��r���V&��pku�F�[zN��fŶN�8]��]��;�)m�֭c�fgLgs��#�ݝ:��%�8�i�+{v���г����c���lg�0����s���tS��)�y/n��Gcs!q��f�F���(^�pP<��4�ߡ����7CO�]O�XæM{����s��b��q�o�K������l�ij��}��8����z3y	�Ap�G�r<r�*��PCP)�&��o2��,RE6�Ul��ݨ�ȸ�+��q�2�k��f�&gc=�.�����>�(B�n7m���7��fe�h��.��~YZ~�'\�H���V7(|��5_�����u����R�/|�S���	i�E��A�d�:�
s���˞J��~��FF��>�r�wkQ��o�흣P�v}+ �-�7�rNX�y�'��s���?\}{�.Pӽ/�|̴�GQS��=>�s���=�\�=�(�65{5��!�ǈ	��R0:.��,�����	�0)�?AUt�D`1>���I��B�����=� f*�j��@��U����P8��/6)�(����=j�~����w{ټj��F���(R�B���vF��]��{[v:;vM[�̮��Ź���{(D?��M�|�g}��fN�>�b/�v,��$F]&r /{m�B7��`HwCpj$1��O�C��א'U������'���wX���	6(-��+��#�Q����p�+�ܱ<�S5*��C�:+���0�,���pq3v�r����&�uiY��F9��m;fܝ�D'/��Ac���WnV�ֻ5�6BU���zwtH�yqݫ�,�Gٙ�O�x���G�Isz������z=���<�G7y�r>{>��i�n���l}��k	�2�����j�\F8��bX�����μ$��y�a���}����fz��)jC��D*�P@>��z�`�^��v�\���������S����q���d��	9�#�:�]w�J[1����9�a�{���zr�������j���t��ϰ����j۱N=�'n'���=�����W*�m���w��j��}���?G�e�ս�ɋ�ܜ�3�+�u�6�a�e����m-��:��7��V���g��F5�c��Nݪ6��$g�&��ŦBZA�`WdQQ�u�+ə�pV�x6�<k�ֶ�XKs�����m��C�*�
���A�oXſG�b���E�`94��7���e[ɹFD{G٦/�>O;�Ƈ��,�=�T��Wt�U��Vz.#�+�����g����@)�bRr��ڐ�B1�q�����[�0�0���CbI�\A�f,�R#�xw"�߂+��[�W���S@�%��<�$wj��1��E��f�*Ne��A��ȼ�~���1:�ex�7i9��D���/�1&|��XX��PJ֪�6l��wK�����+!��êZ{��t��^P�8�F:�}emfk�8���]m�YQ�U��es�S{zwe�%�fU�Q'V�c�S�񖾓�U���=�{}f2����h��0Q�o��	�N�� �a�~t�u'ў�a"�L��N7�Ȟ��*Ź�J����=���́��=2/���e��Mʜ�!�)�ҭL�xɆ�H��U(.~���mbײ������֘��E�?��;�ܜ��rC�.�*�1;���"��������ԠLMϛ�;��UF(��K�
�Dx��c�J�~t��*lv�@n�H8�JY˼��v��s[���};8��&�H�f�;]�(�q�$�{�V���g8]]|�
��^�B�Tj��]�w��#��������"F{��Ѯ�'tMAx]dtuZ��O�׶��Ƽ����=�ٲd���1&���-Z���_��}�>�Rv	<��]�ͯ��Ě�E=b�ߣ�!N�8�!T}��4����e��;����ߠ�B��)�CF @i�!�i����|pӒ(����"��
����5W�C8J�\����"��X�=�#>}���Fu���G������j��i��gs��o���RAB9C�7�xE6�7�b]�w34I�y�7quyUG�^��>���:Eծ�H�������k��M ϭ<�>����p��㛿��;��<��7�v��T]y�Az�o42Q�^p�Զ�e�Y���S$����}�u��8xL ����+�`t�ڜ�����>"1\������v�L��G;L�� Vɮ~���}ev^�%�_��|��ꋪ6TQ�A�{�NǫF���vR�4��'�~��k����-��vDS=���k#=���r������=����:-�[ >�1u�;L��������^�?�`�aVw��D<����n�e��V9���f�[�;�����z[�r+;��E%��V� C6x���v�=>�16Κ���n�	�����پ��밮���J�_^5~~�����Ǿ�9v����.�f4 _d����k��D��r��^K�}�s}U���y������J\��>˞�N���/Sh�H�G�a�N�'�i��4�^us�ه�W[Y�sP?C!B�p1����уމ�w��tg���~�6�.���BM�.V�w��f1�F�������]�9���ꯤ�������A�Y�1>7����x�b	�g��ŀ�7jnT��y����E�3�^�;t-9���(=yվ��֣n<5�a@��:�B�.��c#�<*�+(H���		��xZy{��\.ý�[�����oѐ�N�[N���b�=�O�Qw���[�K$��.)q�����ш����6nx����ӍnC�'#�g�y��u+�Rڷqy�}��}�����_r}� $vr&Ĉ�.�=�;��C���sůp�a��/cb@$
�~�v}���px�4�xꗃ��i��bQ�uvם���7Sv���Ga۹�_�Z����b�E�^�]�:��q<��{q ݻk�n���胧��<�[�R>��\v���}��Sʇ�;.Nm��,x0�����F�fk�i�0!��[���H�aLe���Qy�b���`��A^O�Y�|<����2����F�B�1&Q�����^C��tj�$�b��B�G�s��3k�yn��Ai�Xٝ�-�hGöS���5UX��p��M�\a�f��z&/o�"W��g�7i�$�*4�Q��N)��� �@�Ȕ�y�W�~���>��D��?\��J�w���eL�;��B��-{����ǜ��r��#�u��xK}������	8h�k�a��N��o4s�wI����܏�>����y��7��,�_���g��sܼ���WW���:�{�9����0�I�!�Itϳ'/��̗x�qm�5B��(
}�q�u����\�.j=R��/sƼ<�����mM�;z�43��ϟU��`�V��-dL�QG%�i֍�Fy�n֮;.y�&��N�t�l���ü��VV����w��+�i�wy���f�,�,�U'ҫ1�a�]�z�tk�9�ߝ-}~����5>�C��x^)1�oj{I!tG�),�N!T�˄+�?M���=_���ޝ�V����@u�\���kG��sq�%I/9��([����}W�QȞ�*X�7�����(q�|īg l���쥚�	J�h�V=�kO�{4�8��fpG�������{�ϲq�Q�$�R*����f+�s�qE�KFIk�������������¬{���`���{�t�����������	��J[_{���?!��򷷽yn��D���`��=��I,�u6��q�o�}D�oQ5��_O�����Ik�~�^u�wz]O�w�{��>�]����$�39(�Yy�� �7�.V]����.���#8�;�>��f��tW�{�����'����p������ϼ]� {gc��ׯ��c)�]c�\u�vj�)�.ݤ����X4&��P��*,�"�b�M�r�4�[���ʛ�y���bai�z��lz{1Y!K�++˞�ƷN�ϲh���cѱ3���((���Hݒ��h��b�E�捥�{�{p��z�P�����ҫ'���s�ru�[ x����ڿ�l1z�wqל��L��t� R�����2���K)�^O�~���v艿*t�KN=j75�����U�i
n�i��b1&_�����_��1fo�{*vK�0�2�/z�B3����L�����C�ܟ�͗gpU�o8�#����e�ľ�}���]�/�\�֗����O�*��>9�	�{05C��A�Bl׍(�5h]ث
3D=�]R�K��}w�κ�w�un>[���ӻ.�tg���c�Q�vm�5�j��P�ܪ��'�6b����;���cs�&;.�0��C��9u֨Ŗ��D�9�˴�����9|�؋�u7�=��75֮z殼����&��en��K����}�_	xk����Y׶�c���8�M8�f��%�z�Ĉ�l��%�u��B �}�ڬ���+'r�u[T��+��y	rpr��s��{x��qgv��S��ou���ʹ�,�;����M�S%6�,=�_�g/�ίoh�ϛ��A��fh��Ɩ��o�8���){���NM�S�oj�����6O-ʼ��}f*0�� NK+�o��gMh�e��s|&�C�!U��-��q^�c�<c��"q�f�7����UB<��zܐD�G��Җg���\�{c�,��H��s@ref�}񗐟/|����-��.�� N��=��&�մ
�E�!(�}~ǵĺT��M�Au6����:к����1�8\�j�"2��TŅ쯽gy5�w6��'rB��M��4��*���"=��f��;��oQ�k!y�kN얐�B�V��C��}Ì�:�EQ�>a-���/;������I���"Lʓ��^�nnv��+#}��p��ŋ=c�ew�-99L�":��m���;WaqkU��C�8�4�d�6y��*�'V<����Q�|�n7����s&}WI{$�o��	�!�x�[�{����*�;�(ӊ��$S�[u�z ����=u��*e!Z�6����wwٓ{�����2<8�=�I�$m�0̻}'������eދ]gg�J�'ޮ`�5g秮=�-�����y���&�f�.\ǧ"���A��8�w�Ǘe��a�%���4���k܅�#� �)�4���>�=kgpg��U�ba���~�V]d׽'{|}�*Qi�!��&����߮Es�Vo�����>)�zdbz�Ǫ���V�"�D�4�2�x�����:{_M�FD�>>�|��:��]������_Z�8V��aN�µ�#"rvo��������G�׹!"󟬺�W��nc}����0��B��]��W>��ݬ�8k~5��ZH���6}�(㲲V�Wu���ܱ7�~�*kI��3��j�b0c��1ԧ�Y�{m[�pl8�e�}�ȉ[�}�|��۲jR�%qP��;7�)n�7���vό�`�
xƮ,7���wG~���[�I�ɢ ����m�n9��hN���l��7��=�x�3����ʯ<d�WR���¿�5�4��*k ��H ��T"Q�W"�.Y���}vX�:��X��tn�b��;{q��I��%��ѱn8v�n1`p�&O�3�mʡ;
����9Ӝ���]=�Z�k�6��n�Z^;GF�{<�P��Ɏ*v�׬��N�Q�$����ߦ��r�$&�8�c�R}��{O잿[���Ʈbb����g�vc�+m�XOwe��j��hf�y���ū��%�ɖ�}����h�S��'T�_��b>_CB;�)�~	�f-� ��t���»�4��]ko��D9'�}�S��mn�L������=>散%�T���ܘ3�l��ޝ����u�(��S3�o'�{oY�2�N�5�M8���>[�fw���=�v�{�1�ң�R:?��TCO�O9IK�os�z�� �1�M߾ϛ�n��NE�����DWb���f\TR'ݵ��u�{^y��}x�ma����k���Gh����-�Q�M��j�A�rD� V0É��`m�pO_�\���T�e�9qט�����|�����s3�5Qg���|���}�����������&�t{S$�9��xW�'�OܟVj�Ĥ�:�lI�c�c� 0�����^�3/e|W�Hd��$�W^�.�W�5�������v�ڛ�G�t�1ʟd_���5�'1�{*��RW/c
�{2d�|��G�w�N�NC��N���<Xh`�bN�Zmh�K��=�u^,b����g�����\�5���]�Gc�(�3{�v�ΰ�m22�M��_υ'yG��q�ͅG�'eH�̧�|B﵌5R�,�/'y�������r=bd�vF��I��	c!j���]�Ϲ��ɼz�������[܇��'��^|r�F<W���z�n��]O��V�ٯ3C�uek���4�Ĵ�_r&��	�p��N+�}�5��	��t���uTB��� P�©;h_�`"�Q����q�����D���ǔ�BMp��A��^B�H�2�oO��@�MD�)2�պ�(v�v��V"7|4fN|�za���V�S����u<��U^Y|�S��ӽ|�W]"9�lɵ~9�oFs�:+{�I�'���3�L�D�C�}�)�����sm�͵rN򹷖�ض^G�t��,�Ň��k��|�n�����m�˧$E�d����>��qV�ʛ�t��:6M�¤�dc�[�
�ĞU���Z�D�wǇ�E#	��)7�ה)�=2�R��~��#L:3�E�.z���W���R�l�����W!8�xV��g�e������"���{h�V}�0V��@�{�k&n�����ώy��9:�1�Md\�+̂� ����}��]�Rt눃]�נ�� 5���ݧn<�ٱs�����d�4�"�r�~/6Jbʹyu��7��G�6�:��{�ٖ��^-*0���
Ć������7F����C�Y��`�幽�X���t鹋1�������A����w��-��P���4�E�Hfv�}��q�el�ۗ�V�x�����N��u�79ei�,gp��2�Ab��x��k��n���TlE�z�D5�hJ+*3�/�`+���C��a�i�n�I�P�]�Cx+rl�zV�qe��)3�{Gb�w�mnA��.���P�D`E�
؍Br'.�l����O;��;k|�tq��YLś9s���8&��Z�Wbգ�ۗc۱.�j㽌�.i��i��'*�ˡ -f�w��kU�k����������5����\��ǵf�][/��aV;X���JAkxv�)ܛ�E���w-z�r&�R��;oU�2����h,h�ٕܷj�vK.e�4n��� ��W�� ����J�+TK���3�h��;x�W��/;�h��B�U�Nh�9!ھ���eJ��U�ҷ(��3�[�gy(��fE�s����=Z'>�V&�,���W�\}�`�P=)�fhe$�'��
�)D����������3$��~AV�1�Z�C#pj^�;���)na�;ofT�:�knŷb�l����/Nvޞ���u��Ѯ]�՝�{�XX�k�P�밠�����9Owye��5�f!�N���I��H�����S���ۗݢ�����-<��E���L����x�U�[�22��nc�"���:C�6�Eb��R"l��w'�{�|���f��2:��[�$O�_�¾����c?\;��_�y3u�P����<���57�����#�i��v�ځ�������#����?h��~3>ri�A}����0��W����t��3�#H�<k����
�j���!L\�=�}oWOyV�ՅV����v4�'��F�*�ݗq%s���̘�u��Z���q����b(�opY�p϶i\�2���~���y3��j||��e�\)�դ_o���NP��u9�4~�K�V ��.��rD�+�K ��H�`�
t�7{޽��>`��D�6榫�?B��{޽��d��z���k�O�ؖ���S���먎�*�<�UMT��]� cn�i����ʇ�U�&Y_��R�_�"?-�`m@UU��n��E�?)(������S����C����;� �b�=s�1�����ʤ�j�v��_+�ZH��kt�W(�pPz�)�k�ݫ���ې���F�Ѱ��휼�6G���{w���r�����v�T�	����ŉ���f���y�\ˇ�٤u�FD-�tr�>���To
�ʶL7[e\�xȲw;њ�{��6�nD��=X�v"��o���LA��Q����Ä� S�	Bw�x�<):ng��f�܋8�3^�Ro�^P��0ߎիyA琢+"�S8+��y�l�������?y[Zs��g�l2�o}����&�R?�����Jmֳ�Z��{\��u�qcb��p�;=Eo�/�K�X�Uip}��L�W��y�߄w(�_u�Yf���N�ާ�;��D/r�o���� �%�||}-��\�3SURv����b���� !��=�ɬ���ũ�z�"���=���mmq�����zsCvgE��E%���Tx��m3��,� �����R}>�̘4�C&�I8*w�׽?Q��'P�,�����':*�����:�a3Cݒ;I}���=��䜻�nW�S���g`Q�=<��Ӿ��{'�7�Y�k�gm+���㱀<���{g�²$�u<�<�ݞ�߾�g�+*��"M_;�.>纩�s&s~����;����A���/?*�ʞ�čӕ=u77�*���!�[,����Z��X�_�c��%挞�:��>����N��ឺ� �$F�j�Q���nٸ�!Ё&�7������Dh���G���ݹb��5^f���^?^�\���n�$����;��x��Y��ܽu����Z��B��3����x۾b�g5�˷�s����ni��)A�4#�������c#vр�n=��l-pQr����r�m��u��-�r]:mݷ9\9����������8vm�sxܷm�tnX��+�<�zi��rko\]��zA���v��[���콕M��;��Tc{9[�C�Ŵn����5�<��7:�;�ֲ�1�ݰ�\���[鞳����<Pwk��^ݸS�jI�j�I�H䳍�\�^��8y^���9�^/\M1�?���T�yL��G4}�ٜ��HF�����Q�/��YIL�G{�7Z��#=�y<�L�;�L��� �w�u���j5�We1]�=���DP�e&!��7xaT\Щ�����ے��܇B6u�<���,�;q�ͩw2�_X?����N�X��+���b����ځ��W��k\���1��pa�i$a?U�:�`�=LF��dY�?:?d���~uDmb�ڪ�߱ݑ���r����&�=q�A�?Y�WO���;����!�܁'V�o5��c�ټCH��7�}N�ut�T�
z��>��ݺ"��mrs^�'DP:^@���߇3;��F�y���5�d�Ψ�1�K�j�fZ��S9sֹг���n�@�N�A��´���#cP����s�ȝu�~wW�f�LNoc2+���S�׊�����0�0��t��\�mf{v6�Ԙ�oN���q�&wv�\��/�0v�+F԰Y�fz+�9���ڮ��[�0eS����٦)t�����G���3�;����k�(Ml��l��̄D�w�M.�<bv�F��%�
K@�h��Ͼ��5_�4�����d�Y�˩�>�C�(��S4�J7�(h�{=����=ܼv�.�{�%o���kjZWw������#{Q5o�&��u�X@7��oC��R&*f<3�/t�7� j�	y	�^�Sgj)�U�^��Y��~n���!�<B7횱!`��I/�~g�ͭ."P����N�s�/���L'�<h9��iW1�ٝX����ݯ�ө�5�f��Q��X���gJ�~U����a��r�������`��#G
���	��#=��
�y�ˋ�k|w���c+Q�g��#Tϼ�Ew�z�����%�D����oϖ[��㥄���W_�f������,�p�)}�/>^p���~ڃ߄��|�����L��Bc�z��b��MF�=�z#'��T+n�����3���ζ���½n[nϓj^ua����.V�pa����l����)���S����em}��®i�c��Mg? ~�$�+gHu�bK��̯�]��}�CV�uԋ���C�0ğp�jFE��(�Р���g�@���{V-}�Ǌ��&��s�O_tv�[�[�= F�����<�G�[�g� a��=��Ӑ��t�3ϳ��ș6/o��=9*pwfOn�/G
�b�۹s�9���g�eR�}quT�Ժpv#5�t�;=���xGtkF<��>���fcܝ�3��N���j�LHI��t�{wK��Q�`�zQP:;��6�K�ҿd�Y�^\i�ch{�/�+�w�T�#�=+ë�w�����
O}�W[ἣ��iMX��(P{�q���~Z�ڮ�NS�W��&qN挊K���W���n�]E��<��.��/WNޣ�~X?{ԙ�Y�Lms�c��e��<s�G���Fp���m��4,�\�&�_�ǖF($l��������=��q�������4���������{�֢��R
<�M�`��q��l�J"�	�����0}��s��3ikpeɯ7��R��+�K�Ȣm
�� �ӄRP�����kwE�w1��S�5�������=������7�
�{n�D��Ksb���UU�O^���-��uvx4`��G��EI�..N䐮=f$����`�>0�mVx��}�hS����������~.{%͋�q�ђ��71Pz!U�����3y���ץ\2�`��i����!&� ̘\�]��ńI��{ȚT��v��w�˳��G�N�^���y?'>ʗ5ԼD͊��Q�G���x�d�~�i����Ю�;շ;�~���>��0l@��^u�c���N�s.��KJ��c�I�i�a��/���޵�K|<�W�ô��Y���{j�N�苊�h;b��^��e�ffh�u7Ok9�u蒚ۧh��k���K��B�[���*Sswcr�����]
d��z����Fۂ?@.51^k3�~�ӟ��v���򴓙���߶!�F��V'{��v�¶�Ҩg�ξ8of���Jp~1�"�d<�)��u���g���l�hG�����2���p�e(�u`pd���b�.�$���'�n߽���;���<���XfH�����YC���26��E����[�/��5g�8w�Ni�붾�"V��6[�1�i���,���%�|3�-1uD�9#G�#�r�c�*�"%I|�h��s���#r�B������&�����N�VR�r[Ւ$_��ȃ�ꌆ�S�+ Q�]��u�VQ�n�)�,�\c��q����}��߅��e/�Y,
�?+�ҍ8%=�ۃYѺq��%���\@���4,�{+�:h�u\�\��,4�j!��M���%�^Gxt�*���|'�hIzNy��ϣ=�$��Z�J�����T~��c���:����Z�l�f��"�S^�a'����0Z�b�Kr�xx�'������ۙ���A��O�9�|�z��X��G���]ݢ�Ќ�C��]WF��<x2&`2����
��0�Vo�)_�����?���`����sn7i�����ںM�nr7s���賢���rS=�v���ب<u���{�7fڳn��Cv��V���܌)%����dqR@���
q�
 [&IUp�e�@!���4��ۣ�M���ѐq�mڋ�m��<�(�VZ�vе��eQ�z��]nlG;&4��;z����A�,�:�BF�C��md6:Q.-6��r/��6k�W	��68]�N-옮��x��.�����p��Нh�sf^R��n��v	�n�^CZ��Q��炢��.!�#���W���[v"7g��ͫ��z���60�dv�P@2�H�c�#h�W�ߧ�O�޿q�ɎÃ�-�|j>Y��}�c"�x%��~�f*9;o�u>���+%�5q{U8���LZ��0�	COo�v�N}I\}�*�9�"O�󻋇�{�)(`߭~�D���g��IW�8����@��wuf�7��2!S�������w�ȋT	��K��Go?1�3��,�8���dHr���0g�2�'�w5��K^k�+��f�؈���P1?bZ=����ϳv���@nݨt$��e���іG�nv6�f�O���UK����������7'W���ss��`/����f`ꭨ���U�SHQw��umN(گa�8y�v�������鼲6J_um��<�y�~r�<�k�)���V���U�	��**��Dʶ,��jܠ�dgwp��=��PJ�jw곃�$�&�n�C��-&^N�4��޸�V�W<u�?ZN�AGT-��K�d�w�3��%���uR���C��w��N��w[��3��1��2bK�u|`�]G�T�S�o�|@��8�g�1I��,�IC�h�ܚSX\��7�����Gܣhp��Y9��r�����S98;nΚs��-�!fU�ǬD�'�*�Ƿ9�*�^�q\w62f�NS|�ڣ[�3�S�����oɡ��ҖT���Efp��.X	u猷�����y��ׄ�Nap�v����T ����H]���C�9�H�0�]1�|H~A<��~��7g����ة�g�s�F�����ȥ86"���~"�q%hHn���kAj��~��ړ��W��������L���GJ"O���x�}��;%x�:�`�<a�AO/;�=1gO�̞sO��
P6�撮���?Gb'���C��n��){B�DE�qn����6�E��-��Ä#�S1�_S��P�*�M�=�nE��޹�j��E^+��q��i�.��ý#6z�y��i�x���,~@_�V�$�oM��D$�^x�t��)�\�j�n��..�{n�t݈M�QX٠�v8V&RZ!(�k��%QI�&鰯P��8wM7>�{.��ea��Ҵ^Kɥƺ�[�mg�O�)&��7D��O����>K�h�K7lr��I��pb"I��^�UU0����ʭ��Q+�z+�D�f���wb��I�Cv���'�e/ws˿���S�3� �g�~�f�����۔V�V)�	�vm�4G���vo{<Zdn��E_|B�"A��t�����*���$7Z&@���Y���Ab�Y�]�L����Z�0��0X��L�Շ3Y���u΋�\�6�Ʈ�ѧ��i��@�K�˨�������aE�)ؒ�G�6�!
%��0,��O=�s�j���ۧ��)��f�i���=x��L#i�N�<�(�~Եz�Y��#�/�8�k�(u.s������*W��}$?wT|撃���d���ݚ(ekɔ���;�w��^��D�W0�^������x�L����YD�[���p5J́$d�s��l� ��Y��K�on;�������|}��^@)r�f�v�i�}���#��Mi��0p�Xb#�d�J:.f'q�qf�w������݉��/��5��{��T+ZjF��Ty@�]t˟+΃�xV��Kق^uk��@ُ]F���y��ڃp�q��}�\ϯ�׍�|)c#6��#�]�i;�WJ~���ՄV�\�/(^��m|$����x�,�Mk� C�U�tX�����3�o�n�4`Kp�/��a�J=��" ˥]�}����}u�,���R.!��C�]O��~Ɂ}ްf�VӋ�~�쬚c��Qa�_��E.Q��bM�6~�B�V*������ߤ���Le���-���$|ʷHozF(���=�ɲڮ�S�Ѫ�޵�"��V ]�[xג[e���;���xh��~fmm�+Z��K����*�x�����Su��V
�D��T�]8p�Y0y����w|���g���,�|���Em��ڜ홆��T?ȫ*���B��u5\^�[���x��No�VY�������WE]6+ݘ�K�fvت��5=޼���;Ʈ�WRG`��=��~8���q�H�6v�����Vi�C���6�@�Ѫ;aDo%�p#��&0p��m���Cb\d��Vr�����p��ws����Q��P�Nչ�j"�fG.�0��UX�P��A�e�������m2��r_9"��wS�����s���dh�(�u�Y���
�5�3�s��ia��gŉEM�
ߙ��]q�B<�4��J��'E8��-�\ #G�]}���D@n� ���J�J�ǝ�-8���mѳLmP�D#nshP���d��[<����d����E���F�z�����L�g��	����G���l&���2#`N��-^��\H�"��^T�X��c`Q�ɍ���c�?c�O�'�[{Ҷ+/@��3���Lx�^�C�r��i�>^r��s�
<[,T�I�mNE_d�殝z}��~6PW���
�aT{���*��(�^+j]B'�+/����d�N��J3sW��ϙ�T|����t�E ��
2Lԉ�"�|I�י ۠�QH�s���R�6�׺����Pv;O(�!:���:��x��7�ܥ��U��3z���f��&�:cb�ذw�u�]I��t�n��1�=r'�X� ���Yk&�U�:�>��e���wYnTK��t�0�i`�YD�5�W��u��6�l����z�ฯ��۟�s������M]��2v�D�J�ں麙�4xq{�w]��xnNx�U�y��۶��������L�_m<��S���A�b5Jd���}�ٓ%���r��u�rs�EU�!oaG46D�Dr��Y��پb|l�f;�o__�;L7/�͜+Oziy�]���'o�;AC{����LmW}��Y�\���C�`�3iݤ�R묜�ZN��uk�����3�6Q��b�K�U�ٰ���f�����6:+���r��0�Ǣo �7_n�;$C(���G��m%i���d���a��n��3d�V����&_�3l��=o�unr���_��a���aJ��:赥m�'M?�^�k��vܽ�J��bUs	���O˅�12��۷�n1�9`���	��"��m�:�pw%�4�p�33��CAY$�5�����a��C3o!o*���s�>����t��=yvc��j�¶��Ȳ�p���'J����A��l�� ����O?�T�)�"��Ǖ2t�����m鬫�h���ۼn��HWB�il+@9!�9���>��_M�E�wF�e��ucj��r��B7hz%�rA�������&�1[f�iޜɰ."��l��y�;���؍�Lq�"�������a~�yͮq'7j�v�u�tB��m����۝m�f�l�8;]c�N�=ձuY�K��ײV"콣�@c���8�%v�vE�T'Iդ��m�A�� �����~��� �׋�7n�lq�sq����1�r��6:�1�����{a�F��gM��=�(�n�\�jW��C�9�SS�r(��aL��띧v��lͳ����[`ۃ�Q QJ(��i��"��8"v{M�^U�κܝ9n���&�V����q�tg,q���O�cn<\���� ���4�s���g͊�t��yp�nŋ���������_O�cֲ�۳�=���2�jk±�qV�ڣ_F#�[��]c�?o]�|�݌�\�<���\X^ɸ5�� ��i��,Pn�G���B7u�^ec�����F�q��$;wn��u�;v����,�[�n��Ͱ�p��h��=�H܂̤
�[a.�~딺�EM藺NL���n����i��un�j�PǣuRq��7��7\�W�/.��������Azm������}�~�ڣ�����p��v��{9�c�7��gE��Dv���Xy�I�����;�^8Ǿu���d��-��=�q�Y��~���?r�NB�vkkԒ�]�U%[��n���9����/&��~��i���.X-�������g��P�h����݁�n8�m�K�W�m�r�e�»{��v{f7<�����F�r�eM����D7k=��v�͞����)s�z�-��0�Ye�����'6LG���<��r�����6� �%�a�G4�:Yw-�������w����|��v������O;g?v��|n���a�Pr
��.	�@M�XL����/q�V�H<Y66袴'c2�7.��7ot[l�d���÷Zֹ|M���������1�WѰ�{n���͎�t�hNzZ��������zޫe�lUrՎ������e�<����ua�xZ��j݇f�]<���Ƿ��m��t����ɤd��U�h-��c��a݈w[��NGN��c;Y��mrKsZ�=q�Sd��퇧��!�y��u�����I�N�ݔW�\��?��m��c�ڬg���qh;\y��<Uf�g��t�*rm�Ƀê6�m�:�V��uis+�@���PD�!���aP8�mݶ��rۙ��-AK�#����^}�c�|}���f�\�Gy�T ��_$�'Z�l�&>X��
��3�9"��u�us(ϊ.G��%��e矤Tx���<�]�v���nA4�}&�"+���wC1��=`���U���c�u�O»�	�Ʀb��MX�#hd�<�.mZ������:9�X�D�n8f
nD�'2�2>�ș��+���'ޡ�H�Z���F�����eR�=�c��[��%���\m	��rUc�ȻG���D�]��U�^S;L�ܺ��,GBJ��h��MD�(ۜs�`mo�F��*v�z���}�&�W���~W=�F��u�y{����F�w�7�w���ư����ĵ�y���I�u��\QH��$�@xJ]�3�?|5z(3��7&��9���'����ӆ�-u�~^�z�z�-��F�T���$���ȑ���k����$�31�|Ѐpzvr��I��^a0�îB�8�N��T���Ǯd*<ݐ��y�.tYu�X�-U��R�}ߦ3s���}f��s�W�����)(l*�:}3�(�����d.�^�v�� X�wU��da��~	tu��W��5��g���M�j��]XƲdLC7���X��ֲ8���٘.(�پ�S~�˕YHc��A\�R��4(7KMRΈ�ۺ��Gj�mB���4>��qXBǄg!N�i�g�/���xs��wR�u�o��sf۪#�%ø�V��H�ꀕty̑�q#���_ݎ�w�^���P0�m��!�
��ϊ���dpqe\E�g�';���.����@�,Ɇqt�j���,�NE�g��ʈq���d�?g�d�epN���*:)4�C(4�[wW�C����`�����y��[��Xk��xY�5E}�Վ}�
���ś���N<{Q>'r,�Z׫���)ً�EG�~���,�c�����zW*�^�dQ�q=�|ߦj#�]���ֱ���_�����̞���9r~��`�
?`0?�Lv�fwh4V�挣_s��!ÿ.rYS��*���l]����\V�<^�ݹ�g�9��v/m�8�����3/��9V����w�ܨ��U��У�5��x�����	�Mr���Bժ�������x������^ۛQ��QU@���B`�ওLՐ ��C�n4�U�u/.�v?x-ЊS>�'��j����v}Q��3�`LO[�~���kP��Z����?+���N%Ù�;G#�{�ވ���`��i<���s�S�蛻��ޝ��zC#e��3��͌���sh�z�k׀�����_ܫ��K'K),9���3D�І�e��kn��U�If\�oN���_ٛW0Y�0�EOH�MȾ�Q�|����o���\�a��-�{޿2�X���Vq0��B�~(Y���>�z��/�#���Д{6�z�a#>DNzM*�*2uw?x	ݜ�W��&{=VG�Q*ʦ�g��x��ƞo(��bi��|���~����FF�@&C0�\}�~�K��P��|��vR��{h����3��Q�;�/�t3�d2؋�}μg���&
S���F�D �@��to}}��Ϸ2���dS��d�rH�U��>�}��&`4�����"�.n�q�;W�2�Ȯ�	Jԕ��� ���?��s�:�3E�t���c�s��B����r��{�sy���J��9kDXZ�;k�/{l�%-ۣ���/���Vp��]���N��[�8�~�>&�h8���}u�%)}����9Z�'S��������T&[�7 �G�f4���7�}�,��oۗ�x�������h���C����P���.�{�E��'�����2��M�w\ƹZ��}T �sn���|�t�F!TS���y&��������DI��x����q�di�L�^��������g�n���t��]eMs@ˀ��{=_�
f\����v&~�j4��f�TZ=q(��0�Yr�uN�f�I�wr��.i:q�;�<�}|��⤏# ׇG:�_p�!.��m�\v�v kKI����ӑG��~bF����o�@B-�)��ѳ��)�a~��{��Bb��z>f4>W�2S�3��o��+ڽ0=C���eYf�a��{?Y�|��.����Ul���5�ڳҢlI�a[H&Hj�=lIɬ���nv�ڕzY�;BcɁ2�vQ��Z)�q�P��K��f��sQQ�2&{b��?x�����u�oh�5F����x�>؛rC,�
#Hgŗ5[:nw�u��F%�4+$��D�D��h�xi��Z���l�髽��j�3�9	�Ϩ�F<�/+g����op�ٌ4w{w'g}���DI �P���=Qq���3��)A��#ހ��C�����		2Sj˕��/�Ǖ#�U��D���U�)�*�û�ٮ�\]{�e�W�dm7B��zeoEȚ�>�.5��@��I�|���*�th6D\i�������F���7i�|��|�O�����V����T����,5����R>���٭:���̋	�1�����[7l�Z8�Ns���l1�ME�7���\�����>��rt�� ؟f{u��@�}ף�sY|l}���(IS�ʺ��޶|.P��p�N�3w�XxŦ'}"l�[yיx,��hܾ�N�a���d��5�L��n��1�}-������U��;�-�$��&曲�c������t�qr\��l�>.����Fjv���M�L~�6�qb�����6��۶�;���Ɠnx�d��f���lv�q�7t۞9��%r�]h�=q���RV�e�����x;��Ip�[i��y#��ӑ��*K���}���)�:�nB,v���;��ѶX����㶶����>�ocP�m�7a8h��]��i��i�f䊹�T�NW�Ѳ�c��/pzڞ躗:���c�)>�&f`�����k�y'6�8��]��+���z���Փu^�>�'zO(�>��7�I2~���˵�MG_�խk�����JZW{p×�1@鏘4�����pO�XF�Y�{ÞT\Q�O�hܜ��Ӈ�|Q��Y��[�O�O*��ݥ� �<�)�-?
����uh3�Ǉ�0N-&+�#�#���7�S��<G����E *|���r/���|�w�Ć�v��ۉ�j�р�('�q]BE8��$��z��@PH��PQI{·6�(|��O���+�q��7?S˒&��<�דp����S��^�Ə����ގ��H�9�7����ל�ˏUlDF����8�ڿ<C?'Y��~�O�zZ'*$T���ʬ}楸���D-��k�@����2����o4Z1��BS����W�*�Qj�Yd����6��b5QƵ�#��뭾�:�P�c�!K�A�n�M�Y],�r��'c3�"��fWz<˾�#8υ%���a����ࠕdn�Ͼ�&�u�ѹ�W��
 Ӫ�$^�g�:�����[�7b�9�gO|�B~�:)"!Ag=&����{n=?#Y=ڻc�/ޱ�R�ۚ�H+�K�⺛n�������7��/6�e��'x�Xi��{�/�nt����3�o���1*��:<���r���U57θ�@g�lIaT�9v�r��eچ����E���/��":��_�.w�C�����=�tг���n���u�_yǶ(�ҳ�����h���߷ ܋���c��7z�A>�+�	p;��������f�6�^�}�7cnTA��J�CKz����3�VL�*z�]m�/"��_�U�v��y�*�/�~�*W��߻��x��i�=Ϊ^��Od�&���~=>�+������� W%1ǺG\����!�;���#my�}������b��"�b��w�ޒR�#_�|T���'5���`�r�������J��v�mv��V�`e{v�1m��8-Ə�S��<\kuݢ��	��n���"Q>�5�oﹾx�]�ZNK�7z��udM@%&�P�����=_G�F���$�
|��Y�����LO����3s��.�$���I��z#�*�"��|Ϙ��}���:x��q����~����xfDa��͗C��w�y�/�~�JT��vv�^(C7���ϛ��v=�}��2�!d�`Gu[����6��NY��6#T��j�3|*}��X���g]h�0ߊ׈�K�_EWi��S��j�k$r�JT2�����a�ndB5� ���H�~��+a��ExR�s[+�W_���on����$TW�>4���Q�^w�k(J�r�A�F������RN��%����wZf����I�'��{���[�4�o���K����#Ԓ�jLxwt̬[y��F�2�zj���}�>�蛉@,U9)G���L""��ݞ�{�0e��d{�]����|�o�rպ0��mo7�� dr1*ONzbp�y�'�G�N�Nל~��9�r��ܢ�ֆ�)S*��6����Sl旙N\NMa.��qvov{H�iΐ�᤟v�{EPuK�\�S�F���ڨrA��t���G�09D�X��!��,���w��V,أ��Q�DO�u�3�(ߥ{�]�����#��1s��s?g5�I_�eF�)g=t�ώf"�ۃ+�5<\��z�^.��c�6�P�&}�¥X#�ȫg��b�;��e��TX�.�	���ܷ��qI��m��z������x�ݝ�V9����O��Y�ep�0�����l�{��Dd��m��;3��n%�qH�|1�JPbn_,��]%�}`�O��LOz����Dyކ��gz��U.{q1}9nxd+��+پ��eQ����`τ^�o�s�^��3;}�[E�j�x����)m������f�E���v�40�E�^���w���-VY�n�.�}�Κr����!)�!H�����8���v9����1�H8�m�ܲ���a����s>|=5��4h�'t���`���B��t�����LC;�Ǽ���QbL�1�7;�c�S�����z�P�d��!��¸6�`�g;̎#6:��`�٫��N��엪����UU7"��n�NL�����b�#e��u_z�n7-C����b�>�����q��b�Xc\x����"�AM8dęr�H�h[{W�h{���2���$���ά�#X�W���'��=4�뺥#������=Cñ���J���D5�]C03�j��7�"��I�IP�g;2��bLn����7_ۿ���EK�IH�g�K�}��cQgz���+��Ue-o�j t��v�kqu.��{���@ ��(�)�uy�g��#[���2v��av/3���f�ݺuP_y��oc�Ϝ�b�'�=>�*N���>�,�}ҝf̺�����YuR!�٥���U���p���s1�zЁ {.��X[;�����9<�w9D��4��q��67UQ���]��eˌ��"w�bh���US�Y^��Ҟ�f$�1��Y������[J̲��쬉�����V�!�Ř����;{\��W'۽*��=\��i\��q�H�y��<�h���$�̫&K$
 <��7Q�#Z�B	/Ccv���U;�[�zy��U��ۋ�c�ڧ!=!r{��=g����� ���g��͞V�l��&w��6��dۮx�\�m��KŞ��{�s���W��?��w�\��8��Ȼ����"d�(n�AU�딝��/�|h�{f��\���8v0��<p�+uk\�5�j���v���� ����w�
���Y+ff�{]���:r��v��ک{Am�P��؅�Bə]�+�w�<�U}qγz;D}4�GQ�1�H!��7-!�]TrhY~��e]�X��a_�N�}�,�7[\�}����-��b�o�^��<��t��!��q�Q�q�<��č�0�B�*�=��t'Ըх7�;��J�������ߜϳ\!>����Dؠ�����w���Y؉�2oC�=%j�<[o��5��R����~��o}�)_d�Eu�9������\�D(�V��7w}�T/�Jm�J��������UN���gFp�<A��ՏבM�+������t����ށ�?��}���ѷ繾w�C�qDr���9��D�^�IM��T���8��lY�	�IW6B.e��=r�a�Ӽ��+����lY��GTr�u>2������9';��3�5f�� Z0��y�����%�)�7���\�s޴�1��ѝ����M��W�k&Uש�6-Ԏ�+�i84�b�����q��Й
�}�s&���Ƨ�liZǳDTꮻ�N�:��*oy�����eC��b*��S�#�Wb~@�!��R�$G�m����	&Ro<<G�nU���yW�nc�F��t!�1l��������衕n(9vݽ�\/��%�Y��g=x�2w�S��G��ڼRVV��U��:�ǟ/��>��v'�X�l��������n�d��̱�_e�����}Q�q�{���c``HCe�a��6��!���<-����'�tz��������+9��L.��'�7~��Gg�&4cZ�v���j�"o)�"�#�:����a���
ZgZN�[�
�����]��:���ʟ��}�c���	�kw��O�VC1}K��3:�{%u2/��`[ϴ'��g߅+,!-�zώS�_�2e��~���P$��U)�s'��+9s�"C@/gk��`a�T�pfwd��<�4YgM��g:�}��b$��ģ#������Ӷ��ne!��gN���*v���,Wl�"UP��HHP���w:�9�5��:n]g�"�S����""g2ܾ�e�"�!0s�E�(7��5~�@U'&aL	�}�j�y�p^��f�f����5-�ED��܁��G�5�C��}�O�Uw�`��n��ޔO�Mf�}����|Y��n��cC�d��tW�'{��o�;�j&�׻�RDX���"6BmA$�������?��P|�bb�	t��v�k��'gG�=ps�7����X{���ᳱd���2P���i%���O6��-�D�E�0���蜍I�e�ئ����eX�K�{9�\1]D\s��%سw�u+;ب�ޒ���Ǩ�8�e8.��֪c���v�c<I����f~���]��M����g�y�3����L�����(�뷆����Z����>�A�D�ȅ�t'qH��g�l$�hB�]Y0��:�m�w��pc;ɭ<$�ohE"�DmG�K���X�6��M�ַ�X����2�����J�3��f-����p�71��a�q�Z�.��0\X�]�4Z�N���)e3�N�7�ۄ�I�4.5�[陖!=�x�z�^���[����k��X��fwX�?��s�m�U�/�P�{�\���(U/�!v*n�i���z�*��h7�|�!�iA��`f-(��n�Xs�f����TZvWv�-�w� �@�[�p�vou8^B#
K��)�C�P�`�u�@q@v�G)�V�҇���^�C��Q�>"�m3�)E�0�%���O�s�z�I���@ʝK�m�1�"і��,��ݲ���}�h�#E�V��Wp�:�%��]��$���l���n�5�js2��I$���4�M�oX�jT��c����T��*���}����KIZ��=ˬ�,���uթ��]}��˛Y�Q�w������y��ȶs�՗ ��{f���%��WY���.q����>�:�[��Le�uBo�h���qc�n�`	���U^��9�㐀ϭ�m3u��ET}�S��&B�{�0����B7`��ٓ��O���I�VFļ�3����QɁCh���&��^_1z�BH���"�F4�Q�a��<�͊����Yf��S�s���r!.��AL�6��ldȢ(��_�=R�ޚw�K��x�U�n��}��0�V]�~ucRw��@n��_}�"��=ت&�_-�Fq��k}2a&�`��ts�Ds�z��ԇgC�KJ�!y�Fjq� P	buJ+ .7 �(����K�mP&�tԩ��n�*���:.������#���߫�U%Yr�[ǈ�
��*���-��I͵��"ƾ���KeK*�N��>��Ѳ(���,Y}<����c$��I��}|j�~�xն��|���%�LI|4[@��<*���L�������{��.�j.��uvNRJ�
zԺ*����.�6 Q��{�����x�]a�*��f!2�ۨ؏C2��w�'���E��ZG�RBuj��%"�	6[OՆ�&Zy{ڞy\�>�J�����!���߾=�,od>�?_��Q�J�ql�\s����h�{����� ��H�hηj\���+2[W6��i�Դ�M+l�<7v`�`���O���$�X�����е�	��$��,���7�{�մ���]��;DY��^�k{�b;�s+�L�k`9گwuk�
maG�dF����\W5tE�˛`��z&�*Fy]�!|x�Hs����v���o'� �'�<�mZ`޸��aan<'K
�A!Tb�Xَ�E��a���3z�����/���_5��W�+}�~�R�a��fytu<�ܯ�x����)�9��f=]�p���J�2�ޑg�%�$�,����>9&h��]^����{ʺO�ނ�W�����N#�L��ń�S)e>u�����D}�>]v=�\��C��h�w�:�Vl0�LCl�)Q%K�u�Œ���qU)�]��o}���}T؃�7t�C���;��ۦ���h���t'�F��"2)@$��+�����"�~��k�����%��&10��qt�a�oշ��e��>����<0��\��6!�G�TMF�oz/3`�sS���d��v"\������~���wn���Rl���)^��)2�_pq�]id�5P����/�t۵�'�Ȏ�Y�D�z�U�Uqujwz_��(J>ǵ��H4��ܗ��f�.v2�Ƈ�Z�WC��I��Ձ���\�����Ѭ����/y��]»���r��ycSf�ܻ�>~��uɆ[,�d$�H�JZ��G��)1s��~v���>.�)����{�NܗN+q;�aKr����r�i���vw�����۶��.1�&:�:V���Q2+���я�Q�k�j=.M��2]T�Lm�uM�kv���x�{K�9g�ۭ� �;����g��Ѿ���7:�nƍ877< �k��9g�j�9cfg{rнΞ�9u�����a7�oNn�;��s�.�u��=!!�ݮ�Xk�v�wD2dL[(4)�M��JH��*�Ǳ�w_tH!�{%W\��\�|�s�j3�yq�I��9N��/�����㬋���(����ۿ�����M���-+
p=���z�Eeߌ���]��KdGkR)��1��ə�n���gȌ���wxH�K,B!�}�SP5wo�O���yǦ���|��w��~4���B!�DC!����t�$����c�뾖$�o8���Xkr�����gw~���f�NI�D�	�%���_z�_S���s� 礕���i�MK�nD�U	��tv�q�v|4s�Ҷ��W_[��G�$�ϳ�E˙�J�����K�Py��7��6sZ�����o3y�L�����ȈC�k����IE���1��W��r@��̌�S~Vr����/I� \�>@��Ǿ�z��Oy�����o�˺��V�"�u\P���'u(���' �>*"�fq�����hk�s��#^�����n6�M�C��/�Sdۉ�1G@>������WZK���U�U�\?0�� L/9��	
��1V^�$�SV����G2b�HI�.̫q>����z$Q���,I��I��4�t�n|i�6��NM��_���p�:+l�_a.��ż�!^��K2���:�QZws8ދJP�a�c�7Sb��U!����X����oP��#���0dK��Kk����'��[���lR*���I��u��y/�{EA�s��x0�����N�Ѥ3��0q�F#���@Ê��V9�	�fe�زu�!d,�� I�1�ۛ����ȅ7�=��N�N�>3&͐A|��Ӫ�r�M�Ҩk���ei���
�G�\֦I2<�%n�P��an��t���xh��m&�ܖ�T�B@���|���#�U��j��hە�׊����b;oL�?eߞ�y>�i_���� X��Kͳ��Ϝ�-/+f����|D���og�EP�q6�0���`��zD��C7{k���7@}c�G\�2����p�\k�\s��9�=�p�	��s�ی�u�c�h��^��ɠ�����s�����K�i�O38����Q���A����}�{8Lը��T����q���������XM��D�����<�F' yf`_������X��kX\��S�B����g�#Fy�] ��8'�yŋ(��%��v��AL�D{�;3a�}��C�0�2�i����2�϶<v��G�!\l��m�~��<ou�l�7*���\�ϸ#�s�YmӦ-ًf�aZ�a�^-�Ӈ�=�vx'�|M��ٹ�o^`o'Hp�0+���c�G,�����^����N^�p���{L�k�^��L�y=߻oP�(:Z&�C{���VՖo
ܽ���F�s1eZ������7���%�3�3�~�0ϖ�;��&4j�9�r/ǳ��~����a�*�-��3{�]nzh����{Ӯ����7~��:tz�ĵn�*3������O�u����F��qR�XU�1'��5��?��'���[�eqHe����g<�)�l���e�S��nt۱�����0q��Q&�,!���ˮ��nX�M����x!x�����S�����'��xε�q����1B�&���\Hlnp���q}'� OO_+�K����!��{<Y�.~�=���iwF�E���������j�a���h{g���y�Yu���{66��ٯ�A�oN�A؀�<H�6�sFX�y�3p x�2��;wL��H����>���{�`l*c1���Q����3;��������@����-�[���<�h�V��J�a��Nv<d=S�>�Fo{�<�4���,����}��E�<���F��fX�w�u��ߓ�>���B��JڿG��:�0[���u�^CP���P]�F�jq4��[�V�R�7G]���a�[]�&���}�*wZ��_�t�6����;���B �T�2�����RĽ��W��.6����
̻�]�y�lv֓?jJe�3&�3�=츸�Dd4����ч.����+�{ƹ��D�֊�;554UBG];-N���Ƙ�x6�i�gh�+�B"�j[(����<�I�J��?����|,�pv;���-��G�w���\H��%�S�LI��㕨�rW���j��qrY�p�a��)?WzV�����F1Wg��߼�X�2�&Iy*"�c��=��s�S}^���.�=y�E%��_f������q�N3����x��>y�xϤ�0Q�&�-��=.O=�.�э�S�E8����O�)>�iwO�w������Z�~�u���|+h�e�b<��{�)~C;��s�֡4��®\�y}�i�;Ƣ�2|񽮋�����	�&7U_:���G����b��Q�T�T����J�'�ِQ�)�_&�Bfj�nˣ4�&�r���䣶�J=�U��Un�`,�­��:ߘ��v�G�R�]Zo����bP��$lq]��;��U�`أ&�[�v�T���2�0��R����&1��R׺���Hv����᪶�\<����\�p�����>�H�B(��;�G�<�-�d: ]���<Y&�<�9ɫ����Ϻlo���D��X���c�
�F�["�[3��v�C����n��;9w1p�@jH�k���t��2ύ	X%{9���j�իUm�2��O/s���'C� ��y��vT�km�;)���j0#�ܠs�g�T�&�<q���/ �v��i����i}�\�c��3у/gl�q�xc�ui���<۵
2!�6PB�Fc))�M��D8�
�������;��@>��������/y�e�T���'�{�)+�=6E��1��vw�>�Z�͚L�
Ĳ{��س��x�r�f�,�S-�0��-	�MpM����}X��N![�� o�ϼ��k'�.r.��(^f���k��1�
���̏t����軋�W�ߨ�3b)��8PV	�.[�Ϫ����FT	��1ku�0��N�!�\�����Uo�Ŝ��ޏ\>*�i���L���g�,�&�U�u���C�mH���B�Wx��h�v�Fp{���E-����r�����;��%�{lh����S麗���k.��9�s8�a�ߺ�u8	� ��H�{���/�����fx�@��VND@��g��eo��9Άy�,���6���7R��ﲃ2l�0�u�=�Ya�7��C��ˮN�qu����{U���P|5�&Ei���mхTM�!�����s5��4���?Ez:5ѷ	�����1vf�5G/{��z6�������5]>�F��V7�����;�3����*�_����������n�o'�C�,�ǕY���H촻ʲ(��`�3 ���=k2����_u��s��K��
\�_N]�9��[-�/Xs�o=�8Y+�ޕŮ�S_Q��>�~�~S��dz�}j�ʰW�{��QО�-o���T�o�`���o�9�v�^�~�v���
B�_���e�G�F{�ј#����0q{^�"&2��C�P��j�>ڣ��.�>'T�{�go��`QfHR��W�M�
	�M���˰8!)�A|�i��5���ܓ�+�3è��z �ݗ>�{�fC���v�U�P�Vʸ�W�s�P��A�ؓ>�s�Yc2����z��
KFbH��wX�����%	�*��ϼ0V73�b4��S�է>��T�:���S��
�-�:�C��y�����7[$��寖�ȜErB*(!�����u��Ӷ\�s�n�M�V搻b4�B4�#˿���(`˰l�=]��]���bM�粔��4+&㷫#u�ȯ*���D����x��ƞ�Y/F�l�f�r&�|]<���3y��%6CCP�5~��.T�	3}�s�g�j0FxB��-R$��7{ݡ����$��邩jm/zm*��A��o7��b�f����J	&-�S~���hOհ��]}7Ao�2mj6Ue)w���+^d�[��'���T�P�-?Y�s6`�(�%e�U��}F��ӽr����i7�@Zr�ܢ���*�[}�L��7;��q�������z����(��{zV_Đ����.ѝԨ�ǫ���{�?�4\�	����M}��S-��6:o;��u׈�z"N�LUz�&��GlIs�I`��U�v'�znZ3�kj,��\?<˂����|`lt�4��ܻW�ޫ�:C�yxn���S�^v���V)�ެ�P{���=.��$�c��X�!=����6d������>�Oo7���,%qI[�"$ q�u\E����;uӍ�䝩�c����͌S��$��өgK:�.�ŵy�EN@S�v=]�]O}@��g�6o�k���c|�m%~��!Z��v6Q�ί]c�vGu��	����=���.s�o�ǝ��J�y~�j_j�MV�X�K��9�?T��BUt�4b�F*3QT�
g��'g/s�N��<��5�g,��I(�؋
.Iޜ1����ys�c���G�=��Y�K��Iqw�"<��E�f��]C�7�����7���`��I	)&�D˱Dǽo��L!ｋ�[�1�Vk�/�Z�;�g�L`J�j)a�|ɬ��T�w'/嶻�*�-Fe���5܍�i�OW)ǚ�rٚl�]�Q���9Q ��B�y�wtP>4X�)��A�^.����2l��S�t�y֟`p�������0�PT(a��4b�D��V/�MN�⮑�8����ثv�m��a��7B��;��'5;�
p�.��*��<[22Ov*����>}�'���ҔV����AW�c�f�y��q�[��כ��X-p�Mۆ;p�)>嘾�詪��F/n��Q�%q��Id����M��@�G�VV;�y��ܿ�bk.�=����wn��f/.�tcf�oܳ�ػH�⊡JPG�}�l�<�A���_�μ`��b�n���QNn����i����5e=ٍ�V��t��wޝ�^��1�J�z|�c�zS�0BC������Bw�O��P^+�wX��8�"��=;y��~�}�Dl���]xp}C��;�7��ي�ݨ�5��O}�� C�#?B�:��ٯ=�^�-�]s��� �Wu���NՏ}��..��UU�o��fC:�����i.��:k��[�tN�w[oȎТ�](o�<S�EN��Zw����v�N�*Q�߯nV�f�Un���vʷ|m�y���]��zh@B��j�ܡ|i]7�~�R'�O�#�מ܎}�n���P��6���Z�-�5rf"���f�j��Y�;oY8l���gmB����t ]0t�7V��ei��m�J��;_X����s���i�$�񋴍<�^U���p�Fj�К�L��q
�
����U��:��2�[�9f���j�]弶�;5g#+��e�3�q�rӨesځ��6�P̙�h7 \�\��4\s�J�X�R�[��Xʳ�҂Kd5k5>��촄%���b�WM7��vD4��ܧZ�uȄ�]]�fh=�$��f��Ʈ�Gs�D�4� �H��Jl�v>2cE��W�oD�2�͎�9��Z2��6�IA��fG�L�_���x��F�C��u䕓���i�u_�������yNP�ߴd�ŗ�X�îѹO	��� �3��ͭZ�a4�v��B���x�����Y�짪�,�/�^2���w)Y��4
�ӧ��Q�Z��L��V�1�u����s9��\/��7o�+<�@�2��2�P0G�}8r�2��������՚E�Z%Y��V��X�R������L�0���iur�;#�M �ʒ�Ir��7|�j+X��C\(J���R������U�3�&N���fk�b�i��ET��ص�\�0����&��ؒ"U�6V��w@�8�!Zk�q��ǣ�9�Df%˰��Ļ�ꋲ��P�d�Z2.���v��+��	�-;�Ww,ʏg"roE����,�ɹ��G��s��v󛜄������u��]�J�UJf�uŽ��T�Ѱ`�3[�#m�m���.��f)��v�i�Urʧ��d�&�Ґ
۳R�dn���J�n �K:Q�79�p%���}�g\����b�$�W7���;<�x������f�w.om�5���U�s�T�����lcڀu��S�l6[j!^뺶���;k?��}獓�9��r=�烶\���JYla�uƹA�3�m��%��`�=��9h�JJ絺,��i�|Q�~v>>b��ݲ!�,ռ�]���Glc�^�)�;&��{kG��n�nut��#�s��㷢ǖ����V�W������n	��s����k�0�]l�c���8��*g��y�6�ǆ{M���g���iݹ��ڴ<���8ݲ�o]�,)�#׋o�����|v[�wY����T:���B��Z; �ۃO9�9]���/.Ԃ�v����8��H��.�N��ܲo��ɶz�
!��5=�f���w�>{w����C(QӋ{v��r�S�O��=[:z�gZ�ڻv�Y]n;<��m�w#�v�u\�����]I���ʨ\��7})�{��ǩw(��'v9^�����e5�M�'���M��
�кy�cv7>ܼ<V5�W�kC�n��c��Vڊ:�q��@�oEr"�X��*��,nŤ��u�v�����9�-�Z��E��鎲˵�v��a#.�<?ۛ�｝۞������ۢ���rnݸq1�qrs�
a�);�ٜ;��ڢX@�{=�͵��ۊw���3S���|n�`_}���1��oF�u.HW%��A�@�T�U�L��&�j,��KK�R�N��>��� ����Kn��ɘ@U�r�ۋ>�خM��"Kp�Ҧ��D0�q�dބ6[y�v�,��m��x��c����k]�cl��8U۲$�9�����pk��s3#Q�Խh�T���n[��+?��n�;�t�ml^fϷ%��-i�����n�v�s׏�N�M>�:��= ��,�Nծ	�enQ;m=�u�۴ �wa��o d����ⴀ2������ >4@�n]j����d0펞j�G	�<�ό�殣\ƹ�N:y�>��3���6�VW��oV`M�u�8�ix�CN����]u^�Ⱥ�.L'��z۰�p��7k��"9����I�\p3A�n��Em�	�pm�a��u� ��?s��B�1����=�y�	��Hb˔�(��t+�μ�>�������͓I�.��p]���4�e���tpl�d��c��U;A�X�]��L�0�l���l�0��]�S7��ӹ�b6�c���A�vc�^��xe
���mD�9�w�"��sS��9��9@V�?���v�Q�Y>�[&30���Jg0�c�Ϣ��S|5���������u�ݠ�D�M_;�U�]�c��LERO�"�ۺ��O�n�~��1������6H�0�PSj�i��y�[K�f-�{ӭV��WHoV���b�;e���qlN�#Փ(�8������)���Z?n��j#1o�wF|�;(���7�)�
^FKv��&ӭ���L�
���ٮqYtD^�]=�Z�]&Y����5c��^�{;I8Y�O{�5�ȏ�р.qv����ɚ=�h�W�:��Xȼ�14������̚�b���p5��jЫS4�5��A	��C�Mt�L��k�d7Z*:I18}�H�лHmv�z2X�\�ў��*���&���FԒ~w�)
�P�w���;��una�άs��G�>�j�����;=s��v�N�.��UFDT磺yպ8Ml�k��>�Y�O�m�m�[M(�0�n��<
f�=�ٓ�ˍB�4Y���+o�Y�7�@Y�o/�2�Ogmf9Y|�d�NjSҏ^Y���)[�c����[W�C��/�(Oa��dN����a�D�&:?}���W���FɄ^���$;/�����^�G;2<"x����z�T3{"A(-��%���뻕fhC�,�_t_fnu��GS�(�S����Ӳo���YճD�^g�\�c���i��������5ӳ}�t��f{��w�s��]$)(����̭�|=qVȐ���z�ו}g+=�f�L�@7�
�e��Q��u�/�g+nX���е���bu��(ݫT&D����}�؂�ʈ�3/=�`�*�	g%Vu���~��~���=�Ӧ��bY��W���3��|��K4�p������-���+����G�E}����Ot��p�nζ��V��&���u�g;}��3����(#C�کL����������'�FM7�z��- �J���G_^��J����~f^b�!�oc���������M����E�5s�{�˂$�K�f7�k��l���v\v�wˌ�1�E�%[;6�>���y�f�[|f5���Yx0�_���^n��}��s�Ms�o�}>W�~�|tR����K�ZE��y��w�=���G��߮}��g,�Y�~%���k͝Z�m������H(��8V�Y�L��3U��1�����`���n�t�T��Yq
�����ƾϨ��{ϻ��N�y��O�~���P�T�����!���.[�Ġy��'��K��g����UDܞD�ڣFr7˷4o������О|#J�bC;!�����m43.F�T>�N\s��E���U�К�ۄ�AA��V�v�ڳq�>�w��<&e���������4<c�wy���g+9]R��Ǯ����:o�^��a��-V㺅V��N@"+\��0B�����E<)Y\���1�B�1�T�aP�
z���Sv���@���C/�
�V)UU��Z\��u^"`��ˏo�M��{�巇L��9���W�I`����qK�f~�&������w�h��3��:^ւhS��gW��ǔW_U
X��u�+�c� c^���P�o۾�q*��Iy�ݮ���o��\�A0Rϋ�%̿}��=Ud�;��^��H����/&wd�<�=�+�U�>�b@3k�ʲ����j8Twfhm�}ȭ{:=�z������%D8'
>@���Ϧ����5>�P�k�J����^��W2(I���_2)Rq�w[��8�"u�S�e99�|왪�צ�7(^~�a�Z{#5��&�Y���Ű]��WJ�N�5�������+��Iv^�L�N�Є.b�z���s}��n�,�P�|���7BD9-;��<ˡQ�����
�껫���[N#tr��jښ$zM
*�!LL�4�LUF�ɋ#�����a��aL)�ݽ�����}�'�8�8�8f�y������L\tv�:����+�jZ+I8����/{κ��	x|:ˇ��%v�yr[w�����{y�b
�
`A�R�v�2��ndZp����?��"
�ٙ���.�lE������R
:3k�nG�K܊��!��p���*�Wb/i�Q�+7|�嬮�9Մ@��
z_�����)X��!P���k�f��o���T�'�:0�����h^7�%DY���9�sp�ӻ0�6^���]�ϲ״O)�̹�Bϧn3�M�	9q"oS�b3މ=��xF�䲽�����7,�=;K_���:>������{�جI�v�I��KCٌ=N;���܇5�m=���Q��W���\�vة�[%xA��5�.��}�߳̓��w��D��u-��w�q�Q=�9)�?[�J��b��mR�E�UZ�n�X��v)1;��u�q$j\\�5N��]C|�I��/�ӆV�&�[wtZ�F�����Ӑ`�� �wk���^op|����NW`a��6���J�q�j��6�)�,��΍�ړ��l��;v�"q_�7�ٻ�T�u��!�޺�'���F���vuar{lӷOp%[���yM����N�x�&�r�CMz�������GQ(;D��FH;K,m�F��F�&��k����21�u����"��S�.�M��7q�^Ŵ:�.а*�.\����"���7T�_�O�.�Kn�����U����#m>ծ.6��SjƬ-Y.6Ub�emP�n��[ɛ�n���囯z�2��1�,���7Y�Y��"�{�w��]�">���W����I�']�������Џ���*&!���m��҃��~6M(��z�ԇ��O)�*d����N=���z�I��]w	�(��ϼ ���it�d��3��%�_}}l�QQ�Se7��<�k���A���(5���Km�5$[?a8�&yr͋u/۪}V^G�)���UT_�ڦܙ�&;�e��KZ`��^�z�"ゕܷ���n�g���wϚ��k�w䲙��z_�;��������\;�zx:�#��;f����I��3/��oՓ��IKܵEj۠���.��Ϛ�����#��u�J���w}�Y����{#�GzQ���G�ft�<���ZT�X*��Y4ő.��:f:.y��kc��gXT�m��C�z�L��!O{7�3�55�ؼ7����U{6*r�lWgk���z#A5
r[9��UU\���R~M-_o}�ÀZbb"w���74�OJV(V�x�����]�S ��.@�)��Q���`AX6�Х3n-����hl�I�'c@t(
i�ɚ�"�X���*V;Ţ�9�"�;��u��r^��&}4�0=�>��}،��-g9�Q|0���{�/wQz������\{� G"	��@I	�Vi�|����m�fHbb�F}5��U�hQ�W��C�؝��Y��9��{6\o�	�1S�++껸������1U@�b�;�C&\9�=��L�T���U���<���#�s�x]�h�U���Ó�=#n�C)3U�9�8B���)T����{�ޯ22bE/:?h�G �$BL�т�.��(;\���@x�`)�˅Yw���3�j�A�E1��>s�װ�PD_]�{�x���o�s���O;�~�����J	�)0�D����·�^]��[���5����q�EE��hB�l����537����&f�{��#֐�b������[��V<�}vR��Qq[42�K�J]��,�l8Z�	�.Ga�o�����������kF|E������sc*���S�q����I�Y�z=�ݙkX�jT��3�����*;���E整���7�l$S�$��x���O�7~�M���,���v��Ծ��B|��e&���Wk�59�ժ����ee�^ʚw�y����嵛	�y��El��An���.l%��-P3�/�>�FWX�Wb���#�>�u��|b��dJ�nP��SBJM��{��U>�l�Gyd]�&v�.�+`�������+T�}|�޳��Ϗ�,o�[�M�ˏ�����g���_rrDo�^w�/�&咉�S��;ǖj�	=T���ƤM�4�QyA�lMV��w�w���x�%�b\CSԤ��{�$Z�ӷ=�s��]�$sx*
����|���{R�W`�jQX�iyļЗ��(�Y+#��iÞD���6�u���f��K4�)�]4�U.�z���rm��,��w����>�L��>t6�kWwT.�)KM]x�E�8�1N}���i�z!�࢚�1ّ{7���0�ks�J��t>�+O�[ú|'m�Wa�]�U�Y&�y�B���FO&`��X���s�q�np�:�%���s"���Q�^mĮ�dϳ��~]�>��+<7g���̩5o�÷��L�k%7�i�{,vҸΈ��	�lDCyL��&c-zs ��:�?Vo`�T7���6O[�f(�v����ڬ�;�	_Ә�[�=���d,�H�ծ
z����R�;ǔ
�K�N��fQf�6�;�J�f�!u��=�;%5f�;�{�_ޓdϺ�ME��p
S�
]�ΊQ[4�:]e靯[��k�]*Ez���,���� �,=���(��W��*z��(,�2��+8��|�,���Dr�e)DRÁM@d$�oG9VOf���-�"z���FF������3�Ip���7-�#yuQ�����Yers����4��S.:�=>��mEDW7v�S�����=R/�ȨL(L��Æ��s���o��Co��Y2��g����y��-P�4��O3�t�}�yӚ�B�&��.U�7����с�)s�/c�a�H��j�Z���g���^�_D�T��4���Q����_2#7�lt=�a�W����[�ec��CF�k�S�$R8˂�$�P���܊�@jk�o��*��:�T��/�8��w�+4�`c�Dϐ�D�C錎�����f`��^EG��}�'�3��\|��J��~�
T�,2Ի�����KY�����Kp�������^ә��ws�ۚ8Y�q��e�g�� �aG<~:_j�Tw<�$��G��<mkgiy@Գ����a���kt _@��Z{�DD�tx^'�j��Nѽ��)ʡ�ٝ�*��x/O�w԰�qO.Ŝ�C�Z��ym�;�m�mD�{�.�݌�fV�r���㺮��.�Ӎ�|��,l�.�R��>�q�ዷ;�gvË���q�иn�.z�� :�lPm/=ӣ;���/]�~��=�x��ո�r&�gu�]v������ニ�=�l�v��|��غ�m���,m��	֣l�[dm��{u�n�n��=�Z��(��9��EϚ�y��6���:��b$����b���E=
��ښ��n�������N^���5ٴK��iJQ���5>Ô�ћ�^�;���������C��ln~9�|0�@�#�70��.|��h���W������}���"��,r�%=7���K��}�m�7��1]3��t��
s4��%Q�3�jV�I����Xz���_����y��wMs���W7� �WZ�LO�~k��xkx_������L�z�c��jÇ��k묝n���r�'�5���>��^�3��Ϯ"9y���M�p|�˫;Mtߩ��$Z���E�p7U�&����|�`}��*g@,|��gﺂ�{G�8�dݬ�\���;��A��m��oQq������?�!��ڀ*�1��ٵ��_��Oݮ���Jư�eFXΑ~�V�93�v�Uz'7�}�7�������1�#fb�X��RQ!(����;s�k�y'��ڤ�ۗ���vëfǓ�xe�"X�?KHG)�y�?�j᯾��8���=�8���3�h�QfLOx�^��T���5&�{722"�)C׾�{�ەH]�y�xJ�-8H$JlUף
�y�mF8�j�{�P���F�{^�K~5�l4B�U,�w�͙��{��K��U��(5��N�V���K� �E��	�n�U��%�e�5ۥtK����*v�Wd�:H��v%�y0�#6n���y����q�%������f�[�=���#W��p� �)51�j8%�b`A�-������B�S��[g�ϴ�3t��Oށ4��Ә{Z��y�m���ɟ����l���CɘfǦ7z�zw���!s���7>�f�~�X�ۢ�w�.;y*-���\1��!k�۞s�n��6}I����s�v�Y\����S�\��s5��R�.�4|�·���@��lP�ãL��B6Q̼��TF�*9I3�m�����'dt?K�v�>^�W�A�mC.���+�y4=�#>GΑ���l�l�۶�qv�]���!�#�e���,�׾z�Zk���<��|�__p�2�j�]�Ri����r�_=q^Y+Ҙ���"WRO{��wk���]�mO��J�[�.��EU�(�שˢ��rW���כI�y��P���#�ħ��N���Sۯ8Ghk�M���̻�D����L$Z����4j#���ن����On�Bk���;S鏘�*8�[]�������P�*�-��!���¼�Zv�#��X�֩3���8���8�mL����,�״��x�1[��u��uΥL捁���F��1�-�4썉��+��M�l[um"�޺}�u�p<�i�]
u�E�:�֫nԕ�e=��峴�����u5P��ҫE��5���Ŏ��3���������}3�����Q"�Q'�#7�xi�Ln˻R쮫��z��ܙm2\݂�رi�T�ڇ��/��t_Gځ�r��D��IA�wv����2�)j�`Bt�ԡt+����&N�	�kF�f���8���/UA���#�k�ɏz�B�E��qY3{����u��9���u�ŪE�(�Z��biq��S2Q�Lշ�7Z�ڹ���k�R�
Pa[�vh^Igӄ��hO�Qn�ۗVMԭ^9�~oqX�yu<TclZ4P��e�g�[��]}�G��
ڲ��s�]9�$�s�^o~P��x~��v�2a2�����[X��=7y�h�Ϯ�ř|��Y�ۡ�aӪ�n�\�O������ǵrU���u�	����K��*	��4ӭ���c3dZ6�p��������yu��.�W�x�(s@�ͼ����T=}�
,����c�O�˼5_u7���ܗҷ���C��`�4m]'Q�v&���o��9�l�T/�oVT��i�L��-y�փž����3'D���n���4�w-���;g&�I;�Io��o�p�FrĻ{9�!���ʒa������ڏ?ǟO��b��<��md�w�7ԹO����d�D2Bq�}�5���elh�s�C�1�� 7��Z�����O���K�2�-E�)���H�9J���ڛF�7�0��Jq1g+HT���u��o3m�����n��>��	�E��v������f��r�����V�濨��3��wSV#{3�pjJ�`�#���N�j�t<p�<a�mrSm�#(��gZ��;�NKh�p����rf}�Űz��o�SL�m+�蒜M��#b� ��V+�:=dv��k{ַ+�M���.?#��7�`�ߴi��:� -�R��]��G#���O����3��i���}��&j����YW*[Ϧj��轸k��s�ƽ��T7W>�i���+�-=]CϮ����/	t����\k�M�&�-��&�</�O]�鹜��Aw��TY��N�.]?;�$ܺƞ��A��b�	��6.�a?d�����U���f}]�~5r���^��[����ڭ��1.������i��p�b0����ɚ�H�j��s/95��r��Y3H�|��vJD�gx�U�sν�[� 묽2^>����}���"LsX��r1Z!��9��s��o�����%Z���}Z"b�$�w�g�{{����V%g2�oκ�J�{<�}K��_���d�]�O��+�{�gʉ+��[�K�m�p6�t����c����{K&e��p(p��7�}9i��5��v/J䷭�)��^�����Ù�w�ܸ�S��<9.��-�C����
�B3�L��U���E:I]ruw�2�H�~�5�r�ߒcǣ��ī05c��� Z0|j�H�~��hݛ����뿭m�&&�q����p�aCP�ܝ��t]{F�]����3c�����Yl���������ve\� �G|o�p~�1�X��WR�O�?�H�R��1U�-��z�5�À��^�Wu-=骹�1��7��d?' �}�}up���w�Wx-�y�C�����h��\��\��N7�eD"��^߆�&s�Tl3�YV�y̼O�\T�K]R>k*vR�h�s�DR��+�S
���Oƪd�R{G���1�����{�-�1A"ֿd���c4S��s{3�ċ1V4V�m����8�80�~o7Ms��\��c,��w%$-�B:�E�9\
��uÆ�)�A�r��y8]����P�M4�=�v���瞓�r3���t��bu�\5Q謩1˴̀��'qs�;��~Q��c��mxq������Rr���7�>��d����+��/�s��[-z^t��tgsa�6�
�h�^�������ܦ�YVa�����]�o�> ׷:��ok���g�u�����F�k�u���Ӭr��M��ֽ�6�1�E�.�[�x0pS�Lp\K�M���}�\I�~���W�»1w{n�k]6CS�וiu���@,��O].���g-��U��m�=�W��Ǘ��� ��;���N5)��g�����hu�߫�=�GZ�*�U�7�!�cX*���u�=0�OP��?k��U���˭Y����&����	�)�^:�dš'��Fّ�"�>BwjR���Du�]ϟD���s��͉�Z���>̷;^+��7u�=��#|�	��M&�FN�mN��z;P�zP�eem\���}Q5�cP��93[b����k�9��U��T�!���f�Q��튑�,*��3�{�Q�)*�x�{��Օ��;���[�o:[(%�^f�y�y4���y��:j��{�j������^��uk� �nP^xû��A�h�'��8���z{<u���T#@�S���T�9b
����Ԥ(�v��Kh)~����e�h}�A�,u7AN���ߧ0i��-ڼx_�2fw63����_��/x�M�����4�=��ʰo����#�u/G��������6E�&��Vk�u�d9�E�������N���-�ڭur�M=��ᗓ�<�9/k����&����xV1��v.[��i�q��ڃ~�(���]�?/���T��6yU믮�9����Cm���?u�EC��H���b#�A��@D�)ŝ'@�83y^f<��j L����OF߹���Jb3R�[�3���*15�)O�ڭ�TL��r�ahP�p�M�Sm;y��<��ߴ��
���I:��Y]�K���nڻ��+��*]jn�.g}�\�E�z8Y�9�ƅ�Ω��")�����V�{���3�g3w>&���ֹ�H@�����8��d�e|m_�����:A��7w���=��*Dn�H&��Zsj��lR���ch����ݘqɛ�ˍ��'��]���^�/&ss�d�&e��B4Y�=a���2ey뷩(�e��:��6�U6Rѭ�n��a���o���Dݰ=u52�8N�nao��n�H'x㽝�{>��Cm@���kr%�u݉`RTK��>r�[��u�Ԏ��&�<ؤ�0H=�|O����y���|b��%Le�hA�փ~�����2���o�\������?��;��w.xz5���^���T�O8g5�L'c{M�u+�u���ɔ��}�T���{���yY���1�:5�|��ZV��7FN�{��#Gu�m���r<�Ci�E�
7p
��ɀ��z{/�<~l�{�w���,?k���n���	/��VT{��E�i�v�w�P��'��(��pg��N���ܪ�
Er�o��o(�cfQɮI�w]7� ��@����X��A�Pbc5�X�ǐ�bӞ�;sZL�>Q�v�,8���җ�Y�C�t���pl�݄�ٻ�\uBc�#���l��V�KH�JL� �Z��:�J|�v��O=��9ɩ��m��8Wc���̼[V���a:���"���9y�)35׎����K'߰N4@�~+��-��s"X�ܓI��o������?RW�GU�퓼��g׆�<�{o��I�i��E��W��|�rJ8��s7+�7�L�V*���"�.��4�1w��;P�oo�7\H��+�����f^�d"b���V���V��N�9�����ɝ���jc�f�,#W���e�:��QM�)��ca�<vҎ��������ܙ��� ��hB��A&�q~˿JU4 t)���_<���g$����{���+���7s�0ArՐ�U�`�5c!+HWH�݇vd��n]�+��Y�}�&,��IU�w���Œʈe"��i��/2�D�o�ݪ�xg��c>�שtb��r����7ݯʣ ;�>�IW��~���ʰ����O��"$�D@,3����ކ���������M��C�&�Tq[a�P��AY*?���q揌���u�"B�b�o��Q���6u뫘�}��Lؼ��z��M���t�]v�.C׫�s$�Ь@����Ah�DM���s�qV�'E߫:�׼<!��������gނr����I��\UK��z#x�����-@�xT`�	�@h���.�y��I�%�tz�LOp�K{;ڦ��n=�쿾����~��<�1��o�~�OM�*�����'ť
>MB6��:_�=�}�G"2��w@|��y���
��ԫ&�L�W����X�nz���+�.����l�Yf *�ʔ_fs�-v�X�6,c�P���R�%�t{��=��-8���= �]vͷa�ɪ�D�R�ux�vQqE�U��~��#�+pY�/�C@٫���8��4�
w�E)y����km5�S�ˍT
����"��e�nM�Ql��QS���.i/�9��-�7d���Z7�N87"�7���+):�&� э��5�V����Tu~�s�w�]؜򦗑�@�D�+�)F�s\)-���9����Vŝ�dB<�`=MI�мw#�q�����A�p�ғݪ���.\6����>]��?ú�	�~�[��y��'ɶ�	�UpƠs�n�n�yG��F���N�	�g��H���/Yp�1e�]�u�gx�7\�;ns�� �)�&L˸r'\��2��$i��%�?�cg�2�e��/`3��N�^�y�qk����ӯ2�/��@����6++�bx�]N��&W�\}�6JE�{��(
�٤�zq��S��{rK!9*��n�f�.}Y�]z�w�����nDߒ5x
�^yC␋��$��g�u��Ǿ���.<��֨P�j�Q��Y˸�������
�F{_��Q���ĩ�j��<��A�ks}�9f^�/���yǮt�&�|��ǵ8*�����)��̒*f��'$��+/�F/b�#&:�ԧL���G��ߩ��T��Y�0b�='����uo�lN�\lgJ��AE�qq@ᱶf���{�ه����	>_c:2�9X=�S��:[���>�N�����\�9�]VY�BD��o���Ƿ�Uvyy�0˰�=<��gMuڞt��N��7n��|}���i������>��ת��JtB��'�9�k;D����ulW8
�Tf\.x�z���<�[��ܞ"��?sr�cr�Q��M!����{��Y��'��������F���=G͹�:�gɾ�\2,mj�,\�svVDu�c�3@��l뒤�Ϧn*��F��ޚ����ӊ���R�W{�J���T����{���Ct��NK{ʏ���}R�x���&�O��o߫TmQȫ
�fȏ���k��;�F!8'����}�i��٣S�b�\d�-�P�۾�{[�����ʂs�k���B�+�E�Q�gw�w�<��e��=��{]�P�|n�,5΅�c��奋�ٔ;�z��}u�6�,�7s}��^�;�T���s�$��X4����|��X.�~z~hB��w�g?>3�ɉo�x۫Įk���"K"=��a���/�
��VB��z�c6�1�9Y��ѷ���wW|��A�+r�-�%��*�p����Nz����3�eȹ�-��t[k:�.	߀� ��J��>��Рxن�o���f���dN���?;������|��/O�px�0Ă��Lz�]C��b�2�n��de7��&�o���zW�9�&?M=�Q3�����]	>��ڟ�~يN��sW���o~yI�xe��:�۷D!FF(PZ�\1���]c��z<V'�����'f�b/�-sѕ�S�I��C쵒�f�[0
��h��!s�,�F�5�.����Aۈ�MJ� ��1n�N��hZ�r|;z�+��w��x��̫�{3""���\U�6q�ХV����E���B����<j`>��#��&�/u����d���<�|�e�ؚ�u}cMS�s�n},GF���ZH���~d猬S��Ehu�L a0!�F��^���{����6_@��������݇s�tk=Nj�s��jh�}'�BoH�P�a'I���'MoSa��<�V�;ml8���쵣�{���ƻn�aͲ�����0��F�L��pا�ޚ�n���2���Sw�0s0�Sa�s<�Ԋ��p�rw�]iљrG�ߣZ��T�-g�]f�w��߹z�#��s��M��߰�ՕAmޘ�諹��N`�[�ufr����վ�>��X��>|�{�#^v�zmf�q��@��JA8%�$�����vr}�K��ra	����qNttת�>�c�/3�Y�t��|6.�"�z_?osms5>�至^������5J���o5>;wȱoo�?DP�nc�?�����j.�ʃ��^� �}�.��� �}}_5�&:E��v��Ty�G���N���3k7U�{H�XM���ɮ�X(��4F1*|�[��mmv�����ù�o���Y�|��\�e��j��(�6���7D�EIm�9�o[̭���y�֙��JɀUJ�z�ޥ�{���(�%�e��&(�:����(��K�U}����T��M��D�L*�˧Ruv���<��fuu#�=��c<9����`� 
,�򞣆��|�!��b>��Lr�SNon�'G�L�������y�Wb=��3���V]�J���!D�����kݕ��W�Չ4.%-��;��m�p�7y����:팫�Uہ@�w�؏n�l*�����z�]&Ԕ:z3H���F!& ��HVＴ�E���������9O��I�++ܲ�n���8@���7X�w�bH�Xp�����hV��C�-9��+��y����j���=kG]��p����26��)M"g�͛���P�ǩI�Ė�e}
7��������65E��\Ad�@�I�a���!��S�y���U����	Ȝ�M���[>ޱV�-�:�ݗ&�W������*��岘=�����^��DI�C��.v��,J ����:���׌ԇk��N��u��s.�=\��۲��]岮.e+��p�#.��L��������ߋ��T��i�L[R���8�vFw
-����.�(2��9ڸE�:�m`r��hJ�KkbGO�I���6���)b��Rh����Q�K�����b����#�����Mq�[�Ʈ�1aB���d�UjK���l���-�;�z�2N_n�5Ŷ^���Ón��>SiJ����e���8��ԓ4�����f���E��T��'��娢@P/WV�%��w�����[���������k��!;� w��6�7q/#�[/�N�GW�M� /y)����s[�&I[�U�7��xd<��j�ovv��_����,H��ܬyC�ɼ��X�̽׻�!��!���7Ef��ͫBf���*���_"�8xe�p�&�)a�Wi�c8�^��`e�!L6g54i������T�C(��PH�=k;�54��뷽08��/q*�Lm9��a[zd�M4I[�K�ybM3tg�u�(�V(-��I��Z&�)�� �]G�\����?�c
L6��ufVk��ylh�۴����V1�z�eDl�l��z��n�V8n����A���䝥͝����.^�Nҁͨ]EG���Cm��$O�
��{x�s6���x�^0B�gL���;{��q�M�7�o3e�Z�Bv���:��'V�.�w�>sp�O|�?F�BW!Hd	b����m��h[`�������v�m�$]wA���(�����-�j��4�V��GOnN΍��^fڤ����:��9��k=&X�8����M2�8z�۷��󳏧��ƶ���+ǖgm�'Z=]�9��sq��vF���ܯo[�uжm��Σe�W�����q��v��9{�[����l��Z�9'k�º�nz�x6с���q�]X$P�49+N���[��:�:��h�j��]��M:2�!N-۟�p�N2�lv�Υ麆�η>g��=<���ˌ�<�=��F���r��yړ�0X�v{����mDvj.�;lD�nJ���tv{u�=��m�/em�:��
26�-�U�wu]eV�ܘ@��1�<�zt�s·q�s5Ѓ�/Xn⶝���;pc�v�:B��.;g[pp�@�x�̼����۷�S�M�4;�I���-9��ڧ�ndM�}n%~[��2����m�=��ϐSqѤ9^3�qM</���^;^�O]ߘ�w�g�=g�����v�4�;Kr��z��z�N����3;��9�;�N;�cp�ŭ�w���������8�zx��U����Ih��n����~�L������w�\��������+�<�z�D��c�hN����W'݇s��<��9�7A���G�� ����X�}��l�>��6[[��s�`�׈�.��NOU��6��<�;鱿KgFC�)�Gv)�V� �9q���7������C��������.�)������n��8�b����=���{���k���q����(��[tlwvަ�1�{��+���N����y��;������u+� �:{p����k���q�e�r���;���g�}��]e-�w��한s�g�tgV|�qѸwg������8�vn�i�Μ�'s�y�ΆQ��i<��ζGt+��X{�D1��mۆ�oF�f}�B��s�qq<��r�	�@]<���nŎ^ڃ���s��ps���s�=�q�z6W����%��\`�I�[����v����(y�[�=i#OY�h�ٽ3�n��f��q}��w]�9۶d��A��nd^��v{Epmn�c����k�Ĭᮎ٢0���vm��{e��p��]mv6��5�-o!�=�C���W�Z�V�;����l��QW[��A�E{��µciѬ���z�]NAK&�-A-�s�tMV�[�mn���@qvk#�$Q�P��S�R{ڸ�� ����
��ż��M�#��7<�۳n��x0e;�l�Ӏ��2NH���ടgN�|�M����u���&:�zh��1�Λ�W91B��и�a�h"�$и��Qh�7�,���mП�czMҹ��_��|ܼ�:���^o�B�ܗ��W�`Aw�m�Ԗ�������6��^��s_>+��~`G$��u��f��v��jI53���Ǽ=�:�Iy�lt�����>�NJ�ˢ���ȌǗ� �`���=^�D80���� �ؾ��w�j�<��9�:��XK�s�#�a0ET��M�i�ɀ��Z꫚���{�vPA�}2�ADzD�R[�S�򛥹k:����f��*���K�b�鞾y���;�z�������Z�Җ�<wͽQ�5ػ�ѓa|m�C ��G�o��A��km��� �p�K��,�y���q4j9��{��ۇ�������9�_�@ƙ�u�5傁O�'��m��������(�U98i�^����rN\�'�{ʽw�=��_X�o�Q@�����+�cxP��*���.�d�^��4T�XGe���Sr�S�F>��Ⱦ貉=3;����|��w1�OT˳ݐVm���1����1�/ٹ�#"�'vsF��b�����K�t:�Ӝss�F{Ԓ��'�L�0�9z��jƛ��癑��_V*��,)��<\d���y��{�sf�]*������x�ٿ��2�
,5rܾ��T��	:�'��s�x�1��;�߼���*-����t1r�r�X+��Dݲ}��'.P`g��o�^���@55�#��av�p���{Ƨi�V�Q����zͺ��4(���;3�'���_|�i�BEQU'����'uԡ;��3`쮻\J�@QڛfM�����s�خ�onh1ú�s������X�������%Kש�Ms���О�4.k���w��ն�E���"��F���70����&n���_��6�f�РU�Cm��܋����ϫ�K#-[+ʻ��^�1p����h��i��]�g����on��&�˽�Ò��3��A<+����N]�#�938�U}I{�}ֺw���V�/�S|��2��'�nDB�����Y�+��ʱ��2���̕i*��v�e��Vی�D��bв0���L��'-C�/�d˜��\'p�Q�O��P�5F71��	�Z����Ÿ�4�o�o祡���c
>-̷�˿x���A {v�Lqf2�lF%�@`���}���p+���d�f>�;N���/7��d��&�D6�e'�ԭ,�[���K�R#��v4Խ�N��S��t ����X�qx=~t��99ＴM:yC	�e�6��ӏV���oד\�V�0�-�fF{v:�yS��rr��x��zݸ�}�fn���]������/����ܠ]��x~_��z\CޞSy�Gݑ��o����틊�aѠT-J�ݦ�0`�h%9~�*�Z��{��L�5�u֧��O�w��c
i#�!��(�Pe��l��#=�ES������PI)��[����ů���_���o�ӡ�%�:��ǰ��ڷ�bS���	��}*�^q�:��讴���j <�\_(��p�n�s<�����ސ��v*0 �����s��r�g�ѐ�<��{�͎�
0�p����&aO|O�2g2��Y-iJ1Wt�Y�mXl 9����й'V�3�U��Uvsv��|x	o;F�;d����r���?/��)c�����ۇ�ѸIA�9j޲O��u>O�zT�2��^T��8c���0|��o˅�������s]�}�*s�k�k��{y�79�N��L��!��Ƹ�7<��Vz6đ�7/�V����m�=�<g/]��$����!.^�nR^������7Aӛ���B��^@�8ʾ��sN����q.��nUP�B�og��b�u�W��IL]�
=��	��ۆm���*�[0���{�;��|cy��I6�lh�kr��yU'^;��.\׼��c��Q�/8�0��཰޾�/�K�3I�"
)D2B�����_*p7�V�Na͜*��^D�u�=苒ʈ�(�q�y.T0}y=.��?V��o�ٕi��o鹫��T��V����{���p���,����w�K��H�w��ݶ.�U�ï/FJ%��a�gEZѽ�<}N����|��I�� (�a���Ʋ��H��bk�v���]cv�\����՞�\oU1W[�Kg�����W�7����Cʃ!3�Vl����TW�fo6xbGY�'�Rte��3yv��ץ��x=�z�;�*�u�tk�u���5Ӹ����Kr��MZ�,�!n%볶��[gʧ�7mն�&jg͵�A9;s��������=q������ͻ;�kbrՍ�6��(���kaB2�h�d\x����m�;�5��e�׮�r1Wթ��Ё�$1�)[e8�1��|�Icd��j���}�|8�0����3vz��#]�=n��i-W��8W�N޶q�P ���y�H�v ���t�����9B��r��7�j�o���X��� ]�'!N��.��`�v+g�m���^��{�z�=���p=��U��e�M�=lDL�=���;ްg0��qق��˾��ֹ�]�XP`0�Ln��eW���xP����ǎȯ]��i���}���u����x��F� T�;R+�z9�훱�/αխ���f�db����\���>��G��6�WK�/�bw�r�r�z-�o��~�d��q��5��?g�U���#'御B+�rC��0����jy��ݙ�=��)�`28�<:}+}]��"�O7^��^Z���Cof��iw�sɿ���߮�8�P�(L�m��>�E�g5�O���^��Vr�s�S;O�9w�����L{}�7��gǅ����!�|�]͈�"���@����$,z�o�_͸r�n������;��g.=�8��殞}9M��ۚ��"��B
!
7,�>�v�93KB7����Zk��;.���}��v64�2�Q�t"P����\�!�9y��^�NHN3�T�P�"��PRl;g=;6E�b�]>sWc��o��LlP�KYET�+����ܚ&j�w!�=8WM�W����J�̛`�n�}vֽz���Q��1�S���N����.��l2/}����3o� ���o��7ν��1�:�+���1������9���U�~�lP$ٙ�����<ѩLƻ]I9͎�9�w�͸��W�u�/iٝ�*�ث���b��S꣺���LT��ɢ��2�E$���6��Eђ��a��׏����\�''���	G�/�P��~�c�r+f���K��0燽���?�MI����{���*֋"�2���)�)ϼ,�l'�w�G]�f��}՞9�˞��#��o��B�-̳UA�J�c35&v���Y�-^�����C�ADK@�jEkU�4\�A��݄���G��gNA̓cP��B��Kd���y|׽ˏmkس�2�����/�ˬ��}����}sǳ�gS��
C��wud���v<f�K�h��-�����^^R�����*���o&n�v�f�I>�oq���Oް�Ө%��q]�x0D�>��Og�x[ƍL%�h�̉��T�y�@I�i��ue�)���V�8]=���[l�I�=��E����;�{��������}712��ra"�rhWv��թ�feܜ��l[�8��S��$�
���%e(/n٫���SW�{&�6,)vf������卥�M�nh7�؅}�,�q'�ݽv��慃+�a"�BL%7���8�`���yy�.�6��-���^��d^c��g}=�ܞ��X!����Wk#6��E}A/p���t�4ު��? ��^]�����_C��8MBlg%
w���mw���a7�Y>}���nX���?��g��{�.i�3�#�>���o������l]R}9��(gv�-v�����D�1Ƭ�3%�8�t�	J��n��2�nӫ����� ��՞õg %E�Ԟ���h7K�m�����1���YBuS�&$���hk����w>-<�S�} �x��%C*B�DFF��uY~]�7)?�~C�x���5��v�$���¨�y�JN)L(?mҮ�1ĪA��xD�Wt,��0ǽ�u"$�@�""�p�t��m����J/�NSH_�%���9�Wgf��{<����,����R�����<-��eo��� �- ���i���/�:�v:������|�i��^�hP�Щ�􊁲�}�p�>�3�vE���A*NH�;y3�n�g�&�c^��Y��/��}b ��/��\�����eV���W�b,��BM�#�o�>��W�޵�8LÃ��I���)v3"��H��M�3�ɬ��O�2�t��j�{>��%�y�1�uw=yb`0�KN�Õ6,	cO���輪��5�/���&�U�
�n�M�3��rnܯ��*�f��3N���Gb����ױP�3�/3���I�
#]�]#��d����[�z�t{@�"!�*1���A<���	ͻ�ۜ�5ZVd�RKj, �P��?[�&.:�lp���V\�CI������R7�X�įv���È�2e�{���!A��lz+KQ��o��5Wm��� �(���"a϶xux���}U��Ɇj���GP��u����LbK>�w�|wǧ�br�����ف�޾�Y�Se�ZY32�I�U�����~��ڲ�FY�P��wuԞ�
��Z@��t�{��)x�g�|���?]�=�u[���Qq"�CP\4ͽ��Gt�I�U{|��)�T_�αv-��;�d֊�m�z�Mǟ��?w��{x��d�����v��΁��nn���cNY���n�����W��4�v���ס�he�)j�ݓk
�5��7x����6Z�ѫ���Y=n�7apq��Z8R�v�<�h���e��.�s̛�ٻn85m��Gu�v ;I��u���w]$�,���n��ۀx�kp�L�f*�����mb��`:'�"���宜��kmϝ��x1�{�}|�듞�l������hrkp��m�]��on��:�����o��+��G=�=�Z2�ˎE���d����׳�K���
r��Ы��yz*C1���s7���v�tL�Z�ۡ�����{����h�[��|0����Ѽ������'�sqQgOnW>u�sW�0��]�7.�%�Z&Y*?�o�,��^��x�}5�[3���_�T�E/r*�6�Gy��s����}~�ٓ�7gI��|{���O��!��	�̖�C��^�ᑊ�V�����v,cŽ��褸6�e�y����� ��~�Hz���#����	(h��/f>���m.��)%����>��\;��u�4�4�D+w�x�1�=;����b&��=sNw{���]W�Q{ٚ4��(l�3@����<c�hߝ�9w�}�����XЋb�Ą>�~�f#���+��ӹ����ɉ�B�_�7�cr^���E#��u�M���nٸ#U��s=���tk��9�ӻ��
�n�"�u�������Х����^���Yj�J��E��O�G�9��;_�����u�8R��Y�3��R�U)g0�kNj��|��K���v; )Qh�9Q}:�p�x����P��sC0ǝS �hwwnμ�x����
�}�u�S�jj1��K��s�H��}�~�z��;�z��\�.���Y���0�;�/K��{0x�����O���l
 P ^�m�=��j�;޿z�"��:D�(�[�5^].� ���1�Ob������5�{"�רX�`�$e;�i^Գ�N�_�0�z���}��pMIv�����_N{O�<�l��\� �ұ,^ڨ��� �)�w����ڵ;��S�K>N
�Z���ῌ�t�g}����ؾ��QRo��bV�a�N`s��l�_a��� ������dB�ifu�Î���\��e�,�k�y�ŇGM=F���:bD1�荳��v��3~2�۪b+L!���}k��ivW�g� ���TN�>C�t^�@s
&�"S@��{�)G�e�vϟ���B�AȦZ-(e�ʘ.��Ӻ��}�=���=.&�yw=��۲#���J�ޏ��d�G��U���\�p{9Z���~ۋ�AD(pKni�VeK�v`���UW�M̿c��}ٻ��V��S�z`�)��G��h��e�����y�8Z�����|��U���/��g�5���+��We[�h���5ܿ�2�jj�;�!r�i�П���ǰ�@VE-6F�J�m�=V��v�j� 2h��"�GnZ�S���z��4�]� ���s�b˹u�&�y�]��7������^@3��ޅn����z��ۡ�Å���[k�m4�U��v]c����w%�;��?l� ⒊@vޙ���Ƈ���tɛN�y��/�w *�T�����,@�V�
=n-�i^M��p����Y2���82�s�Icw�������j>��/��M�o�y�q�"y�c���9�gt����&� ���ц�����V�ݣ0���V��9tXo�E3��7��0�����ΩDW+�v󑆹�d\���z��ݥm2-�]p��,��Q�������䏉i�Vn�ޥ�󀓊�i��Eŭ��ƹU�6��o� ��g�W���Z�>ƯC;�;B�U�8Y�p]�w��ݧ���ٰ�w8�,Y�t�����զa҂��e\�V��j�U�Wf�����*ɇp�CY-�R��=[��l�D����y�᮹Ӭ|���=(�8	@�R�e��G����^�_F�<\�6�������٘$�bRP��\����K��[���m�F�97p����ӮUY�x(�f�Y08�>;?2��Zw�v; ��s�� �W�/5�տ�� ]��2�Bzt���I;�IW[���=2!$��E�f:�z0N�u�q�y}������d���"k�^���(|��[�+4X݂�3^��6w�z{4Gz��Y��B�IvCFv4m@��꽸5}�j��e����W�ߣ�O�����HW��x����`U��$��NM=4�����Q�޹u��t�z(��7^�kf��LGʕ���w�b����U+��_JҾ�K����?����(:�@�Z�W,p~77ƖZ��+�ܖ���95����m���h�z =�~�j��\��)����~P����o�2�^��bϨ��O�5�ۋ�"/�Y�r�Ei��޲I��-(�ʈO�,t%�U]����u�xU�V�^�Q�^�=����%Ϲ=��3�|�[wO������G��^S�w��=m�[�<���$#$���ص�cYu☘���j����To�s�}����o=��'���|}O�D���C�6uH~������DD[R�"�a�h�fK�#�<�e�-!70��ν�O�w���ߦl�w����ۼϼ9}�
�B�-�Hݴ�#�������[��i�<Fi�����f�%��L���퓣��!St�f�|^X2�a�{uK������F�9����q̞+�2:B�����&(�e+�ӻ�!��{�3�u���UY��Px}�~���R����Se�t���LflÀ㌑8J��&���.#ro,�s��sع�n���;Ls��ܚ��v��q�-�A
;
{S��wT�	��͈7�X)F9�n�Ci�⽉����z��e���
�y���\�+�!�=�G$���7f��g)�o����U��}\oOw��=�4k:t��Y������z�.*�G`��;�D�rf����+䰂*�v�-��������,���2���:s����z��خ������q�Y���^Ǳz>��:�I�]f/MzP,*	\��ޮ��.=���][����MV�]��i�7�� �g'6����tz�Utw�S���}�j��a/�p'���ny��^zq@���^l��ކy���8��&u���V&�_T�����U�R��\>�n�q}IQn&f�<�/�Of�N�ζ�71���V���o�������:�n����$e��CU�w׎�u:wm�dƖ������C-�����������<S+���9�hݰ;�}�]�r���;k]G>q�1o<����t�A���vK'�s���qm���Y6:1]�{[��6����6��-۠n�O�Tpx_�!����mֻo�ӷ���.��99[�jC�ȧ.���`���W1���r�M�p�}!Ll	�2�����W�&�g:���3r�O ��eګ�e���5qϛ�խ�{v)\�ۮs0x�&�6����0v��l�(��^�������:Ы�]��s�m9������?/ �=e��V����s����
w�K�7b�$�bS~Ċ��H���}��{�p��m��h������>�8����l�P�O�L���d;2��|���Z���ahCP�6�6=0��(�i/�I*.�"�lH�}w7�A��-z�/!����9�Ϟ���g{o�J�?l.���!�_Dʀ˄߮�;t"��<�����jؕ]S�M;\�z���W�����o}#fa߉3��MgyK���4c���􆠹e$ϕ�zf�W���ژ"�D�,���>[J�ﲶǨ��'<LT���n�V��;k�������ݷhzMd���o	)������[E��i��{:�+nI��pBJ󕪨�N�Q��$��3��_����	ٙ��M��of+^��mAP�kB~����(��ί1>�r���TQ�ܷ\�Dw�-���jb��ǥ��~�������%�ί��˘��6��Qc{3y�N[W���k�n��+��W=<�r�"����쮛�Χ2�U�����]��g~�cO\څ���^Ҭm�4�vZ0i�0O�몊
<�<*�gg&��\�}�!"D@27�N���E̸<��>HK;���t��No����y�Zj�;<���H�Y[�'���y��E9{s���у7r����T�~Kh���v�h{��f�>��������߻�z����ú���XN�0)�pT粳_ny[���\k����|.�(f�7��ց=�P���r��[,a`{Oǹ�7�Z���JQ�C�_&&m���a�G7�(����pz*�����ݗ�v�v{c&��e�KC��v���u�ΔM�iw"����\]�nK�W6#��n�����D��`GV8dU�4vWKݷ}m�>��܎d�7����^��f�j߃9��>��֥c"���t�>���<g��K8�Vy�ڮ?����:�����D��X/k�6��[y�uݞ���N�x`vՏ'�����.
.)�����.���iKR$�j�K��}�1wy�5i����s:�;����Rhv�Y�A���r�0���&$��ۂ��w�q�滳��<���V�����r�K:Ġ)���z7��{LԨ��U�^r����v������u���{�+�ן�5���Y�]�W�v�gJz'3��3���W�3B��=���;��E������,����Q��[v�7�Y$��&泚�>�w���5��X�ޟC)�<���=����?,�Um���̍��Y� �yI8{�D��-CI�¨�uݽl�{uo5T��p	��q��u�
�Ѷ-�|�<�qKf�C��*r���]ƺ�a[yK�/4�Tn�����n��[�{~��)�O>��ph~NOgs����T ��M�hK
�L�]�O5����
�1�u%���D����7ض�������)��]���/��/\����Ι��;LR�M�
�.��[�bW�ko�[���c��*;��nDm����������X�^��m�[sc5�Ge��m����*YIE�[���=qze����`���F��&Mz[Ūfz���=������x�Z��P`d����u0���6�$�	^����~����NE�6���°�0�{�6i�Y){�����5�˿_�"�?��!I)���,Noy�G>�ob�7�~���^]K�{k7��C�����I��mnXB�%��E<��5yz��_d�q�? u�zxx�\�ͨ書fR�4�T�� �F�WZi��T#��c5ۙ�k���R8O�ݼ�Jd��6�t�a��X"l����9�sl85U�&z:��/�;��p������ɱW(�e	����lO:�V:�V�ry
��S�p:%�˚uT��ҟCU��(��J��t�9�o[�r���߳��|��H!I�݈�ar��ro�k6�
��|�b�j3G݃
��ԈX��i�W�k~�4fW��^�ch?Z�qzg��.g�����:�6�n:js�Ûc*|&}-��7l���s�����f{��@o;�|ݖ~+�nWme��C'�z�s5�};���Q��צv���!ylC�}^a:F���E�ޱ�{�/��j�~�)����5�D�A�sAHˋ>�g��]1D�h�Ӄ,�}@Gь�qgH���Uh�Kq#S���޸ik�ŝ)�<.o����/  +[&9g�:0b�H�l�7+�H�%Ӻ�����ç���cu�s��cI���0<N�N��nv�1�v��}2��ͭ�WN1@Ɋ�s�N��~;gퟎ��q�ͱ�g�'<n���%��O�h�v�Ioc\Dm�a��VȾ4��x�3wA�x��<pyu��۶W>������1�Ÿv���\���D:֘0��;)�m���K���#y��4���ݓe�������1�\WVʹ���=�=]�+�n�H�������s����x�b��댹��z4�Ɏ���v��!���1�߻|^�s�K�M����"ӄ���Iϝv����{��ʚ,t���V����O���0�p�'������K�D>�Q��uc�SKUslNgJ��-���q�k}�d��؜��y��>-�~�p�6�M=h[Z{����?,�)�Ԓ�ҷ׵+�In����m8BM��{#GE�U��P��o����W�D&��A�f��y=c)d����Ekw�oi܆��<�W� ��8�wL��ky�r�j{���TTof��Rk�ժ�\CY��s{}���g��I?l��)N����fQ\<4�#�[�v�:ݬn�6�7b�c"7��$=�� Lb%q�6ܴPbm�д����7���>��/���.��~��>+�u�{�v����kP����ǫ}��&�+�a��0�B%��w��=Prz}sF��	Vh�G3K��ƶ�̄t����m��#R��i��;���.�ԝ��92�'){��&4�5U8`��Z�b$�m��1.��J�Mn� ]�[���ǀ��t]�A9�n������P��jw�����#c#*e$܏�����t�0���#c���T�G[=~�3$�ۡ��2�s�}4���yJ���/��c.Ù��g'/��뇽w�R�.iP�ɭ�z�\�27�b�uR0�ϐ����뚤��ʚ��u�j���R�5u�쭛�x=��qjE<�SW9�j*�^��R����~R�����/��������M|��"���~����V��n����p�qۋm7<��lպ�vrP1m�`,�o��f�����!�LN��/{1c�O7p�\˯$�r�{J�E��X������{@��}����UA���$�~�<��\��a΋�1y�ĬݓL�~����I};ÐYw�7�}�n�{��+���lVs��y���� �4���>��i��������č>����Ew������{�k�>[��e:��(u5j��w_>˷w�H4����{�b���v�ْ��.t�7���]l��Ӕ����ks�6q� a��<͋��窱GQ�P9�x��nM�w7�Su�b�`牥!���A�X�Ns���fsK�rvw�u�DՐn��� ���y�>� �k]�����{����n�����X����G���o��
�OOm���ێ&�$���d�7g��{/$�y�n�娍��8=�m
88���p+����"�g�����r{�qx[��כ����ЪS��{3�j��}�{��k���'=�N/(Ԉo��2�T3��w��RW}����/-E�7������R;+���^��_,�0�W~��2�kj�^�£Q�_/�DW2=Y�:}E\���<6V�p����:�Y��l�nm�؞{J��VD~)��_�Jњ�uI�O*}�o&ͽ����#�@��q����S���������Z�2�%b{��d�FT��6Y�V��x�]���+Kr��1gC�.�G���|Z����s[��(��rH��=�;����Y*%��r�w[��[�̔�=o�?q�g�Kiε����z/j�+s��a2.���m<91��k������3����z�H�N�<Tգ�r�v]�Y�ib����1:;$����)F>���罝��,И�|}����u�!�P���^�)�3��*��˜���"{�=��=�wsvz4�� o{�=]ף9w�n�p��)^����ª� Y�{��b��M�׊]�݁��\����XfU�u05��7o3o��=����wy�2���[�HUW�{��e�Yےͯ{�Ŭ���+$�oc�:��W�S�`s�_����`�������#�@~7�axR�pn��lkw���S���瞯����Z~��\=��ٜ�+�2%߰�o�B���/�f4$:����G��n�O��$�3��,X�K3�$�1ff���/��Y��1ff?���ĳ/��KX�V�bY�1$�ĵ�X�b�/��f$�1ffo?�}X��ř���X��ř���ř������?����X��ř��������������K3�331,�b��ŋ�ř��/����X��ř��_���k���ř������?��혒�ř����lĖf,��$�1ffo��Ifb����V%�fb���'��-����j��$�1ff=�Ifb���g�����Ifb����bK3fg��o�_�ܫ��NLĖf,�ɢ�q/��?���$�1ffdر%��33������
�2�ϼ-�X�������9�>���w)�R�N��=�Wamkz��] ��ݤ:��lzK{����Z����;w)�wn�%��Э���Tz�O{�x�� u^�B���     �             @                 �       
 ��RS�8t���`{�m��0=�+��m�{� wtҐ�0�b��ǣ�`�w:R*����)�� ���[���Y--�������ԭ��y�t���w��u$N� ���iz�טw��g���w�����ח@�� F^CݼZIU���y�����^��o8u��}h{ �ѭv_      @   4���κ�0� N6I{iy��@� ohH(�x � S�����=���m�vQTlR�S��nc����y� �J ���@�E= ��P>쪭�A9T^}é%$^6�O0z�֫�x  z
mV�9=�΀:o0h����]c�м`5UD�A�� ��(%"����yd�"�����WZ,�4�hlQ�d�ѳDx 
)*G�         �׮تx��޺M�y�Oa�=H�-8��$# ��c��
����n�+���������  z�o � �&��A^Ke
�۷�
����Zc� ����$���T)oy��٥q���k�� ��p�o�b�p]���ҽ�z��Qַ�ݪ�����;t w`�         짬[oo.��{�����޽��y@�-� ������=����l7����c�[�M�� ::�&�f�<]U'�J�)Hr�هy��4�b�  �ΙTW���Ԕ{����EŒR{�w� ��� ������;{m�[d[�x�W�x�*�	� ��(        n��'<L���(��� N��;���-����F��1�� }��n�m�o]����w��X��iքA�w�;� �G[M���q(�\Z��
*�P)@� w�r
��nK�nB�QHy�ީP�>�9�5>3U����|�%��q(��}�x�^�4o�uǀ w���A����t >����ԀW�0t�O_s�3@�;���	�)P  �&$�*   "��jUJ4h �تTR�  ���	JT   4�T���MO���?o��*���?�P���(�qn���󏼮RwMJ1A�����a%	%}Js'�!%	%�	D$�DB��%	%��JJ"#���$�DA
BJD/����g�_��FT�M1?ȼ���N��J.2��m�eb�r��N�EO* "kw��Tw`ʖ�JHZ�:��D��P��`�J�>��������S'1�S���EnPh����S۽Ǩ�������uY52�[�f�ͺH���h���*{@h�;2��75w^�+e���׃����R�4��ԓE[p
�N��@�ݨ7v�x�.E��7`�#ה�nla�4�T)a��,T�����Qڹ����
w�W���c{06�:4[�G�R,�]�2e��e�{�%��iiǺ�of��<��r���Tہ[��j������Qۤ�Q��������+��]�D�6��D�dcrM��̻{P���eK��j̚��ǁJ�����'M{����o`�]n��wQ�����ȅ�+�i*-�Ug�q�D �"vhq��n�v��BL�k��١C�ڥc/#�˅�[P��tlaڻ�Kp
��S�4�hne�*��L���q�͑��Ў�SM)umK:Wyy�����1�I�p�����K"�{�X�a�ˎ�/��c�oskd7�������a5�Op��X���zJ�21긒��&3dKe�ܶ�+eo%:�X����0��:Y��^˺�7s45�y(��`f6��Bβ%���	��_]������ZxEmi��[/c�Q;��ddN��YV��͎�t(���ւkU�ݒ��B+�F�al�vb�<D��CVg�N9(��+u'v����ƺ�{[3#�Άrf㩭�i����#��I�M��X�U�;l=eX�K�N��3SB�0�b�fY�Q�,mE�j��� b��$U�*mdN7i�d��! �.X�N1��;���^�:ܑ�j��f�5E2S[�&*��*�1�2��Tf�UGQ�$���xv��FV�!�$�I0M�8PZi;7�Rn��T�T����>��e�8e�v�t̉�(d��!��R�L�Z��(�[���6�yyX���N�L�M-sbQXj� �'i�M�9�;����%�R���5��,F�4�=-j�v�3�]��M+oS�7�+�Ey�*6��̦(�jgI�O70(���wxB�����5�K�p?^F�ث&��yI*x�i	VԵ��k�.�{(�VI�d�S���e��^0�ұOXU��k�W�2	��5�Kjq8��]�����(���h54��өw,�NQ�x��i�>0��;�]EW��[J�̶r��śv�Y�.�L���C)9V7æV�XvT��6b b�MtÕ�&�ג��� ^�ૼ��Py����m(4v\�i�˃͕�s�)���%�y��@��l��D
̘�TS)X����M�JȔ�w�nm;�.<1৒�-M�p��69�,Z�i�IJ�O^���L&5�k��{t!��c��t�[YSu��f w���E�ځ���Y\V^�'
T�a�Hg�Zxr�n˭��j0QsA�r,��N�`Q?P��%YW5���w?0+�&�
�d�[Jk�� ]dԆ:�����H$��D5��J���^�r����KGڅ3�S]J�5*j]���8��ցJ�([�a��+�E�R��IBV��Efm1SU2�#q�����0�ٙE�z��0�u�'�JQ�i�x+���Fڗ�, �6���"�ٰ.�ߛ[z��S9e��Im�|)�d{8�r�բ�庵nn,v*��wW�	�-����)�� ��g!@�� ��34�}��9գ[���;�E���#Xj�{*ސ�ܖd��vb�;����p��.P{�@�{j��b#� ���HM��Zw5���i2Aa�����4kv��wY�k7p�S2YI͈��SF�m��\i���-u��m>*7$v���5f\����ц�l�k���]W�tF-��'N��T �-xj�*��5d2�*M̨�r3]�LF��Sjm��Q�IWO2���Zd�D��h�U�]<�v*�l^A����^�(A�os -͸��Ĳ�Xܭv�Z� �BYP৏�@��4j�2��+[�%#)�is1ߩ /7u�%�S�آ;{�y�{{9��L�o�
�W���B�7�Ƴ��w-a��U�O�gͬ.�EJ�2b�y���ea�S��R�X*�`��fa�"�����̮K�;��\S��k��[�%���5�
�������f�"�:nR�1�����q\� ٕw����/qJn:��{��x���1�QPl��l*�.b++t�-��#�6��&G�ݹz����x����&Ga�Sx�X���D�DB]��W8��Q�$�J���@Si?��V#�t\9�#Yf�Mlz��q��*㥲l֝٪��6�D6�f�=��U-�S�'����rhT�%Fq��E�������8�R��8O:��-:���u�U�� ]e�b�I�n����GdJּ�[u/4��qd�M�v�Ƶ�1�·V7K��Z'Xd:��##h�����ȭ�a� j�#�HL��-]��n6��$'sC"c��Z�ڔ-1��+#���w"$�4nm3�P7nZ��r��3Xk7#ǀ��V�J�X�Ln�ygXb�f�U�b�Y˼�jE��≩k+ ƝZ9�Kd��"�.�az��F�γ����z�ך����2� �i?83�Ә^���u�&f5�2�����,�G#�ţU�\��-��6	F֐�9u�;,��L���[� ?
d��Y�(2\8��Z�6�u�V��4�B>��XE�m����UL'.�?+k����z=
X5�|��#.�=���r���Tf���t9�'*��ur���m|�]���ͻ���yhJ"F��6��T�^�{��bu�)Y`O�G�.��_dx�{��=�y}���>���֊^U���6x?p���	u��ҝؗ_�dBrӧ��	i!]���RE]����0h:PnBG�鎳/_����m��m@l�B��7��ul}1&�K{X@+,8㩌�v�13IT���uYS�k�dap;�n��=]Ξ͠�]���nn�7sj�H~z2���O��[j�a\#��ym%�VL�S�.IO<Ӗ����๰�$��2IR�鍙�֊o�`�=*0��]p��X����)r��Bۀ��ׄ.��1�媴nRy�Y9%,n٭���J�BhKq���$��4�ƣ��MM'��ҪQ3J�+�ߤgg��v���Q�p�`}�i۞!���dFێ�6����)�����2�&��۷=SF׾M�Z�>J@�E�d�vOƅ<�9�y�.��)�bXc�R�Q���-Ð�F"%\�ML�=T�e|pL����)�p�鈣0z�I��Ź!����7���|�5��
���"Ś��̩,dj�Q7��^^G5K-��qJj��H�7���:��.�b/�a�V�݋*#WxI�0��Z2f����6v�	��Ѹ�奸�m
zt�Q�݅�wB��L�,R��=ɦ�3��i�dT2e)��',�sPc++nm��*#�l"�5��\Rk�o�J�L���5�`lIf��X��������{{��ݖ�#,�B�Y��,�Xm�=CМ~F�L{sB���#d�\�'���aF�U
�\��^EʕmfΥ����[��m��V%hJ��9x��#��ltƩlJ���޻̓����(�kJ����L\�d�N���t.�eeٗJ�\2�l�@�ҭ�����QqQ�Zr[�������.�A[������9NV�[f�
�w�C���BQF#WP���5Bє��ג�ŹlDo0^�ͼyt�͉�v�DԗA���1b��i]cl]���J�4�+s1C��nb�����L�l6�h-[��p��[@Zډ�^��.��tP�T�-��:�8�TCwX�#՗��a����t߄�1��^ �ӘtN�vq�t�T&���ƻz��נ��щ�Z�fih|��ƂvE �3�I��F^V-l�V�Nb�s���k	��L�y����HI5���#�`�ӀM[���m�_e�Ci�%�"v�'n�ؖn�4s0l����. M*�zB�nbVC['�v5�񚗑��K�or��y-��`V�N�����AW$�K�+.�MP��:tK"�I����wi\��qX���ڪU��x�t�:��t谕2�ׂ�����V�I�`��&��yq�z��7e]䊲�����lq���U!ak��؉EZ6�:��QmbS��VV��6�:dd���2��HR��J��i��Ĭf��H)�ʓ��m�Ypn��VխV�NKBE[��&R��4�-�n��^���-�K#'f�,q�j+�DY��E�ʭ-mmZ��sU��r����F�Y�UR/��v��2�,\8���Ʀ��:⫼4�@�>��J�ys5�4��
�r��Z��v�tLEn��b�)��_L[(僗Of�
�+x|�闍d�j�7��/fZ6%�ͩ�݉�י$BZE㲍�7(��7Y���'@�0�X��fV=��.m������Nn�������oר&�6�Mo�p�:5TqܺVZD�H	�I��{�.YXjO�U��S��$�PB֍l����c�t�ڸ�ӻ��l�÷A����xV�V�!![��֬�x��i�&YU��ߴ�0���HK0�t�sA�&�i�㷘p�M��[{�-7��%x~��X�f�؛���� (�*�T�4S��(��[�"��`��h��^�p�E�#���dQn(NI,����Xl��F!��A�%�:0P�i
�u3v50�wf݄Ĵ�؇-Q�ݳ���-e8�ĮZ�j��TCǚ70�ƘFۺо�S1�#1U,�~�>�=h��
R��)6(�j^TT�x,�A���+N�l�DH2JKj����.���*ͧ���LÛJ�6��O�B��kօ��yWy����e�,깗7@���hHb`ޠ���2����L$܋\�reATYsW��L�.��ٖ�8;�q��V(�77��r�8�Π�)���N���U�N�¨��Dڬ1BL(��V��յ���B��h�9t�Wy)8����w7%3�.��\;�rӪŻ�T���%@�8��8m=�Nӵ�`ѿqZ��8!EdmI�N���c2��a{4�..�p��5�b�Mj�[��l��,޵�2�ܩ$řt���A�-3rkҩ�Zc����<�بf#g�3.��b�nnv����nS��(���kVR��jkLU�v��FU���W.��waXq�k�2w�4}�(��۪�,�[J+lX�fȊ��j	,�X� �P�R�Vkoq���&G��.�]j����]�Ky��è]�e�J�lQ�è���ʬ���d��ʭmǧ#w�C+nė���-����T̉*tv�U*��&LY)<��Em�1^�mN��۬n]�Ġ8����%�*e��"SB�T��Y�R����t$��s��h�+p^૆Bp��'5$/��J�nꉍ�Y�hwu7%k|�pe֍%e�,3MЩ�|����È�.Y�g�+���}xk(�	�*����Y��-Ȩ#`=��+!������{���[�]���dƮ�jX�yXs6���b&׶���9�ܐ�G�r<�������qw3%�<tvJQfT��n�=�f�҅U��e��eJ�`
j��dG�n�mk�J�bp�:��6�������y,ʬ;�]��f�OF��h�Q��V&F�铊�l�_������Z/�:{�%�w���Y6��YN�����ǆ"�<�|]9XW�.�����Wx��CC�,�{�ulWcV�̈́4�8q� o.]b�b�p�n"�uf����+����7w*u��H�NOF$����:|(�B�9���[�HV'�����2H�{;�߱O�ߛJ���A��
���6�Pt��'�Mp�L�$�Ay���d�6��i����f��c��SȎ����B�(\#H�:D_=�o	�H!V���v�#*aF�Y��yԿ���ڀ$-�Z�.�){v�6�- $Si7�ϋ۩g��.�TF�j��م���1U�3�M�J�k�
t���q���C�7����p�k�e��ba������`�k�ŕ0���җ�rr��x+B��r��`�Y�� �*�쵪\\�¼6�,����é;�]�.�ejL��o*�f)	�Q$e�AM�z���Ѻn�'&�]�i��6��t���JGU���������na
J34��Ck'i� K��w���8�;C��:.��-�U���6����1�kYt0��eK�3.��o2�n��`!Q�nؼ	w��$�71�{4S�[#��V�Ԗޢ��[l�ʔ�iVK��L����3��N+�[���n�^�F�cB�v��QИYXꤑ̻B�Hz�5i����9D�[X5��9VlZم�����j�R�c/j �8k�Í��e��[��PyӍdr0D��,ɩ�&K�ēLX����(f.K��2��^k��W9����[�I}7�n
�ŗ�Iʆ(l�um}���2t��͜]Q��9��,]�+����b�c���\��8w:�����C�L5�m=P�p+���t�^�x�}af��ʿ�����[[IL��>j��e���XV�V��(|�K"�x�W�$C�XDe3$��G��1�����(>��do�ɚu���R��7dx�����vu�S�ԀQ:�N�Zr����t{�6�c-����g-^�U�#f,Ȩ.C2�r�h�1Z�������X;O�P8��%�����^C)xڿm��~�hښ(X�6Lc2��%^;���:���k8ڌE�ic&�c�wj	&�i�H�<��\�5��ۏp��t�4���:�������*���J��j֬��uӐ@
���x�� 	�.ԫ*�T5U*ʪ��@J�]�%.�6RX7b��d����k��������eem"�!5HPM*�R��j��^YZ����Իeڪ55!JʵUUUJ�,�UJ�
��UU@P�۴ UT�uR��l�@HC2�@T	9D�� 	[Y�}�|G9��<;y�Ϯ
��R�톲q�����m�|w|�=�qwJ�Lld:{q��؇Gos����	�s+�^�����hx��f9-��j3ø��86�c���)3�5"6�p�����l�j�u{]�����v�^Q�x��i�v�gu����]��닌Fݏv���f��]��V߫�?}vC���l�-���^�� �`�Y���y���te�-��	pۮ6�-�	�u�b�gv9FM����/;��\(n��7���=;��B6�;n7O2�܁��\���m/v�s"P�*�Q�˺zy���ؔ�p�Wr؏WGa�ɞ}���.r#�8�.��+�IpS)�t-�B��ۇ�7�}g�p�3Ϟ��g�����y�ㆮ�S�ۥ4��n-<�Ll�2/��b��x뵨��9{7v���uz���'��=����.��3>tHݎ���}��r��ݹ���=�y2��T�m&"8�x�F2bM��P7Y�q���3�v��u\)��۱��.^�(��<^���͐2Þ�v,⭓j�\���N.7@���]�1�{u�#��%�S��4�C����7FL�+�pע��Ύް�5:ี�-cܸ��j��F0���wj9��<ɰW�'G���t���tc�eޜ99�Q#j�<-��u����_Iv�e��]�rqu����+�88��S[{\�]�o��|��\]psz^�ы�.Hv�I��:��m�G;n5>�O=��5>�۳V1<�=gęh���>�λn"�npv��ݹ�V�wIK��M���r-p&A�E�I5!��K��޶j�ֺ��}7vC���rug�La=�b�7�����ۥ���M֣n7=n#�s9�����Ύ�,��@��o7r�սO.nM�Fy���6�p��6ܞ�8p���ys�-��K�8"ݸ�z=v3�	�[�7o��d�:6���n훒�r��{=̮U����h�^�ͱ���u�����as	��w[/ϋ���뗭�^��nN�y��&���8��[���q[��ۋ\�:w8�۪��7_n>��rg�Y�z2�����u�-zjЇ!RD��;����,�v1�����]�a��;)�:�m�:���|�r���`�Sܠ6�m@��G�C�^X��wk�')��a��&۬��8zT�r��m��Il�c,𦇝�W<�e��}�W�����vz�����LOnދ�p�d0%Ƃ��Ӗstg�c\j��'Z+!�<8�ˉ.��^t��o��y]�:�v۝����(��V�$m��]&��ñ7n�wZ+J�G8��u[F[n|��WHz�ם��qܞ�-� <\��v��X��=�ܝ���c<�����ݵn@ړ�\�r������vX�gx�۷ Z�"����ǧ����K�����ݎ������֍k^��w���7km;��X�;{�;;�j��ax���w.z�퓨ݮ��6���i:3�n8�a8ϵ�۩6���붓@���v��#�l�`84���d�5(v@Qy��ql5gI�;�[������T�:#E�����/0�ٻ6v�М�I�A��p�"�;��۫��m�7�����d�#طF'�a��ώ�q��뗤tO:�#��8<죣`�q���^{����r6+�d�n=t{���x6�j���p�X���v�9�J-6kqڂ�h�:��ͦ��ާn�֮6�Y�m��9;t+tNq��[�ɻ[���-���I��ݝڧql��= u�p�|�7jV�n���p�m�M���xе��cus�����������9ݧ������y���7����ݻulu�5�s��u�ٸkƵn�g�c$�v1;e��`��p<�WGd9��vGن��h�;�/!냥�����6I���>����x�4ov�ڎ�b5ۣΉ�Bb �?QR6���Ƃ9��7q�M�;I���ɶ{ycq��v�"sb�r���N���n&��l�2��'�Uv��\pZ�ptus��X%��w'B�O�y��)�V�tN��f�8 A���R�Hy��x��9�g0Og�z�qv��������n;s��l�{ Ԁ�h��:�gPv�k�6)���%i�D�m��G�}[��mÅ'Sv��7�	�츺6��vGV����yFэ�Sk����n�r.�����36�[ �`��{lnbD8x�A��լ����%�n�b�3��j��x〹�Rv�@<�m��їle�w*e�]�e:ˉݵ�u;�to\8�Z�9��=���p)l��5����t���jLJT4�q����m,�rv�չS��g���@�)�ug��[����׎��7\��<�=�M�!�0t�i/-s�7�����)�ݯ�c���k�'n�#�86A;z��\�s��ogmm��ʗ�Iq�\�n[=����N�cN�].�u�]p,�0�8-r(HpX�6��ǪC�XX5\'c�1��h����_n���+f����b����*�hg�m�h,ݷmi���<xerv�W�n{����ayɝh�8��z�۶�N����?��v_�I.}o:�Jj��K�Ýga�`6N�7gnNX�ݝ��5�
ɹu�Ig����m���m۱����	�1���;v;Dn�m`�=����wl{o%�Y;m����"ٮ��۷�}�}�p-+�-b����ynϳڌt�[V����{��K�,�۵v�+�c���0X�[�pv�p��\����0�]k*��ˍ�ڎ8�x(E���ys��ݞl�z�۱Q���WC�=����^؁����rx�4l�������M��s!;&���'��ny��Íɰ��mk�M��\�u�����.��W\�o���L:*z�%Ӹ{y8�l걋�Wh9���cmy6���'E��8�ջn�ԈF�b�>������ل��tX�=M����&d�6���{q� ���2\'������`�<q�n�Ňd�yL�ǻ7�b��8��o�<F���^���u���w��棩��{K�zl]�7s�뗫���gZ�稖ngӹv�`+���;v�@alsȘ�����l�ι�R���r�Z�e��b��87Fuv#�E��V���c�G-]��N6n��>o�5��2nX���Z�n�k���v�;���o�3%c��ɺ˨���zj�1��s����/.�+O%���<==r�m�tru:�76��z\�F�j�S �Z��f�=�pi�X웈�6�C��\����!�v���p��R���.����:��g*�Ų�WMúq�l*v\����9�nv�m����n�ɦ���59v�u���;�^ݷ]oj+���&C!�_!�;�t�t����}v|��z��ŷn��L[l���mWKۭ:��m����o<y8�����6�| �Ln��'[���nV�tN�
�q����ę�6�-�G&x�}�@�u�m X�e׸{sɎ'S�b�c'-vx�j�>ˈ�uY�j�Z��m�ݮx�'��Kn�V�h�8k-�����_g����P�y2�:[�8;n�EÔЎ�3�2ql^2<�j�;/�mSd�x�ڮ맀�[tJYGnݳ�n���ݶ�z��"��N:�^��81��v��zM�O��:���s��<v:E��es�۰��1mb��-9�vm��
�NK]-n����m�rv�3s��뚭�,�.۷�zݮ����u�`��&��C����u���p�s�̺�6�;!�>{z[w:����N�����2�޶C��ͳ䒂#�X�#��a;Ev;Tv���}�oc��6Nx��ܫ[\������@��H�<�(��Cm�\�b�[n;\u����m�1�$VsaCn^��z-m��{Me�c�q�Ok��d�t9�Y�k����6�t��b�����W����ol�냛���8��+�ďg��C
�L���"���Ɇw����^\M��vNF�q��E���krr��e@&���u�\�)E�����s���'DO���{�e鍝lQ㣠D.�N��ɚ�3&ў��n��wlq�Ҽ���֋P)G]�lr�u�4��Wi�!�9�n�{[�qu��^�6�)��;�lm�p.��<���������J(��lon��6H��2��oCΖ���"@㞑���e�ݼo"�[�lmr��{��<��n}�I�`�:lݱ�����ڮ�vc�6h�ks��z��9^�N8�ض�vKZpv�*s�ƻ'Y�-�x-��+�!Wi1�c�1�3�g�68v8�p��QZ��of.�\�\�9@��;OnɎl��ݛ�	n����\<|�w�d;�D5\�m�0]�ޏ`5<�a�'-�ݗ�5�^�v۞��X-��S�a9ً֪v�6���D�v��Mm�3�޹����[�׫���v��8Ng��úwd7;���Zvpb��iU���#���R���&޺���sȼ'\�޷k���v6����'[�N������R������޲�v�;6�m]�ٙ��v��+��c�>���y��n�=���;��q/�]L�PI[2n��u����F)Q���w�v1�'=�^Ԁ�;pn�=��u��MI�@X��']=H���`�x�wVK�q���it��s��8�֧��vզ�������-�u%ی�j�ن�n��E.6���uƄ��<I��9�tn^k7c&(��w;���=��jBnAxw]�m��q��8�`�K�w�a�lK��]�;u&�u�����v��sV�[����$\��ݗ��\k�n�{9G��������Tx�Ƶ�;�wi���,������mל�s��p�۴�[��d�[����[n��b�y彺�v8$�G<k��h6n�a8�u.k�bP�Q�BJJ"#��IBQ�?�IBIDD	D8I$�nT�P!UJ���%�R��˛��"`���"�U��,�.�l��$of�s��m���>��ۜh�l1ۄ���=F�7g�뮸z�t��s�6q��&�:5q �ɱ������r�`�-�z;yN��n�����K��gn�:�Ր6}��6�'9�z�ܝ���+����M�m��^{W��t���Xεɷ�r�.{m���MɌ;lQ��@����k9�䰧m�3�x�HC���+�v�8�Ã���{�0�;���G]�g�7=:��N�T�Ɠ5˄�x�a��&��u.FK�Xx��]��7X.盷F�kc]<��k�:}��Ż-��=Z�_z�D�8;Z�ۺ�'Q�Eq��<pc�IAI�� 
o<���P��[=���Wk�s'>s�.�qD�S��pcl���;<��Ek7�s����厹�;�@j=�/���v����J��;���5�Gg\���6!Sq<�So:�FF9`�>�r�'��â�sؕ�7]��n��O�mX"xݛcz�\�q��l+��G[���$wk��]�z,�v�$N��>A�x�]��b�*:�wk0Y��ܥ��ѭ�z�ׅ�4l��w�-#<��G%�v�9h,vj�x�s��c#r[�8R���ҏ#��]kv�z	�^�m�×�g7�U>�6.��$n��e���Ѱ"N�˶K�g�<N�el�WF&���;��p�yNĉ��Od�!Fή5�x�����溷����.m�<x{#�����f9�5�յ���r�h�nk�wlՌ]=ly���#l�q�m���ͮ��+��Cu�(�!���Ѷ����
G���r���uNGe7C;l���y+�{>:��q#�ԛX�R��뽰��(�v��#��>�xP0Pq����[�u.��3�C�w]�ݹt�^��*`y9�rp��lF�e���*��p�4���xh����讳���^��á�u�ޗ��� o�Sv����]b8�KV糓d���[��g��qJPʊ)���	D(��D(P�Iw���}���fvV�������X룻E�[)���q�m�m�vk�nI�vN����/k�V,���9x�g��Y�ʞ*����Lm�lnz�����g7=�.�S�=�q;ny�I��L�����5���s��:.y��It�s������OnN�=���ۓ�{�����m��5׋dӘ��l�v69˹ ,�'�ش�ɵG@�ۯw�����ðxy��Ȏr�쯎6M����E0p���d��4���JQ?���������o��B�i�����2���ͮQp�;������/�R��"W�e'���mمH���#)�=�+=2��l�pΪ�̸���nءk]ηt(�t�W������$~�{���^|�F�NG#m#�0ma�Ǽ��9��=���T�k�}�ye���Mǣ�T���ܫ{c�U._c��6
�2�p4An�o���2{�R���l����1��P��"G�+`3��Lʶ���z��(wj�ak���ǥRʛ�8ڌ�Q���4�s��UZV-���g�����ݧc!�p41ߍ�6�n�j�_ݞ����m�˃����lX��8�%-!��tu�����3�v�W��x�n��컮G�������&[���J�����s�=�Nu^�5V¹v�"�*w���J�u�n\4y���q�f�X��~��An�����Ȫt��>7�.0�Е��Z'�Zf{޷S\�<���Q�n��Z�/��E�:��dVԣ��Y~�K�[iz�sl1�a�o��A�E��md� �S]��j\ѿv�-��a
W�k-�=~�Xc�a]��ul�vs��r��ឥƺ�'0�|J�����x������S�{��_>W��<E��	��x�ޫ��+}r2;K6Y�oA����T�`�� ��TJASne<�3M���O���%��x�Y�bN��bf}V]D��@׾�KA�5��2���h�h�\�Ve�O�O�G��F�dd��������:;��j��f��z���F�t�υ��aKe��{��ǥ�^ P�����Y$������ ��x�9r�m��h;`�׶�j���ӹ�� Trm��7'j��D2���\������լ���>���n����۹�u䙛2x�4x�hG>��ICp#$�O��/w��fgCҒR��9Ӌ2
��/U)�+]��]B׮�zry^��<������0����p1��u�Ɲ갱;'��b�H3ʟ�׽�[�/��F�*��0
��P���V�5����g�!W�_f�ƪ:qbzJG�/JXrm���������w�)���9S��xB����b�R2܎Qx���ݽ�Zۤ<�i�l��8�s���s���~���7Lҹ��ݒ�v�2f�[���+V��,����d��޶�u�q��C�c�Yj��f+��#���G�Eh���.��;�x.|\އ�qݖ�'�ϝ�\�.�j��;�����2���_�Bs��8��R�%ћN��h׵�A�0��+���M&�rAޱSe=F�B��+~�ZN��"���{� ��M���+lb���wDo�Ġ�:΄#O�LB[�pvY�F:�1��,tު3��y��m�k=��k%k��M5m�WK����VG_��UO��ӷ�9tK��q�����n���N�s}��6iZ��a=�W���B.Nط���2�ݾ�IzS�˖,�ПĐ�	��rOw(uy�kۤ�;2���h����z�{�e�X��=�n]���Yo����rOE��&e�����,-�Y��@�� VwCLx��K5���R����+��CUl8��]��*��E��A�W'�{�_�%`���"AFH���1�}�*�>��
��e>�"�&ov���/�Yq����`ȧ�}[ȉ̛�$a�$n=9���#I<L��sSg�����e�PfMǣ5ͻc�5ۉ[���;[��zLsu:��v�<�ӝ��`)�ߡp	m������w���nI?o5X�Q�c���>�m�o�ٙ���uw��DDJ5��Ap��M6tҔ{'�[��,�X�Q4M���1^�i;����7+4ZJf��'C�^}˝����x3�!�b��K��"7Y���OyV�����g�ֵ3{�kS(���a���$�ɑ	����3��b��������qH=��W�Q�:^��S������{�JX�\��VUb�ڽ�e��/-�k׭�)(���\ic�3ڐ��/lj��kڴ/T]JD�����]�N�������[��م�lo������.<�xv�s�*�/��P�>j�楯C��e��^Zck#gB�i�GQ��ޱ��yJ���c��[��O (�����z����Z�`������bW�e�3�e���g[8v븴���y�/q��ۈ�-�5�'U��G�@��ȏN�GW#�+o�ZO���g��m��)���xvN�v�B���9{:w�	�u�;X2$�[9�<T�9��6�W'n�@X�;y6G<���pu� ��f���u��zs�]qO6�����a�\�1��=��=��҆<���7<���Itnz�3���7��q
�q�f�r8�&���ӎqf����tS�Q>K_X�fI�����Z�;SgZ���0ռ�����4-�a��!�r�G+�ڟ 9��*�t�v��IwH�Ǿc|1=�����G[�[���a
���l�8���
b�ӣ����i�0HY�7#��I5�i�A�vש
��{s��u�N���U�N�41�����C�?I��z{}Ux��1_	R@C�6T�/̈́���n��ل��nv�U�X�hOx��I��]��Cܝuo�igO�V��nR5D�D�;�	&6��}"���{/W0��b���O�1�\�=[�+�Kڹ�,�Ώas0�e�+r�N�}����PVZ��	�F�:�[9��h@n���깽v'&�8��鰧�q�S�j��h4�/w�Y[��K�ݾ�cW�|EvTJ�T���6��z��W��{1�hn�JT�BS2H�0���;ds\o�'pW�d�X]((�vvY�a�
p{@-ҠgdW��u2�k�AD#�޳xv��T����W���ܵ�N�m��,�p�}��]��b�N�jŏL��ȝ�x���p��I.�l��7�<���ή\Xvsz���W�4��u7�=��y6w�>�e	�Ҽ�>��hk%�8ee�k#�](w��D%ռ�㔤Q�#��!�H-ˑ���(��Y��w���Ox*s�v�����$Il���N�v��s�]����o�_r*�z�\n
ή��!2�j0Ԓ`5�٦4`)�>�����q�n-DU�k2��N�W%���}�8�&y�9�m����=YG�l
��2�M��]�uKE�7-u��f�y�f�k��ٻ<�f�,���d�cUV ��W��3O^Y��*�,��N}�v$��/w�e'<�{�*Z^�%vm�\�x����QQ���?�p^�t�����\���{֩��"���N�"���I�������R�T�3�:z�;C��Lj0�\��ܒ��E�;���=20���s�Y�sNC�O��ע��6��^T���hp1��,��C�j�owr�4��U����+Ё)�!�-
�vp���:�wCu�)t��7������Wݎ��e#!G�6�{r_>�5qnנ���ąF!M�=�tWr��+1�t�V]T�P���`<͘����wD����蹻�0\�v���$���w�M��i�J����~�Z��t;1�7����Z�;��.W[�(�e{{�)S�����u�?aʔq�z�b�.��|�;F� ����]Ʃ.�ۇ�C�6ޮ5ىm�Eq�Ηy�)��R*�6knbi��Tg�wٛ�( �c��k{P�\��#���W0�����^)���n�K�D�[8ah�՜��։;��-Ǉ#ǋ���L��t�.�;����>��N������N^O9�L�-���K)���:|���Վ��K(Ae$�z��9��ɵ�$㚯���_�uޖ�ٱ���M�Q��n��6�_��p�y�+��r��Oو��koküh$��e)��+ɛU���еM4���y���I��d܍��d�ѩ!���������𺞧��Q�a�����}�rN.�7$j��v^r����=����TlޱQ��"B�Ĥ �&�+|kE�yx���d�c�udN�dkUX�]��a�5��`bI7~��;�Wb�!
�>%Z�����f���/N�^0�֬�+z����{N��z�&�T�-xYL����@*�آ�'�W�����I+�*x�S-�߻h�E3X��w��{��Z&z�|�|�o˧�eiƜ�V[-ɥ����U�#�0��w�� ��۷�&��Z��-	Y��==�K<����C}�l<�x'g8��ahe���[q��
�H]��pη�'^�����yB�gӝ̆ft�	���T5�=K�p������oJ�a�Pn@�"�I��A�����69^�6��_i���]�G���ie(~�����u�q�h����B
Б�$���Bk���3�"�ǆ�Ϸܘ�꧹�t��Z���X�+����N��)�
�z�����e����M�Y]�x,���|b�3q��nm�u�����«��.mj�Ǉ!��|�_m�۪o%q۱zu�6�j�,�A�Iv��Q�6��4A���cn�>.k'��������Kq�9�����*�ᶒ+;��j��.�a�yr\�	4��Z��V��/F�f����Hv�/c�.1�n�NX�z���0��u����gE��iݦӲ#�>��/on��۶}7e�uM�����&�`�N�g`fp��p&�9n}�K6ȭe�gg���s6$9b�U��N����O�^�w=m��ؠ\b�o1����\�K��a�ӱj����ॼ��������ұ{���a�3����)���]�V�u}x�p�*�蠼{k�("�(���	����/s�>��~���:kV��I��4��ʗ��۪'��<��-����݂�oU�ߖl�n ��D{Y��� e9`�H�ށѦC��̛;���ܯT�����[⮵_��
�XKˣ[���X��Nm�D�Hl4Ti��M���t+^$���	��V�N_`�|��Ԣ{z����e��$��x��݊����_����iF!ƌ.9$�p"[�]�k�N#��po#g;�K��k�9�ėb�rD�����_9̏S׋�=[0>�I�e�Q)��a�h!��r���7�m�#rⓃl�n��Ἇ<�n2ձ�I��ƺ�
n���+�G{b�rQ�h�SZ��q�u�U��w}:R̶���kzo��.�s����s�Qk��l"�2B�z�#E���f%����i�3���Cj0�H�"��/6�6�̹a�,��}�)U	Fլb��kڭ!׽sAQGc�,���;}�w-�w�Ǜ�<�����b���@l��D���g��.�V#n���.!�^��oHd�N�'+��@��O0�=)�MU�T�Ìw�v��+�8Ef�<v��J�~��w�����7!�r�/;#�ٝ<D99*�N���w��v,y�A����^�}��R��}~ݱ�`�˥�ݓ|�3�e$V��d�����ڌ���F�d�ͥ񀈢1�</M�����⋞z�o�9c�WW��g�ٓ�z�ӷ4����=j�����4w����p*�ȕ�*�N���d�Ӊ�ft�K�4�.ְ2�ŵíi.9㶹�ĉ��-���G�e���K�a��ޤ�`�Ei���wڹs���aGK1׌�J���#��[�A���-"MI�B%{;��{eR�&�:oSC3����]P�E��ׯ�ο\b�d;o��@����;�}�4`��-	�f*.G�-�/�dF�mu�u ����0��Z=���WMN�F0���Ib7cD�vʽWkV��à)i���*�;s�,�>�/�4x��p�2����Qqk�.L��Xj�ir^��	D�Đ�[.���Y�ws��$
;�D"v�]���x�����ܮʦoN�ޢw̋���l��[<z��"}'0I�*m�ĳj�r���eq���k�,�zz�ҭ��4�77�X�s_v;y7Z�*\��HڔmvB_'W��:���}y�QD�kn�-#�[��m��[��G;&��r���	��l퉅e�h1=��ը}�̲t��J�^����+����K��Oo��܈)׵�s��Դ,�a���W�VK������Z��e�S,�u��WL�	��[�/�]v����v@ ��ԭ�� �4j���j���b��mD`���7ܬ��&*��)W�t�4����㫖*(j7��y�:���,��j�����0?5:��K�r}$Vi��}B$�򨍺�a��V!�eLLJ���KN�I��ϝjJ�0�6��B��i\ǯ�/��N�W��Y�O��}�d��f�`^��8��u�n�S��gp��:ߝ�n��c��M٫^���3�����f���R�6UT���+q�mز���	��B�q�CY֩:�um����d+݅�w6�T��R�Ei��/nS�t�\l�cV�ڴU	v��&3��α]o+�͓�m�ht=��/v�f�sq��>��v�r�y/x�����#�6�p���X�^Τ_=--�E2�wrb$�fw>R�x����|��E��%��L��/�o�u��ӻ岙�$�^�'i�j�6rn����ө$�opw&:��,)ְW�(��VD\�1D�*8�	y�w�)|'���Ő���-	�5&א���R����0�����v��e2o�^�g�k���E�[ ����|�7WK��)SWm��=�O�/ri �wW]xd�I(UG%��veGN�9'-���^�d���p䪾�D:�]�͋��.�E��^����%FK7�ߟ�;T7~3>+"�F�$��K�RFgy�?i=,V��i�v��^���x��(H�G|�x����%V��a%Mm�땭��p����U�m�g"r_�Y�����ڮ��NӨ�+h�dg���[p�J7�sgEZo/ԅ�þ�A��yO�!����*��8�9��Ez�T�,�	�y��t}���5A[Ys��H6@������?Jb��/f�.}/�s�c���LY�����ݪ�D�]]6k��#�������]��ĩK#%Š��*���V��7�P�Q�P,�K$�B�,��!-F�u��ǁƬ��W7k]�A�>w��^�M#P��h��m��b�(�^�U������ڎ�Q{���&eZ��VE@N���Wz�\cr\�k�����m�$s�lJnd��K�7`�pe�~r)%m�y���$mt��l�'�`��v��ü����6�Ļ�YƦu*�t6�^�ў�Թb��<������9 ��Ǚ��ӻ�-���@��nV�o&�mSZc��6��G�̙�G��u�H�\��Ӄs8�*^r�!��b}�TQ�}�:�F����D�kˬ���>�-�ɮhV��	�*����A�J��a�.B3�*q��p�mɘ-�5�H��v���ֵ���.�]�\h<����p�i��
y7t�s�Z(�_M9�ۢ�ߤ2?�b&Dq�Z1�ym
8"����Si�Oo�}×]��|SaU�7�/,2N2��'�.j뽐�gQ�O��s1�뮗�u
Օx㓵��~Ũ�w[kuKy{Xn�r�Vk��,خ�9�*g��l77�]]��],�-�]S�\�Vg.�=]uVP$�]sv̳�=���A���n:ľ��n�RG>��n�l��,���0�q�8��iޞ���xwl˶I՞Ľl���v�rqnpu�dG�
�ۂ.Q�L;���:�\m�w@�7M[q��`�$��n�@k�8{Uk���d�9���y�j��c���>�\;S��Hz�:�%Sqۃl�\h��s�4m���v���xd����l�v8��bׅ���<��~�7��q]t[��Փ��h���s�ε�a���}FC
�ݺ&��Ҏ�^���q�e3/ue�S8��'�~Uܞq�jJ�V�e[u>����4ݕ�5���0�Q�Ǔ]�`V31گ^��<�F�f�_y�K!M圶�������Α��y�j$�!cp=ڸk��X�{:����j��0/�دi�>��;����U�0!:��d8��įJ���e��+im�5�3-k_Y�\����^=>fFV��)�N@T�hi�Hݫ�`X+�틀I���=���d�t���q���%CAZ��1p�l��"�<x4�ǲ�*�7�ӵϟpjp:�bސt��Y����WXoˎ��Ϣ���!P,$l�'42|F-�=��ɒ6:�gF�8�]��ݞy���;\#l]\��f��\��W?��O��w%J�X���ɖYi��^a��+���Sn������E0rv�N�h���LF��$w���Ľ�S�x��O˅�{<�K�	��U�$nA�nV�v��^Yt��Wt�������:y��Vh��H�g̸sM3����3
jp�JL�û�f���aw��J�{����3[y�h��OA�ћ7=jyٺ����4U�p��d��7$����m%�%�C�S1nj���Y�����z��ʭ��Z��vX����0��u�۪\ Ja��$��>WY�b1nŚD�s�/�A^k�VҜL��@���M]�;�C���y=L��U�͢d�	R]���ιb˧�J4
ډj���)}��y���U���TX;�Adb�lݰʤZ�7�m{W-'oY��[@�b�I#�ђu�����R1�t�a����w&_5��휹��5��|���`����[��U���6/z���7$Z���v�D��҅n^%U�c�9"/�V�^w��y�j��V��)
,�.'"�#�ArL���~��21	�M�9X�I�����&�B"�2��S���|w5��œ 9�L�<�ך&�n2�p�n)�<�����g\=+�|�?YA-ʻu4�堋@��6�I�}h�	����K��ս�B���N-���J���'⁮�1��,�hCp ��Pw��ST���Ɉ.i�l�W����?v�����zM{C(��a��j6�ތ�,fS�e���vi��,͕Y{#	|FSY��?J���6�E��u	6�{,yyj���O�^��U�X��A
*-�	Є�� ��H����Ne%��!wi ^*�1Qlol��㱻��ciE�4v�Lf�w���h�����j�+CR0@��h�����n\�{��v8qr^�H����qڹda+L�Mߞ�]�ϮPGNf�5ЏL��~����� �m�����U�=N��7.xU�&X��[�,""j��K;��}���7Ҭ?A~�k�[�:^�mz��k����X���
#%��V٧��HEc	�MA>QȃR��Y�_KΖ��|X���ݞ0o��e�V�3V���%n�W�®[y0u�uU���f/�\-�P��q�v�`��j�������_Q9l3<��o,�NN��*+ov�d�}��۲����e�]R���)f^㫅�.��fs8½�K��}��X�0���\�J������9�{/9V�M�;�'(N��=��T�͟��:�aMF&�%�K�X�r��t8��¬�G��)m@��̑�c�yDl�Q�J�d�{;=�e����l������!�#Z��=y���bp$�5IP����Ʒ��G8�b�Dsv�Ku�R�nx��=0e�5I-�a$,�p/p�E���i�N(�tN��&Ž�M{<ur>#!�wW�ߖn�!g�l3��c��6�-��OI)փtjcG/��v���(nOlK��]of�κ���c��Q���p�X�9��TQ̪m�g<͗͢^���L�O-�6�|�Y�QrE�.�fd��E�uET�/�9Y��J�M���c}\�"�(9	J�%��@��넛ӈ�oV�da͒L�����l�����W�8+93f�=R�z�󓟒u�9�c�Q�B�
�V0��[ݕ�����7�7}��f̫���	��w;��؃�c�L�_M��y҉�S��^R�F�sޕ��ތN���[��N��G�n�2�-�K��ѫ��n�]u�Ֆ�,���h�1f`�{N�Va�������vN��[�M�[3�rd�`r�����/2��Nx,�>�q�bm�ojm�&PSVv�x7-��|��l���ݏn{Zْ`�[�!�Zl��83�5^'B�J�Nv�ڃ�=;��Sm�;35庛�O7c��b����[u�]x��X���G�p��pl�u�<pn�̥kk�.74�띝�I�t��-�v$ز�G��b�Jcu������0�\�r�`���en��e��\us�6��XU�.4���	7���ޙ��Ag�N��)pA~�}~[��s��u��Gs�]Ӱ,�}R��Q_$�恊8M��r��rc]�����jQ��6in�}����ㆬ�����ض��������dVҋe�fP��uo�a'���HD̍�G�U(}��Ы"�9>�dsɊ�!�NM�Ǡ˞?6VUϟY]���i9i�ɽy���RA-��
���������l�Z�v`7Yٸ�G{��[���fn��n�tNa�6�Fo�^����ʐ���;h>eC��|�JiH��o�����$�#�uN��i�{��̮<6��i�{�W����4Շrէ����ힿ�n�-��	�3n7F!L�X�R���0g��ƣu�n����k&��z���mܗJ�%���r��6��yF��~��=�{�V�{2H.�3=��l��}�w�r�lZ쉘PP�J�����=uP�Q.��e�r�Q�
7p=��b���i��0C(�&�����%<�+���t�s�i��ޭ]��R�_*;� �iVӺ�
	X��F�S����V?(q�o�����=���{�"P�������BЫƺ�����fh�-ZI�T
GR8�o��n��Yb�3淼��D��z�AvE�!i�v�
N��Q�)�U�P�̏�no�<�
��(X��(��<�3;�ӧ�mt��)U��aWe�_���>��9��
����iEu�ї������X(����Z;e��=P���e�G	d�n���ߺ����0��f��%��U_���`��"��ۘqf�Q1*�{�w~���w��j�DZU#��l ����wEڷGVݒ/�+a�;m���ma�ҷg�u�J1�%r^�eH�Ӱx_y�Ao�hrV��C�o}y%Q�ʉ��'R�s�ֱ4��AvI,Q���#|��j��ޟ<<�R�Z�/#�:���,�m�<"ړU�x�T��	�RЄ�>����(�@�B ~0�>�BB;$�ѳg�����ش�՗;۵Xe�F���*�E8,�8�r���bVk���az��˴�˖kj�t)� ���5Ku�5y�^-m��l�+7!�D5�`��k76�R��.�0�E�KrO�`����*խ�8��l5�#y�����m�{΂�=��xQ����F]�$�������P"2�o8���ܦH�wc,L�Ռ�>k1��;t�W�}<f�[�`��;Ƞs�1�}���1w�[�RNW#��������-͂���eX�N�7hӮ�����$��r�B2�P�����&�g�{�����P�g�{�]��^�Z�k�y�n}��A'�:�g�����Z�9vZ��c/�P\�t���(��gKM>�Omw;��|Q��{�qCE��ٳ=��$� �u�X�!�f��{=gj�kp�W-��t`��u0J�m��[N��<��sg�{w4�u�uY�*��[t�ָ���W�9w�uia��B/;������I+��/_ޘ�!����l�z@iYa��l�<b7�ӈ����y3�֨R�@��cCb�P���&qg�B�N�j:��t~�)}���s.���ph���ž��U��C7/��t�TCyX{-'�{h���i3��������?Y
(�8[ky���踟td+Ъ���'��t��Œ[�ģ�W��9�ף��pUjY8s�lN}�~ϟv�Bd�uXBV��,��[�^z9^Es�⽺�C�B!=j��ű") �S9}u�^��܂�RU�{~m�g�f�)9mCO;d�R��R6���Vj���EMoҡl�S
6�
'$�"�6�+=�.���s�7l	}P|�S�ݛЙ���ҝ\�ݽ�)x�!��nIa���,~�v��$8e����,���vw�T}~��ҫ{���[F͗����J;r���8;������4VH���I	�s�l�i�-�B^�R�,S���ߪ���H����?>d6aY`�^�j|�%���{��GN�k�b�p�o|�>�D����i�|�L+!T�%'+9�����	����b�j#�ݛо��������͎���_B�(f~�62�4HN8����Hؾ��LJ˯?]ZT{Zल���y����ֲ��*�%�)"���֓��K��&@/KH$���{�di
��kJ�X�Uc]8��p�3�3�� ڵ�������O���R`hu �ܬR���*��1�-�����.��TT��������僈U��?m��Gy��n�Z�A]������d���V�-��y�C8pv�h�y��u�U�9���!��M�D����w;��X��<�����r�=6;dk ��`�sY6�ř�tp��Y{}5���t罄<v��q=���oZz��1u�E���8� ��m�@}�	��Z{96�j�g@���A��7�4ԯ�kg6_��g5�&y�1�ud�0y���.��$�w�ԋ&�8"Ϭ*��ׇ,���v�QV*/顰Q�$����J"$W�����&�.Ю}�y��@"���r��f���9swZ���o>�Bp�#��>�6�pk���[HR�����3Z1Ȝ�$x��t쇪,�$����\Ҏ<�pJ��&�|N*�7�K�+Z骧�yye�ho*�!�r�N�ksvt�.Y.��"`5���۝���ٵ�d���}�۪d&#=�^d�5BH��yۘP&6iLB�ϩ[�N���jj3�	����<�)��Y���^�^��a��Dv�Ϲ��7w>�f�\�*�]e���ϙ˒���5��{2� ���n�[�M�l�|�&'��{Y��˴߳c HHJ&Y;~��0a�={8��;�c;xoL_M�.xLWU�͹.��{� +f��qM�Y��HU�.[J�YCEt�T��}ݔ.#C��ٛKM�ۘ"�����a���L�Ԅ��=�:��X������1*һl�ƭ�4`�-$�)K��MՊ^=\v8�m�;a�x�E�f�qn�%��ک������˜�lkq���ϜnA�ٴ�t&T����rw�p=��B�£z<Vt����e���`'�5���ػX�t��i���3{����n�wUίn.�۵�m��Ǐ�����"6�6�.�|�Y9u��A�tX�ڈ-��d�m5��N�,po\b���d�v����pj���zl�]ۊ�=�1���S���ݻ��� 8����j̦�C����x{*q[<7[2��x���I���m���㏷}4v#�g=	Hӻ��"���N��ʹ����]��V7%Ӈ�G��Ԯ���M��x};vzJl'N�!��Iգ/;msxǹ�v�g�3�|Tx{H��ۨ笉�(c�/��ksƹ����\[�B�g�xk���.���� s�;]l��#�k��X�1-qc�	�mv��.N�玱��s<�͸m�-ɵ��m<s�ݳ׆˓nsS��;f4��wW����1����nnI�p&y��{���{��w%���
ez�lt�ti�k�':�gi��:No)q]ۋv�{Z�x�v�Vݗ->�[����v��H+��۸i1�a�c�J�j�#�q�B�=�gc��N�{kn�=gv�<l��ٶ��s��۰���׷��l��f�pۉ�r���ϧX�7qk/�(}��b����� ��̸���6�k:���X7NJmv|�ۑ^,��Y]���g��1'G5̜��V��+.ڕ�����tW�6j �;f웮u��K��f������|7czְ
�������k��ן,��j��qݡ��
�L���9S(`�4�DR`�8����0��5*� uy���p�tql��N�ks�9|�q�M�V;F��&�yp1�;e����`#n�\v�v�\�!��,���C���à2: �mb��+\���o�V����� ۤ�v�^&y:����[��Ũ:��h���&�Wg&��Pi�\@؍T&Bհc��箱s�uٴ%�|��o���+vҞr]�5v!�\��Ӵm��<��5�z����d�ܼU7�uY%��0�ϴK�Y�7��������;@.�!.[�����ȳْU܂���(;��7�֔덶�h���uo�����x�m�T��ݜ:����[���[8y�=m�n�jɣ���I��u痶�N�ͱ�	�/�%�>���Q�5�����u�����R�n[����.j����|;�PI
�I�N:�nU��Oyt�d~
HRQ?8��Yi�>֨�v�]"������g���W]����p_e�����NK�ɿ]թ�軝�����τ�S�\��f�EU:��"M �Jx�}`��ҡ.�UU�۫#@4{�?^R�L�h~cX��P����������Cg�Z���L���\��q�*!1)$�S�ߪ��\4����u���}W�^���;8� ��M��犭�
Z�RR�5��d��x�=mH�����ˎk^��V4�"�u���&I�8�>_c��-�||%`p^-g��ZRi
Oy�v��q��n������[$@���@���T���E� ���� ���R��-<+�����C�_m^J�5Ь��q�Q�}3B���r�k}�p������W�嫀Z.5E	[K޷�u����c�uZ��#�`�?Y����W��A$�2�q�0�k��?yq!�|l�C�o��/��wJ��%32���Ë���d��_�� ����H$���a'�w�zɒGw)Ib��W���k�,�
FD4h�/Oi�r5\�g�ޒ�h6���0ιy؎1��ܫj�n:�67�;���Q��l��	%�.��ϭcVG�eeʺjDS���ⴙ���M�D�H����j���
���Y�Y�BR����T�}֫lz{)���ҡvZ����z�Y�Uɀ���`��k?����}��@.��k|�L��K�@�KR>4���ޮ�D"P�l�/����V�O�]p�=�V+��5�'gB�d�꾤־K�{YsMB�8�	����z��ӘΦ����u�'�G��9x�T_�e��z�LTa�:�9�� ��$TF6�J�'���u����ZBc��ED2�dm4{�w��^Z�z������-n[|��
���n�,Z'�_u����T��
&���Qg�'��"��F�u]�U���s邐$�k8�5�.��k Vc�(�P�j��g�O��⏶U
���tt�a�5B�qØ�B�׵Z��Ƭ��V�QDV#�T�ITʤL�Z�4��Vt�|^���j���X�B��ڸXBd,��I�"�q������|~,�h����Jz{֭/e�x⅄|�,J���k�$zk�H|����M>�_-�BTB��Y��y��.��U"i�L�\p\56�\"�R*���x�-4�$*{�ڢz���_�Y\T<��\/�}��"��_
G�O�괾4�$&p '����z/�;�G�d�H"��#����p�2�Q�|C����l��xSqt�j�k�㞛��m�{]�X�Gi����<򚫿�����o:i�
�&?W~�Ĩ���&v��_n�Y�����A[)Ic,�Y
�	O�ޫ]+��l���w��tߜx�,��I"S�V���*��TE�TB�>�d��t5(����5K#���$�'�P��7��Y�\����<�N`!��HΖ+�o��pKx�8��+��m4ȿmb��x.C�.v��-��M����0"0��A�s�rHB�{}{�A�$q���_gc@�l�����a�֘Į�1P�f���޺�]gI�\��t��������ӱTDh�o�#�m��X�c��'4��Y���"��Pr�o2m��7�4�a'5�=[4��{��*�k��;�u��^��#���剆�Oq�H����
y\���5γ�H����4�9z�}�8&-;�Qma�v�U���g��p���>#��"�?F�g������Ω��h����<��<Cq�H_+j�)�#���q�z�%$X��.y?z�+8,"�}u4Ⱥ}$¢#�޳�zSh�?=��^/�Gf�] �����LjG�N�g⪫e�e�蕊J �	���e��w验:t���3G�Q�kGw���\������u�cA
�������BVh�S_KV�L��Պ��U�!�}������F�3˥����Π�FIpe���t"N�Z3W5�v�V�sϨ�ѣ�*1�-,�
�L��L�uq��Z��k�?`ĨK�\���\��Mb4�5�±M�}\���K˞��a�QQ�yh�y�B4-y{�������e!�Y����ϳ���;��ؐC�#�.���C�%1����gUL8Q�_1PB<��~��_4����߶(�$�pJ�wN��uZ�7�����%G�ɻɌ���f���8$KN��G�,��ʵ���a��/�_�>��Z���Ł%"ڿ"E��9��ɑ�g��ϭiu��F���w��q�h�8�t�+iib�߽Ő;u���{<|��O�
k��L?O�6R�E��^"ϯ~��Z+F�#��k	���pWn+�1`����ȓfj�LE6?"�&�I���,�*�e*��ϻ�[D3��P�O�¢O��Z�5z�J������i�XҮ��s!�GD�����m/r���{�Y�������F��ْOqR8�<Y�{8+���[֌�tv��)p�LgJ	�F������u����:tN*U��Ef�$/����.��!��l�#�KV�g�SS49D�T�R��p����c�8�V/c��c�۫�:�>��x�}�.�2����s��x.׻鴼�Kmr�u
�[B��᜞m��r��%	XĤ�.�__���aMQB\K��$Q��o7چ��<��?:n!#,p�p8�9��n�nxƶ���`s�]��򚰎G�[;kX�tl�|J��wߠ��E��iP��}�M���{<z�H]ϹIx�}��Pܹ���)(��]���Q���~�?�K}/��#���F�����e�o{X��FkVH���`��8�q>��Hy�(Í�ZXiRT��N���iW]}�t�]]ko~�?&m������m-W�Z\���櫍Oez������҅s���.���5��u�H���-a"�{{W" aB]�O=N��F������O��1O��"T�6�χj��� ��yQ�X������U�謎�K�U��-/���/�����8�݋g�V�+����|*�mե:�����Z]:��Y��/��p��*V���� �G���Z��I�N�d��SKhK���m�k�E��]���I���I���WEy9\	X+�R�"�&�����:��0�u�U�w:����l�!��G�-�5�
�:��=�Z�9̯j��kN���� �ʱI�h��O)U��7SU����±.�+㜯����_ς���r�JE���ݽ�������/��Qp�g�zaX�A$)=M1{'ڭ)s��4���͈F	6%$�ʰ�'���*(SƦ\-[�X�����A�'Ͻ��n���l�r|���_AWL+<�Aۗ\^G/�Ww�ޥu��L�7�1���s�T���rIǱ̒Z;%���;����N#O@�[FV�='��p� 48����8�����O[��OW/T�F��[cgT�h�z�k���G\go>��ܻ��D���L	F�:�:�[e��(��]ˍ��ٞ�=��G���m��da�Ş��8��dSx秫=K���s�9ۇqV�u�<ۛ��Ó^A䳃��蝺���O����}��_�k�.��+c�Wn6����R�;lj�Ǉ;��s-ʯq�����3\�n�����-����!Q).�b��mH�~??��i�Mx���,�$�����-�dA�8�Cܐ�[�!�
�e��`�X�Z��t���8����9�ի����#b%Ȼ�N��V.�V��f�D�1��2MU,LF���!�r�J@��{��XX�C.������Zë�x�|_���Hk�w����f8t�z�ܷ*��%D1O7�W�F�ΘYDa�a%�H���Ҷr�v�0ś9���^�����;
�]no�^J��M9c�uJ��ыk�R�i3T$o��њ�uX�$-�yKD.��������OВ/��[�#���|*��''������b�w)r�4:Nȡ{�s�׻��||+�Ec@�z����f�d}�:$���ֱ�>>���l?f���p��S���z%�dIj)!?{�r�1/��K��/��P���{{�+~���I��T@{�'L����{_�A|��ڵ�4^<-�څ�g>�d|/Mu���ODʊ�YKn�^��\jC�\�Y{�U���zD�ՋΞ�H�b�[mp�*~��=�MqZ�H��²<���q�o�=Wn�
H����J�A����zrH�˛,�B�v\_�>ݛ߷=8ү,8Js4�&�>�w;I�͓k��	x��xt��ϑ�/�}�o��7k��!j2RpF��!��!���B��6\p��ջ5-�N^��y<�ub]4W�S+#��Ao���_��U���8�E��T�4F�F��0���YS���t{yS��o��m.,4]�e� Z-$����4@��Ͻ���4�M1�(�L���81x�-�̮K �8\��ݫ��G���ɺ���Udզ?�햾�J-�6�M�-�j����z��Ɔ�h������B�K'su]�
ޑ{��"XuT�GY4�f��w�I��Lp^֥��綮�9q4��ȴ3�i�N�K-�(TY�n8w���ig��x+m*�|+ɯ�|$k�w}+H�Om:�s��5-�����i�C(��L�^8U~��p�L�L��Ổ6��QϽ�Ց�|�H����5y�t�q�~U��H������F���So��xH��1�ޫR�a.ϲ��Ʊ� G8ƾ��?��R:�Q��J�5W�;yw���?��}>�<z�3�]K�y�]<�{L��W�a�SL]n
�ǯ}j�{y1�X����Q�E�y���൹��*:,�䃒e��{eEn}ʸ�p\"�����������0�l
��$p���l�mY
m�(@��s���YHL�!e8T)��6���o;�o�9W$f?�p��M5�p�w:�'�{�i{�s�֕�i��K��oV,�������҄����?
�N����.�I�d@Klɐ$��8��OF)���3v:�5�:歞ʺ�h�qkn�����ߟ������t�P�i�Ԋ�&�T�ޫ��X�=����,�,L@_���0�+}U,#u��&3��E�)�?�ŉr��|��C��<F�D �e��RHB�u���TI�||W�S�T@)(_[G��h����n8HIn��8.V*�+]0���Ogk�p���|_�Oy��ڙ\�}̙�E��*��{�W��0�Gl��)���B=�s�8i񜹢:I��I%�xn�������\#ď���]�*��}���?�,��v�J�a��JKu'�<�x<j�Xeu���w�ޫ��h�]i���B�w�Y�d��SyYw2���'��ͯ!�����f�R��Y�7[d�K;���?*�Ը�F�|-v�������]�n�9����wXVJA�y��E��!�b��./_�_8쵆	X�& N{ܫ�~�VP��c��e�"�2D�խ��+�O�p9��!hdK�r�z���+�q&%���_j_5Z��=��[qr����x�5��)��V��vR��𨅴�;��}X��vo�E�k��C!���=�ܪ����" �_�?Ɔ��U��$�͉w1Q
t\y��f&[r"T���(�Z�Y�QE��+-�V�F=�TU����	�~�'�8��?.ǯ>����8଄�4H0K���q�M[�,Vw\���a��a���4cI��cs쥤,]�I��u9�\�`�hND t[�f4�!y�3BP�G-rm��]k�Tq��Q�0L4Ɉ�`Q��mɿ�?~6X=�,��N5B�d���ʵ���i�ἦ&B�J"���"��ܢ�Z\R��C�;i� ��S����rtX�^�X���������EE`��D+��J�ee ��-mP��K�'��i���M*u3U���H���g��o���2{���8�,���E�O"�}��1u����"����i@i����),�&��ެ�>�Tqe�FcI�e��@��f��o�*\pR��6�����D�Lk�z�ŝ�S?"]6:l����"/9٬_����h9���k�#��31B`/m{svȱ�q�~��Wh��B�"_q��%4���S�)>K�)�wޭ\�e_J�HĬL�����=�����"�Y�N#���}���Q�ad�j]y�5�VB�ݾ�������s6~�>�ZW��)=�
"T���$SN*o=����� >0h\m�"�϶��{;V��J��i3
���X2}�����ez�_�/r�y�ni���|f텽z6�ۃ8�E,�f��M������V9���k4����8�\sĸ���/ߊ�FK�*Z�[�L-� ��d���9�BIo?s�\h�_k��N���M�:o��e}ğr9Q~E����,�)��.�� Qw�8�w
{)HS���
Oy�<zɽW*\���(�$
�Ecd)�~�Z�pbf~�VF	�R����m�3�o���)H�-q�B��6a:�2.z�^l���+�\�<Q�������ے��0����������V)��a=m{�u�k��t�	���Qx�W��V����B�%Q
�{)_��V%�������^%�$O�ZB�IP�__7��[�:&J��,赵V�;����u$�t����YV�]s��=h���(�
������0X��q���/�?n�|�����a'�I�ߛm�\��i_p��1l�sZUs�z�t_I����%�z��\�w��ZJի����V�ľ#�3�'�^��w�P�������to�q�rWF��iks�fz�0k�ӆ-�J���5{J̮��x����H%�o'6���'Ⱦ��E$te�.�ye��ӢTs�a"���BW��U��i��^�e%C�mI
c�֧
����T�5Uk���b3ݥ���y����O��S��^D.}y��\Doxa���WmKrN5B����q��Zg[VF���%�&�﹫��p��뢉)�ڽ̜g���,F>��羬]���@s��D�>���T�0�r_��/�}_���蚮��	����8��.ּ���-�`�[�~��	j�υs�ⴾ7�-ݯ*��CW���7ݬJΚ-[�X��G�j��.��Ҋm�%_��=<��S��������e���J��}QNF���yW�)[}XcPrjVVS�h^\K7y�LD�{Z�^M�W��x���mI&���Sm�T#�}��x�"�.}X!�m�LcC������;�/V`�l�:{N�r=mu�F����l󃮍�8�'���l����-
v�m&���曇v^�-�s�S�������knG�l=�N۲�󶭮^u��ZS<J���JO\\�u�r��G�B��s��:�p= �N���1��m
�.}�z0�Խv�7T��+mk\U]r�M�.8�cN����iyCQ�����`��9��뎸�Ǚǁ���ц���������׺�p�-=ֺ�V
e��y��W�[�T*�cp����z���Ia�n���5ߪ�]� �d7z<�պG�R*���)k�wx^�WN,TG9�ـ.J���J�:bt��MM,�dx�-6i�,�(i.0���@㙲�AB�S�;R����TE�׾�V%���Q@s�U\�݅:$�����	F�H�Ĩ����=~�#m��O>��L�C�x[m��RA�蛎dĹ��:Cs5W�Zg
,Mf��N}��[8)�,���+�r����>�wKI�.DZ������q]��p�K�}���qs�w�O�2�Vx�([.��r�_;1��,^��i��22��PH�͸������!�ϰ0�{⮨o�@�ڀ4����h~:KO͠iQ�ؑF��#K��ע����?T,7��O�a"G��V�S�^_"�@gHs��w��]:��#�D'o����@�29}��H�k ��������㑴�>�0��l�(RE�z����X/�Ҏ�k��$
�=���oE��M�5׶W�A��TtU���$�<%\��ZO��
�LRt�v+#=�j�T�m���l��X�ۆ*����ɒ>^�c������|[+�ɏ%�I\��a^62ml�d�u$�6���i`uy�ۘמ�w���#������Je���6a��\-!24z��([�X9��!p����%�|+=n�ef�+�;4w�{��ί6%����X��R���;8�^���a	M;"B�e��HtS�T���0KH�J!e�˳�X����b]7�K�ԇo��8���C���w��Y[5�ˈ������{�t��[ˠ�taF��~�b0#UZR��{���Ϳ�#�ك��^;S�ߢ?s>,�H�8����+K�_%QAƨ�GŘ��7�����Y+3�V���G
r_����񆽵��n�e��|9n	�($R��|��a��)�������f�j�L�)���"E�{m^�l����,R�*�\�d}�w��u$D��0�H3{+����@�����I�s�tCu:YP�$
��z��x�!r�;�Idv�a\�Ϛ���2��%��\m����Ϊ���2�����ˇN_���ʆq«w?ެ�DtO�,��=��� ��_��U���e)(Zo��h�2��}W�Ҏ"��X"�m=寮����︭x��D���P��k����7%5HS5J��ϤX��"��ݥ%�t'����Z�8CN	y܄�����}��:��r��.�'���8<� 8�u��]A��+9�rزJ0�*}�=Ū�㉸Yn��)�%������o��w��
"�&�lX䢕k͗�kYx�غ�.:�Wh�^�qk��jG1� _������ۜ����R�j��?s*�E�G<՜�,B�>��dh�m|D���[��T�(\�dX�zj�/z��"����v��ϗZ'Z�(	H",o��o/�Jp�^+��&9>EO���0���֑��@�Niө*������E�&�=ɒ�ǌg)K��}��`x���WP�(�R�zG)�>N� ƛ}_��z���aYb�\�120���{+0�3]E�.�NH>xH�_��+j����Wѳ�|�,�߱��x0X+,��;���j�9�����Yg� 	�DJ��k�,�y����!}�S���ݘTXg������Ր�� pq��Yߧ�����.t]�S���4�v�j��],gV�9�Q��q��Ϟ�X���a�1iy��ź��Dl�����e
`-�뮦�˩��^=S�;AD%�9�����S��c�V����[ˏ�Gq����:��YvOkU��vi�p�x�rA��B;[s/Y[u�%�;�֢�u�ů_I��k�n�1�yߩ��H��� ��}G��8&;�0^�t7�kT؅m�IZ����P�(dw�^!�=47fb��G!����̕�d���3P�klܲ�Rӵ1d�ѺL-�,�.�Y�j�,s�Z�_`]-iY@(</#t��^��ى�+�!!�^!6�����r�f��PuY�:���X[�x��#Io��H�̯{}��}.�U���3r���7� �,ɝå'�$�.�2��k����i�t�G^(���;���w��cw�Sc}΄�������:���㛲>�\��O*�Tx�%�eFT����ܴQ/کmΧ�sB"�HCj�ڹP���b�T}�*f��U훋��s:{W�[E���ffLd����z����I��*��7\�)�t���	���p�f��zI�a�.��G%'������74�
��A����K��� �;�m5��]�8���,�-t�o���r���ۘ��G�Z����7!(�b�*$���6��b���W�c�+.��Agb[.���2�,�_ϱn��E T�+V<eE�f`�9Of�Q}��7�C<��v���}嬰���͞�Y��6Uѻ��;��E_�%��"���f���)$�%�e�]}��i�f8C��Q@�YuL��,�~���Ӏ���$sJ֐��i�TAI�oW�گ�聐��T�}��������!L�	<h}��^�+�Ĥv�-���������+f��]�K}�����ޒ_]���r�O�{��c�K��JJˆ+:�l�d��4�@�U*sUh���~$B|��D���7�9��'��afE,K��E�,\;��{����}{�#=2a
�ґg�e���}�+�"��o���"��pФ�5�ޫ@�5�h�<�VA���mJ�$Y����*~c�̡m�((R.s��ڲQ{A��s�`m���ȼ܎ƞ�5� �n�A�<�h!������>	�!8��(����+s����]�*(�p�Ɗ���|9�j���a�J &�������y��噔��2��~�p�w]��t���t&cr|)ݺb�~�~�� �
�$�M��{�l��~BxN�2�h���WfVJ��`/�)W~ܱ`q�C������t=���H�6�8�,��3U��L���x�$J�dx�"P�e��b�����p�9=E���XqЕ�e�o��h�ZI�.��;]pUT>~�o���?�K�Ì��3�cr
�^?#�QB	�������v�iB��;��D�{���,��D'�엄��ݯP��i�?w�W;rl9BV@�h�!�EN��@[K�~D�- "�AϽw�	z�uZ�-_SK����j�&}��6�ʪ�JX%I.�{R"a�~�L��;7E8s��Cǈ�������D��H,�$Y	� &v�}_Oܯ�"G�$/�B�`[ �{���@-"x�T����iϕΦ�~�ޤ�~W��m�%�ݚ̾���5t� ɱ� v^k��N|5=�f�i�ÝҚ�e.��S�W���:��e`�!^�l5:y~�Y���I���L�߅�ݥ�K�&ub��KA�P�������D�v�V,>�'��fM���<�VQ~i��U�F�Ў��5��~�E���^��6����y}G���G
��l�ހ{�o�"9���f����X���_z\���i�O�Wg�N!�3G�W-݋?g�P��~P�H�a�ܜܳ=v�r���*�/1^*��nk�Y|Mu�]��T����L���m2(���6aH�i�W������G-���Kf�/e?�ڵ�=7ڵƘB�p��S��~���>�����9��aߛDQ,�=��x᾿cF6wr�}4@S��s�����B�� �g�����f�!�/�e�9Jf�o��$kS�Uϸ_�{⦻�g~kb
m�+m2/m�}���p�k�q���*�#���I���V�EG��EܩA/~x*4G�٢���cyQ�][�N
�=]�iG�#�����ڱ�}IԔ�9&�sU���,jH�Uo���}���4@��=��F��@+��J=����_
�U���/���ZE�{U��e�	uk�=���v1�s�����U���Y%��),��Hh��7}�W�MȄb&�Ga�'I:/�  &�g��k/�q1��}����"�(B$�9mQyr���Z����+�ε"
#�TB�KZu{�x}ƴb�,{d���.���p}�@�O=�M�2�f���O�i�r+�>�s�T*�`��i�'����E2 �[K��w���}���i�����6�����L8{�w�����N��� *#e��!M�
cr&��;d_����"�q���.(ۺr8�_��qj��9֓9�4%d1H���yy��0�&
ۀަo�ϕЊ�A����t\��3���K�@�4����+^�R��)u�0�L�o�Y�&o��8����}Ｆ����%����/.ݔ �n�d
�꫏X�|�nXd赻z���ms��}�������}j[���Q��6���ی��3�6z�\���
Ӛ���h��v��q�7nx��5[6:�>ݺ�n<�Ok9����u���^wH>؋�k�s��BQA��v :��f�n��mJŞB��˱��!���l��A�^I�"����=�oP�[dgr'ex@y�gD���]N�c^ٰ��s������9���݋u۩�s���O'N�C]�?����v�N�hRSO���XD�W�v��3�tX�i|�*.�1��5Ͻ7�8��
�DH�-1W���B�٣ϻ��s�j�SrX��b�s]�~ⵖ���XĤ\��r`�Ro�m���
E$R5X��>8T%!-QP�pe}��	pU꽒�_��9ߞ��i��6ؖ�l��|��{il)��"�TH���r�}�qb���t���2��ϳl#x�;���s�ʊ</��v�#�2�|?b��& ��GM��� �u,n��5�[�Q)B�����:�&t^��,�q�fb`���J�)��	�&�N��*�z��0]y:*s��b�l�"�\�m�� �dX	�'=�U��o�1J9ͽ�Åq�s��P�	~�~2��Ӊ��pZ�y�\e�!]���\Cʒc��k�_��M_;ެ���>$T|+>>��+����V,,X�aYBɬ�6�
N
>�{j��}�![K��^e�g��^�fzn����^g���A$~G.r��Y��kk�<��!Kik�[4�o`)!-�J�(��fmw�Q�CŚ$�!���c�R���?W"��ܬ^"w�
��q��
�>���ڷP@�D��I7<w��p���]k�J)	ݹ"�R�T�};���_�Q�_���dV8~���ͣ����Wgnumr;�9�'F�h4��H0l9�'%1���UUW���0TE+i����2���̫��Ԑ��<���֪XY���b�8SO�3e`�AV�旦}�@mz���Z�����V��јA��OD���tgy�F�v�a��Q@�Ŋw4��A�QD�**���R�|䱊��>k �*��=�j������w�S�p#��~j��k]�tğ�9O"��݆I��H�]^Z��)���_�kveO�^�w�3v�gE����m-��~�b뫷c5J�����]_���ʰ#�pS?s�����Y��lܦ�'m1YS�z�`��"�=jB4k�s����R��|G�Xog�Ӵ|�Y�}-��.�T���b[z��C�*f��!p��U�|�<�8x�'��΁/�.ݠT�Zb��mZ4TH��sՐ��+A
�؊�n}/���_�{�?���K�/;۫�2\���?]*!Q E{Ֆ	�q�#����$���s�_k�s�UH)*��\_�*<E�9$DqU5��=�fҾ���:w7�e��T���R�'�1DV}�Uƀ�p㮥*�SdB��T��>$�D+A��A}3�n���7֗o�u\`!�)8�An$��@/M}�+d�QLt��5Y-֜ےm�Dr��T�[�~�z�!2i�W~�ձh�=7�����)K�7�Q�f���_AS�9�m��.n�$9�V�5��m;je�"�R��=V��L��j91@ሗWϹ<��,��}�d����m�)# �l:d ��Q������Qځٴ+�ק���Q�U��qR�)�hEL�U{���E�n�G���^)lT٭N0�8��X)n�����z�-/�D��VJh��1�f���ɧ�˹�$�igD�K
(V/��ɴv���T��(N$�d�h]�4��#�"�r�~ró���}](X��!����k�p}}�sky����,�oe&Xψj��ebA����+}Bc��o�U��gz�&�FSH�D'�{-pCzB�}���6��.���
�$1�mg�	���)�L	���U�ΚxZ#��rF
Jy^�Vt\ 'O��:���m�(Es}��:��ȉl��Mw��n��_�ɞ!{�r�I咏��4dwȱ;�I˵Z��<�������_A)rZ�_|!��Z/{K�o�������fѭ���g<��8����ה��p��� �gݾ��˿��h_#�k V-8QeK������1l�	M�a���A�^�W�/�U�Vh��C&�vn0m��$�(�4�e��'�z����R|'M�Qcu0��{p�󞴚��x٢��,�g֫���U��b�8��+�����`������y�P��T���jqj#F?L�{t��H�D�	���{���]Y
�\����s��A9������N�d"��R�a��,<|Eߟr�p%�8E
��JV�RAG)���=6�.�p]͘b)��M���]-�ߟn~g�{d&��$c.}6�a�]Z��j�ڊѧ��im�����:���Uͺ�j���]�����u��;m�)(�T�}���H$`�|q�7�\h�.|�u�o&�����H �T�ZDJ������\�ޭӃ�w�_����:�s������S�L�}-��%P���!ƙ�\�z�����hc���Y�(\:9��
EX�H-ř����V�_����.%lY�϶aag��N�{6�`�ĊL|5c@������س ^�m\�i;��#C8O���qj� p�F2�������
'+� �'Ze� k�m��*T��5V���2�
@��q�.bM��=_M��q�u�[����tX�:�����[@J���M
�X�����mu�����1_㢑٘Gh"	�����C1B)�I$v��k֫� �����_ֹF�� %���0��~���6��+�8��;�T���,3��,L]:p�8o��Ԕ+[���uZ\=W�����;�+��n�)O;괋zp,&���C�C���߭��L={�{���U��s'EǲPYBܵ��C�x졼�>���<��Ѻ�-]��ћ��cY�Om�_�?����Y��P��,#���6L�E���FL��cpW�A�G�!P���DX��3��U����b�Kc�mW��'��Ω6�W�.q��,�D)�&/>��� s�Kh��w��M���q��j��->�����3��4yV	��w�Y6���'m�V	�bKM1O*[�D�Q��z&e�9]��\��x7e�ð�ۢ��/y>����$E>	M5��_�ޫXF���51���O��I��,��/k��K:��v��3&o��{� ����{�_�ZrW7����]�i�$�7�*ڒ$��{�j�bÜj@T�hR&1)!Wы�*j�NITʙ���Ä}�J�/��fP!b�¾�s��$�E�|�x�ׄ�Rġ��
,��
�*��o���r�a(]�J�� �]���@m��4�\��$�V���b��}X��+Nu䴜e��T�z�IĈ�E�[���GAj���qu7��+�`%%�N�����t�;����A�܆�D�W6_��Wx�@P���q�9���J�IO}�ip��an�d2HS?}�Vak��!�`��LNZe;��s-i	�,��Z#�i܌R�D�����^��ۿσ��I������P���ϥ�+!{.b����Þ�b^���3��N�
�E-~�.ů�sq՟�v�~��*7���,��GW�?R�����9�kQ��;k��"@�/���?rfB�s┒A�3Q'�!l�	"߈��ŝ|�s՜FG\v��З��j�B�C9މ��h���/����|��Yb��s>�Z؁h��{��,g�̊��+&ZT&&QDQ��ƍ|BTK�)P [`{�*���D��}d���g���K��-oh��அ��VĠ�U�j}R�rV�z
�xܫGQX3�Q~�2dvN�%��)P���ܸ�2-~�v�m���F��+>��7$�^�4�d�+��g9�ݶ�^l�.���uca��)E��3Av��ƭ��閺�ʆɸ��8�\�;\��==bB;�^6^c"��P�m�n#��7=�0�m�1�t)��nR�uF�c�zy����ܻ��:u<�\��ny+8��j�ŋb�M�Վƛ��ևf���jW����v������D$�]�U T���s�s��a:tuʖ�^N6��&���P�E!��u��t	�W=8���p�����v��R���)�$~�^W�?2r0OZ�]��b9�*ۡ>���"Mbr TC_s���X�Y����V�K�4�?q|��>8��l ����^ͪR
\��O�"@=�����QD\T���O!wZ�,` Q�$�����ⵀ.
���5^�s�&���=۫��c*�$�A����0W���x�Sv&!�j��
f�괃Fh!3�pT;rM�C#��߽8��>k��;<)�y�7&y�%��*�G��{���1���%��kA/ҷ&�]-��`h��!5�����W�͗$�6�YB���J3�Uذ���1�g;�㚩�38���#⽜��Y��}�mߦ>7^ 
��������k�W+�)$����W}��IIQ�DN
d8B��(_(A��7��d]�?N�IKӫ'��W��^�����e�ɋ��	��a���,#�|�9�"!��!���,G�����e���s�Ԙ���j��q|i�'�8��(�x)(O�
7'�����J��İ�&h�r�4P��>��kx�p"�2_F�}���Oi��(�����0��VY�`�����	�8 "]O}L�e��U�:�@� �<��B�����ݹ�lJ���Y�{�i���V}s��~�r�H�u4�������� ��sqغ$n]�=U��I�t'Z֜b�rݦ��j���� ���B�1�v^��ŉq������4����?M����V�.q���/KRe�&���RH���_Y�h�p����^�/���ҹ�h��D�O3���p� �e�%r�7�
U�U�c��� �'ST�D���.l��Ak�4��t��{�V����*6��BZ/�o��*Tl����t�7"/����>k�_Wfr�ð]m�ژ���rZ����9u��k渤�7a��w�~k������J�~�5Sm�\u�F�eT�xa��ebY/x�P�u2���䰂�d�?}���k��|��yp���Ϋ��#�$�E�������+:�\��1��*8�p�	���,��Ј�6U��Yf	�I0b���H��L���x��+�k��|��-#��Fz���-����9@F�R�G������r+��!Q,�j�R����,_"4��==ڱ,,^(�0+o��̽M:�U7SU���i�T�<Fo�?oE��U�i��w[#��>�U�p^"���7\�m<j�0
�{)\'�I�m>�~���i��1���Ydec�����[�F�:��ٝ���~��C��4�/�A�a":aD*�g�C���e5"M��8��>���Ж�J"��=\V��.e�~���	CGw���a��<�C����]���${�VE���N%󞫌��ǎ�mav�#��H
�g*�,�pL�X�Cq��PE�"����4>��~��ۮ�^�y^�9Ѻ�]v��ڞ.8�8��\L95v��ͻn���
��5�Y��/��	�	j�%J)�q��Z�Z/���|ץ���zX 4a�o�`��Ջ�Y��i)�X�_ٱW��^��㞒�o6�00'f������/K�\���b��^��Zh�:%4�q�N?)�I2�UN@����\'Z�j��.�	#}�#�R��N=���.�;�5q�׼�kf_>ڸ[<S����-\�ｔ�=�c!��߽Q�n8HkL轼�U�V��ߝ�*�ڴ��/���p�DX�GwL�R0iӥU5YbӀF�1+�d@�[g�X�	���,���"˴=e~��h�Y�ĥ��wͩ�.d�'~��ie�L�v���3�a@U�y�h��v�B��^�a��$��O/]����mu���:��;�=�e{���]xح����t�<�(�I�& ��=l,��ڼ<C��f< v/��"y}_�G[hy�[q$��9/�fbhY�NKB��óܾ���|-��uc���К
���%X��uZ_���>�G��:~���*�qCy܄��\Ճ%��rU�е���U�#8��U]G��9C{v~���?�gg]�1iQ�)!3�p ���>��U��^�v@F�`B~�����Q��_��[{*�������N�RI�q#ɿ�ۭ]8s�I
 0�$��؊�*Ev����VH�Zh��p�m��F%��<�3��A���HH-����0(��\n�5���=�7	{vV�<�(��{ub�j�C�sK�.��0�Dۓ�=�����y�fw*�Qb�0Y��4��L������Fs���*���(JN������[#��Z�:��Ь��q���ƨ��6G���%6`�M����$h���
�R�H���x?R����49���F��.J(J�,��]��;���0��w�mn����*�Z�M���nDT+h:Yt86l�$q�"O{��8.�V�H���N�W��U���ㅷ�N��[��,�డu������th,�R+m�4��;��4�Zw�q�bO���2�4&I�1�M�Ċq�$B�~�B��
J��r�w}�{��|ܐ*�se���?���ԥ��L��r�"8)$O|�e�f�0@�h�O� 
��RK��ӂeu�[�$g��o<��f�������>˞�+��sɦ�-�G��U��~N*���d+��\>�i��q�&��^{ݫK+��֑��TX�w�w���>ʰ��(fc��U��٤�Xk�	��Ky)�v!���T���3G�	���o�3g-e��2���հ_����=s��t!���ƨ%���v��Zh[��x>z�B�L�&Sh�������8�YBAB%2r�Nz��ĺpg;�Ptz��~��?��y_-+t"3��WJO��2�pR"�b}��l�4KKc�MH�J��s]�
}~�,�:>8����\,�w(
�{�����no���&��m�M��Pby�%0�t�*C���29苳�D\��sطTI�t5������M���8���+��҆�H��1�'�[R-t���+�F{� �r�	p�u=�LS�.��ۧ�G��[�+���/�2���l(���H�PJ��J��0�G��@�B��,��j}���8��
Љc�ۼm����9s�E\��b���u�����g��g�_����<KlQ��I�!��=��F8�Q{Ӧ�\"}��Z��|D�*�G�)U<%�u�V-mj$I����v��9�m+�-��4��#�!r�J�Q��o���u�ؐ�k44b��4VO$��������_W�{e}�C�Ș�m"({k��K�;�d�B�$�t���W�߽���4���DY�����gX�+�����/���-���./'�A!��8ː�J�8+�c�/֐,U럫����;x�/����=��W�@�:Ԛ&B6ڳ%�&��>{�9����
�%	t�x�Ӿŋ%�s:Cְ�̜"�eUgWz�Y_}����_���
8
Z]'�1"��.�U���{�p��T�NTҒB�j�k�O[@oZTaٝ���ZL��2M!� �O���o��w=���td��[e�")�is�z��M���a�h�V/�)\��f�h"��xs�k���ywx�u�~j_T��U��Kv��z쌼wz��gi��z��l5C@��7�Eu�!�vYk��:��yf��⍑'�0<����&��Z�����VK4Ψ�&T˴�7$W�/H`V�h]������^}���]�����b�K&_NF,�%`�YkN��OOqT ���=�v]f�bŹLE|�k�;�΀I/{����u<��W/�e��C:�v���V�����]��5$��[|�n��ks�B�D���+�Үc�/�XF�GeL����K����^��f;�{�
2VT�@�s�<���GAыY]�����:����NG7.u^�]檆t�ݝ��ю��ò"~ö����<1=o�{���;�%��n�����:mygK#��������T��bA��޲��|��`�J���+�����9s[2�U�n^�F_l:��J3%f�Hm��+v"�y�މIq}FeJ:�r4a��5(�F��J #ڎ��$�[�h!���ջ�z)Q���wZ�&Ů]Q6VH^f��axW���wd�{RA�� ��XMG���F��++�P�'�����'���o�m=��7εc���R���[F]�]��uY�y�`��feuu:�Q���^������9�`���'��O2*��%uZ6���]]�5�,����/?���:�`��e�EBW��9��XN��W��$�R�!���u����~�=�?���W�~�
�E�,��R�J���5*�m!��J�m��6�G��S���;]!���<Y�On��&�G�v��m�.vhnu��<[]�������H�nȇ��K�r[��ƚ��/�.����v&�ݵ��a��[a��������ek���z����sn�7V�.�N-�sS�q�q=��v�ӝ�\��a|�:�۵ݬ�Q�8�qg��s�x����vN;j뭦��m�[�p�Z�W��f�&���L����������8Yۘۅ7�����{Z/3�v�ݻ����-����X�ņ�y��\:ݤ���Ҹm�4^9�np����vs˵tf�8޷o�3t��q���#���>�R��� �tmŬ4�v;y{EӴT��ѵ,��P�]��yOnz�Ͱ�`�s���讂��r�:�s]��,�e�v��N�	آ�u6v����:=�����'tkq;.x��ͭ�㳃��!.��OSp,t�(e�<���6�oY<$��A ��Ƿ�B:�K§�v-�HB�(ݴ�]��=�p�K�����n�؇���h���O<v����Of��%ܳ��vs��Akr�pͨVr��\����*1��Plv2�����5z�v-n��:5�r�r��ۀ�̂S����L{<d���;Z�8��:�8;�	���W\!Ev����n��D�������Ô�Î�)�8�ڇ'>r]i�7�O&���']B*�`thڼ���c�2#�s��ֹ!|�des�1��Y�J����[Fg��/��v�]s�un����飂���,�C3�<���cZ�臭������u]q�n���O\�i�.ٽѮ4�mg�vݷ5�N���=۶�n���)���ˊ�����s���콺����\qt�D���.�Ŝݝ�X:�T�Z3bN�܏fc�.��q�74T����c�]�pm�`��<1�ƃy�nz�r�(׍�*��A����k�vNT�\ۖ�w����q�lv)��R�c�P Y�<&���j���u�{�� j����j�����)�`y�u�u�Ƹ#C]��yz;i�]���ė�p��#�rǷ9|����;N%;���v	OpF���,��q��-���t�F0֮��V�[�(�ۺ�!d���P�fq�q��k�����\V�)+�1����l��=��x���!�Jݖ�	�]�tUb7���g���V-!�6����8u�mvŻM�X{e�F�Tn��4�\�l,���mOd�k��;�3Ê�i��'��������v?K��ݜ{����jWV{�W��L���0�e�e%>�t�%�oc��Cs�g�E�b}�}���z��ν%���ذ�T��;�ɔ.���l�A#f��gZ4m)��DFpy�^bğ4���@�F,4������y�U�|����^�cɣ���u��c�����FW,�|_ݘ����Q��+7�f��gҡ8�/�m��AA�f[B�#�<ߗf�t����誅������i^��p�������tzCk�᷺�Γ�+��/0`؃ZClĕO�A��r䔭^�30�nw���|/V	���Jx�dR�����3��luΝR���B�i_ot��ʨz���q��:+��3���tN�Y�[GP�!�v�ɳͰ��O\.��������:�m[6W.8N�d� N���r�^�U9DG�o�E����!�y�?bIX5�n��
�W=x�{v��`w)�I��3")��
 �8[rc	o_J�m\B��J���7+�dǱ�u�aۇ�d�Tv�Z�.����QLwz�e�lhIZ�L�v���҈i�/p��"�W�
�<��e��Ԗ�������:���^`��U�z:�UQ玥��u����e���?�[n��Z#BOz�na5Β-YS��<�U�3��uko�m�H������x���	f�U4Gy�c�I�a���%��nD=�"�_�GsO���Z�Dn�^Ǵ��(��s;�6�H���$�y�c8ݓF�ڝs��*RB����:b�3ǻ�tϔP���!*����Ԋ�m��`-�<��^��O�����*M�bD+1r��Q�� �h{��۶�;skm����%F�˱�䍛Y�f}�����%T�8d��#J6su�(�2��<Y�����.
�k����F7O��S��c"��jow��YZ�v��]_�����{W���a�U�15{�=�,x&g뭣d��D[I��7$8
Ϟ�?J^wo�^e��{�ھW˲×|�&�M|�d��M�`}��W[)��0��T��g:xy��o�c�7%�S	|���1�����%�ɔ������ȇ���w�}2]c��JF���*�*�g/��)��S93*<�w��/��s�I0����� r�;���[3���7�kiH�2�y�Uȉ�
�z��]���.���Y��-w�H+t�1��F�p�Z$�Q�w:_�A���L�����W�h2�S�Ե.GnD�۶��������ه}r�Ί�mz�f���W�,yإw�����O�]�b��R�R���;������nt��b������5���n��W��n�uH��\���T�{F�v�M���C���7<�C��L�uڸ���ܛM9�6��!Wt�q��;��Ṳ���sm	�j����dY>��VRa�::�s��(<>�CH�2��xX�����.k#�^����L�vi�w���(C�)R7&X�΁�D�{'��_gM�ɷB��OwwP��ܨq���K4��w� Y���������҂�X���#��a�K%��l�ʞ�(7�����T���De+5�ȧ.MW��/M��il�'��������w{ ��2�5�p��8���#���2�Yxs%���_{6�;]<�{QveFo��U/l�g�B\[�X]W�n�z	�N��U=3g�����\Zk(%�Y�k�^�F�S-�cU��7W)۬�Wܮ����֞�D �F���йx��s���q�S՛$���E���W������%�Y D(~�E�����06�!�:�K��C�����|��f��#�"���*�o)�|w*��*�z@�a`��Ԭ[DK<\�}���)�.�ٞø:Gm��^�ە���y�0����9�>fQ,ofC�m`IH�w��n�1P���{�>��J���z��nI���h���&l�����t�tJ�+!���1�B�)��#�����
�_r"�.Z(�2�ܺN�/vͬ���h�M�_Գ+n��^����ɻ+�"b��FbG�"e2JB) �r�N�z��RX.�������+n�&�j�)�\�Cq.ͼop�ϭ�����CQ)�3�[������^�D#k�f'�rH7�ȧ���Y����;�Xj�iY܌>|%*�ŝ��=%Խ��t���-��_�UfN� ��l��ɛƅ����j�o��Ϛ-B�nC��߁M��V.��#��<,ҳ�;��!��n��ձ��Q7o���P²1�ӣ�3�z.�s�{�l�}��g�s�:󇂕y���⼿�ío]k��P�r��P&�ԡ�Ǚ��f��P��p�b${[�}[t/&E����  ���&yɷd�ϊݻ7U[��WnC9��lx��5�j�v��>�Y탷fC����F�oqt�{cO'I�uut��0L[���݃�ZCj�m/C٭m��n�v^1��o2�ԏ-<u��ўM�km�k��K�x��n��v֧��.��v1�L7=�z�n����ʙu�˸�c�Eχ������w�N��@v�l�Z^�Lvk���#J�9g <�������3V�f�6�wa�2nFˮ5r'ic��a2�f��znt��\�;J�-���A�4E��*Ox�s�5�n�c���E.˱��x�7=�C,��\�뉔�m0�@��̞�3UΫ��s��qT`gp���?t�^�L��ד>�ly�	=���@��V�oOzW�,{�-�K�/��~��&5����;$�V�~�JP���s�H j}�w�s�F����i^ .�_-Q�(�7�G�aߋ6�m7����=�f�*�]ҏ�C��U�v�Q﫻�N�AO�V:��nf��[���x��щ� ���nu�.��=��c�O�u�GQ!*�[��C�<}<�i�M���Z�]�oӲ��}V�cM��jeq�&D�y�F�e�VP�w�x֥�P��<�'�u���)���<�[V6u�����qyު��p�糺6�[�D�9:�����R��=08�a�ޔ,㉲Jc��m�7����!���{]�$nd��
w�K礶U����*�7$�$dX茻l�7�e�xQ��#�-�=��٭�'"�dp�{U)z�t�sZT�LS�f]'
��$X������PoQ�bF{�l���&��,��v�.��"1�ۭ��7�W
� R����Ħ ��Z�&��x�L-�vuPś��u�0U]�/��W�t�M)Z}�y�wk[-{������L:s�����4َ�p�?t�j�Cu�ٺ�y�����u�X���IW[�y�ql*O�}3ڋy�F�_�j��ljW!����fuݙ��Y�f DH \1>>��Wi���Ax��_�m���dݭݹR�qM���s� ���D��pfH�0Z��a/��o�;����J�R2�DFAA�q����r[��u���ݳ՛���x��Tnȸ�����rp�̖Ы	����8BeS��ۢ#�%���$];�m/_������V*v�Q�V3X�Uj�u�Eq`�E(�Ԓ���˂��\|�</O@Oj����9Y�XZ�U˰�E���{��5��a�g�GDz�<�O0��Z����mZ}8��8龧
�5i���Ӈ�̵�X��x�k'*#egAR��{�ngJ(q�5�/G]�]�Vd�󳤻2�ieK��Rzhe!j�
{�@Gu�D��3{�?vvÓ&9�-E�(�#�>I�E@d�w��;Vfv����gc���͑yYǋYBqW�t�B�}~�RJ=���xPzZ�}�����|p��J)�f��ŷ�� @�'b�G�݇�����"�˭��:Ժ쟶��!W�΅D�M�C��)]yRV+�!ԑ��k�ܷ���p{sѯ����}��̴c���^w\�F�{.�+m���xp\���vͣJ�-�����h���-s6n���b�œ��Je [�o��~\�B�<�J��1`��tA>�Qf�:�`�I5��`�����{��ݽ��O(��+7p=�1�r'o�:*WoO{5lW\s�Ό����x�G�z�Q3��0��l�
����s:Y�U@��N�k}�o�90�����(��RWl-0�}��`؇�I2T�E.I�ف�"2ܗ�d{ά���K�m-���y�o��.�Y�}�����m+�e*�]Ce�tP~��Bw�,�3/��/":��78q��m�-�c>�n$+f�{bG%�:56�n��ZiP������fk�J�T�W��@5� ]���p+�n}���}W|�<:6&5�Oi�1���W��~�5�ί�y���JH����ag1X�u�s�2�h�E��O�Ǧ�W����ʉs㱱�u�zsQ!�2�\5=v}v�]����]l��e����ú�����o�BY��}ǳ�E��U�T6�3��
�KʪE-���;��\����
����<[<q�
����2�� ����얭�P?;/�f��}��t�ʽ�^�4e�-2uʘr�t�h����1��4hƄ�ǂL��\}\���a�JE\�K$%�	��/��ə�	�`�"r���d�I8�RU(�����n��C�kW���fOKHY���I��.�UN:	5'��V��*:��	n�[�Y7��}]+����g��t{��E�>/���׀ݜP��-���:_n4g�pگ jT��x��M�~Eo�.��c��ӄ���HA��DY,���Y�z�s�y���Ϲ�=��4o�Ka��>6W����a��wKP���C[#��o�.���C��yu�f�M�s����DT�Jvl�ػ4�F�AWL=�ve��&؝�u�z�N�|�XI+�9I�m��kQ�Qݎ����8����q���D\b�k/b1^����"���ʾkw)6�e�u�>�E� �������ݜQ�u�p�D�gI.���/"XwF��E����]��X�f�V��3����m���*���9�W&��-�9�Nܚ��\>��lV0�3��V�'A�.K/a7�ݎlu���q�<՗ic��5�m��e1r����㙍Þ��"�ƛXE^�z�����;u	�Hs86ʼ���$z4f[R�K�ۉ���u���Ƌq��`��X<t�����pR���K���ۘ�ʑ	y�(��)��6v")�7��
#.�n/�s��B��W��������Al����=�wW*ɟb>���\�T�'1HH6$m�~�G${~�g��n����d�\]�L���[�f.��+��e��g�̙�-��S������X��[L��E��
��~םE
6V*�8�y�����n�w2(��S�dBq�HU*C��P��)�P{��l�O^��_������5�~|�*��-��(Z���2pk��>x�-�ʗ�D��e�λ�u5ݽ�y��x2�)}$	�~��^�̉�S�cX�T������q�N��rg���Q��n���j݃��Mssb���D�'͸�1! ���O�ɇ�:�wh��<�炃8Y�l�c��k(�/�����cz�}~g�7�x���	�%
r7#�9�`�>��������)AO+�vem��Vwf��î|�sZ���n�g��ofޮ-����BFc1z:�B�4���mt�������eksԙ�N@��!ȟ�3.�/�S'�w:�m⻪绊�e��s�g%�Yp/�f2؍�)f�Ae{���H��=n^��'˜ֲ\Z��η����}���-s@�.��G�9xA�:{�A�}ℍnA��H]�;��l�>Wb\!��^����y�6���XA���^̘y����b_D�z\*�`�o�xp����x<�o �-�T����0�7u���*���]ti&Yt��oxM��IUܟ{��+=q��Z�[$�7�'���� ���"��2�:\va��ܮ-ac7jg�vuph�m�:�D܌"B�F�u̽꫰c7�,��~~��>����0��I�Tږ��i��0N6����ݭ� �|�X������$S!8���36�
�U���J_H�L+<����c�E]��@�s/2����G7Q�ےгo�Ʃ��F����S��Y�=�y��q�������h����t��-�n���󯯞z�P�O,�`W�$�r�M.�72��w1���K�u��5W�+yq�E�G�����3i���V��3%�+�t��G�k����K"�p=�����dB!���Jw.��H��7-����<������P�NP�Hrh���W	�O���GgNHSI�����/4_��h-�`�sf9&���[
����v�9�aP��`7�	��bE��v�MqsUk/�Ռ��V�ŵ��{�M�&0hU��(,�;�=Ӊ��mo%�v�]s}�ۦ�/"+�W����hzD��/7BR��k�gq���F��:�֝�Ǭ�QXɀ�9sk�_vxm�Vﵗ0i'���%;�Yu�˧�q]��Oyq��Ɲ'������s�wI}*�tlm_U�ˡ�c�2V���ʵ��ʞט6�x%U���BWz7+����}g0�h�f���Gu��hE����'��jd���;^�o��y�u�^tƤ�7=cɉ��E�Fv�w^�eʃ�[�e��n��<��%�koml��,T�AC��8�.I4� �6�L~y:F-�����2c0.���z
{�x���GP�/]7[���|r�7[,$Վu+D������4��}��\Z��q>Ʒ�_w^���Q`پ�;�"�گO�fدq|uehk���M�V������V���x���fd���9֮�}����(z�`�^&:��*a��݇���G P��cp�EoL�u�I�OF�f�b�+�câ�ɫ{���u��TWO�:������9��a�+q��6hX��u�\�P�o]k����a�A��A�ӎbU��e��s�7H�P�V�4�v�Y�ȉw�0ẗ��>ޡ^+/9pT��Ǎ���{!�n�w��&��\p%{fl�R5�y����)T%e�yf�d��3m�����ƶ+�h�g]�8*��f�v���I����x!���ՅQI���3yn9��}��r\�v�q�?���<��*Ӆv��i�h2�IW����j�y�Oק�<�Mϙ�dx�"��eP8=���*wк�ra��?S��oE7n�4DY,�T�	_)a�No��ߐw�*�HNz`FNe����Q���l R�0��n{Sl�6Oީ<�R-X�������X�zX=rП&�~��;,�wH��?�VՍK1��4WR�{0s�8{�:�2���ʑ�8i�3geg,cfo�H����dH�P��/��֢;��箱:�ᵬ>�E"qN�`��}���ܒ���������>�/�t��c�\�����#!Nd[��~���
e�U�G}���T����6�Wf��.s�oyP�(�����0��ݞu�0���"��$~ݮQ���J*�9�1mM�vLX�n�Bxm�������B���S���,D�y������vy��_�b����F��뇮Є�;t��0vݏWoDsp�t�ӝ��w�7Z(��a ��r�ش���p	�Wc5^�uν�=2tJ�{��ߺW/uf�\��iN���E��W�]�.��v�6�~�ߏ&I�r B06���xmn��K~JV�#�u���ʔ�"��R�;����$+�u�aT��`j�u?�أ�����Ws'v��<Q6�0��S4/N���W��G�(�=4W__���|��췒Yf�y�j�̢\A��{ӽW"����d�������E�o�5ڰ�1�I{C1ap���	Ϻ�_���3!Q�n�6<�*��ϧm;�{q�+��M9j��&��"���JA�e�,Jp�S��u:�R���b7a���z5������r���e*��KvrD�A�(�^�>�ъ�\����Sl�P�&����z�f}öV��9q]��ث�zoGt�@U���Q���l��r��K�����S�ow���� Щ.�����S.ݧIٲ)t���7H��E�@�c�ҍ�u�5��q�K��[��tD�og��2Wr6b޷F���r���+��N�����Œ��Ű�#�����ۘ�����^�=�t��Ǟ]��olV�Nݡ��ڌ7��[v�1s��-����]�c=���jp���t�m�t+�q�9��f�8[���ryy7y٭�ax��[=1��{�cx��l��cl�Yi�\��\Ru�G`�l��Me��fj��P��y �(]3�H;�FnC.�V�]�7���=uY�[�Z�I�٫C�3����B��m%�K� �ȶ�فR�'����!g��{�q�c��%��:=�[�
$UpR��fz�7ep��^+�Ҙ8�Y��HA�ݒr��"����V�W�_�9����8�exz����vBo5?R;,�'e@⦄wQ��}!�&����Ay��ֵ6�{P��ܻ���o�퐄p��}��#F�*�|ҩ�l�Nw�o���V�7�@��"��Vd,B���2I���5�;9�°���z�זī3(j���4��2�~�Uk�9�F��n*�Y����@��Z�Vk�د�m���k��5��)۟�ȋ�2�:�n�!G�5qr�cl�=���Ӗ�������!(��=�*�8Wav�����q���u�*Q�|��=�������y�7�(��R*�ͻPI�Hd�I�f���.����N�Y��DQ]���G���2�塑�����Q8l�,�u��oV�+8Z$�[�oJ�H,x��Xsf��;v.f��	ҹ�ʻj���Ʌ��]��ONs�iʧݲ즱��^k/���R����f�X�b\����k���}�@~j@K���o�WA*�f�I��ڪ1�_wT�{`�,���ֹm��]K(S���/f�	5���<l����Mɳ0�����֖�"��E���ꏤl�v �z���^uK.�v��`.�W�(���C�'��>ʒ��v,wk���ka>D��H�x��!�T���#p��񉹛�|��w=uRy�1]��n�1�^�n�[�gݵ�ʠ�ڨ����JZ�1�Q�ɍ�q�.�5��o1�6�ڪ��^J1�F��$�y-�y�K��1b�j���B+�s�)���4Eop�&sι�y���4�"�o�v2�BR6kʮq7S��ʁ�RA�;��mV�T��.�DJ��A�y�y�]���n靹�e	x�d��݃�/�=�YKaPDxq��
.���9,��z��z勒0o��K��WK!XZu]�P���(S����5������j|�Xyy)�ca2�M$��3��^\մs2��I�x����&����<l�=�Ȑ���i)Ӟ�v��IOG�)C�\��C�#JF������yH�_j�L�Z:U��
�0�
 &�`�t��b��_�ĶϽ��P��҉R�5�k1<��z�4�_�8C�C���_8�eFw��U��k5�c뙮���ܫ�õ؄4
G��M��:�Ҵ.�tr��k��w�|F��I/U����e��wmt����Ogu�����g���b�=�����N'�۪���D����)&A/7�9���^�l�c���0��B��;�{Ɩ
;�c�*}[(PՒ-���xS��F4�H�����%��'첓
Lm��fm�Z9s����k��>���|3�"'zJ���~����>���X3;V��ݕ���r��&��T`�i�J��w�]$�[�.��փ��Ů�@�G�}�[�7���q���v�%���
�^��]gK�����""[�'�{n�'m^��������h�e��Mv\��ޭ�����y���3Ko"YCP� p����F��9�y�r�>4���(�u��c�I;�����M�ū�PV����ەٷڟQs:.d��&��*��Ls|����SB"�I���� ��A�W��>��=}�:ߋ��WN���W=�C������F�ۛ�Wu���o���?}c��pD١;]�����g��;�-m�:^8-�5֬���`��8��ٙ�e�1[(5�u{iZ�����¥�ˋ��.�t��C��޺��|*J]� �����mR��%E�U�8	!G��V���S"���T�����AUm�Θ�z���-YY*���w�\>fv��,ӡY˰I�Z)2H�$o4�m�y��y�^q��c.�񧍃G������Zڭ�6��Sޮ[��_q�����ה�n>L�m�8L$�g���oȿ}��h�{�K-Ԁ�-�.R�k;��?�=ô��]��=վ��
o�{
�X��	yB��rOT��y�4�ܑ7�D�i*�,�4�ns�(̑��]���G���i�����k@��p/uM�}�|1���G��1ծ[y���q���w� wô�� iu-�rC����lT�zN��7������.Ȯ��r�۬���0P�H��dr"fH��S��\��g��A�\kn�#٬q���At%1�
�G/'��kј��v�9k��Q��h�[L\�Y���B���Ig�����%����ltϵ�-�5�b�w=�'�;�%w�ω���t�I:�7
v5��V�����P�;�v���x��j]qY왕�������[Vv��]��\6Y��;r�*�]	�F�mMЕ�/��	�c]	�7ou箟0us��n�7�5��q���uw]����0xnC��(Rwٗ��=-�g�0�{�Kih�l��2���ͱ���ݍC�J�+|�Z'+�[kVX���Z��ӯ.�T�5^V�o�?C��.��y���t�m�e��UߗK���nRA�d��y1w���D\h��H3q��u^�6�낥�۷��mo7��y�:����O�[�k������������D�q*�7>L�����=$2R�+�]�r��/���c<�1W]P�)���W�v�;�	�}{۬�D�^o��*�\	:���5f"&�b�n9�=ݶq V�C[[F=G��CN����-��W��4o?:Pظ6�;ĕR?��a6c�5�M�������nܚ�����;-�����o�	���aq���g�C��t�sq6�R���b�sx���_c���O<'�:��Omу휽
Dg����������p��%�`�p��}^d�#Ges����X$��,ٝ���MZ��[[sDOE�5�v�*�����ɗ]F��\z��
CoH�X\���c���c.�b^�0�eo�}V);kr���ze�m�M+sj,�;���o�{J�`�cK��^�輜_Cl��J���.�3^��sNN�wE1g'o��y��-����U�h^��f$GH���Ϫ��M��$�a�G��$�j���Y��G�Ԅ���-�*��c{UQ}�}�=�4h*�����Y~�8�&ɡ]2����}��V�X
.&X�ė�I��b!�g���O�fM?<���u{F���`���C���|���C���X���������,�գփ*}"��������8�Gan2�ݑ�h<vz�ˎm�W�Z�.BS%�
$�p/r��{2fZb��ʞ��4��A��@��I�.��ڧ��~��u-tw����#������KMI*�]�&9Գ�r����+��R��ʶ����dk��V�
�z����]�}:��9W+�m��.��4/��i��B�!}$�93�Nݾ�����.����t�o5ofm�Qk]kJ�1	�s-�F�񯔫�E��[�]��;]���0T]t���b�N`]��(�GRA��4�͍ێ�:d�F��u��M#���=�칬х���$Dq�I��c�f��j��{����c����ev�y�[�S��n�e�}b�ߣK<W!Je��|�>2��ڌ��e�JA^��uC*N�xt��&3�7����Y�M�+���gܽF����c�<wJ���¬KA���o8�o�,$%J���;'�S�؋�ul%6�Z�w1�%�h�e��xY ��m�<����6��w�TE\��v9yׂ�FR���;�<8fJ��y�N6�| �F�&M͑\�=�WW�g���
�B�q�?D5"O9PS����c�IO�N�t8m����;g�x�nS��s����ni}�Ly�������|�յ�d�ƂZ�=r�qm����S����l ��X�=x�r�;X
�%|�|:�i(�8���|��b^L6N�%&��"I�Uz�в;�k������v���;o19:�"�������n�fu�Q:сQY\o�줩W7.&m�x�we����6�����'u��˖M��8J;u��`",�ڌ��B�N8L�WLk)����fv�럡V�2jhb����v�q�����^�3��r��I=����*M��c�e٬�w��n<j�-i]H�����{���������}(/�d����7T����.�m��3l\������[v6�ڬ��muёZa��MH����ҹ�vM��y�!�w<eEl95oM���6��3]���u������/��>�-�D-���eul��4�Ҥx,W
E��x\�=q�h�����P0�kkf��|�_�s�(����[;}��j��Ađ;� �FS�#�G �(S�=O&0B�cv�����e�ց�2�mZ�C�r��ٷ6�?5����~h%{;�а���ZI!������c�K����MhU&]����g�:�4��&��f��qvOY�ۥ7��ȹ���hVw�[�U�v�3ɸ4�}lD�������E���g�f��.X�}P�;�zl��_V���x�crX�0^��<��Y[�|0���N�A?n�N�\k��r�j�N��<9wڊ�74b=�*(	�ު�W��r���J�n���z�Ni\���FT��;��ЮvU��!�ol��J��J��u{Jw�^��"(��,nX�x���}1�_k__<���1"��(go�����^��,ʙ,��I#�9��7*m���`�+����h���e9����	�A�cX�¥k���U�C"Y�jy��Rŧ�TkuXbȪ��xQ^E���Pj�>�$x�tE�ؿ{&kH�f����o�q��uڕ��bo7w/�x%��}�<��&�}}���cwbu��
�삈	I�mn�D����|�$P[���ۆVaKb��l�i�;l�o~��1mγǶ�Qǅ1�������0l���8�c�6�Hn�L�[�Z�9���iލ�j���v�Ϥq��v�w}��u_rG��N�u����KHﻶ�Ω�mƁ�N�O��-��q�:i]6�`YAu�+�ͮ)�2�Mze��x��ܱ�`���L�J��EEӳ�egC��X~ۥ��O�x�5E]��E�KZ�m7�e�!�F֒��Wwk~67|����w�U�3��1^.q��U��>O�N���l�?"�Wt��=lҥ���N�赽E�,�초y�<�
uf��;�����WҦ����+�k�1@vgݜ���:��a��^���6�̝ձ��7��\�o�����ڪ��!�ԫJ��]�G @�*��L3�Z]�6�U���nc��dL����^n��[�vy��&^I��;���Q�&v��]d�N���l�^}r
W*���>G�۩.�;k����@ ǣ�Ŋ׃�i7j�t.S���:�혹��l�v	8�m�7kF2<�^n��C�6�xu��]�I6N�ފu��q�=8����e2��=���k�����ݱ���v��1�b�K�ַ^�nf�F�vێ2F,�.�t�bK��|מ���'7� �!qf2�=���>{b���cu����<n:ss��ȚU��ўϥ��ӮN97e�;m<[ΟoZ���j���wlՋ�b='N-����3�R4��xoga;p5�[]t��/bݻ�����pp�ݝ��)����:�j9�����#����ۖ�(7Sڇ\	s����u�cS������y�;�؍��:�	�g!�wn9#j3�;v�[���\]���'a�������Ξ|D�^���hy�۷*�ђS[�����rjޛ�{I�ã��M�j����Au�u��i�-.��^��Gks/��7�ub�Τ�p�>�ͻc=��w'g���	]�M�v�ni��t=�k���/Aq5F�;�Sٗp�׌�v.Vѭ:��z���W��ב.M�ɘ�W�Erv�ڶ�yA6M�<�����g���h����/�	��&�z��탧�*��{����9���g�䓶�+�6�N�n&‫"���Yk�C�`9�i�u�1v�/k��%�ҁkpge���y���۰Bv�&'�#֮�Ί2��lGnv�9�v�^�ݬp�d�v-�-�xܵ�s��^Md�mۉ������;��S�3��s�-ۘ6�X�j��J{��=Nؙ<�m��L�>7i۲�'d�/�cA����W6�k��F�3��5��j���k�Y'�6�m�Ά�U�uF�q�:�N�ce�v��`ꜗ4��E�vȶ{M�1� ���$����ÕYؙ[$-�_Xf�۸���6g$�m]����<��P��Ê�{v��.+�WC�{nv��7J���A���u��d��ڗأ�X�Z_[��鷞��n�݋Y4�c���i���N�ط7�݋�g�kHC�]�����q��jy���k�x��9�iְ��<.�z���=�cUyO����x+�X�n�K�t�u��J\��k��6Wj�����u1��t���j��p��{k˺{9KD�� fI�!�9 ���E-1T��?}�;q�����9�?$x���{�7��.5�ߪj�Vg J]��o�@��q<)'dHaQ��A�Ɓ��s�[��S�T�u�v��ݿ<�hs4��lQz:��`�����J�j�8��w�q��oSn)8!ګĖ���ٷ�cG��e�g��&g��%�P��=릤�Vzz�|(f[�BW9�B�mEY�x#R��k�29
�G#jGG�Cݣ�4����o����6�`���U:g�ȫ7{;��Q�x�Py*�g�F���a�9�o�4U����v��M�B�A#!����̚.�8��s�n_	};ϋ�G�s��<�>J�/��=���e�d�Lw���W�a*M����^�20�ƛx��}q�-�ب箩GP�n���^'[���Tv����٠�m��bj%�N
�<�;k��z� ����B��b����I��*����9����t_�o��{)���җ5�0Y��$Ĥ�M��:��7ۜr��﹝o�
�mn�l�����mӷ��a4��c��!{I��R��h4�P',8�+N౲�	u�q�Ĳ��T�\k+�:~���{yf��:V���O_zWs�_]Й>L��:��(�ފI�6ێ�i5L٪��B-C{�:��ܻΧ��iO���7xU���w�qS0-ڃ"�5����e��KXx����<��㪻�G��J�� �Z�e"�^�3��!{�����hYL�l碁���c�o2�&�E���I �W7@���䯍�كǈڌ�^���Wτ��Rew,��a7
�{����_Ԝ�u�G��>��Xq3�)k'X�aRn�?7'c�]j�.��ݞ�Kv]�
s�Xßa"7h�kq��-����4��7)Nt�/*b������g�YU�����и��v(G꾂Ve��c��m��M���n�d�=��D�$m����bF\�K��eI@���i2��H�n��4����}�6���Gҥ{�2AB\��܎mS��v
�-��g �G����m�W���\��lѯ��wW���ՙ������T+��աS6smRB�ãE���F���T�|Om�T��.�(�ƭ�B�7νP�DnSۅ)�gc���KF�����6p�
�E���RT"�����WNW_W�;�tx��73��e���3&u9�ϒ��N���"���/=h��w�:�=Cy׷u��7���FX+��#Qɾ>e�-r��b�K��uy����x3T��9`����5{x�>N�T�&5x�3O���J����-�N�.�v;��\&,��=G3瞼PO]%��ٵ8�+dd��
4�BYg��'���_qQ�x4�8|�-�<�Ә�L��z.�����̙[�1��h;�EO0�G)�N�Kl�0�J|��A�ɹ��U�^վ�&�J��n����bM��m�^�v�>�������bYs3�I���d����|�m�%�	�OP�WBh3}�$O��v�b�Cxf��&�;�wmxy)&[~a��[���蘾� �V":�n�PF}�R�ys���\�#�@հ��뾮�g�Y<$sYuQy*���܇ut�]����jj�m>�����ؾ���j&�֡�������[�w-�H��������4X�v4�Hlt��X��@0I � �e���AyR���h��q��o�Z�ZwU���fG+rk���F�I���I�Ȫ���I�]\JH�����%;�'�ꍩ.jzE��9�k�v�Uϰ�r8��w�OeR(�A�a$���?G�L��`�J�0d�)��J2�t4��:�:i��%~c�(d:�k$2�>ξ]��?C��"��R!�
J!
p�����밫p]��˚�/�Z��۰��=�W�vK�GJ=���Tv����̧��m\�hFO�h�A��ڊL��H��S��D�8�G!�������0�ռIw����7�'���jحY6f��쐽��$�#��E,Or)8��s"\�zzǨ�$��w���t�j�m��̋s����z��D\8f���E��,;g���G���_R�ۀ��i�cf$�
I3�7�|6��SI{��M\�N"��'���v���d{n�	u�ǣ�H���5��R7�����k�bZn�����l���[F��n�U#r�����ʠ2wxD{]m`���42�ٳl�(Fuj��M�rF�aG��9ۊ�9�S�ѣ5�6]�8��+ӛ�؝�q<�I[8m�&�nvx�uagV���q�v�,pvה��#=j����
��bE^Mյ���������4�>{m�M��m�M�<�1�z�������]�
�ps�k�e�gn�N�M�t�V�Et1�=�'naz��=W����t�2��J�|��E�4��;eh�<E�,O6��>�G��n��M;n�y�91z�B۶oli�#۝�ƞ���ta#m��vL��DPJ����Y�����Y���y�<���<�f��H/Ñ5�n�{��ͻ�*T�������%��B�A���*癛N����.����(���5*���j�yxtk���5�m��6w�.׮�M�aȜ� f9#���������e\"���z�*���_-EYب��s^9T>��+x��
6�ir����9{�*2rXf8�{��7��]
&'�����T�i�uGأ=ҽ��~�D}���z���i]ӱ�F��R}>r: �����Už����h�r�)���OLV�	�5���|K�$�8!��̝0ҽDQȰ�{�����Ւz����_'�ꆩ�V .��)ԍۉ�e��!��� �)���xMf[	�$q	���k6*q>/��kO�[��y!}�U�f(ե�P��/4/\�e���R\X�qAe�a+N<��7��W86�U��˘Wu��(����jK��cA�I1�̣ӯ�6�)�}��9f[�s�S.U�t�\5}���ls9����9��5�iژy7���RO(R܈.�92	��tņ
����e��ާ�8z�Í�W�u?.5^���}�I(��|d�?$��t����rxK)h�yI��P�[������]�N�rY��{B\/I���oL����Q��7�x��4�G�$p^��/[�4�Ԗ�K!g)gO�d͒����9އ��Y�ʬ^$5����-������r1LVxV?4�� ,'&2��g���_y�;�C�P�0gtu�W_�	ڸ~������y�5D�pwt�ė�m䕖�����ߛ�����'�ͦ�D��r0q�g+�d�`�9����5npK���m�.�u�!#n=�#B���Eg��!RSή���ݙ�� �oI̛�U�ͼ�[=��y�U�y��� �{�p�̥	�MU �H{v�������c�!�Dٿ
��=H0�VO���lT�.����m�ڡK���*��μ�ٳ�l�ŵ[�c{Sb����c���5���e3�Ғ��ˢ_Wt��ҽ�G-�u�ܤ��`�����9:5g^X�JcSz��1u�y�;�p�]n5O7+v���(Pn�N�s4K㕻�4y`�5A*	{-؝��"���y_v��;*/�����r�QH�m���;x���|+.L�򌬎��5�5x+���B�������T��qq��л�3r	�^���P�ӑ��P�$���fϟ�w:��l:˳��6kE��2C��6�Ώ���ĩ�k�T=���{�������c U�T��mvǇO*G:�[�qF�sSf��Tpum`�O�D�	�-����Q=y��X�@v�x���E뽜�[�a��<�
j��vm�V�2,����ǣE@�1�Y��R�\����j�W�������1�$[ݔwq����Ҷ6��x�gK�.Vb���~C=hDL��ÒU˧�\^WS��!N)���3C�{I��i�H]�/kuWz������@�3�#i9�J���o��SF3�����p����&�F<��� �|s�t7}8�u�w-�f�a:�sM�W*>Z�\�ӽȣ���)vk�@ۺ�N�N��f]���0s�m�U��b������z>��_HVD�q��,��e�ˑ�w4:�+s�]EƽQ�b�6�bu�=�;�2�m�\`A���u�7I���vw=��Y�G	>��V��c�.�W��f�
}���֌�gn��8��ݮ�c�è�U QYk���^���{Y���-,��F�=�~��������^Q���|0��K�ޢKg�����C�F e)'>l�N�n��E��Z����	*T��m��˫�?r�k�*\�+=���}=���h�-�5��D�J���ꬂ�{��ݐy��;u����2�7����L�H�C�������z�u9!�<*/�BơjDd$(F�(�����܏^����B�x���.�􄰟wL�}�.Ě1�(�{���4��ɓw����I0�J��n���o�[/�t|��x_��ݮ��msW��!>t�E����=Yc3�J�X�c}��4�-S������ڄ��J�ܙ�(�F'�p�\��!�ۛW���L�V�e�L�4���8����:#z���I���K@� �'j����캪�������t-��˩�X�qX�od�����jB��\Y뛇�ɭ���������ێ-a:7#�hL�	7V���x6��,ؓz#�ry�3�q�S��mM.�`qۇ7puU�юN��lvx��]}n{vÌ���\絧A���l��.x�k`�`z�G�Ӿ㌸�n����Ǻ��y��\K��gy�K=8��ɧ9�1u]���[]��s궹Z�ZB$i"T1�l�2��P�+����y��"9�z�QO�(��u8��v[67��pv-��s��z���G&ʲRn5(�rU+s����V
G���<.����(;�R$��9�F#�%;������sih���ֹ��U�j�F�%Y�OZM������](�y��,��hy��ۈ�RIwtjݹNGΖ�<��"B�D	1H3�� �F�� o��H�b��d��tc�~Z鄳�A�[hTA25��0n�d����6�0Yb�qO�)��)�#EI%s~�2��{�d�X:��S��~�M��{`���>3ezłl"�oN��ީ[7!�^��K|�1`��Q@�cQ�ٹ:�m��@Ϲ��o[8ݫ=�޻%]�4vj� �(5j�$��x��v`��NԐ�t�0�&WS<�5m���u�]	�3����ȱ�R�&�ރ�:�@�9,���ں>t%��~��_h���5Ն�oԳsV�ZA6]�Y$Ck%C�j7�&��罪��Z�7ťZ2_X/m5׳/)#n�������e���Xk����j�(˜G.��W7���Y���C	��"B�h��L��ty}�[�?$� ��
�^]�bt{��IXu�.��1\�����;��b��	Q�
g�|���Ϩ���7o���� !H��Gl}<S�� �C���o���GYN�R����Oa�!�Oi��O�������w��^���U��G�l-+!A#�FKV撑��������;�Od�=��xS����$2��C�)Ǿ����;�Pr��绨�&p�U����=�`�'��G<����\�s88�7J[���,m��lU�Ƚ3�mE�v��'p�.89z"��p:�M4��������q������MYL�NP'�K�s�tM��pz�>��=�G����_HH5d�4��xh��{�K�P�>Y/LXr�o��f5��w�VT�l��	,�:��+δ�M4�ڕ��i��&#�&�:�.&l�}P�N��ـ��:�
�]���sA�J��bM��_s�x8jĖ::�=yҰi��V�a��v��qn_u+j]���J����T��6�Vǽ�&3�����4��A����`-vt��%�:�:]\1vPa^�iWP=�,1�G�����3���Wu-��2��ϩ�,�B�&ǲ�hŔʻ�AmѺ��<��$�H驣�M]읆�c�]�i�m��g�n�4��S��d��tj�ǎ=M�藅թ�2�3�z��6��o��Q��8
\�#��.���Ǉ���W1]���@<u�@[��̩KRp�0�!�����aLc���e�3��*��f�x+��T�j�߲�Y��RcIrv/Ճ<^�&$7�l��Ǟ$�2�:>m�{�E.s��k&+���p���L����C�*�K��u���D��������0,Ce[�jL;G���ԋ�fo,��o!�⩼6-;;���X���h�Prۣ<�ʶ�ۭ<��
&{��i};�X���]V��v�d��m�u�{���#(�׻/w�u�ƻ�0��eӧ��ō�����*cZ3Xz\D%y1�����lg^e�҇g=��d��8��u���թ4�#*���=�x[�9�Ϧ�cN����0����o���`�A:�LŘI#q�SV�N���V+���b�$H���Z=�]|ॷrKUul�������Buf��ֺ2�S�
��������:��߱�h��Ք�^��]�"+Q2�e�	ڎE�ڙ �ٝ��J������Z�ݟ�����iHy�H��Z\xM���F��x�~�'���ըh!���N��}�� �z�C�9�x��I��''��\rn.������@ፆ�rBNAoސS-O.}��Y�ĝ���,���uo������A]}*��1#����h6�c����$�E�n	�	Q���%ša}��CP�6���m�k)0�lrI ���ɀ���bw:���������)r�].�0�G'w��6�w:R^��UN�����-ůM2����܅����n9'�j��YBw�*��W�F�G=�j�u{2Q�&-*@o�
6#���3��W �#��pK������Y�|�������������krЅ��VR�V���y6�y��[�Ն���R�(Xr�3�hB��5�+ʵ$KF2c�����	��kv�Fmq�f��yz��O�g����:�f��͗�M��f��fm"��Ƈ�A�2��/#�)��Z9�7�ltt������'5��7��h٨�u>�cs��!����g�P���Xp?v�9l6s[�~e(�`���
$V's�+vH7��]KR������I�=�g�$���� 7��[CLr��`�ۨ"�sE�L~��kvF�U�F�Qk���:�t���ݷ'լ�۶�^���)뛮�y�KZ�yD As��1�W~ޒ�����
_B���"
1�{y�k���=*�/i<���Y��)��*B����J�\z��rH�5pw�3귘���z�VF\��c�ٔ`��ɘ�C�QMv���h�>�pe٭=D��5���MO�$��$�E��h�V΂�ܩ�ג[e�w+�1�O*p�j׏��J`���;u�W�+�2�޻�~L��2�%$�Cm��wO-�EWU�d�F��2e��%c�a�c���2���s�g̕�yy��k�'g�X��8���R�8��LOr��AY�d\�TTy�21�U���OA�G�;]�,c����t[���-ٱ�۶�%�4e��8�i	YY�\&)��+[�OA�1\�|�����,gG,���)�6�t�Rt����#Ɠ��En�z��}��Z��fjvj����ۧq��vMT��M�{u��l�޷E�6���t�kq�k�O����SwQs�n��J�I�;-dη���h����[��}G'A�91�p��k�W&z����2��|$�j�4.��ֹ�]��}kj�ڹ��b79�\s���`
��ӎz�ϞݦZ�c��9H�9�&��:�6�퇅n�9�X���c�͛A�z���������p���ꃃ��[�⣵�x���m{k�9+�N�v.��i�sXu&ӓ:�E������b��ZZ��,�R������꽻��߫��w�ҁ#V���q����C#�}�Mnoew�`��m�=����\�Ή/����b��&��u<ĵa&��a�p��S�(v}(Hc!�Tp,˼}�_]T��sP�u$Н�.� ��/y�l���o���D_Jl�X�/�Ǣ�+)�Ÿ��2P��$J��0�������>����U9;����΍=��49K���(<������)��=~۵f�w� �B�p�*]6ޘC�V����ȳ�1W>~�v�jU.J�7���V�z癶b���'[�C4�vxĆ�@Ս���E9ܱ�pt9������s��U%ɵ���r]�=U�u�u�Bv��x94kr�����9
��X�rr�eǼ�O���k���.��["�4��R�]����K��-Pp�r@oŘ�yJ����J��M���(�����lQX4B��^+zWv�c���b��؋*�PX�/2K�²�2O�J}Oa�Ct���Ҟ!�up0�Y=�uՓ�{yө"C/����q 7��h�
��g��eKWv@�[A�! ����8=u���ꢫ������L�ҫ�g���,�������7B���E�lY������8Sq��O�S��ҎaZ��)�>v�T�0����a����������D�����a���i��X3����X~��А4�4bp���H&f�`�]���!QW��,w{/`מf�u��Sc��W��^-5KT�.������Cz^.4�)'+���Zܿ�;[�U��J��c.���F9��C�N��u�a3��-O�R�^2�a�.���.���M��\�;����azOvX>4���Яun�f��S�:>�}m�cX�e�N$2`jG:�(�)�u�K��j��*-{;2=sYS��Ձ�0���������<:~��H�*ЁA{H�HH��Y����]����d�D��@j��_��>��^dF���ۇ4��;T+���]h�	0�z!y�Æ�����47Lr�^v�۽km�r�e@c�;�v�%-fxQ+K��(fFy�N�QHY)6$k�䂗�I����3cF,-Mq�����JƑS���3°G�t��jJ�1O� �vt� &B�p�C�A]r;�n<����˾�CU�^�t�RN�Ӎ�� t�;@�=�ln�U���|)�a�ݳ=�*�#�"�4H��U1إ$�P��r����gr�9�=v.M�<�`x��F���D\jK��A@�N.�%;��w���<�y ��"��%�,�4�y*�Ax�>�.��i���Ȉ��f8�2(ԑV^���w+ÎoIF�.l�F+���=ۼ�s��.�5��u�IDb���U���ڥǋ��$FAN�~�qV�O�2��fˁ.2�}j��D�#8�˯Ed�[R{U�Q�Xz�R9��tc�% ��0�/X�D���x�����+D4�Kv��}�+^IMEί�qv�PZ� ��R�|�vy�?���O�«�1�l��h�G�d\�Aգ�i��Z��5hiJf�+���-ʽ<�5n��I��d�i�ᬲ�_����e�Q⸔�� *62$�l�ͫ��z]�R7�&ٌ�ɜ�ye ����`�N�^���,c�k>κ��w�9��ߏߠ���k��^���mYuz�	9��ay �c��g湓l�P�\x�d��r4K|>Ň��P��sZ�Ew3w�z7P�n��sjAϣO���DPӄH�{ 8�������k���Q�LNU���8�-V�:KS觅� �oƱ*��6{sȞt;E���~��U�t�kՙ�w�����%@���rAz���:��t�!o�:*�*��b7\��kܳ�}�o��a��{^����W�'UeX�E�"M�DÏyMJ(h�z'��YM��+җ�����U<3G²���T�����${��]�;t"���v�ޭ���Ŀ.���-�1�A�[}�-]���^���D���q�ԗ�J{3^ݗ�׻Pr g��%Js�:��p�(��s�����w+6뵕�v��-�����m驝`���n �0��D��곜���(�Ar��nlޟsF��T�5���V��sʴ�"�a� ��kZ����.F��;�6���+�ݍK�i������6v��r5���c�����.K��;=ձظ�4�-����+tv�ͻn=\u�X=8�Gv�۰p�O=Z�ӷF����b�r��Oc�Go=�]]�i�W-v�r�OI��K�3�7^w��:U�C�cu� �3�����Ҙuƻ�n���w���w<��Kذzw��EMˮ{Ã�=ui�Pi@P{g�Ν������1o��H��f75�Q����7��6����7NeI�F�{|M@�˴�[� �9t_{0�ƙ���n񠹗���QP�n�5-]�T}33��}
#�65�'��q�y|�T� ��qHP�UG����L�?n�=�4����m��I�b3m1�~�ks�nN����}��m
�J^�YtTz����X�Im%��Vt�M0��B}��Q�S��r]�����/̭��s���vAP=v�u{�}(9J������TP��ꎟn���Y\Vmz��']$��?'4���$r
G�:�uI�}R�ג�h�ﯫ��K�x�ewM��ūN�7�����N���w��|���M�l�T1�Y�F->ل.5z������GH�xހ�řu�c��R�cV��ʡk+l��x�g9=ֲ½��_ �^���������U�C�^�>�P���K�S�5�ĝ��qw�&AbI�H+���+��rU�����Xɼd�y&`��MM0�������Ob�x�9�Vdm�NI�ܴj"s1��\�װ�ջc�*;R�ճ<���Q�e�z����B�g?m>��mze��i�˨�;��,�L�±�-��Ki-��O���C:-�<qyΝ�U�W�]w'��������t=�ʙCP-�ۋk�3��D3�ƥ5ĉ'�D�JD�pJL�|k0��{u[ٵ�{�~�$Jl"X���-���m��v��Dc��:����{�	yʺ�M���x��(��e�XBGf�˜w�ݔ�gA/�Z~'1�t�n�l����t*�ݩ�"q���9u��ð�LȰJ>,b�a�@��e�;u�l��7Y
��:�kfvv)R	��dF�G�n��������o�^f���S}����ik�TԜd��:�8����(�.�_j++�Xu�������L㗞u��?�GCnՓ�M�=����=$���O���u���߄06urHQ���Y��{��zU]�Q2��ڞ��otx{+�u�Ff��O�7|�m���c�9N_ ^���Õ��#�X�8n�Y���[�W����7k4�
l۫�_A���v��@%�Be�"���WMg�.���v�ޒwm�e�C{e
_��\;.���冠�����I4���8S{�m`��GM�#)��'�3Fk��ӓ�(���5����݋�e�Oi@ei�#ģ��.5%;gH��]�.���NX��nqC�+쪕��8�֮�}�|�X&w���0o��g���C�dMq�"ԉ`����bhV����rZѶ#�br�u��G3��t���m�+od�¬�긻Q'�՞���5
�cj��f�t邼-��~���4�F��yf�W�-��׼�6��� JF"n
C�ʆo@�<�]��;\��g+��-�-���C�]�JfK�3RE�zz�uf�#86/�L �V���C�|a��8�����9h�s���i���iN��x�2��Y����X��]�v���)o��ѧ�QP�$���j�J.��w�_:9�~2fL�I�{�0E�,ک}ת�fE'��^���T)��}�Aili�d���v����6%�3ٷ��.�v
l��
��{%+# oS�:mmd-���B�\@S��L�s��[b0��wۼ�� fy1`�n�IJ�0�kL�`X��A6�Ϯ���R��}�H���g�5u�Ε� xr��^��`�����!;\���8{Y;n��Fog!NYI���+3j��kK'L�vT��bZ����~_�E��ߕ.$e�;��ɾ���	�4�vG��[K�ϼXZ"ݎ���ʢ1�ę܆HQ)9�ҥ���9���[���]3�tf�4��rr��D'�1Ӌ�*���6V���v�����7���e¤I�3��bt�Y˯ʔk*�Z��p3�P_u�E[��z�%�%�p^��V0�N���}.k[@�?�������*�If��d3��E�=�}r�z��1��u������Zn&�e�,�鋣TwA�۳�.��^���~L���c~�3�&"�Bn
ک�� $�rŏ��No!~�x-��d��н�d�W�7��U��Qo6�
������X1ʱ����V���#�vj��=s�Fպ�-�*�t��VRӪ
��m��{������k�t�g ���&eF���[#�)�Z����My�˫6M���ھ��͡���%�n���!ߗ7a��$cvK�g��'o9��V�P�$�zP���Yy��0;A����hQ-!w�p���d�V����)W������w���;����fz{Y�.gn�f�AC2��;�ޅ�bvT�`����Wu�j'g���mQ��$����_Y�1+��J�Y.�W^R���	d� �Ԟ�:��|�����d�b�HQ��4T��%7��n���]޽��IkY#6����	2��˟\r������K�]����p��B_ǣcxZҤ|�>śH�VȦR���:��U#��s��kT�+�G���:��p�է�U|��w�s����d}���5�޲,���a7��ne�JM[���"�U��Ž���tqq�w��'���α����C�6�l�|r-��ݴ�ֽ���RJ.��h܎�K�Ѿ�25X�e�NG�C1�B�۫A�fu��(�Pr��im7��;/r��5V�=_��~�d����Mk�0�	�~�a�A��"�V�S9~���N��,:��kk�y㱨���n�ke��ہ*9�bn�l�H��41�յj�0\dtf�e��tq�v���f�%mf�����V�i}�d*��MŚ��Ž�n�Dm���Sh[[��G7�ui�9�l�d,v�,�Zݥp��6��m�6��Si�)v�yg�ۭ�O���u�l{I�J�s�Z��;ew��N��)K��F.�!EbtCHU5k�
V�j��=���]��ج���ֱ� E�Lt���*%sɌ;����/�!�=���J��l���P��c+xh�֙��.U�i����xݞݧ�ۗ�����f]�m���%]�\��g�-��PM��x,�r�r�v�n^��Xtk�l��6˸Q�;��ji���6�Ag�,>{v���N6�#�sa��c^�ݺ�=��%�i턱�n#��qz{Dk�t�+�Q�z<EӹL��F�gg[%�Ѥ�n88D.4��Խ:�f�aKO&����֣ysa�D1��ٚ��g�.z�P���Ѻ���h9����4H����p2���,�/[F�=�g'VT��1�=�4�s�ێ�!�<`˼�6]��*�(8^.����t��C��{��nun�O8ޗ{?�|���m�����E�'<Q��N�wkO	q��Qڶ�:�ݚ5]�c�뀴%띹�>|�
��L�]��ܜ%�.�ݝm���w�N:�ks�[����q���}[�wma���s�1�!�&�cX�m�s9 _�|�/��ԛgQ;I��;!N��j�>��{z��f^8mcm�G4bh'n!��0�vW�nN�RoF��n�oX�]X�r�E�틀2{�7]�{u�K�����}��v[����$�r���Lp�m����^�s�=g���s���Z���Kk�n3�g����`��t�n�5�u��q�[0��E-���ټՎ=[u7��5�MN۾������ŵ�:��)˺|Za�c\�¶e`�m�����͜b|�օ=\�k�n>��b>ܧoBQ����^��ݝ\띓a\�pل;4�J��E6���� \���;h^I�q��a�7Z�[�]ι�z1�U�:�셷O*uխvm�����;�:��ݚv��*mӳ8�;�����ma�K�TWv;\��A�-��8�60��c��y�g%�s��q�m9`�X<��G^���zzݢ�9�T�Y���iu� �ēs��Q���sDv���.U�Bݸ��f9.\� �guz��vHS��u��N�狅�N2Sv�9C7\�;jT���h�4����Y8�;w[9�·���[q�������:��^�������[5�E�s��or�H���z�<�\�{l��u+M:�;�%�ugzك�Su�V�n��X](��s=��^�M�����(��uI��I��+R.�ٹ����C��yN�qx��]�P�Ӻ��Oa3�>,�PU����),�b&]����#v},G7'B�z��`��_)Y���S���bh���_K���z�ɷ�7Qz�߾�U�B�,�{v�T`�p�s���4��)�:��~�oJ������\����F6��U�z�_"���QY	�����rIo�vA��^��>Ӻ2�=��m���m^�s�eH�{�]{��kg68^�,�n�����?8��$n(�p(J	��ȇ��=\�mV,��a�Q��Q&�Wy'��c
��KVN�▯Z��oQ�
�u鎶�~�{w캰�6\��������6��u�xM9ޞ!ݗ��(\[Y6������ܴ�c35��S����cH}�i�2m=F�O����3]�c'�Ӧ�8���������^���DzGd�ѐ)$�b�~�[���s���~˩g�hx~�)|-s�3߷����f��:�Iz]d��hE$iq)VǷeCY��t������s/���rh�Y}�U%�^'��0��f Nz�ok��d�ĘWfn���UV��%]�F�N�~��+���ien�V��|U��,�x�`�R��]S��9����P��ٷ�4G�N�/r,x� �$d�;��:r��'�,h�>~���8�:�Z�	}Y�K[}}wę�Z}i��]l�}ޗ�$V䃺��s+|6��OGEu�
>d�x��h1��
w �A�Q�� �X����k�B��&Yg����Y��NwW��Bk�5��˻��eC;f|MBc@��y�o��x�ci]j&��1�..J<�:w��H�۳���ۍ�tV^�ۤ���b8�m-W��;=�_�A}q�W�P�U���hR�ɑ��LS6<�A����Y�]`/zYL�� �pѲ�����P��3{�{-V������:S+���S]�Gا.�p:Ƃ�s�޻�_z1]�1Y���[E�F���Q�f�5�_f+�S�[�_]�Z]��b�^k�}�IԼ\�s�x&�Y��p���`6bF����2�\�6e�6���E˔�,�U����lK7{ӷ������������}��j,�	�䱢��Pr)�2U��N�:��\)�p
��y^j��h��Ae�L{���ƶ9�+�Ĉ�i�����K
ձ�
���T����W�U�=U|����U��A�����nW��^I[���GW��*x�Yܺ��.�����ߕ�6qT
�(i����)���b�q'k�b�N�եy疸N}g��	<Y���H�-���.��/�b����!f�/{���o�@�^1�|Q�f��0�*��m�2\��9�*�e�K�f\�+n��C집��'�D�� ��{��ۻ!z��ҹ��;ʨ���nW`olc��=w�����S��mÝ��ʑ��"� �4pKm�<&��6��o��1��(z��ٻ�׃�*�@�����Xut�i��Te�IEn9#�lcA�.y.q;�i{2��$4�ްw��w��A��a�yܗ���N�훞P��{teK��:��+�{���DSHr���X���qӴ5��D�R�wHu�@R�b���T)%b��|=7��o���/7 ��`�'j2ҟ2���y�����v�\u�'=�'G`Yq{8ɨ5tV���(�Qw��!zx򼸍��-_}��&�����(�p��p��O�d�*�
��z��&��e��:ٰ]=�u�P��Q f'�Q�8F�W7�rw'b�f�����{����R�a�{K�a���tJVzWx��m��6i����fVӊI�$�x�#':�)�}3V2�n.�ŃS<�"ˏ1;���vJ�O���L�Xk;Ɗ�Ć�}d�PȤ4�)'$���Jz�W+���ťk'��Xz���Jf.���sS��Hz�D�4Yh5�w}�:`�}t��#�*�[[��$�l�Ȼ���S�cHե������^kvr�<�ۜ�B���h�7۝�����kR��vud��������ӰV[_w�~�P�2c�p�^;����}��˂YK���p�RFz��P��!w�{�pԺ�Cjp(�oX�ŗ�U���&�	�ۼ3h,�T3��9cc��'<���;�9��{b.@*�ѻ�`Ϥ�_w6k�d��ڠ	m�MPm�m����.˰ݍ�{P�;�f��qUb���w�a��t�v�v�f�sf��f�۱�����`��d���B��.�-�:��� y���$������I��φ��<�j��	w[�<:1���k�-�S�;<���ہ��3؊�m��9��n8s��ln5�=�vZ�u&�`��9�87 ���9�1�ꇓŝq]�]�����{ǰ�n;�Lv��I�2v�#i�k�^8�zu�
jx�ץ�-7��n���|4���WN��sȴ���=�国8t���}Oَi�E$t8Aަ#((aQ9-�
�w׭e�Y�o��q����zi�K����5T�.��L�59��L��`+t�S�K�@���N��R�e��9���5�����GF�蟸{���JP�rP�%ft��́z�Vp{���e�)�S�6�)�ґ^�<}롆�Hu7\<$۾�}پ���x#7x]<%Yb�a��|��do���XyQ��s#�\K�K[�, ��$"�'��1�Vn���1�\v�7������}O�ǻu�G���e�W)2��=��y9����x��.s{Om珌���,�e)TmI$�!�k�4A���n�Z�Of�����v�����F�n�@%t~���(�­�}-��lΙ�5C]�竳%e�X_kY�lt�{��r�� �g+k��䍤�m����G�q�����R�.�(���ej}u��eA�q�3NJyK�Tl�q��J�L�k[gM>��|6�ҳ��.�+M�*���g�5c[��<3TcY1�5��g��{c6r֕�=�oe�4Oe�F{5dg�u;��J �T�>�/^�����_O���T"�Q["t*����TD[]*�o�N���������{L:�7QN����;@g��=�~U��ѝS����dtv���ڡ��� �U��uQ;]����\ZIlWN��d���Ž��m�HD"��h��a�|C=Q�1Z�y���h7�G]�S[�ʱa2���zO��.[m�wt�e̦�+싥�e���.�N��0rv�FU�ʞw�-�9[鬞��Vb��w!��:����@����j�6�ۋ��s$FKL��賶�We��D��8wIm��ۅ���l��D"b@�j#1ȁrA�Gj�Re�^�q�l)�-u�wdy�ow.2::�ұ?Y��ޑ��T�y�	��ihg_.>*)Q$�b��Vw��']yK���LZ�Yo�u� 7qkY���fi"i����I{���{�L�+g=���e^�J}Ef��K+D>�MB �HH�nU��+������r��nɼ?<�8����T?��)�"��[�8�zuC�J��}h�Rݹs^N�o"4�kz�S�f�
=:�������ކ_�B��j����`Ly*r~vum{ ߳�e$Q[���|��Γڔ�w�Vۉ`Z�3
�	�P�rh^�ՍP���p�ݪ<��ق��ywq}^'���;]�������PЪ��B�]5�ޙ6���`A|��j����YJ6ۃ0ja;=+�=��1�b�S�R�hfV�K�=z�gj��)^w_���fiv��5��%���*Ś��r8�v���6�[p�μF�%�☮Y2��ɝ۷��m�<����t���WoN�\��e8<\��=�]i�����s	^t���mշTzܡx!;)�ޑy��.'����Q�!4vӊ{
�P(Z(�o���䚧��5����0~�$�Ϩ��S���Y�(�@U�����My�u�pF�{U,¡n{o�%ϡ��	:<�����4���.G��� ��Q�H'��{���*޽<�G���R�-�׻�3W�"�P��#x$HFZ��"*H/=!ڤҘ8oNjz]᫨������!��^W�ڥV쳸��,kîy�K�i��#<UK�k$��r�;�u��$G1��N��zpC��&�G:�72��B�J�P�4�WW�,�C��ìr���zꨄ�x-B��Bn^��6S��o7��M�L�$a�޾��0J�y��W��D
z]M��x`�l����wz
�{���'{�)�'tF�w���j�����@�a�H�u�5�7C�Y8��Q�c�������乲�:��R� )FY��t�\Õ�p����*� c�g�u���$GW�J�}\�>�v]�x�&WC��r�7�j�v�R9�x�>>����Ԁ�&�z���2qe���
��y�w,�*�_]{��,B���eje���T����J��֮?�eC#$��f�_��;���wX3.��Z�F�o������k�%ymD�#z�S���`�$K{�ػ!��`��o_��.��ӌ�s�2.�O[y �oS���+ٙ��=���_�H�w}���A�Cx퍌y��+m�䄾g9�0G�m�e��i�4aʯoM���C�J�ܥ�+{��7�1��4R�<�:��)`����.}E�v�nV"s�4�	|�z�u��YI�75�+Av���u�Cvc�]��1�. �ͺ�B�����մ��)��ӎ��^���,��R
*;+�wf�ێNo<��l��=83��������;��5�;��2�v��o^���v�:��Ξ	u�����8�n��g���wӌ��˵L�v��]\Vޮ��;���Kn 7:��ݛk/[��v�]/��ZV�]��<'��/NS�f�v��/��,,d���g��yx.D��0�����vtDmyz�O�u���9��]��w]���M�6�ԷE�'9ci�c�9��o;`�-DRI?x�l��{�~�c"���&3�.�8�6�^�d�-�Y��W!��Q�H���L~�KDu�/<��$����r�y�44��չ�^�o*�y0˴���@�̎��NܨUPs�/1�+Kk�\bY��(eR�K���_��L�W�k�_a�U���/呲e�P"�zU�}��������й%�	���z�U5��<��FϚ��������j`�����G�|�q����r�^���w���YO�]���c���L���d��	zӬ8KAA�w��[l8�23E¦K{�=�ݏ�h��U�
�^���M�*wa��t���-u&/�lV�Z��S ;��U*Z�z�������9�C��!�š���ktNS�Wv�og�9��h���}�э��ӈ��#�˭��y���[I��񼼓�?��OK�w#QoY;�տ�I��V��r�(:<U7��+�%��W�Bх��& �CD�]�fo��Q��گY�lN�c�u�cխ�I�\��G����I���U4jÝ}��Keptk��O�b�f$�!u�_K�%Z�<N�]��V�U�H���dw2����Z�ON��r!�"�*��;����w=ʒ}�S�����:be(	n&�:Â�mѭG�X�#�*��k-�mh������V%=ϫ\��F6��<�
�$k:��_a��yJ����tk��"=���A��{�������䮬7�y������ޕ��q7ٔ�DG�(_'�f,������:_X���8���2�@�{:U��G��л�V�2ѿ]"���DnAww�챍�OUY��0�3P&,�6OUt^��;����αF��T�,�<M�x-l}�e���v^
��@�@D#�[UlhI�3���+���WhW��k�t�/o)����Z� �ZޔZٶ�^uZf��v��Q���G� ���Bͼ���'�u�{��:��jUʿ�e�Q���Tl��X�]��B%�������w�3ػI�+��r��(BD+e.~��>��)���'�+��[���#�"=�졀3��,�[�f��Ɨ���ۢ��g��D�eC�/a_|��<g9���jdV�\h��`�D��&|0�9��_����<E���J!U��,.=���c��b�,��j��ue]�a����z�f��n�9V;n�UIf�f�ƺ�,H�w˰t�y܁�ӓ�s���gu�C-'U�QnG�XΎO�w�lW��B������b����د�A�[�3�A��wnAm�Ԏ��^]`r�i٩,V��|�~]gip��B6�Ise>��K;Ns�Ja�*��|{p�^�.9!qT5VnMC��Z�}��s���o��0=�^T�H�+Y�:�e��dv�ay�8�\=�=kU�>ɾ@�V�\�iQ���eh�)j*8'.V�O��u���)w�^oʒ�ho%w3U�����(��\ňU�g9$Kv]<P9N�����q5/mD&7U��f�n�)�z���֤3fT��؆E�����,k����KR�\sJw�<����n��8��Yc-�d�Y�R��Z�j�����c�7[����ML\�@��nW�^=��O�f���������5OeF3*�r����7r�6s8��Wfv�q�</�*� ʭQ�v*��6���11Z�ɍWʉ8��5ܙ�Hއ�;Xd���"�)�w`�۹���Xh���-�v�UE�׸e�f�^|��ʹ[˹�����ћe��-�R�ټ��ڴRc{[��er���z	�|��É�M�r�*Л�[KK���|H�Y%���l��
�=�d�K��p�ۗ2�:���v�5�����nS��%_s.�q�:u`Kmڠ���)h��ڗ�Xn]��-Z�-M,��1���p��8]���u"dt�ⶁ8՝=w��_z
��{���蕋�Zk�;�e^�Hd�'M�Kmv.��P�al�I8o�Δ̏��ڜ3��pO���M��
����2�c�G��Z��9cf�%?��j�H��Ε��^�i�)�ErkV.u��4<�8�-FGc��=�'k7$B"PI&8<>��菑�5���m�9_�4T���[f�Vԇ�W�%�����kX�w�UD�="���D;]�
�_}�����?s���t���0�܂k͹���BAT�Gc�"�@�gi��ͷK%���e�����&ҏ\~uQ����q�>�Y�(�{�ҼG�����/�����8�P�66~�#r�q#7���ρ���M�I�!C��W��ȫP��X�"�W>�\��eJ���������0�=�|j��{����ۓ����l����}�6~gﬀ����d�y��@xMh�͓�LJ�t-}��]`�~"�{�<7�e�1�~���I�#?G5�|@�(�'�說x,#w��}M)�Q,*���N����w^�Lnc�y4x�����ze�8DH�Ĕ��貦�;l1h�54�0�`�Ffgs�����q�`x��?��W�+z�6d�!��	��N��n�B����U}V���h�t�DfW���H��U�Z;����Ϙ{�U��������.#z�iK��k:��S��z���(�W�._ [˖vT��ob�U��Ȉ�Oo��a�Z�&�����*H��g����PDa�$N��G̴����?2�oJl덑f��i�K35}��V�K�2Ge�-cI
��U����H�8�ZE�}�X��!��҈��P���u�3���WQg�^�n��Nx��<��b͡0�g�s5گ=�R�� ed+���*���o�k�?�3O�9��;�@=���Pe*�I�]�D���F�g;o���ؓ#V@�*�Q˼���y�ڞM0��a	����Uw� V/���� Hae�ߠ,D	��ԑ�᯼}YP��:��@�_s�@Y�v;;����𧅌#��=��@���}dC��D��W�F�J����Qܺ���Α;ߔ�Ó[�x���>������c��#���� ��@��������(�־YDr�a��4V}uqo! }�3`+34��|6���j���EK�"]��<i_w�V�.�ڪ!s��"���d��z�D~Aϒ���s��	2�w�5�ߵ2Kc�TGHI�*{�k�]�V,���K��-ZK�I�t���S�1Z�p	KW1?G��w��)ng�{�+�m|v0�Q��M��-����j�",�>��DЕ��$�}��XB��B ����\:����
g�A�`B>��ë����Ѥ>�	��䜃�7zW�A#��@��d=����t���V�Gk�]�ic�os2�PO3�����m���%�P�ît�7�ח��0��]�YܥH���cz�#��<�e��PF��4�l���!C��g(m�e�y�}v�G�N�6���:������m�:�.�S�r𫍴��<�r��۵�������@�
�ڥR��Ӓ�b,5#O\A��%�h+۶����+����nS�r����K�;A��c[������t�O�&wX<�
�� �
���]v�f�v�{S�%�n�]=���b��ͺ���1�|ݻxkB��1�<s"7kv}v|�Wb�W��Н��QQVC&\։x�,�d���pH�NA�����^�^#]s���dG�ZD�ʢ&�h�v��<�x���d����
�Ζ>�?g�Oϻ>OV�`�����B�6�_O���'����ś?
\��1��.IA���?qR��g��|��{,����8��]�?^�T���"4�D����7�/����@�_aÉ�vv�@�ZGEZ�*#ED�Og�j�⶗���'���~��""�G�L㙙���EEUp�a
�"+�I*�_U������Dܫ���ϱڌx�?of��]a�ok��?����+�R!� �}c�e�\�@����v��8�v(���$��xT�4�Ê4���?2���;�Ϭ�}��=�_w��Ys5bKI�	ZFgf4J�D/���qC�K���į���-y��J�+n��A�e�o#�/��7��62~	8~9������>3��Ei�r�Zİ����	'�;�>���J��|\G��e�t�(�S_&�/����1I��p��һ�~���:�m����~RCC3�q�v�i�a��?X?B�գ<����9��Y��p��b��R��N��K�����<1�V��Y�ݘ�A�l� 6����k�[���|�q�	`��}3p���b�&%��	|B�Ϯ����� �rU�{ìu��x�q�q#l}� 4�W�,��
�[��⻍�=��:����x!9���0c�7��t2�@Q�Q��@��w�Dp�o�D�;��G��(��uӺ���ݘ��3v�� Ț������G��MJ$m��r�ųDT~�����0Tҍj�g�U�����p�줨@����hZB�I��D�_�V����H�"�ѤkBG,�j�#�e������J���4Eł�:��y*9�!�\�ʕ8*���'B�ރ�E��y��WF���N�g���!#��Aws��-����4��-�9Dj�����g� u�ޖ':���p���"r��D�_>�:T+v�m[Ƽ��N��D�᜵��ͅ�Y�T�s�-�j��[��;9ߜ��vX�NT+����W����e5��g���+P��:�tW��\h��7��o�I������_�Z����[������F��Ă� �*:s��׼�W��Z��ZDUrb����/��X��u�����C/�����f�^��!-T�$���"Zt��;EVY�����U,+�T����P����\��������3�k�m���8��0��IH�o��i �=�`
8~�����m��Q$�$QDr�]��j��p$n��Y���g;'���coc���������>@"��~ö�ӭH`#�y�(�;�J��ӿh���F����Lu%��[�0���0A+J��@́_�N��*!I|D�����Ĉ��0�#�)_s�%�y�bB7�8n4���g�?S��9��y��ː�;����B:�: x+�{ђ����K���LH��,�q�Z���	O]�q"Mꊪsu�L�V-�H�ۚ=�j�i��^[Xb�BH��d�(n����0�U��=���U��*\Y��[#�f�<�:�]oZO�%�I�����ew��>{�R����4��	k��@+�V+�dad"Zg�;�@�%� lFJ2A�!�ꞝZӺ@'���g~sq���V�`��D�V}�\..=�L�4;��h��ȏ��ZdF�&�0,�6��Z4m�!��5X��&��� �z�?n�/vFHd�*��<����S�.�Y��{?]Z[��|@�_��:彾i�X����3��2S�]�k��{���_cv/��+�o���|��^����9Q�9v�� ��{(;����ؤ6�R�x����5�u5�i�wn�Ǒ���Zj����PL��GŞ�0W���	C$��7��k�<�7E}\6��(�۶8�Jd {av@�%x�:_J~����B>(��,_6�����f%�R�Ä���}XeB��l�h�[Sx����IϜ�dY�d����� g�J��/#����w_���P|�Jc��+n���o3��w�bH�a��=���h3�>�Ë <-�@G�!������8���m��o�RW�lx��9����:9���Wк�.	bx)#:�i���8)��?/�c8��2�YQB�6e�c�����!��^u�x������v�X>S}iYj� �̋��݂�X��#ݠ���X�X��!�B��Zʹ�=ߴ�H�=�G2%����/�;��]�<�3�v7L��s/��;0��X���k5���.Ѻ%<��Ľ����/Zu��F/���Yط�~���i�F�-�?.�$�J�������t��U-�������j:�r�3���FR�#[�N��l3����fک�ψ���W��Oۘ�Ӕ?
����Ry��?���a{*����EB��8���1^H�>�n�7�㑀j�=s8s����A�Q���!L�%fp�@dqdx�4�����`_��3�H��\�u�2ӓy�l�l�5��R�؀��X���0�ש-�dW*>T�p�5U3MR�Xp�8�̒��{�倏�ұ���;�}�!o�}E����׮�Ar��5�%	yZ:˂g��'�5������<@W�w���ޛk�D/��=G���̍T@��|F:ŰE�(���L�K���D��z�|2/������{��%ó��ղ����&'֮PS�S�}�3E����6y�P��>l��I�S�P�g�#ğ���6M������i(��W�q�y�0�[��T�v��]������_#�Ȍz��h�uUm��T{x�nυ� J����x�ww���	�=و�cfG%������Ծ 
�U:ɈkB{:O�Un��]>؃j�h���)�GL*!5wwp9��p�\2���E7�v\�TC�WПP����p/����v��F^|6�%��w��f�}�;�`T{{R�N�vYװua�㘜�̻"f�\QF��njf^?�������V�-.���6r���ݺz�W�|��/�gR��==k�p���c����n�k<]��Fy1Y��Y����;rZ�7(���p�{uێ�m�G�ۧ���8Ml�9��]W!ŋrqֲ���]=o�웞pF���d=�[�+q\bM��Oܟ=�.GGc����s��8�<�WCZ�"ڭ�x6��k���֐�a�T�u��7�+5��]�@�f^��5�Cu��7:���'l�I��#3u;l;�د#�&������}o~nw#Ǳ�lޭ�PfMl(�l�m�.���Q|��JՆ��jgo�W��6;4�]�r�����Lp,��j�	�{��0�!d"O�]�B��C6�RG}�f:���t�vU$��u��y�������\�C����̆��$�TpW}r�}��p��p��h�ݐ���]��?]�i���=��J��D�	�Μ]rqT��T�)�U[b�k�~�|��tz�Ɛ�����T�9��]�3n��YHsa�T�G�	��t�|@�B#�CHF�޼�)'0W�^&r�#1���l].��\�5��~���������誊��~� HI}�C��ƾ�Yt���Т7�XUg�!̀�o�wo�|♏�?e�ݟ�n�r�)�١7�� ������K�"���E�׌��$���p�b�H,�lRp���dM�ح@L@��>�I��x�v�mzP�&~ن����]�P�2��n=��cI�1�J����kQ(S.H�}�c;3{��>&���%�� O8)�q�Wc�N�N8��؄��,����-��Y����]>�X�{^����������>=�ǻ�%�T�i��33�QD{���[�P�V�}I"U���۸*���O9J�w9[�k�]ڣ�,������N���Ϝ)�?Q ���d��Q����:Ab��{���4���i�!OD�߳+��<�b�t�ś�ئ���s2��E�jxi���~��(�[1���0l�F��m���V��a���b�^ʜ/�xu�ey���t]K��>�R@{)�Wz@D	=��D}�	���'̌� �]d��L�e�� tC��=�}[a�E��A�	檎���6ȼ�أ3%2����'�VI|M������� $��Y�q�g��زaA߯e|�����1 +����چ���Ĳ@i�q��E�#���!�QB�P&y,�|�{�k�F�/���F�/�J�"ݘo���d�P�\4�����q*r��|-:��Râ߸�Y�m}"[�z�~X�E@Ki�$���wC�e[{>����z_��@0Fb1��V��r^�o����Κ,�U�>g�r����O�vK?�V��_3��c�B�����
�%5�/����"�آ�8) ���{EȪ��]u�v}tX�AF;m�z�e������:N�I7���?6ߺ��e��S_M�i�������+v}G��b�o��We�'v�lzM���/�Y�BG��T։����dF�uՊ�������u7(�Z�-��K�q��x
%�|�t�@Cy�זzg��{�� R c�~gl��'w�rYID@T���_��x}IMC���H��:��N�m�}�K��sE��������E"l&�Nf%����h���zB�젺����ܕ�{2�O(��K���r�t��y�3Z���xTڈV���|��BþUu�"����i�W$){1ݙF`y]�蠓��RӼ<n���u���lDq�.v[�U{r�����ע��?'	�u�	k����W��,>���u�C1��d�v��dģ"1�XDY�{m�00�Z���2�t�/��u�3�p D	$��]��쫆���D�G� ��8��=�'�qk;ל|?e�Or��ƑDNAP@I���-���(f ��@�����>�~��l#�ϻ��]��_�eQyS�l�9��p5�u��ȭ���c����,B���K�Ұ]ǅ��=�n~�	w��h��P��|s��5\g�B���蕈Tp�tv�����s�㭤������>�����]�D�H�}c�H���R�Y{�5�T,�n�����{[�5B�u)�"��^�ռ6�xo�<��!T�ۍJ臻ow�Y�@n����e4C$�@be#83̖e��cH�t�G�2��-���}��r�����NHj�c�R fB~$^ol58'�q�\V@�H����C���@=�ų����/���#�߮��@�� 붩�Y�z�=�f�3��+��t�L�hF��u�D�QpW�T��\��}E5�mbC�v.���;��aB�5��PU/�x���!!�H�I`s�QU5&�
��Zpf���M��/�d��0.��L�yfYT=�d
�2)LY�"����nay�g�m���O׹�j��%��S��]��Z�Yz��]@�̺=�:��	�F��i}�vׯ]^��,9����6(d���{:U����	�U-S �,��F�H��G�>�EY�ʷ�@H����]�4��}wSt^�h��"k�E�L��EQ2m[B�G�*���{}(/z@R6�k�.�[3w6��e�D��gjJ7����Z_#���*�;/\ې�o8x���Wy��gg��vɮw]��(j'l�-�=߬B�"�:&��6���G͡�$��D��B�5I�7v�� D�w�o����Iew(�s�?@������Df*"�
�b�`�b����N3Q T�U�wr�,���B��t���o�F^�˞d}�������P�6F	�!����[@{���I��k���{~>��ֹ�n����"�lW��B�"d��%��?��b�U�G�<�z��)&�e��|/v�����1p���љ[�68���
ϐ�6���"Y�S�J�� �F|�fI%o��4�3޸�j�^�`����Ȼ�JE)��%\�������U&z���9�S��n�%��J4Q.8oS����s�5�_�Ю���`�E���U2��fwc҄��w�Z�QM��������В��������$�DG�BJJ"!�JJ"#�P�$�DG���$�DG�(JJ"#�P�$�DG�BJJ"#�%	%�𒄒���������BP�QBP�Q������a%	%�BJJ"#���$�DG���$�DG�	(I(���BP�Q�(I(���1AY&SY�ԍ>�UY�pP��3'� b4�t��v84�
*�R���F;�P J�ww*����権�Ka�]�	"D*mL��㚩A���Dm�B]�P�����U@�TPB���%�T��$JBT)@ �
� IEJ�U
	T�	(� �T��mR�� ($�*��(U�O���{s��������ɳN�˾�a/=ݱ�!��T�K{�ͯ}�m����^�M'�}�G��w�ݫي���Uwtʠw0�+JN��(� h�����7��eT�n
p�c�+�����c�t�Vkj��[�U"�:ҎN��;7; rM��:��UwY\����B%=�EH)ARQJUQV�K��fZۥv4]aѦ۠��,� ���
s��kT�	 b��!Sst ��n����v7��n�(�T�G�WKk����U}� :�^�PFP�P��T�ٷ\�%Z�Õ	�n�]��[�J,�͍]��o]�X�G��z()#��h��  |}P� JQ!@ ���{��=��J�aAN��]�:�CCš��
��A��@,� ����t�`<�P�(���x����kފ^�7Y�X�@
��aB���iR���A�/�2 ��DF���'w�T�^z� 9��=�B�� =�� �C;U�u� /.�^( �^{�@
l�=���`�G���  �@�j@||(���A@)E_
x�M�]�IF&�H�{��PCY��.��l��-md�m�-�4�5��IN��Kv��l�c��Z[��R�*� UG2����+�@f�E:��Kl����lV�ϱ����zy�64� �Õ��QJ�u˰�Rw3�!+uέ�ĥK� w��
	R�%Q!%#r��"jRP7X�Cm�r�K�� t�x
Rn��w7I���n���n{��ƚ�a޳�yv�%�"*��oZM���G��swq�;�"@>ڀWh� =���aA@ ;��T��P�θ=�������C�,δro��Gϱ� ��7����u֮ű�������^�wrێ�.��j헶���}`}	O 5O�*T�� �)�LIJR�  S�bjUHfRd��TR�   ?�SFT=@  z@��MF� G�~?����Y��9�a5SyNO��c�e�36���|��FO'+􈈅
"7�]����"!DB���	D%�""!DB������
"?X��Q� J"�J"�߿$���?�6?V��[����œ]�C��t�4,NRiҦ7�r�V\9��P��[W7r,ai7��Ul�V���d�LZ���oa�kM��YmX�Ɏ3�N�&oR�u˦b�L��N[6h�SJ؉m]е���MK�Qֻ�v&C1a��@�uT��f�M���˯C5��%,')��u���͍�u�w���+dW�跻Wr�n�nHʤ2Ƨ�2��oY�3v�o��8�Eujaq�n�7����r�捙�I��K��(����RBrJ��h[(|����ȱ�	)��3��7-,c�'S;b�j*�2�.�$�7���q�<W��q�B�3p��bm�_���0���%%������¼Pf��[P��Ħ�x+d��Wa�0cQL�&S�%�`I��(V�eŏ%�G]3=�k$2�0U;m	���^�y���8gn�](�ܡ��I�Ò�hsB#cA>0-��~�ey�'=u���ZmI��{ۛ��	n�=���{˚��
M�̬,�qi�\nN2og�w��O��Pp���v�ϼ-�4]�P����7M�r��a�>Ң�^�/=�nu	�Y��]ul v�c���3k2�yd�t[�9Z�I&��'��ԤO*?L*]eEE����ܢ,�nyf�|�:P�zz��4���v�#j`�t�c����cFTN�:k.�f�c��%�K-�m���N��<�{lb�	*���D6�]�aîO/t�'*�!�6&nnN��j�t���~t�n�	�TF!R4� ���`d�X�r=m`GC���ݖ�rp��y��\:9���0^�X��r��L �Qg+**�P����~�D��[ػ���i�0�ُ�A��&���v�u9ҁC���f��@U��Mª�.��F:2��/�%�N��8cX�:�U�L��XI� ��u�s�`ҁyx��h��Vcڂ�ɪΊe�{vovw��p�k7u¸�˞F��W(ʙ��HL��-g-���� �Mn�f���af����ѧ��+j`���"�ʴ�-Í:�Rej���6\���m�����e��ٳ���k.ֽjFK������.�5LZQ���zؠ嵴
�¬m���~mcwu�nٽ�(��Kr����+���P��k�bubT�*:f^uS �/�[���=�cڽ��0��Ep3���x�,�Nᤊ3d@�{&Lm� �#ŪawW**ٙh���ۘ˻Z��ي��Q�MPu�BrU�qY%�$��(HG1��n]����n:��K9�/f�7;�+KBvL�����P����G ̠q�Z��="h���i�d塁#�CȫΡ������u��"4]�����5��٩����X}Ҵa-j�==i ��w�9Vj.��d�1�Cs7[4
.P!�Z7!���!*�]젉�n�Z#&^)W����]�k�h7>*UU�igq���^6-�X!��˖�u�ܩr^�+X׶N�R�TU�wj�PRl�[ܢ�����Wv%�I��E��(��ܫ�X�M��u�.�b��Fj����z��adiD&T����j�Q�ȹ�͠������S������y(�v��Bö}�*I&a��<�F�V/hļ�,^��I��u�Y&���H|
��5�ȷ[�U�dfS����Of�B�x����7E�1�*C��I!�s�V��ԓ݆����Q��sp��k*�QC������ɧS���|�c���N;;Z��;�{r�kkb1�ˬPX����	��_-�Z+�eQ5�K�'��:ܯiۚ0,��i��"T��p�i?�p�;��{��.=���1]�`���X�2]ŧ-�r��F]�aj�B�Чs��$V�
�V`׃)e�-lƤa�w{[`U�~�Ij
��Cv�=&R,��n�mu���5�����kbW����Ո�:q�Bz�ی��x�de�2��㗹�a� 4"��m����{c]��Wv�u�2�����h�OEhwn��m��]6����kZ0�8�R�'(4�"���A�.�L�
�n��f��jh��V��Ӗb81�R񒷔�h]s)�<����c֠���*V1��םW;e�ޯb�*(C������TaZ�V�c�>m��N� U�ٺ�vԙ�Q�IЁ�㛺+��Rݥ6�)��R������+��}�ޚ��bl��ɥ��-#:��V�q��.��X�j-j����X�t�c���t܈�����tdYD��;�cM]ax��@���]z������a���N��r9HN��ֲ��U7+g�s��`�&��!��Q+Fe#��݅�)<� u=+K<��{#���(}+88���d�y��B�Č�B��j�M�[x)9�&�[Vt��5Ԑ�75׹����<�siu-�R,e�ϰ��Z�������Ѻ4���Ώ�����r��ZsjN�(	qM��S�@-m�b��f*ksQ�g2E� 뤟�t_D��S��UkX�:��m�0�mQ,/L�Oi�9Q�>�y��+{��]�y��t�*����֫�(t8�#H�檊�:�ɗ2xM,Ȼm�g	�K�z	U�V���@r�����������@QRܙ뻽��n���� +%L�+��s0m�b�1�]�fR�k6^	�1�+6����aL�o-�m;{u��.j��n�g9�fl�)�m�	�fvT��\W/$�J�8��HYZ�|�;���q*�����y����r�Y�ےZo)�Nf�Q�(�m�o[yx�f��NA �r�x�u��1u�;{*Z�w�(\Y�4�K0j�����I�!so7M5�u��e
fө.�?����3��̽����v�V#�s0���g)��۹:1Xd�Jr�[��IB����!�9ŝ��yk������ִ�IM�z�A�g��xJ��n��Fa�fn�.k�VhM���A�p��knMw`:�Odd�F��ݩ���-F�5�pi�	C�@iN]���V���4ݛ2�S�����*Z�珊	�ې��a����HV��NX�/FSWJ3�9���^w%��V�]���]�a%1n��j�a��gtֶ
�YmZ�M>n[����w�6���4��Ť�2�Z�SDA�6��kF7�)�N���<f�λt�k�r�ʱa�]�qGZ�r]��;�ޝb��]�q�J/��8��&�0�m�W)H���kt,�gm7yk	l
�gy�������m���5��3�ʆ}XkD/B�kt��%�b�t�"BY���0|�y�VB�ZS9�q�v�����</�Q_U��2�7
�]�0h�9%o9��ӌ�)���or�x�'�;�Jt�
%���*mi�V��-4���6�+����]%_rb�$�MiWP�\�&9ݕҥċ�ݮs̡�6v��ih젎2Ӭ��nd���j��LL�MUi�Ţ���th7w�+�}R��L��Ҏ���әmj{"6�v��omPj��4�:⭗ƯGU;�^�9;�R����7	礔����좂��n3n�����g�VO��r��+n[��ɠ��.gٲ��ʄ��?�{$���ɀH�����Z�l`2j{��n�o2���ך ���CVX��gs��Q����+��R�
K�p�k�Z�r'�Ҩ\3�޸�z����,����،�HڻI&^:� K��v�6!;�})d(�KJr���$�&��'�lwJM\5��p�K�k�],)9i���Rm�wP��4pQ����:9&ȮT%�lJ̤�T9�\%͑��=xаp�έ=�Ά�M笛�U��/bi!�elӗ1:������{Ħ�B�X���A�BX)fV�@�T�
�ܦj	��,�%��"���X�?�!��5�nZ�4m�V	o]��#Hr}��ٚԓH&���.��9��Ť��DI! *�v�u@�`׻zl�se��ym�Y�
������㕧�k`r<�U�J��Ӓ�K@�AXD
�`����#�N��n8�$�T����cdE�v�t�����NsY��kiu.]�^�$7X1WaԖ�@Si��6���Z����	�����Uɵ�3y$�C1�[v�I��� ����J����`٬�/(�Hť�R}����-!�"ob�g,�BJ=�B�.�{���+x�C8�$��^��ӽ��n��]� �%�'BV3�iJ>��D,�����ӆ�<Z鱨��{�@e�=���.�f݁rfLV�0�"�`]��,2����ަ��apC���CA
s[�M&G!o���cדd9É�T�v���H�d����J�Ŭ|B�M��y���F�4D����r�0�3����"��գ��R��l5�C2�1t�"�d�cƐ51TG+����y�Bb�͔$� �{Rڊ�~��T2�h/N�4�kԦ�f|�)_�w3/
�AK䀽*R��Fźve8 �ORfFڬb4(��[�1w�y����%2;�v6O3���V���{*�Hq͗8�u�dq�<��=Ά�H���O �j�u F�6���=uvTQ�)�+b����0��� K&�Nl�E�,G4ʓS`�*��s�j�d�k|�NAZ��P�5{$���v�d���ec�	vS�����ԲcY*��43C���*�#%���h�bP�U��M=���,�74Y�	_0��`7/@>h[�[�*&j�&;d*;�.A�P>�R�/e�����0�=TГɗ��n�5�S2X�V�Y8bj@�D�F�ኼ�}��V� �&��������u��.�v����@y�$��6FĎT�<J$:ܱ�D�kw��nݍ`�:R�!����D��s,;�t�&���[��k��K��&���dF�=QGCr]��y�*F�:����d��%�y
6M˨K��*�v)2�LX�x*c%���Z������K�A$�w.kNMˉ�y��cYl*غq��]�kzE֎Nݟur;�n����=�����X֍[C�ݼ��@
b:��MN���nK;�.]�`5�"ӑf^�u4�;�r������si(�܂]��Sz��P@��~�tp���<�u-�ݦú�����x	�A��M<��_�6Ƭ#7���ݥC`
��w�[��Ֆ�Wv'��T�mՃ��-c.��t�[ǽ���q��>]h�c�n	�2:7�,�c��A��u[]�0�uu&Ɔ��nК�Q]��`1���Ԫ��X�a%oeaj���������Bi��oS������97�jc���sZ��o��+�ܯW��!Bݶ8�9b��k�<�Ĝ����w�&�FU�c�ͷ4!y�4��d��:����%gqZ/9�OB��ڃ �T��;m;ӛ�j�Ӻ+Z����`��X�6�����ZC��[2O�G�\����Y��˫u(=n�0���A��cl|�3�r��U��ԕ�7 �(`ʻ{�����f�xJMܣQ!�3^^� 6�YS'+b.����ͤ�&���2�ז,[���� ��-�mS��nG��cb��J�k�%�yr��FZ��4X� %��!Գ�!�աYtPY�{�$�!4з2��I��?P��>i��`X1�x���+%b�--U ������u%]d��}^���s��V�x4]�7���_wu���H�m��@��h�N������}��' (�E�poL%d`�g:��-���r<��	���4�E�p�q1GnR��j�2L=�����A3��8�i��	8��ztdfKJ)3xq�Ú1��Hð���6�E�!��E85X6}����m^��;�jG�F�N�gma�F�@֋��4��B ^ځ�U�ZD�)�V�e3-�u�J�p%��NƁy^S4�x�_:2�d���Q��k�YH�e8�2��LZ2��I%	4R�Nf%8<G,,��e�v��j�.�NE 13g㵉QZ��jL`����ub��P�&��V�8��/]$iiAu�����e+����n�e�<�k-�se4s��l�yK4�5c֍�(8h�ÈŚr�Z��gp������'l����98Cv�E�ӈ"�S���&��췗J�kL`|�����j�Z0�+J���w.�ݸ��h%ʽ6L�KY���dh	�m��'���lĒ��ٓs�����l�u��zC�a4$�V�b���[�:V2�������`��cC7[7���)���CmM�2���Y���[�&�t5]B��[O"�5hFj\� ��/ԕ��ױ��w��ܲ3Ŝڹ�[ۥf�$1����D�,���P�����C� ��=d)��ۻ�9E:�������IB��b@�U*]e�Bjma\��RiZؤ;2�4��`H��[�^�fj
l�kL��ghj�1ƹ�)��Ǆp�٦杉Z2�2�$��J6&^7B�ϴe[̉5e��a����,XL�6���o$�9��gN�F��kǈ���nЃ�F=�8�7gY�p��	8ic5N���G�c0*k#"h��&ճuWeW[]p���]�:y�)�q�����~�-mf7oe�&�YVD?3�F٢X�����Z�<?9 4�̗�J��OH{��k�Y���Ǖw�O�*qu�Q�h�/R�l|h�݉� �@�<$���+��M �X���5i��*�p�a��T$`�}������7+�7Ӌvn;��N@��;��m{��ǵ���^��Q�Иd2�*#��h6U�!�fѥz��8��{�V�Б��Գ�ׯ|���vC1����QZ���Av��m+V�l�e��f.�;[��
��qKZ�nл4 P�f�҃8�A[l��.�*���vx�v�ˊ�+fHi�v��$��K�um�Qψ�Ɇ�yk�f�����vb�f�(%�[����3�cW�ȼ�S�ێ;D[�X{sڷ2ܝ�8��'�V��n�ᱮ^;p<ܝ�k�f��^��OO��W/g{/>pG6�{g�{����ܦ8 �a�c�Ŏzz�ˮ�H,�y&�ܛ.�4C)٭���p��n47��PvS�,C�8���<����1:������v�5qO5�<q�g��u�ؓW�����4�g��HtcZ�hJS�C%1�9�>]�F�����K2���Ց��\�]��q��LlB�9*.�6���R�)ʃ<nl�ŷ#u`Q4��c*�m���kdv{F����+<�q���Ѕ��r���Q�\Ԭ\c vF�Ekm��v��v|U͎��!uk3ںٖW���h�LM�\K��<��=���2JYLAᬽ�]/B(`�v���޻i7km�U�6�tGnT3��m^��n}���0:ۄ�%���l�����;v�v�*VS�\ZO.1�uo[)�vMչ������I��5�z�g	psJ�;v���D�Lܴ��ؙ �#@ƌ��sS!��V]Xlu4�Q$Fʞt�7	^�Dnv[�u�m�7Q[��>N�M�	�T��V.��/r�Ɉ���st�����<����VŜZ��P�[n¼Nb.�7n��Q8�2��9���C�0�k�U�[��A`���z�<�̹P�Wm-�0TWq��ǉ�7��m���x�,r�#��1	DyY��Nm�Y6���N�^<t��+���7KN���F{�n�uq,��w(�K�e��W���y����Vʵ��[���0�eƌv���g�\G�=3��V���G��݂�y�8���t�]9M��2Jm:��M�>kmgg��[�xq��4(�\�K���h�i�c����;�<���\�;�d���ɺ�k��y���
֗m�%ť#�kqa��YqNl�һ����kAX��h۠#m��v�Y�Xp�y��]Fh�]��R�ʲ�뮫ft�R]�[���p�XQ�Rn0�+K���ٽ�Y�ޭt�k��ܢ��p���$��a`��(�8�oe�dΎG;��\�i�
�Ҵ��D��V�nF��B�&x���13i�(�(�F��Gx�Nw��V�2���Y�q�kh�q��p2X Beiq*أXM�r�/.1uٲ4����^�uqwgK	�:`�Y�@���Q�l�c�]��7����!u���r�:�=O'3�]�"�V]
V�pm�+[,��=����5X:�*��:����xW��BE�����l�R��MWW�r�p��0�,�+�����B[���j��'�nVgI��Ƚ��M�Ѩg[%��a�fmZ:�Yj�fmL��Y�$��J،���B���,�cgQ�z�m1����J+`�'=U6��.��M��k��-�
�3!+kp�ڐFÞs�7��c%�;�;uv�a{Gci��HRMCkѧN�	zL'!�#�wZ�l=��N|��t�l>�,���'mIP�ż��1fQ(����ݵ<���|�r�e�JX�u�rK�"�[F����ι�jZ��pk�I)��h!�\��2ْ�/�7��:����guv��7����3g�&{p�v��d��b.;
v\��]��(�h�;g�2Z�=��f]2� ��-�m��Fm���u:�k�gD�J�.�̀��k�F����ДHkL��X39�c��p�1�n��+��;.4�޹2�����v�d�Nk��-�7^7�[��+�K�ڜ )�<ٮV�-�\���u���)(�3@,f�u�˶!S!��\�M�g��n{K�=B�kö�]�ibXj,(]��M�Ƥ�MJ��:[�s�`Qʗ+S7Uch���ZF��e	[v�p���;��y�t�-v:$�p%��l�k*V�q�e���
��̍�`�f�"�	sq��[C������zi6�6�x]ؠݎkp��o9���c�q!�
aϞѵu�X�3.)2���0[T��ecv�	R�<�a:[,�qntqP�I�X�x�=��35��tXgJ�Z�b؅1�b&�#�76��Q�s=�z�y�K�%���� sɹ��=�p����8NОG�6�X�V�{S��=�ov^g9��*��+͏--̙��\�lf����E��+74���a&"�f:�*sǳ��1ܚ*�l0izf�-��4n�A#�}t7���fys�s�
�R���W&y��3��v��7#��v�hVɘ3Ϡ^w\�I��6�tE��2�b�0[����2n�d]z�B��2.tn8�sv痲'/göOL�#�<"ݵj_9ָ۫�����
f��p#W�aJ��y��F�M�M���S�v-GN�$7l&4�Ƕm��ۮb��u��\Dz5z�)�X���`���4]on�0l vp<�*��6�X��j(�I�:��t�`8z�q��jGW ܎o/�qq̾�VsT�y�.n�n(EQ��l�N��E��\K�[���6u'������w������n�ѡ{-tv���]�����im�K��܇m��1΢�� $�V�{i�<l����u�5�ۮ녶�T�.�X�A�J�Ƽy�2�SX���J��m�D������i`�7	Ӛ��3b^5�y���:{�:�91݁s�W�eշoG�1��냃M����Ý]�1�=�b�f�sB<gc�cjۑ��>������baz��9����y�y=m�K�C.�ku�f+�A����RY��q�û3��x�)�&l����u�k;��[�z��)n�<�Q�ި3�JdK�P�C��љ^�^��c���0�b�m)�4JWbB�
�%]��Q5�������g��7���7�K1���{.��6ʬ���6{si<;�#kn:7oe`M����1����x=[�S�^(�s�ru����]/l:w�]�b ���S	��*�l4mW�MnpGKec�c�5�WLK�:�e��x������m�,�l���W�W[�!�==��quxѢ�s����<��!:uȻ����^�7]�z�m�q�5O+��ہ��3&E9�����S]��Z�.���fMK�W����Vh���iq3+3���3lK���5��.1X6�n:���l�O�ΟIL�¹ ��9knq�n0ރ;݅9��^��n�.��k OOe�6�Ɏ�\�jj��Q`�bA���0X�<�nD�:r�����l�.	..�V�<cUJ�-��)�+R�lY����bhM
�v'ƻmA�4�NWX���F7����7m�{�mr�koU:�o�,�t��m:����C�[vyB�!^[r�n�Cl�k{Kh�p�S]s�w�<J6�`��bh�n4��Zˤe@��֎y��.��j\b��u"B��qI@eI�����K,�؄v��#&,G<�wcv�k�����cCi���GZ¥��Q��¸8�/m[���8:w"�!�j.���������+���걮"�=���:�-��x���v��=m)����;n���m�3�ni܏Y��p����}/\���E�ܼ��8{w&[�ٺ��na�.��s��z�r��f��3p���;[J���}����v+�4v�9u�1�M,m�� ��tOF5�q˘�v���9�yIS�Ð\e�8����8:;�P��L�]�+�����b�ll!�oG��[�5�םc���y(�p�����������Xj�u�$W�p3��fޮ�N�GP[+5c�LD�m�����V�6��`����`�a՗$�i�6j���J�0.�8ts`�t��D��6-+B�E�Fuf�[U8�mԷ�Ps�cط)�h���� �u�ӱ[��.�7�z�d��n�6^�x��Ϋ��0�\�0Q����s�OG���{���`N��^J�u�vwt\WY1r+p�Ω*�nn� 2^��` �lj�v*�<��x�9{�tUq��������;���a�qC�5e��Pi���GBit/_y>���'S��5�1çv�8�	��lKj�m[eʚ7g�$z�thӄ�\���tn�lq{�n�H��V�sMs��fq0`Ɠff��]�p�G(�r�K�̎%�s˶u2��iGL�����H9	�BL��׎l-�0�c��n;��;�㞹�&��KA6%MT��%*�\���51ekb����a"�p3���g��K�8��Cێ5�����e'��u��!��rP��8�ey�7t�uv`��q�qȲ����^��l��6�(�c���힣�����N3�N}���z�����`�xt�ll�܍��ܱ��`�I�2m�B�{���ɲ��]�v��#Śr+��5�D�R�&��j�¡ln��d!t�kaXG]v���#�� }�S�xԾ�M���Ӏ���4h�2���Nd�ڐ�7)�aH!C�k�K��W7 ���[GlcT벱y�<m�XL5�آ�ۮ
��<�)��bԠ�"�L�^M��6��{t�n�'@�n�(da6�նYs,�&��k1�l\u�cz��.�pc�3lv}e��&��BP�����ͮ6ݫ�=�+��E������g��/1ڃpsx���S;m�>��q�'q*���y��u�ڤ���xy��kn,t0�����B늣�{[���	H���=/��WRkGCf�����O
��K0�לW<P�@��T����؎W:9��c��hu��k(n�0[n�8�yl���n����kv$x.��ظ v���r�9l�:�@�VV�h�u�N��-#3�B	
���w,[�JX�L-�j��˽���iC>��l �۴�K��[�&���X�c6�F�F$k,p��@q��to���tO�|3C,���ֽB�ı���#-����'m�5����ztI9�[��]� E�^86#��%�JeM"�������(�0�?�"���
"D�&!BQ��_޿w!�C̓�e�r*��Е��`V�2��K�ļ8<t]�Ncl/iݮ��[�Ύ��i�g:	t�M�uQ�Uə��1�q�y�s��EZt ��%���8ج5ef\M,RƤ����m;+���[A�<�=���틕�nݠvTѵ�Y��ǡ����͋��,�XM/*����4��X��<5����,��p�l�Z�&�ˈ�A�)k��Uز���Ջ�\�f��$�H�lG��p0��hCE�}���b������D+ƞ�؂{uk�������ZrX�ل0�pr��W�h#u�aK�A�������Uv5��p��:��{+A����-��e�=E�z�l>�����j<��v��c�ړF���W�.�7n�m�ӛ��ܜ��U�<�bKg��ňu���y�.'cz�uU͜n��q�v�g��K�*�9&�s:R�2�w]-@�E��!d4rW6S	�1���Q�	��{��/;1�S���#�Y탰e.����s�emq��<��77M�"����@��⺎���s�'4�`�d66��ָ�l#�F�is�M"ˡ�\K9��ƆF��a,�ajKY�"��v�����=T\�ӛ9]��ʝs�$��Q���sU�466RB4U��ڧv��/�����cs���N�����w"%��s�i�Z8�v�-H]�M��:}x�R�V�;xMBP{�@8�s[�m�f�0��@�n��CBbZir��;=�T�1�힐kR�۬[��`ݷ�%�!
&���-�6=<�gT)�0�#m)��Skli�ceXwY�v�1uؙzD�И��ʼ�X�gD���0��n6g�;�\Fd��Q��`�a&���-4�[2�X�\�dvV�[�u�M���;���;f�Dг�	��q���^q�}��c����9p��Eʷ9��w7.;m��.�����X�����o\ms�q��݀:�s8��$������]���(m�<qޮ�n؊����w��q�(P
A	%!D�
 �	 Q�%	I% �(�HI I$	BI J!% �(�I �I(����"" Q�)Q��m�Ku���bq��ݡ,��SZ�]�v�;����;V��<'b�S�݅o�u��r� �`G%.�J��V��u���P�j��gg��[s����)��qlc��ctX���{0�n�#V-&tWBq�H�zn5l��.�RFڋ3��v�fB�3�:ϵs��:װV�m��HCk��ZDZA�ܤ5�4W�fshv���{8���rR����܇Qʒstsrs��@:�G)�)^J������l��.aՉ~7z2%R\,���/��A/9P�ژ끼þz�n� ��ɷK�]�?~�w]\al3���S�[�����;͜L��;K ��Z�-�d�՘�-u��mV�o�^Rk�)��I���fj�+��U�(�P�!D�nF��H���B�`������%���KaȴOx�F#a�{� ��R�(�)��'m����iUhw��g�z������:�7+<��Ҟ�GKݜt�a��iPQo�ɕc` ��R�X����Omw�:����Q�w���q���xf-�f�7�%v��Wp�3\����|s��ͪ�u���A��`��W�w7T���"B�b�p�V��U��.�٥
�2�d�fn�d��;�L�X�u�h���8Tn�몣l�j�'Cpp;��n�F��l��{kW���\X�a��D���-�w�W��]�׏��S�U���Q�ǝ��3q�{{�j���b�oT·Mi���T�<:{1�����Z��9��Dp�ڼdݒ���+i
1���_^]�-�ڻ��N�M<�6I8�8Q}J�Q�]F:��/F��ciu�f\c ���0�6R��:S&y�y��1�&E�	�-Vw;�@o���}��OQ���T�eUy�=�ѻ��̊W.����qonN��woz���@��0�v�{�b��y���}��Ey��r�O��>��E]'�YU�}KtSG<M�d�o|ex�V2�}˾���;�i{���7j�p����goFڇ���ʲ@��^MhE��~��:�T>�Y�ԩ��~!͏f{1����s�����#��B	
+��c,mm��9�s�8Z7�i���û3���.v�G:_9��1Pnk�u����G�n窵N(n���C�d� 0M�E��[�t�V�)�F�z����"_
�I8d�7$1HZWƪ/Z7��	y57�ﮍ<�3�ҹ$1j���ʆDQ�=�.��d���_/e�+#1�;Ie�9m�f����&p'�"��=��xl�I�̝K0�)�)J��c;:��X�+���kn§Y�eOy��4=�^�:�x���*��o�^�����h��\�aΜ�b!�y�fUۙ����{�-���F��Km8�_�n���e8��i/UhK;�G���_vR�(Jj'q��g1_���qav���N�=�u��mi������X����)�K��.����ZF��o�����9c��-0ӌ�T�7���*�ξ�d��f:ю��k���'h�b�0���'�-sy��X.��妔�{wEU<|�����j���^f�"�
�7��H�u�n_������,m�U+e�U�.��W:|T��UB���ߨ+��L���l�^�@��Ǡ�@��[��s������:��~�|�R�$E ����m?/La%�r�b��c�����)���a(VW�X�w�U��D�(խ��~W���P~��D���L�d�2с(�y1�Q���/�?�B�wX鞍/�������e���Q�97���5xi��{7Hy��!I��ʒH�x����5}P�'���V+�P�f
�b�pt��.�Ҹ����Zu.�l�én��r�͢�o���"�NZ�y��s`F�/oN�.�
֒�w���3�.:�����i:a�ȝÃE!�Iu�QI$HԒ�&U8\.y��	X��c����z�t���Y�����qiola���$o�6*���C����>�μ��W�ηig���E��\�z��f�2hm��SY�dH��%�V��|{���W�W�c�c��W����@Y�R_+��sv��]!>��>�~����y�;W>���=��X�W37`ct��D�Szq�}�p�e��`�k0+\>��EcӾ����ܩ��A\9��� ՝��H'̹	3zf��Y�S���hV�!bJN�.�[�:i�B?y�I݃⭙!����Y�s����Q��Թ�
J8��>�#j��O���Ӥi�:�7*T����>��!M�Uo���zN��K8&���	��PW�8F^��F��m�\��Qڽ���Y.ܯ����Y�:�u��n�C3}�t���^Rm��t��d�P��M������}��q��Y̴�U�����=F���X;�e�bs]G-���W�P�.�5ZWU�o9�3�� ����6n���$�Њ�X�wjXn��0�9�.ݗ����gqpV�8L'o[x����HD��y�; ����:hc+hd�]n�Z՚8KHE�Ŗ�:�ZЭ�*�6��+�;���vL^i��m��㝹'�]`w��G/a�٣p����o��>*�%[����R��
O�eKH��k���Cc6�bHUY�r~����������=^�֯�ьNX�.-tK^�6�qI\Emi�VS�p2I_��ܳ�\�*�otE��Sw����:�N�Q�My��zd<}tyYާ�0ٚ�ݲ�8�-��lHa7���[zr��r�[�kh<S皕-g �աЀ��٦�� ����(��=Zn�:����"�nD�O�0(܎H]$	D�ԗ��C6�9K�E^��T+��wm���b�Ζ͙�={+�I(�+	:B;���S`�#L"đ��Z�RQ��w����8�����+r���h��U
�rʾ�U5��uoj�ZG��l����<�w�
,ل�������R%<=~/$R�f׎��^Y�*49�^w�d���U�`Vm:�P��a�C{�semi�Ҟ5Y��`�X󃇂�NM�I���+�l�{ez�[���]�a�	�-���Dq##���ݹ�f�H����ʳk��=�=���R��y�|k����v��}�����֘ee�a���<о�y��Շ��$̏�Oj޾X�PкXp�����7P+�+*q<�CL&X��Հ�Æ����:ħJ���#8�usF']�����Uf3y����0������d���:��ܨx��|je�q�b���z�}p��Ulґ�$q>��	���[�t�����d��B�~ï��xƐ��J�h�j9�w7��+1��L#�]��u� s��ؖC�灔�(����쯑h1���w���Yu �;�	��/�#&�j{�����}�;����6���7	��a�G*��C��l,��I���D���z�z0�ew�$ �7XW��׍1�OC�ܞ/����Φ�i;)�����
�Yp�#-J��HUӴ]��gs+vn���ZL-�T��~F�w}��_K����'s�8�,i��+��d�]������%Օr�Z�&���D�2e�(�v#:4�~'C��;����KU��U
�@���9������R����/m�Ͻ��߯m�Vw����l�u=�ۘ�M�M�[�%�,�(���̻tGR���y�yw�)�Ư�O:=L�ט�w4M�c
������(�z2}~�m��Ԫ�ߒ��W��؟2�I�ٕ�2o���=�Xse���]�������r�;sr���=Sњ^�����
N4��M���V�Zg��&�^v%m׭yuU�-UbK=��Z8��f�#W���i���uy=�fuފ&`�PhI��K|��E��k�nXκs{����햾�lN_g��VB{[�F��_{k`��TlC����XB4���Â�@ߏ������;�=un�W��.���s�bU����F���Ҏ�R:u����s��A��88���C�u.q���ł5��ݵQc��VQ�L��5n�yL��A⾴59w�^fr���P��'��>�L�DR�$���=T]����ۮ��%�0@��Ji��dR�U�f�mR�p���B�oMb.]���������z�(�
gS
o?O/�����һŦ�X��ǜ۬�+WJ�`W��^�'�z?��2@���Y��x��Yxd�ƙ�(Jq9��Wx��[��f��7˪�'��c�����n�{�ӻ�q�'t�2^mb�"��K|^��:Ľƺ�\n���};� ����j�w�/y�)Z6�)�iG�y�ђ6Ne��E�n�Y�k�lgh��%+xZ��`�	���-n9�	���AG�mfEhKխ��y���v-nh��*�����	�˳k�?m�b����4��r���{�|wW4�fq�����O!�SW �]Wl��6�������[c5�&��TD��D`J��)"��ն��/��;�����Xݕ��F��d���c���HR�Y7s��ԋ!�N��oy�ʔRluHCN,�RU�Bݰ���)^z�X�A��Y�4Ƶm^/���L�P�{��6d�t�BK˫T9m��ڄ�LpP3��L-c�[�k=���Ǽ�qB��$�AM�j�ݙ�{V����
z]w�S@�B$rG�V�y��&�2����h�|vN���v��%@M��ww��w����F�1Sr�#Ki�����v)f�*�UV�n5�db��R5h��O[/���yJ��o^;7h��ۮ�|,�� �`�d4�y��w������hѫ������΍���ͫ�q�t=�
~	�K_�y+#E�zӯ*�6�FN�+�g2�ߖ]WX6mj-�K�G��bV�t�����K
ue���N<��&!��[@�̰�	��E�٥�E%��+ZK�"cp�ؓY0H.�7(�L<Iu��Ĉ��5ō�x5f�[�4��c�P�%X��^\!Ў��틦}��c]v (�6�G�n���iTl0�SsKU�����Y�r���:��%z��Ƕ]�듯6d���56%l���.蛞y}n�=���e�k~9�z��L�Yi�h\�OY
�����x!m-�ҥ�Ef#�YӘ{��"ݭ�+�!q7i��ҒZgL�,)ժm�ޫ�f�Üx~�M<�4�lۘ����s���{:f��b7b�XN�*�sḮd}V��
���Pr�cuiQ��-;U�o^��Q<7�j�w��\�L�Ƨ.
v|�/{�(#6�Q�S�������2�/jH�b�i�
I�2�q�tN���V������Wd�A��=�	��`6/0�;� ��hJwn�+\�~��M�1�6�H�Đq�=�&��!��^n(�̕��UY/�Z!%4��U{�P�)���,�r��͛p�$�����^X}����^���J���2�������;Y���4�q��r(g;��Uyk	���F),L=� �Y_<8�u�M��p�S�]�GMc,�f�b�-�c(d��V��a�S�������^��C+���R�q-���n�\#N�5S�TЕfF�p�_q�YgU�/�>���,DD�(q.��9�)<���Fv;��zZq���-E7�o������V�@��]�J���8pu�xFΩ����7B�T�I��q��2�t����Ԛ�Ykz�r�9.��ҫKQ�경��U��fڱ�C6�z��d>�P6�Q��8YNG~vX*��j���J����ݨ���-�2�po3�0�]Ŋ����x�l�M��nƱفa�@�Ы����0�˻痫�OSÌ�u�4�����1�P뎃HourRԯCM��k^=��	^�pp�K�p�����do�����K��J��"���b͗ZW�Q�TU�<���Q�:Z](f��G�k��U��am��tx����tމ~���k~�ǋ3K��DS�04V�aұ������k(�l+�lpl�ъ�l�P�����mMͺ���,y��_?���}��j��gSj���<�f�Zh�5�oƽ>���*l[��O߾�a�W[�2���ӧ�2�Y\��_R�R�YR��[������	x��W��5Wh;S��l�E��*���!�hE!i�n|c�0��������4OS�Z�X��U�oN����n3,�9��f���:G�ˋ�K�dr�m�ˀ	v�.]���W�s"HC�]:�e(�Sɰf�1iy��n�H��t�mqtHC �tp^Cȓ�����RU��NS��%`���#��j�/G<���w-ЧyY�C�n�}!e��J�0�x�1e��Z�W�j��:鄨�۝O��-�fU�ヶ�5�W�02�N/c�@��3�U�zs�&T�q�jSjÂ�55e�4�YV����#Y��L���;�cw,r�8sMQ�W�T���[G���s�އv�oG�ѽ�	�^.��Ϲt�y��n_R�	�V�ǅe �V1�|�u_���.��.�_Z5Ӗ<�z��ɵz`����{�kI��
۫��]+U�5w�&�/{���rL��3v�3>�O 
��'7K�-Xt���D�w�w-��[��Ͷ�Йf�bWu�^�\���t];b�k�g�Y��5ٷ�����cqˡ��$<f7��UW9���>�{�jlo!Yb��S/��;\��jΰ����������n� ���7���r��_���>o/p,6h�l�x��Z�N�e)����]{xl\�J6k���G�O;j�d������S�X���J�ԯu�m:�_�:���E-��W��ņ�Z�V�,�����_�5��K���t���v�fk��,UgC�vq��0oM��m;��rs�j�qZ�90Z ީ[˳k�س�A����렏�r,�(أR'�T9]¹��/�lO��Ԅ�ޒ{0g'�V�0@f������B�U� #��f]��0��n�j�FSFF`-D1���va�ފ�xE�qWg��<�P���EYZ�j9��ԑ]0����Iy�e���5���Ur7��l�`M�𑜛ğ.w"�.�p�!r�:w~��V�	�i�ǲ�w�U���߬d�.42���^w�_�?Z?s����9S�pd�^i�V6�͟R�U ���یu�j��)K�Y��1�V[���nF4�R�@���+� #B���Y0�$	�&w^�W���a�4�6ܺ��l��f�gt>�*B�iA�7_[�m]P��-R�t[k
���ER3n�S���Ǭ�T?QJ�z,���v��Ww�:8H1_�U� ��6�H��9ץ0�[��o����ni|�]�㡊����˫g��
���W��N��}}.��e�^�ż�~�~��ߟ��`��ԉ�u��[���&���Q�3v��ƥ�:#>��w�����8�+�vu-�ˢhi0w"%�����쉊�5�6-v�7�oѬ��*\l����k���i�MehZ�VE�XGu�E���[5�{���mA����&�&'�2O��}ێwjM�fVF��'������;�Uzik��h���TR��Ĭոz�-H�E��Ѕ�N���G�Om��2����̲�%b3Yp�e��]3Q������OX�˝��[�A�Zl����x���L����z��'� �c2Q�z�X��.s�l^(Ͼ��~�~FS+�:k߻�k��V��mб�����aQK:rܾ�F�W%�;̥����E�8��VI�N�ۇ��������)8$-g��S,�>���zJ����(&�S�����*R1m	�ځ^뵭e24�FWS����`аE��K����*G>4M�U���GN�N�M�͍i�]
ڢ�3M
�{l�����)b$�xOn�Tb��OF�R���I�M]`R��YJ��{v�Xl`XZo�������^���[*��9ߧ�o�6
!"� �K�b�^p��N���)(�t��.���v�'�:2�A4�oe�N/��4C!ytf����Xs�J剖�d��}
w���(dȃ �ZZ�,��Ԙ�c�%�ۙ(�:pv�6ur����׷�a�;WVw"��:��mq7�^��XG���r�������i�zk��8����\,b�V�Ԗ��5�����i���*c%W�S4�`�Ofl�\n�G��X��yn��A�`�o=9L��\F��H��l�M�:�B��웂
ݻ��j���ɴxW��$�
�*눲���6�̺�E�iiQ��^ݷ;��ϞӮB�-=z�V�D5*B�HV#)�[������B.|�ƾ��0Ix��fhc�i����9�S����t�8�xjm/BbB�BH�>��z|���о�=�|��h�S7Y��ILQ�u���&��aB$H��cݏ��m��$%���R�9FՒ�����ru3����u��h"~���D�z��x�.U��i������7�N"
*�Q�y]�JI��	�[���[�^+5fh�Z͡��ه�O�5B�0��q�+`��h�x�n��&W�T��:�vv���k(�e�eh�R�)P��7��+�/��71U�6S)���s����L����R��F�܍J���{u:W�t-�=5��!,����|�K��J��v+��4���$��Y���U@0���w��&�7۶:M�
^y������>tŷ�P>�<����1�{��gQ�фRO���^�\��b5D���l�����'W�,��V��s܃�X��E]e�34ոM�ˇuRf�b��cq�2w�Mۺ���A�L������j�Ʈ���7[�+o�WZ� 0(�X���5|����¨E�ƴ��ȯ2��XKv}'*��܎(�n"NJ�2GI��bN��U=_@_Sڝ���!3�{������k��Q��GvN���W]�hߌ%y���2��d� (��;@��w�D.K�4.Ucu��aQ��P���heeu�kD�"˶M��y�c{����0�
����$VW�8Pe6a"#��빟Vz�~��[N�������'ʲR�c��x8FE&���;iƼ��UkT͟�p�U]�S�<�Gݮ�*F�!��
��#�a�Yn��;���F	d�v���&�m�ͽf'x\BdM��t��u�q��$:����2�W�U0�G��o��=�7��8wZ4*�L%�r���	�B�y�A$�&2���5�fC�b�s3K�D�ܗ
ƛ�n�m�nC���k>,�K'z��=S┽��%r��ܦy�k׿�{�:��Ц��7L8�U���e5�ש倍��F��;r�5w�Wu��|�Z�y"�uy%��b�χ�u(�ufp�rR��G���۹�U=� 1��3wW!��{���;{:�uސ١з���8�ֽ$������\ۉ��<�\}F RD�IH���PoƼϨ�Ԕ�ބ%o�.~(8�>�|扷�6�Di���D���V9�j��,���c$���$6�_��uz�譡�Z*n�=�J����x���coi�R��9��ɦ)�#X��T��y"]�3��
��G�W[���rr��e��E�$n����v�n���52)+�ƈm�+5j��f �/+v��g�?n�DB<o���z�q���9�~���i��A�����������<
[���a�P"�1�rI�4sL�f�i'QC�I㲤b��-��u7{�JՂ<"��'�4���Q #��է�\ �3DT�w|��޺�t2mu�/��N����>��Mu�����9bӭ���*���gާ�v]�>wl�~��ߏ���:��e�@��V����(�$,��8�}�S�	8ᣰ���cU�G�bOf�7����,h%/s/o!k5�;�^�i֨����n���	u֭�-+��oRӴ8�0���ĕ�k�֍�ȭ������'{��?$4F�M�����W���N�/��^�'K�U\�%7X�w�M�t<7� 廘���>M
�B�$�99/n�<m*�uu����A��`�yC��H��#9��[ٳsc��i��,8鍆�jUJ ��{C������7`���lt�SK��Y�9�V]������*���^=ݞ+nJkH��g	���8.HX4�)���lg�%~�3Uh{͏ӈr�ny���p�U���%��ǎw�����m�\�<���Sv�ѫ��@ے8�RCf�6B݋�ز�g�t�F��U/�[�����4��["�2Z�N���k�
i���8��p$�N<']S�ȸܜ��n[Y6��f��s%���+�C�մ4���ү�5��lT�k��z�B7C�]�!�R1QQ�D�߈����hN�j�_m�V,�[�ˤ�'H�w�Bo��|�C$�������3H�ȥ}�%xr���ܮa������:\�ok0��hyצ�IAC�ec(��=��ꕥg����WN�}Zm��B－{6%&b���ǁ[6���Yq]ea��6�`��°ô�K)�:�����5�ݝ�o�5��� �la�8������K��ޣys4+`@3e$$w=��N�q�:�【��x�)-v�i"�[em��KnN��;��N��m-�k2Q��f֍�ˮ��y���)�;=t�k)'q�X�QGP��eu�9�έ��!K�f��#8[X��s\k�a����M����j���]k���p�yS肻
UCd̛�������.c�0��H�����1e���)z3g�	f>�S���hU,�d�v�]�ڱԚ�~�n�Žٌ�Γ���4�1�!�Ɋ5#�eQ�th�n���*�VyQ�Z���r�MU����3^8�0��'�\mQ��}�k-3gm�L0F�I����!׵��1]Pe�:�'���:��.�}��ʳ�WG�T����u[��DS��r�i�14`0+�������w߷�}��>W^��/|7��@�WN�I�)��S_�)9���������yZ��J�����i4x-����w����?|AUUL�$�ڏ�M�O�i6-e)u�V��zm�S(�x/����Ùһ	v�/h*�>�s�C�ҭ�]FR2F@D������<;;��.�Cغ0����b5̈́c���2g8���Hj)�iƲ�<� ���ߥy�|�r�-.RqS����ٸ�m��p yG�˔H�cD�� h$�OZl��n�i��>9wuW啪�q����.�L�nV�ΛU�y�Շ+������ġ�N=��djI�Wx�P��n�P�>۱��u�Z�>�>�A���a��jpQ�{��wA�[5�q� ����tu��A�����_����E�ҝ�hh=U҆h��B�I�F�]0��]n�D�.�%�e�_��v�ͺu`�e�tܷX�4�*�T�m��v)�R$�	rW��Ǿݡ�F�s���<l��T�W�vl��"�Hv�qxZ6eW�B������ݺ��Tr�R�2����!���9㺥�����L��R��t�] ն��S�vv��;�7w�lu��um�Sr�~"-�b�ݙ���B�%�?c�"	��ظW���]�ȁo���9�%�Ħ�`���u�w�JC+s������������A\�s.��9��-!��#&k�R�%޼k3�����{�U��;p��n&̍A�%PWd�X� f�w�N���q�[�l��N�����[)�X&	}��v��;�=��Y���L�^�w��ie*��hN&�N&�1�c�xe��L����>��9A�*T�J�u�������*-%���P��i�+�oX�`X�u䄭����<J�î�> l��8P"���Y�ef�N��8�1���)_C3m�b�K�p����[�'�=����Ȓ��F���a���T��t��?VH�Xm���g�<Ak�i�%�U��Uy��J}1��m-3�7v��{�y�Έ�<�ʱ�)
N�o�{�߼�S����d��wbh(�r��J7Q�++�Ѭ���6pT�,���l-���]�λ.���m�BkLcf׏ �#m�n瞃j��t����#4�Wͥ��!*3q�wr ���Y�T�+�L��mJ����*��a'�v��+g�e��s��B���kX�w�0��4�JF�)�n��Z�+_?Z���,�ҳ��殆��^Z�"�����7�
���6����~�խՈj����W�Ks[ie��q�#X�c"[uU���.�x^��`��wJi��ۻAq7fxc�U��&恭ҼF4A�/�w^��(H�f�j8�a,w��[����8�ejs������}ӻ���-+�ٳ]Tε�~uV2ic��w�d7���n�k~�z��Ҷ�йѵ��z�!�i���ztT�����f������w�ά���1˔򶞭ٳfJ�<�8=y��r�)��4B宐��R�UsqH�PE���e��z��n]��)�^X�Wm�����Q���I�*��pbh�ID,�}A"(_���E��U/X�S��@�K.eyF�e�r1�$��-���[�<��8v�曮�x�V-�s�����_N�����ǆ�	�M�D �j����\"
�R{3e�ըQ���w���X+3Ӈ�~���k`W)��V�/����wT��is�ea�7 �V�x�&n���tq��ay{�*_[�N�5�_=���n-�Z@K�o�B�D	&�1<[T��:
�!<� Kھ
��������C`�}�JN�h��-��,�ROM�l��Gg4�~�꬙����Ga�!�F�9N��=��k�������#����]���n�@�H����[M_�g�
�=�ߔ�&+8�Kչҍ�-S �� ����	i��/�w��<���ʾ�J���rha���u��:sf�x��"�����"�982*��I�x���A��̓^�AGԥ�9q��4����w8t©e=w�Z��a���yʜe�w\D�K&)#vr6��e�h盘v�V�X�1�lG��w��I4T��+�>w��$�{Ց��B�� a��*�b|M�}�m���ɝ��x6�^r��N�+�������k�R�����w������&3�>�Lx0���fs���.�o	O;5�o{a��of�w%z�d�H�p�g����F&���%RE�!�:��n��l�9ܻk;�k��iv�y8A�y����ymརWL�j�YLAk��o*;0���n�w���K��:��k��t�S7�%"�W��� �����ҽ�٧un+���_��rýy*�O=k2ٯ!"*��+}���
��S�8���9�]��
Mšk�q��>����Y[���Z��3�����H����KX�K�L/q�����:�W����7�x�k>Ɋ�lR�N�(�*���u�˓Pb�;	��{�+[���n���u䵹9���j�u��zMvtmmAXl<���ї�ی�g�NUSS�*��#��&-+"T�ϑ�O%���Rh/,$�?��qL�*��h0NG8�:L*h��i���������b�/ef;�:�7����=��p�Łv�B���b��Z��FzV�6�s���x���=/��m��v��]ՙ�a�c�Ʒjqw�$�;�������pw�B*�2xa��
�Uӵ�v�lu���C����Q{V�}k6�v���y����#�4�Z��9b5��I�5�o�N8F���@�KW��Χ�'|m�y�� 
해��ֶv1-Ut���.M�Í�h�yM������r5� �XJ����!i-u	�w��Π�ܜ�u��l��^bVg�NxF^�����a�����S��=�z�	��G�U�'W���3�����"�7�G�<���Px̉R�S�B�]�n�G�}�ˍ��^�;�\ء��n����n���i��:u]� ��aG{u��e1�{j�x����Wn6��Ǳ�����^n��ߛI�%p���\^ً�I��C��+�f��V�ک�H�JiYz�8�lF� ��,�B� ��� �f�CPc� @�^��qd��2\�us�4	b ��E-#u���nn��b�.�Q�ZV�+iA�N�ս�]�teib�e�����f�nΕ������>�΢����N����=:���8ܞ]`�n�i6�,� �s��������nOM��L���iH��#Ç6
묘�:뮺�t�&Rk�Z�G�IW DoŽ#U�_o���m%��bO	�
�uĹz���5�[$�Y�k>�G[��^�Tv�h��]������z��6��oQ���˦�Tƚ�-��f)J��9��z�9#�vonhMy"�죆[w%y��k���my�]��#,�[��b��L5:���B��N�%�����4|u�$��"9��`��<ʶ� ��v�;�Kh:Ӯ�O/m��v-�� ��b�m��jI.����͓K���a�m��cgD��+�23�Y;hصGCB�L.�K6l�sZi��&�2�X6V	7kN��(�'�mY[<�&iz�ऻl��svM'GG%�r�ݽ�6�wm���c[7vp :n+�����R����=��d��:	S�����(7g۱l�v�̮��E�ha͡vmB�X�>nI*��6o Ƌ���(B���X�Yds�C����S��j6�0�z�6���2p�(�ήS%��u���{�e�G �t�u�G,F�(Մm�4ܕ�$�}NN.j��5nn3�W�����<��sq�����X2�h���$M��W$t�;q
{r���v��j�6�ܝ�
���d��x64نp��@�luuL�*�]B�7Wqٸ�0��9Y\IC0�&E���\cL��H� �r����P+��
��Q�C�b�Ia��p�x�%v��wg�U������M���"�4Jn��q��v��)6�]��c,t)�XJ;ASYh�ٶ3�w!<���c�Ö���Ժ��0F6�5������u�gE?7�	/lX�>*��Z����ղ�����}�:i��S�iwX�}�]�Pf��'S������>yb~�,榺ȭ�O3 ��̨:+s��3�^]���Z?+7�d�^�,�^�߈���ڧW�	�M�AfB����:έ�ieW���d���oT�r�4j�>Y�d��/���[��b_ˇ��JȷsO5�V(� �(�����zz�w���u��g�t�oX����ɮ�>\]��S��Zt\5�J,�z]U�pGq�Eq<Ȫ��M��Z	����_������b����F�X8���5�܃��3f��w1�[^=k����冩t��ߛ������:_���[-�2�^,d�u�K<n�l�v�I��t�	�=q㷆����4~��� -R���ڎ|x#�7&�\����L���o�`J*������O^��5���nu��5C�
�����b���t��:�`�a�Q���c�\l���������nn*��*��^��U��U�u�B������GYP��ڔ�6���l�n%@���M̄}gYMa@5��]�X.��i�ٳ��=~��t=���z�ٜj��|c~>��AzK/������w1V��s����<���~�+�/3�>K�̯r��a\�W���2�.�L�d=���G�f6�+7����z�gD�1�CrH��6~[��֨�Mܣ6��6�u��t��:H*�^��-��{N�U�X����1�IF5Ex�.�wB���^5�baB�R:��*ȵLve�V�LS"�
Gnc�I���^��C/$g�Z�%yu���}�]�a�����������1wrјT��4Kfd"D�[.H�M�������s�ZNk����b]��X�#,��nۺ�g�Y#�W[b��7���Dv��:_ �^^�2��e�՞w����6�(�o��:�>�4�0'��Lq��i��O���C�w�����W	������ݩ�uc��b�M����eҙ�^��ڲS9E��~���z�s9Ly����*��� ��ߋ������S�n���$��F��.ō�
/ur5��ng8;J8��QC9���TY�ڮ�v��<{Ք�</3��p����R�q{.]���=��]����H�Ϧ�z��!�Y��z�C�l�RN}n<ᤡRo��4�e{Fy�!���Ǌx!�����>�2)9�7P�C��I�=[r�����Jө�~���]�qh\\���KO.���ĥ��,��V�ܵ����Y�6r?������K���7��/2?_��}����"�9�;*��[�1��n��Z�b�*����ݞ;�D��E7����b1��ܘR�����YWUM}e����#�4�X�`�r�����~i]Z�XOڭ�U��#�s۽�F�,�Ê���)&�-���{/1�k��W�����\ef�ݠ�	�ok�@��%л�k|�Bg���q=Y�ڂ��ooU	���HB���T`�t}@^�j'Í�5|g��UG�%z����0ʾ�g^F;��w�OK�ٽX߶M���2�0�)H�P9� ,�0�ׯ"����um��,l)�}s��E�<�[��/�]I�勦�7}��P^��>��3�����7)�3�+<)=ыk��F�՚�'f;�2����n�;���a������zm�]/�$�v�~�K��މ�/W�>���� b+���	l^,;!�ψg����͡8�HΎ��rq��=Z���\����l���.�v�&q�)Y�A�a��[�HТ~�8p����8ꙵ�9G`\v�On-���A=�ꗓ&��:b�]f�QGLe?����^o{�ߝa��i8��c�w'y
2�ۓ��r*}�fΚ��
�u<w&x�� �J�����r8�z{.k�a��:�fe�3b~^����_f�k-'�:��lܜ�l���L˗�L]�lՋ�G���ɷc���4d���9C�	k�������ʹ������m���T��ėz0o>�}݃v��/����c������c����o��\zz��e��S�%��H�+�~8�mLck�ϙ��+&��~ǒ_��V��CM�<j �fbI%FlK���ݎ�;]��h}�w�ÛS~}���R����^�<��t;޼_(��:�}��RT�fﲨ�VmǕ�B�V�[+�]hzO_�n|x>iƱ�'�m<	}��c�˷��;P+β/��Fٚs.X��b�Y"mΥ[w{�i�5Os�v=A��@��m�
*��Ke#��)H�KBfh�b�����sU5�Ԙ';Y�8ڋp^�Jb٦�X�u"�1t�`���Y��Ջh�W�N'�fn�fp�����{r-��2v�>�r��������g�v�.ƞ	��Gl�<9�c���:�n��cb�yR��d�ucv�p�1�{{Z9�^.ݓ��;��qr	����:筭X�̧���Wo6�p��n����qv�3hF:f��j�L��T�.͘X*N�����u��Q������7$�ٮ�N��'5�Pg�{hI��>1}[�{��#��wY��{5�ߜM5#��
�6:�$6���d5�﷈����mڣ����z���`�]�4
����t{Ej����(���"�S��������h/y鑁tc0��9��áw���}�z�����]���C�j�k����7S^jw>�+8qO����ޱ���
�:�C)H�MJM�EpI�7��o��0l3���rVQ� �%'�1]O4t��ض�Æ�J��s��}4l�G
=r�[�|H)�>()���.�Mt�X�4�MuV{�:̛��^�,��D�s:DP<Y'��*̺�U��Lmbu\�ݍ�	�R�AH��ٶ��8�2g���M�8��خ4e�xݶ7N���Ԍu�Tp1���q	}�_t��.���g�κy�zq2�g.��r�6z��<�u�<�+Tt��t3��(��@�JH�:0F���-U�����{B��<Un����2�2��O���Q]�;���Av_�{G�׶wWHrL9S��e�y�J����=΀�����W:{[�����Ƃw�
����GO��'M��튊�XkA�=��ToC�7����������n��e�è�
J;~����\R�4�N��rh^�{g�U��=LE��vj� #��1�"���U��e|[�C�!�ޗ�V�һ\B��'�Ηgs�l#��� ��%zw]\D�Q����{���Yވ׬ցG���i�S:[fO��ډ�>�m�O��ۏ���G���^���HgCǁ�q{6�P6�$9wX9��(���[Xn����3��R��w������:�p�і�+s
S2�U���F;Bշ��%�t]l�E�逨f�	5"�Q�2J���tU��	^�"{�޽�p��k�-O+|X"M��5��q����L�*�7��vF�8�)��&Y�#��8�{���<��I�<����9�5W
�GtG�?*�jn�yz�6�/i��ϯ�wNg0S2�MǾѲ9ʩ�FX6��Q(U^������`��&V�WS&��/bxP lv�u<�ϻ��,���*�N��������cHSd�r]3���B�.�t'=��]�甊�گ�N�}xیF�&%���۰�mIi7R)�������s��H�v�Cy�$���X�A����5�u�b)c3�{V�˭�<�4X�9D:v�1e7>_&ܐՐ\��[��������v6���M.�ݪ�Z;:G���U�Y�����ή�w�=���U{��Sv�:�=��P�R��Z\���$�Wk��M*&Y`D�<�Å��u��iM�rl��@J��������?IZ�s�B9����'��(Ns�*����r�֍��]/���bn7�R�Q{�}q�t\� _5�G�il[����O3�/[����Ƭ���)����n���R�ǳ�_��
��Z�m�=���JfV.nT��oK\��w������||<��տ0�j_��$d�U
��Cd��l�I{�YIzZ��B�ù��L�fR����:�l�f�kP�k���`@��Oo`���DN���o���7n��j[-�Ǧ/,h��"�={�Q/��&e/�N��`_=�@_d�6��D�)VD�V�V�44J���BL�ӗ\x�77��R{0�n���]w9��-��r�)�	&�)����G}�6��W:�I�t��m���R�v�^b��{]��#7�'g:���t��dq>���������m�Zy��s+��5�֛n�]�Ad�q���`�[K�r]�J��)4��&�tq��3�\u����r��6Q�]'k~n�mo��S�����h�9LX�M����u�לk=����	���j!�B�N	JGY}q"�]��_�L�L愿3U{U�9{�Ԓf���6�y��JE/"�k�7U6n���[ׄ��#����O��.��k+"d[�^��uU·yׅ�ˡ���
���m���WJ_�?�;�KA�@�i8�E8ݜ,���Y��9���o;���<�q�2�{��F2 ��Z�_<�լ5׀��_Q��q�����E�^����	�55�����e;>C��uE�D�:���z�n(�i���]$�E���gէm^����^Ï.�����f!,���uL��c�P�N"�X6B`����p/�~�'��--v��]����ջQ*ϛ(��I���������-Ө��t�� l�:R؉b��
1F]4Xt�c���%�6ț����3ek��Lp ��V�\��U��h]����5��j[,����l���(�`rl��܋+qۛq���r�dт^�*+��m�ü<�r&�n�ƶwA7��6{M�=�+:{y�)]��yx�=�u��Y�m���ul�t'FvМ����s�����f-����{A��;Y�D4\��#��B-&x�UB��X1�l����5R�����n�߇��]���v,�� 9?3Q��!���:`+k;Cf���z����ʫ�E
1��MH��FV����ht�Y�8�P���D��}�|!�U�.���l�>�>�?T��hEM��ͼ����3ca���=�|���F�����2��mj^B�������hkI�#�Lγ|��U��v�r>c,$٬��>�y���)�p
u偼�{�*s�'m禿Qh0��Ƿ���d�2v��D��"��$�����v;G3�J�;S�1`�I����n9�I� �
�)}�[β۹���;%ͿJ���Yh���vcI�^ޚ[M���P;K�5M�aEI䟋�V�!Z�׉����i��q ��z�K:ۭk±�j�!��J�ݕ���q�]g6�n�
��c���y�4��W�Q����=�xG����������"&'�$���ҶLڰkVl]3c����K�A��YI��E�����3K���zy׶yx�m���F�S�
���E������&&����J�8�]*ɲ��,nK�����z�FJ�Q�׻�k?-��rgv)�1�w�w��R�<�B���W���}v{���E��	�>�)U^�ћ�Q�#n`Q*8���qM'�Ý�2��ʫ�r��p��f���]�ե�@�l]]�Gm1M�8�2���/^Gtz�}��;�ʺ�m���~�=x",����ɶ3˸Es�n;V)N1!u!"y�}L�]�f���h�a�By��S�β�&;��������"-HTq�ڏN/E��f���"�K�V=�3v�_c�ĥ���ܝ�|��It�=��ROT����%�w�~�}!1u���m�-���<�)���+�#v�m��V��ĉF�ܙ�0�!nH�����n���s��fz�{�;^E2��^�;��F�W�u�<ǹ���
��Խc�$HbE�_6��I 9R����s�Yk)*�5G��]������P�wr39*�n�V�zEk���ޘ��Rg��W���M׽���u�.�"d��/�%���v:���Z�5~��+b�}�Be,aeo'<u�4j�����VVш�'�3��ʯ%jRI�����tF�Zr���;�ְ��v��2%/h���p&�9��,����3R_vj%'r�}�8-=����śf�}p�i��m��sL�7_V�\[�d��m7lw+�׻��
�r�=x'�:�1𧺮�/nZ��7�a�k(��5f�Tj���ww�,�*��Y*Py��;C9K�7s���U:��v������vM�AQ�ne]:@�/&� F%;�j#gp�+k	iQ��ۼ�
�Ujڨ6�-���m�K��kN��u���;�������l�����+u���r=n��bP�z�����ޏ>�;�e1MnwJ
��ꎵ��Ԏ���]FABUc�ȓٛ�+ɾ*�m+(Z�9%�D��cB1u��H�����P��3x<�*�8���Zt��׭�"j#p3Iy뎴z�rѕ�ʤ��QN,w�{�FJM2�i����Pe�$��4��L�tc;&Ǿ����v�Kr�j�[�/b��p�������P�|�5��'os1,ݣB���TV����������MMnel�ml�����SKz�=W�ƪ�fּ��X�׏J~$��3s۩# ;4�S2�=�U�{�w�w��Lz&?R�%-��V�@��{�kp�|):��jS�M�|Q�x/�7�f�y��S�K{և�}��S�uL�ݡ{@2��u�c4��{�R���¤\�'`�]�׬XC7ʡ�\nӸ�(h�^Gߗ�K�����uy2��Û�SV=��N��5�����m��u�w�t|� �Z�ko����,�}}��^�p2.��וhzz���77;'���Ɔ��s�t����a���ʞþ��u�S�μ7t��v��$�4M)��U "[�����J9���hy�A0��q�$�)k~=甍�JD���9ME����a;l{=�H��ʱ�P�8BPJ0M���\���j���w������*�>y��u����v����O_@D�����ٹ�;�g"���>�fn�a!���� ���	|�-��D[��2��s=}�����;�<�V�S�Up��Lw_^w����h��8U�Z8��/�]��з��A��/GY]O:>=u�n[N�y;���3L����)ш��f�ԩ��{�zJ>�
�z����Z�ݕ�1�bp��|_�=U��B�^�U��~Bb�����%�$D��Q�#���]^gn������Ү���x׽��dWW5+B4�D���r�!`��6=�&�N��S�:͵;g>�-��d]���-V\�]��R^��f��\y�d��r��[}��WXM�JWX�)��Udȑ��B�2��DI1��]�~�ʸ�{J��in 	ͮ+;�yo��X�z�k�tI���b�K ~ʣ ��C}{�niD�����\���e#�Ц2|ܢ9"�aImn�m0^i4`�!V�l M�hf,.����BQ��Ն�Y��扩�^�~�ѴD�r����M{���U��~��}}G��h�@�l������U�~
�״��p8Ib�rG�VQ��E�� z���8��ZOq�7�}0c���DH.��wcÂ�7M��w�r�aJ�C��ռp�p��=w�O0��R$,(�*D��iۣ�{�,�=nCH�]��Z���ܺ�*=�`��vfl���$ުK�M{9�U�(�J����Jr4b��n{�G7S�*օ�+�׶VZ�r|'xmv�[f����Ճb��~��2����w�<��2T���8�KPA�*��<�����+sg?�:��&�z�F��:�{7)��j��qmo+�y�P&�:�T������!4��T��9���V�e��B�<k_֜Tv�3�${�٣ER؞��a��N�!"Qu�:�#4�d���;6��D�Y{Jگn�jղ�x�V�m�^�&25�j��Wh{�\���+uV�P(��D�e�
�4B�ʲ���ul�j�6�ju�R5��6X�UM�E܈U�/ ��R0эq{&LO�;r��b�M��Rt�MC�e�ͳV��cS-1]xr����/4��.�#�>;ԛ��Vt����d����;t�Q���uu�˥����\{=n��y�sŶO-�Y���[Y�����#���5!0�Z�4�����"B�qxT#���X�1�CQ��*쫿��~f8���T98���z��e�B��!E ������\��H����Ư��uߖ١�K:����}�JUx��!d���Dt�t6X}u���s*v�ڵם�i���W��W����Ҫ���ΩR�����t^���|����;qR-' !��q�^߅�|.S�W3��^q�C},��^vf>ؽѰyW(��%v��!z
�"z��=���V��+s����$�%��`�$ǅ�Dü�n�UKۘf;Y:u�y"u��Y�����q�3sJW؝Y�X�nY�THyM�{�q#�e���ռ���m��9?J��|�W�����v�4�l��9ʕ��4�{��YB���O)v��V�������x��G�}�{jW�_h�c �1�	k��%�pn��	^s�9]-�pm���d�a?O�g����JE߶,�*�6檻��TFb˒񏷝/,��K]o85�ꌶ��[ʗ��]�֥�{c�ݎ%y�6��R�`!FZ2S���6�	sel�j�X4��Oz�D?��slm,O���0�w��hU�ke��K}���-�����|6��v8s�he�0���C+�jni��u��e0g$�����ўז֢sW����w[t�����֍ʘ����:���q[�]�E�$�	�$p珲�O:tw��o��L�z&�oW2i�z�n��PCS�.�|�B�R�+��{+nNɴ*�Ϣ�B�*	����nu��.�ظ����O��*&S�EԱ���׮$��p��!�p�p��%��y�������ן��{Y�s���	�-��|W��,����EA�#�09�� ��б`b{�el���7^�E��ieng9�ܶ&)�I4H�BJ73F�)��F�qHgR�u�`�y�Cq�X.):Rf+��]��V\���m���u�b��߶i@���>�j�P��i<i�ym]� ��H2���:�gl5��<�S��Y/���2~ڒ��V�n���kB�ާs�L�����?;�������G��Lb�޷vN�r�x�,U�<�ݺ�e�8�1��
E$�s�.��*��[#i��U(��_�;��Ѻ��}dY|�>���ܱ��K�j�.ێ���պ7e���ח��5,�tպa"�-�b�il�� �]B��MKƀ��8:Ru�NVa�C~˱D^��5��s�Gb�w߽����Ɇ�����cܭ����m�1-�s�/.�X�a�)݌�a�nW�.J����%үR�5���\4��n��J�}�QM��aFKq�~�VQ;�UY�9�fB$}<3J�h�+Uw��棽fg��/xx
҆*њml��&;���m���}�@�@�����t0�Ԛ�kQ�<��ntȓ����Ɍv�v��5 ��ʶ��v�A
b'׵/PRT=�yY���u{Ԓ�%D���v�
i�ܹ�E����^�e����tF�b���j���"�5nI*vC���:�E�΂eJ�eK�;�� 7�c��!�u�'ʤG[���_Q��p��т4�h��AV���Q3�{Λ�ѵ~XVS�ׂ������
�q/m;���o?{|�1m(jQ����$��e/h��`�bH�NG�1�tF�'�q'��#�}��,��II��殐���4B�Eי�lK٨�I��^*Z���++Nɤ�|�5��y	�]��
n��t�	�����pn���:�V��'Q�y;�Jܷy��#S6����g����m+�,|��E.D�I`���#��Ue��Sƃɽ(Й�T�9�߽����g.z*y�η��B�>`/���:�tyָ(2#�{z���۵٤q���y켧͈��aB-p��.�ű��e�����k�V���S��]�Wj���%�V	��o��s��/*?66��ʳ!�#��Ρ�lohP:e���W�~������S��̐��d�p*6O����䯹w����p㢼>�����<�E�J�|��(U�=�ןX5�(S��4X��`��y��3e?=�o:v;��+�5�mWNt1���V�k��at���<���NJ�wFǂ�]�+(X�}3k�.H�92�:���ʕ�����da�{�Է��]6)�ԫ���ZM4�-�t�d�үl�8�w�U/=�ϫ3�ub�`M����r2܍��_��,��4�mu��!$�e��6�[�~����������� �7��sߥ�Ό;my�m**�1��ar�ɒ��I�~��r�e��ڟ�lr-�|zޝÆ�
=Z�*q�y�p<Բ�k��y��W9>�
�V��ZH��h�bJ&�n(܈���l��k��.���h7,�& �l�Y6�s�=���i�OdA*/F��9��Qه�h��xݝ���\��G/k˜������RlK��9�tԩ,�ȴe.ustV.n��v�;k4s�ҪU��e1Q���67- ��=�qے��� ,k!��Җ��r;)1��qK[�F`��DSTm�������ѳ�c'B�G[�ӞH��x.ρ�8���z���l�%u����3yw]y����:���,Q�H]����D��w�UWq�-��N��f�Ըoz��X�l�N�������	�Y��]��_��g\����G�7���<(n�&z�g6q�dƕ�!����u�^U�����/u�ܯS��H�ꅮ�+��y�QJ{�Q�&_�2̑���yN���r�N�9�R���c7����Uї�_�Ǚ��x�L����ƵV~G�U��n�ʝ�����)��1�eA_��������>s8���/��Hoq�^�^Č�g�	�u�X�+��e��>��o��
�Юđ2B��%$L�f�ؚ1K���,������Î����������n�
�Β��h��7�ZV�ʇ�X��-����AW�^U����!�0�;�n p�
h6IB3S8� l݋Q��p���:�A��]��~����׀�	���,����_]]�槺��^,�{b����IK[�3������;��M�_|\���@Z�R����[�Ne2Gt����վ��^�ާ����� �U��]�Q(W�����qbJ��It:V�=pP�Ҳ�p�7:�Z%Z����:�uq����)������I�#�����4]�+P,�6��:��(�<A�f@��jLk�}s���^�u��Y>0�n2$p�$��ok�o���.�ly�TSǻ��q��j�u���Z�o�}G��r��o�~�<	���l�R��kG�A��EI�fʓ���l��g�+�Kv���]lN���
`�����z�vS;��B |��
Û�_R�`�SD1��-����A'[Βr��#�v1���%����¤P�7�
�U��!'��uf��w&��J�4��v���m�td&oY�c �M�p���g'���N��� Tn��.3�
?�����1՛��1:�=KV��V�Q���:k>Y���
�ˠ�7��m�W:�Gު�W__��AP'�I#�{b\ѦW:�����XS�׎С8ltFm{��w�Sm�j>��V@���}҆�&P?y���[��̓R �`��� *p�����2?a[��|(�zw�#=EE��9F��Η3�'^Rwz�M��4N����\��e��ڇ��0��uK߶��0��.��Z2�g�λ"֌~���Vl�����\�f
�?�v�/ɪ@n�6@��H ����mzC��+}���h�[�ۂ�A�X멪k�U�Q���.�q��`R�I�h6�pSπ�mK����ɹ���q۱�ӊb" QA1�$u��t^J��f^J�l~޽L�u�_���p���xT�m�{�[p�}s�g�y���е�=әކ�/A�[��0�\�H!����]�m�=�xJ,��*�a����������-E1D�{�వ�J���rQ�}�5\���H/;7�,f�������gee\$Y��t�Lu�:��4�q�E�3������Nʪ�G���^�K<|Uq�P�չl�
�d���,�5�Y����p�(9�Xtl��9�������U-stH�dx,aAFL1����,Rg��z���w�UZ��Δ�8ք�%�UOz��R�U�ݺA��1������I��TCG`7Q0�!("J'#�8�����VKՏ|炙sjD�k����͋>E��UL��{�\V�N9݂��cy���T���mY�R��eUm��B��>���pɾ[�i�-�I~��ڇ�1�X���_��Z�1<G�lE���=���َ�M��YS9��DGG����K��&�����ǺQ�8����5��M\�*�Ը���y�ݿ-��i��I[ΰ������ᩜ����T�Jj��<����?�b;��aw��"\#��pO��ӝ�gM7n�g��@P��t������HԆ,����I+���y�R��\d��+��="xoe\��2��-�߅��ؔ�U��,�0?u��!!�G��!�m>�Y�ut�S��iv<E�Kū��2Z��lL��D
˝�(�]c���^>1�|PC�{��p����)B@Df$we&�L���MHn���bӵ�{ϔ:ȫ��4�����в�([����!f�<[���Ƙc�c�`�N��"� y���nĜ�Y&�5�]i���<����S����A���oh�oDx�z�ɽb�>}u��=b���G��?)(@L�)�b�eӡ^����_`�Tu�V�j ���0j�N�v�.�\&����U�p�����;�t��)���h���VmY�`)H˄�1ߪ�z �5_���w]G��\S��uj�׹�B<��x��Zӏ�YΌ�ʽs���Ws;��c�w�I�ģ}��U��GK~ڷ,���7ȑBX��	o׾�Rr�V���Ud!i����R�ӛ����/�;�`��m���/��m��ŵwPVܡa�K���z��J�=B�R��L�W���ʑ�o���X�X�u�����p��^��|�5n���KM]-e'\]􍗶	S��嶫*�ю9��Z!�L��(.�wr�%�jk�Y�eK���x`1T��6{9��:����ye8�	��V��9n-�F��Ď�k�AYf5Ҋ��X}�vNUӶ�J������hR`@D��2����Ժ<�(��څ���:�����{���[A� �B�R�zV���+��F��Iͱ�No�ax�q�j���#���Uѷ^u��v��Ń@Nk^�1������ ʖ�7�͙IcS2�����K"�X��U�ī�\�����Os;���y+f�]���{{�6ƹrl�P�|0R��wh���圬���Ӎ'��pN�I��X(�١��UǮN9�ט��e>�r������6��U��2#l��l���PJѣ}���}��z�V��Ae�i�i��(��v�>#/Y�2�n*9GXF�:�	��qK�����q��]�a._Iq���㊸��쏣�KB��Q��܏n����n�]���{G�u�(�m+�Ii�\ڽR=y؀��������8����� $�v������=\A/i�CB�]���#�a9��U�t��ݓ`d�Wn��[%������v�kB%��	[G�L8�*��ͷY�%e&el�A`@���Q�/�9�
�������v3$�%[D��#�3����oA�4���n�M�!x�]V;[��cu��l�v���]`:�WN @�'�o=��A[k����q�0�TX�6�}lD�g4۵��v6by���s�����#z9��]����.$�u�i���4̻:���*�[��k���:�42����ڃ2U�ư��y�u���ic���#2��٭�|�k��@���r�XNŸѕхfu�&�����%zD$v;,��:���֣U���S��m�h�mt���!�Ƕ<���������g"�����vP����ݖ��M�Þ���O
B6�笽��y�tڵafkrru���A��
��g��@i���j�db�^ρ1��:|s�[W��9��Xs�&�X��n�c�1-R��-i�I���:���ZpY����v�*�hM�i�����lwO�vtk223d���a��i�8�U9�HH�n8�^0M�6��k���X��aR�@��,Z���ї�W����ɹ&0v�r7�y�<Çs���ع��h�2���n0kvݝ5X�k{$�k�ի���n�7n�6���������ϱ�僺e�.a��mM�m6�6n��Jٟ7vu���5�����v�u��ۍ��ZH�f����������]lL� �\��Lb	��SL���5%n��X�؜�n����<��;�{���,	���`�l��4��y�ogdP�!�e�x}�X��]�V��9�
rgq�[��"Z�#4�[n�M�z�=��L�1c��b��[�Iۓ�`ݗ۝��})�͖ޞ��Q���/q@��s��Ĝ]�����+֏a�)��Go;g��n׬9r��u���+R�q�.\�mש�mέ˹�����.ǣ�ͻsvm��q�5Sd���dwJ;'t=h�ű� ��r�է�i'���b	���ٕ��v�n�c�Y�6�v��4.�핱���r�y�lGI�3n�aYE�ʐ�.���4̺\���4e�6�-Y$�#�N�.��UŬ�#4W6��3����j�e،�/ff'n*�����������vܾ����y�pWr<Ju���c��s�֛j[�3V��0 L�	��:.��^Q�x4Q���co:9�U��.�]4\n�fk�v����p�fze*Ulڲ4L�!9q����˽Ͼ��5YP����԰I�t�9�[��=�������>֟}щp��p���}������]�[-0�Ĩ�~��O�J$n�N�ST�:���d)��M��{溜i�����}�y����E��q�Hϯ��������G¢E�s)Y �����rr� /*r��CBT���ӭ�7������j�#�[�B��������6[(�������ą���^�K����-hH�i�QLp���q�m���^�$]Oޟ5�'WZU��E��ɸXE��7��f����/m�&�/�}r��[R���Yf����z�6\��W-�N�����ܥ���Ә?Rd����B"_�w�qKǥ�D)��P�KM�0�{���q�(��);ƕ{=�N`��8)Y�1P�����]oW��V��4J���DX^{cy>{���fl��g�;�O�no�#!M2�R��f}M�ӂ1�	i�-�]y�93W��V(�{����������
���,߫��Ľ�muy�z���,J�vX�|�>��93!{*aQ�_����䆛qD�h���"���m�t�{W���_�Twn��Bz�gg�=F)5�Au��'[�כ����O
�BU��{~�\:.��d*!1g��{�gċHRG��ۅg��}�/y�+�y�>���L|��s�ޘ��t�4��Rdnԫ<����eҪ�N��)��>B�pL�5�[����w1%�o����̩���m^�ے���v�ɇ6��K�U�L��^�����A�f�U���/�2�p�4ݭ�/eL�l�ƫ��k��w�)Z`��}�g�n*�X�R�N4�#V�9[�����������L���s�I}<��bS��%�ɤ��	p�,
�~��}��!W�g���?[�_�}_L���2�M]�;�H5#j'!�t�0���S-��%�]W'C'����|\h��^wm2&Z�
k{�X_��U���1�$�W=���ԿȊ�A���Ou0)\��l.�I=i4.�_������-g2Ĳ� dW��.h���w��T̺%0�Nff�#OG����x�o�A��+�e}s�})$�=��V���E���1aZ�J�y]�����d/s��^����HZe4�o���h��f�Ō����N2�VN�(�s3]
̹��TaOw���-#m���8�y>|��I�T��)IUK!_��tT|�����ݯ���:t�6�!}�m$�]��M�l=�q�.����H�j�Tp�w��0�M��>iQ��$�����W.H/���\��X�m5Z��������J�׺e5Ԭt*�t*&�]1>���f+����GlR�V���T[U�mb8EB�!r\��b�{��;��*�����±p��~���qsyT X`c�`��>�K�=��}w��������r��%����#�0�__vyX�]8&ۛ��^�)�i�����o;�P��k��T�a�<��μ@+4��{�qӇEǻz���[�����	�/}0�W32��nt�U�9�}9�:-
iW��j����H�Y���"�.^Ͷ�#s�\�����޵����(����"�5�2P��g_���9�� ������yl,�[�!n�y�Z��a�s0wL\�X�u8%�<⟻�Z�y^{ִ���>Ѱ.�C���|�U�E\�4�­��N�Z��Ϸ�S�/����)��b��R�B�t22 ��\�)V��3uf�S�?
8�lnm:x�!o�2�,Kޙ�x%|���>	q{eb#+���$'^��tR�R��*�S����e5Gg;��2/q7�Y����կ�����}%ʒȱ_�b�b����9nギa1"�+�V`��.�s��V4�N6ƪ!�E�R���dudժ�B��|Z��i
���F������{�fK2؂�S��/���N�Xx�j���s��
H��dБm{<�7���M��4��p���/�,Z+<U���J��kL��
��\���|4������7�t	c�4�-Ɗ����=����t�Rꪒj`�z��:�7�j�c�2�n<u��]gZ}{3v0�m�B��V$j;��[=��}�u���|���0�t�������EbVZ"�B���Ր�|��H�q�8�V9X��{�w���_�����_�Y����A�����i��}ׇ���Ʌ��]rCd	��%�4Sq%�2����A��l�]���p��oU��{.�r����t�}��}�cJL�MO��ńyw���M��ID�Ww8�����_[K>M�p�W�;_�&.�}����gk~������}��:�M&�n"�rG�6���
H��V- /o�x�QJZ�k�TK������q*4���̥�pZ<qD���<K�9TC�%��E���'�b�g-jB��Ss���ud�}�6�\�%�U7H�}*�B,�������~ԻƘ��ϧY���c�Ʃ	�B��O۞��^��ޕ��ׂ�Y(J��X�9��6�C-tE� _�}��mJ;YZ�Y�蘵Q_�#L9%��R�7w�;t���sW�d}��;d�s0�v¦&����դƺ���ذ������D��XF���ʌ �
HT�ߍ�e�fW�o��.�~��oZY��X2��O罷x #Zu=�B�$R/}�^��&k���|������[gei��H^�
���ws�s���pW�j�EcV{�JZ`�	i�;�h����M�R~�T_��ߪ�{&*��!%�`�H:��M�U����&:���p+� ���c [���9uvFܸ�߹?Y��?x/k�jvdD�P�"{�5\^5�s���tɅb��2+���p�ݔ����M9��3�P۷��=��b�SV}���w��*���<4H��~1aB��G#x��N������VebD[����\#��|��zQ�4�9/�]gՑ��>�{������S?>v:/�Y��u\h�VE
��X�,�,����F�"�We&%�ȱ}��`�:������9zepc�~�	e�8ܾ}��ǘٗ1���'����_?ʝzD�p�,���U���(��h��E�ki8�����"�m{�H�:p\~�K���:G�G��#����l��!X�etTF;qm�����\4]D�nĪ�[�}��}������j����'�xbg�����_H��W�n����0d����8%�Ƨ{1�/cKJ�f&��&��O��Rh�}�}W҈���ZE�[��_R~���;��k���:��l5���X�O߽����pla�v�Ծ:FO��^9��+œ{�_��c�ֺF�iH�+y��'�y�^;���{9ٴ�'ݕ���i��i3^��-�y���zB�"���VLH����1l�ऌ]��0�vh��*�4S�g��p��H��C�t��va�
�9�F@�>7j�ۯ{@���uI�BK���]t��®�R7�M�/���j�ܵ�ҥP){ɾ�):R��QI�������d�]�Wѻs��\��Z^:���,���1v�UN�ƹ��rv�xgp�9��Y�a{��8櫍v���Ǳ!���_Gsh�&A)���a2��`�L'�w(v�Ѕ�=�;n�zC�6�H��\�>��n��:9N��t�v^VCln�N��9����z���^�����d�Gk����J�\ifkf�v��÷gOaHŶ�V#�A�u[zD9��p��q���d���f�����6������
�������뵢��Q�2�ʱ��"�}��,L�'
�9ST}߉�$��h�����/ҫ̍<�>8j�͐`���rmn8d1O�r�1P���ܯ��s�w5-Jt�eU
GUńi ��5Bd~��K��m}��R�g����?4�)�cVY������-`�o�;�æ��E!mkězF!Hy�B�0K�g�k髮�����Ҷ�m�����;ƪ�	:���m9���M sN��%�Ee[L��g���%���ϻ9Eξ��I�4k���|�,_h8TC���G�Lp���� ��H�k�vEd�\֢�$1��ff�����`D��"�=��i�R�	�9�њE6�@�j^�}��<�~�X��{�t�����bֹ�b�r@c�0�ﻖ�Z��
i���`YN��L߾ޗ�-���*ňKs�w;u��+;�;��M��a�Tl������%$kjH]�w��00Q-��?K;�^F�� �ҡ,�O���p�G'H��	�8�������G=;�_����aYb}�VX�o�'�]��\�L��Rdt�!]�����B�8RB�C�i����Y��5��њ�ِ��Iq*��RY�VVۓX�p]Kv�!��h�̪�?������bRH}�V�O�����5:ݸ_oܥ��Ex�S����K�}�őv�˄�Ȕ�~��W��߫�HھX�|#�2(��Tج�}�s��˅*�pUy��t魳����k2�ܳ�,#ʮzcRc���R/��>�+]#��y����u��6��L	y%ܙ.M/�Ι��5`�;���Вؾ�謻 �cLZ�n�QNW0ݕ�aWT����d�r�q��4��V8n��j��%4�w��pKOK�̠����8�k��+<E�&fL��=�9e�g�is�r���rH�
\&��βfjduI��w������K5��/��kdꋳ��ධA�z�L�9��I�Y1���oD�֓(���CO�j�jw�HS�I��G�s��p�B`%�p��|�N��ͮ{f>�,��2�	G±);�O�9NS�J�L�Ĭ�r�F�7^�3j@'.��~�g���~�w�=��ҹv&jֶڰ֤�}9��E�8X���Yn%����\!�O!H�K�Z7����3�<���o�v�y0%��Q�TFz�ߟj�)5S-Rd˚�ZG.se:Ʌ�Y�+�e�Ey�՛ŉI���6%��*��nO~ڐ�w��/��v���%-0�*��y
�߱���B�1�Q=��f���V%���Ȼ�>�]8.��ܥD���iL�����{��6q���bc
ݓ�9;YA�:4ʥe��)���3���rk�=;u�ۆ��c�4)��i
H�����k�������{u���F�Je\��T+�B��r�a��DY
�D�2��m#yO�W��z/�����Y.3�<�)#�M�"� ��.S��E�_}o�T�)˦�S3N֑�=j�B
��V*��ϝ��޵ޯ��+ӛVFiɌ
�м���4q	���$H�s�1 ���ĸ�������L�>����q����ٮO���:t�U5b����v{YPh�`SA�W�:���um���'s,��v~�m.�y�[dy��s"�U�>p}�n�V:֓��~�K��������_��\Fgh8p��J9����d�[J�	�&���&�&I��%���Z����V��I���e,��+�<ʾ�z�~^!Xīg�w� ����)'�*E6���/�;�'=Q�Y�k�4��<D q�����#)�>��$�����^�b�,�}��Z*}��rqn[��]�W;�|�]D��)�����jȢ�����2�[�=U��XY�|!`[JQ��k�����r�}�8*��ͮ��[iŊ�ʓ���#E?k>]�.h�Ъj����3�]��0�X�V)3�����dB�iIB*��9������t�����1Ǽ�kYN0�Z\߫�ir{=!Y�j���,��u-'Y�N�q�Ƥ��\��魤�$w���k&�_�g}ï���1��q���8cY���kR$E���M���$AX����f�7cm4�� �Y���"��w0��qŠ#EK�ߋ�-߸��ZB%�
��go��vqEn�;p����ɠ�yx�-S��s���/�ztTY�4Y�1��q�Zp��s�%��]��)i�U6se�˚�c3nFy��Y亴�Q4�Ȟ�}��-7(v?9�������d�7ߩʱY��wz�z�I	�|j������ �HB��r�,�=!L�_S��~}����+��Y����7�+�"���SN�uHɧUV��8Gݟ�ia��;zR y��,#K9��a���E���_k��ĸ���#պ��Mvju.������4�We�+���D,�_��b�h�_[YN��Ƭ�H��o����EBe�I�o=�^�Ņܱ+>�O�n���w����p짴�Ĭ��%2,_W&&�u����I)!e?��^�}��3x��"��a�|�&��YU�o��T���b��ŝ�{���bTӾ*|閅š��"��`�z�n�ز�o����Y0ԩf�����>s&On�Y�1�1Q��D����g�Y������`�4�,�Z�3�qc#�W��!p_:����/<�TH�$��S;Xx�T��'�D$z��d����e$��;dZ�>����ґ/xK�rm3��Y��H�s\�a'��y�V9S�8�
��z���zO]x���%�nR헂�8,�v�|��dO&-�n������ϻ���x	��|��:G��v���^:.�G[JO����ڎ����Q���U�]q��'�w�՞����w��J��Ⱦ���S�8Bvԝ;Mi�/'�����j	�A�"y�����>����l�dI����Z*�_k����4���Q#�|��&�=$�P�.{R?g��;�W8�-��n8��K#w�������WmIb�K�ƹ�w���y?i~����e�(�ʚw�޸TO�5�5��ZO_�ٿ�pS��{j��R�s��tN�TG�j�՚���d,1���fo�kE�>	�g�Yb	7/���ڢ7Z�"ϳk���>�G��~�XԒ�Tܪ��������iV޾{��_W��Z�\�t�\ ���*����}6�A\�E
|�e�"m�+���.M�F�k8�RE�_ã�߿k����gՙ��k�q���G���)�_qq�� r��GTZ�5�P���d���8*C���p���(�)��_Q7�Ln��#)��O;0�����J�̿����dQc2vR�;�`d)�ן���Z/jv%�R-���g�=�ܕ�bp~�<9z�wZ�}���b]�o��e���ޓ{���#2�_Oib��#g���U2�[d���J��6z�©s=����[N�g�Y1�1��ap�;jWi����0�5�hy5v�vd`���n���/��2y��7�3�t�^�]ڞ��{e�yvKm��Y2l�D�1+�	��[�XQ��B]�L�z�f��;������f��x:t�5�9W�Τ�r�E��w;�T�\�-�i��eMa�
0!1Y��R�E�v������s�Js����G�\�[���]���($t�鍵����x��U>����I�j�3���)�oKR&`��cmċ{�
����;����E��y���ë����;��is����;9����߂�%${�;3��N}�M����']�k��sz���4�����P��uN�a�gn�	Y�]��D�S����~�ۛ����Cv%�C��S��o�wbZG»i��s�4|����^#�I6�D��:X�"=�sV/"8*��?�o��Eg'�Jτ�{��}��r�*ئ�r�~�~����[aM㎖F#ճU5�b�z$ɧ���-����uʛ�.�8���~�������.��9��t@h��K��.e ��>�rw�[�	3y���� �������R7T�jJ�*i��"��]���8�t��ֱ��Z]3'�����$�H��0��#����D����E���8ԉQd'��:d{_o��X'�T��LS�|w�Vl�H�3��^��=�"�tT~�M���oU$HBI��G�i�P�iT��;����Ǒ������S�/�λ�ߔ�l�'�w��O)��J���m�����q��XsϤX��\�ZFV}ɵ�q�	|e8�=����~��/�-�Ԃb�������4cK``�ΥMs�4���5r��u�ӗ:�j��rS�3�O/?���Y��y�T,y?r~�]/rp�~��GX)����w�`��}ia��p�lF�U���
�4�e�'tЦ�g��ڗX�&a�}���u1�YE�K��]�5:���Ը��m�w�����)�2�)�EX�^ϱ�-,Eb�e��[���>V�/�W=�{�>�P��4���œ+�+����h˰��}@;��Lz_p�=Z�ogp����\�4���N�����ޜZh��E&�T�UT�\#>��jEϯ8�*�����g��xM5b�Ͼ�O�� ���6�Չ��6;t���C?z�?��˩Cn�4�,XC��r��RX�_��\��Q[0ȱR	u���ެJK콨V|-���N!�.7
İ�[�p��Ea�J��֞/3��h�N
��UnQ�N?�Թ�d�P����,4��jļY�}~��{��cKL�w������z%�Ք�Q��5��֢9v�p�O[4�d+=�#�;V.�����	��QʝZ|���|��U���\t[�Ӆ쳔0��ߎ�!ȣ-H�Rῃ���Q"Tr�V/�������ib��*,��o�"�7��hQ���{n�{H�?y�#�¢2�8TL������`����r� H(��ݾ�{�_g�b�i�y߭Y
�5��\V��%���ԙ�����;Qv-Y���)�������-`�sм붸�V��#�T�e=����?�n�{���_�2�K滅�O~�-��dJ�}p��}��\#�J"v����K�b�����7�I�:��������J��۱I����._&��tT���2�]���߿}�L: �l�����ύɲ�,�Oo�_]Z�pOo���ߔ�y��$#jaH�;W��	����#��ǐ��������i|tJ��J��򦴂O��<Y���E�;������+e�?�ݟ�7����/o��*+Z�Vj��p�X�`Ĭ�lpĨ��rխ"u��LY
�LUm�W}�8b�|S+>`��~��T��g�eR�<�c�I�}yj�+�&��X�4�Z��(h���\��qL�4�̕�+�����̂t�k7!32��RE��,=�%t�G1e��Y��#��wb�o/�1�Z��Y<Ler��Fы=]�I[�k��v��8�Ь��d�rT���y�:�v&��Uq�twYZ�̩�P�;1@6�M�����|3�oō,�G
f�Ȟ-Ƌ�nкj��Y��b��u��Õ˶L���Z p)�7�s }�r�9�֫nX����&�fUѯ���Y
zi��FʲO��<����$w:Ѹ�0d�fՁO�Ij�uW�/�g�yJS��km�v��CU�ա�N�Td��Un5�+0�n�F]m�?�L�:��m*w?�V�.�8��ux��܊L$_�S�S{GU�$�7�5���c۴�j�BG[���%�����'�U����k+{rW��\tP�Ⱦ�48ɪ�1��5T����kWC���]����\/{<���I�_��T�+=���T��)����tU)j�a���Ude�DА�4͂h����,�+'K�0FK��h�)�[MY؉���^J\��|�^�Ďi"�顸�^��ע����R磴)G�U�:��#V���hH3=��m��YM�T�˛���/Y��Uz�T��*5y%iϮf��9��:��u.���8�s&��kMMu5�R���aQ�Y'aH��d�c��c�)���X�v:�)�^�֫EQ�����y�2����Im)����A�*�I��I�l��;I��H\�޴
ķ�e��zn����yp�>Y��K�����]����#��n�2ғ��/��ZdiOu|�ϭ��瞀�>7���\�U��i��촨�"�b����1[����dP�+t����}�kEt�Z�-���k��i_���]I=9��=X�}���b讞����WN=mY�U�"�l9R�rC`i>_rB�q@��0dQ<���sŮ�X�]���!Yý���~����[*W�4~|ݖW��
͖�}�O��x��􅇸�E�D�'O	o~�pΜ#�)u0�.7�p��MY��j��T��SeH�J!�F����q�*�ܬ�h�77cW1���ɇ۞LE���U!2T4zc�$&m�������E��"ίLY׶����.��;d�f�
e�#=�ߌ�&�W�:���?����	n<v�V�L�G�߾���:&ڳk&�W%�WW�?K�T�jH�0G$���^hp(��Q�C-#e�F������8�/�K��VV{�(]<z\�.q��w��aS�)Q&	�Z�8�R�����9�,��>��a��U��xB>��zy�*�͏������r��ߤR�Q5�j����I����`�m,4g��dU��ͪ#D"$m�>�蕈�>�خ��;��I�eQC�k���ߩ�r}�H]!T�s��E����W����,_VgŠRiL��\��{�R�.ϛj�5R��U�$K�c�,�1+:��)[�P���y|�%�N7o�����p�D�����8.�S�'�Tƕ[���W�R��~�'ު������^;�$�K?)�a�xb�hxߐ+U3�ڵ�NB�:6�o<�R��fF �Z�qC�i�d�MB�T�g�r��"X^�ޛ���ӏ6�ZG-}���l�EQ{׫�o�-oW��v�M.��e߾�ฅ�¡X��CS\�e��W�^ᐏ�0��)0]q��r��5��>l�*�
���D`��ߌ\��e4Ù*�n	j��j�}�>���|����-���sQ�w��*(�VP�`a�j��x��*��M\�H�)Y��:uU���>4|��0_Y��$`�!]};ګWEâ��sBZ��}9�d�&�ʅ$H��
�$S��\p���ϗ,�Zց���E���<.��b�w\P���%�H�k�>(d�J)I-Ժ�[  p����$�(�
j�'����b��y���M��f�}"����ܨ}��܉7�RC���%=羫K�>%�+��|/�}���sG���{���Ts�ZAk������;��n��ը)ܟ��{x��>��Z������p�\�Z)��²�K*n��q.�S"�̻����{W�\!}���Zh�Z+"��iib�����-s_ƒP�nĦ�b(���d��jJ&7#P���,�"� �m�TR�^N��z�b�������E"
�B�b]>���ؓ�ھ4��^zV�^�&L�1��_0����^�~�
ĳo�L��%�]�xZ뙎q��&���Ͼ?��Θ��u��
��,���-R�}ҥ)��OٿS�PU+3�?�YX�pTk��)u+�{��/��M8��UӅe��>㴾\���Fge)��Y
k���h�<pRz�o�J�1Ǿ�W�p���s��M��z���ͫ�?�g��wo�����^���6�>�L����ᕜ>|
	�!�2�*R��6��k�R�^{&�6�Q�9D��Qs5�U&�P5�����G���"z
��A�&(
�����fw]A�*�Wgٕ���J�ݵ�@a3��I�+Ģ�g��Q��K����=�� h��,���okQV\K�i���:1�\x ��YT���4o'o�M���ij𰄣��K��\<�j��؍�H/nz��4�鶍������V5۲u![Z�i�TsK(� �Լ��{k��ۄւѻY�+q-���34�L���'�*ڲH�f�7n��ㅢ���{��x5�B�"��c��w�.%D}�mӿ��te���������{�(�*_�0u���U��#��	}�w�Y�h�50��L�tR�>�m��!�C�����%C˔�J�/�ϋKֻ垏}k���L��8��o�$P���z`��U)2�b����3���(T%���J��|��8b���z�����?^�W}���N���f�cH�,��Qp��|� V0S���/=�\-�
N	j��
Eb�W٪��؜³��dh�c��:��X|i��]��fw0��ZxӄH��oW.4Y�I����l�v�O���멖�2(9��ȱpI�-(~����f�����E���e������B�e�eP���|��Z�7�L��dO��Hз
�s��C�)�8Y.���0�[�5�m����6��8+�"眷�}U+"����9Li�MS$�,uJ�i �F�)�T ��;�-T�!:sƓB�^�v���x�}��-*85��Ump�j�LE��}X��_�[n��y�f�/���7�Ԁ�p��
N�V՚�?��g���&�R�p���IM�^���A�mYw2�x��'c:�ۥc��"ڶ#T��)���d)!Wǯ�㧺�pr������K_]#�Qg��|+���+#��.�h���u[�{���}��u�9�/x�[�,\=��^G�(�6�-�%f����4ʔ�:C�5*8Gϲ��t܍y��Rq���ξ<g�#W_�}F�5�������+�0��*��ח��i�V�Si+x���)��(r��`U��S8��q��\�T�'�9��󝴽 ��x�t�{�����W�&G��H:,֦{���R�����:���k�^0���߹��Tp_�k��3}R�!-ş1[:���O!,`�q��\��_�k���茹狕�i�Q�ʩ����!��JH]�r�4X/�7�w�}�
��b�{<y�G˨��s%xY��:^�G��k��H�q�wϾ�M��I�|G]K�-�^?�;�b@ �e0��<�_�"�p�}�rs�k㎚)7���uމt�Q\��/[L�wss�D���8#�{XF�{��>�#�o�+�����VWfw:��[û��z�#�Y�v���Bί4󾿏\��H�GV��4KFGN鍰,�"nR�_{~/D�v�����e
�e{�<��O�WT����n����Q)"�G�m��%_��p�q�X��~6����p�����k�{��YY0�v��*�]�1�~C�����M`}C:͂X7����]qme96�N�B���.K���l�-uFr��Cc�$uĪ~�F
����[b�˟���e�ǅ��B�+,^���pļg*�X��pH�﷦%�D]���O�zw�Bf�b
#[��7���׭�	Yb�Q̛3����T4Lʤ���U��E҄	Q�x*�X%��~���8+���O�����(K��
�#;��k�+���m*,�*�-/�q�n,ǒ��������ɵ5Ncu�/���g*�����sа����:��u>�ȪI���%���8��V+�Zi���"rg���Vĺ/���zB竔��M|ػ7�.��ׅ�i���%̞1��]D�a~7J���2lO�յK�;��'Qb�ɕF��v�$=K�m+O�RN ��[�Ҩ:�� �)I)Y���:�s�>M���n8I�J�äabVƨ���n��Ri�s-ƢJ!w��*�ꀨsCtT��-!H�A&�93����W�Vgp��4�5��n�[�Ĳ��n�̿���:�=#Ｒ�B��5�K���������&(�E&⟴�����HW��ub�~׿>��X����/�k��R�EU9t��J��r�Qd+>"��|��_M����ċ�jȲ=-P����~����}��z�|*8G��2��5�,=�������Դ��U��!P����g����*��Y��U�����>�'�H�]��l���e��:뮱g@P��X����[��[J�ذ&lK�`*hD�̬Ţle�B��+GE�2m���&�-�L��T����ib�Z�������$���0�����Y��+��`SI�[�P��ϋ���7�YS�k���L\��G����}8�4]!�27�P���z��.&��)�n��RȬl�<��T{�|"�Ty��@��j{���ڞ�r��%�O��n+����%B���pb��������t_/���c�p�U�W�.�k_H����G4��L\0�����i�����z������wbtT.�#L0��9�p�]4TCo��/�M�Ϧ�JV���
�odS�O�����'-�f��W$}[J��+o�X���O��ԭ^Z���,B/;�J�G��|�L��0�eF�ɤf����N�.��m�;t�:s�v�ׄc��|�&��pb�ɏ�jե��ix�i�MJ�
�ji}�V�g'�lK�K��%�IVy]��O묥3�^�Z��cܿ�&��p��l��v�������֍@̩-�9Ҩ:*ݔI�V�]z~KV�ۃ<}�%����ǫ��N8|.�����fcKO�/����,�#a@�����#�}�^����(��H�#=?e�}3E�8������.��|K��tK�z,��_�ӽ}��ܴ@��--I`����E��>3_7y�JH�ӄtW�ߪ���8 �}�9��`�E��߹j�]���T��bT �%�hF�y5��#0Q�\�C��8�H�[�iaJJ�ML�W�|�^�)e��E��̝��rO}����:"o�{"��3\*7����:\)�*:/M)V1)!]{�:B���<��T�~?~;ȶ��DӅ|�ܴ��K��j�Fy��|�?��1��h����ά�֞^uI�JE���=��\.�'~2e�O�"�1�N\��p�	i$y
��%c�+�Ľ3U�_.��HT�'���Z�3\!$�s���ғ�,Ԥ���/�ɩ�d�)�nk�M&�#�x��웈��o�b�(^��B�	a�w����r��$.��}�V�\�V�.
�J���͐��>-W�4��}]iY�X`����9t*��ܩ����:1��'�]���說�����,�g8��ZGɯN�p�:�(eKR ��8�f�B��J��c�>-pA�)7���4��^�l��o����=?��f���F�J�=Mg�l��T��&��/�o�a�o\:��M��0ǯ{�Q�d�B�w����%~��܎�i��w/���+Pf�ȞL�H�����YB�i|M4��&���m����ac��>�A
�=Or�Q�}׵pڬ����F�%є]�}�*�l:� 0�6�s���`�j�(b��,=DvZm��D�9���K�Af(��0�I�H�ff�G��n�����l�M�&��E�$���์�
䳺���,OLR�	���a�A+��[%�xjgmҁr�e��Fs��CO��v��<�ˋ
�����\ĳ)E8t���#�ٮ6�g�ۑ�iK��[��6�nfX��K:��Eije�bX�:v	��䢶tx��'C�g��\gUv��f���1"�)�����+����F���p��og[�m��]���T�ɑ>�D��%�ϭ��b�h�U��՘%�Qc,�DX��"���\h�����rV��4���'��H�_y���p�x��q��`�/sܩ�ZG ����}�c��"��;�~Ѽ��n~��$+���Vi�N�~�k�G��-��3��V��s]���Y�J�kN�����g>��gk�L�{R� �,�;9�k�F�+ٛ���L��w�|h�}�uy����"&W%W&EN��pL�쯵��.�0]#ﯽWq���4��kuȬ�k��{�~Dx�8N�kYl���*#&I��?qZ\��HTb���d��h����6�̱N�vו�[K��1�����:�-ʚeU4��H%�-��ϖKߧ�ۚk�UmN:��Ζł�J�����}�ϋ���.3�Y-��,�_�p��
M�*�����׹�,�>�a�q�����;�:%�}�Y���G��tɗC�U33FD��~*���L,�P���b�XY�*7*k�j}��G���P�=j�Rs��;�/�{��J>!�u���RZQb-�������D��K1ċ-�;�ZG��ﻹq�;s����(�*e��jU)�y�z�㝌��c&�[�nۈ�NP��y�	��A-�e�h����k��:KֹqN����}6��L
�L_k��>�ip�
�Hh\�m�1¢����&���f̓�\"Hv5Bf��O8�r˘�A�8TFjj�F��������A��S�N�=�����>�/VB��c��uN�[����ϫA��g�:@��j'3��v�	����R�����p��9��6�Œ'XUm��'����ٴ��٦�[�S�e�\���d.�S��31��s�-Q��B�"�q��tG~��r���OVw�}I`�F	i��vm��_����w��Y����}^TxVG�Wd���}����ۖP�8�;�R�l�O\ۄ������/�߲�����N\��>߽�XGL�=��,\�OU[�����?'�)�+�NZL�uW�����
��.UK$@��T�\|t�:�X�Y+,��>\
��L�ɒ�˪1�:I�8�ƴ������dϾ�>�|���|xu����t]0XG�խW
D	��ݛ�xY�[��L� $���+��S����iX�u-�Y(߽}�H_s}�3��ry�ޢ�~�TG�}Y:���a�:�Pg|�^w|�u|�w[#g�}ǔW�7�.�,VF,k�X�b�{�fw�:]�w��+��1��5d+j�w�jļ�g��=��d=Ʌ6���ךZ�qz�4XB��jV�Sϵ�9�N�/#����佃�mkj����hp�U��3�sp�֦�V�\��j��.�A��#H�~0�c�Ǜ�,��ۼV���N,��!Y�9ى���Y
��#$V-��)	}_gť��]�דM*4��v�������7�-I�.[A����r�m��7B�SRӢ��%g [�Y���e�ϱd|-�Y�_ٵ�o�߅�P����A��?�;�ギ5$Q
I3�n�#3ﾫK�����JW�U������V�>���~���i2�ߤ�������^�6ö��3QwQӧ����X���_��TF�H��Nq��by�������SO�����!���,�n\iʢ��Ѕ�x���PW�Nf���
��U�����L���^�����5!ֈB�w�)�'�5�+��s���4
+4X�Qb]'�����8B�.�)�'��[.ݤg8�&�Rʠ����3EG�0�r����,;:����_{�p�ƙh�����#�f��p���P��q5BZX�.���u\xäpUnH��J�iK��{ӟz�\���[�\(K�vb�$sP���_o�\��a��*8���ׅ���˲H�Q�zRæ���狅���|���L
6Dꟻz�^�y��_�Eu8�Y<�,�).�T���0�O�}�LZ%}xi�<�ݛ��8B�[0��k;��4������FX6et��yC��ջk7��2l20���M�K�1q��ۭs��e�2�J�2�B�8TBd��>߾v������6Xcj�Sj������W35�-�ܫ��֔�B{^���X_������[����e��.%$|^�������髨�\/sf���vQ��d��}ϵȻ��`����N���ZD�B�bdO��K���n���d��בGr�T�B���.�f/+�U�#6f�I��^f|�.�>���V/�5����rg~�x��\���ܾ[=�->��cq٧��鄪�K
�e:�a`���$�n��{�%�~���4N\��3p��B��#���mJ���Xڱ|<��♾�j�q�.\|7y��i�8Q&�)����+���1aâh�Z���ן�Ƞ�8��rG`3�i��/�M��h�+O�}�p���cn����r��%��*8M���W��B~p��k�S����w����C��.����^�bY�!��_es�z��1��M�l!L�7�u���Ts���km߮�����!W�)c��^U�B#Vn�p*��Ɵ�7@��oV����x��ίߝ�/Ϛ�DXYݍ��N�7����~m4����i�.q�xT%@p�(J~�<����NSR2U�����wU����z�׾����ʨX*~R�K�����ٴ�����b��$K�s4��va�u�}�ޑ"�Q�՜���z���ܹ},a�@MA��6��e�Di먦��qPO<��HW�V��kF-�ͯϡp�Ƙ��xT*m+*��.>||��+>|ډ�o�+~̛K�%$N)�T/�(��ig����W4�Jm�~�/u�iYD|Y��c�=;2&.(J���D.���
��Jd��:��a���֑"�	E��<s\��pZ���r7=}��t5�_SL�w����TP��!I��|���Ľ��pŁ���\�X���uZ�.t@�\�|�5W���4��xVE���Ȫ�ʥI�����i2D����B�$���-&h�s1V�*�ֶ�O�ў돳~��.V}��3E�>F}�c�{�p���2_1ZR`�,V{�����.N}ϫ8�4Ä*���d��U��>�*���\�S52�7���ݮ_���i�]�t�c�\�����j��_�h�8*���%z�D�Cmm�1�8%���M�x�Vs���+'��˿�M�p�^�;T)0���Q	��o�NJS#u.���3T�|+4�u��
��P���ݾ�p�+"Dȓ�SM�+�"�O��ڝ>�=��M������g�4kJ���ϋ]�HT_9)X�O��,���gGmi޵(R;p�?�˛�T�uG�Y��y�BF����(�B��2i*^��үf;H�Zn��Q�H}=�l�[H�CUw���\྆��*�*�z��e ��ͺ�e3�>��]s]C����|r,�weK���_v���zw�)�ƶӺ#���wW&�0-]^�� B_D�J3��q�b����	�(`��f藩���cXP9\��͆��[R�G���=��LR�� G��h6��mi���ES{ò:���P��)wL�0��m7�_۽+��'#n��,5.�*��=��H���YalI��!�ף"t�\˘��^��(��.��SJ�ٯ`�R�E�Fn���
ѕCԪ�KӔ��f�}[L�;���MA]jc�]E=�iPS<�=�I�ґ�^Pֺ&xé���/�U3<d��{��K�TT�̬�:n�x����b�tdL![�H^��]�n�NN*�ĽZr�(n_Rڛ�� ������z�_]���q��8l};�8`q%�z �nJYΚ�mw��ج q:�ˣ�P�o�[�5A�ԕ��_h��.���I�^�(����K��-��\;Z�C�N��\�UzK"R���Y�n�����mǟk�&�hJ�p'�b�E*u�{P�XX�B�mQ��$����6�N�[k����Q�p`��br6�\�&g_��|omi�����t}���d�{V6����s4T�p��vĢ�.�]35oF:�����׼��%8U�yg%�ڛ�RWܰu��S�_Ε�aa����)��u��"� �t�n�xb��k-gS���N�:Ƈ�:l�*��B�]�mV�h�Pp�5 j���F�[%X�jr�1*Q��n�ܻx�q�'�#D�V�y�����=6�W:��ru�g������P:�vڀ�Sƍ���.���l����J�S.���j+�r�cm�,��l�U�ōۜ{��KnNS�&�Ū}�:�G��"�x��4��]���w;i���k�N�,�&^���Y�B]cu=� /�<:6�cQu�]K.UBړ�8t�F�[͈nj�K5 ��q���v�](9n�:��J��z��M�T[�9���棎z��۩�9��2� ��6we{v�1�nz6H��)[�m��:'t��0��Qչ�62>*���d�=��t��>�2@�ب�K�s��m��m�Q�W�x������C�D&����Χ�;˃���jn��� �v�3\<�Z����ٖ�n�*�ɘ;��0c���9M�N+�Gf��������Ӹ�ڠ7t�t ��1����g8���SV�6�7����S��5�dyE��c�Ǝ62� �LKuѶ��,^(�)e�o&������3�qnYe��v�7j�ag����;Q�xU�cu<��1��}��p�m͢�y����3a�4�L�j�t"��=�%�m��ێ24����l{N�t\��m�{l,i �r]g^�>il;Ƴ�]�a��&Z����z�kW�}KĮŸbu�����B	���+n^(�Fl0��1.RM��d#�b�T��l�]6�2c2���m��:��h6�N=�Z0�RX �aԠ�1�aM�J8�R�I��Nk�R�[j{v񃐤z�K��g�C:�@���g�-�[����^^v��w$�A���Oc6�Z��r����c���2՞�t���i����}�=E����֔v+�)�sv�,FG�ȼQ[�*˘�V$�d�M��6�c����=�m��	�	��p�Ǉ�-����
��m��7B�d�۩ˋb�ONt]n3�<�^�tfMDgz=z�.�i8M�al�ܖN�Ԡݷ�6�m;��w�Ҭ�Se�2�6�Sq�e�ڶ�{S^($P��(p��u�6�V�X�yv��Vs[����/m��\���&e�HMm�!�iP5��t=,���	�m�h��(�j�nY׆�q&W�.���mݠ�ny��OB]b�0�.�)s���' �p��dՇ�d�th�Juwf݆i��L�-�9;�����ز���5Ń|���ҳ��:1�J�Ϝ�5Z��
��F�n8Vav8��r��9���Oʎ;�}g�����B�Q�Q?}:B���Z��<+8b֕�s�#i�����\�JL���g�	�E�	�RIb輏�sU� �7�y���d.Rp�TF����aO�b�tm����3S���ٕ���\�����}��!��i��q)DAa��q���� ߼���N��Mߛ��.XO�b��[3�y�R����]���\�?�z�}���;��p\�Pʻ��k�e�C����z��6g��h�H#��)#��c��~	�{����^RN��i�E7��곁�-��p2��LX2��R�!wx�d^��tTڒX�[s��+���t纈�Φ�\64�*[����Q������V,�߷�k=��^���;��@�D�TM)�����nmX��k��-AV-��B�_k���o��%J���
#;��gN��oQZP�v%����f�oe�.�v����^�]}�y{����ڶ��GPo�5ކι\�Ѯ��+.�a0�IaD�TW�����>��<c�~���յܰí}�xz��V%�=��D���f�8��~�o��+wv�׈��ES��xծ�l��\�{%C�ьy�}�g>�y�}�e�����o�l��>p�#�2�����<B$u�{�#��p��BY>P*��ƎG��c=�]{�f��3l���"`.��\���^�r�W��7%V:��>��.a�0yj��i�T�a���l�DE~)�;����%H�Q�"J��.N��Gu��f�ڣ��'w]���d��4�\^a�*>b/Qo{b�̧:eW��ib���z^��O�qu�(�s��P��he`̥����e�h�aW���!cZ���f*�RN�^������z�_UʪG�fQ�a�5����X��cB�{؅���v>Ѫ���R�u�ƹޕՆ�����n�;��1#n;�+h�BvMWC�g۵u�+�H���"VwuC����mi�����y|$�wF������ iƂN"q`��:�ٞ˼�c�r�5�ז�Ąz�	���ٚ�Q̖Ih{��i�����&)�tR��D�V�}�o�D�3��]���ŧm�z�����̀7��@�ů��g{�j��nCՙ�㐰Ӯ�F��08�pȠ����Un������r���^}��*�iz]4�_Jn����ct�J�w�mw��߼}_�=[6��u�;��yUƚ]:Y��ʗ�.���Av!W+9���N�$h��]���\��z�ǽw��`�w'rx���e��a�V��-���AM������
���X-�
���fК.�`��L����g�Q����;�������u�.�hNgr�B瑎]�v�����չ���%u�/���r�)�{]5m��w��b7;J���wf�~f؏�ٯ���+��v���l���$��g[�'Hy�z��e�P˵�G���7%?
��&Ql�%�q��$v����5���6f$|��a"���Ͳy�>,4=��
yCx�xlM��)�Ъ���h&�ƣl�	f�7N`M���S���޿y�'v��&����<PR=}���ݙ��b1�B�uS2Nɽ�"�|D�}J,�XU�WV_]�Nʻ�г�fmf��ԎV��E���Ƽ�Սr��C-��y�A���c`�\�CI�2�bb�tL����%�.U�#�tY��ף)q�ʻp��	�
�+C�����e2*o�Z��Nu�SX��ʼ)��8���V�$Q��������6Đ�݂a��*��"�f:SSb��LK�-��(�Oz|^��?|w��e(Vz]zYڱ������O]׍l,���7��nU��fgv -�q�nI�^]�+��y�=c�������ܱ[�̤s�H�\���cOK껗-?��}�ﹾ��q�j����.&�v�ۺ�Q��K1��*��yR�Pt�Qm�2��4Y�/�W������:�[^VqՍ�M�������m���1v��v�Y���}�n���L�h+Q�_{u��n�e��Џו���q�F1�GP��}�^��^+�+����8ξ���y�˒�HLd���P{Ә���u;�bTK�W�#��u�^�Ɖ˛�c�?�yV�4���F����;7��?{)�"���0����;�gB��2ZGd�FOn
#��0�8v<�����u��%�nh����۞/'��r-�Y/�Y&]vM�2*g��Q͐��Ћ���gQn��n1\��j*��<��������nm���4�Mј�Mے׈�$q�i�l�b6��Kj�\G�4�#b��&	�m��[�qKv�ݒ5��Y�(=��v����e�5�J\�c���]�f�+���ظ���������O����$��8���(n��YKnx��,�t2�`�S[�`���ὣ�r�����"�(q��[^_����-L%�v���?�6���up���u:�z���w��T��?�<��+��Gs�v��U#�|��*2�J3*AUS�ٛb�̣ז0w"�#~�y���g��+$纆�%F,1�w����t��X����>u�G~u짎�J�ц����✺���zz$�WAx�ʡ5F;ޯWJK��R��y�q��j��R�l��<��W���+��s+��/M��K���Q��۞ז�+Ƽ���ֳfS���$X�;��/#W^���������y�y,��7��pgL.B��ጉw���UN�O�;:��/vL��.G��g_��;؝N{��8��0�Eٙ�۾�͠me�:��YV���*����b<2+K��[����;3�b����`]��t-	f��jX�f�az�n�ovx����WE,�ף�Z|���I�֌K��p�W˱����B�SȚ��t}�&��L!�G&f[p�̌��J�����{%[y��G�z��4�r���E^v�M���̀��lu�]4�7��p���f�W9Jh�XT_ǟ�J�3�O>�<M�&���q���F���Z�X٬�;7�	���^�O=���=Ƿ���k�kTG�A����U����l��j����O��}��Ʋf�g~����E(�[����}�Wߋ:����P�V]�"a:�\�@�hC��k�����QY�ޯ,]~����ގF�yUWn�]�|��!~��� l�I��QI��s�J��
�%�����	^f۫u��ۋ�Z	ݡ�n���Q�Wp��˛ِ�ऴ��
��YT��ןt��k�%-�p��u�3A��*�c�+K���8U�m�]�5�K���Fm�
FH�����
�s��=�	�>�vi���C�5��
�J���p�(W�{����`�������q��2��{]P�U>�fd򓣫ƺ��>N�K���%/cO�O9�ٳs>Ǐ�V�����Q����R3"e0d �#�	yя��43ܰ��$�r����>Zc�)j�Z����=ҭf��oU�|�p�֑����b�t1�l��`�Z�ƨ1�}u�˫�ʬ�C\/W���>�uLM�|�;�bpZP�;�^�ba%�(*u��]A�������5�[��E��OjZ�����R��K�����c/⅞w��^�\j�1�eL(Ms_i�i2a,����n�uN�r��UҺnhj7;�Y�sƹ�����4�5Vk�r�ǖyk�CM�_����[�ג���l�Snf�E�vs� AvpŶ�3*H�C,�^kM]�T�pV*��RE�j��b�����Wm]OM��v���YB -|��v��͚��o1UV�7x�|�k%:��^m2�L@�p��� |ڛ�,+��C!�~��q�Y�=�;��M��fjH�D� ��u8�M[~�3�L�q��L�e4�/i��\��ؽ��2N�����0`�nS�y��Ox[ZY��mo\�$UQ�^Їp�8PC *8���:2�>>H�T匏u�_�{O��ݬEW����0�|/��JnE*J��-2�Ջ(�����D^����r�f��U�h�׽;�4HSY���֊�1�[A�i���͙����Y�y��lSM�p���{گ�|�;��!�7ɍ���¶S���F-c̫�����'����[r�ڂ����<_�=R�g��a6/)�c?��I�i��g�2� 5�5���bm�c�q�		aq��qߵ�dE_����{U�����Y��G�X�!���^,����&�X�o�����c��<o�(�r��8:�I¤�F�I8ϯM���>��afN���j� ��xu�j�H��^<ӌ!=�Om��ʹ�/{Y���:��ҫuVS���8���A�b����2�{\B�9�L=聂vwu��g��?9]���do[{��gRv��)z��P�����6���L�uK��Ӯ����G�r��H=�ۗ��`'��B��/LS8��(��'|P>�y�yC7EL�����̧q��N;���ә�|�kV����X˩�
�w���R��~�ǉ�����f끣|=�%VF<U���9��w6�I�нZ(@�������ާ�Yn�Y헙p9 �z�	K�-�#�K(��wN�RÇ"���I�kA0�M��v�nU��OWa7�I����j֑cչs��Sε����T����@�P��7!�4A�x�n#�֬6��riAmZ�m�(vi�٩s��^Qâ�ۚ4��7">�=]�J)�^c��a��WZD5�9��Ǖ4��L)��}�Yy��#�z*zɻu@��q�[<�6��֞���u�c�WN���а���pɳ(8%�[�X��U۶t��p�ڭ��8���#дk�n3�x97�v����5֯��`s{�z��FV��>����#��n5�ϒ���A֘�*V ��?]����(��l��$��o��ߟ�Ǘ��.��Ou����{j�,�8p9<����k�$6�u��,I�|��:��w�h$M��PS���b�����<�<��י���-��Q/`#\�k2�;�!�r�k+�������$uŽ�`�p"c���0�ϋ��5��D����.�'�}v��"J���a�J���P]VΎ>��Ώ�_���m2Q
���S��zٺ_=�{%M��jY|��-�)��+���ʬ��VFblB�ѝ�lb��'5<��V�]����<h��7D��e���w,�k�u'��E�uںw<�:�byl ��+�T�P���_Hj�~��(>�jM�P�ӟ^�ȗ��SKq0x�:x����O�9�teG����!��]<՛�}k�����T!�1��b�]`�NX2�����	�^ѹ�g��q�8Kִ�"��C{pL�V��F����*e*M�6uni�w����[�&���3�z��%.�th��݊�vv��:�Ӿm8��)����[��%/Vn)�tT�늦z����eqX�zS�H���k3����:��=]X�O<i�_a�L±b7u�:�|�����ןk]������uj�J�):��F͵q��hy4hǓe�kS�P�@_Ay@n����m�b��Yar���xO[��nqh���Z�9����O�J�y�IfT�|������vVf�[����:���,��_-�K���\F��ָ�n��g�ېCDau%���8�k'�0ѐ8��ԩF�/��Vߺ��s��h�����=!w�Dl#޻����]�gMb�zlG~���en:�iG	�	m8�
@���w;9T/��ڎ�a���z���q�25Dk�+�zt��og����u���o���ï�ڼ�xs=�PA#�C-�M���u����c]�K<�)nt$����f��Gv����z�"ʽԭyg�����M9OfZ�*W�[T6�f��+0�ZN)Vսj��1f�[�q��?h��}}@�j���f��v��wk@vZ���{%Ĝ�f�1Mv�}����+�7go�Ið��G�"�إ�jP���ٙ���,���v
�ƥv��g3�� S���/��od����k���-9F� )Yǚn�2qk���G����-P۞�K��W���c}����-�>Ԟ�"ש�H�3���U���y�]:Y�;o��:6�B6uډ_^�*�Cv{�wo�a����6\��������u<q�r�;�[�w��������ĸ��W	��؍�Uʧ9NŃs#����w�0u��)�����\^jJݢШ�Y]�gʷe�ʐ*���c�~uM�����������F[0c�ݎ��agg��v�3���Ż�z*�{u�%[��E�����p�ڧt�<~��:`��	XpЕk�ڶ:�/�͝��e�^���b[j��R>�>0j�`B�^g[�06�]�9��Z�ne�y�l�}���d�7��oa�<r%c���{���I�ʃt�o��Y|�+�n�EB����9+�Z6�&C�(�]]����;�w�'u��Ը���b�Ǫ�jj�ĩ��/mf����8��ah0j[���bC6f�Ap�9������Bͬ7x�gLZ�-�w�D��Uzy�w�m�����H�:��ó���B�Q�$�;��R�}�F%pl���M�[u�"���n�]�c��'�=�Ro<19�����܂~8h�[�|{s�����NP����m,�rfe6��켫��Osĉq몾�=�
וչ�{}����l6����x��u���ږ��s^��ʰ0
8Q�����i��/��]r7�*�KIɡ
Ky�zӸ������bN��{U�zػꥶx���σ㲶�	�j�e���ys���3�uu������64n[s��I\��81��h��ާGUr�r����I���s�;�e����]
j��bX9ll}#�󦵨{hj��r$ą���ݱ��d�gw��ze瓧ov�.�ܔ��XUE.�sΩ�}���Žu�ej�9�fX]��mӺ8�f���F5$��&��#����i|�+��|õE/nI*���eb�:K����
�g�v�x3n{/��T�=�\�)�Ɋ"T@ێ���z�ɻ��ε7��H&�:�Ll�^�5��F��oa�k��������|�	�q�����Xt�/��9%{f��oL��YH���2��B�a�f�8�h$�ˊh�S/��U��|��sz�ڎ*��t�u����6�NT���uw���W�[�j�"b}�9Gv�J�c%U��Y�zIJ���ц��j/{��d|���>�y�����m�b]�����\u��;vu��˞�O,`���?��z�b̺�4�k%E\����:`���+����������O��Wy�I�ڼ�=x�Xt��{�7��z}�;�x������{���Kw/��x:��m���]��T3�:��k���W��q&sX�����:���h�V,���.�g^�NHq��h�܇k�:&���_�镙���[��R쪁�4�k�v#okX���"�R������~�п_{{�|�SL�6T�F�]����=�{�3;��"��Zv���9�6{��2��:	n�j�����V��{l+�L5|2_G	��R6���r���=ݾ�N�ؽ��LL���B^��[j��3:��E:�H��&n:�L���̔1"*Bn�"@�����*�6��*�����
�i����}��P�d\��0��1�Ag���,7���唧_IE�~v�qy�?Z��Bƃ6�gE�{%�ڻe�8�%ڵe
��o8�v�n����,Z�ML�:��3XgL6�5���ZR֪�D�6�i�3Mu�tl���k��lv��c�q7n<�9⽧{sl�׎���=�[�vK���j}r=gz��0�`\��V�0t��[���yv�����@n;[C�vs�i�	�>3<��')掷��5�3���,��\�r��y���Em��s�C��l���NVQ2b�B�-��~�UWP~�ߞ��	y�uW�M���g;���{x�OӅb\S�ؘ��os�j��٣Wa
��_�h��]���3��7M�ƨe�?EA�u�ȇ��)i-/s�\t�o�OVr���Ǔ=�k�Wx"�w~�	3	��3a<��=�[����1x%�����+{�򍇶Nr��ڭ�嚵�n�m:�����1]���Ύ�kV�N����1����ۥ�}�w��b�ZD��U�B�]{u�՛�]��8���-Vp��7�֭��������͛J�]�n�����J����!VGU�|�����W�w^���B����w�U⏯cYS��Uڅ'��v��i�����K��,NT�*a�т��a֩2��iy�n��Rݖ��ō���چ�wt[^:�����*�c�=}�P�6�9�:e�O{�ό��A�>��;����{��4��(�F�o+I���7(K��t�Y���,�N�����Gr��G�5�=|�l����:�5�h�	�+.^QH����M�d>����=�
�kV5[�?W��a@�`�gG�x������m�Yg�C_��G���#	�6�C��tث'{G����h({�^��[����'�](��R�{���g߷`�XEn�z'��~�}%p����&_�s�)��	I�潬o#|����o���xk��*�II�*;�bNn��%0q�' z��0�RFS&I"�����qU'cz��S�'�������5��M�~��8k����,N�']�<�
nՖ����̹��I������V�l�-��n����ts�QH1�"햙�U���Q�����	#��WQ�1*������un��)#u�����U�T�]��^�cp7EHJp�/3o6�9X*�Tn�9{	�Wu}�|&y�KS��@z�X	�N5������LB�+�*dγ�q$E�
F"�[�����:Ҿ�=��hp�\��G&*ѡ���oJQ��vn^�B-�x��"�ۣeM��[���}�b���ݾą+�ڽ�Wbo�n����w[7�zC��]ȓZg�ې�}|���A������M8�i%M�!����Z��n�7�o$����׻�N�m�|���ެ7@��Wl�ח�WS~�WyY�.f"i�ڛ�}��Y*!}#�I�uI_u��]�器b�<����Z+�e2�t����Fuη��;�v��������w����Z�]
SCr�r2�Ji�I�ٔ��q��F��qmc��!�]��UґׄQl) �H�1�-�7=��:q���s�]�Pn|����G��$��Ynh��_g_b]�҃Ҏ�@�NE��!�(V7}��������g ��*���dM���xx/84�U�e�֣>�hobWES|����zJᙆ�ډ��R$c����Zq�W;�^z6�����W��j�/z�����Ŕ�����讙KP�>��jK꒚��w�Hb���)�#R<&�\4��w��7����|�Ɯ���mޜ[������������T�MV�e^��0�|�w3�H*������e|]�z���Q���}�����t��aU5y$6��d�۪���+k}�pRCޗ�R�'�c?�&ʑ*Ѻ8=��e9���=�@��r��Qs3{̊��ݬ�g�G��к	{řո�N!d8�5��W`�ajnw%��46�e��MbYi��e�sAG[�F٣p���}]���u�Zg�0��դs�tL�ɥ���d޻*�_b�e\o?�*Ii��-��r���6�]O=ڰ,�۩�wKm�+�~��v�P�Զ%��f�=<�눫�mx?i�̈��'2���{�z�޿}�u"���
���è���w'=r��><�w���?>�u��I3�t=����[�+��H�Q�|�B
	�R!�.���X�u=[���Բ#�f�oL򼉝�HU�&��h�A}���z��o�� �F>��=��T�{<ϒ��T���+��x{-6�)��r��Y0XfV��jWqz��ɓ�*��V'���'�,򼸦'+*��[R��³bUG�h=7:mi�������g�!�5���wQZA�si��]�:�N�ÙD��o��>m�K\�ܤT�� �u���-�zxP�f�F�`�kV�)�.@D0�̛X�X�!��1[1��Z�ZѶ�6�&ږ1�J�.ܫkJ.�4H�tU�t��u�z%�QM��IH���mR岬�q�+	a�U��``��36��aܖ�u�c2�M��e��R�u��.v��[��<s�K�Y܁ӷ� ��؊�8E��͐��l�X�Y�����ږ6�ܚg8��*�t��bB�� �ژM�`������������l���zV�Ω^k9z����zM��-�k�rCϞTn�mx�g�W\�)�<w�I��������R�UtN�E�|�O��Q�����1���0�W��nz�ݹ���vi�< u���Ҹ�+�zMцGn��9\{!b����n�<���Զ�!�m����d���
�#Og�Y}v+΅Hy��P7�;=t�r�p�d՟�xיS�oV��`�q}��s��U��R�vw����c݃u4��}�LZ�����2��E��1)He�m6��_K~e�{�mUvӿW���['�,��5��� 邟X�;X�S4z������gS��M4�:[uY��nΨ$�˹vy��mQr�-�m��JX�2�462Y>rF�N?f��s-�*�����]x�4�m��X��P�=���=+i�_*�f]���7|v"-��A2��y7�o��6��n�{����l��1�����QU�Ǩ�n�3uW��5�3�
�h*=�S�s"vq
��4�U�'���۫���!a,���E{��#M{r�R���yZ�6�]�s�n�V|lug5&��>�EP�v"rE�s	���'�F�N<��fP��+W�Y�͘��2��e�Cc����q�1�MkI0\��mϳ3���5�ru��
�J��^o�l�'�a��U��*TG��;/�^��v�,�V��i|c�R9��"e�T�v�Ӑ�%o�Snkj#uF������.U�[�*D��/�2�e��ט����|{�2}c�-��W$gU�+��+//\r����i-��%q*����$`��,l5N#�i�����Ϩ�̌�#w:�7�O@��_k��;t��{7����~�Ҍ�x1�h7�{�OHp�_h����d�[�\���P����Q�R�����#3Չ��ESo�{�]+�N�v��Y[�XwS≐bd�$1'�%!�uﯫJ=���va���sUN=:x�u��u^�pQ�7+j\F�Y�L�単(��M*�2��3��ef��r��]Իv�:�Q :a�FR^4�x��+|�6�}c������g�%^�������"SM�]��a�#(9������u0�7�}��J���/[//J�M�_�PtGAV���La�]y���d�(�9�Zy�QL8BӉ�V��0�>��R�{�r�,SeiF����F{�ђ ��u���  ��X�>�m�U��M�!L��ut:w�cAmf���]�,5k���Qۄ˲�-��a �&��Y���k��?nJn��X�^������r�'Q(G?���z��s�Bxe�
��ay�LU��9���nFā��~���=��H|=X(p7�T�����dXn�}/�Შ\��s�_�a�l��
�:��Q�\�zK�U�-[�$S�H���]^�����	7���*/�v_�Z8xl��2����9���s..͔���+�5Rs�=eD�i@Z��5�ux/.L��C�2��P�زf����\�v
pU(�cH�x���o#�^�n{9��0�k"v�	�8���Y�ަ�I�d�l^�u䰵d�>��u�S41|l}�k,�A�I��I���垹��i�{m��� ��"xA�����|n�(�n׮nza�ZN�����QD3��ϡ�� Ng����nݜW�� <w�y+���!a��;XL]#��\쬷h�e�g>8tv��O�<�\3m�`�f"�r��>g��c�}�T�zR wI���ϲ��o��u�9�e��;
e2�j�E�$h_�z��X��bFLm�d�ߏ4�y-ۮF����a���ӈK7V2��nv슟b��{N{EEx˝�ݎ/�PֶA�}٩1��j�y=M�/�{�ϲS��a:g�}q\U�u��R���,̘���n��M�}��Svo��؏z�t���������AGy]�p�4�^]��j�y��I5�{w����N�b���t��$i���O��>~���7���Idm8dQ�vz��mAU;��נluӏ��1�d�}q��u.k���Tm0�>�7]*����e��MSG�� ]~��f:���Y�Z��]��n�l*�B��4]�qn(�7[r���U`��G[�����A/�$�}���O7ʼ.��E��-(����w��K����T��k�zbh��EW�
_�HZÞ�%�@�^!���ޝ��)t��2��#�\jP삍]2�Em�i����ևI��I��
3�ˁj}�����˙��������_wgu��
��z��w�����(#���s$5k���������bWv���w­tXa�y[�U,������gL�|�*KL]�š�`ߴ��Ҝ˭l����Y1΍����!���\/�k�V��ַ&���哊̈�*�X��F:R>�M���	b�6�	#��4��w5�3m��-����0�[j��B����pZڽ�sh �^��JW�M����y�e��<�.�i�B*Ш��b�_nB3@[�@�zw}�0�_j�es�8�X�`��U&ʽQ���мw�-:���f�e��`U՗��<;�'ku���t��r�*b(֞�w�]&�³&m�f��"WwKlW�P��本�.�o2\�@q�6oNߵ��t��t�����C�d�/�4�����1���6�u�r�$V�Ǫ��v��mp�/5���9[�v�Q��So�������jC���M��d������ 4�Y
,3����X/��,.��pnRo���9�JGx��yR��39�*Й��q�o�����hLg`�HxS�}��.��6QQ����:�mz����<�Ko4sI��Ҥ��S(Ó�Zx^.�w%��9�ml��I�=�^�Z�"�{KE�<��q�9�iZ���9�����ղ��x���N�{�:�v�S��sػ\d����^�ih7㋭��@sƳѭ˫��1��gQt�dG�]�G&�2l�Av!�r�̹v�A#ʲ}^��郙�ׁ��]��z	�5�vv�7�|mp���1eT�����i���\&98 u�]��,e�&c���uW��i7D�0���a`�f6�M@;y�ѣ��xK!vy�n�FC���'p��;�R�� nY��Dج���`m���Olt��헛m���*v>����{@�Q�JI�rM3�f�c���� ٱ���"�E�Ft�a�n{x�J�]Ֆ1�Ҽ-m�\S�su�h)Š5��a�^�e�i�;i��C�Z�,K��T�Qbd�u��;/Q�,���ɢ1r;)�lr[c8o\;p�9��Y��&��=^�|�;um�taH9lA�ݎ����ڶ{lr[��m��V���z����uN�c-E�m..�u��6�0�Ћ�jR&�J#��%�{�N��d�&�YY]c�V��9E"񚲝ZŮ9L�:�٦}B��i�+q����{O��n�MmLĶf�c�6!2$d���tV�ޤ.::��ԏ���[�`c%c�%V5����^Y�e��e�R^�����':��֪A��[	e,�[qRY�FU[��um"�FK,0�mλ:=-�v�\ύ�>���9��	��)�;og�B�p(��d$��ءsy�b�w	j#:s���&Z��3UQ���r=�1��^v��ŕ�Z�댼�q�p$̠:��G`�[��D�LׂvNu��0t��M�x|�5��g�]�q��zw8������αU�x�9��Q��6�+mZM�Z�=�M�sς=L{�c���<�V��8�6�u�^,kvm2���C�v@��lj1��Ɋ����q<�X8��tL������)�n�9l�c���a헣�F��e�a��&k����ⲛ<oOr!�8Y�X��k�v�w7K��,<m��3`�z�룦b^	r�\.l#J2hYs��[M[[j�e��8�&`7n�<a��[:6�s�S�6;�q�@72�.��cc���띲�����]����p��/c�� ��;�����Bm�B��hB�ETv�eJ͚+]�iP(�-�pˍw����[�=}�ćО��I*q�Z��{�.9�Ib���w��ѽ��22�W���S��K�ęJ��ޢ�7��_P�>�Yw�0��2[��">u}�$u�W��x��>6��M�x
n��ڻ_���t=@#��k�F�"���܃�_�4T�@�ߣ������jx��7zh�T��i���ԡ����W�>򩪬9tn.v.%�*Q�����Y+=��q�O�Y{�
��!=���4{������*_����W�h��']�ÓE�:}���Q��3-UN�wЃ�{��Kin��.az#�iʻG�����Y�@s���b���Vׯg3ḷe_8t4뭧�oZi���^.���V�Yf�������[�E��jD���%+h���.�` ��%ȐE%�U�&��4;�4x[���U�UU蜛Ξ�;kC�彻��Pt�h��Q�s
��)��z��(�N2�JC�F��+��$`��:+|���f;�cw{#�0=C�:�	��8:+�	p��e;��Wk�e��[��H��=���dp�v���1��YCt佽1���X�Y��c��T���|���
��7��n�W�;~�tK�J29�	��U>c/�μ3��k��[�ɇ�|�g��;Z5���/][����ժD������7��*$�Ϡr9�~�+L�����ڬ�ޥ��W��~?x�c��DֿUB:�W�D�6�N����~k���]��ևh��p9
a4������Ǉ��F��-�o��(�N��=�i?Pɹ�N�ʼe�G�uR�4P�7�m��u"���j�X˩+sMʘ�o��$;o3Ҷ��K�,5�a��Q�,Ā�ӭ:�գ�x�ۦ+���7�"����7���>��'��,���S��&Ȁ�WT!��B}n��𲈷�=V=�N=����f�)0��w�Vf�Yiܰ�ϑ4��8����ߵ������5z�)1"��2I$�?X�{�&��e�bs�i��O^92[�dpqg�g���(���b/
��fZ�ћ�����d[�<ˋ��T��%���Vnѫh��1�du���f�r���%�ʵ��XӜ4-��*8�6���f�s7�!�&oO�{�:���kY�hP�}=;c�^|��fw^����s�],\�YG���w���7�^���Bc�u�'ޑ��eV:h�u-wg�8�&@��,��[h�o;tOUU.༩����u��yKU!���F��@�]�W�����{<��xڳ��<�~�Nk ⺌-���-���1C+�A�y�z�
���z�=����i����.Z��ү�[�]?Kky3�o��׋��50�rP�)��p���c*l���6���$(�4drG��o[���������}=�H� ��$;4��܎��{s��N��o'{�m���[2Vs}��;✬���U��J(�s�T���*B��38�Z�VS�����&�՟n��ʧcս�&òc�iI���l+�������K.�`�p��6�����/�xIK{ǲ�r"�p��<)�ޗj�����֚�EHX��U�N��ؼR�t�P��͌9*0io�ƆoML���<:�P�a��*sF�ޭ>w��_�*Tn�������#<>�=�r$� �͠�<�J���:��L�~,��w�=l@����;����{����z��g������K�}�+6f��}����Qzl-¤p�p�� ��\4#Xԥմ�{i	TŽ��s���&���c9[fX̸MU�'ߵ���J.r�;w�gΧbW������Lt�}���Uܧ�s��;g�D�b�u� �ψsk�b)��E"m4�~�J��Wa&�m�}���3:��J��;R׵�{g^m�5*;��X��uQ�[�zj��[�7����n�+�t��l(IG
	yg+{w�>�91ѓk��5;!ެ�Mf�z�z!;>s�~��z�ufd3�`�>�,D�$E�`m_}��DMf��B�l SX��W\x�mw(��z��}��F�K��=ʧe5��m>0�V�����rH�N6�[��)�%%t�8�Ȫ��]������蔾��Qd'L׷��,J{�{/��B�-��!�+y��ⓜ`�Y��?w���eZjչ�0��}�8cU��h�	?�Q�H'�ʻ1q뻺��t���+��n����W�����i��<Iv:�s!�1iƣ����.i���0\bō���qכY�J����8H��P0�i�3�F�u�s�/@OcN$Z�n=���{=�N��<n}�z��u[��[<=��Z��s�v��$����M�a]:幱����̓�u��6��A���ǤM����ss�֫ZF;`a���Qcs.�����p܍©�s	P�.�o/��<�',�\�nL������6fo�2��-S0��Qُ�O�ϝu���{�����yٌ��b�Q9���m���#�6t�;�w�����p�D,�Q��1	dѢA�ԳP�x���Z
�������]絅4Y��!��>�:���n�u��m>����x�v~۹�(	L��G#����ɝ~�'Ow�;Ki�}JԶ#�#w�he`c�LсvoA��mN6w����67��]cҤRH#�͂p�I�q���un��#�;��l��d�&���El}c:�R�WF�k����t�Ż7�q�0f[Y�/N�'C�w~b��z�ȁ1i��]{q�r���U�����]z�z�U���w��Y��F&v���^PUs��Uu����0�`ʿ[Ъ��b�#�DB
4-}���<FY�ݽs�b�w��ڌ�5��1��)�����Z�)�쳹��O�,���������ެ�tc꾞^�S�C[c��&^T4�v{��=vlzyV�`q��SnIE#tA� �Bc�8}r��h��wϪf���&k=�w�xs����C�kiN۲�2>4;���q��;�K�tu�F�E7/-�B��\�9΍��8��ПS�`�����1���}�ۧ���������Z_/[�����*7�,7�+��{���_��R��޾k�BY��SR#$���ȅ�/.�����?2`��G۷ǯ+{�V;��
Գ�躐j��;V�������f�:���i�F�A�É��8�Y���&Us�¯�.�q�!痙�f�q��욝!��;4=�c�R��~�����u�7�s܃k;��Ef�H�z�����T���d��a8�I!�}��DOsf���~X+V�"9�=�56ә�����n�O/K�*]�t�������5݊W\��Ɣ$*v8M�Z�]�VP�p�:�pH�;&'-���q��)�r\�u�<6���Uvn�)�;l�@���V�,���9�֐e�kv��;j�R���~ۻ�'{)n�_�7U�Gއ�o�|�ڞ���,��U�DӐ�ɐq�{��s��t-o<�+	�$��(kO�5�g���^��@�k���!�W)��g�k�W�aY�y�
/v����;�w���b.�pCS{;�q���%_��[�@�BE�Q���>�`�h+Q��³]�/�z�nQˊ����/��uwi�2��M�Yr@�zPYqmc,V� ��;���I.U�|q��<��}��&!ƶ��/	U��
�����Y�}�E��~w}n������r���X;\ �����
qT�ؗ����C�e9����6`�{��_g�}�0���C��[2� �i��U���ybʮꩋ?K$uDZ@���f�XC#	�\�w圿N�&��<�B�������FgQ�T��۰�*yQ�n���b�&�o�
�G�G7{Һ��}����]�[sF��Y�ʘ%�a.�6�&&��kL��G68���Ym�l�6��p�G���]3�I�^JsgJ��j~��W�?�CɌ�E��f��X�ӧ��ň@nx����6¯w�3tl���S�}����b�j7y<�{o�:`�]����T�.[��@'�Q���#���� Y�<�Yh���ܢ��E�;���Uci�{�(&!�g�[�מ4�f{�C0	M	RC�R���z�|qe��GƱ
#��U���y��cY�y��Z|�v꫕�d?7Xh��?`M|;�������ٌ�]�C/�^n���K�ѻ����Z|�Q�1W�Э�[��u���B�\�U�7�0t𾢂�V�u�yӹ"��.��id����^��e���Mi�6✱�J�LW-�����n�h;�qY[5 e�~}~�S�,���T�~w�W׳1�8{��(ڐ��NItoCR9��vh_Q�.���/"���?O0��v�aD�ܧ�g�]��D�B[�eUsT�C�{C��%֝�q=�߿o/H�����c5��h�5;Zv�n�Sr�S����1�1ʃ��j1� fH]v��)mu��)R����ՅU�����H��v3���0ѻ���گ5�q��ro��wqZ��?g�%|�P$c�H���(<A�Kw��ȭܮu�r�Q����IN��;�=o��	�p�����k�I�Y�['`b_R�;]
{c�X\2�9�7���$~a�� A�.V�@{�|Ő��ڭen��#���ͩ�I�U�cS5��ޙR� ��5�Cu]�!D*4�+<m,{�����L��35z��M7?~��o_oc�✮]��mz�J뭼�Ef�Y�U�E-���6<o1j����{}S�R����5!�Sw�)͵�Y�2	�Hbr����@n���61�;R;��]k��$�Y=�^�U�_�P���_�k�Ϋ��$.�Y[39h�E��d�����ʘ�ž�u�I�2�a^h���}n�".
Ȇ��0>��f�X�n|LY�(r隒�!V��T�M��ǂc�dj? �~'F)[���kmU!�f��hKP ���)&㥍��B�fc�Ƕq��Gku��`��*��.ˋ���5ۛ�ρ���5=kΧ����魍.Xab�KBRh�+�i��Mlj&)u����2)Zˣ16�G��������TMx;n8y$:<9޺ʧrr�pp�"bnd�����E9�U���v���k���XM4B��,�Bu�-�5�|���eqb*�s���e�3e���\�����
y��D�gwm���H7���́�K�H*��^f{�&{��M~ǵm[�2�%X�����Vg�oi}޼�u`�):O�����2�FԱ� �Tf��I��o��-�mm�=��M�݀��U^P�~�r��}6.�3�a�/��e q�C����������N:�����y�k�P��=<r��O|�w�Z��G�΃:����O�۷[��tU�q��o2�y{G)�+z;���#s3�B�|
e##1E>P7#6O�>��s�v2/�u�W~��m$�[�@���A��6Ϝ5�W.�U�k8Ku�e����'t�V��������\E�se]ܞx1�l!���r.�Ż
t���Q��y��_�}��9���8��T��c^�R)��=���I�(KG0��s�W��k��-&�kY�kA1�2�E\���ěl�t!YB��.����RA��<={�2<��h�xE�1"�g����7j�z�疛:�w3F$JH諼l��k��9+1�g���Ѱ�*G��Z����:�_5��+�Ғ(m�>��,%����y�(�k���P~&�?K�|�JTۓ�,�^��W���#�Ѕ��K\�Pa�a�A9�£ٔ�(�����̗r�k��i�+B 39}�T���bP�~}#�F�W���R�ѥ�>���"^w����G��q��]��sY�:��ٳ�|��[;=�����tu[���y���� �Mz�9;�����(�ݗ����FQ�WK�m!du�[���`{״:����܍�w=�m�e�c-R��& y:��k�y�0��g=�ia%"TG53&]�Ȼ���Y�+fX�b���U�0����@9�;�eN|\�Ab�):��>��UuԿ����9��x����F8g��y?u��2�i�E��W+'cK��DˮhVv$�:���z�Kuǩ�AYr���]��'ژ�m�;>�����]Խ����!�o���|ν�|*e%�k,K3�&��l�F,�\X�;1&-FSF�԰�H��fӌ�����������4��N�;�����rmD�*
$�ӝ�b��3�x J��L�!z���g�Vh�e�{�X���
HR(V���u�ZX&!�=u�պ������ڙq�S�20d�!xJ�V�Y锽5�w8��=S-��a�������,���a�Q�.�ʅU���^z�w�-$�Hn=7̛J������>A5]�qt�X�Q:_g���*�N�)7T^�4VB�)��:D�5/ܵj0OZL���V%�_5\/kRB�r_V{E�w�4����qW:^P�Kö��Z�8I��"M$���[�Ց�����S���,!����\FZ�i_w\��]0����o��8^MQ;x[W�;36�)ӄ�A�t��᎐��jᝌ�/�,��;#�������s;p��m]A������g����!�`�<�/Չ��
^գ%��v�>�y8�x?}������{ގ��e�jJ��`���^N҆���-�|Ee�q�r3�� aZ8�ӎ%��yz�"�
�s����t�wl�ޘ볌�:�F:@¨ejShb�SGٺ`��wG/���2����%$�#�Ts.#�w�>�$$�SY�5��%Պ	ق*�6�!�_�ͥ�5�W`��2%+:e˭
���u�|�D嚹���Is�g^��DŸݑ�1�`�&�k; L�pmc�a�Mty$����\�9�XUo�n�����opU�㲛`�u�Ę�;�>z^s�Cl������y�\[�)��>/Roj<�r�N��9�
����&�J�G�;��.���WxS�4v�W��T�:n�#N�����IU�׫9���f)H�Ty$���
vǥ�F��K6n��S�u:mTzry����q\����Kݝ���C�s����)�K��-��K [��pYJ�b�m��)�9�-0i�^k+yə�5��C;)��0���zb�
UrN�t
�� ��[yt��܅,%uY]������Հ���;���}6��6ov[�ۨ���5�՚�j@�o�s����G���\���Sᤊ����u�8��Q�EcN{_�?X:S�ӽ��#"i>uȱޭ�_�K�uA�oCih��M��0c��%�ﺮυ�,��Ҳ�W�ջ�r�F|�MHTuT���j(�
Wzz��y��v��2*�W}�W�u¢=y,��=��W�ɴ�SƼ(V%��+	^��E�������:(�b�iפ�N����W���#H��E
JL�}�Z��c���Sr敤�VB�*[Ie8A��B�׶n0�\g\+U�"HS��5νg���7�.��!>��8�!N�����p�.y��x��LOZVF5r@�b�.#���z��م'�3�4�5��{����OٺX�ݬ ��#(�l��U睰Nú�Z��tl���[�kH�+���[hT�8xA�bȄ�P�Q"Z%���W�#�����QdD��h��J��|kmŐ�;�V�dp=Y��X�9��'c��dpP��MP��kn��kD�I)�E	,��-m.�D�Ԓ�U5K!-"8�b�B�_@Ĭ�]���p�����V>r_;%����	7��dE�8Bﻼ-Da�DiB�;s+�t�s׷^��.81(�%2��{+���u\�\:����jt�o$Q��gk�����ü�I�)L����5.�tK��P�P��*��$Vg��!�h�QB�+�E���mMƠ$����:o64��*�Lzw,�HX�&�P	w�(罚�,:CWۘd.
�l��������jCA\�;�/'�µ�ȋH�ou%~hn�9��!a�E
��MLRD.���BX$�"]"+vc�#D�y�b�#1�B���غ��S�^��Phy���Ⱦp��%y'}��t��Vf�D�%ė�ڇ���k1�Ԩ�:7�_���i����aP���+mmT��d�G�/���f�T.���VBN\P�Q
'ǹ�":�9�Q�s������l�붔P��;���IJ�2�2�UM� ����:.�W^��ݬ�_|.gO��4��*ZJHTډ���UW+��p�H�$p���y�j"�X��BYNW�&�=���V��^r�!��Tܞz�jy��:^�\V&�G���itv�8���A��UY�&Ν������	a�G&��Z�:B�.���X�����X.�$_�K���O��!24��������*��s��݈�Dig���a��[�^��*4�DD�����췜m;��E���L�EN�����Fێ�.���M����.կ�ޓ\��J:B�P���,ʭ��ȍ��I	h��"\%&!h����kS�K��
�JHV(�"\(�ϱ�֘%�JN{��ptL�)��p�&�'U���z��*��iv�p듫Ȱ�Aƕ���bV%D ��z������RjEB�.o�8$�O��I{��J,��*:����sZ��B]"#8�Y[훌emD&G�Ʌb�b���Z\Z$��X��.	[iP�HO��/ŵ��������|�\M��p�I]w��w��Gb4�*Z��N������IP�X�P���	.g���pP�uJ�	P���LJN.8��{x\D���g�+J��(�K�z�jxV�Dvo�7޽�.
0����
&���(�n�u%R�.�dF�:�R��

H�_�7ӄ�t�H�.e��V8�r��y�����u]ܶFY�]#՗��͕>!+R)S�	y��7��J/���
��cJH����k��N�J(Jo�
��
H��uy��y�'�r��S�X�fvfn:Һ]��YO	t��n���u�V��޻W���(wx��y�e�>`'�����-���JX{�QN�!�r�Qٔ޳�ۡ����F�λF�sj�f`V�l{BY�غm�v]s��p�2͋sx�9c�#s��Dƀqm�y���iՅ�be���X.]364FЗ;��<4&�Ep�JA�eR���<c�q�<[u���Em��6���*�s�">=��]���!�[���:Ae�f��B���2���eY��\���@�܉�oEp�Ʃ��CZ6���c3�(cd�8e���3C��
��m�K��ܐ h4�یr��$��>I|D&D2�څ҈�y*��|]��\*"���!U��4�g|�!f�
H��$JĢ�U�y�ԉ��{�T��Pȅ�Y�VCO�pP�w��F�FM�/�!`�I"+����,�5F�gs�y�%��緅��h�,��]�ֻP�[�̙k�����a �VJ��y�b��	�͝�����!X�v\)~��t���f���!pK��+.
Ģ����{˥x��M�w�û|Y	X�8�*!P�9>�zদ�\Le{���z��6~�
(��o�U��H�[��L�K���G�!�q���ۅ';w�6M�؎
0��	s�A��Z���Bdx�\��T+^�n;���B��BR(�,�s�s�}�6275���B�q�|N���B*�~�}�W�m��
+�^��J��zn$�௮0�*w1D`��﹪�xQ�a���e$^J��&wٶ�*�6�$Q$���{��S�	x�89U��\"�䥶�	QDtK���/UuST))U:uU4dI��q�V�-!o��+��!�7]
:+ 3b����Q>�x��!p�V�YH�\�)#���p�O�H�vݐ���.��]T��ۯ�0��j���~R8r3C�^���u�;e��WXo��Fط���]WV�p�,t��m<n6��\�<"m֝H��ꋔ����6p��Y>���:��p��w�+V8�8Q�EӋ�o/l�+�$E	2�Ԑ��⽹��x{���S������VB��Ma%���J���z%����E�RI��G�UH�UKNjji�ZD�JD�(�+]w;�c��^X�ݝ޳�ohb���h�7�jM�y�C���l�"��/nv�z��6��\{Go�����m��Y�jr��_x��Ci'Ʋ�Ta^Y��o�~�Q��
D�EH։���VE�ZB����,,�w��<���/w�k�}U<ǹ��Z*������}�̨�(��<����,RBR1/u����j͗+�
V%�$�"�=����K�N0LK���5_����4���e%}�����=n(���*ӄ�Iv��-z�Q��D�D1%"gW����]Vd*�1�9�^_f�~�[�u�6�'U���Kᴀj0Vᴯ[���%bRBW�ߵ�'���Z%��&(���.nW��Mƀ�	�{����,Ξؒ!�����i&$�rl���VD?^N�R�e��2����(:�JE6�����-6�1Q	ۈ�y��u��gn��׳�����j�5"��e��f[�ĨU�YdxE�����4����J,R%(bK��m
������/H�m�SөLCˮ���Q=N�v찛o	 X�*R��3�yu�#�	���G��O,��i��l���=��m��Q	Q�Y����4��]������H�k�_��T�ճ�iu���.�Hz���"�q�����fX�y���P��� �X�!t���iب��p����ﳼ��z�6��^"9MB��3�W�굜��T%�j��/V_�q�R�#�,V)H�������RBP9��]�C��(�F�4�"AR���f��Qp���j"{�6@B��S��V�\tF�n
:���ɷp��\�j&�{Vo�]�����k��0u�Y��w&�D6��l��gt*J��ɒu��f�*�3^,E?��J��|���yI>x���&�s�9���P��e(6w��-���Ր�[�623=�M�ɔ�
[��Tm?]\$?On��a0�R�2A���a
��)^��W��ٝUN�\��Z.�۟g7����#n�1*!)$\�W����Bb��S�J.��^���+���
9�}w��'��sx�<�\���������;���W5Ib��IiiDE	0b�r�\B�&F���Da}:�\�!Jz�r��}g���iYd�F=�.\iiS�TD��=��a�{��5�*ۛD+"{3�}�f�����8܁��'l$���S1X-�񔹇�tګ����]`��*�tuC�%4S�}��!��눑.ׯ�k�Ӣ������D^:��Z�7�],�>W�a�Y��N��������=���j8�jȱ�w�=Go�����L���s�:�v�kH�`F�'���Q��*<+1�Vg�P�ZOg�-__2J���vEv�W�׋Tz�)�d_p�ԑ�ZB�p��s�9:����8���R J��_#�����r|]�n+��������4Ѣ(�Ef���&�qG!�Zi"Z)�͸���^�}���s�;N)"��}j�Nip�����R�^2[y�KO���dtRt�"���+�J�1��LQ'�IX��+{-�wb����u���z��H��[��W�s�o�q�29ܾ+bX2�J�0��i,y~�܎��UEۉ^��H��+�>f���@3�5�g{�\��y{=;sZ�hQ�HcdW�qK缸u�7m�R��O��b�z��)&6]Ђ	T�[������:QW���ё�|��G	!]�}�%�M	��U.���N)b��Y@�����^֟q(Q���5R�70�u�
�.�ĊK��s�~-.bq�in�(�DG;�|-d��
���Q&QD���ӝ�_:���ٍ��DҪ�9)T�5κ�ٻy܉I`�ݞQ\�ښ �$`���G[��DZ]AU��]�w�y-��}���S�0JE%K_s�W��Yq|q�4�QA.]w������+��I ��^�żM7R��Dz��:�"fL	��NCC�Mf������!��:��f�f<�;��] ��?
?iν4��8*1)�Jk���o�*&�&B�wׇ�51E{�}�K�\�sHRB޸�"�lΩB��324�JNf�cJ�\��kޝ���Iaf�j'���e?.���o�I%ʿb�G^�O]	QE�۪�:�ΉZ&C轲��MP:�UR�9��0��xү�bb�ڟ_�{/F�g��vx�+�����VD��,��ھ�ds��U)��}��_G�ͫF�;K#�����U\�;�!�9wq�qJ"x�|��{��G3Fd�0��=�?���;��cQ�WX���6U�tE�����ȹ��ܷ��fؠ3�OV�"��ʾ*��_��I������JΓj����KE��q�©&�1��=/}A]�}�[�Fe�����٣�h�)a�eo
flb�XJ�}L��Pn�@���z�qv꘳B�e��	��ePk^����ez$py��B! !C��җq3����d�/k<sW��>���bqY۴Kk���Qf��Yu"�����ׇb�,Hg=y���!V�WW��Jƒ�?���^�aY��U�to5����v��!���s�����cڗֻG&�od�ص��e��R',�iX�C#b����4���/<��\��	�<g���7v�gx�5�"�3�ygˁ�j�ݞ"��a���biHFfg�1���A"";���(�a�՚�"�B��
���׿몱t�I
��_g�ai{�+�P������f?�R�>A�z|���s`���b��֑��D�.f���1^�4�~��Hs/���7��m~9�Gv�sA��H](�2�QF'�>qb�j{K7v�]ν�x��TE�"�����wg�v�JV�}tD��YY�V����H��h@���&[�Vҹ�u{��!����׽z�\�`]��[�<��υ;�z�v	�/=������a
Ww�����}"u�έWńx%�3w��=��c��D{�z�˚㴤X(���ߦ:������l��n	�2�I����� 3Dm�m�ӎ����0�ܝ�8Z�6J�dP�m贱_}�E�緕�c�k���0����w���0TE����a�ǝXi����VB҅w���۪lVG�����\�	��`E��η-�ˊ�"�	9�|��ݙ����������ݞ�!^W|Z�>�%M�,����j�[�<�.LSk��H(�!]{4�f�ZՑD���!��~�L�ת�hѺb47Ba��u�*�M%]����Ն��kM��Z8П�2��V8%�M5[���s��x�D�����r�n$Q�9�Z�7ZD�	���7ب8B#���^Ο�M��o��V�e�t����!2vj��U�v���S���m�G�;�0L�B
rB�6un�ռ�j��8՚�3��!�b���+0n>�
I΃*f�wB:b,h���O�Q� ��ٷ���z'���v$P��d+��W�'���f����u��A��$���شjb(|����� I�P��XP�7��-���>7��Ǽ�l;����{���9k5@&]�������=�ԝ�{�{�"H�{�׵����|)����]#9�f�['�z�wz���|�f��WTӈ�6�G���tǂ�(�uX��\�[\E�)4�.Ho�2�R���=T�#*�u��|M�JH�iI-�^�zժ�J�Q�U�)�o�>Ë��Ubj�0�O��Jkbt���mV���b�$X�w�]TKN��s4T�Q<\�١\[�!>v�[`��������N�y��W;ɲT��u�)
����+�"�.ԾzҡH��M{uM��%0D�MU�J�#��
/r��w�3�y�o�yϸ[:�q��
8�.���:5Gd�rX��[���f�G�k5	��͌�t�̓���F!��7)v��+2�R�&�"�خ�6��B�i�!������97���8���g����j�����uy�Vn����K0l`�Y���c�8G�;�TM���{��m3\K��t
���m�w�0�X����m���=�\��Ԭ��"H�s��9;�����[����9�]�+w��7M�R	.Pos�����wU���4{����\-�R�n��RXȯ_��bg��Q�⺅�
u}JVm�]�X�T��C�X�:p���2��Tm!��3v�����f��l]�H�y��[aב)b/�4���������V���0�j��n��jo�ⴰ�:H�������2�R��7�י힧͞�;[;�b؊;�=�V��5Jd#=�Ǹ��~��&�F��0��_�2�$PK����=[>CV]Di�/w��Ӣ�� �\��0���Kr��Op��[���<��cxN��)����{�<B�)[�+��m���کW�;��+�~���
�(�To�����U4���G���ؔ�2;�WI
�o���*����H*j�]v��6�9�s�=�=��s�n�$v|r�@�cF-�&Q!	�rz�ʈKH�P�9�W�N��ڝ����Lo����q��Smig�:��X�|^vg�uAts���-�Io}��+X�+���{y<�pu��Le�����N��/�ay�ټi�}厍���L?#���ˁ����VpR+$�<G ^��+ZD�ʤ���h!��=���wt]�J^y\�s���˴��z��j����a�4���/:�^V�y-�[tJm��D��W���X��5{;�wHgk��|.�|��i��e����(��ʲC��mgO��+o0�y�#0D�N��k��1��9���0��n�
��ID7��î�cq��}G䣭��P�i��	X-|�ۦ+m���٧y7�+���e� �g��R�x�v|q���YEZ�)���>>��%<��"q�$9�yv��z15h:�K������i��N�'���m�FiA�޹�Z>w),�,A	�n����h�������J����D_&�ws�۪Ҝ����+����ʪ��_��}�����jݽ�����~�NT�5�,ڛWa�1��e�-F�X��vv��u��#.)�����2�(���d0C�)�s�_����V<s��Hj#I|7�bU{$�(��2�v��ݛ3��T�.,�Y��ldl�3v�2WA2B
q9
������ŝO�3A}�~�_%~h���Mg{����+��r���h�
j����n�c�Oh�5�=�sD=�EbY4T���.@���͂���+J<�|���(�}��EX�܍{d߻<��
�y�X��ޑ{�M��
���S{��.h�П'
e0��yb�HV�k����T.Y�|�w�u�,=���h��3}�[7�*ķL�];��%�׆��*_��E�n�[����jvI��4�W��3^�ؐ�GٖoxLy`M4��[����PӤ�t�W�R�yUU2����
"'����
"?����
"?�DD(�Q�DB���DD(�Q�DDB���DD(�Q��DB���
"D��!DG����
"?h��Q�#�"!DB���"D(��
"D~��!DG�
"D~��!DG�
"D~��!DG�
"DlDD(�Q��(+$�k#
[K�O �0
 ��d��EW|ptPZ��(P(   � �5@ *��A"��(P( 
� ���B� �P 
����  (         (       @ P  (    @   @|��     c 4{ݧ��<.��f�	���7GRz��w��{j�T^ ;��S�g-%m˯CW�5����M���� �v�`)�������wop�����٢V�ӼgE�j�`����Z� �������t}�}[�uos�{�{of�����Pnw�I�f:�����G�/ov�q�k��[j�JE���i�     �   {cZ͗,w�jٯzޏI�;����K���R�:�F�Z{jkޛ�zN�C�޺��O:Q�'� +С�w���/�"��3jV�`�g���@�㻨�t�� p {�սt�Oz�(��=M�.��ݙ�xU�	=���X�ͭŏov�;�y ������Űe���[R�
8     �  ��ף����k���<� <���=��� �;��7�С�wm���'�Ӟ�otnݴ���N�o �AԹ�7�G]�ꞕ2VklV�Ŷ��4���{��E ��5NY¶��yQ^�\Zu�k�x��:�*�� �^�y��J�x�R�[�x׶W=�z
ɩRI�6��� �P P    ΋cE���:�F��\���2+��=��=
H_|� }�iJ���a�:-���>�l֗�:8�G�7�=�kiJ��^ ��-�6�nwUx�S��g]�ONF�ڶm���sЧ��d�Ѽ����
P{�� >���B��ܷZ�C��7�:6��u�Zx�P�6������h��|� y�B�!�����4kM�[�(z7�k�kF��z;��m6Ɔ����KZ��g�P    �  �톩���|���ڜ���-F��u/M�{o�(N���J�m�n7LS�Rٶ�#��h��={e�8 zoT�8���o�(|Cv4Ǩ}������A�`������燎׃A@ b}�p�A���|��%J{}}=���[E��(�}���4>m������1o����><ݬ*�����ί���R�4� ��?�Ē�CB0 �b)�22�Ri�@ ?L�TR�  ��	*Pb @�	J��4�h������~�?<&�ߕW���{�]N�7���Э�g;3Y��Q�� �UМ��d �BK	H�h$���@	$$�t �BI�$	#����~W��QZa�9�n�?���,Y]��[��ݹ�Άള��l,����-D�MjW�w _f`��0���[ł�st3�-lDu�Čg�:��`c{�����g�7�a�FD�͡�1E�Xq	�5��	��kS�5YCla���z���9�8��z����da��~y�v帎���n���
l�C�L�2�c6�G�$�K9a�������6dHl���I�:�����Y������d�m��{���L�x(9M�]��I�wk���z��D��׊2��ه���!�S�*5u�y�α������޽���9=m�<�ս~�VSգovU��ȵ��(Z���a�l��8��A�����	��`��\ڔ�h��v����\{OP��K8�\q�MM}�m%ӾHEG/���QD�ك;�Ṷ�֎�!c��X����v�m�4����d��W�+m��p�wǠȀT�l6�/�/��+fh{��&��p�5�qsv��������MC�C��[P��޸ ~��U�f�ҳA.ӫ������Վ��Wf�.��qWwT{'s�7�8&n��k&%s�qcƭ��������,鯁Kq���67O{��w8G��p��Υ�d�H�j��H5�;�)^���3�(3�60hU���^Y��N��!f��:�K�@�Tu�K����3.sgh4��<�&J�*�@eȶ8HѪ�-��Ze�kd>Y�N�y����N�ۣ8�K8�V�C���K9�����3�&:\(���pj4z���23{�����lfA*�➬p�˛�#.k��Ҷ^,�N7�#�#��fl��#�eID�Ƭ��B,U+�Ih�>�rm��P�#"*wZ��4���!r�U�al�bN���Y7�Ef�������vӼ��f�|�oͷ��Vc��i��^+�\��sn4yN�R�ⶖpwI%��(3-*�qo�p󥜂cːq��Mܱ��ux6�[p��Ih/��<2�
�.�y6���\�;wo�j��sC&�7�F�e 띄</����Bx��d��LS�S[�Y����a�ڎ�E�r��8<ъg1�4�8F͸w)p�5���t^bp3*N ��D�:���RG:ݓ/ ���8VS�P�xh������\���f�#�6wgu�#�977��{����4
�P/Oc�����5_I�Xc5��"k.[`��׫'={7=���#�Z����6����լ��qG��Z�#T�	�E�QZ�����.��H�)9��1��y](~k�Z�e�ܗ&c
A؂c+ۂx�ܵ�kZ�d�M%���
�茅�N���@���@]_)�1���Z�˔���|;h��[�Ń�?�1�ʅ��AW�Vw�<w[^�c�`d�8)����L|�@�����:;�F�']��H�&żB��/.9*�ܘb�E�P�ˁ'jmd�
3��w��w3˰��~�.]89/e��a�o,Ոr	F������B+��?,�0P:�42L��D#{���v$�wP���,>X�:uE�ֻ;���,�0�d�����d,��74�{q��a'j���H5��)�-�9s=@Uki�����pN!x��7������Nҷ&ޣ����&[g �U9�����p�ȃ{��ʵ2���q=񹤎�Q�	��RY��z�{�&K4*[��rO��!�BS�;p+/���	L�d��!�B�[���q�s{������2��]���a�f�l7R�!��f��P�ׯ
'"Ӈ�q�T��x�Md;�g�ݔ���h@ܻz̄�q�LX)UiQʅ�Hઽ�chq"�:q��g(DP
�-ʱ�;{�.�S�R���F����j�����ky@<N'l��'W����?�=:�h;%]��V��I�;I�:�:��;9ޛ�	f�^��F����9cɓC˹Q(�Zyjn�jo@5�Mꑚ9.�x�9�oY��ߗ`Lg${��n�vIv"��w9s���kXV�3tuH��񛵋�Zm��C�&jR��.��K��-��呍�X跪9w%=��(γ�^O�g�`�F.�n���f�5�z@��m�]]*���nmH��Om�;��!�Ǩ\}4�]�fob�Ҡ��::^�+f<;�g�M�!��a��wI���Fh�nv��w.���J`lU�Q�DVn��	;p�nV�jh�C�ګ�Õ�oI��$�Nv>͝����v6K�Kw��h��7��b�6�t��T
(���{Jo@\�c����uX�Y���fr�F�tB��
HVX�3x9�91��ħ�0룈uDj+,tqՀ�٫��^[2aT�wtj�;�.�X6��q�g�s�1wq�й��
�Q�1�`�qӣ ��۹#c��1��6@h@@4���F�秎�΅�Ԗv;l���u����G��<oO�i�>_����JVE���� `�	�=��&�����J5n��͏tT-���dk,��v1ݭ�$���9r��[�����q8�v����R��L7I:�Ͳ+�n��"���>j�{�b��k�k z�T� 8����V��h��Ӓ�v��7u��B�[������Ò�浔x�\�@���)�]��)!��g��8`BS�g]��ɛ �����N j�����7TC�ϤKs���5��w���y�.mSh �v(8��):~9<߽�������=~��*���8�HB�p��e�ݹ�7��,�x���6�v�z>����<�ߜ)��^��gk=D]F�s{��60�s��hNb�ܢ>��zOu@d�,�5j��n	{���_�r�]�9h}�
	��0��dqi�H�1�����%�-���N	���6n���� �n@\�V��H��n�pLJ�T�p��r4��4z���Ԯ&r�pW8~ajsh%0���!.f��+�C)�s#��lx/p���M��Jd�tݎn_w-�����H94�L�ӛ �:t�p�X��Tݻ	b
v��c�u(g;�h9�ɉ�"&��u氖X��Hn��+�H]R����$��1>S70�53��ާ
�����N�`����1�<��N�Y���)t�x�P��,D�&��C�I��ۼ�}4�6 ^�ۺ�j�f�xa�I�w�3\<9��&W�0�  ƦSw�y(۪܌�mSa�k4�kY��BR��{#�X�d�1ɱ@�aѺ�ץƸ�M~kװ��-�D��D�:SQ�V �_��Nfqw@% ���6Wr��s�n�A���Ú�܎s�1�7p��d��&�խ��ye��yv�Ж�:v=����gP3vw2�l�t�LZmPnu������m��^�۷�%�����&�um�7E̗4n���ZɻXܽ�D�V;o�oN�j��&A��7���G](,㑮���F.а+E�E�����kᧁ�Y�r�b�*�õٻ@�n�q�I��]�X[yV pG��d��HZ���pA�pT�ڽ�N�lKz��u�9�#³�-�Za�Tۄ1Yǽ;񗎠�u��lAD���m9��m��#	K�p�uv%��,Φ���Ի��k&�T$õ�&H)f�w�](-��3�8��Q�#��IB�#y�6Lo0M,�e��
����S�e	d-v6�.\�b��h
pc���mK{Xa���vΓoU���ɲ�j��F@<ӝ;�q�as�f�r��.�7!�&�ov��3��J��#B�=�7v�ک�ٗ�b���=�(���EaHEhۥ��kB{�W�>�E���W�1p���4T�5a5�gr�縝��ǺCٷ7b�:D�7q:�CZ��ّ;�1��]�3wxS{�:v�^��3:A�n^�ut�������zk���{V\�*.�9�����$�U��=g:��n#Ġ�^s���4]jp���[lٜ{n^��P*�ȉ뗱���b+A^:���RLZ
BM�Qb�í�e�b�0�f��e�ڵ\J�$��N��4�ǚ/>�QN�b�`�c�xD2���[�8���rE�J��JGӵ촶�9�J	e�2Gwf��y�R'��y���$Eo;��p,K74�ٕ�	�s��(;8l2v^�{ $��k��Է�^���;��չ�ߔ���)�,�"�mM젼ksvG0d�����A(��P.*w4L`B�mrᩢ���1将������6��/MdY�;۱�jT�9Q��ٲ��T���E��
��еͽ�^�g\1G*�7�&�CUÑ�K� ��Q��?;9�k;�Ϸ:v�lX
�Nor��_`�E�F�-�1U�2�ִ�ٸ({Aw�+Q�2ѣ�ݽ��4�G�=����H;WS96 ���v�w4�b���=��=�g���� �-�$��A�s{o��D�]s�����S�p5;գ�AZ�~o����ƴp�c��G[}Ժ���f���DS��	DoW�-
����a��J��
��v2 �	������}\���a&�֖t!5�W �˱n j�� ��>{�Z�<�ۚ�f]��spm�Fh���0(rjuk���{����|�q�P�����%. ^��n�+9SƖ`����)�4g7/\`	�Fλ���c�-������b<�q��Y�qn��ŧNr�i'8�J�ܨ��p�	��uc�@#Ga`c{�*4a�;�Uf�؜�O�7u�ʔ�ۻ{.�y����++�[��n��ON�8�ޓ�v�U.������T����7�t�y&/'o1v�9��dw5��4�e��Q(�,��f��{��z�������|��:V-�����8۝u�%��jf���N�6�e�.7wjmb��$ ���:*ۍ�DrF���02��V�N�b�����؇�{w������x��#�0�w#�v�\��3�-ɻ���Px���ל�1>��x\��������],c�g�Ei�[R��܇u���U�H+7V�q�/c!yP��ǲZ{���C2t�*c��u0^,�|2���iǏP�`�x�7ݝ��3V���%�U:?o��@�,2��K��v93�N�m��]iN�bq���bYT���ˠ>���a��C9���ܲԶ���ۛa�c���.�nN�$ʮ2��}ߟ��h�!+4���6Y�W��7�'�pH�cyj�%-�Hݤ��9R�f�	}�h���=C�Jt�3���X�Z:ືv��H�z��,��s^���צ=<g=M_n7۲mC�N�۶�I5U���(ۣ���`��A��lwxh#�tM��XNJ��t�<��0��eв]�x���w=ޝđ�`c���
f�f�XX+Fe�w����b�\ �v�|�w4�Qք���ɖGð�J�{���=��"`��B�{u����Z�hǙGb�]�&��8�\��mВr���s��{ڈ��f���{�b��A+խ�ܒ�&d��S�p �>���&��c�C �!����Fd�����ClITM]G���zh3V,&���v�i7n���]������V:�A��s%�Ev29�Q���wj�L��v�4�ɣ��yr�v��nE��`�����e��A�ᎪGQ�Q߶΍�;�/73��q\��ٿ�u���WiI+5
ؙ�͡��P�p[��g*����b[٣]�L�Ž+��^������3�� �-��ڻ���-�ܜ�,{9��� 'oiO^�&F�\CAP�|�!�	�� $�D)l��Ɏ�\��q)F�k^��~k4aiY���Lfiz��uvv=bW��އ)��]X�F���rK50�����d(oa�����LD�f�]�r�ow5P��ܓb�����@����unv0m�S���, $O6f���ǱEd^�AQ���ۘ��g���I�~g�t�M�S�*@k���P�g\c[�M��檲2������I9A�����#Պ0nޚ���=S�����եx��N;��A������Dr�p�sh��ܤ�G�n��`Z��������v��3�ƹ�� $c�N��+f_�+�&wf�U[$�[���9�/Ԛ�/rY�_/�:����&-�lZu�c�<���S��qޯ�b%�(�XO�$4��`1I��$��]����*�f$���׻��;)�P��F���Y��W�`ŗ��hTPZW0�9��$�^
��pl2�ke��9� <�Z�`�$j���Ge~U�.Iı�9Mj�]����\����֠�x�0m��B�-�ᇋ7�
�ܷ�4^��T�<y����n��[ݍ���r�zeP��oV�7�G��\�Bv��Qt-�S��Yt��BF1���]��\�=�h���+�DYWe�C���P��QV[��őN<u~G���y���B`iG)��H���Һ�0�ȽM�W�L[��]GN���]�=͞�|�2`�ׯb�2�Z��y�^�c�	����^z�nM}�.�s�:��{�~�6�N�!2)�NʡZ;��Q�ע�="��ѾP��a�Ga<j��Ð�x7.����P��R�|���Q�0���<Fn��s$��wE5;�.p���5ƒ&���%յol�X��5̛Ӂk寈T�e˔����	���F�r�y��vNM�(��Z ����َ�$��w�zk�-
]�������f�AJ����بL�%��8aI��=;����HDrb��Xtq��Ib�����*cmV=Bj��nЍ������V�F�^����ͳ�w���̚
͏�������mH�l��#)Y]A���V���m:���l�U����[m��m�V۪�j�vkm�.�T�T�(k�Ҙ���m��[�oZ7]��؞on�m��EMt9wl��5;9}BՎ�m�$�t=p���\\h�lVrGe@��,s�ө��ф�OPۇ/�}��_<�@�'��n����tU7Rm�e�S���O�Ƚi��bF���9�=��=ua�<�k�ݛ�I�cv�k8���>��{�]!GW7�w�a�r�;�h��l��";t9p�wv���8�đX�s�;�C{l��7<-����9�%��u-�9�8;t��gF۹�I��N8�g�u[���g��ѫ�m��F��k�mm���)^KV{ݻc��j=�;��؍���q���K����]��a���� U]i��"Y1��/��Jʛ����6&��ur��&����^�.M�K�3�5�9wh�Aω�ykԽ]�U^3�a����7xgcv%��q�W]X�n{W�k��;0�J�7lhWC۬k�h�ы)"�g�M�+�Ol��J�ٵvU��+f��pt��a��l<�������8�,�;�t����vx�{3r0'-�٫t]]���k����L��]�vT{;�5]�z�۴�ʃ��]�D�p���Xð����dK!�m�<e����7^x�lu����V���-����i��iϲZr�\��=� �m٣"쏋�ݼ��=�xv�$�g��v���S�0�9��:�\#�G.�[}'<uo��|� �Qɗ羭��V˳RY͇��N��y��jDf�i;�71l�o-�<�D>�a��V�2����Θ3ݳ��γ�M�1�D��cqrn,�pYv3q�$� 
�g"����Ըt�0�N�������N��t�õ��<�v{/Z��HY�籵���uͶ݉x^y�����c����t�*���]�n��虵y�����7��'$>m��Q�4;qWGQ��m�8�F��l��al�rn����]1V�lm�#�e�.�Yk��u)��cۭ��f� �'Xt	��#�� �[D�`��;)�n�1��=�$p�t���]��w.=����v-ǁ�ᜌ�y��3˭�s�B3�*�Z\��ڻu������lbۍ��s2i�]��Gm�v��a�uCۮ����lmI�޺bz|X7Om�v;��q�cGc��Z��;d3�╭�F��^�4숺�����<���e��<�1��꛳��=<S	o ;q��۱p����y�����Wnp+&���䫛5���;28����/�e���;��.P��ݞ��YY:��v6�#q�3�:�k�#�"�g[@��:z�X�mv=p�:p�nx��4���Ƈ3�	�C�>��ծ�XNE��bR���sV5�'�s�ܤ�Lc��^�'��Tl��<q�[j��w@i��Z�4�9�7���g������q
�U�F��Ss�Sp {�v܌��-q�����+�1��n۔�r6�Ϫ�շ;xu��uvS[on�dL��˻J<;�*
dG��b|��yѫ:I�5���Fӵ�#+��ޤ��Ԛ�WnAⱕ�[�ѕ�:<�Ó� �5˞an�[U���:��V&82�!7����X	1�;G9�W��F�pru���ݸ���#l=&r6���i�v�U�;<�,I�&�.RD�4PQ�ء`뺑E0�0O���l�[W��d��yϫ����5�&^��6.l7.�]����i}�AK��'�n�f#�y�q���	���6���<�g��c�ƴ��g�b�<<�:��q�
��v�Np<h��P{��nL�^�㪟s�pV����l�kg��s۷E�n��'l���Շ�ϧ'<�*񗵽1�8�v8ƃ=v9mf�};�v쎖�v-ۋn��൷�Ⱋ[r֮˩wf�vx�5Uݵ�!^�s��n�h��q�*r��z�y������;��u�:4�ܽ�]86�aΎ�u��7=�-��N�����ϱ�[� 1�_RM�.����P�f�Ӊ:ڧ�w<դ��n�t�t�-��i��=���pM�c���jN�7����|�ri�yMd��a8G��`��e�^���r��^��u�=��Q�ۮ�h_G^���B8����7bP�fЅ��u8�c�k]�l�e�����:�7<��'\uu̹���۷A=8����؇��p��9�0���1/ucu���*���q��x�hAܽ���ˬn�7|����Ԩv��V�sۘ��sRts��5��tΧ���mQ��ۦy����n{A;q����۶ݍ�ذe��}�;;x�(We��#����^�Y�x{\�/sg��j6tv����ԋ�;vf9�\jv�ݮڦ�����ʎX�;�#˒���x�7lkջOc6��H4snZs>%�±����j�Kj�6���Ӊ���v뭧�O[��Gzvܣ�ۇ��-�^޺��4�Sv�H�co6C���觨Ʈ+ϰ30n$�xm�v�:yq+�wDp
�$�S�l�VK�ǹ5���R8�ݧԧ��/q��=>����}�����40e��'�<Z�Q�k��+]�W��h꼖������+*�;� ��lm��&NC7fc+GoWl/*�z�ܫms֎��7�[fkq��S�;�N�a�:�Z�.�\�mx$ܫ�t#�G��:͸��7[��b�2�u\�ܹ7m�>{N�lF���Z^�k�;��ۜ�Ů-��!hd�m�X��FGV9�n�^�ݮ.<��d)���;/	Onyn�ɞz.ݖƥq�,�䭶����n�Y�\M`7�x�s����@*�S���ڻ%���-N��fI2 �k4��q0�	 �͕���x���<�3NP�It�Ի�`��-DU�ui�m���=�{2�.��G2\I�Ob�U����q�v��у���⣶nv6�����5�`�#�^��!�d-A�ۮ"�>���96�t�����C.競��v�.��q�<���n��sÖ��j�b����D�c�������>!��&�w����y�h��;kp���j]�ېxub�5�ǧ�9�g^.n���8��;L�K���Y�h"D�5�˭�F���^�˜��]o&��3p��\Z�'F��1�*�+M�ZJ��j-��ʬV�WF�[��������Instfj�m���r;��D���i4u�,o]����Ś{pAn.Mk9�ܽoUc����p�jy��ў�)^:��ݝ���̜zMq�8wV���s�v�';uQPfٜl�0ĭ�]�SqӴr�%^n[e�)�pz考��DcZ��=���{�8��qu�u�wB5ܶ��K6�lct��v�E\���
�����=��!�ܞ׍��\���8/\���t�<�#e#��=��tv�E[�<qB6]��a��^�����l��c��Y#$��qvux��"{{��7P9�l��rdɗ�s�n策�[�Ն�93v�Ƴ׍8kqٶ��;��]<����Of�P�.�n��v�l��hĩ:����z�v�{x֝�I������9��L�8����[!��0)U���4"�u���&5n��A�n��Ʈ��;Sb|k���WX�$q�WV�y�QD ��9!�L`�M�۶]����ll��qc�=ǉ�.�G]B��m�ڍ�nӠ�ø�Wl��N!N��x�_3Ѻv�x�i9�A��".R'��{vy�,�3R�prm���A��-ε��pOj��$�,�׌���:ڠ{m�����^�M`��uٸf6Uz�c݄��=�	��n��i�^�Q����I��t���\cq���8��7Y����)�%]�1���NS[b*�tCcz�\z��Z�cn�R����R�X1�N��X
�WXs��p'mS.�k��e�j���Ǟ�\r��ؑ��oJ���Z�I�&}g�n�-����rx�����N����78��pՈ�ض9흜�:-�D��ڝ;]��e��'�+zu��D �q6{Dru;��s��E��ݳ�qc�ۇO<�[l��Qٽ��\;>�{h�ǭ��{,� �>���I�mo<�N�[F�K�ڐ�ۮ��Ɗ�D�ON��5#3��ZJ�]m�b���^����ݹ�U��|�vݦ��p���Ccr��w\��zv.6�n�=r&�<�>[c�&��{p�m��^�:S6=<��qY�{���rѝ���Y�Y��d8�`l胩��i^�{�����59��qe�^`�n����4�`�Z(rZ����q���#��!	9m�����+c�A��g�m��]�+r ��fs��5�xN��z�68<�[��D�&�-ϝ��P��m�{k����懢��7E�	x�-�b�g$Rzݞ�P���q��2r;���	c[��6=]hn۞L��s�nx�Z-ikgvxψ�랺xƝ&�������4y�F�lp�-���1g��d��k��66yG;�km��y,I���2�Ԯ5q�;Im���Kד`Ez�Q^���0����j��]��>WN�,��n�q���ӽ������hv���kj�=S���\�1������.���PvB������xu=����Q��t��'	Ê��-�^t�;99�א�9Rv��;����Q�������ݸ{od:�:�)��Xk,i�o/e��ݲq�&�R�i�p1��ƭ͹���7b���=n&N��YNfl[ �y�nn�b:b��u���]�ۮj�s��̈x7hP��@���q�}�7'C������y[�쯎�M/N��O=�1��l�uqK�K�4���Ց�8���n�a	-��/k��Cp�.A�96����~:>�8������{nw\^r�������/%c:�t��]�9�]]�����:=/;��)�Jى������l��IZ#�����:�b��Äv�b۰l��n�ql�K�{x�]r<\F��Iϛ��6�������y~y�<g�!�w^^�xG�E�΀|�Yzڎ������^�n�-s��w]���햳��n��dA �� B@�?I%� ���$���I$no&"]�ML�T�8�j����3Š'�^�75��/mث��`�'�`�v�Ш�s6΋�㳣rQ4[��)�홤`Z�T�0VEbn���;���
�ə���*���`���9g=7k9Z6���C)�����P�l�v���wV���5)6◮T �1�7b��Ocr�롱��X�jS�Ku��b6�vv�4�;u���wL�E�	�ⴥ�8nq�T�n���%��n��^�f.-�d6��$���\&]�ܶ{s�3"rv�v�.r�����L�Gl�B�$�t!͘�p�D���%ۡ����OWfrQ�ob^dܒ�ǌwU��9c���j�m��Wf��̭$�f�5�չ���b4��l�ݵ��>���5�8gb�X��v�7n��'&Wb춥w�<�jݵ�:����ELֵ���v��q��h�CgÎ,._]�g�:1�3�єy}��#�&���ջ*l9�ûZ[u�g�R�O�+�n:o[Q����	�G5�GN�r��ua�nx�r�uЉ�pl�n����9�����[��9���u��F:I��f���x�x��@��qvv�v��i���v^��t��Y�m��Ofk�y��z[�؅���כ���j�:��.v��Mn�zĘ��d.��7�J�nWq�@��ɮ1���2kg�շ����6�q�.ss���6�������p����37S�,��j��즹cۮT=�\��ݻn�v㍨��'���6�%pv�c���5�ؔT���me��3��G)q�G�ݶy�n.Ʒn�9n1�r�]'�hn�m�u�9m[[�q��A�N;Bݳ�Xxy6�v�c�d��ӡ|U��z�q��F�u&_d�Wh�zֺv����:�^/�����E=�8m���x�ݞ]�n����wp<�J��{rEĻ\<��ۃ��\cv:�.���i��7c�����q�@nR�TqZ�P�*� ���lb�G1#����)�X�A��Hl ؐl�6�6	В �@l@ � �B�nb�8,��6X{��m�w*�`'�N����Z��x{jŴ�ݹ�z�[9�k��=nm�@��rn1��fǱ���{q�s9��� �uvЋ����	�g�����v�e-dV���<��b5��vyMq�!ֳ�R�'g�v	9.dN�ǉx+��6��V펍��<u�e�Ѐ��䢔 !����E�M!��U���7��q�x�q�d8<�'8��;#��y0�����w<�N�%#�}K����:[+6�JT�hwf���r��;4**Fn�ޚ:����ߛW*�1�Q�
�P�b߲j�=�iS�^D8J*/�9U�q����vL�2(�P�{��:s-4<i��f��@>!�*K7�q�'�/|S{�R�d*,S57����4��R�)~�*��z��[���������Ee�M�%�N�i��B1�������Ҿĥ�NO�ZD2�E�a�������SF'S/���L��&&BWz����� �LI%bkoz�"��d�qא��]�~3ِrQ����Sl<���2֊��ԯ��B���\p�L���m�6��2�C�;�G]��[Z��wcש�v�x�ٝ�w5����r���o�����~0~���U��2�F�/Z�!ן��E*Sx����qS&�-�t˄� �Lc���Ƥp0��7f�G4�Lηr�����|ߏ\��V��&������7�:���b0��)��f����逇CYj;�ɛ!N���<x�9<�����Irs�z^�9 }�9�H�~F<N,�z`[�f݄n���7����d�]��V=FZ�������_p~9Kע��K;��w�N[��2�P�U�_�F��2�.ͤDHxߖz��N���/�0I�}$���\1"w|r��wV���g����y��p��O�lwT�bhAՄ-��o�v*'��&��}��*�f �1�AnE#�&C{ ��}-��T-N��N���s��#u�ϱU�]*��Wp�A�$��S�,;)�'�SI�t��� ��w��+m�a<m&�z��M�(Yc"��Jӎ���2n׵����׃���rV+�������3�κ�����1���v21�k�����'~����<Sv��#G�j�ޛTY��A� ���;�Q��i�7�¸�@����ItDT��(t��{`�:�J�6�"H#d���ԃfR	��F�CW�#9+y��˽�þj�Nvz��ܜ��e��;��&����:��ݧh\�M%���6)+�(ou�c����h�k��p�軱����hJpƸ�]��k}���� ~�ͪ��`B��Z�'6V�ɎI����\��Kw��=�[-�>r�]��=��F��-,w��M;��B@�Rָ�5]�X� P�S��%H*�p�B�u�.�Ѩ:!
�����k�߶N����$\�}N.�Ck�~���=2�Ә��=�ۚк8z;K��Q�n���vW�s��� �����AY��Zt�<��v?�����C�8�+�L�ݒ���u{1�ÆNtdC���wa	����l��/�I'.Siv�8�B�R�r��1�!D6��@|E]�"Q���˒5R��N���^�IH�#^��W��u}q����>.!�����=��K�&���,�	Z�^��#��}��;�C4G�8�_9�ݙ1��������`��"�����콥��)�:�@t�R_�,m��A޾���uN�=���L<�d%@ÒFע!!�-�`�Ƃ��eҘ�1��G���1]���$��j�Nӂ�T����vV�W��s�6�ӡ��gC�H���u��6�k��,���a����n�g:�@�����fg<ˮ��p#��K{��_IH��PIr0�B4�m�n�\��{�?X����j���Fغ����c�� ^ջ�c�޽��swq�ɫ�n��']�y|�W��I���44AX�F�DPD���`�ֲmг��q��^4N{3n�;i��o���D�����,�d�ɹ��:�l�Ѷ{�ا1�I}��uh�`̧��{�� �;;xZ|1���|�9<��B�P�%�9�H�z�/�Fkr�=£�\��б����O��:����`Oһ�r��Z~�'��S�l�N��g�L|��,�\A�a�A�g^�D�y���@��G��'�TC�9^�_#��]&&܊�M�B��������W �X~�_\V�_�9�\q'w�A��Zx��B��S�CB���ê`^�QҒ�C��0��^�hTz,�8��u�P�3#��Ͽ1=
.#�|�ݶA�*�Q9�����z�7��b�.�v�iٿ���Mt=��o�;
�`uo����\/ߕ����*�d{'�v�r����+Nkl̏d�]����q#[�^n1�󞎃<R!��Zw�yc�Nz�fs�ۇ�㫆U�3��J4��=��gfd�}��<]�5�Ǎn�p��Z���v����~c[�g���`�f�g�)n#�c��ݸ�t��Xi�p<x-Ņ��R�P�a9de�\r��i7n��^�ԏs&ۥ��wg!�w�����s:�g��/V�]���v)#u����=oC�΅���;�N��\V�]���u����l�/=�g�ѳaͻF�(���L����/!�Cj{t��ҐN9E;Iղey��ON�Ϯ����[e�F)�
L���#	I䐙w���dwha���.��#��N��1��d-�qi�#y�&,�6��� cl��#�#�R�������t�R/��:SMz;�;��kx�?��/
"��+�t$r�����9����Yo�E���r@��
T�Tr5#���1~o6�uթW�D!��ќ���]Rn]c1��M�c��oKo4}el��k��lfu�X��hC 1�ɎD�i�)*T3;�<��z�)��o#��>:��qO��[���!�6��G҆͵>{�24p��8>��g�X9�KR+���F��IP���뻐M(f{��y��'�˒�`W��
���q������S���>��Q�=1T���?k*z�9f�����fE�q;�:`l�N{D������n�v��]P���v0�ѫ�q��5�j����~�E"HMџn����f�3�ƣ�>N�Zg�Uv�w�UqS��k�� (���_��F<dNy������	q���FXX�;��?�ھ�S��#(V�I�-W��zO-�"j�I=����,�]:��x�BsF��tFdl�2�:�Qsi�|l��T����bũ�ʲ#	�9C��W�>����A�K��D8׼�a�W�j�z��Y��PxZ�Cp0[�м�)t��X�ϡ{k^s��Ȥ'k�� 껮��Z��JF�	#��S�m��.�ᓸf5�G9I��F�ȥE�+^Mi_����r����+Č�e~���T������o��Z��2	�_)���Xa���ty����Ϙ�0�A�0���D�o|\hhĊ����<��ɩ~@��9�]V
�739�>�%��>/2��f��UWf�őH��D��d=K4&5����u��͞ y��F���#�5/RTčG	���uN��d2,�m����S�`t�ۭ��1���Fas��#_}Nq�Y]���P�b�:�����	��>��2zl(��ך�ިjp�7�B2�il���fR�+�rfg�Ƽex�R�m�����,\h���w�8�����PpGs#n�0lHa��������e�C�K���4�q}I��Ozhf�}4Ï�z�+�Y[�JO�k��>���1�����Iӭ:�׾;�̹����p�9O����KAh�u�̄�>��)7���Ë�6ŖW�d�������'�6�r`�,��qԹE��% >ϴ�ļ������\o�9��0����H�Q�U*�z�;۹wvb�m���U_b}$�A�����K���8�a#v�;̼��u�y�UfG���B0����'�����W����+���f�mÃm-���:���_"d%F� ģзQ�q˝�l��\<�;������/n7S��i�iŠq־���'[9h2��s�+�Z��xY��gMhCsҭ���ؤ6�fy�3a�B�F�	�#����J4������sy�I�L��Y�V:�(��Jq��iRVA!�[�t�UV�(��t��V�uv]���n��B��xQu7$�8��ܖ��ۦS��_Y�ӣ9W�WH}��oz�r|G��̴��: ���랺f�yo���l���C�sAH�E$���Q%[�M|.��{��}]:�X�@��ΤF�ʛ��?+��.�DsV�gp���*Cu�WcIgw�$F7��^�b^�aB����>=�R`��V��\hP��y��Lu J��J<xC'ҝ�]#��K�F�jU���Ӎ�3q��шwQ�L�ov����H~��҄�p�ɜxn�ve)��%��E�SjW>�~�� w��n���Y�t:>�Djb½Ͼ��ǰ�=������x�޵�Ós:�/ b��sl� D;�5 ���OFΝU������O�Q�WgJ��2>��k�9�� ���yL�,���@t_lTcǒ�wv�H�|��c��Q��P�G�G��U��"��kiԹ�Q����0�EZ�"��Uq���C��x���:>��X��V~Wo[@�S�f�,]�0���u��o�K��GQ@�����lk��塷��P� ��l�����_q��po�0#�"j$Ud"���y��W�zW�"�?~�&��v_`�b�RG�T�G���da���%�V\q���Ń��[�-_v����7X�i)$$�Ѳ�f��g��dY�9I�����b�}V9.�����<�;����{�!�"��w�-xm8p�G��}7�o>(ut��sّ8ϰ��y�Y�^��Αz\�k��Y�|���\LK#/Z���7/T�86R�Zǈ>�F|�~�z�mM� ��v�H����ܮ)7��n�� �q��7cvas�x���0yb2�e��]�uI�16�@�K�qQ+�j�=6�Y<b�/]��/�T��Ή����9��
��l&k���a��f�� }/]՛�����/O�6�i�p�l�B�D&ۮz-�֊ζ8�#d+�ɥ݋�1��h7�'�\���ʞ��FOe&����[�|�t����r�+�umezb�	����>�ru�mt�`I��lH�NA��Ż�B=�`�7K�D��:��7vV!�!5}Fw���ad|�^�tN�����K�[�;��8�|q��l�e��:��긯���]1�V�m(��1�.p3n��J�bY{xW����EZ��>8?1<Zy�T��s�"��<��1!�2F#�0ۋ�B!�O�t�+��Mj����g*�6���rZ���u���?T޷V@%�r��.;�pA�bjF�fI��-}�̫���U���xh}��/��]!�u���X��h���0aFb��l���ѕ�d�t,�ГX^���4t4�r�	��K�̯��΂�?G��7�"���(�v����P�g�Q0���ݹ�i�z�}dcXD<Q�W0�0�-�ճN�ă�Sn��kIO[���,�l���ۚu^˷�7Z�[���o$���z�\�7�S4@j�"�m��r�"���I��|�Ve�{6ܡ�a��@�q�օ��/67���Ɵ�FԆ����3�aҼ���A!]�
�s��J9�ZքA�޾YKX���M,|VXϽ�3��^�`������u�����N���Lz
�ޣ���_.�c�[���;�f[h����ک< |a!���ౄ.o��ˊ�#P\\Χ���v][hXiu�T50M�5�:��O���!e���y>G����t�3=�}\��ț �����j�8nY�����tzrT60�Y�&��L�
6�뱅b�lV��dG~���{ޞw�h}�,BF�vGF�����7+�FE����x!��rI	�7#-B�q��,�$n*x�>����:^R>�G�T��+.���d�~�*˹tu����2��ﯤ����Mz��-��ɲh�$�y�z�k�v-<����=�xּ�x9�<݃��^ϟb� ��ep�������q�ƪ�O$(�J8C9;"��t֍ڄ@F�'h1]V���ݫ� �|i	��F�PQ��N}�����U	ie���������և��]���6��s� ��Z�����ڠ�*
g�0P���
�u�G�9�_Y����[�J&�}>p3BH�&H2��!����^��WŠ�ofϊX%��c�����3(`�{��V�m�����{�W%��.�v/X��r����'�[����P` lٵT�'L�d����o����6"�[n
!'N�S��F�:�qڨsyt��p�����T<��8�m�L0��Ƙ�s�A8<h��F������]�DL�/	ʬ6����S_)�
�J�۶��;�kN�m`��4M,���3�Lˋ4�n�lݾ�W�C�R�_��,��Λ�'�W0o7��+ܷX����7�.P�
�b�2��;J�t��hcs���Í�岧���@�����P5 ����>LV$,<��Z��}4`�Wڶ��S�]֨�E�]�&��:[bm.�
�Q=y}ģ�gJ����F��&�]K1��;3��c�������Oj[ T��Y�;���t���N�c|k��OEVMd�Ћ�ϟc`��]�`F���`B����3�G���y�#uyd��jnT=�޽)�5gHs�wuûhm��Nr���@�4�@<n`�ucuh�k�)���£���Nup�Es�i<�v>~W\�v˨��F���3�+!o�O����O���N��[};��ݮ���J�{�^K�ӑ�-n��<�ΓY�}��G������d�p�jh�6�bq1��Y��Ptvx�%�yƣ��SM��1�d{�KG)N��\dݸe�4�)�Q�C�d�A��%���u�����,��T�y�l�h;㽱L���t��k���_Q��u5���� �Y�'�M�����,W�{���"�e?c��m��mX�����4���-������I���P�,�G�G��Ivٺ�K�}�7�u.1���Z#�wH���;I���"����CcQWm��K^.<~G��ёD#K�#��Y1�[0f��|릺���(��2�Xb�U��=�>��|,�Re��!�P�2�V�����N=�.1��9tA�ݸ�r�:�X�w!ˇWn���<�ݫ����#����.QÔ����]\E�{�V�T�{�F�@xH�|Ǘ���n��^�!��ە�K03���G�؆X�7 �ԋv��B��!"�J��Xf�:ymi�n�����yI�#�������7�87���5P]���jέ�0�DH7P2Geom	�#�w9W��As�[?T� ��M�b������~��o�H�|��·����Jw|�6�!>�8h`�|��f��/{&������C��~d���}?m9�߮�>����
3(�/��D����6��/�7���O���l��F��zo���u���˺�FN
rB�7��?	���u�E�f��i.�w�u��2�5f�w<mȪ��9#�V�Q�|�J5�^��Wר3�D*.�k�v�=��a�r.�^w�)��CmF���V��?SC7n�u��oeZ��h��\-[��K�-U�Dc���ql����1bNՌ (�h܊Q����Pj��l���=�Gr{~�{! a�e���������D����v�ɔ��|���N��N/���g�5��)`W��#��!e�dY�� a}�w:�B�����-���|���η�~�	�5V?�U�T7VRS0�����!\A�a��~l�����N��[�(n@y!i��;f�_C��Q;|X�a�Ll�/��'�]�I�8ۈ��߉�p�7��?ټ��@�l3�;N��+�e�Ɯ(a������n��f��Xj�\O!I�収1���t*$��81O�#w����{yl����7��d7�[������=!멎�x1��mP~a�ku -�����E+%]'�˱^@>���q�^�g���zp�]��z@�h�"�fUo���o�a�%�l�����Χé�l��Ɨ��xF�o.����O#�ѷ��#��ޡ��I��ꁻ|s��eGk:&�-��ݱ;U�v�6�w���{(RVM��ln��x70�[l�]�q1��`8�ub���qz�n���X{y������f%|f���b��f�4�W�q9��3�g�^����1�#mv�n��<=8�>�7b����837Z�s���z�U�8��[u���;�;g��4�9�nƺ7n9�Ͷ���7���f�^�mQ���hE)v*�9��U�-ˋ��/i{S�>kG<*ٺ1��h���A����=���S�����y�A�.�wY<si0�OA�/� o���T����_�Ϭ�U�{c�>{v��d;����2\`��I�cD-A�������2�#o��f�	|�b�]�(�!���`�[�+Tg�W�C���^�7�}��t}Z/��M�']o�
!�c'"����`x����ݣ��ueC�?�򞊥/U3o��h�rך����D&����"���'?X�����2�Bd�`�L�jWO�����Tg�������Y��@,l�HF��fz空"��&�Ϳ-�-q�p���z����$P�k��&ʪ�vYIQ���$ZD��5�}T���eu73�`���څ�Aa60|�Si��P�j���R�kFD�8A�%��h��P����d��:��[*�D��$�a����v�u��Wq��>����8�!t;�N���1)E喯:3����������X�P���],������{��q��uXS�E�S
W�W3�9)��ծ���	�z���2�?QaC:v8��Mڧ�3b:ڬw����n����>�F����숎,<�!��@t�҅��Ǻ��'l�1A}�3�bB�짩YG���
}�eر���������㯮�/�}T��%|(��}W8���$�fɤ�@��ec�7Y�5�f��{�1��GY��DRz=�@-K #'9�}�;�Fs�_�0��z`��4�(�EXB�
��7>�����7���}��#�*+�`#G�h�S���qq��K�����n��:���f��t|r��wҏ�p/��-��A�D������;�q�D��EZ�)gxa�D�Q�u�9��>������Y_
!�T�d��vn�լQiܧT�^t]����D$Q��̣���g��&y�n��L5����Y���֩҄vZ��l%b	I���v�D�ozWGv� .�7��QEpC�i���ү+�|,��/�Y�+�P��3΍�o��_e�� �l���F�����"$z�+{3E*5_k��2AG�����Ր�G�P����O�g�\�r9��j��g[���Q��[8B����F
�2�&9�WU'Ąp�]J���B��'gqH�ˡN|H�.]�.i�|�mu�<L3�+]�MX�������@ܻ˶������-t�vrw*�	���T����Nf^˛�^8~QW.��VU}����������c�TnZ��CS���uk:ҕ�T�EN5��v2�>��۽�~����/�E�)����xvf������;c~Mq��Ld�$J6�m�1v��Ϭ�!fyj���:�mK=��;C_�Uﾼp3����LQ���A��N\aҥ�s��*�(W)t1��Lj�VpȦ6�_9���yw��5���N�]�gJ�a��E����ap-���~+�$�i2��J򯬄Y�b/��.*��*[�˔/*�)��o�Fڃ��޳�Qj9(��D��*9�mWy���ݖ:�kb΃+S+ ���;�zW�W�#�FA����xB]Y��3���t��]���<�$,�%�\k{�J��@��vk'�R����nz�L�6��(9����R�(�r1i��+N�����3�P��������P�	�-G�!��C��6E�?b{=�Ӱm��Z��ۈXF���]2,UZ/���9�/,�3�Z����wkwb�8x�'�>�%Y�:�Y����l� U��\���m�_	�El���P]�:o(�{�W�2�y_]BPy�N��S�t0��@l�f}D�z��-�\���P�%��Y�I��}ECa���۶�(�ͫ鷦Ž�'��Yw0Z�7�N�<�Z�{9˾|[�
⽻��8��ǭ~T�Kq�M���4OKq��B�Z�ʅ�-т�#	+De҂���z�t�WF��+h�U��������gچ[�*�l8�Ƭ/��1��@9I�og��;���ލ��8a�%�YͰ�m��Dt��׉�$ l�㊆bg��R���Z"�Ff�Q�#��U:9�G�<B��]��Bk�1���^=��]�y����F��Ya�P�l��Y(o��Ǜ���P����> S��V;LS�')9�{r�,��6d�wF��|�o+�1۽{$�ڭtcj�^�5V�}�/�Α6�S��������Ex�9惤��.����a��\��t�Zp��Ȁ������r��P��D/4��mb��^�Q�k�<��$/Q,��H5�z]QZpQ�M�XV?H����(SΣ�*�r!��|-�C��ΜZ5�O�o��ݷO%��`9r5���H��p�5����r��^�/,6zP��w�N�zs�]~�,`�#"&�t��L�Z�z�o����s;Bk�@k7PM�c.瘌�.ם�TM����U��]����5�d�@7c��=��vmۈ���'3�Uȷ�q�����͖D���m�m�7iNch��nI��+ ��nA0jD� N��u���r[��g\�,���3��p�^9s�cV���Y�m��-��:��]ؔ:�rm6(v��6��j�on۱ƃA��G>��d�>2����E,�vlO�X�F�#,�R"4�N|��'$k�5���ޜk�4!{��ȫ��y\>��M�?��Џ�O��3	y�����#��Dϕ��LF�2G�asS����۾3>�#Z��đ�8�@bӻ��%Z ����OE���b2r6��p7y����o�A��(�M����A��HnExY��5ܪbr��B�zl�q(�DOzX���Az��=4x��>o��VP�b<S�qz��Ø�ҍ��F7��m���<ƴ�4I�{xH��́�mV����Ոd���X�R
���b�c��']�+���b@Q�#��I��J�,co���E���i(�H�(��̖�ZV?H�D�a�`�=V�S�~y�\T�~����wY^�;bv��\�����4)B�h�A �d�u�Ά�1��zc6,N�Z�=�n�)eƻ�^/$r���h�0�0��"�L���É%�'���(o3�W�k��q��J���Q�(�m�g���G�CͨQc�6�k]z��׶"k�	��x穹�����o+�lJ�><m�R}�VE��c5Aj��Œ����/Y��::~���o�c�^=Y�߶��{!|�j�!4K,��|�g���Q(u�0z����A%�Vl��2mc��/�κ�9+�q��1D2�u���{���[_3Ǻ�B$e,*`B��|�m���@g���=�75���Srh��m��KJ쑸]ɖ���l�񻢴׷gx���'漏���O���e��c%khϚ���*��/\�^[�wn�"���~�\}�ܓ�`�|�n#�X��uWد��ӃZ!���v�HaG<���>��7��ʵY���t������M8=�}'.˯5�|�MM���0���<�s�V��N۱�k�s�q���K�i�c�lhJWQ���!�<(�v��+�d��C��q7�!Ev��2�Ҥ'Q���A2Ȇdp�w�P��p��&��a��!8�q�u�RU��s��j�
;E?��1�����J���!�'�.�ܮ#� kW{�@��er�}��d`äC�_z\bq$	�'���H3�/�2��uӲ�e>����.��)�Y)�)�\�:��%���nWޭ�.��z��]ܳ��!�=�����9qЕ��
�V�l��GH=�j��5�&�-N�?��=�@�:�^�F�Zޟ�C�0�K��:�C%cG����������-��~�n�9�t��;EY�c=m�#�W�`�0��h����z�d浹��4�E��Wz�$sԖ��$������@/�z�랔~�K0�sj�׾;��.���(�!��46�����B9{V��҆�wݭم�M��q��Js��=�.�w>�9�y�ʧc�[n���(��DX�)(�B�IS���̙b��{^
�A3yֽ��(�S@v���3M��*R��,��V;
y�<Yɾ{�m�&C�,��E�>�Q��W�]���u���)
F��#�;�S�D/ ��+k����	�P7u�om���:���K�F���&�%�B�G%��#Z�͊�x���0��Q����H[�2�%��ɪy΋����t���Vh���,����G���S�����l+4��t� 7��uWD?W[�R�w�}j������^���g�$+��_r^��ٕ�J�vx2�D��kz���`SW��(����JJ�����#67+5Ѿ
ژ���r{�7t�.�;� �Iҵ|_V7I%��v�Z`�!���+=�|�l�@ּD9?$�y���Iyi�+�ڹa�Ƃ#�~��@Q�db!�x8Ѽ��1\m�"cW�Ę�m��W/����`㴽M�vnEP
�m:,��0����maR�p�q����W�"���W��([�%�KW{�@�gxAg�3%�ʴ4��.��v��G�S�������Ɛ��Q�{��b�/�DgX8���LK�}��#f����?8�&��'��W��W��a�.�gkZ��wA3r8�NI[��2���^Ȳ�[ ���$n׮ӘphT�Nm���̏�6�s�k.Og���a�O�|�]�,��8r)jI͝���N��?B��"�� �GL�eWEvّC���\E}�"8�zM+Y��r�9%�DV|h��[��(� m�P��1�p�Ы��� �!�����r�x��������>���DkW�,�����^>��[�3�9Ĝf���Ya���jqXaU�C�SqO딒�zE^^P��d�ׂTc7��n�yb���S�����Wቩ��U']�����RH�*AX��tr�/�7��{e�C�-r���*�y5T�\"#N(��f�w1��d���)���$���*�硎��f�~U�6=��������uf����rex��w��t�ܑ]�ro������N}��]����q�/+EK���|�����c�D�{+����ג��(��>�7w��1zd�+�x)�_.v&���s��]�z�M1aV	�t`9M���ya�o�VL�9�Ǳ�2v�d�Ow�$h�\<�!�����]v�y�Q�n���V#��-�(iU��e�WŊ�<鉠�Ҹ_�^��Q�cyܹe+{����X���� ܕ���y>Rvf\E��4�������|�0��'; �ԋ�����}��n#&�ŰTC���Z7���wM� ��&s�f���o(u�;v.�<	��{��^�g=}7T~��?<�:������Oj.�2ث���A{��Stk�]��$�^��:�S<:go��Z�s�k������Ma��D�H'�Q��i����E������O�#�%�GZۏs�a�ohv��֭�w��'Ss�m������_�o������M���);��������{��M��b�l��i��D|.t9���qה�q�����Ӹ;D���I�;{�!������%����ʩuZs/���(̑�S�����<]qË����x�� �g�������F��
wfn��<��v�'n��8��NS��P��7,�n5����<�\5�썘���.�crl��R��1rۇ��9�)���5ֱ�];$�u����&u�j�z�v��6��\���=[��.�b���t<�c<�p���	@���۰ۇ�p��]�cD�Q�kly)�a�����k�-���K��u�q�a��4cԗ��c��n{�1�z[v��K��}�KY0���-�l˵���ݒ���=x�:��,�̜^R��n�Lu�8�`���m/]]�u��bx[���[�Xz:��ge��㩎wG��9�'�I��\�a���p���z��������B��i��;/�*�<��^y{\��C���h�����0Z�qf^�h|�=x6�]�{���ة�ܫ���Y﯁�㷳���W`��V7ޘɜ���F�u�a33�It���]�PnAy��gkz��bx#xys��tL>�nշc=F25�j���[����%��'Wb�M��m�f&�ۚhm�sl,�M���4�V��8���7f�g��f�͋���vp��8�1Uix�^�^�w������8o(�4<�M�=\\�&�v����N����y�t/$��6�m6�76������r]u]`8�&�œ�OK�B��j��\&=��<���śv��I��\j𧄤x���9�\p��v�{:��ƘMh��)A �1XR� su��n�����ƴa��X�����{R�=u�L<��M�^J.��1�!^ӂ�P�����1���9���l1;�i��]źۅ#XAk�C�Vލ�����F�{V�Y{�ˌ�:ۧݵ����<g�9���zܞ���ԣ�ș�,�6�kq���Ok<l8�Uݵf��/o[��F���5v8#F����{M�n��f�=nPq��4[��1s�I�٠㟟��|6���,�J�����h�[m��q�A�=P��`�����m��+ű�m��1YM�\��.��`[g��<v�k�vd�kO<��u��Mvz,�7c$s�mYpvP��u$���1�8�@�a$e/sn�=��m��=�{��r�ܱ�_c�Nm>ō�,v�j9Y�ݞ�\}�x�}�����b�m[0��V�GF��Nz�᮱�����<����&�Ll�Q�v�!W'b����=��>eݺ�&��)���t\���QшS5�Rq����J����S��W�љ���8и�)�
"z��(�������^��Pcl��7��-ΎP`Շ��/����IH&��%�\~�L�7�̢�J����OF�����Tf'e}��|���P\UC�{�/i9voQ�|�c�����28����HV[�����4A����\ì���b2��o�Hf^�hWf�����:b��B�G�s��O�X��,�2�1}�ڑ�"Q	H{�fg�t�t5�؃~�|/Qsр����F�]J�S�ˌ�;���m? �J��65g<=~�i�r��nד�y�j�2��q�Bռ�%	�E����vr�n�װ���9��œ͆{��֌������d>4�W,��f���8|�'���
�J�	�wMg���ڄ�^:z�]Z���چ��n�6�|�T)kLMB������Z���;��ZBh�w�߅l��9�����Y�3L���gX�{���`>�q7=^�6 a6#Q��rg[� ��p�l���1�Y��qU��S�����oQ�pf_[&'�9'd6R|���۵��;�D�ܾ�[4pe��9�7��	u���#��1c��j���؆j��/c瓳Y�!�1֮�ǆ�x�|�Y�y�0����0�,8ّ�xChJ��D=��.�NX�W��&0b�L����~&h~B"�{��Wq�HOT���|J�N6�	�$_6�h@��wdI��+"H�?4�O1^�.ŃB7f��X�Rk���\�w�!��b݉���Fd���8�t"M�&���m�?X��	�	��d�j'ޚ��[f��e���.����T�#޲;ז��Ry��)�?n�����~�#��t��b�ʄZ�A1�P�M4�!�
%���=���A��n�0,ra����n�"5޾�(�޵]X��g��t��9t,���n��}R��a#gOCW�$~-x��y���N9@���`�>�`�+�u��W���W��n�/p>�ȆN/}��l}y~�eR�}�ùh�V�����)���㑂b�Ci�ċY_B��ߍႸ��M��K4s�$9�#�r�uC�[ˎxtIzc��q�1�S�c�_�����r�:�>Hhh�zF=选aʓbuETE��{�k�յ��k����@��*-?b���-x���L
�6ZcH!C�8���/���'77�ӣ�Oj�OG����~�$�߯�;jg�^}U��%�%��MglQ\Q����(2�4��.���{s�Z1�3�9Ź��W�c���#��c�H���U��o9	F��^v:��/�Vv}����|z]���)��Q\y�x�bn'��Mq�!���ss*K�8�w��lv�I���mi������p��њ�У���]b�p��=�3wzf�'�
cD7s`�Ne�F���xxw�Hm-�3 ���i��
�>/0�����NY��Ė�}s���2T�~�x)���c5r�E�y�U��.��-��g�=(�����7�@�L�`��WS&�(�5����b������:�a�P��f�]*y<h����ׇ��"�%U�3�6d��r�G/���tf���<J�����!�y�Zl��-����/����Mu�~*���Z�\����[���¾��x��-w@��\x�]���
�����J����i��sj�G&�ލ�G�:	���8���H�%���d5��z�m�	�\ʸأ��=��\Y��5o�zqw�5����\^��<�?<�+��}��χ�|�ڊ��ۭ+���Xs�s��W{�Mywn А��y.�7b��r8���,AV�t�W��p�3�4�׋8�U�ү��?-2�HE��+���5��
38WC#M(څ'!)�/Yy��Ĩ�qb�L��+2�IǊ��E�:"�:�����|�K-��{�g�fy�,C��[��r�@�����*B�Bdmer��ߎ�k�M�w�W���rYС=����5��/��~ƽv8A�{wU��x���d�$�8�jD[��!�W�A��qU�y�s��+�PYy+$M|e��y:�QZ�QZ�ǵ�h�����P�@��Eq'I���N���]�B��AYn���Rf�"��3�<f$���(�T�s��#ɴ0ο�a���^��٭�q�f�������\�뾖:��q1�*��@%]ӦMX��tҲ�b��?E���'�U�����4I_:����pypO �E�{�������b,����rc�q���'�q��c:�t�9Ԭ��vq�
�݇f/F\�c(qx69��ڮۥ�=��`�$9y�Ԙ�x��.�P!Qb��H�4������v{c�+�nݭ���͍�R�"٭�S���I��������c��y8y틀r��D�WHD6ۊ9֡-���C���-��G�z���=�S	�y�4ڵ\�xŋ��;�||��<����U��$�0�{�H���M���;Q���hM�VB�[�U��j�X~e��y�kS�~y��+.E��u�s�br`��\��lIiûA_\�������C�6���+�Q�	��ن�b�0��/˭_Gx꤮����˼�#<�p���4BE�<�D�w���,U����'��V��T�*��/MqW�\��_{%�.�ܣ��VW���WE*n2�L����d�X�Hn�l9�U{�\�s�ڤ���v7+�U�>>�һF	;$�/}$P�Z�5X��Y�z��42���͵	8��bE{zd�������8;lz�~8&x���U�'[t���VU!��e���h��ri4���W �rݬ����sΓ&G��:�L�9��'�wmqI����r�{qQ��ږ��~o�6�3+��m����_s��x�Z���1�տ����X��E���E���S�V�˔r�5�����+Á&Y&|- �{�:���y�+v�����k��B\3�POb
,�y��VҎX٪)��%��UF��_�=9����fW�-4�����vC��_�o�F������O;��W�d��La:2���xl��!�^⤬Ye����TVA6��%*���֧uK��7I���Z�e[Ȱ�Y�kϬ��Zsp�k} ��Hۡ�l~t�x@�q�K�q�I���[GӦ��C�i����͢�H�� �T/�=~3���57�Uғ�����=3wr�R�b�s�u؛H�_T�ڵ��'�ER:���CW~:;��3g}�G0��G��^R����~�#�T�I}�F�Zm�"^��<�d͗�>�9��˃�k1Z*�hp,���pv��!�v�B(Иj(��B��QY)P��١:����cG>n+���ݶ+D����B��k�j��r����ҟ&�߷�I�I!���4�n�H�ȣUQ�y8�R;) ��s싆f�3���������g���C$�W�ٴʣ��/+T���; ��U�X���b~_W��ɡ$ʢdH�$H,i�wU�n,��o�l({��]��[�����x��R��u�X�Ś#(�85�kxy�.�Z�����5���k�ں蝵zd��3��@�=�k��K1��h��M7a�|7=�^�]��!��u��܍�Tq�$On3��yFΣ�d��qn�ip��un:s��0� ��=�{��$��?np��[�;÷���(3dO3r�^��BQH�c�Fo���r��Zb�w���*��Y����-�zz�4'��x�M�g��t�C�~^�c���!�!
w�~����9x1uI!`�llu�O6.�����]9���ZˆF;A��sEOx��I�!?D�3��2�eVn����-�`!u����Ȗ�QGBu7�������+rT��R�`G�/P�'&����|_erX�+-;�Ar����˪"Z%��z^�Ri>=k^d��F�yBk��Y���N�=��\�)bg�uUݹ�)!F�����@�$�#vl��ܫ����n������5D5qA������\��lʮ�[�X��e���g������_��8��I �@�&�y5)Y�N���o��{缂�>�}�_U�Di�̞���bz؍i�R�=�}9xꢶ��O���j@s`�6U��9�2��3t�VnR7&t4�A�y�xhۏD�*�F��n,r���Q�g���/ �k�����/����e�܇⤈W[#d(��[��'��X�L�+����̢�UH����r���Ϊuނ��b+���!
�q_UGMs�c�]w5�7����c�ű�n�g��[v|˗��=](������^�b�Q)om#sI�W2����#<��ek'�k�p�d��7ȭզ�u���~���{]�͝i���v���j��m�v��Rl�jF3�zx9��x��f��~m�� �>]��^_R�r�����V���Uo#7��̳^wj�����M���0BC!���{5�=,?�3}%� �Rɪ0�_U�{�P
�s�T��?wa�6mreoS.��B���qm��r�+�ʕڞ�|��b�2�\���63�
��eEQxn�����K�{W(���:�{�
��B-��q�q\��~���<��,�'�{9�}�MnNoσ�`�����~�~R���}�r�o�<c��h[���xss��^N:�\�3��^^/݉[ys�gjob�{�W.ߌ	*����hn�.EʎՆ��W9��Z�l,�4�2�N��ٝ�Ɖ�RX��coN�#�������^�<���ggv� :uڸlڂθ���n��ƞ���.t��vH��8P�;d�uĺ2��R!�Q��:�g�x�ll5F�똃vW���D�nv�77=gm�n7Gi�3q,�q��;d�8M�Y�踞^ݝ���ۯc���P����OE������H�H����������������+i{��"�TjM8)YP��&,ňn"����n���N�b:��m�I�l6\��b%�N64ʎd���e��ʆF�Tާ���'���}�^�M�v�K���Bb�S���{g,22�{2�c�
nD�r)$2���K�@�y����\���wVF����v��"c[���S��<�#��B-�-���iz��2�n�y���Ur��RJBnHe3z��Qx���0%�'�^�*������(���֗k�z!d9�<���uB�s��׃͘�2Da���X9[j5Xdɇ"��xر=�V-c�{��M5�!G�Y��:,X�#)n���;3ٷ��yd�0�N͓�B�~Q�Re)!n&+����]��ζ�@yRL�����1W��s�Q��g;���
'��{�٦���f��X� m�p��H�;q�b�2FS=v�-���z���w�<�ۮY'��[U����U"����Z�]7�UQ��OB�^66;���̸1Kw�{�O�@���g=q��}k�|���QIl�
Zfm�Nѭ{z��i�j	{��[_ UfʏQ��3�d5��ݔyQE�!Z-��Bx۲��۹ۚtԛ�`9N�l.�� �w��G�w/ދ"�2}5�߻qXQu)j�˾e��T�a&[|jz�c�E6��7�)ǎ�er�:��~6�wB)W���,�؇"�A&wkԨ�BG�ޗ���Ȇ�w�}����ٷv��|Se(�a�L�=)竵�b��ފ��:����˽�T�+W�:���z{���A��g3ɼ�vљ�.�x���}���� JF����/$�Hk+fx�:��̶'�y�I���"��)},�г`�9�:mV�(�� �����X��~���8�:6���f�M���øג0d۷T�ا����n������O����:��������i�/�����Rz�>�0����7S������)����Ꝙ��F�����R9(g�z�h�W��� �\�fC��j�:F���:�ג������펬��^�(����qt4�yA஻���.�y_��9���;�����)J �R�Nw�-6����!�˲��Yk�S=j�)��� ��؅�E�0*[��k=�&>���ƭ�ûc%[��3�!�O*=�{}vU�����֓4dl"�t��z��Nޣ�x�o�b.������WV��e)�{��}�l�s���g�����+v�v=�Cfb�}�#�Y�50{or�<Eu�J�1�wو�i�O7�Qol��9��iW���K���]���๧�Q҉Ȫ�Z��:Mr�AU�5^��1���񔰴�<�nHa�h�&�W���I��+��{���;}n�%=��cDt��v:�	hED�L�٘�f���i��M��Bq�����fމ�t�~��*�ǲ{j�<�h�3��F1_Eu���V��=�1oT2��V�y�#Ѷ�꼸�a�a�2�ߢ�U������*���(s=ئKW�ZE�h�8�X���̓8j}2�t0�Q��v�I��h���rJwk��ٮA��p�᪥�}]*����o5�����t�)��u�fz�p�|���ڬ�i)W�:��vv����g��b�i�5�c�oO�ϳ���}��/��M�s���o�WPoe�nUPw��"�,�l![ԪEq��0ICt���5�j�JN����vM�ҭH���*�q�ި�[�N®Ѹtdc��'W�nY��/����f��+v��5i��`on��u��_(*�[��L�%��Yi,q���W<����ͺ����%�a^�:F2�X���푳��r��U�������.7R'�ޠ�6K!�R��e���@PN8�m����E3z������-����/���<��K�i��ۆ*�n.���-u�or��<�P�����`b%��d���I_<�2?2�	��Ё�]�aY���:�ަ&����n���']�]x��J��Qd�s㶹yoX<(=�56���Ҽ>����:��n1�.�7�x6C����#v��l�zM�r��Pn�j����~�>Q*�Ӷ�f�+0��������o�Y�߯ΒA����om�9�ä�봈|:}\�RX�B��X�H�gw�Wy�y
^΅ݜ7v�����F�3÷}}z�;�:��}�}h��>˞���:>GEjR�o0���qG����F���s���\��Z<&3n��?�SI,Kϗ�XvF<�w�5�[}�[�¬L(#0�g�����t.h�ۊ��>J�dh�����W����M��5ds��ܗוn�����i۾aL�x�ϰ]�������v�ڢj9w1�r��_,B�t�rn3�S�H�|������ǡ���=ɋC�N�#g}�U7�&��Qd�1�Y\1#�W�20�bH���v��d߭�U/l�w�r�7jS^�e��>�!w�K?[M��yI���囔�9t=/��
A��s��.;q�Gs�l�E�d�#u�r�v�!ӊ�e���۞r�W�ᩩ���K��+�zU�7�_�d�im�G
_>ς��l�)����hajֽ'�nJ+T��tp]�	-#8��Fq-"�|�iX�z-0�/��Ǫ�]O}O���ق"�^�����ra?p�j�,���y{�,���_�Y<R��7J|�Q÷j�w�W����ȑ�y�ʄj~��N��7��-u�Y�3exտP����{=�ʓ1��1��Iǝ�D�U�W͖݀.��7���]g%��	�Mϳ��cy�w�:�ܹ�oj����ڵ�[����G�2�z�s�9)HR7*�ٳs��)�=��>U[M-�9�.в�Ϟ�>iW�̊�1��w��ﶎ~C1�����qwD������W~�Zy�[*�MI��fB�oj�u������(�&�ᚃ�J��>�1�'����_<+L��5�xhaJԬUYY!"|�@<�޹��G;�<�g�+f��8EhE` �5-���մ�";����bl�r��[ncƗ��Zݐ�u�Tmc,�+��緹�Ӻ���6[p��p�Wge�����=��>ٺg\�t��vƸ��n��7��7/g #���n
z&�nu����ڽ���;�'���'����x�q��SvW�;�n�X���9�6Ϣ��lsz/h��0k�8v:��u=�d�z6���y�r�ѐA
�t�?mՏʈ����yJ�/.�
;Y\�����ĝ#�O4��X[հ�!z�q�9�<��R4���"l�$u\�P/y��w��a��C�O������>��z*F/��/9�-�|��e��dw��x�S��TRA�����������"�;���g���g�A���k�tb�=��=����*�@ߖF��ԅ�#��/�|�/Y��j�Ö+����ލe�����b8�a�Z�������Ob�?>��#�xH�1�0�oI���d��W��y#(ٳ1�M:�K�!zyƀ~�B����k֝��w��j��!���������VB������#ɽEr>�6�q�r�p����ے���m���֔V�٥#�y/G�P�~�����8s�����W�27���.�N�t�݋��Y͚{�W���~%f�~��VjK5 ���R����#�.૯���G��y4��GCߐ����7Ƕ�4o(Ӗd����v���Y ഝ%�y�{Nr>�ܧz�4���*���r��sy�Lם9vW�"'�)�-��P�V�0��9]��/��������;9w�$�'�Ǣ�*E$�n�	]�~p���d�O�\`N�����9��}�q��[u�R���?*���]v�+�ұ�|"I&�p��������p!(�O���pp���.p[I�S[xKIn���n{�ś�+������0���y`)�� LB��_H����r���J����~�2����4���h.��2��=��l��\�V�4�Vʤ\}����H�#���(�.�m6�	iQ��Ʋ�4f�[n˔��J|��[2����X��� &���??_���T7�/���B�,�s�����̱^�*>���,��WW��/���e��wx�}�H*	b�%�n�x�"����vwC좈�Fo�?�Gf��y��!�p��Y�\O����~s�yǥ�c�w�6L%�Y��Z�%�Q�&y�3���)��}c��B?���5��c��׆\�ķ��E���� ����{p�WRQVIÖv޽6�ᱯ�M,Wd��F�p���{�g@�w��Z�v���B���ܱ��痔���X�y)��a�B2������n���ol��/��1�U����o�n+�!oid������U���?O\��ET�߯�rL��dBAn,�tOWU͘����C�No,�X�]�䕮�Y:䎻ޡrsX)�������+-�rau�6��p�����5��m�OC�3���^wU�nTvk�rƎr�s�TK�{^?6��ZD�s���)Y���jQ�OyM�F�&���@�z�r��
�"s	�{����u�u��Z�y�H�hO��2䛅�Uc�O�V��_�k~�x���)�`�#�ޗ�k�,��{#�v�{w�Y�F��vN��S��#]��#-�bj@�5O����y�n���MSW�f���]�C�^����MӫS��!F�<X���J�����`�؎I"��(z�n���-��eVz,�9,n\ǻ����·	�5_2���y,�Iԥ����b�&��9����	�{��W9�N�PL��j���Z���U7j>�L�
\��_xp���Um�{�"

/1�L"_`5~C*>�T�{�����Iƛp1}�(ʭR��W��ҵz�v�W�]�I%6n}�-Dyn�'(����W5ٽ�IL}���;)�ɜ����~��i�/=�M�#9>1D'̧$K��=n�λm�э�����yz(�[��66��E�M3���NV����h�߽4��;;Λ�ʢmK[�l�_�i�?т1�=H����[왠��r�6�)���"�7���U�����
��wz�g(�����P�DRz�/�el��㥍��|#TLt���|l��<���IB���\-�vj��)uTf{̼�tBhH��~g�sK]�~��77�i��yh��D�ԯ�{h��8\?}m�dp��F�,s� �vJ���Y=gViׂ�q�����$,V�l�!��;9�H`ou��a���о��	�^o��D�䆐F9 Z�����3۔�щ��7�)�w�=��b�,��y���{*O%C�!��]54�5���KZ.���Ǻ<v�f�@�n���,���#'�}�nֈgV�3S�����DU�l�)��|
��e]gc����u�跧`��EU*]�r�66٪MOPݺ:]v7[���k�tn{��8c�Yy�n��s�:V�n��m��'M]�v�rdNn���g����Z�T�HR���O�U��+�+��7h_]��C�9P�0TL��1��]��&� {P�	;�Jn��6��\��N��=�s�<�u�{�<m������<�^'g�q6�Ѻ8�9�9M۳<�9g��SlB�۞����0u{q5/mG�k�b�ۣ�����ʗ�+�t����%�a)��O�W���ߖ���e���o��`���ي������՚�7����n͛fZ��C~LBA��bP�wl�tmߎa��S�IQ��R����Ξ����z�-��H�%@���b���Vgt�!��&�w	�$�$����J$az�gvx�Z){x4�Փ�z��ߝ�W�@#�[�˿yo��oJM�o/lI�\.	��1����σ;�ʻ��d-��t�)��?��'��?@\�y�	�u(�l�py�1s�P5�d�K�B�B�*�%�;+���j�/L3�֬�N�ٞSk��~n�u�Nj���rn��,���,H⎍��� �}/��ds`�g��\�^�&�O��!���aیm�c���ݨ�5�kE�B$AmjBD�����Y �sÊ�c�߾�x��~UO3���{�z1Þ��������w�|$���"��3�N�׶7bG�y�J�{7^y�q�>Q��RE��z��)��ٲ��Ȣv������^u�׻Bla��<J��r��m�k
�rrVu����"jK˺���,JT�S�ԩ�9G�3y`�+QM���6�o��3���?�U<�P��9�,.+�T�>C;�\p"���c��W�����]*�9�c��+�=�ذ�`���?p�~V���>��p2{�8􆺩� HZb�^;֣Ӹ�^�l:����1�A��/�/�[�۴�(->�J�/v��Cb�n"����^��I]U%L��[c�CD�ϳ7�y���#�Vd2C�����������V�n�;⽞+]�V|�H��Kkw���Z+x���B�8.��N��-��Gv\��g�нu�۷��94��C	 �j�>6j���<������ix-Q���ޟ_����Mљ��{�T�˷���wIT-�iuh#V��i�p6b1B�gF<�ƕt��%�������ݭKr�ڬ��?/�T�ߪH��{3L��byt�Gܭ�4��p�׃V:�K��u]E�R�2|:$C��r�A���̣�S�ݕ7;���V�^t�V��Ns(�ggsޗ�;'N�y������o�j{�4z�#9��Ds���{s^�͠:q
���ܗ��^�����.���;�ݘf��n���T!2�3�	e(�)a�{����:��׾�{{v�^�2Q��B���;�Ox�x]4��6��3*���#b����ϛq�"`NC|�:�������e�@g�H�&2qr�����b�V��|-��ox�i7S�Y�ߒ<mMb�N@�	����G;��>��6y�F�kιݣ�֌=dЖ��q<g-�zG�Ș���IQ�ޗH��j�
�{�(X�0�B�^��Ef{Y��u�uߟ/��y���0^�$@�A%n��wwj>�ܛ?}m2;�������𢟤~L)�%)b�r]Ju�o}�O��\�@��T���ޭ�S��qC(�P�[�F�i1�B\�1	M�]�S>�������+"\,��乛}��|띃�G/��a��
��8����0,���K���rhH	�821<�vՑ^��7��:���V[��$��zu�s�R{'�9�	�3�p[�{��P�Q8[�¥4g��+z�����Wf��+!;�/a2�4��R<yg�9N"�}�G`�A*1M���kIy����d��'p�J���V��>���ʝ��m�ً�2z�3�.��A����3/=����ݞ����R�[�m���HI�8�Lz͝��˙���#�u� N�J��Wģv����7=�s�v�fe�:6�&��٩"��$Q�"*Iʛk�Wz��v�ߡ@I��g�|?%Z�|�%�;	�y�>�H��n��ro�O�X$��BZr,�j��@�{D�0֏v�ބ�'���\9ᘸ{ۣ�'1���H���2J�ƻ�����x����K�n1�"Ym! �)��>���uz��J��\���x�kj<�Mf1���؛@��y�x�GE�����"�'Vn�B�u�AD\��,@W۽{x1��K������^��y�">������Vmz�2��s�
�A�<	E�S��y�*��W��<��M�p��5�@�ڪ�=�[�y���z�uK6��,5ќ�K�od��|s���_P��ٲ�>O�)N]�`���!����V�Bw\��M��2���G�?7�L���lYQ*��j����q�v;} �z��&O�{�.���f��2�V0N�T�F�Ɵ�&��N��p��c`ɣ�xg6�ѷr��oW�2ѧK(���SM�)��bv�iG ����.�ʎ@f������}h���˫��١���R�S��9e���u�GU����:Рn,�Y�HW�.5����IKGB���֍�˽���k`�F�;��BT����'|<�[���n��[#�)p�;U3ql�5��g�4�Pޚ��5ʇI�j�����)��KU�y��$�g4�c8u^�뻸�����Xk����!����7re���*3��81�m�j�����/_����y�I���
nL�6<\��Oyܹ(-��_KIK|eno�����+�Y
���'2��\�88��q-����[��^���O}�l�'l,���Y��i���i�iJ�:+r�o��+qOsFٷ��|�",=�'?M�0�����i;�(������A��ٶ�ߟC�ڐ��J�pz�������6q�\^��K=r.�w��u�������
�WCX�����ow3�$z)�P�_rZ!}�S������jŝ*w�꾾�_U<�w��-�o4�������m.�Syf!�f�zUJ�aH������67����q��ag�����s���ҿx�GV��)�yl�/a�lȚ����ý���ۇ+*˭lY�mK�Zݴҳ��!��[f�Ai���ys�sO�g"�-Hݮ����l��}���zM��a�����8�^�];F��ι�[oO�٭�ςp3ϔum�s۷β�]��qp>rZ��&'cm뫻s��nXnß>^�a8�;N�;V����mj�e���Gn�޷;�,W#�;uX��v�I�{N�n�P5UƊ8{/&]�6�l�U�q0��^��`�{f�݃]���c�ط5�N�Rn&벳�g� %��[��k�ւĵ��X6,p�p�Ý�h���5�E�g���7ln�.|&������n�Ա@^z�$��/Q�k��;,f]�k6���ڥ�[[�rp[�V�mv*�oj-��b�&흮[�7ga8�g�������G=x��=��g�q]uZ%�竹��dt��3AՃ�㮃bS���y�۷m��qX�&��;n���t]��sC���c����z�Nޕ��w ��ݠ���]���4
B�9��۞��K"-Æ��]�l;nA9�=xw=XQy���N�i7k��n�񎔝m��)�W��@�&qp�7Ag^��[����9��<>�%w�x�5��F���ۅ����zFM�����]����cün��O����`ݎ܊���\O5uˎ�6;X1Βm�Xݨ7���;u��S��m�z�H�l��8�Y��x�ͺ�e�\�͹�"7a�x:�zls�+a���ɯ츄ΦH6N�����7�Ër����ݻF�m�]�=�'rp^G���\l5u��n��������m�!V�J%m�(D*;�[ܼv��q��gj���z�8.2�����Onܻt����S�6�ٹ�ם]m�H�^�7[�;/C=��r�sƹ�^ʏ:�vq���	��7n�-�nֶO7BPt9�IN����m�u�6���vl���{A�g�E�܅����7n�З	����Vs2m�R�C�l�� j�n�v��<��Ok���;�;	/ny�;]j��#���4��#�nJ9��qv�8��ۯ^jx:븍���qe9'���lގ7�2v�5n=m�V��v�k��ݎ6��v�얔W���w>���l��h�gr<Y�ڠ�h+�=U�:qm�����7#ۯ\ѧ��W�LZ2v�v�k����l��|\��'��7^���P�M�Æ�;��5��;���A �7��������FZ��v�g��O�eͶL��u��zٛ��ݙ:��e����.�s��{QҊ0�H�!�"~Qe7�u�n�8j ���=rkk���K���VZM��nK���u[t�ɤAT<	��F7+t�����t�Ƣ��|���y�I,����y��B���x���fev��b�#��>A����73�Z[��u�|���g���;���B��)��g�������/e�����Ԟ��|����"Q����B[�P�}`' �?��Z�.J{�]���8*��+�����0�s������z�Ƴ{M��Jب��)�9�5��W�Z�c���Ym�o2ct�Q��ty̫�ݝ�dnܞqeA��f<Z��a$�;Uf����m�{\��XM�z�[=���4Wnc�ӳ�����/�]�5�}N���3o�9gg�����w���ޯP��,�ʇ���R~]����f`�bz1٣��R�E� ���(a)���^.DN�pC7T��#�e��K�vnw`v��ۍ��U��g��V��6�4��Hh��ή=��ұZ�� �6��8:e��5�}휗���=B�^�/�)�c��OZ�j����L-А��4 2Gx��T!O3^�wx��BDk��X��?RX�:���	�-�5)�g�a����#���:Do�e$�	�YęV���OJ�ʩ����㭾Y��*7�����8Ad�+ާ�CX�%�/�zY�P�
�ճ��v�6
ϬB+��$�S'b?�{���JyӖ���$Y>��~����>-�n�}󣼍��{hR�f�_�{�X���&������sOG��١Chc�([[���b��mm�=Z�J�X��>�/�=�ӷ��8�X�Pc6��<s�8�R�g�K�1l(Z��a�/{�o{D����ԍa8b�2ub�|i�~f�X�ד�O7�H�6�oA-�=�30RD�o��u65g+n�\ۯ{+uv�&�s�Y��:��,�C+��ҮZ}۴8��{����-����f��R���7��uH��Q��O-��!���;f���q�U^��a��F��T�{F��j�":��ٹ�x&	9 �����:�sXЭ���O�[�U�__��U4;���7��׉�Iq	�)�����a@Ȍ�>���7hE8��(��
Z�g��e�
��!�^�g�,�ޗS�=�<��7C޹܅�n�8h_�yX�-�J%�cG.��kœ�\�����h#Y�����1�9������@�������+��Œ:3sgu5��FS��iތ� �pM�Mݒ\Sŵ=s�mv��s\v0��(ⱩQ%��'iB}�`�-����7��N{U�.vq���r�:�t�{�߼�܍��e�[�)����� �����μ45�כ6���Y��x�y�#{ת�^s��;��������-{�/�G�d�A�����R���B������vr�ܝn��i˸�ޘ��tq[^�=7h�rz��_g��-]{���Op���)
�L)4 ��p�ͯr�if��
A �h^�`�{9ѻ�w��KY2����U���31^��ɡ�_�̍?/��f�Ly�q�&^G=�tJn��\��H��,yx;�뒙���3ngL��K��J��s�>���l���l�^���5s�����i�}	�S̭Ur�Nz+1ə.�z{y<l��\;]�K1�X�TC���Շ<Tw���\6��)�9�͋�:��;�ӎ;X2p(��Zɴn�ʼ���v�)v�Q6�1��gG#b�w���7�P��]��}��C׎o��|����)�RCf����sl���[L8�r6�8��<�����e]��/B^������3��P����OP�<q�b�W�l(׵���B��@�!%��%���L���J��W�}�DAc>�<�\f�{�7v�z%h��[��fʭ�#�$Q�&9*�/�UŎ�ǯsN�����¾뼵���r��i��n��Ŀ*C����%�#�_z�r�8Sq�<�f(�Olu5���o��~~�qZ��i$���p���Kۧ����f��o��1
�CN���V�.9^v�V1��<��9����6D�.w#�z���T��ώ�����3jˬ�����YИ��ɪ���/��htYk��5Ɲ<v�^^(���b�rq�8��9��v�đ���[���nvcȳ���qm�}�p���N�=����� ����۞y�1ˌ=�;1u�oa�!��^ό�W�;����z$�v�ل|��)ǐ��v,�[d�s�-��6�m��[t�N��'���u��'��Kٱch�$����'m����t�ɝ�`�z�����ϣ��y�Z�sE�z7%�[+Su�,����nn�`B	*��(�vBEl�Ӝ���[����?ezz0�*��_���i`B��o��Vx�`�x9NV�.Ev�\�s>�i��@ۑJA��ϥz]
�y��!����;��u�S�lI�iw%�A�ye�gI�����`��2���Ok�Ѩ���"dϡ,�4��z���{��� �Sʉ��)�}�lAAb/��qy{1]����&�d�;=��MR2<�N{��m���,xf]��<�%��}Ld~��pF��K������ٷ���=�{�r�X��Fb6$-H~��H֗xn���f[�x���]�αTK�f���i��}�K�Ny#��]��>����&�r��[�uZ6�@"(ݒDN��^�������]5n`�2�i:^�n���ۖ����#�2�s���<��ۮ�=�NŔ~����s~���ZO�x�5E&��a}��`�y���ᨣ�k���L(�#�5���άϻ�YyԘ:��x�
�eϸ�ﮔ�eⓨ�]���(d��SFu�����Uf�F����k%�}%�<�0����C��1N�v��Tީ���$B�MY���/TЙ�{ޛ7F��������h��͡0��i���u^�K��T���ʳSŵ��y�fO2wn���ܳ��/���.�3ϯBY�xo�?5���0��V��.��򑛭yz�I��ꒌ�kLY7�&o���XY�z���ZT�޾#©��[��Ά@\߽��q� (�+������%��g~�ō��|�;cKyf�-[͕�7����X���	W�c�-�p�M�ڋ"m��K*��OO:�8��\�/���rl�Yۢ���wm�ۛ�!��Ӓ��Wd����`����3������%��>Z��~�.�.U�A���:J-ٶ/T~rr�+�Ca�hCUy��ǟ�+���#��=���{�0�.�ie������o�z�_)(K<�`ѯ�{��H��S\	� e�pZEf7�H��u�Z��z
�ح"�"a���Z�pE�1���3 �Ty���l�zgtGS����+�DՉ.:��x���A}���$�Qi%�w���>l�C��):VR���s)+�c�ǒ,�(\}c-��א�}x���A$竌�w��2R���
[n,��5���I�k�m�}�6Y�>�Iz��"Ė���z;��gaĉ�_1��6~�M����䗝G�c�Zu�%���Xx�i��/X�o�|����m�=s7�CP�Z�vwI��2������w4n;l7Y{m�dV�'*u��IW������gy�Y �GU��t4��F��V�@�?_�<�WQ�(��k�Y������v��٩-p�D�g~���fx��b!�麉p��d�T���Ղ϶b��wL�۲���4���k��]}鮮�d��(1s���<��H���K�vN���۰�^%���o��1T���0ͺ�A�=��mn�ʼŦ@�+���-�ej��M�v��^O^��d>�mqCR��<(�	�^?�W��[S�t�3ֳVb��x6�Nɒ�y����D�<r�K��0�zQ����ʷP�$��]nPR+�f��hL�ز�XٳՏj`� ⍂b,!P�߯�h�~ڽ�)=��W��nM�'A���ӳ�A��V��t��|p��ƅ��$�r@���M�b�M��y�N���-�G�
s�i�8��չÔ:�m��J�a��~&%�C�w���J�~�Y�R��(��z����Z�+;�%՗��*�$��Y�?+�f�M�	�ڠ����;��y��o}�6]���>��c��ق��=	=�b�&\2�W����P�α�3RyGv�^>´�# �$�H�^�)�p7��yUW�fL�{�' J�喎ߪ�OC��#g^����{�L~�F�L�<AR6���'!ݼ��+�l�uҷ�U�2�ͤ}���Z�eH��RW��53�,�����ׯ��ݭز�}�U�^��.B ��cs"�s����/�e���1߭�~��y�ޘ�y)��ڴ??7��t7�S[�I^��˝5=���G�����}(�/wV��ָ4��-��^�0����I׽xh��[ݭ#��Tݺ<�C׽�S��s�nM�{�����ӿn圽V��E�<n���3{;z<�nP䦇����wZ��x�i�561�����]�;�v9��O���\��vHzq�����b���a9۝�ތ3����ۗ�V͸�H�v}��]�w<T]/��ͺ�-X��;1�OUx�£j��;�ɘҒ�&G��.����(�$�7�K���N�fO�W�����h�Ϥ6	�l����F����&6�ܭ���[��:�=�m�<�<���(�Ch���m����y�ݻ"B9���~{$�$�
���Z�k8�`�~�16��,��&�	*G�� 2]GO������I�ߔzl�A�o%�����O6�>��5��̰�B�|��
kژ�2n��ߨ� �"q�J(R��WUUWG~�+>�8z��ǳ9ꦽ��f�D��{~�tp�uW��W/�Ռ)�GNw�D��|���lP~�v;0'/�Y��<OL�V�-��r��cvQ��S�*\��k��!D#us8�j�y�\�èS��3��d;�	�Y=���cp�/3nJq}�W�[wb�`ǲ����k����]�&8T��=CzuMJ�y;���"D�l���\D�NRʜ"b�q�m��	��@-�z㠏mu�� �D�ی����$J�޾�9�&��mN6��ag�7S�3��F_-`y���!��;}*��͈���<Z�H�H�ph�^"���Y����,�X�3j컀	r�,��צ�ձ{��xC�}��]�_M�ˑ0o���n0�w�׵2U�Q�}���0#�����N"���&_t6�U�gt����o�˝�1�߻�P0�U,"�	�W�kї��v{:��)�׶�՜ߕ�)�%�����Q�u[�/:6{b�޶��ڿ1^V����V���f�c=n���:�@��qb��,�Gl�u�e�9$��u�\�����m��A��Hk���}�_}����a�u�z���W�t?b��\�X2п��YP� Ѕ��U�D����}�F��2��3�����py������V��e�^���^D��>��>^Gڲ*ʝ�;ǛY�1���!�`h�H��SU�����U լ&�[������I�s�f�z<t$�(�p~��?P�݇~�x2���S���*�T߻Gr�mלn�����L�h|2��0���♾X�b��h��aO�H)_,T��'�ۭwh�����v�<�䴝�{�ꏸ�:Kg�ك���$}��ݟ)��U���B�8H���Z�'��u�R}�Gp�9���������).�~��d)He��՚/�[�F�+	rn���n��݁�ɱ2����m�bl⛧|xN{�Ĉ���$Y|q�R�Sk5VNj��}&G7ک�@qUW�o���/l��JU��&���7��ާ!�oo�[?���0?`�j�[Q8�R��mRt��N��č��:�yT:��+s�e�U�^�T���ˆBs_��:t�-��ٵ��?v�퐮���6�ى���6�ۨnA�b۵j[Mn�Hs2�Z0p@iHx�|��۠�?*!�B����GȨ/`V�Y��Z����ܯ����?����c�=���M��x依$��靄8��N�`:^��ۆ\�%Ե�&q���(�9�XVK0MO��yAJ���7�tiT�|�����tL�iݬo�z7jY�DYv�劜݄1���w�@��Z�P�FJ��8�غ�X��!]�U���]o�K[�^e*#�l�a�sa8b���^N���י#�6N܅t�5v(��r��7w{WX�x����F��0;:���*S6ya��xk������1'M�����ꬣ<%�`!>�xg��%&2;h%=ɞz����F�'�2Ǹ���5\����v۹�'�U��buU�B܋�My�\��T�l�+h+����P�ڻ9ȥ��/w^+��"8��{k<2���8�:���|�ՙk�]��q'�� �:�fQ�ϙ�L����hsoT݌bļ��ۅ	}�>Z��G�x� RI�ß���a����������q�F����Z<"���jM#���/73ۯՕѯ���-6�%I�t{1���a����V�7e�����K���E/|�_%N��+㱮p���,ɫ�M���W=�D{�dl1Ի$�$�:G��T���}⫹ĹBB��̷�MS�Z��Ϛ�)��2קS�X�^����XR9[��r�������A�v�Z�E�n�9��!�&-u�yb6��F��sep� 뛭���h�pa�׃ު�w׳ԕH�z�u���5V�2�ܖZx���}z�݁U��~���VX,��p�-�u���Ll�iۭ�,:�Yw����I�:{:C<=Ϋ/�v0/�n�xe,�~kk34�⫮�~��Ͻ.kg��b��H�+-°���ڪ�6�7yy��%О�1�f�z�o��f�[a�z�^o�{3<��ŐD$� $��R��7��}����g`�>˯�/\�i��u=gN�Q���y�������&�_���x����0iܨ���V�h[m��mCS�<Ŵ�Mk,.f.yX��y|d��q��;�W�_+Sy̻�p�i�ܢ7����Ĩ0�W�H#��(�ݶ��A�S��+�Du��H����F��MzW��{+��=�}(�J�ۓ\��OD�(�}��_x{�7h��Zm�\#�D� �D�����:�G���� �U$&���[\uqT6q�F�%��ּ��ʝv��z�u���7��^��}��9g�凋��^�k�OnN�Y��J��	�� N��F���G*�ｙ�x2�x����Z;e�S��D��ɺ���%�s����+%���N�XU�d��	�#Ї*EbIf��Wg��ޞ�2��%�iva�|�4�4}�4f�2͘1)�/�{m"ht"�06�n�RU�x��s�k��k<|�Vf{}��O�����Ѻ���cb�l���՚\����rB4��n*�l�6����z�mTz ���ܯehH^�Ky�ͯuﻒ>�z�ye�
�l����Kq���C��e��f=��W�Z�t��*IF�Z߶�ɥ6Or�dkM��]���Ii�(Hjf̅ϭ}�w9��[{�fkHZH2!D"$���&��D���W;=��q�k3N�=:��=\yԲj.D��.�9��;�5�8�VϜF%�^;���cc���p�m¦�ر������u���X��"���QhHY���ݸ��;�ӳת1�����ma�0-�z���R���v[�n����Eۍ���ٓv�>�>h۷k-��xۯ̎�:�=��ޣ]��;�Y!�n��Y�vc�����oc���+n[��̋�(J�0��&E{F��48߰bW�ʃ��klS�n�K�F��]�'NEx��Hb��Hy�7�K��YI0�cErAB�#��÷��O^Ot;jh�W%.�歼~�w�$6��x�k��L����{�v&z-��#�u=3>�(��%b��s�~�����&��Z���b)P�Νyg���f}f�L[����|�t��S}��uH�E�`,"b�,j�J��Om��{��YȺ�Э���
;e�������gy�����������/>]� ����|��0��8��9e�J��Ӟ/]w �=GcZ�An*��E�2����o?{t�o��-�>���տi�/�7�w%�(�eD�!�^ۓ��A���ݧ�����X�Y��8�{mٲ�M�0䂮�JF����(�u6�1c/'/-��K:��zu'�nz7G{N��Kޭ�g/���LD�+.FP ��O.�۩��S�iw��{��������y@[�C~^( rxԒim��u�
�����י�y����ʽٽ��Ua�<�V5j�����%=3�0��Z~Cӓg7�n>��67S�֡���O"�;�Խ���G"9��H��N>��de��"�{p�iIeMʊ�>ݭ5�JIUo՝�����k�6t}�=-��=�ݾe�Yq��Fۑ߻�Vi��<eͱGׯ_u�qf)���	�U{oL�_^[m׊ܞ�j٨1��.%O����L{�T�\)�܂�d�aˢ���F{6����3�S�5}�S׷�]�W�<f�{�H��_�̆��eWG���[7p�Fm�u�L�p�
D�Y������Ƴ���b�-�L��n~ǷѵJ�BQ��!��i���^�s�~{z�Q@�"Ob�܏WƗ�v{�����OĘ�Z�V���6@���Oϕ	엗�Wg��Y�)Y�Q�|��r�=y��	�$��QnaIs	A��f��&��B���Fe�b�S-����"�C�ؽ�ᯉ=�(�����q.�յ!����gGw�c�]j������]?K��v*�nX��ٷ����l��q��iƝ���f\�WIC��zݘ�w	����K9/��1����n@�^5�U��T�n�fuo���2�Tt�Xa?4�)�CuOӪG[!���(�������{a�d���4+���V������a״V����7�x���^I ۉ�$��N)�qU����;쁿�����UiF���X�}���-8�}�3\�h�y�ӂ�~Ij��������O>�f���j��c@��c�з/l��.[a�-�M=��l���F�� �%�r���7��֗W]��ډƎ?j�W\�wk����DA��Ց�=��m��B����3��O��H�Q!R9�[��x��V��;;�Z���Cn��cy��};�^Y�,�${[���`��A�<���w�d������h����7cy��GA_��1(��v̞�Jm�]ꔥ)���?<{�~x"�1��4��^��HTm������p��:WЮ^��:��������wN�	��zÛ�*���}���Z��JL�Y�ݝ.�	�B訴�y�q��pg�G�T��{�Ryw���8�mr��J�3�ަ3\9��r�9+���}�L£��A2oR	��gM�4��=�ǵk7O}8|��pi�"���:"��yڿUU�eӮXȂ��������ygc,�O1�,c�u�Z���=��ȶ�v;c����*ѹ.�������B�_z����|#ɽ�>Y�d��]Q\ו���-��c�� &>n����=U�D)D[_�t�߱b�&��܏Q�Dd)��+-�ܜn�I�}��=�^�Ti����{�����Ɖk�5,4�D���Ч%�k��5��-v(�gq����J=��W���e����<jЁ����� A�~%���Z� �����%�ɀ���J(�4~���P����]�b�J��e�A�gn��Kۻ�;�U}�J}���.�]D���m����[��+����}]y={]�"�� Dgy�}�uލ<F�CmZ�v���y��b�"�uwr^�6��rW��l�lߜ�쳽�]���-�'N*���{H:]�Uz9YXQXmC
R�.�ٷ<��Z�<��£U����7]rI�}'�흞Ϯc;��R�v��ud�O7���z�6�t��εZn���n|�t]��]���'�v���ݛ���"��u����ܹ�۩�Wc��� �n^\k��f.��ځW�N��g^q��X�Hx�^3[v�va��.�gԂ�ݱ��؊�뚄�p�4F�`�ti�F��M5�۵��ݳ��]������u�X��������n�8=]�+�F��[W��j�V�:�ſ]V;oܧ�W{]#:�c��m�7.��{,���?a��vvP��c��&Đ(�I���P�F3�W�箛~ܺ喽s�B�a�a�K���TD˞�}���mt�+Z������3���&B�
Y�-�	���c�����a��T]�b+NJ �3Ԥ��t����}�ߒ��h@�!j�	>ɻQi���3U����8����g��&���=�����{���j��=��7#Qn^����?G ͩT9���M^���+K��ͧ�p��YW^���	���{|L�f_z5�v�TLf�<*O_T����7�^k�����(�G`=h�v��W���n����Ѱj��s�oB��p\�V=2�P��To�9��}������9�+ڿQ��r]B����m��~����*�6V��f��"M��2�a&S�Ǫ5.4�b��d�֧����q��6�v�����j��I����sy�M�X���;dܻݤ��'���Z�Պ;���_���%�-�*�}�m�vk�Z=,s�O��g�T�0�f?=lu����M�q���*���댈���$@��Z�]���Hr��w}�G~2����^c����vo�b�5�+�9�gӷպz��dћ�p4��En83V�>�z�	�~k�q�]��x��^��W}y�"��U�U�W�is�ɞ��^a�f_	����/n|P�N�,���*y�"<��w��.�����p�.�kGg[�}~��>Mw�c�����Ҽe�<<'�"C��On�Kn9e��:��l&� ��2�$9 �(A���u�Ęv���n�Z��bzg9~~���a�h,�{�1]
w�����N���t)�c[�j����l�Qȭ-{�ػ�у��o3 �hx��'����$������B6}~���T�1H�{MMg`r��{S&l��e�6-���,x_y����\����U�x�?�v�1���j'}���>��mw�3-}.sZ�oӸq��Kp�Otr(i�O5MH-ͮ#�߯23��x�{xGOzI�h���)��]{�U䥮 ä����^E�%4mE ����g�y��2u�Of�Z[���Ju��7Ǳ$]��b���ޞ�`��fO��	y�	��E'o��]~̺�0�lѠ� ��B� ߜ�,�H��O����g����w��2N��j���=��^���G,Ӂ%�`�M�j�O]��2�^v&u��7;[�*p%��%����>I8���K+���s�*���7��48vwfJŁ�ץ\����&�O'���9�߱R��U��\=�)!N����(�H��<�6�OK�]o�SNX*�as�\�2�����_�qf�˶��ǽX,�,����I�i<�gJ�j���&FD�{j�#���dZ��Y���G�U�j���dey�*0(�R$ci"�."���gz��|���8>�?r3T�'���~DWC�Lu��0����ϳ�fV$ɜ�H �-t���]b��u��[!��/�m���"lv]�=�l�h��M�Ӫ�y�)�<���Q�NAr)z�w��Y�:�XZ�
q��H�aMx)oF�7�)����������������(����мN�8-��2=�oe7����uW\Z�l[�ΌdT��m�v�źY@vCE-{�}l=�n������tg�����wmy?Yb��c��XV#���n���e��|wܾB>HS���n
��{g��MO/���J���n�ŗf����'�>�S�ߓI|�1��eH���k�}����!0dF�(��ž��{��fz�MG�k,U���ׂ��ٽ{=cnb�����s0�k�����8��z̅'-���E�������E{��h�$�N��XWL���̏|���D����8��o����ۥ��w�o��fUPb6�
%$��T����زAkl��g��g��vqVױ�_� ��5��FΨ�ߒ����><%p�wكEz)��Uـ�5�
[*��X_]MP4��j�����g	^��㧹����������qm?f�^��4&����v�fi����AǺ�p2ɶ�)��T�މg�5����)��B�3����}wԓ��ni����fWF��X��1�4$��G�A��,R%}����z��]���{e��օ�l��=�9F{E:$��'ַW]�|��[���`����_d���t�����zOR:����ez���`:׍޻��[t��G���ٚ�a^��a<^�d�b�w�7������(���/��^�r����?Vz,N�����8_vOx5����1G��v{xg~$$:��a���K��!�.���Sww4���<�:SV[DMX�8K|/�'a�\`����\�u#%��;�H��[���P�7;{��� -	�HZ������b��g	�p�Okg�Ar}9�g+&�`�~����s����>n��;�'��8��t���\+rk��om�~E-_ZW;&��n�ҧ􊵹r|ᵮ�+��fN_5I��w�л3�a�%/�sys�S�^���-�u��ՙڶ����a�՚�3�%�ev�<���r���&$����X�0|7 �q��澏ܖA��9�}:wR�����U���C��]Fni=c�i_jd�:�gX���*�v^mH��} �Ӝ���s.���D����N����2�g�M��:��%��Nh��'?�b�e�����_nc�\�<�K� �3��|�E�d@&3N�]���n�ukWn�y��v{q�k���緅 �G�;��@U��kpy����ͶL�l��!a;ǵJ=���V+gv�y�ʰ�Ǟ��\��sf�۱ӵm���5[��0���fy�cm�@�{��]E����9�s���l�^3����t[�aG�{a�����;v[�i�[7��3����
T����T�@za�4�2c"���/e|��Z�&�s��5Ns;���y���v ��RV�9������>n�<W�mu�e��禙�����ɐ{9�����޷��s��z�r�6wR����F��m�:�M�8qF���5��\�{vΕD�XЁ�$AQ4լ�(
U��9*˚pF��1�g��c��J��!�����j�u�l��U��n�{.�A�ydSV�n��v�l���� K��8u=�������s����'�^碷���[���R�J6��Lx�78�b��ƃ���7k[�:���=:�&�ݸO<�V�s���5Vׯn�H�&@�E�y��}q/�"m�덗���mm�d�v�9d��mx�v�W)P��4�Q�ڠTV�X���25�r�ݻHr;c�����s�����\�{Q:�l`{DK�Hŵ۵���s���m�67b����ۅ�ڽ��FM��qՎ`8�.�N�oJ/#�H{�'��.�K"�����Ϛ���t���n��m+����އu�R�����cl�E\�m�vի�]�[��콰��Ѭ�9��b�ݷ�6[�ۂ����q����0�ܞ��zxM��Y�oc����j�v�`���#it"i�>�W��g<�^�ܑӻ8	����ۗݡnp�qd����E�������m{s�v��X�c���x��c��������uf%�v{Km�4��ɼpE�����w
�-̻�7�z��3�n�uz��}�k��/�� R�`֋q��rR]��S�М��[�ڋ�<������R�V�;8s��s�c���YƮ� ֣jq(�lty�Y;k��BΎ>@烊kYz\ݎ���mnv�by�c��7N]݋�-dn�]���۠�9��ݴ�]Y���c�`��jA��u�'������jg;h����{n86��d�{PH�u��+(�n+r�ƺ`��^}sZ�1nk.x$���1�1�<�H�g��t�oƹ�'9�8���12�Mc���F,�y�yt7�m��2k��hݲ���Q�5̗Z�<��s�D�dH�7�L �r��np��HV3A����h�~�!���6�V{֝�B�y�#ꩼ�k�z��*{�Q9����B���qh�ަa��,̼��T�k��y���[�R
����g��y~�/U�<,/�/�x����<kY=��.Y,�/�o�;������]ly���&���v���%(咼��|5SU�Gl9P�O���݂���T�3�	��p�D��
tϳ���UD�T#﹜w-q�E>���t����Eۦ�`����Ǎ|�z[��g��Y�(�e��.�i5�n�oa����HDn�Y�c0v�kY܅l�e�y��kDNAM�;��܆��U2�3�E��㽉.ٟp���C>�\e�����C��k�V��UKViq�O�:c��eX��|߹k1�E4Cr��k��G0������v���p��h����G�`T��D=��Բ�+��>�Z����5^�)M-���K����Kdu�L�`��Wn���-m�m�ĽFz�L�����JH�&�[U�uSi�)�=c����1�3�K������f�F���L:���S��s�w��9	�Z�.z�f�e���M��s��Ug����8��!�׌���ϝ�z-��'P�h�������X�6�L8��dN�~S9S�ض��}e��3��NTp�.yr�v���2N�;xGn\�� ���ͩ���ʗK�a6���ň�^6��Ð:/{}��_�w��,~��:K����y[C�D2n�gy�{4�k��NX�N�:�>���K� )��hϯ�͈_r�{������:�{�t�5���'���YSUGd����q���Ҍ���E���̞0��������� N\@��,��_�?�pg��@vnc�k]z����f�'���簿���~��F��#I#����l���I�4��	�5X�׎�M��!/�s�_��:�9m�E4C9p��o���W���y��c��3��3Z%��J�l'����G~�;u�|f5l-�½5�K_���2���k`�k�[|z�TIl%۾�[�*��Ѭ�A��B;�L�)v΅��{��ћ}O�w�1C>����AM��]�賬�w<jݏ�[
t��gۯLc�ƭ�o����2�
�ʇ�^kP3d3ɔ2}p>�[�<+��t���v��5�뱉n�&��]�u�KQU
ܭ�S�[4�ҏ�U�p}���oy��vQ]��[+���KFg9K���c-��zכ�F|�&����O���aK<��0��4s3�u�jXސ�߅�4��|��)5uil�oK�k%�Z a��g��ό����a�Y���S▪`��Ql�䯻��F#Z�>�E5L���B�߻��C�����������d.4V��c��=�H�s�O�6KƖ���	��Dl�JbQ���W�/�]��{�f�m�������rQx�G��W�P��
,��������������-8fP(_e5�A�1�#�{�wg~�+G��=n�;���cPD0z^yAU�i��tKD��(���}�lB$Z~�C�Z#H�Z��^���]p��#y2�;h��ͳ�}H���[f���H�i6sN���=�~�����h�grU�ay�cU��8�����x׹��̀����X��S8���\��;��}c�?�}��Ś�|a-�X�h�O;��?�q�Kr$�i���ǈ��"���߷���q��Wp�h�M���Wg�g�ȴ}��m�v���5�k����v8�"�,9˛~a�9Ϣ���D�]2*J,x�5ƽ�?I~����~2��$s�u��z���v���c��<d�v��gO5U�u��=<r�Wj3�\r�+����ǻ[ܴC2�w�_E�=g|B����,��+�ED�"Z6`���_�ꯢ�f�����?��ߜ�a1�U��Y��d�ҳ����(����~X�?/+!IS��*,�ҏ�zn="�i~x{7�ޖ�}��n�Ǹ���rU2�#չ���SD3���B���v���]�-���~��kv��¹��j��z�5�c�/�}�W�KcdwEl���5��2�o��}9�"яst��ɎP0�?_����DXG�K���ɞ޷9��f�q����G���ˏ{��W��er-k5����Z�\3�Am7����hV�$��)�Wf��cQ6|����zͪ���aԩt�@<�gY�\"Xںϰ�cD5ݙ)��;����u��|�C_\KY�o�Ӈ�矢h��aA��Ϩ[FĨJ�4�����ʛ���gL"p׬E�u��7X�ˑ��2���k}�OyLU��Ρy~v�h��!�&3n������� �r�a
���z]z��� �j�%��w���q�3�M�D��,�UL���������;P�u���nr-�P�|aMSp��^������I�ߜ�5m|�h�ֻ���9�6�̸��F�>�Z��
�j"ofAT���
 c��eP��R�J�ܾ�����2����������[ɐm��ٴc>k���(�,l�V}�s��k9v�Y���{��a�;�\����<�׌%��4e��Z1����ЇH$?���2Bd��B!� �N���S��ƌw�]v��b;��F#��?l��m}�XU�T�;k�����j�9�ь5���S^e=�k=�p���D��6�Κ#���0���G[�T8����1��H_�1G�W�%�����SMETb5��r|d5��8)��G��r��Y楣�Uv���%��?ihƈ6���U/�[G�ܽ�,>��ހ���s&�=9�E�ִFԍ��d"���3�?���f3)�?i�1
?��=��9���S�,��o��>3�����X{�(�I_U)ܾŇ^��SX�P�|f3۞�.��h���v�����6���x(t_f����� u/^��FC�_ ���Z%�d��1:������Z�SDw�-k5�w�}��@��#}�aO,�E�f3�
��?>�W&ý�0�o0�j�z�m_g]��\h�܆?����c��]/.���Ո;��B���n�r�Y.�w�>�Y�c#X��Xwբ�&YE���{��{����d��¡�MT��}Tc�QA}��vڽu�"�r<��Yw/�nq�[�v	�L��~���݁�Xj�.*J���a�x�m�M;Asf�s��	v�r��4Cs�Y;a��gue8�)7[q�u��G�9��q���[n�S��♆�h����>�kp�;��Y:<X��"����X�狶��l�n�-�>ݠ��g�ֳ����n�l=���=����B�y�ɬfIݸO]��{]���p��F�#����K��bZ�r�;k���e{n��=U���ִ�p�h�ї�[�����y���-��D���-~2�yH��t�c����{��}��3�kg;-y���i���:�k�y�v�g��\�گ��r�星x����n1�Iey�����G�_��K���yoL�_#�f�K�\���U9aƾg.�̱��t��kD�a-�>�|�q��E?�ۅ�v�:��S�g�h֌�;��њ�':�594G��������4��m5Q���w�׾�F�y�3�Yp��\�����W÷��F�e@Q�/��T���Kk���U��a��D��V��z퇽�|���oy�*]�[R�e5��#�h��-��G�4�0!������͘K8ן�����5�k���E�a�r�v��P��z�ƈy]�'�v/p�����=L7���៕���Q;]شc>m��j�mS��o� �N#��pW�uY�6@�d@�|�E�XKD�C=�_e�e���2f��h�D>�#\Kv�j޲Y��,)�\e85L>�i��o�d5�B�A͉x�5g�91��������.�����u�����5��[�{vKc�i����f����8���c\丸ܶ�0�Xm5G!�����߾�v�d4�6c����o>�߽]�Fv-�5�4C���~�΀�r�ʇ�<ͳ�i5��� S-���bε��<�o�[ET#������B�"�W�箽cU�F�q����*���G�x�C�~P�ת�vNe�X�ey�|E
�u}E,.]�D���[H�ݜ��؋�D6E�5��ٶ��|����0��Kb�QM�⃫y!���y�h�Vl�g+�x�w��jY,:��@:�iaoZ%�T"���}����\gZ����5�P�8�_�������ʔq�%��R�sK���*��1� -��Q�����!�}��~���e�-LU^��U6w�Z:�ٖ�g���Ϗ��-� 7 �p|�#�o�o!O!���z�w���~y�5)$����p��ֺ2�2�f�o�ӏ�������Q��v�aO�:��o`o�}�v����ŴS���[D������r[�9�!��sܭ~k�T-����y8\B־;�oty9=߿��_���+�IWI3Ӭ��O"]�SD5o}�p��;p���2��?O'�O�'�G��s��G!���n�-��Q��CD���_��5�=����A�Z.��dc����7����3���'KX�bl�ɡ (�7=�j��2\y��S��X�9�qnқ��k�۩,�[	_�����^����Z���ݾ3�y���
ٍ\\��Y���ܛ����E��P�ք,�n��,�h��x���q�q���;h�}�;&HX�ۀ�?�z_������:[L���b�=�
 ;�$�ߕ�4��.�<�s}Y�M����gs����!��Z�7W��a}�;�k}j�O�;pQm���ecF�ϣ9s5�Z�d�W���� �v	�ҩ_4�􇯚�u�2Y����ƈh�m��NA�g{�;F{�;~t��F��ü�������	nS�[D+��V�Z�ّQ�0l��)v�)��Az4�n�<ol�N�����,Rt�Ol]i�0jctj.��~ ~=��TN/�=��*~���?�KD�C�d�ﾈ���v�RK�,���>c�)��o���N�H��^U|��k��G�􈶊��]�M�K�oٴnB5����l�}͘h��C]~�h�>L����ow�vp1�='F��Z��J����`����H��F�aʄ\��r�v�=_a0iG����{o�"͙Y��*��S���fnNy��m�*%�t�&\#}w�b�b5��)��3��m}��KX��G־��#��<����2�VaWl=m�:�8�R�g�U#�87��n�g�G:����ꍥ��[�x�~�jf����]����?�Q;$�!�:�)�g���ɼk���-�!���e��k̚�ڶK�
|��	����כ����O���!�Զ�y���k�z̻f�z�՜���3IE�ȥ��e��C�_�"=!�D�E���#kX�T���-q[��fT6�᝸1��U#3e�ɁS�]�����CY�M��FUo��x�h�^C�}�kT���V�|<~� X�+qF��7R*�a�<��Զ�A!�?o�I �����q�s�������K�+�W��k��L�X��/{dkG.-�5��mc�����Y'�:ѿ}|�����W�Y�~�O���Q4�Pp����'���F#����wr� �2n�d�Jl��8����F��.���<�^5]7�Flֿ�қ�oދG!�&��?������y3(�6w��X�\%NT�o�-j�z�3\5Օ���[8$Y��U���&�_Gʴ�v̫3����m��}�'��*�џ[�3�}��"�*�Ռ���ӹ'��ϓt�&�|j�MQl)�e�{�F�m�d���O�����9S���q};��4C�����-����,Ƹ�up|�a�F�_^��,�0��Mp�~�P���W{�U&ձ�N�n�f�n�xnq�m�4[.�82#�q���q�S'CYp��svܦ�{�����=�s�G�)��j��͸�0�#�)��E�!�ײ��\3�����Zd�N}��}�������ם� �����Hc<kY��=6q�3�IQ��c1�=���s_����D�q�5KK^%�ƶ�!G���}�%�Y�o3�\�|���g!o���d?���j�Ɖk�"`�z����~�Չni��Q�:H���Tf����̵?~�G[5�����o颰��mo��Yt�,��׽.=^n+h���[��'4���2�[Eǹ �w��k���tIY�~6��������kR�ru�=�]�>5,m��Xy�}Y��9>��G��E3YL:߳߿~�D�-A�>G��1G��}e�}\�n�+�؎mu�1��(h�p�h�{�Xc��E3�ݸ�E�a�O�P������V��媍O߅��D3���ȳk$�|���-��
h����>���:=״������;�e�z��-C1�L*h��aہ�<��|]�{�Qo��2뒋k��>�E�s����� �[1��h��Ϲ\�3Xc���\�5����>����¦g価O�~ɀ�q��.Y��U���蓃3x�9���mk9//xѱ���Ө�ok�g��!@��x$��v�]�Ǹ��	�sm�l��4�(����:wY�'\nݐ͘��5v6̭���Ōs\���G�m��Y��s�/�����Ѕ�v���y��.����V(n�cr�tM��n;2��ez��`�`�9�b�/O+��v��۷�҇��d:�[����`�Skn������Vj;v��VYx�툽�x�[�6�m�L���d�D�"���%S[� ˩u�����ۙ��Nxn7t��9��b��P�v��ng�R.������=�>��E>��Ó����8�jY橢Fk_}�q�.6W-}p[E9��n��j]{�9�F�:�j\�c_:�{��k�k,ܘan��[�DA�wOKp:�;YKK^����j4�N��Wf�_&��hi&"�����V�_}���I�)���=���^^�эK%����̯����:�O�	k���Mn{�,���4vEX����!���������D�T�u�A�z�^z�U�ULiWǦ����7��/��Ý̥��|�f�vݣt�KSw��>o��L>��TkGn7�Î����n��a6�����C�^M^hw?3�DF�ѪJ�%�`y�]��W��|�?r$�u�3��w��eԜ��<p�e�߷>v��o��e���l������aU�ݽaMQ�/���h��	k�Yن���B?	M(�`��������b%�Ka]��aOZ�S���ҭ�
g��hֈa�,>yp_2�c���ϝ��}�KT��a �z��Z~�⅑���_�k��<��-���/�HƦ��m��������	m0��FӃU��D�Vx�W;F�AA�+ovon!;y8i�s���)���&
p������t�e����fL�*���ދ�}��k��Yz�z��:���ᾶ��{�~~k�Mvc�Z"��V�����h���!�U�����
f�0�p��H��KE�T�8�h�����X��:z���Yn��v��pza���E�Wo�k�{��ևc8:CU�|�k��a��|2�4�M��.w�C{�����"A��<*�]������ed.f^ţ��E5��P�k�?�~���D�C9h�}�����p0��k�����Q-_c�ڂ=co�$�q�	"G�3W��Y��S�S���شk"`떌�.���,�92?~��_?C� ��\0�$�c��8q��^>5�����ֵ��N�����a�kDC�l%��IMth�U���P�R�݃�ս-����K*�w���4� ��.�����qT��.����\��0�k������ڧ�;��b��h�FAL=����y�g:�W����h�ԯ2��ST�g��2�ji�E�Z�d��m|ͨF}�ih�g�O�3�Z�O<w������3����m�5��k�4S�OHlVk��gϮ�7S�o�zq��˺�f3�zV�W^����K��߸��M��yO�:���F��#z#�ҸWi�;�����v�V����Q�k��3�6�oK��ůQg�4��ε��vղ�7,>�u�\٭k=�������[.az=�C���_a��=�0?v�*u��7v������Z��<al�,���6u�4TT����������B�9m3K|5�ߤp�Ɗ?3D�vʥ@Cچ�,�߾�uu�5�AS*{+s��m�"Y�_��Ǐ��N<��;��KD4d�6�=���#��^#��w���#�~z��|g����B�*0c%��ϸ��<~�ֽz�L)�Y��>3=��F���ϯ�h�}�E��s��s�؇F��N<�/,��BV����8	�#;v"���ﵥ=�UM�G�2#K��G�Zc|�/!��6�R�2ui�c0B�;�=�m�7����1��{4�Q�ur\ư��.��zY����殛�ә^�M��.�r趯�85�es_f����k5vuR�����a���g����gd䇦C�n��/Cٛ9�f3
�<�5.��q��|�L��v�1ݜ;�z#+jу�FC:�f�CԌ�1��I���ݳv� ֻ�s��,N��ӕ��nu]�u�We���B�|sj�܁&�\���$��j]u=[w8�S�zz<4|D�z@��3��zQ�{u"�ok��a[#}HU$��]�+�[d�ٖ�)��ړpK�4g�����4����X��C�q�^��w���'VIo�s�����h�/x�;D�eOӻ͓x��n��iݢr��7K����t��E�Z!:��Z؇s��y��8�6��ݡ���ҍ����[{��b�r�T�[�����77N1�^
{J��N:��yVǴl=�2#�J�-Lϥ�&�P������b�
['2�=��gM��7!��t�����a�M��6��v�D��D�� [q�)�R2-U�\[h�9�}"�3ޣ�4'w�s\��J��,У�E�u��E��7pк�1۰vq�_ֶܵ���n]=�n%��R���rR��8�˶�n�D#ϭ0��1��G$�)��=�v�C�'f��J�_i���f���>�Ug&��k��[l���kG=�<��!h�O�y�׳bMa��lA�j5kq�ey�5��Z�K~�S���Y���w�-d���B9��"�f�݋GzvQO�\�a�X]�\v1���
a�<w�}Yg#-�8O|�S��YwS�k!��"��7�U{9\�luQ�2YW4���J=!���~߿}g1�V2�����mMgo����p�e�|n�"Ϙ�����-�z�h���ҳ�
?�dB0����������+�x���m���q߶��
�ݰa��=�m��)�Pgc6�I�s��w�E��۝b�3����xx��������n�KG}��c'&U4l�����о�ߢ�ƈk-�`;�~�«�s��]�vYMc݀��%�湻�E�}
�9�N��5�� Ǝ_�f=4D9%GQG�0�?d_�~��~��ȒQ]�D��n��~d^Wm|;W�w�irÛ���D�����E�:ο:r�D���h߳�_^w�,����yݥ_���#	�O�|;č�(��n�Qf��W2�-��c�>���k5�tћ��9�.}��Z3bX6ٟWy�qw>�O�c_3������a7�O����<~k�Q|�'v>�U�m����K��~�؎���U�J��k�����~�a�]���V�&~�-��,�>l"���g��O%Ө%�j�=�Ϣ�y<�4K�y��.w���E~�ѼE	h:~s�� t�a��1�g�\횶��5ܷ�'8I�����ܶC_��i�H�[��h�g�L�=&�`�bG@ni�����~[�(e���6������CҼ�����#�"�!���ֺ�-�jXS��ߝ�Gݕ�p�g;�l���R�W���w`�:�!u��>�[��~�d3*5�k��k&��q�{��~q�+��a,Ǫ����-�e�a�߀����Q�!��KU�6LY��g���ínt!��k�pv�;����Y�i7~w����"w'ߟ�汄�m��}�a.Z$h�w�����ʅӱL-���L�m�$���Wr'g��f{+yM|�:a��}m[>����Ƕ�#nwdƍ��>)��t�e��� ��#�;�@�ӄD'λ��Z5�;��TN�¸���墙��Gs�-y��E4CD7�r�}qh�r�0��]1���lY�l��}D��8u3}|4�#���j�g�a�m�
A�$�4Y�(�~�����ϝ�=g���Ǝ�"YS�R��}v[W��C-������J���l��>j����܋Ƨ��3̖���a^Q�k���Wе����;pϽ�O/}�D�n\fH�EI|,��@fz�R�۪�z
k��ٯw��1g��ֵ�6L�B���K��Z%�w�^z�cz�3����}������D_��~�i����;�#Mc=��z�s �6�ų�OT�iĶT�US�kU�ߘc��[<�����㸅M�yqɹ�>ߠ�W�5�Ïoޯ�kT�aN�5������h���e�g2��wnZƍ*����1�\���5�;��>@�9��3}^���sx�Ǜ��3��o0�:6�{�V�Ua�k]��V#�R+���i��m���<�a�u�  V���t[�6I��<�nz,�+�nyr7�q8c]�lk�9:�Q�8�˗��z�pl�؇��2��C���A�㖹�m@�<� x{�lݕܽhuɼ��Z�ع���W&%�����zS�������\�[��wk�n����5�7c�r����\Amǎ�v�7X��NI�喻T�(�=��f��}��R�%�� 	0�+\��I�����k�<v	�ݲd�KX���խ�E*��
�uB���\�Oi��� ַ"�|���^In���F0��]��=y�V��f�-��j����v ���e4K�7Yﻜ,9���-��9���Y։`�3�r+{6���ˤ[S��[EW�<�·FT!�Sz\z��Ү`�h�����h�w�F����kD���)�k�}�����Pk���1�j��X|��g)D?a���������!�_�����/G��"�G���`�&�	8c�jG3F�Z�v!�3�w�.c)��cE�|L���ɳZc\t�?Mo�UU{��N�h���nE�!�r$)�*-�'�ae��>x}�SV�z�m����
K`��(�JE��|F����k���Y�|I�V�=�o��[{����f���\d5=���`|�J�NږSD��H{������\��K���D^�eT.��벚�D�a-�������ģj2b�$wDap�߱��-��5h����|�?�މ�<�iKo�O����o'<w�����W���SE<��|ϝ��8>����ڱ�a$8��W���1�?�\���AM��vc&��ϑI	* �;P���i�7%Z��� �'����vǞ��N��F䛳�k��Oim��_����xƿ3�/~v��`հ������2o>�D��3�ֆ��_��~v^g7�Z��nQ��ϯ�g���h�_݋.�_1�{�j�C_��f/������Jݴb1�d�-���ao�߽�ew�#F���2��g�t,��H	#[�{<[�{�ӗ�ú'�y���)F���9f.uv�ڝwh�m]�����CCvV��~�A�#���R����Z�N��)�ղ_�G���1�KD�s�{6*z�4<�ݾ�=�{���������&jF����f�lFUAL�MF#Z�KD�r����7��qd�;h²Kj���s�Բ�<�[O~������־g]�>j{��g���m�4r`!�P����^<��8�!q��u�6�彧��!��F�am3[f����fNF�|�#�羸��[\y��ϰ��q��+h����m���p�=k�限U�!�׫~�l=��E=���[3���iޑ����;��Y�6��Z��,��C�����h��l��X�SU�JF�i\��ŝm�~�>�������]]{�\}�,�U͇_;�L�Al�yÖ����8�j�a�@F�m��g�,�̨h�ˤ[]�5�.�����1ךo�m�܆`)Ȓ%Q���`G�����;����s"c��s׮r�"ZaB���I��#;�?����k^���Z8�.U�g�
=~�,ƽ�E;f����+~�T�a',��S�4cD4va����Z==����~j�)�y�������l��q��0맬�-�c�/�N)~|dl��U\�r'T�Os)�+6����GZ=1�8��
v���צ�}=a���q�ZF6|B=���g������{X_y�ǯ�{#3���j[Ke-d�x�h��f5,<��E��Z%�身aO�=�m�F>:ct4���}L�fy̏��c4��dn�ڣB�H\��!�a3NsC ^'�9�uv��9��\gm��5`�G<ě.Ьf,���Me�}7�o�u��!���YOo�8t�]h���d4w��6�)�Q+-�E�ޗ�r/�4������䷄��6�Ǿ�;F3�
�|��c�Z5��L;vAY}�ѲH��eA?C�GH6+ﾜh��	k=G��ي����ٛ�=}pw~��8�4z/n��V��y�������)%��-3K�^j>��\w:e��di��sh�y�)�kV@�G�}��q���� w��q���p�0��{��a�zz���T�g��;�^��>�"Z�%�vh۲�{~�����7�;�1��9^& �a��\Zg��f��:�v�ŀ���c�׵�-ۛ&� eTn�=���'�(�5Z�.a���fq��K�6���C=�Y��p�frU����oX[�߷�k�wry�LG7��G�ΙL�,=W����
.���%�0���˻t����e��y�5s�"��L����W'�q���.?}�7-�U�G�h��\��k�kD5��-����N>�}c=�x�x� �5++�E��4=y��E�@�Y]�[���"�7%����_a�������y�Op�p�~��adZ��(���ش=�CU]���]gHh�<9>kw�ٳ�"K��@[	��N�#��X�S^z�X��E[j�-� m|��d�[jG@"ձ��[�(��-���<�~��-�jXk���Pe����mm"Z�8)���k����5����$xݑ�v^�)��������!u��ڟͭX��6����T"viұ.�Υ��P�X�KY�4΍g�����lS����Sk�}I�����	]h�B+.V��(�� {#��T:��e��f�����-���X�K����c�ZG�� 3�dPX.�����=!��T��S��	���7=����E�h%��}��k�P4h��,�
������%/��T�܉���n���:����s���q�+���y���c��珼�ѹ���z�j���;���)�:z��!Ǿ��F���J\���E�z~�f��ֺ�k̦[l�����w9��6�;0��ןj-�k;��_����"�Єo�B�å��ߛQ�
%�4�W4���oH�ҍ,繏>�����sx.k�t*�Z�~�{�@��˦q���E��]����kV�\(e8a�s'�k^����m>���q��2��qx�ެ�+gvMs��tL�T������4�=G^���=q蟹�E�f�Ȩ�N_�r��__���5��﷘�W_i։v��^;Z��E;t�0ڋh��}�a܅Ƈ���q�v-��Y����~``�ꍩmv��u�k������!�ϥ�q���VM�;0�T/�L��W��p����F5' ��������l�t�OZ-������D����wվ��Ƶ�k�t�zA��T0�?_�q_��$�E�V�5^���������Mn�)������~����v�,�A��W�ƾ�Ì�O�ʠ��݋z�/XKD�<���L�Z?"!ȇH����k3������̳�����rtia#�;l��Ӿng@���v\�{"৻(�뒯(z������t+�s��l��0�g�k'#D�'�Bf����c�烨�i��u։��`�����_}��k�g9hX�fظ��f���/Z(�
��OfÞηg��SmΔ��1s�,Oj����+ټ��q�\��g�pV�n��	ͻ��{8̈́�W�j����R	���77��	��	(2ڹ�5��8��N^mgwMRv네1��l`6-�B�-t����	Djҙ��_k���<s�vÞL/h��rv��۵�WUmgo�.��vSe����=}��)�k����W��F���J���nQ,��mS>��E�~�ԋa=��	r�Ȧ�{���3sg�8O~�;���!�@~�V}P�cw��E��Z)�d��SG7�c ��j�UW-���ך��J���%��g]f�ʛG���v=d|w�.���\�ݺ��=�v�4C\d�9�ZsϽ�`w��%�P���v�ٿ}fB�Y��R�|�n����¦�A�5J&f%���)��D�C��)�����V�%�ת�l�N���R�h����󜿉6����od>�*�ѭ�k�����nUͣ-nS����О�w��hD�H6a*��~G��[��fL����t!�y���1���S��rSN��o�h�O��-�
���N�q��w�����{�=�Usq�4o׻WO�7�y���� ~�����H��&���8<~�������[��Bƈ��󵣧��¼�axM0l�Qw����qE{�;G9�E5;���M��s&3�7N��ZƱ��r�~��XKֈ��"�D9h��!'&&����~�}ʯZ9ON2�|�-ӽ���N�����wt�9���n{��W�NR��^�����k��]�C>��"э��Ϯ��m���}�Z+�O�[�e�J�]f>�y?az������ɗ����� )����ƾv�{��gг��FN0���ָ����N�P�1ҫ�oK�AL1ۦ���_�a�������c�l�m����r�u)��mC������8�w#Ψh!&n<�x��{s���Dns���ߊ9Ǒcn���s͟)a����+�ܴJ�G������g,�3�~�w��:@l�yV��^X~�5㠏�C?~�S���K��w�z�������d�r�*���-������`��ao��0��_��jvj�,˔r�s~�﷼v�v,�[���}�ɒ�}����:���~��]�x�o�)��y�ӟ��/!6����Wp[-�,Sʪ�ʊ&I���>kZ����;:t�f�����,R���_����y�G'��gz�6ϣ�\ٌ���[�u��N}�ۿ��C�l��ܰ�6flrۅ<���3����#��_T5W
y�Lis�Ϩ@���SЪl��ޛCK�;�e��Gܪ�mq�x�뺆n�>.,N��?������V_*�A������ly������Yn��#]c )�հ�#3��m�=����V�^g������9~�J���kJ8�+n8��_m��:�m
Aє�������;.���2�ł�~�#�<�~�E��?G�t�̨T�Mk�S]���?{�y�c_r)�	v��w;ذ��[�v���/�Y���� -��ږr�h֞B#ܐ�mO Ƌ3�?JsU$9Q#�4��V�9h��ԏd��ϗ�����xδe���?e�%Ns����K]ڑ�S�z�ȿ��}h�����Ӌ�F{7��kF|�!���;W
��L�T�z�9|��YuP�(��.io���^����c��9�2�����&�r���������D?9?x@��UT��'~��M!�0a��2�"� .�J�cl��������oE����3oJ)>�f�nc3	�{ʨ_���$�49j�o����r�2Y�a��o~�e���-��T5�4W�ﰦȊU52'$U��j�I�u�_�
�|�0�6^}��jYӰ9�Mg�Jl~��u���d���1����!�ӟ}�r8�OK�o|�*�eD���D�}�Y�p��ª�턴Y13����z_{�[���M�c�ҍ+�ɞVy�f�&ўܤ[9ߎ\l��sm�r������Y-kt�-�k����X���f2�k���׿FB�E3��@D���w���8���#�̫�Sm���d�|�=�ڊ8n��ۑyu�3�gs�۞;vx���s��i��w��f���0���KF��vz�h˄K>i�o�h�'i���'d��a/��7ƪ���9����g�I��,�����w�^>�q�ܬ���C���ߨ3�}��P:�␶qy�<*��G�^4�K�͝ߞ#Y1U��l��w�X�g!�������ͨg�e|�j��/"c��������֊e5ʀ��8���p����ׇf9l����ڱ���=��O��Q*S�&&�QǬ���E�h���������V#Y<̥���V�r��;�<�qGO������������;�������u��0���������Ϯl݅ǥ��cK����߿-����&Z�sU8kl�V}�cFdi�9��r3C�:��|�^dl��T"]�����Ѭ�R�ʄK����k�־�7�G� �
"q�۴ך���Y����eS-d�3��4_�z�&�o���F�1�qr�^k}�&^���j�ΧU�����i]�q1��=,v�@j�~/�!��{XkZѦ�Q�X�H����G���jLj��j�)����\k�s�,���g���83R�-���{K�ޭ��������F9g.a.�#�_v0>��D:aڂϹ:�j~�w��C��6!�_�"� p����e��sq~�SnH7@�t�E��k�����r]�q�^N�5�����ٚ�j0�v�S��;�����ݰ���9���mq�8Ϯ5�[��S뛅���6�Ǽ�jݵ߈��[�͍i�}�a��}���<��ϣ	k�gbr��l�_�����
j��a����/�-BD�7���<y Y�L�
��Y*�]��n���?r�tq�����d5�}�v�r��
O�)Ӷ��߻y����f�j����E��w�]��ږ�7����C��H;����r-��ɟ�G ��67+rJ����ʃ����m{>س��c�}6!Zz�4+8��F��p����&�������Q�w�^�c:�0���a��D�ϻA��t���֍�������Z�����6�f����b��6��N��Kg�3�"����.�=U��@:�N���}j�)�70���~�8�zB�S\e4K�@zo���=Y��A��~��q�w�d���sq������E�C���t��A�Ӭ��[3]o�_�޵��,=$doܛmu�o��f4[_D�+>��W;Ϣ�ø�(�l�D�aݾ�����5��la-�����/�ֈ��}0�O�5g��ܽ�Fd]��v�C2�U����hFe]"72@��L�����ls&�U�Q�~m૆<s7�)ݗ�C޷�V�C�t�V�sm�^em��贬P��D����#��c�v��ײ1�oS�(v`D��b��nɾ3ˏo����Y5�����1�D�����t�.�������Ww�P�rBU��_�q��XN�Λ8�	'�Q-�aJ��n��k��*����r^ay�Е{6B��1� �:��R�R���v��c�lAu� 톎���q��]R��:��x�������h��p7 r�p�ᕙ{�����!���2��y�{�ʒڏ�a��ҵ�I����3)���]���sw�n����+�t�7�G��`�v�l���ۙۦntw�j��W#����y*�&�v��v�[�i
X�W��0��|�H3��]|���Q���s�e���Ө�	�bٹ��d.���\�1h�1�����#����s��}��j�Gc��PLࡔ�fV�r���0Z�N�>�S#���o����f.�&��)o]���"nR:u9OxEpu.�,O�(ʜ�AY��\�GD\�E���d�2�q�I�t�է�F<>󯔛Ǟ����ح��
Ґ�h��X���3��uٜm�nOv��d�|�������1#|tJ�z&�nx2�ݠ:������{u��u���ۓfye���v�w��$^P̭\��^���X+����v8��t���S`�h�e�b��}���6��$s|S�1�wzd���c�����7V�� �v�ӐA�u�{fn=���9����a{�c���UV��R;b
F9$�m��Ml�4f\�N�O.�`��v�:�Gi^~w�u�l�G�Nv�3ٱrq�;�z��/O+�q�3��=v���8��oX�v�:�O��w<�3���ݮ[�.5v�_��f��Gs!�;��*y��nqy�xnC���q{���+��;�;^�;���P����cvy�;[eN���ݬ��jwjM��a�T#0������q��Fv����94�nwZΆ{vݦ}��ó�{`۬u(��=���<T�Hj�]��Utџ����Z4O>�&�p{upv�kv���M�m�=n3�C�P��cpcq��u��6xۀdD�������Q-���؝���g�.�e�q�Ǳ�ۇ6���B�W�x;�ez�AI�Hs��}��.B��p��E���X|s�*�Ȼ���˸�݂8�c���7i����C��Ńɲqҭǭ��۱�n���`n�y1�u�b�X�1]Vgu΋����������l�=�<d.Qmd���u��m��W��9vrqnk&9�n<�v	Q�q��˧��u'n�0=�\��n�4m$lm�i.�����޺�6�;��.#��w�q�8&s筈����
���8ψ�e뱸s��	�2s�.#���+�':�\6���U�J�:�a.�,��M��[&�9|��ܶe��w
��;,\�74歶u\@��sG�[a�e���J��a�)űMU,�"HWG�5&L2̸�U9w�O4���rh���g�����wi�;7�m��9;a�[d:.T���`�rל�%Ix6� �#P�bY�>�WKƷ*	�l=�G ���͞����[[n�v-�!Ʃ7O8z�;�u�0�m�m�gs��j�ؤ�;�s׷ur/h�:L
/\�ys�nY�;��<F�DMuq�9�-D�ͧo���ݸϪ�%<�s�۷E��z��s,{�K˖�Ƴs����[����6�@<��^�LC��\��������u���m�W�V��0�v���x9Ìmmˣ���c���v��wh,3ձѺ��-��9[���G;,㇬�j..�=��`�v�9we�g�>#m�uѕ�a��=�:�;F���m�3��{I��#�n�q��n�۠N\��;��w/��]���ܼ݃���Wcz�;��ѳ���ZM�Ǝ9��v-�>���j��G1�wLc�9r&�6{i�=�)s�7[-��7g�m��2*Z8���R����\z�󂚶[�
k񗻿~F��,�����[>j���z��C	e��ɍ���_}��t��g���?��4cD4CGn����G��L���G���+`�2Ie��eٚ��8k�L4����5^���ы��=�Ys+�V0�܄S>ٜx����Գ��zԳ�)�Z7+�E���6���ݐǯ���G����E���[�G����Lzg>��}��S�!�1����_�L����Q�?[@�4ӽ�j�5o��}6�z����=:�Î_��e~U��ek�g�2��?O+\9W�O�@}��;m�ﾟ�-�^��x�W�ig��Y�׵q��R��� ԭ�K3]k�_xX�����~x���"��0��uo�o���S���Iju�h_"Gq��>�آ2V܇<+,,��<�J �U�m��D;q�@�C��s�����{әHm�����;�^g5��j?9��!��I����ڗ0���~�/>rE�O]IIY#���Mv�Y� x�۴[�� ��=(8��9ގ��Ѱ�01)'z
�J�ͮ^����I�����L��_�S���}��A=t�=���R�	��!{�,�I" ?	��c�h>�����&�%M����1�N�ޟ���j^�K����}�Y�N&��D2.��\FGz{j.b )|�nJ_7��=�e�"у�7��'
QW:���ii�U'�)��{�����c���Z���\kw��}2(��xV�#�HZL.��e�N<��!K����~ʔ�5r���W�Qރ�<��Y�Y:�.�Fa�^󬍆*9���Es'��
(� �w�[^{��/�ܶ�S�n�f�^P�i�+���z+�^�Ĩ� <q@�����^��}�k��T���l0��"G$��ϩ$�>��\�~XAI.ڊA�d�}�}MWt���R����װ������-ۦ�S��W�=6PS�2P�E&�07��ǧ����nѸ�Y㧰xy�׷�:��
�&_P�bq0ā�$<=0����+�j^����l��#P����ۆ괪.�)�{�ϜҠր;����w�|�#Y �Oђ�y��6�{���W4o�U�~��՞�>�>��n��ߗ�f��=veKf_��{`z��cj�VclOY>*@bp%��e=�{�r��V���n?el}���>�����@�C�Y}��k���^�	��c��0^ε�xm^� �V�#�0p�ǟK�<��V����_M�x���:eU��{ �t��N噡�Otj����o��6��i�=�`�t��ȢrnsZ��)����Z�gN�H�ߺ_����6�]2���-��v9�,U�e����pF[1$4�(��o��^e�Ǎ����R��6�mxIckFv������(���)E��瑷ߗ׏7��%��)�����#�ģ����:i��9��cn89�᳻F��{��9 ,��jGܼڿJя�}�R�jJB���>������U���9l�&Ĺ�F1ejn�k��w�:8}��*!��
5"�mpOٕ��[��*w~���)�9��7�L�SZ�T^�7W�$��w��o05}tkvf®Ew���h����2�n>��&s�ag�Ɨ���\�~�:m����g�w�&�s��.�����q��fF!!�3會m��� �(&����Nu�/uB��ZͨA�AOut,�Yj��ܮ�����U�1��B&*�<�"�}�Ԙ����G��\�������4x�3�u��K�bX1n#w�qНX2�P��<*{�d��Kv9��W�Ϥ�cU�����iߙ�d_@w��d���0�콦:D����x�E��,�yx-.fz�����X�-N+r�l^O����󆴛퀉2���f8�<��6�lA�:�qy�[m���9	�y+�n<23��h��<�~,_��vj��W��J�h�{ͮ��e�W���)#����r	�Sw�$C%�C)����ԕd��x�4�y��_[��g�x�Fe�|�ߓ����u�k��_��\��n񺙙:j���~N��Ď9�!"�׾󫼏���z�˵[�v8�k��5���h���u�������e}�|��RC(F�������z��E%�����~�?a�<nz[���!$t�஽�+f�Wޭ�Y��y��A��M���%|y>(I!6���s:���a�U-׬���VM8��TSW_�����K�>XN�r�8�ŭOqx�4���Ş2�i�H/���SS�ЧQn�l����e�ܹRk1�ɻ����95�t�P�k{�uwf���p܂qA�+ 'i��X��[�m�Q�n�S��Wn�k��({[`��n��ͳȞ�r�������<�9z����n7���Sc:^G=q<���C��Kq'`^.0�s��뎸3m'e�M�X����뫳�eܷ�z��̸(�;,�z��n"����B��"���V���ŗ8�(c�\��ΐCn�z�j�����̼�^�grd AT#mB�X��*Q;p�Qlt�ɶ7�h�7`�8�<��ɇ@qs����Hڑ��Z�*�S�a#���鈩��y����w�X��o�YY��O?��e��}Ml��_&}Pa���7ج`�4ڒ@�rA�^��S�{&p��}]&x��&j�#RJ�^�=�O��z��,ɒ��{*������@�17��$Ja$���<����S%�{5�j���${��u������3����Xg�r��Ȑ�!!0b���N����8JF���|4}���vn��be�ޕ�t�Ջ���kL#8o�os练.��ŗ<o��2FZ
ժ��7��}-�;y�6��nEޞ~�ܦX~y^|�-ؘ�c��s�坔�W�'�r����v���?��v.T�l�u�a^{�B�!R�,W5����x9�x(�yZ����ӵYG���W[3��e{ΰY��Ǹ�S��_������;T�)�ȝ���2^e����::Zլ�KY;+on�5���l.��>q熶A���.��[���`O.j�p������u2�\q�b�̣�+�Ӌ�*1ܢ��Fm���k�t�B�<,��>�3��_AZe�?�u���e�`���<���,u���7��?vYgET���kvI�QYi���S/=�ꚱ��K�x)�K���־���C >��ՇLV+�ԶZ*u5���o�P7����x~�`?*#)x�ݵ���Z!E��R)g;i��N��l��~�k�]�������l�"%�����$�!SFT�w�m7��[�Vq{<�����6<_�߬6����NHn�04��d"���Y4�9�h��^{z���jT}�?B>�=b�d��|I{�l�	W��mճ���ʐ��}���a���q�q��_Z�C�g�Ƶ	n�ϖóe�mm�2�.���rލؖv�M����vH+���Y�x���O�Қ8�G���V�r
S��ypQ�ZVa�F��E:Y���^���e��N+5��X����H�W�>��r�@�u���������*<6@"�y��y��{�=F�_
z��|(������(��0d������>���ՙWU�(W��:��({{�
���ėb^S�7}u"��ݧ��y!����,�Q�xq����C�h�5��g�_]�>����w�d��+��L5z�TK�;�JCG�PׄEWVg���� �Pdp��(��}fӒK�,���w��g$4~]�I�yrP�9
<��}�o>۷W�����X�Q\~�'Z�4J{sg
�����.��h��w����艁���I(]�F��������d��x����;{��x�U�v�+�ޔ0Z��Zf�}�Ê��<��o9�oL?̑�	dT�7.���v�3Sj�;����=���;y��۲v��,@�m��.��JM�Rzx��A4�'����M���W�F�.���2�\������z�;�V6==��C�ќ��������dU�ýzY��	�s}��O�7�r�Vh�@[1��i܁���tm2�_�&:��!���=3,��K!�x��դ0Gn���ۄ��-'>mH��dFޕޙ/�����Z׆c�,uy{��wyj���޴_���ܬʼt�Ō�B�=0����߂'�	p"a7%�������E�u.Ӿ��H�{�V����������mbR,XNd�-��	�	��Cr�f���(�x&w�*%}y���͖8���YJ��v�ő�+ʇ,��� ���#B\�,�m���+��!�>6ʶ��n)i�����$�.ew�vS���h?-��o�n�7�yz�H���ơ�f��KJ���R$�n{���c���ߞ�	�B4����U�Ӎ\I�^��])^=�v��ܰ�^a�u��j(�"$E2#E�]g=o��O�voq�+Lp�^!+{ҭk	�C��̯,��i����5e@�V ����^�;�����/F�.�f�Dϑ����ݙF,���(�.s~��o��h�d�*��ݝ#c�������z��	�j��__�)>�A��$FD�$�[lA1t���Ꞡj��I�{��M���9�ʇ{۳׭��3����&�s@�O�G�NS�B��dBٍ�w~���^�����_�X���L��3ٞܞ��}�Q�w�y���-}Y���5��<=���˘ʙ��N]W���k��5����,/KSGP�rR�i0�d\3��݁���ӽ=D*hQ���:>삔�̵��3돏	�q�&�~̳A���=o�9����r�]�~c�����wæ��V��xp�l��:�`V��tSnIa�t�oQ���o�{)$��6�!�3��sX=��O\O^e����.�jxϝjf8�7n��u��{b9�tv���v�U�g����4m���q�������8���\Gp>+�Rmm�=�O`<��(�cE���,hɓyN;nX׭�Ϡz��6P�p�Wm�Mu���ppO������3�l[%F��p�Q����n�f2�>ݭї==F�x�sj�j]1PDj��u	���ƅP�}��� =�!cZ��۵E��r���y��Ւm�Y��~��ƿ;��U�j�ݎ�P������t�}㴾�s�纂���B�-��U�D�[��~��)P�SJ��;��JKy��\k�+>��l?f�^��?eAy��[+�w�T�����}H�N e������Y�mo=��\��%���f���,��H�C8/����g
�יc\.6z��r��7�7E���N�d4���Ҥ�
(u�G�;�]	E>�X�|����+�]+%����$ `�M����*���Z��OR��b��'����q1/�.��+��ݒn�p�����*�u�G����'�y��~q��LE$��C�;*�4���^^eY�`ap�Vx!Y%�t���*��W��s�k������WΥyڴE�?�&���?��=�k��ZH�|��:�3v�q`�����¾]q�R�=i�ݝ��=�m�/7q@F�p�b���W�1 qۡ(��bv��v�"LQ��u\��O��z������<�X���x��^=����������%ii�C*���~՗@�C��x��������üW��&�w�[��්�5%q����:K���w]�q����U�Et�����A׸+�5�b�Y���+����,����f ���Q�h@>�d�j�����=�c�;��*2�.{�0��|~'�}��:�Ymޱ��XҰQ��z�0���J�%:s���d��q?�nNY��y��<�ͬ,1��O��d��nd�v޾1�"Y̅M�<7��\�+c�p	g4��c��G�#�}�4[yW�a�/��!c/*K���Y���!�U�l]��"�=�D�b����(ۮ�}�����,��Ձ����M!��W]��TԱʬl���ѫj߹�"y���l�q�ԵU�Fs����}z�7/�2s{�:�4�KJ.5�{o�h�A�*~a-)�	�nգ���VԵ}�w�ڞ�kv<op�C�6�������u�N�鶞x�+���	�Z�s-�O�ֱ3+�uZr=�?����~�^�֍�(�TB�B��\ZF�{���œ��nU��"�,)�e�r�H��˝i���~�>|����%������\��*�ݳSQ��p�󂌬�Q�lōu�fo�Ko�@Gʐ��l��3���:��=Kr��H[�֊h~��o&�0�����[�D��_���{H�!�*�c��j��w}ȴ���q�r/�`�
�T��>1o�?WB�	jYlޗ^��k7ؚvĦ��Ո���L	a��(7o�6)~��X��+E�����78�����7�8�>=�z����xu��G5��N�S�ϕǢ�t]��7o�w�F ��\zo'�^(�w׎)�_k�8�ά��X�ʱ���Y�u��f=�Iц�1t&�lI/��/��]yZ!vg�ę��|��^�Nӎ]5w��W��8�nPsŽ�֜�9t�1r
{&p1z.{���;ex��8gMWv�A��օ�
�'�W�
q�w	>�{Ԏ��_�{<�g����瓋��`��Y�r���?!��ܾ4�Py��Lќ,SГ�k3}�O)��ç�Ķ�R�p�2Y���soHT��tBu�S�T��]sF3h6	��=���#���핺�����.��4��,��6!�d+�8�v��-�:���P{�Z��to;F�p�ͼt��ro#�JH�(>�Kި�����>�4:�GjKV�s��sP+4]�|�����$����A�^���;Se�m��:�V^l���O0gI���+"d澟U�ʟ+2���	˰�7�S-�'`3��%1��+k��*�;���I�GKFVM���E�"��t[��dH��Yr��gI���Q�sU�0(��owu��D�~�;[4,�텫��=#F�^�%#{=r&���hBWM%��5^�#M�Rg�v{31O��R�ܩbgt�wT5\:�);�n�Ų���he���Ǆ�B���>�e_��^hFm�̒z�SیE:�X:�c�C:��˲�rM��'j�5���޽�[2\��׳Nz!bڹ�y�[҇4��Wو�����_��Z
.
���k�.��n_��Iq�(�����'���Km
튈ێJ���>�>� �{|���Ƕ���hW��v�ڄ�h��5�[&�-��9贌y�:��.��4q�H�f�Y�,�-��ֵ����U��*N�ֆ4����ph֑�Mc]�E�zKlz�Y�n6>��:��IM�j5��T����4z3<솖��
�)bP���;[���=�\W6/�;"��h��j��1�o��b\d��1p��4&����k��Ў��b%����U���#J�m�CdUL�8�gq�dlx��疈2�v�:w�5��9x�V��T�V@唵B(�%��Z�K�)�X�Z
h����m͐�1��dE�]a-�%�]C���з`A�S�&�
�\��o����TC�#E,J��th
iq� Vл�̋E���Iq�A�V�w	MzRWr_��r�TԲ"�pHօ�RЉh�"ZK�ﴱu�k<u����܌ɣ/�Ԗ4"�)r�m'�}� �k%���!���IkS�睥Q떐K@kT��M#��\Z-���\�.�zW��zy��F3�(��z�IG�k���]�6Z�F[V-��dE�f��`����i��O�h��TҌ Vг����Iքc�|��=�m$k��6.��Ȱ���kIKT�nи�m
����,Sʑ#��ƂZ%���ceg��5.���D��4kKAm"Z�W��~���i�+�ﻑi-`6�� �+��|����ƀ��P4��KH%��&�_�-�W��"�<�.Eָ�i.�N�g�vd��K��6�M���u-��DB
�ǃk��w�9�d8�\���>Ƨ�\���N��E�G�b=�6���a�����E�y�h�H5���`�iS�ֵ^��M}�>+J��*�-6��С�汤S4hVĺ�o�ɰF��,,Tĩ�,<�I+ܩ�Vhӹ�*�T�4Z��m"�J�
z4���}���M�ްF>g�@�ik���6��_&�W
XךR��M1KI;���}^�����ʟDq�?�/#�Lj�sUl���C��<⍮R�݇	sPciM����kn���� NUƃހ)�)��H��lA\n�_}�,A��	W`FG%k�+bFU{�`�l!K�!6kBlT��Os�ɴ���u��{7�ə�c�WKJ�0ET C8�M�{u�
Y����,����bE�^y骚US2� ��,X�^�V�+|� ����NZU��;@kUr�|��8�mZRĥ������ �����S��N_���cIìH�
�#��aa��"0GX2��/{Ǽ�ݽik�I!�Kث�q����@�S�F�X5�T�PKB֜�ޛƍk�
`����i[GvK3ܹ���B�-&eY�Ñ��N�D1/=:���㴉x��%^�h֭�m �zHb\�_���֐EBH���zҏZ^��8B�ԕP�rR�1��A-"]ގ6�k��^�R�'�����iŭ�
�`��cB��������L10W�H���e����8�5�`SCh����L�z�>���}RЌ�9�a�X���f�4h҆S����#ŧEIQT��715(k^h
`���Zg}�-�y�M6�ڦ�R[���n���s��=��K�#�
i���rlJ�Xq��[]��Ce�ϯ��6����@K�l� ���X:LL_PT���e��3IB���9\T�:��o-v�rg�l�S���9�43c���\�twK�\'U�*�3��	�`+za�R�i*e릃�v�7m�c�ܶ�t3��KT:��:X4\9���j�v]�u9m�\s�c��m�]�x�L����	����V���k۷�x6�n�o$Ӟ�˲���I�pr�A���`����Igkpea��Y�f�qu�ըnԑKΏ^�M�b���R�Җ�3�z�-��8�O�Z6mųnn��������'�ׇ+�(vl6�&����-F�ұ�4�2J4�P�&��&��I��ܛN�S���?y��LG��6�M%���/�m���m�c��`����f��iҦ6�,Gg�ٲc��9Q�s��<��%��ȋh�zIi[
������F1ҝ��h�#{ߦ�cn�Q�Բ�I7����%L�%-%u�l�,c�{s�*8��:�1���{\ش/=e0��SD>�#�Hc!�O�si1D��틴,iG�%6#j��h���d'ϐM�")�ҷ5����v_���"7ep$�ŭ�6��ҍiG���K۲*�3�6#�0�Pк�4pn�R��o�$u��r������.qGRƑuꤽO�nб��n�x��wy E��l�9)6,b�Ǝ�$Kأ�!�028T�sQ5��)�b��l�m��fg���1���{�h9��X6l�]�.�w��v���b%�k	�� {��XCJ�	KB�F��w{�Zr�l�1G�݋Qs"�)�X����\{M˨�u[&��Ì/fW�-�ZT���k����4�a��SV��
i8�$|��U�{a=�ٴ#�JZ7����96��M���m+d�)���E�~ݝ��Z�[����d��FN�$��^}������^���	wjxv� �vQ� n��b{A�M)!m�.�V�^M1���5?��Z�����EN�-,e����ĵ�C2Z֩����"�q*j���}��Xv&7v���%��T���+Ӳ��w2�l���L���/Z��߻��L�_#�}r#���)���o]�\}�o;�d{����=��5`�-B��ʶ�xu�ol�Ļm�����m,튶����	2�Z%��ĥ1�8gfn�c����a�A]���C
�\�!�k����k��d�X5[��#�-���_�-[?^���|�OL�i2�.��� �uZ�11J��C���06�i>�e�J����>E��4��[g����69!,
`�q�7�_�W�w;^T�Vz={�"y�u�*aÍ�#������E�`��M��ȓzƒ�{�@r��*zd�zK�J���d�~���pOzu���6K#�޻֮�
x¬�凫���5��)m����\���h��iK��J�Λ���# ^��##:I,i7�ҏZ�������TjI^4��N��M�)��{1�XɈ�*ې�#D�V�s�/�[��폨��ƺ���`5�P��f>X��ŎvWX�{}��i>�i�}��aq�Ɖ�JZ��R-�iz7�N:��}�~~lm�Z�C]O7\kт�jvy��z��ނ��e�v�y��b��Y�n���?1FB�鄴�;>�M����0�Aw����n�(�H-ˏ@��33��k+=��2{^Õ���KJX�����zok\4:�ۆ��@��=���2�F�l@�Q�#��#��C�\))��}�]X�F�E>{_c+W�ɸ8n7'��ʋ��R-�h���a/�۳i7��ї�?��d#��N �z�Gr^�/�J�k��9��*xí*ac���2�(K�	Km޵ǥ�z,u��Hp>k�)�nT��$V�r
؆�E�XN��Ӏ��j�C������T�u|M<�O)J���>*�jڴ��(�+���G3{+�G�Kr�8�{{2�J��Z�ӂ��(��3}���O8���Q��	�u\��EO�5���h�U@g��-#Y��D�֊b��2h�n�-�p��K1�t�iU���ߌw9�u�svo����ơ�c}r�W3,d��yp�v9%4[V�jZK�~��kZ�K�R�h�����+�d�1���ɋ/f��aY��۝��d0��Dj�ӑ�h�[3^z�Yۖ<z�X׫Փjy����-+al#���Y����,�Cd���XS+�	�{�h�2@�Am+cv��K����2_Kb@�� W���A�s9�-���4�wgתӴ�s�Y�����F.��xWt��"�s�8�μ=������N�d"�CU�{�kY�T�QWh��̿M�G�֋|i��)�#�[�޻�<�����g�3_��m��Kt���k�K1�ض�7y4ɿg�T���D�M<A�%�Ծ��ZOЙ]^t������WkR�{��{�!�)��;���>S��>1K9wt,�����ڀ�mK=���G�y�1��.my���Xw�F���! \��8���ڟ6IrCb�@՝Մ �`8`�ns|��gi[G3λ���ݸ��iZ�]U�~~�=?x�G�#��ٷ�v(�8�C=4ۿE�ȶk�+�N�Y�XKH���g�"�����ۇ�R��j��yܧ7����X7]?M調\�Xq�	i7.��-o=�,^�󶔲,��-U(D���;�8�L�R̥s���F$�u�C�'nx��>X�F�p*�M����6��$�E#kw,:�U��ݫ<㣒+&�s�G�|{I�	�'&P���pT�D,�yP���QZ�h}�[k[�/��]�J'NDjȨ����5���*J<h�!�����:�JZ>��f���԰�KD?4<ﰳZ�)u�c��~�Z�����;�2�z�
�	?r�qok7%�)���JAJ�L�j�V�<���g�/�V�3��ً�F޺nb��S�]kHiz�[ G�n|f�����7qlS��{�Y�y�K)�i� o��k�?!��l�4iQK(���o{�����ystK	�W\}+eTR���U�Ɣzm&��d�S��ůnr����V�w�t�L����Ι'�>Od�'k���Mv���P�DC�z�������V��]����l�C�Sr)<i�{�,�,��g�\(��~p�G�H��i�n��G"�s5���!�^��_:��~DL�Ow��gǂC9$K������٦QBʷx���͹ϡOz�|Α��s��$HE4СWx6��Տ��g�Q��^]ӈ����e�G(ru�<��H�ͨ�m7�ڿf\q����>� GJ�[���F&�+zahׯ4�@���Y$y4ߦ�~�f �g�cC�y����F��4X'�[������#�'�H�E�S7Z��#V����'���*��7��D��.�̗|��΁�&Jt���7^��5���{$Y�S6kJ���d��p���f,KBs�ﵷ�&<���NX5\-aF'1�]��9��n�m�,�㗷:���Z�磩���K3�N�	r���&�o\i퇞N3���c��p<.ӶQOvKuE��ى�^z�ѝ9���5W����SQ4�!��'�^'�TBTڬ�v�m��E����c��-���t�Y�k�g���ˍ��]��G�<%ڻ<�qv��N6x��O>��A�r0�3����Q�e�Ż�$�ZLY�r�㕳�ۻ=b85�؟]�-<�D�cmfR�kUI-�&��H�&���x^����^z�aq�\����a���^	<W�ή��3�֛�O�Uw�m�i���c���@r|X��[�O�r' -%$v3/u]Ԧ	�gלhn{8z|�ӽ�����E�n��Ѩ2�k�QhzUc��?Y�����!d.��{+���#�)�W�U��^\����G���́!������5�R_'lHw]7ƬZ�KnJ!�OyP���H.���6/�ת�ggh�<�Fa��{=8³w�ck��X"���ȯ`jbGYC?2g߂��I�[3]BH�p���B���γẀK,���]���@x?V��!j��w�|�}f�;j^�(׸��	�|��Ȉ��Q�y*Cfȣ����z=�e�f֋��չ�j<|H}.Fķ���7��(C�Dm����ԯ���AZDaC��Y��OE�k%�ԂBX�t$W96�˺H�Wl��mxK�,�\�ٶ�GHJ���D�)�/�)���ߚ��5�H�E��hs���񯇸k��4Uh��{�؍���5o���.�0�=��$m�����8�Ƚ��N��m�+e"r�qs����A��o�񻽷t��#��K�5"�m�n��)W��}0��%^�Zua
��p��P!�}h�W�r\�M��[��7R�;Jv����dLh8~X���k�f��,/�N�Ȱ�%�&��N��`���/QV���>h:��%��
7)�*���D�9����4'�|��h'睪�a�a�}�_�/�{�)I�Й������\���~��o#v�tz��?(m4iĚq+n���]���jK�z��ª�,��{į��{�
�У�}C��Hi�&��B��6�G�[ԯ��ͪH"�(Q�<Pp�K�����)h2+���o��J
!8�=�w��������r�m�!��-��$Q����ވ)��U�{��UM�Vｇ��ſo�>�7�ܪr��`���Uֲ�C���xx�]������i�q�ɨ�V� ��uy�@�1�]A/���8F�����^*ߴX�P-T6�j���SO���#�
+��]�K�~.'���5�)�fM���NB[N%!-���a�L֍���ؽ׶6c�[�y-������<��-����*~\@�2������UY�4�/(��{lN�k��c��D�f
��࿰���7�*��,�>��8�\��b���B�Z��E��w�QW��1<9E�죶.]?[#XR�[��	%�۽��<N�K��L�T��'ve�kn�gc��o��*����Im�E��3_Y���]]�;֖-e2����;E�b�$U^ϟnW���k˵�xm�n8Y�]��*����]�m__�{U������Ns�����;�����f���.���:�%u7-�{7�c��b �g;[�ݨ�&��w�}Y��|�v
�ZE��+f��Ï���^�{��;V鋌��\��ZO{�g0�&z8�� �]L�����7�Y�c���N�v��p�!3άq���`�?ο�����?ؾ��o��s������8_cL��?���Oz��thw�$��>�\���
��V��}3�J"�2�A���o��w����_y��B�2���N�mg?�����^�2OS'����8oM�w��c�y<��i���_!����P�H��;���č�z�*�G������0Z��g-�������=�R�b�Rn�E5D�ew�P�%Kۡr�[����FrB܎ѻܢ�ԏP(�}���IVd��wW�{�u�*����?I�te���%�xU�eq�i��vp���nu/�������=]s������
7��fC�
$EO]М���Σg)�����>�!�+�G��{��-f/S/e:�����p�.�m�K�w��)#k���,���-��%s��M*�M1�׃rK5��0��מL���E���<{2ͺ�[�Xi1���8<j8��w3�g���:;����)YW
����dd�B�NC�m����^�T��c�8Vn��	�&�پ߸��o��v\>S|{���z��P�@Ѭ��a��X6!1��mU}�����i�;py]_�e-��K��׎�l�廾9��G��!zj�Z�^�ߺ3Cw���g�zZA����m�Y��Mr���^qn�EU;���Bv���@d��\$q[V�^m,�u��f��r��)�<�y�QJ� �t�3����I�>�z�:�t�֗�7�vo�̑�^MM���W�X�)��®�'����MAr�p����s��	sm�yc�p�w=8�Z���5՘M�����S(YM���I	/�@	$$�� HI~�$���($��� $���$���@	$$��$����	$$�� I!%� �_� $��� I!%$�� I	/� $���I	/� $���$����HI~��Z $���&(+$�k<�2���0
 ��d��G�|}�Uk^�%TEU+m*�!
lu�"�(U!Qml�
�U�P*֪*�!t2� ���R(�XA()*���"�RUQ�           �    �            
     ��     @��c��ݾ�_>h���:�zkl�,�n������m�� ��w�]ռ�x��K���
��zysU����;��{��� ��of���YK8���*�RT�Wf�{˽������v^gU٢�]� xz򧻷����Z�q���[E{�:;ή��ݶ��ӭ�� =ו�8��^K{�y���4�=�ʷ����{<�:ua4i���      �  {��Ǜv��ty�e�l���}�����^nK�����( ���&u��֫�N=�.���f�/v�(��^w{�Z�Sk� {Ƕ��M�sڞ7]��{��KMD��IT�wl�=� �7����g���l��| }��c�����}���wwsm|{=��I�N���َ����خ��6W�E�l���mf���_o/v�续��kto,��ƻ�����u�5aG֓���x@     P ����m�����v���w`o-�L�;�n�{w�K��l��ҝ��� ����gϹO���wsyνoN[u���k��y[�n��wp�� ��ͷ����xn�m���{*��)R#U;�n�iV����+�;�� g�Y���y��ٵ������nAm������;7�N��ݵ� �:ކ�<����]-۞w�-g���=�S{�:^{v�{t�v���j��m<       ��m�ݶ�����=���ݭ��v��=ݽ��9nu�{�ٻ��� ����mq�_6�Y���=z��t��{v�Ir�^{v���3�� ��������zݗyâ@��l�U^�<G�{m��ʕ���Sx ����m�{W��c��Y��n�r�YGU��������ڼ �Զ�;��n�G����Z��������n�i�����l4�   �     ���_ |Mz�}p:��0����${�p�AN��z�������w}� ��� s���

��}g!�>�>��
D�� =�@
 Yo��@GK�� ��%EJ����W=�����h����|�� �P^�� N��:�>��_,)������B���4x���>��އ�wQN��س�_ ���� v��nzv
;����݅� 8�B�z� �~�R� 0�2dJT� ��"���IU@�@ ?L�T�   j��H� 4 4�i5J�����e���������xn��s���)�F��r���y�%GU��W�
Q�"Rg�	(�Q1	B��!�(IDB���$�!DG�$�!DA
Q� (IDB���������i�kF�_�1[�rVh\2������VX�"�@ɹ���\yi��)������&�w�����Y"Ƞ�'��ԣ��!�1��c]Ǉ0\هB�p-lL�Uޛ�� �L�T7��q,��XD�)�i�Y�_�NH�e�5����m��=ܴ��n�im$�*�2�[4��i	t����o!�d�B�n� �J�:���5�>�{�l�]�ϖI�]c�rSy��R�N�<���j��Φ���02��²ًw-Nf<�MC�	u�2����j���6�85n㡳m^2�ۀ�4�E���kh��|�G�����u�Ȫ�@�if��+Tu�`&�t�\XwsQM=n�Z�[5�`AY��Iw��o�;��5N�C�Ir·Y���\.��͠}I�b��Y�f?d2�����
�z�7�hK��h�����E�F�VCx�2X`�*;ֵ;�6VH�ݵH��f��Q��[��4���a�ҁ��n�`Yg(��0�Y����n�ͬirk4D��yKe�h����n���u+if`��q7�4?��N�hث�����2�V�L�L�кyNP�����}��+^�l���0�#���(��Y��:K��< gq���˶UdXQ��KU�Q7����ѽ��ax�7"���<Q�D]\YcFSp��R�◧�+�qD�=�K9[!;$ ������w���i���X��&�����F���^�$s����x�U������Y�T��ǉ�c�E�M�O#�`U�r+͡��<I\�wˍ��X�e�75��2�j8�fa���S47�~D�ڿ�ʳjHj��-�v�7x#2U.dsEBr�m�Wy�^�Cq:�P��ʌQa�o�f+S^��YM78�j�mb{	8M��*�c)��
A޽i��P�W�>����66�VD���GЪJ��lt�u�S�ڋ�����Y�&]; ǝy�v�,�X-]Sq�{K\%��L!i�B�[�9���f�?e�%z�RQ��l,�2u�̨QY�c��I���KT[���k�N^e�51�1���]�t���PDP֦���Ɔ�Q�؆[{S+lf��;"�H�ݼ�{�/�ѻ�`6�e�Mm$ٶ5lb]��
%�KE�*��6��hV��B�q=L齊�#�Lk�^y�z�2/2�*KF=�qSR����l�㽻:v v8�֍@m�u�6���DǩاI��t����.]��<gxV垠��R��Zc�Y��ޗ�5�q,�ZW����,#m�ǣNn�62�`��Ʃ"[�%0���T�����B"��3q�p�;�r�;y�i�Z&�i�}���Z�*�m�X��.��Ȇĩ��f�%۱
U���9r,�z�t�;�d�V�3cjS�^Ԙ�҉"���5U�zQ�jn�X��zX�Y�s9�?����i�0i4�f`t�e��K��t
��ƈ#�cƲ��<Ҏ!�J�X�q�J�F)��ח,�ڰ�c+6]��f���-�����S[8�dsMѫ�� �@3SE;/ �Pk���� ,-ɂ�L���J]ay��\:U]H	�H��`�H�PLq:9XG�3<&�k,�o9�U3>r�5��"(�+�Lb�����q�z�nL�26�Ð�����F�����^�]l)�<���%�l��=m�ws��əW��s^�/T5pZ��j��ܦ�6�ٴ�nŶ�-����҅
 �Zݳ2����:s Gt'�2�i�� �E����%<G"��%�,#��7qXGu��I�Լ���:�����\��ʓ`�EZ��9{Fe=FV�[�Kl��!������(VN�(.�֖CQ�o��7ap*pHU�X��K�ޖj�5����j9cT��e�NLU&�	+ke%(����e<�̴ ��lhd���1�*Td�G�@E�R��O�HD�rᫀ�x=0V�r�ZD�w.�l%��e�#;2����+el�tU��e^����qAw0
+%����r|o��e��[0�=�R��c7�[����ц6�U�5�N��m#�S��w�/S�P�W�Ȣ����Y���bn���t[Em�8n���/)�ѻ8�n�rY<�/S�h�ڗSu�7J���])5ee�TvM�Tsh@�*  wkdg
4M�S9�n�2��j��z�A��V�������!j'��df�e�9�e*c&���u����.9q^��c�҃NK���-��Y�U�(�:�ʛ���ҩ/2S�&���J�Q@��Tb
�6@1����1yj�^�I��QaQ�n
)lM�ŢL�pDn�a�k4�sD7��	y,��X�`���L[�یճ�c蘷X�o]`[��
�9NV�0���sU�x5�^�&V��&�è3MD�l�b�s�����V���Is�r��q�F��x��+V�&��܅��T��;Zx�����b
n�����ecӆbw�z�8�ɲ܂��(�a%��]�ux�	؋8��۷��y�� +o>1�&n:u��&n�XS2Q���Ć�.��2J�ū*V�P��ęm]��4��8�l�n���\+ͻ�W�A�g<�0VV\06�B�IK+`�kv��0�Gp1l�T�z����yK��`c�,�[�k([Nd��8iQB�@�S)�j�ksoЭ�)ٷW[�<�{e'�v*t%d�C&D�@�#�h��H�A���܈�#@7�C�0�1O�v�6��u`�\�Z��rVѭC#x˭�v]����2J����N��"�W�����6���V@����y������� cx4cܬJ�(G�r7V�0�ɦ�8�$�{bV�fR�B	&V��i�,���2��Lի��҈K �Z��/�i�j�j4v3J�$��"a"L��mj�	�l��i"q[��L#Ͱ��nM+4���e�0�U��R�����Zj4��a�Y6X���z����Ou)���9F�����%�J:����J����(��u�������.�=V�X,��$�bGL�zC0�tfL�(F�f��rm�Z@�Z�
lv�ͅR�L��V|kN
P�s�cJZ9-]���tPI�fpT�Ջ�=wq��^fZe�)@��EՍp;���k"r�^���7���m�4�5�L`ҎlF�k���LF@j+˷Y�qS�O6��.�rR�ؤ�P]ی�/>�����#"E{s��v�[�UrP34ж���tD4�ӛ/�jH���UC�U�2����ˣ���{+ p^[nTݬ�]=onb"�ڷx�٧+�K�{��ӯ"���Q"�)	�>�����fGX�U����l��E�S[�i6ۣ5�&Ĳ�j�v^�h'�mac�a�Jf/R�wn�nCq0�_5�&��u�#�0��$!�ʽ�����稖�(yz7A!��ʉؼ�!n�L�O%k�â�� vs5����
��iD[E�5��N��h6�\�Iʚ���,뎥�z�J]:Z��g�[�J�WS��7"Ò�гA�S-�^�$׻R��l�~�EY4�`�#�潢^���ӱv�O�U ��G,�f��G��II
��V���XO Ƕ�m�����VHƣ��\tb8��D� ���v(	zv�?���K&�x����H�c�B�k-�c,�q :nl#O��64Jh
yB���c�j��wA8iA5+4*�%���SwY)̙�i02��!KF&�Xi	e����&���Y�(ܐ؉=Nȫژ��9x0��v�(�C`�xl�wcu)5�Ȩ]fD��!l�ؒ2��]�S�Y�3lcR:&]�̖��50ʠ�f����/nݷ��ֵ��@Ҕ�OY�Nָ&m,��F�H�*���&�^��{v6�3�H����L:ja�2 ��u�ثʆ��b����5�]kXr�\�c�ʌ>#0��D�^yC~�$JNK�	�Y�	&�1��^U�{PSJj,�lt^֛�-L҆R��Mj��)��ED��� �N�f�%xчC��:X�x�c�\s��S�̛��ˊ�Z�b[O,�EGf�srd?o@p�v�ˬ�#vS>�mSJ���#�CATҭ��uy�vCF��Q�5����$�#JZd
�ƕ�A`�!b�Ŷ$ܕb*�2PQ7鵬/�A[b��=x.Y�&���A��Q��V�,�m�r:s(��3j����Iނ���4�GvSԝ�n�앻�jbe�B�t�����Y�6�$D�)n�A��[P�8cֺ±9h�1���H��A��\��V2R�;X�]�m;�AǷX+]3�r��f�ӗ�� ���k�ō/r�r^�,�Q��p`��G÷�)Mm����5��ٍĜ�JT,��s�xw�S&� 6mn�sIu4͟l���o(:Kzh�M�e�h��t⡋^�YC	�]&�f�B��Z�d���T�G0M�ҙ��d�kRW6���ۘud\�^��q�8�h���'f^͉j
0Q;�T�e�n��J�
���ډm�3�n�"§�=�&���4�mc�^ۤ��F�!#�YjemY4��U��M8�[-�R�V���X��R���p�@�u(;�]��]���1���n���t�׿^$�p�{n�[t,	wz�B�+^��n�U����jܛte��j�IF�=����L�6���W�EB����SǧE�Ѵu��x�@�Wp�{g~h��c3 M6�j�(0��6K�u��ˈc�-�Z"�;�ڽ 0����̰Mf�$�Gٌ��k��RQLN��l}��'%��M2X۴Q��2��#;3vl�lkDi�f|Z����aƾ���#"oN��V���aV�r��hw*�����,
�!M��] ���0��Ιz��j�>"�~��;��f Y�@�X�fQ�^��R6�	݀%f�`�l��-�?&�V��e���Q:m�X���^��1[��d��blR���&7�pY��]���h'�J��ZoPm^�:hl��BW��Y����j���*^��h�X��m��xUM�/^i���At��h��O����w,�**�J�d�ŷZ�೘���qXD�>��5�o*T:��nQ�Uw�Y{�s�+""���*l���ZvE�@����.�ʹWc��Σ�3`�	��鉻��EV.�`#ieB��W�.�Y�\���5u�!t�H6��u��-72���!f�浟(�sq;��کOF��2�sd�[YY����+�RV�Ssj��v�ꎛ�:��FH��(n�jZ��j�M���m=�x��wB<`��Zt�z7Bg1��$���
i�ٻN��cqYn��T��b�H&�p�X�.�S1,���6�]�X�,S�8�!U���T��/7�I��~(�����m�B�	�.��8s��5��e6�b��5� p忷�oe�"�L��䧱I�g�Q�eS��Fa4�G��Uѓv��!�T/j�)��13��c�ȯ(6�C��)x3�Vj��Φ����ds�'+1�EѠ`�I�+v�]�Z]��2�Z�̎4�+��vr���L%K�݀&��h	��tk,�2�;I�XN�-��D����l��<�p����z�?��'����5r��&��ń��ǳpѦ���M��ۣLnS���&�J�K�V��ÖZ�(���ˎ�m�ti��hJ�*7��&iCf�[V�ʹzƠ�k QJ������ʓr�˭^^�)J�`��&��HE;"��ց�e7�d0�f�Uۓ�@朻:��VԬ��"K�S�am�KF����k��d�2D]l�2�ܛ���f��j��K@P�z��be�R7�X���Ot����ٕ�\s�{x����!4E� 0CR�l՛�S:w�Sr�+g]�ge�u��%�K�0���ZF���(C�I��AZ`T���	E�V��,.�Xdj�dnW7����x���{[rd(���sj�K�S]jU�7$��!��,��8�X�c�\YM :��l��#�r��v�Fv�5�L�6�p`���`��� ��&�.U*}6��$�8���հ�Rj1o%b���9���kj|�Un��VcT���Iz��r�D�T�ƛ�P92���jT�fE�5�N����5���h���h�4s4圫�٠-�𚚯q��1̡#%P֊�c��#1���S \�Y�F�h��HLܧl��ES�MGn�/��u��wL��2I��������iel�cW�.����"��FC�54������	]��2�DY���i,l�:���2���W	��0���U�A�dزż$��\;"�Ƚ4�dG7(e.Tw!_�&�L
�M�Zܱ��Ѐ,͢/�IP�oL�V�l�b�D����T�w/l�2�w&V&\vf5rjiٵ[o_ʋQ}Z��%�Ybe�Up�W2���C�s�0sZz��M�Cv��.��p�l��'/&��F�#f������;X-3�fU�X��SrB���G��FDr�d)��hi�w(�̣�� ���YGc�n��`�Q���[v��KE���G����5�����c�4;�B�H��+�IN�M)���j
:���kV�c���N杛� ��ʓ&����BH��!Q�il�
ƣ�8���xoT�A��ed��]e�k����ah�zsVk.9��2�x��6�Ľm�e� l��Gs	Y��#��5�rV�����x@�.-�4Zȱ3���7X�f+��wm%�sY90oGnə�p��tP�!"�j�
�qe�̹���Ňn��@����������A�@���:/n��,���|�
��D��%ؗ qV^2�9Y�Zj�:N�Ӧ��r��{2P�>�-`���ëm�m�����Z����;x9q�jrΞ�9��t��:d�/;��ڍ[n���hQ	Ӹn���*�m����u���hnf�l75v7\l���;���;�ݞ�<qչ^�y�3vX�?׵�	>����e
��ܚ�Og�K����k�l��1��n�q��nCzm��8�=r�����lx�n���v䤹5�z�t݀7\�v.��v��q�s��n|��;+�w7��(�p�����1����Mֶ&��8ż��&{9��[���ux�D��8d'u=�����^��N��-6�:��Z�G�-;�:k^�Y��jݨ������|[eG��v�컮�#q�lR�����wM��Gs�D7W*�K���8�!��<<�]�^�e��t��×�m��cl��T�4�����Iӻl�v�ғ۷ak�K���6��Vܞ3�y7^]խ���h�٭����g�����;w���}pd��k���ݞ׊p�۷۫����;�kicO4�XD��v[>�v�b{*��3s��.B��m�N��0�wZ-N8��@��vL�vh�e�r�Jv\�
vχ\q�~��mrE��w?d(����9ܱ�L8ؗ�����ύ�gr�#���O[��nT�]�v�!�<
c�g�uڛ���o+i��N��eɧQ[ʚu�4FM�m�x�+Wc����Ks�����bq�9�$�ٷ��p��̓����n��۞!�����`��܃�]^uԽ;�G�W��r
)c��Vm��k� �/M���u�=ۍ����E�|&��L\p�����^�j��&ݵ���qX�8�]��K&���s=��t��%���є�o;pҦvNITpQ�cnkv���l�q�^�<v4Fr�H筓��:��p��������q�]���1O ��Kv׳��`�{YǢ��ΞW�u=��㋜ik�>�۾�����Y5���NS���.r�,������N�{^7%��d��偈筻	d��7'c=r+�fn<�^��w��J6� �d�*{0�9Y�u��q�nW�LT�pf6z7���p����u���ކ�횻 ��c�\��h�<��tj^�R�8�N ���]�=�x���k������`Ӈ��M������t۝�L����ۜ��G�����`N��v/r���ô�糎#��F湎{���v�ݬ�7-�l������0b{L�c�^�'Ʉ��e���v�������6�pq�;t��ûq�|�mpmbp��6/	���X���ݠ^�pn@�Ɯ�.pl�d;z�'M�*���ٍ+�����fu�69�N�u�Hn�\�YRvta���om۳�b��n��<x���^5�#!� n3��k�QW���:�X�w����x}��۴��Oi����=e�q��c+�[��6q�O;r	֍�撚��vŝ�!�`�n��Qmlsc�Fw�tg���m���^��=n��l�������G(f6xʗ!��	�Ȝ��#;���u)��T��л"�e�]��ݻn#����i���w��v���ű��uq��;�W���^�w��ѵ��;i��3O;��$df0� ۃ8�/jƷ1��ѝ��[�=�����j*���z��x�)��/=n��6-=��.���wn1|��vJ`��]�?p��Q�;wdXA�;�ےݎ���s��Zw�\W�v;r�xu�s���:�ܘ�Oq��J)R����Oek���ۖv;rf�hh�m���u���ڽ�,���;�k�pD��B-�.�v����ψ��s.�M;���z�^U��n-��sx��l�m�è��]�p�,��]����$����uy�n���Iڝ�X��1&a��=�<k��t���M��*���B�ⲙ�L�8ݩ4��^�]��9x�x�tظ�l�۵���7�CJZ����'c4�n�Ӭ�v��fn�N1�lv��ˣv��s�6�1[v�:p����^.3�n�0H%<p�!�6F�J�d�9���,{]v�R�^8��nqcb˛�a��ɭgv����n��,&y��A� ��l��Y}D8�Y���=��֦�m��s��j��u�j��f�]�C����Y�`�۶�z���n۱��kny�u��N��wO9��1u�m�����Fp�:n�'c��ұ��`�wj��4=���s�F���Y�^��e�t�̋��Y��a�����i6��s�c]��m[�����y�tj����6�tU`�æR�p`p��7Ms�+�^�6�t�pn���ϱ��-5�\ط��5�p��������%��TԬ������[�sɈ��Cf{���v�����G;G��;k���պ�r&81��y��}7����<m��i��1���v�kf�A$�t^9�Gm:��[>��^ݳ6s�k<y�j�����"�}�+����u��ɽ����N���%<M�o����Ƭ/B�-�KWHp\gWm�/.�T:�}s�=a�d{��Ik��f�!��n8��+�m�=��ӎ�ۣV��c>5f9���up�(�s�h�si�us<�9-m��S��g�т�[u����+���y6��vxzM��ڽ�7cs`s^2u�825���lq�m��[��A��r<lu����Y�۷k�����b� yvv{B�1oov�n���7V����;]<�:���ˍǇ<gV��!�;�X�(���I�]��cnkn�{k�����z�nGY��:����A�Lp!����r!�9���v��eQ��뮇8C�G�'[���6��ni��0j-N{V6��Z�5�98�#8�A����	�E��<E`��]��m�y�6��.l�H9NlI+���r��͎��؎���va[�oB޻��9i�r^z໅�����q��3�;c��1��÷.}3)a�q%���a5o	�O�����!�V8�[d�m;<>ˁ�i}�'8���=0�f��PP]�Ru����s����]���.q���'7�J��.����!�8;d�VQG�!\�ku�x�=����z0nmc�̙���r�p% X�s���5N��ݮtX޷m���ۍFf����w��1�o	e��e�n���%A��N}{*��C����=��g����X��v|<u���''m\cd4�6��L��B�p�hΉۋm�����|�&����w=r�J�2h�n.M�u�z�C�Ȼ�E��]tA�;
t�P���ļ�����T����cZx'���N�g���]�꛶����� ��:��[N��ޮ��8����8&u�7e�fb�p5��pA���8�u��]��:%��q�ӵ�n ݇z�p���ܹ�K�O�٥�u6��	^�%�L\�N�	Z�����7'�9���	�:5v�x��YSR���|��.<����O+Y2��=v;k��:h�<mnƧ��A���a��k^QՉd+u�;���uۜ�I�aC q�㗱.�pn&���0en��É��!�\`�9�뗝rv�=q;m�H� ���**}P�1\M��H�H�O�&������������;��1�Q�9��;��-F�m�E����vU�0c��&s���u3�qѽ��v�n�&ѣpvwj�Żu�]��ue�66��m�������j]83kv�ٞ�kk#+2W	��`w7mv��E������)ێ�6��vK
cnw$�\��e.��9�n�ڞ�Ӟ��Ɉۉɉ4�N�s�ɶ�k1�;ҥ��d�;�sŷ[���3u���ڥ�u��^�9n���mƧ��xsll���M��s��
99ڞ�)��
8���n��@�U(т��w6"毲�n{��z�h�X]L���R�ɱF|�`�+�g<s����Յ�!t�[��.�����@�E��=��u�- -M��2\�5��=A�=�uV���s֎ҽ�`�9���nz�)ۡ�����.۰`�4���k���p�
tr[�-Ճ����l�aN�KO�#K�,����y1˸�� ���ݷ-�Yĵ�ՠ�Ż��ְUmo��y��a��n�3m-6��Z�1�v�v����9�����f",r���s�� x��a����O\����c[��m�;���W��M�Ogf��t�:va7��;h��.q��m�v�bwS�BeXFD�EP��T!E�E���N�LW[��Ѯ�;D��t����ur[�D��\���цK����v|�-���kg�c��Z�6$ѝb�1��#�T��[��4����ŎC�bSܛ��u�˙�,�`�*p���[����Ǯ!^�J�h��@'�;ms�l���.�O6�ÂK[vbw��<��8����;\q�t��N���b�c�n��í=�= X�m�=m�soo8�$^:��k���1��q�x=gv@�\vl�(rg��f��^gâ���:e���t�W>M���nW5vڗwf�'+��1�c���.�YQ���ۅyS�{'�(
�2��ݻR��|k�q�r�ܗ�۹�3�g+ Nݹ9���qښ���:�ȡ��1۝�8yϋ$v�����\7���b��$�h��]���U�Ҹ鲜Ƕݵ��=�v��[ �)�^���۶��fsh7n�M8�U�9�Y��/��.��=��Z���۱nt���|Z=)�;�ŷv��M�{;c��'JX��<�{����_����7"gÌ�g�0vQ5:^��}��m.�������5o=f����1�b�g�gpm��y�6�\�uΆq�#��/<����#<6����t��]�e��mt��w��ew"�n��[l8ܦ��89U��;j��럣�������-�7>:�Z���e׶���d�#��n�֦}�̧�vQ�p ��v�񧲢r�'Z���;z��v�z��ŵ;8z��,u���˸��N�Gm�v9�GnH���&qݦ��m��c�7�TU8�;!�5sa�x.�����+^�C�y$q�;�T#۷1sSxٞv�a�-�y�����X��S�nJٗ�tU�n��c��q�XGqۢ�ay��r�:懇��>���(J"�J�I(��
Q� ��~���!�����qrΩ8K����/��˽��jq�V[]d�ڜq�;�g�F�c��m��۰�'/[]�]9wn��u���ɺ8��v�m�Ο8����(�Nқ8�;�w]/�d{i綣�3��knxK����9��׌�v�W^�wX����"�8蠪eQ[N�N"�:�;��K��$��۳�vr �r���xַ]�I�vwX�\Y :\�q�=\#[��Nv�������<Cy��ݻ9�;���kvK��;�į;�M����{a(��y�v�l���v�ڦ4�Wh嫓1�.�zƬ�ZQu�W��8�"#�od�C͸s��F�5�n^.�����z7�]�x�v;=YѨ���sƧl��/h�R �;m��f.��6���:�Z�Hm��>ڻ7<�X^9�v-���]�B�zp@�6툵j^Ҳ����YUL��z�q�WTô�Z���e|t���[�K��^���-�ŹSn]'�^1�;n��;v{p��k�|�z�۞�o^:���x6�q��������nq�����˺-�����t�Ցo=�d���&�ѱ������ќ�y����nv^�r����$ѣrg��{n��0��G[M�ywe��玹Ƹ���n��������m�v�ƪ�6���v"y�W�<ڮ�ؓ]ێ��k�a�1����m\.덟Jpk�Z��wp��Ź9��� ^��qK�1=<jݝ����g�\y�h�FY�G ��A��Cl� l��3s7dt�c�'f7���Ҵs�2Q�p��s�]��k��ꍰsI��w=KsKOD]Y�����&oh9��/cr򕀏1�)̧��m�R�c�\�A��R�X*t�3���m����Z���Î��u�m)�����9�>�=��6c��9f�q�t&.׫E��8�f=��7,K��v욻kU]\���:0�-����8*��� �'6�M��n�:w]�����ʓ�;c���)V�(�Q�BJD$�B�P	DB�
!D(���P
"@%� "!(���Q
� �I%p�R+�O��	ݞ�b�w<�6;qy���s�@�vY�c���x�鉭�x��p�N��n�;<>��q��k�:�kpZ욹���n6��[��8�oNB㧋����ӎo=��"3�n�^������S�����n=r�^m�0p�k �Ŏ�rr1�G���@�k�=&�vzU���v�wbgzܶ�6{g	<���NA�s��p�:���wYҼ��78y�ۅ6˓���{(�0�Og��!I�M� ��j8D��������#�`���n5�fOP�0U.�œͫ�,�I�ڹ�*4u��v��洬I��	�嬮�� ��)>N�@�F˿�|��D�g��i��''w��H�~O|9��TE���)�nͿk�?-?\5.��&�����M�)0K���p�Ϫ����m��8R4��>&�'�9O�֬�HS;��'uc��'����ڿ�8��XIBו����
����C�{T��0_o�_|�B�nl�sj��i�#�K��\>���b��%Z�N�UN�&^��TB�>���c���S�;��/������է�&�ȷ)f�;�G/3k�sĶ\ s�e���FG
!P�G����g&��
HRH��sKH�0���P+�BsA%�^cB��8��MXC�y�y��	g������[s�p� ��-�b�0�(d)0\	io�lLLQ��CI��?R��;:���ֹ�>\���,j��O���K��{*ic�>Li:��&��SǮ�+W�(nң#k-�M8��1�D[r[(G[�Nݹ�OJ��G"W=��}]O�GH��M�w=��"Ram���ǃT��5��ΞTȵ�,wظ��V��j+�Ug���k@�qM�}�ڰ�'S-�����Bnrt�� �c�c:��J�3��:a3x��������tW�K��[Ɍ�י�"��^Q��0���m\�,��8e���A��������u���Ҹ�nv�
T;{cdoJ�W_m;�2�)/��mUHunX���\��D�m�[�^>Uo��h�1�q��e�WV;�I��s���M��ާ�S�ضp8��niI�t��m��#�v�l�#:k8X5�tv�u��H.����@��w(d�}rT�Fgfe���d�B�Uڴ���7wҢ����;��rV�1���k^�Q�W	;R[b�u6���Z�N�f�hV+_)3��z5�AU�H*��5�ݮɷH3�Xݗ��C��=���0�xz�{c<�b��]���69�/Kw��3�Z����1�`��ޔ��(C��'�ަ�w�*`�@^px+2�.�/⨚��5%O��*{��ײf�Z�AY]�h߻C��x���S7�g��Ճ�}(���U�̂��L��UY������ �U���twl�
|�G��0*y�:��ə�T�w��5�-,��E����^�]��2��$�v�x���.ɷ��y��$o�����#�8ֈc
v5�X����l�eFaa�WiP7�r���沊�zЎ��]�E"�-�)��ŷ&���	���=I�E�eN���Z���[Y*��Tm�YGmn�P'�����0k���<��|<7�V���m"�lK,(�/*t(�%\^��9ҝ���ʈ^,��t�S��9�W��7��kzt��9w���q��J���;2�ݳ�d�#e�wB[���ϔln����qZ��K[�:��Ky���;�q[Q\��`�*��E���-p�0��ຽ��m�J�;�
߷��%!�5��k���I�_�u��x5-��^��l�`��)��=ANr��u�߳�;�iiR:�)�,��9V�9�Z{]��w�r*�j��A�ޛ>�������A[�o���2�u��o)L�S�2��ۼ�=��W̡]�\�$�]$�H;��]���7���egq�[�B�#����N�yDR)yo"��e�A7�̨�t��S���C�I�Z�;G#����t��YJ�;;\�3M+��k��u�m��v5��X��T�澘h�k��k�N60��8ݵ�f�U5��{w����ϧ�}��eR�2���pb�{]8pbc�7K]�4�"�n7�SQ���R��Lx�����V�G���՛�K"���ep���Ӎ�@������]�����%���r�/n��nR�=뙂R�/s>t��&�\3X^\\�f�aF�c�hl����g32:�<�� ��]7��Q,��l���6�s���J�*�h3m��=tN�F�o,u�.)�L�
%[f��%
� ��8�&��	�%LU�;sn�����ٯ۾�!8%�|Gy�1%�'+� �e�o=ޡZ���+��*���ǈ����[�^{��|�Vۓ�ʴC�o�Q�!��-�Z��/��ND��ͫ�r Ƒ�uڞ]g�|���ah"S���8y(��2ص�%�A^;X,�Mo�{���;��t����N��j����]�TM�w�YH+<~�̺���.54!YB��a�U�E��)����C��PoR�0�n��oj�i��'wZ���;>-����%�����,S5�jإ䳹�v�g���c�������)ڣ=\s��NH�XԹ�9筅�ollTnۭή�Ōc�%A���tt��Cv�[���]��igkj���N�oc:�lvwn�I�& �NyZ1�y���
zb9�	wGH����m��Sv�uĝ7��M���`�&�$ݝ���۳A����7�l�ۡ�L��ۣ�k]=]�ϴ����5��!括�l�,V$ґD� �5k�'��#<)��قv��\���ӏ:�]�걘�\���.���5ii��o�� GF��5���&��x�����7�d!Y\��8����>�~i��~>w��W+<vxI�����!���m�8�)R����c@��f�x�o5�@�w[�4m�: Y�m���y�ξ��6�P�i��C�3�<����*/r��i�a�*����ᵪP1�N���ŋY���4��Cj��D
*�KQ�so(�zkt_t�͐�W=ݪ�M�[��9$z����e|�N�����9�=�fӥ՚0�XJ��6PJ�r^��oB�Bߤ��z��=���7.�Yź=f��k][H�@�]֠wY�
������$P���ܜ�h�%@�H5tQ�=�|�G�q�,�S��;7�T/cu�X��Yݧ���Fe���Tv��4�C����k)��D�z�eyL������K4�ŽVw�B��`�f�ޔ�43�����6�`�LX��r��vQW���1iM�hbC��[���,G�}+O�������^��"�Njޮ�	d���H�g+�#�F�Gu|%�0���w&��d-傴U�ș´��}��W����ӹ <'o�1�y��j�T��4�-��$k�9�uǱݞ�˳R����&�M8�L؅���Wk�g��<}&xK��<��h���o)����PH����J�7K�����y똦�YIߎ�M���f�)V�m.IJ��S;�CHե*�S����\���|�I�_9���"�l���Z氎k7��w��m����~�{|�f�d3]��Njb��I��e���l�5�)e։;�yO����/2[���%WWH*4�۷WfJ�m�<vGt&ݻ�/��n޻��;g�z�0�T*��~��%Y�.�Ӿ��涝խs�H���	�fI4OC�Ol�Ҷ�[X�K��{Zݬ�ݧ�@Q
)
5e*�%�����d���g�/W
m��Oۚ\�؇�d�vT�Y��)�D�4���ٕ��5�>��m�@���)��AMV`��K���f��3n�f�U!0�ft�=ȩe��OL�ٸHj�S!�;���O�i4A�w�O�l�޴v���ؕ�L��[��ڊwE���Q�d.*���R�-���9 ص�WLgQ	N�++T���R�窀J*E�%�aL�Z
�('���1�����kv�u�o��xPG�|��o�i�/��{��|��M�VZ�pÁ7��|qG�§J�-���I%�&�r�ہ����`ɛ�쫉�mx���W	��I������Nw�^R�Vf7�K"Ú���8��4�aUr�A+���8�L���aB��������4찑���#�X"���%OU��/�j��s�JI����,�<̔��Ш���iT��o��C��ަ���7�V'�4�k�J�Ao٧�U�1{�nS�.D\��Y�:/c�l��V^/��%5ˠjkv�eIow07�Ϛ�k��۽xp�6���U��6UY)ӧ]��e_j��!��\���}Wme��ʌ䠏<��9��|��mn�z� �K�O���a�5\�ٖ���z��5D�!$�kZշǦ��A�ww��A�gi��7w:�
Uۈ���C(�
{��e)�m	�Ee��k()՘χ'���z�9����k4�g<��ev�������[Q���.���lj9�Em�L�o�v����F�vOlᦴ�����Q2E/�����K@P��K���Y��4:#���B��\��"b��\�v]�t�^��xlk�;]zM��~�>?D��n6ׇ�n8������I��@�<q۴;�r�m]����I�T�**&:�$�]ޥv�Q����Q6�s59}
���6�!��Q)�w�;�����XƢF���aӣh"
H�6IQ����4+���t��zV�P:7�s�A��fR���{�S{w��2��+��ӽ'Vɖ��=�yz,�K�M�UM�]5u�>Mz6�H#E����&|͋C��v�cmG�$5�ŵe�ue��;�v�H�M"H���Ly����ǚ�u��&%pv]L\�M�զ����"�[Xr_vס�]��N{mN;�^?�`��D�k������\�S��K�������M̷���_q���N���R���u͡�ٿc0 �=���M��Ju��O�:?e���R�^L�-LXj$�����o<Nǵ%�t�\t@G(��n��wx����i�7NM)��Ͱ�Az>T���1�OV��q�9*����9j�'`cXO;�7p�m�kl�rm�4�Bs\ul����S�y�;�`{m`�'6ⵧ�\)��m��� crȼa��o\moi�/]�n�YLܛ+u�vs]�ѳ��ܽ�mz��W]��t��2b�ՙ<�'��H���*�Ɋ��7��k���ݺ����A��$0�#��l-&鐛�S��&�N2kʹ^�8��;n��O8����wO�4s��.6�:T�[m�6��<�I�A�F��eI� ��k�o�r�l����$0=�D�Ʀ],V��cЫo�[h��xss4?�K�+�}!)L���=:��i0�
�ɐ��1�_������Z�Z�6'sN��$���~��֬.OWk̚��aF Z��d2�[aV-ҙ����ѣ������[s<+�7��ЫU����Ӵ1-\XTț�#ۜ��U�I<�+�a$(�X��=��Y��ryf�)�����P%|�{ٝ��-]4m�t�������ϱJ�^�N�E� Y���KaC����yK�+,�彡ސ7�W0E�lcg�Yg<[w�o��w1i��d�Zh$u
S�`N/D���gi9�@��]l�;V�noYνrk���� 6�|�N�(�9�Q�uָ9ښM^f:�%����;��F�:�Ig\��u�t*CA]���V�F�J���(�UZ��w���[*W���+#�1Q5̭����]� �mfN���u�����no{u��rS5��٥����h�·��@� �K��'?lS�}�Ix�{���vEq��ΰ��Ⱥ>/$�R�"� �H�J��9&;��^�\,c��p�e	O֡�oQ�,���ܼ.�f ����h�2�Uf�C)��8�@��&����+V�%�|e)��I�E�8&�K��f�9y��p=
2�L���EX�Vh*i:��U�F��gNh���{*�-��AU�T�]�A�lu�~�zN�2��[w�L��Q8Q�>n��^�z{g�ߟ�	�uA�q���� �k��DK�^�R73d�&�p]���5��R��#j�o�^�/�H�'��"�4���S��~j��[�u�m�^t��x�����ݴ�8-��h� �_2Ua�j?yS�NS[�����2���,
�<�	\6a{����{�1`6������I�ݎ��v�nj��ҏ'҄�B�����l^T3�C�t��_m�oc���Vy]�/�9h�; f�f\�,b���g�
sZ���a�ގ������`њ��r�K�;	<V�U��';���أ�w��UpK��mi�qŧWSK�9����=6;�gr�i:6�e��MΑˈff^�$B��f@3�q����4�S諝U��et��3z���	Il���킹V��v��{f�Ŧ:�3���}O{��4���Cb<ky��ɓ�Ʋ��rd����,=5�:���[��;���E��}]��ˢ!U�2S�a߯tt�a�\!B�m>�vͅ�XVl�Q3�dLZ��;mA�7���u�Ĵ�݈(��o���o$�N:)]��̧�h.��L,��y�pt�!��<�e�0��F�˷��S���U���<%.޴�e6㠆�� �b���S��=9�p܆�G��HY9L��^Nǥ��m��&����U�I�]��p�3+oÝ�K��I]� h�(�����8�;X���y��m��r�V���=�ܫ���[6�Ѥ5�]vya:�v�vT���h
��j���
�Lc�]�sz��.���s�w+�n��ΞY�I�&��e_W7[�-�i�2Fa]��2�`�b<�-�8�мxr$nv=.�Z�W�{Ff��c�Q]-CrR]�S��e�]l'��u4n*�1�����A�"�e�`���w@_l8�s���e�2�[��oA2�%l�D)W�,�7/+�-!#9��p��G\L��������E~BQB��H��ID�����Izj�DE��BP�	'��B@Ȉ�"$IrZP	/�!%�Fg�~U��m��P��Q�j0P�	$�D)��!}��%�$V|�U�����~�#�||����0�U��)z�CB�݊W$�Qi�o��8r�	����FLC�KDu*K)ms>��3K�����^��o��z�3)`1�Z�67=�ߞ�k�#{��MC�ء�V����|�2�|��G�/�*�B�Y���K��:����6!R!��n���3i$i��4)���B���PM�Wdg��-~9�*�1V����j�O�س�jX4H���:�fI�N<ҾhW�g�|T��X,���"a醟vVpT������Ky�:��9�ɜ����ć�,؇s{͙yT����t�J閂M2C��i�K��O4wz��=��H�t>�3����,�waX-'�W��W�V��ղE�+��re�TU%V	*��,�G�anb�;N��U��ls�kNSN����^z�C�Goe�J�-W���_�r� mex��Q�V�����5�1��̧5'AR ���i�{.Ɋ
���J�n�^���:��T��UF��4��P�yFg#�Eo+��7�O5�.�q�&�hR�4Ko�b`{9�I�����u^u�ߨ?k�j���0g)�ţ�yA�2*�s�3;u�
���G!kjW(;i�#�N��ƷoZn�Z�7"��;D��GW]�Xli������b��VHwe_��XT����uxpXX�exQ��W���^��;w��s�Hߚ�`�y�c(�M&�E|�O�}}�QV�U�Q�T������*1��<�i�.�^�j�tLkhl�����﮷� ��"O=.׽�蟌&�%$����V�oQPR�x���:#��=�O- ��{���4�;v����o�y�KHWM5�C�g��5G�$Km���x�a�Լ:���d�W�����b��A+y�Kw�[�y��W���^�����\^��@�*@�WB�!e'5����۲��t�b򭲭�s�U�lSȜ�s{�os�Y��jw���j�wɀ©t�m`�kR�k�I�/�<�����w���������-���X�COz���Uoo4��	xT�w>�9FvG*kܫ�� ��6$��V�,��N��ӿ7*4��s�P��c�v��n��s���M�sS�h��D��5��w&�r��vlu��<*s�sX9h�]U��ۛ���+c��	yt��p�s�8�ZGz�dd������Z���@n|n��v#h��$L��Л�^Z��dv�H���xz�:\'l��<�-q���Og���ľ�H��y�n,'b��p5\�Fݣ�g�����;r��0�v���U6�kÇ����������T�xe�gW�u�f��yp�5L��ߎw,�*��P�+��ݥ�<���`�S�N� QE�H6tI׮�|4�RW���/-ۇ	O(A��Zٝ���p�7K7=��X�����;%v�?y��p�u����A� �������4E+Uh�q��<����I�=ah���q��Y�jqy ��n���t�`��%�Aa����.\ě����}ڼ�x��N�إ��F��g�v�0�i\/ɜ�qx�3�Y�w�W�cóӁ�|�U0�UՕrU�=C=�y�Mݣ�E�� :5��1�uu��fplG( 6�,�\�L���{PL�GE��=���#!����vKk5B�s*�A��wpoQsۋ4����G��<~�貮�$�R�Bp�۝����y�`�[����=J���C|�-�.���U�~�݇;]<�׎�+��tqD��H�B��7-�Ĳ&5�}�p���,���d�;ŝ����I���lss⯥��\����5r#��4��"Й��BJ��nT�t�x����r�f��.�����<��*-�~�j�aV�6�7�#GͿM�<�)�Kd��G�b��Պ/t���Pf֝���SM���e�U�2a��^��w|:nBm�-��\g�]��n�� M�F���)�ܷI��z$�l���mͩ�ɐ-�3^.S;�+��&�:�U}�_S���Ơ�6��n��J�]]t�	]�J��D����[����ЭO�j�҅�5����"�e�ຒ�Wz��ȭ�?l���n��w����i��D��rG�����)�z�m�=Ej����U����{[p�k=��Τ����K�Xέ���Z�nk��z�7}��p�y����j�
��}C`^�ʧk�r�=�܅nG�t�_]�ה��e��t(��M�!�'Sܗ�]7�i�.${���*cV�x��S��+2������������^����y�0R�v��Q�Wh��Q��؜}96�l|�^ʌP6ur���;��7�olsi$7x�Ws�qz�v��|I���>n��y�`��IZi��yѝطi`鮮gV����������K�\&��g�r�����{Ƴ+�b��h��:k����#	�V�� ��쿁Լ�3��;xG=ݏVa䖧�I��j���v��*�'A��癵՜��>ɶrW��C�.��U4��]�
�'�ns�d���ZH��+�o�L<ć���q����<m\�cswT7g9^5�]{�ݦp��������_�����=\��n-��F�7hj��cj.�ӎj��N�V�4�[W�ۗ3�詃�q�5y�r��
�IY~}���#�vv�Z�G*�(�^���e/���훠�
a�i�Uley�R�۞��;�_yJBf�S��=���;�6�{Mo�g;�P��bzA>{)ٔ�0V����l��S�&�+�C%��p^�rsO��
O�%�������Ubg��{����VE���ּ޴���T�֢[��V���fr�c��T�P�Ez>��Hwկ'�KwU�����!g]vr=��Q�Q~��{�cG����Ij"�S�%mQ����=��wE1^W	�$Gl����[�{���Eop���z^��~{l��(Ls���iS ��B�)ee�~X�އkuQ���Ȕ�෾u��S۔�C�,��E{د��z>c��̫|ÞB�
�E6H7��5<Tv|�V��h�l�^w��.m���mv�:A��2	�a
e:�:��'�ty_2vVBx"��=�nؔl�֯��}G8+�|��KyAn�-�(�Q�C��OU�E�ȤU�$�LXq1[u��yr�I�&��R��Dpﯦ�J{�����*a`�v���WD�ʞ����>:]�\:�5]�ߛ�VJ'�����1��wSe��^7��C�hdHmJK|��`���Ki&��Ӱ���;V,N�8�i,DM�����Y.����M��R�υ�l�W>�]�Cڷ}�Â�L�BFq�ng��|������a�3��q�i��E�F�L�b1+�ޣ��v��R��]�u!��b���Z���B�4:�+Ɠ����w�VD�A�)ִ}�'2�
���,}m<�OuA��@Jb�5��[�n[t)��j'��EdO���q��Ԓ��W�-q��6���>��ΕI�� n��q�A?d�;ﴹ��S�]Ĝg6ң��˱����u{u���7k���ٙk���.^�����v�<�'��3��5�c55٣�z8���M�,��4;L۸�N�5��]�R����q����6�;q�Йn�f�f�@l�ػr1�{on�NTl�]�:z=D-á�g�Gg��m�K���Y���Q���]\�6��v�kz�l%�-,�#M���]���%�x�nq���*��"���Wa��Z�ѿ��ӎ����S�v�ok�Fݿ{�M�N~�2����I��p�S���g�Jj��v��i��H'H����vRy�r�G��Qv�Y�nyw��ǒ�ɉ'�-���[�y����yJ���"[���6��jX6�f>7�e����վ�jxWl�Y��t?D-�eԓ>���׮�S��n��o'O#K�
�J�İ���3��+ggy��ӛ��mc���U�q��>��-�/���cۭ��^��� �$�'��F%�;'ύ�7�P��(&0&�����<��_�~��]:�����c��߹PĴS���n�Ўnz�o�]+}��N�>K���MD�����]O���m� ��<�ZY�Exe۶9�܅�+o¬P�����f�خ��LVz�K�="Ƈ�e��x�$��[g{�x��p�+�Wnc�9
�k�I"�6Щl�v���v��fx�6"�X�ݭ���mlݡX%���T�"�V�i���Mm�U7BiT�˦S���:����;�y���Y�l�Cwyi�N����(+7�τជ��'��w�����OyCw�����ZuI3����\�Z�n�(�ŀ�+���yѭ�yJ������f���}Ee^8rQ��^oǺ����>� ���۳����g�ՃV� Y`�zL�qx��̬�I|��gu�{�
�|�D&:�/�+7r�[7딪B(� u0A&�
j�z ���狀� $:��i����s��,�Km�B�4!�A��{���I�}ȧ��uxa�j����@,��:�9a��`�[S:ź!�TH�e��W"q���X-[���d���cv�����E4[��1���!2-�E�58QdW�;=R������cYB�6�z����{�\�L�"���?O%�}��؉-��M/�lfgk�lX�=#��C�^=���|wO`�	�n�괇$�s7dx���M��������oy˜�XJY�n�O�<�d"Jm"Kh�Y��G�lgy�j~Ue�V�7sm��^E8)�
9�u�it�>��3U�9(�a�g���rnF��=��o�t�4Ho��:�^ml����ľ���
ո;���=���]u��E�O�8u%�aS�H��gkMAa_v̊����;�q����H���ez�yf<����ρ������'O����zK�T	�mV�8x&Q��70]���nR=��8]>��s���a��,~cՏif�Ce����n���Z̯7ܼ��d�A`b��W�<�/p���J�D3�:���܆��Թ�q�{k�{���s玼;�eĻ*u��9�
H6�����]��%Z��=�ۃk��"��8�:S�En{�YH�U���ޭ�*C��[鮟Oa��!>�\����'HF6�h-y����ns��Py�ř��X���wd���>9�rOM�mʋ��B��m{����n��cB�4�H
��(�Bt[ 4���D�q���)x�����J���s��O������M.�f�ҵ��L�����J���w[\3�iTUQ�m��{Ƀ�^.����ln��s�\ե�@c�p��K�!��:�F�ׁ�k>��;�\I6!�R"���m"'V�F�Ngk�HS��	f�4��n�%Ѿ�\1P�7�uJ\�a6]�5u-����kݏ�짶�ϻ�"�?�
��DQ6�Ba����;���G�N.�;}�iO��Кq����S:�3.#gm��v���A�gU�
�RAf��\+~��lYw-�\ٞ6˙2�m=nqBq��&ƫ�����\Y�ͭ�i6�q�`$�w��~�{�m�Ď�׻��uvc&���� �<�U��
>�:	ܷ(�2�|)�]���*ۿT��S��p�{އ��z�@-��]�rL*⫶kz�sT�.�=���7x��<}R]:����pt���Z��Z7w&Ǫ�8�]�F]����4�M����WW��+�8|�5~��U��������U��n�f͊�m���G�>m�>�j��U��]�F��y�z�!9����$�`3�*V-�[��W��(`�U;�6��^���=t�A�=��4���e��t2���u��c��/u�&������c	(�"������^��x�Iӝ�\?|z�a�V2\�i.���u��V���A.��^�t�.G|k�ut]�J�ec\�v��4/�b���oK�E�%^�(�W��l�(3��Z�}�1�4m��{�>�+]�R��XP��=$�ݫ�Vr�����!�v��Cv��\c���V�Ҏ_i��s8CdE�\�W�uv(�>��>�9˻k��j�����C���H6�e����Y"��CYܵ��]�p��/�х��x�ټ��k�f<A�[���:���#�j7�h�*T�i�v[�ή�����c"�2�DD��oq�WΫ}�k;(�� L�nC}G2$z���4��\8
��e���M6ߌ"OjtF�O轹+m���mY�b_*�e�.�
�:�ͤ�a��[M�w����h����6	�F���9V��P�����й[��]:�k��XZ��#�b���)�ڄ��ӆ�g��]���s�}��N��N>��W���	�.�N��pې�8奄�����@%x����ڪ�Mk�@�-�ݕ�mS�V:n��D򶭤���8�Y�X���ܥ�:��Z���Fҙk)$�XZ��[��l/y�3H���p���J�Y�e��2js�c#����2�]�"���k��
r�;WԢ�����cwM�\�ֱ�5}�2s;!��D����	��ekj^�/����83�<�]3ka�s4�q�u��Yu�jeE���@�$��̇:.|�r�Q��^(����Փ�\�NX��f5���(*�
;iݎ���c�v8)��)��F&�:^s������q}ce(�"��l�{f7��V<nz7n=<����x��S��� ����N{�;wX�G��)��m�m7om�:�I�Z�t;�Q�"�[n<�x�_n�E�-cu��X*)���:���=0�Tv݅�s����V�W<�pH�����:"��G*�����Q�'hN޴>9���ʘ����r��%"�&F��b����uomuˎ�v�#��t�m�W�X��Q���>�<�y��$q�u�����7vr.o[�$�W�u:�v=�O�ٗm��p��p-�-˸��W]�We��:�09��٤t��ה�0p�.��w��#&0D���vS�;V��7&m(����s�\[s̓&w�v�폜��{�{7<�s�ǝחt;��`۬l/8g��kh��ú�n�=8��\�<��5�4q��{t㞗��p��źݧqnM��=�\Ɲ�q�����vu7h�&�]���aDĶ��=��*����j��k�p��m=Rs�F�-v8K�Fu�\z틝r7m�hX��n�sΏ7\v}v�Kl�y��<�ynL���wmdu���aK�m�t�>�0cZ�3�i'�Y��ٍ�ѕHM�:w;�����z��:��f
E�7n��6�B.�ѳ=���q�n�����m��pqns�����������s�Av��6m���.���	�n^ϓt��m��v��ƺz9�qf[�Ӹ��f�ݝ��2�A�8[8��.���Q��v�a�Pc	˴8��kn���������<Cq�k7#�:�]o����G������1���8�Z5��r��:�磥7bζ�q���O�ф�=�K�7�X��]:�������C���O�P�\n\p�7 ��6��L��<Tq"�s�N9ۻqs<�WƑ����G9Бs���#p��v��z�@��O��b�J16@cJ��+�S=;`-���+'=X܇��	�?}������6R�m�n&#�w��˱A�Ży��v���Πf�tn��mQ�p�����ɭ�Ю�5&�E�t�ͱƩ۩����g��;t�Î�BF�[Hu<���y�rd���uB��vbxg�=�/F���q۲�����Z�d���D�Yn��{<�h<Xn��a�&ͻM̏6.;F�ZL7�xz�v��Yv�룝�:LQ�x�-�m�!���	Nzy�;n��θM�k�\����:�2E�U��3��=;���	z����ƥmל�Q���;���h�6�g&���;�k�jk��j�1zeY.��^!���I�T���<�]{�]x�Z�+�٦�O ��{;ίz��.�F2�')q
.�
�6���R�=�]f\�=�x����(`�����i�!1ϧy����犧�v�\d�;��w����S�?���G�!c!Y*߽w����q{��[ls�6�s�6���J>4h��D�w���b������mI.�>����s�6��n��L��W���8���"]�Y¶*�~j��}4� Y�G�[Xx��	�3����y��2����9�Z��Xp�w�Q���,u{�'�o��w) Z�rg׫�)Y�z��ٗ��w�l����K��^Y��A�e��N7����3	�i 
����nw\·^!#nG0]d� ;`��=t�,�J�Q���o[K�\��^�@�&���W$�E{2�@ix�o�C��Q�-n`�?H���^�p�'��u	ւ}X&BU���Ԧ߻��$G�����%�{��4�����3e@?D��q4Ogu�nʏ׃=��1z��N��§g>�wu�4��'Q�m	���ScO@aHбV3���SQY��KXC&=�8t�p_��>{c�j�X�T�֨���N�@a0[lS�m6�������z)N�l���J�d嫓_V=^����IT{^o|�ֺ'�=���J��,v_����Se:QeGo�U8�L��[aο�a�)������}(랖3��^TW�ʼ�eN�Ok��y�+��� ���~��T��Z�9be�Ӽ�wuww'u��b¨Q����tϏ�s��*0u�zm��9GO�:���>��V#���ޟs�ş���'�-Y�MS�)���}���X��<�eغ���(ku��\�յ�J�d������w�yL̹0w[��+�G�,�[�թV�ou]�(b�3�%b�3$�w{�
�ϥN���bZ�7��Rv�/;|�+hv'vRZ����U�C���+詼G�}{�z�N[�낛����}��\k��]�l�M��/�X�]�{��2����*{�|%�_�t��u��U�<4H��ʙ⻙�������v���[�t!3^��p[sv&o],Fki,�t�w@��7D�Vu�Ŏ�J�4:���@sF0YK쇤v��K�r��۲7������f�z\�K��u��-2ցB�)l�͜k�X�嫯kw�G::��n�om��8�[��8�Ogn����:�z���=�P�De�oe��* r&T�)��gw7�����(���G3�(�R��0�\ׄ���p�Lj�%^�SnfJp��S{�`V�H��.�ݔ�N�#��Dt�.^z�wX�ٷO�	Ok׮�lB�1��e! 2 ���*�<�׷*�Y��_����Hh�\�!���lk��R<Gd�Q���J}c��u���2굔"����-t.�!�z�km�_�3O�W;U�Մeߵq粟�٬z5���������7�vS�ոך�A|����]�7��)SH�m6n��>�-I�;w����G���ΛBΤ�3�w'k��Iɋ�G����و�]��f=Q(gT�0SA�I��^fd�E@p]G����9=�^�YIÒ��:s��̝C���1����P�y�6��rk���#z�O]F��V-v Ч��v]�ڝ�ں���s>�3**5V��>�[V{�yt��ރ����᫋6�{����%N��Nʵ�A��2��w���z@E2|�#�^��.P���@�	كnpϠ����[�0�1�c���돼�g}(����^t���i�"�9]p�bj�H'�x��9����vR5\��w?ߠ��m�5��i��+�B�����/�՜+��Q�ײ�	�������O�q>�_{�Y������ME�\�.�Rm"	L�I���T�/���וy|ҩ޻�������3�+�"}eJ8	&����mJ�S�Awt3�-�`�V��(�lS��^.x�ݥｪ�����2֡���~�N�Jug���y|���GŹg�r�c�S��z�GW�3�>���Z�nRH��J����v҉���䬈+��e0����5�}��g(�*{1�`W��d�<԰���0f�z�����{�S�� ��Pm�⸐[C��6�h+ʊ��;}�\䶼��]���dO�_[���2�)C^}F{Ӹ����u��*|mqO-OJ����+Z��3,��66������N���,C2�^;r�k��ĵY]>�(�3n��fRd.ƇҮd�͜���5e����6�ݷ"����st��/y�nL���s��rt6
����8룢`X �8���um�\���s�im��z ��y�7>H��Xc�n)�E���8���n���"�'��Ka	�s��m�e�B�����Q�_�z�o&]��ֶ�sݼl�Ya1����k���=nv�lְ���Ư87����B���cʦ]��y��PEucn�T�Ϟ8����3%�Avn+YN��*�n9[Pen������3���qka�X/��c�ქJc�w7��*y�����S�����qU�X'�h�2x\��-e��JIT��z���[�jGn�?���
������'����'�v���*�ף�ʍ$q�����0y����V@�U&r�����XRM���xD�q�Q��HbJ�D�wJ��������[4����#E�Q�<�Kb����RA��R�k���J*��-��4�/I�]�q��
'�ӧWXN-cG��+ӾP�	�K\}�^�����n{h� �h+�1���"�ML{O'��^X
�|Z��"�$���w�ʝJx�����h�x��<<��֖_k�Y<�-��k���M�5!�ʭ�W0�X��vM�x֡����Кt�gd:�7]F�mێ6x[2������ܞU�/v��mq@D6 �Ձ
�]�o<
r?��9/y���3^�k�`A]Gf��4v�K�_ =�Y��P���S�W��fz\Q�
�E��*�m0n��ۛ+<�I�����u��r�<L�*;�V�����i22�JA��9L��=�l���mR�y+��Y�u[tڡ��`�1�@#nC�,M��zi��3n��\�<����9�(����w\��������A[�gx�oAz�?unm�$U�h�R)Xr�Rƨ�G�|����=oz�l�N��Yw�Rv����W�Vx�f��BS窂m��eE.��ugݻ=Wq\�횾V2�HCZ�U,����Qbά�[�ǳ�u40e��}H��+V{�T�ޒ���h��y���3�t�c}�V'�[3z�-��s�m`�v�?x o|U�T@�*�ǳ�l����Txa>{��tҥ,�u΀����{�[@Q����t����%��C�����{��3ct8x>������g��!ςd�E���������Ǟ��S%��;(���&�a�C$�:�셵q~mwv+��t�����V#�i��t{����i�e��b9�E'gݖu��E6��;�[].���`8��_��c�4�-�3��B��M\�ۤ��e��#9�>����ڎhU��0�t��T�7GU��S�`]��>W���n��X�,���oJ�G��.��T����؝�a�8{�]Zt*4���˹����L���s�z,�E[!������m�mf��$�v)f��㘥_2�^�-u�NĒ�\�v.Ρ���hj�"���c������]�W��n���oL���!_Gu�Aa �)|�&��UM�����Q�]vV�}���T�u!�,�.b[��J
��޽ٺ}�Sa2J*���s����� ���1[�3��!-��+�ʩ%���
蓑�����M�.��ňZ5����|���q�h"� ��`r�ם�""�����Y�>�'*J}V����A��z���#�u����<�S��s����خ�8���-���s�]l�t����.�XCd�8:e/`B����Y��~�Q�/�����پ��>Z�z
��8P�*_=�Y[�ِ�h�E`�;᭐
t��m��i��?V����v�βr^��y��fn������o�V��EA,�"H�Lϲ����E�{Ǘ�x��s������V3#�>GO��L�ʝ&]�h��N���fi0zݩ+4���!�������w�d�4:��[�'�̀QT'>��B
��^��jH�N��H�T�m�}�A�`���|z��;k;<���)�'dUS����������U<(��c��~ۙ�y:�}����	5���U1XU=��-Zh��5� ud����lmjz9���I0�;S��d����uU��X�̜A����~ݑW��w��臺��G��j8����%���ux�F�!A�����y��Z��:d�Ϯ��ʮ�V(�Ȭ��1��z�[�{���z�^���';v[SQ4�q��%����4q��u�;3ۀ�6��v��f�����tvZ�Uup`!���'tv�<e^\�2��X
�J�w�3��#c��=�f_��b���?,ɛx*��=�NԹB5�0O3�[�D}$�+;k�
��x�tB���Ra����jvR#�y�p;~~[�qX���~�LzUݺhJ2's�3��^������U=j������J&�k�Z�՚{j?�F�1O�����C=p%:�9����l�c���������#�_����X����o��ᴶzhZO��S�	(�	Wa"M"�CX���U]ws��k�r���M
����^~�3녪�D��jx�Ni�Z�>�8no�ݦl���oN�e�������V���X��l�)�İ�z0���;���WP}5�+c��.SOo �^]yLa��IG��jwz�^�S4�5~�|3�X*Ÿ���yG����u�*����^�XM�����ۇ�JQ���ݺ��>�aٷ��׊u\��7���a:V#(짅RFH���n�3ln������n�l��3����q.㬺�7h^۳�gh���7n�㰇%����Ξyh�ޘ7[���ݶ��Q-���w����Ƙ�}]��G�room63�m�k���Om�l��sێvu��8�����㷸��+���c�7g+�Z���q77����\<q����xl�7�c�:�nݩ�ˣk�9w>ۦꢋE��M���=ݝ��<�u�� ��k�wl���c��rv�D)��ܣu������J����۱ma����YY#�b��_�L�MF����x�n�EnSu���{�z�� P��|��ȳ���9�`L��똫Ni����m<'�>���a��)�A�M'X�`x�
#���}�������8t��{eͤ�	9ڽ'��i�Z��~8�]Mùo�l�\��RMw�%����{��CЭpB)l�ko�Wu�7b�A��\�L�Qƣ�g]J���6�2o/Yw����7�H�t�2�\�J˥����}�Xb(B�d,�\��B�$(���%T����ut"�QnTL	Q7���ky���Nn�Õ��3���b��a�w�~����!�	v����ן�m�21�T�b�1��o	�;�<"F�<HXk�w���*�m��^���&GR��EL}[$��I�K#���W>��ɍ%�3c���8���4羋���ۋ��uQ�zN�q��v��;Kq������mCuV�/����V�������R��N��w�*�zu���wJ�->b7X�����-�m���Ʒ�S��zX��+V��qU���Z�*m�8K5��$��x��7��W,ڻʦW��yxߪ�^)���dr��25���a��S���}ۼ�Y��&��*�iC���SKv1�O}HW�? �4��g�p��D5I��ߞ|ݡ�y������vF�+��px{yj�0+����m�`��u��1Y��ca��u7a�l5��/0�YA~����p6���{e�;}l���;J����/Y���F1�c۹����h�7��K�Z6ʍo)UB�z	�W����x̹)�9RmR�үb��;n��n��;�l��zQ��hڮ�1��J���_f����p��[�,�	�t$���E�1�QF���U��!LD����=]y#�V������G�b��;*d:���Ŋ"��7�zn�*���m�GsrfP�>����:�(�s�=q�O:R��a荎��b�9�O<�nq�=����k^�j��X1���߰R5�1�쩢��]d&��z۠��1�(��DQD�]�Y4c�yPG
�f�tBk�[�Yc�̭t�z�`��V����f�� �)��ŭqe9~����>��3Y:�`�	 �O�vJ�Y�d�M�̙X�xu;ѽZ1^�Y�jsS�3�Nȉjj(��-L�7F����#�y7�q2�t��T|z���|f�����Y���6lY�	�칒����s��"���qೀ�yd�ũC{(�ۊmLK$W�[�d��*�y�JA	rWV�1�hv�ؑ��O��t�PD�r��Wf�/+r���t�q�b�F��i�5��M�(H�.GL+�*լ��d������S���N�*��t�&�*=�9Xe[���XkCf����go-�*a&ۃ�Okx�+3U�)�q40���D��I���M���ʦ��˦��]M�/X�.�@�ns��k�����^����H��jw��B��M�ŕh;�F:x��ԙ<�b�s-�$r9�:bj���M�x�Cz�y�M]qU��0�!�j.�
,�ӏ$ 䶆�o
}�}�;\���A��g�\�㝔ku��J$fWm҄T|
�rŊf�ծˀq�(Q��:����뒭ʏx+�71�qᏫjA��-����t�zVW_�uI$ h�RǀK>���cBB^����W�Md�D�|���� Y�*���Sc�U
��=����*,_>4zV�dr4B�gW��Cu��Ұ�h}An�m�{��o����5��mv�s�1�y��)ohG����"Ro$x�Y���BG�1�#A]N�q�p���֡��m�p��m��9�sb9�q*����!Tw�a�=:�r�֣���Z���Ȳ}�o���,�̼�_fH��f��1������ֶ3c*�,wR����1q;ɬ�;�Wdvܭ�W+�h�u,ՠ]>A���g���#����c�"�+*�ׁ��e.?!��tc�#S>�=r��=�ۭ�r:8���0}���>�V:� ����ݛ��n�۽��rK�0 (W�۴�Ǫ�j*�_W����_�}�sڇ_�e��|z�eY���%b�=4�*��i@Ua�N �O�����3�<�B5������G����n}9���Q+�yJ�y�-�m����^�.�*7�-אU\�.}nu�~�fA[V!_���v��l'd�N��>�^��W���n#n�o�[T��J�-��{�bv|��\׽�E]8l�@Z4K]�ymd�+3��v2
h��(
9��]����V����N��E��[����k) )$��%YJ��F�"_ ��?(ę���:͹��[LTHvC8��w���&N����i��c���t+/���D�k`�N�oz���~m �iIm3x �K���Y>�=��&4c��^��|�n
����Εk�'`���vV��#J�>���M��>�+�c�G�s�q��nJJ��҅/q⯇5�*�O;~�9cb��J�o�{jz�8�ioIێ{�������D �4���6��oh�������K�����E��b�t�ma�9�^�n ,qz��yC�y\�.���Z�}������� W���ϧu��Myq�4��yf��
1;E�)������K�����f�>ɿ`�+�4���|��ɛ6���X4�~���#t7���^P�Yl��&mF%E��D�Y��;��^	�C�*$�=��J�V�u�1��"nw']Xӄ�=�M��f�BVD�jR8F�e^Zۊ$rPuV�vU��HL��R���ѝ㓷ʰhTG��,��0�uIvg���5�8Xٶk���zGv;ƍ]��s�°U2��&Z��;ض�5��;��9;{r�G�+E�L�"��-�}a�T)�H
�c����k ����2�;4I�m�ʠa�AJ<�w���&�m|mև[{A�b�����g	��k}˷�~DwxM���n�����ΟP�����8������^�0|*k5�ޟ�k�R21��s��b��:�m��}��}�S�I� 9Ԃ�(v��K I��*�D��=/j�^SZ,S~���P©	�ò��\h��֎h���X:�),D���Oa8�S�N���Z�
x��LQ��k�&���K�,f]�k�����aM�;����׷�T"a��ۻ+҅�NuԡBu�ߧY�=�+5P���Q��\Ԡ�eN�ݗ����woFUn�Z���^�8�\���kb�2�|干m�ŴK*��E����&�Q�(En0���h���o<�3���Ϟ:��) {6�!������f���۔M��n3���m�=���'h�����"/u��yu%��c2�\۞�Q��4�8�Nݻϵ����G�ۑ:�={r1�<϶�Ӱ�ۮ�-�t�����\&�]�ͻ���f�u�$|�m�]���&�v"vtR��A϶5sg���#���v��P#��k��m�Jm����3�_�ۋ�?%�����L�NR�d�Im��֞{[�zZi��~�5=�|�և�1�ο:x*i�T�]Ƥ��I���S���B��R�\T�>V�"����$jh�hYI)N>��
"�N�T�����;��B'Θs2��Sa�(Z^#~8��i�i�Kb�Z}��?,���R�Y��j�Rs��<��U���-׫�(�ݐU���"�u>v|�d٫����_��<�{���Hk��lR��=ꛆ��b��؎���9�q�~5��|%��g2h�8�}X��%X�����P��кs�n��h�5�~��~:�1d -��)�f�kչ/��_t{A�Y׊����ː�����*ֹȖ��I�EEd���V9�P����E��4��u:j�r���}?W���P��,���`����D�6f�S��W]*݉��P�߮�=ጼ"t�����luv{l�a	�����"�d3�"q��a�V	����~�G��c�B�zV\��[�D�T����u'M���G*g�*Q���%�Og�^KP���W�1}�ʒ��Yo�#�)I#^�UDݶ�Ƹ���c�7I�F��V��Fc�.�<$Ѻ�ϼ��%>����5��E{�&\du��2C� �0%Ƴ0��k����;���UR�2�`Y���%gu$D�LH/�S�!��6��p�,Vm�=^��6���S�����8�(J��E��6�rp�h�<K5��M�y3�O�=z�;r��*��%s��ϳz�?Q�a��AX4Vd���B@�H��HH��p���ڍ�|�qo�R��c=�˷k���n�3$�*ʘ'�c�uc 1`0���Ω��00��:;YK���h�۽�[�*�E
�_�X���emP��rSH�%�ʪ}����ۦ+����k�;�.���~eU�H
�u�c�����R�4��u�ޫ�5�V�S"I^����P ?�z�Qxy�Yױx���c��뱺�0����pk,<@��Э�v:̎�z���s��U8��Pe�)�E8u�b�;���ģ�YOA�eU���=��OKsy����.x=K+(��`5z}��OSC�4�t���k�4��t�g?�T�u[����r�82)�Om��ԭ,V�U�^�Q^Z���Ѵ�'����e�-r�Vlw��!Чn��*���<�T�+���	)������jJ|��뫂�MOE�ɾ^��z2
�i�^~n�٢���`דsΞ����ӣ��)s9��a�[��cb!6�v�C��>�=��!k^��M�f���Y�4�`r�8ϣ�ڕ�U��k��6�^T�0ة~X�B~�R�w�H�>h6�4ٺ�jT�HV7�N�[a�b�a�z��h����5V���Ń<d��xR�xt��yO��R�7F�+F�-��
��V�>�ٟ!�Es<^�^ŪH��դ�����p���}��3��M`�C��|�~�w�q�� e�x}��a+$|�����{�����+��*�����ϣ|%�#Ͻ�Ei�m��N�2�{Old��Fn�b��j�՗���poA& �ck�l�;Us����c�O��(q���CZR��#��_����Cw`"���T�?g|H��6�|~�P��`�YsX/[�օ,����{i�b��$+���_ܱĻ0qP�<�un��{�ҍ{�gCP*t�ugh�0S���A���[��(U��~:�	�٬�~w�z�E�=}�������>�[�jZ�'B��kk��cN�g2����j�/J�Z�d8���I�Cy�:��9���jo��C�E 2�y~b5�޽�QD���7@u*=�
�_������+,�y�TF��W3�R��ft2���}Y���?]6z��W�E]�������x;@��P/%M��ٌ��Lʔ'��j�b�=��m���@�����}��r�j��sjbJ��;A=]���`�/�-�R
q���>>ד26�RJ��hğ1���Y��%���[)�R,P@+)0�˼�%��J�@:c�m�AH��k�<��*PP����`=��t����T�t6>�j�zV	'�־��RN�K�ӝ�t�4��X"��,���%`���K�K��g�JG\m�mv-bXWL��`瘦�q<�3)��Σ��;��QTQ���Y�{��g�>�D�ͧ-*��nT���'�1ҳ�|��Ҡw�r����PC����깾��vF��kѿy����V!�Vo��-�8�a��Y���ØhO<�ҽO|��E;�[ӷR�� ЬTj�
>�\%� �d�^��[j��)��@�[���ڏ�u�r}̌~F����,�"����+��ﲥ_$0�xFT�
�*���=I�=Z5P��z���p�}»���ς�� =�t� 8��u��}�f�h�lG#;H�K~�Zɜ2��.�'���L�ޡ���솙�s�ؽ��x�5C{)�U��\ih�Y���c�e1�
�r������U��-�IQ������0&N�eҫ�{d��X3�n�� �>a?s�uX#�N���R��5Z) <�o��9�]h���L2i�F���� {E�^��jp��4��Z�a�=l�a���؝e :n'LM�7�o�B/s��Uj�k�j�㹻�g��C#.�c��߿ֻc
�r�n7+���0���p��8�N�͌A��5�9{8v�[���㷫rk;�g.�:ݻ:{!�t��v�<�]68)�6皚úe���wm�[g�mۜ��6{�T;/GY��F��/:�ٓ�\�po^y�h
���m��:�˙E�6g���9���ޮ]m�-=�:c�2�`݃�ጱPN�UTi��>?e̘�i���'i�(b���v5�:�.,{X��\Cq�`V7�{i�cϴl�-so��o�[���[�����*��jbⷹ�c�k��KP�*�E����ݨh���2{;�]�kˮt��iC^���4)a[۴�z�l��վ��u�*<��zZ��H���j����� =;�Ŷ�t��o�_�@����gc�d�(����~P� �LT����V)�T>A/����#~w7TU�(�΢�����k�����P��c-�w���d4%���e�c�ɛ��;����bBmm�����oM3!_�+�L.{Ԣ��hu�p�TçD�����$��n��Y�܋b
PVTYim�XG�+�@�^��]�v�ک���V��*���t@Q�ޕ��عD��hV�����o�Z�g�[�O��}K��O�	�4C�^�?8��p
%���u��Z�M�u�s��~�W����	�M�LO��;�uΕ8�z0=�)Gm|����2GoJ��P�j��������;OH��r��V}���x��e�V���<t��=�9�0�ms�\�u����4A[/�[-]��^ѼB�ȫ]�}�S�Ϩ��:��˻�}~ua�g�Qb]7�}/�:���M;5.*��A��w�����!�8�l�"�N���e����J<�3G+跬!V�R\[o��Z�c����֪O%J닼��;ǒY�ne�(�G�=��˥�Pe���n��^�+��o3#�p�.���k��`���(�cm����3D[u�}xn�#�銾��r+�kb�{����s��6YG4�»Lp�{��ª�*�|a٠7;!��F�r5N>��>Bo�r�z/�m�7պZ5;5Ӭ
��u���y%zq*F�m��|t���ܢ'fi)��("���Zan��]2�ڇ$� j�Է�}@W�6�60��$�`�*ˢ�~���F�g8�
�&�8Qy7V���n���3H�(LԮ�5���u����m�Zu���*�Z���p��M�8���ܚW$a�d�o.�\�ɽ��ohVְ���mhШWa��u�f�����L?vOm:�Dz[�=e�wb��p*��/.�h�h"U#�4h����X�����%g����=�=/6.�s7	f�ˇ�8���KF�CR�Ւ�y�}y�����ՙ��<iMn�u}1������F��r���N�����*�����k����B���eJ�_]c_2k�&*����^Dea��Ks�^k��\����ua�'yG��]�L������T��T��T���/�aI]��ι_��_Z#�L��:�{��Q�����a,u{G�}�X(u^Q
�4*�m_�{Ε�0Ϋb���<�*�:#�cY��<.��T\��|�Lw�#\�hG��O�� *Ҕ�iqpݢ!0*�y����M�;����T�v��$8�e�]t%���zr]��l����N��}u�:*��p��#遯� ����b�VK�����dZ%���R[+֐c��'[��y�'t�,լUDxA�␩;�?YQ
v�.����eny}L&Xu�q��A�ܬ'2�_�u�+����』7q:i$���Ĵ���MsZ����<o��gO�Y��v}�g�?n�<ڏ=��+�:ؠ�R	j���E_�Wƌn�;��P>��P���*���x6ԓ�z�槖�LN�1�n�Ps�'sW�#xN�<vj��b�O�j��~�v>���F��U�9������Y�6_dXo߭J�E��#�̿�v>�cw|��/�^u(iY!��o#O��0���'��X�ծzB�݊B��b�B������%�!Dp�k6���n��_M-}i�i*���W��B���� r�MTF�@|ɮ��eu�1}�u�N�0Oz/��ώ��o�@��T��)�a��a�HMԫ�M�Y��'.��*�"l�6�!�������J4B���Jt$ggW@�⼖�v�Ub�J���P������~����|�]cW�2�^���	7{��4I9�o�}_OU6;3}G]
��2���A��*���yT����N{��Tk2��dA�;�@]�)��v��b|�D�󺎼�t���ǽ��u>�kod�ǳ2�1�'�+�*�����\�{G��D�S�/A����|r|�֬��l�W�:�z|��>��M�ЌD����*��!$��J�.�i���Tiz�e=�Pu·5��4t�$�c~b���D�+|����2e�R�j�L�E��t6s;MS�m�~�{M秶w7V�-������p��E,��_9�qx6U�Q�W��y�6�i8�����*Z��Sh3c��
՞[ʽ�>{����U�ۜ/��������5}W�\fq��ͺ��
���%]�׀���u���<��Y]]�^�v����W>�_�>>}ao<�
ϴN��d�
��Y;;�G�Y��3�X@<��l��n{P寃��
&�0V�_w�Jg4/�K8�{ҍ@������"˦ I��lF.����bŲE��0v�n�]�HBkQ����T=�3A�F^�n��({�Y(�Y�����*�Z :�����g��?(�բ��Yl��(�h{��ןg�����M��j��绌�'�ޘ)65�b�"���%J��}I�˪O8%E�P�~+k<8(�/Q���s;����.�/���@�h-lL+	^�Zh{��kv��s��	���6�Su8WO������Z�ġo�5�����bS^.i�46X3��9��Mu��/"�π�wH0�]��2�n5�F$0o�r��b˒��n��9��M�L�&f�ݵ`�sx�t�PDFΕ���Zh�Q0-C���$q8j�T�u�B���q	l�����OP���8��n��m�׊�I�/�Ig[�ؓT��!<x���Q��έX�دq��;����ٱ��qFm�:����9�8SZsrmm����D�vj�*u�I-T��re���T�*�/5#��^�u�r\ѩ*�ͥ�0k<M;���I�N����Z��u!��N�A�@q��K&)�JlY�����Y �����9[Pi]l��K�Ȕ٧W��!��ktm<4�S�q�\iwK����I��W�����t+��=Pt���qi��$*TM둽{47�d�u��k2Wo"73�s5݇qB�[��d�v�N`⸽��h�sIH,6��,��X�EBvQ�0S��7rd}��m�-I�Y�G���落�O��<-���l8^?�ŭm��)���S�Q��l�;�G��l�����m�Û9�|8�d�n.��T,V�Wok܃�
͒l\�ĳP]
s�ĻY�8H.�0�:3�.��u�`]|�m���N[��ފ[�ג��i�KY'*�Qǽ0S���qû%%u�Ty$'Nޟ=ᘫ)[U�i%]7+��0Bn��f����$���<yW,���6��W���b�e�'��}|V�%uX���B�.�'���]�{�n��
�8�t3h�\��k���xpЍ��tE�i��N�r�q��rk��ۇ:�z�m��%���f���P�
C�pk�1g�D�_d�g;�m�l �iA;S:�u����%���l�v����ch��W%���r��z:�o1��q��	G����S�noI�v�k��GqqE�a�T�tr�5sqԅ۷��s8�|�u�!M�@�g�F&@hE
�u�5�^�r9���S��\�]x���jz�L�;�X��}�,����Lۓl1��ݻ��-ۏF�Ľ��ts�wC���,�';�\�;nڱ�k�Fv%�̝n۬���[�'�O5�0�9ܛ˸:��Kq}�ɝ.�b�0�lciH�㬧��z�=��ݝ'��"�4����-�"F����,��vG��ָ�g���۔�������������;�Cs��:ܼ��7 ��ݍ��v���̀�.���\c{��\�.n��p�'1����ֵ�u�^�s�mڜ��:�!�t�s��˻�=��D��b6֟Es��py��{\�u�g1��w�F����O4C�4�x�Ϸ]���0s��s==jݞ��O	�-۱�T��s�p�0�g��ǰwX���e9���r;jy=��]us����Fw7B��q��@z]�{vM�n�cm�v����v��.���1ӻ\Y�);��'8�*�+1�G[km�Z60�����A�9��{<n��Q����A&ⷞv�:b�ۀ�<�.�d{p���gb��5<�ƶ�ts�W] qҙ�=��������qN�u�׷//Y�vC;!	��^8�7��\쬳c8<͇��WG;���fݱ�#���]d3��^y.�NS���X!פ�b�A"��]��'l�d����/o�c�Q�s���^Z�g�U��#]�x�,����۷t�q���:��v��1��`�㎝��X��n��p�nwc�;t�؎�#�/���ۗ�lۜ��F%�h���гeC��E���.��
ʆ�R-+���pL:f6�Ia/�e�H��wKs�����n1�<�.o6�ݴ�i�e�z��=��W]���QՔ��=�s��o=�������6\��O\q��I�!���v�t�$��v�][z�g�֌(t�3��-�7h�<p�E�'�Ů8x}0�K����n��y�m'$9��Ic�k��M�ƛ�0l8�뛍6�5��u�p�s���܋F����W���㳸�cn��q�6�nǙ�n�7��{im�&�v��9z���q�k��=��n*N��aa��VMs2������l9;%^�Wf�)�lU.���O�=}kL�n�3�E6QB��V?���ቋu�^Li�u�j�=�Y*�j�ץ�Ѣj^R�}.IA9Q��2�6�����b�Pۚ�01h�7����zS�B��cpস烥�P�o�m<X�8:x2 13T[t�)�����K�������Z��=��
����������~3�2Y�p��9���Ζ'��6ߝ-�ʻ&��0�n���3Ni�R�mL�ו�>5��z��~��sI4�NxJ�M�J����g��Q����#O�yJ��Y辫 ������E�7h�w��t����3�R>�M_�i�m[[�{�,����<��e}��7�����"}Yx�:���չ��Ч��u��"��n��Qx���+G���Z��f;�ٜ���_������R�h{W�P
���mk:mF� ]��;l��{9�}����&���s�[a׶(����z����f]o�x,�T�_J�+M���ɯOn�07پ���饍\F� R�|ff��H&Ա��ֻ�H�-r'���PS�|/ls��"yKW����k/�A9���,�Q�75m\lةGskm8��\��Z@F�d�����[@��ԁ��.��a5�ˀ[�ܶ�.�!�⪳;�Y�iC�T-���[3_�g�g��^�^z�*�U�V֯{|G�o����{!��~ЈV�
�SlO�g�sB��8���}�W��W����[uV+��t�|��C��S���Bse�+���<��D}�� ӛ>�j�������J�q�mZ[L�j��d�����m &s��Ss�/I<>�0T�4���ǺX���2����{ɀ(
�M�k]�Ƶ�eΝc���t��q!��S˺[�"��R "m��^�DQD������|g����6пn����4����[�'o�Vu�P�s׫U1K�E��Ѣ*���-���\=[\^��5�6�k�9]%A$��OezD3ٷX�'�����֟��z/W[��Z�RW@��i�F�3O4�.F�x<��oꕬ��E*Ȯ�T�ܝX���U���4�|_�>�y�-g����>��N]��PH�],K0]�!j�VJ�KL��������>�{*U�r�]�'����G[�s����I���B��鮬w��Q�f��:�T<=�k����O�J����U��@���j�<5��¦���U;�s>rߋa�J�f�����q,�:py:����V6�M5�!�@�j�Sy�f�ٳ�&�nQ,ȥ�)���ܼ����f'�_��Ris��r{��svWHv��WFf*��2�[�HiT�u�O@lu�TZ�=�=89�yd}�ۊ�\�>"�<&�����J��)�ڻ}�]C�`���eA+��}��$� E�ҳ�.�HmYeM:�%����5v%��;��^۫�*[(�cʞhs2R�}$�ٿ}c#_6�<�T4�;�C�{/�"�W�X)ک�Fy��;��AP��[�K��W���̅<YƳn��n��]s�;�4.���At�H�F��u���~�GyX��
�/9�>�����д*��]K��%[fX$�J���Y��1�c�S S�žh3���h��9؞����R�R�N9%{�^��#�:�o�	Uu�wT~峻7=�ա���}����<�X�B�L�*U��C�k#�ҍ�	��Q둑��i*�InB|��J���CeQ���z�������T^#�]/�e������:w��u��,�;W������e����'94���f:fdD�`��]h��z;�PNl�ޯ{ uxM�H���I�m�G�m�Y����b�E´���q���Hi���}�x�N�@^Ƚ��v������=ҭ�nwN��KTIxNq]���]6�TG�!�>�}{ĝoiѝ�on_o+Ǉ��*�&���c��R{|)��S)�^�+Fo<�T���UBЖ��������$uV*�Rz�+v��6��ڞWw�:��ҦU������\��7��+����l�3~ϩ�@����W,m�D:9�n����M�t��<�Iջn.�e{{�;\�׮-�GҦ�*V��+�ꔴŮ�N��(w.tEDjèS��r�>�*�[�^��l
���WS}H=�8^:ϴT	e�.�s}�_*�>eT��魂���_��xuz��ۗ^�s�n�*j��ף�/��}��,ށ��9Z�x,r�v��
C%����S_�#{������\�D���~�R;%&�qZ$ڽ,�3��\ު��]�Ą�LQ�䮞��WR�^P��p�x4����o]xUK��8WZ�.:��;̞�dQ
E��B������7��YBO���1'���8Vᦨ������ї�� ��H|�]����%V�A�Ċ�%�)�{�����k�a�0x�}^Xir���Ĭ��i���d�|�<�nR�]:�:S�Fſm���<#Oi��u��~��r)X�j9��9lUb�J���cαC�ID,��V�;��M�h@��Zz^��Q�a�e�5( �{���$T�9g	N�fČ�p��s���/-\�ʻ隶VԒ��;��D\���6��\�۲���\]N[w-�<b�^�OF<x�F8�C�cZtE3[��Me��xǆ{��P�qv�tbܹ;-��m/m��c/G��n]#Շ��qGtq�mq�m����m4R����� sncc�,u�릍�E����E��ݸn85�����Y^}����a���+u�Ŕ��)n�W3���Fk�6���C�=v��y���O,�;X�諰�n�v#�i����hQշn�1�籣(b�hVi]+\�����q%6fp%��*��z��c��uK�0S��x�X�"4��Y��L����q�u��n��Z��B.�G�P�����-����K���z$<(��j�eAb���mZ:��( 1���YVO�X�.�&��:�~B��PYس�u��n�kj�E�=��;e��4<F醨6�d �WW��u��"�5(1}�*_�U�Q�zU�����X�����^�Ck�n������i���I�.�$'hʊ�%Q��C0}ð�4��SCG�맽|�!�'[�/�����^���ޒ��}�tS���=�뮫��v�����վ� �#�rB%P����S5Eر�]��3s���Kt��Uʵ�b5=�W�5�����?.j�7ٕ0�� {����^���U*4 �_�{:��	�h*4Kh�i9h]nzy��:�g�����WM���n�Oݛ�T�%#%c����}/�垽ʵw��&�m��~��<k�^տ���_+4��`R��V�*Zw�"F���tG�w������/�b��e��9Ji/=�v(\LG��w�ק��
�H4tKI(	�ݘ7¥%m�[�ӈh r�`�b]Ի���p�n����.����tf�O�M��z�e��ݶ��� <��ZQ�H`��#��_mɝ]Nس=�i:��|�^��~y�b���,M�TR!�Sj�IMo�I4��5Z��3=� >�[+��;�|y�����V�P�������~���c��;�{�wr�]4�Ƥ��o�\�0�	�E I����!���*��T��-�ڳ%��9Du��ֿ���#Wu�u�ӓ�*��:�J��2|�?(�:7��7�I������f�Ή�=�5�'V�ð�|@���<���fk�j�<}����.�@^/q���Zѳ���{�>�z� �����{�3�����f�]z�2�Yc�UX��b��V�\v���KlWf{<������b
r)Å�K�2T�nox�>'�ʻ2��>+!����!q�J���p���w[���9�D��_+֒��>�@4K�CM�]��4W: ��B�&[3�����ƌ���s`�����ʻ�k��Ň���,�ٜf >"�L�ou\��*
��${���h�6�B���=�pNC�)*������f�g�S�ъ��Kj��&�wf�z��)HwV^�FY�^���ڛ�Ȓ�T�P��v��VmK��5��n�]	�����pv�Z��&.�Z�oj���X��ݘ�l[ǝu�R���KGzV50�k=>�Ypoy#�S���!m�C(��sz��d��5�Jmx��}���
c��,����X�d��ʬ�z�i�ƅX�5<�f9+=�m:�9%�?sȞ�Z�\�FE-�Z����ʒ�bS� WE]��,�~��g&VW�wU���y'#$�	�`��k��Ƿ�=��%B��֝�LM�k4h<�M����;kH�,���ͱ���uک����Mĝe6�p���P?�[Z1�'���,��Gٺ���Q�����!�<07��8�b��:��l�)�L����S�Z�[yXM6��޾�E�|Z6�;%F��Y1qu�޷v<^��Y���pO��Y��9ڶ��^ _��2'�2tϔu��uѧ�M�]Fh���]��M���������������󕩪��vܭ�xY���1�9Wz|�pq���6�L!{��o��Ң��[643~�t��7wمUs~�͞J֪��-%5Ð[�%vV�N�Z}Z����� ���M�ё�˔��(h(�\v<�oh\>U+v<��չ``�����]oq��F�e�j��h�=#�T�J�jJ�|�#������Y3h��ure����a'|�cv�=-q�֗k�ᡊй?�h�`:	��~e�[��i�ϣ���7�,�uq�N�)r9)��v�C����!T�6~.�s��9!�D}V1Q��;�F��๚
��q���ga�����ؓ���^����:ȸ�����:�+�j�g�T�*�%^���� 8>/-�%�}-j��YK���|���F�z��ܴ�Ϸ0g�a��!�!��!�u���|�P�
F�t�DRE�גo�e�{��.�쫻�$E�Ҏ`��'ּ��ӕ�v��!�^7Q��*C|j�\�n`���?xx�J�@r�rm�h�>Sp||�4�tY��	*�Id�y�ۼ��q�D,�5������e�zM͢�2��Y~w"�����u�V�^���F��k߬	W(ӕ�:Ԅ��=ܳ;�#Ӡr{/��h�ϻ��Z�;yp� :[����|F�LY�39�y�a�Dp��uw�bo�.{�/*'J�Bޜ�~�C����7Y*�=�ܳ�3F�W�=�
�՛��N�w�;
�}L��Qˎ���#�OUf9��F
E��	-Hk���j��MA���#3�63���z��~�;:MJz�p6* e��hmZx�f\/{;N�+������]�b�:�>�cF��5h�8����6��}�U���������*uc�\�/1H̸�����m�n�]��n�M"؋5�C��u�{r�����.灭��}9��ے6�ݏ�+���a�ru��N�*f��`����6.8��=�ׇ$N�����:�ܛ�i�b��3�`ݺ��m�lA��1��%�cX��ݞ���!,�ư���z8�Tb�p�D�������:���i�ƹ'�V|�Ʌk�����cd�4����7k͗���yw8��ƕ�4�)��Oz)��Ξm�DF쥲���k��YL������΁FX��-�s�~��bf�f�8M��9Ǡ�K���=/��ㄨ���B!U�(H>W��)���0)��>4�P� �Aҟ@��K~��Ob�o��֨���B.)QoJ��k�y�jkd]=;ͧ��d�, �H�ݲv���"��q�-|�_f�xz�����vu2��\M��;�*�u�]4*e���i
4b�V �"~n�L����@�W��F�;:	[�u�u�t/,�v7��`�o���~��R8J�E���c;Ņ���ĩ{�ϲ9�}^�k���c����Q[k�����6J����j|4��R�N�i�ζ\߂˿_���Fn�����f]B�NT�
_\̱k՟>0h2բ������g��Ϳ#P>c\TA��x�nRn�<��{9��]�G9���#��|9����Ue�@nDY_��_��6f0��{�Ġ^R7�y��S+���I��]��Dg�Ͳ���]Ժ�8�/f�#�>������&�%k�C�2� w��Jn�-�.�/)�VC�mm�T�1�[WJ�c�C�*-b���#4˭{���b���gGg�k���]�qa9Ӯ�?����좲"�z�MF��W{��t�� ���e�(w���n�]kJ���U�4o�&Ӣ�_Le�,x^z���^�bc��VW��))3V��������C���~ʒ=ޡg,�76�h��UFWx�n�ټR�I��퇥�F�X���ŗ��^ţG���&�?�Qn��/��I�(��}���	+gY�4���I�j,��!Y�:�z��4�:�Kj��#m�ֵ���o�8"��C����;+δף{A���Y�-�-�p�N>{O8�����W��%�T���^L��ǩ�;r��,����\ �cAEmns��I^:=�.�ԕ�l�c�~�9rV�JJE����^oz����W���s3�b��\)
"���]�2�	�黦(�P�U�l�{�K��]��ohW hN��M�c�������K�K:�6�~��2SW��u��D"��|�z}u�O1X�'�E�Oz]���b��|��n�¼U2�S	:�(Ԧ6����6�y`����S�pʲh����
V��ʏG��s'-(XY�j��,lI|:���#5յ;Z��B�p��<��>*)�a��BH<�l��TinFq����-WO�.u��4ʼ�]�DJ��|q5iT�tNq�����1�HdwVxf7��NG���y���W�V������F��	l�rʬcYy\x|+�s*�g�y �w�ô�6�uh�WV,Ku��I�8vz�6���W��CLݶ��d*C+��^�Nj������ן4���9 �Pk��m3�Aѡ]�Wg����:%Ω�4ɷYW�q��C:���p�CY�(�"�����k����4.-ʑ�+%d:V�َ+-L�כ��rN�U]QA疵����0��;Y�м��d[ڬM�F�qMWSbP+݇�R���^Ӯ�ѐ3'.��X#�N��o�����eL���ZZѤ��=�2���*sK�������[X���(��4;X��7��.>®�8�����&f���c�M��:tpl����A�Ͳ+�x,���ϝhi�#�V#�f��o�|2�|���q�K&�Q�H���t�3R�vu�9����5����Fs܋W5�����j�Wn�;N7�\�j7y�8E�X��r1���{SA�xWCAuj�d���(�u�ǝ�%�� 0��NL��	W��7Ge-8�pn�`NQ��Z9vPɺQY�C�b7�R�a�PՎV�$�P��v��X4+���:��t�y�G�k��(fK��j:eM�����q��O.��UX���5�M�k1�E�lй��[�E�Y��~��ԢHIT�Uv�IVĳz]N�x��]Z��m�禳�e�v����%��W��?:!��h�8��eiTA��Q8w�X8;���>����c��*�$#@�X �V�
F�:P3�S٧>�J�*�r�{��˝J>�:Q�[Zo��5��^��q�+Ƥ5��K ��ym^զ�g�-�jO�U�r�*���㎶�u�G�i�aS7az�7a���8���т(m���?���A~���맞a{�|��muL�Y���a�$�8�Iĭ*�'(�����u̺׋¤���@=��lX��9����M!� HS��_�iA\��R��f���h�����}�7i'����QG.$�WJ�z��|�+�;��ʮ�u�B�e�h��#}{���R���*���E}7k�1Mz?��2�.�/3Ƥ���QN������Q��>�nn��z�5��qV�ib�=�O	*�R��T�"_h]��g.��"���=���o=2ǟN��-ת�Uֶ���ȬF�G!�J�J������+I',�|�����Ʃ
���oV���|2���1W݌!��&��p��'S��ĸ>㸙�7z(7���'��g�tk)�9qu�cV�����ń@t�&g=���B�"*���xq��^t�̻!V-x�:w}�[�Cu%�Z���{Z��[��r�����|��>��t�������;+�V���m5Y��|<�L'�E������0L��deL%C	m��g�-�Ҿ�U������2�p�*f(��R�J��EƔ+�s����)�)�&�1�����t�WK�b^�@P7iDH�C~O���H2'�_q�����w~�r[%��!rg���q�+K����R��YB�}��� �@ބ��{�?6j����P 
�N���e;�E��h�y�&`ȼ�q�e�G�MՏW_���u9�>PI�,�y�d��,��+��̗�x�y��
(����Asn-s$�]���A.�����@�v�ʺ(bb��Hy�x�K2��w�!U���.�UZ�{���@���:WSRי�ɚ�� �wi:�M-�������6���op*0k���).�+4�5�o�T�g�#Q^�5���ҡP_��Ȳ��3.]�s �˘�j291!�s
ʠ�R��A�aj�S�h�N��b���Z��tj<�][]��P;�η��B�jB4�뽭�%�%R*�Д��(:|'j����7%�cj�K�(!ٞ���/U��<��Onʻds��ڷ[K�ŵ�C��� ���8�WrEv��<�ݫ�D�*�2��8� �m��4��s�����	�{=��ۮ��<A�B��zx5$Y^ݶ��`�tcG\΃���s�x���Ԯss�	������1�V.:�H<�j,�����n:�)6���΀cQ;m"�mk���N�u�f�ݳ3Y�-۝.�\g�Z�Pnds�i�6m��4��^ᘣ� f��n��jM��w���b�\�vn��ރ}�.����Z0#Z�-4�F^�U��Ob�q��)�V�\�B�2�B�Zms�uV>2��Y+!���V�y�7�s�6׼M���2Z��/u)�@MT�	��o�S���h����H�̺F���g8��^���sqB��c%e�oe�GE���W[��Tf������o%��U:�a"^�b�R�z�O��6* �z��}9z�{�S���{�j�* ��Z��Mv���k�,�5և-:~}N�o=d+WSݏ�&s���j��d��O�S�P�Oҋ>;��I�����I����[������Y*�|rn�+��n|�r�.��>��z%e\��z
���5Һ��V��l��S��{�S�Y�%c�li� ��Q����N�����2�*��Z�ld��{FZ�,v�d��:Jnks�n:��0��q6��-�UPԌ����1���˦)R�i���q�r�w�roI�2�,��'�&��%Z�E�m���<��<�d�N�T�i���-J�}Ħ.����;ޯx�|Ri���^����B���EZ�]8�+Y�����2�\�{����"��@�j�J�gs/V�oz�zH?j9ݕ$c"��W-�J�������e�SS��mӺ�g�TwJ��h�@��t�@"��!��g]��fW�f_l�ġl���eꏻ+z< ��b�Sz��Q٪F��c��g	,�>���̰	�X��KV��ݳ,�w�Y����1gq˰W���=��P�s��2�1O1���ڽ����_����7}YewL��S͋Ա�v4�4U ���grIf��9|��_�d�'ݧH�0�?`�ў�
eg�1O{,�Fu��+_m-�Z19�/	�.�o���W}�yǎ��� ˤ��t�)'yvg���m������Ӯ	Չ,�(4I�\��4-�J�`�l�\~�X>j��`)��5����g���,��ә���K�j	�x{%_PTC��ҴN��˷bf��f�����v׽w
�;���o���}�vNy���^��(;�w�p�!�݃�vfa@��o8���A�i�=bn�7����ߐ�ۈt������(�a%R�}b�4W׸�ו
-m���^�ѹJ�{}���eW7S��3�]*�F=XI'1>U��G�3Q�p��Řos���۫�Y|V�����Ƶ7�Բ�����*>d�Vx王cg���6��ŬF;�(�%�? -2@, E����쨈�Zp��s�e��ƙ�b"����Xj��w�f��W'���\��c�9����$W���Ûs#�k�����YGu�j)����z�|n�6	�Y((��Z�k�zs�[�z�x�O�_Yy�`oTO��K��Q��+�=|�a���T� ɦ:۱��\�������Gn��9�n��{g͡��Ҽ�!KB������Em1�����qʏ�ީWN�:�T���m�ā�Q�oN��R7�Y�uʘ7�Oq���x�͊+9y���#GGaX�DJ�I��n���9'�g�vm�n��2F�
B��zt�'.��pޕkWyYh��}z��U�VV_��ql
r���B%|X!�m13r瀺�l��r�˰�U��4K_{`�XjE[a�١�>���x���;�y�;Z�)HhBp�9��E�*��y�^ѩ�+jT���s�7�ͪ۝�)�0�{doav��SdS9��P��(?��*���:��O����Z� ��"�vK)�r���+��Д⾓z�C��wzl��.�!���k��(n����6���j\=7v�bv�4�>�=~N� x\l�)�*?DH*FˬN�Bً4'0.V՚�w�rM��Oz��w��+����S��x̂��i��bBe���S�	|�uG��aݦ{p��y���h��m۫��w٧��մX��>k���^z,gN��߽�뫌f�o�����V����`c>w�c<�m1ЍU�6�����@��~�m��l��K��g�ϷU��q�9)��K�I��]�s��EVn
{���Ѣ������O$rosVt��$�X4�5*�݋��I
�7���������KT�
J�bl�ͻO�Fܫ�9���5X�F�Fom-�B䃍_�?W_w��.�ĳvkG4��lUl���g�I��e����(�U�J����`U�LK�wOr)��S�R%��'NW|\2�ώo����;�i��͹c%c(/$�׏�{��%�6o�!�_�r٫��\���B�Hږյ�Gj�ų�����M:A�����S��B�Ӯ��WL,eX��Gr��}Vy�zI>��J��O|�~�k�P0�=w�p�uԦ�6%�'���(+V]h�2�o.���3Ve�"�|�0Z��Gd�$�av������&�eM�u���H�:;��mD�i�;�K�5��Cf��m�ok���5�<O�غ�<�Q�ӽ�@�/�ZgT��'V���ɐ��`��KFN��Ϟ�ne���(q�8r��ݓXvٳ��t��up�ټ;�V=tG\�AͲ ]��X��#��٨�N8��l��n�
��׋Nm�9�L��ݐۖ��:��j^�ٸn�n��d�ۤ���s�m�3-�`뎎y۸�G��Y��i�v�@�=�����w)��nӘC@��f�8�ݧ�04] �]�y�!c�|��I1��6�N��Ė�8��AOJ�4�Yc�_.{�����~���oE
eמnX��Ϟh|M�,h���,U��;p�|���TY{7Ԇ�L�M��� {�e ���n�N�{Ӱ���O��sܗy�d�:���gI�xz1����hӤ� �4�l��[#��鏹��U �Z��^�ʽz�Ǻ�+�7C5��$�2�����V�Y�3��g��c���4�_�V�h'I��ŵJn��;������1Qvi�[��G�l�R����2�l�iUs�L&a��|	u�E� ��T�����=U<����X)�,�Z�l�ī=��f{�����nA(���S6jzɱ���Oq��nEI#�iMg�������,���V��@�� �߹<�#����X��x�2��9�ۗ�����:x�HM=JluV�Q
�%��E�ث����E�M:4�U��nIZ�/*�Ok��Y��@8�v��˦w���ޥ[k�S|����*�E��j��Tj*�eТ��i(t=�}�,���|����K%�mW���Ԁ��{�3�҆�u,�f19�����<��9�]N]v�r��ө�qm�~�/ǚs�[�vaC@!���Ƌ�s�>T=[<*{]?ct��uv�G�hP)��t�i7WXG��y��6��t����Y�i��Nm��9�?���y@�����{U�py�v���*|�H�Ӗ�-�_q�6]9m�]`�E2.�9iU��HD"�.v_�M#J�6�{��d���gC���}#��O��J��j����䳛\PٱS}�Ojh� ���6n�r��/:̮B���)P6��yj���o�-���򷷁D�%o�}���[��5e�mŬ'\�l;A�@��Yݺ�r2\�v�q�o�k��䥒F����H�Z�뫪���$��W�M8>DU�ם�6*	C�P�)or��iqDcՀ�����������g'I?zzx�RD P(�g�i}��Em�a�O�Bt�`�,�X}��g��|d�u���ӵQ�-Z񵰊�o^�g�:��j���d����k��KdVƘ�-�KI�A9=[|�������(2���G�R�q���]8�VPWi�[F �M�&ꕀ|{鈩l���&i�Q��w�	�5ʘ�Wjg8��Kk)�=iwͥOg`��O�om�� cޞ�u�ع�'��0�q��K�!P�[\c4[? DS-2Eˣ�?{�v�����D>g�)����޷]���+6�Y>�<��~)N��oe��i�esc���w�·�hi]L�x#*�E���[���/z����,����r�����z�@�knY�3�T֗��y^��[��"+2�2o�|OE�yݟ=az��H6��^9%��ʶ{�Ëٺ; �ݚkN�/m�M[�NXq���� �x���^���v`�f\��}8�����W��9[����2ر���v��a~s��a�<2� �.�-5r�y�e �t��*［����N�=�&��װ2k���M�s7�o�f�)��U�(Z�ކX)�i�
�0�fOIb�lE�e��m"�)��VH��vCp'��+�^��f� _d�gs�.�|ӂP丹�H��v�]�7ַ��
sV�gG�mX�%vG�)�8��G����&U�^=��o	����DY�r��%C���mط��R��(I�N(fj�2�x�yr�x$� ìh�q�ͼ����u�2�*�܀����$��1]�+���L�zf��-u�/
]}R�o9����N�Z�MI��7@%I4�����u=N��o�qQ���m�4k0\�V�,��{�#<�eo�<%��1�;{>���[����2����ʠ��X���=�-O<c�c�.�� � �N,�64:f$���4����=�h������2�g�*C�9������ulr�[���X�\+ǽ�ى-�W��k�ȷ���#�LNR��ֹ����侴̦o|y�����k0��׆�����2x�y��imd�������p���}6�g�gtu����>��4[%�)&��v<Qq4�����+�&�6��~e�I��E�:=���m��7�Z%
��B��-_����XИ��GٴއCJHY*�$���Z�6���s�r��ϝ=4������<<�g,�T�I�;��Ϻ�.���N�6#\��^~���G}�+�l��S્��h�Z@��}Fx��5�!s��He_�RF�ؽ���,��=�U
43�Vc
��H`���߀�\m"��qy�8�*��>w	=a(1ؓ�f�F�����\a�C_�V!�y�_b��ĹG�E��(���wN=>��s����{����"
X��d�
"쎇�ӗY|��&�������B�a9%������ū�w�	�p�D0�U�(�1Ӡ���S3R5�w59�z�QJ\��X�T4[��x�F;�v'�]�����Z�A$,aѥ���'n�]�\���������Z�>�NNL����i��nn��է�fvͶBVZy���&P�q3�ܫ�帒���U,�D�I>&ZPe���2s�#/���[�MXѽ��S���&+���.��
e��I�o&�R��F��4eN�:f�Iuy�Ч'ƙ�2��{�_�yz�-VGy}
u42�u,쮰3:��+��n�Z(��T��ՙ!g�D�S���ә�<Gw2���nRb*[·]o8��a�9����b0]Zk[����E��E�W�!���V�����<�-`�|"19[����3�t��>ԕ^��Wlٽ���4��)��������	ţ�%�%�]��ٓ�i6�B;����Z3n�u�2�QvT�����[r�B���r��U{ qF"�̼�z���c+N��;�T�_!\~������]GY���s;��2n���=R�D�[���т�FJw�{����>Rm�/rY�jW�br��L��<�$Z��{D�&����;w��hD%N&$�yΕ��v�`�[(��m�Z�u[�Z�ކF*�w����1���q��Sc�n	r n��a$�la:Nxu����G�ǋ^��7j��:3{��d�$���ͭ��Wc��m;��K�%\�a�s`�f����(x������r�iw`��Zr���q��>2]/k��.��`͑�6��2.t:I�Nޔ�<vn�鋷'��k\�5�r����-ݍ�V�nǮ�n,�\8��szn�qvwl����Yg�U����h�۷A۲s�rnɦs�n�=b1�y��qR�.wgW��P�#ܻ۴��g��k�٣�9��7�������t�vG+�봛R=9���{�qɻ�r�>Ɣ���ι��.'\Cuq��n��q��"�vz�<O�L�'\�kt��'{��8]e����Y�_n�m=q��s�ەᔝ�g7h���i=a��vjy���<�p�.�m�<�dsBr
�P\u���ϧ����\��u���vdC8�� 6_k��N,���%�
ӗ��i�m#�YM��sQ�s����8���Ս<�ōSU�웵�t�շY�prY�|�-6�&< ��̶������[[X㋇rZ�,�=׳�m��CC��X1���Y����}�_t����Ӽ����.L��ۍv[��l槸�m�Q�g��nH��v��;�]��҇g�k��,�.�g�6�v���x^��[����v��ۏg]����z�N�t��K�aJ�s������녈���(;�w�6�M�����p+�;�I�1p��-�HMu��:v�V�8�ȼ��랓�h�x##�X�n�:�I��s�g��lc�k����oZ�7�y��Y��۵�F��7Gn^N-"t)��i��.��s��B˧�x+����);4u�S�Wta��w.Ɓ���.��0�7Y��	�М��t]��=�c��۬�X��h�m��v.U{^'��s]=�nzѷs��1ֹ26�c��:�#��t�k<�GF��:�-��`��ۥ�7��-��!�Z��%���v�n6�0a�C#�c�|�E���X0�מɒ3�v�vG�]�iM��rT���

�����rE����]�v�;�=m�V�[�{�jrpuٸ��lwg-��f ��$��z�[xִ�۳vI[����s@������������N�㡇�sh�ùM�Ѭ�q<[mݓ^�Mڳ�l d�wi->z���N�^�Q��Ut�K[��v�=F͍�k���L�vM�o��sO�=t��z���.�Hm�Y�����5��m��;�۠��v,:�n_����Z�i�?C��܈��[ܭyh_:��[�~�6c�s�їX��f9㺻�v�]&\sk��U{�Ch�gN{��gUq����	�5�*�-�d�s0(�f?����rF���,e�Oy%��w�Z�Ę҅[����;|�?x�2ݰ������t�Xv��Ԥ�*S�Ɖ$�"ZA7V���F��~;�Ko:.�2�l�;�,�R�o%��_��������(���$���\��h* K���ʥHIi�#U����ndͩ]-�tr������l�7ۦ1����cl7ޛX�-(uo�w�2b}շ=�U��u����G��5ji����]L
 ��{}��6$C�M���u�\��yl6��=8��ui�读Ӕ{,�T�װq�y��}*�M���l��lq[G�KK��o->�rW8y�m�/�Z�]�ѳ�Qs�o�),�o2�����xB$�|���1Lq :>�sx+�6ў��{�]��YFY����{�:5�F�X[	�l0)Tw�A�l�}��'�Fbע�ەuvWZ2�)d�jN�z���}�D;�v��y�Wڒ�$�/�M���5�ݳ'.&��3Tǚ���ڐQǻB�T:,=i����٨)Q���y�d�4۹[��r�7�1-~t��5�ӿa�������t��T"�l��n���,C����+�ϓ�%>\�8;���כ��w*����.����z�v�y�g V�<���5�e2�h��4�7�˔S8�@�ޫ��[Z+β�q�,�V��O�M�ԴFSo�;]�K˨c`�h����'TY���^�\�i���o�&ED�J�Łr�Lx�K��ԩ{�g6���*�ٙ�Hs/���� �ߠ������_jl��᝵`f1Ƀ|(IE�4.��Zd^�Ͷ�Es�e�QQ1�:���Y+1����O!D�WH"�ZZ�y���\Ǐ�{���Hs��5lW�;�A�DD����f��v���=�0�{�X�Bݍ{ N��N3Jl��'B��%���,��s����Cxӳ��~�ȑ*6vM7���c<WY�Ҳ'}ŶR�m�6��o���d��n�����T�wmv�%�
즶i�L����v]�]ʕ��oNԡ�Q�~`u�w&_
1ep՛�u��"C-;����j�bo"�)�H�M�]`-Ʒ~�{�&62� �<3��:��o�7ڤ�U��Y'��݋6���.����u�^bN����������7�	�y��;J�z>��T��gn3.1�����=��d?;~̜w�+M.o(Od��E�n����J.�TX����
F�+	*����n�X���o&�m/��U�
7嶖�a'��ں0��"�����
5��M�>�_�f־"炭\���\$�s�^��W��r7l�zۣtV���
�q�G�*p�E����'9or�k�,l�z����5F��m��򷣥�nZ�و�gr��V���zf��d��Y;,֐��=*��oX`���K(�H� �yg���ɉ��j�����ț4�-0:_���`y=[�L�7FQQ@���!ۡB��4�M0;칒T��ԧ�������d��֌�s^�'���ߙ�s�ޢ]�C��:��/{����[��'�,D-L��U���1�c ��p}5�˿-I���s���Vj����&l4���l�Sڽ��U�hվ��+�8��֭���Y�I<�<�b�UBԾ��(�o���$�}/��"�_4"����j#��p��|t[\oq��k.k�{Ѓ�ޘ�^�`���E��"���\�0X=��甯�Y��1z}���]Ї�M���N���2�Ƃ�C�y����b:H�2W�����3�j:�b��q��e@��H#��D��'E�lh�<�m���+9���9�mf2�5��:�z
AJB�-���E�Ū���~&��j��VW?*ܚ�e4M.��*�=����^��dɳ��.%hc������!���(�̫%Ԛ]�2�a�}�:�q�+�V׺�_{r��l�t��y�JЦ��p0�=�įw�ҝ���~X{�p�J���P���	6���8ګorOQ�nহ�����r��~E�ґ�=�����X�t�uƎ]U�~�mv��HQ�Y�N�oĤU����
I$�h3֕�5��_73���s�qۄ�-x�	��c>�^�%u�[�z[r�z�m����5�f�G�*��fx�=rmڨ�VB��ɍh
�>I];�o���Yl�eԔ�;��ukǪ^oV^�f 	Y����OL��z���m�߭�N��L��]N\�j��� �Q4O��9,C�^�O�������,�T�w6}[����9bu�[�uj���zQ=aQcOaw�V(�ݣ-9m�;<]�E��3I�a$J��}�!��=s��WAs��꩝���l���!�GD�Y��<�6x��Ѷ�nK�3��j�ՍVk�.�b)ǐ��G��;�j��M�t�h-���xѓ$��X<n��@/Zr��c�@ꔸ�͸Dd���2dͼre�ٷn�sv�M��<j��zy�v�ۇ�=��:��g<m�c��>��9�b�n�H.y�[�5�ϓ�[�8LTWF�����]�6�Js�R:�qԚ�<�8��./?lƮ:�),V�!UH�?-���f~��V������1���^�C'�y�����r�+��q>�h�r�W�]��T���"��g������"�$���VdgƃG�Clp�*���靴�OFax��8,�b�W����$ZK��s��9Zr�%Rz^^{�x
��4�l�I��aNE��ݜ��wV���D��}<�JՓg}��5��)���N]5~O<H�XH]�M����k��l�ͦ{2�~j����u~����حK ;�dn���
%�x��&�9��ꧧ��׾d:Դ�3�Y\������[:�-|[��"�s�*A����Fu�~�V,�%wE�OUp�Tב�qN�Ǉ�Vy��.�^�]��.T���%n�8'�AO;a�~��S�2V��񺺲s;���+[01\��]u�e۱��IF��L�eX�*�n�v���߼���q�������]��*��.�+�7����aK튙�ũJ���^x�EMۮ� :)��t)&[9�Է�}�`���}���y�t����"��n�ݼa&�
3e�:����� E9|˶�挵&��lX���d�	3��ШqXg��\Ev��M>����ʱ$`L��u�������̽%��*��Гg����G��v���	ss&�KWw�9z����o����Miw����QlP)(�v͛�_k���(
�tu־2��*�;�:�ܭA�ז�7N����Cn9�J�{>�s����W�V:ZR��3���`����Ӽͻ��:�\��^��A��]潷Jq�����N�{''������}��l���]��,4�I����"n�O��� �o��╖����Y�1��Z��B5=Q���ؕ%3�Z�LR^��G�ɳ9o�8y_"z��y���UQ>�5cCq[:�t���zc�{;t��۱�Bxx1v�uyː��0�hRI�\B;̥�/��������H:�%��7k��9%N�c����"���>d�vx`p��zws����d�P%i����.�Y���Z�ڇ�(3�O�e�خ�m�,�=>{	<iY/׳�d�^0!s�*-��+�k��mf��+�#�J�ɣ'�f����%f��7��!+�K1sSO��~{m	W�ͩ��u'�C&��,���λ�Rͮ�ǲ�S��0����{ٲ�:jZTHI��Wr�2G6Έ4�+闭���h��J�%��uU�%��"v�e"�ԝ�S��i3Ys�x�Ǫ2 ԝ���˙�J\|��x�'��W3�.���hs�L\>ù4		0�MQA��(��M�A�*�.A���X⸄�����Pz����&�G����9M���q��(�;V�F���Ԝ��9���*�ݸ3��%�:��=�2�����O+&��������L��Z6��k(���{y=�q�g��xɤ�߶�~����ޥ&���/)p,�t�^/T$m�O�OK�Ӻt�zU�ܑ�
�ʪ	AZ�:��8*T�7�R�_%ƽޙ�^JX���l�Lϖ^�V�a�VӺٜ�������[�>����myR!4��i�;�~j�Tr9��*_3,x�^ô�ɚ=ޥ�źj�kn��,�[�$����oۼ�Q��zs���]X�E��I���=<T���w/�M3{��ۧ�Pl�6k��h+�������1R�x�=�ze�u*�r�8�n�$�=B��3껌T��Q[4T����	�+KN�}[���η�u�PZ���Yi]�7�Ci��7]�r��.�g�N� r@��E���l�0c�]��eY���1�Լ{+��g���V!��xී;���W<�?x���S"/y�"��n
댐;0�$ӤMV\m��q\�6�0�iya8;;�%���k�d��>���;\��h��3��u���({���M*�j�=�������^ty��]��i��-h��mԧ����>4[H�VYW9�s*���{�M���s����,y�/�=�����id���4�*Dkg���}�:����r�h'�+��	h�Yd"vY^��R���L��*`"�M�=|��D9u}X�В\�r����������Y�{��������EĽ@p�>!INn8�hxr{Ht����w��b��(��:�\�(��A��\?c���e�A�UD�V{k��ɾ��D�b�a�W^$"�	��׈����+�}R��sr����<��y�G_����%����ڭ�Y�wR��MЄ���M���W�3��콗Q.x�Z{�5 �_u̡�>�{R;HG�$����#9��<�^ށ�ioL�K�c9v���m.�ɕtrH�~�V��bMwBѤ��a�6]����F���.�٫�n9q�x�n�Et��U�#�q���xl:�y����q�����8=Mùz�0u���t�؎:�){r�n�&��nM+ʦ���m�O6�-���5�C�۴��R��Kqצ¯	���S���4�L��9[���=v�lΝ��\Y�D ��{LpgIʵ��1/b�qض��"��^�v�9��E�3�����OG	�uqD�:e�����w�+�o���c8��A�{�����٩�����}��p��-rkҍA'fmhC�.�!WdR�HX�QQ�V�ޓeL��[ٞ�z�5��=�^����^���b�[}���D��?j�6r��~=�Y��幕�"�4�ۄ5��tj��(�c2�
�6٬d�����0��*M�VW{ګ����]������D쇧jS�qʾ��M�]T�Ӝe.�R &�
E$��/���u=���i�B��.��U����/Y<�L0G8���U|�XJ����uj���6�
�{��4�����0�M��e:ۺF�)#C��zζ��C�?pƍ���O�S�	8H�ߔ=ݔ��9*W7�~�9]]��O�r&�'hB)���M.פ���m&�9����{��V���[�TA���M��?y�ё����2�ZX>�l����>��^�ܽ7l�M7#��՟]�M�m�A�̺��I%�_�u���C-Z�C�N�z���3��;���b��&v�5��7�j]��]ve���$S�s�=E�B��bXr�{�j�2��+r�7%��)A�z�6�"O3���A�����7^��V���e
D��#��u%��F(��3��t�&�6�ץf�n����;�Q{�������Ԙ0����3g=5ʩ����d�쫝uCo��3.^zj": Q��9z�V���މ�6�0���w���{�~}��&߉����b�燦��$�mM�u���;0z�:6	��P)�PI���*}Z��3ՙ쫭�{4�ME~����읬��E�Yj����/��ꉨ��zr��6*e��yi�8�c�ROjA�mWF*����	��9�sWcs�L��9�����mN�������
u���U�r�w��f�|�p���fj��T�W:挑>KQY�y:!޻�M���{[;���Ys���Sg6��p�Zd���z�ۯl�zL�Y��7��tR�r�켥^�K��@^=��ܫ��G�L���S�w�_;h1�_j��Z�*����	��$������;�{��*��t���;���<C��[յ�$a�x4�PҚ���t����6�iƤ�-�qͺ�p�@vc���"; ��M�j/?n��]u�^��o�O��)i��������q�@��]wsijwr!E�*pԤ���ȹ�W�8�Е'-w!���;�2��"�j��ӡ�yŅ]�����K�js���<�Q{���e�tim�O��,<�횂&�d����n���>Y�t��!������u)�k}��f�٨�����l.�W�	\�޾-Hu.Ӌ�ۭ�������ۜ]�����}��0��/x��/N��%����8���ھ3)�K�F�q�*�;�T��|w�p�Β����Sw�9�+��'+x|}
?�6��U�Zr|���ɜs�醱��Xq�W7T�0��1���@ܕ��-yK-��Q��X�[�6�T�ْժGF��}v�s��]����W�Gp|���%��[��|SJ�5)�or�}�3o���&���d��u�Xh�j���(}�?���kX�q��0v|p�:8'���:]Y��q�C:��U3I�dMN���U2�Q�w�o������5��9�Z����C��ү��匼H_�J�*5�;b�9Q��*\�_F��:����0r��$}�}���q�wEq�aM2�y�T��K�B�ӏM��\��2�
O��ܬk���;���]�Vm�Ǥn=���k={ʸp���Zz���b�.��um�7��a.���tՃ_N4�8ڂ�_���}$�*������W7 5�XU�x_?���y�;��/س��u	�;�� �Wϩ�m�X�"u;l���\��^;�C�{]%����p��#�!��Gws��u�TZ� 	�v��;,H��ڐ����^w�r�ӦE� �ffݗŖeGe��B&���=�㼞mN����]G�
R������ƞ�����BإSQ���I�x��0�@�v?|��mc�q�:�S������ئ��w���[�����S-s�I�Q�q�I�ww����V}��-v���z a�`�8펕��&	ޗludQy̽�5B�R�D� �-��1��M�v<y�k� |�b�?zD�W�h����ѤԵ.p7��F�o7Ya�/��n�gy܏�A<�W,�rJi1�x�w=�ո�?t�|�ޛ��#]�[��_���ץk��J���i�C�Z�}��V�ar�P\S3^��5�|�Q�Ib݉�;�r����!�W��a��yْZse193�I�.�֑��m�*;��K��޼�2�����'5*���=�Or5ľ�uӅ_�vA�{�bl�t�Z�k�o;�@Z ��*(�IHG]G���~ʒV��"p��X����9��9����k��0O%Q����fQ����ѹ��Q���f�/=E�ӑ�i��n1��vN�97XqyP����g��^�9(�����u�x�W��oJ�*��*�<{��ɂ"�)�gڃ~�כt��m�DR�n���F���z�?`waj�Ŵٻ��Pؾ󥽷ꞙX����n�ڿO����������*�L�3�,^�Pi������"��Wy�G�@�H
o�n� �	y�w?x�Ϩ�tf��/K��Jv
��
�7b�����4�V��%<X��+q��wr�����h��Ѥ+[�)9�i�oPDq�'�v�}���flrv�R��M���_�rc|��f����Oo��^ɺ	"�H���ԝ�Q�VW$d�J�Vkk�M,��=�bZ�/9��@& ��,��WQ�.;���)�[�Qf����:�}��^K�I�Nܥ���I�	���"[:�s3\Yyw:j�*�]��)ć��@=�ho��+S�l�Dλ�t�Do�[9���se�PN�4/�&���'��"8d�J@�BZ�u��=�S��� ����$�ќ�'lnK��şf����<uԏEnxv������_8��0�c��!8D�'9��u�n��q�;`s�M��N7/wc��&��>Yad�cj�ް/Mͺ.�I���\��s��ۣ�n��dcqR�5�z^x��۷mű�O\ny�m��Xڄ(^*3�ѭ��a4�.7��F�9�-�v����{s�}R��+���N��y��u�ڪ������V_�������N����9�f�O8�5kv������=�O/%��N��Ҽig��R����N����A�-�`�Cs7.)S`�K'-N��:=k����;�\��<�k6�����T�1��;񞄗]q�W ��/��_��$S#+�Ξ쾵�Mx�D]&��9��@�h�>���u��:3���,�n/YZВ7^����Gh�I�!�[�H��b�׺�:n�c;�FE���65��,����]�-ǿ53��þ��s�0'��oU�{�g�Ԉ6�L�V�^ڪ(����嶽l�Ս^9��sJ�h��B�I���p��c�A��o̵���L�g��.Ȱ}f�VɡOV�����"�ƋH�qH(Պ��L��f��67��5qu7]��܃�K�AK�,"�	�^�V�oO���y/	�ދ>����vpU���K����d\{v�;ۇ�ȆR���b�E4!4["X�<�l���\��UehD�	�w�y�yFHf,ܻ`��Y�/����u�F���鴠�w[��hݖ��N�{"�;���ç��XӦuW�4�ݣ�9��<�P=�M��Ϗ�w��;����crax��JjD����SX�5����&䤕�t��|��9�{�e�ܣJ�ߚ3�����D���U�-���o�ef�����k�]e9M�{�:���2�H��9,�ֹg�]�wD�i��OL>��R��d�AX5���Z�u��G���Wv��%e5�So�洲�qb~�
�8�m3�?s��v�.�����rp���&�l�t��8��d���Ø��cɴ�<7Dr�����lenX�J��"�Z4����n�A�>y
�=
��Mժ�b�u-��5����i1kz� U?����Tߗ;�d݁m��!�ݮ��^�]�sV����樚K̙�&�����Z�����@ke?�khݶ�׫�j�� +I �Vr��޴���i��%MȆu�Cs�t2'�fb����v��9x�׊Ƿ���t�MOw���޷�~��j��`��^R[P��ץ�8���#���MxƇ����Y�����R�+�uz�� �I=Z��3)�q9癙i��]���q�,P �_:#�d���]v��0N��&.P��(Ga<P�����m?
vbw[�Oj�-�(x��ׄ}$Sq�U�g��+5�E��Bk{����n��s����ӹ5��)��V��g�J�^��~X|��8�oY�������c�:�{O�7E"�"£jʻU�����p-P�^��-������x�����jD��z��T]քѓ��������A�eoW9�o�$p�C�I#QJ�n��%�JNV�,�4t�0��
/��e���5o�S�����.糗��o1�g�Ȱ�N��o�r({��i��S������\�b�1�����8���Gl��J�2��D����Y�oK�7��h��홾���xQ���OcSB��5"@��Np�AP���~˺�=`Rd*HѣIYE�"[`7x;�´�J�H�r����I<�ٖ�7;.��\FG�c�yy�kY~�>�rM��D#(Q��܊ ���N�iPM���U��U~�vK�{��ruv�
K-��o-�:��ś�r�!ճ:K��˛�����E�.d�QX���x}�����X�nѝ����;y�hX�ld62�.������n4��zs4�wU�;Sy��}��7|E�Tܩ�BQ�|O{2�x�[����^�k���Nj�A"�>�6ɗ�ϑ�R��i�Z��כ�x��.���g8Kc 4����S�������q[���F&&ʠ�R�!�q��v��gj{y��q�Ly.Î�pt�x�7��fX4m���w���.qX"ڞ��$���H�hoNgm�=�~g̻��f��v�C2�L4}�Q����+�&�5�vdΆݏ[��f2vU���*[�[{/�`��sen�9��+�^P%����"^��%�*�y�C���6RJqq1�{�y�=���һ��kh���Χq�[w�r��o��Q�t�'9�,w�����G���O��t>E��Evj�ɏ���$�ΰ>��a�����#�{L@�0����fQ�n�d�i���I�N[��ڼ�J"�����9�I�AeRn�ۣ�
-�E);�;|3�����9�{��Z�h>m��p�&����F�0=WH���*�m��<���w°>_�ݶ��RJ��?#X�r�X-��;��ѭڽn���-I,
�.�J�)�1̒u��M��K�oGȄÊ�H�`��B´-*�E"A�n�srb<Fz�ݸNָ���N콞{Xz����oY���þ�6qw����vS�pAm�5ٌ�'�;[jsv��錗m������K�	�>��e��OjG۪�s�k�ʝ>�p�=95ۻ6v��4u�n�8��Ip�N���	��mv��%��z�����)��_0�5s'E��g{x뱜���3ӛ\�s����*�B�^�{n��]-ݵO��كq�f;j79��P��2�۳v����G��Ŀߞ��&~9u���Qp�������.�[B�~�5���k�s+Ƽn`;-��y�'w���Y64Ѥ�9�^`ۮ��άF�S<h���ZEi��n�f���{B��i�O	§�\ n�V��z�l���v�k^�8��7����!E�R)��o~򹼫z�N��
4�g��mf߸�P�<�Y[�`������6LRE/9[Зr����M�$��]ի)Z@�g���8�sNiy}o���i/6���k(mD�x�)�s����e3O4���($#*�3�6j���Y�5	�B�>�W��Լz����1��',׷�©�AW��wծ�s�mI|��t/�ٮ��/ך8��|�T��U���웛��ٳhPT�=C��n��v��h��u���&bB���f�ƁYP��T+RZ/g�ɫ[M���y�u��\Bi��f盩�=�v�b[!��N-��a����{gVg�z���������!}v�R�	*�2$:��E�E�w��}Z(c�)l6^�R'/ś�n=�M������uἂ<9|����uN��*f�sU��m]JzxTLS��r�(@;9��V�V���U��I���7Ee�3�?�����7��?vC�1�v��k��oT�����{�:��7�mq���z�*n���`
���3)�iz׃���b{nɼ��l��˒̛��y���ܷ���@��%G�޼�l�οzY�6��
Ha�"� �p�{�D�>q��J��k�{8���N�;�<�W�E`������?7W������re{�<UavF蔃��S7��e?8��m0�qh�o]Zߝ�B��o�r�@l�_;��P��7;yｯ�m�dnmǙ�3�]�tkQL��?�O^��lY��M�l����9�՝kXK�瞹*�L��j�������U>��J��w~V���{+��Ey6��ԵV��
������=�e����|4�lS��R�n��"�(u��j1�1m��#to�:�{,���t��q잸�_È4wb��|`ZغW�<��-�|��=\=z/y���{��IT�0!9�y]o�5bn�{�(֕-N��|�1o���7�i����*�m0�o���V��Ȃ��:X�{kgwC���=�i�ǝN��J��p��z\ۻg��9/L��l���a���)�S��p�H�����Q$z��K�w�4h
�]�R����N�,�tu��)b�-��s�b�a�)r\oNF���i��}���LN�@5�yZW��2\�\2wL 0�E��)��~�� �O��:k�;m=���8iüٵ ��[��4߉̥�pٞ��k���zs�6.���nPh�N���p�[ho��!=�������۶�]vLXpl���M������2ٝ�w�Ͻ�{���Ê�wA[�߮Ю2�mzꗵ�W՜�r�4�E�6���V{���:`�аQM�D3�+��*�C9�x�m�K��K���
�:O
�������њ���ݭ�ț��=.��oAw�;⩭�6i牰�Yi��te�lfJ�g��viR��ă�޼�t����{�Ќ�M�X�����}0^��j�5��ؚ��zl0@H�'�A�I��컔������m�9�FYH���|
�w��nE�.a9˭z*	�[!�$7��y����\�`v&����]�q>X�*��ήQ۾�p�[o8���jsufN<���[�E<l*�8;���߷�N���ߨK��	$]:��a�"j��ƻ�m���J8}��	���e�k�FvH˿�O���[�p����!ޤ���G�~���V*���c��C��#��Om�S2c�dl�n����9ܭ�4P�N
�+uՊj���&O�+u3�m�`�����ʳ�ס�w*j��X�s;�Ÿ%:V�jU;�����kڊ)��i��-�t貛7�V�&��=�G�SV��^9{C����L������b�nʮ��ƷϽ)�9�Z+އDr�M
n�׾���/;G�J�$٣i�?Y+��g��3e�;��Ôn{@sޯf��Z��{�y���2�0���/�SD��I���!�`�HM�.�E7�Of�^Vwu��g=X���)���w#��[Ԝ�nn�;(ʕ Sh�j�pf�w�[[���r�lzi�2�����k��� �vyH���+5���w����]^�F�]�v��|w��>n&x%�q�U��'�}�%M�2	u��FxBՕ$��:ո(��ޮ�F�7��_.KL�Osh�)���PyE��t]g`4��o�.��B:٫	6\%؏�X��J�x%mp؂*E�Ֆ���{0�w�S]�������Ջ�%6��ɧ6�!AdsIVc�����n�v�,)�-�5���w���	+����se�j�m�|Al�u�4Ep=c(N�@��p�0n>�gEj?&�،��fT؈Ә"eD�{�j��˓�v��v�x�%5Ѧq<Ϧr+Q�i��@ ׎P���{�{i2��1���p���@R���*]ps��tm��r̲�Y���9uM��qj���ut��q��P����w4�s�\��$�7w�"ِ��xh��X��]ۂ���|�u���)V�[�6o�bw�w�]���Zq=o��ꉢ+�������b���*�PT8�uݔ�Sۧ�'-g�Q>N��&e��E��X��g�T�ao�\\�r�J;��l�ݼƯ�Ϻ�H�u����Y��]�����P�ݱ�'��7k���b����K���'�G>�/+�]�j�D�eD�tSQүl�F�ܤVn�
���45Y�&�M��0�͝��u�Z�o7��5U����=5�sl"�u}wF.W&Tޭ׊Y��WA�d��i1].�pG�7S���˝7���g2��}���띃E�L�
p��[�P�-�J�r;{��D��'�^�k���z���:&1~ꆷ���|��P�׼�U�HoN��C /m��1���W!�@�*�ĝ�t���_A�Wzh�ݦc���[k>���B�+=����Ƀ'��<T]��y�)7V��I]���K-�����أv5�l����`�ū3���2��Ktz7Z5�a���Gg�Ƨqه��<�Dj4�8jq�0]fR���n�B�%�`%b�nZ�[1�;v�^^+�7u�<�]pW��p�؂ۋl^_GAc�"����]g�÷��o�Z@9�\s�����m+�b�*n=������7��幌���ݲ�T8�X{=�k��.<n�i㇘灞;���j'�St������O�[�qɹ�-5s���5�
J�W�7C�'��bj�cl���]��x{L�j�Y8緗g��׳�k_?G�������i��Wr���g\nڶ��O2���Ж��0q��;��>J�x����'�z���t5a�������;�U���m��[J"������n �Y_�#��uݽ�$���.ڸ^�M��<�i:�q�)��K3�\�x�Nv�m��p�:.�͸q��%�]��ueV&�(��B8�C�j[�WmۊC�����y���;����#kՓ]b۝�	*qm�S�����Q�=O;]�u%��v�v����c%���n�Ӗ.^���y-u�v-���C��s�j�8q�\d�}F���cX������\�:^v�poO4�e��m���\�r��烵�������n-��l�+N�^�u�yԺ��M��v^ȫul�q�uxySny�.����S<un7Cʇ[��n=�jޛ�]����Υ���[�p��Nz�v���Z.N:������؇cV�/��Y���u�cu\y�m2�]�[�<�=g�����7�8�f�M�87<�v�{t��1��h��&�m�Az;8v���H�q�vs��=tՌ`�����/5�'�譡�7e:�퇞V�X�z]�&<4UWS����:�Oh;vic���)�n�+nC�+%�u#=�c�m�%��v�'x:�v]|V��K��&��Ίr���*�gO\.BXmpě=Crv��-5�;Pk�Φ�s�=ۣT]�z8�����u���}�8�c�=��E���p��'n{y8�Ǝ˜8�y��:&�0��i-��i�����l�,���˰�E�eȼ�+�u�n_=m��v�.�\�kM�6p=;u�6��n5�ۨ�|I���.bC��9�wk����o)�n�nn�m���r�Ǭ�p��[�k��VnH;�����[��v�mo\��sk��pE�Q��}�n3�V�Qɋ�4g����s���X�=v�kqڙKc-w�����_�^��8��*iH�nr�<1]F�.�6�֎�ϖWrя�c����$~`�Q-��qB��T=���pr������5g�jY1��獉��3xM�8�]�k�(٫��<��I��(����o���}R�TMR����~^|�/f�X�fz����&���!=k�|��A�[-p7�����ή�)���7�o���_ySM�-PZJ�gm.�/><6�\���ݽ�|\,s0����c$����Y�^�
��I*,�I=���,��D��%*���}���u���[��+��Ed���Y)"�+�bb�"h��&��uO<p�!��b�S�yQ���;|�
[GE����^��m�/gWY�Ջ��7ܬ����M"�m8F9B��{U����G��_ �BdZ�����p��SN"��b���nk�>|�D_�o��t�i���"�����\Ɓ�p;u�Fμ��'��mZCVN�C<;^�]O��E^O5ɂL��iP��M׫j�\$�o^c����ؗ��gޥ���ά�[��!�K��.��$qx|T�ו_�J�W�5�T4${��8^�wKY"q��:/6����1�ֿr~���Rۚ�K���8Y���H�{ϛ��W�ͩ��0��������7�j�7�uU�nR;�#w8�螡
=�Sd9EgU�d��`�g��ۓ���&)�����Of�*C[u���T�ƫ�b��o^By�LJ��%!�T��*�q�����z{�%�,�/7b�Y[��^M�#�2=���:���3���Ӌ4K�ؽ(qEUP��T�Rͦ�k��	��U-.��9>�z@�����X/����;JOW��a��|�+h�&~�6�~�	�c���	T����{�x��{��,O�0ĸs�J��xַ�i���~��6�e*����j��½R�1��7���&o>Ժ���79�W�Za�Va���ċOk�w/��	���B����9��'�e3�qT�LK{�2�u������A�4\��V@/K�0��A�3/�\ʩuHuT���I/[\#����9U괙���^"HUM|�����̽��W
���t\(�&Y?4�޽ǉ��EGҭ�}��t�B��}V��£���)����)
~U~W���I�)*������vY�o:掶�����3�uږ���Н��ɉgSs���M~��Z&pTB�Q%�>�}�W.8�4��J��"1�}�y��j9.E�jȞ5��K��i:�b��ﻻ��se��ͷ{������E ������/��:.���P�m3�z��K�-ls�M6�Q�j�b�4��^��v>5�_g%�����U�{d�>�_	1���0Vf2{1W��V%���]���Xo�H��_My�\4�&��1+����R��pV�"�{�wo�c��MG+~����/�WG���v�~Cp������a)=�,�d�#o��k��#������%���6�:*��7�g=�~�{�7/{�\U7�T����V���WQ�V����
��f#-�-����J��'�08o�:�]��{�܀˫*��u�{���o��������,��5�u4�����Mhw.�<_��e��(�VJcE����)��jE3@���y�$RB�϶�ܑm]oǄKK{�{9����"O�"��� WƼOޯ�d.�(_SεmɆ_Җ:��ĺtKz;'�D����w�}��8/�����V��Æ�.xx�-svh�29���(�E��D�>Z��dX�X��*қ�o���n�{�46��Ҳ�}����.gc���F��җK ��X�]rc�w��J��B���jN������c�����/UxK�e���<���*Pj�.A3I:G�l]�z�<u��۫8��ۭC����
u�\]pZ%�ςԜ�i�W~Y�y�AcU��%+۹���.�0VB�+���Ǿ�j������Y���m��8h�Ζ�m�W�ˮp�*;U�JD�^���{�׾��W���5d�g�����7aFR�"�9kϖ�խ���`�SdK~ｊ�g���O�i�QP��@��_��(^��ZE��%%�K���V� �HĤJ�si��z���bi�<���ڥ�¾®��T����Zg����8Bб�9-Z�q�zW�fH����0XGE�=�7�t]T���$P���}��B���5e]i��(��/����ǅ�9�q������
Ήm4�����y��^#��E\Ʌ�X��ώ�˽�W���t���o�����Z^x���������=�.�D�ܘX.��<�} 0��1U47�4�K��괩������޳T��Ի��o�5�Q��x8�X�=�f��:��򺳺�.��&�����o��-�e4���}���Ք�KL}�WJ7���u��+#��{�İ�4\w1b-���J�Z�믷��2�A�d��m�p��L�љRņ�?_<Z[���B�ii=�K�go���}�d�1�y�jυ/�"ӓ3e�)�!1}�s�Պ��SvB��p��{(��8�)��/a�ò���i��gx��W\������671� ���;vz��cq�v�����ۦ�t����{Wc<�sힹ�j��Oo��_��b����X%ӗ�j��h��������竽wHL�xT@*0]cS߽�1/�^Iw�%"�b>F
���W����)Q��{_�T@�$.�Z/����sQ.J�T�u��5g��1آ*
�C�g�>��]�{�t��W�<j�N�E	�����wŤ�����#�n��!-��C�\}��]����)4���]��/L����8��weR{�̕9��u��*��Ś�N�;IFWI$s.j�,8D�1.���9�n4W����)8�\ܘ���<�xk��{����\>����d]=!}��i��E}��bV~�8�+�Y�Z>>s+�[c0�;GɁ�M�I3M�ѝ5�y�L4��r�7�پ�ϟE1H1��^�s���3�����U�4�wg�w?j��`�E��&����!�Opins�6��˵�*��,�/+�=Z�Ӛ����2ozZdqq�����|}b����e$�p�Yn��YB�<5���{��8�m4B�H�E\ږ/wｧF��v+{�u�]=^���g�[I�s\����[�QBSS1'÷י�>q��I0�"��7�W��f�-?��n���{���d��z��������=.��Hk�SFJ��/�qͥbݹZ�fʵv��t��GRU;�9�*r�w�r���%J�H!�%P��@7=��^�:��l�mƙ�^ݶ;�rmէ��t������P�ֹ��/h��x���&�y���8���Wӻw��� �۱�f�׀�lhձw'�خTq��t�3��\&�\���d��c�Hd;rBL��Ed��u�k�W���A�zŇ\����<1�kp�����U6Kq�݅7��^����@������n�sڝ�yw:���h�꺺�<��tq۔+�k�����\��s��іݭW}߳ݎ��o��/�?����p�s\�T-"�'�� \�&>���Z��vA#�5b��
��;Js�Y�Tw������+,�������j����H^�K���
��[�1gd������4��GO������*�b�G�ߧ�\p�������7��;�JRY�W��;_	�#�'���v?q���T�\?v�*��l��di%�H�Oޛ�]ڠS-H
k��͛��/@� b�T�VU��{�0�-0�UR�\"fe29���ip����w��h���ɍ,�M�C������ϩ �j��d�ޕ�1��v��XO\Q39�8��xTo�1U��;��{x\hu��^²�Y$�Ƥ���{���U29t�L��y�L�b�~�uk�g> �Jjf�}�Yp�n,Z�'�[��=��;]#��%�`�8i�+8����-��b-�.U5͓��|�g��T�<�t���S
M��ۅ�9�v��2��5���,���#���P�ra�>�W^�I�.��2��<+{T�����O��/v=]�V������<!a���>��N���S-1z�YB���L�LҊ�vط�L��7��l|e���I̒�Y2�c���.��ޮj��ǵ��怫�1L�z�t3	HV킒[:�����O����N��h��˪�����V'tJ�R`�kמ�����;�J�:����g5fy�3;��?X.I�zt�nf��	����O|�%Ċ��B�/r�a.�G�lc��D�TVZ����\��:���X� W�w�>��"t����Y��(�\�������P3:�ٸs��j�h�}Z�]�t��Sݰ���.�!�k��i���$�*�W���7�I���yX%�ّ�*�@nB�����B����D����)�~�̹׶����V���ފ��o��R.s�|D����e`�n���}+��*�U%{�[k��M����B�DH߹�,����=�S1)[��4
}�A3�������H����ϮI��wC��Ͼ�x�o9�%��-f?y���㷳} s9�/:��Q�ȓ�ɠ�zy:`�K��n��DO��-X���|hs�x�S��/��w�nİ3�ڽ 8$�!��\�@��e�	����n� �
*�@j�y�^
����#�HT}��G	�Q�kW���+6uZ�|j傹CK)�q�5�`�����UDSC*�f�m��j�X�����J�: ?O��0�?��Ϲf8�5/��75���N�f��ưn���,$@�����`{w1Z� ��%Dr���e7O�<��> ��p�Z}mY��{��WyŘC�AS��j�f)�v��g��z�t�j�(��esN�,�(�霻]uUDT��JS)��رa���/�%�^VO/�x���T�1�D�S�	�et��{5f	m�@Y �!9}$�]}��\�����(�
���m/*#�^t���h]�H ���$
���������"m&zu?�'���� ,L�\4)Ӓ���Us�!t���N��M͝>��Ä�%W���G�O�/�3_^ʱ	�4�:܈��z�4�\����$:���+מ���я�}-H}^�����~�}_G�%��'O����S�ߥr������n���/c� P�zpX`�ft&w�׸���_�8q�|�(T#^ca��xf	s\*#�w}�rfkVu���ޭ�W�m����ūx�t����7K.7e��KfF"�Q���f7w�.��8�����H��l��!m�R�7^�wf'�h���W���i\�kz�,�a��e,�����hK�=uXU�~����b��=��tHO���dNO��%*FJm(��w��]���ߺ�]�}�ϟ��hX�*T��\,ץ���{^���;)I6���ݹ�཭�U\��6+*��>��uZ�j���˖�(�iy��{�����;�߻8�ޡ��ݾ�'�pr t8?��^�T�)���z���O+y)H���T�s&Ր��(��]˅����?���ԅw���Œm�Z��89L����<..5Da�4��}�ZA�x_S��a��j��F�������N��N;�(,|EZ����K,�/PgF�li���+����S\�w��6i�xv^+�<��e�ݹy��4�*:��4~���|w�Q���g�_�]r����*(]mf9�`ċٛ9Wu����4��V.
�c�N��-/zC�w���UZ�����U�E�Ф�j��}�׵�Z����89=�������ҵO5JՑ���Y"G�֖&8I\�=������6��;
��+��ۼ���k/�*18�'�aC(�N]�_��V?8�tZF��T��g.���=q� w�_no�'��н��"Ǎ0S�ց;"?(���U�f����'�4k�� �(��7=�}�:/�"���uu��3�}�mc��v|�3)Qd>O�2��������]y�+K�zus��/b��5��9�ͬN�P�Co�K��{ـS��G՞k��P����Yi�im���G���1���gs��O� ����դ����ded��Ǥ?{�Wם�Da
յ�i�r�U����6����v�D�ᇉ���wS�����U��(4Mܪ6�֍��o?�JV�ͧ�t�����0Z�L��(��N�R�2�o���!}1r��}gǞ�:b�@pJ�'"U����8�o����;T�Ku��Zg�u֔�t(�Tx9�q^	��M6.�m�!-O=����ʿ��v~�����>�[�d}lC���]@�tRx�gҬ���S9��ᢑS|rb�c�oү4ixy=Z��"�ҨT�v<G�����^(�ݞ���q����X���mu�o��jJ�*+#�V�w6%��φ�p�6�}N(
��~U��ƾ"� ����,fg�K��h��xO2bP��/r}��s��m�,p�u��k]D�/��b����rR�}���~sB=/�/�~~*�#-�[i���\�i"d*�}��V� D�~&>��sgɢ߄��>{p�p�j�琳�&I�����ij��\�ƸC��bW��*���Y�6etd.E�ފ��)�y6�Eݝ޽��k%�U�e�|i=�h�cƕziJ}w����w�|3�KbU�R�E=��k�*����+�a��֋Q�����﹧��S3�|%%�ϔ��#��rrE���._��ZZ`>9�}sm�|���������Q��yش��������H�ui��/�a}�Y�/Z�!��a+��UЗ8׸�A�s��0N\q���K�o=5x�|�l���:��;ޭ%�ƺ�U�(�?IƼ�Zr˕����k�ol���ƕic�[�����/��l8���+B�jŷ����T�K3V.{=�N-[�I�qE��B�}}�}��+���}j��ծ�v
ڒ,�{+�.���+ǧi���
�,�:-Ͻ�|'N�K�9P�"g�P��J/���^��L��ɜ����f�n[�e"4E�lpH�ʸ���K�Q�a��;�M	|�����Y
� �bޔ����r�&�&��w_�����i�ƚ�舫d0:;�%��eD�J'��q7qPt���U:xN��a'�Z<��-��Mݻ���_�2tSŵ�8NZ�p7��ʼ���p��ؓv�y���0�Ѻǳٯj\Ѝ��ܦx��$��n��ӹR��ݮ�uq�=�fC��1�zv�rFםĆʜζ��`Cn�
��g\���c�(��%�·V�y��eylM�g/\.X�:v����l���g���\n|Ե�\�v��F�:�m��$��bv��]z���-?��5��oL�VV�j��i�uژ�~���a.iɆ���F�|��o&ł�x%��ܙR��V������Wۢ�}<�8�,��9�v{Q����eVZ�TA涍�7��QHK,�4+m[�q��P��k�p��<����5W}7�|�29�nM�#�s��ix7IL�[b�*\u
q�D���x�/4]�X|G-����j������p�=�h���5x�ǈ�+!{�ξKN�&�UD��D�p�K���RG*�)W�{����s��!Q�(Z�������y�E�ZX���z�J���|!���p�!_r��4f�J�L-����]u�HC�bD�@����ۧ�\����`��b��m�v�h�k-�����=��* ۜ��=8����ZF8^œa��"罺\,�5��8+"N� r����J�=��ZC�L蔪i���f�][L���t���#�3@-�+��_q�ز�	8C�</�jf*S)R�m�N`���MY
�u��y�^��w��� _U��"τ��q�U�R��	z>y����uȖۅD&��_���da���'P�	�ם~��xa�ͧ;ׄ`�O�O�Z%(��x��c���O��F��d�xs7�VT�޴qS����o$l�l�B�9ނ�u���$��*/�Z�����@�IȆ�i%���]G,j�t�)eF�����,��O�1���
 Y"��_A\ͽ��$��?�o���Ǧ�RƑ���ۜ��4\�3k�İ��̔$��Z�*,r�aHIqi��o��Ŏ4������5-_����Z�/Z���������ȞzdI�w6�R����q���b����+r����)�̏�6�}�
f=�ffܻ���[����|���Ƌl�>��U�M�g׿VB��8R-�M*
ci_�g������JD���e4��nq�	p�]���Zs���jo>��a'��p�P��G�S��4MM@9�Y�Y�\�T�%G��	�מ�`N����@����\
�oe2ń��x��]V�EkZ ���ϟ����&�h��8O�޴��rˎi F��4�#�1��NK8��굍8�|F�e1!c\0Vwy)���xKSLuH��B�&�n0\����&�*����JM�����}9�/�p��ިIF����Ұ��iB��<Z�jG��(	!9}�@�^�ŀo�z&Sj�T)7���RN����$�^�=V��bV��h,a���x�Ƈ�ۮ�Ӣ�%N�֡�9�|h��l�6�'-);���Vތ�L�GRo*
w��ir~�lw���\˹ScX��
QHh�U�x�=ߓ����He�B�\�X�K�=pU2}�x�;MJ:$��rZ��E�f����u��Ƚ��~�o����#(|�|d�k�k`��<Yf";����kr��}����Hv�r�OU�w�{��R1������+�����F8,�0�e4Й5[�}[��9֗K"DH��x(��x:�������_�~>��!@x��I$Q���/�B�$Ho�����x��ㆅ�p9 pr9U@�4�\`��Hu�$���<,�`�K����������o�U�!�"9���}=��s��]"�.Z�f���;����X筈 V�}J�kM���8W~�V�-F�ſr���T*����K��L�,��v��n��S�D�2	n�[|���n�����9q��s|d,�gks�"�i�(��&e`o>�,"��LG��c������U0����s���VT�f�xk������+3w��]s��cu(���Fe�i���G��:�6㥶N;Tk
�\�X�5��_^6<�����뤕�N�r���!*�Ѝ֮GO{^��%)ޱ3w��&U��ȳTu:�G�u*�
�HSy�i�.��]W���;q+3�=�y\��*y��EN�gD��\��R�[��%��qm��a�	�{��$�!�L�8����=��Ix����3CM�Y������2������ԏo&��:lo.	ց�J�2�hwy�z�b���N�0��L�Cж��,���t�{
��*��1�wH�`}5kBP�<3oz\�5���G8�[V赯aT��9�w�;���!�12k�˂��KY�m:�5��\\a$ѽ\�4��CV�i�nt9َk*�+i�t�i�(�6���6��΁fScdWzǳk`wy)�;=o*3�������6ɥ�V�����'������^%��r微��@�>����f=��@�+��'ҭٷ��+X2mՄˡgk��I�����Yd]����xcp���ǩ�E�q��0rHs��R�,rӜ�Y��t��7*MϧQٛ;�t}3#p�G+Eq�O���iw�(t���]�2�_Ny��b��u�_a5pw^���&�5�d�t��i���ǝ��kq��]aV�W��Ȏ���d��Wu^2��N9ۣ�Z�֬�R܏z5`�Xw�j�4��Q�W�o^������+r���V�E�1�I�Ӣ;_Mn���t����7��]h"��+B���me1QE�f��z�;S�q��}�U�W�n���%T�����B�ML�Û(��=��O�T�BX݊:J���k��
�BGo��|U8����,�o�����|9�Ja��A�� @_=�V�频���ܪF4�Ɲ1�\�6�`�� 
n=3(D`�p���Qݪ��U,�X��~��b�\i�IX� E4�s�n���tT	I	`�*����q�C��hl>�������`�ְ��ܦ�\�&�PTa^W��_zP�<r�0o�d�&���Ul�_����	g��������ؔ�0Rኽ���,0^$t��8�Y)�@ŕ���d��]~yp|7���i[�%ɝAڅ�5�k�z�u��K]��j�hvzxN�A��H4�����r�${�A&i��?N�ܬ�O�؜M6!
s�+� �	�"9�ެKW�n5M�l����R�����32���eNк�h�&S����Ӏ��uZ��E�\�T,!�ҹN@g/�_�T��D�T[m�[}y�Z)�P�'����-R��3L��9-�o�'��w��� �UR�qB�w��}�����0Q֪�B�Y��h^����6�&v���ܸ��ЄM�R���\ �¾W�=��w[�<{�tι@-�е��Ѱ T�	��4�L_���-�ɹI�BO�޾,�0��Rr+� ���m�,||}�{�qb�:� D1l緪k���Ϲ�k�o*ד>l��Ѥr�~�Xp��4 Q	�m ]���
ϔ��^#��9�hX�D'��sԩ�˦)�T*ыQ��A�!��,�7�K7��~����tG�r���]���#�(V'���S�|iZ�|�&���ڹhGZ�m2��>���z�f �tRo�T(P���*+�V��u���q*X����.�4UG�S׫��v�wF�������j�P<�%򍌻��� �}����/z�4�q��j{��a[��ZY-�׳�ɸh�2x�"@>����z?&�;h1�UԺ�פm�\�Ne�L�Y�i��5���w���}��]60�.�Q, ��}��}��/�3ݮrL＄��V�֙C
Zdq���Q3��^"3{�}o��֨���#�e���0������R1�h�LF��g�殟��Nl�M^1咖8rT�4�n�ɛ��C�[�eۂ�D��g�]�n�����}Q�Je533S���L ;�^6�
k%��,d���������"�v8�Gm�MI�}�X�ǃyڠ
k	{�P{�$\0҄.s٫6�;���v+x{�����?u؃ f�i�b;��g0��1]i�i3kL��n�ۻG����s�]�+�J�$�����)�)Ф
!���"��` �z�sל����PpϪD.��*�w���ﺭw�7&��Y�H�� TQ,`W����3� -P���J�U5�x���j�8aD*���i�D# %�����S,��M���a֊l@�.zJ@���m:��U�"������}ra����N�oճ�N| ���� �Gg�uk�}w7A��D�#�� ͮa� �ۏ�(�$��Q��_<Z�Z�I�eDq5H� Ѣ�1�d�~�����Aʴ��{���&�5Ӂ���&���M�{9ϟ� @��%=�z�E���Q�jLƩB��͈���LX,5$S~���fK���H@G�sڱa��ۭt�Ǝ�/~� i�+�c���y��`�/���՘��� @�IL#�acG��m����K:Kf�����T�Nq�4�'�6�>��8�͉� r��-�5��>�Ͼ��Y�Jo�Vj�G|����|�LAD˂���k0�Nʛ�͔��}�n�񨎝 ���6Ӣ��*_m�{�����o����9����L1�%m�z71��@��J�y� �8���,�u�QVج�bȺ�g9q�� �c�ٸ�Ѕ�nX��2���b�m��\c�y��-;���rk/#�ڞ�v�[�q�s��m�2/�]�|>���o�u���<�5�^q�����-�e�̸]��0]���}D�๯[�Λ`�m��.ջ;�*��S�� ��9x�S����໮����Dm��ݸ�d%��y��Jdi�	�x�.t�e�L�7sks�'9x���� ͙3�eݻe����������s@v�2vq�-��.ݫ��W�y����pa�uUM_�~�DL��ɖ��E�V����\���}$1�{��aM��RH���j���i�nX��S�����E��3�{�Ɉ�ͷ[��o\�șDa����]������p��)�f��c`hř�T��m��l=��mb�K�KV�Z\
geY��sƨV4p`K���,�83>��?��4]���y��6�w�B�8)��l�D�@��R ����0@�GGe�!�����A��������^� P'�ݾ�ǫrq>�5q�Є�������G2"@��L��P��Фe@�o�����g��1!pgnf,b �ܚ �r�MN{�8�����*��C }���@!y��@skA�-s.� ��Sj�����ޫ� 8C/��i�/
L�}�g��͔:mE�#nKM�����fO�G��;���Nj]m03�ϻ�Řp����<M�\l|��
�b3�{zf�f�Z)��52������M]gޕ�>���4i�^)P���u�������,[?ou��ei���E
�F4n�zU�o�~�G>�`�jŧ��,@�;$�y�J�� �*�7�w5�s"oD�԰R�����$'�|v����z��+Y -�\G-0ܕ��XZ4�X	m��皂��C�W#�*#,u��,B�{5f�jJ
xI�"E����F
�ue�u��g�˳z�I���g,�B�d��s�7f�gu��5�������-tO��Ԙ}��m%I%v;T-���?��s�b�Koa�C�V'-�8���in��Y�Y��ՒE��<^��wY��`���vR��j���y��v��hF�n�/?�� 
w�昺-A�	��)���̌m����8�c��ڀ9+:�[:͋��T�L0���.傶�<�fw9�1�F�ʘϖ�9��we�%�RY��/���OқБ7���MU������Y�ua&���	��tW�\�x�E?��X�(}�8�5b�\�A5[Ř��ne2�����O���>��k\n}S AO�j�[K��|nߋ���oU�ƀ�o�s}<ٹO��t�}���\��\  S��I�I�D�j&fj��.�tX��Ċu-t�Ӿ�|83�NEC��W� @q��_{��,]��
�0f�H������_wٽC}��P�۾�k��b���,�sYo��6g׾�ŏ�q�,�fD�[b�X�{������9@�ez�mװ�J�R���\=���xs�K��}�@|6�2�" ��l�r.���yb`��r)s*ϊ:+%�.e\����/���	���F���������z�bo�o���GF�!�P�Ria}�ٶ���,�V�܊Y,N�G�p���Ig�� $���ⵄh<)�����o!h��Ͽ=���ϰ<�sv�}|��ZXH���A.>%>���o��U������mH�b�~n�׳�� !>������Ln���}e� ��%}�8ɻ��[=�Ѧ��y����n�͍v��v�Սۅ�f��nQؐM��{f�����1)&Z���v�X15��7}\X� u�^t"�0&�hA�	1��z��0�}��Ik�s<����A~ϵb]����e�T�Y�=�޸YG7U�Z�.cA�yI�%�E�8-?�s�?&/�nAJ�#rI-���}�G��X���O��~�͵�94������Wq��񯲸x��~i���\U�w�0H�`%�y���0l]q'ޮqZӇ[�4�xJ�0�%
�v뵘��j�t��{=6��c��*��'�r34qI<�-D:�f��O\nT�i'���@�x�O>��iN3���Ԗ#��)Y(X#m���ii�Ԇ��;�]�o�+�C���)�����{�\À,���¦l�ќ؞������tP3��+�UY�,Ѳ_h� 
|�Z?P��qj��H���;�2�tXF��mH@���wǹ�ש�1 X�).K1��i�����V2!Z���Xp��%	�/���n]��<}�yD�V{�Ց���
lV�L�7-Z���^/
���Y{T���SAS�H0>�s��vk������d2����k��8j7���|C9��V���J�2!��7G�n/Ȳ��P5KCM�H�]����ZL��o��Y����B��H��*@����zX���fg@�<y�HC����ট��R���^�o�He"�[Tٔ�쐑)~��.���k�$�i�"�b���É��Cd]JT��C��8!�^�p�^{l��o=�SAu۬����Ԋ���ݴ�9Hr��{�=���&84t�U<nik8Ug>��4g|��E�H�\$[?g����¥lZ�I�Y�"��jΑ>�뜑��sVF�
M�Am-�Խ$����p�^��b &�E�N��� ݙ�.ԡ���2jf�Va��V}瀯�ꘉ����92~��(��/Ga���\��F��(��*�o�Y��*
�_4�i��zU�˿U�	���ؽ�v%-�����
�����$�m����Z+���������Eb���ֻ��؊R2�-�KmVlC��*�	J����5\.kO�(rր{,����C���9!{��v�q��Ϫ����5'���a���da�J��е���ج���{yg1_��|dqF%J���LI����j��v���*�T�9�\���]�P"�X����k����R��J�@^����M ��)(����Z����+S�!e�)q����k�u4��ˆy	Q��W���;�����犹��I�܀b�påTU��!�J�w֩��5e�����U�ҧ�c��c)غ��bcV��v(����0W��;Օn����⢠bf	ӳ�5�O����ᯝ"�8�	fj���
���U�����Y�k��i2\��%�D����;n&ƬEG+�{��^<�Z��D}�L*"[N\xSO�X��_�b����	P���b_s���%���'.�!�>�~U ~\;�ڒ4�%������]..��A�L�YgX�n}����M<y�8��P���N��ߛm���w�'v�7���kH�0����Ő�U|�Ӎ4��SMAt,�к��qoi����]*N>�d�G�D�	���\�7��?n�.�#��(VY
iГ��tŧ��r�a���m8_ywg>J�����i�^ۢ�X&y�>�)��N�Z�4Y�}�������Aͧ��|��*/.`(1�����:̬d���\(�i"�h�Y��p��{�Ӊs�:xV,-	M����,3�?	b?Ɋ���"�ί��Þ��k50�κ�?�'��%�[�C��K�u�<��>�I8)���{��RF� T&P�JQD/���p����=�$s��Ҩk��r�!s��� �m����ᘊk�,*�	qr]�/��H}�uZ��c�}�ʫ�Ҳ,�Z�m��7�l��~�D�m�΋0� C�zv�sC�1R͎ P~;��׻�Ub�P�>&'�X���]n��=k|�f	ID3�������5f�|�es�2����K|{�ߺ�-ݕ�M���P�++wߜ���%���E���(ִF��o�ܝ���AiS����|��߈�����'��L�n���G[Z�T�4��|����S߽���)o��T�����+��RX�i ��a��eX%���
=ƨ�� �By?g��Z,��g�bEE
��9��cY��ޯU��/�(W�2n�j[�R�jJ��x�F�+s]F�do����L�4�vv5��藝m�-���&����+o�aY}K�J��n�VK9�:�Wi!J���n6�r�Q�����f�q]�[]s���y�e�H�[�뷶Σ���"����{p�#���v��ꄴdx;��-2p\ۮ�ۮ{p���nه�εw&�����e�Pd�s�\�.7\�=&�W/Cd�nK�I�)n.����ZA�nW�(�n�,d�]�8���@�,qӣ�����$Yz�ۗ�]��ݬ�ZxM۲N7O,&E���|v��9�}�v�\��"�:��L���bV��i�J�&�$9������;�����x�!9o~��;����Ũ��-`���'����>;��U_Q���,�9����Ϸ��z ;�����+k���r n��i����uZ��b�
���嵅�V*�y�m��hr��"���.B�mm�ȱ�ЀC�2�ӽ�����p���Љ,r���3�x_��2���-)8pJ��v�Qs�ⵀ}K�<�W�6XYb�,f6�1"���\�ى#E�w{ޙ�����o�YX�������k!�Tj@��[�?���F�-8�j�,ȓh�������V�$,��XF)�6<�d�M݊��u�B�o1��d�S��u|�>4�!T�Ż���(JJ�ŀ�7�|p�ܿ;GΛ	��s�W1���$�~�����C)K&�4��A�/�V1*��9�wk�eq���y�롛]ߕ���(�h��ݴ��G�׊�o���0R�=$��|�#O7"��c�/^����{}s}�8+~�U�����B�p���Rt3�$1g8)�*A
�)sK�Eg[V.�fWd o���O��,j�TŐ��ŀۛj��G�;�r��VB�k�(���5��0�H���+�'�=p�}�%����p�^���x�"�deF�g|Q�ƙ�~��޺[�J	�L�Tm]��q�f-�n*7��n����띦L�A����|�\U�U�@c��|���Q������0\p��O��s�|[<1QJ'o�ZL�})���,J����%�T�B�Ac�d���b_o���w1g���<�7�<@��׍p�I�=���5�������x$7C���{���Rb�%�_.�t^�O�7�=�����U;�_E����>֫߶���aָi�F��m�߉̏����KƏ�1J�a�u���l�:�S(����#7��W9�({!�}��τ��5��s�*��W�)�Ml5TY�����||!��1IID� �}�za�iBY�/�Z��-틠in!��{L��ڈ�����Ƭ�ȱ	I{�j��h��I�7P�-x�5�7U��}څd}�t�s�Vc�Ϊ����q"����(�͝�s���,(��jL!�r�
J��<o�I���E]��o��r'���lV�_�_��G�������~�4�7��X��Z+���v��kC��YC[VB�>��'�������O�nQ0]��=�-nO7��s�|�<���}w:Ao�������ȥ����6�Ҿ�\q왳YM��%�k�����9�{M<�XB�٦+��|,�����ﾌ��ŦGyߪ,�|p}�w�� K���ݮ+K�r��y�y�l�i�ϵb�1:E��\�����/Գ�ls�_s���nZ��~dU[r_����� ��׷����p�rbM���3tn��9��庚�����D�z�R,@��{|_H��*!s�1�6ae�Ls�{��G���+(W�z�
<h�O��}=�u�2�/�/����\>�q���.�뫽|����B��Ֆ&G=�NS�`jT��SC�-`��J�ĸN>���s��w֮k_W�ѝy���$�Oo��=�W��>��Ր��Z ���W�p���=Sݛ�tۙ��_�%���p�G|.﷥���H�������p������}/~������H�
��*��oo���8B��)�*y���b�5E��)��/�U���\;�t
�{�g��0՘���SҚ����rˤz#wL�.=�w4m��od\��3�uX!��1rJ�ݔ�g6��k$�ݾ��D)+�s�t��9!Q��RXC6^.4�y���n��9q�Q	ˏ��i���s۱0ܔ�b�.�d-�I
C�}Ϫ�/u1�$w�w�Y--(]n;?{�1,+׵ϯ��"���Κ/��>��X���综���P�l�=_����c��VWs:+�շ�I�U�?��˳��]�TЪ�jBK3���Սx������K��}�訅b_Hoy�ݢ}�Ɯ�lS��p����[��ф'o:��o�ՉJ:B�~�J����3'��L��B�+�'N1�,#}w���O�z�K��9'�8vp�$�ĝu���*��v|�����Ap5�۫�:�K=s�c�ܟ�Ÿ����?#���\���W���ذL��&>
���g_z�,]�¢2>��Y���bGv���Tm5��W��x��q��aH�+
˖9p�O}�u4F;*�'��V�[hcC��U놃"���{��>z�b�ݜ������?�&2�9;�j�)]�£��d����r�1�{w����:*#�y-���D)�r|\,!g�Ϲ+�.iS\�=�|֑���*�R�SJZc�Y�5B^,bRGu��s��.vh�S�����¡M��{t�Z���'�����E��KI�W)Z_!]=�Y�_<�yŉ��D����3
����|�K�>R4�)��T��-��b��~��{��X/ܙ��~/��y��\2�f��__�_�j~`�J��G�Y5�{W!a	����{�Ru�������Dc�s�#X�x��Qz�[�Mu��*S���)�L��t��%��^�y3����
;�}�_�A�{�ia����Q�|c��t�R��TbXi�V+���E
���;��p���]�
~�)/�T��}�h�lo��zGI�v�-�!Y��+޻�I��B�JT%�����j��i�-$W̟
��MZ"�ٞ��������40�k��nÂn�&{v��(�<x^w<�,�&P�;��X�jxz�~����ԋŉY�8����.�pRD�����KS��*���LtX/��v�|p��\����-/fZy�ݮoH�Z����<}碲9zծq�7�{��B�S4n���{ts�J":��2�|��CI�ޡ*�d���o���Μ��[/s&!�_�B�Hd�K��I�UTG��Z��	04���TB���jH���x��_o�H}BZ1n�d&��1o�Pª�	%1�l��c]W��H�����:�E��RB�?}�+�x��R������f��WL>i�rҕ��ƕFMN%���8G4�g��ƫ�h�s����?��U%�-ۙTP��k�z��	a/��Y��$�!H�W[�r�K�)p�Y�a	�Y���yʭ�}L}DU��SZ��F������*z%H��������;P��ErU��Ƽ������B��wn
H�@�gՕBUu֎d?�5�L�gL�&�M��iNT�+ZRi(��]+Q�貚K�d/�P����$�!DG�P�%
"?�(IDB��
Q�#��	(�Q��	(�Q�!BJ"D�%
"?�$�!DG�B��D(���BJ"D~�%
">�	(�Q�BJ"DdDBI$�@�DD(��B��D(��!BJ"D~С%
"?t�%
"?�P����(IDB��B��D(����e5�3��U͘ ?�s2}p#��u@H �cI@*�����U(A*� UEPR�\�:["h ��h֚��(
�J���R)!T(� �@ (        @      P� (            �        �{��'�=#��Vƽw��R�ʦ����l����::��Z7/ �u�!�z�X릊��;g��\��uТ�����8�� GE�����v(���� �R�    w�       �  �         �p 8�tѶ0�=΀+V���A���m�=�i�[֏m�uvnw� ��:ƴ���`���qB�'��7�==+֧2�yw[e��	��@ �    40�cB����T-�0t�����\�K6�p ;��7&�J�3��
ܻ�[ ���P8 㤵�nn�:1�s��R @
!��6mb�.cvf�W �����i�n�Ph785�U���5��Z8����fح�:'f�{�px�f�7.i�b�g���I��wp��mU(Q�        q�-f��]d�5h�wi�ť,�k5����uU�֕� �:i����b�tS�l����V��㛦���p 8Ӷ��gc@�`Q%A-���m�f[6��.�@�� �u�X��w�"�s�.�G6:��K��"�%` 07e5��*QvmˇZ�c�k�mbk\���U"B�B�2p        �N�E���mM����:�@q�Z�ܷhhi�� LQ���(]�W;9[h����m�Css���T� �jl��+��;h(��D�Q[��u�d[�+�kJ� ��R���\(�+��m%T��75*Z�,�JP`  t���F��öe��-�KZ�\��MmJU(�     � �˚F���EV��:�-gH���r�v!� Z�[M�9[,�.wJ)t��`�!��֔U%� �v�+\l���c�v�T 
��T�ʺ���s۠		p���Y����ح�A��+k nwm�2���:�G ��!��DP��kis�EE���m��2�T ` )���5F 5=O$(��  ��ԁJT   D�*�'��Q�  jMJ��&�����c3w;��\	�E��Md�[bP&pB:O�2��U���>I����ef��4�f93��� �@�l(-���II�����	$	'� $�$��IH�!!!!�����+�����FνO�����f�x-0��W��*U��9��G�IR���W2�6��[��۽�MŶ��i�lZ/V
��'�V{�"��̧, ݚ�ٖ�ZΛ�;�ZP�e�y[��)���*�g�<A�� ��3��nŧ��FSf]㫵9���v�J4b̓$���ݵ�rZ9�n⬒\��|R�2���5�ѡ����[CuF!��vʆ�S��MD5X��9Z��.J�M�#���*�&I�T�)�R��k�)m��0�u��AL�to2�I�RIZ(�%�wEL��d�%�K�[���H�>
��N���z�1�fA�#p�vh�����L�<ll�0�������[i�A�ŮU��3q�$�w���oL�i��[�dCj�m�.V1B�����E���`�+E��L�r�3�#U�p^��1�P3.��wYy%c�Y�;�D�a��٪�8)\{���� �dJ9�,��Oee��>uG�g"X�٨Z���m`�3�x	�����[F��
�!cF�,8!��2�ycj��Z�n
�5��d�f�
Ìfm�ddf]�)XV4��5u�_�p:ש���2��j���3&�.����¿2�%P<+q,�����\�}��û�{2���p�WZ���Ȗ�K��I�f��F�Q��ȟ��u=�Ě���U��2�Y�l�I�-}~�+��4hb��P�i".11d��*aA�^
uyQ�K>���z�6I� ��w���a���:�X�nV�+���N�dl0����+Ճ��d,&H�1�hn�2�c�nEa+�n\�&��V�Q�h8��B	�K�kÚn���4��|F{��y��G�TC�����h�Ǔ(��6���ڻkl�4ۢb�m��գ@w]�yjd"!E� 2�x*�u��^n5�BV`Ux7���Jh$vV�%��m�*:��[��ˢ ��>t�h�kۧ���X�Sx�R�W0�b�+q��+3A�t�ma��O���tvKZ�� �	e��Em���Q�f7�m��V/PK�K(�y�zY��-���`�p���S/8����n��h�'�_4�R��b��_�U߯1��I*�Y��
��4���'-дs�1�,���E{��&�C{u��u�hVeE�f���i�h�ٳ��[6��^�e�xC+�Q��	o\�-<���*�F���і\����i�J�a��Y�ˣz�A5�����k��*��{�Z��N>1t��i	�jd�+.Zv�i�(�Ԏ���^���̊�*Ӱ�=ۻF[�OS�B,+�@0=�V��B�c���	9�=i��mno+��{��ŗ`���ӕy��d
ƚ��id���C(�����z��N��ǿ]H�
79�)9^�z�Ay��3�s"�V�t\Gv:�6���PU�@���H��L+)	�#���ɠ���l����jX��d9m ou���U�4��ң��L¨�#��6��H�̬��G�exO���}����#	n��7h��sC�K4�gh��f󉪛ܭݬŎ�ڑ[���&�	AC��j`*���hmiB���'0�ܬ��^e�a�юU\贞6��#5���G#;�|��V��Vǆ8�X6CR�W�{SLg�����2�k��)ejH��_7cp��Y�(^���e�!�ѧ��m�����4r���6�Ïg��\����W��e����W�Z�W�`�oځ	@-+�NF�e杙�����ѳSRqQ�2:��'P�������şD%A!oT����5����< _�b�XQ
t[�Y>�Jx�3<� �&%��- �v���f��Qw�p>z�Վ�Z���.�F}�(��[�Pm���YZF�Ȭ^�R���YT�
�x����W�ƓNjc� �Xj(vQ���1������j�S�T��������w��yZ�J7�������X�[R���
�3
Ցh�����<��-�8�c5t"9p�z�y@I~��{���pv�'I�++��;��^\[�� 25��7m62'�nz�̗�w/HS��!�t�$��x�5!�
�Ն�jT�f�4�I7.΍S�Ǳmi�(��ʽե�Jj57$��ѷtW�v�8/[52��I꘯t]��4�nm3yp&�2��Ym�Xb �֙[��j�X-�)�EF��̩u��Y�ԩ��N#m諭�#�����-�"�)ۨ�ύ���L��.ʒY<���`��sּ����\qfQ"���"��2��U����b�Vh��7�^j�dR��J�v��{�+=j�u0Z`z�Z����ٳ�;�f��!��@�[%r���U+U�P�0�}W�H�֕Ǒ�g���3�6O��m�!��*;w`�J�)2O��@�+�r��8|��YQR�2���׻J�ۈ���PM�v$�ՀV%�`�sU�j�W[��ز� �z�.������b����&��4�ec��Hs1TN�Rj
��K^�[n��Q�V�֘zw�,7�F���snZdK� m��`W3,2�jZ�B�Ʉ����2�A�rV��,��u3D��74]��t��,��輶��٫�*t좶P�ѧ�W0A��ìg�/0В�!q�9��U�]꠨]+Ӹֹ#"��(�b&��iS@���)�����o~h��ǠC�>�uc'�3@�i
8��7�5�Y�5+P�wMJ�<�\2�V�#w�&U��;��]I��iG*��aX,�t�^BP�էl��v�V^V��e<���� �]�ld��!�y�eZ�B�������������#bk��x���ځ:$7��b]�2`:�)�0����x�ICl�M5�GG2zB%��I�&xJ�4��>YXJ쥫31@F�XPw�Za=ɷ�5*�am�2S!�
!�lPm�@�������7"�o^`�-S��l[g���!��hT;s*f�i3����%P�W6(�,К1n`�gj�*���f	��#wHMT�7�OXr0�^�2��o,�0���~��5�3�q�����K��Pf��.��j�Y𚧋Kk��Vj�rlc�B�VɏQ	^c���[2M����4�8�i�pVM$�un�cSwe(���+�fQ�tp��&+��[%z��Ei����M�#9��E<�S(F&e�ֶd�û�����6�YQ��fb�u�]�	��mŃ*����y�ohJ[1�Ɣ��}p��]ZB�,�G,Tf��Ͷ>z��&��N�{�r�V��ؿ�0�6�g���9$Vؿ���O�t��][�øi#[�j*�9t5|��a���a�^#13���7ײd�@�[K6�r�Jf<��~�m5uwNJ`��n�M�5��ɕt�F�%�i��q6�lԱ�ՖP/1�m��Un��lp��$�WO~̤��X�r����fg��O�3Q;b��L
;���	e! ��>j�Hq��'�񫆀H2;��I���- Uh��a����E�5a�7�\���&�Y,f`���|!���2�֤������! �iؼg��Z�cq��=r���3w ��^�{k�M�S*j�0�Lm[����ن�]J��� R�R�6�6��{B���7���H00m�b�����O�}z2K�8^�e�Q���t�*��G�Ã.�B�K��tV�����o���{U�������ɴ/ts��'�S䓍�en����5�G*٬�%}�^̦�/-�/�]���wv(�,_s-�O;���'rٚo�I��(�5:w�R��棹�!x�4�'Vs��o�ט�1i$�=%���pĆ���I�)pZ!^I:x��lw��I�QW�w�K*���'OB�R��f;(�S���uV��-Y5J.��x�_�->�M��N�V����Vx�:URJ���j��k��Nz~6�i�q'@\�|4�3�|9��8���tZ�0���:+���}��.��JS��ٕUmѭ�o��U±�"_ϲ�-+�ֆ��s�	�M}��Mmp��i���"���.�[�vUҫ]�NI��	v�G�ƭXF�*�bY0��]��V��kL�DR�n�'{B��+�.��t��L�4h:̨�6�ʽ*��a�
��+ޕu�[B`(# �VAYm����6#o&L��m-�r�S��R�+n^�赸�x����aPyWg1<-4�N�Z�.�M,`�D��r�v��eܬ���6-X50�r��:��V]�z��rc݃~���c+E�4j���Vn�4�0��Sr�r�����(Rר�MҀ;5=AX�ne:5���J2�p"lhIYѳR�mj�J+������4���p��x1���%*Q{m�X�z�ܛ�.ݜs2��u:H�]xx^e!6+z��]�M�`���m�Z�u�ν>q#��A�*%��)(M����(�%@�a��Y�F�R�� T�����?^�X����b6V� c[	�N�3uSt*�+��ʕm�E,�n�P�x�_y�.��l��x�.��Rʙ�^��}a�x�NV����R���^,Uc��0m�ĥ�$St�YmK�2���E�t<�(�i�@׫#s޲��%�`��B�VSȍ
��u�]�fk ʏ1��]Cye�^+ef�kq��[��/.:�.sWMM6�B�5�b�q*�j5�-RoX��`d�B�Z�'aJ1]�;�Vȴ�����(J��)��n�̴�F�P�b�N�2��Qw�XSo�B) �)e��C �Y�8j��A(��z�2�o�S[�ri�f��(�5q��m(l�Lʕ��R��5��h��![��d��c4��쑦G�dTx)��1ya��7W��+��	z�8���iݛ�R^�[�����u��D��g��/�Fɤh$����W��t��q̥tp|v�,�@��[E�6ց ��� �=��/*(eԡD�h���Sf�!+�o]���y�hM���FQ��Eأ��RZw5��ݭ�c/!��@�(dXm�Tۤ, 5yҗ9^�]��/�p��4)ݬ��OT��p"l4�U���R�i�[պm�;+8��xu
�)n�*��ڼ���c�r�".�ܙRQU�������D��\�a4`Vۂ�l%e�<Ѷ��(R(oe�J[��腭��R,�U�J�4�Gt��'>�ʽ��}��)�ꙉ8NV�3wp��5�t�LV2��˹x��^^�L�$k�nڔ�Yo3^HYp�n`:����Q�;pf�opB�ʙF�Aj�3Bvv�r�b{vՖɇf��kUfA��")Ͳ�5n�:n�GA�P�'Y9t��O�eL0I,mj,�oM��l�(�Ê�� ���Z%ӵ>k#J軫[j��:�O���Qi�®$7�R�у6==Ne��&s�X��ô~�WEg�;�}M-�Aɘ��ꉉ:609ڐ��M_.[;߮Z�թe˛�<��z�#���+Oٙt�y^1�^���T`�	���Z7���jӮ�y[]{��b��0!L�
�j�6m�`*�;�̑�Ey*XX�fYDY�X�ʲ`�Di3��������m:��Q$�&��$Y���7&<��mk���]��C�N�ow.��5�=��[io@}&�ln���b$r�!+)�2�X��h�:P�+�g)e��N7IX�Z�C���\��
ʍu��,ZG/�XZ cfR�'�Vi�j�(Y���A���~e�Ҥ��|��T�qA�T���-�s�r�k��xݰQ]se���U�M��1MЅ�[���,Y��#c�5v��"m�z6*ڔe�iv�txo`�����-	A��w�6H���i3r�m��X��H���1�'��G�$z�v�̬GT�72�jN�q�[z���7+i)���ɫ�e�Id�*�Xf֩nф#�V�w�ɟ]�&+�&���JY�%K(
z1�g��	(�7A^b�T�&\��`XTBV����̰�J�L,�ݽa��b�A�&���Vn�ڞB�\���sec�݄��d٩s,Je�B�}�F'���<+�H�>zwD�n��/�݁�΂�Ƀ%A�m3�md{Y%���M��d����A�
��Y}�&���X�ؚȆ��b�-��e���FmCY��1�w���R����2�5VaȰ�z����sD;��3���EP�tE[�Wqf�mL�����r�N���MD�#7K�(�P�Q;�M  ���wE�N���f�)lu�t��7����go
Xt)6���Le ��[�\+�_��.Z�a�c���X�;bܶ�T��۱�����n��]���6����ĸ҅`����;���{ �U�l֊�
y��6�!�����g��.=je��GQi�]�ӡ@�4ȸ��]ꅯ��LU�oS�z�vcN���h喫m'h f�q��WH�tb�[ۂYsA%3�H���ͦ7Zw�b6���!�PJ��hW�
�{��'�))�b40Ѡ`(6*�mökFK��&ۛi�m37%���D/���\8�Ah��xtn�h-'q!ۣuղl�ݎL}�*��SWD���A5l��@�b0�M��VFN^х=[Y[�)�&�f�*�՘9��v��o!�����4Q���o^�LV���t3&ڙ��+5F�,�Eҵ�k�nK!����X��h��pL�e�w���m]ൣ�+�n�h�c�������eu��H�Y.���d�HX`���極,����V f&&��hWtL�^ȇ��bъ�j�n�/oe%V�kX�mI&z��l����@� �Z��l����+f��y>�4.��q<A�(ne�v��ͽK�.᫷�����^�Y�\�����?�R�jHw-\��J��:6���A�8�d�OE*Ԫ@*�US��0 W*�T�����т�]�J��!oPeLe����U�tlQu1�R��1�uCu��q�w\F���gEYNz�U[�J�QU@UUmm+��UU�h�y��'�����'kRsg�S��:����d��α���l�P�^�;�pu�����M˨���N��ޞ�79����h�k��cE��3=/=xoi�v �_:�5����g�4D��ϱ�s�V�۟;�(^ݿ6�Ϩ��ܭ�����AhY�ɺ�n�-ޅ���[�=�1sÃ=�����[k��Eӓ��'sÚ]��b�%R(�T�$��cy�aqH��u��nڱ�u۰@�7"��p��=8η�ܚӬ����������c\hZ�f��ܸ�r:6\�q�Wayv{��Ձ�n4+nnrr�;��l�v@ӽ�'����X{8x�NR�Gvۍ����֬�n�zH�ڷL67���]�<2s�m���]�����/mۚ�m�W)Q��[���%v����M�4e�r�[qf9���;�.���Eݣr��+�d�&�}���KeD����ƫ8v�+���oqn��kܼO{��[N¯]s�ً.,�n�;Z}Xܨ����ݮ�k;s�Մ��Y�n��'rN��W�����[;�������۞�S�^�|��0�j_e��y�k���v=+��2��N���c�z�v��m=K��،���98�d�\�+��՗�݇�Y	�f6m�����lcw8����ڃOd��=u�׶���1���LtZ��s��<�<��u����9$��nN�<�۳\�]�gC����`��݄N���q�ǵY�v+��ۜnwF���c�z݇�Y�n�q��À���.8��[��l�b�����m������� �Gmڗf����2h�6蝵�5�y����Vl�ۛ�� Br��rs���]��r��������R0v�s��Pkph���x�^���^��θ�M���<ہƷA�f�Zջq��t��s��ל��Gd#��z�s�[�y��9"�X;5m���q�K���.��[����GG9�&r��oG��l�m�k7�@K�k�g��ۤ�m�A��g��Nz�A���U�ݙ'�8.C��m;��e�r�n�9!<�Y��۬���d�6���r�O�s����8:���r�xK�[;��Z�n��r���8��{n3�����kn�nx��7���#�Cѳۅ0��	n�8�ƀ��.���*����p�i��Mm�ڷn��s{;�x���࣠mgv�.��A�li�x��Ӻ���z�F�s�����^�:�^��i�դ1��s�ly
�;\�t�&�jݷ^����l�vP1u6y�m�Hc�k�ݫ�t��ź�����.ؙ���\M�>{u�hsɤS��t�ra*Bfn�kh+ax�U��������iz+b^����J�ݎ�s��v�90�tG6�b�/X-���q��1��ڻn
b�G)n��*��F	��{��>^��.�� g��1e;���5�9�y��y-շYɞݳ�w]�%�`��\@6�;�ˀ(��pō��p��;x�X1�=ml�]\X4v{�6�m�u��U���� ����f�Ü[qj���)ٍ�1�=s�S��퇁�d� vN�x�Zw���nr;K���m�[s\]mtl�03z�=N�39��Ln�E��7k/A��۞�u�n��a�<	=�nv�����N��A��ӈ�8]���{r��n�7[w/bx�s�O[���8ym�2��F���8q���3ݞd�k��v�󵫂����O������3��xT�]N��8+m�X*�U4ժ���Z��]�v��8ݪngir�^��I�=��/s��pgp�z�@.�c�t�k2&�u�=pS�/��`�صՠ�+��-�ϸ�W��ɘ�˗g��q�0[k�v�u�꛱\S��T=���2�@���]f8Ҁ����3lw<��;�/c���r�rr��Ӵ>݃�<�ݶ�V���8�Zvέ�vK�o<ү����7@z�����;���'E�.����m����\��n�f�ڰ��e�	���\mt;��/h���63��=B����;��]��n�zĶ�gev��;fs��������s�P�ܱ����g��NW�k�'bܼ�7L��4���kw<�gb݋�V�Dv�{]#�9z-�vg�;�;wQ�l.���p�wd����G\$ki�nw�ݑ6��0����7��[�r�u���gp�����ٞ��|��m�;�ɣB���c��v�e���[d搊;S{;��^�UP"<��{{3	Jp�Dk�(�;�m�����̖s���v�=��7/����%��!�;��v;�����x�6�]�cn4�X8�G=z���˱�i��{u�4�Sb��JZ󝝑�nѭ���WE�xۃ01k2,�tUݱ�/.F�\�G=�7lǨg��<�a4��ң�Xs���.Ͷ��'^���y8��V�cB��۔::ִ,���*-�{s(dn{f���?@�o���'N����z�\<FN��S%ͯ"��we��s��v1v���[�����{xxz��'k]��`�;3ɷj�UE������۬�!��������*YŵӬ[>]��.m��v��l��{���}���ܗ�ד��nZw��Ӎ��6�n8ӳ���ȉ��K����S���~�}���d2�H ��Ŭ`�-����8x��yg7g��x8�c���;{m#U	�%�cMY1�dN8��e|`��� pG$�	U �3�I8�z#z�Su��<��W]{%{O�[u��X�s��˴��v�{dGUb���m�H*+�gٕ�nݩ���سt9�
�._\GB� Üv�v�k��!]Z�m�y���S�"G���o�;��n]�ӷS�y��m��vv��~�۵� :��u� o<���Ǯ���2W�"+vR�AR�c�B��b'n�h��u�۹����[N-�6�ӓW�{[U��C�9hˎ��clk<6��`B{��\p=f�����v�+=x�x,�u6�9:9*��r-��mj��Ol�˽�����F��ݞdu�>�7,��M��ѫnx`D��������Ů|�޸W!��E���v����q�)S�<�^˃j��s���w=��;�L�8�B�v��ݞ���D	�F�N��uPn}hM99ܦ��l[z0p�5�ғ�2=�[Ֆ�3��j퓌Qv:fR��-Jmt���]Ƴ��f;�1�:I;�m��t�A��:C����u�^��Z5r�ӏ����������l��/v��r�m��;wMlm��gL�;X��j���;��Ԃ!�aӉ�M��ãFn�X.ziܨ۪�P��5ù�ˍծt�1��!E�89� ���R4���8��U��˒�7Sm�A�85Sq�wn�G͢8�r��E1
Y|D:���
�Mq�bB۶�� �������[u��]�����㖹�m<n�9�O4��rng����u��=z��3�t#f6�Ma%�c�O6HJ,>{B��8�z,�9M9��\��F(c���_cv�����ɔK8�'^=�<�N������ہ,]��s�3�ܮ{�l]��j���nC�]9�n��>�O]k�6�t���q9�gn�7v��x%㎻X9��<�lI���l�ťk����Y�֮8�%�������s�9��x�Q��s۝�/G\�z��N�1��t9�[�Iۑ�O^Ǟ�������\�Ϝ�x������q�:��t���e���������Έ��+t���N�������胡n�a��ۋ�5�d��c��zVy#�rs+�i�:��m���pt��G�k^u�n<l�FOspe�k��uYy���aoX�;��k'1b$1fșf}�1Ĉ�pg`Ť9�g�vpY���<�.�h �z8��n �
mt�5[/&:�/ۅ�x7^�㬎��7�s�W)���3u�a�;C���u��8*om�}��m�ɬGg�w␺p�:�Ll0e��Y0�ݩu�5�Љ���w���;�u�w7K�e�����ղ�h��u���vv�ہ2@'=c&��">n�oR�wS��6�)�e�Ǧ�k�lC�VgJ���:��BG#�R�e�Evݼ���ݘ[���Nջec;OT\�ޭ�W�s�M%����&��u�͂��"N��gY�=G�n׎��k�s�7mf�O���l�9��U�nw��X-6,��9���e���#o��Ź]�'�<]���V��d�ݎ���.ݲ��9��q��^-ß4x�3v	�y��GB�<���.�u�������������;V9�s�$c���\��{Uv���sӺ��a0������������x��2ܯ��;A�8��;ù�'D�����j�+]�Ń8�I�19!���=�a��Iv�ۓ��7\	��<m��;u������z��9���6r��Ŏ�z:'�5�hݘ �����g����f����hr%Wn�1<3�f���},�tmy���.r��ůX�0=���g���a7c<��3�3�-�rmã~�@� �c��}�/X�tu��øݸ�;Uv�m��vN5v�����q��n3k��tn�m]/�mv������g��ϝn{I�;������zԋ��z� t�¸�=�PC������������c�}�	�ݛ��n�Fe��n�/K��k�{nπ}�X1��v��f���j�m3{v��7+�q�՘���Ԃ����L��uu��]��d�z�]��#��G@��N3�mǶoa:%c<��a�ݻmd�G]͇Fmm���/n ��y��|��U��!�O�[$v�����[��^�9��ڷ67k*>+��:.����Dј�����"U�81����i�n�8����\�W'kB�9%�����J���h����!!!!���BH,�$� 	$	#	,$��������)[jPN9k�cu�N\']g5T�Ig��.a��ɕ������{	��;Օ�g���ہp^.�1�q�>�z�X�m��݌���˝٣���gu��i�+��g2��W)�]�JVe�rf,j��q��{m�ճrI�g�<tq'�a��Q��7b�����g�c��^�<1m烎Ѧ���1ӻv����g������,�C��N�ݮwK�%��v�\��)+�Cm�v���on�ڹ��'J��9{r�V9n�x�wVq�'[���;v�ۙu�ݫn7c���na�vòrl����<l`��ֻp데n�d����t�s�n��sF�R;l
V�{Zғ��H�ggwƢ��d咮On�1�M]�#;�9�ۗ�����wn�f6�8�]����z�f�lc�t:���-nڐMt�3����iջXG���<g�r&�m�ɋ�5���V�NL]��,��R�v�{f��Yq8n�q��amv�8�c�n��å0�W;z�׎x�h�ŝ;��f���-�0�-���<vW�-�����m�t"��.*�8N��nݗݲ;7m��t�i/([� ��ɹq�F���[�\��v�w�5����[���c��XG'l��zF�\u����j�O'�n��;�0Ŏۘ�9�SG�yb��6ѭ��v�cK���\J����ѐK��^�<�s�6����QI�ѹ���=s���Y�ݽ�m�5�rl���s��i�D>����&��D{��5��g:؎Z�1%��ڄ��z�벆�nc�#��Mk3��]�yc���ڛ�Ak�A]q�6����]��g�n;�q�7�@�dzi�^݌۲�V�n[�\�qTN��c�m���7cn���/'x�����e��N�'�Uu9��˳��cnr�v�y���7<��,���k-��<�6ۣ�82=F8�^�4��Q�{uK=���@Nt��;u�A얁7&��D	x4�{�$��� `@�	 Y	"�!"��`BX"�;�������>_�;a�{n��M���<tgv
L���X��N�����5�x�k ����*v����u�]���6�a�׵�q��n��wF3v�&�ȂL��3N��C�s\��v�q���0��=�<�a�p<:�[o\u�d��� �����Aͳ[m�6��u�6��;Ƈ{/h�q����;�<���.|��ng7!354=�f�{��k���v����ln^E�`��7*���.�ɸ�n@��)���!X�Q0�Co$c:]R$��]����p� �~b�X6Ϸئ�}ͼOS�͇������&Kf7h�o8�����އ¹=�f�`�~�"<;&E������u�o1�iCޒ�����P\����5�k4Xt)��M�~�=�Žz�����K<������N�~g���g0.���R<Z'VoJ�0Qȋhg�.s\���	/3¦���Sir)_��j����{=��g�G�k�%�����l�����br��}5�L�ڡh��&PԽ�1���o�C��޺3��#N�&2���$F�x�-�B�^��U��'�br̹k����cC�Wl��^�V����Y�A����n!}�tF��d���Z^ʖx�C���j(��A�0�N;@�]�;`k=��R�m�ď�l���T����W{d:��bKK���S���V�Jψ�`��7xUP�B��_}�L�7tF��̸i��S{.e9��YyW��Jd��p�����誈�vyOfJW�o�z�,"i����4����P�]J�~����ց�^�{�l�<���u����!�4����N�a>]i
O����;ϯD�����������<f����?��T�৔�<���ǆ����fv֛����C�MNe�>n��0����0)�L�H�f���o^�uｚ�Ov�0�e��ﰙ���M��a���>�$r�KFs�}���m|�����3[�?=|�Z�������s�T��7S�4�)�B��v~ͧ�P�·�j��Oư|Fl���i9�&�'�˚a�]{f��x�by�P��}��co9F0�<��_ܿ��7�����_8ɬ���>@���%����}�f�3��y�Y��)B%ƺ��3�T�j����40�V"��tLa��6~k�k���L���!Ͼ9Y�}w�ޠ(��$F�W���1�f�}�]�Mz[����x@���-L��m�}�,5�[�c�b��68��u�s˷l�EmRUJ�*#��iq����V��X(k�㝭_�P����ُ�/R�̼S�a:)�#��S�g���\����w|�2���V�u
����Y�}zK����Xt�P�uO�ڕ����e��m��d��l��/���z��߯�"QK�E^_c´1�h"��t��]_}���pChy�bb��\�����S��a�����+�ϪR|��1�gj�u���:~�c��ub���ԕ��t�ylƯ+p;�Y���)1X�>�l�O��8��Y����^�x�g�PI���z�C�kk<����J����}f ���\ʳ}KuU��y�]�;4��>ۖ��"�ż��)����-Qy7ۯ�}��@�y���G��Y�)�[��}������Y�<�W�
a���Oj�,j�(�*�,�g��a��3D�=\Up����7U���ѡ���U)�����q��`q��s�Ϫv�ڽWi���������㣽*WE~B��
�|���M�*��Қ�y+��eQ�Y�����wtu��̩�_<�u���+2����M�}`��0'�m�W���$���f8����:�ٴ�Ne@��~�w4i��}������/v{�9�����UB��HAI]���fxώy�r�;�c��kp\zv�۷\9{jM�
E��K��RC�9�I2���ę[��q��LN&��\��ET<����Nv�+=��R{O���V���T�>B�]W�o��Y�N��a���-��&��ww�V�|�"$e.�ƾ�����|���K�pvET[�Yɏ�־��	�O������נ�yD�|��a�_���8�Ul�(6��]6�^��G2�!�q���{դn�����~獽�?��\���fF� �*�o�_��4�������zO�q������Wٗ��0�4o1����뿽����%���ϛKv�7��:x�^�m�����=��N0��%u6��L�)�L}����	Ut\k�hs�Ӽ�hr�ӣ��i-��������Q<��N�s��|�6��6��U`�B�y�j>̄h3��JN�Բ�[F�yY6,{��Y��i�6���әpf��GK���{�h��W�ض�5�ڲs�2������J� |����m/4?���u�.��k�� ��wu*��b~������U9�>��p����}d���J|�KC�q����n�Sڠ<��N>M<�nv�I��:��٦y�s���56VИ+�T���vW�L��l�e�r%���y	��\tm��Ғ'*Mwm5�n�ov��{U'�!i�ɦ�M%}T�gz���=�֫P��,��4ϝ:f�k޸|�g���[�b�l��2�+:̽�y�Z��~H�w\�9Tc+�t/ѺŤ�.�(��m:0�*i����^���"\I����R�
��|��J�o�}��-��� ����d�4����h,Co���v�!�^���N�����&ݳ�n���Y��f�8��ۼ���bLa ϖ�B��x����Hw��nk6%0/_k&�^U'u��z�N�EQS��ڲ�3V��];7[t�+�]�2O0�:��w{㲲���z��u��wk�k�����R��=���9�4�^��wZ'۟kz�VͰ)��㤤�9�`b{\��T����9ޕ*�}^�4��}��.Y�X��-�6�j�ڕ���Vm]�a��߽Ou$�lIgu>o�<c��5�׈|8�[����M�n���q=��u��>��u���Z��o�&��Ė=�q�����_�ުI�-�I^�:I\����U��
�֊��P|'
<E�d�Ź��<nK=�gel�5����0ڎ�����q��(��:�Sn��\�B�+D��ͻ� #=a��Hp�I�y��qn�M�j��0�yWh�n���s�#��.7��nwQ
lz�wn�]����u�b��ng�n���UzN=7O=kEa�n��t�'Z����7[���\7go/��{.w"�n:�9☮�m����8,p���V�n��^��8�{	�p\<u�P����dr�9�8�ݢ��f��C��l�si�!�ڢ�s���!���r�A����}��ǈ��R붎�^ݭ��M���YZc�����	�U�������x�0��j�y�h1&5���وR:��8���R�~���U����O��:������*�L�>yU�q�o[�C0��Lʞ�qt��}��:�2��Pe���m���F�"�m��k����V�5��ƹ��J}7� V���DR,7T[�jÿVs�yyS��fP,)&�����|okU�޻��d�u�S��]U�)�UyiM�0_�Sכ�4�3{��{�߫S��Zy�H����5P.�/�ov.�Sl�������%?}GY�~A���|��fӉ7�7���ϳG��v��ƚr����q8���+מ��k]��o�S�w�YW�<�m��r��Ӿ��#7�o����m��m�a���V=�_R��/M!�(j�b�X��u2ec���E�<�d�n��*�FO�I��9���X�C�U0s/0�f��q1��I�4�:s5��7�&���������w���٩O;�Nn��n�V�1�,�}�j��:�j��[n�x}N�w������Y8y�q�\r���{�[5%��-�I�m3����o!ٸ�z^���L��3٩�|-�
c���4��]Q��~�i�{~I���U��f���Rߓ�P|��8���r�=h՝�����|���S
������ݾ1�g�����pLC�3��ح���	�@o������8�H[�&���������Oy����@��W�f{�:\�{�:KN��΋������P��[��F�в$�	:q_I����76@z��-�?ga��_��Re��8��I>v�VT7u:��s��jÌ�q�&�Za��zg�O}E{�����﮻��e�l�n��i�-؆�)3��ssD�KMq��&4�s��i�}�$ĭQ���7iUz��8,U�����ɭ��eP~"
��*�������gu�y����h5~���˖�bÈu3(�w�����{�鶯,����� �緵5澮>'��?^�3�G���,�u���?{�;�.q���7@VRϳ=���ԘͲr���bf��u�u���ﹼ�u�z�O����Qr��<�'�"��"�+vP�]QoU�n��^�N;k=`���8鯛\��Q�\v��v|�sCY��P�Je&�w+��3l�+�傍U<g��j�5A�&{Z�h���m���AV��u�W�Z'�b��r����v�r\h}<&�;�"�Dq��E#����V5O2)*���D)JE�ߚ�IW־*�ׯF�s�5�
i<�'7�d���6�����Ch{=g7G�u����y޶s�lܜu�l�v��V�F���O�v��%iG�r|��qNq�+r�E\�/&�)L14���5\�랺�����y�l��5���u-����ՠ�v�Í=a���'
����]޵�L|�q���H�_]ۜ�a��M1^N�^��iW�\hk�ٺ�IU����:P_c4�f�Ҳ���Xq�{��Xn��u�|�TJi�{(�f�a��]�9�O�{C����/M�SI�KN�� ��"���.YF��l�����ԬYniT��7����jkw�����B���hw�mznQ�M �S�U^W�z8�x2c�b�+o[~O��nq-�Z(�m��h8�MU��5�]-�-�^^�f���iNQ��u����P�4����q������ׯ*(b]߾�M��c=ϬB�;�l�6�i����[��N��?���^�t���
���^cI�k�k�s���X���7iAW����$>5�Ι��{�l>IO���}�t�5��n�^�,<�3H|�W�>����z�|�&>�`�ZN�f��d�k�1�D�&�+���_/1ﴱ����r�Iaݳ�s��'���͹�p�u^��+{v��s�<x=Jp���2� ��%]N'���'j��N�\waN��}����'Ϯ�Ő}=��
��c���\?W��a�N�>^|^u�B�O2��5�^�E�Щ�����q슿����J(�b
V�Y8��U�
a�ڶ���k��|^�?!�����:�eN3���0�u�+��M1�u��lB���&�^��0ޫ��2[+��Y�ot�%��>c��ة*:��P �^"���_m�Z]�y�5d�)�u�L�1oZ��M�<W�f��7�n�����u�n���!�i
i7��ՠ�=�{4S&��!�/����_V�4����Q#�I�8ǽn��;��{���V�e2귮��^��ow�ۮP{��Nj�<��-��*����ǌ���'��n�v��B�~`z������Y8�e�կ�7d1���$>
�Wx�;L��Dhܤ�s�R���9|���lX��X��If��Ee=�eL;��lZ��[5\d����U92�**����)�l�k�v$4���>�.��)�9����\������n|�T����@n�����ü���2�86�����WjC�n�Hw��۪���A�)�~k�iP�)�u��.�0���T�ײ�ݝ�6\�Z;^��݉1����s���Q���������o��������{��Zq�3K�@�?W�R����ޤ�xf$2�Ϸ������Ek+�f�l�s�i'ɤ>�Y���� m�4���Ggޓ-s���A)�y����.��.�<o�dCM�wU�{���绣̬*t|�c'�[��4�h���v�QOk�ތq�k�Q�w��O�JM���_��/2��/2򧒝�Jd���T~�5�S�=t���ӈ}�o&���m;��:p�k_����sf�;U�ѥ|�/��F�o���c8�Oz�O�r��t�X{R؝V�D�U�}��/�|>s�z��Z�︗-�|�j�vu'�{��՘�Lw�on���q�ͳl6�T۴�x,�}g��:>�T��!�����=�:���?^�B�������QЕH����9��h~� ҉�yr|��B���n��GP�u_��a�);�o�zus}�r����O���6�N���A���u��m�xkI�U�	~_9���W��*���^�PS=�Y�*�lz(�=�Yy����	�M�uc�mû75ۖݡwdя=���T��Aq�gA��QM�ݳq\Y�5���BI-�B�O�5��^;����Ѹ��Gl�ۭ˶7L�.�R�����#�kv!��a������o>G�c�,��ׇ�ɬ\��\܆��O�v�����s��=���ݜ�������Op���w��jSυ�N�����;j�lm�3`y��6z��1�����uP��8��8Ţڰb�Z�������mf��Ȯa���WT�܊��"ɢ68��jv�9����2���Þ��Nv����l༝z��e�y��A~B��?~��5�Y;�����\�O�޿�5p�t�ʚ��4uU���߮|���e�׼ʟ0P��*��g���
j��9G��Ѧ3�pq��j}y�L��2qv��J!�����0J��T��zi��[�X�UF��{(�f��-�e�Sl%'־٠�T��2ý��M;C�[sw���1��z���M-p���Z���,��}��H5ƾc��X�ق�C��O�P����^Cl�q�7�\�����8cm��1�5̚NU�r��%eM6ɫ�t�7u�P5u�S����9���uK@�J�k��Iy���L(�_��P�{��TJ��em��{�o��i��H,�C��~�x�Li]'�9��>;νr���q���M��GyA���w﯌6�y����^L��o+1֒ue�Դ�ӝV�,T��ULob���w�i����8�>��bu%��-��������4�*��e����@S=���$ἵ������5�R(� ��7$A�tq�w��gn&��n�'���gn��.��b���g_��sڍ*��}~K3��Ͻz8��l��O&�[�<j�~�':�8�N��6�g���=�7����k]+�������u�uu�r��k�o�ƾ�.>r|�����*����sh���д�i�}d���k�Ͻ�>J��fZ�����%[�el�:�*^�8���^�ym�Y�K70�R:�7yD5��7ը/^�j�g��H1j����i9�n��Rc�����f��L�|�L:�޳�V�u��S�r�O�=�)��_xS����V�B~�V�c�rG��k�2*9h�m
���_��cCB�����_���Z�i�����RS=�^$���{��z���=es��]��2�-4�5�>���M%%򡉦�hd/�o�[��_���D(6�P�˳Zs\���VÕ������M�yGy,�M긇�VN���}�%�d�[��oqӶ�|��{�Q�V��湛����ٳl�o�p�>�ÿj�Wl�(���̸�i�.��z��5��a�6�eC�vי�����k��<׮u��]g���i5�)<�wz�h/���KK�k<�~LV^�co�Ud?i?W��b���wi��a�=�n9ՃH�.<�צ���m��:�Ёs��d���ò*�Q4T	�B|��>K��C��ch}��6�����1-1@�;z�רf��[ʐ�j��<�׼'�^��wf���(Rbk׬5z��Ӷ{E����ת�A���H)�I5_X��r�N�Io9��hRo����zx��4���'&3_}|a�T����kz��ׯV�q)!�L+��T��<���wqvu��G�4T��.Ӥj��/*��R��0�P6���)<��_��gq��z�9�ˬIT������Ga
�����CJW��Hj΄�������f;��oH3��1A��V�%�­c<��)��D5�v�%5ь4*p�����y�ȇ|�'��}�(gbo�&(I�.�g �W<:e�+�r�f�0d�[���3U��M���0��m���/��m�����%%m�)V]��Sa��![̼SM��Më��e0g��W6g��K���Y[Z�0��Sz����CVM�]-7�n�P�wD&�o�\�Ďuꃅ)�G����C����.�����yEn8Ӑ� _sG1Q�����w7qu<�;V��o�K�IꠘE-��I^ʱ��$�ܚWa�wR�j�h��rd`���;�х�sj�]'H�.����f��Z�����D]\���ܔ��:h�|���{��c-	�����'d	J_VC�vY{f�n�5�n}�E��#��4��{U_ǋ�#o��c�����9���^�=,����B�$��-�6 	��1[ ��4�)H�����Sb����&d�Ǖ�&�9Qf�/TP�W�8�W�`U�-��.V*�WK�N�\&b����fc�d��
*[q���v�
�R�E\�}�ݕy� @ɳZ�S��0���Y�k�3o��ʙ�[i�ˋvWw#9���T GL��Ӟ�+Ko�qz,*������Ҏg��^ee�ygf,YO��+����$ɓ�):ܔ�Zx�XLnz��uk�+8{��1����E��KKp�p$�ʻP��繐�v�^"�L� �b������J�דoW]�x�i�������t+���G�D�0~�:�L��� ��bs�W��³0����&�)$��$9TAH,V�
ATAH)�]H�o���p����H)�	�) � �~e0����;Z��{�I ��$c%$��ʣ�
H) ��� ���RTA~@�� �����4AH(i�e�=˹>�S�D��R
A
Aau�$�UR
AH)>B�:��
AH)��w7�
AH)���Ă0�
H) �7TC*�) � �����w��������*���R
AHe{��'���
AHr���R
AH"AH) �*���S�@ZAH"II �����v�i�.�������>JH(z薐Y4��Q)
H,� �9TAH) ��b�S��RTII ��
H_��F������RAHv����Ii � ���]}P7�AH) ��$�/]��O��
AHg3�{�RAH) � �RRAH]Q�
b=`P�R
A@������bJH) �=��th��PR)��Hr���_��R��s0��R
CUD��P?%$$��-���Rַ���)1
C�) � ��RZAH(f��� ���D��Sh�RT�S�$���o�����5����?}i���7�XV�^Mg��f]�:�eC��� $v��m�r���9�e�e��
AH)���� �:�AH"AH) �.���S�~B�TA
AH,>RC߻ߝ삐R
~@��$~�Ii �5Tq�
AH/�T
AH(JHn�<���v�X[
H}z�&�)<�!����T�gn�)�[H)J�i���i!��
AH) �s��c�$���{�V�%$���{G��ܔo:�RM$>Iˢ
AH) ��0����I� ���R罣@bRAH)!��
At����RP�R
AH)� ��n�R
A��ZAH)!��pmR�fQCv�]f� ���D��R
AHUQ ���FM����T��� �>i ���-!�O��h��Ф��R� ���;��~7e��M]@��B��J
AH)�h�O�Ru��R
AH"A`5T��) �>��{������R%��D��R
ACݢk(����aI�愂�R
AHj�:$��$�����F�) �꧘RC��As��
A� �����;ꖐRUR�R
AH)��u��)�) � ���Pu�����Q ���D�Ì)1�>JHj���R
AHn�j��ř�\�fSYyF�)$��(Hv���X�^$�') ���ʩ5���R
AH~��) ����Hw��ս�Rb�R
A=�nLH)!��
AH)�o�=\aI��� �/��i ��{�h�~II�M$M��D��Rb�D��X_�5�����a����Q ��) � ���i �?s���d��R
A
AH):�$.������ �̔�D���Q�
@�RC*�H��
H)!�_?Q�?%$�ܰĂ�Y)�tAH) ���$;TC�y�$�� ���H)H,��
Ag̚�����G,V�����p��R
AH"AH. {��y����Z�1��`�R
A9�ޯ�_>�{>��R
AHn��������ik�Ѡ��1 ��U�Q ��B��@����
H/���� �N��
A�JH) �+=����R
AO S'�P�R
AH)� ��B�
�@� �������v�%��$���u4AH)+�o��p!��-%��R
A��
AH)� ����U}^���zL����~�{�\]����XV��e*N�ҢM��@����j�ȃ���-yt�f���j!{jӘ^O��w�~of�����- ���R
C^������RO^XbII�̤�βRAH(VQ5�AH)��N��R
(
AHeT��I ����k���-�.�V`�fp��R
Ad��]R����R
�
AH]T��H)�

ACi) ��B��w��_8AH) ���ꤴ���RM �R
R ~Jw��i��) �5TCuAĔ��!�Y�����������RC�����=��&�$;ʒM2J��נ��)�%�
d��!�	hWh�^� �����̄7�-�II 9�ۦ�F��x�Y��h����a��=�1����L��&�Z���˻�Ɗհ���m� k�4�K�)? ~� ���U �7TAH,4�2}��Xc
z�����P|��
Aa���)�}�D��R޲ZC�P��1�\��]0)II ��큫����ͲRAC�)��U��������AH(i%$M�jZAH,�$:��D��l) ���R
��T�Y1 �aI淽삐R~B��O~�vwv�Zu�D��R
AHj���R
B�) �W�- ���R1�����)7���%$��R�V��R��*���X[
m�I ���Xy��Xi ��w���maK�]V]fa�
AH)!��
Az���R
AH) �.�E�AH) ����S�RC����s���R&�L>aL�|�VII �9TA@�RAg)���R
AH)U[@�� ��9����:��R
Ad��ܢL
H)$����U0�~d�����) ���R�I �7�on�AH)1]� ���R
CUD��R�$��P<���j�8��0������F�.�wگ?���AH)� �L
H(x��OW��N���R
C�D���R
AH) �=���ae%�h�,������
AH) �{�%�1�����
Aa��R&UE ���ʢ
AH,=����k��&Ф��@�Kgn�,�%'�
H)? RAe�RA~�p;� ���2q��R
��r肐Y�'��=\�JH) ���^0) �2���Xk����}�o�ߡi�M$��R
�}tIL
i �����t�$��]��@z���D��R
AH}TAH)!uD��@��H(RJH) �/\����)>���i�RCۻ�̤��R
AH}TAH) �m��Xu�&�)��� ����aI��/��K33*ܬ��R
AL@��*�)��U���R
AgY)���ԛ�e�����z��w�Ă�R
A0) ��RC���� ����) ����I!��
�N��T`) �.���ʠ����I �7����
)�֙)���Q ������Rn�i!���B�
��
��
AH)k�V�AH)!�
AH,
i �.���R
A`cL��H)�~��}���k�I�R
Aal)!]�����3��$����Q�d���P�h���TJB�?n��`r�N2�
~@���R
AH)�]}�m>�ΒѰQʨ@]�K�F�����
AH,�� �5TAH)!�
AH)�TAH,�r�����2�������
M�����Q��\��Rm
H) ����肐R
AH)�ϹU]�ﵟk�ZAH)�7�{ ����R�) ����II��
Aa���R
AH) �5T��`S%2�
C|��h��P���h�l�� ���RRC�vAH)!UD��j��ۢ�
AH) ��N����d��H) ���R
{vG(��R4�I ���RTAH) �:��_1�cIX�x��Y��Ppב��t��
�P�)�>�W��6w��w^���$�ʇ��k n�k�o�!zV��%��e��T��>�_F�m�:l��P�l�vcv6��1������J�mv����,nk`�;�h�9�q���{9���\q�\3<V�
w>*���	�mpݎ����]�-��I\��R��pR��ܼ��g�v��E�c�[Z�v�f�!�ݼ�r�V�6�Z��Z��q���m�y^�юN�A�#�WkS�A�����\��1�.�띂�ֳnxySQ��h�<n9u��U��2g����s����fQ���R
y�� ��J`[I � ���`]ԛ��R
R$�$d���ʅ;`s���{�
AH,�e	�"�����B�RCuF z肐R__pld�)�XRC*���������������ϙ;��٢
AI�) ��ԫ��r�TO�~�=Clߨ7��ۮ��|��u��$�>�=�]!�z��K��N�E��s�}��$�zM'�%�V[i4q�=M<HSl�ϊ޲v�go�(��3mr�)絭:��>����ǯ�(�����_n�=�w11��[�'v��ʐ�s�ٳ��E|Q�����P�ʣ�s��U�%���ʬ�'M�q9�6����=�R�y�(4�v����kÑX~�H[8��᫾j$�u�q��yg�W����g�S�{ʁ���Pj��jeT�1-�f�F�i�+��^�j���[\v�[�_wqc����[/}����_5G���o[�A|�;�Y�P��ys�|���4���i�W�]=A���.µ��;���Se�s���x��;����ٸ%X��)��;�[�mn�j�eX�tn��K�f��2���j����b�j�믻�r�,��Mqt�N�9_f�vq�4�3�[����e+ԜLR�<�gݭ3ɽn���IN���^�~�'����}�r��܍�Tl��ʭ�i�8��$������F1g��Ў\����vjo�nm��!���'.���Ͻ{�i�-�ھ'P��}s���ur���4��R��l�׵D�}�Ν��>�G��}Ahb2�{�:5tB�y��զ+�ן]�f��/(��ˏ�UM���X�?���k�ھ�7�a��L�<n�a��j7rx_\�=;w��tvC/�;���85�Úf$u�����
g
�P����1W�ɧ٪��t������4����H���Ҧ��v��H[*���r�R?}r9[@Ӽ��i>�����fh��o~y�w*�}�>D�N�nr��ƉX�!m�ruz���O���:�zϽGS�P�)��n������ܱ����y�駧ٶ�}��@��w��P�io���h6�1�'��j�^��4�q�a���)��ꆖ��5tV)u���[f�y5�i����<�X{�:����Fߐ*�y:��ڣL��[��ђ�����|���Ow7�F!�ɍ?$��~�}�so�mO"���|���&3���c^�4kϳn+�%M[P��y��O���&��)���!牿�p2��C�[=��	⭤.���5�s��k4F�����;�3y}a���w�ƽ���j�ǡ�#ER�U��Y��Y,+ɡ�;����i�YY�+Ek��:V�4C��j��^9�0�֫�l[�G�<D��E�fAx�O'SC��t��~�oRu��LCJL���o��}��&eL��i��{zm���Ǚts|��I�uo��޲�Pě��qX��k��5�_2�)���ǐ�Ja�ʩ�I[�6q���{`Wzk�/�u]�|kYL�2���^ឩJ��,����s���'{�sΘm'��o��|��~�o���h}��R��#�U��I�!�wY��q��J}t|�����뵠Ӷp�[n��4�1��ه��[�<�I.���Z5%��SY�����ej*��k8]�F���q���G8n�z9��@����׻W/��e*��2�j�7G��{�f�4�:t�6�i����
�Y�����ۼ�l�_^RZA#A6�`���#�
�Fyo�g����u���B�J}�!�r�oUs\ɞ�t��L-���w�`Zw��!L�u�i���w�W9)^���Z!���7U���URە�WVᗙ8ͳ2W+mJ�a���@]���C�ǀ���w�f{#$�}$���z	uUvN����Y�^����DM?r�C��pb�w	��m�/Tc}W��{�.�6��� �����
HA�-z�yS�]t'n�Y�^M٤��${+Ìc�V��L�+W�}k�4��>��/�]V�ٯd���3�Fi�8��}�ϯF<i�Rm4�u������Շ���y�kSۻ�����ě˳��!3�֍C^�O#$u���Ʊ����d��H��*���oɺ��)�v�`�}^w���gh�]��N�ju�IhZ]5;���ȷʒ�O�j��!���:6�ϐ�3��Z>�`�q�~�~#��YЫ[W�F�k������+�<��%�(��$X�cI{N!����q*ҙo�6%��q=�QO!�Q�i��nW��:��{�!/��+-ʪb��h������>��l~���S1
��/G4j発5�����P��B�0|S$:���'�1��֫޳oݫm��`y;��3B�o̷l�դ֨�5�{3�4���jC��������=Z�c-�>�K��^ ��Q]5ޜ8�s��LW�W@Zt߶g��i#�ܔO��3u~�����Sw���2:�[���r��]
V�W���%�*_#����JGº�g��W���oܩ��|_e�Ֆ��*�F��6�]���m<��/�������Ԫ�񘪪ɿg������J���j�;f��5ut�����!��3�bu������F�|��5��Rz��|�\Y���w��ژBYZ��8�3��n��O$����\���'G,\b;v���G��_i��I������P���Kx���r�f���D�T�'����,�-s󖪇�ל������𽥕6�V�n╕�ԚCWF>�RS���}�i5�)1-��ٴ�u>C��C�s{�[����y�Y��I�b�9����{u:�Kt�!j��\�Jf��(��|�3�W��և���L��� �ڔ���UR�1^Wi�e���%V`�����5���G��ף��9[�ӈq�3l�z��%Lo%��h�\�.^�K7T�e;��d��q�j({U�j�����ݮ��}�<�;O"�M �u�\}|~Z��u����L�̭��i�
v�٣���������9����g�u-���d��V�:.���<Pi6��:���{Z��aֽqh���ܯ��r�������J����컺��^�Xz�ӾU�j5M6����I�;���3MAz~� �~�b�{s�Z�ۉm��\�lG��ȼa����d��Y���<����$�}F0�f�iNe��IL{P�c�s�[�{9�1��IK�t���E�j~~Ύ,��:��3P�3Ew\�F�:�Ə]ӹ�t��q�ڤ�a�Q��9so[3[р��SO)��_�i���	>4�Av�/:���qbwk��;Olcu�헖3S6�M�H:��L�q<�W&Ґƣ62l���ʮEx�o!���������v� ��T����Cz���{�Ս"��C���w�x�Mӻf�e8{u'�8v�ۻ&�v�S�[*<�^�o\��<���� F�Uŝ��9�M7T�Ѫ�s�ٺ:�l�kRC`���qvDκÀ�*��܋q��q����x�W��=��0�4�w�;�����n�O���w~~紆~����q��[��j���iI=�Vn��|Qb���p�wd�pB�Zv�h��C�"{�)+�ȥ��>�b3����~�^���w��m��YE3u�)t^eV]�cUy��t��oZ�I�:�s~�e ���Կ��l{��r�f�Bq�-����8�����{�<�ݻ�/y����)膐����'r����f�}¾u���xO�_�p�!��O�x��R�e���<r��(�Ty>i9�!�]�򡏹G����Ն0���\]T��N�;��}��u[�|�c��ݳ��a�2|�]%��pƟ���:6�ˠ�	l>�e&��$TD������k���z���9*w,Uh��*L�����6�5�Y�PS󈡿kXc)�՝d�Z������5��C���y"���_/��q5�)�r�)�i���M]},K[kwK�P��P�~�.�[a��������M��
@�����3�u�=�X��W#�����@V���ܥ�~֯�9ʶi���c/��v�fQJ�ُ�S���F�E0ٺ��y:��=rmT�I%+b�����|	Wg���k�v�[g�Hz�\�ܷm��g��9&�#��VaI���ZJj�͢�g9]���j
�Ka�Py19ڜ�o��M']�d���n���_y�AN�����.���i����/i����0���_(q�M���]�vQ�U��Ve膒�9ti1��˂���J>��4�4eg9qqX��ފX�l��nV����A���$�"����V�}���^���>]!%�H�r�W�^�7�C��vM]�G�T��LXZ'{���q9�>KL5Qq���3~���o/{���޴Y�)�ǝ�=�{U�7u������!L��o�Ʋ�䥼��'�ؓ2����g���}�6���n!m8��������8֊���麃�*�8��|5�ͳ�I/�I�su�TM��6�����6��!���
9r��8�é}����k[9G��z|����V�M���?U��v��3N�� Uטڎ3ޭ�P�!�8��x�KU�n���;�zjߙԗ�Wf�>�?4�Ś넏P�b�E�Ȣۖ�
"k+�P�u���tN����>N!����}�f���/Ri����5<�I2�}�
�{&3i�檚�!�KU���a���~� W B�h�iC�V���;.��N#�_SnmA��]x�ݱ��H�rT�؂�k��m�Ƿ�%�5�_��m��'ɮ�O0��n��Ρڢ.=E�M:f&c�d/+�t�����q��������TS�c��o��C��{kT��H��k,��F��+�({*Lb��߸l1��_/�ߍs�?Oe�m�M��|�����!�6�t�$���:�]kնN7t�&���wx�xeZ��̚Nh���w��u��}=o�{ky�w�u7��j�Z�X��"�N�H{tz��M'��)fЭQLY詺Ͼ�H)���{��E�����i\ssm�*+����n����Dw�R�B�0��gDGG)X���׹�nHYYԒ�Qk6����Ȧn���k�>���������~z���C<������O�hug��HӤ�)��G�@pby37�W�>=�{�Z_j�2U���y��@�T�T�CǷ���o-4�Ku���E���q�N�\�gɽ{�;�w���LMw����;�R�<Ii�u�h�3+�|�%=�:����5{�>��+qd�Ϭ�����S�m�t�p8�E��F!N�z��N���٧�L��գ��<��p�.�@�TP��:��<��Q���J�ch'��ql���>ȩ)�z�˅��q#���}��m���R�7��O�����i1x��Iy�z�1��w&�RJMn���0��l�q��C޾n�L���ѣ���]t�R��׶�w'_3�l�H)3�t���Ʋ�o3/PYz���je�����+�u�͇Н�^��]94]Qܜ�nz��y)-��,g�3+�\e����w��d�)�RWٛ�i۶[3��\��Y=X����j��fi��Mު�e�a5ʇ���3LS�):�$��[4��f<q����U�V���ԩb�����H!&���˔����yX�������q��RSq-?����v>q9;�4aHU �a�Js�N������|�~�g�����������.IY����>;;|���5�u��[P�~��\��Wr��H}�b��ze�|��+�+t��Y�x&i�#;�e�b��e8�&���7s}�X�3Gd�x��v��M�d�i����P����ξ��0�5R��F��u�'~�L5��.��Mƽ2�l���i�F�)�] c�UW��V�\�3L��n;�+7��R�|R��V�W�ӿ���by�L�o=���PR����E�N?a��
�9��=DV���a���?]��S&�=;�x�:}"b`�$T�ѷ]��G��cgK������e^Ⱥ1�Ks������y��d��f�P�]i	4��Q7ܖ]d�{�[_^d6γ՞�j|�g��i�t}Z �<*�_���н���`��dN��Q�wte�����auT�*JW��&�#��[Sj��~k3/�b�V}B�a��I��U_$uu�}^�;^t��bs~�C��aT��M2V�cϷ_z�_2
��r敃�{���v]�� �^k{���D�ϫ�����rzs���n�b$�F�)wƒ�bޫ�K�������9G�4�&�S�C��[�;���A��<�}��j��KKO���o!��-��׶m�~��|��s�r�gܸ����e�n�P����-T�̳�R�2�ۦLk�N�U[�u������Ij��x�L:�i�T����/�oڢ������m5e���*�z�7�!��n���ڝf0�޵e?]i��#0Mѱk
*P��^��C���l�>��N���o���/;Zx�%�dJ��sEy��W�v��Al>��`j����|�^�IN����1��tɤ�Y�z�����gܣ���Խ�����9;Pp��7��*�c�C�ݹ���ƴi����.����e�U��w���mi\�VwGj�VI��U�����7�]��K�]&��L�׀�p#���	��<2L#���K,��s*v��>B*�/+�C���1����bΙ�*R�d\����j�`�{].WR�*���^���,3��ٖ�$�G����m�&7wLс0�߇��)�ꢫJ^���򒇕`���I���cvv�g����SF���&*T]���c*:�I�*W�;�u�1��u�=��j��gv�* 8#�6���5P�������1zy-Ѵ���hPz-�-;෵nA0jc��I��q��Ό٧+��ZC���}�f�s��T����M�o���M�4��\ޡXGm3�7]K����y4�9�mt�yy{�5�Ʒ��mhV�X���-t�Nm�W�gS�\1��%���u5���
�uч)�|f�AkV�G�.�@Zѕ�.�[��r���<�VmdN�u8<?'W�u���H�~h��[{hl�D���}�����%m����дlN��*m ߴ,�8��x����fۚ��ǀ� �ق�4ƫ�؍�;"�1�u<����dP�淮��_k�c#ϟUȺ�G@�P[v���yC����/����>)�{�N^�ź82�E��;F]�te�Xñ�O��fuݵfi�fw,��7i�*I4��ɷ�R����|J㷜�!�oO�gH�dRJ���B�V��۲��c��P+�c�UWp�ݺx��9�G�۱�cg�tg9�7��]�Q��_�x��Gd���0�,r}>`����{S�W�v�ۥՖ��)����Ǧ>��Ǿ7֭��ז�۸�.��r����.��[���[�uu�v��nx����Յ<n �|���۝b4]�1��ey9c��c!͓<]��s�G�i;6�c[N��_&6cmp+�7&��96�Om����YzlF�^�x;y<�V�ޝ[�5���gy�.]�l�1��8�!n�F����5�iy}����/a�M�>CX����K�Ծܻv��U�g�g^�倻n�r�Gm����[v��8�ֲv�'v�<��tcK��u�3vr�úq����v�qgJ��B{v9*���4`/��DM�H�M5G-�ω�Iۇ�#+�k�]�[Sv���:��P�)�N]Ķ����w�7nq<��U`�t)e�E�j�]-M.��q�u�;6�۱�q�������7m��=k: ͷaL�\Юd7��^Vd��Ɛ6G�t.�k��G� ���zAݜ�˯;]Ãn����]8:.�gn:V�s���
�crWi�wc�m�d�燗ďj�Tsȫ#�+�aNl���s׶ն9n�h��v�Kmݎ�n�����ká�V,�˜t�юC����lE���1=��'q���۵�8����π��u���t��X����qx�68��<�S�[�9�֎d��w(�V�p5c����k�8�ಛ��m�����rqnk��6M��'����i����rv�uz9��d�9���{�ZC�i����{/k��ڽ�Y�rn�b�;�N��&픍p{YNvbA�v{i��\�C�d���&uqu��x�s��D4˹c�rb��̵�:G'ً#�mlV�̸I�)�pu]���j9vL]�0V�p��Ac��l�t�b;rs�۰�v�[[cZ3�,aF1�=�J��{<q�\���H�	��2����山�Q��Oh3<�N�9��G<�u���-L��(����x��֠�æO����.`m�⢟4�ۇ�
�ypN�Q������9���N�&�T���Y�����Ƶ]�3�x�f5w.�J;/X��۱B���8��n�j�]q�w`��X��v�	�P����j�\jc��V\�	N�xɉ�]��{&s=�L��mc#�%���ss�c�+l�κz:�[�Ap��{1�6��s��݅�Mf�.���Uy��>g��Oj��E��O?sn�z���P|���z��y�%z�^*Zi�M2���q�9ߊ�<�kܑ�M2}��HS�|ްҚ�i�z�˒����Q霋W\Ӟ�q��	#�	��}���ǜ�}��mnն�ԑ��
��6+��*ˬ&ǒ�T�3�\>�f�C���_lճo=�&��5�
mĴS�k�4��2�w�����^z�X��汷�����o��&��t�}�s�:6�]��)A}�N��>I����ÿQ�+����:���i���9�?Qi��{�'lP{��ꫥ��{=�;���<�9����<�N�ͤ�n��׷@�N�kTZV�=�6�_s�n�]� ��ki����8���zs�W��ﵣ��8�-����hz�f�Xϒ��ݠ=�~����ͳ�|�Xy8�&�Hm̭��[O0�-6������O���׵ύ�����>d��l4�ʊr�x��9Uei����'Y�z�&�Zg�z��1w���d��~M�'�YIWG8�¼�ȗ�z08˘ت"P�\�,��^�B��ǽ}ս��y��㜑��J�s�{~��oQD�OB���EP�u�s���{ry#j�"WprKm��r^ܮ�=g�Q��
-&g\}4nA��Z̆����>���b{��o�گE�ƞ0���V��旮ޗ�˝,���峖�Z'{}C�]�5i+��v�Σ37��!�������y}S�i^U�Kg��.:�.�JXwTްV5B*[�3�[ȋX����%eʽVA��@���ם!ׂXR�a���LP���bQn�팿>�~]�W�x�f��Fߘ2J���_�o�"ڂ�l��#q4�#��V7F�{�G�*���A1�������I	�O9��h����9��nY�-�r��T�.�y�L��@��Mܧ��]X/FT�+�f���2k�w{��7J�)k��`�8������{d��Ѹ�|1�.܂trT)hN���D������A��;�kԭ��X����V?_�y��5A
Kz��c�!̱�ݥwt��ޛ�O^�>TkJ}.�ƭ����pk�$�B�p&3�����7/=C�v��͍Ѧ��(�E���$��>�[ی[�u
�4������^����\;�ƃ���.d_+�.�/ƌ�LJ����0�)�I"Zo�y W���Y�-��4c��pe���Nw)wS����������ȇ�W�,>˂��H��g�+��mBiR$��)->�g~�Ww#<n�f j�{���A3k��'����K�UĐ3�m��ehW���Y�Xj{���l挟m:5������������A�/'Ec�*W�/�_>Go�~1qS�n��K�-�n�y���%\fW��z�캗�k�R�o7���Lz<��N�.��t���<��\���֪� ϗm�x㩀�aұ` ��r�^j8�c`�F^U�2��o^c���9ػZ��pQOf�S�I��U��^U�|�V��ՈP'm�m�!m+to��t�Ob��y�;q����wEۍ<ܫg�;�xG�� Q�������X��s{����>�G����߼W��[*n�im���OΖ 0���^�n.�ێ������*8	T�� )7ux��i��=�t�B.�|�����ѽo��W����5����4�K����|y�b��Z*L�5�<}滶!`&R����}�\���,�|�r�g2�f.ݻ<6�qyўb�xC��5t�w╙$�
�3{:���_����= �P�΁�
��>s�gZ�7;Cp:L�e5re&�R���q0}�e���q^ϗ&��⏏�֨-�ӗ ��=O:cՅb���T!�)+;�_*cCLjN�7�U���:��p���ۭԀ�fU�f�;׳=vt���-����+hdj"8������u�H���z��3W��C�cV[��u��RE���y�1�lm �]�&]��ގ8��=�r6�ntuGkU���
ㅍ�u�:@��On�����^��ۭ�y�S��7e����gܺ=���������}
�H�	�5�w�/7o!���C�u
c1c�e���y��to��\�x"��miu�' <��e5z��~�D��(�j3A�榫��)�T�Zj����<P�ދ��L�\��{Lxꢓ����HZ�e&v{�>ך���M˝�j^�y۩�hC����Rm�w-��V��*U��+k+=B�/3Jx���}l����M�(��T*�X�Q���]Wõ��!����茦t#3��a}�X��v�_01�~~�}�XS���-�'o�3���%W�Q�u1�:�rP����/5�{�o93K��Ѷ���}Y�N�o��{��f�{�Z��EA��$�`����[w�.m_xvE6��%�����7��ns+2G��c����$1�ʹ��p3�(m�J�
}�m-�|���~~���L6�[����|&�i�6W=�����W���Z9�Q�ϴ��Ә=϶�-��e;����=z[���ݻ�q����v�ϖ�c���k��&2���d�ZC�n�^�q�=���ݛ�����	�l7[���lq�{v�f�;w�n7^,d82�c��[����i�CcI˻V�����n��V@i퓖������u��g==�<�9���$]|�+�kX-��sm���.�&�n݋�ۍ�\��ݳ�3ΑI�_��ڬ��eOQ��D�Ļ��}�d͙D�e�ގp������
#.��om{����)K~��J��'H��( �m{�l�!�~�=�9�Ԭ�}����%��W�;�襟o�8g�%���n���d3*N�n���i���l�V?lv���pM��7
+������Y^%=�N��s�6ĥ^��n䱞D���_��Y~��Ԁ�S:{�u{�pn]?���O�����F��?'�Y?J�p~��Iβ�S��}3.�|�U�]Ӗ)��/zm#Ird�ۘ����[�+�a��䴮�DAD����V��腴f�qR���A���-�׳ܫ�3�<+�*�wcR�ne�M���޸��{0�$�t���w�5Ҧ��*�,�:twg��#[��#�Vi�3��Ԝ�!�'����3H*�XB!&�u].����}ݺ&yh\.ONs�P�@&�g���u�ש;�D��L|(�N�d��-J��C��Y��(�A?6�ƀ�%^a�� �ژzvZ3/l��lx�˹F�������]^q��ei����8e���5�KYvp0Vel��=/��ڄ�3S��\5N[z� q�K>�{�hm嫏�X(�����?�1�>�ϓs�q�MGjw�1m����E�@V/R9�͘�ʧ�`-2�������hئp�ݺ����&�E@Ob�,�{ݘ����V��lDy/]�{�DS�`�f�zǅ�)k��y;cs�z�m�~&�F0����U�2	���n��]���R�T�S���Y�GC֏z�Wl��lR�Z�]a*��h��E��o��q���v��>�
��wF*�wU-һp�}��n��)]�̬�8�x*x2{��)ݭ��!,�:����7�u�i�N'���d�J�:*4��n��u�vq��{�b�[�Ϟ���w'��%{ ��H��^��3_
�(��^�^����[�1qښtd���,9��ex�SXuR�e��䃤K⩻�hM7+�:7�=ʅ~�O�A�)�zv`��zz�����e.܎��]��Bg�>W�1�Ja�.���*��4e��ٰ��~�t$ 2n����Mv�7�ы��X���k���q���~hk7sV���}�%R뾺�|�=a���u�V����G�%}:� T��P[��2�ӻe
&����cT��+Uj��^��m�$�3�����V ����,�]��kY~�gu�>}�)W]�0�jT�҂�5҈�i:b�D�%�l
[�^�wu�b^�b�F�l����NAX����^o}�à˃������~6'��U����FS��R�I )�x��VV�xj���dmDQY���ٞ3�͋�
>�1G�6��yRK�zm���]�oQQ���-tt��%�-��Y�0��z�=Xy{tk8�����n:Z�˫�	�v�*�Cꤔ����^=�d�k���+���,0[�=�$�s6�+K��=R��v��^��̎�܏=x�����\qw��Z��%�Q8��E���3%���^Aط�n��#�wO��/h>�p�[�r�F�ܥ�~��EvsQ�_21�s9�+ק��i������S�F��弍�]
"�3Y�B�aTF��K�J���W�[�</�4[w��n�J�V�m�_�oiY�(���lV����J4<��a&C��@�]*w[38Y+"�qoo������i��e�������b�������7�ޑ^�z�hu�3���+�� �^S��P{�m��9���T���k�w�Kas��G�3[����ԫuϸ4��ѭ:}-�����k�hݱb/γ�_�:6>4������!��c��:�4��Mk�.���Z��wW��#%.�������9�,�Po��}vUU�V�@�oUn���;�-�����]���6�i ��6��c�n_%�I
i����1������{�+¹IΗk;؝�*��1K�Y��o0���rsك^�
�������t���-E��ƬuA���E���A�E]߁n�-��d�����}^bX���A�欟h;ĬY����´��[�/(���ו�Ngl�����
�}؆4
6�,S�f�{+f�_*�):�mŘ�� �=	��z��u߲e�zWWu�������������tQ�u`��)S�[��32E[�L�M�%P)7tl�EW��\�ԯܵ�Wۭ8}��_������YH��rV%=٭�i@Ng������<x%�W����n�,,��(4��-5��љm^�����±�hv�xʵJ��ޯX� �2��>CU�`�-�;SO�t��*�6B~vo:q�a��-�����n��^�X�dgwˠ����3L\���כ[�jn�E��ҹ=�0h�Z�3�mC(�.r��� \	��H[���HPg�v�[�qo<�;s۵�c����9��^:�.ʓSu���t�'���p<+O0����M�c�)�s�Ѫy���_|���w��m��yݻ;�s�m6��胍��N��k�ԛq�8s�,sF̼�w��w7�s=��-=�����Ή|[��sB*p;��;2�9l����㴥�[um�8z�i�Y��i�,b�×���=u�f��ƹ�Ʊ��Ӻޑѳ��ґ�[��n��u�ډ͂�V�.��/]�S������\�?,���Oך�y����#nI�/�|�ޏ�6j8{�z��W�WS��86�Wv��x����b�`����EI���]S�ubgs����݅��M>켩�A|G����;ݡM��$�f��G���t�eN�
ً��*Ｒ�sÅڻ/�ߟ��7�Z��R ���б��1~����.�]�K�)S�z�O���TR�ԎAn����G��i�ӇumT�T�ؘ��;7zG�<IR��>�ګp�!m�
uǶkӪ4��ř�����Q��{��<�yVP�\�l����>�zz�M)Lu�X���N��v���Ɓ��D"�N�=����*/?:2�џP�t�q�oؔ7�����x��W�%���C�{�|��)>�V7�=��흅�\ͩ,Y���
��*��f�(����G�$��0���k���nsn.��&�{#��0�gY3�f�<�7��s��t��vޝ��>I����n�d�f��=��|wn�d�gr���)�v���
��(��WW`��^f�9k���hHk�����wQ�fx�yG��b��[\����U��|2�א�ٻB��Ү��x>���kW�#�~�*��g��5�׾��#�{�zZ�l�^Z{�n��db��g=�l�WK�{}�d�U���Nt��qA�oLw{���y^�0����Oeb�;���V紓�}Z,�s��	��}]��X�y�F��$��TG�)�/wj�n�O^������f���߽)}���
���̏���!҅�y*�r�DͬY��,`	�)������0�Ӌ����.M� �����uɫ�6���ik<}��{Ra�/��e�ʉo�r���5�|�Y�/��Ș�������th�S��h&�z�m�]U���+���b���kl��g�va:66�#��w-q\D�E�i�[N�D���ȥ��w�l]o���J�J�ӧ
�O7W�ˣ<�G!׌<9�yz\bp{n�R��V��W��+Y�)q���|���TJM��u�^&y-܋�U��7g�g��*��/h���ګҳo���J�Wٺ�#!��U�o09��ܱ\�>ӣ�i��X�W�u&���(���h$�W��j�f�V#��8��|l,���(�uU�v�t�Fn�j�cR�W��W����f����5�n��Eo���>vZ@f��ذ��wybKVY��r��N��́��A��z;���]hU�{�cF��8B�t_Pr�-��t&u^���N��R�}̚8c���;gt�p���H\�w%���C���t����uqu�tsh��/9.�]��9�Ğ�fqW#B�s�A�p����bg�w�i����N���6,���z�Ėw�Qz�n���%=m�@5��s����,���3:A��n����,cA�H�ΗS5Y�:��3��Zv�[��	uhE�՘��y[�5@��ǻ;�T�;cG"�V`@�&n�*˭�`5ζ ��a�����Ƕ��F��8�;�u�|X3��Q���Ũ�eM�v��N�تWQWg�噡M�f� /�<S��񗙨\+�񩷿���4-hpÔz���dΛh��>ns�݋�6w>�]�5�u�w�rna��Ģ�>Q+���kJj=��1Km��j�d���봡2�:���8��(��1c��#��F�M:
�K��t�����Ie��G����.��N�oei��f�1�7��:�gzT��x ����y^lVh��+|�v@��U�|V��h�}���wt �N�VlO{L	�Fs��R'���3~D�ܻ�M�f�r�A!�f����4�|����ws	����'K��C�*(«Ǐ��w�w��#a��6+�*ʑ|�T)�|�yQ�u���s�s|�Sza�}7���j%�B���i����n�)�/Yy����u��o��Uo(�ι�7���|��b��wP�� ҇�U�׾��n˿p���z��nwW���ei�-.�b��Ȇ�={k^{�E���+�{���!]I�q��ĩE���j5����e�,%w���֯��6�h|�^�8�o�� �EmG���(�Ka5�[�۪�:c{�n��.$*6N3����� D(�}�y����vg��Ε��m�'LS�>��W��G�e���r.�]+�tn�.礫,�=�R���<'+�A �2�hI�;>���w5�ݵ>�zo,�/Us�Ө�L���QYA�O���>0!b��ٕ/��p&߅u�����-B����Ǭ�ӧ.���U��j�����>ں�^�159�`o Ʈ�9G'w��T�*ݓ�o��mvL���	{���|������}{ަ�n�7��ؖ;�uiV���Z\����9k�_���Q�^3�+����]�qK>��y�w�d+F��xE\�p]+��za"l]1""^^lڰ����W��Ժ�,�3e�0&p�u�*x^N��On�� N�eMvs7X�w7)�XG����s��l3�{���ަn5��_n�z�Y�s��9,(
b��S����ؘr�iY��V�Y�wt��v���2z��o:�@�#�O�J��99R<���eZ�XH�����m	�v�v:����Q��N��U>~��)%���l��;x7d���s$ǭ����6������/8&�C�-u�J�{��K>}01~������簌�h�:���*ꇽ܋+�mT��/�j���D��)���&��n�+n&Z���3.��q�~�wNz���W�0��l�Ζ;���*�/KEd��<K�z���ԏs�}b���^{��ǰ1J��s�)��Ca
4M��M���e�vmvT�`c��&u1�:���x��4N����فv�c��]�R�sV�O� ��O/������o��4��o�S���Kh���``��^3{~C7�W��;cm.{V��ee^6K�ðo��n�[��߫���ZN:l?���^�7��K,�%V��ϸ�<��ɽ�w��s�.Zc�"��32m���{ڏ�������(
�u���1қyR�nJ�:���PN��g�1�ftx�(/�ptW���FΗg �^*,m�i��NV�鬮����z_.�36�])&uex�e�c����}�׃[i4D�ʕ����;d��{��.͒���kk�j��u�7���E�#v�ێl�.ޮ��A�a2v��ܡ�;V���ވ^F���㷝	��V-[���yf�v�GuAn�������Cf��OGuz5��x|�<�o&޸�qI��M�೵����X�-���Cr��oXO�>��s�<'n�~�����ˎk �t9����t6��z�ƙ��i���X���A��<��s�뫍Ƈ�!*�����Y~\���Z������9����/��υ����g��Kᗓ*���f�R�Z�*�[���J�1,��;k��T-�4Q,S ��o��S����+�7i�K�9���t]��;�������&��k�@��2�m�e�~ܔ�r��g�����a��������x�"�nT�렳��m%k�睼�p}N�ޫ�}�1g|w���T��.��ܮ�!�/���
Y���v[3���~��]�oqIW-r(*���9��Gz���6q�ˮ�����Y�#��po^a���^�b
�X~�ٕ략�>���.�$�6o��{�XN�����*Ry�aE
�)԰	�\W����9{ʠ
���5l�[�����ի�@u�d��k;�D���q�g���%�n^�U|�ó ��c�o1rld��č0Xk��)W\i�ș��Ýqr�q��I�ͺ���f�:��P̵��+%��%�ήp�Y������f|m{Z��ϖW{<��4֨��(}C��)�Ԫ���E?���m�z���w"�S��{�K�n
��S�-��
2�[��OOZ�������چ�c.���L��]�Le��g�v���Uv^V��R����D�LI_���\j���儬{e.�@�9�x�̤��if$�k����i�����~�̑��G�B�t��8Wf��W�l�U�n���D6�>Ž3G�ƊQ�A[��y�T�nx������g*�qӫ��d5K!�m�ކ�Ŧ��{;��wZ�ӪV�Qj`&ʿ��Ȩj��43~�+~qߖ!*�C.0�%l[*��7)�UM�E�Cw2�_pw���s�-p�ѥp낰S���Sh�R^,��i�8y��p��b�WWA
�t��c@O�\�n�tyfC9�*p�ު�3>���L�z�%��>޾�O���MSi}b���0������(%� ����<�V�8�7^�C\:���^#�̜��7\�q� �	-�姧kݳ�2sY���;>-��^Nچ?Y����v��^�O}����C����七���yZm��J�W�{�����U���T���
J�6w=':�yjyK���ή}1;�\�Ls�T�اo���;8>a�0h07O]Eg���}�,eZ5�로�\7~������(S�j���R@]�v���u�{���{�t��s��=�^̫Ero*�s-\S<֔߈3t�ecu��r\/LN7�emn� ������%��俄N�x^y����[G��y㖏���� ����5u�#Nm��^�3��&`hjC��z��
��S���Sì� �I8�P��'�af���e�u�����r��/��"��v��淦�:�׈�c&��A^�s�M���t���x��j�Ih��ݏS�eP�תy��3�4#��uY�J__��׼=�=(���N�c�2�޴��X{j����p�2�d��9��Pׅ��� =5��S+2�_?J��>���<�H�� <lRH��<4 ZC��nkv�{��:ח��l��r��D�*3�t�`��*{�dZȑҡje��]O�{u���Y�Du{���! ��V��ԑ{��K�UKU̥a
*N�YY�p��i���I�m�5�)��*$&���5I5��eA/��p�ƌ��}{Ɩ{��.�O���b��EOG]��7�I����_eIgݞ���u�ރS�4�U/����CR��^-�v��0~���!oca\�s����=#Y��
'�r���O�zS�9���.UZ�S��͇�k׫�+�lƵٻ!X�n��\����1.j����>������ޟi���]���s��R�X�{0Ǹ�v���6��^{(;.�_h�F��m ���h�p)<u^x��,�iY����ܛ�.2�Vt�Bh&y����̟f�qq
u��Ԝ�T��nE'�j�;{�hT�~M�c�U�q�hZ쉀�����r�KU�T�j�����qDײ�P����R�Y����.�]O���������>��:�n�L!}��ehU
�M����Qr��'WC�Om�IN{3��wc�bg�75=Oo;�ݣ�Ν�p����������yI�&�[d��f�R}�'t�eO��c�%�*oH2]G�7B	��R�0m�9��}�jg���v�����P��i#Q��K��}Zř�mk�&S�Ҥ�;��z��_̕�ԫ{7{~������e�O�)��u���f�>C�5��m]ސ�����u��s-Ԯ����Ԓ~�绕�Mh����M�%}��T��M���=����N=����V��G*��%
W[����s����Ǒ�{أ쫵YP�e����5�*����EK�{t��''�U%e���}q^��p�B���`�Y��Yo�<7��g佶2�����b�b�2��ڧ�ln:�-e����?֗��"�վ�%���Z������u�_�5g�Jx-��%)���3�wk��$Sŝ�7������fV��sG8!�]M��PB���b�T32��U�-�PoP�]x�'&L�����X�Uf�Ӻ)nm`��e)�/ɽ���k�޻����i돊���-��c�1��� .{qu���M�k��n���\�;d�C��8鎸+c���u��e�� A�;�Iϥtn&����"�1p{:�N^^��s�u�����^9��j����h1�p�gg��$7[s��J��9�,����=6�]s�P}�=�����/o$n7hN\�c���Eo.�2/.zZ`���� ]�V�y�l/�]c6l;k��e�!����.[�u�j	�z9SBuk��pl\;0yݻZ�;���J��[a~����`�?�`�ϧ�O�r����Y��a좪�S_0��r�Tr���Ƽ,}�lL?;Y�)g4�{�J�Ò�Mr�W��t� Pl�(��e`�+��f�.��W����E�3RfT�ǯ<!�]3��f�!�rh��3�P��*��}t�o�KØN,���X���dJD��$�%1��	B����������c��V���z6(��W���0g�]o�+C�Fנn�=��j���<���U.���q���;�9���j�*,r5$�ʱ@Q���h�拑�Ji�����J�BT/1{�ި����*A�^��B���;��(�#
���:ez�S�YM��:���~�Kܚ�dR;#��B�-���o6�>f�ｕl�F]73~6�*��0�;��_n�U��wH�3,�6w,�"��}ͽ�S��^;��ǎM	��gW��]���p�R��o`���v�\�k1�G�=Wg�l��K��aN���cfA������s�v��4�t�wݛؼVګs7{jS�-�'%
���%>����{�n��5��nQǷ�,yN	�u���u�"��	bZ(QZ�s/�ڙX(��V��� QyP��O��a��ȗ��M�j�ڃ�G���}}EZ���P��c�2�7Iٷ��Yۘ��1mQ�t,�]�Y��<tz�)F����*���f�դA�{��]V�p~�N�o݌��)*�y���eM��i:�~�2T�ǯD�]<���MT���?;��),�{�B{{<�75��nrQ}��Y0������C����q��mU����<n��ͲR�*ž���5?m�6��8�!W
Ի0N���=,QM|���0t�F�JX�������-���([��^
�ת[؅mO�Z`J-o7��[�z������	�"#������������zQ�rxQśC�bʯ*�8�ք�~�DʷOry9J��/춲��k&q�I��y����}d�тn	��̹�Q��:�����jC�+[d�D�����nq����2�����9�6���=��<�y��a+G҇>�ee��+Ɋ��>�뺰Pa�E�v��N�F*{��7h��bi�`�8(V � �h�MJ�SŊ�601���O�Y�g���^CPxZ���<������z��i��ҧ\�q��YywS�[����s~N*߇y!���b�O-���uXR������c��;+3|�ܰ��wج+��Sh�ˀԄ�<u
b�뗔Y�L���MV���x�[47-��9�h���>�>���F���ݣ���a��©j��	�+�2��M�l/�/�7�����X��9Ʌ ��7���dX-�&[��`��nJz+��%��� ���n.��V <�tˉ�`o��Y�|a�:i�QA���2`g��糞�oۚ���<pS�ɏ�*�U�.@�%�RH��t�6�;�-w�;�*Uߐ���r+:��f��-𥚘�y�U�^�B��nW ���e_�L!F)�����obf�0|\���uF��C�.��'a�:6�1�@�L���[�[Id�n�Pn�R���ms��UBT��*�$lUk��<�+C�^Q�$��%��M�?Y�����u�y���e`��+ï�ݿ�B��#W�2���6u���Ѽ���J�:�D�����j�+�|�^{m]^��ķ�Q���z��{vut�X�^)��xD�s��ڷ��T>��{Tm��h�n�D��*��}�r�}l�*DG�|�v.>��sk~�d�����D��>�9G�b]=�Z�tp�,���]e���y2�]�p\=���vjyR���c4�R��9���ܨ�oz�����	T�N+�ww��|��H�3UR�����*�vR��>y���tV��/CN�I=�� ��V�l�q�8o(A�@��[�L����<���޺s�d�?u�Q�PA �*N��|���n����2�V]K��#}���}}+��3=,G�k� kx5}2����^�u-ٺW�*���÷<,�U��d"�$4��H�T+{u�)�1�2�N��ۋ���wgsv�ӛz),�T!��ƄH��^6�����>�f���'�fyW�n�>��l��Moq󬣖]�xM�V��~�@��g-N[�*s�L�w�]�Rd%N�i��N�W��[�'��'�.�;���f^z�a�R�H:u�fP����OӦҿ�;���'dd�U���V���o���yj��g�E{�|�X�$�H�6�JM��> ��Y�yR�ru*����J�]�n}�%Yϴ�]�e,�	I=����T���lUpȳ �,��ad7�p$:i���ӧ�.`��>|6�w�-����W��:Leg�5�����R���;�ux~F��
�����Ca�U�|���Z'��`{u-��1����I���xz[���?�_>L�?��߿~8�����k��)_���-��s�D"�.������5s��V(qB��S����UUr]��>,Ak����]b�7Spd��\f>�:�1�ig1�݄*�����u����*��?	� ��ƻ GM˨m�ez��	����:mI�����iC�F��
̠�$*]g��,��"���"��=*uvZ�;�)yWBL�$�v��B�s%Y�}sAJ�Xb�V�&�r�>9gͼ`=�.�G�i�E8��G5vc�L����=��E<}�[�ٙAJ
��¹�:@��&�7qHP�ٶ:wh��.����
b��9�T�o7%��'�}�KY`��?l*�j��V�me���yd��������Cq�t�>�5�Ӌ5��K1�s��]��'+	܈e�������2�*ns���3W�]D�Kn�jv�l��4!�:3���(�i�U�v\��8ḭm�/��ub!;]�޳vb��Y��{�E�Ѵq�'�ʶ��.�-����5�,>��h��8,��{��p�ܯ
J*��}F5�&{�Mx�(��Sϭ܄�3̨6�%�+����Ib�)h��D6�_��^��j�^skWZ۸x�j�N���p�u`c�\nPeX�A�@�q��VU �4.s�z�T�������ٚi=���f��n<�M]
��Әsgi��F݉�u��s8����` )$].�<Ã���Ӣ���+�͗��y�W��^�9�@�3\ͼ7���]d�tq��4�K�hf+��٭3-i�.Wj��m��s.���6�$�MQ�bԤ� �V(iG( @�P,��$�!0u;X�=F���Q6L�8]���v��\���r������p�\m[HN��\�����9{u���X��Mcn}>$qmv�4�q�Ƹ�u<�m�;c�����׺{ ��G=��wI������sv�'kE/��vݬ�٘�=i�N9��	�s�� 8��q\t�M��hwY�K��b�u�����yN�-ό�\u��p��q����<��A7Wu5���=,낵�/hR�>�`vi5�y�g�5Iݝ6�]	it��]D��j7��Û��ɜvS��d��49Cla9���eGJ^�u�^�v��»mٷ��ϵ��k���'��m�w����s���մیspc��s�i�=G�s�\�[�i�ݽ��ձ�}�:�n��]hiH^�N���:�B���e�M���dg=���S�w�6��O�����GX ��S�=�|1���ηvm\n�'���'K�76V��=O��uV�Ø���ǵ˶
񅝞R$ݼꓳ�3,��V�
��7c�����Z�y,�8�ݑ_m�+pf^EzH��Z:�Ij�ó�kv��;fy�:puq�v��wS�컚�ۻ�-�ԭk��-�Ӽ3����<R�^x���݌�pnջIn�t\ݗF��RdبS�䍩n��_X������Cl-��7W76vGnͻn�ヮs��]�I��k���q5���\�1飣�7o=ۡ��Er�[sĝ�=X�R�\��h���hEݯX����q������Sk�n��!cvNy����%�w�6��DM5{vm�����F�=�]�� ��u���a�镑,�mX�x7���s��n�-u[vS�Z�e�N���6H�k�g�%QT9<��x�����k��m��l&�7W�5��;�W����7a+v6:�ŜYw�Ghqh��n�=��1���5u��<g�������� �w������k9���5ϕ3i�t֋jc
������]�9��^�q�kR+3cf�g*z�������p*�����tu�՝5��\iQ����7۷�%�)�*�2�kl�e[�4k����8�w/:��{Keݭќ�`90���Ķnḏc{s���ܗnssZ,��%8`��$�1vܪ� ���
fc��F���k�0]�W����1�%�R;���@E�o��}�δ\ �rm��'^��QZ���n7�1���,��_ɿ�
Y�gU=j�5}O%t�ʟoj�_K#=��T��������j�!�����5W�oV�z�U��+t�b����E-��	0h�ѭ�+A�#T�����M{+]x^y��S��[�W�þ�a�E yR�ϭx��0�Aܱu�׷�|�פ��������|�'P4
�O�i�t�.�rS���U��ҝ��>�U�-4��#��d���e"0wY���[���L����^�|�h�޽+S "ZQ��C�q�dǃO��oc�sQ���b��̩��ޕ+C�'e#��qM��<�/)X3�M+�3���,�]r��L�C��.�uݜ���5�����5jZ��s�V{>�o�J�0ܿ9�B��r�J�@A�u
~��e[��������b�	��,�]y2�c��b\�ܳ���J<h���{�r���K���C�Ld8B9�� �-mױ�;����Ci`��~��گ�񄬋��J�4�p��қ���~r����Ƿ)j�	^�%�Mn���0��+=%9٪V�����X�YC9"G��-�M�y�L�[��/��4�2�a������C�����~����X��P�%j�ْ錗z�8wq�F��!��K��qX;r�M۬f'�����J���{��N���.���ϲ�QZ�,|�d,��%2i3�9^��FI��F����whr�K�a��q����ң�$�x��:�;�a���F���?A�c����>�OT��=ؑ��c5YR�P�۩�©ã����ά �!�~��������{@�;J&W�N��}�ʮ�Xf�)�l3F�-�R�*�0�i��3���*π����g��~#���Q�8�*w�u{����s��mO�F�)q�c{�t+k6ɞ^��X�ߌڤlѺ�O���|��{3�ݓ�(	(���_��o�y�����+�EY�u�Օtr�Mmd����^_4����T�*`w�wW.�r0��b�9����Lr�{6nw`�Ÿ����VP�79!��=d�Y���hٚ@��K���P�/��P�+��}S%�o�wc��]쭿�$�,�ng�9S��q�i�u�٨��Cj�qB���g2�e�&|�7\��������"�V���iv{0_��H;���6Ej��[���cr��9�]�^�x�A.lyc�j˵,���h.kW9۵�G�^	U��BYcn�����1��zj;~�FC ��W�o�n�� ;{�8��w�یq�{5��ĵM̖R|ȧ� 6�1�~%�"��Rw`鲲�B�K�x�}?W�2�o�U����wD,�r��v�,��ܩ1TG�� ���I��U,�������'��P;w�Qў��WW��
̲���v}�3���DQG�5�Mu�5�R%���ǫ[5}�6����X}�Oz������i+�JY���i�v~�*��>�9���4��v�	�9�ʕ]Ơ`�,}��z72�����ɜ�_�R�^���P��l�ˉ�V��X�n��Iԟ�}wǑ u�3�͎ۧz�Q��q���B���7�kƥ��<y1�ͳ�^��?��ŕ��PX@}���^�����:�`M�L��{$��N��>�j���ϴx|�a񩓚�֫�*��EHP��ڏ��4��CNe�S��D�|����-�{<�}!b�g��_yl
�2������?u�[�I�pe%!�^yW2�+��$�=>8﻾�D]�Uk��J:�[{���Y�r�q�J�D�^̙�K>]{5w{�c'�mp��[c��ׯ��{AJ�5�^���|�˽�v���r?7c���>َ���|X.�-��Y^��V��#f��ʟ!1���i`�y���O;&�{
�j!d��v`�b���b,��*Ğ��}9eܷf�AK+��)*�V��.%|ts���,���2z����_.�Y�l�gW�&�U)Z�)m�s9�
��^e�q�V�xh[Z�0Բ��$�];{�(�O`�݃�{{was�t��AX,W�}�a��?C�+U>$�4�`�ѥ[W�i�m��*�UG`�,�㔍���g���U]�]�n�sփ۶Us�gm^^���4SW�V������	�M#Q����un�ӲT�B�+�K�+y���xQ������5ziߦU��I�a��o�GP&*p���s}־�1��xࠪ��ԱV0��K���Sx�tΖ3	��9�������)>�[B�ƪ�@�ֳޯ���Z�#�ѭc��-�8����Z��%7���k��Ow��ٱ!���2��� o��W\�0|=;L3�!����X�b����5� 4��W�(~�,H��	�����`��ъ�1�M��|jqrx=�&r���+W����i�j�� �s*�ކ���k]+Өj�t�����F9͜<��U!�J-u�~ЫQ�4{����lj0,'	S��p�R���:�L5V��/����h~���^�EWee�i�Fs_:����s/|t��-oF�qԭw�7�{G(V@U�}o7�a;az�s1:�B��Q���:��l��dm��Y9�K������V�rT�1�����[cp<��vD������<\sیX�Ş���O)t��&Ę�\�n�デ���t霏^N��
�v�<�����q���g���ӒG�Ƚ�p����pp%ǝ˺��y��7��]Y����X��^�t���g����s<�S̠S�t��+է9�[s��=��a�{ALn9��l��'�fiH�s�8��x�PyѝѭWg��f8:p�N�+ў��qs;c{���V��^vR7 >�	N��X�������{����}�HOY4b���8����}��ŇG`�y�~ש$�^ �u>}�]�=����߸
Ϭ� �QI5��p�{�T�^c�pTӿ{8\��_�Q�=��4�  �7Y�[�t{�������pm���5�}BT�>@�7U�	��3��mŪEi`�Z�hf�]q�w����~}�)m>�7|����ژ��UW|�a��W���O��*���2�V��e��p�Zd���E�A���[H�٘{4x`�9����~��b�����G�hX�@��^sO�fh�Z�Q��o�-��uJ��TƉ�~~�}Yu!�<R@�*�
u����[:�����LS�m݋����%ڟ\�[~��(������L���*��A��\�pU�KK�,������T�u��Z 9�E7tT�nڷ[��̝"*m,�B`�]�Bv�H�6J#�N�ֺ���Uv�fwj�f�n�3��;��M�k��v�M4/{�0�(�Q{�/�Rf�nc���ѥ5ʎ���y���K��:5���C��)ⰅT����ߔ�C����g�����و<�ls�2�Y9�:�ohy5o�^�.u��-gc�!�X��)�ol7����xeE2�=��C3�ѣA��X��u�.�g�w���M��}WK���>ҞP;�W���P�9u����-�lj��o���Ը��h�w{�_���Mdޜ��o�º�s���;}6��ռp�ro��ע*�֮�����ɵ� l���K�g��"���Z���imU�����}vx����յ��b�d�"�1��fHU��E] ��˨a����ٛ�y�J֭dΏX9.d_^�~u	�����u�8�m1����o��Y��ֽg��j�ΰo�+�����+7��~|v��&X�3���j]�+1M���:Iy����ᱝ��W]y��q����_�����������y3�8-���cn�����ܩf�.Ӽ��gk�(y�5r�R���}�O�`:,���|i��4���.���!����آ*�O��KR���x\���V���L;��_�q����϶Y��)���A�T��(,�Q��(�޾�uq��5���(xA;�W_.�'����>}��6~W5�j��˻*o�K�ԯ�~��)�������r�j
���(�֩}��g/q�w�n��VCY��j�v�����QW4���a�^�kDV�����l���V#=W�i}�/M�!tvB�s� U�ʴ������Z��VMwD�m=��|� �wc��M-�ɹ�)?\�'0¥���>�7Vm�Y�"�d0�U��D(�{���W���1&Z�����#�*?q��8�y��K�b�.ii7�2�)ԯBV��T=�6:���-r�KĐ���c�Sy�SFfF._�Cߺ��meW�Z<�N�:��%����j���U��C���W"V��-4�.��*�ct���>��n=���'7b�,j�1H�l����lmkulZc]C�9� �d��8י��5�<޵˪��x���Ob�>c%)|�r�*��������jCY-U��:����A��9�j��ujz3�5����S�kE�r�S�;�'Zu�0f�u�m�x(�����͔�2vs�w֗�n���Ƈ���^d�T,7u�~��ʗE����+��0�J�Yߧ�/��{�]g*[��>`�	�&�'�1��̰����]ۼ�&��ã���1_\޺�X���aH��c�X������ ���>vg�� ��Ԇ���I�餜\��E	BЫU��۹zw���j���p�ڱq��@�n�m�h��d?AU=����u�w��{+�ag�4/��P:�����h�T��ʖe�����ʃ7�8�5���m"tlwլB�.i��7�Z��T�ɫ5�҄��+�a��2���W.�EeJ-}���q�F�[��g�kg�����;��n��������5��}�7��ެr�0}]x}t�fg�`$���!��Y��<�ut�lh��m뮌�z�CItu���<@��1�=��������tuȰt� 3~�Wn���TpZ}ӷj�\�?pT�,��Ώj�f�E*�:�෯6����
�Os]�^�Z=���	��׊��)ch��c絧�s]�����Ycí�C�!�yږN���{*W_����U-�w� ����%G���R�j�z��D.�iwU+�W���yl�?�1' ���eŧ�M��[^��:����y�,�i-�'��{�ocWu���[������/e�Ub��#��F�X�j�VG�Q0�M8�-����i4X��=ܮ�}�{Nlt��ݶi	��t�E} �j�����b�Q�2���C��o��Wn��&����Q�z"h��N�i��;��<*����<��o��j��S����ׯ}�C;O¸�Ei(SX����R�|AF�j�ы;��&Mx��y�U��K�[�/j�yym1�����޾��h��E�����/jOhj�+}�]��Ya��I�pH���g�x̯犥ܨ��ʝs��m�qk[�a��)Z��y1�s�w��p��x��h9v�^� ܜn֞qѓ�\��.�;�[�Q�<�OsV�Gc�|��\�\:����m1��g��}��n��9SK�xxvz����>6��f��rV��n��;iݱ +��Yr�=\�y�m3c[��\v�lw$��;F;.�'��c��.3��G!�<iS����p�!���я
t���خ-�Y����A�NU��.��^x��S�����[@C[GM)���5�
{ֽ��T��E&����
"�I,V��7V�1������#L{׾=G���N�@@�H�&�k��'ЀI"vP�������O��r�g���?^�ٖ7ݝ��MsDBd}r�V
��X�Gs4Ϩa4��İ����:�Vz�p�˒mv�8�@
-q��l�7ŝ箸�V6}�|��}
��5g�^���f�X��n�oT�,7��ӎ��Η�ٻ�_bz~�Y[��ز	�$$�U S��[N&)R�lz��unt��]���]֬�ܗ�����`E��%CSi�t~�����������Qrzʛ�=XJfs��i�A7a[ {]}��4������{XN���я��n^�j/5�V�+��7��@[��Hkq�N������t�M2��y�=��8یr����WM�m�K�Trn�p'i�'0�nlM�.87\��ư�5���pP�mw�prw"���3�4;+9�A�u��o�R-��5�b���}b��u}�}̥бQgO=��P@#L1�����N�BW�O7�G����ɥ��h�������nWt�1���*MT���C�h��jiW��q��l��k7����v.N��Gw�e=�vD�����o�vꂼ��G�q)u��	
L�ws�m��Q�N�Qo��s(���������E��^,��q� ~�i�&���e5~�[�q��ʕzi3A��7�ٰ�򯑫����(��,����w,]��J�V/e�(/�0���.uzƆ���;E�M�����_���ʱN��o��KX�rp�OUMd&���ۊ^�|�����3��`�YZ������	p�N�`Qd�I������S�ls�6na~ݯVы�D���U�M*�s����R?2i��
�������yҎ�4��{=�3R4r%�Ɏ��%R�)!`'e�m��u�7@�۩^y㠴v��.x�I�v�.�i�tB*�;���k9�}��5sZ�z{P�A�i ά+�z�}]�S^G"���޶��{ϧ��R7� �:�5U1��+�3�NXY}��A�1��tP+䓦�T�L�״ֈM�e]�̩�fut� �ERƾ�;����ci�Y�O|�WC�xù�
�������^c�^�=�����������{QS��mYn�g�J�T۫0g�c��;�(���*�W��2�������ĭvT����erÙy�����j�ߨf�}��"n�l�&�S3���1b�����]'#��\t�ee���/V�^5H�@���i��o��t�Hɥ�QhV��{h�܏�)��t����K�w��Fv�~>:Q4|.���W����θ�ֽp�i7�-R;��	�ԅ���c,�I�z������k6M�[!ۅL[��mR�/����uv�G�崝�R�]��C�|�����|;t�1J��z8�<��R��F���̓vP�8����J�8;�*�.*���̱� �X�1ᘦ��qH�A���2�MnFl�2���ϧ���ZN�[�ϊ&,�{��aMǯ����v�nPoQ[R��φS�{��}R�֭m��F�m�I�2�	�w)a0��L�V�VW��5O��+}�&-�Q�y� �i�B=h�k�1x�Q�:�!��g6�0�,sp1�-�}}�4��Th����eL�Yvٛ�.�Y��V���p�a��n��g�Q��D�۔�\m��s���d ��ena��=)cje��V`������I�զ�
J�;�*�c7�u�z�rӯ�����<����#q;VϠ�J�w���7�K�/u���/k9a}��%��i;��r���+����kc��e��h, u�s��I���us�����ni�%[)�SU^V�z�2��[�g6�aT�7=�Vk^;��.���D��A�Eǒ�E׵*T���W�A��H�t�'��"�zO�s�6���FhC�;U�Ε�S7P̻w[����Y{:��z��
�w �ڂ���<<��ӸU���h���p.�%гL������&#����O{PJ�~�<�,��q��0aC�r[��s�VF^Y�ޛ��yܲ�2I��,�9��Vnk�i�����%�@~YXz �#8�����u��$X��)n�Hr�j���"/NQ]Guw��oT�\O�yl�[�k���W2��$�.�i�D��7^6�vywmv�:Ƅ��Cuug���xU�m˝܊�kr�vq���ߵ�>~���G�Fh�ݭ����2{�>4��;��x=�Y��c[�X���ח���Z_��]�Ϥ���׼�ꚁH�n��E��0���/�K��T?9U�
��Y�ޯ
�4>0n>~����H�Jy�yg9��u*�W�6��|m�k�͠l���L��E5�v�]��q�L�(�;��>����� X�ׄlv�Y���c��n�Wy������(�rQ�WWgr�T��'Lb���x�^'l�x�Z7������tы�:��Йŏ��z��ژ�4k���O)c�ɐԠg�����u4`k�K8� �-�;��=ۻR�]\n��[/v��g������e�NM�.ݍ`�κ���lU��*�Y^�/z�����^Y���jjd՞��$�-���#9��{�;�O��0�#J��R�u��v�4d�������0|�<%�I�o��w�q��ayKs>����N�F�y�3]O���C�3�8H�q4�V⒝�"n=�H�l���tmwk�������k���>��Ķ뫇њxE��-�o-�IC��v��_�w��2dnf�(���>ɞ�^��� ��o���n9".�+���u[�ju��?O�F�0Kn�{��0!��{�2�c�uN�QLH*���Ӻ7^��IWܺ���+��L1z׬�p|E���d��Yx�˦��^�
a34��wյb-D��YZ��6�{��r�+�v��4���[U�8]��Z�J�~�h�6�����Qխg^*"�j�vZ�OL��v
&��E�o�@�*�E�2"y'YwDFnT�[�^���lE��Ƕ���9y��m�����ZU��W��k�Bx�
9;*�
5^^_?I�q��)Q)4�u.��]�ݞ��"9B����L�՛�ή�o|È�ȼj�AL�^:ܥ]��-W`�vT��� ���Ds����!Yz�
'1��uٍk�i����&;��b�YP�- ּPU��Uu���(���U���}ɏB�j�,�O�κ>�q�j�+�#����d�*gq��Dܽ�,����>�l�Y����m�ݹ�z.�V��f���n�y:�X��N��XK{/��x{sVV��z,�'+�Xp�>ݰ�ѻ&����/]�l���+��]u�����v�K����E)��vtsp��va���-f,��ngcm�&7��2�<���N\�Y��63IG`����٭R1�ou�HN0���[k�ټ�k<F#��4Wf�u��(��#�m�7pq��{Y�!V*�#,���]�n���(��e�J�VP��ݔ�[z�+��"��#�+��c�儆X�.�׵�g��Z�8��J
 =i�����r�}'u?�_uus3{�k�i�wRu���$N��V��_��vk��X>��G]`��kE�+��,�\�&UX+�bU�����u���S埰G�x��B�.��G��wTU���5��xM ��<�X>�������c�W��<���d�O���������W�R�}��-��ll��p�ԢT@�������ݰ��o,��������=;{2�w�oχ��Ō"��ֹ�����),��!�C|/?ŏ2A����\���i8�ff:]�;���G��]�c72�ӻu:��
oUA�A]/�5���tntčm.�=�x����ݶa9�7(n����spsv�;7L����R2W`���qX�Geq�h[I�?>�\�0Xq�/9L-�VP�k�N�3~���h�����/o��3�}��^����c���$w�
S��B���0�Jb}kE�FG�K�gB.�ǲ����qݍ�+12�M��]IKˮ�� �#9�mf��4�uX�"�x�[�@�y�p�.9��'Y���/Kw�O*t�L�A���{޻^��Y؞|p*C΍j�����V~�N0e]]w ��H
-�,}a�Y6b���\� a�t^�/�NU�i�S�°Ռ����w*������]r�C1��/��C����Z4����j��s�ㄆi��i�Ω~��4y�ODf}�X]2�`��=�]{�ʾ2�!Wgڕ9���C��1�L��51(̠ʸ�b���>�V]w�F� ���B�M�8z�*�	ACO��*��^��t�	��3��1�Sþт��S.�2j	�bZ��vr~^��ׂ�/C�;�=U��CG�p>U��],��:�[�|t�tb:��ǘS�6�v�wI���Q��ݻ�{=ϊ�9i�b1Vl�RTJ�[}�*z�7�*ͤi������о|���f1�<lh�=��^�0�����rr@�9�(�"�n���u2��[��;,���7��J@�ٖ���M��t����Ue-�;ו�^�b�jMY�Z�?.G���'A�M
`ߪ�s�?e��?�nh�^��4��I΋.�Q����5��L���N����lE��++3h���'��̙z�:��z� :���zj�͆+�Fp�W[��egu���ĕ�)���C9�+ʐ�ee�)%<���.���ͻ�wO=��m���B)i1h�]u����F�[J��6��q̕�
�5>o���eP�������|��ٔ�mTU�G���y��{cU�>����TՔ����"����c�]-p��]OU$i*V���y}v���S��4�]��mb�.���ՂN��̶P���n��5��%��N�+L9��\�����N����y�5ٷ=��n��v	�M��Q7Ar����ֵ�ۼ��׽߀8\4ٯ=�V�)�(�o�V��*�s�4���s+�	�ZZ(v���Ϣͻ�PJ�{��
h �^wW`h���n�t���9�Ld:��Ğ�'R��ofX�*���n���Oo5ٯe���y�1<�3���צk��Q��(O����.۪�h�R�,W���Η�>�G�tP%���ަ�8�漏\S�X}�j����>���8L��S���3o» �4X@�70"�����.�K��[=[c�.9H��Gպ���<� ��[�=k<��N-���zV�V|��e��r�q��x�)��R�L��nF�P�3����+u����9���YR��}��wpIGQ��bYn�aV|��JZr؅0|��go���]�,�&=�{̢�2q��KJ-�����Lg/|b�\���{sz����Ž�/���<���џ���y�r������荔8$���+��k#�S��V&��}/�~Ϫ�o�)��t�v���L�)���H�q�;������F��@�C�M���?��'��/&��u��FŎ����4&!-+-�o���Vn�U�&`��z��-n��U�A�b�Gs��}��qF�������!ԥ��<�3����� /lr=��z�u^��J����L,��i��`�Q���De�=�}���C��d�F��������$�U
4*�K5}��(
��nk����7�~�#�iѲ�S��s~�@��A����QZ^�k��̣�e۱Y�`$y" 
�B�6ȕ`�?+�'+���@�fͫ����	ư*���h��9~��~�����'xxQ>�k����v9�2��:J�X���X��R��`�Y�Sh�z0<��>x���.��	�X��tߒ*��c~��z�����c��쨺����,�@_�_�rF��y���	��?:]�7�e�����J���J�^��߄�m����FG�aSf�IС�ݩ�k
�k,��~��h��P�[Aƅ�j��uݹ���F�������e۳өM<G6�u����.e,G[a�F����/j�m��<;�qn85t8��uv�+��� ���=��1��Zk�!� Gpg]]�z�ǵ�� �w#����1���*���a�6���l�Nz��/���Tv�۴lf�����*]�JRl�b����y���R��P=qqq8�2�֎�\�e4]��N���n�ۜzM
��/E�۷<<��a�bR�4���ݾys����f���^�w&�z�Z�o�+�E���6��ȏ��,�9�:B���{��� E�E]�⃠�$&�i �l]g�t������v�V���FU��k�%w�<��ڼ/��>(D㥷���M�􋝞ٍ�14;��Q�ͱ��׸�4jV:
���Z�N'J-=ON�+Q�=�a�w�ڨ&%ti>�r��쩺��`� ��W�np��4�)M���m�+���|�8�j��ƌ��h�d�����7xpS��w� l-f����b�g�J!�Gb=y�j���)m���ؓ^��Nƍ�5,�B>�^��`��%R��[~QQ�]�'��΁�""\]����$�#�y��2ڼѼ/G)�Ul�h�s�{�Vd>*9J������ZH��	�In�yc�awl�����h�ܓ��v��E�Ȥm���n�"�, �A������;�|�#(��A,���9f�v�ʵ�1q�g�&��`t�
 ���7�=�]���^�y챽�_OACqZ�+:��ת�Q����؞�f��z,`"u��Vy���E���y��������:�9>���Z=+9W\����R���7i�7���g �;һ����q�*wN��C/��鈩����As�{��*KU�je�;��_����rkY�S�c*�ڧu�Q�:^;t��Ct|��v�]ܩk�JD�L"ZM����OƧ�f�����k�l��)M�De���v����OZ�"z��yBd��X�.��t�G⩤�iPI3����K�J��*��/:����w��@(.}n�|/��N�'���pW�&b�X������ܹŽA�Q+z�����pA�h+�V��j$8�S{�3��Uc�5�bf �������8w�]�ܴ`�C�o׵��ڳ�%��k��Oa�y�l�=_.�jp�U�I�s��PfN#���7q�qg�Δ�z�.�3um[�x���c����bƠ�	`w�������_=��u��KKzf�!��N߀Q�V-=G��*����,�ZL���Qw�A)�)7���%rQ����Ü�;hN�w-�`d���~�^p��P�x�T��z+��o�f���7(�����V����,�����jG�`���9jH�����hҫ3(��ھ��UM��%����q"�+."u=�������,�p�����4��v�@v�o��m���)��D'�gT�q�m�̓F�ޖ%ߪmK\&����t��x'68���ʷ��!J4*݈moyJXh���j~�g�<��a�Cz����VQ��g��.q�������}����O��u$�ү�Q�57w��Q��K�U2M![�_}��4,��z2�К(|/��]&)d�o-{�54Ե��#�f�7�R���ʬ�]��Zv��V�{H���qj�����ɵ���')
���ť,��mn�f���Ƈ�F��X�m��t0�۸�g�YaL��b�M�Y�JfLR�Y��f*`Ƿ��x��O�>޾�����@K�_7��Y�4ó����Ƹm�at}4�ʵd�8�U!J�,�a7��9l�x�t3������
�4W�p��ʼ�x��x��[S�)��C�-a��q���V_�lP���k�/T�]�H�B�ChjdL{qr̲�X��"�O�1�v�Y����%Do Cf�#����/F�m�qn�V�us=��l���B�k�u�1ۺ7�9U�:�q�]'���%��=~-�)T����{V��ao7@��qv�9�;z��v��硫E�ց���0I�z��:s5� �~��V�E �	����g������t	:����RG>~	m.s�J��f"m��έ���J�~��xT8P�R�
v+���?��7�]%��.�@>�Q��߁��y�ޡ���P���� �qA&�EnW���]6sm��x㐫�M�F/j��/ۺ�ޣr���{m4->
��9h9P�R�l�Ͻ������i\1$v�G�k�<�4_�<�ef7O�wn��eh2������Ӭu+�5���޹B�>�X��(Qd2Rg4xH`-$���z���5u��V}�n,�&dR�Zb������tF^����|=A�S<s��Cǩ���ۃ��%�mKEͱ֮��g��yHkj��+ٜ��J%��:xx�����5�8׾�6j��A�kr-�R�1]����X=P#L�D��M���Ū����Iӽ�D�����啕��P�3�-�ՉH)�otʺH��,����
-C��},�W�n�[����伙�hQ-�E$�̞�+N��}ۧte1���&
��Z=�->�u.&�(�����F��<2�̼@�����폪Q���g����-�l�R��0>�)��[�^���(���'�49�B<#+(Ox��Ay���hffY�����v��~�y�qgp��9����DZ�9�YgE.�{�V�*X�5�����*u�z��5�b�	�p�b֪�+;����SwEn�]���3�Ѿ헹��ѡ���m�r��j�RJ^-ź�l����V�\W_%BU�Z%�ȳ%#�K��t�	�k~��'�]:�UmVݑ���vh��a;)0e�3pFw�o��*)�;�M�G�ɥ��w�nz�ަw�BƻW"�pޗ+N�v������Kvj����l��dV{�j6���R�u�)�����R�d�#��q���ݓzi٧�
��H3(������v��u�^L�U^?���(�"s럖�}��t���T�8��[�K�U�+w����T��y�j9z"k����\�Ii�oR��6�ݱ�b�0P�{ӭD7`=4R<&	��o��#�vV��Rnœ���U�k��.�]c�i�җ[Z�J��0����c}Q�b�uX�e���+�[L�4�����K.X��a�z�R�ڵ���J�N�vM��ճ;�"":��S�k�.��j�٭��4Ы+�	�\������t�è�&穻{Bj����lx/9O�2ۭb��ܙ8:[�ݻ������Ce�=�<�}C}���?_�����vqn����f#N�����Db�8i,M\�oۃH���'߿ꪼ����t��djG,��Ҷ�fB\��!=հ>o;pmkay#����ǲ�0S�s�yw=pv+��c�d�����3�8<mse�Q�i�cnS�F���v��+����uu�+F����󻋚�4gu��$w\3�g]�r�۬x���Gl����]����/5�"^zy�k�N��^�\�㶻ob��
s�Q���C�����n*�p��^�����gi��Ⱥ'�Z��N�\\��z�U�����G�ܬ<�mƸ�]q����{j�Q�yL ���<�Ʒ�{��y�F<�۷����tE���a���v3�' ����-��6x㹭��t{p=p�SúۄL�nώ���쇍�D9yu��:+>�\��F���cF����;���1��`��PfT�=���R�6.ģ;Xpr�v�ᚌ���E��H�=��ZݫY}!*�a봪:0�s��F�Ǹ%ϙx�!��63�Y=v�ۉ�W�cr��� ]�p�z�l�-@;md�:��R�'d��-z�y���l(��׬�l���hIC8��c)EkB-�Ď^��m����S��scA���y����x���۱���G`ǭ�M�͓:\��6z܅qeev�s�����]�m�87��[�c\Us��t��4]����n���눺��FC�@fĹ�����a�	�\�\����8�v��]ls�;��.����o��O=�]�-�9�βs��n,�Wl���Wcm�q3�h� �J��9�nlXq�+����,�#�|������ҍ��k�k�8�Q�K��&wm]�ۀ��JÇ���d��,iL;mk����N[F.���և�Mt�m�7*^��v��m��n�pc��R��q�C�ۮC
G�;�û{hS��5�8ۚ������ͻ���ۍv_M�����7������Iď-����xk`�ñ��o:���5�rܼ�j�7�۴��6t�ѓzC�/T��l���-m�z��gg��:u�sב�����^4q�';�n66'^���k&x^�l�콷G\�v���;a��58��crwݎg@�<</
�Q7��D4�� ��s��rq��
q���^�pr�N�6���R��9�^�*����n�F(�� �yü�O#��w�8 .y�խq�,�S�[h�c��].���\V����G���/E� P����ivh�c7v�R,���������;	�J�*���4��ќS꽏^�Z���1�m%���v�)�:,��� ;^3mܮLy��v�V�ac����	('Aʚ
-jX��񥂳���cY��lz����p�ǭS74�����[�=�%��.����������TU��Ziz�V[��eǁ6P��Z�W���d5�5��ʠU�='�nQ��z�e�/�X���$}W�r��E�db�+=��P�4JU�o^\ռPe�B`[�n*�GǷ��R�ʼ0V��6>���Pf×�ݗT�{��p�	y6�Ǐ�߽�������C��E:��/��ϪJ>�*��G�ŧ�Z�s������zr:n��6G�6��:��Q�z*�Or�Y�LR�O�����<�+���E��t���V�!����I�o�<�7=&�FPp�'v���=����.:��.�Ύ*�u9D��k�V��S�g8>�aV�yOx�5��|��U.���s��
��p���)���)���<��\�2��OY�,�|nτᩢ�Ю��j;y{z"am�=c��L���(5 �����o]m�H�Ū��B�Z��b�mj�n��fwU�f2T����v���Η���a2�E�^'�q�]K#ݫ�j����9<����}�7�
�bd�XF����%[h9��8�{�ccz��eu{��n�$�6�]�����e�������֍U�~ �j7�5(@�[��)���10{��f�r�=�M�v>�V)����@Ft�y�W�Vj�'��wV��U8hƣ��"�z���ʏ��L�VZ�=դw%F�̒�h�����hY���]ۻ1���4>r��"���%��f嗅�pOT=�O���8��B�;��,|뱾��û{��_|���b5CVJ��t*����ʞ����#[�<s�|�t��\��|uc�a���B�̶>y�0h�u� �s��U���M!Tf{ʦ�Z	��g�q7ʞ
��h��f�<�vc��M�(W�]R���V��i�[r��4V���l���{��9��a��M�K�,�2G������[D�n�Wa^l��b�c~�U┄gб�E�}�SX�@v�K���7��Vyc4;�/�b��d}�<n�t��*Ziˌ�׹W�e-W��dy�W�T�I��F���7
�5yd�h3Oފ��f��";4��k>��D+��ʐ<�޳疜Y���WC^���/ղL*���7 ���:���I)|�&��S�ψ9�x�`/R��]m�ۃ�G���b��yo�s��n��eH]�^fz�U_n�s~�?-�k�`���$���iR��
��hkژ�|�J*�rz9��Yp�Z�b�};9q�����^� :�LX�~��Y~d������K��R/pα�A/�������)�c��1v���˼��X`뭀�z�y�BS�.�P��gk~�G���Jw��!vkj+��V��ͭ�q{�c����I�(��.dL�}^�i���ð^���&L$ �S9HU��~�αeՍ�nԵY֫�Ө�'V^mݦ�|��X�q��TT���V�n����$.��YX7���	�-���*�@QB�d���X����k���ɳlZ��w��kY�����S��Ds`.9�Yˇ��m�e/x��?+�Xܰn��?�/ȭr�	e��}gs�lC��Q�յ3i�,A��y�s���̓FN���zu��xR��l! ��p���n:�_aK#/x�'
��aٮ#�/^��F"�Y���3h��t+�ﮰm9cBP����2u/z����+w�H�=c�"JL�*e&2������eE�|�q�B �ܭ�`+>�cw�Ǻ9�=����{�|,פ7p*��j=��C3��ק��1w9��b��ނ��(��t r�ʦ�e���]�>�I��g�w^}���+�NC��^h��GQ��m�[���w����3�]X��Q���s�+��NӁNFA��2�])�w)+Vu���Nw�Yꬆ�z��w�y���E��J[VV��i�v�ܺ�v��[�'c2���7/qO2�O��n��������2g�rs�z�c{�z*�3zUu:𦨯�o��f�{c��~��N���,b����(_,Q_xs���_�7�=
ͳL�61y����?�<��РĴ �MJ����ߞX؏�0���~�g���KlE��9����Xf�E��y��X4����W&���
�ݼ������R��a_��ح��5J}�sKD��>�W�rm���V��{ӄ��e��N�36����dbBx���r�ͩ)65�̽XƮ[�s��Z���D�����ĺ�2�;�b���Y�u��kͽJe�S{�7�I�++qR�����b�s�u>I��R8λ\��u��̖��{x���u��͡�r���d��WX9�<gLmBݝ���o%}=��_v��!8�dv6�F̞=)�7��:aܷ��(U��4'Fk��� �=a:�m�#����x��F�ex�Ѱ7�������/M̍ډN�dر�:��c�9����tv.29Ͳ��3��9�E�Y^�`��O=ni��[��vwf�ǃӻu�c��	�v	�yw=9��n��=F�;��h����UǺ�t[Ojǣ�iҳ��:�{�_]��pX��{B�8Z�b{=���lh�7-�}{�^���~,º�{�X ��#������C�s|�������b�M�H���.��t�p�?b�5B��;)�!|i�y��6�s�5�ۄ��e���h�����;󠘠E&�k.ng���gl{�	��b8� <��Q]C���b�#�v�/'�S��H�y��Z�Z����T��@���������^̿v���oW9K���B���=Y
���ɜo�񛞂�e�����(#�|��e�y��L�d�i&S�� ��6/ت4U�Y��tw�a0EEg�ߍ���˫�j��0��(��+�z����`�*E[�xT��TΡ�w�ix�"��յ���nHۈm�(Iw0�vإ2�+���Ƌ�7gY[<r�mx������lKT�6�y��v�qQ	���$��%�xJ�,[�/'f��߉O��ǭt���6��^�HM��:�s�a�WRn�A�*-6rv�oF9�����������JҬ6���^��L�����ݞ8��mĕ��m������s�a!�ô�Nk��K��(�+��y4_W�<�5��;���n�kq�4#�䯧���/J˾k7xt�
Yէ����Mo3^��%�HФJ`m��2?3���z<��,�m�
��>>Um�t��*	I�R�����,gv��by�[;��:/͔����o]9Q��^���P�������u5N�4 �
��qs��>v|�ݼ��N�h�T��St�]Im��"�6(�J�	S&��*{Rii����{�зأ����2�+}��?[�Q��4\{d�o�9�C��S��"���3���Zʿ�=:��v��w�>qz�oI۰����ɹչ�!���[���KUQ���!:�91Ͻ{���ի�Eg�D�^n� ��䚽��dI��{>����bY���֧�Q�x9�Z��z/��R�D�)�{R��;r��g����>Er�q&/�,J7\Y�=8����˯W$���'����Z(==���nAϹ����p�WA�-;������S ����=��(���e0 �]����N�N� �� K�>]���:Ym���">i��h�>�)���w33�lKZ�=�N��%6��ثƺnP��S)b�x�ʳ� @e��X�� @:��6�3�:�v���q�=�����6wem�{Z�"oةW_�Vӽ�>+/+wx1�!��x}���3h�E{��席�," �%��r �����W��x�/=7i]�u���e��3}Ϟ�Z�4�lvc�`�����[�J2�k��[[[Aka�8��n4^ۯ3Ƹ�Ƽ�֑�/<v��G]'9Umv�FQ��j7yw�{ݺ�y��<�y�M��$�V�EJ�M���g�?XC��`e����x���T���/)لF{�k.���!H��"�LL�Y�w��`��ng��~�w�U��4^MXρ�w�C0q�5��Ѭ��/r���]W�{%���F_�XEA�f�M�i��~Y�c��{^y,���q�[+J�"�#Ɠu��ᎏv��ڞM7}�{��v�g���noK@��DC-�{%5�fT��W��]���'n�A�y���v��,+����_��u�ɮ���.�\�X���^ĩ\+�H�t:>l7~M��j+�@B����h"��4�\���"��[����E�
�,�ͽu,7DI�Gt�w׻���P�d���aDҢ����H������3=6wfq�G����,�g�ݠ�|\��t�:��M�����4
���x�'�C��Ǐ������R�54۱�B�*F��������C8�n\Űv����[�:4.�r]�����4~E���k�ܻ�;#ϰ\��'D���z=��M�����'�L���b��@^z��-!��y��8��N=M:� ��V��]hcW|�yW}5u	�yd� )r�}�7S	^v(�\���_d�HX#�?�>�;hל�{������&���ln+��*��	B�p�F�>k��=��t�>4��[��R�箢�����+��lR�0y��/�˒�74��z���`��ИkGPZz3�ث�����X���	��{YS�J��e#&�.�}^�����;�`v|��V�z���<�t��:E6���8��3Dq�:7uf�K��g{l|!���γ�~�l��E�j��zO�ʱ��1���Ez����~�� &,`��n��E�u�
)��qt��#4�g_(:�恩� �B���]��ĵ�p�ʴ~L���m�����Y�Jk�z�����o]�X�]��Yy��⫳{O2OC»����rtYΕ���d�M�熖x�K6���E�n4�b�g����� <F瓂pͫ�=Ov�d�n�e��:�v��:7��b�8{#�9�O�q��*׮u����tŋ�p�tV[��9�n���c8���p�9qs�ǲ�s��р{V#��8���rm|���<��5ֱ{WX�>mgW%��#09>����v����K����e���}���	?���m�@�\�������rY�ȡ)�Nf�Pט7j��GJ�-���SZ�����?E%�V!4:I�qS��*\��~��w�+)"|9��x�gj.�*Ug\Nz�kq.Xۮ���Z+����zn��ko�IHx��%Y@��`QD [c=����ݏ���Z�����G7w�G`U�n��!����E���Ċч*�僴��Zg;��_,V�V�:�)9�aՈ�ֳ��s���t+��n��E-d��|�qy���WZ�~�������.|����[�Sxd�f��jg>��,/����X�%~�M��~�֫1۝�io���lԳ����4�KݴP�9v�w��P��J�9;guf����� (B`�ɺ�Y�}U��`z��ni�5u��=��v]�û`Z(V�hKe({|�H{�A�=�m�C���֟s���c���f�=�����!S��#kVZm炙W����5�}=]ⱄi�G9���[��g�әN�\y�mj
5"�1E(g��3(�<d�;s/2Q/���TXo������Υ&D�w�Ë�ֻI�6����-'fȺ��}65�P0J���|c�U���z�'��O{l�!�$�;�D/*b��좫��H"��bͤGt�xܽ��~#ɷ@����PU�����Q��%X���G���8f#
{�YW�[@@?o$��[z�>���:��gC��>ٌ�^���xY��>x�]eC7��PR��u,��]��'nm�r"��,WDRoN��TCd�@�-�˨d����7ם�X���j�\<i`ᱻ��k�Q�z��ͽ��g��]�+��]ҕ���q��pJ���4iP@���9y�[�^,�7h�*ٯs�&��Ewn�ɣ��;��AD%O��!&}Wս\Tŀ��wj�(����7`�?3|��:EǴa9�0�Q�銷yŌ��>�G�Ԁ���
�>�Z�M$L�v��J�����>󗫺լ�c�|�����.Z}G�|��t/��&�ߺ��$��������q�g���j{ף�-�U�TI ���~a0���@���1�ΞW �}����w�q#~�<��޴���ڗ6��v�ni/h��@黭�]���"�p���+,R�uN2�u�R؁W@;o��bީ>;�T[N��c�A$���/ o��Ξc�m�8�e�XU��T���6��I�iZ�������G�w�ʚ�Sn���%��
��t�[gƞ������5�R�8���\���Pj�S���NoP�mAb�@�h�R�V��N�+�o�!;)F�5����c�bρ�B]$TSR�	,m06Nڻ����5o,���է�^���,�k�����i���2жdw^6�M�n��� n't4��;�n���Je�eyyVAW/��[�dk\�������s�X&��q�а�Qɫ���0�6vs�9{g��˸�3n�w3>w�a�wd��u���i��[Uls8�#2ʧbzkhL�f�ܾiY!K�A�6\�9˓
m0��.�H��	,o+�</od���U�g�ߒ�^A�^uu��H�'�E�R��t�ֺ���×V��-��/:D�ojz]'Y/v�e�O'��祙ۣ��o���G#�$�k�?k�����a$�~X�� X+�T��{l�U���R�-mRV�ҝ=aȧ��f���]��>�oJh|������1ؼ�->�M���V�r��:���Ya�}�æ�+�:���w_$&	1*Mvw/���4�y]7�/��7��u��kw�����o4��Ŝ�Ry�2jW��e��0�b�!�@a�Rgo���Ŋ{�t�<ՔÁ�)y�wջZ �/s���mVO��z9V�-�ڒ�e����Oa*��G�T
�*$Q$Wc$��
�y�uB����_V-����Uw�������ո׼����a3��]�$%����u�ih�X��>d��(��������=#����G��exD�s�-�l�mG�������7z��p�֋���կ�ܦ��az��A�VT�_;��h�C�w��h��|��]�(w�����M���0��*?��w��+K�%-r�X#3��B�M=fj�����臝$#�}���L�����(Q�:|������	�Ƣ)7��˭\5�_c��<ܬu;�q�=�Q�������zی<��mh�i�I�C�"��=���:�]-$�\���3���w
�q�0d��}�nܜ��>�D�޷~��1�{(�=|PS�{-��vR��C���*�-�e�>q�\�	q���`�FWf�7��'K'����3EYO
و��O�ک+�Z/MҜ�m5D*t�4i�ו�����8�zJ�?f>�1Z��"������������J�W[�CE~ѽ�Xk���u�>��o�V��4�Tr>{Wt	��5���wh�!�pmn��ݱ���i`���{�W�@x���,���=:�v?���x�;�6�v%gm��*��uz�ʱ�k�0nN�^���<��
_|86؅b, {��Ѿ-���V3���]�{v��o�e��R����Kb�ׂc��i���=6L�y�ճ�&��F���rTRJ�@�};^΍������ɨ�
������g�M(���f�t#}���Y!_���Y�<�ܶ��#����,��A�ԁt�����&{�!�Y�7VMr�ʉ2�p{�x�X��>���4�a�g���D����2U�����|.+
��N����
��}���^V��ٮq.5վa����|d��w���µ4�'x��z�ؐY2�>�e�����%�b@��b���PT��ƖE����a6���.���W�e�Qň�f(M�f�۴5!�⌡ey_�k�ϳ}�l)"�A�R*�l����oms�)^r��7<�ڻ�eÐ�4��ա��Wd�u��Oro�9H��/	���(���2�z{jv	��U�s�꽰��u�ܔ�8^:�������-H6��m����ssn<v���^v�m�v�ɚ�L�31�/aFzɝ���9�&�Ⱦ��[�����N*��n�cj◉%���v�V���]�O� ��5ӫfV���!�O��$aWY��X'�b]f�BKG������j�2���y�Β��ks��Y(�4����7B�_��ݘn\��hc^u�o(��̱�ս�����hP)�f�P�5
�����<竳7u��0�\Z>0�{�@v���� �>>��$�f���0{�h��,QEJ�4M J|7����/}(�KC'϶%8�{6T�L��WoN�^'�W�T��ƴb��hI,��E�����hQhM�~�cZ[��R�t�V��]-��n�wc��/ҕJ6���l�[�g�:G7�<���ݎ�ˍLsv4|��ӯ�Pt��|�	e	��y�(Y�g�{�Zo���nU�~�t��֗���*x�<���tސp�,w�E�[�w��L��G/lk��p0�C�W>��e��\�]M�n��0knn��C��
��j5Ӽ1� E6|����ug1���N��$�����Q]#`��v��{��+�=]�����c6z�����y`&l�@
��:�D�	�צmeY�g9z{}5:�cg�7@pF���JRYd׎+�s1�<]���b����e�V�Z++w�oWL��\Xl��x��q�Vb}Lƴ��̣7,���]��K}&���t�!���2k�h�Bo���wzKf��)��2��ݞ�B��5_��� }NvTD|(���~��^~�]��G{B�N�L���{�%�|-[�2Doi�G����Rx}{\8�5{1ө��Z���K�@���];��5(��S7���{D^~��w1�q�nV�����%3�R�رtw|]2�=⟟��^ar�
���e\
�E4D��X��^W����=/N+�Ҽ/��[^��i�{��0&z��
��h4ۅcc���^!<A,�1P��ѥ$�u[
;��	a�]^Sd�=g����ͻp��q��rT�(�mK[&&����Ts_<���=v�z7���#@����&Ȩ�n������3��C�i��<y��33��^E� ���R:�.u��D�����8��*tG���4W-�u>qȎ���&Fl�[c�aK�=���a��a]����@�-�6���j�y�N�k�!��Z;-}w�ymmn����k���U������$<Z��Gucq�Cw�r����m����/ѻ���a��X!�Q�慃��yeͲ�*�q��$�0j��"8����CΙC���*I�M�.�h�f�7(�Cm��h4}5�����5��]�0��˸��nf�څ�l44���Ô~`�T:9�I!�D�Q�6J�.^~���;��"x����;,)i������b��IE�C�<��ο7�Z2�zB5�,*W���Om�T�	"�����rA9섻�ĕ��W\�<�vn��:7���<8fm�����_���~z'
����]��E�6��Ow��Ogt�z�r���[��B��w���X���v+j�+V�*��4H�/Փ�-\\��x���gm���/)�K7>�&a�jl��zOG�B�N`Ӯ�6[m4l���,`��tM6ﷺ��9��b� KB'l`ڝ��dto�u�}捽���3S�]��ϳ��Gjn�&��^[�}��L٠T@E>>˛�+<C�+����߻�Fz>Q[98v���i&���O�t�e{����[�ߞ��Gu�g啈̿39:��u�\��9��q��̙��<�Tu�Kͧp�vu�n{�~xF��4|px#b��r���w��Y�/WF_�������:*��˵X�)�S����o�\��|�hB��F{�;���e��|�X{�t�1%Wօ�W*H�I/���=���������H��v�Y5��Ź��n^��
�v٭� �("DS)���.�/V�Ⱥ����l�)y>:��f�{�� �A9%m�$؏�ׁNeQ�+�Q>�E�4�  ZjL��Y��y���fO+�ʝ�w�5�D�����N���\=��%��O���M�ꬬ���[�_�Wxd�|����	:,:i<��D���M�g����by��M�H���y�Z�?ZKޓ��N�n��*��]f��T�`�`?N#��?ew34�$��	h�$f�Ӗ-\NOX�Ǘ7���y�Ze�&*��v��Y���.��{ޤEmA�h}c3@�g��2=c1ׁ3�|7�T�K|C�=5��K��+��r�G��`�����/2���^BP��8�Ʒؓ�A�w@n��:P�V�W�`Z���{{�m�'����zt�5�֯	=�'��U�̍d���J�Gw�@/��yIݗ��<�l�՚&'�Ķa x:Gs����� (�L��;//f��痮�H�u��/�qt������.p�[n:���v��J��l�{M]�[�����`d�I,lkV!�S�����5�������.;t'���u7� Nw7uq�S�����`�m����!� ��uۛ�kֹ�n�˗�w�cwc��w ����7@8�ݰ��l݁8�U�)7�5O=zG�=�;�vvzqڍ�MV!��xN����ph�����ՊmX�gu{-�3l�W-��/�c���k���]��+į�7}CǉI��T�L��3������낌��B��,�x�H&�A�e����&���f��;Yi�%bƀ�7��(ש�R�Q: f��H:s����w����[ߑ�ə�Y���8JY���5�oD�fOSK����RƻW*�ֺ�Ծ�9�{wy��``"�"HL�.Y뫱:m�A赹ܬo���@��*g7p�kk)�VX��DM�T.���ZC=��	�A�@&��-󼈗����B�Q`�6��#W{�Wec�:�&+��]�3JZ�AKr�A=�Q �^$ͫ�{��#��_?��+��ՎCMvPn��c�ٽW=�x�aԗ��)�j���ggb��֬�����l�|��޳u\��0���G��Kݫ�7���.����}W[��M<�Z����A~q�05��Z_�1�U/Ωz�~��*RSC+� ౢ��4p˕�Ŝ���دX��U��Ѣ��%�gM�����_׫�]�W`RX_=�#���R̘�)a
�c�M��ʰT�S>���s�� �R�o;7þ�
�!%)%��h��0_ev+�;�yP��򩋽D�>�����`Τ�k`�����'įr�^ٻu�]0q^,�SB��"�R@�^�����w��gA H��;��}���]VN|�����U��WE��w'rk�'=��·7=��g�#��6B��d�w>���f��C]W}X�b��5�f���gku�x�b�P���6�sCНLjeD�����y�I�c�?�j�pYn����$�qm�é]5�m�]�fy;��l����B�ҫ�˝�&��w�T����s�Ѐb|rE{TU�`��mD��܂W��Z���j�&B�5K�@M�D�^�F݉�l�߰��x�,�W-��>���w�Y��nw�L,q��>�)H�#�$���co�׭��k5��>D±�曀^��:���{���u��T`f�~;�vnA$�;q�6}dz>�@��k���36w9s��i�o ��{��D]�ek��6�r���:46nΩ�ڵ�i�E��V�D�>�P�����j�m��ֵ���]� H0Lb��3�@Ű�C}+x���,U�ɪ}����	^,���o�*�����/���3���D�mmUݵf�kc���C�`e2�5�����	.���껜�7��e+�! ~»Z�5�=^�Y  ����ڞԦ�fp#3w�^�ٕu����Vym�x�>�A���s�|n]�g��GJ9����[rd���q�fyѮ���˩�_0�u�ȓt���{�2�.�H�fzx�C~B^d͠�d�}�y�fs�E��G	�7�'��Q��'��v`��<��<J���$ht��ρ�K�Sw'�0�Y��.�eK�YH���-������^���xQ�f���Q�xʤ(�߯ ���9<[�i����Oul��y�{�ֻ�JUu��v{��x�z0��8d����6N.����
��֔�L \7kÄ�֍Dû�~{��`��ϼv#F���]j����hW�f�OJ�=I�Ee�i��]ߞ2碤�N)�u�Z}i�׌���|$�; �V�a��&��y���[mٰGg��ˇ���z|�6vQ�ˠ�4�=5S��XZ
IFs�=�Z`��!��r�+��w�ޡ�u.�zA.%���}�_��}X ��6��̓�SnK��hq�[o�JȨ��#��qԑ��v��p��bn��6��dm�i�� "�<o���/�a��Ԥ�2��d"��)�=%7�ν|��w���%��Zܪu���ޫ�5G ��ux<��	m�}fh�MA�ᛯoR�'.��.j�>$��xy��Q�ɒ��Np�ܽVx�m2��**�g� `R�A�-Q-�ߵq긲�ŕ����ɉA]�<���)C7]��پG�N�x��J����y�x�5��E}w�C��V9-s˚�x����WoQ��r �攫�����G��V��-V����l&��DJ�b�+�����
.fur.mOX���""�J����S.��{�cA[�L�9HmH�7��/eNHl�ͪ��<,
�涜����j�쯪-Լ<�KW��z��	y����۔B#�\��boZ�.�u�(lU����w^��ə#�*,95dN,Z���˺R�i�h�8vJ#�WL).�e�S��E
��z�Y���sX�Wm��J�Wj�Ц�y{"�*�`���j^�Įj�j�m;���������4=`�+eX���cv�əu2���}�<r�WÎ�����*���3K�qn4�֩�YF�U+T�;��WhQJ�{e�Q.�c���g�V�2�"�cow�a�'v6xZO���L��=�fO�ޞ1����^�\�ntcw������9�<�!��)]�����d����EnX6��V�2;�_#o��P����t$��t�e��� e�d}6���!ޟh�����v�0��v�<��Z�ҹ+�͊pat/�N�v�-v���zvc�V��Kǉ�&�r��l�R�����^����zCSw�vnZ�ˠQ��`��2�'�R��N���;�2-��Mq��]Qmto����'h��w�mj`Y� Wd��ݭ��
�٥�Dn����n��巗r�j���1��e�k����VMN���D W$�˽�j ~�7K��[�&��,Bx{�҉�۵ך��6��l�c)�M`Y��H��]\�X�*�wY� )�!wt�@ڧW��Ks0��f���a�n^��\����.G�k����U�[��c�i(����ŝ�Zd�`?B�_�n\'<��j�)�v;8/4�n{@�j�ϗ���ۮ�&�m��v'W<�k��%�6�db�k�\�ג��@�6ڂ�S�W+�B2(��^���1�{y�w�cW;���n9��=���g�.�);E��Q�m��-�OA�l�s��ي.wFs��|���v��&�M�n��k�"�n�t�̑��p�Ĥ3��x�j��<�1t���K��5�+O���/3s�9�`3ps�g��9y�㒷��l�nqh�"^w#j��������F�dm�q����s�ݞ����ݐ�;G�#�����;\�At���٢��-���uvמP	-��O6a�zw��=�6"`���ڮ��O�:�
܍���.��{�ڗpb���H'�]Wn�ujBԮ�
�]�x��݅���Nٳ�b��6�s1h}��uiKF۶�6+T����G^�q�=�ewg��cH=�95F��=���hf�n.�{p�n���n�����얳���T�M\Qnܾ6�fڷ70�v�ô�ct���8���˷Pnw=FnW��:܈��m]��l�V�{��ճ�v��t���}n�c�=@tk�.^�7\"�룎���:t�ƹ�Pp�۲��۵b�N��'�T�a�s�]u�&��t7Z�'����:Օ1���pWgs�)o'=��S�]��fNC��K�<��C�3�uۍ���yn5&�����I�!Є�O��o=�[z�<��듮ʗ	b��E��ǣ'�=s���Q��Ƈ�=�<���nM��9����N�˧�ӫ�Ku�x�;�#;b՜9=^�gF���"s��!�������S��4�iw�ve6����#]/�jd㨂�X�)3(��t��5| Q�1W83�k�������\tu)��q�+r%�pK۞֏&'�f���8�e�(��9��rA�;�#v���gcN<\h:ų��(��S��^�p�L�d뵫��+���/]��Y��qk��v��^�uv{i�>��V	�ՃX��2m��7n���l�ܹ	����x�tskO=�nhm����]pv�z Ճu�<M�;0i�XDZ3�nA����9���`+''��Wj%�b�s�q�����&\-��x!��uY��ճ���ݑ:y*JTz�U4��3;\���8�E��rƸNG����v��i����M���C&=N�69�:�vv:ö�\��[��a�o�.[��aJ�R{\�N���.��EA�B>�}-?_7!����b�Zw<���wJ^����/N����[Z��?=��TY�v{��u%Ӽ B����r�{���^�>����v�WH�N����/�7��e��A�v���".E�+"�Z38P�GO�8�8�L@�L��fdۘ��./]��Vd������dІ8�m�)��N;���/_�t�|<�7һ�ڤ�0h$�Y����̼��]�l��Ͳ�O���X	����f���`v
5���j���2�ܼ�w �Q��V�;�/W,��(V��_X�A��7�<���
z��fp Y嚱o_gx_��Ū �/Xw��Vl�֥��\�}�ג�0�T�ՒZ+{u#�v+�����}�`��E�Q��=� lS�V�˞SD2�����s�a��v �c��dy�� �=�*�?��p��-�n{���qLˬ�}�>�����$e{{�b���g$K��1�j=�S��O{mֺ����k���P���{�.V\�eق�k�r4H��6�z���w��D���-�n�?0ߐ~���9<s�76Y�r��y�{v��]7��^��hg��qVhH��آC@��]�}̑�׆���B޻
Z��3q���Bdl�՟G��b�Z���~�U�:�h����-�e��Y§���;��>����sʳ�Z�vg3����d<��w�k
Rw�o����p��|d'�hל�+�u�SO�M���߼��^�y�8:N�g�u����A��c.�8=��"�qΦ��y�Q�JD�5m/��:߸o����������QT:��ȝ��B�Ξ6�1�rnL�D��]���uM67A��uv�\�{5���	�C��ޠj+LM���������{�w���#,�s+�qH�y�%��^�<C��&�>p'�^�B��2�����K�#�{g?��:D�y/"u��,�����1���cG+�W2��Z�7���J�":���g7��syk61HF��G��>�	<̢���ᦇxƁ�|�מ��rz�~�m� �p�'+�s�y���ؒ��C�;���sH�7=�ɰ�f��1&&'���75,���n֟Y��^�w����I�t�<�X��}��0��HS|�?���?-U��?5�ϩ�,��krҘ7��2<r�	"�M�Q��`}�1m�b�k�/7�`s�{��ޖ�)+(]����8�IM���;��n[��S'�t݈��-�+���{��ѥmgR��*���%��^�b�Y�{[o���/<�㶍��իjކ�쩭�i�$2m��u�#���{-m��x�u��n��'-roG�)
t�X�x�Xf��������V�oǀ�8o{�D��`z���xP���A�9�&^���&{x^�а>+~��-j��U	��OA����3�,X����v:a�}���G�%��s���,@�b�:� ��H�@�UU?�)��C����ZWW�H����Yk���O��%�ڽ��q̄��Dv��x��ws=����֢*V�����%G����zJx���vj]F@���Ѽ���	/�̙{;��3�a~�k��w����X�!
�Q�#�-}��E�'r�'M\�tTWB���a��8�]N#I��o2��*/�����g��u���^�VW��[�W��3����+d�\���e$=�m<�/q,/`�zDـ�B�^�����:�k>;����WQa��j��Z��/k�GFc���Lc�]�)���w7F{r�H6�M�:�Z��z��v�g;��
T�{3=�T6[uk1d�!�	P���)��{� �z�{��pb�R�4Ll�o��5�L2B_~Vkt�"�v�Oر��XǇ[-�yA���^�� ��P��NzU�ֈq~ʛC|MuF��j%���u.�}׶������2Q}�U���fZ�O���=�TW��J�ʌ��^�=��j7��ECMoP@:�d2g6wL�h�0Gͮ���������ɱ_+/�Q zz�~]ب���xD������i/®W"J�H�ڰ�kiŝ5�������椓~;�x<ϵ�@�I=�3��QYG.ڹk��-&0ۯ 2�*m��X(.�b�4�w�H�/(etŋe^�e@b"ĥy;񗗖bT�dG���9{��FŒ�=��N��\�X;��unnY�q���h=n۪W+��[�L���{��*�:6�7`�s�X�	��s��՝�m�</cnx��+����:�mfc�qv�4F"X�!;:��p�ƌ�ڎ�tt����^^���2�E�kɞ^gl񷣔�8������?y%�u��ȞV�'���ˌ\�-������]6���wn�7��ݱ��/9_]��ԜOOfN�;�Yً<[��%�7��i�Jʙ.-]s=n:���)��l�ln1��^������?w����hnb�ۥm◶2�<�����B�E�7܏d��Ѽ��֭j~ˬ�����#C0�ޥS~u�>%�ڙ�<&��$��z=ݯ<�$Y2��Áim���d�g=Z��o\
���7sp�%m�r��FzW@��i^�U7) ��>l����w�sTZ�ڝ�F�(<��b���w�+���Y�/����\�6r�o���k)���ʽ�^'NV&;��o9�׼�'s�u�V����҂=�3<�������[���(�8=vxn�f���J��F7n�/���u�@�}^��D_��-��4E헭EL���([*�����n�>Ȱ���1��R��ӯΧS-x֚��cď�
���a?��n6�x�m�#n�;L������2���r�❎�)�
�/o��U{G���a1���9�������!S8u�a����L�7~��<���ki5t�-��4�(6�Yw<�T{/�U0�4k\K4t�c��O}��
�̷X�r��ʻ�9��Ν���Yd��ަ6��pw2�Uuy�S>�M�,��3Y[����f������u���>�]��t`ۇkդ�<��u�6z������)S��ߦ�rɕ�Q8���gd�5H��vE�-���_<�F���s�{8�5��5
�y�����@��n�����I�o��˜�� �����G�Sͽf��^ܨC��)�t��[-?��}u��gɬ����.=�O�s>�pf�گ-�q��,[ի�Q�\q�{�l����a�A�sO 	k��%��������`�<߁A���G���},�@��&ruu��U{�����F��m�[$�Q���9��W�ہ^����:�gG;�ؕm�l:�@��mw9�/.^n�iw��Y����#4�Sސ[��V���T���4V,�{<����+o��|�@��$oՐ6��>�l��\+s�h��pJ�����ԣ5�O�϶����o3�J��A{�RU�Od՜��jt�ɠ�*G�TE
G~G��Z� B���i�*��G+�}�<6ٲ���v��}�egw$�4aə� 3j�.�8��ҋlVP>�{��w'�&��e%_�r
S|��Hz,R�n�ۭ�Ttg�Ou�����菉�҆q:{|du�˛O��W~�I��ڳk|��*<M�{�8i���j~�Oq��w��Ճ�R�c�F�U�S͉�WS���x�kWj�\S�3�4�$v���3�vg$��C�L���i^T5��$����;�fZP�>~
o���-Wؖ���F*l��<�F�Y���(mh��/�����v�;�)�s��2��+�ض]u�����u�mB�;c��w�xnkY�#�je�N��2�s�׽��+e�u��t+���|���Y��9�E�q_	Hs�O�m?�߳�r.�wB��& �[�~���]��;ݾ��>��+bv%��ž�`�ק�a~CجK��zT����J�ׇ|34�I:H�n�؛1h��EkS����7g,�|'ms�yV&��Νם�sR��D�*��&�^�\O�>��~i`��;f�Y��4� ��^���d���N�݌�s��<���z�0��8K~��] ]�$V��)W|C�~�����)�4��4�Sł�0a��]�q�׫ہ�7o̘x;o�/��6%�Z*���/���	Z�ژ�g�x��G{1_�Ln�1���IY�>��p5;��^�{떩��&%G�v������	�p�Y�k����;�.��kpOZ�'n�y���+�[����\Eʫ���ϧ�?�o�ºָ|�7�gOk/vV���{d�wO;����gWz�Q������zi��u�>iWg������z�`�)��xG�����ܭ����,e�F�/���q��J�^�z���z�z*>636ľ|��^��t�a�="�S{R|�XT�&�$��p�uü/�7:����022-�{��-��J�i�֘�_3�[���yFZ���8�m�yZ^��G��!�͒E
E5|<$�/�XMj�F�L~;�-�*Ec{=^�1 (.q^9�;{9{ts����б�w�)����y9Y�4�q2�c�MݓZ��φ��E�,�u��k�L]@��vx�[h��\|<�DN��t�7�������QtN�q9�J}�^g<���Wy�c³�&^uepʜ�GXg����[��F���m��ٝS�ưh0�̼1���I6�P�E�`
 ��[u��ϣ�tn����ݶ\l=s�O��:��gP�nsn޺�]�8;u����^���eX�v�}vƹ�C���V�S�����އS�[=bv*z
�ė�hM�Nv'���F�6�[m��'r5z�;�l�vŵuцv�' ��Ѹ�r�v��َ5�`:�3q�Mqٽiܓg������u��i^-�mu���5�:0��س�M3�ry�9��Е���a+�f ����u��H���t���]eY[�. �e�#)�o7X��K��� ���S��ݙ�wG8ܴ��*溨�@A�M�o�<��^96�rWi_~��-m-'�����b�~n�η$ u��G�d�8�n�xLov+�]�����E��hkf�u��9��:�җ��wY^^[훯ڼ)Ka��yL���L����ʾT����p^���u���^L�[|�U�(.�����~+�.�a�@[~�o	�h�U���l��P�w��?{�W.�N����_��٪����u� ��YBWp���`>��˖�����K}Rf��Qރ���Z�t)�o�*r�����Tw>"�RU�Mc�[T��VS�"H�ݖS�����c����-ټg�=scI�l	�Y覓��������-��B*���p���s�{:��Ყ���Gz�BU�Ƴ��<�dS�Pƨ��(Ҡ�t[y{֙t��{G�׺��Wy��q⨩�g�.23Vn�x��d�Lv�y��2����SV'~HTtR��T�6Jv��ʄ�y�����@��ǛYkk};u�����r�Nr}5��|�R��Ϸ�7���M �n�i�4A�\�����e�}���'��G�x^Q���]U��Z�[~y̥K�l�|k���Xgl~D
�r��eyl�5*��!Rw�u`�`�^�G�/%sA��=��LWp=���^x��+'۔�K�{��9rx����6j��z5z�Dܞ�l�$�e)n���btW&���k��;��25	�z�π���\�|=��4��Sz)�MM���`��VMs'�B�m$�֓���7Y�R�� ���k/=WZ nە�ØI�5H�;���w�";u���|D;��':��E�h���]8��L;3�z�V���L^i�A}���Y����x�%"��V�:�{�ƫQ>��'�~���~���hݯ�k'�h�H$�y�~��>�׌�u+������4p�}�$W�]�i��﫩^雚&ei�����|mS6�N���h����jw/^q[Fey)앑����~�[�	�s�1>�ɸ��ٴ������ZC��`���*�uv p�˝�w�q�1dǛ��Ț��(�w.��gX��c�-{c���9y��̬�.��i����
Υ������Ӏd�r4G?��/�(�D�h�^ԅO7me�R�,l[��^%'~1�x�7T��-�+����E�T���ݽ`�b�yW�[F�Xt�d��5�����S�Q輭�6�����	�U��kw�Y���~���ѭpn��o"ھxGM꛽V�wvJ�V*ig�If�4P�M#�<���J��6f��[�����E
�k�֕���r��݄��in���Qp��S��j�_K9}��,���u���!�c�P�\���eo[�^_b���&s9�s��c�n�f�e7��a�Tz�����sz-�/'5u�����]jwt4̢.�L�z��T|���~j4D4U�Z�jop���j�g[�T�skFX�����t���b�$�޻ڄ��-TjVL��)˟f�Vi��cpVg=7���n�j��u�UH#��/�u5�u_f�neKə�ҝ��AϬ��;ջ@��r��s�ou�Ż҅ޥwJ�k�Ĭ��xQP��@���<�0�M��o0����@��mT���w1f�\r���r�_M��'/vV�fx�̏p�OB�]z?fa��N��Bf�]�`���Kn�̔��FT����[x��8����a��<՚)c�����k �ʽ�9ؽ�8,����
��+?z�,r ����g���j�}���5�T.v�ѕA� �k3��0�Fx�=�*)���_-W�Za��
qy�7��!*�8�8�׹w�Z�N�����5����}�/�S�iٳ��h)��0�-����u�^7���xQ�����Zx����o|&���}�N�S�����T�f7/��^���|��+��̻h���3�<sh��A��/&8|�����p��<�vnu��cH�����6�����ƛL�^{Ϛ�6��������FmX��'�/R�]������ُۢH1�5g��ޕ/7k( 4{��x���n�y�7_{eޕ��뺅c�ݺ�m�W�Ԋ�
����yLfvr +c���뽤����Tt$�"V|�ho�G󆹋�U�u���{����֞�+s��}�����ex��Č���ci�Hd��.Wn�s<�i��ӗ��h�i���Tv;�(�G��i_]�(�#�-��m��;ɏ*pi�N��;�%��xZf������B\�l��Ŝ��qZ*�lд�g:���k]�X�5J��l�M��+t�O������D��O'S�s��hYԯNǦ� �*�]!���32_H�+2��fKhjlE�� ���S��o2��ۧ�n���H*������Ʌ�]V�:EW�+p�W����5!cY�].�q���gb�HU�_A��Q��'O�$�;RmZ���v˝m�-��r"�]n�`�#��^�2�
딦����U��dJj�3Ⓣm'����"��N��J�{S����4��f-�G��W;�u�{��V ;�0��C�9�����Y�� &
�l�|�I$h�5�r�OZ�Ԕ���x]=�kyR�34�9H�\��b����bLu���u�.(����/
����A ��I�����Y�+����������n;�g��B���2נ��e^y�!��CW�|4;��cV�լ�og���W�ޡ���k��ۿ�Qc�]2��` �r��l6]�u��p��We�t8�=����Q�W�߹��}�tG��� �f��䰇W��`RM���M��WR�qH�����PW��t�]�ҮJ��ϻ
�T.�ǝe�{p�Ca��X��9�	G�Z C��A��gsU � ��I��P� �kz��^ev"	��'t����Pp���({�`��-�
o�mJ�h�^^�s'���dUv��.w���m���X�{n��&�]u��k��g�)�<�uRgn�e�ZmYFzn�]�y��\<��� ���'�v���%/T��ն8����oU�.��]�Þ��d.4H��nu�����c�ul���v���\]%�ޫ�I�m�-O>�KԎ15Z��̋<��ݬbt
��O=k�;z�mj��nz��-ƣ�;//oJe{gV�ڵ��:�	�Cn<��m��Y����Z�v���{7)�l~b��"V,X6X�������w+�;��/y�
R:N������\���䲂϶�� ��� i]M���ˉ��u[�Fn[C�{�q�1�79�>��v ��<x��M^����ֳ��O����ZU���9jsa�%���;��+%ž`r��k�ń�mX��tǓ�.~�-�w{us�?=y�o��l�_�����PuN��"��6�)A�d|���ݳKڮ�H;Q^j� �h�m��ê�;X{vN�~�IwW��7��>�C�4G�s��|آ)��1[�f��!okի˥a�>�k�4�3�gR����%��"�
P���΋M!�o��M>Ow�ڧ�2��\������C��Lr�b�}�O,��1[֫���^���I�����h��1ιu��A�eɐW�=h�29騼����ܝ�X��6̽v�փ�U��T��=�#(!������8o�1ر��(��K1
��7w�78
c����װ�ok�ǤU胡�8w��VF�-�E��]���r��!':���0�'�nS�+cH��X����/#�!���c����;A9QVW_t��{1!�����R�k��[:d�����/��;�3�l�,>t;���>���v�IaW��^
�tO��ٔ�O-�r�]�r�J�(�lt�q���������li��\I�a����r�>L�`۝�
���y����6Y}d��h��D�k0�n��B*K�]*8�їw��t[�b¤���X�\ꜙܢ�c��XZ�҅g,깼�Տf��I��l_W}�R)�.�
)4���OJaofa�䆵H���m��L�2��E
�}�ةZKgc�2�/�f�Z�ۏ�ͥ~��:W6�n���ݡ7�ݶ�H-���v���m���(�2W�n'\� &ʿ�x�̔��������������:�x�'1q�k�P]���wq��ft�e+2ܾ5㫸���W��5 iS!2�n����d�Pm�����<�U�%��\�=�EC�|��>�h|��M�4:_���<7s�.��f(��'չ����	�-*@��D�OQ����l1 Xஒ{C�|;'טWέuidjx͆Pȯ���q͵���6H4G��
���X{{��!�W�+^�!�FiZ�1FW�<����`W�hNQl>�c+�x����hk��*��A6Z@Q� i����
�4��/m��<g9�ǣ
qC4��<�Owi5Iszׯ����=����X67����+�|�ӓ/2^/��p"�| !�XAm]\��^����)�X��'���{vvZ@xvi�i+]�U��
^���� ��F7�s�/׎9�^��G��ׇ�vv�w�k�Z^C��N��gg�jU[N5eR�}hP�Ƥ	��Q�ǂxR��_F..l6��z�[G�=e뤺�l/���6�w>ܡaL�L�<�gnX�bծp��L��(; �����`�2bY):����<w6iG�'7��G��R?U��Xus�1��p:��a�.������n+�F�&�
��uB�_y�"��)vw����m������r�Cӂ�,m{��9�d���ד^�Û�շ��|r}��%��g'�`����$�,uy��Cj��ڕx�TPE�koZF�N{Z��X���� �ں0J#v�uM�ؐ����y�<1��R����W�K%e9Zj����76�r�?1�� mv��J�cQ>ވ�Oe9��������]]	�,���� L_rV��r��R��4�ўS��ָwpo���X�v%����Ne��8��:�40X�׶�������ER@�L�V���JʬhI��ss�sx�k���{[x�^�ױ�����wOV4t̿�=�\��cm��.�0�h艧���<�j�\W���~z]N�T�/��|&c�HT�!h�[v�j�������\���OK[��^�fj�9��q'|��x�:�F��r�-NxWQ�4�b�M㲇�Z�V'�Kw��mb,�g�n���:�wm@�$�+=�3�#��{7�{��'n��)�:��f]/+լ�v�VБĎ����m;fK��xW!�?^7'Z�Ľ��V���2^VR�P���w����w�鄹!G�i�	A�ѩ�7�g%y|��{(�^:��*�4�
�c'Eo��a捹(�G�o'i�e:����WP�q��Rq��SF3�V.�5��r�)����L�7�use�e;��焎J�;�� ���bP-إC��;gN��Bau��h�����oD#�{����G���fɟv��g�q�ru��tp�δ�`W���S�:Ƭ,����>8�\�5���y��#v�@f�ٺ�=u�슔u7)gn��}��k���_l=0q���zsn������v��hܾY�M��ǈyݶ�Υ7g�;�8���#�+���Ξ�ps�L�z���'�����ȧV�/Y���:q�n]Da+k��k�w�r۞ހӸ�S��+�������s<qf������"�~6G^Z6u�#yzx��r��[�g�>;���k��>I�&�� *B�e?�!�cc�o)���d�g6B�)�m�W���ۈt=�ռ��/嗓۪�RKǀ;��e�/�2�Wr���ܢV��H�Xm�^��z��t�^6,T"�d��v��G��Adu�Sf+�2vIH��+�K�8�	ne���YT�D$�d��_%Cu�mfm����ztOb�gcS?G����¼5i��x&kE}Su���ל�m{u^½�R�M�K��Z-���`	;�y��*��/���YQ�.�V��i"��ʣ��xk��6"��/(�
Yueh6�����@�v��ܽx{�,���"`���$ۘ�ݹ����t��	D���ky��N]{��7�<)�s��!O���8ڞ�>��n��Ì.FL���֋��r���i�(�Ej�o'�[�c�y���a^��-��]�H��	[�V��h��ut)/ӣnf�g:��!�vu��1��!�L�܈T��N�.�� �딤H5he��Jl�6���|��(E�˙�u�j^G�!ms�z*!ʶ�G�X�O
�.���h��t�e�I*H��n ҚN�g[�^ӥ�x�y��Trp��B���h��+^y��I:׶H3[yf��\�RTe�$�Km���d�����[��x�r6+ȷޔ��6�u�G��g��R�h�g���n�$ƪ:Ƒ���O��@F��5>
45R���3��˖"�w�pQ�n*�_�jt��~\��z_b�7u��L^1�W��3�K� �i�wZyt�A�u[e�81�q�x���N�������b+$*�sG�n�;�F،j�n{�Z|�`�VWY|}��#iV����{ew�[��^�^f��3��4�d&�h����;+�kG�� 2�vn� z6�W�>�!�ד��c<��oS�h���;����rh���7�&��Lr"A���;9����x��n��F��̠��<��\�mmC���_.�Ciqxt|�w�՜�j{�wٱ�\�n����T�}���M�Wp�[���M��B�\��1��oy���D{�)��.��D�|�@m]�U�)tia+�zғ:j����dyz�{��U�-3��m1
�b���*K,-(�1��fݞ���W ��m2��oi���w��okۦ�f���2>�S(�ɬv�J�:��=ã�f��`l�ᶩ)�	z�ozU��Ǯ��M�����m7���ip��ʭ�hNA(�v��u�gs�AY:�m�`�L�Q- ���SuSV�=͏������7{95��<�{s;|�	TJ�}	�V��z�L$�'�����J�I�`r�]-;9��Z.�{|�s����0P~�}MK���EZ�1k7���eu�
qٝsï��=AP[�ER$)��)�Yu|�jbU-�Dj�6����醦�v)e�H�櫛��&�<�����	QT� ����<�5m�72v�u�a�Z{X��j�t�]���:7p?QU��O��i���u��T����w{v,�oD�"J!������,�jժ��ǘ��{ވը���5ot��ɔ�~�/+X�$+e��*Q�(����̝��=z��\	�VM���\�稒ph'\ft��{�Z��U��nM�mv��v7��eㇴY�ٹ��l\�'Bk�kүSn�8S���{�<�Nۥ���h`9y��&oP�s�����x�p�+-C�]�I��5�sp�c{%"�+��m,l�
j+ �gyΛ�7[g�t�'m�4v��x�_n�1.z����Td5A4���K�f�m=�y0Q��(����aF�M��$ݏsEx�+�o���� D"�{v%��k�hf�^��ȭX�D�{�YT)�K�����1�^ߗ�iű����2��r�gb!:vX|+Z�[�f���v�VԸ�R�墹`��t¶�f\S-WAim-
Gl���V��λ�4�"��xZ6�T���+Q-�6m 0	�Az�Z�54�_����諭����I I?� I I?�$�$�	$	'� �@�x����$�$������HO��I I/� $�$��II�	$	% I I. I I?���� �@�`	$	'��I I?�	$	'�$�$�II�f(+$�k"줏�׻� �������c�X�  � �a�U3e_;�9)φ=+�ݺP/�<W��hP}�u:S�>�fiV���2SCF��'9VmUn�@��fԦN�nܩ͔4n���   ")�@RJ� � 0M2h�����BU"0L� 44�����=UT��      ��5R��F�d24 j�*J�  0 ��
RBA�O#F���)���z����9���AY���"��$�+���2�V�f�[��Y��8�af�2�M����K)QZb��d(�2�{l�f;��7�Y�6�@V���?��i��[ο+^6=:͚�r���kOK�]�q��r��q��ܖZ�S��$�� ��6�q��Z*Q�Ǝ=}AR��uu�t;v�0��OF+�����n��ͺ;����%^��L��Qˬ��0.�,oNd��͕�bZ�.��4�8IG9�6�	M��F�t⎟u�ӶH��h�.�,ExE�óGJ�Xh7����N�Yk.�Y�.�n���/��;	�����F���b�:--5x)���6l59�CM����)�mچ�K��\lHC�qJQH�yٗ���Gs{�R�%1�9�>��ge"���L'�$XLkt� R�W%� ��v4��y�T���G+��ozt�@:_[V�м�֯/�ֶxgK��Z�7�q{ ��?l��?M�,��	��B|���N���_��=fs�#��3�x��ٸ�i�(                                                  ��(               �                                                           n�L��ٻ�D���Ck����ͪ#�(Sh�[f5I��.-����L]LY.�' <�������6�ԍ���ܖ����9��M%�A�J��m%��-[����L�С@��X`���ٙ�M.�J�j$����i���\kl),\���Yl�,�M z��Z�M7i���6�R��6������`SV`������̹�gI�5��5]3�X�k(���\;Z�l�	��v����.R�Mu�$='�K�׭r��$+�9ulPU��}]��}���K���5@VeX������e,䜜�w��}7�����       (P  -�           .ջW%�QKx�@Rk8��ja����̭(�5���0E]�Isn�ڡ)n��rNs�����  -� �smں�	�8>xZi(	L��2������.L��o���Nn����pO%�Oy^I0�m�Feovg���^��{Tkm�&o�]A�L��Hբ��K���8c�P��W�ox���N�m6�۰��M'm��LW�&�ySϸ�ἒFҴJ����zj�����X������qǜW�6q�>��    I�/8�fl[k$��M�Nw���K�n���<��Hє�,�3L�:��sI �$,��U�q���p�=���N��rdz��Q�H��%�������l�77&�f�U�x�W��\I�L<<(ӷ�ʹ�ټ��ث�bg8�8Y������ލ�L�Ps���\KaNr��y��bn��}��)��/U��z���=�;���s� �!�  ���#u��ݵ�t��t���{�Cꢐ�}�ɴ
g��՗�Y����6�T��f�����x�3Z��̺���ܤ-Nw��S�s;�{N�n�����&�3hWjX�P�*�����֐��U�s0�o��(m�{�"<��ŏ���wW��:ؕ�g�
o�u�:��.�F��~|ظ�|�k���8�0��ߏ�q����_fe����.$^��&���)���k�*͡�b���|8|�B�r�����.��#��m�2�)��x�SH{��t�Q/^�ҽ���l1��X�2�wt�s�[a�{ܝ���`    �2���J
��g9��)�E�"����"�k����lE�E�C|��"�"�ff"��H��,�]��*m��x��{�������dW���T�F��jAJN>{��Z�
��Ka[��߽���g>��߼�N������.��S>��1�vm;�/!�$NN��{�Uu�שܓ��Pz�k����XfP���֘�Ux��w�qμ��F��]s(��RO7�f����ͬ����p<y�ת��S�+&���u'/W;w�˔�K�?F~[�������Ϫ�C���=�Ə.�G�>��ځW�y�PGl*�������i9tL`������Up㷍�N�����|��    Y�,�S1�RS���p��$��go��	�{�`u-��통E-V:LC}�z�儉��#���B �3����˼3\`�c^�Hc�����oiI�N}�Y4���뤮�OY�y�<E�<����[jm�+��b��������u��{qʆ:����S�ǾW��q���||JI㼳�y���*�+g����}�bk���Ղ��������)=~̽%��u��M�)��y}�˼ˬ��(f�p�=�i>g'i���L��=�c8�\�k��q)
M�`�P"!����R���L�	�S��k�{�u�����q�{����w{�5�I                        �A����8u��Y�بR])F�%%�@f)�:�ƺ78�ٱ%[j[B��^��,���    ��wnUuظu���U�ٚ��%9�͕_���mLi�C���6��P�=��$�L;˿9P�)�AH) � RC~߷v՛ˣd�����R
AH,
�ZOP��$���D�S&]S�(ٿ~54�R
AI�(H)�R
C�Yd���N2k������L��L�yS� ����A`[I �8�AH)
�XaIIL
H)�e���R
A�8��������U��ͳ9�9r ���$$�N2� �2/��XAH)+t� �CuD��,��a��$�3l��Y���_{��ͤ��Y)�����Q&���AH) ���P@�HOXy��a3�U\�30f32����������x^ ���FM��`RAHm���R
AI樖�e�L��Z�̦��f&bf&b,Hk�� �AH)�Y�����R ��)���&$AH) ���X>gפ�����3��^y����9�|&�����:W�KB�ʸS�3�eTuB D1�V� G�=Zd���׭��m�  ɖfȚԒL���C*�k�fz��y<�N�o>4�;Z�{TRi����Ǿ�8���w/m��\.no\�@��;��8���!�iO^U�{�.[��N�/>�3�PS��m�}���.�u��Q�j��G�<�(D�"&��)�ױ%��9W�i�������F�Uי�ffcwy�Z"ɾ{�&��;��{�ޤ!آ�1��CN3.X9u��מj6	��}��x�c-�|�'�u�e5�@S��z�Y��y۲(f��-�x�ɾ���ߎ����ߝ�   Kv_W&���Q-�l����0R����4���YI�i4¼�oɌ=I��~1N�J�c9�k331����s��C���K��a�~4bu�<k߬7�񞤷��xLv�^V�߲��A�)~g��3/*����\����)���7s}�;�f[����?f,�2T��f���t֮��8^�ͨ��z�>8{��P�SN=�,O��m��U�����;�P}m�V})���K���m�J!����j�O0 >)A�d��<|g@K%h�~��O$�   .����jpJj2�m�h%W>�yTq�`Z��\�1�>&{m�m��i�b���n��C��T�s�u5`��X��:�Hb1��P���£-L	v��9c8vq�d�`���ϒIZ%J��v���ffo�5%e+��U%xm�x�EX(Z�X�=M�1ĆI�:���vC/�}��:޻�:��g    6��g���T
d���lJ�F�˞lpÎXR�K�T��Æ�/�7sL؛�Pz��3Wng(u]���C~��^���I[`�e�u#�Bro\����1����'z��<��mAm�T�oL�X6v޾��.�	�eY�R��>I!aR(K������<0�a�WU��t����ަ��f��a�:!��c����y��w�Z8�N��yӞ��f޼�-�                         ���wm��+�����6�؛
Ɗ]mn+�M���HV�ە��4u��6��6���s���^�����   Y7kR�)b*Z6@U]o�k�e�|'���鯆�4n0�����.{����I��.Fomb�5Sg��r�JG���)X�ɞI$���Ļ�;�|
��%9��=������9��O�֗rI�H�]3ą'��.�Q�/Ηi�MO$~yܠ篩��6�O�k[��w75�'�EUs:�d�����������    OVT�fٚn6��h"�E{�{��90Cy��J����q�N���57��M�3r�ug^Lv�' PE�n�ۋuTV)IB��cm@H5�V���9	��YpkFʍ�wwm��[��u������:���Pw_��f��)�oG;�Ǔ�g�lÄ�d\�ё\�gE���]@\a��SW�ǝ�u��u�f䳯    r.�ݛq"������mS��d1[�n�q�ƳY��r�U+}Ch{Qt;��m��m"��Z
�Ӱ��1W&��-n ɼ˘�3\�p�m��TH���gi�GOW���-{��YV����+!Bd_@�Lkˍ��(]8Ø˫[�Pa\tH��G���p���A��,�U����m�f)O���6����a��n	��w�p`�W�C�NﭴCL�oQ�uﺮ|�.t)�f��J�����"�cm��  6�K�YuQ�(2�%��h�R��DlZx�z���Sb�צ�P(��sm��+l�kx��"���҄��;<J���>I.s7���e�U���t��e��
���1^�'��������IE*�M��,�۬������.s����{آ�z��ڀ�	�]㧡O'��8�i�׌�>NP�fz����*��ڦ�m�   l�g�D��Li���m�)�K�Ƕ�=�ʰ��MP���Õ�ݏ=]>�t��RM�p#=>��TTE�^�ܹ�w�wY��	��sm2<�u3Y�\&��l������X��ԑ@IJ�r��1%ű�d�ڮ��MF��
���8��5J��:�}�[eA��}*��s���z�0L
|9��$�!���ɞ����p2q{�ЩXz`�6񌁗9��Wg�u��g��9�]��{��                        �nc,�K���Ir<��0h+�v ��U��ʀ��s�-�*���vK�n�y���    ݶ�m�+.F���ʭ��l�)�g�ۚ�V�O�w;{�;�ew�O˥�k[h�P��qxdo*��g![�/s`!��l���"�ɺ+���$���\�o�b3�A(݃����,�77Ֆ�l����o{��\�x������5TܫH+���<<驴l�n��x��rn9�qѵ�y�'��x�ϝ{�Ì޸_7ە    n�f.��7L��Q"(YO7|ۻ��m7f��ϝ�NRmq�m��,�b���9@�j۪��=/p�y�{+�g�Al��I`��yl���r]NL���k��1��Kv�<�����"�V��=��&��):�j)�qBa��1���l��qG4�7��쎽�Ӥ2�y/��9�x���}��    l\���M34rW*̵��;v��W�q�Z��2���1~���F�l��&3�d9qϺA�άm��Ï#9�n�-��I�UX��f���a@�91��keO\���|6���X�*�45�g5e�:��M�Â��O�	g�R��#=��~�m�����,�{���1Ȇ�ɹO�h�7>��T!�[�鶚)�3�^n���׽٘xY�Ю���u�\[�{�m��m�  ]ۭ���Զ�	T�
�S=�ؒ�X��d��j��d�$�ul��m�Yh'�y�\=�P��s"T���U+-K�̛�Ҿđ�0��t���L�y�Į�;!�g�t��y�J5��%D ��Y�K�T��+��w3f$F��v�N��g*�Ͷ�i��y7MP#o����L�one�6+R:�d�(�oS���    ە���Mn�+Jl,Ny����͛�L�)b̮���wcm [�K�&&u.��VՐ}��<� �q99'��+y��60��lr�k�Z�|�4
��iw/+�r�V�o�3�4(I��.A�7ᣱd�x���sL����!&ATj��"�	|{����i{CT=ȋ�\I>*R�BvIy�����+3�V0�x%��Ǚ�;����z�8�RN/`                        +R]۬�efC8ɫ�6£�.nt�	�KR�һ��*pytQ�]�&V��\ee���    �2nQ��i%�m��H�vq���zgQa�J��y6y��,����H%I+9�6���I�6܁e�<F�N�tK���i#H�D&R���{;x���q⸻6/gVH���(5��z?$��o�����泓����(�������.|� ������׭���}N�&
6W{�6o�8�    k��8ȴveW:�7�󻤻��;�$�{0�Ysvo��.��i�ʹ�S����0���]�s̉�uj�b�L���E[m�a��ev�+����{�%Fw�9w��f�悲�MGV��� �K��"�n!.9f�d�!>�ha��*AR6�I�ޤf�0du��� Nlo)m�ަ�v��    ��Ha3h�*z������Ź����Vt��Z�ݣǦbmhi�ST'���-�gv��f����I�9�rfe�����Gp(�đ�U�����ܷ#ϡ� ���I���
9MM\�cx�v�:;xiI��wC�H�i,7*f�e�^T/}�m�N& �z2�I*(�V�qU�*1dLc�|r�p���a&����c�é#h%j�Z���3bW�`�������u�ý-$�   VL�$@�(�%RH�I�j��l��Rq=q�\��f��]�IM�.T/5͆dm�l���s�^�m<(|�|�P�L:u�F�{r��(R��"w���ُRI$m%`��j8����m��8̹�vL�9mn��J�*�A��K��@��8Vn�� ��:�wvo1&��\�   �Z�FZ.f��]�Pr��U�������%%�-q��Ќ�Z�D U#3�r��Q��J:�{�S.��܏	�K����i%`��q��Έii�yK�;Rms��IY
�����Ùl�o'm����,w|]m��C��$@) @��V���{��37�f������6+�"�(����X��{C��/���|>��p[©��Zm�� +�,���ӑ���v�m�-��n���U��ME��-:���p5�y�3�V��O��Sn���덲�q�,-�6�'6�vr-�n�V�:Z[�~R�tz�}^/�/M���+�C�@��/:X^{�������1�e������/D������>�/�,�\Q��}z,ut%�7��KE���ظ�'2�}Z��Zu۽��ff�9yg�?�9��@԰����
�yi'"ڽ�c�n�z��>��k�����15�\������K�:˙v�P��?�ɿ��
��?~c��M�<c(
��-3�����@�z���<[����/���>��NJ~E�^�������x�+��Y����=��GAp_�� �vA�/*���_4�5q~,�a��&��~�NJʧcj� �j�C�Ȓq�̱�-��~�s�R+Jm�йq�ln����{��.��Ծ�t�^�gB\��z�OMS��v������z�����v��r����_�:��_}�{j�ϙ�@W��[��_���K���x��u�m��X3#��U�����?�OGꞟSV�k����]��<�tw����\�OgIv��������izս.�w1Y@W��cg�-�����{����5�z=�~��Z��:1���K�#���]��B@����