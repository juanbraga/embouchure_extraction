BZh91AY&SY,��˝߀`p���2� ����a��3�"*
!��T�UT|-F�P�f�4$P��-�T�bJ
��+F���IIP��ReL؊����)@@TI*A@ U	�IPPm�%P
�D�*UE$*@��IT)$�#A�*����ER�J���j��Q��ch��靛�����3j`�E���q�;k�ͣ��r��U�5f�E4����@(��qq�Slۗ\`[��Ɖ��4���%�n8��GG\�-vI��F,\f�m8�CY*�����s�R��ـ �Tl� �UEn�������ˮ;u��Trd\�:�c��`5�۫s�)%p�v����v6,���;�ð�[����-5v�E9�l�T����R��Z����'.��Q������`�[�v8��5;smúv�6P�`ܳ�rk�ۍ��	a������6���@�Q�f�8�;�8�V���Y;��t�vj��wV�������,�i�,3i˝;�qڮmZܵV�n�M�������H�JP��9��X��4l�K������`�d\�8v�7n۷4殻�.���m��i�*6�����Q��r뻡f1Ҏ�օ%��"[��Y��\���q�Ӊ�]]��w6��[�kq�8�F\q\!�sR�q�c��dn���v�nͮ��;q��ݭH��&�`*�*�T%L��.T��9�:�p��U���rj��K�ӭ��wG9iLAwK[�se6�lu0���v�a�.�k�ݕ۪%�YaJJ
��\ήwm�qŎ����g�k;s�I;U�	�`b��eò�T�)��3nf
�6ۮ;gs�+�VZ�e*H�W[5�\즢�s�ε� ������9�!��2�1�l��v�\���j볫��k�6�z� S�)J�CC@#F��O�bJR�0     )Mhhj{S$�@�PڃT� JR�0     )��L�04�L�4	5	J��     nٻ���n�h��iR��+|
dW,/z�L'(�+l"�e5�&�DQV�j�
�*ʪ�*������EZ/tDQV?zEEZ�x�(�����U���Jp�:R����8�𙙼R�zWK'��
n��Kq3.��+k2��lPd(�BN�yb�b��K��/r�TM�*ˬ��DU�yB�����F5D�VJ��Z���J7��1*JCz���1����0�ku��l溒�I�/�d�d7��Q�g+R�A�]��41[�c�V�b��47&�PQ�x�/i�hLݠ�*��!H",-�!o��o�u��r�Ub��ǚ���bX.���L��U��߰��E|A�n��ӥ�1Ҋ�nC6C���e�anڽ�K�[V��,\�h�L�w�n|���s��+p9�"�WpV��xc;��m����Ӎmm=�L���3y��H��	���C6���� Z5�Ø@A����	�h�oX*�K�Xi���7pM��ʥ\WM�.��6κoo쥶�qG*� ���^���Fm�T�ӪUXb@튛H���U���A{���VL�!�y�Rn�˦��7�:v�^�B�YX��d*�<4��[)kvn}&U�˕b險�����{n��hmॵ��kD�ş!Ki3)�-��x)��:FF�y�(+�W�Q̲�4���r�
 +TI�6̹A�h�k	Z�X@͙�彭�i�T�?��6���T``�6:F�U��0e�)SM�{�7 ��5��IE��Y(�J�Wmd
��[u6�U��r��ő�ٚ�P���r��a�/C.�3*^�ǎLI�[� ��;��༊��E��A]���U�[�d���wi{W�<1�{W3�F�u��t�Mڏ���-댟�����Fh94�oF���Bs�o너��z�N�+��nX�vTEɇq.f�rlWr�f��p�v-Sw���sN�JP5�!���Q\��RU���"	`���#�4�U�݉�dP���PV�b�En�I^��+Z$�Ы[���.��F&q)ae,�$��uZ��y�Mչ��n,/.km�y����F�Rۋ6̙(Gy��g\� ��n˻J�̅꣕`d���7�G�yQ�w!����FZ�R�t�]Gt�c����j��r������l�F�.��0�sb��x��`��6#� ����)ar�\;b�R���Y�ڀ��֩��7q�յ�����%�fd��:�.����We�V,��AǢi��+���P�q�m��i�O$�FJ�)a�կ$9@<K��ɤ�L�X:�e�5�٨���^D�3wc�2���C���KNe桔���\y)f���Y��v�`U4�m�[N^)�zv�c��{�f8	"�k���¤*m�(l҂:����C
2�v�0���.c%0~�;v�[N4�ОDA#65��[��J2�M�J����st�z�^�͠����!�`�[����J�CW��Y����`��r^�Z��0�xM�C^!x��Yb��ݖ�ХH����9`�,X���@���rŘ��LZwSܲ�W@� �j	�T^=&V<����h��b�����H��v�cKZ�U)�]�i�K5�	�O*���XT$`��v����s:ګ-CT��7Xɀ�t���32iyi	P(XT7q��c��CrFhۊ�4� ���բ1Xہ�f�,YdhhM��*,ӭ�J[�7 ��)�E-� ˦�v�!�����mV��Avi��q�)���LwN,�E��2��F��3wS";wX�mPԥ�V��N��c�3�rM�m��>�yJ��*���t&hn܁kJ⽙M�F�jl�[Y�z���W�w`i�%�,EV�Sͅ��b׸�ɗV�\#M�M�j5T2i��@� ��rC0�p�;�tBM̛�5�8����s5��j�[یl�(��t(#∬�[h-Q��!��B��6��j@�7.��6-���g_����yZ��jCj����nH�FU����E���ť������R�%�zr��;�Tk1�V�oZ�@-I�ԉ�+j���sn�Ց�P��ܪ،�YL�`�����X�F7PR�,�G�j؀M)^Db�NhJtelELU9Q��:��A3�͔aTT\5�l��P,2�A`�Ӵ)PD��M!J�����`c�X�娈b�p��f��f�DE�B����s�Ί�8�[kYUw�7� ����1m��I�	��kN+���N���|w�̼(��0QF#�,e��������c"������n����PѪ��ާ��'�6hYX�s�(@�(,%+7?|�;7)hOjiw�B��yvbU�#2���2��~%�M��i
dZSl�5$�r���mv��pl�+&�tV��=ρ�P�6lA �` W�,��ә㋼����NpS�	��Q�a��L"�.@*�%k�j1�!��v��!�(0���A �#�hF��@�H6��[��Y�QG5�0S�.�lR��R�M�h��*Bmh�Fhѡ��5�j�#nLv�����=ɭ��ǁI�d�,�9u�h���a��h�6cN;r3h�W��h���#�赪�]�f65;۠@ҭ��ӑA�iK؎�m=t���onS�Xb�k1C�K+j��(U��7c����~#+m,�Ok�@F$�EI!�;	�逳�#��U0D���0ت4��b�`��*�;ţ�e�i�Z�AZnEx�B�ݬ��W�@�R��3n�l�*[�^�҃5R.- �&�a(]
آ�����bdQډ7#w��< ��0X��DU�PH-0)����IH�R(/R�i�"�����l�
�0��Aj6�t��u�Q��]Ֆ�q�qdD�v��j�|)�*��̷�����z�ie;*�^�-@ވ�͕p��W[J`��]3b��E0Ұ���y�QNn�5p�wO�$����,ςw��F�m�����Ыy�Z1�cX20���,
i�)DU,�YʡL)4���`ky.e
dë�H�H�W|�2�Tt�
:�F!���t�T���H�H(p�vX��K�4S�{AĠ$�Y�-��!Q
�ʷ����T��$QD��qY��07D~�~�1�\o%"�I��j	Zݱa���vn��a�sN�ܬ�͊�D��$��+�0TJ�x��ܔ���he;[��Ԋ�eiǦ4*���̙/	�up3�`u�1Qb��hI���J�FSw��9t�V�A�(S-e��t�Ee�pb��	Y��B���ܶ��zS"Ad����ֻ�vo�M�T�ևT��a�
�� �����Qp黫ԍ9�7�Ì�$P�@!�]�ĶAIޭȵ��GԢ�嚟(�B��>8�#�U@A�̂aQl�Ϫ��b�GN�ŷY��0�؛�ԓv�ԡz��4R�;Y�����0S#kT���	�f�h��HYn�l���6e"S��$���.6�-�M5��j�� T?��X�ɴ����SV��ئ�d��ҕM�y����`���ݢw�N�+iit�G��Tђ�c�bd���]�0�L��v/u��
D���.^h��e�/p<y�X�E���1�+l���JQ�nʓr��[B���I(�*�;yre�$�a���٧Z�ZZ�`ٵX
�X5d+A�q��J�,����cm�e�K"*l�J��v��D�	\��7w[���$ƣM�qR�d��NeYd����CS�!�^��")�î�^���VG-���ccUw2S&�V�B���m�)���	��S@;���h���):�q��^�؞[�w�O��>�<g�'\��.-�Y)�����͡zE[pf*BR��Mn	�4��t��l�!���]�B�8��sS�`X,"��-A �`�S	H���QE��ѕ��g5�]]'m(R0+:dV��B�ںM
�2֗l�8�j�e܆S��B�[ʕ(�ڰ-�o`ut�4�w���c�qАTi�h���8!"�� ��1�K�B�a�v�M���>V��2��� 9Vn���@�� �&���ۖe�N�F�۱p�l�
���i:��ok[ʡ5���Ɋ£�Q��Ӎ`��er�ڵ.-�HWU�99���q�3-*,�ՠ�-"���(7E�7v&��W���BkZŹ�R�K�Xh� &樅J˼�֚i���W��&�2bw�4�%n�qXո��;���7�x&�+%��h]ik*�1��V;S�G� An�)P�XB
�%�
��:��d$�ZV�Y0|�%�Pn�U��@˗PSG�-֜Tr���}@W�}�lPͲ��I���Jomը�TX�t:�AaN�(J5��
L�7��ZbEd�X@��]���1��� �c5�1c٣)lʹ��񼩉�x0*��K,�o)X���'�~�����LCF�!w��V��IE�T�5C�dL`���.��^���	vv�	�eJ�-H�fU��k�][�L���g�U��(U���j��rdfKy˨̠�A�t�\,��<�(hK�lU�/Y�hk ��OSHm��6/Ķ��P��}N�(�ͻ{Kb��V�a�K�f:؈z�A�pkF�����6���
ᨉ̎�Z��Tj+���(�,T�{v`a�/n��OM���wU@�6��d��bG/r�#J��`�]K�{h�X�V�e!x�>)%�8JD�2�h��i�u��D환�G2�L���֦�����fJ��aݠ�@ Ԧ��b�̏�]�HV��%��*d�1���N�ڱx��F�^Q�l���V�n���ǉU�p�����&s[��j�81ލ��Z�;-T/�)�he��rKl���,bWa^�
�lӦ%,:�Rü�ۤ�d[5�9,Vl�b��3�Zq5x>�-鹟;j���m.�P��i�ް:�P�n�o��/c3����R���Յ0���4�Օ"��K2���|4�"�;[�(n�qBu$�V��nޖ�B�d`5���6�6wk~�op�-J�WB���m��ۥDnT��gjC�Xz�z^��૶��̖u
Zg�ab[d̄�oH�S���#v�kr���:�$V�С4�"�s�g���$�@��w7J���T-Z�7bRIJ� ����͙�\�̥�93A̺y�S0k�kh�Y�p5AԷ���8l(�1Q%n����(��Y��ڊ�P��E�RJ�{�}!��}�M�td�.�j�@�J�8%�� Ai<�s6��[6˂f�
 �+F��5���\�Oh�Y_;7.�f���.�o7N�"�Gf��K:��W�!-��×N�Gl���3�,��.�љ��R�Z���ε��r�Ʒ�:۬J��A4~D��m�!e�U
ЙT�m�B[�r��֪`�R���4�ũj&�p�G5��Ҟ&�`"�K�)�/]j�H{�	�$$*_̜�� �u�u`�+,���i�
��ޤ�[U�mЃ�4�$��QD�+�4ۢ.,Q�Y,V�dU��J�����e\D,�(�@4���"bl���,X Ux	$ <6XO��7�@��;x���X�3V�75ZN�b����G2�EHn�	[7��m����-옍��#��%�J����S��ƽ
�P�F�4&�5�#��b[uX��w bM���z��(�Sj�0UX[������d�閾�dJ��Y��
V�ӭ��aܽ�ulXuh]�Q��cf��I�9FV*y�Ģ�.�D��Q��)t�â�Z�rl������T��*��'�EbD�j��I2ҩ@ ,$��)H�L��mM��tl1��ۭWp��z��x��mM���ca�"6UA���(X�S���Z��*dsi�+s�k�r���)��-�/J�ɏ$�D1��B��p�	(��㽌,�uQ[���Q,ȢM��*�����3R�gXUmTVE
�^"��KR �DVŅ�����X���-!{&*d�Aq���f��t*V�G�/(�e�ٕ�w�2\�Lm�S@���%�؃O��?�T��j�Cq�ħ7N����P*f\z6�QdU�	R�x�-�S:��5�����(i�:6��b�ϑ�~ a0P���VnQhl�(![{����K�����I�����n�*&�m�):��z�:h飙F����F��XE=��ԯ��F-m�As���6�B����ݸY�9[%��aR�k���(с5U	��Z)��tm5�O�]�x���	$f��9*�d��cM ���j�W�cu\źr�����j��Y�â\9��F�֋1a��Jc�����˽Y.�`��Fm���(kW�z1�-�EJg\���j&�6.b1��;�,@�yb�x�)��l��r��,b�/v
�Rҧ5�kkpej�J��V�F��K�;Kq�%QSUC����L]����u����t@����b@��m�iP���u��
_niS�SF�W�jX6�A^%����l�����b5Q��-d�)��Y�d-J�t*�6م���	���+��[���C,���������

�v���vJ�߮��4.O��U��_k݄��-��kr�wjS�yB�S�;ݹV?�!�]M&L�ٶ���v�� \��ù��yW�l�7w0HF�z�Mk2��Z�܇Q����Q�4i�r(he#�]�[r��6р��&�ք�Iv�Kӻ�Lz���=9�����5gZ&�-�,����4��:��g�����.gO�g��T4����k�)m���n�KHʍe���<A�mv*�܉׺�#k���y���6���8�_3wt�ֱ�]$�1c���E]d�0<j���Z��*05c��	�r�pÆq��3�l�%J�,������]��N[�y��i{�I]�{-�f��춦хZ����w���M��n70rw�-��I=��Ÿ�q���;�%)����6�{���-k.T�@\��ZR;�Z��(�Lz�L��Bʲ�z�/��2s��ȱ(�ʗ;�=ov��;�i��j��Iw��ra-u\����%N=x����%:g�����d�/:q��ڈ.û{���P�T&l���m����
��׳�2:>i�K��d*G�M�[��1U=}}�W}�lͮ�얖�*�s.W?��Ǳ_&�T��o�>p�w��fQd�Zc/MQD�oxˣ���
�+,m�٩��ɥ��6��ے�s"���1�sIn�KvN������%��F�݉srI9%�����y�]C��m�~����K�a�˔XoR�|��uZ�������m�2�CL,n��ͩ�N��k΢�'j������r�-���J�2�8��V0fEt9oH���z�w9��{r:�5i6��9N=��M�ͺqǘ��;�j���u{kK��ꐌ�aUw+j�ĸ8l�Ozѩ8�dZ;z�Ae�]���\;/>T���vs�	3w�H?�QB��{Ej��3hwH���`k�Rn���ڜ*Lʬٙ�qx��|^��1��+Y:�N�n�붓R��:��Z�]�tP<����.�����p'wop.S�B�/woX�x�]Ho������]X[�v'b]ǒ7:��S�+tU ���D�̚�n��7��3���CU���33&4��%���-wG�̤�\�m흑������k��&,�9�(p�y�j��y��fs�td���)�ksb�&�,J)��ۓ�]���V2`�2�]+F�]�ݛC\r�+n�zv���\�;=Ȳ�H�9�-�V�t���R�[�����܏�����d��J�c�O����8V�|�hw4���N�ph'�\�(����V�7o���RK�ـ�`ï7r����N�I����gm��HT��Ϩ������Z��9ذu�Q<)޻��D��c��';�S+�LY$uyYV���BAN���o�(�n"�J�LU�cU�����\��ۗ�2�c�y�'N}�6]���G,N��񙝷z�5���ɶ��2�C\����LG�_Kԙk��l������Q��	�U��^ud���]�7������_^�C�]=��	�Ʋ��c8ӳG�`������Y.���}��j��ỂjF��Dj�kS���w�����%��2���o�6%��nE��M
βZ劻�����،X�oue�kгP�$T3��1�H̳j��Z���R��f,�9�v�LÏ���5Ǖq��%v)�,Hr+�i����R׻��c�34n!ݺ�1�;�[�k����;�%��5g�k�4ӧ�j�̡G�%���;�:��X��FZ�b�swt������]�;0\�Ӳ+W6��6U]
����A������nmT��D���{��7}��-�7g�=��Xᝠ�+�5�	�iX@I��-�����o�ݽH��e��ɕ���iYe/{g9�#���1����}2W]5�=2���v����V�=f��f�@	����T)��W�*������]�S`�U�n;ۉ�:���V����[���۹�k��#�k�,Voq�i�ݢe�{)�M���"��}�����jzRܟM�.ۥ�֔{�	|�n��^��ի���V���z���W)�wE%H˥����q��g,�]�>5O�oV��WD�7���4{*5��c[ �$������o7C���FEV�KV��պ��κ9Nws�<���Ѿ��ij�(7���J�W7��5.��%��mo(�j��s��Ėd�Nճk������37h�]{��wM\���G:8�)*N�*=I(�\�n6�DZ�5�DӮ�u,Y��r���ɛOyvĵB�+��Gw6����׊�yNΔ';���7"��m�����V���l<��.ZJ�@Mot�i#�X�ہ9;�'<s&$�y�8�T�`"�{�و�K`��&k�l�V^�.���D[��Y�vԒ�z(3�2���y�o�dsS4��u;�gjj[��gfu9�uEEȯZ����ҍ����4:�^�P��ow���.c�K]�\���y_osګ9�!p�`c���]nѪ�������-=��b��$}&6�I�냲R���m.KbKZKZO1,���j�v��U�[����CQT.z\&l��t��oWD.����p�33�X���:��1��Z�,VH�����ړ�N֩	}����Ŵ�Rt���5o��q���-�(���.��U�+YgG¹�A���W�359��yr�ft���U�yo��

��]��ơb�u�����(#/kdV���~ �PC&sK:�C��켴�K�vp���ρ��� �;�h��7����4��v/2ŕ^P6���Gz��J�e�蘠�����2�F�� �4�Վ����f���{v��t�ǂ�R᫦svt��i��nÚ{-�7�q�m�����&=�i��I�晉�B�����EҬ��.�%�>������q-�-�ff�h��e�1���
�Qq�]%�h��k���̵ȡ�]�)�2�6v�N�r�wh�
�L'�Gg1rŏZ��P���^��]}��F���e��#��nWoZ�?m��Fwϑ�] �6^���_��B�V�.�/N��ެ��k�I�;��K{�Մ��t��t�H<���&dfvK�6�/�;��w:�����+�� ^qӤ[E0#]g.�t�O0X��-��U�xܒ�|l�:�:Q�B���-��upan�ڒ�̴�$�HaK��}++7Rvv�a����G�%�J���^��,��Y�Y9��v�$m��篊�3k�*��nmt��ݹ[�t/��xz��5�s3+n��V����e�M� u�0�a�����wXS�pn�GA��;��x��ڜ����%���x�<�P��}t���{ڐ���=y�9}q�j;۝��:S9��L`�һ��oʁ��d����r�sc�+���osYo�yG���qy���&�%�Z�K�ڜ���N\�������r���H�H�5�#�0M���1L�ݏ�����Eu�Y�[�-��2a=��dv�n���al��S9�����FfYe&t��\6eB�v�uv;�{�)N���J�f��<D����7x�Ρ43�\@�n�ˣWL����cs��2��Ż
�9��V#T��d2���؍#�\��тr�n,٥+�ʻ\���ǯwww]���-{���/w�r���K���(-�-�L,���4���f��#ږ���G/v��pr�a�����u��F�ڋ7tGf�n�F
7�f&9�i��t}7i�n�B ٚƳY��p[����BWR�YYB2z�2���]u_�^u֧��9�ybxꆪ��U�C�]��׏��}>2��v��"`ƛ�H�3�A3kF��m���+n��WI�q�+�9I����=Yy�#�ٔ��ŕ,�&\��2�W�A���0g&)���;b�9o.K���ׇ���41�z�0����ꕽ�i�*u$�R��b�Ĕ�uwx�D��Zf��;��2(�7$\�P�?�a�o+mf��;I�\���kN����+�S�%>[	�B���v�gFeͪ��rC���wٜ������X9l�w�v�^��ZT��+�-�p]ѧ9Ov�U�rMJ�}6�}�)��� ����P��!v-�͘�L�wj�T
�r�,�X��ܰRm/�1�V�vgWr�G�|��s=�5ۇ�u�ܜz��o��#�79�il�t��6���C�#��p�ԉ�Z9;�^h
�%�����׆<�Y��=�8)n�mP���՘�b�$;!�o0DM�-ܱ��D�N�����7di��U���|X���XN��>Os{�����.�V�l�	Zn���&�8�7LL؉�q�L¦2�u���z�۽p�� <���O���\j�m)sj��+D�n�*v�}s����7;���޻̚��)�3�uwGE�}�	OVҤ�;5/R�jlpTK�Ǜ{{�h���s���b� �z	��(g^���<5� Fʸ����J����S
�5dY�q���%�ҕW��,;�x,]�u;��6��i;����g-��0��R�2��/iX�:��囝��t�ԼB�rZY��:��c7�� @cu���\/5���7E;���UC݌���X6)�X�׵U��8F��0I�on��TQ�̒��r3���~W�Ĩ�yۨ�$\����s�@D���3�hӺ\�|�]��F����ؠ����Y�>�fa1>ͬ�1J��a���f�ow{%�p,��u��E�y�\9j��R���n�8�����c�4�V���]ju���G��P4��T-�ђq�-���T-|q:!��w���Z��gf�lx�0�\X��蔍�]u��
�H�e���o�U�r!��x��p'h)4 �[��˫m�P�y�0��&\Tܾ����󵜧'����#�9/��D�L m�t9�� ��@9l���-<{	��@��������v%�ͩ-ve�V����d{�w=��r5�P�ʘ��{mN����5ن�����61�6�Uܗ�ϒ��t37rh��%��e%���[��'�s�8Ϟ�m�Z;����!�צ4���&��u[s,���%�8�mQ��Ǒ�nN�K,µ��.����Ƀ���MU�'1��.��[� i�P�)4JTb�C]K�F�ŌR�ܨ�h�=e/1.�n��y�te�w��b* ��_�Pݎ�]9j}I�G^�,����k�DvR5n:�$̥r����u7.'������v�S�z6is����h�'���n�Rɓ��R��>�p���Ԁ��.+�'U,�ns$α7
��9�35�3P�V{����{����C�!1����쑭������nK�;�t�Z2�����X(��gbG:�;�h�9#���9ܷ�mr�'*�ej�&��W󙮮-�|s� =�)VX'�8b���j�8?�mL����+���<��L1^��%5��V�;����eb�/nfC�Y��2e�a]Ra*�5����D(�ު�2�譎�P�4���9�	���Lc>	V��m�m\�����m����N_�eWC�O[�ݚ���g0�a�+J�`f�ù�V��VJ�[�����T�W5p�g4}F���',�k�vX�����0TQ�ky�3�ev3�iYH4���++���u����d!��2kZIX&��J����ݥU�i���4�ǝpTë&��mO7��u��X�W�5c��ei�+��]ͽ���������1���S��(�@fհ��<��㫎��\��½��o�o�.{$ͼ�X��͡���o�-
�č�R��B��1�%���W�kY�^ewS��֢�^��n��]@���ȘE�5��-l#�:����'��{�m[zd(wl���f|��ξ��p�u�����W���xw���T�;�X�X��G�m;y�I��N�����;��ڗRSz����9\'=jӼ�c�k6��E��a�4��J9!�]"�nWg,1�N}AX+��d�U�S���޵�0&Fa�3�\ڔ�yΊY�S{����X���!ڴ���L�ռ�e���+j��y&eY|0]��._vSQ�3��E�m���y�P6�n�Ű<o&p���ݵX:���8�H�1�A/tz�!�_qDn��u�X�7��C�����ՙ�zs3� NZ�5�}H��Qq|{n�kf�S�30=G��yW�hr����;4i,y�mm�7���K
�0�;2��:EŝNd�/�]�ln��_^N�S	�˕I��;l��(!K��u�]�彊�wcX���6�H�$̵.=����m�AR�	�;0Y�M퓂q7��1���&���оHZXr�s��;�/�a��t���w�%�v:]�3l0	��2�{��v��n�B� �내\�&�H�J��Y�˹�E}X���h�2'�I��c��޷8�D��X��F�5�*nCr�0c�+��o�����D���5�� ��4��^(`ݣA+���T���R�ݔ'�J뙁��|I��ݓ��rݼ�V�u�iY�Ȭ��T铇�Y=�5�B�u䮴pp�w�mW>&���U3p|;��7�тsvz_9F�#��AOV��eu5��'N���Z�E�e�a��Zq��X!��K*��Q�&y�MI�6z�X v�uώ7�2�t4����uQ�LyL5��R����ެR��B�嚱Z����W��s8-��4SSWI��[!��^:��+�*��Ա�ݕ��6:����h��Ӝ��i��F��N�72��Ņk���__��z%���W]A�	�vV_:�Q�u��]��jkx�nb��&[ϺJ�溕*@u����K���s�+3�������Y��%Yn�����=)�(��gI9ic��c�N�}*��]k��nS�tZd`�r���wA���e뷣.���������vi�3�Jg�O3*v����ա�ΣH4*��2�>�����;�g��y%kC]E����*�{ϥoJ�T����a����tҏ�l�'!��]34N��:m��Kɋ��S���a�p1'H06�l��6F�3�vC�д�R�����n�7�1��6���2�n�KO]��ۍ��癢�s$Nd;��aT�����:����9O�K�4.©�V�WL����d�\��u�A��tYk�[F����P��g`�}���4;�s��#37�Xh<�k�4M��*��-��6Nm�)�ݫ��d�Y�ۣ ����nle��=	AԤ���z��X �˻x�}�곎 �Q�����'���\�Z�V��.$k�	�iv+�*5;w8�%�E'���ւ���Rc7��7�n�sn��p��x��d�$$]��TUU�����∢���U�������!�ġ�|i�Jg6�9t��_���v��6��Þȝ���㹆�nu%��9��j:k��X�#N�I�.���
vV�h!��XͶ���;t��^��RU�kR=}�G.��#�r�l���چ/�J�j����5^�������[��K���_
o)�;�z1Ӵlޢ()PYȱ�S�F�ܓ.W�-35\�s�t7����I ��(�On���ݜ�Vv�j��wKLj݆�:�uYX:v����7Ζw�im�:�W'E{�9uj��r�]����Xm���s�����$u��y�.��
��8�6B�=Gg�균){��TF붠�͸��΅��Z]�&�'1ʪfgoc��Y\�IcuUjM�f�w��1)v��f8���eZ�֞���.]�{��{�v;ծ�d���;�hv�����_�.�g�L��룈}�'�m��D����IW�]�J�`�Dn��v3OhH��𕙭�
��N�W���O�[죖����+��
b;�:9:y6� Ji22���薤;fQ|K�X�p�gU�%1��VƵn���j�u����V�b�0�cj-3j��ÄD�����R��p�3E^�=]u8;�Do���:�{�VL�2�";3Z��:9�{�.Kp�Eu@$n��[���A]��9��&4U��:����O�$	�9��<��Vty�6��L����v��x��ٜ��J�ut,��Rg,���+�v�އ+&���s�|�gu��V���}��}�}��J��@��"ˏ�)�5�D�.�Pq��+6Pzp��;5���V�+���>�]�����T�"�s����Z��k��v��DĶ�Og=�y�gL��*X�S26ER���Ŏh9�7��d�R��)��+��״��wm�Ղ]ɗ���:c(� ��䆔�Q�s�M�motX^'-�c:�?�q�_*�u.v�Q���-'�z�j���pv	�����R*�dE # ����{D�d 7�r���R Ǘg,�5}7����e0����Q���nѮn�ꒇJ��rg�Y���8����x�ξ!�>��kAAU��<6waD�P���s��Z1�Y����,�WP6�����;��]6�E���� �x���Wv���d��NR[9���	"�b���A`*�d@K��o�<��VG7�{gNV��,��)���皽��u7>���nS䱮���O�-��71\�@�i�\G3e'���:u�52Ӿޖ������}��?�0�q���-�k^��ޭ�7�����rb�䨧�D�uN���;ըԕh�P��x"�6{7e��f:0�<����)�u3��F['�}���{#9�}x$k��j^<�]��	���l1�{	2�(�5��y��o�����u\��/5��)
��ْ�w0�7/Q�wG���.�n�P쥪fl��O��M#�DSo�K��h}���#��'��;Ǔ���z�[9ۄ��Q�[�خ�d]���,,��nU�p�n���2D���Q���9>'&��-� ��u�ՙ�� " �b�A��`$ ��
E��o.;U����qYv�UJ�BE}����G��F�)��ǘI"� Ns�Ms��n����枌�-:?m[k��}��t���v��/wbq���l�/�7��K����\p�W`�r	Ӭ��I4������`��f�hnWV p�co��Jˍ���>�������`��]
ehǗ���[�r�0s���;_M��=V��YĞfٲk�#%x���Zϯk���_Y*Dm��
�ء�)���Gn�)��;�f��y��p<��oJ���Vv��ց�R
���1z1��rUd�<TN�T���j���ɳ!��@�$���uQ����@n����v
��4�
��{�n� ����Qb�E�$@bEE1AE����
,��7��y��޳�9��}����w��oj^	Ч7�ֵ�R��V�Si���:��f�ݛ� � ��G��Q��s����:�*��	��-�����v(�M��cb�A P�v1(Q�17�l�:3%^�︗��nN��$t��9,�͌S�˝���J�[��|�]z�Y�;�P�u/�M'.��stu�C�!o�F�+��=����ʭ�g�k�8wb �FAcV �# ����ѭ���|�~��[Z�Y�*�����vn� �j��䠽ܤ��Y���nT��a���1��q$r�{,�����4������ʞX�W=N�,m�C������v��F���8j]�F��vH$H��>�*�"��#Y�޵���cgs���5O_ e �X�9�/CptA���^U����Wu4��]��`ns*��>s�j�5t�آ[گn��U��ħ�Gƣ+kj���}�W�;f���E$��6�%V�~�x�+�S9���Bb�nvefbw��5�˓���WQĳ�A;o��c1T��N�-u�*�U�24tN������m"6M�R��_>�"����	y��4�,>�#V��-������&Wϝ��ٷ��z;��| ��n/z�f���h�����n
����N�%p��0N�P]Y�'�l�X=��}S�U���L5nZ�v�ܼ��rw��  sE���'i���Z����+�j������N�A���K���"���Mɘk��LXF�������`����d�m�����A�c"�PQa�Ddd�0aA�EW«Vq�-��y]��ѧ˃y�1���;��[xW4sYS�a<>gU`[7B�Y&�if���Rc/��b�B[����f޲�[R.F��BDE+�*�����f`�ak=u�V���x��N�#rWF��{ۋ���)Z��`���Wբm�Ç�:N��w��Ѝ�WAkj���W�5q���RU�κ4b��)Zu��Z� s��ʆ��+{��;��ٜQ�<�+�u�H�E�!�'�]���g���	Ӣ.��qH�|��^X���f
VsFړtˉNKM�6d����ɚ��n��^����n� >����ro������5�$��Nr	u@�Յ��M�bvЗ�F�,�� ���������7��ݼ;��UE���*����"�$P@�d`�" �0F�$@b� +��;�]���v����$���`�c�яv��Ʒ[�V�I��ܻ���Ju��k�0"顼=������룵�S�W|+�oK>����*�ѯ�| ��;6z��f9�㥝y����D�=���e����uݽ�u+����V"xh���!�g�7�MD��35�VM2`�ep���[�mE:�𖦡j�������4!��ᣩ�N��F�kn���cs@U�z�[":u�1�2٫��Wgh�",�y�BC�\�3�s����>ޤ�އ�9�!�WN��]\Cm����a�ۛ�a��4��A�jV��嬫�N�eRοW�WմvYH�QPP��)�q��(>雑��v:if�dd���X�v]L:���#("�EDQ"�"�`�"��Aab����]o�$9G�_n���}���٣޾r��p�-�Fx��
M��	���%A�=��s��np�v#)�W��T�
>�+�C��v�H$2��G�Dq�q���F�ƃ��np���[a�[KK��e;W�j7�B̛�nN�,e�*����^�����X����TA��b��QH���e%+����#��ŧt�F��;�i���[v���"n�Һ�	u>ASM6�Q��9�Ɍ\v���k��E֝C�7��3}�Q�=Z0h��%jW<��v�W��Ҿ��7�C��D�c�J���nS��$fu9�^>�]ƒ������e�.�S5���]�Y����[�j�?���)Of*H�^�vv��8��N7x}�;�m�5ןάQUD��g������P�Xv7����@��PdA�
���$P�a1AQb+�,AUU���f�"�,F1��2���Qb��n�S�z޺9���$�Y��b���������k�b�ԙd^r�L�֡se�(T��\r�d�z��U}�*~mz�W=��J;��@8��Ѯ��T//3mH�����x���d��ޫ�ۺx�.��i6{]k�I"�d�Ĉ����s�Hk|^�Ƴ��}�[��7��H��T�[��oF��u�w2��8��sA�U�t�=\7�雫g�;
�xRA��	�)Ј��8c��n]������mǃi�����u`�y����/:p������j��)J5���#��W����D}bZGͼ~׽��
ݎN��䷖��:N�\x�8�*eͮ%&��s���Z��T����ZΞ�f�HȌA �HU`$FH�d������r��r�3�&Ղ���?�>����t����ͭY6�Ī���������U�;5��|�.U���O.� .l�eKb'Bڬ�;{*�}G���q�PvJ�I�K{z�57��;r�	J���\ڕ�_G���Tz��p�Gt�A�{�2g;y�Ï5{��@�p![��{�M�W���O�����si袑���;���ޡ� }���9�S�C{S�pv��p͓+i�N�oZ�3'K�B��z!(��ŵ��B�ٵ����t����[��)Se�orl˟���O�k5��;�O���`)�]{��N�N�J�r�K2�z=����}��W�߫C��`��c����(O���>k!�� ���:7���v��p�ƀ�{S���1"��� ���( ��?zяpLھf�UV5�R�> �d�<ߘ@���[��{��a�5�������L=lؠ�2�=��<�V�6Ʋ���w���b#XӔ^�x >��~;��;�Dﭢ4�I�U	�m���`��>V����F�׷:8pǜz�D|&��+�oh��gk|�g|�[�h^�Z0`�!��*�((
�	�oԛ[����M�O�y���-���8����O�ޮC/��w���P�@��ٚ#�N��vOM��f�@�C�gWB�e����`�[+�A��������Щ[>G�d`��);��v�Sv���U���Pz�u@���&�J�E���ԯ6�XG��طi� QV�c����)k��쥻]�왖�B��q[ά�MnV&�Q��>T7�#/><���|tb�;���ܠ
g0�1r�w��%H�n(�ݽ��$v��d����m(#�)�g�0	��"D'ЊYڧ�,�X������iWn @`��Ȏ k&+���1��W�T캮��,��*� ���Gģ�n�UK�e6�DXkl���ݷ��x4��s�N_3�s���E�ZFw�cdf]�8+���
Փ:K�|�P�\n�,�:젺9�V빢���V����2[ĝR����.���|����C�"e��������6������)Q�W�_lpy�a�����͋!���'�?��w��I��YU��uF�����+wx;7-p��Q��L������e���J�o)3e`�R�i!�̪A�[�AK�/1��Z�ZJ�"R�@�cd��M�	��	 @���:������l*(\S�@	
��#5T4�쪈��V�����2�����)�/�Q]>Dڰ8+�B�ȓ�!����Gy���q���%?����₠
�*��!&���Z�E"(N*��;Iu��Ԓ�� y�5�s��ݬ��c����V��Q�Ҥ:�앻C8#�����y�w����"{v2��&S}�Ѓ�s̸j�}����]�>�����V냼�u<��G����nTcs�0�UX}���Č�j���y���[�YnŢ�d-�֗f��RcI��uy �/�5���rX�B^_t����_�]3r�m��(V���r!L���獧�y��a��^��@��n��:t��[�U;�K���̌8�q��nU�l�,2���Z��2�f�����V ˙on�s�W4uv6��1�� Ū��U�å	[{uѫ���Բ���D��vQ"�'�
�Tz(W;n�d�x��fε�Wa��w��%f��k�`5��w�2��B��NEL�_pⓉ���u`;H,/�+���B��j�9�`��ζi��T���/��M\C�1�0��m��6m�; ���S7+_wT}��2]@������\nk��RS˲u�c�j��][ش�G;Cj�wiOyT�Ξ�xn����ii��+X�d(�q�v���j�F�h���v�o�-2 �֥mq���Y���B\�nʳ��ʸ��e�]�����&v�����.�:��˻�Ím\ǣJ˱�x�×fGQb�mft�&Һi�8���^!B޻ܬݒn��b���.��	��+�7l���D�RK4�J����
yLJ��j��%mM�e�4%yd��%���.�l�Y�$���d���8,�z�-��]��1駭;�&5f�i�ތ�s�Gp�|�GU��z
���k����Ǿ�>�=��$�i�r������D�s=�7��f��i	7�s@�����7DW@�����l8a ���1��'���Oq�����긪�D@G�ˁ��������d�*(
Qj%�IE5H�
d��X��Xϻs7���"��F((��菢'=>�PwM9�NI�逛5c�-J
:1x��6���#7;W�_n�X���n��Rx1�iu�����nlz�����*c��\�F3p��}�}+���C�)�O����1�В���ޭ��&Ǻt�U)Vzr�G�޵&���"X���}P�Ǝp*ym�f`��;u�_3.�ֳzv�X@|���PH�I����=zM}̒��
�՚/Zz=e�*�g����s����#����L��%�`�{^uu���¼Z�����	�{�-7}/���ևz�Hk��c��F$'� |1���~?n�\��h�B����͉qW=����[�m��{V�.ڠ���^-�Ä��I�{\�Ĺ�@��:��JK0[§��j����R�ЦeX��'ޯGЏ?+`��^i�5c�1�g� �,=�4xE�xA �E`�d�� "��q�Y�r�ǯ��""�
�� �P�k��舌5�>��S��m��4Na��]PV9.w����7As@t�6�.1��@Kr�N��/*������.�v���_J�ք�E.C1{{Pܣ�yϾ�����;���q�
x��^˫|���o\pn��G&�Th�$�c�{E��7P�X���ҩ�]7/Tt."��taȱ��2ti`v�)a�S�
_����DG�3�0Q��e�[�MZv%�r���	���Qo,T:�гd�>��
��Y*��c��p^�Y��	cثc�iq^�5h�3'�S��O=��Q�X+�G��C��RU���.$��sU���9wi�>׮�뺹 6�HJ�>{D�c�a��Q�6�Z�賯s�E3l��W	$��Ha��}�]�+�g��6�����{t�`�W]��]����V��	Dc��8�1�C|��������Y֘4�!p?A&

	�TP
*�QdPd�Ĉ��`#
 �)TTAdR,�:��ovytk�E��f���]�w!2�{��¥R�������UH-U ��i*UF*��F��L�ň��b�**L{�V��+<�Uժ�� Y}X�m{�A�g2���=b�~�1�#e�0�/x����f Mn���37ǋ �Q��w�%����G:�+�e����%_�����ٌ`��sD6M�M�����}��~�F�MwY.I螊x크|��[������V��o8�+�C��tBKg�����ǯ�s0��69QJ�V!8���菾�_""��c�|�X���U}����č�����5u�TX!��Z����J�M�>�:ns`u���N�)�����U�T*(4(�q[�o�+K�WJ����X����u�m�Л@���9�S;���;
O��ƈ��7�Q��������[ǡ5�b��'�8��j���w�W=+5��!�H�C����wi��mM��=o�4g
6T��s�8@�j¢������;}t��Yۛc����,�CF��$��TN���/4��7ET�/��c�nۖx��ߴH*����k�I �^s����pND�EEUUR#0�Y
)"���~엯ԫm
{�����!ֽ��CM3��ď���_��8v
�G�$H5�1�{G�cv�@������7���=�L\�d`DAP�ґػ���FU��/7�D�/G�}E�e6L�@:6�`�Ns/A�ʏWwfB�o�	o�!^�Q��f��q]�;'�
�OOrisn'���d.��}:�ƈ=:nm��7�d����}$w����u���������Nz���nW����q�	a["P�;-Қj����nKˮ��UX�ƾk��ג�O�~�:Q�4(�r�'�&dà*��DG�x\��~�Z?�<�f���ӿ�Vl��;�d8��U,iq9�{�{�"�����vF�诙�U�\~�e�=:�+��n��ʾ��H�D`���"#H1UH#AED�*0�!�,X�>���}ɶ��%���)�)k������+���p�-����S1�b�S�WX�Ϋ���Fܸ�Z��}E��ٌ�r�,T]9��O99�=G�WF�ﴁ��}_G�}��T�3\n[ �\סi��E�Rȼ�Jc^ZH��y$�x�u�9_��HS��n��}�jr1,|VSO˨���B�����J��T��3.{?��
��S/p^�C��?ۖ�^LX���3/'v��:p��|��3v#\#�O�;Eϫ���ʁ���L�n'���(���OכY�����,�q���HOP؄d`�AA���qPs|�8����̭B[.B�f���\d5��µ��P��'��wp�r�T��}��O��3��j�k�.9s���m��c6/��gS�g�P�G�D}5;�1(����مʹA^�˸"�^v�s�f��o��+%����൭i������=q��e��w��5���!<9�ݳ�,n��bQ�;z��*DR"� �����LU��9�W}k�9�gܬ٨�U���U�b��$PP� (��^V��*��7�7jz���l^�֙��BN��+8�kD��ͣOs
�k�_V�g�Uֳ�5Ty��]wS"Gt9�T$��E+[�.ގc9
��nA�r�g��ΏxS�0�۰m�~߽đ��>�ǔ���n��D�7����ﾏ���E�qҨi�-��<���3�*����_e��F� �A�Z穞�ք�Q�C�e�T��5^T��Q�,�����=��!��v)�����~���ˬ�<�VW��`)3��&�<�@�5������ZA��t7z�ltqz
�d}o�2c*%��e���T_p�p��us����(l�H������hc�ͬ����菾�]��r��?eT��$Zo}T�dᰄ0]9�ّ=`�x��.�ђ�iWh,���H�C��圩C�|����c�].���I^y���=�,��I�	�b���F#AA�Ƞ1�$Fg��N߯>{�c����9��������0n�`Q�=pԈ�r���� �� �妺�4�ܼ�8&�r]�x#Jp�A���V�bA2�I�}�y�0��60e�(Fu�8Ww�&�k�)��à7���]�C�������8lt'���+���N~>w����ӈ�/t�ȣ�s0��m9gc�~����3�3>���%� E�״"�TL"�r��T����x�=dE�����7*m�ѓ>���� )Vz2%F�}N��[Ɯ�v�>Dc��1n���~��&~� ����V��������}T;7z��b��-�]F��\on����x�U�Ѫ��4�='�=�z�߷�5�	���Oe��Sɯt���kW"�c��}���%__J4���R��TL�9d�f�^#�֧&8�1���
]�s����QN���zGq�h�6q#f���;c+Wn����;d~D^?��~ 0DX� �T`��=��������%�W|��	Ί��F
 �,"�G?@�b��O��ۢ�m��G�z��emfa���fw"�ل��85]By���{M@���22 ��������� |���׵agG8^��R�`�����A������Ԇq���T���A�]����Õ�b���������Ws��s�EoN�<�)㦯=��pgI��=GnK�>��D}�F� �^�V\d�ro{���	��ü	�� �E>M-���ٌ�/��jDe{'�-�4!�ۅTy	���'���$F!֫���n��	��h|����0�45T2
B�!(�j
��I#TTB�T����EZ��-VM�����'B�:V�j��� �]���5+C���'Rt�]Z�,�/��Ǻ>�z�P2y� ��º;	>���h�d�}[~�/ί���c����}D}����S�3�&��Pg�Μ�\i���"��cc���O1�6`N�U���;o;�<eB�٨"-�Ǌr7:�e�T�j��ׯ3UF:��d���a�v����=���I���Pd0��E �يN���k�n�l���̜EV,b��I���M٨��/ɩjPC�
�-<[�ī�\�n��c�d텊�b/�Y<�Mկ�/�Ig��:�p�i��^߹���h澐���\�!'RE�E�����_>��9�Usg;����r����M}g���c':������u{s3�siN������bO����k}g����{Z��7c�t�ub���*��ܟ��<lȖ.�a�Q�+$+�+@��<�ifl��¶�J�>����P
G�<+�12�B�0`a��ҨĦԝ��
6@�w���z#��c��>����|�.��R�ȧ$�u�/:ꏆ����eM�#t�78̼�C|i�BN9�A�88�x&�+���a��ڿ�>^�O����Xk��B�}���>����ѓ�f���b6��	�]�r��~2�������Z�i<gdj`�������$�;���17r��^/m1�n��x�<+>��ۘ	;��B���,� �UU�0Y�XŌH,@	�|�����E�����K�o�26O�$ͩ#��S�םt+�����/���gd����΂W#���8]+�#T
#�2��b���z��������WŴw�}�·W*�3�|���cc�Ǳy�~�$�d�'_��Ѽ]KJW��f��i�u�\�8N�ʚ+��mp�1�G5wrg��!/����k��e_\|��;8ލoz��X�p�Y�ۇ���xd��z�vM���3����W1���]��R�ܙ�g��1���t}���W{��ٸ���F" ��*��7�~s�w�W��gǫ�N��],�����F�"6�!`�'�T&�;��x��CK���9HV��R������d�����t������r<Ǫ=�31E͐����7;�˷?t�L��gЋ�Bu��A|��_�U�b0y�,�3��` $�q�>@�\�f��c�PV,Y"�AdB(
�2]s���WoU�v�=���� �����߮�Y�������0��Zg<���C*������X�0�9�����/dpn'�3s�i�_�{n�����7��42�Go=Y�oF��w��|� �!�:u��>5�rv<�27s����C��LXY6`�R"ok�P�}��N�etz�����|���҆y?6=���Fp�$��׌̐�bw"nK�lq�Mf����E���*v_S�G!���x��*�����nu���ҭ�G���hД*�һ�WA1Kcop*@���ˮ�ꆍ����,l�r����Pb�ӆ�W?�J��*ܚ��;ɳ6���J�>{�Ø�5�#X�շ��qq�Ƙp*����++��	�R���^"s�c���6T+�79�Ѝ��0)I}�R �xpQm��a��:�U�y���n�
u'6��X����@Ď�0���14&4R��R_F��@�

��S�·d�&Up��r�Ah�轂�M�Ц�F�]�X����%�CX�F�˔z۵Ye�E2�7�CKL��Ǖ6|���V�^�>�C�p8%�ѽg ���?�(+@ l�N�oՅ7p�����u7���|&�dP*�RP���]�@�Ҫ��:�E�{u�e���jq��A�Tn���^���ywd~?\)�Xd�A�1�f,|�Y�1P@0 ��'�C@QH5eXɞn�S�6US��
|T�P�f"~?	}A_���f��v�|�gY���Bn����Z]˴�D^U�ft�s�oroY������dPoXD���L��%�r��X�4T a���nI�G��z���}��c���-'�ҧr�y�5Q��e�6���E���V�dĐ�*�:�N#�T�9-��mmX�m�+ޱ[��Z!�@��+Wl\�vȨ����t�i���F���:K�.B���]"ۜ�S-��l8i���n%'�/g���9�G���f�����4W��YLa��>K�D��,�H#R>���晝���S�2�%�6�>BH��x��27��sk�7��m˻25���2�5yr9�r��:ⱇ+����@^ͩ1������;����	��_�n�J�xcsen��<ea��������e��mX���E�QK08�8s�Q�k,,�爌������)aw�W�3�V���j��>�{�N�������΍j:���:(�;W-��݊����9�IӬ(z��2�bvVD��ҰƠ�}/�:Օb��J��o8zB��I��Y�Z)n�k{���sq�$�vN˝j�WW�Z��k�c�2չ�ժ=4I�vޙbY�QP�̒T�~����#K�|�|�ǚ��Ȟ�3��;�O��8 �[:e8Uob��&y%���x�G5�Ȱ���#>n���v�C�Ԕ����d�7V�;[����/��a�B�4V}/8=\�+�|�>�[�Y����lS75��ك�:��1m���p)R�s�3[#�7�"�k����PR��\u	ٶ�t��1]k� �mv�0��.����zB�t=�}Z�h�S����E��KۣIÞ���s�G��S�փx�)r��9(�bL���ͻk�����U�"X
WԊ��蒨�.��_�(:9f@\7s�i�����c�T�zz��IH`o^ֿ�I�)����Ux��e�'��#f��~'��[Pi�{W�t�k3mx�va�L�{]*�lǱ�����oY��5a=$�BN'
g#A��8~�D}�2.�������'����#���"�J���6�N��DZ3-��V`'�MY�Ӳ��#�P�ǎ��,�biܼ����b�Q�:Ea2�^�{�e �$�?:�����W�;�}�w�ӭ�
���(0UQ" �*�gs^糯8sѫ��c޽:�n�)z�3p�K8>���a���\�g�K2��U'I�橡������F�7xf{�R눱��>�"�cPZN�{K��ХO���#�ty�%{e�J]ݓ��N#Ը�5T;&�H?B���LΩ�kh"0e�̡�e'4��1U�!��t-�IAF$QAQQ���F"��EA*�X�yT(�$Q�*�� �Q�@�*��UADH��E�����UE�P"(�U
2D *��D��� "��
���$E�Q*�EAX�ﱜ�z��^q�5��]Pn�W9t�0�vv���l:F�����F�1N���.�ڊ���1Ma��jM��GA>9D�G��Bs�(s]�}�`����5�~}�䑮j�
m�dJ�Wm�t��*�tj�ʈЬ��R�I^��pjU}�fwj`�)�c���OjqFJ.��Xj}G�u�xH3��k�0)�ً��c�TK�7�������2d�no*C�s�L�l�p��Ⱦ�I�1�S�u����/g[ܼ>��^ ��G�RMT��S��g�!��b�EF(���*(�"�Y
1��,g9�r����k>�e`��e+;a*4_��6b�����N%�\e��d|�5�~��1|N�jb��{���Q錋dU���X�c��GzgѹI�LTi�F���>�\/Y�E�;.��2��F�S�z��&gv��%��g��M�r����Wș�����}*�>.'N;���p+�dM�9�����iUe:} �qg"� $|0A@PE���A���Y�j��,���`�|CpR��
�|� ��>�c��ݕ��wfM�x.�ge�ʞ[Y��憃�+�x�9ך0\�q�������+"�7�s���@'��X((k!�9��@I<zf���R��j'��8C�	�^��C�u1��O#3�}$�i>����%�_f�mם������׍sﾼ����(��X����(����X���X����b��qv;�i=�tf��������=�������z��C$�TX��+#	!�� ����:v��ˍU���?�1�J�U��S(�D�X�95̌��B��=K��$��=;�[�E�j�;lw:@ٵF"�s��6��,6!bl	�Q�썞wJ`�D��.��eR՜u���ߩq�O�DG�\yez��0q���cǹ������tj��(^��
�^�q�녕'َ�Jbf�Es��<Z�a^�-�V}�󈲌�r��8|�tsO���>���=}���}��6�f*��D��X�?`�=�ew�g}l���t�
*> �V������:�y�9�_�ݼS�S%��s����r�+vF�*ǜ}U��f����h˻���cL-Vy��N��@�4����{hM����b��|>`n����kl�J�Pñ��n�`I�q=�+4��g菾r�~4�w�`��T�P�fA�rZٕ�8jnb7n�>Y���6�Ⱓ�̜|���4��nX�Tǔ��N�G#��P���"vR
>����yY#X�����cWY�߲��1�b,TX�cȈ8k\�W�����;�y��szo��P}�8v����a�.OM����A�('G0�5��4�Q�a_{��Ӧ��Ă���O���~͡���=���}`�x/�䕨st�al�{+�$�ͣ՞�>�4��Dqд��=շf�	�7��]����t=�;(�~\���g1���1EF2+�+��!;���_{��)�g��эT&������/�h}���f�%�1�j��q}�̨]{�2�{��,���ﴊ�b�;Uq���c%R{�7��y���>�]]<�`G5�{8
���B��t��+]>�y�&�-Pk:LFG}�~��)���.���Y6Ten�Dƀ�D�@n��ʚ��}�����Jmq�>��w�
�8�@�/T�r��1̈́��8V�I�������?0;����SVf$E�=���/εw������u~�ۖ��/VDAQ��"��TDX�QV*��
,H,��$�A?U�����E	3�P�s/c 򖮢�M� }5���2�x��	Y��6/^2���]J$��dn�)Qb�%����pF�"e�6��`�i8�ܵBӖ#����Jҧ�'�Ք+l��g3������U�g#N�:�Ђ���-�;���or��l�+D35]jS�xś!0�oE�&'u���ɪ��X߹�n���$�d�og�?}}�.��{ّ�0(��{����X#PI�������	ZY�x܉����2���q��-5���&�ǧ��X$׮oz9�}q~�,�;gk("j�B��}T� �B1�b,Xŋ�����A�����uc�S}�mE��WF�ñ����y^o]bbaV�vt5G�m�Ϸ"x�J��;%vv��t`ky˗�vo:i���&N����?��M)���ø�곈$ǜ:��Eq#E�m\f�A��꧘5��N���G!�8mʉ�.��=��ׯy��f"�� �X��H� �ۯw�O�h �DE!�{��� �`VD=��9�=N�]|ELq�K��X^ߵ��xQ�Fc���tD�Y�S�cCqQ��)Aa��%�\�f/��]֤Ⱥ��~5G������Q՟��:���=�>C��aB���ǅ�SJ�;,��M�3{U��sH����t�=�����|�J�Cܼhf��<B�����ө1��d�ü<�0�G�sG��k5Ǧ!�7<fnaļ.�tƖ0�)�Z([�Hnm��#�_`��ɻ�	yu+�ʏ��f�8�G��9y��������#}2L�2�����>���a����SK&8Oǩn[�>�o�(��UU����w\��*��b[iLC;2�M�շ{�-���vr�9+��x7v�(�P���4�p�Q3g���ѫ��^ud�-��|��������n�^���2^�N^Э�:�U'��d���U�����x�*��>$��#" E	"
DT �cN=������*E�dQ@UB,$A��	7���?y�dgs�nl��Θ���WX�֋���ED�,��U7��	�7�Ǝ��NȮ�*$w�	�7����`h�!�ͬ�w-�V1&z�O��>���]�s}�&'�p؜~=����C8u�2�]�r�{��N�u��0`�\=Z���:�9Ӻ�Ft�BWJ�a���Hu��oY��a�� Ө�QH�*�����/g�5��w�"��V�ބ��?'�q��n��S�q���x��?P�y��eI]��V�`��]б�7g��FCm�����*��ﳠ��?U}�Q�%��>y�1��d��tw�V̷'���L��s�ds�L|��" a��$�	g�޽�o{Ĥι�{��X�=Р�ǆun�s�4w�.���]�\���XU�",|2t�l�7h�����ǘ��Gq���1�SN�ŮW]�,tB�H�S���]�6�+����}O�S|k>Pb��"�,1H�"*EE�DH,X��;U������	|��}��.���u�\gY�q]�}��Ap!��E��ja �F����)�ՈV"����w}�����~|e��e����\��
G0�X�T=�G�[u
]˓��[�\Q�}�d�ݬѺ�Nk7;>�l�e�,���y���kGd�
*t�W��P>���L�^�2����"�{<���^3��b�E�F'�>�3R�5#�q��G'�%��uZy_p�
e"��k�"Z�o�̅���H���et�p$��%r��+�~.%>��éB_���i�,X�|93����dwv�\��������wà��t�F&�S2c��8�j7����{Ճ��>/��i��,�0�ܾ��$Q� qY��^��`�Tb���YAQTH)$D"1TF,��E#a��}xǱuE�ԋ�6�V��/�0-�Y
�(	p07�4��v�m#�u�,����}aЁΰЙ/!s��[�ؖՂN߿V!���)��AA�  B� ?��#�!D~k&����Y)��G�Y�k���HG�y�n�I�i�?`m�I�D�K�v�����'����3�v>�,qWn�������>�Ц2}��E��Oz'��7�,d�WOI�T�5�C?96�����1��9��L7:D��������Q��Z��gHᦽ��F"$X�T��0H(d��o�]u�sƻ��B���19�>��.��1�����<��ު��t�n[p6rl�УmT�z@|O�� yxb9�4��3�8�����E�X�=F^>>�
��M���1C��ܦ�u����g��v0e�,V��+{.����;�K�<��v�F�!�����X��#����T�����1�Ggu�ƳHS�� ��	1x˧�c�:b��RH�(�E�H$�  �$X�"�@Y�\ߗ}���ǻ�9e��RԦ��1��r4챎�U�!��u���sV�b8[Fko�R�h��}f�[FCӞe@!�)n���g�)S�������6G�oe�<�Y�:�瘝ܽ�ez��Ό���՗.�B�|� �Ȅ1�5�j�n��sEM����>"5�>���ʍ��,u;��5'D��AӉ�GVr&%��ו7�:����"K���oL�A�xL��JtT��&�W�P�]%v��v�%J�W����nX�o�ޭ��|?!�}D H��C�����ޢ�$���)=�Z�hq*2ms٣!X��+�|A����&�M�Y��p�R��R�S��o�wЧ��8\��m-�)H�7P~R7��}�g�>�BViUu�`{ƥt�A\���3޵0�{8�	�;�'�ε��Bg&i���ո�e��lh��t�kP6�׮�W���P�7�	 ��**��F"�PF*�<�Sy5mE�ϣ��������c�H����ɥfx�*w��-�_|�^�w�mT1zUK�Ѣ���0 �����Amib�4�ܣJQ�V�KB�
|���]�qu��G�}$�8𘮵 nt}Y�p!Yo��6��ԥ��̷u��T���WX�3�B�����ѷ*��D%�*-i��%����Է���tJTDD�Śjb�jđ����(�3jv��45$�m�fq��f+���� hM�i�[;��q���L��X��t%¡*�!hÊx�d����=�ww�-6Ů/;����?|0��� �i1d�/^+��NJ�)�2� �AfhY�r�H�*ނv>�b,��Fqc��`K�N:p	gVF�i�i���
�
�z7wrԸwi�@�o'lq��N�	b�6�hH�տ�度�[��q�>�Y���T+8�X@R-���Us:��В�&pn� �BU�W��n�����5�ьv�H9L:Ć���9�"^uuJ���ҙL�cAAI��2�xM6��	�)��g��D�P"�R���m�I�O
٘�  ��;\�b��R�4�3uQf�q�Ʊz 	��?
U�tZB}bFG"��j�j��T!CCIwW-�)�s�+�.cY�چ�6��P(r���G��/�C�A"�Q�R$��n���j`�(��+Z��5Y^8�j̕��t�����	0���hYY���eP�&OI�P���wuk����~�$H��톷H?l��w��.�z)�Jy�mU���ڜ��N��)7B���R��S�n�ZM���:�Y�_X���N쐀��좫O@�=)���٢�Tn�27���'er�[�<��9�º�usn��;�7+m�ڳ4"w;�j�mtV����$BsqCFR	F�SV`�҂�*YӽddTu�&�)p��U�Ż����%IRJ����{�۩ �.�K��wGt�̤C8sv�P���V��әԳFB�f��7��/�u�۸��0VAHld�ֹk6���%s~v���e�6�2mc(vՌ�-��[�_��GOlSk�"�(a$�{T��eU췕�v1�60��3�|xi�N=���o���m&�JMG��h���:q�6嗳sEr%7�h��F�t,�px��Itq�K���U�wX��*�V���o'��/︴�b���N�Z.��oj�*ε�JW�\6��F���|�5��E�����2�N�d���[���u��U�v�-�mC�8��f�l��h"z}�c��vR��)+����׏$÷��� �=&V��;�ͮf�t�*%��sX��(�tʦ.��}u�s�o*��_e��YYt��]Mge��t��./��ӌ��c1M��Ԟ�1[ϖn慺5`���z6��<��a�Ᾱ����E��`ݝ���]6�:��`xx=9�4�\��Xݳ���ӽp�[=����vM�+s1�E>�ñf/�U�H��VM�"��9*��/,�{�:��`Cf�"j��D�L,��EG��퐵��N�@\��iu���;S*�kc�wس�^kMiη���u ��W�/�bb�bV�Ϸ��3}�Z�K��*ߙ�4l��S��׏k��}�H�H��̄��:�z��u�AkNu�=F��V�V9B�����x��;� ��띌KWh�	����Q���\@�/,�fL���?J%�ݳ|�wS�P=&��x0~�͔b�+%��U(��5�s�7L������]�Xc�K� r�%}�������=y=��Ә,"*`�mB���y���]��G%�\o�}~�e��Q�a	��%���ո߽�n�΋����",���A3}=e�ig��i
��X�����kdb�YBB*2IdU��E!()((0X�@�v�!2}�W�΢���I�ݢ]�͑�r��5��`�1>B�+7�%{�nN��s��z��/����aI'��LV�g>�s��sJ�7=O�\�.�[b�}[��j�F��"H��mZ��7��#�L�]�f\�Xcb����޾�VS��K	�»=-zE��xmK�!��m�?7r7���Q���1S
<ˑWy8���h?u�xU���"���>�h���eW8����O�7��5�E����/�D=�t�f0�<Z�]��R�����z��M/{��,�;�� ���
H�EB%k�x�"2H�W��ê�X9ҡa� DWz�+4��
����^Q7�?�V?�ݑ*�{i���˓��ؠLGwQ����:zUP{Ek(#R�9���>��2���
��>$�A3�u�+�<ܨ�LƎ)Sc"`H���
ȋҳ��h>�S:��=��GVG!&r4�;r��^��[�f�ڵ;�_�xZ�I�Z���g���Dc�����$�� X
@X��ԅT�{nwL��eK�#S�(�ْ#P��	�?��BRu���tqVP�[*VZ��w�h6F�#���@����o1>�⒇�7�*�{Z�=��6�N���<��E�,�e�I=�y�)�V+�q>jm��u��ʰ�F<<�eu��`㮜B��(v�I ��R<G=����q8W{�;�A��_����Yw�"���;�s��N�y�1'ǝ��'��$�+��(���u鹭7Z��*�
e�W3���Ye>3/Y����ވ��}>C�C�b�u�y����3�q�vD< �Ty�����o��Hp0�y5��.�cg5W��nxU���&�9�&���_/W�!&���|�����~��e��*�ު�/eU�H�5|;�B�f`���$�LG��ص�]��;�sp�5[?Pk@��Yp��8���iA�sWxq��E��1D`�P���`,���>��f�~0�u^���0A_���% P�DH"���Ӌ�E�GoD&������8D\:�u�k3C�z/i���9�$D2���1,]����WONϒ��Y���i���������}�M�𥣽�{�}�}]�7X��(�6�>��1?wi�I���$���(#:]閇Dw�nQÇ�]2��a�s�{`�`N�y;e�Q�R'r\���ev��v(��^���6ߨߣd��eD�E9������#8$&vE�yu���w;۴'��7Qb �y���oF�����QR EBV
1�F ����Q�/��n󸅋�K�N���u����m��<�P���@�1��z�������`���BWLˀ�Hl >۱���t8�:p�y��>��tF�舊do ٘�2�jE���~�"�<��/f��k�+��_\�m���	��E�
4���0�^|��pB,�G,�~ � ��D@`��T_U{[_qZǮ�u��b���q��� ċUb�y1�$�y�U{w���q���q��8�F��[���@ԋ N�޸rjY�O�>����G�PEƭ���U���ް��IS��4�dt����DL����\.���W�/�n��\�ɝ͔fN_X�LZʉ�����H�+i�>i�*�O���i�G�R7�լ��[�M�o	nJZ��Gg���S{��zo��N�mp�/�:	��ـ�Z�OS���*.L1{y�C:R*�M�34ְ=����cB.�ys�)�z��Ԟ����b2�m�\�-�5�w$<�d���c�y�n��Ϝlл_@���pqjԑG����%ۼp%����pj�\�ݪ�����6r��e�z�W��ȸ9����ꤼ��T>��_���~��'�J�Y�2H��=-F�9�0�ȋ���Φo��B�Aم>bX��O��D�]/V�YLN���Ic\#�"�0����˿�O����D))$F���.1U���Ҫ�b��DA!�q�>�_�}�e>j�{��x���� z�s�}L�4ǲ�hLo3��*{��r {��o_� ؏w�2���2�C���ʍP��Ѫ&D(�od>������*|}�!Pκۜ3^>0#hA��w�.ܤ��c�|���@^P��|:�9�d?Y����O�׹�w>x� Ǜ�><&�^
m�y�Y��J�݆�Ý��:)��g
s"��^�h�\�enI4c�ո֞��}��-9�;Vs�����M��"�a8���;���H�C�������}�C�O꯷æ��b]e#��ܻ.K���Tc�U���1�lU�3���;Y�#�H�Wj��s=B68����D����/�%~尴�	�/��W���ܣ�}|���
z^?L���a����ؾ�Twy�E{�p�����iy�
�}��l�c6e4nD����!�5���g�]�����Ⱦ�ul�H �EPX��� �dE����* �$����ɫ�{�{���#�0$c	(+H,�w���|�|����>s�g�0*f�-�+ ��Dv����jvy�g���o�db���}�)ӽj �5Bcm�za���9V>p"d�c�~�>���\�����>��Ő�1��[8��qD�!�x��Y��]_J�g����Q�^$�{��׋j�k���w�oӘ)��1#3Ҙ�4t��#�9�@;�n��-�95Tƒ�X���*`��P�A`��v��1��ETUF*�k��?mL'��~�Z�=��vh�폮e%��b\�&iN�k���t��*�+�q��8ӎ���!���ݽ�� � :�5�?h�ޕ���B���
���:��>8�&?x�'�<�}����;�}�yh��C�d�^A�#��������lq�7�ï�
��O��dmtפ�LA��
�����8e�o��
tv��}��x���ް�P�>�~FI�����k\弫��X�QDE"�1b�L{W\�����F�Y�^�gy���HK�a���ҹ�z��׷2a�G���὾z�x$�f���:��
`4_�g��$:F|O�\���.��3�f3�*:4�,�-}Y\��A���� -P��K���crb|��!N�1:@�4��Ψ�ء
7hջ�٭uڀ���4�y���%q��\!1/�8(���"\�����H�'6[J�{��t#�}Gvh�o�������~�<}�V�\J����_W�}�S���.=K5+�x��N���ʉ��;�炶�9�Q�L��ͨ��7+_��K��rŅ�F�B�[i���N8O��r�Y�Ə�1�^�^�^%X��Ȃ,�'�+/���~��5��)�)�1�D��>鏘�蘗�>���f��MM�qӫ�7�(o����R&������O9������14md����h��A�x^�k��A<���O�c��.�A2 ��k5~�^�PV0VD`��@PX,��3[��~����Y=f�[�^mq�d�5����̲Ќ<���:�}M�ӯ{��Q�l�a���r�M�b��� }Jrh�d]���#�*{l�j��3aX%�����C��~b,�9�ΎOPU0�����,۬��''R�)E鬡(dMZ~��FN�N3�mz��u4rc�bC�gb�h���.s���;Jx(G������(|�U*�I@H��)������wY��w��>��W����ܻ����k=D��h�&��Oj���Xcl+'m�sgy�CKH^F���?  3��}�8J�'�o��u�Iݮӷ�c���]:�m�مT�j�k���qU�p����\�p��dy�k�"�@�ܵ�fWv�Vm�ë43[q�+{z9�1ޛ��ȧ��/�Yy�bI�(K�?}��b���|�z���ʪ���3G��,Jf�]��D���w���y|�w�Z����4J�|&��T+�_҈4�q��ba��u��tB ���DAd�(AF$P�

$`$`�AG��+��y\s��v�CވED� ����|Y�}>��Ƶ�c�/B�K��s`�n�^�Y������(���F[�n5s1<���0�Yp�t��vu;u�]Kݵ�((l���Hr��R���7��	���Ϭ[�*}i<nF���%��V��M�u�P���>�~���>���|�6��5�g�^��!��EZm��ׁ��:/Ц�e���r�aG��??׹{��a�ج�@��6V� 3,��)Y�*S!sلM�q㺶�(yb�11�����.��g%Ԃg���K3���c�|s�i˩�G��yRh�-��i�	����>�Y��Q`a:�Eh�8A�.�=I;��[*v=r*�ė���3{E�$d��t��>(����l
���|:���\�^�9\P�j)n�i�n�IۢpB�p/C���l9)��.c��d�;�&�J�P?'�'LW{u�\����3��,$�~$4{�;�>��f�����jH���$F��"��! ��D�U�D"+��k��>������^�exm�1,�!��Tg 5�r}�&Ǽv��������>ahC�Ό���U!O��|�'��4u�l�� OЄ��]°ќ����ڬ��/�����m�}�dR^�\�!�`���Mj+l�=�Ǩ˗��c{3E��G@���?]3���0�)��3*h[�㜽}>�J��QTF��#(�J�!*��ϳW��덚��'�'����b�2��^h�;LT�k���l\.cҽ�Mz{��	|5�Ρ+դ�_dcʬlV����n��)��%�/�!�w����^~�|-Rl߬l �/��R,u�a��2s]���T9鷌-�O�`�?=�u�`B�J[�\5����s|	Ђ�}�s��	�CL����w4�T)\hɌ���y�����5�f�^��U-Ö�L�k��DHF��9�$X�h��-�q&5a�V(�\;+l�ӗ�&�}��pH
�P�f����w+�vL[�Qٚ�^�d8@�+��B!"�ی<��8JP�F����aI��Hm@6����r`�C,�0!c ��z��}����ۍcGq�v��r�5��+I���5����/Xu�I�
`��AF��m��C�������[]������S�>�uY�%}���zk@#/�kY$��i���ʂK������־f�L���#�b˲r�KuC>Y��4u�8u ���V�<
x
_�*�\�9	_Q(Gd3P��V��l�8m=>ВIRDZ���D��v�Ք
P| �I���6E�u�M8m�7�����pw.y��/�4�@��R���YV�@�ҭ*��,�:ޫMs���JH*�n�v�1�%��t�jR;�l@�i0�:W��(D������9e�ے�9�@/�J������Bo��?�UFgO�uE��E+l���C�O�A�� �_V�cK�p
N��׮�m�N&-�\1�̦�,�%�l���Χ˯��P�����AAv�v��ES�޾����:JS����KQ97a^fI�bʡ��%!$�����Y�`gfM}�_Z�́�J��':�q�j�\⫪4�}!f��J�	r�[�6����s7o{�d�}��5fZ�ۗg�1p����(����0���f�\OwX�r$�m��u��ѷ��W&���T�ZR�P�Stu�,h<��-�ȲK噋u�����#����tY�h����]G ��4u.��nT�]�^M�ڵ����M�l�r=x�V�Cy��bt���p2[[Ǌl!)8L�{x���XIE_Q�m�e�M�{*�UQ�Nw����-���H�wv��Hk��PQ6�eR�.�Ձs�����=��nndO�KG#�o��%�s���,��Of`�I��	�)�T#Ku���ېfܽ��+9� x9��۽�������*����G1	�M�So�hRA�ՄT�Ս��m+' P@�0��[�������z�Q��Q�wx �"�	�(�9R ��u{ŝ�AWa�(!9��J�vB�䣊��1�mzA�nҾL��{��8��.Mf���_D��˻����9��S�ۉ��I�5�T�F����1Ѩ�W�6�#�ht�x_H	d폝�D�öw�C���PD�/8�՛x�
��z��QV�)�6�vs��bF����i:����h�W��Y�(��bM�ǘ��:7ӻ���i���j��X������⣰S����eEW�gO�������Y�xf�nf���**��~��}������-�8`�\/���٫t��,�Sq��XA�ɇ#�����WT�:Tj�V/5���qy�ݓ�xx!�R����G^l<��~/� /V�
 2) �$��1# (z�SV�"�F
�@b
��0EX�H(��X�U�[��'�DO0��*2�M��
{��r	��l�c�2����.���%{��e��Hr2ax�p���7�T�z�Wen���Pճ��Ss菾�dM�2ܛ�<>D� [#�Y�vR�|*u�B���-κj������mӅ�8��'�W�����(����kf��1�K)߲�����|�<��E�A � (|�G�����LH�=l�O���o�;��(]8���v��+��/C��o�Ep�>�*t������}{��q.@�D�`Buu2�9�ًWY:�hc�=���#�����lǕ_�b�]f.����Y&��#���`y�i���{;�������x����a�~�e�ƻ�͹`�}��0�R1>�-'aG+9h��k�:B5���7�Yǂ�V�ncU�4E�V�$��:�U#�9V���=]&�3髣ӑ��ޣ��C!SLB�(l2E�]�X �c��Y
dE����q�w9�=��3WU1��)H�PET�őAd�?� V��-;�uR�H�ؠ5ł"��
՜ͼ����.�먹K�u�3<F��*��d]=< ���.�}믻���PC�T��<_��V6���}�p2��79�$��Ǽ�2.��LK��)�2g�Uu��vt�����[�ĵ�s]:bV�` ����;e�3�K��T	j���>�}�SK# ��V��ڕ�'�4�� 7l©N�i�g	��/�3h¾S��t'�����t�Ȉ�D�W�8�f�pe���1d�zT�r%u� �\,�k1��?Hȟv�'����o�����sM����x��k_Y�J;�-�aL���\a��h�^:Z8�9N�R%��������5��$^�:��
o��C�N�y�=}C>9��3�W������I$	�Euj���4,�mր��vo��Z��_@9��$iT'o��j���Ws:Ƈ��$HĀ��~� u�n�Z~�o�\K����"�"0QYV�(DE`H����du��}�f�������f��cG'j��ѼM�D��}���=���t�L���b8ش�!�`�<�d����B%�`
��}�n�)zy/�S��UI��l�U�M�)�FH��}t቗*�9��dɷ����~�/�Z>��&y�EUөb02g�56C��*,$>�s]���x5�u�qZ�{��i��ň�F2A�1��"Ad�=��"ὯO�(GN��f�V���y��4E�јK�v��gV�;�o �aY.E89�l�ϓ�+�m�C�\S������G�8C��.tZ9��h�}�R�����R���#OM��j�W .oo�`��ͧsZ�zl�2�������ͭ�ͺOmJ�]t	Bb�D˱9�0)�˺]�k��X����'X� ��d5�o��o�т�ȫ"1E (� �E!�����!~�k��pע�-�ԇ}����CEly���Wuп���t�S��i��]��ͬ��Z�9hoifkg�z�*IN��B^wr���X8��=�F=���&���<-�K����$�t~Eb-K,�'$=c����Ŕe{�C��lӏLEm��I�Dk�RŌOa@�v�`����=7#ͽRM��� �sT���+}�7��u�R!p�=�6���������f�����Pi� ��t��txk��r����w]�+a"�=�x������;�cW�{2-��KY�gѫ��@DJl����wD=+[��^�f.���nLW�ǕԽG��(!F�$���������]�s��B�iU���J�n�2;FLK2����q�w������iJ f;���@^�"�;��K�d+և��W��.���} �`�~����k�y"*��`#FF0�"�+=׵�On��<m�u��¹�$�� �@�5����t��]���wGm���	����Or�^J$�}�ց��{3By�ϒ�ym`�M��*�2K�jl��B�^�ޕ�f���4$!����Y��Q��j�U��x��G{����8=��	ωm�#bT�t�a]���j�����X�l���݉�������k{O���3��u
��47�Q�<�v�<��W�
��Ѥ���~��x!Z�Q����l�1m�\�ɲj4������k��&n�}��U͒J��"B"H�!$XQb�Y"�f��?{VM��ǄO�kN�L,�z5��K���k�LZ��x��8.#��s�@�i�D;�8
��.7x��t��Zy�E�!r�3Sﾈ��#$��5���� 0��jk�b�e�v�"j�c��"*e��W@P���DÁ�с��ʆz��9���0�^�҃;���4�UT�8�ٝ����¨�U(IT-
"�*�d
�T�BT�ie((�)Y���[߫���z�=5Y����++b#bEI����"��1TX�TQ`�A�Ȣ�D~�9�u�V!��i|�|�~����x�����7y�Vw_8 ��7��+���vT9=|[]Vܱ[/����B�	� �z�Iw��u�����kl�}ir��Y�+��qrs�
��5<F���Q��w��z�1옺]�br}�B'oej�_����C�"�Ʉy�CaM�fQ����$N>=,�;��g���v��j�튊�BBCU����X�;̽�w嘸��J��$ew���=�S�_���]�	5���@D��3��_��j�eo�˓���$DNw���"�u�8U�9�a˞��-T'?w�1xo,�_xTܥ3�:\�{��NJ�	�sg�<ed�Р�~�"#�#&eg�yFMF�>��6�L�f%7[�jʴc�*c��0����Qjs�ֽL��*-n�t�@�zu�#��)!���+�\���G����*8�dT_��cUQ�@b�(##0 �*��
Ad ADd�b�O}���5��xȣ��GuX�+������zp.�]lV�0q��z�✳�N��{��R�VLl�%��U4�r��糌ct_k���cC�Cl��~��������]�R�UrގT��i���0Thޓ�gEZK�&ҼZ�0ʚ��yr欓2������|ew�3���
�����L-c�G�&}-rL�����N	Z��d@w�;V�N�dX�ȳ|�o�Z0�j���*'K��T\�OݔL���ֆ'f���۪��o*~��$�����}���Ͻ	�A^0ʢ4��U.2��	�����*�S:���(�6��.���zMB���`��nHV��S;=H�-��|5�;ԍ��Os�߄�������q���I	���W=)�a9���$�M�"��.�ŋ�Y�;j�iDS]C�R�8�6���h��|t��F����n9��n���}zUQQU���PU��ۮs&ֽ�o�U�g���y�y��(�F2�D����}�wOv�V׸{��s��7z�\,tըk�Fײ�d�#�P�Y�šފ?zm�Aɪ^'ř��o��O����ù���=+}%����۪�}kvu��5�{�c�ْ`E��S��ג��z�UԞ�-gu�W7Q��U��LWJH�,H8V�pկ5�":�˒tVf6՛�:!N��������Z6�\�}�k^�M聏1�=ך��)1g5���O0.ݪ��XՔ ����#�A�WN��`s��P2H��nF�����0Q���B($a�B9��{����g�c�˭�ّ���إ�&&*D����r8Z���N��wo+�+K������~#H�������Wt�έ�~�W�.���l�,�_~|/ޕ���˝
��Z���n�.Lp���zQ�]���#���hEI]{�'WNp��<��� ����37�ٜ=�jEЈ�x��c��J�ddPb�E�(� ���Z�'��{��O~�����`�,c�F"�D�b�<;���g�T��ttH#և[���t٦ ��p+����Z�j,�����iO����k��lj�n��tn������4<��8U_E�"<E�_�>�l�7<(7�|��f����}�TO\�"�m啭�u���A��al��,p�R��)xP�<�+s�P:�)V���mg�,KZ�s�⻨;� C���aUh\��E!Apj���|�=��N�O���?t���ĭsNa)�'�V����]��a=��E
��g�D}�?G����}��a��k�O��	��&�{s������p�Ҷ%�=�s�>��܈�G�~�6n;�>�P9����UK��k.������.��n~�}�p�`�3���Cs/�q'ǜ��B��\I��(�%�x[^�X<���>�����@�}����W+f��֌
�FنB�^�K��'��[�6������c	 �E�`�H��+"��Ȣ��,(AAH����Ǳ_�Lp�%�����˶p?ZX\���Xd�]G*O5ƃ�+.��;��*x����x���!�[&��fgf>��!5Feq:d(��DD?o��!a��6J	jC|���S�_UL�V	�Y"%?���WH�%��ѷa��Ic+u�f��ꊁ'�$CFu�=W��q���]�ɔn)݆���02��R�����O��"�uꬸN��ɜS��)t��Gn�����u6�y\�ݰ�]ܨ��M�m(S���5�'���>����{wk�}��0d'��󈈏m)��&�ov;�Ʒ&���/83V��=%��B'o�u&hM�e{�;����Zi�=E�\�9�G�{����WD�Ik�G��P�7�}M�_"׶w��X���Uu���'���~ك|c�YO��כmF��ZS�vrV�}e�7*[�����;z7��ӭk8��*�"�cd��PD�'\�8�u�z�{F�xg���B $�`��(�$>Ƨ�}�`�7+�o���)��v'M9��Z7{s]v�pŠU5-�yu2M�?I���������|$���q���4Vo�<�Uk�!�ީ����G�B3w��ђ}�z}�%��;�<8|�����,��!<:��y�oP�����Y��,wW#�O�c���'A�{�Q��T}
v����'{����ǮAA� �Q/�2
�0�|�ѽ��Rް��I���8��وo"'X"Q�x���~�`�����(q�p����Q��kR?�|FХ]�t˿�?Z�p����K�p�f��2��kos����g��]�C�,�5�F�����5�$���c��`�����3p�]ܞ"R$W���mt��H|��mW/��p� u�ƫwj�3��߽دZ�}�L�@��.���"%�����!ג�m�R�� �Kw<��,5P���.,E��D�����)���v�oUڞ��s+F�n�@m��C�A���i(���6�o)i�k1vY�Y��Ὀ@`�QU*ŗ6��W/� R�/0ʰC����<�w������q��#j:�ƪ��3*��f�L�_]l�tM����M����{�+�pQ6��W{�1��)��v��UI-D�	��'w�H�t�(D|�8/��2���k*�)��໫WV#q*-�h*ot��k�z�n/�޷|֪�v����Rn�3R����e!"'Q3�#K�A%�I��(�n�Z�]o a���	��b61Q}>�8t(A"#��P}�V����!"��m��xYЙ"�ҲG��I$A��
.�X��%�&�\��>�WK�muj�>�k�
�)�_]n�U(:I� �5���]�ʽ_T����Ux�1���
�WV���[�t�D�7��Rv`J�i{gm����ǩ�U����ė��YCT��pz���4-꩟>a��Oq�D+I�ۻt���J��]k�h��9wvQ����ܨ����X	��G����G�p��B�VU�\���^ӎF���v[���#�J�=�X��̍����̻Yׇ:��[���%_=�}��ު��R�q�������L�F��ga�s���3yN�THj/�����,����d�W���5D�I�[��wt��ͻ��z;�l�����y՝y)�H�=����WuoJ꾡}����:'v�HN����Woj��{5&,�:���T���K�{����x(ΩĔN��&bu������*�vܞ�4[�6bʽݵ��5���-�Q}v)���>A�+������:v�S��H�e��-����Qo,�]˩g`��0SU�c]Y�Dܐ$x�iD��(�G"0��r�*5�L28�`�:��6�8��]u�pv+cٻ"P@N�Ed�����}��%�i��yR�9�0�m���T��H�M�w�s�Zʁ��.�Q䌧�;��'R��f�gj+�Qt:�D�Q��f����2nP�:d��ԡ�u����&��8��3%�ԬG`L��:(!Vi�]�'źʢH���!x-3A��Xv�;΂^]I��˔�̊S�خ�����ᵄ3��I6�7�`Ě���k���G:��#J^ټ�D����E!�\:Ê��Aӆ.NA����j�:J�[37l�F8)�!��eu�s,܅�I[:��n��xs[(U��i�K\�
����]�T�;ב�aV��C2�Io"ԨT�;W���f�!#O��a��@�&�I��N�o���7��E��k%Ú�7��|>lu4����x�k9��#����fSہ�Q���q�b���!��/Q�c��3	{����u궋X�9���vr3�����>����/�M�� V7���j�����ŎX��d��F"��X~�	�pw�G�pz�k��4�	R^-�W�[����GcN�9GF�Т/�gYen�Q��o[#�q��+��c�2�~���r��[��꟫��o��xnM9���,Õ@M�{UT�P�>��M8U�7uUSf�z39���{�>�_��jd�k4x��0M�kEinv�B������j�>�+W�>���!���gG���9���L{��}��z���Ǽc�������m�3���=��v��q���c�9Ш�N�{��zl�J��/:�OV�:P=�W��^��f>o�(��.$8-�A0�t���޽�����0��%�&�i�rA�bskf�$ 1�)��"&�ȗG��u�o�f�j�ۗ�zY~�@���ɭ�#P��:�:W�2zc2x��W�|U
�~�p�<k��ף.���#����p�9�Ȭ�gNu���]=ƑDTb�"�dR
"Ȩ��X�QD�B��c#޺�k��k���/�d�E@�>9����q~�Ʃ���o����z^_Q�B#(�Y�q٦�h�}}n������0�������*یvrLO\��>��%�R�C���Z��~��Y}R�~�`���[><��]�	��b��Ω٩��{8��٧Z� �:}�^�?tL����18��7�n�|��JdGM��8>�IM�޻�<�;�I��T�H1���� A � �H�OUF�c���?��3o�U?�A�
�6�`c3},5O2}靇�Õ��w�{�`,�a$$+�_~k�{��E�r���unNU��C.ʔ��}�iM��2{s˔�4��c�*b�� ����0��5͑��J�V*�Պ�D�y��q��=eϧ�-'����
D�"{�ޯZ����y]�|��D�ޚQ��'��7
}J	���yn��m2�k�MŚ���k'X�;�f!h�&T�dK������\�Ҟ����>��PE*2
��AdFIav]�*I�7��fu �B\s�G�5�	Qc�E��جw��ۭ��+���N7�xM�y��'�� ��w�bڃ�5��S��ۊ�t!_����d��7�vٚ�ғ7]������WԄ9�=Wgˢ�����A�~$���Gĩ��bլ�8����z���L��'��9�n-]��oUYEPz_bU��t<مsk#�/���X;�N��)����M�$)���:�o/;ڮ�@+��=1}�pf�Q1�dǬ+B�K�� �"���ݪ�P�̺�=*T�l�5�c&՛h-���F{�t��\ȏ�|>���Z^�<Q���\r�d�^��f�l|�MN!�w���2��n���4��X��zv�v��n�M�D�W�J��vE4nF�Q&���DH�ʠMp��x�Sg�P�*�q^��z���0d�aTU�$�����P��q95ze
U�S��Ы��b_e�/�9"Be���b�*�*#��D}���o�.�OQ��X��
���AB#��9�~�E�c(u7f��tGOeu�9����i{"=�����5`��Qs��O�d�����"bbj�!d�28̂�U����Lrg �.���ǰsæ6�:�� ��ZrB�{t4����vG�ՠP�����g��a�;�������,�a�>�O9N:��U˕�^7Y�}�����|�VE�D��H����_5U�oO�����������ĝ{�ϳ^e��;A��w�z7C�Õ~�e<��3L+�W�,f]���鋨�x�y��\�Lܢ�w|��1�� 7u���2��]�X�>���f����%~9�V.x��;y)��ܷAktAqW^�Rl�P�p�mRnM��m��d�]���)dj4j���4�H�ݿL̍F�a"}�%]l�j�ՈA!��
j�Ʋ��b��ĭgZx�]8˹��)��^��Hb��慿{��vU�y��R(�X��F0c/k�s�q�W��� �(�U��2D��1`� ��b��<��sM�k����y�A��H}�'ȱ9�Z5C�O�|��)���Pao��=�S�*\�[�W��d%���4�����V�n�uS���L'RX�����O6\��P8h�NjU2l�Y?*��=��9��F��+Z44���4����~�1�>�F�/���=�����@��9� ��f�/9u��Ư=���EF"O�����s��`_��P~�slo�SWI�/�qȐ��R��b��0q�	J���>�G�=O����e���u��s�133x��! LmJ��Bi��i���s^�����;�$z��yeϥ��g����v�U�r�鏣E$��{�˟sX޳e��՟ۚ���̮��\Y�m=�n�)5���'���!�n�lZ)h�Q�v�����m#���"���5Rc�s!�O��C������D/r8[|�k=���固*�{�`��,Ec$�d�X��Ƞ�(�H��L��V]���D:�Ѫ�DTE� �*�EDF1b���c�&�}kW���w��+��h�!�AÈ:�U�zJ�b�%M��7�/�K�Ț�4�1%O؟�����ԅ��-��.2�@}��U�v������|�����~Ӳ��;N39��E��}Ӆ�����=��1�+~�����K=x�;��@��r�������E����Ӽ��ׯE�[�9(�􁼰X6ۧ|�1�g��-R�u�[x�HҏD�sm�3�)��K�b*rnYp⸸&�фGE�
;Kĥ�[��sH���^�_�׷�3����|#7���@�ة".r97���@��F�hb�Xr8h}Iم$@�uޏ\ܵ_��[$!n$T����������zX��=.Ym׆O�'m�F�#��`�s)Nr�>ۊ�g��7��^p���<ޱ��,Vt(Y��S�7M��2a�Ѥ��ع!Yf��î2��D+��Gr
ꢪ0�w����` 2 ��~�q|��TأV1��*���E Fɝ����{{�r��E�l���3�.�N���(�#K�'��J����_s�����TuH�R���<���$Y0�U��_��:��`�f��G�#�,�G�"-�{d��틊Tl�#�v�f!��1"�48�=2�G��"W�]/{�SL�ެ���Er�ܙ����h��
���e^�f��� *E�0�,� �D}p��t�朘�	���ٕ���?J������&<���v�w�C��>��
�T"�}�JD#&њ��i�C�D|��:v"<��b��|>��Ul����S�V�Ⱥ�Ǝ�rDAzl�Nb�iF�Lj�
!�����P���%2et�[]=wN�;K�<�|�{��w>/WIx�ښ� �
�0E�� `�@$P�
	�Wk��z�j��k��<�5��۾g��kqzK��\i�#9��S��l�����|�o�f��X��V{]���]�l�a��ij��9߻�	=	�1"2M�T<p8���s�˭~��E�`��6Nu�5a��ԃ��E��քu{�g�d3	��y��b��0�^�����G*�y)ht�G��'yB�}�Ч�<37R )~̪C�p�X�y�Af��PJ��w��b*H�n<�8ץ��ꯇ���pV1�����',�DȎ������(���� vzTM	;C����~��$R�sr=Ģ��T6�w�}@��
SګѺ�55�>���u"i`�Y��@�o-�\C>~���*][į�Sq�J1-v��Ī>���F�W�T��F��e��6��C��s�7/�a�ˉ���ʩ�l9����:�(E"�>s��
9�����w�E"1P"I��������w��~�J�����S�n�O$I��H� ���s���yG������?g}β��H���.��eD=P�b]�a�Ӑ���цU���U���_��C�M>�D�SEJ�';�g��bVq�w���:p�3d������T�4V��eʫ��W/�8)�6��`L�<-�%~1sp��ĸx-� �_�������˄N�V��<�hv3"�e:�Y
TO�>�Ҩ�x�DWz�н`�닇�acU�Ro��N�V����D��,^���wKɜ�a��׫'�G��r�b�78lE�\���xx��Ob#�+8!��"qЅo�Pb��H"`|�B�kۜ��~D�����J�/w�3V[n���8��{C�>��m԰���l��@�e��Y�<�4�n�r�+1���U��d�g�}L�	N��y+�i�ϻ31n~�̬��2�<�1���3t��uqX�^��G�%U�;^���N��1��fﺱ�3&�'����vQ��v?{��M"Edd"+ Ed�y�����E"(�d��,�� ��ϴo۪{�w:|K��ݡ'�Vr����ɧ���{ۿ�� B>}���Ѽ���G�1��բb��Q:\�) ���u��)o)s�����R���T�!�wff��J��H���8���.oS(c�S����ˤ���e6E�$�P:!�ݺ���u%7/������gtT���g��P��>Ĉ�"���VP��%��G���2g�Q�c�#ڑ�ω���9�z��>s��}���݋���]�3�M�־�
�(�EA@�q�ٮ}�v���"�8v��u��"��B���B����2W�Xh�w����^�`6�fh�,*����uW
�ČY��3sl\����}�|�}g�j����9c߈��H(M�Rb��|.��N!s��[7�&����"羑��~������3U �����Y�x�a�����:ܥ��U���E�DT�U�_����xU�ι�l�q$�Cw�H�z��.UL�-��ǧ����"�Be��`[Nf��?�V��B�~�J.�$)���rK!H���M�B��a��o���+�3B���bKY�����3�����z����q1�^��
���;�������*�U��)�g�&k��t��̒Cś|�(Y�)RoM�u_Z��f��(^vM�Y��SX0����Qݓ�Uv|���-/n�J�-���J+<%X��V�aE:=�^�:#�дӍ2��[W��7ÇYC�d���b諩�x������S7DR?�*�h�N,�R��]:��������$�|�Վ��5��W28�mY�QS����S5W���pL#�ɷ(C��	͇U�l"k��s����$�I)H0#H,(q���51�Ǐ��u3.Y�HB���9��p�ZEm؋)oG�~��W=�-s1L�$?��3O�X���w��̛7��E��sΝ�o4q)e��*��n*���>���^3�
�A��D���ˆ(bG�_@[IJ�rw^s����N�A _St^f;����d�h0�"��aI� �%汬���*�k��TX�4)�	�_l2�����+
D$�O�I���-�t�Т� �Qk7XL�E�������0+"�G}�Nw]�ٍ��[�taA�!�1?���-��N�K��b[���(@KGiG./'N��P��u��5E�8��)퉻���c:�lZ�yϜ�J�w��E����x�P��etf�=y� �wnU��Nd����+��w�7[&���|��yO:����\�]}��J}����z��_|9o�\��#[��=��U���L=6�H���h�e]���s�$�Oq��Χ=�Q6o�ESx]8����ܶ�)s����J���*%�[[��۠;���m�K���k�z�;��b�2�M���fǖ�.��t�d�'��wK�z��m�]�(h3·���y�
X.T-���R�ЫVo�L_+�3c��WKyh�Av#8��t��;�V�"�n9��&�n����<����p�/:`WrJ�p��$��gv��V9SZc�Pm����m/쵅��x��:�	�5�r͔�
���#�+xeK��I�f�W��h�&U�tr��v��Q]1�c���Yx�iz�#K���7��+@��g�����[u��nu�z�Ǡӡ���i��uM��3��ë�"�\I]:��u�c�J�+��^�&�\�|�_]��"aS� �f�t��P���ľ|�^苫�2�9\H�ޚ%�<��{k4��W�(�Iw+��{�h�l�+%ӎ�Z�G��*3��&9a`�͊m=��gE=%J����J�6����ϧn�Ö�7�
��J�{�D1��Ev�Ŭ��7]����$��9�c��˳С"�;8�N��Ƿoz+&���ñ�|��*�L_p����c̙�0�J�T�G;l�k..I���b'�LE} o�'Q쫌��0���y�%��Oﾏ��gֈ�َ"�tP���j�s�9.��C�t��aN�n��4�̚\�@o�=��no�
n�~�r��(kkH���"3���/���&x_� �HQQE��""�ׂ��,���g�nu+��×�)#�^T�N�r�L���FM�1�]�R�;���,�
���;�|������A��{޺^갃��gfIR/f���x�aNd?G�}@��ϧ쟪�Hv�;Ԩ��$�d#�&�=�i<��;ɐw�N*���j��D<h�t{S�Q @ �J"" �0c�w��U���=�ޯwZ9Zû3y�v�>~��Ȣ�H@Y3 C�7�n�秫w�6���ݴ��G3']� �\;�ƿ@��?B��·�8��� w�����X��y�ڲ4m"���eM,!���j �+��i�|@*ﻳ���a$;��9�U?�࿕�rf��0������ʴ.ı�g< �S&>�;}:R�Wb�ar�!���w�;q�QĔ`���@��o�w�Q�nсSfsVC8��1SKMO���{�θ1��\�Jɋ1��`�$a���N/8]kw�Mo^���o7�@8��0��b
AB�߉%��>�6��˜��� �lF8htӗn������m�ډ���+����?F��Ƌ��7�z�����~��W�F���OI;fT�����j�hQ7+�mﻒs钟_xQ��X�#3*���k\�t5�饧�^�4����;�����^U2p����C��-bl���
?1H*"���&}y�o���iTV,� 
$Pc �E�w�����=�﷌y�[�p�z�4Q��]��F���sl-.�ҥ�΄�zUރ�0��S�Q+��s�3j�<O\aܡynL��ЇP����o��}�(���b���/�.8r�����^���)�I���Ho2�����wC�wjmc�O�Z�y)˩K���]50 ��8�NΑ�w��M���T����2�zi�L�џ��p7���<��_�.i�N)c������thGD�`��+�5Y+_M
����U���E��0!�})v-�;�jķ0F 08)���E�lP�:��F,�����}kjt?{a9�CZL�1��D�e�?8b$#��}UYz}'�@�~�߽1�u�R��˹�P�z qY�X���Z6��X����x�<������'"b�Jb%�(˲����k�/�T�%_��x���dc"$���)���=x��}�5�ow]�����DG��ǽ�~G�G��睰"clG�O��?y�k�ýI{o "��Q���s>`�j�g���u�O�ת'����J{X#P�̈�[c?��j{d�S�=�w�L��e
ՇB�D�Iڛy�x���C�4��W���|����Mx&�@>�X�
;��N���a�j�B�$�f�A�T�I��.�M����,�(�ߡ�֑*�h���;ʬ�*;Nuf�5��V_;ʺ̣rp4-׆/��oN�t�G���'q��ɳ�q9S�DY"�$�Xc:����U�����k�kC��V�.��j����`v���I[�*k��!�t%��T�/k��iT4���<$����o,g#7Z��s:��Ь�߷ۧb��}�NfN?�7��L�g�?��?Uo��\e΀n���O)��y��i�zaWg,-���T�V&r9��$��Xi���S���T��V�^vo*s����j �9E" �`F2�>�������o<-k���u��/A�,�,QU��� ��P@�����N�N�����3w�F� d���{V�q^ alD�{3Қ�݁Ù�H:��h�ܮ�.��������Gǚ�+���߹�C��P��q��qİ�&r{H0_.5U�3�q+���,GdI��[m�C�F@��_�w�"�)�c?�67]�ݠU�^�+�"�4���EF(2*��"�D���EQEb(ƪ�LQJFSPD�,��^>�M��q�普���ng���BfX�I}��Κ��$n�NN�]�����9=�1��,����&�˫2��Tݥ:�����m/_������@V�]��|_/Y�Y��@��H���$J��t,���(�Wg�u2���z�}&[��R"�����U�u���u��&2T!�4��g��4v� ��m����[�_���:M�Q�>�F�-=�C���Zq!���Ӌ��Kh�LMTiz�H�R�G-�Y��T#+m+�2�Izi��1������q� ��e$�d�*,:6=�L���R ��c+�������o��7�ٚx����3��G�z�f�j���oy{O��:�w�����túz��b����Ob���v }�����fVA^%lM�{D8�}�HsKO�35��3�2���&c��+�T��s��8�n�0��}��B��Q�&.0�*���G��}�/�ot�"F֡���M�ć��}g�}������U��@P"�$���8�5|\k��g|a�Տ�ڋT����v�SU�U����*���ź�H����)��z��ً.�w>��mӬ�:5�����Nȗ������嵲�ó��=Q�a����~����+*�Oz������; d��[�g��'���|���969���&�q�e�_�����g�& �[�)��lC0v�:?z5�h���|,�G=��VZ�ޛ��2
�EQI �
H�
s����8��{��Zې&�w����� ��f�ѣ��ś�ݻ��"YP!xN%[��X.�\��JVz�����^��J���8�x�glgTF�O>���r��0�Ps�:�1�Ä�]o�}�x�����^?�d\G�>�n-�U:��
��*�aE���˟zuR�~�ww;�����[GB�y��e�I�?W������|K���o0����FB"�����f��߈ퟵ���s{H�4�i�c���VT�Ƿ��{�-�{���T-xh��ۭ�9���Z�4��՜z��;1B��l���i�7�\�!�+����;@�bbv���8�;ݶ�.q�@
U�^�*M�ܞ�dD���M�+��}r�h�]E��/��)��sv�¦/�ĩ�^�>�>�_�uVq�Ϩ}��T�f櫆��ڋ�9|�OuY�?^�04��:�&	(��+�����fW����ה������7���CX�RMF,����{_{�㺧r�U�SPQ�+"�,�X�z�5�h���G�[���b�����ؽ���6)�>��2WWS��k�tk="ڨb6�.2:��]^�Y\��lc�}&0W��� G����s�xR%ٹS��rB���-�kE�깣IH��~ۗ��h<��o$E>=Z�T�N��ԙ�u �~�qV�_?P������"o�����Si��x�ךг�Zv1�w?;�]yY��Jρ)�n>�r�=w37a*S8�EC�t��&�
)$XC�8_�c}��w]fˋ��+L.<I�ݪI�%�`���1"�Ϩ��7�L��ʼ��:��WQ��1��M1n��|t��v�a)j���;�1~�K�N���f�#���}DL�=IW�k�rz�p���J�|�]�JU}��d�A��� Oq�����Q���>٣D�y�����yn2B�L�
	r�l�u'Q0�mW�b"",c�c>�9����U�(� �315IX~E��jK5�p�XNY�R.xix
�F0�`(a� ɱ�e�p��/�g��i*\1�Aʲ�x7F���Oj���C�ޜ��~�;o�]�,4��~� s����z3DQʫG�@V~vlL����7�?Gᆻ2�H�_99��d��W+��<�m����F����M��J�� �p\ŏ]5�<0H(���AI�U����~UEp'�V��/k��u5*�����1Y��1J�qgf���>��w��?�e�"�:�n�F�G
eU\��!Ld�`.Ou@Ǡ���P�B(k�{;S���c�_9��u�D6�,�,o+f��1h���%���T��M��c1�H�mL�
�ނk��W�>$���<;MmC�
7ԙ9���|%�4�׊_��ֵB3X��{�`.���c)k��ã	�$|h�=�ٛu��Z��vyJ�"�/c�䭖V	����T`,R)$Y���oܾ�u�^+�����`+!"�a"$$}���G�>n`�z��z`���G@�.�����9G�`��KcA�Ѧ4,�Z�{�<�����Β׊��4f��?T)׽�N&TԥPom$�e�dG�>�|a�3K.dД'�\{B=��i����dKږ�Qy����qS�!t��W5��3ćي��*͑���~�(l>eS|Cʯz��<��Av����>$E"Dg�IU�S��.�����ai�5�+6K?�9�����u��<7�|R�:������х�u��t���=O/H{s��Wӈ�nA�u�9�r�`F}�|o%FE������~ҟVܘ�&��,����9+U���$�E��  �S��W�H�+��Bq�E��ӭ���s��.���Πvb�9އ�Y֙mU�������3�Y
N}�S�՝��z���A���Y��?;���EW�p{g�߰V�2{�J�'����w��k��=ʏ�f++EVkTl�s�'s$�"�����k	���r�����"�EQ �(V �$�
"�L�n��b�d�6ER*��U�r��.V���=+`	.\���YxĤ@�#�s(G�ʃrK��)]�*k���F�;���ۇ-&	�`��+�z��������μ'�� {�FA"]�|�fT*���69�щ�-�%��wNZ����tV�Ip��G�M�n��+��L�9�=�zںt����-�<WY�"�nQ]K!

�\�ęyI]p|J�_x��;O7��c�q ��6K�Ǻ�[�K�V��BsYb�YtDG��j
`����<ž�`�p��Z2�vq�x�n�L�%����`k10����MY�UhQ���h��P��HVA��Ԙت��7�0���ߜe=�|�ۈ���Z��D[Y�toz�׹��P�][�2`���n��:�J(%�5���p��jR��ag�|�e0�+�5.]8"D�(^�X��![��i�j��U�VP��ݵ��+��z�ߐ�8+L��2��r��SY��e#5n\�����xb��O�<��}vF��@K�@hh���no���W;n�x1�f�ZF%�$��W)�?>i��x�	���1��h�>]Z�[��I�}��Mj��4�c�1Ҫ�U;:e��kMhҊ=��G�� Ź�Ds�zmY���w��������6M�xo���t3�W�$J�?2a�Zm ��J@-��r
��{Ln�SnY�xԊ,��X��o/��1Ů�S��W�4� F���}��0c�H)UT¤b�R��p��Ѿ�����4rWYih�W-�v�JJ�T˂eET3t5��&,�|*�zf�ܠ�e P%��D�`n����*uU8AC'��ҁ� P̬�B�J�T|��nT��T�۷p��.nZ�]�VM0nc��n�;��-��^Ly���l�stt�Ǒ�54�,-%��k��n�2��U���D�G{@��-�޼���h�z�+E^� �9P�v
�pY��q��;Ǯ�6�.d�@��u�v�ζm�2�Α�%��4�I�y;:U�m66�A����v��1��j��m�|��wv I��ܪ�+��Cb�f�:fs����Wr*\�m�R�N�����sU�=��VY�*�{�ցdc����s�<��J����M��]c�ɛzB���<ʇ�7}��3I٬��~y���w�2qL�Ʃ�df�+q���+�m�^��ڲ�|yD�iq��ż�����k��J������0�vȺ�f�uv�l�=\h �i�ǹ�8�}݁U�t:�GWTת7e�i|������8Ӽ��8�� ��wmB�v��R�x)�	��	Ԇ7�X�^u�����Y\]�����W���g)��Z�U5����칂SV��l�yR}�=�+�sh�suԦ�ˁ��'��4������gJn�-_nα��*yϕܰUl87E�-8Ɉ�T7K�~�"'�c�#Z���9C�1�T]A�,�#Zz3I4(���/&��U7���˩�]�j�ѿJ��5`��45�W\����FJ4���3�;nѼ��T�|i*ˮk#�2�F��K�Y�{�����л���a]\�y�:3�iE����Ž%i��+�E�cwa;0�y��8�0�ؠY\�
qZo�Oe��Խ������'z��ԉUæ�k6�`�<��w74=������y���H(*�{�TW�d���ѓ������Ĉ
*,X
@Y
�}��Ȁ�X"�1H��&g��ڷ�ULh��lq���s���$[6�'�X�����kt�{���+�z�6Ê�[���J�n��;��,qrC19��g��s8�u�2�$/�}譱!��.B��s��I@�ǉ'���I�P������zu�KT��E��fhkdw'Ї>Wʉ���׹�0w}�:��{�oG�mH�`$��	I ���ۤ��y���p��>Hyc�ݻs&�W%!gI����{͟��ݪʩ�jΉw�z~�Si~�<��@�>�E޴A�Վ��f�z�T�G�� }��"{k.�iiϣ����������lC� �}�p��U>�!��+�����=^������`���
�k���s3�� �AEUb�R�"�`O���c5���dy�[��˔ep.I��;�ݦd�dpBֲ���3���p�<4�D���T\6���\��F	mouwqU������5u�|H�����d	�'�i|��F}�r?U]jy8!9i�r� _|9T��F�5���Oz�#�	��x/
�ȗGw��0\��Pd�\�٢�xܫ*��|�_��Y�Ǧ6v�C��p�F^�q��o/��t�b1/���������B��H�w�|t���� o�:-�<�����e��r�өym5>��%�i�r���B�������}�z].����y�����+��w\jUE�H��h�S��S�C�s�K���2y���V��.���K�mƛ�3�K^��1�3�9�D��r��6��u�d�v7�����idO����k$��Lt�_���y�WJ^0��Y���pKs9.p_R�9HI�D������>j�/�o4-
6w��1�F()QYX�b�*�"�"10DP��FA�A"�F

H1`�,F �o��U���5ݶ�ۼ����qn��q�Y�fGn����f<���rZ&�#w�s%^k�ޔ����$9tB��S��NA�Փ����7�.���7@0�:
.d�E�k5ڬ5�~����P�'�1��#�`����O5�-Xh�t��۵qVj�P��}:�4�y���YuN�F�[�=���+�8�hn��ZP����ƶ���Ư|=%���z4�F���I�m�j��w���[/�ϱ�c[��k*6��|�(�A���PTF���dh�I"�Ǧ~�C�@�n{Xp�^�������wP(R4v��r:�̴z8Ǣqo��Ȑ)W}�?X�!�vk���wC���}Gd;�3e� �/�DC/�g*8�/m��)Z}����Rq�u5�Or'��3۬�S�J���ss�u�Tro$79�_�6B'=�)��*�o��^0���WM}%�<1"�""E
� EE$"
1AUȋ$���$Y"B(D`,�Fy//��{f�}���veG4�$i����By:����kB�陸~�>5�ZScp'�-^*�&�w�Lͻ���{����K�����P޻���jU��΀�=ϯ����k˛l��(�]/O=G���9�Q��[|�LR}�0GH�zRx�cf�S\���9Ҹm���`Qݏ��}��5���zE�e�R<Ù�I �u!��CG{d'�ǭ֔��B�m(�T���A�?	(l���|�}�5]��ؙ�����r�Ʊ�������$����$��>�A�P�^QC�r^h��t��E{D�s������F��z�"<��=����812���5�૴��V��~��9��� �=ދ��e~}V�l(���n����c�p3���U�+�͈���:��5�å*�]�[4�=����A�_��F���uk1m�l'tn�aE�����T`�Q�X1"�(P�������ǰ<�V��w]Wy�$�$���f߂��U7���~�K5c���1�.��D��&'�E�ț^��cX����9�՞{q) �v_;��7���!���Mђ�jh�5pmt�+^�}�U��ls���;Kg<��|[c.P��K�+y�k/s%�C����rk�x��-�_�"&�Wj�f����r���`�'�I����KC ��s���?X޻'.S����z�v�["v�~	~@��m�Q����\��UBM�<n\��x�ѓcr�UЕKOH��	~��������؞߾��HQHe�)��1م���MR���v�TT۬�������{ń�!]�%k?\M�A��;5t}����u_h��hBv�iMP�ܯD}^,����dz�L��M!ە|(�LX�;��=Q�+ʇ��,�[�p�4u��;�!�Jt&:��-������\�Jre��i<�P��U:N��w����A���+I۾�{���q�!�b���"��H� �1c�w=�i�pqλ(kfQ8-����U}d)�R��a���jsl�U �ip�4��g��fG��;�'��n��>k�S�0�*��PXV l|sν��_m���gYݝԵ��ٝf.�b�;�d'|� �t���\+�[�v��m�]�gQ�d-��pvG�g5��]S� �d��^�A�͊�կE�β�nk�*3� ��[�z.�9�泆�%�Zl��D\����o��b=~=;0��3���p�k1S37c�K��v�5���I�͙��X0�U���BF! +^�~�G�5�_t��i�[�D�eA�c�7yQ%���_&M!t�%f����'SHf�\��nP���2��Պ{L*ݻ��gfP��@���a��2}�6�'E{����+x0��-�-sLx�&ϴ���fT&�0"n|��@�ۜ�z�F�G 3p��sEM�-��1�؜�g�\)hE��F(1Y,Q��d#V��"1Q��X�
��Q
��AcE���ֱ��T�}���N"������`�A�3�S]'��Y%�K��'�y�!ׄ�2�ځ�>�S�N+&3��Ն�J��Q�n8��&g	�}��\�3�;�*1��ĈGs��f�� Iy�n���Nq^͹1�j�vn�F���̧���Ij�ߧS�UR2��d7��o��Cn���P����\Ma�at6����h=��t�v���K옞f����w;��#�#u��Z��]����U/��ȣ%kE{�w4y�}�zw�O*���*ІPX'��߅A��[	�C�|�x����:7�p{w!�v��Ax� >7V��8��2�`x����Kt&N�� ��3<#��U��Wpo}���D:��%�������}���d������b�V��-�NT�ad��N�vG�PU�u�Q�ϧ��Е������p�b(�H,���@P����w�m�u��߱ݗ����/3߾�~ ���&�|hx!�4~�?A�r���Z�L�*˸[k$(�c:@*j�{�I^�}>0��+���~��n�J+�-<&��^2Ty@�O>�m�?iYY>��/E��c�r&w�V{g��N�f�s��v��J��E�t[�����N��W�'�Eay1��&Y~�J��i��p�\�ӷ:n��v��}v`�����uF4Z���7�\,J���2f�=Α䪛���������Y�����͉M�zJ�&E�
����K �qb�D�_}��P��3~߱�O��`�;�}��㕯�_3�뎚�W(;���cW�gL�s�%�s�N64��6v%��KX|C���x>�=x�xܼ����mn��v:�v=�D���byό��_��n�D��{`�zk�ʹ�yN�7��Kj�,��j�u�a(D��L9i�2�G��T
�Z<�T(5��1|iN�&��'ҖJdH��T*U4 ��!HF�, ��k���:��ױ�kW�E�P#V@P�����lx�ٽ�:$��8h#LvWW}��נЧ)�m�W�+ﻼ/y��h��v�`vPZ�xUx��O>���
lb�{��+���[9:GP�%����3+�6fc^��]2&k��J�;j���b��R�K����[����BA��zXW�ɖ�E)�������1��N��oz�����4����}�о�C[xB0;h��Cw�%Pq�ge�v屃gϵ���hn��t�A�;�'7vԘ�g��[Uw��'~����E��*�q��P����ND7Fә"9�;Y��><�����2=��{��V�ސޘ�cl	T/���U��s��O5ENs�n�\u�@������W���_�Gj=����{P�mONYqj�˙�b&�鶐9	Ztw���{ʨ�ߐ����s]s�}o�)c�e�;�I�����7���4�Ǯ��b �Ȩ���"�E� �
�E bF #�R
b0DF"��H�,V#ͅ�m7f�w��/vT��"�B��Ӹ��ځ=U�XQ��$��<���Q|=g3]]� �眑{�^�� ��_#s�D+����t���3�ڣ��^����ɡ��9yqFYx��֊�Š���D.��q=b��A�
�LJ�N��u��4#�7����\=�KLTm�3�K��<�����3�Y弼�?�E���r��3GՇ�}~�M
�F.�ih�Ȉ�
(�"���TaTQ���{���w��n���﹩B�`跉�Υ�7uo���-'�}R(�8u���8r#ݚ���˛|j�إ*��ER�����M����vg���ػڋk\��z��Y�J��]>���D�`9��#zK�%��2�1ۦ�39��t7�p��_N���}ދ���~�����h���։�<
6/�Zn�[�,z6��������s׽ZFĶ%aS�R�$K���9�ty�ȱ`��E@VF 1�)AX��"@D��$����g��&��W���)�V﷗��"�`
5 ����gΫ�f3��P��+�ToI�ށ��Д���vrp*��
(��lCu.���A뗣�[Oe��]�D�Ѣ}�Z&�����{Bd누�)�|���SH�;>���t�:����K�����'��
�]� �j`}���3}x숹|ٮ�����<}��"�Z�u�^�!�c�#���J�;1c��0��C9舟�+#��@׹����xB�sU}��uu�M,�]k��Fc����[/5��6CKqV╵ݕ#��ooe]�
���7���˦̉��N*K�{M��I!Cy�)}��b�9��k�ذ{5ܶ�d�ϐN��CUKm* 8���-Kn�<ϟu�O)y�"�f�'ۥ��P۔��|��G�"����4o���n9�p������X]�
Zo�7M�ס�l�f�VT�84yYn���D<�&��G%:M:�Z��^�*�3@aH)i�i�o7-UPH��/z����?��F�>�f��2�].���k����c�u�J��5SC�,�*q�q(T$�5R���]@�Ѕ0 �1��2]"��r�*�k\��E��2g���-,������������A�E:�����
\,@�vގ[g�F���P�|���X�D��������W-�b���ګ�^w~�%�H2.��m����3�f�v���Y&������A������
Ƙ��Ϝ�#$�g:=�]���B�@��V��w��(q����ŝ�mK?S�Z|��ʄ ~�$��F��DnٵM= �a�|�	i�4ej�)�W��d�n<&�&���`��(6�!��?2(�%G,m*�7���2���.�Ջ�T�5�%�b���(@D������q��B�����]�d�1vȇJ�xe5.��+����fξ����u�t�s��ot�ׅm��1�b4�f�������Y'���\r��Q���F)�p#ٛ�Vo�F>��,�3.�`��)KD�e}7��Sr�N�cF�w9A;4�ZΘ�����u���Z����້q���u�x7�"Bv��J�.�N�m
���X�{�*�A0��do	�h\��2>�Y3+���3&�a�sIWd���'wrH��}�*��u�hl�#��r�op�@-�l�S��]���)��S%�J�7��5F����X�+T�<� ⮏���ݶ��c{p^9���`v83+ �o�)Q�����KwI����.��]�wS��۫�sw5ɩI�v����f�\/��.ٜ9u8�T5��M<���u{�
Ҩ�*���~P>�VrX)�d�R�\ռ�S#O3rn��=�ڸ�ێ-�o>bC��PD5zY�J���k/��uwЇ�K�ޕ�)f��0�N���*֍��'UXжVE�#Y�?��������f���N�Չ&�dt}�x�:C���.�tKA[DɌ
����	�ܵ`�
��]�ɏlz5���kWKrb���u���V��c���;\�`�a}hf=�]p����Ǭi��^p�8��8��۵g��R�A�:R�7��{�{�2�u͞o��97�W8��a���*ɂ�/�i�N� �:H/b�Y��_Gr���G�u���!�2�`G�Cݵ�_M�X�;74ዛo�UF���9�6��n�c�#'T@���2u'[��̖�މ�Nbm3���R�r��s��$��4p[=�4.�6�Zx�R�[Hw���c�F([�A�\���$�����F8Vu�]�u6��F�c$c��5r�_��r�{>5Ց1LP�˅|�ԝW8A8��B�D�A�0�[�0Ȏ�v�0�o�a�-���b�fq�s^}<z���R��1�ţﰀH�,�k@����3�uG4ZTQ���(VDQB��W�D ��j0d�"|F��9
����l,Q�~��g�z�1S��X����3���A��ئh�;6��\-��/��nSa��t�Y���Q��K����a~cj��t�P��Ӷ�����D�l�s_���M?H�+fW?S*h๑���;Rt$����k֚�ou�n�MV�Y u`����ßG��Kn5���GƱmҟ���es��2���n������z�<G��^W���y���yN����Շ(h��
�/�Z:�b]\�;�i2���yY5��Yj�J��sX���i��%!�\:ue��ה����-r�>�܅�r�n��%!����^�;]��;�ƕ���}��~�$.���^ ���p�=��o�z��`,��N�����&�!�gsj']1�]21�c��a��0�S���ٔ3k/|�_t�*��DE���`,�k^(�u�����&0T0c$ ���of�k�e,_P���!
�$��9$��n�p�Q�=�pi�=���� �5��,[���ezo���r�_ekgx�JO,�_2_T�3C��P��|G���d<�՚�L��]�=��v�K.Ϩ���4KL�qe�ܒ���A	� �V5�i�"R��:0gi]m�";�Ts�sn`|�Ȱ�{a'3�V;��7@�w?JC�d��6A�:4��S%�@�.!-�ۼ<�$���t��}���m�\Dˠ�ފ�|�j�S��=����q
� `�{��{�G�vW	��vp�A��c{M�Ǹ6�P���'Xf��;�Dl�(��n6/l�v�/��:
�#��{Pw2���;�69��A����G�n��3~�ϥ��r��:4.݈�{Kk�������;�&�V�5.������?O���Y� �A ��
H��H���)${�ǌ����޻�����˻9��H�Da# A
C����~Ʈ�W�n\�2�`	�99��qb;��o�O�(���T��G�pw�Ж����R5���A	eU�t���}r��;��d��d�Ȭ���~wK�*)@5�;D5�.�.�b���[��՜7d�yZ"�/�F�2+:�~�;�����/��ߦ�Ԑ��J�ED�!�{;�y�2�.}�Wፎ4%p��ɞ�Ǿ���gnֱ��\���g� یT0���7�Ϻ,�J�3���'g�5C�B����F����/w�� ����VWI9*�xl\��]�c��������#��ՙ[S/%M���NͼJ#�s!�'{Gje9�e�6B�I���(�x�Հ��mb�NH���`�/��UєVs�I�6��(nzr]oK������*�A���y�f���!������� �V�QX�,@TU>���{��ky�U��2Sf�%������<;V�U����P�^������!<�щ[��h{�9���ɆI거�<�����J~d�A^���?#����59(d�M!Y�uw52�y�G-��}�qIھ[S�[P�u�s�T\���G�U#���W^�� �)�ܞ��s���s�:�����P���߶ec8�^|���͉�u},�頏�/z=��|�;7��^���������mLv�(����;  Q | ��{ƽ|��.��d�xEh11�قvpIY�ctr�R��􀝻C�x)5�N���9ث]�nS)jΧ��bn���WFia*�,�p"q
��%��;æ9]��5��L����QU�Q���w^;�=�Q�Ѿ����IHC�y��9�OAq}���}�`©�w]{
-�ہ<�d˫P�e�&�	��S;����qP)�GJ��􇻘�H>��#|c�S���>6c.�t�t]�M�@���Ff=]6�nT.�b�
zz`5W��U���l�z����k|g_J�dA@�D@���1������:��q��Yl�����G3j���)M�����*e����N����\m�M�O�O7DT����Z�o[K鎟�z(�-��V��}H�uG�n�R�����R���Y�����1�o=���=4�R�NڂD"�0F0@R("�cR� "#0`+EX2$�UV0�$E�TdEdX�+dFAP�Ab��(�H�P�pk��_��L�޻��h��������}�#ZA<��\Y}9����A�w�%������z��W^IG���O.���g^�P
��>�/Z��Z�5]+��n�W�T���!=�{�t�	��&OO${����3�X�"g%T�L;4�ok�ع�C���6��4f+��CU[�[�� +�^g��NO��7�b���^T����C6sB1gzTM��>�D�|TZ�Tn�h����h�2�������]�v��#ᵟHxky�s;�����s|�&�M���o�8/{�VWbjy��<�k�ӏl�G�y<�P���z\�pܣ7�)^��m /gd3h$�,�g����%D��H�0��j!V�H{�J{���d����j��V�{AA"�X�
���$���2,#�(�D��1QUcV1cA�*���� �>����S�Ź�: &����c��a�M�Z��m��L�Ӑ���I��h�EDA{g�p�V_l�u�;�>G4ޫR��75�U�-�.���S9xTk��!�r�T�C���wnћ�4�m�ժu.'a�W�4<OOI�n����l��eUaTE��	kcS=�;��ʵ	B]fl�a�<�N�����}�!Ժz���A�_Aٻ&���w��">���DE��ѝ���R�]R%*�d���7{���}�G~�����<`j��u]R�.彩�Iv�*�k�����T6�ڏmR��٪/�U�eU����=���'K��ۇמ�奔C��@�}jM��bj8{�z�l���cH(�R1���X1TQ5��k���gy����B � ���d�*���޼֫������K��R��� ��2�����CvmC�X��;��א7�����;��ݰn�ܝ��Ҟ(S�s�v߻�o6�Gk����,����R:�%�]�]��̟t�:�^юS��=���z]f�6ӡ{_�����;m����U�{U�W]���O�kQ[L�=�N[�a����3L��OA�4e�9���~��T�?v�w�����x4���ń���oX�%����޼
���r^�+_I�u��������_M����t�]QCv�8�*�g�{W�̧���\vlt��ϖV�>�騲b��#����F�vN4�˃����x�Q�(vb뮔��'�'�����β+ �@����/<3�'�Zn�߽g�E��(�C� |(W���G�-���^��ϗB�����<�^���+6qt|b~����̌�٘<�3���
Ǚϕ;���ͮ�q�&�]d���UGo�:��k����	h*��i��ݜ6����qM$$!���L��5^Чz�-=�����	aݡ#=фW��z=c��/���f�]Z��S�(t0B�pY�j�s�#/s�vγb/�̌�:j�Ԅ0�R���"";�f��q��N|�:�*��l�&̜���l.swJ�$ו�p҃Օ;s��(Z�΍�dI)(LR��%(�{suJ41h��b��*$�\5�x���{�E�ռ@W�{�T�fb�pvL�Y;����ոgݺ���Ǟ�>I$3 8��1-�(("
1E"�Dd�d�b� (��p���w��v�qf�Vk���<�^n`�"�V����/���l��.¿�j69_I߲O�SɆ�I�I@$=�V}����0�y���y~�ݼ�j�`��;6�s����,�H���~=n����b�|d�_=���v`�xs���k��gIY2���л)Q�_�0ƾ��|��x�������M�ۙâ)�ENd�k����濸p��t�����ZUx��D�;�N�}�s�w@i�@ADX2�U}������<}]�ŉ�H5$���W��2��꒳f��/$����K7Yk<�#�ef]y�듎X?_�� �L�!9����O=����;����5o/9�c�]ha�pƅ��e�դN����}���;P�>�� D� �DU:�g�Wn+5Y�c׻�`J`��7�=RK>�9oUj3���ò��S�����|b�;�����<�Գ 6f�TTM՜4v*L$��jD���f:��*�Ak+��R^4��ek����2on�r�Ҩϧ� q������N���PZ���.��\�'XD� �:��%؈�K����a��ik=��j���l����r���r�Pl���v�t�Ѣ��˶��'+{h��������tk�U�A6��0��:�;�`�]N��ۻۧ��yyp^@^�5]i�����.[ �_cA6�u���(�X!i$�B���0C���&�#�<:�gfLxEV$�R�7.mn�D�s+�!����}��*�Ф�(��"�P�e���2mA�֑l-@�Ij�����u�"��,��Dp�N$���֩��3AXM��I�#3i8�wL�2����o+,�Cy������c���p�[%�ܜ7( Q7|��$���}�$�[��b��O�k��&S��I��+Y��op;ڕ�gGu�����lBi�m0O� �@�U�m�@)>H ~h�=R���(�B��b������E�(��AF�ے��"�A�zڡ2�r����D�%�,-U��b;UE(�*q���5��j�,���&��	)�����`�]���Zgꉖj)�(�\���\W*�a�w���,��v��$���\�{s/ �B:�9��JnPі��L�i��w�n-�a֌�T�uJ��D7WtZϪm1KsL��n��gdo''�y�}��CQ�Xk
�L���n+��&�����-\[}�Pn9�)8��_Z!GvGuL��޾����e�{�G�n���书nf�A�(��qs��]�^݊��ɵvZev��o���P����B��LֹD:�*�$`�u�KU�ݚG<�Y�6�ն��{�����(ʗ#�&	\2������W�&���Ӈju1HP�-M�лt��\.��[�buc���ҏ3p�WX��ƺ}�Dx,ҝk�T'3�f�I+9�Yg���rv|-�๗|�I�xk���� W5D�ڹnc\��vH�2��u�'(�f,x5\�c l�t��<�7�Χu�+������dpno�jܓ@��[]������[�B�Z���Cr�Ԝ��]�oP�������sק#G��O�-�c6Z�8H�z�΋E���#�o5�V�û�[S�oG˚o�U:�L5P5(�3"�õx���)ރ�1	��
�pa�ŧ�n��m�oû����ekTV)q����	��K�'Jk
1����JY�{3��a��T�h} ��!��#����>#�/�\�Y�p��ب����k&d+9�R�{n�,Uuf���F�^i틷�g����v�Ѩ΍S�٧`n�oV09�g7��a���YeEƃ���n=ī��m��h���%V�Iχ��+�r���o�{�d�#���e�T���~���"��ca�����6��6*Wt�0��WhiIU�E��>���	��Y45�w�bL�m�6¹�q>9��~r=�@��B�<WW\s�z5=����=ß.B��߇������=�F��+�>OJv+��XV��CE*���Fv����N�҃�4e�u��D�Ş��e��ӄ�"n�O-׻�Akݔ��I�m���.J�ٺ�7�a�~V̏k��ߖ9�]ީ7�sM�����j�����}Փ��^��;�]��lbDF#�1A�RU���C4�����s�2��H�t6�^vԈތ��:ⱭzS���S/��+�Ȇ/�rnؤ�uf���R�N����U�:�u�ݪ� >��3�p��&�����f��k��bsE[O��Y�l�M����	��3{8��X]7�&c����]��!ɮvl�k:�k�6U����zZ�>#���R"3��}O/MW�O������ö���W}�dR�3wi^���7H��@T\��liC�m�po#��㜹���#6��-=���|9�9ʍ���뵝�LN�j7�N��˗�
�1�d�u�@��ZM! ���U���ٛʸ5�WD}�"tp߫�>�PAa�)$�Uw�
�*�H�I��$FRF	+�x�~�^���f���w�7t4h�2(�*ge�l��v8ɉ;��3�hi����<�uйL�	]u)���)���Q��)�L;YQ����G�3R�Q)P�_v���R{��ڛk>m�U���~2�		�n��f��Ò�HZ#��Ŋ=�\��;dY��@v���Yp؝&�W��s�����썹��j��3����]���r�$��RI�-U�(}���R�z����<`�P�b����{���5���y�7�=8�[�]�V<�p��6 ��b.�i�["��}��qٵ�j�.�\{�X&1Y0��V^�V.�K�x��k:���:��.M��Y-]���8R@���e��m���1<��oc�ڋd0E��UE@"��;�1�s5½]�uj���DC���v�:��n� s�9��KZ�)��ܔ�T������=��l䶻 8m
l�s�qec�T�l%3�[� o<�9yRXO��.�>�fG��v9[F^<5��}<��7�2b��Ҹ�J�v��V����՟f��{�_HN�d,b%b�,EQD�����QB1�cTU�QY"��б��"��E�Ȳae%1UQX�.��* "1A`��Q��UD`*��U�b*�@dX#�hw�ۗ�eZ� ����k�{��^cL�3�@��u�4A;;2ј��O��ҺCiP෌u)�.a�i{��*��ic��<�.Z����~�D#*+i���;$w.ዎ�blFVX~�<>�.T%J�ԣ�=�7�xz\�Y����X��l�������=<Xn[=N�Tl��u���{D�etƨ�
rL8��ץ���U*�f�p]3VoP�����>�1��%\y�@�B���V
 ��Q"�`���(}B�Tٝ�/jZ�ݡc��_GK����8תzO����.y��4����T:����o����֩Yq�69�'�U������P9F�k���Z5Q؝RG_'�bXs3������]'�^Q�G��Cq׫uZa0�gYНL�L��X�A$=zý�V��s�Ϊ��N^�Z��AI X�޴�zƭ�q���f�m#�Go�a�Wƺ@7��^��М��P�uq�B�W],%\�(���)JJX�����y�W�����\�h�G��o��Θ�S2�g�Մ�w��T���Kx���}*���E
����Sޥ�F�Au^���9%Ŋ���%��_�Fܮ�p<���ݒ*����P`��	���������;�����X�F#b�� �`o�����`�PQdDUA�y�c�x�����W�ԥ��x�Tٍ���E�ǻ��cS̭�֯T@�h߳��4�gKYV1�жJ��"�S�r��]�'TkU'��.C4��M���Y��q�.����4��C-�|��[/w���w�q�
k�sX����""�\����EUjͺ�}mA�Δ��P�B�1�Z�m�Zp���e,$�}���V���W}��{�v��l6ު���W>v�] ���t�\q�θ1l�WZ7��.�8t�\@�5e9`�GS��3p���%��׵iXW��o5�N �wCj)6��5A�5��a�b��p��|����=�a��V-��p�L�-ƹwp��DEQ�1��A�Q F�ȠE� �����)� ؽ�`g�}nW-*�R��l]�]6rũ��N�KJ+�`�k�W1[T�+��r�^	s��bye�G���t�Ʉ��9[K&^ƾ�zP��ʼ;h?Kbe�Y�ٙY%	��X����o�V�>�p
&��]x[��w�m�/�+� yؔǽ�-���:�]��Ъ�f@��z�=�YL�r˜7��-^��sV@k�ߏO[����x"~}����M����5U�]us鹚+c�w�"y/�T�e�fwe�������m2��EM��t[ԫj�묦���o��]A�-���O�2z�&�JV
�^̘���6��O�eM9�U�����E��h۽��{y*���<�s.M������0�V"	$���������b�cX,`�y��x�9v�Up�}� �51�.A��}$�]�~��M��P*�y��c�v}Q��m���z.�X�ˎ.ڂ�l�i�S��	��y|�z�u�\4�enh�v֯�&�,�w�"�>!�gF�^��s���!L���G)�}��� �#Td�yO|�s���kǻݼ%�4��8;9�u�9m�k����|ѯ*O��Or�������D'�1_}�cMW��UV�珏_��[a'(_y�geK���NLt���K���d�.e��åok:�tpwk���
c��٥�;��nu�����<X��:,w��U��aw�8Tr�=��6�Z��c�ks�������] ;��E�uꜫ}�L�����K��	1c*,X1TPE�TU
Aa �P$��x��r��஻�.H�y�����GM�a���7{.����1ъyX�PŦ��cq�`�����KV�3�ؼ
�Ձ�X�έ�z-�DP������0�f@���uqT���	���b�>D��E�ȗL�w��Ρ	�L�9�},���݇,��&��j��Ȕ��D�]c� �����	L_��_����Q��ùA�1K�R����J5�b�(�=��\��/����Ln�d�+�Po������/?��@ ��$|	&q{��L�J����X�&�n���6"7qк�Wv)m�`N�J�v>[A��䉱�Jt�B.hh
��_Nܨ���Rn;��=:v��ԧԺ�����˼m��G��� �Ab
DQd�#�E����/����|6^�����">���'��v��9��m]g�����!MS���!��ݛ��z�<1��2�wb�i�EUv���\Ы}Ց����:�iǻ7����`��<*����i�~�&�so)B�������=��
o��y����p�w6��`�AbE�0���k�4�9��7�fu'	�t/h�m�_�&�:5�m��ŞOwm�4S�>7�^U�ħ��(��VЫ��b��Pxf��I���<7�H=Kԋo��Œl��s�(�7z�q����������1��2�F��-���9ɡJ���On�,<�7��/�֞��}�+o��cn���K���ڻ�Ƕ�3�9�f4����ÄΛΫ���U
�'+ʻ�����Q�|n� b�c����]w���"��QQ� +VAag����D��v��`Q[�Co����I�k�+ۦ�\��n�J���6Ŏ�]<S���|T�v��[��^� ����eo�W|�'���e651�<����+pLt-�ٶ) XO;'WfUw�Ɯy��Vo믇���w�l�#���/6;;�/0��-ܺ��Kdo'���B7����۬p굸���oV�p�'K��S��N��Z9��]�r����@�θj�ô{����/^�vx�8͸��s�h��5y�ժbp�ɜr�W���Lk��y�� ވ�*Ҡ���������x|�U��AB��!f�\	$ ��H���>�X/!Q8QQ��.�N��S�y9bY�ˇC}'^�Ԯ� @@DDkǯ���U�∊*�v-��;=���wDQW�,���i ��|{�(F�q6�s�DQV EAt TU �q(v��"��kqueu�R܎X�"��q)�*���m'�o�O�|�EZ�oyi���tE`U��P��*�o�TEnM+��}�+BՏ�	64&2�0I(���m8W�7��DQW��J`P��>��Vx�DDQV���E^v�;W\Dl04���8���Ю9���*��� :�Zs��uk'�Q�p�(���zV��U�w�l�˦��?��e5����G��� �r 	 r}��D��T��i�T�!z�ȵ��[46bR��(�RT�Rlk5K(�̋[mM�f�B*L�V��늫lm��P��a$Eҕ�@R   ��,mSd�-42Fl��Cm�L�[mB���M����lJ��bŋ5���c+R@$��V�ٺ��;��jcDڳ��<�;���Z�ʤ��Z�{��h�{ϼ�G{W�Z��u�O�����w�����n7�� ���t���z��wz��}x�|�/w�c��xWj����w7!��ϵ���[[���������ޮ�d�d�lVfO��6�>  � }
 ;��    A� P   �   ���,_=�:z�=��S��>�}�x�����}�o�]������/nng�����}7t����>���Wla�s�
WAj���R>�=���o/N�����������{��� ���ﷻ|N����������{�qǽ����lI�[���|�v��{���]�ϕ<���s�ڽ��z��b��t�)�.���������4�|w��{���{����X{�����k���{��Gw�=���U� /��y޽ݼn����ǨT=�w�<�{=�ݎI��s})��8� q@P񭕳���h�$jy���(�w�=�v����xz�=c޽y�J+�����w&�Vs�G{8���������{���ǰ��=��vy�t���]i���۾���T��e�y�=�u�c&�<'Tbݸr��^}������/��x��Jm����>l=�^�n��nw�vS���)�lյjڀ��-5M�	GC�}�{�c��u�u�n��w_A�o#8w�w��F��{���'CV=ÎǠ�wW�'F��áw:�^�����n�-}�J�#�la�*�b��F���Ǯ>�y�ý��9��^�{q^���:���<��`��7v����/=P��O&�n���Q�gG{��.㆙����<�޽�A��5��B�6�b
i�:�廳��˧E��x�ﾞ�����}Ϻ�>��}rZ{ع^��t�<�5>7p=�}�^�=��.2��a��z���wﷷ_eq��=��^�iL�QL�Q,��n�S����3�Ϲ7;�����y���q��۾}�N����q﯏t�㳫]׸�9�G�G��9���Ѿg����|���5ǳ���˞��}�]j}}��| <E? ��J�   EO�RT� A��S�2�*0   5< RJ�   E?j �TѠ   �Q ����)�20b~>ߏ~O�>�߉��w���j-�c�/pU�Def��X���<�l:�����H���$��K!@�C��I!$���BI*!�RHI	$�j$���KBHI'�$$�����ǿ_����Y���o�l��������V�J��֫�2����#��+�ڙ%ѓ)�\��o�N��ՙr�h\W�Ĉa.���-*��F�27�m;�q�9��rV�̷2��-mD�̼wQ[��}2KC�fk����N����6�P����U�wg_\��nr��i.���u�&L�)atT9��v�+uM7�l#oT��5}#ٖ�t���3y�J�콖;sXt���FRi���p��eBo7(2&5Ӭ�)��b�*7��1��2��2#���,�)4-˗��k�\n�c��m\u�p�$�Y��rn��Np����;f���)����m�z���+`�e[sܬ6�(ut��y��Ԧ�WY��z�
KrwN�[\d�9%z'�&v��wZ��pP�Y���,�{M����t��n(�س�〨����-��+��
Gy\����eI,�2B���q�x����֞��,�׍�z���t��Xc��ۮ�aō��C��P�,�u��Y;�,��wi���P�%����u�Hd�ʣí�)�`�M��kCg*VV����h�O=�u�m��Z��U��^Z���Vɰv�91H�w����$�}դsG�u�C��nK�ɦ1�vzOgH�̸ߦ��ӕ�"�ӭ����ᯮ
O�1/��>��ݗ�U���8�1fۜ��K2������V�z�T��>�����csy=�w}SjĊ�ԩ��]�7*�o`mP�*霺K����i>g�òi�>�/�+];/4B�"���>�ܩ�2𬷾w�u�k�N5��bշ*�,���cw3�k��w[��X3�	j��C�Al\A��Π��EÁ9V&I�zZ�Wq�J��BSvVgZ9��Gq!H�6�a�-�7/���xn#����u�A��(���0�N��Nd��f�&�3)5�[�g^��fS
w!`��/1�5���!�O�n�^kC�0a�υ�d�t��#�h�rwծU��q)I��,&#����U��%T��R�GYI�h-��=���`^3,�Vf�8�9�-9���oDdu�i�M��Ѣ�&:�Z$7z�r��6ŋ[�V�Z�m�#���黩�q��1S	�+F7A��jL�&l���oU5�M`P��.���x�^�jL���|�`	XpsIoG��e�����ݷ· xuS��ҝ+�}r�W������4J�i�jWp)/����y��S#2�_H�_��E�����U{hd��n�и=$|[�H_N�����#�qc�ZV^�/`�i�n��U�,��!TvVd�0*��5Y}
t��l�ޟ�f�
Ɩ>o�YsQ׶���0�������Ո���I�3cqmiB���;��M镵ᆴ����V���X�,�ܭ�
��f��t�ܣ���W�s{P�̨��Yӟ]������/E.,����-Ѡ�J�����F�,��^���o5Ǵ���ҼG7�vi6��"�n^X��[L�K"#�8G,��*ݗ՚�略�$�sl��ݭa����[q�=u��rͯ�.��x,�U͌[XM�������k��U,�ǚ���W����V�(���Va��s�7���_p�/��j��@b�m�]�Gn9��ݕ��A���u�|�J�*����
�.��y����Z�X�t���/��)\����#/�r��NZ�ͺ�	��b��<���d�f��$p?[+��U͙���4�ԑ�A����5{�Ÿo�<�Z(��Kk�.d�e.�릓�4�۽����ژ�U�K�SI�6�E�|h\ҥ*S�B�$���kݬ`ӇE���"M����a�K��/w�e��zIM�����%a$ˬ̡H*LI[,
��Hb{]��ys!�;;{�*�l��c�m C��$�-1�ẹj���[�G��l�f6��wjyce�uܚ�VS�'������^dY6B�T���trZ6��y(:��U,NkTˡؽ �C{��vfbr�!+R�c[����T`�]:���Xn����iM:�$�#s+�y"�G���b���V���L���Q��D�Ŭ�*
�>��f��CL�M�!|�滫�\W8;<�ws^��6�\T`,�([����ڤ�5��k�ҽ��%6���,�wI�g~6���(򂁈ww�����)e��7�-hae�T�m����^���=c2�틣f'3XE�w`�+2��(�ȂLV�n�&��ܰ��e�ul�w/�u��fX�$�L�V�I�������Y4��ި��H�R
ޓ��O�Jak�f*��P5�aXiV��r{7q\Ux���PHk#D�oAU��y�96lڶV�uf]�p���;<�
3 ➡NL4�j��T�jt��smՖ�0�*]O-�1���.��ۘ�n����������ە��T����q!*�I��b��&��Ս�A��*�R�CH�٬���4�� ���@�I�Ïr�Å+�96�֊�iX��=�Q�XĂQ�����l#��t2)1U:��\	��i[*3�ۼTKq��	�w5��˱��M:9�EM"���VN���jO���hn���÷�7rf�Ȭ��Y3+3�ݵ���4��0�5&'�l��4V�vj�;u�Z��m4�Ik�%�(K�i$�G"�ݚq�*�LW�hN+ԑY=���(n�vu却q�A)�ALbGL�;tcuI�ؒ!����� �K�ɵ��pY5[[oKʂAvkm��=�w��H�k�r�\�Gr�� bʼ[��b���3*i�A�CW,�G�B���pV�K���.�FB(+��+���K�FK��nǸ��eܫ�3�wx��{��;�L�J�R1MY��Qa��q��F��rPYCf�m��6]�kb�&�a����q�P[Wh��4�\YSD����P�H�Z�PY6�8D��P1�73t֔��ۃ(&O1���@S�C-�&(ksJY7=vt�&E1ʁU÷{p��B�j�ݜ�5B��v��lM)���f��5Ir��*A��`��T��۳�Ǥ��Tjγ̏E��/Ml^����+3���jӵ&Vv	U[�be�&�����V���u�5�%��rP*M&� �w�;V$��V��l|.��=������tz�d�jv�T�8V.�}.й��V	}���Ǹ�Y�����eA"�R�FSfl��p���_0�T�e���=B'b.�ǘ�v\�n�<��8:-Ҥ�Uݖ�z*�\;`S�T��
zsz��9��7W���'pa�h�\����Ҟ�p�R'�fr�S��+5�h��HmU�^U��2�W-��8vt�Mإ�+�o�)m�N*���V#�/�3��D�+?�����)�R�w���nf$�`���W5��������h�[qrA��Ֆ&��IӔ�nl��S^�-)����,]�En�|h�II���I�����2�m��j�1�f���*w*(eLjNmJ���o--�{_W\ފ�o0(%G/I��ø�[Z^��$qn�\t2	���x�oE*>�d��,�׳C��őn=��{Y��w1T�+YU�ԣ�)�4�WfI���ںmf��۸���x�4��ΰC�h��5Y��
��eR4�XP=��Z�[qJ���V�`��H�8�(945RۻWi +Y�l� ͧ�EP/l�noK�bG1XKr*r�F��*´��Rݗ�.�5��*dVb�N9���6:ʲ�����.M��)m{s-�b��/��<�e����4��(2U�U�D�jǯZ�;�Tf���4���, 
�(���c#6,�`��(�U;b����n�In�$O �԰v�ݝu�XM� ��Ӷ��T�-��Qǹ���'�7]zV�P��N��� \2�d�	�}G�/F�_�F_	�b�|���4^X�E$�b�B���V�j��bV��m�v%[vs��(=�X����0YwvDOBy��VBsnjk)�	[��tLNj:�h%mXH������2�r��+�كb:����R��z{�(�̸О��$@^F���"�1U��?n�}���Y�髼U�%�\�޷V�� \T�lَ��Qޒ��\��1� �Vn��%�5�P�9��-�9q�Wb�zr��45�����sq�<v�޽*b#�i��*�G�W��.[�(�>ު���'�R}f�^�6���j�u�H�n ��o$��Ur�N��,�H9���*�,v�L�%�2�
m�t��T�*����h�*f��k�[�]ӛ���V5��3fe�/d�H��VƷjI6�v�՛s����fv�rN��GDm���]�c�Kw4�^
��!�qF�joאD	�����%��x��R�$�,>>"(2����[�#N�	%̡��{�2��s	5�soo\�h�[ņĽ�F�?�c5������#��q]^d��J��p�E�ۭ�X�M�a-��ٕ/-���eݼ�)�z��Ƀw
cZɴ�m�v%
ZM����!��H�̦ek���MX��3aYzN�>ߣ�s.Չ!j�����`b�VF��!�u�ҋ!�QݨN�b=sZ�V9(��6N��H�4�`��R��fXgnrLnZ��IYX��'�^0D�űhy��"�O�kĀ���f�n�2�-:�q�Z�8E	w��K�&�1$���S3,�>����.�>�����SBM�^Snk��2X�$qյT�3�j��x�� Y2%}�WU���o�7k��`�U1���Z�b��V� *6W�%���tk�̰N��I��JT:3+fu>�]�b +n�lWg:�1lw�>���"5�m������f[DYÜx#��%�lUE�nt��%>���K���Ԧ;�CL��Ju'n��@�:ڛ� 2bK7Ԕ]�����fCM��ib4��[��ƀ��[������cr�6��Y�H�tF�l܃V|@�uG1��vs�ZHm!����w/�C��)�(��defk��jR��d'kI�Q�ZC�Re��s\�l�d㱓��8C,� '�����f�G�B˩�b��F�R4%��I��oN��������v%�ۚ]wxi��j���[&{uv�
v�CN�ĬZU�<��佑&���dF������b��tZԡ��Sztby�X�N�����,5 yF՚|�a�7kmW>/r�F�ģ*f�s���鲦p�L����?$���n���d��(�V��ll��yM:��۬y�n��Z�;�[�.n��t�qK�U��T�e�u!y���
J�M��m�s�U�e�¥,Q`m�g����.L�f�*J�I�ebݺ�X��.7yd�<)�C��y4�+��$��9��f��B�{A�`�+{b�� �(jX.�`S	��ٚ��7*��fX6�����K2�VXT��^�d��㵸��B9`S�#Sl�L��IY���2��P��̐5,b���]�5�ѱwd2�ɟX�0�j:��+)F�^�k2H� �E��J3!�vQ���vjڋr;ː^�Z���VP�3t��Cɥ�����7h����ښ�Z9B\i�̎��V����lfѽ�����L43+0��!T��FzC��Y�d:U�flY��p�չv�L^��ZLj�b�Ba�yX�bXu�v�d����XX�q�t�n�b�r.!����v�{�cS�DwU�B�L&]&�$lAy%$�)۳���`�׺t=��4"4�j6�����Wc��פ��i�K��`+D��Bv��pnu�F�h���ٞ&��^�qD)��F��w�-�7�X�\o���[��H�0TJ� p�炞Zf�-Q�e��K9\,�N�n��Ս�I���fY�p�S]1���/�U�;����u��Z4D&Kλ罷�$p���Sn��bںc]��j�%�v�7�È�9���:�z��5�����HP�j����5��ǮU��5Zl��1���+p����E�v�0]A��Ԅ�4tmt��N`�����f��=��yۮ��A�`��T���h�9Qo��Db��*�ha�4��VXU^9k.��J>B-��ј�XmP�`�Z��M`*0�3"�5��3w��6���M�Ú�Ccd�LF���"�t�!dl�ρ y�U�p�"،^�����Il9�N<ͥ�E��d����a��:�fl��"b)��c 6��nk�m�ن�p�b���E����0	A��\�6�ͺs6����ӹ�Kxv�������{ ��I{�U�`B�^P#+veXkȲ��j�U �������f�JSB7eՍ��U��f��Bhy%nl�qnn� �^�>	��P>�N�P��J+�6�[�CIzH�s2U�╝:B��t�*��U�������!��&�hU[Rڽ1�Kf�P��2-�i��jSֱ��]����Ć57Q�t���osM$�Ԍ�+���ө�k�I�k��/T��`�ưh.��V��ʍ���[�����h��6��Z�Ƃ��d:+l�{v74C~9�1�2ĺ�T��V���a�(�&�dڵĞ��^Z۔��med�k1G3n�v���0]k�|�v^�x	wՉQf�t-,����t�fK����e�qn��o�G0�M$�ɬ�q��ڙ�K�7$ܽL��+M+>�Wx�G56-ӂ4�rXk)��򢤈�0[ٻA�O^�	�BJ�^䷤�ҫox�`T�U�l��r�7(T��iU�p��� ލ��`�
/3 �n��b�
A�dfm�l�2�k-{�CtI�W.:&��ۃ^E��+ �Ǖ�cf˦������.l{WDY"nH���|���ɢ��"���mM7�X�Vi�l�CV��e��X�dܒ�Q�-��sZOL������Z&ip�	�St�t�0���)�DG�ժ�RE�4���Z76
��$֖d�X`�ƕ�2��Cک�����f互	$�I$m�$�Fې�$�I$��ܐ8`�I$�F�rI II#�3�Ddm�$�I$�I$f(�m��&I#m�"JFۑ%$�I"J6ܒI#n�iG$IBd�0�Fl4��$�����BdI$�%#IH)$��ӒI$m��a�ӑ$�n	��ےFHj(�1$IH�
I$2@�T�I"�Fے	$��	�	 m���$I(@�q#m�$�%"��$�$�L��$��[I%$H4�h��m6#h�L�InI$�I$�I$m�m�$���a��I$�H��I$�D����$�IRI$�D�m�$�HҎH���ܒInFL�8$2G	��n6܄Ĕ��	�InInI �Bӑ��I$�I	�I$�I"JI#J4Dq8�@�I�L`�bB[>�� mSh��
?%��H�m�!�BZh2�a�l8Q%�I�zOK��d $4�" �BP�#�(�K�Cb)�#-��`�0I�i��Q�g�0��l��L�@p�$�4�e ÈF��BOƌ�Q$h�J1�� �a�����!x�
,�F8�"���!F	?7PQ7������p����+ɺ4͵��}��c\d�jmR������i���4!M��v(CW��K���|�8�clHBjKO�$}�H���f��!�T�ҥ̤��(*��������;�D�νl蒷�T���ٵ�Q��NQ6D̾&�Rc̐��(�W]m՘�����֙xIq�vt�,���)�Ko0��S��e�{R���H%�
Q>�1��9o�Ƶ�)֎���5Y���U��$�lեb�͝�zH�ےmJ�θ��]qE��Vc^i� ��.�ξ��x�����[W�9��XT@�í��y���.Bl%}LX�T��F�.`	��/>C���x�nR=N�2nU�#�F�!�
ܚ�&;WN��Ѭ%�D�gb����ݓf:�h�/��Pq�Ze�йp��)��G2F��vfA ]�5�S�R��\cy#{.��1-��u���"�q��'5vL����fָmG6��J�v�{�3D̺]���\dZ]����/��3{�Z�r<�.�8�H���i��t�۽w]�7�7��\�aiG~�FcY�]ګ��jd����(D�H�{�;�����z���TJGT��K!U �,i8ZV:���mv�pز�p�h�,������V��7.�J����%��F�Q���un�$]g�f�����w���Q����Q���9���ѫ�+���ԧ��b�l.�O�H�gjl��cFVA��.c�~��=���g�z\����-���T�pry��
��[W�Qeꤷ�H�L8M�!;e�H�v�7�w�w�ze�8�H�ܫ:���F�a�#�jƫҡ��������
4!9iWX6�K�)�6J�X��9"�K���F��TE�*��޴Hj	�Ex�dYB4I���������v*zX���0|� �b&��Y��r�e��z�8���[\��[�}������us.�s���!ە�TY7KvA�S#%��S�.P�.�+܋p_!�V%D�1
�:�m�p�-f�])�e��������gl%;���i��A�]vp:�&�فN�wI;$���H?#�̱�4�|�+XJhw�mv�b�Q4��Rg�C	�"��{R�w[�I{�2]�%q9MK�2��I� }3T��n]�X�/�md訥�Ǌkׁ���QҝWh�@����0��t���������+F��7�	A�1R^�rM�p䧨	�y��!�q�0P4n;07\v2�8bl��}G���m@Bv�ݴ�vmh��Fc����Qc���hQ�ۣW�e�vA�AUA]+��mN���=xB�L��7�}XSŷ�zt�*88�x-�݈��]�4)e�w1�3�
�d��yu�e {�1+t�@�@kj�2.I㥳�T�u֦�3:��1�2���É�3�J�>��통\���Ϯ�ly�fkq�V��e ���ȥ�tU����rE�����);w9�I^ud��2�mi�}��V��6A�:薠��n"��к�t�ʬތF]�a^�/o���PR��zY�x��T2n�<�΍��L�z����� �t��EvbN�nP
2���	n���z7�6��U��>r��E�!U��<w^g)%ϴ�3�Q2k�e���.�v�\�.�b[�G1#ּ�%z��%�w�T���td,-���X���Ƨe1]��h�ԢOG���8;�5:#wT	�hK(°oVc\�Lt���e���V�w /+ �D(���zz�&7:�G��SS
��L�O�"� �Zɶ¥:��sL��e�$�9s�fn�T�2"�&ޘ�U.�'�����W+3&��ThOsI��oa`0z�N눁���e�y<y�z����E�8�h�������R���l��O����^5�;{%�r|����[�;y[�N2qjho��GMZ�o@f��Op�;�9��ũN��!���mn�O@�I�^\$���`�2���3e��'2+����r���=������1�#5��7��z� �+!JӃz�(a�����b�E�hÚ�E��+E�E�y�c�\�嗔��K���n�%�2��t��,�V�Q�Y�!�}e�6 �Y���ʃ �˰�!Ǳ�ʖmO.��m�uȉ�©�&:�ՙK#�9P_;�`Gw��>j��p�� ��^j�=�D�.�O1Z9�ur"^բ1�2+L������"���0hL�n�r�<X�7���L�'+�j�A2�!mD��E���!GY{f+4Ɲ}bD�Xg/2��!m&�P̠�;΃ddi��u�#c���^��N�f��)���B�n��>���:�,V�K@��@>NtXx�e��y�-� ��쬎m��냧(rT����B{pŶ�*gv�C9!����u�8�4+�G�F��>���Y���
$V����k�9��n錦����3M����Q;����g�vN�ڏ3"�!.�r��3tgd���sI��3�/
�f�n��ol��c1bZE����b�s�ͧ�5���k��s�4n����y�l����k�	�@�1�0�-�b�e
p����������!Lf�ɛ�u��O+#���m���5���3㚉�3�[��&�S�XΤ{vMl�8��]�WPݓ�LCh�w;�	Ȣ5���$ɑv�I7���ښx)x��n��]Z�4>��#""���33�m޿�a�Ǵ ���ӕ\e��5�[jg\��C�C��i�"�0�͒��cp��`���^9�v����B�-�h��k��4�ke�5��l�gtQs2�5�.Ȇd�Y�䊧m�遪�R�ܚqhh�h*,���@�=�	T���6�h���Ǔ���QM�f��f:j�7���^5zn��R�r8���f&v�l�:����)��v����b�K��#Jng��M��s\<��Cǜ�C��
���#�U�Z�A醃�Ȓ����W+�S����J��9�JU���3f5�^i�lT�+m:(;��'@s���a��B��W�YFk֔�ގ�N9�,�˚����wV:�*(s��]��D����p����آ�k�M
W����;�H�.j'�,�8�{�`���
�E..�$j�sYn;+%���X��9]�bx.�\�+n���9؊��#LLN�R�֑"�uѸ$��3v�C;��Zбr��PA�MY�_WF��C�&^xe�%��T:���b>�h���AA^m��w#A��J�r����@�*!�\��J猌Ǚ����.Jոu��v�cKIJ�<��Oȍ��v�B��fep�=R�r�LlQ����[����cI����ʇ3�`�P�_P�T��x)���L���-+|,$\���c���L�"c�!�_��Y���Չ�)����B05��ǝ���.ŭ�Qbu2�.4���*�.���U�Zc���Ό9�a;'nt	역��mКAf�ü�G�AM�P/e^mk�N�ly�#�b[C�[���:G[¯�c�ԯ��:;D=9��9	;:��}w��pZO��, J�����N�2D�YGF��6�*�->��W.�Mۈjs��Ĭةe7���T�骝_"������������0ݫU�����ȃ�����L�!���ת�KF�b�M��7X�n2��W_�B��j1�W��֧�����W�1d5w��'U�l�q��tQm�{ep�	�曬�l����m����4�,�*h�[��%)&RUԻjѢG_���f=8���3T�A���K�j��ҕ�\|1piX­�\W[;ĞhX1檢���Np5,�D��A�����1���[�]���A�X`xQ:AU�{3ve��$���dJ@��toI;�f�S,n�φV�%SU�M�ؑYͳU-�y�C��t�ja��8+k�gC���	N,J�Gd��A=b��͜�����C:�D��S��=�RKko�S�]@�RH�engU�%�s����%�ñB��"��ˍۑ�7����4u��{��o_k�P����J�1�8N3J`J����hگڅqKWP/�Z���rA$mٱQ3�����K��R��E/4R����q��d[h�����l:��O'i�2�g�po6v&B�v=0Ƒ�Z��/sP���x���Q�欕��ّ����W|Α[L����y�غ�Uhb��R6�L�[O����b
52*����a�;�R[y&�N�i��xtX'Է�Q��[�ث����ӑ�_n�����V�koa�x���.B�-���d[�8�9��X���F�E�uی���~և.�zư��z�J;��(��d���JyC;8F�&]:yK�����]���}Lq���嵜�7�$�R2���k��jۺFq�B�A}HT<��cEh�����-���gr�\ʫ���ْ����ň��3B"��r�z�ƙ��;�KHD�L��y|b�0��ʕ���8R�&�=� N#���vN� �{���7��V�\F|��٭ކ����9��plh6U�,��,"�F�H����im+����왻�Crje�a�5
Z�Y<�ӢE:���J�[חx��7.�ͩ\<��xE�gڣ�_S���k�[z�n����%��������UU[rlU�<QN��t,*q�Sw���`Т�{�m �⏈Z�Uw_<U�W�e�o&�҈������{O�G0ɇ*�80��V�����{O�m�*4k�'m���e�Z��Я���H�Ls-�t��Y������]c��!H��] 7�
Ҳ�pĄP�ɤw��G뾔��Q}�t��X��;=+r���k}�vN ��ID$�@o�f2j�3^�q(�U�3J������,��Dc8�p��cq�A����I�^�)b�J��:��rH��%x��	f�uѬr��}�M�oX@��X&�7X���3A�hv���n��c*UM����"��.eRgb�RD��w���%���j��:�o	��1���2���6!�WK�ݐh�H�Gwr��e���Q#Z���ۖ3`]a&��6h3([лh��V
�-
�����v;�W(���!鵳v�`�l(�t�ݽ� L'UH�u����� /b��6J��-��Y!quiy��{��2�*�Gn�p�=��v�>�\+4��a���(M���L���P��`i�9-����Τ5|�"(����p����˴nG��4v8r_=�K�b�� ,�i@^uT�&HdT����ɉ	W�M-��Ct����&�vn(�]P� �T����ɚ��1;�X�P;����'1JTP�*>�(��ฮ��#��m)2#��ꄼM97}{��eL�=0�͛J�'WwBdo�3�w�un�$!m���4x�Ĭwxk��YL9�j2冹�[���4&Vt2}�A�������b�� УYi"���|����BV^��\�R��V��
n	2_AYBm���V�7��A��M��ޥj��4nKR%jx�W�����[BRv�g]훱e>�zA���wô�=�yx�Q����j�!|�캆�Y�[�"�M��׎�{�����P:�Jڼ�j�
�������������Ujdv�p&A��yjSP��]ظ$��R}uwd�mb�v]�%8�(�k8Y8kC�.���+L
�q�d�K���'z��� ���\�������5;��������@�9�Y8bWH�1��.r�:6=�(�|'Ǭ��P�-JL>�2 +����:���r{ ��t���ۺ\�C�9kÛv�4�aBHd0���`c���YPP7I�dc:m���(���v��;5�Yc�8E�SZ�)x �(�l�9]����|v@
9/ge�}ʸh���u��ua�f�"�+-n��}FA��-i�a{`�<5jL�;�k[t�(��%�����F�ͷ��������PH\�l�7�ֲ`U�xPT�HԹ٭�m�mv����X��`8����5r5�6�`�wl@���Vq���Ei��G���-�H(j�ؗ���p�����F<� �
�.�Թ��H.g�L�`�&��ڡ���6KV_�"mu�e��{u׮��ʣ'�U��Z������4	�}mR�h;d'� �-**�%�1���9t��I����}b^�����.*.>m+ҽZ���ӝY\4-��t���b&#K1���a˒�=��v/( �nT�B�b��
Ă���t�a��
ANB����*Q$��8	Q��7{�{I7������faD`3D�AF�e������"�{]���I)��3�2�(�ѓƋH&餚3��Jt�.B%��"∡4ҁ���1B"p�YP�a�@DrA%�!@�L.7xŷ�-U��� �BI?D�$��KL�����$$��c�.�$	3vIm��a�#�6�I$���_�mHˉ�L�F�-ēI�R2�Q��D(P��$�I2(�m$ےH����A$F9fOD�QG#ny"DD��"�mA�(��e�X�(Xt�'�D,��Ŋ����JT(�K���c����Zer��,c��i/V��u�3�<�d+6�P�$ԧ�r��"�ZF�\Q>Z:�JEa�"��+���h�]f�qi+c�h��b0и�q��4y��E<I������"����UĂ���R�5���Vqu,�l3]�fF�8S��KaR�X�c`�+`9&�'e�'N�l-͆Ӭ�1��$Ź�V�km��>��@���.�eb�"<ǗDk���Z�K�6�n��i.))��s왥�M��Պ��^`�����:��:TEƺ��[]��
���H�ց�ލ*M{s��)p��qͳD�=��
/:I{����ijA�,����g����K0���	�9n�������]�*<��'F�S���vL@}��������Vͺ���QtM+�t+�l�$!c^ói�ك��z��j٦�-��a�z�C�Q��B��:
U��oR9B�ue<T�r����:x����<hܠ	���A�3�W��ݥ��-@��P�"f�W/���6�Y&s��"q�Iֳ��^{�	ݕYV�ܡInx�2���ڏ�x��(�p��t֕�v��&V�<x֍z�1�[�R_]���2��UH�7��l@n���4�y�]��yp��meXr���{I�O�ȡJ>U)SF�P�ܩ�4��"&5[9�	�!��T�ۉ���)St�tv�辈��xT�lS�5��#��ܵh��m󆣼΋�e�=VeD0Y��
((�!E�H��uv��X�K-F��9!���Q��R"�.#�0"�J �F?xxxx{�ޯ}r��܉�����D�1@�eL��Z�ߏ�Sv�6��� Ѻǣ΢�W��6�f7�U��.�1
�m��Q��Ұ�i��CK�]ݞֲ�	Ҍo+QЎT2Ʃ��wh�Tl5�!�KI�y}1���S����2��E�qM�M��/�Sjʜ[�?�@�˭�mי�P�H�p�:$o>B2��I��'m�O'�C��N�f<T삲����x�Y�}�j�>h:�W������ 8^A���W����?>���3�q�����Z���ׯ1�0���=��D������K����w�_���.V���=c�$��@QU[$���jN�ީ^�fy\yuDq˸�|j�8�.{�w[{@EDI
��f�-OW� .�I�}0p�9f^G'?C�1����)+A�,cGP�Z�sWCI|Q�����ot0g{{F�؄B	����=�m`'���x�P0�`�va��l���:-����w�}�3�%Q����:���k��{�>�MԳƶ��_!>։Q�C�:�޴X8��*���z1�"���j��������p�#��h>c9W!�&��@�����%T��R�s�{�����WP�o� �)(�F=P�EU����U��F�z���+K��Z�G�upd!Uz��۟M�b�'c�))�a�]�d� ��,���T��l��>��~�!��������{�D(�v� j���#B����RZٗ}��v�-�Rm8�*}����nI�|���Dp_�v��L���,3~�L��}�*g�ӝ�o�<������F�JB�`G�>��U-�r��H���R�����P���nחu��)����4��ڙ��<�k���B�߹� �ā���?n�y���vQ��Ge���A���c�mc��W*b�z�/�E��= �H ���W� t��s��� ��!�ٹ��i]��|tD0]�� QUrgʶ�~�� ��e���{�`�J<^ߛ���Neq�]���ONr�`�DH���X�&_���O�)5e{���Ϣ.���J�vѤ�a���mz^�;�M�Q���Z���Z4�J�;F`�u�*R{�龜���>�}���������Qv�
ԱwA��@���YC��H�	yy)>���"�������f�m�Fj�}����b��j9�1���*���`��6L�b��^���w��Nn�ԺwnW�i<�]�/�;qR�KyV^j��սӉ�U̠u��N�z�8� ���g؟�!Y[�E�W_u��t�i�u�c��A6��� Cl6�����l9J��_Y��G]DKޝL�t�fL��,Y�f=�r����L���99�Y��;n�D�8��F'�A�k�k)_U��Y�<C���X�&ߗ_���Mzt`�ia�Y�W@l}�%�$'�@N�o�G���{��T��\��wQ1z��[����x��+P��L~�Ռj�}D4��QC_˖Q���C�ݸ�w�Yo��c��#0��-3���fH{������]h	�^��*��KHŘL��+>?u:���p�������R���Tzxl�� ���J� E�bK>��Q�W]N����`J��,�t�,N|ū�b���I�Ur���&��Jp�]�����Y�}2�dX*Z=
\��vX�iX ���^�?y�� ��N_I֢�lz�i�Ơ�h��h��������V)v��{�7�U:�o�n1�ڌ�+��E���E��A7T
"a����2(���" ��޷�s��5�x�B����|��C�+�	��*���S&'�HP,Eͭ^Z����Y����o��& �E�W�+R�v)����I�Q�!�'8� Y�a�oem�>걚F�@q�	�<��@�f��F
�+u_˦fɵD4*�9Gs\v�L�r�>�E�Z�zȉ��
�'M-�W�4���ē�'-�M���%r�1xVo0þ]��9��(�w��@�ێѶ�J�0��_%�M̫q�R��n����r�:AxP�zU�X�g،%[�~?p���)���d�(0����[�;J�A�P�G��@�*�b�/��dՅe�������뭲�KQ1m#U+�2W@�!F�L�;B�����Q�����tz�B	�j���:f#x���n�2�
��A�3�^jSwq������k�®�v�Je�����΁�t�kx�^[�h�2Ϸg�nާ�}����D�hQ����� �V�6/���%>r�tm�4H�AbŘ`��)X�X0"��7�{=�S�Ž�^;l���C��{;�i�+�4'�$�s��^�#U�A�]�|���2�>m�_P{�4�Äp�}Us��|\�:/�6��w�Z#F����e��.M�g�|ښ������S�a�C}�y�Ì�Bd�a����;�՘��ա6��>
��RD�p�DQ%�F/5�B���e�����x��0ΪuΪW@u��F�`���Ή__nñn�?q�U5KޡkUa�^��1��&J�Ր�Lֵ��P�M��-�]ڕqlv��&ҡݎ��(�=�m��A�J�����G�T"��s����-�e��A?c�9��%����f�h#���V�h��o΅�*�����'�'��( 4x ke���^���W��&�5� �@~0�(d����� $���x��!�	z���/��a���N��>Y��7b���
{}x��3"����jϰ�zF�2��h�7�W���<~#�CZ�kW{�-�mne�O��u�h��I��[� 8c��kV�l5�?F��W0 |~�m��>�Р2��?8EW�Q+W����<5*����E�����oFA�uT���5 yո�j�����/R������N� D���_mA���D�`�,�h���W���}�?Do�F#�IL���P?�>"�����F|��х�u�q�B���j&l$ ��Z�C4�V0<d0��"��N�,�q��CH��|��?K��OR�	��0�=�S�߷�,?�$7��J^2�~�,�#�:�$m�&|�Y��G�@�!�@�Hu;~���I��Z���4�Awre����]!�O�m<�q�b�X�@�|]D��A��5��1�){��Z-| ��7vx����}z����Z�qw����U§��B8ԑQM5.5x>;�4{v�e&�ݬI�Ò]hU[g	����A���@Q�b�}��I��b��iu�u��B_{c�y_�d��6߫�亞��C�����c� e
f]�R�e��Q�׮���Hsڗ�w����0mL׺���}L�t��3v�~fo�9F&�˧��vn�v��9	֘��F�#�����9��'q��'V��}3��y����#��r�6(a�4���tCpl��!O�l(23��߫���@U�������#$`�b�)�����E���7��q�{���rt׼L���8�P�Ac$�w��{�q��V�B��[�k²�$ܝ7u��V�=ٱ�]�W/�U�A�(D�%�SgW5����ϱ2׈�ڌc���4�雏��B/j%I�Ij͈��I��kG��C���֊�N�([�F��ㆁ��;!}��=����|>�)h��H��}�g�]/zQyIą�,�K�7�/3S�/W����S�
�!�f�(-�1���2�p�:�D��Q}�����N�,]��fte�a^�<Չ:_�*q�݊�&\�q�߻��}��CQ��1rN&���(��d�U�&��f��r�{7��(���G�g,J�s��b8��)c2)�Us=�d��s�����-��~\t�^�Q߮���Ї���s�)˭�
#I+��ݲ��9�����=�$n�l���3�Ho/Q����"��=�wڣd�K�ɪ}��<dñ�.��!B3p8!A����֙�P�#?D��a����;wvw^D��J1�Rc#B���L�
�g(���{��o_^Qʎϴ�1sB@� x=��⍚p'�E�+�c�OPUR�^��S�=|����戞s��Pq���>U�&wh��i��� ~�����*��ָ��C�r�M!eB�3�E��<�� O[��߿P��ˊm[�l��((N�IOL��h�;5��^5pS[�48xxW���	�N�8\~�g���G]Ja���'2���w�@���;�l���{tu<��ݧf��421�J���]Z�U1-�X*&�kzC-��PT�o5���<����׼k���;���)TQyK�(EGR:��a��-<��R�b������MD��֡˵��\��},>��n�j|��ų`&���� �7�� 	��$D�"�(�����*���b�Zε��K�J8�A�i��A;��<c>Cmsۄ�D�u~�xѓ�@n�B���:_֋WE��%,$��S�8�k,к��w�>-�*p*��BDb_�c��lRk�>��kw�_,q�y`p���tlM�#+��G�>�$��G[ü3=k�M�;]�X��-X�;J����W)�Tn����*�ԁPT@U��we��Y�",�DX1�!�`�=iH��� �y�u�W����9�kN��A􆯚��8���+�v�/�5�^��xG]=� �lh>K%谡V��������k^����e�x{�8���|��z��4Gcc0܌	�X����m�l�|���9��V8w�\�1^�Z��.�B|!D�r�0��i؛���-2l#f��������ňE���#��*y��ۊ��ۼVI2�e)4���"���MP��{x�"ynە�aX�|Ͻ�M� i[wJ0�q	��hB\mH� �F����~nuF����5Wb9���-�<=�䔶�Tef;�ݨ����W���ȏ��҅�,q*�Q*�f�l���3M�MLK[;�Un7,X:�Qt��SkuquԕJ"���A�f$����#)�WK��i�ʠ�$��0�q����j���$������VQv'6Y�t�?�r�00s���ud�>��M�F��
�ѠK��MQ�� �D�"x$HB�OV�^ZG�2�%��0ɼ�4���6~B!�6��ˏ�#����[iL�8�����"o�Ǆc�(���#��>_�ھ�%��|N�C�S�VA\�$X�o����ouX����|����w7<�;j:�ѭ}�Pg�i<��ؑ�s�x�v͆��]���Ql�ѫ��}���o"�&��ؼh�E`i��Zs�r�">ް)b���I�7�Y�,�%�� �BԈ��Z��E0+�e
Ӗ<[͙��K�~��V���aK�x�v��l��,.�Z��&�A�}���-^�ڨ�E
R�$�Yt�@���p�r����ҳ]�40��~{�ݔv7$���6��9Ɲ=AۓڌZ*�2�NQz���O&vvOS�=�ħ������%y��G��4�2`@�!�׫�53�{׻�V,�ݭ��3T��>���;wa2���c{3�=6qè��ъR��M�&ݾꥷ'�&��p�3ou�r_9]��[Sg�#�8�c�Gjg�a�U@�GlX1��#,�ٽVf�o&�7k�������pg|5j���l�>�����]��E���bϱ<Oo�3�uy�Ac�W���QZ�M�{�wP"}`�c��^��\X#0Qcd��U)Tg3P�D�HV�
�΍�76���]$i�P��4?vV���&�H>�r;���{z�|sǇ��
�����j���lT&�4o��#���/7 FBo����?����*��j5A�b2�Α3�*@uG�F��0�XᄮBr�d}|^�Ѧ_%Gl}��6}�^�aGVۥ*���W�@pi������#< �3��c�|�Sƚ'5��=�s�8���[Aᩌ������.��)�C��T��@Xw�}�VH�=x�{݊1|v�"Ȉ *�� _�7�(���B�T�ŏZQQ?h�=�u���'�m��x�ဍ���#(�5t�Xf��b�%�L����f>��[��G��d���a����M,�6�n� �H8D���CV
.^h�"�v��X�'v�Z��c�n���7|�N��D�E,��G+��\��eٕL��H�k�T�
��{������]��<��<E3���Ul����i���(ο���}��m&6��Rw�b�p�H*҅��c@V�qNq�
�e�9vK�U"c�|GT$cL�>�]��M	<LU�t��Q�(;5�Y�3cz!����J�oӻa�of�nÙ+1+�j��V��<3��,];sȂ/zCz0�0�-�ZZ������A�Πo�8!gr��A�mkV�>�oN[�lֽ�.� �z��ŭ�,WSw�����S��3���ߺ�=���hj���4>��K��VT��U�]j���*cdɷJ����m�l#,U��������@����V��Y��[����X��(��}��Zؼ귕7,��I��5���f=��\GJ�P��rB�V�هu]�ĄG9f��Ȃو��
"Ҥٮvm8�`Ž�%]p��.�ܙ�Xn����՚J��o=��0&����CL�$��"ڋ\�k ��W �vUZ"�(�h*�h-����c�N���)
=�!1P3Ұ�.��P���̏mm7��~$�b6�ы?.�TF�]��ɔ�����3N!O��^oC�wk�:/ӷ�p��H+.^�����V|4T�c�":Ki"v���Z\�H.�Y{�(,8��	�u	�.�.@��o�u�[�[�����;A�}�����{ձ�Rl����/ep��.�9��zi�~��_l��4���f���'Ն�<[�s��GQs�ܝ���3(��4-�@Jͷr �\�y]�G�6PSּI���եNE�IeٸK����-�v`7ȋ����
TqthV\k%f�˺pS�:�{�iC�i�U����c��򄮕:��[��Kqv�yM��������JԚ�m�u���%5�TPP<A YnT�cM`˖�+=��G /Lɩ,�����1e2����G*�˃l���[6�N���v����K�2.Ԅy�Q'(���E�ki�r�����)��Sm�N�{[��k��s}lXyoxu	J��[��gr�\*~j�����W�z3li�Zx뗥W\yqVv'˩�m�b��I����#n������tӺ|[��C��G9��ݰƷʷ�S�=+&�}�Aq�0���Շ�-{g1.x��í��C����~��~�����O!L�'{����+� *����j�ˢ[�D� b��%v�a6�0ǎ{g�aa�h����n�ea�_5T��9!�S��3	�
I�i�����N=�H��)�o4��3���['[H��ؼ*Av���b�Hy�m&��۔-P�q��
m:���Rs�Kb��y�AL�RM}G�a�S�N���{�����a_TsF5������
w�@[�al>aI��i�-��\�}���L��Ľ���[`S���Jp�:`S�a�縓H['�� �!�4�5(���S��UHq>B���a��I��TX��T�0R"�]���0Ea:������׎2e��f�����)2�al�Z`m���:Hq=����-��2S#�
C�e����ؠYhS�F�n��RIL�g�r�L)RX�Z|�![�{��h���T���� ��,Q�(�wI'U����~@�U���}u��`S�8�Y����]v�(i&*�S<��öM!he%02�u�4�z�,UE'L˖i�r�sah):��T���>����l�c+�ם��i-:�H|���4�#o�R[L���a�0�z����X�(G�4���W}�8��N0�o�I�Y�'۩��u%�6����4S)�q6�:o�s�����ĦN�O���h2�AAALr���3ڐ��P�e�2�HW��fM+e!��>m�S&R�8�OXn��-<��ٔ�jC�2�/tMn��(���~�1~�����0����#��g� ����N2i������^*� ����PQN( ���#�	WHi��)5ʆ�Z)��|�UT��4�Ň�(r�o:tY��/%ED9$@ @D ���%��[>�B޴�(R|�������E�`i)��G�N��i!T���[II��ҙ���s���f�
y&����2��z����{����!�8��5�r�0��SHn�)�������S��g���0���L�:ڲ�C5wI:�éH.���MVlHf��&`D�h�@�S:�Ld'ćXB|�2 ,6ݘ���c�U�݁L���j���e:s����)�i�U!����˓����U`���cF��oV��3pri��\�\naίUX�v�e�S ��L�I:���B���a2�8�a�~�>��0��N�?bM	ۻ�y8�(O�R��<�O$�g.�%�u8��3��-��!=�~�~���[�X
d��d��	WP�O�Sl�I8��%8I�T�ɆW����N��AE�$�8��P,1�X� �c�`�
���g�Tyj����͝(m����s�rͨ���(��i�U0�o�"$A�TY#3VaH}	-%�����-<���S6�&*�l���yu4�Hq�
���T�2�UG�2a-��(,Y�i'}Ai)2�@����w}��x���� |�Va���q-�S�&=A��	RU��A�a���h&�a>`��R�E ��&��⪉�RAf��C>u�B��4�$���o:��k��^���i%"�"��y��̟6��� �>��ϙ1!5F�v�i��P��m��+�Ru')����� �w��J��`Y|�-�RO���xz�z׫Y��-3�Q0��
��β]d��qZ��0��u�U�@a3�h.ꈡ>d��Nm�͵�Y*u%'S�œ�d�Arϙ�a���C@u
=�.����=�6�!L.��He�B���o�6��>��C)���!�
M'���G��2�E���<�Cɖe�
G�%��q�E���8g�Ǔr�,��-�w���f��k��|Z@���S}�i0���;ڒް)�Ï	
|���B��p)�!I����Jd0�}�`/�7�i�-&�Ro����D���W��7��;�$���&ٯQ�iH
N���E ,���KaI)��}�#�4g�!hu��!IL
w���ɖv�W>Lu��$�GU
H)���~Ű2ȴ��ѭe~Ͼ�{�C�u�*$Öw�@́��8�і	�쿓I-�)��l^!Q0�_�d�a�C"d���e����1��X�Y��8�\�<�� ��Py�5�-%}S�YX�-���K����f�ӿ�׺���[�tq:�T�8�q����]�q�]6��L	��q�I���tIUº����n�qG��Q���3ͫ[[ˤ&����a%�}�Ю4��:0>�D�p[�/3*���S؝�2D�Ԏ3�(�M�vF�6��ұ0����$�4�^>�چ$8�f�A��*��j�4��B7��QdU	Q�E�/z�Aa�J��{ y�C-4����.��o���)�|�l��}X`ZR4�'n��R��r̵TS"ʹ�I�-�I��$:Ӫ����������"���"�H�/�PcDUz�5�k���(m%'a9�2�a��W>�fXU��ʩ>��P�:�C�0����D�EV��
ШSH*F#$��T�bq8AKB���_k��y�Z��q�B�M}PӔ���GTC������i�KO�������{��a��<�?0׫̓5RRa��1��C	>�R&P��}d��œX�\ a-&ٴ��<.��u�0\�O�A��>o��HGO�E�ΓL���>����&���L��)W}���1z�d�e-�!��y
b�3�@e�ʦy�Te�~�u9�60�E��q`bI*�QKL�Kf�ZO��|���u���g޾tI2��QT6��m�����@���	l�f����٢[�Ke����E�
m������5xv`��m�a�@�ա��UZ'c���<�)���õJ˵�O�8�����R?0�L3�))<����,)"���6�l#����i�ꈡ}�[>Ich)ԚN a-�~�q���:�p�x�дD�e*Om�y �E
��ɇ���=ʚH(M���u�]�`����;�4�;�z�L�V�a��n�m�Ka_}cʓ���l꣉)�'����ϳ�v�
a�T4ᒾj[aH5P�g�\����|Զ/�;�8aH(�r�Cw��m%'�R[!��e��P�ul��� m	�P��i+�Mzϸz+
�DU/PU�o�qn�1����I�e��
g��y�HL	�Qi�f[�AI�y-+�>a�.�K`������L��m-�I䴊e��KUHH|������C)nP>NbQ{�w;��ux��
e2���j�������b��S�[>B���l��Ĵ�a���/�5w�������I)7��m���n��qv�a�іE��{��@y:���KCi}��������u�A�@�U����(��U懤�Oo��NS*�%IgD*���+�����;�(^���F�m+
������/�OP��XE�=�H-v�_�Vy�͠�,�IMn��d̕��ZO%��
z�I�ZL3���a))�Bd`(��B��Y�d�$�
L�C�I�ZAC�B,� �P��UE?U*>��b��X����{�s�s/���8�ٵK�A��L��~�wɩ��PE���6��,+��L$��8�>Cޠ��(>z�д���ILq�Y�e����]0�תةц�t�=��_g��+�H,
��Ä�n�Xa-�IlQ�*q�l���A�,0�wRٔ:������n�e�i�!�� �a�:��X��ƈz�u��g��l����_/9�yﻭ_���Sf;��h�B�>���(�M�g2�Y6���)0�T��u;�Y4�
a��*a����A�	>f��4�
N}V�B�q% �u)6��{5����:�y�0�+֡��- ����(i%']�Z�PP��s�5�8��I8�I0��O���va���é-�fࡄ�2�|�̡���L�S�
t��g��]�u�u�ߤ�9�1��C��>i�Cl!��e ���'P�<�1!]�l�p�̞!����RcTb������e!l)����dJ|�8�Il2��G�V�u�"�d*gg���+ӂ��ۺ)�q��Z�2�I�KKI�)d��x����[ ���iT!�[&j�h��Ag=@_���i)'RC���n�!��-$#�1��O�!�E��O��J�F1g�S<�a��3�Ri)=�1�p��D�����6�F �c/c��ȲFL�dMY��� 'i/��L�-쪥w�����MI���d�0�/�-6A�G�1�]��bj�|^DG���M�m������I�!&�>����/f��Y,�vO��V��@�� ZD�1-��▐[�1#U���E�T\�H�Ѭ=��[���a�z4Jp#ĘHZ9B�<�s��*��jZ;��v��U��O)��/:��|*�	b�O�L4[�9L��k�K�gt������ﺨ��>��)����zK�;�4i�}�X�h��W��a7cN��T�O������!�f�����X�Z_���H'L>0벼�@jI%ݷ�{�����8��æ�=B�>��}4ԯ\�t$�W�~M�_���hf�9��}�v�����у��"��_ 7�����V"��������M���M��8\��H��U�F��������ؠ�]+9 ���<���>���U^ul�"�DEW>-(�d�E�Z�9��שUzq�F�ML`XXp J2�84�O�f�"z��Ԛ��l~���b�����Wn׽ kU0��$q�JW��10|s�lx1�d@�q�����|o8ޘ���}�l��3@��}+��L�t�˓\��h�~L�\l�a�1�2|������5_���ڶ=��-F��X~M�2��7?|;����^�yކ��T�!��T�` :���#�0H���Ԁf�v�żo����{SF����"�ꔩ"*8C-��DEt�)A�O���QSM�v�d�
%/Q`�M��k�+uݪ�����n�wQ�X���`�	dC�G���)0�N�F�`�mT�T,:�ٕYAO�vF(�G�YR�[�7uK��O�l��w!���$@��/E���0,�2���+ϋ"*<ʵ��/��o�:ܻ�J&%�mex� }�ю��)3�8<<ˈ��>S�o�UB��$	��L�hs�H���3źT��ln6D���|؍��fu8J���)�:��Xa����	[Q�0�����>�|"���680ǼL\X�Ƹm{�Ej�F�YP�����t��~糰���U}T����\}E1f���P�,EV���c|���[Q{�1G���R$|��(@��&+y���t,���Q~ -sϫF��Ro5,��m��[��"Qv��*�O���~�V�n}_�_��B=�w�>��G�MQ��id}Ȑ������J:ˍeɛs������f��O�m�C��֘eo������*�S��u�Ec���$�B$;�߯�1T����ȬAy�6a��� վ��Y�#�zf/�2�>n��c,�����
1��<�pC�ʉ[��� �с�>>�Fw����On|��Y��7@q��G�6����EG19p�Yj&da�	�x�����<�^BX��i������i�"�h��#1S��
@�:�֞s���Y�Em�P�~��$ð993�ڴ�h�$��l^:vΒ㐂E�]k�Q>�3���F�1tv�j�P$��dj(�d���`��	$�������$n �U��R����`�|HO�����R�0���.��z}�9\a�3�쏾����U@F3w��p�v �� �U�p*�T:�����W�/LF��͝�1a����������Q�D�[/	Zz�����>��N����v����h�`�E��g��&@�ռ���S��u��u��_����ãu����^;p�x���|�mP��$OٹB�_��ħ��|y�{:�{&N{�10�5v�ru�59�b�$kԐ��ԚG���������w����+z`cwf �X�+��jzFFx�.F����G~>����������-ēPs)���X�~X+��^p`���[�=�u+�}{u�H���ATX��{W�z¢��W�>�՘o��2�O�2�*��0�E�&b�!���`�W~��P����չ�ks��+����C�*	~�1��	:�ki�۟���Lh��׆�	�Upk��FV�
qGFDvJ@��L�6"G��I3�'�R�-ӊɆa>�a_Vj�����9`I�M4�(��o��bR=�c�.͙�c���D��[��r�l�.3����rME�%K�Mc��j>��,�����9���� �N�5��TT�dڻ~_�����<�([=��R}�"jC-�N�η??��(D��	�'y{��d�X-�q�En�D�Z|!2겨H`Q񯏫�}˜s^�cZ��|db,DF,U�UD`UJ*TH�T !H�JJ"���y�9o���w��汶s�"Dل%y��L(C�=eK��*�1h����1����_k{�U��_U���_�sC����L�LŤV�О��0��<��^������F3:z}G興�ex�[Q�'�'��e�Y� =��ׯ{ܬ����~�#����}y^�\m7M6�E�Xc|�/��}u�����\w~�+ҖRR���O���	]��iv��>��=��OW��}�k�Ʊ[����X�X�B#X##�}�7����'��o��cv������|�5H�A�D,��X�>��w��`�7'��w���ݛ����^�mL!�$ݍ�sT��p,4��y��2ֽ=?{J�w��Qꍬ���~z,x �>w�����@�����g�DæC���_A���x�?C�\�����1�z,�>dB8�-S�Uڳx��Thi�׻1�Y+�;}�.l)K�������\��5��i:PEM��E)���9���4w�JU�*יs��ɼ}��@��N�cC�zvH�}�]�E�'��n(�"u�l���4ȸ�y�m��
�4Y�|�yqu\�1�K��l�0/��q}�w^I��o���B(x<R�µLp�;u�I??j�]�_1]l�����P������KY2�ax��[9ǃ�Z�R$:� 7M����ֱ�:�d�D�PhA�̲!���z����L���~����<vpG0@�����&J��}�!�+�5	H�V�����~���n~���?�^ѷ���u��������οb��\�2�זӌ8������/��W����zr�anm�����	'��h��ƪT�"�JJC7�S֍%H#c���c���צ5�ᅛ�j
��@��uL�8R�@��$��%�X�@t��Ó���o�r������>�k��o����g�=>:�#>26R&�O8�ݽ#"�N�fy��p~�:N�-���v�ٽj���޾3���>B�m�3T�?h����s���%��N�*rgc��O��>Di����un-�׻�],Nd(�X���t3�A�P��+0�&��1�@�HKÎۓ:FϡՓ�e��$��S�p ��'�����F+��<g���};�f���RCb��Q��}���qI\���}̟I!�H�FA�%r�TyϾ��>s}M}B��>�_5�M�M���ѫ)��'(זEP��'n���7
�U����r�����z\�[�C@wo�>�ə�9oC�i�5x��",WJ�i�Xh�EO�dA�*��qos�5�xy�_v�2%��S���~��Ȁ3��3��s>��~�{���DPD�)��{++p���y���6����p�<x|��7�������w^��z�3=�{Ǭ���V
#)��QUH��-�Jř��x־����Q�z��^a���R@`m��G�^�q�篗G_W���Z��s�����5��=j��FE��)��"�z��XR��͂��>��R��$<"�ĕ<���77{�X�F]-��Rr�S^��:6L(��`��r��uB�gqM�/w��g�Ǚx���� �����?%�4~e`ʐ4�-���ޣ��ފ�w�|1nTk�Z�����n6|�a�@�ңR���ss���A�ܓ;:cC3Q]�7H�Hɚ����V=ʛp�U�0���Z�����F��m�M2(9z�'�,�2���=�d6/{Prܶ��,K��0+�eh�Pa�j3�O���d����ٞvVN߲��ͽ��t�f/s���(
0p��&��`����`�<��@�E�/��~�^x�e�y�r�H�#`�:{����6�b7��o ˵CF�J��*v�4��@��
�m��6
a�.��RZc ��n
�z�Wv.�����Y�Z�,jsOL�J����뵊��If�ݷrs���[/�4o�Վ�Ѕ��D�w��aS
ܮ{��+[{��*dsil,Jr�e6{X+]JT�s;�#�s��xr���J�U�YĄguhI+�ud��"�ox��Y�:n���Yr�DFNs�=�mɳOuӀ��Q!{F�ΝԠ�+���vt[�b�L_,�eB�J� ��HxgSx��0j�
��te�t�n�.��]��i9�3v�HJ�J�VX�%Z���x�f��F�6��eb�vV�\z��]��/��h�~�΋����O�:P��_8o@D{˱B�4h��
�/��]��sw�3� �u�e! �6��2���]O ��=�l7e���N�vR�U��KyV�d��ˮ��$��m&��F��ƣD��H�R(�.BY-�����'ɒ�nEh�$�EJI�H�q�	,��i �J9$�(E�
)� ��$m�����H8��(�l)�[0�I3���^Ub+��"�[C�b�%��fU��M	G�5�����j��C�*k�SG�1Y�fX藬P�pۡ� �F���J�t�>昧��꫅��T��=)�Bf)Ҁ��J�³'_>��L5�֢�ժn���!\�2*��ӛ$�N����Pf����[s"ۈZ|Lͺ��h՝\,B�,#歊�ʞ���ӓ;�ѲE��3�
�mtd\7�Tx��-���ȋN�8m�f�C:���e	)ª�u�F�B�E ��X��F�T�Q�5iݗ�"Q��6�V�ꜷV�2�����wH]��ʹ�*���7~,[��o2�k�t��9��ū���(S'U������tPV��uj�1J8P��Ǧ�WV�6;���2Ⓕ��q�1'WGk����.��Q�'*��;%���vKw�ZQŪ���a*N���0��{4K�"��s�]t�����簅��� �y:+��W�.��d��9��\v�%�X:�ps>��Az� �*�������^��\�J!kP�v��iEuY�K���'i쨩�fՋa���0�5Ą�^[;fY�wl4�RҊ)�b_U�b9y�s���0�:<����>�g��ThuSr}ìg(t�G1heC�<�s�0���/N�Kچ�M6H�j��ʭ�r���5����֪cU�S�a��<�/T�\t��C��
#ˍr�1�T��������ZH��\�i�O%��%;���i�GYCRt4������g.�>M�u�%��N�-3A�U	m�Z]"(+-7P]�iT�\(w\�˰��$!�"rH��I%��P�I
1�Z03<��I!mD�
D��	�'�J�F	���}2��m	�I�
��.=��y��էy\�ܜ�Z;y*_��U$��$Q�B(t� 6m#�.ན0��We��Jɤ�ك�,a;9�׬:ۮ�fz� ��I�>~njM"PGE��f�19#��J��B8k���0�fڄo+eFg1�lq#�|��Xa	v�������s��E/���`�b�>�31r��;�Q0���5��s�G�g�IT��y��^�;�q#��T����<�1��~0��p#���pO�\9�sW��;�p����*$�� x���>�mJ���[ՙ�y�>�W���^�v��ޙ~0V���Z��c����W�.Ix���|����I�B��ܿn����3��	���'}�.�}W��o����8�yUԯv��CR10���"�ʣ �a�#�_��dB~��G�Uoӱ P�:���|?(��ù���"�u�ã���NQ[b13��B6Ϙ�m��c�Ex�;��^�������O>����uM!*/�%�j�E��A*�z�< !��}��
��ַ��6�`�=䏨>١vb�`~>�A��Q���i��?���mW�s�I�qgʥ��b�һy�^�=�Z��QB�"���1"��,j��R��6�S	J��1X���͚����QVy����	$�9�EEE�F**�������AW���9`�ݧ��<���7:Qz�:�MTaNSӝ6+Z'��N�}����
NZ�ua�Ơ�R���b">Q�U}��R���R���l����g��>`杶������1��^�*x��@�E�$1�`;�G:"yCDPo�y{�=[p�i��Gw?ѽj�/���*�OV��3`s�)lt�� ���3��!��狲�^�?v������O͏�6^� Bb�j�!�Na�Qg'�$<B�� r?>0w�o��D�G��Yi�lǣ��~T�[�Lb� �$D�EDb�1UQ��=P�H1b@�� � ��~�^SA`��[���-�J:4L1I��j����E(�hM)�ҙ��:���$���BS�L\�� �_\�����+�U�ų-$F�tLϛ�qΈ�!U8`i��}�������W��E�>f��ҳsV��mxL�	��F�4R<_Wz��<):������w^���z��e�~����S��ƀ�Ŏ(�"��:��a:��t�'~��S�S�nf.�N��}�3���*H|1`�Bj�@�����5㕆߷���U�>��;��h
��Q�m��~�s�W.��c����#1{Г�z���뜰'7E�����Ƃ�2�p�L�{��8���!yr>݃`)1j.nP�D�f��x�h���خ�z�����]��P>0 �Pu-�[��z4h����V�|�۹ţ� �oؠW�9�*����#���o=Ҽ��w����/i��׊�N���!��o�>�WY}X2�{�}��Q�S8�ޕ�71��_�#��ٔbQ�_ |�)>N�,�k�����	$����q��Fzȏm�?T]�d����n�d�_Kq�a���GpV
�Q�*# �2�� E�\��Ƥ�F���IMaB��#:�]����1�l�{z�DwP�Y �Ю0;ّ0��*��b4Bg=��"[�~�������K'S��0r*�=(B�?o�ps󏾏�=��=�0w.�H���ӛ.r��7��Ba�{�tT%�f�Ȟ�?/eō���;@·0�M�����έpH�mza "��\�0����٩A �_r'|<<�#�ʮ�<K��?g����� Ei���4|���fd�����#��㾽}w�"�y�{^<�*Ï�%p!�p���8}d=�Xά^YW��<�@'�׋��/{������*{����Uw{jR�>�}p��<����sw
E�����W=׀v�dm�ǹ_̻�]##�سG=l}X�N�PH� �=���:������b6���L�����'��u��o�}_M>�+�9������Hb��s��=��uDUW��3��*U�5R
NP�,�^���p�#����9�`3e�6zxA�7���e��g|����}��ɳl�>ǏQ�y[7U�>�����U5�$��s�s�5�V�F_;�{�
,F7@P���DH�#�?k>���_s��_*_MU����k����K�Q�򑦐0k'%�<�}�Y�^���-��"�̋���߷�dLY��2~c�diȅ~�G�}_�I����}�"ǽR�\�d}�,|[Y��◮���
��q�+�0*4���wb�i^R�e"���>�NWH�!�z�woT ��(/p��5���/}7�����;�4*�!(Ȍ%bHJ�k���d�ef>�����<���������u���D��o�c�!xȟnV�3(�|����K&q:��\:�m8�6�Ah)��E�ZH���Qɟ;)
���g�� ���CP5��I��Q(�IO�8Q�lB��G�
�����U�N�4=ۤn�TǹνOd�
���!����f�3�<$����₴����

��HM��PnRk�W,�m:��ҭ�ꛅ��R!��$�&�lF�f,�D��J6�J!���sG���Aь8�l�!�~����sS3�� g�]���Q7��}�.	Q�:�x�����?�Q뉬�EM����5�C�/��˼'�ԏ�G6`!70�}���y�˳}�8ȄT�s�pX�	T�u-�Ǫ�f�R�mOՊ�Q�{�!�*�����T)�2 0POT��S�r��	|�`a}�%��d�ƌ6F�nAW3�g�\�|��Q�nXA�+�1��F��V��
����lE�����������\��U�V�����j�����ٟ>�w���!����1���{�)�zP�����6Ϝj�r��f�ǧ_��!ݖ�`�]3Ä_E�v6���}qʸ8#ޙB�kN���f
[��s��<�_�`8���09�8,p#Y^��A$�o�d&�Q�$�Y����~G�=^W+��Z�U#
Q=�YH���MJ��0�SO���Ν �?n�w��s���P�fu�c��=���Xڭ�1��v G�#5��Y5��$qcGو��x��/v@�G7��� �
3��e4Q�r�2���)&rԶ)��fsǽ��v�w�x�����<Cʊ�u��r�L���.x�3TCK\���7ϣ!px"��>+�"7���v6�S����6�j�f�,/޹q��`U2DF����W���$N�͙PBlN�u#|ť渂>6X�' Rh�`
�CCW|;��b����p��O��5��m�D�/�R*�j�U�"Y�f�@�����������
�4_ﺇ�c��D5쏾�h�+�Õ�T�#��s��BW/�v���D%��ʽw��1=���)~s&=�p�k���Z��޴��F�1iL�7#���{��)�#kU|��~�9"��H��(g��������y�yt�Jc��5��u���,]kl�ΐ_�Z�p?ք#+�;?&�<���}���!F��;��oq�����/�c'�8��	�Β��S���*C����#e��48fԿK�u/ M������=�� a'����|�`�3Z����?1>+I�u�X�.c����!����8�<j���}X�y2ҁ?.8��ǭG�0��>��E�̢)�j��=&}����	�s��ي#��d��!��c f8@(y�?t��I-���L8��!���0Ix�>H[�G=���p�f��h��#�c�⯉|�uڧ�2���|���]u���S�tgI��՗+	�.ՇSl+�.t�Q��
�W���K�=|Zh�i�m5.����I}~�aT���@�Xl����3B��k��裾��1K<����<��u��Us7�{����(�,�WfY��~�ۥ � �c"�Yv��+"����k�c��x]S?p����(lL�Y��f"�=��"��R����>���}W�1�c���ӣ;Uv��U�D�;���ra�]<��$3����ڕ���J�I�G7"�J�W�� <E��ߧ��c?,"J;4��Z��Q`��ܴ=�hňg��Uٗ�X�jS�@�o��e9=��g*���� ����20�:�c�2�"K���-�;�xDP�����!#�Il@V0(���\J��.��l�5�i)�{&}^���\� �,ld��Dt���o�0�6���F�=�i��V�#�??K&bmd��)�#ǌ�jbǭux���o.4�u���>��Ad���OF&c[���M�;~�nʻ�LeTx:��`ĄT���1���d��t��)�B*��ā,�����Rq�g٠����0q�D���:�4>u;�S7���W{�@��@Q��ʵR�X����n:��:��/9���Y��(�=Ғ�;Vا�i�b�G�i��IO�R���c���^��8b}G�L�=Q�>���޾���%EE�"�QPTEUUQX*�b��T�rY�F(� ���{<���v��菑��Y��p�1�XJ���DԱ(Ei�8 �c{fY��e���0� &�T�Yl�ː"�65*��،��(��������x=}WU���s�I�H�<1��u%J9"=�T�g����}�`}[��i�1��G��v���apz0`��(DyK��VÑ����Ʋ�����Ʉ�Y�(�н�z���$|��Eߔ��؊�<J����ە�`~(�&K�a���0,�I�=��!�ӄb��Y"*��"�A�/ݚqEu���C����C7�߳ޭ�����P���Pц�QUC�Nʯ��j� �FET����:�����ۛ�z����"����bY�/	��!Ʌ�T�M���S��q�Ng�kݯ�}^��x�?�<�q���jL��p�X�;��~��r}y{���T�w�μ�� �՟��CS__?Hy���<�1&h�ڡ�2��,MVl�F
|��U��CTQiŕ�s;��u�G��������/^UkN���b��e��bN�e6�,�4�	�b�S﵋t2P�+Tg���K!�[�#��b&NQ�bYhb�GXZ8.���x�3O݊0
�~}u�N0��9@��MS;�ĕ����*����9ְg(�����ƭ��Q�I�9	��E��<�
>t��N$1�5(�4@����+ݕ�)��g���h�������eH����'QC�qB�lF\��c��P��:�F9�]&6�b�P����7U6��.����3�|���7flx���~B�y�GB�.�I����N�Q������U��__��|�F�>}o����\˞:��`M����d�ђ����ѽ��j������a���]pL�v��э��J�k�ۻ�=��DT �NRδȤr����7O��v��|��#F2g�P��-�~�:��!�n�!�����]X������q�|4?��@�;"�Y���o.�|.6h�{Z����~~[���X��<��h���t�R=D4`���Dp��驺'�IS�����4�ء����UU|�/��A&��~�K%���J��8xO��״~B�i���!���}3�t�u��:�h}t�y�H�{E?^�i��2=_BG�f��ز��C�M�W�JCSL���&�XE
���������*���u�g��iQAA�Bm��?W�G� ��ð���g>7��̛؝;���ކb1��il��K���VJ�r!��˾w��u觴ަf��{�9	#(��C��eL�<>#��D���3����ʄp���w��a�v;�C.8@�4�s�V)�sC��ؗM�Q#�c}�2�ٙިN>��/"�dH����>dY�a֙����f;(�vH��,�Z�W��bP�Q`�1�*��.s��1q��<�yR�
�`�^s��Ҹ��%�c�㵣��W�*i�7�0�{�W��?U���@*0��E�U=�a@ �M�ⴐ��^��V<�����+� �{�*����nt�b4D�"��]_����m���lIﮡ��QD�M�r�Vk�f�|+�Ic���F���w�}�}���πWvW�`Je���n���>�b8����z\�;nF������|��.�&��N������z�Z#׍o��9o�M�{��������w؏X�F ��ș��*�"��U
Tx�����ww��b� ^a'��_��Ug�__~�M�����p��������?8GP�ą�\w�C�+z	�n��c�2��&�/�
?*DW�e�=��䐷�dȍ��N���f�~��G_]wq���ݕ����D!yu��ChckCOH�?P�K(b�,(g~b�B��6r��~b��W������$�*tUvL�:ج�.���t��*e���[���ݥڧў�QA���7.�3���N++ �ȶ��-�8����1X*�x�	z��8%�}pH��*�]�qB��-#d/y�Vj�:�Ķ�=-�M�[$��rU�w� (�
�����)m�R�R\��.��eb
3�а})�*$�c�X���n�z�c�wS�Wm���e'�(V��a޲��$�����Zut�=OBph��+�O��uȮ�{ =mܚ��C����u��͆ێ���v�5ڭ��R�����Y�O��2��]�G���6��}A�E��Ͱ�obU�A:ܔ��v�4-h����=��sY�PN*n2�(�Gs�J�s���T�I�W�-��e�- �c���u�o3�6*mkuҔ� t�^�BK�],��0I��Lqof���$�N�)�W0Yౌ���6;ER��Q/91@�Y��pb���s�ț�k*>��Nb��V�Y��%��^Xʒ"�.�*U�6s�����0�]�hVX�H�SB�E#�{+9"� Fv��԰��5�I�1!�[��6'�c��F����:ơ��6�udu�,�Mr�K�2����4Hƹ��!�{׫�9Km�&��O �e�n��Z��j2�K��&��c�U�^�Z��Q��.p��Y+���9����1��&5�3�h�DR�4�E���㕻���R��ɳ��Q�cl[�\s(R�]Xlhi4�nFw�]�Aj�b6A���-�+T�Hn^wm��h��[��4�wQmG*��rT���l�E��<�
]�������ڸ��U㭏�}!u�=S7<,���lw�=��:��:�+I�W�r���N&��'+�P/��Ry�e��Yj�CBU�}���RC}� *e�*�KmF)J#�/����>�.���y�l��7���`H�5���6�J�ʙ�o}}�R7�ӋJ�y��cx�}����kIȥ���']����rYR5�ܰ���ݙ:�b�Cb������(c����@@��u��Ã�o����-77���Me���cV���i�I��RZ�]���	�;DG^Qʾ-<&�8�0�W�Gc9�;i��]s�PR��}u�O�?�Ҭ�c�!��E]r;=2!���Y�.�������VXE�{��{��&�9�3g�"d�'H\} ����Ue��9*��hn�Ħ�p>�g¬W��õnv��s%�u�a�D�0ʋ����9�>0_5:>Ty�cө�^�ߤQ�� �}~$��θ��9��~��ԟ��-��}_P�P��[QD T��P�k���Y�K�S ����t(����2��qE��#�gѪM��u �u/������|��� ���P�䏼�,'ƹ�EL]��A0��(C�n�z�9�ɼߪȘG�E��*&�g��wU���~�>u0�蠀�*<9�W&�{�$��^�i]�8���
������=�py���W��k����j��@c`ğr�2�-���5����gK�8�?<�e�#"�DXŀ�P�$~~�>ߵ,��I�f�U�,Qu@,P�����>��%�3"+z��d�dâĤg���)u�.���Ν��!)�@P
a�>�d���Q�g�f��Wһw��>�� ������Rbt�8�=��Q��]�U�]�����Y��Fg]3 ������c�IΎK�L��g�c���^�k����}��	���)�);|� �}F<#�`�����omX�kbC#W��=.�u��Hh��K?nc���.]�5H!�<G�
`2��,&��5ZhYP��p�x�wV�{c�SF(B�n��ۆ=�86�L1�y�o������x9��>��Qdd>]�l1�dO���iNW�tu}/|�˷O��z �+������T���Ḣ�o*�9�\T�w?wN������G*����#Q��N#���D�u���߼1q�G|�Y�p���w�^�!�w����ʫz�!�7C',}׌�ϔԼ��W2��+Jα�]�aK�i�o=X�� 
��R�²���*���}���3*hE6�� 3;��a�ʇG}J���F�ԒTCH��A��A ���C)h
"ֳ���ƛ����bl��wb=��h�c�$G�/J`� �b��Wj�O�'�**��w���z�Y�]�]l:%J̼�ci��St.�}F3]~��*y$�UT�P<�g�adq '����}��;�c��G���F�[`C9�qB�$H�	����Q"K.��$�֦)t����PK"E%p���]t���cg]=���V���ꗕ�/I���KF��i:eT����b�늵� �A6��5��)	S��Ӑ,�Y\�AGE�/%�)"Y.9�I���2�H�C,(x�㢄/��������k�;�O���*�楦&�%LP����C@{�Ǯ�S|�X����=��|��s�p2��D[T��B���zC��#�0U�^:�O���ډ�E{]X?G�cʖ���r��[�,���k�$����nn��O�X�mx_�nm�r���M��θ�L�>�6��e�
�ϕ!���{3�ef{ިct�o�[W$1|J0�:ΊQ}�4�J�&�2�=��r)[\�
���lgtԳ�=�Z�%3�^\*<�l��q�K��mn2���aOc��_CR���K����V��<`|��/����PDF�*z�Ad$a䨰DE4�GN��s<�{�3�Y2�I�5@�~y��|v��ˍ�(�8Y��6Q�Br���6O���O	-
��M_��1ᮬ��M�X:+���|3yU�x�X�,B]Tw�'��U°�;�+�h��z�/�|��;�8C'�މީ���;jɣ�C˞��۷p�y$��A��^��^�ͫX�BZ�ӄ�,�D�J�#UA%�Uon�W�f��O5BTG��Cki��R�[��İ��\U��� ���"��K����K��������q�e�3􈰹���9IaP������%cRoY{�@�:�!؝����I>\������8!Xmb�E���イ}0}B���U����"�SQ���R�Ǝ��c��R2~=Y��@��k��3F��VfB����|��[7r3�q�p|&ZĭWr�����ח�kL�����������\��7��@��ʙ�Ƅ�⚩�Β��zG]{.����mA���b�mL��48}���u���<���~�܏@ĬPc UDW+�PR �P�H��ʟ�M~2U�<Y��0P��,kUؖ���
?�t�ӭ�#�B~^���:�$q�B������}�w��x&w����ʺn���}��X����g��yM�N�����0i�wNo�B��60�z�ݫo\I>�*���Fφ���#:�#Ւ�b"#�@����k�mj��{��8>�6��=��'>��<?�ty��g)���&�#t�I�I�	�|ɔ�f��t�}�]�z޸�Ӝg}H}�����<��u�s�6�d��U�-��#_Ac�y@-�E��:�L��
�f�r��أQ-i�	&��w���=�R�،}5���T��|<��n괊�i���*7�wS �I�I9x�5��~�ݝ���0#�_{+���#�}��i�
K�{�v��{Y>��F^�u��K΄��@�Ävd��x�9�z�{Zˈ>����u}�8��W�Η0NI:�C�{�G�r 1׳�*s��ۇ�]����hdM�J̯�2in=����΄R�!�V�Zg�����q9���2x�`�,0�,"o�_F尾r�ۙa	����Vk� DU	�f�O�Ok���,���`�b��ȰU"�7���{��ԋ�@PF"�z�>�~�{��]��Gd���gȠjc j�8w�?$�����O�i�6��:L��[6�׍��&#��J�f�7�YN��f\ĳ���c����9��i'�>��$��8�+M#���$_���y�\Ό��bՑw���-���C��꺀>z�Ѓ}�B�1{8�#��Rt��0���*�GgX|�L4���	��RS֫��降��<�s�$Ti3�ܮDp�|<+�s�t�=�]ޫӖ����=��6T[܃Mj��C����J�tڹ���Ί7 ����YW^,p���F�q�{������}t��{���I�~]P�Z�o9���WN�P��|q����U5���vh���}I��gT.��{!�UC����)�AE��^�P֏���>�����"�x��Ż����|=U��,�]8�QD�7��oR��/z�x�O�R�.��Yl莣oe���FPrt̙���6�/�tO�I@���+��[�����5��;�����EEE�i�A�щ3�%"������|�>�.wUl.,��1��	
��k��1�^eK��Co�Y�?�9�F��Q37b��m�wM�v����Wm�!X������&�^Ym>�t���>e�����Ʉ'�azm絏����cݾ�Y���߭�/���O£�z��ז�:�ͺ��t�KfN�U�����=���_H+M�\�{� �#˻.-��
�������.�~}X��c�΀��������z���DD8����~߼�X�x�qT-PR�U`�"(��E��i�UF
抎�f���	�����%��~u(L�5ұ�7����W5L�K*�V9���A���@���\��YL��!�\r�g�Ckn��K�b�hw��ՠɞ��r�gu�0�"k��,`���Z*u�Ʉ1[����ۙ��e8{GCēT�R�aqg��B�VJ4w�o�+\�.v0[q��w����dTP7rI��R�N�\~zl�
']r�V���-K�47���~�9�6uUW���>7�X���%Dͷ��Sm7��=�@��(u��8D%� C��,7+�^I�Ø�#��P�ʼ}���yu������x���-)<.ӨZb��/\����*���@��.vg�P��	���4�Ncji�a���gǰ�Fp��D@� )Ĥ���1}���*0"'k_ZؾNe�'Lh�·*c����$��I0���|}\�nꏵ�ř�z>假�|>2|�n)K�6vhC�����c1��W"8*<�نL:0u^���3:�Ƹ�����G���%A[�b;ٕo�3rb<��>�%�W��>w>�K�T�~rw��[q����.�y��Ү��E%W�N�7(���נ�"��ܔl4ڤ�B���;g|cB�;s.؛&Kn�E�+�a����qL��?'��gN��'�$���!��2xG��Ҧ<f���#����WuU��>�>�r�`M��ߪ��mx$�<�P��\w;�K�3�A$��Oݦzr[O(EGf�NyDmc��wʹ����Y�fn�˱��6�B�q7���c�
�V�*�����T&�H^��J�W�*�{����k�m:�3�r���m��>�w�o�3H,C��QsʶkU����\��]�o7Γ�t�z�pU���������xV�6��]��n� �c�ҷќ+]5{�*�1d����#p�꯻��� fB"~鉔"�*���g��b 3�3����|ߞ�9����Ո�� �����M���X�g�j�g��o���W���}��<��]Q�w�M���N�oV�ȑ�ԩx�M��Ĉ�������(����0~�?Z���+�w'�Q�b-�:���E������[��{�K���Ԕ9�+����d>��"N?'!}74���B4��n�Uۏ���b�*���ʪ
*����h�*�B����W^�r�p���B*�9B�Pt�<�zF�a~yY�*����ܯyt������������q3�a�1�Z��y��_�1�r�PRa	��X	-
N&������ߕԬ�9�`�����m=4.V<��xc�P���F�..��$�CsNxv{�/�r�}f?;#[�MA��%x}}�%��י\�wU3�m���N}�e��7�f�8�0��|��^oN��Wv��HFfjvW��L����X'ӣ��ڜ���� IĞAX����%? R���!��1����{uY�Ą7$����=_7���
}�=:k�h��7�@1ay�g+�"��{�p֌��F�WB�������Z8�Ԗ�pY}�W�3f)O�w��<�}��\���k�^~����s�Я2�Q��׫�>��wK�����aܫ��Q5��i��{[�]iwr�6��U��q>h��W��������~^��]��Iф���߾���u{e�˯��3�;�٢�p{�^��F�ڹ�9�3.���{�f�9�k�4�ְ���V��M4v���ވ��|DBa�!l��e���ě�c皴�xle�m�B<�4
�pa˾c{�0f�Q��!�H溗t����Wy'4�kW�j�"Q��LF�I��p�swS���!��C�������Z7���5���kq^n��f�s����գ���_!P��ih#�]���,��N�Q6���;�j��L4!���
3��n/��s}�s��Dh�<���%��əy����X�"��!�X���E��Xc�^a���P{k;^�#3��v�V��Ƶ�	39��g~��I��;��G{d���x���
����Q��z��P��ꭅ��舂X�Pc�)5��z�[c��z'l�ȉ�^�k}]����ǽg;2����v������J����s�r�]u�&WS�ߊ����c&���k��<�ۅ����c� @ G�� �#��z��9�t��7��SỪrbֽYϯ6����`�׶�k��j�aE� ����Ѭ���^���'o�]�������ӱ�[�`U_�R���5���\C9�=}?�Pl��%�qmm̬���q�,2��\�R�W5�NoTP3�6��]HGYc��s�b.���w�����ieF�7{��&U�K-e*�:$4�b�����mV�h>����� 9n�A1{F%;����5�I�;�N\$�	m�)�X�G�7u������s���gG�A��j�GbIZ��$�f�����c5�r���Q���C,d9%�y�.KiqW�j�*�}�y�8�����.�\��v�Mv%$��#j�J_X��9�Ɯ���K��i�N=���U���Ϩ�7��~�k\��\]��.̗�k��O�j�*pgr�L�\���Ч4]�6z�*�F��b�U�ʭ�,E&�I���343��#����;F&�<2-ſ��b�m��8�vh>�˕3�	��P�N˔0�÷���c,<��*�`Ko�8V���G��\U�y�pn�l�}��ݝ�;��"��:�I.��Ρ���3ni2�;]5��
	b;g9Rܦg.��MM����7o��}/,*��p<��k���!Z	to�Q�*�s#ެ:�EP�������ǹܰ*]X*�R��G?7Kkk_VU-KD�L���2@r�(Yk���`V�u㹘�5�1��-�٦`�X��T)�*�
��B�}ECY:�Y�ҧI:��yH-�{+�̩۪'���q��d5��X��0���Fڅ��h��m��m328fC-ƔƉi&�,�\���3͢�H�ZJC$��I8ےI$�I$�D����7e��2�M�\I&�H��am�& �,br�ҁf*�#A8�7L��2il���Ũ��GB�^�nA��3!pol�b�Պ!���2/���1+��J�kZ���m��kM���G4�b�3(�ֻ$�'-�K��3�Fn8*�W�j�/��2Y* ��*��@���D"e�{����m�h��-%x��V��pP�/V�9���2�$�U��b|�9�t�T�6R�UGM�Bc��6�}#������O�,�+��&�9��%c�Qv���ә"��EO���/�:�[��l>s�6-,楀����B�eb�3[�V�V�~��*o��URo��2��%�1X,�k��Ly�^�J�	uq�Y�p���C�e���e�����	���d�z(�j�r�q�m�<��^hGiJo.׻�I�GĞWE(8iU�[[oVTBB41�?ZWo�v_2�/E�eVW�1�m�eSѴ y泃#<{U�uK!ٖx˧��i��g&��!�!Xj��is0Tټ�-+z�t�㝯MLpWK�FCEi���{5)�=ɕ�kf�ev��'���P�/���Z�b�6��:�Xc��	�j0�%+-���
VnCP��Z4�r���9�7�Hgs�W�;8q��M�uツ��=�#��wl�H�'V�)�y�ٖb��^�[h�	е̞ �G��w��޷��i�l%F��+q�W�!ެ��-9�uIȓ`k��M�agb����^��]�!̛&w�1��F�aEBP�aYH�1M�t�w�,�o���a��Y�yW�YG����m��P!	-����5᰷��$���8�Il�"1�$0F�(HQ4��"�J8�@�I1�#��-���4X��|�+�R�oc��.c>���ҭ�y��J�Z-˩v�i0'ۼV�L��u�v`G{��	a%!���(�o�5�䳇��TCFk������!�E�u�EҨ�bB�7BB��A�L5*����%fM�ҽ��Mzä�l�ɌB�~�}�A{��7.����ޫ�{�C�uM�r�{�w�[�L���_�}���P��������y�dԐ>�+��(H�ÍkW)
dUI�0H1��M��
,$`�]�;�^�+����F�=�ճ�t�����C�f�����g�O�م}=DP�`�^}�9�^�z����{��4��OH�Ú����w��5�DAj��y�-;�^�E�~X�K�;ês�.H}d�u�l�����=����l0�V��h����w�Ƶ�t�Ctʫ��J��^F">b>�>�|""-��>��։}��pWl�-�=�n�����{��y�8��>�/+���;����������Г4ff�z'?-�1l����q~�-�#��}�=[!t������u�L���+^�6%��{v�&3'���T�v��_̆Yl��D/TK����%��݁�.������bh� �S�T��9�{���|P��3t�C5��-h�ͤ�wB�{J��[�=j=tAo+X�#���ϴ׼�b?Qf1ϻ��<��꽸i���E�F1AE�h~K�ȋ���㏶�����,D��b
 �F"	��}�u[ 1�����'I�x=톩ǜʵ��V^�xm���=O|u�Q�o^���O��2��zǹ�%��\kmQ��-�j>���s��࡞�X{��zj��9�/f;}ڔ�=�@�&�k��{6�s�U�n�]��s]�s���qN��t�����߿~����n�����b ���̚k��H�U%yv�H�, ?:5���k[�GON�<H�e�-N�
����jg�b��z2}��9w~��@���oP�-�(�oӷ�)�o�w��蝔� �3c&_�rĵ�n+W�M�SK|2�S-k}��D��.��b<��>����#�>���j��Q�{TS��$6w���F�k6�$�����>����rW`�7 ޡE��ڕ�nOǍ��s�aи�EW?lنf������T6��J�]�>��خ�����>�A���I"Z�1�}�}�g5��E߾�m��T�""�"�R*�ŧ��@
�j����
�۟�?O>�~����Er���J����_����Nw�����m���s��IGh�����CZ(؏���%�/-�-�fx�>ͭ��x����T���3|�&z��J�2[ju�b2�>	T��~����3L�Y1�U1v�����ǂ0���Ny��p}��l��뗜g����u̚R,�	">#����|�ӆv�wb�x��HɊ�Ƥ�8<X���w�{m�~]���b�s��>]#�����=�?Fe���-�"�x�~�����0�xw�ny��P�����;t��R�1�T໽~��ɷ:�_{�>ؘ23�X|��e��V�R؞k�3u^�O����Crע�X��뫂���[���s�>ǽ����#'��I��T� �,���CL2u����R�-���J�P�y��6\��a��6�TV��x�D@xY�b�g��|K�ͩoFN�v=��SS��a�jT�����˻��Xu��q���E˝Ժ�c{���N�E�}^�ا�eyt���2�Ee+�pt��r�[���n�_�EWN��so�ڗ��:�u�Ս������\u��\��]���.�BND��%
%�_UQ>������G�{�f���N�f�Zx�=�������W>�2�o�o6S�2��o�u51�x��B�6=�ETO�y��_z=ʡ���X��v���"!}���0w��)E��X��[�~L�Tt���޹F�+��	�m�dy?Qٍc�y@��W��?�����C�Sǰ��+��CZS~�q�Ьn� ��舂������z ��_VO@>9:jo��"Ղ��_:B���]�G�༡{�(;��U�zSeL7��~��锊�TdYH�`�D�q����s����Z�c�^+s�돣��DDC�:dB|�a���d��1���ۜL3x�y�"�ܲ]T�^�g���3�ԳEZ�5A�}Gޢ4�O��ԒH�M4�P��r&X���R�.�����J��L9��kT�C	�OT`�Tn�T�c�:p��ՐLS�jQ�r���#X[,m�5�{A����rE���ݶ0�T]�j�	�lkb��dB�`T(�0�����&�&0SL$!n9�m՘5A�d&��c�BO�RՃ̺=���uݑKq��/�������u#3�x���T��ʽ���pr����}�m���������+���`��cu�IŎ�ƶ��nb���B(|�衣&x���3�O���x�v맕y���]+�#ȼ��1�9�k��Nw����"D"�<��0����3�s6��U�v^�Kpƥ�{�(��R�nD5X����߮׭�{��9�����o{�]���3puwr��X���7���Mz��,��H����t}��e�_'���z����4Ƿ���I��c�\G��n��5��J1;���8���@���u굅�f���U�����>�c�R��,�))��{��3�ܴ)(B"(�,2*"���K����1b(��]f��`��/w�%�J�>Z�1xn�y׾��������<Ⱥe'ޢ��E$=�!��k�sc��f6=G̎>���]�n���r�AY�T n4�j,�45<�p�@��W4Z���ŇVޮ�=��[������<˵�W��(�DD�� %9��轕�O��W!LY}�ڟ�H{�V��iU�s�[�|�t��6�ħ�*��o�7�G�����K���?dn������o~>��>� C�!!�z�/�_s��SZ�>Q�md�]�����^=��]�%�	d���@�n5���>�suu�2j~�f��B��WJG��" [Z�����7����!p���]A-$���zհ�Vl����!�y�߹-~�
FM=�k�`+@�����ّ��^X�GNf��[x��g�v� �_�5�^.)���U���cX�DAAWj[EAc��"	z߻Z��?�[��΢}Y���(bJ��W�ܕq���o�����-̝3@e��^�*��F�\�]ö���X�L$����a�ۺ�h7��G��}����>�O�Zj��ٟ��9ܼ�J{ˤُ/>r�B>�9�Sg��)��`:9d�ba{2b��[��|�-&��UUKN5��Ž'���������^��]����,R^�_v�e+��������=�}�/�b�5g���{�g��z� �~18���q�	
8��Z���zk1���-�])r�>����V#�..��h���ɬ�0  �ޤO�wY~ɘ#���̋���5���K}�8g�V�l���k5\���>��tv��1�חn��D̈́�D��O���q���d�m8�$Ay���߷;{{�گl�m�s�7���k}�k�5�����8�X��,�T�P �c�Z��� �]����ꡀ��q�і<lĿ6�
!;���}���v�����o�5h�Ҷ�^뀦�_}�b�=y������x��UN�9])��2� 8�kV� d��岻}��x=ɇ��a{���kܭ;�j���2� �P�G欁��q�D",nJ�Tv��M���B "/x�3~p_�ݽP�����n�v��3f��v��md����xf�W�P����J|�,ȓ�>��	�w�ϯ+��`���z�����뗰����˜o����(Ϳ=�~h1�]�}���=���q!7\'�݈��Ac�ο~bB$3Ԙ=uiD^�lk�\��h�©أ�t��Ba����n^,X4�tv�ך�c�ߴ�}�[�k��9����u7�	y����h�`(.-;X�o�=A{�w���8��g������{f��>Y��W�d�瘚�Գ�}��_|�8��0r�=K����K��Mp.,^z���Y�u��Jޕ���rg�2Ōa�dE(�D`��C�����[�ӷ�[���~�g��=��`( ������� �H ������îf���x:���mc�Y=�q4�e��U��˴�Z�˸�U �Gx0fAd����bA�qs��G�""8ۍ��*�������C�v���3��*8}�:���e"'�F��T�a��ȲW*Ri%f��M�^j��u�����q�e�Y�@�(i�I�H�. ��$i&�q�0�
���J^�y���V��8�2��X��VP_h �����.�Dɑlڊ��h��L����wF��]x��w��%*K��,���ШH��2s(��	\a�}JZkSتn0��$'a�� �2���A-˻��)��n�T݀���Oަw;Щ�.:�u�ս�ە��SL�BV����X�Ж�� �!����ry���߶��:�how³�KO����M��U>2�W�Я���^.�Wm�#u�Y�.���EG9�D�ɗa�긗�;d����V���k\�9�8�R�+��p�ӭI��}.;�Dt��H�0�~�'(ݧou���}Kϳ��g�;�z'j;ǝ��Y�N����>������
�DUA�͑��  ���m��m����8W;hI��L3U���!-M-���a�~��_[Ֆ�b���c�s�]xTe?~Cwʹa���j��M.�q�QZ#S4J1���(���}�mE~��]-}�Ѻ��ˮ��o�t�t���G�������U
=W��qn%M�7>]\�O�}e�U�a �O���@;H�*�M��ŏ-�["ϼ<Ͻ�neI��Eu(.��m�W\��[b�7�����MP	�M��Nt��qC����}��T�?�y}�Ɋ�����ɑ��D�D"�Q~�	�����o��%�g7���S������g�ԥ5>�ʍ��/.��9�ו1�D��hIu��,;>��H���`l��_^,�|4?�3�D�Ozu��	�֪݅�ƣ����;ESU�0����&��y�©:�p���8 ��6��(���󕏼�D$X�#������X"D�sƴ��/��>}Y��P쐜�]�t�<������y�-�$B���_X��\+X��%Ӡv	P�M��n/��~�ߚ^��G,�����q>���������2��W�{G�)T���r)xG�Dq~�{A��\9Q���$��vk�HO5]9x��kTq���)E󛎎�{��N׭�o����J��틆�pU^�գ=ۑ/ק�B���ȩ�f��+�A��3|߸r�JO:���]@�Ŭ��P�nM�3���+�)ru:�R<�ϓΙ�ܖ�9�!�<+N�Qz�	�R󒞚���@�Zs"d�;u�}�ﾧH�ɇY��h�f�e�����|����;.��a�ĺO�F�x2�%�R.��g� F�$1n�.�*�c�ۭAF��p3^��y*.���JP�VJ�u-{y��po%�mq8m�~F��=��D���� 7�j+$���g��o8�		�4y]�����	��ԫ�~��G(f$�ŉ��{#!��	V��˸�쐳�鯆].�yN��z��n6z�/giPI�d��
�=A^3���S�^�LX�yl}�l�ɇ
Ҹ]'A�*�`d��H��o+���}[���3�S96r�$�l��ϯ�9?�D����?.��K�;�Q4�h�{Z��q�m�1�������]����n�nr���(%)�vy��mn���ڳ�3�%g������u	���l,ٗ?��6Q}" �f��~,y]H2�;F�6�]d���:�z.&'�ݴ�N�A�z��h%I�a���h=`P:��V��>p&E?�B�墂k\�̘��9V�֊Z��yw}��a�Z�\�=tO?h��q�����3�/�[tT�C�3�K�"G7��5�,������x�74:��gxɃ͵w��~���Ԑj��	1w���h6n��0��={z��A�&Yo���l��Iԗju�f��A��m�֗+;��y�����s��DWr`k�|;f1�U��O	�J���߶ �΂t���g}rp]���Vs�j��yk%�<;����j�C�p�S�L��+���T:m.X�Rv.��Y�F��r��Dj�S�b[����;GB]�]�X{��OuEle�u8���خ5�;{�^H^��U�0�R�gd:�o]s�YO�G���q�s�n$��6�n��
�s�=k;���le
����6�7U�p�9�n��5p����E�S�Ƃ�S��hd�7�f ,����f5`�rI�����ڽl%�����ݑt:�yI���0��s4�nn(n-�*ݶ!S)��N�E��}s���3� &����MGS��hޝ�0Ʀ'�����&�a�P�ǻ4�Oe�8l=܇���,�WM0�(�6�n�ќ�J�Zҧu��V�{�ju���w{�<���0��.�.�o�#��X�Ok&��͎���tC�x�j�}�X���;�Н���;�����{.;Y�u��܍�̗- ��q���rTK��s+7�Z��m}��i�xQ�/!��i��m�������)��y��s[D7u^� ��7e4��E��V�+:ud3��r�Mݞ�;�-�QeelΜ�3�j*����+�L�辦r�����Ti�n��;7h1y�,�~��<�9���o�<\�ޝ%��Q�}$F����*I<^8������[>�����)gͫ�{���_}HJ{�*�t����|�s{�J��Yl�K�Z��H�5������B�Bh��r�*@��q�7ٸ�w�����F����k�g����TX�� ��"+aETI�)�e���u����T*���zQ|5�Y�62���� �J��N{9�1�v����M��(,��kr�!�^sz��_�T�����o�x��j���N�ռj���fsQ����U8z��/竖�Fq��^�W�Rg�U^�����E��ǾJn���2[�]���kze_�s_e�B�����������"�.��ז�N���f[��?|�DY��ϼ�D{�N�1�j�w��j����H �	�o����J�����v��W�k�d��c��m$��݉h�q�krFbr��-�.�꾒�����/.��TPȴ��I����k�CеQ^�W%����=����6��S�{]�ii��>˽2�.aͽڭDzL�0��&��ϯ����m��+%H�%|�l�qAķ{U���f�?7�3���o��D���fӯ{�U��_G�~�M�H~��{���o���JH�c):�1DU��"�!�8!c0v�������N�?`AX�FF0��}>�v��Ƒ٧��<��QT�F�(a��j⵮���Z}�`�v�9����dO(�\�n[�N|��g�s��X�~s\���}u��l�w�����t�r��M����P
x���Z���%R����.t��ti��5Wޚ�UO=I�w/E��w�>Pe)u�[���'s��p�1{/�פ�yd���1H�������_W�,�-ߞ�)j%tZuV���::=U��VEW���)�����C�0��������?=�3�[/O�n� {�t�ҭr�H�i��nI$�����l�#n���@]v�Z��8ӱM��wU��uʆ T�x"I���EپS��UK7n��LȌ҇d*��b�J��L�l�㦝VH� �x��غ;�Kn��%�9�B)R���p�IHBӈYN��5m��b�Ǫ`UQ5"�:v��q<�}j���<�i�c�s7]�c����^�j��� <�������c�$u��E�>hS��'"s5����T=�{�j�ทq����̙)�O��O��H�����X�Y`�"�a(b��UU�/�F�w}5KTI�_L��{�����B|� ���v�{���g��y�^y�p��;Ū�L7�����tވC#k���6�0���QFH�f�˹��>�su(��J��|-<�
_q/�G�>��DzUg���w;ąd�ݛ��][��zK �B���Rp����ª��|�ݘ7�����ہ.�{G����}��u�ߗ�;��+�gZ�Uΰ>b��L &@�l�k�%�d$W*�	�&�?�����xd\���l8~/�*xm�u>�^Z[U��8�3T�.K6�����e�zA�z���N��F?�=�?p�h������s�٫4)Yݡ�T�4ɖi�f��
;۳c���]�j�N6^�T�µ���[@5b�䞓�����U�m9����ڹ�ʻ��w{�n����Z�tG��\|��l�}��yv��!��_��o����a���A-oYmˌ�F���ӟX�J�ׇ�"�':�a�}���vy��kִm�C��4�Hy v���������}5�{�c �M4���*�p�l�� �x׏��`f�/&���T;i���+Ow>��D]�gR��x�w��)t���7Rg�gTVz��^��S���~���#�5�}��[���ӯ'��^��a���_fw~Fca��6.$��X	�%3�<M��D����N�dV�ޯi���dC�d���V�s��-�pֱ{E�.��{}h!# �`"fd ����X�*a������Y�_Js35�n���{zQ;4��W�������s�4�4z���w��!@���Z�K�`8lF��}�2�1�k���>�$}��8�i���>KC��l�^Jq��k�]h��Ov=�����@�|��v��fa$�g$:/҄��v=���!d���:���B��c7T$��^�i;t9G<.|���ÿ����h���n��fF��Boe�{߭�<������}�3��J��9��n��    b�QԢ��QH������ f�uH��@T����YDF���;�_��}���3_K���//�9�G����zm��>wf%���o���w#�+��jF^�C��N�	GDh����~����	�D{�@}��c����}��G�^������_������Y5{�W�����_����z�;;��s�Rv��]�GC�.���h��1mF�;�ӷjui�]�
���AY'�e���s�W��_n��w�;�n�oӽ�WOT�!�x,b��u���=��Z��۷�ޘ��Ͻ�}�鮽�]�t��Z�N
���/t�1�������jK菈��/���ğ�Ӯ)o]�}������vi�M�>fi�$B�x O�!�S���U�u���9�ю>G�D{Ë vtp�g�C6ꁇ7+���qK����odۉ��G[�ږJ�%�r�`6�we��9�̵7�-���VR�l2��B��/S���u�;��<��V �A�����)����Q�{�{�o���߽����u���__C�Ƞ�R)��"�|~�>�N�;�+���#V��Ⱦ1�ߺ- "T�
�"ꗕ�(n�~|�� ́1u��I,~n�9��H�em���7#�z/*�����������o�+٫K��|�O��ҡA�5s�>�@���}�dT���o�oز��~���#��#Şb"{ѩ����S����V�q2o����%����`����W��/y���v���DDC8}+���y�\'_u��@NAP߽�D���忆&3.��~_�Gcq�z�Nf����7�)�7G|Ԗ�ǘ^��U�6�U}:�7��jr�%s���ٹ��z�W�Vb�on(��,��撻��������Ri�:��_$�ä*���X��u9~�Wo��G���x3T�����q�b0�RNY@��e6S�%�!u��}�QJ$�R1���yo��Ӵ���F[HeRD&^��xkM��l������n�Q��@;��y�\���yi*<!0�͑u��a�Mj�X�$�	H"�*D�i�L!2���PmX���$N_*-Sa0�D$��k��ٔr����c���������!���P@db@Q�G�w�j��<,`��b�b
,/_U�bł�'��y�YU���^KUk57y>zn��L���u�yWc��rS:?���OW��6#v�����ns�P��}g�⢑�����{�D}�#��]v�L3��������>�t�f�?ws%�����E��[H��x����L��O97+ʴ��zp�m8̿Z�˳���h�v8;y[F�$ ���3�I�w��~�r�>�]�+�E�����7���PGi6����=ف麟�r���ˋQ���/���JX�E�������<p^�"5��}>�խ�Yo>�(	SNnlǽ<�g�`y��JGt䎘���Y���2=�|�O%r�cQ3@ƪ����Nn����O{c�3�l�ֽ��*�\�s���{|�٭_�c��j�e$��S�T�%=i��:J�m�c��ۚs�}���do��un���dX1�@��>'� J�஼x6�7|�ޞ��
j���W�N]���(봳{w���q�W7n�U�n��ľ���Y� "}	����J�S�{�0�-�E���yu��<�}����9�����K9�/G>�	�*l�gM�s���K�U�ʸ񈏷�i�Q���%�B��(��9][�8W�f��9I�ݒ�`���u��w�@����oϳ)J�xy�w��0e?�S9�,����D{ﾊ�~��A� �r2T����u֌�}���ऐ��>_,�"��O��x�.����'��p@�'�0�*�_�&tp���O�w��[�zN��S�7���Q^l��3l8��} }���x�w�WkRA��T�]�ެw5])͊�z^w1�/&<�y�]^���@̣&j��yZ<�E,E8c�cl�Z �I�H&}���̿���M�}���4>c",�2TX(�k?HLgoy����������RJ`Ke0�E� x~"5���_���ɣ7�7X8�HJ�u$-�N_5��o|���oX7�v;�Q��Jͼ�J%w�8����nv���\����{n!��/���|����Z�Dz^J�#����vzf|
�s�ٯM��W��q>�os'[�Q�������/2��mK�)��c8���h�l���wAH8VȽ��*�ۛ�!�#��7�zfO���\�;��Q�'����}p�dԈ�f�H6h�P��g�7EI#���׀�� �`�"Ȓ3~���{����{����vW�+���{�W&�T��8�n��۪9[�陞�<&�ɶ�_�8ZT��SiV�v��OSpf����h��nUz��18vk<}�[�yC%T>�P$�P��5	���G"�R�����dv�ų��>x�u=^��l�^\Ykw���ߩP1Dc�C��3���g�s)QDA�A� RTY�)��Q������︭���f��#�Wz�����*3lo�!���>�{��𔰲�Z���߃�]�s/����}���D#MV#��v�jVv�^��.M�ݺa��)��t`<�o.��t�kf���99��}x�j�4϶/W;1~dw�·ͤ��v���W�>G^k���V��}w�P}ki���~`J���ჲ�<����m_���ӝ<-��j1�����~�����Y�WS�<���5ܰ�zVj�-�tnn<t�-��m��Q�}��>���{���;�����8��3��0_�Э��;^��s{���M܁�<���mzc9bl�G���]]���1՚�Q�2`=�۬�}*_�|�xOt��@���f��\׷=���"O����*������[0:���r;�OG�gkR�<�f�!e���3*���������[<É����`�,c�Ec�V �`��W���u�n��I2�Ȳߡ 㲣����c�P�"���]���>n���.�mw��))�[K�E�·+aK���tjͩ�=��S�᳙�@:�*p���5|p��+�D���p��C����v�×�/z�j�,)Q&������jTW��npG{�j��d����>T�cBU��rW�-p�=���.�1aE6C����`7D�"q��*V�!l�!^��3��\�EDq�f[�ux��Qu��n��̈�P�3~E0�7����в�=nN����<�z�D����Wh���ȵ�8�Ҳ�+�����^�軭��=��n�lP��h����e*f�D�����Z�C$"�CT8���̦��w�E
����ֆ�S�!�[*E��l����`T%��v�B�^�Ne�m�.�u���/� onIi��[�{uw����LR�.��լ^�v���vdm�F�}��������Pagp��q����j&�XE����m<ݎS�U��'FS2�k�7��7o,&�C�}����;�~����B�N�֢�l�ڙ�\�B�6Bbs��z+谙p���$�psղ�]� ��\�J�<Cs�6�1�oS)��/ 7�Rb�lG�7I9�}�B㽎�h���Ǝqn���V�*kb�A��_�r�R�N�|��L�q�ٺE^Ay�J5��F �FK���9x9a7���(X�bTF�;;6�ݳpou;[Q�j��b{MYC�@���N?R����m<���ȩ�[.�!݃�v�i"d��T�9-��m!�N�$�	��a�Riȣ(�S,���$�"�-I#17I��P�Ò4�H�H�'�8SI�[��n@0���nE�0 �nE֥.Հ�tKX��x�t	�r#wvgX1���M5�TD���z�^���щ�傣b�r�	U�:��s3<�Rr�BUR���N��p�OuVi��Z5��Y4f"d�%+Nt���z{v��yWPI38Е�39���Rf!���ړ�v�p�WJ���ycy�Do��Uuwm��d뛮�bw��sN'}=(���NF�7Z�dۅ�X�ɼ��i]F-�RЩ��,��o�}�[�!Q�:���r�:�G6�w���[\Dꮎ�U��B�W� U��(C�Ի�(f�q]I*!��ěy@�uHg �,e�y(e�2�D��v�S^͎��7Rvm�3�k��v���F�;�u�������8��}�7ʌ�r̜���5�:�h**�o����^s[K����v3l��0��|f۬M��[�.�_fc݇�:���8��U��͕��Ěj�R�V�T�e���*ﱹv�!���b�5ɕ���g ��7R��C���޼ڂG\h.�����<I���VU����%�d1X���u�鰃R����+�=���f@��'�Y;�6��,Bz�Dj�N��K9���9�K7a��.�BGP��=@�]
�J��y�\���KvTJ�K����z ��`�Uf9ia<oC����ն�Aa��b�o�5}�U1cQM����s�+Pt��+&u��=.{
'��	v�q��[��^�KQSu�Nt��X���(c	��{�%�;�+Ҏ�Q��Z�;S�y��z�i�m�XE��4�ݲ�DU#�<�SoJ�[����a$�x�j##Fb]UPP1(a`� DD�"2�nI���(F}R3a0�(�JE���C*!)PL��Ue�iL��b���f����e�NVk�d��щڝ�)�X�6�՘j����=����iV�@Wg[GP�o��q�S�&��Rf��0�!m�uB�MRN0T	�A��2L������ t��Zl�0�g�:���(d�dx��>v�/k�^%��U�S��f����z��ŵcW��sz*���(L+������7v%������k��A;���ǽ�&;u[M��� �*Ȣ�PQE`�'�U�������ssګ{7�yS.����;�;���Q%�Z���av�'�1��0��}��"��vLH�v���yC�.~���KdN��u�s����z�>�t�JԽ�۸�嚹4��>�}��y��?����ݭN�Q���K��'l'�E3�����KAd�i"���[��A�;s}�w_x�s���<��W~=���r*�( �	�| M���e[��ٷ�L�D!��@�MS�t���0�v����š1Xl�6���,�j\���FG`q;��_rlW�xxC�~֟�y�`~�_�
�|z��R�����(N�uW�`�S����@�CW�K������?�'�{�ʿ�P�vܝ�&>Z�>m>��4�۬ŗث�oBrȭ�c;um���\u��t3�;c	��9S�KUe"k�E+}��m�����&�<�\o���w2����Y�����}�c$C�v��ws�g�Y�;=W��z��~�kP��em�[��s�{��2 �`]R"���{���/!ʰC����l����'�����]�X�צ~�
S����GG��\��d׷�W.1�p�V�0؟GaJ|����tv��LT�}}~�p�u�u�p����.;�>�O�{�]�K�T���fuǗ����i��{��f<:H2��� S�𢩴l㍨Pp3s
韫�nK*�x�گk}��� pb�ʩ'ޒ��o~�e�(#�TU����1"�
+��9���9����y�2���}�~��r�~�A�/%��>M/��]ے��gУKgG���[7��Z��0}j<۱���-+��>�!;�5f|��]�:[�ϳ=��'��˅�a�_�Q)���NUBٔ�d�x޽���X�a�˷�	����2 ���yw�	��ZҚ�k �Ҝ���me]�ǔ�
)��X-)����߶[�Z�(��Q���{*�5������������w.�#�Ÿ��O��������r���"��*�!�{��.�eZ�x��bk��f�������Z����Bek���o���{:��w�9ϼ��C���>����t��[����[����(��DR�)�5��r���H �:�	�ލ��2�v������i�R^ht��I��3���<�򿼝��[i��z��	�y��;��/��A*2*�������`*�����>�>��!� ��C��g�SSv3yK�f|��=�ee۶a�P d�;����4����,�۞Q�[��=x�^ɾ���'q;���>�}��P���Q��.*~�i- ��S����o+"��S>�>���6}{�>}�B�:�L�dۆJ`�dR����t7�=ظ*� qZ���qj�S�-c�M㣺;=1>�+5�o�bYa"�ofV���Jt�ԥuwdf#?XÉ䉃�G4��G�zǈm�TR�Sxo�V��:}�k�g�A�+ٕ�7xw�{_g��{�@xr3E�[�J��ڐ�n}F���?aG����uS����8`w���@K P��$ЂhN���#��К�{�sj7��#��so6_��}����sT�ǝ�/u9����:��G�s��;g/=�m�-��;��9Q �#B�:X~/ y{�r�V�Wp�~T/������7..ʏ��}]�,�}��|�a�rC7�w욮ku�Y�}��ب)�B0UPV.�X� �:�Zǡĕw<�x���о��4D�o�f]�v�~��^�ޑ�Չ���=��Q�+��'vڳ���|����f�S�x��r~��hKp=7@/NRM�}v�H�^:}���i�bK���iD�CYO�ys�z�'
=)�O��'U Eb�X�4��J<�^.[���kS>i�T�PQPb��D��A�IΚ��X�L���yLٳ��\*�De8bB�$�I�>��aVP�CQ�\qnH�k�DcE��P�B�K�*]d�x�[�F��v���ݔ�X��ղN����E��-��)\�u&�:��D�ev豶�0ƥ�lmk1FX4��ل�mM�E��:�Ύ)}A�"��I�s�`:�lX����i�m�,�v��x8�C�Lk��-�C�pd�^(�����j���u��f��W{U)��J���=�����vob_ �yڄ��z�!��&��t�2u�Í$��d�>�M^�cΟo�R}�UU�F_���Y�#O��ꦹIM�f�v�L��=RJ��֋[����b��Q3\�Y>gA�;�����Ƒo�ݼ[�s�1~�k�|{w���>�>��nW>@=p��21�+@�R�$QA`+1���{�AbSB�~���o{����c���yA>p��p[^�ێ�o����������Y͊qa��(�����Ǔi�����v�ǐ��������^���z�/U�):��b닜��尧�1�<eU��$�u9�h[�b4��^:�.��?gw�J��}��<�����{1>��[�7�j;��z̮�Y���G��f��0Mo	��# e��w�J�7��!h�O��0�U܄�|�1V>P�W���t�F|��Fc�o��χ���=�׸�E{֯l-�}c%���<���;�n�d݇p-xٔ�q^���]���뙽i��
1�M_�����r��Wp���,�ly>��{~^��v5(��"9�+V�ȭ���v��LD@`�B���ů��~�ݭ}�)��Yb�]"
��K���s��VlaT��g`w�׭��/&�W�멅��c�-��\��r[��/`�} hN�"��"EH�UbQ(R����) ��]}�g�_�u��Ͱ
B |��$妵ϼf�c�ӛi���vh���ˣ��>����P����9�.Ї��M�b�S��Vy�e��h"'�����
�$��D~�\�M�WJ�ƪjS;�� 6��}A�;�M�/K�>���Y��x�c�D�S��u����('�����h3�5��κ}Y��#��nz�8��;r�C��#��A� � �AI������9�m��/�$�LL���=3�pq��o�/~�f�p�B[�
 �m$���<8�̀��Sv��\��Wn	���x#Ջ�̂ד֎f;ѧ`��wUs�0U�0l���X������Z�:>�$t/rV*��ӛ�_��r�?vz���-c���h܏�j����BV0�{���4���	\��#3��ݱ���%� �r��wHN�ê�%|də5�1�G�:���j��[�5g��g��1�^�����=�����dd������ϯ�W/_4r�J@D�����j��%��E���uSh�*���@�W�*>�B�Mș����c�mE>����+ �{6�V�mc�+��W���>�;�l=U��V�,e�(x<<�{z���^ux�7j���g�����<�����keMG�}�q�Z3��ɓ�*�{���p�u��^����}7�h�zy��V>�e�����}�>���!��Y���	
1��+�:�����v�W��WG���3����i=�oG�=�11�58���� �����CL�N>�|��s�8�^1¶M�Y����Rm���^u�{����`=�X�n�&g0��}:�L�8VK�\t+��wlC�<��ᢌݚ��g�'��9I�����������TUu.ϔ��|��RT�K:/q�u��׏���"������T��&:=w�4�UEI1jCO�nh��-�:	�M������S<�My{�i�a�;NF�-q�����"�"(��@+���1��I�1f�QC��f��g�_�Λ�J65sW����<
�5�\7��׎�y07p\���-wo��Q�O���ڒ�G����v�����˷���k�������%ע�����N��u�^�7�e��9v��ϵ�kv��F���ӽy��s:f&SC��y��m�Z�S�|��j��q���s�|6��|p��D���ϻ﹐ԫ�����|��q^�������F���7�{,���3>/>#K�Ŧ�	��k{4X�F�+��,���W����{�	��$�$)�4�I�q�?4H�jȄY���_�!��un�x�0�߼6���I��!��m�E�!�כ
Oiݧ�H�\�����L%Ҷ�S��'�l<�B����)W�Kf�H�4Y� ���!�Y'�e���� !Y�Ī��!F�!W�2����dE��)��U.�Q�WW���$��a�$���ܝ5n��	AFd��|�֨}�zZ���LݾĿvwՙ����K���(]���2�\[K_��$i�͙ﯾ{ʬ�o\�n��DR(�VQDb��b1B1f�|ֽ��~5�w�N���"���F�~�Y޿=����99�'إ�����k]�Mco]��(�|%�TW�f�Bj��
��>��V��M����?!��v~[���:���a�^Ģ򿍋m��̅�~�s>y�Y�nv��4�³��mҫ嘇��t=��rb��t㣔4��ݞ�5B@�k���+=���P�b���O��o��sX�x�|���
`O����k_Q�!�~z:V�8�J.K�P���O1 ���3�5"����r��:�R*��s/C�|%\���w��1ǹ~G���N�s2$��|��F��n���bT,�8���u���	�l'*��0�!6��xlS\�V�!Cy���kq�2P�a�؏�|!�@{H��g-\�=�}Y�����Ǟ�������!=��,;2���z�Li����wFy��M��o����mǓD�\yP>^>��n4|��Rꅊ�(�?�m�ע��>�<Mk;�{S�u����EQe!QPL�(�~j�B�@X�,+V[�=qeL֟Bs�}�TԳ��Ī�ik �A*�OpO��ϻ��.�bU>�o}\�_�]���.��^E���~����S�JΗ�����`�.��7�:�G.J��9��FǴ����2��{�~�À�����z�W�Yt�	�y������`��oBG�UG꨾j�'�M�!.��B� �~T]������ {?o±����1dvmgaՃU���&�D��A�~>�}�RK>1���WWv����Ff,������K�+�-��=�1�Ε{�T��g�`0�>�����pW'�~��y�76�a��H�9f�K���WyB�uX��=!�yFtc���a���!��w���"����J���������V d�P�0�|�i�k�	Y���e���Η}�;"��cS#�m��ߡ�͝k�w���Gpj"�81�vF��y�[v����N��T�GT�nlc��+AiTLZ45J��9��^L�=�g'�_zJ����X�2�}w��l�e��*��X��v�U��uc-p���'4>�5�o�{����lm�&��A����d]��t���A)!x��]�e×X�3�Ȩc>w���2���4YSD>�+k�.y������]�{,u���!YF��B�P���f�Z쳒�d7�2�S�An�p�_��n�}u}u�0�ac�"]����8�v$����|�7|6��
��N�h���v0u�:֧1+ZB�uٔ��|$��%;wWv�fLB^�#,�4��mC�;M�7$�hpQt�N]��+�Z��s�usv�F��)d���?�	����{r��wCfi|�ڧ �{Gm�*^�ʗS��#R�-��=�R`�aK�-��G(*t�s�n�8^lkc�XEY����L�sCt �"]�m^W�,$<;E�Nm ������J�o;EJ��P��*G0�,	�Z[]}:��У]�w]�9>&��N��$�JlF�<d��{��P3�um��q�I�փ�)c��WS˟te��&8��,��U��v�)�(e�j�Q�q�{7F�&������f]�-��� ��2�8�7��ڜꏬ��A�[/%-�Ǻ�bY3�a�0�)_qV�:`Wa�=�k,�KX�\�Kt����;6S�6��_膬�Y�Z<��ܹZ�2N�=�Cwc�mc��ˎ�t'E&��������։��j3�|!�����j؊�33E[��կ._�f���� b��%��1���`�Qg�=�K�_E[��cw�oF��NuJ|��%iy��	tb����Ǯ�T48��t���w���֛�Y0��=U׳�\+4��r���!
Z�^����TM>�r�<!\N�5r8�}n��*����ǪUȾ���ҭq�{B��th���ʳ�sC�JȲ:͙PiM���4��*u����tBp��Xm�H~Z��B!Q�1����wU_|�^�Xל��<U�����C�n7�λ�:eJ�[tUq�*�5���Lu�T�H���1�쥵i�ֶ�z2~qG���h�wS.c��r%�r9�l*���QJw[�144O�nx�LV��9?�dgC�U[Z�r�?L��	���N�1����j"�*�"�5R��,�5�72  D#�����]���(2���6�i`�h�L�wTb��;wK�5����i���:^Vv���*\Y���Y�C�)i�}UT��q����]�5W����?|xd~�?8�@��qکI:g��~��hQC�%�1̽�[��[ZܳЈݫ�^u-�����;Y5����h��/5ߟs�����@H��E�${�}��ڈ� [��Ʒ���%r�pw'\I��t���^�㬵�M�hlJ����5Y2����m���>��'�
:b�&����c7������S���������m�h;���m����������Y�({��[��]yS��!��}�۽o��;����4r�$�ZB���!��()E4[�꾤u������Φ�D�J*q�\�!m��1��Y"���nu���A�Π��]Im�@u��.wD;.�p��a�$MYYQUU��q:���s��,{�b2)Y`���F�^�~������_��ZJgr�䮶��̗��z���g��Z�̜����V���x�2��5�X�"�ƕT(�]#X�#���Q6�	�܀�ŷI���'A��>��d�����9���=�Kswn�zq��e8x��-��v�R=�}�ִ�wJʷ飙;�p�ڸС+Y����}�|����|��^����	7�-@����ʵ����|�V@�F��jؓ����9�q��q:N�T�b�!���X���`##��;����tLq�~���~��w��VN����q��f���}]T��}ꬶg�N����f�c��^sw��/�߻�N`׷�O΅�V�3��˽��X��w.A0��0I��{�ｷ��5�������f�-�ʪ"�)-�J��f���4��E���]s��b��+�Ը�<|i A>��y%iS1Ĕq�⑶�nHC�1I@��5U�c�����h`�7B�@pY"L*���ؑ�KA�|���{�0ŹgTk�NM�z�.,�3u�Y0c6*�l2���]�]>5��n]�1Mx�r:�B���r��
2RNo$��n��ݘE�L7UW`F�d���qF��at]�y�z=�d;�s�1g~�]�|���xo��>�|�r��}c�gً�S$�|Ž6��k:3ａ��WW���(#;�n��#eSX����;����ٛ��\��.��r�z����T����Uw�C�:�7�\�͟��kŅ�Κ�}9^�mz{���Q�R�R�,Q��1��G���=�Q�;�>�Ug��^ԣ�^�2����R���p{��W%T<�v'-rJ�;ql���9O1u�wt�^c�'�ծ%�L�KW��9��I��\{�AL�{�;�%G��|2��FK�^���o�߼�~���s ����"� ��Ru����"�E�M3PD����u�y9����8װ���cc$`�,YtP�ATb" ��Q�ܡchSR+���7�|�F�dz9�-ֲ�,��Tx�N�V˹���[$�uA�%��T�-�q��}����U�8��Hh 8�S���d�kf*=��kU�؅Niu<��*ZoUK�3N�y��׹�P�2�d������	�s�e��m��)��ڰ�S���^�	9W�^��K�%���*���{ɸx�[/��W��ELn�_�ܻg�\��8��e�yEo0خMG��LU�b��')�?9���;β�-�v��T$:0I���l'��ٳ�}�L�fu睮�hW6tg]{������w���U[�����i*�A���+�z3�ï���;�9����w_��z�HW��L ��:�j!�oćE���@�,�/p�%v�e^��5*�2����
�<�z�gG�=Σ�5����z�;��{���g�"�	���X+"0`��a@���%+0Z����4�7�v��w�G�F>�����b���[�����=>�|�7_]��Z��5�S�c��׫=+پ�y���t����!�u>�^a�[(�J�R"���s;l#+7'L8Fb4<(�"ͪ3ksq�ԣ����I���L��9^���h��5q�����V.�Q^s��g�����6�VV��~�����V�B�����ٹ�b��j�������ҧ�
�p^���v���ӧ1�u�P��[헗WQ
���۬�S���8��M�}&#DFWd'���p{��������bȅϷ]��E0Ӆ%����N�Q��TL/���{ɑ/�z��W�}��S/�@�@ˎ�lO������\��^�j<���宐��(�u\dov���ܪ[ʽ�
s�zG���Z(��Z<���V{ǳ=��\7~9�vf$�S�;��Ћc����$�P��z��_����8<�b���Q����e����*0�D���~ᏹZӬ<��y�܏>��<���X�7�^�����Y���W/��c˺]��_�>＆i	�@k-�a��ZS[�}5�u�5����)z�2C,�'q ���ΗXN�kxŸ�FToJGx���a��4\�v2��8R=�_G�d�����~�e��w���j�i�c��E��fNCPM|��C�����B����=T��C�B���&&&���������D )S;�:+*������綶b�@QFHb��@�2��v�j����rN���u>�E*�lu�_���5;ѯ$雉���~�s��̏<�yֶ��'֔Fx{т�1?}���Vy�I}q���w���'�,dě�q�!���w�o��y[����dkS߷a�O~R9ʯʵUx������G��(`����+b���
�Vcr��Q��fQX#���=ϵ���v�!H����Z<�qJ�z�{c�n�.ȵ5�Sv�㽫v��-UN�NAAh��}��w�ϓ�N�!R�����X�־N��~�����pR���O���Dγ�e�R{�H�)�L�ʠ�4�G�������Ͻ�2�}EQ�$E��bB\�&JP�_�R8 &Q�v�H] �F��+���&�\pu�5��	l�]�A㙁r1D�c)+� O���&bP�7 �s(�7r�8��Nse��޲�l\a����hA,P�cu�$J4��E*��5K��]�L��i6�$�B�)�w����I@C�6�I_��>���F�wt�ʫfuɼ�q�k���{��g�O����V���eq5�=_{��G�f߹ѱ��SX�Wg��Z��w^��H��=��f�u�W�^�jg�뵜��%T����J���a���n�&"�ng�˿e��͙"�RcӒ�yz=/��a\s����13R$�F�9V��i޺�Mg^�j�uMo_��[y���w�=���c��j"�b,H�T@��E.��E@�N4�t�y{>�$��+��7|̉��޴���d_���z����bJ:w�)�=�j�1��<~��s�sTy�8r�x�R-M����+4��C�S���$Z��N�~���^_��\�jvn�_z��?q�=��f����$��7�O-�>9�t���1q��am�����eD?�d�hSy�6�	<�p���:�7�:[`O��NH��9��2mj�󋡶�X��D�mek`%�nW`�$:u�6�,��T���ź{����/�w�՛^v��N슷�>א��{����%2g~�~���z$��z����G��a��J�o8���ks~��%��~��^���r��;+��va������gU�޴T�M��//M�^־��g������F�p+��}�ls��XX���M�/W�FMi�ϫ�T�ΐ k�ov�-u�Zۃ77�n��]�n^�oN�.��֫}���\1U�U�х%!L�hY�����1� "���_�r�
��KǅJK�/��]���W���l ��V>15<��v�Tkj�#����~���;��l^o�nb�e�>wUW���P�.�mX�Z'����/��t����G{c�2�m�^���ҫ	��O�՛v���Z�2l�wN���+�V�n^V���w*��! "#DF"#0�C�֒I���9�#����u�Pm�T^�jG/q�/�eJ�K��u��o�B|���Us�s�wm쵴��8gJS;�n��p�Ｆ�\g{�U~_���ȩ��������y�.����W�z;s��mM4�uo���gϫ��}�Y��	��#�n�..*��7<=?n��U�+���
b�^��"LDt�/��UK�����̫���z$�x���+���9�p�{È�R"�'J$&d���n�I��s	7aʞs���y(�;6���NW�s�ky�}��*�����H�0AUEb(
�(�FcPV(� |i{}O�c=lOt��݄;��uh\L����F�B/ѹ�~�*���Wgtk��E뀽��oK��J��kݳ���0���G�����\#���[���wj_o|>���Ѫ�{�?d�KI���ѯ��,��+7��ol��dή(��d�r�B��u.""G�<�	�>~<x>JT��.1�"�X��]�nKUuCM1F#�
�JC{�r�y��ޒ���$"+���P�(�ww9x�}��w7zЧ,ʷ�o�d�hi�6�(��Z��&��.���e�v��*�౜��{�d���*^A�����kYt�<t�N�Ê��j5���x�ٛk���7��ݡTl�H�^�,+&�x� N"L)0�a�������Nuʍ��_S^k*�x��y]YW�z8�ۖ͞�㡾�݌b����@��>���2�** 0b1��F,D�QE�H�b�A�Dg��]s{�~�{�k�}���#"=}�9ʡ�_�vȿs�zNv
�򧖮��L�p��f�_�����G��W;�Q4�ۿ�y�Rv���u���Һ6��~��7>߷ﮃ]����7����W.�������C~������+�|�����$�ﱾ�M�un6tg�=���k1W���'fq�c�" �`�`������������>��*kbu@��O�|�l̳��>
���3��6`�u=�W�3*��P;��/E��#�i�QJh�tA�SO]�P�ՠ�Hb<�5(-9��/�b
�����5ס�U�r#]�|�ҍi�w��/abQ�ؕe��qa��46��J�/�k��]�*�
U�:y�[���i&��NY����fX�^o�}�O$[�ɤ%�{�R�`�eR^�X�l�-���S.�b��N���6��+is
v6^a�)��Lc���!MBcCB�)gm�����ʮ�
Y(F�^�o9WK�c+�f��it=�&�1)J�.�B�T�L�gp�x��)Ĩj���$V,۔ �.Is{����� V���օm���Vӷ�5\:�k�R_1܆Nv'E׷��L���,�5�.4V]�I${�a?wةU���o8��|9�&�V��6�_m�'Y�4�d�Jљ�q�^>����R���z�\�sr��\��ה-��w��J���hd�Ct�<�(d�f�	��J�M��|swLl�ۨ�u��\iL<QK;�"#5+����D��C��ڗ���-�yv�t� e췩�q3B1�H<�dUcn�`��`i��%hab�lb 2���E*��hC[Q���8�]�z^���:��E��B���o:6Y��NN]dܿ�����ټj�
<L�e��N>4�,q�Ԉ��m�$mģ�F����-��>�I��!�A2$�L�Kj)<Q�BRRI!)F�I$�I$�6ܒ8�I��i�#FO@�)�F��0�	�&�d&a	[��!�bI�d��"�?B���L�b��U�Y�DNa�5��U��ٱ`�;f��Կ��>fD�ѷI�����j�2�.#���^�~�m&��8�ۏq
H3/yf��ɽWdK�Ps܌�������q�h*�J��V;Vm�fR����^��E
��x�d���Ù5�Bc�H�/N�����7�鐰��s�M��wˆ�;�%f��T�C�MTywr�
GzV*R-��#,C��9�;U�Mռ����s3���S�:|n��B����u^7E�7�D�2꽩[�wr.iA����2bj��y}�E:;HVr��<�+�:kW�D^ѿx�J�TZ�y�]�YM�E���i `}�Lǒ� H�1[i�5��U]
8�ۂn\��;i,E)|-��Ά�:"�vކG��e<�c�8�x㹧/�Lӂ��`Z��L�Ih�7�e���e�vok�ˆ��#5d���pV|���^� 0��X�7�Q���.=�iq=}�㶭GYC.� p޼���݌��)ݰ�7G	4�i��[!pY!V�����}kmf�き�[K�&7|��N ����u��aCI諯i. _.Ŋ���-I�;��Ӯא5��J��7j�9Pr�Aѯ�f���1k��vM����Vrz`r��ciX����DAl�b�ִFY�y�[��Zf=�y�*�ęBkd����6��vMW�QPA�W�(��d8�Ɓ�����	��p��*��O��T�d�֑J�+��ݘ�2����>�HM��ۅIݨ=U]�A	Q�,�XAR�b�=���G�ti�!q�T0�Ta�����q� H"�BF�h�Tjx��^,��v�83���Zxf9IP�i!L�T��}:���� XƷgM:�XR���o����(n2ɲ�K�H�Ŗ��P��صI!JZ��p��|�@	7i�ܚI�F�q�v�'(�r��XP�1��U*�ev�H�иШ���A�D@�Y��6�<N������r�Y��^N:�כ޾�\��;sј�Dvz����RO�_cjj�r�w5�k���@��Z��ƽF��c�g��Nr���yyk_Y!����`�]o�[�՞v��g�؈Ȩ3l��3���_�������DD��ۓ  #�E�:�zOZ��W�Ix��I��l֒zg����1�SZ�޵��������X�߉��k�^k��1�+7i^S��_�+����X�9O���p� �_�/�y��>YQ�Soӧ������:�G+�w��<�Q8)ojT�]{
7ן�~����/�A����<�,�[�]D�ى�}�h}N{�h��
��տ��M�e���rc�yty����d�>���S�`W�n��.�n�o���_��|�`m�ϐ4�	�'q��He,�L�rۼ�˶Ɵ2�R��!��#\e�m�&���]7;NLX�S-mٌ%*��rsr���w?N��7rI:*I�kϝ��}�c�}�e|�}����$]x<�������41 |�c�6�t\/m��r�6YP���fO���{�"H�}ҹ.��_{�T~�Y���V���J��R��Z��*+_;���w�����,ꠈ��� } }�	���~��[�<�V��Wb]�O���k�rgT�i��e}���Y������}z�����Hn�y/��G��5�+�����Z7�-�4[�)�W\�"0H,�U�_���9�;&C]6RJ�ٛ���-D���Mk�!�gf7����]���'{���ܯ|J�y��o���\�3��1n����=�I��y����<0�s���է6�>�*��O�pmӍ�}Jn_j�;�{���|Hw[׳�.b`�p�͞�\���T���}I�C~��]�:ɤ2�h!�kC�a�9B�tO��}ً��<9�Ѐ;��������������ӫ�/�ςU��8����U�ˬ��`�������Ɗ���[�����k�]쫍�}n�xҏNUt�.o��|����u[�{������C�WN{יA��Q�JVԔD����_�kn������ޮ�B&P�"��u]s��ߗ��ڕ���z� ~���=�����-�����lt����7JF4S��ܐ	�k�@��k�F�ŌV���]1�m�Lv�ö��6��yN�p�B����|�ѳ���~'�<n����ߞpjZTВ�J����I���n'��磗v�&y2S�r�4W�T���㣡�+����W(�(���}��$��A� �0f��w�����R;�/�����|���շ(��P�z��F�q���}0�����g�U��w��<�Dv���k�љ�B�ٸ�`�t�
��u����3�ϸ����1;�<�v��-�z��&YX�u�+zs��w;1!�Y�Kf�
�G��lH�
;⺤JE�t�k˾��i�WjTw�J!�$��u���zΔ݇�u)3�Я��"�����\���ϧ��ي����H�X�o����� ��I���7�۟���$�S<#̬nk>��g�!z�w�.���"�*$Y"m��;�`E��|�YP���ˠ@-Zy*1�B�ۂ0���B�����(�b%��dF*d�Muu,W���u�u�d�E����������w2,xt�_w����Ύ�J���U>�3�^7h�o�f��(+�W�ݙ5���d�{��}�ٮ��3���� �T x�M,7Wf�f�l�j���������y]cDq$[T�e㟔G�d�ʃSC�c��8hQ�0T�����+��� T ���37��2�]�P �[N��ۼ6���^Ħn���Wa�9Lv6ǂJ[�vR�ַQ�;���-����y���"�f�����A���[6�j��������R��(���\^�U~K`y,O�0�yƫ��V�խާ<!��|68�Te$�e��q�$p�T6S��I>��+��&�7Z;R4h
i �iL�u�N²��h�S�{<�XuS�Q�n�v�n�$�]Y��&�ҵ��6���-�.��(�C5	�yR��)͡PM��QGE�f�E�LI1UQ6n�Zþ��	,Ud��qD�IW���0,�R�V�J�7s!�O��Ȼ����g5�X�Y"$�'jS�����J����?}��Ӹ�ثMf��8DA�����KE���ӂ��ޙ���󛽞�'�Qϵ_{_jBG��}�	]+�7����9�M ��w���vS�I���y�u��ҟ�G�G=��%EH�FOU2ً�n��<9L��H�虖2vj�o�vm�b[�}�����w��`�͵���EW�r�c\�$3ۏP��^��{�xG��ښ���"R�������|<�y�*!�Y 4|:T��$�~�+\2T��Ӛ�(����!n����& �8�X��w_RF�xj�;/ݺ�'];���;��o����Y��~��t9�_�-Y-D�J ��ϼ�{&�h|F\UTES@}��u0+\��6�|�:��>�7W��>�Bg�y3��N�=���
8P�?a��;"CߚfoﴍD`�Fj�m��~b�xaP-$
dR,��)&�����F(*�b��D$�O���le����.��,���	QEX�$��=ln����d�`
� �A�uk�
�T��3j���\�A:�i)�t�I���y�63���������=����a$:,�������s�c(?���CY���]ѵ�����n/`�� Fٝ��jO��{]ƊDi�S"Y�?��Շ<z�}�ׇ�E�^��չp��~9sإa�7��ri y{&,f�� �S��T���t���f�f��4��ץd�:H�%� `�����w�'��F��,y��*`����$_WvM�|͎i��w-{��7�?!����@:ie�G�d�ٵ���ɍ�%͊$��qwM/2��1J�Tc.}����m�Q�P��(2�҆��t�e��_${�M{+��ꮘ���{ݽ4�@K�*}��~�>���/°80r8J-�������{���\��=�X� `ޚ�7�6�P���2b=���H�ޤvc�O�hP7u�G.̵�q��@��ⴲZ(J�>�ݭѷ9�}!hCMk/j���YE�U�ᡛݗ*$�)�j��H�,H��Fj�]g9��+*���ȰDc�������������*�+�o��7޸�i����v����e٨��Ђ'^6�WZ�93��6�vވ����f\��1,�c�C��U��5?e�3��+�D�P3x���g�����RL�C֮��1H�ʙ��+�L�T߶�f=Yמ�U�=H�F4Y�+x}l��7�!%��o?� ��b�L^�����m�-��x5e�6����]gmD&�.��Uu-�����!�����M�1� ׃�+�.�]PW�(쎽}�=uv��B����>�j��3�ӓT�eK�
z�|7�<D��A�	��'�BY�=Cjh
�j�� ܦ�7���cV�͵@��2�B�FC�D�f/\ݖ&�����@�W�Kf�Z.njg��axՠ!oX���7B�LX��UP��&�sdMY��T@��j�{ݶ�=���W=޺B�т�;���g�5U�0�m<��w�QQ��q���TZ���P�{v#.�V$<����o>�u���Փ̒),���5<51l�]=R8F�`�bu|%!�m�f����)
M�W���g���>�>��Dx3� ~��wh
RW,e�N�;��D3oMDI�(m�J=ׇ-[��bNQJ��|�G�E}w3�(e};l���)��w�3���F���#��l��P����K���f\0m�/o
��k~'�k�53��3��5��$(����T6v��6\�F�5W`B�2Β��[���K��Z��;q_���]U��e #j|�g[�;w)�\�]�rs#���oz��g��'���dy��5 �7��}�|K���ܘow/;�)y �>n�Z�N6p���BK����
u�����W�F�-v
��6��D�B3�����[S,���{�YxU�����Fp����ҭ:l���ې�3����R�eM}{g�?�����~�H�:s���~�9u^��zts��z]�pﭿ���id!I7ڰ�Q��d�����"1�'�-�X�a��t᧿Vo�Z���9� �Q*1wϱ0
�u�[�ï��bp�<�f�ƕ��d��Й<�{��_}>���G�G	`�h�g�S4�kZ^w��^+vW	�d�%  .��K��F��A�$�6#%y�m��NB�F.�z��U�FeHT5X�GT&(-��ys3�X��hk���g��Xy���[�{��޴��X��̷��^���n:����e���X���Nr�^���j�7�b�K`�D!-AK�@�V{U>����]8���W���p|;�t�$ �oJQ�����{�
����>���sQo�A��z��<o��.O2o��hw�u+�����S.���<`���w��Z�Y���ܹTu5G�}Thg�9�;NN���U�u�:|޺|�UUW�u�7��4Ou���Dy̯I�;�X�]����r7JF�t>�w;׎˘n����^\X��=>c���W��N*����5��(#�b�<*C�b���ӸW��/	o{�y���-R�=zk�^������}=�B�rC/�����L~~��=<�{o��1���C�Ƒ7�ttGu�F�W�}�c�od�_ e�:j���9ZKP(��P�����4���v�_p����LM޸d�SF9���kU���Z���2��p������?�O�Qz$eZ�3���r�=��+|9XY���ߢ�}u��x0���:���5TO�Aa�|D>w|�O^����,�U�X D#��y<i�껍��4ƹ�{s��2��F��+t}}W���g0��X0����ٺ�j��0ɮw���캒:��:��F�J�7�5{꛼�iU­>��D�]��$�G�8hŷX�G3�埴�L�N>nי�Nz�uZ�ﮟ/;st@�$T$���lkw�l9N��12��;F¥��i�^ڰw�_O����,+>��AH�{t�lv }
Kb
��κ'�ѡaЂZ��Α/!d�y#{W��2E��q�`�]O]��픣O���h�ˁ��"3vP<�7�aN*�Y@�T����� ooɢG�t,�]*jh�3*�bf4h�^ C���3!����o�k��}�f�yDc"""�b�8���*���w����Ϲ�s�_�yE`��&ϪP�#�����2���xwz@���������z��]����\�A.9�Lo�P����yݲ/��b��Mi�hZ����#�㗶C�ѻ쎻���������$kUdmD�ˑ	��G=R!��=R ��^?e�/-���ͷ���ڗ�1�@a�x�0����Nmbw�Đ�vۓ[M�b&sͳW�gR�}�U���S\+tX;}�-U��3�Rp?"�N����[��ϯۚ�ÁD�M�W��]lV�(���^_V�D\(��c	R��}eɆU�iǜB�S��BE�v��v�/��qS�5��{}���k3�]�(�8�o�N���%djY��6)�h~އ$զ�����,�c5�6�\����䦹h�
q~Pm���-Ɲ�l�.��ٳ+!ŇQ�K2�ɏ�W�p)�a�)E@\4�l#��]�A�{gccl-��L+�Y� a4����H
�ue[6.l�I�S���xԊʪ4ruv�t���L����i=J��������1�/h�`��Y��E���o���b6�r|n�6��1Nw����ըR{���x��:>�WwM����e>�<����v�FBo��v�*(;B�T䣏Hծ^��9��U��[���sǝ�7mvr�49�e��0������z��D��ۙwx��zA9#n���.�ܢ4J�À�w���������t1;��D澈e���uS@lVɔ�vk׶�,]2�)�|	��O���GIJ�]}��^z9�������`/.��Ml�s},����T����졸�>���U3�:E���łX��<�kF�v>M�J�t��D|;/��V��:cX�+r��m n�K�'j���t\�lo�[F[��n�[�K��])��`��~��t�Y��	K�����S���f6{��J�@��f��^�b�I������r��̙��7�]�Շ)X�N��xT.�Uv��D��3��[n��ҭ�qڒmB�]ݱZt;�b�k���+K�7�^L��P̮��j��ׇz�U;�5}���jJ[oӶS,<�'s�NQ�ً���h�ǀ��-��M�zРܝV�%�"]�EΥ9!ͬ��k(r�F���^;��5ܰ�`�7p뎬L;���k[��;�H/n�#������H5����He�;����p��kyP�{�]x�]��[�Gs��<�z^<52Gm�[fq�^a]�Y���|�.YERu��[²����Z�sL`nm�d����u�
�n�+�%gB�޸0��α`>�]#ۙ�}i��Yk��7&�y&jY�v�� Y}�(a����c�]��k�5�]G&=?�i�si�!��������p��&�̷�1\ pu�c�gߦ�ه�e��us��/��������=�&LvСKR�D�s�R�`���� ��g�U�2�w�'��Mc�X	<��������;�c/�X�c���um�hm�˥�����85��1�{	`Ϗ������m�~獂JZ����M�͐BD'PG��r��p4י�{�_����?���z�^@��d��Wp�C�f�?Vp�x��wӃW$���Yw	���i.M|gS����t�Q7Q�\5�޹Z5S/�4kծQ��}��;�.�Sw�o�~��]��A@b��*�E1g�|�;�����D��\�������8�R���<zrT7Ƨ%#�ܚĤ�w�G�eO�[0�J�~��#��za�U�Cx��
#�2�����Q�6� P��g�B^��k9������/lw����("��~ ��^����ܽi 9H#��"j�=��!]�ݷ��xJ6�\�#����=t�ƭ}(�{C�j��z�Egh�͸:{k7R\��5*p@N|��"j2�΍�tE��o��{+�(+{8�*<�q��R7�0�����ǎz�<�w�������۳�]��B��T?}Gu6@��b7���Wa�ƒ,��Cc�����W:t�/���~ʳr��TS����Y[Rě^���ª�`���3�>X��x�����=��&a�rL��=J����W��� ��΋�ڷǸ�(5ϼBP_�c-neoa�W�,:%�ի�'r��q������ּg�-dP�$Dd�s>�E�������D}̗1*�I������>Ǫ��=&]>����?y�$�^���ubN�]J=o���5�Dv6�(S�ꮺ���LH����`�:���J�ϼ7�-tj#GZ�J�#Sb����ٜ-:��eeUhjS���*��VO�ҟ�5&�,���ݺ�3f(pO��s�d����>�8(�u�5����q�a��uyr'��ch{OؼO�`X(wL}K_V%��K����n�Q1 +EV��ډ5E��p�#�!�8�h��n��ڻf+2�Y�I�r�}�����4�I�\J��ӡ�m�h�W�a�9�ke`�n�h��'Zld��(�!��� ����m���Z�k)�	L��R����iJe�MF�>Q�Bi6d� ].���1C[jB#���� :g�].�H���6�\��� �!�o�}^x��P�ʲ�� w��t	c�se9Td��>���~A��ttU��nzd
�$��=7��6��N���>) 	{�}�Q�OCK����N���e[�� Jl��z���6|>_R�8��ʝ� `��ޘ;2��_E����DV�LY�w,�K��؁�l�]�|��A��`��
EEE$W噾��B�n�0��"G�w6�p�]u�,̕�0�Q(1�%3��q���J��1#-O��\�T�����%�E3��E>��`���v�s������y���k��,��J�^�K{7Ҡ7�y�1\�2����C( �Pt1��`�����[ z��^6.���>v{�엞K�d�oKz���V<�e}�b�Q��	\jØ��������h�!��5�u�]�Ŋ*�Xv�EAA�	�(TAA�S�EA4�m��� �qZMbq-t�]�u�5ݼ�3��{�m'j���� �yT��E�(�ڨňmp��&c��3p�U�9ܾM��,�R�9�8�H�6����t����ʱ%i����X�������3�)lk$=u[�2��k*�|��.�/j��䛠����N����%E��,�Lvm�n��<{]iy�~����I}���p��nyV��`2ǽ&XE+�ݮ슋m���s��Z5��1�mfL�1���tBmC�;��)c���Mkވ_�r��M�ŏ#�;�Ge_ou�� �
> i�H~?��4yN���|0QH#`�(N�TX�����s�҉dX�Ƶ�{��{���$���)�!��z�������"����3��ڋ��HQ"W���p����9��U��).&���F�dg�H?J�5������ٶ6L���HܽJݺƾ_&�{0�paN�Ѫ{���BB��/A��~�[����Ǧ���M�{}���x�1�R��*f�,G"�Nz��<Xx
s ��5��w!��p۾��^]Ԛd�h
$Q$hTy:�e)�>�Hfr g/���m�����I�jM�=�P���z�����{���#��{�cGS7I��V�xq +^�>�Ȳ��9:3�7�e���M�ُ/8�ɑ��NU���/$L�B�.x��{u������J���F���=y��PY4�牔2xk�>e�6OT��e��:�H��tZ��ן�;#�<e��Z��=���J���@`�ِ3�t>1aߪ@�d�O*c��ʾ,�V�g�[=�D����yo���U�dp>SP���\�d�t���x��� �,b2"1�F(��:޻Us"b� ��"=�|�(���G���)���߲k;���L ֲ�&����i��Pߧ�����qs��F�ˁ�[���TJ���.��-O�	�`����mՊ����m�Uʥ��ڱHl8.a^x��m���f+ێ�=3(�YRM�}a�H�!*U7k�K~���/D�_�%m�v�x�>�4i�����>Ub�޽���֔�����{��g^ca�Õu�ܫ���!���Og|�QC����5�=bR���r���]�h1�I)�󜺎��[��^��|pS�}ݩ��� )!����B#�TC;�*蚭���W�
C�~����c���[��Q��Ƴ��´�%�u2m��Q�4F�L�4�gK�r�÷��L������{��D���w��	�1CE������2'�4Gxd����~�����3���mm!��u]�d��Fj�C_f8ͺ �����.�eR�'@�ךG Rx��T+5�w�p@3���FuI�U��k�s��YJ��M��(g[A@D�ws_k�5W�1U�m���=x�9���j@����e'@8�����mG�/RwK'����I־T�o}P���~����w��(	U|= {�>�a�E�4.���7YW�zg'g�Q�~�~^2�B�P*�@bɍ�� �.4#Bǲ��/δT�(|+{v��c��PEs9E�B1g<�����7�������(����[q����u�x
"P�Q�^���p�����HD��H\�u�:jm	�1�/b�Yq<N����j�ܝ1�fUxg8��c�c���q ��q�V��:������wz�G��OzΑ�B�i4�-���E��J6؄���-��mnsdV�s����:�������J5�^uumd��8N�J�d�f�ϓc��ˀ9�ax U�r�D�B��Zc�,�0�*�*>Β����.M\�%-+� h�]�J�"�jό��a���D��u\����E[!���!�CZU�.\���LI��=_z��r��P��h檯1���ѱ�3���߳2��+���2��(|��䎏�v���������F��,V.��� ��d���c9�\����]��`$O0�hUU&P)�40U�j\#��ޱ�sY;��+Y�D$�G�c� ��̱?R$w��o�0���=3JO�ߵ���|9��da����^
TȐ)�*@y���1�z^[d���_lv��t�̻ρKt��Q%�D�{(K��)EJ7g��[\;���� A o�d ��A��"������>��r(;5�g�x?�\�>��u��!��k:��z�{�J����sm�:��.5��D"�@�.�s�>=]�ɠa"�1� J8&'<�	��0���~� t1-��uC����Д���1����Z�ڞ�P��k;����
�c+R�9w��_���o<�������Ci� 7D�}��*X�$s����(ά���� i��9u�#:s7�\�z����=�/
��ۿ-��hA��W��6��Z�%L��6w&�qL����(k�R���٩���������G�����RKl���g�V��v��ȟ+�OCJ�5�^��珝k|�N|1Ĉ�Qn��AAV)�L��>��} @�]]�ʶ��pL��Sh-�xF��B�<���u�wTW����� ����ǖR�W�+��<�������KgDz؞� '-�B���>����_yw��'�a�Yr+�j{j� c�{�W�@i�w�\j]_Cv�oo��ɾ��{���|`��t>��z��>˨�T�3��)���ey	�N�"��+~�(jBH�+�W��-!��N�,�Z�P=��j  ��Z�~_o�g)P���U��|��޿V��ąN+�0�v#!'��b�V�o|�ԇ�Ԅa���^3�V�r�<�!�N@L��E�+���]\!�ؕ�{;�^�)Y�Q5 �VRLS���1;Ε:�cտa�m��^��HI�ѿ�M�wR�}�gޓ`I1|�S�Vr��#́#y�mn��7i7�+���	E ����h3;R���j�6��뵖�S���d�v_o	'���Õ��߸�#����A��q)*���N�#>��^3����Dbv�v�Q��Dy�����*�:�u���v��ۣNZ�!Ёk���_0~?b��������\�d~#�O1�FhΟ:7���Wݜ���1�6���_�+~/�F�<m:��3,�ZGQnj��1X5����^jML���D��s�YT�ک�xS&O=[l`���}!������jN������P)4�Z\g��1`��Ah:ľ�ZC�{q���(9�����w��|�:���T�� d)��W�n�#Ԟγx7��z����q֠a���`�	�
�E��s�o<־=�T�wk����X��~�鋼�!W�t�C��$�+	��������s�u�\��y}Q
7e�2D���H�阿ڟF�-Z��-T՛�fh���r.�
fq��dץ��Z���k�^`j�53��=Qsm���"ݻ��t��f�-?�R�~5�!�K�4��0�Y�-�ss����.�O��F,UF+�9 �J�H���$��$�H�ӧl�N����9kkK
̶�9�P�� �m�w�C���wlí��\o��:EӨ��1oO�*������~6�Z��8DV)�̸�+��P��� �o���}O1a��?�.'櫂�MeA�!���=6$:=)/��!�ѭ�7��ڲ6"&%BB�
IF�Պ�[��%�6L��D�q�V�ג�P`�Y�f�)��d�z��� 0,��֔�����r5��g�7w!��gA�{a��^T��O�H��ya�͐b��ə2���!�za��X�)��M��	�#�|��ۺ5/>k�H_��������
�u�
���;��f�/X>|�6�+x}Uۻ<5;M�� ��f���9Ϙ��鲼��~%�^?�O��;�a�]yu�l��(�j%~�]��}5%��$��!ɉ��5y����� �}V�j��,p��e\Ɓ��%�W��K����$$����I������aBBE�B��$�00	'���3��$"�I$ ��I$$��c?�=!$�$?�@� ���!$$�_ԒBI??�������$$��s�������l�h��$$a$�I�@$������$$��s'��?���I�'�~�߿�$$��g��I	!$�����O��$���M��.I	!$��7f�y��L$���OΒBHI'�>����$$���$$��{�?^�?����$���K�~h?o���!$$��*�HI	$�����e5��\�*%� ?�s2}p!���ҽ�tT�M���ْ�[imm%
�D�]��6���m�%�PA�T�4�%R�%m�JѡB��Q���ųӠA�|  >�(���TP
AT�����%D@�P��(��!"DQT*AUB�U�T�H�� H��IE"�P�TQRU$���ͧ��/v�jx����ݶ�Ǟ�v�-���5<��|UB����Փ_}�__n�[o-�mV�ܺ�m�vt��uOj�nz*�yސ�rݬ�������Qcr�yuk�ݷϻ��}�[��!A��|[[]���&��>��K�K޸褋�Gz�Ē(��yPR��IEv�<�(Q�n�S�B�z�UE3�qUђ�jT;;�����I*��$�(EP|r
$�2{�:I#�X��7$�J;��{��H�U�����ID�븾��J(�1���$��I(����4QE+���'���(�8��h^�R^�����+:*>�w���s��IE;���T�(�ݜ�cJ�/,��{:*��ΡEZ.X��(sސ�]�I#s�^��Q�tU������O���s�
(x}J��δ���
�RJ)@��T@$�)��(�N�9|F�H�Џ�D�y��(����(�n*Q������袇�c��>��Y"��ZNZB�$y��T��IIX�y�kB��㢟��]gF�gD�|�Q"O}�>��QH�}�y�J#㢒�1�ۡD��܊��E-QJ/�O���ݷ)�� /z�k����$�-rژ{�N�zۗm��vW���C��J�*���%E*�T� 	��UK�����w�=��}�t��z��U���w�ꅶ��w���k�x���m��w>w9�;���T��>��V�qu{���:�ܮ���o�m�o��_U�K����Ҿ�Zؒ���xܫ��>�s���j�}HW;�V�r����í������c��^Z�b�����R�z�T���s����\��g�<��nѵ7��ս�9���\��ݔv�$P��/ҨR�R�AB���(S�|��U����vV���m{�k}��}���]����k,���� S����o{r��\���=�ogZ�w�;�/��O}wO}7eE�}P*�/��:w|���,��^^^��!]l��%Z�ͷ�{z;��s�����m���$P��}�9|��e{ﻣ���s��>�����<l)J�<���*���)T�v�|�U���}�����}�t��A�ϰ�Em� 5O�%J�  ���R�  4O�Ԫ� ��R�b�� �4�*D�R�~�CC���)Q��@��?����.�ppj�z9�B�2D3���μ��[� ps��@x����s�� � �'N����N������N������'I���s�s������~���� o��
��s��A��/0ɷm���UJq�n�5R�6��k^d���,ӂ�	�f��Քb�=�fL�wOI�sl]�4��Q�P�6h*��(�4��R�1'�	�z�pU�of����Z�����7�Ѷ7!W";��M�)Ӱ�|������H�����u㣟
$����y,4. ��nC�����nꨫu*��������{�q���ђ�`	�v4mcא��6,���҃N�m�L/)�A���"T��+4n�,*'f�;D��a=*�0[��;lC�2���B-�������+����"�HGWǍb�y��P��9v�奘�
�"�����T�ѷWB��9�Wi�s6�#Y3�N'X���ػ��.L֭�hk�EH��W��d��Y�g���
�ӹ�iq�`��t�Xθ�s��191��p�X��U���K�.����Sa��J1��]��	����H.��q����m�y.�;�6�H��Y2+T��P�j�-2�`�^φ9�P���An=��f�USfaw�7GfX�2�ti6r�ڶ��(N��=ʋQ���h'���P�Y�\P��Im�wCds6����*f]�giMʻ���n�j����%�H����U��i�;�����C勋I��J� ᫑9���ϓR���
Xp^�@�u|W��S��H����}��pm��Y\��w+����e�f.t):�K�͐³��^ovNop�r��T���2�4�d�>��CoE�}�j����V�Xo������))�ʉ��fe�p��!_G̋N�`!�@��p=��fG���i��+r�Ѓk+f��*P�YY�kvT[Z-�`Z˴�6^����e�Rf���1L2���ͽ�e�"�ȩ<˧��G��d�SkaC2U��+��@V�0i75��2fY̮��q6qӠ)5�AaT6;�5����ژ6c)Ս��z�7�;ܱ*��װ�Z�	B�v����Cl�R`B�����L�z�7\�"�H7�R�!�V���S2�,�{��\L��YmB�9[Q�cv��LVcTɩ��R	2�cu���	��W�%��MAt��b�Y�ʸS!�\��gM�p�0bܚU��={{t�v̙�h=���9�`�� ���l�*fM�w�7R��sSfjsB���Bx�kBS��-�q�ǩ���sZ%x8�]
�޵��d����H�f��pC1�^��c��`H�M�W^e��ͽ�tآ����d�v.Soz�-��j����<�u7�p[�Y�v6�J���<D˷5 �F�V�]hn���슢eCE�at�f��Ε���{r������ux��@� iAOL�[c�[j��4,UYI�7)Խ��v���`=�n`��X�I�P�G�
e
J��|��������NV�@�(֒y��4�wYЛ�Ӄ:�,�+ڡ�J���W���'*�ᶝ]���mˌRp�� ]�/>�4�FK3m�s�[��\8`���x��A˸�J���1[bk!%���u��ċ+Z����p���2�i���i�)^�f��AM�� f�Y|U`��b�/W$��Qښ	l���K��8���tl�)�ɴ����hT�j�b땅�`V�P���/N8�ɛ�qb��5��1pe^U��!RuS�.����@P���X��[Ǚq7�;�^��y�,)��V�lb�Џ6��0xh@�l����sm�kbi:�ͫ��%xnK"ə���e^�V0V�Kզ5i3T��sG'.n��o	�W�V��Z�Z���*Z*T*��v���UX��������q�yW��k����ke�nY;�ە�k�z��k]ec��j��'�n��5e��Ç+ifwTgxS@.�����I�tdU�S�u�v�7&�&�	�Ob��Z��!IѬoD՝hY��F����>:	
�ʎ���_*�(��J��f�X+mfZS`�N���,���dD:ԩk ���R:6[����b2�c��a<��qkIѠ�x0�u����lj�p�$�Vt�rb�eҧ�u��
���e���g� r<p�������f�ݼۍ���ݝȭ7n,˰p�&2���"Lҥ�n�w!b0���~�2�X��ݥ�X�&��ؚ����f�����R˖�[9Fl���\�(�H���"o42��6�r�)&�jd7@����++^1):.�f�n�p�L1l0d�,���-��&�7j>8\������2��I����{f$4�tV�y\E^i�SO�$�n�T�Q5�*]�l�9�t�(��_ڧ_�j%V��s\>�h3#U�Yk�H��Ug��>Yv>ICw�jZj�Bx*�:0�pq�:U7���)�V�k�P�a�vM��*:�5�x�k0�A�4�'a�`T�5�Y]������kڗK
�٧8곸/�:l��{!�!���С(�7̫D�I̖�fGkr�0 �1��uB)͓�z��]�Y4K�:e*'C8��bu�7�Mo]�ɡM���u;��LG�Yz5U9�N����r�	��[��x]2Lzn���-pğk�V� o�uv �����q��y��UXP�i{f��eV���5w�F��7ƒ��A�&��۲�gn�yc
��c�.M��n 6��쓁�&�5���Y��F��Qٸ��32�^�t�w�5��)+��ޫ
a�2=�n&���)6om�t���-�/6�T��*��Mb�F�5���4��hf��B�������1BE�&�
4�V�;ICVlФ�{����X�5� �F�I�e�/S��d�LT�B�RH�R�*��su �ݻ��7XX5�;Kp�Uif'�-^^��e����Ƃ�'3A�����4�8qm������L��J�y,�t�v�����,&	ҩ�-��Aܩ�(�D���f�M��ׄ;�mӠ�[em*�E*��+E���4�Uxin|�6�T(���P��HZ�c E!-e�8��Q$��e�k%<��F�9��k��Ecm�4��t�Ra�Lf��A}f�V �L��Z/NLڵ���O��U�T�;�/]+�#�����Y�#GnH,��g35Q�L��.ɈZ����p�k�n��(c(�2�ϳV���h��\`՝��&�SI��ն����-p�8,;8Mjԍ��t��W���e����
������C0h�)e�U*).'VB07b��(�@�a��Yf�IQ�E�	!S/)�m,���Le�3Q�&�N�l��N���6vp`�؜��r�P�R���ci�43���[��ҵ+4,8$iU�rθkkg7��l6a����WF�����
ܱ���m�Ė��P�ti��L]���
9j�"^5�"��)��c&�ŭ�!�w��VQUSd���q���AA�9��v�7KE;�B)�z3S����w���;�t�_wYoje|����h��S��Tlm����R�*Y�4���=K�{m1�e��l��F��yR���b��ɖ���qާ�v�,�Re���;h�6�a�o��B�6�X����pހE��la�f\�{WS�����w#��z��$�XA���|�0+s&�B��M`H�V���k���&������Xv�C����kCYKU1�^Q{�QCE�x�f�k{�L�4;R���"ʧ���d�36����6
�i�ᙬI$%^G2��9Jڊ'ۛ`i4��i1WRʼ��E֑2�A�u�y[mn,�jS�B8y�����4����"��#�o`W(5�D�i7P6�C5�y���TEd�%ɘ���sWٺ/R.�L+U�ʆ�h���HZ����d�ٻj���O����7&�MZ8eD�N1�L�2�fR���UK֑�5���vc&�k�e��:�P�����B�oV���O��\��� Nu�UHKF
��J�6��q��]+!���[1�HA�j�:4.Y/]Y+k���F��LT`1"t*`m��̆8�p�
3mL�Xt��!�0jWT���&��6���f)�m:�|q�=���Z��e�ɥ˴�V�HM�_$o�˱YLf &������n��*n���#��A�o��Z�ܥ��ù�kK���(JC� ;q����@��x��h�0���۽R�cBͽ2��k�8��lr�T/tU�j�R�xi�ns4�L�l@u�ꁕKz��ٖڌY�lX��*� 4������`�%n�"`iY�-���yF!H�2���*�F͛p�#�!���]U�aq▨�ӻ�/d4�ѿ�����ve�m-�#(`���<�Oi�� ���&X�ޔ��TX�ʁ[�r�d��`���Ð��Ǳ��ښ�ac�t����[��VjcNdnP��56�FbT�@���D�
����´qԹA�z��О�b�,��aSl����1�@r�z�J�˰�m�Y�.�^�*k4r�m�*�f�� Ɓ�@^���ԩ�r���A��K�X�`�ز�ob�z�$܂D�a̡{��w��eJ�C�Xun�[v15���m�b;bĚ��-5�]dg-[�tA�T����H�$�ɺB`�iO3U��ݚƴV:h��6ܴ�)�yb�K����5�V�YY��n�0�"*U.5zj�Gj�X���Ŝ���y�*/)Q9�J��q
��Pm6�Zj:�7&͒��e��*�{u�M��0���V/nޚ
��GwF��(�:�nK8�Xt�tb�X�F{�N�O�+����U����ܩ(	d@;�#�N�����i���W�A���d�䭫+���r]3�+D�9iŢ�-��1�4�i���kt�d��K0R�+^泅3e�ط0ַ�96:W*!�b����ʍI�Ǐ���=¬ف؛N�YIv�C��{l@U<���N=���H��nI�
�i�Z5!��7���߀�l�TM AN�Lwch^�6�u0=��cVc�}"����'6�	�:�V*Ӫ�.'<�w���An�aAL�76e6[�KL3d�7��3!�q�����uP���XΜY�,�YbSxnM�����h��a- *%�a��=dK�6�n<�.�_	�*�.s+d��o�w�'sE�7��$1���`��V���.�C(5�:.R(a�RƬ�C���mh�"5��V7�x*č gT�J;f� N]jd:���q⼿pY���%Lp�S���Sn�\�)�fF�R�0�p"9���P�j�hfM(�/��\k:��;F����� 8P������� ⾄Pd��^��@�͎�ˉl1y-h��RЙr=w!ǪJ�-SRfei2}x&S5�T�*^
o
E�eATI8�7�M1Y{T�=U�J\���V��3A�B��6��N7#���h�l��OAKvseУ@�<$@�0hX�BpnҸ�-���E�Ii�ml�t0���mm�j�;�5V6ed�-+մ3p��!�����&�(=(%��ڴ�ǐe^������u�6UUdr��������"�<�` �$f��U�!�tG�`ycU4��=.�PdMQ7R�!��� �^MH��ms0�NT!Y�[B,C)f��N�zs�d5�_P��ɳ�3�Q��;x{��M�;ļo���I�nw��S�[G��(=�B]m�M�6�f�	P��B�&z�OY�+^������x�� :�C��Z]�`����'/tʬ���=��.ב��}���-%v��}��UnP7A�d[�Q����,��?o�V٥��f���UlH�r,�jS��_^�5�L��fUsQ�4�+Շ$u�K5+ H��u9�U��ʗ2�&ʝ�@�+5���V�ݡ�[��֔�lk!������v	��R	w|[z��5ꢭЅ��)l4�Y?�������kpT٣lI(�F�)�f��(\B`P�D��a�C�i�>=��W��V;#�~��\�K�d��KyUEN4)
�%:��`�e�=;6�	��B>$t�Eҍ5�p�����_U�sfk}�8�hh�V��ځ(3��I�Y&�v�pi�Va{�Ī��%E�	{�wdڴh"�e�7nQ�^wW�uښ��uM��,u,p2��{�a�(ӭ�+;�:l�sz��QV:u�}k3V��P@Xʗ�o�I�>IC3n�j�T��1Zԫz�uDf|��뚎�Ц�b�eJU�yA\�iV,K7 <2��VI�
�Uƻ\N�욏�c�L׭��x|�Hx,��q�^�����c:-oM�)W�4�mN֠�X�.(��SO�o$OM�ѩ�̮��X&|�`���f�Տ�����RV������l�6�k|�;WQ;*�om��G4�»F$0�(v����w�H�����Eо�n�]��'i K��T����Z�cu�l[��5�v��KU�M��rZ��s7�����/zk���Aւ�+�F*�WO9kX�#(V,�J3�.B�kg���+��R�U��t(�V���5S��hy�y�ݺ�P(��j�^��i��a�,�lݹ,\n� �J_�]���׍e�{�b��w�)R�UIb��=�A]B�7G�����n��Y\�dcuhi[UXq�C�Mȸo^<N��W)I�i�:���=E�Q�C��MA��w��0�&�sa�V���Imѭ�2�B-jSr���J�(L7v��)^ޓ�*�.��dׂ̬9�m�5�b�e!�Un�@F@TviYy-�s3*�m��îX�#d���[z�T��^Tt�ʽM��8��i؞�l4�t�Ю��I�W�i�Itn�� K2��N�D�t��A1�R˸�k[�1eԳ������i�g@�� T��#Q̷�n�8���i.�0"U�w�X[�^���ƍ�q�sB��ǰ�T�2K���fV+-�{�"Yr`��v�����pAdQ�A�6V�I��r�u=GJ����:i�$�j�]c���,��iV�����_��U*�UE[���NP ح��j���SK�,UU�j�����6�	IejPV�j���n���;5�Yd�܎����p�r��UkpUzU��U�c���~�W�"���^���檦��q�X8� fn�&�u�u��ZU�U��@j꭪�ꪪ���A�o���������UT
��`�U�����ZW������ @*�K�gN�U@UmuL�;=�5r�U@j��]�ԭ c�j���w�̫ĥ8��9��S]HKʁ]\��
k)nJVYPت�\��ڤ�0#5�	 v��z�T������y#�---lԵ,��A�y[�n�mx��.R�$-k������(�k�:�l�Be����r�=�����&���[��ܵ��L�5���#u6�G�*���w:�vn��i�t8�^���3��`]����B$�7Yk.q�<=dUl�Yg��;Z)��@�:Ȋ[$��\�S�S��*A]�+n�qp�!g�\He�P0��k#�;d���df㜜rF�E�������h%!,͊�&اs���k�*���v��r)��Ld,ģx(�ۈ8� �n���n���X:q�������ړ�sn3�m{��κXв�P�۳ ���Q�1)�J�>�9�]��.S<��Ks��+Oi��xە9MÞ������x�aں�=&t洼�������=�����xkF\�n����{�e7n���;]�U���fjp���E���#Ka,�7��Ƙѧ�m�!��vKL(�����J�/�����u�7$�˥�;"��n$���13�t<�Ȫ�kQ;h�݌GZ�;x��W+	��.%R��eG��:Q�݋m��w<y��]��6�,�V|�������޷I�U�W;lZ��[<�]��������e��;G\ѱ��F�b��Ո;l> {N�%y�S���tb�zٮg�Rvd�y�!��{��N��nr&m��]+��G���B��Vr fnqU-���=q.-�L�5���`�:��6;`"[A�.�|��)	6%� �4�
�P"�B��.Sk�.et��M�����it1ƚ��n�������ԋ68Ռ�m�fb�ᆺ&]mӵ#����Vn����k�T�(0�-�v����[���e�M<���܊F��� R�%�2�[hm���� `��mT�y�Ĥ�^�B`�ެ���,v ݎIw&�4�CK��=���pqX�����ȼ詛�]i��ڳn�����䐞�GAǎ'�gt�/#mi�΅��Y\����i画w7O�cin.7%�t+/g^M����Y���1ёq���S<�ǎw���.4��#�I���5r�@�>����3ַ*:���m�L�A��:���8�L�٘�D;9�Ĵ�����5�X�4溸\��9�<oQr67Q�]5���â<)��vy%cl�`z�0�xs��0s��yV����+����mP�7��]����d��uʜ�mV�#�;\�8�;&�I{Y�絵]f��\ �מ<v�ۘ�B9���!�`����2��7PWO[w\���ۡx�8�<�+h�>͠��ᅊو��\��ٚ͋� �SV��S��^ܛ�Um��R������C��wc��3����v�Ba�����:윧nv�%����O7����.l��^ Q��4,��]u�;m7\�cJ@�so�6!>q�2oc;��o	Ҵ���^��8-�=(�R:V)Ջ�nu���N��;���<\�8�nԢ>�u�=Nݒ#��γ���ܻz������Y��1&헠e�X]a4ҡ��Jr���Ut���9��H⛔٭r���O&��O^(�r��yu*������'9Ѷ!`M��e5pd.eڨ�sev��g��\r�S��5��� ���U����y����@w��}��AR����SF��v-�kv;qrñN�N{j]�0��W6��uR6$�ju{\v�ާq�Zy�q�e��\����g����k��5��n�x���1�����SK��@�,t����YJ��q���n�̶2�hB l�m2����Ы�[��W\=#�m��1����S�9�q6�Q� �=+�#=���z+]M^`��I�0��t�m�W������7�
|k�U��=q��7g�Z�m6^�L�ݻ)���K�t�L^ ث*���n���!S��څal)mܮ���M��^�x:	݁v@�.m�8�k�UIۮw\O8�X첌�7g&�ёP��zd�v�i�cS�ں���r;��q%����m���@dmDX�h�"�A� ��T8"﮾��`6�[�c&�U��n�`n;g��Eqn�Э'$qk�g�ah�[O�Iz�ٝ��X�RJ���Bʲ�,5AiP�H�4a�b�M�`�S5���V���g�=�yٹ/O �|��^р�HC��q��ͪ;Tb�1S����q��K`\��E��6�ؕfH�j�!6К[Vck�H4���z���C��lS���8ݓN���}��~��]�0t�=n6Œ3ȯ a��;�`��B���]�=��nöZ웮 ��%��&�:*�U��qv{Q�O��1nA���L�5hǩA\�)=����1�Ie�dxv�l9�������B��.�S����Ө��@k��BD_o<�ų�hͯZ嚌r޹^(Q�ۮ����5��#R"n{��:�yI=s-�4�҇�<��tv�����m.㉖.&-8�9Vvg���'*�B\cH�W���74�À����܃���m)tF��)t��l�j(���آc:��� ���W+�o�o��Y�A�J���r;d�/cZ�s��ϗ��'YK>̗2Y"��{u��x�؛�䒊n0����H;��A�nB�K�JY^�fF%��:�N
˛�8�4�;��K{���4q��6wq�ǘ/f8�vc�%v˵�P�)P�V���d�a-�Ƶ�庄�6du�f6�ڰ�`�e�b�̶Q�p��K�iYbdA�2�rnG]�&�nް�ut����t��ی�o�1���Զ���CXd,7m^�^s��]��C4��֖ۈV
��Ơڔ�#D�j��)�Վ.g�[����M���6�⍨�A�*B�ܭ�R�ԋc����k�6���Y]\kY�>>���p�/3d�a����<����3��<1�M;����V��������Xh5��	��|}���pd�6����|��K[HU�C8��9�lve��h�:�N���p8��79���	�3�6���K9"�T}��m��a�k2!u	�&�I��(��(����GB��b��3��C6�ȸ���f洶��ⴜ�ۗ7F�v�-˚7nG8��6�K��󮤩�[�.7�s]a�I�hd�Qy���k�WK�ai�+i4�Z� ��ܪp�K�sU�oE�:�:�-��@�Z�]��z�@h�]�����e�b�8�]�|��kfu�cokWv��8P�sٞ�����"��l�x�]�V��R{��tf�n�54c�s\6�u���{[�R��4�=�ڊ��4�$,�pKD�[Sg��ţ���Og����2�lwge,JY�-�`a��i,�͵b(=�m�yͩ��٠�&s��|H�c���L���n�a;D.�3Ӌ��r��M�ۑQ�L�]�ђ��j���'=�0t7>z^�8��t��k�'��D�����l�{i�����!煙M
��¦�x�'��=���^w1��|�s�<�ܴ����lD�
��R(jkh)�Jfݹ�&��:�	!,�t��0[C�i���ر�0귣�ڀƸ�sä��AIf"�k�t-�x��i�8s�-,�jF���kr�ef��`��h\Y��"<��e��)�,S����š�#�3�gNxZ��Oe���k-���]KUp�8�2`u�۲�[���s�n7*lYNч���.$u��s��H���
��o;2bg�b�\<��-���e����9ֆ4m" ��[6��\=ta"Ʈ�(l����l\�%�˲b�r���������g�We��X��v��Yc�]�<b�{u�Ϙ����=h��e�S�͌�p�n'�ﳻ�O'���5 �0H[\����&��ڮ#![�t�Pz��^t�SQ�8��,�ͦ�8��vے���W��WE�l4u�4-��aR��9��nx6�H�ew��5�/3�^3g����x���0�2�R�٦��Z�a)	�Eb�h��me!/P���0�5.b��x�X��Nk�}�d�v�4��|Ѯ-�_����$�5׀��qB�°�,](V�R�3���Yx��D�1=��8�� N1.ֹ8�9�7�bd�V�mC�K��ut`�&�Y���V�s�J�Me��c6u��Жi[��#��3�3��������[������j�����5��S:n��k��V�ݯ.����wT���1玛��e��ǜ��㶀&t�`�̱�\�Y��� ɞ	�]�c9�v^է=�m�s�HW�`ꎴ��Bmՙol\�;�W=I���c��CX��HJ��d����I��	]@bR�nqh��<9�g�ϲl\�Y�f-Ѱ���
�n��zq�n��=��擜r:�q� 3�R����G���F�"��k�������{Mӷ�zF�X��>x[�-�Z����H�K�5����=:N��Y�EU�4�<�Μ�줰�a+�b6��7��v�*���h�\�(bT���i�ٺt�k�Ԛ���k�$$�o<�踰r�F+�����%�tza4�e�y�l*����m G��n���<C�9$�nl�S=���Ƹt�V�n�/I`�9��gv�Ka�4T�&��h��3d4�v�Vْnݴ��F�Gb��֝{&8��8�9��y��B�Z�k���ݕ�NPN��4�ہ]��D5��e�Ғ�v,�,l��b�V��ɼm�mPirٍ��Md�*:Ņ#�,65	�33��t#�چBw]j�v��<��t��F��	p��Tr���.g����M��k��n�'t���?�i;�N��$�Ӥ	;�t�?�:I�wwq�;��wt�������cF�b�()�����+dg`�_.��2`�6*4,� R�U��$94tg�&�]�i6�M�5�758�a1�kGo'..�k�J�d��ۘ&(��4�9a��Tmb��a�m,8��6hYbh6YeQ&�������y���ܔ�\���b��,.֪\��	�bU���*�pɊ�e4@ڞ�񶫷e��!k]C�g��}o��U8N���OCk�Ȓv�m���s�����X�5u�mJK2Ę	�z��F��,�.qxP�e�4-δfhQL�$���0RiM^fY�]�WL�M�ݣ��9��-^wb�7tۦ�۩�1�N�T�]�SL�	�2tD\���p��e�]�Ks�mbVSC�׭;��s��x��mò�n@��2u�=Fm]'Y��T���h�nA:1�Wa���+C�y�:��cG����)mW[X�q�SEA;R5Ci�p+��h��1����V��a�5�\Q4K=�݀ e�J�W�W"g:�
ˎ��y�f�I���aDQCZU�����pV�g7gLλjջq��Kke�#B2�^������"`b��:#�s���f���p���0��O/[s�9N��M��w��ǰ��޻ ��Xy0�I�:��Z�w�M�ܽgLnӮ�6��#���t.;f��D�nq�0CW�t�13���%�zY�`��e%)Ɏv>0�kO��s=��J^�1�=/�<S�ma1uy.���[qu ��=�Au�#=���<�z&,G:b��'[�Y�8�g��3٪�`�6���G�x�Wc]�j�Q�WAS�3�ۧ�Σ5�Ʉ`�\�Ku�b�hm`��Ě��5���)��b:�k��V3���q��;f9�:��y���q�f;n&�;�]i�h6W;�Y��8[�:6�"܆:lv,Z�vl�ÎckA���D�I�%`�V
��k���h���.�;h��ыfN�!�ms�NrWj;r��'�r��1ۅ[mI�� ӓs���d�܏5ƃ��%���q5�ҷJy$��;�v�Me���@�ۅg��tv;OX���ӫOiҙ���F����ɜ����*�N�e��FX�D\٬�	��S�R�̡�g����YJk�	��[�&F�0�
ىֳ/f�/r{��,#�sv�֞�wA0����hYRl�W�A��]x�m5e��[�5�ū4h@6�ٌ��F�;D��qu�y{-�k���g]�N� �^{�8�h��Z�-�j1�U��e�e-�9�k��)��Jh�_h�ӎ���c�?����\�W���Ñ�Y2������<Q��)e�zVO�u�%��b �c�����)�܍$Q'$�op(�Gl�
�+XQ�F@��ֹ��Z�z+����?>��N�ȳ�?vk����7����^�,tqz2]wE�#d��N&T18��!�E�h����4#HCk�!E_*�mj�Zs!�Տg�����nIBF�F m���`�0��1��.��B.6R	"�G]��*w{�g��}�S��ٮ^n��U��H���GE�DP��A�� �-okw�D�;���MďÍ/ a�~���M�np�#;Oǋ�N�X��TC����>l9>k7��ya����ɕ<�E�����*f�� �B���z^��N��eD�D��ܼjcd�z��c��{Z��a�ח����a��0�� ��)��T��v�М�>#��42��=���� 2���*f�ٽ��
�84�S�vJ��0�E�\>p������H0�Ή,�W}+��%!(��A=�ln�f��L^읁��s�;�poS���ḯ�IQ���Zm�H���X���2��5�XO����<ؼVtc��E��b�sB�� ��~[��M��2+��TF��>�c��f��,���Z�mᇈ�|��f��_��O�j-��Y;�bυ�4�D{0Ua4j��ck�eh�~��0��ܮ]`9�/D9$�u͊U����퓵r-����]3J(���u���S>���P=`�k����{�*np;(#-^�&����܅��If�+�9���v�Q� *u�I%"�$�4+y���\��֬az�#ǘy+�z(�q�1�7ٶ�s^�`D�X���P�jY�ح��X��GHX�8x�{yx���{��q0p�cR�ʴz�@��cf�{���/yh������BD�^�%ԕ�P_�C:�����G���X@˕c)��VyP���J$a2����i��6�$��`�أ廬	����-P"\W
�H� N�*�+N��멼�]�w]�M0D��['���"8��-�A�-�G�-��k�pR��y�I_�c�;\/��Y~���Qܡ�6wz��t�1p��gr�Y�8p���oh/c�c�ҤBQ�I<|�;U;erx�`DXzR����ƒ�ދ�Y�����[LF�6@���IS��U�.�z�=&t��5��F@��ۛ��5�o-��UWM	�.��e�z�$�z��X�P�7M)^��ι$L�X�_a�G����0��c�7݇�/T�ܽT������G)�����X�{��nK��>�1�`��=������	8�����z9m��5�f�bz�c���Xs��I��Cf��أi)¸!P1y�Od?n��
�=��=<x1���fԪ� Y��^U�o��`���`��"mX��12�Ij�ڐ��w�twf�3M�!v"��i�"���n��:�g,ػ�!�6)?�]��w�;��w�"���=�c�����17$�����>��¾��`��>�Ob|Snz�{���
s�i�"&E!�`�:b�>�&���<��4"$-8�P��y{�� wg��v��LT[�Z�5�(�/(�K�#y�����؏�U�/�&3o�Z�9�F4�xǑ��,�o{��3�{����6��E�6]��v�L�]�شQJL\y��M�W�Q��\S=^�=�Ҍ�)n���j(�JI��������7��k�hѥx��e���7�=��ky�+��ha�#wn��~�������l���p2�!�S�]�:�c�W�p���v͋��E�q�[�zP�!�`rI�v�/��=�6�d�R������ u���i{���M�¬�,F2w'�o��:�z�V�"q�#�7#�^�05y�ߠ^�q�g���ޭ��]@��]ǹ��|���Y��JپI�s��9e.V���{���d�D�#!��H�ިqR���ƒyE����G�Ⱟ8h�>�Y�w�9�<��	�λ�7��ۺ�_qe��.8Q�&��b�ݓ}w�����	^��ˑ�iʋy�9��A�=�Y�"N�#����u�5m1����M���0�д��"�J�����*�0;9#s��W6Md��,����v��<����9�s�o/�pc�,}l���eY.��*u����3��{�#/R2��wR�ٛ�hW�����7��B9�����]Yj�K�lG�'T����8���)c��v�^OY��<ױ�s�:֋
�7JZ����D�,�Z�gj�����J砼N��i�0z�R�V�-��K�ݼ���`�׵F�VO6�ͺ�^cΘ�iZ���ܪK�̠��y�Pg@i����&�hl-��#6�.5�0�gD������ɖ�����n���PV0�f��!�pFQ�B�耲�b�D6� ]��s%�Sl��n��:�&H��%�6�Ǭ�fu꣛v�"۵׳P�h@��M8)�&����\�󭫭�tɋ�H���y��]罫/������,�z� ~�"u�Y��V%�š��$�����Ɔ�
6M�����X����(K��!V�M|q��Z����yq�x�u�˺r߯I�S�l.�{"��ZNK�Ӻ�i�9=f�]���묒����n��pŏ��rw��~ݨ��e^^��NJ�I%(�[vFQ�I���
��f�ݻ�a{��6����e}�s�Y���,v��V��C{��s��E:��bD�m�$�Vz=�����7�3Ѫ��/����a��(�n������V�IXj,�=��3��0�:!-5�&�����.8����b�\vBn��C=n��rm�+s�."c.qH�l�6���M���Z����;x����mJ7O躂�iU��(l�M�/ޭ��q��!绘���kK�ce#�4<Fe?w�n�������5?���ɶB�A�=d�p��jvl���K\ߌ�s�����2��meh�E�d�5�Q����O��ˁ�/n9��V��|/�V�T� _&��Y��K׮���Bz�]
��$M�C1��<�DC�!]��F�5Qm�^�癵o2:�.�uA6�����[�wޙT��1.W�����RJq����C�y[��^Ӟ2��>E��%���x�<�y9��)p����{��ŵ0]߫��$P8�P��u��5ӓ�gK�)oYN��ޫ�-��	������ �O�M�����>��_��2:2]�R[r�Y�@ىh�0��r5��N���;*�G�\ei5)ڱx�δJq{u���FҎ8�0�JI���Y���rf��Jho_o����׶x��>�@��kۋe]��$mR�@ UE$��Vn1nO%�����F�u�&�(�q_>��-_���5d����Kb�^��y��3ɮ���bF�nDUmq睧}����~p|ho���Q�|n��tEW��2�eꏦo07lC�j�Ǒ���B�7�ι%w:ͬg��,e	��8`L�ad��^�9�#�:�0����
�VW�ȷ�e���6OI�{'�z��+���1�I*;�Hj���+��%���\)��d{�ϵ|�2n�yOz�<�jëCo�a���z��׀�pJVh���&P8T|�i�pR�rR�m��Y-)�R�V�ߵo�V�Ei�x�3V.k��i��!m�H�B/�$T�h�:|��q�e۔�=��t��;�ش��읬�SHi2�9-�~�]s޳j��v2�Z����t7��x��ڙ���ֈ��������<�Y�vOx#�H��i�ɲ�M��<����f��/c�j>�Q^΢_L� ��j^!"~�ޮ˚�Y�!r�R#�Ol�-��D)���	oz�F��{�o4k���O.�G���}{3Քp���8�՗n��V7�69d
�/'h�!���b����^�OV���Ww�y��-a����}�<�Q�N�s���icKԣ��9�n�0�:��j��!�R�2�K�]�3���ڒ���+M�u$��&@.�}\�"s�Y��k��W��3�NU����<��D�"$��a������;	��3�<���KS�ȭ}�^�B���^~o
�tm�Z͊��վh�O�H2�ICK,���\����n��:m]{jc<6V���8+B��N\ UM{��ڎa^�0V��y���k^��,;�-��c���e
V+H�^2�E�q�hcX\�u���Fe�����<�����O5�dp"����$b�k������o�wN"55-�>�p�(�����S���ؘ� Ӻ|w�7�[t/����;5��Eo ��9�Ȥ{�]��9xT^\��Zp2���u����[��#�ܧ[����6�e�ܟV6'���ܨ�B�N�:tl�Ib���m��ǂ0 ۔@)����:�}�=����vKe�s����i���������y�T��Ռ��'�d\�Z�=�u��z��Z���r�Me_��t76.��(��	<xr�h8���0�F���[CUYӛ�M����Hn&���[��O*��.�
�u�s�ZEP��]�g^�6��W��a�7 $ц���T��m��a����kg�s�Բ���9<Vt����ņ�ҵfV��n(	���7R�FݣmrH�`.�b���'<i�F���vӭ��0����+qXd9�ǿ��{@�u�	o`xU�&�]�^%y����{w\��uذ�g3l�2S!�5���h���:�o����=�v>8���]J�cWb:;I��k4�l�!�&���?������p�to���o���<��Ȗ2W ��7�܇^���0fa7l��*��.*�}!+�󷙹{���CI���ΰ�\5�b�����u�w�md��p,X2��y�rp�d	���a�)�{$ųi���衃��k���X�ž]���H�a��a��?^ï�¥b�|PE+6�HJ�r�d��k�ti�{���8��J�E�����y��&2�e�u�w��w6N�D�y#AB�x
����&� �U�p0_�p�[K�������^�~sa�z����:x["/k�e����x��dP��km��D(�"q�m.ͻ][78�8�ww$��f�8�P�睱m������q�y��n��l��`v��Ys�L��x^U�s ~�U����ed���[�
CB��d_{ �D�II�s<L{W�T//פ,�o��m�a���u=HV6��bC-�%���5�.R�96�V�<l1���)��*l`����x�ah��h�2�Y��:����ʼr{U���U�;}�S��~���s#U��.¢25P2[�J��Xڞ�k(5�_K�.� {�IӸ�]1[�Z�䪬�'���l��I�!� �g}�I�WU��k1O�<�e��ɞq���ӕ�V���NJ������	ֻa{<��1I EF�"�OGn�{���s����7�V����~����潊�p4|w�c�?T���۷�OV�(v�bw��ԄC�.�f�z��U�;r=x�{�[U�݈���i����	�iH��qߨ�%7ޓ03�����H&`�◥���-��)�:4�������ǜ�g���?0`A��I+-��?�ﳭRf�osɑ�h�(�MF�����������.�Ovp���Ae95�A^E��
`{�J�fD��Wn�*��ݬ��u�t���V�����G}{pt���OƖ�8��cT�4�ͽ�P��07̾����&�Qt[aqvN�4:+p �w����J�|0�u>�;�����%�{W���H	��0ڛ�<��yJ򓘳V��x&k�2%0iQ_P��+�����=����^C3��P�l7���e�T����t,cܛ�Ja��=n�M���)�_ùoR��3:��H�Y��:A5ϊ�u/+8ɈmbW��іf���ĎI��M�6&>7�*V�� 6�+��܎�J�R��YEmp贴���0�38�[�4�r��oo�^L]�|z�o����;�tM�M��K����x�.-P��H��|�s�"�4N����Ն�Q�hDFS�Z���b��qL��7���vBD���ά��;y}e�%��>��L[������F!��\\R��mjƤ+��^�����Ў'b���ʥ��FX�/k:�n�eLyV��G�·ٻ�^���Y�ճ��ut��`ؠ��rA�,)ɸc]�9WVS4�`-Xx���wct�Z������U�
���$�S��'ŋEJY��u"���$�X�$F�';n�ޥ���5i�5���r�iQn�t��R�(�$Ɗ��07'X�M���Jzv�����*�Ŋ��t���;�]�P%��\Sjf��fd��E�[hc��s�u��:�66Z
��)'v٭;�>�Q��%Ւ��:s
��(Ӈ�}J|�C2�
���%����n����Xy;^7c�1K���T�(Z�g"Ǐ�_��z]pME����n����f�tQMјz�F�朼%uR=N*�oH̬�
�xn�zW�(�m�h'';�n����}K��۠�c/�s�N�H_�X����.7���̾�=�̼y�M��ٵ���*4��L�a`�>K��:��Q�݃��A���$�1P���`(�Qd����v>յ����+�>���L4�K�b<ǔu�C���9�ݦ��zY��&2Pq��,�N��T]�e������w�{+� 9���}6"W��׳4�G}�R��^*#���s�NΕ˻��WC *��-#5�m�����5��}[:��{�i��]�K'z��t�x)�y�\0��Y��r>�"p�0��I�0�c9+#ٚ��.=;�s�#��4��KM���(���`7:/�uQqnZ�����nE�7kd�8N��dB���bv.�"��T�ǳ�G�2�)',-�m@1j!ũb ��M����nߥy+f��q��GnШ�������Ihu꫏��Ǫ���BZ�{�*]+��9��jc��m`�^��H���t�B���ڗm�n,#l�ųsL6c4��Kڶ$8b����eӵ䒮���.�p��]jڶo��z�cio�;~{C�`����׋��ESw%���ׯ�T6l��&��By8�]<��V�w>C���E�K��8�*�%��u��&2Z�:�/_mO�߽^d��\�fM��L�
J�An�W'�Z����ۆ��6�Z�P�ӱ��|�����vͽ�>����<�x\�$�p^a$êڿ�<%צ� mE�>5����{=�	��3�v])�t�w�s����=�Q;���Q��90��J($���d6�K=Y���E��lܔ��^�μ��dV�7l�}�{�S��i{$2t��+e��E�pT��D�MO��U#�ۡj�<7Z�wY��d��ǡ��}��_/�Ɏ��1��S�V��������FX9.�s'k���g���Xfm(��e��ʐ�u���S�*T��w���u��t��f�@���p������Y�cju�L�L�Z�g;�[��c�����غ��0�u;����<���Ç�����x]�;��]�=eٮ%\p\W��;���3�x���Kv�,-��q�qYB5���l\Ue�#[���x
$�u�7b;�]"lez5�:+\����uJ..�$͏���M�����Ԏ��慄g<�̡
fW��!޼�Y=�q���g6�\OT�򣒶���G,	d�<�ʸ��g�<8F�D!a�N�P�_&'���b��x�������t%��������+r�����-e���Xᷳc{�G�F&��P!`�#������2�i����'�����t��ϱ�>�#�.;,��L}���,�=�j�0�B���D�^p����Nנ>.���y��f��e{'h<���o�{C�Ś�3����F���{�mjC�D�R���&H�)Mԝߧ�^u���`�⺱��v
~��&�)���Y�`�9�蓶,��:�ٛI���۝S�Y�UI�di�jDEDp������W��d�W���8��N��Qs׃D�0��QŃ�>�@�}�kD�~��rM��uԭ.h��"�hܨ��n�ʮ�t��sd��2��D�i	3ȯ����a�M�ϖ���I �C���9�I�)	\ں��,������C���}�\��];j֢�dZ7nٶY�F�e���rx�O+g��b�������;��ul>�����z��f�`���F)A��n��Vo(�c�V������-,�8�c��=��j�ǐ^U�
&��R�����^�����z�Dt&~���Fg���,��ꏭ�,k9�Nﰂ����^OW�H�
B�#A J>��s�5~�=j�*�N����act}���Lj�Ο6ʧb�;鸧i��ٹ���r����$���-� ���2�6\Ѱ�,56�H��jE5�ac��+[u8�DE`<���M6���E÷��c��>�"Ój������Efxv��ˌ��uTՕ�:=��h3*9$���n�Vݚ�eL�ʁ�Mm�����u=�;	?�>ha�w��X��bC6D�=�"� Β��_'��Dy.��<�|aX:�0E$�FBr:�7B�BY���,h8}aY�A��{zx�j�C{ؤI��N
�;��[f���p��H����la]�`�3vl�(R��8���:֜,�t5l���}��̉,A��sG��u��S��GӔ�d{���L�!�:�@G+����ml�{ߤ�/��%��I��[m�_2_C���b;^{,u!m�ٱ���&�+UJ{>��ae�f�n�_����Sء�i���O!ކ/=8���ܧ����$��u<�A�@�aȠr$r'c���>><�E��􂬍5������3~��qE�=/����D�4�r�R�7��%�tَȂ#�zh[_I�����Nx5����p�W���t��<��3iaf��Bޕ�ѹ��'5 ��KA1h����������~~�M��EJ���D�>��B�E�I��$�D�g�n�'U����6���~�S8ߖ}gM���:��W݈�ur4ݠ�"��ߚ-AA�E�����z�!!{o���W�@A�8QR�HҥQ���vsW�*m" �E���E"�8rL_�g�:{�4�aW�,q
S,׳�0�BB�L3
2I��~H�5f�Q�*��P�^"�)�$1J~�z�_�P��2��c����O+�����;Վ,]��b$�"b&����\׌�A֑d3_P ���a�P�B��!_����+<Q�yâ��ȣ���%9�_?5v	���r�Wk�jN���Y��Dҭ
K(�I^X3��}R&ll�?X������3j���^j����`.u^�	f�1����Q�3Z���3�����Eh������:Z�=���Q"�A��s�Rdo��J�>��b�7+A�26,�{������#�}�{|��^���n��e
k���#�"����i~��Pm|��|�B�3�=z��찴��4յ1��t�	ζ.���h%痴�;�չ�o�D�t�1͎��R�&������_)��d)߾�|�X�H��X���V|����2�=:G�����,{}�T񙈋7HYz�++�T~H��"�z������"0F�8���Zf����O�٢��<���\0K3�A��}�"��#�9.P�=�Ve�"�*<B
۾ȢC!Gw�ꖅ'処�w���F�!Ɛ2D�qN�n��ć�,�G���-�h�n$ْ�F��Y5��ώj��<������ڊ�^^#p� �~��1ISΠ��4��=#��DJPGK:U�,�9����m�C�rڡ��Ba�#'-5�lV��0D%�Y�C{�hw��)!���l���"k���H�}���H���q�#>��Z�d�ECH���U�ȼY�1�j~}a���dE/R�q^0�᷅�i񱼙��PF���zǢ�ӆ���H�"���}����� �!��
�Ǻ߿hy~�٬)���ݿ*)"w�\xPy&UH`m�}f��bA��Qհ��t��˭z~{��3�q�4��W�M_w)=/E��N!#H�b �1�FT�����<B5��s�F�U�0��b0݀��!iI��mJ�)��I{M�����t�j��#h�Z�xC<U�2.b�Y�����m��>kI�1�Y5\<�wl\��c'[���Cr�#�t�D�{��u����z��䅮w%�����V��H�lh��y�l�.%fn6LJ�n1��6�]� �vy��v�;Z6=X�\�g>z�W,u΁��K>g��^��x�����%K�֠�J\ݩ�e.�K5j�Yg���~�J�`#���:�uQD��=?/S�f����4��gn�f;/�Z��t�__���Z�*Нo�^�c�F�-A�>8yOx��DN9�)#pس����#����M_c���"*����~�CIـ��ӱ:�x��w�۱a_G4I�yj�#+�Ei��$ߚ.#�_N��{��J!�H��n����""I�q��7��8�5홏�U�
#R$�ġ�g��B��~
�]��Y��{3]�����7/��臸ĵ�7K
#}ߖ��Q(��IeȬq�f;κ*�g?�7[�E�gL��gd(K�߼��:D��nğw��
=�RG3����wo���~٪�Ӥ����d�:>'"��i�W�J��X~� �,�n1VY��'�t}�c�o����o͙�6в�/F{=����a#qN ����<��DϺ�"=c���J��	��cN A��W��jֽ��d��1�=����r����s���Ma�2ݪ�H۳~τOy�~=��W��A\�Xh�/P�����m��6I��irDg�����V<��6���S���7̄NT>/7}_9��VX����#�ȹ_-)b!D�FI��;�+��O!�%�-�N��)�=O���gUmy:��Su��ŢSт�����X�6iɑS�;Z0 k't2���{$N�MY8%��\U�8_\��î7/����^_v+�0�;&���$C"�"��;d�B�L"R�:�X+���VvN�|>"��(��M��ħMq&�v/R0�4�^h߾��_,��:T+4D{�l�s���=����|�b�n�T���-�8��]B�|�=���*��#�jC��}O�0�E0ffs�:d�C���+\)�F�K�w�,2��(���4O�z(`9�Qd�Fȁ}�l݃�}�M �]����!���qKHe?@���F����03�����X�h.�g?m�q�4�~��l^`@Oz#t�����]}F��rD(_��4	g����DA5�~Q}�H�Q����P^����G�J}���U�����fM��Ƌ�J�U!���J&؉(K��2����Hp��t��������d��}�g�"�4�KT}�U��% Nje�;�M���2��}&���� Q
�6}W��a��Y0��D#��'֋�*���Z4AӘ��>y�}U/����Ag�+c'V��N����A�'Wc���
ˈ�\�r&���"�sf���7}�|j�&y�⍟_XG"b�G�Ɯv4�!E�L����|:ZL�4�M���r+�%ƃ%x�;���^�sd��BM�ح��`���b��j�����5��H��wjs�1�Pa\��VX��`ܬ�#�(I���U���-
P��2��O�]�KH�o�i*<��j�q#$�6�t0��}hDs7��蟣ʼn��b���`ʚ,�O���i��ɠ���%ZCR$� ��Bq2,��ޡ�C0�]�T�*ȭ�b�Ja�G�D""cH�]�\�!,�e�J3�M�Y9��/S�����ΑFZ� ���#��,�ϖ��o�2Db���!�{�(s)g��'V2���Ѳ��Th�~������Q����z~�1uMvq�β�آ�7<�7]�{X<I�]Q�`�Բ������Y�D�$�L_��y�/ۯc0��4~p�Z�zY�(s_I���,�ei�X;#yL�]d�`i�n�T~�Ύ�a�����nH�`��3�gʈ��@'�{n����9GR\����1DT�g���x+�P�e-h&�h����V	��4�&�'���b�l!~��8s�������8'�+����
8�:x�e�h��E�Ȓ�MA4��_o�]�~�^�ے8���H�7q���A��,�}�>��ڊ~���DRD�4yg�*p��P&��^$����tu��z��x���f�wW�gH��g�(ǑvC��E"��@M/Ncd�����kƯ�z͟��N2+2����@�<֜��p�tL��z���%����o�V�n푈�@l���c4/�]?��r�S�G�D�S�G�(���(Q)��.EC�2q5iFF{���Gԑ��u\;��<�z�5E#�ye*��{ׂ��+�><|E5$Fn=���}R�hi�O���I򎿨!����z��.�A�r9�A�rb8��Ф2�յ�m\msg�9㮑�H$e6�z>3U�a�f�f��/�o�i�dQ�$(���E|u
8gn&R�Hz7ڨXyWcdxT�k�|d��`�}�7��(�d��L�^A8��2���HM����f��&����~4���%^ �}�2e�f��o&�j�;5���P}�}�Vu/h��c�)���V��e��~#�ƳsS�O�}k�K�3k�{>���3ǽ�����mI��<��=�Q�k����	#t�e}UX\P�����O���H�r��#B)0B���ZZp$�,.I���Ԭ���5�&�3��4B+�f{�G�Bo����z�E�R��6t�D��qB�#qI���`�<�^�j|�_���m$Q=���B�qdB��g:|a�|��<aex�]��$_\�9�^���}Gu��O��*6n��~1+Љ��٫8���B!#U���+�#�!�4� ��}M�u�}f�f^��>{��6��@��t3jK\����Gnv[���c��6�_l&^��tw����]���ckw�5��|1h����]K~xथ�oT�qz�zI����;y�U����z�/N�3��Q�4�r�[|�V�B��;�����7�+r��*�	p�U��%;,/�D59JV��'n�S��9�]�&�w��a �>�'p�&r���ü�"�{��0�q�̩B�	�_eZ���Y�I)(�b�+�5	����w��L��N�,X��0��d�T�!�,�B�dl/	�S�8��Y�����^����R���5S{nI]�W*�\���4��M�FJ/z��h�(�5
������1'����J�����a� �_��*o�yP�Ch�.	��6pꂕ�N�J��i(
�uj�=ۙ)�'���gm��J���%��eA
47p,�a�����=Ų[�p�H�k���7�������T�i+߈�E�nʣM\�㰵&mĳzat�_L=l`��DaGjq�I��'������eE��qȠUuzU!i�3��y��n�uI��2��m�.l�i���r�U�F,=��d��{�\cF���v��N�+���� 9�]&��̰1�էp��w�(MK�����+Y�LU:�cǁ�	�0䆍���Q�G(�gr&.�5��ews4�h����O��w�����}l�A�[��m��(.��fX�b�m&�)"�i)�:��1�<�3�۟*u�� �eY ��;B�hΆ0���P6�e7K��%�kΜ�u���uo`�Q�vCգɇ�����]�wk�B���';O�0�����V/��Y|�t�Mn*�����g���K�O����G#�U�zRE���������u�"��)ݭ����y�S�]���R1�6$�]
�����0� 2َ�R=C�4���6�.��ff�j�;^Xtc�vV�e�el�+���84R�M�urC��Bbdll�L͞T�+�80�ρ����}���\�"no0���(˝Ld,���� e ͣ\L@�bK�(��&�mn�Ύ�s5�Ԣ���t�;�yN޶�Jϙ�GmӼ�j[/8���B˥m���hYƐ���C^�H�P̒�w,�e\ن�%���Ɠ����i.�&t���Ѵ���O��M�Ye��Ʒi���I�vQ�K��.bb� �qC��%�}7y�ujBr�n�H屷N��PH�e�k�p�RgP�%���S��.�1nHBf̷sMCǰ&%Gk�����8a���2��[Zq���Q��fMv�mt�Hs��v|��d��v6�L;:��H0bCgE������GR3#v�$�+�H]B�B�'�K�;4�㣞�����{j��;�����
D��F1,�Z���4+�	AS$��jIs�1�����S��^��y_\�sS�/�u&�8�n�^ۭ�Z��W+���T��M�7���=z;Nj��] �lf��]5��<N������7��S���ue�z�Smِ��m����=e��G��{m�����.#�)�]�ʻ<��k���q���;�fs�8�h�m1x��1�CY�a��v!����]�R�1���ڑЎMe҂6�Cj�]a�t�cl����q��-�Q�4l"�dTۭQ����B�ЌjG2�u�2��0�U4�B��k,��@Ԁ�CZͯZXBR�g���l⮘G<���pw.9�E����m�+�X`v��]5�`�Q��pj���#���p
�+71�tn�6�e�d՞��U
K3YSgF�;Hm]���Q��jv(�a�uW��wZ�yC.�oF��&;mec�^�s��-�{[��y�D�+r�[���X�<i]������kZ$�z/m�)�P��s�I�ѷ|Oɱ��ѻ>��:"�I��Ǝ�n��K�e=;d����b��%N725h�C��n!��u���@��|�3U<�֝�Z���Ǔ����ol�Rb�?�����f0�r����(�"ȃ��򡥑Z�g��U���MY٦��z��f�BgJ<Q'v��(q�&�@:�-a�Q>h{�$@��cN���A��Ϸj�&�U7���~AG��h_{�:�Hg�tѦ���Vw2b~��l��LV�x�t�Y�?������\!H����2���i�%��:Qn��60�`�Q��=u�Eԏ>���5�#�̃^�A`\D����(�>�9�K�d�}��� �"�4�*��q�H�(�����DڬJ#(L/^�B�"L��-}GިYb�di`�"�ϲ��`��CL�n�O�1�pC�~ؾx�>�s�"�t����(A�rB���OM%z�}\�����\��zl�����Aq>١��/��$���8�H�� 4:�(�>x�[�ܾ����b:G��N���i�� ��6��guX�纨�9���5�7�9��'kt��Nò�$*$Ïy�營h��_ۿ*��\C�4E�E���u�dH���Eg�M����;F�đ��i����vF�w<r�#	jD;�x��d���0��3�����a�!ϫ��M�/N���AC����>��{+�
ww�)^R=���\m�D���r�Z�oZ��)y�~)d$g���~)����O� �k��V4��>�H��"��G�Yb�5���S�I9�({�COd���G�|���dgL���}�$���E�
���yD���h�$)�CIԌ<�U<Q�ޛp�(�_Y����_Xi�#�R�{���~�����Ь@ѫ�y2#g2+5�6�:p�`��z��6��qH��9���ק>�����#׊�ދ��\p���C8A�*Q�U�#Τvg�(im
!(���r����z�:U���p��.�]ϾoB�(Qr(�H/�:v�$�������u`�-H�T� �W�z;��ʞ��g���:B8Q#S0}��ƻL}b�da���!��>�#��H��c6�X<�r�4�������,�:��fWA��R[H��A��.��Fonv�&����q��#��# ���-�O�o�I���
3�[�������_z��t��4PT�T�V(#�����f�V�F�"H&�=��i��4�n:t��޿fH�v��
���r�V0u�~���H��U|�^ӝP'����F�E�En���*ބE�"ui��lݴ8����	_)xE]�f��Kx�.�!7$���U�H��Y�2���vF�4�7�@Y�Ƞ�x�2x|*-s�1��e��:�Rt+�).��W��C�e�u�١l�|���qk����,:��`I�.���u��mͺ"�.�����`�Z梃X����OP�ɥXG�2B:A��߾�4�4�u$O~���IA#�d7.��Դ����<��4W{�J
�T��>�,�-|�i�~٭4YF��D4��iA>���s�ʓ��֏�g����4��x���|E��RaAi�څ�$��:l��+���f��+�'�N�N^�D{�ln��CO�d���~��^2Y�jU�E���וx�h2.�.��C�bc������6'n�����5�OS�8��mp6��Qe��7\�k�<�m��bu��H�$�=�	,>!Rk�~�������w3��+�/zر%�$q��X��+��7g�84�x+��KHa��L��m�d2(� �F����:�L|�P �1+	�2�6F�ޱ�zCJ<N�Pt�����z�P���#O��5v�*��6,6h�SM�R��u�-��U�1��<A��O�:��(�B��X"�7�cH-Z�\��H�B���zm���fr�y�Ql�P��xŅ�a��I�!'�M�Ǒ �X�?^=<�����T$����IV!�ȝYyڭ8]��6`3ۛSYgi}�
$�nM�{-�׫�����h����<D�皪���f
��B?��І򋞞Y����L�}��d��-*�-e�i�[+V�AS�pS�Q��{[ݔ�Y�.�>Af6�y��e�}5؏�EPA�I8��;��@�3$�-��[��ԥ�$Rw{�ml�i!ܠ�2W��k7��t�"��Y�Q�0�tY^۵CN^A��Ѿ�d�j�+:�B��'�=ٲ}�L^����C�0L�H�:צkR����7=�l<-!f�+��뎷`�l��!�r&�i''�H�~C�#d{�Ӽ�[���Y�7��������t�_g�b��g��l���g�H&���|���Pg��6G(��~haR	�(�fJ�JJj������w�;�:��D�M8�]���}�A�ǋ'�}��:�r��0zB�>��a�F���}`����H��ڽ�)b$��f�A�r� ��E{�m^�K+���t���t�Z*�fm0��Oȇ��6;��x��8j�۶�#��e&H�-�(�}��ԌD�h� ��xI��RDw����~	�ƈ����/��"�
0vo��n
?2$�ǽ�V5��]���k��k7�����D��d�P�=��uXs�5$8�:F��t�l�W�e�N��\�d)FӖB4�UB�UU�A����6B���%��#J�A�ϲ��f-<Di�5�1]�K��?O�˼�[w�h�j�u;Le�kx���FUǩY�(�/��4Uw�;�iȬ�lؓ1�bEy6��YQ���i���FЌ��ߞG�ۗ1�7/^^t\������\p�����0\�rW�Bv�#���D[>��rn^0A�^I�nu��Eͷ�R�:�iwY�eږ���ͳN�Y�vٹ\f�J����\��bO�9�e���x�Bn!\fc���t�{*m���q�+pomWk�A��Y����6�j8G�֮w1s�ݶ�ܰ���<㱷j��vNu#q�+?s��=����t�s �{l���޼�΍&�ZrF��s(l݇/����w/�*�u�\�GUf�n4�������V'߯���~?�Y445dQE1���}5��� D��ٳ����c.<)���p�հ4���0w��J?Ja�G�[���s�^Ψ�f'$(D�b%Xe�%Q��r���͝�KI;k��[<E�ǭ�o'іMr`��2,�j�7޼6<���	?qD���M�҈��=�z~.P�<���c�
e��&2�R<8D,����X���lm�ե�A�c�#�Ŋ�8�PD+�W��3�S5��ȃFȼ����l�"7��gK"��Z�Vh�� ���9e��r:��x���>�T�w��x�D���l����<�)Y�Xp��y��0�6w\(�CW��Cy4��P�T�P;�AdG2�`d����4�4)5
j��5�.�_\ID��'1�#M���� ����W`�DQ	l}R�W��M��zk��}��"���A���Xt�t��v����A�"��%�<{�ݵ�IZm�S"��HYm�6`&r�d��f�)��|��ZR�����ѽ���keA,�]��������Q>ͨ�V�"���A��!E��b���Y��n��/��r��
�b"��F�����C�A'm�(�nȡ��ߡ*
F6�,�%s�����V���1j���骫P8̍���̥������#$��N��fn�GE&PyN̗(fj�[dY?L��f���˖J�����4�l���ʏ0��>�ZBє���q\|��As�lX�z>�p9/�ɼ��պ�Ȍ�[ɟ�)���X�~��	|x%)HDIn
�*#O��f�_����!��1�E�Gy?I�{��{X�.*�#�6Q�~ɯ��;�)D���~��ZDM�H�5�����#��nIlH�4,�������=q>|I�y�C�]���E��mx���+�PA���,�޽ŝ$�T	�=�I{������c.o�����I���>�~)��M@�
T8�4G5JfE�~�]�9d�w�GZc�Uvȏ���;�m}p��_F!>��AjdAց#�/��w40�$�c�.a������Te��ZM!�A!H㓵��E���F�ݥ��θ�y��dݳ�ӱ�pM�[v�z�Y)�{����<N�d].���ŦL���E�n�{�_w!؄�����~T��5y�ҽ�o��4����\C�j�Wϕ+�3c���0�1r&�I8�n!']b�D+՞���$��ߞ.>>��J~y[s��Iov8��a5ӑ_q%}�JH/޽�!���3�\m\�$����@���^�R�51�a�b�i*���"g���CƱ�%������%�75�ZG��x���}5L\���5��`�5^����X���9�!�2[t���;2�8H�+Ǫ�ujz�ٲ�^*rhu�	�/My�B�rE��ڇ(�~��A)+J��l�]��O���[��[��sPJ�.�-u{�m�"5�!l�ؿ�?p0�Ȧ(i�z�|���=��6~��9�v�RU]�L�yW���b`i��ﻅ(̊)CNJt�oB`�H���f[�z�Fj�yv�����|}�N4wVJV!����~�Fm��4�'}n+�O}�	<Q���b|7��'ZZ��q��a���C@��������(mS�j�n+z��.B�\6�@�l�y��$r���B�HD�ܱ��Q秤V/PR����voP�d2!�������|�g��z��N�d����5�ϥպ��4��a��~z~�.3 %�� �x�ʊ!��a�*d�=5�w������ω�.�A�T_�:(aިA2E�#��b��Ρ	}F	����ŗ���ty?:[�"O�s믙֐�F�1@�N*t�Hi�,�u������8F_@E�G���A���W�M���;�S_D g�ذ�2 �E"�{&�&4�:y���c�(fi8�+ZPa+_'�+ް�~��h��B&�$4�6�2:sƢ����#�a�҆�^�3�L��Gz͘��)<�@N*�CG]����D�F�n��#cb5�\���|z�lh+7+F>6���Y���s���i���l*�ʂk�K�{3rV��G���ӤT�`?p�@�06�������Di�Ϝ/c�hID�t��E���G�pptEt�5�8�̸g�!��EJ��B���z�\ʽA&��H�>�=�|<�>^��E�ʄ#c�9����l��b�<1���b�K��cm��d\�{]�8�b��O���R����D��H�kU$�"�}G%<���|ρ�$�!�uފ��o���t�ʻ܈�B� ��E\��Q�F�.�#�	���7	q$t/�#��B�q������n���,��I��8G�/�h3F��$Y�>�Ẅ���,���Cھ��Ǟ�Z�wJ[}�!�2������e$��$�d3Ə���R	]y.(cJP����7+���)l	0^HI�Qhi�s�ث'��^l�T2(K�8�ـ�����><�OH�^7���0�z$z��7��<������ឋ��Q�(Q�@�/��%� �D�8�z���Y~�q �nzL�/^1�n(q�+#őC�SK?wǸLz؉�
�
p_3���`�HQ�_�+�����2.�Y�Ef?�Fo�|��y
#Ě6|G�ފ5�j��#���>�gc��B�~S�9X�0���٪���)������Tg3����1sy+��f0��U��%��'ak�9A��U����o�v�����nÎ�+5I����$�B��4�iyM���Wr؏���/�����Ԉ���
��r�!e��%�3��|y:Б�]<<\�<��]���:r�I���q������dǀN�s�=:���ѷ�u�$3U�x殶r-�ɭmm5��[����bfĭ��;�R���]��\8��M���-Ÿ�kB������g����m6����c=V��V����m���Gk�!���qq�bQ��<͋l1pY��7]T�I�������e����
j���IL��������\ՒY}闫	+��	�9��P��I��fLȁ��,*���~"Oaaf>�c��-c_Q�D2.�f���0�&[���x�{����I(�dz'�ϮP���Y^ӣ�P�PFk<�9�diFȿ)���z:�P�_V؀�#���s��q�턶�A񼂭����F�w1��$q��I8�i��Ց�Ngn����Z��?{}w0�d��П8*ٙ�?V!��&h/TG!1q��I�+��҂{�q�F��|CF&TᑨS:�A�f�5�WS����p�E�~T8�Zl�}&Qs\ww�+�U��Y}�컋�y"-e��R��Ɔg�-Z��h�$��r��=(�V�Iy_7��p@[,�L&8��hq�$������7�r$�H�УU�K8&�_����B\}�_Y���D!L���vߕ{����=䌋�J��qo���A��\��4`��p��w���f���KX^'�vz��:��<<N5��xd�ݧV����������?{+�4�6DdN�"��zد��#A�(��޸�5�^�vUu
���w�(a�&f<G��E}�)RCլ�"ϩ�(@��$��d�AB���4GI�%#������W�|�xԭQ�k(�����jn���pu��O��6mfv �醅Զn��@si�����i=��!�U������_]�P��$���+6>F�\ifNҀO;�ŋ�<pْ8�0G���Fۨ��+���c��d���̑8��3#��<�$a�C>�{"��V���_i��Պ�:B��O�NP뜂d{��U�~��%��a�j���vCH��#�rƑ��"�|D�*I�*B��b��М��8Ժ�)�Ux(���b��a�:C"�PC���AfƒN,0)}�{΍چE��aӛ�����7�����t4X$������m�Q�BPM�vI�D�j�t�v�}��V�:E!�I�����Y�o=�%W��Q��If�7�����0t��̟��k�#�o>LB͖r�}�X�2�c�O~7j�f8���.��܂
zv�z9��۟k#֫��7#���.���)�hфGZQ	u"M��#�zo�Y�dQ�=���.6t�k�5�3��qvU��ҷ�������i
��U�'Pf����SP5�w�-AG	8�W�v�5�1�"s��k%<���z,�ٹ?a�j����$�H�E!�^�P��O��(�Q��gۆ��Dc�������(��}��%��-�q6��7�TC5e��E}z����҉��o������3_ �a���`1Kӕ�q�yGo
y�x�ano�h���O����j�g�-�����.̠.ͨ�~
ܻI�8Cg)������n=�Qd��,���k����oJ�_H�V�QN�ثkg*n\E9��=`TΛ�N��M� �pg%)������s��������x�W\��[5T���b�ȫ�K{E��4u�O�޺#]d]��w88.�t'b���d�`i��s$��W��wĉ;0�v�p���qk��w*��<F��{&��@�0>��X�/��(���)��S��8��X(�P	|��:�u7�����';��O����y��Wy���m�Ɲ�٥ho ���T�Fڥ���G�<�6�C%mvl|�+��M�m����6��O�(��=� �ʍ�G�k�h�V�Ȼ�fk�+���}����wX�戵*�DyV��L��vIi՚�{�Tɳ�g�<����F�(�L�c�W�ۙ}cN��o ��,Q����Ӕ�fG���&����1n.��pe�:.��N蓚n��&���Wp�l�-��ߛ���\{�t�z>��!p�+��p51��6�.��`���Kx��;k�������7$7��uǛy��n�|�k[�b��� Ta���X��9�ZkߡY��t������H�qv��0j&n��R޺b�|]��cӽ�f��}�/Y��(��Cm� ��:V/P�Շr>v
�:j��`��ݬ�u� �����$���+7�jŝ"�Y��rP��=�����	²Q���i@�)�d���d\������6;5�F��y�0�(�h8��>�=7���
,�|��Cr6��F���$=�JG�r���O��,��S���tH�q�2H,t�����J���e��eh4"�	�=���:�y��c�����o���_o�(3�!$n�=��J��Z:xQ��C�W�<#����z��Q��Pf�i��QJ&H��C@-�6a���s���b��ɦ�>���{s�+A���)��Eϒff��(tֶ(�?Q��*��H'<�"�܁������2���a��+|�&nh��_����	���� aQ�C0�,�di\�-#z}�_i�g�O��ĕC"IjA람�z��$j9aQ��a��rYq�#ܾΛ�w%�z�3���`d-Y�����L1*HІ4��J���{'��i,�n
��Gk��Y���N+Hq�$�/���������d�J�B��g4�������e���A�p���p�P2�HZQ1A�&�5�빭g��c7��Ш�L�l�<E{�s�<9}Fr�4T��ۊ���I�t���7�^��R�7H�s��c�8
����>�d� � ��P��=��+�i��w/j�.�-t+�]w��	r�7��z�A�㧖A��A����'!�����=6a�	Z9_S���F�|��pf''��Ν^��#H���G������:�0Ɇ�8D�ۆ�8�](�E�$��=�����q��18�l�B���v���=�dt$�̐DgtZ���H-T�i(�%ě��H����^���j���q��2�����e��Ŧ~�B}Y��b6ĎF�Ǡ��4�A>������=:E�B!)<���T	�܄�ِ�sHgI'~b�>ʯ�a:������ cF[��Doz�}�A=DY�{.h-C$I��!�}j��D��^����y�m.wNZ�Dfd�1!�H(i�F���@�(ug���E!�B)Q{��Aԩõĸ����ht��wE��E"��(\��mߢ����[tzG�H�����`%CdH�#J��H������z���3o[��|Q�"� ����B
W�M���H4Ϸw�?B �0v�1��Z��~vkK�0�u-KPfxg�@�B �Ɯt7�3=5���쯣�t量�(�}}Ӳ1+��Wfz=`�l��$Q����5��D����`�=�08E�A��:)���]�U���|�2�m6�9R�$jd+�
�G��t�䋔����2���,t�K$V����_ǥT<:1�!$�E˝:��]D8b�����2��&W����`,/[�x�us�|�&�Vۉ�K�(\�n�:�\���"���Fa� ��B{qX�����b�(�2�>e$��͉㍵�4 �͆��h�)�;���0��J��65Ǭ:��6\Mk��F.�7�V�z��m��,��SDl��l�0��"үn��rp/$z�����Eu��H��`笹�(Mu�za7ugv�����fhλ[1ñǶod}�ƴ��,y�Ja����ٸ.�i@�r/��OƏ>c_�:�M}�y�Zzh� ���kќ����G�C��]{b�������W/_�k�4N/���;�D2��J�2y��q��m4�d��x,�Yp��=�zkige.b%�u���)�%�=���=Q���H�(��dW݈�+�dn/�޶+�g�&k7�r��|��"{�o�I��7dx�8~X��uފZ�Ej� �/{}j�����p��f= ��e�<l�;�}+y�Y�G �2''�M���$PA�޽<�gH����a��)��<h�fv���jjy��MȄ��&�t��l?h:l��zج:Q&O�K_`"�9z)�Ȳ�`i���tzk�;�(ף�GGN����a��I"�i�� ��B�^��E�&V��/��h��*���nxأ�I�Og�_znhD��ca>:Y���*�kB�4��D_��~�E�٪o%$M4#a���͟<=��q��<�̴��s�.5��"��c��5D8��zw���V����8���k�g��vC��G|ع�[�z�G|��}�8g7�P��v{���|�!�i!��}�پ���6PE����(Y$�$_��$)���p�:{�Dt��y���Zt��=����=S)c��u3��X��x*��5����i������a�Y��mZ�V�8蝔��
Ln�&)�)�3�O�f�����9��k��6�2,����vp�ey0H�:��+�ܵ_�F\b~?A��ѧ����Dmg�x�`D��d#j���D4�M�7�~�xIgvb�ԜI��nz������S��$?LжO��Vl١e�'�2E��}r��4F������Ĕ����*���YZ����=��֗h��^d���YN�y�p�$W�w�b�g�~�Bkc� ��}�	7��S�8W�خ�}#�\���y�^�C���p�mI��9Y��O��o�FJ���M�~��q^�٫�~�Vx���{}�+f�a|����բ�n�dA��>�C��߾_j���F!%�D(���z��~۾��\�@��umuu�����5���1�ڊ#�ˏ���J�??h~y-��!����%8���������e��>��Eغ�rF�gA���o���l�O�_�l�ģq�j )��dX2Ck� ��vz7��S3�SN���ͤI>~��s�	}qy<NeLP��Y����]��Ej	��N���u���=�=�t8�p�'-H����ү"�͡Z�.��ڨ��WDHq����i��&d�Þ�>�u=꘡�pP�Ś���;Y�W�� nru�E�S{NV��*��|x+�VqrN��33X_V�%�_����oGlm�"��Dq�x�z�U}�I�1!GH7��}��)�i���xA��2ݑ�c��S�>`�������U��k��:x_��Y0�h�$A��SE�O֯�8d�^��oxo�{���d�z*A��C����"J@Ah�"0�s��Q�C��
��w�vY�B=.B&Ӭ��;/_�Uý�>�#_�3>��B�d� ڛC�g��%ad*u?2L�"��?�1ؗq�e��&d�8�YD�43x�]H�c���Әڟdk���y�yu� 0��E�ԏGz�f����2��*昔<��l���|�g�6�p�C�����4.��d�x+Sjw�Q�G��딎j�N�e���f�($!�	5X�8G��o��ssbF�Q��._ag�BvU}�
g̋*P7}^��N��r����v�K�S����eG��/*�����_{����<��ʁ��q�����lC��l�����'�(���{�m��)H�i{u7���m֡��ݐ��Ӈ�0�&�h�G��~1�4�M�y�N��DI":E��a�Ǽ�o�y\z��F�����p�Z�$�Jn|��U2�	�8��M4<��/���'2��ソ����q��1�q�����{�'O^�G|���a�GJ�˷*��w5�s�e����{)n�����w��MkC���"�����+����	��,�&�&���W�yQ���\�D���\J�G�zNF���(:q�yet�	|��u>4("̑��?u�z*nrN���l��wwR��3&#��H��qC	�޶1���gj��"��+v{��ќ7n0RgGZ^*�MC�$^�$�?lb�Z5�����%�Hd�*z>�{�z.�|���6�f��d�[3׼�������{�g��"Ǳ�E��8^`���Z�0�<p����`��Ƥ:p�BXE��PϾW�=>��< �:`�#�N!�})������"��U$�?S\j��+ފ��u>���z/�u�M/�ۣIAw������'��;#�ۚQE��}�48��5$i���b�㔨�ǁ�p��g����xP�\EZ=HK%���Y�3>(�{���]��>2���f#��+#OCϒ�n
��i�*u��x��_Wt3�}ٷ��;�G]�Bpȣ��<x���<��ִ���w�cNK��\F��=oc����6�L)#�$��<6Fw�eO���X-}${i�$�S��k�J�X��I�Y�İ�$7o���_f�l��{ۖ��f�Z������F�R	�$J񫉻gv�N^��ƑWO����(��%�ٺ�8�C9�S%5�.i�tY(�t�вA�!>�k�vv�
\�V��oNY��v�#���9�n�	��ڦ���r��X�j;��b�l�pJ�NЦq�g	�se�a�Ə�Z��C�i0m����5����v9yf�����c�	0��v]{j%.�}2���X\皙��ɜq2���F����cT�$@v�H[��5Ʈ,��M�+���!0�:v�]r�������V��� ��6쉳�s3um5v�l h{g�)=]�6���,lP�Yu����ˡ�������1蟥�6�����x�$���3��4,�0��?m��ng·�oս�-��H�j���A���LP�R�-Q({Q�� [1DbB�qZ6t�k�X6G����C~ż��r����t���kݗ��~ޙ6Q��?z�6+����#��̍"3ۦ��Fz=�~=�Q��N���v��j�1!`�	r	$���x�>"�#��Ɋ�4�l��8f���b�p ѭ��iI������H�,�?iO�q߯��Z��c��Q�>�[d�ӑ98cJD�U��+ʏ;���G�w#}�c�D,q�=޶(`,$$�*�v����;��h{<�#D26�<�Y�?F�:�u��;j+��9��Q��D`s�8�� 䂰�@�4���W<~�D3&��8o"w�@֍��9~�~��\�iz%�B���B�� �R
B���۞�QKfmx��R�bҷ�*N����f��Ђ8�xs3M(�Y�:HA��Na��c�#Tsp����-H7nѨ"0��~Y�vE�b�ކ�������O}��9���6+��Q68��>wz,Tu_��Fo����Zz�0|D��񮑽T{�_.-$�����($�G&/K!V(�k�"�o�_����Ӻ��/�e��	����륗���F�R���e�ǽ����pڹ6���E]3����35��Gg�~�[����b�f�Q^���fG�)ٱ>\t��C����{5io=]�������!�!T�-}E��E�����{���z,�P	&su�����{��rV�V�N(��5��C��J��g���deP��G=�*�8��>�L�\���(��*
i�CO6�Z��b��B�[�xӻ�~����VMX�<h�dY�o���ȓ�i����x�x�}o/Ei'��Ut�t����ӄ���RC\��-s~��C�$M%��mņIFh_Q����V�����Y�_Rq㖃k�^���2(w>�����2�~�5��|�`�Fg���D��B���c�8��ӷn-���&GL�K�4*b)i{]�+���\���\q�Ś��?CD�_Q}^��K�\����ڼvf�U�!&�i�-�~6"���{T��9HA�/P��qVK_v�
	b����QD��m&<�E|�S'�z\�$jW�g���ʉY�*�*~��^1�/!��'��_/S�2D�ͱ��_�횳�8�r����*�a�Y@���e}$���ж�3�)i�K���D�0�2Y�����U����?_!6���g��w�f�8�9�s\����Ui�o]"���=�kWnX�hX���V4LӢ���/sc���t��TA�������d�=Tv�5�g�Кy��R�(��'�ɮ�y�"���b�Ǌ$��@��u�����"$�#�;�Y�/�iy�]���Dכ�>"H�A�#۷qC���*���Ѳ�<�@Ï�F�$x-�/Da�[�F��j��#E�gyz��ѲZ��FY��t:B�荔�6{��_�ӕDAMA����)#��+�����^(,��0=��:����g�#��8�����?W��[��1-��c�x��T��%�256�'V1H%��N�ؑv�^z]�#۶L.�]5�,�mreA,���
H�Β~�M�{,���γc�%R�N���}�40��(�Ĉ��15g��D}`��������'����3�4���Z~���I�.*"�I�#�U��,�G��(Q�U�������&Pގ�T1���?]���E
,����~��ٯJm Iq�_i�bpaYc^LD$��BR��A*$�͡ؾM�����h�k��Z�����g�Y�|�"f�&��u銃^|���:l���f����}���Y��aR8�d�NI$jō<��g��Q�:8���׺���;�Y�=^xh^8�Ζp�*3�f�pb@ӳ�#12���\z�1�\x ��1ý�m(Q��̝�U���o�0�^I�DG}Z�a��˄+�7*�������]�Ir�����ҳ}����j�>#�<�����_�B7"�q)
fʯ�"���6H��j�mM ���t(�^z{67�J���a�!�@�
G�=�'fw%]�����$���\�P�P޷g"l��r�T�;J�,(@:�Id��L�8���CǩCWD��������r� ܅խP7Ctq{. ɼA3�9�ݒrr��҆�ԅo��P�L���I��v{�X;�BǺ vfB3R#|��|�mW��ˆ�O��C�}�&ʐL�1�xG�G���#�a�Mg�!P�k�gX����"\AΚ�_̉#�>�{P���2G�2pP�A�EZ'ۆ�;�V�����O��x�����R
D�*�"f&DXgI��>]�����̴Ş8b�X�t�l��?j�`0լ�v���%�7hq�(5��������L"�}�ur��3��JhJ.vP��<b�Ƥ	���>"�#��u.<],�ೠ���cL�T�����=��5�p�x�8�E��[A�0�!�NMf�S5^�9��׳ʰ�#��O�׎����z"6ʁ�����H�-��	����_6�آ�3N$�7�� �x�8#2�*�f�2x�Ã"q���~��$#��ZYDe[�Rm����(�8D�>�D��ʨzҊ��ɶ�Cz�50zJ�ۼ��y�U�>�ˎ�J*�qGv_o9$�SlqMQ�"��Z< z�4fZ����z���Wr0M�ݘt��sw���oT��x%u�f^uk��^��E�9c9��1%�����8�A_)���q����n�6�˲su�m_gxح�pw(	�^�q(��;ԜKh�M_Z�2�ễ�g�;����b�
�I��?�7��GI���e'�WMP��Oj��0�Kui=Y��
n����^R4��0�L��*��9}n��t��Wf%Ɲ^��f��A���ݱ#WRΰ��u���;w��HǕMa��0�s���U��]�k��U��cdK��q9��uP��ٽz#C��7�S3�Y�!�Q��YP���5]M���\3\��H7���{Q[�θ��Śe�2U�;ǎ������ަ�"�r#���8q=D�.�h,E�%6r�f�">�/�;ŜȊ����܅�u���,eJ��[��ݙ2Ν���)>媝����[7������:���V�Ͱ^�6eX�ғu�7o����=�ӱ�?���:<�jx�R�xh�:Z���"��粖2xvo:ޮ�έ�Ũ�ֱ��ɹm�r�� �:��4��[����*����o7UMXi)�;Ý��E\=���J��B,�4��YH�CC�jIW$8�J���a�;.r��ƞ�-a�#�������Z��V2!h���JS��loe��:Bv��W>��μ�9f��i�w1_�׀8*��bC穽��fmqD�n0�9�����=J1�[kJl�jVWX�T�QR���֗�-R�N���6�w��/>�ø�6�!KM/�BͶ�ld\��!����v5�g#;\�hT����\�a(
��LB��iu�Y/���0�q�J״�Y�tn}����1K&%�����ZXC�љ�7\u����xe�������.�������]��7k�gs웝r�&�U9�^��kE�nB.�3u�B޲�J���2]J�-��X6vx����!�s6�f�����-���i#�K���J�u�)	K�&�2Ve%�%���ո�=8�`{sDxF���=c�����3�%y��0�Y��M-0)F,U]��ի�!�uX"8]�
8^��@�m9���S�V:#��y�P:��^Y�*몶^ D��V���"����7sŌz3��ζ��i���]n�m�N�v��)7F��i6�p��d��ط�ͥ���k��Kq�7;��U3��n�8:֔|��=E���ؑ
5%b[�є!Z2��n��Y�y�q��y�pj��˃j�U�q�\+@�`��]�Z�okʩn��qa�9��]1��2:�Ilgx���Z�5�[\�v��Y�:�!��jv��ι<�t�+�AM3u�d��C��+����6��c50��]e�%�֏.�ٷ��u�@��%�mq�R�uc�<��9�YGf.��m�g�ZO$b+��u�Z��[�����v��Li��H��b��&cR����o:ܶA]����6�#�	����5K�m�%�f�.J�`�2�� X��{u$�nњu����s��Pf-�-���,�7���6��r)a��K����6�e�1�N��eXJ�����R�ŷn�d�0�;b6�J��l&  hʨK����&��Iڞ��sL�#̀�\<�z�t��؛����1+�v��:���#�.xc���]��s�-����W�d�K���W���D�L�y���B��*8����U�ӵ��\��P�:{||o�F�WlR�0�Ʒ����Ļ��,����`i��E��N �q:�܎ۇ�t��B����i͸�^�q\�-4vt��\�c[֖@���C^pmh.�9n�w�����f�.�nio[���^n:mu���q�AV�Ӥ��g=���=Q[������\vy�W�i�jE�]u��͝�g��6�R�P�I�vc;�Zy�n���9��j魕�a.t!Eƚ|F��^���8������.wa��s͑��)�Ak�^N�#څ����lE��Y�����u�_p"���5h{o6(V۵�]:;�y5��cR;�5�:�����秛�-Dbp�D��fe*e��$#�7P�U����<��<�L?@�]h^��@���v:Q�Q�|hm�jN�L!��V��<�f�������������!HRTe'�X�G��ixy��<~�m:�(��v���F�n���Q��|C�n�A��x��p�z������܆�vMv���T��q}B���Q �a���*C�4�ie�����EHJ��:O�����M�G	4}��"��9��g��r�w�X��B�#�Pv}�)g.����뼟K�X�<J#P}�P�H��({�D[-BKMb��Mj�O:����>�jƚ��(�!���M���j�ײ�1�"-��a���L�8�/r�d�c�"mW�Chn�),?C���I� ��EuM���m����x��lލ#���5μư����6�a6���ƚ/b"Dh慓��/��}�����~��'��{�6�~���6#����>����ە�]>)D[�Y�+�?Un5pޮ;P"�F�t���I#E�
fb�7ɵX������熰�J�������+)�@��t��\������ȝ�]�EŚ%t�A�m�L"��٦�iߏ��e\j�\��+Z>y�<6Pu���L��y�bş{�!�đ�ڳ�ǂ({��-�@I��z�����}�O�mi��N��Q���a��M���J0ա5i����\���VQFȁ^�܅c+`q8�z�r~>�z�xc�ug��x�Ə��Bq}U��Pp���v��,�#/:>�DLeFᑆ�{�g����e>��D��<"��#��k�\�����(Z]�a�����\]�O�(Q:�&�u�F�#gz+H�,6y���t�}]O���D�#���PޡD���g�ߝr��|[��r��z�=���p�]Ѡc��]�2�#^�����T� ρ�5�+i��¡|�x�hd%�H|���_b�dH��������c+�ڔ/cB�5;aٔ�:��p�Ԅ2���뜾�ֱ�
��y^XT��ٓ�7:A~��ڊ����Otx�o����_B{"�$�&T�g�aP��Z�t�-��v8B���<��(��휟+:{�&�f��
d�8"q8h[A�-�f��xHn.+��V�����p����Eb5��
ƃ�I���L����Yh�kb�;o:+s�aA�R�5���$��~�+_���"
�I��$��fG��K���ƾ��5���S��{�U���dT���UCRu�u.蹎g�zi�F!�s/"���\��F��h��=�x�LG�QS��K��y�q�SI�K~d,HN��m�G�M]�=��-~|�	�[>�҃�q�Ty�n>�
� S���f���O�Y�����2���yU���M��r�mxJ�5�y}x�#��K�(i��Q�2!� �>F�~�3~�;������i���/S`�w��*7#q9	M�|鄞w���X_�ܙ�p`ά�*,��~�q�*��)櫲5�$��a�t�\~ց#ԷP��j��C�w!���󓶢�}�(452�^�răy�K/"����qIv�
N5� �E��]���T��\\������d@��aB}�b�ob�G�ΡƸ��dN�1C�_Q�Qܾ�y!��ES�ܧ�v�FhB7#�EU�>k�S�B����]w�(11D��T,�P��C��QX&�\��ئ�h���B���UY�D"گ���u~�P�wLi�4=���\�P7�m�i��4:|R]<lo�zc�F
��Q�]�ԏذ��d�!~~��Y�4$��^�dι��㡜�ERJb.�ݥ��XY� ɤ8����ɫ��~�(���޿4y)P��L��_<_���6�1`���(����k��~�BZc���5t� �قQ���1c�� }��+�w���w�'s4eU�ϣۘ���o)#O/�k�����|�K6_Q�H8˛["咭�fnX����\޲R�������qL�"���G�u|�]Y%�Z��Xl��z{�+�/6�><p��ϢŖ�:~�C�U�ޘ�ۊ��rV��:Y�3c�ߟ��O���O�!�����Z�p2����p�A�k��~����L9��\�2˴jJ�K6X�5N#�e��1��Z��R[U��=��v$��S
$1ľ�iZDG��.�<��-,�CΣ��>��.�n`a�D����������}2�QdN/T6�����h,G1���~�(@��
"�#83˖GNϝ��.�Ϻ��6����%:�)}1^�ƍ��T/quD�#����(A�B����N>����\xfm[��?�z=hu��>��8RjF�m:�Nִy��;�>��hx� �!��r�(.�E27�IeN������~�#�;�k
����
#X��>�\���q���<<y�Ȑ08�nCqP�	��]�7>8!N� �w���/�٩I�f��"(�?]���|�
9w->��p"&ϳ�s�+�O�=zǍ��B���Ė�*D�P��nF}�!�q�!�I�_���t#5���FU����m��+��!�AY�HW_{U��몁�A�DS�i�+��A��#������A�.������U[�^�w�N�LRPo\��GԐ�]t:�-�g	��cw�i�j�#T뻹��}']n������ԄD���.��9����E��M�#�6��l=nǐ�6W�m�.�Q��'�q�r;�;�Фb(��J��v�Ofڱ�Z����^-��E�2���1�&�gQ��0ggT��լZ�4� ��"�%�3�r<q�8C��jIXZ�Ңd�%�:���t��)��`	���Q���nϙ�Gr�v� ��R1Ziu��P�b:䍳8)>p�|;��T�d-[�:�����F���[�d�7m+N�K��h���D�RHg���?� ��V�w���|k�Y��zhi�C���:o"&`����(F���繪Bψ<����v�U�GN��(����(S��[a���Ǐ��D3�i�Y��ߵV�:��b�?+�~�}y[�m?y����lYM��:�bZB+<�ł��c�2Ʌ���<򯯒6��҄�x�L�D=�x�D$�8"qH/��WL���=��۟;缱$x��7߲G������.ߣ��с��r|M�Of����x}7��u�؂/)�]!��6S-"�l�����g��,2oM�����+�zNl!���b�{���o?l�p���衧����&����" u��ae���Z��3�WKX�LD
��RDhi�d�)�P���:��}�G瞯W/�.F�E�uP澛q���熄��f���f�$O���=�A�<C�#����܄!�+�o�|	RDĕqGwb�7U�;[mmiW�ۓ������<��6z`�ʐ�jE&7|G��ȴ��fF�����q2+ޏ�Z���mX��������sf�}�P�(]x����(% ���c�΁��AĎ�	чs#�Z�F�,����h���@d+�5�inVA<�hA4-`�K���/��UF����J-�һ_V�-���F�v�xM�H����P��-�g���3Wɺz_�^~����7%P�_Q�'���q���q�C����w��@��v@���	^4ٓ�b�~�h}BqF"q�q_=�����H���g�*��2�$�Gͩ�������@�|���./�yV#gˌ��%ߛT#�>���y
:F{ۆ�ƙ]q���<�����DmF�`�ԍ��D"�n#���C�m�+�N(��nDb�=qz(m��*�Y�S��!�������Ї�5��m�8;Ͼ�z¡��0�9����x�"��Ƣ)�Q8�H8����,��~�C��[VI��I`�w�Ue��Gwޑ�y�	&Ѕ��*Ɵ�,B'P�G�~j�4s�#���+��}��ݫ�V
7�� fW'��!�\\�S<8�k۝��������On��cI��Ĵ$����~�׌�z �3�џ6��󎁆��TE�B�Ϸ���XCj�u��]�����F�\��:F�f9}�޵T# ��u��<�zjt�A��1��i��e�ԇ0�ya����xd�"O*�\_-��an�����ch�z<�Pϋ��Pp�����Rz(i��,��i����诳������F�H�����Ir��}뀨K*2�f w��������y鿙8��;��jx���5B����*6�ќ�����V�H���W�R )aj���R�Ֆ�u?gb���u��jP�bI'>(b�:Eha�5�lM�c~�R�}(��:^�Xt����{����Qށ�����
>���U����w u4�͠�"��$�P�*%_��*?C>M�NzG?"�}����Qhi�����E�4�Iҏ0t���=�,q����H�c7�Z|A]���<������Y�;��i��$z��!Rf#qX������Da3���r5q�G�Db���N.��)w*�_Q-w��H>��<x�z���zث,�#�E��h��8�_Ƽ��ԯO�����B�q�(�F���;Eru��7�P"�;�Ѱ]��gMQ��FS� ���#�P�>�f������3�b����k��@�;��(:}sۭU`�����-���@B8x��"�K�_޼5�I�cֹ�0�?��!�(MȓI��#����<h��>�^F��W.��x�?/K�Ϛ��6�%��.�J��1��lPp��L�Fb��y��:~�!��9���ҁ���=_wb�7!� Q�ᡧ���~b�׹������_Y�K�xk�X�p�G������h/'�j�SYc��Y:�Ř�������KZ��?]ϭjɂbApD�]� ��[:��O#��'���DP�����~lA�f��������x��� Wy頋! ����dip�T�n2-{���54[��I��nW�����z��h���r���*i�\ڸ���n!@N�ر�l�_��o�?E!�w���{��S%"i�8w�u~��gH{�aPg�#H�7k^u�=ތ����s����B�����z�4P�u`�><����o�>�)��{Q<h�w��g�5�!���	e��F	�6�@ؠ���9�^ݺC���n.y���T�N�D�a7$�tY����i��>���k�C��-�(�N{[M�7�#�{��w��l��;C֭ �>�^��T�b\ءg��
ϊ	���4�U�9�g�z����ؠ�e���Ī5&:��蒣c�.
C��(3� i��f�]��6/�BZ�!]禽��������o�J�adNz�r$�j&�D��X,�4j��a/�~�c�rt��75D&E{�ePM}&w�4;�7�Ч��A�d�[�Q'���CH髽��t���`C��F�2@������j��w���Gky���S��/��D]禾>��I�t�~��}�ü���ENһz�@������f��-1Hidʬ_zM/�LJ� �ԍ�����,�v�g�/��t��"���V/h��؍ּ�P}C��:D�(���ݕk�Y��B��V�w�P�kB@��gey��}��i�C1fU��|�9Z,=�#e$[�!��ԾT9Sb��a&��Hgl�n�죮�{�wW��-4�Aq������yW�o����8^������a�pZ�`U�p>3�Z�����3��9���JE���6ݥ)�ѧN��%�sl�զ�'<�t���,�͊�V�;�i�5��rv�˶E�,�A�E`�ۃ�N�p���R���OBi�q�e�M��p� b��eLc:��3V�m��K�I��1�!��L�k	m˵*0XP���i�͛�3�b����)ے���v�\�n��[��U���냲mF�I8P�H}�$����ܯ�# _gcT,�&��\I �2���5�>�G����"�Ӓ�S�y��Ј���|4�]�$*�h=��V��<GM��*��Ӕ`'0��r> �����N�jՔG���I|��O��b!�b<��ՄmК���&[�_c	y��a��L��=_z^⣓��}k����p�A���^j����0��l��p��ު�P�q$�s�ܪ�hYk�d���~�_?��Q��n}Qy�������a���ݱ�S��"�}J��;�|f�OD�1!�| ��"9��tք7^������=�7��yQ��I��n�05|�D-"�6�{ۆ�KZ�%���bۛ"j�^N��Q�H��eF�Շ~v���X�"[((��0ǙVr�3� Ρ&���i�@�B�F�̲D���]����$���M�0Eg�Dй͐�j�Dm��H>��#ǁT�:����ٞ��!xyɚ�<���R[�n9��e	�!ϱv5<-�pG=,�v:�ñ�0�J�6�k�nIћ,~�������~J`�ƈ��鯵�2~愖Fz�%P�~������}�A;���4.J�+x�m29�2����(����$A<�G�م�p@��2�
I\������޼�ӆ�՛������M�������i�#���5�0K.�:r��s:9�^CWv.��:�r�fR»�(�X1�^-�l%IԽ�F"�A��C�<u�����k��q�(�BΑ�b���N ���~��v�. z�Z�S�������$�7w���p6�M�
�7"�d3�Xr��;�(i�Ѝ$]��E���Z�E_���c}�A����2�k�㵸��:G�}��b*�����-#��������r8hY��c��{����32|oF�j����B���� ��1��B��U��	*n�w*��,���bn�W��Ę��Cs�sY2!����ԟ���h�>$�D�-����!�CŃ�q#�;�sZjx�?]�'�b�}���(���
�|&�=Π��#g��~zk�D�B�ދ�������p�hx��������A��<Pŗ1u�%kn @��l%r�Nƻk����^ݥ�U����U��j��M�}�>j����{}
1�H��H��XK�d���	?7�7W޷�P�w�n����Ć�_3�6ײh��1�j��	?un���5$1��rGΜ<�U�n@��s60�56=� �������R%zh٢:���L��*��q��+��h[E�Gl�<Fm�>���K?j#=ש �1���3}k�8�7$nۑ�4�B��n���{#��T��cH��H���M��8gH��
�/��Sw��{&�2�	�/q�·x"�úy������e��n� ��
9@dU��Gv�K���mL\|��%m����`X:zAY?n��͹��ɼ�:�4��X����B;2�:��غ�+͖z��Z�ZU�,�p�)Mg��t�����2ؔu�b���(��T��n��ihLR��4�3�]nQD쿸��T���z)��o/F��u7߷���K�f�����;]'_l�ΥƹBu�6v��#���ܵ�,S�\9ֆ\�X]Gz�N�^��ֻ�C�s;pC��	���i,������:j��L㓒����PH�WI�3�1K,�_ж�e�4�f�P�����ޑ��T�
��.�cs���n�N$�Vr�V4B�9��$�S+V�ĥ�۳�J���� W
�2\�E��W:I�`Cy��G��9H�j:�o��������t�H(��3&��,Ct]�h;)�*�օm��5��1@' ܸɤ�2�MfK���L����w���0Cnokc��'*��h�ׯBˡ�7weAhK�8}������6�eՋ�0��r���=X�{�lv0�۔���ݏn̻�z�ɨ�s\�Q`�.ܗ�&4�Ʀ^r4�ť;�b��zN*�n�F���yP�ˆX���!̊X��k�4�}��e��#e�'gMm���5x����m0�8�8�+�{]����r��R���+)9[�!R��B+� dt��t�:EB�?��4�����3o\�d
���V����=J��">��8aDR4�(���������-���r��SE�^��;���Tu}w�au���P�X1��,�5=�lV�I�G�Y�Z
�Y����e�?m�?Y��
�@BB�i�n9+��Q��ц����]�C�w:����}�:�5��5˯��6W��d�հ=�T�c�%�1K��y�$�Cm
,���ML,0��О��e|P�+C2�6�R��f��l�����#q�i2�k���E�i�=��nY�5$^�M�J$�!,g�G\���r0�3���*2��7���C���Ʊ;8}ޕJ"ȧ��u�C���=>��Pʢ��"z�Q�[��I���Y�d��G�S��ƛ���lgŊ�Ox���|�Ś��nH����#y��*���R#%�,ΡS���s�3���P?x7���A�q|��m���<A���GHF�j���zG����ayx������3���6<<�����X+���g�x���nΟ6n؁����^b�i���ӤF;��*fJ%FRQ8k�򓭞wre�\ꕡ��G��Ev�*Aʽ�8����:����}�N��E��Nm���~ܸ�~�y�.>WN�z�׮�0����`s����"�k58"W�R�rXg9�V��Mt1	/_$Π��Ce�z�YW}T����ODϳ�g��f��4(�ȳ��?ZxDD�+���2��{��4�g1a���i�t�ʏ��4�*��.P��o�uP�_M����H��<7�hm!���Y��*�sYG�񌨃��
s�{���~�ޝ6b!4�+�ٚ�k�H��K��h=�&2]Jp�W[۰���uC�2�M��N>��Zh�Ug
"���V�#.����c��%:=�&cfϚTuT��݆((��>^���F��6��<-���p���'�j�+MǤ�EHSLB`�Ŗ4���gO���>{���{���_�߬���~5�h�H���ʻ���������Ƞ�.䍐�r��G�ފ�	��,[��Z0�:C���0S&$�(�RI/��x�zBƞnW�ݝ0`hm��XF�@ǟ�M�,٢-���I�jI��T<~�C������\�P�+�-�<���b��Y�4�4[�X�2�4�ɿ�����OE��+��\�g���,��걶4�2�JjD]'�ޘ�e����Uo������%�<���>��(x}���H�%�#�����<�|ƞ}6�P����\�.�G����G��,���<�A��(@�(�!��ȭ!�'�w!�����/\�1��)곕�]��3N��ƹ3��}hK��v�K��8l�u,B`i8X�*Eڳ(��Jc{Y�d϶�8�#Uh[��Բ;��H�h�i�'t��zK�/�ǈe���������>�vTf�,14t��@R6��7a4��ݝ	�SR�6�+A�s��l�v+W<vrgs�Y�5/)η8��cD�̲���ub1U�b]�rA�����i�!�bb������S ��=`�	���.v#̼��-��j+r5F�QD��]��b2C���fĤ�ݗ,��6�v�:��.@�!�>^��M�N�m�ά�]����%v�u����$p�*�4��"�Q��12*P�M$��S0�ahg(��S�B����鱐Ch��H���6�YӤ����n��dq� r5$)C5�9���ch\�8Gb�eT�eE1���Q�C�{���|�Ϫ_�z+�|�ZDI��h+�1B��F��E{�3}���1t�m	�A���,�����~��d�9!M� �'2�!j����w�N}f	6B����v�z�>��8sQ�^]���(N��C��
3�l��.Nۨ{��RcH�����)$G"r�q�7�|��v�~ͻ>��c��wW��-P�:Fˏ������>������V���Lt��z�?Ddzb;��s�ƾ� ����g	#�`JH�2D�iȬY�#ut�dKW�"��̟�cޑ�1�R�ZNSӺ�"��"Rz��4/o�⇼�d�@�0���b�����*!�1B�S�>�uGu�|��\u��l=;[E�r�&�)��pcN�@��2vC�9{V*㉩y�&̟$M�q��g
l�"u2 ���f��BHe�l���*fT[��1�{�_z�����8���?20�99�Ƈ��D�ʑ�%��4��B͗��������"C�c���\m�[IY�{�6mn큢����iu,�F�)�bwe��s'G:`���yZ�2i.���Qb.DӼ��~v��duC�C����:��4�~���"i��|o��V�H�W��k»Qc��#�#&�$����^$�f���!��T=�q"��z>��W��k�Y�&�1;w*zvq`�C����G�(igN���tS,��CmҪ�;�p����X|D��d�#O�[��.K`�83����I���@ѽD���P���1����n�D����lr·��UH���Ǐ4���X���0�)(�5��"i��>Ϧ:åRF��:������3Ր��Z�~��À�万j�!��C6�垞��ZB���V��7-��<��,���)�>�P1�@�a��˫w�s�3�y���]�����l��]AѡM'#(�D2#p�YB�r�>��o�6d��ٳ�C����i�P��+~��ݦ�Eѵ�7cY�'j>V�b�z!�Y�(A�0���00�1)sM/��͏��m�}�|hi�^�>���TSH|й�.��J���P�!��;�vha�-#sѤ/{���D-����{V��$��f�ጒ���\J���#�DW�a��K;j�N�*ϻձVH]������U̛�
�c��T;s�R4ɩ�D�hV����*��0���f���
�M	�������*-��r#H��t^s�1^��}�L_f��ȓ��L��(�w��$�x���!�]�n2R�q��(��ս�(�w8�{�Q�u|lx�&H澺C���_h"�$Y�T���T4�b"��[SZ|N��VG�����<>��R��H�)��H�ij�4�,��MYD���f^�F�v��g�4Y��x���3@��H���ZB�A��4_V\BkH���W�*<-r��#pr��q	<��N^�u��zl�\E̻X��ݙ�b���"WG���ܔM�������(��ڵC5+B�m}�j�z�W4�Dŧ����@�>5������9��Dc�����G�>�4��_������B�RA4F�>6EU��%�~S8w��祬>=Œr�2Fe�4/PFM���A�yᡥ�4fdY���j���}B,_��2b�dT�h�w��s
T&�i(c��Ӧ�iiD3�}�:6D���F{��_b�|_�3=|{b�="�I�C�|,20�e���ȧ7�5��C="��e�����˅�)�;���Q����P�W�V���O���SRt�hY2���*.>��l3�`C���|ȃ��/� k8���TU
�0���v)�^��S=�"�wa�2�H^���o a��7Z�>����v�^�����5*��~��>����7z�.�2�����9
M�/�Wʏ7�(���2�P��D<�M[�;#�����홡	�?x�?w�,�!�#R�#���Q�Rf�|�ӤF�����|�F���b�Sh9lZ�k�4f�8qJ�Aa��^���.ɸ��1(�2���+�J�dg�ػ�꣺	Ф^^�'mۜ�D��I�5�f�����&dl1�^vjH��j۞;>`��F2g;�c��M����B��o�:u�鉪�k����B� ��K�ڵm����!���V�ǀ�=��?	r�.%�m�ގ�-���<2��&��BŠl BHlr��c4o,l@i#8��d��˺y���՟vOqg5٥\vK+�t�7^^}ٍ��l:�������>6�<�C}"h�6����Aᢀ����_b�z��^~�ǃV��^���q���O޷G��5Kq�|w*�ܩ���6Ns��v�I�9���F5�U
�� A:-��a;��`=YK� �i��3�7z���=,� _�k��l��痱\lMY�2)��س�]��̰�&��̺���Y�F�fv@v�@{�|�Yݐ������7[gjLh��lV�D�w;�8����t� �����v�k�����{���8�,�خ·�9�j��O�=��]�k=��1!�%�v���砨|���V� ֫`������-��F��GN*|�����-]�ΰ��U7<�Vt���h�l���͟1q�������3+�C;���������'7��|ٽt<�%!&�R��V�*ڰ�����-@����3�͙�c��p+
~��J�m7�GU^Q��蒆�q?O^gh�bj�`��&��mB�l��,��S�x���T�sPg�:�U�i0��׻���x��~~�;���Wܱ���Q�ːaJ�:f�VcŴ�$�{�味����v��~'�:�9��|��Lot������z5���E
ȏ��D�"'@�Ky�gy���������~�����+��Y{s�)\��b��{/�C�"RiH�!�p6��"�f��iQ�YU\��f&��6����bu-���tT-5$l��+q�=�R������词�Jʻ�o�^�^!��$C��zy�v��q3$/��L�$�6(�6�EZ�����9��|�tB�{B���@br1�h[J����ے���s0�k �1���X�6�Mf֪�>��BB�r��V�-���u&'��������l:S�o����G�p����3���@a�@�.���	��m��~d��|qRI�г�Tu'u�F.��=�+�*d7��&��5�u�� 9���	��M��wL%�yz�'��蛛fvx�)���IQǅM��Ԗ}���9��-��c�B�J}vh.�,�P�������kF�\�ݔw��1���[~�B����/ye�ˑJ�#o��x�j6��m�|��a�n#q�g�t�YS�@��E.���Qt���'��".7��r{7�}a[�����M�x��«��W�+k�S(�-�ϫ��SתQ�O'�ޒ0�[�������|w�0Vt��ӸXw�9�`�.j�\Y�Mi�Þ����3䲑YA��U˷��*~�H�qƃ2OI�s~�jڵ�	�,�5qg����|�ӣw�(��u�q�P%M����qYIpOb̔v�ad���Dj�E�N�+r�v���s��vH�~�7�;��KcJ!��� ��V��a0���G��t̑�{5�]�d�y���֊����/ *�ޓc֞�h`��h�o�ky]�<*`���EBX��!�Ś��˵�pt;,^�>��:�_)q�`/[<0T���vG\PN��I�ᏹ����P�(�Vomvew<�n|�T�ۆ'����uv���v��ڸMCS��6�ua�@������7~~~���d-���k�$��nr�V�U"�g������֫�ªy"	|���ֆ	F｛"jIƘD���b6}=�xg�u�=��=�<�������eQ't�.m1���ʂz����$�ݔDm"H-�o��Y��>�?.��s��P����O�s�� =��L�g�yU����:�:aPți>E$�P���Ј�ɾ��n�j(�>��0�I������&`~��m��]���&^���K+���u��17�w��4
���%q���w(��i� �Md��4T�ս�M�[�w���y�C)�T��PD�(8�B7�:�
=�3z���f��58������nzK�$��Ĵ�w�Iz[�'RW]ʽ�M�]v�	mH�b��CU����K�#����ٺ�.�{[�f�Wa�r�d�t���^���R��o6��w�na�뾵������ok��l����z\�MH�)H���;���&��7t�_wo�MRעb�.��7��Іx����3+�������RH�A�T1�q`��_�a�/+�}4L��']������xt�ʂ����L�a����Tl$(��"�C�94s�Y71�q�y�q��O�8W��F���ڲ�J�<�l��\�sO�7"6nZ��=���X<�!%�ԍ%��;^�c�n/V����?G�����=am����.��=s�!;����n��S� o	^��[ÕD��/��n�Z��n�c�N�J�N��N9}ײAS�K6M�E�X�6�[��Z0�n���فu�]y@*�Z���U�`F�C���oH.g��J�'�Η�����gbhW�/8�U.��ᢇ�1+�7t>Yg:�U�fv ��u�.��'�^�-Π�i�O� )L�j[ܯn\��$a�l���(N���!���x��"��ͼ�ƞݻt:�I�Axl�*f�������ݝ2�0Q�`u�Å�>��U*��\6����<�9���ǲŭ�Mu�ⷵg=�Y����U83S�U��lS�$�캕*�"��N���*>wt+l�b����m�[r6^
�W�u�BW]1H�*)���X�
o˔�v�ئ�Ρ�#}�s7i/C3��N*���QeZ@b��Z�Ÿ+]N�xbR��WV ���0���|q�&�Ƞ����vE�\C���|2އi�g�e
�^��9q�an��q���
݋��O�։vI�}6���6�|�����ob�p��Y8.�ܬ ����/��@kҷF�d]D#Ю	jl���c�ie��G,�ln]�);��+��yor�9��!}���c8	np�Mcb���kB�]�P�������}P��ɧ�M��f�k�����ӗd�3x�h
@gT4Fn8�TR	�yh��8�eAs6�-<���øqө:��\�/I�L"^.E�0�yo�m]wbR�w:¡����`�ک�h��M�܏�l�Lglh)G=����y�]�&�r)2J���,�cY���mсGZ���R�|ė];�G$�B��0�������ٰJ������ki�Xg�R�rvG9�ŮװN�,5���\�w��z��շC�c%��v�7�˕�5�iM�z��9�U�z�ۄ;m7f"ƅf�B�
�B8,�l˲k��V�)�Ȥt;0H�۵r/.�s$J�L��8����;E�j�rF�₌�Ͷ�.�g�i�:}8z9��/��jTie.��g�Z��1���u׈3F%�S*�.m�C�,�s��㓷�
���T���ϝq^�-��{�՘�A���5�j,�f�&��)�W;��3�v��\�&�(�a��5[�f*Jp�F1��<��LC�f�F����j"����y��n��>H纓	�������*��]���|��9Z�%�f[, Ypa�R:�s�8��F�ź����nCQ�';k  ҈�7�1�n�n�f��$��	6K����V�A�jl늬x�,,0�i�&����;v8��g���ؚi����;5�X2�.΀�	KsH�F$�Y�R;i�Cc�������h_Qۣuچ8z�V�<5����m�0ݺW��a���m��2p��v��T�kX��۳���&��H�;9�^�1�q<x��cbz� Wn�tE#��w=��[�R��g�da-����;��[�M�6�z�'>�!3p���A4�9hf{���O-�p�8�-7m�T�v{&X-M���r>��κ�:�mZ]Ak�S˅�n�]�D�5B�73Vմj��V��0�c
��o:�hY�(lkt�����GolF��5�c�K�nLq�b�e��g�I�/]��Y��4ٻd^�)���P�U�Tu�]iG2�5+,$@Z�P���<��C�f�.�3T-q��ft��Gk΅N�\
�țm6&�a�qV��s�:�۬���8� m@���hK�ڴ��n&1��K�f���`pl��@J�¼<&�wj[�^�gF)Ra� ��u��IZ60c�����#.]e�4�I���{��K�Evr��{\��5��8�uSغ���U�F8�ׅ:pb�t��Շmvqg�>�[�eڭ��8�km��/.k����.���a`i�2<n
��2���6�g�-Ԛ�����T� � �-p�,9��QԈ�.��Ѯ9�z�\Q�2�Q��p�L�%�\�q��m��@Ʒ�s���Τ'<<��8�r.��	����`���Y;RG��t3j)����j[]���u�q�T���y(\��RA�(ܙ������,�J��O��WWZj�t#����J�l�}�=�g����9���ADd�&-�W��y�ٵ�J�	u��s$S�y. '�zj����{Y�҄�jL�����8m3�1
�f�����$V�ۙ�j޵���r�Y�<��*^5����=�6矂�,Hci ̒8�ӻ+M������:�9,�u#�J�-Ӯ͘��eD!�=���)�}�QB��_���~{���3wf�#�l���s���N�5mXt�����+�x�q�Y|��g�EFP�9!ŏ����er��=�ö���K��a7�Y�h���|��س;zj�F잤	]O���a�D�ٖ���͏{˴��o�lS{����*mm���[{��tͬ��S��X����t?
��ݼ+Q/t2KW�YQ�z��/o���P+�ZYW���Y]� �/h��G{�������6�.λfx�(Ʌ2��)L�gu8b�q�8�^�yi�5���s��6�=�
D��\���ZD��@��v>*�CBk������ݬ
4^�	�#���b�/k'y��1�����u�&>����a^�L�6x��i��2In���m6�k>ߴ��-|���e�w�I���X�^��C���>���%-��6��f#�9�w]��F�VV�YfԚ�!Jъ2����L���fn��Fa�W��m�y;��3Fyyn:����o�y<��0��x_���������b�!I-+D�@�K[����	��u9��������N�2�5՜�Qx�+�1�.�݄�����MBYI�x��wz{^{�9:��Qk˙j��`��@��������(Kn���V�2][=�w��g5�S%����5�Evsp�:y\+hh��To�tRuFn�v]��skռ��&ژ�<���8A� �*�C4�^c�P�"�l�q[嶟OgSqiq�y��nl)���BP5���}�v����Q@ZA�*�H�O���0þ���ٲ��l�Cg��jz���9_x�j�{����pSq���me��������:�PZ�A�,����/�zu��"�y�x�j�rsvqh��Z�JԤ��H�DΗ\�F\��k:�<!y�o&|�����'niU;Kٔ��#׾d$ٍ� !8�7f�~�۷��fMy{������Bjn��m�֫����|�N7���3x�̆�Q��"��D��G?c`glܳ��{�V<"׼w�����*̳q.�KnP?zL��۹}ǌ�yR�I�F�	$��3h�����r�2��l���Ư���x=��d���K�%�N�
�Yz��u�p"61�3��6��&���������k��7/�L��%͘*	�	�b��r�2W�7���G#4<��cH\�B�Q��IVz���U����D�s���-&њ��}��{G=HO,����
�2��y�$�y�f��ј �e.0���tg�D��������7���m������d��Q�wƗ����0�"���h�?[j`�d���G)J�����7p�9����,iyu��'�%�

2�!���G|��s{w�S���b)��%�9�<��>G���r��t��X�����X�:_�N�3Ȝ�[1�s�2��w���~;Rc2�ϒ�m_x6��F�罕h%��C�\@�������S&3N*��WG[`pB�z�TD��Rk��揳���t�ɽ-�CT����@�;Y3E^ݏd �OœQ��9�����{��c���]2rq�u�܉��G�Jlk7�WY�}�����e�y�Ū�PS�M]�h��W��f�
��[���!��	[]�r+�b`Hn�eH����ӈh�D�.����~����a��[��r=M���狷R�콚��kt���l^�&:���ru���0���ǡ1�����wk<������;<���{��ףڍ9���gQ��srr����v�����\�Lq읰Pz�9^V�:��y�$�����5nɧOVn^y*�vy�rlf��f��%�h0Ţ:Wu�[ڛ����_���i2�f��v�-a�;�������gmq��T��ݲB3(�b7n�n�u������:n^�^��]@�;�W����/�����Ϝ��~�1U�=?Eg\W~2�D����׷�������7X,�"|�M�>��_E}��?^	*W�?k���<d3%�:o �����{��*�� �r('#�Q$��sB�z;P��j�zy
k-�,X��~���������p���y����=;5F�
%I�aMǳ�2�W�2�ݔo�l�k��γ�2V;(��Z/���p�L9���U<6/z�����t��R8�&@dIĶɏf�wո4b7iJ�^�j����w�FlQ:>����YYHWq^�6�#g#�Sj&���n���OX8�R�'�O8mqɈ �s�V��M	Q��N�2G ��)Q��7l7@8=�s!X9S��kEeab���|}П�i��[��i�в2�M�%ۏ<מj�X�l�&)1��=������(����o(CH6U�Tf��p�x�#w:=�̹:�`�m��K�<���!����Xd�T�`:��B{	�]��jY0��+�	n)��Ȣ��������k	�ޣ�(%0f �7t	�7(8�W��X���}�1[�j���B���?Iix��`֔ȫY>º�a9B�nL�0)W���v�k�C.�W���]�gP�·���Q�,�ם=����.얼wi�?x�F%tJ)@�{�T��3�����Q?;�B�e�z&�ڏ��{qg���Ӟ����`�W�;ډ{0�̩jʆ
()�%�x�D��d�t=����q�U�v\�
A��E�!�&bp�!RO]�k�ⲍ�e�¢�~b,sGy����S���:�M��V�XR�^y�b���,�౗D�N?=�~��`M��wa��@�q�rc,��魻�Ӷ�Ua[]�܁F�����8�/J�1!B6��7"z8#�o+�緲Qڥ��]ױv�Ɛ�'��l�·L[�4�C�����rr�|�հVb�kZ�_q���)��8E�o�[��#<�D�ށ����yo�ך�2b���5�@W�&� ��HZC�nK������?w��@��\�geў�5�QF�ߘaKܛ�}�]Ӟ_f>,s�M��lia��x�(���OVS�OZ���{�w=Ef�b����.2��0<��4kSs��Y;"�9cb�^O�I�!�z�������8y$�n�c+�d���u�n,��46�`�q�͚6��c��l����x� �~��=��U�%*��;?0Q5�Jd����}6�<�ה#D���
%#����[�/}����|�u.�;�����:j��:*;w�꣏��S*�O���l8CQ7wṷ��>���z<���`��F]>�T��:n��ެ|L@c�mL[���0Q���A�J���Ӏ5�'Ӱ#⯱CVwO�-�w�hy;qÆp=%�Ӿ�ѽ�:ݻ��9�u�`p�$H��vn`�fض$ȵ����kz�����n�Yտ����,m������X�,�����R德4�M�#�7ewe\��Ǻd��a��m��gF����^��,��x��T��������W�e#�&�1�uWjf�7}'��yCV��)z��^��u�G��u����N8dI�dI���ts�l���w�==z7bk&��)�S�,��Z���ݎ�8"veh��VM��J��J�M�y��;����yW
�D�E�vd`eB��Dǝ����U�mu̿h��`�t�Y�Y�#1Đ��������ͷZ{|u���T�ޡ�LF�1��Ju{���Q��pZ~($Í!%H�;O7u�hyf�η���]�lY��֫aN�Z�uh���Pzv����Г����0���Q�J�b�s!���d�[�j98X���x��c�^:;���^*S��ݎ���װ
�w�b��sz��.��BVQH�lo�5�n��\h�\2t����GR�Q��*����4�I��xܭ6)��[l�4N�aah�bTl�%�kr]rMcy&m4�Fht�r���.��=��,����ٱ�n��JnVs���v����"��E���p���+]�&އCn�<��c�6�v㮠n�>L��ڷn�G=��u���]��2�s0Y�!�14�-4K�����������.�]�}�*!qn�YZ�p��.9���I1s�����`��
r,�P�<x�z�+ְ::��y��nb&������$'�M�tP13� g����r��Hfnd��'A�gW`{��ǽ55�C���oO�C^v��B���9[����C����q{;�-,��)��ϻh�w��+�t�t�x"�b�o�E#�=����fM����w�0Tj��P��BqM�o�T\�ޮ|U�v�p��OQ��&��$�F�#�o�vLr=�C���p��v�Rxx7n�-|rX��=�#�� �"3u�ِ�����^��'I���&Ya�Ȝ��[���>]�V+Pd��^���b}��}�On�،�_gj�h3i0+���j��H-&BQ�B�)�ÌFa�4q�Kt�Dxsi vNw�s̋y�6ܼp��.E*���y�X���nYR/,�]R�+s�6ɡ�"W�A�h���T��:y��k����`nY
�H"���}�_My�S���Z<h	�묜f��3�w�	(Ӫޫǡ�w�ݛPԓ��8��Wu���8��Ak��X�#��t�n�ScN�J�c�{�7�G7��ջ�bۋOX�1�zy�U�+�*+v��V��my������R���$ڛ"��c��P�cz:u8�J8��N�8��3{�s��i��]�ݾ�Cd`Q���M�F7l�X*�y�����<u��]+�\w��2���oܼz�܁Ff���ܵUU��[6~�^)��8Å���H������B�d��gޞ�{�}�����'~� *cq�\�����e��j�����PLtNt%��ޡ�Ɩ�Jc��n��.�p���c�5Iы*����8�u���~jmcl&o:N�0�ő�=���ʂ���J6�[Ƹawt�#�!�۬�紊�����p�8���{�9�3D�iz�yQ�~3��i��Pr��Xb�j�><��Gw���Y-���f���Zف1q7	�I��zjK���1��y1�����g��T�
�{�������[9z�I�G҃�B�O�]�r<��5��qo���ܗ�vz^�U�����e�Ⱦ�B�-å�3+PzX6^&��`�A�kT5^m̋v����/5��+7���ckN���`�b������;`��I'-�)��7��:����fC�#Z�#�c�4���GEZ��p���/�'�n����@�xl���;��oz���&¦ 5�<��xݘ��k���n�w�B|2���C}ԣ�)��?Z��� P�dPu/�[�v�,��[Fr��1x��`�1f�7�*PNB�L��ZYu35CDe)�ID��w-�u!f�Rm>��-M�KEm����	���`��h.��G5��XnMilJ\���>*��ش��<���7��ja�d���n������Bw6��ķ��l=B��c0|LFĽ'@�zӈeK�=��91I� (�*�-ܙ��Y�&r��P�9�jepy�"�y��E-�	=LSE�.d$Z+#Ien���;�����V���N'�!�}�LH�2��͖�;��y�X+^vp���3��E%&�3ע�n��H�p�:�Ô�Ka	Cȴ����>�yD�T�����HͲb���q��ù�񑯈�DS+�҆Xl��)��{�V��TT%�U�-���M��Ӛ{Խ�r���w)D�1���З��E���t�Έ%��*���k=K&*Z2{O�;F���MֳE���˒�6��n�ꑅ�;�K��cF��IK���5��T4QV,�*����v\��X�J	�<iZ�����>�f���ƥd�5�5�9��dC����D���.��i�S�y/��|�Ui{ޮ0.�@��@g��:��>��A%�|���B�-O��D<����H�q�nεm�OT��^�E5�XM^-�d�;C���AW<��[�M�¬�~v����׶��t����Taf/x�VE,ඖ�/��t�;��O�SNĈƤ��q^1~gס�̃RD��	K�8�٫�,~��Y)��Z��x�u��N��{��MC�C�	��(-LX��}�_�s�^Ŏ�zd����(��i��<��`n���׺�Uר�	�["H�w�V�y�˻3C>���b�g�}��~Gʘ�z�t|����y�(/<��.�VJ{Ζf�p_I�F��6n�ޚ�6�]9�'jfs��P���d6Iâ��E췆�������}}}��w*m{.�x{I�`�L��x�(�H1���|�0#�]wd2��;z͞�>��T���hzl�4���{�=IpY�MsX,����wW3����s�JgD��u�'u�,�ϧۓb��1�����U���K.�����m�4�y���{}�TVU9��01{�j��,~��"^����J�l����5���衵����F��LU��l�%'Nڞ���/o��ޑl�HE�{A�b4�HA���B���T����^�<��4�pk�@O�_���/^��x�_bu�S��"1@����mDTI�ÉL��=�Uz]8S���Ϻ�Z"��b'|����0��5�!�ze��n��7]�}�k�<I^	�cl�����G��u ���q���R�=�Y7;�p\��O�V�.��-��ݭ�W��r��Bk��Sx�_\���{$�6��-޺��=��ë4E�BkR�>��i�5.��R�0D��k��L�+nV��9��Bꡡ(���"	BP5�=q�ю���1Aq�.3-M;��g��g��\�n]��<���O^<ѓ��B�oA1��d����H{x�Z�FŇ&���ϣ5av��-�#6�VlB�k2Y���&�=w.Q5�h2��e�i��6"髍4�ip�7K�D�M1��v���9.: �n�T��9�[�vC]��`�S���hZ�s뺈�i׍��.u+�j�WYw�1�6,�Yc��iI`��A�����8{=Y��q����х�z�v�E�	����']c�$w}���$��[N��:�"��^�T7	�)u�U���7�N���cy4�R����:�՚��亸���䬵�h���C���)Od�:�����B\I��w=�}�kv�t��Q�cxU�O&׽��Г�� S"�}^���w/����ƌ4��HL�4ް]z��}��w�%!�s�N�|��9���!gUY��l�zdH��짏�E������$�Zb8���O�t�Y���r�>���/��\{�ʼ6�j�wt��*�C�6s#��Y#�
�u�$�wc��^�c0�	Fq���ۭ�q̌nzz���1%BX�g�&�R���Y�e��c��#p��0�=��KױmX��{. -�N��OXu��ù������ �����#�d�6�MɹT�v�c�c�ž�ǧxa��9���7r� ���r�bq�l��%��pR�)7Bب�T�f'x:�uå�D�ѵ���n\�0#��5�8Uzy=����Gd^��K�oh~���<n�,��������i�GZe�yeq�C���ÔkU!DL52��^����w�,�^��b.gD'��40E��s|��1��ڽ*����i���z���o�0<���W,���x`{��/�0%l�#q����^_�ͼ�jG����|r�@+��^?V�/b�e �C��9r���`�ٹYJVz��m��ki�\ƈ�Omu��qa�kh�D�68��v�c5�z4��=�kp�bܬ�~�gr2���F,weꡡsI�{"���i�/꺕4>�p�ӆIjүVg�
&�Uv��T�U#�����w�=�^T��ir�����J�����w�Q}3Τ�݋�J�����r��]ܬ��Q�l�4ൺt��pu/c�.�qS���om=��K��YT�L�3K݊�e-��@8nz*�͓*3u��r47.��;]l��ָ��A���]D���V�ɫӎ����c�%���+Iz�Y���q�W�S2֖�c�n�b�6E��V��;�N�lI����ޖ����0}�9�o�fk�f��Tң�0;�Z���<6���hj�y��B�m$2IY[W7<��]�.�"�6E\��<�(y��k��w(��M�ڞ����Ѡ��|�/���!HD\�bY��k�2��hvv\��u��z�OI'hn��(��b&J*H��U���[�T�\��=x���I��y3(�XM{��X�^Z��d��J�情Vyz"�p�LF�RKo3�^9���k�v�lF���ܣ:��eNO<�y��ۗ�(?nӽ��SÕE���+*E"(Ff��y�
G=�̔X�n[�o�lQ����V/���2[�����?&Y�}^y~eFTQCQ"rj�������eZIY�F�4{Ə��M���5X����|y^����t>�o�Х��4�Xm�dV�Ư��0s7Ky�|,}�)���+�*Z����b=��՜���Sme��������.�F��~�}��m���;�'2'RI �6�<`k+ݞ/�٪�}=u0��ޣ�X~���>sl������c7��.-h��m�6�t�֦[,㐰Dl��2ҁ��>�fs��+]�nյW�e� �H1���s���H�*F�ũ�����#s�j����zn'x����Y�`��4�^M೚^�ڭ���^��bp�!*F����m�;��폋	i�7O$�<�C0Ļ�+����&��+��o��rTk;�-����jh��hH��B�E7�=9��*l��2s�iD�pg�����/3g+a����G�;
��@U��U��n"HNE�!āxtu�Kܜ�7�3��#�f�Y��n����&򌄹<��<�S��ꢼ���*���D�ܕ�[(�w��e����ա��U�=钗�sF�zc<���Et�֗��1q�Q��U��}�bt�ӕ�1z�ɍ���W7���V�@���cI�5�H�2�u��I3�8�8n���+�Ϟu���KK� eؖ�c���ꪷaݲ��#1���
�b"�m ���dw��f�R�dl\>�����ukd��fN7h�&������wi��I`hV��xull3gm6�N�A�Xl���[A���u����E�ܱ���;u;�����}��8���4��21#F����0�s�^�]��͞s�.�^4&�o^+N�\��nx5�J1�"bQ�v)�U��S\c��F�"dv�ch� �����b�NG�V������b�� �i��?�̪~�N��Kh��٨[�j2�6z�EI��"�j�?�K� �i�ֱ7B�FH�nG�蛄f`��mz�Z�*�X��A�]��W��+6߉��/g.���u��g�Χ2��*��&/�Ƈ�i7P�����2ѥ]�����y��C��|en^mp�Z�\�����Xl��#���,Ȭ�3{M<�1�(��P4�j�K��ʍ�r˵󅖹�(���~�[�qy��Pg�K��E�݄�¹z^q��m��*C��Ʌ`^�ǈ�����[�3�]�kN��r�m��q���q�y]¶kh���X�=vӄ!i�Prm�[i5��u[g��K�Y�k���$�A�nk�sή2�	�$u����c�0�nn�{�&���d���5�e7]�@Lom�ƳRF=�e�'hdi/���% I16[K�տU�i�b��h�r�,�Lխ8f�5㛔6f�VVV�}����`���J46��\Sn�\f-6�O*c2���9KD�4�/},#�c��uɈ������/����w׈�� S1H�$��s��/Gp]�S}؏�B|W�t����Y&5<k�s'���8X;���I`Dwi�pޔzW���u��[q[�յ�0��A�����Ȭ��x�Q��
<�qI�+��#P��24��ɮF^<ZN��l�8���\��k�^Ə*��{����YW��c���ҏFl<��<�Nj���L��'�l�kf뢴�So�����n�]�����i�1�Wt�8z���y"��IT4���n{�o�3[S�X7{�]!�9��>qBo[t�*��u-�2�6��63Odi�	iƣ*F��x�jb����.k��R�,v8�š�2���]{aG�JnJ/;�����H�J'�H܁H R7JX�ai�o�,ծ�/'��|��5���.�9Y�A]�^�)[���\k7�9oE���P�-f��M�xV^��i�32�uvv�}nĔMLtͱ[��]Y�M�j�'�;���|�,��ZA�JH�M�{���/���7TzFR��m��*���&3�5��Ez�Qu~��{y���K�|��a�a��n��^�ۍ�zs�	�{��L1�C*�g��Oi�7ko�xǣgh�K�٩�;���D2S�+C����V���C���Ŭ��:���0l�x*�&!�\\-�&�0�����QF���.�ɗ�9����
����o���.�{}���p�0-�`}ۧ$؟���e��P"QE���ItzoU��^L�v�3�	�"8�h�DL}��>�Ţr��h��Y7�B��g	>����0 �-B˄Šͭ��bΙގ�Lf�(�X=�Odna��w4���V��
�eOh�����
��i9q��Q�}���_w/��]I:%��{Μ�P����Ǵt0��ŷ�M� e�.�.��˴cB�<��J\1�6�i|+a���qYW�À$)�y�6�;���Y��4Lt{��-��ݢ����{�@ܔv�2�O%!�����$���QTo	���{���V8OC��ytr����^}���'������jM�=<�ަ]�=�,�qϠ��E���!!�����{o�W[��s���7j/g����2O$8�QH[A0�&H}����]�ng>�y����<�yJ��x��xw#�ܻ�/ ��U�%� P�	L��ʜ�<�hу�[N��܍�U��XO%��yAp��@�'��{�c/ë�,�M�L4֦�j	!n� 8KvKb���~�ԥ:76g����=��w���u,Oզ��&|��͗�����x�
x�l���1�8��&�'WhM����'nU��45s}�NA�w���%� 7��Ce���j���]P�7�ޱ�t=+yJ�ly8�1(�q���"�����>YԦ
�T<v��[yh��N�R*�yJ��d�	��[k��s���<��'�)Iz��0�U�n�p�x�7����g�"J�m����:����g���jk}�����Fu��6'�����IЃգ��Y0D��dy�r���YА�����
�a��X��x!�V��0vue�<e˃,ԗ�pb����&��mT�ِ�h��Me�Y�m�ޱ}�gU����m;�ax��7�1 ,�g��5]I��z������>{6��u3]1��,�m^��9���"�`����KF�>�$��fk�+��W��L���B�
"�e�e�b��\�ú�e	��P��y`�TN��/{1}�� �5����L���e#b�eI���Q���LջAa��G`��&
��C��Z������f��Ӱ�Uc�i᧔U��Q�;D637j\�L�v��ٯF=��&����eu]��ò�Ԛ.���v_]���f�斁
A�9p�,����kM���,c͚��B�AA�m���![�Qa�5�Nګ?57�B�x�Mz����{��s�-Yo�)O��2�b�Ms; 4􀁖C�$�(a:�7"n��[(TR��Vd1p˦&����� �:��:hu݅IM��I7�#CzP�!��gml1�-�9��<��d�ΎDMѧ]+&��Ҋ\��X2i][���9g,R���7�vt���E+Ʌ���(VL_E���A�E�D�O����Uj[�-*��b�\XX Dxw��v�f��9kH�Q+��!5G-YFl-�V�0u�M�$�L�� ;v�o:9gvM>8�Ш��Y�j�Ęl0*��˜����s=��\��l�`:0[*O;����*V�z8s��P.��x������0�j�к9��c[��@�����nR�,�rǈ��5ֳmĖz��3ɝ�@�JV�]�rS�`Rm������3��rZ',8(�b� |xYzWD�=���ŷOn{Em� �l;���-1w3/]C�[C�%v���89�l�s�f��N0�%�֐!V��&�a4�jk6�M�Ƶ���y�k�#�Cټ�m�Wm3���>=a�	�c@G\k��8ܤCB�K@%��	��U��g�8�H�
��3�Z��x6^݆<;�aԒ�D�� ��56 �7��}'V�p-��.y˸7l)��=&��uٲ狓A�8�70h�\�k[B�Ub��v��6��Cq�ٝ���e��`'7:כ3D� fgv�ŋ��6�7cr����{t�f�sJ��>U�K��>��m��؀&	R{`�]��Cݙޗ�ƚ�l�X�Gg\�ݛ����R�v�������n����%�4�IO5������nL3[�u�t(Ya6x��슛Z�n���Ad����b��=����i����=k.��7��]j���o)\8��wHD��㦙y�C���v��65��7�ku�N�z�;`.�p���ee��/`�w���uK^�,B�{dw�n}�+9G��`ZW;.�`�;$�)a��.�ϊ��ѓ��=�7<�V��f���\eS�'Ha����8�<k�'a��q�O�`�[�^�f�-��>��Lq��y�ۭ��ku���4�Rkۑ7nq�)�.�m�ӽ�i�m����94Zv�6y3s�*�m�.�<�v���" �NxxyF4����au��1�`WȰ��9���a6+;�M�����=f�5�ָQ�:�������6��]M��C*cY�PNBb}�kR���7��nQ�r+��&��V+\�m�o;N��٩+@ J�J�����kMcHD�Ҷ�+t�ayz_GD��::���v�:�B�Q���s�/Z�f��[�S����܀XG'^�]��0�M�F[�W�d�4�UB��0��F%�ֺUg�ۏ.6�h�>+�㫓Ims��a���#[��@Iɰ�n��uz4f�N|�=0h���7vc��SFil�%Մ���=s����Uu�kC�n�W��j<��ا��~���<~�	��o�q,��)C~�o"��B�x��f����)��-hz������!�H�I���r��V�}�44^dq��^*t��jݻ;+m�eD�f�P�}u(f�"J�,eV�d�N�KnRI�	R9��tb��>�=-�Q��W�KCo,o�cԓS�[�F��J�I(�~Dˆ?xv�zR��p��VQJ�&L�B�-ڧ�:�O��Q�YY�ţ���۬T��.�a[^����i)��Т=ͱ�$�Ҵ��Y(��ޚ�������Y�^��0] �=�gU�{e9�*\��v{��k�@W���F��Y7C�s������N����dpSS��7c�:ԓMT�s)n�Q��ɮ��_~?���^���:Ǟ�;P�1�^�)y��:�k8	�D�q/ĥ������0 & -������l�n�l^��S�#�{����0�#�V[��V� 7/���Ѳ�J�c�XR��"D���u��X�gk�җJ�e��<GZQ�]�T�݉(e��I�=<�<�T���:������KB�CW�Lv�E���W�EF){�7��~�t�V���U���Շ�şITc��	��v
�v,�t0�Qão�A���&��j܏o�.��Z�q��r���c30����96L���3p����b�����kd[�|h���kͣ$mD�G�,V���4�Mm�1�(u��&����9�^�\�����J׾M_�����U˓ہ����*o��CB=� !l��&*���81�T�[�sl&�8ڎ�kW2��:�nˁSy��	e&*C~�m��Z��1��<�{W���w�mN�>��������I�uսs�w3�`eٺ� GȒ��a���,�5]�o�l�5L������<�y�=)ev�~3mHL�<�VP�5LUb�L�Uԧ28.R��u$]�$�u>o�g��Yz����K��i_�8zK��w2�B���vQ`RD��-,_v>�T�4=�e�fZ�Q��N�T�UJ�wV��y���lHp�(�P>��{P�0��x�6 A��f7u�gn,�~�tdW.�Z��q��uBO_�e)y}��VI�:kA�ⲩ��Q��~%k���66�׎x[�8�A'��7�����^��u1O>�L��b;%��J���0�c��#�r��դ�F���U?�q=��י}z��s�9vº-e�Z�պ����ӱtF��f}t���.���Q�F�a��)ԗ0[�҆{��U��C^{Տ�����x��%è�!������K��B�
V��Ny��*B��4��N�y�.UOz�[�{gK��z����A���P���Ƴk-�:ɧ'�>��Ǯ��ġ���tg�P�HJ.H5fV���}$��
���������Bv�Ɇ�&�k�
��mZCo]1��u��z6�%&3*�0'�����k�.����Ҥ�c��뇑��h�,��oө�����v5�V}҄8
��.4vr��	*SA�V ����V0�n�[��/إ��7��ܪ��@��f�iJ
��m�.������W�*.s���v�^A���DC��C.�[�}��tY�8��7�l����jY��m�2�@ߖ{	�Z��X���g��?tg�ӵnzZ�'��SքwcF������y3uۣ�qUX4аK^<�ߍ������&[����W``��r"::�^s���*B�w�qt���T��Mٗ�w���(�0�I��8�^�H%w����#�����n�+oH��Z��u΃�4�5G�����}2�>��n�	�J8Ӝ�G$�o��V���46�x�)f�y�J��pC��T�����KNcM=�Op�ol�q������3-DQ1�b2F띝0�hX7�����jr�(um�����U因���h3�����<�|9�**٤���S�<Ŭ!,6X�5$ͥ+v+����ׯ��ێ]0kL�|f0����<���ClRW���Jf�g��Rz7/��n�8�X�ɔ�>�V����@��i=�4,ŵ�܁������!J����@iJ��f����T��}y5Ә�d�N����I�$H$F�n�Vܨ�7Z��ljC8\���WBhKI-��C]z����)ՕL���[B-��tpn���sJ�:�ѩ{nj�v{{e���>��â��܌�)��d��멺�9�{\�2����-�Y�ה��T��q�#�3��ٝ�}?o�m����v,�p/=�����g\��qXv7p��We͎@��x�q'fI�:����c�b��iu�]�&4&&W(�F��Nb����n�S�[Z���C�	�R�^�����E�0�Q���16ß�yK��gɬdP���noL)j���*~�^ ���`B�7#�B��̞+ڵ��T�RۋvVE�ν���Q�����-��ȟ��߽t�w�d�ݫ��޽�6�d�n���\h4yvI��t�MU~�3���ˆ���z��O9_w��%����>2� �fd�ʼY��4�����|'^L���#��R��d�%"3����T�/sP���_J�w��s��o������@�˯.k/&��*a7�"�;]xz��*����A�b$-��^���Wid`{}��ȁ��LT�x���<�~�UȷWy3wZ�LK����N�{u��h�c>wن�X��%+�0��,K~��>��:e�H����P�T�X�5qI�p&$i��22��xuA�]�ô��T�˯\���♹5��y�����3�rT�;����r�A��YP�+�|�b7���q�Ȅ9���:hov�mnՋ�
C�u�܃7,�;l�r�{r��R'[�t�A[�c]"�l]��\�6��ʂ�����m��c�97��c��N�= ��ࣦ�/e���(��v�wX���ƥ���D���IQ�A��-/�^��=�]=�Φ����Yϓ	n��2���{Ȗ�O1�$U5I��7Eh�H(e�Tb��H^p�q>3�����o(�Zh�7����+���p�����9�εZ�hw��F
�[��T��[��3<��;����q������b��7��%'DY�$���Ķ���W�R<���BɸOc�y�ϵ�Lrĝ�I[!�c]<&Ϙ�s:�J!s���,LVd��[�������w�}S� ����Z�ɡAF�N������6���.�v��$�c���U�!Y�����/h�w�L{���{։�Bk5k'�e���Z��y7g+Hw��;qvt�7pdDA��y�1k�.-�RI[���l��*�	�(�������Us�xf�3ޣ��a�1#v���T��1�M�Ā��E�v>�f�e�4���H���?+p.���������v8w�̳
��6�s���AH�(I�u�f�I�A$�i��ݒ�m�F���ZC�i��6)����Ҹ!�rM@�1����`��u�Z��,����m�1E"y�J�IdCz禜�F�[yQ��gk�Ca���:�i�qõ|��=�\��>�?���>�3���3L\�L�(ij��m�9��Iծ�`[n�xw;s]�gy+��)��l�=T̖�u��T%�MF�S�:7de��ِlJ/5�1g]�GΨ3�s|�+�Ͷ��#t/=%�$2�N�k�{��)�-�t��W��[�^؇Q��}�c�`S�f�y{V��1��F���X۲����C! ��"�~���4�Ǖx>e��^+skmu�f����ezZ)[5��Hr�)�&l�+�yӾ���h�!��6���j"s0��W�fyex�=�z����8рFlg-.{��t�7{��Z�ҽ��2�=���w���C�~y��yh�g�ρ�Y]ڹ)gm�(��Xlã��C/o<'D0z�l��id ���[0�d2c�d�U�z�zV�eGc|�ք\�F��8����z�Uz�X9��J��ͤ�'NY�&i���~	�Z})ת�h�U��]���F�Kl%�L��j����g���!��8���v��/fa�ՖF�y8�Oۙ�����u}u^���|�X�~�=r����=y�-5�~���q0�2DSrK��y�\o��F�%����.i.��j��
��5V{V�5�Kl
_u�Ev�o�`vԑ�f2��3�ba$PE�
�(��"�G���v��ڇ9@�+�W}0{�?YM�ޮ>��r���u秫E�kN�-��b2G��%����ğ�QYH�'珼�p�X�˶������
�Zᝯ̛u�5d~�{�{=q_����i��R�
�#8��]NY�PB�yBbw�z��y���/~J��Y��z�}��1z����g��
i�Em���v���%{[��l��4]>��آ7yk�����s����uMae�w����jͲ���q��v ��3�t�������щ4�!�P��"b4�.�A���㭛kd8�<�q�"㫓q�o
`n�6筬9�,��C�T�Ь(�9. c[����7���^�蒵���	-�!�u��X�5"MEt�x��U��;�����rmJB�m=�g.�:�������>V��;p�˯+���ۮ�/u<������\=���/>Imv��Im��h�Yx�R�|�jr�O3�{�#�%�"�]^چ3�8&���e;mp��莧n�sS�n+\ŋ�hY�-��vn>�>���ܠK��n���!޶�U��鹷�5c��EB��͞��c@�����u�c������H5�.�-'$Q�$�FDrʲ<e�C���{s3@���g�*A+�O�ݾ�������=�� K�ֲ@�ܸ�𡻖s�@R�~l�ͭ�D�N-9,#�� фll�"G��_a���Ys�I�Z��tD	�qԝ��e���W`�uZv�A�WP���,�6#e7d@��P�9���&��}�B���@�o���3����I�K�����2c��*�2���(�}��c�8㜂9$��礬���,h�-R�z`$L���C����L����vkR#I}�J[%��)u�˺xrNU;�"E�F��H,�Gt�rŊs�O>����ص�ju�<��[�e\$b6����9��C�~�v��a�1QW�a�4Ehb܄§+���4��yui�B#'�9�(ʐ�d�RRK�{����5��4��rg��y]z��_��ڙ$ʴ6��Jq_n!�d9)v�LY��۱�լ t�W2�	Ɩ��
;Xx�V[j7��͕��	&e6H��7J�]D}+�����-`�w�K�Ҳt[�s��ߺ���>���ؽ�����2�>~%Șn"�!nl��kU�	~�I[���*#H��r�b��!:V��Vl��Y�P�a�f�H�g1�[�@���ƒPS�F�Z����@[Zץy�����Cכ�]��XmB��E�i�~�\�N_�;��Sժ���c��2Z����j��~E�
%�Lpf���i����UF>w��n�v��۬����(�҉��{�g
�vjR�}�L]U���81$�v�#��i�E'����\;��#�gj-�u�_/k���z˜�z	�aaLD`.!���o�9�?�Jw��~�kqL�˩�?bO�a�c�|��=�p��%�[C�ٹ��d�;7ΰj�}*�<��V�3�.H�N7"6���2�c�\HWH#q"ׄ�,ۤ��):{�,��5�A����lACPQ��Q���N�h���������Ă(�L")�%�:�P��a(gVh�6$؄�P"��z��(%޽^����8�ޠ�t�7G)6^ǆ�l�=���8.����i�]#�%��TzV^Y��ԣ����m⍛�u�� ���4�=�-G+��e���~|"�� �˻ח�U��zi��!�sR�9D\! ���V8v�mu[��n��J�v��}�͒-�,�	tr����"՛79���|ܺ�>}�.�<���8����m⣜�a�f�W_�d��E��5�$U'%�8wE��իv���ϵ��ې]�cU�Q(�YZ�AD�C�=F��*^e��CJ$�PF��ZNo�Gd,�6����dcw�i����ޮ�Ϊ�Iq���v��8;�
7�w[|�L�(��lp��j�n��g4��F��S[�����F�)�&����9[i�b��Ͱn9}�� F9���8��r��U�o_q�E�U8����T��K�U�v�<'L�`v��%�u��}iLb��دw�=�O�m(��$]իC�Oj���atR��`��*X�1���5��6!�J���ͅ�Y�+��KIn����?[��n��z��W���o���w�歝.���KeP��\� ۙ�bfI��y��V�ܴ�'�jʽ��қ���L��}��K`��A5˥t��#ȷ)���P�8Գu�P����nPst���frt���%L6 ��V�Wu�2��B
���&��\�P�y�C�E�5��d�`��IvՂ�n�!T�U��p�ٽ�QT���W=��LU���朦XWH��^r�uڱ�G��>�]f�tҊ�r��^R�Q���Y1�T�\*8��K;���ӏN�����s�}����Z��6�ޓb��^�%���/w}=�툻SJ����R��0��v� PFO{JR3$5	r����<�0��Z��B�g.�>�Օ��v����my��k��R���u�,��d�w,^܆���j�bϺ��ۼ���Md2��(x�����L2��p�=�E��u����ݥm��]3u�N%��\p��C��Qu����!��������x��Г���
��wH�T�Z`�X���O����Q�

1@�;~��bRp�"�H/�C�Gqb�;7�1S���c��e_Nf���U�̘/c`i���+p�fA�`3��;��LwBr��gawԐ��;ly.�nA$0�
����e�\�/��pѐ�y�����<Y��s>�u�'.�{��*!���]j+g�R4�$[֛�Ib8�[�ygG�w[�:�`�\6q��DP�Z\X�2��	�����B�����	>Z_0r�L�p�҃e�	.��9ӫ�/��`���F<=�*��6��������yu�y�@=�B�bb{}�n��R/"�s=�[ЊBv��a�V*|^�9$�ȜNE����D#�;��吹�c��w"�J�Ws�t}�6��7�^J�H:D�Ɛ������f:�R��. �*�o�q��s��Һ�lG]�B���s�n.���L��b��7b�9n9���Мq1n��b�/\5_��~����~/kUyW�ƞV�9��^���t�ӳ��{���.��Bz��r�3}+�=C�2Fz��[��P6#i�p�U\G�(�}anrc�\]�	��b�U�NG�[���u���(�}�n����#��D}[�)x3N�D�V�L����^�!Q��LB��^�;�Ζ� �(o����ʽ窷�4�ܺzqW�:܍qraxً[��4��p<`iQ"�nx1~���J@T$�4*��Ԓ��D�wn�.�k�PTb�_�9L���l
"�ńVT�MX!�r!�T��gR,��D�422&�L�����H��H�)% �8,i�鍮�Tl뼢��q�|:���_��\G�X�9�(n.U�X�"
w<j�-�#���aM�r��Ѽ���b�ah�rF��X~�`Y@ɯ6�:����TzM��3jS����d1��#:�L��aH��!���6�mVQ��尐l�d�H勵�8.F����o���{?X�CˮG��#^��J�nn܇Y��`���:M��v��t2�p�x�8��m���Ce�)e�bu�a�و,F�݌B�ɹ�Y'7����� �,�#���]�u�A�G1���"NDj��$����#���Ɓ�] S��J�(1Ϟ\�/	MFhѴN2s"�G�c��)�V Y_\��W���%��m��W�M�w�츩&�c�ܓ�%Hx�h��Ϡ��*6��{���-q�H���|}��]9���;���ʹ]���:P�؄׬��D&��c���QS�E��Q[V��Fu������}�5�*�n�����^LJ �N�]Ot�|t�Ya�=�0���D�a���*H�Y.y�'HHC*{sX�e��!]s�e����xp���p�ʑ���g'�
[��;.z���a���-�]���#2)R0\�n,�ɛ�e��7�g�o����1�m����$��B��.�1�fR��,���[h�y�3<���V���v�㾱��
1�\*8�a���\�)_S���K���iS5!����<]o�P��,�(x�J����`m�v6���9�$�Q@tǻs�=	಺qFSI�
M�`��ζH�>��۾Bu���Uy��C�i�nWn��v��C ��$Q���4�o;�S�Yr
��
�c�$�ܝ����yW}|��|��b��?{>�������)��WLΆ*���	���h@�28o�lp�;�K��L�Y3�r\zxݬ�:.�`pY�����(";Θ�"������\]G&_-b�B��s!���`��ȷ�X��_M�J�TC�2���^,WY�9z�髏��`����}΃:diqQ�'Ϋ�H�nl�W*���<��g����[	*�IH����κ��W�w͋��
!ì[
�~�Uv^�d]ZJ�$P!hf�M��ϫ�iV1G��\u��^���OMKt�j�#�F�.CB)�ϯ���t�o:(�<��{�_:Y��r/�)Pg`	G�7�}[��Kʮ�B�����WQ֮>��[�������{]؎Hb0Hb�fg6�<����x�`��kCB��\������LQ�.��M�=c,J�<X�dv��o�<o܎���zq�'��*�@�H��$�AD��K���,(9#��b�B��z��G�Al�n��b}�����qg4��M��>#ő?{�S����X_���8�p����[P�s]j�gO��qQ�~�(ao��̌�(_���H�I!s�6�:s��;F����,VW7B�H�'�d]��i�r��n5��de���{j�#��<T�H�^�0���,�[��M��A�0�6�-�"�D�a�f����� ]������#3��)fx|EE�E��"�������OFS=�C�:h%�l�i�b�i:y\Ѵ���P7��Ц�t���)R�=�M�����7��oydD���ݏ<�����t{!d�5rT�^`�5w���f<��.��W`�4��)O�o�a��͡Zv.r��;mgEꯙ��|���A��b�5���"��PUa�kuv��F'���^Sr�o&�	O{���C�<�i�c&3����Y�:|@:��%�Tx���u+��)7���/�����ִr�d;����L|iA��4V>9N���8w�`�4d�g�����^t�ٜ�����l9���H%��7Q��[�@�b�ŎN����ʞ�8<��t(C,?ez��2.N����E����7�n� :@����������h�uN�Mx���@Y���<Gʟ_��b8C���b��4�sj4P�v�{�+�^��5���O��~�/dŮ���������P��tŁl�5�fk�C���T��Wa�s�`�Z oi���6CH$�#xD#SJ�B�7����SG�׻�(^�6�ˇ)���:E�d}��M��@|@���[l	s�ycV>i;.Ϙ4
�\0��2�n*ۭk-��q�ةʝ�d ̽{���2BO�D�f���Q@���,����}�,Nj�Y��Mg����R�Q�՚|Ppm�Ec�Сy�c MP��(��P��(t8ͱ�h�;��7��jL{J�fdśȴ�Xd.m�][��#��g���,�̀"�)���AF~�̐(�-�+p7g:`¼f�m 'U���<�/�ͽ"��&�9����c��J���|#�o��^�Vj��CG���V��zK� ��~"`P#���]nP���TIn��(����\�P��ec0���͉����^���'���T�d��t� @kᐁ��4s��Z'�>K�zJs�+�5ڂs���x�p�g��+-��ع�v�����fC�K�wz{ ����{6c�o�8I��0ekD��u���P�y��wP{�j�����}]�S�O�e���1X2�jUi��I��)�DC#���0(�.]{ޒ���1Y�B5I�׽���ë��G�{%r���xEΑN�=.����<�����m�[P�0T��B�'U��d��-��8ڌrQ��"�a�̿d�tv�m�3՞=�,��O��e
@��G�w|����++n�6���#�B�14"p�3Vڠx��n��,t��E�;vֲEm�h�t�^r�����<�z2`�Y�%��4�+؝dD<�Ӧ�<4���w/ j;p��9��Z$����bN��St�X:e�p���l�)v�jޮ u�h6�ќ�+�[���'����z��WM!����7a�ML2�qp���&������D�Ň,S��%;0M�T�8�Yr������aH�=kS����wp��l�}t���4q.��"6���Y.2��ef��!-���ap�=��͹���t��n�ؖ�>��"���Ѷ�I���Cqe����i���5�12���q6�5��ƃ��\��{������Ɣ*m^@0�
k��Z��O�_@Ƌ�koi�˝�k�I�ksy�R��&��-IR�H���2���;F�=[7Gj�翛��>��9���#wZ#�b�=�;�k��$_�f�i֚�wp����C�x�4�<��Uy�U�l��iȖ����x�{_�
G$-�-�T#EJ?���}�x�� �t7g���6���c�Lf�U��.
�7�L��^@ռL�,��-.ݠ�L���ỵ#2��~�r%r�rI@����҇�B$5������71_k��i]�4�t}���}����62E�&@�ݘ��N6:['���{4l�`��O�l��@�ɔɑ�"m���;�,� 1��]��Bq�lw,�!+�E���x�z�6g�9�|����(i��ra�b0��V
�h^����ЭT .�`4�|�Pd�!Q�BҒ`�0�9�XV��l�@i0!�����7���j�tyD�`\DP|�yW�:��!���dip�<���p�%"�@0����i>�8��e�M:k�;Z�������*��k����.h���nXLB�k�eK���ǹ=��B���w�<@�;�U�dN�!�#�r� �.B+��-2�
v�+��Ǆ��Iz8��F �yX����;�s�==��_�<T��JסR�,Dp��(@,��s����b��/R�6;�G�f�fafR7rܦ̼�oi��|#��YIn�d�y��s���c��Y�|^�K�)-�ܩ�E�3A��y�ζ�n����OÁ��1Z�"�V ���'�D|��x���p��8E�����b_��5� Y�wSt�κrNM}�$ �R	��RDBq��4�D�9�ۻ�p����4|��P?3��2���A��|��<O��CC�m�߹�]KD�d\�����A�At����G�~ft�'2|��(�+*�H��{T�Wrڜ}+��W[�8�1������xTb�Vb�zJ�5BO$�P:�Tl��|�!�E^[_��N�����9Ӎr��!�azʅN�EH�U� N0�.wۆ�6��e��rȾ�*���{��4XYUI�d�����������(�0���<#'����X�੯�8D �k/{���ghmW"Ė�)8�gk�hnܳU�s�X�i�6��m���X���e���Lm���P�W�������d�C�x���\�Z�������!�/+�뙜ׄ�M�{�-A��^��#O:F���y���8��99��pY��'���J&�L�Tq:LpB9��r�<�ײPI��C;=�?p�sxD3��Nz�vP9��a�:@��/��߳�t�D0@yf�9q�b���lw[s_w>�w�i��~^��������
I/��n� 2�(�� ����x���[��?!g7�O@�͖5HP5
�p�I��{��U��o�ʟQ��ZEl�u�����Y/����!G�[�s��_j%z銝{��c>�|�/��E �-!��_u�<g����� �z�M�'#9&L��VlGᙺ�5��j7��!�f��+��x�#���2��;�\#���9��o:�0�D�l�U���b}��/�Z�m<A\��� ��:5&���p�$pXD�@HY�H쾥���M�Gu�X���{w�ɼ��\tG-�Z�zP��Cd<��d
�g��`#O<FAls���"k+zZG���n�F8�q ���`�5�W]qR��PP@��<]�;\����7D��8��"�{�!�b�Ѩ�W�pt�q,9�9d�nڮ�A��y��@�>}����K_k��D�$!��/�����N���:x�!��#��=~*1p����$�<d�.
<���A����}]�{tcɞ?y����dD#���9z�!H�G\s�҅�?	?�  ,C윾��K����1��|ug0y^\��R�E��[��v}�����5�{٢�0�x�0�f�����ë��.�6c4}D �|8��o�f�܅�4�Y G�ৗ�@s���O,����h�C�R��B�nI3�t��sa������z�<�<z�(��,�Q�#�y�<�~t�O�i��X����kNt�Qd� �_��8��K$E{����vi-58@���x�,w.ͯ���N{��D�yST���׆�u��/V�^狁�A](�����x�8�o�p�T�sf ���=d��Q3l����Π��G�
�9�xk� _�T���k|x#�@G=<v�5�Z�r�9� x�t�,�qT�I\���pB(�<����w��\��t�T� �,�p�޸1�F�Gz�m��,)\��,�k��%^��u�1�Z=Zk�kf];ڝ��������	;�:|���oo֫�a�288�zQ#�~��s9<y�G�x��iʯ:"�O�X��;����#��y�#�	]���G,ty��pY�Υ���e��<V��I�I^��ӿ�z<�'��쒸缕���<���x�f�8�9��n�s8�G�\#�^� {2P��r��2(���Z�dt��9Y`n����C�<���i�Ҹ֭��i��LwOe'O�@��^>u���9�u�Y���2�.P�f� ��f�қ��cC��N��H�k�a�< '�zJ��Jbt�Od��'�C����v	�pP��x9���B��\g��� ��oo%sHDs�G8�G ��׭W9��	���p"4�G8;~�9�9�����G�~��k��[��,���mE O�aҝ'�ѓ�������fQ&�J�ˤ ��g����<����PT� �.�ks�Yt%YT��Ob*]��j\�>��.�O� ��9�� ��9���N�����:I�wws:I�www��$�;���Βt������N����?���I�www��wN���IӺN���$�;����I:N���3��'ww'I:N��gI:N������'ww��N������'I����t������:I�www��$�;����$�;����'I����1AY&SYg�	��ـpP��3'� b��)RR�TR�֭�$HT�H�kUR�T��*	U*RP�T��kAU ���Ͷ$�E"�T�J��J-e}��*��J�� 
�
� $PB�P� HP )T U"��AAJQUA(��)T�$* Q�%@	P
 P�D)ST��ާ�*N,�BVq�N��6t�m��(R�׶�W=�B��=���e������]�u{VV�� Y(�\��m�]Q�Z+�F�ms��z"��ܪT�sР7^�J�
����Lm��Z�PJ嫶U�w��{������ԫ�w=5�N7\��mr;��I�@�-d[oyEJE*�$�
�@P�5�{ۥ^�*㛬%m�7z��K�t��=���z��V{����U;m������o=�^�KU�
^���n�W�J9�h������ַ�m���R�W�{V��⫶ڽ����-R�����Z���U�z�-BU��w��b�=��)w�꽶�b�PKa�ފ 
@RT$ ����U�]��x��cHN���m�4{���[m���T�����8��6����G��w���ӥI�<SzZk�]����ZEe� ��nD�oyǢ�S�Rޞ��\n�m����W���ۉʧ)k�nQ)y�y(Ό�eF�Z�%^��/D;��%*��v��T�H�h(�m�=�T(�
*� �U �)6�\Yב�D���M�K����K�I%�Q��� ��I�U�$�=�/6�^{���{h�EGj碀o(�M�9�H��I+�CMh@�U\��ּ�=�GF�<oz
�QEYe/Y)qEɢ���D�ziw��H��ǞRJW�����q�׺���'"�֏Z��:����y�D�o5�P� x U*�� R TP^z�E�㧑����q�'�GE�:D�<�S�*��Mx��PS�]d�s��٢(��n���dJ{�9J�Oy�"RU��B��J���mv<�U�<a��4 �l�E"�8��Kf��;��B��QO7� �R������7yt�C����m���]����,i�i^�py�\�0��k�w�N=�b�k@3����
��g�m��t��  ;��{0��Ѣ��h�A� S�0��" � 0L	����`D�2�T��   ��P)�T   5< �*��C�S��O��ƿ����������q��Kޞ���9�p 9�ru������  s��,p 89�p#� �s���8 ��9�G8 ��8G ������?��l��R��ђ���m�کe��LCe�u�!�.9j���������c׊��ݙ�od�b!�����PN�!�ș7u���;T+{����q���=�u�;Ѷ��{g2FG�s,�Qf�*��eM���cǻ+�����n����SIm��L<�W�k˷�['��Ћ(� (nc9��!��C�j��U��A�{��	��J���^���*���@��Y���)��+� ��SCFTN�͘[ڂ�r�׆��v�	U��"�Xݍ�Y6/fS������6��g]�&B�9N�ܘDD��YV�VF"6cSS�ۇ8�&�m���Ҫ��K���E1�q2�^��׷�����B
�<��zk5],zj�䑘�ݱl�$5��T�2�D�y���Fbg撘����=�!/DջV(���d�؂��hm�_�#c��4�z�!Z�-d��T��T�"�Y���E���rƌD����h����Օ���#l�Z#��D�
�[���PkZ����r�m��3!�^+(*ʌ�ŨP]'.���o �&!	�w6��"�#���4'*�{�ǡʊ���tD��l�cɖ�ynj��Cn���Ik�'!*,�U��2�u��õ�c8��U���8��{Mh�d=D�`nJ�,�ܱ���(�M�rK��Ōc��pm+Ȗ�1��0����^��9�(*�q,˘V�A�&����"������t9el`��М�#p�;Ш���SR%Bb�TH�\�M�:uKJJ���J�%7ubwz��b��i3�sw%��/dZ�L�D��)�GN��iVpϒ1�j-�Z7+i���@���鱀�2�1u�v����TCe�\7�O(n���Vԥh�Ǻ4�[Լ������ɽ��b:��0S�.E��Ea�Bˑ�wW%�v�/7AשU֜m=ǭF����r�u���9�`�E�Ų��c%�A��;Օ :�3wGdP�KI�mS�^�T)��)*.�,VI{r�=A��LX��.Fν
�iV�����HG �.�e9�o*�ęyU�U�0\{f�[	T��^�,��N�ŏN�l��ʎ��t�\VS�E��zu�ػ�b1X�m�N��60N�tS{�%��5��Wz�k*Mӷg	80+��1*��-i��:�[�4G^=��9mU����i �z�ڣQ�Na֖�&�d�t2c��{(X��A�wyiTh��O�|⚮�}X�|s!q��H�[e}��cb�li׈`P�ՕYc���i�ӝ�|v��\��*���v�.iٔPZ�Ą>���N�:�6�4A�u�J�ʆ(� ���&�N���L��g��k�� �Ӷ��E���½l
PK����`��R�#����Nbկ$��yF���޻8]�M�s�V"�5�n�N�ީA��
�8R{YQ*���Tn\��m�*e�xS�5K����Mݏ#꺰�T&<��q@�#.�]��J�n�9x��]�$m�5ǹ�t�ي���F�nAT��f왥�-�u۹)�5�1լd�v�*�HK+����y6\��=9k]-�Ke3�HE]X�|y�I?	������f�歨�5��]Mj��:�qʍLX���nn:�BB�vf�Ct�ܐ3Y�Rs10D����Y%^Z�C�u7�b�;3��lp�CN�/Fa%��Ց�!wwx&��aM}�(��n��*�Ti�%e�M�,�,�8��fC���Z��f��F��Sɥ�;tt�x�Lۦ��F�й4�m6�v�!�b= d�7I;Y{(�CdɩCGY�%��xV퓄Fɫ5�$9ȴ�^X���!���f�Kn�(�p;P�s-j8����S��J�t5�e@��o�`;���dZ�6��bd��X��h�FV�iF@�4�+X��q��he,��t���F3*94�w�/p�x	�/IMې�c�#t�?@P��Ve�L3�dv8K�Qhސ�,�q�N�<{��6���қ��5��L�C6��Ʉ�Zэ\8�a"�ݥ1�;@30�̺�fIi]�����^�x�0j?���,�X��`&�����y�S~ʶu*fեgq�L�AŶ���1Q,[F��(Ѹ�+���B�$M�R@���tR�izS'2�Vi� ���nfJ4��lb�f(,�[���Qn�jf�uM��M��>8����y�e�$��8�k55���v�ʰ7n�+�7� %9҉ٽWa�<N��f�I�m�OE��+	WZ���TB*N�K�kF`å�b��Ǚ������l�F�bfb�M4��o2��j�%�hݡ�#��QSaz�\�ܚK.೩H��rib��9)���u�"�:i�;�%G%�Sg-��e�{xbx��heӔD^U�oe�f��wE�q�L��b�ŋ{.����ad��KwN#�·�J͢Y�Ve;����1���̧]m=�H�I�N�jI�w��r�W�-5����/Z��@R�z+B�k@cMm4�9�9Q:�O5"�u�v�#j��n�c�B-}�[VܻkEt�YN��֓+a�+oh���,�38l�{v�2[r������CF��&�]�;U��ӕ��|�5���k
{+s[���P�RCnf�����$���c3�&B����un�&�ޫtM�XÅ�����V,V���L�sib��@��pV�n\���I�v�ԅ�����R�I�Uҕ�Px0V�ocj����Tɑ=�Yl��kQ���7�oI����n����WY�Y���p��GAnE��3,Gi[u�W���V=�芥���&��Ӧ�`�Y���{\t���ý�`����(�WJ�=�F��]�B��CTF�,1�yv&q�V��;c8�ݪ��Y���SE���-2j�&f�*�fʐ��Q�p�z)mV�gO7�Z�~XE�`GP�e��X͉V�զ���/#�wܐ�1��w�N�Մ��d�U�[NI��d� ݄%�N�c,��m��eRФ�l<Ň�l�&��؍(e�7Y�n�*�VU�u�fedR�ςGJ�Z*bt��{73M���S�Y��)�0*2n�̹��HKASֲlF�B�U�3^�%{E�Ȋ,Gsf�ȩ!�à� ��D%ynb�um��Mgt��rmf�:�,��9��Ȉ'U�˸�.�i`�6H���h]�8(C�,�e���7B�n�L����m!��ÄVݥ�doD��n������,��ˎ�6�K5%�ۼ^cl��I���T�;�r��n��w#��D�w���Om�x7V�+�[k)�⭎���ڕƛ�+ne�PLx�! �Ƃ�&Ǎ3.ު̺��
B����X&��J��F�AŹQC�E�ܥN��˳)�m��7�G����ٸ��/�#�-�0IH��I�F�9EG�7V��n��GmK��b��.��I�Vz9!Z�����դ̶p[.ӽU4e�y�ژ�w�܊5�պgmbD"��f�1P���7��՛�X�,�gSm�%sm�� ���X̬��QeSZ�N����cV���*��y@4H-�5�U��.S�Kbc4���G���1���൰l��R������ʁ֍�H�W2�41Í]mÔ��������ǰ&�X>e�ƥ!j�7	ݡ%�Ȱ���t5,�3-�m��z۹���ej!�jI��#�r�o�y���N�e�fC��*d ֱ[�z���Q�D��n̕(@�6s7A�I��漩��Yh҆��oV�-q�q^Ԧ�$8㫩�sT�UT�طF�]E�V�͋����i�q�3t-і5��6)W���a��xY�f꙱
i��j��EoNV=�Aݬ,Uŵ����mNH�3&���jxs%2:h�͖.��Z��r�b�ĉ.�ЧOo�-a�Of��L��M5z�d�PX��F�X*F�^H-Fr�3��˫�3�B�F�����%dGnޡѱ�� b�M32*Xt9	.��	U�xv�;d?1Pb�J�2U<ǐh���MY�i��]bÐ��1Д��ڵX�-ay&�b�d�h�V���2�9S�UQ�����xS��Zf
F�l�5+��ٱx��n��1�f�0�sZt&�ub�J˄�3���������/�K�'V[Ҩ��i]�tt��tB��<�����x��,��ނOUWh�N��{GF�e<���}]p���X-�Ç��d�^���:��	oAT
��p�&�h��%h�3f�iil��yw/lc�1e�x�f������wH�e	F��)-���h\W,Ҷ�`����m5R�Owj��sw6Q� �i�Ҕ�ۻ��f�ct�f��dSP'!���ǃEL��/�дR]�o2�%�Nٸ���{a�u��/f�L8�vmF��v9oYa#�%G+]�0��E0�Y�e!�ZK����n�z��>:fK�b��,c�'f�˅9p���)
�/rD��٘(j|ր�`��r���%��K1n�����"���ܤ&�wv�hi��G�*���VMj�kj��+yMе�I�A���Ǥ� Դ��{q��Cb+��v#4����v��{
�Si�ub�Vkf=�-.����D�P��2g��;�0p`jQ�i�*f�c��^7�~/2�D�B�m[���2�P��q̪��K㽒g.����49}�Զ~u�ו.���HK�=U�<�C<���	Q�S�[�:q���N�f*���SMفؠ����c^�X@�U.�:Ͷ	;Rf�����[�*�8�A+'�m�|�.�Νm6�;�K�������5��l���C����k͙�8�n���uA���%�����:#��A����UX��e��F��BF��%�C_QWuo�Υv�_mǠ��=�l�S4�ޡ$��+Ww�+�͹��ܩuV�-'�d�g*�0ȷ.���fK������AK���	�Z��rR�c���e���Xp�2�ɡGa��>\�܅V�\���e_GI���s�r�"��јjh���L@�k#��U
۷p�*T��%��&Ό'�9�*�!��hM݋UV����3�L�/+&������5���Ne<Ņ&c�������S�
����Vu��F�2�-��0(��@�ƢoC�er�s9X��%���i������9n�u[F�Z�jf��j�BC�Sv+t�g	:r�(���i��}U��+s^�z��"��*�:>6��s��&S+D�bR�M����j��[B����Mr����L�ES�:YӨUe�kj��Ҵ30H,�xs}����ѻ7��pXx��^&g��V�Qv�ː���� 6�����G:��#��:��(��;h��`��"�tڠ�;v����[��D Ӱ�G.��T�2���1��s x7(^-�*%`�Y�q�wdf��*T+"6�(�x��L�"Qɸк�.�5��jj���y�5J�:B�o7X\9�����M��Z�.�2�Y(�Qn��Gקt�B����M�Y���`ٕ-S�o Y�	���>$�{��P��r�*�PD8�8jah�
Y��%�A�E�ڗYz���V�e��t��z��l���t���	���[���
5��W��U5��t+v�ym���KEjiDF[�Z��u�ˣ�.�f�j13��"Ln���p"E!���;��7V �K�.ڸ/TհZ��0c1ֈ*ZOQ�	(ԎR��O(b.l��1�]꽗{�P9�c���cZ4v��%\FԄ,�6�J]����p�[�Ksz��Eβ�k	<5�A�XR8.Ck{[��ui�r�����_;h��(9n=�\�[��ET�*��5[6�V�b�W�PZw�`{G*
%�F9 UZt�!6c���:����x�^ʋv֊�� ��n�V44�5�1כ�^ JpZ5��˺�C����ɨ���O�W��U�]�Y��侗
K,;��D�'N�#!�&��Q֞K�e�V���Z�c�����ctq;���oB�EkS���))���[se��� 6 ��[����B(4k,���n�nj�1Y��T/չi,ǉ]�	C�<��%�]�x7���7&���V�d������^L�'u�Ȥ.����hVmq�jɣ� ����f^c�1�z�a1e�*쉁;��xeە�G	&l�������ff>嶺����,�<=e���L����Ӫ��ŕBhMN kQ�żA&(\��i�����1�a��3j�$���6D�;i�Uz���T-�5�hf�X.�J6�4�=�l)D��퇷xcT�-n�S0�R�j�CQ6J�.<���F�Ě�5�yp��ʹR-���uby��wW�Q!�4*�ݎ�-:�g^!���Z�̩�8�ʠ$�_ڳPU��F�j���C��:�a!�ZB�j�Uå�Lvø�%�EC(�ҏ�����X�m��5n7)��b�6&gm'P�i�a��K�G2�xn��(�����w���!�m�֬�@K��TL/oX�k7tyC~e�EՋx�����R�9�M� ����e72��˭�7���MaG�f��DKu�Q�b��G(ҡi�P�2��N���ZYW�1v1�YG$�V���l�%��ڽ���n��8�J�)�V��P8yU�&��4������L����Z�-k�mA�v�a��v�M�D��O�B�oF�Y%<����51%WZ�ὤ6VƋ����s:a�rw��:��J�&��h���oI���j��L�κۚc�����wg�H_���lO��T�֬�n����˓��@d��Y��������v:�{
YX39 ����\�c��ؕ��&�(S���	�n"$�
���-�u�:�o-��7�f�F[��n�h�U�ЦuP�b�����
#���2�ݴ�C6�p$gc]���ǜ���Xyŋߪ�Y]�����GAv���FbV�j5(F�Baw�p��)���*���P�m)��v�������m�6�m���lA4Ŷ���?�Ͷ�����j�*��v�T�V�{KUT�0WdA���Ut ���uUr�*�R��@��rϬj��ڶʶԼ�)��v�T�ۍt���ۮpnvy��u�Nҫ�������媥Z���mZ�V��i���{U���[sq`�%�]����e�R��P
����(��z��s�5���1h�4�b���m�>mmO?�}o������Z�a�u�dz����=��iz�[��1�N��:�G�kf	3�d:�uR��J�V�+p�ZK<�r�e���MI�(�b�0�Y��]�*:<X+T� d���HV��$M�Ħdt%�Nݥ���8j{=&+I=�<ST1���i�U��ݽ�_�8�uƟT��9z4;hMA�lg�:6�vٽ�!����jc�C;��x[�Jj�S�Ѽe���u���bl�S3�]�Ƿ!3���,j̗�-��h�,�EbQ�gk��3l�ͤlliNNɗ�v��s�%����,[��V#��ku���ӧ�j��>�5��^�Ƙ�eҍ�f��>�S�suמ�16f�+��c:K��d*�ڛ�\�my!���(g	g\�TM����������lC2�W3A,9f�2�ۼJ���I���ϐ�Wi;<�*]�n���[=��Q��]�c2���C���k��7��7	�W(�ԝ��G0��l<��F�n)�H1�,�Y��K\��eix�\����0��SLV�t�n�sr����7l��eg�:�;��3��q�2��
i�v\q���n�X�tk:���tm�|�	+�wq��=I�$����7<�s���'Kvϳl�ٞ�7V��<l�i�<�n�d��~��N"�y�s�wG;��SVy᠞.���#�z�_nL=�q֎^�ľn*��xN�b�Zٜ��r��of	yCԸ���ێVڸ��.}���7k����օ��o)��C�F�
1�e���Ÿ�����z ��$�
��#��"h��KJ��T�q۲�A���;�4�&�A�=���Н�vZw!�̳ih�� ˢ��5��H�'�ӒH�[Y��p]m�"냛ϥw0�]��{xY��qm��U{;�Չza��;���E���#�Z����9���j�^X�j��csTwk��<7YʮӞj�F���2�FQR3,��v֧<��uvm���e��Lg�E��X�m����-����`i��dݳ��Js�����N�� ;$���'���y��n�/��Պ�۩�^4��D��K+�n/pu�ú����⳥x�=p�![u�9��aq%��5����zצ%ۚ	���2q�F�y�{%�����k̜�t{�v�t]���'v9���-q�'D����suփ���%�cLhna^i��4�J�Fl�G�.%���f[k��H�^��t�n���:xM����^m�t�</h����[�������<d�Q�&�h4��M�JJպ�m/bmnxg�v��n6�^�	��5��z-��	�ܗ�����\�9�tA�
5�nEϮ7��}r��-׭��s�wm�=.�ꍱ�S��<m.q�H����!��t!:��,q;wI��k3�$:�٦�Kd:)4�at1M��ȕ	[.�6���ǡdl#�vw6�b1��lc.�%Eɵ����Ď�mmY�Q�\����;{rr&�9�E�\����w���+��z�]�5��s��c��Gcw��ӈg�ah;H�a��r�K�MH�̊&&�2������
r�v�`��Ϸc^�z]��b:Vh�5%��!��KvF�H���j�ضkX��0]l�^�h}�Dq�N�6V��ƚ�^'m��7n{N�87��N���������xsVlYA����%����{i5%��n�������0v�mʜ^ЇQ~�>�FwR�8���.���'<��V�%V�!3�5�60���l���@�v�c�Ϙ.��3m�Bcb��9TR-�����|�z7e��ѐ���~�g�5���f
n.۲X�$�P�vmugZ@�=���T�*bh��!f.��(��V�0Rh�Y�4���2��OI�ӷN��N1�3h�C��Y�����8��~ή�T���G��a�./\R�:zs��$b��6�<����u����b6�v�l�s�)�DmͶ�@�1Ʋ�qח�����w2uy�jϓq�e��>��L]h��}����+u�F���Ν������q���:�۞E�[3݇4�Ύ�m�KUn�.9�ѵ�zݤ�kf�X<�۷�����ȱ�]&��}�#���
8�`��6�Ha��Y���X[+��F�b��j��y�y�)��[�ϝ���lm���<u�z)���5�+�F냮{��"�.�ge�3�5��p�1��t����Lu�4��q�Ds�"X�ј8�n����y�U�ƓMͽ���퉛Q�c��έ�Om��4Z]mYA�Fmf�P�傹�N�C�Ky�ܔ�hw<z�Q���=��]��rt�y�҃�=v ��h���z�p�X{���H�G�I�p\�v8��'�^�9;\<� +�G+�mIIt5���;f�o��;�AS�`}6ݲ�6���k�I��p�5<���P������ݜ^�P^�q���6x5�Y	�[\�]2�:�v@�qzq��I�/-75vT�j\8(0������^f5�T�P4&8���6a�083��t$9�H4څf��o��l��m�#ps�pC�SV.�[9x��c�Z�������GT k�j���yl����V��E$�{t]n���zv�od�O	h�������JP����5o��r	.��N���j�8�񩀦�X�ʲ������جn�$v��Ev:���]Ggdm��tpe�\�buz���"܆e��U�]�g)���O[V�w�����C�����!��3Ae���Z!V�n:�y��-�yg�x�}Z�s���Վ�z;#[�.9G�[jU6 3���7�qv5���(n9��7��2I�9�5��/gz��w`M��#�:;$��N�p�s&�5��c�]��q���n���m��m��q1��=J]��ԇ�m'3.	F���V]�p��%h�ns��w8#��5;n�U`�>^Y�Ўv��;gqn-��N��-�d�\v$�¡�lՅ��k%%�������`:R�B�]L��;�g�SimڄlZ���b^��u�0*�3�.�ΌqG3Kf��5�h��D�!��z����<;��2����T�ɑ�5�LN
�mT��zݰ�%-���u��m�t�7xf��m�1a��fO5��āyU�y�b��r�ajĵ6wU�
ϕ���uk�	�����sr!�#.ܲ�Y,qx�1�0�UB:�籼v��q�q�<%����؜�����Y;m\K�{Vt�)�b���;4i��9��p��D%PK���Y����G��
	��Q�^g�/	ӹ��֋++�\��<q]1�>�sj�tZ�k��Uc��#u�ڞ�E�V7p����{Y�S�oWb,]�a�[�F\$���6��;r���r���N����a�Yn�J��5�jDm�Q�66�����D�$f㱘b)W\�B ƪmi���Bmtr��q�u�	�'C��hQ}����U�-��OOuIě�ɞ��<�\��K�˵�\h�],\��
	�9�Ά�:�F)йø
�Ή���7k��Q��-��X;�[����A��쩽���C��g;�-�cu��t��n{k���wC�pn|�Gm��@���g�]<O<��u�o]\yz�p��J��VͶb�Xt�Y�� +c̷1�km�7q��Gl.�BD;[w)�0�-���ˉ���*�i
���J�����^m�Y���n�_<c6z�"S�&�ۜh�)ڸ7���E��3s�K�٬б����4�G;6q�+�7cv��X�Q�Q�=�֫l ��z�N��j�lK���j"��)h�t�8���Z֞ob��+�<���-L5а�(R��,���[��&�S�O=`�x7Fa)�u�c��]Ƭ8��qpw˰ݜc3���cN�l�k�y���N��z}�[�4���jC=]RO������;ٮ�5[����<�<g�Vuv8���3����xG!rWE��1++-�e�kM5�U+{���S�.71�Tf�v!��n}We��pG����0�[a��c�v�&�L�a�3������^i��Ђ�1-v�)0&͖�ao6Dp�夵"QQ�DNVi��
kԉMX��m��Ջ6*�p*ٙ^\�U��<�i%���X��g�n��.{\�K�0:���)+�n:�6<��B�,���7G�=rp�C7k�m ��]+�e�3r0��+C%���B���Ce�؎��Ѭkr0ڸ�Ţ	t�NP^l@�V��\��pp�F�-қXQv�yyj6�S#�w���3%�4h�M��Fj�f�fu@��VZ8��<l\���ٵ�i�1�7<N�ΥǇv��v������'������-��6�'2r;m���z,w��o��y줧az�����֢!Y�5�b@���̤�gl������z���Z�-���㛮u��sE�K���vGhM��*s�T	^��P�G=f4�y����ٗE��s����l�̀�:�=-�bP�Q�2�'��M�v2t�R��f��4�i2�r��nbG'
mf��%����n����6SY�3�j1(�ڐ��VI�Ie�@Qn,`
���|�=�[��gn��\hCn`����-��݋��\R��Fk�.0ډ��b��mA���fYyvna�-���N������XD�ڀ����+����M㗷[==a۪᪻w���<���Ss�L�}k/j�*�f��[�n�6R�fa³�󦃳]���u;p����T ���*�2],�,UpF]�RX�`�9�Sd��r]qn&�b���%⚺�k8��`����ԧ����=rg���/m����;/����v�nq�ŸH3,�gml����-�:�Eӹ�����un��2���䧁����F�̳1�SF3K�w-�Ȗt��z���F����=i����mw��*{n���{m�'*k��^�qU�{���9�s��#� �s��͎����  89�s�����I�s�9���s�rI=��CmX�˝M�Gm�ʨ�E�E��22�GvW[Ǹ=��sY��s�!��82�f0�5д���m2in��0�f6]cH���"�PG�tn���1�sMv�J�nR�6V�\՛Wv��*�ڹ{8�e	�彀�ZhK�o ���*ۃ �5q��^��P
��XC��;�u��7m�r@+��yX�l�oQ=��K�oR(0m��B��0��4��4���l&����wH-;������N� Ū��iÝs�b�vx�v��_k/Z��ո��e�Z��s�;����p���[s!Xi��ԃn��5�Ӟ���l� ��f��;�w����I��q��ݢ��nRڌ�j��:�7��\�%��ʉ�b��z�/<�g,4�S�n��41�yȪv��.���X#����Y�ǧ��k�+d���tR�h&��rF왅3��:�m�존nF:s�g�ۃ)۳Σ�k�e���.稴I��O�ܼ��/g2�T��)��8���t箁��v{j:�霻:yN���`�s[��PU+u��]�Y.�۷\�/
�N��ݺ0��aO>ڸ{m��:�i�mfCK�)�4ʓRZ�m��<t�f�����ǆ��i�0jn�`
�wl��u��ݠ-Ÿ��Q:m�E3ۗ�Kf��v��v�K�vv穑�{#u�^.Ki���\+�Z�hNwN�I�n����.��vN�	�&�y�4h���n۷Ӝ���H#�����yݍ�O�7$�O6n�kp�|�6l���T&��F���*1`��En��z�ۗG]m��pY���u��2)��*3�E6{;��y�7��v�����n�e�V�[���ٓu��FMm�m��&μM�MF�[�d�r��{q�Q�����wo^���������e �l[*����ΖBV���҂lͤ`���X�ȕ�3:^���tZ��<v�GE�h�٬0������]�g�*wY<�=+���^���צx�g6�7��=Tɣ/�;Fե�GClFt�]{Vٰ����{������ޯ�o�tT6�v��H�gk��(�֔��Jݑ��1��ĺ26��%��`�Qe%[���x�gT޼�v�}(�Q^tE�p�=��ڸ��K�
�I�:�oZh���^ˎ:��k����v8ㄥ9(%su�J�Y�G�(ԑ0#���[��úݯ'S�Mm����V3x��zsV��ۮ�a�f��0����C�sκ����7]�s�mb����m�PR��Tb��hF�R��iJ����҂@��������5�Qȣ�\��+�t�{ И_U
�sV�Q��y��i&��}�"gn%2$�ׄl+��b�dZ+�x�c��ݨ����2
�]a�!�o�%���5e]W�!�.�D=�Y�!�Ѷ#*�������i~���vC6d�����"�"Or��BooWY�#��,��e�rN/{��rB�R$ْ��bW���^��.�RM!��a�?<S��ޚ�a�[�1_�nR��Go�"�)��@�sz�CY�s��G@Z�fT�*.���[DA���OX���]˰`U$[%u�����:bP���Ʀו��&�J�*F^Z��(:WJ��!rk&�!v� R��xi��c�E�ί\�������Eo��`1[�Y/a�e
�gX��H�]�"J�����21`1��"rH]#����S�ӷ׶E%1۽h�P��A�v5=�b8��;ò��L� :��bZ��9,X+7(<V	b6D*�e�3�%�.R�r��AZ�/u3ׁa���0u��!��>��y���3p~�L�ܭE����%�(�EIY��=�}f{ =�n��C��Y�.���v�VD�]��}��r8Q��mH
&)e�C�<zzzKYzou��������K��ʝ��`�p���=S��N�jv3�!F����8�i�T'"��7�:7w�f�峬B'*��YB�`D_fu2s���Xo���2���v�o�1	v�G*E��q71GS�����ҶfA�s���x"�c�y���mm���L;m�<;,�)[ven�S;��A�rw��g��6Ms�Y�r�f��R��۾5�;{\�ݳCF��$�h����*2d�H/6����=h��
�a���n��E����[A�ޔ*���?[��Zu�n��{�7
P���8�o%�l�wՖs���"��>j�4/A�����`[�_CK^�(ԗEˡ�(���vÔ��+b��yXD�(q�=��q��#��Nqۡ��\��������H����)#�Ep�v���f��F^"�e�g"��j6H0Y��Օ��p�]̼��Q�Q��{u;��[g��dŀ=��|1��ׯ�fG:z+���(HA�����y�C�=a���",L7�7F]�ű�'�7X���3`��OM;����:��;�|����5��m����4Q��=][���:�w �C���-?�f����P����I�I%��Ƣ�~__���r ��������ѽtD�{נ��i�+3#���w���SL��b1�`�1Q����#H��
�\������uq�~����^�v�y�
�^P~Q��{�Z�+�AP��ّ7���\=�mdѸj�=�X�n{�ܡW�4<��ͱO/{9y+ ����T��p)$���U�c��=�^U]n�y�������4,�#6_���k
�5C�f�B8��Wՠe�8���a���g})W�k9+���������7���t��+�kmn�L91�K5�Ge"���/#:Y��[�(������@[* �����z�P��X�;īąd#��\�\�7����wd�r�B��������LA����ˋ�4��+���ا-%��::���W9������޷I��\���Q� �b�*��N�cd���J�g�z���+u�7�d�(�E�D}�t����wFF��c���dl��%�[������u=���2���=z��_{˶-�b����*�G{3Ɔ���N5�i��F�r2�7�C3%�����E�-}>u���0uC�u�<�NC��0��imᏪ���#k`-H�JE-�v'�vF��=p}��hw�Oj��[�����;�%�}��d�h���N�#�{�:���ҐĢ-��.�0nd�˝��d;�e�I��$�=2��������z�_2��װF��J��*��gx��O,�&��DP�c:*!����p�&`����f[˩���m���66�f���;��;���)9ޯ�{��^&U�6:l�t��0�YlG���sOYyumlgDq��QG�{94�kv�rm�馄�4)�3YW1v��yY.����w�; u�=u��Tۗ�^gl���疽^��S��=����ܶ�p�g��=4Gm���^�0�*�`kR�~m�Ԍ�ѹ��<n+�L�#�*�ۉ�y��{�9��6�l����%���68Km�ic̷B]�\$�滏a��bw��:Ҷ`�z+�;e��Q��q�n�8Ӕ �9
�&�!�_e��9�aۨ�d
��/�m]-��d�
���&$q]�~��F��(<}�(�p��$oR��vg�T�
>�pX�+��cm�x6�\�a���;X��6;bI�g&�B�`�!!@ÒI�X�����*ջNxGv���ohM�_ky�{��}��}�i5�t|�$Fb�H�q���l�y��"�}�ma�����`�q��CH�]�T��[]]�V�
���a8��&&82�'}N:,ME"pԈe9s���MN�r��7�n�d�������N!�$⒪�n1v��Nd󣤽��C\M�5���V��jE4an��f�-�c�.��f�g�xד���e�6�5������oz�f�˝����vs�=K3ٷ���!�Ԓ�7]ew+��݇��v4�Q5��rq@��*�õj��Y����q�`�A��u!OR�cB�[�~��k��7�w=�/w&�>5,���WE���r�bAr�&{�ݷ����JT�z���*�ۡ����ꤓ%�X�� �ݴ�Eۖ��TTn�8f��v H-Jh`�ٮ�Sq��uD77d�!&֟x���K�Iiț��(t�$�;���X�u��綎.���HDd۫��X>)��7�o�G�'bFc�f�{+N�L�k)��n����b<�\��ɍ�{y�Y������r�� �a�E`J3���s[C�\ø�kAǯB��b�݆V���f���16�����p���:D#�������eoW7J�ON����\#5�JALõ�^��E�N���h6Lh� B){��>2�yGj[5���a��Kz����<��<��KY���3�i�[j�y.�^ȻS�38�r4�̇1�}[ҝ��E��sb�NZ��B��v�b����C�S�����]��m1z��H鲲(ȅ�K����]��-a̷z��lff-�m�j5�PFҰ�ҽ��8�3||�
�bq8r�[�;
6����,U'�]=ǲ�蘘�m����^�����t�w����#"i4�˺z�]���z�^B��D��cp��:��O������}���r`yL��Uv�x6��F��g�/m�� ��I�u�-���vv�y�6��=�o)���uT��61�.ډt���|�/ߖ9�[&�{�JY������u�ߟU��[�y���k�ǌD��(ݴဎ�=��>�˂�o5yJ��伯b�:6�3�������eu<Pϔ+��A �I&Ly;��̄vk�>�����3�EOY�������7W����WO�"P0�nA�\�u�)��Տ�G��
X�~׎=ˀ����h�$�ٵ�h�^<^:;	���N^]��Zs�Z�V��q+:c�{;��Ǒ��g^
M2�gL��z.����R���{��D�+�c�y����A�$�<���7��q�' $�{dtO]�Z7+w��U���`��^)���N�N�����G��.���X.��%lv���%�W*M	�6{u�v��}��N��8S	$u�	b���ˣ����&�G�]�ͥ�)�6��&�G�zõ������FH�N�7��S��ొ����.���A&֝T[7*yc鷳�;����	%��"j�0M���%NFa䗽���~����'z��<�.ɸ�,�a!��ͫW;�T*��w>���p p�ڐk�Bg�R��4+{�3��Z��l�c�u83`x��)0��� 
8�g�y�/�2�/+4�E��6���U��PǫtWU��3ܵ�z=��t�ӽ��X�1��E4U��B��˖��k!�M+��!KG]FmwEAyd^�gk	�Z�p6����%�"R�u���9K�Ь��.p��)]�W���-�L�14S|.H��q�Ȧ���%�*j�\���Luy��@9�+��/mԱ�k����]�t������v�q�����ݢ�N@�ov��T����m�0���V�H����gt�[�Z2��f�;�^;t��s�sŻ3՚�z���m���ϭ�ˎ�E/� W��+�:�[���K5�b�Hq�v{\oW�ۈza׭�\���A��c���mE�;=��m���r�eT���5����/UuS#���ǖ;!`�9��BЍ��a�$ bFd�u�.�ٟ����xS^�m�+��\��Q�஻>@}�����ނ=�YX7o(eeA jAY֦�*3�;�o��坚��ng{n���{��WX�T�g�f9�B]�!|�L9K���
D(�B�8�c�T{�a����z�}S��z�!,�P``�&M�3�=]b�J�9�p�խ�H�M�RG#�����-���tХ=�����I�9��	ɜ�"�EJ�7��`�]���׽���5�|�NW||�N#1�BpH�;œ+���޾�2T���g=Cf;H�{��[ݝ���^���l���ϟ�'z���u��)뇫�a��#b��v�&Z�9��`l\��˳�v��;L�1����1f*�.�u��Ɍ�޶[rwQS8DG�Kھ�U�1�Gn��%I)�u���{��n����f�t������cs�9�7�!�e/�Y�m�;�R��լ�'!�E��/2��_֟CM,�x1e�%wf��Q!��o�oN�t�]|ū$;.�njzj�ٜ]��FVh��ڌB�tL��8����A�<�K�~"_�$�����iL��0�U��ި.�k(#O��2}L�#�H����\����d>\|�7F�ks0W->�FW��ޗ���
 I��AoN�ݜʡ�x�$�J��3rn�0��;�����u��=�5�����y��	.j;��:��ד=����{��'�ͅ�[��x!�^-��]y὘��s��Z}�c��=qv�KI�c��9#*0��Ivdo���5�D����Ğ�v'(O,�������;�& �!NB�d"l���ɡ��4�dГ]�Sa\���N��{�~4/&˹�uW��x�G����NCYs+ �z65�u���`3������p�C�m��mw�K�M��\c����]��=&�ny\�HO���%��`�,7}�A�XOmo����qhR����YЈ�S��T9Zƪ��핣lv�o	Lv�67���fg]��^u/�(Ceot�q_Uk٭{"��˒g51dNNIJ���kS.��QH�c��
9*��P�����R�J'l�IL�g�C�Ia��Y�T�k,�o�x�B�g�n�L�@�eL�Ct���)�O�Ɯn���u��Cav��`v��ͮ�ךGi�����Px��%գI���鍈�{eη�g��eJFXC^3�q���uL����p]����u}��j�`��yg:�����7jV�	Y����Nj��j����2q:�i�|���ҎZ�c��E��Y�xl5���.����D���a�p�3���EmG����ڮ�`���{�q�Y�w��؆VeE�_<3m^�ɥ��r���zhd�h��q�k��-n�cK����
%c��v����z_0�T���r�[����T ���z!��)}٨ e�����|���Y��m��d�8�+�r_K+���6����|�9��M��b岍K5��5�>���2��B������'�+h�09p������q���v:�*t�{-�z�I�{�+2�-�z�N�����K0���N-�
�2���ʳ6V��Y;u,�._\ �Q�О�3jҼ�β��n+���U�I]չw�rFD��_u+ݪ]3p�M��1����D壯��]��V@��T¬�4�x�����%�3����x�WE����������<�j��4������\Dþ�ڱ=Ӂ۞�Ō�����P�QS�{]��[��oױ��E�]:���igt[`���k2��y�p:�ʎ����~�$	S0E���a�;\t&͸u����Rnn��ua[]t�.+��u��ߍ�����k.q���Ff8f'�0��ⷣ��OA'�������n�=�9���H̎L�XY3���)WH���{��f(��*���7�νS*�wm\�K�y��#%�	p �ųC��b�����#�w�2�O[�^=����)���#_{�)d��`� ����ȸ�:������ޟe���^�z��C�\�̬$��l��}n���s�僅]!����j�x�[76�u@3�9gTW����Ý��{r\fu�]��(�;���q7�G~�m:hh�����d4Q��*E$[l؛�3�=��$�v�[�H�w�}�N�zr��{ZҸ3��U�~s)�h\��ilmsv��i�4�;E�b�[�Qʮ��Õ�"v�T�5��G6;6����h�~S�_�뺰^FH���a�W2޾��K�`���\��TɌڥ�k����r�m���a����X�߅���^GM���]������Vb�k{�z]ڄ��gG���ȉ�df9	�z�>]n��8fvzUXN	]�µ��7:�ܺ���gV���";��h!�#r�Nu����k��{H엧�ݾó�,����(+2�3�n8(r�_�z�y�d#���L?Z
B�Q�s�e��뗙�6�ҠD��3���8�sf��1�d�u�w�E.�2Lv9O6�Q�ꗶ���N7y�OL}��Kƭ��5���ֈ&�����˩;}MJ��=xWM���]ECa��Sc��[��]���m�j�÷]Xz�d�<q�kn�3��LGsJԛ<�	A���[0s��m�՗�Kt�Ö�0�ɱ��wK��X�۪x�r�7B�d�J+q�PT@�܍Aֵ���#&�
��k���uk:�d�9꨺���������'p���v��8�p5=�q�7�qm��/V�V�9m�C��c�9
�E�ه�A3���Ӛ�=�������%�����a-�m�gy�.���79)�nB�H4?�b��^Y�q;�։��X�*gM�9�崫m^V�+��Z=�%l�"�=%����n4�w��b �Q�jV]ok6�Y{��7q�^7�2�X�&8����|V�Y���%7��"�{:,��{&�KOC����M
���EU���&��㔦�3�X��q���	�pS8ͮX>#��ɇ|��F/�o`���v���k)�8D�w�>�&C~�4��n�C�1	�$�Ż����c;Mj�5�ٚ�{d�eY�o]�2'!�O1�;�eo��d�H7�lDT%�����.G��2��:A2��ͭм���.B �c��)�I�p�̐���D���س{�ʪ�����7��T�vq&��zi͈+3.�^q�l�����05�9p��9��YfΙ�uZ~�8f��T��tEs,��f�ﮱ����ޝWk�^�-Ŷ���v�8��@�b��y�ָ���ׯ�n/Ca��4��ޕ5Bs����Kb�ȇV�C�_
�� ,��1A#�>�}~�CK��k��M��9�|�����y�i��Hm�o3��`0HIa��
H=�G{�:�`a�چ_15:(4Zl��TS��oߧ���eç�[�f���T�w�n`E�*)#�9�oޛ�)��j�$�w����d��No;���������F�XgZ�x{�}E)�Kq�3u֛c�u�.ۉ�Z<���G/F����Cs�j�(YA�$R@�H�^N9�W�X3�����#9{kn��y�o���p����xHN)���Q�/7����"�ױ]�«Vܛ1�ԏ>�s��/eNm�&Xx3}���~��	9#FI;���{ΆV9+{s�3B2p7���w��ü����X�Ć�y��,��v�<S\.[�n�U�al�u��*s��9�Z��ަviۼ�eǒ�b�C��"m�ڷ1���Y��.4q��q�8����ˢ�Ψ�@��7K��AN���}���ѳ��o���V�3�{/v8i���3�<�q�NC��F{�^���U��q��b����%��{bz)�����Ik,���u��c���E���*���\p�n7k�e|T��p7��v��.�As;���mA
B8��9-O3����*�s)m�t1n��'�x�d_΢���������@�{V��M����"r/��j�O.�����\�l^��a������\�xo�}~���>/��q�ֽ��E�-Ɯ����Y�SvE��n{����$x<�e#}�)�����5�m�+����#�n\��О=�m�ٯN��]��3x�u��^�kЭ^�KeJ�R��h�e{��SwK]Ο
�}��.�Tv'S]v��̥�T�t����/����kr���'��EԼ���>��yO��	ɦ1�{�v�L1U�߶��%��~2Ip)��.Cv��Xw}�z���펆�A��eɞi��S��R�l'��]5{�pg�{P�M���ZI�C
#�p��+��G����^��nv�$On!���_=���B�NM���G��.�{�=b���s<�� ������ �G���ɂ8�F/Z,�Xl�ё� ݰcݽ�=�,��.]�OGIW6髏V9���M���kC%�}7d������*���.��肃��\"�6�:����m�w���#P��[����L�ƾ�v��z;����^�ym�!h� qA#��h�=�y��E�w���f�پ՚�S�}jk�D���g��5��[}���
8�-����Ȯ��8C��;��!�#��.���l�k�v�y=՚���������Ϙ`w��u�b�d�p�VW=�ǟL�w�rFɨ |����d��8�է/��/��e
�Y�7�B��>���\�ݖ`�u�රcj�1H@��oW���;M����sbNܷ[�Y������9 is�uS�廙:;����L��4n�4���X���e�3;c�Q��Ct��]J���l ea2��`h�K�n�zK����|m�p=C��^	�����2gFj#V�8 h��;-vKnҪ���]��97sQq��9-Q�g#^i5�Om��q�%qe8����7B��q�����	j�[4�+śfgG�tm���ܕ͓*�Y�qnr�͓��6��*���i��0C�K>���U��v��+/��.c�v{�h_�,�4��:�Ժםk3���}��e e9�NCvX<�u���.�
ٺyVC=ޚ�2^N�j��s=�NuIձx�v��jޒ�GL�Csv����V�:v��r��N�Td�Z`��箨�"��N]�g�84���D$pܑ�$�ͦN��7c��=��y�ocL+ݏ֦�����-���֓�z{(��1A���S"A rF��f$P�WUս[�U�t��\3�|�8���#�y��a�f6M����lkB�ŧ	G�f��(XI9NrK"rC\e�p�����{g����3��z�0�b��\�څ"�
4\�;2w޽����X�n�gu�Q�Y��8��]�W�&k��V�d�rF���ܒ�Q��wީ����gz��WfV���ǃ͇/���o�A���CDԨX�N���!�*��t�T��9��Q;GHvW&5X,o��b�c��z��#�z���;�E�E���m���7�K���dM�CJ&��G<���_u
~�Yŏ<����-��+�5q)���qӶ:���v��Ir$[��#7a4�fL!T��:��p5�=��Eŷ{�|�D��((F]D��2���C{Z��'#�P�c��w�n��o=;4�\�}H�P~]h�Tۥ$at�ͮ�,�/.���O���m�$:ݕ��i�g�m�P�J�N�>���9��T�m��v�l)4Y\�s�#ןgm�i��WSgk]�t�璦��Z���v�ȼ�N�\��.�S�R�yWi�:�
���G��"���)�XKCQok�,!���gޡx�k�-�VΎ�)^xf���X�N�
@�<^�m�&��$��p��.w��8����^��2�9W�ǰ���ІB�W0A���5k��e��j�o�
�ZW8[x��ȭ\��(P�N������DE���fz����n���'/bn���������M��}��D�$I���p߄9���A�j�\>/���[���� b	|}t�G^OGg�ұ�yG}���`��-���|d�Y~ݛ�Eז���E]e�f�oNk���e�n��K��H��������߲>U�߸���[���ZK��w�WM\n�Ts��\7g��=��틆���e�f&#j�[�᭕L�ߍ�ˉ�����]��S����ω��f��\�����8����x��\E��PC"r=�mn��{n\�	]j|�+�{t>�ԅLx�(���qu���н%��&�W����,3N7"r��+��Mݒ��;�\�v��"�;�&�.�l��v���G�#Fϼ=����Ɠj���l�;]`�Lq5^z빵nѸ�W��Q6�gvYag(9����]s�J*�:��ci��	��)�y�
C��������(�X���q�F���%S��HAw[q��"�0��ΪZ�2q�g�p'A�L�rN�i>��^���Y�@����J$�7�3��Ev�ϝ�*,�t����qO=č���\S��޹v\��;G(��6&:�):\�۶y�]v��t��>)����;�W�]�e��6+������d��%�\$�O�C��u^�+ײ!�I~�n%	�%�oo����qE�������S�(�m3��m��we�5��ظPe��
�����H���%���J���5os��c�X������ϝ�{&w�~����f�����h��+���>�@��5e�E��9["��6�N��sVc��DAj2$��gT��=��	�@�p\1�q�q�(w�<u<i�`/h~���z,5ck}��Z�D���
�M xPsE��F��p�(�P����oF޽��1�g`�vЍ-�Xo���C&�5�k�oU�ޣE�NT�и-�B<X'Y̥%+��ҏ\��4��//:�r1Q�� a�9W�wJ��J�1X��e������k|��
�c=�R��o�]��Ǫ�-��-�8�����UZ��wEW ����:�g3��v�
�k[�ii�S�P�O`L���nX�ec-���+�aa�QM\�f�`�H9�k2��屺;�.�7'wo�Y��kt�� �}XS���əE(U�f�^�j��Jn��w�	��B�v��� ��1W j�^����9q-�΢0�@�F���2�[�o�>��3s\�w�輔��1}oi�	kͽ�EU�0_K�o.�H�L6m��MiM��)�[�2)��Ps��pL�y�p�[L�nT�+
av��OWNj}Lۼ��F�f��ʍ�gt;�SQ���SQ�������x!W�����΋E�f�)��E;ep�V�V�oF�����LTk��B>�!^d�t�
� �0k� �z���Lc�B�틚֖gF��;kX�Ftox��C��0���3�wv�1��]r��n�Dw.��1q����rv"V�hWu����7|졗')vb�{�w�]Q��t�� ~��I�](���W�(�����F�^e�r[1��Wl�&D��"�zEԡ<DM�X�%�sc6�XT���;ot�/�j��b�+N�Ȼ������E�iI���Z����m-�V-�9��1sr��5��֕Q5�m�^����I�Zv6,)��d^٭�`ym�R��i���݋B�P�z��u�O��n���\2��b{%r=M�9ͺ.3ܜkrtfuj6`��Z��Ya�b�E�-vcb�L��h#�&�#9c����<�S��n�v�����ͨ�0C��)&t$5nv����G��Ӷ.C.�E�%�ɣ��M��̸��v��F�#+�����ӗv�2��jן%taT*�h���I�b4�ɢ1#J�F��	̛r�P 6F�)c3p�nx�3��*ŶR�#	�����)2"\��m��V��f��	�r���.y�mJ]����ڃu��0�m؎�\p�Y���9ޱwa�m"��^�e&�
ѹ�6fm`�vbT"G�����{�9�0W�&����ن6��9'�s6儶2�xK�YD gl�
D���i��Ǔ�دi{���Hۈ���P�U�;ء��tu���.�cB��2�c�86b]x�6��ni(1��n���uMm�c�W`"�-Ɨh��5Bn-F��uT����h��aY49L�Mhب�^��腆3�\���n��ƻ��i�{{�p��歷rT%=�ƃ�F!�	�0���.vwG19�Gi�,t�F��N��y�G�.�,���B�bWK�r�r�G�q�6���(k�4vݏ��b��L�\��=Hw]�"&���r]�Oz�+�.�ݫo(;g�����֦ݴ۳^��Q�l�x��ܾ9�7Bm���z^�n9rem7:fz�4;�������׵���v��g�Lk�K�/�z��:�α-{�����Ͱ&�㙵�iX���۫�u��8����g���"`�%1T�X0-찄n�^�֝*UM�p5��6�50����j�Ӡ��<�9���Y��9ӠR��ͮ�����dm�mm��YͬSÓ)mEqV{"�7N776����=l.�����;-��+sҝl��X*5b�;�ͅn���59y��)��c<=�:�,��:���{3!\e�{i�� �<�u1u��o%τ���@�F�v��s��dds%tҌ�MX�3]��V8N����v֏�<p�,,�t*��y���
�c֍Bm=��'nDCk�z�m��]�)A���fx8�k��7���^�ٜ�K1���n
S���!�����nE�ד�yl;���료�s3]��B��h���;B�rj�gx�6,�8AeJi�2<X�~W����y}1k�-���]��\��;�NY͌=v�y\ګ����2{�x*y{Үڸ3z��˖�z��b\�}��v��&�/JV⮲���P(�j5r��$�J�G:��F4��ֽ�S�ڲ�Tw�{qm�~TR]j%u��O��܅�#qFrb���W��+:��&WSk�ìwʑM>$r�"�O]�5&o���x��$Z��\e2�p!��X�I�F�r�����d�U��>��� ��w��OP��7Ž���&�mN�{�BH�2B�rH�U�������2����ț���Z��!����y�w�&��ݑ�����p��Rс�x$���*��gmF4Ʌ.�F	��ۣ��=*re�Ji����	�@�{�6��R�䃮�.N/�;ǃ5n�e���Ix�U%c���|���I�ۂG����������!`����� �v�ۺv
����?[[h�=FD6uZ�g7$�ŷy�\g���w�U���=�T0�ˑnwAPj�p���*O�+Oշ���:�Ђd��w�	��6�g7`!��,�P�	A1�/+�z����赇��Y�cM�������|v�8Gk��ӱX{��g$*H�9�A:.a�k�t�qS�f��=�5f#q=�sהp��������kg�P�3��BTNˌ�׃MUv��Iy@Q��Ě�:�_ ��]r]3�F8F�}s���}\|Ծ۝y�X�1��;s6��j��m���=��uӘj�����X:9���Y�&J���;��J��iG&��Yྐ+�;̺�F���SL���K���<�ёA��7Fn¤�L;�e���&�j�;�$�(����XU�9�R-8tS���.��5#����3ܽ�Ԧ�&����n�˽���tʭ�>�|-�Uz�i�|�yЭ��]�6�𓍊Kc���sQ��sn�&�ۧ�E}�a#D�.��S�/�t�F�X*������+���ލ�^���Uz�(�=:��z�<�&��\r9+#�E�X�G\^��k�W����{s9g�/��OR���ډ���P7j�
0���� ��EI�2�͋J#NЧM!1h�k��˫���^:��s=�;"��`�V=eC���2�W	r�ةn�(�JS0���ѓ�ո�;S�6`��n�ֺ�hj�sėl����9J;B��-==�.��q7�^J�n��=��K(�xf�mEn��fd��d8dJHo�:+�.߮J͠�����Ne�me�ol�[�N��F���Z�@eW�]�v�b/i10a1��,J�Pb��}��;��:���;��f�;)�gѻw: �Kڱ=���A|=�Q��rC
nL�s0m�Tv�_�o`�����A����Z#��U!;~��b��N�q��x��=�BuzYcUu�`�j���'�����������\ :�B��M,�����I��{���v�bU�e/'L6$aIqS�Y�[pu�Y�!ܡ;wt��z��K<��{\ d�=홨�y}ro��~rЧE�lX�㮭a2���1�l����=�w<��e5�[�k5s[��]������)�z�Xƞ�����=���31���˩�z��b�*O/,i9h�H�$�eY�>��{V?5J�t��a��ʌ%����e�/���`g_{T%�~�������I�Yj&�qïs�R~���"Ȼ���Y�,{g*�fN�3��i�Sm����&	a0T䍹�FR�Ժ�I�.�̞�W�M�Rx���R�n���w����d͞031\	(�q87��gN68Ɋ�ۢ�e�I\�GvE=Bqy����Ê�&{Em���,��,��A��"�aX�oP�����V9�:�c�q������,����`�, ���^��/N��9ۯ�j䟫�=tVŋ`:�� t�z��}�j�֪��2��jrƬ�=�'ny�|HO[��ٳƫ��/V�yK�r��=�<�s�-��3���ܜqӡ4�92�7M�b���)�4�hִ��%e��*�hS��9^L���y!ˌ`h[��Z&��1�Yf��N�q�L�8�Ҳd�P�ˋ�<������3�i��JK�o\OP���k%[�97k-v;.|�v�'b�e�#ԙ�9(�W}��}��LE&7a�K���䡟z��S�.�ttt<��˦�>WV�[�IR�y�s!y��gԓX#f$"8����į`K]Ra�}}��~��XMm���C�݊�,[�z�*���x}���j���񶡍��G醝3�~A�·8#�Z�\ͺ�*U�4U߯*L�&V��a&�C���Ɯ�M�"�+���.і�e�X�[��7��V�a��{�Ѧ/��k��C�=���1?�-R3#��	Q��զ#�jj�̩����l�1�)�����\]J�7d�wM�f̡gh1�2wr�{�7��I�j�Wc�����cgu�kv��U�[wi��J��S;[Lnd+����\jaL��U�%81�����W5�jI1�����`���*ZtJ���[�*�U��nå�ؼ[!�d0TnI5��+���V0���K"2���b�kG}][�����tu�` ���g>w�.g�.l��5����*c&ds�W\I��w:%�+z��$.<�j��]ښ)oggY���̀��uf\�v@³�X����U���c!�"NEZ����}s,�,U��z��y*"Vy��w=�����;�^�{~�׵7$��
5N�G=�kX���b��i��։�=���e�����ז3�9��&�׶<�x�z~p��MI)9-U���]�fq=jMCnzU�dd���N�v>ŭ&���Q+��˿m�6��K{ucMb�Xs�J#]���x�6箚,V�4���1�Թ��{T,~�к��+�6}�=ZO�����Pխ����/;Y��յ4�����Yj).I�����z`�����:�K�>/�آCo��R�ʭ�|C�,����^ĳ���H�BDpH槗o^�yk�Yy�9V�S^�;F����,�8�2�׶�F�;#�	aL�R�7�k/%�2�L�ec�\���`wH��1զ����o4|����	/:f�e>�fsyЅV���Ҝ	1-D����ʥ��U�2U���o���Y��@J�q��t�{��_s�&"�qQ;;���l�)�s�8(��	�&ܙt^Rgs�mc���Y�(� Ѯ�c��M��~��b�j�p�;���R�����Ѷl61���C�F:D�:N9޶��=�PO���AǢ���ms��ZLF��r=�����!����K�# s�ފ��;0�U�)��H�e��a����EL�Xr���U'��{.:-$=�b�"]<&�I�16H^�Cbc�hQ���7*�|�����6���ɂD�.I�Y���ʫ��]�0�v[�~�:z&��|*�n����{�[�5o�9��b's�8s,��Ѿ��ia>�{�7��E,�����@�����	'4s�u�|�]���z�9�v��
ӄV�C*�Q��̹pt/+eܶ��g5ӝ��x	���{���Sz�]� ��rM��c���|A��J���lȔ�f�E�;�~���߭�F>]7��J��w4��w��f�~3*kq��b���6��T2/�Q4�ݳ�a�f��ee[b�M4���8ܱn͹:7g�ˇ/9ə�
p��A�&�rZ��C��A�i�tPDY{j�'�au!��ޓ򻽭A����
HHm6ʐ�fQ�-���I�gȳp��L*�H:t�o>y����G�"�/N�ߵ,���ڶGJ�������/?_��	�*��z�z���V{v2�����!����/aې�fz�n ��������N��;���нL�ǹ�e�d�y =��;��T�YD@i�]r���37�eX��)H#�7,8��v{��DP���ߘ�X���g3$m�;��o�Jo���ǜV���nn����W������Fři92�i��E�P��a�ۛ[�%�ů}4��9#�T�2������j�p��Y`�6�\0l8An6⮍iu�r�Q�/[����L�u-ĝ��X�7;��磓#��ox�b�_n�׎�D�*"qcsT��3GV.ڶXͰ���Y���;u����T��uzM��,sÇx���,��uo]����q���8�rݩs;8�ւ�����\��<K*���Y�7�T��J�[Δ�¶�� e�f����v���ᝋ�*\뜸�}oI���]/]a�p�aF͖�m:�2ǧ0�8�2D�l���ʂzw�;X'�~�J�Yէ{|]F�u�s���>���hl�}����"I��9N.��W���ov3�9G�����7Y^cs�dNd��A��˳"l��֊F{"�J8p�Pr8�Y1���=�$��y�va@a�	
���tl!Ω[TΞ�p㧽���Fg"�)%�
.j66������97���䙕jȒ������{�.b}�����,���C.�s�k���c�U?^aGVWRk�W�����a
7�t�O�o0��k�5��cC:\��u�v�����ql�&J1>���Ɩ��1&ܙv���]ƻ1�{���M�o#T>G�lJ���S6^�bHά5w��t;]���&"$rH�Q�v����ML�Sj	n�.I���#��Ͱ��lLӄ����2�3�z��B�%�F�V
�"�T0ڸ�u�FV.�gj�B7�������gC��g���}��W(��=	�	Z7w<�%���Y�X4�Q�`a��V�?y_��7?J����m?���n9���s�ԋҫ%�n�dI���䨳L� ��c��&c�Ƞ_W���9�o4�z��\��s���t��pd����5hY����xm��PI S�8}����}�o��H�Obj���?Q��7R[G�ގ�xm��ά��+�-�d�Y��qu���Ye��;��xD���n�z��l�3�D(������t^��W}t36(���ڳF�{:kP{̱�4��z��G}�l뫂z�)MHc�(��bf�מ깜�'UW��Ǫ;���u�X�{'�;={6+���ח����Z�ot��g�RBCi�c�Hh���0�P��;څ���wTJ�?c�с�+�F�wu���r*Z7,Q�<����B��j��zC=ڵ�HZ�:n�<�Ze��kǚ#��++-g��X&��,�]5��7즎g2�֨t����v��Я��uq	�Ioe,�+�GgGp�}25�h�p�wwk,�(,GڔR���l���6^�N&K�z���=�ǳ#Lh���ݺ�Á�5�[e�R=���l�R��G�r�&;fp:D|^�+m���mi举�3bҎѾ�or�&��(͔.\2����5RE��"�ݺ��ݙ8�ЕRՂ1����1��
�Ѳ��o��F�jY���w=/�f��W{]qo�ʶY:���FA.�1�B��1<�hí���˻\�e���2�����۔ʛ�&�6�9�x�^����y�j�U�j��\��`��)�]�ō�n3O����Z�|֪�[빖���a����Pwk{���p���N�0̬��EC��,�ͽf���R�a�f���9�M˛"̸/�Y�ulƯ�&�ن�\�;�uӒI��۠ 7�l;Z������oF���y%�D̕��HI;c+n>8&�����ۡo�q	N��ʽ�=�:��Sj�Z��l�{�2�� �����æ�<�Yp�z����P��D*1�:!Oek�x}Ʊ=��nM �=X#.^���v�hVw&�\��;r3��w�yek&_j��F������(�!
�W=�UĹ���D�x(���i�]����j��"g)�l�;�K�͉b��`�vd���J�ݩ��N��m$�ux7��^V��o٧D��n��K�� L� J$��OR`�{�~%��N���򠋼�EL�/R*�Ap抈&*�c�;�6��I�)����"���'R�=�Ɋ��Xw���]���77��Kz��@� ���Ŧ����������3c-u#�YnI�뛶�q3�y�ܗ4��s�h�,��3�^L+r�$N$ �N
ɻ(vza�ARƭ���	
����o	:/��щ-�-t�;�GE��	�$���RrR�=[^�c.1l�#Bݜ܍���x��ӝ��ˎ5����j�l:B.Uݢ��Q����qH"q]_v���<��׽W3�א����!������Ԓ~~��lC�w�[,�L�����b�,-7���tO�L��{�Mn���M<϶
⧑�y�}^��C��JT�td��K�GK)̙ջ�n*c6)�tV�[�'J�6�q]e�\k�v�,�1��m�
���o��Wk�GR�M�5�tF��a�=媞=�=� ������6�&�(B��h���b͈�sP���߻��9۩�wi�=yk��f��Zy��'f<s<<�mr"�Xm���.��.�ͳ� T��%R���X�̝�qIBk_�������rξ�z��!��	�nL��(�����Vpx���%�w+��������Mdڔ�=e!5�v؜��T�wG_p�G1$nH�sf�y����H�=��є�=Wi*9����%�s\��ln[�(5b`J�l�#n����ȧ�}�]�ݭ���<�����8�ɷ�58FG��&��گyF͐�&2�p�d���w��ړӰ��1U*Y�5t{z4b�퇧|��*��-W��6ʄS��5(:_����	�}d����J�B�,�*,����ەa�ʡkCr]���)�qom���N�Q�Ĳ�[۳*�Q�infv�a� �[j��e����R�vx��n�)z,n�� ��G\!��๝�;�Bi��WV�f]U��;���V��n�W��;K̹D�1jF���ۻ�c�"=A�#5�	��l˭���Φ]��VƌcR�!�N�{	�磞��dx�;��r^�����>8�Zr�i8�Y�pG5ک��:�:Yf�(W%��fբZ� �e�۝�!r]1t��[k	v#��O����m��<��t=֖���u�@��J���R@�#qo�%<w����5��w���������Sǈ�����,L���Va��H!�%!m"�eʕlPS7��"�d����jkC�t�����W��!���D�s��%��iA�}$`�$R8�MI*�ɂ]��Z�ɾ�������LtC�(l�VeL��c��HK,��q�z`�B*�wG,9=c9�s�8�k�?P��E��&�[vD��B{א�o�Оļ�)�R�nI�{��o���Kt2�D���z�Lq�����to,�����<W���1@�N�1;�$*�w/�6����-bm���+˞qb����-�r<ǯv�_}6W�����<�L�B��3��K�����T�䗁�=�1�u�+�^��r5	%	*A��ʹ~�����U�º�l��n�&%D�{o���U�az+��VtY}p�x�fj�3�+B��=�㨞E��\N66�Xs�G�a]�Y6V���k��^O�KɃI[����,�
��/l�a�Ӊ NX��M�jFdn4��&�^�q:�#;;^!�{�������[G�]��Gio�k�ɬ(ᡵ�ҤTLFZb8B�"Ya��x%R��R���#a`�뵸�~�6gIE��&�tp�];�x����yl��gy�&0)D��A��ŷ@�׷�^�9r��f�Ⱦ/^���%s`M�����d6�E��vxzYE3M��l8�|O��DlKbA�w-`��B��-�� j=n6y��Y��Ψsy�$�S�o7�/��y�^���`��5y�u��ݾ��{BǠYݚ�K>Re>�Ňa�D���㽶!�:����P�)i�@?_b)�Q�����8�'��\�H�wS"W"���S&�D����JE�
��o�?,�mI��ͧ.x_�OR��=t��.}�w��3N���ۭ%8e���e�ۚ!u�P��I�e���^)[�!ZL���vS��m���;���æ�{]P��'�����ݳ�h�jr&؍ɚ#�lʥC�b�>-�k�ۡ@�y���J�[�wǽ�Ey\�Z�T�{c{�tw�>��G�HL8Tڂ6�tp���� ���M],�<����A�J�1�\r[yHq�74귷�!�Q�&�RR�����A��R8�A�{x��qMhL�\a�g���R�.T�ˆ��z;/
8�������{���q���\'r1���;��%��1UP�.�: �q%�	R@؅��Y,�i�[�C4����t�u��*�����z�
��t�bŨK����G�"G����H�G%� ���7��V�vv��r��m=Bik&J�N&��m�Qi|�pO>�CJ)#�6���C����7;����S��N�w�7������zQ����߱�!��0�E�}׋2��p!�8�0Ĥ�߻hu�	a0	�y�9]* &�t�X�r�ќ�慒�<�Z�=��7�� ]~j8	����9�C��`��=�����:Qe΅}��T��,���l{B���;���zN�ty~�O�RV\���"k���'N6�{8�qQ�\�wj�6�=�����\l��)��*$��39��59�}9]cC�#��D���K��t�S�nns�z�'��X�4�0��$�V��7�郦�fL������%�2��U�~��;����6��^��y�=z�}V��@�n0��G�W'����4�v�U_�$a�h	oKk6X*sS+GD.��*�Q�rZ���[P�c��R���f���Yࢩp���X�ߴZ�E��{O4��Vxx��%���	n��F�+�=����U2gn�/�﹖�����ydr=�~��7�[��2� ���(Z-%y�f���n�7a�W��+|"�O�=�}B�Q�'*#�O�W?���
i]N�].�7�ֽ{@���]]������{v��F��Աk�=�ogB���E���p��U��fFh/@J��ExK��^�r�x���6���lp뷄$塭�>�=�{Y�k���̌n7+5�r�ўy&ϟ]y�_[�Jx�.�u		�`�Z��֒Y������/�[	�6�΋pK����t�'�;"�c��c���ε҇gC�pݭ����M��&���c4e(k�3TbA�nf�\ru:1��Yc�Žr&�"�t2]e��s������b�;�ڝ���ܘ��
I��N���OR�iתx���ԅ5NL�y��o�Q�RS��=f6�i�����(q^>��X��:xgN��K׍�r$�3r;��6�W]��^�h��;��L���A�xU_L��ۚ��C;Р�����Q�=g-&gW�P�"��u����uO�M��g��c9��uj����/˷��M>���&6Z�� �RH��3�]���FV�5*�:6=���ݙ�{�k�����nxk���x򷸋���C̦���ى���ݹ�`��q�^�Ups�s�r=)�M�wQLT�6�����UёQZ}^x�!��dOo��]]8���{3_f��b gC�J�z��Yl�b&ĒraR��/mΠ��f�GD�n�N�J	�tVk�]�����I�K���m�j�����QZ�-�媁��u�m�qT��'a�n���\��u���=n(�^b�X�l@��PI�d����Q��GLF�yv�]ey���h:��i����&���=�x����PH��f{�,�&�I��E#�1��Q��v��ޔ��C�U��/f	���[�*�eΚ�0�&���0q\!�G$)�ܒ�r[��M캫��Љ)q;[<jr#=ʝ\���gNL�Q��s����|�u�S���]٩b���9v��=uvR�����Z��벖�W2R25$xB���Qn.��,���/V��=�Һ6�gԎ����k:�=�?9&���Q��hlWly{�t�]�x<�M��4��b�^��cD;���4f��ZE<ۤ�o�4'?�J,@s�H��\˷}��v�UN���J���]0�6��g�7^���θb�i�S��w�,*�,��c�ۉ�퉪��=�֯3+*���К�җp�ך���j�]=�,:�����U�/�}^`p�č@����`�����x��&f>Ź�)�VEe���n�� Q;��w��{H�ɗO�����d�B�E7'F���ߥzk$Ժ`#K����wb[~]Y�qg2�����o���vt������Z�t��E��E��j��yrY�J�6���:�7��I�6M�ה�����Is^)%3���E����T��QM�������wY�n*�m��#��;���c�$���#Qǻ��}s{���ӏ���~�={�ؙ{u��
4����^�6���ayT�\4i���P���`����h��.R�N�zc��R.���p3��в��^Ҥ��(S��i18�����Q��XKHr�,\�-t����F��J�����͜���<�y��F�Ǚ��:��m�x.�7b����TL�@�_pYp�;m�笐���8����,+�_�gR�ݝ́Ls1��:=�"&12E����v�e���ǻ8��O^6�1p�/�#��Taܞ+M6�]�`��#�t~���}�u�yn�u8�=�[]��&sVc,�[T-IhA��f�Q�L����'R&c��w_�Qi���bx1����`�-�ޞ�$1��t~-K���0���k�L�$m��Q85�N�ߎ:n�EnP���rY�ŵ�;�l�f�S�z�/i���RYW����Q؉'Ffnn��������)��qyzL�C�S�e\�H��.�W>�"��oQ�rF�lƜw�����w�T����z���+{���V����gLZHK!X㾗�|N�Q$
N#�{�C��V/%g3��hr.ӌ6i������6s�z�����S�+���=�j�uT]���d}8��4�����"�A�z�Q�˝��c�fJLwu��.=n�&2�"��{�ً��J�	fX��d�Ѯm]l}�"���ƫP�9��Ȧsq=����Mc�t3/w��H��w���n�t��n�"��U�X�`e ��ͱҕyq9g�oQD�L;�I�ۚ&wcy�o#y�N�����|�;�o{+7��7e+4�Z䄍�B�j���r��u��kx�g��R
��;��!�J:�kL��VdFR���i��Cr�����4�K	cù�����L����Pu����NV*ְ�z�n]nĐvF�!�@NTt7�0iS7�h���S��VkޛQ���V�ɸ��;�9<�� |�@���K��f�s�u��%��7��d�X�e�e��LQe�ǳ�_VB�u�j�s;�d��s��_$���n��7۬g`O{#������C����T��������w�9M�Ek{)�mm���d�
�B�+�s�:�N+��{�����㝫[�F�5_mSm�v�;�(�����Q)��-��Ă�Yckg�d�ה��rhF8t�MM�C3�=:�k�co:�љI�H��	�ᛛ��*	��vZ�76��/gAE�D�Ww�������b�-Ǯ����N�_Q�r�=�n�{;In��D�q�1���82��7x@a�܃t�j��5�3 ���!e��{@��:�oOp�/H��_�t�Yc��W���rs1�+��ԨH����
Ţ��Yl�Dd�	�i&ݪ��KFL%ΥFlgakn�-���9�S�]���!4�<����0^{�c�'6�|�����\�ڸ��Ù�m��Ec!4`�U$nE��j�#\X���ӫa|k�%�[ٽ�Z�ک�֐�V�^�]���Y����i�:jy�xv����U�n�u8�ݏf+�pL�ff�M9�����q�"K;��:�W+���&us�8��Y�n��Wgn6�ͺ��V�\r�a.6�Kz-R�^���(��%��Jϰ�� �;m���rm��.��6V���"y��������٪N3���;�/#�n��p�]40�36�"k��Tk�񱻓ϛuI�D�����/�mK���<�N�wm�<�@���W]vs�A���鳷(�ٵq{��6�u]��N��p;����hvk�_�������9錈���/+^�v�:ye&���f�	lK���u�ޞ'i��.�N��G[������[�Eq�]<nۃV��_\`��	-��иvcy�
2��2[u��ܮn5�e��q�vW�06� �q�3ŕ��2���uO[j��]lJ�X��ɹ���r�hu��R���U�5�z�N�L�@1�av�d�l�����C�e��bkְֱv�̼M�qr���^�����rZ�#�2�r��2��[:���!`Ù]m��݆+v뎻sϮ�F7��(��(�1D#��Fᕶ�\a��BΛbNy,���ˤ6:{����e���QЙ�k��ݝ��'gs�l���Od*�l^�@v�ۃ;��cJ�����u�8ѽe������/�v��rs;C�>�v��;�ǶZ��e�	�&�c���o(P�y�g=7�לn��ѥ)���r�d�1ŎnFGn&��¢F�QЅ�ʌ�(9�8�8���D�M	�˹�ą<���.�k���w	pw]�1�)vV��cpkCu�ݝ��L����p�NL�<����u�{r&�^��q��=kl`���B]�Hk��9�t-��9K�c�p�.�hz��]NE�G���������&b���fC:n�Ƭ�*@�-[7	itf��n����,[.�[�V��R��+n٭ϰq�n���l�i���YF#pY[:�F�#][1�+\F�O=.-���;�kt��Ϯ�5��ͭ�p�Av�����{WC�q۰7�xC��ͽ��x�nu�S�b�̓-���X'4V��smԳĊ��f�q��À�t�R%/e�<i��]���X�ܒFܝɎ,��ەOz�^uyM��z�C�-xHya�tf��b���nd�\r8}���k�'�U,$c*+���V��z;Mͧlr{�jJ��:}ްed�שvT@��x��,o�d��P�Lm)fRDD4ן�W�y��5I�b�B����Gm�aq��}�z�樂*4gNq�n-�[E	�cA[
M���淲v�3���6�v��R�=���e!k�C�_�v���RE厯x%���25!���UBy��%6��^����M��ʜw�({7g��2#1�	$���a[��Ԁ�)4�X��6�S��洴��4b�T&�%�ź:��K�+�,V�n����k����~�~�媮.�]з��ckD�莡�/�$��!s�L�g���~�z���oH%�/��fN�R+�g���'k!j��e�����h�9���7����e�ǧ�׮0X��3�kk��Ӳ����R���t`�۩hqW&h�e�=������@������\�y�w���_}�巽���S}�_z�lDQbr5vEf������ݦ�s�V�Ik��AR����{G����rm���w+�v(��H8r�ҹ�	�]��	�ďo�x�L���]~z0�t��%���M�>��r7��")��!M�㆏�-��]�ͼF�EEy��#T���o����]龙6�^]���<e�>����l�P]�t��e4�-b$am�i��4+vK����b�8D,�X%s�RlBb2HS��Z'��~w��R�'�{��os�&iE���E��*w��ޝ�[F}�'P��#jD�r,X��zxf��qh�6���/1��b�ɼ��^n�:�Ղ�<�Kηwl^�*6��K����#���������{U��?i^�:J�yk6�l��N���H�l_�x�՜��yX��gF��c�U����{�dM��͔��5�ɽ%��Op�IZ�B�� ��g��8A���-r@��I���%��}`fk
��qԱ�3��M0�~~x+2>o�O�8�x��Χ��u�6�Ԍ��7�K`�ˁ6"7�׳|g�f��L�s�����f�RvG����� �P���u0^[�y��w��(L�1�e�����9�k�-Ø{���.��E�n���]f�։�s(�M6aAd�%��ښ+��Rj##_��YhI�U��#r(�njd�^ڪ�\�G?�^M���-��o7Uf-��u=�~W���W\�M�&�jJ�9,v�qO�U�#H��1�<�*��Y-�JFF��LPWgx+��{�B�^�`�w O��c=��Rհ𱽉�d18�Q�6� RBs�n�"x�U'�my)����]4C�>��u����9����R��˝1-}�:ꤥ����S�����OE��E�J���}Z;m��i���9&7[���s5�;kU�N>�TT<J�NF�,�	N+���.<��{-�h���-�7;��٫���[ Z��y���½��S��{�;�:�\��S.�6J�����i��&�E͌8��,G@�r����.���se�c�ɹq����{`"W��o6�vρ���2_Έ�c�����t������N	$��NM�8����g��q{l�<Ȉe�1sCr�&%��(3-�������K��Ja�(i���Dz8H.�-��J�X�{�^Y��_��_d��RP��c�'&Ov`�{��3�hC{s�l����j8��m�-�j��v	Qeduq���E�)�����9\�w�� e����Ԉ�Z�! ��o���Xm�"a4a�}�񭎊c��WT�T���ѯ�u?�(R��=o%� v9���w���d6�j��or��^�َ.��M0�m�{����<�rm�}����l��-�����O蓇vs�ۭL���A�]t�7D���F��k��t�5]�c��1B8��0�Qڞ)�fsj{IFz�^�M͍nzrA�ۀB`ӝ��#��m�
��f�G����)���X�vd�BWW��xCFV��Q���hhl&�Z67�f-ع�\f�����v�P��60kY��:ȳ�E��&M�<A�*�,�RԚ6���,Bvx��3�K�F�[���Enq[�عƲr�7\Ÿ	*�˖36䭖.��pk$M�6�"HZ�G�~!�|���Kx瀖����;l�6�Q�����]��.��P��M�"pe�j�_��,b!���*���b��;7����)�zz��)�}x���Ʃ�2��4n�f��e�S��c﷉��-bu}S���DS�=.
�E�ξ��b2�ݔ�|a��i���X<<I{�y���dOt�lsN�	-��ʕ�7����tg������dl�H	�8�n95c�;���ɰR��/��}`���{2�\+2�����JAD�iFO�Xe*�9��%��n�r�{��4杸��6��ۛ��\a���6P�`��"q]�͗wܯ,9���̅k*�޹Q4#;�nj��v��~����"C��ߙl�
@��Cw76�x�����t52����P$��:��*B��֦f;�1�wD�����X��묘�-��r�K��a��v/	:Kw��ȅq1J�Z˒.������ÞV;]��l2�0�t��L��a�N6�t�7}�I)aݍ���9�LNE�}A��7vic�ˬ���a�P��!������'�aJ�K�4�RP�W�oW�𬹳a]�W��67�A�}buSݚU�vx�yB�PƤ�(��.��u{/�旻�jH�������m[ŵƧ$HW��4��^�F��l��?7��姚�f�d�o�ے�Ҳ����:���&2�ۡ�s�\V�uۦ7Wg�ZzKk�J�h)�j6x���cE���ܛ����
�òW̥]x��Z�%�GI�v�H�锥}|J�AWd6:;��&��\��8/'��zy��y���
�P�Gif��#�)c�7M��! R5"�����{|��V:�D;=�����{�=�F��@$����}ٗp�1T���;��G@�W��k���9�כY�W��f�,����8���	�U��R���Y;���G���6!.�F@ԋ�\$�롪��X��nW���^��[�;�\+j�����{�������:��Y���k�]��er��A
槌=];i�]1u��?_	<e}ɫ�4�3z��czd�!�Y۟}NFg�wW+7d�L�8�Z���\r���[9ݸ��h-h�S�kZ�P2muL�����h=�"�َ��k�j8�!5�	�G�!���$V��
�r3����8\Ddp��C{�E�پ[�7�L�O���$<��c������ΐִ��7Z�w��!B�n6䁷zl)a��b���tP��ޏ�Reb�[�N�4����e}��]�gtp���1"��G$7��>J@Y����x��U�]�1�A��J��r�rl'�f���Ο{M'�ݾ��j�;.�^��*�"fY)ޞ�6v�Ӡ�nv����X�ܛ�֩�^m�2��,��:���볕V���&�fBXR$�pc/;���d��B�����u^��؁$/>^����h��)\O�c�$?_���ӴNK]����Нp�Y�@�l�]�:��!k���n��N����6�jI~}�
������3��|�ο�D�c��uG1PU�|�0y'�����"J�6�<�řc9�����lNҪ��z��{��~7�����u��{��m�dC ��n{��&�9�R��Ԃ5$��5i��VF��Ҿ�<s3d\.h�~2��֩��3���P���G���$H�.Dۏ́2Gnq����ݫ��{;�2ti��h=r9[�#�?IV�z?Vm`�~��`�,$��0�H�ܙ8���H�|��Y<@j�mZs4B��ν�m�f�7aD������c^�t��h�݅��7�@����D�ӭ�O;ێ�ͷ�,ޭ$$�YpQ�ľ�s.�2��qn(�FsNG����O�Zzt��ڳ��JI��d�����$Y�tb�f0u����!t�.B��WXF5l��n���a�����pN#ϵl�'H��z+�1y��R��h�:�Ӹ7>!�i��^{W^�ۨ���vw`=ut[y���q�DGmx�L�f�����W�Ք�7)r��HʚQ��H��UmT��!���nUM9t{6�8��^�#��*mŎ��`;b6�K���dqNB������8A��˷]��7��̉�h�3
r$�P�ڍ��r^�`�5�Mگ�(F�<E̐3 8�|�����;��"��\ͼ��;��"��8	��]\�o+���Y���z�K6�߮#��'�=L�;������`�5���]u�C��#��\qI��R��&R�uuxS,��+@;
v���_�M>B�G��~��'���!qۉ�[�
6�1�.X�0w[�����bk���f�	瓭T�/-�H*�,f?w��<����ER+�c��K�Xմ`GMHv�5�>�ǚ~�M�=��o�޹��P�Wr�n1�=Ƽ��NQ���-�)��+�H��.9�x:��ݞݳ��2l���W�v�bHK�5"�(��ެ�,B߷��Gvw]tNԓh�E�}l�^��,b/��z��8R0)��W)9�z��Z��9������]��Y�4�{�H7 "P��
\�,FF�w�D�V���)�JXqݨ�qڛժ�Vtv�ɵ�+�"�L�#�O+p���x�4,ݒ]C��m#$�Qܙ�q�E��ԑ��﹩�-�FD�����##��,���Ϲ1Uk�9�Ҫ�{�����bfcp�k����s��&��?W�G�FbE��0���߸-�YN�v��Ԯi��{ ���8L�^�Vvl�^	�m�	R�)ŒL���~�lSʤ��L��FeA�ou��	~�3s�d�x^������&����EP��3�NR�Ê� c������3<�׈R�n͎����.�P7mEFI��쯟���Ųح=�ˬ��^"����q�H�2���VM�t3��F��	Q7NJ�SU��0f �#��{�;�zF�)�S9�C��۝*�0a`�Uq�p:��n���) Ɣ����\�E�E_�P{���=����̯��vW�ɞC�W4��2���+���p��e9���6Cڳ��)�����
�0�ͬ�8��V������LfI�s�NL�B�v${��r�|�-$�����՜f�^�E�_ì��}[cT���ݥ:��N�ctJ
��A��
�k�(�,m�ޙr�[�n�%��l��؈Aћ*.�{���7ٳ�!ژ��{v4!�5�-�w��%����i
9��J����mR���:��s�ܔ�b��i����4^Js_:2� Ȩ����s7�y(�=5��4�p��ڗ�޺gHgN��-���l� ��.��غFW�͖�^��)M�3�o�2zo��Tu����{S D�JM��D��we+�Ƭ��ٹq�ۨL���%m�ԩe�d� �����n&��^�T��]�1�3v�j��Z�[]$r�'.�BĬ�|T�d#�f�ZWm���wq�+w��dY��	�א�旽\eMU���������v_\�X��h$�>���\�wy���v%���՝�Z���l�XɅuC��`��Ͷ&a� ��NΚ�l��v��f��Q����$�Y"띲T;����J�#4;�G���4�ܫ3��"Qqʹ���6Cֶ���7^��'F��Oq홂����*i��]]��ö�9��B��/NpCG���a��p\��_c�k���[��n�F�;`�WMq;��vx/*�v	�g�;n�9�H�N�8w�v[�PZ�%.Ws�ڿ�C�eƐ�+r�+�Rλ���5t ���Q�)����4|OI�V�Dx\��$�t�G�A0%�A�eUMZ<�j����n�ء��ko�x0�v�1��w�k���ك�9��p�\1H�M�A�/V�Y�Ĕ}!�MdL=W<�Z)��[Qw�or3��xC�쮡%�����n�-o=j����\j�ԯO@�zm��I�z5�Ǩ�c�x�wbF�L`ا7v矖ydܻZ[�֋ý����#���jU�~yŤ|�,�n��*�aW�JD�q��9 �tD<��i�]W���̻��V'�we��3c���Bɻ�s���8�QQ5bk��x]�i�%�	��T�2r�T.���\b�]}�؁�H�r�;꼹�VEfz���~_2���A����aI�]Efj>��a�v>/���Ի�;�&����ʙ����D$�X�븽��{��w9�\�X޽��s'l+�x�Ֆn_v��V�є���ȉŔ�h7&i�<��e�O1k���/:��>�OQ�Sz��x��� b�~�m�Y2Iݣ�}k�+5A2<^7����h� �v���'�L��{	�g�^�N�xi�Oo��]�hV��e�r���\��]<A����	�A�h�]��i(���̮���u���ܫ���8�^�ha���Q�y�Aj��{Ֆ/��ۢ��y��I"\�	rH6��y�_�yV�*�{N�^O�v[�xD�e��j����YXBc:����}�D�3.�Ĥ������A�`+��撚5o��P�(]\��Vo\vǴN��>���V�]������2�$���	9�4�Z�_)�ͫӏ_;ko:a���V�>�d��6��V��K�1���L�m\���|ׄ�#��\�Gd�D(��<��֗m�q�
߃��7n�n�9��}ڡ�c�r�DF�V��p&�5c\�b�u�)���;NRU��\�g,9��F�p\�j�|Q����OFw��;w��Lt]n�y��w�ge���h��;��v�q�c�;^Ϝ�Ŵ/"Dw.46�!Uءt�B%x���!3�y�tM�G�Gծ�7�ն.Md�da�Œ�,�րYy�[�2])ͅA�䥛V]5��h������s'f���X���r�h�7:��΍j�Ŭh=g�͊{N��W*��	�*nk�N�dэWS1��g�\��-j��X����W\r��šs=�ѓ˦������g�5ngv���O���E�䍦����!r,٦v�u�f�e)f{�K�F�վ������\�ŹY���32<�s+M1����8�rӐ�;���H���Ւ3�l�~εz+�GEҼJ������yF�Jذ�_�w���m��fI#nI2��Q林hٜڴ.{�%EX���h�g[�̝ľ�C�*�����h�|E�Ԓ0EhI!ͧr�wX��»���e�j�K�㺢�)kC}��l�n���(�=�0kj�Ω���%�\IqI2I���Vkz⋸���| 0��Gsɨ�;���Cb����̂��N$��߱�A�PO�Nh㗮w-�]qɳ/3�6��w!lh�F�iX���b]��vc5YYZ"�tu������ʫou`��%k0a��ob�t��g8�4�+�������$ �����wl[~��h���%V�a>�%���Kޱ�d��h/,h����l����SB;W:��=��ݤ+����g��u��أ;\�V3�kv`���>v�5{\s��ZCZ��t�z����C�mduN9�8S1c���#9qF#�m��ݩ�[ȘA�����2���.�y^��7Nnw�cn�߼�ɻIn;g�V��2$�%�hc����+�!�պ�)�U	7�mض���(V8��S�����bj�����߳�	"�M�$RC��㝚�6���࣬Y��6�k�iX�\z�zn��Rl��Ϣ��m�	�������8��o� k	��E�%����v-�f㙆��M�[Sq���r��;���q�}
�R����$�U�|~��Ѻ=�}�cن��e��{��R_֦?���of�^�@�^�#�	�!�(3�C${��C��E���Cn����c��ه�z�;���QQ]��0mgJ-��4�˓��u��`�����8o([������ξ��^�L�"�x|g{��Si��O2��s5��-Q��b+Е��bQ��#G;�����r0�Cp��!�t7�X�l��XR��/]�VՏb���=6���/�q�����̩��8r8�v�r;A�o�mS�^dZvVI� �S�˂�zT�e��cMe�vY��oh�Ɂ���:$L��HA@����ԯj�
�y6�M�pd�W۽7Ļ7۷��>|���D'�r��*n�� Q�Y
[tَFzH�����^�K��%��bK���vQ�>MWb�!;�T:��.��0h�p�~���O[�n��h�Ŷ�l�I2�������2f��;���n�5�`�JO�'!��	�C�����opԽA�v�u��H���k���/i�;h����̘��T}�A�{s%��f�Ǆ�$m�#1�k��z�:�QW%2�f�1��$��7�/g�#l�0wk����u]�U{�U�r6юI#i�(k�@��$��H��V;�3k�V0E2��y�t��ͯ�l�s��SUf�Vj����"�Yk�hk�=7=����]�OF���gcŕD�����{�{����k1��GwZspj̴���@�Kk�IҎ��W����Sʣ���L�ORH�$m�������bz,���U����DoH2LetUE�/H�K�a�{���}�U��f�5K"4
�eO:�Lfv�і�cD�w�����N.��+���8��uU�r������S2E�n!�':�La�������Gi*�����5��C"˭�����^-{�}HO%�A��۲豺�/�@����lFb)��1��ӽU���%#��L�������,Y~���z�?W܄�0{���3�&4�T����.�Ă|�g9}z����F�c��%4B-4�t>�;)��D"}��g0�zxZcT{�<g������>�4�7�}u��Q@��(�5?|�^�GN�:�9���}ؒ�C$p��1�,Y�Fw��|kES,��>Li�.Ђ8��{�e���?il��~�b�l}��|l�m}��&>�8��\v$y��|wP���܎�"!&�f4J����<��s��Ղ;�m�� N��A+�R�\|���J���gH�H�C�q�y9�;���ڎ8QD�VP�[*N^	Gg���	G}ci��iLںj��(��'� =�Tv�նI���5!�h�׆W\ab�:�q*V��k�5�`����Gug.2�[N==%��z�@ܮ�u�kc=u˹N9�6��8l$]==qv��S�8�M{ԩ�Ư/
�ml[4�c��ʄqu�&G �m)�٢dK�������Q�X�}g��s�콌���0�6/=W&��s۶��e��+H�e��u[6�j�.�+�+�+�X��s�[oaڷ^uZ2���q�������i�x�o`���:�p�;+�:�"�6u��e�,k�z��=X�x��j���[7J��-���/s��<�_ ��嵐��0�T�1��'�iFj)
(]��4 ^'
��������t�_WC��~'��?���ֺF��Z�gw="1Y��/޻�*Vi|г|6����MJDvG�>}?cF�F�'p�������$�!�Y�3�e�"� ��4U�����&�P/�
a��CL�}Xx�>�i�f-��H�B��?���=~���
#����U�]!1��0�`x�BHmT8'������#���3y���;ea�v���<%�kN������RLѤI+�|�y���E���2�쏬����.�^0����G��tW�*�1��P��<y�{��F�Dd��#�������`�8e�yK~�4�ڕu�A�7>"m����i~�A�D3����%#���{h�:#b �_if�����������mc��O/:q�:�s;���&�[����;=�]����ݑ�r��Ғ�u�33��@�d��^��^#N�2D(Q{�V����*`3�\	lnz�f�Tt�V^u�ͤ+I4�0�?Y~�Z{Y����L�)n
zzl�N��Ç�2��c�ϯj|��s� ��E^�N�yj�;�3��%����`�b]�v���fv����xwZ�3��r�;C���:���{�j{�Ci���/B��yC�?Y�z���@�C<�Eu<CS�$�s��p���=>ύi�j��o-@��L��
Α>�P#L)Ȥi�\���9�id;Bw>:��M�jd��ޘat��k�&>�tt'���y���I�Dn�G�&}��#��"��=���d1�I�f9�5g�#��_�G��1'���ٖ0����r�O�(�w�[诲:�� �x��^*W#CH��x���"�Վ��@��G�;�Vu�����q:~��K�.�2����Ó���(a{�gv�rhve�(a��G������n�$aҍ��ze�TA[B4lq ~�?_��κh�k�,12k��N2.���cj>�`G�[M�u��ѹ���O�W\.��0�̑Ǿ$�Q�ϾKC�_��w.ZV�pɼ��ը3�����-]���� ���ʯh���g庪vRY�_���6��;q�=OH����(�~�4<{'+�s�O`��?A[�-?�Jұs
�O.������X:ElB�;�T0�唜Eɲ�}�H�)w�Z��#Q�\΢h�H�d�뼦����Y��iw��4G�t
������55"��S�,��T6bE,�s���q�D$��۝���T�Y^vt�*F��&���74]�R���M��L�g�V�"k�
�w[S�����D9D�#7��Dn/�q���g�D}a-E�L��I%"�#���¦��@�7���G�?o��͑���Ɵ�QP�̌~�Cbab|e�`� !�^��"��a����CHdݰ߲��#1Ț��r) �i;�d|g�Cy��VF75��d3�s�h�v����5��!H�o�1���6�\�:C�Bw�������oM�����u���|�D5��)�K��:^Cor�F�nԺ�z��� K�`�r��ܷSt-F\FDL�h����,��}��L��Pf�1o�Sp<l���u}��VߺϦK�Di$nz�Y��X~T���N_��R�diDBM4�9���!G�����4{2����ɡ�'�՞Oy�f�gl([d�{�,��#�k�5"�����)�DE�]S6]$��������8b�Ɏ6�r; ����y`"��׾��?!�3��ɉ�T��W^� f��K�}�wr��>>>"�.c�c�GO#C ��#,��p��Q$n����i�# iGUR���[��9B�U��G�,�{�u�P�?.����/�������:��J���]���;S�!��Q:�nc�Oz�Р�Uֿ�BV+��&�li���4ŉ� ���N턣Dн��FQؙ`���]���Y���O�x�Ύi�ƭ�tCbi��B��q<F��.�;�Ҩ�49A�0Xy��8���ʃCD^^D����4�V�{+S�"O��\b�ު�,a��g�G��x��(���W)��+�5x̂� 7,��Q�,&�]�7����q�ôX�,񨁌�HFb�����gP��|���YȌ��L"gD2"��b;=�����)rc�H�~,OYH:YC�j��{�l������d�\�_+<�yjb1@��ȐT�Kt�(�!���i�Vl*�����m�CŞ}�l��\���"������G��H�&���߶"���}>bp"1��=1������)��*$8)�߂V��X�3Pr�A�}vj��Iha�����_Ӂ��GL��bA��wi~��X�_S(cAҤ���*�t��'�dt�oɇ�� "IrX�7S� �wRH��*�E!z'G�u�<oV�?ML`	���0���/�fU^�0��F�@Z��xг�ɑ���A7|j�.ZG�Y��cal8ьc1�k�;�(�v���R�a�A���
�FQ'��}���!R�=0(�;�,��蒅�j����<� ���a�#�s<&���*�h�U��[��\Q�B�[6��ܮ�Dۭ�(I�k����,�fud�N��5b�����_q�n��*o�ս�wqN��_�n�:�4�0�nJɬ��'o�G�*kTVͰX���Y�T�I�T�����Z #3xH�'Ze�x"뱢�̵p4�G��R�/ ����Wa�*(Pgl�njoU؜]�ٛf��jgfI��~���Yw����I���5�ŀ����
Wpr�Ū; ���_P;�����I��d�61Kw��ј��\��kޖ�zf�����h�=L�)m	�X�/�H�<�J�;��w���pC�[��+7T��8�o��&k���-���Poep���@&�͂�0�����������3��Y[��R�������-tt�D��^�,YS�jەu�{���ֶ��M��`e�WG��)n�tf��s��l;��Rnӄ:e��i쭾�f��A��YBUV�F7TQф]}��ru���&�Y%��Ε�.�ngõz�,Ú�&��Mw�m�R˼��t�`��Fl�;�����]����L�Y)u���LZ.���
e��9���)�:F!Rˬ}Q1Z��]�1��ҏS�Tj�̇z���[�بY�{.^��9X|���=���^P���ǧ��<{螇�e�ϧ7�;�Od����
��o.��I��
��>�r�aE�	�M��vA"�;݈����N�������r�X�2_��oD��p�M��s�[�Gcq�c��W8����ra~�g���繵�]2����p�6�K�k�u�p2�ΫR�ڀn��x-ȁss:ӻW-�ذ����{6��f���3b5Ã�#M���\�׌�,X1)f3(�y�oVLa�k��:�6��tE�;K�R$�J��.ci;�mm\Iu�gǗp���)e�gM.$Q�V�F����y���e�1s�td��s�>+ir�힎�1�*\�B�A� bK.Z]tݶ����[2n$��Ŧ&��:�VZ|7Z�cn�[W���m����`���%U"1�������m�i��Y�G\l+��X���$��`Krqć0�[��@jԔ��J��l]{PuE���6�s׍����+7l�ۯg-�Ks��B��m��W:cs+q�'�[n	�Ä8J��|$�獚�3��lcUY�����c;14K�2���\t9Ǳ�\�ݱn͗Ѕ��a}������1o����x(�m��V��Z:�W!I�D�Y�\&7�^�`���!*����n����J��;U�4HI������W-�nz3�p�:�l�G)���g����W���="=��v�T������X�pZ&�]�3�c\��5�n:N5.�̓r����M�ۍ�p���vݶ���'n���td�42��7ml��}��Y�׃.��s��fn�����k���ղ%��뙲��F�]G&IF�;��,��hc�N���s��,85]s�:��䧃��q��3ps���b�e5Q��<��kb�)�U��&÷W�.{uV�s*clٲ:�,uvyr�DqVͧ�m�tmf`����U�:�84H�#�m�m�g��ų���9��^8�A��j�m��#e��@%�h2�Қ�hiw/��d��w1�p,n�Xe#��,h���F�>{����=l��5Ġ�C(SA&����e�ƤtͤÈGEr�D�@j�������W:$����V��m�:ΣяS������"�!b`�[���Տ=�ekf{Wnz��tzI��t��Q���Om]�y��q�셪���79c���E_�E��R�<]q��f�N�;<��x�ܤ��,��������5)�]1x��&f�62���G5�����z��Q<d��Gk��[�u�n���ˮN-�k������w���Ac���V�X�g����I��b�qs�8�.�k����iO`�=��{;=�v��I�i#�og��If�#���7"`vM#��� r�;�枦[ ��D��P�]�'&��֍��퐶6�RyRfh�W6b��k�u[�v����z����z$��`a�¢�;h�C(Go�?:^���\!޺4
�Q���6d�k�a�(�>"��cO�Z�%h/���".�SF c�R�=����a羛f���F� �Y�q0|yE��������g�`Ѡ`�Wz!�������������B��y0��{�Q<.�?!�)�T�rCcڄ.�/$W���o��!���K~R���ڦ��5�0���/�ƙۺXg�G��FH��n~cX�)�ɧ����k��:ݵ���9�P:�+��t4�A��52K�>�����DYz��F�<X:�u00�א�v��PC��qf��aE���|
Гa@�&I�`�](�6F$���ƃ���aۑ�C7� �tI��_����*���c����u	?a	��_�N��>/P�y,Ar�%�byu/��D6y������\w'6��p@7=�Zp:��n�V��n�ijs��j����G�q�"�|hiO�/�_,���z�����C,�s�)�� 2ځ����ow�`����)ك�Kb���t Y����m�SQڅ���ϐ�V�"�W�n��\$e���<"]x:���e���m����[t���wtP��Ԝ*�l)�����B���)xn�9I�B�utsv��H��r��M
��`���]��]��$� �K��ɯ,(����}|V�F��Ȑa�;�\�b0B�J"d�ًş�8E�KG��
Ѓ1hy�?��p��CHK�Ҥ*��D��P�X�G~��v�!�!�=�u/�o��\�{����-�f9��\,���\{�r�|/�L�Xi�T~�9pΠ�o���CLZ�Lq���V�^�&�æ�b�Qh���8뼥�����:GNbe򇁱���@�`�ӊ�ӟ,<��ӤAH���6:Y �k嘍	����:bP��]�!��2;]̛0eS�{���c�2eA�	���h�8|D�Fq��g��ӈO��9눒��;-��AIx���H�4��)�����i�\Î�+���tц�]�n~��Ekǌ�@�7��_��#�jfP��,,_Q�����9~LR�Q:V��2��l�2-K��tZ6~@J~dc���8�R ��6\��z����{)�!�T[>n��!x���c�46�-�s�����
9��2������d8~Dw{(�j�ba�_a�N��s�.��jK�{���K����vw�ÇN��Ho<�&4鍸$3�:$щ��X��ND���Ը@Q�����կs�<�e����m�J�}�����ƺ�^ԙyE�q���5CX��n���P�_vEy�I�� �~���O�:G�V!��l��*8+�h��;�P<���f�]n	?)}�CM�@�b��_Gz;���P:��\E�EM_��RW����5��v'��\��7 �>&"����92QϖT(����jB�64��H2�E}��E}����G(4sh
9E/��\׮!���Al���{k41gHg��.0�yC?�"!� �&��N�����<�ݮ�лUƙ��e�ݶ^�`� ����&N}�ܠP�F��+���80�r�����L�F�˞�KK�
!}���)�W�&,"��N�G��:�ag���@&���P"������77:��>fݐ����}�o�8�q������\�:`#1a~�+���Y����.���(�T�k�cOΐ�󕄍��'P��������#ƶ�k�N{{sG���E�����Lш�$NJ������p(���[�ƛہW0#BoU%����:�'���M��#"_���dIi���_fz0��Яs��B��I�$6:G�^Ǩt��.Z���y״���k��Y���V<Ɓ�˲�ϾUΑG�B�дh�#�C����J�S�m�ɕy���O"=y��g0���v���;��e� y�i�r�<],�]>CNE��{Y�%"<�����.p��F'�4��y�,�-W�n���M���c��~��b���O!�y	��ʓ�l�!�嗇�aK�"�/�2��)O0�(�\N8�lIe����Q۸ۓj�ҷ>�[�:.��z�]�RhdZ��bX2G$3l��g���S�e�^��~6~\AB�Ou1釡����Ԓ~�+����P��w�YP�pW��Y���GktΞmcP�'����E$Q���!r
�N��1g�5�Ŗ�}d��{3J��;W��׻e���(���gꞯ�����d��f|��"u�BK��}:��<�Xx{G��Q�0�q�80`�(Ҍi�	�?C�n�g�Q`�O��N6��bީ����$DN���hab�:Sh*.&D���������W���̍r̓����ʸ���]d��'�80���ztϨa��c	A��G����A��@�~C�|(\t|����&�r��!pE�Kdf��5a�sS���7po���X��m{���d��ጟw���<v���`ells��h��X��0�����YGg�"�q�ug������aZ	��B{�ъ��q��T�}���SqZzk*��E�a�R��ÝGt��Ն�w���[�Af�\��ٝJ��S�/� �Qp��T��Zѻs��;ynݼ��75+P�P[�s��tJV�;�2>k��/Y�N*�ZdwF��ロ�K��wg��s�{6�Cz����#�T�82�$��'�k�;k� ���p�)��t�N�t�mۦ�Z��|�z�]�5P�]&*�T�R���v�St���l�d��G����Z[/��!1��:9�v�y���q�����s�k�]w4�f��Q�Z�um��e�q������;\��k������]n��\����~?C��%��=�u��0A����5���?��dt�X�׽0�B�R����`H��|�M_Es�m���d�?��IVn"�� m��yy�<X����k��\�w��0v#l��^6wPι�,i��r��J;מ,h�T��+P��z^�S�:~�6��B����E��"���X2L���NB�w��G���!��������Q�1 �d""�=�^��hBN�g�P��
`�Ee��H����}P6&��}��\ޡ�:E�B��!
&$��AE7��1�diS�'c�Y�����}���mY�#�Y��J�A,|s���������j�B�J������o3�����W!5�G���%$�	PE 2A\��;ߠ���l����y��k�Y8 !���Q����&V�H�:��2~Sy��<}���N��7��Ԏ�y���y�T��!��C�E�;p���l�pd�>b٭6�tՌ<.7J��eMۛ��fn�]e�QR|M�P�yDE�w���/R4y����9�0�Fm�t�ǽ���g��,GN���#�ۈ<_@��/N�x��R�G�}-6�E��6�w�*<���rk,ˢqo�w	��ڊ�e�3�4%{ݰ�Z�:̌>��4B!���A��(@�b2����t�n�A̾��K藈����:=��ٻ�xi�v''�y�ǁ�(�'P�^@��0�n���?C�(iz�:�D��+�\<k��t���ג5#mȉ�Ӓ��di�,����\�K<{��!�u�B]��dТ<��z*��s�2���1(q~�K���� �q	j�Y��%��0Ѝ$$�G}#��=r��&��_4Y��k�B�h;C�nW�����$���t���������G�]/��V��#����c�F��,�\#�x�q��JO�&SC4E�L@�'��E
'V�'�,�H�H�����7�*��0�E�5am����"��t�_w��h�44����Ӽ��Dx癯�m�
He�39�l`'����kppnͬ���m��ݔt��]n���-������d3���4��z^6`�4��x�A���3��}���(���#~��I�o�u4D"{��U���Y��H������J%���~��W�zc��w���a��c��9֑B�4�����-}:�V�YE�ކ_L���:����l��é��s�0a��D������H�Đ��#�(�2&��B�QӍ	Р�2]{C�H��?�ܯ2�3SB��%�Կ���ޢMwd��t����D��J�{Հ��&�s4������V4��C�V�@�Ճh\Vn�<�]�Ц�4:��#�%ؠz��<Hi~�Th��I]��q�R�4��4�h��1���u���'���Y�X"&�ɉ�A������0�{3�Q�l�s��im`S��.ӑ����C6Eݗ�*a|p�bn2ӗϺ��!<}C2{��YFQ�R����M�s<��E���32�a����HY����ώ�ֹ��Xy�i�,#�} ȚP2��/6ݞ��ۅo$�gqvP;s���!���A<�����vj�0���6!Sa���?���-B��ע�:���I��	��bF, �͘��=�X�*���6���,�"�}s�����d��$�
ǁc�D
2b�C��="�H�L�H�����O�l�"��s��"���G�*��G�2~XẄO�:.�\�- �!�vH�7�� ���,�����i8n"��2!D�0��6F"�z��Q����=�c�ԱZ��Ys���t���c���1�ח�J��D�����x+珧�&A��"sg�.�����1�!�;�����������:`���ç��RI6��z�W٨It�|D
�4��kꙹH5�O�>��b������\볗/��KV:47o�!�q���Dj hg{�W��I]wqz�&���ۘ��m�"���0R�0�J��Whh�$(#fܕ�ޡዤx�<��Z]��*x��$���"@4�vr��ׁ����F�"� ���C:�gH$p��LߵP��/�XX7����F�/o��~{᣺�<�qq�v�.���������ԇj�Z-�v�W�kl2�N��j&���>"�c��ʬ髦2К��H=��/��9�v	����}y,G��'X��lsy=�<���{�������s��C���d�P�!r ��IdN� �#o޸i�^�6U;tiJ�?(�~S~�ī�������V�)Ti�CH�E���Z�<��V��ʯy�g}v��M�@����o�s��0�ncޖ0�B��fA��x����Č	��Q~�x��0Ԡ��,-�����,�{��H~����3~?�[�6�(�m�c�RVGM�uo7�Z<+�t�>ۚ/�0�!���
��v�ru��9a�n�I"Nya�e�u��\�%���p�;ccఏ���,C�4Ȍ$��2_�u&~�B��n6;��X�S�I� r���5�CC�odKȯ���	\�:D�W��D���C��HxU^�f���ю>�Ww�N�d��kW�]X�	�$y*��,C����U����{,��p�s�N�v��W/��.n��A�R���VuV���IV�8H`���+��J�N����c���z�x���;�T��q���6�&���"��MM�f�xCK�pM�v�vm͢6�R޺뇵8�lWu�z�'i��\jv}�.�{�&�b�Q�d���R�K��u\�����:�hv7����&���<��^�`�y��a���)c��ݺ����&�����4�i��N�Ѭi�{qZ��M`t��ٲ��8zmמ�Oo\�j۝�ι��sx-^/n	u�C���u^M�۪�V��{�w���,�6Xe��~΍�N����]z}(_{��/�����+�#AU^��,�4��َ�6~dA�I�|m@�r)!q�|ӆkQK�^��vAަD:�_B����ޛ�I��in �vx��c�7P�c=��ߠq-}T�a�Q��j��"O��?�Q��#�Xm���z@�z�H���EQ'n\�Di~���.��>�.�K�$i��*�r�kMj�P��.9��Q���1#bÅ���茂�$H/�"vh���&��(+�'ץ�#M��|���>����:d<D_���U��BD�	�0uk�������}��]+<n��H�L�e8Ӑ���FQ���\ӞTG��.�+2yk6
w�����?T7���D�a	8��Xbψ�0�4Y�w:?�~�K��ަ��ZmKf��n��*=�Q���u�zPl�m�j�
�F� Њ[�rm(鵹-�y�������m���0D��isWVߓ��(���:G���n�B��]��gl�;��t�,t���g�����Ш�$8bQ��Q��i�l�+�t�)�{�
��������0Dˤ���k�����{B�5��]��VӀ; Sr󨗡���JgF�f%�p���`��\�:u��G���Y�DH^��
��5��;�\V������"}O������|�#A���˭z=�(ᅊ?t��'�8�!��s:G`B���X�#$�&��v��fM�D�hr��[��E�����ؒ2!7p����EiB�b�jg����8�� nAc�bu��S���w��X$�u`bN�x�1��G��µ��$��S�AFw���f�4}�=�1\�S*̲��.�K�r̐�Qhs~�}�[���\݋���'���lxQ%���v�$t�6g��F��:�(W��$�Z׈������@�.P�z�= ��}�|�����j�>����{�(�mb�L�s,�`t1���a�';h�sǮS�k0uu��Ѹ���.ձ�������,�DY��ʹ��{��%��d�Ũ2C*B��B]�d��F����ø�?a��������O�:F��c$W���nQ�\���n�����a�T��}�6<k�F����#�g��ݕ��[�:Yf"�y��6�@�1�"{7��dh�4P� �!+�0<���"	�n9p���i˦߾�C���h�}�Q�e��8��K�2��ޟP���~z��5�KF]!�q\i7Q���ˆ��ݜ��J�|:��`q��§�R볋�u�X�2��W'+�ͤ��]�nV��X,am}�l������r�GYч��]�;�hA32K8��H�@ժ׋R���R�'�B�:.��:�UJuH_S*CR�$�V��)��fa���k��rg%��U�ҁ�aސ�S�4/32�k{rÍl�+6��kz��Eq��FZ�}�l�_6���!ۮGV�iyd`�Mӟq[n�D��b��a�CZ��6�!�]gh�.X��X\vu�v�A�6+���R�a뙯�mw6�y�k�GB�YM�y�L�n��iCw��Ze3C/j`WGػ�;]ǆ�F��}x���S�TIkL0vo���u$^�ջV�:㺋Nw:�����'Uh͡����S�{�&D��-pXޥl�S�YJ����L^J�өMͥwq Cº���r@+U���,��i�6"6^w.z���}��]d����m̭yM��F�ŚcX�:�����[F���i��(ӖD�Wn^���r��w����Y�E���5���B��Fb�Vw�v-�+;/mK�{JV�$`��;���@�UI�\,�J2�SU��qv�9�V�u���w0�Gv�<ŧY+(n�\�X&>�|��'O��k��EՎ����mJYzth��&%˫2�|q�m'��w2;k�\�)l��a�ޔ$����%�|�K$f�B�.�HS�����T��EM���wB�%+#�ާ�-g�y���v�(u$FDҏmr�|j��N��/8X��:�D��Jp�pX�zQ0�;�!Z�k�`d2s�\����d^/�����V�G��(�SxXX������`�"zFׯ6h�#�苝-4���>�ws�G$�ӆ��G���50t��=��C��Fr5�_ӻ���C_3�G���G�1v��3 �/�w-B��#�dK�΢q���pL�aY	NNE���RCr��d�c�,�lN8��Z�aNw�z-�����j����k5�c�vN��}��`rz�(��ڠ�73;�S_w�=�"���OƢ�b'�|�/oB0C?Y��}����(��mY��,羘P�nCc�3da���z��gI�ܠ�<hB%��~zl�(Wו(i�p�$w7��!#gڑ�V�s������]�&hWh2�J�	x>8I���q�"�G�Ӧ�7�,�1]|�aHe���W�;"��M�tYڃw��E�������99k�BAgO'���|���w	ᗣ�|c�~��VQ�@�L��:diVD~I'���Fi����|�����K!ZXc�&����m-_]����xlr$Q�4�7C�p�&��T?X�T�ĵ�m�1R�1��Ad8��56�]�$�p��N}t
;Z6�����T	��ll�����w��ߵV�G�����(�%/}pA��sN�y�1D3��(}�J���/W0��� VX�H�3�_�Ǹ�"�"��?d������2dG����4�q��H���:S�x2�P�����c���7K��ȣ��w�mP�le����v��6#�G�su��J���zR������/ଆydOg׮����DoS6x�{�CO(�?O�>��s�b�[H��H��Ew���,"�!��S0Da��"Q8*�����߄D��R�uL��A'�㱤?�}�������&���;�z�7ʈ�&�F7�혫Ї�o��o7 ��K5���Nz�/�mT	������x�O��Vx��F�{�*B̖~�B��$.���-#]H?}P��J^�(��
�X�D�#J+����UKx�l.�u2��/ n�
8�UΜ��ﯫO��7����(]:�wU>0D}+�*g�����	�(�܂��&��2d.؂�F�-��H��!�e���E��Ȓ��c�k17@��7 ��6�L"�u#{ס�:F5���F��)Ó��{�%�%d}D�,�Hk��b�ft�4�D5�y�Y���Y"�L��<{����h����gs�i@�+��ֶvb�B�������Fu�bs��@=]B�̢��,�^i������6/�FgFwU@��\Eb����1�`:-ag������k��-��WBQ��T��q��K�ls�/�
�@Ss�v��Tk����q"r�3����]]�'�=�!b-��Ҡ.���9h]Z�t�G^<o/6ђ�hT�s�Lm%p�XSV݂�`ێm�*p�ݗ����S�L5��V�����[�<�x�LV��f-�*[{+�.���Cx����j��7�ؔ��d��ٹa��v�J�ƹ�,CE��ZB���gv�Fd��f�Lȳ����h��1�3���+�z�����vQB���P��2&VF ؞��yll���P��=��.��$��3����.D�1��0)$��1Yg"E�\w�}Ǡ2�![�����#|Y>�x*�Ɗ:~�:���姍Z�'���d7y���$��(�7�{����C�k�
D#M�c����_<[�]{�a�p����b��l�����e�daA�R���Q$K���#{ے��/��(�*�Z��T�F�L�����>5����(ah�3.g��^���_N�tP�:C?`�"�+�UE���8Y&�bOy���-:M�!B�H�y�Ɲ���W��E�xU���P(�b8܆Ş��ȇ���Ͼ��4�:5����͑�S9�Ｏ�ղ�?�z�񯽱�5��Llq9���p�s�د�����S�����~����Ց����Ґ� h�
DK�v��C�9l��Xv��&�:��=��䓭���Dl�AQH�p6��%qYj��u����uqT��B��$?f�'B�-H:~�C{�e��	�cb��1��|��uT�����t�"B�>��cňم��m��aӆ��)�(��VX�W� TF�>|C�mR��^!9z2���Q�܄��f��5n�u#�����[ь>ǎe�ғq,АL��I"2��n��I������Br;�{��x�><|DR�A�w��ꂰ�jQ�޹���7�9����h����4~�$6��L@��P�q���:֑Ӻ�����N|E|��\|ƛm���&Xz�El� @W�&�c(�3Auf�ˈ�$w l.}��R:yu�iK��߂Q9�\�)>>�L#�X�9��ݚ��{�ք��yP��Z���ӳS��`qF�(�'�ŉ���p��}v@�A�;�{����i{�)���f�A�Q3�)�d�I(ih�6E�.�۾��,��Y���L�/Cq`��
�Y���Q��z�`�^�p8��N~q���?!HY�(��+�'F�T�_<��9��xW�x��{R��M�x{E�<B�W3�Y,�X�g�is���O,[/]\W5w����w��0`Yf%8=�,Q�*�41}d{��^��$�Q"�I͑y��
Z�1u��}���a_"O���X�
��4�G� �m}	�#��n
ç���dT���W�|બ�nIN*#C2���@����Lw�c_W�b��Z�0OH��C�Bb�8>�44�\�9�;HY������*	#J9Nb��;�4��Ͼ��4��r��_S�n������^8Ta������b�`�Dj&����'.����쏆��v���2 ���S��wN�(r=���@1Ѐ��X���j�����!��Z���CS��">J�n�^��nV�"��_��]EI��Q"��RCCM����:|A�c����ee�]�8�D�?L�_��fLb���'���C��iGy��Jy'�}���K폟ք�@��>�sI_G JH��8󕨓K��@�*r=V�1�F��1IQ��\-ӯC�<��!x�-����֚ńADR${�0?yi�&a\��L+<~��ݺ�C��F21H,H�o��u�:�9۳��NR��7d2M=j��bye��f�Ζ����<�����߽�k�"ۈ3��?K�a,��1�e?C�d�/�$A��t�����ޯc8d1������P8!n2�u�iύ$�Dv�����cK�j��qC�4�����"��gA_�~�,�8���e��8z�nuj\���+�6��{4�="r(�i��I%�!��#��
C����;ıq�0}�x�XE%�B(�X~�9�3�{���dI�n�ب�ǯ�(a�� t�:�������0�E��FH/�(���9}4�U��jD�џo��'��6 wϙ�oث���(�zE�5��r����Hi	��w<���.�h��M�W/Li�˖��Z<4rn-�=��֡�F�X��LQ�r��N���u�XmHx�����r
�jv��� �A�a���t�7q ���CM�0����y�1D���Y��^+��]�͎������͞?T|����&��F�z���te�ǤQ���"��u�M��͝��2��b�mGk�9�^۲4���t��
�X���q<@�����}�����q��&8�y�RD�A�a�~2��j�:��jp�a��'��Dh$�-"=��B��m���];�(�ɿnt�6�i:]O˯�%S0Q51�ӆ��@�Ӧi�a|>�p����e���Y?-\Y�q���ā��4�����o�?��7�(a5���r�ڸ`�WK�Y�&������>E�h�#D�nE��=]�͔�r���\�vt�B�9.>� ��_��� Q��E��v�~Q{����GHG"T,�j��{C�4�4���E���
�""ZE$�m�C���Hak
��ŷ�GB/۾U�����(M/��W,`?N!��(t�y<9�Ha���vti�{~u�-���B0Ќ^!�`@�{ARA��B�E#�t�a��:�a:�z�44�ErQ}W�@��U��XP�����k�}��f�dd�9�F����}��#C_kS\�����˽
�yX��3.���݃�� �H�U��uTY�V�.��P���v,r�at�7�sm qd����ʺ��gb@vR����u��ymԈ;Z�j0�a�s32bect�3sw��.�ViWj�pm��\C{�rz�:^������5��ZAe�%���&M�+Rz�<�䞛�q�[��Ӄm��9��{<�1X�9���e��.��
G?�z�J�9���Uж�!�b�]�p�;4�Y4Z����:t,T\�h��u�㳮�]�+E6��dfa�1xƫ��WWGf�[{+�=�TZ�V^��K��p�al�v�t���P���,�Z�Y5�g�㵭6lyx��_���:wߴ?��8/~�#�Mtf�!��4PS�dRO�Z|I�A���U��MOљ�託�ޔ8� ���G�M�8~(\!�L�ܰ��
EL�
R	$���g��Q�ڌ��4�Ud#4�G����R��P�=�����*��c-|��F �Q��Ȭ#H�R-|�>E�C���k��#k��e�N���H�2��A���EYp������	��'�C����/�L	L����Y�T�b���6`�!�D�%�P���Njԑ'ڙ���!_'��{[��B���>v���:'�캡P�x� ����c֧�.�(�NN{wS���C
����0���R0��>* ����X��U�t>=!e�Ο(5r�l��S�Em��pP�>8Gz��m �����i}:�U��^N����E��'�s�ȘBy�P�+�g�:�Z���CO&5�f�o��g=�?�"�jw��&`�^��R[��1Q�m�7��T�-͛���(�A��j��"��g��,��p	K���9k�Q�(��;v��WRO:.}Z(<�z��֯kBAFH�fNu{C���JHԤݮo�|�q�0�Kv�O~S��>;�E��S�8��ux�
�~��H֭��,~c������W2�Jf7Y�63�`��L�6}�
Ru�r���Σ�>�tq�K�2�VTm�y�F4(�>��a�JX~������t���I=U��X'|c��1t�s��:�d&Hԓ1_i��t�D&��G DYCھ�@ϟ�?��e�h����p2"�r��8E����U|�Z�i{���@o�9�A�ۡ��"�nN3�J�Վ>2��+�r��Qg��0�7/���,����$�8�ǽܷ`�6&�����f�������o�Uu�!���hϷ>&'2����`G�M�dt�"��?��,Ʊ�ۣ;i�]*dn�󬟞ǀ�4�`��1!}k�<1d��>�Eo���A�PA�u1���eo�����>�����T�y�kvm�Z���t`�*f��lt����j��:g\��IU,i��D��6��z��"�_o�2��������!+,���{��w��o�f�X���t�!b0M�1kb�k�-V��m(�&(�RE|�- ��0��P��pŜ���V��+&>e������C#�i�Dy@�D�b�"A�C$�+z�..�i�3�7�^�􎞃�CR�P��j#���"��d#�6�a��c�j��;��
?@�{�}g¼�.u�х�ٽ���l��msm��ӫ:���]�=�0�Cu��F,3;�u'� ڬ=|Zǉ0�]+to[Sߠ����c���SCH���+�rԫ#A��YoO�|0ωDc	C
�&ۑ_H�[o��- �>C]�h_����8�!DYm*�}����Xh�f�	Ŝ�~�>_QGWd3�
#!+D���4�u��4��Ǘ��ĳ����+�E\m�"C~�7V����p���l�&~�<ƛ����ޞ��������y<Ty�e��}�����I�Ծ�n�k���gOӤ1Q�'�mUΟ5�N2a���6#�V�����mŔ�g=G�fR���v��������D��v�߉���O�B��Ls�0��>�����1GuA"�2֛0e�>���=����,�����8da�;�=���ya�amdiDb!$NJC�˲4Ч�3�����#���T�w���	}7�8ա�~��Ȏ���<xR	{�z��.6Q4e����˟�7;�D8aG�ϗ�4!��81��
T�PJ�T��s���4��@�j3��(i�%��QP�vz�Q5Fdv\�#��׌�0���?I�{`_���އ�iӇ�5���&�f���R0�I�CDav!/��K�T^�	g���Ipj`+ެg��όj��	�W�U�L2�.&���1^~�T��܊�5l�;N�����2�B�Uˤ7�Yﱩ)��1�����fuuX轔O-�'U��\��&r���7	o㞓�Н������M���c$�9ӆ$��8C�����������y!�&E�q��_���Ǎ�Dh�A���t%��J��3DoK�u8ޥ�z�|�R���,�8����|���],vф��	m^\�YQ�5u�T3tU�v�v���A�j�=%;Xڏ��+�'��J"�����P,��3$F���d�2!aD�� wo�1Y�IR�S��G�QhE���se#�H`R�����~%2W�B���1_iK��(��炆 `�;0�Y
�>��my?�Dl-!�G��thz���LI��4d�h�ϒ:QwUY��+�WM�̒�鯼��ME� �6\����6��ԅ�������N�t���']1�l�ZXx�F��wC�+i�f��:G�2���i������b�ׂ����!)#T�"v���.r ą�di�|���� � ����?��?N�@�p��#����r:�$�p�=���Q��A�A�}=tIK�z�g�䏈���*ATQ�����k��wi���y���>7l$)�׽D�9�$�ce�&l��):X���Tm���)<~�C�+���kO>Buq�w��b����W#H`� ��@�ix�T�{�����P��{f05���[�M��o��t]2����*kp�C!aK����ؓ8o.vav���Y}�4�<�mP\Xp� m����c:LRvk)V����KJ�����F!7�*=��+9�w�Dn2`.v	}��֭$���8��7/�չs�I�Mr(�=��c\̝{-;�,S�n�U�̽�yT-��I'A��L"u�
�3��8�eĭ�>��4�Ub�B(�7�gy���Y���ءv�Q[�����1�;[�R��UhC$r�w����d��;��Y�(��Ոn�[Ĩ�0od%l�.���r�s�=,� ������v8Z��(+�6�y��A��Ŋ�&4u'�
��:�zqF��,��c7��-}c����4ޝ��e�5�4�ެ��n�OV܌�U}����}ˢv��jo�V`C��+ze(���in�����E�!�iX�[�G#75mKCyh���k����m
޶Cx̛���p
�M4�ɜ��*�&�O�
8l���3v6�YǼh����䡑(/;o���7�Cn餷V+���>5�	�N:�|�}�t˸�oeA�._��P�zb�ݲ�������N���{3N��m�ǎM�5�E;�RVO�yb�*G�G�+���r%K�TR�X���N��$�A,\� I[��֞����;��ZTe�s.`���8�_X�,�"r�����>�{|�A��#��|wwn�7��:�_M�]/+xwVsrU��SǛ�w+v3`�����o��z�;���3f
��6K����8�3G��t�����+�����n��vTjm���Cur�3gq���T�3sf���}tL��5�Kb�ufo<<������¢ht1�)g��Jj��nݗ��aт`�k�$�P�%ۙ�c�t�ݏ6CC'!�ێ}]�\�qִ��y�K��Μ��T���v]��8,E-�u�6y�TzL�x��n��@��p��w}�h :e�e�:X�cn4	aVb��
d��!�CҏK���&lP��R��`Z:k!"�E��q���h ��lIf�]���d{\+�SZ���76r�68ͬ�,���������bݼD���8Jh�0WF�W^�:Ffy嫭b.q�uk�z��m�<��&��kS.��m�\��ۇ^�Z��E�hs����v��6L�kvϳ �o#{���1\���
:,�KZ&fF�im�LN��n��x���ó��b����qçt]"n�Y��(��=�A�ON�nm�u`�ebmw(Ѭt���c��ɖ��2�b�66����x�9(�<�=�S'��C1d}��%3��x:g��;�o.&�[�x������z|��S��6m�0b��6�Lvz�g�N{��nf�٣��e��`��\W�kn���Imk�\>��]�Q��Ͳ���=uɞͮt75v�Y�ݗ�k<����q��i�1;�tj6�틭ƍ��M���2V���zU;Px���A9+6���z]��z�D7^�=�
bvM������!2������w����z��n���C���0����M�s@��H�R<�6�������Kn����-g��F;BNz�]�sU�rF�.f�%j���*lq�ܶ:<R��`�G`%�H�����\d9�XM�g��u�X�g�:��ͽ�����{����p{V�-�7�����k�����C۞�O�Z∢�TwH�����9�^��s�p��"fTB϶�]�6���F��0=�]=��9��6�#	����m���6������m�n���PI�G:5[�s�Ͷ�03��n�g�"Q��;���t"��kD�m١ť.7�ݞ1;0�����bu�E�i@�!���. �y-�R^�6�	���.j����bZ���c������d7J0�]��v����j�<(e�:&,nas��7�w>$�<m*��ox�CU����б���]�K3LyN���:.�]�s����=Uq�h*�zQM1��h��V{n��^�8�,iy���r�;�J���^�ٳ:i]�i��5�]��z};�?�O��,��(i�d,CM���j�_���Ņ�ϲ�g��..b�(�3���V�4�(�-IR���_�C!��Ԏ)����}t��fc�_��:}��9k}�"P�$N_Z�e|�E����O���f~Hl�[C��Xl"ͼf��G�>��H�ΡR��Q����Q$j)"���xh�?�Dj�쩶I�f�$�Dh�͎̟C�/#C��	{�'�=��ނ ��L��}?[�����ue��@]�xХ��]�1"-BL���0#-YhP�}��`d+����Z�ʝa�ENϾ�B����R��.Bǽ�j���5\AeyϘK��?V�;��i�~<�C�@Ѵ���h:Mq6��0���.-D(�\�:�aY�"r>�o����:��V��_`���$B�(�z�j��폦��F�P*�
�{�����rP����PZ�W�g�A�`�����ƣ�M/k&�Qc6Љ�v\�J�$��}Yq7�[fi�m�2�:�~�?��|'����>>�5���"L6��tA�M԰�E�h��b��܎��Cߦ��.��`��>$5$Q��_����i�Q�E����u��@���7Ο�Gx�l�|��m1Z�ѻ��!����%~�R�Q9wh�Ziִz�Hf��%|�gZ}�<h��1����z4i�'`u�J��kYj��Y�7v�)�0��uT�|b�wj���hbʾ�6Q�&	k�O�z�Р�!!#��e�0������Ώ]�Q��4X8~B�x���AJ!�'%:
��:���6F����_n�6D�O��
�_Q�`�3���� �J��/��4�)Q��,am��N!>VF�({ؔ@�1%RG�<dVh�o~K0����"A�}^i5�e�
'=~�/�� 2�|t�0%
����ݏ���9@�fd{�u���@Xx���8h���0!K��p�]�~'\<'��XY��/�;��ѪM�⅃P:��)��_����q���ݢ$mfhzM�a�u*t��K��U��3���6G���o���p���h [�0�e���F �\�
;r���v��&+3�k�8�v 7>[�t2���c���ts���������MkP�f~1n�ʾ������"Lӂz�T�P��P��o>�@�:�P����40���8�,0D}b�/)������JCVt��WHuQg����tEv�4"Eo���qDN��JF�
��ȌH���$��X���HԤ#P�__�[,i�$f�lW�	0�%�x,|��3%)"�g:wh��$G`L�A����,i|�Z��9)��4(�!FM�6�q�<�_�Ey�p)&����p�`Y:�s!"J�w4��F��+5����efB%�t��Z�es��sq���:�"�6�
��
A�����E���Pغh�������䉏:lyf.O���*I"7i� �V�ֶ����(u情����_qF��_ԁ�S�,$r���"�뼘ѫ�?	�GH���FPþo���3q���_@����"�?��i��t�5���|xtsߴ�bO�F2�b�L��[w��|ڍW�:�Wרe��qf�G�a��$#���\�֝ζ��(b�,ɌAu_�i�u���R�6�n��͙m�z0mo/RB�s3�)�t�f���;��Fx�t��I8cF$��z�eQ"HW����:t�拝�Z�G���,L�i�5M�&	�yߍ�dz��˟�m.&#A�3+����ZR3HZBy|p)
FZ�9��ִ|C�6\*�^є�g��ȷ��A�����|g���S�Lr�z	F����칠��0�H�"��U�5~�<:N�q�A�Oƥ�����9����rF�
8ʒE#�f�|�J�D��^�Bt��x�ä3n�(�
���T}q2��G�󥛢,̉0$9��Uϒ�,�0t�nX"_/ho}�4�+#���z��I�a�(�,�K�cg��̶�?NêI`�3��ʚ�~��B�6>�Oo{e��i"�Aq
���y��z.���T��d��պ�j�?Y��<G����1|�W�:wMdTf%�h:�D�;�)V��֝&���ЫvC�'.��&&c�B��̒2-E�)դ�t_^��$ 4�#>:�cD6\`�I"Xn�(�"�>��Fs�y�\|�q�|B�_�Wa�<�$5t��l��=�c@s����`��4._�w(�<bcJ��B��X�o<п�EN!x�m� ��6�&r�ƍ���ѷ)��7��8q`H-8�%8��e�&��q������.~z��"q4T�w�<k��0RcR&��A�e�2)�e})iJ�ʓ��H�A�Ⱥ�Pj���D"uI?<�Z�Hڵd��EP����3-�HGi]�>5DjP�{0m�$t��+��] ���.U���R��0�����K��@�R:#�ya�����7��>���1M"� �[�<<<�!a�Mp]�����{y��q���{t�z��M�b���=Y�Q7�&�H�OD_`d�9�d"�1K�*͍L��	e�����zGN�9o��'�s~g�m�S8fŻu=%O�^�V�<���{9������曆:���u	iO6
��EY|��6�����P$o^���p�`YCN���#=���[�y��0�!��C`�x|���R�)#R�N���@��L�� ���U�8-F7�aj4v_t7��`��qW�'c��#��?J^��2��ԉ�������V��#1B:p*�J$��"��מ��N���ꨁo��؋_���]�VB�j�Z�Çm
�������t�Ȃ�4*�Խ�X�pi�-��I��w�w���,K4mgق���� �^qb��w\ի�L�µ�Ԁ�a`^D�N�n��:�v&9�!�.�Җ5��,L�I���qũ�"�jY����hø�[M����4c��r�����F	�)b ���bM�N�N_#��X���Dz�[�HzݮU�k��n���f�0�ܷ.�5�N�����=��P��q�ݤ�[j*�l�s�3b��2���ۄ�6�m�����ng:��θA�s�t��7e�F�^ޛ�ۅG��H�Y2�m	�>���g<t��t���6-q[f�{�@-#���?\�Z����?f��!'$I�F�"h.I��C�H�&zC8a�3���1���s����K�}�l;"w��d�N���\G��VaF�s*�:���K� ��NDi�$�|�^���F���/���u�v��6E��Y�Y��9�Vht>�N��HKF7�$�80��*#K�d(�gs�Ac	��0��Y����H���0zz�T���f��n�;�ϕY��H����2s�%!�G�"�Hi+h�e}
�J�BHS�9&s��!��3�J=�ʥ�`� ���tNl0EL	[(�,���<"ח�"ȃ�Y�7 �fa���4�!aҍF���ꬊr���`�8�|Qz�	'�3f���1��ےQ&bBJd̋x흌�Oi/oV���4d�"��V�(�Db����Sb:�:p�4�W4�w����$F�-�b駌#�4S��0�4���٬Ws�y}���oSnD�P��e���䢲�ͽjv�`�T����;�n˯]Xh:ζ�.%[2�����|2z�^���u��`/{p�w�"�a��N���x4F_�T�(kЄHDO�`�7�����u^��m@�L���.�#u�1�"��}�i9@Ll�����ۖP'|DZ���7��5of� ��g9�~C�]Ѯ�ቜ�|[M����s	o:�x��*�mY���c�ދ�:�X�[[�z5��_f^B3M���>H�!y*�W5��Hd��	}w��L_&��	iF�L0<��W��Pw�H:�,2!]n��&J}�e+V9]�߃n��5
PG �t��\�c�+TU�8�}��5��Di����g��>��At�!gهǋhH�멠�����g�H���u��tF��w�~��Aid��흒2�AI�5�`�2��z�ey�@L��j���(����#�~4~\���a�쏙��i��}��U���4��UUA4U�C�+�������L�4����������m8�1jC|��)��v��	k=�T�}RC!��3s�mҊ�Kq>�$JE��""Ԥ/�X��������=�O� ���Z� �F|4��Wf����ډ���-!k0�BkEŭ&�f�����v�ːTӮypI���.a�z
�33'E��S#�D 7��(i�%�F�7�!�����C���g,��H�6C�{�Ü�U� �ؤ!�LR��ܹH�H�%�� ��m�	�pB�A�%=+��;��q��~��V��*C3v;Y��7���K�D4�O�^�,�"��DR�@��Y��d�R��Pf��ɫ����ܦ;楶t��y��+�"�1/��\q�q�YpP�B��I��&^�g���R�����AsW!��s!�v�y���\�j�^�N�7S�Bh�ǡ�%��+�_u������P�X/1��w/>�i��9����ŢZꗉAB�7�����n�;Y/�"M��C&�E�7E��R��0Ͼ?�	i'8�p�"�t�p���\��+���1ޓ���.�����0}���c`E$dB�(��C���P�R�yq��up�|t����'�ݦ��@�)@��C���'��"��9/	�TF�E�9w�o���Xx��i���|�Zv���,�������{/ɊH��OJA���t���A�L�Y$>�"��꾰�d6�p�(#RnQL��9��T�х����*��ӷ=�����6k��S&�]���=t$>�Ф	�����"�1|� ��x����&�b�fCA׽�4.5���c�\}�K�1y�z^hC�������<lK6��8�4��cH��e6B��+t���&�w����DڀO$D����Jr~DF-0n����c	"Nj`�_O���Z�0I�A�ӯ�,��K�W}�⤂.F\e��,��;<��1��z����,�"�;X��P�������M$i����x��0��t�g"�P9�~��͒p�������6\����B����n�2BTe��"��oٌ�"i�;��U��${z(Y��$��!/�X���M�#������>7g�L�!��W'�&zekxY��Տ��--�Π��C�2�T����t[g�A��@2ջf'c��ƃw7۵��Vh��*����]!KN�6�0m	��6��)#m��%�z�6D'�<Ce��1�cL�:~���d�}t����t��~U�:ь�K�a���To��LQcM�,���Eh8OR&�,0zWVI�|�>}>��,B�R0�n���,�v�%ջn�M��ښfa+��\����bV�Zh]-K�	v��}��=Rt�}5�7@��>�?J���*#=Z�,���
F/�@Ro��,U�/.���o�(�����0<��� �}�n�[=\��H`5X��Vb����A�&�q_:wU�>��	č�}0С�� ��b�H�'P��Đ����Z|�A�ǈ�5l{�v��
dB0}՞.�4�~�c��h�Ξ��V:cr"[����9%� 6F��e�:��S�����Ɉy�v`b��I��Zh�;�r~�!�~Wd�K�1�R,o��m��C�OcH��3��~�Ϡ�!���(��/I'�?wHf7!q�>��B��l]9�"Βc#�{�����BC���Q�o���j�M�$jJC��Zt��U�u�!}�h�4ZD@�P0a-�ԍ��6:t�#� �������*N�����l�<��d��y������:>r�����EI'}~�@��q
2@�H��P	1�=���f>ˀ���D'���� ʹ9���mֈʂ-�����Q��̵;�a�ﰟo��\��wڱ3�_w�2��b덳� ��i��}8����.����>���:�KrJ�����+pl<B�o]��0�:���cC�<��	=rn�-ˣ���f��-�����@ �f
�,�R)o��v�xm�\���N����)͊6֣�^1��R�VyݣvR��7k�h�[�؏��� K����smZ�%��ų�#a�it�xՎW��s���`�;���ùy��b쏦���f����ڸmUsRv2���Y�����!B&�`�T;� ���r�<4u���ӈ��1Ƥ?��������Bq�]���v	�f��cS$3q���\��p�$"�+�r�>͚"��V�4��+D�[�.��4�&��3�2~^�lFND!2C��à���#��B�>�����V��Af�$��a���?I�g�M��oŊ��!Dづ�g�����|V��`"ElY��q|�B:��x��< �6�rN�;��ԉ'�]׎�4?f훲z�����3g0�����&��h�	�K=�_Y�E��:����;ȼ��$��XY>��Eg�i�R�4�'�T	�ixi
bJ	ㅠ��=(��[@�ɕ�;���ٴ�,���OVCh�	� ~�st+�f�"������H��i����E�Yk���}�
8d�{��ؔn�����=����y�
�����dڵq&�	������`q/bg�ԙ�8�8�ٰ,����6g�Lx^�,!b	"��y�ײ4�E���0�H`�vs�:�+5E���u)%\�:�t���KÇ���O��g�фո�;WFv̀N�YkG���0'}��4daD�+`"Z���Ɂ�y\b�@�iւ���b���VJ�!�2$�FY�"���o�~8_'yY�xFw��~�]��c�Ȝ���Ӽ�a�I�r!_�&C�.��,�a�6~R3}%���=L��r�����i���c��:�v;�"fJ�Ң��B�lZ�JGVo �nrJt7�����0�#1��m�K�ڿ~�V��2��x������c��LsLI&����GGԡl������l�Б�g��#���4�5�0��+z�&�&�QHlf�TR�i��!;��Dm�}2e"A����"���Q�\tB3O.��Y�c(�<%�<,���vM��2�H�X_�2$���إ�"��W_,F����P��9��:WM�7�~�(ƴ��� }�R�P,��5�,�.���|�0��"�l�H�ٸ�>a�d(��n"�}?Qف�G�����q�#��(�F���y}/��]Kn�����CL��M�_ϯ�)t�E x�b\�T}�7Fe��^�<�+� h���$I�Vx�`��l�D�(��ϫ2]��=�;�t�N�����k�+����)#�ն^3 ]�H��9�K��
�3�J��έ筋�&��.�<�K�0�g����~����[��G}b"Є���;K�EqM�Xz�ƨ���&�S�.drD������ѯ<��P!�}�c1�Y��zP�]�x�Z�( �W����i����Fۡ�kt�w����L�Zl���6Qj>�����t4�dt|�#;�"¶4�;��.�
�˥I���=����'<Be���^(�!w?}��� ��O�]~s�!Pf�(�-�	��~��	,� ���p��ӶBG�|�,���}�,��j!L�#����c*k״*�=�E!��nh�t_�)��A}��a5oSPe:p>9���μ������{OK{yY���W9_fg(�p��`�.��f�*m��u�^S��*�E�$rSiH�=:�������C�c�k#D��s����a���&�o�N��Tw7��o Ya%�GwQµ�*��!+q�A��w���U������� ����J�bY\xn��X�w�8���V�O���XԔL��y �}�-�F��_JW�pvU��ŚN���K�n�������G׺FQĩF���G��V�]\ʼ1��,�����NľQ��,^��
�z�E�.i4�LSOgVXٕ�X�q�f�gY�;3m��թ�Ft�U�z{Wp���k\�v��-)[\GZ�KS.�ֻ�qV�Y��4M�5�y.���uÒ����k5���Y@k]e�7re[�/O�W���w(Р��>�JNc��v��if�:��>ZNE�}���_N���r�]m�V���3��T��|8lc�'H��/o0ŃD�K�`����h�c]��WL�[�k�5a�h�[��a/��Iŷ�S�+p-֊j��Mnf$�ސ�Gw��.6I=�x�[Ojp�P��[v�c
�d�j*5�:����_^�f�@��
I�k�h��g��=&ho_C�u������6��w˴"L����HCX�v(UҔ�xdQm;+^ےU��eIf�-�szt�C��gk��#��f���Dc�C+"r��R���QI�A�eq[a����ȭ� y�f�{	l���WVv̼O.']���^����i�5�H�S>����
�T�U������D��1�H�=����FO�iD0��K���jDp�)$�'P���H2b�K�M�o٧����o��Jպ������9|A}��Wd΢� Ҝ/F��@��<X����_iw�����6�����0�CL1+(��|�I
�B�-@���.�;8�s�6�{C5|ȋ����t9���Z��jNt�$�ށ"�/⼅����V��
�~�(�Y�헀� 4�̒B�xB2	�ןz{n�5�Aq)��f�@��7,\�Z���nL���]�
l�V��[:�������rda��HG����B�ӆ)}��Y|`��̇@�؂M���妫����Ƕ-�'�z��k�ĉҥ!_�I/������L�̀4BLE��v}��nk���{Ϗ���O�����_��5d�==��oG�;��P����������Z�8Q`"�)�zwl�HCHB�,�#|�ʅ��<���Q�w�D���NL���&�R1	�����G9��!
���W ���,Q#J�*-}L)D��D��g�P,l}Fl���9���@���xw�]#L�i��/��/��M��H6!B�T0�����ϞP�n� t���6D������^^�;V	ԯ�*��(Y�~^�f�4��&�0"����V�F��km�b������F����V]�Q9�[�X@t]��d�}E�ze-�y,��e�� ϫ�Vbr�DV�$�n�>̵�Ď��ρ�D�s��L�@���H]e�u�q����x_�����D��x���#I|D}�$�&�P���t����r쭚j�ږ�����O}�t���2�B�M���n֑��Bq�#�j�9	�|����G"a\Ivvn��-�xq��t�����u���5�+��c[�u^1��-��}�C�I�u�H}@1�!�}��^������{!�<���:#��<BWHv�'�>v|��E��E\�ۡId#Iמ.�C~n$�,TYh�)F�~�\(�ے잡,��T\A�u�}/�9��G�5�t�s�N�6\_M5`���S�~<�(>(����^qv�6h�(���x^{�u\:F��Ľ��lβ|�}>s�"	Q�x{�ʙ��$�� �,{h4�4>J�/'D�Vd�؂,��w����%�c௾x�^�� �4�9�gnU�12M��:Q"��xK����'�)6z��gJ}~�Ƶ�����i�p�F�NR$�S��-wt�t��/v|�� �%�&�aJd�{��X�i@�9iA9� ��}��x�jC���` �$�������O�7M0(�64��i@�>�x>�Hx�Q��-�pa=[�p�I���Q@���_�ܕcL�D��!Č��{�e��/~���� H�(�6��ȃ���b@էU1:��5���}W��P���t�vW^�Ƒ��m�U����7Vl�q��X��<�����	�48��z��\��XÙDn��Jj�ږ#X.�b5nN��0�2L���դ������`�ϗٞ��!Yq�<�hY�V�ػ4�fΈC��O�ts��g:{!s�8�U�=�:;c9�+�Z<�S�h�=�x�*�7v6����l��,7�[�ۣ��8��8�({m���+���XL�E"�'^�ef������O#x��R�����3��ǻ�i��ط���]��=n��7\�VM϶�m>ggV��\,��ϯK\n��`�������ێq�ٞ{e�&�d۞�-�:���n?����N�ʚ&�����єI:�z$��}�<�i�8��b�^k�T((K똉=�.�À�h�L>"�$�NrN���ϯe�∖�b�r;H�}�sA������j���5,a�l� >� ��`^���o��5��B�PSL8g�"�{���:���ې���� W���U�D�"��.*�>�^��i�BQ�"�p���:#�z17�1�>�[��M�sp8j��1�H�H�,�	h>	:���qjXQ%�����E}�T��(0l�53���*��t8&_����Z�
�"	�=9�?SuZ��KR$�힒�n�
w���Ƹ%��]�U�Jϸ���	<�Z�ڪ��xu"{�"v��~���7�,!<�� �0A�=���Y�$Z�͖�&<�x��F��jG��D��罣����������t��tȄi"����W��k]6�y>'��_�>���L��M�w�G������捕��zs��X�p����TX�M���5}��#�imt��į���^�+�. �	Ĭ��]w>�_w�o��?P큎�Mu������;���nJ똮�ɜp��[��v��H�N4��A�t��xD'�(�D��XӘ	��H�9��Cr�~ύ�$�y�	� }\M�M�H߯�a�+p@gtw��,��#PC��A#/�l�gR������N�!����¦�Ku��:����'�H��&>Cݗ�t	 �O��߻�<7�F\Kq�"��u���UM�z��%}�Z�wX#ba���p5!����x��+D�J�rTκ�'%����ތ��?Wք�D���ٽ>D# >u.E�9״P�#e�1$D��I I��C�.�Z�����z���dPՉ���z(�r6� ��ݒzz#� H�(0���vN�+]�2�I��1O�.������Y��6T�#g�g�<��0O��l:�Љ5?K�=!@��O�f|�xp�x^c��z����w��ۍ�!jH�J'>�'��@r0������a"x/w�E�#�F�2'
$Zb#G��FP����:d�MJ?�<]lQQ�RD���Q	e��Q���'�n]�������S��;g1
x$&����7�U]�ڭ�o'�>R{
	��B>(���d�Y�L(1�>9����ܛ����w�O�:Ѳ�2v�?k޸aܠ��a��Hĉ�0�h���V!��ZF�$�+��	���H+�U{�n�E"Ñ�RP"���g�����鵍��H�6v,G�xƠ78�|Φ,�Wk�)��<'�p��_Y�d�B ���VԳ��6�1�lN���d��~�vH|���6UPL\��"�=���/��CJ�J�bZLC�`�����KDaA���}5f�jh���|>�9��҈&�}~�쑋pT�~�+��C!�D�t����<�pO8l��=0�q�<s�v*�{ �D(�iO>�Ϛ����EkMX0��Hv`,�:'��o��	i�e�/�K�P�8_8mxXW�������I��	-"uW�U�K@ِA��?�2ħ��3�h̬�`�4�R��iS���w�nY2����*6«�X��8_o�ae�ꅍ�ޡ�N���1oB��:���H M?�f��b��IOÔH��p��~�������r�`�FsżH�+�>�4�!�@d�H38H=;�]�H=��}c���noI�C���{�����l��s��F*�/��ݒ	; 8D��x�49$e��,c�lD���)"C�TW�@��T��j��k�Δ>&D���ƾ<���ߛ�K�.�V�v�x�H��x�1@�D��k�_:v�6�E�$�c�K0(��þ�b�xH��r��Ä,͖cn����>�cti�!��K��Ay�5�=��,U|V$H�?Rt���O�p:#�zg}OM�_h��2SZ��˔#��jޮ&��:�ـ��nR;J��x�yhg��P�9!�O�;��:��Ϡ���l�7�.���(�
뀐3����W�����H� �HEH�*���Q^����$�}Q$��0>:Gv^�`n�PId� >w+��������k�.�l�s����z�'lHu�G�>�tH'S����N��
�#��.aJ���`ކ�6��Z�l�p�#��Kߍ��C}(�!���I��얆�a/�\��4�Y�2M�,4��d���y���+t����;��A#�`I�m Nz�UC鷣ׄ�<��$qq�v�'F� ����_]7$�H����G}���m�y8SJp�#����sw�c!��ӈ�=P���~���_{Ň�n9���p�%�!����Xy�E� q�7d�F��,���R��9<�^� �C~�W����~[��T&��x�q3����r�_:��N����$�Xe2C���TV|"��|��H1�,_���o0:���7:��-�r�η�']���N2��d$vV�Lә��[�+s�4e޵�t^��u��K7;��۷�B�׋��x�e�`tX	y O� 
�N$�j�ry�������M�ls[�}����� ��'+!ؗ�_�?x����d��x�.I�^�h�����o����b�{���Mcf��l��N�8���K�tU��6 H8�\'���[V�'����kg�	��I4Q�,�	7Ul�~$0{v]��!!@����g7^k�pvqW-v�l]�����p�f�n�b�B,ڮ1u�R�5�{�蟺�G]IP�B%�_T�ߦ����Iظ1u�o�y�p����Ϸ�va��A8Us�r�F�y �ۿ*�Y�;�ܨl5Ƞ'�g:�/o�V.�45�g-
0�qq�DD �{G���BgU�m���G�X}�l;XX���`tN9��* z�֧lH1���AJ�{�(P6>��@i!���
)B�wD&}r��� {$y-�/� 	��� %�	~��� w���P��v�"l�?D�������"v�!q��}���#SJ�s�;8��S�z�lݩ��~�~{�	��f2��\6Uq�r̄�ϱX�W��M.*r���!#���@@��E��@�w4U�s��>(��g� yԁ�ƚ$�>�udp�(�_-�I�';r ^~?>|��8΄�t��>S�ci�|s�@��>����K�4���r�JE��}b=^� Kp�&���vOs�a��ԁ��y*�	��H�� ) O$/qz*��'��Ό- |P�׸����������ҳ�gi���!�ȳ	�@�4�>�É_�ϳ�����- $E$O�:�ںvތ2�]���1�~�V�y�� ���N��U�j��+��������Z����vϏ%9T!ds��A�$D�1�$lom�@oz7i+���_~�]�TV]zJ^�^w}�٬*��K�p�ۖZ)����K�V��d�����ɔz�+�
>�»uR��۰C�=w�#,(���6��Mu�9^�[M�������r@ȃ�R¶a2�P�bR贚�h��KV��󳟆�;�����;	s�êR�`���p�Jn+��s�u�n;[
1��x�����N�Q��A@�\1��0u3H�=�㶭�零덁��H;[/\m�zc��8y^8וڝ;=\MCy\:G��ܶ��ڹ6�ږ�4�Q�q8�g�v�ن�-%�X��d,],�]sEkl��zG�cϢ�g5��0K�3_���~����'��x�#�q~[�Y=J����\$�A�>���`�G��8xl��8�#�p�jB�+�����L�s�'?`��� 3� �}�+��XY��� O��p���*�!ԏ����GjЮ�M����<����� I���!H�8^q����8(�F����lZ^���"~D4 �Vn1矻���|	��H��I0�F�8H9 `�1�K����~�"e�4I�\,p|�q9��u�<�g����}�'��;���mԈ,=���ߒ�����l�����[e� �P䐞bFD���j�cx𑎁8Q �:�	R3���Ͼ��邢eE}�	�r����f�iE&��S���c�����dD�N�	��$H�n|n���d�A/�ƸG�{X���;Ч��3Y�ͲVHĉ�U����Wݗ���?���t��
 �,|q�"A"�C�W�hp �0��L�mp��ʇ�:z�h�"I��r�Q>u���^�G2�4�i�\�`ghYS��t���7��NA|�0�!��.H���m�r���!�"!p863\Y<k��+�_9:����/�*P�i28�P&* .׽+9�G4�C���TGiw6�XޠF���a�֍��:�סl��-���.�h ��y�:m��B������&z�%�MjՋq{�i��`*  +ޙ�;� QE�r���hQ��(��B�Y�ׁ���������HlW9g� ���Y�Bp�C�x�Om�(�#⡙~ Ƞ�#"$7��s��c�� "��s��\�\6���rXÛ���j��\S��s���f�1�Dޫ���f+̽�d��ʒ��oW&l�y�ڳ��4������Z����ʥ�'�q�W(�	�f��5s�X�i Su]y1F�da��,�5��_�s  i�^�)u�~�\y��p�O�3E�N��[����9����������='��~Y��O�N�d������� )�Q&��rwO�!���Mf��i� xz�p�P�$
\U�9�$�}��?�!����C]�����3��s"�S�9v9d�W���h=`Y�|���^_�pX:y� 0x4�SD�.얪�"yS��iw�m���4�y�@��_E���79��O1�������S5.v��v�sÜ���Q\=�����dvB�d�s׀x[��H��T����56�����\�N"@�����<��9�6�� �.�z�c�̳�Ĉ�9Dl��r��o"ġ*��.C
L8[D�K�l�P=��$ml�AcX�y��
5*��ں�,�Ԯ՗Z����'�t):;�����j�yb���\��@|$�v�}�i��< i��'b�/�3�rS�٧��@�W�O9L.a����G4�.- 4��\�8�x{^!�Q�\p �pF�#�Grx{=�C�*Ͱf��ݬs�+x�` ,"�3y�%c�(���
3��x}��\��-<��(<����sء<��<�je�,��~�� ����-w���t�`l�;i��H� !�>� ��"#�W>�$� t����Y #��� �u ,���z)��f��Gp��Ū�@���.Yn�В��@QjC��W�6��ghؽ�|�������F��c�ަ.�j֛��x"��� f�/���Ϝ���<x��G#�����^йΜ�C�N|r�I�9#����M���S��1�|���@�Y`a tB�oEr�gu��^O)#�s|����0�@Y��#���=�Z�r�8��`�y�as�@�h�|$�<���di�^;�ΐ����_WtЪ!p�<g�Z�9��	ǯ��_>ck�Bc\,|4�0������d � =�r�@|Q�
<�"���dq�+w$���'7�O{����(��G�~���=n��s8!���H��#����C��#����G+�Dp2&6"��?�����+���y�g��3��5�´��R��Î�T�ufۗ��Wvn:n&�n:��tpi�̨�dpu�is��.����8AEQ�8�@���hpOE�5�@y�*H9g��y��@�s'}��*���q^��󧃘C � G<#����{����HHD���<���,󋇛\����qB�F(�NK�<xz�9�P�9g�������)�ԇ{��n�pp�"Hi ��Bhi���g�����G��9G��p��j�(��C�0�y� �״Wqr� �8:a2�^�V��x!���s�h��ve-�B�K[�RsÜ����9A�h0� ��8���\��+$�yg�0u&� y�G�z�sH��di��J�g�r����s�v����$<x0�;+�i���9�ܪ��y��*�@�x�o�|��ƃ`��
H��@{G�x�NK����pt�QH��T8,�s�� (�	
�����,��| a�����Oq��@< �a�9G���Drw��<n��o���p,���6q,$�P�v�t��Hb���M��@J���0�+w�_5x�yB<�W��<�q)��ݰ�A�y�-�P s� ��!�:x!x f1:?�O&�X˦�ݻ����/%e�9�39� �߽+��#A�y�bC� ��]�P��2��pr� (�x9���9��W�p��� �" ��4����f����#���q��pi����p?#z��2D��m���3��3X�)mY��V�Ei���f���7J�f��т�.��;�O	���9���9� |DQ{s���$�:@��\���us�Y�� �8~�J��W�]�
��������sZ ���\���G�����qw�+�S;75��9'�$���s�Òs� #��yP���K��e�,��G!�0�pQ��7��U�����g��O �9�Ds�{pp�� pQ���r���Ub�� ptUT�̾�4:�@�9�y��p#��ў�"F"�#H@��Rs���t'9NOy�LNN�m�zW8 ����s #�G9���J��0�pQy���k`�� 
$�s�U^t9��xO88(�Q�\�<� wkʀ�:G<���x �
~8�N@�RE@pa��y����%\��]V��9�m�h�80�g����������Ξt�x8:x �5�,��y�� 4���CL2��l��ߥa � "<�<�e��&(L�`��\�0�ǀY�9͵�<�z��9�<���~��5R�u���Ƙe��!�jg2ｕc��8 ��9�� �s����� s���8 ��9�X�  s��?��  s��  s��?�s� 9�s��\ �s���$����I��Ns�����$�s��?�9�$��9��� s��Ü �s�C� �s��pp 9�s��p 9�s�p 9�s��p 9�s�G8 ��9��8 ��9��p 9�s8���9���e5���R@`]� ?�r 	 r}�"A����֊:2�@�EP ͪF�B֔T�m�kRP��T��kMf��٭5�h��hiE:99e�7[wV���5*�廸$P��         �                          �        :>�4�K���ն��l��.}ܠ�,��v�oH�S�))' �z���� r�Ck=<�G����w��^�t��5OC��nx xt5�''�=�����;��UE��   y     {� q      w� �     1 �`    y�7o\��΃��K��H����@/\� �����=�]Ѷ��=��;�U�����MM�nWM �z�*���`��        +OT\Z���l(�����{�gg@��hcͩ=^�u=p ݊�+����;��ʨ������q�˓����� Ǟ�4�q�y��ʵ���B��,+��ZKŪ�k��۸:�/ ��*
�-S��
��<�ҍ�q��x��AJ�����u�޽�]� ��ٕR���b�+�rq[�ݍk���ŕB�����         .TuKnZ9j�Z�5\M�9�oy㽚�V8 ˶�sd�h�\��m�9�ٱ��j�M7 ��j��Ö�Mr�h�Ff �A�;�њ�w4��j� ;�Vq��57;�Y����{ԥ��7vV�h� ;]��8�͛m���'+8��+m�i�R�H��(�        ��k\Gq��K�wl`�ڻYk�B�َ rG,���m��v�Y[s���j�n8]6m� �鴷u�ճ[�T@:&Ɗ ښܵI9�\�R�P� 6�U5ˮ�iW)͖�u*S��ju��p ��cn]p6k\��c[[r�t�7v��f�J�CTS\        ���<��ˆ��\����Eͥrҭ�t��m�n ө4������mr��e�\M�PYs7m��\ k��[���[[r�If�P�UˮUmYq��f�2� ']q��U�kqp�d�cGL�.A�YS. �:d���W�֒6�M.��ƛ[�{{�+R���������IT� h S�i�)U  h 5RК0��A���=�=�� ��4   j��T�P� h S� �����1={c�~���y���w[[馶y�6���qmc|i>H��ӡ�	�#�L�o�_���P�ֳ͖=�D��!AԡA��P���%*����\1$$�	B��EQTUHZ�UUUUO�1���cj��܊������H�QTiUTU�U��L��ߐT#�5i?X�{��{�:�ߵl{�A�am�8������t(ø�ot9.�\��dd��&�K����tfGe���I�BҬ$走�Nid
ݙ+v�I�N�%�����ٺ�oyȭ��r67q��J��n{��da�*֞>{��Q�0ݽYX����xpr��<1�l�^�P����+>)J�@۵1��Sʹi��Jagj3�h�4���6nЉ	!�r��p��6��È��(�
S�x��M9EmY�wem&����sV�wm�]V���[0�֡ˣ�>b��.?�Dt�}U�;8��w�͖G"lR��ȏd�|�U�WA�Hb�13E��w�\;�N��o�?i�8�`e�XRm��5\�wó�:�+/-��`R�V�r'S[�ir�nn�3֍��F�d_:�Խ#6[�m�M4��&���-��g,ja�c�TٵN�Fѧ����KSv�̤M�ºQ��ɹn�6�s,f��E��'3#��;�|�q�w3Ht��,�ah4ST�!Ŭ�R��B���nA�X#��Su[�26�Y�+p�Y�*�Ԭv��1���1'8*�	�f��툺u�b.��%��q��p�V�R�`N֠�K�Un��n�0�4��c��Gs�"����o�n*�hYYB@sϔ�nH7]���ӣG��q��^��%ԭט����Ս[μ�@Ź�:�S]�u_eh����W�m�?���-�T�&!��N΅6	�iu��f+h���2����ǒ���ɕx�e˖�5M;T��\H�/�x���(]�}$f<Ȍr!z��Sa�C`�B��=�[�&��Q�2R��F&�۶�uA��\VV�p��KN�r�gZ
��G�"乻f��l�t19�J�f٦0*��͙��H�.���%�}v.'���Ne	n��bf��w��d�Fýyy���#�a�3V&^�ۭ,×���)�Yz%����j{��Nd�+�r�jU*B��1/��*9�[0l�;h+wJҪ�tCNZ�Q���gKJLn��p������+
��iA�,!F)ױ�"U�`n���`�R�ru51{	��š_���:���`��ܑ�'%$7TS7o6`3snh��6��m'^@woc�Q\
�ۥN�5�V��&�nk��f��y�K�˘ۥ��E�ܣC1͕5TwG:�NU�P����Y�9gd���Q>����x'�s�[o4Dp<cm�E�>LP<.�INnR��f�^]������*��sV	����T;P�a�#m3*�̓�1��e�u����{Fa�i)���D֘3U6R�c+Т�����r�*@�{K�n��7GAy-!IZ��ܰ���5��L�nF�T1iBU�z��:��SE-&�{n��R��/M��D�@�,P���Z�b�j&�J����P�麍�+Aneiٯ���W�*4m̙RΓ�*�9�e��cuq��r2.刬L�&��O1�e+a��IÑw�����[�҄�^�Փnm�(����HhH�f���*Ut�������X��t��ٻ�U��Y��{Ya�ݻ!*����G��0R̘�4U�a�iS��L�Q\Ff�!Sj�9&![k�f�2�ˮ׽{g!b�,
�2袍%�
���!p,4�`L*�A�a`Y�f�[Z>tU�킄j�E�9yZ(�R�jf\�L���9u4������Ҝ�>�iտ�!Ți��)�;F�UX`rƖ1'��VE�/Kƕ[�Y�`&�bd�2�����K2�b��a�9�@Џf��ۗ�hG�A�Iә��Vʛv%����/@6Na���@Wf�<m��p�t���v,��{�x��2p�_�x���ݩoC:�0`��KA:�`�yf���/rmIE������V�w�R�l+���C�,��&u��L�.V;͆�/&m8�������"�y�蘓�5����3�5[:�R���P�\pu1JJ���,9H���./��
v�%)*So�;�ZAчvh˪�{�M�������b��nHC),s�T5��}��0bDb=�@27��w��f����k\��������׮��4r�ԩ`���#Ґ��&�e0YX���w�d̈́E�e��X�i\kP���KK3p��n:�Ku�5���­M��m�`�7P��:�q��C� |g��*�h{��vV�).�lרn&0҅��Ȭ�Up�l�z)�y���D�8��e&,�,R ���{�	9Oiv���;�=�A��^�K q&��$�&�M��#vFKV/E��Hgx�����n�ؖ�I�����-��m�m��{8}L���̲*V�iV�B$x���Z��h�ϕ�L��b
n s���-�-h����-�bn��ɷ�襳j�=PV1�Ym�E��6o`���m*Ɂ?h��U5�2nǐ;��S�&�e� ���N��94#J��ɏ@b��S�d*�yjJ0�!�H�R�)!MV��t-��>.�^7��i-E�l�汊���TBi�+�l��L/3n��X&�2V�oVR��!�qBê"Z'.S��z��$�����JzQ5 �[a�$arѠk�c��j�"E��w�iV,�L%+7J�EQjZ����.�M'h��m��F$6lC�᫬�[f�'�[{+h�'�fG
��`
+o�<�j̽��V{9
z�o�R�P�]o���2��۬��JΉ[a�:n7�t[yW$��\X>�N�=jVݺ�"euB2���	�tJ���Ъ��F�ѻvU��G���^,�h&�5N���M��.��'4=�&��f��e�*)�5n�"�٘m�a�(.��n]ѧ�#6/Qh��s&�AYt�F�8c����lm;Id�B��c8Bz�d^�������N`�$�{�ہ啗�;Gǜ����m�#���T��ei,լ�i��eS�V2�%�T����tw$���^H֧�q��K�rlku
�����P�'r�2�9Y��yY@�Y����:�AmU��Xw`"�eF�{h�Y֢�-�--fꜺQ��5���wh�5*�	��'e�\-:/wq�0Eu�(�[�,�	ad��/�+\�t��A*�e9���b�D����52�)Hj���+\Y��˪���SCĝ�-I�u���+���:�wC��N׊֙i���5���mu��eo�l�u٭��t�Ϋ�*�wE�'b0ça+/w�����	a��݊��)�'5'������X�{F��x�I��V��oF�X���n�D_��,!��y�i$�%�i�2�������x¥%Jԅ�+�9J�Uҫ!֌����x["��"�`�����`Ze�}r�A��Ux�� )���.��o�X�l��OPcX'B�ͽA��l2�]U�� �65���z^����K=-A'����L�[Sd&BX�f��Zi�bteۄM#M�\�'���l_�N���h�]�Z��<�l�oe�KKQcbu�Ehxwq[o�Ӳ�S�T�f��+c%��Y��%�;/��,]U��*��/����>�Y�>[��R;7*i8��$�5X�F���r�%�L�)#��\�As(��^��.�i��\8[�%�՟:�,K�~�>��pw�_1~�C����=���5�m*��������E�jHhLЈ��ZR��U�&�Cc#��A"�N^KrRDd�TB��QQ@Ǟ���-�|>�0
��2��iꪫ��������P�y6/T�B�Şf�S����e\�kv"���S5o�-����G]�U��e�Fm���1�䕒m˽W��i>�܅�xu�fYQ5z�
��_Ufm�_"!Xv�J���M�5�
�~�TT�=&�5:�mVnU�$d\@p�b$�ӕ�q��l����p�Gզ�m=&c�|:�u�a}dV�E`��Z��m�b��s��=E˅p�8]�ݠN��K6յ�c	���)�L!U�)N�Q˨�YM���	B�mԴ�\�g��`בֿ+��H�7�.˾�XL�|���O/��w�p������8��[ݍ�G�Wԑb�b����5�k�9G2"4��Ŝ�n�[���k.%_���ѧN[�@w�-�Պhh��n���[�M�Ҥ��Ym0�l�:.]�;vβ�����X�(fNJq~F'�^S�C"�t�',[�U����֝T� ־e�l�ai��L�I�{L:D쬭�/m��3L6�2��*y�nm�o�2L�/�v��X�����y5�5���ҷZ�i[��p�[��F���SsF��ֻ.�m(���9�T���g�=��9CZ6�|f,̗&mP��#/�p�@/�L�q)�)��:6\�(2��U+P�adǄ�[ �!<�Yu�]p=�R��[�vLJ�۷[u���X�0���u���r�ks���0����; �a�m�YuoY��0�5��L5�q ,Q�b/����]APڛfr'�%R�Qq�F�o#p�{(p��V�9�����Ybd?*0��ј�E�%v�c[�Ĭ��E��L7�54jЎ|�4�٬�i���#�ѳX�/n�h�N/��s��N�`�2ᦲ�5)V�p-�`��dM7/����Ȗl�z�Ϣ�2�R�Hȼ ��,ЛP
!��J�͖�n��� *�2M��ۉ:`�je��Y��^"�j��]]��Kd� J��V��f��
c�f�m�L(*�*4Ю���Y����p�pA�+w�$�\�i����sr�Sb/�E�]n�BSO~#AO&zDw�H+�(��z��@�㣤	�(���i�0���zi��=�Vn'm�NV��ሠV��j�`�F~s�4	WB��[��)��L0���nAcwn9Rd�V�F�
�T�F���z�\�0<u��%�2$�"�b4�fڈ�-7V��Z�ͳ�;j�2�5�E ٙ3Z'+��5)��j$bN����_��:W;�e"�k�ٮ�\�*��c���ӹY�LJ��*��٢��ު���׻:�v(M8S�K��ku9�R����m���>7([��t�S���wSlİE��9`�ծ���kĞQC7��t�m�dVH1��9���n�۩2��!v�wv���g2Z=�jk7[���\w)���#6�5��$s��E�mwP�ܼ@��QJ�cמ�UB�}� d&߆ɑ̣5ٴ���7]���kCE�2��&mE��f۬�tDMN&�6��B+6LS�In)d�u/i]�V��J����Ka{`Ɛ�k3���g����累i]<.��ړ;YLR�ܠ:�畜�o�Q ���W�y��ʭ�g�6��WGU�Y+.�>J�4�P�u��}�Q��;�u_%4V��2�;(����Q|��� g�1�%dO3x^ݤ>����׽U���3�A�cr�נ��=�=,���"s1X@Z���e��_�tLr��r㿵���I۩�F5F��mm#^�kv����}�4C[��
��	u1��C�ϰW��A�A�ĉPU��F�}��
"��[`�lqj� �ȷh}��7u���m��]�PIhs��DϽr���e�7���k|�}���נ��Q�qp�$��<���t��AS�����"Ok ��n��6g��᥏%`#qN��C�s{S>����ƒG7��T��+�>�eqr��m���F"�XܹoP��u�ۜz�����*��e�:�`(��;m�|�X�dyt$���~���/�B����g�����6l=�49ٺ�`g&�����{�4;J�����L}wdK����r��tv`��[�t�Jp����ٌuѥSM����j��,��=1A��;X^79Z*�Y��5�A���l����#���&�H�&V�G6 �o5TF��V��������.6���S�J��v"u�J*_2���
|�_;��c�f���<h�J���8ڭɌX��ڕ���((I9u�hU�ķ�����ա�pժ�~�Ϟ.�I�=����f�54�KXuV�V�l�6�I-c'u�Cg72����MM��܆fSw �F�u�!�#�wV�h�]b�=��:t�m:��B���Τ~ֺ�N�h�5�n�|��@\���>���������nEu��o��@6��:�O�dw&"�jp0,i�ѕmޢ����f����|d�n�"�.��}b��K����3��E�ǹ*�ߺ�~����ͶQ�����`�i�m\a�*��YtI��n�@L���pc�$�є�y�m�q��VfT�X���u�����)��%����9n`��?\5��2�����V�eYTm���M�жE�m�LCfe*��IJ�Kz� ���fi
�c�u̽ڄl�S��ӬR��� �4MA�,m�Fܭ�sL_��?}��
���מ	bP����3��$w�<����)�;��W��ye�`�	�2��v��ctA0iV��Pr���{n�-�����:J����R�iW���o� ��D�)^�8�ϰ�Nf%�Ƞ��LYk0���h�o�T�ʚ�"�ӬOE`F����Z��Gmj�5
!M%a��:�*SV��F�,I��H��
�LGY�!�*�L�f2�y�6�M��i\�b��-�i٢YHƞ�����R�*��Z�����[��ǔܥl�˫�G�f�LJMzK�lG�^�iu"I�0洚C+�b$�M�%It���>�k/2����c\��5k�;��E�h*�e4�Ǳ�}{�b�w7Cg���>"�䣍�#qĚ0��)�����E�
������ꪨ
��V�$�UP��B�y�M6ڥ�n�e���V��iV����
�	���KmR��G�[@R��]�j�kj��j���������a[f�Z�������Z����MQEKPU�Q{ ��Z�i^���Tv�h8W��[(�UUU]T�U!�z�X� �U-���>���d���jHj�eU��RUJ�R�H\�U]*� j*��jU�:���V��UUUU*�UUPUJ��UUJ�R�R�T�mU*�UUR�UT�P�Z��^�MruT�@@uuPUT�UOZ�����X-�)V��"d���B�-URD�q+UR��WKUJ�W*�hW��UUU@URJ���.� 4�WC�n� ��[MVw�%�K�gT���U]UWU[t�+ge�R�K԰��5�Q1�k�T\��[E[Jp-J�UJ�X�%���`��j��Pm᪩	��Vݪ�Ԁ�Uz��CE湑zc�����I�����P&z6�h���p������6$Z� vx�6��n��z.���Z��7p8չ�v�a��kv��{b;��Ů�1t/*f���{n�R<�3٧v5�p�8R�us�e��If�<�b+�{q��qę��yA�·\mн�q[tq����-�튰��d��M/�s��c��Ku��ō�o'5m۩��-m7)I^6Ωz��k��c��v��nrQ�ކ��7��m<!;y�.�n7@z���e9/)ax���q�����[]�0��c��ƻUr���Y�u��מ�N����76�;��w�=;�xÎ��Di��mچN����TEqѵ�q����J�s�f�e�,s.��M�n�o/k��e�pv�b�}�rnܤ<"��%w��興�gX�l��xi�pA޻nɺq��tp�{[N�N���t�J�1��R����I��ܼ�!�i��fw<���k&���wU�d.9h�J=p�����1��7c���v֛mۮv�z8��v7d��]�uV�pM�]YR�LGT��V��ó��� S��y�����\�������ߓ�ݾ�;)��`M�n�vC�bޛ<v��nN�e-ױ�➐$�ϳ��,��uv����"=Y'��ۯF�_ݯ��m.t&���ݎ�[����Ͳ�q�ˀ�{<�V���pg�����w�W��0����!��X睋f�q��Wk���ƞ�q@l	��.{<vn�2vዝ�n�-�,�Fpi��I�!س%�%�v6��Wqvm���V�x^��ݠ�&���G����n����wK���W�XIg���t��9�ێ�낋(z��Y����x<�b�ݻEV���toc't!�������m����p��S�\w:��O5ٞIѮ��;n%χ�4�۶g�6͆97=�h4���7���:�m{\��:��x9�IM�f�u���1e��`1<��ɷD�qv��C��x���m<]�Q�,�)
�	�-��Oi�;a���;9�ݔ�8�qL��Éͅu�dG��9���b�7%��Wu������#����B�'e2���s��/K������ufN�,�<�\�n�$�-^;��H�m۷v��݋]�u�H'v��nu�y^=�h����^\봖�n����v��nL�{���q�h��<���R٭kn9�����q҇��v�nx'�>����^��:���sy�ģ���L��J�{3�;�׵[�=��8�ِݵ�!0:�`�ۄ�qV֮�]��"��؎��A��=X��p�9C<�>^���.�;��n�;��/J�9�v����.��Hw`w?B(����ދ/WXSon������q:��-�v�f��p�Ͷ��k�X�8G=�U��щ�;Gn휷n{<�'Q�uu�c�-ڶ��h�80����(�gS�~���NG�c���I����#u�kX�nL:�=8���X��k��v��)��3t���-�ru�2Yz���fڮ�h�ō����0�;ur�Ͷ5���h����n:���i�.7l�6�îz�ÈFU�u�a-ë�n�F�;�﷾{�KL���l�Dw#<O��;��b^�Wi#g�5��v��v�^��[����56��5��[mv�d��p��vݎ���t"��9������CZ8�r��W�����ڸ��Y�t��Q\<mO\������v�����u�by_c���X�6�z���w�g���v�N��Z;D�r�6�p�a�qg�9�tʁW<y�FC�e�x��ܗgz��٫�������o��:K���7e.lj�bC��7����Jr�;����/'m���u�j��<]E5vOm��8۲�S�7A����y�����wO�\@Ýˑ^m���e�o(�����5�S�{������v����������KcnG#�ێٳ�nwp�X���s�/Z��:��.��.���u�'��,m�]�];o�ݚ�N{V��9ェ���]�t�t;q�v�uG[�Þ��pts��]�y�RoG.�v!{��������f^g��d��^��QvC�^qpt�3��ӎ݌n���k�z۰��ٺ�ѓ��ܖ��f�m�ٌez�pm�7����bt�#ۓtN�u�#���ۮ,Eݜu�R0��|��pV���Z������]��y�v��lj��õ�8�:k-Ƚ�`k�wn{f��vUݥ��ϱ��:z�e`�Q�Kf�1;��ۛs��Q:��qj�nu����F�m��&�2�f��W"S�����y�������kZ������͹4��c�m՞j�{m�밸;s���V΂�`z�u���{p[�wr\�dyzӷ����&N���h9�<�����^د:�u�듶��W<6���ڻv����=V��%WY���<�����6��*v���[wiv��&!��aش%��<t
N�v:��5�޸\r����j1�sٞ+�ѭ���q�)�vqulj{]��P����c�L��<��v�<�X�Ng<<��dn'�y)�p��]��ll���v����p�d�vi��������.�F��6��<9�q�k���mTv";����� Z��ɑ'�!��v-�e3�kawC\��rnҘ��\�i���c���XN^o��q��[L�ľ��Z��n6Ů�s�� ���:/�:Hz�0���g�zt���ȔN[��}&nn�㑞��k��b1��|�u�nFn�m�eU�;{uNg��7l�͒��N-��۹���^x@�Ǧ������DM�[�|����^pm�t�z�U���	ۺ��;g�ې�̂{gm��\V�J<vx6���mVl��f^R9��m����^�nt8ϳ�v���������Z^�FW�:zmu :R��5��l�z�h}c�ێ�^�N�y��1�Rj1-لc�f�n=МAmB�+����;q�p��#��#*y���ⱣH�w!{q��;gp��v�9���.�*[���r�w9�'��I�4v��Afq�[�^vL���.�;��5c�&3�&����E�1sE��f�ݑ��ݭ��4���[k����9ݺ��{��W�n��<��+�Ӆ��![{N�z�G	��۷#�Ul�c����u�s��a{�q�r���k�/^nD�ķJ������\�8����Ol����Ƶp����#�7=d�>MMqk��;��X�����N\)YZ�&���ļ�'Qu�8��'����!gg
s��;m�
۞^��g�v�{�v��y���X˜h<�]�a��\�,�g��5kW6WA�5��7<�:��j�B�G����n��9�˼���Dz��p9�g�5dۓt��痒��H��r12ơ�r�p��L+��U�nƴvy�zŭ���X��_iu�y�� nv,��Nb��wfZ��i�p9N�������#sl�p��d��]���l+ٻ���و��cZ^����u�a8J<�ק=�ӕ��r��mέ��K�=sl=Cy���9:�̽�=��V}u�m����;)�i�b�9:��m�s�Y�g[k�L=�zoF�.����{:b1��3���jq�7d�y���X����\�FS#��X���ۉƯ9^�	%#]$
}jC�n�&^�O4�u�*�}��WB ��`��xA�b�6\�te�x��͎��{���>�{n���8��������;l����vwl�k/US=��c�ԑ��^��gQ��Α�m�A�N�4UtY^;g$�uݼ�7��s;l.Cnl����)N����ƛq��ԃu�ˎG#��#�7qרw[y�K�K�n��a��vNp"��C8��Vl�=��!w>˺1�N�Gm����2�ny��۲ams�!�ι<t\������{a�۳�tz�6m��Q�n]�u�vK�ی�&�:�Oks��Kp�˄�ۊޥ載��H4��拷[]M��䭢͞�v�l����|r�[�L΄��y�k���%���qƺ���I�gnǝ�2��J����v����7��rG}�9y1n�|�Οe��N�)�k]�۹ö��n��d��g��Ǳԧ�/ <��b%�]��te0K��#mn����s�6������m�qӌ#ۉ;d�ە�̪w"��ڙ%�eJx�>1ck��Dk	�WWI���o���]��%�=s�E�:'�Z�Ym�zW��㸓��RY�Z�v����M{+��r::���y;���;b9ql7]�g\a|n��qI�\��󣝈���Άϝb�D0���\]���7��Л�����!��q�*�ݰ��{u۬�ft�:ls�G0��WnMr�s��<-lp�Hn��v:�&ynl;�x�:�R�닎f2�R���w]���{E=;ۺ��#K�h�絳�Rۭ�h������}?;��j.�\��D�]���g,�;h ���g�M�������l)�d��F��\���]J=Hu�musљ�R��NJuƌ�Em�ow��{��,^�5��"� ��r�� �R&�u��\t�m��MY�v��;��IJ�����*��q/h�4��D�T峣zd�ب��7T� �O3s�����VV�UU�H���l�9��5���I���f�6�tc��M�<m]u5v��+��8��:�Q�������vѻp�>ۆ�SQ�n�C\����y��q��Wn�i��V4���M�����ܭ�ꎺ��N8���Z�r�n�0r��=nշ���[�X��gzt��E���j�KaܻƄ�	��t��	���Z��ɐ9�������9��u�s2��':t�6��Yc9���j۝���[0��Z�r�_=��g�G��J��[�k�I�8�/�n7��(rk�1e�&�����s�����v�+t�nn0�{g�\qG�����^�֪��D�=�v��\�-��v�3�Pz� ��=���xMvܹ�nH��=\޺kt�M��f�ڜ��Y���v�3�mF�u�u����<��,��m)cq�4���H^��n�����qj�臵�sgv�'�N#sz9z��h��/��0���8,�%ra9u�on5+�n�Lg�4���{G&�L��[�+�k�.�Z�۫���O7�٩�Д�J�t76�n=��s�7YnW��[F��Eb5d�c����A��˛�mq�;�����:�]��v�*��=9����^�'���'H���=���!뒶ٶ�Vv<��F�(|m[���'3vmf�6�;q��{uc>�v����:Y��=v�u�c�G��ƺ���`֊�E��9֣<k` ���,ok]\�s�z��4������#�:ۥ��ŵ��I%ΰ\���H��	x�h2mn���qnY��n5gnvC[���\��9�6�u�y�y�#L�Î�:;<c�'m�s�q�U�WV;�����Ȇ���#�l�j�˕��vA�$��N�k��X�U��]��8�o=΄��5�(�At��z�nS;'U:��r�O��+�M��G�����b�a!8EU�U}z����r점�KUKd�^�ʤ�z���˝����\��X]gZP2=�bnf�w�ka��n�)�;��fo/6lGV�ٮ����^��Ŝ�
��۸�n8�!�aܳ��b�Ԙ�^q���v��0ے�q�q&Ƕ�=i��m��w
(/,,:;<N{���Ż���{���5���x���J�-��7n����d�ַ��nܻ��6���|��qÃ�g���d���63���y9.96{\�M�/��E��q����?XhY�^�r("oY�k�a{�V�dQ��9>>�z�>LI��w[zDSP��;���}0Ј���V���D�/܆S!B���Ј��^�2.��N�
m!n��{6l��;��5�c�
�+�k�Ooٚ�v0Q�^1S$E}��ɣv�@��h$'ܳMA�]��@�$6�{�گ'�4��w��I3<4n���,��-������a7%F*�/�]5�����мHR3�e�d��ޗ/ޘi^�SY:����IH��89���?vu�C���*��k=�ٺ����҂"m%�=e�def\H��b"��Pᕮ�飭�v1�;�Mmi�[�9 ���'��օ���w-3)hi�����
8� ���4Bʕ�R���u�'C;Mq�}Ĉ��Q�&r�B>���:Y�p�2�s{D:�0롵�Y>�߬�rAԂ���F�~���1b���9Ǹ��vA�A�:n A$� �W���n���*�����X�1{~���$DD��x)�:�c��i�e�pZ�o#M�l0`���A����ڷ$a�����gk<z3���N��SWAm��.ܗ�wp���nE��"���g�팓���K��c��hw"*4�Jd�kޙ�����d7�e0H4jF
(6�<��őj|�l�q�1S$V{��]���i3$��$��M��DZ�	ſuIB� �V5_>��Tr[�Y�U��	F.��|�|�f����d�IԛӐ��Da�&����*�X��)��v�'����b^� 6�;k�$]:0)*l0H�}��A);�"VB75z�'$��ndnT�}�MN ����u���P\Q7�6ř��]�0�R<b}'X);e�H���:�B��d K
XHC����� b@���L��c��1 T����5�w=u��#J
j2$[� ����p�A��A�j�#�	21��.^d�7�6���ӿ�7��N��g9
�2�]�/�vR!�W��ݒ~��ZU ��IkD�],1���4�hH~D��?�³�T=��������Ҧ��Eޮ�{��#���d���n1H�1 �I1�����_�[^K��l���4�iR�k�o\��ߵU\�"y�	 �1� ~��|�fު�dB�!<�F�Y�&�%�="�x�G�H�OD!� ��	u!����Ͳ���mA��K���s�ɫ��q��2޷�[��q�ú̥�����Yӓa~����ߤ��A��d���w��������$��$J쑺_�$���h#T��y�!D�5�خ�A��"�#R+�"���*���/{o���SI�1}����m������	v�`���fm�$U��Ԕ�{�����hjI�E�pBM8�B����E�	�e��-���M��4���ƴQy �"�J���f�"�A��o���^ɴ	�ыԡ�H�g�Ġ�8��-��F�Wp�j�ޚ�4�#	�R����Y�n��Z�]�Q,���ͿW6l�c୭����C%��%"M�f�:��O$,��tefnR$�*_ܖ)B*�uK�wvIy�f�%{�� ����S��FFT�Z^:�
}�s�U��b*&"��5h��dDa�FIN1@�(�������x��;�߽�~J��^��c\��.<��ҷrG���B:pO�U �Yf��ά�I ��mYd�z�t��ȂF,�b�0�ˁ�V�H$�G��6K.H�i��J�q6R⨠LC�m ���(�č�5�$������=��M|`�Ι齯%E2u�nȷ����r�S�ua��z�MH:�s�kn���5�jԑ5x���xz����ND���w�*E�ͷf���ښ���K���՞ݧ���y��3vG˔�r6�y3�O$�OH0���6m�vW*w� ��ND���Qg�>b�M"�����6Oܐ�g\�I17��g^�k>����� ܻ>b���يu��E���*ﯡm@�1�M�F�͝BET�=3�����3Ҕ}�:�X>��4.{��}(�KlF�]�e�j�V(f4X%�H�L�H'��Z�d�I�[V7�1bA��k�5���p��ʧF�{���;�~-߮Q��=�ѳ�o�ر��l6=�ܛ\�0�0#���� \H���{o�?"D;��6�҉?R��R����L��Il-�}���,[�&]�\	 �h�D&���h��MJ�u����]B"p�3J�x��R��:aq~��׭�eA��5�A�30��z�R�/�0躠A��{��y
�lo���ٺe�0�X;��VN�-dq���L���u�����l�ٔji\^>�t�7�E��f�5��G{��3�9�@~��eN,4���Б�s3b�e��E�m��{~�^���G'B�MΥ^w���ӽ`V\3��>`�7"f}�:�;�˔d�Td��0�D����3�bс���A�8����n���M4I�ß(c�7��s֯L9�� k�0q�x��_Fܻ���n���3~;�����d�F/�|�����P��ē�;�`��A$�I�_&���Qtl�U�L���h�恨�2���NA1D�ԉ���`�� Ȃ���b��X�Iy<P�(���Ƭ�C�����s�<F�Ӝ�
���%��ic
�3��:�&w^�o7$mK���0S�^�
��M�����gp���m�+����%�6Ō�̽�{*;�F��o__���+�k�����J��^�t��d���6U�)�~�$�d��W�:|��K���S���!v[�M}��[efS��"Ș��S$�I~�X2�J=��IA��mB)��_K��|�~L�KNȍ{D�o^�og��-Q��L{��ٓ��x7|-ߣ�H(߱�-[�A|L�C���q"�a�K����\�Fu�8��gJ�gRrEzƴ����͋�����v�"h������4� �D+h­���Q�	 ��AE���!��cKKi�m�5 (�=~o����[��y��-6���hb1�4�;{rEف,Y�ޛ�vou� �G��2^Y�J��۰��J�V�����Ȃ��˺	#��gT[n������1�rn�>sa���s�|OQ�L����6l�c#ˍښ�N�t9�\n�FǓ!��GV|�[�cU�8�]5��i&9 �8��ƣ�/\mڹy��"C)�3�Ѻ������n�����<�� �=���V��{oZ}Jv����[�69Mf�z��k�[l�N{;��ظ�/�n	�����8�.N:�Dvܯ���s��3�E�ފ8�x�f����~�%"T����2L���/��'Ƶ��P�$�"L�B����h ~+p�D��1חJ�|�����	&�z���@�{���A�6R���(B����ٍ�JB�8�6��N1�8ਙ	�?��<lǛ��5��8�I#�����C`C	u#i�Ku�Jf�t��c�d�^��x��|9�#c�=[[�&H���R�d��	��r?��p�N_1f����f�"�{���_��V�9"�sz>�y�-.A�5s;�{3��+�$��!�8��gJ��u#-�Me��y)�T.8$��IɣH?D(��k�Pc�%�ַ��'�B&Iʤ��pAN��Y/[!����d<��O�H<`��k^\i��	���k�H9�a�
��C֢�"'�)��@�)��(��LT�*��b�B�.�Q4E����y��	 �+���X�֯��	�o٭�H*���i�d�U�P�\'�`�&�&���g��c/���6�a�T�@�'lgm��+���)���nx�s�m�I�o8��6q�$ENOX�.�����ΌY�I�~F��(ń=���_2�Q&��Q�j�{������a6,��� ���wE_�u(P%S��!Qi�L�"�^p�~E$Hq��t����?�������hK�6�BQ�!�
~�"26N�e\]d�c��8����E���������O�QIA�,�zŝ7��	ܮ�$�G|�o^߳{����F1��t�8p��弔�X�� �(���Fi��=�HT|Ӎ6#qU�Aj�i)��Lv��g�e��
=��g$W�A������dW�����4�S��f�4	�I"���mwM����q[4�)�	˺�l2э�H��#	8P& �nj&c�=�(+���n����.;� $��K>$�p�����'��njڊ$���9#[ޛ@W{qp����\?:5��\�'L�/P�H��E�"��)��(��ч	F�����x4{�ޟ!b�<^�0����+��ҍ�;�
��t��A/��-�7�?\[���@1P��2J]uh���rF�pn���'���h6wx붷�6y�!jF�LE�I �}��
�6��εX~<8�r�I�zU!�C����`���GP��E�ƅW����zoԝC���~���u���e�Mi��yd�l��)&e��@$����7��P�;/�c���{p�A�s@��v2�\�B��_
1Z��_hu�  X����C꾬��<O�ʗ���"�6���J�)�� nv, }�:����Z�#|���>�R��}�*)7L����bW����*_Y�%�E��Z�if�����L�}��?�w�s��e���X�o>�P)�L�!��y��X�#��мC��݌q�$�Ā��� �2�$�R;ÄLR�`�^qN����s��(����շ�eȺMC1b@ن���ꨙ4l��D�.��T�
���������b��)	�(�,�p?��hB�� �B�}��%	SR���<~�A��j�"��n�����iɫ���{3�����K{����&�~��ٌ:�:֠֍(�������V�퇥��`�tל3�d�K�J	�#��8~�� �_
?]M���(;b�o�0H���:���ʻ�lik�}8�'��ꫴP4Gm�4C��J�\A��Dx��H��)e�T_(�R'����0�{�~��t3���!	ѳ��#��)�A�Y뾥v.�+���DO.�(��:}����ܾ�>�,-zLp�܉�s/r�cV�pa����kE�v�=�r�u�dv���r�'��aJ���/�����ҁ䀡s�P��I:�'��!@�rG�
w�ۏ����A<vց���~[�y��n�Yu�ow>������>:j�Y���̲*���>]�����K�ˮ��机�սW��nْwb˗��ƵqSl���@X�ǃ3Ti�����@pb�D����<ʵМF� Oj�	=`�C�#��~�L��!���
8v�Š=�F�7���0_T�C�y�ȓJ>!�%q#z�
!Q�1]���`C$���J�Y)e���%�DX��:��li���\>Ρ�y�XٯnGa���	^��q��g��6j��o�>Í��'��z�:�Y��-"�,�݂}������_2z��>c|������+t�4�zs Y�@�վ�>X�8�H�*GcӄD�K��:��E��
 3@Q����^A`F�A����@��@������/��������'iR�7y�D��.fK�^��	+�c�S��?t�6�9=4�yv 0�d%�[Ef]{��<C�ؕY��qZ;���(��B�p�NE��.|K�#e�0ԏ ֛L��Y齏���ƈL^���4d��<ja��\rλM4?J��1�y9r5n�5��`M^�،�o�:�0<v� 33����Oi��DH0���C"B�5�?v�ç��$YE<&T��{ٛG��b9+�޽&��˱.$D(�.����H��x�i�gf���C�lʨ��Y�բE+
{z�Lv�
��f5��ỊԱ@S��4v�����)�R�t,>`�d ���[}�����Y�[��,=�A��}��]���s��=��$�;VɎx6�ǷnA:�v�C���ap��s�9��Q��E�qm�`�o\��l3��G܉�(�bh4Q닶��׫��kg��[���V.Y����Jq�����؋�����μ8s�u���7mq��A��Z����݊w�Ge���@��շ�q�v� ��ۣպ��C��m�g��E� �[-���<���9������� U���c��楱��w�����7wJN��* }��aԄP�|�o�|��?\v�U�,��d�+����,(��!DC���x�>�B�)ȓ�I �K�"USI0KA;~�����|�wU���+��#b�b��H|�Qf�wV�3U�&&CG��ma�Mw9}ܶ�È�(�.��(�nNB��
$����)�ܻ�-(a����(�)��+�^ ��'f���CCKo��0��5\�`�ﵾ7𳊘-H0����,)n3�I� ����^޸�Y\%!�����E2��>�e����E/�Ω@��7�Ck���YD"l�B$j	��0�K�
�N�!ia��9T)#�0�#LY�LF <ޖF��2Z�!������'��Q|�#O�a��4��g��
oٜ>#c㦾�|��k��Ej`����
����nqw5���r#�����~N���|�[6n|#xwA�\�j\u�:����6�/h�u�-��I#ˏ���I��V	��ԏ��b|��1
8N��H���:�S9�ͳꘜ���� ��I^�H�h<�$YC�m��m(�q`l�gH@ҌN���6��#E/H=���3H�E���x��� $r%%ݩ�]�Yn��Ú����T��p[�
}AnbE�:��oY��8@(Ũ�Y>g+C�}~W�.���3��!�F]9a���'��j}�����n�$R����˟��I3%䯕Ӊ׮5X��������,z(�����I��Ľ���u���Z�fz�ޛ��?3d��#P�ݖ�����Y��4��ҏ���z$�(�Kf2���t����)^�Ӝ�	��`�Y�P��?$���:���odh���4�=�^��Τ]*��'9���WҸ��8�T~0���`�m&�|��\�ID�>4vj��.���٫���"�H_%G���{�/}�s�>�j�D���J��`@��أ�P�H�? `hë�E���	.7-}3u�S��ʈb����zs�U�;�ps="���qv7=�:��d�KS���+p0�ў���5����`ц9y&$-�}�� u����~HҚ�^���/��:f43�n����6��!x�E�ZYW\�;��D��n����C2[f9	n00�VF��M��|k	��J�p��=١)v_� p�!�
`��	���s�Rsh@�0bD=�N#���(H�Pz��f�7���u���Y-41�~w��Ϸ~k��j�=��+�'d����6���(����U�D�t�w���׏���!�s��B�SQ����*�����x`��/[S`f����q�ا�j<-=���}�>�զ�L�ʸ�o�U���|�!#݀��7��|M<�V��oz٭�b&�`�Y���uN�ufcd�1u�`��ٗ�A��۷�2�w*!M�}i��|�2�m�b4Jr �;��ko^Ľ:�f��kᗊmX��ޥC�hC�Ow�r�������� �����0��N�0��Ҍ�9[�wX�.=�ÍvH��E}\Q�Fh�K!��}ד2�=ϫ�[��I�uo�v6�hR��n����y$vY0����ZՅ`I�3d�*�;�ưHm_Hvq[c�(���[��VEc��N��-�[��*[/k�<y��u����݇����p��ZNҢ����(+���M��[R��;�,`ScL�A	A,p �oM�4ïd�Dh�.����t�P���0����j.Y��� ev�ƒ++]�[�Hm[1�T�ڜ7E]�7��Iܝ-�7�=�/o�����[�VI�����[f5�j[�ϓ8:�p�S�V��t��$��9w���W�(\��9��ʗ��"Exʚ&p\(:*a�/����k�o><+Y%n;Pڍ���"-{���L<ш��]��"(Z6�vV��ܓ�=�e��r��q�R���u'H�uM@��R$��ܶ �	�ע�V��eMi��6L]fej ��,�����ʭ'%�-������e�J;!B�F4u#KE�F�5;�}�����h����J7!B�-CM�
�m,J�D�h�~�Ψ�[j�Q�
��D�em��(D$J�4F�h�F�s���2[y��^9��(ܔu�%�e��B��0�ܿ�I�o�Q�jC��5����8�Q(F�mDHэJ�Gd(R��m(R����4P��=��F%Zj�r��#mgy�Ui�4F��D���]��&���^��P�r�d(R��M�J�B%F!��\K>��-�%\B��~����e��@�k䴡J(R��m�׮�nB�HP�s�����2�Ke�Y���:�(R�kH��Dh�����H���m(Z�U�f~���h�]KN�bQrPi�B���-(R�K@�߻���o���Bѻ�:�iB��	�R��Bэ�h
)D! ���"�%ZP�ߺ^����1��(Z���fj��h�(PԅjB�(Z7�~��J��A(R�>k��)X���h�F�MZP������k^�}q�&d���Ju=�-=�7�O?�w�c|�^=�l<�g��su-���[�0�2Ʌ�Fe��B��@���-]ʭd(R���m(R�J�(Z=�濎��U�Gd��m[�H�%4���Y
�h�[VѭJ-(��߳4P�
|�ɉB�"P��Umh�B�d��y
�ߵϦ��P��ϯ^��3�捍Tj4~h��˅
Q�H:��1�m(R�����~��G�"bj��!B�-4D�!�J5 #C�󽽳2幒ᙒ,��tm��D��(4u�!�1-(���*%F4D�J?�MҢQ$��f�E��=����P���-4F���ZW.�D�h����Tm��Q�̖5�T@�6���J֠Me�)BѴ���M��}�_�h�J���ZZP����J����B�
�(P1#G�~����_jUZQr)B�޾/��u��h��D��(Z����-�%�s�f�l3���338P�G�+�"P�B�-��Mu��F�(P'ж��߿:�mwR�҄j���bP�i�%
W��/1���G�E�mV����B�-4D�k�W.[A����'���r��h�B��A>$B%Fs^��ƣU���^J�j%F4Dn�"P�[Dj\�J�����hH��#GZ"P��?d�1�%�E�\�J$�
P�;פ�}��L.�e���Fڮ��J��Qm�%
Qr��`��w�'>��~+O��m(Z�@Z����@o�-"B6�iz�K�%�([�v7��(�"P�
A�~��MQġx��([Ah�m@��i�j�(Z6�մ�FO~�f���ڔcDM D�8r�(Z1�%
	E���gr�����^��^�4��e5~' �AY7N�H��YS���EL���FJɃ�S ��٫�� _�sOs�F�T�_Јx��?&��e������J�J�hƈ�J�Gd(Z��IcV�4�iG��_�+.̍�ɖ伽)F�4D��vJ1�5���ġBҢTB%F�k��Q��J;!B���h�Z
D�����#F�#hB�7��������5�Ǫ��3FPVҊ�B��F��&$�� cU�s�^��
B%Ui��@�ڢ }p��5T}�o�M@��V4|�F�� �5U�nϯ$3�w&m�\����n7Z���'Wm�s7[��Iۺ=Svr=1���F�Ӱ�͓�~j�j4�p�J��e��
D�B �1�4cDh���o���/E
P�|���[V�D�j�Q�4[X҄J9!�b�P����vl6�(Z�iB�-��)�}��J�4��R�"Q�����B�B�_��=�'��m(��Q�ܢ4F���3r�J��KJ�LkZ����}����HP�
t��m�)B�/�j�1������O�Ļ���!3�H�v@��ZP��ї(��h���R�&�(�'߷�5F����-VC���߽����BѦ��)[�;!B�-h�B������J'9�-J�R)BѦ��)B��҅�����/tq(R����Q(Z6������D�J�h��Ƃ%���^��D�h����T���,�:r����B��DJPR�HP�G�?q�a��f%�/.�2j��
P�F�#F4D�J9 m*%F�#��%���h�J��$J�r)B�4bP�~H�^^�nm��_�Q��58���ޥi���4u� s�_g�4�8bP�
P�q�%
P���3@y"T��.�j�ҾB%A�-�mյQJ�±�-���j���ܺ�J�~h"F��҅(�
Mh�Dh6Ƣk���/���8�G0��́ԉB�ֈ�"Q�P[��>��Ouz��Y>���J�J�h����h<�D��UCr�$ԬhġJˁhfB���h��д)D���ٛ(R�	����(R�(Z:������ #G��ݚ<J��-��"��۲���w�|��~h�DJ��g�k���D�h�DJ�#U��nQ�DJ���Ҧ��)��3[��*�L��#���^;�J��ەmTh��-��(R�J�BѦ��]���wUv~��4J�B�ֈ���)B�*�4F�U�HQ�M��2��B�w���Tm(_����cT�h�дw�bQ�.����ƈ�)G����B���|���Q�Q~�j�Q�戔n@R��C�F���z�mcU��P�CM�a+M���V��B벂�4��(����'�d�K�;S�!�.�ٕ�,�D�{F��UA�5�9Իv�u��W=��(�V��=J�ڠό�k~�ՈAX�	Ƃ)���R���X�M��k���;��G��z��z�6���9��]�+��zE���Q���������wP�gv��7X�X9F�t�e����Jĸޗ�嶶�v�#�mv���nO\-;���[��髎�v�\"���wΊ���5]QU��=��^�=�M�-��8��h��ZQ�"F�_���vt��+E��9v�\M�c����Z�Hn����I%r�;�n/6��7�E�<wUN�q �\g����;�0�����
P��5��������J� ��iB�i��
d��{�ɪ6�)B%
P���д��3v�YB��h�[Vд)F�~���B�(r��i(R��E�F����Ǝ�D�J"J��k�6���|����}��}�P�X�#^h�@:�(�!B�#E�F�h�Tj~>��4���qJ<���owV4[Dj5Q�戔��!FD>�<�f��nErH#s�{�>(F��F���r�4q�%
b�,7��KF�#F4F�lkz�\��[4P�"�E�/�?�9�����G�(R��@�F5�U�J�~�Y@�f��ת6�-!�P�F�"����0�Ѧ��[�O�~��B�-h�B�#G�(Z>h�B�f�>�9�U�����M^%%Dh����}ww��U�}�����w��j'�h���q�����e�ˉ�`�����(Z6� D�rPq�B��>�����P�D8�%
��h��?:�iB�}%Z�.���DI�[hġJ��7�i��%�m�"P��3E
Q�(�DJ���P���>������~klC-(P-=p�$(R5��ϯTm(]��cQ��-h�H�v@/!mc\N4[F4D�}��l�B�-4D�!�9*\(Z�U:��(D���F�����˙��e�.��Lɰ�ԡJ>��h�%GZ5p�J���O�2�´�-4D�J7;��h�%q����)B6�F�5h�B�jB�%G��~�<J��,J�hڡ�+Hj�ZTJ�&IV�-`�g�k�h�M�r��4u�%
Q�6����#Zj��E��;~�n�����?�BP�Go�t��J;!B�)���܅
P�D��Ѷ���-(�=��s �e�^8L��sE
P�u�%�"P�G�LJ�;p�r�!6��}���Tm�j���V�*�0h��D�P�v����
P�u�4}�wY�E�M�mm���f�hy-(P��КJ�(�
�j�F�"P�B&k,J���~��iB�r��
P�[Ff���Q�P���i�&�-��5V�{?}��>�f
P�|�%�O�[V�A(Z�Th�(��o]���B�(Z2��d�������Nl���*���k}ΰ�#j�j̠b��^��m��'��C�ݻa6�^&�l=L}���r�"P�:ߥ�B�ƈ�)_ˁ�!B�@#mKj؂��Ur���Y�:�+���"b�r���bP�ge�4��J�j�B�y����J���Zj?\���|�.!�iB%�cE�ZF��J?��]�J�=]�~��|�m}>j�ġj�PJ�h��%@�ݕۅ
J�y���n�5<��X�#]j�P�[hZP��-#@1ƍ�F��j��ړ���prdŋ%ᲅ(Z<�R��;���!B�-4D�J(P�M��~��A��A�H�FL��Z�VQq�e���v�Ɖ9�B�������F=mC:%]�S4��f%"6��J�,ّXw�;��]��}��rg������)�``����4D�j �|���f��.���-V��P��*��4�iB�nB D�h߹��Tm(Y;ܠ�(R��M(R���h�Ѷ��D����6�%lB4|����_�ѕ����W�P�G�|�Q��J+�D4�~����I�d-�Ȍ�ǔq(Z:���UmF��˭�4[D@��B �)BѦ��AϽ�j��?k[�e
u4u�&�mV5�JzՇZ4�nB�HV!3�9�(Z/����Q��h��#Dh�|��׼���'�]�i��ҿ!w
�Ac\N'2R�i�D���͔)���-��҅(Ԕg�V�-h�X�B\*Ģ�(Z?f��Tm�jU[E�v�ZQ�O5֋C�P�B���[Dh�h"P��?c.��lo�e�f��Q"h��%�ak
�Aƪ4Z�G�8x��6��(�@�����;�&�o�(F��{u�h�h�D--+��a�@�Th�Dh��6�D�_}��E
t@�t�:щZB%��k�Th�%�)B'� ��h���Q��~2�)B�֌�P��J�~;�O]�}Ͻ��6��(R�7�ڷ@~�����E�D�j��]`�-~j�F!m�n�ZQ�
�h���.K�/$��&e�4�(Z:��58�Ʊ�҅*!ۅ
P�m�:ך���h�B�-h�� �u��AlJ��#[j�P�P�9��������}�s>(Z5�sn��P���ʯ5#Dh�D@��!�P�i<ո���V���fh�J��l�h��J�]e�- ���Q(�
.B��~�߻7GZ�(F��F4>�ZhġJ5f/�5���X�-F�9��==>_����T���0��$4�6��1��׶H�ف�푓��>��}����.�SY�˵����O F�5iiG$(�)B�@̊P��@���~��:�ġm��
�h�5��"� �)Bш��责?�{����o#F&� ��@X��J�h�DJ��C��-�;�4��P����^����>�TcA8�z��ۢ�(� \��=����Їequ0q�g%���Z�ئ(Jd�5cJ>j�г����%p�������ɓ!�&���o)�H��ek���_����{�&��F12!���ջ8O&�S�!
�4űܲ��]�IZ�y��Z�pĩ��[$�
$�����^}��e͢R������x뇚$xAf���0�z�ٚv���d`[��ͦ��p��7�.��8�nS�2������v�M%v\ܗ�ӂ@�#x:e���G����ｙע�u�z��p�>y�7�Q ����%$r�� �)Y:r��<P>
�����TZH�������������7��m�Ö�Tlg�"��2�\;�bW����L1��"�a�ƑVP'���	i�"	4���4�E+�DO�׵��Y�Q�{UX�d (�5�s�A+T�bur}jdMR�A��Wز�d:��GZ��r*1��]�	h}kk���'�a>h�"e(�7m`m���B������W����q�vb����6�j"�a����Æm��!����k��N�	�\A&��[����B��0�Bޮ�@��YU/8VN�$M~f�6�2�� xʥD���`@�@��m� b@�)�SRH(�� �&&aF�?t�Wg�q���,�k���
P��� 1S�%NTi���Ӏ�qD�?P�������7��q)���h#��N_��a�	d�ZY�A��pB�d�_�I�I��1k.AS������Qϳ��qklGa�d ��l���'����)k��Y(�1��"�Y�ic��2�J@b�D�ԭt�M�܍Dҹ_g9�8�P�j
�J�>�x�\s�����T_U��=m�OX�-�罂��?p!�7���^��y��{͆i䵬���ꇍ�5l�T
f��Ҭ�t��Ը�%�[�I�m^[��h�3h�$�tG��L�`�3S��e�$�᱀bX��9넚D�ݓ7���4�~&���O�<0R��C�G�@�Wt�<"�,�@����u�d�f��X,��{}ȡ�-Q��k�:���g�J{jz�H�`���jݥx�/c5��#D�N�V�A"��`��m�}�2+���`=B�E|����uf(H�#	��:�T+��M�aY�M?���?}�C!� �D� ���22
p�+Ĳ0�������Ŝ�b�κ����0P?2^��q�e��N1rA�}�p�v#扠Q�\�a��i�^>�*�-��@���R��l�$"7,%%q��KLim��޽�O6�Er���/:M'Jdi�}B��D�"���Ń�)$	ĉ��gzqK�g�L�,5�_����!?����6~�(�������\T�6�(���0�d
��8R�f\�@@A�e_Q�L������!���zo�~�ȇ�e�/�xk�9}%� $�A�3����¤��(�`���1�;~�B؜��>w���M.z�V�8P� ����=�`�0�ڷ�I�ob�yu1"X�隚E�f+ �]�yWvU���z���kVnv]��
�FU(�}�[jx�k���P-�d�3[涮���=�g�W���n�~o���R���)r�T����h���c���s����p�b�:S��%�\�*�KJ��
��ڥ����Z��f�.�Dz�|�.Zh�=�x�*Ϣ�Ѻ��7;�K����Lqs�[t˱Ʋu�;&;���3��r�s����Og�Tn��1r��,�!	��=n�0v�I��{=�v������nZ��\�]����sǁ�\i�[���ؤ�I�nã7n�{6zTt�Y���I�r�tle���g�࡮gT�+�h���m��o����|�����w�H��:�N'��tѾΉ�/�,v���sه}��:��'�=��W~m��E �Ј}�q� �M��`a�i}���J�+�}h���[�q9h	�O�-��� �&@��D����ؼ'��7LP��&�,^�i����+ĔЧY����]���H�e"�pP�2y�
�	��do\�J?
(3Mt�TZ>ٲd�׮�C	cL�y��	��#Â��	 �6��J?Jș�y-A�✍$P*E!bΟ�� ��h�=U,�_1�[����(�eBbbw�/P;x��pc��O[�q���	�C�㘪BM�u/��	�L6~{�jG�$!(6�NE�� ��H��H�����
,����\��o��On�ݛ��/Ͳ	�+�<¾�C�DQ��w+�~C�Ʌ"�b���>}`o��hD�*%��	n';�U/��gb���s� �{n,{;�=��&٢��߰���n�cߑ�+�Pů�hk@Q��^�pQ�1�:
�KH�gj���%\�C:��#4~dC�iGR�1!�4b�g7bfI"�8E̻�w������B�g��`} �#|�,f��9�:��,er��ft�`�wn#/!8����T?��d�-�f���l�%���0��nu�/�0Hsi߫B0HoB�u����<~U�~��]uN�S���߽�R;.Y ��/�\o��0����+�jXf&D���t��ğ�HLq�8Qg�[����~�ob����� ���e3uf{�8�Ȏ>������d=��6}�l�h�SI�{�旝�x��ED�=��A$����Ȩ]��@�"Oԗ�Ga�/�����N�<G7�(LC7�}-}}����?B�g��;��{4��^�nb��vuX����e�8(�y�^d��/n��+����E���K��Yʴ�L�B�*ꀭ�����C~��?W�� �
l�rY������{n��w��ԑ!杻���H�I$S(��8
,���t����\EN��BN�q#jv�E�疞d=a�>�8�$��QN�Ju����'q�P�7 �"deE(�Y�S]$��2:ɣD��|���K�)H�%[�_f8��K���x�Q�-}D
˯*�S�4��A"�A���p2Ԍ� �&�@!I �Uɽ��U�[��h�.�F�����H{�oG��M�\�<`G��=�7h��L�"�_&�]�&�t�'1��W��x;h�"�+x�p8�RB[�8��?a@�'�*6v�_� 4�,"4�?ZB~��VJz$ ���� ۬.uP�s�<)���7e f�
f�P�Kd�E���nnlůI��,���Z��i��K����H� 4�����=��1�� �!��Mf�J�P e ��%�1H�B�2�JJ@.�Y�l>���P�Fr������о\N}[)�ں�3�Rv\��jR]猻e�?Y$�o)"B�{`d��-�s�B5D�DrT~�"��;��%ad0��fM�N�4�I�39$T���So]�Q�$$SRS���N��nan���b�!D�v�O���\8�IKe�=�o�ò�� ���������B%�2�PA��LQk$�'iûqv��y���s� �8z�{��3�-q)$t��FA$�t�4�Y����F�f���նnݕ�b�$����4Vuҥ�@Y�!l�O�:�����D�Jz��y�-k�S�r���|`EA$m�1�C qL�ER��^��!�L-${��D� ���S�˂�a��{3n�L�1Srm�T�v�`
��G�_��\���R�R'b� ���S2H������O�mm�L��7��눼d���������H�uf0�Ɓ��q��w�����1~�]1���7�Ǭt֗��7����d�&�����RN�0���1�j�8�F����'�?w6��m�#�oۚ؂܊��ɓT����J �^�@�G��w�X�g�{�]�7�j�V�dK��8�/3nr�}{CF^%(����6�C�n�k~�N��ޚR�Ʈ�)1�#)0l�i��Ƙo��F�Dԉ}Da���(��<�up�	��\H0���ws}���H!��EI���N�R�q�,m�>���d�����DB@/������;�W�2��ש��{`ض=��l�]!�\)�阭qP���c�<0�`���"X���q'f6��{�Xq˛��Ig0��M.�\������b~&���A�޲�TP�:��/[0���j_:溛b���K�<蘣�Lp�̹�*"Q'�"w�ƅ������0g�E���`5�����o��l�z"�13�iq	k܅�Y���u�|gex��id
�&��l5	����Ѹ��+�h-�Y/��t�n����&�z�1�4��	�{𴕟���e��ɋ"�@%l�T8�gM�d�!��ܵJH�j �%��F�ICA.��9@+�����9���yeA#8��P��K�$�6RG
��x�~�j�B�@Y���r�`屋��Q��E�YCR��ui~5g��"B�PH���������&���j���n��A������a�z��h^ԥC��%t�dTL�����z[e�"L%#־�mZ�.o�Q"��yp�>��*��F����y[/s�4��(룢=R� ��`�&�"S3�.���iE�w�$�s�:M���{�ڌ�%��@r�z<f��k&��n��t����dU�**h�ζ5F؝zv��ȸ��飀�7u
�BWb! �[���gC ǩ'r��G=_Q?4ۅ�JC�P��.5c�s[P�#w7n.Q��e��B/H(v�an)�)_R?\z������[u.�9Y�0�L~�W�b�Aj�Y�n`�O%���R�;p��`��F���&��e�uhu���Q�DC���uݎ���n�Tݜ3 !��v$��Ŋ7A�f�s-{N�RŹ��{x��[ڸi�y�cl�{�P|reJ�$y�$��zى��.sek6ˆ����4
i��Z
�N$l3���*xkC�:}E2Z��^�Ǭ�ĺ�T��������;�޷�\/��|��3$:�FK�˙�e�I<Gb���{s/i��5�y��f^�Z�.�#y-�;�[�V����h�n�Ec�D���Ѣ�TS�@�j��bh�Qfh����z�#��"����m[��z�^M�ɴY]]��,<i���
B�>�VU���j�pʎ�'.��b�Xi$��57� �gRK�8��XKm���\��ܩ��Z0���q��.���o:@F�r�`��`ǀM�S�3�B˕.,�5�4��Ҏ��cv(��~В�C"e��l��"�m�j��� %��`PeZ�j�1�+U��5�D�=
�*��Z��sfv���HnóѴHt�r݌�c�&�7l3�~zB>��.��Us�k��ה��m��/��b�r!��� �j�9v��G{�s��u]��ԕ��kv�ct�pb���lv6y	�Gv��s�:� wn ��&ws˶���
s[y1�kn�ݞ\���P��/\+ػ3bݫ�7`�퐷f�懈�Sui�,�2Z m���3�ְn���Em��u�0On�{[�Я�ʨ�8��i��x�aʀ�]�:8���L��Xu�1�6{6�ٸm�k,��.�4ڌ��g��'i�=����x�
�kw���ݥ���e.���ӻf.��'\-��+��%J��\�wI�m�8�\������n�3]�c�^����N�u�6��m�W���JdC[u`�:�7'b<m��N�Xmf\�r���n��Mg����;�պ��{v4�a<��:P.{J��خ�j�7X���Ϋ�E{��*vm���v�Ί�gn�X���v]˃g��"�n7,a@��᪭��v��i�W]�}vG������<�;Y�4n��H�vn)�{ho9�P�zŇt\�p��-C��:˜�����}�}�9	u�u�x�m�גf�ӗ�&�s>�I{lH�[��i��c���M�bf����lE�p�q����Ъl������Ӭ��x��x��;[Jz��ݵ��U=�;f����q�Զ��A8Z�ɱ��,�s��xݥn��:�[��yn���{qjza�p:ۦ�]��ݼe��mN��V�7�ۛnq��`j�cG���ë+�GS�8�zz��u;��y�G�yz��j��q5gU�zy鋅��ƣ����a��/8�~����'�2�[�Ǿ�|�l�m����9tE-����e���stOmlX)H;Sۋ��%�U1rs��ۇF�7^ݫn�':��rs�t���Z޴-�/���;���Л������-�YΑԒ�`g�:��{*c�-���k���\�Z�ӌ���s�g��zLx�k��V�r���{le�=v�ח�w��Xe���a���B���dǕ����؛����`�qN]�rk�n��:�������qc�T���`|�x�=����F&v�cImv��76x���l�0�:L�h˹<d�9���x���:�<u�����#�������'ٔ�n<n��m�1�ݝ���݆8-�jcf�6���iHI9��� ����f��
�  �e�+�H�Fa) �I�ߟ`Wh�XCCZ�H=}�����7���(�,��H�믫PZ6;���z<?_��oH40�nF��b�@��@�B�{��15Ud3\����P��ۗ�/`� C� `�}/��l�f������%	�\��=�9�����7�ρ4|�;L%�˃k���x]u���y,q���vh��:QEz�σ�Ʃ]:��.EO�v9�knε�'.-"�jVܒ\�t�l��d��B?!i�PL_V~M3!�	i1� D��>���,�
;��(�N�R6�̏uNW��͒p��@�XG�~�Z��P$��h�����c��kڪ�ĆF/'���PϜ$AQ9����ʵ�s.�Jמ��3��'�_1��X$�5Vn�\��sPfI �1��D��Iً,s��t ��*rԑ��B���FM�I�F�Ȃ�9�6L�'T���\NS�#�{	=�y�j,�[a�Gk2��urt�n5p���Қ��h���G�F��$ HB�dms=0O�1ȡ��@P�@�Yt��7gD1D�RT �jg��*+�a������l�:�;�(����&�w�x1��,����>$��'ˊ4`h~��T]�>�g35]���VU����]w��9݉|���l*�u�3n�6��U�6l ۹�Î�)��u��y]G�ډzXyw?8��~����M��Z} _��*���S 	
OV���'J/�{R�����)&�𭰳���d�I0QZ:�&h����b/'"�T��<��>���VN�zc~���噷�����X�t��ޝ���#Ie�
$�VGc�[1an(�M���]�L�dA#��U�%/��C�>@Ѫ�z�ϴ�?ae��1���P��?�6QE�ǟ�t����C��F0�zĲ �&�S^etH!1��)Hh^$�մ�?Et��m H$��g����U<3tM��\P���İ���*�t*dWW/}�V� �� P��O�nf�C��!�����n?n!E8�+"�P3��^C�+n8�ݴ��F+������h�u��'J8�pmCk����=�vH�D��d�$1
���?"�`����H���}�e*�a���[��W���q�E��$�m����͎��"Q�I�"�}�ϛi����ɓ31��Ey���y˵��x�nZydF��a�h���$�G���X8I�A�D�w`��$���4$l��^�@�?�1�"��umE�q#��)��'A�E7�'����D6�һ�K�Q�(H$����V@C�^��h������/͖1]���R�J��Ǌ�g;�-FZ}��,/tVjs3
�EΗ��"��9�}ɲ&�r[q#�z�vu��7��-R��RÍ n8!4���3�:�kH��or����>���ahG�����>���b�pW$-"���=���|�;m>m�{�y&�Ut.�=��r�P<D�{Z�JQ���������N۱}����v�~�� �@�N@A=�+4�����f�˳�O���s~M��d�bDI$o~s]�n���]Ů}x��g�Z^l ��
�HT�����t뎗'�<ny���_n�5�ͻ�A�V�T�@ �O�Ն,B3"�=�M\<�@o�hx��C;��9��^����S6����A����,�e ��p�Z{����"��f�td#���}��AIH��MI�Y���4,b�����s��~%�H���wP�L4a�s����i� �Ze �]?+�۞�U�{VV�"�Ԉ8�B�=�BAP5**��������'�$�$�d$�l��g�T�*�C.�9ߘ�J��>A/\��f+<a6��a�G��1Gj�,��"L�W֋
A
%	�ذmtB����P������2��r��E0��N�z����D��1}�\`��<�H܏a;R�D_��;z��w�9;���!*꟧���7@O�Q�x��4���w�lP��t�1�=*��L���D�<��%}�0� �H�#l�d}o�H�R6#q���<�I0�\AD��q�������-l�u�=��݉�ZF�ֶ}��k��jM��B"}"�E��W#�g�f�p�����ѣI�L[������3}�-�Z���0n��Ĵ�h5����k�ݻ�"&9㐩�<�����M	J�R2����$�m�M�A$޾u���oZ#�&�߯+�Ԝ�HI54���t)pU׊X�xx~K�b��߮���!b�DE�������b�p����;���oa�������5D�$:���;Q�����񲐶�U�]�J� ���A�����b��Ƅ$Hۘ"��e��� ��1P�V.=�ဓ�z`2D�i�q)$t�T��TH�C���U�@)�Iu�=9�:E��,�ƪK��=�ځ#ͲL��j�<[ֈ���@���!��C$jFi|]o��$�D��$*Ic?��0�g���ɻ敒'�|�����;64�B�v͊�0��*��*ip����b���t���Ż�~�6{�gn��������ۂ�����S��j����&�.N@�����ko}1�-Dw/K���oWUB(��@D�QTX"uvM��
m�Nv&�����]S��LT�D�7��G�����Q��|����E��3����/�g���N�䬽j4كU�m঍drc��L�S��&l;�,�~���"�"bFQ��ln��c{<\jEI.$5h{^�k��yK:�/� �����C�<=����Ʈ��CEf���vR�c^������ϣp;����+�^�q\)��k��t5F8eƹ�E��5�HxѺ��;�<�u��_�:���h�/]�W�̱pn�R�a�Z�=�)�����Xն�ٷ]��f�;�>s��^u��(��fH����o9�ul��ci�v۪�G;Uk�ųV�٣���;H��YV 1��;��o�_����D�D���H:Q�gy���Y���H��H�(� �i׻�՝�{^�����D�H��(�]g����x�$Q��)#�Z��-9���X" X�趚NH� -{ɡBU�H��cWڕ�ɻ�����#�i8�A+ݜj��O�RFA���h�͟�_m�k�����T�$B�h`��n"�J��YE q�!f�";����Ҽv��X˕��צ�������=��[����y���֭ȭ*q�u6���w���t���v�C0�<(y�N�:_�G��!�{����}�Y��(��ءx��4��a�QD�]�\�M��;�H�ܪ �E|4��Ď���V��yo��B��#ϐ�3� �I�$�k��~���U5.��b=�Rs���zs	�Wu�� "���A]�~Ĭ���r�5����Fײ'	�=��Q=-`(K~�|AF�о�t!F�-*Pwg�7/��z�s;�����ә\콹�J�9�a�eŲ�{<�[���u�on�Re>��4e��GJ4C�S�h�__@ڳB���k���^rj�^S���A@*��EZ�d��0�`,�vr��M�0!?�T��O��6@����?ǧ�N{�X����Σ+>&���6�q�vˇ�C�lSW�筸����=�k5�cQXj�)�-�Vcٹu����?&�+:�ݛZ5D`!R�t�H'J V!5�ګr����ΔP��ǝ!*�2���(i#�.�/�CQ l1	I�gܠ�>l0~%�X�LUiac�w�0Q�"s��擬TGSݘh�E�� ���b��n]��_Q-""���]>[�ad8 ��q��.zx� Ȓq����g	Ċ G*�Fe�ā��YLF���Fa�03Q,��a�o��	b恥O���B�,����,�L�?z�a}�k�T3�&� ��EI#��u�!RD	BBT�8,H�5J��*��ɰ>�� �n߇��u{u�i2T1V{�f�;�.*���G�'�� a
IR���]\���>b �rta��.���=29��:��g����Ц�ؘw��-u���/c2߾Q^˸7.�m�Wr�\�C﷿Ml}۴�#]��K��S�Ap�>��W� ��0��2&Aw]��R�����[H�U	=�(P�30�7#w��/!.Ey�j��.��t/W�$�R ���Y&���G��N1u5d'�o٣m4�Øap�*,�g?r��+�;���]����ON7��
:aܻE'c�g�q��a��d�����a$�%�����R�]�cs������{]J&�8���5�!��SE�Ȼ҆���P�#���w*c�V5q���ց׃�03�3if���x�YƊgL�T���2t+�]7n�s����ӛ���qWp��^H�_Q}�Ư�ҿ$~&�����@���bq�g�t��%
=�浮��t�~���b���2�V��:ؗ�>�g�&ȣ�B9 |�q���i}R9�һ�s�0�#�U{�_$RD�F �@��[���q��HH�rP�A<ӤվB�\okḷ�?e+ 8w;�k�}�6��j���4�hJ�a��ݎ
:Q$d_"��}O���|�M ��h"X"�9�O,� � п���91� $sg��m�e�<H/�G�y`.��g�vU�q;��`m���[��3���7ȏu���4�B��4%g�[�腝O#& �)�KM�OW>u`�����`��Aҁ2^WЌ�1�DLb��w�K�����Y��2��א� �`� ����T̃'���gxx�̄�3��tk�#8�������(��P$ZDf�*$~��b��ԉ;�Oŭ��Q�^zx��h��ps�KNB/���?��O�F�5�s�� B(ޠ��`[���`��(�,�<:����C<1��1�볝����	�u�rFm3��}�𳀔V�)Q	��vGF$
$q�x�8�i�ZF�=6sP�E��A��L��T��=��g!S�Z*MhR j��"��"|A����Nq�=�Xx��	CKc�Cud��j�'M�[��$w���ק��H�i^���w'j����E��I��j���u��&ebo�pPU�T-��q&lф��� 0k�߫��PM,,��$
 �Os<f��Z �� {\���Y0��=ת�Xr��lĹ-'��w�|��1Ws��$��~.fp�|�2�
6�B�A�O���C�,���s捡�v�y��F���Wn�3κ�Щ"����N!���I���8������@ b��0Ѯ��	���''�u/4R�E��Lu�7��D�il�B$��3ƞ,Wk���$8P|��J��l�A������ ���b}�׳~��S/�$�^�$�
<a]��`���@��M{ӰP�0'�ā �I w݈�*���vi]O�$ E{�2�fcyLsr��m�t��bE�L�{��H:w g@���ӕUJ��*�d#
5�Kñ>�pd�I�zBu�Qo��'�����~�}x�Q��'I�WЄ�.5��d��5(xy5}S��:��u
vV�P�̟{ً����Z]�w�NJd>�z�$K	!Z6��&�r����"F�!C��o�l�0(�r�oh����j#��/����x�$Hi$�K��U�mW�9�����$j�Uq�H9HC�������0R3��K1h�G�^g�,ɨ@;�6��+=[�"S�^�ڂ4֫*uf!���"�T����v�d��w�z��Mr�o<�O:r�;^��j���c�gg�����P'�Uv"�wd�=�ћ��1����O;P����qu�[����ܥ�U�螧7l:��V<j9<�������.y����ݷ��vDD�8,��c�h�ew����lu;6�}����;��q���N�B�����!C���v8t�v���5�ݠ�e�n Í����o�<�����h3ۏ<O���n��`ݻs� �{=�C�L88n4���l�sǞ]��8{3VǗ��%Ws۸4ہ�{V&G�$Q_/fu��5<�m�t.���E"a��-AO�d�x�:P$n�L��V�\�f�n4�RCJ�e_>��;�H��q-�>�a�[��\��e��y�$^5�^�y;��DVx�6�$j2bG�x;׹��4ʏɔ�jE}�sJkp��kL �bSd��j��c5͸��7S~%���f�W��G3���DZ�XE���{����'���N��r�$La�M<+��ݨp�����6�����	"%&�'&}�1��Yr���^�"h�yv�)�B6����Q��<����UI�Ο���$��D� ˷F?g�[h��Y�{�ށ��u$`��o��!����@��v�H&�@ "�'��b�2䍸��Q@D��LH��ҝ�����;kb�7�1+��s�{滱�D��`�u�5i�(��w�����k$��"����H�ZXW��Jj��	�N_OO
�ݡ#�R�4�+d�� b�K�{w`9�ێρs�,gvӍ�t�DXƸ��O�߭�/#"�'���ZN<�̆�u�d���Y$Z"c���@�M-i����Yv��kQ���QRh)�]*�J�LF�=�%��;a���x$�.�ͫ�}8�C�LTL��c~�h��8����l{�9��lQC;�J�dJD��:���x�3Ka���� �'}���K�*�Az�5F��-l��S_Hd�����O��?��$V�?��:��d��a�
��@�~�Q&��jںލ�Wt�C���-@Q�8��5��GN�,D�KrFLv���8�b+K|��9D��6��", &]4�n˖׻g����"m��ɴ�������r���� (�A}~�S��`����JO�MH&jD�a��L#�������D!�=���e	O��fN��	��b��W�r�=����7}�a1�s��q���߲μ������!��4��0�$nK�~ �l�!�%ڷ#W߽��H��:ιK�AH"�g��Iç�+������w϶�Wֺd̍ [>(	��ۙW>���u`Ht�$�1�A��l:c���߀薻�;,�ym
��>vI��c=���]h�8�7d���ҵ?�l��q@�N1�<�Q6P\|�"���YqbO+]?{z�s[�d�nq�be�l�kݝ,&��W��(�,��#~�؜NrA1�������%�E�"�Ibd�L$��Lur̤j�8{����G�~߀�	4���s��"�1M/��&���ś) i<��H�c�L�B���X=�򙄐@E�F�9"$�(�s�jH� sq����OЏSk��e�W�&�B����d��+k��T*��t�N��^�2�|�:F�$��:�k��<�+Z��ʌ�`�m�p����)�w�ە�ۅ�����noҞ��p%`�^�X7��R��%��;�A��N�����W��N�l�Kzf�����&�bw�k�HU�&8��nu����iݮ,Xi��#� h`h��{bD����Bxk��B��B֚��WY�쭨^��1cs]�N-Z�3�n}[�����7�)��)kn��Ɍ�Y6�輫�5��2��.X�E��;v�V�n#*;���k]��.�V����\�:�mm���OT��R-�r��ώ�v��w0e�;ԯ+�}%��� [5vUC$����6)!������R�yic����yСp���Q6��*��\]k��1��:̋_v�9�]��[3�]o��ۻ]׸�N+oj��g$�{�%�6�i���'u�T��dS�h��}�խU��������u�yi��JfVv�S&��[����g4���Y1�2�c*Pؗ�/����a�֦������k�С�k\c�0n�r��a�W���::��Q w{b[
T��쮿��f�뱭������o��r�%N�gn�p�ly'1q��^��QwBv`�|C��o*LԀ�HDh�n�
���-����{��R���
���0-+7�^f�GWu��#E����c�⹽�J���mӗ��H���*]`��8�� ��pE�Rm��1��k�We�\�d��$u�IR�L(2^����A܄�|YW?�;�Q~�A�vY�a�dJ!D2A]LK^��4�-!EVu���뱚#*��r}`!!B �s#@�#���N?��W����jw.֚{~�پB9"����>�ܮO�wKj����@��阃5�N���6���X�/~�y4(�=�U�w�fC�3۽�ʶ�"�`���	h7ְ�mgѷe��ծ,�]��mr�ۦ㶥m�q&�l:��%Ҷ���~�s��r��InHfm�{ه:�J_Hi1no>�`�i�I��Q�����y���5������&��7gЏ���{��Dl��(�m�śĢ��D����R���w���4�2�pU�ם��\�2WT�B��~u��C!��4�"��It�����磈҉�]�m�0$���"-��U��ʘ���1Ae6��ޘO�o�lз�0Y�۵X_J_�Y2�ǻ�g7�F�V�+�]ΜVB �I�-�f�W���$""э$K��V��	/�.���+�'�=��k��>w��C�|�4�1��oٜMw��5�5�������l�H�8��F����)�\_�:ًV˳V�K�O%!{�.����qi��yev\�i�D��'L���k^3��<��3��˗��'�x�m�lj�h�)G�� �'��JA���!�zyqu"��s��ٙ�%���T�Z&'1�st�p;��������;���:��zW_�"�l_^�'��D����+�Ƈ�+���?�q��QqjK7i��lg�tj�E�mǮv2� �&�6����'Ok�$�H��Y@GĤ�#��t�����!S�:���Wi�b��Oyv7��Cޮ��f3�w$�T�F����Τ h�l�35'�e��"�M|�PxR4�P%�5V~&�d�lD�%�vv��y�_6���{�t�Թ �|k����R4`-�~D�E�Y]%t��Dm���l�ﯥ&�D�G_�P͠h�xHԈ�v�d2���b�JH<s�T�K�m)�}��;7�R4��t�q�V�`� �s_;��R@@���6<`flM94�1Þ��2��Qq���S\�a(R��EHh^ M�7d���W1��"��>�^��Yc���.] ������<�1?sfT�D٣q�H�=�0������<o6�S7�"�l�	�!�{w.+r�����̽(��)�QZR*��҅�"�D=H�"���jk۰{�y$���٭��40E�uT!uI���HI����5^���w�CYCY�ձ2������tU��r� ��KwT.��,F��� ����e�o[��$��\:���v��*��Yo2�}�n()�a�"]�SK�S�@�uu��9x���ț�;k�i�u�����kW�uum�(K=R�v�N��sZS�:��ƃr�󧶐��L6��N����.���7Zݎ9���K��q�(�j���;C����&0X۵o�me��g��lt��]���:�-ظ7Y��)�$[u�}�tr۶H�i�pb��Y�Vli�iy�x�<`�X�(h�WnM׎џmպ&�ě�5΢$�e�K0��-��I���]-��������Cf�o��8���/��;dQ}f�^�ҝܔ�E�Fu�Y�g�����:�|V� 
z;� 2Bi\	����_Y����dF�P��M��X��k2K���\$.Anw��J����n��s@@�@�{�)@�q��J�ϊ$��.U��cA�D�Qg}�Aha�؊�̱�U�֚r�O�0�p�o���h�-�����{/�nEZG��̆���w��C�h�ѻ�iM$l���$H����%v��oz�9� �l�rw�"���m�S.I(�p���M{#C��Im����w�\~��H�A©��Ψ4�\�g�JGvV
�iA$Q���\<
�CsE"���"7<��,�!1�$$�E�>��]�L���Ch�Iw"X1cW:��ꮮ�bN�V ɢ��A�n�����N�j���nA3�o�x�0�u�I	��"r�i�ys�}��㏤z��7����'��ˇu���wkq[+��s͙��vGr����u�v*}��XXIb�Ҫ_*���vN#i���]`�rK׾��s}��iG���X*��P5��e�pH�"��������ܔu"m�@�J��:�B\�0��PD�40�G��H���,�N'��gV��Ã���4[	g|hK� �g��j�fk�cD�
�u8����\цl�q�h��]2Q�-��j��(
��Y�i�M^��j����g�/+��$m�޳B���x�I��7��w^>sr}ur� ��"��@�0�3�b@cN20���(|qCEm��Y�h�0/�M��}hQ]ꠕ�ʟ��Z�\冼Ǣh��f��������߾�\��'$b�`��t����0�f�nK�A�Z�����ǩ�ڕ����Ȫg!���MH��dl�bF��"�)��;ޯs�W�#�_B  �ň��OP@�)׍�2f&�^I�1��K���O��N�ɿ�L�FVB$�k�%��z��������F���^�t�{��PP�J��_1XJGA�����/���I�t�=h�I&XQ$$��`:�]���ܛ��V����jrX㗰�ٷ9��Ba�x\���Ǿ�W!)r2g�/t���8����٬.̾v/�TdFLH'
�hy��ֺ��͹�D\B"z����/�T�$�{7֘ODi������6�L!�}�ǁ�� ӆ���A�.bO�����LB� ���ݙB����c
4��E�����ViSR?N�XI !Hc����TCkvD��_='ΓN(�]I>ϼ��'�"X���#"k��"̚c�63�pȮ���F�2�a���\V��wzJ��`��M�zqG�:S���Qjs�2��Ue��C�������i�IAH�h����j����lA�#f^Y��|,��)n?��O*LH�F�(%ط&�J�\��h��$HM�cN����{�k!@���
Ť�F���:��
q�b�9��$�J�� H�.�8�?H^�|�ABC��d�X8P&�D
0�a�t�a�YD�!�uf-�9����.*6�30�;؆�ZƑV�(t�y!�^
³_�q�H<�����y��[�w¢�S2�d���$�dx��C��I3j�-;zvL�Ŕκ}��r�pr͉b������ٿ?_	D�`�:��yάi�ia������V\P�2<J0�k�Tfap�&���?$]ʱ�O9��ORHth�����n��m��E�2������G;>�4/Y��<���w��cm5�_u�[]��I�JFM\oy��d�Z�$	Ԥ �E�U��d%��˽��i##H+�y��R$��H�i8@Ӏ?o��E�W��8����]T#6{�LW��@��_u;s\K|����+4X$a�I�ۍ����8;n�^I��Z���E��!-H�r�q"�\
���h�y�����?��� �Yf���>�^�8����?g�澤/JI#�!=Ocέ�t�\�Ex��`@UJKTV9��Eº������ϕh�C(���p���p�}(�!����?Ƽ��t������r�f�h�w�v��Ă'q�����\�
���j�o30��AS�*O��R�+���銱`@s���9V�N+u�Q&ȳ�:Q$=A�]`����E��V� �why�jH�	Pi�l�H�a�=��>&�m��P�"%'
-��V�i��t+��6�A���t]y�&��lh�ڡ`E�$�����:l�M�E3�3�i�{�i�!ۍzD��ַz��%m-�3˺0����F�);ģ��tA�dԽ�tl�$�Q+f�I.�A�0�R/�=kջPI�^�U��G����޽8Q ��2��x!G�_��0�4�,d�j�2_�9��	p�M�L m�0�y�XF���c]Q֌���Ʃ�~�~r��m��^�H(�H�F���H���Cx!������H5h�4v Nn�f�8�k�!5� ��7�W���W E�D���K~�3������#��Vn�ſ^��`���N(9���P�S�71ߧ9*C��\�m�����n���ņ( u�b`7�!4����&D�I|G��C�c,��nA_�	c�TJHK�wN=-�� W��T��g.߻�{���(��O᜾����LZp���hade�c�`��e�3X'"w����o�{��Ggf�!�x��Ah�))�ʖ]T9v�̻e�
����1R�5w"�X�@�uU��͈W�I�E��\H[`�)�gG�igv���<��|dnۀ.6�xh��w�.Okp����n-)��?Ƀ��ɧDol��ڛ��v��6��ik��\��X��Y�N�n�)�Fu�[gi���q��l�Y�įZNb�c�<��iۜ7���l�l�{k <�OIҘ랇��8�^��v)M����페�p��{&&:su�w?��ﱙ�;dXq����͹��]���ݥ���d�5�[���`����C�N�6�2f5�䅱_L�$T������e�F� ���gyc�B�,�V;;4U��]u����VoT�g]q������
1$P �U�}�[A�e�m�B��j��GG��xL ����{���P�u~w`��Qԇԅ�}�]q���0�m�;�;�G��&J�ުu��� .D�XFCfI���l�C���m�uag������A��>�Gψ���⷟�5 D�g�l�Z����a#o�z�5��cG;C�{T�n7jᙉ�(i(�CL��uc�x��{�}%��[m)�g�z�����-��I}�%�E��G��f��ek��o��3Wg:�'��d�?Z�D�"Ϡ�6��	Յ�D�`�?��E�Z�B�~DRA�f���Y��<<=m�ZY��,�f}��u��^B4��s����&I��ݠ��v^����^M�@�6�]z���g�Z5����}ɩ���\lj�1mG'6a!�O�ﳩ�61�_���x�����ij���v	K�H��D��B���?p��s�lG.M�2H4 J'�A~��٣|�y�ኵ�:��R{$Ԑ�$P8~�X�4�)�]{� 6B��wp�:�]��껵�j3Ӻ|�ް$n�u�Ŏ�B4q�g ��+.r�]���>,��-
t2o%�L����Z�_Qg,���������7�������G�C�7�T��+�ܣ���
҈�Xw��E�[-D�pU�~�HX�г_����(��Y���$1�/�7r�CZ�o��ށB9}���^�[�S�	�t������C;<7��#�L�"�j&ӇG)^�����f�S�lemwzr������B�{+�)Lw>������9��^��&�!�l�:�S�#(��r �9"(�/��eY/�֫�o����S���OX�tk{'�Dk�R8+�v:`�T��P|o�^L��[�(ر����r��u�^V=�8��;9ᾺK�9Gpd\L�0@��RL�D��t7��U���*�V7u�����b��'w�;\<t�� wۣ2�h���.G��pS����Q��ƾ��VPтFdµ�K��U7P��w�ET��z"3�=Gu�L�&8QZ:c�Q���Y�����GWv�����PDrA�v۟fA���V�G�G>��{oy�v;�˨�y5���n&��;'hfeK�����d�݋/6o)mJ>��v�׈�"�x��]�q�0�X�!���q��E���O�@�b��QH��e���'�_k�+��j%�seDQݦ��}ʭh���ʜ�ꘈop}��mx�F+aH!�O��A P�%�-�Q�=�����AV0Dc�ޛ|:{FI]z��%���=�'lRL�#}�\��y[�.,0�Q��|���F��2�T�$�T��z��������@xL�F�;n�b��� ��vS�c��C0�%��]��������^��H�>�T2�,(N�|�.�������f!-s�[(�d�.��S���W��R��2X����/�A.�ꇽ9b]��U֟9GPX��t��F���㔷E�!�E��eDB�&�E�'c6�:�]s��e�a��=�sao���V��MۄԬ"����b<U�ݎ�%�Ď7)]�u�w@w�*�r�-{p�C&�=_R��U,ao.�x~�5w��{�y�D�'��3���m>�@3�����Bټ�T�5�V�}c��f�n7zy]Vc�Aٚ�Z�|�v�W�_CT�?�~��I���$.HՌ+�{��c�.���}��d�ö(�%���͏Oe(+{Ea}�^�c�g����g�/�kE8"�݀�Hsq;�<��d��4Z���WD�/���=��SU��r]�V?������"{ϬVF�����B;,�p���rb��s]\hu�����kW��}!V���e ˄�f8�Q��P"�5����C4-m��r��]z�d��/O�`��Y�w�R��5�՞4��z��^�$U^�9���&���f�k�wdA ��YZ��J[��d�o��į1@�zF���v.or�5!��OH�`B�v��?,"�a�JP��[َ��`E�h��I��[��4W��gҐw�Lf�ȗ��:�~Y�M�Ce��IF���|�Y�\/�����1D* �*E��]�d�{��|��0�:�{���ڙӾ��CH�O�WL��l���c%� �z.i��|ӣc����Q1^�*]7<z�Y���I��Z*dK�cSS����c^�����%���7nb��y���eeMa��4%�ܤ�ի���k6��N�%�wXN�ywZ��� �n*�Pv�fe�эb,CՃ�;�`ږ�:�/�J��5�`(<���9K9Wtpz�gV(�c�+�ݓT))YvE�ă�#uc�5dCC��ঁm�M;���z�5�&6�΄f`� 8r�)��[���u����$"^�7{;Fܽ&��3�S�sp�glI� K0�v���:p��6�V(Ѭ���0���'�wF��������+�� $WkY��݃��EB�Y�B=�M�u�Q�-�CG���^ވ{�R�Y���)���2� ����1oV�����wRj�P.�ԩ�ªij�m��:GS��Ҿ:�tv�-Ӯn<����Gh����O�n�@��x�.����h��w��Wr����͵�@gq�O�8ff��6n�L櫍f6*�����yݏ^lXi�p�񒣺7O �y
�J1����XeE�h�^�TbȆ���b�r���Çp�Lo-L�XF�!QT6m��׉�U�|�V[���K�ن�u��#N���m]�η��l�γ��f�W]:�p��Qr�뗂�]������Mmw.�ڐa�j���u]u��t��&i����Rk7�x��:"��7�B4�>B�^�j�^���,�q��(�JInDZ;$M�cS�����	U:%�����%�-�@r� l��J�萚V	\ԍvQ(����j^��%�|u��ݺz�!�p��U#�\��k��/y�b��e��Iu�=��� 펑ȗ;���p�/;v��Sn��c>:N�r����r�ey�[����v�ۃ�.ݻ)cq�x7N:|��B���q�t��ָ=������f�����s�;�{F�onMU#�T&�dm��<�u�:.�.�F�ף�ݵr����1vv8P6z��+���ݻ[������K#�]�\Gv��^(��n���h����Zb������qG9�m��8�k�'�n{�۴��mx�Þı�S�8+m�}v�s-��!�ۣ���N��#��n3�۰��;\�ד3`9.�υ�ϰp�rY9��Wo@n�ɍp�k�^��xر�������x�#���v��i��	�z�g�ى�C��O&3�X�v��!��Ƴ���ܕ�fzϰr���zѸeh���=����� q�.Y�y���aLn9˛c=/n��5�
���q���A��1�l.�qчwnGn�����8z�S1�&�1�\zx#t����j[���v��\"W�병;c��[�]�{j���a<+�9uv�M��1�3R�dp�������=��pyy�&�m�dغ�cn����w'grۭq�n�v�ݍēS�'����]]����s��[��s�v6*:�����,�83ƍ�+m�k�x��ݛ�n�;�e�uӐ�G�s�/���v6ݴt��68�}�5b��m;���/Y�<r����:R��n��9K��u��n��@�۞0㵎����O�8]]��H��v�m�	S�N�[q[&�ێ�Ѭ�ݻRB;7;�Nv��/��$���41t�.�އ�pcc;��q��<E�m��b����g�nyx��-����y�ҙ1��҄�FN�E�B��q��Ӯr��p���OV9����Ru�Úy�أz�#�G*c�ۙj�l��sgk�=�dݛ�M�'���ܻq�c�l�.�v��3X��X�P�w(�)�dE#'���g^{^^�0Z�*!�ƶ�j��L3��&c�Gn_`n��y9C"���jp��Y�5!�H��u����!�SV6��3�����㍵�ޭνgs��\0<��e�_]s��n�^�c��\1[��N�O��;s���a���ݲnv�������=��vSN�:�vm��;�Gr�ۓ��H�@�"qIȧO`��T?Y��-���=�9r*_t�����	��m�_���F��Q`��R�h凣QG��l�'��������TtN2�]�I�_i��`�C6�F��/��;;p_g����1������d�>�\���ܗ��}�aK�'H�A��$�(�-$�`nj���U�$4B?m��k���c��|��*#�#���5(r����꭭��jPfq�>�X���S�(������h�w�cwT���>����W�i�Uc�;ZԠ�)
��)���[tR������
���'fW<(3��z^���K[�j*�U�.Ѭ��Z�g��8<U�%Ċn"�M%Z���;�7dJ�\)f��g<��\eݮy�t�m=��Bb,8N@A����w/�tӔN�S�5b3����Ý��sybY�Q�^��md7׳.���F�g��H�EE#��Ӈ>��^*a���^V�c�0S��%,� �P�i�]�C^��D�c��Qu�|*t�Yy�pom��c�Ō��]����T�δ����G�&}7x�7X�=�z6�������ͮX^����&_��6(QQQA
bGx���DQO���3���1�|��f���ӗ��݈�7x�$aq7�ϫAͤO����\K!A�������vř���cnS+�j&�Lha4��W�d�n����D�4I�����w??w��L���CC��=�Za�B�H�qG%$�8`��vp����R��,B5p-�ʽU6 G�_h�Q���]���Դ���~Hn,?���đ�g����:����k�59z��=�u�\ek����-�|8����FԒSI[����{x�7Ƈ�"WK�wD�kP��7��W���wE�md�Ӹe3��3ܵ4Mm�dh�)8�1r�rmwW�e�Yt5�t*t,.�!~���gU.�gn{�zb'��-�۫���]��B3oʑd����P��;�U�A���36=��$�mg����Y�ż�	�
L��9���kd�F�m���C���q'���(h\���u���+w�]�q�~:�Dc$��mkҲ`�	��N���ȧ���P�0�E�r8/:X����"�fY;�ۛSz�3s,1�5�����-����GA�Krk�W:�Y��Cb��YȇH� ��i�(i�
^wܫ|r(�mq�1_X�޴ʳ]钛8b84��D�u�@������Ēx��FD'�

!;�0��#�}����j�g&T����Y�	��v�:q�T
*T,G#�����q���+}=tݾ�ϴ��f����si�g�����J�UyC�`����f h�%"��3a��^
�}�D���o�@G>'���V �g�>}9��X]0���]�(�Q�|/x�0AAH8S���M8c� [�ɘ3m�%/:�1"k���W��0��΁hy�˼+M����Ļ���f]a�/x�L��@AN:��dHi��y7�w3��[22k��p�Z&��-���l�"�����MK���[�z������sirN��=7wr�4]�-,���[��ڳ�]����b�]׶�4���?m^c5Ԥ���m�\$۲�Q��ᚫm(4kw<t��0IL(Wڗqp.[�ۣi�y��B΄	��
����XI�����َ$1,�"�1��ڝ�չ,�0 pkz�:�s�[4囁�Y�zm���M��qt�U�}3c�˺�g�m��]��4��r�8�z=��{��X�!~��毊��$_�'e6�!�
�7�WV��"	jpb4�э��d���z瑭�+��B�?##��/	��X[}��_r~��$ß3P Ԃ���:�t�`<;����~ZA����S
���P�m.�s�ciU�d��2)�$x0V,������X���^����G�����u�[��d���^�u�f�㿁8!\�s�C�dIц�-82��ln��_g�P�5�'�)�㦩��Q�!�\�\�a�bB���e����"�+���}��ǳ�S7�wJ�R���;ȷ�@m%x{sM�qÙ}&�����u	�6V�wكf�'���b�j#��	��&��펫��R�%�s C�F��Yc770;�\p	�`�C��l`�l����Y�r�sTv��Ѹ�ٽrɻEq�@c�y�q�#>���<!�-��u�9ڭzy�;`C�������Z���Cl����,�k���r��6�e��W(������m4�)�u����]����r.��7*�9������ݳ�;�:�
��ڌVs�����9즻/b:����{r�GQ����N��
j6�R5"rp�xv��Z���V]B,���]H��)��!O��T����E��|Q��#�pp?t�2|��M��L@�-�~R�P�48�E�V�~,�<ז�qx�L������2�v\s�QV�z��Gߌ��/6�8 n�eE!NOu�cE"Q��V�T׽�h͈g�	x/�O����aǜ�>�p���z��sO�eⱁ@Q8�A&�H�g�\��9���!��;�W�_`s=�Ӧ��Y�pfִ���{���$?Dk�x-���|oU�\KX���l�#��s�Eu@���Zd�%�Ǧ�o�9y/Q�Vw��<���ύ����k�db�d��[<�Mu3����Ȅ�R$$m 
(�t��=d3;�9M���ϫ\I���m���N�9񮹅P�3��Z���<>�ds].ĩ�@�$���w�z�wq��q���´S�~M��5���UP�BC�H���yW}.����cٰ�.��ѻCΘ̥՚�f�w,g�Q8�a�
����'�3��.m�4M�Hۓ�Զ���);"(Gr��@,ۆMvKѺx.f{��"���ꌙ���A"R2U�U�{i��[t��J�̊�{z���<I�1뤱�v?r�HV]��苍5�8��G'�L
�r�1�W�����t,xx��'�puV��O��Qb��?k���o�C��~����\��,�QCޥ�$�P���M�ʏ�k����2Z�Y�3�/r��!ϝkK�}�<��0a[����6�3�K;m!ޱ�m�Q� 2$�E�c���m����ٮ$W���; �Gn�����u���p�Di8*G���ﯱVH`��q���:����]FF�՝~�ԛ�W%t�]��t|�_k��ObHE �H	)�4�����g�~���Z���)�U�VQh?���i�@G���#o��/AN�"��u9Wc�B�FT�z�T��N�B�_)9H�q{\^�*��;��2*�� �b�J��R��P�6�i����{�(�ra��a=�X3s��i��L�bǴ��к��{�]D�yu,�\�so���j�o�9P	P \�2W���5�^9s@������A�v���z�t��y�)�X9X�OS0�:��HHbPE#�)�D��׮��,]\?-�Tip��BI�>^R���M������ :tE=��ye����4�l44��@�q���vu�9ܖ{PQ�l:枙��gm:�:�������L��#{�q|bJ���*���*Lc{�X�-;]���,]�������I���9(B$M\�H��kj ��N�=z�7rH�Ø�!/A]��֬/+�/����3Bu�}���L�\�~��,��U��pN�E(���RKn��o�}�f-鋎�yX�xs��)��Y�7��|絟LMcdD��1��d@�10���9x���ci�>MKΨh{T���c������!���y��4����3�E�ν����4��?�\M�o�t�o����Q:먡�gb��K͙b��C�������I����z+ji�f��籋º�.l.�Gn1�H��3sMg/b�}�5f�L���gk�]C��L;�|v7ˌd��{,_5���G�)�C�t({�d�$��'�0$Hf@q��k0up�M�W'=�jH��غst�mۇ�����B#�ٹ�UC^��� �T�6nX�L�ǥ���[�.��	�ޛvp���\�6x���A�7!�b�0�F����`���z��젲ol��Χ�5�$�jgg���p����륨���_�N��P�$�R=�4\�.�w�2���.�/챁W�:t�^.�}�sxJݦ=ƸI���k�D�����!J@�%��q�FXM}���g���hzCT�^���J&���C"�1-m�s������;���g�d�(፠މ]Ȱ�B��8�U�R���\�t��ͳ�De�~��O����!�3w��Q"�9A��!�_y�V{�g\��ffSB���ޯl��onST�;�_E�{�*�ŷ��9{����U5ׅ��c1�+n��f���іH)/ډ8��&b-�%������y-���;�;<n�m�s��$ۭ]��z6����c����O̼;��G�8��eEx���N�qrC�s�.�=Y{�)s�r��g��GE]s�z�RF�v��m˺q���Mr=�ب�e��0��)�[��䨷"�c���ա�sh}���p��v�s��:�e��>O���o����n�WΪ`c�#�x�[���]�26A�n;�[zz��:z�mu<Fr�&FTl�d��|�7ˠX}+�;Ng!��O+aF��NK�ڟA�:zGbF-��{6a��z���Wh16���!����_�
V�u��ߣ��9�A���-yOQ2H�^ҧ�����@־�/�E�N��ӵ�(P�w�b`�JQ7�����ePCӲg�c5� ��W���\%TB��gjm��f21�>��Y���4���S�7	)�NT���,�
���幇��R�~U��<<4�k'�fu*���#Z0��W�ۮ.�ҟ&�6����D"p�P �᳋)����l!�UUyt��2�;���ؘW�-w{��gi#�����l��nQ��e�����Ȃ�{S����mu��;;�nǞ�ݗDg �%�^F�;�����$#���G�<�}%w+N�&���j�b�J|��,>ЧTv֬�SMc͗"��L[�`�D �@Hg-O �İ��FQ�R�fw͜�dP]w�^�s�7�r[wER�z2���*%�wtM��)&6Ws�Im���n�5��Se)���R�G��|�/�� (��{�p.�r�{Ҳ`k�����
]ba`�6	HL�I]2Ɋ�ȪD�DI9�Z8���L���xi��ޯ]��M��-}�/��� @������
7$���D���l�7��zI|��*6���d�~K�朳FqN�tk��WhE�[ꔏ׽yV
��-�HS�n�|ΐ{���G5ig��uRY�yP{|.��0��]�5D�M�_1K����m�Q��H��B�O�l��8�r����d5ŷ=�xvL>22�"�}�0Q�Oi
3�щ���I�K���3����h���g��U"z�W���A9�ڡ���i�۲r�D��!޴�!J6�.(��%庯W5�����X�]����e-�5�����]j�c|���u�Ǣ�аi�iJ��zWZ4(A���F�,��\��w��4?E������n����a��7�bO%�Ss��˝�ak�++74��CJVV��$5�D��lP͋�nN{�t�흩�J�Xi\9�*݁��/:�R�LeBv�$+�Z�m�pK-�y��X�ޕ�)���7�([Eo�|��JVt���<rD���K86�f]N��[Y��N.Cw�w�+�VfQ�RƂmzEЦwj��4�3W���1�h�C��m]��ih�����u�{����]�,kѶ΁��:1/�u�_�K4L�t�}�
�N�Çz�8���[r�*�+B��I*�0Fי�a�p�4�]�F��Z�h<�����& ͢.���=ܱu�C]��2����x��p���
Γ�:�Z��D����6A1n��*��?o�xb��\uX�E�S�<[�`ي��J���SS���pq	�qe�t70�S;y�ŋݜr�v�6�ʨ���3�X��W!;M���lL�יc��$,���j��mn��w%�%�;ͼ��AVl1����j/�4՛*��7�x�q�����.�B�m[VGM�����[�G6���Cf��Oa��H&���(�'��lP��㛽a	�(��g8�V�j�(A�d5�6��<���&W
5��4�Ɍ剢�ªuJ�uo�-&ڱ��/����	�8u0ڻ;3��{\�����U7p�a�/Ui�9�1��t�B=���+m�=��a7�Sӵ���R��%�n���w���~�	��v���9υY���:�o^�C��#3���O�I!��5����{��渘����L6�R�=+]	:��`����G������Y�U�:�Dq����g�I�T���Vf�GI�Z=W��?�����q3�2�l�ɍ��0�m�;kl9F7;
�'InINC$-��B$.9'm-�n�ҫ�xP��d �nD���t�UJ�
�f}}^Q��������`'��릂�k�5#�Ip[��8�9t����V7�����B�$��x��!��~�Z�Ӕ����c�U��fu���{N}�{�*�HY?V��6��]Qw>�X����]u9b�2�ҕb������U}W|����l�Wc�8,@	��A�:�R?`���g�@��K�����Uz����4͙O�G�9~��4�
�v)b÷�j<��wC�F/z�z��kk������a����8E��Ʒ]���ֶ����y��g�Ye�p���bt8��X�� ���7��ty�����{D`�wJ�J�;Q���s��1r��z��M%]� ����:�����``�"��E����ƍ����Ʒv@�0\c����7]��Էaڷ��P�*�9J�,��>FxvnI�u��p�s��yצ�)�Lƚ�6 ��1�s��dC��}BD\1��f)ݲ#��������o;ȏU�w�R��Z���rW�ʛ%�uȏ��ݛ���:Ͻ��2ZS�e�Zp^�^4	��3:����u�Zӳ5=�'P��|���k^A���&�y�9��ysJT,0��Ɯ��(��E�Fe/_��"']w5�t"F.���@ھ�
\��5dɮ�����}=��ҵ��l��^^mC�q�&BO��/+k�dS�q5�;H5�:����n���c�0�:��vTEe��L!�����������^����R��c[���e�eέ��:j������&3I�����;L�kz���ڒ��r�7�����~����q�8�Ī���0�#��殷�2�'Y�g�����;n9�y��Z���V��8��m���Wk�vyx3\�z�{<�Q��v#�8�M�n+K�'up=d燓glt��R��r��x��
�؋�U��+���/<���nݮ�p�nszjp�m�v�ӮNۘ��54v�Ӟx��JO5>���B;t�Z����.ݜf 2��l�y(Y�k[9��ƳwC�-�:{	]zI��8X:GcʧM�)F\�)�§{ݏEk��������{�W�~����_�C������O�m!=6.��	Id*I+sݨ�������4t�ڂ�ir�k.^=R�x�"��v���ꆊ�^��/�E'�Gn�T�ޓj��ʘ"�}��Q9Vēݵ����x]���j�ںB��@�&L`��ary�T�wmݗf��r!�ƝZ��wpl�;�qW]��?o]������K�Ƒ���F���d̲�(�C�	�W�O��8S�rܱ�g�nzs��Y�4�m����	�}�Gz�ú��k����Lїl]"m��Ÿ�8���!۞s��GJ�;N���:�pL۰��<�)����}���}�(�nL\�?7���C6"q��\�Ů�~]g|���E���,��78��>))B�%%y�L�b9���i�v=�/"v��G�ֻ�mp�)W���lbZb�U����f!�	ӥBSD3�{�Fju������k,���du-Ӧ�e�r��(<&!]����]�s]��H��d��ذ�&�ʅ&$�#̫��;yu��=��+�W�~�ة�E��xbL�����޵���`f�g��*��6�	!��p"T��}�Ĵ����]Z�ݵn_Rm�*5W\U��pY}!.�U������>˃�j��<���OE�_s���J� B�
F�b��{)Ľ|�:6��"3Y�\(�Y�!�]������Z���f����;v��G� $ѿ�]�Ȩm��ب}l2C΢��.b��r��v�m��b��>.A���^⫡��&b���V���v��ԫ4d���\a��pn�Z���m*�( �* ?5 ᾱ�6�Uڝ7���Y��_/��^��*����w��vp����zw;F��]�t�#v����*R7]Ta���_K��!�/&��M`�/i��k���r.n5r����]�sYsD���Q�5W:�u�\���͗Ba����u�.𨆇e����wp��̣��ZI�;���u�|!�{)��|s�"�&ВN�e0�����2�wE[�`Xm:�o�g��ر�_�0|7ubာXz���y�ws�0U����ܙg�����~r�tb=��&ul���tަ��*��Ehm-����v� ����r+�s~upgË�h�Y�Y�6\�'���N���������x%���p�e�l��+J��u��Ի�'�˚��yx'����ػy��u�7�gXC~�ȳ��E1^�AƚQ�A)b�o�W��}S�2	��)u�S�p�o*�X��^��n��ׇ	6���~8m�2-���	�dF�9�q�*��zӾ'3��!y��ˉ�����*eʲ�]��b>�Y$\�k�ǤeC�4D����������_���Oj�XTk��k�0�[��H��6�m�}^�b�%�$�z��Ң��\����+��
��g��r�{5R�ۖ{i|����V��7��F�%ZLS�+mk��<��p0(�B�

���=6pR)�����W��f^�(�q���nd\��ھ�x6n�&��ޏP�^���"F$?Dd(aSݘ�mz���e)kg�u�ln 1ڨ�s1�����_nr�Q��~���*N�#����/���d�@s�������O�ֱ۶Uߝ��I���'��_R���hD���x
ڃ��="�����vƽڕŪ���^G~w	g���?=��?H�c�e�RMT��zX���FeL�ïCN����`X��r:��<�qm��k��q��øY�c��$%%y($��^�s���xvZ�G[�;��19Z{)���U��.�ٺ���i��~?js���/�D�1(M�Yy>��?ar�&�{=Yk6��S�$u�`��e���B�7��x'*0�>�몧�;��u���a#�!Wl�5�X�Gݖ��cf�"�D9euouk���MӖ.�5g&qg�c�/he<bvv��2;��U<�e۬��mr�'g���'��F���m����k�����dl=s�wq��p�nI�cb#MbZ2��cRr���۲�F՛��s�9�q�cv�Q�conγ���V�w���ۙ�Iu�(^w$9����pNݸ��9����������^�J]���hcb���'F��<6ܶ�����:ݎ��Is�9,a�\@��<�@����':�^�k��"C�$�ף���<-ڎSŪ��,�P�9$��t�o���T�O���\5!�̥F��~^����TW������k�2i1@�$� ����|]�
���{�!4��&���]��VԒ,3A�2�^����z@&�V����{��'>`�d3$9v���W�`7xͩ���g�2�ތ	�|��~�'>���v�p����^Jɧq֙,�%B�RM�J�Q��)rI�3��w(�sҰk�j��Z¾ �D�V>�4IU�M,��H8p��T���&9"��/�u`��К�f��^��ׯdmf�'F�W]�������L��*��s�:��dɋ���Ϯ�@9(��K[%S��nnّ�鶼v�I�XU�xN9�2\;\�3v���z��+�>
�̂#v'�1���ڭu��v
�V�5��y�Y�X�~H�b��S߉_���YM���6�f����y�^�j��ȓ36��(�۶EdI_-LpOww ��nhy�V�/�p
T��%���`���-�S�`&�¦�Fˑ��;gIE��ܘ�ưT��	��~�U�M����(��bl8R%]�A	#�U���t��3qU��=��qCJ��R+3v�-�Jkiٕ���$L�TgA��n9m(��_�Mڙ����aS���V�R�ut�������`���+b�冡f��SK"��Ƴhx��m�J)�`/ ��ty¶�_�ą�Ժz�L�������t��2��uj��Z�?"���Sʑ���q�	zM����n�A�]�P�e.-�v�ַS�1N_\���Y�f���Ջ��$D��os��7�+��U/+��WY���U5��LI8��fay(_�!5(�S�`�z�������,.>7���a�G��
W.v]�{�ڽ�<��i}�^O���2Fم��pS������.R��k�ԝ8;=�iWL�؄6e����6�8$��cI�]�\{��0���'Wf ��Gu��y&���[nC���>�+(m�r�!�θ;$����J����bC9x����9���1�o8�"8WwJM��Ț�����^��.�ɢ�qfUF	�{U�q�81��8q�{cD/޹�$��|_#@Y���ֶ5�Xn�o��h����3�\�&�mY���kS �?n�"i퍞p�.��fs�G8`]^n�ݦzE��0�<aw:�cm�g���߽��YB��L}R6Ί���xsZ ��˲~,�oeab����^Tߚzp��ZBҢ��n�laű־��z����tߗ�wU��'1���5�ڤ��n�u@5j����D��������Q2ˁ�H2A��
��r�e�Cmu����@���?n�� �d�[}�o�}N��q��(ѐ��`̛s�������#؅����J�̟�1u�;��:N�?�#=��j�#*i���	ݦw��nX�����{.�l�ٲ���k�� ��VQm�5�)���o3Fi�%�@����:��y=�ܬ3�=��9���,�>0G�^��G��gc��-��nS5rHP���~8o�4|o���\�)���J�tsU�lf/{)+�7P��[t�7�=�-�C�ѻLd�*�ű�'cyN�]�q��&8���Q��%)��K��}���.�Y�Q�BwC��V�3�i>)�k����~]�Y/Ox+<��B�RJ�WIa
�F_s�4v�8�GLԼF�	 	�{�ד��Rȡn�n��-��8��+�����!t&QXL���(㓨�[>��N���F&{�9�[/8�Z�\i�s=o4k�n����	3
m"�p�^�4������z8Rzt'S���q\-K��a��Mԉ�͟i�8�9yw���&�C�Xa!	��̕t���ydש��Ӓ�^K�ȷ���|�,��{��]`\6)߾��H�� 4�W�P��`�Iz�b�ܰ��o2tؘ��d��k�7oH��rƁ�\�Ȟ\6h&�z=I��w�G`d��D�����wN|�z�(��V�w5�9����Iٜ�n�:��f���tƜQ�
cK�06���S3l�[X�d�5^����}��볊T�]$�����B�N&d��{���x��OMJ}�Q����Y1]M���M�Sa�X �o/E>䳻���sN�,��%�S@m���
�x�6��o`����vev���;.�=׆VȲf^� ]S�	���ų�of�3�T/�K���fSV��.�m8D�6�M�	�(�6�6�5���>ֲ����wK���)gQ�������3u��P*c�� Y�V	�ҽ�6�=�1��`������u�|����JK�]�;-���W3���e
��U\�H�c�o���&���y��\��6����nd.%gqa�.��{]�po='��^z�1�y�.�Ȝ�ln�v���r_v�"�6i.�������s��s���u�]2q��ԭ�����l�(�wҚ7���%��Nq��@3�Bn�S3�%ڰ�ɳ3*=x]t��&�M�OfϏY].���v$Z`>��w%��z�%nʜ�
9�ފQL�c){�8�r�=ϛ�A٨t��Xok���u
��g�d���ϩqߜ�X�w#T�k*b_F�#������i��i�nT�YCzNyV���v8��K��%"E���-�vd��j������UZ��`�<UUA�H[5n���cY�l)�����`�'jj��B�����V9��ۇ���o]�������S�C�ƕ��@w�]Y�v������Y9�\��ҫŻ+#�݋t�a��o�u���(:�{��F���k�U�ӌ/����ɷ��s�6��cs������mtu�ާ�b!���f�VnCYQz�9v�g����b���f��=��0k���kn��cF���R��u��Ggih^���n����w��.�a�+�yu��7��\�w>gl��Ƿ=r=s��uC��[��s�-���{O#�Ȧ�p�CnۍՔ{F݆�G��b5Lg8���0��gۓ�=t[��ǭ�mΊ�Y>�v�7O]�����]�<�n5uns�;uۜdu�GfG�$����<�Q ��l2��rm�8
��X�u˩û[q�b�r���X�]�#���(WV.y����rN9"ݸ�s(�#�ܻ��e7��؁�/fç�v�(�%�V5�8r)&��[A��mV磬�v�`��۞�C��6+�'�rq�\�0F���ڴ`N'��605m�ȝ��^�c�]X��gX8��l�1Оd�ezrR�������<���ј��z��u��:Ĝ�Ӹ#���|';Dm�cmc>�݅$�[]�v�(���y��.=���n:�y����6Z��t�h��sws�׸<�s,'p���l�;8��o��sl�*�#�{{Y�[svA7H�v[�uݝ�;�y����j.�L{s�kK�<�n�]����Ϭ���A���۝�rq���NPw��[<�1��.6�z�s���D�ŝ����'����s+Ļ{�m�n`f���Żr���͙�==����c��a�%��;��P�᫞{x����%�,��ɷ�sp��\��7a������u�e`���=���]����vg]�?�s��~�#�
ʦ+v��Z���쒫�8w"��ܜ�f�h,],�՝�J���[7Q��k��qc�z�dx���z���Q�l�̝�]�/^D�.�@	�*��.r�����.��tU�Vdܯ'v�iV�7jsoLq�7[��rnꕘ�ZM���ZWOY2��q�-T��v�d�"�Ş8���b:�������^9�4v�Oo����|R�u������v+=Xx�b����d��u;�{\���u��n���+��m������ҊM���G{u�n��@�޾-��uJ�½�/�+1U��D�\�1P�'���Ԏ��Z��8��k���s�=�W9���Dǻ�Wu��+�-�N�_�-�
�z����\����/�4�Q͇�28=��.�M��C��0��a:�� w*]i����������CۏSt�\�p%%"P�X(5��L[�#��P��`+��6�L=�UT ��1�!N]�����+����]�'c��c�� I/�
Ҙ#��uvydÐ��WP�L�Ъr����-]\��5�k�׃2O������E?��Tu�v���sHļt�nv�v�.�u��m�r�̌�j�Li����AYc�3����w,�����b���+�<��L��Ų��OG+_ّH��[k�$7q#�/ٙx�;5SN��u� "�L��0v�C�ٖMv�Y�b�p�ȊIk�x)���_4�X9R�wlŧTi����R3}��qґR�1s�=��/o:��r�y_E����x_!�o�P�̎!L�.��UxJ|��"�m�Ycn0:{&S)t�y^sr���u��1lU�
�э�@I�
�]���^��W�q#=[�oo��b���Ӻ�qP%�Q��Yu�J���)R+�_h=���N�L�$҉'	�%f@�,���y[�6<��w�i��]�­Ór-�J��N��,�'���q�U���7�s�˴��e�$��b��b�W�ro�8��o3c�s�{{�����7=�J.�ek�$Tl/}�N����qa)�ż�m�}�#˕-����{E�b\P6��>���R��AeI� ��i׵���4a��N��X`0MgQ����$�U��V8���w�����d�V�]��fm�N�k�&�QAm�l.^:�W��A�A��s��3�q��<"ź��<�2�k������h����/�jG��c1ԙFc��/9�ո�efŻI�wn��Y��������J�*�E���&�B�H��n�2`�c��J�8"]��I��B�f{��M��"�Q�ڳDMU���7�"�eA"R�{���H�7ݶpVM���}�&N������/g��gԯ坻`y�f�?՟-��U'����� I&A��a�
��n�#�{v�h�]�,�s�h�����m����rD�ʒ-��:�޾�����#��E��NZ����Q\v��ow:�M�g����Jc����%�%�S�3&R�o�)�Y��2���ɴ8+o�ʼlz����Q8��������>�D���Uѿ�?-౤�������D��a��)l�[oL��΍�^�g��ל�[Õ�.���,�N�zE"&g�l3%��Q�c)��/��ٱ��I�#�)dl�y=�/q����Hu�k)�"�W�brA�<�0�m�
�^5d>C������:�T�*]#�Vn"�b�r�*���z1yPU�����/+>z�b8��fο��1�UI��Hp3��XQ�!�M�2 ����m^p��̛�Q3%1��[(��CN$��2�����亂��BD�1�M����`�dq��8�Iuޚ|e�y�
�`�����$�L6X1���2��S����(7�J[ܮ��elo&*.��(4��Z粰v����(-~?�f�q�*I5̪9�Nџ�g�Xl�<}�����O��,[Y2k3��~|��A���m�TqI��'� \���Y7���UYŁM���������u�g�rgU>�)P��g�kSI��r���A+J�A�^+�;jŻ�wX�|���e�ؠ��<r�}�����29~~Lm{��Z�+~xZ2APF�1H3�g����s�"Ld
L��d�U��7l8�z�&+m�Z�8�j&i��\z�V�� P|��y�ܾ��9D�v�d޹�X�m���ft[�I�-5��2U��c8o���7��:\f�?���c���3�қ
� �g`���	�.
̣�u�.ɭ�<�M�u� ��7hs�7;�ܸ�:m�9���qnhݬ8������k��U���x��Ctu�l�E^�ӱc>��eLlg5m�J�j����������=�����cVg� (��-ܓZ�my�0n�a��C�z�S��<=n� 9�2��zqm;`9�%��v������^srY���.�]�F;<�|�������<�cn��N�g�����j3��ь�$�#�$)B�g[�r��«�瑫��k�h5�m����U�ҵ^!���DAA�\)�Q-��l�#�@��ƨ���yp�{5X��!�"�Ȝ㪟Q.�Zj��j��KM�M�(�4�P�	)��g�;9�����;%��}��s�)7z���0����GX��>��$���9�X�i�}��~�ǾeG�Y
���S6��]�gc�2�G��<^q+Է4P��b��2VȃQ��H��+wq\j}�Q�񍋸�V����ҕ�וE7݊��n�IS�p��w���D^i�7�d�=�c�(;<�˃��r�ӎ;5t�:�4�z�㫶� N�B��ВG`�Ѓ �u!Qg1��uۋ	҇��ku�w����S�$��OVJ"�:�S��ș
A�TL�#���%%-�N��A5��d��fy;�n�dq�/+篵�,��K*����wg48�²1�+�� �����m��J� ����Â�ɷ2s��5mf�bn�����oZ��A��5Ƥ��Ԕ�ڌ̀���닆=�U'1��C�FÞ	c��V��u��<IS��o����T��PHB4��ʽh��b�=��5_�/%�ʦ�,���b�J#Խ��B�{3b��kw�J�V]���ΫM����4���f������w�v�_7wz���V#�SǢ��F�ق�Ep���uB��y�;��<�;�'�j�B쥎pjn��$��n{n�F3�=�����	�7k`�������o]�s���:��ح��9q��k�u=;�{|�n�P}<�YP�LR�L'�GM�͖�E�q�g
�˚@��:7�j�F;�C0�a�n���Um4�^�'�W�V�1�)���
()$�N�z���3el�s޿t�]>޿51�A̷���A^�x��N�VUn��g��E��e%]O;&PfU����4��5�^h�SokO�z����ӽ�5پuW��ۆ��D-�A�Kq�AUnJ�TFUZ�4s.�/x�,8Ĝ�-�sOS��9G����;��\W^-{���hĤ��#����fھ�.�T�s��;j�����;�A�^����J�9g�K=Xw��j
͕-%�!D�N�Ɠp>�<ݝ�����Rv�nSv��V�\��)�Y��9f3g��%	���+h����/�Id�Q�q�����x�8�X�}^�"K�ĳNV��7'��r�E�D.D��;�t
=ӗ�֭�mRi�8�,��)2��N-�K*RQ��u���-b�-�[.ms�j���I	�
AA�c�C��h��7yg��`���G�mܮ�yVdl��k��-�;���i�q݊q��
#��#�յ�^ݮ'}����t���\�)��]�l{ґ�(�;(���Cg^�G7ikJ��cίJT2��v:�h�"��E�-��P��vuZJ�X�e�o���9W115P	n��
p������)dѮ\i�Y��#0'$u����Y/w_*��K�Ջs��i���Q����w6�)|�����s�KT�	o��������8l���N�뫠��\a�ok��m����m��.��Pu�� [ғv(��`��d�N��)�૥@��Gv��ҜS��R�Q(���P��U�n��y_�T��o���P#�Gfz�n�nl�{��86.$��eh��ݘ�n�t��j��+�g-V��/�Co'�P����@ӑ%Q��v�m�5�)��-���|0�N�O�Ӧ)����qa^��w�������m0Ϥ/ AJ>z���FI˦���������K��8��O��k��L{�b{ـ{�]EYrh��Q`�/��H�* ��A !IG4O���'�t�K�h�+���ul�u�멜P�^T��Nr�m��yV�{�0��?o��ե��-�e��i��:xٝ3���r�b���T\82^d�s[{@Dۍt�f&U^�(f,�Gu3JF[J�-���5[�h�3S���Eͻ;���d0sn�;5�;l�wl,nqYp�A �{f��!m���u��v�;�v�.��܎3�� �����m�)�pv�h����|���AǕ78��v�s�ݦ.�1�cF��<��r���q�9��PƤ��ϒu�
�5�N���CXt��q˥�2v.��8��հu���Qm �X)^�@Z��q��K��_�ζ㱄�gus����"n=�������+�0:%��=�.;
ů߿�ͬ�f%��Sn�����K�,��}�N�S]�h�&�cu�5�ϴ��QLH(���]Ρu�dփ�Q���TQΥ�"�*�d�L���wl8��'�R���ˢ<^������|�J�L"�H����T��\���0���6�3��Eʵ�Z�h������˧T$���Tz��$3��1��rL��G���L�]t����޻~����u���d�{�^z�v%�oq�f�t��4y�1|dQ&���ʝ�R��G{�5�.{�x�O8�-��jR��FY-�k�^Q�Y3���%�گ\\�v�ܱ�Sx8��������I&�c>�r�ttu��n�ܠ�:��5�7jJ�u�U���qƲ�MJ9W	{��81.�}�!���N�
]��v��f�-��%d����Iʞf�#ݩ�==�^]Z���iߵ��l�7ȬBwsog z��D�ʖ��U�Bj����nb��Sx��^�ג��bV�.�N ��V���eDӠ�P[�Q�{F�Xa�X]�SY{���yX���0�fM4 �yx=��A%D���T�$�����ىV��O	����~V�J����pȞ�erfoe��G3�V'ol`@��&�H(໔��a�4�T�J�A�Y�v�N�=��ײuf���j�@�ڥ?)ӓ9}/�m��?�J�@�(�f1��K�
��#�o���/|��#�ӵ������=�p.��U������yO���xZ?��0��n��\\mmvj{)ݮ���2�9�r\$��<�#�Zm�
�u�'\��h����Ge!��^;�J��0�Ot����_u�5�6;{�u��}&����,���
�R8��w-����S���k�٭𕙓��&����9�W�t�a��,���C�WX�:7��=}�Ҁ�Ɏ4�N�y{�٫�n؃+b��ȵυ�����X���u9���.m0��|GnV�+Z�[yM��r��(Ǽ��/)�!�k�8/Od[�ײJK.�A�5�-�w*;�W�Ȝ��쳌r����l�]N��iUf�<��=�>�p�&PәE�/C�#��_V�rf2@�.�w=�w���Lx'^b!fLg�����7d*�V%��i4�z7�yiTH�;�;�iD�z�0���$��X���iZB�����M�Do�����
&��m��\�`�)lu���]uk��<��j���� "�[�E-Tӳ.�KvuuH�����r����-TN����pD	�Z�*��$���[�n2�t$�++G�����&)<-hKn���;d��}.wb���|n�ݠ)�2�t����Ⱦ��܀r��dn�	�ū�2��Nr��W�f�v��Հ!�@�^�K/U���XV�ؔ�]V8����1j�%;��W5nŵ��DT�2ɳ���v��ҷEk�ۙ/@zf�h�X�3�����3��u�p����$d^�����
M4�!���ฉ]��b�W7�gQB��lzo^V�4M҃o3gi���YZ�n��5���}X�h����G���3�Pk,�ʗ��>���A��;lni̫0P��G}LJ�4a�A`�r^�f�u2	���b��v��Z�r�?f�s�ݓ��o`1�x����i��;��m
�,0�|����l���l�&�
�6�f*7��>�����{DU�v���z/&�絡�Z��d�Ҿ��	����<�2P�!ܓtV'�7�{�Oe���ą[j�Yу�ˑ�3l�����t{�Ooh[�����]* H��!A$�)��R�=���`(5��ϫ<7yÚo!����ܹt�V�/u���`0ѭ�=��#M!�	����Ÿ��A�����7&���l<ZIa�xv�y�DdH���A�{�i����=�7]��y�w��VV�Z���Y�&�;1x7�u��4�*���"_��2�I˕)(�dU3�`k��c�oZ9S��yK��T���Z�܈����q��	��n�:_\�����䏆jCWs�2�U5��^�B�����s�m�qՇ�ޱEq����jeeW2'E�Ȑ��Q��<���^g
�Wp����b�]83[ߺ�m̭	��o4�p6��Q7�n(:���]�F�v�ǽ���޺ޫU�82��k�ʁ�1����//,-�N�r6j�˵H<���N�4���z�@��R�!����}�C2��<\�6�pܦ�e��N~Ձ�1���=�|�
�]S9|��T��k���!��mȈn݇�c�v�8S�x6�m�8ΐL�Ń���Y��8��+�ʉ�)&��bV���i�����W5JwNԀ���a�=ܰ?uX�?g�M�k���ᄢcP1�}��؝�=�pܯG�6jx8�sE��-oR���g��EOWT�vw��a��:e𮌛���`�N2R�Ly3gt�C�L�t�.��"�Ju��5r�f�O�=��iDS�ˎ#��zswGN39��x��᫨Qi�9��;{�&��OT��{Y��@o:�T��V�+��5;�T����%*٬Ҹ���_k��&E;ݝo��)T��S/c��BZ��8��Yt�c�w��<�^���_r3�6��&�e.�+�����.�]*C �u{��f�Uh�ưG��]՛9�q*��������o/	�ҙ���n��YJW;\t
�*x#��d�|���V�y����e�X��Pݘ�oQ"����8d�����P���81�=���Δc�qO��y�	[�	��Rv�c��Gm��;|}�ܯ�� ��>��q�7>5G1	+=����*���7�UXw===ve7�#n9_m�q� ��.P&�X�{�`�k�r��ۀ��;Ԟ� mO|>~�Ѷ�v���Wufԍ�����-�"�������3�����Ap۷U������>�1���Q�W�|-�Թ��ʮ�{W������~�s�ص�x��K�����c�v#!���	ȫu��U��Ƴ�Wf�;[&9A/\�[+Z�g�����{.Q�x׎��/+*�U��22bq�䝪V���F�nL�����,ţ�5*
(ҏ�P{��x��}��tr<E��N&�H�����`Z1��٭��ܫ�ɠj���g��Ż�n�ls���:zޓk�����nD[F3�!���1�7ܳ/$+��%�7�`���Ksuo�Ѯ�1�T�iJD�2�6����2I&B��"a-@�2ܶ餺6{���F��q��𥵀�t�ێ�^`�~�9/K�I�},e.��}cf��0�'�\�%�6pR������.P1�|��#2"c�^*�>���
��C�� ����n���P%�S�"ry˕�
������%��Y�c�}�n�GF��)���V[Y�v�Xy��:�>�qУk�-?!sc�O'W��Q�Mfdeh�)����R��9�mC��D�R�^��j,W}���+*�����ܱ����t�;����p�칮>+����m#�NI3^��"�A����{A�1o(����>؝]���6�H����I��|\��Kp��"��+©]�X�ߺOcvEFMOe÷���V���<��EnU��!�3:٤�i��4�I�T7����U�A��:t���*�N!*ŭnӪ��A�Cҝ���sU��ߨݿ�݃&d<���ͣܭ���#N��=����ڦS���$��Mp"d�p�48���<ݮ�@�[�ݜ�ڵ���pZW*�m�[�&�l�`�C��v�	6���������{=x�>*Rήh�2�+k���:k/I�sk۴w4���X�ŀ2����C"�J�/:����٪\9��7y�kh'��kN�]�ˑj��B�t!�׸X�V��a�c�׼�$�Bdj2KrV��t�幙��V��v��=qD�����������(U��O�z�.� s��9�$$&R�����ˀ)S���+ȋ�]��F�^.���z4{�����;:U�=5�X�p����AqJB��ywOD��=u�N��=�yx�p�r�ogf�cw���@S��"��ӷ�F��q�̓f�<���8V�X�qHFf!�{L��2]͚�v��u����b1�o��p�%�.�����k;Ź[$V͘���k�m���m}�\��QS���1y��J�;X���%����v� �#iZ٣Gn.���)�h�Hf�:�%�s�Ut�b+oE�|'ZIhn#RH�N:����ɼi
�7ۻ~6��2,�gmqˬ];\8������+�z1����RR�f�n�{�H2SV�������n�w�����k����aNFmҫ5��5;�H[���CS(G��}Q�JF��'���i�w� �R_B�L3r�d�m�����=�����qϻ���{�p����������N}v��+r;�q��wM �yG�vk�g8�d�ι��ȼtP癅(�D��P�dN��LH��co�^A���5���9Ӑm��lW�TP�F򛸼�A�$J�}�f��l�q+G��ٛ$n&kTP��v�7do>»6�V:��Avtvұ���}��<:mkD=DIM��A)���(Ⱥ�ҭݰ���1̭6� /qTWV�9�"6ˉ�����r߈춘��>�U) ���2(�vM��qU�߇��sB`�/~��Ȍ'���
�v����"f�z��v���I�"8Pq�"�8�����Ԣ`�ʳۻR�[�7~�n��qf�ܨ6u��ݱ�
��$�=�)	l��^�wn;A:͉���<J�:�2��sף	6��ޘ�P��m,̣���t��íb8�_3K:�?�\� �//\-UuJ��t�򱸮��:⍿�q�\/o�B���ݘ�g�ݛ���j;��s����j��;6�K��s�9�=�:ƃ��c��l����X��6��Dxe�v类0Y8鸎2^μ�Go.�pq�b�#��κ@7Cp �]5�g4��h�=n2E�&�'���]4bsӮ��)Vi{ێ�ۭ����;�vͻd�'N�X�+��?d����ױ�5y��t,��b��u!��z3�sZe�-tNF�)�Q.I�տ���U�*��t�K�U�&�J���@���'�2���j�u�w)a�UJwŦ�IF�I$�]�AlS���]�u=�:��Mu�S\<�5L��?�q�Cgc�Ew��R��^8K�a��1q���$/�IP�m)v׌}��/�&�c���l*ݾ��W�+oGW�K�	���B-8�b1*I����+'�uj[�Sw�A��[�a�齄s	i�+Mko0�Tp���n�����<Q	��Q	 ����Ṭ@���NTMfQx�L��ǆd�-h�sܣ���4}��r��y򏫧�a�xY�)���G$���V�ٙwO=�㗞
YLvuoGl6��n;{ɒ֫����?)#𽻛,Υ������Y�s$�Q��Ḙz�n��Gk{����������_�+r&�j܍��e��������+�٫u�S%�׵ĭ�;@O�e��)}�h��^�9C;m�6+�����ȷ��؄�
�HH�st=���f̖����珖*�ǹ�HY]�g�rU���^n�$�;��I�Ob�n��I]�a|� 
Cn�<���ro�U�څp�)�&�q�cs���d��s�����a���n+�^��؍�^+VX���ɛ�й������u���ר�ώw�� [��.8�p�&�'��_�o�MBz��\��)����i_}9�����]˓��~��s|*�X���,2i�"�����N�m���k�kq�xՙN*�ŝɮ8��L���.`p�Î6��b�HNw��z_u����";��٬^�E艹NT�Y�#id��Т�WG�A-�m@�F�R�woMh����=��4-�⣻{9��n�Yv(���Gu��[T׏�(�E��g�v�_�1��f���b-���۝\~�R���{.�!d��c1&�f���([�KB�W����e��4��Yn+g4�p��Z<������[����V�&�a�N����G9�m��8���q��~ǙʻԳ��lƨ�����A]�q��J�v]2��}fe�J�c*5p�nنI�d6��J������-��a&dʉ]���x|}�Cȸ=���	�ry܆�a��\���
J� ��!D�p;W�:ɫ�v,`�٨�P��Z3��L��O���N�#B8�R9!�<Y�=������{�si��EYͮ�a�.�e���y�{}1ry�A�d� S�7 1�	�܉%o2x7N7I=7z�YsxȂ�3���vY�-!���R;��6$)��s�W�6�I!I$˲�i��3���{��Ý���O[5%��l+˒���;I~a�wĎ-�i&�%H-�uޯ��j�$����-��;�e�R����p{x��	{��:_u,�1�Y�Ę� L����W��Fp�¹dn�-5*�Dh:��2��b�LZ4���=�W�����v���#�:���0T�L�����3��0��5�j&~<��ɾ�ۗ�O-&�kݖ}� �������C�^��ې{9�u��u!��<��ɝƍ[�9M��vݵ�\7H�]N�_���Z��`�4w8f�Lw�i\21�޾w����"]�g�懧?*sտ����K�jC��^��Y7����n�A9�f��esrj�@�-NgE�#�t�K�C��t{�z�!$M1n8�nY�T�'��f�ǉ����4��b���gkމ��w�����fc�~}�p��$G>J��ٰ�{���x�C�WoL�,���/�?}�U�^������d���P!]+�u{�㞗3J�]}LRKʁ�n,�z}D��'�^A�Ę���a��y|�9�vJ2k�����U�U=�(�D�=�j"����m���=*C@e�e���e�K����U����n©/1���R�ݙ�.chx���\����u���ޮ�טt�ޮ�OM�3U���������SW/y��Q8(�m�G֭Y�&�{��L)�ͬ�yd��u�+قi�54��f���9+�u�w��˶�90{w$�
�f��/uc{����v��`�U�9ö�k)L¢Ep6�QF��Zo]��er�/fج�թ�)X���T�K2p�{�p;��m���X���AQ��vfI�1��9�����u�{9����Ç�,�3�r���[�2��Ѯ%������SN��QY�fwWo�=��/j�k�V��o�(��cy�bKR�ޢ��P�hv�}�f!����m����Z{>G�����F�'[�.���DB�Ӣ�U��(�I�N�ع�bo6�딶���q�o�]h��k㽍)�t��h�dn�:R�%:VM�5�s���F��ťͼ���
$ܣFI�IPa�K-`K�5��Ѭ��K9C@giz$��;Wά�2����Q⯥��@��V�t��º���(&�SW7�ȪȃY����)�/0u��űW�r���F�{3�\�!��,m�.�46���+\�Z�����Aa��f�f��۫�}]$�#�V��MK�~��	�+��Q3z�r�A�D�KU��e�S�����>�ݘ�m��(�hwlcl�U���U �(�J�UT�of]�4mD���c�U��0b
���H�Rm@5څ�J��Vͳ8I�Y+�� �91�Ru
2(r7F�m㗰]k>�ۛx�u�j���}}�7@{n_<�Im�F��=��P��>{�qU���'�z�2�c�V��m���,x,�x��2v\��re�pOZݶٵĚ��0�zvwgJcaS��8��(��kO[ܾ�Z�=�'Z:#��\�8�M<�f8����]���<䇠.!���l�nGk�۫n9UjێVN�8������aJ�aŻRv��l������'a��qƞ2�+u��5��u8�x뱱�W�cqYTWK�2�$�w9����Mj�Q,��z����k�{]�zi]����r�J��[�@|���v�V��-<ϟB��[ݗ�7&�%�0�9vwM�v��NN�7]cl�ksٟ.\�tl�^pg���\�vy����69v���ܨf��[��]�W�v8{v�`:�u����=���Ὂ�b�Cc�z�x��TN�.y���W��\�8�3��'oQٞ�W�D�v�c�l�s���i<�e��n�n粚�|��4? �v�Z�=��8�K�pu�h���f�{n�׃�Y�H�n:�n���]�3�W ���6���r���P�>�u	uW\���\�8�tL���W�a�;�7��ѧ�]S�Z��ݝ�a�����=p�Wt=��Z�u��©b^��Ʈ��:�΍��2�F�����nM]k1��L{3㮻%l�\�rǠiG aٜ�+��h�;d�@�<����5�;K�	��j7>��;Pc`�sD6���]�Ӽ[v�z;k*n�_����k u�1v,磇�K#�7p���\�܀ə݋v������t�
�&�nc�k�!�1�q�m���Mo[���H�����9�f˱\%��nt�!�j�/p��5��=P3�vw��x�띸���.;���F��WM�=�uu�nP�ec�Ͷ8�\�']k�ڲU�]JN��(�Ӹ#.�n���k��pܽH��;r��9���@�xB��5�v���ۣ�]�l:�P��I�ۜ��ۊ�ݰ{u��f�uV/H�w��ƌ�L{d�C��������mEv^�ա�뵡�1��R�����Og�nz	�m�x܆�m�1˱�@�^TҔn��組K����$��a&�$",Ip�#n��q=�g�2�삁��,��nm�ҏsՍ�cѓ���u�y:�\�@)H�P��}\�_�}[��l�Fm��zڠ��r���!�w���ηb�7��aw�FCM��h�%W��|Y�0Zjh;�mkXw떗�l3�M^Z �Ǟz���bWk��;�wp�K��¤q�$UV�t��X.�!ur�h�<�܆�L�DV�
A��Q[&M���[�J�ܾi>.%d�@Y���j�ǳ]�.�`:3�m�v��������7�D��<�0�s/�x���Hbf(���8��v���K]�0�L���>����Gf��<U E�N_�����-v��9A!+a\]`��v�ֻfŽ��6�W)�G|�Ȕq���ng%].��gf�{�t`�K�u_����c'#�G�6^�b�c�/{��r]\�T��q��PI1D̑��3%Ҙ��R���TԒ�d���N b��*�ŢyS+NևEV�f�{�d�F�kݾ�c�z�2�T�Ӎ��3�-ܭ9y�"���j�sL�(}�z"Ø/�{������9m�mX����Əu��^�vR)�N
׮D)(�i�ґQ��5ߝ��4������Qͺ&��Yv�ך�_꫘��f�~_���!F�p��M�{�ur�x����槖�l��A\�jR�.7D�����f��=�ĸp��h�90<Yc���z�o�t�K/ �׍�Cqm����>{=��
��zC+`���+�?��7���3���ɻ@��G�����-�Y�f��4�i8$�Sd������i�yvj"�]��fc��M�l�kDf�^ޓN�;]]�<����P���H�!lD���yTK.��~��4�]�5��f~m��j��B�F�i����=̖�
���M��f^eݏ���eD�*�L��"����UlfK﴾�V��Im�Jsr $Ez٨\��a`"���b�m����:�'x'�˽�D��VUL�f��u1���W/HS�q]�-�v�1��D4n�,���<\��tJ�c���!q��Ekr��r�ۙR�'�:ik��{�*R��o�nV����+�j���`�td���܅�Q��&H��L\o�L��C�+��'+��z�U>��U�'/��e�1���4z=�b��
�֦�@n��;v�p�;�0s���9b|�4�q��.6�{/�A��1	H�JZ)Ȼ��$�hz���t]C�~fx[�~����0����[�]�3+�{-��I���M8�����Υ}��Z�z����{��s6x�/��mY9�)�.!�ǽ��'c�z��YaDY#a�[��8��O��n���vR��!G,��o.�h��)��<ӘyGZ`ƴG��"#08�-H�ɶ0��e儫����k����m��_9�=���C��Ms������t���Or�#B���@Q�$t'��fRQCq�?<Zf ���o@Owq[���	�V�g���+��:�,����|�ixD��[��x�,������"�4�V���,e���'�֜�'�Wt����ܬ�������x<۩2���RD�%��%	�Gct���Ƹ��[v-��qq-�v�=�ڤ�s]Ȉb0��lgUQ�;�Skb:�o�爗�pˡw�m3�
�|ﯫf��{�Ѣ{�㐸�A�RDS����/���믗A\�mnb�yx����bco�X���Oz�H=�G�Vu�H����L���$�i���mOt��N�)��K���KF��u��$g;+幷���m���	���e��֯���,FN*J�Ǽ�z̔c�ٹ}�E,�C�*��k"�ar�>r�vf�=��6�-�L������iTmZI��NI4LY�f׶5Xł�n1�R�Mp�Պr
5�/�\F�zY���u^E��]-(�Izt��D惸jSƮ�*�����-�״r�c���EgG񆅝D��Kީz��j;L�m��N"�I���y��tv���$�#���e�a�:�wF��GC�냞/�����u����8��p<S��>�����-���\qն�lJÞ,�'E]�'�rt����<㭮�8�'2i��>��!��k��D�!̇��l�&�0��l���v��b�u#/a�z�v�^S�ݍGn�@�^���Aюr�[�czɱu��C�s��<�ܭ�,:��Gg�3ۻc�;V똍�@��A�B0�)��RN���~�֮��'�yU<Md��ND�X��K]yK�q3eգj����i���#1H�/F���us���>F�[2��y�� D��{,h{���O-̒���ze+pW<'m@�bB�I/fe��u���n�����3��=r^.<`�>c�᳼y�ӷ]�`E#.2eK�E�'��S`N�
IPt�k-�|��b��G����Ί��R~�Ց^Ŵ�gcz��b�x��Y��T��ILb9j/n���{�m�x�>���B�nj��(���u�X�Iޝ �]{,S�H�ݝ��L����&H�t��-g*��r֌���*�ɋ;B�=	��^nz�k�h��<�;̗�x�#)v��s�If̈��c�^��@G]��}tnU��(-�J6�BKI9eX�UC��E2l��e� ���^㙯лymrRs�	�K�ը�Hz/�b��'3vH�CP��i���a洓�DhY]ͥ�\��\����v^*��K�ՙ �Nh�"��\	F6�&ҍ�joF=[)h��u�_��c3jƮ>I��)��������9�7� ��b���H$)�~{�6�wp��f����E�4ByIH�*��Ky+n����8�����I#G�� lO�m�vk�$���n`y���^S�dLkh��I��X�\�ηsg7}~��ZZG�}�b�$����0B�=+�o2u�Y1GE��5ێ�f9��>b����X� n8�6ܝލr���2��;��s؛���
ꨨu۝j�P�����|�7�C�mHC,6������5좶eT�s��]�����VT��{ɬnk��c�5���fʍݫ\��K�_��)���un���"{��k-J}����y��˾
�M�;�Y9�ku�ݹY#z�-͑���|b-��Sq16v��Me�׭Vd�0(�Y�U"��g4�D�ꚥ��i�v[��;�޼�Xa�T���I	#�E�c�s�+T��Q On���oGD�1�M����t1�Xu�3ۦ���.\p�-7��^�]g�#�U��ٽ��ٲ�땦�>�U��B�v{:�Y�X�9���9�Q=ͱmgN��*��	^�9W��x��;��m���C�l5M�+���W��~�ލ���Ĕ��bb�k��uܗ���W緜={hK�D�x����9	8%%m��v�"�q�����>�ș�nA٭��"�^�wyS{0޺���&��^��T�|��I��7ᨉ"���${��(�ֳ�+�y������xz��Z;�1�j�Nl��m�fI^�D�D(ځ������K`y3�����Ʒ
�&5��k+��� �̙�ʸn�W�g�/�U�cR1��P����e���;4,��Z�T��~�uη��{�n�tl���Q���/0K�{�]�vՙ0�&~Wwg�喽U~d��U۵֗V�j8������S��Yס'�j�=�jnj�7Py�,�1���.�_R���hԣ֭��:q{�H�}�8bz��8$m�0��I0ϋ��=Y�5I�<*m��]Ռ�H�<;��U�<�`IR�JJ!#	$+ㄠOw��Z�\��B��Awqf����6����W�/���R(≲���2Es���i���acP~޺��9�o���bWbbN����N}�_f����D΋�^es�x֦��P��M${s8�ϕ�{�M~���%�l`T�12�ɖUp�j�g8^�I�X���d_lvW D�e�Ӓ��+��
�ү��^`<���F�u�N�k��n:��N1�7�Ǒzx��dtw�`� �bq5#�Q������j�}ٴ<|�Y}Z��U�8�y���o����t�1�b����ƫ��,>��i�u�e���0���G/.����c}�ہ�X��ߚ�`�1�B�,�>C��Fp��2�#�T��Q5��;�k��â ���^1Ӈ+�%��;o#�\n���8��O/Q�����ŵRA99��F79m^�g��y�}n�����;��c�;pd��.��n�g9ܤ� v4��8lh���[��k���qDn	�#��ۃ�ϻEn�z��7n,A��US�����[�u��O7LOYg����;�4�,�!��f���2�iҾ���=��H���XZ�'a)�^�v�n�l�q��(Xl���r��~_��/ �`�wo3?s|�녢9�up�t�v"�s`%��
1�Zx2yܞ�w
��������+R1(�����M����<��t����f��{PX��� �)E�GY���	p]�ż�śO����wy��FU�M�yeOU�$�y��HI|�6B(^��v�O�Sw��"�������[��<���Dw�<�}:
B�J8�n�_^P����z� �RF�I��r<�wS�|��\��^yLV�KC���m�"N��CT���Pw(�u�x���77�T��E���ff��Q��nW�9�jqE�㨛�1�N;n�����%Z��'c��=V0"P�]e*;EĹ�`�z��S�����V�F]�ySU+��xs9�"�dE+RI)����Y냤��#&�w"�w�Cwu��Z�/�Ӿ��<*���qW
���;bf-��,'�i^ν��a�;�|�_p��\�"�.��5o�&:4n-s�y���lq˛t�����M�>j(*Iap��~�.�!{�q��-��u��L�{��/PN-�Ws��hk'�nrBH���i��@%vgye��~�x��x��E�;�,%`���>�
���׫(S�g#�ٮ�|��p�8�c��v$����D	��ǆ.�������>�k<^xjy���N��x����=^�k��νʹ���d0�Q�iG�Q������ql	�M�n+{Y�5vG�S:�v��anS��ą$�+S�ߝw�FL+���f͉�5^�>��l���������f�o2����ِ�ڎᲰ�����fl��P,Ѿ���(����MOE�C��`��$)>�K9L��*II5'��z�`�ɐ�#�	r=�Y��{�9Y�l^a�gd�V�˶5�m0��׍�]�U�J����`n��X��*�bo0\�g����t�t�^JЂhvj���I�L7s�-�����]V���f�٥gT�V�#C��=�����ky���k�vh0֡�!<yKR���)bA�u+�����n�x�o���քMr�����S'���va���֯`�O���ʰ.Z�I���b�q��["�H*���c�
����f��l����)��eq�o��K't{��vKz_��)�WY���P����T��¦�W]�u�2`���W"�f��SB�F��kK��W
��#���JɚU2�gv���ÂIj�cWuxtel|Kƍ�2ek�{�Y�Fi���8�O�£v���ut]�{h��:^�KV�{�VX�`�
�55�H+Oؠ�s��	���eD�G��[zC���|(����Mը	�b��&iE���V��Y�w1d�YCm��C��t��	X���e�3�4voXL�nN�]���A��/T_k�ٚ����,|�\Է".!�6�W���Li�D������O��w��<�JW+� �n��N�5`�_'���,�٠�4dJ�\B�Q�7��H���2���S���Bi��z@�(r��{�wK+��p��L�fʼ�T
ϕ�Q���8�����4�`�n(�O5���@�(��H��t�V�1@��n�yh��4�v���O�SU�|v	l�M�W=�;�oM�3P�+U��{���F��V�DO|��ó��{u ��.�ᵚM�;sZ{;��n�AD���q)&��N|��x�	J�yW�KI;=r�gc(����o[��k�f0��/����KB����G�B�f���\��;k-r��<�Ӟ���(��ahwqvьs�f2�(�R>���p����u�����G��v<4ޑ���Lx0�0ϕmW�7���E*5Ts,�5Ϋ�X�
��gE;\-�O?u:vn��z�ؿ,�w�,��� � I����n�����(������K�W��|���W�J$4��WQ;T���[#�8!0���^R�T���u��0:��fG1ps�������o֮;��r�s܎�j��^�)Xj��W�aUl('�F��I�� O%�ن�ǽ�vgׯ��cիe�F��a�<.!��Z��M�i�N�e8���Æ�ZC2�1��������@���,_7Zyb��9}b}Va�;�ץh���b��aO;}	��1"�m�A�-���D8�N���p/V�{q�mA�:�F�ܧ;���=�̗t���k�����l��KY@�z��hf.�3��/�np鷴�P*���3��y�䔅I�SmŻ�J�Q\:�m��h��s�w;-��y�򾭊c���휁%�z�<��<�����y�`���&`���i%��ΨOo���ۀx����8������M�X-�8]���khX�^F��TF�PBc�F�oM{����Xm���q+��h���N~o�k%8��S����ݞē21����)F)����u��[�P��VvȊ�pW&5F���9�K j�����wi���o	�vz*�Gi<�n��kN#!Iwf����;�Zu�M!��C1��;۩(��u�N;���uz+e"|�I2� !��ʆAiA�s�"���l=�˺z�n�;Ҏ���3� y;&�q�x�n��
�{M;���a���+�Q5q���;N�n���##�sܼ��p�f���rn�t�4\ۯY{VU�pyz!lk�ϱB�ۜ4m�c�s֎<�F�&�+���ٸ+lůX��ֱ�������6���#��7S�v�O\�ؼ�p�ݶ�nŵmgsd��ۊ(���v[+Y6OCp��wq��Ƀ�]�3�6���X�t�3%#��E%N����b�_mu͇���8��t҆4�_YZT]˲r�����"�	A9&�k�)�;�����_aܯ0�`�|+ݒւѢ]�{�K9Li�\ݱIw���g�pF�p7LFⵧ�=���~#6�uܶ��64+ᡍ�k��O��7�m�]
G���@�	2�y���5= KQ�0��*��Դ�|�8��v�b�ɺ|����jn�ho�����v E�Ą6�r/��B�L+೥��An>��M�ޟn�E�����$=`�� ���-`�^��[D�i��������ֆ����+�'6��;�<�p��[l�qb�F���3#U�Ӧ�%��6��7�n��D���Yc"��?k�$n�����=Yڵ�*�wM�M�	bBSF9,e��]O.�]q�#O����[&6B�U��iUYt�D���'��C[���_`��`Od�m f0F2i�v��D�&1����M���wL�Y�w)U��ٲ�z5(�yv
��4��µB���]i��zk�
"Rn#P������xU��v*��m�E��2{�x��1u�N��oQ�Z�AЍ�P:��	�#! he%��^L��)��u1�v�rU��xQqF�{�2���^�O��"x�3ҹc��n`q�rX�"/�|���y�¡p�F�6�~�\T���NU�^bw�h��/���V����KWnx��ts������rco&��&K���N8���<�����XR�s���w���K4��~5�y9<��{w�NU�.]������p�MVV5������p�SDCi���ݲn 统]�����ܫ��ޓw��;�;%���J�[�ޒR��Ď�]�.�)�!b�-�&ў-�Ҕ�^�-y������36p��@�g�J��X1ؼ�,��\��I%��.�:摷C�y��T���9sw#�+4�<�-ܬY�E�|�E��wNT��g�ծ���DA�Q$�J�{Y��A6J���잳xaݥzx��״wM_n���.�D��L�~�'^�j&�iA!jr`�=����4��w��7��qfFM7^�yM&����8n�1I�k�<�:��Yÿ/��{~w�����Vs��/s�8
�ۇ�5�8�=qƭ����^��	5ƛ�"%��˲$�?:���μ݃���G�ӑ������`\���g
ZjT>\��E�2���3*E׺a7�,�����<}3]dz��<�yh�5�r�P�k����ӹTs�޾���9�-1&''k���ls�Aן5��*���;�.���К�or��x�{0�\�S�n$���4����N��A�dq�5z�ٴ���*�x1�7�K�-��*<6oT�7U�� ;��m�'%n���{�����;��9j�����[��9T[Z�Lae�:,ӡ��u7�ߊ/.U���/Ip�~|u��	Ș�VJ�U�����ÎD�t�]b#�f[�o�/�*'��e�^���%�,�Z2m�J��T��c�j�qBZeɮ����N`�.qo^�S�Ƌ��
c�F��,�$�ƃfBE�g_�`�N���F��Sރ:���̫,�:*�	z��]ٖp�a�E%�9шDcI�I7/z�T씫����}��ª�#��e��ԋT�:���]�F�W]9{�t=)R���Mjz�lz�I��Pb�I�-oҗ?>w����C�ٷ(we�K�� s!K����@Z\��)z�6�6��z
0������03�zזh�j�ֿYC��]�����Wf�gl��6����/�CT�bWm�JF�0A�N�����*�0��1)5��&�j�}}�i�[��j�^3�'{s�����#h�sg1�>�Z�uB��V�Ǵm���,@Gh�⣕�x2X��)�����O�`k��d�F����oq�f@�((��ENI$�UT͒u���ld��5�]Ǡn���#קF���.�/U�؍t�\1iK@r!����m�n,[>h�17�ɳ�Z導�'<�u�6�c%��]� ���#��`{G�����mθ���l��p�e�;���\�硋�m��:0D�S��v��֍k`��;r\���dx���ێ{��u�8q�UYyB�'�l<P��C��=�����.z�++<j鞖��؋���m#�Dd"d����S��&GU�Yܘ�y���}O���"]H8;�[� �o�$���2�[�Ce���ؗ-$q�����(���e*��6�-����ߪP�T�k�j��M���������-�N�ބ��5��`)�ݢ������j�)d,���˩���ЪF�#�:�Xda7N�����nhUή��|b��L2�n-�X߰Wo��"�*�����	�XL1��c�������r�����W��1](��w@��ί��=��x��_�v$Q��CޯO˻�R�$��9$�?�.�}0f鯟�.3�L��|�,�i���e)�2�'��,{�k���̇Q�ђ�_����M�H��n���v�X���[�+I��R2��՝`*��P{7vv��I�p��7")�M���7QCEI��KNM~�C�
#ݟ�:t�R?�Clad_w�;�h��0�}���'3��1�pF��C0W?}�xJ������Dv?���P��j@܈$���j���D��?��O�f�G��N�l�lIY1�]�ǯ�Y��r׉��}b�F����9��݆&�X��Cvmf+!�\8Cn+m��.o#��'�^��u�����B�-l�����K���L!!z����5Æ$Y>s�����Ă%��$M�0�$���F���u�����(x��@ rP��,8S�b�^
@�3�y��]_�����͜��&�!>����'T��.�ӄh����`bBP(� �_�gE�7�Y�蟾G峳��#�=F��W 0$D����WƨG����Y��~�C�%15	����AM�/?^�$iq���<v�"��^���RQF�)�vIԏ�Y?a9�~�´T~�L?С��cjl�p���p�ن��l<Q��
��E��b߷��da�lH�Xa���KG?��!��L�ǋK;�*�q���Q�yベ�����9�G���jcv棗�E?�������m1)�~�����2�P"�����Wو,KTU�h�6���0�+ɓ��/�{��4A����ݘG��6G�~Dd�ѐ��NEb�dI"�. w��6,����u��;�g|"�ے������͢F�6LO����%k���2��G�W�,��M4���c?v\�Y���E_�a����A+H���8��^� u
0���t9 �K�PY	6(��C��*� ���(���$��߿d_��#dm�����ѷ��^�d�y���D�h����S0�KFD-��e�ݝ[�ᶌ��Uݱ�y�A�2�9E�*��� ����]���#�n/��h�?w�M�L���E�6�8��1� ���|8A��3�����+z��mY�iTB�w�B�	�|�Py�N�����p4[~r%�e~��C���*�my]�:�R�fa����R2[&8�I�r'�� ��yL�Wª8z��1���@����yN��"@BC'�(H� ���5C�Lh�(GS�0@s㓐����G������H�0~(e�dI8�{n�pZ��喚�c��*��Ӯں��rqؐi�rRFE$�4�8�#�)
��I��+�$X����s��\`�)��Cu0���⨉�
"�d����������ѿ�qY�c���O�>�e����#�iȳ���)�9�����(~9�+v%A�+��4w?rw��(!�DX���{�z'��+>t�|A	U|����tAq�tJ�	3�m�s���������s ��*�t�H�qTi�h�#�o��k�Zl��z)(cA	�����:>��N�Q���}�)@WV�p�cDP���Ƀ8=HQ�#M0X?��֙�1_O��7��̏a�w�>�o1B/�<r�B�1��������+G
p�?o�r	�~ˣB����+&�X��@_B.��۽c�1f���bI|s>��e�,ޙ���'CU΃���;�@����+V��9�v����b+���s"�I@$vr���=���ں$�BȲ�8 �6�9�tb�w
������tȡ�"��ۡ��j����utj�y���	�(-�fb���*�x@�$�F��g��l�������<����2�;1���d�.�;+�'f^�K�ͺ�M�V3��R�ZIo�V�M`�#�~�1CF�0L4��t!����F�HU�#g�|"@��S��8�U_eIQ򽏆�_L7<!֌����/���2��_�+���rTt?y#�A�ɣ�Y�fO~������w�oLȏ�!
4{z��p�a�4"`AC�����,�:���sQ�� V����c��u"�4�����LjB�nDK���e�t��XX��/?��lx��d�k����~�v�mT�����T*{w�OIyʆ��q�u"�aտ�+���t��� �~���T@�qD#�X�!��Y���yx�~����-#�^zg׋�Xhc͒i)�_�]��0�	Q�vh:?:5\�Zw��~�1��X� ?k}N��W��7�d��H�{sԛ��$@�L ��X����+�8K����p豢$Ϙ^��7���}��1z� V��߰�V�h�߾�i6��%uB���>����%=������������ %P�P�� � �7��p���UA�̡A��z���
>-?��ߏ��=>�_:$�*D&)B���1T%��O�B����l�
��p�Jk{�(5(Ps���6�(爒\n�i��|gem(Pt�(Pr����ל�A�P���z�g�Fw��r�z��z��~!UH���?��d�Mf�	C�VY~�A@����~��}���|                         �    = @E!	(QJ�	��@ ��   (
             @�QQR@    A}P7Y�
������kV�US��gU^����P��=�Uݺ�c����u��:�
E=�p��ě�x�v۽x=����[f��u崗����6]�
������[m����)U�w�Q�x�]i^  ��(
�   ���+�USu�V.��T�s��z{����u)]׫F����*�n��+�Ԫ�;�{�@K ���^������]�T;�%�^kk�y�5m绫�ko=��
��5[�T@�z��m�s׭g�w�^绯b������@�JR   PR#�z��޼���oU^[��ڪ�\{ګ�H�/��޹����[��O4�����s�@U�{Uk��z��{��m��=�������ս�1�V�^�:/Y���n{{�*���v�y���u骹��*�{�R���W�{��J�� IEJ���  
��B�=�J��z�W���xgs��{�@G{�[{������6׽{��ls���ٝ��*���==iW�p�j��ޯk6��ڵk�	wz���=kgzΊ���ѯ��ky��*�U�g{�U�=븩Y��U�{�uW�� �I     @��U�]�^ӽ{תZ�n{:��z	w{cm绯-U���{[�w/cW�{��Vs�@W{ڦ���ǽ��z�ת[��[T�]���* JޞZ��r^����^�y�꼯=�y�/z
��[]뼽R���^3{۞֚���ک�  ��iU* 4   � S�i1���F�`�&�*���R�Pި�!��`1 Aت�b�#L��F�#����Q6U*�� h� !* ʓLJx�4�OP=F�i��i�O`����������:�����#׮}{���
M��* (\�G (
�T@P2������D@P+��ӀQ@�{�Ң* }_ÞD��O� �T~�4�q(&� <�(�@<aGH<�^cJ�iЋ�hU�t��
'� q 	�q ��C�H��H�͡Ut�T�t��M�J���AgCͤ^$��!�̺�QM" ����0<H��4��̦�Qx�� ���@ s0��*�qq ��(�0��Ю�ѥѠ8������HD45�P!HPP�t�ATRm�(Z��
��	���kV����N$+U�����I�֐���)I���B���
�@Ѫ)��"%�B��B�62��4�4�U)AEHPP:Jt�ѭ-lE+E[-Z
��(��((�J�M)c�)h(&�)H�(
��i �&T���J��lFi���RQP�&�БQD��)(JR+HP�5LTąU1Z2TV٨�1E$H�ITU1���4��J�S�(:���4#���֤�:
"*jf�j 

�b""#A�������*����� 

h�ֈ���2hJH�iWI�h1R�P��AZ6�1;Vq�P��9"�b
b������N�Z4�SQRl�""D�EbI!��"���X�l�gEUiӣUZ��D�	M�M(Ҕ�ATIE!��3EM&�PD�PP�hM!0`(K	A4��)R��"�ӊ����J��(4�aIU�BP�%���(�!h�ZE��&(Z
60DB�d��Ge�lIZLC14�e(v��QT��UV�"Zih���I�aB�sI�*���D�"]j��
$�:vMK�E!B�(R&�*Д,E%IAQ$HhJS0��TPRm�(-�ZR���C�

i։�Z�ٳ�6�� �AF��RUSDN`�Y�)h��C���MF#laf'gU�K�1N5X"q4E-B�0[5N�j���.�$4.�`�" ��
��H((����(j
��&�i(��R*��hJM���(���tm�ĄC[kN$��&�B��	���֍Ris���p��c0N��i*ml誧Ψ�X#b6�DVt����ch&(����ӡ�5D�M4DET�E@Q1V�����"Bd(*�f�T�������DM1��M���Z)5@�L R
Q��(�H:R��J;b�4%и���6�Fڦ�*�]�"hZ��#cA�-�J�ULM Q%�6�gHڵ4F�1������F�6�ӡ(J4��I��X����t�%X��b�F�i&
u�-��%:
�j-[!�(h�ãHkN��t%	Z�Д�-lck�H4&�Z0%4%	BP�%	BD%	AIN���BRPP�$N�BP�%	BP�mdДh�&MV�5v�hJ�.��3:4�c!�bJ�b�[Q���h���ڤ�ERE���(J�N!(uZClj�jZ΋m���E���V��`'b�Ƶ�bkh�LA�ƌZM�Vvӧ���h�)1�m��.��C�Clb2��Uiqm��	A��	BVf,ZKV�QhtZ�[	E$���N(v�md
j&��"Cl�Z�Pi4�&��-�&�Ek1��k���Z�Mk�h��Y0Z��D�Ѵ�h�Ӣ��l�2kQ���RN�#H����"�R��CT� ii(
���)�i�h
(Š���9MX�)��H�
E�h�P�	BP�%	BP�%	BD%ƉkBP�%	BP�%	IABD%	BP�%	BP�%��`�(J&��"��(J��(J��J����XД%	BS��f5�4�1pcX�6
��I�ӡ(J�N��"���(t�J��(H��(J�����J��(J��(JB`�i]hU�A�1I3JRUP$��4	2
�F ��h��(���Tm5�J
(�4�h("��,m�M���эi�t���%��Ҙ�� �Dӊ�R� �!�(��P�ɠ���6��!�*��("��k@iB'lP�4����WK�a�F��Jh�@��D��+BP�%"U%[����BP�$BP�&��(M	�)�&�
A�P�@�I�SY�+J&�N��]tQh��	�4&�Д%	BbBP�%	BP�%	HldJ�cR�P-(�"�+�@�&څ(@)h]($�li@�����SDm�gQ:q[D��d�!K�EXs3ɠ" i�H&�h
t�M�+III@SI�h�(Zh!*�)���f�mV�ء(X���N�EDLAI���l�1@P�ihCm� �kQ��ŝ�Vƪ�g;P[��DC�J�Q�4�Z��P[R�lkb4��gLMP�65Z�Ӷ��4`�Ӣ�m�RmlT햊6֌�Â�LP�%6Z60�ք4���(((tA��)"�c�X�2Q@�;j+A�4�i(�(�����KM1K5L�bt�N#K@M�Ѫ��(�M�LQX�ղ�M.��բ�	ƋXѶ��pf+Ym�!BP�%	BP�%	�J�К4���a4%	�-�5i�ūhƊ3j֒��(5Q�E`����&�$��mDim�M����.*(��Q�i-8(КӠ��Hlmh����ht�#h4DR�2��Qc1�F�X���c0gb�a��T���4�	M�Д%	�%	@clE��F5���!�����Efˠ�Z�1��b��(J�M���Лa(JDP�(4����ˣBD%	m6��4gZն�,Q�����&	h��J�t9��C�)hJ]���%�(P�C��PģV���Ѥ
�J�$�i��	t���b�Ji�(����TADi5��EMQI��:�D�4��"i�JZh
cVƗJAI��le�N�6��F�LDUQ5MZ4- P�����̊�����?i>�Yov�������,�h��|v��|���Lm����~�g��~���EvW�������� *��UE���   �U@TU  -�M�T U UP [#����nނ�� 
�j��j�m� �uPOT��e[   � m�UV͡�  �*P �EPJ�*���U�T
��
�JY��UT��VȪ�     +( 
��R�*�wU` B���J����> 
�
��l��� �  26�F��  �+nm�Jl�6���[��q���9� �m�B�{b�W�)�       6Ŷ�W��E��6��©z�9��zU[8���+O4�Ѹ� ^�]I�*�n*<p��<W�l���n;���W�����|Ul��V΁� ~;�뽊��n[q�U[hU
�uD
T ��%��*�Q*�=T٤R�q�lY��M�� �	�®��0� ���}U�V�{d�����`�݁���P;6�!T�U9���U� �P���#���Ԁ*��1�p��P  �8@x^�'*���8@yYC�a���7���R�.bp2����18l%h���m��� 7Ӹ@ �Ui�U++R��U*�;�Z���T�        �6�T l�-�VǨ��k�  N ���� ���d    �Ҁ��UT�U   6�� dU*��*�ڷ�U��@� z�Q���m�oS{n� 8A�6�j�[�\���W�8�r���j�Bpu���zU["�����v�]EZ`A���m��i�g
��e���`�UՔ�P�e`ʧ������8B�@\�)�S]��V���NR�"fA��s"l�D6�F�rm���J��ں ��֨����nD��%�,Wu����)� ��� p @      ��� *�j��Ai7�,m,�U�N�l঵R�Hn�M\���lֱQ��  <�' c ��*� �����}�М��S�w<�#<���vrV��0�]Y�,���ZA�U�k��Mz�͞�.`����{����V�;�:s�^Ww��۞+E�6�e''3�6�B�C��. �R�
��j��VS��Ϳj�� ��C��^�e�R�j�{)nʮ��4k�j�j�uMfU��Ux*� c �l� z�  '��t�� �������s��1�g� <sq��Il���.���qw����U��!<;{�mv{��(*�Ur������o�l��۽�m��
�lʚA�� �[Ku�)2�Tq��+��g��u��ճ��&Ij���Q�]l��<wg�d�5�T���*�R��@N �c���۳3l텗��	���ݝ�J�1[:���
�Y,�4��
��J��6:�S� �&8�Sg�]�xަ�d�lx~�璨�U{���_U�Qv�����oAB�T;
�ڢtN��Z�Z�yQW�{�V��~��eޑ��&�*�Qy���y����3��w־S��1�l�ޏ	��3p� '�������U	�ʁw<*���諭Ψ9j ׻hN ƶ]Z  �)u������1��[mA�x8;��v�YC�����ݛcӋ��n0jj�ym�)��Q=i�Y@�^UjSd y�Q�;���{��Tۻ���C�
��UV��)�gڤ�m6S&̪���z��47nw̟���+]�[����]�K5�@j��V\lunZ�Q��\�H@��vA�#�B��.Z����+V̄�3�0��n[��W$vݱ�;�z�Y�7\y�k���{`<�Ҁr�l�,��?v�wzz� �a�k�;m���=��L��?1;�dj�h��r��c��6q0M�    @ �
�e6gs���gJ�uLkt:u�1���F{���u��J�*�4��ɳ����zP�Z=n��e���*l�*�J��U@UR���yږgusT��  P
�i�uY@�Ql�=m���������u�T{p���N�[S+�A���@*��I�RöJ��l�km�m �n����5��ʂ�ˁ�%�L	U�L̀��[DS�r[��O�hݍ���ys]��h؀ѭC����B�AY.+"�6�̫*�����TP�ac`��أNf���@n�̀Ƥ�c�d��8�,���rح��/N+���'`;r�q���[U���%��A��v�5��ƷS/�Eqr��-,�S��UAEW8�7��9�vLd�9ݲ�-����Ɨ "�7b�ӬPv��K0�� ��=�-�(7�]*�g��VP�{%�t��q�v[�#�hU��m��,r�2�l�L���9��l��K��zU�W���]�FxM�	�1e!�[��m���ݴ��T�� �k�����W��e�$�̩�'5��n. 9]�ƹU띕v�q�.W��U�O�b�Y3��6�  �ھ�����#)3��`��<��[m( VP �-r���UJ�*�oN(���� T 7
��n�u  m�@��6�lv�n'{��  ���f  6� m��   �
��P   l[&�n6�6��?1w.��qʹkvc%s�jZ�7�s�0m�=�V��Yu��     U@  *��
̠      U                                  �   T �� *�  VP *�l@ݬT7Z�U�e@V��  <�  �*�   ��T 
�n��{������  @ 
�Um��]��Ue*�u�����T��e
� U[wY  �
�UTb�  T    z��w7h  *�          T@ �  @  *�       ;� V��@@  � 
�N`*�EP w�+*�n�;�      @ -����Ԡ���@��B���F�*�R� lP*�T*��@�6�M�d�T �  ;���
l
�
��ΰ
�   *�� U�;�����"��	���L�\�T����n�w�韷cg�ՠ               �          P            m��  
�                   *�    @;�@����Y��U    
�  �     �            �P             x        
� �                    ��ܪT� ��    P p  
��|  ��ٳZ� YJ��U^����   � *Tn"��sR���S(  
�me� *�m��l�@ ��_          �    
��@WV� تp@U    *�f@ *��[ � �ؠ    *� @  �\�-�@+mAT     A� ��                0R�T��               <    ��  Z  �
�����	��8@x m�p@8@x {��Tw *����                      P�            *�             Pp�        >��         � 8          
��           �    � U   n�          ��r�V  ��  ������@ �m�AR�SsT *�J�PT���(@J� 6�-��� �S�m֮{*�T         U
� 6ͳ�ݼ�-\-�QV� UeU \mV����U�
���o;��n�  ǜ��w=��M֙��6�  �m�{�WOf��               PU   p��     r�;-����mu��O
�J�U �EJ��v��� m�����m���� P         =�k��7� ��*�      *T       0*�T[ l@  9۰U0�+W;�{b�]��ks��s��(��ʂ��}<a89���������#�>��/�C�|���������P dU;��c%AR� �T � :ʀEPM�T���Q��'b�n� �:�v���.b�;��TN��d����k�s��e''c;`�VM�8�
�uk� �V#X�Ao�k�E��]�  +2��Q8  
�Tp c-��{�����ѩ��[z�*`�����Eɦ���N,��5P C�mV��]�/T��q��p�==��ٜ<
��=�p��Յ]W��]�\�u �8I���M�U�V��l���p^��r���<��8*<*�g�Z�N���]K<X���uP����\uh�[v}]WPV)�OTꀜnG��'�;j�b��lvj�.İ���xۑ�� (��ģl����$�X���;V1u��*� [K�v�T�T��� t�R�x��*��j�wn�SaV�w�Em�����V�.��撫=c{�q���g{tk���n]%��,r�mںm�͜�\ŗ] ��
�*�@�[f��
�"��Gj؁�r�Ln�d'�2�ćnīU*UTp�xm��-f%s����*�n����+۹� U        �J����U ��� x��*�ت ���  *�  
����2�*f��N�*�a��ͪ-�� Um�\p���  *�   P    ��Sj�UT@ �    <    m� UB�T��
��p�6m�  T+%@�T�� U �� UU   w@    � 8����    ª P  � 
� *�� \� �+(  0R�� *mlVڅQl���� ��0��G:�J�w�   @ ��U*UVeU�  m��@  -�P �n����~�_>J� ����9��jX�+r�]v�zm<���j�[v��Ӹ�)2�m�VӺ,��䨺����5jv�$R��մ1�K�6����I���N28�Cё�Ò'�a!��l��q�M���6]U ʫl�;�8�sgT�(j�m;���6��UT ��^�`T�Sa� ,�� Ux�-��@:��m�mJ�LjjU��ިЩ�T��y6Tۓ���ll��D��� �< H��W����)�(g�?0�n����a��!�b�e�p[0}	��**THVFKk,�ן_�;p���(�aV�7N
�{A������8�u߳�مe(0 MY_1�<|�@3��Ɔ(�^���UdC+`���.���
 ��a��F�j�R��š����n�XU�y\�A�7&�,V{b�Ph6a��I�`��B�*
�`s��Ab��h�7N
�{AX�-F�i��U�r�v9�;骝�;{y���e�۹  �Z��M��m��pv6�m �#a��nbOE!Z3/o�l|��}�Z&̈a`@�h��ö5#�c�1J��c���hR�E�+C*��h�6>��nJ�45��Ey�n�e	!d��a��+&ڗb�V�T����X�)�Z*ӂ�<
L��@*	\A��L���=W���Z3/j+��Ɔ+�i�֋�
�h�(���a%,`2X7���u���+�k�����$0Q�� ��-A!�_��|���%Z����F s*+�Z��̸M�P霏k,�c�`*�j�T�5n�-�%U��T	ku:���>}9���z�Ժ�ق�+Q���69�|�\~}k�ج]�Wl��2�TbC����p!��U�Q�
��s"�+E٥���� ���"I6R��B�%�/��kH1���`|{���t�f�!���zl��w�$��� bv�2u�}b�>W���au}�K�Ί�1�Ʊ�賵�E(�-"���q�`��
�Tt�S�� 6*#��X�~Ͼ����'��� 쩔�TY����Bh:���)�۫e�V�kj�d *P9�\%]UQ�W~o��}�KE֋�ExZa`A��V��W(.??���Q��ֽI�Z�u�	��$�lAw���M�j	
���;�
��!&P1��̺�l�D�AJ�M�YB��%�b�V>2­�pU��N>����
��,�����QZ�VU��w޾����,A��*��Eâ�Z``A���v��E��?ak�n%$ -��6��G���Oj	����;��vfg`������!m�6�@gs��9Qإ�p�կt�]�^�*ke@UPmTKɋ��9�S��wZ:+ P���1�z*ƌa��Ǚ:��F:�q�,n�J@��Y#a�PxnO"�"�]��� �e�Iև��4����+����"� en���5���E�^j?x�R�ע��OP��A�ғ��B�w��̄�Ɯ��+)�x�_x�u���^���6K�N�V>2�/5��8��r�����m��P\�G�*���0T�y����vW��,A���Z.��V���m$� � �m��y��[�P{Uf�=��( ��Jݑ��mR�c���掰*��WOc�gm� �Wz�b��U�!��zر����ûI�&Yf��@�����eO�+�u��M��J�@� �fU�@ w-��eOTw��J� *�(ح� ��u��!�AT[!�z�n�r��x v`W�>��Z=�v����m{��2�F3�r����H5T�N�m e�\�"�M�TMP��
����,h�Z�E�8(��k:l|��PHpT��F�U��v�`UA�J�9���a�#&��\FC��xؽ�F�ܭd�B��G#�c\y��q�@��i���0xA�����+E�^�p���W��d�[�E���7Z/��ZcT �
��mʸ)�6�#g�����#�"x��4<�I��tb���'���hbIe�h�m�.�`�^���9��1�l(n]/ ��%��=�&kU�r\�q�!:�H�[aT�m݋,��۩�9�m���/<��_鋕y�~cB�y}aP��#�Eh��6cW�����ҥlKK�
�}�}�����,xV^�Z��������Lh���^j?�:y�J& @i��>?��P�+E��w���%�Z���c8�����ח"��Ej�*�p}��$Ʈ
��F�h�+C�{i�B��ڨ��׀�c!��$�*)�Z3
�ԢU}�Yu���X.��j�AX�1;��h��f9m$u�B�v9q�{v%z��=���f�w.Ȩ�l�m��w�tXHP#RcQ�N�<�p���<>���lT�w����1:��>ݙ�VY �GKhRËτ�_<x���Pltw�*ƌV�EA!�WOe8�ǟE�s���-m�G�k��OcW��0��J7PX0�6ӭ���_�<hx�^^z5��-��M��t�f�!��0P��6~b?��A��9�!ZSe4PI4ZA��� �{Y�Z-��}A�n��pV(�d֊�C��_?�V�r-ҭM���7a���@З5�L�l�ol�-�d��m�w��"�amn�j�:�q���
?d�Px^��nꈭ�xiQ��>�	�/>d�]k��)�88�hA��A&5p!cG�Z�Z(�i�^@f�>bzʂC�����,J�h6KI4��SW�hxjI��A���/E��� ���TӍ���h�ƙlM��@%M$�i�,T$6*��X@o�Ca�Px^���F�x���Я ��3�<��[,�)$������t��>��Lj�<6���ӂ���5��}y3��-��%����n�uA�K��OP��v�[T�J�T�l	�cq�+N����2u�3�w�&P1�u�z��Uc��}[�V褶JZJ�|ƺ��(�6+Du�)���)V�46�����h�3I�)��l6�4-�PX��"/���Y��б�I1+��h�cY�n��եH�Z`Zi��w���M�A��<��4<5$�>�g��3� i��$�Ȫƨ- �}�e���ث��U��������o.6�D���� S�k]���^��h�񮠳*���Ag:�m�?��|Ͳ���Z�Uz�
-�[v����0�pK�V�Ue�zn�A7Q�qcBD'3΀��9\��������Yې gs"�T  \\�T +u��Pw�Gr�l��eUP 6ǀmT �  l qS2�T�������mmT/T�%���)�a��J���� �g�l1�����J�����*�5�j��V�2 []e�Ѭ}��>k�X��0�O��ExZ�ct �1A&5��aT�eJD'��ɭE�I.yE1o�V��d�� ���$F%6h"�.�E��� ����h�A��U��PHlU�{*�C���	�-4�j�mR*�3����{A����H�N�\:+��
�?��_��V�*�1J[m��e\Ə��h�7N��f�>bzʂC���q�+�
іd$�h$-$�j��V�6�u�-��^ow;B+�[h 6�V	%��@ʘآ�U*)�P1�u�u���^A�@�LT^
�F
0�5���lܵ�*	�I$Z4��[���s�[��c��V���Q�PX�?-$�C�ExnDM!t�l4�D��AX��N�<4[5���8(��k�c�'��$8*p�p�S	RM�[T[-5!���I��A���.�+:+� �
�(-RpT��7L"�E��m Q�˺Z�D4n�K�{� 9ov��D����e�p2�U[�����8�:7q�(��2��D���J�TP�Im�F�:s,�m�+t�6�����4�WPS0V�UH`�+r���c��2a��$�- )؂�W��G<��І�m���?WkLag�:t��a[�bR$�I�I'L:i]AX+p�F��R����(
E�tu㐎2��/���'�#ǌp<G�4�=����<�|�P�%%�M/�Нnwsݱ��q��@ȴ3o���ߛ������{�{��u	G��� s%�M/3�/v�pN<{�^9<&���J����������K�	O�'Ri}N���.D�).ri}u�!/6��0a�CA�� b��}P}D}���%	BRw���&����%��Q��ԝq�y�߾|>a(J��&��Y�������w��&��Д%����^�i|s�!=�	n�n�7�?_j����n��`{<�n�o)<�,pݭ���[����T�� n��d�1nh���q����rPO�^��y㋗�%Մ��Ri}N����nD�).�iz�<B^,%�:���2w&���J���:�N<&��Y��Մ��������{�ϯ�̿�#u�X�O��%	BRu&�׬�	Ͼ��w�7�(�I�M/S�(J:;��d�M/���%Ք��'�n�~8<&��Д$@`x=��{����G_���������:P����_����>|�x�]��=@��{�s�#���x��XJ:��OS�u�|x<�	IԚ^}g�N������w��&��������Y��Y@,���FN$��I���x���4���M/S�)J��4���������٠=N��;<�ʔ�riz� ��5����=��rh�)JR���~���2 3@܌����?;�y�Ju+�=w����H���z�x���r�#ĽJ=w�|nU�#�9�{��CL4���}�}V>���,m��l&�N�Mt���;r월�nɢ�~�:�eYw@� l��6��*��Ҁ4�[�w�n�d4=I�=΃�<x�ZR��4��y�R�e(��u�(x��4�Ҕ�)C߻�|������)GRRi�׎����)G2��=g�K���8#�۞y�s���o
Q�:�{)JQ�w|���G��R��QԆ���	�;�Wxrh��x�ĥݔ��RhS�#��<sGS���>���/��x�$Ҭ4�$ZLP4�<+܏2��^����/>r��r��{�ߞ9�z���/�۾�|c���̚�Ҕ���x�w��9�'�~��X�%��M�Tq��ZR���п� ~G�?|	�q'�LO�R��Q�CCԚ��N<q�ʔu!��M�Y�R�e(��z�<CԚ��JR���{�<@w�~�(|bD}���fL���m��UStM7W���~��Gܕ�T�e��w�C�M��JR�}s���&���<J]Xn����w�]�wk���k�����O�O�ݾ$�� J��*�c9�`ݕ%'c#*ޠ)�@�@�	�������7X�Z�oU�E��rR��
jm=@Sfȵ���2�T�b��[nA諮m�0�S�\U���e��c!it�(����UUUUM��m�d�  �s
�sc���m�ܪ�UTeJ� 
� f� � � �PU
�B���_�-��۸x
��	]ʪ�.]�g���oK��v�kj�li��;!2�UJS�b��'c�����k��_��G����ZD��Nt��$0č''o�y�H�Oj�B�0�$
'M��a2ZI� Mf��H�	�t/� q x8����D'I��b2����?�X�����m���`6��r'�8�˛^�%�OyU!��,q"��@� 9i��<m�Co�~�>����dc�����D'ą�abܐ�FWgexĭ"N$Hp�ѹ*��bG
>�=�w��#x��Z�/l��+Td�t)�,q#	�@��v����I�䥰n$I���&:���
kH�Q��q����2F	�T�H���=��q���Q⦥v���*	�T m��+����YPba{Ͻ�y��j	`�05�*�B�<2	����>��h�kEh#NDI��$��>��luiZ�F��U���j�]K���c�*�Dn�b�`՚�>�%��e6��+Fa[�c�*}�(��m#M��΁��DN,I���b+�5����	d� ֭��츎F8����Z�QH�V� ��-"x�ʨ%LTlč�$�>(#j2�H��m�y�@r���< �@�g����G!:H�Չ�H�3�g�f'	 x�;�$�D�)�XRl�p�7d�	�&�*����B��oh ���e@ڴ�=���j$�
"���G���W�`��T����>H�'
�����!�x`��sZ֏��v7,��qQ��*m�~゠���4L�x�hz]�H H��_D����o��� $���m�5TmN�j�(��>H���]��$ "8�@U饦8'��h��7L�Dµ+A�RU2�nZ��� ]��m�#ufU�Cx��ܑx� 	 @l����ō$2@ {Gr���DBD��J��˪��
�6I'R'�A$��Q��$T,x�>'����� �������"uRa�R)98�^8{b��$M�mq��z6۲��� ��9c�d��I�
�JM�d�7Fw����$ N=v		x �~��<�)�ZּkЎ�A6R2�U3M��"�����/H(���G����꿉YY���Fhz��ʬ$ ��-�s�<q�G�Z�` 4�0�=�8d�H��D�X��GY��H�Hh-�!i%�(K&�M��E`��נ��`3�v,i"� �Ǯ�'		CD�u#�L�QH�E#T*7T������(�G�$��y#ԍ�onJ�� �B�!!�Cx��߬�� �o�������H��v�q��v�ی���ĭ�ÞK�Sz��bTWRU ݸ%ѧ�[>leؕ��7�H h�Wb��DBE�:� ��'�wyfY"*<HD����g2ȲR�a����m�=�}wČa3��0 ��Z]�w�Y<HFz�Br� "5����
~�� ���͑��?��❳�<Q0��bF4���JJ���L~'d�<HdH��M1Y����T�.�I�Rm��AW�z�\������j
�ペ��H��Q���%�z�}q䞓N�v*�:P+�qč%Ҩ�E��%�m#8�]�Tp�aG�sk�$��%yU!���&�&����� [h [h �-���w6����`8�ꭶ-�lxu�e17(@��5���OL���;�;����G��������+���\��)U5J���1��T����``�n�c{�Wb��Mv6K]��{���ך�@  :���P� �6�m����nѶl�T�P
�mY@
�P��`� �
�UEP-޽m��[n��;
��t��b]������wAu�vB3j�;�B���� �Rʀʽ ҍ�SAj�j�LK�Tx�t���D�1#�c�*��K5�g�1)*��s���u��S�)���,�m���g$NЄaw�*���U����f ����Cr�Ʌz�Ok�K`�H��7�s5�,��:
��Mt!0�k�2$<�0�!^H�i8y�rUL(�W.m{���s��Hv"�(I
�q�g��#z�cyz��8��B!.p�R~�B8�Pxy��
�����ג�I���H�g ��� *!Ȑ�@��y�y�$y'RW]!`p"��@����H@@��~h�T�R�[h���Pq�P�<?k�U�U�r��j��W�U�tX�b 3PS"�tS�_ �@�.�w����*�B@@Ȑ�BمnX�	�@H�C�Hx8�giê�@�I )��$�!�Ǽ��)Dc�֟!�G*qs&�?D!p��Y�VV�ET �,g5��tW���gy�8�$�C"ED9�s6/%� D��$�F��`p"��~��5�봐v�
ۥ�[����ҏ�tĉ1"p�$�U���6\,B@@Ȑ�!l·,`�;#o�3٭�Qq�D QZ>IT|Q0��\���ZD�W�R��X�x��z�ZBqฐ��޹~��4n�@C�$�Fԥ��+�H�B��l5[�p�Y��k �uq�с��Pe��G}}o����K5�g�&%Q�Fg�?���$2$TC�!`�'3b�Y�H�~�g$������\+L��޸,�$8>W`p9i��P�$ā�]I��`�@�D'I��h�@�Z�q�>����`���Kd��S�!8H�J�N5��`�ݪ�UƸ_�>ab�1��c�
�h�Q+궀�x�c\yQ�c\kإ��PHj�v9����uH��1GL\̑G5J�-��1��6mCm���xZ�4 �
��NĮ�����2/�Xz�鵂x�Ρ9���Ģ'8�5U��V��sR��Uwmۖ�F:XWh�5d]j{y/����f�*�<G�L������<���yMr-Q� ����C�τ^kGӾ�OU���F���\����˂ �� �ݼ�ў��'k���]Bw���` 	)�v��!�@�.:���@�<���%6�i$�@ �/0p P x�d,i  wR=�<<I��-#4�ꣅ	%��� �4bRa�H���-�)Q)�,Ā$g���^$44ƌ�@� 1иn�	:������<�ݳam���k�,�w��,����;���SPF2@�UUU+)�B�lx�r�JM}m���a���N4��H` p"��,n��>��t�b��Jc9z��4�Y�&B��@����\��N�ư}����t���[�qݟ���Ι��~�o�-��	@�Y)`B�����>����Ѝ�Q������F��4O.Y�!�>��`�$�&Jd��!�M�"�蟔�LvO�Y��=w5?!�m�;~���$$�AM})�d�m�	/j�����]�>P��x����זm�ηY_�}� }�Yj�Mʛx�{� @ Y�hVS��6�� [�F�  �xl@�*U)���� U�/TM��O=m�U�  �Ѯ�V5Qm�=��Px6ǀ`k�=R��<�K�< <S���n� �=V���lT���� P����� � uUp�� <y䡦����^��(8�W�D�K�Vx��M$q�2�׻�x   ����u��u�����SڗV<s�wa�.�T�yT �n&��wz���	�*	Ӏ�k���M��۴�g��aGP:]���/+D]T���uP�_��}�o�ͰU�-r�Ҭ��9��S��0\�Z��^��^�	�m������.��Ԭ����5/6X�h�c��
�v"�rҋ1�y�5�鸐/G:L���gDUUR�<XN���Z�t��$MC�T���AV��H��P�*
�U lf"�]�*ط#N�Z�.9j�Hvܣ�j��aԼ�c��vx]˗+���.]	!,����		H��[=v�vʰL�W��Ь��MO���|%�V�~�[����`�UAe;�r���5Pj�        U Un��*���eӺ�TlX� Uz���      �kjJ����x  ��ScmQT
�p�u��f ��ܕ*g�ր  �    �     9��|    x         U*��*�S`p [�TU   ���U  ɶ *���     s]@   TU�*��     U �|       6� ` p � u!S��Ql�aS6��A�0 S�j���ʪ���*�$  Pë�M�*��ڍ�k  �Ͷ�  U �-�oul���T� Y���.�ː�'�;
�W@U[��r���Sv�OIn��~��<Ƿpl$�D$6>0�)�P��d�ͱJ�B�;+��.r�Yҝ5���]�ݣBf���u��ri��`zZn��n�wvT l�+(���U���s����6��6��*���� *�U �   � �l�'ZUƪ�,�vi�`"iV5I[pW+qnv8Y.�U�qlm�0c�=�/T�� �l�[X���A�>��[uد����w�_��ʱD{U�}1;�;�F/W���i1�j�;���a�T(ld���C�.@�\!�"~S=1�?QFB{���?!��Rڰ��^ŷ�W�>���BJ[]	Jqk��f��_d<���z�\�D!�r)��"?a��������AQ���a)�|������V(�՞S��'b���3U���e��Yh�00,k�֑^U�ُڄ?x��p�ԉ�L������2��\5hqv���mʥA$����jn������]�]� �L�l ll�.�n	�	�tEl>`���AX ��ru�p(k���G�>2S�A����&h�l2�.�\�7Ӭ�u�o��|��<dsj����ny;F�q��+�逩BA�,�Y���^j�۬x��|��B�ʸE��^]��쵬z�knι6�8� [m�6PW�Y�+òY�/�8��f���AX ��>N�\�ؗ��<�ŷ�M�� 2s�v�sP�u�u�u���H���w{��v)���Km����6F��^�g0�n��qU�[m��  
�j���a�Y]4�qx��1�Y��"�ʅ�"�FO�^�!ٺ�L��.��ދ�h���V[j�R�z�h��z^k����郎O���,�v8�<|w��,��v-jכ]9V,)T���x�t�� ȇ���j}P�]-xm�ن��Ǫ;��G��ZBj���D0.��5��ns>ٓsI�����ͫ�n������c���@M�2���{oT �[u&:W�PW��=��*q�0w��u1�d�U�#m���^6NU�AҀ�=����5҆�J*����?Sogt�zt,-�[t�Y���^k�^��X�ѼU�J~�2!�v�\#�q�S��m�Z���]m��f�Y
 2�P���<z9��dt^7�'c����Q���vmǻp���T�J�nV�H5^�&U�
e\"�tO�S=1�"a�:Ğur'�!}�o�\4D>�{��2���#��-k�_^��i��B}C���F$�>�Y��ys/�!8�Oz�����Rd��%��ݑ�l��z��)hB0�Ȝ4D>�3�;�r�%T�u4��Ѧ����B���:&�v��׻�s{�����@إYYZ�m��3��+R*Y��9�L��R�����p�����݇bּ���і�)ik���p��-�sK��ǡbS�PD!����"�X�
s�D8^��g��B�@,t�5�ɻ<K��}��l��܆�O�a�58Y�{_s��k\z�{�R>k#����,"�;.�\d��P��&Z�L�ܕ��3�����Y�����  N�
܋ք#O�[�w�n����V!a�����ɑ�C=V(���q)QYB��P
�]+��2�`U�#��Y����* �g]��w�v��� i��0�)HN��1���!����1g-�`xyr����;�$�����n����B�U�3T��v�`Ip�ʎ8NwN���`  m���mR�*��=��k�4�l���[%e<6¨ *�p1� ;� �*���U
��v�ƫoK��(MO�X�ĝ�8�)ˎ�6���Ag���G�N�ml��/��@��v���45�����j�g**KU���8�B�7!�ɑ�x�1�Z�N}=���"v�]v�E#��Z�Տou��*
�QR)��D�T���9�s�2ܓm�F���I%��
�PxVӝ�_B�AZ.��W#yf��=���d3�����֙G{�%H��A����B<���ly�v%�Ԉteg\�g�>��I�|�"�eRm"�4*�;*��~�=�ړR���ɏ���e��U�n@���c��[nlm���;h6��m��*���ȽP�E�`����Sd����Oe�/iN����n��F��<��'�7򒬌E����+}�/s���m�k������iw5"�Ǌ�]ȬV�UoJ��rB
�"e=�k�rc�Do+�0{�X�2,���Wj�槞U_�=3�u���� l +cB�xG��:U�.�rf����8F��ήrdqn�OU�*#��R��6T���JZ��qcC]��=[E��i��\�z�Q�=j	"N�dq���fA�}zGA�IK-V�ln{Dv��3�8�7�mUw*��� ��J���� �1��[mRs��Ʊ�c
��9Q�����0��x�v+�E�h����Z+g�0�e�(�I�I ��U�[��{�\+�#�{�Wk�<^�L�$B!�9��F�*�F��[�v��h�
N+Y��L[�dY��rc���ێ���X�\���ղ����Z�P�L(��i�b��[j�S�m���\��D�#̮0���zv:��<w{Ц�I:- Wx������W�^4d�֢s�BOU�k�e�I����7�������i�U���G\�8.��F1f�A�P(�UR�� �B[�㤖��I�aA^fN�,kϸ�|�FŸ��/O�<v�M���NE�wy��XH�ٛ�#�@��eh���j��#��K�6��Z\Km����!��-#̮0���?l')�jB��Y,q��5�5�~��{'5�-=B���t�c���U���/�Ϥ���'�#�V[mmIKŭk��ry��m��_j��FŇ��"������xO�~��8ܨ�,M�b�!�p��_B5�R���(7,B!d-.TW�����2�Mm�0D�Ã�����"d�ˎ$N±�K��j��IeZ����$���P��
�lvU�n��M���c� ;�{��}#Q�-����R���2�[$�JKk]�{LPI~ڞ�'�06S��I&Р����b>W�R����{çR��GT 
$p	6m�˦�9�f��w^^��v��ử�?>^�}0C���-"H�d�(Ƽ߽�)�rd�%�6�i�	/��E���;�+���N��(ԎX6%s[K��JKu:+�`���c�w{�燘ߞ89��ί�<�,�o �&\(�%�(ƴ��D+X[p�UR615t���{zނ��[���  ��<U ��;��*��ة�lͰJlP�P   6��N ` xJ�T�l��?��ª�� �����C�e\8y�e�tk��w�&�O�A�T���[����5l�D�i��M��	߽*m�C״|�k�(ɞIIk���`H��� ���-4U�rAN쳡�w]ދ�e������j&�tRm��8!Ѿ�6��^�̧-�ӻ)��]�T�����I��n��m®�+�vߘ���X����DA-2Bl��d��G���n����]�^�O��g=�4�a`J�i6M�:����k��$BҮԂqR���U*�V��-�Ӗ�E�C���	�����Z���7n=մal������n�������]l¯�W�m�!���fmH�Ć�[$���0f��Z�foB�!��Y�����d�I4��Dٞ������X�yi�ák�o�g�� ���
�a�=�/����̫Vd���/�>��4����(|�II���[.��ѼB��q�]���UGpN�+"�h*�US��9c��g2������W��'�B�i��b�ŧ�k���35�r|�u���_єe���]!Rg�gy��}۵n����/�R����p}��Q$�4�E�RMBސ��^3!����������X#�   ���Z��"�z��$tW��7�~���7mx��@Y*�^��\~}S*��A��}p��,֟�fO�<�縱��f�*�lP��V�iD�3}��4Fbv�O��G�9��vt}pE��Zf��I"�&�"R@#Fx;l�/.H�Wd�f����2l�
� 6�6��فT��wU��^�O���P���)��pN��W\>�QIΕ�p}����b�9�/�u�h6�D$�m&�j�C�h�ԇ,���O+�E,2�p/��Qմএ�|2]�D�B�m$�������FB_C{��4Fbv�k7��C�ݨ�tݝr"�:�DRe����R��C�p}���R�
l�����T�'5{��x6Q	�����mfC�����u{W��Öt|��W��XeIľA[���0�R9�Bj�=��`�n�W��۸���Wm`�����3y��w��T�T�Ve��?"&���X~���3��=���?fl�2(��]USa0�7f��/�RҼ!��V�F]��6g��؇���D!h��M��%��_`^�W]!R]|�c�&3������_�EyM�$���M4�I�	U��
:�pRG�>6��A���.X��
�,)��0�i$�(�n�C�qWR|�r�<)��G�V�*Y�*��`���m�	U��"P��1��[�  �`lU�s�m�%[T͠��a8ۀ{�՞v�z��w��j�<n���ݩI��S�>�2�UuUP�Jb�G���dc��n�t���AT��4���`ʻ� @, QWTʨ*�-���Ws���m��T�UT �p �� ��` ;��UUJ�-�ͼ���l/T*�!;J��pV�cc�ݫN08P4��[JKUw+ ��������ﵷ�6M"�n�Q<�?G�~����*���ƳyT�Y/��d3c8D�����xX�̉�Y��R�W�Gf,��H�VV�p�֜0�7��"!hp�4V��I1I$I6����
�Á�.�U���N*�
�QRs��ɍcWl�W��bb�E��XT��,V°̱���A� ����0��<��xE�gz�[��YP�l-�Zu���>ku�ӊ�?����Duu.��(yL�b����~~ґh��������('+��"���U���� `�)Q�m��{�(��E�m�h'z3��)b��/�]��l�U�ć���g��VP��KKkn�{'�cDx����F�yo��b�"#��;�5�x��w���r(��Pe��`��^�dYʐq4d0T�}��>ꓨ���C�I�y�h��B��U�i9wWnt�e���to<����Ͻ�R;�50���-V�,r{}݇�5�'ģſ+�Y�W��3(X�ǎ���\��B0>���W�!sHC6�U�fJ�5l�(�iGQǰ��b�T�)�B��-������!�u�}�yw�"��&8�Uˈ���Y�Yc�(s'������F��
�XsZEZ����b>!h7%�U����>*�p\��X����H�+���e��i4ʺ��P�R�AV�����2�fE^]�s(X�ǎ��^�IX�  ���7e�ּ���ڮ*�[Xc�*�6��]Al�j
�s���z�\[> j�R����i�~�,�+s�\!�j�\̿���j�}׼V��s��AxT�$�Ir��WmYcc���v���]�܊��Um�&���������Q�[��%� �]�1��w_aWP[*��-h���CyT��V$+
�;č�۬,d�ZR�����X��Ӓ*������ط�X�:l��6rw��K2�+����mn�)y�xEⱲ�᭻R��rz��cr���6B�r�����w˒�h�uJ�n�m���{���V<|d�=WJ��@uG���ě�dW��RI9zEi`I ����93!��=1�г���;�? 0��*��f�ҧ���� ��Z\��EQ�P��;�g�9\q��s ��~�
�JNwkm��v^�xנ�c���%K���x�l�?D8knԸE�ܞ�1Xܿ����/�$�qF8IT-$�|�C�Y��cֺ/b𞘪�g���'�����@.>r��{��`��ɐE6I:��� C�z���]�����,Ä>��*�O�7�+��l��5?\���!QZ�
�q!����d�w�ȅ�|Y�/���@C��ٗ��!����n�&�- �rJ�s��=|il+���x��p�>0��xK���iAx{�x��q�*�f.@I-$���-�S�M�f���J�R�T�i�d�ecN�2�tY��<{m��q�tL=kj ���ˤ� /^W��ޝ|�� <�X��ۜnA�U�*4-��H�r�.x�D˱�Sp�F�-!M�=�@��� ��w�  p
�ɲ�p�l�P6ʪ��K2�*����  � ��
���z��޺�0���7X����7Ob6���xX��+��T�PWR�+$�*�~GξV��$Mi�%;��Z����^}�-}sW�\"�w'��*���|G\�b�D����ߛ��0 ��Y�u�����~ �(��C�T5WQKW.}8���dK^S�����ж;i|E�ܞ�1Xܿ������y<^q�ssy�-�v]3�f�ij�h`2�@�mNv���}.f�������b�s/y�m�������W(�FP�-�JSb�D��÷�J���{Up�2�g����N��᪺�Z����r��m�SR VEƑ�n1�ۈ�5Xݳ�G ʴ�j��誓���u'u3���@�o"�|�K�Q�Y���7/�|a�½O��A���!������VRH;,l�8����5oo��z^"��/�)�=B�4f�ȓ���I 	I����%��Q?y��Q���E�#���"�������dc(e�j�?��ߋuܶ��xM˞�tK�y�W�%U4�D���t���t�q��Kۜ���}g��ˤ�H�%$PAB�]�!�K��ch9&A�U[]� ml�̍�zҡۉ��mU1&c����X{�et�U����Q�/pI{q'����%�r+n�黢�j˾��3{���w/o��(7.\�ڀ��#m� eL��s5�st�79.��䖪9!\nsרD	����$��4U=�<�0O.oU�^�#������r�>��ߏozI`?�u�*#Os�M����kR�^�۸����Y��L�����U̯D�<��ŃK���	n3F59x�w`�f�m��3���!\��HR�����~�}���_�ϴ�5X�
��s�+2x��cF	һ.�a�lK�A��%V�sϯ�9>dw����[��t>���Y��+�ҹ�U��\�M� 2�I������q�2�eu�X�cj:��e�Uu�z��u�MV��`$r�h���Tj��[������6a��/�_�~5X���pd�wTƌ�X�G),�J*qfÐؔ�;/O��k��@C⠹꿛[��t>���z�]zY6�	luI�ʣNr�;p��{ :Yi��gg^qd6ٮ��h݃��"  +��̇b_>oz����5p~��6ts���O�S�.y����f��o� I�$hd�D���ުe-��i�be��~;��;�/ƫ����xv_�@!@���I �)�z>�F	Ӳ�qv_�ν>?]��dW���'��������`K�Z:�H����_��-�r~@a�)8~ز.����Ύ|ǲt�D��r��pd��))y�?Ǔ���O������Y�ZJL��������V	_W)��f�9���m*0��@�v�   �T@U1��J�U-��l�T 
�ت'Z��v6 *�uT�<�l���m{jz UD:�m�U����3� �� <o%D곯U�{�X`#��-�s*���������w  �Ytx8T���  �T=�឴��V$չK���.�p�V��|���)P�1%��{-  W�-щg]Ṹ '�@󺺶�r6Þ����+1���{�6Ŗ�m7T�r�[wh6�x=T�������k�aq�dv�[RX|��mԆ�un�½]�턭*���U�sڵ�K�tR���i�f�s8�#r�i+�$z���^��1�M����O-��=���q��"�;��\q�1�yG�X��e�N�薫@�7b%X�7b��U,�u�0*Zts_���Z���n��n/a���w�wnîCʳg�t��Nz�z�]���'��v��y�'4�L���\��sV�4��{6� k�F;F�Vι�N%˷vʫ� m��*��Ѷ�Sl;�z��dyg��oG_�� U           �46�*6�TN �csTxq @  U *�Vڠ���� �M��@ �[%V�P�
�1y��R����w�  
�        �
��P    �    �   *P *��[hT��eU   r�@�� UP+( `   �    ����]H*T     U     p�   � l l� �� -��U6�6ǀ T�T�UT�; j�X�)�wQAf*   �[[��
���* 	��T   ���s�m�D`
�� *�ĠT�A����'gj�W�nF�
�˞����CL混=%�Z��<�xl\���vYmS6pNU����Uj�;�6޶
�!�S�9j�:ۅ'��Y��Gv�uTK�[k�߻�ow�  
��ƶA� Wd�ɲ���6�ݶ*��*�6�T+nJ 6��NUmT �U)q]�6m�� �5U�k��*���2+d��֝˔^�n�%.1 )S*մ��2�c[ �X�TGI�Q�g�����������'Nˮ�ƨ�s�C���]���D���l�n� ea!hƀ��_�=���c��f��-\�� 0���?CݞG5o������J�� �ub�"ĩuzY�Ɔi5����O7�?��Z1kR�e��~�
�D�,�E��d���U��l7�u2x��cF	Ӳ�qv_�ν>���]�W&�A�m��'>ؖ�����Z�U�$9�������U}���z�l5��϶�퐡
[D�ז��s���]Dֶ�x�n�o`;��S0	P��;�1<c�\��y�S,mGl8˅����C<.���у���uzK�HH!��)$R�w.	�8��М�c�X��|{���ݤ���슻]$�%�m
{~��g��"�U��Wr�Ww����)]֕�^�Ӵ��S.���N���E����%�Λ::\��cN ,.p^�~��3I��>:)٤5$l�T�E�F��5��i�bm���eq�5V#����s��>}{��-�l�dRe��5�I��*�����`�%Jt�vVA�u ;��F�A� JY���JL��|��X$�w�6]p�+���V��Lw�>0��T�i%T�VDF�K�9ȗ^oJ�p��<�KΛ<9���3Q -���1��'�~�em�9h *�|�!�q��a�,<�ICeE�Q������{'���ݥI�m�!I�U�^9�쭆��TL6�1�g*O'�~�J�o�g�Y��G� �$n�C�W�����󼟖�M���r⠻�Y���cbf� �uVޮ��Jl�9�v:�(�.zr��*/bj�i첫UT�*�Q��r`9�,+D�<�����=?.>��/��b��Ė<~=�U|S_ދ�A�$ j꽧T�¯��Ӯ��l-8*�|�(�LP^C�X[�Ň%!#� �N~��z^M����@��*��*�@�,j�P9�/�澋1��"������q}��=@X�.����n�W��g٪�>Y��i�ſq!��n��m��$� d���r�_
��0=�ֻO�����K����蓚�|ך	�rH�^�� �����S����1�V	6�;��6��U
�L���9�iyt���[���%���-���S,�vȘ;�Uȟ���)T�#qn)��5E*��StPTÿ������=@X�.�)x����?U���+��z����
� �������g�&��d1|&���x�LN�D�.�f��+�6�;,�j���a�k�t�[��� ���(�'�Tw;�Ț;�����e�=n��-u���� ��p]+��v��'y�}�x>�se� �� 
�{VoE��J���ZH��D4UU�qh+`�����l�����cl.{[��f�8l��
���.y��#�Z��M�,Z6i�D��{b}��T4#K�P�H�P lwM�
� �\�UM��U<l��U  
��   p� 6� w ]�*�6�k�ٰVU�c���7�V�U���Gg�tGl��W'�9X�6���[��8*��e�h[I2}�'�����n󏀾}�}�v���R���)2)�{�W2�D* ��L����;��u�]�������: b��͝����a�7*��#���8)n����
���pUb3`���H�	$*%ޡ���o*�m)��.��C"v�#�9d��7��I��>i��@"
e�p�w��n��u��r�lv{��X��=��%�T�(��E$i�`�]��6�v��n �<�Z�M�QPU������ah�`:k�??>���Ut���J��}!v$�D��u��P��	"�e�I�A*r/P�<{:-�#='V���X�G��r>�!�M�d��%���r����x��[�6'^�6w��ُ��A���D&KI�j�R��o>
d��is�m�����b�3��|w�˶�\�)@��Xؼx��w���x�H+���>�B#\x�0M����"G*&�j��`&H��3���:�R�ci݃jXi &��m��eb)vA�Xv�TQM �۸0Tq�Hp]K�WP}��خ�V���=4Uٹ`����!$�EPm���wX�7��@�;�8}��j��b�|�������fP�42�D6��N��3�'�ؽk��+r\,�����q�ϗ���O?=�7k��  󒣜����=��`�q�ۦ��s֏��ww{Ź�y����G�� Ul V[�J�>l�3�
B�c+��7�GH�+��D,����Ы����\��L�@��S�8��â< ����o2�]J����UI�T6�z�������W�*�֊c�Ƕ��l8>b���?�`�~Ƽ���vǉ; d�i$�7�GExi��v*|:|�G�*� z>�62�E!�[r$PT˦[m�J�����Cؽ/O��j�%�����dW�R�7�tvH��?jନހ�$�Z�[�����g,<��Xv��cH���h����d�d.c��'R)�D�M�ؠP��8�X��������펠�Z��&�!���:y��pF�B�����m�guUm� �T���`��s(4�"�ո���Fz.�签�����5�'�~wf��a$�$uJ�����r���w6��ܼ��=�k�}+�Jƫv�K)
�(m��1���o��Z'���!Aǫv����]�h�K$)�,���;�b3�x�m�ݯ�{�Ξ�m�D��+�@ -Ylp�ޭ.���8y�����Ϝ�}��UT�J�Ԭ�J�A\��N��ʬi�U����M¡T��s.��u�m������	�$�;�㡏\K�\�g��mZE��<��t���.����m��*�F�����δ��V����S�H��gv��s{@ ��*���AUTm��Ue*��p`�T���[%ͮ��P�  Wu qT)m�?l޹�
�����;��TpT������=U�^��Y�Mu���-ր�� ��F�|[V�JӷOܳ��S�۩*䙵+����s!���[��` 8�u�5�5;�����+C:|_I�ɚ#[�:�`����B�8Т�h�d�w�28�]g���Zh���D,�_-֕��h��%���i���#�T�5�萙N�it���^4C!�N<.��x)
у���C�;h�>�9:�G5��>���Ә�����}�6��7�
���캁o���ߏ���U�g#�+Ӳ��9����;��#)����;��pU�^��J�B���a�}��W3y�V���_��gy����������di�.F�)�l&R	6�L����t��2,<p��!�d>2���5[!z)
с�eU%���M$H�|N# ��Gr��<0�"�Q7�_�1ՙ��^h~y�w�J�#$�Ri�@����kS�9���&p�ϧد�צn���Zv������r�u���<67o/4OoZ��KRU�}�4$Gl *�rH���[Ŷv���2��� -օP n�j�TlcL���m����ϝ���?b>nj*c�P`����V����G��cfRK	m��D�
f�E3��������0�������HO�^Mc�.,���'�swm�Ų2�B2H��`W|���+Ex>��z(|�	9׾��>��&4�x���7��hk7�;mq�6X�T�澿�`��x)
у���[��2wO��{�� ���[
V�{>��s:z9���b3�v�����zwy+I6�a�2�+�:�Hel��J�q��e�m�ت��ͨ�6E9b�.�upd
KH2 �����צOc�\�ܝ�]nm���yu��SA��,U
m��Q[,���S����qn{@�����zs;�z�T�7j$��жG(zn�;:lk��z=Žײ��G���c�~��ں� kj�;�8�s6���v(c���2X�Ks}Y�BI(�!&�i*��l�͊Ի�}]��OJ7玑�ux��%4�`Rm����� ;�s˲�ˊ����8 M%���V�D�H~_/��\$)ǲ��ե'of8o���-��j�s4�F���J�����]�?Y��gJ��-��K\��7K��Ca.@�(�[m�I���˂���ל:�m�݈�v�}�s}��(*�D��,�P,k��y1<��qBG��������\>��s�VǶ)���0 �S�R��i������:焫���o9o�9�'cm�� �+u��Y�҃)vX��+��M��56q\�/n�� ����+�x'z�*�m�ݯ]m5U����^eʣz�Y�����{/]!hۉ�%UmT�Pލ@��>R��k8i�)\�Α��J� ����[@w)�U&��{���;��m��
�Lȋ�*��   �U xJ��UUm����JZ� N�UI�����;�8�m��z�٭��/[��@�U �fٱ�z�~�y6�%CA��w.�\ў��7R=͕3e��X��}O��L3�I2��m�A*7�LT7��y�K��|x�d*㽉��x�6��0��yw�	�n�B�K���և���=cy;L�#c�||~�[,�����gl����~�lq��mAG$����A�ڝi^��AZ�����,�SE�6s�c�֙B��R��ԥ����P�������hkϯ�-����tD��>��;�,Tk�;�[%�%��0��r�*�
\3���=��Y��]��{ �m�
�"�� ˥L�l��B�n��a���|�-��O_F�J��θ�+�RDK���2�L�E��sJE&�bz\;B���Zu* ��l��mMl���N�9Z���r��=%���26�ب0A��Ȕ�G�� ��=�k�+{��?���}1X�3��잱���#��^>��!��������%-$h�9ֺ*U�W�fB���vpb���J�,T��u�އ!���L6�i P��ڥ��9����nz�6�Q� F�Uj�VP�mm�i�k�i�����Y�^*	�o/ZdY#���ɍޢ�S���_�FB�|G���d4�L6�vU۱P`��:����AX=/����X���B��V7��6�k��Y�E%�s_^��ˋ&GxG����Ep����fe������,����5�y��^��c��)�B�f�B�i��xӨ*�=�����L�c��0��c��C#����{PJ��ag5���7�_t�v`�E󜻰:;���𹇹�-S�n�R�m�.��-&��8�а]�x��3JN�/e�j�pU �m�g[ݳ�II[L�v��?w>���g<�/��Snԉ��vH��8D�V��i�t���lR��vk^|Zl1־Ŝ���A�"�9�������#�X�#^�k�K�o}#��m���$h���28�����&hEz�n$|Dp�G}"����Df�Ų�"�E'�  1UqkC֮���_�w���=\�D!ڮ������P���h&����$�RRIH�d�h�X7�U�L�F��Ya��[�=�:��A^�&'^�0�X+Wy$��_��������7̼ɗk�������; �U)3jj� ^�4E�z,Z[��w����8u��>���Ӛ�j�3Q(3���dY�/G}"�w/B��lRR@����}�Ϧk}�V!�*t����ɑ�Hr��!w]�zT�>�i���E*�*�"��U%^��8#ò2''�Daz\�7\k����ڈIA-�e��}�������t78+޾÷2�Ry�Ecq��#�����BH�R�'���}��d�Do+��Lubf[%�����y���Zֹ�fN��ZI  w�	��w�ֵz�v�Pئ������� ��,*�����hՌP[[3�3�ԼQ�P�YU5�b�|�(��ùh��E1��^Ѱ�����enwT��&b�_���^��ޯݙ  +�T ��  N���\���m�� *�@ ��  
��U� � �T�keC������6 ��ˬ��r�I�����:��y��5;�*�CJR�uR��/T	d���keL*�w�#��˄[R'���d�Y#_.��D��#O��,23��v����Im���AH�G�׭b�y1�{��G�>�����!f���y��V#�}g&b%Ȱ�d��v�;vD>"��z;�!�tOd�Do+� >���E�El��o+�|���|��Un��)KJ@��NkZ��ì�J�G����`�p�jE��s�d�[]k���vu�k�������ʤ-N�2;��h�K�G@g����\W�q^�1�h�����>��zݐ ";%qʎ�*��ڧTJ����l�3U]I�F��U@��v�^�=���вR�5����P�Ӎc�\kx��w�x�FD���#�^)��b=kE��ml����2s��Vd��B���z��#�q��L�CjE��s�d�Y#d�*)�%M�M�j�E�!����[��bT�ЍKLg/yiE��|G����
�Km*v��h��74�Y�<WJU�v~�4��XD?R'�X�7ӟ@���$��HR�c��8����j�j�-#J0f9p�G����E|E��Q�e�-��<��R-�UL"�n��1�q�4�-���ې:�ce<iXډ1�Z����B7Q�cf�T
�SX9�'%8_v�r�$����帵o'�����&[+���R� �U��'�B��ng��)�])V�8��"h3�_D�F�{THf���i$I��Q��A�fbfZ$�cy_��eu�!@���]����"k�����9�[[���sX��'��s*��<F��*�D��#O�r�Dg/rz,J�#��o��j�Caim �,�͝�6/�Ǧx�w@��D8V����ԉ�t�}����&��,���]�)U�EQ�וQ�r����I6�-����]Yl��2��� �.m��ϋ�7fo��7�O�L/zԱ�zӋH�����
��q]qȠR�)i#D�9϶ִ�W�W�R'���(X��p��OU\��B4�G��ز.�ĩS�TEm�j�Q�k�_^j{�l�a�滭�8a�^+�'謈p���[R'��؏�i|�	 Yl�l�vn�`�-z+�(F�.z{}������mOYD�����h���ۗ;1Wx�J���C���1\"�H�)��ňY�}�?(F��{F�IRh�Er-bUڷj� ]b����
����p�E6
�;	��W���ƦtYe�p�j|M��p��؃��XG�80�/���VD8ow�_jt�������n����}�b|F�����B0خ�p�:/l��5FcLۯ緸���	
mt�;��8���\>0��]��*�/0��/�.ԉ����'��h�����Ie [SD�y��kϸ���dlSSr#�;�Y��D��_5է!�^�Ϧ��G��Q����
0�"�!��s�CjD�W#+r�C��S��w�<P�6+�\,��ڳ�w��ݒ��  $  Z��*�leT� e*� �P *lR�UUT�T�Mf��l[ ��� :���u!�B��eZRL�Z�m*�a^Vvr�m� �"p(`�
�0� �����T6%��`�
�u]� [ Q�  Vڪ U*��^�� n�u[\���ɩ�йP���N���g�YIys�g�� ���z��-��X��p 
�Sj�͚6�+���yM��{�cx��Up~����]%�p������rݞ�骮(�l�T8� ��Z�wyG������O /K*�8qH�t���
�%��G��
]��ܞUx]*��T���g [��D�"qh��Z �z�]j��׈b�Fg&�=�,(������V�1^�X#@���&��3���v��m4]����od���[ ]UW*���.RP -��,n9�x�61��l[=C:���T�K�c�nWժ��۱�k��B��&WJj���� Ը�&��ܧ-qke,���G&N6xըYf�*i4m��n���n��7]� =�]U]����F��t���`*�         
�Vųkp�  �w��5P.ZP� ��  P  ��@��me  �m��f�,ڥePT�r����sJ����  <     
�   � mT     �  �     *�*�@���� lL�    ��l�` T���    ��  ' c;��� �pUU    
�P      P T � � � uP�t��6�Cl �K�� ۚ��oq7�b��H    ��M@��+u�@ � 
�
�UPt�n�;�|/�tT M�����ݱU^����1��=T[!R��8�(��5W[n�]j4��*T	��8�W]ӤUy�+�ɱ:��氪�n�Me��j�M`c���{97�g�6�V;�H�[[��]�զR�  ��UR���[UB����m�� 6ʪ����d l� �� ��
��
�f��@ ۻZ�Ъܥ�����rȋhԞryW6�׻��vB�As ��X jT	\�0i��L:TP7°xx=�z�q�/����ˇ�����Ey��Mтb�E�݇��7�%��r�([l-�Ŭz�����_D��nEt�6,��������&&:/x'��/*���n���]��x�w@���!÷3ήmH���J�.�>0��\O����F�}�G>��5Ғ0)`���5�;���ԋ�!�޵,t^���;ܸl�=����W�a��/4P�j�i6�UU$�4�Ћ��<^��B�,Ä>�yUȟ�#O��.#g�"�'�sW�{~�����
�d�Z��y7�wUcf3����#*�q]ږ� �ګ��iw�[X"�� �nYś;�l���j8��V;�O�Y����w��OUv�}�*�ׯ�f�'\��@奡]%SW�<P�6+�\,��ڽ��9F)��:+�qi)�|a��U��WY[��o>��Z��5=��H�R'���(X��p��$���}�x�|k^�3����-�)d��k���w��j2�Cv�XG�8aX�$�\�s��)=������UT����w��:Q������e��-�8^�b�"�+�RQ�[$�N�}.;��beY�����;�w@��@m��U�ഗZ�C�����T�0�+���r�C�тb�C2,���,B�8C�'�Ƚ��|𚃰��ii5�}�nk���k]z�TL�ݩ�N�F;�O��ZO���]�����p	�j�ӺB�r�+�8`�]0������Sz�1Z/�ev"Ç���Gi6H6�uT�ڑi̬��E���/yB!�V�S*�ȳ�z}ba��ާ�Ke%�+�����ןuʧ#b�]7(�.�a����t^�6|�U5��\�L� dM�~�%�]�+`j�A[uj;���`*h �R���5R���F��s���mF�^;������c;Ltw$[/�^Ě��X�[I&��l,�Y��k}���z����ٸ`�0����_�4ia_�D�)�;sjKJKq�2�^�-�u�NG�(�^�v��Q6X%6-��!:iˏ��K�����V�EBi�~՛�K� �`A��f�/A�5�|1�뵺���,����������ڠ�Xi	tv�ŷ� �l�	�i 쭪w  ����ou��|
m"�M�T���V\��/O5RZR+�[ɹ�n��ްk�(�h� � �m�ȥ/��e���]F=U��ogR�q����1����
ҧ"�����G�og�2V�6 V�U��'d�Y�z�C��!�$W�Q}�,9|l����F�	�:)��T($��~�]��fB�r��X��p��O*��_a���F�5{9S�Ȭ�#���Ds�>?�ĺU���/�*�񇈼V6z
��Q��7�t9�q�K�-߾ah   ^YZ��@��
���J��Vr+�͋dp��/w�o.{ �s��玌Q���j쉝we�m�"��j��gg�V���N�&뤅;�܈J���[v��s�1�k�ݶ�~�⽯\�@ VU
�6�n�s �S�����6��UT�P � ��P�����U�6� � ��U@
�m�݊ . 
zĪ�m=��I��BS��g\L����Cq%R�����eej�gm��p��t��n���n����/Ƚ�}y}e��.*�/��`�}u����h��������}x��yl��w'�~.�	�|E��^V��bx�����+?xN��0M Qd2�i��и0T>żnA��x�C����\��T��k�^�j��O����v��KJH �f��R�NE{θX������:��,}x^М��"���%S0�m�J;�3!�HU�pX�5U�-�������n��n�1�E>���M��T���"�펙n���m��������� N
�[eG�m��e���`ә�����Ś����ǩӿ���J3��ِ��WS�^?ޛ���-������%�~�G>�j�;�Qe@Oo�p��=?C�~���u��ׇ�'���R$�a�J&��ڗ��fC@U�pX�����������[�̔�0i�[���t��,�"C�'�E�_a��֘~�Yg����9�X�U���_oV��i�n���"e\�׏�^�U�d�!�n/y���r�U��6x�b��M�~������A����`F�k���O������	�ڝ��ڧp�]�mr݉`;�I(���
�:�s�^Y����������~:���å�s��`+�7����KI�� �j��C�7��V&+<t��3�"�����kL?_,�*/S�����6�Im#F�
AUW�fC�Q]N|��e��^�֠b���w���\�W�녈,V��� �� ��H�a���]=���n���>9\���W/�В���<\k^��"�m��q�wg�~e�7�������xS�݊�g�S]�ֽ�})ݶ۶� V�H �6O<;�Ph61i�rU^�]��d1l�ofʒ��q�^��Q�����>9C��V:+�q}aT�<E��ҍ���4(;1�����ɇ�.H��m��N؆�6B�z;���}��MpЭ��9R�AV&��ReC�ۦ�$�����A�|x�{/�͇u}.�������ץ̫����y���3پmb�V�@���fϼgf��.�b�&q��o�����x���:dy�t��񢂤�l��E�M����z�JU��6a���ye��X���dl[��x��>;�����i�*���a`*�q��O����&�viP�`�
�[j���o=��+%�Z��C���O�j��1��]�#���|]'��k�<^��V!o_�f�G���7`B֨����t5��M]�5Y�g(p]*�q�!r�讧*�zvkI��I�Mҿq���f5pU���.r+|�0�b򗼫�.vK���n&�А%J�ж���l��<}{�9�Y��5P�θ0AY�t>�~�U�Bu`�*��_����ƛ-���Jj���8C�'��D���}q�l^�];kBfƑf=B2�lW�����7��U:ز�� �l����X��WR�(R��;6�3�S�n��;���7(�,p��mE倫�l�vv�j^Z�t�=��j��c��h�x�]u�G�8�PMQg6ݻm'M��
W+�؇�w`$6  
�P
�� <0n\��Q��wm�U*T
�� VP��*����` ;��U���m��m�j���@hjX�10�펤�`.�2a�[6��L54��*�������e�R�0�?�+�ڭ�E�_�\�s_�����.���3ήmH��En;3��Cq�^�Vm�E�,�Y��t�X���ep�:u&�1�\�Xo��L��
�B0���UPM.��3�ۯM�E�JF�˪���n.����G���������A��[B���x�g��C��"�X��y���ގ�mH���X�v~��Ț�(Q�I�P(���l>�_�gw�ƽ���(f����[r�CxT5��u�wσ���~Jʫ&m�\�eN68����z����խ��]�,�ᶠ�mUj��E&E-�i�I:T�9?ap�1\"�H�/91Y?Q��'3"W"v�?\�|���}��޶ӑ�փ��l�~��P�OU��y_,?e8���V;�^D<~�[Ʈڑ<R�CE	�A�K	����z]s��!n�%�ȑ{W��$X�!���[���g�����hs_\#�U��/"D8n��.�D�L��d�Y�|̉\���30�B��N5iK
Z[9��f�����ֺ���)�bE�*�a��#<�wzW������s�L� �(�-�aY��T֋c&�������w
l 0U*�Ow@�ӝ��a������=Uҕn]��>#cR�*��n�%��轫�x���0�r&
����UM**�����CH\�K��a����Ȱ�j�M����?%��P�г�����(0 �JNfN�c��3�(>�a�yӸ>ʯs�n���J���H����|a��e�]$Yi�l�KD�"�+�p}�C���_�Hs�a6&]��?l�i���q}S%��/��1D*�[���k�׏����ծ��g_?3�/���*	��̝�3����T�촄�.�-�҆��C�s�DьZ�u��  Vurִ$���u·$���kX���n�rf���(>�����4`�j�����u����;�@-�VU�>��w���5��hpw����x��ʲ!��-<�1#����Q�E���_܆'�tXּ<\�1ƭw!�{]��6~�nK�r��Pd��I&�`�M_�l9������p�S�ra�+D^*�p�H�Ƹ���&��@N�U  YD)N�4Ԉx�S����
��x�t��y����Weyخ8|7��!����A\W�el���bU{��ot� ��@m�����3���m�lt�RJ��/bFT�p���3Ƙ�\ �ڹn�Vv�n�.0��"Qm=vX   %9�Z��˳�_�.�^R\ʲD,��p��ܪ��0�5q�����ɍ?� J�R�@v�\G���c�j�"S���hn�J��Ph|�y��	3���E�Rm��@����"?���U�q7S%����/�uv�4J˷�μ��F ��[Z@r*`o���o��&#����9��8ew��=x�K�M$��gE����F�9�w-�1�r�+���*���sj\����� �[V���L��6���w.���ۮ��ѵESH�C�I;��Xx�RЪ��KT/=�ހ0���n�k97yIw6w���  9��P  �۲�*e���6�� eUP .�P� � w   o�}���� Wu;��(b�ۻݎ���A�*��-GM�pp��ĄN�UV�.�(YB�R����k�բ�QRO�?����O�=ߢ�3����\�S���*�܅�8*]gSA��6m�M���
��1����C}}
�`����=e��8+�A���ɰ����V�X�K��Ov����q�8+FCk!���l�s�]k?�V7�:������s��x�x����Oy�zG����L�ř���Nj1��?�w�ZZ�r�N��r�8�p����+�f�#�B?l�n^�kH�*d�?qgi�i&Cm$�9F���.-���p��i�o;�'s��ݹwe� R����؋pZU�܆Ҿ#�N/��4V�!cצ��f���"�0Z�3��cAg�}̂ l�)&(o�����"}΋\F6Ӈ�6Vi�lޑ��&X���ȩ.���(��@�澿ë=��ܜc���:��Ҽ��UL�����U�ӫbFG�|�Ƞ� ��>��R�$�t���+U���u�����|�ӭy����Z�Z���R����Q�Ʈ�1�WqptV����E��jbw��h����;@Y-��Ļ3�7+m� U��Br�շwEwRݘ*��.y�E�G1�A+NN����\�S���l��!�Ph|;���ƃ�����W|�|-R�-��-p9�ry�=����c�ɤ��G�\�Z�lQ^2^�X[�D����%@��8*)���ђ�*����\
���\y�ߌ�5�`���j����u��j�G�u+��pp���Nw�ب/�׿t�Ϟ��A��p���-,+�야��ɺ��1/Ob�C��%T�q�UӐɎ�(Tpinp��A�p���m<P�
�J]�v�VյQ�� *����g�s����3u�U�jC���n M@��ڢ�-�I'S͟P�����Й�`0�\�S����9�Cc�Ӽ�M��m��IM���:V)}<��:~=�IzU�?J=�p}�Yt�q.�`��@���M�QWZ:lR��12��8>��mO��	5.N5!���2K, ��Nc�y��`�?�><�3���h�U(��q][:����$��p�E�@��r8��fj�&��Y7Y�:@�(���� K(�ӎ��X-�/�m�dVD:_���:��Ҽ�R�e؇�o�A���u.�\@��ň�	t�%�Y4L��<t��ƚ+U���z,}c�B�pV�����Y]�=���%�����X������9N���h�}BLF�V5T�޺�s װ�zEHR�[�������G�}�����+�4�S.�><l�8,��l�f�b%�6�6Zh��2���j�I���;�ƖV�#�z@�9�vq���3�t ���������މ����W%�U�*���c͂��y\sv�E�v�tn��P�D��'U��t6�1T�Y����j��p��!�Nb�Ɔ).:u��T�b�8+��q����j6�8mg���jv筫ۛ��  )ݱ��PUU6��D$
�ݚڪ�MmAT
��EPj�*�lxUm����*����YCgvۭT	#UJ��f8�����#c��	2 [v�J�[yUwr�lB�� hK�ِ�@�
~��*��?(X��4Wtw�5�a��/Ĳ����zG���J ��It*�` YA9N/1�A��#�*�����j�4�|fy��7�T��xd�P�S!-�����Ny�y�=W~�%�q7="">la��Yǹ��x�4I6��8�-���ƅK��P� -ү�kH�=�XY�y���,-��H�9���X�v]h`�a��S���v;�6+F�{�������D&YH�( `z.^���keC���ܓS]�[�w  ��JFvKm�ZP@ �{*�9ŏ�-�W/J��੓Wp5gM">la��[_S�̶�됒��#v�J��/���1|n����*�>�Yk3E�p�k�|�V[*����ei�%;�<t�C�������)�|Q�^݊�M�ѣ��sAh�	6H%�X�GJ�Tʱ��	9\�7KH�8����G��
zD:F�~	
5M��l$��N�zޠ�x`�%O_�hH�'���V��I��RAB����H�iy"��3��?.=�e���n�� UK�
�L]Ի,!J��B����3�e���P=���:F��L��5 saA�b���"�-��Tw�6>�Z;����:��p�U���g��p}�L*��)�Ъ"�e_���i����3�\ov�Cjx��R'=|�$S*�IPmX��?l����N�����zۼ#����X�9*!IqU�D��$�!'W��*�u�*�u���Ak�iWK����r�%�2��'�(L�6˳[�ưs��G'ewm�
kX9T.d;mV@m�� ��[��;��T�%������COH�}liU�Xs�g�3��da��.���SN j«d'K��N�f,�Ŭx�D�N�GEh���,yh3�xty�O�沔��[hWTP8��lr}N0�d�y��C����4Z7}���_^?�.��K�@ ��*֑f
�M���f��U�t��ƚ+T�,H����h�L4�R���I��a;�92ȕ�+B�kxŻ"K��������#X��جR������"*�htMU]�g� ��ҕz�nF�A, �3�������6��6ơ��
���{��ix_)�x���A�2�BP\�8-}x�nU��gEX��U��%(�W1�+����5�:�� BRRЍ8sϏ��\pX�����Ďr���>�Σ�k��ck\��KF�Y,`o��l��=W�Y�ghpS%uD��K�_w�í���� �����\��/��W5�q+��)��ny�1��=�Ͻ�[h   ��m��T�#�ok ���m���U  TJ����۱p�V��l�U�gU ��@=l�C-J�m���o7�����A+.v�\�' gW-� xogw�kI�z��P�Uw  ͪ`"�@��UVJ�6����$�+�U�nѫt��a� )��:�Q2�mR���u���P  �V�m����w@� ���9ür��/ש��U<����¨��-tCe꠪xc; �n�-֍ܽ�d.�y;`��U�
y�ۯ&��z�^��pw1�s5X��]t��ԯ+/9�*�l&��;�g�{ � �6��8J�-^]���Ҭ� UWR�)�Gc���2���9��r3�ƶ�yYB7v�Q�HG�膪��y�� 5F]t�;J��3ճT�����[��e��U@�B`c����kk�{4]�b�xl�m�Mi�c�m�e3e�]td7\{TV�T�m���8f>;R�n������X��gP��[kD�y����Aխ�*��
����Z���p�����   P        l���ASd �.��j *l 6�z� [    *����@Uk�  5۪�U +%U@��n�@���hn��     U  U    >x|Vu@    �   �    F�T 
�� lu �@   �*��  �@P���P    �    �0P��<U@  ���         � p �@  
�Q�ڶ»���  �r� �[@���ۻ"={P^�@     �U@�*TW^�@ ��� U   ����WԨT�� *��Wr�i���=z��ui�z�[ e�+ƪ㶥�ސz����U�P.�����(�՝���\��]Tz���a�0ҕ(Yn6f�f� [�7[h�wl���!cyZ6vˍ�K�L5UUTU����@ w-�Ee������u�R� +;�  � �tU@m�Tʪ�Y���6u�� m�` )Q���yUZ���{GFq�\[t���a�;w���U*��RPuL`�V�i+)C���?/|=[�x-ױQ�h�ۚ�%+]�	�U�c��w!�+f���5T��u��TW����哮�m� �#,��������ƌ��w\0A�EWעƊ��E7�������������I�!�>2���GM��r������4f�5_�@��#�!D-��N�����|Y�5��Yz~�en��z*Ƌ��ܮR���J	 �1�ժrl��](t�^N�v�uzݱĮ4�U91cZ��;��]�U|0|­�����{����]��w\0h�r���Z)���T�\�I�h�H"ګ���θ)
����Ex��֦�(�����H:*-��4H	�����'+�����+H-����*�x�E�"�STl:e�hYDWN-iF�uU��^��o?F��u�7�l�T�b�V��"�	��l�����K�W7T�9���E���cU���0XҭN�����-���.��f�c'j�kè}��N�v�*\�)v� ���U����T����%��F�sA�W�Y�d�VH�i�63J�`�R߅���0l:_&J ����`�C"�q<&+��H&gC:�{5����n���0� "g%8p�#M��+�G���^�$����k�7��Z���,�mm�
8Zi�4
v�,�W�G���Y�zG��t�D#N���<G�f��J�.�4�LU�4�:@}cdy��xMV>Dp���wu�Ȍ#:�U)��*a�ڷlv�\T�U�c�Lpb5��ڸƩr�UUJ�D)b���ϝe̅����l=T�20�6B�V���[ן1�<���cU���Ro�E]�  �n�̎�{�Ŝ?������|y��W7���K��#���hXUٻ��t�ײ2m�@%v�+�Q�L jx&  Ԕ�~������ɫ�9�q����<����wǵ�-"��IKh��9��%e���X=����U�A�����)�j�`(�c��p�q�@��х'�.ͭ�+\ \�۰ݻ͈m�M �r���7���#g+xl�6r�A�4�E�xx����:�%�V����
��_��ś��ƙEH��corI�Y�s�u5�ܑ�UX��l��)r�q�h�ϳwL�{C�P�$�/D�Ti"�6Z�Z��h��ԽJw>��5��\yg�l��c�]�D9d-,cqW����mnʝ-{�κ��mʝ]�j:�>I&VZRge��UW,�
�= U3�v��V��M*��@��.`颫�ݑ�n�.>&Ӹ��ˢ�/Z�k�yLj�*�զ�%el���62�f��$d����k7[b3�)�X^Y�*&9Z� 
�k/�*UGp�T�X�;��l 6ʪ��+)�  
��  ` ;��~��
���AT���������Pn����<���tv\Gi6U(9�g�Vu�� em�*7ymV�ub��H��@��g3:��9���]���|w�G.{:�{"qW��$0URTꉠ[���&s�md�~�M33��K�rL������� �KeB��%1%��%I1A�p�*���M<"�!���B��i�.ʻv*b�C��`����]!R08'��!� ���rg��?
�i@E�X��ֱ���>a�q�>?c'�
�`�jN6@�`��k�Ak���@��r��t �W9�wg����tQ�U�qJ�* T���X̕�~#���:2�#N���u˙^�()�,jVRV
t�S�*x�L߯5�5�發Q?��h0 V9B󈶸ᜌ���&,0��z;��8�Q2�D�ƬA<�q�>=��U
۶�#,���־k��t�Ǎf�b���I�pUك�s���=5�],m�@` K"��Ʊ���l�,T���y]AV ���Hx�+�F:��i������F$H��W�Gv5pU���$��ȇ�����>#��]���ȑ}g����Yء`n��c���9i'����t�U�6�� N c�-���;�rWd#r��?��4[�q�
�C9�f���T5C<�5�L}svl�����$�[
�K�֖a�'4#���8펲����V2����Q����n�| �e��*	U����������<����HA��r^��Abd8�������Ңn�F�9K�cX���'�qx�э4~dv|���,��_>5��6c��
�!mn�)y�
QNVpc|���������m��_��>�5�9w'.W`s<LmR�w1���Zƀ�@�͊V����D�Zl�؇�ɜ�/OqV͵��=���fv��خd�0\$����L��Q�|x��QTjP�f�i��3����a{u�&���� 6�U%�����[Gd��<p�}u/����6eYpX�5X;P�	I��)��	����AcP�:�cEX�K�OB+���)B<w*v5pR<��+� ���8�>�53'S�b�U��3ʮ*���u1�h�׍q��o�l�B��m��-׃��]����gE�u6���a]Ԭ�*V�U��⚠YZV\�__�Y�x���,�6xWv+��e�}�l�A��g�����6<�H�MRMQ,5p�|dp�c��<p�Ɏ66�WKee����wb��V+��Y�=�������5׏���[�udCf�/S�<�⠊m���b��X�?��yo��IJH ;o4dC�W���Y�W�y������?����ֱ�����cҔl���MIE�*
�ٕe�Z0lr���bD��ֆ4U�.��p!f�w~v��������jڕeX8)����c]+��m�J���P ymo<�qvM5M��ͼ����7�
���玹�2�U9%A�dplR����uQ��'a�v���3khL�Y����d��K�ȝ[r=�\@ �T��[aUT���u;��� m�U@ � �VR�w 
�`6� �T��^�����z���]�� 2�k�b�&yr��|�����Cj�w�s�wU�\�D�=b`Fʪ@�����qq�����Y���-�,��D>0��9z;�Xj
��q�U|����$pP�C�%+��������f���]j{����x}O#�kA���૳������v�e������_�g3�m�Vj
�˂�l>
K��AX ��	Xz
G���	�Sd6�.�i��G��Y�2k���:_E�n��f�ӑ[�b�b<0Q�}��XkE`���́B�$�IAsX�l���K|~����tLƇ�Z����,�g�u�}u#;�� G ��Z�y��4���d�C�P㰒+�um�H �+3%Frl�)r7R���~�5]�1�s��!��R�+?`��!hb����n�`�+�$A+�4�M��E�����X*�N�f�݋$����o�r�ޛO˙[R�iA K ��d�f����.)�u�uΜ�v-���]�^�DHIx��n�ti̗��es|���P�2��C3�{!0�t���+��KKH&ė=�	V6Y�.�ʆn:�3'S�Yro�s�S�������-U�D㑡�V��zi��]�Q����w�@���  �G��1�.o�N���>"ȝ�=��+Z~�(�]*��������"9�Ar!�t�CM6ʤ�m	_
�Wg]�zP������A4��P��dx�݈M�@x�������m-�D��E놐8�8G"tqc5���{|�гC�4��s~����f��,r�� c�w�:Ayv�*���d2$���+@3����#z��V:F��*�!��@-���e�,Jj|�Z�\��s�U��u&^��t+6�N��!X*9��A��;<����YG������5:W�vғQD�9iVtK��`y(��Ds]�K���`����ގ�;ΐF���VkP.��i�����m��R�}?/���i��-t�kmU!���r���q=��1��:�i��7w��[SB���4ٓ��� ֖|E������Un�*��@��$	�D�BI�YM
w�GO��-	p��,��d{Zx/+��!����^�C8��$[��@�_:Fb��e^���K�W�y�4gKt򀣦�[����n�^l�]S�ً<v�<��N��g�wYZ�^���J�R @+�Dʻ0$̆�5�XM��D���{N���7�h�˧]f�h�tXY�k�?��X�x��[%��@��WgBS�0����\4~5rxl��XW>+_�K=�n�([����&N/�:�J�����3��*��Dx�=�����֖���}��}���#���$��е�Mޟ5��`S*�dg/�jyU����}�^�����1�Wf��J
��M$�,7sO���݆૳�a�*u�G���ք�j�³TOM�����uX��In��VK<� ��hgQ]�^��[��0U<�k=�'�޼^�5��/G:���5�����+sսs܅`V�X��04X�jq�n֦6<���θ�_�|~|>. �b���gMK����h V�b�@�R�:յ����l�@*�* �l�  �� ��0 � �PVM�@�m��R��Tc 	��5­W*�V��Tqf��u��;*^99�F4���Nw 
��̶mF���hX"/�w��?��c5x֠;ύ#<�o�ʼ��i����p�w��sl�%: �r��<Y���M5��E���^7���w���ӮX�Vk�Z0+?U"�l�I&[$:�1���<1��b(&+��ެ�*t;�Ѫ�/}��2���m'Ty�\���k��Y��X[�q��u�w���?/�U�l}HL+( 2��zE7�:R��<Y�Jxg�d�,�_*@��]S0l�Ga�dɍ]�@��Bx1�ή��m�P.�P4��U����[v�.��-��݈lȀ\֖p�xU��_c�ޫ�Lh�7,N�� ��>��Ȁ�I$�M�I�g�^���VkF�aҝ�\l���l�[ύ��!m�b��U:SW"�aZ_F�pߔ�*�UU�>O'���S���W��+�<� v���;�����}y�E�?z$��,�GD�y���C��Q�v���Qn������qS�G�����y?+��^��X�q��U��Q��Ca��~}P=-=l�nx��b�g��<񖷭�tV�P��R�ۛ�[Q�A��d��\�_�:�sW7bZ�(;1�������Z��>����X��|��D$[$�A ����P�*����A	m*��X���Ȗ>39���:Z��A��N~����������u����ܨ\Ao�FY��\>=���ܻ%���4PUb=6������H.D:'^cw�����ʘ�c��y�Q
���B
 2X^.r$=��W5�֦3%�����q�#y t����%DV�q�++Xxu\vˆgn"��"h�X8�m���)UV���Z��ik�����ؖ����s�hl���Y���j[&�fA����͢�E�ȇU (Ӆax�_�x�\F���mZzI�y�[�N��R����JIl��Nj܅Ӧ�����f�����ۻ�ɍX�������n�F��ώ�0����2��-,)k�&����v��&I"���Y�wq�ݼ��I&[%/������׫N�-�q=�� 청+�F�΅Z�V��n�lq������u^���.��%�t.�'������ɻ�R�b �@+�nn�O��w�s�KdI��n⭳#��t�L�)�i$�e�^���E���;�:w�t�������+�zh�g{`�!QdL )%�1��͜���o�[����+�R�����Ci��5��Zx�p���E A ��I �)�/��4x��BC�hdpX����a���ϯ1���d�}ݻm��(��Be%H
`[f�U�<k�1�컕a��n������v���6x�5�ګ�Ƕ�ݞNa�UԳ�$�y,���-�k=bV�4�(�E��`�`�)^����F�f]���^�nm�x� S�m�Px m���&ݛ�;��l 6ʪ�l
��*�w   m�]�J�m��j���r�P��w�P��^̓/'aCr�nֻm\[�cT*��䛰-�@��U��h�*-@�ݹ)RUT�߿:|C����C�òZN"Wt�L�?x�� �c�2!�:��u�0��S�sx�X��{"֡���\"�;�Ʊ��\l��]?=x�q�679Uqm��e�|����'�\?Y㖪tb>#�Z��cEX>�z�X�E�o>A��l��d�Sn��y,/�y�+<p��Խ��>�q��(X�.;���X�a�Ȝ����b��2qc�f>��[��ta,Ih'?qöd�E����N5���f��J�h��	X�a�=7N4�����ٳ6��W{�*�b�T���)H�6�lf��\��,0�������x�&+��a��|�f
�����X~z	$�e �!��D��c�04$�|)���}]e�<|C�j\��~�}�����S��^��d����5���Ǖj����x��pфx�L��0��ۑ�kU�����{d�`�� D������T�)ȷ?a��J�p�!�]�d��B,Çk��ꨡ�SY��F n����5�Z�|��d���R)�p�dY��y6Dݵ.E�^��������eC��V�p�s���Ԗӷ���*Q��puJ�뛺� ��������>}=���֖�8���Z>�[� �	j��P}�s���ȨYk([l(^kW�vy����S1Fi��8 �D�*�b�_�7&�x�����6�m����(qy�Zp�8�,��}���Y�b�C2/�Z`Q�dh����A:�l�H�I�yJ��^��+H�,�{t�C/^Ӕ`��I4Aj���u�g�v�y����pAT�&,�ϧ=�o¶;c,
; T�rG�-��]m��q�RNj-�@U��P n[wV�@dn�-����
NkK_���ևgF��P�)��W%�pU!+��o�1�pN�D�I($�HE3`}GM�']K�x�yX��i�U�ek�@�yV�1|��ϯ��yv��CN�nA�;��#�ȕ�za�{w�)̣"¸�ª��b�]r��|*�"3) �I4�H$US7ő��\�2�>+�1���OӁ����/�䗤x�2O����Z6+mEb-'5����w��o��$�R�����n�1��$&�V�	���vf;pZ���86�%��������*�6M�v��wcF �d�+�Wŏ��}����\��-Qz*�y�"�$>5)��!��o�M�+qih�@BNnϚ�2�*U��-:l_O+��3�Pѣ�1@Ɗb*� �6�D�KI�U|l���*��x�z�0(�+#�ڗ�3�=��`
/�
�6۠�m��qAgf"�b�=4t���I���m�N
CF�h�4A�� ��I]�`[����W�(�
�uAp1^�W=����x���\��#������>@���Q���x�?�Ȝ����<sp /�U����'�D)@�XUWԀ����@��"
<�
#��PA_Ǎ��\{���9 @R�@ �������~������_�y��������}�������D�������Q��R�D�����������'�s��'���@��u��ӓ�����������������@��0*����$*�
�����P>�π����@P?�7�ѿ�����_����xz?i��dw���DW�q���/�����}�}_#�������8���
��Gë�����_�(��|�D��NO�@ED|r}�"�
�7��k^k������냏�p� (��������
��?O����s�����{�y��w�D@P.��A݇��Q~�����~߃�U�}������߸�}~�=������=u�}���J"������>��������^�=��ǥT@���=~��=xED��՟������d�Me�͸�	~�A@���@ ܟ}���o� }  ��f�M���6��n� c	v`kMkg�vȴ�����^p 6�nv�,���Tu�8��N�U�v�N�x�'fV�-�*��a�Ԥ���Q�"l[-�0�� �   ��ݝ2�ݚu(V$�Xf�J���+��0�+W�     ��Bu�A�݂�@��z =(:��qJ�d�}w7�  � � � 
�B�, �B�lP���\)$TUID���OYIW��E+y��A������<�:��x7��>�klz�N�w��[gAUʷ��A@����z;�����ϻ��l2��'��Nm��={�x��������xz>7��I��x=�B��}�����W9��F�u�w���w!l�y�����۫{��ޏxMU4$=�ƺz��-���k��
�W�m�=-�Y@ql�@а�n���o�k���#��{<�=��U[��V�j�P�oL�����7�q��C]fz�^����Z�v����zU��k��=7g@�]�oj��	�����v޽��;۸s�j�pj��o{�.���$�٢QJ�PT�>��mt���E�;�y\�������m禴���:�����zj{�R�f���i�t盞������,��{km����oj�v���k�����T����@��ɣKjP4@m��=:�����׸ެ�a�N�F�ܭ����
�W�w�/b�N�n�ν�W�w���]�U9���4����8y�zU:ɛ��px��Z�J�5���*V�DR�>�-�42��^�	Q[����y��(�-^p�oq�ww�9֚n�E޳������;b�7KW����͠w�=��Ɔ�c޻iJP-Ǵ�����%v��՚6��>Ru��sN�e��۽��*�ǽ�����43n��� z�)��ś�g��O{'�v.<����酳޹��{+�^�y곻=�N��z�N�b�YRR�f�-j�K����{�U;�=��מ�v�,����\��{��[Cַq�mZ����g�o2��Ol�u�-�ۣ���j��w��ч[����zg�V����bMh�ٶ@cv�h�q��{��^�^ޫ�[��pi]�o{�=����^k�G�ooG�ul]����wj�V�����vU��{��kF^��{ݠ�ty��i)E�5�=��t��Z���u[j�Ǔ�ij�GSO\��ݮ����xEu{�G]��7YV޲�����5�;Y�QO��ݮ�׽[�t�k֏�1J���>ܡv�SZ��Hv`���I �U�]��!1R� @ ��FJU@ �  �?CF�U%OS�h���5J�A��&C@�?A)U40d4�&���$���Q�z�OTa�~�����������1#���bO��C,�W��9�;���Ƴ��@�		'���������!$H��!!$�b@����?��HI?���		&!!		'X@������?���dX��$Y��"���#_��o�7�����@�(Ad��?��ƻ�ĩ2 �JDd�B�dm
+\�#���5���%J��[nJ�,�4�@ձ̦�T#�&�dQN�11U�E9�Jԉ��j6
�����%d�ՐX
A���#$�Y6��NB�IY �i9�4����VJ����+H,+J#+X�(�P�*k�bA~ ��+��d�������2�@��~�4��,C�04�4��!�cl)�ңm^R�7e������ �Ԡ��%�=lb�%X�B��Z���EA04�bB�2{\ޮS���`m���!�2��q��J�(�C�B�*AdƲU-��A`6�g)��H)��))��Z�KlA�1eSB,���AIR�A`,��m �QYZ"�j�j�*b�j�V���mY14�C!�
�T�`VM3����m�X11���)�S+-&!���
B�Y4�,He�2��f2
�!�
��1�VAIY�LIP�+d��*J��
����,�+
�IP��Ă���`6�m ���2�P���߽�s�9�I���kۦo1fPݗ �3(3#C�ZDne�_�V�Jv��a�?}p�A�v�j�D�먋I`�9���z$�S��E{����+t$�&2ʀ�H�z�L�?|	�
,X�b�&>}��޴���
2
H�F(�DUF �3;w�Ή�R��l-��`LZeZdeVi!�C�"�mVN4T7i�/�`q��2k���w�n���uv^k-)��6�� �:�G�Q����׃�,�C��數�֌�7d|!FԴ�;�V?�K����&����Q����yV���]��\�(`����Y@3R�m'x˴�V�re��v��i�m
�4ʊy��hQ�X��������# ��EQ��TUAW^�^�f�Ovk.~9�������bK����hd|�/�0���e���%�?�"�OE����{��%��.�G�w3W�}�f9�I$�"1T���gG�3ì�����o���nl�+緇f6�?��z��U3�-f��X#�벷DԚt��Z1%��Ǖa�#�Z*�T"��<ww�y�W�'A�4�@� �j+f�9TX�R�I�{FQb���ݒn'Ү[ʠ @�gF+�.d!�ti7Eɘ
�1�DTƥ*ٶ'�v��[�sF��""$QDE�	�Qf/'ŝ�l*n�i۵��5Q�9X�ګpZ	�I��? %G�cUQa��UD�EԚ���"��^ׯ}}��\�i!P�E�Ϲ��{����d-mBp��,��/}�vPAPX��{����7��L��ͼ�]��z�k3VJ̝"Ds�լVu�A#q�����R ƪ-���3	�b*��X�b�X�� ��PP`�"������#W����n��T�(����T&e�.���{�F˨�^�;okj��9l�61K���2�����
I@��mL��wj4�вj�=��8�[(k��ֱަ�{[��uw�k���$R`dR
,E(2
�R(���H+A��� �V<h���H,UUF
� �"��F,(�(�UAETQ@X*��""J$DR,��UX���*�TV"��V(*�+DcA�bm�pO���Y%v�in�V�ږ�e^%1�d聺!��Q�f������w`�#W-	�nĖL�;f�x���XH�Q�_���4V�:�7U��(lК�N���V���Q-V��0G��U�ڻ�����T�rFeˎj�kYz+6m�v)~��h��O�+8he��c,��ɉ�^��%ݑ�)tp��R%�vƬYvE����u��z&MZ���X�XnT\�O0١)�����XAJ��r���mѱF���Aʭ��m��>/*�"��9a;�v���iU�P�#��*�W���z���$@�r@�.ݍ�b7Z�tsr�.�2)�to^����Zq~G,,��Hj̆	�S�t�p:{gT5`�@�1R�i=5��թ�N�:�U��7xl�4~!˂<��'IV����)��)�7 �7?2]�*͉Z��A{nwcoI�LQ�D��j�:X�̂	X�n�p�nMԒ�cV��VC�b�w
������U�p�ea�r��ea�Y8wT�2�AS'z/TC@���X�!��Rn&Bj��ٶ8Z����B�[�v�ʳ���/̓�x�w B��e�{�,6�ҰQn�1�]IZ��/U�#uh[�X���.a�"�fMU���;�J��x�"m^��w{j�i��<�Bࣖ���}>�)m���4��e��2+���;�����'��=.��K�hHq �q�%EEQL�R,�b�Y,�b��Z�b�u�XX�iP;lErш�*���
$���l՝�V��b��Z��yM�K%��QD��L��#v��S4��2�Ae��%�);��7W�1 ӻ�a	�JtJ��Q���u���Μ���L��C5,�4�7����R�
�znQ�cK'^��ml[��a�˵�m
�{& (��0ҭS�V1�n	��5���r	��rw(�ٻ�9H����Q�[4Y�Sr6�GH��Ez�X�dʻ�v��t��Tsn<e̼��^!�rXiG%�Sʤ���P�d�8Tݡ�t����._GO�*���E`t�+r�����`��0�R��Xˢ.i��ܛM�r#+(:���ׂTɻXf��Vb�,iq�/Z�n�0�r��Ut�8�oI�g	�ʅ��ط�S*&�cx�����\D]�b`�&Rę�b�ǆ^��Vo0��.u\JC�X���W����F�pJ�Q6���m<h��Y�<��'���i���rg�:�ڴ���w�� ˚ɯ��PH��ZȄڻ���E�Ğ;,=l���-Rr�g����:�S�8,
��ѐ�O$1�3ɤ��a�#օX�X�r�Tp�'��H��@�wG%�*��v��m�$� ��D��ԱU�Aam"���
aQv��!���s�ֽs�ֹne�T�2I	�o4�H�XzM���o��ʼV^�����n9uB=swc��E��p��fʽ.l�ZB��+�zᗲ+Љ��hJ�1'{D\b�50c6���+i�nZ�U:�~z1V�I̙V�܆
I,PKrl�E��. �Wy�|yN�j�0�҆�kU2����ׁHWL!�
��QV5Q�*��t1�Tc�QU�YH�6�)R�Z������qX��
eI�RHi#!QWl������Hy!���
��M��2�!�Xv2bCi��d<��d8��!�$4�W,4�mJ�.����N'7`pHi�XxSvX��U�6-�Fy
"��O$
3�(���N���!�x�H�9K.�P�TRh��$<�'XT<±�`�-���Aa*M�VHy20FA*e�Dl����S�p���N����-@4��@����Bke׳4L74�a�N�&kw6�+�V�0����+X�*e�uj*�
����O���Ӏ��%�m9��f��P���yF�$t����G{�AͺuI�2+��B�E�kA�^]�Q9M���dFC�UZ�e[�[��ݙw��������bq��
�)�~`a�R{Ul&(��MU-Ճ4iUn�J�J<ז�@3u6�	CU؛c2�w[A�;z��V�5.M�)�i�������ِǋc�>/6���yר�q=����yu��ĪEDX�b�lELj(�5A}�{5�:C�ʫ5%h��kW��Z��Ћ"�ƽ�K/w^�l�Q����YI�lF�٩�c��]��);�T64�7$�z��u��^ܐ�jhC�6�f��͘�����
�?��APX�qZ�F��Iu�^;w��.&����B�^
����	�uU�Ygb�}�;a&�4�D��5�5�\�������MF�]�ޒirħ����Vn6�=T֋�Ve����l�ҍ�>�� �S&��(�]�F]T+������
k�!����n�j�ӻEѭ-`Jl�$-�9�H&���nd�wi��]��aՁjK�z���EP�(.�����5U�B�,$��h��Qk�)�;�G2^Q�.d[��������.���#`㴨��˄ʩ��[��ٯ�&��AQ���)�iE&�h=N�X��aq���,̫�4�6�J�kT)���4��b�#��7P��.��Z��)`�����j3a�Y����Ap\6��[j4�5;-����,����1�Ӥ\"�e��I�M�O�W�B�^�V�Ô��;ᢡ2H��e���K
�����b�r�I�d�m�j-���و���-�����~$�
�������,��H��x�TEU`Ȣ*�PUED#��w�ֶ�{d���le�'I�E�b�,��/�C_�<��Ӗ�y���
�A���S%�m�Y����iT&1mjz��*�J�?���s�\�nE1�DɅm[ۢI����t^�U\Q�61��N���Éᚌ�o2n�R���ٚ4ِX�9wNݺ*=w�ԕ�]źoi�G/,1���+��l(=%�]k���{�SC&�N!QH�\�	�d�[W-ba�xC�f&��ո���V6⁙���9��̿��"on2�i7�(N[B��`����fY�j�9t�AA�Q��So]L��uT;J�Jx�Zg6S�J��2��c�֢9
�7e?�A't,�Ѕ�wS�m͕j��v�Ƶ�ˬ{�FL	Cח7��͆NC�2�\)YWTh��0�m����Q2�n�"�ҳCokU�d$�8��l�-~V��Hu�P4�m"'�S-e(�H,�/~���K/-ػ���L�p(q�2S�Pm;
�ɚ���+ ����Z���ӓ(M��컂ʂ�Xp㣏�7e�I�5ZD)�\�f<�m�Ш�f�٤ɨ�Jbo%h��O�^~�
ݪw�7�I��"��-d��n���f#����� "y�6�`wVCLҳ��@�d8���v¾I�������6����X���sNffwzu����@2`q!�C�d�q�J�,��� ,���H0��a��1�^6��v�`£ɪ�
�N&��c$�șv�5�P=EՖe;�V��
b~@N`g����$K-n��4�Y1��"�̼⎻�D������>�b!�|o{wi���RӼ9��MEL�Ӂ�&溷�[ȃ��F���EY9o���
M�W'��M3�@�3��d��u�R�]���Z�pi�j],j����a)�|9�Wʼ�烾'L�/�F��[����#�6+굽�y���!n�7�$�u��\�#X�MmX���7���D�u'y�����ΰk}���6��D(��b�u�"^������CJ9^��y�lr{k���n�s�K��Kv1�]��n�d�čl���4ԧPfk�2#ڕ! ��[��}u�a�b�ݦ�J]3�JHd]j~4��vM �� �T�M=��CoJ}��3/�@���}k��.Ƭ"����t��i#�9�����Tj>d΂�LӖ�)v�<}�Й��,;��\�x�."l�ۀŽ���p���5�	�֭g7�WS� ��[��oe�w���!�f����N�ؔ0��Ve�������ǝ$z�,�yH��P]7Q���v�]����t�B��5v����sn�S��6�30��Ո�ep��,#N]�͝�-�yID�"rg6)�x�^�w��ϩ�쳹�s��&�$���)�W�R��X{I��d�Ҏ��ŌdNU�K����s��r����E�Éw:��'\���ѱ��mE��j�/��;���q>�$o8Y��ʍ�<t;�U(�<�c�P�V����Oc:z,w��u�:��*jfoZ��wAc���p�#Y!�/Uq�Id�̈́���Ԭx;������=]��.���z�Q��'h���u��}���h!b�<&v�;�v�Dr��Q�Z��ڵ�;k���D~��ׁ��w���<���[��;��ֽ6r+�=���r@h�B,k����k`T*�a�fӫ��b�pk|YN�_A3�y�HC�hr�k3gfQҁ5���qӺ"�c����N%u��v����i�;4EX<  ����ʂ�b^�Sb��J�.�ˡ��uRY���kn^~����p����1��{2Q�����Y(�7a19�w>�2v��XA�[�����%Ύ���6Wغ���J֛9�q�b%FuO8�EU�%���#�҃0w�Sb��8�ۤ���A9�7I��	6�7���e��`7�"��1D�U���xQ-N�ض�y����	f�`�ͣA��4Ů35T�4����vss�2U���5)K�����ժlN7���lb�C�0خv���*�;yZ�V�|��|.F��>V͝��l�뉞Yr��|�wO�����g5��0l�H�'%۟GnI���td2�XS����ř?s�=�Х}����sf�|8��퇹�$ۙk6�g;�P�:��ioFIk�^ˌEuv��}�������.w]�FQ�m�w��]��5��.�RT��l,��R�۶"4k�4�s%��Ålt��ƻnezZ��K
�PWTc��������G*��yh��q��齊��z|X�g[��S��Y�6$������^Zx)��yb	�ov+��"C��#Rn<<��ɕ�:r7}E3��!{�ײV�iv�aF�R��FA�}�[}@��:َG�@�"��Lv��?�X��rN�����m�"9N���=��DXS������vG9l��镛I���\Gy�`1U��5+�:L�%�ĕ-����u��R�:XQ6Xݜ^t2��P��b�N��b�H��f���0�|3,�iV���t�+�o%7	rf�S.m���~O�]��ֶe_[1sݩ[�)��!�U��<UY���^V�(�%pɸ�p	�ĺ������L��]�eJ55P7�F����n*J��2_gP��7�:�Bxz���&�<�K��QП�ꇔ�c	�iX�뵉z���]�)��\Y�K�\$m���ӧݙ���!��wz�o"�Q��ۜ�hm�Y�	�ަ%��@�ߟY�˩�j�n���6�&5GG����*��iu����OR�1���DŘ����6 �LQٙ�ʅӺ{����3)��W�6���P��>{�@"ȣ����jՕ�ѧO��|7+hv��3-�����ԫ���ݗI�Q�;(s�䬨.����JÁ���Æ��	��׶�װm>W��n;p�g����.����V�����G������+��;�u�_�6��P�V���Y��Z9㣥l�|l� (�ot�0�*�'�E�������0�0�[=�ா¾��N�:�>r�yo`�	�w��|�mv'��r=[8�K�e�gK��gM-thU���)\oN��Ke�W��1������ܔ!���w��vY�A[���m
���-�1"���^0O��X{�k;����^z�ç��]!��s(v\Hr�6%A�J� �ʶ�c{=ٗ�����SJѬYx�����R=݅n5&���gǕ�wp�#�U�wzK�����@�H�� ]K}���XwJ�� ��2���.��2r+H���@;����_��Mf�+y4I)��a��.]T̕|s<:�UT�a��j`Ή,�J+7S���^�*&vk�ZY���	�wyi�ku�`���Ue��Q�Pi<����5eH���ɔYL̫�����Y���E�Pf�x�v��� ��;Nٹ+���jiWvүe��d�4����.���f��R.��E{p^o:.����+f�f������d�o2���RO�x�{�	ٱ�-:f0v�5a9Gx힨WrY�eڋ�X�fԺ]�ڮMq���
�9�&:u��
��m��Q�������Y����v[]�
�
wM�1�غ��읋��{~�u��\#�wk���r�g�ᓹJG���ޭ���ԏP�{ۜ�;��WCId[�v��h�b������\��բ�96q∢YA��q*f�Qф�ؽŊ�����֚�;g�V��#�w��*a�;ɻ�P�����W:��Zh��B�P�w�(L|�{���t<��	��ә�6�y�ʏ#ܳ`�(���rP9����[�`�}gn�ް��8](�zk�СN9�R{�0k[�Z�7H�k,�YtNA1�Wa����e���LToN*�#H�ֵ9b�C��̠t��]`��
��H��T�l]N��k��c���JRN(u.Q���>�͢,ɋDQ���0���%L��X��K��x�gX�E���բ���.[^+o�L��0WR#���94"\��|\�n�3��s��.���0ld�Y}c���RKsk�Y��@�D9
5eN�1ٮԆ���7\;.<D�I��VS[o4�[L�U��r�����
r�4�f��ޛw��}�yڟfwf�]Z���I��� �
ڹ��d����u��ˎ�D���z������o��X��m��w-�B����PM@!9@�#����ь�N���k�T����xVt�֠@��Th��Cz�ֽz�[k�jN���[[�R25�P�e��������PE�ܻ�P�U��6;[+ �0�uPf�\�o.�3�зYr�P��:^J��nVv���m�0;]s���l
R���)ھ�o����ـ��[y���=�io7r<�ۉ�׎����lc&�    lm���ԍ �     ���iL���� $m�hl  ��!�H�ȚM m���  m�      m�ۙ   l     6ƥ��  �6       �i6�ܶ� lm�   $      6�$��s-#Q$��dm��4!��           $�                   M�6ā!� �H    � r         " Ā    m�      	�"m�nm�
��lm�  ��           m�  R cm$6� 6�lH`   L�`m�              �`              ��            �    ��       ��C        l  i    l       ��m��   lm� m� > �  l m�l m�    l     ������           m� l m�      �     �8}��~�_}�d%��&��G6��,�W��}�����;��rf��z��,�� ��k��'�#��nɜt�7q����ڃ2�5xw*;�BJݕ|��I��hjN]��;m��q�W������)q��olǌL;�8������,���gӓ�Iu��xX쉼ؕr��&(�f³�p�@�L�j��۴SȮ^y�������2���,�hj$�-�&-US+���vL��fm*�Iuɢ9׼�j�]u�!���iWe ������B���o[�t�R�m�iD딋���$�IX��Y�l�p�M�fV���|OT�D����@ȫ���P�w�+Y3件ۈ.�;��`�w��O����4�T��9J��=�V��m�J���>8�-l�o�'�$���ejh�庹�ؙ�m�v���u�3����v����7U˙����&o&�H#�	��;�n����&nq���u�ܴ��V�Q͹ӂh���2���b�����9J-���nt$�emY×Y��-��}όNUQde
0|طE{�j^��������t"7��jo�p���Q�W��Vý�B&���r�ա(��|o@9��>ԕ��{��T�"����c�4�̺c�,e�`�+OiDʻ�@bT�%��*�����&���l-�*�P<VB�̇f��	�ձ=��w��w�:u냳n��)�^��V1��_i��A�P6�;�"};�����u2�xێ�JwP�+�ngΎ���:.Y��7���:r��&�[�Es�"�W��l槛h�UY�ݾ�i�eq�Oz�6n����}��ݔ��ނA��*s���Y�嫳U6�Q*�n�M�Yn
2��J����5ܷ�xPt��+3�ݤ�ņ�����A�{/[���p�{���κs9��9�6.-�Cs�L78�%1!$��	� HI�āĤ-(�P�'-��7����72 L�  �m��S)��[clR�4�!��8s.e�@�fs\�A-#L��2�S@����:�L�oh��M�#2u��w"'6o�b��s�e��h�P�����L��pW�:��c-kƯ1�(�	;���h���F�t��U�^�}ӮSy�%��AXy�6���:k6*
�r��W}�[]7���M�a+/9��-�w��yX޲�>��x�++-f��:0���#��� ����r>�ˋ;�1�İ�������4��;�4�i+��ړ^��x=�M��Q�V���:��~�%j�*���N�38�Z�%�ڣ0�Rw��L�Y0�	dۓ/QG�>8GP�:���lA�8a��ٝK�1��D�_�Tj�6��T�    �l�nd�t�        �L�   @   �` lH`�M
U� C)/ta�<INv����I�������C��/��f����P��~�J�����t��K�]uۀ�\:]3�6-��a_�b���a��4�^R$M�q��3/�{(�Sa�GyΔ/�h�٦Zu�`)�]��p�Iὣ����;0�O��t�.S��7�fX]��K����,��k��K��Q��yv�_r�9µ�[î��[r�Pc`�\�7�C4�j������X�r�c�ǹJ�)CL��t)�R�[[����sk8ǧw�e�Ƿ�@Wc��1pmp)vň1W�3������'aɽ����v%���؅M����O���^j�`]gl�
f4�`�$�B����u���t���\�5V�����E|a�6������d����j֨���뾝P��A��E�)
:�����cA8d������F*����gX��.��Z�shڀ������iu���7��#s���$|��� ��1\�+Xdj3oQl&����&���X���0�I�K����/j���������q���|�RwWw�%�uq�\��3�V��P79S\c��ߓ��磺mS+/�����ҖD}+H�0��@]5�Ԁx*T����-�Wy�}&A��o�L��,�vR�1�`�壦,�,�;َ�w��m���:&�rَ�^j�/��0�)]u��iD
�xwe�	nؽm+w�H��m����%QU��ܮ/Y�7id������P"����B�ݢ�;�u��.c4������di�L�>�'F�Yݱ�5vcݶo�<�4r����8��/�Y�me�.���of,��K_1���إwT˭��[�&��[Y�*:�_v�KO]N�U�7�is��q���&T�n�I�k�5�34���u��v�e}���k�AuVP�a��+r��WV<�!)1�Y�	/o&�t�ՌAy�ue>�ଃ���������,eTdFQP�D�^��Te�Ղ��N��m��QVӈ�Z�[D��W1�|n���X�;�p�o��oB;�3O9A�JV���m����˼a��!�yz/L�O_�x
�����^t7���*&�4xk��D֎8�vA+6;v��樬����s���]����7S��yFd᝭ɶ�:W���o�iR�L�f�5�őm&a�W��]dyL]�dT"��R̬{S%r��Z�O�[/���Ew]��R��me�{!��m����H����$$�?��6I$��$�<� ?$B���$'��$?��@��+ ��dm @�!d�$	D�I�$1!�w,���)$��	R@4���}�HT��B��y	%- 
0��J�,�>a*@7h@	��Y!�� B{V�!� ,VB�FH��1�}Bn����&R@� I{d&2q�����ݔd4��?P(ȰX,�����dd6���d��'P3��@�	Y�/(���ȡ8������Ȱ�]�T"�A u��哌����``��-0�i��?Y�{�$~l�q>`g~��i|�MX$�ff�Hf���Vo)��m�T{d�WH�"E6�\��ӌ��O:',�Q`aP����Hm��{���J������u	ěa5��LHV�e�\�Cif��1(�<�!��C�҂�X�Gt�w��wvJ�VLO�d�WlEb�,$�*I
��
���ɧ���(���ɤ=�4ȳouu�I@�*AImZ�i�h�,���e���C}��,�E�B�ye1�Wb�DYr����(,ա�VB�>J�W �}By��6��i��Ҫ+�d��.]z�<��Y���M��MP�5�6�i���Y��r�4��RЬ��v�2bg&v��g�i���o��L*"}�{D�f�8Y�AAdQ=M�qPwg�]������ղ^RT/Kw|����'6k'�fR��o����3t<�5aS�s��c�m��=N&h�0{j-�'��N�GT���ϭ���d�6�f�S�]�I��Z�fv�0��<���4�Im*t�[c�c��lc��0�J�]V���mF
�f �lP{�0`��yg��켧�/u��gos�Fҡ����}�\�1��1'�TQ��d��}x��q�_=C=j�:��U�D��]XTY��]:�W�s��v�hE';t�(3ԥ�m*�1�S(V���E��P$
(��*��\�Ϸ���3�& ��0����h㬘�b��+6.Z���28�p�wn��7�g��s��O�����/R�e]��p�<��i��xh��2Zl�B��00Z��b)����}��^�3g-q<��
�����3����U�WY�t\�֧�q�'.�B�.�* �NUR��kK"�[�t��w��*��d6�Q�a�AboY���m]?e*�q(�=��뵞���£5{i>��ޣL�5��o쪫���M�hST�h�]�*(�$��"p�����#�%��ԬT�>1
$B�ٲ�ڸ��
$�d���?7�C�� �V�Q��[#�t��S���a���TA�Q��c5�i�\�/��$Z�5�9�lA��R�)ӫ �<x�1VӋ�EXN��WK$�I�4-��/�+�Yx��Y#g�ĊK���:�w]��I0DH�e0Z��@����Kc��E��VZN�J�zp��$P��Yj�0��e�V���2�Է��M��;*/K�%�!Fm��:k
g��B���}(6��(r����
��U�Y5:�h�*B	�(ڢ�4E�2�<gI�b'ۣ���pi�a�c��M\����m퇴`�4�޼6@ؖ�|��G3v�ʪ�ZBdbDB��j���r�'�6#Z�"�)Ӳ�H|n^��y�W(�HVP��E��,����
�D��9;kk�č?a��k2��fY�j���"���V�]���}޴�iWX��G�V���a��,#9�@=Z6}݈W�h��W�A#I*��Y@յ����y8�_	 ҵUc���R�aD�b��.�&iF��J�e:F$��q3X*Z����V�Q��ͳ�F@	�*���E�_vc�Agǁ����E2���������Dn	T��@i\�%a/�ΡdJ%��LY�祑J1�lƾ	[�iJ�;	=զ�ā��+U��w6,��rc���h�l�9R�]�ޒY^�|��h1���j�ae�Ǖt��Lz]e�2c�G_c�O �EB�\;fj����K݌�:厚QV��n>�����5���P�$�
�i�6>���o!���M����	A���֙���e�q뭡��'o�\������8Q��\�s�wm�	�E��DX?]�C\��lʝ�7>m����[�
u�*G�4^�X���$���D�UB����آ,Y(�j�w6��6�ƞ�hUPF`UR��C��D�zd��A�4 ��f�J���-;j����hb�����k��f%�� ����������S ��BaÌz��5:P��&�?$!��A��ySs1�̾4*�S��D/�b/��lP�r�;ʘ*U�okhKd
:�1ְ��j����/��b3Ƶ��\�{䡨�
jZ��`G.�T5P[T)S�7��.�n�Z�К�7e��0�G���(�B��������d��C
6��QWmX9�R��!��^ٱ(���1���#C��UJ�-����@Q�Y�����ľ�����������E"A�ԋ[��%Ź�� ��n�MYb�!T��h[7v�ʢ%9i��aʁ��nU�� x2�
"�Ѳ�*>`����4c�i�s�����q9d/�4m����S�rA�N���'1Q��w&��u`G���Xi�̉W�[�TL������C+���-Ee,"Mf�U6�q�Uv2�N���u�нCm�.4�v����\/��U+��,�#�pV\5B'l��(��M���o�#�e�԰Q	j
�y���+���m���A�	����fDj�UR�����{rZ�Maئ4�u��P���-��q���m��,&��� �c@]��j�|��q+&Vi�;r��f�2Œ�G�
���&��V��jO� (�a���'n��*��69�e+�Q\��"�č�ԫ0�LSWF�Sa�W���ma	_JA�6�a�-��Ě�������ʢ�^lhP[���2�L�!ٻQ��pPp=���F��f$4 ��ak��q�i�)���_�Z�8NU�<W�B����t��а,0'��7�v��kY�YRS�P�	�΃�h欃3�}^k��w;}��q���`�		'�?��n�����	����X���bM{H��T���F�B3z�M��qZ�wCG�<���R|��S���,��rl_>숓Ռo^���;��P���0�ɽf�ft��p��Y[yd��|��gaZ�q��X4�w��f�V-�w�:N=9���݉.�S�{����ov*�x����B\v��8sN�j��P�H��C3�����i�wn,�e=����"X���B/�d��f�����yim�Y+3�72]ڨ�Q�ºB���������M�t��z`�:J�|�ɮ�Of��P �TLf��of ���8�J�y�����b�X�_w>a��2�mK�ۉ��#+�ћ�NU-���V�7��	�  i�!� m����6� �L�@     Rl   �  r`    �M�6�         m�   �` L� �`�  6�     :D��Y��X�㝮�T����j�w��lm��[ܓ�Mv_9��7�n��\Gb�a�׬�\�x�NI�Wh+C+Q����#O\����GL#m�Ө�萋UH�M��.�D�����(#'va��ށ�5+�ή��|�!�hSڻT�8�z#M�&�66L
�3v�N���>f���*nڻ�GZ)�<5ܣ	�t�`Y��iz�$q�� �wri�Gtc���G`�&�n��?=��u�u���Nw�Y�����:7͊�0�W6�MR~����ez.�Ѥ��A�ۤ�}��   /ӳ�C=����u4��9��w�Z"�]��k;�\,�̦t����륡�I�R�[m�6�H   i 1�y%�Yn/�I;`�d�o&V#pp�n��Y�Ê��㷶�o>�8\����dI�>@��@�6��@� �3NI�`HBH��I ��H2w�!'�	4�I$6Ő;����'̇ �5�a2kz�$��Y'7����w�y��i�_��2*���(�QE�*�EX���"�Qb"�*��)ct(��DU"�E"���QAb�
��cE�:j��"�(�7�Q~j?5EUTTEEA,U�R*�EV>�r,TV0����u�F�*�E�b"�TE���V#A�j(y�Q`�,�*wW_�T���F+RR(�QPb
����+Ab�'�t�Q���1ED�EP��|�U�"�
�Sz�����B,UQEU�c1ATDdE`�TX�/;�ҩDQ����(*��Qb�@E�)DH������H����ϒX#�r�QQDDE�Tb(���#�j(21b$U(�����`�I��,E�θ.�U�O1��m����"����S���Eb��`��Ĩ�=h�DUQV,�PR,Db�?�E��7Lb1QE�B�QE<ƕ ���E��:�X�*(�,b�lU�*����b��1UAQTcmTX�*�`��;B�����f***"�QTQb�*�E"��e3��QQ��V"�1DTUX�Ec��5�<�Qb.���b1VV��ưU��*�����TDb��=�;�" �F*��)4ʤA�I�@$H9%]�sn�m�R=��v��_ы�ʋQD�EEN4X�D>uy�$�����h�PX�������+����b�b��(��6u�TEE`,��}h�,b�m�db,QE'YY�sZQ�TU"��A�h �DG���KJD�(�IQMZ(�N���;�,�,X�+�e����A��X�T�J$X�X("��",U\zɉm`�������ur�1TE�D5�Ć[�APQc���DR
H�����]m#�g���z�A��EET�-X,U���ᨱEX�������Z�,�Ԫ��
*��(��kh�F,L��
�z��*��X��r�����0TQY[`�387X������ª�
���hE���b�AE�ގ�*,b��Օ������*�Ҡ�(�޹�W��{_h��u��ͼLTD��1`��Ϯ,u��hTb�� ���Kg-�D�?w{�~J1c�SV�'(X�5U�=F*>tొ'�T�EQ�~�1b�1^��T��'ԧu��>�~j��n
�����
�	��O�D����}�bĿdN��L���E]�V��eb�DTO[�c8��PO��Z��*1�lw����j��+Ԡv؂z��,s��Ѹ�4دy�^l�v��NZ���b��
��T?%"&k��v.�U��F"�=s͸�J3�i�p�� �G�)�$W��6o�D]Ҡ��P�T�TEG��"��Q~�T�7�mբ�")׬ĢJ"���dwi�~��E:rOw�ѱX?��"of|�
�('Z� ���D�@| ����{�vfש(V Uo+1l:2����Q13�Z���ݶ�!���J#{�b���3�0����b�l�f�oSJ|���+�_��Ң'��FT?e5ZVO$�*Ŋ("(�Z���k�ѨH �x���$L7x��y�vo����v^{��� �A �]p]� �\�r�Q�*
��+��U~ߵ�L��!��kK?��Jsz�&l̨3��:�j1���f��Ў!\�b�b�ւ�~rr��w���6ٌG��m�^��[W�B<P9�nn��<:���N廳�-լ�w]:���/�;5p�,G��3�sC��ǜ	$D�Qܧi�.s7ݸ]�s��{��d]��)a���u�7T�kRW�A �H��"�UH�6�*��L��*���C��Q;KG��/�٥k�`�߽���(���S�ԟ}�_�����v�D������EQ�aEb�m���?v�c�U�wϧ����go}��:|�I�M�yf�cG����q�-��QG�K�(��7���щ�т��AS_�ڸ?9"+9|���C~����?n��{g-V(�{y����M������j3j�������aG�&���9i��U4}s/̚u�PX��elED}te�����SK���*���:W,v����u����2��k߾��E2۴2R�_q�C�8C#)RO{(��fpSy=��vot�)���"�憚�k&�%QN7�h�CJ�#�e��m*����<׉>泖��U�a�m�"&Xp��)�s{��ŀ�_���IA ����Sï�bt.Խ�����!Ӆ2�vu��:�v��f�4�_�9js�߻��g�V*��}����k�~�g�_�eX�y�g��fZq��!W��ưW���	���dʞ�2��1髻��]���1��t����C�w(���4�w5�;ݳֵ�ձ�濾���j����+i����;�����iX��ߩ�k��k̃��-o^8�,��m�Tf��T��n/H�A��I"�0G����䪳�ry����w_�%=�V��N�c��h��0\�������<�;Jfڊ��E H���Ltr/zU;F�����`�w�y��3���(*f;Ѥ��f���"�*/�Y�S�T�3�ٰ��~�߻���).�G��Mw�nO'Z��i�����~��Q#��.�M�^�4��+�
#�A>��4~�Qa����V�*��w?l냭��]}Cb$�v�4��1�~�U�9K��M�Q���W��n�o��B	"����O����k�[8�.M�'�̟4��9�>�O�uڧYD�g�T�i)Ģ"k_�4��+" ���F\q�!B�h�"�+��a`a�K�sRa�����u���	���YUJ`�3����6�n]�ծ�/~�JƓa�����-�a6z��e�y�]sd�T�Z=�D��{s�#;8�ᷘ9+PQ��i����� ΃Fs�5�r��p����^�R�#�c{u�� O�v��~�o�A���j.5MS8k�md���}�*�j��}�ۓlNY]�~-�q�n��׍NqY�T���ت*&�R��|{7���ٱulPS߯����Z�S!$��*#zz� jD$-�D���=u�e��~J�믵�Y���_~����M��л�����#�$T��N�J˧����_��F�	b<#<�2���PV�����q�O���m�V���E�������E;��ٶbu�`����v��K���}
ʤub�C���0�H��@���SZ����S(FK���G����g�A|O�P�Y�F�?%��]Z>l�{��e�y���oP�
#� �u{�(��A���ǘ(C!C�$���"���'��6a�>��s[??px,���_��1�K�U�;�2E\��N/,/ڹQ=��*}6�EI$np��u�cמI9].���}���ؚf��,G3��L�*]5�?F�g���.O߻��}e���sܫga��Xp�+W�l0�a�6�=�}��4��|��|hY��־#�~'�}�z�yZ��T�����-1����ك�X}C���8���Φz�5���Y{X\V��Q$����ϋ��9C,<:|��ީ�B�Z���^w�����-*�7�s^֘��n�/r�>��������{y�ʝe>ӟ�h����?��G���n�ƃ��B�v�#�}A|�-�~8���D��7��6!D�l�MwT\Lr]f+:��m�:\u���"*���u��{Wq6����n�(Ǟ�.��H����-�.�'Y�x�>�S֪�9����̏��q���_��U4s	���������hk�(��-(� F��Ѣ�*S�V������3T$X�y$�z{a�&X�nr�dK��)����J��(���aW�#���ߢ@�Z�]'�7�&'����ּ'&��Ep�uq-��b;�n�!��\�ݹoaA�z��ϗ� ���{�h��*+V��;���8O�~�m���l�_"�ō�$#���T�Q��{z�!dZ\@E:�����������N�uM�ܠ��w����+փ� x[do�`�����26��"�0��#�A��A֐��uV��K�^���T�2$�~Ye��� )N�"�{�2YE����'�H�>,�D!�P�͚eV~��Ώ��5�~ʌ{j��1����~�!�tkZn�e���g��{׵�h���-_a���#L����?+�6�W�qSMzw_�;,E5J�2�o�6�}�ַ�s��+:�w������lqY �V���6�Π���n��_Č�ǒ��)?����͵{i��Vs�׷|��C�"�zI�&,
'z֥��7���N�z4��MY�LqW��=��i�V�s~R�ͩ@e�k�P�����}�����c�_K�T��$�d	j�2t~"s{{O�v�����P#
���:#�P���wd�Y���1@|��Uٞ�s\���u����I�>�F,�����\�_߳����>�x�H��O��a��Њ�.o,���vw�Q��(�#O��퉮k�5?2���[=J�����]��n�;����L�4�6!���P�����<I^���]J�����':� �BbkB���j��}8�@@�y��	"���Z�E������~����K4�k�:�Vk��b�c�MJ͜O�ok���}�d�P�H�l�l)h���1�ݠ�h	����Mj�||guv�y�n��ľ ���^�_H��I�]�/0?�Q�M����u@!/�7����L�+����8VO��]�jU��D���M\����݁t���N�[3d�����1ٷ����ml��:�z��dܥP�61��dk�d@�Ne���m�  � I�����z[1�v���{���u>v;�Z�A�=]��"�ē��iI��g<|bT3k��Z͸��{ݚ��X��?Y�Y�m���i0Z~9*�|���"&Ry9�
_'�����s���]��ɥ����k�rs��k�r>w-����`�B��z[�hx��"�=aY�v���|(y\#���UF��yn�|oH���������|� bƉ��~?A�$�-/-�����@Y�D@�Rz���a��t�Nd�y�E^y��[@�AŪy]�+��J��_�qy�N�ʈG�Iz��M�~�V�x�@��׼���*O�iעÃ�����{�B������a�]u�z!��h���Q�v�m�)�n�~f�í$d8�P��O��؏kk��巹'-�:B�"�6�៼l��Z 1��y.HK�b����e5��>mG�"Y
�6���-6v#�֟���~)����<�P�*ՠ��{��wƩb=��5;t&(ƿ��N7��pCF�8^S�N(Ί���[�1fC�V���L@{�>�������F�&y��L�M�z_`��@����쨡�9�`�z�x��$Po��f�v�[��Xv��ߋ����Dl�5���YT	#��D~�X	x�3�g
��Mt�Q$�n?��yn,���>���y��]����w�!�y�>8�k���h~d+iZ
�=��D5o�2/�sΚ�V &�b�`�����"��7�BV�=[aO����߾�����Hq y!	��y�6����@9E�@Ą��@4��@�'P�a�@� iq�^���@�Br���$v�$���@��u�Ha&�!���XO!%@3��Pհޯ�VI	PI��XO�q�H}�� Ձ	�!=��Yﵭ}���I[M ��y�WD�V3�HSTvs�9�Y�y&�*M��s�D��0t�B���۷����� �hPV��Ú8t��"�\��6�����IP�1mRɴk��5t	����~zrG�;���k�X��x[���9P�*xUtL�a"� ��L�_Y�bՔ6��P;C� �� ���A�ʢ;�({�O���~�{v�8qw�G�A"�u�Z��!a�Lj���ۑ+1аP�d+4�o1��I��N�?1�Uy?U�1]�D�/v3��\Ըד�_�F�b'��D��CK49?�&��4ҭ$��J��a}� g��x}W���g���vަ�����~i|����^�ʊ�7�</=�	��3�+�"�_;^3��k�� �5�����]��O�ԋ�ƕ� 0e�'�~�_P�� ���Ӎi"`����@���4�����'r]�*^�>D*$����wZ�:�М�s�w��� �(Q��*�-�޽c�f����L�S&M����n�Z+�1TO=�IPK��s�h3�oc�b?q�
���7�=M�,"��XT��k��lYֈ�R�%�i X�7w$�o�{���p53�c\Cs*����D����F��b�
�*��G�_�1Ly�:���A�s��]�<�����u�Ͻ�y޼|�7��Nť2�"ʋ�h�l����_(�R�ؘV����#0>&
s^�.���%j�~��M]�j�;������ ��^��$��,��$������@�9���I�gQ{��k!?z����S�ٶ��h6��N"��x@7�ހ�^�;ݛ��X/RO��=��0����٧���k��~��?�~9��Hz����4����ގ��Ix���\ �������̣���2;{��h�*��^��럣�A�޾yT��[��e(S$�8�.�$;΃���̿��\"���yy�$�z�1R�q���N<�^R.�N�S�#m�,�!`D\�_�|ѡID�H�CE��\5��=O S4)���׶�3����<i!)�;�F��M�}��h�j�:�F�&��廣d�jI����D�הL����8��^�Y��kѩ�C���g�P�pZ,����C1��|3��<Z�ɀ���ߩ�+�7���
�\�UM�hAB4���X�����,څ����6l�~M���!k�$�Ƈ8����m�^�6i�nW!Fk"�m("��zh*4�lˈ/r��"��?kS�.v�ֲ(:�q,�.��Q��H'ެ�P���3/v���6�?�-P
���bhRceҧ+�	 ���3�e}ƀ��b�(D�b¯��X�g�w�gܦ��N�$�$/��.��Y�D�	B��6@��vE�v��̘��/��5������7��)ӻ�����NS$O&	����%��>���XCHe2��A�ÍH�/��^�0*U�7>D����ݱȕZ�"������$�G*�g�Ki�Y"����T���* ������8��� �\��.ad�i�~�v�����e��7�O����a�ͳz2��궲�ə�������M�P��WKF�(�w05%�z�c{[�{��x���Cƥ	�X���!Մ���H���L�� �y�F���4������
໯�~�X�}���a���<y���ɛ��ת��l.x@c�ܻ�i;5�E���^��E׍_��^2�� � ;��2�"RWO�
{3(3�
�Y�>���cܓ��A�v:�=�M�5�n�,�mA�@@���T�Ɩ�7ޡfG�qfͮ��u`���3���˷j�TRn!ZùcK��_Y7t7O�ő󩎁��{T�ճ/�("0���CjA�֛9|4]g�a}���2�e�:i�s7)~Ɇ$�l��6k��Z�Q���48���#�]�Wu
��7������ş�[�z��O>�f�]Q�U�u�c<�!�F�Cf�}O��0�"	�/u�b��n���"���9��3w&ë��qaw��u��N��^��=qE#�Pq��W���t����t�d���>D�ch�i�$���d����>Tny͛^�{���De{}4]c�t���*[��k��"��
#��O�hU��i� ���|Ю��Z�#8��M�$v���HI�b�=� �1��Gت���L�Mk$d�݇V��~�am��a��������r�?��A`�E���@��7��wze,�Ez�R����D�;TI�49m>���˭ya�3(���Z�L��#`ެѭP��/$f�W�˖��ݣ�:�1k&���ҢrZ�����lV�r����Vaպ�U�|2��7(*F�w.R<5��:k����݄`��nF�2  6�      �W�l=� �JH�)��p�ҍ*x�8ggKؕ���tm(C� o�5��:�Ưn0��&dk���~$^ۡf�@)�[Wܳ�IN[Y���b>�^{����Ք�`�ɣw�R�ek��s$�Jh*$!��vv�e/"�ܦ ����f�V���<O��4��1U�||��.<~��^B���|���� ��9X��N��ZkG��Oi�96�ʶ���8֌�*;cٔ��~˺��������Oǚ:���/$�Dw`󽿢h<>�x��[��x�P�#���^�WÄ��t�����<�A�sXF�_�o�B�\J�(u�N�����/(gd���N�g���@�@|wy�Utu֟��,^g��������+:w��H�NWvc��3��^��{�
�[��@�Q�b�+^0�N�%&����ޛ���'̆��o�q����1�w_d�y�sb���89��|��T��;�t��s!�1B$��s7N������-�M�ͺ� ��֍YA����ޝL�}��x��U3��|L���6l�Q�7�_��ʞK�p��f�%��$%�V�Ϝ���$�5U��TQ�ށ���+�=�H��Ũ�Ra����vU~ۚ��{��#���|�YA��ɪ!-�SN:I�u��;j��+�Z�݂���<z����V�⣊��3�q�q�j��]��Et��¹�d�yQ΢�Rՙ�����GX���[:_E�m���^n��#�X]X�o5��_��7�2��k��WJ�� �+7ޖ0pV\�B�Y�v�>���["Q�����L��^��
g�yf��1~<{|<�Y���>�Z3��V�ޞ؝U�Bm�Lr�t%۸�:u"}��NɊ�y�~(Gՙ]�⟲#���{a��B�Ϩy���eN�����y6��5��U��%c �����{o΂5ʝ���}�T=L>н�K��Xld:�u0]�k~~��N���E����{N'=U�4�ȢI�Y_3u�wM�DXfٴ��jE��mz��4�/$����̣Ƶ�JϹ��F���s�[�ٝ�7�89�K�D���b�%o�����?���u�4]���/�'8��f�!�[�M:49 lm�Ȕ�lO2��tz����
���܊r^��F���"��[�	Γ��u�:�=��ς�)�&���Rm��������Q&�^qhS�Jyv$E�Q�D�h�*�&�:7�9���6���~b�~�MͿl����c[��[=�^��b9#{�؆Í���*�a,��dS��z����L	�:����^����:V�d�.�Ϲ�589|>�?���``N�T 'NP��!Y~�  ��G>7��Y��8`��fjU�Z�n޺ڻ�f��g@�$R�'��;WVj����յ���}(:9h��&ε������1ed��u�rq�k{��̥�4�����gC���˅ޮ䰣��)��c�J�n��%�D'R8d��d9H�o��r�3��H:�ZA��:��W��o_v����d�����Y728���eB�~���L��0X��q@�h(�#��©ƗOxw���gDW��/ذ�{Ԛ�|��J]Y��ޓJ����n��Ή�)5�*�yR�1}�
����[K���*��V���a�L�;^sj�����x'/�E�����S{ka'��hͳ牻l�D!STU��>�o0����Αq�R�sԖo5��W�"�HU�	[Hغ<�Zr���t���+;Aἂ���'sswMBǼB��~����A��u��*K�ݝ��C��7ק�4IJ�k���drޮ�h�}��f��f�hc&���]�E]�� �I���9�f�`�a5�n�s�xs�����]�j��v=��YRt!�k:p�R�X��\,��2�\�;ۡ�L��wkw�ĸ�@�}p�	�q��ڝ��lO6J��|En�_P�Q;�r�U��d�RWНi��M�`B�i�7���n�������*��k���[zhk��Ɗk"΢�D�4a.�8���U���`ce�P��7N}�%�(X[Ɯ��R��cY�])�B:��n,UӍ�5�Z�Ϧ�]�ml|8���#�f��/�K]��y}t����k������k�;���h��y$�Ddܻ]ǖ����ۉ!gU��N��qܷ�oQ��ؙE��.��q�Z�[	���]��SJ�w�֫X6fe/�œScA��<r��㻿�����s���
!# �
9wuq����'���%�7��|ym�����gC�aU�i��~'
�HFqµ�vդ�v&�Gk3Um�>��LJ����/�j��juXSV��S�U*�TCS���ڼ�0�g8�=�4�[ w:�����}�ڲ��{�l?f^c#Xx2J���N�I{&d�Q�ú���[�3��˝˵n�f�ui�q�'��;�/��:�K�{�O���=h��sy��-�8 ��ͺ2/�@ʩ�,�,�'�=����|ԙ��{��r�1đwJ�^�x�o������?dh�c�f�_ab�O�]: YW�?���~%��9�ceȗ'i�n�1�����6��*��>����-�.�O�>���#.�g�]�� �a�p���X�K7h\˗�t���2A�Ez��9��d-��!/��.Ϸ��ueW$]kC���	�1�1�j��.y_f�an�������
Q3����.�߱fE����J$�l�d�W3�܎Y̚ohM�pbYc�8(�k �Xe�

�ؚ/�f~�P}�E��KDN� �g�zF;IK١������>��6`6��<��3LWSwt��'��F Wz�Q��k�#��ۦU�+�B���o��냭�4$.y�7�<�q6Pm�(�O�=�j=!����JFDn�"^m95���,KK�x�Mf�p�+�����1S�)>�����i��t�1�&[׽X:�{^dP�^i�>���Il�q:)0�}�(ԣ�X]H����?K�aYF'7��+S��tm�U���I?����[����1�����.�8[�Lƣ\fG��O�Ò/V]���UA�n��'-?'@ϼ6}��+x��K��qAGd���}�U�l<��V�0D�n���`�}�f$}*B�0��}�+����=Uq�4l8Ȁ'ʲ�"�;A��	���jvn�+u��r%��5U����v�x�.;O��r���]y��6�����f�u�:�ڜu��89�U�]��{�C�b���"����:�GZ}�?�TXϚ?h�s�ۺ������{'qt�0����d��+���� G5�D�L}�Ŋ��
�K\R�Z1!@m�f�_l��؃�G��ٹ��=-$���&����ky�EK��~� ���6�P�֜E�fǕs����.;���od=���0ŷΞwM:���B>�g�����
�mb����D[\4�;,��3�\�7Ԁ�=����.��2,��S��y�Ҽ�2|�Ɯ۰�z�����2T��
o*D��.�Hc�MAtp?o����,��&��ͤ�HUB��`����Ǡ'�;v�Ί�^r�	Q뎻ʺ������3S�dff�s�V��u�"$�'鲹ٻ��~Q��|z�U�	Fr�>5��+�Gn:�5�dA֢8�,W6�Vz��v��Nv�4�k��Y�K��w\�]�a��1W����W�Ɇ�P�R���}2�f�׫����
��ٙS<4!�Ԯ4���!"n��E�F�^��5H�zq���)f��0�]��ܚvn�X����0d�.��zŏ�uB���hw	d]˂|�Ix�#�5�*;�2I�*���(��k�����rm���~E����x�Xb�B{
?fM&2y��&�
�R�>�}ϳz҇��?RT��\�G�G�����ze1U[�η9�.�zY�N��K��5G������/�������`�w(N�������ׅ
_��@�?t�����|;O�¡�i��T}5�41�w%]:V��Y�h$��$��      m�  ��ſ� �$ե�P��n�)��[�ʗ��qM�ݡv*�������_'���'�y���g?nC�8�S9�jJ�m1)ϰ4��2m7�Nv�v��O���D�?�?�ڲ��A��Qf%Da~�`k���4�#�R>Q���g�	����#���s�&٦E��L���~M�+6o9��$6��w_���*���h�ģ�qV�9��:��L��ԝ����M�&����K��^���s{�RP�T2�t�#/������{t��C����)י@���Oox�LjxLe��&��uii�hAc�&o�8�`s�}��
�?R�N'Z����î~��ͮlL�߽�f�0���I��I<��F:��`�B���ܑ}ɸ�۩��WA��划/ewSc#�,B�Mz��Y}s�H�2gU�'��kc��n� �������B�ma2*7��쿳$�(|�ϝ!��L4����]�k�}��&j����B,q�m�����S�og'%Z�]Ac腗n C�C�:ϐy�����i���cFw�Ηz�X|�a��4���!�ovAI�IShM�<�o |ì�,ٜ��ϐ�)�M�I��'��H�x�m<���CkQ&_��55k����-�:[�<�U��ń�Vg0"~��}N\a�F"�&����'�J��ŝ�f����w��gg�S���>��� rJdC�Qgo������� ���d�����y�J�G�G���q,Օ<:@�X�Xj�a��q�u.�w_�,��M}�>N���(=�i���S�Ov���/S�_ Ȅ~�n��n5��ߦF�B��m�Iy)��ADu�����D騌3�?';gR|�@�o7�M���=�m�b~z�:����6���
$���6���o���H,R�̿$��a�w��C{��<��=�dP�1n+yI�9��٭z+�R��A��������O�?�����M�@�|�'����!֠,�w��6�2��k��`{t�,&}�_�9	Ԭ���W����6�'�Y3�2a�\���E)$i�Y����wՋ���!j��	Yh]KР�=j��S&�¬��,fh[�L��5����R���D9s��c�?�f%��G�o����뾣��oM��Dvw6k����rs���֠�=�.���ک�r��T��K�E3vgG�����h�ٹ������w���A�}���~8�?�sP?0:�����'�%C�����'�S�Sy0�m�n{n��0?������M��B��O���|�C��?	P<@溾'��G�zY[�]�u��������%y~��<�������&���~ўx�z釒~�B�4�}��WLR��g�4~��{ Ro��z0�Y:���a�Ȁȣ�::�z귑���K�/���C�O�L?�|�`}�g�6��S_Xz�3�|���b?�3����m������E����gWng���0,X���#�j�ךaF	��o��s/�/(|�>�P����/��9��������o{�8`�ݭ�ܛ�"���P9=2V�쿜xn�ۋS9G�j���|"F��6���Tz�GW�؋�̹��6i�	э���n�nz��O�������C]�ûdv�Fa��u�3b�:�;�����p�[�#y����Q^ԁ"KpZ����RgX=�O�l7=H���J��m����*��]eyH0a��D)��q�����UF=��xv�:�"n�Ъ�P�*ha�6��I3;��/w��'�����<�__����-���X[�ޫ��ģ}j3�S�:�4G)�Ou<����c�b�/x��Ǻ�Cs�yEf_ϒ�~fAELݦ�x��}�ׂ�/㖫�@�v��;�6� �,v��B�͞�c�
� 3�"5ԥI��B9� @��yu�q}��Bٹ�{c�C�O�ܰ�6Pٱo�޵�����(�bn�e���������u��T�;n�$G*І>�MKk.%ȍ�:jTF(�G(����6<�5���Goe�Ŝf��UO~�Տ/i.:����pG+E�����SE�Ԑ�M���n<�1�Q���Y��.r�Pc�p��s{$!q�%���"2�2gk���v����j	"6D��mG�m�I��"��Y�J�W�E�K�+��SuH������V#I��X<�]>���2�$�6f�܁pD������SJD��=
���%����xFT��gy�ў�n����t�:�`��6БEWk0�dכ�ؐ�v{��������c9R�BU�[ �tv�I��H��9	>�&��h֫O�#UWWul�������,�t�N�%%-�C��(�B6�v��]_*��N�
�oɈ���5įgD1���]R1^W-���u�ȥ���d���
�b}aG�\�U������'����1��P��z��M����E]�s�P08aV�����*��� �n�e1{=H�p��\;�~����Z�٫s"-�8��1f�fK�f!��:����EF�>��upm.�vGb�@����-ю�2�y$t�{��D�3�v� �n��e�MT�=�/������_��N'��46;Ф����'�T�s�5].�P���W��r��Rw�u)黃q���7����E�[β�:2?z}[��W|�;Y��U#�v�:�|J��8��H	�=�U�����3W3�~��|tfk���~	B�2�Z� �iE���:�6�i���5Ѕ�'ЯL�M85%�k	�Mu��`���&��7�U�3��τo��d�a���Gz�	;��f�.�%pﺄ�b��|�C�9ͥV�7�5��;��.h{�v7&���C�Ϳ���D�T^%lWl�=����ʢH��}���/F��C�BeX���O��5�8��ވ�A��?���=����X��i13�2Wk�;m��]�2���z��/��>�K/�PNb��Z�Ш��L(c�ﺼ����\��f�`�ϫ�F�����~��뛜9uΗ��2��}��@��^�A�]�k)T�UO8�3mPR������x�{�IE,�Y�>����=�"zb�1�,)�[;��U�����q^�u��}�&}�iOu�Hd[람���"*�zP;2Ǯh� ��B����F�pŗ&�5k=�Ov��O��`�@�6��U���pvE�wmv��ה�NuY
�3C�+\�e�=�Nȟ�[�Û�?���/�L����z��?(1��{�Ouw������$�̥�"�U镞14YR3�fյ�7�YQ<��ybSg�������>1V'�����duz�F�b����&���=�QX��e:VA��iҥ zPuv8N`�>C�GF�s5\��\���^�<E��DA����r��.�F�j2�5eG�F�{`���z�>y��|�i�%>`�����tx�� �G#.��0��z�囑���~���1l]7�[��b+lD�N�$��yd�ҽRD����H�an�2�`����ݪ�l\ΰ8���}��]����q��W=ƻu�_G=H`�s-��4�       A�&?��VI쩫�V����K[�A]�$+�=�I�O���m&�D�W�Iu����ExsV3o���|ӯ-����ao�۝�"HYk$�a���␝N8K�o�f��|+���Ayv��xxW�`��gc����H����a��0 ƠG5�m�����c�Z~ۘ�u�
=��KP۟	=!����AH��a/\�F�p�����$v��r3mKH�x<�5����spM�D���і�e=[�_�O	����	�f��*�S���Ia�6��N���bp�QW�ݪ��|����=ڔ���i˞�|&Ü쫎���hY"TlV7+oLy���4�9�%�}a%���:ߨJ���2 :����H:����b�X��\Kg�Bw۷d��QӘ/|�cz��7�(�ů[|��}UT��6a��j�����t+�-�q�0��t�̣���c���^���䭁���F��]N8�DF�`�Q3�=J��?A��+cg��Y#�'��
?be�GVF|1~;^1P���G�_�#/ڕ´0&�����7K��{�?	RWW���p!n�̓rU��?rU9յ^�������):���~��.���ws{~ɉ����bä���+f�(QU��Qg-����y2�}ֹ)��u���
���cs<��Vj���w�gq�ֻ�ZCr踫��+z��}�f��K��Νu)q`\�lΒT�UH!�Ly�N�|�\^e7U���u��]C]�k�Z�F�N�R��vm��r.ŷu��i���F�h����;h�(,�t�X�3fgL�0v��4Fg��h�6(�vrTu쭗�A��*����ݚ��ܜ�M��ќ< �G2]�"H�h����ĳb��iI>�����*����9�j_�*��QIS��lo�֏�Zc����%�{�"剫Ӟ�"��3��U��/x��E1s>5��bLYM��D��za�zY�Z~T����sp�CL��S�=w��� ��s~PD�,v���iG䐏O�Y{��2Y���l�.�]1�u������=p�>y'"�+K�.���=�h����έ6A%���&_f����-�N�j��^���7��*�Lz-��Q$�ҽ)vbvH�U�*I�*��)B��q����)WcvW�n��'�!����f��Im�,��3S\w�0Ƙ�4-S���:i{}E���hujy�=�N��-�����q� �G�#��ܭ�uR�}z��$��F��X�`ڎ闢=^7�U�by��E��X�9Ub�Ri�Lg���]my����e�I����fO�͘��	q����k���o��u�뢲�`pK��1��s�c.�c9J�O�gو��}��O*M�yϫ�l�}��CU_�����q<��;�o�G�ۡ��-��ю�vgPU���˾��o��eg�]��_!]��>&^mE�T��<%�����j��V�sqh8T��pt2jZ���ᷙ�MXjt�KU��Z�.�"�.9�Q3&s������w~mU�J�\ݫ�m	Ժ��a� Vn�O�ۤo�f����h�9���.8�6R��m��=~��$�B�~���h�..�e�k�5�b���֚��T�BݺF'���0�����"-���en�����Ѱ��a�6vX6gv��omg��^�
!㾡��(���"\�5@����\w�E�*{0��ϝ�WQ�fb.N*�fb������L����fmd%K��|�W�W���ݷ��Q�whNl$�ݯ��r�LăD�v�����S��t��I�ll ����wO~�-��M�\�ώ���T�D��H��
�<�vu�cy2'+��(�jB��x�U+�*���J������ɒ㻏h����b�. �~��x��1D�௺��bm��3F<y8��[��=�FyK�P�k����=�E��]�j�v�6���4q�D�Q��'�mߢ�3y��3Y$A����g4=���Ѳ�vF�6�2i_���������k���u��snO��d#2���ࡋ���g��@}؄;�S�����Ff��DH�W�Eb2g:�֌
����ٹ�=8`�k:�R�`��=�����z���\�C?]mˁ��M<��\���D;��"x%i���/a�X:)�)	5/A�Sɼ����2ط�r����1v�S��[�/�޾������he��M=.�cLi�[��O[�k/U��-�ܸv��â׼�HȓK�n	��;����Wtu�D��e(+�d�	�H�� ��bފ���M�:��Lѫ�i�+��5�����)-�����P]3�aj����|r�#���7�/�q�oe����x���j�^�|���Z�~K�$�������ϠÎ���D���Pu�TZ` a�� �Ɛ�FK�u~9�7%����+����I�*-��L�����B�0��y\���7cՕ�sl�P������fRD@]	��N�����[4E9U=f\#YWq�n�c��I�U>xk~vW�Ju$\6�S@�^�X��F�o��|y��IMo�Y����\�� ]u�Z���f�Q�靓��Er^�\�fg�} ؋R�}��ƻ�1��*훛�Zt<e�/����qr�Uy��l�r��t�V�A��l`��=���r ���\+�m�<`u��<�-f���L2h�^�z����'�6'�y�̚:�̯uCZ�Fs��!��jH9����R�>��C���V�^�Q�J:>f��{�ݚ���mo)3�|Є,@F{��&��$,�^����+(��lx��oS��r-@��hj:&y��
���E�whV6_�j�C2�p�
�a�/whN-�fn:r�H�ëzv�O��:ż�}U�GIC=A2�i���k�P}s2J]Y6�]?s�v�۔Lg�x_f*�ݦ���u���&W�=DLf/�
��0�|��ި��t��@�9Z�]8�͎[�1!3	���Un��ٚ���4$� ��9e����kw���9Sv����#t����G��fH{��q�
�#*���֌]����iDU�t�]��������ď�N>s�{u�x�ƶ-U/D�n�ɡs����нˑ]��P}Ƚ4��d��Uf���y�QT�Fo5)E�l[��2n-N-��s&_gpU�e�U�e��޾N���8���ф��6�ݱ 4ET�s�vu����cm�_^Ump�Ds�g����5�{l&$�Ą�&�I_s�8몔�|�D��G˞�T�_i}��+<���`5ݢ9�q��"���栞�y���;��J�0n{%�>k0q�i��A�ovʐ�;i�ܐ���T�;�z�k�Cn��p��`
R��H�f�s���w�w��v�\Ds�]ND���K0��v�SX���w,	�i�#�Z��\X��)c ��EJl6����Ѿ���:s.�v 	�V{Y--sF�i��~y��Ƞו㘶֛�ud����`v��;�61ø�7�nIj��/�*���J�v�їݦ�ݠp���W}-��Fd1�Nlŉ����f]��р��nk�9gfr��5\h�W�ݜ?����>�]�}��W׋���M��ut�uX�a,�������@��D�;e`����B�K��̬�]����^:�X�L{n���YnA���ݜ~�}4V�����g�!땆@c@.Q���o���-��U�f�[��}7��s�+V�l������I�S�;|CufE7�j�#tl���[#���7��,iM8̮o��ق4� ���cՙ�1$�c���3�=)h#6�,�_�-�G�%Ӕ�R�1m��O�L��rV�)M1%�F�_[���fly�1)����w�Gƺ+�Gm�}����SֺZvwz�K�ə���fSWkH'�F�&�c|�̊�wY�A42%Xs�����ԍ��63D�}݇[{�5y��Me�U�7�T�e����ԧ�f���.��t��J���F����������3%U���z�9X���3��sx��͞��/A�4�cm�lI6�4�`  �  �`�   72&     BM�l�6  lm��  $�$    �  �` 6�  �`     �             S3f�+�
��ӧ�O��L���Q�a=ohd�,�,�ݼ�vT��	���η��J�3}�z�:��9XW��pl�PWTg�z E>�6U� ��ze���L2�I4I�� ����b~sy��5q�:�z9?<�ͥ7�Xڦ���  I5*�/Gfen���}�^��˱� ]C���ұ �WR�����ݘ9��1���tU���v��m��=�����M,��,�+6ͱMت�|�Ӹ�e�y]���lw�ɎӣǑ[�K��-�s�Z�5���c3���D}�U��,äf�5:���r�d#Ig�m=�`�y��9t�j�Y�3�$�$�s3#m��`     �`��ٌ��ՕJ-�J7@��v�#r�յ���#�t,�  P۫���������.<�bV�~�W~��YG�h��R��#Q��{w�us�y"3qs���uI/��m�E���g3w�/?� �����Q^   ��MN*�����U��>[YD7|#k<q�#`-�vw�MF��P� ��i���?H��ϟ�a7W����ba�k��R]e�=����z�i���lvDR��m҉���^�b���y�bj}-�۩܏�#��֫ �v��u�T�<�D�����>���kU������@��U�۽��)QH�7{���D���y�7X�g�f�^��M�1n䖔��;zN=5�.���4��/���].�'Xe�
���!���m̮���J�A��f!_���r^�xr#��/�f�E̒`zۜ<Dӭ��m_=�8]�n	�Xޛ�Po�MbUi*�>���Ꙧ�&Tr�`ڇa=�a�0�r����n�u���G�'(ι��,���1�j�j̍�B^N�,�nK���Z]�!�4iC��zمRm��]����uj���9�۰6�^�������V�K�UP^H��a���Ch��䞅�J��8���{��9Q��R��?����W�\li�R4�8�J���Lmp�����>�ʑ�PBTϧ�\�N�1j�nCNuǜ�q�kf��.���Mm̿���Lu�D��l��M`��⥅Z���<�vU�y���c0����+52�bWC&dZm�馜{��;3M�Z��!�����������;g6���jW�ɷ�^�boV*��U"f
���u�`S�����r�}���鮽��J��I��V`왌���5]6�7�\������"���d��dI�I��3�idj�Ea_w^fJĝQ-��6��1�ջӚcz��Q˻u���B� �7�d�t�<���d8��SD ���p�S�T$��7�t��iY�T-��#-?0^�}SϺ��\���	xְ������M.u�Z��N*��"���q^�MJ窵�P5O��x�-��BV\
��E�?�s��c�܏*� �.���4��=�Zc�֏Z�� �].�Q�~��U�e[��մ4l?�r�}�x��|�$i�Nx������k�;�;W����h*�H�*0��*�H(92j����6�WK�)g�W�b_��	x1��kJ7u��đR�!Ⱘ\�^;�PV�e�M˧��|J�-qe����OJ,��O��[�-_��N�n$��eh����s�Xp���)��KDrMo������ir����*=L$F��X�-�ȮRFJS�m���tr/.]�����7tA"�R���@��	��U��9Yaq�ȱ�ٞ�����s��B���k�|uS}�]��3ꮫ������~�$܍�#j'���3�[�1�"���V��-�G�팥>T�CI(Z`ŪmM�N֧z�9�l���7.��F�RY�M��N��vҸ��tȡl���9��=��;N�_	YJ>8��#�V�;��)��M�,��"��h��P*�i;�GQΝH��(�1vM+E�O��}�TWg;n�.�5˱FћQ]ƕ�O%㟳��`�Z���D.U�J�x�M�G��V��׺�
�
��D/�ហ>�ܨs;5[K� ��T�w�B�-^g�`�(�L�jeݐ��{x��W���h�$�E�����̷���|&L�5��>p�e,���s���aS�����94�-�yij�Һ��5EDN��8:�C^�[bP���s�^�K`����AS'ީr��O�XiOz���M�:�q�y�9ib멹_,������@T.��"�}��oC6�ZNݦ�� ������f�|D��<�7+T�NB.�J�4�N��ם����V�p�9���b��3�VEY�O�?W���Y������  ��*�?����Ϊ��$��Sd���0�M9�C�15�T������P�NL����b7sP�Q�_��,{])��<���X��p���g�z��Uh4�h1SM������	��\�M@q��䪞�]�{�M����Y9�"�v����z����:�[Z46�ԁa�M
��.f�L�QwR�"��G���A�1^oUF_�4��	Q������ܗB�a�yP��!��fEߞ����.�T�RV�^Q= ��$�J
�x#n:�{����q�>�fk��n1�������W��#R�f�-V1�r��[��W3���Q˥�˵�}Iձ��n�+fN�y��T��iE�&A��f*Q�SZ{W�5�)K]��8oFp��C�I����8wݕp]@�JXF����tLV��⩐tZ<�'(��_��q�ZO�E�-�����; X������x���hbQ�>����φ��{pE]�xb+����gV�U��+�P0E�|�ۑoU��4%�y��_�wF=��+=p&y?���!�����JO��t,�����c.*FT�������]N�(CyuU`��M���j�ʃ�]>*��e2z���ϟG��}ы��x��ޅp���[�T��\��\L
������kw��G�u�X���(���6l8"�j=����]m"o'��~�����^_���O�����'g[�g6��S'^^�k�i��/;��D���J�A��Zw-a�u�ށ�P�1���������)ꈞ���%%K^Rv��5��'�7Of㯍Y�N�3|�0C��I䥞�.� M\�l�d�a��a��IJ�<O���r:<��kr4˩=/t���ȥ�y�>�%��m���$����m�[�ײG���j����ͅ7g��7��.�ˉx'"��-c�j!>#ue\��P��[�d绱خ�qK�A��޲�%T���x�Sм//��hw�n\�%����{����:1�[�����0�b�"�0è`*��޻��x&��ִ���S�e���;;�4�J���˩�#�3���+����{������|�$�b	� m����  ��h�ۚ
�F�彊R�߮7��S���q��%�N���+�v�y� %�4ꇌ�h��ʃ�ɚ�]��J�2���<��M��� ���z�a������.�tS7��)��c�2���M���ګ�Wy�n/��uu�8�'~��NrF�y�Y���A�c��.b��L��ʌ�m'�3�i�|�x�{�\1�P.�@��L�y5��9Tn!{,`�1��}OMx�+�}�)ĳ>>��`�S��ZP��d��5_�~=�DllaR �ʷ>> �px��j+ݚ��z��J܇���|��nEM3@�ވv��_(�K]VuPfࢆ cZ������Q"���،g�����hnC��x�y"��!l	��AX'O�2�]��|wjC������KOΊn��x��e Px�IX��({L�]��S:��m�M��u�]mP��q�����|&&r���N�v�>��iX.��P��z����!-�h8���n���r���}n�4V�����͜�>]2PP`��蚵n:��Σ��]l�7m�m�i8pb���w�}B�M(+�P#������k����]w,4��Q�Z�j�L����<ЮҚf��0�6m�4YuԆ��Q��mGB�W�*��<1�f�*
e13j�����T'k�*"6�~!�rb�&Q|��G�9M1��U�a<ƽ��B%��cM�S��jӗC�e�ǟ��5�殞�3��We��^ �Cw��B�-����h9��ѕ���x���=!�?a
h����V��PZoz���[!�Õ���J�v�$+���zdQ��_{w�/��~*�UŲ5�z�kFldV�L��#����-n���<kMf�;�X��1ea#U<�k>�`8�k���ދ�L��y(z���w��E.�c����ݷ���Ws�d9pX&��H�u3@贉��2%�)�>>�۞ٹ�N�Ծ@0���eԒ<	��B��|����vI��`���Pu��E^T�IVx����N3Qs����uU�/�e�G R�)3RRf��l�C �P�3s��?Sn#���_�zwݺq�I�u;zw���m£��#4t!�㧕�T͔��y���K�w/"�z�[�z�����J�]�&��]��ͥ3��K��ǇǃF�(,g�D����d�9/	�ݛ�l��)d�:Bh�Uq��"6}6�m�M��KT��jq$ߪ�;5nZ� ����&�I-�6肕�AF_��"\-���<�o���3���yO2���_�T��gBˆ�����z��	{QZ��ʧ�	ʉ,��}/ܑ��$��Z�fn��y7�.�h��ɜ�<��\hc��c#�yGA�� �[{2��#gm
4f�R�blUع{�0��Qicx:"b
�ynx��M�卜��֝3ZQ����IS��}���ǋq��(�j`֦O�&U4���l�>�Z�~ҫ��@9�c󾿽��o^�|�l�J|����=u9T��L��%����ȝ��W^�{o��c�-�/n���.u�7S�|�o7�HQ�]z��5?E8�X�=��v�k{��1)��=��$�n�\Ω�X.�4u:�F�� ܵ�m`��U\é� zx�qc��k��A�u��Y*s��f�x�s��Nnҩ��/���qD�X�2�:ω�ZX]��n�3��=D�ܧ��uP��q����_�iWU �Ȫ|��(@f����E��fwաEg��#:d bF��t�4h��|6�I�CY�(��c��WF+m��ԡz�d-G��%Y����Fƕjj�u^�~��_�Ԇ6P6���U4���Q���nҘ��ow����]b��������;��/�;=�^^�MN�٭��W��T7�1&,��@���4�g^-bjH-�&<������J���z�]n4o�׫hH���@苶�F�	H�XBK�ݿ�:�x@�j�yݩ������h`=�����x���n�T�/�?��u1%�ʪ���Q�	��b'��f�UŜR�<X����� ��O�+I�"��RDη��_�EN"�)~T�.)�`U��L�5�y�&}�Ϊ���Os�Z����Ơ�y��%���u�uHy/}��Lǖ\5T�\��5�ʞ�D@ jDr5S.c���f���~�u*����3�ǛBn��q�<�\f��([M�D���7�|_[pI�霤�L�	��c��O�0{���s�f��o6���Î'6V<u��{ơ�;���
͚��M�0�a�dG�����:L��u��JM��\�)��{��������9𮐊��9�v@��D�ɱ�&�ٝ����m���fX�:,)	�]ޯ/e	!ꙡ�k����DR�J�q�Gu'#A�����S��ᗑZ�ob���6�i����]ޭ�+;7.t�`2)�繼%�ՙ���c7�1�S�.�E�L�8K���硑�K���\Q�i$��W�}w�fa~3���ټ\UҪx
2ks���Lj�^����JZ�����@D��2�����u8p!]�����!x-�Y�]&�u
`�蠼��S���{1��[�-r����ߦ��|�`��S,��U|�y[q_�!���^Y�+!�W�o�z�\�Ha��5��3�|��70�^U�Sy�ŌB�;�D��w�Pi�@�^�D��yd�HD���3pK���yθ��%o��Jd�`���s�9]����e^�q7	܆�D��R��gs���]A"3m'I�	Ҭ�p�����p��c�Eo��hp���1S���K����#�"���g�7���{�]�Wn!�Qo���<ۆ����jJ=jc��� �iH��>�M1�xS�{2w��C�ƕ�Lz��}wS������d��[�n��>�_wO�ț�fK��^�ʎ9��C3Y���it���^�L��*�=�[�K��yg�)��-��{Z��o�����w���~����<�޷1w���B�s	{AP.K�p3a�"J
9_eE�+/�7T�s82κ�:�f�	��nw��W�!F�B�洃���n��ՃյV�����m��l ��l �M��I+S��M@�`P\�(/37�
0xUR��\ ���3������0)�7{���HrRhkϭ��D�*,��.����V�E��W��̅���ѵ-j��]�񚅦Lٙ�M�[�Z��IB�+[^R�F(A�x�A~F04.�NW���֌-�*#�lSfs��ޘ}�ǉPH�n������aa�.�Q��y�YZTt	m4�Y�/� ��c��Q��D�C�&�h�dۺ�쪮q]�R'"7,����'�8��A����j����P>��UY�K�����	n���_Q� �45/� ��,�kV�,A<;a�ZB�9��{�LK�,�G���W%m#7�nw���a�KN�"�K�&����C1��uMy-���p�k�/Z�JQm>G~N�dzx߷����̏*��
0���*�E^*�us0��^y»�X��jH��m)	�3<!�R���ڥyMc�9=��d��>ƕ��B�9��fga�z�e��cj	��l�)��O�� ԨQؕ��/��������j����ʝ�}2� �1������=��۽��kn'����j��;6C� ^�J�/�$:~bSܵa�����}t��+�	�}�N՝�{�Z�_,e!��/� +w�xݱ�r�������4���JB2�h�	�n�v'w�ߧ+�����9��ʴވ� �t�o9Ӕ�ս�Y�L��O7Wa�q�]��7+�ީ�s(J�Tv��϶�`�w��
LYKP��ge�'���gjS)z�EE|7k9������o .�:��<��r1�ݩ��₉6�/�gV.��I9$���:�l�YB�4O�n�3�����/�U[�Ph��jC2}�,����n��Old����U2�ׯ �d��1�qIe�n�m%_�rL���mr*��(� < �H�ώ������\×Za����rr����Je?\*���L�v.Jnؑ��x:.�]u���uRD
D.��#�X�r6E�V^�u�eV
�S�Q��R�����P�n��O����6�GH�$ ���]ʸ�;Bsd��f�%����P��J�DuK�[�\=<��.������t�_���4�����LL��ɨB�ؖ�T̬�wb�b/٤,�:T�\h�������p��� du\�]4�7�FEra�pn}W*A�m!�rC�Dqݱ^�⟛� 6�ܪ�o�J����c��ԓv��1@Ů��qPO�ɬ'�rM�����>��~����4l���Ϻz��1u�)Y�k�,nz���A�>IؒHC�"Q>�O�v�s���<�V���޾�q�e���9��!��?�R��P�]%|�׵T�~1Gcw�� �'0��uYv>�5/:'�y⸞�@CFh�,�}ʑz,�T��,�-�YR3G����[[��}��
���K��ֹ�]P�n1��AH�֨[�ű����K _o�Υ����/����[Me[L*v.�(jݽ�b��RHe7��8a9��7C#	Jk���N���x^T��l�e)օ6�Zj��,�Q���k��5�q�Y�Z4�� � �y��oeKS\F=;|��!�kR�\�nw
�:�ꆝ���;��hbm1�¦�s4Ռ��ںJn�V��P�3�V��u���LF�ւ7Wta�Su��Gq3:Ҫލok�J��ލ��[6���'���*��\wgCH���{����x]4VUq�(4���͙bkd3��1�'5��7I'䃖@ٞ�G���O<�b��[ڗ*Ɐ�WAQ�c�\�j\���f;��j��zƳrWe�ys��|�f�!��� ���<���S�]wV���٢�����low.���䴭�I%�T��_�0��2�N���̫F�w:IxPլ�����֟v�z�v�7[��x�0Z�f��<�юv�������h�!�V�ӵh��yB�_�L%%mլw�px��eVM�X��Z���VbKi��Ա�+�u��L1��-��DH�|�U֚�*��G*���]�jx
��t�]��q����bZ�1�{s{?rӽ6ZF]��fV!����F��Q��t.����=�m�ڶQ9�Yd�q^�YSzdY��v�.\�$������v�A:Ž͡���ڰy���1A�*ýƭ�I���]��j�i��#�%5��q��v^�2Euf��Й�uq������_^uA�g��5$�Ǉ>�����:ޯ�Pik�̷.��Q�����n����k�u����Ŧ�LV`��<�wU���`/�-gl���Df�\R^�]]�Yz(T= ��C6G���Y�n���I^<�Lǌ�w�����LD���PWV�	cFf���%u�I�2g�h�O_U��Ƴ�N��޹˜�49B�c��Q�7+mS&*��_|�m^�"x5[�8v�B[����kX%� �����}a�u]�Eswl���`�&�i��xڔ��`K,I��㩹Y�^['L��M�l��:�f�O��˙i��!��+7]�:ݻ��ΞLɒ"v5�K��j�H�eN(�\�ɇX����v�9ڲ����/s��}}J��9pn&�s�BhTuU���,�_Z��&ؚ�lٵ,�;x�	W���� ݱMp2��#�Q2l�a|j��3��.2�uSݏ��)�Zަ��y^�Vm��Z�y��-��!vMɷ��̰��z^�gV��c��s^����X�SV����a�-ċ,7E4��ـ	0�����DsEq �Ս��� >���
���׻]��;�
ݱz�(�
���Υ��ݖ%M���:�\�#-oL���y�Ndk)�@&�ڃF�$~��Σ+}�j�������+�ʨ�E'��|y�=�n;��f�1&ma��ȕ'9J\<���Ӊ,x��C��9U/3k6����)�$��Y����K���$�B�F�J�YV撰v{��]�ؤ:I��%E�ƀ��$*R�<+����o��]�9�ܺWt�0�V�e��N����h�;f�3M�'s�	�$�7-3�|FעOJ���^53���w���w�3 2�J��zn�t�f{�U� 2���C�l2 QW�f*c��Wa�y̐o����O����1`{��&�a�2�Rw
�Dkr@��>����v�1�����%v� KQ�"�n%��K���<C{N
�+�ؤ̤O�{�Ǳfs�n�9�s5�ڙ��P�F׸�qs�m$�P���bL�6)��s����*{�61�p�8Hݵ��o�{�`�Y'����-V�}.-�8[��!��]W^�F�Y�X_*��A5�8OA��"A ���_�����{��<��o�.H�H%��g�|��f0��y �w��������J��1)r�K']U��{�8�<Pլ�~�T��2��LكT�TI%t��룸�eVԡ����㇢P�ା-��hU�U���,cu�g�و�'p�/�a�Ӑ�}��a�֎8�2�8������ylÃ/�[�����ؤCo�vb�o7���_	zt�X�TT��CۖZy�P:�DL靂aC��I�ɝ �ݏ<��K*��u���<�-��G���VU9K�f���V�ԓ��c�D�ޙ����ME���Q�:N�#s%Qj����Ũ��9�33T�G5e-�!��
�>�W
��q{(G��E�S4J�;F�V��ʛo���Ϡ�Խu.�S�Y�x��I�(�O��Eݐp[����V��l����Pb�s��Ȓ��ܟ.�tC�r㊏��s%bS���� �(�Jbf����O L�����u�n�z���c
(/�
�	�����4T�F���*~Z��n	i�r�g����}n�i��!�Ԧ2�`A�-�߳ՃCݸC��{�a�/]My'�Mͷ�B�ՠ�|�����J�(�M�p� �ϟ_]��[�.�l��/���{��@�~;azp�)ty�|�d�:j!C%G��ec5��F1uoO_y,[�znE"�J �8�� \���}*�%W���f2�m��q��+l�;�T��/�����Ep����ʐtD������>J�5�}:T[f�C���~�q9�d�ߟY��qޙ�s��2�[N�Q߱s�^@��:�+:A�0�=�n���7/.��D�G�K�pK�F��y���V��{L�c�E[ɥ��s�>��Y}���U�s�Ғw<4�J����̕ð5}�-_�{Px��.�������(5bI�\�u<ʢ�L��+god��U�7;/#CY+L�k��z�	�DŸW�1e����CY�e�
A��&@ �m�     ��T���r�|۾g��f^�2J4���Զ���ePw=��z����m����Cm�ӞM4���I�"Tw�ǫ��ۻ�d����l�.���3K�^%#:V�K��u�i�=�P�eW%��հ���\�M��"�1�-Lx%�y�B֣��-��zb���'�_��t?g��|�z4�1����<��A�}*R��m�|��:!Luԅ�"�˗�P�[~�N+�*�ф��9N��}��G2̸�h�CG��X��]=C6xT7��T`��5)t�S�-ɤѿť�>�u�F
�<q�y」,,8���,�6�{��*b�W��0h�p�#�O�eM_b�Ĩ�n����=x���~D��J���"">FGZ��{eD��]?A��2Gz�k0���52�U�C5mi��W@�gdn8��5Nyu㶴[���P�4�x�Wgh�=u'h��1_�OY��o�������Xf��e�em�;Њ�}=�B����L������'�M�[��:t����H[Q�8����>_<�r�n��2HJ��Kʞ�;Lc�1S��DB4��~���J�R��Ӷ>gī��^ع{z�xݣ#�qTfO'���	���u�����pJ��me�L��~�p�%7�3�Z��9p#A��q�����}U%5�@���`bO��Iz��� $�[�φ2�7��Ɏd��<�R�'w�w5n����o�2��0M�|��FM�T�3^��}�i��x��ПSJs��H�K���5�d�x���ײj*�k��s�l�&��6!	�xI; ��~&�J�l�=����T�3�Z�U�Z���<�;�Dd��C�0J1�T�N"!A+'zC���h��+t�D�d�f�H[�n�{��8��fK�n���L3��5w)�>C�E4��J0���6���B�33�O�FT�+�oَJ�8���F8*-z�,2g�!���vo f��x�/z~�2)!��i�P��ɵ���D�ޗ9'��kA򯊍QO�D}����Y�{�l~� �nv_ݦ)�;�P\*:�GT	�rgb��c�/�V+s]��v���Rzt�ھ��ay�fmӯ��J��q�$����sd|�A����3W@c-�j;�1'���Va�ለ<knM?���������;���pX���Lj�	=�����S'	TC�f��-5$�C�1Y�S�x�ܓ�s�֊�!qyL�f���*�9���@ύu�����Fj�hs�)�ݨ�WU�m���'q�)�2!�����c<��hHr��>�5s��Au�y��F�NBB�k��}�?1��2ߘD�:M�r�U�IX�ORx�y��a�.xm[�I�i��\��3g�9�۹�.��fo:�1���4�1��k��\�vc�b�:�/6g��v�)3��{u��ԓىu\8�֦��xҠ��]G�����x����ML�Ա�@`q�x�<�������)���j�1%�n@�:u����w���M�ڨB�Y�{O-��������fiq�1)+��'kB�o|g��ap�E`rqL�hN�ٗ��>���n��Тa�/�0چB�lx�>��(z������gWYf�3�b|��4��������S��K�N�ܾ	}��N��B�y��c#��KVO��s����;�,%�zU�k�d��$�<%;�VbE���c�/��^ԟ��6`��^y��$o�F-v*��=;zOXT:��1�L���$������N�%����?u�����q�����z�/�����K�DS�B��4('I.]|�F��8�">�ٙ�t���>"Z��6�L�G�(���&]m�f�Y������+�3精�����IEv��k��Q�=�2P䫦�U�^�_Mb99�a�p�lm�5H��`�͌~�� ��_[F���W#��:<ۃ���=��-�.�.��@���E�lx���^�F��Zک�¦'���f=EX�����w���: �w�>��5y�2*�7og��v����]��bR�חĪ�iv���=r���~Ie�v�H���OP=��KV�l�0g�\�,�m�[Gk���huª�]!p�j��U&j�v�H;v�J�䚡���yt����l�#'15 �QK^<�z�Ǡ��л�s���N�c��Jo�����@�������77�8'}�l1f>���dȤ/g��fct�#A�8��u�JT�k�s�P�գ5��0Q'r��n#S.���j%��I$�p��9C�S��������A=
%>���C�L8�ԍjz�RY�TrߔΙ��_�@�w�K<vC��y+��t�#�f�s�ۃ��:4����Z\�	�0�-vn�����(���iˢ�qO�
n�*�%1M=�M��OWϔ�4�:g/�׈UL�_N��b=��RW��3��o,�c�'��f,��]+�.
��<�yU��\��{�\|��sj1�J�4#�Q9A)�S{u��G�s�b���(L�Q��`��bGx��H�ꔖ�|���Q�u�04�E��J�P^h@a��%��y�p���i�@De�U.��k�@�EN�����u�#�8�ވ����P�Mv����>Ψ����t�Z6�b�['/u�x�MarOP�����E�>�5��-	Q�i^�f0왛�R�H���CzmggL�䣅#X|V[�F��q�{X��w��U:�z4�u��P�/�K=���CL��s���L�S�_�e!M�w�=nPAV.�B�Ic�b��D�T��;JY"9���9̨����ȕ�� ��  cC` 	   /����T^z�,���i<�*Fҳ�縰*��Ƣ�H!�iAm�υI���&mi��0�h���^1Gx�Q�Dmmo;�ջ���GTk�T��ߚU����G28��*���UOf+P��]eLs�oe>��$�7s3p�G���si#r�U#�cU47�h�+Zb��F~�˸ύ�۞�Rڌ��1W���|�o%{ʹ�/V�
�~3Tw+87�s(�q������O��'�[�A�jYæ��w"Y|%C���/��'�S:���h����sfĻ���e��Fw��=
�=er>�ez��z������55�yz������Ϗt��-*�cU���av��}]�d�3:�Ab�:���O�����#w<��{Na��W�Rޣ�n��Y�z�PW�	C�<���R
�53Ք�MB���c=�s�qF<*�\I��P��^��ve���h�;-:��
�W�
�춰�� m���8w_#����|��l*�/#�.�
T�>7^?E����yj��AV9���;�^K,S���ƥE���V'���7�R�j���_��X�RL/�WƋⲡ��[Q=�i�GR����K^m�
�E�.���棺���������xt/!|��,UwؕcB�9(��1	��i}�YE��&�m�'zy�+4�gL��و�z��܅X��7,�y]%б��oep��S��j�y�J�"��+r�1�:���t�d7�b�޷Ȍ�g�}H����G�z�`Ih��]遫�� ��]���jT��{����1��t/D|�a龕�������(.��X�^>�6F$ǟy��,�y!�;잢���dh��2y@���lE�~`M�\ǖ��Rz��8���x��[OU�����]��i�B#d��ǉ]b����<��c�dt*Go��w)[OLdۃ�&�<ȃL�Y���˨g�6%G=�E���'�dFZ~��"���BGumc���Uh11��R�m���r�,v��
�Hk� %LLJC�{�"}/i�ydQ=�<FȶT�@�gȞ�g��G�@�zP�`��;�:Z��ag�ƭ�b=����A��7k���	3�ѱ�]�ٷ��Qz�=]z:`U�l�X=Օ�޹�rO�K�b(fGg-�1�[�/L�L�e���(
cut�'����w|��=,*6p��'����"�����:�޴UB4L2#`�&��j�Oí{����.�wm�^�i�]�R�_�]v��@��aٙ�"�ܱ�-]ok��ٹ&A;GS`鴲s�r4����Z��1���1�j�r�A�YHܾ�D<����6w�C�E
mA۷/he�-F�@;:[���J�Ʀu,���݊䯪��?�r��FS�4�̌X<}�(��G��]�Qc"�`V�d������R:��Ё�2K`ejm����*z��:7�6'kVz��"�f���N_�-�Y�3�x���M1�׷�E���U�e��̑���ѸU�3�BN6b�e�D_�ӻ��MZ���N�Mga���CF%g+�Vx��|��c�Y�������d��(����:8����pL٘���� ݛz��/*��#�CF�՟���h�p�?��J�+nt|r�J-N�y�w�ws$�%z�^�c�O>U�`�V��B 
`Ӌ	��Zwll8����U\�/�W�F>�*���/����S-L��L�X�?]�'S�jQ��T���n�B��҇|�RpT���%Ŋ�����Z1�N����T�{�sģ!����&?gg�~as*Iv������7=&��s��j��9�iSɖ0�ޝ�T$���Zp^Ekx�\I�Ĉc���f���c>P�V<
��n�%��ly�΄�v��Y�9��Sʊ�O�\(	�*l_:�2�*+ ��r��n�9&��,8k+��m<-^+�Ȋ����.��{����4`�zH�+��s���psGz㭬�����h���7���7���L�����2�lcb5�_v\�%�B�jkt..wu&�
ӂv��n�(���[%�tM(ʾQa�'�F�5�W�k홋R�3�����3e�s*#�م��ć�5�Z��N��X�!��U�x�-gϏ��l��i�e���T:7,���X�yQ�u�w<�:m� (��N����m�c�֗K�hN���n&r7)��z}n����Wy���o��K�tcbH�q�1�U���sJ�WU��KAqM�϶히�E�8��{�bQR[�����`���������c%q2���DG�ܦ�L�z�8��=��\d$ft��"
�-�^}V F䉨R�zǦ�ꞑ�����Ҏ�7��2���}l7��.�H�����eʂ���.H��=6���E{�_���	���1���tWWҪD��2DQg9��e�n�w���mQ�����.}�8o�p�vL��|0X/:�>ŭ���wW�볒+ǈ�8zѳ�(�oM͎�e�vk��}�K��,�<�,˔���[�Y�z$��cbϱh���v�P��1��Nw��͕��:"��3rA�	E��?}"�KM��ғ/�|s�
aɼ�]��D
O-���݃�ۊ��\�k&s����X�%N*�����m;3*�V�SY����ڍe�[ظ�U�*dװ�w���#L�eܥ�t�MXy}UX��QI<�v����j��na�	�u"sj�ZR��r�o��)��0�
<i�D[,����T��x�C�-�L��d졂u�i٫��컣�8�]sҚ�}LWJY���v0�a��zy	q�ȭ���u�;c���Π'��05/���v�=wUԹ	O�#�gQEe��S��p�j�;%��u����Y9��~���ygc�p���檒��iܑ9Z�kD��1�7̜k�VQ:�Jzk��ٮ���K4���& fK����U�Hrk����Ξ�s=�i�,�}�v��b	Zʊ�p!!��o��J��ii�+�99�vX*�������'�J��n��M�m)'r�W3���E^��P�����-LA�8:��v�� .R�����8#��zݫx��~W�;���I�x�1�����Y��l�B��NWz�t�j�g���9�� ��tE'ZoMV<`�����1.F䖳�tn����|v!uj���qhc�,���DU�a�j�N=o.4Z���}������©��h9n���don�ځ1*�¶�,��)��i�v̒K��AH�z�t9�R���[8q�X|Ӑ��MP�+Dgоg2�aAe� \��:���r��S|�1R�^��W�V�u�?�"j^bդ �N��	�����j��u���Z��8[�k�\���6��G�Z��J'�m͍� �B�Y�a.f;D��Y��Y>��9�]�פvW{�=�b�~��i�s�r��.%z�%m@�9 Wu�2_,�B�foP�*1,lڃ8�������nk���Q�L72�&m�|�[Uu�Nu�C߻��e�Υ�L���㙰�q��������<6Ս��"�M5*�R�jVՖ�����>�Yg;ծ�K�q8�h���W�u7��|.�>y���kM;5�yw-����\�,Eoq��sf�WTX^��b��ZM �!�m� 6��m�   8�I� ��ƦT)�R@ @    � 6� 4� I��`   6��`                  m��     m�m�+�o�v�"uԂ물���ZO=�[7i�ѥl�fɹ�p�n�)��+o���1t���]��q�b�jl�����g�o����97g�s���֖�Ղ�n�W���	��0l&ZBP��L�%�:g;JX6��_^j����Ĝ�g��y��،��Ҝu�x6��   �����J�,,]��Q
Fm�������]Bo�j��ַq
��Y��D�enw�g"�P��R��.�jp���}7��gqؘ��R�,�t�̕�,e�v�$r��<�	��:��E��T]\�hg�| ��ӾoI��Ѓ���q�/���u�Xڵ2�t���`�3��[���Im6[L�M��    �46uU~�����P5�N+#�n�4MaA^�S��eX�k�F�KZ�, mβ�$��𝁔����te�7P�8cmY�k�a�p��lFn�H-M7Y+�SM�x/*����{kf�ݪ�Ѕ�m܊�[ӣ�7#2�t��$�.>�_�mx�pi�g�s�n�g�yUb^1�>��Ց��]��X�7������&��G(yW_���;��=�(\�>�~w~J�"[��)b�n8���>�5t)@֔�]��ؼQm�d�w<eM����lfT
�ѝapb=
�'�9k7*��3��{�ԑ�	�GݙුSaR����㐲�yQ"˘#�WZ�6Y�Ǿ���,�)yǯ\�5�EF��9�q�Ii�Y���F} \�������D��(����^�~�{EuW�hH�����:5Iz��H�2��o�y�
�:&��eU�=8�ZHNζ(Z��5΅�`����֨����`��2cXA���ʥ$vu\��������/1���X��.ޞ��{2�Ƿ�+ii��~u�����I���R�꣧���UT�� �"ar��މ�b����%fCOkI��=�*���`Û�gwvA�6҄m�rK�Ƃ�ڭ�8e<��.U�ﯲV��P�|��,��u�ܗ����:ek;�+M�Zs�=�l����n��z����@to[�qW��׻V���	�c����k�]ݾ��^�#(��Dz]�Ӻ�\�6BŰ�cQo�3\(K��$6��|��g��5:�*�����%�*�u˨8�T�j<��$@�R��&��;����ݩ{����/EoѼ�?t����8�Ү���EJ:��Kۤdj�c��h�7��2�������KҶ��δ�ޑ�D�x���(<s�ޘ���$�:��sU�u�&��b[H�G��7тw�VR���)�`B����U_�.�?n�25"25s�2���{va���{;rc2ϲO���MWBISm�6��vw���/��yj%B��կ����NB>�k~��nF�4�=rt:1�s��-֪���"��i�
̔&�P������@蹓���r6�v���G��92.���(J�j��ep߄>��&*����Y����8�"�����XC���I��}�g�&pʭ�;��pT��)p.������V�����	�#�o�2֔����'ʛ�^8���r!�}L���hG�k7���A�b�VM'��_��Y�IUE)�r˸��������;(��܏�mȣ�6���WN�5���}��l�w��s$�u�M��%F�N<��v��ʼ��<��Q�Z��>7k�탻�f�#kg��I� EE�y�̹$��M�CH�p{�Z�^Te�(�pK�u7;;���������TL�a��+�Ns>�� �Q�7�|)_��b)�9��ؿ��P98[�!$�>�_n�<y�|����C��>���F#]T��N1��:�tGZ���K��VO���U��깂&8V�f�WL���̫�l �!�ax�gہ!ە8JJ�f�%(���,���>s5���h�]8C^'pՋ5��A#;�7�.�������9���0ȀY��+�"��!�>Q�z�mgl�d�*~����Z������'�a�qMqR�Ui�b^G*}��d1������cL�\28b��ّvA���]��t�^�o��Ð�2�շ�xu_{A䶍����ڽ#1go4�D�O����֭O*���4�|X�8&�(;�Ƹ]����F��9�=ST-��Rϣ��Wmk� �_N����Ř�$�ǆEA��)-�ƀۅ�3H�E4�D���5���s������>9�1k}y8
��D/3�NI�=���6���/m���j��t�f%��E�7w9r�����Ɋ�0�p�\9��v��Ij�K���a3'�JU�c��&��op��BùS��g�y3������O��r]q��'��B�&V͝�ޥ�7���%���×�:k���f��#,z}v��:/#����;� 5�bN&|L_M�&K��b輛�vJۺ!�"A@� c�s��@���G�����MC[�o�%,gM��37�'I�]�}��:V��):�K�l�jU����C�����Qq��ח�Sѭ�GYH��W�,I��lz��ؒ�Eӕ\���sB�pA鬾��o���&����O2�0��D{�)D���h�I���C6G�+��]1�dn�>��\V�=I(M�N�`àU��PU�qЇ���a�
�0U�H�υ���V�˥�ڀG����H�e�xM��"N���+S��VÓ��5��t3���%4 o3�v�����;UAn�ڼ�1��oQ�Wj���my�
 ��=uX��)N������q��k��o���Mٯp_n�d�ө�ev�{�Rc1]I��o�	L\�<1�ҳ�޳9U�8�7ϴ���j7(��ӆ�ڍoPג�9��Q5S�}0`0�0�(��%�m�I�h��e��5�W��`a���ws��2v��VN]be����:�]�0;x���*��UW}ú��.���6��c�(��ޮ���rtN��w� ��$4�26�      	�xUЩ4�;dL��_Wb���ر w�ed��[]�r�'�aCC�a����TL-�s�$9���W(�9�6�%�W��C�dT�
FYّ���.�{�0�7;S�JV[7W�k�Kt�W��z�ұ{F\l-��_~&[�ͭ�m�E�џ.O�E��U'��(�������L�3L��(���z�M�g����𥪢r���Ie{t+��K͢�6	�7�)��ܹ�?h6�l��,�۬���$.��oE����M��o��V];�8�ֻ�p�fԌ{�~�+�p��8�J�u�l��Fx57ˇ�'�k<&�r'�\)�>�	�r���(��T���3����7��\)�K��	�P�U���?�eg�DYhX�;~]w&�6�-���l���l}A\������Ge����^Hk 漢�Т��um]��ҧ�K�d>y��������Щ� 7N��5����^�mȫ.f;4)�D/R�u[�۲��&���W%'3ڱ��f���}p�C�\ǫ�gY��(���u�����#wb���ҧITY�g�:p�Z7�Ǫj,�4��R'�V��r��[&!("q�YeQ=8�/���T�M��st�`�#�
��M��H.G3t�'#�6���ݏ��|:��3��t�|�7pݢ�uO�sgm�K�s��9�hά3�HM��m�۽��#Îv�;�b�D!;<�&k�u�	�XF��~��U�r=����w>�´lT?���=��7f`��y_��a��Ղ�C�aΛΟT�x�\��zoB{>�b�2����i�̅c���(.��ǣ����nO\4�<g��%�Ц�-֯T�o�	���C3���a�W�n�Bj��z^�`]xkɱ�G`��XYSp}�O7tߪ~��K7�$���ڎ5��+�;�����
�����{8����MR$�ʶ�nr�F�"�Ι�-q},}cD�2� �q�ʾ�vթ쟈)(I� �����Aoi�\$i��s��k~;1&��ϯ��\η&�%qHP7V	���Ṉ��b���&�h4OUWK�P��g��X�Oz�A���y��}�찌����$ h��g����p����R��^�oٛ��}�'�B��R:�Ǘc
!��DO��e�n��
FݐTC���2}cA%-C~섺"�.&�`����G��f1�Pضl�O�k��`�n�Q���Up�3b��]`�N�J���/S�����;�O5&��w�y,�K�`x�;�Y�\�wr�D�Pޛg6%e�}����w���l��͜4���%��[y�o��"�'��n�|�Nl��=�J�ޮH�ؼA�l��rC�����>��z��y� ��[�����I�9�5[۰�eI�(��r�ɂ����{�mh�v��c�9j��c�.��1��Uk�����a�������W��>�c'��s��z�j
�
8�tz����q����b'gK���`�M5�K	���}��Ƕ#�/`�vO��Z�OF]G��fFT.��0����Z| -j$P��Ԏ� �3��G�]N������ޢ=f��S��\o�3��ypD���}Ni��P�x�D�q��}KT��%�@Zѓ�Bu-�nz��,L���B�)N��;K�mz�^(��cj���o\#�Q���o��3�~�n0ܘG�|��f��<���p;s�����+���[꠺}�����t�zi��i|W	;s�ݛ���f�A��>��}d���0�o'�A�*�߭[ͻU�����W�H��2kcj
K��(�ͳ�f��(�g�&�������Ӳ�#F����}��1ײ���C��,��x��|\NmeN�y~Z�Q�v\*�wv6�N57�	�TEF��B��EwA�p�2��|N�v��]��zR���F�GK7k&�����R�\;���G;%[u���u�ק�/���̈�:�s��q�	��+eUx�S��YTgp͊�¤4��6~�<�f_��٨_խ�3�j�j%�Wk���f;��=��<��8�1c9�]Gbo~�7�]4�q�ޕ�YK�U�SB��A�{lטȪ�W/�Ǚ]������@  )R�~qU4ƁP�C��+�c�-�|�]*�y؀�[�5�;��r첦�j{�ڵː��>��C����iYC��9�\�p�i�T͜�W��t-����u���2�(�[�<]��m[Vb��'�K��!W~6U!g������]�*�éǮ6Y�ڌ`C�g혛ވ�r���9���^�;������UҁR��9�y\����dP��`ԉI���g�F.@����}��~ߐU)���$�r:�O�]]��ׅ+�m�lf��ռ/s�Ǟ顨��׌A�ta�Y�ݲ��ꐐ�{�V����lh�k��h�bs�W;5��n�z�<.dN]+�u��P.��ïn�e?y�]�w��*ob�*���������ܮ���fӘ~��7jx
*<�n��g��z_���U＜w��ˮ��ٵ�k��5�#骛q���8��×^�\��6�����
9�����֬�4�ə�˗+%^B>�-��]��w=�.�Q]K��z-(M���M#c!���3��	%��s, ll      *{��]����{JlSUTvn�������ȉ��D��.�}N��$���$�i������軧������3��#T���L''�/}��wqɠwa��C��0�q�[����=�L���}��c������/��ݫ�7�l�셆�=9�o�B���~��綢u
=ʌQ� �y�D�5�MwtÏ
��W�{����:�R��;J=���Q��F��؟�tyᘸ&���R8�yF�C�i�F �%w�2�J*խ��C�����tS�N#G���Ż�}0��z�u�f��C�c���.c�` �v]���>l�n8,�"�Q�T�}nt���ƼF����~����[0[x�yV�kA���S�������eל�z5��Jx���rE�-Uz�S��D�P����<�\�*;j��X��%�1���mͯY�z������eq��]����/U%��k�t��I��.fUZ��!B"$m����<Q�pD�9q��
�BF�®s�!�r�{�NLRݔ.T1/$t%3��㱴\m�|m^9&ʀv�����ú����Ϻ����b�?��}jp��I
��)����t��v\)���\�s`(P�/Evnj�:���/t��j\����ifW
��lt�n�1��e�+1��w6/;x�	샰wf�_r���2�a��'?��`�bv�1E��V�'q������ly��ȏ����e��ȫD;,`�Y�����S�Y���ٺ]d�z=�q]-4��=6E۽���"���ng�z|�h#�2��c�&.&�����܎��T�
�^�lid����ݒ��K]���#3Jƪ�n}ހ(�>�$�)�3B{�Y�$���V�ei��at��J�iпtx�S�_��]��|��UAl������J�z_���\qX�𹜻�4�Vֻ��qZft����hLo��/�f��:�WB�����F��ooԛ��A�D��HY~q��|��f+6��\�/2��cp)�_/���1�.zk�w5  �w*�^(�R�r�'Ӟ9�mp�w�5��C��qz�N�'\7��,��ţ���+X/���;2�
�9<������*�C���x���چ[��Ex+�c:�������ǯ_�MK�Qt<�4���_�vV�P\T#�;dYX/E?T������Hg�7Ȝ�xbcaü"uHw���A-�jfM��]�v��bX(90�a�%���el��"��V���b�\	��Ib�:�M�V��YT�4؟�e���C"��D�%��s+�Fp#��0��X<q��rN�z��K�E�sl�.{�r��3:�٠��bل⷗wP�n�s�5Ya����<��	���{���+n�B�/�S��]ک�AiVE��
�[�o��,w�W[(=q_Ls꩚z:����A��"��T4Uvo��U��7��5�T<�0��py��gQ{W�r��
���#/��i��᪨�aV:���|s+E�)EFoM�۸Wf��d&��k������	 :�y 
�vI=�g_��� �v��T�Ƥ7����z��]��<�C�	>v�u�p u�@ۿ���� e�a$���Ӷ�g���^�CL��j��|0����I�S�j��x�E���䓃�9�f2���1>a	�{Ɲ�$<��޲@��� �y���m�����> ]/��s�m")��F%�	 O�q�V|��[���_�<����/����D.B�&�;��B���L�U˩?���H�<¶�FȄ��K_��I����Ց�lk��U�д5;_!��ҩ��Kj�+X��w��
$�Z�c ��í����S�AfW����ƻH���KNݤ|�3�!�
'�wt��gL��L�R�{��HS]�.����٨C�HC5�欓�a��,!c�{��\�k�' E�Kl:�> ��@�`y�'RH��6�s�u�t{���s;��߇Y�X@����3�Z�}�d�3I﹅���^S��{1��iSO��k���$ێ K�_�#�*}��k�Ǯ�8I��@F�]|����@�x�Ԇ:c'~̞��ڝf�Hm�fq�Oе�7s�H�`���t�XM�������|��xO��^���pG9��Xx�Z����� 8��۽~w�W�Y����[ :�H�0!��1��B��_}ܟ=Bg���,����[3"wyvL���/s&��b�.�C9c�gk�w}��vl�{��V�|A�1�:�?-�M���;�	�������r�"��t%mZ��|��<��dq�ks�84��y/]e��� Gq��9��:��A�eD���F�V�S�ѥX*VWnj��uq��u��7��y=X������-J�ʡ�0c�AV��:��J)[7��e�w�Z/��Gs���݆�A�P*pE�r=������w�2b�O�n8����Ƀru�Z[�*�(��&�\�nE�j����ŝO�ѰF�Xh)�H[�4��2uJhG@��&HuE��w��ٕ�&8�)���9u�X�v#ؑ��8��G��M��ٸk{��4Ѡt�ؓ"�d�����-��[�ˆ.�v=�hn��]�+^IXKQ�ǂ�ٚ{EA�5@�����f���b��a�I�Ό�����A�M�7��L�Ɲ���WNC\u���Jк+�s1is���	(d�}ӦU���.�Ρ��u�K7ţ�Q�
9�N�e�7��5<p�u��Y��mQ��n�!�.`|�@���3jRu�@8ݺ�:N�|������DR��@�˩P%��R�I#ۗ������2#7NΊ;���4�
ʨϬa����E�`^t�:�[�0�b��}G���L�G��6�ӎk��&��h��4Kk��W�~7~I�N����6Wx��Fބ(I���x��ѻ~1xgFo�F��J꩏iT��O_��:yB����ڧ�[� �E��3/��"��c7(a������~#n1�.E�kE!鈃��z�<��C�ꋏ=�!}R�Ps�8�L��{��(�Jxʅ�:�.���A�Zg�:�(x��#+Q�+�v��Sg���Ox���t�n���csP�E;�,o���/c����º��ª�s���3c���S�|��@y��"5��E��j���'�z�j}?M�=�t��F�<���>SC}����S�{4�~�jo|e��P�q���tng�%Gy�Z{:��_Yc�|�F�T8|F����Wf+3}է>�u��囌=����Í¡ŕ�����m#K���W�b���s�����i��S����Z~=�����l��-}W-�N���eF[\W�
(�$ѱ�8܎���xdg��;��'�C/�76r錓&u(����25ƺ֧s�JA�����n~�����"�ϴ��#GG[��m��Mi�-lZM���w�I
ڸUn�%?�{5�RC�)�dWkd\�[��E�56n��Wj�;�}��ٗE��1F��s��s���&ӧ2�������ls�z���Lǂ ߃�=M̡��v�h��BtB�|�N�8�YW\!�L	7�YTR�Z�9��=��.��$��F�(�w[pȇzo����tue/��G��$k^�0)�m��ץ�:�z�� �ps���q/����K�۾��ָ�9�{z.�)�x؀�L�|�n[����g�V4�����z񫗥lW��K"��C�]����lB��8*N"�\u��:'M�v�]���{Ok)�fE�f;�=1��;��X�s�u��&�5��3���\��46C�DY�c�����QQ��B���V�=��i�}�[��ý ��}����b��ܯ@��N4G��S[���T�vn4��a�b�k�/�Ϫ8Y�S���YP���P��Q���{:�X���o��|��{�vNUn6@� ����^�U�(qx�/�!��K�Q�λ#̘_+����o6#Nv������e�'=y��
jj��������8�5u��~��zZ!��z`�sb�/C�3���y�]��N�?dc|s�o�g�2�M]��jB�F�$:&��"�<'\�#ҷe��o�M\���T�A�}��w7vn�\Om�{�Vs��n�1��t�tC�Ξ�"͈ͬ`�"Z�n��^����s��8�I&�5�+:2;���9��� 6��� ������ ˢ��OuO;�k��6�l���F��#7��j�-�F��^ff!ð ��i�嘵��
m���E��NC��S�q2)#�`Es�˲<�ܶ(�^A�v��ӸlW����ׇ��!���JȢ��Э����)����Y�P�u�m@��4:����U����x���|��'�F1G��Ѽ�D�4��0����%�@�����U��X�4*ڷ�ӇL�l�bw[Qe�W%�/��tv�&��b�֦���哖�_>L�ǲb�=�H�o����"x���}�&�>~������UUa���.��m�=Ϊc <�f�O�q,��>�O�^ Á���o8��:60�}�������z���&��;��}*��M�=������vpD1�A���ӎ�G�޼01᫔�8��:~�=�=~�Q�\�vì�&|�֐�'6c��m�4c�˟$��m�kn���z�닷�x�ÿ��tF������U�Kk��e�_m���6���R�����y>���<z�e`�v���^�)������5l�y�����{,wm"�Q�7���c���ڬH�g����!}z��W]p�[qt��H��j�o�"ݹ*�i3e�]�E滍�bu�P�<�b�:3\sǜ&�ɷ+�]2wу�����:��y�ҕֶ~9�Z{�᝽�\y�������i�R�N�:�r��#P�7߰d�t��OmjL�5��1���m��[�_F~��wU���}�7J�~��ϴ*a�)�&Tzbmn����{	��%q��el�48{'�E�f5p���C}�e��|��Lt�`T=cC;����;5w]}3=B��+$�U�~��Q�dq�=�#�+��hENpܜ�)������u���}㞝�4����8��S q���Gj�DUy#�c�K#�Fx�3�avyn�X��L����ӓs��!�����p?ܶ�j�-(�V��^����Q��+��� K��i� ��Ԩ�p��u�rW�X�^��1��-v�?��>�i�T·�O�wqu9W��_����ޜ�U����C�=��ܑ�O����������x#�=���N��pL�\��Hf�,�K�m;�~9a�M�\l0��~f9�W6�;�U{�X<����`��7�t$"�u_z�/G1��r:��R��㗢'M+��8�w��_����!jU9��-6�a|n�r~|E�e�7o"��Է��x�a0.����r�$��:���v�;S&���la�J� �C��G��)�<w4o^�yTt̾9���<�Bd2��8�vo)Y��:�b�1���
cͩ�|8��8p��3�Bɡ/��Xv��l؍��a��ޢ+(ȼ��;�c�c��u������^:/���^w��,������ihc���upx�D��2˷������t3��K��r�a_�>˸g�`���e|.�˅�jc'OػO���I�z:�h�jA=>Խ�h�.6_�+m��^R�����F_i��^�*�K��Q �e��8f��!�G�HǙo�/F��{�W�.;|ݑ����j�;>Yv����gT7<�tx"��h�(ՊE�
;�K3ꊢ�s~��fF�{�$N�/�*�M��E�B�F|L��;m
Qz�<�J�e��o�Ȭ{Lc� �sY���X�p܍Ns��)�@PH?k�j�łU�PsT0ANP�:��GZ �K�5��4�0.KOeu~�)�\�O�E��y��dQ\����zt��/G��ȇXV��|���`�\$��ǣ'3�H�ޚu��|�(O**�YQ[>���v`�s����+��R67F���w��I�N[�Ȳ��<��J����{|��J8��Y峩ѵ7a��p�W�&�T�ͭ	��YjF4���5׷���-�Ւ��K��ܗ����q��u��+��}���(1K�D�J;�][�V�y}�m�L��Y��;��/{ӂ�/���z8zZy��F����3:���dN��cV%U<<׎�FWu:&}t:�Bgz^MYf����c9=��}�.��k��]y�L�%���d��<E�L|Ɓ�����U�	\���yZ������/�ۙD��W;n���A���dLO+�}��n��_�+�f�0D�Ryp��X���]�F����@����or��ؚ�_\emnwT-���`{=�c*𻽷���!��h�1�A lxt����O>���{޳L9[*߭o�J�V~#��}�������[��z�� MI4'S�7��'�r|�h��Ĕ<yu_���x�ON�;���g9��*�bR���O������x�u�D_�:���I�)���7�&督�a�b�������s�z�?i/�x�i�짾�:�ڱ��1Q��w'���"||j��Z/\Vu����O���A�=!Ur·�O��7K͞�
�����<��ϯ�Ѕ�W�{lNP����a~UM���s��V�=��>B.�i�E�2�v34V0�����3q���O)�k�:sRMG����!)H.�t�0����1��[�[6r�a��:��9�Y\����������nl:���NI � ��m��   l ,KPF��n��'y����\�}�h���;��p=[δ5�Q}+���EP30�a�s�Ę��<�mO�ԂN\�o2�wN�%�^�T�{�]L4��t/ˮS6gr���</�ᑈD1n�Bc]�$d;�=ѻ���_����hF��ɑ	��]��8��U�����l�Q�juE��R�YaT���&�P)�7YW7��M�0�DF��3���۞��5��MwM���b�F��\dJ��u��1�Ǡ�7�F���k�9�u���o7F�8�c7��}.z�`�K�u1CX�LV�'[`ȏ�U�������-�n<�ڞ�r!���~����{��6�felXg.���V�x��u�Ϧ��&����l���WN���>�Ϥ���{���f�
X�c0�ި̊��JKp8�8R���'R�Tq�x@���갠��*m_;Z�u� ��m�2�6���-��뜘�ࡕ��I.{z�o�J�]�;$;1n�X���;���Й���0���V>����C�=�<��z��L�V_�d;��o�v��P�2�����[��F�uݹ�������}I�2�cڽ��u{8�L�]ٝ�t:DCK��Fj�P��v����|��cj���3xv`����N���z��Y+]ˆ���Z��=�G'K��T���y��^��נ�eW�ْ ����K����r�+4D嗐�g��QT��is��J1��*�M�ݵ"�J�y��`M����	�EPL+���=k' ܬZ\�zd��쵾����1T���sF��P%�f,�D��켇�G�dlLxM�J���x��'�SP�Y�M��M����?w�x���!���y�����?���"bw���v�C��O�v�<��p���Fζ!���:��f�S�z(���j�i�<]a����8��H銰{��M���\:��hs��NG���E?��1~F�h^^ڍD�����n6螌8�nh<_��]��w!(Z������ȓ�`������wd��ǎC��2	�-�V�ZP;ڠ�����V�t3�\!^����=/������(���w(�hP=���vǤ��=���uDT�K�=i�s��Ɇ�mh��s(v�0œU�/��^���ٯS�ߌ�75�vt+	���ܤi��H�Ǧ�XC�5�������JV�HMѬ.ħa3�4�n��m� U����׷��AND"ɼm�t���#]���.]fW	�&�W����V:�Sj�y��l^���>�7��N��n���]`�,wS���qsyi��=�����~�W����u>an�у��lyza���|\�yy�+�Ja#����2�U�
����w]�ay�C�:�;t���qa�gUwE֬��H�����|�'����R0��1��b�M1����U����P��\���բ�_!2%����j�Oo�A��
+�z��ݮ��bl��;1G=�Gi�%��H�`"9�)�'�P���m��˺�\tMT^�yV�5,Җ�d4���#G���dL�ꎺ������`�Z��_�c��-[��5�h(=�����9X��W�MNF�S__0��7<r��OJϞm(8�{P�L�f>��1�"�PGV��>?o��h�6�]	n���eyI����R|c�l��>��^Q<� �s!�YsBvؗz����QSj,�'kԢ��*�C�^G+��>�+7Q�Gng.j�],I��Yn��Q2Gu�mt�,��	�jU�p�8����9^j�ܢ�=�o9��ȣ��H��T�^[Z�D�1��'�A�9}O���P5�f7���Z*���%��To�$����*;w:�54�r�ʾ��v�����]��a��aT�Z��j�p,��u(Z��b�VJ�3/���������fS���d�5-���u�ά۾�\��S%�ԧ*t�5;�P���м%�k��1�_���k���䲛r�����Of�׆�b�c
+����yBN4D�+j�Kˬ�8�ڑVy-�2�U�dR��u�����Vb���q�q��.���=��Ҧ�r�  W>�D>5pj����UTd4#���]���5�M)�@��R:����w�}�����;�g�~Ұ�w`�"7��˚�u��Սu����M�=�h�]~�~�0B�5�T?{���p���e
�R�̵v0���<�x���/I�p��0;�}�YCi�*�}�0dGCA^ᵅ���	P~B��6���ͩ�v�z�+���P#v9�[AF�l>���}���Y�ã����*Z�j>�#�>��Լ9sEӜx"�;����W�R2��ޓ�fٱ5��J�G埌Q'���� ���*+��x�%��6�NoyJ�r|�L�ٶ$�Q�35ѐ^¶�	�S��O�7��v��liH#C%JʢQk��i~���rLB�)�7��&��7N���]���Y�����v�^IԦ���T�	��3х�Vt�.=�g���3�e�'� q�ߡ\���"U�50ƴ�s ȷ������HV����\�Ue�X�� 6��H� R���cC�D��͉IoQb�L� ���̭����?dK,yO���!�^8f�����WL��V>�H>�&�s��W��IO����ՐA��	t��UHn���H�7�`�wN[A�!�6��uww&�=�6~��f;�3�9Z���0��=��G�r抴�s���V�U��[G��z�;��l�����ru��~���vHd��٘�ud&7o}�m���@�����I�|� Y�]]k NF�.su�Υ�[v��|Q:�ȑ�>�6��З����@|�����޽BQ��Y��4��B=����;�k��~�}�޹@�@��Hŕ�1Y�31�q��P7G���K�d�	lJL���jC�bD�8�}p�綟i/��#uB�����nNu��3��	�}i�c�}��<�̀a ��npƊ	&Y�IխsC|G*�����:P�Yb�l��VÙ&����Վ[?�i��B���[�ے��@��9S�.�m+B���7�����x�́R��� N�@���6����Y
�&�e��+�m���V����;� 2nRb۩Kg=��aUU��3i��o:�� yU4���8Һ�����8�'�֘c�P��Tj��u=_q���q��*���F��V��PE��Q:C��4���&�N��u��}�-�e<1��u���4��wW �v�Egn����	�DP�F��C�d���Բ�m��rm��j�n���y���7r��Z��c��7��Bxm�L�����A��̛�7l����6��5��a�,�L��+�ܵ��%��y��V�Ox�ɻ3�Q����i�՗3���z�)�ܜ�υ^v�c�˱�ɍgC��T�����ՆG�k烯��ڰu���"���^g7��T�V�gZ9����9��ư�.I�����4�#on>}lwV�-.��f�]��V�9���:�<j����r��iݼ��[�#��j��7��6�ƽ�J�	{������Z)�E����)u�L�h���ګ��I>#�y_q�>]�i �*��\��2u���9BN�Na�O��V���4��Yڬm�����ԍ m�� ��` � �`9c@ �r      � �`   2hl  m� 	               ��l  ��   �      2*�c.�=q˩H0c+Kڙ����L�j��Me�3W~؆wX���V�3c��h��e���;@�ǣw�v�yK�C	E�^�8� t"��V%hP�	%�	�s�#;f21.��\dG�n�����I�U1��d��^���eȫ��72� 9� �GjJ�h�û��hC�ri�,Y��\�J������'���%R6-#B�v�����PĩlĻ]���#�u,���bvT`bhyf(켢v�:B֡�8݊ D�eI=�c7wz%�M�;wE1a�QM$��W�����~�t�����WB�Ǿ�U��*orZ8������YI�M�+7�;lkz�2�d̃lhli�6�  M�lV����6�X�I-p���d�ާ��S������Cu�m����
.�n$�*%x+3��L���Ԇ��~�R
|��7ݺ�(�s(�#��giB~Z�{�F�Ǡ.-nǣ�h;�Jr���q#��e�\���7�M�n��*(R��^12m���.�W��+GB}C��p3՞����P��}�����g4�=D�Q���<����"�m��B������	��u�4�{"}27�k�7���uQ�E195�sl�c&�5��s�Xu���:���}y�p3��H���G�K�O0�9��^�����[�6��<��*�h�Q��*�WH���@4��ۊ�S�6 x�o5t�׺�w�����5��T��W�#/:�#E�,�$p����^��$��O(��K�J;��CT����nC*,Qլ�H��x�Hѯ,�� ̢�\b�g��Ľ^#�4�d�o
+T�|����-�>0ו���F���#���b��V2
����T0�6#?O[��t\����	�V�F��b�F��do�Lx���/ux�}�=^p���������e�:�����$P��pv�29��{�J�\����A�Wz����=�t}Ք�z�^Y*C��En�b���a��&�]����0�pb�I5����m�t4ο��ƅ;�~"N��<kN��Lps]��W<S/�sOvMΡZ�Gί���@�o�Ď�z)a�}���1<xX��7���¾�s�mR��9�Z:d۠�$���>5;3
H�|+$���'5�Ă����3�8MQ�k`��Ϛ@g�ճ��P�{r"^��~[� s�9|^��)H,P��qQC��S��1󏾖�Ƶ��&�xF�$<�`��絲�8r��	G�����-��s Lĭݙ���y8f��18b���a�]uAz�Y�9ZV��7�������ƸX��L���lc-M�,�Gu��<U�����6�|7N���47�����b�My�8��n�: z�c��z�t���y��v����/}�ḫx�\��T#�������ҭM+�~��������9�:���W�3�c�8zq�u�_�>�x�:)���>�Ѿ�Q�H�$��i���J!F���ʽ�_�2��k-�M�����Vj����;N�Γ]|_!X;�Eg �/M�wq!/��a��Fc���9��f\�e\fQ`Ή��F)��]ڍ���l�������J`j)&�m�����>��ۉ$�f�b�]d�S��]�n�(c�a£���c��yռ�' �|��O}���'���ތT�ɯ{L;���˹�V.�u�}�xx\��.�N������sq~;���x:�&Im�|���,��h�Ȫ~+y��6��Cv2��Yſi�)ׄ�γg�qg�B����qq��B#*�d��,�$����u0k�V��k�S��y�����+-̶� V��˿��wpi�(�.rG}���V �?E��媶.܊�����"�I���eR�R��"��i��0�$o,�al����핂�l߃���S�ln
8��u���U�IG�������y,��}2��h�U�,@"mH�Am��JR�;n�6.O��-�:��b�g���&^
�1"�>�����0A��7����v�t-��A�1:G
�X��Cᩭ]ޝ�h��0^�E�%���Ѵ1n'��DFs�_����w,p��O?m�;������j��h3�������w�Z]��+3`��]KW[M�=]��C���/Q���YD$�.�����x���5K�����
Ք;R�@�B���κ����V�;ePVv�;qo`�"u�kVʻ�����l�w ����.=f�V�-Y��.=/�m@fyvT���/g?�Pqھ 1C�E��ox���Z���aWr��"!޿.����Tz��ά3.6s]��s��Y��f(:�x!�0+;�n{2��6sX *N�~S"���Kiyq9�b�%��+C^�]i�{�U����D��w�+������P�`ݨ����4��p��GFuK;wNt�[��Dlp�ګ v�����D�zsEz�;���Ͻո�٘�b��Q���4�0k_����bd�aC��ݴ�%W�c�3�X��M]�E���+���ء{���*��L�u\�	��k���O�s�(=�t�S��]@��*Q��-����]�|���ש}��/'����Z�??]�.9+��:�׵��5�4��;墷����Ӄ[֤��J(?keɒ���z=��hD����/i��T�[�X��1�+��j�cf$�)1���zR�Ŏ������<S3��"�z��U�kd4xt��|�!���.
���!���o�AD�)���;��V�ނ}��O��av��s7qΩ�l�������Ck�Ն�5+���u��G�:�va�4��r�{��޽��UL���gao��2A��U;%�h!�r5%��.#@� $�    �`   T��v���xb��YF1Z]m�F%�Mt�.ĖC8��Ӡ6GA����-�Q���%k���=��ꪣ��]/��M����=�]�����l��+���n{a��p�_F8/�q��^��g��Ӽ�O��^�jמdY��U�+jqU�<��*|�5��)��#i�b���
��gظ���s{�l\Pf���fܵx�z�L#V�z������5ۛS�+�!L��:�ζ�Q��S�@����2c���vJP���K#{�+��_b3>�Ԍ��pg��Μ�ʁoۘ͠�0��X�����i��p�8n��
�<������&�OV�
�>�ἲ��q�2��=��J�wb�Y�rrD�W��$g-R�B��``��^��5��ꍶ`6s�XP���<�f0�ұ�8V�6\�=ǎ9��U@�3
q��*+%f�H�M���t`.��&sޜ�f�b��8��JuE@�����D;;E��ƟK{'��W�=7��L��e�;Cz�[ �Q����Ǔcr�d�<��"�@�(_ˎ��槙�b�y�z����\�-��Xj&����$T��O�pY��X�<՘t��6&��k�����.i�*�\p��;շ�h�K�\���V����Qz�!:ٴk�pju<j��K!�Z�(�\�WL"��J��ԝ%쳻�s{"m�<YN=��k�T�?^��7ý[u��j�Y�����Cɾ��p%~-ʅ��4z������c3�:���͞mֵ��2*Ů�o����L�/ΐ���Gͣ�W���eE��~$J��]z�7�y�^9?�G�����t|%ﻵ��n�O6�T�[]�<�891Y**�̻)���j��;_M��u4��O7���e����D��3�
�W;��nrk0%n�>ք���:d��<��[ӎw-n�
j�uR�mR9^>�	m�Z���m#y5���D�S5W���.�lγDJ"5�S, �z�Vz�W��*t��j6��c��\��V(����pu�{'+k������r���=r{-��)��W}vO;~�w�l�<��f5}#�;%��>�!Z5
n�����+/�����/|+7��艹*���p�����3�/�Y��|:����X[�z��ׂP�k�$Y��)�SF�s���W_��;�X�����k�6c�Yn��R���:{�ͺ`_�9Ǖ�e)[��w|�(�.eL�MћJnU<��i���Eט]�#8J�X�������G�9{]��5���eN��h-=g:��Y4�%:dun����d��G�Ue.��<�d�к��-�drn���4t�M-G<���.;O�^7�Ȼ�xGL1��Q�\�M��t�x�f�i�ٷ
w���)ڻ4@ת+k&�h�1c#�o0ձGA{`_���:)�r�0gL���hn*a�N�Ա���J����P7|_��JY�oԣ�=��^H`���~��x^�9��h�;s'���ך�}������F����1�ʋK�;ۊ�P�;�;����|�y�K�[>�,�튀<S� �ˇk2��:ߨo{v:ʪf������)�ן)C�͖6vrn0��6a�Of�)�Z���(��<�E��yfFmdva?L�S-@շ�\X�'�c�z��,?�����w����J1a��)W�������X?_ܲ��Յ�1)���a�Ϯ3D��t����i[�����i�Gnf�g�R�����=/�Z�M����`KMn#㶺���Cɰ�.��n�t�%��l��={�*9|���Ji��0\q�句D��&uV�����fN҈�ȩY�fùػQQZ����z��� %N8j#�F�/�����e]G��yV◊�Ƕ�<�����gtM���v�-	8�Lr1��X1ɜ�	�v�l�v􎳉,�;/�S��x��ݦr8��4.̵�/'MCzm۬�(�`���t��ǐc����p����>���|o�֌#�3"��[$!1F�No��}+Ix
�NY��>�grW�}
��\���t�b����g\�C=�la�w��7JF�L"���L,�Ը�FBr�J�	��*�����&�OG֙0C�|c�C��={����Q�_[�~�8}Z�K�܉�t]��/Jm���/}��]���ݘ��g'��󥸧g&�5����1\�8��7�)��o��m���ډ��F
H�%�x�^�݇���x2�_W��Q;��hF=�|h�`J��'��znw��<�lr9>ϕ��;.P;���>�Yُ��4�S��	�+�he]�[��>o.��N����W�+�/�=8���#�-u�j�ڋ8�uGuѻ��<�T�����Y��E�{ǫᐾL����}�fK�7 �q"���.�K�u�BkE-�8r}ǐ`ܭk+�ס=����^\G}`"ܳ��q��<&����^J�.x���س>�m	�Ijq|�p�1�=a�.�w�D�sђ���ҽ�\Q�9�lg�IyL���[��F�]=G_N-�b�{�!�p�`F���W�E��oi�˺��MY�obt�������g^B�kEN��L�ot�W��P�U�p�"q)6�B    m�  Eb�*�U�9��o**�E�iJ"u��c���wݔ��1�ª�	���UP�6c%^1�̃͜+y���l�|+���=�)8�3���B۴�2�����W��S�������F������f�٪�Ѩ��Xb�W���.`���A���ũ��>�m����*�������{5+N�f�����R_G����I�6�mc�Ձ�G�x�-�-Yѝ�F���O�QƢ(�V� �K�L"��b3���/=!̛��c^{b�hsw-���zĝ�
Q:p0,n��z��j�ܓv=f"��W�]3�������/�U����+lE	d�;��Rƌ�$	��Օε_=Syd�3�.�RiB�Ι��
�+O�r�p�$y@���:G��VB���H�����9��F��5�;�s^51Ir�Q�w�;��5u�{�'��#�`�Y�k8$E��<9�>*��H��0�ۆ�@P�)guc�Qz�P��P�����0b��G]�ͱ�,yR�/ڨg���M����Z����F�Fb"In~n����3+9s�sEH���xz�V�T�.�^��3'��&ц��eT+#��"��,>ӗs{�j�������Y�+yN�Y�R�11ל�lK,��1��)��D��l�=n\&M�3P;Mk�]e���(������(wu�WhOK���C��L[�9]����E����M�?�'�1s�,��lF��2S0�Ή��c}���8|2�vi0�lX�2>f��&h����<�'*$�^*�ؾ�=�ܮ)-�3-z���ᓡ��;G�5���ކ�w�̩6���_v���(�@^��g|ֶ���7.��&�m�=������{ѕ�n���{6V@8�#~��>��Wl���+L:4}�ƥ}����q7G�)A�'کQ�.�3�z�n�
X+��%m#�<����N⫫�5�����T�(˵�K��DZ6�������֔?Gv^RQ3Pd��75�$�m�)�:����o���9��G��Af�cM�GnO�]���{�3W:a5f�Bդ�+D,�n��z����Ꮽq%��3ރ%�d�'E�z4`��u���_?��}�{�%ݔk�R�ָ�#��d�<�S�tV����  F��X���N^^Tץz.c�#��Mh��4ћ�vC�K�|�����)��}���η���sԯ��hTY����K�ؑ7۪��/lY�uAT�gU��i3���%���ݼ&���u�#��Xy�[T:+F�f��-��x�WX�1PJ��d�P�Pb��/��`�p���{ZN�FX�ӑ���ܬ�{\�7�Ip�G�G��e7H�N9�0 �lDڮ�����r׶���!q�hST�;�=�C��^i�j�Sguu�u�m�q5�3I��a7�]P�]��X�b��v̾�]���9�}��2���`���a{��U2B��T�r��BZ׷���A�cB�痳N#o�ERV!g���'�G4ʫ���g�nԱ�<Vm�0���&���G�彊�U����=��W�3�_L�څ܇�5^�%���ڶ�UQ6�f��h�٦kN 壪��F�2��gM=�F��gj�#VeM[՜U\�jj��[�.���][���C�Աm� �!s�,�=�u�[۽SeZ�ͳ�ç��h�yP��8�6fԓ:�Y0�%�Fژ$�4�2���;5ݳ,�"0��f�I���Ӝc�>ɋ.Y����5��[��!���9yw�.�(�t�Ǧ>����劬�1>b*��cb��$y�U��Ө�@����5��;�ِ=Ӵ�&7s���O��Y��;����\v��7�prp� k5��or�X�*P�9�jQDT�@��r��WG9�[��\^a}>��:)'3k�}�σuEҌnM�wR�S��Px5�ۼa�:��6�ݚ�vwu�r"�j��W!���R����H��Hƙs��o8���;`��t�Ws�F)�u�9-��z�s�B�@Z-��oQ��hK<q�0�`�۹36�@��X�k���&c`��"�������!�b'�U�X2���y)��qWT��"�2G�(�}�<�{í�ۜx������]{�P�dNS���;�ӕ�{�h�d������-v���C<��{^k�����8����Q��V��i�>n�M`b�J��Zt�m����Q7M���F�� �R�tv�̥K5�f��a���Y;�k�UCN��8q�ү�Fm�2��������j��=��nW<UΥg[���)�F�י��q����nP�;�����T�g9*2������qٽ���2N��.������K�7�9\�)�6;z}�X��F��C�U�6��'Z1&&e�Zz������V�|��gj�"; �{�����\
:�Aa�K�m��{+FY�����H���Y�fN�|�K��0�id��Բ�8G��@y����ɍ�GwF[WyT���}}��3G7��V���o//f��@�v�6z��j�"���+��CSkB�Q��eۋN�(9Lc)�&cH]����]�7P�z�#���gUK�&��Y۪���s4?�轴C����tS��1]�S:mn�}�[rs�~��:*�)�����0�S�$=ʷ3�T����������|Fdn��s�=U�*�iM����u�'cry��-
�d�z���M:��eZ�sYu 8��n�[#�m,���~�{�w=�����xu=�C�8�PC:�`�8����4R�G~�F����ʕ�c����@�9��.*�����YLmڝ�bJ�i��=���ؗ^���ޞ���X������vGz�b�EZ��	���Y[�큶X�FZ��}Y2��p�㦻�T�[H/��kɥ�)�yJ����C5���f���JJR}���@�x�������C!yD�-�[s�j�x�����J!Lfp��K�=�����t���y�:EL�0��:!Q�~��'���ta<���5[�{�gn</�Q!D̗ho�J%��buo�X�=���-Iy��J6Ӡm^��������W[��oc=��Ϗ$�n;3Sb�����R����gM�������|��M�-u�.�؉0)����JV������C��]c��{���{}}֓�>���c!� ���|�r����t߂fJ�x���7���xVf��6G~vO\��sUB,mg�w7L�ym�����P3�z{˚�N�����wgA�[�|U���̀^ɹp5\h��^O�}�����h͔�k�Tī�Y��f0�pί�U�t'Sf�Y�}u��T�x�"e)}���W���u/�a���?g���W�ԭ�Y�[yH�?]E'��O���ki)�j.:����n<�b���U�;����.Sݽ�+����j�
Q/�й��xiV�YƸ�>;9��;?�D��O��<;)�K{�t�dy�4�.�|��r]#��2|��h�Yy
��\���]ug���(���S��~}���@��mt:&/;�E�lw�����=����s��dwm�е�sN�Y��n�n�s��=il��#�w ���A�&�q.xX��U��lI6�\Ȓm�����l    X<��?\��]�%�	�H9�!/ׅ�[YDnfH���FP��N�v��n�2�uєp(��l�t�[�v/��{��	[��-��Z:}f��G��_U��>��>�y��22t�ϢĸOEu
��뇻�/������
�h���?g���℘1�����Ӌ��	��	�~�5ml��L)����P�Z�{M��]>�Ϧ9��$����u�+���J�ͣ��F��X�.�y��*��ʴN��`X0,҅����kdQS��-&�36�j�s졝��;�ˁ��c�ew��^b�jL9�<wxɡ|�)��W�V���Q���w��C��Z}���"|�4�]��t�����-�Y�gU�c�m��t�>�p����.`맕���V6ܒ>6�.EZ�Ӟ=Ǐ���k~i��$:��+�v~��5�+%vR0N{�iW����Yt�w����E;�|w���8��^K���n���;*�>����k�Z��sZ"=�˙SO�,���|1�F ��<��-Պ��sL��5��H��I�`�|�������dY�����Y�z�Z�}M{T��Q���M6_g�W����e���]�;y�`}�� �<����a�N�yLt_W�R�p��������Q��Ip�;i�KD�=yz��0�)kػ��kt���Zq%7k�ʟ���+˕Л�tF��T��h{�5���Ab��1U.����[��2�C3�#�:�3���T���Bޭg��	���������=���&���l���/�P�g:���/��D{���>�[����_v��G��xp�d���Wg��ב8��[������נ���w덚�m�������a�FwUm�J��t��F>�^G�z��g�����^�ݘD�gwO�|���	T٭�H��o£��}ޏ9��=e>̄7V��U�'�����H}s/șܳ�\MɌ�Y��H�ؾ�ʀ���Ϣ�������	3/��z �;b����^�3(�����n�Э��O^P<r��z�1���^�W�9�������^���=J�\&���1S���aԔ��ٖjJS����%q��bD�����ɶ��>�o�y��7W�(\םF�*>�5N�Z;qu�y�xR���2�t�d�x�5�F�d��.�H/2u�*Pu�r'3�\���1��H��ޯ��7�<��93��7����
v2{=7��z����������D�C{��a\�f�,m{
^Z:_��_s��T��E��^��{i���.iG1ւ��ɿ��3���݌g5u`���G��¶��NGuW@Z�@8J��m�i":�ͫ�ιpv#v�|���d�&�V3��D;�fs6�-.Γ��)0�g�c�lk�O�=0zb<L����������[
]����y
�t�B��Ǽ�f�vȷ�� ��P�=Qo�\,3�ն�*�X�J��k����H�Vo�L��9,/����,+X�J�Q��l�~����T6�3����4̟n]�����4s�p�?��o�X�u{ <��\�9 �â���uϨ�U���R9�����s3�M�t�V�$�Es�}�s���\TPt�5s���w�\�{�v�%CN�*�-]&*|.��������徙GWാu,!��4�v�j�;RG����s7S�e_��z���sR�ݩL�'����/VQѴM�]~�<3׈�Ķ��]�B��Ɨt
���&�v�D���2WEe�ͭ	N��_��������*p�;��cU7E(p��%� :��3<;��6ތ=S��/� ��ltuy֜�Ŧ.^\L�Qn����4��A6��z�>�]t5���ꧬv_tBr5b�3��V!>�����_jy�F���CF����]�<��9x����]\�9�)u��K[�V6yC���݁Ky*S�B�sz��t8�j0U���iQu��Go�����u����:�{Z�z���5+&rbX��g��
���ﶎ�#��T6�]�����E�ei�V��*����v.&8��x2�a��ϵ</f�D�bw�>���9�(����U�?d,o04G)4��p���l+�*}���})�8kuo"�6>��t��S�:�c�ޮ%��.4�(*�J5��J��e�M�8qr����4I�*a�aV�@����G,ܒ�-��q��pc�}�կ�_�o_b���s�;9�6�r!��&@m��m�   ����u�Ϻ���&\�&S�b�(<��;d��������T�o�ls(���2oN?kd����A�y���9��Fw�D���
;b~.~^���&}Em������Oq�{�xk.�.�s>���Ds;���Ah/��~�m{��T�+�qӗ�����$���7몼Yf��P��a�K�]ك0�Td�v;����.%ڼ�Z��E<덕B2}V���zڇ�Lڲ֚y�D����u��>�c��LsdX#3X�pB����u�f.3Y�1V��/�Ъ�N]�h�WN����]+�@A{�	�_׎����br(M�X�K�Ki����>lp��sU͋����9}z���5?K���JSw~8�ۏ�����;�&ylvլo��k�PU �n�͌D6Rm�L�B�� aU�r�3ϵ�+�\���p��v���M�:��ϫ���b�/�H{�7���8K�VG�i̥Ȏ��{���Є]LrK����as;u���}ܰYͯk+*t���r�>4;#q=I���#��NK�5�²j֡�3j��H5����*T���Ö4�/�w]g���{ך�����Ly�]UMb����=W:w�*���ꬤGn��{��f��HbU59,�B	nr�7[Y]ѲJʲ�+��Xkq��7�!���Y"5�_ �,���Ȝ�ykrb����dr{��_Y�($z�c�F(�
�C��[���j��>�ۉ9&5�Ed\%��Go�,W�]�:�޾U��*�W��+'���[0K|"/w�������z�㈭���Hd��*�����i��%o17v[�����m�=�}C�^�f�V<c�3�w�V�O+���f02$��'���m�@āH��E��z2(��@���|�g�ނI�De�Uz^�a�s)GA�N�.�z���l�1�xVS�x+nϰ`a$�*��g�s���C�>VL�]�˿�o���LZ��-�m��o�����T�xT�anqy"G?���DZ�kI�ue� ���e��3�BT0� �vE5*��;g�s�}ni�b��w�#4��2�2�;;����^�M㺏[���N��U	�)s���h;Yx;s�#ew+.	��gqԃ]C�/��K��C[��绅n�2��;8��úsy�hL.�^�����fW.]n���v��sq�=�r\�d�����b���;8^z�][�W�~��ΰ�zgG�r0�͎}��±����De+�ݍ���Sآe'���+�U���9G!ے�KҷU.�����Z�g�Ey��B�]����[��]��ޭ��FyO�y5�K� ��݉w)��ys�T#i���l����fD��'����M�x��{�h��G��G�:�Xj�ѫCN}�]o�=���a�#�Ëwt
dR����S�_[�f��rȜ���do�˯zm҂Ŕ'wl�{�}�>+(1���� ��^�s��=k���\��ٴ�ԛ}97��i[V�zg��J��N����x�P�G]�*L�Oj�ti�>ģ1#U�=�rߛ��Y�{Rq�\	q'��8�̏9Uɇ;�����7c�=�8#+�Y�3S'��`��e�Z[�ٙ@KR��b��x�9�*%C��7�t�����ۺC,�o^�j�Xif��7?6�_/��b��ܯE�9�1�wݯ��R��=$ڜ��`�$n��q���k�.�~��=�g�{��{c؉?.�4�����"/<�P���5���7����L�Fmn��[u^bӓ~)����%7C�  =J��ok��q3o��߻]��.R~�=���=�d��j���jl�I�3
�fr�<�u�s���z�^�a��W�&8�C;Y5����፿Sٝ^��s�m]��ʿ�	�g�6�1�#�=�3��T=��3���2|����7k ��?��񬽗�fՌ��x�p{�n���b�n�������,̂���=�|aQc�W8J�����1���t�^�O��oo� ��y��W��Vw���
�&���W��+n&0����k�;'���S|2�:��V����������
���w�=�ie�d߅bVv��wS�N��}���Ԣ9�ѣ}�Gz&�o!U���<���X"]�i��F'��s�N?�G�}���f���vOwr�[e�B��m��t���Ύ�VYqWU��WB��7�j#��s7�*��ʓ��IC5TK-�Eq���F�4�L�����rha��9����0ê���R��(̆��y���f�uS�l+��j��[�N��|g2�P>ry�)]+v������\�1p��Ӌn7@ц]Ҍ�ԇ^}����B9��Ol���7*X�^l%F�%+&2Vk�ī��I��36E��ІmfC}��@.C ��/��u��<�l'.��X*��p}�U¥Q�z-�:��ƻ�p�q6��E���g,:*��bk�SW{71>v�u�����f��J|Y%q����7�����
�xuK��V�f�G��E��$l��[|��6T���*���W�kw����;�;��wM�}u�D&q v�롏�9�5���}�՛��v�2�gu��װ+�OH�J:ܧ�tv,DF�z�M��=�&�Ĩ
�V��P�*��E�_>��y�ɺ�/;v^p��̶���v�P:ܽ�-^~m�J��|��O �"��\5��ĳ�k:Z�݈@n�M�"wD��ۮo��h��5b��P꾆�+4��038�Ӯ�h�o��Ìκ���u:�o+Yל�qX�^���Yӝ%��4�ܑ�\�%H�1�r��1���+����˔�u�=yr��}ܬ�]h�}�ndy��Ce��f�ޏM�/|�V�V�eIab��fJ��sv��\��NEj��?=����C��}�6�������
�*5�Ju�f�nsB_X�5���N��a6�B���ln��ᖰ��X��]b.��NId���s7VB	��u�R��o7�;ƚ��;Gq��f�3�T��ud�x��yC^��l���ɧ��1��0ӕ��Պ���qێ�㣻�o-��4լ�����f*}��ݍ���U�깏��6���Lӑ%f�+��Ղ���:}�Zuc��(�Ģf�%i!�vO�w�F�X@�B7�4��s�n�2�E�k�
�p�no^;.[�	�]�X�-��q���=�|s����;-D��	���� 	d� ��  6�4�0 �m(�0 �     ����m�m�    lH l      m�    @�         �`6�  4� V8aQqO�rJU��o{1tfWS`䂮m�V��We�}]�SݵP��z'\���ߴ���[cGM5���,��R�kk�s@�,$V�=rUȒ,�M|f7w��m @m����l�M�U��BKJ���m4�Pxr�R�Rl���Z86mn[f�|��0�0 h_��ۨ�o�����vD���=�5���ͤ��3q֒s�s�-�b�ƣ�R�Y�Gp̋I66v\�*ԫ�]q�[�"�#�@$t̛�doWU�n��˱�U����&�9Ȅ+#��AX`���y��|>�ﱛ�|5�}�5�f�y�݉;q�j�82A��u@��q�^4�R�r   m�  � r�.7��nֹ�U:ɘ��pS�X�(�V��iW6��P�5B�r��J�@��^�ۥp���ٽ�2�;�S"�)�>}g�{잡���pn>̌F���ww���;u�����	�;߹�$��x�A��W�ɦ�?�2?f�eQ屻H	>̖|3���v���7g�;�w׃������w���R���=B�N/;��v��=���
2�/��=�J���U�VN�ݾ�J���"��n�c��s;�6�`�-�%`K��Prb��������ߟ�P��l�y=.'{����/�!d��V���S���=�{>�_�y�h>P{��jO�w����~~��{�[uB8S�s%����_/�]�|'B�S��;N�㸵}��ɒ��ߓ�Zļ׭�L�E0� �{*�_�˅?I_:�{�j��F͘��N�;nJ�O�5�� 	�6�aو�����J��z� Ɲ��p�E�%�Qyn����W���t]���K�������wc�W8\�$��-����)>��
�rEϝ�wP-�v�v@0�q��/� �!��Tp;� ݼ�y��1a��E��:��FU�\s�54~O��ި�[��w�*:�oe)����zD� �wRs�w-^�T&�X<�u_�f�]`�]���b�K�1�$���]r+��w�ijw�<�}="ܨ�7����r�o�~�u^�m8H�'!�ܛ����)u:�<����<���ף:�og�e��Ԝ{uMFjZd�'�F��%�4��l/�y��4�h��>(�~���vO0QC�r��1P�*�����j(��ʼ�' ;��5���z�N�k�M���x  S�uSN��:�ϟ����Ga�L����ҍF"���;n=3g}� w}%�TNz��$|�f��=o*��.���FG,>�E?I{���,j{r'�^Nm%s���	�2����ö���lV�9@Zp�\;�/,�AS�y��@�m�ύLV�ڞ��)>��<�z��`O�$犚lK�"�d�y��5��偍�V�d�hs���f�IݻX�m��.�@��I�YZ�k���f.hC���X�hܜ���jjRv��U /{%���Pc�U�fY}���"�9v�y��F`��І�{�9*F�ӯ���OjZ�x���$�sƺ���o�ߣ��}f�{֦l�,SiűB�zOK��)�
���p�a~����VO�<�b��H�8�e�7��N0Ўx�|O=�O�k�1�X�����q�Lyӿ.ܡ��{����8y�܄�^Zߋ�7m�Cw/�З������ER�@J��$�%n%��~���}�yYj��F̓����/r�i]��5��%�����m��\JWlH��
+c����Ȳ�O�}݇��A�kv�ǜz�[�#>Z��	�wA͍�9�����"�9X������׃���F���7>%ax�^��Q����s�W�>d!!�&P>��P(Q��r��y{�ӭ�	��e�����L��]�m��c-����I��3�۬�>��|*���rq{ss�[^�Z�κU(�1�s[�"�գ��/��>��T�=�ѮEd	�����:���נ�䮛�S�E]X���`�;�S❳W,C�i-U��|���)��1�dwa]㜆v╒����Ӗ,	�Ku}m�5Z�Wl���n�v-�ܽ�|��k��ԣ*F�fw�{��.:�������|�v��zM���I�7PFէ��yHwXr�v:è��}���$��T}D���B�7�*�I�E�䥠^E�C+^=&����}���6��C���^[����̡�ȸ�����8�hU�=�󮑓�[Rwrn�W>s��f��z� �cԧ�.��]Gc�9/�?e-4+G{sEo\wb�A�V%z�����'�YT63�_l/�z�E{���z3;{�c�-�7��e��t;����Z|{lU�H���K����"��J��+��uv-p��)eßZZ�l9~�^�R^ɕ��M�߽�\T�R����Φ2U?WG���D�Q�Lt�M��d:@E�z35�r�(Kͯ.0��jo�gV�I�l�j�v��0�2P���#$�uv����_,���62'f*�����mn��+��{4�+�y��3�i�j��3k�jE	-3o�]�:�Tb��\�y]���=��	�i�حn�	�럱G|���x��K��p��V�F^L�cl� �d    m�     	:����|wf#����N����%(������I������ 7:�h���o��#��>ۑ{x�1��ޯh�lm���'ʫb�%^e��j��s#[�ѵ�7ӯت;[�z�}Ӣ�Z����-��3�s�Zsy{���NR���v���g�f'����Yuj\��߽tձ��q�]#)���(��b���d.S�����#I2��OJ���4���g��⻾���p�KZ��T+�D׏�T�(rײֹ��"��9��AE�+4:c���%{z�{*sӼ=k\��E� �]�;�Js8e�{5�0�ޟ,���u�w�Y_`�ޜ�a�ίn��{Q#h}��^��d�>�W��T��@�I��:�^:F��rF����6��\��m/��͹��%��3=��ңQ/EWz���Bȡ޺F>�T���[��n�㵙C�j�m{�'���dfey�Lh����8ߡ�����Ǻ�%��	|��)SC�fq��S�C�gG��qHT�ݑ[�����S�Lu'���e��~��zi�z7�`Q�o�o��N�:�f[*'�xZ;ݝӨ�m`]����k��)��GW,�ݕ��<Y}�-ޫ;�{����88Z/P���������߮jU�@�8�_}6TCe�{=S���I�^���F�߹^	�#�+"�����aY���:������zJ����B���[��8�3�:�/�2�/��F�H[�7�?b� 7����Z�>�gh�ALN��c��g�sQo�=��_j�|!P�k0��LL��ĥ��U \hBV������N�WVsQ��I5�S��+S��]8m��J��V��ުS�9*���c��^���x	��$�ĥ��
�;}M箵�l��i�x땉]l�R�w���C��/<c}W��d߄��tv����V��U�k\C]�1�\�˪�םKD��k�wds��qNT��I�¯��w�5�>[�}�}���S�H^�G��:��9�v[]S �>յV��ϖV����%�ަ0���u�M0CKU�{X9v�ͬO-��k?l|�$�ѷP�	�@�ݼ�k�,g+#�:�P�tVm�٫�]S���e�Nu����;�U������_�/�.~�Ǳ�ڷ#|Lue��vVqK�����iӅTK��ܣ�x�4g"�4�=5�2#v'#�"���Lj빇���Ύ�����'��sO�s޼��g�e�u;�D�7 ��{�]�g�[�C89���qY^�c\{Ʈ4��}}�3�^���œ�Eh �Π"�RªK<ޟQ^��i��>�J��S�n�H:�Sc�b�r2�jX�!t����ޘ�u���Or�4���3�]@��:.���˛r�Mb�e���$�yn��g�!���E��_���v�\����X~����Flޕ䡹�qұ����3dzn��i}�+@�v+ڙ�h�pَ�M��*y��ۿU4A=��^�6���a��\hsn�����f�f�Ʋ��3���;0�V^���>�0����b�x-Y��c�{�g�;3��hNk��2u�#�ۘ3:p�K�\����ɤ���2�Vn�Ѷ��6��.�gm�r���]\�ڢ�7^>(u��pVwrZg_M�oKw4���qEC�T�0���s;�'yH�#[
`�Z��K�������r���G����ힽ�9�W[��5m��*�m:�1�Ž��,F��^������a5�:j��6�i�e!'�3'���FHW�ӇqV����x���E�7������N��|�߁��$�=���Fz��^�s��lmF�r��U�m�U��Q�XPzvӚr�HG����7�qL�y]�5��&� s#�≺z����B�N�����<�1�E��8��9�Q����f�d����^5yO-t"�,�s���͔2{�A�����S遌'p9��Y��P�����b��Iw��v:��i"�V����f ���aU����}�i*��\�+��ܪ�3��� ����\h
�~_p�<���u29��������.���c��ǻ�c�ᝐp$Z��Y�^���u����Q�F�
�>�k���T%����\�b$^oh���ɀhGb�+(j���It��L�Ym8jm��8&�trݦk<�����6�|�������� $�&f�m� im��   %�+�"}}�5G�3�8�p.��ܚp
��Y���m�3��H���)v];�3�k~�F�rp���޷���KҔ /���-J�ީ�Y>>X��.��P�F��퉉8[�'7j�+F ��¡�ss�B>�y����k�vzC��x4�kp뫌'�Y�j6�{l�Fn�z;�U[�,_ �J�/�O��O��B�Q���Ԣ�n�����S�{�u�l����ػY���W�m����>�*�ͳ!������;��=S�����s��5���Ο7�۰��'t�T��1!�d_�(1��қ���a�ɛ0�U�f�V'�Q&緰c�1Q��j-5h��'�>��<
�q��� �8� ����c���B��k$��&��/L��s��m���|}�%��4�=6�J͠ƚЅ���V$��-JYWW�9��}��ʎ�����7�v�V��Y(1�Y�W�Z�ξ��Y4�\��!��N�-�-s�gR�����hY�
�S�����Z�I֕2y#����f�K6��<�d���]�R�)ʢ�bf��R��=�Ml�Ab�ShJe:�"�nDr��I;1�9R�|�[��E��,������G]�P�6�G�|5o���􉽛PŮ��z~n�m!�&��ϲ��ȋ�\UN,��?LI�["�SD#0e���T΋�l�W
}��)��-����|� ��<w^��H)5�4�Z�>b&k<{�N\c�SޱU\x�k*��ǯJ��~\���*]��Hld+��r��ݭOVl�8��y�h���6.ZӇ.�_S�*����psk��݆O�WF�r��uG�`V�d�ʏ+S�n������D45�w:���=!�j��͢��7NRΠ�\"�V4r�����w�������63:2������P�U���q~1w]�\�k���L�B�{�c{�{�2C����34�z
0��D���������X{[3�L��.��ZJ�y(u�ᶗ�蟓I��7���/(�`�c=�d����2��=q�dXp>���[[Al��c�WuM���6�޶u1��y����0s�I��U�@�n��f�i�k�j�[���us,c���\f�
��얱J��\�5ƗM*���vc�(�sr+��໻��Cj�Eo�y�(�fP�/0a���pD���$I�S6I�)']DK�`9Gv����02���7����p_ov��jf�x��:�-�ɧ۝�tr���`vp^��v�1;.����}W����[��D(�e�0��ɜ���ݩl?ot����#��8�U���ԠU9��-��K�%a����D�x:�l2�� �9_�{�~��"_6�R��k�r�j\��J,�NwF��Mګ:�C�jeA��w�ld'��j���ݪr����'����۾$����9��jm<�8#[Ξ�n�|�Jm�<T��Ris�zfʃ^T׵6^i��)v���J�k��p�1M�+ޞv���:���̌-��nX�V+i,��^w��ڷ�#-��R7��@ji��V���^%۔P-7�OO+��ы;�l��E����{t�׍ע7gg�M�l�d�qZ�\�2��X�~o!���=wn)0 �XPUP���w�ű� ��1�5����FFwjF���h��]gt>���|��EiɌ�ԧ�f�  ����uX;�.�Hw���r`�Z���jṅm>VGL����kR���sz^�n+���*��%���oٹ;�G:9\g/���e0Ⱦ��v:`/���䆥��l�(�ôꪬ�*0q<ر��֢������/`�/|0u�귛	4��b��a��
��}��8p�����r�*���#j�5�}K�"HfP�_v��ɚ�]�5����7�4 g���`��k\qd��Օ�2ɊY�y'�@�I��9�FW~5�C�ȝ�ԙ]��wV+L��u��2s�qM3K��n��cʆ[���3rˆZ+����7DJ����0�[I�슐gI�����us�`a��)��#�u͔��ˏ�@�on��tU]�Z�Q"��5Ɲ|�溌a+h(��{��k��b�V#߯�	L��3�R	F��m�:�AvQo��K.l��wВ��6�9�;M��Z�Z�8���v/���5)[p�=ױM۬���;�^�	�i�R��;mpޚm:�c�#���ش�7.��8g�v�ߥܣ�F{�,2��uʞ6�t���;����/妬0mQ���Ȍ�Kt<}����P5w֔$��d�� �(����42�!�u�C��]7J��wS/�n��	Ηױ�nR���>��W����o>���=|M����1��*+M]D�=S��L�s�-+Oy��{���Xݝ�]��G�>u�%{/ɨ���aw��Î�@��0�d`����ǡl����&���P&�������V@�ܘQnW���f�i���ΰQy3�rл���־��{]�+#5r�Zy�)�v����>����Ij��J�m��t^����T�ۚfP���6���;���|<hz�թ����-.��pmJw�/�����g/RF��?6:������p+&�盝�F�b/��.�(:�T��~6���v�jB�YX{�RD��p���I�FUL�}ƃ]�iͶ hKˡOl�x���|	��YR�'b�Cf�>Mҍ��{3������|B��y\���[�-���Zt���q�6�:Z�Y�gR?�r��n�u���]�3���|c�� �M�y0}^s�2i+����^ٝ{��>�ˤv՗�/T�#���e9�]�}�4ipNV/_ў�7�����rMtsTI��8�`<��*.���WuӎUѸ��R��vB�Y���CMI�igcb�7��l�f̝�u�T$��3�+Ǣ�����~>�Υs\���<��٤�����V�V�3�N˼��"~ؒ�w+��9�b]{����?Zu�NR��/빝�b�]{I�X�M�������G�`��.x0�����i���*�O*�{�Ms�1�H�^Q�<�G������W�{�t��B�g}+��`l�[���=�����	{|ш��c�yPb7~��	j�[ZҤ��o�/y���-^��J]Y�_V��6�P�+"hdZ�K]�}K�b=��y0�A�T��U�5���w�z��ļ���X"�pǸK3YԆ�/zsEZ���Cl��;K>�%�Z�?|*�Y���D����=��8;�W���F�sx����ɍ��w�/��O�k����]n��h!wg�fj� �r�a����:Y�+�攙����$����W���b�۪�v�H��nu��pI.�mMFj��J9��$32�� 6�      2��+��v5F���RŖo/@6(��A��-��,ܝ3���H-��ɺ4VKH3���D���AK��-r�K��v�ul�ڹ��ȣ �3��l�m��}��v�UD�\��p}v�ۨE����lY;զ��sߌ'3~�_R�[���xΨ�{j���c�IO�H*���x����G�n9uo��"d�ˌ�<oǶS���3�{��"�M�y'�({��hs�g��h`��~���㌭�N�\JW�л!���@gy����Yˏ|r�o��j�|"=�5ꞁ���M'��*�.1I�km��j���c����~���@ת�Ǯl��c�N7�+�~�Z=�{�1��}x���KK�>O�4��n��}��S������F.wh\!�Z.uؓQ�[~�U	$iz�̛��0�R��ں���ؙ�W�I˥�n�~���tު�j�Y<���|+���Y{�P�����5KV	��1�k��H�K��a�r��q_���^͑u�N�m�S0�����W����&��\Ls�ж�]��E�}�$�0ڛ`�Զ�/mJx�5ٕi�Š2�.���cP��s2�nqV��bvu�9ا}`��m�ew�|����E��GT��iR�3S��{����Uا�%q(M͏>��.���Re�'K��U��}P)L.�N�s���J`w��gS#f*6hלr� �\KMg�"n�^l�[��+Ñ��lV�S�g+��Ry�v��}���������t\Uv`�P2/r��K������/s�_xۧM^���u�霓l�42��b̋zl�n�%WP�k���Ex�ܴ!�/6����18�/��C�=}�;�5��U���?@V�d}�RF��� *��M7o����dmU�W۹�m`����	�T��_�f<����q��z�cĜ�+���<�=sߢ���	�U�^ݵ3c���V*�I�eXʸ]��{�rj6}^�F���#ۛkP�$[��؏{bݶ]^�
6u�>��[��b�w)�0JY��s9ݻ�&��oxo��	z���L���C��W)q�ĸ�Λbt)�,����zQR؝}f믙�HE#ێ��ܠe]v�g]-wU`
����4��wˇj��hN��]7�E��rwsY��{1~h?�P�J�YWV{��[�t�ԕ3]�ag��,�~��jB�Kz�?��>������*�kظo(�����y�%��ey�,�̉q3:w&��l�Y���\��n��j�P�y��f`�玿\yķ�*D:�DM��~ګ���PI�j�nm�y�K�&Q�R��W\��7~��j"6k���;T��>S~��5j���~���#�A���/L���nD���N�£�z2��ə�_dw�,���7�F�b$�%j�ʥF�tw?l龪ŮA�5���:���?>����]L_���V��)���M��yt{�O^q�#��|�՘"�8��+�T��aN�ڷ��Qs���?�f�j��	�cqܝo�E��͇��%"um&\�L�/Z�u��M������s�*���չ{u����1����[���DN�ê��p�c�7����y�AG���/fޡ��d}��=���)_��g�zu�Fq�P�j�S��e�1�5��6����v��z�tI��2D�Lo)t�N;��d��8{�F��C�z^����u�5�u���gU�SrZ�)9�f����z&�ƌb�86Y��1s�E���7�j�vo��v�g�_��W?��.�v�$�>��P��������rr*"��O�+�σW:S��.^EOK�$�� -!��-K��s�mtK��Jı>�֢�;im��#������F�2��b1xO:��O-z�!Щ��ky��ukp=W5$80IΏL<��,!w ʾkv���~~�bBvz�۫�}��]����c�ա����8��R�Iy�b��
}{�yA��R�:��c�8�n�e��9e�I{El���@��(�ڄ��T��n4�#�x�	8���Sԫz�T����E��%����u�����uo�G�_�{�]�	���V��i�nyr�&gM7���j:\'�^Ҽ��W�oi����ۗ;�r����w�F�ep絜Ll�V,����&$k6Ǽ�squ�V\K����!e/UP����j�l?�W����X�ň�ͪ��~��'*h'u]�^��'lD��2��-����p0zݗsU.g(D0!�L��`         ��V���9�5��9l�dk;��b����:�M��ۭ��s�0 ��S誢�~�S�7����л���U�&��Y�?�	1v&��՗���.KޔT)��_�*'��*}��K�Z��[��s	N��0lW�����%����݄�۱������\)�)�l����k�1׈{�5�}�����E۞�:de+���q�>9�V�Z0����u-�dV�+t=n���t鲎�Q�=�])�,���b��vE�U�ŏF���2�>�W���y�����,M�A�S>z��9��ճQ%��;a��#d3*}�PQ6��)�u�EK]�r���>^�m\�w�cW!%�����){�^�[�s/2����u,��cOF�J���W��Mh�^*i���U� ��m���娑Y���t;}�3��5����!�+9�����Tpҫ���]�Sy6���3*j����̜�����PR��������}���d���h���=��^�ϫ���s�R�s�ÐԳo�n��D�S��9˶=��R#��c�fVLN�#ȯKv�b��@\���c�oa�y1]�ջ���66���x�\t"��;1_M����U�[Ǔ���,��u}�S{�1	�֖V:��Pj���k�G�>�w���1;��Wx0��W3�%�E�yύ˺%�e
Ź�|��jtC�������S�>�(�h�Z��k�Y�,oJ��a�}uF��AhǍx�^��W�;5�>�)o8���6��{H�x�����Ee�xs=�F���}��yر~�sO&i�"��[�jI��Hؚ����Ρ=���,8�mж�)z�t4;��M�Yx�k�7΀ē���Q�������+ոV�ۤ%������^z�����ͭ�4f)3���r�=<�M���i/���a&��E���nU";�c�x�g��Y]�S��z��M��kg�������6ϻ����O(�nOhw}��?�����.}�pB=�B�z���t��z�2�
������pq�v:�m��i��vE:��X�$`kc=B�]�Q.��m'�o���Õ�����}Uw�5vظJ��Oo0�k��Z+�z�Fi�t`����x��<u)uJy���pn�2�uN��~�qq[�������ǂO�|�:}��F�!�ڪjjK�Ѷ��8(_�sp�v,��o��s�*8!�۔ϺGj����/�Zת��쬋���npW@�XR���j6��U�5��s{���m�v�?���^����fp��!���Z�_�Wz����Wbg>�"��sW�L�U�=�.�  ���r��%�b�����z��.�;&\�J�q���wQ �rT������	��se�\c|�eٰ�X�\�ɺB-Ҷ������B-�W����@z�zzv<�Z��eL-Q}�߁�L����s	X&*����v����eR�W}-p�}�|a��A��=o�Z&첪��$ܨ�z*+�`�#^{cЈ���Ȼ^U�Wy.*�5~yK9��>���?Hw*󚿫Uw�F"ϻ$a������u�\X^S�Ț�ߏ�o��}j���V�73�L
�~�r/]7�.�q��D�%:��V�Ҿ�1�ze>2��j�U�zƷ���Ge$�`xcs�r;���.H����lH��c����{6-��i�6���6�5w�7N�Z�sf������U�ج4x_�����ˎ���I^�UQ�B�6�*�؁������y��u/B>�׿����fҠ8xD�r��&�&^�v׏Sׯn�<���ӌ��s�>ތv����QvK�x���u��0:��)g��2��r���C�[1U6�K�ſ>�ϰO��W��wLo����4�.N�OaH�*�q�]"�M�v(�m��1vk��y�_�k(��/%ϔ�{y%�W6�DR��<Ҧ���^c+��8竲�)j6���%J;?|��E��4o\
�wo#����yG����32��ʥZ9E*�G��^ynm�� �g
q���;��`��������>}ʧϑ�/�R�%�]	h79AZ��Uʆ�ŢF1���f���բ�}��ʷ:6��ߙ\���:�|����{{%a��ޢ���q@�c4�����qC�t.$j�<�#]���)n�uU�&�����:�K���kZ���\^0�	�T�Bs�6uݫ������Jb�k���.�,N)�7�-�n��B�<鋥�9��7���_Y�v+�D�y5\�N�v�L͙��1�C-
Cie���E���qh�v��;2��v��a����%ݨ.������Jڡ�|s��Ý��UxO]�M�z��n$K���wv-W��Ž��Y�<�f�6_,��˦�U�ؖut�k���O����!!$��� �?��,�$�����Y	Y Hc	BCI $!�@���$!��		���B$$���� BBI��B$$���?�������� BBI�������������������?��8��J	2��9y�+Ƃģ�-Ge6��I:��������r�(rZ�-�dj�0DJ�kV�i�"㤭��W����sr�Bc��4�Hj�Rn�X��eg큱in(����`�3u,opK�h�*GZd�)V3v�^ ndz�ӎ�!�e[9�\�uKCn�$�  t5�J����oT0��0�A^�9Gu a.\T��w�[LG�򉲞d�,[Y��e,�.��lv���Ձ�n���t�X������QXZj�\5�+C3*Vp �d�`r�{��w��K�R�a��,C����Cg]�mXs��ݴ�xv��H� æ�]/�T���ݐᶕ��Z2�`,�M��T�fj�f�Ef���c@&S��b�{�5r�C^
�b�TA��jز�B����\ ԭ0㺳��b-kU7��R���e�lԀe�\�S
��t0:H��G3{�K�Vl�G7j���q-:��;���dvF��7w[G˽�I�d�f7�i���@�ZR���P�v��������R�sS��h��*�Đ�6��ԏ\�
���LMݚ�Ԫ��3t<�bc��Lb	��V�'"&�,L�T�xZ�ax�	2��!7qq�8t��qr�4��������l)���m��-'�rŽ+(�j��6�͵����(��̺��+@��d��/n�iUe�,�R�˜�74
'kU.���N��M�9�%nS�
�dd�⳶�ǷZ�N�e��Eh�]Nn��M�M!Zj�^c��YZ�nr<�Cz`-޹����֢gtٷ�R��*�w9@�qG����Hr8쥙k���4aݷ���nI��������*H0X��a{e��)���Sm��Q"ɸ��l��r<(�I��S-�ut2��m���*̨[�L�L���;XLP<��h�s&cHI��F�*��Ԭ�e;�Ѫ6n���Ձe夣�ǅ���	�h�Cemn|%[��1�KTL-�A��t,�iރ��GJ]j���kA��	mL�F��{k�R������P�AWx����wVcT/�fG��a�
U�ͨ�f��ri��c����YB��y���l7�`�X�D�FLWF�CHMt��ٸ��ȥ(�&�$U�WY��T/O��xѲM[�$\�n���f
�M�"j�%8���X8��GH/M7���9�h^��I$�����c4o�.��4C��͓Z�7o�s#�d����x����iPGn��ٴ�&)H!�\��ؼ�t�e]]na6Qqq8�h�x��7b0�&�5�= lV6C��bضQ9FX�b��8
�q�@�Nݦ�]�YcTE�Wz
��"�ol�Xn��ui�v�fU�����@]QJ^���b4���ІA���Z�t��\��@�Y�5)Yq�J�`m֫R4�^B���rޫ23.G1c�;�P�hO23�ᐊ2	���������T��~�a�X���Y�Ҳ�0��sӛ2��WTYvYѹm���I4�wt�����J�I���s(��/
������*6�V<w��Qܽ�VF�T�,8��	a�r�Ԇr���H�/!nM�h�{�莄��)\wSYI��_�rJ�pH
��[�R�-�����$����w�9����0���1j�7b/���S0-߷0bk!�wv�.�mI�q%T�	�.�-��5Y�X�n ʕ��wmK�3�� L���{�K���r���awP��dWyM6�[��ӟ̲nU��X+�E�2��b_�b�Y��T��uQ�A��/J��l�?U�$r�n�^,"���ek�h�z�V=�-Zq^��Ɗ��MV<��E���M=wOp���G%}��1�FMݏ\Jd��u&��N;��/p�:�h�R�efD�Ǆ٥�ͻ�+,5dc.*{Z�e-�X��H��䅳m�t,u�����I��M=�ӄQT�c@ᵲ�6��Ե?)��۸�Lq�鑴���$�a��t��R�@\�[��5 ��l�ɀS���Ts
H��"�:@2r���֩ޅl��[Z��n���p�/��n�Aj`�g2���:1�t��w��	�cK�#录.�p!���(Ë�{/Cۡ`�a�f�lR"��nnn�n�D{w/ĥ��f=�E
�e�鐰ch���3���T�ҷ#�zi]�Z�,%�.2�m����� !(࠶��cʭr��u��f��-e׀��kÎ���U��	PYEA[/�Z�Oۖ���'t���Fb�ɸ4�	j�9{!���2��Y�w�eS���y-�xm�V�9c7�F�f7ADKv�#d�ٵ{4�6Tɏ� PM	e��˒�!ԛFN]2�T���c��Uʹ6�p]a"D��H����c�A��e���W�����}�$�	 !	#I @ 2H �@���FI$�,H�I 		$ I	$`HD!$� �		�O����������_����@�����x���~��@����� BBI�@�����H��w�F�!!$��l��ߵ�٣AO���		'�O���$$��!!$������������~`@��������������k��s�?����e5�[#�
�� ?�r 	 r}�$��J�Cd�m��jUMK-kS��f�F'&  ,�l	$WlEl��m���� �kbSLFSEX� �I Q)E(JQD
E@$S�T�DJ��65Q
 4 q@]$(R�T�UQDEJQJ��%IN�     �i�t�ݴT5v)v�u� �*�JR�UEP��Q!I�      �����(.í�� �}�

��5鞆4��ؒ�vbɝ�YWu��l�[ܯw���{v�]bQh�m��.����+��-���c���Vڻ9Eҍ �P�mۮ݅��*H]�`{ؽ��)TQ	4�D��B��@�h=@��

AA���k�p�$$-����ǋ���:A�w��6�#vj�K�m�]�*�m�Y�U�!��P�w:r[n���5ݷe�3v۶�.�ݺ6�ۦ�ݺ����T*�JKcRJSe��t�v��iT��uvٶ���;��R٪�UZ�7wm�e�e'u��i�ksW[�jn���mY����[]��b��:g[e������j���Pu�uUv�ֶmH�B�(vʓYA��c׍����.͚fSK��cQ�[)]��֨��[vs�tȗRhej�me���ݮ�8����)����U)���3X��jil��ij�[�S���R�QJ=��(k[S��Z�L�ں��k4il����5Rԁ�Ewc�3L�Z �r��U��cZ�[(�V��Th�j�U=� ZWn:�J�띈�T�W�d�UZ�� Ӷ��HV�;���6�M�Uj��ֵU��0cIP�-;k�F�li�j�25�KZ�X �D�of�d�J�����SmCA�I �MF�k+6d5kV�kj����Ѷ��v0�m������X�Z��j(�"Բ,(��	QBH�**��T�T�J�ˠd�c���X@�M��گ[�{��,j�n�+�n�:Wj��k(k56��U�L���hݎ��i�u�*��Ի �t"%��)(u�eT��{:�MSX�3F��0R���5 �)h�m��S(6�ʡ)�AA�6Sfj[5�V�LSZ����D�*���KcI�gBOl��4��붚����`�QWn�;�͊���5T��m�S���ݕ9L�[kT)4��ɢک��(dU��Jj��EW��p*
�T$���A"�%���@E? O%J�   "��I)U   PL�T�L��d�����JU   ��EU  h &����F&C ��Gf������4��1$aЕ�a��w�����ٷ<�sy���}L�ϲ��g����@$������HI��	�	�� 	� 	&D?�$$��� �c!$�d 	'�����T���)?ٟ��fjc���}�W�]�R]�Ǌ!.�u6^1Y�(F���C�p ��gݲ|��H)�cC� �5a�i'�����tvg8-V^��z�a�U��xPH�T��� ��H,�R�#N��-װ_kz"Uwr�� +4t{}Ŋq�t?;�zZїP�q�y']g ��!�ڵ��I:֌G;��g_�׌8��|�t�ֻPP���v���II�Z��RҢ�"�f��6��Y�D���-QpZ�����銂리�p�8�P�RҁP>jTMd�?W
�HQ#%v.E]'�[�B�ԻK/���B���Ӭ�`�8#X�w���?}��srN<�AH,:�H;�ɈV��t���Y�>��AH)����G��;�(m�2\��;�)Y�,��]�wr7rE�G|�<�2:��H(��5+�zé
��@�_��~�O��y�m5�rK�'��m�N�r��܋j,2�o{����}��:��7����->���?�7{���*�/NF�*�V�?��1�R����}���`�Rz(hT�U�gF{��D��8�^+	�*\�wc��*��߈�?`|+�gG�I�q)B��3P����E�KrLeͪ�\*��'됅���Ѧ5#gBE�yz�B7\����s+�.��`�Di�u-�3��ͮZ��u��r��*��vŲ�����U�B�+]�81Ӻ4�E��'F��e�_����0�UZ��0���*�U-���ǘ�QIn�֖m�Z���ǒU�Mm����5��(!���������4(Сt�	̆j���*�Ȗ��yu*�m] {(�߿A���Zҵ���D:Y���Xк��R����
�PW������eS�~sQ��a.N5���ޛ��t-�t)��39�/���?)a�1�_�d�k*c /�<���<��
e���J�K�,q�v�v���������@�C�%f���9U��M��3*E�N�^�����TY�s���y�^8�����ݙ5�!���gw;�l~�!;_�U�cϝ�_���=GU�w���T���~�?>L/���k1��m�݃��!�t���ꩣ�h��ׯ$�Z2��+���sU�թ�[��
p�b�SUX�����k�Rfsl�¸���H+����f��F��|S��
��%W�BO
C�L�ɸP+*N�!Y�P�3	�(
�H)!ԇAB�����h5���ݮ�3XDuK���n��e�.0������z(RZ�tw`�N$V�ڗ�P�ռ�a��Ū����ɾXa�k�����Y<����U٤Ո���B���"	���F(n�A��v%9���ڬ2���u�'Y/J���X-b�%y����4�J���.V��"��G[�6�؜��&��*�I<�H����Q�5.�Yı���W$£Ϣ!ajU�/����|q�s����s����}r�E�����p���i�B,����*�V(*(�G�����f�sq˕�+ǥ��`�*V_�b=U���x�</-���D�k�?W��~�����٠?fcz�^L����?Ldt��3�}��3}w�d�Ćm��^�9O9'RE�����d�n{��s̼���^ᚉPYx� ��8���r/���bs,��5'�g�!Y���xw,
{M:��jXlޭ�*��͊mW�۩�E���2��*�",E�,"�R,&���XF"�EQA�1T�3,
1Uyj�*�"��DQb��
+_�S5%�8,7Y��FŖ49�YH��54�
�8��qLWm����9�faR[)����hf`�((��[��c��ýǸێ���n�VŽCV�sn��uTj-�#-$�5���ID`�(�Q� �V
EV/�m������W����[�<�*I8�y�����i���4�D�z�BQ@^n�bB��u֋l��v�W�q�� qP�v������iT�w(�ד*��v���T��g
7@-�d\ k��w��X̙����;�h�(��nL�k��]X�_��_��fD�8����Ň&��-h�b�ڼ�4y���]��A��!�	*"�������A� �TF@U��a�S�LN��]J��,���u�&���x�z�T�AA`�"
ň���Ė0dEV"��1RUX��DEDX����0E�EdU�" (��P�F�c{h����+��B("��Ȍc5�����
,D"�b1W�
(��
(((��V"�F$QTb��Qb���0QA*0F"*��P�%H�"�DU""���TU�0Qq�,Tb���#EX
'���QU@YE"O��y��s;̢�l��+r��v�Y"	YK���Q�'��t��ʜs�My3/9/�%��i��f
��+�Fb�6��'�l�.;��-�������V݁U.��ƅvb�����鋒�ߴnd��UN��ڻ�l��q�M�5�N��7��rE��l;�J��d��!�ds�s�;�e"����#��,3�'�X��p��LÀ�y����^���\T��Kr:W!��$֛Z�j~�O\�pa��1}b��Sh+S(1w#�B="�p?^]dש�)�I-L�^��b�8!�R��^�xbђ�[�^#osUKs��2�O�a�J����i]2���ب7.Pu#Z���eѰ�9�q
ZT�23l[{���uxr6�^6��C�������6�3Y����an6��j��N�F5K�om���.Sn�ce1N�W�_�w���o�Yl���6��8��#���Ep��e�:b�4p��](�m���΄�t��}?r����o��wz�����I�����.������k�6�*��7[���v��.��x�[�Ǜ���[��R�2ѭ���#P�`=Z��c�X�K\+`T�iն%��B��lͨ��5Rʳ����z�hwM*k
�l�4m`���e�0�\zIE=��Q�(Swy�wSu?e+{�/u0Q*elAJ�WW8��3c�h�+8f5b7����������Q3-�OF�nm�
�Y0m(rf� �Z"��_�
�]`��V3���z�{�zk��=���lr���/�����HgK�R�<��eq�� 
�w7hs����:�ʔ��"��'
4)�����Rgs-9 ��g�M�9��6��d����5w���WL�w�z�5� ͙P��j�	�I=T:�I�f�閉iP��n��}�Y�b�8kl��"��ʺN�M��e+J]������jq|.�,�K�����j��=��v�SqN6��81�{�q������;y�>1�jE����+T(���⃧[27�����d���̮��܊���	�L���9�Q��oFL�T�â��.�����#CjQ�!Ԝ��]f�Y�DZ�����Q~���XG�N^���2l*&�<v]g\;��������h�x(�U�-\W���]ʚ���V�3mac��m�?1c��ē	�)����|hiK��>��7� �Z�\�<�`i[�J�/���)���� ��G�҅����De<���^6��֋���,&�ԙ�\�es1�^�InB_���?�l�J������y�t�&�7��.vV��*�u��W0���J�ZY�V5�pf���Ø���wq
nl�ĭE~�e���)�s��OE���T)l���ђRpֳ�C��u���;7\���q��/g+]�p��w���wM06�oQ��b�W���w_4�s���w~�jAH)>j�.�B���4��5�uyi��MA"��3f16\����o�B���Q��������C�y�����Qdљ�X��R̫gC��E���w4�?�۩�&�Y��)�~�4�sk�x�ک�]����5�)+�����g�1ݠ�\�ﱌ?�+�n�TE+��n�vm�1[ӸiZHn�f[�V���U2��(c�mbT-�)��* �k+c��6� 	�n��Y6t����I
v�JG^�x���d��`�.��h�zv.��1�{��I메������j�"w�e����x>>��^�<Hq'Y�-B�u+'�*ڪR����YQ(�JS{��r��۸'b�}��\IY���}e*��l+UQ-(�?��/�PG�,S�QD�DQ��J�����	Ԣ��QV�>qQ��9ywze���]�Ȳz�@�a��9���n������9���qW���f�����|�g�پ����)�u�ԇR��C�!�z�~���o��1�$1�e���'�~HjCc)b��
3��DU�R��aF#�b���� �{�{w�j��uܲu!�2�k�9�o;o-Lɺ�݂��
a	v�6����u�a�V�� �(O�w_����h�x��V�`�P+?��R�Ɗ��7Y��<�����t��N�3��r���f]��K�TN�i�Cf[8���ǷF����x� ��W�����ք��o\a$�������wR!��i=G2��lb�ˌ9w�AU\+� h����D��eNZ�#Z
�ZEr�F6�S��O�.�����0��76Iʵ�g�6m*GR!R
AH,������7���d��y��b�Eeo&�n'��_�ʄ��Wvť;�]�`�H��H5{��[8T��X:��AOv�#����jCoc���tn�4��FcO�j�O��]*p1�Ŷ�z��D�N^+�Y
eB�Rn����HP'��
��`��E��:��,�Y+v�k\x�djn�M������+ەv��o"����%�-DV��i��Ow:ȍ7�j�!�Hx��wOw�1!R:���A�X���bő���刂��۷6�.�[��aդ�?#�ⲍ��Vݰ�ګ�lX����)������2�%���6%�� ��z-	wsE��Ɉ��j�@��[cZ�q,��CdE��w[��q���B;� �GO��e��-�#*�[��cu��C�ō8kRЖ	F�8̡P䅪\�=�z�_X�̫�򒉖�ą��������8�퓩 *��?Q�f�koEm�coQ��%8�Y=Md�����;w&e!Ԃ����t��Vj,���AMN�Yn�u�LIK9[6Q�GjS��|�Ǿz�'�<�C�R�Z )R��=Hu'��m����3G9��3��OP���&xxwޛ�r�ܐ�X��S72�V��p��j=p�w�2��y�{���G��C�a�GtU�P��:��!��h�W�Z���*���E��0�l��^]���v�5�r��9�1D����S{E-�T�~u�C\ݗ0~d1LX�;��ͨ��̖�ĵH��ƭ,rf�H-�x��?_���V�kU����C8�������~��m������Im��$�%6�I��m�D��e��H��H�-4�-��`S�A�@ I/Ͷ�D2����M6 m�H���("�%�鴙E�I
$��Ci��&ZL��A6�I$���M��m�	D�$�m��M��H��m$�i$�l��i��d���Z@$�d6�(0��	��m��m�D���l�j��V��a��r�W [�x�53S�s{V��(�����ED�{��N\�J�;���8҇w����P
��H�r�P�:����Y�f_ �0�jk<�Fa�i]���
�}l���T��\��}v��]��[��`4���}�G�umL�Dc�v��i�G�*���7�Y}�&z����e�;v�,i���lJ�1��{y/ZӜˤ��[ Nu�[B�ʊ�Μ`Ȥ�ہV�M����j�Է���؍oS�{Ͱs�x�f3f��:nܵ�*�	��&4^w*������Ǖ�s�a��у���
��;�x�1��w�n�1��z�l�����ko1��qz�P.��nvJ�Z�����U�m�E��.bpuk���{}5�2��Km4/,�\����{���i��nRtv�Uۣ�,���	���q��eE����_$yM2�PNH�v�%9��o4�)���ibG���fùǝ� �Kܓ:)s�T�qWW�_n�g.U�N��K�U֮]�2��\��2�U�{�ftg-R������$`ht������x��lH�Zep�5�Hd�1_p*��ݺl�WY�4�X�Di1�ϭL��&<�n��s����m��˘R�o�����:�geh5=�!�ad�]��Pck:�+��E�+�l�;�<�ə�*&1��7)�et8��"Л��{o�Aݖ�98����.��3������NOOe}���ݺ�ʔU�K��wm�^Ѯ��mr�Wt��b(-�$�����އ�&�U��yS�t`TC+��D�uܩTML=��º��V]3X���8�l��މȤ����Fsޜ*u7��%�
�s��rr�Ѵ9�{��Zs�b�u|%�%t�qfk��-�%]�����e�}O+��.��h��u�[Db����KV��<Ç��]w�c��/.��з��y�7oC�cz�����zc��;�Ǧ���.�ֆ7j�������S���62���X0�\
��{�n���L
�j��CWn�bv_E1̻�����F,r��ṶKnu��9�Q��.�$����gu���:��/�[KJ�35�1`�7�Y�υ�N�OU��:��/)]v���N�TOM\eT�v��U������8�i}�U�ㅬ8Dy�����}y�%*��JJH��X9�����Y}�{6WT��o�hC�r�`��u5s����E�Qӳn�p�z�
�o
�3��s�����)��b�N��Ԋ�#<l3�nU�;M��7�%j���A�؀*� ��=�����k���m\ّT-ʝd�ܘ��&�[Մ�+v�{��;���#�;�¢�jSwR��m^�[��f+Et�����J�J���E�^��U��	�fv5(�C+�]d[1+�'�i�0!��obƅ��Sr�����ՅG
a-ηB�t�Ⱦ�6ڥ\XӔ������x�i<�36��'Ԁ}���S� ]�g{��B]h�Sv�+b�
��o`1����3���޹R�������.vLʖ����|�
�lbGA7ݵo��g�ܗR�k�W|��W�ԃӺ�t���m�i�!6�@��ذd�t���!�y���!�:��sh<<;�l��ON>���>���[���'>��$�[���CjM��e��"��L�!lz���J��@^�uwu��.�l�P�sR����o�s��P4�\���m�`d��{�rl�m�|�����I��f����ܧ*Χ�eG�b��4\D<�]�_`�,��N�x4���5��ei��2 f/' �549wi/k׬�OoU�ƛĭ��n�u ��l.�rV�ز���6f�YY�Q#��X�)��ƌ2�7����e�Xd0t[���� ͩ��0u�@ݔ*��s'�fZ�qY��y�Յ��e98r����H���C����X3��Y�b�������ή��%ԙ@�a�Wd u��;m��Cv��^^7}+��X5	��gT�WE���k������ QҴ2��]B���W}S�XkOt�êK���_U�[Ҭu_@M�N;��k�V�Z�.�v�t�X����q���n��*�\qtȏj)�z��U��,y��Rsg7v-~H�f�HfH�	�
8D�w��:��1�GU�g�\��dK����z�n�ZfẄ�A6����8�:�]�D�3�g�� �������:��)�	��OEu�}'&.�N�"�����ZQFuaCf���/��� �@1_1{q�v�W1�Q���Jf�,�7I"�j����.�\찐I;�2�V�~o���T��cC^�Q�0���nLd�T�,�x6�a�v�f�7t<;�l&Sg����4�?���
�SՇ5WV��'.C��&�ͣՔ՜�p�1�{�#4J+����d�z��/��vC5Qo,��:ژ�4�V@��q����WfW>�-h�K�V��0�Hm�N�/(LX�09Ȣk��zpf�'Rj�6�Cs�K8s/���]�ДP���m����r�oS4G
U��Rg;8v*q�tvjU�EZ�ԺQ�]j�_��K�y8Xtc|�I��ŝ�a5$��NĪ];ɐ�E�:aY��],gG�|.�d����W$uq7��we�%��z�]N8��!W�ʤ4�5rB6���w�ka=|��w��t�33�����9�l�7%���\�[,�퀪� o�wX�����3E�f*=o0VX��q�rH��5��z8]'H.����k�]�
0��mwY�]��k/�{ ���7����R����e|�ݼ�ܨލ�b��m8�y���}�C g{0�1����9�;l���)$u��� ��e����M<����J��esS{��M���i�zC�wm9aq��C9{�R���	�G9I��}��"Vz��*�
��O_��մ���ޓ��e��Wʤ��+����*̽E���rU���gaٙg�=9G����f�n��*����b�[h�D�noF���A^�ހ4����vM�c���Y|m��I쑧�+����vX�t`*
i�T�]���W-A�o$§ge�ߺ�z�͊r��H��!��crްN��R�1����J(�wgf�dA"�Q���t�z�vr]�]?K4[��ݗJ��v�t)L=*����$�F��N�/M��^��,��ALLK����]r��խ�`�6���*-���ʦs��q(#D�*�hV�q�yY~Wz�XA���E2���;sd��S�Kh.P�Ք�)yt�`B+O�FZ\�ы�:|mңK%��-݊�R�	R�p��9ԹLP,+v�we�N�ڸ{��SS�h��N� v�H]��\7j¿�ɨ޽�ؐ�����,��U��|���.�U)���&�-��v 
$K����ƨ~�M���V�?����"Z�
4D��$�Y@u� g�6�C)��1� T�-Kr��-ۥM�Z����n$H��P�V��Z.�A�h�x�X2��"ܿу��k�İ]�ꨫE���[H�,�/�4f+l�?Q4�rf��I���Ts�p�)Pª�*(��-��v�j"�A
�
km~:%*�~�n���,�[�	J�g���F�F�j�+i�a#	F����A�&�� �L��3f�M�����RUtL���u�+��V]x��we*�*i��X�j�a:�^�lT
��ui&��60�#�tw2]L�;��S\��vح].��]�w.�5]7�1�c�1��5���m�WB�s:�%�@�@��l6�E�QD
�%N���L]�-�L�m�[�����L��naL�w6���rsܷM�u��2��\7���0v�7E1]ݻ�i���.�k�-5�͉�n.W)]����D�
�Z�c0�̹�p��/
9�w1n�m�4�U��jfn��3Q��wW7Ki2�%�m�hi �H���V����Y�ӱ+�U%���c�*էau�خu���GN�!��(�+YƇO"���o,�*f6@S�y��?J1�ott��os�uǴ�����Q�f��Č��V2�����Y��<��i뺉����r=�&��1�믞�,�ۯ�܃y���P�Mh�ַ]ٝ�W�G�ͭP��
.�ũs%�wS{������l�HF�_iP�7:��{��)�J��8i��a�WF�Z���}��Cƚ��B�r���)l]n�v�Ek��[��hBL\(W��Ku�a� �Nm/����]����8�2t�r�#Ur��.�*c���i�3K��-�as#�A9^1(c�9�!,�m[��jV��n�+��v��T��*�'=4+olY���(�&��5ZMqƜ�sk&�v��M�Ü�g9�5�=@��X�@`/hr�*Ǘ⩥����M�rҘ��s�?A�q�Oy�}KζܦvP�z��nL1jk�x4��̄����fnm �Il��y\�Ć�2������fa�-|sx̋�8]`dg��;��M]�YP�3���M����E)���X���I�w�h4eԹ��*�mͮ���;�y��Ꮑ#�b��78%F�"�f��/خR*�n��y]v��fyI8W_C/��3��S�\-�#+7�Ғ�62��t����]�v���ݽdv�\X(��1j�{�mN����ys�wU����C˪�Pl���+�olŜ(U��xr*�\���K*�sk�-	��\8%�,^�7��:č��\���:�����v,�+��z�r��ڷRWB
`��1�פ��b�u׸;JE�ՙ�_H��nJI�\�P�p�8��]t���Y�m>�9�)Ay�呗������9V��n��qG!lC����oNmb�OUJg�ee��<�.������{�V����q���9=;��$C�3�������B����ww�b�{h	ӹq�7m�,��^`Z ��tr�K�����NT7N�U�q+)\�gK�����㏹
8"��]�g�eJ�߲+L;�4��*�<�N�v���اj�F�J
��bB�T�'Y�s#�H�c�%�Y��b��7գ�GQM�J�|^��p3r���l���z�����'�=�Ⱦ�R��R�oU��sJ��5����9�Q�/^	]ċ?��/tN�'mۂ�Q�W(�-��!^��o,!���ܵ�IԽ4"�)��@P�#X�;Pw�gasB�ʎ0����[�T�p���e�}�,i���':�0h]*�g]����ԥ&��u�n�6�Fz1tU�2�m��a;�_0��|85�����ʑ�M��0Lv�������bd��S|uʂ�(F�g5��bMԆݞ��ku|�ǐE��Վ]�6��F�ugL�陛�������9���ܟ[*g�7�Wb��%��])��6Ӥ�s8{��,]���.�縅�f�t���a�zΧZr���Җ%±��v�3Q{F-˧[W���r�X(](;Z�Mv��H�;��f���v���Q���,K1.8�K��v��d�&p���D��Ao(o2ܪtR�`�;sU�H1�+���ܑ�QEG��s�� �v���*��'��e4�ܨ)�
�̻�f�<��	+̷:�&�n.���$�m�3f<[X�E�Wss/[�s�ՄN�O[��s��ۖ�:������F��]֨MX8Y ���Js�T�oqYئ+(C�l-���y��=��t���{[n˒�ئ����]g+�%d�QhUn��,z��f�I[���[��b���G���\T�;�c*5ôVKj�oEot�o�,�^�YE�wN]v���˽�*]B�Y���nr�@���%�"�v����j���n\�e@U�O��7[ ���J�)֦��PZ�S�!N=���-�y��rf�{/���*�:�����Np6��ޜ:l�;+�j�t�t;�!\�u�mv@�G|Bz�m��Ae��s0����p�9���|[�`��G�0�2���!��G�z��n�P� É d\B�������:]˥m_ý��w�4cC+`���L��G�1�*�;�ͥVl��.Cniͨ�/:�+L7ݼM�
d�X_=G#��e���YYM�Ew]<�Đ���خ)�®�:�U7vD�o.�ˬ��{W�J���c�m�c�d2�f��+b��'IJ��7��	;UvCƀ�[O����+�D���Z��ǐ=���r�{ss����×Щ�>���,�GB%�1�z7����ͣ7�^:{L�hH�?�Sx,+$l��-��4�{t,`���4sE��'�"c)E��hE�� 뵬Z��e�}Rj���}�R�>ͥy�PD��h���6�@vAF������۲TB�U�ɲ�n�s��+���m��(%�zb����j�Ur�e�j��T�/���E_�d�C7�]u�.�Z{�_.�^����`S��j�⬮��Ϋ�b�[���[5�>hV^:h ��v��қX���p�r���%.�fc���5�5�Sh�ve��3���d��9��N�N��ZJ%���X̼s���c��@�7"YB.&����2��\;��}�.2�7���N�)w�#��w�D|��  J�� BHp'̀�;@$��!%I��HE��Ra Y 1 J2 ,^P$��	�v�!����� �H���@:��!6Є*H) (BK�!��1 ��H)$�?�!&y@��[	bH� � �l�|�ABq�P�u!�l�ya����"�e������@�j@5 ��<@���$���MIͲGϲOYd�8����B]��(!Ę��N!0B>�T��Q�偌�_2KhT�a�̘�q���e�s�I�<�@�P1̥��P�n�:����M�&��̝�M`T�5>S���2c8���u��I�R)�{�d{M;f��1��!;��
�L��d6�S��<�!]Hc#�g�d�|�E�a����,�����Q����N�&�C����ԥ��$�߬<A�0�yu�#�q�=������+�S��6��ԝf05��YZ����9��]I��>�%=�͔`|��_��O2`���1ć�)
�5!֠[CP�jaw�xÏ3܇_��$����9��g2�'2�2���
�2����Y\��2�S��'��:��"1Vj3�z��3�OSXu�SY\g�xoxM��8��ZO9g����!�o08�%q�ݥ7�r����윖3�nyù<AH啬Y�[��ML���L��2a�¾�o����3_q������C�>NaO�R]�.��z�m�ɿZ�֣^��fCk�o�;�w�8�g�����S�h`��Է�ΰ���SԜ.��p��hk�H*�l�^'\y�Ow�G��o�|��>ϳ�1���Or��n㹾Sw��Zz�����z�9C�ffq�=����Mu>��wmkY���1<��<�O>����*x���c��tr��;�3�3�k:�F)�&iq����N%�%��)ĩ�q_�h��h��1UZj�+�-]�4�J�'/��g�U;W�Bk%�u���|����N:�ۜ��b��q={㫘fg�D��(�����8���Ċ{�݋ǩǎ�����_��<���}K�5�)��u�-F+��:�_|��k�6T�(�����y�
�h��R�R����z��0����=���TR޾�y=߲j����]Y�G�z��S4WCK�����P�_��z�I���>g���1�����t��@~Y��d_����_�S���]��(e�*�fr�(Cb��T��ݳ')���q*�o���͊(�x0WPa�$����^TC�;.�ﹼ��N�����K�>�p:��S�n�N8�~��y��gl��Ȥ�d5�!��	B�t��Y�����=G�7
N�O�L�}|���w1�Vu�E�Z�|��i�x�����9O>�/�ٻH�n0��Q���ߋ�i�ǸF�����^����Hإ˼9�d��̞&#�o{��p�y�m�O\Q�y��q�gϬ�O{�6��9l��f��)�y�˔Ϲ�����5�7���a������NٞP�$~L�j���֣AS*��U���Z*�4��@C��p���X֨b��;�Xh���k1��3�x�/X.^��֊�[��4���7���� R(�����bq������N$_F����1)�.:��x���}��/<�A�������Ni�\�>��O������������+UOqr��V���1=p�:���y��-,����u���?R��
sJrr�9�T6ܹ���i��	%
�h)Ͳx��.3���Q�T�
�Sr�Q�Xb�].�1,�p�XC|�p�-k1DP�!�)���zjFXj�n��� ~��+��Z*��Ӎ����@�)���P��IУF�8�5�m��V�Y�>����0\׸�]�9�b��MW̚a}B��^^��U�����OI�,Kʭ�X(�A8��)�6�u�w2}|�q��ۊx��kZd���9g����L�
�T��+��ݶ`����pT��^4��_f�<80(yR����A��Y��P	�kQ�3 ���V?:9W��^���!�;����SK�n���z�Lƕ!�/�����.��'�j�hճa���](��R�<C���oS'9��PĨ+H p�����V4�=f���V(�0�
�2����UZN�G�!�T�^E����<Jy{{��)h)�)�i���@B��V0S�ݹ����ˌ�U��\��(�[����]n�Q6)��Ŋ$�v�2�Q���tk3�[u�R˗"����T�9 4�"�|���D��X�JV�u����J�k�a�&����I����*��9
T��bpā�L�۾W�YG��&�%ܺ�b-�f�'F�ۧ.�U��
���QxUHD���,
�\�:�f�+�-3��2p�(���W��9�}���ݳ����e�äw"�{�RU:��.���	�ɨ�� ���B�� ��䂅\�`"�qB�]������n֊r4�hx�VJ�LR��[!�'�`GYWX���ʵ��b~�:7TR�	�f��M[L` ������4ĵQ�O`��T%!ݚ�B��D�W)�� :�S5�B���MY��S3�E a�%s&b4��ҹ��$~(X��PA���w`R:�;j���HЩ���8�k)�E^�sb���H�2.��T\%`H~�-Q̛1TZ��1���5]����.�反�}����]<�㏝H��
�/!̢�%,����'�/KQ�M��i�N��Ӂ��:�07Vlc���;*E�GT&�1�-+׹LPaP�1��s�O�������{�E%ʠ�&�q��bfL����cz؎-�M��R��H�]1bj���a	r�L����� ����Γ����c�7 ޯ�5��Y�h�e����0��܁M�v��pՏl3�٘X�XK��ك7v���2�k'.)����L�wH-�ܣ�Y��T�=�٠��h���sM[�IM��PU�m9-�ݗ��Y]�*m�l��)���2��*���dG���.������y�~O\d��!9s����w�j��f@�߆B ]��!Y��V;J[ծ+��MEi�\I�=ԅL�3Q`�2���p8�ʝ��rppJ���Ǚ�\tJ�cw�іpg9`����\�.lWM���j;t�WD6�N�RK.�*��Wg^#�'l���B����C2p��B�<P�7��
[�țj�P��������MU�$a���wA�� 0]�G7I��IzMue_N8�^vZ2�7���Y�TƥBpӺ�*����|�5Û���ᱥ�mYm*8�b-km*��A�V6���c�U�]� �����+rAO�Nw����Z@�V�v��t�ov�F��_NpZ�Y����:�{q�a`J���Oo�7�`/��@	��]���Fp���b����Y0٦���#n)rXˡܲ-鰁�<����.��O����ݙ����*⡷�ʠBm���;uK�HonW�ƍjO�8}�6[��r'��fVm���9W7yk{�?���]A�-��]��B;��\�������"�q91����e�Lj);����1-2��;pާn�!e��U&�v3��=ŭ�U%�LruW����X�\]2�S2�ދ`�R(�JVX�Ļx���`��!��O׎��5gu��jP��
gh�lb8�!`Cj["�o&͵OjQj��͎h�fV�7j�ɸ�J	�EAs(T4Y���K�* ��w�VCY2)V��M�n���u5(��R����˺BGVke�Qt�iA�*HV+ijZO���D[F��^���體��r���קn�;��6��B��m���(kfq��p`4W=��3w�ӓ��с�k:�[Wk;��}��y�0^��B ����YB>t�eO�������Ӌ�q4�rޒ<��٫�M��G]I�CX�':n�d��$Àk�J�U+�;�>�7���FQu�1t���㲸sɦ:�1:V�@W^̓1��[�T'E-;2k��Z��3]ߦ���m8�N��bɻn�΄�V��9����ky�v�H�4�vnu�򹰹�"�Q� [��}"��N�Y��Z:�n݂��v6۾�K��=��j�����2!|��n�0���o+����ë{����.~*�fd�r�%@�ysv1љ[+��[�e���Yv��X-e����Ⱥ��R�<�7�^<�U�9�%.��7}zμ�\�����Y���̏�9�_w*|���S�G�����*Yh��v��A�vu8�f�w(��`׶VZ��3K�<���-�Υ�mƟg�w��}�M�8=olS��,gh9`�<ze�ʒ�,�Q{Ndf-�c��4Vz	�:�lЄ]��|��[K���E�rI��v�,v�L]����z�kd��'-,N�]�����<ܵ} ��+j"�K�E�Wdf��B��ү#���S�%��*g��vNcɝ�&T���#�Os��>�����Ɂ I����U~���r}�����gX�jֲӀ���-�Ξ�
t�rޢo�0���C�����m��F*cwz�Ie���Jroן}�c�?�I 8���0	XH��N!$Ēx���@=a!ܲ�B
�	>H�B� �$%HIYT��� VH��,���Ԅ�dX@����LIP�� }I�8�%a&��!���� @�"}������������"�V1Db��k�TF(�EAQ�X��"�UF ��S�* ��9kQDX(�QDX�"���⊢����(�(*��UUAQb��.YAPTV(�*"�2,b1b��J.Z�Eb,V=��YUDV ��ȶ�F �UR*�
�U�����[PQ?k翮vu�"
����1UX�**yB���Q���TV,AUD��IEb*"�l�DTb�(k+8�Pb,Qb���$Mh�H�2�DTQEQV0EUE��������¢���*��F �Z�Q���F,Z�&4DV(�"��T��qE��DH�DT�F1EUE����DSƊ����D_�Q��"�x��b*�b��.!DD�Tr�Ŋ�Db"3�USY�E`�"�0��E#�PEH��/��GQ"�1Pu
���j��(�1VF"�ֳ�|o>��q��xg����*���U5+X�TE��]�TDAĬQg�ـ�e�m�yKUXZ��"���<h�>��W�EUEF((�؞��(����V*��%��jTH�Db�PX֫�%�X���5+��`���PY�҃�(�PDb((�L��(���h�EG����b��0DA�,�ETAA��LQNYPx�T�%z�u�DUb���6x�1A��EF5
'樈�����b"�j�=�AY�PTE"*(�ĭc�&�{����(��UQ�UU-�"�"/��3���j��:]��a�P��i�G���F
"�q%QQ�����QUS�{�WZ�D ��PX�X�H���RU�����U�+"�\PXͥ=���X�Z�*"���i2��>�DL��( ����*�zՊ��*E�>�UTb��6�zs0�2�������b�R��p�1X��Aƪ
�����q��m{kߙ�DE\�}��{�(��$�"B>�$����.�6�����9���}s���|pQb�X���8Ԉ��b�j�
Ռu(�AEQ[�r�S����N5F5�Z��i�AJ���ED�Q��UNa���*��h�0UDDO�(�F(���?�;�A�墫�X֨��J��M���`�g�w%5���L����+*,��(f��Ag�lE���b&��;ʣb-�1�
��)v�������}�"Je�n�e�[y�U~N�G�{�����1DWԯ�?a�<�c2ɌǙ��R����֨�*�c?85���Կ���+��QQ�x��1\��,\K�ܕQ���V9}fF"�T->ݘ:�
���+W�����F|���(����Fe��"�YLj�7;���)�EE�ګ��ณ�s���
��^�k�>�C�A�@P�"����r|��G�E�B��[��ݴc�f �[jʇ9���1�T�}lQg�P�yg���_�1���lĢ;N�DG-A���mk)���Y�>���QcmS����8�X�k<��q�n苴��2���A3�s�{��t��7�7���ew�G��Q!,S~�ٔ�эo��W���s��f&EQJ����׶�~JÈ6��neMr,��4�*��ۛ�OԹ���DUQQ��+�����W,�N�+(�Z��|J�/�sI��/�I]P��\�f�ڻ~���{�s���?
{e"�Y[e��.[�sv(��2d�^�[8�}�|��ˋ`������~���Dx�,��\/p���̣�����("���aWA����wG
8|F&�\������/�~�?]
(P��$J7݊![���$��߶�LZ״�Cs�kD�`�R��S�TG~�L�~�����ܢ�jQ���r�e[6�M�fZ'���^[���i��51"4kA�6�5RJB��+|��(�r}}x:�N���8��?g���O�(�z�m%�e��W��B�+(+�ӡ��ʹ/-uvk�k��	�Kl��x5�4eY(۔ ��=���B�fu����,b� ���S�!�:2��r�!�!4�@JE �#Xg~���1���â�l��9*�/j�
��B������=F�� ��h���g����3R_`x��s
(!�����Z� �k�&\�8Q`Ķ���C����	�J��T�Zݸ��G��0}`��R�n�5sK0=a�Z����7���Te����w�}�{ў��±A�[s�S����|�o���p�'�ʖ,�o��QW�b(z���E�|��3���#Zv�9��Ǩf~�s���쓌x�W��_>�g)�6��ܙϿn�TAE11& �FҖ�1O�(,*	߲w�K�����a�+���m5���٠�u��5]��f�+��Q��Ľ�^��Qz��h�{�1�A�ryi��)�1Y��G���rł;{��PGm���8��ٞZ,7h{��*W�C/�"#mE<{�_����fF�ѧ3��X��D� @�"�Yk�*�@A�^4�D�_o��C1���ƱG�"��֪2���<��3�9<�E|�P�O~���,:�L�����8��a����&e��ז�R��T��y��sW�UD�
�Nf)����yh
�e���]:�-
���?x�@f`m��):����A�xCZ����߷�g
��H�f=�u`�,�i���~�u]J��Qzy�7��~��s�s7Jǧ�Sv�c������+Xf���Z�-jTF�"$5@~��T�'���<h���������5��ʊ��2��Ϳ�ɍ:�PX����a���c5�7�s���LH���׼�1�l�����o�^Z��Sa�w7��Fi�Ȱ�gY�G�cy�#~�79�������6�^{�k���
�
��~q�h�M¿^�E�߷;l�*Ofe�M��m"�Vm/��/m��F���n�-j>�g�^}a�^��_.?ng�}�oY��~�4�eL�40'E��/y4S�u�n��S��b�G~�-௉�ϻs��Y�UY{���|��	�(��z���es�3���M�����s�����,G�f���J�\�3X|�C��hq8�!&�4(�����/���uހ��JT���C,E�G�h���#�
u��wr���ٙ)��fx�?y�:�t��]�N}��5����������¸�?P�޴��;��~�i�!�7��J�mH���6�7;t���0<�ɩ庘�r�~�"�ز;s��jC�Li��
#��7(��}�9�s���ŋJ��/䩽��SĬ���p�*�z�忳���]�!�׮���/]��<��up�n�*榛��f˰�9��P����&��O6b�e%Z��UB�
��}���eH�KF�P+�m%����37))�\3n�)�AG���P� \������qn�"��h���ܓ�*��P~5�k�P��O�Qn?�j�x盜a�y��W��~qS]qY?w�vfC3p��%Ls {n�F����bT����>���P��0�D8kkz����a{������U��3���u+�_�7���*��j(z��X�����A
�d���D����۞|tJ��3+�q�Ұ�y���y��}�\5�B+��GE3�ݜ��}�N�OB�%�7��
P�׳Gl�>�)|�Q	`NZ/�?P���79qK��y�L�Grb�����Y7ډ�>(����Zۣ��������D��Z���[�mw��_ֲ���\���MK�0���;ֽ����!�_��7Y���L��]15>L��g���m�9ޟs�_�?76�?�Rx��UC�����pS�՝l�����RDp�4T ~���ۦ���5�f����ջ�ya�:�V& b����dD6)_<�{��5Iפ痬�H�C�J����6�޻ٴ'%;yI@~e�Q������'����3�8�E�<���~�:��ZO�M�)�Eh+6A�B�o���\E������D������>;�/�G��RfW�jޞP9��v.�C�/<��EQN^e�SZ��ߟS�wq�������0ϼ��ܥ7n��N����*a�o+>J����R��TWx̊�[u�o{��@��{�ח�=��o��5��3��+~Z�Eُ��'S?{���y͛�E��n��w��M/�َ��a�y�?p̦�3�wf�^0�̳�Y>H���]�o�9�忳|󶬫�y�H$�@�\����}P��K�+褒�C޷Du4�3��oj3�v�J!v[B7��hI!D6B*�B�UԥE/�\F�ls�U�z�Ү����.�V��(U#F��qJ�^X|�3��J}Oϻz����L_٘q��'��i���ݘȧɭ� a5Y��5�U��_����Oy*sƺ�w��Ň�m�k�t�z"�Unı��[ϔ�e
.fdn�`�	!!�]�"U�L�0��\ୢ7�4��,�8���u.���h�΃$���ᣅ��'��-���{�2�κ�9�:�Զk[�oT�����U�6[�k�v��;��^Qm�p����s��[N��S��X4�s��(��(/�z��/ɩ�6�����8S�׏8��)�k��Uqq�gϻ�x���r��b����W��=�R��\+��U���������.���\N8��j�;��x��8OZ]����R����"���P|��u>)�5��֛�˯
��rT+$fO{��x�����f�T�/�Y�3-�O�O���-5�(����G�*�;=)�O�/ʘ�PUyͭ���oEx�'��{��N�q-�[�@0�[F�$�>������8��*+���Ы�wW]�I~F�pɯ�>����Q,�8�"��/,��C�ۿ��i�{�%{\P?E���XC���y�D U�`>�Pc���v"�x·���I���]�6+�Eɻ�^�\�H��Y�}��?&���2OI�~���hq���� ��t��˿��u��Qp��]�%_�i��'v� ���3G�"ζ��UN�yˑ~� 'L���h��(�.UT���aQɰ��,���x�ᛘ�?F��2;�~�;DZ�,�Zn���,���ɳ�0~�5���?S3�&������L�U6���U��fh@�]q>��OY\̛����w������}�t1֤�lpy�<ѹs�̫��M��OG͘����yy�1�U� �f-�~�f�G�wXG�Ly�z0��GƼҧ@ r9����v����	�B�p"��>5�� 6��6���F�?vV�(��T���Mx�3ժ�o�o_2��>ԫQ$���=�
�>B�*3$R��pa P�x�jKۯ��ۼ_t��ʋU�
����a�6������B�V��ny�:��7�ُ��J���}�R΁w3.L��	V �|���"]��f�T�{Շz=׀q�#�R���d���3�Pr�mHW`T2:�*��5��8N�3�~�+��]R�)�T��Lֽ#:����۬��1����ሸ���v�D��O02�� ��!������?*G�{5Հ�>!&��,����.5Lv����~��E_���չ��`~��|����R?5��5R�H�P�*���Gz.t�0�� �lc/���Uj6o��;m_K�qy�ӟlt�P�P�D"�������҆���ƚQ�/(ۙO�D"7�JD�t�c�.H��X+oѵ���#.K*�7u�H�)k>���j:%]1:��ٝ"�����
j�h�"�:ү*&Wl�	�c��P��x~���:fM��[*�U8v勲K���?R�כ#ax;��>�;�K,�d@��y3��.&�+	���b��WJdlJ�[�_FX��EРMX�����9R����]r�.����6 f�F��-֒�p�]�T5�n.�'�1��U���(d���;�
* ����d�Z�6�Q��xy@A�z���v�{�L��h׬��y,��U@V6˺��?ơ����l�K�/�P��P�:��eX�l�v?д��Y)���{��g2�����;�U��+g&	�}n9��zB�B��Jv���(k\��U4,-z������U�&�S�Sq���N*K�	Qn��/�tO��@�5[�k�ׇ�z�.�O�c��Gj����˕JK�V�[�wu`$��.���]+<�@�n�a4 ��P#����aE��[�P��ܓ�(}A�@>��{�.�#K�f�B�5�J�َ�f2���m��(w~sG��S^���Q�\�5ϸyܮ����@�:�F�RW��߸�7��>�o��� HH��V:�$?{BLd�?$�~d�$&gs��u�@�ք`B	P���:�� 0	X@'��]��I<I�+$P Y�w>|:i�}А�Y̐�Iy��}��=�ϸ@	P�I
�@1 !Pk�@���@��\�y��@�$� �=�$��P��	���|�&J�F�Ү���Uhi6�/k;X[ƭ�"a��L�����!kkh/�m��\�w.Ѻ�җ2U�[�J��鹑���F7�ܙ�`��peJ����^�ov��ϗ��Y-��I
S�&�#��*I�v-��?��uIb*�y�j��q֣@V�X �G���K�x`����M�����r>`�:K���w��gDXbT�!]�.Z�kʢ�̽�J�/)L��2z%�_�١��/mV:>�� c���nŦ�;(k�^���}{~��P�v��f�$HM�_�m/���G<ޞj8n�:��n�"�Pk#�[�PX��H�S'�_�fWs�#i��\�p;&DX�H��T���� �Cʨ�nst/�R�A���R�N�7��Q�` "��MW�.��B&�� W��;�A�=cϭ�)��=�2m*���]�{j�Bk�י�4��|�����BF����m����R*,�5�K����S������wqc~����H��4h~8�+�`�Go�R�.�0^U
�Fu���5���L�5<�z�B��إ��(Gr�y������;�<�E�^�R[��4�q��&���t�,t����#�ON�`�@�G[�����c�
Z���^n�
#&~��<`%����~9��;ʫ�5c��a�9��-�
�I�醚4�x�\영1ή��G.S�	�,\K��U�B�/�t���Z�]����-���w0v�?3K�j��>�:�6H���zϮP�h����~i�d"�T����J�G��x	�z�\4h
��Nc*��͞�gp���(�%�q��T�Q�hq P��K9;�R��L�"�� $��j��`#��}x�0�d1CUr>F#2+	�&Ѣ�6�@)O})O=d��ר�}G}K�N��!�M7?G���gg�V~���ş}wܐ��	{pk����;y���v��;�_}N�y�Ћ#�2��BhD�� ݲ ߾�w������>W�O5̲���X(���T�R�8q��*V����a
�ʹ�iCkwy�ʢ��H�y4�C�IV��d�=�R�ӹk�eݰ`(�]*S�V�JW�"�ƽ5�k�����c,�JD:3N�b��:�o�d:�H���
�٩\�t՟=۹`a����jy�
��G�<�>��<j�F�׃�;���R����k,��a6"�3i�vj��5�����J�~�_-�������F��7)�S��*��+|�P�;�YE��Y|q���93":��OˠA� oz�T�clЌZ���k�����:��;)C�Jr�ki�H->�.��8��ܻ��-AE��
$����������O�5�.LL��b	��7�W���ȟfG3 ��9(P���< MpP�^��.����V�*&y$ t<�:�X���� k<�������xd�E׳�˓�t��?z<�h ��W2�`����Z��Lx̘R����LF��ߖm�ܪ�+'l`���Ӕ᾵�o��Y�ry�y@2P��`�a~�WZF�k�����ݣ�h鰏����S2^^�km�mme��*�Y7b�馐�r��(Q��=ks�b��!���������?�~��I����ΩD�MJ�q��n����+Պ-E��mmRL?9��33>Sw� E
ώ�N'>���l����42�j�[v�y�vz~S�Ӯ �����z�b�T%��y���7�*U�Ȋ����p:��%N^�-*�[r�oz��t�6�J�P�@�c���	����<��n4�{���z>�{(z�����ΨTE>2�㮾��X��wk0�75m.��6�$Z��q��q�ׅ#Υ��{L��*{�0�xl��|볚�y��m��tJ�(�&v�i3oP��nPl|-Ռ�=��{�3@K�Up��٠�T@5P��3��1݊��uҮ���u6��w��}���@�b�v�3��Խv��篶��H��UAq��r�xV
U�;��eۿ� �$qT�����j�A����zcjH�ِ���qV�w[��,�[x��;x'����A�RgJV�\�S�z��qDB���ٮ���__0����AhYcϷq�g�s�w�?#���#��	�#��<��H� �[�Y�o�7( �'ڐ���/|r�?ZBQ�s�A=�ك=�4�y�t���F<%����:F���?���6J�W:-�������_�n��mj�L��N�g=H����T�Im��]KJ�� H��fz��4��<��)u(�cG+���"���J ;(n�|��k���ӣsO�v�J@P������Ӭ��l�s�P�B���/�\�B�+��!·�o�6��8W r����Z/w���x{��Wwɾv%M�j�
H�����9R��ʏ�@񤏇�g�t�;5XȬ�u��̟��4�n��D>�E�9��\��G��m�~��+��S�A�ޏ��fILq~�^��'D�*�5��ȗ�fe֤�;�/�g�*�B�������~ͷ���h3cW%�{�r���
�T�N��W�� S~���^�~��|�����}��˥Q�胳� /1���<+`�ŹY@]g�ޔ���/���M��?��m�1ʝ��="�a�M���b��NPۮ�]��g������.��+�X\��;�v@�Ƈ�, ���wkbf?�j:z�\���B.��������`�D�S��*B!P�nRzu��%u��F��%Ǉ돴���7���N��ٿ�O�X���e�>2�p�{��ˆ��[���8-�1�I�<�A��ݹ�o������G0%]f�*��+����sd�VQ�S���v�_�@�p�Ϊ~��y��xk�?j�����\z+/��-]����Q�902F �SD�)/�#��ׄ������j�{�*_�l��^Uw��կ5B%�L��3$�)��F���.��}�����"�n�]m��F�
���D�6
<v�����j�7w꼯]7N���{K'�~RϺ�6�%N7PU��>�AU#L¥�o�̪70�*7�ۺ:{N+Mc�b뮩�a��u�1�����ːu?
��p����	^M����OHes6�c5^4�eȨW2f��$ ��JI���"c�r`Qc��l�1rL{��r_�(,~`ةn�]Y~l�J��R�����$|����u�d
��O�,��嚠���M:_�	SH�%D�9���N3[���n#<��J������[�GH���`cگ���8�Q�����[�%.p����v��$8�l���e���"(G�;�c�sa���:�e-DU�$�^l�	��moX}��y�zo�Ë.u������JM�g�����RIX��7��+7Db&]\��p�r0v�t�R��]*sخ�4j��(u��I[I:hN��v���ݕ8��T����+
q�ڶ�q�n�
�͈t`[r h�'��j�7JФhH�)�S��|�f�x����]ݾzTHES�,1���*�o'�ʀ�wەM����K�(�^��U�e���(��Z�J�F�"�4�o�ٌ�	sMÖE=Z�����^h����<*��i�%��}i��
�UCt�䀚W%��ܛq�� *yAL�Fgb�U�]���mbٱj�0��^�&����r�A̱w�UNKe��W�,Wj��t+�X�=mr��q�ܞ���088m�.��(ж�W��V�Y�zzC��g���/�U�D��C���#g���\l�p>1�UUc�3��r�]%
w҆z{7��p�a�K,���m(С���H�ٚ�"e��ࡡ����\5�x辱$����-�L]���W4�zù}��o��&��V+�G;��H?��g��՛��B(:pA�x�YW<�!"��i=ː��z ���D�ʞTV����zXG�*�D_%��j�8[�÷�����L�5۽��vuߦM��;e�X�P�?�ފ)|GUG/�3׷��;���K��*V����t�rzhPK�]�fߔ�Z4����s���q�R�����B#O�h׽r�c�	�Ivm��Ml�μ�*�7�	W@�O�#��uRH�����Ӡp}H�����=g�F��[�㓴2�$�曄-U;).*�!�/P@x����}�&g���.Kz�����d��������������rD��"�]8�Ee�p���T��{�w�L��ՃE��]kX�&J"��]3s�)���?�kg.�+�ޠ� �q�G�����n+��Z�g2�к�Y�J�9[�rnw,�[ge��c��\���z�)�O"��A΅��sz���W�TO��Wp�����r���f�]���FPª�5�]e���V�G�ى��q��9ws���g%Ƹ�(��WV8a�_�u7՗���8�0���hM�c4�ܦ�OiL�]�U��we������;��$J�.���n��Ο
JPWu�����	qb "�w�yei��i�592���±�Xs�Q�C��V˰�}��.�@=�D��O���I�6�(���&�y��o;b���Sj^+�V��ȳP��;��gT��+.&w�{m�X
u�����+x�\uʒ��4k.�m7 \�.��RHVڛU�r�"��7G�+��}Eڭ�a�a7& �\,%�Q�������]��	�I0�a�4)��MҤ�N�m��m�Ja6��ʝ��)=�t�#c;1�nu��e�b��&n�Ղ�9�-�Q��Vs6=;�|ץ�P�H��Z�Xa��.��Y\�9�-lܦ���yc#Q`�����"k�o�3�]��aĬrF���
��;۝�;�'I��������+x��y@X�nS���ĮЯ\�����S/�vp�/����w�Tb�s<�p�{*��{F�u��k��Z��a���M�i!�C�o5ٌ����0���\`���X>��t�N���U?sE�F����U�A�6���ee��w�jӘo)7:	oQ�%�E���Y�]W�c���B�Ɏ��ڒ#�vG���Vlm��Yd*w����Ԛ�d
�.��H*�d��ĲT5���M0�+JPȼby6ژj�m�N��<U�0��]�TD��ӻl���ٴ��4�i\ɵ�s�7JW
�4�G[��K��jd�;h��!��Lp�nrFެ�ٺ�z���\3�n�Ri5��Z����hs/(0��]t²R/wS���U26���7��Gj%��335���9ɑ���1c4��­ډ�������#�Ҵw��۹�it�����*������4�4n�e��?s��i�o4$�q�Q����"[�r�`��%�	��T4z�� �zsar͘;\�<��=�<�Ko��h;'�|$��csy�<�4,=̔�����4#���ɮ���ǻ�Ŵ��_V?��UW���nZߺO{}�虠u&]����GB9w��mR��Sz7����Yfs]�K:�<�=�)MFύ@(��G�*҉O�`���_��߆�S�>}I����u�
�����l'�d��}��V���q���0������118�S�*}���{lש�����?aX��ϓ�5�fd��.Ԝ�￹�~��W«}��K/gd*8ie����s����x�"+�3���3+E�����<�n٨x�'�f����z�xϓ��13�㎡R~q��9���,�Y�=<����0���ßfq�������c>g�13�8g��_J� MG�G�^����#�`�y|?�߽�<�5��ܼJ��
���{���B�����2N����LB�����u?&'�Ϟ>���Tr�-��C�Ǉ���4H��u�f5;����� 
�dW���#�ݿ���	�;u1Y��^{��;���E��ɛ���uMѾ���խ+]�D,��3,?�P�͡�󍮠���R;��Adq(�������Lb�|������Q?���7�j)�g���LMh����ܗ�߯��tC��5����Oyx�g������51��b��cz�b�yU�8A^��JVϗ}bK��ԝy�8���o(c�jJ�����:�L����|�����Y�f��m�ק?d8�<�$�\g��.��:߷�R�S��8�yG*�<����%q;���<O�?0�5�d�"��b�}c�ד����$��/ћϹ���S�Nmc*�?�����>S���L��u�ܥc�J��[߯���Y��]�*A|Ab%��>�QE(�Y�7����q>z������'���c_\C���:����5�g��s�	�1=O_����>5���}�v��vN��b�]
����@��c�q���4<g�ci-���Ұ��2"j^]f2V_7ۡ��)f�R�>�g�;���=���*���_쒦2��'�׉����fD�����$�d�~���x��I_�����KB��]$��3撥(�t
x�&`�[����R|�1�E���1�q��7+C�����`��ܤ�g�������E��?����$G�f���T�TaR|�r�s�M�2gtLh�}s5�*����V�9$�:�}=��n����q>�h��-��n���"3P���]a��Ԙ�R�5�M���3o�*vوn��^�����958�u+"�ԧ�r��{`c�m��y�S��<�5����g�X��Τ�f9%�[��6�'�s���q��ϫ�a����Q5Q����~�>��B*_�w�o_������{m�n�"��XW������aQq1
a_�w�ʇ�U�����\&0S�w1N5
}q�����w���l:����sy�~C�/�}���Vwl�¦&>�����@;�?���L��<�+~U�)Z�h�u��-�H��xhd咟^�k	�� ;��u6��v"P+�p�
cJ�-Z��sw�<l��ջKdTǼ{��r;��S[���)k�8��ի+��M~�V͔�wg߿S�_�ˬ����%b����m���~�!���߿���������;��׬��W)��{��Ĭ�TNfJ�r�!yx���a�̓��]f"�T���Iƈ?Y�Y�g��|C��ckԾٛ ��q�L�9�~������ z��ӓ��(%�Ğn`���8Ł���yM�PQ�	�1'���*����D�w��~���ƪ,-����1E"2����/�U�?D7q�ކ*{���_�OE�����~u�R��*(V^Y�Y��<��M��Y8�Nzo�P��\|Lg����P�����p�P��c���OS�^�6���������g��S|l�VJ���O�G��C?S���q�qۄ%2��\6#����#�@���C�Q�ɫ�Y�P���ۧOs��o����%O�f���z��1�g����&��Y�ԩ���N*V0��}���[b�R��%���7��3��I�����~�U<#�;�;�_Z C;#�t(F?�J��qyi���d3��v�3?��d�]g�L���:�m5��d�����
G�s?���1���������<N��^8�� �nDu��T1��}�����$��׉�'����x�}a�$�_:񛡯�V�{|�{�t����J��@̳3�3�C�?�O�7��������c5��N�a�q18���1����9`c9i��k���7i8�8��[�ӏT��d�ۮ�P��}����}�����1�����v"1q|��0ȏ&ȵ�dA�J0���?�>z:ʍ�L���'���Ӊ�O�M�1��>a��s�&������Ŭ�n2���.�J��C�P~�qh\�SR���疧���R���?5>��У�9��A  FD��Ձl���󛪝2gK��|����S�>�
E���P1��}x��r�o���6�����i\���>�+1�ɉ�+�� �z����?S�c
��Y����m����>�~?��S���X;���1"��h�b<
=�s'���)ʽU���<O�R����SS���=�����1��>J9w�߼�|K���e��[�a�}����ˬ���;�����\@���P�@ǍO���^fEP�2������&5<���Ͼ�UX��*�
��o1�/����
��|�q��K�rq��'��_��Ө�g��3��3X���{/�Mb����ܡ~��T5�A9}T�E�U�9 |G�GmM���I��߸8a�%jW��}�!׏P��.X|�U��E
�/�����q�ǝy��1�L%�_'ǎ�mN��gV���ao�==�����ɪ��-ƍ�}�I��9�R�@1�Lu�D��9f�"��?6��)�iN����Z&f�O�*�_n�=ۺ�=Wa�6q�v�u�y���>��<g7v�!OwO�)����2;?}�:��S��iw%�Q����_Xc���xw�|@Լ�sn�����b,�8������G��ٿ����M~g�8{���1A~uA���lG� ""mA�a���n����4/hn]h������9�d�J��3ԣ1��!�1��_��(��&%B���j]��r���2bW��繞�� ��=@֥<?���?^���1�����Y����<��{��*�}!�~�9�}�{�n[�D@�0!�ߞr���DJ�$�)��(q�CEP��1=q��]�>���ǩ��LDIZ�S��J�����x��k��U�����o�&���b<3�#�q !� �!��T�����z�7~�\h��!����!3��"��㩇�W�!�Q���ç�q�
�
��=��ݢ�W�-�����>�j����3��:x�V��!�.ϩP�VVg7t�ؿ'�1�'.�c�AC�`@��h�Pwu��[�=�+��G�>��R�� �1�C���<NN2W[�?�T��שϼ��C�?%A�p�L��7��O��K����a�8�eq't�!���b��s5���ۏ��C��n0@��H#�"0H����ȹ:��Hc��5X�)>��F��(�P/���*�=Lx�Y��Ό+Y>}7�N�E�V���l�?> m��1���SY\eC�y����'��2���MN3��
´N�g�?mԬB �>�"�H��3J|Vvf����ȤM���j>��6~O<�c���u�R�Qa���o/*Uz���X(,߳���7�,<CX_�br�&�D�៰�1�凈_م�����~ϙ�{~�ĕ�����Rr6�`��fm�D������0�b���x��9���ӾPD�n�.[3�����a�1�3�2.0�g��Ry���=ee�&}d��ĩP�������x��N����0~�a�<��n�C���|�:�����/ճ����xp0 >�>`Ɉ�	SY��8�S��l��������+���R��RS牟�*br��{��|f8�s�L_�St�^����x���Z�l��=I�و�3=YaD�dߺ��7�B$}���J$��(^;�Qx���R_������T�e2�����v��n3?��,���B������w�{��k}I�Pޞa�c��u?=�����rx�7p�?`������Ut��[�eJ� ﱍ��	�Z�%=�� ��E�煹��P�6j;�,f���(�ړ�SVwxfs��\$�����3���om�c9f����L伧��=<ҥN��Y�͹�GH�$C�B�
�TР�4�T�l!��B���<z�L0/�\�C�l��O^hk^���f~�r'�}g>����M��
�a��������bz��>۩S<�uf�����}�����~f3>�5}MgW�L��&����٩���Ӊ�XW�����ol���,�P���?{�Q���Eh���?�z�+N*]�_�{���?�E1���o��49�,?7�%�}���OmKK5���������2)��}�q:���������9:����f�DS�7SW�&e��C���ĻN%��!���5;�γ?���tD�MD) P�bj"|��c��ב�r =�Ez�\�T��x��KQ���]w*�T�߳!�;�Y�q1?�ݧ9z�C��Orq{C��̾o���%g_�|�f�]�Rb������.[�9����%K��������C�S�:���Xx����~����nݪth��C=_?p�F���C�㽤�e,5�b����q��)R�لr�&'���\OY�[�]����� .2g��99�������QOw�N<O9g��w<�7����8��n�b�����Nk���}8{��&s��磝>4>jk�B�o&�#�
QV`�r�m7�0�?���j�W��Ƴ���!�Y�Xy��j|~�L����ju��|����|��x�<gP���O������Xu�Vy�ٯ�|�@���/��<���O���O&�EuK���wC���Q� ~�Կ�h��|g���y;F�*V)ÿa��;mDq���n���5??v�G����3�9s ���|�8��:��i�yï���1^�jel����?���9�\�Cɏ�13f���Qw|յ����}W���4�~c�O�MLJ�1ǜ��q�뜿!����x��[c��g�}�Rk���3�É��M�,�b��y��Y�k�hsi�O�wj����3l�P�Y?���d8�'�q��ܦ�yW�߳���T���Ͼ�><�(5�0�#��B �jɸ� �xl��N~�4<h�~:��YzRn9(���AB �@o+���m`���Qr��V� @����<�g�+
�*A$���	t�rn3����l@  W~�=o���f:vm/	2�r��y�G~��L�#b�Л��<���i8ś�?�Ш�����Ǜ=�#���߾�J_'�Fʪ$�������_��?�< g�q׭j[A	sh#NM�������H?��=H���4������9l�4�5E3U�L˛IV��IL��r�̺����sfG��5W!\�G���ykn��|;epW�"!�G�:�osc��&�QK��x
W��Z��?=�H|�e���&*��x�~ɇE;#ID�i�7+ �Ş�5V��s�&�%Zg�[R�Q�/�?$�q4aj�����|���+,䊽�{-fe��ݥG��p��y����[֢E��/�x���O���H��Q��r��գ�ӕ��}~�H?�Tʤ)Q>�}<%�����k�O��y�����N�Yq-%���1[(X��'i q�@>Nh�$��b?�w��T�Z��*�Q'.���/�w�?�*@��*t��X#F���JP�s�t�W@��芟,Dr�W+�uۻA��Sj<E,m�;	���I�v���ؾ�F~���^nw�;������)����dđ{⇳�ǁ� h�>	&��g���S�{}���G!�d��Ge��7��+�ㅤ�{:mc�4	{�e;���a���d%ꝧU��@cn��39�t�O��U!�Ń�r�Up��,'r	�ɪ<�u�Qަ�U��K�q�آK�����\�otK�du�k 4Sφ6�&q�Xp�=�	ɺ�ti�L��޺��LAy�
pY�<�g(/���.�W�I
��k:a��H�^3>YO�t,�/�@��f��:+g�?(��z텊C{��Ix�1�ϲ�H�<4�v
x2�g�sk3�>�WMi�+��]e���]*� 7�^J}Mգ�JWݢF�Ud�]@�ۼ��t0�.��c��"�MY�2�]��q�3f�*B��zdޤ���߲�����;-���"q=B�-�{{��=�D���f�B��W��p�d���L46�k0-��ԲjW�{=dY��e�N�@9�Y��	mf��8�Ճ�g]/(ߑ�8�1`���@?����/{2ҏ%������%���Sur�X��K6�p96X������po�h~�{6]�+������k���X������B�dv��
�{b���Q��fx߮�d�[�VF�ˌ�#�N����?M�	�����q��W�s�eDx+�������^�=)'����1���ۡ�����s��ą؞�ڐ/���� �F��M�0 y�EE��_�8�,�+�y�}���Y+����ש,�n þאߵ�C�ޗr�	(/�6�].��{�6��
-䒵u%��a%P��
���[�I[�!
:��1�nU�g,�L���M��T��!W��֩m)P�z��C�-���px*��_%-�[t1�"��Qj�A�X���&��~�Y�8!QӨ�"��P}Z'ֆ���W5�p{�ÿ?��2R����ճ'���k�S��*̣Ж��^'~$G��jn��K��2I#�:ҧ�6����֓ݏ;q�����{�{�	hrIE��(Q�}�gj�:�*��Bg��}屧�*Ay!W��D/M�8�;Lt���r�l\g�Y$�d�3�Ԋ��n'�r�UNp��۸a��yKe[<�x�4�w.��y�U��a:ޖ8.[=:�
F6���/���(�	}	꙰�˞ɻ���Qb�]+ݧ�;��\�o\j��:@�}�\�}퐣�k5��j�*��@�����r��
����5\�F� \5/�;o�4��n�i%>@��@L�r-�<�P�݀|�y0�5o�(x@��F��b/Ί�z�:��+���݇{쯨�O*�rO���̲�|���4���Ɛ��(��U?H<g�C��"|ī<��7qQ��%>˨�_g�)���Y��YD`R�ȵ�����o���{�1B���%���t߰��j-�Ŀn�^�sw�ج�Ow/N� Bv���uC�&�}�eϞi;�.㓕��P_kuӇ8k���J����6k�B�2E�`T���8�!Ď[�·]�ac��ӣ����~�*�w�D�t���h7���@�k����Ȝ�}^?�^��ȍ��>��͍���k���4>�i]��Pa�ֿ3Z5�>tƃ��ߧ�#ze�7�jڅ�[O�b�����]�ۘn
e�z��QG���ך��>����1�L���t5��[f���
��7m�X�=��P\�&����-�����.�Of��W1a��<zA�A�w)�[��>��\k��?�(8��ξ��r'&�֭��������2��]�C�iP&�|�%Dx���R���f��Z����݃\��	��:��vh�����E��yQ8�����q�q4OZ�n�[�*0!��p����"+�|'F	h����D�
�LN���4����}�Mxd����pe
�)�ֆ�� �s/053i0*Q��&M�`�L+�k/x�Ï~"L��L_r]�r�rY$im<�H����� BS���l��O�O��c�?${	����z�3��W���� �.|+�*˒����&����f�m�ޚ�ˋ����GzPc|�)��r8��v���8�j[�����u�� �������])��`��p2�f�ꎲ7��f���ڃ�[C�h��T�����d�d�j��}.��8u���-�xT����=�r�򥟧�Ǚ7�R��JhK���������J��N,�x9U&d胵�o%�Qq�>e��G�YՋ~�q��d�p��D��96�e��3b�;���p�r]��З��O���W�J��a��=EQ��n�vo���hu�o�gk�Ƈ��j�b����:�S��1�����{j�D���*��C�f;Є���YYZ@��T�7�.<��������<G�KMq�8�)��ܛ�1Ɨ���o���������هDhw�Yw˯1w�ik���p��B�c+ǃe�|���Ϯs�,$}x�ϱ��6�乹�q��Wt/['��!��=F�%0H4M�qMYoޠlS��!��Y����[1�B7�+yJ�co�W����,� ���$KS�}Yo�E���u8�����_���M�!R���F3�b��y�������J��q�y��+�!Z>�����9;�/�ܠ%�zvj�g���o;�]u�x���@��+i������XO2�]�'q`�?����wy4�9�ΩO�{�N;�x*�A�ܙ�4���G*u���@�V��0���h��@p�a��\�x[��k�s�J����pn郛IN�ڥ&3�CK�ߍ�p��w�k��J���W�r~�}�͎��߾��f����0��,D�Wo�����ۭ�� !+�ڼ��rk���6Ĝr�+�/�T;�Χ��/1'>���CC���w��]s]$����d��ɍ�4N>�a@�/�R�~˪����`;��X�G�.Ǝ^�o�3Ҝ��9��!�)�L��.��*��g��MΒo�D=˿�L�E�B*D�O5�����c&`%}�E^�=��#�~_ͫ&�a���×ח�� >u#Gl"�5�د� �u<�弮��0����f��ӧ�[u�ұ�J�r_���j��Ǉ�������*#���l�Xt���kܗ����a޽dVN\m;�ڭ�cU���o���}yҨxXOlM�}5tW�L���+0��H�j��/ǜ�O�$/��Pї(��s}��'x�J�ZSW{��[��tZ�%}�畳#��h槦�Ԉ�[FB�՗Y?���7���|�ϐA%b�Wv�^VrR���͡Pc�?E������0��h�\M	Å�˯�OR��-9�����Dl@��=K���>:+���_
�7�B�um3iE�k����5�*�ܻk9��9�h���R3�gb�-{�e@/��YQa�G��H��	OJ�-��S�5v/0#�R��ag�Uսw`а_]��6�a���cw9��{�i!/ �q-����f��>!�*��������	�T���r��ÉVfA�W��Lh)�Hr{�Σʥ�@]]!93���;Lנ&&ޗޟ�f'k��C�D��������vvΩ��L��9�ïE�a����$k�\��xL��2O�۟�ջ�?I�����P8���H󼳝w�4���7�a����K���4h��u�1�h`�U���=.��|��<p�\���6�������<�>Y����W%���׵91����(���E�~=� ����!��h�.�Ș��q�R&\wv��s��	Wdҿ��XCr\��Ӵ��v�U�~SR��|r]���.�^P^;�)���n���Z�ua��y�[^��a��D��_S�5ƻ�Zu\�A����|w��*.^I�p�+֡^��	]��˜Jx��_�z��}튁�T#�6T�	����*߹�Q�Zί����:�x�k�J�I�󰤶_��z)�(�By{|�?�-xm2c:��(��>Y>�Sζ�/ �����M�Ӵ�R�5���A���*(���?��U�]��v��
OQ�pu�����x|�l�ҳ�y�'o��*�`��!��|k*�P��h}"
�^^�ӫ���_�� O�^�1��$�u���E�{�
�\�KS��+�^r�;4i�eqkm�dⳊ���A�O5aMs��j�^��?9u'S�)���lڽ���4(k��N&+8��Zf<�7�X���ѽ��6��uFe>bEBjIjV%/��+9�K������6J8�E�e;��vӕ��k��y��ub6���u2w
#�#TFǷ�7ͷF���EMȇI�n�����ZG)fK_杪(7Z��$+�β�_*T۽}0�{R��T"�sk���s4U����WXSs�ncC�@��ͻ�?۽5��F���k�5Տ*����G[u�r��[������N����F�ް��c�Nj�T�]0�|��K��=�U�\y[�����r�>6m1�Aݿ�A90�\�v�ٿ�Amİ��%�TP 3����M�淠�Ъ���\��x���� R�e._�]����%��
i��C殶P|uP"��4wS��}�.[�mZ��:v��������!�}��s��{���v�y��4]H/�����EO���NM��Q\�_7s�j<�v�S�	g�sE �w+�
���.�z�A��3��Q�*�%]��LFCu�V\�Sw����)�]\����okN���0�.zl�׮�w�;�be�`g5õ\e��5[yҷd�J��f;�X�`/�I�[�3�[Wٝu`�A�� >���.�ӷy]�?+������Km�Ph;�=�J�΄���Y:�u.�FK��k�YܶtQ��Y+=h7׈��3���nd�iej��3^��Kޑ�wWm�웖�t)d�*�B�sW{�x��gv)�]tܠ����mN!�9�r�%�5��Ĭ�Z�� �f}鲬k ��r�,=��X��5~3�)>��+��M<
K����6Mmֶݘz�j�Z1lrf+��mڏq�Ĩ
WΝ��u�F�:F�i+��� ��6�׫�m��k��]@k�x7{��fb�N�-�;W�I���Z�i�Ʒj'U��;Y����ް��{ky�y`Ʃ��K����$��g2�o�[��3�ޮL�N�/T
N9��p9I�.���5�"O�+���Vt�:v�j�a⥰]�&۫O~~f���C�5�UE�In;��wN�XҌ�/p�N\�����rKe7ǺV
�y����೼g-e�ph1cy�51mj��LE\�.���!T{~Θ��FQ�a)h�}Mgk.�V:<q�&9�pنڎ�YZ4�.*�v��*u�Yø��_�.K�W��Fk��a}�YN/�U�s{�$t����%K#ke�f�U�dOm�;;�)m�+���L��P�+��V�/��L�:�}_��U~��	};Lv��޲8a(^����f<�d+q �k[ǅ*�һ�I)��:�Л2s �]m��_�1�.��$��*�	~���x���?%����h�
�wYY�~�O��P�g����Z��# �e �7��O���l����F_��4����F�}�e��)���t��u��*~@���jc���k�^��Ec6Ʉ\K��{Z6���^q2:�L���/�v��*D.�t������Y2�?�����|�>w��ɱ��B�����[Gx�S��ڈQ����ֶҊ�=��<y���̌x��3<*�ѱ`F<nAq��zO�я�Voٿ�,-I*B����s+���?9�#��:�����(,~R��A
�Rݚ�L�d_@Aa`��S��,{�׵e��<�xyGH9Ƈ�P�ۑW�WP_3�#������o�=�<������sC� e̮z�.-4�[��	/<n���a�*����%_<��U�������\��0خe��V�Z��׆�S4q�����A	Ly8h6^f烖y\��B�W0�Yܻe�\PzT����������D��F��P#O�*��+�c�]��u������Sy�
���O�h�o��#��%�^��~E$i#��A���L��a	�����s�=��������g�pv"�- )�A��0(W��sb�G^�uw��q���h�����ގ��J��H�V���ؚlɼ�6F�)�����Qҡ�}XBv^=�,ItH~ѲN�ה�s8�BI6�4�%%M K��]�S�T�Cih�Ԁ�aA
]3
�v��sv�k����U[��+W�QS��|79*Ϗ�E_z��O�=KG2�<?v[�;r_A�U~���҉����>=bU���q�̡M�����(O�v%_
Ұ��t6��oQ�U�*9��8̲�$Cb�_��c�|�QԖ��\���K�ڣL��t�o�Z���kE���::��K�Kƞ�g�KC/wM���D�<'+R��`�Y�{�r����U�P��/l���$ϡ�Vf�}i����O�C��8'� ���������g4竝�#;����jy;�~4&$>��E��^�>
�$PƝ�Kk4_-��Ux�~� ��C'�y(�����K�(_`��j�4����"�W��2�
��k��:�|,2�{w0�D����WO!=X�dԥn�Lf���<�ʆ3����1��W���qQd�P�	��vpغ�(}��I�������XŲMI�;;ܭ>�P�F�8ϡ`�}�pm���3]���7��u]����<M���	���~��j>���=�M.*�=�����`_ڴVᬆ��dp�ø�3�j|�u��q-mFWH�������Y�Vz|=��#]9W��֞:�9���������|i�Se�?�D���T�ח|i22�ϛ�����9e�^!��W��Oy�B; Oo�ܭ'rLZa?�](Y�gf/p/or� ���+0�/�����Y���9�̺��<�r �s/L} ���s���o+:q���q^ӓ��,�8�P`�'ns�{Vξ}�:�C����.�|��M�zS��?�V�������j�����d����D~�������Wk"������7o��ڀW[T�Vm�>^�"�[竪h푊\y����?]*���h���ʄ&k�!�r��]�^�yn��;-9S��$o�w�zK��cY^:����Jb�i?~�W��[�͊>���]�3�鳜��/.٢vj)F�a���g���wb\�w�feO�h+/Ǵ��<K�U����&��w�����c�#�/�d� �+��};6��߮����|�����y��߼��m�z��U��*	�+�z�=)^I��J��v}uyЭL/
$Qݛ2���*祎�M+eF*��^��ΩЧ޼�E��w��(
ĳ�>|���P�F�皁�����-�������\��H�c__szC}>�8́��\[l�I�ҬD��ia��(*��(3���>]:cg���kjΊ�(�(W��9K��;���>�b�1u�`e�d�J�Ǫ4���t"��h�s�����.�@��8��"�I%�Ə����)(�ݦ�ߙ���"��DʄѭLN�r�տ�x5��
�P?��u7?�,��y�1i-ܭ���BWqkF�nK��������\W3d�82f��G��Eukm�����[1�}���%$��9e���X�a���j��8����[��}�2/C�dX���}��V��l]͎��(���X#�{l�/�]	��![C�K�p�ן�o���`�r+̙�������F5za}��w��='|�X�_��y�Eug��@�Q�G���<{Ӵ��r��(�}�{��_��)_��l<�#�M�fX�h���Z�Y31	RD<�|I348P�XKg�x{�U?pk�Bv	fv�>A�^�o2�Qh*U�ᆉ�U���j,Ѡ�rK7���}U®m#v����C�.�b�%燒3�;�Կ�{w�R�S�௎��;�K
���l|G���ާ�Q��'&.jăQ�J����ٰ,���"ƽ�6L�eۺ���>�5�$���5�&�OZ� �*��:N?��O��d�p�Ŗ{�U��x��%�%��_� 	�r�#��
dT��W�Qױ=�+:䓙鍳��v7��=kr9w�t�~S4M�����L�:h6[����u[=@�G�\>�<i{�� 3�����]�:�0�?��*[��o�}n�Z7p=�+͸"�C_�U��7ϲg������(�����O[�`��?h��߰���E�����U�8�=�О�t�3b�p���;��O���e<�³@6ǥ����ߵ`�dY���j�o���~9�r�^t���gu������*l��L���]���7��oj���mE�(��5&\�d0Vl��k�J�yu�Sz�vp%�-ɸ�7���]��έT�q�~��x��7�<����Q���m,�$!�W\[�wq9Vy����
G�w�u���D����Hy�G�n�%6��Gx}$�����=�Oû-�U&IRO���~S5�_����e�r����3rd��Y��vZyB�N�]}"8vA���Ւ#���+!���N�z�
������I3�oim�{���d��B̓���Pc����0���^Ϭ�g�p�Pfr�]g��+%\{�ޝ�M)_��`,Zs��'n�$r���N�Z�b�hEP�1��f�����G�3��l�)c��y'��ΜW�������'�7��2�F\z�#@�c�fϪ�T�^�ꂄ�����Wt��xP�H֨�Pu�{�EŠX�$�H���ױr&��s���{��� �N���<q������/L"|h�x���B�����d(�M�2�Rk�{/(Wъm��fxͺeݧ�_׿{͓��N�5_L�P��S~fw̰����G>G#dݟ���sC��1뻞����T�r��9���@���!&�03��Gt���WH��{&�(O��i�ee=\�d��t�=���H�� b�X-�C�(hS w�i:%o;�U$�1��2K�5��L�3�7�a�e�C�n�za;a�h��+�Ӄ�Yf(^n����vsYYu`�J�<�s7[㏖j��\�����[�%�I�Ot��w%K�3z�hw�C���ec�eo�y^�?,�7l��D���T ��V�3�r
%�R�'�n�-��p��:��YGm�TP�k���}�r���c�;��J������,P��s���.z݀<Jً��N�g�%
*�y\��5ٙ�? w���=]wL�Q��|�=[>�[ѹ(����]�lƀ���ؤ*��M0Q.��Ȯ��2L[Mt�хg�<�G���ə�C�4�i^F��q#�j�ɶ�ƫ��|o�x��d���G�5��Р9��\�����+4�}��D�g]
��ЕD���� mâT�$U-�H�>��\�.*�[>�B������b?�^��2�-�� ��}4P���~�V���ѥj���`9������¾R;"`y������'��K�F��һ�������,1��i,��W�X�1�a�חdG�B�Y�¶�,ϱh�)Oi#Ur�ެ���-9Z~��Qkg��'��h<;��޼����答�����~��T	��mB����Wt��o������N�2(�myzP�A�S�ø+��q����$2�N?Iz2�獌bG2�lDw7>~�v����fn0O�]y�<��Ƃ�F
z�Ll��xE@T��7w���^��
�I[�T��͉M\ЊC��uw��Ok�d�>����p�+�ݺ���{�M�86P�����Η��H.v��p�Q��-{+�N۩�/7�d��{�-u��LvL��g�[:��D�6)u�*�15tR��WV�.U]�x�Iؠ��Üe١�ۺ��\��k;��!���r��U	jn�/o�=v��j���e��pW�W�Э�%��hU�0�Z�^H9}�n��|x-�l�-}Ƽ~_ig��������]�cϙ���p��yw\�̬�H��
�~�	@�s$�_"ԊO������r�_:���嚽̠|���'3鵛��yQ�| s�����ڿ\J�Y�y�FDP��W��u[9�6��I�;��|uv��ɴe]u��*��)��}�I��Ւ�u�x��~d��}�`b3��{�t��H~/
�򯘣]C��,�S�g��;�*2�X���O�T�{�O��Kw�o��8{6u��3_��X���0��#r���FS����,�U�����'�RK��>�� �Hu��A��{i�8a�ћs��׺c��;O����7L���T_	H2�׎,�x%��{=�]y?��0l<&��$���u�h,�y#�'[4g�)���`�9I;mP�4}��s��]W|}�	�wq��F{գp�|���ۘ�<�rݷW�*>��%˲v[��kOf�y�{bj2GGn�h�t��e�I�<$f�Z;+���k֜��򻿓�m�v]�ˮ�4۫��cq�PD�c��-z�ع�W�]�.`~��O\o��~��a����#@V��1�f9\e���T�ܻH��gz����琱˻";�jJ���qЦy,T\�L��E�cɛǻ��U�)��h�X�������7w�P�S���D��{1\F����tD�f_;�;��cSv�%vX��W*H�K�w]��s��\e��UOH$F���B=Ģ*tWNrN{j�S�s/��	n�D��v��)$��ٰ�ʢ@�d/*oޭ&��j�D���Li��;��g:�:S�uP�����|�K����fEC�}y�T�IɡQ&5S,�T�N�	Lhb�Gr�pV��̵E��6A�>	�}9�x��S���PW�ٽH,��hQ�Q?w���$dd�j؛�y��`uK�$6xp�b-{;�Om�f1�hC.	��o�|}�k���������4��`�+1��hRk���>;��W� ~b�0�[>Mm:�����	ݲ~�>5���|+υp�y�}Z��5
�x���cOD�(0�?f����I�x�W�f�9>�9����ɇ������ �*,��cYy�m�H�Y��|�����>S�Ζ��|����o��*����P�n���Z�������5�#���x:�F�b����\N��^�><gB���z!�r�z�%�}�-�w���Z����^����ӥuc�d ��l���?X�ze��o������A3	��L=3�ͺ��քuHPu��o�E:�7n��$���N�i~jzt��5y��_Y�_OI���bxw�V{�����L�j�Wu ɗJ����3e�����6�oiG`��K^:���[$URU�+3Vڄr�c�X3�!ӧd^։�f@�G�.�٭�@,�}��uՐ�9�q��5���4K��9 ��3�5UϦw=��Ь���(8�����,+*���
�b�vO�"H6��x��u��!ÜF�V�)T��^���V��Y������E��R�^�+E�KM��|�I�Wڻ2�͍]|%�[FT�2|絻�����e��|g���~^���lUxu���)�&���G��5��L~��g-J�{gk%��c�NFy,�uR�ϊ�3���C�T>�_��O�_�%�h:����e�~U���6w��i�*,�+�����9�W6�?��y�)|���^p�&7�[���k3m%&�ޙ|���x�!��k�h����O�@�����Ta>���$��S��}�{� ��:Q���≦#��~�m6+7v���⌿����a
�/Q�߆?e�"�wj���X�u�����V;~�ΰ}����~���6�n��T����+au��#�����Ļi-vz�+6����"DF/D�������^�5_y�O���둲�C/Hq�|`C7�X�}_fG�Xy��L��O���7.�Z�����'$�jXl���t_�I��d�h�;�]�W߸b����O�v(���
�>/,[��a�iuC�u;�%����O�n�SfQ�F�-%CF�qԖ��0���K�J��h�蓼����;y��6)ź{S���b=cv�8��"��
�Y(�۴�5 ��eӤv�d�l���������Zn���{B���x�o\6t��c7%�<P� ��Vm9��ۗ��8F_����f���DHE+���i�%�}+��ϿN�kK�R�x|+Q����b��Q91< �z�L��<�xuu9�tvS��o�բ`qBs\�߳��!������~u�I7a�f�Kk}�F�d8�g쮝�{v�Hꉎ�Jw0�1	��瑱���5XHK~H�����@N�u�(�~��I6�"��ᴵ����.A䆟���*�tήQ��iӺo||��l�ֱ�Ѱ6U�f�kR�`�����r-p?qB�?�}���p��V����KÈI���Ugު&��t<yq�;ݒ����j���r3P�Q9��J��׵����R��&�w]�f=S�&`��׹�1 )��oڠ���5�[��!}3dױ�ϭY��SZ���
�g[��P8�|{�}I�4�ְ�_CZ�X�����7����E?��n�*�i���=��I[�yMګ��F��^�{��c�HE�I�J;9vZwY��lW��G����fq�{��oTz�4��$�d!��6ܿX�3.�l�}Y9U�q\�~�<lK�ZVtƊDGm��By;���R^݇��1��~9�-'N5��)�J��3�&_\Y�T�6��,n�;&۲�ѡ�j>���/A3�jBb]�ن��n[S���w���v������V�3y�.l���f�z���%��/V�\O��j�1w�2G�adI;f諭�?�Do�ݖn��=���6W*~���-�.�%l���o1���9�W5�-;�L��LG?]Z& m��wCp͕����wm������n!��st;�B���f�dj͗{X�2q0�g,U�l'��/(ؖr�5�S��q5c8�t�5z���n�˾(�em�+}������^^�wVVo�տ��^0�c9 �K�Z���"�Cˤ��):���X���_�%u�I�q^�ֶ��W15]�Y��K�?�-<����MQ�T+M��k���9����k̷t&(�d��.��eЮ����(� d�^�4|5b0��Rp���hr+�OlXۧ;��-��j��y�y��&w��:�P˷F�������z��jN|D��[����
T'����j��n���jW����kڱ%4�m$�K.�
������r�!u]��20�¨��=.�R�+�|�ܻ�e��/�o���j�D��YU��d��k�),��&/����n�՜h.d@;�Ф�oq9�oW~�hsa�V�n(�IeTeY�C��&ek�勚��J��u���5����B�b䦹�h����^�������6�Rs�E��]7�+����u9�r���oi��E�r����^����n:��-��bYÎs�K��gm���j�>���D�&�K��,�����Ś�hӠ)��E²#dQTN+{1`=6��(+�r�M�Zx��p��k榅�>�R��um�g㠳��` g��,jv���Vqn+�Z'�U�Li?݉ѩ����7/�D���ю�9]N�2�6�_�A��(1�'4�f9�7vbC+9�䧔Y9�MG�R�<�tYz��E���y�������
.�%�lj��q��[9W�0�лys���}�n���T�t(T�b���f�Y���@���7�:���Ț$�vA�{��ͮg0�5���cWo:ĕ��fm�t�y��f�OTkR�g�t��
�zc�-li��(�j���b�,v�I3�4�%��I���K:-�k�����i���]�m�j��m&��<�L?�(QpQZ
Z$�T�� 4��Ih��'b��@�Ҫ��M�f��R�i��i�׆mi��n����T��7��6[s-����.4˂e�0e��1��֮�a��:K��Wv�Q�Ld���fVH�	eˢ����oE�z��G�ץ�!]]d��#��J|k(e��YwYڊ���Oz��9�&�T��!���%���.h�V��μO(��ǖ].�W{����)�fN=V���Chu]�}�@�q�Z$޼5�Xsa�9Md�[���ǲ�Fd��z8�I�C𮵭])|��ŷʯE'/���Di�{B��N����f�Pjɖ����XW�+�]ڏ��%l�])��L�̼^��8��O[��}4����$�9�/���h
��_/e�p�%_wmu���]��%�r��Ww�1+��n5���;'*��N㴺RbQ�ܰ������M�Ɲ�L�3Z����Ԅ_�V��щ+|�Å_|-h�����(��cnWd�gM��*�s��s�)R��8k98���]�s��G���Z'�'�Qq�rfB��?[)J�)��幢�_O�& �8Y..@+�(��Qӎ�{���0��Zr}q�L���ܼ��܎�vK��5��g�$b�����	�U=WC�g�<["�}3~j�=����n]r�u��ߗ�o�������N�+X�c��쿲������vEQe���&<#�VS�7�AD	e��1�ή�h���#2��ծh}�ͨ;�w�mm�~����b�_!(���z[��C3<́�����Ag�>��8�m�2�C}���#�a4<K�{�������η%B��g]o�K��� �y�^��c�h��^�U^7�9u���r�$�K�~\�z��Lo���mW�G����K���lT0O�v�?��@Er��G��B�J��������?5�,E3A���Ǿ�j-V����!h��_+W_jn~�;��T櫖�>սh�^�F��*�?�m��.e�����E�^X�930���'�w/~@mW�_I�%v'Nb�V]o���t��4�$���mw*%W���*��{��:���$\��=�ٛ�^S"�[
ol�m���8�*䘘��/c����z�۝�=���ܢ�U]X /dH^��^�.�%��T&�[<�W���L��X��j��i[I�O��������	qЂ�F���d���7Lx�W�<�������/{aR����X��t��˵KNc��Z��tp���ދ�T�|�
ZI���q�Z�\6�ߒ�m*��L��ֈټ�eʟT��V{���Լ9j��J��k�|ӯ���`�^{v�u��o�I۟�N��\+�6�O�}q�s�V<�t��g������]�2�|q�șq�N��}jl��%�^V��Q15��`݁��ެ/�?�;�����z�����˱7�u���j��qC��6��ǲ��+�("W�-��B��5�����/�,nm���Y-�� �3��	A��φ��T����<=���(&�h��-e��eP��ɟQ�-S��ב��c�0�ȋS��o��W�/U�Q��}$x �W>l��� ��c�2>K�1��Lc�R�KǇ=�'�ok~%�Vx��l+���Os� AΝ�u�n�H�\��/}U�,������@|{۷��U������������������.����ה=J�
�W{H�.gr,I믮�V��j=�\4)�c]BS_��,U{�7�Qw-�u�������f�Pa�H���WOV�~�V%Tz�塎a�*��q�
�=���^�w)�]^R��^��e�r��\��$鎬��޶9�n�Ž��P�q;Y6��F��>6�j}2�TLh�:��9<���9�K�-��2���� Z�RF���]���Տ�)&�> /"l��5=�=�vRcj� (zOT����̹�'n�u�ފ����4�K�;#��\Dvc����g-��J���Z��~F(1�yL���QmeG��sM�y^<�|id����(��f�}��,'5 <Y�S�}_.Ҋ|^�m��k�|D����<Cn��fŌ\�>��2G�cw�Rb�G@�C�����xB�_/[��J;"�e�-4��}�!uf]���E�ۦ�F���oǙ����__Y�}I�S�f���~5��)Ty�K�i�;���i+c�c�'RM?�s�����ǹO��&$�I���(�GCA��t6���N�S�ӑ����e/x`��O/w�;��M'�x=+&�&C�Q�����<8����S���׭������h?;� V�N�*9rS{�Xzg��}�0��`�$���s�!��0p��	�S�y9����j��֘w&hS�u�{v&��b'��R:�N�A���x�8A����tN�]`8�_��>{�ך�ש���=�n)�;L�A�8�5^u�ɒ7r��Q���]lc��6�\�N���`s+���a�^@�d�N�Y�{��O���SQb�<�F�X����C��2�l1����#�`�B�L�A)$�-��n���ك���we�tN�;a���U$�f��J]��V��>eO0�
������k:0/���0!���;���<r�ݶ�}@b�TMl�C���&�4D�ͯ��g¾��WbP�G�^��s�)�:�=���{/��9J�,�L�R�;�
6�`���\##W��4H00h�@x��ﾇZ3����:nH�m�}��f��Ó�BEYa#y���׷םf���&���8<H�w�Z�=8Qy��j����-��y�R���t���t_Sw��aq��=?G�9܊�T8�I��#`�sW�.�v�ǽٔp��!M-/~��uMW)���˾�6�9�T��F�.5rAz�/�����^m���������J�iC�lR����4���6��J~J
�����f��ea�>s�Q;�{���U`��'���wyt:��쨇�@���j����@<q�Ԍ3zV��[��3�����7E@}�����sRa���O�8y��P�/:K`�<�0߽��ܟZ�^��V]]���'��]����_�V\���.�c�2�ڝs�W�*����'����ɒ�x��o�c9�ᙸˑ>�:;9�Ȍ��饝#Z�&'��1�\�/J�[[��,ɚ`L���O��?��s%w��4n��v���?{�0�r�e�c�Z{26c��*��{����@&���a�4sC�&s�ܳz�x�?!U��[�����Du�m���� ���V!�����Q|��(Gb�N���5�P4���:�b�������k���{I$�0�52������:�*�|r_ŭJoѥ���c�C�-K�'m��z(Q��Н^_u]��K&��؞�EW�`\f;��^��'��o�m�߼� F���ƕ��Gnv�x�,-����o�����y�'���ot�9�+�k���q�S^�Q�1"��׫.R�IEB}g2�nz�T��b��c�L{T��Ѯ�F���3n��6^����|}L�N���.ߑă��h��3��ڧ4�t�=.�n������l������9�Ҳ6L������yۅ;���t!#����Dq��0��z� P�lh�_ޑ�������3��zqSc9���5Z���oZB;v+�B=ͅ��pSOL�ʫ���8���t&e��t{g�b�~�ԊB>����Η��z&��*�0W��8I�g�eH4{��+�め��ԇ��*�ߺ���
;�Uc>�+@6�^�%* ��~�V���d��VqS��6��e�f ti����s�Z�Uʈ""r���e���|�k��]�����w���2�_�L�x.y�6�(P=|�M�}�ܮ��'�£mj�Եued�PWTW���q�n��|��1ѭT��'�3���V���*k��bu ��uP��rl�U�2���Do*o<�]�s�AZ�Q�u&�F�HS'4=��v��tH1�G>5d�[}
U���V�<�ʊ�X������5:�H=#���N�-���I��X�2'����w\�$ u2p��]�5܉ҏ����-�/g.rulM���x,41�|0�3���/@����BY�h�9��_^�Y�:�>s�.K-L���~�bH*#�����X5�F��&�.��4;iVcG~x�C�H>����W��wQ`�{ �B��(���|+<��IJYVP!��3�C;dIZ��.Z���w�.7O���)y�x� �d�2��y148MHn�L�T|�FI�;�Wէq�;�z�4'���N��o�FJ��O�iv*��PB��%j����5o��x�2>�-e(�S��˓7�{������q>XܧK��ݣ{�����ǔD�}�}����X�鑄p'_�Q����C��������_bT��X��[>�q�s�5��񛠉 z�۲��1�!\�j�,#�$��>��L`��
y J#;���߭��泵�%�q~_Z�E��>�[��jq�!��|�m����3�^��7��?��t#�G��cT�O:j�v&�(=�w2��=�bf�r��0#j���ᗙ����@�g9N@�c�hWdSz{��q��/(��i�\���S���U: ͜w$�Gd�!|��ywB��T����\��/1@�lh��N�Wg	2���R\��?�v���ƏY��3�^ǈdNN�NT��|6���@_��V��v� �e��S.`�}]� ZRF��������hZUY�2]K����m���V�������vc�tԷSŜ�)ֻ,�?�c�Xk�b��̱��O�{��-��x��y�ݓx�f��p ��������ѷ��V���H\6O��?<��	��a�:��2�e�V�i�I/�����26���(!���u��t�}����5���RZ�G��}�E�>�B���+޻s�h�Z�HY�}�䗚�G�����E�W�2�	jû��N6����Of<�l-\�g;���n{$�_�ؒ�C�Z��`�}q��Te��b����s�!�w���<���Y;K��9�Zg/1?S ��0ɰ��6 >�r���R߉F��02V��:H{��z`�q\
<2C�ɑCPS8#6|9�z@��bCY�}�|���C���EI�Ch�#��]>�8�O����}���7��T�������{����>>�Qy:�*|f�`��W�B��m���	���U�[0�nxz��3.��=S.���Ro���cT��NX{�^���tF=�v�h)�d��fm�O��c]͘�f���v]�ᣤK�̌�'S�1Q����:��VdR�s�5⃰��,D�*T�o�Spt˓f�6�]�ݛ��7�ޜ����]��%h^�Q����ޖ�O���p�4�]
��O^����On*X�N��&N���2 ��K]���%_��Y�J��x<܆n���~���$	3Z��yU!�w���e��H�D�ᒽ;)��#$��ޯ�z\u3{4{{\�9�q�ҧg<>;����F�2�uy{Q����':wS�{X� �c�tJ�Hzo��k;v�^=��*>^��aw�پ|��?f�ߞ޾q���z�T�9�I�:��f�{��W.��t�w�'���J7��{��!���<�Z�}��=�L�}�O��Ϸ�4�>ߵ�}����������~�����J_�/�ƕ���,��٥�|6Q���g̭Ǫ?�u�G�OK�e;����p�ލ����P�i���=ښʬ%Ӳ�d�'}QQJ8����Tu�wl�>�����@g�/�1ea_��P��D�v�:�ʮ�:<�zWg�g�ʭ���	���:2����w{'��c�G�&os�H1.lM�ޖ��'�]G;�Ua�<�H�n�N��U��^;A�iV�?�x�-��D�?n�z��XV���}�]���mcy�E$M7\m	o�֪�<4�n>���~�Y;xw��֮m�S�	f�,��t�F�iW,8��{]D�)m�-�W�`��.�����YӗUzU���_�+�j_Z�.�9�B�՟J�<Zy�s���3�j�rM�Ծ������{������<����7�Ev�|�o"⪴��ĔR�U�U��xڹg�dO�*z[헑?P=寧��r�-u�]s��.�"u�Ɨ��皏l3]z����-O��`�_U��������V�=�Wp�E��^���ݳq�Q���Wza��7}�{~oPǾ�G������:��:�J�^��UV	!KK�D��P�.�|�;�Q�o�z��<p�D��F���R^K��{�;�}�;Em�0�]	ri�ca������a�F����g�mF�.�+q�ύ���,��#�vT37T��+�E�ƽJT{�រ�8��ƥ�)?F�=dc���b뽂�z~���˳�����"�o�����X�Y�%�p.jf��/�[�0&���}U���l㊱Mf��]�T�S��{�m�]�:C��]�mEL����'�M���it:�5.W:�wf����{����%�Ew*;�7��Eީ�����:V�ө˩K���qӓ.!��;�sq��uL�m��!����۠��by.̨��zԻ�}�>�sa��۷6��yO|�=�W\��~ϫ��������~���󫫱^��=�W�1����D����y���+��-��]�8;����>�b��rxcy^�M�rw_3V�3�#����-��<�R���	��.����3ַ~�a��o��%8lVT��ڼ�ҳsdD]�m�z�cB��"i���57[��U�A�	=3����Y�.�/��ǜ11�詣^��ӆS;w�#���37��Ŗ���3�x���֎EF�vn�gr�}�d_�����+�FQ#�
��?U.ʞq]����rݷ n�<� �������iz��Naz�9�*��*X�F;S�"�w�&��>�s�1�'��T5��iF穀m[aq���T�W���S����|�ϯ�
�ּ�Z�k��Ǻ벦;���"h�=��W/�-�n*��������G�x/����Jz<}�C1Ѩ��v�u�@2�Ki�����ұ�r"�t;P�b�
�nԭ��Q��S���LTCMT�[���:{bV*��=R�;ޭ��{�O�Y���!�ڷ���&Ә-&�c�nF��@-kx��!=�u��Y���\����L:ˇ�3D䭥�J�k�����3�ڕ}{�$(�j�2��u|����z��޽Ͱ.W.��)�ԛ %��Y��/Z��ڍ��l��wu�dF���r�r�!��,J]�GC�6����)��k�?���+N�b�=���-�o�mv�
 �e���rO�;�x��<<�k	��U3r�٘G8��Ӯ�go�+ԣ���2 �Wɠ�TI�ETՎ�{W�ћ����8iX�.�i[Q��7�ɹi�=�I���5��ggn[�����=sig'���s(LE�ݏ��;��9O��}�Nt�M�TL"��j����
�qn��I���&��E�:\w��d�۫�fV;dA�P��o@(5����jD��쒪�\q1�{!G{)\oQ�*ƈ��-�	��p�.���͌��1aJ��u.�xh%�c��՚��s�bW{wm�O�΍��P�#��O8�f�sy]r���Y͋w�b�_k}F>=L5�vM�w8v.r�0��E�;"����d2��X�H�na[�4mc���.`���V�9�4Żn��̉��vFR^՜��ݕ���խ�*[&���L̀����ں�lQf�p	�\ʕ�]���6s]�i�dȭwi�yLm��+};�.ө�u����.��.��+y'K1�*�Z�k\5��e䮊P�6�cU����:|���͙&ޒ����lt:��]���Ev]#k;���A#��Tw���bCH�_j�|m�Em�Gn���ԗ9���������� �g<Ƿ��J7�g9t�xdx��8��\�BP}Q�ZkI���uٸ�d券�c�,j��C�-���Uǜ�K�~��4*؝�]̛�;=VWH��;�2ۄ���u��t�ݖ!��u�|If��P!��r���ٮ�[-��C��m�D�@����M���Ϳҥ�D�Z큫볚OR��/�c�	��<�ӽa�۬�nu��u�ΗW[a{�e21E��=eɮ��w�'>�aW;q�)vq ��I,�h��=/2�ٙn�rx�B��,��*�lp��L��6a��1�û���Y�M@P����
�E����n,6-	�hu �$p�Cx��q��W7\�����\��'7x�
̘!���d���.��w�4���6:i����e9��3��~���|&Z�g�pk�^ ��5�m��\y8����el\{�����ݭ�����w��Y�[:�����d��4�=��y܅�\:붳�ǌ�нQ�>��d.�wi���z}k}�z�w�[��W�Y���}۞NM\W壘�*oj���ۯ��6�#��.�^��<w�t'��vg���&�L������जG0��Y���an{㒰��x��Z�2;����^�аM���fk�Vk��u���8%���z�ض������oz��v�<m�p�G��U��s7�Tz�t��ӭ����+��Y>PCZO[G-.��j�5���.u7��X�T)�M��9�3����D>0}���)4֥s�]�}I��	���׳h�ԡ�GS4	�\�ϳ�|H��|+@2��H������l~P���]����ϩ���K�t:�>��Ǿ�Hv���S�t{�싱Fj��Ր�o{��m��nT� � �h(�	�V�c� �_����]ޮ�f�u�Bf��G�A�3	�Ǿ@��W��C}F8z2�Ç��(�����-j���y��n��-�*ʙ�Am���0N�׼R:����c%M�L�k8	ZO����wX�v����Oݧ���3*�\���`����Dp�$ 'L�ʤ�j��T���:n� �m�#������8�û{ ��Ӝ��l�&N�k�^1'��i^9@���a�|WO�]��m�����Ρ^��6�ë�+�V=���J=s�X��#i�7�!g�[�|]xm]�31����zٿ%�bg�r�v.���+�l���Y3�>	C��6�4����7�"�?Zג��~������Ty�G:v��Ǻ�m�<US�C�mϨ�7Vq����\ʷ4��wVW|{��T5}y�zL*C[{旟~=���ً̻��2�վ�@��v%tEvw�j�Q�Fbf��sZ�wW���o��Lg=��%�]�G���&�3�gq���y|uVolan�;���L�γ�s���p=�<����][e����ϱ��e��f����:|����'ޚ/��KI%���彟_s�W\��>տ_w��3���3�}p���]槺��O���βՍ���Fh��{�fP*�ӬC�Ǆ���_Q��Q�;�_J����=x��9�j�V�u���-�8�B��z���v�Ь��lK�xҤn�v��+t.�`�Q�[���jwJ��c��fv��C��N=�sgxg(����0^�b3�+Kmuou]*p\��Z��Ҟ�[��ܖ�O\��d�j��;|{�K��Ξ��DOԮ33<XW��>�-p	�>�2/&i��͵>���elӏD����U����k�d�`��N�=syM�ً���W����|x�xx�]�|p2;d�>�C�����}O}8A�8wη$�ٻs��Q#S��T&�=s�L�#vq����U���|����9�àm;'�_+s-`�,���>�ˠ���N����E�l�����#ޞ�>�,�SgI���'+zԄ��߾���^�f?���D��S؜�S��z��#sÄ�7�T�5��Y��V�w~k���o���qͲ(��mgO�.=����N�\7޺��T}4�I�6�xN��ep��냋ຼ��Oxy{ӕrn���ss���3W��{�ٱoL�^o�ՠJb�iy�+B�D���}s~�z��X�	����Fg�]dW�{Hj�&r� �Gˢ=%��vFvk3{78��ٌr���Wz�����kCN�V�xt��[�S�[���Υ��+qWV����7�����1We+ �d��v��Z���]�*T�A�Nj;�Y|�<3��G$����X�/{����OU�p�N��Y�}B\ċިZ򹖑�{tL���7�|㮮��o>b)\~T�W�_{�
f�=�N�� }���ב^�y�u@^ڭ����|��K�:o�"2�N��U}<;��b?d�q�i�UF�ŗ�4��V�qe�����r��=�q��fs�U<���]��w�h��:��EQ�U]�k�w��H�>��}�*%)�*�-Z�����¯�	*-
M׊�KccIn�eLʰ���+��q��I7�ظ�=Ad�NO9�B�b������*��5��Fy}n�T.�su.:G���	4u'�b�\��:?���x�̏���߿^��ɷ�#��bj; �&8�(��}��ʚ�h1���C���b2����{ԇ�<\�����FSǱ��n"�M@��D�1���>
�U������m����f�v�f��P��L����3��}b��ޙ�"Jz:V���u��Z�nT�'{Z!�H��=3O*Cb��M3O�=�,߲�m������V��|6e^{-xό��GP�\KW:&��7۝����a��\�ff��ƥ������e��|3��jl��e�R�s1ř���_�7]k���:©ӳFh��ь�:D�Mq�
��><3�tx�<��l���^أ-��rtC�v���F�l�'�8C�a�=կV���)E,�<.�k{
�^�J�V-���]E���S���(����d�s#ׇo{9b>��QeGK�P�nyU��߫����)W�}V�J����O��u��Or�ge�-����c��?�BZ�\r�m�ןe�����y*��u�JOJ����m_=�&�uڱ�	.�o��ʣ=��}��I�<��C�*�W=~�̧L7��\��@��ˆ���f����`��qJyv<^��O���Z�C���o_έ�^��tڮ���e�y�y{�*aw�_	�q�]gkB���'1���]��64{�#0��L���/�Ҍ.����K�=����@����^`�U�w��w��J��7�0��O������~&����P>��qК����*#��6}2��'<��"�.O-�}x�����y/���-��qx�l_@�ܮ�s�yGs�,�e4��Ig!����,͜4�����D�1]�)��Ex�ޅf�noj��� ̃h�,��N��u�x�Kle�y@:���Rsr�����;R~�͡K���H$8�#I�_�k��"�Yd�t�d#Mc�6���3!��\	�r�|r���L��j��J�Qu&A�m��ѧz��1���?}��g�}��0�=g���o�L�ʇ{ޚ�
�*�}s7 :�&2�PνGݚ� ;�x֤�[Y:�grɽ��p˅lgD���}3]xh����L��VFw�/�j�vN#\��jf�)XU �4�1�^Ǐ�j=����C�j�O��O܇x{�I����"�뽄�%�áZ�ye����v}�W�[��]H�����ϓ�xz�����ٻ�$�)��� 7&�;��L d��3��O|V�,��f���޵κ��z,,���S�ʡ��ۑ3����g�kX�y��g��"8/������Z�ε�ܡ�����\�z�fwúIE5g��O�[�A攺��S�`������/)�0�l�V<�����`��~���_׾�����D���Mγ/������RLUz�G��ך�j]��'~5��>�޷ل��5|�N�-���X���7�:Y�
&d�B���<S�ʯ��K�[啻���	��*C��Վ-��7Zd��"��sE<��T[8+�tV�[Ut5>��݃�dPX��q�̛�����b+�;�R�]|�e�P���8�{����Cj�����e�/&�ÿe R�W��[u�-o�_�E��ǋ�w(���R�Rc!9Ҷ��%J�h{�� �_Y����W���8oeu��N���m�&u��	&'�=K2k}��ӏQƖ���1��ؓs�ף-���i9�c+�y�}X�fZ�'�󚞃�N�Y�w���cDvvT���=#ۙ�m	Y�<���S&{'������~��m��c��&E��َ�)cF��p��8�KM'�Id6���#6Ԧx����;20f���Wv����� �C��A�[��׾��rk��io�uO���O���y�k,L�z�n����-=�}cg6,��>�M���,ғ���Q��2�c�������5=�g�G��8c��f+�z������<�	�1�ޙ��PՑ�kǖʗܫ�
ޡb3|���G��˻�VfGxՀ4KK^sjH���}�:j�����W���������bk�?}����hVqu�s��FC>��)�k#5�\��GF��mZ.��U�rj��H��}�՘��XVn<��ޒ*�ڰ�^�ڏ^]s���*�bb�t:�,�x�=i�{)�� ���Lx0v�����r���4�x V��xa2vrG��rӏ�;f,��{k��W�N��o�z�&,i`=<#�{z�,Fu��ٕ�h���5��9 \8s[��d:\s�C@�>�^�9�Ǿ~6�����-f<�T��Gc�v;��}dۅ+pJ��M���=`�w��}�Z�}ZgI�9{�B�s�_{�8��w�b��c�cPO��H�.̞N��?.��~�/��ٔ읛�>P��mgʣ<���?�S�jf�`�[O8x���m�+�W�8�k|�Kz�s�̝?nn�>}5�Q]~�sٱ޺�����ieg����V����˷}����u0����������sW���4�&��ď.ʑ�̼����/�cU�Y]�s��LY��n���g�u������3�4ՈC��h���s�.�z#SJ���߮#�w�ɬU.^�8�P�n�a���D.�%(r��s9��zz���n�ނ�o� Z�Q^��ӞV]M����W��\_Z'b������k�ql7���sp�Lc�Nu��W�hȚ�v����c�1�kX}�nQ�G���p��x|��ԩ1�d̹׭��l��R��.�7:���`�H9ոp�yKU(��f�K�����9��:f�5�^S���M(�e�b�.ے��]�����ߔ���J[���0���0fG�]���;��0�	)�������°���ٛ�$4���'{�]7"�W�j��w�n=(F8��W`&���[�T�3}���W�<��*���g�*Y�H��t�^���v,Pj���Q����is����|��ޝ���}��pb4���2Ig����l�By��W�5�un����6xw$�M��K�7v�݋c���1v��yЯEծh�#_y�6���������ξ8������Y�7��?�c����O�7f����th^�Bu�GZ�*��7��̝�M��qO��<���E>v�i}�"y]����y�y��d�i��M};4�%)�.�gջ�%\=�2��]GGi��(RzxRhdu�r��l]@r�R����>�R�ݔ>�	�����sY-ͺ�5Ω^�٘��D�*�V�,g��zp'���Sv=�;�Ւ)�[��[��cc�z�+m]���+��ė6�o�5�f^�e^�(���M�]�����)�w�m^r�F���RI�)]C��[��6���;�)EM3@^�����YfJ4�Օ�%@R�N����2�9�TKC[�4�����ic��(D�-�o�j�T�M4��gQ:s9.��A��+�Et �����
wUl�ec���9�*�z7��%~ʖ�oڦϓ�1�1�s�����{��|���7�۬���F/�wE��@��W<�?O��ڹwBsE>��9Òϳp�MuBa�J������2ehn��X��	��J�+m��F+T6���.���V�z�<`��V=͢5�_e_u��=fc~E���sǤ��P~dĝ�g԰�����ﴇՑW\:��N_�3N�~�m�y������ ʏwS��m̓0pϖu�[�k^�~�$��_z��dn����MV���8���	�{Y
�v�}�}į�g3��?�J�S��J���֯_���ơ�ݹدF���jǧ�I�3`����LW��=��s��9���5,�U�Ī��O]��;�F1�8/��=O���w�q�_}Wm��?� ��4��m��+��Z=X��U����Np���E`Ψ�I|6��z���멊ǈ�m�,�7���&��{2V�w`ԣ}ӣ�7Q�wƕ �{�!~,m�D�a�^K��t�˙��Iu�2����Pr��Ñ3&��
�ҹ)[$a��Q���C�*�5�M1�� ��ˋ��,���gH W%-ʾ�ޖST��/3�3���Z��{(I�Qպ:�i��oWu�Rȝ��4���]n�޸s8��n��@�<��x�-�,X�bg�E�Wׇn�:��ʒ������??d���xu@��']ɋOVp�fl.b��]7]�7�_�QӾy�s�iuԹ�x9e���>j�qv�˶ݹ[�ekC��9�e���~�߫��A>�������'R��=�-H��efF^�#��.�~�ߪ�]�U[u@�W�}ۙ�����<>�d�gْ<��'���>���`�]�_y���}���H����;r�vt��3�I%a�q7�~�������{�����~�T!<Bs��c����~����y���� =���^O̟�r���`fw�}��>a�I	{��2��q	�6?{N��V�9��:�L�����;�p��!=C�|�ˌ	�f@�茶S�����9���X}���<�B�x�'1�ߩ ���<�g��=�^��OX@��$紏9�{����y����~�@ u�Z�������5�HS�|��f�f�oo֫����d�V���j�]�{^�*:� ��	:�o뢺�F\��2\��,*�)^�tٙwW��~�J�[��v��=�u�΋�>ș��e#?~������"h�.��f�uj��B�~����)�]���V�R�(�����-ۃ7j���Tiؿn�W�x�������k{P
�Y���go��ϝ�ǘp�������6k5�B�$�z��k b �!� q�J�����x��)���^�4N�q�!�I&����}���}����$'7�/9�߰}��<�]9�w/���s��ϼ����$!�$8��jx�@��� ��<HaKO�l'�ne���rC������_�&+i�m��-�	�`6贛tD"�m6�m��D��$+v��n�ʝSa�!E��4C+�"�;�}x��+�n�pԡ5��1]���6�-�X��񩕵��)��/x�S�8�9$��	<���������2�%~�������|e���frW���o�;W4�Z�:��ՂP�S���W��\�S���a�ofV�z�:���i9a�.?:����挬�4���i�G����+v���6�8oh t���Glv.R>Q\LK�8zI��t;�	9���$�F�l��Ďf���zv] :�]u��ۏ$�]��mK2��{�/9,��vD�<ּ��z*N�� r��NT�����Y�XD���YU0
��H��q�E���3
�$[���Sk�)�OD�Y�ʸ2�,�G
F
�T���ILC�9T��.��B!O֓��r�I#=-� ���"�Qm����)�*�_�:m�n4u�tݺ\���-��ݻ[Gn�k��+����w-+�m���W;kx� �p6Ͷ���q+���ߟ�2���3X��~�� 't�{�Q����QrOT9����NeEl����
�����Π�"j<���jTv�̱u֯�R��ɴ�]F,G^<������=�����W��wt�:��v�Ӯ�<qM���p�Wx�o�,oZ|j���B�ʍ��@�*wP]��vg+��U)ٖ	�B	|��@��{����Y*�MS��ڬ0]��D�)VR�3[��n0���[��zt�}Os�TV��mk�n�c/��U_��K��G����z����u֯WIAnQ��ܻR�9��NN�]}ݡ��PxR��!���Pbܙ�8�'L}��u��s���7��h���+܍SW�E�;-o������y���K�7���A��Em��*�b��2���"��nnŦ���O;�^�m��fv� �ۿ%�s=��]MN	�ѻ {X���t9�}���_�#e{���w6}�����뉠�]�
HG֫����K��z����2_')v���6^{2��Hchz^��z���P�u��S�3��{��Lf��RL��9�-�Ǖ��(=٠ٽ��K�u�^�W[re'���r\�6�}%�k4�*3�_����#��;؏�S�=�Z���ݫbfpW�x���[[]lw��W�k�lҺ���8��Z���>u�8q�s����z}�>�{w�s��g�Pc)�{��}�Z*������+
��?E�ѵB���S��W᷵��}�R�����}�c�?�p���z=�ラ��Ҵ|F9a|�|y�|�yA�ͺ��L�\�h�U���(����}И�
Ӯ�s�w~�y��A���V3u*n����������S���
��s�-)�c�:��[`f�����r�w�0N.�=9��Ãb`�nq�WkK����ܤ���0���ґOq�]��;�x�j}�O73����a���t���=����E�d�3ʌĜ
g͕��1���w�j9A0T�W�9���Z�^����ǿ}�7��}����̾$���o�;������s�S��P o��:����7�����>�a=��|o���u�3��?��f_��Y�����獼�_�楻���o��{�M{�5[�������G�_���sW�����"~{��.��pM����7��5�D�<��-�*�h��.������w}y�s�w���:���\9�7��e�����坧f�T_]�|�v����uԩ.�$7�SKf��]y����x�Q�U�$��q�F�Q�*ӛ�����I�ۀu�/m��ϒe��i1ʅ�=Y�:����L��ХGr���&y�z�����_�m+���CB�=-j0(�NN�������.�8���o����/p��҃mu�qy$�'�3ME%-�KyҔw��F����s�4�f�J{v���)�ծ�����{�j���`n�;8W,��F$�mkj����xs�nӼYK�i�s�) �q�t\�����{�v�w��4vn�K�WN��ie���n�ar��ܤ�UD�����)�u���.����=z�Rg_.����T�%�d&ܚ�O��� �un�_Վ��]2"��9�Ȳr�be�0��E�FG����:����tV���Ϯ쑜c��K�!svVk���I����
�Q Vb�0�cc��ݼ�}e���,y����r��/�j_e���+3q�3�Su36}(&��;#x�_��ن7ÄŻ>ɱ��Mz{�o��J�WO�5�St6*��>�B7�~�װA=/;�5ރ*�Òr������v�zj왓5}r�~j��Ӊ|�vş�����n;>G\{���\#�����Z�h���l�ڬ�M��E]X�|��;�W�̋�D�`����{��f����(:��ܗ0d[���\��HW�D��Oz+������=s+��k.�I���!t��#�~�D�qJ{����R��ؼ����R�P��^�GYBs���{]�����ǆ�z�ғG}��lU�˧����{�f���6���>��AC�@��DF�B�z�N+.#1W,���j�J�8s	��aЮy���7���]\�}&mBJ��-N��/�e]D%4
P� �".��BM�I��'M�I��v�n��Z�R�U����*T��*��g-�掟]��g��;|��7�7�݇�yԼ3C����	����՗k�{�Y;_wb����wc�fʏt���hR��V�[~����Y��֞mf}<h��ޫ�7���/S��:��� �����/;���W�R>A��O9���ԗ<�i����Pf*�C�9۝����#gw�|�j=�����]�wvsKخ�R�
�����J��/,����O_��xA�C�uW�{��ǐ8���z�U��~2��p�z�`�"�/J=��&z�r�M�+����t��mvª�}4�_�����^�n���V�6�]B��%z����7H���k/;P�����������Y���	�����瞯���d{�z���fF^ؐļ��e{�*���߇�{||T�zmı�o'�*�\:��#|2g���wﶶ�l��I��U���E^�xs��p��WU�k�_�3�����lK��o��;Z��$��mv�uҳ1�"���!s�Q�ے����a����,�-?���n*�K�y�}L�ٷ�s���$�Z}���G�46�党���e�nB=��ro�~���*J�}� 5*.�b�<�7�	@)�ǩ�R�qk��:������o�vV��T������h��������A��Y~��7L��b�߫;�&�ۼS⳱��ûӲ;/�1C��:����͹��g�춷9�!=�O'[��d�a]�k�&���ԉ��˟k��ˑ`��D�X\{�����%�n�أ˸{8�L���Z��,�";��^���P�����=N���ԯ;�񤖬%���ם�95�
yO@)^4T���ep�	ڽG�|g�羛]F7z�_�#���y��26�(ú3Tit���&�0�k�݇�z�Q�*?�V��3��{�3{ٹz��o�waJ��wQU�wm5+�|�y�z6wA}R�R��|��"���ڽ�0WU'��r{RוF���'����q�;�T���W��c�s6���ĳ�˪�*�x�۶O����z�P�����r��}���}���� ������&j0GU1�s�� 
k�!D��цn�.p*�KA���]�W�ljX�v-���R�՝�ԯ+��@��ES�*t{;��5���r���G�́��U`y^[�C��]f�y���ri���T-)�X�H�Σ��}Z��ґ��[��G0��\��HI.𱃍�5x��E����T��i�Ib�]��qO��J.�`�����ʻ�~��9�JD�l�{���ۊῺߓ��>�Ϯ3=��jw��צ:�����?jCd�>��{�g�e'��vB�}=o�}�O���%lxq��J�v�����v.��@�Jp�3�N�/\�Z�W����Ɗ��s��\[�b�9��Q��:����0*��gȉu`�������F~�ɓ��k��bHM��!v��~�>ｽ���3��TO���{=�O�N��z�����튌[�f֖ F�6��#"Z�Wk*ko���.>-)��>�ʟ]�|o����NyY�o���Y��B�"���)o��|U�[Y�m$�/�C:��C�Ŀ���[����a�ُp;w��b3��̏��$��^ᗧ�s�#ɾ{Z�ׁ��b�߲�s�&c��S��/���;��"UR�q76���n��>����=E��mҕ�]�p��Z����+�vN�s���tæ̓��~��{ �1�
��r�>�ݽDh"{#�oV�Xp�^l���{��w;t��R��v1K8D�Z(��ޙ�u�4j��Y7�qG&��jl��m'"��]·`Z�A�>�W�/`�=������0�N���*�uȎ�oS���=�[��غ)g���L�?��jEkz^�Ӱ_(;	�^�[ѨI*�������W�X��o�g_*�U�x��prkD�4f:�	������[��u��\�j���L��J��zT�o=(��+��������-��8�8=S�zx�:�'tҫ�7y�N�w�^��>�.%ڟ,BP7�����s��|>E]\;[�<�����\�W*�ۺ�'O�����8�_{�
��w��MV�O���]���i󼷉 �Z�����۪�����b׾�{fo��/�C�R��A+/�[��@��uvqۉ���Ãr-%aM�+5�R�Q��vz5��?	�8�Q�ᱬ���UҊ��nX���
��w��¥t��<P�����i3������-��Ϻ`i*�t��^3�}�����ϊ���[.�>p�_2}ڰ	�nF�[��"+c2����w�f��v�rVj�þ.�mx,�;���v��Z=����s�N=���8���c�ba��t���'�Yw�>*��آ�,���t��kM�4.l��+./w���(J�yد6v�Q��?�ξbe pT$�*'3,����,C�ZN'�D��XC��WoN�s���w����8v�p�q�QW��hУ��[f�hE��u�n�9�D�*j�+��۵���a>��d�aZ�1Ďx���'���4P��Ɣ*WGs2X���%NjG�M�#�=�H��j�|!�ӓ��|��>��z��kr���Ϥw?Et���7�K�~ߢ�7�no�hP�O�׮��x��5�(l"�>��r�ݨD	��)�U����O�b{�����u��ψo���{�[w����ܙ��e���U��z4������{+6���U����,�w����=���Sq�{)�O\�5���c;�3�q�}�o�Fץ�F/�R���VOAZ�e�������~�^�v��O�{�oWMx�]x���t���.2�O�ؖ�d��֯ǫ<��U�[��Wo�$���u�b'*8��g�4���3"c�9�H�|>��1���~T�z�}��f�����f�&��Y�qek�F������qu~�Y�>�0f,YY�{O�T�O�m}.�_5ol/d��?_96�'���]ɾ��{7funDl��\n�,���>���<˔��'��EN�]\��}]��F��;���y�Փ���[�y�+0[(��R����B`���Kv�9�5U��9���ۋ�6�TU�>��������q��~���ҺNZ�2ӝ�|B��{\�{�8&��mf�N����W~��y���1~���T%�r�A}���z�ۦsw{t��f+��:�}���T�v7i�}�����7罀dX1={ɇ���eu�֍M��v+��<g٬�\yR�`}[ݱEGr�Ye�(�A����֥4b��n!K�R_M8�{��� ?�>�G�x:���Q�Q�Ѿ#�O둆:���E��ʝoz}��>��:9�.����dϒ\��1��^��^�K��N>�g��8s>д֫��+��&	�O�l��D���y�d��l��+'p��`�>��
�F9	��3������F�q�a{ά^���ޕ袳oV��J�~¼���bi���5�q=*���}O�9jw��t��0�-d�$��[�l���L��ᚠ�wr����z{H�C7{��s��?���
�~�����~�����x[3'����z�̺0�ĕ=8@N�S 	*��2v�c�Ȯ�U��K������)�)��΢-D?0w,p��۵�`]��FmM��P�7G�%��9�9��tk��x�ʾ�&av��33���|i��^�#����{f�`7���"��}n�觾�uw�=*E_��]Q�Z��~�Q�����_��bo�&�'H�ia�O���5����S�l�>�.eb���w}����a��Cݬ�N:��er�s42���R��/�	�/G4����F+����Щ�:���-��ڹݍ�7�t��^����X7:k�u�pV��|�<���qu�!��W�xS�n��z�m����4�3|�m=������������`smI���?H|���`%VH�)]M*���;zU�C⽇�+C����������]"��^h��P0Vl���b�i�������������A��ocΪ �^͞ك��;d��v��TY!,��cw�U��Uֻ�!b�a�� fm����cN#WH
�\�J���Vߞڬ�t�׽�����B��>���;���/�eW{�.�z��̌�
��a�O��=@H��U�O_�!���.��~6�]9h��<zcBd}��Qv^��v��vq�L1��#w��֕�^b:��t����:���v_]<|���q˙fw0u��!�ɣӖ�+�n9�']<�3`Jo:6�qd��4Ѐeu&t5��S�x�I��J��u7h�U��
׶+j�;�7�n�o��|9�gx%1�W�R�^Ǎ�Y�3�ob�5�҄%A�8"]X����ߙ��V���l�sN�,u
=}9E�����T�(�ݺ]�S�|5ʋ���]W��e���^^��2u�O�ޫU?�̆�M��cޜ;ٵ]���ib�VQ�7J>�tv�a��O&n�W�^����n�/ԟ7M�L�b)�nu>�ҫ[2Xp���Rr�E:}�?߲�ĢƏgQ4�ħ4K"���ѽ����9+�]�37L%4��F�]|�:&o��t7�-��Eq��]:�~�_�8]ŢҤ�/�^�He3�UW��9y�6��ʈ�^k���}��@�	"�Bj@}�)���]&\�����o'��ѦD�ءP��e�r��L�N������V%�ġ6�e�b�Z�̭Q�m�4j}�2�kC����e�x�g#���r�ڝ@h<nv��U�f��2͇{+�kX��xj�f�cV�g��.G1e�3�ś2[ݿҲ���3���0Z�E��]�aN��$�A��+������!=�������m�}s�����!�^]��KU<��Z.0���Y.�����\?�sU�;\�G�-��MclCtQ��U�gQˀ�V��Yҧmr�y�+��$�'h�P~���C�: ؔY�Y �Yn��Q���I��-��'/���qC��f콌g'�^ɳF��]�t�Wu�q�9Z�rp�O/4�5��ͭB89ӄ����Ɩ���9A�α���w �v�sz�kU7�W�{4ğ��5Bd��!Uf�z�kiq�Z�ZPY����Y(���˨�5)�$���<3��jD=�`�ۻߙ=�e#|�Y}�1����~)���/�U���j�fD% +�>�3�+�2�ܰ��YW:�^-DJ��Ă�1�� ��-ź;t��Tܙ��݌x^�}��e��2B�t�/�7��bm�K�z�o_V\�yJ��k4�6�q��B�d�����I*9�\�U�����L[��s9�bz�^٥ίP���V+k-�qcgQ�l9�P�D���nQx���ՙ(��eU՗���pP���*<��}[�)�3�-�Y�v&�gJ���Ӕe=C!��ޯR���'�ߑ䌸�:����!�}u��Ωxf=�a��zQ�:�ʊ�B]:�Cf��OpM
t�|k��:��Z-2~�-V��{�mT�w��-�X1�#��� ��(��ɓ�܋6�K���
|�U�	��ua���\E��D}��߆��4�<�^^l���B��ѓ��P�s��V{D�#�;�vm���s\���*�]�ǭ�E@��&���.���,��у*�#���2}u���X_e������w�}ܵ�<��z��z�ތ�����Lr˼�4�<�/�HyR>�'[��
o���K%Uᇧo�1��L�X{+:�3��s����G�wG���Cce��{=b��Ӕ�:��_�0�o���y��[p��
�+�O�2�6�Ͻ^�����x� ��~�(C}�{x��fP+�=4�#���^�c,c"��B�F��y�1){��z���9�woK�Q0������G�7:&���+<��}u�x�H���vO{�]�Enڬ��[x��t5
���Y�K=�DߕE*eI��<���W�N���ƒ����M���ݹ0ˬqY|hU9��b���{mR��O�qIkI��Q6���2%ח)������z����߅ř���v��H���o.�/۽��g��K��g3�	mv� ������!x�w���e��� �ҕ@Rj��:��i���c�`��e�7<��i�އ�;R��F|���JC� ���ӹJ���<���f-c#�L]?&�m�i4F�@��m��Һ���c��k���F�.?mh[�u÷$.�stsm�fk��Gz}[՞���w����(�=���Ao���b���T�8>�r�SH>W��*_��涮,����]��|�M3��1����z�N��"���pmft�v
���ŷ�4���%�<"�}�(����+/G_�Y�.���r��v�ώ���%P>��*|/���kI�kw�خЪ���L��9�^ǔ��+�Nh[=!��U�I���Hn�ƺv��t�} a<�������a����Ӟm)��D垚1oh��N��1�h)]B��!O�3s�����
f��
��u�t������>�P:to�C�U`9�p���]���g|.m�xdo�=�۹5p��.���}��u`��)F�=����FG�YK.pğe�1�Q�μuiT�>F�(e�{wJ=�t����]���J�{])��o^�ֲ��Iy^G�4�o=��ƣ�wn�W�q�w�j��h3�R�t��}X��s��ʛ���D�'7&�\�>������G4d�GM���5ܹ��u�L][����C��(Q�`p�r�X���HR��$�ۅ��ꚟj�V�2b�U�<��-IV;��O���)QdZU�
��N��`䫣��s[Su,5/�}���u>�%sn3��z�w�'��v��d�f|q�Ղ��ct��I*z�6�eK�^�,_�kh�o9_��NS{����a=�#ٳn�+��Ц�#;�]�fDp�fwp'`�75�q>��^g�3����ǲ�dNW�{$]�S�?�8�+�U;֦^��nEQ#����ܞ�C��0���W���˸��U��~�/�ݺ0�@�3QObdpI�>�4�(>���Y�r<�j/����_��\��ʻ��yj�i)�߅m��6�r�q���h������f����Mev�V���~������?�{;�]Op��m�%��~-�Ӿ���ҕJ�d�*�J����H�q���A�ur]�=~v���g�	��=�_�W�^�� �뗄����{����3��6��1��+��)����W�4׷Ϫ޸��c{�9�}�I��L�ӟ!�t�l��f�vD��4���$T� ���]�p	{�$9velE�O�x@ۻ��@i�#�s��t5*L;����R�ò����;:�[[P�ϧL�����nrA�M]��e���+�b����]���{�I�� 㴞F���y���U7¥	�}�#����Bt}�ҋ��_k�]Յ��cM�g֩����/rc��*��5N��_��gk���DO��D���%�f|����Y�%��DzÛpB�z1`���avS�+�q��Ov��_O{3��J�ۺ2���o~r�3�o���J�XF7�)2;
x�*���n��O���H�|5k��J�=������ʺ�01�xZꌨ���\�Ed��]O�|#�،q�I^��C�����n�����T�.��s5�?�Ϟ����G�}����d�ޠ��W]JW��)O74~�%u��Ε����z��9�KƜǆ{"��*c&9l�|+��G�um�gynR�U�3�R��^�Eօ5�_f��ʊ�^�/����0mn��t�b�O��i`��ƒ�GWz�N����85�9�O�-���V����C���@]��^t~>H����iME�aǝ��5��+�Z<���;������]"�V���S�F�^^ĸ��͍�=�hr�K�<̜�[�*���0�Q��^�kh[O:���J�V�K5��JN�]5�w�[j��h5�p��RIf�a��޾λ}�3��8+S�����[Vv,�ӓ�Rs=yK!�f�K�����f���{(�/��ްL\�Z�~R�V�w���E�dy#��>��^�{"���9�hZ�*���r��M��vxΌ�'gm0r߇�&)B��nܸ,@={�s��Vfy��p��O7�l���#��Vd{����i'fq�}�Uxh�K��R�"����7*Z�}�3~�g=���٨����vN��y�žΐP�Zܾ��������.uA��W���|Jk��5��h �w{6����s<A.�'*\T��Cng����n3�+��] �=%j�7f��U�͏�W#��^��`O�'�S<�Y'��L��/ev�k���{�TU[M�������
����b����C�F4)������>�Oz���j���k|�..z�\�{���s�����Ǿ�|[׬��d�}�V�_��o;���/n��=0m�J?q�}��Y8�~^������f��<�*�z2T��Y:�W��[�:oR�K������9έ-dYKJS�՛����RT(A�(@���o��T�Ѝ77����8���z@\A�P�ȒX�VF�PܸfY�m\k��*�R�"�C{��<�R&u��Y�!������F�V�t�\��a�Ka�[g��Xݹ�Wn͋,΂����/��{o�t��3i���%�S��T<M�yp��77|e��G�ňƷ��噴��麊��+���Q=���l��/T�i�{�L��7c�g��I:��J�����`We���r�o^v{���ej������Ӎv\G�M>b`�e��l/Z��w��[���[Š�K=���i������Z���虹�5�]�v���X�mw1?'ȹ�lږR�����q&��]�g}�Dw��h�����}��Qģ�G�z��?0�y=�w]��aW�6C�\�?;_#�+e��.
��<�2){a]��mK��J&�R��]�e4��ɡ��kb��*���H{Ӳn���	���1Xz�x{�Ĉ�ӼÈ~\f�0;B7�3����d�Q�/��<�?9��pԟ�g����/@���F�磘y����O�S�:��8�K�U/O��U�=�$��*�Wo
�w�=��p�X��U����<⭥@ad�a�_f�+9�;�t�V��N�Ċ��w#��9�-�H�e��&9�`�ꄞ�)�]�RUҁ[ݴ
���ە3Gu�m�Ⱥķ;��Z�7��Vs �Giwe�U8�R��TnyL'! 6c����oU�꺘\�[=P�������3��Cp����Q�b�}�=�.��ic��wgz �Y���]̊ٸx#ϐ��B�����x��R���=�^��v�q/�Z���������t/@�m��\ϳ^w�"�G=�(�	��N�С�uLQ�Y���5�Z>��M�J���['V/)^�����,�q��Pt,�y���U>���On�ת�����Pk��.��N���ޓ����N?er�8,ʬ����g=]�z�Be���SJ��s�Vх{��]���#����+n��v��ʜJ�bRGOn�T�nTWl_����������_��͕u�2}�	�s÷���*�����{����|�K�}'ܯ�ٱB�Q5�V|���Y쥑�v�.Ӱ�9n$vӁ�7�N�/�1C�;��a>�1���+���j_y�ͻ�.b��͵��\.����1nn	�[�E�-7�H�c���E�~Њ��Ⱥ>�l�@���f},��#�](2�ObrL3^�m�}C�l����$esB��0�˖�u���z\o^e��|��w����_i�#V�d̦��w���x�����x���$<e�x�q�Bs���[��2|W�}P-���X�~<�*g�w��Ua�j�[�O�w{V����TTM-�=��{�?e�^?`ʍ��S_�g��X	��~� �3�q+<k�^�=���N��&P��{5�׳�=��2/*��_ܞ�@��4�`a�_��+��Rz;��%�^?a�ẩ4�(��}w��ٛ�b�~��T࿹8���|�:�_�=ϛ���=��z��U'I���}z�W��rn-�%Y���}�Vg//�;£���m��G�i)�'� BY|Mmݫ��_ה;.`��]dz]��/�]����ޢ}�r`G���.Ǖ��( l���*7�̕;��x���L�wd�a����]d�ۯ��w"� b�J��z8�f-�k�b���&=	q�YC�y�_�Zͱʻ%�%����x,�iP@���f![�V����	pi�ڡ8^ī�h�Cp�y+�����()CE�TDV���OTZ��ɀM�:r���E�*o-oJ۹-#QBa�.���-��Z��D��Ȧ:�3���[œ'R���iM}��}�]�Xn��~��7_dZ�m��>�>JW͙���\�{מ���d.�C��_W{f�m����rQ/���k2G�E��P#9�54�Q~��'/�� T֫�eW�2+���nsG�l��ɋ�d�޷{}���W�c�$T�Yi���ۆ(���ы Aε��i��{]��S�:���.���%��3PC9�G�.s-ߧ(\P�A߿i}�3��˿|wJ��O�+b�.!qY��_o�r��P�%����Vq3�<7�3]���ߨ{��W3'�ӻۼ��ʊs��WLf���y�=����2�l9�pu���ɡ`t����<�\[fiG�v�~���H��)�ʪ���r������gxv߈v�o�~��c����yq��P��<�=�����N�V]y�.��Rw�瑓�g���t�{S-j�Vc�h�����0�VE�s;~��-��x�0�ʩ,w���������/˙�f�İRV��9�j�^>?�*�h��f��W"��t�X��_-�\�s�f��ѣ�d��Ch;Z��:�Aݡ5�**�Q9�1ܱ.&�'����yպc(B;B�b���LԦs�8X��R.�c�(�"��	ˢ�n�KA����+#�9�b�N�s^Nyɺ�8y��bz����U�����~����)���C(������ּ��mX�!S�w{�]nΉ���������PuK��y|����EH]ە�ݮ����5���td��k|fZc��{�ؽ�y�:ef��;7�dz{�5����VS�7뒌Q�#�����>��y�R�g���g>L�tɪ��-r��$����=�F�?�^���\&1i��G������՞�����z{,: ��ܒ�q������$�Ջ�j��� T���ޝ����Kv}�*�\�_}��-�SH���L�1�|�eǼ�᪋�N/'�3����c�����3�*�ɞ[���.�E���~�+ �\�TN�B�#�>WՓ�&���*��?x���>���y�ފ��l��>��Z�f���6I��о�����=�m���-��������¼c��jm���T+���{,{�8�Ez�5��= 
mH^R���c��:�*�O���l��X�R:��aIC��E��UC���H툶(��'�+n��]�8r7��*uNt��J��ak����퇺1��X*cS(q�so�_�hq_�^�W9Ӿ�SJ��]���W� ҥ��)�i-���e�:��EH�V�e_mrW��f
hqB�m�%sk�RX�u6t}jQꑻ}�3�4�b�қ�v�����.s���{]�ǹ:XyR�]rf��F�j�-h
�:���TwW+M�ً�g�K�(;�]��{��w/������X6�dW7H�)���Y�S�Sܖ��Q�L�.��u��V(Tݫ[c=fWfo
}ô��j��+���Y#�a�KP9t�Z��VP��i�'�/:���R�!��r����\�ӓC�m+�o��h�W{0�,U���ZH`�&J�����w+tRIu�klY�����_>����sYG��NX��9ͱ8���#��b��i�vp8�c�<����WYlr ������n�h����E�*�T::���l@%g<<��M�}1=W���?<ܠ<�1\I��s�q�gV6W�׌�W���Z�ηwR��i�贫]Z����r�1��#�pj���皱�3�B���pp���h�chKÙ1e-�Q��'vW>��HUԡ�՞��k�@�TttA�L�RL���o���]O6�� ��n�ҁX����*K��n*�3-� I���v�P��}j�TW���Dw*��a�7m���[a\�jY�1Ѐ�R�W/��;xj�SD+�ѢQ���U�F���qrY�m�Lm�5�m6�	2T�h���d��-��I$�%���:9��o)>��Nu�Q����lѾ�(���g�f�4�l�M�8�n�9�<XNe��""��y36�G�|YĻ����ihu��~��d�m=�@�y�)�ni�:ɇ��ֳ�_\�^>��cR�U��^\�������Zy퇴�9E�2��IW|]��+�u�5�q���5�!�jS�e�9��or�Y����A/y��ά������2:k����v�@����������Z,C���Yɽ������Es��hgZ�Y5����I�{gE<ܨ��}"j������Kุu�ε�L��V�в,�tU*��(�z^i�=�"�|�.nu�h���8�ʒ�/vR�h�bcBU1� -|� u�Y�ޒO�W����� &�m� *��6$ U�K�	$�f����y��,Wb��u�����g1b4)Jf��(�)Rl��L4G�LěT��$%@�d���E~ESt��iI�����
���e�#��|l�����D�z*{kJ��"z`�TX����_1'�r��j����!R�����-�����ِ�R���Q��5��C�
d~�ż��4�I4zvjΜX�p-��X0^��|�Lu�(h+�ظS�7��eQ��T�3)Y˗n#�tfSަ:咥G� l�6�.P`T��T��-��qS�ʓX/�C6�vY.�e��tb����B*퓺���!i�"�G5��$��Y�B�,��B�`-�6�a���UUUS���Kp3m%G)�o�&8o���:ġ'XڀJ�ݛ��1w!Z�Ǡ�B��4�p���-j"r���2���J�7�q�����:%�#Ls�*\���:��Ms�H��8Z�~ģl#�E���!��N��^�"�'޹ܘL��cw�pM�MU>3/�(r�t�wj�1�gs�{-m�F(�S�Ṻ�!&ѢW����u*��|8��S2��\H�5��OG�w]-���y�bY��~ದ:�q�9}c��3N�ϰ�}��W����j.7I�Uή����+��i��������EL�>Y_3���>p|�Ժ���&jlcޙ����P�L�m��:]��pDK�=�ٱ]�S��W����#ʼ���o�>^����
w�j�=ㆤ�trzd�lo�Ǌ�+CJ�Q&�MWJ҆��uvѭs9������k�Jũ�7^�!��N�����j|��G2���zX�8WT���W���7
z��Qs������N�9F_��z��=557ܮ���z�ԯ�iee���=��<���s��g��]�����=o(	��}�ne
t'����v�~.��ݝ��w��5�EL��y�:u�yOaCӍo:�f�N�J�C��Қ���T�Z0#�t��\�kU�^s����.����{��ƭFx�s��q�+�E���x�	����B�8�iT���0n[<���VJw7Y�Z$�`C$���o!�g~�����=��ɗ��� ����Ѹ��c��F�2c�O�ⴴ�u��z2��ػC5�&��#�]��.f����o��F���Iv4��E�^D����GAhl����o�����򷟪#�=t�d�w^'�Ŕ<N��w��ʏ�;='�� ��Irul�^e���}���:�q��2�E��-��|:�g�]�,�F�9�@�����e��x�ݍ�]�B����v�9&8��!GX��}k�t{h��Q#�5�����5���ʫZ�q������ꯁ	�+8�����>̉k�7aW����ܞ�*�u���&G�3����}Zg�_��5�J{��JдS���e=�6���!��p��d����4}K�Ubӻ��K�MbQՄޞ�3Sޞ8�������P�����+'��Q��2bǥ|*�dY���;�[�m8vC�����,�c9unﯳ�=�����A��'n���9�0��9�p�.4�U��]m/Jf&T��A���f��`qH�8�lt�ȃ��'U����^����_��w#�b��I��}�-w=p��V��SE�}��K8�o8U�0��f�칭�
O�0��*V��Ω����3���%ɘvX�W�b�����$;�x���n��Á�J}r`͟��n�Y�c$��W��-���0oՑKٞ��3�T/S��Dt�2vS� ���Ix�����<��wy�5���\�2ؚ�y����v��u��v�����z�(E��{��TR�=�RP�^���_��Y��|�ig��)LN���Q��=酙���_U����J�p]{���T�$��3ň�y�_w�m	�T�TW�%[}ӻ�$b�|6k���Ƣ@�}뎪��Is�����t�=}��^;��r&k���{�S�sa'�d�N����g�zW*�!eHx/���i���K�=�>�����n��ۉ��[;�r��Z�p��z�,WK���]髃�a�	��f�"��������%x��䖧��P����R~�.wn,55�IX��u��L��>����Ĳ�
^��ު�����oyY��f�7�T��_c��=>�Ep�>��;�ڗ'+����o�)��|�\�_Upx*l��w�@}�[x��8P:��$��0p�rbx�P�x���1���<�m�o&�\�b��e�X�]�mv�G4�=�Q�5�ʸ+:�UwYK���w^��a�+}�u�=�pg�ns 4���7c��R;9��C��בа�.�WnBЂ���@H�3;�E8�u�\�p辎w2��\��Ć��E���lv�;����uN��R�P�("x���[��y���)����Q.�J��L4�V뤠�]�s��P���qfg*t����unb�̏��{I�^3Ʈ��*�����1H���ٞ��̷'}�ڥ��x^���/A��r����$Yr���u�G��AP�d��Z-U�̳���(;b�͟� ��}��t�N��TU�UN�1ǠU1	���SSQ/aUp.�����.g���ާS��0�;�~[t��\P��ٯ_/����L}t�,Z
?lU���{���=(��J�:��y�����^�/}훇gb?25/b��M���ꖘ�>��^���u�l&�g������[��^_�ʑ����sc�>1�D�{|�'o���q���k�h���ﳃ�=��H5�)�/35O�mӖ�4�@���D����\���>s�z}����M-�H���d��=�̻k�������u�/�ߡys�W���r,!��tU�ٛ]nz�L;�Թ��C�=�{�}}�=뭾��K�P���� ������u�3��{O�ڧ㒗5����~�i���!���t���ƅ�g�j�������{�2�{�>�K���
��X�N�vi4��L\��������gm�2���h��MCG3J񮽨k�-�.�]�Iz1LѬ+
�p	�G),�w���q�:�]�da�����ޏxE�y1w�q�J>��-�wHn�k�=4*�YbW��&r�?J̬ _cV@����f|b{����A�m<�7��
�|oKA�X��={�T�y�ah���@2rnsH��R,��;ʳX�?PH�������.�|�OU����5�S	��x�"^p�hLtvx;��w/8Ժ-l�����]���9Go6w�OA��#gj8��������D���.�׫8��t������f{�?�\LYݢ6L��½;��f���Gvꀏe>�����S '�pi{�0�����$��{&�&���y]E �ḇ�3n����>/�q�=P4 ��t��8H�J�7ٮ�~/2�.5�~�5���#0k+�]u�Qw���''�:���u�m��y�S���}�rC�T��%\U��ܛc޼%x�E��I���:O/�8;�nդ��v�ˍ�xMe���Dkb|:,3⣌�;u*�c��ʱX����j@UTyC<{�7�b=j��G`|%Hڙ�-3�������EM>�L��=�u��|�|ĺ�~���{I���ۦ�D�G�����n�_a�$��V9t	�;[S�^�U�z�����F��c{[���ɢ��Qu=���d�"��̖9�.��=!<7�t8[��=���wt��4f�E�r��v�G����ͨx5O�/���l��GN��2<{�zJ�wѧ�π�U����~��h�7a�	j��]z�Ӎ�eT�M�6:&��'u�;�Y�Ǡw*����g|��e����j���ϱⓍ}�3�u�v w�c49�U�4�=їf�k*$^����z���u�d������g�1�W��ù�Q�ה��=y�e9�l�צ3��X��ŇU1dt�;=����|z;'��{X�{jl�A:J���S�� ]��>�kJܳ�4�����W���3�I�{��_[7&���h�}�Fg�t��y.��䕙ݗ@u��v���v��ή�a�l%�������cM���pF����#��9� Ȭ���rܙǴ�f�V߷��H�wn1�c�j�4�)���Lۙ�!���WI��U�W,�Y��̱�����MX�������U�S������p�OE�T=�>���o��g��}p�F��V��x�])z����:;��I]���z��
�e�)�8~�}�mz�1`#���UWULMFXU�2�����,bZ��z�n��v�`R�o�wAZo6�u���I����ih/#�͕(�wLc��k�������][:u��\����.��Ԇ��R��:U z�l��M�БP����ۖ͞�St��]ZqXo�,��w6�J�^��G�-X�����j�3�����n2��ߢ��+!�
_���+%�s�����W�r��S�?�n���m���l7U���e�������/�*5t�l\n����$qYO�}�{�}��G�Qs_K�a{%��d�_S���������\�ʮJ|�ø 0���p6Ћk��m�Ǭ�gR�n��ں�~��x�-��Ꜯb��R�g���+*$����}�L��(3ˏG���x��?o�:U?lέ�uހ$_A��Ci�G"\�(ɱ����}&乷��O���YxGUӮ����z�͋�ۋ���DtM��N����y�!�E��z��\��H�4���4�N��qy[��!|��LΚ����7����{.'t�Π��Q'���p��z�D�5����1b�AF'�6 S	��^�����*�P���s�,���g�������Ҩ	�k�t鮆��e\c�R.y;rX�h��u8��:��aB���}q\��Ǉ�-[����	��ȟT
�+XU�V�tW����u����duw��(����9��/�cP�ف�@��s�X�8��w}ko$��u:���̽������9[���s����n���4̩W�f��f�7HJ-/��T`5�M��k�[�9]��������J��蔆���b���e���B
�e�!$��a�i��2��]�2V�,�(�ÙW�T� -���x&q��3�99�	�Zߚ"_+Q��o�Y�O»_{�`{u<�9��/��4��KZ��iܛ,}�,/�6�GŴ��Ǭb�V���jb��U=3�
�>���OP����3K/\�h��A���`�"+39����u�� }[�ѭ��v����G�n�叟V�FPh��x �Ĝ�]�M朄:66I3�z�L�LO��h��n�g�7���M���#�^��_��JπqQ�Ѵ�n2fay��W�Q&����ģ}�;��4f(�J<'y}{�y�JS�����~���i�7>ڭ��T$�g��r�����������w2�?9h����8�#����m+Քz�f<�[��9��VA����3���񠹩T��!\
���:���ٹ�Ҏaə�<����A�{2<��ٔ�uC��T���DԮ4%�+����.7[3W���=�0�W=�d��Atur�\N�5�|���� ��9ُ������W5�m!Ә+fƣb;xI�h���.9{��)�X��Ǧ�
������3��zf��U&�Q�vb@���U�{W��o����̮�L�9M�.Pl���ú��������`�AN]�������u�ë��>ƻ �:��"cy����bc�mLuy2qX��+�,��u@��S���ݮ�8��E,��ה��VƞCʌ��E�o�U��|$Phz[��k��%iѲ=�H��_c���Wg�/$�Q�z�ס��x����d^�4�����8���:6|+�<�ӂk�Q����#ʈ�{^���;�n*��N�{el�5i\p�1����?)�E~2K���~X�n���&^X5}7�|�g���n���3ޏrc��^�U�m��0�T�ۭz�)㬧E���zk�O�ݴ��^���Pg�e�P�:�O_iu/�ᐦ����R�v�N�+26���x��V{ތ�P�ݝ�6k՗/��7k��3
l���O����u�A�C��d��a�u�ٌ.&}�/% _]���|�r=���H\q�JUS���9cvү
��cM�SeUN{��2�3�4�,��l��1����[�&�-�;C.���p��gk��&(6pO9�q�V�o���c�S�}���Qi�/����5B��*�3/�z��y3>^H���0m���24���>qv/�ב'Wj�r��w�Ҡ����N���g���8<��[��*O�p�C
]Źk� *�8���v�ܓO9�NRI���bu��4��W�]Uc7��ιϷR�9����"�+j0=C!���N�Hn��$�Ǖ���$;�~X�TswE� H'9gޟL���.���"�7}x��]��I��)�Hc��on϶��z͇�}��xs�_��͏��WA�#�'�X`P}�i�w�\~���e߮]vZ;��,�:M�]P�����V���ϱ�%�Z����#�����4j^�ۘЇ� �����NZ[ӝ>}tʢ=�V�`���'�����Q�N��8���4��y:/^���?/OkT�طw�|k\�9Gݗ�6�dGy���V|�'�x�$�tRL�{7j�P�$�����m��y�k��AW;��^ҩ��.UtxO��?_�=���sn�?����aټ5��nl��&C�
�H�[�Cا��ׅ�Vdml��`��@�3`���Wцݩ�L�}�g�K��3:�L-x�@Z�����`Β��M��nˍ�UǺ��v��YD����1�&bq��(���vj^��J�e��e�N.9��h���ݶ�w6x�lvk�'p�0TqgH톾G]�W�v|�s��oT�2ٽ�e�"݋�k|�"s�K�������!��L9Yj�goV�C���X�D�@���f��c%�kT��?C�PyО�ɕ%B�8s6��NU�ƚKڝ�9W�޲�-oX��7yr:-bxy^�WY\���c��{y�eL<��԰���@��!Q4�ͳN�ѵ\	��p:;י��D�"Gd�i[ހWh�<%�rX��[T���шI��2��X$��*u@q�k�����o�'��Z�\����V��S�U�>�i=�ln1���J٤��ez��<5���u�gs7!2WdR&# �V�sMB(w�f��#�G{n�ĤC���Nw�u �_a�o+cf��oSX4��a'��7���|`�˻�flX�(E�;p���h��Y8:���2��;��s��OlTlųO皭X����ރ��LA�
���9��X{��n�ɖUJ'��AS��n��ø��y��-b�}\s�aT�tr���N�+xKzU4�ͼ�/%�;�^v�y���ioh��Goܵ]�$���+!�4p���7���;�6rQf�[��P��:\��w�T1�x![2���.��3�f��!�E��4��1�����J�^���̝�h�6fF��7;<�u��O�nM�g�*�i�4N���E0Ք���0Mޠģ�n��T���tQbf038ǵ���^/�{�;���+���h���j��.Gj��lu��b�kT�ܽ��wY�Z:��ܦ�_u	�E0�F)FT��#۲N��$���!�_��뾺�)�[ܧ��t򺔸�헛;����V:{ۋpIٻ�,�gHa��2�;ɺ"��Ǽa정l��3��d���O{pѹܒ�8�Rfg5|��sQ�����`��rv��\���gY��Wn��V�TY7��~ܒ�3�������!�P@���J��{	o$��7]]����\WÐ`70�Ӈ�(��6�����(�+09����r���M��Q:��)�XlS�	{[�u���vuT:�|E�]|w[K�I[�;�`W�^��=s��s�"j�q�Q�3lK��z�����t���b�׻û �#�(JǽV�Uˬ��Y� ��
[y�Q�WmZ2��q���:,�:w3p�Ւ6�s�	niȠ)���'7��kS{F���
4���������M��a��oc[Qr�i���F�1�w�F1�+�7� J�j��hNgh��,�뵽������]�Xq􈤟�]Rf��0�w8�\/6ެQc���f�AA���y��;'+�z饔�n=�		ҭ��ڧwZ�����.�X��KZJ����ߪ�~��I���n�zb�W19����b�tF�J+�8{tء�V��c}*kͳ �3!']NH�6���ʉyU2�'��n������opy�{��U�g�j��Z�cc���)-Z.]�}�~��{,Y����rꜼ����S�X������ђ[d���9�����ҟT�/{_]���㥝���QY��g���YQ8m�oN�h\u}��}1����YV� ����F8����-�1y�V2=�Kל�	A�����gzd	�̃W�E>ʌ��&��A�U|���8��!�o�瞞h�W���`ю����Ù��Z���>5�W�
{3kll[>d̗Y��a���׿���$~���d��/~�d]W����}�ZBߥ�s�߾32���>nV��}�R�	�у#E]X��n��dG2	���X�ʻT�X2f��5��}��e��^���38R'�;k' �X�ʧ�K�~���,���>@Z�j��[߳�]'̟
ν�����e��h`^h:�↗���8;ծy�g�~f��J&���x�Q#��M�#�!COz�̡�>����de� ,�+c��7�/�Mݫ��;�R�� �+!���\�r�u2�ݓ� u:-+����d��a*�`.�&f`�ɻ�ܝ���q� ��fN�f�%F𺙔���xs�3�\��sq5-7.�����%��gH�vG���7/N��d���-�_N���ݱ��};ʰD��Χ:zk��㥇��G:DY����Fy9.Y�z=O���j|2��l�!o�\,�o˕�␁���N�5��R�rH���j�����[���PV�k{��*�˨�a������T�/��3�;����
n�y�C>�A
�U����71�fd����u���1�ڻ(oz%ʋ\����һ�6�������|�����X��H;�����O��T�j7\r�e�
��u���/]G<l�<��g�V����!#�~Ħ�o�:b޾�Y��5Mwc�a�Y�۟�ڭ�P�̏�����Y�6����,�=�Y�u��>�Mq�7�|XS\��[�X���z�򋸘{���/Z�r�����p O6C�I}��R<&+}�@C캅av�b���㻴����^W�͢5�W�~�+�DO���	@I�'�b�$���VT�n����yW�fou�1�zZ�g�r([�����FԄ(5���Z"�:Ц�2���eߪE/��'���Kj4�Is#1wt�8��=nr���Z�Zy�Cx��r��jɹ ��0C����`�)%ZO�V�R���������[���_.�9К����h����%��3%��s�n�0�j��З�;�<��-��=��$T�<�]�����Tb2�b��w�����w��V)Se���5{	V+�_f6�߭����P�=���&{;ˮ��z,�y���R��Q�TȰz��+_u`����g�v��E����O6g�9� i����2�h3�[>��Rs�<��˿]�'�����N�TDMHY6�s�������@����p7o�:譹Q=
��°븼�:<]��'���lD�}�������KEc��V�oy-8b��c'Mו�rl�M����5܋]������9@��+et�}�7G����H�>�.����Y�9Xy���7��*�{�&/���$�Z��Y��廋H���sV�gy��A�����U�BQv0/t�c�JK�$��]���	JEw�>�H�gfGP�5���\2�=\\�G�<��{�Wpb˘�8$��k�쏼����g��lh�t����sьl���iw�pi�� n�?O������,���c���X�?y����L�!�fAu����h�\S�1�ե��vo�%)vf>)Z��X��:�����v�;�����e�������]:�=�u��{-'�q��+dݷ\�'�S���=�>���*k�� ����W������)�,O{j'�93�|b�`L<\E��v�q���#�7��I�κ�XceOA[R*�*s�%Ot��R�c��Z��S.��e9Lc�Q������9��p,��K2����7�,;�С�8;��a��_P��Ł>��V��Q�nm��J��a W5��=1s�O���sHʎ�B��{�����{������<᲎���e{��}��瞀oi7������(��:�i�У��Ah�#��דp}){s�fڕ�4th_�}����Q�K'���q�W�F�/��%���㏇�=�DO�>9yʄ�1�Q.�a�C
����_w�Dw�s�V\�nKGg��<��H��~Nv����`�������@8�#~��'���^�l	��:�����2O��7u1�zR�u��R��2�<Øg9�I"��"}*D.����T��K}sB8螋�l{=糪�:���k=��$����v$L�o�cpv*U��6?W]����~���g�Y���ɹy*B�)^Ի(5�S��Ymk
���}P%uJ���QK���|oQI����t�׼�Ӽ�mWm�WY�6�\��5�uE�#�W���5ˊ�w��B�=���q��Z.uپx�*Yh9��Y˰t��naڵ���~�-���Ŭe���W���L	}�@yekM�;]1�68�;���=�k�tϾ���f�������p��(+��yp��ӬyU } xu�٬�q)G��nw��:��)&�
�J��+~}����W����4����c�fWH����N�B| ?x@�T�|W���A�aP�2}��=����B�UB�H�2�Ϥȋ�ޏdy���G*�ݰW�J=��Q�`6{���q���秆��c���1,׽}���%��m������(Sy�1pˠʿ�Wc4�$y{*{��n.4�1�OoUjrx�E��bz|��b$+�ߢ�ܗ�h9f$�n�;�%��V�/3�v#eU;�j�M1���ژz&�a�1O����Nt+��(��\�r��j��K���3�x^�Od�~�!L]�����h˺>�b�����{���"{��|�׃wX;0�+k5:�G��D\{f{i:�����AnU�b[w)��#�9��;��?P����:|XX��/⛮�n�U�����mI��w��u�W��r5�M����k������*[��IO���;6�wX2���#޹���{��F{��u�t �u�����Ӥ�m(cF��)MY���6v��ԩ}7��Δ���ֶ���-���B�]A��IA�b�!��iHQhS=�׶ԧ&�VG|�fd4�6�왮U����>������M��X�t�>�$�˙~�a��2`�ο4|8��:;��yH��rE��7ߍ{[5�$,�ٽ*��]�"�u?0;�}�>�땄�0uGLS�Jb�9
S��^(N�~��'iqm�h&�՗�w^��w_/X��٬��d�KW�1W�}&�K���j�~�_��!�}��dfY�3LПB䳙#=�V]̉�qX���|�.���xŇ�-��~���=��%�G�v{Ǫnd[U�+A	�:�Ż0�c�I���ʷf�8�U�F�>��=}�6�3Ǘ:��J�lvlD��m�=E���䆫��={��g5~١<@lȒ����:Uԅŋ�w]
������L�R��<�V���/OEP���	e�_��w4�IX��%�/գs'�(���1����&�z{Y/wr�s߶[�w�;}4�y�=�y@3N������K��Y�%��^���u�\�}љa�O5O��~ޥ:�2Cf�����qk�0h����)K�{Yt�|�½J�>����̃��4n|#W�0����hbk��\����f��*�����t:��'�,�Y�.(_R�xk��2��&�Ѽt��;�=�!B��}p�$�If���o��w�]�_V�=���)w�9*]R�8nm�����N��5��C�V�g�!Or�z��3V��E��;��J-�������(�S�pedV/@����WP�����sǠC��N���́��v�ʧ�j����q�+1m/��=�{&s÷5��HX��-�ç=����|��T��8�{��)�Ov]ҿ^�W����H�P���]�]0�Q�.3�ף����Zv.�'}����֫�%bL�a��,_S����<��Iv�	$ɕ�|�7~��|٩���>.~k���.�=ؙ;U�W����6KG֕L[�֗��h��¸G�}��� �ˎ��*��/��ʻK^~H��� *���*����k�:��ǀp�߱�Kjk]�
33˹��'��{�m�2z��GȠ���X����o���0���h�WӋT�O���u,_]��5J��?0dP�J���8o�=�E��~���*y�qS3�[pE��e׏���>m5T�b��:%��M�KF���T�����ntp��P|Q�(]��|���I� �њc�$6���J�i��"��5ѭ�U��� ����U�&���va�F&d�v�HAys��v��)!t�4yh�.���"�_�f�����v�ۉ�w3j�d+����e���F�)��跗z&F�wT<����5�����RC��>wҦM �߷h��/�sL�3��S=��빃4�o��/8ĳ���l������j����`��>��W��-۟���Q-���uy|�08U��ڔ	j�5s�VW��x����uS��i��7ii����yX3�[����!���+|���Nh�	T�95QҤ
��~��ڌ�R���3>�ʓ�pc�iCҸa��c��3;k<9�z��3���Wu��Ϸ���,>�]=��,Q����#Tl�c�@��xW3Uc�Lv�e���Lt���:����%�v�����|BE�?_E��In��ªio��=z����:LuQ� ���]n�]�'8���׉�`Ԉ��G���2�J/�c���O(���,ə�����B��ޕ��v����Hʨ�x�8-j�X=��u&��g�L�7����t H��g�Mo¶B�B�B�|v�M� Ÿ����Nބ�_ey'�s8on�Gy�מ��R|>�����N ��3�0��k����V\�?~�]�l�L�2Ts�M�qI+3j��m�LA;jE�m�2��厗����N��o���ܜ�頇�gγ���.7�AE(o�*�gH+�L���M�Q�tDD��麵���*����Ц [@.�s"?tp�lJߨ"g5�7_a�s�4����z��׽����,�@&���>����=�}w>\ح�Ȯ���Qx����3�)l��q�#?(~�v���R*����Y�����\|<�`t�>�&f��Ak���t}$E��\V}�dwX�p	U�Wz:�L���ؘ�mu���x$>s�Vp�_G0q[��#���N�R�p�5���0'痊g�[8��2l�ڐa�|��Dw G���Z}|&�(��
��hU�G���{,E�� ԝ��wz�u�Q�צ�R�(���uOP�>���}7��D�p�?�#�[�7���7�wm�S��z�.��V����� 5_EY�r�_������^�X������)��{����e����#t�Ǘ�]��"�^�A��ꄮ��y���50��T��^��%5[ţua����wۺoF���F�^�E��ܗ��<� =�g|�sԱ��Ni�8S��v���_����ʹ�w}=����_WbF��2�|��r�x��ͱ3
��|4�KKFL��1���]��;�r��$�����$��,���4C��U��]6)�&�T�FsU[��U�>���_f�4��s�HL&J�4
j�6�
��ʢ�E����������z�`!Kmiܩ�8k5�1�6.���罫�}Dm��x��,e��Y�r�|Op���5q-�t;�b��l�W$���&Kejuuf^�;�k����n5T���h"�-�6��ы=���*�/�.?�t��}T�u�HD�VÒ�\��[��Q���� �b��7�h��(C�~{�s|�1�@��w5��R]�2L�(��_���P��a�µ���ќ�c�A����W�랯n����"ߦ5���>Z>���
��+c�k��)��~�{:g������ ��	h�\,������־��><q;u=ev(�� %�⼸�\~��+���(���is}�#Nޛ�`�	~w�P���]��y��/2U�U���x���z@z�N<Ƅ^��k����( *�wBS�0a���DOo�����|-���G/7�������� �o��h��Q�O�M����F�0�SVٞ��̎��)�z��l`�,go�al�s�=��}�nc��Q��k6}�S���IU��ܫ �R���%�2���s��<�tۢ�M%�̔n�`��Y��=���1��_9c�:�[�7 �����q�坜f9��:a>|.�+Q��c2SGB��t|��Jː�u�"�i��%kR�:�VE�Y+7[cX��������T�������,�8��pl���#gF�t\�yg;��jN�⠳.�ȕ�jb� �m_TC6�������9)WK-M�w�q9K�������	��%��D��z'k���*���Z_07z��ꀗ-f�=��������%a�1�|��)v���G�.�])y2�:��������	ʲ��{I��,h��g����4���rs)�ʝ��F�ߩ�U%����o�>!�������޽]u�VY[iiT���M*��Ks�[yZ٤�b�]�xr 7��15s�3����56��[�9�6����U��̛�&�[LZΒ��q�
��4U����V�ZA��nwr�=��ىvDN���8)�Y��6���1[�ӗZ�T��F�u%������R��k/��#�V�S*&�mA�ڀ�N�A���oQ��FJ��ߍ�	�qq(.��lIX�\�ݰX�)˱sV���X��\�.���5^�X���](��*+��m���L�K<�o/v��8��].�r%�HoT�d��>�i�4۝WV��=�*�n��եs�Su���Yͷ���$4�w���w,�Ւ�K=N� e�Ҫ^R(䝒�c�,V�+U��c��i������;���-K��X�6��@��EI�5�[��x/4jt�%���d�S$�C	�I4KJ�M��M$�m��m���Z���Fo�Z�0k`'dZ��)Ivq�k��rأw�u3u���LI��J9IC��8��u[T���J��#)�V�V�:Auö\�A�`����f���9Y�jpu��e���i�P5/��� ;`�^���u�U���5Y�tWo~ѕ�,o*YK�ܦ��::4�O]��1���<ré	 �n�7x�Np-��3�ɑ�ѩV��7'�4>�û�.�PٺG1�\0�{M)1~Q��Z/��Y�gwe�RۢiehA�R��V�SG�y�;7�(���'i�ݢb�*�&ݬ�}JЗ/<��R��۳{��j*)�a�� lr�!#�p�������]�}�.��\Y;v&T5��N
4�]F�rW���Ĺs�{K�iw��q�5E�3u��n����g.q��)�ֈ���]ʊPH�0�S*��E��w(�D�b��6��SE1r�,(��8$��̨R(#����
�}�ȥv�I�������7F�����3��nP�W`äδ�������yxL[.��c��O�8�
t0�����ު�CYG����*�Wb4غN]X��fj�I�&�a�6���I�"�W�Vfj����;�C���"��ɮ-�p0���z��<O�2s7���Q��=�-��;�vo�D�L`�z�`u��H¡�2V>��g`�v(�i�����j���]d�ͨ��s��,J�R��W�hd�Q�����m�Pf2E��-0�����s௝��T�:�$�&�X}݈ó[�T�0 �9e���=Nͅ��ޜ}Ԋ�vg�Wʈ��w\#��ݩ�@�/ǃQ�Pzj3br��c��7��(�zZsoq]4�6W�ݷ{��}��>Բ���b$*�����pV���ƹD������VW����[�'�;q��'� �޳A� 1���f���)���O��ͯi*[����H��m{�����t�F:��/������F=�x.:��|�
^�2�����t;��������ƆOMJyr*D�^����'������05L^+�/^y �&#���>��vHQӂ8�z�ᙏ8TuO((��bs)�S6�L(~�5�"��R���1ma��^���팩�bWɒ%O��Zͧ���	x2�vx�Z��h���'~�Mt��={!_��(rd2���v)�0:��� և�xw�s�Uݘ�~��@��o)ni�z�17Y��>1V_����[�m��l���Q�Ӈd`�Ǔ����{��������R3F�Ġ2�f�(�R�/�m���Gf��O��^���6�\���|�u\���U�ɜ��Q(�j�G���Vyءw�*i*8s�����*9ɉ��=;�Y�w{[Ԃ
��V\���f��=��3��L���70�Y'm�]rI�`Y75�S��S���Mzۙ�?�p�wيO�t"�#�?lbϽ>��-=-7�ԨzPé�(*l�hЛg���[�*S޻#n��C0=�h��6U:/�ۃ��`/xJü@�tĠa��_p=�d�K��VeS���o���}�M�s��f����>��4s}�^�mٞ>�P�s���(o�i��k��G�ֆr�>�n](=�*[����)V�m�����L][��)Sn��ȓۜ�ٹ�|C���=��"�	���k���T t�s�ay����E�2���W;ɬ�乭�����lX(<�Ϲв����U��{�f�d����B����Oc�v��;�d�Ɋ��'?wz&4G�����	$:����YT!g�R�x:�ޞ��h?g˓�Ub��lY[b{/N���4��+"�}�ב���z�>��S���k!�dI9ծ�d�AQ��fHY�R��Au��a����ǻ��K������ᖻ3��=ץ��y5���}�d�3ދ���>�����besv�q&gT�|�B�$�,T�a>���IO�8��kG'h�v+t�CZ�{ Y�F�a{��ɜ1C��՝qf�%�]��K��:�.����X�]7;[��ٔ�\ʾ=��k�4ѻZ2o;�H���:�3�m/����3�ժ��{><f<�11Z�c�H�_�O��w]�������j.�eT Q����U�gk�y��2U1N�ͳ�5�e�o*����>�?���R��.�t{���2��ӗ./��;�꿠�˾2�[<$��=�hYU(/V:=�ޛ���0�}�w��.b�zX}3#F9��{�;��p�lS�S��a��܎
n��C����l�0
ΓґO�O�]����[3K���ٚ�)v �A���Tcg$�����^����{��G����S<��x�ʶV�a_u39��y=�{9��0G��MS�<��n<Y<����2�{6v�>$��p�WLnM�y�*���{&s} _.��a�(\tgP��h6�f�vQ��U'[ЕǼz`�O*�O��sc����1nǓ�Qd�0GNt�i�����=�AVuQO��	�Q�UѴk���g�:����}嬓uT��f��F��ĸ�b.�;ǟI��d*�^z|����zq'E���+߯�u��c�G�Y+mR�5�A�j���ua�]�X�Ĺ5��j˹m�i�5)\�6�Ӛeљ���{Z�A�(KT�i]���n��Ƒ		U�kx�F
n���ٚ�hC2�lom��m�lfe�+	̻Z�.���T�U����zS�\����n6��x����jCd̮��V��ڑ��^JY흏(�U�r@�KҰݓ�W^�F�z/�R�z��:�qB�p�~���v�{J6m{d�YGX�ʷrg$3�ee�����|��M�w'˻29�<�}��X���Zٞ�=�@j��~���/k=�����쌗�c��O����U_T�2�G{�*Z�hz&.��lV�/=4��J��$'/��̩���NΓ�������������Z^�|�V���Y
�H\�q���thY�4�l���ueYs6l�=�{���sE�W^Um�מK��g��Y%����I���Aa,�K�wMV������Wbi��S�9��/�;~�͍��^UT0%�}T�$DI<ǆ��~��pퟢc��di��ݰz�IS>���Ry��"������a,�5� ����_dM���{.�ȷ={NV,ۿ���?�%s�c�ϋI�~	���� �(9�:��>+:Fb���u0��׌�Y�G��w��}伹ԩ�:�M�iή'���S�����t8�������)�)V.����f�	G�L=�S2S�*�e>�+ŁY �0��uT��X��w]uwq�]��ƸH�t���۠AYA<��B���KH=B�V��U\a�V���P��N�ÃTw��w�=[�yur��+��R{�����ϔy=�O��~�s|�ԣ�� ��^-_mbHL�&��&7���2x[����ʏ���c��Y��F��Ң��aR�ag�;��%�}s^����11�>oZ��Hcl�޵�]�a*�&~�lAƶ$����N�X��ޙ��v��U6(�EY�W����O^Nx��Fϭ�}�����}�[���ا\��g��@/%�
'��;�O�L��6H^W�m�p��x.Ř�>.}0T��gү��S�n�%x��؉�&��X]M2 �^��f����V��܊�ߚ!�_g��`�>��P3���ճM�q`3릮�仼��l �J�Gf���r=�F����v��ӫ�NF�9��wl��5U�k��N��$=/�YC�]������2���0f�O�3��^���ϩ�$�Jwg��C�L��e#��+�&/J��5�1,�ͻ�R��ٻ�L`�C�r�FN��_[��|rQ�I�!�\?,޸�m��}��k�!�xʤ�ji�{'FQ̛;j=���;��)Z"�M:����9�eY�33���H�#}�¦�^�V{�ޫ�u�J�=*��cޖGM���Y.�_!�u�pm1;���䏳;���Mj���*�t�'n������fsk�J��x�+rk�ή����{�q����x���}re��g}3ˢ�8w��p�n3Ԣw���<1(|VӣW$g���{JW����K�dG�H��5^�c�P��C����p�A�l�}���z^_�ϗΒ&/�gs���y��}���c�.��n'3�<�H�K��n����w��0�WC�#j��\��W��;U}+8JwUz�x(���yJ���K ���z�s����pT�O�ںr�V�u�]��k��>z��ޢ�}��� o	/mGGzzRI���;�b&��w��L�g��9�.ݤdbUvr��^�=<tK��qZN�\��y�ˍe��n��,��}Q>)d��,řI��8:�}b�e��$�巾Ž}s��Qjz�<~��@��j��:�7�3��!XK�^3	x���R����o6�x�pp���Y�?=�"�I��9�0��UQo�c����~���g�J��$���>�>G���<N��ՠn�o2ϴN��(�����az\׵����v��L6�F_�v���S��@�l�u)��`�pia�kWM��J[��r*U������G����N���I/���͐�와夊�9nfq�\�����獙H�6A��i\zWk����y�}ƅٕ.W1I����d�3�!��=ܖS鰼|0_zU�MU���;/���l��_}���e�[�.x�f�{VU��_L��a�X�s�\�Ь��`YM\���x�p�5���i��W�u��>�S����;m��mO��`<n��#��.��;��v>���T@���;�5��<a�^�-!7�����^\ω�7k>t{�,G?9���Ƽ��������)�̔	�͚����Q�:3���בv}���U9䦏����/�efGl0�J�`��W���+ٓ";���{}��^�Dz���Y��#����:[���=>��^��w)�sx楳�'ýy�0-�h�,D�N�>T������1�MR;��������`��1�+P���|���|��Z����7�N/��e��������Ї\f;φ��'�#���'�����߁�>���S!�9&"ObTrg�}�.�F�����[����3�H4�qǒy&\��7��Tc�%r�~}{�޿����f��|cȕ����=����:}F�JnDq��X�޽'5���Dޠ9�8,�.Y�J��YnWc�;��YY3���!�J�!h?ɤ�o����]fnk��.�Y�Ō�.P�	��_qY�42�_��,
&�'q1t��$�L�%@1��l�hE��`&V�l��SѮ�!1��4�N�oĎ+�M��՟E,u]���Y[�|������������O����_l�?'ug��2�dꆂe`�DW%h�_uG��xLE����r����*'�| �����&Mػ���ks����e����n�?o5x�۬e�����0s�V�Ł}(|�9kn{�6%}�/Uؐy�h�����BF�I͔��O��^{���T�ُe0��������������}y�f�yL[�����\n�y%�V��(`�k����lTn9���+�2%/oR*s%Ԑ<�P�[���!�B����}i�Ǜ�KO�n*7#���� un������ȳ�/���u��eV2�M�ۀK7ɉ���#R��{��C�X����V�X1��y�{���6&G�o3�C�Y��&�`��Dk|��0*^T��7'v�zh��0VNX�����#l����V�v8�)���:!�]�Q��M�:ܩ�N�����^��Ć��h9��=kOFQ���g��N�u�����ً��v�u�zɞuܸZ�z$��w�����<�^NJ���e��3@�嵽[L���\�9;n�b�ܜ{���5�EV���h��e�{՗ι۔��:�\�>r�]>v���X[��ӻ�}x�;H{�Z��s�װ����
V�W�{t-O3J�:v������yR���㤜/خ��@F�I�L�>��/��o��W:��*�ېT���*�n�z&{?/f���@giV3&�ο~�0�A'��$�߬�u��|�',���x�~W;T��7?��]z����Q0>���r�Ϣ�KKEF�1��]"��[��<��Ƽ�=�,ب���.�ɝޞɘ��-��#���}�.���`��i��W�˓�W��X�/�H�<ʟe]|�����{�	��%��)���W�QOd�^�|���=��~d��
�A�Ν�W�U�{O�ߧ��̼�U7`��37B/�&f�GU��2���)Hu&N�7yV�xV˪��6r?�>�]F�$�K�Ǩz]� M{���/fv#h��i���5��z]����#�b�G�G<k��[���UMK��V�;���&v�P���!໗
�t� ��>�W2KT0���I��V8>g�}�N�Ě��<��v�Xc!Tz��pm�����^�g��j��G�dßq�6:����d���e�	ů�P���}��
�`�����/��l���6��vDWxj�J�e��]�N��Z�[6wS�VI� ���uq\��������F@�%��o��s���V�}R�������c���G��_�C$p�>�)_�yv<��_���U��a'{N��O�ƅ��3�{G-��0xrv�6�a,�ǻ���8Kڳj�pP�N��Iޞ^n�U{��qq�P��ٞj�Q�;���V���3~с��;e�G����R�_�w�g�k�F�����:���2c&*FoR3�\pܔ�+�Q���J�}ON���ﺪ5j�:/Y�=��F�ùb�L�f��4��~�=���۹zwJ�t�]�fJ�۞]�͓<эNN�������?z����p1�`��=�z��¦'�&qO��/�P4�Г��V��e]o�����^Y>�焼����>��~�����֙;�m�9�l����J�^�[��1\KF}�� �wؾ�����ԓ��f���U=�#�t�e�3��~K��5����!K����T�{��w�"���Ι�q�a��7脼��v.�FԨh��Â�=A��hT�By3o���]:���H&z�J�G;�?eŗWl:k�Ё�Q-��y#(��9;������C��d"�.�[9ro��T�d�9��W�yb�]���P�Ԋcmn�s$��J�2��_"i�ꠢ�՝L����ڝF�݌[d�� [�JAu;����X�#���
v솤�۫�{����ُ��x�4;RRzM�]Wv�}OWn��:ఎ�؟�'u�am͕n�U���d���]J��:����l����i�y<���bl�t���#謏xleS�Z*(���q;$X�Z�{.�Ij+7iH�v��D�^__h���d�O��>s������y������I���@$������� @�B I!��)!!$P ����I1��I �0 	�����������$�$����������@ O���g���Ӈ-}5����b�f��슥�1UWtvY�@����[��f��� V�b��h9��P��� 9M\�.&J�F�Pe��J��YM��t
���1���M�݆���D&Ar;�r��v�u�[V�n�N�nnE�G�j@�a�,c�VwL�ו���z�toj�I��Xzș��F��Ň"oe+In7V4�R�ª� �ݠۺ+H�r���RcxV�b���ͱ�5���(��7]�"��{b���RG�.i&�)[zr[�a�ܑ6(c"S5��5�*j�R���헍]l�x��˒+&`����5&�9sw1����GXE�� w��5�\r��&q���0��
����U�J�K����4S,V�6�d�����$NM �r�v��)�g���`���[�����=�u������e�sav˟�j�p�Ҟ�I*��u�1yu�t��@e&�Tyr��f��H\�(�r�p8�Z�oi��dŬБ��@�D��)".�e�e]�J�-�6��ݜa�����Q)YVw+B���K�eS������XSK:l!�Dhֺ�5�����.�\��YG0Iwq��Y��j^[�);�j���i�@R�'dW�&�n���l���?^�T���E*@�#�2�����k.�	kSV��Q]"&n%e��pb��$8��э���Ե7]�t�%dNmj��f����5	��u5݋B�3Ji�O��6�T��m��l�f�G7m-܂�V��B�YH�a'�Y.Kzh��5��Y�@J�Źw4Ɂ�r��)'�4V\zL�(�;t��\4ŚT�ڸr�х.����6�SN�@C5�5��l<�����&�.���9�-��Zq-zhfn�LJEYL=@�aV�[Ʈ��-�3r��x-IT��b%jӠo^c�0���]��hH@u���3�h�5�6�X��̤�ԫ4�5a�kR��ؠ�b�U�D�Yt�ah��[+���hU��5��W���\��4ӥszR�����xU�at��tv�:rkI��A�����/5`��'Vf�SXq)��6�,7LT�[ ��y�u�+q'A��͹��Jɓl-zi�Ǣ�b�����7�٢)T@��Μ�(�wE�0���~شɷ�K`4c�kt�`6p;�VK��ZO2�a�J��E������P۬�ݷ��H�`�wmB��t3��dk�B�Ř�T,m�F����nZ�zU�!6�Ŕr�Yt���
���K����7��vʋas ���{(���
�	Ҷ%��D�Y�tZ���ed��rͭZ��1ێeEk(�cm\9@lyX��VmH�ĢN��!T�̩���"W���Dja��@�y0�wX)ڕ��"5�۬���1R�ef0�
P{��CX+U�ݖ�d�bE�m@�l�7A���@�ԑx��CA4.g�r\��y����n]vUr��N1B�TRޛ�Q�(�؀�)i҆��`п`����[aIvE^X��h�i�j�J�M�0�j���Ǒ���Z�TGD�X�A;Glf�VݺA�4t�Pۊ��J]YVv�X��oS�)�.�t��*L�Z�˶�3��xɊ�Ǝ����w��1L[�j!J�+C�]�Zض���-��@­�F���'�SI��/.e�v�Ƌ�c�ť��,�u�\����
:h��П����r��U�Z�F�J��y��h����44����w!�R�7O �uFRц��Ռw�eT�aͫ�i���j�l��Y�`U�j�Yd��;�t1�`J��U�I%Yt�؎%B�(/jβ���Ɗ�b�A�E8��l�40���wk]�#�5�H"ДZM�-B<��c��0�	1VMuw@bd�rV�bl�M3�L���xF��?Z��To"���-��g��D���D\b \# N����9lҔ��D��aN5���щe9���r�����U��#�6��w�2l�X+	��Zuj�x��I��l���0E[$\�Fr�^5�i�Y�N�5U*z�X5I��l�Ad�ofVK�<����Ղf��DA�Ge)v	��:���ڣYW.�ɔ,,��r�2�Y@e"��51X�4���ٺ��݆��E<y[��AqnSZ�K��J`�kbV��*�k�D� ����73[�)��ǅ�&"�K�6�s,��/Dȡ����=tv�cJ@�H�EneK�J�?1�鐠ӹ��+�kfܤ�M�-m�!b�rU�W&31j�Ƣes$�&,t*]��A�N%��o�T�tn����K�Q�v�Ĭ6 -~�IfY�z��6l�b��`�h�Yd���,<n�	[���ذ� �m([4T[�/47��G�y�b)¿m�� ����LfcI伧\?�K�p���VY͂��Y�����vF���J�]��4�k40��3�n���%A�ݴ"��k܁kYX�ب�Չ�I�Q��kle`I9�܉��e2l���֫FMU��&,j���$�ӄ��̷w[5�&�ǳ.�6Ei��Z��B�`�U[/Lk`����ь�wr����˰_�M) %jݔ"��u��A[A㫐�����w�2� n�)L�DY�*�Gi)��5R��h���4��C����*M�Ȉ�d��0 0$#$��!@����  �D$$` BI @�$$��	"BI ?��?�� 	'�0z�M�� �"':���� "F�I�@ O��H@ O?�܄$���a������4�@ O�� 	'�O��^�@ O�� �~�C��g���ɧ���I����_��_$�%�@ N����b��L���#hD�{� � ���fO� Ā}��� �H�PBU�W�ݒ�(T��(*�v�(EH�TQEP()$UQ	 ���J�R�%$�%R����|ҕ ��U*"UQT�TRT�*�B����*�����	*�*��)I!%�H�����U��{��e���>�'�>�{�ꪥWڻ���^�����z�}.���K�5��{�J�!�{/{=�[RO�{�:��e�:��2ם�P)��w*��D9���;Z٭�U)Me<����EE%$ ���ݾ��Z�����������䯾ε����O{�]���hs+j��w�WM�b���}�����F+��f��}﯉��������O3Bo�y=vS-6��q�%(�yΟm�RE�D��J6o6P�ڽϏ�S�J�^�,�������t{ ���S�SF���n����j�i�3��{���T�л����I�;�Ƶ�\��ډ�e�y����a�tooJ�z��͕J:��*$��d(��H�@ $R�Q|��uz֭�ͭy��g�P(O;8�f��E����δ�;�"R�|Խ��/���ݛ��i{V�������y;�l��*(���T�|�)N�������My۷�{�JkOK7��-�l�fT�uޱΦ��k�(�����{���l�<zU��G3_{u[WqSi�iW�U):˽�HR�}��U}�m>peW[y��1��,������{����{�u}������N�-73]�UoO�U)}���o�{X�.��@B�kJ�Ԓ� �*�JD�[�����ʪ����=:�fK�n�xl�9u�i����S�ֵ͏����gL����(5����y�U��7��9��br�Ն�ﾐS>�����m�s�����*�����Y�'�n�[�RWF�uB�������}@{�������FŞ�q"J�������u)����5ko��O<�=�Q>�GN�5K��=�|x�����K�T�s�-���Hy�.�w��ka)$%JRK�>��Q(U*O|n�A�+R���kj���{z�}d4�9q,s�{���ޯ`ʵ#��=g�U�ם��r��]�{�٘yiv�^��ă��v������'"��m�{w��[mVӐ�V�J%T����k﻽���w�R�_^�w_G��\[�s�oq��|][n�����O{=��@�ҫ#/��]�����G�D�w����6۷��m�����m�}��*�尿���Z����T�H���*�RP
�e��m5k���m�[�wm��;I<��먏��K�����{��=(�뇡�-y�(�d{�;�kW�D���{ޞڂ���Uvg;��my�x�!1R�L@ hEO��T�   �?L"T�J�41ت���!����S��eUG�  OF�SL�H���G���I_��� ?��Aw1��h��}���ﾤ�~����>�G�:I$���{�I�I$��ӺI$����N�I'ww�N�I'ww��$�N��I�I:wt����O�f�n����������������{�����5|A>�m�|ռ��|pl@͉9�w�z��~���ݣ[�`zե0��4�k��JI*8T��v�'�$�6:�{�1u7 ẟ���f���eҕ��2���?�,,:1�����GXȪ5�e]n�o]&LY��7���(�D�6G!9�p��뱳0k;ڑ]��o$���0�Pak/�ȳ�Z���#��N&�.�3����{�x�d��i�Y�e��4��&��&#ܞ�Xr�O�'3�[��� ���0�X��7��83�my=�y�V9�=2d#&���K�?�,*�o�����
q�.�o���+rT�w��=�`&��_�;Id�o��o��Z�R2��Dv&N}��*�e�JAԐ�vA���l&���]mSa�&�۲�X�\vM�f�X�\��ַ4��'��%^aB���%�b�!F#X2���1c�(;,m֝.ouX��w;���3E���]���Z��Q�C��L�K.�����ܧd���(���|�s>4*�Z�a���`���3�|��w^�C�z��{�w$x<G��g����\`�;Q�y!媴!�,?�G��t)�6~��r��I��k�N�w�2�`�P�b�Ж�ӄ�Y,ҫ[�- T_���c-�3����V��(�W�`SGL�d̤<+�Ow��KX�i~�+�{L���б�B}���;m�.@�5�/6]��;.�3'v�09&;��X�V!���M�����b�aSWp�ݤ�Q��b��G�YC��Dg��EU����XD�%J�HuwS�B��?;f�'��ւ�Q��l[ѭ�T�hg>��fl��E.Ƒ��F,�T�/qSj�:)]����sY�2}��(e0�RmV�78'�)���"D7(L'�
BU��Q,	��E�Sk%���{u�r��$�I@ݜ��#�]1%)Xn�w؆i�u�������$gpM��P�X�ȗ�x4��i�+��o�[���J����
h<�2�~/�ּ�ƞ٨�����&�Td�k��^Ӕm!�ml]pN�N��ӥ���ȦfL��D�o$tK���)�wR��$i����	;�𙌩���&͠���hO+UI�Y�I�غ��7��.��
�2f,׹�0�e%t�@l���ϑ+��a׼3���^ �
�:������������8P��8wh���5�-��eh;�7Y{1U���a���	wb�����(?f���x�I���������JN���n����Q�w����]x�?�ރ1��ے燭�\)ĆCL���뜪ϋ��/��v+��	�Wh���.7�[�_ �.� SD���U�@�C��=��ғp���5�u�z�=7���Ȩ�1�����eᶵD6y͋�;$�ݸz��X��g=x���i��Wn*��Xw?r���V�9D��v�����4��K�e�X�H�E�bl��GB��|4b]N4z>)72z�a����jIY��9Vͅn�6[�� �[�3�nD$43�
b�-����Z�naX��L��f[����b<�ʗEY6h=jNћ1j�a�=,:U��`���ʻnĢ��ש\�`-k�v��K���,ۃc�&��ه$���M��x7�g��1sL:��f�I��&p�#�v��N$fe�=JM�\Y�%뽱a��A*�&i���N�!�F&�V�Fn�wu������E�C}��g_�wq�?q��]f�<���k6U�j�7!Uah�׫Wb
�i��ɩtһ{��5�����5��:/���Ffcָ�q3Z=+տV�Z���u��=Þ@��,��
��C��8�S$�WA�����V��zE�5��!�I�N�ٗr��:�EFMdN=��#e|Ovp��U5��V��nk�B�\v�N(�+0���B)V&S��$ɯla4v�$un��(�X^ܒ��@{'�X�x�Q�`͸"�N�'��̲�;�`=����P����sz\�aE��Բ�mD�����c� z��ԄрU�w�X�0�,�&®hɶ��}�v9a:/f�e�EQ0ɮ���'~aXs8D���׉�G���Ƃ��N8{�E��cAr׻�W�� ٲ"p̯;{������ĳ� ����뻞����0�M�כ�o��Rtt
}�*�_�t�U�͕$ܞ��T�;��y���t4d�A�޷��'�Nפ;�=�dg�����82V]p���W�+o(�͡S��;T�{:f��͒`z�x���s>|�R��<�,�:�퇂��@��D�k*M6����d$�u��ٛ�͚MW�S���q�ix!�DLÛB;wi�rJ�,.�%{M[
��N;L[�5�fP���י�D�9J�p8��72ǚa��%��x�c�װ�,��h7�^�Ʊ��]�4�ͩzrj��$ԩ�]i����jK��^���C�9x��h�ӌrH�.^�\9�j�&?�X�]i�oj��␬����N!ӄ�3N+��m�_a�CB��x�h�f �w+2�&�l��n��"
6-w�����0̀���PP�u��!�
Ee�	!��K�5hl���E[ۻ������^s1��ۖ��kM��3�i�(��z%��+u���6#�lk�fړR�2����������QL��,,��E�ё�o�nx�ڣuD}h������.rX>>S��*������ʷ��v�Bq%r���6�[9Ks0c;]N�p
��RB��]!Π4�Y���{�������"�� �F];��?8"��y�	W܁0���e�wA���n[�14i��:ë��4ar���cE�-r3��s&)���L�7k!�-�ˁu���c���c��y��16P�hQv����K��{�`�7�)ڡ�ol�#�h�a��xFrD�i�=�����[��G�x(A�����3N9W9c9�0Q�˧��p�U�&�ԝ����R��}Bt1�8�O˹S��EW.�`�F�Ø;E{З�<h��Ƽ��n^�zI̧���PI���~ڻDp�#��Y7�/owx���tt��'��\��9��y���x�|�Ø�Wz�^�T���41�Q�]�GT`Pm;c�	ʙw$� �y[�j�4ʍ�;�k��q��'���v9
`�`~�'l��6��*W�3�խ�Q�m��D����e�a̓7M����P��IIW%a++�K�P#�=�e��B%_
{b��V�������5����u=�wN@�l��7�0��ܵ1�/s��#-?����t��U���
o� �ǔt+Ӧ5��lVNo��+Ʒ�L��e������p�p���η(��V�����̏
`il�e�:ґ��B���+�n+�Į��ok���c�� ҺRbM�-F���F��=�jy�HWqבp"�,�n>�qm�VH{9��X�+C�=������]�7���秈�r��:�|�@{7n�I�t�".�P�@�U��Laɤ��,:{mZn�3)�Mk�R�����#Nˈ�"<�t(�a�ħ���rI^�!+����G�%��f+mFC!�n�ᏹ��ع�,
&��r�`�4�j�6ۭǉTnݫ�!��r(�ߊ�ܑ`�r�ܘ�1�Y<正�����-U��L�SiH�j��uShG�c��&Ӱ!;��z�&a��s�1��&R7v�;/�G��id(��Ô�񾓎�Q=�����d��J���Z9��K���*z�X�
���w�ΫF��].6�ͩ�i�v�ό+������y�=ۧ��)",eє&`�(Tب~[:n8uz��y��w����BJ$ގ�C�4nS�8���-ف��U�ۜE���Plà����au�.f׵��n&T=�n�uƗӱb��+݄���-�S��7�e!��.���\#���f��u���i�����3�5(�r������/`Ȃݡ�8\�Ž���R�g+x���׼˭Ƴ;Vf9��'���S��F��r
ē�l�ͧ%+��NՐ7�a(m���@oSq���wn����N1�.�-��2QטQ���7(,�$����Hk9���� Jv`	r�mЇ|�L�".vb͢x��l'S0��+FB�G�����`^'s8�эC�E-�T�%Mn`��Y+l�xu�WˁQ���v�F����`f���P��Ms8^�&p��4�Ƞ&�"(�^����I���+����m�d~��$�k���'7N�P��tK�����`#)m�n��4l��pT�i��Q�2qu�i�;Z���e�=F���2e�0k��e/��}�Hq�\��g����J����vA����$��\	SAɔ�p�+cʦ]��w�&*^B�[�
�nU���z�)S��ڼ�h�Q;dԧ��e����@J� ˳���h�I�:�(�(�&𵔉��rD�bSs���r����q�v�[17��N\��(�Ի��O��X�O���.G���M�TBo�3��}{3O�`�d��7ݙ�(@��u�1�۶��Y��&e+):��6h�1]%�0,����f��1�]���ӞO�ay
1$ʜ9�Qr��>�{3Z��0b�'�[��T:����1 L���}6]	z�8Jx �ȹ�.4�eJ72���[,���Y�%�'-���Pr�/^�ȟ�ۧ��h(�A�*�+�(~t�:r水��Zl�+X�xh ��.���x�(h�>�w�h����VXM��}�?���M9��=NNE��5�a��!$o4u��n��zE���]\���o����r>:�jSt,�*�Q���n�	�eHl`�nA����T�����V���rb�-�AN��sNI�G�*e2�\�/�VDed�[K���T�\�h�v���-^i);f3bb���M9���SIRy�&�¦;�]H[�'+�!b�gwvr]�i�Zm3���2e�N��4l�+!���!�3�7��t=�ιJ���v��5;�63Lz7gf^�իY���&�̘�e������Cr����4{�v���Y��D�O(�?`�Wb���d!M[ՠIB&�j<Zm�7�z�f��E5=׌��	��<*HM��imqsP���'t��Ic��f��-��'J�-����
4����L9j��%XZ
����%� 7��P�E[J�y�3���*0��s��$��v�y��}�Zs4�!{�KŃs$F�����&f0�tcm�q��W*���l����~=d�
�ą�c~��]4�Vő�'��׍�ˆðJB�{�ŭ�s�o;��P�qsz�2T�?ѣh�Т�Ur��p6�U2���E�@ی*Ć1�(�i��I`����13(l��;,}���o)�Y%�&����x��77�-J�x�aw�r�{�U��M�8��fJU˘nv�X���ɓ�ڞ*�\�4�:}�,��ї�d��ZՉ���<���d,f�[����.�¶#�z��j
`�S6�˅����ƸL�e�M�	N��EJ�`��F�O2T"�Xdn�e,�n�Q�B9v�嵒����p(øZÃ*x:>Ɂ��d�����#`��k�}ѺqU"+�;7�ѵ���q��j�K�F=�뷆������Pِ�!�� ���1
S�0��j�I�֟w�f�dv|��pK=c��kOF=������F�e�͞p՜���r�O��z��:wk)��*!�A�dPR61͗)��x�~��x!wb�ǡ@�o�
�I�ڹ��=��ܗM��<���r2ұsw��i�Ǻ�F��ժ	K�.��2�[V�Z�\�PE�K�ï���l�%��Usj�7�/az�6v<��W����iFK�!�;F�W7V7��p��9ߎ��)*9�6��3�0x����� \|q$�y�维gkc�`�!��;4/�2'���Dz�.���l��ҏ���eӼ��61�{�F� ����EBfUqʵ������n��^@u����Wn��J�m�Q���tSr*x�i{xj���6��xk����W��ؘ=�� ����.��@�������{W �L��(��OX�]����9��D�!
����k|*W7o;x�+2ȋ;���r���Xyl���ƻ�:Qن)C�w�
�lr�f�zӰ.��]�Qס��5X5}��	�՛���;µ�+����mc��%&x=�R:�����p�;�Xso�<��ˎ1C���i7�ұ&�4��ˌ��4[��)�Pn�Ә-�7��C�A��bkt�M�6ږ�o�����;J鴶˃x�B�D�S���ꙇff2�Z�P����GXL�Ե{/�����NjY�	��t���D<a8�m�`[
��x
<fgS�K>7p'7Sh�YBl�No- k�򙶰%���������f�`�^7���=Zq���Ƥ؇�[�a���Ҕ☧F�f�Y�rots��c5��x^���L�T����]��Y��@5�v��^��	�@;V]VE���!��W6jn-�2rf�bٕ�Q�y�m�
`���h�8�u�>�M=���Դ�>ss�c��I��ظ�J;��(;˞H�f77d�rܙ0��1�p�/�v�^�/H������3;�h�<+�]����<F��2��	�S�a��]�-�L$�:е�y��eX)~��a6�v��cR��]�Y&���;�>��~חW3&�ocV����ȼO�,�=���Á-�}��2(V(�k�D��IM�E@���\aT D�\�A�v�����6�ܯ*D�@7<ٵ�����ɲ,鉝��r�䂁T�cK���Ԗ�*���J�UU�H�U�ʠ2�UT�V.P�eU�%�6h�4EnJ�\�#��lq�l!E�F�sq�q�"����Jm)�;&�%��%��Rel:Q�P�Yz	��,�l�˷�)�ş V�gq�0�l�M�6��G#�q���=�5/�0^yKn�X��Yv�+�-h��r�l@��T,v��0�jM�^U�c�Nب�󓤄M�9Zm:�d��Z��砸��w��h2�a�Ն�ܝe���2{:rݺ���
v{]�F�gc8Ɨ��/P�oQaF��m�,t��Bk�3K\��a�{F q��Li�W�0]������1 ,�Z���n���3{��G;+˷*U�	Kl&j�pge�Z.%�����^�.��1i5�)�l�, ��2ݠ��
�s�q�;�uOkh�k�!f,X���LQ̨YK1�p�k]�Yt԰�k�U�F�v��Xs�hyt�3�F^6�!�5A&�����R�K�x-/���u�#�i�Ic�P�Ħ���9��6K �6�ّ��^9-����*�O8A���P�]���nz���_!Oh���yɯlj�ט:�Ǝ�G0�	�q�틛�N�e���g8�#(��.�q���c�qTۙ5GU���q���SGg�=�����4`��4�-t\�`S�4\�ׇ���;���v[n�bۭIc	����XR��ɣ�n��Y���q���Ҡd!�b�V���%�8,��Jm���k-��	��K�cnJ�D	��Z�chtŸv��9f��4b�Q��gG�����R5Kz���v��`�v��Ksa��η�(.���S{:uq3�*�mn✳5��9.Hk͕�d���iR�]�Z;@b{f��Gf�L��Q�T����$6�נ�wPl�н����i���]�(CJ����f��刘�]8bْ.���L�U�f��r�1��X��nw:���D��KΞ�0q�r��pud�O�F �pn ���鱷\�y�X��Q^�AE��!5um1\lh�!�n�z�w��d�7��9㉵ƈ +��۫���4yvY�al�[�$������ �'e�ב��f�ˢ]�4Zsf�6�V4��l78�dG�c3ڷ
c�C�nx��cun����۳�G6�%���7���ћ.���V:�.�LM+1��P�ld�;��1�޺�l���Fp����:���-k���p�ۮ�Ộ,�-�\Wb#+�H1�̨��+	�.��Qn��%݈���ȅ���q��\#t&ي(�/Fg�(�(����6�7GOVcB����Keq�L�\��銦:g����f�'E�Xv�C�ʫ��1��C�\�h�"�;ZM9Y�U�^v6�:镥���`1�4c��^���\�4�79	�R�70=P��@�㮎m&:�^|q�Nwcg�F\��J�(�p�Ef��)$���v<��p��(��R;�ZM`I{m�ڴ%��,�/In��g- �u�e��C:�طXh�5p�v����7m�Y%����Ƀ��6�1�)��*и�� J�����s[�����nS�gC�uĢ=�g�����&b����Dhbl5��9��l����8���!,<�nn�`��d�6��q ��6b�ڥ�In�W:iK�ls���ݖ���˕��m	�Ye	S]ٻ��á��rJx�9]�3#rܬ��tnth�%Nw	f9��$h.��rnÑv�9�t�ط<��kq��h�Ѹ([�:�:�[���c�p�*��I���]�.�P��sv��	B�[�a͸���3@6P0���T63Eijk������<z�H�\i�aW7Q`\�3�XK	�]��e��x�hUaa�iq��$ذ�(�j�뵃m���D5�7l	�BܻB�ˌ��J]��2[��p������k�p��7'#m;��'���m�;�m1�IC<�ӳʆݍ�Yt��]��GQtc�ִ���{r]� r�L���w�ЦNK���+�94H�q�p��НpM�%���Z�!��fK� @5�<^îd�pŔ��r�Q�i{f�Ic[��wn��g�'^z�����ۊ�3�@ι4n�F�`Z�4�!.�Jɡ�e\�6���s�����,��&Þ:Iu�\��z��|`8M�v�+����s�㢰2�b��n�lzʻ��\�5mۧ$�{u�r5��v�k<^w�P��ûqn����y�z��.��f�f�B�zl��pY�(�%�SEXg�R�:�8v�aܗ'�2�ۓ�q�v����엍����8dH�1�5݅R4-Z��)�<:��!Wkp@q�3+bU�Bi5�K+��='Wf�^8;GB��]�����f�1FU�fK�2�����w�V����%�Ϟ�s�t�ut3	��7i�;��ѻ��:�6�r���f�\8��ݑ�Z�'H�O`����Cp۔�9�ˍ���[�N����ی����ݮ��)e��[7��k��st��i��8��Xu���n�Z@�4\:]�A���n�2�]NF,�v�q��H�r�V��ZY��3&
�!;�w���	q�Q��Ǻ���-e����PBX͊�Ƃ[�`�@U��܌Oe����h&���Q\�թ4aViJ����(�a.������ƭY+\=��l�Ի ��62�k�@�T{���{J�mv0�
Rf�Ƕ��1:䅼Lpmx1��X�� Xk��e���˼��Vgo9�n#�cZ�!n{]���{0H!CZe�pr��z��6��g� �[oGd0�M��ӽ&5�K'\��n9�{;N�wF��Js�����=��81��jܻ�˹V$�C�mK3K�̧��)��glv���@<���rl7��P��tl&�����>9*�۶�A�.K�
P�(�u�Ki)o-��l�j��#z65(e]x�����Ɔv�U�	���ɹ$^4�0�FV�8S�ks��g�1[v:�)͛d@�:mz��%u�%c�]��!Tp�n];��k8�{(�xNgM���Wi���2�۱Lɻa����=N	��n^�eJ:�xL����،��`��J:�.е7� 	�Y�$�PY@���@� sZ� �n4��{7k����`�$:k,�0fL�G\��ƺT��	h�b�i�=��<eph��2�A� Sne�n��3s==�����bhƍ�t�nu�8�>K�l.����t�fs���ո��©��P��aA�����YK'[���������F�Lu�9�mֺ�$I�:�%Vg��w\pnĐ�#b��u�0����\�=6ܖ�M�N+����$��mm�Uń,"�˚❂ɆD��ڲ֚-&�;�:I��<���Z����'nH�r�ӂ�v��l���I.$u���ej�s��G�x1]�ݥ�g�#`Y��`ƪ3J�PԺ�[�9�/V��K9�;>�6�m�W+�n�r�<�b�ô��V=X!3�k�m�1��kqX3g�]��͉���Ye�	^���ReƇ��S��\hgm��.�p����܇5u͔��׵������h��4��x�iӺ��ӫL�:���)��K��GMHXP]�
�4���n�Dnc����ծ�������Q�9{�,#���M�q�
�8�k��q�%��7\���=�D���YH�iN5�,�d��T��t���meD�3jyacۨ�r��@��ƞ-�A�w\��c���l,�;u��`nLn ��E�\F%wS�gp�;\Y��k�3�z�@�8mvwc�|y�E��H�] pF\ˮVW�Y��Wk�RX9�03V1^q��A�k�6�ku��xr�nER�-���!ٽ����H�YZ��K��f&���⦱8ٳ����n�!nwUoq1
�Zn��<捷f{p2H�i���gx�.*���긘] �^㶜gÍ��s�� T�F�![�	�kq�<3�(\�,:Q���N���2�a[���k 75�#
k�aU� �bFh�� kl��lonN��g�c'Rz]nc�lb�C�<����<���Q`��h�r��BR�.ռJ�f&(���/!����QMZI��v��9랢�ȝd#1s�{ �fn ��K�ݚ�1�����vY�w%[<!դ�)kh���h�����Yf!��(��Œ�v̫�vnrGk(��'��vC�l���эC��ptu�3s<�GB�n@�Y��xJX�/fY�Y9���se<��9�x1�</kp�d{]Y�j7%ѺR�@K��I�Y�G9�vkA�e�r��\�^�n4�\ 	�d�\��'n��\E�طq�s��@"K�̩+�� Yj&�Į,k��<�Ԫ�<�����	v^�z��\'��۵�F)庹n͏=�rҋ���60΋��1��£�؛#�rn��������ܐ����3]6�TF+�"FV	�,�&��+���Z����0BWa�&��v`�競ݎɮDް ��5qy�p^��]fH\���Z��c��ϑS�s���`�7CF�R�����HR�1N�Ke�8�q���ɶ⑵�!+�u,S[�Bn�=(��Wa7q��P�a����3�.�э�	��d�_cg.:KC���ɏ^vp�N��/\gwk�q.�R��Eyѳ;4������Z�&z�vi�ݥ	m�&��wn��ɜ���h��\XVWR,�4s�Ŋ[��ӓjv���t�qe#'.5�/&ss�Y��y�؜<�7!�e����%a+7G7C�lz�l�lu�FUt��GDm&�+�e&��n�r�%B[m�2�RR�$�VF��5��֒ͬ��(j��-�f3R��
WM5ɶC\���=�#�l�lp8�F�-GA�/c�͇qe����Z{hZP��B�S�zN�Iӻ��:O�߽�Ӥ��wt�:N	�$�;��t����ΒI'wq'��t���I't���t�:@�N��;�;��t	�t�;�t��ӂI�N��$���N���:t�;���I�8$�t�8:N�ӡ�������?
y����0��-�qRI����v���ľ����.�C\�;�~ȕo1
�l�m��i�
`50 ��i����]޺~E��A=�6�a�)�nC��Q��Y1�f�U����>�l��4t{~V0��on�Χ�<{'��VD4��EA[��4�l���p�gm������D�ܫ���N���˗�|�V+O���5������}'2n�<���P�����P�t0�)���2�6I#�>���f�Vf�$�dS���������!F��6��tekXC��*�e²<�ń�Ylm����o׻��\V��Qy*%�gn�a^/����~,G�ڦ��Ej��Վ\�&uE�k`F�h3(M�1_�s5�3�};��2�7j��'�g�d��1Z~���{�Ի����OeƏU:��iњ����J�@>��P	ZB�(�}��mz�{ܶ����<f�R^ؠ�	��ݨ�[X���P~�
i��.4��0�F��u*���ݴ�&��C"F�	��Q�����&V����$��T���4�aۺ�͹�"VI[�Y��a�����2݇
ۋ���j(s[���t��s�-�m&��=�7��Vң�O�+dNU��f)Q�%�`pQٹ�]��e�ݠ3�3<f5�!�	ɺ#q)����	ZX�-��R_�c ɼר�G���x��7ciӶs��F����c��:���-�����+�4�d���r������]{!�t\��sz�z���q�ke�&ѝ����ұN�Q�:��$���k�8�.Ƨ2����YR�L�u�-��#e�'Ug�!垃e���.�����T?ѐ=�>̹ͅ�lJp�X�o(m��^����Ad ����5WF�hlx�>���W�iڊ�(�;6��ՐC ̝�tTX��}��Ѝ�=������/\gӵ��'a�C0�d�u��F�؃Wr������x��Z΅�"i�����/�[�K,��Icm��Dk�"��x{K��tuЖ�02Si&T!��M-u��:3I�~�~�a�3#� f��f��h^3��w'lE銻[��T��wB��MH�h�u~�6�ˍ�w��xwT^�pg'.�}~��C���e�d�Fb"g'6��N�]-^�nۯ],��z��϶E׆'I�5�ˆ��+XP�2��ő�76����}�X5��߽��;���~����l�2�l�p�ت�l�wVNт�����^��4����H�{0�(�I�PA�`Iz���J��z��œ
�S��@ŷp#�n�["ZS�g�֏X�F�}��OP{��<�f��f��lj�I-�?Jә�|�10
t��o^3��V5�����x=��ڌ٦�j�ً�|�ڽ���J�z8|3���kgn�b�N��m����`�v�zm�!{WY�vf;_�XL�fd��#�Ⱀo�!��y��[�H4�nW�&��&��C���،>;�0�j? ��f��˚�&&����j�MPЄ��! �) �J����3�G�PS���;jƣ^4I���>���2G����~���շ6��pT�jO��cdN��J���e�L^��t�-i�KE8�pu�F#qc�9/|e��6��ph��fvvvLN�Fia����8Z��N/3׫E"ζ�f�f���s3�鴥��Q+���?_Q�7�V-2�GC58�~���ifԊ��.�fw��{�D�&�,u����%A��M�u;���\����aոP�\��0z��P��;1Q��H�%(�^�?u�xk���&�پ�K�u{}>l��=.�=��2g�.g���M9�q��ү�T�9~���Jw��өo�<��A�!�D K��@�X"��������3��{��;�&�T�� ?/�Ϋjy{9�z�V����k�_�b�7��vZ�3���U����z���w4@H0@p�:�������o|��3����>Z�cmÁflq�STԵ�n�5llv{=�3E4�I0Rj�����R���[�`��R��	
��\흵�M��#X��O1/��;-��[)Kwg��y�c��w�s.h.�X�i�a����z�G%6��W���ŀX��c��c�P�[�`H���A����L������e�O��pg�s3�B��~�.��H˿;�Tzc�J"X�⃍�x����!e�	i^�w{��YL$�pQH��U3G%�c�P�I�xn9��WWԖK!��d���n�8왤H|��Jt[�����M��S�lm-ʪA��E�t��[�z�ԟȢY7y�n�;���&�S�k��w�U�[��ǊLVz��O md7^(p�+��%�����iuZٍn7w?e�����8��I� 8Q�b��1ĮU��S/n_x&�����iq4矌��tM��ܛ������f3F�U��nz����q�k��8|yͣ��˼; %����V�׏d��^��H��Q��T�%n7�Bt9	 <���vH�j�.%��|k\�-Z%4�n���A�����٨I6��
͊����7��5��~�3�cT����?Q�ә�"��[0D�Ű�����P��>SJ�C�3r�f�P����˶��Wv8��Er��*/.�j'%n;����ԚJ��i�0�'ej��30��}w#��-]�wc��Y;L���.��!�v����	����'*�"��v���k'>��0�cm��v�[Z�m�/�Z�~��f�#�����d��N�{��^K���.�x�[@{9v-�KC\2ϝc��ȡ�%�V-��a@M6�'�EԒ�9{Ƒ:+���;yf��
��9{uw���O�{^�p}���#�q]H��=vsf�񍻟<X��ÙJ����F0A��E7�/k�H/N����7�XXY�k�}&�mt���bi��fVs�E⾓�?[���m�ey���+;�r#O�`��cM6�x|�;���޷D�qq���kУr`Nb�m$�� �1�d�n�m]/8xN����ڽ�nݕ�Nwg�щi��;f����0g�T�>�L�إ8Mm!��f���5k2~9>ɏ �n0sbZg��	"Jd��YW�}>�k��;�w�F(��t������R9�=���y����1�
W�,�y{�9{�����L����O���p\{���5��$���C�gP��w@��kT �;{C~:��7�2V��Y���w��D���gZ��x"S$�q$z���v�ѳ���ߒL���Tڙ<v��g �7�*ɳ-Yr�"���٣}��R0]�m���d=�.t^��+�QQ��X�p��,��~�=�e?���` ��(�( RoN�u�ݚ2�pd���Ml�@�f�������5��b$O�Ү�����V���u�:^�t"(%�8���;{"�vd�����Q]0k�E%M4�DꩦeɌ�F���s�`,�k{CMrP(Bօ����<�[��S�Ź0ܸ�� �s�탲O=��޵>ݲ�M�]v3М�R�2Y�P�a:u��d�'���Ӿ��87�9�]�|��Lol�)��-C˦�(`�о,�n)Mx�MQW^�
�ԓgKWI�l��������ߟ�k.�o�(�^��Kڽ]�El/ٹN[���A���^�p` 8n~���/0 �ٚ�$Л�u�7�����~[���*��ո�
6u�9�ٷ,v^�92��a��bc^f���C��{l��X[(�ؠ❽���0J[9X)���`��͖w<���i$�`+�[#3jn߻�I��`����X^��ŗ�ab3��(:^�Kr��o-��o?F�Z�Ox�\�����
	p)�^ƏRUB1eee�I��Z}G$��=����U4�ڦ�z���uޖls,�8��ޛD��K�d�7Y0hی��#i� X�֏��d-�ZK�I�����M/zs'�Pi�~>T��������Ʈ�����0n?Bo���"��[U�L��E��G;��.�/T��w.�g�ce�Q��q���:�������\��αӢ�p�N��ɛ2��-����J�ݮ��O��W9}n��3�A�/�L��{�8�]��ZM�c�/8qE�[l�c�������፿��3n��ٙ�C/����W9�on��Q��n�&�P~ű�}pƻ�lLȩ*4�	(����m��-ʹ�v�]���iK��V��nT�J|���Ｋ�c�R�>isWg������5���5����{�'Bg ��*q������ sP��ZUj�(�j٘���F7ϥq9�΃��BCD�/�u��W��w���=�ǳ��n�}����<ښ���{*J�~�p��N
��MU�r
mT�,��u��֫ğ�i������z�.�^����V�|ϙ�|O+ ����7���)��d%�FM��䧨|7242��L����HҪz��gr��)��U�ߟ�C0z�w������3���=�6�`T�R������u�|�$`��'��^kTe�:v�u�^��jfO{���Z�T��{�{��5K8��c���X���/Rךn�5αn�k���B��G�8�IM��]�Y~/=�a/Aњpg�$�/^��`ra��D�7���\vȏ���ۡ�k�try�/<�A�X��Ǆ�Э��5�l�C�=��׈�vt����k������Z$ƪ_V�N����G���+����8���mk���ή{Np��[�N�7��zOwpX;�eeV6o� I���^k�E������}&�ӆP� ��R1Fg������xG��-�[�G�ۿM���N����Η��wb�T�N]���&��ʖ�c�	�3#j�3q��@E�4��
V��W��ob;uj�K���g:�Ü]i�'il��|��9̯$��9��zX��wm�O���V����0:r���p����̡9TF��f_�w)ߞ�Qs2y�F�Im��:�tl��b�3ek���zk�V��<��~�3�q˩��PDQh�;8�Y��3Ϊv���h���u����t"��n�/ M��W�����un�Y^���}/r����y�9~�;�cO��(0�!<>�0�vbp6��'}��ݛW���],]������"'��h��q��.�cq�aũ70<�C�6���3���*:z�f(ōܪ;U5wS�/a���G�S���ל�=�z(f!�S�����݋Y.
���1�wzb��|\�BO�h��g�{+��%���*Ѹ��ޯ]ں�%}���[��ϰx	�h_/����j�ǘ�`��k}�������]s�-�Ւ�V��^�n(_%�����1p޴:a�d�3?L��D��|��g��Z�_��O���lhŽ>�9�[]�9��*,�6V�^��$y�;)��=�c�H7�^��-
J��Y:X���Gp����K*5�ŭ���Cpi��/��&����'��w�|���l�5��c}^}�&,�ll1���>�뫇�;�uaÄRe�P�R���q�fuf�t��؅Q{���5�-��*j�m�����R�U�w����Tݫ9��^��D���� X>��(d�h�0tU��U��54�k���RN��1Q%���lG1��=l2�z��nk��ܹ�tm-�%�<����y�����5��qeS�Uv�ȓ���5���g��j���N�e�9ߕ6�<,]��^�`�@PPŻwst�c%}K�7Lj�qq�Q��\J9F�D��1do}���;<}�ycb�C8v���W�����E�CM�kƌ���ň�e+c��zc����Ʉ���K�%x�I��B��s5H+w���+q�����&4s|�ppq$�$&������{� }������߶{�d�b���6�O�z����V��V0�q�Ȃ��Փ��t��܋�����>17g����*�Z:-͗ CGY�����cH��˞���4�J��[\ɤ2��m��9����ۭ�2�JA�n-n���\��n"^;p=pg��{�q�-�\�h��/2d���}���ye�!!��9օ���H���ٮBׇ@m&�-� �L�X͋2���7`XKH�4��٣����7'��\��78m�d�Y/<vx4%��.�B�K��[E��ۓ���qi,����q�Jg���6`�Q����^F�\L=k(���a����l��j-�mA�:���׷cI��U̟3��^[��J����U��������WK!Ӽ��A<zۍy�^5�N���Q�Y� �E��4�C۾nM��_������t,�Z����z21"a-M@%�7c���u���nyKYr[!�e�&�@�^������}}���6iX%V䗞ta��; �^�{��7��+���?g9��BI� ��g2��W�jtM^h���w���"����^F�޺�jgo�z4駉'�u�b���\�ڔ�i�Vd�T�9'i�j�0�(�� ��다���U�dd�y���,�|�S	��q)��o%�x?�K��,�Lۇ>�7:�j�< X����ALؼ�5�.6����e{�k�M=3ٗ1󭻃=�]+��=Wz�\��C�1�crS������U�P��v!N�3�
+a��?MT6�W����X}����~�R����6��-��`�4#η藿�Q�uZ�[�ӡA�
�x�ۜ�� �F��3����h��Dd1�^��E��W\9����oR�vf�(��`�8��EK���-�����B�s���L�d���R�cr�CMbe�f�ΐ)L���	��xr��{Z��lٛ������5?p�$�1!�2su�gwI^�RS((�P�v]�Od����v��\BS�;s��1��麚��u���[b��\���$�]`I�n�����薑�[�<�=������hFWS"�"��:��kxwov�m�N����}��.���k�[{���*����&*��fJ�'�6o)�1������z6��*7���RK���,�򔙽�u|� ���u,���"��\o2rw�>�o�ֽ����mT;B��cw�t�ūJ!�pZ�r�p|�����-����z��t@�.���w�t]�_��A������{�}V�qg-�[�M�ro ���{�Hl���ρc��vm�^G�U�Bl� vE�Иe��2(y�2�м:X]{�*�n%jXt�p�=��V�C��$b�<�pk��d�b��J
���&����p}���=�*�z�!X�����3u~ѯ=��c�U�LV��]
�*s0����e$�I�fj��n2#�d�"i�=��;ƚ�7�N�|�#������S�b�}��{�6�F�a��$���7�0��(Ⱥ�C52��6�T�}	Ǐ��9�'���y��C�W�p��Nߗ����9�sFL�|��	*�Ѷ���t����:��Avj�I3*�cg�ti0=�5�\e�f��r&76%[pe�Xe-�vY,����X��KL��L�LlYHqxwgf8��s�D�]@tj�͍���!lPa�S0�8�I���8�tm�KYf �ō&�b��#,�����ε9���y��Z�N�4��k�=��v܇�^�V٬��4!5i�r�؈;�-��q�n��J ka��zr��"|�V��!a�v��Zm	vu�9����>-���]�p��c�J�EsX���,���Rn�{1�����ۧXz�f���p��[zJ|]��m�rq<� pxwnt�k��;	���$�+��bР�r��9�.:�nL�p]�[�\f�{a�$fm���"93�֙l�8	��d��F�bm.��`��GLE����=��`�]��ZF`K]*��nA׬i��;%�7%4եz�y�sګc�G�/m&�lh�'t�|2�sVV%d4q,�cI��oN8)����ƌ���y\B�59��X͛��5.����4�j���m��,���0@���.F5l:�^[�k;M� ݋2�a�\k���Y�LiaW��m���cb)���2�ˋ��N��M��{���=��
��;����R�2H[N#�m�hK�E���#ԝ����M�6^B�s�����v�`����\�fe�Rܬ�V]���-�.�X̌� ���Zq[+cv���ڪ.=(�$������� ����csm=Ɇ�$���ɶ��x��q��YI�g]�ݭ�ra-E��ް
T+��x��u��^�0;� ���3�ۄ9�&3�Uݨ��wlRkt�u��큷��;�nKv��7
�(n��͐��Z��'=!Ƚ nEܼ�Xd��\����E�%�`4�:��MK��QF=�P�$��BlL[
:�0�͒3��v�YtmR:���#) xW�co W6�\�����ꭺ`@�;��Ѐ��	V�k��؀�S�G�� ���j=��]��Z��x�ne@��t-iBl$ū�ܨ �^a��^g���c��7'�X�A��!��o6��;[�aZ�v� H�u-BTWK&�*��B��#��d�yX�E��a,�1;�]N7�LT�������}��6�?
>��) ���t*,焹��6��l �˿F�y��A��%і3g�{x
�/	��M�M�h	��3x�޾��0�bϻ��K,Z�Ne�Yq���=A��Fd�S�B��{�	���^�#Vݐ탦�Sy>3�׋^�Y��.ߒV���K�@�u���M@ ��Wh���͙�8��=�T�z"��p���{��뗌淣�=�st�{9+��?�OSeC�{�f_�����ŗG�qY�e) K�Cp�\��U86Q�^�W9W��;?x�0��L��u B��sp
����E�2<gd��������S�i(�}�n�$f@�����IIqW:{�g��2i9N��<_�]�\������;�3�U�/,�������#��k���M�P��������U�/�۽��������ۭ���F�W�䢈^K'uW���ɻFa����}��麀^��b���u�+N\9(*�#'z��u�307��b ���N�)�����Y&Fd=?O��ID�(pU��z6��M��#��7G�c&\�P��P�]C4zae�z��^�u ���@rX���\7�`�n�40���TǷ>��|�TB
o���t���7������,ߒ�o�i����f�ʘ�
d���:��sn�nv�i�p��܍y�{sc�a��cA���]7����oK�c\�b����/�e�^������'�y\��d�`��41��o�H3K�k��uS����N_dhzGz��01t�<���nyձ�T����V��/,ao2�`x@B�>
��a߆��"����X����_�³�pz����AF��3�GmM*bf;cY�F/o=���bk�K���������,��w���L���͹��(*)\�7�+x���<���T�egm"V��v�K�8i�,"Jl6��a�ǌ7�2���Nog�#��V+)��j���Ϊɲ��h�	�=���6�O�?Y��\��,��I��a�Ӟ|��	G�-���u&�7y6YP�I��Eb�C�N�x�{��sVv8�ʳ�t(���F2^������W^�}��fl�݌R�5�i<�q(�3^p}���]N#�̩�����՝�s�id�����;cVἙPiˮ�2��!u����zz'��"��[�5�w�S��d��:C��u�V��i4!��j	� Ͼ�ڊ�͝��L��}�����$C�~+����֕ںc~����%���b���s�V�����
yJ3S
�e#��n��G��B��h ��_Yf�׸HZ Ufh(���1���~UE�W7�Ҋ��6
[
+͹�O�������ﲧ�3�����X�����QbY����e�W��O8mQ0�]J9����K���� �x��&Z����"u����%�筗pIsƯ��J�b�S�x��5��� !�C��*p�֕�3{ۖ�㛊�]��fjoE���!u5SZi�W˯&h,O�CX�%�{[*�f�M{*Xwy�t4%À�=�Y�\�V�\���J<;,�ZNO�j��/���q�(�_���~�����ԥO5d�&i���$3��$!�7:�-]w�7�8�xB��m���'�.��y7�/juT�\��q;~����W�Qq�3	��4i�ޚ�w��Re{�Ɂү-3�q]SҨ����XtN�T��)V���w|���!�+��T�����@�n�P]�ɳ��&ǣ~��eiѩ��W��p�K��}�-��c]��6VLVZ�*\w%���b���@OC[F�ev݇���Y��pN��D�ĤRc��e<�ҭ۰�V�n�L�!��JHj��Ya��]F&ں��ΰ J�FRd&@�g�N�z�{{\-B��o	�"lr�˂�.�ۇKn�
B��_��o�F�Ł�N�u�'r��+Չ��1ɛ�ls����9�5��;*�ۆgEǐə�z�0�"a�6���v-�%l����31��I�U�ηJNGrq9������`_���?��68��(H�++�
�]�p��������K�����>\`2�"ۆ�&g�Nv������.�]I/5 ��ЎBk��V'�;"�t^TT���̛�k	j6�������l�S6�.]>:O�6(�]T�,܎��Y���8l����{��5#Nk��^��{B�d�q��;�3q����=����lq1<�� ��D[9֞(�m�&�$���F�=��j��e�/�x��
�l�� A�|��{��mϪ�Re�u<�7C��S�e������K��i8';-_Ϳ3��/����P�۫nR�}�@ӿ櫯�Xah�^Z��<B���i{X����:��(��	te�'پ���L���e����;G2��
��*(��U���y�D��trc,X�Q�ё@���I���:N�cE�4��^�Hd>c��2�?{�99��>�K��6�*�R������Cl�?_%��L�A>��br6�E�Gf�J�5=s>�a�ܙ����P񌫻�$�����&�r�x|deI����#�p���u�sN؍̔78���ft"��_�3/3}S��C�ōUtL�3�7��f���ư{%?YX�3�^�ӿ�u�7,���r�xs@�J�Ӛc"������\j��}������sٝ����#�]��� ���hd�Z/z���o���~	vxC�}�S0k���!�aoWQ���ܣ��G6�i�$
�ȹj{ͷ�95Y��]
yo��{_	�#/�׷���j]5�"�bX��(�ŠiX�T�L2a8mBPP 4L�y�!S��@����dBx�S���s!�Me�f ��5�q.C+3�w�ú7�΂K$4!���ԑ�|�oo��:/��܍�={Q��j�2�^ϕt����'e�s�N���&0MA���%�qS���I�u��k�P,ƴn#�@��V8��T������N��n?W�B�AW=t���~���{�v�V��-��OJ�+��_Z�r�v�t]�&��@�p�kb�a��8x�/'��BL��P�Ò< m6R��!N4�iN�.��v"��&�����<�e��K��E��4�`�mv��Y&gӳ^]g��t	��ō[Y�B�a_q�qI�e�P�Z��;6*�	J�F�Y�W�����y�#K����6��o􄫭����#0rj� ���"71�յ��)�q��\�N �kz�E^w̘jI�L�I�4���O/k��q��-K��Z������,h�h��VS��-��P]�v١�]�oa�����S�aA�;=���i�7�:g\��RK�du�Q��e�A���w�*�g�P��YW8G#C��"fY�5�æ����~�Ov��s�/�����.�\ޫu��NQ�?��]��?t��/%�XwF�����ҭ�sSm�F&��EǏRL��Q�w��=ļ�d��8t��uׄ���:�.�6�M�T�S�Z�ٺ^��'4����o����js�	�T��K��ɗ�:8����Hf�o-�;�*�ޛ~�i�������+�Z�]��d��"Vb��{a+�i�7jk3�^��7��چ��;��{�5֏a���1�x�STJ$��~��;F|W��a���L��
���>�����3��5�����W}���O�]�9?0�α��\{�a�2�&�E��7\տs�eb��>�g��*}�n���=��P�p�*l�OE�R:�Va���e�����/��1n�<�������)�p�W]�K��~VKtb�Ɏ/ �.���Og	�=��h$Ä�#QD��h5X�e东o��jt�`�m,S�����DJP�E0��i��P1�qb�E������$9���E4�m�aT�������k�T�:=g=;�r�Z!H3�����.�>U�=&��x��e�z����wo��f	p*���)A�4�t�vXw&�}�9]M�F�[��ד�-U���U�ߎg4���i1�N�T|�}�L0��n�g���1O޻��R�W{]�Fl�|K�� ����e�&����x�+�c��dm`��)5; f��:����)ܭ �Z%Fr��M�ŴU8��]�������q��.��ʝ%3��+�ڋ��C��\S����i�]!ۜ풴Nk�j�Phٽ��Q/�޾D�Fn�����%#KY�A�s,�y��$�4�*j<s�������X[��	gm)]�~���$����{w������1��ॳ�	��[D)m�O����;\�\[�O�J�����L�T%��+#��yg�)YևF��Z��i�	y������o�>�染伌� �17�8:�f`rB��aN��᭾��9c�n��գkg��5��҄y2I�(�=�Ir�;�,d���_=��i��A�M��� �|Fa)La� %
i���kr��s۞.��ic	��b����޹/�}�X�	|���	N�a���!�,F�"��t~/����g:H���m�e�K���N��i����h�'��nM.�7�Wb	<Qg0w��oǚ�W�Ѿ�|d�-�$Z~ڿ�U���^㼺j���)N��{/#����eo�a[L�CA��3���t��کuY1�=����֧�Cq,]��̙;�a}aC�]5�L�Ws�c��x���1�ef��z�G�_��Yy}�g>zRPD4b_b�3�@��Y~�t�-mi�Z������x�Iw=�O񟈹��5� P���V���L�w�W��_MP�O�l��Cn9W��\� �ƪ|�~sf7@�Ҧ]M��,�H�=��fM� !�a����6�i4�%l�״$�:Y-�f�aAb��7��GC��J4��H،mIG]����Meқ��Ia���v��3�S>��ef��^ڲ��#�;=�ۛ6;v�,h�V�h�"5���z6��o{1��L���D�K���F4�`ދ��1�Q���s®�1뇤��m�r]̢�����Є
!��4aA��?����\ښ�~3��Ea�/s�5վ��<�LP�Ѵu�{2֬�A<�iBLMr%�����C�~��Ge�{S��'�'���t$�!/�=^Uz�wGR�$֯l���аF�GӻQ�`m襎�}�sM*q��Ƀ g����.(T�B\�HCa��O��緖b[ԥ��#yӊ�k�����U������B�@�࢓PDbP�g�O$���n�<ޒ;c� p pI�	��L�v��k"�.�d�q^�J�x�g��4'�`ʝ���p�M)g��UG��[�Ԯը��6��	���f�<���ս��{8�|A�!V���z{oه�-�2��L�{�q�g��tԜ����bB�r��J�D�e��n1T����Ϧ7�@0�'��r�ȿOSt��9���=�Qq��ݞ���_i��cKe�ú=�hڟ:�o�s�sL��(V����
��3{�uu�F�� �O�V�^T�G��h�p�l�#%���*n�G��B�b�[�������qU�}x�c\�HS��je��Nl��D���hf�^�td��Q��i�k�i_���F�K��l��J�o������=�*:6:
��Y���'�:;�u��v�1���XH̲���gE>;Ư�������^HM��������yuo"z��۝�+��$#u{,�M^��&��6Uٍ�����>���'
x^e�Ү�>�㵛�9�]V�F�Օ}}�\n��R���XM�Ր��绐̣�r�/gB�ƻo��$�%���␂�� ��c��ؚ$�խ��z.�i^l���l�F�r'�qIq�X;u�S��;�㊬Zs���s;�6s�*N(2��?'*��M��U{ۧ$R͊�9}�v��^pNM�Zm�$�5�o8�on5%�rq��מ�YЮ�����?/\�ݼ-�=���}\�Cr��'�np�-jxf0Z�u�B4��x��H�*qSNz�e�T��ã����^Y&���c�������/�弻h�;Ɂ�����C�wcy�l�%]���3��Ƶ��g_��L���)>�k�s�a��s��wEe��� ��`0\�u��||����]OF^�e����nì��@ھ�O]��~_t,��/�f��y��^w8�ؿ8K3IG��,����	Ό���$���Q��{Q�Ehٮ�fg{�.��E������cy1�Ǘ��D�KO[�=؋݈�߇��&Xo��9��.�ʜ����k�Oq��>�8R���9�k�^�xe-�i�(H[���x<��ۺ�2m�#��*x>�:�$ �>��܇<�ݹO�a-��[4�6]4E!6{�z��-�ի7���GT��HO�o�ج����b���ެ�״��nX�r!g{nz�ı	əd#ԕ�Ũ�ͷP�����<!�0��ޞl�).�ү���.�/��7mOwFu�S��XFwm��<���ô�S7	mD|^��Y��W=쁣_���$(�<q0�Ir�ͷ�L�`t%��h����}�}lR�e A'��b�Nܞ5M��sy�yg��Dҩ��n���D��K'��#�z�m�a�B�hكVH��;��`���z2�KQ3w�ߍ)�;�o�>3��Y]�1���F���u��mod՝~��w��[3�֘��8E�9�{�f�Rw6���2�e"�,���/ҥ٣��%#h�L0���T��}��H'�T���-�����z��v���xN��vh��ȓ�#�#��-��fU<բv����c�2Ȇ"��to�V�g���Fr���U�s� ��ެf~W.|�\�^)�dԀHm�#d3*��:G��(γ�G}φ+�K�vmgb��^	Y��%$�먹���90`��p�= ���b���w�w�=<��������zb��,瀰�X�83������.ù����N�}��g����Uv:s(�q������Qk�,���}<y��)nd7F��ܥ/���q���~Q ����|����1�U��9�����q-�M�\$���$ٔ���:�o�i�9��7~��7�A��D���݁6����2�w�1�j}�>���r��~�5���@�!|S�y�o,����Ղ�{�U���lY,�*�݁��妞̉W��elL�0�n!��3<أ����r
y{��<+f՚� �����Q'���߮�xR��Z)�
�wq�XW�$,ّ\qjo�i��փ8`�qpݖ:X��Hy�.����b�=�C̀�pù7E+���G���v��Z��#(�ܡ�1��ض�sڥK5�����E���v��vv���nK��<j�㳆�D!i�+a5�3�uv~�E;NЭ� _��9�kq��i־��Ǝ�����Q(;N���Y�
/��6N-^��y /ɐ�ʻ�����t1m��h&+ʱ�B�5���;cej���[V��"�u�Uu ú��+ �m'�˯�v��C{^%��˽�������{@#��n�l�"��$�8k��t�變�h�'n�r����SvgtS�N �l���X@0�)+<�]<��W7pc���,��&��Ӕ��;f��w}li���\fY'8`要؜YX�a9�Axή[C\��9pgk�D�TR�jj��Ξ�7��8ﯰ��y'S�æqo��M�����U��<X�p�P��yz���Z���E�OlT:�p��mln�ٺ�� ���}�-މ����% ���c]pcYg)'3C��S	�]̹�/��hᴞ�õ(�j����:�:W�H]p���ǑS��S�|���хU�C���
�^�#X�����K�C�S�ݡ�-��]���n��!��_�������E�+7��l��p�?s�3x2iw��SĦ��U#s�4Y��.ީȻ#ӟAة��Oל�+�=.����\���,��0��皽?/J����*//�1Icc�v5<�RQ���W����`5iN[q�z�q��d<�!E�ɚ�ء;g������ǹ��R���1��2�훚$Ü��əڜ[�(Q�(-C�C��js����X�^؏X[\�B�K�fgm*�n�.�Dj)�\�m��ZQ��e�RB��~.�C���DS#������>6����	�pK�Zݤ��Y5c���"��lpI4m�k�A�T"J�H吊�˥���HzTK��`^g ��|%�;���t���Y�Վ{�gع�W��NN�1ٹ.�۟�}��P�нݐb��e� x��r���w:�S��௫=� �&}Y7!��M��F�B���Ȋ���K�L��L�ˇf-�	�&��wy�����'�>�6��]�\�qww�hU���I�)�uҠ�ʖ���#���u�e�{2*�
u���1ů�NS��"����
53����|�-�����G�{]�<��V�ÍZ�S�%�����_{�K�� ������h�&o?��W ?G��7.{��]���J�~�(��y���|��Hg�ۼ���@�����H�� ������.��k�B3����33�g��Ndd�ޕ�u�鹻��b��<e���Iv*w	n՗��_�p��m�X�Yf�Ͳ,�ɫ��'�����ƹJ�����?ͥ�����9���L]�l]�pL��Gb�u-��������isB<������5�����#�;Mː��]�F9Ls5��Ny(�qs��]8L��غ��B����`����U�c�m�]��'�<�ecYl���J��[�;րt����=����0V�����69�B��g���昤6�ˆ[y�{S����ʪx�e8�b����qف����Y}�����ay����Skڡ3U�?/%]�ͫ�f{&{.��
D�%=ηK���̒ ��D2y�h�;T����y�n�:|��VpW�J(I<C��ie���8�I`�^ފUZ�_z���r�N�B��P\�S����C��=�As���t�����E٣��ω[m8
e�ߜk���0�y'5��/t�-8kP�X��k�F߿��z�9�ح��X���x5v2�v�E����l���$�=�gv���g.O�G�u��ꋾ߸L"��r��ޘ�p0���@z��~�OX��2q�1Z2c_got/W{c �y�H�up	������c �59M\r]�����36}�$��7,vȫ���^f>�*���>�7DR��t2u������V��3�ȏL쨬��#=#�\ -�H,w�H�����%��Q�پ����.��@�qY`L�몙h5=ؕU��kr_��3C�ݢ:��~!i�t�_��{��jgn�`fJ������̷���j�M(D(�1	�f����E(#Rkd`����x:��)C�3���n�x���{w�v��yWi�5�<�%���ܫu�6����|tR�ev���Z���;2��A&�0���F/���]��#����)e#����9tBC�I}�s�Wh��4��d%����_?k޾˙V�$gz>��6R�լ�K+�&��Rs��s�9��j�^<��M�/coޞ>�^�ݻ���P��°��{ܭc׽��<+�(}^�<�k��t������_��B���\ɐ�h,�V��,����UL��0p�#L�{������@�à��d��1�-�8��ۮ����Ivd�dyNЙڮ톷\;���>�ﻯ�����������'u݆�o�0�J׃�oF���̜��:��0�[�� lf�M�&��r}��u�H��LXf�3R�������+[�H�cJ�+��ki�NF��S�H�P#i�[��VJ�38=���y+�VC�ݴ>�sϞh�V�c��m��;�whg��ފl�'��A��[V�T�/'c�����s�&���1�T�8�d�~0w'=�VD:>�k�'�}�g��3�޹���[-�<痳3�7����oDI�ɸ��K�w0��a|ӂ�
�{]��I�\�}��1x�#I�Ι%���2�8a[�t:�]O'+xB&���GFh���f�N�ӄ�FeAs��ʇ�Q�vH�De�L͛��n����f
 �(w2yD�p�p}=G��Y��gz]Q�]� ���kԾ��j��]�8y�(�p)ؼr���r�W�Th���Η�oz�����~�,��qXw�w�{g��Sγ��`F)8A��'��j�L�vMZ��ܜ�Ic�E�386�}kh������S;V�p�X]l�됍	�gqGe�3���[hi��zw�7g���qS���'�L�6n�|�>��?)��Z��[��5"����a�L�(R��R�<U���N�J����>�@E[+7r��8-�c��}},lͫ��q�}���7J�"��zky��ݾ����(�؄6���s�ũN`]Kb�b9w8v�&���a�y3���޽��u՛�y���+2�ʶsV�U�:�j����g�	�*�N�ǜf�JV�{����8�O3�u騺����%Р�@_+U4@��Rdb��2�M{ˢ:��y!�t�n���i-�N�Y��f��ݻ�:&�w ���4md���˅O�X��\�f��0�eWn	��8����"�.�C��ou{�xg>��H|V��~R�	���+�`��a��=���o~7���Zs��n��g����'͡d�dt&-��ZD�5�+�
����=7�+�	l@h�a���ź�fׅ]́�{��=���7�e�+^G<���Q�
}�$P���|�|pw��p�@��{ӨRz�h�#�����mR���˪M�1�ЌI�s�Q��pEk0�L��q\���ު�2��p5���>���R�[����j4����&]`M	��If������1V�rs��DճY�1	�7n����{�OR�-(���䡟LM��<96Mg�q���>�w�����j��q�O�_	����[-�6�_\��,B��C�'�v&�7ٛ>�1��'1i#W���27�`��=CԶs�P���݊����"!U,2��	�.W,F�Hb;�{s^�U#Џ�L�e��g�+1�S��0:N�Bm��ٍ	u*�W��j��/��`�1���`K{�RS4b��BF�k?����8�R���8�,�sV���F�N�"�!X&oj��.�=y���,�a����&p���ͳ篃���0(Y�����ｫ�|�'1��1g�W���nO?�4��]B�v��Y���|�k�}��"�l7�/.$�kɈ�cy��{��P�+�yy�f����o��⛎���Mx��Ǝ=S�]�s�k�<�F���R�P�r��it*��c<���L����3��t?�B.��
������[y�#�h�
�`���H�#�L�����J��sYz=W��]B�o{�n^P ��q!�M��m�9���M�ye�㤲�>���k��r�������Ml��nm0 \��r�ƈ����)��}'I���'|��'��5��ct�H�MH�8��G1Zg&����f�+[��Yh4؂�?L�������b��g;�_������M���"�-�	�	�47ݞ�"(g��.=�	3�7�9�K�w�?c�TwF�i0�J���7�!����K���U=��Cr�ɛ[�8�9�ySl0dݴ�f�&׀��nO{>��,�j�\k<�s��՟M��xɴq��N]�MB'���$KB	�TZQ��r�^%�K��vpg#\�{	.�Q2e��~x��=^���O�
���'��8@�~V� )���I���ٺքM�g�`/;U��7Ĭ=F���q0�Rl8j+������ݙ�9g=�M�PH�F�z��2y�b��W6u�@���[�����ْ�E7=Csv���k�dѳ��a��ɿ���3��hDv�����XW��"�cY� Ђ�A4ɂ`�Ym�#��=7�~j����8
��ΧW��v���+��]hM���A�=�q#�w2�9�s���ʛ�j�i-!����p��sU��1N��rώup1�NzQ��=�Ta|e��	T*	v�F=��=q@uicf�f���d#U�۪�v;A���X� ۈ�*��!Ǆu�s� v�� �vP�O�U6��'�����n�%J��߽�q� 6H���TF`����H7�&�٨��]W���Q�3c�n	A�
6ը'���c���a����{��Y&�Xmg��,��鹩Q����|!:œJH�	�!l�={�n	��T�v��ӱ��W�I�$t򶒪�_0&���`�{�bs�FpQ�(m	�LvZT!��Q7C�?,��7�dik\�|�������q@a��3��$�B,e��Ů�+�$4r����U�_[*\ =;*;�{��2a`1t]J�5�EY>�=��h�F�61/�<�M}�z%��8B�34v̑�P��r*�pv��{:���W��.H�T�%O�*mĎ�^��ZP�M$9!��93㜷 )�s?���p�&�ozKB�_��Z)�(�x/n��U��=�yr��juw�S�wٙq^t��d�	�UcRJ5/��ܙ��.sܽ\Z����+}�U�ݦ<r�c���^4
��Ka8G<������D��L�w̠*D�̴��b��3NlM>�12����ǹ��pRi6�^���������{'>SLwC�s!Y�/OҋU�4�>��t_eߪ����ů_�Ubhl��S��ͫ��>�~�r��Q�J{L��'L.����p�7j�CK$5��A]/h��w��.�g���wF<�n{3��ҋ*�U�]5�p�B�F8A�Y�f2�6�T��!�?*���
�w6^�M$�h������Ԣ��| �/�w�o'�x�x��y2��E,��QTz���P~?�*����v�꧹(�~�Y��G�2귻� �4��C�����7'�^��򮪭k;�[*�w;��P%9�͉�ҍ��� ���)u�9�n����e4G[�;j�-Ŭ�ͷ�ClF��>��Lf�a1��.�)&{�v/a�Dz��%�vs�:� ��|.9����vg�r�V����1��@��O̒�!�6l����_��X����(y�D�d�gS��4�B+��F�����,.��Y��ڴ�N���������!+54&J]K�lfwD�������I�+�*^mɮ��2ogǟ}�1&�C�]��5?O��_2�1[�UȺ.���:�|�^�UUF�����_��ɪ� �b�'�f��G�-�F��U>�GF�6Rd �eCS�=�04w��,��#��'v߰����7}�w	�N��D&h�vk�5��Od��sּq0����[;`K�}�U"` �CoI]]3�]�V���c�&B-|#�qy\��ds�����pd䔓�ݻ|�؆F=+��*{o��;��[Q�h��qX���:�t9t�9��J���h�����,�����uĮ�U���͟��Ȑ�M�ɲ�X���3>���x���IoN��pBT/LWs�=C�m\;���4uR�^�e�m�kr�l�?Q 0B�� Ϸ;���S�I���W��ɩ�6�gjB��I��>�ٓ~�c�թ�/l�^!��H<Fjר���_�^���S���l�687��l�{���Kq>�pfF��e�w e�sy^-��cne��o3K�A����C��yC&
b��l�Ʉ�3���1j:�m��Ĩ�K����geK0�.:�k��l�@u�8�{0鮆KxŤ.V�t�Ph��*����k_wn<�G>�=�L�%�ֵ�=�����]�3B�}n(ீ���^�V�>��lV�N��_�~z�K�� �nn|4�ǡ�pT���|�*;1��<SU�4�$[��.���� &�0b�=��9�f���tN�*3���a�*R.�s�U��Ӑy�mw�?^ٟ��xxAHE>*�C[����=�{孡��.�&�����Ћ��U5���QŶa6��T���s�سf�հF���������ZJ�{9H�&+�U�5a�n(uqk6��cZ��d��]}2��m�� �ٛ߀��QK�\����4���V�q�R�vxE/F���ȷG���:y��
r�vo�A��4F�$!_ԣ��!�n�uy{�k�ئ��m�81�nF3� �A/kiM�w+{�M�H���4zk��P�'�R�E2��ey���(V��a3�<5B����u����k���L��m��$��~�Gr95膽3`�
���\�$���>�B��<qn�l�Ne����Sr����q�0r<L��r�˼Ș34`��)c%��2�6�Aw����Fh�M�	M��!�l�Cם���۔��K��p�뿹�U����(G��fLt>@���ݳ1��aO%���{'6�[�)⭅6��M�m)��i6��w�X��'6&wi	����戍D��飔�%/���ge��ĝ�������z��!eu�rDu�|����<�����y�� ��X�����|Ѯ��B���_a._Mݼ���&��7�_GS�ľ�����^��z,r�a���>����~��Τ2��Օ�Qgի���ʴ{Y�n���fՓ{3�@%eC����m|}�`v��ɞ(�f^�o�����m�s�XN�7N���ZU�C����lؼ�}�#~\��^�>��Kn���`�(yT�w�~�@s���r�^�Q��ב{�؈|�e��6�躹C�H�kc�N�w\�����6p��]�8m�q=O>� ��ೳ';��c���)�4x-ٸ�Y����'|�l��@��Y��~�i_�n�p�=r��.f�g�x���dP'l���ֺ��;��Mi��Y���q��b��D�U^t�O����p6��3�^V�s�Y֨��8�tq}av�Mٞ��	�=�ƽ��L� 𝆖i�^(���+NFV�=�/Z��ݗyJ��>B��s��ܛ��3���y�Q�8i�Uun=����wdǽ�g��"���M�9��e�#j�b�f^
Wl�/��E���d�HB&9��G��]�7	eX�Kx�����SW,t�^���棄ӽ���h�l������b���foa���<>��y��L|�{�\��w/�K�;�|����9�F��NxzV^W�/x����O8����Lm�Z>׷�g^	�
���t��Yf}t������4�榺�y�&�$�x2rGuѹc����YCs�n�f��6����:��nk�g�6�Ƹsժ0���<6��|t��33s�ɛ������-��9F[�H�����Fk.Y��M��fw8�ۖ��{q���#��ŔkI�b��^C�e!�ܹ�l��]s��:�n��G�P!Ҏv�B��+)���;a��n�� �'�����M^dbY�?/ߧ�����;ʊS� 
�o��E\���6�:�3u�� �`2�e�h�U>��;/���Hyen
|�7PS2~�Cғ���^<�'�]ݜ������y:w��j�쌚�/r*�9R�'���A�me��;��^G�۳V���������x2�i6�E�n,A��O�M6��^e�;NN�u&2ca}os\s�Z�p��g��9�m\Ec]u)9v�D/s�����ģ�-�M�Y�X��Ox�M��6YE�������]�l�a���TUL��f瓊H�[��yy�0L��2��}7uq%(pl$��;G��<5�f�ym��>Ws���׷h�B0��m��w>3څ��������2е�@�C�����
D�;���z��>��8I��C!a����BU93�;�a\�h���&&=�2�f�ܖrs��<�*J���ڔj�D���G4�p:�"��ق^��� �)�.�n�\ �x�$_z�+�u���Rm�Z)�H#��3G:ӫ;���C���)��0<:罓�� �u��C�2#��1��= �d����uf4�
 �������𝪷L)�0B���55�R�Y4���I�ۂ]���/�4J��S<:��Ň�*�.wO�˵�{u��R`Q�]c�O|��m�w7
�z�0|H9Ж����#�{�|�׏)D�	����Ё��m�έ�O��
�|�ؼZ܍������k����+��`��4�Y�;j�~��/"]EV���z�gx�y�#u"��;��J������ߔ<:�'��Z��7�x)!{yW�o���?O)u�g{�s3�L�v�o���cV#�R/��ώ{/���{���u�5J9,&��cR���`�>����ܗ]�w�Ǖl����^<�]H���5d|Vs�>�|���; 9�V�lvZw
��3i3-T�8�Z����w��7u:)S��ulno�o�P=
��Oc���v���O������I/4|"o��4Fb��������a9yɼ��Oc=ՒS;�V06��.U롼�=F�E/���!\�㭿
�k���T����]�0��a�b��M�`��g=e`�p`���5Pe&�@S��lJ�̱��Kx��{1��y*34�S��^�
����*�@��g��.�Y����E`��?`���7��|�K�3$m��3��p�,�]gXSE�ck&���*]����s{�u�;��]�Wn%��1s���-;t�譼��N��;��3����{M�Z���{xm�goj	�x
�b�y��i�x����]:w��>�RH������=������BDi�}AԮ��-型nw>�6�����h��ۂڏk�vz�˓���'kb�J۸G=� Q �$���n���p�m�)Uvh+�BS�W�jb�h�0:7��<n�lvΦ�Dr�@���v�n\�]"���]]�L3��i9�r�{.��=<]��1�d�-����h6<l�+u��WXtO�qM�`��)�vO������:�]Ƃn�K�l�]k���[�|t� C�N���^��nݛ���va��4���b,�ZR�
�G���u5��X(z�۹w.=>�E �x����v��Ms�rA�0ڂP���5`D�\P�N��\n˸:�F���n��k�95�51�D��՘Mafݬv��+�$C:�b1Pvf�v�1z�kW,�zm�ewd#.��D)y�"�ٰ�2S�&PFp��H��U�.�7��b�$c[�c�����R��!"0H���C/R�6l�!]���x���{n�/e꣪݌�x����s�l&qr�|�[o=:wo3�#�3�C�9�z]����J{v��i�^Վ�8]�L�]�]XF�g�`��l���3��
<n:�^-�s᭠��	�u�݋���v��)�N7n�/;��d]��C����q���q駝/wa;lkÎvs��]BNn���k��LDj���6oB�+gy�1۸0v�����Q�f�>�p�����l��s����h˻D�i.����EuV���.�K��QmhfV�ݭY`���Ц���]CM���SC�nQ2;�].����;�؝��	�{%��l��wZ=�<�l���TH��v.�X�1\���8f��F0�G^8�:�)r�����gv6x��x��i1�(P���W%zˠ�B2��eЁ�A1٪瞵l�;�`nK��z��3T�\��;,��0�4�c�m�a�WB��
1�{�;6δ���î(ir�y��:y�e���=��S(nu{]����b��ԛ���z�WBvǷ;���z6v���I9#5�l�g�cx�(�m#���� q�Vŕ� Q1�5
st�0 �  a3&��ݎ��]NA��t�{&j�;9��;؟^v��32�a�����>���Nsx�s��jP$<�=�kU�ӿ�Xf YF[�C � b���.T8���"qà[�;srDI�[>����#��#��*�"u�wZ�'ЂխeJ2Tg\>�n��Sd������ Wn�Eu�}�7�%�����?Ђ./�'��T��fnS
:H�配P�\uv�~w�*v��F�<�jY:2}зǳfn2*q��D{�*BQ�^�#�2��ى%�fP��HLql-��j�;�:C�P(��'�;���h��:C�W���u|e1"%��%������[oT�74S��r�[Ҿ��(
�l[���Q*l�i�S�q�pׇd�
$�r��f:��sc�R�,��I(=����1���e�����7ǃ;m���������FL�=3qZg�Yu^��}�7_1�׈<G���V�yL�&v�P�o�����qP�Æ����$����;�	>�L���cq�J����μ�KQ��dƨ���T5IIVW�9視�Nfv�n�x{�|fp��IU~��~톀zj��G[%>�9W�"�٣�qpW̸iZ��b�3eM.�1�OKD��M��.^���b�t�*v0�a O��lT��� I��KH�ъܙ�̯lJ�s�~I̚��}�h�p{ �~Z_�|�rm�9��z��8F/*fE�5F#�ȱ�b����Ϻ�e�� F��{w���^w��Ϭ�s�^=�.(�����.�?�N;&r��i}�=S�pxo-�ك%�BTR��r���v������І�a�X ��Gq�f\�/��9X�q�ԯ^�8Բ	��cA�}��l\㞜}{f�!�(5�-��r�Lon⡳��ȷ���Q��ݷU��)�Gr'�(�)4�\P�ἃ�dE��Yq����\d�)ra��	k�G-c�z�Tζ笌�j��
��F>[��*ɼh'�T�i��/{7A�m�F+�≆T��g��� r@��HZD��`�ɘcB������A%�y1�GG{xM�O�am@�bbu�7����QY�w$�Mv#_T�+�^'���'�/ʌ�k��)����,�ƈ�s�tj����i���yMn�S�O�r�cQ��}}�"os:�
)}l��s.Q�T,����R]ܫg&�����B*�F��F�{B1����W��:�ANs\��s R6��ab�˫�W��#K0�"`�8g�Ճ�8k�W�sB�)1��F�ad�lʤˎ���i�$i�F�fĺ[z��T�$�%����sX��B����~���������6��3�GD#��E�J�%m��9���˯�����os�[Ig�t�̖8d�;Ƭ��At ��(M�^�5����]AG餢Ou,�����r�ǄX��.��i!d>�4'������|n���i+�|{5'�e����t�<���o��7;wj�3J�����E8u͔+Rfr��(z��>;T��G�¡��J�1�[j�s�(��헢�������ƹ�j�@�i��J��5������3��3����'��� �s;��={7"��<*jԢ�ۓ�M�C����x��	�u�eUg��V���g,j0��>s�S~�޹��wۼ#)�P[	(XM[�r9�١������"i�(�n���,Ҟys��w�oڎm[��2����Nu�#�C^
�l���<��a�ǝq7�_��W�U��͠�Sc�s-�Y�?5qBD���E�z#Br������2�.CD��r=�9�^��/؋+����0%۱+)���U��O��r�.�%g�G$�ϳ��#"���+��B+a����d�Q+���N%�D��y�>�p���/fɆ�D��z[�w`�2.6w�v4%�����oOM;����|��w*�lX����qn5���W���~�߇�"�Jt=���,���,f1��^1�>��Ts�9#}�?_,�/0�7�/�wxFg]�C��K��XY+
`������:~�5z��86F�����{�W�V��oV���h�d�5�Ϯo���D»[;,
�є@�����>�ac�qX_�(�l�-�/E���@ށ0�b
pIw.�1���b���@�����@p�ŋ4��;�X��>5��]d��g�_CE�A��p��j:hE��P�X��/7��SG�q@�Y��[324A�+'m�Ndv�L��)��eX���Ѓ��&M{k��wtQ-fk����CD�_�T0Q�+��iϏ>IM���X4Nм �N]l!�Ԇ��{Z�^�<��9S#�K;vJF��1��6��xU�?vs�y]:x����R[ł.�b4B�Sמ�9�}������:��'*���Cc���է���0�3j�C�$�����T�t1�_�����`��^�m^�#�m�2�\�6BS%�"��2�y����nT���,a���(޻�:S۪°:�"暗ZM-�9�6���d���A>��U�9k���ob�`^N�����*Fhr�(����ߟ��$o��	 ��t}F͈��z'ֺ����V���y�'���S����1�����3@��!6�A�����k}�'��sPر���s�=j�֋N�f����i��u�B�9�Z~#	��e��?t!��¦�r��Q�}�1��S�񱪑�Z�h�W+3]�c:a$Bp�..�c@uI0�!���!R!o���s(��>�3!��!#��}��6�������&aks���{K��&\T40�p��7��>��~�U>�ۦ"I{���㐙��	��#��k?s\	�ۀɇ�f�ɴ�,��G���7s�1"*s����$	m���f��Bp�0|�u�	���.?\YE��Oc�gV6���������_Z��Y�'�O�eL9k�x������!!C�<��]�*�f�=���N8��e����5m�ds7v��
�j����GҐ:(���O]�Il��j��i�3�5a
�Y�̐���gq�@]�h+I���!y��A�݋����� �
Nx*(�!?�Qm��=�t�ď��~ʦOʻ����]��Ɋ��������V=���g�&E�{$̆k���ǒ�J9h�"ϔ�P�9|�Uo3��r� �R��F��Q�|Anu�tvf4|�{��s��ޗ�~TDX/�"R����>���c�YF".	�F{*�AL[�1C����cE�}���w��f�`��t�t�/�Zv��:�+���F>�G��{�4fF�r�Q�i��ZY}��}������������כ+�:|���$	��B�Qxj�܁��L���cu�Ux�|�Q�S��30�ʲ�6#r�ƪ��������L��gJ�D���]��^��͉�M�砭yE2J,��PZP��ʼ��>�C�/��EjۓG�62%ߨ�G�Q1�ɬ�p��� *_lI�g�f��N;´2	bה��5���&���P\�꣈�����
}��z�~� ��S�������۫�"�1�KLL�%����������fE�]O�]">�E�8����������Q����<M@ngg��F�x��m�KH�M��c-Kʽ��L�U>U�웩�O+5�������ڎ>������hȽh�!��>Bɥ]}��"eVs�Օ��#����<͒͘�aY�1|�.ol�}�$�mt��߱5��=�@�3�K "���B�\�3\��B]����(_�n�������ϩ׆��:�\��f��o�zJh(+/|ri�:M����ظf�U��a�M��e������ BO���b	^�E�y*]u��g����V7/]Dx��o*�;�K/�?h;�[�X��O�֤�kY�^�&e�NƪQ����g	���F��;G3���۹��}��%К."�R`��jmê_ �g�*h��B�(?I�w@`_'U4)����t $L�a=;����y-�u*�k�"�\�v�¡rlie���ܫ7��H�N��۟��
�k?h������V�q����v;��s�ŹFyy���Y>�,#�{���5�,t�K3�^/{4VTř_2�4�u���.��zs��&K��F=��Z��N(�W��U��g:@ʙ%��Uf�\�M9��U�
���Z��*l����e���e�Hf����[1#��n��H�C�&m�k|�a���2��6>/L!NI���H���R��Mԃ��B%͖�F��믖G�`t���.��0�^��!���{(�{,GWfA(
�9>:~��9Q�x�k�Yp�c���x-1���9xso�aG�eȉ���s0O�H�սxB{<[�ԙ�\�!E�S�������7}B:�3zG� &A/���K�$�0��;|[�{�&�aB
'P����R����|C[���A�B�nn�1X:�9������uM�������K�2�s�h��	%��i�B���_a����Q �63�]�_v_�E�Xa��"�*iz�m�D$c�������c�Ez�Q�8�fi,���H�Uv���׬�^�v|��ɫ0G�L8R�sy'j8���vwB�� ��n
g1�B���+NC�qK�)V݋�i1���J�Y�s�A( �E�L��v�B�Wa���]6��Fe��f!
�6�@��"�]����(b4 ��_�B�`�nu���b�86����W��t�7\9{'�I(�?�-���߅Y�p%�M�����D}�h�F9̡v#/��Z"YbnTɏ t�ք.L�BfT!�H�>�9\�l�\Y{�|�#?I�n��[J���G��E�&`�q�C�9n�+���uY���>	��E�QGǣ��E�*:#����w�B��s��L#��*a�X#.�"�V-�F��ST�w*s�����̤���ѽۃh\xչ�X|oMaJ85�~yiNT������Ly����i]#աY��
�YG�me��sX����'C4!�|�ۑn'�U}{=o���Df} f����E�{��w�;g@`�pȏF#!�J�A��}�~���S����E׹�;�9��z�6�f|�G�=晊ev}x��V��SN�B4"3QxA>90��޻��������cw����Ffm� }��"��	!!6"��j3rƓ�n��Dň��]C�9h�q�� �r	���)ukQ����B:����`wd�ʏ��d��`G[�iF|r��ӗ���Iz�$ɏe�d��ny�]D1~�.�~%�a񛖐��Ĩd�xNe���~�LPxXH�nv�/��.��3jm�iU���фd�6��H��� ����(�J��Q/�<e�#v~'�pDhٿ����}��IA�#�t����?{2"��e|LZ���>�d�>LG����<&"��UB�,���.
p�H���T>ɴoe�bbr�Er� A���:K8����V�E���z��Ԉ�6s	��N�u}}��[�~�=0����<�8��#�4~������0Ȇ�ْk:8Ci�`0��0G3L�#�(�6#�c�N�;��􃙺�P��Kc��D@��f�ȗ���9�G��D`R�ro�ЄE� �v��ٶb����"��\�tr�m*�ء�H(�����<c;�8�� `��>a��m�Ҏ|�����i�,o���L�����.M}�}Ƕ�C�cΚ�r�4�� 7���仫�5q\��:T�ۗʝ�"|�igXpeoW(�	!G��]��FWAJ�C�\	��С�Cŭ�V�����q��PY{C�Ź.;v���r���H�@�S
�Q��vv�-��YEη�E�hE�1�X.ccӭ݅������ �lumv{�C��2�Xõ��U��9��qs��r���;���F�<��g>s�$[��I�t-�Ûu�*�`�/h;�����	���r1�����+y�e�v��]n�^F�|�q�p�<�M>U_���I�u�q~�b4���+Lų=. �Pƈ�Ń�g�~��DG�s.�9�z5��@Q��}�//7g��6���8����7�
����H����rɹ�e�?pE$��J��v�u<��G���D�7',��U~SW��������G�w�����[��P0��m�p��i!ھl�S8�@;�e�4�2#�8���7�`@�[,�(��s/�s[<�zya�f�t��!anK���#n� &@� 	m0wb$���� J�Z�VZ�00�����/�w60>1��d0*[��ʃ�mEl��P�AH";*,w�_1>O����8�|R-��f0�?�q��Ro��\�a��K2Tq�;13��R()�cɩp(�J���"�^fE{/�WϑQ�8]�a�L0��/TM�x|DP���A���{�6�w��#�aт�FR Q�W&,@'������^�z'5�3Y}�޹���1p���ݹ�,]V�C%п2z������b�8bAJ��Q������g��І��3y3����!�/.�m��wC-(H�Cb�"�r4"B��[�Ue������Zb��w�XVb2���G�4���������R���o�yƶ'Дb�����,b����1��|>�/��F�m��!��y�@,ÈMɣ`�fd/r�9�f	�H�D���& ����c�쏗��HJ��~�@wna����͡@�����y_e�w(��P����
��`�R���	�{P۴�5np�+����ҷZ��,��G%��}-�}Sʎ�����4�9(n�ɛ*dz7,��~��ZG��Vn:�C���6aqbۮ����g�Oـ�EC����!m�C�e�N>>I�o���� ��b��B[�un�6�s�۫�l�rYkrI d�Ǎ�1�{vŰ�A�,n��ۼ��'^1��� AV�OP��"�_sl	e*뽗�Sq��OѢ[���*�3*xצ���  Fr�h�L�Zw�<g�����{hDfg���O6�Tb�	�K��Z��
�N���}刈��`��yw2���*M�9��/9����pH�"kޫn��aM��������:#�M�a�a7�(��6X��g��z��!{3���\1X���a?L��z�c9�A��ˊh��>�)��C�̟d������L,?h�nQ����T-���P*.x̋�`a~j.W�=K����	]�t�X1��ٮ��Lx3�-ɿ�>�^��n,D���T~�1~�q~�dL� A�c�9��8q�_�=�����vۡ�F!ܾ��0���wE{g�"�p�~c�c��9���Gtos��@��hő����T�H0���� �Owc�s��AD FX����\�PCr��;j" �ߜ�!l���
��Z����Ai�쯶<T�{��_<���,A����'4T�U}�U꛻�:�N
L3��&-�c��"G�+���꫶j�(V�(�.:;�G6k��6`<=�������d��s��h��N�6���yc[�`{'�1
"75�]�<�����g�+: YQ�~b��x����b��|�V�c���cN[iUe�gW�|�д�NScQ����ޝV�*�ٷJaP��&k/�p���xz��N��	Z7K���ym��If�:�g�W�����
�똚M?��a�8�K��
��uGd�B�J ���PEe�"�_5DC8 ě�U�R�߅���-n|��Uw�yx��7����=�͜��Oaߟ1�Q�yڈ;����!�>��fc�-.BP���![�3G��Ȉ ��P��A���6�L��{�W��H׶c��fOMӿdVȽ^��$�%шw��.���J��*��I��%�s{��$Vs3">����f��Y�M�sA�ݦ��
��(�o�;�
���%$�i2�˺<�25�tl�8-������������ɪ��"����2�s\�	��(B`Djb �!ҕk&|"l�{'��/�M�R���0�z�;x����B!C�����]~黹RP��(+[��hX�W(���<�=�En!�&�*hA�2TU^���8Z4[B^�T	���8�˽��Y�m!5�5\O���7ز����@�A��)E���d��#,��轻b�i*(# wӰ�=nyQA$� &H_���Oi��9�me̳��諵��DBp!�4�@py�P�;�N����qł\\p~�?k��1���SE}	�=��{3�v�fTA�>��aǽ�,�s����"�Vn����M~����,0� 	E6�4~��+]�Ra�T�jP��nvFo�}2���Dĵ"��y�8|%9�w���H#D_�'Ԃ!z
���,}������O��؋��R�w`��hBpZn�f"�X�9����u� �˟����MvٺM���q|�8��FF,��ޤ��H�Ӗ#�7ɦ�mܽ�U�V<�[�s�t��V:�F���x���t�F��1u�Cv�p��_uy9S�+��^��[�P.��Q�ٵ2dQ2�G�w4)d���Pl���16�<�>Gz���}�x��uj��}��'d�Sz�im:	���]�y^��#B䢥<��������O��ɂ����t��ܖC��K��ŋ'%��8k9��2����PsO�v {s��	ǥ�ˊc���w.��$��3]6��,�1���\�w6��ͭ��^�V�z�Y0\�/�`� 3'mq���"K�Ckn�:�ʛ;�*ن7�_�va�h[���fە�Q�EM��B���-���y��������c��읗ʻs;f
.½N�����҅`�7Hiڕ�e�`	eE�����prr�M�x�R�X�5/��S,��õǗ�Y��I��s�+��<Y�h��s�&�oĂ賒��7����J�Ӆ�<��	o[���9�v��݇s��D�.���0]Qړ�IJ���T����g=��9#�{F�>ϗ��>�0�12)��@"�owg�xf�ǥ�fa��ğ�2m�O��ۺǻ!�:��8̾���m`�	�^+U�{��	ֲ8�7I�R=��=XJ��W��ӆ,<��҅�n㐩s�Yw��K���4֪w��o0A�1��p)E.��B�o����$�m ��14m������{*�\�����0���a��{n���w��~�-Ծ�8a���̧Oq%"�4VQ�|��[ԟ�G�����p��h�?<��uo+�@/���4h`�g�����q{2׮����A���I»9���5��e�0���uq�?@�
���oV�eB��&W�Kp�_z)[���Dv�)���mpX�GB,��M��6�Ü�����@����K��/���ـ���M�)D!�E\�W\B��G��&��ME�=½�p��E���9���N;�����r�y�khdxze3�����=���"؂�2ڂZ�A�P���j5v8��Wwe|-ۄ#�l"��gj3��oC~K?���c9����;sϒce `fS�c)p.����V�m@o�R�~K���1z�J�?�ǧ}���`��j�1��{K�*&�ր��`�5�+
(0�f^�쨫2�"4��ɂ�2����)����������n������>=��_\����XKsz�R��q]�yo����'^����{й�~'S��=����ᬺ'���9_7�mI�qp$��s& �F"I�0���U�b]��zp�y>�	�L�XT��˭�"��#��2W�a��w�����+�&�ޕ�+�\�W��Ӗ�=���w+M�NBݫ��C��!�C���$,�}�qL[
d�W�E��Ϩ��A�������*�,*����gAy/$��s*Җ>�X�Q�X«w���.�]w�uY�%^*��Tڶ8����s�vd����Xĝ?�7�������fͷ$�<t����X�g�Qx���ő�]n5�^�<��*�C�m�ll��v�V^�����x(�N����!���O�m۟i;GBݞ�9��Dx�u)	�5�s���)aJv1�IL���e�j�j�҄f&Yh)��ƞH&u�g���[�m`�:cg5�>���1u� u/OU�S�n��Gv���Dw�5-���������eMx�I�� ���}�of0�+����O��B�U���}��?��a�F}21��{�^�[�=({���$m�5��D��R���T�*�s�b(A����q^��w�'��|��cF��<xl��^�]£�Иw��#pt�]�5U[ ���&Y<��Jo�����=���h#i��1O�p�:(@��8��S���(�l�d ^r[<�l���2�������i*���(�O҇hK2��� ��ekqz;*`
�=�?c<��p���:��}N�1��Q���)5��
����	4��w���qF?,���Z�%'�~�u���i�J��˩bo�2���3��2�X�rD�wf�O�iQ��ǒ�*1�S]n�v��pL �h��^wI�/.^�7r�a�*^�dR����f(<�"%>��[�ɲNm�d��gA��mB8u�Oi<����}�dJ�����Td�M��~���m���he`�P�mN�*}�x�$��pYu9�+%峟���{I�3��j�`đ�}�d^�DN��b^�\���;��O.�jYL�wv��D���uf���#��>��*�� b���"����g��y��&�ق"ro4#�K+ ����nz}9�$	�n	��y�u���?@���s�_��E"n!]��y[�r@X�[�=�2Xz�fQ��v�/6Xo��ұD�ط�^k�f7ڐq�6��ל�5�m�#����ِG�L�ͳXY��y&
�!�϶M���l��e����[&�^{&����0�
�A�oǡW�g��$+k	wŰ8NG�,dö�����A$�F�Îg�lx���V���j�\��
Iè4��cd����Ͻ:��Фx1����n���Y�g�q8��9���X�1|�wg�3�ȯUe���'�'�Ja6ɲ;�SbT�H��#2��yDb��@@/ڟ�a̫��(\�CT�FgT��c5���xZO��K@��r�;�;'�sS�ڦ!�Bi<u�fא�aqPm"��(+H-�FNeɧ�1�r���q��V�4�7��ıM�.�or�~_uk�d�)���"��^��!=�6߼�h�,󝴍�R8� ~��C��9��a�P��w�3&��w�۹>ϗY���M�?s�ٱ���Ј��8��X�/��s��>ɫ٪IK!��wk���c�/��b�a�g.ܪ��������ۉ�Ld���������/R�:�h��(����1���j=��3�Dd�U'2P�[����:5 ��8v$�u҉�@Z��zlM�X�ՍB��C�p��&._e�u�D�rp`�M���O�xlN������wr�Fx���j�cRQ�-(� �$��@I��"����Y������h8���	�	H��ٴ�p��0��2~��z�j��!ގr=m�0��b�.�TЍ�	M+MO:�͙���.$Q �Vf��g�_?z��)5��Fi���ʴ
�c��U��}�Գ�g���K��"q����g8��t��~ڛ^�
9��-�a��+�K^]/�z*&v��dT������NV�m��X#	�ֶ<w��z��a��G�Ww陇)D8�<�8`����U��"\�P�~/k�����Ǖ6\P��l&��ң	��T�T�n�Ͼ�����ϲA5�2��"ї��s����.c\��4���F�kxs�胤U9���4���mF̱Kz6Z�+�>�˩܍;��4	`6�������.n}����#O��t�sLs��3��Ƿ#�j��d�F���0��t$v�G
2�i���N��א��G�Ǿ�;�C#z8�P �`��b�7G!ڱ��8���c��z�*�2h�i3 �Et�mzsxLV6��MN�,�${]g�{�qb�5ȣZ8��o��Db���,� �ۙ���ȱ�{S5ƻ�߄� �P���"�l�v��w"k�c9�f���l���H� �a|S�ify�����6�G��Ҹ#4<�2a��ɾ����+��Uj9�dA'r5�B�y(�"Y��S;}�ժ��-��4��uL�H�Tnfu՚�B� �Z)$
}�y0�\��)	�e<�C4�0!��
Gյ�}ͯ?K
`[�s��Sj�fD�@��}޶�g�"ҫLf�E$���z��7���f�T\��ʩv224�8)��.=sȆ��M�=�̰����Q=���T�r��J	���<7�-���:�� a��hD�]�?��#�dMxG�����ˁu�kmg�qk���{y�0(���'�p��RR8�nۮ���~�fk�	����bNs�5�+y�C����d�F�F,w�n�2Y~<i����S�x�J}���l�B �e�0���<Z(�ζ�.�od���-���$+�Ԕj�{7�3c=[֖��V<��g٣���4����� �jz�h���=wJ��S��hJ잓j'-R��`��J�?+�9�l"!�Ŋ�#��a���].��̩�H�aLwVzۤv�r*��	�^��h��������o7�+�C��r��¼�A,�ov�yg������Ѳ�v�EM�	D�ٙhik'��Xp|Cisι\
��>0�����m���Qr����y0o�%�R�l��y�JB���(G?߮�&�ƏZ���
F�.t�>�8�G��!g����F0�Ex��V��ac�}���u�=���6l��&�wD��g�誮���j߭l*\��˹6R�8��﷯R���Y��1Fv�����==�|�)�֣�:e�nc��4z}침M�VaK��'#zX�1�[WLFdw.�YD yuY9s�1Գ��u�a1�0���9�;�ʊ���J���,Eׯu[� �p�#�1#��&ď��\#���4�3������$����J�ؾ��u3���h2T6E��=�0���F���z��=�ݛZ�H|�y,�VP]6�|?Y+���h{�ob��)˧^ؒ�	fZ�Xѝ�QÛǚ���1k�8�1�*��^>z{���o�ǚJ��ه2�W���R�a�8�U��t����ZVc���\���7z�7��3�/6���e�m�[��ѥ�����ۦ���U7[��1�v`��-� �#(����7XK���컃p��jLF�v�%�/m{4���LrYXhh�)�(�vnWfǅ�^.�8wf���&��ηn��1�9��	�27!��ٮ��n^�v��J E�d�����C��X��LV[��!o�&%���v���sKwS����h"�9�b�g�jE$#��,��T�{��1⺫'�.�Nxl����Up�gwɓc�l��x�[��Ч�����7����.����k�╸��B�'���`�0����mL2b0CX���hP��G*l �mUd�x5Ep�>���)p�����Y~�ڹ=R� h5�	�!@��wRp�=[�d�F�����<�l܋����v�o���f37�(w b��Q�}�Ż^��~�'�Tؤ��*W�e��WnH�z6uF3�����n}��V͟p�He��A0Ϲ�]	h&-,?O=�`e�R'<Ԝ�9�g{3c�c��i�f��h���y60r[#H�F�r��� �&�&:� �ފ�ʄ�0�����R���i��ܙ���pS��8�N����d��zdU:}��,hۜ8Ո4Ӥ���}��n[�(�8h�$b7͟r~x*��N���mF�Z3���w����:ƻ��'��0F��nb��Uy�p1��)�e3�]'ћ��4h�)NV���(����}w�L������[\��L�\jq����=�F
�ͪ3�ީx��+
s���/Q�� �JXH����3kz�8t�)���8%���a�ӕ�B�]�(��ٻ���t�#�����њ;|�|��e���?Ng����4<c�y�њ�l����sJ�	}�|_��JH��q�ˬD�e0�X*b!��~���._eCǇQ7�o�5��B�wG�Y�s����	���hh9�}Z�
pwo�`���$�h�i������-ʆ#��Ȅ@+@Q��!���e���hUޗ�-pF�惂Y�֐,��1^sle;mzE�ˉ��`�s-��l�Z�$�t��#R�����˪8��u~[ �z���糶�D����M�7�{�Y~���sv��u[������h"�ο92�PT���7��ٌx�ax!���W�w����ޒz�[��h+)#~?0J�}������T�_石?�A�:T-7��@�� ռ��{�h7�q�>:��,�oqtr�E�y:����7x"b��ٴr{��uʴh[�]���I���y��?a�^��1��.�^}5�	��"��Yy���v��Ezg�]K������D���p�(�9���C*6�g�v��}��*�`V\̏��3qcU�����f�doI��D%���q�@��x�\,I�e�c�JWf�zu�E��s���w ؈l6�*t�2s�p��s�Dr�۩D�N���ٟ#��|��Z~������U�zr�Z�m��÷l8;�д�I1��u�Ň���o@�eՖ�ɰn��B/ު���]�7y}0a�6@��i����=����̮�w��YZ���!�X҂�P!����{s����K3D�Lv�=���ĳq��,�F+���C��}���%�挴5P�2}Wf�4J�3*��w\	4n>�2��g#k�
�ށ�F��B��d_��r�T���bl|ȂC=A`����#P[���M��_{���w�m��]��wL��&�o~#y ���(p]�+�Xy�Ί����N�H&�!�Fҟn�fl3�yG��A;�qF7�t�G�3wt���'��J�=~�v]�q��?!y�z'.�ٛy����$B�	&�`|�4�p�V�˛�klx'���{��Z�������+-ǆ�K�#&Ҍ�}�n���`�6L,��B�����	GOw.�vfgǦT@񎬻�,��t.�l�
b�]���17��r,�e�A�g�+������/��uw�E]����Ǫ'�L�}C�14���d�`��@�Wɜ6�sO��oy
ԯ��Uk��(�$4S��hvD��������>�Dؽ��[KO<�����!7��`A��;�w;0��~0�W�<t٧�at�Ƃe=ν��3OaT
}�<tB�Z�j����G�b$�J��X��AZf��j��1�ڏd�)^�=�ﴒ:�D��F��^z=��v6Ό��ŧ�5����A��p-����0R �}���OofI�%L�?�㾻�g�_��S���7+�+�'>���`��^�	�'���rh���{��z�@��#�4�*eh�uYu�ʿCD.A�f��@X2����5�<ҧ&:���s�*p;�a@�y���b����a�+�qx+G8Ee�Y��sE2P�XiA�^�B��\�ʟq~�	M��(��δ��a��әu�@���/�7`��K)��o1��s�˖�F�G�s:Bݽl8��8f#�]�]L���}A��ۧU�VK�&�}h�TӼ��3��i�{JWc�w�C��*��(������g�������
֘�[Y�$�2}۵p�nz	�K�`�Aè�y��j9!<�*�����+V�,�m<޸�y�#"�0��(n�4������]�I7Ĺ�mF[GϪ2s�]���zh&*�Lh���Heug���.�S�
2nhI9�[��Xd��m��ʏu�o�{�����uf�S������,��Q�k�ɪ3�:C��zL�(Ӳ6�}�j<�XgNS�V��#/r��tO���۶i���U:[B��v#�.;��J��6,l!��}n�C6�����^6�gŋ<�Ṽ�g;-�I0Z��l����3{���%<��p�ӹ�x�<Xκ�\4Y��oO���#8�}r㉌���fب��S�wG27` GB`�K��b�4�k����qY��zU)^
M��g�Iw��˿z
q7�h1�k��Q�85�&1恙���KfDn��Xq�f`�[W��vri �j��}5��3�{��@�b]�����,<��_�K{���5!�&��J�>G� �ٛN�6�4�"+�B������慗�ZI����1��pO��J�����8��ISY���|=�� Ja �؋h!�0������fb��9��c���]X��_��9�S�~7���pZ�"��S��]�vä=�K��7)�>&��J��PMJ9q���,t���<�T�E��N�ή��^0 7��)�����n�Jg�4�&�vo[�(s��&�c���j��kD��KkG�=n�Y�i��l��I��c%���[�nn�s��+:1�����=�:m�»�2F��=V��ys�̀�������k	�6&�cxveeI�"G3@xy<t��>�ԗN=p�4�[F�ir7u�,6��Vz�)U�Dq��bֳ7�?��u�v|���Z���P>aWWf:26<�p�J�O�t���Hb)ő�jT�_Y��.z��o+a��R�Q��z����p��F5+�֜�٨�� ��l�G�qۼT���P}9��4��^���\�����4Se�J��9x��:Ua��2oy�M���������aܟ�OAD��0�G�����<��ꮗe�u˵lW��r�ɻT�������P�zm��T@"��"$Z>8�����r�Xs< �2k��9�}�,���DZd��3�� g��?:���V(w$o@i|[�IhPpo9�8N�s+֤��q��};sB����4]`T�_С��W�V���ׯ���k��Dl |��:����bW*_fU�h� ��;�ou�D�y�ˇvJJ�6b��r}링ǫa��d`�Q�~�����������Jȁ��1���l3��>���Yޯ[��N�I~�i\S�'|W�t��o�s�a� R��B)�l��j�V{)T�MA�$��5�[�F�ӾP�1�fkݘ��{C'��F�f=�B�i;�#y[�:Pe��U���9QD����#��a��ۦ�3�w$\2��,������Z���NM�0,����y�b'���|�i�/��ب�1��H��PA������M�W��"'�=���˒D&�]a�HH��b�C�Z��2!ǝ��J͑��Z'%��kQ��K9���3:��2����nw�ۚ�]��V��9:᝹�k2�/Z��}�_I�3}3E;��2�nQ�u�3-���E�c%+8�y���|�\8�C���3�)
�۹�y�[���������G�����h��b�x2�-�ݶ<m9��~/��Z��)Wx_w�?���+�O��r��Z`���v-�T�1N�������`�I»�췏_�r(v� ��J�a��'�M2�=�<C$��Ʋuǣ���o���yu��gp�HY
���=(6�n�!�7:ќ_a�����^xĚ�h3S�
�����RY�����E��)9��eκS������9鿟[cͽ���o��k�whI�S�F�i�x!�A4�ٔ��)s_����ll	�gzj���𐛾�|�͓Jd<�C�Z���Y�����_CP�ky	���[�����v�*qZ�v����1��Ҳ��J����c	Q�)�͙C}78w�tRy��No�e�����s�z�i��\>���7��)���!���':�à�ǩ��$�@(�+16�|'&p�Y�K��]gm��zIݢ䦗<š]6@�yF����߲��3��^٬g��.@cs!h�.�=4��ܭ��}�O8t$�k���z]����[���/�����~Y��N�R.��zq��ҷ�o;����v:u :)��e�(��Z���gi�J%4!��fx��N(�k)�;lj�X�IUx���'a#�ݴ���	���z���CT��o�.�	��.�ct.�����DC�Ǟ16�4�V#%����Yr��Hd��\�.�=k����Cc�f�k�攚b�+�Ŏ�Yi5��n��Fz�`��z�����y�Hd��|f�<�B�$���G6p�h�Zf-��1M�b�6i�� ���۲��F	��.��5�2�=s�C�d��U�i��zr�z���k��F�����=�8�m��"��Z�Y�����M:��X��7V�E ���l0"�%���y}Z�Ds/Vk���:�ɑ�&��6^�apC8Be�wZ��!x4��H����n�5	�A��a��ak�#���э�f��%���|���:�pnt1����C��諷��i�7]ff�:�iK��2u�A���\����,�+��t�Ӹ��]�n�|�A��,�ގ�4t��N� h{=7.6.0�z����ʯ�����a�rq����	&ǀ�fz�F�v�;��gҬ�=���+Y�j� ���ɉ�y6����b���G��r�p.ɸ^B��Ƿ&�]i�C.�v^|xAe7l���8٭��CD������X�dӵ���b��Д̷33���iI��Y�`�a�ڻc�E����jy�nj���a-MYFY��[����#\���v��莉y�d�L�-!��{	�k�GMxq�Ή0<˝�)���0�ZQt��܍����|_*�B`�mg���d��8غ�qC�^v� ������\)�	�#,f���e��D	��mعc0q�x���j���5�r�{p���0�&a����!�v�Z�WrxT�m�^7c9y1��#��v�O1�C�J���Q��f���].H��3��	�B5�S:VxK�Y������e �]�ia�h[no�8w���~e����	��\�{x�5�b {vMaۑ�.�:�-�g��u�_���]�vx]�ǩ�$�+��T�|(<�M�8 �0�6�^����;�nҕ��Q=D�g�hVp��)8(Cm�L"�5`[R&�u�53g��.���s����z��Z_P�����}o����9���9�ސ�z�<� 6�f�>��6��f�X�6S�Ħ�N<��j�5��#��κ4l�E�m ى#�	��i��]��aq$ڽ*i���e��1ȧ�� W/�#,'��Q���n��[�F\ܟ��o"��!�o��s��������*�Y=�饹Gy�T[e�i�"�!鍅�2q����IK��?v��a�Pe�F�����5ѩg�r�mY�qZȗaњU��Y@��X��;�L�y>���u2���-Y�q���
�CV@��`Q����rR��g�{�8�|I�����cU��B�q�뎕��%yg��G-��v��)M<�h0)���\���Ӕ���<dIL�&(C��Ք�;G!�a8a��E�7 �#+�<�k���Z�*l���Q�`��i���o<��J=�˅�$el�s��t��U~1������s_)ڦ_���6&bx�̉A���싴�'x,�mCm����s^�/p~�[������� ��56S{jq�v@$����K��n[O�(��m�m�5�j��Kr��<��=<�ɍ��{�u��u�\����\dP���z�
�����O_)z���YxI�W��$�P�g�W�m')����=-�]��z�m%#|<�cw%��+\���/^_fQw#�ti��kec���&w�
�w H��J�˻����&�=�OP�8L*�`�b�\��̽��q����2F��Mz�a{�T� 6�������a�ͦ��7�'Tq�Y y>=���=n�r�Z��~��u�8~���� ��%��~�kA���+k:eIB����I7Aå�*}��^�f��Ҁ0
�ˏh�����O�� Ыǲ���F�����o_<�9�� ��[DL�Nss!Ud���l#��q�����1��S1�>ں�Ma(xb�%�j��k˓Nfg��郴��ǂ(�㍿n�]�a�'d�V�V\��,�,K�v�k_i�Q��/k���/����ba�Ga�y��P�>��)uc�vW���ST�T�=���[u�Pω�<%r�:�}=x�\P�����c%w�A0�/S���\HK��hw&����]THȭ�|�E���g\�Q�R��x�׭
���;����ž㓌�ɡ� �Fώ��%�۬r�]�嘬83m�*"$���X
��7�ܶo�<�N&�!#V����h���"�'i8#���٬vr0��-�4�w��T���ۚcs��� ���L���G
���*�.�A�d�2뻧/ ��A�=�Pc��c3F�Mf@��s��"1sx���y�2!,���ճy���u�Ӥ��B��X��{�F�Rj l6<1u�M��n��_�y�^��>{t@a��ܫ��L��zN��L؂a�Ԧ����;8v�k&f6����[D�zu���>�u��Z���:$����Y3��n��{ی����s�{}Yr��p[�:������D�J�$�[�ELw��El"H���yE����R��f�ݎ�(��!B`tP~�������3�n'`W�C�Wu����1�>;zFo)������ 1PhϮ�����@
��8ֵʳqՈ�ˆ��K�s"*���S�sb�O�p 1��I��rr�P�`�(���x:w�*���J��>��$� ��#.��H�i64�웬�7��O�0����g����I>��l����AOe^y_�4:p�e�w�p�կ�S]���5g�s4^��d�j��Ō����g>�b�� ʙ���B]XXXg$*��1��E�6�j`y:���.(y��B��0���+�����|�>�t��+��J��,7���t2��D�+�8�oU/UoWe�.k�|���9�m�����!�̝�3�]��&A���Β܅�.��2 �I�K�+�c�1IIS�rO8�Wǹ]���kQ�`��z�پM�2��aW=��"�][�P]�p[
XE��D�M[��3�R��p�Ѣ$������T��^����2O:HW�G���:Y�G,����oť���F��jY�|����sy�&G��d���z���QC�p�e0U��G��<����܏���=���O|���"�F=>�ݓ�}IӿǟB�A���ˇ���{|�^�(.c6ޞ�>�L�'��z�������3�'��ܨ�<\��C)��rsχ��[��74vXݎ�(`�h;m1����	U.��%�f���х��v�+�ь�Yx����G	�K���鍣����#i�q2l�2���.�6�8ܗoE�ٙ�;Oq�/9F�B��,9K���HQ��*�K��ط(��eƊY���=8�OjS�[g!s6,�����mhV@BVY�[b �n�f]����8�.KL�s�X�>���`�%b�:K`����,g�\���H����E�䨯������i�Q�S��`8呉
덊�7�]o�p�l��̙\��n@fo�,;#;�è`ʾ��e>�\��سA������������NE�Y�+Q�*I}QUF4w"W"S�RI�����z8�������r^¹�m����sYP�@�HJI( � �oLۥXs���ڒ����Ŷ��A�[34���������{�}k��cnևR3��d*FE].��s)0z{Ш�g1� ���ލ2ٳ{:�h�of��pX�4�*��;j����y(T�h������Q��3��mz!�����"DFZ�����-\��.�|T�a�CI��f����Q�O�Xr�vm>��]֑Zv:��p���8�2+�}�>�59��v;0��A�����/��R<��E�CW�0����`����|V�����%O@{ҭ�d} ���"�bi���_lo��pa��E�Ejюa1�Yv%'c�2�X�3��s��9� ��dd�����z1g�� � u�G�h|\���bO@�UwQG����P�-$T�t��y�8��ZP�(.��Xz3�>��!�ƄOOW�+�7[z�Lv�& H��o�U����4��_��,{��^g}�M��O��,��',�������4խX�8�/�i�k���1Xvq�;��Y�y�.�&��*�S/����C(J�+B�v�����W�����C��1��X���<T򷶟�3b��}K�C �I�t����Ga�.�eZ۽|����v��|��KnRsA�
n#�.����[�v�U�%��U\��ᵇ5u�V�a	6`-��g����s2�����Y�ޗrh��1'}������N�"|��s|6D�}W1���!�I����� �JO�-FA<2����"����?JA�"f��RQC��?!�����a�K{���Q4<Uuu�i�3:~=�.H����ɺ��vR�c��!�K���������	��I�b��o\ɿXN�S&����� ]���>�c���(�N'��n�3����=��@��>�af�+&�(8�R&�R�9�����d��d�c���4�bZs�f�2���M"7�|H()�T�Ҷ[�
��Ec�������-
��]�*-Lx����r},�U��0�cP�+4"lr'fD=�c6.E��F�N4�B��ju��3:�3|E�Y��oo�M��l�)���	G���Y��º��j̉�gM�\Ӟ��I����W/��r��z6_��X7�z~�\��b�Zԋ�{��V��Gݙ��GT�
Z�g�}NFg��Q_�.�e	���8��{[��1�&K�T���~� ����v��G+�#��B�-���+&���q]\v9�Z�Ba�
�ݥs�#Z�f�HD�Kev;�%sV�l�z�׶j��N*A(�z�2ۙ�@��������F�Y�7G!�2���W*���ȃ��r��;��΁����qm�׼�@���P�υ]�~�#�0Rn|�ߌ���߶o��nH���ĐM��iº�L�{�g1���w<��[��(R�c�(��rͣ�B�=�um\���v���n��{�՞�x���F�Q�뿶��/�U�*�62Њ:���Uv=�@�0&��d\F	S�����a��݃��Ϫ��g.�
���oyߎ����i�.�L�rwb(�ș�X��Sc�����s����ڨ�H��k~�_F���,˅�6���9WsT�s�ގa���~Qz�|V��R��y�y5O?�)>�=Ċk1�����a�>���V�z~^�B�F�=��#7;A(�N(���&�Do�=�:������[���LƔ���)�kn˽_� ,Иx�K�4����[��ݓ4�gS�����,�����E���$���6�A:�Irު���2!=��5L
?r����1��_� z���m$%<s> ��	���f�O��Y\�M[ih���H�:3�z�u�K�Q��0;�3%cz�n�ыI�G�j�{w�z��jT���{��2*��[�gA�[�˃n�!\1�=�Co-���궥r9k�$B+H��ZeW����^M=gw��w
�*���MѼ�=����'*�t���;& NSF4'�Lwe����4�4�`C}E�j�:��f�����H�s�R�v�)>��7<pbN���<�X�S��ż3ra��:z�!l�8�)�+�=���k�&s͸(Rɴ�a��1�v8M�t��+�\���v[�$Pؓ�
}���n�����vl��H���9�u|G�Y�LiϺ9�)���L�[2�I�ԄwQ�.r�v�J��q��5rx˯]⬼�:�����܆�Y�T��O-ݮчĬ�^
���3���� r�Ỿ�٣��;~�.\�l8M��q�Lb���Vqo���xfv�����B���������O^k.��U0�)J<�r�N��X�}�e�K��|3gė�]wW
���ĢzP��&gٓz�Or��l��n\M@쮉���*_r����dd��{m#ztP�\���{Mn3���4d�l�����o<z�V砄8�j7	�~�[[��+k�y��9z��7�w���>>���B��G,�X>H!묝E���e�\�^�����a��p��ۊIrO,��B�T:��#���7�rcq=jjb+��Ҽ��Sױ�ӟh��_sy�ɸ���p�o����	Ꜻ����-C�E���{��q��ޗb:�c��~��=R��5]ǽ�`a��2������ȸ#�;X���3.��kj��r%���",m-�m��0i\�a&�.�NC��`��3��0��1�1����og��"#���i�+��r���f<��f&�_d�BSӪydf*7VzG�l��Ɛ�ȇ���n�����Ɲˁ��=�qB&$ߌ�-��(�ƘV�i,���]��%�ѭ�$��Pf�0�-K���(��4η�BYc5m�[DLh�R̙�
:͒��'n��ʱ����E2c��'N�6ϗx:�레�r�������m�0ڊ=�2�*�osn��x��[r�J'(��s�&h�:�KJ�ƹF` P�^�e�n�U*\W:�v�ǯa�[``r+ϥ�컜ck���8���<7�
k͞��v�>=��W�0�#8o_�����GQ�D�)�3fu�wu ���.&�=����j[����'�������-�(�j����P}��"��#�~Xa��������jf���	�,�<�r��㨘�޵�'{ G/������U���켧����ƺ��}��3%��:A�j0�A�D�ˌ�=
n���G��6�d��<;fY��>��foR�G����Pj�a=�	:|'��w��{�<�I�ͽضn�P�۞s��O�Ogi���
l����Q<�R���}�Ūe�:�4ML�zS��y�3$�)E^��:��s*�v��c<���.哋`����*�Q�������С�6�ff�&�]�2,.�a@���_B�Y�r���y�//�s�׈O7�C�w~βD���FǛY��v]��Z�}�0���;�}H)��{��R�[�T(�z=<R�����^�a{�u�_�Y�{{O\�μ'���uN�3����==�f�p���4hy���UFQ�Z.mr�y�s޹˛�oȨI �d��F;)�������[�� ��$i�)����
��H�ӛI�v	���������7���냌 ���S����)`�EIB��=Y��omN���6��ADq� ��a��߅�jfꩪZߞC�����H�����0Jh�n�:J��ymV�[C$B� ����	lJa��Z��I(:"=��h�t,�s��\�p��1;���N�uW8k��}����8#/�O}�k̿����B^�n<E�_:�"s*o�j� gn�pr2�א���o{mm���AAp�i�|��f�S�'+=����%��{�r�RҠ+�Ǧ��k$��zkA�o��P6Nf7��Ny*�l@����X}���i"+��FYu�As�08d��c��J���t��T�o�d�u�v�;�b[�+q���u�.g�[�d[�n%�X���^�-^��0�Vcp;x�p���ːVO7��67��)��%�{�H��!j��"ski�Y���:�K�b�X��J�@��X옞{��f��ތ�=5��wZ�oM�:��.�k}�GA0 ��8C���z�n9�M�s t�g�E%�3�K7=��->��5��Pz��Id��8��d��q�NY��U��#��J�ͫ�ۋ�:n�5�"&��ܪ�K��-0P%��_]�;�)�����F^'x��X?��V�O�?pXP!��e����&�s����'��1�Wٱ���(PKA@D���sm�M_|Mu*��ڑ�<������H�C6� �M��.�! ���U���z61���N�Mb�ׯ��=x��Q6,�-���5�>B�ei{<�;��#� B̕
�p�/0��]���~�櫕��x8?8��T%t�R9�fs1��F枤�4Wt�fd��T�L�$��q�}�:�ӭS%���-or��3V�<��w�܇F�1B�3�vz��{�ˋf��$]��j�uv\:�w4�\�W�Q�5����O���umL���viH�C-=澝�i��[���k��X�\��y�*s%g��O!U��.��� k���2BP#9\��X���+ט���1���*��s���Oٝ;��9�;�6%Tϩg��� .�R*��K�4�{�N�c9�Ӌ>��2Nn���aB����1�]	�݌������S�vuy�e�0��lX���K�d�k���}yc��4��8p�sÊg�nn��4Y]ƥ*��*{���̴���+�zT�M�f��6Sro���H�����5���1r�#�I\B7P���c�e�^���us�M�,�tJZ_guw��J�M��0fnSZ�Y�)��t�ο#���R|��9%1֬bXWnP�X�3�i:���A)��2��<ڼs8��˗�<邜ʤK��u����c�3��'#�/M�y�i��_�V�~x[��߂�P��+2Ը�jb�޼�q���,���P��z���k�{7����L�5>��ͦ_X[���	37�������(�w�Ӻ��h�a�IYT��zw�1�z�գ����`�l�h�?����k�P���e�Gk��+N�w3ra�"ʽqv��w�(,���3:�~����]Vm�;R�j�%4ӊR��B��ޤ{�X�t�O`̙�{��k�l=�݇:�^Mx�]��*��tҵ�����Q
�R��M2hn��+Aw%�U��;9�D�w\�VV����0ݣ��9g���5ՓgLW|�"�/�/o{����܇��;Z�9��c{��5�'e���I�ͣ�����1]�_d#Ə^ֱ�5UH3x�L��)�$���[W�ǳ=&"�0kB�ҕ�sHE�g;@2k���L}����p@~���x��/Λ"rf��h��Ԡ���"Ӵ�<�,0K��=BS|�{��5��y��3m2q�.#)Fw�^A�w;���A?i�nؘ^x��
�)��RѲ�9,��s) 3�P.F[��'b��Jb��{�ޏ�N�"��)���u71�����8ϗH�e�Rs�G�fվ�\�;5ʀ)
����1D@dч����YG�Gf���o���uA2�so���V�����IL�P�ͮQmtƵ��ۻ�4Y	~rC�;�R0,�{VGo���q� ������I�۾·�塜�-��#sP�ճ��)�K�*�X;��G��v*M���m�q�d��݃��@CxpXLs׼�&��&���V^
	K��;��-�y`S��ߋ�>+�/m,K'�;1�f�0�Km��ʮ�u���C�2iO*�6{��z5>ԍyt�*��˶��3P/� �A�D�Mj����2���g�hZ���ٮ����zv'y���{����N��4u�g
;�+����!R�	&E巸ۤ�*8#	�i����èMq��>�f�x�S���(8*�m�T����/l'�����c�Ӽ*�Onc	��� �>�9ƷnK!N 裉w,��K����J
P�F��K����]:���i��|0�@���� �f�yG/�\m<��З�ud4.�e@̡e�a/�tfwu�v��J��QYG�M�JB�(w��e=���'Ĳ�׈���!�*mtK��$U�ql�&�E��$���_��(�nOm��5�-�M�g>�4pC/�$ǆ֪����X~���1�݁&s�i3(�)7}��c�����t5n�e�OfːM��e�q�
=~TүgA���i}�E��b=������A:����>|/���q�f���Z���uWw?Z�d�<��\f3�Z�
�{���_�L0�`!�$��Ot���``2䰩	����ٖ�E3�R�,���A�aa�j!�jO�ve�il}��|8��US����|\�������g�r;.��mnx��b���8kKb�J��E��8�b�"\/h�m9�ay����u��Ա��YJ�hR#uW%k��8�˱v�ui�h3h2ۮ3H�|�xy�v����InІ^s�ά�Ƈ2���g��o'i�XF�t��kG8����
uU���8����[��`��y�=�m���v硳���ƍ���3���5��eڋ�:^�<쁲E�M��C)��- �:G�j�W~���<�^�{צ��3�5�ݘ���oY�]�B#�|fj���_g�P�h��-qT0�ǱC��N{$���=�_@�޼���ob��)ZN���7[)j8q�\}Q�,Vx�2�\�k �%��Y��^�rFn��A�!�Yܽ���K��ۊ;'�%:���b�8ڹ�d(	�2ꢐ�����
�Я:w[o�k7gA0e�N%�AjӚ�y�4�=�i`N�u��zD��+�	T����s
(�}���"Z��v��Vem��lr�Tq4ل� �3�bI���\������+]'/T���}��0�D����k6���l�y�z�J�q�����9����=�z����ݠ�Pi�S0�:���՞��f�����}<�f�ѻ����7�w6���I�oTzw8n{�oV?c]��&�獊nL��"j�[�/n��ł�WMV�կ|�:5���q�I���z�ٙsS��m�G�Sf���uez�����ba?My�{�7{���O>��uW*bz�ޕ�nd��5���tt$�" %|�H
Ya��}Nt	������̝�-���/6�Ibj8�/a��^�:����X-��'ӵ�%H�]m��^���s���qǡ�\2-�)o�������hܻ���z�V��\�����F�5�v�,�a�S֙�ߠ�Y�k7���sj��1�]���Uʲ� G�Be��Ms���`5>�L�މ�}��!wp��,��4`�� ��v�rF$���I��]v�k��c�k���,"�Q�0���r>����Q��ǺT
��M�T2懪�Ș̈́����;/���Q��k�>;ǈH"�)8A*�zȮ����Vv{�ӫ3���زnf*w��v�!��~�̍@Z��Ӑ/��"+��[��]�}�<+}�Nm��2ˡޚܕ����<�����&g��|󙗻�x�
��G��S����1Kd�(�ϊڅk�fL/.	�x(����kۄ=��l�9=��s�S���GÄ�p 	��c����\޹ͥV�8�V���s��}�]���vz�X_?�z�g{^X���3�܉:1t���@V#Qc�v��;=Yt�v�DhE�C!����VPԼ�`�p�p�l��޳d�-%�V��w۽����-�79��syS�g-;��N=��j{f'�����h�[Z�D
�̫�8n�jo��k2/�Pr��P���3}�soc+�A��;��!�W������@�d�	�4q�p�]3�\�)��ꍟS{8j랪g����y/}�[#�V@�v�*S����B��a�_Ot�אձ�7��yt^��Q�N���j/��.�����*�(*���ݲ�o1�yo��#v{ְ��s�7�#l)ϫ��]},���sc�+���
���[����d���L��B�77Tw��F]�o��M����1=q�;Q�c3j�ٞ2�"�<g=7T9y9��rj�ɥ�*� �>�&��� #�u��j-�ri�x��~	ρ�W����N��8+��ԍs�G����Wb��P�K|yqɝr����q���л����>V����]������SP�p�N��XV�l>WU~���g~G�4�Jb��_��oǶ�;K��P������]�,^u�5���Pe�ݰ�	��:j8���w�����l8$\6��W\g�㙏v�^!m�뫾���5' Z}�o}vkL����Gz��	]6N��@c<�y	�'��bVr�h�y�S�y4=��%rIBH�>����v�w�j�1��S�Jw,�#@�2Rd�Z`�55�[���a�b�]f�;[��z�_G��ھ��'wt��iUV�[}/�O���:�jԦ�1Uԡ��Ζ�^\��o2 �'a�e�0�Q��>>HR��[t�޳&��(��z��
]�g�0�Z)l�l�D%�R���~o7:�h�ٓ�N�Soz�{n���J;�K-�B*�/d�o% ���P�$W
fL�zꏙ�2�%"���9�*k�mW�o���!g�^���ϥA��wM>�ϖ�^u������=�N�J����5~�Rπ�-+Uy���Un��u�"t��2���m���µ㡊�S��S93y�K���E�CD�B��f�EX��c�Q㑇��:���=Fy��Ӓ=XWlX��NÿU�?/W�s/|��?�����x>u֨)����k��^r����i7	�U144܊�m7s�;�7��	���`�<�jDX�c�.��v��S=�i�vx�ŝ]�3�ÛX'�a.g�O�C�����r�hz7+���p�)���O�eMz�n�\�xN�5\3��srcz�����+	ݳ��g(�-���Xܜt\��y���9�u`�	@�foթ�*���I�7��aL��\]w�]�W�\{��D��F���nkwT���.
;4Z4͘�)V��cA��(��؂,���dME{IB���;�f�>����aYޥ3[�4��]�^�P�n�:Z;t�%Fm����R�y�a�D0L�B��Wb��]3ݓC�Cc��g"��'�񖂔wv��9k�:���N��������Dy� ��=�i����l�¾�3�x��Z��7�<�7	�Z,��"Tr�)��NܾBV�����M�y'==X&��=���Y5�r�<O)�zɹ���.w�.���������&��~��2�v�y�]��!��c�
�qBǰ���~���KG���ȯ�g�Z�x<-�۴m�[�I;'knٷ.��E3�[t�0Z�y��Nt�l�ے�}>���:�-���Ւ�l{>��G7�v�m�c�1[*e��VU�uZ�sĭ��W�n��X�*�鮚���JfX];5�1nLj	�w:ż�[�mˍ��y�8��p~G=|�K��:s7[.N���0�2������P���h��5�<3'8I��s�8{���N]M+ߔr��A.D�t��dd�0<��$��$�̒�e�z�F�h#��V��8x����9B����.���¼="+v���%FU��^ݚ<z0���#��WO\{w�6~a4k�)w�J�2^`�j�|%; r��p_��9����rh�)�g�j9�$tG�9Ǜm��-�xÄ��f�K��ө܁�7#��]��Rr��5�ș�)u:/ݹ�~�c��x#�؋�eߨm�ք���(Sٙ��O	�uuxA������b�R,`�0�����7x��CQ���[4������s����s���%,��4!d��d�G�������6��#ׁ�Uٞ�q����emM0z�=��GR����9� ��}y::}}�ՐZ͛���r��Y՛\�N!�kۀ�j6x��sq�L.uq�v�`�iδ@�X/�x�
6��X{9B�ѷ��$)�K��li�J�����\��l�e$��ܓ=K7� ������s��\4�"����n���ї�{ᬂ��O���s7�֩�]��T����,�{X�K�Xd?F�FF�E��}��T�>��f�TVi���oV#�M��	G,e>Vc�Ö���*����gκgq<#���ޖ�'���	VZ���7�74Q��h|��6U��!���HԾ���3w{���
�v|�?���ZD�X��V��G;�;!n�����pR.G�8nvOc��G��O�:�T�\&A>j��ә�s|LU���PV�9YO��ۙYs{mϊ��dhi|	hCͲqe�5lG��R��}���� ;r-��p�6}����Uf�{��(OY��{��)�jB�3��eA[`�B�i�G���l0�P����5�<&.��OX�{S�1�׹v�h�a9o��z4W[�ˆ�Tس�]��F�5����6�,Yw��۞�v:d@4�z����ټ��:����^İe��W���b���yfe��J6iz�l��Vi�vrfG���|�&����!	�
A���9���,��w��9�=y�֯g�}{�ب��M�����J������CN�G�U�خ������ܝ&��tT�,�4��S�.v!f�P��J`�Ef�OQ�Wv��se#�qE����Set�4�  �@$[syW�L.�%�^ȹ�u�҈%��n��ϛ���k�-��&�r-5��&o� 4I^���bF�|�&ѫ������ȶ��w���rP`��fr��#^��T����hJ����,�l�H}���-�ZR>��{�I��{�3Ng�{��ܧ�1w L6� �0����N*u��ufo���v���#uA���OC���4��(�v�����u^d�#9��R��Qv�ϕ,k9v^8�� ~�-"�ޚ������/��w�_�BY���]g}&��S�ߊ�+�/A��D���� q�����I�9���I+Hq]�c�v&rfRȟ1~(M�q��pӄ��	��EF�K�C̀���u��/��d����t;��`��p�
��\I��s�ʽ�/<w�K�'9r6�6*�q���Elb�u≩xgІ�i�(0@�߫&^:���͞�x���2�n�N|f>6�gnڙk/���VP����#8�5wM�S�%�ٙ�3ش&f�wtתNl䃄�"`l߱���Q!�荖/c�5~�O����`[�l!7�ڙvP��k�L�k6�tԑ�Lı���HIP�i2�^�k���S|r�"�HÕ���05�A��*���{^Q�*7���@�ttOb���Y~#��� �P��;�vgNA O��3ٜ< b����L(�K!c�)�:�9~�K{�G����Fu�^�����kEMS���罳�7`��4d�Y�85� me�T̅�=z�,�*G�^���x���1�����v{���=��G��]�:��t��~��J�0���vی4��3����Bu�~�j��&y?f_�h!}�l�J��D�ޙ��p��q�"75�M�t�Fr�}�}�)z�q�[��9��t��H7�	�m�|f3�^�e��q�7w�|�.���wYX�UW	گAo�����Y@� �;��C`ڤ5�y*_wa�v;	(.�h��in�M������o}����;yS5Nt�;p�˨���S�rq }���5<.��<��aɻ=�=�'2��؝i�5�]X�Q�H2��$�Iѫ���NE�s�Ľ����[�R��~xO~@��Q2ZT�-�F2k�uu��5��Ў)V-0p`�Pm `%�*��Σm�ƍƴ����y�=�x�%�	Sh-�A��,R ���~F�uU�'R;
�O���_�s��,�P3ީ��N�x����&�u�nM6���[c��V�!�k�=�@���y�z4�RvD��s�M��5A��0ZR���X���+��v��>��^�u<�j�}U;N|s��_N��E5W����+qd׽\T�������^�'�2�f��aa0��M�p���q��(��ۂ@z��op~�A{/�*�֫��� o�r�\J���3�׍��ᠺ��:�	��� |Wjx��K��w�jގѱ{qݞm�T&}A�˭5�����D��ק~Y��vN]��c7�Z�vx�#�f�2gv,�f�!H�A@L���G���.�*�g�� ���N̦�^�[M���E�K���4�ze��s���&Wpsl��s����]g:Ԭa-2Զm1���^�&͋B]�L�|�?��\<<ݘ���==���X���U�ލv�e^��r�t ��/'�m<5��C���h��j0o�e%@���������b�������?D3�Y����+��iZPa&�P�9��1��a���٦��x^�Փ^�Vl������N�����b�G���k���L��&�Pڴ0%�w/n��ޢ,�6</�Rtb�c�81}2MP��dD���c�c��Gj$u֚f6&��i�zډ�9��J1���L0�D8l��锶��Oq5
_`9׏����PS�]p�Ge�[!E?K�'���<�Sr�լ��m�eeg���׀�{�����ί������a���Bg��[�q�~=R6�=���1֯X�Ԛ��ڽ��e�����ߪk=3�B4Y0Z�5�s`�,s�2��o=�|o�+��-g��CԦ��6]���jZ���*F��/��gy���+B����VkqMql��_����*�M���x���Y;���YK��a^V���Q7��8�r':w���]&��>HDv�: �S�I���h��O>E���l�����U��$ �v��GP̙t��+���n���!2�bI���qLuZ�|�Y*��t �bF��CϨ�hˬ�"�9�� �uyh�:���a.e�ĵ5D̻���.m7JΜ�Vs֎j�ZU�����R���z��J�#����z]�=��-<��-�Nf����ci�L�b�w4z�#�^e}|��}$���q���;�=��n�aXv���y�=�4����n]u����ԝ�߰Fvn@��=�1{�9/�3�N?7 y��+�o~�(�sr�t$�գxCc3�3�K��ұ~�
-T�};v�ՇtU6������N�;X���ޱ�W�z���2'��pc�Wx�l�}���Xn��}�a:�?�*�W��w{@����z, hq�i��Y�����AЇ9Qzܚv���[k�y�7M�.�����W\�$�<}iC@�`����t� �ྚiü3��p���B��YrMق1�/M&g�ݼx	��	��K�̕�x�o�&�7�>�夤�ܵɩ��h���e���;�w S�ڎ5s���6]N6Y�eZ_�4��ޙ���[�0@죡��lr{X��J���U��`w�y��]mp��zd�5;��nt��v����gU���8{���1���F�͏��^�����D��r�f&����O��gkVC7��W�*�Q^L��o.��V�{�c�#Gr=��9�#�x�~�^C�,��ܰ��6������g
�C�)�C�=�N�&������S37�p��[b��sƃc��|v�:T�,^�t�E��4�!$�i�m�����C<��>۶� 7HMRY;02j�t�vb)oӞz�ڛ�]���f9��nۯ��vs&x�ce-x�cB��s���N��\��y������Z�Hƻs�Wn�v�zs�Ϝ�>s�]�լWa�9������n�kʪ�6m(. ��ia1�eŎ�1�s�,\7�N�l�ʚ"�f'���H�'^pwB�8��%��%烰5�T=2�̄m8m��ӫWb�rOl@F���j�Gmى������j��dݔ^���t�k�9@;maf[L6�)BB����e�Z^ �*m���NpsѺ��H�8����c��f�fN���Ҵ�'%����Q�������',jК�ݸ&���3R��5��j]ۮ,HK�2�9��ti�i1������6���_4���^�7n�m�9�9�'F=O/�����y҈`ت}��o+�{q�P/Yf�zm�Kˁ�%�R���X5���D��b50��8x���=������
8堌A��i3�3)g�`v-jt�c��Ĉ��e{A	�nd4n�ͽ�q�@����r۠�B<����ƶ+O�mZg�t<]h,u��S�����JS��X��U�53���>�R5�����G���ϏD�9LZ������^9�\s�M��vGu)'u����wdHN3��zu��=#��[4�Y7��P��L���1s����"=Ë́x����nǝ�l�okp��]�ٱ[��L]5lc�Z��h#���.�tW�Mn�s<��#��y�����b9��Z�-�2��,,�Ǐci0gd��\������6�T^\�XcYxf��=0%�Hh�y��Ʈr�p��qna�"�b �sh綉il-�eݱ�söh���8@K��N��HV1���l��#]��4�<̦G�j�c2ݠo�|���|	��㞆Ia��]<TƄX8�S6��kU2ڳ�]�K-���09���n�*���l����;��[���s�n��a�s��,����M&���������B�ebJ��x�'�ϕ$��6(d~���vwQݪ��:9��>\5�HϞ��O��� Є�>i��荱�ӌ���5"Ϫ�k�*���6U�:�=�_~�}o�t�G�gўL�d]ef8��=�-�u�A4�m��\�٬s����hǝ]
�Ke�e�
�;ϹBЌ�:�>ڛ���%1����3���/+��c�$S`����V�������L�OQY��ЪFI�h�oW�\�ᝰ�F0� AY�4P���*ܕ"	W���h�3k���D�9X��iҢ������7�T���� ��Po��޿(c��,竣T�}~���,�0�7@���WC]�2{un����n�!
�d���|ڤC>�����bU~���5u�P]ޛ�����g~řUc��	L �l�*'%1�m�~w���9�����ysz�YN�痺��M T�'c����|I5 ED�`y�e��w�6�T��r}Ժ�/Etݪz�9�
E�BE� ]��4�.�]������7�Ά`�7�K�� �(��%������˨�KG,�ْ���h��!� � L��u*�9�q�)r��q��jٟj�$`U=��g���y���f��c3+��ӥ��2�����l.�k������ڜ����t]�z���3�zVz��?�]��ol��4��T������*�0�ợ�E{5��q�x �sj�!��,gW�?�0X���M���گi�q�xۻ�<�{F�`�ʼ���k�D�&��n��2�`U��0�|'�sܑ�fMu]����y�uC��s5*�}�1��%$��z���A���9vU8�,�����x�O��S dn<ٰ4�u��j���ydw44h��8bRko9��\�v����)�U�˺�.t�������,����٦P|w�<��7������o9�	�vea/��^ҙ�dh����0�,��_�L�Rݚ#�mUe����Wv�KH+��Ww���xOӀ�����/��#
�m���S�^�s[~���/R˪Ш:���ԝ�ޓ��K�a!��E{]�o�O��g���<�fz��޾�Z���,B0�,7�oF�
��܎����3�Jʻqr2��=���������x�Tq��T�/]w��3^N�2q�;����p�G�c��Hö ϟ�����B�Zf
��ȥ�*�̴2�I�{9O�u��{=b�������j���v757�w/9!g���Sp���P���|Mb���.��sAj	FZ[4$������^��c�ezekr�ibٻ���Ćv]���TMi��d�ݙÇ��d^H����8d��qL��|�VZ<��Cfܷz.���K�y�#���2s�n�3��j��g���B���9��s�Is���	SQt,c#舘��p=�`�@8I�.�,D�ӷ�����d���{��r�}����"+�7V���V�ӞIj|z�f�»�m����w.[�lH�Օ���WB�&��N���(�����;�*�9>�ܵ��x�$��+�_�9ѷaO/"V�m��@֍eI�������w�q�/�sG���ZkgyT$���F`d��rn�&S��J��3|���+�垆)#�� "ЄPL���kex���l,b�����mtGF39���߿�x�f@;&JV�ں��XT��5�����N�t�ˤGd�[��a����>�e��J��*�(�[B����3��na\����h�ƻ�3��)5���zރ�:��zx��K��9��޾��N��5R�xy�íy�]�sw����H.:Ԟ�5ؚ�׾���J�ԙ��*-ۋ�_%�kLO��^�Ozz�E̜x�ܩ��;�;W���	ɺ�VN
�۷���Dr���@m�dM�zd<��#�s�x�§�Y�GtWU�W���t�n�{W����.]���Cx�_nV��N�e�&t���(*ݘN�͐���%@YSxnm,��iX�eq��$OA���|�o3(�R]�ʊ�-�	XgX�4��8���T�6q����m�l7'��ث[4 *��;U���h�n�p#�ݯ=�t�^�Y�aOkbY��k���`�D���H�Ѻ%6yغ;S��Ī'hʍ��o����t�:����$�Tu)�8ݮ ��i��k�F�	Ѻn �q`h�b�dΨ�-"��Ԇ��B<I��Q|��S��u���CL�.�3��3�h*�c]lN{wa�&A��3�i�d-�ٗ=��U�B�X���!�K"ׅ��e��,�d^�ɹ�y�{{_��\fd� �2�*��SQ]��b��Y�룞l&�A���WW�t,v��aR(���>�eA|9�S=c���ig��^j<Am�-��cy�m:f:;d�ˁ� B%���H8�Î�^)\.����{��u��k��XB���*�����J���1ٵ�/*Õސ�xuZ���L+���"@ά���Z$�oqP�4���Y7Vx��c~��1���g{�ۣ����^j�O��%��lY+ky��:2�$��>ӂ�Gj�9�,0e�I����Ӎ�w��#�/��-�*�(�Da��T���}.A���;�7��;[�4/4�<�6�
pb���l��ܛ����<p;����7
�[LG��`X!�v3��q�X����ب��jz,z�C4�J/�*k}ĭ��	lBl[%����
X&��7N���s��$l��ʵ��J6}n�4��j��J{��Z�qn(`��ӈ�Z"��紲ň�f/�'�rk�y]��u_b�X�Ý-R|<���[����	���|��ef'��I�Zh�'�㌾�ziL\f�B�`($�.I^Ra��WN�l��
�9���sy�<i*�Q0,��5��u^�`r0q
&sq�{�x\bc�����)��O�t�U�^E#'���ۅ1��3��7[�sM���^ˡ��.�g��΁^�`��(`���:Q�`?�@q���f��<>K���+X�8��9�������3���߮��8<��F��PtlE?{r��^;���h_d��t��C{�K�� �pH��w91p{=N����y��U��Ӽ�CO�v�i�ݥ���2fNm��;�>j��)`��Ӣh�<l�9]�� �/x��9Tg҆��1��%�a��q`��ŜR��I�� k ����V��iW��x���Ȼ��p�P�Z� V�5QG69ښ�ʕ'&���Z�3v���y̗|��;����M���Y��ۥ�9�ϯ��,d�%��/K�¡ѧ��X��Xx�X�\�~3�w]5H߁d�=W*�G<뷔;O"F��L󋑆��V�m�Q9����.�?Z�+w<�cRo<�9w`k���웱e�KLC�ef��^��,�����G�ݎ��D��ե���z���CэU�Ysg�����X�R�Ϙ���c�H>�+�m�tk��$����)��LE��S���{��˺�0'�����0P�4�i��F�;�(֛��c`� p�l��Y�Q{�<ޮ�>�2���s�y
�\?T�I�~��#<�ß	O�='n�Z�4�o/1���g��G[R30�i��&{9P�{�R���d��Ȕv �5�
4�[��15.xΡ����M�R�L֚���s/vǼ�53�b�i*�]]I�NK��{�n3�DXg��d����J��e��:�4I�xeY�B�ns}�� ɭ�R�{W�O6�)ꢲH>���5�w74�.��	��(4!Bh{��껏D����x�L���z0����L���
�;;�Jj-<i���X���@��*͝g24��ݻ"�y�#yw�_��U��bx�T4�0¨��Lއv��4G�-zP[�U՝]����u�w�q��y�N�ϩ�X���c
h�i�Ǣ�?"1`�� 	c'{�o�v)�x�� �ɥ���F}��4��u`�{sd�Wܧ��� ���)�>��Ug�����6�`8*G�t����/?"iL��M�k�M�_�#AcȚ��>�����]��5=>��b�ڼ+ޮS�G��~~=�zb��OBe0�MApP�fm�5N\�{}����[�IV0.�%��Jf!&��W��\�[��^���DN�ٯ�C�^����B|�&��>��[&r�D�x2�t� 7�0X����2q�����#O�l��g�|/��JO�	�RV�آU!@y�c�]�9�t�e�(���'
��ţ*�Jכ�b5�㯏1|Ü�Op�o�er��+'�
��c0��b�x�M�?N}y��	�c=Vo	�����L�S�[�7/-9f<Ǣ�s���1�X��g!�5��.���V��+@Mr��c6�r�>��CO�{���;�O+�T�
�T��g*�#�u%��ۆ���u���wv�b�; �'�ñ�ҡQ�)�};�S�69�̸��ۢ��qq��:�g�Y[ZM���3�Eʱ�*���0�1���f*�h��N��Ϫ�
��o]�+��w<.�񺽕�����I��6ZA_�6��0�޿X�T���ا79�8,ǈ�J9U�=��pȶ�/�>;~����'�&�<K�����P�I�uT�w��$�pLB,��OO.������I�.^�V�2�7�Z�P�xN�.�Fh���|�i�S1۫W����ʆ�Fq�Α����*u�2�ܧ%�n�t�S�J$�}8h�t��'����u�||+���=��$n��Q�C�_���2q��!4Ƃ/'�w�]˙���К�2�
�S����C3��{p�2�N1��}����J��=�a�1����!p�l��*@�20u�`����ivfcˀaK��9���煎���Л�8�O:��$7��8��<n���lKδ�m�0�\��-cv�Iy�)s���`�Ԕ�9�EΛ����?w�� R=�6@(;�=�����/#�kp��l:x�c	F�/&Am�<���N.;[�vиJ��y�$�����==7=Yv�J�MӞ��!g}�}�V�}S�k���P{kh��'u�Vj�V4=^W��G�{����9��@���ڭ��~��7�[~�1�	����I��v0�Oȑ�M��&��	J�Psa���m�J��>z6|�a�>�2;��u�wwǹ�PM@Pu����n�l�����ѧ�r���(���A:����{��{\<r�E��n�CJ�:32�Vk~ݛ�l�(R�~f]Nfky�ǡ�n󗑸���~�5�����!_�%���+����!&RIᬐ�1����=�י��S���#`���b��9ӈ�Fޠͩ�3˕�k�����YrI8�#ۚAH-��L�.�@�7���D��ݷ5�VBKƥ籩�)�)ի ����l�+	�1�܊=���g��V-�g�bo�8;Ѩ����*XMQ��?��É:��}�d��ɹ4��n�d��>$}�]=��-uL�Rwj�Ϯ��&i���[�F=N�uU˭��("R`��9Yj[-��+�k)�U��F���kh�
`�CQ9�2�Q��zf�'�c6�w-���d�s1������`/8Vn���y&�y��Ǐ%YsP[r��f���ll/-�z�EJ�o�0V���*sH^/�p��ΐ�U�xXлͬ�?��� 8(�҆�x��q�H��k�p���C;p;���_6K�wG5�x�s`��5Gjˎ��m:8<�-]��6�|����Iwwf��'�b#"�O��'z��;�Y���u;���l���xpwL`S[7�������i�M�$�L{yL�]���b饘de\��-l�T���!S;��+؅@أ.Ĵ����9�^��O/\�z=����&	�I�.�xWA���Y5Io���˳[���rɝ�C��=����1s���zV��[j*��L��Y��n��/V-:��w��jw�D[�9�$��d�ҋ6i����G���+��2s��۷����5o.t�+�aܙ^s�֮�Ж5+����^����? ��v�b(�L��gwp1�G�<�+���%\��f�p�ʰ���i�q���-��2����Ŧ�;��	�0�q9u���Z�Ʈc����X24�HtH"KTlcB�Vc�*e�8�6U�5�T��8��}U&�� �L�Q5��H�u73a%#���%�����6�絳���l���j/':��x��wz�D�]g�m˪��.̒�=,�f�����F�ѳ�ʻRt`M�7���˴,��K�:�꒯5c�A�r�v%;��-z�u>D�[8�¸��r�[#����~�ljl"�E$�$�j��s����y�b��GF}���w,��L���L�;Y$w�\�Õ�FS���]~��N�6����f�V������oՇcv	i-1�hHr�u�'�g6����>����#w���_�����'	�g\�O[���8���
�8�i[��2�v $��dմI���뫖#5�qo����8W ]NI$��pA�
:�V��;���|����%3�� U�i�ٵ��m/Eh�_�rf�Oua�������_G�}��@��$Z �>`����:��޵X9�]�q
�l7�5�Y��92��g���K۹��'��N�U+����*2��"F���no!o�3�{�GZ!
d��|�6�q���Y[�A5�(���,Ձ�!���Đ5(^\���+��[m(cJO.�u�kn�1PB��Ӿ|��c�`�~��|Mz}����i��X�*n�g����n[��w(`�<�ْ�8������ ��f91�=^��3>��8:�'[tn��Ƹ[�E���Dܼ�q�A�w���|G�P|=��Ԁ��ۜ<6S���dZ�e�~qS�p�44n=־�����ԕMF}�e#w�oe�������;�I����s%S>���{�d�(��\�ht�]t��р�/v���[|�l��дt<3t�Q;M��v���/�L�M�A�g1	��0��B^�vo%���m��=�G<{�9���n�'��������X�X���bY�~�<If	��U������Yd|#Tzi\k�Bȝ���+�2M�X�.�����(�x1�-C=���x�X�uT�K��:�0�=6�7|5�$��ҳW{�1��"�2w�kY^��������.�A�����
i���e�l?\�'X��eq�7u���%#���-8���޹���r���Q$���.v�:ۢ�T7�]2�Ln��G�t������v�Q]B*�(��wa9�ˌ\5��S/ST��=@�3/'�=�4U��}�D{��2�9�c�q�b��=��'���ܷ��\�0qv���ni@��.��5����t>�C�^��@h���phS�=���j�Nk=��2�҂�;5Ν�qu�D�"��~�x�b�sQ�=T3����b$U�	0��p{SjW:�c���W�o�8�N ����퟉�k{�]��!ld�~Ȩ%��矔�rL���@��5sn��#v�<u&����8l�l��]n��f<���&���1V��z��-Ͷ�V�oj�鱬��k:���Dj�ų:��N�`��^q��Y�:�a�yV�0�jy�çr�_/VJ��E.�k��cZ4,�E���m��7E�5a�&���~Ɖ�}D��H��a�ʾ8��W��CϽ�5���z� ��9��u�8���R<*7ؾ���绐f� �1�eȞ�Y�;��ǽ�!3�����]�#U)��{rۯ^A����F}{n%�������PYlnL`��"�À��.��6���Ϧ�i,���k@�*��{i�wgT�����y�n�Ó�I��sr���Ʋ�D2K$�\L�Vx�vjc�`���{�_4_u�����z�ׇ�zu�K���-�CR4�<��@�E]δ�R�^a�������#	;���Mx�j�Yۅ{��{"�i/��m�#������b�^kܢ�s��E��-�BX�ʡe�`k�lXkC4_��DD���@
�c�E�ܟk��+��1;����t
*emӓ3J�^A��ƀ���d3�TMp@t�9�xu�'f��N���S%ʺ�^�Ґ�u�Nf^�^<��!׽ٞb��<'�g���\�����?���s�v�}6�Ig��A���J��X6�mm?g�e�0�N%��^�I���\��ov	��Ex������(��$�-��wX��9���j��VZ��I�1�W:���O��a��("��˨ެ2y��opcmȕ��5�T��ƿ#V٠]��g�cR�"F����Ń�%��m��8�� >^�[�p�r�VnM��E�7���A
����f�����٤J!m�B���lc���FkRP��`�۪�l0X�n5 5f[Ļ�\6�M����E>n.�=�S�r>��NEն��3$� �s�5�@���r��#���9�zqI$` A��4B���*�\8�^Ǯ=d��S��R�J�I�)�̵�&������Lm�����췏�k,l�1�g}��S���e��gE@��"iX.1e�O95�c����G�9k�*{S:�>�~�·�,/��Ͻ@э "!��4�*:�	��sᤡ�}��ϣ�����*��7<��1gh7h��1��Ӫij� �A��hCթq�}[L7�u��s�>Ր#���j���#�wc���0�5uᵦ�5�d�$� �0P��/�;\����L��ᰮ�Y�����Cպ6��j���$�a�X���d���Lӯ����{7�f��+Xm�@��,X	b#=ޜ�fkX͉R�ʛ��=����կ�~yvQ>5�T�(������d/9hݥ�F�A��X���pN���C�#���U'�b���0�-��'/wdƙ��Yn��w�yZ�:�_ӡ�0c=����i�S4����w���n!�{�t�Q��^����t��A9�(N
w��v��(��?:J��"�k�x	�°���7v�L���}�'�yc�>T����7��}_C��tm��=�~����{�+���+1�(����SU���$�/��j�sO�{��׼��'n����Fe�?�{���J׽�p���t����o)�E�"��w)�q�O&�����{K+P��w�%S���T��K��B����:�8�\���\���\�Y7\�1��A��m�{�_@��y�QenW���G��TG��}�Piv�$�]�o��b�	P��FFE�bЋ�b
i]�<XaK��Vs�xl�3�n�w��������o#k�[lg�T�(��oG�5M�<������;��*0����|�z��-r>��n'Ջ#��s�`˜��*t��J�~/����jh�*�;��������V�-i�f���KuP�˩�U�d��-0�8�,5=��U��ly6K�>��X<vb���O	�c�tc�A���̥�o�r@lp����|3!������G��>F��	'0��f�98�J����x�U�L�kH伫lC�o�j������˟��M��^��o�yN��U{����0PS�8ݏSSW��4��
�j[pT�K+%�D]��-\� �a��D0J)6�e���[���P�J�����%�!ael�R(�a�K���Ϟ���2�R�/�U��|��i��'��
�T��ߵ�#<�k�؀�G?¶�8A�Ɵ,|���^]��^�F��grhx=�#��~�9]N�'!�a���k2K�^*z{'_������!B,�N48��2r�����pܝ��9�Y�~9��S"+zz�	����^� 8[�t��lgz�á_uz�+�0����M� ö/`��7�N�}�#��Xc�LU����ޚ�!�A�!fKټwk
�6$n�B�f�z�^9�#�˲oԨ���tn�&�g�Κ�^\g�K�,؝eP�ck=�A�fA��88�^����X�ڳ�>��p����Z�_��rF{����(0�m�K��5��y���J�U	x;8����=�l\�ޑ������]9��)�Y�8��L��n7�&�7x��=ː;�v���t�����޿
N�)�,��,_b۪�[a|U���B{ǁ7_�����xQ?3�`e����KY��$�erlU�":f�7��]���䖆:������}n��W*�&��X��f=�0'	v�Hfc]<�G��ײqJY��nz�n�݇	��4a'�O�E�����
���c�wdn�8��NF�y�x���r:��S�S�<����G��~9�:Ӛܽ�3�GB	�`"��;����nO,����^9�sn���܋�Y�t��O�E�zu���᩹��w(�;�$S��ٷ��Skmn���0g��/�1hA1��=7<lp��\�`��z]�`Ws�˖`�oE�w�='�51"����O��eb���SQ�7@e�	lC[��Tp^NzLr^ �G����i�o7}Y���`���֕h{Mx�5�iv0�W�&����-�c�w)m�0�J0Sb�'}w66�5�go+v�I��#<�4�;3<�؟kt�ɠf�Z���~^4l˰��U����K�xHY�,����}�#u�6O�X<ܳ�Ϫ�͑O�B5���b����LT�Ù�"���,&���fŞ:����ہ�=����+��ٯ�7��X.���[�BwT;�YOXwoL��+o��^w�.���گd�h@ƴ[ ��a>��ɾ��ܳ�n�?<�����l9ga��o���.��zR�U��=áU�;����p�QY���fI�۝2�s758!�_� ��.��c�h+�%���U�.�u�uߍ�[.�1�.�wrފ[�g1A��Z��T�p/aѓ���g��x���#�\}��.���N��l�a��mA.�Z������έӵ�%�Y{��֌�
����I;��4�3fn^��M�6*���gzK"nu4�<�&��Q�N����W�J�2�^̠,d�&�w���	+����6\n����? Yd�+N1�z��Ʋ��4 ���t��G`��/��&M3��Ƥ�ok�8X4������Ih����&u�����r�qveT�@�6�nk���� �Ṗ�;��u��_��n�\l��=6法���y�O$��Gnw�p�Y�uk7&���ȐVlL����5�i����m:�g\`v;����I�p[�	���vf��2y�:�aϴ^Cw��v//�����^-Ծ%��L0Ϙ�q��w�+*�C�4��v�N��P�,����r�U���/���4'�>�v�7,z7=7k�V5A��l틳5�	Z��$X�&��P�:��˝5ى��z�y�~?����VoG�&,-�%Y�e�]\�-���4�B#�����6.uw;}���f](=��P�q���#��c�M�2j����@*����o+ I��/F�k����܍Kb��R�ZF��g#�KO�)i��co�{b�W�����a���{�w�gj��^Ɂ�#����wR*�;Xdn�/O���	���M:��sO�omݻ^k�b���غ`�b�aak�J�8z�����-�~���� �͡k�V��^��x��`//ԕּ�-xD�� �?��<+ixQ���",����{C�/����P��j������L'gt,t�V��~+f$l{�P�<�^�kӫ(xY��	����*�IO'�[���fcd��^��^���8�$�R�沩��[�Ih��4��������1jc�vn�\9�܈9���e]?�)=�Ko�����>v�\,���tQ�g�!�;����#3)6�6 �[�.Uኯj�b����gv'7w`��Am�R�hB��]zP��0/F��Y>|���z���V+tͣz�G$E����̳�a� G'�4�,� B2L(_��+Nf��]"��~g���FpEJƎ%[ݵ7���YeV��{���z�^ǷX6�e%	���}��!xdŪ
(�-g����욘7���[��q{.��Y��a�00
�����2��� 8]�ʣ,df���C�hf)�w^@����=��\65��|�T���ʪG4�pkJ��9`畃�F���v�̹Z��sݜ�B Z�	h~�>����(���g��N<��^gl��v�l`5[TL�t�� #�Uk۸�;�m5�&v�L׍�u�w�_p�Ǯ�Ø=&�U������I�TD�������c��I�����l3��{��N�y!X:���g�����:�c	����_^wy4d���h��gA���/����h�[$��*�=��T���^^T�'���㼨ӓ&� �Qm�S�IQ�YO2�ٽ`u�9^�c��u�k��\�-�O_>{���K�^բ�z����X��c��M�\ԃBHl���Ԣ���2ۄ/� _� <b�b����E��
kDkEbt@i����!���]	M�Zw��Ws=���(�]�Y�p�+��L=���ln��Yi%�z�'�`��*89u�C/��s^����t�	��ʈ����3����r�`ʐ��r��p]�K@�^�B�E쇫}]��D�X����f�Q�w���sӉ6�d�@�<V]��U�=<� y�uo�]Z���is��o�0���^(�i������ӈ[CCxz��٧��,%�G��x�W��u�\K����ٝba��<28{:��>���K�.��gK��pa��[��5�C@�d*�.nkws�J��,�����ܣ�����<��}k��vq�g�{+�8�z�j➉����iW�k�%v-6�����鮻Y� �c��� ,C.2
��4ƃ��=L!�y۝�eA4wW�����	���@�6��m�W~=�cT;l/gs�[�K'.�x�� L��{��e���a�-l�{mx��\��ǹ^��`��~hlP@�e
��3~�l�7��	�;��½��?�{M�X���'�Y��Ή�s2�V�ۅ{u�g�2��3z�||�탭z�u
r��zk�Ꞻ� �l��e�N�2��)�E��_D$F�#�'g�5D�亝��*1��w39Bx�b;D���y�L ,�=�y�����;ʺtwc�糂Z��m���*Ə]hS��\CP�����V���3�*�z���T�:N�L�֝�)V?MwU����I�5y@Q%~�5F}������L��w8Dg�v{�,+gxI�Y�k�����AY�w����oԽ��XOޛ{��q�YL�X�L��Z�D=�
��A��d��{k1�����p��:�H��i|�����~"@�<��K�2A"Fɩn�ٺCt��fFipj��],m�[6Gj=0�޶������֛zc&xv�:�,6�:�e2a�x�m\/�ß7��7&�d��N߷r����)n[j�/,olo���W��$'����T�cW����hm��xmњ���6
M��Dh�1Zt��z�,X%��:�>ė�_��i2�+���d�Y׋7�܊��:}��&������;�4�pJ!�׳K�.�����QD?mde�r&7m!�D+��SD�A\��HH,w��nn��š;����8�~��@qS��w��l4�#D�@^�H� �����p����z�ȳ�{Ќ�+Z�8Rg
y�*z���2#W&��c����8�H�c �����*��y�6�-OŞ�ɻd�q�16�8t�{�/���.�����`�5����9�c�㎻v���]1�V;cvv�Cr�c쉓����c�ε����Y݋�dk۟Z���6�^�������$�����4��t6v�$�V�3�,�3t�qvH�WR�GX�0�ѻFX���Z�h44���3L�Y�cZ�����ێ���Ƿc�X�{��2�}�I����h��,{1�x�*��R�w�<�+n֪9��wT���>60_��������'=:k�>�8vq"�^Y,�~�:����{�V�=$�w���7�UzV=�&:ǺC���6Zϛ���S���J,7E�Z@>D�#�wr�v�	����o2�K�����W���4��ke���L˹�Y�Q��p�q����0�7��-�^�ڶ�	��EjH������S�Ǜg17�}�wrL��nm�Ά���]`�����J����L�f���E����Q�-0�Ӣjn�h��ԃ96��lhYyqqH:.�{�XS��w3���=`�d^#��S�a�D-,�0�(���H�G�v�S�����]�oR�뽷�Z�h%��j�9�	�;�'�Fi��-=��vsV9^�X�
{-��m���T�| ��0�	8
,P�##
)L,�s�ջ4�m�7C�	c�c��
�'���S�M�sA᷐-F�x�6�Ĉ��j�C�2��W��sx����'t0S�D�3T7,��*�7\S����D��VfE�b ��vv�1K�5�ðӱ���~_��t+���{Bި���Sܯe�*��o�)߶ A͊��[�Ciw*5�Q�ُ�<��Zg��Z��{�ɜ�J�u�ڑ�|r��w����'�aB�=��⌃ő���%��ް!�`~����,�Z�6����l�Us<'>����3�&b�g�G�&���׮�쩥��Ϟ$s�w�ny/5�pR�
ci�Inw%��t��"��z�)������2�{��<H�:�ä���e�Ǖ�{0x�6_UKν�_Jl�Y)����|���#�_�x]k�"���驗�I��A�7���x�O֯�[yz�y}$,���9�s**�*���Vrr�r�N�*]�J���mt}��O{�X�^3:<�Q���)'3V�)}F��Y���۠����5;�j!��IAʎupqҦl�v�����ҭ��d�u�v�X��S�7WZ��(�r�g䳷[�ҐQN7I�H��֫�+�۫���4h}�kl��� |���l��N�o��2�]l�i�F��
���$�:��og���u8�m+-��˾!��ֶ�ue<�6��A0�.�����u��VÚ<�+zN1+[�V�bثw����Y1UZ�������Z��d�P9����2�1����&�4�Z%�y�s�
oc�Ou�7�cڒvn��1�7yF��%��?F�ս�]��M���̏7-���.F�/^������ƷYrJ�\�0���>]��2<��mkN�HI	�]W�0�D���wH�X;^x:�0U6�lFwlF"�2��S�0���`�n�k$Q�����;Î)���%x-�a�������'E�;���İ�X�G��s��57Ǟ�M�n_S����GdN�<L �件�7e���t6��ᠦ�q��l���̥h2����5�UL١iLlk ����hP�˟>�k�f�`���b���/J�5����ƌƘ�e���ͱ�՜X5Mnс���'F:�U6��ۦS/;��؞;{��]�θ8��m�����Y�B2�,�Һ]P�Yl�q�sJ5)��_:������(�y�r�a�q�ҳh��.�V�dU��(���[c����mvwY��ǫG�R��f4��-�z^c��'Dk<Xf':��6��䇠��s�y$���\�$V_<���Ȍ�F0��Y��ӵ�F�[�]R�Rщ��P�6s�َj���!�{Y:�����l�s��x�D�2t�n�v,
:%��(�	{W\���.ֹ�8W���W6���#k[H�nM�N��u��[+�Fmڜy�Z�9z�L��#�vM���[ݲd�q<v1��nBj#�7����X��."�
LX+�e�.������9p�^!Ǜ�y�Ю�`�l[�)dH�9]/kq�0�fj�sq�����,З1,؃-��:-�T�����-���3Kn��އ��vu�pugoe���HFV��Ы��r6�=m
�B�Vdل�JHl^ml]��/�'8���հ�-���O�9�R��g����������^ؗx�s�1�N�wg�c.@��SY��;v0�\��nGGk`��y%GՍ���q$a+i[N�M��\#� t�pZ��O+�v��,�l[�7L�]	�̧��S�Ű�i����X��Z�W��������tlv���z�,�2��5�.]��ٷ'Wx�G&x�u�E�k]\-�F�8ŞY �:�ݹ���*�QY�����v��~�U%��ʭ���\� ��jRday��\�
d���bU>��0�1,$NF�+���t�.�+s\uB��r�'+�q�1cT�0��w7rk�A��<}9�%��5k�M-)�ͻC�oEdќ"ۼ�꫉yf��J�Z�ո~X*���O�易v�Pm&6woFӣ�L<t�ƶ0�Ƕgr����(��9A��A���]��ĝ��AF�(����߂�!���~��=~�OA���Y&A�"���֢��y��ۛ�6�z`37=u���l�;���#w���6	T���l�/.��8P��|�[{��R�ZyD�.pI�C`n��f��:�t
�o�-55
��Fnm����0��� �i�YQe	�{�Њs��z�W��&=y�[�sd���;nwf�j�a�D�ڨ���?{��7e�Do`��m�@���Mm�a'K�
 a�lx�I�UgRsmK�dgs�?�o���vB<i��/*�u�܃GO�����#��団1�g�B
<���ҥg��v
�-�T�3h��`�8�.�k�@�,6|��I��������f���ƀyD-k�<�K
9�*��]���)���LI�B�o"sy�V�^yΒ�k�(n�$�X4,֛"	��l�V�Ξ�o�y���w��W�L�d]��G��F����[YS5>�S�i�x�I�^��	��a���`Z6	��2,/TZ%�R�:��WL��G��IM�7���r��rv�:C͈iٴ4&���<�p������뜚u���l6N� ���Q�;u��a�0Pb��؝�B]�~�q�K�hv���1b�+�F``F�;6��>2��[;Gr3cHPZi�Y-A�p������A ��X��1�K��~��Z�������]���u�����7��Çv��D<�嶅r���ECp�!@7��DNM�fD�6ū�2N���0iE@	YI���`�(�0�#�Efʹ4��y Wiu,�WD��y����}���?x�-�ʃ=�r��������+�]�]��j���8����z��рb�%&Lهv�f,�#�yRY���,i'�&�i�(��Mjɇo�4T�����^��=��m�1���zd��$�%H���6���YP�d�H7��T㐡l�K���r'|K�X�w�C,ě�Ϋf������;��\����3��M�;G��1�=O
u�E���7ً���dÅ��=.� mo_>~e�xZ:�� B@�[��l
j�]0!���Pzg��J��qK�3{���ߚ���i�K���T+@rg�>���� ���z_VI��N�H�����g���3�#<
����7�uMh� 5�$�� -�q���-R�����SR������<������iЯ/���śhg��ｅQ�&'����ʃV*����+2��<	�@�Ae�Xӆ� R��{� �ԫ�s�ۘ��C�O=�}y�_��4��)f�,��i�k��fT�k�@�pa��"�D �	���S��v)�E�xp�/�u�{1X{�;�{��ӕZuY3^^�ѡ�*�Φs��(<ma/
��(p�N��s�ż��͛%�f&;$�W� ��s�ޱ�Ɔ˼����ڒ4Mku�wV㬪�+�p>7UxpM�2��\J�h��1�����k�5-�5�w3��#Gi�cȶ��_�A��o{��WP�E"b|w�,l�MƦ����j*�[ �D�u��+K��a�d���7�����m-+}����SCY�"&�!�h��c�y�C�q�םCS���~qЙ���j��&��;�n�+��eOщs{%���h ]���k����1)��s�qu����..}�<��K�ɷc�x�r1L-�E���W>u˚��>z��ӓ�j��ChV�VY��х�Yv&ZL��:褧.�Ζ��H;he���79R�+�5�a�5u�����[@�<\��ҟ�V^I�Y������3�K����9MnW���<s�����W/[��`�Ŷ�b1�v3��{�<!���=!W�%�XǦP�.����<:���k��F ��*N}�e �'i����B��9pɨ��3\�>��.�(=���w7[&���qR\���x�\yt�{�gؘ-�
��;�2$qaW�d��-�j����4,^tgc���nKcrAG ��.�9�m��Ů�ƹ@42�ul39m����������j�/�5^l���>eed%9�c(B�� �yR�
�E�v��3��BE�a�'���ݺ4��|먵b���g70]��j�Ҋ̌�@&��������qe.��RŪ�i�1���b��ݞ��5^���2�py�׈�z���<�i��m���f-C�)�-�㑎�m�6�r\�z��T�.-t8ї8kb���7��If�^]��3.�y,��:�\�g�����|,���*�n�6TK9wot�ͷ�����,�nJtK/l���/K����t��FX�xrGnq���fu�Z����ۚα�s��},-7��#)E�؍\����u�KM�U]l�3�5�_�xh��3|S��b��Ό.���YM��Gٍ����1��\=�qS�"�( ��_K�e�*�=�Qc^\:��=xPWuշA�[)����b����c,����Z���T\��7}z�R������	��h��ǘ��`�����g';,�9c+.�9Wsy�}{��
�K�w�
B��_7ذ�6b�x�K�2p-�h��'v;}�n�w}���,����?2i�[m���s!��ce�m�(�0�9p�IK��le�Y�V�^'�S7pr���q߳�"�a�an�R
��6�9
R����?v�6Om���|5���A��Fc�ʅs$:8v�X�YI���qA�q}���ð�bI�����Ɩ˪x���zp>�'ך����\�A�eu��`�zH���3o�\�:`E1��b�Ш�^���l�I�d���@�*�0!{a��g=��[�O��>oq��˱�{|�MU�����<u6�-�HM�ߙ��S�D���z�p� �=u^g�Y@!4m�Q����	9u����p�a� �h�2���ⲇ�Or[<ޙ��K#��k��7�W�B](S=�-�S��r���&��?�T��.͌��"�c�{����v��hwAi���)�)/4�)��Kw$�~�9�k�'o)�2Tylna��-E!�q���r�U�YWK�;�$�
�Q��V�ĳ�ѧ�v��8���wG��&�3�v&��l{b�Z��+���D���N��	�Z�]������Z��N���e33D��4���?c����F���'7��U����R~QR��&Z������3�w.����V���m�<l�ۂ���η�y�ف	0<Ç�N�6#y��w��q\�9�~<�;�\�
����v�����Y�-������{��d��dLO��`���J��ng�pΫ��nfw#R���oa���Y��kr�w;7��G�6x�̣W��\5@%���si��N��q�s�QB��x����9F��u�Iz��0.���r�fcZ�;�d�ŉ]0i��Y7Yr�B���{J;�Ɖ��_	�G��8 ��~8��s�SK}3}|[���J�?�$�H��8_�*��n�^,�O�(�'�V�4e��72�o��c�g���o�b���{]�O���E�)�XT����ݑh:�{�DW���݃��q�=�`ŝIr����uA�4�;����z�9	n�\��xr�&�˝�h)ƫ��|R4�^p3s��>ϯ_T4؁ll��suy4�6��P�t �>�<A�m���x�m��:E��z#}���o���u�n/(}�g�@�����W��w-���yx���<a,#�e�c�.{���W�nF�[�=��p�2wfX���խ�1ܷ0{�˲��Ł�
�ڂ�3�>󰝇���ww<S랬�o��t+�{ӳ�ں�ǝ���Ww.�S]���S�bU��Ri�@ܥ�®i��#�p}^��-u���6���U�� �gd���zM���A���R�	�vo���,D�[�[T�тv:�MfW�z�洳�ekԎG	I^%���A�F,P�jE���h3m&�>�A7 �ۃ��=�V=�7+�v�,+�;���δ�
��Ð��޴]f�2ل�ƴF-�*3��R,s����*����4��0�� ��z븤�[g�rc���{ Nx!Ύ#<�=�x�ۥݼv�Ĥ��m� �KZ4�s��a���G����GZ�F�x�)�	�Å��n�y�s+�4M"�z�iZ.����p} n�q�٬��FVV��*��������go)�[5�&������6��&L�(F2�����u�(�&oN[����̼O3ica���|�hIo<��ty�7���0LK�n`�(�&_8 4s`;�m��tf�(!�˅n�̠��T12eO_~��ᓡ������v.�=��y�/A��w/����<<^q��M����[��������ov����6_�Y�0���]�9lf�M�:t��k>q� �e�&E��zK�U�w]�����;H�<i��f�f�_f��cIձ5�zq��:>ma9/)��t�����,c��o��,B]�!k{7��z:K���7+�fKKr�}�ж�@�:�gn����8E��g0�sk��G����\�G�2��V�^�gw9����_gv���n�P=2�=@��<��".��)�����|�&�mC:��[z�W���Nlc���ݪù�Z��m��֡,�w�0�43h>Q�[�r��K�s�ϊ,AE���e�*pn�T�1v��}ut]��V�ӠUg x�â7�m1^�l뱣�m4�U)q��B��خ!�N,�Ø ��d�ݘfN8���󧪻6'�(�(3�_uv���q��t\���|>Ơaf�l�_�&b�[+��a��>����;k�U���ܭ�d�Z�9�3 ]qW�K�� ue]
 ��Wqj����P�|�}��GL�J0VJ<�eV�#���v��]m=� }ڵ_���7���o4q4l�7�+�sS��ۆv�ٝ�,ޭ��X��Ӎ�.ѫ�j��?:=���n�ǱϊF}���l��X�*�i�kz�򁘖��}j /)Mܹ�L'_~�;��^��s������KN����aE�7�C/�t��cEb8�/2`.�>��`����f$5����n�a�!���#"KX��6�����X�X4[--d�ߌz�c����4a��yy"I�̥}�`<�ҿT�B9�,��mL��$:#�7�ؘO0g��2�66�9�s{މ�Ær�[Wg�}w_��kcβ��9��ӣpv�X����Li��}�D���X�E��֩e�#�=�Ri��gk���~���}ݰ�5�{�,�N"��;/aM��?#ys�n��MΜ8N��6l3[5goV�OzP���4�Z{��f�t�SZ�@��v��yI;�	�WB��2�6c��`���htjo<��\
�5جV�1j��צ�`���e�x	bɄ�(z�`���6�{�Ҽ�ۺ2j�ϘU����!g;J���z�ɝ��]�S�W/)ɖ�>C)�"�p21�T �U�x+m��5A`z)�烱�x_w���q�rA�b70%�,/���ҭ���kn�޹�6iܚ�8�Gو_{�H*����y��kc�-ܣ���.�(��c�F����x!�>"��E���/�uc0lz���HRm�ɝ�3n:�O/�;�������7���vC&-�!�AWr�?��2������������$�N����I'ww��I$���i�I$���I$�����I$���Ӥ�I���=�I$�������$�N����'I�:�$�;�;��I�w�wI$����N�I'ww��$�N���I$��׺I$������I�����$�wwY�I$����I���gI$����N�I'ww��$�N����I'ww�t�I;����d�Me��I�}�~�A@���@ ܟ}����   4(@J��    �` ;����k�o@��� �
 5"O��{��� �'C�((Pon�O/`    f��  S�   u� 4    h  @ 
� ��@ h  �:�   ��ϳ���z�n���w�Y7}��q�ϽϽ���;���6�޻�wO���|e���u����6�=������ʒ���w����^�/om�U������_}����g]M��ݶ��J�<  t P P ����=  = 
��`  = {����   �.��K}���� � �������������G�}K���]�G���=��=i����E� � ��a������z�۔|l�{�^��M�w��}۷�.']sUQ�{�=�=�=�:>�z�����t��۽G�޽5�u�{�R{k媎�.;��4>�=Ǫ����ow{����t����5���*�7��  ��GU}�j���u��:�cz`u�ob���>�}��ûWG�˽��.��En�v�l��F�{�$죽gG�>�����N��t���B���c%T�     �wc���w�������/g�zV��뽂�>p;�N� ��� 4�[:t�Þ�t:��<��}������  ���^���|���� P)���{>O�w�= )�w���`��v�=î�F��+}�={�os{��N�*�    ��]1���v�ݷ��]�Ĺ�r�{�x�m��ہ�Ӭ{������˶:��6�=;�NG��{oV��H��E�   �w����wk�q^F<�6�}ξ��0��}���}:�o��U�E����_{���gp]u���W������Ǜ44�"X    ���z�>���tGO�ݳ��m�`&G-:7��OMt���7����u�$9�mm>����ﾯ_]}�U$ �� � ޻�k�i��\޹�=�4�v�w������n��o��ݜ���/�^ؾ���>�Ծ���=��o3Ow�UN�����{�N�jt��W` "���R    j��	JTG����&�'�U)�U  h �~i R�@�`&"��MQ2*�    JzD	*�����d�O������j���F�����k_��_�.Jvz믓4������>�((� �œ�@(��*������P ��EUQEV�EUP�E ��((� ���� �

( ?�'���?����������B-?W�m�Lf0"��^12���c�X[.	6<sJJ�n�nb1���;M]��}yY�A[
�����Äy�W�6�ݛ���*V+wy�M3%7���5�KT������M�x~�-�Σ��á��T��wr�re��"�^e*�3w8T��<k4Ҵ���t��٥v�V�28����W�P���}{8]X��M1�x&hR!72[�ZЍ��ܟ;˪���u��<��ǹ���:۪c"d��[NeŦ�Tx�JY@�nf���s!jT����,���=�;�U*�2GCJ�T���;w�r�/�~�jQ�V��MKR���g˩AU�g,aF���GCx�i��݁��b�EUkȣ�N� ���34Z��v�7�]�]n2���ևuJ3"Ij����F�pQL�7�m�k7Y�΂K�p�,_�yd��GK�{/��ڽ̷�	����˅?�%<���7�����K�\dU���-��r�*�ӷ�yyo!��S��'%꫻T�%*W@�]���*���gK�)K�Y���Coa=NƆ;�NZ����͎�fWp�Ή�c�f�����I��u��k&�	�ħ�Tv�US5ʂY���p�A�WYX����9v2��,���6���Z3����+\t�d�s������.9g5{ۢr͑��0�Ы(*��tf%Q��e��5�c�尺�*SMB2񯜋��a�t�)�{�
М�u�Gbә���e3,f�ee����Kkj�b�7L�b�z6��~x]#B3m�ݒ�T�%�]���df��`�ܛkR�1<��Yī�	�Be�,��&�wH2)a7/V^��xSi�'+U(L�՛�]^h�v+�7~ي�_�.��:N�0��(��-J�겱,b����*]a��٩����ʕ[/����*9�&*�	B�K�ț+
��eh�l�u�r^��5A/h��wWn���ͻ<�WQ�����b�s��Jɦ�)�!���ģv�������B�7³�ӏ*�*��u��W{�!f�U
�Sx䑚��e��%<�[�{��!{�[+�
�*�4��bب�e�n�3P��+_eѢwi�S�]�<�ޗ�ْ]������u�v7�����U�!{��f*ڐ�^
��ɐ�0v�������z����μy,nR�"�X8����yYs/��l�$pfp+ R�_i���l��H���5V�302����h�J�-NZ{�+.ڤ�j�����.����8�7�Z�l̪z��;��k�6e�L�n'�A�w������v�u��Eއ��f��(�_إ"��
��c�s�YdUnbw��+B�;�go-T٫v�Q�J
���t��L��e�����A1CZf4�n[�U������N�Ow�ȅ����&U�7A���'X��*n���͚6��ڪ����`�]&�w6�tv�9��-1�_D�ƫ���V�֨���"�1XX�c�0)qnEWz7X�A�XY�tuZY,����46�\�m[�C-k��H�ۄU�v`6���M��sE`Z�_UR����b�W���TV�W��J/�c7B���w<��*.��s.��IZC�K][reDDh�OPt�Ѻ��EF�2�J�E���<7݊���m�	QˑA�Y3I�_f)4��DƄ��vР���G��F��JD�T��B��0Z�I�i�6�
�2͈����b���żj�%��]�����1Y�H-�/Mh�E�mkE�z��3Q���U�m�0X�#�g(�/e���oj��J��wz.�����B͙t:�э臎J��r��w`�|y*<f�!R��Wٖ�ki�x��ɟa��P�F��v[y/���h �oq�8�$��֜Gn��=s�E���]�X�f���7��c{��UE��(����qgTTr���Ečv�C��xq
#GZ�+���S��ȱ;ћշoqt���0��p��[<³���t/2�X�݌<��������1U�����ɐ敋,*w��X��[�nLv�tS^�|)thuW������J�t��Y��q�M�(-T�Z�O%���ic��6�9���u�a�U���믲���8�̂Q�h����tT����^w;(��]{tĪ�6*�>��0i�%ۋsFL��+^���-u+�BjɼV¨:��dqEw<�[�6�v�~���&t����w۠�@�T!tR���x%���Y��_R�Xf����2����`_fJS��C���a�s�C�X���X���v��#dѿ���c1��|�Wj�k����
�U��jK���bg�<G��vXR���w�l��ѩŰT�9�)��KU���F�PXe-�b�n�t�1�P-�*+ ��Wn��b�#x���N�X�x���\mt�ƙ���B�TDa��ֆs�#��]��u�V,sv#C�4�0�5搰Ţ`[��w�ŕ����>�r�m�F�X뽅�q�'6R��ن��N�^mࣗX�"f:��"�Ե�"A���EU�T�L�2��1��x��X!�W��UM0�"������?+�	�0�c���U��ffkL��]�i0[h@
�Wp*D�,e����^L	�f�Ӛ��(	�ˠ`����)l١��ҋf�h1Q9���F�j
�f���{g)��ݫ;�5�#���Im-�n*����AM��[�u"�ݳ�!<�!�3�m��}����@� ��dȻA[����DT�M��M��n�8w!TGY:���(ݸ��_]X���������6���WKt���3���ר)�|���v���[���Ү:~��7��o;n�¡Q@�ܓ��hu1R��!cp9Wv�-�z� "NLX�6�튺��Ej�>�;���0l�3$Ɖ�b����B3��C칬� y��J��+��a�f{+�O��*��q����5��F�����
QA�k��4Nc5�j��٤��a�sl�KC�榹�O��c��ݎj�����W8�3�S1�j��I��1�G#O��(>~��Ug���PNB~z~���}6g@ZC�;�{su]��k���к�:��zŹ�mFF�Q���/����t���oe�S�������WÆ=f����c���u��x����i�g�(\���{�I�/{g�ںE}��_l�W\�s9Rb��b�^��v�`r�S0YƇU�GC�_w���D}[N���:���KX����Jq	n[z]����!]u/�D�=�0n����u].�]�}Ԯ�}�3k�ׁfE�w���\*a�ȴ��k7Sj�����G)�nd/���6�����Y!�L�]ChmuN"|��ܷ�*M�U8��d|�:�����.��披"	E���[�Lnm�Lq���/CZ�f�ڣ���W��ϲ�s]�=�����g���Qd���KH2X?Q�����k��s���¯UD�P�"�f�b2�Na`*ӯ�s/����貋R���{�E�wwxJ.�iv⬄E�2Z�CEȅ���D�H�]�;ܛ���X�,���k3.�b]I�r
	!�-	IQƃ7,�1St�<wtMj	��m������%�i��j�\�
;'.��W�c�����3掫�9�C�E������}%�Ɇ��Ǧd���7*T��䑚��Ӗ�-/u����em�V��`�\kr����r^gJ�*3V��h��e�ZY��@!���c�ʧ��+*�E5�iG�[�pv�9 �mZs����Y�0�c	������l���L�>vy/5nPUq\x]�w=S4;���"�M�s5GK���jp۩r�������T̼Ŗ���)\�8��G��(����i5k��V4ꫴbʹ%���]T*}>5Mi*���!yP�9���Q�ee)7Ϙߎ���0�4qܗ��9g3�%8z�!3�*wT	���6�K�;jM���E!d:?8J�TA�7%�y�Vbא��U5���T#����Y��i:Ov���[M0�e�v5��Nu)m״wN�ؒ�V�F���-��᥄ ��$Aʹ��Ue�7��X]F�r�$	.G@��)\~�p boN�kHhLQ��ؤ9Mo�`���[�)�,:#Ɋ2ۘ�Z L²�xf*,6q֫2�N��MG��Zh4�A���R���Q��d�����)h�ARJ�԰e� �+>/�}-�[�u$`����N��M!�T�\x6XTCi�kW]��z�ki�c�r�wvܨ�YV�[e�Ӎ�H9v�\��JR
Ӎ,��̽�p�K�	A�Q�i��te3E�	��(�(����0�̓	t��qKA���0��%�ae�bIct����^ď@EiV����ҐUJ�QV�UEAj�"j�"UE�KcD�m*�l%%H�v��bՖ]T�n拻���+J�	DH�Ɖ"�e"R����[t�.�%��Lm���q���2n�+d՗[ː7"ܨ�c2����	#J"f�[ic-$\�K��q�3rf�IE��1��H[J
Ҥ����Ż�"ʆQa,3y��YRiW�,%����|�&'��᾿O��{S.]��3.��Ȳ��SII�B��\�-��6�#z���jV�6N7%�dH�Î%�R��х�L"�Ȥj٬˂�y�|Ջ)�n�'�X�wf`��l���.fȋ�k2ћ!k�&�]��.�A2��D#Dx�D- �m#�.^��u�_33��j��vf����La.黰��!*2oY�$inAB�m������[Z�1��I��b��-���}�����(Kn�U܌�8ˤI��T��C���m9(�#��\"��)bMYe�D�`�XB,�)ԫ�r�b�T����EZchi�c��<�CY���mQףz�v5���O��i[o.�Y�l����S$u��L�X�M9�
�����P�:ۉ���)f\1�j���֯5��w���)#sXL3Z-����Щ�.�F�Ad�- �M��ˊ)t�C	wәvccj(��2X +Cщ�V�$�K5�懈z#b����S@��P�̽j�YXEd���Ŭ�d/PS�"�L����Zn���K�&�&:��BEU��]�->Y�����B�����#���X&i��/S)��&d���&�5�tEj�Q�;�%���7�}�U���n��m��rM����P��y+f��):T��;��8k�n� ��g�&��C`pH7��j j}.�WSG�J���<U[嘷u9�[����fe�A�V*��d*�#7��[�b�\t�uL�f5$�DL�E����W[ӷ2q���֛MM��!�Ӫɐ����j+oͻ z1��5
��C&UL�d��ɶ�Q��(&�@!g�#���Y��`��B�Cu�j�Qң_�f���A��_� ����g2��.[�Q�`ڻ��yx�R6�t�b�rak&���c/h`y��QMp�s[�m��7��/XE2`���NR��jeE�'�O��X��a��#P�nY�x�eMH�� ���S��32�����Q���)@h�P�ܔ�!F�3In�U�X��E*�E)�j�j���M��jIN�TF��P)9�j�j�SP��B�1�d���DR��҈��T-(��2��:�f���Jrk��[Wk-.U���7y�W�l&���n�&��i��6��[̻9�:s7}���m���%�f�!;w(U���/�F���	�U2	%"�d�xh�-�2kMj��B��K.S��wM*ҲTQ��%JP-���(�儖ekU��֩�[DDT�"(*�(Ԉ�A��AQ#I%2̶�9sFɗ�,8Z��C���f���D܄�[���Kl[�HC�v T`I|��M�x�@�紑�ڭ[[�~�&�4cB:,�Q�b��i}p�D2ٻTWћY6]R.�J��EJT��K����@6���h�e8��.óUO(:���*
۴jL�f��{%[���"E4�Ջ��:�yt�#�ճ��aT^B54�g%KMv]������`yt�<?m���,UAK4�:�r���|l�I0�n�W��#[��cm[�fɱZc���6��ѻ}�ζ���c�`��.�T+ea�����}�;f �0���ב=�Unv�F��}SE��>{��I��|�W�V҅9�Cwϳ����5���S�lq\;�3N�֦��d#Z��K-,�*'��8��r
�{�KLm��
l���j1J�q��. ����I�k� ��ɼ����>����)T"�z����0�ؾ(�8'X��.��4�2�f�Y�q�C[YI�m+��pn��N��*tD;YzE\�8�k��d���CuOU_mL�t��N0��J��V��eҋ����g+�cS$�-0E/�����joId�|%�قZdi��Pݵ��v������B�ۭ�!���0KUN��Z��u�hc�¾\_E}u;y�]hI�����ڋC�	�P򽙲=��k�S|���~����j�_R��:�f���J����_ի5^�XZ�~#�q�(&F��wW2�#*I�ѹ�ÚT�Q2�yZ|�fg�8Y@�e�KiQ�7#�m���ߴ��k�m�Z&�7_/��s!Ԡ)c���T�*0f��ٱ@3I��8�oCpf\$n�+�y�����PJ��	)k����v�5�f�[��AM��m$�๛�v%�7#��-����B`�t�/#f%�UP��Pd�Zִ��Zִ���I%ne�u*���t�sdr�P��|ˠ�h�̷�F�U[FЋ��]�6V6P"	!h�ZPh-��R�m�D��U,]UUUUJ�J�UUUT�UU*�Ի;5Q����x�iV����K����UXElڪ��E�5f���  �#*ֆp�ҭ\�U��PZ2�L�(�۩���N.�AL�`���欒h ��6���ꄒ2tR�ܪ��c�Ȣ�S�s�A�N�WK�T�qo:K���ڕ�=�8xg9�R}yT��#YL�(�#*�+JJ�Q�`+��0J�,�����)�"�UUUUUUU\�-UT��)��*Ԫ�UR��UR��l��jL��d���PE(WP;,�"�l�G�q4%�a��p*՝�O�Ɏ�հ�m%S���]kuɮe�ppn�Si�)J*54��Nĵ���KH1);�գ��	����5R�UUU##qg��M�j�G{ b��M�����x��Ҵ�^��������R�6�Q�0�*���|>|s�
��Rv�8��W�!g���gV�W��FU�Y!��Xlʌ��rP�t�����S`&�UuUUJ���E�*��������Xr�*��9j���U�mUTQUU*ҭUU6�����D����UUUU�j����ꪩ��b��SU�uUUUUU�j���q-UUUUUUU<�UWUUUUTQUV�c�
yY��R�%�Ҹ�<p�u5	��p ��ʭU�U#���k(�Ԅ�*Ҁ���x�z�ƪ��U��vg�V�e�l��VS$p<�7>�! �}���j��ޮۺHJ�������\(�!d���7���f����SoG&diʍ\[r��$��d�l��	�r�l���.��VM��8��b���!�{�,7<9��n�jw�����u��s�7�����YΚ��{F��m�C>�-ŪAȣ�������n�Tb��̛����q�X�{�q=8֍n#<�)��ƺ��7V�q���ܓ�̔��z`��*ub��v����嬔i�v�¹ss�0ŸnE�3ڡ�{p�툵{�&۪����ю7�w#������T���=�nXȅ����0;k��e�Һ�������x{A�6&���nvD��=u��t��ۄݳ�3��d�Wp-8�m{!&{t��v��5V������[y�s�z�-��,�����8��d4��g�<v%�xuw�Ͷ<vRI^\�n�q=V�8ݚ��=�8[Fw=����V��v,pl�5[���1���:��<�-����4v�j��I�ދZݳ���=c9�C��$�ZD�)cR]���#Q�˥�$��:B{#����2��U\��Z�)�.6J�-.�*jͷm��E���Eٴܘ��;lcr拄�M-�r�R��h�Tp-��Ղ�m��=V%�*fN#�Dh�t�jNyv�z�!L �ܣ`��?��|���Ml��I"7;Ki[U0M�9؇m�iY몬v�3²�m@����u@[R�W0�v�n�c�1��*�Z(��,V�����Č�A������$�����vmZ
�;n(�Cc: 2�5U�_u2*�e��RP�N�
����P��7hV�R�=��-��hѥ�.��:'���m�Яz���s�T"A�3���'9��p�	�gl�s��탬�J6���n�P�,nyM����/��n.S%ё�ɻ;�=l&��lvؒ�ݶxE�n���^x�욭�9ۄ�]�W�v-�7WWo9�������	68�F�&�[*I�[l~�#�iʂ+@w�|��m����wx�[w+1d�B܉u,�S/�<��{K;z�����u��x�8��⻱�d��Su��N��5�i��:F��fx�Ů۸4.�!�;�\�Ǯ:��h�7���i�w�V����tc�Sd��x۶���Xwu=�F�=r�;��5�;�:�T,�qcv����;�rN�r�>�6�l�xw rXl0��f��WWgcC�#8�tq��W�Ѹ.{Pn�>s��C��M^�ѩ7[M�=���\np���=����l����J�M�pT��
D�7ͮE�{�%J�P�;Y-9��a��t����g6�rk=��s��T�r��s���qDc5L�[
�΢�´�4�\�E��|Lt��pn�m�2O�]&ژ�g���f���U��4��ѳ#�m��ÈV7ILvn-�m���Jd�W\�L�.�M��g*�im�W��i`P�����C���v�������rn���:�q�Ĝ��V�O90[' +�/@����ދ�r����v�Ps�Ů�Nvooi6��NMNm	3MN�XD�6�-&�N�y*F��Rm�J��l+9b��Ŭ��`h��l8ìu�Z�	����+pZ�Tl8�b�n�=�'��nۆ�Nsfʘ�K�GNQ�mq���sѸ͜�͗�S��u�bd~V;X�v�A�k��vܣ� �k�n\�i���N��G;p�OI=f�s���պF���d/]��� j�ͻewmUr�7:��є|�T�c�	�:9kIμt{{jnɖM�R��0�V�q,��LB�E�N����=M�vG��9�۲�����ۨ��ڠ����ĀpRQӻF��mn��د'M��gK�������(��#��g:�wNf�T6���������G0���:Pz��Qďb���c�����Q��ۛ����ݼN��:n1�r�nx��m�秶�i���bLA�r�,n[��ǻG`�z�@��u3���k�ی��5[�8^gE�grM�]kv�#^�h۰<yy�׌�sС���Q��Z�ݵ���GF���hx�n���m�t�ͺ�yG�X 7��N�َ�lb�ט��w=oa�s�"�z.����!-ݳ�� �;��^�m�ka�1����v��[�y;�==c;/)�p#�9܈z��ê��2�;�@�]���� ���p67<�9�Ń�-c��<On۶z�ݻ�w`�拝O;nzC&^�a-�[e��ceݷ<r�n�Zָ�y.0X���@��6�uBȏ��+��ܝ�Kw��ǃ����Gd�������oi�v�&v��n�ɳcW7Ok���gع��V��^��k5�9wv��5՗�x��ݸ��.W<|^N�'n��S�w\��O=q�N;Al'�\���C3*]��p�����2�s#1ny�%�1�@�o9�)�s.�m����Z�nu�J�;a0)mm8'9�Jm���9�r����.�����uL�!E۳�in����ܛ�ã&���1�6����<���/Euʇ�ٰ<O9�� 8�/Zyk�!Α���b�	�V�6Ϙ��R��u�{W�������v�Xm��Y3F(���i���"GC��w80�sl֫�YI�-և�ΰ��Q�lY�\����V�SP�#�����ͯ;lۣpx���l��H\'dEKXۛ�����6_W-lv��ͬ3v9[�a���3�˼��u���#�Ի��̸�-�Q����K�crl�qa�U�(�$���.d�/̥=��u<��9<[l�s��v�l7��X�N���]�l�}����q�{r�7c����p�s�ӛ�v� y]��=�i��⭻WG��8�`d�"�3��Ah�����Z4;�+�����c���9�'m��/����kp5���u�s�^:����1���r���7>t�\�/v�r�1;���s�n��-[����W ѣ���Gv2�	�q2&-��\2�q�t��؍��]�v�;i���SSY�<<�m�;���z;8S�)�[���p9��7g>=��DW'�:�V;s��2�ݻp�)����oew8v�[h�ҦR���^[z��r\��]�]h���殱Ê:���7n�(!�������v��l �`�5�{)�Wh�l&�v�[��ok��c#dY���0�$��˫Nw��;e9�"Z�ԞT�*q�N���;*��v��T[���kv�v��d�x�l���m�tgV�uplq���9����}n:��%S�"<�w:����z֫�(�<'�v�ɈF�<��gc��#mr��s1���zhSV�S���(��ݲ\�XS�!�B��v��63&(�8Kƫ��v(�1��/7���`D[*d�~'�()�c�q�i��s�'l%d�s����j
�<����n�z���^q	�w��G�Y���J�����������{f:��Z���=����Ɲ�r�잊�-�M�'��1[f�qֶ�\h�s����G���g���iD!1n���vu)E�8ݖWMv�ۣ�2v��]��]�:0oLk����i�z�N��q�q�o�ۮǇ����,;�,��WW[��Ϟwm����Sق�ݶ�;V]��vmLv�3������m�I�mݸ�$��ܻ�ku�!�s����[��s�x����$�,l.�������8���4�h#�=�)����=�#�1p�Ļp���D|>k|>t=x8�y;F�{G@t	=�!�n6:#u�vܮ��#q�m���Id�e�3��E�u�2��?>�����mN�pNn^�pe�"Ѻ@��P=�kh5R�uq��<m��lg��WMS�1
t�ݵ.ln���I�K�h�F�KT�]chu�9�O{�gW���ŵ�q��Otz���m�{<�x��f�����<۰s��(e�n8..�v�\c�8�=R�&a����;~x�Nڌ���y��nq��Gl.�[�*���X#t<�Y7[Hq����c�5$���g�L�qO�949t �Vۡ�Wr��./@�h,��8$��ڞ۵�+���<f�d�n��t��	N1��y$�!zF�X�H;t=v�/<�tn쎨1����ގ�qGn�j���y��#��W�ҷ�r�Rs�4m���7Fx8������|���6�`1���pl�z�on�p�٘�	Ψ-�a�� ���T7�6���ڑ6��L�ꋧm0�<�u��lѨ����sJ����@��^w�'8֧�ەm
Z��
Ύ����l��=�K��wVP��;�y�-��"ܴ�j��0�X�m�Ꝺ`�`�틢���Y��Wom�'�pu�;�4%��տ?�������h�(� �B���UAAZh���E �K(�AUC^��ϥ[�d�<ʉ�M۝�h��K�pV�35�R�!e�!�G����]�B���INj���d�C��n�Zyk�޸�tLC��hV�U���TQj���.�j����]��m]J�mVS44��h��[�H�#xC��[s�F���C����k�ia�m�G�mhC(i��(Y2�u�d��eT�evM9m$�T3����ۏ]��R%�ٝW��G�a�&iˡ���gu�nUl�s��̂��\��ֹ��!ѧ�)��z�(���2�ݭ����uI�`���#uL�V$�e�"(K�\��v��յ�X-�M�9����;��SIf�t^��ɰ1��17$f�K!�`L��5�s��66��j�L�ݜ�.�71�u����-���=3�a�m� ����WN��q�Ⱥ�K[���,��%��t[r�h��<�+�Du��(�������/-�;b쁄�Cl�+i;n!��n�-�����|�{ޠ�բ�)h��j�*�h�B���Z��Z��P� P
�(�*�Z�
��P��Z����
?�o�!�����Q��W &�j�F���\NvTW��#�l����9p��L�9�q��ָ��3�,ݰ�4��lej�C�[��c�<�3���J����{���˻e�+��v�/e{���R����?����Yy�0٫�Uj�K��K�Tf�Q�W�$��¡���AMCmc��o�����q�Pi���*p��^r�b'bI4	9�,�to��˕.�Eã�{Pg4��� ��Y^�[��&�mG5��c�UM�"4�TJ=F�vС�]��*7�6+8j�[�3nN��^��#Y�b�t�В�/�}��vIbD�׽������)e�;=Y[���WӥU�y|��f�H���na�9�t����2��'���Iӹ����c��JF�
7F����r4�FZ��B;�ԛ䀣.��M����T3
T��.M5k���]�|�p��fGZ�����K!7s���^j��X`����s�1@G��z>>C���E�P�rlӧ7L		�6��G�TPI�z"�Q�3���k�fN��I0R��$Cl�]�/q$�����}8���F�\�q��R��Qzs�Qs$�Z�3=-n�9��`쐔`��`pNt�]��om�Fw@���ӳ�D§�ٮ=]�x��FN��$��QL[(+T�T�͚��hо��(7�~��<[="��(�q�.��Pԃ/6������P(ٷ;�y9����C�d#0��b��>�E:;�wL;�]j�^�!8wpl��v_�����εζ�vk��V�ۆ-�S���9�]�7�x��m�:��<�eݚ׉N����Ign��H��x����۳��"�IG�Wֆ����r�j�M��{{�;I�:W6B�5±�-�.�3���fܘ[&��H���~�5�=�i�Q�29��ȝ�HI���&�F����Y
q
���>{��ƽ��\֓���7�E��g��o&9���lW����f[8d.��yM�2f2U��2�\�8�U��S^�dzS�����kG}�c�-�^����1�i���w�a� �����P�N�������WsG��8���`WTV�mCΐ!���k���I ŢG�aR����l� '��'#��fG7���c���:j佲���{�6b�/�j�S��_�bk�{�5����\�
�b�1`�cX2��r�.��I�����!*�.�5pbvPz9��E�Rd�|�S��|���*�'/�����]�=
�q����"5@�$
�_In�#��Q˕s�F�a��ֲ��!�^��F#-�ұP	.��L�$ d�ͮK.�-��~# �yyB�d��Dv)LV�I��\ƪ� j�K��)�LԠ>�﮷���:c�L��$[�|Г"Y��r4�6L0������B)����
ssD�vh0юj��D���1�ܾ�S޹���*�x�MH�\�4ɫ�}����d���&�2C������]��Gu��"oUo�~�+�f�;�I�3c銩Ъ5��3�1xg�MCa莤��_(/뭁�AUb��5i�B�)�w��j���l�K}�.Wu41Nt�jL��s^������SQa��D���hQ��hNeNU=|�� ��.�'V31�}?I�_^qy���]�ImYnVd��bv��Y�n�xo�}�m�k�n;�Jsm&)�lH�P�f��lU�+��>�l�t�o��)�F�i8BY)�H��6)���h�тh\e�yP�.2�m��YX��ʸ�_�Ѥ��d�2�"��-��Ŧ�u��e �Z���㷬(��MJ�$���]�0�$Gq�n6y� ���a|%��޳ܵ��/2V��n�o�N�Z}�]mri����dy�D���w	]��:����I�45�uRIb�6�*�$Hy��m�,*Lט�;�N�r�M1n��t4w���d�x�]��s�����k�m`o��]�qt��ac�"���{��=6��r�S�-�譜����\�r�!:�=q�썾*z��kE�_�l% ��K�B�/@ ��i|T-V�A�H�W���3���6�{��K���Qֶ%��^��1V��s͡�z�M���`�����̳��;���gp�m���՗��Hj�D��Y����h��$��&[�η��;��e�kn���ɲ�"C���]>�<��5TN�;���-��84�9�xk����0�rA���w�(Z��p��\ʨU�r�|����C����qD�%�m��/J��s=�RT|�K��9�ϰ�i���o2�ម]���꽹�=~���uA��rb [u�s��Q�=W!"�j��|�:�Gv�
��\3��A�>QMs��Eni�-����ufL�/K�芏�F!1U	_�"�KY����~�}�y�,����.$����}d[��"�ɞ�S	J�v�e���ep�b�e,���Һ�-d��5�6���M����0(�3
F���ǔ�	!��{oS8jl9	-P�����*��Wլ(�*D�R��!�i%�`�v�X�%�r��+��ok;��)jڍ[!]OT��U[T	=��Rq�;mA��ʚ��^�}��@5��<��v�=�9�tuE�ܸ�-.4���鉎�'Ǳ��.�#awc;E+��[�ju�k�����$z2��|�o�7]=[����� i�&��!9� �%#���)]XL'�����е�0b��B��|��Ҋ;�=���>�ȡ��
fc�M�P6Q�0��# A��\L���I2ҫ�4/o/���ϧ��'{~�hc(�]�O3"t�{	�[g��f������tVѰ���
A�u\�c�E�9�0�B6�3'_S�C�j|�#Z���70��m	ŮX�iE-
�B�y\n� a�N�P"�/�ۉ��]ܸ���ǟ�¾8��^e��0�/9����K��!s=�N��Q���9��t넉v�HI���IF��Q���­]�G�\�o;���絾b;a�]�˼���l �g*%+��쁴G{n��f��o��XF���w�� ]*z�Q;*� �[��OP"�ځ;v��֤y&v9m1%�[�r���a$�0�(��	d�OM)��9��3��r�+(C!}\	4]L>S0 s\���2a�"FF�ЭF	l�� ����h�S�_ŕ�R��k���02�F_椇��P1v�eVK����Wέ�UG��&.��]��@:v���,�g���nB�,[>̦��;n7X`]��c���u���<(�w]���=�Y��xp�����zVZs&އ��K��h�0r5�reC惆�xE�0��W��9�#��zѽ�ڈ^��fj��]{{x
��f��G2I��7c�=E� m5���!#P였��48�jap�x���X'O;��e���!@��ȹ͞=ᥚv�I>�<�|�$U��?I����oo
 �R�J��H�1F���I�\/29%��{3���rl�b_NE��o:N��{�9
,�o:^��Dz �C �%̬cO�`c5Rf<�������y�^�XF<�Y���y�'�����N���$0��F���"+���- �^�[�|��-^sXzhje
;"���ŝ�Y�ڱ�&�Yy�O������E�|̌��=>���%�k���U�E� � N��JGKR ���h���gǻ�D�����.\�C�\�q j���@�PV�]�*o1��p:��2��58�5�)�.�P�=HCpj��ߌ<��T�j�`�������G��Y)��=���6m�ir� $EƑP�7��V��p��u<��YBA�ѧ*�e��G��}������v���Z#�}x�D+��h���������'�p�@M�
ۖ�e�i�R�e��}��D����ٮ��Ǳ�.{e���y�ds�O|�����&�|��^� �}�h�nTɪ��P@�K��x�8��	cD ��A�
.����4Q6�+�!5ynFw_
"��D0�t�P�=�Ǒ����_\l7�5�߬a�:���n���M��7���z��+D�q�x���\b�Yۮ)Jz7y�'ݨ:�6�}�᱒l{��z�L�<�v�5�W%}�N5-j��lH�T�l�g�a�S��?chͫů�P0�Q)�r#���t��SfU8�'�G��O[Q��{����y��al��^�:a&;�p���Ҩ[��-�ۛ�<�Ѥ�h�;k>�Y�j���,�9P~��ޘAi���8"�ù�d����8dkj5�4�[�d�����W����tmo@ga^�23*vSkϑ��x6c�q��O�L (���GD�7�
q!�+�G4��:+g�ER�g��"����n��lw#�U�ҭ�T��ࣤ�v1��,܎�L����r�Qiղ"�|C�X��Q)@�� �f��:�h����ގ�:�R�8��I�A���O�WՊoPq��Ck�mHu����f�Ul\�8⺊�@ ��3���p-�$2�8&Ff��5=#��Wd[#�+5���;��6��Y�t�s�hd0b(p�`�����6�q�B>�_2�;t�h̙W.r[u���NwMB�߼�w�%sI�%5�c�#H� �7��}8�f9dK�7b�dB%�EQJ�r�*��D�Ϊ��p���V�O6�![#!�����l`�q:V�O3GU$�R���;V���ͼ+�i�)%E��p�b�-�L�@��o�,��%�L�7���|�ˍ�-髮!��%Lm��(�2����S9dgQ�k �~��Q��y�<|(��
�E:a��Q=�Gy���8�V|j�:/�ň} �ĺ7� �C��"6�;ڵz��{aJ���<DDU�7��}@f�qL�!]��+����N���U�Y@lS���c]j�$��%L�J�!ӵ�R�¢ޥP*{8��qJ&�[�:���2��t���ݝ�mv�/���`��uV�ٜ�p��մ�t�9v�&����3�m�+ӵ:6�ܸ�L����r���L�/���?h�}���m�p��<dlĊ�Afħ�������v߈ml��b�eJCw��Y��<<�*��,C��0^�Zh+fQ�0i�jPC0�u���s� �o_C�]
$�E�2`�|�$���J�o9P��	�y�r�ǋpH�F����������Syk,³o�gϨ�7�T,B8� �WY��<��Z~�Z�f��4yKX50�wۧ	�ώӯ������S��,�RAme�u��6�۵�ˎ�|����h t�N*���J�jҫ:�*V���܃��cj�z��.��
����S�8[}{ځM��t1.�6F*�a�XL���ˡ���S}N����S�ޛ�+�F%�Ɉ��\3�t�U���"p$����#�M�[�7�s�7htewTK�g)8`�y刮�q����.�w\r�2𿱯�������
��y7��F\N<9��̛��q�Gu>���vg$�-ā{���ҷ�JE5G�JӸv&��ٙmC�@/�Hzj���BD��.��vj��{�{y�V7g� abR"r�\�	?J@�V�UPNG�M�e�kw.ݏB�&e��\H\g=2q{�]�Kp�7�ŝr&��a�N�k\d�t���HL�Z��0j��2�Ib���X���n��Pg{�2�h����'9�h�DQ��W9I�b��VԶ�lm ư�F2����PP�j�;Z:(j�*�5��
��*ph��E������#05����V�3re�-�c#ԛ�����{ϯГp��/S��{�����0UQm��y7��b���ܱ��L���W+1�9y�Yr�\X<MC��~��O'����5���~�m�]�D��73Uz�7E���'c!���&�A"����ɖ���:��v�{����#rU�������m%m;�s׆o2�MƠ�(h��n�a6�Q��A�L�9�W��ܜs�������27 �-±�mD��J����әAjq�L������Rt��.O�ș�(���(9�ͦ.b��2�|��A6��{� v��������A��!�,�F+<D���;Rd7��X�7�~d+Ԇ����@Ki�x+��A�����!�&oN����{l��
I[�(Ud���P2=뢾�0T�C�|yk��(|>"�[{˾�]S^j�g/��XU��e���s�m�K�\{ގoN�C��VX���!\0�݂�m�;�u;e�F�S��۱^>���E�Y-��ɪ�9*�ǯ	��v1���C;fk��]@�cz�;����v��ō���.2�z��LŮ]7V �/��';g�����˗Cl௧1!����]���n��F�e��'�|�p�z؋7��._{ݽԌvY�O{ʴ���:&,�ۘ��k2�A�[����Y<x ���s	O0�I�j'��l�[�o�d�,��A��	љ�(�8��ܻ�x�x��Ъ�5h�rwjε�;�qu�9xF��DULc�=t�����2����W�\P�w6�]��-_O�|(��W�-���M	J
4 ��P%R�TUU)AUTw��?l�c~�oOG��Q�Y/���=�#O�U��'�֡r`fV;n�6ɍ��Y��J���x�˥��U+䘵��2�������/2�F���##��.��m���U�@H#�=p��4�M���j��E��������8m㧝^۔ݴ!���pܼ�.�6�e����	�Y:1<�nnK����ܡ{M�.Na� ����k����f5��[l�=7n�i^�=srk��s<�6�y�n�@ޱ��xz�<�����j�{ O�5ۂ�O�Gk��や競<n��{D�9����ƭñ��g$Ѹ�z�y�wU�:1�ֻ<���x���Ƙ�
�݁�UW��^�on�]���v��\&Y^��hMƺP���s�7��6�����O�ۭs��˸%�)X8�i�Y,�*Ķ��%el%Yݸ亶#9�]�XۧӮ�H�Xv�<c�μ��ܜ[�Z��]<�3.7qɎ�/^}w`�Vը63��v�kf؞!���Z�7 0 �FW��t����d\\q����'U�8��د
>ݺ���3o+���Q�:'qؼQ`�x^ݮ7Z�Q��&�ۙ�{c�q�p{<�����6��<�%�t\;���F��\]�<���e�rh%�P���O2첿8�C�Zd����TC.U%"_�xџe�}��Y��u��J;!B�V�%�|�ί�Dy�c�ݥ��̽�u+�ܕB�i���}0��2�n{I�5����9˓v������Ӵ7��+my����b~B6Ѵ��Q$+�ܕm}�k*���B�'�@�TJ���&�?_�m�;�Q��7!j�Qr뺫�Q���s`)�9em4��џ�����O+U�?�]Lj�v��kZ���p�!5Ti%k2���.-W��Ks.��j%�J����K�U�y�\Ə4F��)�cAm�i��i�k/l�7���ۣ�ژ)��^@��Ƹ�KbF�ih�DC�~���g/�o�8L��*$V�4lh�R�����.�1����y���葥�0e�m��p���l��e���d��F�j�~�҅����E1����:n�3!V��s#p���hu����D���ٙ��)��T�:�D#T�({�W��X{ڃ�;JSͥ
Q$�\��rV'YvXs>����Ld�m�c_%�J��d�A7��Hj�j�/�n����Z!r�Bӏ��)h��%�Y���fU֙+�~���GemǭJ���H�YY��Q��r��W�ʴ�����)Eɤ->�X�3�º�����F�v
Hƈ�� ����F��Y���	J���v�w�d���J�(n欮�{\��-*5��}r���j���DhĊ��YS32�Ԫ�i%F�"kMZ�{�c��5wU�L�1��V؇��7���|�Co�8�h�Djڨ�j�V����Yp6�DOk뭸����Z���/�.f���m��}�ƾj�6�D�z}eaﷸ�9���)�Z�Ͼ֨�����{)�����Ad�F�RAY
�E��˖I�a� �{���{�/5�ǩ.Wȥ��B���-(�A��j���;zq9Ƹ��(�mV��Tj%F��K_���bѴ�mۦ�>h���Q+cDJh>�%|�Ď������eC��A�J����ģ��Ҋ�?��{�]F��S��i����~�߈��l�5B��W
Z�h?$�Q~k7+Mq�Y��7��yf괇�E�ĩ�F�|�M� j�Tk����1���j��@��[��LJ�D��y>��k!�	z�C�)A@�4�,���j��j�������$t�n�'eW�y��xg���
��5\T-3z��y��<�����lm˻Q�,1u;d�v˙��n�e���~J��J#��J���Q�׿e���C��V֕��i<!�5SЍi/]��f����-�iڴ+#\LJ��|�Х��E���m��]��I㿹�A��ƺ��5%�/�Uh��z塉��|k�6ݷ?V���$y*�իG=J�Dkzﰯf���xC%�дy+� �Q*�"P�P�Gߵf���ˣ�(cZV��9���ᮥ����T}!^�^~��9wUhuވV5B��/Ҩ�r�T����+9�_�GH-
-Q��j��vm{��R�Ů�����s3A��'%���?~�w*�+���1�;��c{�6�\@�GX�@��At��W�����@�Y�*��M7v~�\�(O�a�Hp�P��|�~�ܯ8�������VMY�3��U�p��j��ZV����S�,R���Z6�3�Gg���L2�emb�~Od��ƋhP�U�ʭ��V ����3���:�5B�A��>zZ�~6>����!~+���2��[V3-,��}�j�+߿^���4�6�����Α|��u��r�4bk�d�~�׮����ƌkj�D�#F!cFo�����j�v@ƣTI*�{>�����~Mw�[~Ku���?y��\�W�Z"|�D�U��J"+������ɲf���^�!m�f�QҦ�-+cDk�}�Z5�7y�5D�:�T-��"�-zx��>�<��Y^���5둭!�cWX�ך4یC橐��A�q�ڡj�IT>�D<�+]m��<i���B^���X2�m%�bW�K�Ѥ��1+�B�gn>��@���K��� Xj��.�T�̸��UJ�N.��aJ�α}S�l۾����AJ�.z�]l��EqJpX^*v��MB\h���g�H,6.��@��EmA=5�z�s[�ν��n�<r8*���lj���9�%]��[b�0�:w=�]�!Ye�e�\%ݪe�.�fg�j�p�m���U�xh�
����c^]?o)@ƨR��Q�DkI�5��U���˪�N���Qh�WnU
Q���8�}��Hoܜ�U[j�ig`w���[kJ�r�j~��Ѭ���m��`��=��34��TNn��5hi#B�t�hG~항ߵ��-��\�R���_��+�D@䋌J��R�W~��s�k
۴<ߠ{6sٹ��P��J�5�J�7zJ��m�kH)�EE�9%P��F��kW�X���U�T�E�th�Q�j�E߬���G�wvvfK�����TI(�x����{���
���V�u�������2�I_|�Q�*)ւ�TKJ�%�_ji+��:�WZ"��W���TEK�P�X���^]OsyF����K�T(MM�C4k�5Q59��2~��5�[J��(�䶿4EE4�j�%cJO߮��~��ޫ��f��W�Gi[B�8���U�\V����Ĭ���7r�K�������~�F�PD����w��93�:�
�-<
�6�ř�̱�[j��޲�v-L䯝rU���V�p��h
���}
�\ϵAMP�\B5�u��u�w�Y��9-��$M!���q�[V�C�k��7ˮe�ߗ�g'C�
������ե1����hƢܣ�+b�Z'n���zh���͋B��%-D����M4p�~���nkSSTWmqR�m+b[Vմ�c�H����
����Ӊ�7�o�6�����h�|�ٗTF�Qxѽ�����QJ5%DZ#]j�D�"{��bq�q�G�I��h�B��U��m.�j�E�,��/?r�<8�S%��c ���睚#���V��������y#X����T��)����/9�uXѡ�%�UEE"iN�X�Dh��Kh�E�KK��d��V�Z�!i����<�[օ*��拚����5��hh�Dk�~��?X~�7��戛�d���j�E��-7���n��wFh_d�uQ��(~�i-"�}�^�A��r��+�EE�~��_��s�~H�Դ��$.Ө�壣LT�sk6!�g;���7�D.F�[� (~�G&�Wl��=f��˺�oY�-/&+o1�o*r�q�Č���x)���2ڹ���q���7��PCg�:�8`�H��2�W>���̘A<�qm��eԹ,�`�r��/�Zj�P�i��u���58�!DOʕ�����E�hEq�K���M�4C6B҅(ԅ\C�k���J��&7�W�����cr�G�k�i[�.oC�TR�!�KDh�=7x�x�kwy#3Tm�M�D�ҋ�U֬O+U84A.~�#��0Z6���+�}uX�B����s�o
��ZtQ�y�4lh�Þo��[G"�=p�{�X��٬�лB%D�j쮡?J�4����_���+��~߬��/_�jڴRIQ�B�lK��$k�啓��D4i�Љ_}*�Ҵ|����[���l�v�Y��V^Ef��l�p�$�v�<�R��{�75�ю��4�[�1%i��nQ�k﮶�s.δi��-TZ8�˄h#F��l��W"��J�o%Q�j�Z7ߵ7?r�4[]��ް�j�<�������V��T)i�'%cT)?Jh�v���5{K/1��Q���Z�mL�i���E�9%��vi�.J���ZЁ;(�U���V|���g8\ҡ�
��b��E���w*���Z���jW�YL�#]kO�&v�#VժvJ-+����Qk�ϡ[ә�Ts�|��^E�H������U��E��xFa�>��z4h��4#D-��8aU�p�yͽ��ny���p�_8���-��EE�;%P�F�O׉$��\M!��h&�ƫi�iZ���R�k'�|տ���h�]k�6�hD�6�T-�vV_5�Uh��޹��_zq���J��ph���Cކ����5��}�*���E��+i�ۺ�zԩ��a1�~?������gi�)_[��#Ũ5x~M&٢@��Ɲ��[1s#~|=�I3�\}�I��iQ�'��$_�)'&�:�E6�b&��w���G�.��ݰ̰��������D���i/�/L�yϓ��P�Vd
��a�%�Q��#&�]������ځx��3;T�Kuu��pm.� �{�W0��Z[�x]h*��˵6�6Q95���I��Y�:�Ɠ-���r�U��XaES-.�Y+�r?~�Z���9�-2*�ޒU0���6�ZTM��ZDD���	���
��V��͹�M�Y��'��(q��l�Ĉ�[���m����a�u1e%��Z���UY�2#�`HEY�,���t�6���[$�����J�@}�,�r;��I������ox��K�n֨��F;A=��q����2]nHUcA�
[mLD���6br1,��8� z�M�ʚ��2�Hz�q,� j
�{ft�2�������ޘ&�����^"A�Qr�~��f���T�0y̌6�G2�i�Sy	7`�"%)ޜ�RۣpuT�]E��V(��'j��S.־S����u@ �Pm�^�	Y"(�q��U7��E-G#��OxVUq��#�vk�ӛ�k����h��G���%�4�LBS�`��*��N"�J�YIN$��N%;df���}�\=m�oY	�:��:�nT��o�*��E�V�mn��&־��n*��J���Rvgc�p�Ԥ�o޳p�)e�=���ۖ��c�8����F�o"l4*�7tͬ���z�r~^�=B���y(��'�T�ɂ�0�K*����I���r��waD�$TbC8d�{�x�*r�׉	v��a��H�dP���n�Ϸ�o�0�/d�vZ1��>���́{�g�y>�\˔�SȤe��@,&G�0�c������h$����RT���Y����Ι�m�z�A����k���
�����\����NV\�X��O(��8ܙI!�&F��!@�7k� 	9<�W��e��f��C��9��w��y ,���m�����8��MZP H�H��G��>�0�iI�	t�/G��Aբz�h)�`M Y	��$��n:�����F���U% trW��l<H��rs�u�nt���L�������I6m{��f�$�À�`w��uZ�k}34�s!�����ë�9����rD.�0�JEΡ%˶K�<����?X��q2�<�����B��m�etJ8�@q��d�^`u<��J�# �Ț���
��!3�1O�%���	��~&�ͦ���8~/�n^���^I��g؋JKe�!�
c�*�`�W�o���*���Z]�+�ǋB~�{�m�PuP|�%�R겆"(H���'�t��&S�Pr��}��[��*J$�dY��W7��C����%�E�l<@g�_�|�z�vjU)����]��csqgl�{8v$#�6�����{c�݃\��sq�����Xq�9.3�5�  �ֶ�X���r��|��%c��t�CGH�8�-���&f��Ȧ���~5w	�~ԣ��\U`�I*q�^�p�[v�RLO%4ثloT�s̟_o#�L�" '5[i��s��G�h�C�H���J���t�K��4�6`���u�I0�Bf�����f�����pp�RI�|��ZP݁���	�YE`x������zd|kq���}��C{�{�j���Z�1���jv��4n	l]���QT� ����C��AR4	ſ7AQ=�b�K�g�--���j`1?\e�rP�Gm@���[��陡����7��J�#��I���in�3��T r���-���`w�rJh�22�	�C���\d!kr�@�y�y���?n�.z��03��cԙ����E�T�L6"iE�wS>>��*)�'��&�����%�L�����t
���)dX�$M�[�2�����^?I@���(�cX��D����n`�QM��y � �U�Ɠޑ�������%l$>�v�7����(ͯ�d�KӶq�1�nθ���}X=��	fU��G�fM�P��P�-� {����k!���$Ҏ���?M��L�wD�H�i�ԺS'�:4�A��`�1�\���um�0�T���ŨW�|_�F'�Ĝ��#��Tn�{.�� 3��5D�ʧ��i[N`��7��ѽMj6�ֺ�
����%�[bi��b9�a;c�<�La2�^�f-���\
w���<-�@^�2ss�]��۴��?ߜ� ���:Cq��9��ͳѵ\���=�\�\;�l��{��~J����j����y!�x�"�'Pd"M�[��\$���īޟ������N���q��$�+U���"��x��H+��JB(^�c�j2�A Y$�Q��4`*ߩ���p��Q~�����n��I0�W�1p����L�>4��'�
���0�T $	���*�H�If�Nk3d��ω�c�z.��d�\�j��ĈLo酔�\Y�|�s���-Ӧǁ�:������xЙ��ĔH@�%w�f�R!ť9	9�w{&,��}*S��}]���"+��IGʳ*���)#���S�v�r��给�34�� %ǅz�vlLjj(x��.Ir^0}WR����	_g�}�3x��;���{�4�)[k"rTw���9O�����v6����Ɉ�W]L���[�4{���O�-D��џSq#L�Y�	I���@��U�ܘ(�e/l������@*&�/����/;l��G\����$�M�ʨ���;��❫~�m���),���Y�bj(�R��+�]A8a��(��u�;�w�m�'B�J�b��ٯ>��J0��H��}3��	r&)Q���:I@Vvq���F�:mK��v�uL��{��m:�1�,
�ݙB��ɺ�5�UX7���ٻ���
p����Y��c%eq��vV>�p�rg>�F�K������ "����zJ^i�Y��~;�IrZ'=:˞���;����hp�Nā�� �DZ�5p$�XᏮ罭��k��{���vH<&~=�����,-�9�i�[��y����ZSD%x���'2_-��%��On=e��܂���i��{ڡ��n���+�9	ٟU n�VW���;-����6�.����b{���Y)�:>� @ʹ�O��Q@��$�aZ7I��l�b[7hV��|�zp��ydLxF�R���Iw3���KM���G�Ϝ1>@Ӑ�z\zZ���<���~��۫�x�*�/&X86J���k������x���&w9�k��sS�T޸,��EC_OT��{7|=!�ّ�3[���B��(l��'`A'�Oz���e�Z,%�-�=���L�d�I35��zg#4��P>r�L��Kщ8i�e%�_�{y|�� e	�7�@V]U��44�B(���|cB�ao�_��m3��hƭ��dUA �8?�x�V���{v�t�����*�>��w��y���`N��O��zf� �JcW����.�|��~�B�\�)R�1t���s�n`m�]?x����"=��`���Q�'x<L��s^�y�z=_��a���Kls�/��v�����$�K�k��l�:��B�0H�	%��Q���Vo��
M�����k��߿o�Wܳ�d��t��/.�˹.Y1�7r��_�s�� �/ݮm��������s�7WUT��I�D�rV�L�$�A�OĎ߽�3��7��m+fz��A+�.	5��?����I��6T�t�DZ�����
��nF�3H%�[t���3��LhKrC���{\O����Yl׻O�&�'�A"��O����孢M�V������I5���d|\��k�|���&(�H0	'7�zk�Z!����/�@FH�{TȂ�$���_U�qg�T0�I�0SB�xK�ᒳ́���I*$H���%��xy�/��7;~�9�G7fw/j��Z�p3�i����=�?nM�����/޷&~Lڟ0P����DWIg���@쪨�@��Wo�Ew��j���,Y#�/1l4��0TlN@>3��o�^��:����`�Ҡ�$8��@�ږ߭ɓG���@:J<�j�G������|At�}�p�21���;ךI�Wf���&��Q��Z&h�i�^@��A��(�?��-�T�V��8/�j�w܈�`�]���4�9��N�����J�ܥ|�U��"���߽q*����hŵY�m�}R��c=�t�uOzfD7o�ݓL�������8��}uC����ė�-�x;��+ �<�/4>�[��^z�	{yhv_��8���XU�]���Ҡ~Ӻ]��W\O�S��\��rQ=$;����E�
����t�a�1���U��ʸ��2th�*�Cչy�����3�}�T	��\�`��6�؜ؾ=C	�N� OwJA{N��s��cf�&����JFp��7��#�>�""�WGݓzEP�Zų�E���ٻnE�^�p��4���[dʠ�A����켵h��s��Ϫ�s�Ʉ��b�������4����ܒcm���Y{�����R���9��n��ʭ>�+dL��̵SuL��ͅ��9�q��Cd܋+M���j�!r�u*�!5UT�.U���UUM�.�j�Z���T1�kv�&��u�1�'Xn��5�p6�P�Ҡ�LV��i6�*��Q��TF�n.D��ڵ3�7P�Xc<g��Y��vҬ�c�/I�$�4��#�]k]�0�w�=������l�O+�������f��v®ф�=-�r*v�ld�.$+ �%\��#�gI�ir!̣��v�j��r;@�[�*�q�ۍh2�
&�[�9]:s��,�<k�	'U�2SWϝG|~V��yXB��LR�ìlRx�E�s�ݏ]�ٍ����\.�9�vw�[�0����'���"Nу��q��P8�-����.Z������,h�7nݷn.�x�[o2[�hi|&ᝳ<n]���^ۻVH2����������<�n{g=��8�A����]��]����>#��JB�n.�V�(��W�հ��1�=[;L�1t[2u��Ǎ���Z;]^��Ժ�a��'Vܼ�Y����'u�J�ٷU�y��v�q&�757H��l&x: D���1��k]���(4R���z��rdb�������Zvϔ�>�МB!�o/�z�"����_RX�m}!S�IHG�R�ݽJ(���p8|�B@!����V�p�r�4E�豶K �_y
�z���sR=��Aoz�ז� t	�eN��KX��6�q�������h e����������,fWmEL?v�G�ɹ��� J�{�
���f���e@@#٭����Ў���"쬋�T���,5�kTz0%�)n��Ԣ���퉓� Y��FÉ���
����.0Io��sub3�]�1�#�E��p~�١ �f�W��Ǖ�_�m}�>nd�\�`��H�e25��.���}��K������ʥ�:�&M��L41236�R�]v�a4�6xr�I��f;�fԏd������!�f-.�Ha���{�i!�vl��3w��K���z��]E�T`�A��|H1 �-�B0��%�4�����z���ju(�P��V�����揆�oB�7��BGy����E}��N���?�ݹn�OV�0��n �ܖ>$rW�>$�7�����͓���oq[0���4.�8��{���K�g>'v7��M$y�u��?	/ѻ���_ >�e�N7��#�m<����Lr�л��}�6�}�a\�1����^gD�޹��-����syE`��e�0�9��6˫�h$L���o\O��
I �� r�Ar[���f\\��n���#�.+��oFX�4�'>���sş]s�}��;�F��:\Hv��v��r�7g\繁�B&�ܝu��q��z�mU�>K#�$�]�L������{+Gڽ	�r/g͐C��&݅<ޤ��$�h6�e�JF1j.z�c�j*�+���6PO��$G���QÆ ��n�eB[_���V�ãl�l���x�	X��d��I��@=��[!u(T#|&�W9�\�c�%-�S�k��%)  �?�B��dP��Z�\��Kq��<�Wc|�-u�9^�5�B};�^������N��D��2V�T��6�J��YH�
O_O��I!�6XQ�VX�C��g��d�lc�6�	&%��2I�m/T�l�z����C�6z���;+��O��� S˹�a"|D������̙��i�Y�P;ܯ�	*%�	� _���c^�U��1�t�*6{��e�j5����B�l7��a�m���(q����OD`s+�n	�m�Dק M�FI@�?2�1]qۮ��۱uq;,ES���3����o�������+h)��.��,�C����5�� �n��]�#}���$$���u&�ރ\��/���2�f6*��:7��+����6h;Щm���3��~�C�.�Š�"L7=US�'(�Q~����@Y�~)��x�
L�7�NBw*��f�$�mLM�Y��������@7��Y~	 �	�9�i#�B�:꫏�&#?8�6��S*�5�^��T�4P���^e9�
�X������p���X��[�2`WSs7N7��Ο���>�u��m#�%�T��]&ϫ��6�y�m8_*�D�F�@ks4��AJ'8_���}�o�T"HQ�V����C��6�e�P����WLs��>L(�x0��c��z03 �nf`|=�Q#7�-\@�������9�x�
��i��cM��������U����`<���Ș�ɵi�;h}TDO!��x�}���|9��c����-N��Ww����6A��\	̶�^����l���Joy�P�ݟ/;ĺ1�%]N��~V�)�(uڲg���B�SP�-U��Wfu~��	�Ҋ�o���$~i)�[���̜�C�}��$	I{�1�ѶVSI�-��1jOz`�~��|}�x�u6Di�S�yǗB�Š��ܺ��[�_*����>�l�qmv����ڡ\ l����Zbs�II?W���G��4d^#i#��u�6��U���0V3�e�
d�gJ휅\RM��s�#���ܘ�rL��]�l����k��ijL`��^k^͊*r˾��T�p�%���R��r]ʹ}c�Z�p��~����Ҙ�Ӱl�#�p�n�k��f[�ġ�d�l����V���)���]�-P�������ɨ��uk.'�'��dFz��o3��5Q�"to|֪{�aL�_�cqi(��� ���Xȩp�,�x�r�n�L��+�=6l��%��\�}S�K�����;�wb�N&��'�L�
gs;Y�ka�I�$r�s�eh�jC�v��$"Qu��%�ݟ���}�(%���6ǣA�tql��PZ�\ۦ٪��r�?{���ן�H���6�"��~g��w~�7�Op�UQaBY��N��)��m�{g=~v�h�b�~2������sob�G����p�$E]I�������5Q�����і�f�=s~��P��90��O�a�K�$�/1i�-SY�>�X��\��&�k�_����G�U�9刳��quQ+&EW�kμk.��a �#�i{��&�t��I�֦9ꩿ}���H3�`a��?8�F�J���9]p��ߗ>N���s�2�$�TL����"��C �Ndi3`I��?�~��k[��bC�¼M{ͳ)F��Kq���j�\�*)WgGx(��!��&�}3T<�'��K�gC�@7dZ�j���dG��G���oM��q�.5�l�ݧ�\p����|��(tܠ�I���K�aU	I��c��`������&FA"����_����]ꬎ�=&�@���c�ۘ���b]�f)�b����M���2��2/ �N�:��ś
�4׈��c�x,6ЦҢ߽S��rj�.��CI� �����=�~��C�;���oŪ@_UUt���s3O�oה �zgk.5a�t"Q�{�NA����0A}-� �m�H)2����U�SJ�Z�3Bud���F��O[r�l&�O�&#��L����lc��e^y�%�ʶ��p�#��0��'�|e�m�����5z�<��H�]O��u����Ϛ��Z&U�#)����{3K�|�a��i��z��qci��0���u��2�5&�@z��I�_��l���j�ٷt���%���f����e��?
��D��O��Ϗ��1�i$/}�� �C�B$�sl_�(����:���F��u�?:��
�nܡ�g�kR��l�;Ru#9�d�k��}x��mߋ�~S�{Cqս,?xb��QV��$�(a&	3bv��K�j��%�ؐ�tP_X�8�����K��چ_	�lN�6bL�p(T�ix�N}X�"�U��ѥ��H�ѝ30hB�&�&u��b�����*M�T�)��:�jr�˸�7���6a_p�F��$V���ux�2ʽ����#��&�����!k�{v+#��e:2"���l����tLt ��e~���`z�[b�,w�r۳I���9^u'�ч|T,0@�FvI���7+>�T��1��]=�{5l������-�60��/ ������F�{��W��zѶ�1p�#��d��퇣q���!�ݱу����������D���0#I�H�� ��@![Kg��W���{ߤ㵼��9n��&�lov�Pe��D{�B�0�Hl�G�����}m_�\�_*�#n]e{]�T��b_�oں0!�"�l�r�a3�.�hF�$)�L;�ܥHV:��6�
�nu�Q`����p'�.v=��y���nl�E��4b�(v�V[��ͧ�y;��y�lxM�APz��zz�g��g����:��B�R��3�P���4�f���3B�|��.��蛠v_�zЭ ��h���zL�Uy�[T5|�<e"�om�Ë�u��J�(SM2��'�|H��Ѿ�7]LU��x0�5�laj&u(019���6��ג�X�K����t`���7�zx��gv1.:����']�!�j��F�޵���k��|�5�J/M��g����Ve��ݖ̱�Q22��9o�~_z��=<�#�+䍊H���Etg�����|�����k��B	�F�)�
^.a�����0����-j5P�Z���9��7Yh���1��s���ɴت������4 GR���P�=I I�:��Y�g�.�=F�t�V%$t$�f���j=��`��Ҏ[�]Lu�����U���&2	����7&5՗l���&o�Z4�$h#
�UKr[��
�?�&N�m�\� �F]6�a���ˏ:Q{˪�
;U��$��$�<���}�~�*�;9�A�i?��WrU�AE�F�)�����,�B�l�!��~�_��G����&ڑ�ť Ř�%����鲟�b�{]S_�HE��c�azь� �Jz��WP�{��v.�(�Y��6���7w�vل�{�9���ߩ�P�~n$�@LU�k�^�y2*�}M��BF����:��a�m]�Ұ�(�f(W&)	ӍHN�`�TGW�6���x��pq/�e���m�h��-�>��Ci��I1Ę�@]`�J��3pm�k�u��,K3��	 ����sv��q��<۲C�ׁG�Ҕ�<"��$�'C�V�,�Z�k�?���nL�Y�DΦ/]�ߞ8�v�KQ=��@hU@� N�|g3zOL�$�`U�Km  �H������TD2J&�a��N�v֧�WͲ~8Hj\�>&ɬc��u�"`��+E�ﶟ�+�O��x�����t�$��E�8��q8��mP�T7O�ېyZL�����EI1�9����[n}�GՏ~4덶��wPj|�D1V�Oƿ�A�Xi,x�I=Wi�U���6��I�E
�
ԡ:>������+�5���?�(�aۻ���3I�$fnR�4� /� ;�5r����_d-��f.�770���%"��C2�����R~1ڐ��9��bHOPt�(�$�'��	Ty���I(�>�B#P`�	u<���H`�5Q�(�{�3�b��������f(�J̕�)���)� "I�_b�9���]B�g�!�҄�ĒM��(�q��C�0:	x)+!R"�Azڍ�,��"�({�w��K���2\�m�6F�Xԙ�ZŐ�f*Yr��}���y�e^�Zng�j���J�}.�E'�_�.����|G�:���&	1�[��7��x (e��g4o�K�U��촸�ꓳ���V �,��+W^O��ȥU���,�������o�0^Iڡ'�U'D������pc�j����
�nI�}�ҪT˯c��AGK�Pم%�~��>�2�*� ZH�����dn�!�N����J�lRkA����w􏿬�X��LʌL�"��1K��55Gm�V�\��'5v�ȉ���yJ�ȨG�|��c�ג�8(�"`���̕Z���P���+�X��*!I~��"�e�L�F�`ܪ��= �N�T�Η�0��᫾=C^7�5T /_h�`Y�y[��br�N��A�EyX=�M�D�QJ����s��I���-���8��6꾇�ݺ��K�������6F�Pɐ�b�f�
kl$���M�����}�M�f����?BIzޒ��lc3�1�}�U��^2I�-�-@�����8θ�Nt⶙�?i��[GA�x��c�O3s�+�.��5�kÌr�w¶	و<h!n^m%>%��;M���!��b%�"UX0�����F&����F�Z�d���9$�#�{b�꺡�������{6/]<9�a�"�c��Փ���!{Y�w>����Gt�}�Il�O����y�4��v�H��8x�"��F{qD�UuR�5Y4�\�T䉭ͭ(�Y��sxM`a7$cq�p��أ`e`ݓ�M��	��k�;�5u��g�
(��x��kg�=T˂���mN���t��ٲe�ٗ��n8G��T��|g}�ǚ��
P+C[�pHC/����]�,3���}s{|tR����u��4*T����J��P+��F^C+��N��+
��Z�bc
	`Q~��6F�����g�܍c��+��Q�Q*��	�d�����Ղ���K�(����2b�o2������c��Ή'�����f���n�ٓ��Q��m�)�����i�0��Y�=��c}۔��CcX�N*��ۉ�����}$��r�:�F�"����ؗPK��2�y�2�΍㉸)8�T�.٩'��V�����ÍF��4�fkO$�'	����~5�-;��?_4����0��E
|��j�}�LSn���h�"��{�z����TÆM"J��N��Yn�S���5I�q󑹊(�hг��:ǑK��[*L0��D�Py���%M�x2�%��`���]WЊ�>�$���-�f��[)��2��d�s�?(3.?1�z�͚Q��;��m�,wa�;^9��3�h��迕VN�YjsZ/̯���Ә��\v�7��@k��s��z!ݖ��J��\OU�Yx���]�xG��nu��D�ę�6�mXiם��'�q�K�5��-�u7ry��F���c����� ;s}�?|=n<y�B߳6�(�v�2a�uI��L���`�q)/:;���r���*�*�N���[@��-�:�}���Yز�0 �d�b)��M��`����* ��_�9���������Cy��r��U����昭�cDS���n�[E7�G^��~&�ZbلV����I��I�1��9=�7��&[p��O���"b���\�u�b��F>1�q7��V.�<��B��Tڍʟ�N{��ZD��U�"�V�t �`�Pȃ9�u��3y�C_��O�&���K'�$�6�%���M���>��Ȃ*b�#�Cn�f�P����߯�d�,L�2.[���88��Z̵�2*�9;'��[x�W�=�3��A�`�S|ҕ�'����k̅0��n	�O�ˑT�;�1�"Q$�yW�,�e�½�2ӎ��T,&e"����H���}��I��4��R[���&�5�<oFb����~j�	?g�&��áͯ�ۿlP��9yٓ@^�|A��]���%]��%����Jn�����'�5t
^ȡ�\Z��������F��A!@�ח(��X���/𧓯�w��@���4��M���:ϕ�G[>~��2��4-��k�mܝ�Zy;�:�B[M)I9�*��YW�fk۩����ٝwkr��uM`XԁU��lщi8׃j+��^M߫�����w�;
�ړ�6r�g�:ΩD3�M�V���<�`�Fl���J�bf�����{�o�����˹UFP���$�x�gP�́N$v��cX.]�V�����us{]�x�s�Yk+���xF�p]g����]��o�c�3\�k��|�SCIPg��8�?=CVIx���Z��"��u���.�b(6.i�L�Z$[l[C}X�fo�<�.�z\rdр�u�q%<G��ta��ZgF���0�]���a��v�]OOfp���P��3-��u���%�7dV:�&�^���r�����,]K�ڔ1.5�V��<u��e��Un"DWX�V�8ɩ���*2�ƙ���Z�d�t���i֪�k5�Ь�'VKku��j��t]Y㛗�>�U[0#��6�v��N.\�r�]m����WJ7:N��n���݌�Fl����>�q9}������I��+�Z̥�Ft@�-�Ӗ⭂�q�^=m�	��f\�	+��b�ṫ��m�n-����j^�q���#����f�z@�sk01=ۢ�KZ�a�u�	�.��k��=b^�Q�^��8�$�u@;y4�qW5'SnG�oIc�n
u���e�n���6ۇ��5���1���w��pz=��c�[e�z�<;���8ּ��{77�ݰ�;lN�ܱ�@L[lX��*��_�cZ������������ƧZs�Ѯc+��מ��:��۷�ni���88�
��Éֳa`7I�A�vs���9m��t��47k�^=u�9�*\a��I�m:o1�F�����k���St]c2�0m���hI6�т;v��Nw�<u�Woc�$���I��3�b�{�������11��	3��c��<|hܬ�J�s	n�h� �Z��ϰ��ۿ�fo���sR$���P2&���ǚ�X���&���ߟ�>�ilw��4��E"2�:��$$ �S3�iW���ֹD��0`���dk�����J|=�6�W�BiY�Ssu'-QeJ�,���M�$�!����R"��ۊ썁�=���85^�%��2L�k^����'O��
��p�
w�i�ױ�K�ZMcG7�lV�kFm�ڛ\z"4:IY
7'�"\�����(��.)md�|�5v�A=�UD�8-q�\(K�� N㦶j��Q'�D�ʃ9�K���!���W��EGG��m�x޼���o-O޾�wQ��O6�[G�x��|�tn=�×%�%ilu*�[�*��0uj;CՖ�j�._���5$\'���o��x	aV�����qj��˄�Z�	��hB^W������^��6�6��j��'�m�J�H����!�֖|`�ӏ&�8%��H�9�����59����đ?�t��'��z���'��}(R��2#Or>�g垼^�^�den�dB+"b�5-M1�Հ��˞�֜fB��С�_@)���%��&�z�%�j��.�H��o�:�*��3�I��ƴC�T�
�b���Y�ȭ��»E�Hq~��â#c��С����-%���쉇��Dw��-�)Oĳ�HxM���� �g�bA���z��i�p�5�$����E7���E#L~�&J~��T[����֕5R��9w1��{�,��։pTCaY
	��c#��z�}��S�z۸0e�تg.2O�����7껸\�u�	*To�(�X���v���4�ž�ʖa�PL�=����}?�f�+��� ɺޔ�� �����'&@�֔�Ŵ��2r���y����N�tz��FĖ���$�Ĥ��L*6�q�ZH|'m��7[�����Tkž�Ù�.�K�����F~E��-���I�~���O�du|U�M�4��7=3,%㝊F/&�	j̿m)�J�V�4�Ym��\��^��^?��r�B{�?\6)g"�md�H6Ъ3ј&@�{��"8�|�l ��N4�)-j�"�%|�ߤ����K)�<�����O�t���S��I�IԽԪ\�oRB
�ڻ֩�oԟ5>�b�g��MC��ƥ���mú��kw��M^�����S�Ͼ&`�񃤹U٫ު��S���&ȟ��_�-�
�� �s��Vڪ-�H][��zw�E�!)%��ܳП���.��k�B!�N��7}��w|i�\�:Sf�Khʨ<�n
�i钽J&(�Y�����m�,[�(1�B�����]����Ka���v�����g�보�U�˳`3�޻W*�ex9"ƤsM���{3�����klY9J�4��9�F��$K,���L�`���?9��G�b�^H@Q��d��锪�&���̙�C�ZL�IOV{;�d�c�Қ��K���EI�=��l&��Z@xA�L�[ym�,�M�a]-�)�`�1s5c�I~Ue��ϼ�2gR[䬃���>Q#o�J�P�O�p�%ԓԄ�}j��*����%Cc�������j4D�L��{�@ j�BXc�V�K�7*=R��<�4�շg����$�Ҏ��b��r~�'�����`��G�EL��7��I0�t�M�6�ēIQYP����$UT���}��>�?Svr�`�r���"L6KH ���s�9둹�2�)��G\wB?��?�
�m��ǫ.ֶ�R�ۗ3��ƪ�h���y��\;�3��j�'~�0L��	��so�����6!�[^	z9�Ut�D�&�;o#���R d��IjZL��*�g��4`�1� [�Ϝ�n���mD�}M�8�j���ҨH��I�ѭ<����FÃ��B�	$�9h~:8����{�n�Ja.z�����X�BƠM<��A&2[~�R�����lXթj����7&��T��%�Oox�w�6eJ6��Ty��.��Es���t:��k�dg3*D��]H��*MG�k�~���"��b�L��x�!Sk+9��X����
��r�Z���qҝkc�`��];S�N�]�Aj xCtm��K禣Sˇ=\�ܿ�$R3v��+���[�K�v�od�Vp��Xw\����w��N�=�P�ɖ��d�6e��_Ʈ����c�e��2�?�H�8H�~r���j��z
�H�@K1�O_�*��(��G�-����ͯ2���Fv�Ƣ�6��}�Oj�ԑ'	�{<����!�HK���ĕk~�Kt�E����[��H��>����@�3qH[��Ǐ�����8�g���H*��y���)~���ZL�_��~���Rk�N}V�8���jj|�;"�K��Ӂ����ի�ɵQ +#���t�
C(R��ދz�5cW��)uJ�*��c�C!�~+���) 37[>V$EL��F�ڦ然�3i�4H	�[-�Lp]y=D�]E��ā2��i�dd����Avi�	ld$�����F��]���V5��\��pfz��j���cuUki�w=��.c��p�fu6�~It��m��V�T���Ķ�(�ʖ�.���R���n�!j
SwUU�!{�ŢT87]�Io<����}O,E���&8���P�9ۿJ��}	#���e���6~7X�W�-�;
gU#�N�����eu��W�M�Wk�T����	�>������Z�~�R5��\��2C��,�2�&5�[U/��-o�y���JX_����3��{�Wn�F��S���)i:kR�$9�n���󻩃>��Al1¤��TɄ�>^s6'tL�D� P��%��l$0n��Ӛ�Z�	il..��(p!�T HM�W�{���zz���(�9t���74�$��eTm��&I���Hi��9�dy.�7�}��N��o����<�e�n�XH���𕝓9���d]����n �l�5=����%y���ف*��콹������wP�߮���%~I�$��ȜRK�$$*ZH�;>ml.�H���(䌯0Үw3/`�yu�9���]��X����H�&)&]�x�Iq����⏽���șV��|�묗�/[�	�
+�TM����%C	tud��WR�ɧ�ޙ���Gn�&g�K��s���m,Ü�%�H����ta�]%�f/,mc�{�S>��7�_��a?��P��ު��S%km�B7�bL�����c��U̒�{=Rqʯ9�c�(�\�9�籒����J'�]����K&�1)����b'�U>����Q���bR���͟.֯��=�>l2���'B@z�o�S��I���C�"�q��=P����}�n爔}�[ ��x�J��>}�֠H���H�1�n��݄�M�d���7��,O�(("��<�\��zd�U���f��`;�0	�u�΀%׺���m>�D����Y2"�d ���Tx�̨�F�*��a�)#��P朘aX��	7
��ܔx�d܃�a8
m�r*[A�揜�Q�v]WH��e�K�����&'Z�Z� d�?I����/_���^���K> Pt�ٯB(��D�y��篴b��˳i�jW�ơc��,����\b��됹�g���%��uu�X���'��_]�b	4��P��u�D�oO�RP�D�߻�ګyȎ�6	�I>*h4�~ˣ����[<��Y���PD�a*������|��V(���Mm��4d���3^�j��O]T�rb��@�XM�Y��*�A3�$�n~�q�P�W�f�>�M��)`�A�>뵵��"@^�����6�nE�EÝk"�qi�ԑ�1whlc������wy�����m��MO��B��H"t>�ğ�7�@��S����X������8�c[	P�Y�"�1(X���^�g�y�v��	Q ����Ct���K�� ��	.�����]RͫZ44C	BA��~o�e�B���K��?U���M�EQ� eP\t_�v�G��_�<O��w���#p���+-;D�
�G�&M�\���_7&pWl%��z�\�A.Y�����IK�0����y;Ab~��fG�~m	j�@D����Mg���9K��ą� �>��9%��?~���-���Y5�̲ae�W���𼁲tN:�
���!���q�iX ��8:I �Y���
�R�+��g�E���^��8W��=r⸆�jom)�Ǥ\��p���=�a�[q���M��۳��z������k\*d��\����Ƌ<����#S.\�Ad�+=�~[�[\����VԘI���lXn >��ӄ�*p#>��-?w�hמw�f-�bD��+�C���O'8%U��K�D�>��;vT��n�%&e�#zF/�Fd�_�]��=Isb�Ni���N`J��i���!�Ŭ1�&o u�T�P���m(���:�ۃ㑄�Ķ����ʙ�S�R:�������5n�W�d���t�	�)�YlЙWG�S�}��y�Ƀ��Q�M/|@�j<ڏv�;�o����c�!�K5�t]E&�&��["�~|���:7t��,L��
��Q U�$�Tw���??~�Q��.�Y�����a��f��m ��2��$����I};�ހ�a��@�R4�SOzʲcM�r����!>�n �����z槒�
��g��2�k��_��"���$�	��%M֏H�j�=k!�Y��Ģz[�z�{� �y"�j\Jc�F�6�����!�'EPTiz�>G�W�`9���i��?$2|�|����4˭�	����s�BO�|�� 7:�d�q��tS53���g3	�%�I�cv������ <�S��0�w�D�G�� ���J<XT���O�vm/E�'�`{v�@&c{���՚a�ۘS�g�R�����>�%_�v��L�(��F^vKr��v��c��=��t��n��,౷#�l�:�9�V7>��K�vvȮ�6n���<8��v�Z���6�ۮ�1�yڑ:��6��l�I\ݖ2�*8$�,q�M|�o�2��>��-�*�&���={�KIlA�(ҕ�
�m ���WC)�Ə�z&\�~���sQ~���*���c`l��1=햀�M.�S 
 mHq�|��$V�����$;<Z���� H�5��Kə�{[}���s�m�̬���l׷�e�V�c�@s�«]��i���I��v�rV�������w�k�:}F'լ� ��>��8�1*�"vv����7���|�*F�CY=�ҏC2٨���zgb�����!Q#�P .��!7���߸\ �8�%���f��e@	��(L��K����\,@1��cRپ���a���|�>���L��CWn`�{ۂ��V*�F�k�@��%���Bn�� ��}�c��39�B�(�`�>w^��=���F���U�)Q�+��'�+ʰR�9��q��}�����Ap!����E%���Y�H0NmJЏ�xk�`�`�'�������ޟL�4�yIT%C��ws���J��j�*��G��hVe|��ǥ@��0{�g�����&�ԘB:�D�(��eCh���s�J��x\R�ۮ�ݎx�����kLH��f�A�ቁ�1U��Oa�!q^�w�&-|!��bZ�ݓ�B+�z�87�"�E(Q~���G]G�6��}]���84��j\�{�O��1о~�葽�\�^w�	�H�qp>S ?�Co5�f��9� i��V|�E�ķc��94�D�io������/�۶�*r	���\�$-LX��P`㝏6���Ī*cFzTUd�+�� ��	b~��r5(��"��bO��@}9N�Cl�B~���2�c|�2� /��&��2"���B�18ׅ��#�I�A��i��W�9��/EU�3���y�'@A$ʫ��z�f�v���`���:�}eL��6)M�\W�oy	g�zݒ�����z;�א�	�����&M�Veu6�C�	 U{�>�/E�cǼ'P����6���<�ݨ�hu����`�� ��d�ǂ�F9֛4øWك��DA^_c���ˆ��[����k՘�\V����ۭ�un�6���Ӷ&N�Z�m��<HԀ�H�n���S!U�^�7l�5ޘ��L�8�(�3;م�� ��:�*��D�*b��%�w[ncˠ��W}�F<�&(�UԻ����!\{L��5t��ɑ;a���0�k��y������3��>�5�F��Qx����X������S�k�d�g�s���f&��:��ɒ�L��-�ٔ�X�7���+F�ɖ�M�
Qj�@>�2=��l/��8ͧ9�Rą�C�kP�1�=�-�frm f��6@�On��9�:(�WꐲeZFs�~���H�zg���p
�S�SD�|�I�GJ>yGc{��(A=
�b�9i�W�	u�)�|�G:���9v��!HCKI�~����zЄ6��C*���q���lr��i�pɝ�����-ݣ�!�^��(4��-�M��P3�^�Cy���{b�8٥3s���Bo=� ���9N���gj�����L&u9"m1Ov�C�
�P n�R�TxO�aL� 4 �S����h�(o�i�S)���@���0�c�1b�SS�}�z^�r~�=Ղ�?V��g�`�6���7������L�����I����	�Xc.�W[����Nwcx����5%F��T�:p����c��O���O�M�7���	�sN�ك>�+N�Ό���oO+����n�I.�],�"�;�=��l�8�X1#�	�5E��n	�����f*�#s�;�;�Of>����J�{�\��å�$E�����?J�@�,/x^��eAY�=��vp�`lE�䝙�\�3J��Q�py`��"���@��ӼQ[V��DV�zf����[�N])��V�����Tx��#~��߲nc&���S{�]j�(�B�6q	�Ӣ�z)6��R֬����u�n�b�We�t�4������ìW�F��Jwx���T�68vj�CW,�f����Ѻ�����Pu��s��|�Ǔ�9�#8�n]W�r�쬋�R�UUT��Pa:S/a���<�Z�Iw`*��U&F� 㶀W���Ǻ�˸��2Ӣ�Z��Y%����������VU�iV�����lL��%�-fw7�f�S���s��;fL�\+̧dv	�avP��*�%sl�s�	�`YA͌j�yzJ��[�U��+HR4�	�֔�Y�c�j3)tK�M���(����Y����[e�s�H�vLcm/<����0�|WZ�y��y�z��6��r�æ�Lv�C���YY�fX5���le#.v�ȜNܣ�\���ޱ��2���������w93�gٶvMq(q�;��h��n6{f4έ��v��s��3�xx۳k��5�'Ü�g�m�()����x�l����uY�\e�-;,��v�q��;�b$��V#��7"�q9.q�u\*ÏGn���	[[�N۠�M�Dm-l����(r�$�'��m���������'�4�S����mj�j�7D���V�=��ܝt�Ek�v�K<��]�/Gcq\���Gq��ր�iG[i�:4g�m�Z�ey[�E����s�챱���	���C 0��u ���� �M�I�"����Қ��SYe�}�#)pz�����ct�AM�o.�v~�\)�ɏ��a<�5�Qk�16S9��Xx�A&MF ��)�����b`>W�����@�Sv�)/My��`P��A���t;�\Clh�����Xā��'�p`�$�D�_Ď�"O��zS�X��S�$+.%�a���U�18���C%���ΒO��{Ftiv��='�74�X�P+��P�F�ϡyd�NG�u���k�K78�Of�t��o+��½���q1!���N�tj����,8��q�=G��W��ؽ����%:�ԂL��P�D>�Q���!URE*y`��mW�׳�"���B����������qkp�J�^�1���.1#y��mg�`ǡ3�A'?(f��緵ٿN1n��X��Di� �,�\iMy�7�\��x�3jm��gg��2 0g��A���/���P&;|�+�B#�:�I����v|D������O�@d��U��"=��_��P$�����X��Ʒr<�Wv=}1�-�B�+}�j25O�A�D�Vb�[��lXA2�)���Y�뢕�y&v�5��D8��܅˻�%[֨0�&�畽�9�ٺU983l�z���ԇc8z6}��J����k\n�8�*8·@��o7c��[����*@�	8�n㱐z����ٛ����	�^�)6}����:ގ��_�F�Ci����TLk�)�Yك�m�ՎT�bf=��N��/����\:\�`��W�B�#az
*���N��CG��KP�f1AEUi":=m{�kϺD~U��!���DVR:^��Ļ�g��|��m�����,��S0t�B*8�sל�'��K
JٿA*�[��6����1Tn[�g^�E��11�~~pL����"G��׮����S�aL����F6��zH��	���|&Moy�(�����ɞԀ8Tշ�>�̆2�B���G����z�&1�A�x_��	+E�:�TN�m�	��j���v��c=X*�]X	�����4�7j�(��UN�D���M%��x ��R�馼�����Y+7"�ȏ1eK��=���T~|T���9C�Y��M�t�q$��,dl{���X"c�{�u30������$t�!�x	���	�4�F}���>��ț��̯/��]�!T����(�iЂL��*�Q���1��A�+�,���],�Ɣ:.�]���ch\�d��mN�fkܽ�=y&�S�����%6�Ve��.�S���Γ}��[�#D<��#���I�CK��j9��C���I�lWIg�5=|��0�h��UPj��8�V]��J i_��Q���>�1o#a˓��}
G���K���͂2:��-�NmɘD�L���V7xF����C��0��N���! ��a��m�Iو��9�DZIf�m�&'��t��nP;�=.S�'`B���V/L��=��,���6`u"���n�h8q��ò���_*+ڸz�(@��L��U~0�%���b*��U��0GA�aF�	%t�g_IB=��l6�v�AUw��.텧yӠ\�'��ᚨ!@�P7����lz���<�"R�\�L��GA���+X>�O_Y�S�� n�7�i��m?�m)x4�J�f0V��l��{ɐ�Ă?�EZS+.�*P�A0̌d�N���~�bc������t`��ls��55���wz�O����<�JVܵ�q�e��)��
�rea�;(��z�+�?w���O�p>�����{l�'�75����`�8�5~*��h!�*%��PzN;���ѝ4W�J�o��`Tsh?t��^P*w;I��{C�u�-�sЋ��9������ŦE���F$���m�L���&��/}�v����8	��� ��G�p��O���{է2;6v-�W��o��y��#�b��Ӣ����w�����=�/��#0I��A��B��:#�)G��pkYw밠�ꙶ!�B(G ���}�Nǅ�0�o�8�vCa����E�*LX��ǹ�$!U&	�׿R��!��Ws��w�~�^�,T�P��8������>C���Ҙ[BB�ȢD�����ݘ<�F�l"�&;	�W]Ix�⎹��[��3��[��H��۲��ɠ 	��
����b���^�r+�j��f�p�����oe�O�!"Ia�`���t�����ɢa��I��9G��w�ZB^V�Ӏ\V��n����OuJ�f�ƃy(��ݬ��0V`�*P�(!�0�,*]a̪߳]��O���6�P�04j�_2�0��5�X\�=��4�g�[�n:ȇ.��K9�V]6�d�i���d8���Vt!���\tr"���梸p�v^5�ۓ�@�i`U�*�GDTF�H�(�RF�ꬤ#���^�.�m�W�;+ � 3���	"���틻.ܟ8Y���E�w���+n+W�P����m5�p��O`�(f�5�'�����
�"����rt��T�\�#ϵ�����/�<�s}����P�נ8Խ��}3�m����E�&oҹ�Ewg��jO9|mv2˽��ҜO��	)Q�A�L_�"AuR�@�D�-s�{y����
�)���:�ټb���i�q~w��o�$($t@� ���<��96�6e�π���R#�wp¬���}������&`$C(�w�
��zp��EDʘ8#�032�ǜؽ��
MCn{'3�oQ]�cE�o�>�IG�~8�~��#J�Y�h�#�[dc��r28�|�9���P���-�{0������j�@�p	w��D�8�U�F��1z*4��b9�4R��N�?+���A�V_�{.��.�m�;���k��&-�,�W���א�{~BMR�ㄵ�.�4UXoi�+�O�;y�N7O������מnu�{kr)�̴�Υ6.�pv�{[m�ې�lGW��x�U��s�D+;Z��]����Ř�e`�H�2�����v��Tx���4�@��f��(!���"�m���Xݩ##��h�̿F&`��3;���nb�%��o՜�_�LzD.AsPx�p(��X���q����^�od܎Q�B�l�|�v�QU�X�@�Zή®!�v���$�	=C�pV{6�Ë���Ն,���{��������.�X/�c�
,��<�~G�Wp�UM&k�6�_B��}�L��W@��+;�<;p�Q�yh^>r�c�(0�4�xG-����tEC>�|U�'/M�YP 2R�M�"Iwk�Æ��˲Rv{$C���,�	�������Q�ޘ�$y^eN�`�2;��f��:��Q&6�FO����Ģ#��#�����J HS�Thj+��Q7�(���)��'����)�8dr_��]糑!�p�幃 ��]��(�:��#� ���N'�>e��;�a@2[AU�Ǭ�Ί�3�2(D�����"�E׼t� 5����3V>��}�c!�����1n����Ї���#�ge�FT� p����"�^z+�MF|UE� J�?�bV#�la�b�/T�%�0U�ٙ�ES2L2\X�@�ѹ�f*l����"븿p�4�8�c�O�hQ�����1g3w7��_�� ?�*������,*���1�_�~��z����mDG����
f������ ���� kކ ߼I�`������
�ɓ�oϟ�p�۾6^�6;F�ڪ��U�	Ex�z�o��ӟ�`�f>�$�*v����C_"��s��殽[^��=��&_1�=x9��Kڂ��ɚ�[R��N��na�	��H~�l�ŧ�#Âo�D$f���@���skĸ)�y��Q��sz>��<��U5{v�~�����v/�
��8!+(���.;OD&33�E�u=5f�]���-����� Y��58�gx��M��Q�bo-��ӲHM"L]ߋ�LC�`Y�g ��Y+n���6\N���6-uf�K���#�+���Jo7_�mA��z\��@	��7��C����>P��x��z~^�OE��X"K��F`�$������r �C�^�6�!���LKRQe�Exp���Q��s�u�T�;�79�
XHBj:+�6�n/dz�����r�(2LqUk6.���l�Kb�@��k�8;m�i�R�d���T߼�Mz�1���zp����1�1�}��W��F{�:��!��])��yx����X�p������C�P��m���v�tg���#�T��A \�z��GZ���v�` A�k���^{�!��D�a��SLx��B�����ys���=��.��;��In@{{ ��@�vc����1d[V��z,�s���+W72�!�&L�xd��2�3�inf2{�{>_�K�v\���?g�j.lt�xN,��:�N��Y��IǄf�ڐ/sb�ĀA��*�ݰ<�����N�~�
���|��{��� ���
��2�ٽ8����\�S�{��@�\���5`� }N��z��w.�f,��V��mk��ᢸT�S��S��ɩyZB����x쵙��������i�y�,ݛ g�p*El��A�6����(�]�;C�:�p{Q��r�l����-�7`��+F�n��yR�b@�e�pa��Z8�c�+3޶~�ɨS�Q�}xs����3�8'�ϸ!t8ʼ��^4�3��>��O�+R�A0��E�M�]
Dg*ק���ciH�oɋ���@��H�tO���0=����9�B��ԑ�S���ψl�[��D�����X�xCp�������s$/LX�/�,W�]��{j�!@�Z�5���y�1�|ˌ#�(�͛�,��T�'q}�k�Gl���d������s�:��Nrmg�f��z���%���bf�{qK����$�Ӱ�]DY�cy��3�u O���y�^��)F$��*��8�@�I�⋕�Q��D[�>��
{W�J?Y��"��u/)�6 X�z��g��� -�Q���7�v�Мp�Tx�b����������@���dC�O�VfeA.ٗyf82.I����޾_�)��������K��0
���*ДN�a+���o��!�ʓz�?�s&>4
��j~�z9�2���]"�F.�c��O
'~6��%��v��0�5' �X�(WQ�g���bki�g�x_<�i4]=�zM;�p����qJ��A�Gmؘ�����wT��#��]�m.�e��B)�%v���lOV����wE�kp�ə-$���s���Cr���-�^�XN����F��0�=�:9s��71���|5�X�a���ÉJ~5$B"�K=�����00�cZ0QWD@^~��}���VO,�����;u]"����4�f}{�~�K�3�f�gXY���#9��.2�, 
�,�1Q�EQQU`(�������k��o���p����T1���/�������sl� �K��t"Z-�=�Dp�3�n��-��6�s���m��tj��dϕ��Y>������<�^e(����zS5�����C��m ����Svu�����6.�3�O�`X������/Z����CxS�xB�>�]�Hĳ��;$.��v@�,�b�ѱ�j���jsw]* a6�<`� ��+���4%�X�c��sԋ���S�x�A�zB6ܺ~u�%���K�i���^َQu�����Ņ��_�����A���DXJ���Oy�<�XQ����Ȟ}�+.c�/�;:�e���-��ߵ�*�uw:G7{c5��.��j���=�|J7w�V�ɼ;U�Y췮P%�̉v���(<�&�
���6��@�b�F
((�ȹ���)���R���7]f��uk,n3�0�h�b��)���y��U��IFW���nb� N��B��$���.Tc�	*v�_nI}�$ž�繹��UG7Q˜s�ݑGP^�:qy<��*�����LD��a�^��"�et.��a�=�:<5lĶڬ��8�6}=�����a��"6���B(9ӝ�p�6�zP�L�7��&1z:�H�����߱i��g|j��=]tn��:��h}�����z��]�Y��^Ma����,��懩Ǿ7���A�.uۘ�`��s��R;f��n������K���̕�X��b�M'g�|��r�m��nɰ�UR�j�jUt�Ȳ��L�I�`aʇ� �t�����-ţ��p�3�ûm�4=�kz#a��ڬŶ�����HW)��|s�=��9���n��\��s��n`���V�Q�:+�.�un�=��?����4������^;�n0#���<�ѽ��Fn6^�1�`�X:=�s9g�n�vuk�<�R�A�4V^������;�c�j�0�ض���1�]�88�3��3l�X.c��7/l^=�GN� �9p��ָ�ݎ���p���Od1"]�fb̤���0�Aj8fݱE��V�N;�n�-ᔷ�NJ���bۅ�Ii��C��m��\֋��n�l��]��6f��؈V�@/�UP�m���e�l��Nom¶�7���V�y�f�9�� L�tv���n��-�q���sڵ��G��S#͎��v;)$d��z�*#C��ɻu�0��6�ڸg��[���^�1��=�������m���G9�2M�Lwg��HR*"�
�n�,�����p�eq#�g�WG9��A�ߥ��&�:"l�J☄S|��>���\N���SPG�0L�Sdc-F�a/�{�Px�#~\Pշ|�v͆��Q�a��%x��y�n�5V "�����ﶼ\�RD"���\���1:�h�ީ˟_o "N��z�j&�໨%]��r�����d��y68�=�$$ \0,�&|p� ɓ^��\��N�	��f&���s�<���	�+���1�GQE�s�f�f�	+wt�iƏW�7�RHL��B6�����M�hz;�:�
|�V|7x��	_��&f/AߛLV��u�3d�2����1��}~Q},�L]�X��K8L{�u306����^��8(�m}Q�9��{�a%�eܾ�y-��ǶrB��G�Z�1;J ��"���Z�s��	����w��o�xѾ#�Q�=q��&4����&�4�r&�;[fo��W�9��$+�\�N�ʍ�f�u��&��X��/D%`��o�3�>�U�;v/��Iǽ	�W��}	Ϸ2W�w�qջ=Z�?v=������	b���31�b��
&�
57l���o�f_��墸AE��p�q�}\��t\ř�����{1���8x��0��7�?O�Yо;�%���_��(������M��96#5p�z�[=0k�>D��Uqj� pD l��W��g��Gx�&{��E_Ǫ�W��.����ȧ ]���㴛N:<�!׺@m�DFp[ۏ^ �D7�&B� ��|�]��O	�o(p��?�m�*K&�˕�G:�}��}{��C6�{��Ƴb�~�����6�/I�ԋ�U^��ɥ�r�Ʌ���?M����~�]��͂!d���bCJ<��5�Q����w�
L�҄�G+�,�G�V��V��v�댩�j����޺����/!a(�aBK-��9�s��������^C�f��fJE�q�Q��&Z8��Z�`�d�����jnf�{r��V�f�X�ۖWE{S��vk��ٞp<�Vt���ZC�	�vۋ���u��#j�) $�TZ�@~����}�窬{�q�P���ɨ�Q� �(�90�xy)w�A��Ҝe��{4�M�#��}�%B�ǈ���g�c�`8G`[@��>�����aSH�a�>�:>������!4�����˚�b-,�&MW���sN޸��P6a���Q����T����QЪ�HB@�12v�#B��A�t$�3k�$�	�ֹ\���}�^�� ���<�W�.q�$n_���ۀ�x:w3��nL�D\x����>�/��J�A%�@ďN���.�59G�&���.$G�p2�E��VB�-��g�2J� B�zv�B��x�k��.\)Bki1�Sb���	Q��vr��!#;]��p�ƨ��&lF���~�x���l��AA�R�h�QnQv�	�	��\#������K>�3�߽�1+�oZސ�e��l(��"�N&����ݮ�ֳ�W�U�H�&F:)Fz�w�;2kw�=P�TZ�{(	��H��;��28{85�v�r��gtl��$l�V�dB����콺vi�EtPm��v�7-'��N%�j���I�u�zw<<�i�s7�5ۇΜ���A�%�3�*�B㛎��8%��Z���IC�\�1r�zٓY���^'˯�}�	LS��KA�'�n/��t#fc �I���ǣ`B�{�d^b����ǅA����G�e��c|�Ʊ .0��%H	q���s6�a�^�.�P
E H�7	����	��v�ٌđ�)���.��H��;E���|�g��/a�=���ѓ*��F��cz�5��^���W�n�p�2�d���*�����"�-6���DC��Ŋ��C�-��`��F_�8"��x�/CB�P���o�Y&:C�s�'����2hlmH�*�h"�P�p���R�7� �r���C��Ņ���C���ـ^�1㰋(��=�2_�U��gƁth���ἡ�ڪ���O��Oq�\0
r_{ܸE@�PALyE�s2�_Z�&�K�8[�#5�O̱>:��|���i%Ї�~½o���LR�Ȝ���0�0�� 8v��E�]�F��=��Q~�e���G���Xi�yx4<���M�[��4|_�7����3>�/��^b.�N�(��9�P�_�c�O>IE#�cƄr��y6ڤeU�HNJ��YU�+��e\{��;ߦ �P��7>���$�
`T�"�}6''��'\U���ۨc��7X����c���YB� ��$OC�]�Եz��0��ę��#�����=��G�����KM�}�6/#�q��e0�|���ٸ�`�fݑ���:.�,�.zO�}�2ҷ�/�uwL�n�m�ы?HA�g.x)�>��E�]F�x���.�Q��@]@
�|�N̯j��������xa1+��"Î�h@�O���ǥE��O{)y�p�Bלk��׍H�[N/ �8'�f:�^b�<3 lj���Ûf91��-���,��w�4�C�2����w�
C���$�s��8E�#�,�Af��H�>:�m�8���y�K s���Dq��Y��[T��{fI��}�t�"��l� �,�l�&��Q\%�|��#�?IwlՌ�^gU��+睘����M%,A=/��ɾ��N��]a�;ځ16m1���M���O�]���^�����#��}��L4�����Dϳ`q'��@�i��"ᏻ�߻�f��@��@��ܓ&9���.e�-s2�7�7w</Y���-�.��p�~��,�%�<-]��Q4L��<��[���/�A�^܂�l`�}��<vr�lT"�a�j9�r��6z<�������B
�tU������0T��������.�� E���yޝ˨C�BH��fb��۝�U��"R��׃���j2M,b=� @3Wv�P��6�{��=�b㹆K�u��M����L͵n�ktM�����I3����͏e������z'��L��fk�-�.L�yx��y��2��9����p��B�`����M9�H���h�q�&%ހ�o���SU�q�{J ��������#T�)�X�ȱ�c���h;_�d?N���Wx
*Q
n��1�� ��Uт��:7.`[��#�ߟ���K+&���R��r��	��t@[�]۴��KۜɅ� v��6]r��ػ]�8�;Z�q���+�V�B���v^f��X:���yGW�{Fr�%v��I��d]��ɢv�w������V�G1~�83mi��}\VN���> �5u�r���H��7b�]���1�	4~������AN���>�UJ��(�
�00����@��b��{{x��㰌1[y>�\���j=Ҕ�>S곦<�#�*���x��f��L1/��\��@�_4���&3�v�Oy��w$�-�\.O���ʾ�PA���4x��{�ߛ��&(|'#R����FV����[���G�)ב-�0~�m7���q=n�N"w�Y�i��|��3gň�����4
\�&&$�&���	��<qٹ����ǫ���m�G��	o����Y�df�.H�I�]��3�$t���U۸�!dz�u ib�쇎���V����1�g�E��S쟚��l�����N���Ǵz�p���k9q��,�mep�-�lC�ի�"��R1� �َ�.�&���/#�Y�k*�b�5�qͩ�ނQ\�zk��4�ܥ�e� �pX���6���V����۬��$����b�dZY%_R�E�|5�����wgE.�ݶxvS)5HC�s���V7i��776ۗa���݇q�<�j���R�g����k�u�{HJn�e����yJ��lx�;��\��]z�5�qH��&Z&K��Z7��C�f6��3�(�;��R%V���j��=]U��>���a�� �7�mL/��[�*�I"1}n_/�����V�y��1L�ٹ^w�۹ ����_��]�h�T�B��ō���oi��q]�(��\��b\�="�"�����z	[n�� �B:Fn������i�/�̌�}vͶ�6�A���+��˕J�"~N�{���\N��|;++��ډs�,���d8����0@�y��<�I�1v��K\�I���p�(���
��R8G(O�Z�p�ۿZ��jMe��h�!��l�a�WE�圽�@p��Ugt�>��ށ�nvp>�m�}�=7��hp����X�P�2r��>��H�~�K�V1�Eƞa���'����
{DcZ��xkT�����M�E!z_�?z�M��0���"6Ǐ5P��M��C�8��б�qb��o�?�B��!��T���I���S������ݢ���1S5�)/@�65�cQ=�!��k( �P����ز�nXW ��F��[������	s݀��(�+L%t�~�բ~@`�/�z{�}�]f�{!�d��H���]�ݘ�t�g�J�	bzĕ@�
�e���
~��nٓ�7f�&Տ�ƪ�?"~׏Ϫ=�C�������-r�4���l��g��y=J�`Gt�"��~�;���w>�؛{r*�
�)F��/��:Y��.W!�k�!�ԃ
��p�NQ9���h�Zxq�pw���\l�xۺӓ��ٹ#�H�I�L�Wɋ�W@��ui'��	��E���u�0�.Bv�,W�I;�{���p�<E�WYd*�������S�8&G��kI�]]�r��k���kg�jMee-%w���w׹��S�Y7k�I-��2�5d��s���/&KLf`̿w���w}\��V6r��3�&��?�M���z�i���� ��`�=�1p�N���L�oEj��r����W����=�.w݃+lXK�i p�́}p�X��������nct�U��,_j�Q�sESNT�\���78�%|*n���#!o%ߦΫtm�mٶj�m"0R�Q�A�\!������El��p-ۄք<��<����ίo���Ѝ�� ��g�MX�%� "+i�.�/K�r��h#��Q���R��~��v����lrz%�����Ҫ �>�l��q�����R��8,�_��F�l=���.�5��/d�	R�M?�xr{�V��5�D�=��
�;r@���.@��q��U��c��\��Y�ZH/b���'��p�T��'*��5���m �y�˵��|3-�0g����<Uz�{ĿAvDL�tV3Y� c���� }v���ee�����UxUf�r�����:B�T�c�)q�U\ј�M̝O���U_�Y�4m8씝n��yv��`�+r����iip6n�ٕt7���"������b��f�{�upj����lw�By��T�Ck�T|֮�L�C�Ƶ�q��]]��u�mjgD�7־4OmL����7�ȍ�v���vYBgm�!0f�c&j)*4�3-V�R�o&iD��RU�[�Rg*.E��
��m0]�ɍۗz2��v��q܂��sR�*�v�:��_�s�o��T
l���;zur'�T�w�q���X���7j��/��y��Gn�m��*T�_X��P���W�շ2E�NWI�� ֡@��o���p >]�|}6���q㬬�ʡ���Y�]��gP�w	�6���}C��H�f>ҁ���\�
����|���Үu%қkXf7FJT�T����Fk8Èj�+	��J����h����u3K6���=���g/EMP\�+Z����RSSUUP�UU6��,��n��URFu�v�v�v���r:�r��R�]�� GH��Z0Yۛ#$�:�8#9RLXƦ�Uy�VUT�M�x ͒�1��n�g�F�4��楻I�l[��
m���Ƒ�\쁖R%�Iwc n���i�4�'5��q��pk�xΆ�m+�Iq�{Yz�_L3��O[�hy�-�c�=��э��h�qX"�Om��N����V��B�jM�lzԔZ���	���֞3�d���ݶ��˶컆��B�c���Z1��x@v��7[k��n2���Ul;6,vG]���5G7j�M����D�(��3�Z�ɺ	����8�("��7afꀶ��u���3��zB�v-P��k�+x�q��f�I���=�f;d�4v"�Yٝ�(�UT��ur��^@��6�2�M�!N9s@6U������u���ݭ�˶6���{<"���<���CNp�$Hkx�����������k�;c�ܗ\�ƻq�v�������c��A���w+��GF󄣱�&�p|RG�i�n������a�;.����d��pu�5�dڄ���S�}�x�*ɠ�L�L��]�2d���՝��{1�%�d��o�a�PϜ�r�	9l�-�m.b��lyy�goVC��7ce�����b4�@g����M�Ka8���h#�.�ZC#�]�b�*�q�#��$�
fȫ���&f���ݻ��>���"��|=J�p���"����˶R
�i�b��}0�F�W[�c"Ƽ�h�!��}QW�4!�����{���or:�����d�ݰ��Ie����1�p8�7kF瞝����5��.i��_n6�z����]�4������>F-a�^��w����0�-Ѐ��(ӥJ��,+�:�m�X'p���ͣ)���.�-�w�����"�Vpﶵ�ڵ��]Gp&�%�WY����^����<�I��a.s�Ս{`x�aݭ���C=��v91�H[�%��@�tv�S1s�5c��6읞�<�мu�:��5��g�(g�nu��T�99�YpYka@��BFm�ww�$�]��x1����)�t��.�A�"J�J�h��f�5��Y�V��v"�Ý��·.����_n����v}�|V��=�Ut�-"���׎�[�6K���P�.Ʃ���������BY���2�=B���5�7�|���q'a�5
H�	
G�����>��#G��A�����8#]�^�<��#e�����[a�\j]�/;W��K&�#���@X8���K��s0r�l�ǁ����*���9�h��5c�՛f	�R?=�%�mo��s�)��y�����_�0�.r�3D�$���}u���q(��a��xF&�íF�FUJ�K�P.Lg��G��3]:�'��{�V�˚��0(����U���6������r�d�����`�����\�b����{7�+�*�f��=��J��]C�kmb5bQ�[� ؂�������>�?`w�`d1���"�`�}Yz`�ʎ*��x1M=~�/���"���C.�LN����6k���jBӮ�&��G��8�.v��������n��\�֮�����C�P�DȄ��e�v�4s�s�	g��X:t��`�J
�{Ϧ����I������u�(U��zn����L2+�,��e�L�L��%I]|����j������!���Ӻt�yf�80��:�E}D
�NhЃ-)p��_.��uvT9H��wESz7�����@�i�k"���]n�Sh�ACM��XV�\��=)�m���a4�@�`�DF�B�|�Tu��k}�x^�5���o�Cğ/Ӻ���@�.�	KS�t���*mi���1X?3�h���`��_pN�����0���^�X�9M���-/�f�a�4�j+݊	J)�3�����Ѻ��3�3]|���u�h�� �uD1�:�tt�7C�e����@?�����y�͠!M�pPɽq�f�TX��t�{B�S+�ͤ�N��DQDS	S;�1��
�/Koѿ�������k����u����ޭ3E���v���k���x<�����������G�T�׵U�;�jWK�pJ1�;@*�!��tc]N�0�Ej�Oh��&��W����gWY�7�nd8h�u���1��^ɖ7�����y�����Q��/7ƣ+V��B�*�QH-��֚����W.��m��i��x8A�t�\<�c� �E�
����6�42�#Xd�F3�U���&�`f�V���8��Z��Qm��Y�,�D�3�ᗵĞ%��\A	4F�A�YÍ�@V�Tjj���mR[���D�rg5g�u�r�l���9mfv�4q�]�^gy�m��s�4�0k��i��%؏a瀓s[���'g3ˀ;v��c��I��k�4-�Dި�n�5�J~�����)����o'�����a}5�������+����4�$�v�vAPyna��P��M�u����1]f��`��R��:��Y:3��Z&�<)������\��d�RF���*��M�=�eHM`׼0�(^�Ԣ��2�9���)j�fb�S4����v����F��fʹ�*�0f�-Rp�v.�xr�+da�v��z�3�J�O���:�mj�G�LW�xȋ6p��w�!���v:��B�:�8(>��g4�-7�m<Ԋ��X6/�{�VT�Vh�M�T��t$��S�30`� �� R��}��NS�u�t���mRo�M�t����9���e�i<R��p�7ؒA�РE|�`��-�ԃlMC��n�[D�V縄�'���ط��z	}b��l�����������l�g*vdj����h4�Mqc��6�KU<��=m�v�t�Naڮێ���j��T'&�vv��7#_Og��
;u�V�=�]n���X�e=Ɔ���<V�Ss2��ne�mP(�lh��n~��߻OU�G8���¾W��#k�.�F�v%E�t�X�[��F۸;�0�"�I5ԣq��HԐ>pDM�ϖJMeY�m�GNϮ������ڵR�2I 8B��n��Y�9#��d��ls�B3q�F���v�u���A�m�Bmme�bR���U9�IIhgC�z)1N�G��x*.��sfE/ii�4���i��Ӟ�Y�*p4ui�q6�k��sL��f��rVB�B���8Z�L�+&VLĖe�3���j�5v�J�X��7H����!3�o�a�J8".���&P1��|+��
�/�N(�c��=�ł��_U����7��_f�x	j*���)čf$-״ĺ�E�U�e����.�9R�����b��۔3�BVc
�wV
M�O��L�(m�%76���\���Yۃ*�͐�˨=���}�=6�9J6�zob�ꄡ��ap��-���{9�&#=�']'V�b���4�R���o)eD*�@�G�qE;; K��*+�\୹�!���4�M%��8 ��z�|��r� 9�U�Ncsr��]ҩ�"���������"��;�3W�f��.Œ\L�$qn�[m�=v��pȐp�Gv'�>�_�����)��ǘ��֯a���[���N�\�otAU��������J�,0�+�����1��)VB�P,;98c�"d�O)(l���kX�/bhA��7t0~�*`���,�E&�~��l�ǰb�����u6w�RM�����ky����ZQ�ay�o������0��-,� blT�-���&��>dªMhm\�9�y����ݱH��^�P`L���V�#�GK�*���m�Ί[�AT+_*V���K$����
��Jq���9�����$t��.��9w�2�6�7���~*��H�Ǘ:v��/q}���L=a��=l����ȟ�B`	L'@�1v��>�&�e�z��^Їb�L�9�I�%���	�[���*m7��%���%�H�Dб[�[�Kʪ� `�z���y&�˾&(��o�wK�qm�h�|ʾa-i֒��_�� �_F�"�{0�ve�H������@�~�Y�i<�<v�B�F��v�kB��4	��~3g�W-0�d�r�%�+B\�b8ӧ�t�k'&o��yT���3����`���qbc�;	��?3p\�j���;+�{ޢ>�?_����|mQz*�Bx�Sޥ��
ӥ��?���]`��D��P4A����<l�|g�~᠊�������0�ꤊ���DF���ظV�+�5"�jUfA�d�F<꽷\xk�-�m��S�G�N�:m����z|]u��
6�.�k=<ep[t�6묌[���W�����;i�h`�ZM��0�FϷ��p�e�.�}?��3����Wh������>��g�Ku<���A�l.��K�T/d��U��`.B!�Y�G4�f�d�'�±���%S2pD��m��R�ױ���z�pt�҉�L^C�MO��{�V�*�@��U���=����	p:�mٲ4��wm����+�Osn}�^?wS�#���L�nQ�=v/V�Us��������:�=?o="D�j}$�����Ê��^�O�����Kl���_� ���;�s9�,r7�9+���L�/�T-�+a}��r����P��������p|�5�L�!.2"W!4�VZ\C�����X�1�γ:��U�(�gN�ػPG��~�"U6c�T��<r�E<H(F΋ThkP�.#Us���׉n᝺�g2�S�<���J[(�{]�wf�$ql��7�+�h�2����C�h�)
��/7��I/=ͣ��w>�{Ny��t��v#�қ���%c�n�Wl�V������£����̍v����]�d�l���ୱlK;�ugՖ)\��D�g���&_o�FL�dB��c��N��94��듋&'���D��qQ3)&W���c�E������앾A@�50��}j�բ���pLdfBt����`��<}��._<�$�ka�8�F��e�)\ �`X����1k��n?q��Tө���k������t&�гȇ<���o��-��j�軓< �mF�S4�_K�:�>1��?�ވ��ypI��p��oQ�;��s��PQ��V�"��Y�Y,�#(@���ɬ�̃�k���3��U �������^΁���♟WN*5�{\�a��ὺ AQ_����6�3}k��ț��5�~�:q5��`�hQ1���ͥ��n�)܆����!�c�����`/��#�%����k�j4X�+ @T��B/n��k�uU�Xva8Szw2�������剂6R��C�8����f7������ѻ*}b��5Ruv��a�c�W�]-���>�����q� *����UZ�ӳ#D�ӈ��/�{&I�w4{܅�(VW
������f]εYW��r�s��^7��N�5�7ڣg_t�#�$d�Ǜ��z��h��n�i�omR��T��akЫb�/���p��vwVo��9�'l��A��kݻ�7/�o�&�R�.q�s�I-��2��e��F]wm����;�ZP�=���S�kF�ni�?Jy[UN�E
����YT+�Ed`���A}�4��^V:^%����OzC��>��I�f��:\h��.[�kw�N�L ��͠��8�̠���D�7��/S�kJr0��w55�\��w~�dD��;$��(����h��b��'`%�U|�j�j����e�v${�����0"�7m����q����V��{�5�-ð�ۄ��d�-nQ�|&ĳ�<i�nlgN�'.5���:&���z-ɸ7
u�M"��˛y�y���p�����\����;-gk���	ܭ�r�>V;��=,��J�%�e�pp�n���mN2���qri�s9�=;�(8ϗ�b�9��B�zѐ�98n�k�����sj��X��^6�=���s��ƅ�o�_'��|۵;è�фs�M�8M�a�[��˶y���k��W��-c�����Ń�ȯ[sҨ�w��א�?���1��ˍ�宮�Eؗ���Qә!sPN�tF;Y�N{���:��&��ǭƶ7]�y��60'����a��8���7T�j�Ԙ������.,��Ğm�^�]��6���%�l��"Z�)�kZ�9F�w��twg�c���kG��g��ܧDНm�{*'.8������VKx n)'v8���魻hn��m�%*�w���X��2�re���s_�ￋ�ϼaޕ����
�}��9��E�-�j�L������^�"pY��( e���$lY����=͝���H;ѱ�:Y�_1����w�;5]�J�t���:V�h��1\�-!�Y�p��fz������z��U���Q'+w�Q�����h�������va��ZqGn݊��ii��n���c���5�N֝����{[�s7�A�זy1)u�5��u����
�nS~��#^ﯣs����P>d
�N�S�Y��1�NP�n�=���2��d;�l�A{�
�
��f�:=�!81mGT��E�[�`�'����-��WΧ��q�b`��0o޵¤h�	%�~��xri��v�76����
 ��X��֍9�A��YE�ڍJ�_U�M+� �l��U�M�ut!�ԯ	��v1�a�%FZ11�Qҩ�f�\��߹�fw��ш�B�-�W��t�����d�1�~�v�d8T�~�r��)՗��^!V?�Hڌ��#b�:]X��`�&��*��:�*��]��q�S�nl�Q|�yټ�c8��w����˸2���l�o�s�$�E ��ή��$c�+n,���]�g۾�~��Ğn�����6��W���w�Cv4��jPP�)Fx9�����4��]s���~cL
$�1��45�:������ ��d�Ap}�! ���޳��:g��>A02���,1�Vd�S2���
`;�	��s-ק%�^�r3Lz5T���m��}�q��_m���	nA���u�d4�I�m��n��h����P~�<��M^�<;��y2YL���<�VU���M���]��p�8e[)VsDeryW���v�zT�kira��q6�6�$�u3��n�u)):� �=�H� �:C�+�������8�K�)�ԙ���CWFz�7'	gs\4��R-���1�[n�zmv��:��t��D��V7=k=h�8�c/�^�1n�D�n�sf.s���o���[R6(�Ыe_L�p1}�
�W\4�]Q��fS$�$4o��,�{�s�?A�J�I.�d\R�uV����LBoÖQ;<�S�Ŭ�$a���Rn�wCm���J��ܞ֓���Ŝ�a���B�f�jd"�}���o�[ȎH�K�8G2-�r,,ra���y�5��뷝�y�*t1�iK��VHn���BU�T�*�a�����[Ś���9�*GmL�3~�&	�������̱�� ����,ֻ��/S��������铈9[X�n�9->���좔XsT[����b�vU�$s�6�h9L?�tu�ѝ]6k�9nwl�s���>z�k�]>Dr�Lu�E=�YF���ۇE�M�;��{����r�V�y���.����myַi�O�;x��q�ù����F������\�N6�\�5�\��܇7��t�H���8���<��9G��Ϛ�������5D�W2sv|uﾃ���Ü�OV�pa�Z���d��q���ٹ��"��K!b���hO�ZΚ���dE��u��pL����̴�R����Ict�"t�7fޟf�lU���&�C's#��["���ф`�FJ3��E3}��i�y����4r�)qj�!&�mStq�[��&��ؑW<(�b�����x����s�c�sM���ö́��h�-�m0���T�G��7��fZ�����x�=˼@��a���(�*�8�� �9�}��W�lM)����wKy���p6�n�YMM���6�g;��	h'�[[����ZHYSV�;RIW0�Y��\�up�J�n���?�5��,h�Ve����Uw[G
������E�ƺ}0h#�#'�������KN��S��b���*T�7Y�s�;]���[�I�꾗��Ц��A�7b3W4/&��$@�����:A��SV�nŜ)�L$�o���Г��x"y �
�E��p$s6|�nI܆$�����ؽ%�ZW�2=�JȂ28��K�#�T��FճS�߸�d�=��Tv�7���h��v�u�k3o���ø���w-D������5��G�0=ڣ���J]��f�7�9ۗx��n,�kc�Y�ȰԹY^;�����71���t�Vp�;Ia�B��a��7��6u��^m�s�$�Z]y��9M�f;D�dН���Aژ�`�8��u����gWTQKNx�aH��b���8�72'+s����1m+7�P���ʡn����F������ɣ4 �@��]H�9�V���O$0U+Y��JP$Z��cіV�Y
2��ө�N(=��|�̻6���˻L0�`�IWɺh2d�˄�n�|��B��5���d��u#�o�n�×`{j�o���H�a�L�Y�w-Z�LA3��F���P[���KKt� �9�kY�B�Nn�e��b�f�xy�zڤ�XN����3S4�n�P�C�sZ�[TWy5q:��Wާ#������x����,ʃl�r\K��-�#e�}�ǵ�M�c3��������x�>�}���vSyy�*���{��i7�T��"�Hj�<�c	��;��"���;A;�}T�f�ܞܔDq:p��v�ɝ�'�S_ǰ����.����ψ�t�Us�Q+�\��d��mwmae��L�h��U����H�������=u�`;p�ʐoX�0[��9�Ys%˨O9.=G�Rr�����n,7<�m�0�+ԁh-<d�
qõn�س�� ��۲Z���L���������c.x�����Te�ż��i![y�4��rUHRE��kP�Fn��x6����
.��QGt��6	A���n�,�m�����bb��*�6�S^ԸU��i n�=�U�JR��rJ�y�y9�.�����R���ske�K�y�&,���R�h�ܳ/�][1��]�{�ڦ���-���&�/{2�eȍ��L+�%<z@�[��4�����[uH�s���s����#>c�K�1�L����/E�:v�\�6��L�H�A���\ј�u������_,�p}m.�ε�w�kk���ys���*\p� ��]H%�Ȅ��?W���)����e�&��Y�O�;Gt�K
�����E��z�T�q��ǢR5j�X��Z۸�M�;n8�h��c�9Z��]ø<�r�x��+ubGX.���q�v���ڢ�.[�a�zI�X������sb�v(��&.ܙ��+�Q4�qM�6�%M8�=p�}�KT<�N�Ւ4mh��$S�D�'>�4D����r8f�bO�����Z�)ZT2�����s˦��wJ7����@�p��i�[]R�)"��mjYnZY��̱��<��ֆ��f
�7|R�싦�Tiz<g0U#���6�k��u.�3UՁ��p�������ƣe�QT����q�:�K���S�n�K#5�{X��a��'n[���XD�?�H�4�L��V�9`��n��qb�f��a�١R�����Q� 2M�æ,iûY�5���$� ͹���J��������7Ç�:傢e�Hi�̙j�^�i�����˻�
�K�YF���������Ʊ+�'H�{E!T%޲M�X+E'T�,F�]���{Y��O׾�����m�p�C�.5b�^�K��9�û�0}�����,s�@�Zw{���6�m��LSN�fA�ot�Ki/�Y��P�N�c6�n]uE�^���De�p3��UU����|���d��]&o�Ư��l�,̸�$���Ğ�n��l$Kӄ��ʰC6;a���ckk���̢`�(�ٽ�Q�8���	B�Jib�
+l����]��m�.���!}��m��ʅO��2��m���)U*�(2J����lW\��a�Y�rK3�X}9�3�=��C�e�X����������sݫ��N' ����a��y1u���y5��n�z~���Ș��a����wee���d��e��$�c��u]%9����Y�䩟v袦�.�/���B���o�W	�jة$
b��y�b�[��s+�q�T `[�6�9*.�Q�Zػvn1M՜f�S��݋e�$R-]���	�����+�Y�ʡm:�9,�أ�{�iTZ.�cMȣp�\4[~�}��I#!���r]�;��S�,�����f��S��2@�*���oQW��;��!��N�oJ�x�k�VM��	5����%����q�ፉf��u������9myR�*��&v�Դ*���1�N��\�q�1�\�S9T�E"�I�u%�lGM@$I��^+�V���AЅ�D�Y�d�ŭj݌U�L��1��V|]�r)�L���MQ�9׀ѣ�7y��J�ƬIZ��f�br�(�B��\wU-`��R|�Z흕g*�IKf�B1{��1�LVvL�8��;E�g�M����
�3C�?��g��\����ܟs���ʡ�����l��B�ZK�=��m��d[���gq�בj�h��Ď�E��eE�����e<�l�|2��6��vp�{��\�t���8v��UZ�`�Y��U6hn��_-��Գre�r�n	�s{����Ή�M}}��LɥT��6�:�7-����E7
���7�.�ӭ�f7}] ^K�WWeFv�U�<套]�`�鹛'�(�w���V���{�5�b�g/ݘK���� ���B�*��s���$l�o_�
�y`�m"���-���㢚Ր̬L���_JF��0S.��h����VQjh��Yj�%Z���URX�*�T)fF���8UGUƅj���Y��J�8)�6(&�7OH�-s��v�T�CCMUJ����UT�J��WUUL>w���ŻD�-Q���
�<�s���d�:��lk՜��UH-	�95�R�,D潓��T@,�XF���?әݮ�º��Tہ�vۉrJtm���6��[S.�.��e	��@��,3�P�n�rf�8��ŀ}��1�]�e���:m��V�1,���vP9CPԓ[K�Mاf^��ێ����m���k�����\�<�١���y�;\M礽09[���m��=�����m��ꭤ�m�lklq6�9�l`����+��{='ͮ(b0�e�b"4��Nn��^���i���[u��]�<�i�䕻nu�iۙ�P���p¦��'_!J�u�Tf-����`�r=t�M�&5F6�1�)�Zvp��.~_>[ �n�ψ�퇵5HL��aąJ��l�z���cc��4�/Z�wPr2�A��wU7VWd,�.w����ԛn��F&s�L�&�Ѷ��ɱ�ݼ�n�uA5]<y��㭸+�3�mFE�n�Ǣn� ���*��(�[7Ov4��8m���J�}5�E�{*/�)�u}<FM���uR��n^�]5B�46.,{�{+f�&�^���v]��ĭ�> n�'{�q��$�u���£"�j_y��tuc����'s vg����c2��3t�T[�b�܊��MSh�Ok'u��V�9yK���L��K���.�Ҁ��& ?�zs�~����^@�Ow�A4._��D34]�#nV���$���މ���b���GZ{4�wuή�F�
<�i�Y���,U��By�����S��6\K��c�yc��b���Be�˻��[��c��ts�v�����&�Y�?%����1D;��Q������]78�:��STԈ�n;��V�YT��U&�.�:�"�v�mǫo>�r���Ȃ�t�]UH�{?���''n;h�R.�F��2\�}α�L���-�M�t����Rl�[�lmj��{6��g[f��ㇷKrx�z�F4e�TtO9|pc^��m�[�|{���G��G�X�w���� �}��f�U@?^�\雚��N�(ԧBcw_#�}�xEO-v�`��;�[�BOo4��&�y�v]� % ��Jxfa����f�qf�*��Ӱ)i�qJ�T�ؘM���O�����%v��nl����e8O.����B-�9亓/�m����\�r[ʠ��z�Y]ͼ�r9:o1;�j��2�n�S�t�M�� �W�I��r���v�ב�2BY�����d
�	kiӱ�؁�L,OMZ�8���Zg��H9���3B`2�@�����x�=�V�h�h���իpsj���&]	���K�q88Z�KI�Z�4�(� �Xob�,�c�ks��䎌Zol��U��J�]���9hnMN�ڨo!��f�p\-w����۵h��3s�nhKɒT��e�����.�j���RQ��V��ay[=]UOn��ͧha��;�^����W�tn��96��FW;kmO'&,p�#�yq�OTH{����FH6Drޕ�^����l�#�n��-�s�9��/p����P'��T����5El��[��p�10���:�C�w/}ݽ�j&\���\�^$,i�0����]�p!vM�iE� ��`���:���N	�c^,TH��fqh;�z��i�����z��aI@�T�ӽ�*x�ˏ}���I�v�u�k��w��X� ���4A�����XN|�﷮�k���1c��33ዑ��-P�,+���w��9��ιOGu�1�����.�X�PF��ؔk5D�O���YUNݜ�ê֥ٺ�m�Ʊ�]�;��r�ִL	��t@�%�ު��*�2n7;�x�_b�rc����D�Y�m�VU�;�ӳ4N6D$�!�;^�x�m�l�MԀԂ�Ov����mӍ�\�����-D�:�h���nL`�ufW%\�

�_`�y�rx���7['���ۛCw�6Lr�6����S��p'�Hp	�$��R�	oVɬ}���2/�{�ګ�=�#yS��D����% �XF돼-]9�5V6��Ob��q�����8�y�qɉ2f���ʐ�r��z5�t����E�C�b�(�d5���q`X�l�a"�Z0q����B��Ҥ��	�|��vb]G��fh'l?J�e�{��]�6���ݦ�:�,d#�\����s/�Nͺ�SDH��e&Cj�v���\��R��B�n��J:]�]��X���"GQ؜rpٵ:���Mq�mO9.85��i���V7X��I����):6�W���󣱰�=t�53llڸ����Ԝe���A(!�
��u�7@���G%[��7��j�9�]��u��^�8�m�O�A�@�C	���n�,4��pd�ӹ���;F��[�Ïs�}�Օ^E���%:�jzҰp��5=0g`��H#y���;��͓:��;i�!����:����LڪT8�(@�d��Wݿ,5�|+a[P�R��W%/��V��(�I�}����^�z_U��%MwM�df�#����7�)x��P�Wkj����;z���F��D���IDŲ�d��}�&��t�0�k2�kէP3����0��e%�փ�ӄcql(��%!��}�f��������l�B ���7�=zxxEn�"�I��`�Q8�'b�1B� R�9�Cz�&�bϐ6M<�.�Ff�ԫ9j��`[;1nk};<��i��lq��pa%�&6����8��&r��l��4{ �G?ϝ|���|ד��Lq�Z|�Þ뭸�&3��옭�x�;�L�n�!vB5˕�-�֮�ŋ��\���[rh�u��ϯ�gN{f��EkE%�yS��D�5�["������,[�+C����L�m�V	C�V��0-���x��,u*z��6ۄn�V�9x!(W�S\�i�b��#qK@�^ݔ�%cv��(�%�|�v�a8	5��6VcvEn�q��&�ڱ9j%���}W��s���x��d�X4�U�V%��3�T%���(�4�]��3r��� �m�cS��]�&W�7M�&Z	]����9'V�� �DbΪ3P��Ĵ���$�SG ��mj���Ŋ��%���"Oq��#��x���ޜW�����	˞��N�$/WЊ�R�G7eB���׹���Yqe$��vA�F���$j}�f�D�Zƚ��BU�-*���f��o�!r�d�+y{7�K[I��/�t��7B������)���Y��]��)��/G��sU���q|Bd8pKKn�.Uu譎�R�0�
32�����U���4��!o��a`�[�!"�o�z��׷�
��M�q�'�,�H�	�{� ����;g�۾�����j��r��=-�).[�Ƭ�d�I�gqΏ{�KrF�Iڐ1�܀1�b��q�+@����|�},�g��4��ⶋ{��;�-��>�9��nU�h����<��Q��X&����u-�ðC��B�w{oz�i9��AϚ�uU�&�*��(zo�V��ї|`r`¥���euWJ�}�l����9=�U���d箽�ϰ�Z�m�����[�9~V:C=��?$e�a|�����!s��U��ŀ2%MV��۩"���r�h�4�v4+�B�+b�W8�ͫР8P�sQ:.�&�P��X��"F�WWo�wZF�k��/d������5�B]xNP�>��5�N��l��uF�b�s��j�힒�V�
�B���z�E ���]��!����Q�� M��԰�I!�7���S�%EQ��1��&�����nN�s��yv��[c�%\GTl��Zl#����x�D����+L6�R}"�M��/a�߻���{q"d�T��f�"#t"FOQNٳ1�qǁ���jky&�R��O�e����UUK>��:X��k������i�烪��ЗD�]zop�$Km�^�]\���� ,	1q�sI��q$�#�K7'K$����G+� ���Cn~P�=L�,�lܳW�_*}�|�v���P1�v������rf�c�*�)%���$�U&�t�3�ݓ�nh�	�� b�ڈ����)�-���p6����s�j`�����e��<�:�%dqڹYysr�J����wu�-:�#��;7s;�A\2��%�vA�D�UvZ���m7�X��E|N�5q����Q�u�a��g��+ǫ�SBd!�iY"�E�3�S{�*8��܂y��G\n�V֋p4�	�U���0��M��!���\�;��G�ܜ�s�p�v���Jh�UQ����!BLF�����̛�@�a��OSѫ�!|�{�׌��rQ�㱬��fmn:�.'��$�:�NEj��=�|���$'�KRhT�����5\�e��z���a{{�#�`���-}[�l4���M= �Ց`��p3�C�����0�[�!n%�x`�-ӿV�D�c��o�y�=��(���6�vcے�'4�{�A����7�}�˗��Pi�,;�6�z�Ģ�1*�uږ���=��-Y���kL%w�oi]�EuE�e���FiYEnۚ�粞�N竝�=N�E�8Ɏ�v����t��v�tz�n����oL[�{\�m-��2ttXm�mn)pXd�6�D�V7���c��<�ܦ���:����~c���p�`�f$�u����	�,i:tlW��Z�R��tS_=���<s��P ���|z�}_�ѠeV�,������܊�M����s��N�wC�Ǽسz�E�н����������m�3$�w��q;)YK`�,A
����e��w���������Eު�Gݟf��*f���X0cC�����u�cԪN'3�1�����rt�e�=��լ�>~��ɞ˸'������بRQ�]Q�F��;<��Vv�:4�/�{loI�U�#{�u{��t��	��kEOU](��S\��'%��+b�L@�7����ȱS��h��9w��p���Z�k����AĜ����P����k�BU!!�T�qx�J/z���A1���}M��Ug�¬oh�`�Z�Q�I�cq�w�u�{�ْ^
��YDk��dWU��w�/7 `226����On��laa��:�_���k(�&f�[@Z����v/{��㫙�%Z��^�P�2��(�[�-]��f0����ު�;b��;{�+�:�]����31B^���.9��3[�,��z���*:�XY�����c�9������v3֘bS:w���ۉWr�ۓ���+8��ܺ}�)��5���Q�F�m`��`��CL+.fn^�s�O�{6e���'�/�M�gs�7�fÂ����/o';�]Ě�2����mg��� �OSHj�K��h]�6�k
��vQ�ۺ�U�T/yK��h�\�N�WQ���{8m�Ƹ�gRK,hr�aJ��W]N��
v�"eZ�
b�E�M'mݻY��n�pe�*9�/��J��q�K���70�u��}�pU=�C��u�b�P#:�ܼ�;���{8"9�����X�ٳ�N;'g���m�t�t����nx8�]t�6n��v������g���f�<�-��J�O7k\j^;{&_d�o6�u���N;�{v7���`�;������Ί3��-������۝��{l�.��7<��X3��ͱ�G���Ln�h�&-[V���\F�&SIh�f^&8���qc���p�Ԯ�v�m�8��]c��X1�h'F𲣞��$�5l]�.��瓷n�L��<a3�.�Mnݐ���W�+ڗR��n�h�ѵ�\Gv����\�c�y�i�����Ol���5Χ�vq��!�c;�l����;��ŧ��\��ڴv֮���pu��s�d$⤠��Z5�v�j�S��a_n���7=�v5`�3����mp�:.]��t��͎N]q��9DzWJ-���;��T!aK�|*�r��h�?{�^B̓y�M��-8���T��!��7ؤ�=�6����?�q��~t���x�&e�M������8�]$��/�-��&�D��3Ġn�ғ�����b�Be��Q���[Z��NV}��5��N�OS=�L;��	��^�h�y�8!t���l���؟n6};i둪�3�x{�,�ĸ�F���G��p�d�ev�|�ك5ʲp,����6N>X��M�$�2����G؛�#
� N�ܢWtl�����1.�FS�ҫ�� uJ]�2q𦶬U(E�]mw޷��5ܕp$o�t�*��Mtx��Gj���	�h��\]Q�P�?��&t�Q�L:G��k���Mv���~O�M�UB�a����\`%��0�;=|��:��u����T��,���XF����+���e�b��W/8P�F��Ln-�.�/a�����6.J�K5i�q׭
*K ���;�dĽ�ИE��D����Ց�n�?Q�Z�O�F���3��k6�F�lfx[W�����R��#���v���n��pV���*��4a�L�C}"=��!�U
��qǣ�н����u���G�*h�9vI���1����>۾�y��@����z�l�g���Ȗȶ��0���W�%�L�&.�'�m�{��KT�A%��I���D]�{r�b�ѭ�.�(Ճ

J$��D8Z���vU3^^��a��8�����-��D�q#��\k��� ���̿�5+R]�d�����=�[�c���A9�`��ݡ}{�k;��9C!
�z��\�*��9�/,��
^��!�GB�d��]VeV���S������]ַ2�����U[UP]J��۞g�eՇ��SF���Cs<.�Px;<���u���b��Ͱ������ve�p�L+r���E'9�f;k���]�n9��zݩ�6n�B(ʛPU9a/�R"�i�oٽ��pH��WOr
��+P�f�dR�;��O'wCڙ($�f�IY2� B�l�7�0/�nM�8��y�Qof�ռ1�rs���{�������\UC�3˫�Pe�����A�]#;T�X�� Z�p�ǖ�֎��B��lp��gn둄c��VA�R��~����r�ݶ��.!��a�e����cRP�5[�IS�N����.<ۛi]L�y�1&�)}`sz�!)('Xv�,	.�ى9���n+��b��F������)',e��e	����	T�Tg�ed�-H��x{-�	�n]Κ6Ǆ�3Ɍ�UE;O)�{�8�I�F�U3��TdwtL9��C��xN�ˎ ��\����H8`^k�VW:��v�X<�]#���i�eQ�9�A��Mo��!��n��d.��W�r��ݍ��rv.�H�<�Mna�<ݶ��Zy�b���o��ѮeY�w�|���q4[b4�dr�K�����x����^u��m��aݷ��<��>�pQ�7�݄yz��,16���8�HCNaQ�.
�TU�g��x�h��qq���y�4��x�a֊'��=pJ59�T�%P��Qv�F�TS;��FF�p%�����ң�GB��Ի�)�D��+͵��o���]���n����K��]^e�rLzo�ٶ������Z���/��IX�dm<��h��E��So)��1j`PmPF�(��8��(QA���{F�6��8�Gix�kD��)������k=%3��n�Ι�j�Vܗ� O�����u���]�W�����^�;�W�5�I�����F�B�Q	q�Q>�����Bn�z-��;�!�֣հ��4�k(k�zGs֮��i���Ġ�1�B��Ƨz�^Սn�y�����U!K8�w{�J������*|k)
����P�#�:�X	b�}�Y�V=|֊�Ƹ���X����yM�,��c�Wڶ���t0gִp��)�j�[x�U��"m[�m��7l1q�[������jN�$��P�p���T��$aWS"��L眝R��̼�ɨ@�	����4�7�mF_��+1���3�D�0Z���r�I
Hн�𭡔�����Y�Q{ ��tݾ2�hB�#9P�J� ��L6��i%0����X�����-�%�n746��욺ܫ][2�\�D�\`�o{�����i��� �t��s�K�[�G�x�,s���P4E���Wz08���
<�Y"�C������1(YW(����/�-�ü�[�X{�v�J/V�z�r;��R�C�{$���Ck��̩y/u���v�so�7<>v��^���`�#����Wuܻ�4'1�㼓���M �]i``Af!!F�o����s[�<W*�#	v������@��[h��w�;�V�]h����`_+C0��Or5�S��OZ�ڹ�oD�`�y�llfP�k��z-���ԫ��[I�jŔa)x��n�e	A��S��m-f���[ݘ:3T�T`���r�z�!Df���v8����,~s}w�۽��6����rj�qY����H8|4&N�rހU��l�&6i�A������wS����r96'D���M���T[�Ѩ�|���夏#�01 X��Gq�����؎3�!"�*Po��'At�<���g���͒�a��<����پ��v�y�B�6�M#���C���0����9kn�19���nF5ZX��=(p�F��r�m��8X��cmA�3{�����5c 
�S��X�b�-��Đ{�g�nwI7�`y�z��R���L��ϯe/�7��cKs�B�G�>����
؀*7[r(Q�HW�*2I5��0�ƅ�^B�&�H[��7L:U2)��E�`�cs,Z�Q`E����[��ڝPPW�W*�N�J�y۱�CU�q��wW^f��y9�niRA�L�j K&�V�U�ॹ��p�WX���4�83Æ.�:�Ż!��b�Z�Oc�Y��;��x��]˒	���7T��ۏA�0e�m,m�SPں
	����vd-亼���27s&F9���NY�Ը����p#Ek��(B@�Y�V�H��㙮��"�Y#�҇W� l/
�w��f�
f;�h�j*�֝�%κ"���&�p�zڔ�q�\�E%Q�����C3F*�h��+�Z(�Yk0U��	Sn���Հ�z;,أ�0FQ�܎���7�R�҆d������&��\U^T�de�.���������x��3ȲY��tq�Dv��ݯmJ�M<�����5L�"�����RP;`ƎV��j�~́�\ʄ��e�SZ;u׽�O�Qs�%�9o�G�\��m���ʮ���U��
�!� sZ�Av�K���\�6���i�������$�p��rbC������s�V��4Ҽ���+<,RkWM�!��	��b�$#zy��ꮁ�.��$vP�����!�ژ�B�-<�OG����8��KZ�����z�D+�o\kJ�+P'Wi�T���VT6�����{��i�j���8���m���7���d�wO��7o;��%P�"�sj�;vz{�Xv�,��{[eқ�����k��D��4�˵sZ�ד�i��\��v�s�qc�!�eH]�����3/,�ɒ�w����8�����<#AZ����TUx:Z9N��}����<ND�i���ĎΔM��~�l�]>�P-�����jZ*��p�8R�Հ�����l�e�9|g�_[�����<��ʩ�/���������X�C��H�#n3����y��qz���c@���ȱ&2�ޙP�X�`<'p�+7m�^j��������#��:�Ϡ�r89n^�&����7s�����8��z���"iG������F��C�8`�%�nA��f)u���L���������xÁC���	X7SPv�Ϋ9j�t5؇���yhUuu�A��n�b����B	��0Qۼ�i6	[��r��JYbR�*^��`�[�1<�ڋ�\iJ���u��v9�]O�������\�	��K��Tj1��`�(
�f(<Wr�ol�%+d/x+�|�2�+��i�7u��Ά�ۺ�Ю��j�"c���˭.�Y�{���V﷏:9�'0uz\M��0�`�S1�m�j�h�����E�V�NĀ��f��K�\ݧ�ħ^ۂ.2`����;�M�6���R�Q�?N���K���j����(D��n��p�
K~Y	��;`T�(�p�\s��Ǿ)8T�%�a�b�b�4��W��1���iK�M��&U_2�o��������S�d�1��#c��'\�wB(@�Üu�S4Є�F(<0�e�l�[��/AB�d�.�����lYX1�`�ˌ%� f0S1B�މ2k�O)b��a�]6x`�Xֆ�����'�r+8���Y�U&xZ�df⫪ZO�@ɗڕ�Y8:��d�_=g.�2��w���ޜ�������O�ݠ>f���i;Ȟɦ���[�i"���ZŚh(��� �c.7\k��n�v�A��{���]ϜHp*�١�GЙ����H�\�᛬<n��3�9ۈ���5��Vyvݟ�>I�V�,a�V��0_Z\�`B��P.�
�@lb�8�G�2��������c�ڕ�C����8�巏��Nr�F0D5Wq��2�_���3��;��3�Ԍi�x�֬�kΧ�5��,���Au!&AZ�ԯ�oָ�@[���9���ζXB���c�	�h�qc��$`�U�W\Խ�A͎��`��.xJ�0 �$t�8��h8an�����-7��������T���i��"F��T���*�A���N4;-=����L���54�F�7� �H���������HS-nu���\�y|�N�VL��K���&I2U�&c2)�{Wf|:sp�/�g���څ2�Jq}���{�έ�o������v;�v�~fl�x��)q�Ӝ9m���lr�=]T>v
�sz�� �n,J��u$ ���u�{���.��2�^����(������ ���UAEU�!UUTW�䢊�(��5EP��U�PQZ((*ڢ������*�����
*��μP ���� �PQ@�������((� ��ƿ�����g����UE UQ@W��P (

����� ��_W��PQ@���O��>��PQ@��Z((� �PQ@��P s��tPQ@��.�λ��eP ��� �_��k���� �

( >�O�������wE i�6���n�P D�PQ@������d�MeeA�dх~�A@���@ ܟ}���7���P[ �}�mmA@�k[)Fĝ�     �M�N�P�@�N0�h	!�n��c0ww  �"�H   (     (       �      J�� (� $�  re (P  �(hQǠg`�c  ����0�t)݀�@�9R�U6(>��    b  (�  �*� }�޻�m��\�]i� �p��z����.�!�#N�q��� <>�   

�B��4�ӣ'@U1UӉ��\�F���q5Qn�.���p��j*�ԌVXQcΗ��K˻k;���} �}�}F񃮸����Az��;Z��H�\�է��&�q���P�   


�T������"Ҍ[�7�Tw�"��C��1�`,�F�M7;����Z�.{����)ꇹ�֭��:��ɋ��p�{׵��V��^x�ښ�]ޭR���     B�� B>�ڶ���ڵ���T��]U�pԖ���x�u%�gM]:�n6�۞��wm7,
���>��y�֣W.����@*Fz�m\��\m̭q����M8�G����{u�կ{��kW��UN.�S���    �	P)�mj�j꫖WF�q+���F�W��j۞�T8��k{�%#��[c��8�黸���lܹ�j� yH����7tZی�VZ���T�{�%C���9�zy�<v�;��Ŕ�� S�%6ʩT� h T� JU!�  S�j�U i��F AتRE&T�h�l��  h M"I��	�40b~$=:}�̟��?��}�o��;�{���Ͽ�! � �$		i�� � �� � ��! � ������������✩�@����	Md�pM�*��V&%��)�8v���H�Ν�������}>�����a%�o���/��vh26��*4\�.�w�a���]B�+Dƛ�۔(Wż�+�E�.5U�UT�U��DлީX��!U�!$�33����Tu�l豅YU!�y���-��E�a�pˤ 5 U��%�� �X6�	L
D�?Z#�e#A^��(�B��T��vh�$�?�P.q�v�����Y��S�n�K�s0wf⠯�.�?%͛��Ⱥ��ޠ8q+�bvDt��A.ʹf�̧Pd���B{�|��ӔA��,�5h*�HҗL��#�������R(��m@�n�pWeۉ]��\�4E���?_۫����c���*�`�.�T(2PVS��$�w!��7U_QTٮ����5��l�����d���(UU��d'P�T�@�Iy��ʳ�8�Ul���n�y x�A�n�oWi��ۼC��c�V��Y�V�oN̰3_�2��U��B�N�Ӑ!vT�c��Ac��Q/�Xd���".�3YNZJ�vN�eU��@]�F����y�{����o�<n��b�kN?<(�'!�T��k�lVh�A�ޭ_]Um�ON�čX+�5]"T)\��-_�1nf� ���&e��w��Eʃ",�c� �C wjѼ,;��c$N��h:	\&����� A&�"J����+��:���mm��2�҉�T3�����Y����B���(5�`��m"��Q��4(C�f��K`ٌ$(c�K�w�4�0CxE��JQ,e��E0krƻ[�m����V�
�6*�ϯu�i�7�pe��j�X��ꪲ��"#���U������s2�&n�]�m;xr�(�7L��L
уU�N[�
�)LJ��T��aO6�q��R�F;9B���$"�4��-"I��≅/lJ�Y
����I&�)Q�0��T�+�V�9h����LHe]��f��2�&�;n]�j*�'��Kr�Q(E@�n]@+uR�%�ˡ�s
%��W��gN �7��*6z�kY�;A]cx[C��97�am���!�XB�Sj&�8a*�[˘(SjD a�j�����\�u�5�����՞�sh;G�6L��R� �s@%���^8sꈈ�L-��ׂ�Q���%��f��*SH�m�
$�,f�j����&�l��fɩr�0����ф^+���c�m����h�na��j%*����;vN!lvx����ژ��f�QV
q�f�B�2X6���/ν_c����nU�}�y��<�E���Qn�9�ÓhZ٠��G�q(���y{/H����;���sm��m�u�m��D��U	ᵱi��TAHZ{AV&eк�wxR� t�_Uo	����2)IQ(�[e�1����h�В{��4�&9�b%Q9tɽd[nVL�[vr�p����v�;��|�Lr��Q�d^�c�U��C)��,�h�ZZ�qE���.S钝�����H��1�D֨�m��4}Ьa��]3Z�!�U�ɷu�BU5Hq씣�p(�%d2�]�r�)�6��QB}Kf�X�X,.ł����ٴ\���=��6Kq�o�rg��7[�]�
`R(�d��&���(���VJ�gj�������/��P@#�0�$*�kT�cI��4IDx��*��7�n�u���KK$RjV����w������J̙��/c�^����}�,>1���a�E��H���t�F�c���&���`�w�F���S_�*P+wB�śP���Р���Q�@�T�M5N��b�-m�� �̊k�l۬���\������<aD�V2��U�U%h��t�e�6�`7p��q�7"�-AH���i���(��3!�_DD�ז�j��M��5�kwwx�h����N<L��<��;JUe�db��*]|~��-4�)R�U+_�řAb��ؠY���m���x,�+G�~2�A� ��)�n��3*�j�3��xb$1�0��p��Y���8�nӚ�\��-�]�ضQ�sS�L�Mv4�fiEi�<��_�������P���b��'�f�ɴ��j�D�#`�I/�)����4�B�N'��}d��Pd�D!RT��`�5-ӣPSA� S�>������oa3K�������PC��'ܹ�b�~?>�|��AQ��,�F�&ꐢ.��l
r�EM��y>��]�aʑkpY.����T����"�7�8�w����L��G�h�^:�{�W�rڕ��I�8a�X�X�����,g)ETH,ieUT���@V P`�j��EHH�,� ���*(T�����E-*�Z��*AH!%�(�*(����X(�PFj�kX
AHZP*��"�,�l��Zж�T����Q�cm-�e��2,b��lbZ��F#�FB�X"[QUQ�P�X�+JTR
Q�(0R)ETRTm �-�TTU��� �� ��R�B�
�+"�*,��UaUF2(�`��KB��V  �"%@�"�*�J�
�RVT�K%R+%�X����� ��A"���aPZ�m��D�%��PX,�AAeY+b���J4DF�PkiAka[h%��kd�J%H) �,"�H#"� ����!m
�d�m��*�TX��Em�
��`�d���E��BXHTYT EB���
��jV#h�UIm�($
�U�2J��P�T�`,��#U�P��YRT� ���R
�H-d
�*�j�
��HT����Q
�HT��R!XB��
AH) �*B�*B���ih�J��,� RE �,�AH�H) ���R�
AH)
�� �����R
AH) �!$0jڊ�͹ � �C��<����ن� �
(�����ő֪�������ERq������.郈�1��r���&L]<�F�a��n�U�������5R�nB�!DJ-��
Z���ppGF�Շk0��ڍ�-_g�B=�k��~���T+ꌄBa'fEY$�$$B%����v=���|Y��[��v7�_@��P�80!���ǘ���(ρ�L�
܇r�X�آ)r���Ǜȼ��T̅�,PM)�X&u�lj1��L�X����|i�XÔmmA���+�g�/;�|i�1ڙ����ZT��t�ɀ�wtɉ�mÌ1m�L�k�U�$4�!��l2����uŻ��;��7��¼�����H�,HIlY�t��Ib��U/����tݼ��]��7#�ࢊ��`VJ.�&]7\mV	]p�(���vp坟]}�#����D��%�N����g/)Ki\�"b�.�	��`�Y�X廆�*�(,",kU��2ZWZ9KR"��VU� ����%0�q|�4��룻��71<m�B�#��XeYb�j��PV�
B�*Q%H,���a���TW-1R�����4wo7ͩ���bs��t`��G"Q�'jq���_������8ʻ���2��n8y�d���׉��eo�y"�ݹ��L񱒸���x�s�n:�L��V�Z�B����AHT���`*�T���H) �Y��RE`1!��-n�c��p5&���H��)"0��C[�ى��E���a�1b�ej��\�
����Ȥ*B�D-�0R㎥.fj��)h*(bYKV�.���R�7.�LjU�s"��,�m�q�� �=>��L�1%d"���i�2��� qJ2�*"�'�)r̆Z"�Yb�[��1�\h)rౘ��̕l��pR0��-�W��<^n��F0Pv�.7eC-��\���w̜�(��0��W"��Ai��)S�뽇Z�D��.\���	�o�������J�
&LZ[��\8ˮ��9ŧ}�;�B:��v��m���!r��hؑ�Ww30�7��獓{}�o���܂�;�'A�ڣ�yY����
�u��Z���
J�n�����)D#�]K��GB�9��P8+e�+��� �oT�e�&�e�)Р��F[���?Tm6��QX�1�fV-��w�j��5�E��DyJr��o9K������p�PS4˂�V�-��_^V��EEA��g��{p��=��{z�7۫Oo�@��b�*��[j�P�nf	-�� ��-
aS�t(UB��R���Ǖ��h2�a1�1D�
3�
�u9tG��3��lP� ��x ��ˉ��Ŧ{O��E� �R"��LQ0�!90�2Ы�d���A.�N
�q�i4�v���Ef�i�qX��]V!Y{R�#�[����O�#�QZc_g�
[(���n0F+�e�l����r<!�yU@��5up��e潼��yKR�`�W���Mk�6\z�;��^eMԦx��O�ᆹ�;��)��m^��<��9��VᗉZ�\�g�w��eD�T�HrO�q���E�Tp��"m9�x^y��n�{wR�h����+�X�"���ł1��R�PR�B���J��V�E�Kq�wsZ�)�ܜט��͉]��v링��Y�N���QM�4-)T�F #.�Bێ�Tt*�³j�;�Щ*��IUA{A�d���J]УBE�
,A�rX%Y��ڨMb���5�[u�F��=xUIm:H�K�-�mMƫ-|�<�sL�Ng�ۢ��8�>Q���`�%`?�2������6��)�Lbѡ[)r�+x���B�1�՜��*�!_��
� ��	7y�YN�D�B�!�;�7)����.���Ub+��vl{������YN���w8��;n�1<ؼ��2y��3U�@ӧeJ�!,j�%�.��	��E %��ږP�"�iA���.���y���Ms0�Qq(�e`�6�qw��eM/&#r����#�4�و��(R��a��c�c�t��`��lc�r}�����n���s8EU@�V��7��DPB��e�)]u����(� E<�ƾ2�Hd���Wb���L|�r(��
( �C�w5PGJFDŷ�X�%���[�����ׂ���"�m祬h�����0���ph�`"Z՜�k�9��ܼ�r�����~~c����|��n�܋Hl�܂TR��-�˻0[���v4`�/ej�`��j�3�G�b�e��]�ˆ��jA"r� T8��ܺ�d���]�߲2�Ĳ�є��f�D4m*{?^U
�s�!՘3r����]c	޴X1v�h�p%�fű����=�G-i��6fQdUi&ꪦ������wOd����TRh[�#���S f����PlW؅��h�t��h���� �
,D,�v3-���t�Q񍘛M��k)>z�qv{�e,�)[Y$pQ��LV\��<nnЪQVNŰl�k��ܭ���)g�[!Z�i"����m��"���m-��R�������K���`�o�p@G	��'L)p<�Z{s�4��$�(96��&:6�<oAȦ8䘞����i!��B%��	���i���d��,����k�2Yb#(gg5F��	��D�Z��كh8��C X�wQ���d9�fV'*�\��Q��u�T��-8�ƺ���R`�\X��U�"�F���j�ݪ���P�n�P   p 
������   �
̡� ��C��� 75���5UJڨ��������n��N����@-U#��89�t�#�l�՞�M��b�fHrԦ�w�������-��� jM�ynqe ��*���  6�P�J�v�SŶ� ��   � �� ݶ�TaU�wf�%k���X*�v�Kʪp�   TQT       *�   T
�*�6���� +3( �]Ԫ���*T���Swl  �[!T T�7�+�W��d  �  P ;�w`*��� ��m��I��F�͵J���*]��RP�f7N-��n-��c����B��k���/��Ӄ7nzη�s��ڔ(�����ʮ���� *lT�8��UA� �*���r�y�y�=��-ÐA �&Jۍ]#�PAx�&�*�"�ɻmme�����\�0�0$:�t�=Y� 9]An��һ�"l�QY��C��K�����㱩�;�ҳY������v얣j�_E��Ҷ�P�4Gn��n8�����b�ԕ�9��Vg�Nڤ]�rl�=����]me=,������U�M��7�F㪚��^T��&K�a�H�{A̚��m�n�[.��-��U��+g���z�,x��)�u*h�n3���nx5f����+�9B�(��j''Wn�\ۣ.l�[�v� z�3���d���Vւ�ݓJM�����	P��mv��17,��&x�qі����\���C�d��`�t�p�5Φ�	N�3̊�7'i��!��`���T�:�g���Ix��LQ���6�y��Ѻ�)�C�xyG�PϞ�ϳ��q/���ƛ�e�\��;ܯJ�Wtۺ�(��d���9����d
�YGF)�m~~s��&K7I��"l��s�m��B�x����,��^۔@����y�]
����`�Z�Xkj~�}�G=��\�tŚ�@N�a�V�bؘ)5��*���ڐm�ٶ1�Me
(m���j�U"Ӷ �3�m��x��<�UVІv������:��gkG;�Dp�X�.�97щ����\)��8;�|���Y4��;�n�3�AÈP��q��A�`�P�G8q��6�ejy�v�;+����a��:�"���������6ɋ�4@8�+-����]�l�*ᝎ�@�7HB@�u���u;:xF{99Ӣ��j�k����Dd�ۮUf�
���`ܸ�뮭���][�p���PR�+��g�଻y�{&D΄�ѻ�-l`���Z5�g�mgPݲ����E{SU�c�8z�8Q۳tF�Ҝ2l ��7��'\��Kk%�y��2+��#Oo3&T�kewM���g5�x�� OG�K`�,������+�.�N�R#�Y�v�=�f�w;��t��rLy�6��b����.a�I�v�nY�bD��nq��e6�d�9;|�_�j���e��.F�C�˜KUm�60��4ţ�jKY�[��k���Jm�5�4*��Ǉr��,�hq*vi��.��1WMۉa�@MEu�p�廳�;�����`�B��Q�v�m��q|�m���y�݈��
�g:@�Y��s�n�	r9���&p;gL�:�IQ�H�M	�,ܗE�"i��^��Vm��Z�nt��r`K0Z8f+KT9 ����y�6��ù\���a��]����[��&mfv2��Xr*ڳ�V��╧d�R:ݪ7%�"��S�F.ַ[l�6�ƶS�DsJց�#�*G�Ƣ�+؅�S�=��Ӌ67���j�5��pm�w$k��G���}�;���s0ݔ�v�bVA[jϞRx���Lu��x5���;��c�N5�x�*K;�8N��)�.��n�n�gj���j��`���۬�M��c6���U4�k��$�����w)���͍�g��[�b���r�\����i���
Nn�cY�g;��H|<k�A��iM��#Pۈ�W���k�s��'-�����
�Ah���|%;Z� ^��7[8�m��m���ٕ0G[�y:�dX���{c����\��s+n5��-\.�"r�F�L�g��ˮ7K��ޙ^Ol�h�Q��\�ր5�x��jtr����6�`s�&zLq����vܐ`
��<N���a��[���mk�8�����<�f�.������kb\�����
8�n��&��2�+sG��k<�Z06r0��V�(�ll'�ә�b��.\�&zWu���-���Oa�g�6�"�cVf"6�.���o���Ëg�R�Ot8��Q��:&���`�oa�a�N�}����mRڣrn[k �lFȾK́�t.���S�����I��X��"u��LC�=����Sʪc�7[���,����$dІӣPۏZ�-�D9l*�@�f��>�v;8;k6�j7N�%��D���f�<�:|\󆭻V�&�-�F��ֵ���7����~V�Nͮj4��W8�v.�ri1DE�Cɇ�l�ey�sW{��k�J}S��k+�s���^PTi�#�v痑5��t�ρ��G-w1K��v΍�H��g�yvۆa��p�[�b'c%�Z䢭֮�a'�Lk�뎵��ïm`f��<�;�P�a�2��3����w�������o\�u����&q�N�Y�ܹ:';F�z�� �fcc"�ݸ��n�{E;��U���=�+�8v3��@��;jx����sC�<��{BC���q�gӞ�e�G��2�͞ �5��[n�F��h��4#��ș���O�۫����g5I���jG�_��mv>���q�d�;l��v�v�`a�P�D���S��D؊c�r�uݍO7��Uێz1��v�pwd9�;'a��7��Ę\�����m�aݬn���q�qHd�5g�^wdѨC��u�=�W4u�:;X.��7M��3��X�M�<�ƍo󐜑ɵ+��׶��+`�Y+�=����`z|r���",��v�������UѴ'f��� KȗiM�k
�h{���0�l6�p�n���cn��uu m�[�q۷[��xGl��m�uۻ�t�.�p#l�����^��F�v�d'v%�;�`��۳���ewi��u��FsR��pe]�+�r����<�e��^��zN��%���E���Ͷ�b�6Y	��c�i=�M��aI�
�q�l����vS��d�.��h��H�9�ݦy��/Fn�%;ˬ+ɳVЛc4ݫ����|�u��M�{*:��ss���s�)�lٻ��6z��m��Q�O.95�%��䱗S��3��Tv��*8�@�YFU�yAUZ�j6�^���-�z8
�m��d���U\s׽���f���w7Z�]�u����u@�    PU
�aY@   :��aN�/-��l@  N ��s��< <U�c *���� eER�UUlY@  ����J� ��k���6� ����۞i�݋m� ��Ҝ4G�+�bD��FV���]ou�Q�Jɽ���45H ���N��2�uS,r����<Þ�	�9�� U@UOAv�T)0;=�l�R�$q(ۀ�vږ Zx&��=�[�#)�JTY����� �       
��T��	UIk�(�ѤA]#3�S�U��U�ж�Ӏ1�p�� �p
 ���   ߷w�ߠ@    	��8@x x8  ' c ����` < < ������1�p�� �p0;�[+�;z����( �Wk�����`6���	�g(k��ݩ���#��r�̪�U�]����P�P��v�d��U<
]@gW���~��*�f��}�zn�-&�3�jz݋�c�j�֮���@��T�̨@O&�lױf�T @d   ++�lBh'ӓ*��pb^v��$���Sc[2l�  Sj�Sb����:s�����Uz��AY@ *�5��nkl  N5��ob�m�@ N �g�*�ֺ�k��s*��� T ��^�TJ����*�Z
�jUhSˍ��AT �{J ���;ݵ��iYnYN l    0 6������L�� �T � @���֚��;��/:8�#�jqJ5&m��̔Z�iI�@m��'n�9�]���r���"4k�哉��,�UC��� U� VS�xT��ݕ���J�y�����
�܏T��ms��1�l�ɔeU:f����                     �                                      �        P[ ۭ�  �m�� UU ��l��        �P�A����T         
�T  *��     �� �T       `              �v�  �                           wi��n���m(�E���������XI � �4� ���$�� ���=�҆]w7nmHN�Y�v*,�X�wb�\�c,%uKv�Cųv���L�0 ��n��������}�@/T*���"�^��*J�X��vu���v�� l�̫��P@ 
�檬���l�iX��
]�W�\�f�}�<��uU5;:"l�ݍ;�b�@�cu��\�b-Q����ySA2��۵,�8WB�tt[�ܽc�;��pG���n�S�T�\�����rOj���8qy����ͭ�{0�,��^Ec��&���8�����Ne�m�.����Nr���u�]��cxK6�%1��m�u1v�\�{[AۚȻD���q��I�w]���S�v�Y�܃b����m�dL�<���@�Bt�����Q��WTmn�G�[�֥�s�̒����,���.��w�q8u�.zqۉvѷ�<�����@;��B1mګ]���6�.өb��I�� �p�[�,f�gTct�Q�hY۲��a���tc:`��ð&��&�Ob�]�i`֗�m�5`�I�2�Z��6-���-h����$��upE�$��ɗz��`!:W��δf�z�����-N���a��]lgs�nR�c�u��g�;��,�n�S��g@������R�3��Ŕչ��6��v�lH�\#sz7X��n�ܧ[kcqs�Y��+�*��ڦxg����8z��2y���N�:���b�ӝc
��J��tW @��UR�@�wYG�� c*ʵ +m@*�n[k1v�������z��v]�Z�0 �M�ݝ����p0^�=����1�p�� �;��O '*��r�
���n������mR�Z������yF^�*�Բ�Pz�x�
�*�����zT��P*���fP  ]��玪�·ճ�ZT�����ۻ{7�`           *��� �   �  
���    8�   ������\��rׄ @�I���~&pF���1���0�aA�z�]���Uw3��.��i��0�M��M���̙N���*;d��9��=���k���&]�hym��*�p�x`��Rj��9k��[Z�Lnp������[u�u���!�n]��"���]�c�z*��Ī��n�㵬�u��x�m��e��N��: �6���c[�˵@ Ul UlT�{��G@;��{`�e��s�xϳ�8r��v݁n]�w�(�L'#�gc���}��k�Hg�q0t������E���"�k�k�J(k�\�0a3�n2Κ"�8殊���=1ej�ޤ����������0�%��#�HZ��?�����g!_oJ�-i�� ��5yA9��4^�.|��É�9����Ο���ب�e��	����8h�Τ_2�%6�Gt,�Z~:�����\�q�Nz`����/O?>��6`iD��.S����uΚt��(9.1���u��AUР72y�P�ft㍴v�xP���r���-� �3��H�g!voJe- m2PvaB;�i[�Dq����.����;�!kǼ��Α���=j��d�Fa�i�z���c���iA�p��H��5�Z�ӄY�������,�<Ő�5dgR��A0Ւጳq��a�@�r����jaB1��Z���p�v󎅘֑��%8��f���e6QzaB+��s���!kH[��a�(���TF�;f��h�X��L* ��
���ɛ�JEL FX�K�"g�;�lK��\���5�2��.a��Y��cXE/S:t�!sWE\E8B���KD�
蜬�$,_4?C�{8ɧ����a�\F�;�q�"�F5���,X���W�<��d��B:9��B�kH�h)<0�!�QsӦʋ�!�#�Q�D��"��Lkq�,6�IHT�֨�8v�0�B4�Š�:t�6Ђ�k��igN��'=r1�Y
2�Ø���\*�0�u�#g���4� L;K��g{��|���3��7Gc�l���h�e\�I��=s��˹�; �uH
����;V�K��2���o��q�k��f��0�z�/"�GvPJat���B:�#f�\�5�@�&I#a���Fr���Di�[tT��[�0��Dn�B
4�G	7�	�i���t�B/f�j��:p��.cGZ�7�Zx�g �=K��g��`�`�!E��%��H��n��da�Dn�>R��kH�iH<0�!�A��i�g_[l�Ԉ	�Ĝa�TB�����F�U�Di¶�)�2�3�çM�È�$[k=`�������q���lۦ+ nE�֦�Pg�c��4�)e[g6�Y�e�Q�B�5�Y��3�H�o5rU�Qӆr�qB:Ց�
��H�<��D��P�	g�Yl��QƷ�h1�0���1�#�� ��,�w)"�a������TV�gM��pCGZ�5��t�3�����#N{`�!��4�`cQ@��H�d���GM���(���#�t�B-�j��:p�Q.#GZ�5�.H�Ƥ,2���:E�4�iqlΆ���!��1�4F����u�k泷��@�-�*�Y!�=z�t�n�m�){�Z�Ye]��VP9�z�'�6$��c�C-նM����y���ni;m�fe���=/�۟�>���t�,��g�NƷM��xi8u�;v�e6�� Hk�<�9�u��0�vr\�������5/\�\\��Ul@ �n��[v�m��nx�<��
�հ�:e�$*�PQqb   :�  *j��'e�9�1�l�G��9�6��mv����qv�\?BOԶ5�as����X:¹#���#e�u�49�c&��R��֨��ɹ�"��*=j��hk��Jn3���Պ���;l��Q�V=ou�!�OE\E8B��"08��ʄa�VF�+O#CԸ�6c��H��a�{�c�ύd\Y���"K]t��m)$t,ƴ�4^����{���4�>i�&o&�t�39E�]nT&� �Y+�Z�뾾E��ִ�N�!n�Q����g����F&B�c����Obw=H:x2��h�㎹�z`���۳�`Y*C>0�j0�	Hۮ"��0���dw���4�D<x�4c�/�H��f�z
�l?�l��q�M�-�,��0�4�F�{��#N�1�DG��"lE��L1I��.�:E{�Tx�4ٛ�T��Z��N�!f�Q������΍A�Q��1�ּ��`Nqtᜢ\G��#x����a��i�=��"A�[f(�"�F5�_' ��#joF�Y�ih�i�d"�i�0�:l��%�H��Ŗ�$�В6W�.���\lt�����͝��X�m�m���B:Ց�ԋ�a�(���֨�8i֓0�B4�;�:t�#L�ѢAjC!Q�B�kH���Ӥa���5\E8a�W�#�Yĭ<t�>c��V�d��J�yӭy���+�H��lމ�8æ�Y[�JcZF/YE�Y�ݳh2B�A�Bm*�,�>a�VFoS.q�H�Ƶ�=j�ӅUi3d#zA���Yb����"��=�Wk���Ӥa���5\E8g(��#�Y;����#�&@�����'���&���.3��쵂u;skj�o��@�S��c0k�"���Di�U�_V�d#�7�pqgM�/��,ƴ�"���7"A�L�0PM����o��0�:l���B:Ց�x�8äQ���=j�Ӈ�.x���$e��Q�ZC!k���:h�3H�[XEԎ�#
-�kMWGN��Ѳ��d��IZ����^��<:F�d��VF�4����(�ط��c�ύ��ld��%nH�^uƴ�#]������QJat�Fo0��Q�D��"��<�-4�Q&�N��n��ֶ��<�!Ȕ��X1���/Vʀ�a�*���Z���j���4�Sm)�2�i�І:l�7~�[XEԎ�#
:��Z\M&�7	.@��"��3�K��do���0�+�Z�4٧�_V�E�u��Yġ2܎F�a�D)��:��0�z�/"�-���M��sc
:Ց�O[��m�[	�$eD]q�H�9r�֨�8c�3��i�ћ�wh����-�03 Q&�1�����jit��|F��doB��:E��`�yӭy���N��:�� ���A�m� \J���mR��l�b���܀������8�[E��e�N�&���W�κ�ݰs�ۙ�.�N;��v���n:�n˗,�����@c�ִpfs��ݹx��7KƬظ�s��B��ġ�q�N� �p����s��5l��ݑ"e�P����zk?7�տ`y�x< <���:�9:�@ilpSae�@   �Uq�D�f2 e.Q�ؽ�]�U|ujӲ��xz\�oX�X���6��ם@9��)4*��챗���<� �Κ"<�-г�0�ZO��MEf�o1\�RLd��-ŉk�ތ�y6v�]u�6���i�wBt鲲pX<�Z����E��a���t�B/g��8��9D��!j�ܬ�x��Y~d&2)]n)-,mם,�6T�'�H��f��a�Dk��%1�#ۉ$��,�vw~"�I8.	#j&��"Λ(�����Dou�t�<k[�֨�8UV��2������' V�Y^n��n\��#�W`ûT�q�u�=C��v.ָ�������ı��`B��E���֏{�U�a�Q�H��0�[�E)�qӆ�qB:�kk=�B�Fյ��I��۸����,�c[���t���K��a�h��� El�7`
y�0�S�E�#��1����df�i�0�a�*�Z�4��M��e�		�
4�i�i�ˁx�m��G5#�H��ԓS�����ٌ0�%Ȥ&&5���;+:�]w�沧��\�a..}�cm��E<L��mZ��e.7�#��6����[ʮ-��g�2���jn.dI��~[�M�yA�Y�~Ӧ�kx��#���{�s�:E��#"q��+�%�T<a�M�{faB0���t���
,���jGN�#a�� $F�m��������%ܖۛ8-���� $XE�
Bd�I"�F"��DYT()���R#QE�(�UT�2"(�U"�F"�dPQUAEUDX�(�H�F �b"łłŋ�*�U�VEDcEX(���
b���AAEU�)U�E�X�$�A��	$"�E )�"�H�"���B,�Y!(� �E�Dd(, �"�"�
��d�$���
,X��T�
*�
�"����`�������(��T�,AAbE@P@F,b��X�)DH�*����EX�*1R()b�1b�E�QTb�+#�AU����
,X����,QTXU��cE�
�X�A`�PTV
*"�EF(�T�
�ő<I��'�{�Z����	�П�I�d����O��� VXVN2�;�^�����t�ɷ��n��
|��8²u�!��y���q��d�*C����{�]��zʐ���r²n�ܻ8�����`VaY<eHr�~s���r²wlć�R
{��n6��]72�ts�<a�
��T�m ����g�|�+'߬ć���a�
����$=��� VXVNm���3�i=@�:²u�!��w�@��
ɻf$=� ���f�~��D�&��יn 9�+[�r��n���u�\�� :�2�TUUm�YM�3pLrn���B�u�!�c�fJ��}���ćiH)�a���T�ϸ��)�`�d�ىԤ���t0�
��*C��S�
ÿg�|�+'߬ć�R
u��²s�~��pv�q��\��n�x�������f$;y���8AO�+0��eHyi=�>�40�d�ىҐS���{�v��*C��S�	�M���OP�a:���^<���n��k�V�	�	P��	��	߹���u	�'P���;�x߬��򔂝@�=K���}|�x�Xc
�ͳ�zSH)�a����֐S��W>�L�q�黮��0�²nُi`��
ÿe�VN��;i=@�1�C{ϖ�|Ϟ�P=ed9~y~�H)���'w1�H�w�`q'XT�Y� �����'���훇]!ӫJ������1��K	�I�����>�P�d��ܰ���4>MIԓ�'�߭͒q�ܧ��'�m��'�XO%a=�����z>\Y�ty�[<�]Fĝtn��<���;m���65�����UV�&����㹛���{�d���: ~eg.��8E=`T� wl�C�,���~���>aP8��v�<`T��u���Y����
u�Rz§|��s��AO&0�m��~�F��y7t�-ͮ[���䂝a_-�?[ �{����wl�C�Y=`T��.B�u���J�T�>[vq���AO�'XTYR�9o�Y&0��I��z��~ƚ\�qsp��|�x�u���;��|�'ߩ'�����	|����N��d��ܤ��~��o�'T��[#���3�|��Ld;K �X'w��\76��]�m�5���-�Sֹno�W9���)���
��������$��Rc
�ݳԲ
{��cv| q���
x��}��C�~�)`������K��]]ێ�3��C��)�
�-��;�ˆ��T�0�ed?[ �{����*��{K ��
����T���AOX&!]�>[yϩAO�'XTYY������i\V�A8�37r�*֩��	X�����|l�0U��pe�u������e�x8y�+���9� A�	���*�
�ۃ�.���p�(�]����b���Z�y����iͲ
<�҇Yՙ��]a\7!�:�_9��<dX��V�g���U۽�i��T�@*��y[ٹ��mݝ� 8��*M��Q`�7m4m�^�n��{�r  6��  *��v�osU�D��u�<2���Ngغz�m�.۶½9v����U����9�n��n2�|#�*LaP>�1��K ����́ĝaP?�VC��)�����O9
���1��K �X'�>��߹<d;l��0*G,*6�d7��ٻ�$��Rq�@�+!�
}�S�ܣ��e[���s�<H����1��,���*O/x�@����
~`T�XT����C�Y:��: ~ed9{��9 ��
��
�ݳ������uׯ�or����Pn�d/7�1�C/�Ns��7�%3~���9����ws=�}���\��)��r�4��j!�E�m�GG%l9����d���: z��r����AOX#��f2�d����: |��v�=`T��}k�!P>�f2�d������~s�<����������sz^�Ԋ�WCܐS�I������)��|́ď��f2��S�
���9n�P=ed9l���#������C�R
u��
��� �ϼ��=@�����1!���������v�v���@��]�V�nɆҽ�p��s<N���4���U]v�+v�[��8n]��u��<a�����AO+_�o��d����򔂝@�=aY<��.�$=���@����m���3��H)�a����֐S;ـk��v�H{JAOP+�=�/��7nf�弅d�*C�H)�`�d���g� ���XVOYR�<�g)�`�d�ىԤ����a���T�m ��
þ`��VN�f$<� �������k��r�mutwq���!�H)�`�d�ىy��wt�>@�8²u�!��~�f�����f$;JAN�Vq��k'��ZAO�
��
��$������>���f� �e��3Q��Lv�O(bw�=��gD<���.s��7�%3~���>{��q؝v����z�̶L�6``?q��kp�4C�xl\6q���'��j8�40����V�Z�b)%.�(&���Ҹ֝��w������e�sx�mm�b7�r���u������BG��|��H�  u�:_ �h��+���p]���q���m<�\�������D3��c��\���1��)(KtR@��$:�?�N�GR:�NʭH�D��Y�ʑ}#,rR�
ظ�A���g�[�(x@�GDB����Awƌ�ׄѣ��g������AF�$
��ݟ$O$q#ʁf�H#�K&�5Z��e�9��q�>|�c��7�p0C�y\:��Ԅ��#
78��n2f���z�M�8���|p�/y��$i ;B�`�xg��_l*	�u�D"i�9h�nƁ�u�l���F� �]P�.�-J�v�J�c�Gk!	9��zɺܾc�o�������������w�.������r�����*
ך�����4�"�Ĉ�?Y��-�Bd,�-ϴ�!Ʒ�D���@b)F���s_��`��o;��[���=dCw�	�R������:���z��|��ޢ~����Ie,�W�Hî�i����%�u#�i<�~��(xC�?do�~+��ޤ��VI#��w�!��&��D$"x�#{D�<H�@h|O?��=�zNs��y�;1�@�$ֺg�;pnv���k���&�d�H�g���09�M!UWF�u�)y�KmR�ǀ����g8����nV�?���̏�����,�g���臽��������J����o�����~�	��s��8�g&F*�!�`|f~��-���7��䇠~��:X����~�5��0C���5=|~,�v���ǁ�������T~�Xj���"d���ۉ@eqHh��[o��D�F����Oi_���p�<!����m�m�F���Xq��|!��~n�u�p0A�f��Ϥ臂�;ϧ9�}�K��~�0>׺�lB�~��A���^fV��-Fy&�����R'j�\�\f�Tī�kn�SOl!�Y���m��qDm��Wa:��$�c9�C�<nņ+u��}}��:�Jv��s�Wnڸ�Ѻd�k��fL�p����F�M�U�\gi�aq�ImK�޾���]��P��tY��Dm���nx?��T�s�7i���Z[�g�v��  kklU �ۛ]s��8��2K�l�J[�z�l]n��b3��8;���l�(����!ّ��JO���9d���``?�s��s�!臁���޾?��N��=w�=x�k9����vQ�+k��Jܯb�\~ª����T]�~jJ>AFA�i��7�rɂo�r�8%��/�D�qƢf@�l7w�#���s]��7�O�=����W^���j�_3�:!�����+�ƻS=��}_��%d��?�pxtg{N��x~�ʂ���]��5m�t�  cK��|i%���ʬ��>����v6��vN�~�	����pA��Y.n���|��k���9d�8��f���tb6ºs���]8&�;h��1�9n�Zӎ���Yv������Bm���6V)��7n�s�����˗C���fY>�n������`>�|�Nu�>��~��c���K"e}��7�#���於3�Ş���<?teA�]�	.���;9���UD��ф�m�;�5!�Έs8��q�h`?í�;����?�s>o;��n3�K�u[W�|��z��m��	[���o�rɂ�7�pn_��[��<!����r����7�O�<�o̽]z�yV�qW`�j�DN��cv�<�:�_Y�ԍ�K*�}O�B�x�ƭo��O~��s������� ���V,ɍ�9]p��=�;v���6�PY@K��Z�UJ���*�v*'HJ�;���'n�(�Ā��/!�nh��aG=lFu�h#�#�:�'��#i�%��4T��%#��U�q����<�;9���Y0C��q�_��g9�9�x!�|�5�~�2��3_c�2�d��Z���%rX��.H������?a�:�M"�F4�r+�<t�w�!ma�bP(T�j4��#E��)M?qC�/��֬���C�HçĘz��43� ���xSA>~-�q�y�E�o�El%�Y���?iwI����ۡ��yŋm���X;6WkZ��{vІRuV2q�\���nڻ��a	m��#GZ���)���{��=j��C��0�!h=�_�F#ۼ.Xp!Q%!!�(Ymi�}绍=�3���	�'���-����E8&�Jg��=�/զ�ƪ-�^5|5(���n��*�x�$ka.bT��n3��5���[dt���I>�R4q"Y[��{2I��t���_=���m��i�|��gl���YZ��Һ���\x!���s�խ���������~ 3v���8E8@$K�Th�@@ƿ���x���h�M^P�U� �\s6î_!�; ��L
�mV��[����+IF�u���?��6�,ױ�AA|���ޤm"YU�y�ʸ�Co����9���Y<!�C��϶��+d�0����?q�w�����m�.L�q���'���:�ۡ�|�5C�����Co'wZ����e�$�|��g,��7~��t�µ�2�>��"��!s��]�֗�no�!T�	\����j�)�8�Ե���e��|}�~"��Fѐߘo�� �7�D�	2'�@CqT��B�kO٨vR/L#G�RJY��3���#�|e�}�������'$��QUb��EX*"�(���,�R)�V,����d�IH�
H�EP�*�R((H1�QH�TTYU�(($ @ E!"�`*�X
��T$YE���P��B)���H�$����a,�`(
�,b��P����X(a$X2
(�U$X�R(	�(UaE�"�d�����*8m�@�'�:n����we�h���`���z6s����m��m�`i������nL�V�X"��X+z�U��+*�E6��� ]2���5Jd����6¨*�{e��  P 
���;�ePs� � ��K�{����F���x���J��HZ��J�V6�\�;����C�s�d������ۖ�@�r�\���.�\���髗Sː��zzN8�ƌ�/LG���N��Lb����8�6)6���bI����:�4O�p��p�>9��U�3WuF@�cbQ�b���;d"���i*�1�	��T��h�76ˬv�[����#��v�8as�F����8ݳ[`q�U��
�:�3�����U�)����1�exݎ+���Z���7bs�6Q37h��P,�ĀI�{[�r8 rTl�jݺ �s��]m3�d&p����2�9�s�[c;��*�q֧kv�b��]�{U��*B[��v=��˰ d��9tKmڳ��6+'Z+�h�XL.=�tG&KYv�'X�ctbc=cG#��m�m�9�s=u��복u��C[aA|��u��|m��ظ���݈��k&a��kW:��_n�b1�=sa3ю֘�ݜ7i:ێɤNzx���S-�~�c���+���8�uMdy����Q��q�h���mc�lQ��uNθpt=�`8�Ew-�){ ���s��P�ss�-�y�؞�.y#�r���VV�;�`a�slc;eࡀ[m��  m5C�P*U���AU����wwwy��=Z�(D�Ѻ����w�� 
�k�]�<�� �� 1�p�� �p0^;c�GW�Y���Tp� �T��N�m�{��؜¨+�w��#,�y��Q��[`V_U =lTm�m������Q8 X���m�^���R��]� �v��$             ^���  �   P� <  T      \�
�~���m�gf�37F�j�*[Fl�&b��ΝSr@[��mun�݋gR�~F�����gF:م�\(�m�F��������ܦ�٬��Gi�6��p���C�as���5���f��N�Λ��Hl\�n!��7`P�#A �ޭgǕG��k��獳�^[���6ؕU�����gm�  6�0
����h͖
���� �1�L8@\�wgn8.�厞Zಀ��R�UU�c��S�v��bߟ���o��������mTNhЦ�4ٙ5		��o�dS�������#��+���{��ͣ���n24�p�4Q��
O<H�X���p��.���|��g,��tse����_��Bбq���5�s����xC����R�8�n2�23��C��������!����m[�K�l���U��={��yӏ�`�vܬHĉeTl��X�PD�J�;�D��|!�!���
z�mZ9v�F���~�3����`��ͤQ��^8B�(��'�$t�7���x!�"�&��[�7%+��Yj�8#v��X^Ǜ�k
y�1����nMH��3UV���u�7f'iv�/���o�n3���q����<�}��}g<�3����?q��N߄?~����k�Y�����_��e��~4x�5K�Y�J�G�G�|+��n3�2`�_�<��t����e,v~�[��0C�C�X�ĈH�@[����%m`Q��q���z���40��:�$�,��ld�H;u�C�}_j���>�q��o$�q����?g���l�\~��i�i��2�Aȡp8�5������pq��t�C=~4x�3��*>;H#�#�m���I���|�gk��Yi*��6�I0񜋲]r�;[��nrDt�����nn��[zA�*
!IeV�n.<���o��xC������7���NN	�F�
��0��͇�[B���>����oյ���x!�'=������f�jv.=��ӳ�o��`���rk�Ua
Ul��	��n2g��?C������2y�ߣ�]z�|�]P���C�����YS!I\�s�C���z� ��Ō1��q΄�8d�1��M�L5��ƭ�m)�Vݰ��%��8h��A�a<H t_ 4l'��>�����p��gf�V�Ǣ��jwB;i%�~h�T�T�9�Ή��s힯l�d�"�2 ����@]`��4��yI�������p�!Ù��7|ܟ~����|x�`|!���[z��8��փ��k��X���c�<��}9��7��cb���4c`h:O܎t$A� �%�4Ŋ&�����9��t��8o��A�ix�4P�AD-����L�>_j��|hv�q=�X�V�GISkh����BO44d0~+�C�ǆ������U��ZB<���lz0��-&[x����4c�Ж������1pch�Ђ���ďwtBnueNJ7!�x�8��0�Y�&�P���ֶ
�4�]Mv3/�E-U[n3�Ԝ�d�ml��"T{�λ�J���cYb��~�}���`��1{;	8Pc	hʥ�>�;��9��x���BQF5ܸ���3L8E���O-i�N+�F"S��1�܂���E��=~���F]r�+g��`��~��1�GYN@T��8y�yD�O�p�������N>�*�ʎ�M���~d�&/��Q`�/$TK	��ě%�{|}����n��9f���[G� ��$�U:~]ؔ��m�-�$�����e�XԌH	��T΁[h	�&ԛ
�F�<�8�6�5ֵ��m���0&x����j��^n;a�)��gs�a�=�|�qD���nwN�ָ���P��-�@�#'E�NA��O=
������x�won��*gt:���⹶�謥P ����y���6�� 1�{l�z��Z�,&��+�p�v;������  ��U
��Z��g����+��h����^'x�^��۱�-n��j���35F�4�Dی�2 �*Bb�@U���{���H�,U/�-�pc��+g�?q����T]�
�q)7!l�b�?Ywx�2�E��La�#[��R����P�Sy�R�g�]�Ud$R8P$a��F�#���uء�����#�g_du��D;�^n�qC��2e"ْFʌ��5�J�y�z�Ĺ.��.��
�PHO�gq��U�,H���E'<�hv���k]kٟ��4bå�Y���Jܴ�����J�6����=��wn�̗���s��p�
Q�B�n "�U����Ib�FʅG"i�لa�@��W�a����U\�(�[Z{B�y24��1c�Gen�!,��]v	w��ĘdY��Sua�Ђ0�u�3����N�^q����b��C(���� I��l�uu*�-"YU��
���?����3�F��C`8����N��z�V������w�7��ٻ[���7�#M��
<�8�ďuϬ�cd�#iI�MVpo���-�v�����t�z�@�!�  /L�n�A��08@� U��A�3��-i�g�rq��4�SV@@�)g��Q`�`��ّ��j��ݍ���ˌ�p�Y��il��.����7�6�@�����H�~�;kn�2�.�HC�#�I���t� �AǨz��r����1�����ާs=��kj��z�Y>繀�G�$�i�q���uq.��N�Ӕn�DH;c}�n�x�dy�����m��oY�&x!��	&�T�h)�?i�I.���q7���5g�W_�n���0�.�x�-?i���Eҹ�8����M3�m������NS8u�3B~�S�\Х=���"y�2�^[RsG�������+�yΕ7����b�M�mz�u��t�O���͚ۧ��пA!�$�nv7h#�#�ve�TI�@�[KǢ+�d� �����L�C�r9[m��>��o����rТg{��fsy��g����ߟN�A��6n�#�}'D?~w-m�o��9��$	��$�D�l\x��n{߭o̡���o��������'9���mݮ*��<y�GYG�YP�^�m��ۗ��`Q������@H'�@�0 D� ��%���8�m~��Eɧg5�{Q�$��E<�d�$�D�sd����tC��}z>��p���<�}��� ܎~~N��?:��\���\�PtM�'dXtl�үY:%[�l��v�m�&w���8�lT�=��Y��H�dY�z�sO�F�2�\����5��5��֮_#4�G^?��g�ovɟB0��撾D�D�c�E	n�r4�q�ik���$����)�Fڢ7z��wZC��JZA�(������q�e�O�E��E����wŌ1� ^$G�{s�Q�??�ʈs�4̍�8ݪ!v�SO�����?Q�Z��aT��7~�����gjU��!��5�ˇMV�]0Z�m��[�k|����]A�0�
�ZƦ��-\ˍ�%)d�$�r�����ڱ\`�Zg':��xx�g�]���ai�`#T����톸����m�ra8x��֋V���48]�ӌ�"N�{���E�ݕj�r]O1��5]Wwt�=���*���Rђ�X�!,�zl�[כu�l�T  �U
�6�=3m{�5T|���b���\��qa==�znX��4�3����,�U�CísC��2���� {4s�L��	�>f]�����m�@v��2f�b �P��#L����^�)��G�2i1���_a�Ō1�?a�����	a�Qe�;�В�~���_�Mڲm%4�/[�Nj��3�|�dG$�)	qDk�E���� N�*.�2�L|̻,���Px���Dpe�D��N5�����=���;j��d�E�q[+�ig��,�4P#p�qȊ��ώ]��w���;��j$�X��g2k�M*�5��eD��-mڸ��y���u�{���V�~n��i)�}�,$���a(�"S�sU���m�>TY�S"U�pi���L�X���ֵ�Ԇ�!�b���*����o� ��dou�e�����ӏ�]����9�w�� �r��J� {01��dĈ��_�$����u���v���Si�J?�	4�
�5����sU����}�N����+m�m���8�2�Om���<?��snD���.��m�s��[��P6�f�vt��来ضU[���
�֊"��   �"wx� �@��g@ }�$I�;��  
���ٍ�D��o�É�}������$�`-�ˉ�$ ���8ix� ��B   ޴�wa ā�c�kn>1H[.4EI��ċ�ZUG�UU���מ�3��?�Y"�H�E,$QdD �B Y X�������U``�(	 QQEb,TQ"�(�$��@�	�F,�b�X��(���b�d`�@Y Y@ � �(�`�)$�
E1EEVEX	���Ͼ��  �W�KE�$ d��$��]���r��z޲�L��1���$�Vvk*�R$�H��y�$���o�y�ӟ>��m���ԑ��`�	L�cv�$�UA�I$�R7��	'$���!:T��D��J,�[m����ɶF�
ܶ�FZ�[��l���J���n�<tZ��g��W�32����',�6&��쩇{��x�54� P}�HV|N脀  z7�藒$�Kk���I$�N�9���S�����2�m�m��{��^��`w�L   0}}��$ 8�9+�q��Ͼ���x�F)�ƥ��Q"��g�I$���S5�ݤI8�Pl�I6T�Ń���I��!:T��[m�2w�~���H��)���m���L$��@�(�� �%�B��wD$  ѿ�oD�H |M��Y�c��Ydo�m��2rG�Е��D�oع��U��J[m8I$�a7�xg9�m�p������DR�a�Q��I��Pzɟ5�(ˊ�{<g$�l�T�j�U۞�k�t;j���?_��<���ϯA��o&�A_=����*�d�I��l�$�H�O{A�k��',�[Z�]�z�Y0oc���o�{ss���n�m�gC�����q�6�m���,P$��!c�Q��֥iM%���Q$�t����
�pm�ې��P�6�/�J�m��7� d���AaPKQ��6�y-�q��·��_5��6�m�۪���m���]������p���KGl��Fq����ه8�2����cm��}f{ps���15[m�:�Ӱp����u����-�s�y�B�(�`w ���ʷ����1����ԛ���5�N��'C�3�n�ph�N��6��^m�1�巵na`��vy�әm�bͮGh8�rl�n��?iO��������� �Z*�;<��l��]l�\�nG��v3��<��QU���D�c�%Kv�.o{Y��8@y�?�>������D �*���e�G�  9� P�mݼ�l�n���a�Z[��-�v$��}?|���AB��lPm)r��ֵtd�s�W2lX����UW��v/=��Uyo�|�^qU_[��dĘ "@ oS�'� ��Im�j�������m��u�����#IHT��  A�,��6��Pm��37�G��������,%�����m�A����z��w�Aib�G�Y$�Iݼ�����q���R��n0EI8�A�Ě��I$��MYVn#>�f��٠�tP5
��%���gua	��P}W��VF\��s<��f;�(��� ��
:#�� �=�]d��hl�)!�L�1�BK@m�Z]�:頍j��k���a�����e�#O˻���d,Ԙ�}�5��C��!r��aA�����5oZF?�a���9s[�nή�CNH�r"�m�Ӯ"��^s�������4%/U�=ovs�v3�%�b�7m����ky���4�բ��n������a2I@%��Á����Y]>A��{��ʢ�0���EZ8Y-v�]��y���i}l����+����a��i5���hiGtr��jΛFg7�ߠ���pc3��x=<�*�Kႍ�Ԕ�VF;w@���D�i6���Hu����r3*��;!�`��9R��39�/�Ǎm�dSI��Z�r�K��kb��OH���Z��di�]-�;��}�Q�O��'�8��G"S��+���~�O�kf�nq�#V�pa��-?7�M Q�E�r9Q�����r�qY�N�~u�=���)��@���2�UD��Y�g�M?w�$�d EQk��Hkh��:T��%��y��C�;j����T�y��D�R�*���j�Y�� 1iOH��sMWbN�:��#��'��ⶑ�Z���UJ�~�֖e���r�Q��k�.�����#1�P_�Z�@hvGT�����!M��HK=���6vW\��-Ք�{�j��Yv��N�U��b�i�)�8�$��T���(����A|�-����_n�9��疳z�Z�,r+#�������-������i�����o��7��g��?{���t*Gp#ѝ�\u�Ě�݉�k���l*+�յl�Ce�y�c��<���lZ:ʭu 
�)L U,����@i��_��d��-�����3�0����))����[���W�@/U�}G��q�5o/�Ŵ�� :]��o���j��,��s|%����w�q��oĿ�Q����e>ә��&�g��"�k{X�C�%��8�~i��\�Z�@z��@�^��)���gm��~�{�8J���)bu��v8���?x�����[���W.�^���q*�Hռ`�W��d���L�gu\ײ�(p��*����Cr��d�u�nzl�ۇo�W�`6�&N4-����j�9�+�S�;���l=��'�If����)�;I����Z7\/u�:6ڢ���c��v���L�cv��s��4q�<���4�:��df.�o3�M�<KHMS`&�i���ԗ��]��ط����:]��Oa,�u��  Sl�T*�3����wj�:�M����b��v��/G>���n���jE�,�dp�V�-�'3Z������/�ɳ��dzC�)�>Ү�/�fY4e�O�s>[� ��o�L���{�9K]��t�Zy�z���U�)�
��O-��t�S��L��{��wL���C�f^v�k{��|��L���~5=�@���GJ�ڣ���p�g��V���m�l��Y�Ew��(�$r�y�}�.���~�3���U�5@3����V���P_�\��������Z�#�U�>S2�g]�^��	x�#Ѱ���	��lR�LNEk��l��s<%��-��|N�]�
G�@]��N��@Y���/:���!� �VVR�*A�K��=�4w�{c[f�.����A��������|��h�T%�)cl���}���j�]��^t�W�)��w
jF)R[@�3ڍ^�d{s<v�fR*���~��&
�4A	��XQ�)�gt1wwq9�=s����������9�7&� Χ�u�����i˚�%v]dM'�UV�n\�d� �l�h�R���1f�k����K5z�I�l�S&�T��>]�~���o�<ծ̤Y��56�l�lEnʩ�~﹦z��a�ކd}����^�el���2Ax-N��[�_j��,�T�e��ϛ�߲w�p4v¨1�,rF�6xn�wҶi��,�2��,�r��S=<N�j��!6�7&n),v�}��c�?9뎌���.�2,@f�vδ咺/�-� ��ߋ ~~����t��U���t�W"�t����Qm +Z��n��R�Ii)y�)������	c�i��Oq�����AFgY�.�}�3ḻ�)=SEU�:R��x��_���P��s��U����)�
��O-��)h-Da(��I���KuU.��@qd=��n���= �WE��ʖ?5��6ũ�W��Hʹ���4�E��ŧ�a������S�}�;�/�f\�U�� ���N|.um�3��;�Gl[�0y����
f���@]n������/U����?_ ,�_�����޿�t�ֹA|����֔�R�m񅸢q��$mFR��<�n}in���_��?x��w�n�U��.�^�������iIq�������T[H�9M�1|Wt�s �]��{��k�b��2M��
�ׯ}Џw�m���;������:��͛��8��Q��)b1��I�{�w�;�Ug±U6\���翺�B����fSq1i�Mq�u�E�1<��(�y됱��`N�7a^v1��HM�sN���V.�s��R�F��쨨U�UTR%���+"�J�� �A��-t�]�mP[j����@*�  6�UCl��Tm�$�*m��wu�ٕi�k AU*ʮ-a*����Ӈ�-ؘ���t�xe��f��Y�ۍ���b�im���uɷ\�*KqIm���.�r
�z��O�Y�e��!�s3�X�8�뚔�6��l��Đ�̔�����{p9wn��5`C�c�C�y#K���ǎГ�9Īh����}%�������$��Ӌ�|�d�T��g�u��7E@m�:S�Ƚ�cB�Qg�.����̓l�Nu���$i�����u�ض�j�sѹ��[�g�L���!��n0�N�7]�ܜ汸��%��U����<�/9����]�t���E;X:�$pa4j�M�h�v���6+�`3��ǡK����a}�A �L��d�W��5�92���.�y�nȆ�Aŕ������h5�&��S��NRx;L���"������C�ŋ��g��7:�tf�j%;q֦�J���p�]cV
�pc�H�댣��)�0c\��W�y�s-ү<�^9^%�� �s� G�ݹ� aۆ��1t�U\8I%œ��#9�v�E���Nܮ��Wm��m�7mtm��$:3/z��,��v���N(�v�ֹ�e�蝜��v�+C:[n�fl3����6�.�.�J�-� N  8@U U@ �Xo+n�m�n��*u`���ۭ���l�^�1� U\��u�v�` �  < ������W���6�-���.x|�<�M[lQR�T�.$���U����U]�P6�{<�@wL�TU   < *�������z��wZZ�ݪmUR.v�ݝv&�X   �        ]���i* TP  �           筊bɧ����B��APz}-��l�l����s˝��Շ!Z�X`$Z̪<�^&��ݵ���N�ڷX\���s�n�ltW[��r����X3�`\�N�΍��Z�;fCnw�Iș3R[�º�;j�kqc�6yzv��"m�N��{W&3�=�;/�Cǲ�ݲT�UJ��l<���m��s��]��dZ�y� LĻM�T -��}�@  �m �TQ�b��Șӵ��v�`�i�N����NӞNS/'eսԀwy�ή�z{�$3� �S�����:H�wq�����+3���u�Km��8�/���V[#]}�O\
e���X.%�Lf��(��O)�ԟ4��0U^e��;�V�ʄ]e �a��8Ō�-�jv����>�j8B����5ϻ��p�s�P1������ў��w��c�l�F2˯��K�����$֫�k���ۗN����B�c�&�v���J�l��FU�d�.c��"�19~{��^�٩m��LxR�̳�j������D��i�#��*�Ĕ���ߩ麕�);��M]}�§����;`[.��=����ow�+��oFr˯�rT�D��4^$�H�辷vbUvwS}��)t��%u�~۷M�"B&�nly+l�R*�Y�^��"}̙ Ryg��Mh�h�֭r6JBF��L�Ԧ�}��] ���.@�Z��*�����\�E,m�_��Mn��p�=g����֑e'���� �-X�u{}m}$��j�p�_Gf4l� f2�`���8{�l;W��[gP�"���ϩ�c��Ii8Sm&��X ��I�|�&��3����_5���n&��-�Xn޳��zYp��K�_{��}>�Ŭ&�K\�Y�]�B��z�:��3p�6w��=����2Q�ۣ�-R��<6*��m���y@wy��:=�k�*ӭn��>�ѣ`�Բ�"ts��G�g������S�>�j=��)��x�%�� p6J �K�֔�-������o������o��R�/�kvж��}S��TF5��N���Gw3{i��,��l<xX�Il��k��}��p�ûy/?C󋃘��@ 4����x��[u�m�Սɀ���%��D�%�4� y��]��lO8�	��w��w��U�[��e���o�[ˤ�.��IGT�����廚�쾾��������<���Ξ6�0��2�2�i�w�����t	��K��ӻZ�L\���c&�lH�٫x������n���Y�_�M�*I`��&���[q��\F�n
WwiQ0���IJ׼�{���M��uz�h��j�\�u�U]\쭵q�町�7WSsVܓ��=[��hs�:��[gˡD2�ݗR�:�A�+����.,�LM��E tOF��,cnwk��Wv�8$�mohoeջu���Ӗ��1���ٳ���\�=7n��рuhm5���
�wW���l��1����#2����)���=U  �� �U���Vۇn7 ��ٷeѼ��+!:�,{I]T9��L,ʽ&�M�Sa��E�~6l7A���{e�'�U+ѡ^n�|��ɍ6�N���w�;#�����rɺe�F�w<ڙ����B��ۙ������537R[j�׾�Y� ~L�R%`!a?}��u	#�w殅l����#�D�n�� 3����e$�0ɼ���{v�jL����p�>g�&����#mX�$���`�������7���윦U���e[rH��X` �h!w���_��� ��E6���wYܗ׾��E��Q2�Z� ݓ{��w#e�J+�KRj����~r&�M�!�7�D��+��}�f�/-���]m���~�P|ZL��Abh4����-�J2��
@O��.���DJ�&�E��0 �ص����c^��>�wu�eZW�&\d�Kf��n�cm�7[���mս� 7n*ɞO7l��d�r�g\T�+�u�n����1����=�Z��{�f漬����U(,T�,I [a.w�q^vV[}o�w0/yw6��0�����i�}8�OU�v��	5�xw����d��A  H��)$�n�)I{�Gӹ�'�e%�Nn��7^^u�,w�l��i4�r���Z�QإD�/��l�ё�H (d��7������-����ݝ�`շo����)��U�J� �Ue��L����/����?�]h�}3�y<=�c��j<%�����U^�܎�ڲ{�&{x��$�@��h�hae�����nE���W��nGd�R]� �KA��,���dخ��s�MU:m�ݻ��I����&b�0��X�.s����n���E(�=ɓ��}��N [i\�0�cv/�ۄ�'���ۜ��;`�Y]����nJ�m�Q��Yml,uT�����{!~>ϣr-��Z���6�vz�	)2^&BI�PB߾��֙6k�U�9S�L�tۇݧy�y B��L?�6�E��6n��r{}x�U}�c~V�Y�Otx>J�p4i4�2�i2��fs��e��}�m�~��w�hU10�xPl �@"�;u�,�[4e�M��߽t��Lۘ�a�k
��ƠJ��x�[!J9�^j�(���V�ڻyu�Mmpn1��nk+�ja-��l:�.�=f�SHՐ;sl9�	ťǣu��p�����g�.[��=�m�7[�j��R�����>�s��]I	���3���y�ƞ�׷�d���8[��ݻ{�YJ� ���G�܀��� 1�ܶm�m�9aŒ�N(�cn*7��  *��	V�51��S8�#/]pf�؉����s�����=`�[F^�SrA��Vm���)T��a����a����}��Q�<z��a���T���$�`�m%�r�ɰ�W���y��\ϣ/��!r/��U(����~H6�O����r+j����i�\w��آ�d���)"��3nz��i�/�v�]���o��!p4����	Ab�Z!��f7\�d�k"���5��6p�3�V�=$���`�! ��kt��P�va1Om`|�%뢚Ԃ��1[,�~�H�԰%��H�a�׳6��{���cU\"��e�OJۈ��  ��I�O���fW9�>�k�s��{E��h���1���},�MZk~R�"l�|��ϹD�$ΧRl�&�ĉyWov���k�߶���GaR�E���5%@�g,6����'�ہ_s�u	J�9p{��ԃ=�O�y�dn� 1@����Ȋ���*vIU�[{c��nk8Nz��� �u�J�٨QR4�1�$���m8���ū�������#�|���o�	��q�Ll� )5�}�p��2f���~��ս���Ն�3] ���hrPp�r߾6�֙=5�*���߿~�ٟ��5�q������{���V�@,K@��w����w�7�t���iF�=с�X���i�
����A���������"�ٵ����4T �<�I�γ(��+�)cq�iһ��7F-�9���h�,B6YV�`]l��f�1m��[
���~�h���}�q[�s(�N�u�dVV}�oԃ;w˷������Z�э����(Jܐ�R�f}��ÿq�bY����:��w:]�vK�M�4�E��;�r��J�^�[4e�M��%_s��� <��$Y��l�9�x��j��+��d�]M�9㘵��sР~�6Mv�`��.o�p0��e��w��	@ͥ,:�GEW��-#�q�YI4[鍙`�򓞲!�ړ��;Q�������d9���24�i�;ړ?;�v畉(�vΣ-�̂�H��Z�!	$���w��,�\{R��{_����!?(lO���}�%:�t%}(��O*�k&����P�qa|�	$J�I�m�)��^ҙ���;s�ĉ�e림F�1@4��  �l���sn�P�)ur�+�޹[kB�'QH{[\�I��q�^�ٵcbmACƹ9�u�m¼(s$�j�� ��gFю�9�+ўId�k��m�)��P��<!���E�:^u7t���lڃ�[��{ksq�t-�ua� 箾{m� <�ST�];�cK�����oUې   � U<���w�6���{m�[Y���;[Q�X�i�ţ'(-t9��0Sۖ@����{-�ݲj�H7�ߔ�E����h�f7+��G����ܒ�����D�1�rF��c���$�B��(��򓞲!�ڞ�	�ce�"26Ɂ���˅�n��|�/��AG�{�۞V$2�фX�%�)�%���2ϔ�}��梻1\V�=�-�>�`��!����$����\���N���譛�[!����Vjlq}e"%�h!�ܢ�m���9�7D;΁���z�`r3�<.7m5T�\�B�
A�F��3�M�y�1I�D�����r�;~�����(K�B��Z+NPC���$y4[����۽R}/�/{�2σ=\�HӃE0	���L,�n�w`K��f�.�����񮻨�̕+�?��	~-��q��ݪ�.W���k;���}M����;�sk#
�dS�n����bQV���s��)>����Wp�?��g���ntmWX���<qd�>`��ۓr����Px����v�7N%�Gk*0S�GW:m��Է�� �n�v�:����2G�ym�
�B7dahlzٽhIO������j��>�ds>�'�ϤKD4Rm6�/��Ag�{��<�HUY~���|���3~�$�c�	�����GW9ʀ�4���"�*�e�n^�c�.��E���U̧Ml�ZJW�'j���Etٙ��'���9#ak�����J�9�zƪ��&ދn��+��h��̪���L��~-00'��'�e��_Eo�3����6$%g,��r�q���%��9�诱{�ю�,J�t��ioE��n��
	g�$�a��-�Jx�wö��D�+�V+g��R�.�UAr���(�E�'̔�2H�`���3��73w9��w��⢹����'�x�!�X�86g�k���I�P=�j׳����[��s_�3�#��Ń���A����\-U���K���8,�-UU�\��%;2��L��7R�����sQ/��r�j�n!����F����%+"�>�Q��z؄��Io���r�]�3ؒ��s�-jH'#����Y���������8�z4��2Z�dm�
�+�$J$g7���S+��6P'�ow��=ڢn��V�l�D.2Y	q1e�
o��v۰y^�O����N��{�-���ʂ-/� H-��8Z�:�X3�UWi�S����l�]��.�)�q�
Fl��v�ƳJn�d3pbg�v���O�{c�8q/uغM3������aڃpu���X^���ϱ��[��3)�z�'< u[���9�j�-n���s۳�g;K�� ��Ӗ���Mk�L`�l�b;���/�s���^r�;����H  �* *�Wqv� ƹƱs���2U�A��T"��;�s�®��4=�L��$r���Y��$��Ц}��sgH�|�w���p�7'���ލUF�\�Z����%�d�o~�2��EvUf�	e��E�9����Or$�L�� ���B�[>�B}�Nߙ���82����[�hM+q$S��	�fr�)~E��z��^-Q�_�]o�'��D<���%�h���حȔ�|�����v�'Ͻ��o�"�@"$���!��95�`�v�7h�JCN�Cf��'Yj��O�Q/�	���TO�]7t���*F}�s�D=ڢ�����q~$&�x�R�I}�����Q��h{���ks{��z��J!9],���߾�j�}����R,��ߜFz�A4�̤���A���՛�y�����5���+f��6�����p��ɤÐ�����!�˗���p���m�(e������'X��@�B���%�v���3۶6㵂��Fu�82�!3vh�;Hu��wsZ9ޯ�ÃZ�o���������^��.�˱Z�L�}4i��-���#v8o��[�}��ڢ�j��;i����e���8�OvC)&�H3�MU][ �3髞��|~S��KQF{l�1�t�NRE)�̜�o�������O_]'����Y�(�/���!@�p��d���_+���v�V�����;S�+H��*���T�&}�|��P� z��i
ƺ7H�!������mk�f��S�,�\Ie�v���9E8�yY*F��ݶ�W�������w�_)��6v���iר�������@� jBZ�j�8�K
aˢ�]� ��c,��<~�xO:S��u��v�R���%$��sZ�Ʋ����Qu,"���0���l7�����<�)��q���~q��vHKQ�#�y��M�b�\F��:ons�,��Gw���Z�sB�C���j9}��\�IGo�A�k��ᆘϴ��">"��u���YK���Y�%i$�H:�1su�������'�rG��׮�>yf�2�Z��m�X�]���inh�C��~�6���Gpמ��)a��S��.�mXJn+#N���!([�l�Ye��2������֫O7�I��WK��v'@ȽWJ�B�G<jl7hBJ2��q}��p�������������>�p�4�}�n����]jg�lV7
FI*��C�i�<'�)��:˗��kh��]F�������_5ޗ�1奐R*�X�[9�:�?����y�f3�m��Y��1{�%-�?i�8}���o�y80!$��׼�ww+���m���������5D��[e=�a.�j�ܶ[i��SuG�se�wmD�Ql���� 
n�r�Ƒ��r*PlJ���M����=l��m���   �ؠ�iSq� U����^��me��A��Xj ɮF�	�){iM�K���!�;�w�m�7e����jZ��:�����]�mF����6ʱ���l3��q]���nb�#��m�y�n-���Ǻ���۩��/G9.�T���[c,�Wc)�k��,F�e�[��'=��k����
�\	�mm��nq3��5��e�vv.�-=ey�=�^,�9�%�$<�Lْ���t�@Ϭ�lsg�6��Y���H����9iM5�m57[���Z�9R"Yx���J:��TuA[Y�G��6x�ٻY�==��踸�˳�"q&� �Hukv+�!l��>�]F�ӻ<��o[V��K��dz���N*�ץy�P�u�[HZ커3�<��N�y^��<��něn;D{ث���W@ZἼ)����,-���	6^6��O�Aj��f��ӂ I2�����sӎ��ke-nEs#��6kX^�;%'=Ӡ��za�c�1�W��g�0g�n�;5s�T�g%��x�28��v�Lػ	�g���Y���<W$���]����r�h��1G7���n��Xkm��66�g����㶘��Ø�#w:r��*j���Uۅ�a�Y݌���m��m�oQg���PY�=Vܵw@�[ p <6��-�uh!�����T[.�:��7D��!���P!��fR��*�� *U]��m�[���瀪  < < ����{��Az�U�n�[Fm��K��[F�s��U�
g�g�B�w;�l�e���A��]Tث�3�l���  c
���8�B��k иø �@2r�r���ּ1˖              �
�ЪU  �*� � 
�   �     
��ն���k�c9)�yQ��-DN�����-��޵�e�!uaKN��b-q��H�R%ˋ�HػS���gb��a@��dq�\O��xt�+�0��&��>�Qc&�m� �{;S�4��L�S��u�x�\<�Į+x@����Nt�Y��볈�{6����	�� P� mkk��c�v�P��ƶ�rm  ٶ���*�;��(��<^W�M`���k�یU5m�{Mv{c�����Ɖ�v����m}�bL`�S�B\��t��~�(g���~����3�?���;x�2m���S�'�f��Glq��q�lk�]�do���v,��a�.#9T]�^��Ǎe�m_ai�>kw�q>�����*�@�Y�`����8V�,��R�/��N����+(-l��0g�f�&j��e��l�K�;���ܾkD]w7=N�4�b����3����Z����{epv;*$VJ>~|3�����(����O���z��>��/7G,�Ǎo��Y��l�8�U�X�	�;Y7'I��r,b��`W��C.um��!K`��*��k��#��'�p���D��
������ӆ=�����U�7����k�/�kC��Z��-NH�w+��i����I�IsH��;]��S��<2{n|����P(�l��CV�#v(�5�������w�v�y�\˶�i�<>��� P��~nH�)(����XsZ�Ʋ͎�/˹i��!��J�������w�{�hYlE�����˷�۠g�{۸����!��2(ܣ�d>V
>)���݄�S��.�(@;
�v坅훧�N;P�B��f��]��U[[�ɓĚA��RX�љ��q�2}����o�Q��h�i��3�qw64_�29"	'�:L���9�p����K��XG<�\�9�@����8W�p8�!��l��fW��)����wNP�g������~<���f,��cƽ��U�Z�N�j���_!���=��3>�	8ѐp;~��a�y��ǭ#��֩
�Q�Wlk�>�x{��
r�M��4A�K���U3O�� �37cBTD��h�S	���^����,�p��v4�bԕ�[⮱b#�-U[v���)" �l�s��{��O�n��iJv�ʠ���4�f�p���4�1(J���N��ly3�N�]�Y}o���s_%L�Ȇ�q�$@����#�nn���<O;�������"Kx�%@�M9�%��;��7_*k2E�\=K�m)w���iIJM,����h8����y8���*׺�;yli,�$��;m����c-��,9�����ޒxŇ�+�&��J�d�;^���cmHL33*-�7�����+6�^֒۟j�3\����u;(Z���	�>=p�8�T���%]��6Wz��ͭ�T��5�k�#��6�
H���(�Lf�U��P�@/U����#V��/�������t洧L�uX�N��Y,��D�����?ƞ��-�AFgW?]��O�OaY���!����h�I-n�������*p��)�
�}݀��_q��y�au��㿯?��m�Jʮ����u5R���Jkm� r�pjէ�&����k��۱�tt�e^�2���h�;Wk��3=u��<m��7A�e$����Q��v�������g|e�xu��R�֮B֤�O�;=H��A�d���7�	՞�6Kag��d`�UL��������`�ֺ ��lC�ݺ���7n�@ �m  
��w\�f��Y�up�ݳpPk�Nq`�=����a��B7 f��8\4������_5"-�n���{�uخ/��=�φ��f _�8go����Z������bI��0�{�v$UؾӅ���!�j�{�`��Y;��j�����o�
C����*���w{�ƫ�t���K�0��/���iE���
����>�`h�#(ۑ�����*�21^���;��Ỗ<C�'s�2��t��D|��@`	8H)ϫ���龍��0��=@�]��8d�JY��	����S[�Ф$���2�Z�����϶1�6۵��'�(�Xΐi�qv.�:j�[vD��4�BK�w����{�w���3����c�	j&��Oq�)|�_������m��F�w��������~�W��_#(C��i��-}�Q�@��,���I}bBd)ah��Fo�Oq�:�oh��[��[��:c�&Y���h��K���M�҂6hq�,���6����	�?2l�0�w�2E@7{���RI�L����[w�C����({��I�{ʡ,�G���{Z�߱0���%���xK�-s��@���|F�s��6f�c�
�v.$�6M���݊k�[�~dΔ ��8d������.��3���6w�����s� ���M��JX~Ԯ�z�A��Q�fm���9zS~i{{�}��O�~mC��K, A���{���T�k��̸̬�+��^����;[=�Dx�޴��b&�P�b��#��-}��{�C>��DB���nx$y�����B�}����!3l�j��t�<�ƪ.�n<E���D�W�sp&0���	��D��G
%�\�`�qƫ�NN�g�5����n9]Y�K���}QUU�d���t��:43]����{�/P�R.���M"Ȼ]�|J���>����Ϛ�=Np��R#�n�m�$T��d22{�Q������jϘDV����J�i����ʢ�_req�M��$����Kh�6���?��I�e���+�Ҽ ��(��Y�Ŕ���݇�Y[
�#��}�)3������;��^���]K�V#�E�v�w`2�W�l�r@�$�Kd�n���Y�*K�Zr�1^��w�~���w$x����1_���!�y��-Mƚja�q���jwe!�s�r�֙´�c2���Um�p�z0���l׾�����	_��3��������*z��a���9��z�jky�d���7$m�T"W�e/��`La��{]�H�����o�ZgϘ�|�Z�I�#2�d
�[%���3��}v��y�]���c��o��1z�R���O��<c>��e�&ts+�h%�ak$h��?5�[�s��3N`������.��N�9���x��SOS�7S�v�$�]vڒb��!�=]�)g{Eꨶ�D[�b��7sжf���ﰍ��1Ի,잖��� ���
��T �ݍ��y�Ǘ��sJ�j��j����8���'R�^ã[9��u���9���n�ɀL�% ��؋�,��ҚN�w;�#m�#e7���1��2,t�n�=6ڗW'm�팸�hG����$PcՖ���P�&4�{���c ��=ثǅN���)]�Zw`3�ݱպ�p   6ʪ�P����M�{m�Uۡ�J�X���u��;�nV�,��vd��N�Үݑ�Fzct�8�@��8���{��Y��u�2�����<���ӕ�+ij}�N�Q����MEJ >�e�ឭG�/_����v���g�� ���	Dqص�t��FY��O�Vxg�u�gq?����pZ��"�Z�@T���]KO˰�aK�v�Y��#xf��5�᭜�1��*&���L"q7]��qS�!�♶�sHG�N��򸶖���+��S�kz� �	��t������H�l�ͭ���U�6�<��e&&N��*��dn'm;J�P��g���{��/�?.��zzȀx�Fv��Wb�\@�i�"�T]Y#�
 c���p�����s����m-?.��ae_��Y��_��"�誖��,�L�B��nP���<�����t����t��quW\��#˽hP�*��Y��-L�-�F���c^j�o7a�3U����jaˢ�O��O���#}�E���0~�s��[("m$���u�~�<���D�+��[3O�x�#�W�|��Շ�8U6L$KI?�k39R���F�ț[F��1�A�9��Y
n�zy݋��U[,�&ynrb����f3�c��^��1�b������0~��ܪ5���b���[�p�56�)�RRC<�.�g�s<�qD��_����?q��v���Et�zПq�Fq��0@`����]�)q�<Lbz�_{ޏ��8�@��}�c�8׵i�{�0�S����9
����H�e6�|?A���{���~��?x�!��f�Z�����24�Ot�(ʠ8붫cE�s��u�Sr踵�d<?D�S�3�|+��������א�	�Ά��ڂ:	�-H������c���ڢh왛���-��\pÐ�i@�B��,��Y�vi���^+<3�FI �[�`R�n�r����uvVձ��+#�k�W�oĝ��~��ϯ�oB"�l�����a���#]��q�O�W�/@i�8��C �z�����2����2?.�ܕ�i}��w]���t�z�('�A>23Q6�H��]/J���>"����Wb�\~��F��os9q��^�5"sk��(�l�rF^,r���0�#����Uܰ��Wzԭ!�jb�߾�9?c�V�w7"rD�ظ��+F<F���O.].Qt��SX�0K��kl�R��2�Z�>g�:c���x�p�T���eqӛ�$d>��v�c^k����E�m��"�e$�C��o�?4�~�wo��
1��~鶪������f5��-�0�m$�Kg`��QP��H�>����"��
�Ň�8ez�iy���65��������c�V��i[<u�?p��!�EN��~��n���zw��Eţ�a_���c�Ot�5�~݋��:���GoV�#$y��_��U7m��Z��kZW���of�O�?�-���m���[�h]�\=��bj����YyN֧#�2�����C�s;OyŢ�$"�=�v�Cֵ.F"3=98D޶�[=���]v�a�B�vۜ�2�v��PE]v�%��O<�7�])�4v3�����YPӛK{j=��g��	θ[���mtl��Ƞ�˺�]����  δ  U�}\���[�^9��6���I��ȡ��-���\�A�{.�T�@�Wc��"e�.�3�=���+�/����0�7Ҹ�]�Ӈ��a8�iQh���:��f߯��2�1�^�����`�\�i��ė4�<A�U�ӆE�0� �3s�#��0�����1��E�TF�*���B:i���A���{hp�VVFAсh���a�q�ߥZ�Ή��f�0.����#ᜡPg����G���1) Uذ�6z����6_����1�b�QJ�53�nt�4U��msMp����.�ے��GZk�-��#�{mKL��`�yjU�E#������%�H�1��k6my���#�9;S�2au�;�ќ<�.q馶j�0 �`�H
P�dQ�C��(��pia�O��G�/|��,�XF�=L��p(Jm��mh������8|5K��b�����2�1�W�T�F𸯪�C$��6�n!�9Z�O�QX��熎GFE/�l1]�����9���W-VĚ�@E9�!���|D#v�xcXE{�#=�@��k\x��T[	%�����c\�Q���'i��=�6$!�!���Wn��*�Ҕk&�7\�`*ó}߬��~���E��J���\�I\E1���ӗ��Z�O�[smm�q��Lm0��53�yǈg�G)1�de��7<4r:0󕽃 ��jR�1K�F�u�TF�1׃�B:i���A���lߞ��Ef�H��s�� %�(��L�њ �j�������4�*���VF�+��ߧ5�Sᱎ�e��#�iv��פ�{����C+7|^�`\��\���[���,6.�&:�ײ�F�[�W[��z:��3�i��m�b�v�<�R~�o����\�Aj�Ov�ͬy��s(�a��6�q��%r�k�z>��q/���k���D7Ӭ�X~���פ��:�
KNc]x�=�����F�[����5����4Vn����퐤�&Q���-�__��F�ˍcQ�{�S֨�e�y��3����"}�B/�[�M����]��5�|�?�oeZ�[t�Q�3D�_?��3GݸF��q��������e;��CQ���:��JOP,C�L�*jjU۝Z�g�ݮ�2�E8�V�Ϯ~�+���k}WY�2�1��eil3þ<C>;ك�U5m��D9�k���W���r��A�[�w�8x���Md���L0cE�l�l�#z�馚�(��pqaޜO��B\��x!��gM���o
A��l�v��4u{@���Mڗ\�F[�Z-u�����s!�|�u���lh����C<4Z�_���;�r:2)Ipdų�����|�ʄ��cj��f�����ڦ���uF�M��q]���ص;V%��;�ji��Dv;SeCa-n˹`�$Eh�ȅ�c"l!��1�d��F��q����ɇN����K)89��@�.h0��Yn.�qi#��;Ͷ��]ڳe+kdM�m�n-i��;۩v�^+r*��o5��v�x�5�2�]=�	��Z��;���7GP  l  6�={=�n�f&�6{��L;�������� s�j���yWB�u��n+=6��_����Ddou�4�ZF������)�m�
AK( K(�JA�T���k��D+��?��3�䪈���<^���Ae�!J&E�4��l΁�����0�����9=*N�W2�k���H��m�'7�y�T�#8�t�S�ȃOdou�4�ZE3��V5�Y�[$�U1QВGZ�3D�������ዠPg��{ ���>o��4@ю�D�)�lm�r/�{`{u��8��5�x�Ԗ���Ayq��\�o�ټ��6��U�F���1�b��Q������^�9�����ֽ��Nƭ�"�����Im1n�Iߏ~��v���8S]]dA���;�ȚcZE�;IP_�YL��KsFx1��+[Fh�9ׁz�u�#��i�WZUذ�6W{	?O���pd!9�q㰻��k�R2o�eq���;|�@ȳEopE�#�5�E�r�$*����q�ݓ"��J�ќ<�C��͟y�ֽw��	�E$V��mR�׮��3����m6lp�ϕs�opw�v�*��ly`Qi!��p��F���<�<��|�x�<F�FW��8l�ZG5�i��ZZ���iC[�����ʜD!��5��1�b��O�N�K�3�17���T::B�J59��֙��xg�::Js�����4�"),�{��	)I���8�F�|��R'�g��
�њ8dj�����|�<j��S�eE�W%r>k^��K�V�њ1��n���Z�{u�*k���sG`�� ��Ll�"���6�ָ��8��T�,��F����*����v�C.Ə���%�B~G��7<3�ч�	83�W�r]�Z����}X���A�A10��2"O{�A��Y����4��o �$�Gh�e���ϛǉ�$)4T���k[9N#H��\L�V3�«��c4]�\z�@�1�.|�p8�f|�1�Î\i�#ٜ g>$s/�AZ��s��GF�p"�P��n�"Ln6�{n\�-������cY�OS�dY�$��RE��8�4�jݻt8�n��;�W�a�e��ۖj�ۭ�ulh��Ut�1��1�/�b�O^�^�'j����u�6���Q�Tb��O�Ke��k�B�Uq���;|�h���#��];�h�ᖿ�X�A�PHZ+`�1��	��p�O�pb4>�Dx�#;�za�4�B��q�I��E��Anh�wA���G���tt���92Z�^DBY0E&���ל������MǨ���Df���w���~�����������O\X��U�k�v��Z�8�nq��>��ь�z����Z�9b!��[<�@������F��Nst�����
� 
�nj��iAT ��8E��EP�� �"&`Z���d:�tl�ڨ-�-��a�t�AN$0�E��51���b�F���[h�#�-'&N�Թ�w0��Ʒ��%t$� -�XMm���đ�9h�I�V�l&J���$r��ڴ���k��+��9�IN�0j���M۠���km��vyWYH:���� ��֚{=�u���L��vX�A�Yp�n6:��:lZ��,=��H˷[w,���-��պ�V���N<��ю�ڷjF�PPue���d��j簪��ۉH��ި6���C`ꃪ�T��	 $�8��u�E�6�,�z�&q��䵇�m�;�����YӸ��p<�р�-�c
��v�EC��r��X�^��I��t�½,�0;�-̛[�(������(���֐ҼX7\L������0<�چ*�z���og�yg�P��qul�|��� m<.�]���rqûYuј�9�"gո�:v���u�e��i�9�t���$ܺݜ�[=t�v����^0ck�f,۞7�3��щn��/��>>s$�7^N݄����=x[���6�6���Vy3cq�����/�۞��͐����Z��g��q��㓏= ؗ�����3e�x[[*Y�gvڮ:��  l�b pTx j�WV�uj�PlQ���N�#Ӣ��ٝЄ��N��7Lq��UU�  �[��� <    ' c���8��7�#�#�G�]p[�ɕ���)tthA1��cq
�R��+�L�Mڤ6kﾾyU{�9� P@/f�n_M{���g-T�ow��]٥��   P         U  UU   Q8�      6�    ���p��u�]ܮT��)��-+$�k(�U6�Z�
��Q�\-�Ų�K4E�ew�;$�&-��E�Z���nmQ���[�'�ƌ���v�vŹ<	�#���\�K�e��j#mq�D����(s�f7gk�g�Z�5�ȝ�ku;t�l�cu�2`�n%�^���	S� [���}Qge��1�wm�Y���`3� %��eYeyUj�5v�^�  -�� ��;):��iڴ�ok)Su��������.�b�_dbq��S7_�����.�<�F'�r}��~���2�M ��m��lA�ByFx1�i�|~�5��C�8p��s����v�1FԴ
Z;`���:�W���sZ�\�ZY�/YI�4A�t�K�3|;����N�p1dWg�/�������AN���f$�c8|�'q�����m;�BB08�nA���?.p�����I���W�M��x�ƺ�߷��0�����2X,���h��ݮ�1Gm����b�MI�X�^w�M�m9���_������@x�x1|�h�ev���@�0���^cX��G���-pP!k � F�ᣔ�>G�\��B�yۅ?�5�1J��kO�HG$�v�;#�f�C?-�"?Q���Ȳ��`�0��{�����<=Бʭ!e)m�r�4�g��O�"��������2�E������_���M6F�
��kr:[~����T� ��3�~^��(x�g�~�K��F{~��������nȹ	��^ڜ����v���P��c< [w,�.�Y[R*�#b
�����Lƣ�i�?B7w������0qG���ɿ}"��QE$
������_�mf����b��_�Cy���0�d����H岤_x�����u����@Ȳ�,���]iܣ����#q"�! V �xTmW�C;��P#�~|���vo��?27w������J��"�2H�3B��;�ԕq�����~���<S���{�~�����=�t�2~���$�A۶Y�/<�|rF�n�܎31��`�R��iWn܎�H�d�'h�����/�~C*����Wo�d��e�����A7q�,�ӑ�_~�o�S�?n��g�#�x��!kߦU�=p�ڊ#"�����T裥�U�h
��ޠ��{8��H�I�Zh��w�ee��jd]��v�=�I[�9�I`�dn71@d��_[�z��I���Q���{���ƺ�\� �b��%6x�6����Ӄ-v˳X$��Y�e[��[�G>�%�O��TB�!�~��q�x�0��U��E�M�+�8�,��QD����\I��#����|=-ѣ���7�{mۧ͛4���z}Z�Ph��% b���gָ�L��R�:�j��g@8^?�� ����Gj����{�y{ޫ`�d뤮�+�oa[,�\}�t`��wL�!l�W7��,ٹ��(퀝U��b���콲��s�XԵ@@WT���p}�F�ū��vζ�X��{u��<�]C���]�ɛl�t�B;�0wj��I[#�'�<������1�q�s[�����Սѭ���.�=v׆���<:�%���4n�a[�qvl�BO�����p��A�Sm�Ok��������vR�a �Wg�uC���  �1T� �����1 :YK����U���M�y��؍]A�G��]<�6W��R�5Q�D��n�"�Vs>.kp���g�W.Z�ɿ\
E���`��x�,��%U��6m�Yv��b��sY��>�-����+����l�zE�gs��`����j���_b��U+���(Z^W��)քv~�/�<C;��� ǧ�<G��J�yY���<X�L��i��m%�d�.Jt1���C�0xmw���e�ep1�;C���KZ�)�-�.�=���N%����2-X�TS�d�-���]��%�c<T�Anh��]ϋ�?h��󤛹i�Q���
��2|o֒�c�:��"`4�m��E�h��ï��k�b�vm� ��_L���[ ���h��Ph�0�e��nZtQ��ߪ%���ޥC��fF*`�lt��xe���P[M �m{F�?xE�'i�_���~b΀n奊8~u����wԴ�(���ibl���huۍ��`�=I�?P�2���4A���0�c&98��� eWDH����؝dx4c���Ӽ���y�Wm�%b6��iW��C�Un�R�#�'dk��u�㻚��+���o��bߌ��	���>Y�ѓL<��Ѡ��X��O������X�W�?AМe��������<�A��!����H��H��!��| �o�84~�A���ch}v��~��4c�i�?xE�L4<m�E�Q`���>Z����49�(<Y~��-N0�v��p3��*�<�ݵ�vW\�ֺ�Z�����,�bt)y�Γ*�]��o-�d�Y�63��i����3�J�c��B[����g{���7{A<�sr�
�_;������}�����8��^��ډ��a��2�4Sb)>�<�G8H��n˔�=��j��Z�B��ȣq�R(����jy�ݻZ�(��?��>~�E�'�Ҡs��4�q
�!ee�����r�c��n��w�������qXaS��a64��ChƬ�lA����1�>MG�A���y�4~�hD~����A(���"�7%sԤ����^��'�;`��q�U����v/m�}6����У>���)���>�C�(��ۣ�+��[��y���\wf�'ݔ����>��e,��A��ܣE��ޖ���Q�{��g�>�p�E4 <��1�7��t��Ch��R6��� ���b|?A�et�����ii��Z|?|t1|&�T�:?Q����]��y��֍���c��Z��+���E�'�E٢��~b�]A7r<p�ް�"�ޢ�܅$�DK.[۹��S[��Aڕj�6ⱊ��fƙPg�Mۤ�@u��:�N�p��g�t�!P�Nj�^'l-0+�E9���xw]�6�F��,9?����^]�-�K�5��	sm�q��X]c8���0�+u���I�u�nv��{b��nۭ�T �o/\�ڰ�y���V;vY��ec,�h��ݕj�9�x]׷�  Sl  6�.�;wk7Z�ӷ
��:d� 뺟.�(�(���9�B�䪪�.�q[�M$Y�ߟ�����~o������g�`��}i�G�Q�r�v����k��Fq�g,=|i6�(�1H]�ahE�?�x��;��iǴ���>bt1o�ge.���G��:1S��B���!�!m����l�����q�`�������~n�J[G�x;4x��^����`s�e�5KU��4��2׻<L�*?x���pr�E��q{��֏��F5Ҥvf�	VM-S�XI�Χ�S�a|?Q�����Y��w�E�����������?PRg��4��Nۓ`��=ks�)�;�3ڭm*�e�d媪��)90���q��h߈v��^�i��Dk�#�M����=<Fr�]�m5^?Q���\�I,V�-nJH�x��^��5�%��_`�;~����59�M�5�'��A���M[$�KHm��s� D^�8}$����}Nو��
^�1�@(�ePT߮��7��ټ��ߤZr�R}�)z��T����$��a��2���֟Uw^�}*�m�F�__4���9��r[���E�3ļ�ԲQ�r�v�v8X7g��v���H�92��XJJ�v���y�
��2�K���߿�F��g��(�Ƚ@�����c�Y��W�,���Є�L��	�v���vewŏ�|7n�B4]�������֧�?o�\,y�Fj ���mnK��_`�f��U������w��� 0<�'�aJo��a���?{_��U��TVO����>�k��C��#����ސ�!�x�'�1Ա���.�Kcd�� "�����{$�ך�/�iw�,;n�Z4����뿱�]jo����:��VH��ѺN�Tx<�5��k���R!���*��"�`+".������>�<�=�7iI��c�Sa&�z(z #��"����&ԐG2�������Gh�g����Fa23ޯ�K?��Q�a���m�Q��8WdT�N~^q������-/��C���@_��h�����ܙ@�P	b�H�Z�|K�ύd����úx���f�>w���i���z�j��b�C��i$,6�c`�p�i�����r�A{F}��e���pC/]����7����VƟ��6P#��I��;iyNy&�*7�˶%���ƥ��*����AB'm���y־����0�oY�������p�J��)g�G{|�b�.6�nH
l׈v���.<�8h�f�����?
3�~�}�����˪=������-v���f�,�ޠ���J��fY�3��[R�F���;vQ�3���Q������I��-W���f�E��NheO��ݰ�z�g09Bp!��P>��@v�V�s|~]sw��ji��9o��Q�9uv���6��=�_}��GX��Δv#��,
�T�K�W-T��z��c�BPGd�G9�\�m�M��"�V���\f�8�i.W���ij0���#��b:��e�[������w3�������;0nl�}��m[l�ȳ�mt�S�9���'p�.^�-g��Os��u^��m� k���Sv�� ��`��V�*��I�
UYK�v;�@  �eP*��ۋ�݀v���g9��q����Ѯݖ,��	:�ɓ�"���������)箌� I��q���R+��g����e/{��_y�^"�i����^"���2W��8�����O��rHM0�ՅTЊ�0ߺ�P�Xz$�\o����T��K�~j�ޙK�?����{�}tz���e��݊�� Ad���M���Y����o��ep��{L��9����?�E����Z�>ӛ���4������j��_�ȣ4�/V�A.|>u��,
�n�\v&ӖA����kvrm���z�WcYAB�6��Y)v�F�r��D*�sŝ"Z��K�?����T��3��(�FKE��cj9Q](�b���~^�k���?	�� ����«0���~�ʷ
8g��>���m��8��,��h����l��k�@�^r�vg�G��wε�33���e*v�(@˯��s}^t3����t�j���~?.����4��7���c�n�]��!�� �g.�.��?��Мg���U�Tt:l��D�P�+>�??�g�� 8 y�`q˙�:,l��uNC���۔!܊g����Y��h���秔�/�����{�9�h�π{Fn�3�~�t~�
��V����|&sz=nx�W%Q�k�{O�˨eYG��s��Vs&��p1�7�g�%w�-=S��o%#+��B؆H��Ǉ�S��Q�"��G��h��	ǭ{N��޸S�W����F�V���e^�S��]`�p�|m����4W4|���O���\�?P�c뜓lQ"rEl���K�s��3��J!��A᢫(��r���5Γq���B���m+u����X��\uD��`��-�&a��Ln��e���FݖH�7�Z�����N|����xd[?]�G1�u�\z״Y&��e����VJ�c
��Χ*9�<+����S~��qvm����N6Km�l��ձ쯚�����@���'��3��,�~ ��'���s5<��m��n�ҋ-�j~��}i6�Ke60���7z�cA����7�6������O�����AI
�	@G�M,t�k�V�u����ܝ��n9��`'�P�Xe^�Yc,���RBʭ���w��G�o�t3�{�>���Т�d�ِ��!�1����MT]��/=����|�d�!�ַ7~�OG���
�-���R��:�.����~���ˤ��#�y����_��M�ٵ�2��%$iaO�:?Q��y��J�u���?P�1󔣿g��>�p1�ə����(���n6�!֟����B�G�o�N8f�vY��x������w榑��}�[�Rs��m�k�m�E�8�*ժ��I�rp<@)p�jۢ�6:%gg��.��@��>�}�����j�1Ճ��F�c���QX�%��u���8�zu+��n8�]��t�&�d���Kb�v��u��ˢz��Щl����9:h�Lk*F�XIM�6��W��Xש�G��k�����gQ�	�%�8� ��9�u�}n  �0 R�Uv0;: $͟@]�-��έ�5�N�C�.H�U���B\�[+�說�zp��s�d.Ż�������������|��V��:�+ݨ��~����@��J��$�ϊe$�nDq��e���|~�F=��ZE�e���4��ChƺԎ����h�����1�����0��˓�9��4�PD~�4�c�>}1}�1���1�MT���[Y"|�]c��֯�AᎹ�g�~��'�Qv�I|���<�݃k�v�d������j0x~�PTp�n��?A���U�b#����h���4eC6%Qd��L*� )a"iw����O;��vJN8�R]�c���܀�=�����Z��b���4��Ba��K���4�Ǎ3wU����ۊK�����Po
+�A(b��Zh��~�f�(Wu>��N�-M�Ο���ni��K���_ͱ�<h&�#h���"��O����tQ�����x~���Ʊ�6��U+!$A+��u��Y���Yk��o��Bi��K:�柸��u_�3�k����Z)��Qd��Ο�{���j�7�L?jWI�Y:l�{�m��H�Q�[mH"�pD7mW[n��M���ŷ�U�ۍC-Ӳ��x�݊U�rE�&wOt�+��ߛ�s��̣�fA�[�]�����U����D�x�G&��Ɉ�1���ْ��İ�ڵ����m���?3������{���V���q���\��֜?W���:D=���׍,��r?�N<�8|"�q<m��6�,��Ч����\���E���+2�.��0�i����ﭣǶ��u"���I����1��N?
�ϰˏ�-�cc�d��6H	�p��[֥��kq�؝�j8�ٝ�`�2�p\T�m%�()]��d��3���Y�����ۉЇa�0����J�C:՝�epe2���j��4F��&ڣ��q]���ڮ�2�@�G@��j<<?O��\!0A'M��ͣ��<.�3_
37�����GARQ��c�y��,<@ z^d�i�
L�+L#M�Ӭ�0��imi��e��p��F�p�o��χM&T	L�x�)��"���_R�m�!����`S�ϗlU��x)4�R�0YnV�A՜�q��n}� Z9^93��j�Y8�m��Ze[m5�M�j;V�irG���XPQ�[�_
34zA�Ej���T�gL#�޸؉(�2h�bm�b�����ͦ߆g�ɏ8Ç�-��C�1t] Șp�C��9^0�e��Se+{���!n���o٤��C�Qb B�^$�h7/z:Ń�>�ap��4���|~�����(�d�FL�%~e�z��pc����7���{�<g�>}�柚������ � �/�d	?��� @����@���$"�BpaĐ�@� |�� O�$ H{��y���� � ����@�?���g�����@ @=����������G�� @�H���  �@�HI�I!?�I$I�����hx�g���� C�H �?�����@ @9�����@�{��̄����  ��0������4�  �@�@�?��N @ @?���oL����i���?ρ�������-`@ @<��������)��>�$ ��/�0( �� H ��0�/�        ȃ@}A@�            ��     P
@        �	 ��Ԋ�P(              � � � J�P  �Ȅyꪮw���s�^�=��Uݺ�U�"�{��qU3��C����:��Ȃ]�UM�ꪭ۪�  {�@:�� hN�A, �`h<� ��M��w�6R�n�<������,��$۝)zˌ�l�.���VZ��שA�n�Y_�� T��  !K޾Lm�����{�[��m���o{[Zj��P+�"	w{j���R������ڪ���Զy�!�Z�{������}�W�W���U�����^|T�]�U]�9O���S���W�y��U�!]ʧ�������޲����m������
� �  UR	w^�U�w=i=뺕.�^���z���	�yx�{r�7����oz�{j�"
���[��U������;����T�����z�����5�n��U绋���b�8zK;��^��C�wJ��U_}��O�� |  � �  " ��F�q�T���)�W����{ۋ���� �{իo=�y�ouv<v��׽�^���!yީk��{k{۩ﻇ��u�>�Q�<B	y�V���1���Cծ�w���w��S{�Dw�X��n�6���z�=�w���� < ��  	@�����Q�x�ٵ\�z���N;7<Dހ���;���Uw���[�J����ĭ��z���U���W�w���i����[���Q��z�n{��s�Okx����z�OB��{��ʫ��oQ��� ���UR�& �a�~!6�*��   �~�UJ�CzB "{RQ�J�   ���TLT�Q�  &��$z���i��=����'�������{���h�y�=�� @��d3��!B�BB B~��	� @��X���$ ��	0$	���E?��`,��E"$��P
�(�*ȱ��AH�,J��`�����D"ȉ@PPO�)���� (ڊ�%h�#"ȱAUJ���TEBJ�(��R������T���+�T�
��D���d�R,"�Y"!Fڀ���QP�*��F%��"Ȃ(���R
�E$�)"�TX�* �D��Y� ���"��U��X�R1H��E�,��[D�$T���F��AZ���*���E����H���
`�#U#(��Z�����eaD-�E�
�E�)�Tb"X1��Ecm!+ ����$��+�!��?�8�4��2�Y�TCI��A�jm
�J$�!�բ��J���`q!̰o�8ب�B�,q�.˨�8�����ҫI��
�̠8�R
CĆ�,�M2͵d��A�T������Y�SS�3i��l�1Qh�*"z�R��'<���]0��ŋ�s,�8�X
�F���Ch}�|�E��ȺMf�

P�Lg�M"�L1YP����P���5�2��@�i��c��C�4$�AHx���4AM$8�d�)7l���Z3HS-�*�Ax�E|`\��@�*OY)����qm�Ć���Y�>�*aR5h��)y�uJ��%��T=H)Hq!]�d��%J�RH(�U|d��DUlHm!��x���UbDգ}l4�(��7).P*CԆ3Ԝa�uh�+$8��4�`��YlEM�>���hX9 �%M�)��Y"ũ:F+Ƣ��H���*q!�¡A ����-Kb��ejT�-����PiX�Hi*(m���R!�{JɌ5��V�ef'��DDU�Y�`c�(z�L��L����CĆ�$8ɉ��8�I�Ҙ6��a����
�Ć��Y4�%$R����ԬQ��11F9JȪ���KV��"��1H,RT��R)���b T�HV���PXq���P�
�\aP����]4�RIQ��,b ���Y �QE�(���b �����(H��� P� EQdY@�DdU�XE�XVT��T�`��B�H,"�(EX��%V�dY
�4��!��:c�[��sVc��#�/����e,r�x�]X���\����ΙiW�0��z���5����Z��ks�oVWz����n��H����ͦ�n�����}���/�]�2��Ԣԭ�+5K���*^�t�V�[Y"��xi*��6���Ycb�;m�t��t���k�!��x+V��4죚��8<������X/m�
+������?3T)�gCdj�����4	ݭ�+�ߗ��^��I��C�4�6�0�A����u$���=���2��������5[�d���LI����$�G��6K�W~�Myz����>���8����xi�I*,^���t�����߰^���T��ZW��/W�4n��Хy�W=��h{b�+la؂i�ﮞ_А�Ԉ��2��0�N){t.*8�2��a�^�7pr��9\E���E1@r$��n,��U)��I(��BײP7 ��Q�Yx�jz�Z'Z��b��i}�.7VR9L�-���TQz�	� _
H�?	�}(VM�bd�s,M��ɗ�[�t��Ba�I	����T|tx������p��;�QQ%x�諩�값2��:�ć��%��_�rh�4Q�`��ۮ�i8h��} ����Ml�<��>�Y�1"V[�"��6��no�^��i+��P�x�,RW��5��h�E��ܘ:�̻V���Z����~��o�_R(����Z�]�|�4�Pg����E�U>��TY�$���4M�J�Os.�>��F,8�GIT�G�(=�U=.��N/W���l1�x!�R�^�Vj�Sʭ:��w�H����X�Z�@�A�J�s��}��s�J�RM	*A@���A�R�R!R,d�$1��Ve�-Hi1����4��ճ�6s\9<Hi �6�ąH{�C�
�R
B�E(UR�D1��ean��QAE �(Z�""��IY�bE!��<@�$�m!��5��H6�L�a4�IY�K�����0�J�&	� b9�c&�*[Lܹ�(�&&]�ּ��vdC7lDJخh(k(ٜʖ��{��aRHo��!ǂm*`��dM:ƅ5��B��E�3)���fZ/5LQ��3(S-\Bեa��kP�s)�l���EƊ�9��hWyQ%Jaje�<��2颹*�Q.�̹B����a����\y����2�ڢ�2�SIU&5���n�Qf��Ab[ ���EU�CUDqY+ETD�"�a�7��PP��+4�ی4�eI���E�.��dwaǄ�-!��$*C
B�*B���ͤ����J�)7���RH)!R ��HoT�$*B���R
AHWH7z�AR!�
CYH)!��$�HT��R��AM$4�4�\�&�
Cb!���d�@�JZ�W�ٚ�
�
T�1�CI$�+%Z�Q2¢�\T��V)�6�Ă��AHT�� ���Rn��UH[HT�HT�H)!�B�����P�$�RI1�2"**E�$�PY * �H�IY	X�XDT�R�Z���n��$�ke`�Tb�%�*Q��#(ʒ��R�`���ۡ`iU�	B�dQT�<I+Ci%`H���Q"���d6��`�h�YI�T���QBHLI X���a]��-�b�E��$P�<I'$6��s�4�)fe�J\`
Ci���$6�R��C�!�R
CH)$8ʎ7XS%d*CQeHbB����
ɉ�Y<��v��P�$��6�ąHbCԆ�H|��!�Ԇ�$=Hm!Ă��CI�/���3�����$�0 La�  V,�R�,!
�$% �Y�P�1�@Z�ʪ� ��D� Z6��ҖV �%d�+`�S-RI U�������[#Z�TDX����(��Eb�`�B�����J�"�,�*��
�P�� YhQeB��I��x���,��&���
&>!�1�J�*��w��n쪕�J�I�-5-Rӌ+%�Vi�Py�1���M�R��-iS-Tʾe���WG�<��&03)%��y�O<���y�x�;߸�c�=q���⌬(����h�8�XV?e�M���C�E<J(��Ȭ���2���U=̋�%�\��*a1 ��S-UY�����-,Qw� kAC�ppH���=��{��su<
�X��#�����|֦�v��d�HTSA}��e�̾�0�XR]d�:HT�� a$7�!�����PPi
C��Y���QWĬe�֡��v��*�z'����)���c�*O-���Xc
�V��x͉��Ar���B	�]�Gt�љi�9���55f$<Lt�iaP�rəX��*��W���cPY�TP�!�����4�D�Z1S�(�1�������:t��NEZ�C���r�Hm!Ă���l1
�[��0ޒ�޼�M�1���a��գ���
y���%w��@�����(�b�d<Hx�R$*VT�aR�C�$<f�0�<Hhq�l1
�_�s�1')���aX�%T^"fWS��<M��5�^o[4�+�%6�������ɤ-��
�V1���*C��M�H�Td�C�3L�����$8��i�����!�6�$���@��Af0/�FO�<D_�����&�`�6�H��_2�5FGvc�x��&���QDYF%�@$e���3#�U��xb"��m����Hm�q4ؙh�.Uq�*�B�V�#`��(WY~hET@PP��L��S����N����^��V�'=�����s ���5�H2��W����Tک�[� P2d�	����_*�r��
�֪ق��$Ԙ�8��n6ys��.#�չc1��{W 煍:��g-�h���m�X3��\]�����@���ɞC[�f�q�ۖ�eD�q�1mfvCƎ�����m�ћ'l�K�������v5j�y����l����[�������n0Ӟ�$[�˭7��뉝������s���ci��V&vc�X���&K��!��x8���Mkka��kҴ+�mf41�ұ�tm�3K���;�tr��ŮB�{\�:x8L�[Q�eƆ���n�ŭ�f��n�;sb�r���d��\n�u���U]���nq�6��`�@�9� {*���1���2��%��S�L��	6�)�����t��:�l�r��슛�W�����Qg��f���wR[� �
6��rcV�t�B�p�V���-����r�L�qt���n�&6���c�+<
<�ax��j��\S��%ͰCq��琓J�)��v�t���suCi�v���z�2�=�V��˚���;npv�m�\s�e0=)�e-��\��֧msl��q���{t���I���g�.z�����;�mc)�ɻ!8kZ	rSc9��N��;]i�wg*[f����q�lQ0n2iR+��_>ڕ�.�s]�d�N�9�S�\�{�C��l'��t�z,�0o+�g��kjS �;�v�=�ƶ[t�Ak����o�9ȶ98���`'��{n(v�v�ڸ���N ��A��dr�	mfˮɷh�[�E\�!�v�`=m��k"��ڙx���� �&��pe��*�6�ɬ����J��p�yxwcaݝ{y�z���>�T
���m�Uw   U ��U��TU
�ʹ�ڪ��T6� *������`Q�l� �U
�l׌��l�8�  *� �*��@UU��QUT*��eUV3mT l ���*�,� `P�A����+mN��mT�d *�  
� *�mZ���`C��*����U� m�@mP@.�� �Um��*�UK(UU�����ڶ�b��`�W����P����dv5V��UQw�
�Ue@�
�
����˺�@�l�6�R�ntE��@)�PY� 
��W���P�
�+b��     T��U�
�U*�@U �U6 Ȫ��d �K.ݠ-�m�KѲ�A��  � ��0  �   UR�l� C�l���u�;�*�3ql�T�� *�P U �*�J��*�    `T
�    ��j�̢�ݕ�)��Pw   �Ncl   ��U	�nM�����Puk)TU �@T�O������   *��T +(�<V�ڪTR���@T��P�AT     �T6z�+��WsWm P   *�U        ��J�d U *���     	� T   ST*��+*�
�       �VeU  f�ͦ�l��EP     
��  
��*� U PP     ڡT*� S` Ud � U �T�  *�� @U*T � P   R�
�P��ب   `Qf�
�@     jU����*���\la�uJ��M̅v[����s�:�X���vh���zI_.k�����P�[%d��&l��;\d��N��f��U@�UwE��l�vJ�׶���`�i ��y,]@�i�j*�n���wj��`����T U*�@  �{����@ &�ϕ�mgD�	�*��B��A�����T0�VZyy�S[r�f2�]���aϑZ�&�q��:�*�;�e^�  ]P�&����YWe��o[���9n�<����J�`�M� m=9�̬`  8Ca���Ԧ�]�  'V�#��ۚ��*�1�ȭ^�f]=AN~G���[J
�D����mڝ��*x6dSKԪ��̶�W�5�s���}� �zb��-�����lTl �w^��-��PU v� �� P   P*  UU�U +*�<*�m2�l�gd������.�U Tڀ�&����V)C8]�u�
��
����g�k&M��b���S��0��A�S*AL�֥�P��jj����SZ]��D����|�v1DC�`t�a���z��8����Kg���@2���h+��ѵUUR�[��Um�m��oe �E[Ume�u~S.��U� �����en�*��Y�*�l��7v�4���u�ˍ��Y��U�N-vp�i|�v5��d~EȠ ��Z��dW`�������Ō����UR��صw)@vL��e�+mA���R�Ij���ڧE��g��ѓ.6�ܡq�gT�!�a���t����d^8�k���'WA�l���;!�r��v'�&*^�����۝�`�v��A�j�h���6ڞz�x�qPPT� W@[v^Jr����=5�4��6�5¹Nz�Nj����pfH.�4Y�ny�rv-��rͶ�&��-%1�C��Ġ���)me������s�m<�(J@�Aģ�� �69��n(qD�Im�ѓt��sźު�U,���R���LlJ��UTUJŸ�ܚ�Ȥ�=��SE���h-��%[�Cn�U�Hl ���A����̼�7(�����"�O%�B̩ �@m�{p*l� 
�ܯwwk���6�<ж��  
���]�ڇPJ�ű��1y3��w{z��  T<�ߺ(��   *�w�w ���   �  � P�׶[� �*��R�S�5=!��  m��H�z�UT  ��   6��  
���k�U���  +(���b   |    
������׹q�?w������  m� YB�d      
�    @*T*�m��p�          �|  +*��ʼ����UU VV�l� U@  *� ��  U@����*�� � p��@�@cnR��ͭ�� *�   ̧��;����6���f]�@fF���jTֆ����I7(
K���wc��(              Pn�l          l            U�                   U@ *�  U  z����Um݀  *���ج�P��               {�            T        � �                      *���@  � ��    \ʕC��     *U 7��{ ��T+�C�)�TU�m�t�<wU̞��*� 6�P��    �>T           �      �  Uf��  UP
���[� *��q�� T�            ��p�ͳ���
�         �>                  
����                        
�6�  e        UAT @  ��                                 ��                                    >�  UT   P   *T�                       Wt      m�   ��         U
�^�u�P ��   5��ʝ�� �T    
�W�     *��P  @       �TC�C�;����P� 
�  T ��[{@-��¥UV�d*� �VتإP� /f6�e  �G7����z�U�����8[.8����m��T  Ws�n�UP�                   T �     
� l�=���v�Ψ*� UU 6�T��]smJ��j�   lR����V��m�O8      T
�    �-�cl
�Rp�P      [         d
�� U T�
�l*��Cl�U�Seޜ �pu�������$��! I��$ M?�	���@���̸7��vxYYe�e�Űci�zd�E{q�y�^M�5��pK������P���lr۱����u<n�s�#7I�Tه.�6�VA;c����t��K[�G����ӹÓ2k$b�q����6P::'=v6#�h�!��������a;(:BA̧.^�k8�s%�[FK��,�� ��0z�r��yG=��鶅PVP *�@�VQs["�*+%� WuUP�������*��mbj�M�vڽ@�P�j��Sd U*�e�V�^u]�bp� ������R�@U ]՚�P-�k�Tw ��PPm�液 )��� `  *��h� ضm�    @-��UEP��*T  ��Z�x�2;�sWf.����6�y�x�*
���V0VP���^ɻx��W�I���S;U�B�)YF�-����#��K�c#c@u	T�M�@ �l�.³�g����<.[����輝���/\��R�Cn*MN��誶�Ά'l���T�4���j+H�!�nŔ�Cm���̰A��t g�,k�y�v�vZ�s��xGR�̠d� ���%U�����\{��n�[۹�D;�j��2�T��U\� �wu��PUlPc
�+�; �  �T� U{2�fEUP �� [`-ݕ�ض��u�@       `   �mn��Qs  �         m�� ��Sg�*�(��)�U    J���mJ�  �Kd @   ��   �P U�             
�TU� p  � �' u`��  �   
�.��P� ER�w{���8ʂ�l�    ;u[e�i�l[:  z�U@
�   Uk34h�b�`B�����q��a9�|uN{t����m�8�q�2Yv�ݍڞ�U!*	5)*�p�)c;^%\`�kj�m�`�U \%Cu����[���@�)�sT��2ZvR�5�`����������Б�ꮷ��.Bʵ��R�wm۔�l�J�eUPͨA�EUP� �����ح��Usm�� =�m������zw]' q��2�Wvy�<�q�e���aE����+��e�vɻ�%Y�U��k��Z���,n���h#��)�ύZ��(~���4(@Pj��Mj�ܹy����٩��z �aǥB̈x�j���v\�mZW�2
��m�{q�������~'&��l6�~�5)n����)j������d�#X"�YL���_�q��B̈Y֖!�Q��	7��B���-OQ�����s���l��V�~�^2����a�?CgI���ՄSϺ�����\7dH6�-@U�KK�v眛�����iZMEԶ��U@4�$���sX
%T�߿��}��{�Y��f�����C6�;�ڇ顩H�t��|��6�%�n�uD*UJ�����l{W�V��P�"Ŵ�����F���r!�_,Cb�kʏ��R��E?��ϻ͙�~�����+�Z���<è~�ΓQ1�Z���ڄ���}N�i&Cw;�C*�ת��F$�P�_-^9�?7�:n��7����{3S�O�A	�?��b�'f����LR�\"�>:\���!�1T4dC�^iu����G!D����B�;�nn[_�[7�����:�e�UBjU��c"�;��%�A++uW"���-OSц���%��B0��+L#b�31�ZE�8hm�R��Z4��҆s������w�rg>�uת���"�|��mB�4aɜ9w%�{��d 
L�_��&h�M)H�dl_SQ��Y��QTl_.ߦw���&�&ow�|e!r6��x�������9���N�����Ŀ�-#2��ؾ;+%�TSj���L;�,����ؾQaǠ�Y�7�]G��C�y'�_-BL���ɫD�U�6V���ƗF�۷n�3�E@҃Kd 
�W�U�v�g�i'T��RuT!��jx���iwE)H�dl_SQ��Y��[�6/�_L��ٛ��.5� �Ʒ\����ؗ����lؕ�w�_+[�153�xgu���73�6��?\aYa�6/�3u�YӄBn1�|��)�
��#|��^�D>7��`n�T�U2ꩥA%p�����K4!������iwh�H�Dl_S�Zw���\d��2�-UH.\�o����=��#8Fb�K�\TD6n�U�2����=LB��L���W;q����c��J�X�j��N��1����ͭ����wUU ��(-r�\�����~�����Ei�l_)0�H����cb�E�Q�q�'&s�N�)�$,V?o�s!�܈�ER�j���,CF#����j�f�9�W'f�s�������T
i���*�E�>5@����l7����3�^B�!�p�����V���5�A-RI���b0��lK�Z�0�(�0����it���l_.�L��۔��P*F���rg�\�G��C���B.��Un��b0�v=�:�uy3S/gorUV�A�p:�m������㐳>�.�k��eM��lJ  W3m�ٹ�N�t����e����
�� @����&�g)lk�V������j�iw�Fx�cY�ۙ���ORv�{vX����;:M��@��ª姀m����R����N l �R�l pAT  �ھ�U���P	$Tc��WQsP1�jH#!*�V3�B��r��z�l2��UJ�
���Ԩ5)��U�1��N�*��7Vl#O�K�����E�6��Zh���/!qQ�^���T�-S8�j�ܨ����:��^<L�+��]�����c��:p�(JuT��e��D�Ll_(��{BΑ�B�?�T"��p�����IO*ن�U�8�zڬV\hۯ�W�59�c`äz/�bnl!��l�hH���{{w^Frf�~���
��~��pkrD4v���e���S��4a�%�/�:Fe�"�Ca.�i"JmUJR6��k�k[�0-�nc;��#ad&���VUv[j� �c����S�"Μ"q���l��BΑ�B�?��!��)�"�}�w"�I2�&�[n���S��4a�<�J���Y��3�"�����(��$_C�m�I;Ul����#93{��L�&t��w�_Yا��h�dK�b_�t����tY$�@-P+�������L�p�:p��6/���:F�z~�������D�2
�(����b��R�ч�5<j�V��;���a�6/��-��Y�� ����L�Sٹ�j�,	�jڰ`����K)!n�l�@4� 7ymS�;���U6�'A����:�gH�^1y����͉[�p����LCF"J��ֲ1���Uu���7;ܼ������B�gN�����ȧ�*t�������5I'M���dXD>;y2��.�����Ȇ�8G�����KH��1�����v�������ht��,��e�6/�XF��kM�#1z/qYٱ+|���V����n�:5M$�Tꘆ�6F���T��2��|�;��,��!�ؾQa
����6]s�L�գR+�YT��8[n�2�B����@6�[/pت��)"��K-���#�B��}�Y���e;�]/�/^�)p���_�W�58v��%m�"F�c\E�٩���p�N�t��U�,#a�u�Α������lǙ�KM�4��IPJ��#-|�lS��4a�6�ؖ-#�i�lA@�(U�,��ZhED�E4��M�A�؂�ȧ�T,��.�PȨ�|v�e+�] �z�)L�hù�;ߖ#��,RH,u�W�4�����H�A�&��F������
,#a�u�Α����
5L �N���+Uy��]	���Q-�� !�a�R�UJ��J��i�HJʪAf�u3�R�ˎ�H,[�1l��Ve�KH��r�vg;r}�ޡ����7���t���lAEdS�:F���2*"�S�.�X��m���M&�[��Y��tg�Rеx�>�q�a�6!Ni�"Οj�Cb
,"U�n� 
�m"Mr3�7��ߦ��!�r���h+[�G+ki��wjI"�
�P��
l:�!ӄBn1�|��*��\,��.�W���~|rc��ܤ�@�ͭ���a�������'.�#H��3�KS��JD�ʲ�FҡPHH�J����ko]�
��  *���=�<�;�q��JY��
�R��dR���k�4k�Af�7l�;c�3���@Zu*L�c#u�P��@;�aʭ�7�F�UT �� -�U �  l 
��������wO�mW�ll�w6mn9*�BQ��7R��Y�L�ѢNG�k?7Z�U ٶ�h�k���U ���3M�wy����p�CSƯ�kH��5*���:rwT����K�0(6�W(����|�q�m�I�r��{�h�_+Zd�P��6G�{2�V�,	(��:�[ɛ��^F��������|b�*��_a93�ޒd�_��fv}6g������[�1p�CSƯ�k�5>�z�;53����p��9?*kJ&�:N�t��U�,#j,U���������lܭ�FZ�Z��-�?Ga�ޭS1J���V�:�7@/nsnGaj�j��`�U���Ra^Si�RN��h�dm�/�KH� Za�3l*�C���cb�K򆱖�FF�:q�4�o�~�5߶��;_^���4a�=O���"ϋ���9)@��h�٩����Ǥ�E�>2c����ڋi��f/E�����G>�_�����J�j&�FZ�Zا��h�dm�o�KH� Zd�v����+ٝ��^�5D�2U�ԳGj����^��K˪��<�/vu��u�E� �d@�imJl-T�됺�����}�eݦd 
����E��c%�T��3����kk��v!t��U��Y�QV�;3s���8V\(�Y����gۗ�0��L��h�6�د�"��_�&r~7�)$�И�U#2���;���z��<������I (Y  �`�$� ,���@$P�Y$�!E$$H�"�����,�� � T�
���H���`
��� (�`���� H
21�` ��X� �P�� A`
@b)$R=I�'�&��4l'�	ua?Oi���;浹ćm �+���*C�}�m�+sB���k-�4c�:�Xm�d��!�����l&�R� ��
���z7
��*C��S�
�`�k{�s�� �h��+'���湫�
u�X,��1 ����3-{�q�s5����0��d�*C�H)�a�s�PY7�1 ����
�Ϸ�ss��AO+��wf$>�w˧d�a���T�- ����h�X,�VbA���a�=7�:���IA�L�+V�[l��n�
��$�ڠ��+(�m�f�ۗg�k2浬���>eHn���,�㷎jm ��
u���d� �9��>@�%��H;i;��t�a��l�� �+z��7��Y�m ����+&��=˭$5	��+G�~n�}�mߛ���K嘐��/;�vAN�VaY>eHyi=�o.��Ad��� ����;��n��T�- ��	J������~B�~\�m��鶵u��fk5�]����&�B{��n�>Bi��	�;��}�I� ��������_"� T��wf$>�w˧d�a���T�- �uϻ����N��u�kZ��M�Ă�uf/͂� V�a����;i>@���a�:�~��x��=^w5 ��
�)/ٌ6�)�z��q'XT2�[ �'{�Nfyn�:�V��e���n
>�M���zü����M�#�A���/n����$�a=��n�G)��I箾�P���a=BO�����	Nが�R@�֥V��{C������o< 0U*�\w[mݡR�g��;��{�~����{����@�����6E>`VA@�Y����)�������0�ed>�AO'��5
��ٌ���)���
��}�9��AO9`c �g,�~��ܖ��0*A���~��g�+�{i[ ��n���.n�d� ��
��,1�VC��w$�A@Κ�sSl���)�I�
��*A:s���В��k��w�+�h�3F��f)�kF�a4�|�o�$�w�w	�i&j�u�z�}���f�>a7�^Ry��5��I��������}�����2͐S�I����r��kM��]]c�֍ u���
}ۊ�G{��p���)�I�
��+!�f�]�)�ld��>6AO�������@�+!��
y偉=�{�Tv�d6ma��yϴ�=�ZP)����w���n��w,9���}�;{aRm�@�+!�d��Ӻ��A@�ٌ��d��Rw�� |��v�>큉Κ���h)�I�
��+!��q^�5F�j/fn9�� ͤur[A��쬻'q�	�c����*�
���]����@H	�FR�����A�v     UtxjL��[!kE�Us+Ur�9��F^Kjb�3��UK��=m�e��mnհ 2Gu�U6�lv��2w�sqeUP��Q� Y�T�  � �*��Up��W�/��m�S�@<����C,j��P��W9��1���:U�
����� V۫R���z��<n�ֵ��s/��&2
~Y����)�{��p8��*�Y��S����y����l�A�d����@����f���S��1"�@�,�C�}^�����
��VC�d�\��t\�.�K�.f���]��E������)�I�����@�+!�d��$X(�^�����S�
���VC7�tw �ݰ1"�@�ٌ|�u癣�ߞr��{���턲�Aj3_z��������9#�l�^6gv�<���,H�.�{Q��?5�׽3>�v�>큉
����չ�2���U�.9��A�d�R| x��'Nw5 �ݰ1"�@�ٌ���)�o���ĝaP8��}l����ď;���;f2� �X'����k9ϭ��I��3�:JI|5��Q�8��r
u�Rm�@�+!�
{ײ�$X(�1�~l��0*O>w���*YY[ �ݰ1"�d޺��78�z�
q���d��!�s]�S��1��d�ى� ��}��g�W5*�1"pKTOn�m���@����A��wB岠 ٭쳼��k.�����f:ї`q��+&�RZAO<�c������ى� �P+0��׾t��C��S�P1��d�Y������:�Xm�d�*C��S�N��X,��1 ��
|�X?}���Z�n��)�i����AO�@��;��H?4��@�>aY<eH'Nw4AO�@��;f$4����|Ѱ8ì+'RZAN{@�7���Ϭă��S�
���|���2��残u�̺�k78���
st`�Y3�1!�>/vc�
u��
��T���S޽� ��ɚ�� ��������+'YR���v�ċ;��]nI��'Ϯ��/1֮i6�m��m��r��WS�8�zi���y#�eo�frG�� �n.=��O[5o�ݳ��жr6�# $���Avم${�q.H�l�_
���$b^H�Ό���g
=�X�K�D�=�XW��S���)�H�p2���V�+u�����[��+oh8J��`[fQKn(����y#�v��dH�H/��@��6jGR���ߖk"�vx���*4��~'�n6�r�u�]�������Y|��F_/+�&$}����+9���ĳ�ng$}m����h$��F$i/�,i�1#����$HH�s2 �dک�(����;lܰ���� �(0�[UC0ĉ��ɻ��ԋ(�G�H��7m��܈��lč�N$}��L����[9y�^�~$@e��m##d��Ǳ�(�F$OvU�fF�$|Q��~y�$LH�6g?�C��g��d*RɊ�U��V�[%%��;�/V�=[6��SmS¨w6/˖�:�YIZ%�Eצ˝�N��r��&���3y�$HH��䌍���L�����JU�nT����P�_iF�q��i�Uk��"<l���^�M}�ר��4E��:��mD\@UJd&Mzdm��n����rjMTdl�z��<��Hĉ�u�Y��A�{�{՘bDĎcqƗ�,�B3L�v���W}��QS|��:�:���]�N�aF$m�Ԍ�I>�&d��ڪ�7*����LH�^�\�LH�=��jDč�ɻ�V�YGR8���VdH�6Iį��ﵻ��c]C`���\����6�g�u�g'%*��U@�f�Wvw�$��Z�5;lm�vϹ'ɲKH��䏟��t���0�]7��<Q��H��\�$ď�5|�6��KY /�Gz���N�>�N��>�j"aF�޹�����Iv��;U&m.K2ZvIvم
2rm��X��p׭ճ�	'���Z��OK"^H��Vg6I|��X�1,J[7Гz���f�~���"Ƹb+m6�[ւ����E�M=#֢�B$Q��*Z��0�y�i|��gm峾��䊖����S�K�ϊ0]��1/%;��禳�8Q<Qĳ�k�䏱�K��1ڨ�<Q�}n��n��e��	�0��37Da�[�Uɋyy�L���ӿI����UPK*�;�h	9Ұq*�V�m��� *��*1m����U�ٽ��s׾���ݻxi`U*s�]s���le���Q�ZC���T˲�rMK�7c��� �m�PU*7a�l��J�
�p   �   � �J�T -�ݳ`�]����X���|4DE�TkY��ւ�.I	bIy+:��J���+�5�Xv��C����?x�|Q��7����%�aݞ(�(ļ�|r�9�K��.�8���7�u���-Z�چ�������Ö�/�r#�
�⍥�y#�{�TH.�0�aFm��o�Č��9�Ymkq��K����nY�yn���9�A|�Ҍ�s=�pļ�H�3��+9�e�K:�㖇���`a�U\"����5�zf���z��!�Y�Z4ʄ9C\8��H��rٿi�L��nY�}��Fɕ�	BBQ����(��l������(�Q�[�OR̉[d�����3d�F�伬�w�"ɐBvY;,�0�G!qĚ�Z�TZ�۞��
۷=���F��4�J� 
�N���I�S$��|�$g6H7\{�<Q8Q�j]��+3�$͟e�Y죆%�D���<^\w���OK7i�zI9�@PIU<�H�$��c�U�"�2RBՑE�CL�C�W
{P�C��~����Y�ő@n&.��C�7)��ɳ�ZQ#��r���6h�aG�nM�<ȑ�l�_�܈��l�(�\���}r}�$1�8�B���{�%FaD�FK�o�Č���K�sNbZ�c�
����g�|{(����9�Ok��fr���UU����sf�'�8�u���H�$��c�Q�x�irX����Avم
=������I��;wf�h0l�UR�<X:73!S��s��cP m���2�rBKL*d)�zY>�ĺ���W�\�A˘xQ�^f����D��d���\l�D����,ȑ�	2��	=T��*�YqMIJ:�K�S~M�<�
&g��j\H˘H:�T�p҉ҌK�^fд���Y�o�gņP�%* V|g�%ĢG�R��.�����ͤe�<S��TG�l��P�Ɛ�4�lF��)�Q!�Dl_(�CH�Yű��!�\r�g�{�W3�Ü{�ti1j��h	`��}w�w/�2�tzz���:�f#�|�Wp�=3��_D�hV*��ԭh���j�D8-���ͷCV�� �R��Uwm�#��Q�����s���Ϧq����ψ�T�PdB�(�G5|�z�~��L�f|w�!,=(6�Rԅ�_�!�ov��(]�R[K�1Ek���wW�ﭩ`�UɅ^�s8�n�.������qW��ZG���Q �l��A3�.�ı#��Ao�6ߒ���B�R�ŃM�zY2I>������BL�l��]���0�IjG���k����(�H&�O<�H�$����4�m���H�*6OI�#%��d�����\��� ��aݞ(�(��8w�Y�� �l�FU�+̀�i��ʒѪM�j����n�irgu��x�;%�UUUJ���� G<@Y�&�O	�M%��d���/�ٲ��33��dH��$���͓�y,H�~�&A	�d�����l�;R�F��AW��>p҉�D��w/fsd���⌾��p�IjG���/�;�MK'��<���߂Z��"������L�C�3ܬԞ�I�ui�hu� �l�D�G���$g0��X�^���s���$FCpm,Ʊ����8�������+ڳP�^�[�k��`<�2-B��
�*!P!l˯Թɜ��u垚��_�)��D"��vтU�p�89_���[BBC��@$P�U $�	 ��H������2)$P��,�Ed�*��"��
�`,�$Y $ �) ���IE!$��a R�E�(N����i��[�cuJ��0 �hFٔ{�uڹ��0l/Z�g��r�����$�rP83I>�i�S��v�.��p������1�0�봉���Q�x��X�;��Z�:`d3��n���:rg/F��፲��Of9��κ�؃�V[����;oX�%uZ���m���M�F�zx4�0�aet�0��~k�Ͱ�UU@*�TT� w*��PU6�T��*YEꂨ�Tw  m������zq
����Y��v6�b��R�2�˸���Ul�@  6�@VڀM�w d�Tx������@*
�� )��  QT � m��  ���    
� 
�� 
�� 6�@���߽ok/Wl�����p�$�+ʵ��{<� UBNC!�V�
�ZMV�I��t�vwJ�kh���vh
U��v.sӶ��l� *��*�  �lR淲�5mm�W��[��v��Cn�.6��4���t�uU��7c.D!�u�� yv��Z����5���� s �c+�6+s�0�m�hwv�][[Vp<p��9�F�-�٠v��i�']�vNs�ou8�`�-��.i]��ϻ�UQ�w5��P*��Sa^� ��n��8�P ���   �M��  �P�U�/Q�k��l��s�X0  �        � 
���}T            R� �m�v�l��ݲ�*�    F06�VR�  \�      x    e  m�       U �|       *� w  
� .` � ���� Q��
���4����d���P6d    �> �T
�J�V߰  T�d   J�-�z������s�)�{F���nB.��z붞lr�Q�U��=|��]�� +m,�6�m����]���ĩW�P��lm��w`a� 
�n�mܪ��+w /���\�D�*ɴ��
>��֣Y�sw'���U��.%�͌H�	]�B"��S``w\ƺ��6��6)�UU
���e 6� ;�  6� w E�T)�m{��[l�Ͱ-��74��![-��K:]�v,���0�de��Jb��[[yV�l�~�6�`��jf��jY?ĳ5���Mꎞ5��=�N���.� ��>(�}��s�&K��_RI��ERFUEf(�IĈ�;Ƭ�l�_6p��;�d�KR7���:��sf�'�$�߶��ϴd>s��f�H$��AK\��jOK$���s;�d�!9>(��NԸ��0�u�x��4�xQ'�]�B�*�T:C���jA�d���q�����/T�PdZ�ܝ��H�$��1ڨ�<Q'�����]����NK;{�r�fQ�-�&k��F\�A��n�Q4�O"Qz^�q���_�d�&�ԍ�d���/���zY��\n10a�8�1
+�U���N����g���w�wQT�U*�E���J���9`���~�oA&��@��:M(�U.�|- �H-#
&z��K�s	]5n�Q,����k単�(�h��������[ά��#|�9�B�#E�Kz��H�$K��͓�K��6rOr ��2�"�K��&F��d�Y��J�a�0�r��n�Q4�R�Dd�=2�H����擦��[�{s�����0`��.&���k}������Y�͝��R�֚6Oq.K��>�[$�#*��Piօ�����R�m��m��vg������L��GH�s�yO�{ʴ��4���Kz������A�Qp�$U�
I�J� �S�7cË��X�;�*N�A5UUR��#J�++ ���4��T���v!wI�iDҏ��+����A��f�J5.�FAzS��L��},ﵿ��I�Ā�e^�����>����W��(�(�-������6H:����x�ir^�gE���iDҍ^ՆbY����j�ɯ[���L��}u��de���Lw�͒�sGJ2�c�Q��Z]͙����X�H�D�F�VF�\�h��Ɠy�l�w���N�E�M<��+��Z�h0օ�|�ł�j��G_Z6Ќ���dFv~��L�5CJ%IHى�2������%�;��;�>��R���6Om.K�no^���¥Ba��V��XuT�����{b��n5;w)�[[e )���e���U�E�I��7�26�K&�q�v���6��t҉e�R��ª����:Q��g��K�l�l��!$�&A��֊f�l%���Ju���͝�d���Tl�(�\�w0݈]�AiB�ƃhJ��T�w#�q��Z�u��ﯧѝ���u%�$����y��K6�T/yz��f��i�۔�V/��^�h�_2	):t�hah�i��^��MZ�"d�6�j�}�Ԝ�i��͡l��W���Ժ�~��r�E@�#�g�=�Ϯu�>{ڸФt�*毗�'��v�"��������)�L��XQ1��Mڶ��6���X��&��vEA�+2Tm�ۻB$���1ʢK<���ч�����&^����`���n�w��{Vj��^�fA1�Ɋ�
�k޻��~������H�Oz�M��MZ�"d�6�j��]��"��/J<e�q����b���P�ʳ��x���Y�{�G}כڱ�H��NU�!NuW�<��F�y��E+ؚi&�'3��H=5W�]2�x�s;m��R�Uɐ�SV�W-Ǻ�F��L(�����;���ۮ���.�e�{�	uSRz͡��{�x�n�e6�M	�ט�����(�y
��Aɥ��]��]5Y*TN*�]K���w�B�ʹ�m�۸
�U-�*�:����s�N�p(��b�Z��e^���Oa�-�ޝ�p�U�m�B�Nq�z���� �� 
�V�����;�T�*��P�t *�l��   � ��
����EN���i��@Den���E�mF�6��c��+�{jӇn0�e����C�)�uV͍V�d�1q�K�������sڽ�:�rOv��r);��]qosoZH�� �m�Z�uU��)<���k\x=�L���^{w����
c
���yM�}7o�Rzo.�7"�B�������v��ｯ*a�(��۔r;[׊%�K��uR���D��_gʹ����*t���C-|�]Bu}jd=CިW�h	LLC����9����_d��A��-�j���]�TOu���*�נ8�Y��@ )��d�C���06Lz��@T�H�"���D��r��lC�|��(�b�&��$R0_���(��k�ngw}ޞɁs���S
`V��lfU�+�s����yp�[��%Qn4�o�3�\;o_����uu}jd=C�!_���w&t��/��b���Jcj�6��N(@>�Ǫ�D�/)�D�r/�o�@H�f���k�ն����!�PP�A����f}��~չ��e"=�)�0+^"ۍ�U�v������lq�e�KUU[mAt���-` r�� 6�T�I��j�T�e��V6�Z�|�x�uV���	�d!��j���S#H������_�8u	8("��L�9����c�Z������=��S��F��}��fw�����Q-k��*�N�����8�"j�,�Ӱ�_*B"�e#蔪~����bl����aS�{֢�u�~��Of���Er{;�=��N}������-j��բ�jLځ{ik�:�J��ǽj+�:ߧ�������,�+-��m�V{ufۥ��<Ix�;9�i�ڥ檪�� U;Oꭵ��m��߮3;�����W��X��U�df��:�R��秲e����|�`�~h]uB)��c�|�"]�����B=�)+�2!dH�s����Hwia���qp�%���;�����?��L���!�/������O�J��H��,�����[8ʅ-�]vg&?\{ݿ�?Yʛ*�k�>�q�~d2*�i���O�}r��Й"F��#G&Y�}];?i�T��_x�.q~�q����xϦ3�;�k��6	d	�����&����k�E��]�Շv�d)�U*�2��Ѫ a" �i��w3�S�]3I��S�LO��*s�R��^3�.^�(�����T�5�r��YљW�+��(B��s�%^��|���6Y��L��r�� �VcAI%Q�T���Dg��Ĉ֟��)�S���N���"�]�6Z(�eѪ�dU��w?j9�LyV���q?4������8�%N1��ɟiҚsKq�I&[N����R���yYٙW�<~r]EG�>��W�#�b�w#E��[����݀�S�ܽ5y��%�v�Q�P�`P�T 獣j��ƪ��T7�=R��Ԯ�*�@�@�@�z���Z� ���` �m�ח�LZ5�%����G&��[vmW:�0���[��Ii����X�+u��`��*�� 0@+mEP�U � �T��@5ؿ�ϒ�niV�P)Ñ:���rR�g2Ѫj�����B5�$��R�]U!K/���UL�g�QIfA'�a3|��տOܿɖg��n�*���C*�Ї�yx�����G2�%D��[���gK_ﮧ�G;��4�t�h{i�Ȣ2ym|����H�:�Cu�i�!�<�}�׬�����<�QٙW~[����������T��Z�����]���?1��(������t«O�!le��4�$�1%���ޮ-G{���jN�Z~�q�������?3��'qY0�`�n�%tULo+�4�k�W�w���n�]ն `͋�m����r�ϟD8�W�ۯ����y��}��n�379ޘhhX���B���V}��rU�O�k<�~d
�Z�|�a�-{�3����;W-�	�[b�]r~��r6�?w��IJ�60�����3�/�����_ՉTx*�c�|��[_&�������YU����~��3�d�������5����̼䯽����Q��������_*_���;��Ë�n�R7 	�ɔ���Q��NI8ゲ�H�lE�Ъ .n�nc &H�HArf}?s����~�gN�!���r^˄}�W1�V~����-R��G~'�v�:�����y_&�������YU��{UI�b��Q��W9?}�ft���vfj~��S�n����`"���@Y$Yd,�FH��E��I �0X� H$HI$d���I����$�X
IB(A@�H("�B(I,I �BH(AHH) �"�$R(����!"��I (���2��Qp�������37y���f9�g3�~���j��%a�տO�ג����0�����J�!��^"w�s	����d�b� ڵW=�'�J���5~C=O�@���k٩0���o޷m�6�
��:��R�=�����Å�PI�����V�l�*�C��%pm�5���9�\���ՙ�S���?-�C�Q��d������hQ$܅lJ�@�'�fk��`������A��ѱ*����ʢ!��XE9m6��$�m�W{�@��k�^�����?6�����<��Ma��$�&�m �&g����^O۟��q3���T��,��?-�Cڨ��T�4��J*]~���w��O��w7�?�w?N��@��wL*���(�Plm'F�jTd��nǎ�:9;��P�V�V@� �5н�nօ��߻��WH���m a�I��O�Xk�������{��%���kQ��_��� a�y����U?adG-J�s5>���"1-Y"Z�Qr��߾�[�6����b��ji�>/���N��*�ck�-���O�L�ufv~��:@s.�J�h�G������3-8dqPKKk����Ϲή�3��:DY�y�����)P��"Vە�^j�v����d;;`�{]^���	N�P-eٻO����e�g����.�:���UErq��u� �*�T�v�Bwj#K��3��ا?n� �[{/[+'4p�m���l�=i�R�1BX@�H�-�[ U �f�{d�����UT .�� *� pT � � UU�T ��fٰ�Sg�QT�z�ۻ�v�"�㹸��j�bݞ�娞W���)�V�P����][r�1�
P��~��雟���9���I*�~��6���ȫ>���>?xz��P���1�h�,����'k��"�T���#�o���Y֪S�g�S��B��X�܎�3s�8ѱQ4E���)��F���A�?y{Zs�990�v8[T���0Jb��D/Kr��4�?9.��g�e֛Ϟ��|��� �@�,s RZ^�lױ˪sם��6�If���vZ��Q��Uݳ�gzO��7���(ڪB�V��
��GS��Uڿ/��]}˳�����s�s���]�j�N�b��ai~��d�wJ1�;;(I�亅�={R��~���r�"�S��A�Vx�Y{�R���>���ZW����M��*�A�������R�ۭ�
���<_�c��m��i�Q�� ����[�T+6nV��29��x��s����Nq�"M��f�%*��i$p�m�+��W)�؍��e�j�*Y[j��v��;��N�j���o=�,=��Ӵ^�[�-G�������wL�m��N�����}R����D�XW6n^���L򟦺L"֖� F#x����p��ϲ�������.Eq��BV�[��)������w�m�9y��ɽa���9������;�g�>� ]�k$j�$��;.���֮Z�e'�wf�ymΊ�X���.ma\�٠��ۦ��ک��@^��Gj�"Ɲݝd��4���w�$-��C%� �����w�OzԪRk�^��s\�*�\���{ V��F�����M{G}^��z�R���+o���Kt�Tm&�h�������Qr����W$]����o&�6��d�z��
�M7�a�9�X�N��Sn�ړ�)�l��^�w�ۈ6����n-�۫����N�n�*s��J�Sy�Wxs}������ �sBҨ�u=UU] �˘��i:&�`�T������L�
8��
P��k{�Y�jt�w=�\��v�Wd]��.�o&�5)m�e&�L�x�m��d��,��c�:�=mב5'�]Sgh��#�4&V6�Ɩ6��8q^+�-�8����v��;�o�oou���\��-���\����y5�@��2<��_��w������B�*���u�k�/|l�Nn��,��c�:�=mב5%̹���)kOQ��e�����p��vNu���@R8�G��r��+)T
���+5��QYtC��0�ؼ��n� +%U*U�ó�\�:� [�������%~S�l���u6���c`s�7mNCC�S�E@�%�^r�2��Wq� +'t��p`w+(�*���[��  �U w   w �UJ��]x�b�=�PUzAۖ��ڶ�*���R�ۅr�y��??|z��B�¶X	V�d�P������A�qD���_m�\��ޒ�g�ܜ\v�v3n��͝7G�8�l���)��\���&����u;�������nM����QN���w�vo��̑9�/,��5�T������Q���(�k{���u�I��=��j+�ȶ���o'|��q�Y��'��S�ĩ��y+QM�m]����l��R݁mA���ۤ*�4ɺAuD�R��8�x&q�t�pvd��D�U \[������u�]�N��]ۭY;�i<�v��)x�ל��x���!M�ր�)
���7�{�[�k�j^�z�ޗQ���M���2�0Qia$�M�����N{��Z�-�}��\�ܞ`s����:#`���t#��rT˧6�z�����;+������šb�m��8w9����^d��.������5ӛQ$��|��Jl��Wl���Lv/6�v��sE� `���52��^�'�jV�cac��w=��y;���s�ej-�'}��\׹��Ŋ�5@RH�$����ܕ2�ͼ���޾�g�n�KsԵ�Ueh<N=�o��ù�'_�m��$���M��Wf���X��1���=f��^e~.c>��&^z'ｭ���u��	B�%�4F��Gk��2���`RZ���%��6���Վ}����0�3�_51T+;�N���f��z���S�J�۷m�xlz����RN�:_��Uw�:���Sܱ�&��c�8��J��dTbS0�Q �m�����x����axN'Ӟ��]��e��}��z�e�	���ʭ�u�[�eu{<:R�;�)-kkF���~�)�F�+Kl�/����/v��^t��.���������K�r��
�
UFd���n��[6�h�����.�����LDc�4a@y{H����;n��ホ"s��M�xU ?ezάT�1�aō�s����&����||���^�W����M�%�T���Xc}g-�9ӽ�^���^t��/'xM��(L� �\��}����&�\�w�-�ٸt\��\�g6�"�	�y���&������u��4���i�Ni���>6}����EjGD,�$Kl��r3�g0~��M��6���C�b�_�p����/��GG����w��~}��a�<<��.ˤ����gOlu�������{Un�y���̇Iŭ�̚:���ȓ�������r�j1�3�[/g�N׎�׍�K��=<O\͍����pVmBn��c���Y�+�g �&��[g��sN�QG�v�ѹFp�H��5���N6�Ks.���ӭ��@�'F�[�՛��v�\�����T%X� wn[*��� ��*+(UY��J�Ux   
� �ڋ*���zuEPr��l���T�UTI$Uo]�.� f�T �1J����  �^@Um��{�� � ����@�,�G� P*�*�6�T ��ʀ *U T  *�� *� U ۽�v1����TvL���<6]V���6��
��{j�����]�61Yܘ��0*�L���ؓ�`��zyZ����iT c  ��UUt�i �S��$M��:L�y�S7��ӷn�&�
����UZ��6������hB�k����Vu��W�����s��Tᝲ��kul۵h��/	/H\��]�s�a�^�t!����i���eb���8�YT�u�j�6�w�w��=�����^m�ې5�`.� < k~�7
��  R�@  *�(�
�  
���ٷ�� Wtu-ҽS2@ s          j�[s   <    �    ��U P ͻ��ƶ�
�     Ve Um��  ��@     p    6)T T      �          � �  *� ���� 6͊ 
�   ۛP  ��[h����Wn��绨�     UVL� 7� c��  /o2�@  *���.vu�j�r��p��m�C�+s�4a��t�R��+�� z�c�U*��T�Z"��B@�H��T�V�ۻ[w�@ UR��4��5�z�b�R�r�ʛ�J�f��Q:��ͷc����fݮ!�nW����{��4b� *�l��;��TةP eP � �P ` x��UJT�q\� ��Q��VQHoLiV�� j����m4&�J�. ��� ��Y��ٶ�̐��"S5K���'Og����>8d����Z� v��SPl����iX#%-A,j��g�m��_=��~��{
h�%�O:f��f��S�o��)�keeR���;u��DC� <l�զhZ�����0�%<�d��[H'��Ǎ���@3�p��ϛ�����o4Bʈr�_���i�I�4S����8�yP�y�ߴ����U{�<0�w]\*�{pƫO�p�#�����Cmp��d��*��q�s�%*�j�jU��m��ukFծٕ�I��=��=�X�ey�V����C�@x�ݫL��|�Im&O*�I.���6Z��ɦ*��W�ýݯS>�Q�}ｮ���4�mT+T�����{Oc���4�LW��I��꿸�����=��+ċ/e6�'5p��ǁ������V!����zh�E����>�C!���4����Ç~���b�~���k�7��4Y?x�,>�������)<�S��w��<��ʯ&8ւ��I�tU M�����juV! 6:�xp�g��U��;t�-�H8�<�]��~�%Ƙ8�XZI��(ӧ`��4sU��#�eث�3��! (QѾ,��Io؞ffV6�a[Ȁ������C��n�O?o>�N�H
<:J�� �@�v���6��q7�{����h��ewp�����g���Q�t���4�t�	���U`3����n�k�ݢ5^?t��7C߇3ƭWG�>@[���$�g�-AYQ���U��a�^���Ե�fQ@�U*���ӧ�۽���(둟�s<?_٩ϳ���2n������ey���Ҥ�+$^ff$�y�t����%����-o���g�����Թ��M��@�2�m�O=�OJ���@�l���5�f5@a�<d�W���#�UR-SǙ��-'�GN��
;���AᏫ�gtja�^C��X��	��G�)Ī�PS_J_�����n}s���g�In��º��]ޑ�8VCJe�b�Qp
��Y۪8!����z߻���PW�N@T��C�9�f׈⁖����3��ͤp����+�0�#�����_m��F>��M�C�AF�X�߇���f����u�v��2�@�W����x�Z��s�J�n�eR�M]���
!��ө^�����#���%O~"�uh�eu�s	T Sm����?Xn�_e�i��ud�+�0�#��v��oO1'��F�*���N{��>��<���w/�}���x>-B�(Sd��d�i�
B3��s�\�ՙL<��9ðq=����UMF��P۹��g@��U9��z�qW����R�  �Wz�\��?{��U^�-�x �d��g�w��f�9Q�ۀN���X6�v�s)�v� ����͝��@ 6ͫۓ�6�ݺ�m�@ ��@@m�;�l�l pUUR���e^�m��VWj���=1pl��I` VU"pR�n��<���j�r��s Unj�R5�0�8���~w����=%~��.�s��T����i!�Rҍ��y�9��x��u�n��wE�y���ϻ�d���F[UXQv�Ї�l	�0������0�.��ey
"ݗ�B��m�D�
U�~�4D��0����޶~�(�ޏ��Np7��wg�MRIp�N�T��=�-{d�K���x��{�Nxۋ0���l�Ik
�Uk�+jۭ��s�;#d;����7;��5�,�. !���ޝ�C��w)o'�����Y�w$ۉ&�F"�3	�q�1QFv�Z*��vJs����d={��w/�
��`������;r�^��s,�2r�8��w��_2
�A.F����^j���7�O{O��P6��x�g��C�6[�.��F�)RT�SI�Z��Αd@�u���<E?i��r�L0�Ǘ;��ϋ��>�tm�^B�cG�S:��[�ܑ#�a�u��m�
���m+$q���+h���z3;?z��'����bW�����-��8G���xa)�*�#�&�	��m��{��>��ca0���+�~������������W�����u�h�`��ckb4M��J����g�v�aS0gH��3�%�"a�7�c��-�������2����	��t�y��!�����K>#�[zp,Kh`E�m��=��ҥ�W�#��a�sa�"���"�|t�l�ca�Ҳwޱ2Y,����m�$��UҪ�� ]��k:йm=�g@UJ��f��73L*uTZ�C�C�?~��C0�������Eέ��F���ӧ��l��U� df�3S����h�ɩ���ֶ�|1��t�~c�D#=7f��e��^6�Oz!g���V���P�W�"<Y�K�H�2�Ǧg�953��-�#�.�j1]?B:mӸ�M#ǧ֭�C0��A�cڝΫ��]��$�K	x�c
&�o@O�ߴ��w3};�c�V�S��;41�7���f����� Mm[[%��=k�2�iZ���[ m�m���'����m�{ӿu������;��wr�W�om�Ǯ�G�l�D-$�8q�k���w!��j,�����9�z��3�>{<�\�H�ق7�i���4��{�_e����+2T�^K)�!�8��g=}׻��i�;�{9K�e.�|��Fs�N�T�SXV6��3v/U���o��\2v�o��y�-ɱ�qU�}���	�KpYaWIj�[���;FĽ�4�t$0�U*�5J�T�eRS`.�Խd'�����&��6����  W�[T��8]g�ߞ�[w.�J)R9a�\l��(�gKa��g9-�#�s�) r# lһ4�UU)>����<VQ�UU b�m���  +��*�AR� n+d���`�o#�ۭ^�����h�-+HUz���#��ڞ��ݦ��M�T*���E��d��`�N�;Gk���ҋ09=�������}�s|�� ��}TYR��e�ى��GN�k�D!�xf�ǣŔG���p�x����:N��A6�ӧxC#M��S��0s�U�8��d{M�ͅ�Q��i=/�R�#	��<�K�f>��<t�[��L#J����t��W���G=�W���,�M�Y��x|zDs���Q��V�#�����"�8{�{n��73�{�rգj
�`2��U��\	���&��ݖ�n�N�R�+���Ҁ[2d��V�s�����m#���jU��L�U����{M��٩����]�=��H��TU�V��=�r��a�eG��ψdQ.�����q��隙���������ma�?C�Dw/7��ǤJ���Ȅ3�ܭ6~���b��s��?�Pom�X�����Q�kɖ�ׅ�l>T�t��--�D�E$�l���2v�	��s��h�Ͳ���|讋z�Mg��dd�lh���z��wg��e�,��T j��T^gE�CD� ��?7;������+H�ҋ��:":|D���p�!y���jg�R�\셅�.Z�����C0�ͷ�G�(��)p�x�W.^��f����aG\��U@�Rm#�boI���=��f�tݨ����@�>�~~o<�:�z����㡦�"�͝�Ӥ(��i i��eQ�*�dx�	ZG���f�e��������_z�d�HZѐ�D�+ǉ�z��v��s��G<m��k����mn��C�F@�g��ר��C��3�-UU[�ɶ�ػ���� �VYT�9�O���q���2{��5���v;�Yq.�m4,m�HHa�:+�X���w���}ɯ��^ۮ�r�^p-2�QI�C#�W�o�x=U�r;u���)�r{�0�[fK쌪�$u�s�w�6+�n�|��!��hx�}��C�T�X�mV�{�w��f�ǹ���u�����}���I�rj�`��V�waj���F�a�m�Tgv	�6&BeZ��j��� ��;e�?^���U����^[�q3ꭜ�n���;Ǵ ��(�={���μ�nW�3]9��n��.R,MS8�l�/w���h�?J���i�oB��Ǧ��':�X���8�׳�����,�.C'��f�ǂUl�J�V�"�(����z��'y��q�	T�|������+�� �3d���X;�c����Ӯ��T,��5UU@l�R�q�VٰźG�����˸��PT VP+m���o4yy�ꪥe�m �Gg�4Y��x�naێ�����Q��g�¬ݐ�����ZU�����T��m�� ��f* �  ڨ�PUT��x�M�9luP[6�j� 
z	K'[]���-2�*�xӳ����og���� N�R���A��xh���F�x^<�Nݡ���;�vm�g��-���zpՙ�YL��m��0n�Ӈ�������]�>"9���DB(�}�p�l��ǝ%@3M��kLcZ)��6�=,�8G}jp�x�e���x�y�*�G(�Ol(Z�����`��=ɩ�׽�6D#�i��M#ǧ��uh�3�-�G95,�f��|RVQ[J"T��o�E�G`�!��h������o7�O�H����Q�X�u*��Q�hT�ʢ�U�-^�����ef��h)���iPkb���iRI��<#�L�%[\�v��s��G�Oz림s^Γ��ڑ�ع ���Ǒ��L�M~�;u�d�*��;j|>��w�HSd�\�aAL���8��Y�(��*G��I=#�J#�tvY3�S��=�d�I��AU�Pn�DB�˰�:\bU���=3m����#�w֧�G����I�ƚA6�ӧxC#M�f���,|{*���{L�ͅ闋K�x�7�ɷ���R�P r�*�[�Fw1�L��)��Y 
�U��%��Զ�c��<�m��0鲣�ǎ�C"l�0�*��VC#��I=#�J>}d$ق��)Q�N�u�gf�'�=����DB(�}�p�l�jr��Q��x��(�3��ER�A&�%5�ٜ���;�p��x�r<Q�g��"�|w�o��ͥH��'���R�G�m�O��}x����R�Jc�J#H��.�mC�4���zns���m�m���ۮ���;�a��M�{k��M�9f�l���y`�I��h0S�U��M�捁Z�c[8�5�]#-cu;�p�� ��[V��n6��")�ss޾}��N�u�sMx)r��J7�zH���vS�4�HcI6�b���E#���}5��Ҽb�z)i��M�Lx�DiWC��z��﵀_��[��[P#��na�=0�U�0����dC�f!���m(�C0d�ѭ�+�S�1%�$�m��8kE!�Ev��:Q"����j����p��>Z�2�pҊ﬛��
�
�Au&z3��L�6�E#��t�Z<+��ƊF�F�{
��edwQ%O�[��6ꩵ��*�[9GN^�99q���$�U),�� �!�D7]��Wn�ߟ�����P�¬�G�|-��0�f]����_<�Q�.�0\y���%&��ѭ�>�V�C4��ך:t�8E�W"�3*�ʹ|=�Ӵߖfi7�nu�tw*U�R1
�.i�3�y�+�P��*�,g	��m�S%a^g����5��>���:�WM����������;�忒�lX��Vұ
F�2v�և��F��4R4�+�^h�Ҽ�H����j���xD,:�9�8������8wTͭ��rYѭ����N�Ē�M!2MU��nTs�h�����*�ٶ �   *���l�9�i�!�ءU[���V;	�"&�ګ���\�I��n�R�����A0W*�R�ͪ
��ø�wwUJ� lJ����   � �*U�R�ïM�6�m���*�ĸ{q쵻.Ҫ�]u������oF=pPZ� +m��z�wwgzG6�$����G���
�eCM+U��I���X�SB�Ӷ,V���ޝ��X��6ł����A��¨i��#��*"]��P�<ze�r���S{�Ys�I����q����q�s�iM
F�2v�և���Vh�i�Wn���y��i�ڍ�T�C^��\�=yנ�<t�e�j4����E,��=�K�K"��vmOx�E����Z5��
���F#`=���gH�8;��!�����<xh��K�E���ӫl���Itn��9���6nUݼɋmp*��f�=��{���:�*	����:a��"#1N����0d�њ���F�����"�A�Z���,��ō=��"��:D�S��ǰ�G����eC��7X�zH����}�^5�6�����Dף?e��+C��_[�OԏBn��N��ngpמ��nj<֯j 
0��#�d��i�*;���#uzL�idS�
mѭ�*Ĕ��
m�Ǚ�E0�E?R.[�4x��"֮:E�S�U�m!���(��P�]�׏��oZ��5R���edb�� <���cdX�
�� �m,�m�{����̌��XAw<��;�=�a�W���Z����U�ܓ�IICX�I6�FcW���A���2��iUCˇ��"�#�C����SB��l��,�-��[����u�l�zf�Ef����y�aw"�!�]����rn8{=I�҃&I\,�V�^ڇM+��פ�Y�{M�6�Фt�&.!�»�kE#���k�lj�kT&LIu����73�{Q��8u�C؃"�Gw1ʇ*����}����}���`�[E b,&���>ndCz�nݷ(n]�fJ��kkl�^����p����g~�W��G/M�5]�Qt�Cw:mB>��KeX(�[��gf滑�^ʇM+���4R�;�'�ͥ5H�kݚ�'�s��{@Y�x��,m���G=>�ޔ�:T\"��]4ڇ�j{"�Gw1ʇ*�y��֎�$�Ji����E<0��z��-�5H��p�͘=sw��5|ϸ�y�n"�!:tJ�⓴����EDC��͕W��h��w�N{�[����ߓ�^i�s&�f��kuqj��UVݣV�n�hzݳ�'�m{�[h\�* �uD�ƄƸ�Q#�uٽ\��p�����x}	�)�t��E�t�j:ġ�L�zfޜ�ĚKI��!<͕W��.����{�=o3ٴ��`���!�,R�"�zW���9HR��YJ�;5/o�9�hB{�:Uw�7�p�ztd�eC���wE�,gf����{-�!+�*��
.�+i;a��n�O�|��G<>�ޔ�:T\"�t:i�#0���ŋ7M���^EDC��=m��0�\�vb�S釽C��=�Jj��	���B<�� ��*Ӷ�Zְ�[��u�u��A�혪l�v�.�ӡ��;6�ز9��6Vy8<�JjŐ�Y+�����&�ø2����t��l��6���<��ʧ��yܐ�=(=d�6␘��g$�p�d�n���>ەm��"�͒�m���jwP��D �pA����/��G8kƙN.
�ņ��9�^<׹�PUm�l��I��^�TP��m�U6¥@�mT�  +mm�������-�=�RnĪ���uAW��=T���Y�{�� �  *��* ��  �ݲ�\�-B�*�v�T*��U U ]���P �@  *�  U x Y@ �UU*�  U �
�� ��w����nwolxGvv�U!�)��M�p���ڮ���ݺ� iX)���ge��UU�Z�SR�K���vK\ש^5ʀ�
�
���sommy��V�d�(M���㴵2�
�t�9�� #>��Sh�`� 蠯#VP�UJl�8xmz�Z�����Q/Z�l�"�d+�9������kN��M
{m˄�sPML�R��<�f����t�m��[ m�����KpoT;�Z� ^�S���wfz��E�
ݺ�� y+whP T]�  {p�����  V�V�Fص�C���k��   � �      �ڨ�   �        
ʪ�U  l���j��4U �� P @P[   EP      ��    U          T         d �  �  � sUUM��� @ k�� �
��lU�1����     @�]@m�Z ;�: �@u�T *�  �Y��a�ie�gP�'X�]�V|m�۠�����s�'tK��/L�HR���+XǛn����uf�J�����*��
�[��;�+k��$EҨ����lc��9=cn���ZfT�n΍�5
�Zch�l���m��UG����6�� eUP��SP*�*��   � �UJ��?l��ثj�U��(̛�����&����Ez�3g��2]�ۙ]� m�	@e]�������X�^�F>?����؆ʋ�I֝qg�[��w�Y�k�B�!��bs��~L�SØ�),�LccE,ýB[״��;a��n�O�|��G<>����f�����ג��#� �"f�8a]��2!�ws#L*/Z3;��:a��s����}:u��(��i�x�f�ȇL��)�)���W�b*/�����F�|���+"=՟,�� Dm@RBU5隝�W��JƊY��M6�6��#�d:_�#ǅ{L^���*�wT�)�O��I��@UQ��7���\Z��y���Y
V��]�U�u=��;3�U�a>w�����1����=��M����aQxۇ�Z)���βsx0&q�o1$�[
��D�p�!�4�Jt�a�U�h��H�7qæ⟨�����!+�[��gg�]���^���n�X�K0��m:�#�`q<������K\'堶����\uٜ0���V��E�Q��0�]U?G;h�̳}�ۋ�7���6�[��o��f�mA�5�=�;�>=|��̋�9�z\�ʦRB�E$K�h�*�@7�	��R��3tU[p�J�T 5����Rܩn-��T�f�g�_]W��"��m?C�StJƊY��A��i�P���s�/��<!5������a0��"7�~fE�Q��0�\��k3��{��1m��B���O��zй��N�t�[��_#M������qH��������2^6�i:w�2/�-�h��.��E�C�n{�O��T����a��H]��,�F�ږ�zi����q�y	����(��F�z}W�D<*-"�t8i�5�{D=r�Kc%T-�h�8%V�]\�<��7#P 6�T�m�UZU��r����߽�C�'=�yyuK�}�M�A�5����*�4��t�,*\ێ)o��<◯r)mVwGӷ���#O�ے�*[ �e�B��I.�z�-X�����^�Ե�>�
^�Bd���W���:�5����]}=���=���ӽ󑓙���X�IU���,B����O�}����նW��NP��$!�J�
 `5U�K�Nz89�n��Զ@ ���\�{�%hL
6~ 7�_G���ӛ��-B��i����;�*��y�a.b���S[m�2KUJ�8T_pO�C�H��z�^E�:{�[u�Yҵi�ޱƌ6r�݅�[2+U���%���g7�#�O��
C��-W��T_xLuޜ:F�m��4m'M�l�����:\%�f�8|V����R�="mW�i����N��ٜ�������#DU [a��|t�<��*/��2|F��������m�D0¢s9��A�N�p�Dm�M7C�u����nG1��Żr���&���uUH�*�g����k,
��HM-�ew]�Q�*��R�����  �u�vPh���q�z�-� c�1�{M\ �����Ni�3��d�	�(���t�;��;���M�R� x�@��U@`��;� �TU@�V��� 6�� ]u�[�qJ�h��Ň�����@x`v�-�^��t�`�Pwzm^��ۯ{p�J���U�ë�����C�_�7
����ݡ��
����ݍ؆ʋ��v�ۖ���Udu�N�� w�ƹ��p�x���W��E,ýBp��������� ��=�R�6�	�����@o�{��t��J����e2!��]�����^SJ�N�UT�!<ͱ}|���襘{�,��5}GF�7k�>��_C��%����Z4i���o�t|��'{[�횕}��ce_C�+�/^�Y�z����k��kE�;@�q�Bk�m��;v;[�����T�
�[h��ڥ������u���{���޿�;Ξ�h��a���3"���!�E�fvY�j���\�=vr{ٽ�/��Bq���q����^/��ܕ��}f^�#H�RIU6�TPe_�a��Ǜ�2/����L�䢼͕}��u�_ݜ�;��ʨI1�cm�W���z�᷻N�����}�=�a��a���+~�"��]�i�q�q��Đx6�ɚ��U�>5�kl_C�P��X�Fb��p�_Q�ˊX�y���U]�ej�v��׮��{W��� 6�J�T�B����(hM6&1fú���0R����)����2/��^��"�)x�e_C�5�\�L�e6�of%��67�}���z)f��^�-��\�M����ǿi�M�\�� �fj-�u�S������E�f�7��aF��ƶ��=��/��z3������R ���H.�x���rV��4��4!U�0�bV!Ң�(��tȇJ�tbXIU���i<)b�U�>.�ʇL+��ע�aޡ9U��S_p�)ΛP����x��k�-�e@U,�T9�g�=����5Շ)�sP m���,�[��& (D�5��vn}�^���K��FCL�p更o*���m�pµ]�E��?�d�MZT�]�6a�!�}���?/��<��!�g�hB��"��W9y}Ǧ�e�Gj���M2!Әmj�\-^-��Wt��Y�z��W�iM}�m��%f�m�,�<���A�X{�0��ũJ�
��2�����.Ѽ��|\ڹ�(�T�)�v��e��߰��g�;>�:_i�U���ܕ��8wU}8{��$q�ūQJ�T�Z������g�y�W�=���ؔ6 6�T�m{m�\v�0,�����MK������N���o*�,d�eC��wE��K;5��w^�gɆX[D�u�U����zW�7�=�L:{攥h�ʋ�����a���i�S����ec[ʾ�ƺ9Ǜb0�!9B�tR�=�7�5\+�wrV��4�^��$�'��Ǎ3�a��i��X���c�a��.�7��2ž�t¹N���8�e��%�k��;5������S@p�J�W��=�4���J�
�p��h�!�'�@���헍n���#���$��I=�x�CT����*����f�]N�N�+��R���k��T U*��w���W�ڧ�k�bRU(�fVݸ�\i�.ob:�*c��ejL;��c'i�fL��v�8��/������u<l��J� �P �`� ���` ;��U�-��lmni 
��� zz���f���"�ѻϏ=���qmuc��� X��٪���eT�6ö�`�]�[�?���a�~ʼ�Y����}�a�	��tz罽����Y�8�ۦ�E��9����8)V[��׆3'd{]�x�ݚ�ݹ�G�eK2���7��v6'5��o9oUWM�x¹ܟ9ٚ������т(W��b���c��L�p�h�D4��f�W�j4�(yFw�����e>�S���@`*�ڷ^�w=?w��٫CN�C����d��i���_kў����k'��GKU%`R�2�V���=b�.&�d
�ݶmڥ-10�[� D���o�5?j9����P�q]�z�����!�m��SB���.�s�ɣ�(I$=!Q������bFƜ+P�9�T<{���ͣy��pr��P�y[ޮ�����K-��[���N�{�=v��+�R4����B��)�E4�Ѷ���K۟L=����0r�\���g��
���CH��ak�m�tҺ��zH��{�#<�6��R8l���ϛE��T�$�7Ʊ|V�|á�i�:V�xTC�\t8i��6��CH��ތ�_�V�e�D ��)JSV�@r���b�� S`�U���[T�HW �5�\������Ͼ�2�0��Yy崭B��N����)�zg�����>W�a�-E-��viQ�2�=��P�W�=�2!��ʽͤi�j�E��E,ä]r��c�ZtKuU@��\7HB<`ex������:=M�� _�^��m�i���~����׳�ڀ6����	(�ۚ���v�����<�Bou�N�zG���/�B4���t��^ʂ�^p��m��C
�Hᇦ	�ǿi��2m{�~��9P�!�܁^���<��oQ-,ƃ�f�Y"��Z��W`��S�6��*��٪���eT v�J�cu�� ��oI��4�͇Z��0��~��h8á�YӇ��7���6WeQM� �M��1|p��g{��BȇO_e;��9�6��8��ou��B�a��RJ��d��"�Y����3)�E0��;no�ȇ�6��L?[x�}sS;7:{T���Q�d��^?C�)v��$S�"����0�~ӛ�c��gN޶LI�.�l�m�R-c;���.:4����F�!�C�v�����y���������w��&�ݣ'U�j��{d#\�(ݬdwb�G�,��U@
ogu{����V�X(���w;3S���f��q0R��SLo��D:FI�60��� �e�<Hʪ��u�\����v*�m#��]�I��6�\+�p��C���s���Se$�cH���!���Z�:!�Q"��L"ʣ���!dC������a^]si�B�D�ꕫ�ݑ�>#g_�±F�^�����S�a�m���ϻ�z����h5DU��{��{�Nl8�U�_���Mٱ�T*N�(V/��-9�帮�۝�x8G��;�&ⷌ�s��mj��.籱M��xVMݶ�b��x8�6�U���mV�T��l 
�#!� �P�6S`�u��J�AJ����4<S�T�gO�\��ѹWs;3%V�8���j�
�J��
kh�l��eUPT�T 
�@;�� ��� �P m�U����R�� .�[N�lg�YJ��:���l`�c7l#�n�Ψ m�T�JU���c2M�T��?���l?W�Ѹv�Ed~u¡��N��+"73��٢)�-6�M1���4º��<�z)ᇤz�Ӱ�(F�^�����S�SO��`��	[h��Yٹ{~�Ӻ�a���=�H��FAz���
�.�|��S�S8w߯Ũ�2��@\)�FƋ���
�0�H����t臅E�\t8i�i�Z�I��p ��l�T/"�!����N��0�!��=���=n�saMB4���t�t�-9���o��*�H -T�n�]��.��(�ln�;3�;��6�y��^R���<M�[Hᇦ��D,��D�x�am�Oj�!�ѐ^��pµg�<
F��!HIp\�z3�S;��V�#p���a[1&it����QYZ<���$�J��*�t/�E�p�w�Y����|E�W�ۃ�sE,��=]έ�5��夒�4CG1"V7���X�8E0��o3D,��Dɵ�:a6ާ�i�h]\���0P&.צnv]^�Y�Х�t�O*p�P�6�r�G�>Ȓ�&jrn_��{�[B��
��Q^���^��3��z'9y���d�Y@�i^G{^X��0*ӹ:���ߘ�4���0�/!�7�i�ݣ�y��0�-7�v8ه�WP�Z?e�-�m��cͥ5�����!�4�Jt�a�vm!eE�&M�a���gp��h0�X�x�[ʴ�xtd�i0�R�7���a�&�S�b�p��i�����I����QD2&��N͟R���
�H��p�ҜR��-#����}��پvk�퍑Z5V«}S7�V8kk�&���
%&�Pk���s��؀���m7Usj�IXEݧ��;n��� `�)Q��mV�Z�V�_�<����z�M�^����wnt��w���N���-���*tۡFV���l�?^ikp�8TVG:��L#Jg֍�Z~��9^$�X�M��!���4º��4������2��R���P�l��C��+�+n���,O�q���
��mt���WSڴ�����G+T�OXߙ�dJ���F@U�"�){?{�C��x�]X�it�<e�\�M�gg���R5 YM�mQy�R�>f�øq���z����ۺ�:�겓`�TkD�޺�������i�LԅulF�h�L=#����SP�>�ɩ����}mK-���+.��7!�o�YQt�6�L#�����i���+�0­=7ͷ̒O��KY��8�E,äM6�6�#���x�4î���,���iO�QY
N��Ɓd��3	��m<0�)�.r9��˧8Y�y�s���>#\��|U(F���W33�i�GfӤC�kF����'/�xT]#$��!=�n����M��7��R�-p�2Z�z�8�W��9;�]��s�޷r�- ��UQ�Z��l9�@��Y^j�p�M�2��EP�� -��.瞶��nN^��U��d���a�p����%9�u���g Q���f��S�5m��$��R�U*��0 ��m�ܪ�R�
��T   �P `?���*� ���mm �2�{���]�.*6V4��Tl����T޽۹X�fE�P;$�07P�n^�
�=�o��4���G�h����rW���2�X�<t�h��"ΐ��i��T�.�rn^]L�����':�5Yt���p���x$�A�0�X(��7]�������q���B�)�)�Gn�,�.���8D#����N�I��)���#ǇFQ{��SR�=cE:C#��saMB:g��ϧ'�g�W�ŀ��,���,�5p]�ƚ+U�Π�F�E=[�#N�}�|E�W��x�%UZU���=���g����w{����
�Yfƌ����h
��>6!�0�'y�j���cG��Ў���g#//�<��ͨڟ����8������^��#ô�{��SR����!��%caMB:g%<�H��
��"��#Nm�u�Y�=S�8V�#�AP�"�c��VF�7��1��5 8�^�N˻��n靈�Pp�-�m)�F�C}�2<Y�,R�"����L�Z��*�\�r2��{�M�S�H��є^�#�Ժ/X�K����e��ˍIqcl��F�+T���yMM�mf�q=�u�Vڻ� ��꭛wI��%�[FȍL�eof};��<G��mu�Y�=S��O�Մs�ٜ�M��e�ܷ ��]O�N>����z$Z)�8D��:^!��{����̟z�]�3+b�H�.�8|z]�F�A��y�S��;o�4�pw��A�+{�h�*���A��lh��t�n�`��6s��:�
Տ�i�ᰵ:tBL�78�x��������4���Dȇ���̈́i�w��E<0�n��-x�}_߹r���iCSH\��j��s�۱���E���Ъ ���VǍ��4�H�w��X��O��^=�H��ψ��{W�K��h�-�1��&�3S#y�g�ƊY�H��
j���x���كɚ�����F!�T��̴c:!�Qi
�C��F���o"�!�zx��4º��e��HN���2���6����A}�"3|�R������腕H�Na3�
��l �ic�i�gyW'4(/W\5�Be��JcKݭ������e���UQ��nV��ݪRY^�rL� ��U�S�e]��eP@Clf�J��@����B�Ŷv��O^�z����z�o�ׯ�,,.l����z��N�zE�{�
���M�p����ͤ3L�x�R�=!�N�%YB/d�9�af��z]:D:g�W�ia�+�h��t�n�p��l��%D��f�vns����Q�g��~R�r�{i����H�URZT�mUapS�7��۾{�ｳ^�I��z�E��n 0�� �[Q�z�kj�"V�<l9���o��J8�ynLnt�U�ZX�wI�]�[�˳���s�S��:�lO=�՝���8�ɺl��wAli[4s�Sɭ��&i5�F�6:�=���e�E�ٻE2vI�t����+�ZR��Ԉ�ՆZ��˗R�;^Sj��]����g���c���1�Sh4k�<��F-�T�����R��U�  @_|>P�VP �d���*�U�֠SbV�lPqT,��j�]�,��G	l��^���i@��B]�݀< +*�  v�̂����̅ek;@U��lmb�v�v�< T � ��*l� `  ` *��AT     ��e .gkv�V��;&��AaU�Y%��9s�OP  �)�\b�]�šjˬ��x��=
�ԫbT+����l�z�%�]*K֨Ê]� �T ��m�Vn��� �=;����xV�l�f�L�Raf����#�fs�@P��d⦐ؕ�8�uD���u��V�lq�R�J�㤁wN�5I�,�%T%K�M�1�$�Wss��x���C�|�?��*�	�ܨ9K���Ý�K�KT��f��w���a��,�YdV��z�a7`' �@ +ul�T�P�  wM�*  �
�Bm���C�����4gi�  @ U      ����dq   � T �          �7Z��ʬ�     ���SlP  ��     {`    *�   U    ���       *�� �  � �   
�ͪ ��  5� �r�R��A���ic�R�r�   � ����  �vڠ  ���T7�kհ��ۥ�ݹ��4���nf�7b�Yх3�h�N<VQ[���uS<��ol�k�&�uF�J�� �]��f�`��}��b&�6 
�wv�zn�3�����xGN�ٶb���ׅOt�\Wu�v�fֺ�6)l�gf��w���R�@ cU U�ld `��Cu����5� U+�� m{>	�٩V� v�uD�;`��E`�λ;hةvP  V^��]���w8�6额S�+���H�F�M���͸�FgOw�%iYW$���d?9ƍx�|y�0֟���4���ds�E��S�tQe�i�I�,cag�����4��홊�1N�zE���:a}W�a�鹶�^"RÉ��i�[H�L�x�B�=#�Na=�u:Y��DoV�4åN˛ ��Z
๬�gf�w��a�å��!��eq?ώ��o~���c3���z�VAd����	��p��rn�ӽW�����YAU��	F�)�q�����M���z˚0�h�y��0�81�lC�Ǥz;״�C5Ѩ$�a2M�-�x��xG����v��pɶ�p�#����f����,�L���!���1��p��E�),�[��#��u��<G��9��as���M�Zcx�XΊ@�-`��t��ߑGw�w�Y���]��6r�L�x9\��
aVk3���:���L�ѝc�daݾ�b,�=�PG���2�|v��K��S�UU�HN�-��t��@�6Z�����eeh�l.`,p�i<��i=��=�U�������d�#My���x�u�1#x�~E�	\T��90�N�z��u��E���;s��[�7�,��U�,c$�m[��������<FR�{ZD���C#��
� Y�c�mF�������÷��3�0-��!����d�#My���x�;����Eq���7���������2�<��X����AA�y}���ȏ�~���mקi�X%`gP��m2��iⱻr-�gj���J�R�mU�tX�1��P
হ��=�������w<����.W��Pp)tR0�����XA�Z�u����/k��������/	Vھ�L�n�}�w��MQ���Sl��I��k�w�?to�z�r�<ϻ���M�΀T1UR���o$�е����K�&Jr��nv��(-�b�JA%x�N��}���V�QG騩Ϻ�����%�n�4Ҳ�[]8�3�p�s�l,U�CS��V��+��k�@�쉇�
W>�^Ce����i�j��b|u��lB(�}��r���G�X�hRt�.�����0ȇM�y�dB+��͓�ל�w��wlw�94�)I,��+33)n76n#떾L���N�Ro!���w�N�k���b��+h����c�����B=���R��h]ϥΜ��,PU�e��7O�w8uN��_��ɳ����j	FW����OuV0��mi5�m��A�{q�q:�pvV2������6�.�qLV�+�^�a����6\ T   �>�kRg�nWjWmb:=Q5UT�Iñ�;�F�te�l�v%��l�Ը+ܦ�m�l+(�����f�eUP���  
��U l q_���� <Vڶ�jPVR�Uz�w_��ݕ�YT�.W�n*�����n]�-�[r@�HR��mr� r`�^[n�v�~:�y��k�J�?{���_{����0����F��y�z
��WC�M��z�2I݁���_�"�N,x��+[�Ф��r��m���dx�ݢ��i��r��JD�6�Kx������,�ٴ�)e.������K�)�*v��|G�����m^6�%�i��+\�Hdx���mC��7Z7�Ȇ��Cw�p��i��E6Sd�HX���vYᇶ㛱`�=���T�,J��.ʡJ��V��RL�XX�CN=���(����q��(�(t�
v�s6�C�5�^<K.���I2��!���s��]��>��y�:E#L����wP��q�.h����|\�-`���)����#�N�mC��WS�2!�܊�6�8i����E,��!_-�c�L��<�kK"��o��x�=>�Fyh�3N���h���.	C��S�.gT��(l�D�f3;>�׳�MZ�>0�Q�nO=��崲)e.����xvD��&���]�&��&�k�-��gZ�������s۵S�\�.�JʷdᏝ�u�����b�a#�e.�mC��WS�2!���y\�<x�P�8��:��M��G�)f�j"g��8�=>���h�3N�B�*ߴ��!v[�� ےP		���'�'_f�1���6#x���>!�O9�G���
��ӓ=1��=��-.T��,R4n�7���lF]�4�ݴ��̉,�/�{w_�ϣ/��d�	b2P�Z�ھ�\�u�"����ܞ����f�=Ͻ�ϻ��Oek0L��1ʴ[�Q��%qc.v��z1�v*̀��R�X�vlƓ,+`�UV[��5�9���I�y��ٰ]ym�v��k���帻��-,m��y���k��S[�Ջ]�v�^���U�z�x� �!f<M��8�-~��V�0��\L��P���"��å��/�o��>M�$��o	�UN��:�Y����Y���fE�J��H�4�ˁv;�_q��[m������h�Y�w����P��m8E!�CW�a毴�L�C4�ݷ�����߽ߣ���&�Aqf��pCf��wϛ���3��=�确��R���͎gC`�k�S4'��[��=����u��M/Vھ�Ml^=$Bώ���p�!dˌӦ�a��U]+�1}���7������o�dC�\�NWϞ�׻sS;95��a���E-��e_S�+J\�^�O=�-�ӭ
F�K�ci毴�`R�h�i��m�8��Ȋ��u�����;��}�_����P�!�ђ�m��|kh�k"�|w�9�x��R�&��%���Dqw�Z}7���ny�3N�d�7�|F�(��'}s3��JCH��5���[tny�	�,t��&�����[,���UUM�UV�0;H�Z�8�h	2([*��Ғ� �*�*��`�ڍDK'�{=�u�U��=�FQ��X��ٔػ;<`���U�xu����g�����k��6��Wt��6��Ul�U l d  w �� *�o欯��x��68�6��mܛ���x�6��J�ۮ�z���0/=\�--lf�@�Ues��&Y:v�U �����E>?��t�W��h�w�L=��崦�#M��1��P��z�{�31���*r��Mg�jz}=�zv2��.'NP��=X�D<;�^�ʆ+���i"j�)��E3Wdq��	��U!�sM��-|u��j�qx����V!¢F�'�$�.���Ga1���y�Ȇ���;Ǜj4�!9Q�w�L<��崦�";�T���[m��IҸrЇ���)i�n&!eD8G\U:Y��Ӟ�Q��L��34��-K.$�D���p��5���\j��d m��QZ%��ˮ�M�v�J�M���<x�UC����9hnn1ZU/���!��!������g�s��A�AcI�f|Pmh��D8n	EVˮ��]��Gu�O}yFw����]	%1$6�ce��)�vS��]sf�>�-����0�θ��//�@���i&q�i��m��Q^�N��㦹�M��C��7�g;���,I&Ynz5Ec@���o=-6	6��E�y���!�s�뛙>����"�F�T�]��{S��~���]$��x� Um@*�J��X�6��Ie��T6]eִ��6Fb߿k�Z�;)���F�
s��0���ǈ>C�F�XM�M� �m��a�D�t�y����ӣ-�ʇH-M���"�C��\@3��(����T\�֮rgי�+��rZs��o��  0����W�$CM~���}����}�m-���UaH��.a�n���h��'wj�Z���r���&����ٟw��'�bڊ��<ţŕ�Ȫt����,e��P�j��^����= ��a1�����M���owsrܛkE��Ãh���5@ ;��L{����d��ҚO`�L]CǇ��n2�0��nh�Ҽ��Z�!⫧38�!��L��a%�cyæ�^؆�Q��<��r����p���yv+Ӗ���)8�Eq��,�q��C�-�����;�x�|��(M���N�/g�l`�KAdh�u�ϣ�=��(�3h�Xf!��pOU�!g���V<p��u�N�$�&�l�CwN��v���p�כb0��7�=<hy�հ��舨�x,Kx=l� w{�[U�`P�$p�($ʴ�VVU��H �q�e�-��SU��ú�O�FU�xf[Z��� uE*wP��:?c��SH��RM��@�kmC�ka^h�����G�Ǣ�1��zo�+��\�4I%�y��a�֎�@�J��":��^�޵ԯ�aZ��ްӖ�;���$1�.V
)�S]�W�s�׼��4�ܤg'p���v4�Z�[Mp�������IeaM��G��v;��V.���X���*K�.*񘆟���u$]�S�S!�Րv7��tq�-�T��WiF�5l���R��Sdz�
�^��h���wJ+�R��wgt � 
� w���U�i��\ܫ+*@*�T��<<�m��Bs�D92ͣL[X��f�bmLr����c��pUm�S�6��d
�J� ��T� ���� �
���{�6�ݮ���^��*���Z.�p���Z������+���;�w�U��N`��@ 6�m9�=2�A��Y��GC���cN�BuqfD<uݣyæ��ն!�ջ������/�Z�O�5
�aM|=W���CN�Frw��
��Ս4V�9�jXH�9KF�h�^��n}=�+�����,�:����ޖƗ�� ��a�V�k���x���~䇼m��BuqfD4�u�����	6���$�[�v�e����}��ɽQ�l)�����l/�x���Vo��������GaImPl����[@�}�ŵ�bM�s)� 
�oen����%M�]Pv4�Z��{�2!��|�r�Q}c��0±u�]�/~�`�l���������=�G��ѧ�8=uh�=�Ɯ+P����f}/}�>2�*�h��o��x�k˾"Ε�6���GN��J����s]��ɩ�~@#l�qP��Q�4���ƚ+P���Α����/�&�WåZ{1qm��Se"�%�����DoKb��_	��F�1�s�=�=��tC�D�t����k��7�y���2qʻI��eeZ�VVU��l�z�%�n[c2��a1���/%�y��G8�i|WW��5w�Y��\��iM ˾��Y��I$�X��t�t�hʳ@gǅ[(�
AS���m]Oj8=�V� �Ց@n �zf�%��.��Řh�rح*�fᆴ�!ï�<|:�g&���P$1�m,Ɔ=𨀨J8|GK�h�D>6��눳�j�|u�ƌ>!u�ce�׬�Udh�d.a7��﮻73�:�R�h���v��
AS�g�p������%@��*��8L3v�v�ٜ��j��\�d �P����ol�K*� �ƺ߮gc��u雀��*�ߩ�"l�@3�E�I�N�$���ĵU�\u�Ϧ�J�! *�s���vzz�ǙX�0�A5a9��	)�7�qh[�\�V���jV����e}�dy��O4�aa��/3
I��vڸ卅/ў�N[����v�}�αd�8��+a;��k��U�IP�U�����=SKju��M)e�4 �T-�-kt�;c�tlHtl-�PUu��Wq�J�o3		�V7���vr�x��s��T�z\��y�|�q�HجT���^��vڸ퍅/ў�N\�mSj(�a�Jm��o3��j��/Ƒ�	�NƑgN�K:� �G�bp�Y�4���~d�e�P	��ss;9=��n�A��K]Έ�fϻ��hi��)VäB�%�Iq�[Ę-#�f�F��[�� �!qT�Y�=�u�A��/VڇH:��r�-���cn�v5h7c�Ź����m��{P<����n �z�{�vfP�;�ST�w69mw@*�K�;���qT UP���D��l�Ͷ��+R��-*�q;F25�r��ګ��:=O�v�Zڭ�Vc�G�
Z����wk���V�eP6ʪ�����P+( �  l qT 
���[o���`��V�T cq^]��θ�ӫ�z���㸫�{���V�T p��wl�Wx�ʥ.c(�m";fFzkw=�l�!s�Y͆�i�� ���B�B,Ç��� �,�}�H���m�i"2!�꺬�#O�A��H�H�1f]��9�J���"�o9cH4��h�a�ka��&�2��a��c�x�=QV�;��QeBh��x��	:��n���S��2�v[#�7�7&7
"���5}��-�)ӥ����VfG$PX���rf�w��cNW�[����71Ⱦ��ɥ����O�p�=��#�ʹ&@T�V��j���@�k�5�!��
�ڨ63@�Q���ܹ����}ߛ�me^��uxm=W�E!�xm���6a��a�hȆ�1"�0]6�m��ka�t��U�������"�aޡ�^e�p�GO����z}��X�FJ �*�g�3�S��~5���8C�P��j7��"�O���9fռمa56�$�mjZ77Y�Ox�K|���)2�|����<3�Ś)i��c�
E�у��� �Z5+Mz޹������5?j6���P�Oz�5_n������]�5?Owg��V R�@0�։����x4���ܡƼ��� T6t�N��4�6���<���?��~�J�_;��0�cz�fD<f�ZD?a��{+���@�׽q����zj���Μ����6G��]���"���h��zc���,��ƒi�3E���6��NP��^N����[:��;�OM�zO�a|]~�*�8Fcy�7��������Ԡ�ym�(^���1n[{����&�[y�Zx%�;����]KڲsT��Jt�~�b�[f�s��M�����-�-0QVդ�� Y��F�޹w���� m�� d�����[�m�Y6j'�}��zdtc�D"r��pڇx���t�~���<��b��nv����F�)��E'V���X��u�;z�޼�ip|�S�,��բ����uq43�]2鶩�
��=�n��,5��z	����i�S�g�0�P�%��t�~5۔�%D�M��)�_�$^,d�V8�O��b���NU�NT���mQ?�3���/�1�L���n��=����rܬ�-����V��L�kt=?zjS'������J%�5D@��^B�t&mj5�V�*;��� T�Mv�b��b���2J�g�w;3�7��6�|�y�O�=�%�!����w4<��N����K�	=��PR�em<"��įӺ����)���Bb�!�h��w��9���beM<i�#�|-�[j�3m۳�0�!:c�zs[�%sm�I)%Ŕ�m�B��&��W��#0z�pȇ��f:���v�
�4�^li*d���
j�u����ý��zve�$J��j!�+p������'��#���$ � �! ��H�  �[d��FO�[$d�!c$CHH��$			:�I k�������	������������$ ����_��������� B	 $"H�0H0$	! �O� BI �?�� $ �������N�?���@�! ������	��H$ &�@�! ���7�;�^f� @��~� @��~d�������$ ����?��nh���a�������B���~߷��PVI��PT�w�\27� �� $ ���`��  � ( ( � h 3�Z� ��M6 �Y   P$�0�64��)G� 
(�   
  �JA���E� h P   	
    �( @ ����  t   ���=�w��:6 3�����O��l}�} ��>�@���C���@qG�   ��  � � y � �mB���bsס����}w>��-{�zV�s��κx��Z�� I     ���Яr�+B�7;�A��=�t��m�|���]���C��N����a�� >�*{��/���޻ם"l�{n����:��m�ϻ�5��:����&�ֽ��{�'GN 60�m{���Kw��P*�    @������soY�W��0=� �@��7�f�度��i��K����k�n�k]��ٴ+�� }U>��+�����>����
���<v|>���;]�j���
�=�]^{�
S��@�� � ��z���wCE�8���B���vw��bj�j�wז��1�b�CT���P9����w��r�=hx�z�Y���֙�H�����Uu��Wָ���qiѯ|> �����j���UN{t��=�)|�P(�  � @�>��J��u�qz�;��zq{��h�C@�-У�it8��WÀ>�r�ެ^�zӋ����z��x }���Z�o{�T�������z��|^�������;{�Z<m֨qwj+b���~M!�R�F   ��
U2iF�@ �*���T�FĆF ��@��U*OI�    ��5I'�UP @ zSmU( �  h�<7�߷������v���&n~}�<< �Jb��k1bĖ$�%���f%��f,X�ė�K,IbI����ŋX���K,IbJbĖ$�3ŉ,I�?���[����V����wj4��}��Hun��ȵmkc�a®�jл>�V%K����'�P�XB�4爥Zb�Y�qY���k�Ka"�Ս���r��ժ�)~yx��N*�h��"#n���[���J�ּ�]�o.5�>ڨ5o�˕r"�W��D�٥��Ey�X��]CU�.��ٴK����U�B��b��+0$��4Y%X �|���L�)�	�y�.oN�h�w�S:]8qa8E��
9)�^���eogf��0y6
��e�/�c/=�eHe��c}�dp���La���_[�{�mk��*�,���X�Z��SP��#���WA4���d�z�Z��ͳ�FX����� Hbc���M�>�ן*����>������O��Y�ǌ@��TlۣeǕ%���Gu��m҅���e��Nj�A:�:�n�����i��'������b��L�)��,�Ã��-R����4�����T����=3:�����{��FckF]V��/e2��]\�88��rF�`�'op@�v�BQ����R��G���o��D]��-��H[��yt^��˛�MŖoq���A@H�#Xk-��w.�OhüJ���C)*���7^-k[3)�uwl1*�Ϩ���;\�j�
�P��%�
Q�8=uU����/*��$W�h.�[6����"�$�IG�Ĉ�Pe*
�`!��b&&c����^:7tC�tv�h�u��6�1�cISeԫ�u�f��6N4���P��6��G&"h���څLn�
�lw��n��TN1~,+ce�D:�w\٫���I�����ɗ/vѻX/��E�xS�W�=ƌˆ�B���A��F04P�:hāR���E.8�QǧYB��fe�i��["=k��̒ŧU7O����p=	��Qu����`�y�@�^UN�rEH:�����
wx3.ӱKu
5����&]�v�oP��h��40�i�Db)���t�D���w��Y^&n��R5M����r��T:.єUTJ�{p�`̠�\ǾI�l KL4���������p��f�ڊ=�@l��6eJi�v���k`\w+[!�4E3j�7dm�!�vըp����=�3�2�طN�4�Y�L�u�Utᔣ������pV'�p|� �-"A$���XP5�P��Uu[EK(�v��Iٻ��$�&��;�!٢W�7��lTa�A����P��J4lU�T(33me���u�1��/�|И�z�˴Z��&��کD
 �@�G�O�)F.Y���W�Z���+�c��Ĵ�Y�=� a٦H��SHUH���V*ah��f?8��@�&���	6���˶ˁ]ȭe���d���%0R	�;�'� ���Ģ|@ʤ�xg��:�f2�g�8C��h� *�5Y5bY�)��� �a��yj�]Q˥�EVf{�yVb�n��h�0cT���A����a�G�%Ypc8�F�D�
7Ik�i2��A�m*W����#��g� �F<LI0Y���i����7�W)T򻥵C*��4N#I^l ���*��^�|�woJ��'�;�dѳ>��̧Bz�b$|H"�(���۬}�%x"�> �I��� �@1Q;i��%���	D�C���9�!_�C�ꮖUF�����2-d�	X�nj�Ulb�#�1�է"u$(��ל<��
B��R(��]hW�M K^H�E`A\l$�v3ښ*�`�M&��v����h�^oj�V\���+�Z�ʖ,� �PT�If�B�w�^:��vr$QHQ�F�y$!�:l��2e#�)a�@ѝ�k�\�"	�d�#��r�+,���j(Y��$���n6�$�y ��t,;/n)��v��ny��j��:o4�=2�!)ʼ�$"�Hh^��|�P�(/5I$%�C3*�H@�`��1^7h�Yu(J�JS�JC�b���L6Ȥ�=1�w�v\�s(L̒�E�>�f�;��k'H�i	H�:��މ�*�<N�/(D�����I��ͤ�a�1�!���a0�4݋b�ƝUUТ�{���E&º��d�r˚�L3D�EFX���6�ɖq��E9HJN@��0q6���cb��@�0݈Ҳ�U7a̒�ha��nx�D���w�Y��7%r͒�G�7n��sra�h�mB.�U���1
Vh����v��$���=�e��?	��Y��;nJ�bx� 	���Bq��d�61��G#P�����*���N���q�9y���:g#���#I��QI$R	���f�:�"q�=F�T��9���m䬺�-�<Hk!Y�M�|ɟ�ذK)8>9�8��}��|M��Gr�x��&86I)i�:�+�^Uэ�	��Lڷd5Jy���S�CeMY}ւ�ȥԍ^�2�
¸�3���(q�y��cȱ&�Aq	�� ]�x�m|�L��q8�D����gNx�YR��]�@�7���^�h�N,�`��A�>1�	�3b� @ŏ��A��b�fb�01,H%�X��%�LI1b���,Ōbf`����$aMk�%ԧ�W�g.�p%�zM�0`���c-`��Aw��i^��r�����v�%(^d0�G��Qu@lM���"m1  ś��w�n�x𼇸^��.�}7}\�k,�fP;���t���2M�G$��3%L�/�4!q�3
L\�t�>5�%�3�@��@	,�&�Q��e11��f$�����13�b�r<��b@�2��X��bb�	1&��P�M�ӏ��wނ��9SA�x�������b>
 ���q���R�X�pz����
D<!93PX�1b�f(Ƴ��&�$���	��H�1�31Bx�`,��!��
H(�����s�Ye�M O6��Kd�I��1F#I�cl ����o$#	!7�ܞ�W<�Ŏ��)��|<� �I(BQ66�X c�6�i&,�A	<Q�4��5Ka%(��U�Pt��#fg(�J��� �����I�Ӷ.$D	1��E0Q���!�q	�� @N��	���X!tM(64���c�6E�-M��q� B�?\U`��i��bB]�� F4V�b0A-����m�m�)�Wq�-x��e� �0��J3��蝇ӓ�=�w����D6!A����p�x��q�L����2S>H^��hU�1Ci��R1(FZ�M
^Y�h!�%i�ܷ��S̟�����_~3l�Nbz���q1����o83�pI�(Tp'�Fc�/��
쳵�UA��E�y �J�z1�`�t_��[�&uT9�K+�H�w=������P�fG�s+.[�:ո��}�n�irR��v��@���Ù+לp݅���[s#ۂ��aʲ^�T4s�b�xM~�!^F/'��z�`��������BK�%��ɚ�GuX&<N��Z�ŚX�egP���c�v�!D��$�� I��D�&,K@ &bb,e*J���K TcN8�y�1B@	,"X���	f �!1��(��nfHFq��*&H��HQ��)k)S�)CV!NdbH1��H@���R��,H
�1$�A�/meI ��,���b#ĩ;"�K0��6�r,��%��H,����i @� ���X`����,A��'��� �h`��ǀchhcb��;y�yC���e�e�M�����<���3JJ��C�5]����1(f<H��C�N�	j��$��X�H�q�\6c��j@SA!#�W� ��CL��F<�lb#3A��$�i  @��@ Ly����#$�тo�"q!�7�!0"��`a��facW�EQ.S��jp*(�"
~���>T�Nq�g��1D�hh�����ŉ �a�A��3 M��nH��\�q;��:�b:��k%�IF؄b� �rH��$�X6!��! �$�@�ŀ� Y�j��[�R��1`$5TL�Ą$!$�H33'3�9��� o0��cIHF#Y�6�LCxXɈ1f ����Ā L�bY���,� A �h'��ř�,I�0a�Č($� A��Ŝ310�����hb�f`�+`�,A�F�0B� �hƌ�6�x�1�<��H3�$�\倖C��H3 Q��r/��]1r5�� C�"4�X�J^�;�N� łm�bM���K�a�L�A
f�aHR�IH�쑾I7Zp�9��ށ�U�T�����$F	i�(N;��	��IB:�Ƌi��r�1��nbb1�0� ڍ��(��������i1qٖ0�M�	 @�b;fd�g�/�ؒ��C�W���JW���J潑�@��2�DnÍV��8��;l��V.���
�hpi�#��N
 �
�b#�J� �	��l�aD�A��)�M��;���5�Ѩg����<%�T��eгK�,��6�b�LW�|PO�8@��4���1���$>�-�I�Iu�v\ʤ7�3	�{{mr�kvLB�uX�2�mP{zH���*�5BcW�*���b\a@�6��n^� ֜7)�1۬�UVU�(i~�K����R�!o[��F dR�Z(5��D,tT��&�V��n� GN�4�c����76�m���j�U�4b�]��N`5g<�e�gu�\��kL.��{ob�O�|]�X�v6�Mӆ����7�� H�K>7��	`��������O�S,�Ĉ^@��jx�F܉��}O�]"P1���XA��1,P�,�6� �`��@���b`��fOm���婠�9x�4]ժ��s��:���tӹ�f�DT)�j]�'c���+��j�*�>���Uxs�A�M��j���u^��2��	o��6YA��}m�	�b�iA4<�M8���(~�8)�>��&4�`&1�I�	�( X,��1!�>���Ul���R��Jw�T7�����XQ�����?s�Tb3%�q̊EBxă Mc���iw����m]?={{g��z��^���CAF0ܟE�b�8�r%"	ڠ���!#`�H��01``$�6������ȁ��$Ts�W�Js����Gd��Fm��0(2H���� BF8�]br�	����a21����"[�:�`�f��Wwk0b2t�a�6u=�bI��׬^�tT�n�IA��*��qUU!Z�I6TG]NDtV�[�m�Ꝧx��j�+ƛ1c��g�4�2͂M&�K�E�ǔrA0ZL�0�b��b����"�����%mLYz��Q<lEؔ@�X��U��Q�=C9G{J�!E��A�</��9�z����d�H�PGE1Â�k�!�t^8�ă
�:��l�t;Qn��Z�#܋�/�MZ�~��ϘB!%?6a�1��5bTm:�!����LJ,���"�c�6��N�	�&ݮ��C ��ʢ��{�����j��U�#��S1�I	�
ZV�p�%mJ�^6�T��,�T�ӽ�Z�ge�]�f�]m� �U]�j *�&�m�k��g{j��U�E� ��ҨJ�.j��³��c96wB�\����,�`�{W�`��SYֱ���Y<�C�UwU* m���l 
��ˤ�� [oS�@*� U         *�      � �      VPP  �@  ��*�X}�*�QYC�MF�N�ŰmX��Pn"��w�l{���������e�
� �Tءw��UU�lR�Z~�bSԩY@ �[���@�Wu��D� �   �m�W�����;��     {�-��B���;*T��zap0  *�T�m�wV�N�����2��yCb��)(�(��
� �PY��^�� �1����n�c<y����lsUUW��کH��FW�]�h��U\fF;�y]��Х]ճ��gs�S�E
{�����s�]���on �:A���*��qC-@x5JVúxU   x �0	�   ' c ��n*���;��p0  N ���  �` < < ����m+�5     �        CqU����;�Tj������&��d   R�A�ݮ8<P 0�     1�   ��^�-�R�� *���    � � �      P��        P 
�  *� ��` ���eU��� ;�� =T�@ @<U n C�  [� �����ں{ePb���y�OU/[lʪ�����Y�ҭ�w �-���@ ٝ@�T
�b������ $޵��
�yU�h�,�T&ⅠR�   ےUK���)��6Ͱ� *�rت -��� ��U 1mnwj���TP  @ U n՝��P�-�         �6�  U�   m݃���*�lw     ���   /R�l^��B�                      ���3�
�     *�
��T *Y*62l�U         ��M��fʣ�}��U+�lh 	A���U+         �P     �BqT �aT 
�b�3j����  wM�1��c�������.v��mU8 /�!୽f�ݭ��n���Vd�KTJ�;c ��v�	�E�VP{w���3k�����S�і��o��U{����Z�=*�*�oe���Ւ��   
��   *T  nm�� �@*�P�\ʠn�^^�\���,���Q� ʢ��jl�6˙YE^�Ӱ[ m� d*k�Tڙw9�lPw��   
l�@
�ͳl�jW&UV��V��O��9,�D�A�*Y���띜�v}u�7,��]f�7jU̺�1u�ʛ3�R��|pe&F���>�mH.觧e�m+8��'�yv˶�ؗ�[���,�c��}��V�E�ۢڶL�Ƈu(�,h�{Lh�c�j��Ʃ�TF3�8;���R�ζ\:n�Q�V)�"n0㮱�ZvU��A�!�!n%�ƶz��(/U,���s�+=b��3��Ɛ��]i���G��:�d86Lm��@���7RǷ`x�g&���ݹ�A#��,��\�ט�;'l�[,�c%�aucf��ۣl�"p���l	�Vְ�t�e4�Ycj����j��F^��n�9��=B���U�1�^;���cg�ַ1'��$�5�]�Q�+�VY@8Ѥ,�gx�㓚��<[)������1<i�����Ɍ�@��lX�U��0���\� C�xwz�kr]�wv;�k�9B�ͭ&��K��d9�k��T�FI��:K�6w\u�y:�,U�0e��.����,PKSS�-���#l�Sv�1��)1۶,�+��tK�Ri)eLԁ�ɋe[p�5 +
�6�1u&��5��շX���*�<��Ȋ%����*fR��-�v��a�t�Mr� �dx
.d� R;�v�Vnm�}bck6�Q�nƍV�E��@n��w�2�K��`9#����l�Pl�Ǧ8���N�m����͹��Ns�Cd��ͤ\ʑ일�Q�s�%��wi'i�����A�i��ѺHn�/j��F��.K
�F����A���u�ŌW�:z���|+���}��k&rr}���z���t�sٍ���\X��N^n��q�֩ݽѮ��gɹ�n��q��Ü]����=Y�x�����ۮË);�6=��xS=5Q��&n����ӂ��=�㛯'p��nt�T6X)���N���cO,�Lib��b���/7T��"n��n��μ�h����.�OQ�����C1�E�W
L�{��X�"Dy��50�6�G�A�YE�s�[�[��r�B �p9��5ɛ�dV�u0��0M]LugF4j�s��"kc(������AZ\��y%���,Yyt[s���ڹ��{=kf������u��!��m�0x��v��e1��a�Hp���e�4�,;h6GF�&��Aϋm�l�ge�W�+�e�� �c�OgV�e������|�s��c/0n�e����v=<a��_5�-C6l z���8��,�m�(��;J�v���fA�MI�����8+��ɖ��F؛�+ā:���B�s�qrZ8C�!�#Z�ޓ��<�������T��v�:q\��bga�GC�`k�����ȫJ�c�`��dLT۫��pa;g�gE�{1m�<s�,d�7ks�:s���c�C�� �gn�0���赵;a�ݹ��e�7I)���3�՝Usva�Dܕ��r���i��U0��p�{�qM���m�u��@�m���=��j:��*�b�۰�L�q��5�w��Si����rb��;�f�S���)}�����7�&f�i��T3,3v3	�i\z�5���N'���7U�;[�:��F�����]��l�}��|lYԛ2�9T��Q�)��q�R��b/�om���bZ�]�	�;e����ݦ���3��3�/�o���̙f�M�Ϡ���Tj@�)�ݏc�cuM���nG�����X��>B5�ۧk+�vW��:��h:�����PY6�J=<:���#h�'@��mo���.�-c��C 7��;p�g!����K͋��qmɇF,���m+*6���Yg��1����j��W[A� M�r�f�
�q�M k�m����tβ��Í����]I��6=�����8Ջ0Ԙ��:g�u�mg����DK�\��y�.�jxv�+��k��;�0��j��IPB�_(R"
�
�����z�ٕ���l<h@U�����̵֓�gPn.�"L��Gf���d���]P�w�|��nL�,���9ܽ`�nq)�ε�%�$�������'RF��tn�"�O���[p�m�.Y�z���c�P�^]�X���I�;�cQ�p��R�eې4�ɱ�wc[�����g�:ݝ�gY��ɺ�jL��f60Y�n�sf�����G����"����;��^�x3�����8�C�w"�Zj�ŗg9p����bpV�����i�L����J�n���e��g['ns��Uۭ���kF;1��ZK���
ɧ�ոlګ���cg��n�U��ڱ˫�N��cu�ɭ�4���N�;x��M�����B꺍�nV�n����hޝ��\����-�a!3�\Լ�4�<Q��۾�i��c��7�H�n�,gn�.Z�nh��M�FN.���y�i��M��#v�Z��r��ڹ9��9]t�\�bΈ�0rqpumӌ*�B*��ħV�/)���Y�lVi�����u�J�K�j1G$�QB��SB��|S��۵����m]�x�x�z�2{`q���)��qVkz�v��qd��g��G�Ev#���q��,c]M�P㤎H9ڭ�{9�������tnNd��Q�a��o<�s6d6[+��na�1��i��{+�m�G��S"�c�g����d����`A�:i��V5=��E�f:���72)�;ug�Z�a�0mɹ���3��y�Ӣ��ָ�+g&��NNK�����%X�:4�6hG�ƴts�wg�6q����.�)�����:$!�q���猖�%�u��(��s�$L�xz�q�H�l)^Nƃmc��m�]ې�T����(��S���Sj��ڝÌ�o�����?k�`;H5eحLq�A�n�퐱��b;����S�C���@��6�����c�B΋`=��䊬�l5�X��.���F�m�F�\k'm��ֹ���a4Ƒu�F�MEm�s7��p�ifJ!�rD9Lh����6�n3�i�Fc�+<8�\񺲼�N�;[��n�uʹۓV�&δ��Õ���6��`��/��lkr@��K��Y1�I޼[���9�Mѱ#9��g�M��j��f��67v�ܒэ��=p��EG��)�f�qϝj�-g�Ľ��av�#�C#��WuN��mu�.ִ��E�.v�� ����v�萉Mb�7S��s]�um�;���86�V��^7b�gc3��cO�:��p`3,�:p=R�@s��"���]GI��q��ڠ�fک��˴�@ˤ�Zj��vc�����ݕ�0�F��v��퓂�NP1Ι9�AFT��i��Tݫy\���2K:������h" �K��bpW �Z�U�����T�sf�=�����۴�f�z�zX(�y�a:J�n�Ը�iR��.����)�Ų.�˔m�I,�r8�m_�Y�$�%�Y�X��9��,I,_�1,X�Ĕ�H�g9�w�������c�A��t��$��VȪUU=�6E���(�v�5@H
�P    c 
�Pm��.��ʹ�|�ʨm�QT U@� x*�Vj�V�� �/g@<�k��u��{!'c�[ ��Sj�H`p���G c[. �*� `*�(��֥P 
��
� �    ��l�*YKeS�we��
� �UCws^�6 �;� /UT�P �� � ح�T��`U    p �ʩe  ��[ 
� `2�n  һ�����&m�ڌ(4g�ћ
��UP  �U�Sc�ZC�'�U��׍��r����a��۪-���	��<=�vJ��j����t���-B`���a�rd�mښ��^��Fq�]��dX�*s�9Mv�����Ũ��Z,t	���Mmm�䡅9����l�:��Rc�����_A%LwnG2G;=hy}I�5��vn�<rvAW6��
�ɰ���`��C���;<�B�V�ͼ�C5�^Le'�Ol6=n/g�̽�T�3k��$D�h�Y��Z�l��&�n�۰�WX]�\�(�)�jҙ;z�lg�m��Y��n ���F�y2�ݴ��	����]���c@�i3�������&�8]���[���X&a�Z2$��<)A��O-�cE�nS��q���4�N�U���be�8!�e�hv(�p3����{u�c2h�o۳��[v��a�r��8�q��%!n`�B[��zU.�����fP���,v��\�/�����8���M�i�����<
��6�g�����hl���úS�dm�z�Xq�=�[�dT� 9K�r�[����Z�6��cC�� ���,WU>���ˍtI/=K��)�h�T�Ӷ�p�y{�$s�%��8=6�a	ɵ���d����Z�k9��7dl�;���q`�@1c=�1�RhM�;�����3�"V�]���7+g������x�%�3l�zV�
:���w{��(�g�胲FG]�Km��
:�lz7\ڀ��G'͊6͵P*WD���� +m@�˹K&V6��9��*ԉ�·���8���Ug�7E碛�����V��lR<sxM�8�\��"�	\�p���vǣ�d�^���+I<���&L:ѻJc���]=m��cҏXO'gqƳF&Tl%�"M"Y�9�:�t;=����ݶu�XB�К�{ǝuˀ]��l*�m��۳�
�x���g d^<��`v�����Q���
�3�ݠϡ��Su
��īW��T���Ն>|M���B ��eƩ��Uޮ>㇡S��8G>�g{P��DU�>���r��2@T�"܄(�
s��8e �g�K��5�9�5��h��M�j2"���hida�6�t�rkh:#�>��[Ʒ��ȳ�W/C��{��(�ق%�XD<@'��\�Dޣޮ>㇢S�Yl�ԵM���;��?��jٷ �*��S�N����H�<�^�q�p���p��wfRf�RZ�KQHP��j�p�O��&j�,�5����2�y�ܲ8����R�����6���*5�>�G��X�L�:D�]8���Zw��a��ܫ���å�/����pB.B�rC����Q�<�7T!Q��Wq�Щ͌�ӄM�I���mWw��L�<}��&j�"�U���锃�����~�-?�Va5�!�M�xO�L��݄�#��cłE�C{����ާdq�q��j�А��I$�]�eev����c�I�'m�k��t9��[{3�fh�ڗg�qΕm0WrI�gZ�C�7h=��XE"�G��dn�BU��"��(��it$�jF�"ɑ�]k��a�+WZ�P��q�3���8�B�� C��^Y����	�A�f�\�w=��Fˮ'�ܙz�ZE6B޵rdq�%�8��]�6ځ��n �q SR������TL�8�rh�1��"Αd#��7S#%��D�qA	�d�it��1�ɑ�[�ʚh������q�;y	��w}���N߽���N�ҭ)2��KՔR�����PKn.נ��&{h��g!V)�Hփk��Ϯ�^X}Ͼ]�l��0�]q>0�����`��,�Ƨ;�#��Zo�I�l�"�LĤN4٭0�k��8�l���ZEDȣ�w!Ə#�*�,�Q����������Dw&Bqoz��tٜ�;�#���T�G�O����#�|-s*(��b��ZD�ȣ����#��jȇH¹u���;�#eQ<+H���[�$��*H�-�ɑƈ���igH�U�͡������TL�8��h�7��E��ӁG�@���Ju�=b��{6�[���&�ѷ\z{d�p�q��Qd,,�dVG#K��^t]>������A��Ѧ��t��Jsɑ���Ni��V��v�qĄl��e!������я6�:B��"�"���r��w&Gt�Ye `m�D��%� �"Λ<jpc�28���Y�.�^�dq�q��7�iG��Q��-e	k^8x�No�,�B�N�#u2�[��!�fr3��L�8Bi��!�* �n6�i��V.2�COƌήU�:L�<ƾ�Y�D)����(�V�ma�9l� �M��H\�ܺ3N\-T]l��K+R�����iUPw ���ʶqQ�*NVW���z�V�ۋ�uY�Y�I��� AQ�Q]w7��kc:�<�i�=�G%��:�Â�x9��[�ukOCq����9+iʘ,gu]���Q�6���A�Ҹ���,��1e�i˲V�ε�-ǯ��u�g���/
�Թ�Su����Z�Wi`�b	䌊=��MtZ��[R���\B��2�������<�Ű�S�Z��EG|G���	��˔�Αv��;#�={�X\P�fG%����V>���sk�mm�im���Û��ӆQ�}<g�J�f8Grdq�:�'4ÄV���COƌɽi�"���C�<h�ں���
�
��-�s���)�Y"�<��N��.',#�+���"�:����l��ِ�!I�8�8�[[´���Eb�C�<l��xՑGH��t���ᚵ�="��]ڞ@*Kn�O,�D��yq�i9�3��/8}[�,�v嫠/E�q������!Ӈ���o&G"�ssL8Ej�,4�h̛�֑-2(����D\
lm�An�]~�������C�a\��|aɐ���5�Q�dmu8;�#�Oyc.4CL��$��,�k��8�8�ڛ´���g�C�6F=�UdY�,��r���r�B$�4Grd94��qt��Q�ɑ�[��Z�+	<G+z��IM�=�V��2(�|y8�ƈ]Kz�!�0�\�>,����Uͪ���ߛ�~c����1@��VV��<ai8�����>.��ۭ��t
m�gc�1	)����3Pf�rhl�}�������M,�j�k�8�8����ZE�Ȳ���6F=F���D��H�Yt�#A�dn�B�Y�V��=ENCy28��E�4p���.,�¼�J*5(q�8�Ƿ�֑-2(�\�8�ƈ]Z��(�W.v�Grd9�I�\)F�A�#Q�,�7��ɑ�Ȕ{��Αv�ʢ8�l�N�ZGk��������Y�VږּS���o�Yt�#A�dn�B��o�H�N��!��p�خ#	��iC�,�+l��v@�r��'nG��#����t�;���OS;�!Y��;��o-��ߚ:FZ�,rc�#�uܕi�"�r��c�<h�Է��"#�a��-X�BYQ��n'ő��j��ZE4F�S��28�CxM,�k��G�����͸�I@$$�������G�C�6B;Uf��dh:l��ʆ�V����G덋�s6.]Eĸ3����7��4��+S�x"�Dq�2oCZC�æ�`��t��lL&RA���qHԐ՘t�+�\O�#�3���Y�DN�0w&x��q�Y�.�]���ڑI�#0r�T����� ���:pFH�L��xN�|��rv�i��'��p�8��x�l���ZED�|��4x���U�:E���7S7Gm+q"	�F�,�#)CZC:p�(����#�`s�8Ej�U��4G3'tU�KL��Q�l��q������1Ş4B�ޑU�:F˝�őܙڪ�itН��_y��D���JVR9%-m���:E��J��#����kHv����uu���U����j�"BIc�z�r#ޘG8gB�����wL�+��"�o*�P�Dq��Ԋ�P�m� ۻ /TP��{a�;ܪ��;��6ʶ�U,�(��W�m�Up���oY����/�+.�g�s�����/q���ݵg]��΄��g!�vz�۬)�q����-�#gEC��sq��c�y޼f��ml��9�L�G=�����k�EB�/����Z�7clNgl�]�i��{p��n^;e4��Z%°�����R���V�<�$�EC�M��uF)I�z��6���c(��H����+��0�L��c����Wpä)�4��i�0�²�&���l��nb1��b$��U�(�b��صI8|��5�#Ord"0���lh�JD��I9#���:E���3S"1�it��Q�ɑ���<�:FZ�T�|I�' �q�8ћ9�"�dQށ�(qg�����ȇH¹s���;�gd4J|e�Z��"4�0V�GM9�#yx�GxN,�j�G�����5�\L����n����j%U�VX6��l��;4d��8��ö�(��kn�ڸx`���u�1�	l��d��`��G���o�Yt�#A�dn�DsRBit���ɑ�GY7�#fD�"Xi¹�VwV��nM��桇L�d#8a�����t�(�4�6�I(�M���;�#k��u�Y�f��L�8D��gt��\ǈ�e	�ybP��H�PD�"�dQƻ��G���l�Yt�#A�df�ː-��7q�Q�Ѐ�$j4�q�;��5݂>�g7�G���gI�vsg��[;���f4�2�UV���i��^̻���A��r�ja�F��gĒ;<�+Q��\�q���[����t���"uq���:h���Qh�����}q��8�K�h�6WWq�!�D+9�a�dc�2���Q#
#PĐ�`��,�'�H���#�3o���]X?��>��`�H�bKb��f H1`,@�0��0 Xf`�1�� 3H�!,�b3$%�HI$�	!f$$��`�0` X��A�f 0bA��H��A����  Ř#1b�f��,�fb,İH0,HIf$�%��3���`,� ��b	�3f$�bFf ��X��H����%�ś���s�g�ŝ1g�ŝ1p����|΋�X�pI3oft�,S}f��[m��",%���$�T���ŋ��@���T�]oft�,^mb�f-w7�T��X����I��x�2����3���� ��I��bfg��NM����f(� ���g�ОKgϽ��b��P˹���-133�1b�k.�&b���qg�bŭ�@�$��񉙓{�s:,^mbD�1F�gb�����-L��3<c/ͬ@���T�]oft�,_6��f#��g?IS�1�fUUͫf.뎋b��{�2ݔ���x�3g���7\k(B��sո��bfg�b����	��n����X�h�f/���X��wN,@�I3ofx�,_�X�s���K�-133�1b�k/��1{g?!�fi�X����I��bfg���m��Ղ�Eb�s:,^mb�$�P���Ŋi�qb�$�T���ŋ��@���.�bfgb��� ^Lůx�>b�g�b�[X�xŐK>��q�xK:b�	gLY髱ɭ���Ge��Y�1,�?	e�=WxK)�>�_i�$��,Z���I��	�����L�L��X��V�,@�I3LL��X�6���I,	eu��H���񉙜1�o/�I��'���ŋ�k/��1C�8����|�όbŽ��8��$�P��^y���Oo�v�%��L��X����$/��n�Zkn��h͌�<�c3�1b�ig�Y�.}������1,�/����s���8%�M�\Y�,�ڀ�t����@��"�o'bڏ*�UrØ5�����Y�T^�Ol����ݱfk���M�p�UU�]X�uXs}�b�I3�L��c�w�� ^L�L��X�����]IpŦ&fS�y��D�1oIˉ��c-mb�$�_�L��j�ؐ.񤡊�����O�b�K]P�i�(8Wň�>�LK�k/���.�>�b��� ^L�y<L��X�5�U��LL̗��\�y����1x��όf%���9��e�1g�Y}����Il��VZ��Ś%�ş	g<Y>��/�1gD�LY�,��6�ş	gz�d���գ��3133Lb���ul���S/6��f(�wih<�8R��E_1S3Lb�[X�n�{�����%�� _��1x����1b����,@�ZJ����c/�X�s��R\1x���c/6�������34�,Z�F�/�&fs�{�Ka;�Um��gE�ͬ@�ƒ�U��j�-��1t���1��� __iR\1t��Θŋͬ@�$���x����~mb�4�1Q'W8���p��1x����1b��W�td�T U<cT��F�]�1���m��VVZ� 5Mvڗ3�T������\����_UX�*��X��m]Ȝpc-�U^ ��v�En�d+b��+�aգR�i�P:�lҶ�+����۠���'�{�����ڒڗ+7�RU��nX��;�������������-%
a�:���vq�խ�2��:&{l���<[%�P�ɺ��٪���#b�ܺxq�ؔ�	�ݕ�Sq�s�!u�0f�n�t�Q:��7[M�gq��P�LL��ŋ�� \�~��ėL^133�1b�k/�4�1{�~Rsfi�X���D�1t���{��s:,^mb��ICoft�,[f��qb�I�����c.���~z�W%��48DJ��$�b�� ��X����$�Z1S3Lb�[X�n��1V�d�;��gE�ͬ@�	&b񉙝1��n�ň�ICofi�_��ڵ��z�co�((��n&������i"�lO��G���x�"#H�t�1!��i(b���׭��r
���("��΋�X�~L��3?ŋzNk��u�����34�,_6��w�!�%��L��c/6���IC���1f�ŋ��@�I3L|�ݯ�8�~����B�D��8傜X�h�f.���1b�k)����ይ��ŋͬ@�$��^�~|�L�1�mb��P�[�����:,^mb�I3�L��c.zsd��u�����34�,_6������:QJ�e��6� �%7��	�	�-�F��"JƁ��	�=��6ڮ^��D�R�!ėLZbfgb��� _�4�1o��� ��X����&b�bfd�wNgE�ͬ@�ƒ�*� ��X��V�,@�I3LL���~mb���%�[��1��X�xI3z����H
�s34�,]mb��P�[���{�8,^mb�I��bfg�1bޓ������1V�f�ŋ�� S��K8���&ft�,^mb�撆/~�c��3�1b�k/	&b鉙���15�l��d��gE�ͬ@�u�����3:c)���qb�I�����c.����2��b�x�3�1b�k/	&b�6~|�L�1�mb��P�[���Wt:>�rs�#s��XLcL��o-[z�F��WW*\x�6V��"�dQƸ#�6GlV�#�^.C M�����:F��7S!H�it���ɑ��u�*�GH�C��I$��$^AI%U[ �[��aL�sՐz�`n��j��V	'k*�҄��V�B����y�����"`��!�4�Sٺzu��y_q�n$�E�ێ@�2�,{}��8�[Hzd.�9��:�<F�+k���i�Ev�%���`�CE�!h�"�J"���h5���4���֗�f�F�#��dFc	2`\0:�4�ŦP(a�a�-��)�F�d�!d2$���|G���a�`X��"a��'F��:F��1ڙp�Gk�qFb�*����t�[Z��Մ�m�\��7�(&z{u��
��y��6=1����GVR�u��KtQ��-�}	�TEۼ���h"��L�����4�a��nLp���(�q���ӄW_X5�ikMQ(a�a����%&D(�tB0�E��\kv�WR���g�|}�Dn�GmW�H���g(;�#M�(�Y�#H̓���\H"�P6�J-����bSq�'��DQ��Q�H�4Df&q��$���ED�$P��"ΑЧ�f�t�[�iFbz�5���ٯkH�3���F�Q��FԠ�΍�j���Zl��B�.{n�Td�ш��@��������v��t�+�\L27S9&�*��:}��3��jH�7��1yH�{�д��$]99.�5�:Gr��Z�i����L"E���s0ੌM̸�#Nu�����_���9H�a��n�Do)���E��G��9���6Τ[q2�s�8��;�8%L�������T��YK"U�ۣU�/T<!Qʖ����Xa�o�a��n��_)f�´�H�t��F�3V=�A�Z�i�
^`�p�ij��  {U�{Pp���������S��w���R��um�e����0 m�lJ��\Ԫ���N,��%�*&Ԗ&������U^ۛ�;;�DD�9۴jy�}���wP���s9�i.u��kn̩�e��d�F��4����(ٍ�f�u!��2���i��8���m� J�l�ͣP��y>˻�n�T�ԖQ\��Yv��]b*��i-�t�Si`�vsd�q��nyi��1�q����6~��F���0�i.�9�t�v�A��z,+S��P���ypJ����#�����ADfR�-��Lq,]�w"���r�-L�����a,2�㥑j���6s-�8X�io��P���J�"�#u�%\��G<��\B�D��ϖ��sz��NS��i4�X����+K�$pNȷF}$���j�)�N�pB��I�����+0��gr/L�F5�i
�bT�<!KHOLo�}��{j�p`����Us*�ܒ8���c���on�aA{i��n��G�RiSTh�[c��9�����>#�CҎ�0J��xF�"���G��5΋J-����[��KTl��d���3V�w(�//|��l��;"�fh3�}���~6:ہ�-�u������W���=��HBȑp�ɛ�P\=���-��N��ݚ�ܹrX�P�:*x_���\ҋu�{{޷7�^�zn+҄��H�s"���T�y?�Q�����7���?]����f�#H�\5W=#�EzF�D�p<p����5�$�OI#(�NH�UUT�t]F�m�-�b�b�ݞ5��e��vܶ�0�n$�qAj	"�p+��\t�i��*�)�=ɕr�G|�|Yϧ=~����wi$.�ZP�1�8-Zi�
QJzC0�Us�)�-XG�9³|EꇅNe�%XE<#sܔt�R�(��J�!u�Jx]��w3�Rȧ��;ư�#�FR)��åGHӡ���R�
 <Y��X��Gs2!"�!�o#�t���*e0���M�Q��
#$i��y�ݹ��6a�D���0�9��$p[��Q9�Z./�6�e���-�L�.����۶3q����õ��n�̗�81�p�X�9�T�L��7O�5�^�t�x��mY�)dB3�Ӿ#Z�t[5M����H��[B�u�Yt�?m�v�}���쯯�U�l��K�1����x�*l�e��5�^�2�7H^���zGL92G��}ח��v��!Aj
?Y�4�6�=�j�x�▬��x_]��|.���v�$O$���l�dZ�<#�)zF��!L="E�ca@�!�vV�	VOH�g8���Ӳ\�K,�Gt���w:N��컟6����]�\��`���݁�ZM�C�3�9��v���"��*��a}���[�i�=�x*|/�>�ds1,
Ǉ0<�*���F��8e�h�VN���3O>#�V�\B�E�
��G�
��M0nX�\�]���^e"�)��K�4��y
a�fch����t}�n
��
A��q��j��w��۵%v�->�ְ�pANִ轷�I4�#u
���A΋O���7Gr�D�~��F��8m�P/k�ӂ�/��Ψ|/�f/�f,�_����PU�^�V��0�*�I�F@eio�@%��{n�޴ j��   P  �-�dGR���	U�\�,*�Sd )P  �Ҷz �w�Q�:�m�_'ww���s����r�^��.nl��ǀ8*� U	��B�p  *���3�
�r� c�P�  R�
�P
�v�v��sp�*�T �.���F�{��T�m�� +�6� ��6�Kd�m��    ;� m��U@�(6+{`  ^j�%GU@*��A�b6�Z�,Q2�BNȐTU�*��>�{��K���a�T���
�'��8{e����N��g�q�63�N�VvQ��SsP�1.��-��p�im�U����$u�lumǭ���m�vu��6��%�e�S"����]�y�t�3;co�ɧ�k���n�n.��L�.r�턛l-��\�1I��1C��k�=��lD8��pZ�*;s`{2�=��k]k�OY]ͨ6c73��M<!jl�1�<�ֵ���-fwNx�	9hLMn�a���`Hvv�nX�A�c���=�A�i�Z�8�m�"W�R���nLv�nw=�v�u��gb�r1ɱ��g����l*p�;�ٺ�]�2�ۏ��F�g.�`n$en��Uɛt읖�Cú��:��\ڭ�58ۖ��W��rbw	��7>�T+���M����z!����̊��7Ba��c'=/�������#d�;4<Xժ�u�s��v�d�A��f���A�7���p�L�l������Mn�3��`������\s�<&��\V�{p��9U��&��]<����jݱK��m�vݛ�-c(q�s�a�yk��n�l��m����mv �9�L:�%��WV�Y�n�m��s�N�F���ufIN����®�΍�jJ��ILswL<��Y�n79z��F�WZ�-b�������c�br��{!:eFx�A
v�ي�kh�6m8=���ދV����Xಸ���ƕG4c�\`ةec;zt�-���CYX`r��\��j� /ln�OqWGm�S�U�e�w*�B��niSu�l*�l �KJ:�2(&cZ܍T�����`mI���0�[��O�\퓌���vݭӭ����;М mW"vy�y��w>o��8ݸ1�1�H���Z�e�8wh���6�g�J��pj@�I�Ʒ[���qu۞&q�mZs��ٛ���Yy)�X��<�����g�\L�������5��!��m���g�n�6��.��NM{;8y��{i�V3�6�SÙ�c#�,���߿���͹Y6��RT�|G��0��1��lbI �ǀD��D�7fW�-XE=#sܘo�ެ����і���#J�l+���D��s$*�Un��D�t��|G��t�҈�a۵5�"�.���"��2%ް�8XC��61���Ⲍ��-@͔o��XF�r��Z�<#՚�>#�[Q�s2�)BZ�i�{Z�����k��V�Z��zC��r�3�9՞�CB�#��������ժ�U��"�Cg1��-���]�6�e;���a�÷lVr��;Mk�5P�s�9�Y��^Ϯ�T�<!Z)OHf�t�8D���Y~���'�G���+;F��ŵa�i�rbf�+ڳ�Rȕt��N�5�#H�\5	W<�q+W0��7:.-����ku�rP���|m�k���nl�s���3g�]�5VXŹ1*���v�ۛj��D��jf�u�T���"U�^���j�3e���o12FQc�/=:eҰZ��zC�4ʹK6�"|��B�E��g%jՆ{go���,]���.�l�[+l4�s;�ez���q�.��u����k[vԑ�5+�x,"��l�ޞ����tyg/H�}A��V��C�Z�񷻌�&�-?
��;$�2G+n�9n����c�r�8�����[j��8F���V�{�2�QzC4�Ter�e����R2����BՄN��E⧧O���Մ/�]#4�%\��P�r�)dZ�v�"�"�f4�<�v�;����J�i�P��^���*��׵��\�T�{^����d~,� ��Z8
m��!DC�)�̛��>�:D��f��ڇ8��6�oo����鮷w��j�9qt�ʁJ;Q�����]�H7�m�nޫ��:W��U�ks��R���EM�~.�ni�BՄN]I�6�xt�аZ��zC�T���Mֽ�[�rZ���ZyQ#�"�E��q�6�;����Z�i�P��^���j���#{���l�v�[��b�9��>=��j��pZ~��.v�{f�3vݛ6�x����l6CD���)�����KJ/$���+�U���͞���W���r|����8�8Nfc,ٲ{��W��ٶ�5�w�e��{��nH��/̔qffc��L����\;\[�e�[������d�u0�l�l �n
jh|��soyϺR'g���q����mʮ��G{�nۥ�U4&�H5���6�6s�]�Z�x����H�oZ��]�
%۽^F�[D��ax�2�
ח��M8m��k��^�Zmn�s�-��폘Y�<��q��m^m��D�����Qm���Xr�^��&Uv�z��m���,cletR:\�^m��B���o�Hf��e���mZ~�Y��hֽ�SD#�b��m�p� �x�Tp�%yS���w\�/UW@UZB$UVBj�m�R�k��A���
�VC�T�=��T�r��iorm�u:�ҽ�]S�um5EKe!k�nb͠�Mlf�VF�s쒕=[�;s�m�W�K�m���h�ĆN�9p:�֎j��;U�݌�*{��|.�Nٰ��C�g�&�:F��G�6�D�s��͹2՝����=�GlyZ��-��������Ļ��yMt�%���3	qlVP5��X�G*˶Y�äL���ɿ^�{���~�[��n��<���ˇi���E�B5�p���q"0�
�e�:)Fj픱�p����C�F4@��B'���!�P���s0��XH�Oj""�P�yFl"�r�^�-�#\<wM�DsU���ŧ�C����I�^2q��ZRglw떩1X�6���OI��n1���](8f���� �v��y���}:�{�Hz�;"cN��_@D���& H��������pӨ	jUp��sn�/Zf3��v����s�g�5!�cN���dq����RKU��8/�צ��^�w�o8��"�q�vD:��æ��������{z�mR��6͡1P�3�"�^���$XG��S��J�k�a���h��D�L�at������*�YYk`���o9�Hw��
Ď�Bx�I)�yܪ���"O �
'���و-ھFو��v@���]�i�l=���iD�)�W�xbDɘ}36�p��b�Rw�K����l�U�ﾨ�%��)��6��h��q�W��9���D��>V�,�u#&a=+��I:Q�������H��%Y�d�*eVM��'�l�����K���e��H�ՠZ,�����&���Ʃ?D���l<��d9��k`���&�~���bGf!�����2!����W��?jE�B��a/	i3PX�Tnĉ��6�敦���K��|��H����:I؎�R�����V�J�L���;�i���Z:2�l���p֖�R5re�Y��R!֫�1:F�J��G`�G`�I)��\����ٻ�gԊ{�e�[[N��vd7�t���tR8F�؍Ďfw���l�M��GHt�)�	���C�R)��6D;�����~�SΨj�op�/	J�U�
xk`��0F�L0��D=FN�ܔ9��^ݛ�T{1q�N-��8lKR&z��m|�H����\TR�4��'R6��iZ�H�Qɗ�f���}��A���ՙ�b��K�xQ��uf�3��^H��̫I�R>�a{nn�-H�Q�[cq#^k���`鵙��.f��.ټ�#ĉԏ}ȷLAq(��D�J&$d�1��F�HԍH�y����z�������Љ2;c$-�Kޚ�kg~�v���-H�x����#ǘj�qQJd���4z%�bR�O�6dR�&\��"nJ�p8���G������o�����͇;ǫw��MH���o)чjZ�$�+L]F�C=CS�RY	�i3�w&��a�n�ԇ��pE���1��D➘���*G�0�WR1�e:F���lLC���4�ń|�:&�i�[D���("ڑ8��VF"���\G���BF}E����)�"�W���;��ņٚ-�@�^}c~�_��#�ZD�DS��BS�<�=!��f��;g�����Pv��CCf�����xF��Y�^�2.�f��il��"�&ٞ�$�e�DE���#�7
h�6Dz��qE�s�"�B�u�q�{�PqƛhƢ�H�T5P1��8w6�]�Z���� �"l@l�mN-�c��U@�*�x:;��:�|1�|�gt��E���l�A�͹���L�c�j�Y��&��wY�l½����.۷��=��5<�9�,��ٕu9ܝ]�m�� ���ӒnS��S�Gg���z�'l�����UYed.1��|�r�<��M]>-�G�#cg�SI��h]l��5u+�3��խ,2|�n��[5�Q����3��n��W,��F��VD2�<b�߽���t���I�E�Gۼ��}�%�	Y:/��F2/ct�
'GG���\�Ee?�q��Qy�ӤY�^�22�`��i�i4a!�q0�����0�ݒB,�l�w:���Бg�����Uv����|.�8�"�*0��ծ��#�x�4ό���,%��TG-�.�ܻ�w�]6l����k���O�k��Q/����1�v5Z��f�46�[�6uɰ������Id�u���3���!�i�Tb$��2��">h������Glr!f��d@�y�,���I�:����t�p���^d><{�x�'f���G����a�)�$��Fۊ6с�Z}�oI=ƈ�D}�_��W}�M0����6D+/"M�@�	lI�ЁY�4�8|0(�����؜"�f��Z�7BQ��)䕤VwBE�}E�k�����g۹(l ����s��� ��~���R�MST�UT����Q�#�<�Y^�=\�YGc�]�βt�
Ε�ΟJ�k� ?6q��{A�l͆��5#�.���h��$�ԍr梹���[����Q�[A5gz1�:2�$�H�O=&�.%�� �gZi���>l��R|�rɼ"S��_H~�y��w�� ~l��������_�ffbIHo�+��$�F ����R�$�D�}(���u���pB�7�ސ�|�w\��$�ԋAOJs7bD�%z�:jGP]KR:��_H�OR27KY���%e%+�X.y�6���͇�#sY�D�II���� �-H�H�0��G߾F����,��-,x2�q-IGJ����%��Fx�7��&r!XŘ��ڻMR�X�ZR3�~m�n��O�'�u.�u�Z��$�ĎIwޥ�O~��p��1���u����&�P| ����+t�V��%L�k4�OR'J���$��>���ԏ]K�[�ζ�bFKi�s�9�̀lۯy�7[ �wd�����o�>8����s��}o��=�\�uV�KKp���I=H�u(7|�$�"dך��#�R�G}U��H�N�rK�F�-H�}����v.���\}�������% ����>���o��,�� ͝iｬ|� �a�yK�SL�<�d�C.�ڰe\QOn,�{A瞅�b�=���F�+L�f�c۫�f��H��jD��N�ĉ$�#�]8�ĸ�[� 6~i��>8���w��]��P�r��ސ�>m��Q$�H�g��R$�H���P����7��}�6��� 8��q��B'�3)��̳���m����w}�����U(L�q"I=�f�&��$��ϛ�m��^�w�����
�"D�&+��jG�.�ĉ��.����m��s���}���Ϛ~��l|m�+�M��\2�-�� >����5���� ������=u(7bD�&My�i�G�.�Ԏ�W��z�.R�� <���UAl��ƭ��O�w8l��NyA�]�jT�� `z�u��r��
�/Y�L�����.�mf�[k�+[v$�5�l�ˍ9�ț�
�Q��/�k�Nd9��ے+�h����s�"yn����ꃦ�{�����=�.v�>�u��z���u$�XӸ={b֪��3��v�}C�\����Ԟ΋��X�<:5� �U	rw�����m�c��؎�0��<�9�==P
��a�����"���/�����KR$�$��"�5�j�&I8�-#�D}�� �Q"I
�c�L�2()�EV����d�-ڑ�F�O��KMH�云��)��MH�#���#bZ��G�o�[z����:��l�`��}�SN#ĉԏe�<� �(�ԉLH�0G�W��y�͞l=8��Mv8�p�c�P��o�z��w�~~�@����z]���r��4ϗ�~��<�Lr�U\�C���N�>?wҒ����=/5�?x饻~c�_l;��e�Hݝ�ʶ�d�LA[�ú!��<c�T�M[p�xsv{;;��=nm0�$ZnWt�1�����)����ޝ�O�"���C���8��г-�N.x������^=,d��D=#<��>#��x��?a��}�mT��-�Xs�Ap�k�.C��e�4i��z\)���s*��%%�)9�@�Ze+�H���"���+�̸�dw}�&<u�E��B/A3����x��ʸv�</-YsD8a�>��x��t~�����ت��H��dݥ(z���M�gj���],H�/��"������i�3��8���o,��a��R%1�p�~r���t�WBp����o/1���m�;H��u�Kᇄ+9Y�t�8^Z�i�?��o4]<t��]�-����6Em�����x��4��;M�����a�tݥh��xBvT�l�d���X�æ��6��xD:^z!|x}3�"������:]�#��ٰM��}y|�������#L<!���ᇤ'fQ��[_�l���Z����Xl�� ;kl�f��@�]�1=���[J��w&��F[jF�l$�j$[Q0�GM��҇<@��iL�D�!�uS��><>�s[nIA�7l�`ܧ3�<pW��w�H9�k{K"/=�+�c�Λd�R��"�4t��e�)�:}\�m#��xa�t]��i���i���~7U���*hP�#��xE��q�W@���|����@�h�i��ۤ�6�)�U�i�o��L��Ƽzte�7�p��=�����NzJ�ӤZ�c�Ѡi�������8�T�W@!LV����[��q�B���+�2ޭ��7^q�s�M��q-�E���H�^�E�M ��x|G:���:@����#Z�釉�w�p��.��k#�
6��RK+9�]'�o�"����i�g�r���@��|.u�{��G"�"�d�r8ʹ����[�9�ǧr\�~�:E�����NzJ�ӤZ�v]<L���X�,P&Sp�鲷�'r�����q��;�e	�,���3�Ǧ�|�1��
���/8L�~�zj|��.���i���.���OrZ4J�i��ˡx���(��UUb�UI[MR�ɺ���&��w*��{��eUP
������@m���b����]뷮j�-y{"�m�x��\��e0]9�1�z��AZke�Ȼm�n�Fn-͠���Rl��!��5����]c��4����<��l��t�6-tգ:ͣ>��t�c���5��n�;X˾C�ËB�SͲ��DG/��p[�]gg;6�|l��a�놠4Gn�rYef�������s��,aL�C��h��M�:zn`3n6{<-�^2������j7��@���j��G5x��z+ߩ�N�켨�|&�ޑ�+%N)��ӂ�����%���Ÿ;�� ���M�#1oa)��8����~FI�NJ��8E>���4�2����Ke��ٸm�3l)*���Y�0�n^Z�TK箲m���Zfo�m�EnV�j3gh����m6��4䒼�t�W��4|xW���i���͇O��T�F��~�۴٫�h
�N���$.Mn.۪۝�вu�!۝\�-m!@V��A4q�i�f;N�8|xa��;�8a�ڭ9mp�!���7��v["
��U���p���]�ŧOW���Ҝ���x|�[H���5+���$�M���pç�/W��/�U\�W�U�DfE�uC��͖�H�����vˏx�m�T|v��V��(~��p�8�Hf�l�S�۾�{%wd���(�K9n��\n�q��V�Э�Aͭ��H����zz6=���\k�z^��7m�n�
����i��7}�saV9�e�����ʫ��,5{��TiI��,��K1droG�Q]�|y�f��jr��;h�s5�h%�I$^�Q��-����
���IM�*.�|�#	H�4�X1Za�eK;�p]~ᗂ;r�۩w{��L�m�1�m�/"�����}����޸�Jy��ݬ�̯�wͺP�U��RZV�Q1�Q�n��y9�vy����%�hvA�<�w�kݶfI(��� Bc�ǩ�����c��[��z��.��&���Os��oU UA�Kg�1�33
Lm<?n��mGi��t�-�Z��J�k[�,���ڎغ@�g��XE)%��Lv[�3u��^{Wg��GA��\@;\�W>��E���4ѷ1��Iq��L���Җ��7��p���+9�����?z-��o1MO��kf�JR�!�Ed��u���&7(p���?[p�
zeڸw�k�]+}�מv����O�ֱP�jdV�	V�J�F����Rӷ��.�oS�C]���m�=c�I+��7.9-7��K�����L���oe>,��H��@>�έ�����˦�-`[����b4KN���uw˧!Wjϩ�O�$��.:z��o+��{l�$��Q�@Q��앉���p��5?Ch[H���f�Qf�:�'�_DhF�-�co~��~�r��ˤ����W���t|t�bDڄ!}(��3$1!�E\h��n�%= i�sE�sOx�.x��'�����D��\Y�f{}��_�`������a!�6\s� m�m�V�,��w;rf�ପ��  U  T*�@6�뭎��@5�H[&�6��(��< < m݅S���56��R�^�͍R�޹���2�ib8��\am�8@xn�c ��< -�P ��{.��N�[ ���� �  �yT-F�U�V�	IUeY	����ʀ
�t�1��Ъ *�@   �jV�v�    :� 
�͵ ��*�� � wj������x��k��wu��@T �j�8e�$]�5&��K ����5�W��LGyw#I���u�n}s��׀/�9ײ�A�)"ڤ$�A��U
�JJ,=^�]��2���ma��4���eډ�8k�l-����5_.����M���(ֶӷl�h��n�b��rm�$��qÌG���lat�lkvJN��R�b�=��xg�W��.r"��狭t�/*���5j�%��v�m�\f��6㘠H`�\���w��<�ơۃ�"��B�ض*��V�A5b�g��"o[V���^d������$�;f�s�-C������Ǖx:l���j�љm��Mt�o;f��7Y(5k�/���×��\���e�8�̹��e���6��;5��f�5����E�s����vH^0F4�H�t<���܊q�����]���e�!�ٮūh}��m�
4�q<s��Y#���u�f�kmFu@�MN�زt��k=��K���۫&�'$ў� �M�1ط�v�|�#��3X*�OkN�1���ڭ�I�gB<j�6#��ʙ0Rv4kvN#LidklD�m\'OX����<AGh�kg8����WmŞcpv�k��9�I�펶zB�-���4ZuΡ�/���4� �iw\�S�5�1 �b�Yr�-��m�Ym6u={k��xp�mB�drh���`Ζz�+\�l�\�H�
�;���mO%84j�Sp��N%b�n8�4�5X��u�ƍ�r�3e�k��������@^������7Vz��̭�m���f�%B� �QEW�� 6��Afm(+�8�T66]:���N��:�;�[r�Q�Ĝ�9PP�]�:H5�9ɨ�ܵm�ob��6�K4hԠ�F�Y���,��c�;<S�W9����;^� �H��,�-�(��-�ld�������Zb���.�%�3Ӥ�x�n]��Yg'gv�j	��U�Uml�6�pb�sڞ�g=fƸ��'�v��8�vM+�xV2�`ŉg)����w�?h|t�%b�qP����-�xpxM���ʊ����8}��Oo�g�x�')�H8-�:~��c��={z�vuŋ��6μ��>�ww�W>��I	�yDO3���P}���x�{��#u�I*��K+9��@:c;?H��ۼh|t��Ǣ�T��G���/_����T)P��l�#�2��)���x����.��r���4���o�H9%�?J������#1�j��X)X�Y���`�[���;���s�	�I�;�%��-�: Ʒa.�:�c@G�J�$X� ��[�����Bz@�Gv��7>�'�6ِG#!�8�n��B�ʏ�����m|}բM��[�yk�Ė*S��7�4������T��)�o0o٫�]7���Y��3h{b���oK���m��-�y�m?Z����4|Y^�]�� ��WƏ��m�S��;��:dQH�q�t�s�㦛V칤4�:�5Nx��c���f�3@�ӧ��0�m�ݼ�(����27��I�(����:k4=��Lm���܄�P�%��N-���g(~4��NH)�@���M�ߵ�����v����;+��L��1�����[p�OҪ^9F��O
�����h��l��3�wM�m�B��K��ZS뫅���tz?n�4���y���4@��+�o*-�f�L�8�1�\
�w���ݫ��~4���P�~{T�٫��e�M8�e+�5k�P�����L_n��>�7h߇N�}U��0��W3Ie.�L�T�$��
�L1/h���I�^!�xv�z놗��a�8�N+t�b�W�\Y��x|����8G?���L����9���堺�O'3@�*�2�äEk��	��.W;����]=4�$�+%*����x^�����r�k@�/�K{WO�!����ʽ�o��K�0� ����mԉ��UKH���|@T�M��}�,�<���b���5L4&30�Ȋ4�n8��Y��g@3��\W���k�^ =�"Ƨ��9��K�wSEL��u����]��s7]R\Q�k��<p�tzi�H:U��c��Sm#�?g��G5H�WW4F��Y�U����0����y�����EK1��B�W�V���SݤB3�ӈ��?gb�C�E
�T�É�%�1�ףt0D��B�W²���w�-�˿A���um^ U�$�n�h���x]�n��1p���i>��[���9=*�;�MGsX�V411�����m	�Ug{.S����>����HOMcm¨ <k2��FcHe�[�U�U� �  ���nj���P۵=�ݳ��yR��m���&9^��콘0������Y[��Ɏ�Ϣ�*]�nmv�9y��7�28�Ŷ�odΕX3�j@y��U���	��"D��y�2;+�Ŋ�;(�W�bۭof�����r�����ׇk��<c�(��]����٬M�*j�wBr����MUR����rs]��c!	�śʯUNw
i�S<R�ǘ���l��ܓ�[];$��+.��l����%r�m�ÏM�9��o{�˓�{�FW����k��M׏'�ײDBˍK��W���Zd��*��ՖZ4R �A��/�k�p�ys���� �0�M��gz,�:�T��Y��ȍ"[+9��/���n�jK��Y�%�E���y��y�vM��t(f���w%�E�R8�`�Y�ve�]smɝ���|+�g�vi�jͼ"����.�m�7��+���Z�mv�����2Z-�a�-o�����A`8�����j�u�]�,����U�V*�rR9C�Zh��f<%�d鹣-�O�>������9��Q.nxKs>x�&�l?�l�s����6�-&92(��4{˅k�:%����k�{�f5FXAԉ�9>���]=�xa�^���S�0z��:�xӯy�����}���m�L.T�lڥb��VQ�q�]/�nM��I��4.۵��v}y5w5$��*�crVZM�H��W�H�x�����Y�M,{�ΑdJ���<FZ�/�G�҉�E �nU�3���vsE޿��~�9��ݯ����|��bq����q%�-��V64C��L�V1��:B�����H}Q�"���Y�P�`���i,B�C�80�x蟷�i���p�?#�];�s&�~�O���#�x]�[{Q]�i�`�s�t����i"�9�l#�P�(t�+�<~�����x\$�[oٵ��r��UUR����n�1��a7q�S;������h��T��,�Q���*��"�����F�zf�jc�3��۝[O#qt�S��}Ëq!2dd�\C�S��Z"0�
�ʎ��#�g�za�
�l��Q�ȵ��n&�I��7�E�����.a��^F�ȇ�޷�a�{e�w���-ް^&�+���ѻc��O]�_���w�E#=6�\J���Uq��+���� �AW�uOg�d�2SC�'���]�v����l�	�m�e�V�PC�vr��k;]"���S�:r�=��0AW���j�nE�I��&��v�ɸ�Y�O�Vk���rk���a%��5��q��o�nJ���S�9�t���κ�+�Z��^-#M'���|�ݳt�[��χ��7��d�Z�H��/�8<9�I���~�T�'&�������z��m�Վ��a�������/w��˛Y�nL���MKۖݜ�ŋogZU��]�u��+g.�V^�NP.���
�ڪw*���^�;v6�S� U� ��US (ꕚ��`䲹�kHA���V�\�Y,����a�mQ&�
W#��.o��=�v�x]rjt�z����R����	ێ�iɳ�ȱ����L���$�t]��:Ys;�p�7��l-��7j,�WN��{j�ഗW\��[���������y�UV	����\=9����i� 	)\9�6u���,tz������̼R���1K7�!JO>��{<nA�S=�ɪ�m�*�ead �ϼg��sWM0�Յl���(�����Ϩ�>z�ƞn����Ye�э�V�ȇ���̈́q�E�������%w���x\'�ȯƋ�>���p�9��h�^-7z=u{]3��oK��Eb���B4úB��"[��.�<��,��5�7Q�HN���~�aL�M,�Յm�PitÏ��l�Y���Mx�����Jm��]ntW��ϳ�nJ!(i8qO���3r�s�+^��8ۉ����0믇�ר�6s{�u�p�,ۚ7����%��~�3rP���'`�V��王㇧<��EO6𪘇�D��i�iSD�a:z|�s��%E��,�xP�{k�1x��S������)�饑���`�8|S��F�@UH+#r�x�����U}��黰u�]��Ӗ\���H��6Ғn+p�Y5'춹��5K����l|�|
ԓ1a<I�U��U"�4<�&�h����=�bx{nڣ�������u�� l��Eٱbߙ�!�d^?�x�"0�	ϟ����F�����X]h�i$�~P4���:!ag�ytH�~�1�\4�9�y���"[x���P�-$����2�M�ēm��!ᇤ\��l?B4ɻ~4i/�f%��_�No��M:?����L觾7�8��$������"�=�eOB4Û�=ZaK~�G�_�=���SOm�V�D�D5#�=8}��f�g��Ms��o.բ�S���wZ+g��U�X䀇��J̻��,�v�v��ΐ}1v�v�6h��d�M$�:�X�9;Uڌ�q[�zɩ{r۳���m�ě_%�ĳk�r�2�����?o�GW��O3&�t�+ZxI-<M��+1�v�e�Nf���oT�'&��7�t�˘�xCc�
A��s}rQw'_�����9A�n\�G���։1�}�$6V;�t�R���WU�|�|$��Z�Z��C�N�"mFJn3��eM���w`�2h��j��g�����Ҥ�;z%�y�E	�Q�6'n5�O^ػ�-�n�];v�����I$`�/(��xS����|���ҙ�K�T���+S���Y�`��?�y�&��^8m�����Y�M��c�����{"�3���x��z��+7R�0�Q��>.}�uR�S=���-��(2�8s���{h�o/��*7g=m�5����w�����:[��!��UUTU/ � KW!7j�w8M�9�6�J�PgwWt�P�c��� Ul��NjT�(�511�v�2�`8���+l�ٝ�Fv�\����l��{Gojw3�1d���s�Ξ9v���icv
'k������q!t�]='"���X�s�V�Asة�	�s��s�LC���r��#r%�u�Ѐq��q�h��-�`�PV�Ju�mc�Tv�u����D�g/c�һ��BE��.�0�<K-��kd�ɗ0Nȷ�[\�n)S�p��u:i�oU�%6��rD�t�QxẮ��浸��	�Hy"��Ⱦ�x��ݧ�gT�#���Z+(�"�^>��D�:��7e.a�۱*N�ȇ������s�l'��I$Q6�����xa�-�[Ⱦ�p�����,�ݜWE#L=6𪘕c_p��=���i܂4�5_<Eb{��SЍ4{{H~!ő
U��B�:Br׋y���n����B��:檕v����ݬE/n�6�oXfi\����0W�/n���f"^b�	+�#�<O�Û[X��&��K7�}�*5�y
%��e,KIL,O15��\f���r�s���s�j��+')<E�q�Cl��g�d���R������dx����~#bȂ�Cua�H�E���8�m��.$�r5W��F����q�w'��\x�>,�6M,���=�8i�s���ݱ�"�K+U7aY̢������#��!T���C�+�kyЎώ������Y��>-���6mo *延�O�w�z��|a3�Y��훴�z�&�%�2���l��q��E���w�`bՍ}�.����Y��%?�:d��|o�N��Z|_���D8a�Ks�/�*��a�$YՓx1���Orr-'�������M�,�?�ci��d�ܸw�"[x�T;��/tn<��䷕}H�tCM��l��-e6�q��rx���)��)�T�,Y��tޗM2�ϟ��!;�^8vo��+%��-M7�P}��`��;�7���y=��]���o����;��"�4�$����2�Z�sD�8�O<�Wg��]R��ݴlͨ�q�#^^~���3u]9�w��E){{�4�{Օ	�����ޡ��PLؒ��6K��'l����?W�$Y�ٽ˴�i�o8ŋ5v����I������ltV�O\��-�t��mCuV���E:!�9�zr���H�Q�]���uM2�3I6�I��<em#��fn]�:�{e;H��c'eã�)n�mC�YP�ӿ��p]�.ba�r_l���ⷕ
GWs�=�ƛ5K��4���_k�k��7v�h7r�-��$Um��^ۗ駕t��gJp���x֨��ն�������R�.֊����'?�����3�L��YP՘h�8G5����ִ_���c����QI2ŏF��ά��^�8iWM�|��p���m"��c�2����%��@����}�^nJ/j�sm�����e^����˻�g�h1P�	�"�j��ٚ�n��d��i�սѮ�_A���3���w[�T�λg^{���<T�eѭ	u{vҖ�8i͹������h�E�wʽ\J�6�%�[P U[+n⢩�\v�j�^�IT�l�U7v�E��SlVLÊ�-����Sn֍�DZ���Z��U�A���25kpE]��)��jbSp�(l���۫���;n����l�mO�G��ֱ�7W�Չ �n��f�3H�RW`:G�z�v���	!j�{:��y籕	a��mXx���<�gSh[-��4
�Ym��kv��e��1���Y
]�0�Z�nۛ��g;�q�!��t�nI�
�J��,DR��D4�4�t�=�mC�YW�w|V�xG8�e�ý��������|>����Ҧn��Ѓ15��4�踘�=P�u8D�oVzw	N"\SmCZʼh���6�+7�֘ѧE8G5�ʎ�4�5r�Z���{oGi4�3r�ߏ��	���`�*Х�S�9�흨w���*;"��]��ux���O�}���������B%,Lco1f`њ��8�t�6���n�ŋ5C���p��Vz.��:D<.�7�k��V�V�)�4�Ҹm�4t��i+HBV#�{�٫�ͩsp:�{���HKSn�,��\��eZ���
���+9����⦮]P�>���4m#��]�ת�t�gf�;/'z?���9�m"T=�82�����fݵ�e^*;�S�7�JG&"�$Z��4M�,���~�n �qyq��E�i����8ċ5x�u�$A�=�E�ÃqH��!��p�o���]��;��?�в̬�*��ۣqygU|������ f�k���;g���E�:�zF�mH��7�י����}��'�M�������0��;�Rc��g˓��p�K����8v{^.s�2�����qk��m3��Ӽy�{��W_[ލ{��mçwu6w]m��8F��R8�<nG�{��o?!;ょ��E͕�ux��U�#���gyW#�t��~8�B8�x�kBE�YN����y]��gT=#x�;H��7�e'idC҃��T0�Y��&N����;�*�Q���|C�-GyWM#�布�$Y�٪Q��4��G���+ʓ��RTH�8�\���5�8i�yd��S�H���Eö��YW��{7N���v߻��b��6bʵ+>͙`]��9.����v�=�v��]�-�If�f&LE6čWNȶ�t��՚�0̗O�r��ꧤo�i�j���^{�#��Z̶V(s����6mj�ʼc��S�O:��ˇyW#�布��Vu[��I6%�H���AcH�OM��1�Vj��-���M�s�'E�]:E</�q�qe^9:#s�����G\\��i?u��2��U�H�Syv�j����Q�_W���}|so'�Hdp����������t�zfͣmC�YW��疊xiޡ�V}_��a�6�Q��f9���
�ǁ���Y�����:4��=�vy��9혷i�夵�!Yr�ihm�9��N�gSg�Q��4���N1j�T���i��~s��t���s�I���U���3������b�tS���͆��������:еgSc����)�b��(Á�L5���Z�����r���w�ˇi�)�oڇx�����ŧM9��Ͻ�ER*U`�CyWM#��s��WZo�ZF�0��g8ī5S�����9�Ǥ4������@|ӂӥ���7Z�YW��;R)f����Y�U�H�Syv�hZ���~ |>�}�{�J���[��v�q^�Vªu�a��ޤ��ni\nTe�@      U U�]�̩�e.d�ʫ]@c��T1� k��*����^�c;v*[&�M	U���egG���퓩�J��H��x8 v�`JҨ UY���̀  �@    *�@�UT���Y�wj���Y�*�	T�iV�%eZ�J�` 
�Q� @���������   U�  UP 
ۙP�@ � *��T��j6�m�i��2�H[DLu�Q�Q�r��T@J�8r#Sƣ*�v"m%��e���s�o]��� T�>�fۢdp�Z��^�a-���u��K�����̀���0;>$Ԃ�E�@�z#�;l���uI0r���#K]u3�آ�vt�N8��n��yvZ㗩P2�7-g��rx�C�"����[k����i��e�Ex�:)������z�s�uЏu���g:{:�B|R�S�Nڐ6�t��.��3֎����F1s:�a9�We�d�nv�;�l�l���q�֟\n�q��]�>�a��=7��7���<���6+�b�ա��̑�Ռ󲨑��۝ь�V��t21�1P�b�F0���n�َ�=z�t���[Q�ĵ���5@�nш��b��i6(��ɒ6��[�1�L�Wmvp���I��whڎ�����h�^�5z��#r��R��k�-��aN����^:\[�j�N�܈S��e�V5ִ6A�jxN9/nI���]��S��=e6�۸Kq��y�)��ck�}.�[��x6(;;�vsm�ꬶ�,ʋ&ɠ�f�|m�a�Yp�s�75�u����c=�ը��9�s�5��Ý�u��t��$��xK�v{�G��im�!�8r�pp�p�#q��r+݋A��v2��Vnib�!�]3(n��h���\��J��]�X�QE��29y�w�I>�����el������s�Sq�5h�h��J���"ڸ  {8z
�T��N���g����ڪ�TGb�eUP��]նw��o �p�qU������j�oa+�e瓕�*��tݝ٭�3�N���is]���t�$�ڙ����V�&J�FV��趕у���g��۶�%�D����m\>W��\ۍ����$�5Fgxĥz��5�8�Ws��m+��W��q$Ru��,흆kb�YV�a�c���x�	��D瓦P�x��6��\b�y�fО%�\[_��>:fm��VuS�7�Q���>^R�m:E=2�nm�wUk�6M$y��1,D�ʤ�����?5����w_�E�u���~B՝O��m#=3h���=?��v����Dj�폚t�w���D�N�O��!��j�x�c�Ӣ�4�vege\4���%^&�$<h��Xoi�-\��WBp�i�윣E�z���(�p�9՞奕���z}���Ԣ�X������O���Oゞt�Wˇm]4�����E��c{��t{��6��5#�%U��B.���vv������N4��C��H���*�hA�Íy;����9��8i�s���:t�x}��6�ƭ^<�k֢�~�w��)P�b��S���쫆����:E��O�M:}���oU=#s���#z�䤌X�fbL���%���zfͣi�*���O<#�/Nںi/%],ϯ>?����	 s]2��v�i���ڴSơ�
��p�H᳗Nl�.�M�{͍�Xqcl.��d�z���?=����>�ztR�}}��m�v��q.jec�ʀ�u��he�V�*�\K�`_\�ͷ8��g�y�I��X�_J���s�^��;8wW�H���v��pڼcw�h����;j�x��/R���X����x�V���4��˜:)�zB�u8t�p�o��8/�NI�,xT@�X��C6�ǔ\X)f����EM#�M��t�w����SN��{��0^Km����x�Q��H�Tj�\4�z}���#�U�2���:g�$�b��W';����K�:Y�U���N�0Ӧ�+ŢU�*|B�]Ni��Ul2Y��m��q��N(�5m���α�a�����,J{:�c�
�f)����Þ?��ܾsNNꮓMW�*�vY��97�!����%"��;�-ꙵ[r����֊\�[��λ��|�y�%�6�PE5���{���dsݭl��#����[�[��)@��h0a!��,���ӓ����O������G����H��	&����ڶ�fjͪ���Z�Z�ݭ&�dD3!)n�UV��2;Yv{t��6�����q�*;����O] �3���8n�[%7~7���#�W�
��䈏I6!�HA��|yr=���D�V:G+����zaʸ��0��l���m?S�#��kR/�uk��~�<M���ˑ[�L�]?tټ�N�j�W���L,�o3D�x��t�a��U����cƚmc8V��<>nQ����^3.�视�#�oR�U������-\�^{G!�UQ��Թ�g���vu^׽T�v�a������~�Nz�g�X�����_?ޝ��d�*ҩ��U�'m�{��.��x.�*T6�*UW{���_��l�;�JJ�T�3�l{e��3` �3��k�8bT�=���(ۮ�K����:��֪76��L +�!�לHb2k����mk�����qp99�m��:��[����\;L�a�`��
g�;�mnk��y6�qnj9P��z�v܅��l�#�[-��@�5������E;�K*Y݀��uTd.�\A��ca����8��[�:㮥d��;0���R��ȴf���������M���u�
��oAS3�V�S�P�0�Ź-B�*���ts�u��~����l��]3.�臆�<��sߟ�8j�����[]L+b��!�*��7�a��E�OD;����g��ބ��:V[RÌ�B��3o"�%��v��,��Pͪ��O�7g.���R�j��L,�m��ō
�TjUd��8��n����=��b~ط����j��/��h����1
��5�z�VЫ+�OS�Kv]��݇"�2��d��7O���32��,*�1��{:�~eڈ�o�ڔ���7�afz��������K�y|nn�t���۴	m�UY�3���s���KŻ�.`����!���?t��]�Z�7���d��ƨHܣv�)���;�����%N��x.Q����NYx�|���l�D�7���W�����r�gWO̻Q��R��������ɭ�eo�>��E)�X)m9��<�j��;O�:r8+[<�1ix���������?���#e���Pٲ��q˴���S^ώ��L�1BRº�iUűmv��K���O8t�P��W��o�/��(�p�/��s�돴���q�XN�JH�m�]��Ln�h���}C������K�!��,�z����d<p�5=�h2·����h�2�񇽥���<�w�g4W�r8+[<��im�
�������q��-�ZJC#��a�����Q6ӧ���0�쒥�b��NZv�3�t�8�luZ@B�6��������ճ�i��cw��w�y�ѳ���*&�������[����DL��Õ	�zV.Y��0
:�mm�N�'��s�b�6ӎ��%�-�m���J�W��z���z-\j����L��˷����N�����!�(�M��sg��Ԟ��)F�qڪ.s�e?x�޺^!>W�	�!���`�Wj�|	��"�,�1Ѕ����~�ۺ�wLҜ��[<��F�f]�O/�y��vut��/(μE�c0��#i�!j�X&�߷�a�=w*OD��S��~4�!Ϋ���g4�8}5k�m���l�Q�k���t�A�R�=�2���8����r�:еu�)/�ae@|f\I��ӨV�VVT Lq��&͂SN}'GBA̷��_��q�sٻ�\i�q=(Z�������ӟ����|��-��zc�F�!�(׎K�z)�x��J�C/&�o��gWO�.T�C|���`��߰æz��/D��S��~:{�~w���v�\u��m��4�'�V�y�t��
p��C6*�T�����i����]�Cf��C��f$�,~�29Z�j�T���Ӵ�C�O�+Y��ONz^�Cx�^*�HEV
h7!����>6~3ެ�:�X}fJFC|���c<�~�C4���ʓ�*�v�Y�k������UUUw�5Ք*�;���\��O�6��lU*T 1���6m��_����b�*����W;�ԥ���P׎Ԁ��8�V1�D�fƶ��]�vs�ۧ>-k\T���Q��-��,u`��P�q�ˇ/W`�k��,���[����{#�&4i�	��)F��@T��2#�/Ht��f���H��ŧh"$�Z2%�����ۆ��	�w��kjG:vK�&�gi�Yg�['gGP�{��l/n�$�5������-e������Ǉ�C�W{�����x^z��چ�V�x�Ti˗z�T)�{��I*"-��I�w\a��ӹ���s�����:�Tޅ��!��EEBC�k3l�=S�d���������Ȟ7�_�����4Tӥ�彲Kb	"-��ec=�5O�\�.lC�Q���v�����؇x�]9����������T��&Y(s?Ƙf��u����г#�/D����.�}u�~C5;�m��ڈ�䎠���a|lz� �.}�:糭���V{tƱ`�dGkk�W��"Q�m�ϯ��o��N؆�V�f1|w�0�!�9Q���NW�>;�}�~{�{�d����"Ƥ�?����n���T���
��eC�NokIm<?i�YC;�x���:R��sBgh3���4�oo�I��ҿzt�<T�.ӭ	WZn���Ӧf�N�WZ��Q��3<�X�m�Pı���s��+Ӵ���fѶ��U��|V�xi�P��(;]4�7h̸���_���6�����;p��i��m*z%Z�>!r��i��rs����O��}�ݙ�1rl�l��sf���)�`�qpq9�<�N#�s{�M��`�u$S�vtS����O���{�;SOx�i�8��x��]�Z��o��|-4���kn�$�XZ������O���6�mC�O���ӤS��F����̓.h�M=!;jM��x�(�����gB#M��mw���?� ��ʞ�׫����T���K��pu�&�K
+�-���N�ǅ�6��C3��-�0B�:Bjs��GJ���p�V�~�	��_1��;H�O�m!\P���6���GM�s�a�!���ð���'�ed�ɶ���V���ݳ��xYӸ��/Cb#���e��z'X:�U�����9��Ə#_��Ň��O���m�½>�Ft݊�f�SP��O33>8H��cO����ͥ���x_��F�8TZs*�)B0�	�Sة�x�m;��[����A���gט�y;��6�h�⇄^i�p����Q���x�o7N�$m5��2Z��y�:��ʇ<p��:��#}���������<t�����qUh�@�>-63E/=![��i�^z�im<"�3�#�E��b�X�:C�Cߏv|nY�D6�*���W8'�l�i�
��pY�e���=�H��K���M�gWL#�^r�8D+U�W�S�W�4R���/�l8a(1��G[QE,-��N���n��¼YNG�駤zޤ��GK��C�8�YU��DEA&A@�e�W�<6sr���=!NT�i�p�[���t^:_]�W>��vN��u��GRhkP�:B��~�ү9v"��C�S�fѵ��P9���M2K����<򾜹V���8c�Y�{[y�g����}��J'$�9$�B��P E�ʕF�0P�J�����%V�*��`/T�w� � ߞ���,�T�����/Y�5c9�V�SaL>�`�]l�.L4�����\J��D-�Y��%�Z͹��;q�CJ�*X�j۵�3�q���xs�)9��S�	�\aټ8�6Z65pd���B&�۵���jS�Q�42@�YXF���hL7�r�ֆ֥��!��;iw[��K+F�U���f]�3��0]���\�u�R�I�q�)����-0RO�櫁����~SF{�zB�K��p���R�xD<>�WZ�Pr"J�d�S���ᶭ�4-!�HWU�T�:U�.ÄC��:hp�<p��6I�T-T��-$~8-�m>#��\,�xn���!�x}�EZ!ᇤX��� �ăư#��X��:a\dg�#ǆ`�O��6�m/D,����a7e�m�B�Im&�[O�K�����M9��X�:B�2���G
�.ÄC�i��Τ]Am��(э��]�+<�5X�8]�c�p���boZ�F��='/[�`8V��tܜ�D,ä]�h�t�8n�S����[Hf�q$�(�	[u�I_��?}�WJx\,�O�� ��F�tݪ�f�Y��{4�ڙ5�2��$�������?�".;q��3���_�R�:E�\�O����m��jt����:hp�a���4R�="�v��#�����Vϯ�g�ݗ3L@Ɔ�m��3�m+D<0�m�æ����|t����<tzsuX�Xd$�MR�[QE�mY�ѷ@F��,tRCv̩��6枳���-�ݘX댼i腘zBr��L#�z��[O�K�����M��E8!��k���u�o
; �e|���{y���5�6;Ӣ0���l,�8W���W'd����/7�t�#<+ӕ�xa���æ���!�i��gc,�m��D�7B��xٛF��C�����i�p�^V���!�����V���S����&򃪨�Ui��5�yy��G��{'������lb*Uj���X�`wn�=�1v2��k�9ޞ��Ϟ�(�g �ak�F#��V��<�mt�Þ�ɯ���wY��Щj2ۊ@�iDb�o�&d#��xfXp����a+��+�3��q���q�Ԑu�J3�O6oJ�Lg��ٯ�!���|@i�:fq��q�ͷa0`RHJ�4x���2�p�4ݳ����l;�����zk�p������[�e�/1�����)�t�:xT�f[��\S�%=���@i�$�T�m�qfg�`�r)i��n�v�X�뼸|G���a͜�v�tᲷ=>xYTf���o���|^Oߙ����*�S�!]V����{y��緶IU�*�d�������(��t�M�Æ�혝,�xn�Ŵ�a��
J�S��JnF�q��g������F>����Rs&�a��m�腘zC��AĂ8�m��a�p��T���YC>��t��4S��0�
��8a(]=�2�FG`� 췞 �p�M��S�fѢa��K�B4�f'Kg���K�J}K�SC0\����g|���p����^�����˝�3q<�Um��r�m�sإA�
����>ު���6wm�w^�i�@g;����i67.�����Fɭ;��w<�8_/�9�؅ֹ���H���$,��`.�Av���S�3'=9.�3���R�w..�9���kv�6"ve�5�Ӱ�Y<�VJHΥ��(�& *�#��;�t�MzPݵs�T��\���7[���c�(�xw�|<��n��gۑ���qJ�l�վ/f>~#<)۟�G���;/(�xa^O�B:t�I��a�d�I���2C(#�P��!m|���QΝ�V��<t�KƦ�S����D�$��n��-�S�!�t{�o��P��,ͣE:|t�b��!Vk��n�
�%\���w��a���N�F��oN����}�������X�-u0p�s�5��ݺ���Ǥ'�_��s;#ka�</�կ�<R��\PЂ����Z�L	��v�ش'�5m��9k�U�mE�9����]���W��Z>~�y�.�NÆ+��a�\>��:4B���?k�����QX܇</
�˅��xn�ͤa��{fU�Ǆp���u�N�MӢz�Uh��$��E�¥V���0��=,���K�x�+�g�xG��E�2'�m4��C0�sk�
Y��l8a*�,�m��������1�m�����d�}Q����v�m#<3�z<t�"�@�.�Y8��[h��ԅ6E-S�R���dغ9�fG$�kXć:��kW<��Ӆ�����o�.20B:t�OFF��e��Ϗ�:t�>zF�L�۰�RE*E �4~Ý���C2A�`��Ȯ�N�|.w��^�EɵF9\b�[
�v���۴h�C�2�C�{r�l�M����	��45��d�XY��zG�R�>#��Fx�<DN#��>:o��m��~ҍ���=-jR�$�ŋa��+��m:D,�6�6��3]9E(C�!]V���*x\U��I���	��[�����t�.�К�WZ�(�A�h �<{"�K�S�۴h�C�2�K���y�i������j���ӊ���1��m!����N�xa�
J�,�!y>�G�
��#aa�����2J(�\�U8�S��?sd�x_���a�!��J�m#L:nl�p�K<p[/9&��X��G��x*��.ږ��M��4S������lq �:�H`�vr�M8{�}��W�����G}�}�w߀ƶu�����B�j�ۆgoPs�6㉭�zU�J������9F��RBӞմ��Pz��򧝰�u�����^�����cF� H�kӧ,ä]bӰ�p�����M٢��F�t�6��H��ř�+0��M5��itQ��!��ô�a�^�)�=#��t�B�����=ǖ�2������7E�
tݪ�e�ș���vf�f��9XR������Sm���/	����h�xl����>�'��K�f,ŋhsh�9gum\(Ck�UR��v/Z���Ou��A�*�lR�    U  �j���mǡU8gV�
lU��	�wT�p
E�<���x
�{v�U]���r���#^T�;+t&�*�ޯ�<���*�w< <����� ' c@ *�}��^�@�Z�@ �`��Y@   B��@ mN���K/1���V���)ђ�p�[m�*���EP 6��ZU �E[Z�  �}[t� )P ;��ʬ�{  � ��Sl��FͤUe��	]v� =J[��oj� S���B�j�Q岷�jY�Wme@�Sc�W��nݳjEᇪc
P/E6�3�W. ��gT�Jp�������W4v_j��pFr�·f䱥�!Y�n�X�	�7;#S��Klc�H���pd���LZ˵��7"+�A�kR�V^��n�l90L[vAv]5\r�_}q����(�����F�w*O�v�5�)��'���l�m�:1�wm��䲤9d�-\�1���S�����g۶�f�c.��t�Sh��87=���V��X-�h�j��m����7@�GVV�m<qz�j�7
v�tš���4.әM]=�lq��9�;m[=n�<]r��t���9�lm�q�@���6���qH���*�������C���8��=�6�S������@��5�"���Yl�3�s��)ۗ��hŋ[Sm��[1]���uf�z�5�|c�<r�S��Adz^\q� ��{d;$iA � y.��/����u��(�mk��e��Fia�e	�-��J��[�
 m�Ja�8@ƣeջe��q[�-��n@�i�cQ�%���v�헭���v<������7`{˧�����M-��=�.���s��rm��3��*,��X��]b�tw�e$��՛\s�SN3����`x�+�"���:�	e�s�)�.Drsm�e�TIk2�0`��B�ܿ:�F;on����t�;�/�L�v��C�q��۳��
�ik����V� ܹ��� m��e3��*� m���R�@�Z��q[iP�ت!Jtd9�5U)��!��v���-����&������uꇶ��<C�7�v���h�O�Z��f��4�fz�7i�Y��4�=�:����P�ۭg&�E;��1��!e�]B��`%p��0����$vĽ�����8�-�!�FI:g۴�񺍞�-��Y�mmR�&�H�����R1�ym����9A�F�s;�Eql�v�G(�\�i��p����ӱ�j\�=�\���<��M���ٶ�(��V;Ni��G�)��:t�o�;�鮭�4RϏHSn?`�}4]d��W �VBWeG>8e2�^�i�M;v�,R�:B��;��l��^:o=�m�c�[m���t��h�<!�ip�iw�K"��;Hff�����r4��;_�x辞�����T�OG�
����0æ�4S�p��T{�b��W*䶍�(�B�l+�1���j�6�]����O�mt9
��$�;v�=����xa+���nI^�i�R��C��+�Ѱ�G
�L�n'���	�D$�6�G��ޓ����e:<t�#,������La#�Pu�dn�"v����h�������:/M���3�����{gF�Ƒs�W�,ܝ�{g�^�v����\�F��,��;����T�x���Qp��%�]�矬�;�����x�:���#�)�̅d��������o[z�5UV܅1K�Uq�Rݖ��Gn[��Ƿ:�^P!;�u���xwnz��if�4���Ј��V� ���m��4�!Ӄ������!�M}�J(qf2�6�X�i��24��AVm���t�-9��#"N_��m���X�ζN����k;��ҽm{�C�z��;�8Fݕ�?i
SAĖ\#1�����Z0��i���#�Kf��CO���-#���ϺGL�-�`m�Ec	c|y�<E�R��a=��J{�Dn��9��p��7����d��T�R��9jnq<��.{]�Ӷ1�;=Jgb����6z��n�q��2�*�*�&����6W�x�+�׽<h픽�#��Y����m��<o�4�Y11��_{<`c�˫}W���۝��w]��� �\p
�8oS^�⛘35,�xK:�%��0������$��V~���Y�:��R����	l&ԈD҄�$i�N�d���š^�>�Bh�|$�ِ�� -*�mV�W���nl�W5z��+f�մ�6:�z؀Y�c��|B83�x��p�!�ùE�iG����Zp]���X���St����t�͡m<"����vq�|
�;��i�۝�Q$�C&^co���Wtki�ut;[O���k�i�B�]�D�����(��Λmi�x��F���ܣ�7��V���l(�~n$�E0�s;�'����� ��{�M��̈́��?w��QWl�Jl���ʬKd���n�i��^Z��UT+(�T��J�p` ڠ�U�|�.�՜Ŵ�@qڛ��@�gb���݇�b�.�`�T�N��Ajlp!&�8��N��U�m���jI�Ӱۑ�=����';�^-vu�ш�4JK�;2�K|TX������+�v�˞w��Dsw!;ls�qa�bYފ;����e��P\�1��o]����@�@��L$=�^FW	���%��,hr�m�lno1h����DD(��)4��>���[��b�6��s=ո���v�ѥȴ���I�Ls�ٽ[���<[N���>��!ݻ]�#
�TL&Ў2Ae�r�z�=�[�E�$s��'߸D:^[^m�o=<��X
��9@�o�..:����u����#�M��Бt��\i4�:�:,]0��K�K�sO"�gi�ަ6���!��~�*�O���碞�C�R��H�ڎ���a��N*KJɻEv���6�(�kFN�=�b��,�r�@	������n7)����"�Yb�m!�xn�
�%\4��*�t�U�tQ��)Ҝ2�V[a�8�ceC�T�g(5h�=�x�gif�Ҧ������ǒ�ͤp������n��6���}4�W����*��U�����Ѳ�ު|v:|�S����m�Z�m<x�;N�GKʈ�P�t��W�3O�4\�*��J�Jt�U���T)<C+�Kl1���u���P�*zV�Pj�Ny�2�Z���#�M�������M�{���[*�7l l�m��7!�����0�tq'=�vI���s:@,����`�˖�;g������OH{TN�6�ާ�at���}�l�~���Ө7�U+�bt,�H2�g:iޡ�)t�R�Hg��Z�Vr+����i�.h�L="˽�������'��,ʇ
���H�M۵a�P�O�5,�x�N\�i�H�A�1�1�*��&I_<v�������4])e�Bb�F��'>�t��#�M�.�2�E��ʇM Ư�{{r�ۈ)�=;�->�)�Q���h��B���y^Y4�6;�N�Ѳ�����&�h�%�bw9��q��vRS$�S��,泯6���v�5��6k���nG��KY�S�Ycq�Ӭ��˩����WWG�����{O-�Jm��0�a0\i����oR���&g�;�<�n��H��_��T!�}��oei�\�� �]��4Tӧ�-�L=!N�fD8W�!;��f�Fʇ<6�ζ�,,���4w0���p��!�-y��H�SnU��O���#��6r�b�0����3?3�8�eH�eN1��W\ۡ.�)��E=���h�X�K�w>�L��i�,����1,\�p���N�Nv^-��|g�:!�z��-�xi7(\�J剖���iε��wۜ�CNɣ)��zB�\	æD8}�����C��q���H)du�N{Z�E�5/�!���R���GL�ˇi�!���j��.p�<l�?̪�Z�,�h��xEبt�*9��ӄC���;j4�*�3D<><��s�
m0pfu�Yo4Z*HnO��_=:{W4Xi��tC�p�Ϧ>�p��C#�;���9Ъ 6Q�z���k�>'<�w�nz���U����.��0w�;��eR�����c��U��>�t\��3r\hX��7
�g\�)�V�0,�ӨA��Z��']�`�\��/8�s���9w�pq�l)�m�e�n����n�6c�k&�!���W��Y�c�,s��f���ĺyb�H:�m��@fmvt����bv��'э�/h: ���f�@lT���\�6^ۄ�+���n�2h�K&�')�jC��v�[���yO�K��hl�w����zMX)�Ox�mV��Y�t��*�xеx�g�+�m(��dA�P9�=���~�ڴ��7|ht�j����"�o��k�^��8�&AJ�R���Ӧ�����[O#��g��Z�W��a����&�p��&�u��K�	,Ł�if�9�7o��xE:_��Fڇ:��yB�E8i�!����N�GK���h&��ki�B���[H�K��ūM=!鰺pʇz���۬���~�/ߜb���e��+���@�����Vຉ�7<���E�	]��]n+���=��#�kB����������N�Y<n�ɹʸ�C�J�܇r�n���COǹ��i���*V���TWD���*�U˷#�&8��C�G�ǽ��=���8��� �PB��9-1�9�E�t�Ff��l�&�c��3�v�5��e&��l��>��8o]vN|q��{|���=����2ڈ�rRD�!�����f�V����:#��_�����Ρ�8'�w	���+�X)X��i�dW)ɜ�nA���弡F��1�H�0+�Յ�Jm��wA��߫��?#�����gFG
���Бd�
�G"�Ab�!�����
�`�o4�i!ޭr�p�x}�͵�:wҏ-��;gjѧ�g�
���z��X�`�k�i�6ns8|/۷	�=P���|>+�߳����?o�����������-L�y��s�=�vTk�9�]��Z0��z�֍hH�[�Y���~{��8��Hh�p��3)t��U��t��;9��wT>;]>�#8�������K��M`��nqW�v���7g��m��m�;��	��^˺y͍f��lrRJ�߽���=o�-BEӖh����"X�7G���/}��}�����\����Q��*�V�D9�ڴQw�|y�`��v���k[O5yx�-�H0���,�G@��p�|�@Y�\,��w���q3������ϝ&����)4���|s�K����mDg�{˧9te<2Š���a���#�A�6dC|��x-�#e���!�(C;C��#�C=T�l?�����|;����m�fʙ�si���nS&�(8�sMι��iƞ}���Q�_n[��cx��y�{���v��!�<�D��=_N0桘���������$0��m����!�P�̧�����������t�����Q��E&�`�V�z�$��æD6+�|����"ꇧ�9(O�0����[�rC6�·�����wN}}A"��]U�2ͬ�p��{S��]��P�6��F$l�[pW�
:��7��C�8�����~�l< *o��ޓ���;����Um�1Wm�P����T�t򺸕O�6��0�*�gM�UK��Y��w6�OTATol����J�fz��EFͲ��ⵎ8�3�?�ro�~�]-�]IӃ<�s��͞�۩�.������bM�A3�� [��j�C�ˡ(۷O7,n��W�Rvr�n�kW��㹀�&�v$�N�stV͗�+dx5�y�x%���&��v�΁F5�A�V���]��
V"�6����Us��[nn��j���/�;�N-lU��6Gk���q�s�i��H��_j��%�p�"]�ipKP�������[E�"��U	U<��e�.�H;�l<hH�o^Ջ@���kD���[�f"�X���ř�2!�.^P�Os���]������r������m�[�h���������l:dCb�/��@��s��	!�u7�.{Z�����W�>F42�n-��,w*�s�H�own$���_�u��q6�m�\V���M��lb�p�l�`Ɠ��H]l�	.\em��A4Xk2�H�a��k��.��Os���C�P��]ߴÜB{{�E#3�R���w>����^�	J�ї�f�7D������ӤM]}������7� 3�����!�x���B��a��+;�%v�ϫg��s}���d��CmM�-���Z$\0���~8|G5^Z S���9����_�@6X�ר�1��*�d��=<F��Z}��f�%\4�ښI�R�33@)e��9@�[����.�nB1���I�����h����U+�1A��>|i�Ֆ���K>r��F�x��{��ZCJ'�����t�����QX���mm,�WLwzJߴ��,�:-Zi�)�_�|.�����f�?J���-�B񷅼I�gikǧܻN�xi��ʷǇ�8,�<a.��g��3փ̒�
��Z+KU��|4�l]N�p����o��~��󴍤f��x⡍)����I�`9uH7m|X~��mkidZ���ߙ�f�)�jc��_�~z��.̀�cJ�m��l]]6�x���2w��Q7�m�N.�ɌI�(�l�e�Z�Z�6�&��o����H�C���F�xi������?x�O��4:���jFX1)!~߰���V��T)��t�������M"cܝ���E�@�&�k>7u�*�!��힌̓�2O�&x{��$�2	Q)�@�ի��û�M]N�f�>��\���!)"G�8�I�:��H�x�otG��oFU˖�{�ix���rqڶu�J�������&���1שۇ�ո�;um�'��:�2��c��\s5l�-�������퓍L�{�)oV�)rN	�2Aܹ>��V�s������Uk{�W^�������T���uY_|y��;�)ů�ZD:p��UtJ����p�zF�o�\G`Ƃـ�G������������<4�-!�pӤ+�+;ç�t�{���[��޶�,"be#�����c��Vie��g�s����i�)�v�����9N�J�Jx��`v`Q�m:�ս��*|*�ta�l���Sb�A8*�^�@� �T�[vw�]Ƥ�J�+�J��ր˸�6��萲[A.�+�+ltg-f�%���F=�&J}������<��<�9v��^\����t�ŵ�G�-�^��{=of��E�0T�,�L�gP6�|u���۵��2������w2텸�9�rb� :<r����:J�SnJ�<�iB�����C����lu��f��VB�4k ��P�T�T�+�,t-��u�ÿ���f���8mi��V�&_���=3M�sD��|C��H�RÍ`e�a�"��z1�D,�[�7��d2����Y��C'-moH�t�.����?��,il<�$XT�����n�b�#�GO�|�J�)��`�m�̑�, Ԃ��0�>���h�!]���)r��xޡ⸳d9F�4����t���XJ�m�^/�p�'p�O�+'LB<t�ݬm�Q�T���W�>9���O�hT��ڕ�"�l�ȶ+[��q��!A���\v��nB��gSF�`:76A㮣�7�
G�n�-�������#����+P�d��fD:Vh�fA���O14�1�Z<=��m�t��̼:<x|{�+��څ#NV��T<s��;���+�-*n:��4P���N�q��=!���D8T|1��,������O��}�Ћ�E�cÜ�C���V��L�<T۝[Nqs������O�q1J�#Ò�\i|R,
�����s�zsN���FڇJ��;�[���:�ʺi��5����D��@`C:^���m��t��ջ�����~��.
�P%�s,�1.L��<�w�B��~9���zk�2�9��[�38��B�}a)�������eD��Ж��su�_���ˌ��Z�I[[ʸi��s�a�!"~Ww����N�|���@�-��i�C�K\t����Y��g<�Nӧ�9j�P�W�n�s8x�~����R2<�'%v��u���qipϤ����[��9�3}�L9��h��+��;'�n��˸vᏋ��N��4�cܣa|BD��������aU��l���M��r()u��Y:�`������Jɬ�a7�Ar�+*晧n�J��z�x����*՜�;N��z�h�PާV�}��i��\��G��;��v����9y"~O��/�O���f��=���i[��KD����6��&�BOƟ�=�~�w�W��t\[�^�>ݚ�?k�[��H�2�TKZ�y�H���OO���c�8��s���|y��.yo���}t*3/�>cgL��5�����fv���j�6!�缻_��i���⸸�d����UJ��Ujr�#���vb��sq�u���	��U��{Rٻ)ե�%�����P���\t��B�eނ��>��{ӹ
��a�6�3=�:�|۪���G	a9��0�����R,7Ga�m�S��a�ㅟy��uw���j��	BIy������Շ��{w�0�P������E�	�Z�%"�!�?���9�X|E��8g��\ݸ��?3�D�\:{�Ѷ�~c�����9�e�x��nzi�/���ka|BD���_��Y[���~�������������/���x�,K���,K1b��k1f%����1q�D�,ı��Y��13�9�fbY�LI,�Ř���sىbĖ$�����bć��=�<< ���������׼�� o�
�o����/��sŉ,I	%�bė�3K3K����sŉ,I}��>����bĖ$���������K$�%�.���Y��h�f%��ىbĖ$�����$�%��+ŋX���&��l�B	�������������:�{�xx��������#���g�A����ıbKQp��K�����sŉ,Id٘�� _����(+$�k ]c5���0
 ?��d��0j� �TIB����l" 4@ *����H� * �i�"�� ���tV� ��%}�     z          :                       `         ����p�!�1A�0�=7  ���[�t�c�����@���A� ��`���O�  � ��`    ��S��{��eq�ҭ�����Խ�:W��� �^ڶ��=z�4�-�+-��y�=5Y�  �       w�zjW�Δ=w�꧋����c��  ۭ,��}��W��ַ=���{|� �g�Ͼ�mM˫�9�u�Z� �UT�0��w�P�j��s5N�p ���s=^7����N.�V�          �y�޳{�w�j���z��}�@�� ݩ���^�x��*��h` ޭ[qn�g�{�x=���� �µ�o��W�;���!�+��Nڜ �ҽ+��W�q��k���U,          �z��^�,
�8X���  νj�ZUW�����U�-B�� #T�-�T.Z���CULCU�� ���-u��Uu8�ڞ�|�M ��Z�y�������[y��5������    �      ��qj�j�V���b����=� =��T��z���O-^{��Vw� y�5����yk�Un\�qn�Z��}��f�>�O&�9��bt��`��� �uN&��^�:(�޵Zq:��8j��M�J�i�M5< R�(  ��R�O'��  E?2�O�UJd� #��UBmR�  4�$�ʕ&�� ��<4w߃��?����Gq����왿�< ��'���IbKX��f%��bY�RĖ$�%��ffb�X���$�fg���,IbHX�,ĳϿ���x��"����UQ��cC+��FȚ� ���!Q���,bbM�1� A��a��� ��&�(�f��	�H�F=S$����#�6D �c��us[?����Q1m�$fcLc���2
&�!V>5^�cM���M15�bU�n3u���8�&$�flB�n��@ !�&`r��bf"Gǃi�Z%���:Sl2�������&a���+I&+xn�jљh+pxЄ�A���L��& �G��✙L�����X4�Fd�!���п|�,j.����1L�7!�Ѽ4ę�@�ɠ�X��01 m�1���o��b����������	@ ��m� ��q�*5�!��6��8�&bf&bA�#J�QW�	�l![��m #
�(�"Q�O���KȤ��oqe�z�]�;�yM��� �؞1,����Є�lPD�����Г�h$��"�������0Lf1�i�i �@���v�C�6�"���s��2��L"d��H�"f0	 H)�bA����P�O��
O}�k9��-c؄	I(���
�M|8��I~@��0m���9$��m� ���h�Kh�2��B�Bר�B'�Ame��9����~�&��m1�آ-��0�وQ�!Q��B3�M&f7fH1V�)1�	�m�"r";_��,H$7��>�q�|bYmڮR�f�	�'�)	/(LJ��V�ZI��aУ�Q � Q����m�Ɯ�+7T�kl���ui��l�!!kJr�6�f1 FH�m�����L�MD�\ `�$S�A@0�NlQ��ڿ���(�&ݖJ�X2yr� �Q��M֘T��1	 �@��A��4�(��Mrb	�uV�:���x�#0GY��e��F�ۥ	 �P�ֱB ��5��� ��'�m4(�I�&�0D��� �j�d�LLq�n��6�6��ۥx!~j0� !Ƞ�clCL@�l%�&A�!:�T���0�^ˁ�ң�B7��Ix�KP����x �i���Ǜ2%S7�Qvԣw�d �!�� L�Hm1! �1��b�*c���1&����6�F�e	IS��P�΄���%�|V��ګI�e��D�BV���6 �!
8�[�!�F!m+���S2�(�1��90�D��Q�X�c�-��і��/�.c��B\��m�4�-��~�GY�(|�O<�9��14 *cz&V4�'dQ��� Z1%�&o$�����\j����^�c�^u~П�8�`��&R����E#�[G�2 ��$�1�>i|����@Qs.[83-��� qW����e��M�A]�ݕJ�S�5"��a�3��>>$�i�1�@ؘ�i��x��Ph���9��q�*��lM�� Cj6 �  ,���1��rq��~"�kVc�g�Mf�6�ڍ1$f1&Lx �Yv�w���������AF�x�oq����o`���v͏k����ZB�X �o �DZ�B	��x@J�'0@&`cM��آ02� �<  �F�m�Q�7m1 X�u���w���5���а�dr��-��,��rh�j�n!�&>LL�2L�q���,�*�.�!ڏ�HL�مxՁ�6�g_g;b���0#LHF�o�yu�d�=c�"���),R��lxgW��I�	�#8Ӡ���>� ����ϧ?=���g���\TB@K�B�dco� ��i��,�!U��y����L'&�9"2	���RƑ� N�"&�``b�2F���`d%_����5"�6$&�&�<A����N}����(~���c�cx�Z��U"��RE��S�q��8�us��r#0	� I�5�p�h��oU�R�=��0u5x��MƱ�	8)A"��(�K��Hm7�<���e]Ae_N��ط�ԅ��O����H��}�o'2&��@�F1��F7�x	 @�1<��Ĉ�!�����P& Dq� T��ۗ_5�)p�-2�p��*�@
V�b& &�ق31��� M7���a��J���#��F����b�F0 0C_^�.	tT@��9q�b�̄�M�e�M�D"AH("�+i��� Ąu�;��� F` A�	1&��E��
�� �B	౰�6�@��"�f9	��D� z<����'X'��8�<� lBb���K-tDB��6�ѿ�_�����#
ѧң~g���5��Vs�M��Z� ޢ(��8�^IL@E�Y�/U�M�P�H��'ov�|���Su�(�VYPp�@&�n��F��*�5��R�?e�a��9�*�4֫	ǯT[��e�g#�����MH�Mb�N�BM"ܹ�xn��
���Jڙ�mn�_�;�Y�bFD��4�>���8'�hkڠ�a6�*T�\WyE}�}���#�Ǚ�aɶrr�;?V��6��NAGb�1!�@,
H�������c�̀b! ����4�b@"Q�D��i��]���y�)[6��BC��X�5(�:c�F�6�v���x��8���BNF�x!`bi��Fx��ݢc�^[%b�{�H�d{8Y��_蝏]q52ȉ�(��6����P5�%Ɩ���n�MJ*����8]��� J��!�;tk,=�@�hPh�D��fQ3<c��Ӄ��#i�ƚm�)V���lVE�.kc�#f�×,��)LC!��"F0�x��8#�"z�4Bn��1�UxVލ@�0lbT�,%2dD�j����L(�l�͑���ڀ�-��8l�Aq�pعSz���MZ�iU`�)�8[1�bz�r�4oL��y���[`��e�M)PR��H;����Py�0�HPAj�9pUK�� �a�S�E���"4�r��Z�IJ�j��C>ڰh�U�5`�!T*������^��6KR�ԍ��N");Ц�T-u�/8R&�=�m_Sj�[��ܧaU12c���[�R�,m�b��^Y�D�
��rD�4��%z��у�A8�
I �1U5�UJ)���)+�1��2�y1�2(��:����k-�{"�d4�5!1181��mȐ�/*�Q�S�O�j�:�ɗw��@������\5���QD!�)Sm�^3A���F��RHB@�! �$�@���&��҈���x������Y�fK������cof�I!��~�������3��ڶ�IC$��I�X�b�11&|�IPk�����C��X#	�FD�=���l�A�vpښ�Կ�&� ���Q�����r�ӫk��9�ܡ[�GW�(!�����Kԕ��F��-"
U�QC�L;��bU�UbTRs/ׁ�F�ŕ�)ڂ��lQ�@�KPG��������&$�ň1�j:ڔ��������?^T��CJ,���(3%�WP��,\�DTÕ� ��ʱQ%�4�$!_6���q����L��F�b3@�`, ��0@ @�`�͉1��e���e�QHٸ&�Xh�t@U��'[o�w �d��`��ZMb	N&�p��ZR�KN�q�hdb�7�n�e�&�m�'q��3n�e�f�.�G����֙U�{� �u���5xar����1��9�!lbQXس�82m��wl����;l�r\rDQ#d(���L���	��#M��"�<L@�fM��P��:�cD��1���z�"xv��`��6\��p+�gMH� �Z�l��]�R�4d��-�\[fE�U�H(��R+��J�+�L4�!��5�r�a�E XVٹd!Ư.�V��rd�����HyH���*��KU�0!ڪL9��@Cwn<�Uw�@���"�	I"L�h+x �Z���ρM �A�w�Y����d�a^�T���bF��3�*)v�A�땤 ��,Q���կ1��	�X �X[e��"�oI&& f%�y��B<8� �����e`k��;S��)�=�}��B\�i\�A��F$�b�$��$��ehI��%���*�����	��=13͒u�9�������@�6�C����۰�r��&Ě��J(�Kq�a]9H�X�l�je,*y�����&u�FM���z�2袆���U�#��%ͼj�KA`���b�b��^%F,
b�X�b�
��Ŋ���H��� ӭ0N<���:�_ ���3�$!$!vI���8�֛^ D��vc1Ƅ! `��i��
���5bP�Kb�@��&�M�j�dC	 ��`�@����(�n��[�+`8��5&Ƈȡ�#�Z��V-h���>~I$�1`bH�h�ڎ���01$#8%�B MDc�q8�H�&�o9l��C\C�1�d#��+��⿶���B�p~�9��&��1 @��˄.�>���J�%"z����dP�Jz�.���[�6�_�Є0�FPP�,��	���S@�c/5Q�P�P�^h��cJv�dѤ,�H8�����5��� �j����/�s���%6�@�*FTh���C��'�;�a��I�!���e�Û�[�XѭP���ۑ74�u#d2L`�#�[Bν�Ef�7�����;,x� � �l�"�%��Xm4H>T��yTI�-�$uJ����m�#(ůES�BXji�IGjl���O���Q6�w鶉�(�ZB�\������J�m����z�$�0�)�B��Q�KV�})�Ei�j4�/UXt���A�U�1![W�o�Y=�� G<�%5NP�Ç9H�~e����d�����C9k�K���}T��_o_+n-�lޓL�"0�Vꮐ�H�⛨m�!0Ofߡ��__��i��B�F��a�l����s'��h����Q�ڷfr��ny�s�g�W����9X@ �~����ܰ�&|�F��#�� �rE������i5�H�6�<i<����8'ßU4x 2��<q��l��C���[[A�#m84��ȴ�h���a�G�A$2hoe=�ܗU{l՜u�^F���e�-�\�H����h8�����V��.�z3����X���+h��-\�e^��Sjdi�.���`k��fI"A��њ,_[����4�䂥�����|Q
=��J������i�yַM�Q#e%i��q&��!���N��v�������@�pq*T��(ӡW�S>^����F��"��*����Fs[�)$e4��EQ�A Q꡴�
	�X�.� �Q�2]�wo�7}^�I�)�Wcs�k�L*�'3Mp�1]�6�~�&�R|�b�H��¡h���-ˮ��.��س�)�+�f�6E���V-�+{��wOI�-�:���[k��V�]��w�P�TJ%B1	��4)Q"P80u$��˶HD|���i.߅i���vhMvni^6��r��U��v��!aX��w��7:���n���b����D��bK�y�st������2�#iU�Hu���\��A��ꘕlL�h�L�ZN	�}��Ϲ�� ���9��țWWv�}��5�T0��c[Ei�khOt�]d��Ud׵���CWg"�n�آN�c�1\�d��r�Xc�^�S�n�s�4�[��nI�	�t ��@���H	$e�n��n�,�-� �I��ـ�`�RF��J�l26��b�S��M	�y�P� ��M��
�pLH�"
�И���F JG�5��A432��VӐ��4��4����4f	1�&��'��'��H�!Dې$ �ݪ�C�� Y��FM��(�8e �io9�50h��T�ZEj���Z��]��gs���vv`�-��H���A/J�Leo
F�>-�ڎ7! �`dҽ���.	���)��C_�R�Rۺ���2�X#��`W�FА%�0r7M�9�:6:�i����"1��I+����a{@M))�Gf��%�B`qI3d5R�WnԸ�9�!���*�G���� �L�$Kt #*QJ΄&Wf�*���T-�i�d9�U��'f��5;l�PlT�R���T�vׅYT�I����L��Vؠ�T�)ʲ��*��Um lD��!���%��e[�V��� :Yæ�UR�X��`]�&Wm���i��,��E�n�YBk.�v��*�;�͙�T�A�,�Q�T��h9�j[��TFQ���R����7@$MY;<�@[5MJͶE�e�*5�
-��@��T3�B�mV����j��Eہ���c9��--!D	-@*��=�@Yd 8��6�Ό�' 2��f����N�X��r�;�JJ�T� ң@��e2���@T�US"i
X#��Ԑ�h��`kpT��Ы攃���	VV���O�(ԴV�HMUT�J�,��v�*��;T��X���y�%y,ƍl�v�WA���U��Z�P��u�m�tR���'y��R��! 3jB�*�E�j�[SR���tf�U�Z��&�btT�f����ZV[T<b���W�_��]u5:2�l�0�E�k�+��.2M++!-UUUJ�6��P骶��(B����ł�P�V�vZB`,�W)��:�Ի9�&�[UN��t���N��@S���ez�T<��p�Ed��ACa�f�Ɛ���IUUUT�br�rr|E7Ut�f��+�� g;0	Q��ͪ��j�JT��UUUJɝ���'%�W]:-����RvK�5��r"���g�����e�u��ō )�$�Aa�V0�{G[(g��EvEM����E�j���E��a���5���K�L�ևT���Vԫ).fnU���v��zy^��-��R���UJ��X4
����54���jj�%�uR�U@'L[tt��KQAD�7[l��,�If�&W���VXUU���n����c�s�kI8ܤO\�v�j�.ٝ�]�a 6-9�ۊi���R;pi��>l�6"ݻ2����+�Y���3.�(O[�Y!�W��<�q���lEn��[�	�3�P������4rW%s��UUL� cxv�Ӎ����
�8�m�٬Xu�rv�+g�P^]�vC�۲�����2����H4�r蝂��6ӸY��2o�����$8�Q�իa�c�*��JY��;!ۘX��B�q���}ۂ�<�;b�+��9a����QV�eݢd���Q�5�!vm\��"�jygf �e�7jmd`��f��ֱ�V�i\��]:�)Á��[DuZ��g6$$hV���y�]�m��9I������� ��3r�Iv��\��k�L&�N^k�ϏN3S���C�ʀҲlu��uJ�)��>/�l��6ò�;u�%����tX�2�G��[K0awkIv 70�)�xĕWp����R�]P�l�S�$N	��IL�`5���m�Q{����+@��M!+�\�#����7��Ơ�Q�Q��3��wZy�MȦHpZ:ݬDm΋�S���e䛩�Uz�,�Cd�kc8��K�c�N����;o�V��nV�����&���[����9�Kخ8x.rΫ��=�f��x�9�\4��*�g2mY�>-�sv��݀ۙ�p�t��*U �ntv�f�kU��c��^&ݲa��Mm�zvW��6d�݈tOi�rn)���+�֗9�ܖ; ����.��cq~����-+��s
�/Gn��7lw\F�wܱ�B�E�:-<�Ɠ`��M�Ba�G)@t9�4����6���8���`��e7ZG�d�}����}�h͕�n¨؁&�Aup�3�)���a-K����X_Z��}/lY�q�'���'!�5���s���Rl�@���X�����/-�����c�+��!�v���X��V���	�ݶ{8O[��+�;�`{l��n�I��7M68�D�%qFZ�ZRR�n5��e�H;3�덱�X�śm	J���f9�����Pyq]̛km4��֥#�ݎ��\F6�[p�p�]yzn�\,dx�҄��ل�96�[s�Nҙ0��
�v��)��z �핣r�S���T�PpP�=�^٭	����ݴ	�5k�[�	�`[m�˖�d��̾��]�ٷ��8k�`�r��9�4�6�U�*�R��볗��������`�qg��m�[<�W�!��7-�g>lc��c�&-�gGn�hI9��v�Ϟv�I���g`���@�؏A�ų)����ѹ�k��M�%�v���)v8���˜a�VI������κ��gG&�	q�%7v�#����Ӆ$���k2j�@t
�QE�U�(zn�H�Stl�hx-F��'�=����U��=��]�%�����e����Uk���}��w!1nn�ӱ����po5�x���h\�n�k�0z��<��h��9A�ܘ(��l��'aeR�����(-�*�Wq�E��J�ԛI��mUأ!�t�:\�v�Rp4;��p����Jჲ�p�1�N]��'��es�q��Y\����4Wg�YV���c�E�lR� �>��fN�8-v�R�7&v㓋�Rs��Y�ɺ\=�	��`'��y�Un�9`wms\����T[���<uȌ[����;v��0��B���lge����k������qeC���-��$�����\�>ۅ.�c`
r�a�oY�Kkv�8���"�d����Ur=	Ӌ�g3���Il��x|��U��؀�]8�v.���f�̋���ðz��]���ɺ�{t��m�4hM��^	J�)��p�Y���`���zCK��@���,�v�<\g�
����N�p�Gca�^Ig����[$����[���!V��ڪ�י̙�mQ���{cr+�C:�ɫ���A��,��7yd�ޖܨ*��LJ�Oyb#��v��q�f��U<ఽI���mω*�<�����9�Ht݌��t����Χc��l�'��[j�F��b����
�e�I� (�".��p"�6�J7w[9m��2f�s�g���l!�S ��� �n�ѥD�΅�95�g���т���n���Ec�A�2A4���K��D�v�%$]��]g�8�#)j셥;mh�˞���aⓇ�1�R�N�lY���F��z5f<�%aLg�p�ηF�8�D���tTOmfێ�톻7O;9ٌ�
P:+�׫�-��$�m��b��ӎ�{dͲ]=n�^�n{x��g��an�s`�GO8�`.vvK&6�ֻ<ڤ�k���Nj�_�ur*r�(�G�	�4�
`��l���£��f�2P�]��8N�2��FP�u�$lq[y
i,�۵)l������Gr��p���\��'%�:{[H=��l�c���E��pn08��:��#�i�� ��qWh���qkX�)c��\ޭ�<e�6��-�١�]�;/u��|c"��4]5�4�M��2 NuE'�k�5//��n
��+A,=<�$v���Mͬ%��\L6�q�y��jwd�P�!�iX������`�M>�j���O@,�%J4���o��i����E�{G��RK��F��;v2���:X4���;/���H�]p�O7lC�z�議�5!���g+��We�5=�(��� �ej�.97m[�=�u�4��pr.�r���n-2�7�q��7|�K�'$T�k�����qf���۳���n�㵬�3wY�{]�m;N�����A��Ŋ�(lS�f�&綶{wHQ�[#ce瞶���cf.s��f���u �M[X�����P2���]Z��:u��� Ŷ��*��6W/@ڻM*Ncm�U.���bu����,lpɹ����3��f)d�R��z��N���$�.�v&S+�#���Ѷ�s�@�8F���ѓ]�&�\{Q��rҩ�\Vf,�.ql�x\=�U�X��m��s�)O]�1�*Ս3�I̕��Y���"s��,�K�Ld��"�FŮ���Ses˴��&���۹F5���>���q6�@��Z�d٦�����m����b"��wtU��;����7Y86����]���V�a�E�C��i�[jOr�g`��m� +�ܳv��FD�!H6Ѻ��W�l��M�ĉ���1��l�s� 5Q�εX�mι�7T�؂Y��@�pU2�kN���s<7��ѭS9��>��t6���-a�n��|}|h�\+U�NL�q��Uw;"�Q�9��5,�C�m~;m���泮��4ӭs��S�2��I��[Er(���:s��� Kt�����d�
�s:Q�`�����ﯯ���)'@�f�t���VX� �x���۔J��!�gnFxm�S�\f4z6�.���5q�nRcZ�ܻ���]G�1y��q+<k�4<�HhZ;��`b�v�	m�m9:����J��p)-.��P�n�m mU]HMT͑j��������j��ER�-R�J��UU)-UU) ��6͝���/*�8��J]AM����u�w�)۩5�ͤ��g��<��87i��`�(X���c [��	������j����E�V�H�/m���M���3��� WN$T2;MJL�8��K���:8��[i�UUT�J�Ti
�������VU�U��-J�UUUUUT�J�UTUUUT�+UUUUUUUUUUUUUU �UUT�UUUUU*�UU)�UUUUUUR�UUUUUUUR�ET�]C�&@D��\��UU*�UR�)-U�
�Ԥ��DUUR�����V�����j����P��UUUUUUUmUT�KV�J��rT�UJ��5EUJ�Y!x����#���Z��>z|�N�]�V�),��Ykq�u�ԄԪ�J�9�,UUR��UN���j����Z��+n��j����P��������*�KUUUS� �P*��rJ����X*�Ns*�Y����������U��ZU���������������V��������
UZ�(6" ��Z������U��T�)!�LlUUUR��ԫUUUT��T�UUU*�UUUUT�UUUl�ԫUUU �UT�]@ͩ�	hԑ�U�6�b���`nڠ %���������m�UUT��Mju ��UUR�%]�Ւ\�g��y40 D�^xl���6(C�s�^�bY�f%���ĳ��bKX���)/���>�:�T���D���m�U�6-UuT��$�3:8VS��<�'/R�Um8��\�C���m�W=UF^
�`Z��T'�6�j�`ېVL���eB-�KU�U,9�Ul��5O�#!6��%]��	mrͩR�s��˚Q�eZ���Ť�V�Z�8���A���Ӫ��5;3�I6��[�;$ܬ������`P���a��q�:Q�iV#tqp*k*m;,�3��v.s�aM�nL$qb���klt��s��v'6�Y��ږ8{ ��M.�	��q��jR8�5��7N��� �ʙ#(ݘc-�'\J��؃)��x턗3�6���Z�#8�\�������XD���8ζ�w\�p�t����sk/8 �v��8#�y�=km�������ק#n�Rڗ�!�Cnٛ� �n�y۳�s���,�&�c��'�7r.�{Θ�f0�{6��m����u�ȝZ3���ˀ�d�/�3�L=�o%��\ܔ<{��:�������ifhte�Z��90d���c���=COJ��v	@9q4�r����x{+��m�^M��h ݻd���w	���.�:��۷"m�NY��.��^�yb�x�۶Hڲ��F{B+mM�Cl w=��M�6��k��
�Q��rF�u�UuXr���M�u���gm�u#��l��+Y6ݓ��IH�Ztj�f��ol�\�6DE�=��1ʸ����SGjk�!���L��œ���8xݵ��Tv�Ŏ�b�z�h���.��ݛ�����R�c�Q�uj�w0�n6;#��x���;#H��GAJ�Dd�N���������El���d*�G��b*�)Ȝ��l �����v�\�q���R8�ǆ�!�=��a1qb�]�֕�8+J����کI���d0wHZ� ��UN�d��*vЁ*�JV��������j�����mUJ�eej�yZ�j�j�(��ʗ(�@��[��U��8*���P�*�zPe��Z����W)*��HM:A�j�ꪦ6z�]�7�uU5;uD�	/�������u��;��|��F�3�90��p<ĭ��DwW>QQEd	#p��NqvxԚ�86C��T�C��U��AK��zz��)��ѸK�fM����:īۮ��X�m��1�84�y�����\��I��;b{X�$�V�۷�iׂၵc!�<��֬�
�n�eC�jyd��ٰ�)�v�N���j�z���SS�\�p����j���p^��=��S��6Tȏ8C˱����v�.��9�r;��.���r�&�/��L�O�D��B��,��7t�"��Κړ��/z���Qq�{�Z�X�&c��I�0�Շ�e�\}Ɗ�k��dP�zqg��	=
�\}e�Mð%n�%��iӜs�������+��OZ��9�ѝ,�"����q��G��$-�dc�guaE����h9\}�O�m��c"�guaoUd>4]���Ѻ¸�nRYut���q��4�Nȫ���\�C㚬�g��c6g�am�֥�ʃ�q[ P#`��֧�\3M��4�uFL�We�u��V�S%�h
ʪlfXA�u���V��Di�O�z4B�]����q+�:Y�a�i̄�"PN�JF돸����(�ZF�e�H��oN��,w_*�.!��b��H&T���2R�)�t��X�d\}�:a�i�ՆWq��B��v+#x�YmH	a��T�,��P�a���sMۚD�4�L朎z4E��z����+�G�q����
�3Dy���f;�dYg�hy�e�d.�q��]���|��8f���h�c�ɷb���1�%��I��i���0ظ�G=���i1@TE�/`�c�눸���u�8�����c�qt��:Y����q�p֑gM��n�p�\A6`F&��B�EDP�xN,�-@t�Gmqp�Z�="]'h�Et�Ϻ���R�:�dv����V��3���a�w[u�Qӆj�f��dc&�i��,o�P��fK ���VG0t�u�hi���[c�<}�cCME�a�>�C���ӱI"�"FTnEZE�6|���C�EDP�xN0�-r&�qp�b�="j-���2 *E���&��5O<X�+����'�v��-t���ݮvs��OF����6ۄ�#�AƏj1oP��iUh+�<}��$�.��t��P��+e$��L�P2#b����.�i�VG5�_J�44�[ˮ1�>zΞ��E�aU�$�Al�$e(x�9�6�qx��Cy]�#��e��H֮#�/�̩4DFH⎽"]'��I<}�C�CMŤa������r`�n��t��B��`FH�fOg!�d=�i��K�|o������^����ou�8�����?t��S�\�œ����l�Ë{��˝6�kmvq��ӻ��]v����7��-8�EB�2����s\x��:��*�,��B�/�A�	şe����B$���`���VG;׍�F���L�zAƏj1oP�qih=Rl��s���?�I~�(��b�W�+i�5v*#��MJW���ج�6`�|����Qf�$:(2L��"c�<}�J����0�ˏcA��v�24��x���XC����F�PIqg�hA��;k��_c�^M5�y�Əj1oP�r�gg��X��)H�Z6J#*fh	����ݫ���$v�])ǎ$:��bȘ;nU���pG\�v����l=6º�mŊy��ڈ��cPs����#��V���7Lml�Y�;mc�Г��x-RI�1�ޢ���?������gs�'
���E���܍�ܯ���'��#ص�fv��a#� ��mD�Ѭ� bQu9V��]uUmVY���<y�,v�� ���W�p�aX�}��܏�ɓ�u���nys.+u]p\�[�;��kv�ÌK9j��`��bUp�;DNXxϼ��n������TFj�TFgf�>���ǱY뭾E�I� E@⍹�8�j>�ͮ�E�����5��w�kx��Au�9!��06TC9=Bo	şe��H�#��*�W�!�����H�i�'ѳ�"D�Sݪ�4ݺ4�ZFI�g!���\C:p�TF�t�f��4})<u4�0�$*:�Ӧ���t��w6��N�\L�g�|l�p�!�e��A���$`~�7gf3gSx�n��m��
k�ڠs$[q��n˵A���#[gouF)DZ�V�gMs�3P�ƈ��	��m�N�(��8���w%z�4y��L���m؛V���k]!�?'N�WN�|�w!�q��\C:p�����&D����#H1@�+MJX:�2�Ξ��}��,���6Y��ŝ����}�HhR�M�c���e��CJ畵��<p�k�A�p��M,�mBuqGO��u�)r.�*2�(�JCM��B��G����q���4�ў>�CU�+��Nt����\*C,c�mط6G`�WaҼ�ڍ�ڋL�ї-�l�AhΘV.�)��Q�������]4���c��7���f�K�^����yu�8����.�Vш�P�<�N7�;6l���}c4�24���yC܃.����e�e���Ԁ<���3��=���n�;u�i��B�ю4x�B�z�kH�L�]���0����=��\�@d���#]1z�������Gҕ��ǱYp��\�����=$k)sI8BM�%Ia��b�j-#ŖY�Z��6�24�҈x���Y���}e~6��˵dDs���GV3ڳ�3�MO�Y�ڮS�����[���vH�l B�9LW}v�9�=��ㆷ�<��Hi�����Y��
�]9_��/�����n��*væg!���눇N5��v*#��MJ]���dqüs�,��Ir:�44�\z�1Ş>y��5���>�\{`����:l͋�@�B',&��B;U�j��7��ϲ�'Ws}������֛�!ޑ�Ə�L�IwA�Y���O��gg	뱃���U���;Q��Qج��NO�\��-2��lp�������]�(d�Km���Y�o,;uzֈ뮷<��a�a4\�VG3��J�5����i�0���0�i���<x����:�;��<��j6J�ȫ����\���Ǣ�(mp�a�Z��.k�B8�۵��z�i��V}��j�ە���E�N�|�ޮ7����z#���U���(�!��ب�w�"8�$9�ACJ�Gҗm����㇪_J�5����k�-��Y}ָ�mL	'
s���SSH�Ϲ��q訊o
�Ϫ�'��M�fl���[*���d��!�*����Xf3X�XΛ����z��6�/0��u�x絋N,T	�t �Zt]t�[]qh8�;f�rh�1n	Ue^�Ԙ���ʉƗ+��ܑ!9:�R�e�'36�b�#�"Cf��z�t`�����ˎ�nQ��hM���ŝ����Wm�k��vu�n��"�;��Z���-�#u*�W��CHrͤ&��SLp�ԛi�#���R�GE�7mW��$Q�9ٗ]�:۬㗥�sI��������h��}�\��ݰĻ!�,���灝��x���Y�YW[}6�Y'��L%1�dΪ�G���V�o�����8�[�A�;>�� ѱ���ۋ�y��o�v2�?kA��eU��"���XF7�qg�hn�$!#IFX(ș�P�8w��^���k\�1Ə`P�P�qihl'�<}���f�$�J�DG#u�QӇiB/P��Y��h�R���+#���ש���ٷ��� �!v�v�є�-ڻ�=�7��m���zB��7.�ŕ�aƴV�W�\�!�
j�pq���臨i���<Yg�h2��5l�x�	�#܃.�0ר�B��(H��A�V@wy��콡ʱהCMŚi��q��ڌ[�8�ZFÉ�,E�I�z�q�>�Cw\D:p騅�v+#��MJ]���dq�]9$��Je4�,H�n:�44�\{�1�>{�����0�����q\j��Gm����Tf%%0`�!3���A���k������u���Һ�V�DK���Z��p�)LqV�q�z��W������h24Thj�:r`AA����E"�t�h�]ou�,l�t8�t��Q""��:�i��{E$�8>5$abt����O�s{7(�6x�Sdq�O�h�0�"Ν:}�i�86LĹm���giՓ�NM��x����A���� ��X�@�f$�b��@����bI,�bHK1b@�,�b�X��!ff�X f,XffbH`b@�X�@� �İ1,B1$�bY��b1fb��I$a�� ���� X�,@�b0�X��� K%�1f��	b��X�����X�BX!%�HX�0��@�f X,Y��b@�!bB�`�1 H3�3$�,X�,Bĸbͧ�����1d�,�?�������w8,@���f#�3?ŋ� ���UZ�eRZ�/	&b቙�1�,@���IS����1��� _	&b�|�vn&ft�,@��f#���ʻ�znpX�bD�1t��όb��ʪ��$�F�L̟<��h� V�A�N��ܬ��jK�.�������I��ӗۉ����,G�@�$��񉙜��znpX�b�$�G^&fO� �{ӞpՈ��1S3:c X�_���-1<L����� _��1}C�(�6U�0k�n��wZ'e'��.x�+�m�x�k��,�r��Q4`«<I/��{�1�a�Lfg���\�b:5���1t����1b�%X�|$������אX���zs�R\1t���ň Z$�����sq33�y�Ѭ@�$���3;x�*)dn�!�l����I��bffאX�gy��V ^L��3:c X�>��%L_����#�@�L���o��3:c X�|b��Yz{}^���if���Y�<��y6�Ћ+!5,�Ś%��n��|��qgD�LK/�� ���|�C ~!c����pI3LL̟�Ab����X�xI3�������w�H�8�h����z�ዦ&fmy���$�^~�������f.������j�w�$�����@��x�ŝ��k{N�yn%�gLLIp�f �@�bLXw[�<��R�7m
`�{�	.�y�h�gL����~�%��4�Θ�ǋ�K��xu/E�3}�fg�:������,��Y�1g�~����܀��̐�&��=8�\��Ђ�y���i�On�=�tW@�gjhd�M���f{��@�Ę��&$�1�N�U���S_W��F�1�N��KE�11%���1�b�|s��/~y�~b�b��&-����b��(,鉉.k�f/��е�R�J�l�� ^13[�kf _.��h��/C1b�b�?LLIx�f >�̂����ӎ\�1b�bΘ���c#�����=Z��<Y�p_ �T
���������4�Yx�2�w�7{�7^,�����廘�u�gLY5�����&�4�p�ė�fb��u��:��P�GG��tĘ��'��R4�
VFWl[��/���|��z�����xy���t�ė�31v򫘁~�Ġ��&$��!��1�/Ϸ�gLLIp�f �@����|~�ŢK�<�b?��_�LI{�~�)%c$�;-�s�b���P�����{���x��LLIx�f �@���%�Θ��漆b:<��$Ş~�����A��~�Ġ��L�Ӓn�@�bLY�_�fb�����_��UU��mm���q���@(2����F� �Hn��}��֑q���Dn������V����څC�W1����69x�3g'k�V�m��6�dU�Dޝu�)�͌y�A���kcsͱ�H[p�9�͊n�^-z�F�����ڷV��ڢ� ����]�s�Ho���U�)�VG��U57P@����9U�j�BV"o��_q��#"�F��v�\�w<�sӺ�ț�E�l���m�ɠ�5��&�]���O2��g���,�bbJ�<�b8<�
qy��n%�g�LIp�f �@��Ġ���Oq1%�C1<��$ş����}�۹�1b�x�x��漆b���қ��xX�7���o}en)QK+%�
Bs���d:3��^����6ސ8�6R�0���%K��TM���/ϵt�]j��� ��M����W�������N�Q,�ڣ!��8bG�Xv�a,�ʢ�-#5$�T~��� �Kc��d��<3�E��	�ϝQ0��GJ5<%z��jD��Q��#���bG�9�}w�I�.�q�������c�3��l1#�D�,;30�U�Qe���L�r$Ir��8&���ϊ��o!G�r}L��+mi0dU�mN�ʝ�#����ۙڠ�sQ�6֥���U�Wn��N��q�^JT[�f���'Nu�����������a���A��F�� �BF����,􂓃H�ϗS�q�S�'j��������!l�7hj�0ID9E$�W�!���7�,�4x�B��it���v���g�r��M�U��p�D�hF1)�����)i�9�h��'����G���Y3ҷI;uD��d=���l�����o��Z�'`U[��t|�������`~�
��UfQ���"^՞uD¦U�����8u�́��=�Y�E���{pݺ�]���9�X�N�{l&�=�n^������
ڐ��D&,��-��Y�f�?$q*�<�d���ⲛ�̬pĎ�a9c�V�!�ɛc</
�~︿�P������7����m��s�:Q�O0��$�Fqˇ:UZG�l���JH�V$킙�h�;E����͚��.�t�U�YE�b���.��^�d\���[���Ot����,�)B��D�q"�%ř�Qč�Yܫۤ�H�V%\̬p�GR$��$�'G�Ό�g|��'�����W,F�6�^�8xel�aٵS�a��G
.��{��I'1����#J�ߡ�|TV����a�̍��U��D[v���΄��=	����AӞ9�����m��^�����C[ =��n�ԋ(��P�$�H�=pʱ����6�r�pKJ�n���*'�u�5�(�ZY�h��.�̍0��F f	��B�A	BD���ejMy#���	$�D�P9��L(�E�K˱g��y#�-�=�� �����GZ�!�Kn��K�ɀ�͵%#5Y��H�L�&am�:��� 6|�}�>�FzF��P�[9��?6u���u���٥��P$�H�-4��6Q�GR�������l��'�>7RS�h'�e�*�m&����q�g���0�mp��bv�P��Bvq.2��P���H�D�|$����QiƦP8I'�:�l��
6�in���F��Z�7��nv�7a*�$����l���i(�GRs�7I)"�����8ZG�[�3Kr���H��Q�W`*�TKd7́�����{��bE��7��HĜ�:Q�:����"N$b'���!l�U��̈�F9j6du�t�X&�^�G��-馱#��I�2$I�%a䔷L(�g[��r䱪&�Z8�)��#~��Ag=St���'R1ꙎUybG��핺I��Kު�О�bG�_ݽ���Uf�����F2��V�Ћ�i���\1�~���	F�&J8Kbٺ��t.����ps(R�N�iQ�0̄��k-cVs��4���F˱��wی��>{\/��dr=plU�����3��U#��������`҄i�Ö5�;����t��_Br�=dwWW�!)���Uۅ7Fŷ�&@j���<*�J��+G�2�I��54��9m9��0�d��=a�w�m��Ϧ��cђN�q�� ���&�
.�6ԼE
X(:��Ǜ��xg͟���l6y�p��
1"��F�e�bRUR���Z�p\������`J�le(]qf(G��շx,�k<����X�GR�X�3	e^�Qi��9$�����[M�z�;*�-�s��kg�ԫ�y"a]͜(�o]��"N$cn���#>K'�VF��N����p��h���w|-</���n+i�.T"qI�j�yB�W+�a���;��~c��0����F.��ZD�H�OrFo6h��J�9W�t����U7�eZbGR�X�7C����3������cqIv�Z`qr�XM��ں���hM�5�����sn����hM9�X����F��m�|U�6*�0���$^�Yi�s���cUպZZ�'1��IU��K���D�a��	JGvIiAe�`�z�!a��<�j���B!��ߟ����C����B�T#.�z������tĵ"O�6�L�7�4Q�%���+�M$OX���:P�͜ó�=�҅W,Q���Un��ܪ,���fP9$ď�V-�V�AH��#�*�H�)���{�ݞK$�Fo~DA��i8�AU����#>K&zV�&�%���^4pĎ%$�nf�ݪh"�1CQoo1�����Pnv������p��.S�cW=2f�0h��8J�Y0ml����a{��+����o����H�S�GJ2��n���I�F����٢�$q+���ݒi"x���=���eID穇z��'�9�L*����H��fQȑ&$O��rB�L(�E��yVZD�M�~�����i :���ǿ{�{N�چD4����Y�#����Y���^�a�C��BH`lB�F���"�5A�F�awP�:v+�(���J9�B7j���b!-��q���Z6�'�meF,�-'`��"�7���<Z���14m�
q,���nwcN���X �h��oc�����;�1�A��<����!P��C;�YC��?#��L�!��5�"<oS<�i�>=��F|�N ��JP�Q#�b�fc��L{�뮸�ssW��`��SȖ�{ξ�޴��!�1|%wͺ�$�{�D�R�8Q$��z�r6�Co��y�:&�=X���vx�I';>p�D�Y��(��.�8�����~��������}��!���VU+��y�<�%�S0�+r��G�1�$��eP�k0��H����&�r��F�>�y�F��n)�"r�0�ʛ�rWn�%��mV����1��%��Z('n9ӷ,nX����p
�l�G}��4�$��[u�I��������6�wۡ��H|3��_&}�Ԫ-��RXo�͇�ޞ��������$M��޴�]�i"LH��=|o}!�g�������"�&�l�[m� ��������:i���`|���x�ڣ�H�H��M;��]3�oX��Ԏ�4[X�n�\��ճa^9���z�U�+���W^G�yu��.��?��2�dNPN�R��Hak���qvq�r��2kD;�Y5S�B���������ǹ3+��Yt�3 j��h��n�BHu(eIzU.�*GZ�W+���#<���AUI�h,ǛŶaP�2Zz��
��&F�� Y��W����PQl�L�hAؖ�B��5��U�#;l��n8ٕh���vä��+�2mK����YZ��˹�tme[�W�VK�H���V����45�\�+J����KH���Wg-j����P�!�!��;.��Zr�&`�+�yՓvs�ա)�kLdPD3���"�ϴ�u�,h�Ͱur�#9Z��.�p��F�6� -�b6�F;l����]���1x�<E�n�(Ǵd(Q�<�u�*v8�g:�k��Y�yf���֩��K�F8�P�iڔ�Bs#Tǂ� �M�msI-֠�CL\��y:�#�T+4�uz��ʏt��Y�b�(W��{�z��Aݏ[���q�۳�����q�\]w�9ڦ��u��'�o(�cB��q���I�Kgn��͔ٯ,WF����+�{n&�b���tt��޶���;.8#���qY�m[Ok�Pl�:w�]�iC�z��M:ݻUu�n3�\d���8ּ���LBggc/dæb�n6La�lJq���.1Z3�Y`^�E�����8V��c�ŋ��i��b;4�Dt��ϖ�u�C!�ۛ=���>����'l\[d�ۨV.�9����E�n�ݵ/7Nt�t9�W\�m���m�j�����vD8]�^Ln�2��wS�Gml;��}v�L�Rs����򁉲ݸ�6 !eՑ�;�,mŹ����F2�r	�۩ì����km�[���� �V�][��;v-��a�ѓqq�/<���X�f�JV�ؠ�\(&3&�����.�cp:�*�^���S�������4��A�m��1=�/����vR;F�Պ���r� U��)�`�EUUJK)E�����GJ��Z�Sv�ue �j�j��Z�����@�YZ���'�R�T�UN���P�IX
���F��@UR�1@T�T�(Oj�����U����U�:�V�v���ݪ�Pl�<�n2��$MT��[��lm4g���X��%
V�V��8@��c&,��Oo����o����I�V�6�n]�sI�ᅺ��Ĥ�:6-#�2�m�g�s�t��KGLyi���R��.����d��Z�A�n��[�B�q�[�#IήN�n]'xƶ!M��ͬ{nl�c
/j�p���q��`��Aq1X��ہ�v�k3��v�k�D@q�Ld��]Jd�<���YX%m�*����2k:㠡��d�wg��]�ݶ볙�	�5�q��mtی���D�;CFx6�q�&e{'3$����p�����(2/U�q_b���mٙ��W�G�<��&�%�K*�z��]�B�e��BY���8��'�H�*J����7I6�'R%�ܺ8�QҌH�obۭ�N$O���n>EB簙��;��6�'�9�K*���G�;n,$ĉ�V�Hot�G$�&�M�E���oһ�Dղ�!YlզSߑ�ӽ|3�wX�!&�'��Uʞ�bD��%p�C�ݓ��d�s��d,�Ȝ��Z[���a�Λ�֙���~�^��&�r�PF_����M�Iԉ����f��g��y�ɑVN���NqGc���\������+^�z�^܎�5 ��sH���4�<Wf��j�~�ރV%���T0����$�3	ejMZF���r$Ii�	+0�Z^oW���QَUS%�Jgݾ���8~�#n�j����z^�&�%��E���iI��L(�f�ZWhu���s���g�|�t�<�l�aeP�3(ČKR2�ˬ1"l��ҋ�uQn���<���wi#uX�wUJɵwvr$p��>K�[·bGR&�12ϕ-#�4��,l[.eC�?�K�߭��SFH�1���\��X���۷���7+S#K�:�!Ż���=�u��V��SvJ{g6�N��ZӞ: L�Aj��t�u��A�3�nԭ#��V�wz-:~�}W|�<�̨l�1�e�P�t�E=Y�L�?��������7M^4��W�*m^CX�=�JՐ�/�^�X�ӧ����	��M;���T��,qZ�Q����#<�9�VD>9Y�!pT7����X!���b�Yjdk�2�ƈR2d��$�w��u)�o��ދ�i�{¹����1�v��D�0�$#��MT����x�C�Zu���0�8��!�ZS1g�c#:X��U���N-��ܩ��m�Aٱl�9\��0�)�p��K��:E���[����T�U�Ŧ��2��X͖Fyd2ج�t�gL�m�kTbo]`�L:GT)kS�)u���D�|N>��}z�'���i�dag�@���3%;w���HZJ�Ы���Z��SD�d#18���z�p��;!So$Y��\:�W����*D���%.H��,�i�O
X�-H�pͬ��#�Ð��a��_L�Qqw+xL�D�%PIP�F«��0��Z��ء;=�DC���׭d�暒�Gնͺ ]�L���yX9̓��`�5�vݸP�-�pbɣl�v9.�-��p���(�'3�Qx��_(+�.�ݎ��s�vB�^H�T#��'ƨ���@�eX�j��U�4D9����Y��(9b�"�m�6�0���$J��CE�~N���F��r�yߜ��'�D:a���n(G���p��\�}�f�Zx�zoPx�r���UX��G�+�Tx�cO�M=�v��7�ڻ�?��pR[\R�봘���T#��J���ȍ{�����#:X�������E�z�.z�%t��%l�=�-��A���a�m���1�sR��]u�Z{�����'t��p	���ql��,-q��yꀖ'clv-���ݣ�g�v6���c�����+�Sx=��y���
����93����=���%t-�Ikc�G�/$�faƄN�Aųl�{�e�������+����h��U�5FD��UT� �4��m�3a^�%���0�[�����1�غ�n���:�@��o��'�3�]ƶ�f-S�d��tN�A���,��^l����M�*	���f�P�cj�#Lϲqdo*���B'F6�-� ��5�FF��k1Yd..�"�P�j���#�{�|-��t�=�*1
IcDT����g�u�6�#TYs-8q�Cky[�2�Y��#[��!��HX;h�Wf�v��=��w�~�w|�q��k<N[�i�Ď^��D	�'�6���ֹ�㽺�ӇV<Vumo��o���.J0$
�+fьg[Gn��S��j����b��ʰ։iDYd �2}&�;\�����=׸��#�6f��;���c`Fz@�(�FgU;�ܩ�uû������[��ޟw��-�_Ob�VƜ�0]�1�e�����DsY�{
~Y�0�fX�UI�!i��6�f�Ȟf?؈ұUk4���Iy�M�4�l`�3�py6�VYs;x͑�g)�ñ���*�6�Q7M�T�yw�{�qQdd�m`�ȽN	)^�!��S![_z��_G"�U(������j��!��¼���M�֙��w5*�hI�6,�@t��"��+d���Q?#��j�#Mͮ0��yV�B,�>��{������:��p$������C��]pʷ��R3"�FZ潉ߥW�D>#�ɵx��L�.���ꉵt-��Ы�l���LN�6��0胥��qLP��f�
,��q�XD"eb4Gy�DE��*9_"�S��>#�.�8��&G�OS0��<�aO�Y����W�B9U��
WZ�W�w_�x�̡E�mW*�(D �k!���S���P��������6��*2e���q�\\�ٶ9���r��З�� �n�Xe�ɝDY�Ÿ�̪Z�>�~��28��*���w����0�: �c��W#j���"�x���)*�Z&��NXD!�+��M��pM���l���6������#����N�S�#
ءka��g&~C��s�R�x��У�_'p�ء��d��2��+������� Z�(�-��x�Rn��;k�>���CDtXX��o�"�^�_��v�;��V�RX�p�`��/S��\���wS!kƼ��W`�CD.d��Z��!��R�еD�<���{	VO����[g]���R��ݵ���;VybD�f�L����w�[,�[K/$���?!�k},ww���J��9R@bm��.�P����t�%+��9wL��i��\�H��"�m5!�0��NdwZX�F��k��Y]�cI�h$ɐ�ȉ�yt�L��u5k��fݓfX�^�\ĉ��F0�H��}øty&e����u������i�����(eJ� J�����.B`�5l��"8�luM++`�'yh�j��ʙ�KG`�TNQ����<�xn���ٷm�e�Gjz����ݭ<U�������v�ZAi�����1sv�ut�np����X��v"dL����[��=��6:� �nj�٬gK��6F�������W=�54tWlˇ�Ga`V�����I�]���9Hn5H���%��x����2q�&v��VܔY�9L�pym͉�n�k����E���MU�Bn��hw7=���߅��ߊ�m�S����C#2? ��\I�����3we�Ҷ❘7vMf�k,�B
/Vyn�iOv+�]c�����̫����N4�f�R9��֜goj���gh��s8�J�y��i��q�Y�æV��^�̺A�ۙ��\[ܹ&J��Q��`���O"�.���mV�{u�
��M���ij�Ӓ�m���6�;�����Ǳb�Kwiٍ�Q��ub�d"C�*#d$�w�m��u��N��ژ�����]�h6�J2L%�Q
D�sS{]h�3M��9�] ���v�Ƙv�e���2�����3hn,C8���v,�TZ�,�B���%"	9գ^���k!ޏ�w)�x��zX�g9ݿ���M�ӥ�U+r�%�X�0�5ͮ�|���=�4�;�v�u�yG��X�g���;H�tv�%��
q�}��΋�]ղ2���Xwہ�����J�r���I�"M�
0�n&
#�J_W�_Ҽ��tt��i�q��!�c��8�H�:>��M�P����E����=������7.����� �|�c����#S���OC�����I��s�@��g�L�V}�V���W̅�l�����[C���L/�-y3�)98k5a��"Fb�[���3�GA��f|)�����YX2&�V
�R,��'��\�q���ۅzf��
��Q��s8�t���m�XQWmVM�Y�1�X��L�«pC��Y�Z~�ޗSz����@��¨�Ѫ�Ϭ��;����./՟q��p���BǪq�ņ��T_HTi����$�8������Շ�X�i�R��nJ�>��n�KO�]�Ѳ�,�$$�"����C����q��tt��)��g�%�����w��?x�ijT%�J�	�(2;�ţ��zX�gA���>3Wc�i�q�F�m�r):s�i�U�����z�tI{'Ai�H�m<qu�n
����;��6Ѣ=y�O���������s�x�����{��v[��Ϸ��ƛn$�(\lJ�13��+�"�W�v��GO3��^8T��'�t��^�T�r<��2A�W���Mz9W�ڳ�俬���sZt���W��k���J�2NL�?2SVȪZt�6�?"'n��>^غ/�t��P�k�����*������^֖~�e
>"���v�̍���iK����I$`�!p9�:'�#���JU�a� ��!�WeT�DF�V(�3DN���׃V]��3�E�am��>�[�?m�cn�,����J)k�Nm\���卵��h�X� ����������L�����[��q�}��f�����Y�k�ղ�bym��7���2l�+mu>��db�1;�,ݣ1���n��l8�9YPslY�+�yj�ԷuCqKUmUUB��.��km��hS����cm��	�w�_<v��a���J��p� [FЛ�v�$�~_�_���
����7�L�t�y"��俬�8��5���c`�e���(:Ֆ��^>�w�����r��\|`~�X!���t��}�y�/ ����|p^)gT�oF��Vp��Eqt(��(w{w����s�Il�&Y*q�[^�����UE�ΐ�̘���4�36�M2����TZN��$���&Z7B�V}e���M�x���5d2*V)���<�	���l��j�Vl5l6����VtR�v�=W�����#
�t���P#a$�=�8�i�s�:�v��<�<|�ӫ�:�!^��z�=<�8|{q."���Ԅ@IU�׈dXNj�l�ګ���8!�⛌ݮ#�9��h�F��D�,�T�Ud��c#��L���dJ�V�,�q氺�JF���a����W#�O��r>��EyշAU�,+Yxy��|�Z�H�i�����/�B��jz��EZ��^8!�ψ��n���|Fv�Z�(F�m��mޜ<�d�V�(rr����9���t�i��%RY�#	(a\l�͜��<�nl�,��C��r�4Ȕb�Y<-*�|�޽O�����8 \��j���\�����g\1I�*�q�;-�C9�,�"��Y��VIWu�5U*,X�-��]s�𾫳�:-;C��ּC>8)�,�iqV��z��p��{{��ETm;+(Y���G�kȩc6C>��p;dagO�v�T�"
�md6aW!8	T�صJ�YV�kXC>3/jd"ˊ�17���p����W��n��!��Q��]@j�&:�ʻ=>]�[�X�<[��guȯg�������NT����&s`��%�����:p��=ɫ��:��v|S�0�㮳Z��7E�X��ڭU�D��
�;,��^8t�w�=ɾ��ә��8͐�yp�����u���|��xJA��8ψi�\a�2���|z�*d#-6��tvt�du��{�<�^��z��q;F�v�[�:C�|�Mg�Y�:���z�/�i��Fj���E�:]��7D
�� j�����W�2r>��Hy2���^/�s�ʺ�l��b��g�Y��N��nH2�(9��&0t�޶W��9헒7]}������'-:I��]��c]�b�U

�8���#%ec8Y僤
�/���S!i�|����C�#��
D�
�#��Yn���y���-�C�yhɪϨ��p�Vj����~ޜ:-�����G��w$@�9辇M��26�j��N���|C�&��j�Ƿ\���ȑo*�<TVU$�jD�J�<h�cz�->_�V3���X9į"��ʙ�O���������,vKiU�]^8x�|"�Xڿ/��;-�D�|�aچ��,��uo��y�9�a��m䑷m���b�W�W�&]͵X�y��	�9�X�M*�\��DW3'�"�Я8��6M5���o�q�Y�Z8�fsG:�<�:�x6�v��
wc�͹^lh�v��۶�eؕ�7��N�m�`:�nУ���şE-�ѝv�d�v^G����x쨅��BUb��[�筝��#�E��fcI���ciI�v6a��V�`��VyV�����F��4��[x:���Pm0(�c�|Nlp\�K�=����ѵ҅������	�g6���{�{�n���^o~��_C�X�22�j��Nׂ0���M�������PB�R�H����l��3�g�Y¸v[����T�#-P��^�g�����e�6MZ��dV��rb`���l�Lj���{��#���4�9�9UH�X%#1LǽT��7�[-v��}��n�}|]ή��W�CR&܈�[��F�ڬ�^��s�ʺ�l��c3�g�Y�;�ⶾ���X�Fyt#�P>;�������-�v�vy��܄�9x1Iժ������-)�n1H��V-@��4��E׹13O`�L6B�-��5}�A�لC���F��U1�����w!�������C�x�]LgO�%����V$՜E�;�����@����W�?�?rz�ɿ?���:]2Z'�f��E�zI%2�a�̶7Fnչ�ʼ³���*��M�+Q�m �nc���������T�J���7X����$�) ful��n4C�q�zY�έl���s��]������D�%�[F�,hB�2<yT�j}:��r�}%;�]N��9u����	FԏԂG+�5�	����c4��;�n����+:���a)#�4ʁ��e��U�k��1�ԛ���:r�;쬽�x�(ד���E[�����LT����\�wF�]_J����͒�,3���
Ga&����^(�A�����fe+g)^;{���"��+;&��[	?��u�J�	w<��`�u/�]���:�hyV�;v*�h:� �F��_���l��{�u��zs����j�sY���.17��\_b����Oԅ��������:yL�_C�X�V}v���"U���.L���z��΅z0�*H8��7%�Ǿ3�{���8~�Q�gC�jt��Pצ�i��j�]j��9��HYI��H�ש��~]��!�ǡY/W����]��5�z��u��|p��ǯ��.RXյ����1\_'[S8���t�����t��k>�]��<����0�P���uUj�lJ�]��6���ku��l	���F�n�m��Q�V���<q�YGްU
�a�������f���~qo&7t��<(ur���R:��i���|>�Y�[I�Ņd]���tԘU������\�0C��B�^6���7�g�ku1m�H�~LR�Ww)�������w]����3�����3�}�s"Ϯ�r�Vި�L�p-�#����㇌�����|��1�W�D�n��a㧅ur�W�ٱ#��\�[q֚>������t��)_��.��bl��~<"�~��/Y��� �g�_�$nH��6ӍպB]�Bz��J����eZ��h�>��UK�gq���YC�9��3�!�SU�J�@�)FГRtJ�m��F�cYT�!e%��S�heh
��TA-V��j��� nݚ���X�h���#*�Y[B��J�����J�"�e�ToaS��@nS��8�ti��:Uv���ML��n�v^T�
�D�:�,�&�eN����-r�5.���t;=F�T�f��Ź�J�E��۱@jGf.
��bUc��$1�V�XSY�4�N��mV��6\�ٵiA hHc�[Q��]z��^�nv��[h̏%�V���� l�;u3i�]��nG�|W#���Vu��Ut�z��D�׵ǊI0y��m��M˛$�O�Z�'=j7�\p�T��i.��M�mbvk��ݶL���n6�V&���J�<p����"�\����z�vԔ��݆ðv�� �v՜�Iq����y��sv7��N��$f�m�N�y��\;�+&��d�Y5��vѢ967&��˙n@� Y�OFz�Ia:{lƽ�����HrlG.����U�k�to=Q��W�#��jv��1�ق:��ђGe�m���;i��#\&�v�V�<	��,e�/KJ'W&��a�ϛ[��7.�c�祰��\n���������8�v1�ٗ.R�=Ԇ�;K.9�+���d��G��nm���u;�me�yh3����lv�I��;��sқq�@��0�!�m���L��q��3��6��0뮐�ĭ��1r�7u]��(�=`&���2m����hw7mϰP뵪v;B�G���[;I�S��-�m<�δ�M�PSM68�v3�ڬa9�d��Yݕ�烔��i��*\GI�+�m@���W�D��6H<�<���ݻ{<B�Jd��7��Db��@Z�n� ���a��$���� �ѡ7`�̫UU*�UUTUUU]R��J�HL�L�L�,�ԫQ�U*��DD�6��@,)�+F*��^v���T`�z*j�U������J��T@UT+5UJ��t[ ��b�
�Wi�cc+mhY`J�mX�ƫS�fٻ6����{ `�֝�li9�ñ=�rV÷��ưc
̤[/��',��Sֽ�Ŭ�X��ck�g� v��!�&h;MA��\N�힓=��\�G�sG-۞�i��vNS�{s��2nyݳ����^�����aL�k�:v�k;-�2+.����y��Ӂ����1�����j�7P1@�<p�-SN�U�'E.���� �s����=�^�v�yl `��J��GXlvx:޵Ë���5��"�tE�H�)��~��Z�/���y�:d�pCV�_'[S8��seg|���5���@L���k܇�?�Nl����~vdŜ����ar���7�}�ۚ|p�z?pq��t�X�T�!V�_VVq����׹}�Mz����\	���S"?ZWB���*�#��%g)��g��N>�U�����x�q���W����:~�S��
���T��f�^z/��r��}����L�U{:a���*�r�_x�jU\?tY��L�	��,�l���6 ��뇔�z�+�÷��m�0�p�`���ت��"#�IH��C+�飡�����An�u����3Iu��l��D���1}�A��A�p���_G�qݾ&�se�5Z���ޭ�r"�e>��VB�2�_e�߽��y���{���z���:a���*��z��%_X�n�T����w�~}�8��O�>_N�y\S���N���҃4�5{M��'A�H-����5�KJ���|l���J�kW�n��5���j��>>������
���Z�� �𛌺���{;�6����<�1���B8,/���������óOo�L����;ƾg�Ƴ��X�p*�t��y2�I��Bx��I#�����Ź����b�ϰ���-���_X\�,���������u�����y�m�.r?���9�0�z,�x�Z��c�~���M lD|X�@�D��2��g��:,4��VӇ국��yf�Ƴ쥅���,���&PI6ܯQ��I�Y�X�|᪶~�L�W�`6y����6�����-�.I���V��]���G5cMv��$�Iū>�(��s[/*md%���b��D0�G�����wa�@a��k���^9��?qT��-�~)��a,��L��z���_5@x�����z@�M����+�����5%��We�����~���}�	��U���ۊ���W�Ȧ����d�̈��$��r�rȶ��?�UZ@V��%ݠ(��~��V���'�� N��R��Dп�Z*�<���8���^���C�f5x���M�fz`�s�oh���(��23&������l&�'h�Z��3�v�nݬ�O*�T�r��8�
p�(�z������2c#i6�T�+���>JY�^ :��:������� O:�p%ʇ�\��~W����d2+��`�r����M�km����F�%f�Uy��~9���P��!��P<�k dI&V5����ߔ�����%]c!�fL�Y�@i�fLd#�n����y��z"�7�GE���vS0H�24�ڟ��m�]�fByt�7I��<-��8�j8�m �b�*Y��@+(.��6)d؞ʮ�(2��fm�M��L=��޹^yG��8:r�ۮ���m�S�Y�3ӧ<ݬ�aҪ�����F�;zk�裤;!�l���/:4��8�Ll�rV���W���m�k
8��[=,;���m�l[�e�=hvz�mYܙK[1lV����WE#���=��.IQ�WeW[SSm�8�Z(��������S���rk���l�:�g�N�+�ɚ���5�.���3���ؗr�Ӷ�Y��@�����;��Ɔ[[c�fu�&weM�7��xyrI(��b��Ts\�<��3��˽U�{��_���i����REam��{�>q���ʨ����2���W,{�j�ZF��mqZ�&��)4�� �e��9��#�H�&2w���#�9�_��nM�k�/�I��q6�R)�w_nJY�u���M'on��Ws]λ�$[$�i����:��Vch�j��1��	9�IpP�0ca�20sQ�>�w#Y������{�6�2�uQ���^U<���D�M%	�'	;���fu_�z�tp��Y��{Uop�y8"%�BF(�E'��pk�^�ާ�Kqk����nʶu.�,�)MC��;Z_A6��No�������Vx;��>�D���GK,deL�ɫ�8+S�E�`�W~âAP���z���N�]�ONP�X:IT�*���ֹ5m��=�q;l�:R��h^M�.�M{h�s�j��"P��
��i碽y����|a�8d�g�|]ɷ�E��"�[�h��Cdk!�� &(h;�p�fL�d]�t���C�Yg��Szi��,��>��o؎�tM�UTl*���-ͱ�ag�1ײ?V���g�:��ǌ��)|�5J��w�ag�#��O�����i�7���|j9�XY�&�H�V_�H�Q7))�d��������znH���T8!���ÙU��#Ǯá*��rZ�4�a�^G7lJX�-���5�8�{M�A�Y��=��t8���%6�q�r��J�D8a��yY���vM�L�uw�.��Gߎ�T�ӥUB:����q����,�7&28�*Nq��J��Ӈ�8-��@�	�J%UU�氍"�mL�����0"���V}T���˫!���褲T,Zp����Lq��4�/��s��U���ϻe����ܺ�LK���J
H�e���cF���a{Z8ݹ����=�6�L��B�ܡj������Ilf|�[ۅ�yA��8\Ի5BV`&��m�،�!8aNa�}�Y�YΧ�No�����+��\�\"�2'n.�X7�x�އ������������?=��Z��\fGMN�c�V0R�t3�M��K�œ'�FX�I<�Osi�s�,��՚՜�}��Nֶ����L$AjB�Q�X�n���n��՗ѭgo&�.�<ゞd4�m��<��;C��lT���� )��A����ܦ6n�Y� .��A6�9 �ZJ�������vgHW&(�n�E��;`�M+�r[�����{z��:�n��7j,%�
�v���U���ڐ�s�,gkI����b��<N��� ]�;�vC\gDYhOL�����Z�s�;Nwb��<��F�`�S�t R��UnQ��-R���˰&0Q�s:֚��{t-v1rj�hJ�u�/i�[o��H����P�[����ͤ�qQ�:c4�ʼ&��/''����q��7�U+n�x�����w��r�a�3�E>6��՚>!tڛ��.�����Ƭ��"�����h�aO�>�\h�mUJ��~��VCG��>��}����S��2�	�Y�a㧜��kM"�K*���~-�f��g4��k9��h��1��Tn(���p金{�����oo�~�a���"��nh��:*�T��}UЫ��@�Xw/F�x�^|��c����<E�s�<���+��������h�p�2Jϑ�pi�x!��'˷�|i����^edmU�%m���a�z��E6s{ �G�"}ʸa�Mx�/��O��-�РlR�@�|S���zj�æE����i���g�'K�V�(|p������U+
���h�����s�o&���ѭ����k�(2�N4�E�ެ��c[y3�uyכI�<��u�}�����r�;<rdzF�R�ɤ8��5ǎ���v�gh�A� ��D<�2Yq8�##���Qt��A�#�C�c��g��1�<FG�?{���q��Nrж��7�C���_uY��:nL���溙�d3�1�V}t�!�ѷ�4&�v�-�իƝ2h喙�Α�|:��A��[��3t��(鳝��o+,�3�"��E ��H��6}-A��Ydi��J������[��~œWp�҈��n&D� ���|d�)�N�J�vS��ˮ����_}4�1�<���yn�]�mX�i۩5\c�{#k�<ع�4ȹB���)k�L���TP&
�w�5�}��F�e���ɑ����a�ȉ�2"e�a�Lأ��-�Lf꥕xM+P^	�kp�\�%���a�&$Փ���sm�s����՚����^��M�ɷȚl˭��H���Mǩ�x��j4��=�TY%�")&Ke����Y�ٴ����t��O*�ý:Nݶ��\"4J�H�A�Rٜ�7
uӁ.�0�ڷ<Z�y�9u���[\��`��r���G����]k��oU����:F�,B��z8`�kM�j]r�D�mn����Y٧�y�x�Jw�)��0Ɣy���Kq�ͼT�W;�c7J�/tk�a
"@Y��#�x5��3�=����v�fA�V;mhky�I8[.2#I��N�vӗի����w�{�o.�9�1��d�ؙIg*��Y`1��d��UV;�\�[��Y|.�`s��^�����r��+N^f�
\����{F��AY�ns���ͺG��{=n���M�3γ6�;�طd ���,G�'Gv]�����9��c:���[�V���ź��#P����5���;�����m����p-�{$�Q��mUAK����l+V���[MT�Jڻr�X/l:9���'�ʣS��;��X�؃�f�8�mkN�&H+3�=cQٍ�n7��'����U�3v�j}��=wǌ�}�5�/��eQI��!�<�ʿ���g��6�3����Ί�#J��Lg�kܯ Ԕ$t��B��Ы�9�ύ�s5V����Ɍ���wA�y�3�1�V}t�Vy����]'�ڋe�W�t��K�7�t�+�Up�枦3��0����c��Vp����P��e%"n�6}-A��^�#��
�o�bmY��d��g����:.�N2�I,���[jh���v��[O&�]cx�����y�L9R8!P�R)]M���P]�u���S�=Օ�{o���m;��w�Z�*���q��B�����z�<hn����ٺR92��$8���F �I�M�ǔ[Θ�Ы�F�9�r��>����{�WN3��d�i"
�Ί�#M�9&3�5�����Λ�5Z���������	(��n�J7i��w��t�gW��6?��ӹ.�l��pw*�5e����W�g�g��~�~U��V+�]����)�ɭ�3�(��.���n2m��)P!泍���Id����z*t��s�}�����\0�z�6ҽ6G>�_���Y��O.FAZ�ۀ�H��j�æE��e��X�&3�5ܦ��rE�/$׫����[�vĖ��F�v]񧁚��Y�3�n̋!i�eM��`�>#���Y"��+v����HآHeHJJ7_F��\ �3��Əm��Vt�W0����F������J�V�]�n�B7���1��6�M�K��{!ǪK��b�QH�%\�p�WcA�ۭ�X�a���gY}���5O7d{D��-�[=�P�������Ir����ٯ��2T�"�SR��D6Y�!h����TA5U`�uuY"�!rE�l�i�c3�XdagK��V9��diDX�a�>�7�>l��a!,o
���&��n����a�C���x\,�1~���>�6��~)b�mAuk"�"��8=��Y!���^.��Vx�#�Yv��N+4��dMEm�V���-�/Z)�}�Ud�Ȅq�2��#yg.���,�֠�Wjd.�%���$�Q&�A�7[��f�R����~�wdJ��['��T�+)��b,ʨG_?��+�W���w�Yt�.T�FڑYp�����H���t^<�x��7��l#���^�b�!a�ŃܷU��ɐ�o+�қ �>�i��AU%J�4�-��}Q�7�ӥ,�oIݕ�w���/o�{�a�?R)����H����v��M��e�s���u�&_3c?{{Ȩ�{��j����J)Qm���!��:�����Bg�k#"��psY��D��^&�-�wj��Z<���^u�nrO�r��Bl㦥6�B��̙Gn�R��F���y�A,�����*��we�V�sb"�&�1���7n��:���3ŗ[�sW���u�v4n�cF��;/����v÷Vu5�v_1��-�6�s�:��Ls�C���C����Ec���jVI��y��P�R_m͵��Jɑ�۫���m���l��Z��JJ��ө�"܀J�`9���)�[s��<O\]7���;���6q�-#��0K��j�"�v�fl����FRq^��6�Y�GY�)d���ύ��*��׽~��~��rDL�U��W��Ě�sY��!hk���l�~Cgǲe{!jE����S$�ح#�:[�]8*/u�k�؄#�`/���@g�o#"���Cy]��i��v"��$�35j���"x��2�3����!JE�j7(�l�"�nUc�H�qr�
���	�p��Gr�Z+�W��~#��V#[���2�~6�d^��VȽ�w����~5��'=iG&u*� �Y��b�8;K��l��u��ݬ�i�O14K�q�J�k�����ë�o�dC�Y��1��!7D��(�׵H�~�uxZx_^���;GTu��-XY���J;鐈E�{Jd#Hg��kfB.��N�nY�D��FņJ����l{�=�����/�{�0I���a�z������i�3Y���%$"F�i��w}��#)H��&v���!�&8�D?R%���U���ɖ�2�č�bh�
�Ї�B���W���%��D"�W=�2�3�fB.��e�Q%�J7uu`�Z
E�qp@�b�x�����h,� ��`u�B�a9�9��y{6�R��2�0䪒��u(�o<.�l�nTym�l��)5F��Th�T���D��!���y�N/b�'W�ȇH�#��G��rx�Q��e
Ux��s���~��b��S�8���2�]oT��C�3�ޜ�)e�dTdr�En�[��7�^�D6F�\�Y"�P��dʫG�Ƹf�F�t�b�"(]l]-R�6��`qn+�x���U�#<�I
���|z�z�B.ӊ��Ž�1��]�FB�P.�x���Y.2������-����܈�Dmրk.�b{7�-�Cڪܭ���"s=���S�<o�ɁŚ�.!�^L�L#<��yQ���R�J�+7y�D<r�B2Ԋ��yl��0���M���q�2�Ät[�zy��r�+��|-<~:��;-�qx�����Fy`�%{���"�����LR�$�Q��l'aQ���\9�+�x��s!��a�4)skîs���D𶕫���f���9�*o�/=���Ckb�Fڑ_��%=X!���&J��^(G=�t]@ұ���,\��h�u)[��&��dJ���/%eU�!�<�%� �U�J��]Ud8C�y1��B4��ĞV[�b�qeU�#|�9
��
������B��ʨ�%�|.W�;�Sw�:a��c���86��h��l't�dC���:�uTj��ڣh��qn���u�!��]o�Vz/���Fb�_��&y`��>#������L��7�w_����b�p��bb`ޥ��0�blV:-�qx\����ǅ����SQ#�T&���V�z,"=���F�_�1�`�L8B�q�q_�#�ۙ��/}�>1$��?��?1�Wlel���Iv�	fD�VTC���.uL�f�fyMZ�U�g8�ഓ��\DLu M*Ʃ�1I��GT��
ZS�U�z���]��"�+J�Z���;L�q�K��b�US��V��,�ڇK�ڍ
��Y��WmIEU\�S qi�<�y�Rg!��^��1ms*n�*���@�FT 3m;q�@� �l���z�l*��Yq&������� b��26��9�h֪��ěX����ڳ.`��2]�-v�)l����)�}wg�m���e4C�2�g[��h�Ov;E�UZ���Y���4��E�)�N9g��x9���Ú7I�h�!�\h��mn�'��K���q������΋��9��|�<���W&��������!sn��Ц�ܧP�9�96x@ݨ����.�����n��ɫl�m#^ɴe�Yc�G�7Bu���V�gEvy���6�rN�5c<��7<	�6z���jƔ�f��`6��N�;�kK��gc[�:����t�ѱ��S�iҵ�h��Ajސ症�mt�u'@�����-Z�HG�ցey���'j�A��";� rӺe� y4=�+#\�SGc	4'3�`��a9Q����7h�q�l�*�Wnf�{#f�ex�Ln�3�۲\���=Z�V��w2���9����Ce)ۛv��a�s:��}\��m�zQ�ݨ�޺0�w .���Z��m����s���� �v��l�姶yu�&+�`�/:��$��Cv��yE�6Ύͭ���r*hQ4��n��H��Y��2�m��ف1�\��5!ӑ�`�s���wNsS�U]��\�,��lԪ.��s�ƻv���SÈ��[*�܎��f��ԣ��8�����j�,`����S�����8ȼ��4pJT�T����Fc�$d���h�ZU��M��T�RҕT��UUV�*�UUUJ\Ŵ*�P�ʵ*�UJK�\�e�4��m��T�T��R�R�Q����lKUUUUUUU�����cSR�U*+u�햭2��
��FͳI�I����j@K�ek`W�
���)=n+����CVrQ��N�4�N^�5�N�R�h��%�����X��Ż=I,����/=��¼d}5�ΐ�7g�v��pێ�Νr�^�sOQ���y�@�R5u�'css�V���HFy�4�#�N�i\��M�ڱ��"�
��������Zm�u��3�+;3��Ԃ�.�U@�3� 4�d&�T�:pru�<�Kdq��N6�k�zh�|��vz���7�F@v*�^��KWTmХq�j��YS*,o��|~/|o���u\\C���FyW5�Y�D>9G�<o�����s���k�R6�kq��*����>!�SUd��B8�J��:-���:�!a��جt[�b���..Y�)��Ѻ��=]�����x���m�B6ӊ�SoVtÄ.��|<��{��0=���8n,p��5���Z �
���n˘Y������t�3ʣ^����C�n�HתѥVj�R�VMWY�R+�܀�Vl��ɒ�$W��\�W�lLN����i�������ڒG(��b�#&�՝u<����{v[�n1fL=T�O9���\�H:EF5j�Ȭ�W|����
qy�<x��U�,"��א��"�'f-��㇍t���N��$��b-��/b�x�s!�:-��VȆ��`qf���cד!��.ת��%@*Ȼ&�Ti^N^"p�����-�Nł0��bdY"�P�;&U\8D9緫ޅ��h�R�X9Gw�����͋5�E�6��-�a/��̞��;>�-��Z�i�c2&�N��F��=~��[�{c�ĺC��0CZ���}�,��$-eN ��R<ݶ����/j�#J�=��;�ѫcvlu�3�3�2	i#����ZE-�㇅�}��|�"+!;B(ȷ�r��CF|&E�-���3��(��кUU���톖B4�☓�9�E�6ͨ-�a6$�\���^�|Et�WF��!d[ʘ�]X!��d�������CDC�X$��!���V��R�UU]��-������}W�L�L#J���j�Ő�2/yn�/~z�S��^���8�Z�����U��^�Gqb�p�E91;|Md#L>=�^�\^#hŊن���P�k�IeZ�g7��0���>z/�4s��Y��[nNS>��.Ѧ�X���nH�ڿ�׵�}U��C�X��3{y�\
��oe��'�F��q�̑0d+�����T���f���Y[|�����\ު`0��0 �"[Wǧ7�'N���ݾ�d���˩��=��!��6I"	��ې=�*�����7"�ʲj8{{6��>2�I	%�#��9^�V�T^M��s]l�Q��ڥ�����hj.�d�RM� �B6�M0dWkq�0�]�%77D���Mу�Ϋ��q@�A�m��E�f�}iu��z;�<쭮is~zؼ�W}4�\���B���J�ի�
�`�n���D�6�,�j���Y�}5f�B3Sk֩����H��l���@�pF�e9[����+��!�$^�ԯ�Y�:˘#W�����{zi�s�o��ۭ�*��YAɼ��|n�V2/j��y-�!F�̊�5X���b�a�ʴ����K�ܒ�jKG74����;��{�<�S�[0�=�=�Y�}�6�![^��m�����y����WM���MR��e���8��+v�)J�Z�]l�a���:݆�v1v�Mf��w+��9-��"�]��!��I5v�c�al�ksxD��t=�퀑�\�s�}[s���&��&�nڋӟM�\m#d)�eŸ��o�U��=p34��v�v��-�����q�b0;-�=�n I{m��tu1uU[WUU�W:W`�[Q���&Iv��F�ڙݜ��w\�֎��*L��np�n	��\:��v^(�U�"�⚂��P�����m#TU^��6D���ʵ}��y�f�g|�1����gO��0q�T��1��%�-M�w����ܓ��<����ر���^Yp���g�[%dj�}���0���^)(����U���X��g�^}��(p�s5�
��ada�߹&��Ο�9�XʭV[(;mޙ�w����,��W�����������}�������_��!iUe��i���BLg?2�d��|j��N3�kڲh��!�ψVz�wF����X�Gh��6�M��+���c��nN1���01�.�{Kp��G�<��[I�^F��8�U��/q���:P�n=�_�y��K��L���\r�^[ N���*�곚��.n-�g��jxb�`�K6B��'��83��6~�]�
0�]QWlj��t���wۛ_z��<{Y���L�3����Ռ���Upl�uW#$A%�[kwW�:~�{�߼���q*���k��}��>�ӕ�]��}�=1Ũj8�[b-{�L���ɽk�x�ɷu����L\>�t��&r��/ܜ��ݻ��B���`�8�;.�0<�4�0��	(�U�\bie�	�T��dQ˽4�qߑ�)s�N���>�M��T3���<�Y�|ϋ�rhWAI"qG��PqWo,�S�_:x��bM�����J�����ߠU�agOw��c��W+�
�@���_z���jم���2�9��(�ɪ����W�����:h��uj�v9mn�[Y���h�>�zL�W�,�<�:n�ןOU��â����$OͲHʕ+I͋�x�2,damz�\;+4Y��d�qU��mī�#��U��Eb�U��thw[��m� �ӌE��e�%���F65{rN�	��� v�k��2�eM�iӇ���W�|�y��fFy`nz�=��n�k��+Ե~���nJ��n�x��-���U���F�p�:/ykt�����s���s��{��r�G����wƌ��N%.y}*�3V23j��a;0B�>"�Ug5z���~	�дj�
�,��w����}��>�ӕ�ŞW�F��ad{�s�Y辇��:�BP��$q�t��R�>��>6~6Bg$�k־ӂ?L����D�_г�����rH��B7$�˹Y�X�mv�]��Ӽ�WO:�XH���ꕫc��#��E-�^�����9��zp�7UI�S6/��eMX��M�bهd��?����Gn�vVɽkm}�l�L�=���xRϰ��q`�{UE�
�m�Y�p�U�V	��vnɺ��ؾ��9�Wx��M�b��`�6Bg���}��zd8D���`IE?@�be��AD�{�t���{Ϛ� �3���U"�9�s)iΊ����~���r���B�ڶ�x�n��Ex��ƙ�tSɉ��K!�L>=B)���f��x����.�]��;@����Uj�b�l�H�`G%Q�6	:5��m����P��GO,`9tH�[.��V��\���'���klG
��=I��\c9M�B����q�I����u�n^���;ݐ�L\6 cnGk�5흹�iM�KA[9��UXwbu���ak���%����05�z�$�\�҃n*�٪���Ⱥ�]J�յF��;$PuB_���%��g�d�X�en�@�<��&��@>���{m��6�۱��<�G#h�Z�6on�P���ߟ����X'�ު�D4�x��[u���"�*bmvY�0���s�4R��$#]]*�Q�Ax�rz�;�/*Nu~2d�^{=;�߽���^lp��&Զ��B��d�{���.z�T������*f9O&��~sW������@�m��;��Wx$[��#EL6�0���$�Vz!���]�#5H��Ã{0���!>��k�TԪY#N���׌�����淖�3B����灵����'~7ҝ��Znv�]	]q15iTj��n���]d\����KtPu<�Q�Zr7I�p�	mU�Kd�E���Z�g��������-��Q��:Dbd����1���3�r�删�26'����!��5`mn�hx����0������CO�=oe��#qH���JH��RX�H;iTr��4O�{���׈���2"E���U��0����x��NK�ñ�:��8��ɛ���4l��V)ynH�XH�>"عd��G��GQVj�_P6HTmQ4�"E����5���B)����W��/�#<�E=w��O�>7�g�|�4*ԴR�V�j��¯�t�KW��7�f���v�-�g�5�����Z�
䤶[������W��f�0����d�����)�d6D�yl'4��<x�;���q�A��B�%��?��.?'�!��Uڤ͋��x�����޻��o�Xnx��N��܅v�l��������<�>>�԰m�5\}a��fbI���G��ڿ������[��O��t'�$y��N�m������]��y��\��"0��\�5<�㓞����环~n+$�U#Ad?igŇ{a�����W�<gO�gb�^?C�deg��[�㔒��
V.�X	�z��Ƹ�z&eN���5Ƨc��U��f��W@�˕��cj��>��M�D6a���6�?qu�L�͵�:�k�K>.�S�!�R-?8A�3j�(%f��c!���e�u�!�C��U�}E����ڙ�C��7-�<�#���JIF�jvأ���;��2���O�
�a���Eu��g�}0Ɏ!�!��߲r��ˍڭU�ٸ����E�C�����j�G^T���O��i�����{_|��GX6Մ�"-�!�N!�m\�?i�[�X�D<m�ʵ�Qmn��L�!��2bB��]�v�9���<�`N��f7X�]�7ZYƳv��˫���B#�I�	��5x�� ��ڞ��ߕ�&�a�><1�khx���xΟ��t'hҤeE&���8�����ke��I�z�C��~�J�U�2<]yS?x�+��#�h�E�eVʦ���O�`I��ha�f����ֆ��m~�^�;׵�}��Z���j,�w,�t��fݶ�P�4�?<g�o��B����ã���k���OY��-��"��]طu=jLsώ0vU6�7�j�}^���w����-%��
ے� 73rGY��keH�s�\(���
���.8����'j�يU��=��Jk�c�uk�C&���C�ϵ�8I�/]a��v0�vɹ�۔���9vm��7f�cn��=���
H���dm�q:�����m�m��퇧�1+�aT�#Z��Yx��;�r�L�FȔ�e�� �(��f_H*ު��4�?u 9mF3;<$<�HT�=j7%����\pi;=�����pv�k�����8��+������*���f~5��C���~���W��hsqVkZC<^E�V�R�F�VYV�;�5�Ӌ���p���W�v��~g�V��!gņ/|U,,��
�JY���|������3�;ƴ�:W՟Y�t���8!��>^�\��n��X����p�f)��a��\]it��9}�8¹B>w������-��Q�+e�νN76m�g�x�S�[/:Y��6����/{�3��Y�8��A$j�ȆUԑ�C���ӗ�����p<�Ó�=���h6�8h�c i���p��E�����8�\���e�?Y�q�դqһ	�Y��z���xu���d�VɫƝ>|>�M-�"��1N>���H���u����v:'�1�'�A�PR�c!���ܬ~XC<rj�k>��iF¿���><馚�(��1���_���+���|���|t�����εD<�z���?i�����f�I5
L;1�j�[w)�������N����.#Lw�l��ϸ�5y�i���BbTN3��!oo[	��"#��=�����J�"�ɸ,�:�0��ێ%�Iar�5kjFK��]��2�}��o:�L�=[w�a�w	�^t��p�Ti�ɶ���#w������oL�H�.|D<|n����H^x3��5��}!�ؘ�eC��>�𯞻�x�&�U�,����qc�+g�0��� �J���I���"Μ;A���t��W��hsr�Z��|~�Q�$7O|�i&�m$AqCn>��C�2���ݤ4>+;-��G)aŴW[�tnɒrƎ����;�o<l��v;����#2�fM�ŸS�.����&G�ٵ�r��o׺W.��w/[�;��bA���L[kiw�sͺ^�o��[8�MY�f����f�G�f���i�TFbI�+��V�}ڥg�x�|"v����	��?q�C������׼ʴB�"P9��j�����m�>��䯕z4�N��[�����g��Eq��"t�-{����:�|~���5y�i��T�QuA��Y��<Ǔ����\�$�V]-�Nn���y��)>��=:�v�?W�ʟ4�.�
�g�o%���R[y���?�>[���ҍ���C�����X�F�)��?3g{|��H�QJ늢��E�����������Ǧ�>���W+#N�ܧ���u���c-���u[&�x���|�JkH��LSO�Ì�tu�YӇ_�P�
���}�p2M���X�t���7)�ߦMYw+Wt'e���t�Mak"K�e�.FWi��3䦑�Ӈ:���M 3��u�#��xB�K���gU�U:� [���˘��eH��Vr+��v`�ifU,�7e���Bh6�[Sv�i�WZ�$u�Ȼ�>�Ě���Jv�vۃ��^M�0��=J��ӑ�]kv��묣�͗��t����b����pf�Vׯ[F�j��9N�w�2�ۭ�J�n�b�c�7Wm�!Θd8wjŢayؖ[`z�]�F�eL�[�]i�Rj��5uF�M���Uѳ�A`+��(�^���ܻ�׷k�
���;H�Z}-h��v���e$T��Ll7.�^�-�I����oB xS��K����:=��g����5zX�����P-��48GI�q3w�^�#N��c��Ϸ��_������<����K`*�ޏ_���L�b�J�D<D�v<Q^XC���	A���`�y��h�j��<�/���N����������K���e({a]����"P��8o8�<Am�8�\��O����w���Ӧ���+�t�O~�n&�-$�aiѤ��ю����sE��o;��w����g�w@S�m�� 	&d�m�k�u1�� t휥�S��aщy�"<�6G���-ނ,Dnu���w~��Zv�{� ���k^}����2����q�i{�G�ci��fz�0��;�%i���+T#��4���η�OξgH������>��Z�1�X!���l�/��׉~!��|��^>�x���t%����G�aR)�xvޑ�c^}G�����E����ч�n2[+�݈;zs����V�)(`^ې�;q��ˣpⴌ�:�r� �e��G��O��~�e�7��"ΐt����p�֨�q���"�䛀��$G%f&}�}5U�D$��ɺ��#6�ZE�����L�/��,��	"�dR'�
�?WTF�D,�eK��2�`��nQV�{��?���d�+�������,#�>SO���gIZE�8t5�~����)ޞ	�;`9[l��J��?Y�[��Y�ɹ�Ϭ�I�t�X>6x��Jȅ_k�$MD�p �uL�{V��Mv���(8�I�N��ñ���A�R�ccaG ;.4
K��[�3�4Ĵo����;�#��<)�~8~��MTF4�R�aI�RdF"B7�׬�K�ał,������q�����0��it�S~��d��PL9"(����JjȔ.f����f��3���[Y�9Js;R�3����T�E/(��[�Ro���i����ϊN�{�F>3-��G�a˾8~��&h � �,��_���r7�{l~\�9.:Vd�f;Y���'�H�P⧝vL�(]g�x��ڸ/�^2덭nWavc���xŎ�MYF���{�ws�G_&xoD3���ܝ\�9�|�i�d�Hۊ�q9n��:a���m/��/:�٦M�Y�Y��+�Q�E٧�!;9+������S��g��xkY��8[�T8!���R��C�||���i#��4E�7�?3e������JfzS����׏s�{y�h�28DR4Jr<��T絸Cܗ�
ڛ�a/��Z�{��~g z_*U��q�Em�,�������R�*��)(�e	�(б��P ��%-�q�J�WHOU:fP��dx&�IP�j���I5�a���JJ˜��'����������A�ژ��6��(D�u@T]-�y]!��.�X%`��ʴ��y%�UV���rӮ�v��� I�Ļ���5�sp����U�]Z�&�vbe.�aH�͢��Ig�<��;���s�c[Zz�Okk���.vɢc��HZZv[E�c'j��21��1��l�22nL��*�āe~�m���.7BkFG�_,�4MnvB\�jn�Ǭ�a��<�]��bɶ�\�:��rźꤷ��y�L�q�k��#e�ѭw�ܒl��ɢb0cq��1nZ�7;\��ݭ
n[�n�B+S2��Jؕ��rJ��Uds����X�+s����S��5��=�Z��2�����7n�{v��ӖV�N�&���A�n�y[l�@�����=&��m�й=��Cvw,� {�XULh�z6�Hs��P�<7n6�P�����:���¡�ѧ� �quF4G��lR��;a��AϷ=���.H���؞]�����-�n�R�냋��3cn��٣ U�=E�q�y[$��39��Σpn��\Լ����@��ݫZ'Z��'Y�q\�[��x�ۊ�1�ۭ��q�VݎKOn.9SS�z��zy����<Q��#���
��q�����l�l��쥑m'�t&΍��C�J-؞+n"slq��g�� %^�1z�'0�[�cb�;rb�B��l���瞥{<��8s2$	�9�R�:l��F�~��v�1� �p�G���`ե�	��F1�Ԗtc�����ԓG[;�p�d�U;���1���.�<a-����U�0;��U*�UU����X6��d���$�R�+ggV;U���]�P*����Uꪪ��
V���m�;�I-P �U6����UH:��-���,���Z�%V�@5UU[M���U��������iV���Z�e����	��D�ԱZ1��j�N�)ͩ*2R�AE)5�E�{mP˪i� ���h1;O''h\�ey�2��L��ػn�v�m�n��{mъ����c�H5`@���`�Hi�n7����j��W��6=%��\��չuH�U����������Jw[�t�ո2���<GJb�9eȀ��i��xnN�`��u���Jq��:jBe��Ĥv�-�WU\�����uC�Vڗ3<�㝎Cn ��]����pD����`\v�Z.ƭ�+#�lm�ՙ����:��ڠ�����,�j�>��[@������O���O����~��Fݲ�G�������e�Ư��p��spC�����O�~��Z�D:�j��ne���O�j�V}g���K�Ζ~�-�8|F�S�w�ޙҟeGp�
@������E:f[��<p�e�?Y�������׹O�=ޙ�je��y�V�C���RU�G��1�V��l��:�#>�T�l�!�%9hի@�]X�̹����-ngm&NI��#�^� *�����l�:�<�΢��Y�}�~�C������em��x�Gj���g��W���*N��ѕ��$�T��q���\��Di��(�#E��r�>��羱�Z��H�Y]q�-g�~�ĸ�B8��T��H�$�|~��=]�u��/<ǝLb���6�z��pAB����#�r2��?tz{h��}��mյ�q6�����E��q��A9"���;�E>.���C����9e��,�2�#hl/� �7Wm�[��g��籢����]��㲄v�A�1|#��{�~#��*e��8KT��y�#�h���"�M6�E�㡤Q�SՐ�A=�$y9
�~�|딈�e�M�<ЎU�i�.3�C8��8�E:JLB#�f@�9��.5*�`����uWuS���ApF���#��Ȅq�%�H���a��D���8�M�}��piC,0����,Y���ϑ#�9kR�-�ٙ\����c-F�l�iP+:��7.�;dnHۦ�]	�f�
���NJ��_UB0�0��0(�}\��g����"4�!�)YP��B�mՐ^���U8a��� �#��c?q	p.e�x�EH����$٨n�ݷ�GqP�5�N����Ǹxpy����4L���\󻾒M��rs���wl�ж�/��VZ-��NB�DU��d��x4������+�~����U���D+�+��;[n�o<�\�nV�rj2�y�2��N�9q��ӅB�S���#x���Ó�L4Fw~' �!���`�GЇ��+��e����TQU���W��=診
�*������cvx�w�g� �^�v�#v��@���Pr�3�et�����h���Oo&��M�Q:mW��"�г�����W��������i��*�u/�$6 �lǗ�|�[g��F��gQ��A(�$��U$|��c�iUuNӞ`�t�g[/j�Mps1�F���k�I�O5�ݜ�����9�N��a���f�a�;g����nӴ�;����0dͻOk�8)�t789�%�Y67k:��v�i48�#��lg�m�����ۄ�E�vN-rZ�hRm8ҹ��O6�:yYٹT�$'!���Q��q�������=��uK�ӅP�]�v�	T'�Hƥ�jڪ_�}�w�K�a�cp�mt�]qbNI��nh��]���� -�\���)��E�٪t����[�h��v�{�y�1�~<�	FڝQt��A�cukK�RJ������M�W&<.��wk��*f�0�m��t����Y!Q��J�j�t�1ūM�vئXm��Ad3�~�.�\����Z��(��X�,J�^Y�G��1�!��Q�OV
!��	���Ȣ�2��ڲ��.X���ơr��!�|.������Z/�;�k�E�gS̲�4��	p��c����p\JFE�v0��$��uu���Ʈ�y�7n\��m�B �����Z7"��+��G���zw�=*����a����X�ٶh���!Z/���O��S#v�";*ދ������"0��I���)�T��6D�N	�h`dYg�Ӕ|M��4iX7wJ��#H�5Kg#5W��l�!�<��dm�t�2\�"0�����ӱ5imt�!7�E��{�ޘCkJl/U�Fp���madi(}�zC����}���"���S��y�!�M8��L��pv��t��$�t�F�Q=Y�"ӕl�F�0���DA�����Ss�%�v'L���.�.���f�1�3փ�yz������Ȣό{,H��4��\8Y���da�l^��F�gJ�O�u&ʤv�qY,E��?ӭz��d3|򕳄6��d��20���c�>��_ٍ��W]��oJt\(rmc"�g��5c#K>1³ل3����M4F�Ft�A�#���,H�����6C8l12`d"ό{,q�������GH����F~��KJ�22I��ue]�dQdRd��D7ޘe����ɐ�
{�k~�9��8�B3D����s�b�%n-���X�C��C˔��g�G�OU��E��d07 �j߯߾�C���C�es���ee�y9�{1��q��q�R���R���}�7�׳�'�?Kq���i��V�)�3�TM�6��-�
lM;�:Kj�>"���|h�#ަ�#M�O6�xLA#	R2Xq�E6P��`��D@�h�4x�6:=�dY��3��Y�}~�n��iYUE%�/:h����aFE��X͐��"�>3��:-��{���c�В��k��M���U+�1�&*����q`���8*�aG���Uf#kkrZ����z�a��9-��q/Ռ�,�a��dC��1�L�dx��4%ZH��ȣuK!�¸=�024����8y��`��[4Ym����0�x�/e��Aƃ$8L)#�"���~ӕD|l�|B���A��T	N��ȇ�J�]:~>�W�O�e���Bɫ�=�C��\8Y|+�CHgNoՌ�,�/i�M��N������8[)m$B6�qdqf�54�h��k�qx�]�ۃL:Ep�8��Y�8�4��g�B��,�ʲ��+�-���'qr-�2C� ��
!���=��غ�ny;&�)�&۵���v�T!ù�Z`P�j��%�E�M'���պ�n"nXی�ol%�E66��+�gX6�@�;sVs����h�2�Y��}�&�;�!�ۧ-��7'E<�q��l2�Q�0���[�n�]�++@ ��7UTTh�XL�T�5uJ�K]-�d����:Su˷m=�"9�-���:���۴U���9��:]�
xgʀ�����!�;���i���n�i��=��"0����d;h24� S�!�:-+ �Pժ�D��H�[d��S����U��2��R����^�ߐ������E��r���:�&�Mܭ��v�ƞ<E��fCv�#�9�+g�ZSh��"�:��0g*=� ����!VP6,]f�#�X������+�XȼL��!���1��;�����R"�\+,�_y��|�*�Ȳό�,tVe��p�2����Y��B��e�!�y 2DS�5r���=�=)���)����k ��i ����9ӴVgZ�f�;���޽.7A�Oqg�����2/Y5�����;���*�HR�f�"�F�ٺ��kH�l����rm?L��K�SX��sg��H�*�.Я�ش�*�es�%�:�t�]�Q����&�[�u�
�����6��{&͚*z�[Y}c��\�:hH��g;��z��(�K���'&�����-��]�bG��{6����Ak��g�T��G[�=�Q��囅wX	Ϥx�z�%�F�g�U��%F�Q+rF�t��/ア��o��<\~¹���G4$&�*�ȳ�K���i���F=���uWD2��-��j�4Uiܭ"DS���W�0�"���q.T%V�݄��t���*�#y�>u(
8Aã��o�}���Z�,! �G�+��g��.���#��rH"1��. �g��y�"��q�g2S�����dR�gH�˾i�DBP([���|���˄q���o�8U�8��ƱN�}��.����6��m�d�G��Gf���G��� j��=N��%I���lX�9E����@��+�&��_�z(!��ͮ�J� ���E�;��f'��ء�H���q���y9|<k��y�U.4c+�4Bq9���8`Sk8��� RkB4m]��@c��4����� =0��C��P�_{�z-���b���XEkE�E��>8/}�k�����h����9^a�N��Yd���B�!6"�@�qgH�T;��X|,������3<�V�����c4~Ф���/Ovqɐ��Ѵ�ۚ�`�gn+=���oHx-�Nʶ�n�#j��������=�N3"χ*G0y�,�����dJO����4 U|I�º��m���&|p_�_�o|1��M4EⲶp���L9�|M�`��)��cV�|�Q{��J|/�X:OVx�4�\R�qk�ڎ��,��y�a�mUmV�B[�9^.�@g�!�<֜d�JY��Ks�����xa�%-�N6_ �iBQp��v���,d�de�;k-�� �:D��L���ɿ%4���>G)\�Fp�Y�\�/-=j��A�U4��8\.j�M#u�8F�-���������Xvm�U�Rx�P�v�W����g��g63�'�^�`�}I��4<�r^�ѽ�9��v$T��b���zP	��L��)d#QIO�5֑7&�|�n��+�!8��s&�=� ��3ZZ���kzl��ٮi�4�7C��Ю�8�K05UmUAd+��W��iw(�Pq�qy]�����M�3y{i�wT]���;jT�W��Nwr��]��A�AmƊ8�F�����H>͌�?J�|��@@���Α��o���>^u��ܭ��8�w_W�!����Y.�����kW�A������c2*χ��}�I֗�����Gj��8�L5_t�K��������q��uЙ8���j��J�(!f��%ZWi;���Mο"y�v.���l����zo�<_��;�Y�P2��G#�~�Ƶ6&�`Y�=B9�֯��=Y����|�����O�C�v��M#��:�ӻt�6��ͧ���jS=�Rpܐ��f]�\��qѴ]��߾��p4�ÄU.�^�^���i��oC�ԙӂ��|�jV7j�*��.��M�)���VV�U�W��p=<��V^� Czqg�k>=�:Ab�p*��=��s�R���㶧	�0,�x�1���0��!���U"J�EY��-�`l�q:��g���gb ������e����ƹףX].�(�'�ܭ�;Bj�I�3�v���5���ߏ�Uî�t6P������Sv��� ղ� 8��Ν�8ۯ+��u�#���]���c5.�X�hZ�X��c4~�V:H2r6�Y��+^5��;S>�?r�3Z����K���![^ES�o�կ}&����Q��\1;g׊A�޴:k�G	�-�D�"[76�����{��(��t&3X��~�U��5�62�^���ON�6�b�6��%����f��f�۪ǣ���x�s6���8���Onx��O��lr	����rWI.��*{����3�j/[�J4��c����zp���̦MB�ٻj�e�mٱ���n۶��:�R�H��mp<�\k����09�<s���j���@Cf�L�>�AZ��s>��?;4����N������V�QUe����T4q�]r�!�_�v��M�s��mY� %�A�� o�+6lUUɰq�����.8���W��幧u�sK%�Dn�D�9������.�WT���%Eȳ��Y)� �Ѕ2�l)	�5��>��U��˳�t�ܡ9�~��9U�ٵJ�RHS�^n�s��X9 ��U��y��Unz!Krt�	em�٭&u�#t߅5��{�I�q��e�E9Q�P��*��p��l��4.�Ut����@q�o-�Uy_8^ʗq(�����b��Wh_*�x�2���E��U�di�&�桨��������LlTP�]y(R�9!��Y��O?�c�(��Y4�S0�l��f��kP�4��T�������1��I+��BYc��S����\�h2N����O����3�)��ދk�8��?^�����)"�;G�5[i6WOeb�ZE����vn�>Kf�R���¼"የݴ��-i�F��!�]����9I�2']`�@Av���=h3Fc����-��udӴd�n�ǍY�3B\.���̫��9���6n���u�E���w��K���ܻ(.���#��d6����Zz�
��:Cu�5�r[glT����  ��WX���*Ձ'�rt�&r��u4����u�TX�)wWV�=��n�6�Q�a�<r���K4�ê�n�k7�ח�~�n�dx�2�Äz(T��7����$�c��ZD��9��!V.�ѡ��d{��oH�3�����E�f��z��p��(q�f�?a�ļ�F�������U�c6G5��`�QgǪK�d2N���i�]|F�OF����vi-��S��/q�x�O|.L�i��8�Q�p�q��:�C��;��8J�KWc��k������f��#M�&%p�C>=OjVB,ȼS+�DC��"�$�I�� (U6�\��4���p���cq.�͔�//qۮP��WU�T��Eٱ���"�$^"��%+���(4M�!��:yܰ��d2�����~�H���6���"��p]8wi�]��?�\r���>#��L�Y��.�p��_�����JƜ��K��8>���"di p\4alA1+���޺�J��~�n+��C�"a8~��}�p�إ���?q�0J��p�s�3eVE�|z��bqD�.�v���`��)k�)�Q������ZfC��FE�[4�e���N&H�N�~y�o1�D]p	VuЬm����@�fx�|�k�i�M�̣�m�Y���,+�qƕ*Bҫ���甘=d C�H��qȸ��q�͖F���J��~�Ü'�R�)-�[m��Oy�����5<l������P�Zq�!���=���|[�)#Zj� ��*B�`�^�x��yS6Y�l�o�� �Y�^��Ny{�R�M>�{=9E7�V�nL�n]'m�Nz�ܚИ}��bJ�d�Z�TMW��.��O&�Ų�4��^�nϢ��/@�I)�����=����%@`Bdj�(B�R��Rh�m�J�`n�����6ɺys�K��gge)�ܒE"��Ֆ�������w[,��S6Y�E�o�H�VB+�,+�ľ��8�*�4Fǔ&H��n�w��j�)ׂ������^���g9�G�Ʃ�-�j���Y�Jل璥�^�qN��J'�Ͼ�y��;��.V�<��+rS�������@��Ӗ[����>0���0�6@�����dJDٻ�Vj��
�Y�R{jLڧ��BI�[����'yd C��D�"�J�(U���;	���f[a;s�3��=���{1fшv|�̭����la�t3�����&|~�Aˆ�#b�!ҭ�@���dU�׊狮�,�����V(��n�f����(�'�M�E�_Ƈ�+!��X�ae���4͞"�;�أm2/�m�oM�����i�9$ՀQgH�����t���˰iP�
�J%]�-U�8�)��9��X��E��`��a�O�/��\t�w� 8V�d���8��S������,��L+�\p]�g�:]s�޺/���$�%�/��$�$�%�t�$�%�/�%�,IbI�$�$�%��bKX��d�%�,I�1$�%�/�KX�ė�RĖ$�%��ĒĖ$��$�%�/�KX�ė�KX�y�%�,Iq%�,IbK�RĖ$�%��bKX��T�%�,I�X�Ė$��,IbK_�,IbK_�Ė < ���e5�x� x���?���}���������� �ܡEAT���<����w+�3�A�;v��+{E��{\4ӓ&�l�p��Z2h�����@���    昘�0�   L#���Lj�J���0 2`F *���UT�	�      "��U U2d4 ��ѣF ��CH������#LM!�A@�a4��MLM�ɠh�'�8c("�O�>�P���&�����E���dY_��d
���"H�"E@�*(ʁ��Aj(��x������
�����f�EE�P��,��\6�섖��;�kZģ���{;��0�T�*D�9ᓦ�:��2�M��i�P5������,�Ĝ��rR�M]˖�T �l�'Ʀ��[�[���A�{ �!��UƢ�@�I�(e��_'qv� ���OF9�/5�Ǳ�pz��i0�ć!�a��gkw����Z�|Ah��(�q֛�)]1��,�CNI(1��L@��m�7L��r)PC)�Be2�� M��PB�
"
���6��m���h�Ua�d�'��Ij(�B�[J�
�����tȂ��V��B,t��NJ�"m��-�ⴀO�8�)�+��C���1�v����f�֑m��LbI�I�)!�@���H[�姩76'�P(��F�R��D�m��Pv� \m	@��մ�Pe�4�B�� *BB�0B�#�ڀ!n7l��qM�����l`� BM��H�$q����F҅;-��z!av0�l���n�X�I� ���%��^��i�A10��MM��E2�"4�X�p�A10H�����z���T*1�&�"�P�A@��CBm��!LT"���m1�6�c�kRP�p���*hH�um;��	�@&�X��U%�U�#���O4}PXBŋ �DD�5�"-����G1��hJ,jm��_G��V�\Kx��m����S4���h�B��UU),����� hZ�r��@���ل�YZ�"h$�j��j����UUPR-���b�jꪪ��*�7Yʋ��Z�����Pq�U��5m��*�Z��R�Vm�Y�=� ��[6&*�"�*��	]6-P��L�)T�uR�m��gӢ1���`V\�pmT$�9`���P���WnE�8�uij��SlH�Ȼ2�!uڦ.�0�.�tc#,@#�T���c�իٶժ�����0���`'�57lI	�e�A�:�����i9&�MŪ�8��CA��8�c����٭m�$�2ȗ�ΰgtFD�4�������h�P��<�Lm�w�1�Q�N�����l�ݲ��A�h2ੲ�IÞ ������DV��@t���n��雝��Ies5�����97n��m��u���]��T:$�o:�֮���"E\��Q��ݭ���ޱ��̫l�kf�se6^Y��c��:���A"t��ܩ�
�Y�z���C۰Iy��BZۊ���}=����.iUA^�5��^V��ql��G�/���h 6訣 $��Ѳ��M�����m~+���pZꪪ�6��0԰R�� UK�l�j���ZW�WI V��jx�/;[e��۶�m\�̦]:�a�'g�:����ɕm������|�aWA���:�ZH��śq�oo;w��y��^wt{�Ͻ ô�䋀v3���e3��snt'����H��/��w�������W�s�rdp��x��|ˏ/XO��<^l�5M�����Y�K����r�8��|���3��Zz�?��>'��|F��)�M'Ji����J�!r����3�N�Skq-��u�q\�e�ɝJ��RD\Gga%BH�\d{|4ݯ�/3�5Sz����%p��[�v�iE��%#5i^�i=]~Q�m�p�c�7,��짋s��_��oG"�ecJ� w5�P�dԢ%�҉ns�����m|G��A�I�Lm��q<YJ�0��axi'�#!�|N�8�.�HB���z^��4d��t�v6���9�xSv���i�dQ؂��׳�ء��/+�(bD*E�S�R��+8��[~�}tׅ�}pwX�X�e��E�NΞ/]���>�On���f���ǾC+qƩ���D�I6�%��͑s��l��G����+X-W�%�� ���`�D**�Z�LVu�U䨈q��UoAP�5�K�6�� R�!QU��*�7�UX���/|
�;��2(���r�8���I�U/ED�#PA�5� �DB�U���\�p�g�l���A�Q*������wO��'�A�ԣ�Q���#�O�f�	%)��Њ�Km���~��oZ���p Z���V؛�@���1G��ޤN���H�U#��:H$N�vB���bl脄����>)�_ڼ�/�i{��T�)��z%R"q!����
6�"\�k��|��N>$�����M/)�Bu-����F'"zN��@H�[d�	l�=�'伐$k[Ll��$w��D�o��V��_�C���6�;+�J�h=mz�]oM�3���}�]�G|������B��$�*�Z���U���mq���*��MUҭmJj�8����M2�9q��e�K���ZA�3q3D�����Po١AyId��k��Vl�-l�g�ܝ0m����)8�����;ׯ���״��Jl�k��3����i�c������j��{�g���7�h����w��y'�m�0�wz�[@�C߫�w�gw=��a7�n(��=�W�j�T)&&SE��,�n�+�PPP]AB�����bel���rՋBW���J�X��pLI11WUr�EH Z+
PS}��c��A�[]�B������&&*蠠��hZ*�o�.��yw�����H"b{䉩b@��r\��Ǣ���_��{}|o�P	*�M��F���PAՓjqָܕji|��|�%���'䁥
��d�ɡhI11WE�Wt�V�anHF�$���beB�;��Ix�m� U��)xT<�V$�����gb�^P�B����nA$$��G�m�GmݭR���
��(-�&*AUɾ]h�*�+�S^x�9�E��VB�Rݔ���SB��ȫ�eD�����"��T6�TI�%A$qxX�����H8�D�%@5�|b\��A=P*@��LP��ȴ*@��.u�a$$¢Z%Lf�� ��y�����T�J��d&6�EeJ�,1�k1���:�Ys�q}���V���qX��fˤ�:޵�5b�:��P���6��]6�q�-����v����].!�]��ꭵ��x��h���u���v�� �nrDZԿ���4���ҠU��*��R�*��&Gw#�
�魗H�x��t. cJD���K��v�Ȼ[��jl.��:U �+J�Qu�鵬;E�(Vu��Uҕx�����r;�ܒ1�vp��]�|���*�[ۼ��-A�}�q���#��C0m������S�$��$��8���h�}v����Z	�1�����k�X�p���$�$5�j�z������q�Ž�c������F�p3;Q��?̿61GL��6��ru�P�h.a��}�~L�/N;h;���,�������<�ދ̡�	z\rI=�5n<b��}��E�?_0���5p�"�߁���y�5 ���sz9���ݪ�����*��)I$����J�̕r��Rv�U��t�T�J9Y�WRPu[c\�.WR��&�Ɲ�L(�	
���L���Ki���b�*���˔����mûW��Qmq���g�'��l{�Wp,#�sv��Ub�	=��C��V�d.��o��+�o1޸�vE:�
����9��-��e�8�h�Y�qr�o��R~޸����p����:�%�ݝ����봟�9-\�-۟�h����t�<~��4ZNE������n�v�nSv���݋��.�v�-�	M�����}����Z����j�+qX[�E��B�o�'@�=���^dy-�.��%�V���<B���#���?5@MUD\%7�~<E8F��!������q���И܎��-\�u�&�Y��qui��/w�����o�w�gs8@8ݯI=�I�d���"����z%�a�5����lp��2Ga;'M�y�f�Ix3�%�-k>��+�c_G�ϓ�g��e�b}B�k��]����2Y�x!ǳ���� 1�Ĝ�{v��M'����4)'�(Uv�����]f淇�{�"�}���i�K�3H��7:i���"-l�7y��~�	���3��M�1~%��<rפ�-�)��-|x��4��/�qdk��-�0�����ӧ�dg�z�B!��<aW�:k�x�~�q��̖aŽ$���R��&�Q�(�����)��.Ƭ�5fo%CF���=��z'��_��DK���	���;;���T�����j�m�A�æ��çFh�szXg2V�>hɍX�փG��g}�g�7k�O�h��<N�����F�p�8h�nd�<�[!��J���|�o�o�HPS1��Ԡ�+*�ƴ� Q�)T�H+��@��A f���v,k�����"ێK^�'mGh»$!���ˍO�3�6��� q����Kq���kVo�ׯ[`�vv��U���93��(��	�,N�XZj��6zOg�v���حw�н��7{��<^�ݝ��0����r=�xu��b�}��𱟒�:bS���N������k��/���2_e��>�mڷ=����|��Z�mF�b˳��n��0#b8(Bd�R-�&,{�p��E�� �4`���F�b}݉���G�Ge:Kބӵ
p����9�T�aJd�M�Ψx�lS��EXR������5g-"c�8����O>#����+{�֩�	���x��r�4��h��f!$���q���u:���N��}q�vUXd{�ݯ��3�����VH�	@�m�?Sv�&/<�)�����K�۽t�c�gR��U$����|V����3f\��8#��ulEܸ|��xp¯8������<{�X�5(5�T!^,Ss��G��yg-"�ÍŲ��M��CΘZ0-@�_/C�<Q�)��X~'O�![��F�M8tFu��1��C4��}4ڂ�LS�vּl@�_���8CʛՆ{n�����1/H�-�1��FՇ�c�M$�8i+�3�ߙ`�x��S��H�;P�L+�Ʃ��|�!�F�Z��e�`s�A	�NcHۆ��8�ϟ�4�2�f���7���\	�@vL=��&=���'Ji��mF~.�!v:t��3���U�6��D����Ӽ8ݬx�6p��v���0쐸�>7k�bǚ%#9if�i;�����-i<R&�n$����*'h��j(��jN���npc�e U\�*C���svD�mV^ӻ<ݷ���&��n�Yr!O=t���.{'6��8��#xu�9�9۠(���]����߿n�޽!�֛l1�Vʩ9��n��������n�[�/�����f����=:Hi�Ѫ�*4'��/H$Zm�\o	<x��8�^\���G�s�{�yg-#<�N#/%�����+l�Hλ�K�N�yN�DЋ�(��_}}���_-2t���Ǌ38d%�I��B8�:]�z��%�<�#�$����=��
nפĳ4JAüa
 ^�V��I�O�#|B��H�90�	���푚v�t����+R����	���>=��(B�8�s���ym��)5�����E妓��4���!{�K�h��HH�rljvA	P���[Q�p�d�d<l�7�<C<p����j
�1Aȕ�.ɂ��Ǌ8�5S�����:N�Ӡ�T�b[�'���.�_����B����`z���o6��T��j�����Oϣ4�T�g:4�#�3��XҔ����g!n8����s˷-#�P�R�Z�`���Q*��!x�=&��E�'yx�s\-�A?�J|Fu�[]:n���!�:M��JH�&�4���~�
n�<Q���J����!P3�xAM����f�jV��ڒ� �~�	<�!e|B��$x��K��t��iY���ͤ�0����M��M[�{�;�D�TJ�+T�?q�<����
|ꟿG���P[�����!k�>�d��LO��x�N>�E����p�7����m1�!�p�l��M*�2>�
o>���h��se��a��
o;0-�Z�U��P@ RA@�  "��Q�����N�>~(�v@<���a�`�+�:����EBW�KBB��(�Z���` КQu��'��R!tK�P�z��AQ� ��Wݍ7οp��+n�Q>u��=�D����V����7���X�ΑH dWR��_*��� t�<m�>��~�^�TQ�
�]�G��u��=oWP~�� 5	�'O�v"t�؂u�TQ�����'�� �0����c����n��J�"~6�dLt "xϚ f;��Ѳ&!�~�=Ӿ�PJT������*(�
�D���Lb�Nk[����4cԊ�;��1+��ps�f��(s�ț�r4roa_��_���`�a�3����������8@�f=�?�/���>��/�+H�>��^�� d@�:�:�/�G���
�<(��Ҍ��#�=h�h��O��A� �h�Ȩ��>��(uPa�"$;���hD�����!Ȳ��.� �-�4���%�yy��Eh@�`�B%�8�\P��7�,�"Gkƅ>&QGS���P�:QG���!�s�~��~=gp����C�窝h����P�i�x
y���)���:�QG�t�\����gө�W�OH�w �, �^�Ah��N�_G�Ƙ����t�@��΋�-�t
q�J�{9w"s�"'����Rꆈ��E����0��=�%���7N����+Ԣ\*ȝ���/��%'I�!qN�! �܊�c���"�(Hhs)� 