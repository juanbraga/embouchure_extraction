BZh91AY&SY�^�En�_�pp��"� ����aw�                   �                                                      ��  5F �` �,c@1 	 ��  �!��(*VG��  �X�P��J�,  MR�-R��j�VZ�U���]�          �R���X�U�qTb4R� ���"uC�V-U*� �c5J�&���R�V0�*� ��X�R+�UX�R���EW  MWZ�T1�*�c5U+-
��          ��X��6V6�UX�!` �u��Qێh�e�J+��*� wU	ŉUc5R�-J���+  A���խ.7WV�q���]�  Ƌ#U]q�:��N�           �WZ����Z-Uq�B�  ,��V6�h�7v���*�� �UN6�X�*�څR�R�V  ��N,��cjX�R��  �:�rԪV6�U1�R�����          -T��ԪU��U1�R���` �R��J�cT��A�  �d��Ъ�UTb�U0 �lj�����h������U` q����1uѭ�꫶x t��?@Mꪩ� �4F�hT�$=*U(h2CA��   @   S�ڪ���TѠ��0@i�MJ��	��D�F�mL���H4�b�T�  �   '��۽�����o��o��z�^�/W�W����<z|z~~�l8�_n�ca�ll�o��6#l8���6�uن6W��1���~^[6���U�|�k>v�]�0��9��u))�Z�E�[)���)wmӮT�L�Rȫ:崙Jۭ�U2�Z�+Qk-[T݉2�L��IҪ�N�njY"�Q��M��e*m�����&t����*`Jd��j�Q-m]�L��V���ʋt�j�t�ʳ���*��!hD���L�W+.���M�
ĵ2֚�S+SS)���+Rj��kU[�L�R�i�L�S)���L�T�S)���t:���qڑI���L�[Rn�r���N)�2�[���T��2�L�jԓS)�ʡL�S)��2�L�S%�e2�U�H�Tb�&���Eh�-�(mij���bZ���VͲ��Q6[b�)��ZT���j�Kj
	��Z�f�-hZ�GQ+)����MZ�)�R��52�Jڜ�E�UJ����e,j�ȥVS)��emJ��تe+%�k+iS)����3�t�V��̭�e2�L���kkH��YmX��d�VԖ)��X�S)��j�-UQ��U�&"�IJ�ٲ�Վ����2�jm�Ӯ�U#��j)*�)��)�e2�L�S)�ݮ�L�ڮ�L�S)��e2�&S)��e2�L�S$�e2�L�S)��d�L�S)��e2�L�)���L��t�e2�L�)��e2�]K:e2�&S)��e2�L�S$�e2�L�S+jP�I��e2�L�V����s�L�S)��n�L�S$�e2�L�S(U2�&S)��.���)��e2Y��)��n�X�+;�2�]2�L�)��e2�L�S)�e2�L�S)��e2L�S)��2�L�S)�e2�Y�t�e2�2�&S+::e2�L�S)�e2�L�S)��e2L�V;���%λ)��e2���e5jd�52�R��S)��e2L�S)��e3�t�d�L�S)��n�L�S$�e2�L�S)��d�L�S)��Ύ�]�,B+���:e2�L�í�t�n�L�)��egL�S)��2�L�S)��et:�7&S)��e2�L�S$�e2�M�)��e2�&S)��h��L�SRL��l:[+((�mR$Җ*T�gL�st��M֦U++tuZ���趙[wlۦڤ�h��UjԒ�]�QYQ-��RU�Җ����m��[f�l�vS)��2�L�S)��e2�&]��m;Ws)��2�L�S)��e2�&S)��e2��e2L�S)��e2�L�I��egp�m�)��GL�S)��d�L�S)��e2�L�+n�s��2�L��:�v�Y�u���ev��S)�e2�L�ML�S)��2�L�S)��e2�&S)��e2�X���]X;��b�N���e2�&S)��e7u��L�S)��e2L�S)��e2�L�RJ��GY�t��L�S)��2�L�S)��e2�&S+����KWN�n�[���d�L�S)��e2�L�)��e2�L�S)�e2�L�u�n��en�Ιɔ�ۧZYL�S)��d�L�S)��gL�S;��7]S)��e2�L霙�)���sRjVt����[ws)�ʡ�3�S:e3���+(�S)�Ι�)�e2�L�S)��e2L�R�U��2��̦tΙ�)�ΙL�ws*�T�e2�L�S)���e2�L�S+(��L��S)��e2�L�S;���e2�L�S)�i���e2�L�S;���e2�L�S)���e2�L�R��)��gw3�S)��e2�L�I��e2�L�Q�tAuN�L�50V
�V�4���:�+u�[m���Y�ڌ�5`��j�ms�����՗:��uq��2�f$�(SV��.�Z��n�Յl�[��:ڙG]�f�j5m�1˵X�V���gj�u����[B���Ee��rn�]vg.��1�VK5Ӎ�M�ZȷNuwN�t���6��ef��:fۦ�Θ��Y-�wr��v:e�j�Y��Sw%��:�s+u'.��tj
gw	VrefVu��u�g��u���.ۦZթ�3�S:�N�l�蠭�2�.���]��.�jMU���m�*7L����Iݝ���tt�el�P�GZu�[,��[*�ښ�9�ݎ�C�̭����ۭ4��u�tI�l��n��t���L�Su�e2�J�M�NVt�n�]ݎ�t��&�u��L��gL�S:g[)�uS���J#��������=D��$�4��I!T����  `@��YB�ם9;�w���e6�Z��2˻�^�j۵s� < Op �>��(       p�       �m�p m�����P  lm��w�f���is^�omP �    B�N��@U      �  �     �c�^m��wu
  w�<<��p�@�v�( ' c*�6��j�kt@x x8 /T�` < 6�+��]�/l�p0  N ����	��8@x x8=�^�  ���nm���Uwv��{7�M����WsÞj���sݶUA8wg�\��x����J�u��ۖ�8@x x9�<Z��=�h�3��������6 OOv��@� �p0  N ����	��8@xP�` < < �����U*�N:�����8@x x8}����l�4�`<����;�0  N ��   �@  �0 3�p0�ǣ3�v����8@x x8  /,��l��ޖ{�t��8@x �	�]Xw�����|����qql���j˫QY�| N �  x� ' c ��{�' c��P  N ���y�k��8@x x8 �8  ' c ��� '�<� c��8@x��	��8@x�`> '
�y����	�����w��1�w��N�Px x�	��8M���gk^x!�t�c��wc+���u����  'K{�����p��cx�žW�z�T *�@c    ��V�R��V��m��� �  -�l x ��]���@w6��M�wu^  U  ��� N ��ʠ��Q��=��2���n��*��*�����ҭ�*� ;�  U �K�d   � 	��xQ�ef��Y�^�`������   
�  +2��@�  ��Ϳ_~�@             � ���mݴ���Mܷn�  .c�m� *��U ����+�Qٞ���1�r�m�}� �l  ������w
l�e��
�:��w>�P�>=�Խ�Xv�wm�]O 'U`=T*=��q��Ψ8S�u����+({;�P    .{7Z �Ͱ x   R��    �     
�      @   Su�۵�  ���͵Zc���5�      [-�    VPU� �u@  U   �[P U �    @sl      �;� �;��:�  l U
�e�p  Tw�����@  ��[      
�� <T 6�m� `  U
�    �   � p    6�����l   �  �ݾ�      *��ګ���Ww=^��y�zN���[:sG6��r��6��b� �  Y@  ���W8@ ��]��*�f�@�Nn-�k�J�'o( ��Su��v띘�TUTg��z��Vk���6�fvOD�� �  *WD  &��R����jo;y���Hw6�    ����#lp󺻧�૥�w`.�����9ϛO]3b����rzmۏ6n�*��m��ޟ~����{��v�U�m�e�V�^�EP�q   �  8@x��`=YF� N Ϋn���{�wZ�^��w[.�[h���wnn��     �^��    � l   �:�      ��  +�
� 7`  >���okwd                                �ml��J��         �}     �                                                      �  *�           �>��                          ���        �   T       P             �      l
�  �}  T  �  � �                                P       }�  �   T      �                        T                      l P U �
�                            U          }�            T *�  6ʠ
�    � 6�@       �                *�U         ��     �             �           �R�   � ��a��   EPU� �����*��                 @ v                                           �  �                 ~��    �    � ���   p         *�                            U+-�uR�      ?A�     �                      Z�P�                      m�kj�  �       ?A�                           ��      �� ��                   �             ^�V�2 x    AT         T                  }�    �                 
��                  T�                        p                            
�T                          ���}��                @    Sd@ �  T   �R�               �y @  *�@   � *�*��    ��                 ة�[kl  �  *�   `EP            @          k���< PS��              *�*�    �@��\'{���zw;�  @Pw�^�m� P            U        *��P `�{kl�k�[��P�U8@  ��� � -��N ����	��;�T��p � �     �6�` < < ����P�TNՠ ��"p6���p [;������ca��}^L������~�����̓^�?w�w����'=���������<�x���w���Y�o^���+̀  �5� ��n�` .�   [E�G{��w+��݄�`7Zz� ' c��	����o<6�9c��1�w�  N ��;���D�� �=�*�(�xx8�_4 ����f�: <9⨜����^#pN �;8�<�xUn�0<+��N��� 
�Vڨ�g,t 6��m��՛`7qlյ�K���  ��qY���[\�T����
�)6�6�l��
�  �T<ZZz�*�b�� [hT-��d   ��  
AT =Y��g5�*��\6�t����{���ؼ����΁գ{�y�����t���y�ղ7-�W�U;\�e����'�w���S�m��       ���T
�P         
�  �@        T    
� �      TTU@          EP     U P  *�`
�    P @   w    
�mQ��   �    �   �   @  U       ��@m�   p    U@�     U P   U  b�T     @w   @        *�             *��*�*�  -�  ��   �  VP �   VQT    U[E�[]�U  U *S�� ���6Ք
�< <�گ�>|������wѕm����{dv�|T4�9��\��z�-t�c��Z�[����f����Ub�[�;܁s�)R�[*�r�n�m-6�s�5K����y�@6�� U@ V� *� � Q�TT ��
��;��T *M� @�U � �� P 
� UF�<�\�^�l �>|�S���m��i�$�SI�H$�D���u]�U��[j��UU���I�X)�h$�y�S�0���C���c���P���j�N
�,�ʙab�/^,�q
GJ��E���$�qB��Rȧ���#���O�t!L6�H�a�<i��r?\����U�V2�q�$m���^s����-�<���B�祤?Yxzi89��%�ܐ2��ͨt��zr�4�6ƹ�"�^�H�:��FE0��<��i'$mƒQ��YL���܎Rȧ���#���O�t!L6�~���<i�t�x�i�m9.nIG�P^��v��@�m��Ql�¨*��]e�n楔 �"�������]�^�<�3Oz����pӄ[���R8s�d`ӄS��$�ZAp��m�"��R!��y+�AK6��<�x��G���/T8E<>��2��Nu�aN2TnI#a7�O�x���)>7���O�%�#����b�mT���58ۍ��$�xi0�r3jE=>��G��i�P�b�Np����n!H���ae�
IC#�G� i�S�r���i�5�lRͨt�K�,�����c�
�8E<7*���V�^�^�M���q�gS��^� ��PxU*���
�U�g-yܘ*'$��ّ��G=��y�O�x��b��܎Rȧ��K�
G<05Yn�$�&�nI!%��0ڇH�.�M#��76��S���yHf�u	�)�S���D䐖�m�X�y�R8pz�@���奘)��:k�إ�P���YO#����KI(�nI#rrj"�^��H᧼W��}L4��`��)�*~����,�x}g.��rH�m�܁��~ᧇ�:�U?`���	�#6�?S���yHf�ue��"���{�om�5vml٪Ԁ�� �e*�� �P ����ܑ�����m�E8i�:2��qS�܈a�ܴ�"xgMy�j"��\M�đ��*6�qe<4�S V�����α��{Ŗ�2)����e<�)9�P��H�-��	���O�,�x~�a��J��p�E�Cv��r�DA�5�n6�rL�3O�x�+
0�j�Q��*%{j]H��+V����B;Xhcm�ے6�IȠ����U���8}L|�S�x��2���ze������+�D�	Jw��=ɶS�l�܀;��*�t �6¨*��[R���r�QT7��)�t��ds�������y�d>>"\SƚGO�W���m��J[��G�m�#�C4�������(~4�0�ۑL#ǆ粑!aƠnI#n(�C4��%r()gǄu��e,�Y�L\�҅��U��Ef�3]\BGn%R(ڂ�|xGF^,�����y��G�|e�H��t!L>>#���A��R�I$��r�GH�܌�����yHf����<p��eƚFҸp$��H�jB�rF�ż�G���l��'Z�ѻ���U���=8�j��;���lVM�u�P�m���[��U@ e`�k'p�wx{v����wh��۷�����    � �   yT  �UPl�PU�*�P6�� 
��J�lU ` A�>��l�m��W��T^���j���|�l��[G�����3张�x�dڨe*��m��ɰĒ t�)�F�Hf�ԮE,����r�����M�Jp�=��6�F�JI$�8$c)4��qAL0�yRͷ�,�x�n�'f)�J�G8k�鈴J'$����@�0����q�i"r3�����yHf�x������ViF܎)nC^�R0��L#Ǉ�ipR!��up�N�:�ʮ\/֒c`���$�n6�rAX�<p��X�G=2܌�$���K6޴�h�a�S�6(}���~�p�����m�m����Tl;�+�J�;�*T wn^���I��n%$�I"�0R8i��S�R0Y�x�H�[��T0�z}��G��i�U3���*'$�&ۍ�jE�P�m�����z�F�-,ʴ�"�خEU��g��2����[�YNG���/T8E<>��2��Nue���a���o#����j&rH�m��NGU�Z'$4R8i����j�1Oi"r3jE=9�׍���4�RH�	�R��C�q��8i�</�
Gv��p�xm�a�H����QX��I/ħxV�[�j֞�@�m����Q����
�����s���]�RF[j
Y���{Ŕ��8}L|�z��)ឫ:�R8iά���L4��Q�K|��rF��7S8�#���#��)������p����)��)��<i�p�넳J6ےI$��g�"��r���!�{�<'�S��#�(~7�p�j�������	*��M�IH܅��i��\j
Y�C�y��e<4�S ^�p�x`�Ρ��4�P�gβ�HܒF�N)��т�,�q
GO��G+��������x�E���Tz�L��`�8�F&P�#jJ�ش/�� C����lY]¨+)k�����q�m�Hm��GH�܌چOO�{���=��R)�N�x_��R8z��%C
i(drH�F8E<6�,"z}���mC�y��e<4�S8��C�S³=I��TNI	m�#�1��s�-�dS<"w�^��B���{��Y���^�pR8iၪ۱�"i5#rI!B0�0ڇH�s�� �#6��S��^�<�3Oz����pӄ)�A��TNI	m����q
Gz��p�xm�:f
D4��.5,���=/x��G�����_��ʵZ����;J�5�i a�^�U�R��wc�+�SqHܒFے1-C�S��ѝc)4�V[�ȦxGG�/S�B���{��Y��⤺���"I��r$G#��E�1L6�H�s�� �#6��S��^�<�3Oz�������I$�@��pӄZ8���R8s�d`ӄS���L�4��.5,ڇH��
��L��q��)YO#���'�"�곬e?S8������w<��S�!H�����F�.5M��G��}.R�Y���;A���s��F}�0��O3�{2H�;;�Z�ژOk��}^�c���p{m����{{
v�v���\�v�&ʠ𻪳[n�m����*T[`	{{���;��'xwn�j�_3�|��l�      p *��  <   *�� �
� 6�p6� � *�� T
�� ���  �� ���<v��v8����N𭫰U_m}���u 6øUU�UQ����
�������zj9$&6ܒE��~�ޡD�4�p��_��R8s�d`Ӈ�=��`�a����H��7�F�q��>�#�׋)��^1;P�<2՝c)���n6G�>>!N��#,��d�ےH�e/�R:|or9���{��
G<>"����x�.b�4���R�R1��d���=�0���{S�<��S�����eB�Ý�#�?a��B�1��Hۊ�H�OO��S�}�8G_�S�Oּbv��<xe�:�S�3��֛	0CĔF3E��rP��l�� ��گE��������b2&R%(�n6�R!#�:��_�t���sş�����pR8i�6�g�C�_L7�i(��I'͵����ϼ���y{���P���g��������UG$����#3���O\�����{�~�W-�sמ寧���24�RI$���bמ����}ܫ-��G�8;o6�򩎘�_�B[l�d!���.b��b���ݷ��-�/��@�{;�Q�%6�2G{wl��r�f�MIۭP�� �e*�� �UJ�ۉ�{Vʉ���uKsܦc3�ިO\�����{�~�W(]��D�$�q�c���-��bמ����}ܫ-��G�</�#LPF�n�I�Dm����g�ڧ��/��33&K�M�L�K��)�w:M6녆�v[�&�&n5ۦn�~Dt�ܒ$�q���	����~R>������3hɣ�3w:f����U¦M�f�&k6N�:�L�Ι�fn6	�k�P��~Z��^��އA�����n6ڑ53pɬL�$��
Y7��7y�6���M]�Y
�7�q6��v�%�hɨI�d�$ӈ�d�$�nɻ��`ɻ�|���!���X*�=ݬ�l 6øUZ�*���dU�l�i��a�)�%)����|��}�����2n�f^pɼ$��P��4��u�5�n]w036�ˆK��l�꘦m�L��>���������$���ے6�M�L�$��&�t�ں�*)3`��3&��g͂�tۮ��fl��p���Hɽۼ�i3f�f���fM�Ô�d��" """f`��I�6c�oy�7N��fљ�ntMx雼�f�ɷ��"�&Z2h�>����������a(y�q�$q	:��fm4[�m�L�.�˘�R{˷b9��H�\��p}��#"��]T�Yn6ےF�h'&{�q�Gw�Ĵ��Q�o�V
��&���U���X3�����o��!iG#I�2��^���PC����lY[j�
�������2LQ�m�$�A3j"�f�>'�^��w�ȧ�}���-�#�.���)x��|�B�j7$���r`�a�xA�v��Gt/4Q쩾i[��eC���s�x7�W*��O��q��d��2��(]����\ט��E���;˰��R8iN1K�j#d;衁��J6�n	� a�+�g�"���|M��;�܄R�یNսB�ҹ�Ԣ_(ܒ�fF$c ����l�H�H��.�9���=�7�+{�P�!k\zr�gڒFGm�JF�e��7ӝi�%� s���k��w��N �aOm�����n�>T�� >+�u�w��@ض���-�w�z{^��]������=s���<� *�  P �     �  Y^�*��+( m��U  T m� 
�U� C�}�k�*��rܹ���kKWűϖ�u延�t���浺� ��ݳ���̠;�*T^n:�����1@�x����\��?s��O���c�T���q`�+�y�L�U�k�bP��8[m$������1e�{T﷗�61m�_���;�i%m�$nC�{y�{��y���ٳnU�weYm���#�݈+Q9$I6�nFd�ۼ����.���c��ڏwƶ��SzL��I$�Hd�n������r՜b��=��������� ���!N'�櫽�<��ݶ{0 ��U^���6�Tz����.u�we�O���+x�浆���K��x�*�5o���w0R��C�rj��#�H�%ƣ	�Rxn�#��t�zo�Cj�Z79��[�窜B��_w��bm�$��ےHq`�+�y�L�EW����8�Rb��z��)��"�I6�#n6䍴�ω�w���ܵ�]��Wz��k+��K��x�ق���mKWe�D�ےC�b�9м�G����o�A����Y�qϙ�r����t��]�F[�ol�g�k�U*��ǔ U⪯E�P�
��-�kl��;�"Ͷս9z��):;���)�W��`�)4�".�yo�q��5��HKj�6�-�3�O��7�>&�ޯJm�\��.UoA���a��*��7��I�ۉFԑ�&
FC�;������=�7�+~��v��z�F9�6�U6�l ��1�$����F�<Żz��);��#�)��<�&#��DC���!�+�e�q�$m�؎	�@��n�3�O��7�>&ջ�6�x��*���\ֻFLK��r�S�m��m*�zt6QAT��
�+2�pJ��ʹu��mo=2iI$���`�^�͘)i�w-s���^h��S|ҷ� ʇaZ�yǦ"��D䐖�-	|ͫ�Z79��[�窜B�㣻�,��}O6	���H~/u��J7�E��0�;�kXy*Ɔ����Ws���*ơ�{��{nZ�[Exu2�T9$I6�nF�˫�CH�ўcL���U��cS���Gt/4Q쩱�#�C��:K5�I$����CZ�X���aF#2��1�kԻ����5��OdZ���{��i����T�S��ٳ���S]��0�ª��*�� U]��u��ƃmT���U*�Rt�ݸy(,+��o���˒�{�~_�"��%��2E���o�//=x'X�y��v��-��;�CO�9$I6�9�|���-�R�^\1v�X��v���Č�(ۍ�#l&�g�<��`v^�|���f1n[.H{��j�L�FY���-���)�����{'�q����ׂu�睾�?o�����{�M���䫣m<���ŴN:�{���Ͽo�U��d �3��wm��aܶ��	��=�=����y@�z����P
�
�m��lYG���ۅ�9��_9܀U      �   �  wP x
��*��@ �` *�;�T U  @ U
�  _k�� �r-��n�ԣ�_;ӥ�o���P^�W�P ��U���ճt�ՔGs��]�w]�)�U���w����Gn{�܈��r�W�˂�]�_��p��m�$�I"��^_���}��C\�#��
UcXƼ��Έ�k/�f��p�up��<Q�m�$2G3�1�~}f�X�0��uص����J�U�ZGN]Y�0a����tB�j7$�$�s4�:C�w
g��7܏4��}ʌ�v�s�h��0�#������ۍ��$6�
xG���f�C^w�dŨk�dw��J�kו�Э]#zL�@�E6[&9p4L*(�M��e��V �� ���QR����p1R$�P��i��c4�#�w�U�����nU�C�=��{b�<j��1�귫H�\�c@����d�$C5β<vIcVƽH.-s����D��y�i6������)�ײ)L����"�ɚC7W��78���8G`�jo�ˁ�>��Sj�y^�U�coۨ����$���I�i�V���ә*Ɔ��ț�k��a�V5#�7�X)�G��_Ci��$nH�b����k��+T�<��K�5ԃ
y���5�iG��I���uj���e���X�ެM�p����
�l 6����.��vh6�F�H]]"���&����.�#X���*o�ˁ�>��Sj�y^6�dn%$�F��H�i:Fщ�v�����V45���&o�����7*��\:�=q4��Ē�����5mx2Uw@Ʊ�{*յ�Y�X�:G��Ńǘ�zF:�֞�#l��m�܏4�#�h�Ȏi�<7�)ںp\�M#�vnǛ�#�J��4�E��p�ےH���Dx���̓4�c@�%y�x��A��hk;2����M��#-����#hI�"�mʧ��7w �;��ދf�m�(*���l�ޔ�eD�q�$H6��!��D��`��V׃%Wtk���[^yp��Q��鑖\M�[m�$B8�x��ֺ{J��r�)E�c^x���i�WN22:i!��^��RF�!*�o������ʛPם�x�+CVƎW�ˏ5�vs2U�c��S� ƠnI#m��<F�����!#*7.Z�ƭ�J���ƫ�V��b�t�H�6�Q�$��H�J�Aq�n���).�x�g�N���}��w���[y��{wm�n-s�<U�Tl;�+ٙ�;�*TN���hƤ�I>m��1�;�c˪�y���6��;����+CXƎW�ˏ�
N��I$���l��f��p�d���k�_�ܫ����-y�G�xĵiG؉G���ĚRI%J�UR�[^yp#��5Lk�ů<��Z�{lhkʌ�5�y�� R�B8���d��"�ӃfFGN��m/M��ןY�Sj�yR��sX>�[��2IR(�d%r{���d��u�io�_�ܫ����"��B�C32d��;}��b%L�ʙO��   ?��U}m����z �� 
�-�޷v�o��n�� n*1�p�� �Wo>{vצ�oc�k���w�7�y^)�e�c ��U< �z�r0�^ <�s� <��v����۝ �۵�V��8�c ��' ' c � q��<���y;�7�{|�^w ���x{�j ���߻}���U*�E��ڠ[&0=�^��*��� Z�( ���   �b���=U	�¨u�wk�^ʽJ��W�؃]{��    `� �
�U UU @ *�@ꓛg]�@� UP\�Y@ V�C�n� �������طw�����m�6�����q�wn��T ���y|�ܖ3�p;�p^�� N��      �R�  @          
�       VP       �  ;�                  >�� U U             �           �  *�Ve
�p   �    w   �    
�T       U  `   l    �@      p�      [�� C�        �   @   T     U            U   wU  @    �
�T� T  *    *��� ��     {�� �Pm��qms ���8M�e+��}}�v���a��ż�Zc7h�ԯ@6:��v«+�߿w��ߨ�������S���Aqꢮ�6*`�Sl;�`pws]{����m���ᶺ��[�<�@  @  ;�* �@     x`��� �w�  � � �@� 
�   �  z���^�ϝ�۽�Gr����r��^��5�� 6øUUUQ� 
����2�ܯvh6�F�m�w�������0a<ţo7��R�^yq浨����>R��1��Ĥ�I!�G Y�p�-9)T��]���k_5�m/M��ןY�G�qm�L����$�n7 �Ahk���W�pt-k3%X��0��S-C�S�y���!��\ʁ�mk"(�-��
9��xFn�jޡ�t���*յ�.<vJ-[�aqk�d{��	�v�K�"rH�J$Rq摤q�*2�XBֹ��B��z1�-x�!�۱��CH�Z{�I�ڟ ��u�|��h(n�=z�P�*��[+e����m��l�����
�
��k�dw��J�cq+�`Fd��ř*��5�̑�ݪu4�m��nH˒f����U}�dS�0��%W��5��W�V��u�z���"��K�\�����ł��jj{l��ܨʇaZ��ˡ�;���7���#�l�鑖\M�$�I1��uN!�x��E<����ձ�W��е���cCX�MTJ�Hۍ$�pI�F������jG�)7.Z�ƭ�y(�#Z���0�gEӽ��Zi�a�-:���@��m�� 6ø*^̥P� �PUy�����e�j��~w��޼��מ\y�h�lhkʌ�w�c^<7AܚC;�M��a�ۍ��!��k�Ƥ}�M��ןY�Sj��<*�c9��\�5�#�[�e����#�)�#H��.=�F���a�5}�#ϔ��-y�V׼��^��)+=K���������x�/]�R�Rh�+v��o�����c"���a8w7M�����#������a�f�>��1Y�b�a�޸�q_S͓��H�J�"���%�]:�w9�����yY@6øUW��*�� U^��h�z��I0����x�#6��3Hh~׹H�<z|3w��U��.�< [���I9$nI#rD�g�p�G�3�`/��x�׈�s�"�#os^R]��TNII(܁��G���}�9���kXҁ�7��5�a�O ����kQ%�7�I"��&k4ܮrG����U�+|�ė�a=>�����ɩ��NFbIF�M�dx����'j�#������x�"�-�/��t��u�rn�|�],�״���s��@�wUz.j�mYAT[;�������uWu#m7#�@���Dr��<xwI�>&�N�̌�� -6�yj����A1�ˊI	��$�G#�<y�g���iy�W��k���V4��_5mx��"�l���q�$m�ܙ�6��w������N��<G��0���<D> ��:Z(țd�ےH�rל�y�h�o�V����5�y�8���mT������E��
MIq��e�Z�E#�G7�X�b���X)��W��k���cK#�d��.eoU����=�Ou3\�O�u��� Nv*n�ϴ����UR�)��@ws��[��( �k��^�4�vzoZ�w���P�    T6�   x�  �    �*��� 6��*��� 
�l  U    *�Uz��� ����j�����W����+["*�ж�Ѐ�� ��VeWuR��N��&B�1��H�a&�4�"����ri�u�b��%���O��X+7mWX�<r/h�[셦�n6�Q�
D|�R��kZ��E�J�y0�7氏n���mT����ԒI m�#Ǆ�ݏ-\"�㣛�,�1_R�f���r�����[k�QΦffF�m�dq�
�ڷ<F{��܂�t/nk�=ᱎ����,��СĚRI$a�#S݈{��cޞY�wos]��;�_����1��X��!1��m�ÉUl���+(�w
��Q� dU�(䑲AQ��-�����&���n�n[�������ɷ�u�޶�n7�7	k�{��5ʏuo�=�f�Ao/�wy�����rH�m�$P6Ƿ-��S�yO����zyg�ݽ�vQ��#���n%$�I ���ܷB�ۢɯ�t۱ۖ�G7��'���u��rH�I��I6���*�{3wxF̬�V�r��w#ջ�M�&�*DCA��ש����]�s/*�U^�el�Ք-��U/[�T��Wu*�;�٘�/-��y��:��9G��[�-�^[��@���"�H�J$R��ܾNLs�;;�����l�.�,=�Ӓ8$��ے6�r;�{����a��Iݗ�d"��z���z9�X��1m��Q"��V�v���;��C�=r�z�N�r�Q譖��Iq��l �U���kչ|���z����tv����"�J��M�؍�ݺ�̕Wul� U�
�R�w PUw;��]5P�����{����9}NvK�-���NzT,���*%'�F�m�$e�,�;=r:�����W.Z1�g���q�e�:���gIq�ܒF�-�!����X)�T���69cX��P�5�.(j�@���Rq�i"BL`����4��M�c���X�{�p��V5�x�q)���zH��i(��I$�!c�5���M�����T�Ծ#�r��X)ᧄZ'�����/+\D!n]ͼ��w]ҫezc3�( ��U^��ܪT��KOw[{T�FF$c)��U���CM=�o
gz�m�c�5��D^�_<k�:�31:̉4���$`��H�ux�sD:k֨a�6�kϰܩ��\�`�窯H��¥�7�N)$���M��3���u��vƵ��ɱ�\���ʛf��=�
xi�٥�6����7!�H�n�#��Gx�S�)�U���S��mwdZ�Y���(rƭ�d(�
��"I��r$G4��xwN�3J�;E�R�=j�SaƼ�a��O��Y��%�!$f$�($uX(u�۬�*Z=��x����b7��w�8buW�Z�v��-���!{eT*��mP����y����o�+z��5ת�gu �      �   �  w  ��x
��;�U lm�  �   *� 
� *�l�m�� >���l��t�W�_7�Yu�J�A@{�{��4�
��*��[+e�����}��uS{oE{d)�$�3�s�?���A�g�O���3]��e��,v�=~�2�ƥ�y�XM"j'$�$�o Na�O="�8��\4�^�O�:��"i�x�S8����q����-��m6�K#V���\��x�D[��a�T*^c�P�*l#י8L��v����n�fjfTL�X�{�r3ԦƱ�d)\者�g��V;cZ�}r_����[m��#n6䍴܏4�wW|�r�n��G*�U�ak�U�U��iΫqi�HçM!����,8�^8ln�67U����� U�
�R�wT�
�0��9j�U*��C�����(rƭ��P�Z���ȷCT�4�eS\�=k�{E&����P�܏7T�G��qf�=�8�T�CXǌ2�tG���y4��:w.i�@ܒF�E52�X����ʛ�����m�C�=h�Y*��l!�|j�J��C��qj!��F�m�H<F=>��ŃL⺇��H����TmC�!kC�b"�Q�]�9x5��ԒI#-�#O��\�*l"�ן-=�cƇ��Shk�B�ΈZ�z�9S3M�WUλ�Z�UlR�J�l;�U{&ʩ� U w6ӷ�w��UW:��V;cZ���4?>�r�ƥ�{г��p��ZY*��l!�y�[Gɡ�3#�GR1�xF�����~��Y�I�P�[�7[ز�#OM���$l����i6"�cT���`�*��1�U�2��+"�C2də�.��޸�a�?o^J�\.<3�]e���ƓR(ډy�u-k8��c�5����4?>�r�ƙ�]��7��ӇOHS۠��Q9$I6ܒ(c.��#�.����iΫnHj���A�hu��ԚEX�����U]G�����^��UJ���oF��m��]�l���eKm�<^F%JF��$�c�e�:F���"�S�0y�Ms���S|Ed-#Ǝo��O�Ϋ���z�qI$I$�f���M��c���̸Z�x��V<cZ��ʾ!cC��7*ljXF�+�6�ߣm��m�H<�Diç�m�Wtk^q��V<hy�ˬ�CV�:�w��b�C�k�@��#5$f$��1c�5l��ً��=f"-��0�#yT�1�Z�a�7�VB��Z��Fb�6�nH�	��O�έ��@�c3��e�Bֳ�^J����5˨p�:s�F�����1��a$�=�̖]םn ���*�C� *����mT�۷*�о�w����סr�*���%Wtk^q��V<hy���	�5lz�TN�S5U351S32�L�Z\/5&�C�5l�tl��Z��j�F����k�ǭU��H�.&ےI$��yuN!�xՇ�,x��`�3�6����
W2�����y��H�� �Ik���m�$���!cC��f�X�0��.VeCC�1��d��ak�"�*Ǎr/��K�\j7$���nF=2��,y�!y�4���z:6�_���QniwWur�p�h)$f4�Q�R6��2��m���6-0���� ����.f��ݰp=�8A� ;��E�1�]ԛ �� �
髻���ӊ�Vͭ�c��      ��   �  ;�  S�� ���S�   w � m�AT P   U  <�^�W-�MZ��gu��u:�WsgL�W�� a�*��@U`�6�w#׻�[ʦʮ�n�1�U�2����C^}����-63Ԧ��1�;!J�\-k�H�M�J%$�I"���ät�5˨p���ܩ��a�\�ʆ�lcG*�Ujޡ�t�ΰYA6�HKm�"���Ƈ���;CVǮ��E��^k��)�H��f���H�Ù��l��jF�B�9�CO:�nl$S�OH��7�n5��쩱�C�q{JmsX�����1�ӊI$JF�m!�O�"���V<|ֳ��![C+7"��|�xK���#t�]�HJO��ȥe��ʶ���޷@�m��]ʨ�
��m��l���m)@�����25�ݪ�V<hz��Y6����^|dZ0���+��j�VB���j�I6�m��.��4��0�3�I�:-Sk�ǭW0ʛ�+!y�ʫ���ίpo���7�H�i6"�񝐥s.8��g�̕c�5����!cCY�ScR�7�U�4�D�D�UBM��ȈӇw�E�ռCH��g��x~�)�ꠤCO�[ŃO1n��9p�q'�(�-��E5�Y�0�v�_���!ۡ�aF*��\�>�)��yuN!�xލX�D��a���/VŴ�������
��^�R�w Ql��ۥ�w��0w*�33UV9hy�q�QHj���Jp�����xƵ�Q5�,hc�����$m��iD܏4�wW|����8F4r��]�l!�y�_�X��E�d��OJ�����iFQm(�"G!��B�Ri9cV�*6�_���!ۡ�aF*��\�=k�x���8�i%-���CH��r<���Σ��)�5�x�cR��Z�y*ǇH�sL��cP7$�I!q��8F�>�r�ƥ�o�r�*���%Wrޡ�t���1�xF��e˱� M�[i�*k���5]͋�����w W���w ��R�^�{k�*UZ�)L���=}h2-.��H���yQ�����]����i�>��iԒI'�<$i���%;��.��C^}����-v �R�CXǌ2�-�:C�Ć�$�F�m�dR5c�5����!cCfQcR�=�\�ʆ�lcG*�U���j_�U1"Y��#	�<#Ox���x4�:u��ȴ<�^jM"�,j�r��W�#ON�ޑ"-�B[l�"�4��7ъ���1�Z�a�6Ykϴ�T�����z���<`\�ٙ�sS�=Eh��h�U/^�OZ� U����*��l*���wZ����[o&�"�fjaZ\-k8��V<cZ� 뚡i�Wu��
��j��qiF�-���A��"I��@���F��w�6U�ƹ�E��Z�=}h2-.9�a^U)f����p��%#p�rDr#��O��)}WN,$x�OH�7y]P�or:�9�8�.��RUTDDEL�UU ���zN��2Qfl}�o�{�����i_�m��m�!��u�����q��W_e��,ޤ��Cy[��"PM��p�Q� �m���哀6(
���ۋ�	�l)�6��n�����UwTͰm�u�od�J��e��X�nw[��|�*���ݞk�_ `�     l  T�     
�T 6�VP�6�  l   6� P     ��U ���ߠx�ru��^�W^�z׏-�ŝ �l��߽��� *�p+=J�P� 
����u��x2z���(����o��O~����^@ߩ��~7r=׻����$f)#n6䍴܎�������;����E�z`�}����
H��rF\������"�mܯp\El����� Y���T�j�n5m�ӏ\��������fR�D���TȰ�O
s��L�*&ےI$��y��G�����,�{��g�Z�;b2%y��5{�d��ätͣ[I"Bm$��&8d�0R���swS��Vڠa�U+( ;�l w$�0%���n4��$�R0�z}��ScR�5�R]C\���U�����˫<�i�s�=�P·��$m��[���C�����(rƭ��P�Z���ۡ�aGki�Z��ģm�x��ç�Jwyn��C^}����-v3Ԧ��1��"��u����ɍ%�I$�H�k�5�ꂸ��}f�M�K�B�FT4;c9VJ�tk\frnb��*���U4��X����d�ձ���ȴ:�^k(X�>�j�Z;��Ͽ�����S�xeK�;���UD��p U�UWtU�lm�T[;���b�I�I5#rF�0��po9%�c�\�*l"�ןi쩱�C�[w����8t��5i�$���I�B�:�Z�q��xƵ�PW����ܩ��a�\�ʆ�lc]e�N����nI#rD$c.��#��Fy�4;ؾ���=~��Y�N�T�Α�vq2�*'$�&ۍ���Z�5;t5l#H�fT��c֫�eM�VB��=�69h{�>�L
�H�JI$��$�ç�]��^���g��c�5��"���|f�U���pn��JI��=r0�m���W��B�e�S�� U��J���T]ϙk��vh6�e~��[�����k�
�U{��l!�|j�J��C������c��A�hu���k�	��MUT�[���Y��#oZ�u?p�hj�F��̩�4s����C��k ��g�4��ۍ�yK"��]�z��öQ
W���Z�y6<cZ�˨p�O�p6�+[m�ܑ�r<���ʌ�S��w�����b�c4��s�=�Zpi�OJ~�jP��"�iH�ł��j!�viGH��ͩ��![��[�2����-ǲ�,�E	��IH$bj<�������Jm��� �����l���r8�i%-���COכ܏)����z��öQ
W���Z�x�O�ӹVi
0�P7$�I�e�8~�����Hguw�Q7����|&�=V�?]�3�4��s�n��`�F�m��Q�?i���X)�V���f�cT��{T�Z�����CV�4��ſD�1�$�O�x��i�N�#��8���6�o���v83Ԧ����R��P���ZĒIm�ɑH�O���"����~�¦ƥ�o�r�*���/��'�ޡ���z����mI$m������=���-t < ���T���ޓ���   ^�۪ݸ��� ���c �
����	��8��w^��8�6���zp�� z�W��	��8@x�U�����=� <� �L	��γ�K�x��招9�Z� x8���� ' rp0���
���� �Zg��. ��^|�@
�7V@m�U�ʨ@x\�nV˅T�u`N �3[�
�l�V�  ���Ԫ�ȥv� �/l�]˖�l􃖎sV] ���x�    ����݀@@T    ��]�6�P����� *�� 
� �7η|�* �˹{���|��;�������D�8C{��P9��M�����os2�md�xz�ocۭգ��=��9;��+d      ��P  
�P            T    � *�    �T Sl�                    QT              �     �  T  x  
�6ʠ ��p   
�    w   �*�    * @    T  6�   
�   ��      ;�
�   
� l            �        �          �      �@  7 +*�    � P    T�   *����@/f@   T�X�P�xz��  � ����3�����b���{M�P�۵SԨ<uh�7q��3 <�#qZݶ���^�&մ�P[�W ]�n+��6�PU�������^�x��Z����-u����        ;� � @ ;� � �B�*��*T U` m�` � 
� � 
�R�*�T< ]���T�������l�*��vr{�@�m������6¨*[k��[ۮ��{�N�j��M*�V<k��_������A�k�dwB�RiC�5O��ڇ|F���{�$E��rHKm�0摇uw˃3U|>x��2��+ vu7�Z��i�NjǬ�S4��Fۍ��tkY�^M�ֿH��1����T��;��B��3�i�W�=��rH�m�$P6�]]����	�3O�:���Ӄ�z�H2-s����YAC�5�R���cD8�n#q�Cr#�WH�Ӽ���0�#ةs���Sa�5�û�,�o{�5M�S.9i�mC��u;Վ�@*Wt�W�T��T[.��ѯt�06�e������#��s�Lb�������GU���4ҿF�%��zC�;7�C�;����\����M����U彫�0�Ƌb'$��15U��w�^^\C]��.g���#��r;��m�#q)$n@���/�v==�:��Ny8ǳ�u�}oJ�t�n6�-��(�~^�{���C�1�U��z��׹A��C����N}<*�HZZ%��%�"h�v�ok=w6�t��Tl;�+�@� aU+]�d�leU�M�ߜ�@G�a�_5o£j����ڻW�S�OH��	TM�$�I1���8����vL���ޭ�y���6�����v��e<4���-�1�n4��%˨>6o9R�wйQ���kì�[�l%���zU�ӝY���t8�nI#l��x4��@dZd%r����TmC�!kC��Xf��ݽ$�Ɔ��n6�o�ߙ��0���q�]Qa��Ҡ��ߟ������~�*0|��)���U:�^�@�m��� *���
�U�j�P$�n$���$�H�����]���۩ 3NTeAa����X��EDTnI	m������4�V�^l��a�Z�C�����(rƭ��J/u���6#��{�&�nI �sZ���E�K\�=j��T�Ed!�>��Sc���#=Jmc:�,mL(mE$���H�y�#�Vq��äk��&�4?>�2�ƥ�{йY��#�i}�D��F�7$BF3uwak���*Ǎr/�a6���s��,y�u���F�Ѩ��mqG�E�z6�k��Ej�����P
��U+ԪU�R�*�y�'7\�m���bH&]C�i�0�#��p\�dR)���G��q
G����4�4��.V5��7�I#��$#�a��<]V�H��1�#�}7N]C�i��YHf��+3�7���NFbm�����hhzׇW*��l.k_��cƇ{˰�CV�9��E���B�Sڝ̳�H�%�e6p#H��Vl.��4���a�v�\�dR)���G��q
G���d�(5$�Ĕ��$�(�9շO=�H�o�C��j�z��V��X�W���j_R�[1-MUU��u�l[�*8n�Zj�ص�wwʶʘ�8����m���{ln'�A�����@]ޥ��[� Uݜ�u���]ٕN����wPP  PVP]�   <  p   �� w �� w���� 6�l  U T 
��x@��9*�����n�k���-t��ou�sw[r֫@�w W��� 6����	 Ò6�nH�)ȹ��{�h�䆆�5��ʯz��k���7�����׃H�8w����m��m"�uhyp��P:P��yθ��-hh���Cj�\��ȤS�;���&9n4����Y��)7{�L҈Ӈn������I�Y��M�Z*��\*T5ة�I��%��H�eȳHgǻU�CCC���W����?�����~�ߒ㍸�mH�n<F����<a�]
P�ռ�R�!cCFP�D><����M.�Q��D������Ա�@USb���TlJ���͹9�M��Hx��4��N�#�9�^k_��U���{J�y�j߆�uZ�!���J�$�F�m�dR5j�5�:��,hk�˨�j_t{ЅFT441��\��A���y��Q1�I��0����:����F���hu���P��������j�ޖ�*'$���hEi��=�2)���o#�^!�:}��L҈�ӷNv	��p�.���i7#I�nH�K�;�xT���R�gnө�uB�e�]E��~{��T441���S3��=��z�qݹu��om�W� *�qT�R�T;��UV�s-�ս�$�$��#��/sۢy�ltzkۗ�N�-{�ܚ=�(C��kLQ)�H�Җ�������+������.�����܏V���˭��D�J7$2A6���*����,����"��s��e!�{շ���l��m�2������J�\/5o|'dX���M�jߞ�����M�D,��D�"R@��8|G���˨t�<4���յ~��T��c֫�eM��^k���_&Si�㑦\�%�E���l��WU a�^� �
��l�z����$m�ܑ����F��L��fv�� �u���uZQ��
r��S�]H�ނ�m�Km�#q�2�/��/ ʆ�lc^d��25��#�Y��i�-ŧ#=6����JEm�[��wP�4?4��س�Z�����CT��E��-s���"FYq6ܒI$0�#�/�t��yidi�ۧ;�Hᧆ���P�gM�!���:moI�ƛq��-D2������*/���v�eCC�1�q��B����i�p۽m�|���ٽJ�*�{k^� *�ت�� UaTVgu�k|�q��)ST��msV�롆E��Z�Ч�|�3ʍ��!kC�Ƨn���΋�Ma!U�7��Koxt�N�#�.�sZ��eM�Z��{J�sX���j,څ#�(G�4�JI$�"O#�[�OT0�z}�^E��i�P���DiçH�'�;�)+6���J��#I6#�ȳOӆn�8)i��dZ0��]
|��c<�ڋ��=y�����e��RH�	C�D4�-�-s����"Ǘ����*lr��v���`�p�¡��-��II�b{�e*�������mR��w �xx�)��k�U7{wx��� �[�������{ .b�Em�;���n�[oo*���9��ٮ�| m��     S` T�  w   
�T 6�VP �`�
���@�  �  �@ *��Um��v��k�F0gv����=�4�����������z�
���R�p��Q��H�޴��!�K�;�X�N�uZY��;��s]P���geE�R�����hv�5�.v�D��HܒF�H�S�!H��ўc5�C�@dK��[笴�L!kW@~:i:�i.��rH�m�܁�R�=b�\��>y�}eK\�=j�3x�O1
GO�w��F��ec\,�dI�$�H�r@�R8i��,څ#:nq����-�'�E=>�/"�C4����d����$�Q��̈�8t�G*�U�d.k�W�V<hv��v��|���"��-j�!����uU5V��n�Wc����ß=�m��6��@W��@w U��V���m�;�Wu6�R�v��g*6����]��4:���:��];��oj�l��e����q�S�sy�y���A[nt��/�B���S���В>Hۍ�#l�����݅�P��kì�^fB���~�cƇn��K��[���,��d�ےH�q`��#&�㦵�GF�_���\Pվy�k��b�:zD�a�'��J���y��k�q�69hz�Tm(�k<}ɨ\�ک�s�e<4���Z�Iq8��B�*okm�����\�
��*��F�UUJ�έ;ۗ�� ꉅ|E�=}�eE�R��Ǜt�lc^d��29�~�_�X��;&e����m��M�Y�Fzw�0t)�5�GF�_�_U�[�ʞz��8#�5$���k�="S�ʛ�sZ��eM�\$����Q|�><6���U!���qT#�D�m�a�!���:e���XE=>�/"�C4����!��ʲUy��1v�D��$���#	�<#N���4��Z�C��]
|��cЋګ�5���G�&BL�A(T��̒���q���u@�w��UWR �������9$��f@�Y�a��X.j��ǭW0ʛ�sZ��eM�Z���`�p��4ˬ��r4��F��r��|��V<|ֺ�U�ms���ʋ��݅�P��j+��bjeDnIM��E62�q
G�����kAu�y���-q�hh!kUB�c�;�^�IH"27���!�2�(x�Z�(jڿE/K\�=j��T�Q�ݻ��K#H��2���D�m��%���ͤ�o,��,��C��{ᗸ�\�s���ېƛm�m��+]۽��o]�.� a�^�U�n�U�g��v��ծ�U~w��X�NSr�_v{�^�YAu�� �'w{��3YB'$�&ۍ���/��*�m��'��z�x6y�ԑ]�ck��8̉8ے6�r=[��/y�^z�*����,�w����W��WD6�%�ܑ�$U^r�n����ixǷ-箌��7r&{�{hz�a��q�ډS5�B���*�`i��'�WI��z�Ѩ$I$����q$�P��������ø���^������ov���z�1��mwR�m�qT7��y�yR��V+-��gl��<�=��vu��uv��{p    �  U�   �  �P   �PU�U �6� � m� @�  @ *�U*�ez��l �U]�w[3,<��ٽ�l�Sd�[=p �ت�� UaTAW���P�t�@rG���.�z�6y�l��$y{���ʅ�������m��J��緛�Us�;�e�m�����:��l���F�Q�fHG����ww,�ۛ���snz�g� �4�ģm��ko/dau3��8��e�h���k�[�sa�<G$P�i%Ĥ�I2D2�0^'v�tR,,�f�֊�g���Ŧi�q�!"��e��#���;��T�S{=�O/T U�<*�Cl E��Ή�m��P[j�)�U��E�)X.0�Է��h�V(:�汞N���k�2�S2�Jm�Br)$� ��D#���dx駤M;��j��X��*lr�5�Ɏך��n�g�	�RH#m��#,�0��sP�Y��;��tR,,�f�֊�<`wT�)�M#�5�&�P6ےH܆#M��[�
�U�ƹ۠V�y���C��H�t?4����X*'$�&ۍ��f��)�7�!��f�G���T0ʛ��k��69k����v����ݻ��T��]7���Tl;�U{)YC��@Uݶ�זm��7�I$�G
G<>��)g�xSfV��,�x��u:)z�m�Ef���tk!D�&���.dDS���uM(X*=��ЫK�u���=t0ȵΟ5�xx��B��&e��wD�ҍ��{��±ifo*y�Q���*Z�=j�Sc���}<�&�s9!1�䌹#�,�z}�]8)i�u	֐`�SfV��,�x��u:(G�s�*H���I#l��G<8�.-(�E�M(X*75�ЫK8wy�A�4�úxq2�i��Lq���������j]@��U@e�ATw[S׵;��ƫ��W]G���+�(Í�]=�zj{5S�F��dt���&�7a�Iq��,��?R8}.�<�dx��	w#=>�)g����2�GJ�^�!L��nI#l��ϙ8{�x���H�;�!aF,�7
pl���p�nؖ���m��mH��#��3N�5
;Tx�f���5I[���΋�/���eB�j6�
<dx���OSc�����*o����L-+~t�x!�a�{����YM0C�H�K�3$�Il�)O/T UUz-���l��l�1D#�H�m�Hm��<4��bR���������[
0�g)�S�����Qr&�fG$�8$c<xG�:t����^t�Pr�|��}ʻb����
���H�m��%�)���g�4��}Z�?<}��4�<zg������V[��i(�Q�I����u:q��r��{���f�������#
7$�&�m53*��R��FM�=r����A�;����~�o:�����,�^
��u^�]ՕT�yø6�WU��p�����ދm.j��*�z�������@C8�k�T7��:��j�N��=��!�[z�� 6�  P
��   �  w   U�T ;�VP �m�T  � ��  *� � PT<
����W-�m�Tp���v��ums��[��l a�U+�J�;�EJ���>V�Bq
�Cr+��Q�UV������:�v;�n��u��D�m��	͝�W����{j1_n���v�.���cDϛm�ܙ�C����T�Oo.�^���r{�JM��RI&$
�N�E���E�U���ڶK�s`з$f)#n6䍴܏� p������ǧ��S�~���
�m(�ī�Z׏F���MT�R��Jw��*���� m�p����
�mYATw[Q�׹�Ԫ�(��<GM[����=?]/���C}Fq����6�������q��e��|�Џm��/E��>�:p�Պ�;]��z~~صF�.4��I$1)&S����w��+���a������F��uӄ{귄�mƒP���#��v��:n�f2:Y��t<s����3�{o���#JE�� s����)��|����yyM����wý�&�l�`���h�q�S^���
��UU�@6Ք��l�dF1m��mĤu��^5�tt�=yx�½�w"�;�O���s�hE|�KR�I$��< /m�3�k^0�"��Z��ܵ���ssZ�֡N�M���rH�M�������v��?<u�2���[\
u�,eE�p��l��"�jF�X�	�T��~O2��Ƽֲ�ʛ�8�]8)|zT��Lh�B[m$�k�����Uŉ>v�*�H��սoHx��;w��������H�[oa�G#�m�ʪ�n�J�ޭm l;�+�J�;��,�S�p%�j�l�(�zf+

��U�U�Pv���q���o3�|FwC���r���D�$�rIrE�G��ۣ��l������c�:G��ܻ����,�Z�)#q)$�8Cp���>��<F���2����c<D#����0>{�0���H�IF�&c#����s��}�3�g��KZ��aw�=j�����m��I(�x�7�w"�#�t��td���McQ�^c^k_���sU^tJ���k���m�M��o��w
�����6Ք*���>6{�r���s%$�G#��1t~��,G"���􎑺njO��n��"��pQ�"�$m�ܑ�s ���v�1����n9ӂ���^�L���^#u�V�M�[m������{h}?^r+�w�tO{��g7�[�LnHۍ$�e�s������������u���=#sJ'rIe����sw=9�y��x�<���mkV��W���>\���*�V�ۻ۷O�8K�  ٭ml�<W^� ��T����9�m�����A9�ol m��=|�^J�m��8Վ�p�_;5E���0  N �7���<�>  �'t@x x>'*��9qղ��P1�p�� �p0'T�� �pଯ݌��;�C��{^��{m���6�mQ�
�pV��w��
��U6@ƫh���m��  ��uݴ[!T*���U^�k�M���O^�N�m��T     mf[�]� 
��*�T� ���*�u�u� ��@  U��UPU �V[�˨
��m�M�z��k5��Z�ۧ�݀������ۓj�kٶ����*��A�c�ꇃlp;��A�w{���l�     .܀   @            �      QT        `                U                  *�  U         � 
�l�Tw    �@   l   �     �P        +u� T    7    -�      � U       Z�                               
�   � �  P� �    *�T      �     *����@    CU���C{`p���  0���(���Xں�'���wwe�� ؠ*�pU�7� <7����[��X뻵��*���m�=��s��1R��͛`�lR�wTܮ�{��.�k�gR�_  
�     6�   x  �@ �� �� 6��U  ` ��` �  � �U� �lR�-����۶��y6��m��Q�ҧ��^o%@U�mT[ j�E�U���6TM�m�����,��#�0��Q�`סEh�^(ŽS�i��r�cP��I$e��t����N�J�s�j;�o�Rh�y����	ĵ�$�%l�d�e"���Ư�SZ���_?���a�rּj�<���x�7��LM7I3#�F1���{W�\h�Wu=4sH�`���E���ï7D��
��!-�H�V?��ꢩ�cXԌ&��sZ�|eN~�{���H����_4��cM�oDꪷG{v�m�d؀�� �ffP� � �n'�j-�eڥ_���k��B�k���r��SZ���~��������F�W�ľQ�$I6�m0��p�F]�0a���i��i�l��y����4�|�FG$p����[���n��~����8t���w\�H�t�.�<����L�-F�$�q�Jp�a�z�O��"���e���P�"��jpl(�kڸprY��RF�³3<#��<p����W��b�yX.4]+���
����n�j�8�|��XyUIݹ�, 6øUZ�*�� U^�˝�o3e1�D�I�R)�h{�f��:xxe���Ϥ�kֵ<���5�k�b|�I$m�ܑ����G�<�аR��or�R�f:�r�uZ-���Vc�#�ƽ+������m�$�'��L��a�rמ5mw��^fB���~�j����u�<F�G�#t�(ۍ�#e��ϙ���P�G�ס܋;P�=9ud��2�5�:t���e��rI$��#�+�R:}˼�?a��n����H��1>g�C�h��!��~���M�1|�I��ܮ�m^�[c��w^�R�*�qUW�ز�ՔG7+3|��UR�Ѣ�c=�0��2x��1t�{�dx��k����5��+��V��o�8%ґ�$��A�p�6�Y�>�"�����;�e�#Ǧ�4�M��5q�m�9�x�!��N�)2��b��E���)h��bޗR�f:�,����"J%$�H$��S��f:�a�]���U?�wި*꧎�P�+/�-"k�I#I6#�F0`�{;�D�.��OIf:�lj��X^�/��<7	޾H�$�2G"e�u��ζ++{k[H��>��+ٙ@w T�*��u�ֵ�v��	�~���v�>?�x�,xމ\�V{��b��Zۺ���ۤƾ*'$���I����ZЃ2��?�����Vן��u��p_r�#Ǆa�7`M�m�"��a`q��њ� wۨ8<F��]ŀ{�p��}#��W<�h�D�m�$
9��t�.��yn�#�k�O�M"!y�zq�6����b)9#q)$�@����>#n���C�r�WoX,����P�î�pJe�M����ކ���/o6�' �85]�C���M�m��ʽ��e{��\û�]�VP��x�oa^��b�*������{���\����wP       �   �  ;�   �UQ�P cl@ �o�~�@� T �P P�B�� m��7{��y�T�͗hUM��f�f a�*��� PU�l�k�.�ک_���۽���Su�Q~�V�*|�Q+�#`�ş3�!�+�4Ή#d�#h�2�O�
�Y�C�x��w&���^��#�v�S�B�Wʘ?kd@ӒRIr30[���_��{�7G8�7lc�����$jI���rF�J[%�۟e�*����=�+��V����\�A{v$��d�ۍ��>g�C�YC�?p/J����ӗVM?S*��4�G�®� I�C�#h���m�MT��8�
��UU�,��ed��%$&�?G#ND�,3O8�#�ܻs�j-v�'���E�z]KI��˻8�R)��K�j'rI$����:�a�U���U:������������#��g�?3��Y!�uF�m��M��
FF���>g�C�YC�?p/J����ӂ�M?SʜѢ"�f5$��#�#���딭B���]�xj/N�E-,�y�-c�ƮA��D�m�D�E��~Ww��#��U���M:�����������Ӭ���������x�����v6ͯ^Sg��T��핔pJ���Ӽ:�&�1�$a�$x0�aݹ�ࢣEһ��i&�
�T`�TZ��z�C�SҦ]�&�*'$���!ȳH��غ�CC�����b������*mC��?n����H�V��f$Ԋ7$(F0i��<FќYH�t���3��dh����­ז�z�ZX�\����	��!-��a!���p����ۚ�
FCӻ�0ڇHw�����Ѳ�rG����3��pZaKz��I����O��0އ�:!H��.�<�xo���G �۾-�;X���`�ª��*�� U]���ލ��j�^�.R�Y����
Ww:�R�WoZQ��\*��?>̲��|�c�G��TD�N%$ma31���O�A����E㴜�(\I9��)`�VF��� ڇ���0�Q8�M')ӆ�o�xt�����S��^(htt��ԧb��^�!�H�mĤ� ���F����pR8i��ՌA�0�5k��W��5��2U�+h~d�><�2#m��rIs)7W��}ۖ��x�,�>�ֻ��V<hw���D��a�҄���	?��8�'������e�P ��+�W��f�m�PU͵�N��޻-��W���^�s���`����£�:���u�q�w��O��.e��4ç�)���e��nJ���.�b�6�y��ʛ�=��Hv���\�C���5���;c];D[�d-��d�[q���p�>7��Ʊ�{йQ�hxǍ�S�!t�,��<#Nug���.5rH�-M)�5lz�h2-�����=Ra�����P�0���r�Q�M��o0��<#|w���4�y�u7�Z��Hv���(�K�\wB������߮��.Ggp���y�S��l�"��'��cN�A8mۻ�{�eOV�^妽�Tǁf�k5z�noR������l���w][:����6��Z�s�P    @�     p  <*U��U�*� �m�T  ��[��  � �U� �ohU�m8�w��������W�����-6*����qܠ������6E��iN��,m� x7���{�/��˅����]�³��j��T��"Ѩ?U����g�i}�I$�$�n�*�X�w�~0Sh_�E�u���A��cT���Z��5��H�&�nH�2�D;��\�ɧ�i�G2�+��>�n���&��D�_�Q9$%��N%s����ql�=�r��f��ӕۛ��%D�˨�n)nH�B�f���7,��͇w{�7qW��=��|��� �2I �H�e�nsqz��wv׫ ��U�
�l�UU]��Z�9]��P=�w����^�!�z�{&S�;�������F�H�JI$�(�[��]�&�1qy�$:�Oq��fPXn�VC�TNIM����y�����ݿ^�YY��*�� �&��WBjө�nf�e�2����ƛh* m׬
6|ʘ�(<@�?�Ω�SUM�DUT��� ��&
���M b��!�x�b���/5�R9��N�����U*m�w^�T;������VPVM���t��md�P���������r��ra�+��,7ƪ�����ʠ���i����m��nI"ů7wܚ([�@߃��4Hau���ӈ�����n)�sL/ݧ���3T��5�&<g
�R\!�\fB���6�#iD�nI$�"7P�|j̲Ʊ�{йQ�hxǍ�S� i>ތ���iέ�#RH�6�m���EUMZ�=~��Y�A�y�jީ0�aZ�\[T5L#H�j��Z��.�����;�ms�U���Ԩ�w W�Sd;�*TN����8cRI$�G�F�t�DZ%�����t�T���Ǖv�-c3�r��.��+�	ŨG$���l�$�f�:V�r��І��������ʏm�C�<h吧�B�k�lu�DE:����uR�x��`4ګCVǯփ"�� !y�5�1�[�t������lI6
��!-�Hr!�D;��\��1�Uɖ��5��{*lr�{���'��OM�q�m�Å�ԊL̺U*���!y�\fB���C.TWt!���e�cR�=�\��ܴ<cƭһ�A��������p�
(�j6+�]��EPm��UUUQ� AW��k��$��i6�˼C�;��<ŏ��Uhj����dZd/4��ӧH�6i�6S�F�6�?4�w�-hzT5l#H�졡��\�n��C^}����-v8��e9�nIM�a7��p�ừ�LŤ!�\^B���C.TW�������!���-���m��Lm��mcA�bhv�mxy
{��CZ�j�J��C���f�[�Z�C��!y�u�!<m�$�D�Q���8t�;D�Û�t�z눸T5l �e�P��Z�&[��ޡ�x�w�(Ċq�R�2\�(�1�u!6�c�<�ly�ֺ����
�cN��o��h-ݵ@�Էw.՝��P kb�lU��-N�תʷz����o;�       �   ¨ p   +�6������
� p �}�  *�    ����J�x+��k�;�Pn���η��;���l�Jn�ewUz.ke����-�S]���Z��� _y�O�|r�
�,��R��}�\+\^B���C.TW������-��6�-��$��!���!D�wxǍxy
}�d!�~5_�X���i�0it��h�����nH�75��Ԛ�ƭ��!kC�*���i}�4:c֣�:��sQ2��F�0��n��4���#�,�=��𝡫c��*���!b�^E�ΑӴM�.#mƒP��.��4����cR�7йQ�hxǍxy
}�d!�~5_�X��ǖԪ����Q3>�r���۹Z�`P�\5@6ø�J�P� �PU;����,�ch�CVǮ�Y6�uB�Pk�c���t��p�z`��%"WM�#�$~�m��měy�S="x�jZ���r�*o���v<��Z�;|r��9�#�&���%�I$H�iät�%ʊ�C\��˒ƥ�k\�ܹk�>|#t�괍#�ϼ	�I���ET�5��;;
�5lz��hwQ�t�x_�4�=򣔎O��-0�ģI��7P��!�]9.M"�i֫����k����ʛ�-sݏ*4V�8t��m�V�[rj(ڒO�mJ�'[ػ�(�w
��Q� 
����޴���L��ߜ��}��k�d+��t2�Ey��z�e�cR�]"���2)ᧄGu��8�m��Q�ST����:�/eX�w���U��:z}�w�6rΫ��a|�6
��"I��Gח�z�+���[e��6r����]��[/F�9i9$�Ϛp`�8tứa�L�H�`��!c�5��\���CC��˒ƥ�o���`�eD�$�q��ɘ��ç�{^B�tYk_�W�V<hw���S�5oOO�n�`�8�P�L���I�����im��m*OY�6�R��UU�s6���m�mT���۟
������߮��o�L!����ŵCT�4������(;�Z��i:�����!�����Hqf���^�B��p��D[�:�CX���c�5��\��t-#O�]] ��⍸ے$�f�����r��r�������CZ�j�J��C��;
v���\y�b*�:���[m��bC�Kź�H{��Ӥa�ɺ��Z��
���i}�4:kѷGd_)$�DKln�u#Ǝ︭[\�#UxZ�5�*���5�w8�iGO�7x�D��b&���%��[�ت�׻�eUa�^�R��� �
�;���k4� 9�����!�4��9�R�w�xK��"��v�A���
GO�Fy�E3�ߩ!kht6ۍ$�m�#�}��K�j!ޗH�C��Ts��ON]X���uwW.}�1#��$lH�����2��ןi쩵s̍U�Qhk�T�4�V�H|�N%�Iq��d�$C4�#���aOy"���)ڹ�<%�q�O�=N ��x�#��������29$p�#0�g�͇��H>�t����K�R!�w*9�H�����}�7��wm�����ʋe/j�Px���;�R��g��-��]�z�1�p�e�Y�����ݞ7����T -:���wd�3��*�5u�w���     P�   �  ;�   ��
��
� F�@ � U�g� 
� 6�@ C� @=V� f�w��;�t��ٶ�*�i�� 6øUW���6�l��m=i�����7��ޣ���=�\�+b7��{�\,7ݗ/"�qtOn��H��W[{���jF�D�84�V��87s�f��t�j�0���O��c��m\���ȧ�a=�Q�ܒI	m��)���4�w�_�Z���GpmU��cR������K�N��n�6JrH�2F��US�!kC�k�j���i}��:c֫�-�ta�ϴ�T����Yz�Q9$I6�m��4�ç��b��B���+��t0�S|F?��s��4�����e�>AGe�XnVU+����`
��UWt[+e����w;��I��-&\&6�n6�B��{���/qa��+ҋ+geP���_�E�3�u��Dp��I"DĊG5���t�$��?;�.[�2�(htǭW&[���ןk�̪�Sm��mFr<���ޯ	{�`�8t��Eʤ:�CX���c�5��Jn���O��+���j6Km��I<�ͅʏm�C�<k��S�!k�~�cƇ{��;CVǯ��⛧-�m���ź��{��Ӥa�U���4?;�.[�3�F�Lx�������Tu��n��쭱�T;�+ԪU� �
��tu�-��nIl�d9���4���#��Cݏ*4�hk��EʬI������L:G~~�69n4����=P������m\���>�ç�{O!O��5��E�U��_�h�-�L@ܑ�$�0it���Kź�H�\�cV�]w�k�~w�\*����zHM�MH��#L:xD�p�takϴ�T���ǩ��-[;���4�[�i�wŖ"ID��IR����t0�S|BƇ�ח%�K�B�G���5��)�A���ߏD����Ϋ�s�z��������<��,�a�*��6UO �ʹ����I#I6�H�i�4�V�w�F:�h!��B֤�#սRa���i��7yL4�i4��H�!�F��g\����-�ф!�>��Sadi�W��аi:x|��|ӊI!3315*���!y�\^B���C�7�,h~}yrX԰��.T{nZ0��`݁6�Q��7!�2��ҵ���
�m�M�v���_���u����Ӥaݜ��H��$�q"[���8F���	�a�]�ˏZ1�U�[��C^}����-v����W���u㥼��U��Jv�7� Clm��f�6Ք���=X��9i9$��Ӂ`�8t��ՌA���./!X��])��^T�;d�`��qF�J6�{�1�7�Ӊ{������X����@Ȯ�h8���6Kq#ٳ�nj6�w�ꐊo�:�gX|����TD��������n��H35O`�0��D����E#:�O���n����L�DUUD)�� 3NT{nL3ø^��mx�@ٳ������O��d����6ܑ�,w�mǻ�  �{m*�@��1T�;iܖn�ۛ������7 c ���+m�ݶz�t��^�P�C��(�ض��p��;������<� � 1�p��y�UBpu[��[ Op�` < < �F}�8:��p��� ���x�N��;��O}���Ƿ��x�ݻ8�Z�m����U�6�.�G b\��خ݀\�6#�몀 J�  ��h*�*T�E@�[z�� N���犠
��U   *�Us��M��� U 
����� Y�T�:�  �� �{��*U �U�� �T���ۼ��nM���z�����v��@ΥI����Q�wy���+ʀ*������@p��߿@6����n@     �@   �         T          *�       U�         *�T >��                   �
�
�           � P�dU <   [`    �   �T     ;�        ,�  @   r�    �       �      C� =Y@� 
�   �       �          T    �    ����  p@      �@ UU    ���  *���mi����     ��
����öw x86�����w�V�pY��^���qY�cZ�;�����fD�������3]E��m��*T�D�V���AR��ٶ n'w���Z��{xn��ť�d{��{vy *�    *�w   � U�  �]ClGp
� 6��@ �M������ m� U*�U 6�z
�8UJ��Um��[۶�K�H�OW�����vM�u�T�w W�T��TWx6��U�T䐆���E�?�#��3N#C�j9HZ����ڡ�a�:��tǍyO�&ܑ�*\9��դx��idv<��E�c>�T�WX�W�4��:fӚDI nI$�Ԑ,�[C�ח%�K�B�G�-�!OtZ�x�B��C܋�k����S.6�R9$p摇OM��`ӑn���t;cV�Oa��hzT5l#H���Y��I$La��%;�z�5��{*lr��cʻE5�x�"-��1n�#�x�"DjBd�BڈFwEV��ԥ�l;�U{%EQ� `tI8c ����m��"I�8t���Jo�Ƈ�ח%�K�B�G�-�O�� �V�i8=�:bfB�P�ꪦ���V;hw�lӱ�c��@�n5�Q�C�5oT�C�#Z�o��B[l�$#4�wW|�s`�Lx�y����������-v<��K4�<0;����$i5#rG"Q����5���V;cZ�a����h~}yrX԰��.T{b����'S?LLRI	m��)��ŤtໞC4�s`4�UcVǯց��qר���C��m����8Ќ�⍴ԑ����� *�ت�Ql���e��w[g��d�m�$nC�n3�WH�ӂ�5CT�4��)���-�фy���y����Ws�-��n$�n6�nC��c��*��� k��vƵ��)M�����䱩a����f*"1$l��m�&,xt��i��o�����V;hw�g`��ձ�0t��n����
�i���$J����8ƭ�I�;և����CV�4��)i�O�;�m\դxޞ������JIS2�f�lr��cʻHv5�x�eʤ;���d+��t0�Sa���omݷ��Ϗ"�-�U,��*���-��z�J���*������#m��n6Ҏf������o��k�<h2����k�����vvL�0��E��\M�rF�%��K�ֺO:��z���kC�\E �;�|�.���8D�i��ˉ��nj��:�a�5��{*lr��cʻHv5�x�"�R\b�fE��ֿ}7���F�Q%�n�����4�a�.T{b���>�2���~C4�s�=�~�Y.5rI�H!�j����:C��#Z��t;cV�I�;և����CV�4�W���(�31U��k��P��7wj�m�p{(
�p m�U����5R�ʈ��:cƫ�n����=�69h{��]���<|r��8���l��-����F�lH�N#�w�v	��ׯ�.K��G7G�-��S�դt�s���:�H�M�$�ӄk����걪c��@�n5�I�C�5oT�C��hz��S3�n�Ù�����4��[��:�C�<j����6��OeM�Z�yQ�;�<q\1D�i�$�6�I���b��GќX;cZ�.
U|E�=}yrX԰�z)�����O[w�(�R9,�\�(ް8C3ݧ�xn4�w�����V���S�c�w71���]�Qr�@�/Of��s���  ��*��;�2��nO,�{.��k׶ʷ�vy�T@    s   �  � *��l �\��w�*�;��m���B�  Tl�� �`g��Nz��*����)u�Vۺ�@2��t *V�UU�EQ����ٝ֨�i{V�JcF܅������87�yӄiΫ9tC�D#`��K�꺯j5���ca#�D�m�ؑ�v���г�緛����2��c���=�c���g��T%�7�I$�G�G��R����b�2�|�0a���1����.�ͫ�W3�����D�m��&,CC���S��#��k��,v��c�8P���-0R�Z�C�A��M�[�%�"�wQ���4��"H�����CCƧYn�A��y�B���ۺ����/S�+�΍����WB m���J�UwPTN�=��ż��D�m�����^{��#�a��!R�b�fE�|�0a����cH���d,M�rD�Q̤3j��ش4;h�;�29�v�_��m:�r��4�F�ZRzٍ�#d��NT*�hsp�t�t��T�θua���[��ae!��^^1��U5M��m�ˇ6��R<owܙ���^t�|�5o��J�:���d+T��{�4�P��I$��7W�.eI|Ծ���
�lZ
�������������w���۪;�V��m�n�^n{[mP�� �e p m����	��m�m�n},�=��;�h��0CH���G7WH���FWj���;�F�IS���:w�XG5��{*�rVz�_5�[�t��1]ZB��Zđ�m���B0G�cJo�Ɔ�j_to�
�j��i�6��Y��Ӟ�14�)$̎IH�N�:�.����񂗊��<��!�D����4�Y�k�rHKm�"�f����.n1H�|7�W��r�fiDi��7�,������~Un���^�����-���� *�ت��*��mYAT[;����6�n�MHܑȔc����{�`��p��������d�s�3�/y}�F�BwN�����i6��՝_p���,ӄiΫ˿9�"�o��V���L��m����J6ےH܄C����H�BR0���\��"�!��2�^��}�ݙ���[����TNIM��9"9�}�AL�j���3��i��z��H�HG�]�����ڍ��6��f
~d[yՕ}�m���q{n�����M񂗋�_{����mm]}�֪ݫ�o��'ymq� C��T��T�]�]�o@�N)$��m6y�!�h��#�Wԋ�E)}��.\b������}��������6�nL�y��v#�a���� �b���+�F}�8m7y�WԍOq�d`�l��rIo<B>�̈́*ܥ����Sy��-���C��˿9�"i�����m�a�����_U�0C�!��	˫�!�Q	�0���\��"�!�ZIDۑ��m�!�C�˽_t���3J#Ox���g�D=���3��()�;@:86H�ٱz�6��Ϙ�)���rw��8ClF����E�^m���� ;���or�������  6u�C�����wWy�q������nk�U�͵ �  
�   m� *�  �T  ^��
��
� F�   m�lU��*�� 
�J��x-���l��]�۽���Ǫk۽�-�k7�����ª�� �m��l�$$��n4�� ܁�/��G�<C>���;�)�/�ά��;w�4�s�=�腴�j�$Z�,��4�L�V���L��{D�˫�!�Q	H��/yno�I$z�n6�R$�im��-׶���;J��C܎�g�E�mC�ykS1Z���GZ�%�I$6�a�>�� yu}�W#���˾CD� �S��:�;���5�$���d�$[6ro�"�{��w�>�k<=�����X䑗�	"��Xq(���R;m�� ClUU�EQ����m��T��Za��&��I$&(��s��x���g��g��������D<�v@��8���d99�u}�D�?a�>݁���H�G��=��P�/ �S��F�j�E����yg�0z�i�L�w�>dC����^��z_!��]��#`���$�n7 �Fsut�!�U
���Fz�CC�<�tlk���W��?;��o�����*x)���o��5o��M!��@�"�!�l��R���F�fG��>��U��S�����S�o�g��
��YN�PT;�+ԪUWu 6����W{����U�S3�?�lA�߹��vun�;����3ׇ�$��m��I(���=��T;ֆ��P��~�{`,�4?�^�7�z�G�|��n&rH�m��NL����Z3{�G��V�4�T+H��1A��;M�˫�is���o$m�����s>G�\�&�pi~�y�2<ֻ\_����b�:橫}�����q��m�$����qn��f��O�{���w�kC\b�U�?z3�R����q6ah�ڎ"�2F��4�omM�b�޻n�m��� ����p ��ܑ���ZN�.ux����c�{�ܬ�Q|�5o��M!��@� LPi��ҌmĠnI$�c��#꺒�����CC��>eƑÂ�j�?i��"�m��q�ڑ8)�5-[�lC��Z�k�O�{������]	�==;��jjdnI$�H�\�<jN����X��|�v�Tv,�#��X�Ni���=�H�J6�&�a�7N�#�p�G�ǹHgǤhy���Nn �a�k�ԫ�H��ᕠV�*����o[�T6�U]�TUaT-��m���N�G$�$YNOLۿM!���n�C��Z�k�O�S��
V<k�rr��Q9$%�̌D3H���,�x�<��/Ο���ܫ�s�r�j/�cV�Z���e%��$1(�8i�r�)�c�T��k�T��K�ք�w"�!?S��8��D�M�3�?5n��"��\��PԵo)x*o]�x_��O�l���'��a8�{�5gz����+�������SeӔﻼ�wv;�f�m�Tx]��\�U��=����<M튣�fx6	�w��S����[	TwU��;�m���[  �ԨVڝ��w;��wxn�[��{=]��n܀m�   P �   yT  �U  �
��m���b��l Pp 6�ت 6��0�P 6��x �m�<��ss^��{{"���j� �F�O2�T��T�R�T;��UWv��7f�mT�������s��|Q��J�<��Yܻ�b�����!��zoF��m�$l��o)L���C��\)�<��z�"Ǎ^��D�9r��������CW@�NII(�M���}�7`��:F�wBi|}՞���E<#�[Ş3�x��i��Fm��F�ɹ3J#NSF�;���wA*���B��C�X��G�W�F�����nI*"f����U����)�<�Ã���N��[�)��r����,���-s]m�[��*����e ��
�P w ڨ;�e�ڻ��Saa�X4�ڼ~�{>!�tM�3ut�=`�&����Y��>8Eﲒ�L�a�ےH�qg���۽ɔ�)��ޗ+Rv��)ZQ��5.SR��Y�Rv9n4��4��~�^�!��B��s���
|�4�iDX�zf�F��q��HۉO�i�a]>ݎ���G��&ҧ��+���R!PFu]�%-L�6�m��Q��
p��2/β<��m���rmC�������<Қ\FD�6��q��R74U�����sUw@
�l*��*��\-Pm%�H��)=�N�G�f�M{W�΍���h����U�����$���d�$Y����t�4�0��"���G��&ҧ��U+��|Ki����I$��C4�>=��^)���9E�Y�8�@��re(�p�3{��>�P�|�qI$%��N(�
pڼ��*�C�X�a�7�/U_5/�6����S�f�	��Q��Q�!�ZU>	JΞzⅧ���<�ʇ�;�0ig�x�f�|C>�Q���(�~��mvV檎��<�T;��z�J���T[���{�A��6�rA�WO���Bi|y��^9���;E�Y�8�@��re(�p�7���H�JI$�r�?w�tANU?`�!��|0ʛ�/M_5/�6=ש����D�m���3�L#��ƈ�J��E��箽�QC�[�O���j��^�8u����Dǂ�|Ot���is��Q����Ĳ�[�Y�8�@��4�F�I�䌹%h�Ҍ�=�OX2���R��5�j\����8n��G�����VJd��{�-tm�[��ۮݽ�yZ 6ø�� �m�����V�UJ�^�SW�K�݁����:k��S�\y�Zɫ4��ze��M?7�������m�$�X4�ڼ~�{>!�{Vlup��V�g����::=Ixdr6�Q�3
f��~��n��xReCҏ0]^��@��e�4�.%�I$��~�o��:=�y������w�ފ�my��m�(ۍ�ԍ���#�����ig�^m}��+:5���CV���q���[m#�4�p�'�U��{�����R��V� <s��nӻ�bv�M٠],���n�� �,� �n�T1��m���On���wn�>^ٵ�u<� U      �   �  ;�   <� n!s ��
�� � � 6� P �p>�B���x �*�^��y��g���r��+*�nV��{M�@U�UWt �6¨*���R��\P+ڷ�������ϏXM�	gw�i�Or��r�M�w)Zp�����k���m�C	��#ӻ��\?I\���9n��>�WH��\ ��29$p"��Ǡ}45���hx��H�+�j�AmC��Ll�B[l�YH�ӻvR���~�E묏���Zmy�<�G>��7[-�ƓR7$����L>�O�F���<�����:B<<��:�Ď���7��B8���Y�&�E�z��vz�PT;���U� �n�Ԇ6N)$���I��t�/����ҡag�xQ,�h��ř��?\�����%�bm�$��D1�3j�\���=et��V��z�m�{��i�O�*e�*'$�&ۍ�\����� ��Π �I���o#�y��s�#Ü^����7$n%$m����C�d��tO��)a��Rd�z���rؒ7%I!jg�!��ve�>��T�a��Vm�B9G�Vt���je��o\"�*�m�Wg��͚�J� ��
�R��
���e۷tG�wT����#�h�`Y��;�A�z���p���a�6�<�\?
�=ȋq�!1��$�R��!�sw̎x�M�:~��U��������tv���[mƣm�Kr<Y����7����5f�������H���/r�C��z�Η-��nI$�D#�<y�x�����H�9N����.Yܥi&c�ԹUKxTg��	���q��e�t��u�����<�̎t'������۫W���0|�fSm�z�Nol�yڨ
��*�� �6¨*����ڜ���"I���#��}��i��������P���M��A65���q�ڈc���m�"��B7E���=�̘�x���t�`���R��ǆݓ��D:]JI$��ϼF�w��N�_��!�',"9��< N��#�9$�$�p�#�����H���v<Yׯ����'/�V�^?�O�UK����&��IpH�i>8}�$ t���z�L�멬XQ�ʽ3K������]��4�y�=�����]�k�wT U�<-����
���.���|TNI	m�p`����ѐi�|0ʛ:1��4I|Կ<�B��s��f�	��Q��Q��k)�C��=�V�篬�CJ�c�T���^j:���e_n�Ll���$�n6�rA��/u�%X�?=��vM|���ݑ~yk�n�&R����"��"����I&I��zX%'aܥiF��Ժ��q������/M_5/�6=ױ)�.)9$I6�o3��CL"�P~;���v��3O���O���>��,�=3�{����{6����o��l�1���=����
�3cϸٛg�6f��flfyz8ff7��s�~��6u�6fo�?��~^������C�o��?���������l�|�_o���/�`�����1���������ߋ������1����?���z?/?$��{��^����{���]�ͳ��fm���Ͷ&3�Ff�o��z>�s��1��_�{�g���~��~�Y�6?��������y����?����>?�`�ýO�y����{����1����|~?������zVE2d�$̒�O����J.?;�X�&����ca�_�ῷ��ca��ޝއ=^���>^���1��}���1���~�+��N��//�Eآ����_�S2I2L�*��������}��o����>�l>O?�yy�{6~?�����������e5�2ś06��� ?�s�m������ @                     ��           >�   �J�@                       �        �� � � � `	 $ ���  @� ��ڼl����P(� .���c  �7@ �iAV3@ V3@'�          r�(� ������P��E= ꩍ�15C!�kחT�� i�\f�Ucwk��W��J1��(� R�X�U:������v5Ū
� u���v�s��J�6P�܇]��           c�+�0�څ,`j�  �Uv�m:�mE,cJ��-
�� ��caz��Ucg�I��V  �Icj�U��=n0h1   	�cz:MPb�^��z`        � gT,mOq��ڷE-, �Uhc�k�E�U��U+� ���mULmB�.����J� n��8�Pgp�qj���zN  @r2нe�Ъ�ڥUb�*� �*�      �eUq�u*��U�\n�U��n��� ��bӦ� @@ ��AB!�Ӑ��thb� ��T� 2 D�;
c`_  � �? �*��@ �dѠ S����E z�M    JH�&� ��a4#M4h�&��M<�T����jT�@z�4�4h4�AO�$����di��i� #���T� �   �NwU����w^<x��.�8���"�#�y�Eܛ�T�j���H����~_�
ڢ(f|3?m�"�,��%*C���g��ɤ
O���4�ۏ�s����<l������HsB������(��x�!A�W���Q
�Sld�V����eR�-eX�	&��m�l�X%3|�YP-�Um�e+lB��"m�X�F��T6�e�[`5�I�)S|��7ư��k!Mb�R�X�&���Kl�Y-a�F���� ���T�T5��Sl���J��ԡm�Y��m��B�&�)kإ[䣘�Q].�[s��WW�˳�=m�mlF��Xѣch��8��4UL�TMI&�ElV�(��5T�	BQKCQ��(H�5��������(JD�����"`�#Z�MM4M24˥4�BP�%"P�)BP�%"R�JR�BP�
R%"P��BP��	BP��@	JR%	BR%P�)BR:t4%P�4�LPLSKJ��"ЈR%�% %	BR�% 	BiM"P�%"P�%�%	BR�BP��)H� iBP�
PBP)@%�B-%#��hZ"GBP���@�h]	�֑4��H� .���B�UJSlш�m��M1����J*���I�)�"*���*J��"(J������X�X���MT����ГT����U��&����Ӗ�����&����R(����b"h�mb�m�T4�6lZ�b�֘f
jb�����j(�������HF��F4��MERLPDTAAAL;(�*�H*HvUCD�MM[�����E�5��f#1I14S5MLĕX�*m�QTD�h��b"(���I��j�)����*f(+clh֦b�"���E�M����X�AV��LD�����F�m1ZJ���[kZ-�ֱ�4:t%��Ȕ����Z���:DhP�FBle"
���	@�@�@	BP�	BP�%	BP�%	BD%	�(M	�4%	BhLBP�%	BhM	BP�$BP�%	BP�%	BP�	BP�%	BP�%	BD%	BP�%	BP�%	�%	BP�%	BP�$BP�%	BhM	BhM	�M	BP�%	BP�&�J��4&��(J��J��(J�F�րք��F�К��6�j�t�:Z��;d4%�lIZA�+�Ka4�t6LN��6D�6t%	BP�$BP�%	BP�%	BP�	BP�%	BhM	BP�a(J��)��%	BD%	BQ����4�:Z$�hJ4���(J�N��J��(J��(J!(J�ҥ*�hLM
��T��QJUhZK��T�L:ӥ�U�HbBP�%	BhLBPД%	BhJ�Ж�hM	�4&��4&�Лa(JBhM	BhM	BD&��&�КBP�iv�P��КBhJBb1F	JhJDД%	�(M:BR�ѥ�)����	BP�BV�Д�J*����%:Bh4�IA�-��"�BhJBhJ��l�BhJcmDBRPĕSMb�*��)-"iB�)*�(��cX���V�6�6�[.���ˣBR���%-[	l��F��mI�*��$�*ر��H�!h����E�:�%Qk%1�D���j6Km!�T�m�4�5&��5E����E�S&�8#8Ѣ��k1�%6�-���@�t��E�)Z h(Z
@Ӡi��(�cBP�-	BP�	BP�%	BP�%	BD%	BQV�hJ��J��(J��4&��M	�(JBh+k	Bm�КH�&��(M	���ډ�P�AN�&��(M	�-��1%��(J�Д&!(JH�$�hJ��6Ω4�р�&u�����Z��H��(J@��H�КH�&��J!4&��(M	�(J��	�H��H�%	2�Д%!!���(J��(H��(J��(J��"1��(J��(J��J��(J��(J!(M	�EHi��(H��)4��(J��"M��K�(J��K�ClU�6gF�-�4X���ӗI�kIƊ�-�AE,UKTk�#ZF���Bi�К)t%	l%	A3��M"hM	�4&ڀӪ!�6��4��Д&��J��(M)E�[���l&��)44�ږ��i(
�%	A�Д&��6�Q�tm��Bh��(J�Д%	�Z��(M	�JBP�%	�(JBb�*\T&�Д&��(H��)��M	�(tКBm��(M	�Bi��h6�P��Д&��)�kBP�&�Д&��4%	BP���4&��Bi�4&�����(Jl%	BP�&�Д&��"�К��(Kd(1���6(�J� �l��)� i "�bm�M�Z
h�F���J�h�t�i]S�t�"D�T���4�%�(&���Z(��u�q4�b�B�Fȴ�J4��P�Sm��h�--�(
���4�˵���"h�@�5������8���U�qh�bb�F�Q� �
C@R�U	T�T�TT�QTΓkSDU	٬���"J	��#ANg`��*`����c��Bm���KIb���)X��:Q"�IDN����
6�S�J�A�%i�̵M$TRR�І��4UV�ƴN�U�բ�J*����%X�&
B-%"���Z��I�6��D��E"R%1TE6�,�P�Bb �*ll�\՚�Ubͪ�Q9�h����M[8���Q��c`�X��l�#j-m�9"�&"���h��'C�N�BX��Ϊ���R		�*#Y)�ƒ��QVډ����PQ�5��Dm��٠�ؤ���`�L5��j�j"v��f�F
&H�**�� ���*��
$���H�`4U�A��N��Q$"Q����䲯&Fr�4*��)�z ��_�[�����ce�e��ۻ��[[�L/����틴���/ᔘ���Vo��%�?����1�ґ�e�:��W������;i   �e��,��    ���^��ӷy��*� 8p     �   ��      �`  �1�p�     '     p    �}    x  ' c   	��    x �`  ` 0�*�TZ� ��n+bC*� m�=P�V0*�� N ����  ��8   < <      �  c��P  N    �        �� '      N ����   ����` ���   	�    Op�` ��  ��y�   �z�X�8J� *��]Pp�����50    ' c ��� ��m� x�'Z` m���W)C����p5P x x  cU ��z���w6ͮ�u����]�ݴ�*�6l�7�
���m��������펷j*��YJ��vMz� 
�*�@����P<���s�ٷ�ϙ� ۜ��+���0�����d6t[@�<���5�����뵵OZ�S����^��:��Ww77��b孅N�˽��Wsݸ��.Om��̨�����m͵r�{���ow�����*��כf,�m-ٕ�Wv���Sm؀� �   U� �.n������ �evh  N
� 6�e�i�7y�O*Ux x8}����T�����< �;�`"� �� ��  �_U_k(�� ݋l��ꊢ�U� �[�� �[n�wuv�j�ݷn�R���zb��ER�]aYW��d�L�uۺx���V�ku�gz������7-r�`�[����/[��]�z��+�s�+;(�  O' c��P  N ��Ux �0 Ψ8E^����Tct� �uJ� ���ꀜi�p�� <�q��	�ʧ/Y,��ܣ�Z�QTb��8t���wx�3�۬ ����0�`��Gms<�2�z�yֳw�Z����{�7jחu��k���2���l���vy�j�V�]v��ӷ������w!R)ka�+,���U�um����PPu��7\ۺwv�]j)֠-��!f[5�F��S��7kP5�孞�ogws�v��U�����Z�b��T
��   '-���[al��U�=�.nךk��*�ױt��M[����6��
�x�_U@�����W�  7;���  ����m�ʨ
�R�m�wVR����� �[��l�M��̢�sE�¢�WmiTAu=�Ǯ�w�n����in���T�aCwm9�� ����a���+������ݺ�� �U�;��e����U/Ov/wcv��wO{9u���L��޽��L���V�[m�VR��ڕ�M��闶�b��C��w�jӅ[��۝֣�eT*��d��ԪYk��mTض���[��\��Zgq��G�v�v�U���;c]uQ��;�f�T*���S��� �� ��3���j�l���m*��mm��ج�d��SlQU�$ܜ�:����ܻ�U�]����J�ܫK]��4�������V[�[m�9��]ޫ<��{m��;s]��y�y�ܚ�:ݺ����]�m��(�2��ԖB5�:o4��9�d����ܭrܸދt��u�ݞ�K5�b��[˹zڋ�����*Q]N�A��n�ݲ����pfZv6ծ��+�ݮ�i�y4۩�Y�vZ�A��nH��Z�#G,ݳ�{u�}���u*�l�[�m�U�b���$	t4��[�h�K��������+7Y�陕o�A6r׬`+�m��?\{�n���77{��w��i�Ƕ�����ʜ�j�y�-޻1�̯r���y��6n]ex�6��׵Ӵ�y�����������
��1��/l��R{�%*���a�.ZFS�\�l�^���V�u��9݀d�ݺv
�P֔�׶�s���mif�wU9�[v�����j����6��]�6V��v�[g9M�Y�u��V�n�k�n�*��s^�i�) ܁%˦��[�Q�,�%ZXٜf�yWum���ٳ��ڀ Z��nяu�ǭ�����6�z;�5��n���ܽ�7o^�۹+���hc                                                  �>�                                                                            �}                   P                              P@� *T     ��T*��U*  n�T� ���  T m�� s                                      �    C�  ��   � � 
� �       @                 �  U   
���     +���P�          *�                                      �>�   
�             � <          �  PP  	� 
�       T  �� �8�J�  @?A�U ج�        U �    �6�*��  �  U  �  *���N��m��l��U  �pl�� 
�-ֳ�ۺ��-ܫ�\�T��״���                    �                                �               �P         U*�     ��     �`     ^��� �x ���  �l�     �	�  �     �                  W��  � �   ?U}�      �                      �                            VUP 	�       ?U}�         � 
�     U
�V�;���-�>m3*�� }W�� *�     w
l <      U �@
��              ��)� *�    �*�l� @
�  U     *�m�
�T @     ��    R�                 ��           U    T        P  0  @          ��         �              �  �                          *���               *�l     T          ��                ˔  @      U,� z��R�  C�                    lT��VP �@��@ �  �U   @*���     *�u`  �   U >��
�de�d+(     �+-����.`�[i�½*:��v9w� 6ʠ U� �� U U �]z�Å8�;��lUl�� ͰU75* T 6� T    �)�PA��8oM�˛�[�՘����6z�L�� <  1���ûud�m��ms,�ٷ���lWqT +��wm����>��=�[�ͳ}�����~�b�RX��}����~��C|��\u����ڗ*O����;����_������u;[9��@x��oG��   	����� *�*����	�  	¨��  � �  ����   
�<�*� 
�Z��� ��6Ԫmi*q�*����U��^��kím��Z�3�l��n�7Y��[=@z�C���� x�' c\'���R���R�ݽ��p����wt�k(�z�����%T�W��Ob�� @��ڥk����v�s��m�=�`�|Cmfm[�v%6�w�{';n�mwJ��*�mĺ���e[�p��)��,�&�����r���-�*�C]@��c-�vw��UE�\�Dꫛj<̓��[ͦ��z׮ս�Z.[��Ҫ�e���o[V��[�����ދ����eo9�ku�E�[s�����ds��W���JU]{�u;�5�*��ۼww^�3m�7���ս�����<         T              T            *���6�*��       � �  U     U��P          �   �   p P�U  *�6�P ؠ �w����        w   �    ���� 8     @ @*�         � U   ws�Ъ -�P   �T      T       @P              �  P  l�  �  e
�   *�� @� U 
�p� *�u+̀[ ����@Vڀ 5mR�� 4�scuf �'_|>����$��iy���$n��A8�   ���)n�]��S.ٲ۞�i�6�GO8z��xR�S����ݵ���wl�tu��('|wm��ۼl�[λj�6� P  U  .m� ���p 
����rp*����� 6  U�̠ .` � P *��ld����6�F��=���U��w��k{{��%+
#$I$��$�%2J���UU���{�[�^��!{"�גU�fcC$�5���=Y��[��m��
JI"I��@�W��O�A{{Fb��k6�*Y���[�����6�m��RH�����08m���ZsZ�9�鍯ey��5������m�[m��MĽ�ڿ<�[[v��|ѵYG�/c�Y�n��f=Ă�Fۍ��i�k��n�W��A�[�/oh�-�MfօK7eϲf�$�m[U�J��l����: �6�U�t �7PUT�]e^.�n����q&܁�y{�}Q�~ֱ�LnVQͥ�5���n���W�5,�pĤm��h�ٷ�j�{e�~yz���n��F�e���f��-A��a8�m�����V�G����G���,�o����h��k'�[$X���m��I����nn,�þ��?kXɦ7++�Ӛ��Y��K�$�)$�D\q���{EM��n��j��|v��n-�F�ef���H��=ީ��+�w�S�u C��T � 
�[ouk��ޮ��m��Cr�S݉���ͨ�f��G��g[pn��xUk�9"I�ԍ�2kU{Z�f켭ۍ[/p�<�V�&�ܬ�[ORD��2I$%$�n[�v��:��[�f�{�+}K=-���յ�~t����$��8�i�-�Q�רlz�v'�3�6�ջ�n�W��l$�&$�$�r@XNA�{G)h��<[Z�f�V��q���G��՛rI$��hF]�Q�IR$U�v�?�� ��
�P x����um���*l&�!����;7N��9Z-�g��[�w¶�{mU�f��
-��$�n4S�kn��AuYF{6!�Z�v7�3�6��g|�"��m�%�a7W��9��36m��Fm*ͭT�v^V��q���5�\�IFFܐ2�c�g��e��u������V�ǾH-l*m�m��nF��_�V����9��]d/ٱ�Ż�c�y��$�$�&[�\���og{�V�����\ 6øUU *��TE�͹Q��־X��U�,�n�G1�<q���ø�{j�mj���KRn�n6�j4܎�^�ۨ�<[��{�,֣[�V��P��zd�[�.�m� KVm୔����+VU^/,�O��C�6A�X��[�%��m��j,y~6�ŗ�ۨ�{,�km���qh�Ś�S-+���RI�&�VU�n�w2��G���d�ܬ��t�ɕ���_{�����ߠ` <  �1�p��s�SSގ؜�cw�oU� m�)5���e�I!j���
.YV($�w$�ŻX@�����@J�<��n��w>c       Q�   �P �' x-���UQ������  �@  QT *� ���U C�+u����Zu��}} ս�ݾ&�n���犲���wEꪀ¨+)�U^�{;ww.��*�$������Ö��6����ej�˵���.�yj�.5a��JI$�7#S�ŏ3�f�x���u*�x�+}��Y�d%rI"M(��lW�J?nK�ݸ�e���c�hc&�%eyR���f7��Q�w���t�׳�t�ٻ�Q�Z��K�{{�e�z�1���$�nH�q�f���lCj�n�o&g�ͨ�n�ۥ��{���$�D�I\���m��d��g�Z� ��
�P w T��%$�Br7�IH' [w�r���U�h��-z�dv�^��T{�f�M�(6�$�rB�1���vn�[�fk�6{=���kw¶�{mP��:�(�%��aG�ݭ�~�게�z��ջ���&xVmǫ��@��[�D�mƁN,�e��m��oh��a{h'�[Mf�^V��je�bm@ۍ�rF�-��=[��cr���ӫv��t��g��Y�w`.F�p��.I$�����;�ܧ�t�`�V� U;��*���&��q�[m�!�F��]����۵���]
�3ٱ�իu�y�7O�6�T�n6�!)#ջ�n�W��3��ݽ�7Zȫ6�ћ�s�6�M2�#i&�Q��	��w�ǫVLnVY���mn���Hm{=3PH��cm��j6�͛/Հ훪Y~yz���i���Q��ڭ^ֈ�05
��ܒ8�y2�&mG�w���9��㌭�=����1튳o��I$�$m��3��PF��͛���� U⪧2�� �:��*cm�m��Mo�kҷn;S/p�L��>�����������)B�29#-7��y-�^�ñ�kX/�/V�ݭ��Օ=��A��6�q9�Z�v7�3�f�z�}�n��첰k�7ojc�S�Zr�jF�8��D��꥛��V���w�ǲ�[L1�Y*�f�i/���$%��	�i{h���l�{Y��f�ñ�cX/�/V�����~�u���슽�v��̳ ��
�������ݭ� �e@�NI(�.VQ��ڭ[�ə�+i�[��n����e:(��Bcm�"a�3kh��ϲ*ͭT�v^
ݵu2���ߣ�^,a�a�ۉFۑ�bee��V�����k;l�xv5�k-{5x�Hp�$��q��[[v��w=iVlCf�ݍ�{�v�Ż�XR@Ǭ��1��i�/Vc����;Z���t��2n�t��Dp��-   ]X  ��m�ǂ�Uu��~}�~o�o�=����V�|`�����ڛ�](O�헶��N�ҫ=)�wJ]μrw{����ګ�l��k����U       O   �@ � *�ly�` �T S� 
�/lΕS`` ��T ���*��V�s��
��ݽ�� �֏:��Ӳmmλپ����l;�U]�NଥPV��w���$&6�a�}8��c��/wt�ٙ����:3^l[��-D���MF�.CUo٫kl�=�Q���Ӹ��OOLʹ~!!*6Kl��4�}����z�n�pn�ћ�3=���n��H-F�m��j4܎����G�Aņ6w���ӻG6ڣ���z�g�l� nI"J(�mk�ôב���յ�t���͈miX�da�$�BZQ����]w�뇴�^�� C���qT � 
��Uw^�=��T����w�7jl[�Ǿ��zV`�|������<��?%��m-JI$���^ӛ��f��Z��kӫ4�������kJ#H�3[�_&ܑ%a�#�0�+sS�H��Lô�,�(�~�U�Α��ƥ��|p��jLȪŻ����rAZE�(���>�����6���~�G���V�
E�4B͸�l(ےB[nH
m�<aDQ�h�t�F�Ԇ��Ϗ��\u�QҊ9���4|~��/���W���p��G9��V骽� \ø�� �* �����9q��Q��r���ٙ����83^l݂a�jQE�f��gH�ö�m�E6��ےb��<h����it�7cdx���<+v�iDi8v�9��񳵴���FԊI$�瓣������x���sh��s�ϗ��ᖨ()����P>��Ϳ���U���A�� ��یդN|��=�\�MS�j�͝��\�wj�%�m��՜��ꓙ�ޚ�M�5�VP9
8��<SU�_a�-��L!�FZzq���\J?�r�l����2*<F��]�)&U_9�+����6_I$�$�Cr([���v���w/j׷T 6øn�z���6�l�ե�u�t�ڥ:�����㲧�I���:B{(�FFrp�C#��G�뎅�KCþ�ˑ��q�$m����Gy�pJ��(�T�!��8+VY#K�ί�~g�M�M�d�ےC��En�LަF����p��<E����Ї�(��7����|��q��@�%�{�\J���~玀O$��<7�rt/�aH� ^��(���GJt����/��Ԯ3��i��E�5�~�K*(ےFRN:���{.Pdi[�O�Pa~���Q�!
n�g�Eiѷ$�I%[�ǵ�|�u�|�n�zq�9 C���ދdU�UU�*��m��U*���Uڅ�=��Q����L�?Q�w\�y�������#��߹�Q�W�������Z�L�E��㑺>��>�R��?}�=+쎅��/��s����|�|��G�y�q�'Hw'�aJ�#�w��7(�#�w#�/~d�o���M�m��N����>����U��>�������J�������J<J�#�}����'�r>J7�u�J�#�}�Ԯ��#�m�m�q�q�<#���r;�߸�_=��+쏰��}��䇰�#�/��>s���W���~��#�/�a|��F�y�i�rHKm�ܒ!_|>���i�:�y��9��2?��>��=+쎅��/��s����|�|��G�=7��t/�aJ�#�-�]��w�9�y��9� N     *��U�˻���nK�Uo�m�u�������ۏn����T��^�7���:�
��b�j����q�ޗv�����s��f77+��       [`   <  � 
�1��PU`+(  �P 
�   6¨ �    T��G݊�{�ʥU�����c ��[.ݥyn]�ͽt���>��+� ��AQ޺��pW�m�#rB�o�����~">��������+��(�+�?}�<t�p�u��W��w�Q�W���o�9�_�}g�� ��a�P����Lm��[�Y%j��ҽ����ٵ�%=����H�27$���hUVe��Ό:;��Ox=�4��t�\y��pt�8�F�m�a9�{l�.X����zc���L�=�{*7���c����I$���N���wV�ګ��nV����[�A��/��cm�d�HJ�H!((�7��޻m�y��� 6øUW��*�� ����>5��U���~�_���}�0�*��1B�Ҏ��pa|G�ݩ��3�sEk^�܁%ܒ�.�����v�7�����Վ�e�S�������W/3n��.��ԉv]��\�4Qr��S,}Y6���>\Ps9�)�	9�8��P<��2�g8`����;;tԑ�ܒ����b��s7�t��@�Mӭ]�M�Y��ܮ�)��䅇�q~P=��	�䫒@�IkRK��Ŋ`���~���)�N�VϮ��D>��K<�)�7u���rD�H��zFrI$m#?睺�M��n\/=8 6��[j�[ d�V�u�<��VZ����ｻ��>\�}���)�>�m՜���g9�����9����P+�|���0�H��IwwrIV�ޘ!�1|���n�yH�N�����:b��|��֮���xN������R��w5J.���Z܍�����@�sw�ޘ�L��ݹ|��>]�k>��M蘾�KٲK1N,S������������ۇ:�<'˛F���ŋʛug�u|�9��X��8'3.J�H�r\�I �r�9���r���!�1q;;�w�R,S�}~��:b��|��֮��������� bu^��^˜d�i�� a�^�P��AU���n,�EX�wwvIr�w�qLX�g$,<'$�(^go�1b�!�5߻r���|����4C�1�}�}tʄ����]ܒR�gS���;��:��C��p�T��	��Q���@�1b��M����:�SVsm�6\�]ܖ��n��V���9�8��P=�[��9�:&./0��=����z���:b��}��1Ѳ2]ݫ$�wAmN|�D0N��m���C��䅇���@�g2�zbژ%]��/��{$<���@��)�I$�"�r��e^�ɰl�HumL{�y��׿\�mß)���7�\�@��fͿ����	����j���smlv��ֽY a�*��TS��+ڻH�$�"rH�m���9"�Y���!�J����׌��V8�<x�u��YB��fƤR6Kq$qVj���*i�#H�F3�؅}#26G�>?\�R�6F�-�aF�F�n7�9��6W��(ipѷ�kbp�#kU)�O�C���Ȭ��[���F�rE#e��U�(��B0���ٳ��Q[��O�h��7G�����[l��r@�r��dy��6~��i�ih��؅Yp����0���aH���$�I$�@ x  ' c �*����u귮��Rsl=��zm������M��y�w�-�Y{���͗�v�,����T孛���kH�%�%��\��J-�        �   �  p� �t�ATwB�8 `  �  P T P *�Al�UUn��ʢ��nm��_@s�|�{���z͐��
���W�v��k�;�PuI�:��f�UY&�����x���V����Һ��Y�V�-m�0�G�U)�O�_��e$�*Fڍ�$�G#8D<u#䳻=�&)�ՎeM���)���o8b�'T�ݜh���~�_���6�nw�	�1|��o���"�	�ϵ�L_���u��SD�:�/C�vI����].@����7r�C�������ޘ�)�yM�~�9�)՞�g�]�uL^�wI,�8��	�cOu��IrI$Hǽ1~P>P�͸s������}s�)�ՎeM���)���o8b�(�G����Ii�����m� q�z�w�k� 6ø�R��
��n�rSR�l��$Iwm<��sk{9�☸��6�p�:���{9�����@ꛧZ��4LS��f��!�AR9$��M$u/$wi�g�ǫ����ޘ�)�yM�~�9�)՞�g�]�uL^��7�h[H�jF�1����|Q��Tyu@�B�6�̥8&)���}�ށ�1z�̩�Vp�:��noҥj\n���I$�N���L9�y����P<�˛[��'���Tw��)��>ןkޘ�(P�;"��q�$���:䍔u#i<�tb�i1~S3�yN/�����ы�'<���H��%P`��M� �A5�y��n�ݻ=˟���4 ��USb�uQ�U
�
�wv9�u�Cь���4N���͚�f(�LS��ל<��|�y�p�)�1O�ջ�Wd�H�V��\�5!�7�I!NT��8c��b�I������7g9�)��n��
S��̎��)�}�Ԣ$��wj�%Ɔ[ޞ_���u��R��qg���]�r���7y*�R���׽<�)A��kRK�\n~2[9�>��w�ϥw���c�Ig���J�y\�����v��R��w7�	)����[�%�e��@�yz���o�)��fμ��ײJN��ݩ���˛�g8PqO/�?�_� m��4ݷj���˹h ��U[�+�Puh��u۽٦�\�KaD�p�:����������fj���Y�a]�S�򛜕f)k�3��'��]܁$���ozy~R��M�;��(�V{5�]w��<�\����E�(7����������ۦ����%�%�9�P'��߾�ށ��c�&�������.�@pM���G5@�>]��%��%ܕ%�����8'��̣o�S��Pz�w{�_���u��R���>��^y�d�H�^Kw�j�m6ےF�L7+��Z��͜�
��v���(�i]pPkxkcK8@������wkv�l�NVW����v)����eܪ*l�i��n�\�r�we�d����v��R��>_n�������i6�8'v�QĹ"	4Q��P@A��$m��2��5@�:���9��_.a��xj�qJT��a����3:�w�P��㒉��\ +wwwRK���8���&�J��|�}�g^���J5|$s��b��ufn���(	��۷!r��.I"��"�s�).B�v�r�.�(U�u�b�	���~��@�^�}����\)i��CX->f#jE��k�2�wy�����NԐı-����\m��^{���wy���k�B�(7D���[%�r$э9)��I$+�-�܀ � ���    �  �x  ��*���  � 	�     � ���� �6\i��P *���Q��-����wV��ٺV^�e�{�s��x��;kmmݍ���kb�Ψ W�j�Wp�����+\�eUN��
u�^���w=�^{����mv�p�UA@8@�v�nx6ӂ�=�C"���w3ݜ[������sN����n;��77k���^�Ȩ��*���u�V۝��]��v���.����Gr��ʶշ���u#m��ʹ�:ݙsU[�۲��+*�͔�;3����m���v�mm{]������s��n�^���s.����-��R�n��n�n��/wt܌��3۫�>]�KQܻ�j�mml�_,�ol�^�1w���w���ev���.���ot����{s��[{k�A]�� �MYl��                                   *�P  R� m�        
� U     
�C�z�          T     T   �  �  �@іͥ.��[h   @    �   p     �Y)��       ��       �     U    *�T�p�P
�     @����� VUP �  �                   �   �@  P  l R�    �� 
��TT � �6)e<U�Ϡ5]���] �g^oOd�ʎ=^��֡ϟ����}���ߠ ꡌ  � � �*��m�VڝK��Ԫ�c�'z�R���������}#׭mJ6m-�J��y����M��;qƜ�e�63��{����j�]븹�ՠ         PW�  < J�]��
� �R� �  �T  6� P @ �*�� �+ԩe�zAV9��ܞ�ۻ��vë�uvu ;�l*�uTF� *����76�$�&ے~Ԉ$�F�}���.�=S��Y�V%�����ޞ_��>6o��P1N,�ٷR5u$��I$`��]�I��%Ilk[�1/)A�/8>\P>P�n�9�Pk�8���y]�E�q+K9�F��7$�'$��u.�8'w�8{$Ս!�'7g9�)����s�pL\^a��xb�qO�g4f�wrH\�Sr���/�T�:��.��	՞Ϧ��@꘿)�����8�P>��W-j^KPD�G��٢���$�&I.H�l�(�Vz�gһ�i���͆�f)k��&�^�<��|�y�p�)���o>�rIwwwiz�w���o�͞��{I���w� `�*�쭕S�-��[dݕ!��jn���Տ�&�C��uq@sz�.��ovq���b�]�{9�i	���7�aE,��$��42��W�OU���t�_���u���!�ug=�Z�@☿)��eX`�_(�T���$����%����HxMw�b�Y��~�ޘ!�Y��,�-qLzsx<��|��̓���K���#%�9�pC�}[���@꘽X�	�ep0N�(o^p�ܑi�7~��sTZ:��ZvO�$��6�nw���1|�������������:{���k�߸::��Ǳݼ�{�tu������� m��ݶ�mW�NK���\ c�
�+(�
�S��[�z8~r(܍�$T8�t��Ԩa��x�'�c!��6%m��AְӂU�(����*t�˒K�*�8�t��͎��G��Z�@�4V澒P��V��O�
�P|�r���di�ܶE�Ǐa2n25�><�S#�Dv�&�#�=��&�h�$��)�B��h�Pi�������?]_}���^ϩuy���#�������)i�nHc��̊;��"ΐw;���<d�۬����x{������ǀx[k�H���Wsl����n� a�*��TN�6�T[gwba(X�I$���`��q��B��B�:KdYx�&��x��s(�6@މq���#rI��خ0�"��\�Ѵ��#�z�j�>#�ww�V!�w\M���I"I%�9qG)�j��ǌ�e�0�)�u�h��ǻ�q�j��CX�r7�I!R$�?Y�p�7ˊ0��o��
<3�a�=�l��_Q�g��C���$m��m�ܦF vj�&�?x�*nSC �0�X�,��[y���#�zC����q�j�q�sz��]v����wV�Vʨ�ATU9X�޳ؙ-��	��H�4�+�0�[�\��2�H�	Mˬ�q���� ����D�m��M�@i�wh}%#O\a�x�!G���@�Il�Do.7|E4Ah�q��RKr���σ��da�n�bi�<E��H�0��TC>!�m&[)}��Km��n�q��xْ^���̩�3��8�Pw9�8p�r���������F�m�"nGXh�#Ǉw�Pa[�_IC���0i�Q�w�� C��wO)$�� c   `AJ��i\=��݀�Pm�����'�]����zE�������˧��v�lӶ�Wr�ҕ������_˕?�Z)P�}��T      ڪ�   �  ;� P7Zl�PU`*�`�U  �e  �@P*� @Um^��=U�܀;��f� +�۳R�z�����V�� \ø�J̯�q�*
���2��ݸ��m��@�zD#O��?�]}G����> =�LM4G�����(6w7��A�I�F�MD(i�;��8G��{Vq��m��0�8S���G�xA:yC0�䁘葆��z:�q0I�X)�u.�qx��x����?F����m�$.*��Kg���&L���J�ՠ���\����0�M)$�6�C+�d[��{�+3���Y��ǃ����7���E$�E"ۻ{�j���۞�|]�-��ڻ�U]� �w �+]��_,m��T�$j�zDܺ���{Q~f������`�Q|�n)n&��̥�o������2`=�2�x<ާ�����
19$��ۑ�c�e��cnD7��{�+3���X�w1��R7�I$L(\���.t�\�H��]}ޒ{.�����!Ii(ۍ��rN����v�{o���.[ջ�N�,����I��#m5���u���qԳ��� 
��UZ�UOPUΥ��]��ۺ�~�T����6fQ�Ǩl��t��7�����a2�O�i�"I��2Eմ{��C�<.EE�rڹ]�ɗN��Ƃ�F�n%$��܏G>V�qu'm���ME1��Q�n9uUD�P6�d��r6�n.���������T���>��F��pػ���H9��8�mF��kw���[^�;�����tr׫3f���t=��$�I$B�N2�J6�:�:�y������Vz�J�� AQ�M�A��m�$�������ݺ[YGwC�2��MC7(�c�6e�jD��L���mFb�2�	ͥ���/o����T�OCs��ѧ�:.A!� PF�M�
�B,�����g�t�Ռ�և��Z�<ӥi����Y��Z���q��h��6t���뎴��<pw{VC�3�*�er��i�JsH��,���I|�)/%$�2�q��gH�틧�Q���U���oוǽ��=�����ؚh�|���$��$��-HKH�͕�{�� ��U�(
���@*�	�F� ��nH#m���V����1�Y��c��3���{V3��4��O�V�#Mu�و -&�nHc���#6f��Y�$۬g#ǧz�,�6Wo�+H������E���m��M�(qv��7Ϙ�6x�ˆ�e����c"�>#�=�:Y�9�Z�\��ܒF�-4+�"�ǵ(c:C>2	��Yg��X�ψ�����Gϻ�5$��$�&ۍBӵ���R	J�Yfa�,q��2K����<pwz�q�4��Psh.rI$  \  ��1���)�Z|�ڻ�T=���<wU�j;�<
gjy����Օ�}���^�WiC����̖ܻy�����͵]���yỲ      T�   �  ;�P<
��`�
�� � �l  ^��
�� U@ �  `*��m�E��[� �*V�Gǻv�t�[��{���� �ClUZ�UOS�}��j�W��^�����I
p9%�x�]�ЃO㦈[���G�v�Ä2�a.j�F�|{y$J��[�D�m��%*l��&�8E<�H�4F��'�9�޼�:a�[���$	.��Øada\�U���R	J�Yfa�,a��uw\u�������! ��IM�i�o(G[��	ZE���sP��2!�,r��#�r�C��� ��M�rD�%��H�����~�DC�!tZ���F���!�����E:Ou��$�IFZ��m��m�Zݶ+T C�<�U ;��*��Muv���ꩵUZ����g#
�W�CH�J����0��M9,�Ɋ|ɕZZm���T�֗Hi8;��q�lq�Q�v+#K:T�E�a�!9���Α��Ԛ�2Ln�$�r���!�l�X�����2��N��k�K=hiUf�B��|fo6��m�m����E>9[֨q�܆�x�8YW�����<D:T�Tm�����I=�F#F�p8���6����A���N՝���UI^�x�ȃ5q|�����I �InL��\�lw��������U�F� *�\�jW{��hm�]�!��dg�y/bD0�{V2/S>��u�o���;�f��u�+����8
i3#�B�q
�do,/�SpqYg��X^5��g#uW�*s�r#����p��n7"R6�-��tu�������������{��w��^�u�HP�߽��y���qp~���^]��o��ߧ�S��tã~���b,l���`qx�CHX�jFyu�{�!��3ڲz��!�1�DC��z������$�nIi�k��4�+7Ϙ�:C��I���FY�sV�D8�s�i��]�M�9$�I$����Si/r���篝̀
��*��E�Tw
��m���f�y���6*�.�}��a�!�Y��jji�d�a��<�`u��G��\{�s^;/��CN)$�&ۍ��JE�6V��i\W!�,r��#<�佈i�l�Y��bvE w��D��6���L>!F���kPdiY΢����0qt��޵P�/�Q�w�c)8����m��5���>�<N��B!ҲJB���ji�d�a��=��qt�㷩B�&F�RH��7q�7��}��JE�6V��j��!oW��|����/��8�U��I$�G�u���lv̻�:�j�k��wod� w R�.��x���n�\@e�ү��W�i��!�;�j��F���!��.5&*6!Y�;H��m��j4�T7���0�������U��膑��W�L�]f�4���3GS ?
FܒH�n@�K�4��j���yx�����[Zl��!j��!V�+�"��9%��6ےFԄ�^�,�8tP�Z�E�f���r���[P�5�24���q�7��rzCQ$�nE44�:|f�T7���0���f�:E�~�Wd�r#��\)�TǦ4�g�~v��} �  N ���pIƫڪ�s�AU�i���{�0WU�Uo�6�l��ܶs�\c�xy/n�J���;��[�n���n�=ڤ        �   *�  � T��*�p
� M�     U� �T P   n-Ī"ۭTu��l�|@xv�xݪ��ٶ����m��@l;�[|�S� 6��n?��ۉF�D�d�6x����֚�='m�CD8�T�^�xYҟZf�/���L��%�I���#<��{�!���Ռ��ϭ�!�!8�C�֠�ӝn]�A�� ��n8�q�7���0q�P����ƢC��l�dn�}u��!dq���|�8L%)����ϭM9,��0���6�c5�2<xIڲ!����
���Θ�#@V�ܒ�m��7���,�[�ڮ4t����!�C=�!����m�DC��;󽿯��� J��z�7��w��:|�o]ִl�ح��UGp�
�7���D�EFܒF�,�5��E�X�E��.5&!V!Yg��X:/�a;�i��]�wbE?��D�m�M9{��8�U�r�_��Z^��]	����=b��!-�۬��qx�侮&)2I#Q�T4�:l��"j�i�C:-4FyG��!�C޵ZD���f��q)$��q�)�Dq���XC�}8�CH���|�i�X|9�OW0�3��k^*s�+���[��f���.��G�
�!dC��d4n���SNK$3>!�a֗Hi47��I$�	q�����w/�ӽ�T;���T7t�U���i��U-�/����U'�VFt�4��5�<��C���Q佈a�x�BKn��h��n*�%�/�`��ج��ҵCZ�#J�u�p���,�{��)e��r�kr[��~&����[4Y��)�3���(�Qiz��t$i���LԾ��q��M�it��8w�\uő��Wu?!(24��I�X桨����r,���~�0�n�$���B��k�q�#-3^C��h�p�]�rE~B>/{�\l�兊�]�IqD�j;�z��5��l[@�w W�T� `�;v8�T��Y��!Y��sV�D8���E�7Uy��3���"+<%+�f(i�nU	�J��2LtH�g����it����v�d4C��I��/#K:T�M�k��,�޷d@Jj7m��QHEq���(�^�0�ay=�X��Lא�nZ5�4�q�ӚN��t��w֤���I!n8�q�7��I�8�:t�oZ���_!�l����^�-UW<b��x�6kgy�~"ܐF�i�5�U-5�6-�!�a���OX��X�#Ǥ��,��⻩�	CH���3��I$�H�m��Uh����2ھn�� 
��*�����[��d�We�[Y։F����!Ws�q��_�mt�!��Oj�E�f�NZ!�,�%9�����"I��e4�5ő�QY���gH����V!a�䚰s^4G���3"�:�C`�F�n%$�H��1^"��Ef�fa�v�Tdaӧ�eo\��w���Vm��ai8ܒ$�n6c�A�[G���r���v�M���][�;�K�j,���6Kq��U���ʆ&���9�@�����o��~���%���$�I$���I�!��`A ����N{3�p��r�J��Uὰ	�n�]Zw{�+�!ob�]�9*�NW-{=�e�i�s��8R��S{/]���        \�      �P�TS�Uz���  m�  �
� ` � P
��T T����� �*�� �owUz�f�n�<�^˘ B������ �
����q��Um��T�?!�h�jg$Ű�Ӄw�7��w�Z��l�#���R$ۑ�Ͳ���<2>�G=[Bc��s%�1�c#B�qB�Zn[���fۜ�$X���7΢��uAR=.�I��u#q(�����o�휙T����#M4-SH�����x����M�OȄ�nH�M��,�#�;�q֖G5�����,�Ri=�#��jƎ�^S~��Fې&ZHS��$���y��������;�+�@� `KN�eUa���w���~����뎴��K#ވ�4t���+\k��0�����:Vk��+U��r*�7C����+z��O
�4���4��.����+܇��V�ssH�^/Uf����IrI$A�
Ӧ�������2<zN۬��qx�r�b�24��IdA���B�Oy2��ġ�9$2Ghd8Y��%�CH���u����yp6�"!�!tZ��kPf���r��Fْ6T��+������L��Q��c��8�j!�;�6�F�I\�z!�8٦z�FےI"2H[(ۉ�Z�.�tx��m��]ʨ��
���e��.�I"��we�!�+�p�;�%���$����xIڲ#yx�����Y�g��PvB�䐖�l$ȡ��_!d*�v�q��W�mt��/'��i���m�DC�C�G�0Ð��H܍E5��E�\�#!�\jLTlB3,�����\���f�:E��v��6�$�q��b��x�6WY\�Qiz��\di��M�X�b�v��Hqx��s�)F�I#%�t4�:l��"�5D4��
Ր�dg�\��"X����%�/ʆ��I$��a��|�z���׳ܽ�T;�7�U ;��W�*;ӱ��{m���>�z0��ڇ!�A��s�J���Pu7GN���T7���0��
@����&�m�٭4t���y���a��v�F���ji�d�:GI6�c5�3�oO41$�Iq�)��K#5x������4vNbb��(���"ydY�K�u��o�m�ۑ2qW-i~Cވ��!{W.5��X~��4�^����֟�a77����H-��o+��Lk�M���7y��臏�dب�#13MM9!?q�d{~�$�H��ې��'��֝��l�]���� �� �Q�
�(Kl(�n6�Q����CO��ꎴ�3W�{��J~�EwQ{�Y
����GH�]{�I'ѹm��l�^�(�����u�TZ_��7�?C�H~�]9��X~��4�^��7D{P�nIR8n����޵C5x�Cw=l�dn*|�X�D<~�2	J����o5�%5"z*���+ۻۧZ]!��ޥZl���s�����]�D���Eo%V�m�$m��)D�4t����Q�um�i֗��������7�o�������|{���8��}��m���ì��S-��    �x��1�     c ���<��p0    '    N p0 �   c <m� P
�U�J�TZ�om��]ԷM�ۻ+(*�mu���n��m)����q�ݵM���z���� �aWD*���P ��w �[��*��v���:����|�6kk�p0W�]C�A8 :�ⷔ< s᛫�N�{:��a����� 
������J�;���7{ȩ\�U��f�YZɕs�
����8�گG{�U���wR���j�Mݱ�����ީ����w-�����ol*�jb֭uݬm����x��v�y�z�&@m��{�2wwn��9Zê��o�y��w�lv���X���m���w�x����Sa�ݹ�;M=���ݾ6�o�融Νֶ�f��޽ލ�                                   m� T�Te;�          �     P    �       �     < @   *�  
�  �  n�6@� ��ص�   
�    w   �@     *l�    �  a�       
�           
�*�  P  �  
� �   �   d P          T�     =�    �  �  �  �    J� U x   ��
���kKm�q���� m݂��+(-3B� 6��Υ:�U�S����ׯ�8   < < � �v�lL�֛[T^��^�[��Sb�Ur��㸼�<�n���)i[�un��u�Umۻ�u�W�rr��]V�      Y]�   x  p  <c�UQ� U F�   x @
� T P
�UP-�ʥS�zm�<𮯛� ��W�����f���]@JTUU *�*��m�V=��n���M)$�#�{���X_N���:roZ��_��0���Ət��v1^�<~�3��%�$fH�M�Y�"�i~]5Ac,�'��d5���I�XΑ�x����?i��!�Q6�i5"���3W��d*�v��"��k����0�U�KZ_�7��:G�y�ݡNIM�$(��.֟��|�q�3V�����:^�T3W�Մl����v�rG�T%��JI$'�r�l��Q�Fb`�SNAa�a�$���-#�vZ����\��I#a��E	�E�W�����y�onz -��TJ��TJ�#���A��ā�z�o��[�f�KfU_��]n�uǊ�>C^Ȥm��m�����O��v*e����o��L���ͥ�k|�e�� ��$�rIg&U/b�1{zimjgdŚ*nn�Mځ╳�B�IH�JIa7�m���=���Y�cq���v�u<�i�j$�%�ܐ0j�ug��.K��[P�5��3��1\l����iϡ��;�I$��@����!	j�JU$B� �wK( ;�l*�:��9Y[Yy7���}���4p���Wc�_q���"iKŶk�(�����X�p��-�Q����H>��\l���r~�Pp�]�1�Z^��i�H���m��ےF�fJ� 8�z]��%��yz}Ǝ!v�|k�����+������tm���i%��6}�֨o/�}fa��]��N����H�J��f4���Rmģm�S����;�=Sw�ݕ#�g]L.��=�f����t�I$�HE�6�m휴�ٗu��v ���*��Gp�
��6���޾iޛ\A�5jc��s�=��5���jd���Ǖn��z} 1�$F&�RG�6C��A2���,�9��ƢC��l��.��]�W���:�B�$ԁ�#R�q�v��Uf�4���4Wu�Zj!�x�v\uő��Sл�*E�6{{�#p�rHKm�����|���Y�FyG��!�C��i�FZӾ��i7}4x��.=0�nI#���P��iVo�1\l����F�,��9���Q"��a#3_���~ ys���uv�]��λ��m�� 
��T۹+2�r�
���n]
ܒ$�nH�q��!�8�;�H�X^.�[	F�#&����0��]q�7��\����q)$�DЎ@�aE������B���P��K�v^�diۥZD���v�W�|�RI"I��TS���8����q�.��4���Y�b\j	�V!G_H�8�_!�::��H�1��M�A"�?r��z!�!�Q\#-q�SN;$2�0Mێ��C�����l2���!1��E9+�#yYOB�@�aE�!����B���P���7e�F��>�ߛ��5W�� k�1�p��� �۝��-�.�nm�V�]N����ڴ4�h�֢�w���o7�l,��n�fx�ko��wO+��ާgi���w[��m��=z�l��0      PN T
��  �  �Twx@�*T �   ^�*�@�  � �   *�� 6��[nbwm�}����Hu�]Q�X��[�;v��{r 6ø�� ��S��{yڒ�_7������f��r��a��3Z��t�G_q�7�é�8�#f�k��b6�-��I����l�v!�*����3�3"�l��ƹM8��gH�5/��R6�I(�nGzz[F�y��ҩ�^�X8��>CK��5D!
���hC򥛚H`�I&�n^�D8���i�#5q�!�h�D0��bӘN��>ߦ�iҳ_�iz��$�Hڑ��t8�"�e.����EN!�/o%g�"fEF���r���=��]B�j�m�x�����-��@U6+j�@
�*T��*]7���c��	1�#��dt޸at��gnC�8��bW�V0��2a9�j!�V��M�ܒI$m����B"Zܥ��z��C7ԫ�KX_��7�#�i�>׎��u�������.�E#q�#ya}ԙ���0�V�T6/�q4Ї܆�b����Sn	��$���M��"�k���C!�#���X��4�97!�@��dQ٥w0a��	JE���o ���v�C�%��I�B��=F�Q�"�kI���8�f�I$��g����k�G��{9�UR��SLU�p U9��N�A����J��|�{��Bc�UQ�t�18{����*��<��TR7�II������)VzY�'�ɖ(�v�9�Q>�t�n8��H�IIa9켳��i��3C��#+�Ѵ�P�iÂ���a�B�V�R'm��]TDq�P���yC�b�*t��C�8��]84�8p�oZ����<F�����.)$�4�l+�"�<���܇��eoR�E���%���M�X��o?�???@uv�c�M^�s��aw������`��@�V�U-���4�RH�	������Z9��>:|Tߘ�AjB��ڭ4p��Ѵ�P�i�+6�d���6�m�$`�"�"����-a
5��qT�|�q�7�\:7���go|[�JF�Q�⡼��<D��"�?r��C�C�M���3\�,��0�����$O�q�$��GAD0�>{�{���߱{ž�ty�]��^=��B��Э4p��ԑ��ۍ$�1d�0�|X�=��-^8�����4�0�+���6F�s�I w�c�|�ooomv�l��޴n�@+(m���@�
��ֳ6ow��l�m� Q�E>=[֨o �:���U�Vz!�!Ҝ�p��+���&Ki��m�[N�l��+�㠢E�v��\Y���Z9�CH����!����'��+�ȔI��2G�4p��ݤ�P�4��C}j��h+C�9h�p�]�p,C��:�
0��"16c�1\l���Ѹ4�8p�sVQsx��f���^z!�!���|J-ƒ�F�8n�����K$3>!�b�+C�����d4F�h]p*E�6{I�$O?6ܒI     � �[Y.x�m]j%u *���*�WO���]������ZwN[U��<��f�6纖�W��:����z��9        ` *�  ;����܍�P �R� �  +(P�l  U   �P 
�z��T���<�A�[��uM��'��.�u C��Pw
�pU
����^�2������7�]lx�[��V�:Eyn�u�Q����d^��x��!�!�)R�qH�R(܎54!�Q^�|�C�8�K����ǌ�5`q�(�8E���� -��m��n1rW�"+$4n���0�d�a��<�p:
!�Y���U���@�\�hT�F�RI h� T0�8l���C��St�TuQ�+�v��B��Z�X��"Z
׷|�+�E�$I6ܒ�RDG0��ڇ�8�+�*P�t�B	t��(��սj����DW\�I$L�ҩƦ�W[l��Qӻ����UN �J�'u�ou�ʻ��U㇈�U�y臈�J��f�{�w��;��n��g0�H�2I	��8������]��߳R��Y��ْ�"�Z��L�(���m�m��A��H���<;z"8���,�k�HqT�Q�q �Ua�����-|�7r@�Ik$���ӭ|T�����N��C�C�M���3��]g������L�R-��m��M�g÷�W#y���ap�Y�1��դ)�]��G�*�kzI$�:�yh�N��+m�t�v�r�
��U�ƪwPUT�[�۾>kOP#l�^�Dq��C�j��h+C÷�h�Q��p,\F�(d:C�[�"n�m�$���j&kH��ǫz��/Sx��n���^z/�ʫ�f �wo#��1�$�DJb�<|F�u��(��>�j��@iz�X�M U�u�"�+��3PZ���l;)4䍷l� qV�8Eyn�u��ӧ�XȽAj�b�B�mC�b�(��L�ѤI�$�C$q
�Do ��q��1�XAE�*a�x���d�r�l�uzH$�Iq��!��w^��ݗp����{ d<U�� � *�����{��Cʪ�f���{� �L���c$۬K��|��#9�.�"�<��2?�I�l���9����i��W��'[�������{��;��~>��t}u}}q�z&�E����n0��
��+T����Hq��x�x�f� �C�/ǎv�_&vb&6�RI$�RWw��x�t��Q�Fb��%���M�X����箲"4�%юE$���n0�)ƨap�Y�f��S4;[2^��f��
�Z���gI �[iT�mm��g=�������@�w ^��@w�Ts]Yyg��JH�c���z׎r����>�|�u�#�G��:oR�=�{(�k�$NIM���H�vb����=4䔝��f8\�w�P2�/�PC��d���mFr>Oxu��yx�ӻ�n�cfK܊f���e4
E%�ܒBP��Q��햦Hz,P����(Lr������N�7J6ܒ6�	���w�R�eR�]�d�'��Y�fH\����;wb��� �8@ @��u�V�ٹum\��ݯU�-׻�UkQ(U^�P�T6����۳�5�Yޖ�e��Ҳr��m��Ի�{z���zs��        ` 
��  �  ��(UQ�   �q�  �T *�ʠ P 
�J��U*�\�ٵ/�n[�P	��s*����u�m���or� 6��+m� U�*�����ܷ�n�RI#l&�o�~�돗p8T^��=�f��z5�ْ�i.�n6�Q���^�aw��7
�!�C}�}ҥ�KjH�rI��;jo��u.�w����v�2�Rl���uo��@�UU�UUR�R��Are�wo��u�� ]��"�ⲻ~b�#HS
:�i4��Hc�Zh��i��:}CwVq�i�1�DC�B�C��0���Ͽ����G���=�Չ�ӽ�� ��PxU x U)�p��HF$��َ8�q�;�C�ax��!�D�U���r�y�8��Z�}�$�R7$���qHY�J$<�P����+��i�sn�#��Uԡ�X8l�w�j�1���D�m���w��<B{�ڭ4t��ݤ�C,��=8��CH��Z"0�%b��0ۉ��F�j(��DaWf�B�� ��(q��1�X$B�*�8EZ���8[�D�m�#NJ����R�E��%�D�6�`�a}��qdw!�R�RI"e��ݗ��[�E����w ��*�� �m
���V���u��tqX�,鲷Hc5#HO4;U�����'z��Nm�Y�"�>��4C��$�$�t�tg�h��u[�B��(�t5C�H��8�x�f�!�$:��̹%�)�G�O�w^B4�p�%U��fm�0ID�:a�J�Fg�5��I"I��(�uő܁�Q��Q��~c5}�iL�s��Y�㫙�aVVc��)����m�a�ZEZG�oDG<x��j��a^�R�C�H��E"��?��Ns��͚�۷s���]ݼ�mn�������
��
�ww�D�?����m��Q�C�#�9���,"��r�u����M"��F�$aӧH���m[���mFr:���֫M����Q�"����#^k�+M"��z�G�1��ۍ�|�g��V2/P�D3��B趡�0�W���Zl��&�EUH�m��mDᡤQƼy�Z�܇��h�8E�~Ÿ��#N�=ޕ\��Q|������1�ے �4���6��@a|3��i��Y]�,��B���z�
�nͲ�N�s������n�_>�< 
�ª��U ;�`+)��.yhU&�I���6t���:��ѻj�D������:t�����;���Hc�M7#�H�n1ZU������x�᝽j�j-e��d]���% �û9�	%��a��E�"5�������d�aA�47۪���eu����u4��AĚ�F̓��}˂�a��+�w�φ�>��j��k���>kN���i�)�d�HۉHQCC�w�Ϙ���K���woR�լ��V'|�m��I$� *�8U <k��Ê��l���b�����v�' m��c�KΣ���\�㱳���p�r�l��떽�����={�6ovn�;{y���     T 
�� � �  � P�N � �)� l   �   m� 
� *�  �x �=�%D�{t�`5����Sf�{ýe��� ��
�� �* 6����=\ʆH�e4�����Y&���7���ܷtg8�m9$�D�m�)Ζ�D�|�1X��<ēPI�Ni)�ݶ�RF��FTɞ;ʗy���1�������f�#A�$��n$R7S7���g1k٣g�����@�7�7�F�nGc�Gh=UC��F�͋�サd8~��ʿ��<X���@.�i]�����c��� a�*�{��5S�*��*���wy�OnDdmƈN*��,vwS#�?�[��so|���:�|������s綏��vґ�ڍ7(q�Y�����[�_QaY����f2E�>?v��l�܍�$�6�r
�Y��֫�t��0x�>8S.@�pV�g�k��A�zF�m�"��da��;�W��d�wS#�?�K�
���V���]Ϳ��bF�m�١�Y����@�q���[ok!�-O2��I$�D�h:�^M���7��m�ۙ@T;��]@� ������l��UT�?������Ytnm����UP�|h�;� a�7�IrRI$��U���dr��#���� l�/,�4x�_*]@x�{�/���ܑ�h���� �(x�o��l���i�0���.��"��Gw1#0��jF䑲�u�"���Hç�61��,���U��(��ҕg�ν�@�$�rAm������x���ڭ4~��y�"�OP�_2!�{;���Ο�-�m�"}wUG�ۻ{�n/YK� a�]�@��P�j��헻Ң�G	J)B��Wv�B�����||fI�!�"�5���s�TP*�ܒD�m�N:�,�4Vo5>�x��d�8~ɱ�4�g�z�;ϗ1��NI$q�����g��ܲ4�!t��V��s�a�է���C~�ht����$�RITJ�F oj��(��>�(`G�!��웂�+�&�aw ���S�Vg���i]+�V��������(���{�'��;���� u��>���î�y�3��k�w�؀��UUU*w+(*�m�b�gL9$�$�nI Q�`i���{��E� �(��8�!Ij�?CeG*��#��~<�n�m��j4��"c���J��yyU
#��5�sHb��d{6&[)}h��%��m���0�C�.�/V��^Q��}�sM�#�0�6ے$ӑ��Wv�G��w���o31wpv�o�sm�Kur�m�����&�hS��!� Nk*`��	·9��l��՝-"i[آf=�O �\�   '   �   0     Zm�<<��` �   �  x��	��   ��� �� Up�� �y]�˺�z�V��U�[*�k�����:���r����rݷi����ޖ�W���Uݷm�u <U�� �*��W��#ӋI��{{���vٶ3ּ0 ��	ʣn��TU�;{K��<
<��]�)��ˈ=��ʹ6�{m��-�=�J���k��3;���+.9.�ضB��[�	�cw�wm��Q�ww��ڪ���Jg/^����Y9�iZ�:�+�Sq����m��U�<\�Z�Wu�=�X/l��Vq�ww7F^�ح��^�٫S�ү6ڶ�=�q��ݽSzv.鶺�v��ۻ�\�(���m��[�yk�2ܲ\��Y��lf�ys�^[zwz��˺u�`                             �        �P��
�l       *�P       T N�                 *�U l�PU T0�C��J����u.��   ՠ    w � �T @ 1���� ��  T   *�                v칀 � l  T  �@   �            p    
�            6�  �P��@     �� _*�  � +t���u� ^�T�
��  ��{q� .�m�X�������' c   < �
	�\��&���{ �M�s[m�zz�����Us�����:�����뻊���j��r�-J�݀��e�Ѳ��l       ��   ܀ � x Ë`� `*�� 6� <   � ` � 0� PwT�o6�J��μ�����;�M��^m�����z�w2 �C�������UQf+wz�l�qfU�w���ޣ�t�gH�,��_��U��u�Yh��s��0���IhImI$�ED�8F��ܫ�#O�sV#����qp�ܻ�0�#�rʑ6�Q��Wb�g��2L��,�<f	7F�}L�6E���P�0�+s[C��4�JI$���#9�1�4�����iE��K�>6_�o�x�#�AQ�y�䐖�m��"g�s$x�I�r��G��9��N�X8�=��{~~~�*�]��CR�Zv���5[��y���[{T �U�PR��&cf"I�n(�"��x���Ю#���ʾ"���`�q4G�{2��>"��l&ߘ-�$I6ܐ��(�"��s�(-w�f�ǈ�����[���s2�gSI�HLm�$m��R=�#��p�#�Q#�x��(X�q|;z�
#��
�D&ܒ$�n0�Uk��.AF��q
H+VqE��0�F=Cja��KocN7�6�R���Ȣ;�[�FE{9����y�������n�c��8�~�p{�v��NV����b a�*��UՕ� UJ���xw�I-�ڍ��aE���iF+���G�G�#��r��G�Ɣ)�QD�rE#l&�G	#��F���.)��y!Ij�#��ęy�B0�Լ�_�7���)�1x��e�H�'E�`ć�{���a��=X2�+����\�\�F�T<A�,��_��U��uz���ew}/J�v�`Wƕ��"F����ےH�R1@�E�޵B��;ޤpqx�Q�C�<��RAZ���,�?  �l��|��2������ �����E^�PVRح�u���d�d�ڎ��Qp�]L"b7/i��H�$kj`ć�{�J0��ӔF!���l����Q�:oR��B�y���E^��W�x�6V����$Oq�ےFی:��M��6u�b$8�>�X0�80,F� �0��a	�D���M&��Ip��æ�>�2Т0�꺘D �d�^�#�Dvu��E����M�$i&��8�
#�E�J��i�6nҡ�1!d,��G����m^��0�ߝ���HNnwj��*�^y�n�Z��6Ϯ�
�*��*i��VǮ�-����!R;�D"��?/�x�#��bHa|#��a"p.`X8�<DRm�_+��$JF�e�С�bC�>��a�Q��sm
#N����BB���20�Fu$�s(�n)nF�2��aW��1B��iE���lͥCą�^i~#�Q��l���I$I6�a���t�6�DrPE�q�(X<�g÷�P�0��C�Ή����I" ���Y�j� ���wj��"̓*�P�8�|EmH¡+��       �k�p�r��۳ue^�݇��vёƫc;���תm��G��-ݍ�/m�ru���Ӯ��Uk�����m�{�6����GW{�       Cl   � �T KdATw   *��  wP P*���*�� UP*�����l����_ 	ʧ;{v�oV׹�w.�hf�`�ª�UATm��+���6�q�$�D�m���L�6E����!�Q]�*��Ҙ�p����x�HYA�Y26Kr6�f���Q\^L�C�qҜڸE�Aҡl�#ӹ�!�_�k@�!�HLm�#����.XS�����]�&���#��ՙU�rTCM�rF�.jf���Upܒb���½�T�GWS�c���n�m��D܈�ۉ6⡄B��\#�QVr��P�l��9�21.ψ��=oI �I$�HÏ����Zܱ���� *�q][�+d���`�-~���n6�Q��i"χoj��q�s��i�IT,x�Hq;��XFi�m2J��P6�q��ux��U��+'r��l�#�mu�(�g>b��vj	Np��q(ڈ��"��z�#B�/�x�*�V������8�A�����1#���r�B0�,�y��"χoZ��x����`�4�J�c�䇈�%Ȋ�9$�H�h�U�a�u9��ǌ���(�KI�זag�i&�����w���~? ���-r���w����� �� ��VP�*
�ދm����iI$�)qТ7X��0�>#fm*�kC�-��G��N�^׵��l�HA4��m��U�f �Aҡ���(+
!�i��j�p�cG���r�WOLkd�%H�V�Q��lP�!�!���V�O-�/P������:AR�w=���dQͶ/�1��$�l$�4#C4_�_!B��An���(�����{PZ��{E��T�R��4Ñ%���)��4�x��+�e��Aҡ���((9��Y���T(�j����$�I ���޷m3{i:��{� ��U�
�l
�PV�ݦک\�n#C�X�]�Ѓ:�|��x;W��do';j�!�C�Ɍ����#�>&6�RF�]J�G<l��g�{�]!�YY˧#9�Y��<vf�3P֬��V��F'$�&ۍ��q��n���!�C
�TV��Ar�����M+9���:׊黋��rZ��B�*�do t�F�g�{ͱr
!V�j���'&��C�r���6�-��m)+H��e�Y�6<DC��]4Ì� �ҳ���#ya}��E:fN�$�I$��k��s���n��;�wn��>d U��_k{}�`<ATZ��ͽ�ڙR��S~�����~�a�����.���p�r#�����⯎��Ҵ�M+٧$a�22�#�Ii�iv��・-W#yx�{Q���Ε�Q:-2ЄV9Z�3�H�*�#��i��d�ڍ׹#��ɐ��ϭ�2��L:B�T9Z�+4y�6FrýT��BT2$�m٫�����5`qx�C�������U�=zJ~�ST�p���5��S��m�$m�#�?3����aL/���	=��9��а3�8WIDX活��w�;���^��  <o`	� 
��ת[�#==�R����sm�������{�1�ݸ�w�ws���w��8f6��Q�tWk����b�=�ۻ����1�       ��   @ �  lv֠UQ���0 6� Ul�_~� �  @ U �@U���J��[��� ���m��^��/Ku۶� ���Ww�Y@wll���*������N�����D��߭�z������%�>�`��~�
s5ӚN5���6B�T�����r3q�3Vә���t�޵C5x��Sk�,��^��d�<~�1�u@�Q��RI$i�ح"����m>?3�H�2��5ds�˶�����y�T�HM� ��؍?�in���f��yU�6G�rV5�fߦV<�XH�a��R(ٍ�yM�3C��7˟3ݻ�z�m��}y�S��8d�I$����ujmfg]���d m�p��UPU`UVe����w��uڨ]�~~{$�T%�NQ�}%�NU7�N���SC�4�eH�I$0�=�6�o2:fT�k��K��#ڬٲ[nK�j���$JI$m��|�r�����<y[zs������I�����Ruah�h��I�i��j��_��Y��ɮ�rK�;�Ar���x�EB)Y5WwM�"Ⱥ���t'm�����Wܷ�������J���h�}#m�$��;'����]N�n��{no��U����ẑ���k���ʡR�ν�ܼk|ͿL��Lx����\�	�yM��V���mbG%�[���[֤�z<űl'��� �pu�.J��!Smģj4�i��vR�νZz¡�_�M�+<�l�O���Qz���x;U���^]���H�!l7$�I �׹#���ui֗���S"0�
=P�9h24�l�Y�q�
�F�m��j##48�:|r��P�^5�*i�0�7T�K�d�<D:S�HM"Rӱv½�p�$�A�4b@���6���� �� �R�T;�*T7Z���� �_����w�~�1�)_h2<xIڲ#��L�G"Λ(n�b�g�Emu�*�(�h�����^\/���8�>3MӘ��Lחo�(�tä(�C���3�úW������wq��8Vk�;�lB0��c��8�UJEL5�F�~=��^?q�[;���9 ���-�C!i���B!�!��
��A���NՐ�/��а24��_ ���l��jF�8С���CU��
g#<�٦ߐ�C�Ɍ��ϭq3}���g������I$�I�����;�u���1)r�v ;��UW��*�� UWw�W|ƃmUWj��}X�#J�+�!��.5&*���=�j���z!�s����.�K\�Z�-��fH�i �r#��]�	�U-;���0�ɔ�+�28蓵d:C��z�nFc�9$I6�a�F��gN�"�X��BX�j���Y�i^�#��n���kK�tH�-�.H�JHڦ�U"8��D.�\kMD4�*�j!��G��Rb��,��sV�ƢF��MZ1�$���qHZ5�Αv�j�g�"�R��p���5ʄCg�����_!�x�	u���G�A�� '  �w�m��t�nyU1�ss������lQ�������+��Q�g[���Q�ګS<��v�n\g[�wfĮ�oub�u�=oc�      ��m 
� x  p�U�6:r6���� l 
�7�U���Sl  U  P  A�j�k�Wt{�n� mm�K�u����lS��v�l���ql��
��-�wv[�5�U$�����#�/����CH����慇hB+ ���kK#yM�ҽhB!�6߉k���@�Iwp���+�pא�2v"!��i��A��s�J���X_u7GN�ڑ?.#n6�Q��T7���0��^:E�~=��C�C�M�B���j���0����h�����n6�q���#�;�n�!��3ڎF�t�"�c��Q���l�\ÆϞ{W�n]Ee��2�d�<D<q�Y2���.&ߦQ�H]4Ð� �ҹ���Hqqw�n���ܧm��m��;�kם�{\ a�^�e��mT֫w����IG#t8�:|f�s���|����#uu��D8T�T-���ѿr~6Rm�M��uDi�O���aLh��i�~۬f��S{FF�p�1r���M��K�K�I$��Ê���+˅�dql�ڧդ\ZY�^�S#M�6B޵Ƹ�4�37��@����*H����X_u88�t��޵C5x����/�Nv����F�+�l.a&�iI$��B������:F
�jada}�뎴�3W��{�(it�Yw��H�H�q(��ն�v;���up�Z 6øUomTF� *UU݊��oPUm���:eDx��
Ռ�dg�4ޑgL`�Ld^�h�4�eΖt��HJ,eܗr7i!g4�a\�Mk�p�Յ��8�GN���T3������U���կ�%�$I6�h����P��h��ٻ�lke�n��׆j�TF�\N6�RI$��4�:��͈3�ad,r�g#<�ͥo�B!���ɜD���f�$}i�$�$�iS�S"0���r��۪���Y�9q����:r��P�^=��{�l�
��T�s;�v���n�޻[� �;��]ʩ�eQl��wm��Wu�f���i��p��<Gi�.bq4�*�ad�W�Z�w�
��b9$IFۉ�U���^+A�Z8Yң�E���ՎV���dg���7�5�i�ŧd�Ikr7n�!i��-�e�t��r�W?T���.5&*�A8Yf㚨�ABE%�[���T3���0��^Y���z��~�J����L˕A�Ҵ�5�_�i���$��˔��{�~�::����x^�޺=��c��� �+/P�w;B��"yf�y�$�I���]����nk�c�[�� *�p�ʥW�@ASλ�j����=URI�_j#��t���	��d3�a���rʠ�ҫ�D0Y׌qd;fF�m��2C���dޥC�W��0��^�U'goEn!�4�S���U-;uo CM�ܒI"��dxM��O�8;��
#5YX��CH��=�A��ش�]��6�M���R�8�H�'�W[R�#N�n���yw�?������u{�w�_\u��������M&��Ip��Q����`�(����f���l�#�N������;�￟���V�< c ���[jYmlk˵A�Օj�
��U]������ۣu�d��4��6J��wd�^��n�5����1|��l�       Um�   �� � � \�v� *�����   
�U*�����  
�*�U*TJ�UTp�� nyW�Ǡcm�׶��u�m��6�j��m�UwP�� 
����w�m��UvW���}���~_��aFM���i��vZ�D?kv�����:Ax���1$I5 nH�1�C9C�!�pv�H�'�m�������5��M!���	��_i�(�f�	�_ܒ�m��0�HiUf�B�#5x���E#�6���_k��J:E��iq��G#p��"��z/�Ҧʡp��˵ʄCfGd�
��A���NՐ�/3ƴ�U�IM)8"Λ+��o*/��oj���+�;��ܼ~�m�}\E�^��':I!�9 )��)��k�mtSw�m�̹ C���Z.j���*[k�iƃbmĤ��4��N��Q��[\�R��<�wU?ae��5`qx�X~{,�k��JI"I����GH�O9{�{���l��4&�)iz�m>#�<x�����#ǯQC�H$�4������F��Zz¡�Y�eo.bÊ�D!�C���)�z�=���o�~��.@�Ir�$�8�:�6�2��L:B���H��Nv����X_u ��(��;R\��܍��mF���r�|�����H�Oǽ»��S%P�Fbf��*�a&ͻ�;v��jW����{n[��.� *�p+=J�P� 
���˕�۷����H7�7�<s�.:���^)�=�`dm�t��P� }��BESL:D�^�;$!�ډ$�	��qQ��+fT��C�g��l�������"����+�������k��7M���3C����+x����^?>�����U�z!�!Ҝ�!l��˵�9���m�䑵��������G�	;VC�8�S{Q�����N�"�E���zQ��f$ҒI!�3���Sd��z-?C�朩���ϭ�}����C���J�UV �T�{oj�{^�����]����pw
���S� A^��C�wwr���\�!\h��g*A��Qӧ+x���C�)�������N�����M��B��$ҒI#l�خ"���r�ن�2��#Ǥ��h���{֍"Λ<��i|dNH#m��q�C9Q|��x;U���^]}ގ��i�w*d#-3�\M�L�!��Ջ�=HB\J6ԑ�5��E���2!�Ƥ�F�#,�8l8��C�>����.קv@��Ĝ�$�nH����x�t�r��Fbf��*�a]ML=�<s�.:���^:�&�F�vھgu��<M���^�λ@P�ت��sU©YE���6��يm$�I8q�<x���lA���C�X�X�Ǟ�&�l{:�۩.��d)�D�m�$��U>���K�)�g��P��v�ɍ��\�'��f���)5�.�T�z�^�u��49�[�;�wl��.��k@����$�&ے0j�L.i�f`Q�ؤH9jH��Z��}]��Z�U�͕I��nH�%G%��|-�eM�\�W�W?T�1�(�3�Z���vF�s��FM���N�7mt          �   8@  �{mTp��=��  �	���� �0  �k�  ��;v�1�p��G���USdr��f�m���g�ڹ��3r+w��[Y�Q��<�[�n���L����
�
�e�`��S�� �
�*�YE�;��;�N�xN�ٞ��NɌ�+� ��O�o���pu`=�j�|��'����B���7YWM�v��E��v�w���X�' oq��ݻ��l*�]U[�J��Z��-��j�ͺ�[%�@]�k��ͩ�walf]�.��I����j�]�Z���l�δ��n��V2B2�m2�@�K��.+iRZ�t���ٯmҺ�۹��ݵa"�j��9�h�U�׷�w�m�����wJ�m�n�kYk�sl���׷a���[n��(���;��ڤy�ܵ{��=h                                      EPU *��         R� ��    6�U              z       '�
�   ��  �� U*�����0   
�    �   �  
� Ȫ      P�T�         l 
�T \��P -� /}�_~� ��U@ 
��  ;�         P � c         ��    P 
�  -� 6��P    PT�  J��� eO�Wm�>� 6��کT6� ����P�kv�3lwx����ۄ��p�  N   ��UuN�sʮ-��m��pww3���n�2��wm'Y���wl��{���6�Nؼ�ڷ���ok���z��c�=���r       N�   <  ��x �TVJ�PU�+)� �  �  �߿O���� *�@*�
��*� e���ȓ�c\���W��=���V��T;�+Ԫ p�*����M��d��d�ۍ����VE��?�3�F��3����^&i��iZYZiW�_�v�$��"��0�p�v��A/���q���)�T,g+/��y����^]�������(�m���G^�dq�4�>�"���M��"0�	�0�5���g:�d8C�o$	Wd�ۍ��MDqt��o�k�uO�#uW��Y�D:T�lN"�iz��y�
m��m�r�a�&R�2�#Ǆ��!�:/�^�5�Y�ew.B���k�$�H`���I��u��EK��͛�ր��U�(
��l�r�f�j�k�*�3���Pl�Y谈|m�ʘ��Lא�o�`�L:B���24���ZP�[�������4�Y�����,��p���^#�x�8Y��g�����6f��j�%4��l�خ"�3^Q��a&R�2�#Ǆ��!�3���{�it�S5>nEI4���!�4(o*/��x;U���^\/��',"gr�22�5����X!����m�q��RI	m�f�R������1Q�FY�p�qi��FN�h�i�}�I$�H̅��e�f�ܻd�;��ݞ� U�Uk�lU<AR�z���K��ڧNS���E�!ҲJB���j<�!�!��S�x���U���^:�{�rH�m� `��"Λ=�A7��q
�����)�z�=�gr�B2�/�֭c����JH�b��J�<l��L9bdi\�R�C�ԜL�\���N��r�F/��!j��$I+qsNWz�c���_�ӣ��U�\�X���i4���7�k�|opT�"�n&⑶qW#yx��aV�e�*E��QB8+V3���Pl�U�TG}r	$�I�D�m7z7{��u��� *�px�̪ w PYs�Uw|k�2���u�>�;�Y��-�,�HS6̴�ҳ�D3N�|M�5/J��%;#�$�$�Ff�r��x�}�8��.���p���!ҭ�"���j<�!�"ۇj������m��q���i9ݗqd8�S{B�F�t��aņ��,p;U���^U�����j7Q����ʈ���ܩ����y�tä)��k�:N{6��+����k
aF�F�IH�f��t��o7�Ҝ�FN�p�n��~�=��J���e��i~|�~w���;u�婃{kv��8+����{( ;�1�`,�R��-�ܒ6�2X������i<$�Y���L�YҜR���])�%l$`��wwwJ���vC�4C8c;�2�����ذ3�)�^o���쒄�(c.�-6[�1Zh�Յ�RsH��NV�9Yf���3M"�?j���4�]���%�\I�$�H�Q
�*-,�΃L:t����p�>��Zl������,��{Ѵ�&D�6�l�3�|Dpz���,��vC�4C8c;�2�ig	{|�i��Ȯ�}|�nI$p� ݈ 0 
	�+k'���*��9Q�� 1�lQ�m�ڪ�i�U)�k���uK�d+=�5�ȴ��dnQr������ŀ       ��   �  ;�  *�Mhm�lUP �  �  U6��}
� �� 
����n[ٶ
���Iz��eKl�|�+���������@P�V�*�����nWVɶ�ow�׵I��	��p�+z��+M��������`�+,���/�Vg6ʳM��M�$����c��`�4�6��,��>����!��U�'�
p���I$�"pVdC��Ѓ9a�ȎV�<E�I�6C"3�S8��+w��%��NIM��R�#M�3>"��ת�����Da��0{U�l��9�(�%��
3B"�?��dif�&�T�Yݛ��Hɴ��g�Y�7nI$�H"Q��V�W��z�v��>l�
�� �Ue� �:�#�_1BVT������b��>4w�2 �TY�&8+V<E�I�6C"[H���i5R&ʎVQagI{|�ih���Y�T��U���X^�qFf:0��\�-��kW!���!ҽ6��T����di�&�T�Yݛ��H}��͕i��m���V�k�=�Α�iL��id�!c��Α��v�
8D��v�G�b5rI#l&�u�Di����*'���r���ghËл׫'�Բ�$rI L��q��ݭ��Z�]�� ;��o�� � �����KeT�(��y��Yyf|ER~�΂�l� ��D�*��:�W�zG#rI$�9CH��2m5<Y�|7}u���VSл�VdC��Ѓ9QgH����E��Q�ԍ�(Q�%���Gw�di@����L0�._*F�!l:f|E����`e��R	$�i�3V��!lL��Yf���0C�*��,�+��ҋ���6�	�؍��n4+��XY�ap�L���~�y�Ҵ�3U������~}�]������ 6�������:ܖ���z[��m��]EQ�[ �sfZ�"���E$ԍ�".4(g*,��y�!�֍�����#���:K��|t�:�d+&'$�)m��5���ܮ|�M�����̍�c���e�����KӖ"������7m9x���P�EEe������jYg�63/kM����W��ʉ�"I�䐨�W�C;ڵ=�~ٚ�
��kw{�׏�Q�.9�#VYS�4��n%$m�EԪ~dvæag�s�o]
#ؼ_iO�~�}��e�����=��ٷ��7{���;��{�R����UP�U@�
����W{��d���rIf��'�������Y�ER��dc�"߱�e����I������6�rP${���+�6F�����<GV����!��ގ�~�3Z��y��I	��eGXDkŞ%����#r3ş�޵�j͑����̏�~��8ۍ��&��e��m!�*��Y�W��AY���U+,�F0�8G`�-I��a�ۍ��U���}�}+J#5Y[
�A_Q�n� ��,��TB>"Z��~)F�2I$�I � *�0  8�m����v;Uz��8�NWwm�h8�m�cw�]�z����T/f+нSŶ�2�So:;w�Mu��go=��9+mͻFvm�        � T <  �� URq
��;��  
l  ��UUPT ���   V���-��p��U���R�%�],BYP�!We27u� ��
�� �� �Sm�x�UZ4܎���~�d�XD����`�0�C�x������V�#ua�&W�(T��P���D6;8��VY��(��T��΂�~�
ըL"�����i!l�ۍ��FP�4�6��Y���^�ҍ��➅�}D3ٚ�ڨ�����b�#%ݤc\�}r��9���v�WQx����0�=H=��adGy��c-�v��n_��p^�g�o)Y�5$u����9�$�)�F��fY�q���d�Wr���R�Ҫ��UEe[�wv���׳���k`�l7k1��w�4_����d+n
��g=�W�A�䐖�AF��E��pQA��Ksw�����#��5e�����a�<�Y� ���F�M�kK?Cݶ�֟�W��)�ȳC{����
#���s��o�����_ŪJ�����4��Y��s&A�a��#R�6v/7j�O٪��Lt�I�4��IeIx�"���TY�g����.��G^4F��j>��^,���$�I$���z�+�7-���뛞��ws�U ;��:�U]�[A��q�
UP�4�u�0c�/5�;���+2zٛ��TX${5%$��"IFxC�s��dib�'ѫ,�L����F���g7kl��I$I6�h�/8�A��K+=cE�$���a�s�u~c��+�(4��gn�u�Di4�͐�6�m�d��}�g�}�CH���t�,�T�z�O٫NI���4��tZI$	��K�W����`��{�6
�^#�/W}>�x�]հi~ߞ��$�2�L��d��q/]n��'c��r 6ø�e�;�Tm�.�T?�nHۍ��*H�ş��޹Z~�VVº�"�
+{��9QgH��A��K{� 6	,�m��M�x�Gm(����#���F����^(���k�?f��[�|W��n6�QC�!g�v��<����!�E��ѡDi7Z���6��2}��$�(��4�6o\uچ��Eu�i�7Vy=��%iGR[�Ѓ5]��L��'�B�q(�h�СGH�����ҏa�}ZEE���u#M�3؆e���� e��U^�����K�ẁ
��*�րGp�
���g��ۡ��I�$�B�q֛#u^)�_��bnr����x���"�?���B4�ǽ%r8[m��dWT�PR��C,�nm�F�#�7q�!��Nh]���"u$7�(�iD�rD]�8:-�<D��B�,��䞱X,�D�Q�i�J��4�4G>더A�9$%��e#f��Y[9ڭ6F�S��!�����Cz�쭲�O=Ib�*9�H�i��2f��dl��Vn��ި�ssEu���,���ɂ�I$� 8J�P   ]H]�gw��ޝf�9���Z��-��<�����μps*wy�o(�ӫ�kmsmݭ�m⩫j�v]K���b�-vަ��      �p     
��  x�؅PU�+u� m�    �ت G���
�P  � 嵳e�ZW����n�weۼ��v���X� Q�T^���� 
��[m����2M�P�&����~hX�Wk���^pq�%���@�Ə�Gi���ٺ[�zW!nB�n%$m�-ʯ��4B�ƳT!��<�����
�CGE����W��obM��I"I��m6hC�U'�������rk"i�b��ҟit���v�t���JHR�T�Ĥ��r���<��]�V���{w�g+����Rq�%���@�Ə�FkT�K�mF��ۍ�Tr���uCĻ����4BޥƳT:~�����df�j��>?;�L�$�H,��rt�ڪc�ur��� 6ø������ �ʛ6��-��/�����>?c�AQ;�Y�׍���+T�*,�ͥ>p���L�CH��$��܎�P�H]u+�3V�}E{ �?s��{Uڇ�|�A�H��9sD7��F�i��?�9�iF��P�5�&:����h���C�{��$O�<D-��%
��(��tt=�|~��>"�w��x��k�dM"�x�3'A6Km��j&���#۽q�p���R��=��B��g�n�c��_�������1�meO�y�����]�f�v C���� U<AR��m�(��	��R	$�4��]��ξ�V�}Dp��>l��(q�<@����D��rDbl#���Ņ���0�yܨ{��>?gK��N{�.�l��)q<I��I$�(Ȯ"�n�^�)�Ä{w�:�P��} ���F�#س���i�3��p&@�m���=�ݪŇ��V೤K[�ށ�����O�H�n�k����a|�ށm�"��\QCY� ���#د�	��i��9P�*���}�!�*-�������ol�v�:��ڦ��7{� �qT�� ��{W3rH�m� i�ٯ?y���U,�ͥ>p�n��]� muԬ(�b�'{ltF�I��H�jF+O���\ �����R���-owz^4~�s��*-�uy�Q7	NHLm�#��U|0�o.5���ާn���x��O��M��ʇ�W�>?*�26�eG
:��[��>ךȚER�P��S�<c۽��r�H̒Wi$����mƁNV#س���^����Ac�n+<~{+�/S�z�g�w�/�ߟ����{i���շ�{�w|�[ ڻ�
���� �m��7 Af8#��#q����T^�
�U�gÍ��EsVY ��� :G�o+����^���M�#m��n6�n*�^P����8ED��K� k�dl��fū3{R�/�T���E�$}绵�W���PZ��ҧ5��gs�dY�2�'�ɕ
���m���nφǺ�i[�+��t�̭�F�g�q����m��*����z:��C��>���;��h׍��=Z��Qf(y�����   
� � +(c�gZ��;�n����C���f�n�
�z����[��aua�x-֕�֜6ƫ���.��t��6�v�n���:�˗w�{Y�x��      �`P �  w *���7� �*�  �  u�@�  @�A�  ATڠ*�  m��@1�����+yz���]��@P�V� U¨*��\�(FBl��I��x}Dg����j�O��uܠH�/Z}EwAZGݺ�Az�ʇ�����7m��m�Zj��,��G^4~�k�Dkŝ%�ݡ�#�x�,� ��eZ���iI$��T!���Jz~'�۪���d]S�"4�V��>>���Ӓ�m7#5�U/\�c�����?G��7�
�T�+�u��J8�J)�/U@��I���n�G^#�������Ud"=}� �I$�(�0$�,�ru����F�� UA��T�UK2�l5.8�D�J�������P�_��ѩ���}��^�>�D[�dY^XD��I�H܎4�F�GسY�h�^����3�/s�:�P�2ut�H�/Z��ц��I"I��e¤�����+ڄ��O�C�����Gۅ�"5�(Ub���7�6��`.�����s�/���[�U�(@�Η�)RII)r��#Oݯ�5�>Ś��*���{��"�;����_y�� U�򪪻v^�/s���׹� �d�Ī�]m��V�7��n%$���r�~^������+ڇ��o����f��^"����-$m�warIr�\�q�lv�����ˍf�F���v�Q�^St�4��Ab	�Q�m��r:��B<G>�����]x� c�iK1B�j3�����'���a�ۍ�䊻T#J#Eu�
"��i�z
~��L>��(p�o��"�o�$V�&ڍ��i���|s\�#Y�iB�~��r��y�~��L�I$�BR���ov�g�k�ý� m�lUU� *��TVm�5^�֞�§=��	��^��g���ަ��w9jf7rZ��I6ےF�ME�����wvuT��|t��������ԇ[�M)$��Z����o�kƳ7R76�{�q��Z����cNII�\�'�Ky�v��5��ޛ=]�ӕ�8jc��Q�R�Ai4��I���V��|�3w�>���0�]��w�k#ݽ �I$������={Umr�޻sl ������� ASe釫n�¯J����>���pydj܏lV�|nTǖ�\���s���g�MF�qH�m99�4=�k�������s��[�VN粯w�Nȑ��$�r@QnI}|�GE�[�gNx3۽Q��ݮ�0�=j�s���I$�"ʒ�۫����6�3�+{��w��g>ީ���m4C��$I6ܓ�C/3;H�r���c��Ks=\zSz1�k�N�t����c���r�Hx�����l����yYJ
{�pΆ�">L�*:	�
6dR�9!M�e$(�[pҪ��R��%"�o󰂵�ROf�ٷN�[����*�eE	q��z:^��>��?ˏ�������=�������~���(y���~_/W �!��c*��������uiy�N���Ծ-�{���"��������\���]{�s��=��������()���!F*�e$(ĤN�(J�K\:'s��"�z�}��o7��Ǳ�t���s��"��N��߆�_??ٷǗ9��wk������ݭ�6�"���������ß��(w�C�������J�����g� �(q��������������N;6���ڨ���yt��ꈡ���3������gol��X�O/Ouk�*����|V�Σ��TE6��'_w��S���3���F����yq�z����ߙ�����9��"�&;qϞ:�,s���:��::\���H�!��wG�׿C�J�������y�w����
�2����+� s������y�>������     �� �    ��X ��\r(QE�㪢�s
��w9��УC�`tQE�-3����Nv�۩�(�gw*�[��P��ÉWu��T��T�7*�\ ��n�R��r�W-J�Ҩw\r�� 8��R���:TE��JR�v�T�s��xh    �&��` &	� UO�4H�%SCML�C@2S����Thh44bd��b�Ǫ*P`LLa12Oت��@ 4     �H�4�&�Ɗy2j�������$�ORy'�~��{�@	#?�퐁$'��H@����	'�'�?��p�I�F�O�I��'E@� I���HJ�@ I5��}�w�p��z� $���
��?�?�4��~�����/�т��A�4P��(
�E�""1c"�
(+"[#ib,b,���`�1����*���XVQ	B���T��DV`��dX�����@Qb
�*���UT
��%#h[b�-Kd�"
���
��R,XAa�(�,"Ȭ���
�%Qk
0 im�,�Z��KYH1����b��U)P�+!DRکR��1AQ ��`Ȫֈ�#"��EV�QdQX�U�X���R����E"�FAdXXh�)!`�m%�1�E�(
�
(5+Q��1b�AQ*�V%�Q`Q�b*�E�`��Ȣ�����mZ����
)EdV*,����J����(,�aY"�X����X) ,�AV� �Ud ��*���)���V��I�$P*�*�P�@$"��V
P!X�T�`�$�P T���-��R��T�eH�-�mAeI��
�Qe��`�Z�jV@�[J���)XV,*T�[,�Ҡ(��ȥ@D�m��IP�Z��mJ�mRU�*HVЕ
���$U��	Z$P��,��R���)�%dQH"�� ŭ@PAQDdPY""�R���� *��T�)F�"�
�dE�����O��&Ji�C���w�{�q�{�w�����{}�j����vUAl�T*���m�U  �;�wUP� �4��:��� @"Y	� ��
��>
�YA�j�AYyV뒂�cj���6�v-��QR� P�   �  � U�wn�d.���b��ʠ��j�S�|��|�5�;�Y,�7WR��T QT[+(V�U�,�uQl�`
�T    
� \�@ z��#]����2�b���m��۠lP�le
��uT��l�U ���UP��]ٷ{�@*��R� UM�Z겁T�    *�P�� 
�d    ���   R�P �  �P[%P ��>|��PU Ee   UPU �U  U   P     TP    *�@ @   R��*��l�
�        QT ����̠ �R���07J���   �Um��Fd����AU���+)R�f��ATAY*� 6y��*�Z���.eP T� *�� m� +( Y���  ��V� U ��cb� ��S�Ul�Y�Uz��UU
��o%�m�`[  
�|>l� 
���U      Z�] U
��k�꽀 �k=�VV���V�H���c	S��vX��9�
�m/ ��Vs5�N��0-��0�*�xcB:���F�HB�[7-U��]��۸�L
�ݢ��Z��H&�6��wT��̫+˚���p9`�	�-/,�k��b��`@%K�$�����뜩A�����ݞ4sһP\c�{A�p�b��[��.4mB��r�{��_�m9{nr=cMUUP �U*�s <ٶ� �
�ޭ�m�� ���  ʭ�P�=n�d  ��@   �݀ |�|���-� ���]�ݏ�����Jz�r�p�'Om�L��nf`y;��O_�B$���HBI���z/����E"+��ü{�����v�;����|�HJ��i�Tꢻ�0
���P ��Pr�o`�l�zT�ezٳ�U�l�鶁m� P VUP P�� @U      U 
��lTcd�U�ʬ�B�@c` �ۻl��QT  اr���A��wQ�#�I�i�r�B��-�a� X���y�u�Bu�Wu�;����P���Tb� -�������z-)i�@c �X	P�  �@ez��u�c��u8��>w��S�\�ʹ7+���f>�6Nm���g�}=unC��Փ���m��s6�|so�ww{��;νcٽ��
��Xy�c����L̳�}Ɍ��6���we�����J6`\3s��Ϭ���7�C�P�m�kt�'=٨��k�b�Ny|�]Y�g��v��g�����8���f2��/{��y|���u�ϙ����fی�5{�O �	krfkk�r)Ǵ�jNe'~��
t�gV�q��J�ɜ�.]1wCS��X�� W=+��ub��v��R�73.��jc6�c�0Y�Y�h,-��(`an7$�K����19I�����36��Ԝ�c����_XO:�jk�u'~/:vt��3���15�_9�HH�>�~��fe䓺��UP���Yn���e�ua���f8N3��'��&�C���K�'I��)3�+<��"9H)�'I�=S�3a�c1�2L�����`*��@��< YEe�ԪU@-��zʲ@��9���
R�T�x��޷t��Rg�6,�2�S�=s�̸�a��1Ԙ�z�<9���P�Ԛ��w����w�je �^���W*8���hH]}��nf�Ѱ�]`����9d�]a�s�59�C9��_��r�}���a53�}�۽wgӉ���a���}g2�eJ��y�bc˘�֮}���AUm���-�ְ6�v� W�u���Lx����q�*nY;MLf�z�y�w:`���/��!�(jyΗr擤�b}m����L��������|H�nX���ۙ��v�^��N0Y�_L����y|���u�'S+��a�:��*q�v��S�Iߍ�*�'հ�\`��d��n]1����Rrc0��f{wV�����#�.t���S@ݦ�T���˲v��Ͷ�bW=v����]�P�(js��MLg�9��׾���YS��8���ά���Ͷ�7Ǜ�M�!��s� *� U
�6���R� �<���[��ҀJ�����מ�ݼ��<!�(js�O:�M:N W9u��eL`w���^�S�I�51�l1����,�W���p�u��������;N8L̳�g��_��=��p�n\�4���s(�N�*y�N�S��36��1+�%�p�<睭����551����<�쩨ff7)=w�f\N����c�0Y�^�3���̶�@-�d1-5�{���Lf��z33�9ݕ1��L@��z�ٌ�&����!ކ���a�
��T-*AH)� �c*C��~���R
AH)�}��Y5� ��î�1 �'���N�������wa���N��X���zI'�~����ٛ�������-�)���!���C�Y0&�'-��0Ԙ�#�m��kVĒK����O\���	�Y$�z��w�=0'l�
�u�&�	��	XN�I76���`Ld T&�Nz�8���}�s3��u�nj~�{S��UUM��w6ۗ9��g�Rެ	XO|���t�N��'l�
����$��	�	狀�t�8�t�ā��'�$���@�y�� t���d�q	�	��
�w�&�	羯y�,	��T�Nr��d V�����O~g���dbRAP�r �P � �����)�������G�O�j��暪���z������ic	�LH`L`J�v�=���Ǟ�w2�ׇ���̒$�`�a��w|�{qd$�;�   UVF��L����*�uG���y�=�:N&���q��:��Β��9��C�(js�Nq}�'I�
��a��S����Ό��
��O�� ���^�Ox�t
�f��`���<�¡�(jsη���;N& Wͺ�{��>/:\Y:�2{O6��51��y��׎0Y�_l�f�P��W��I�t����^��^����K�]O1mX�����yGH9����33'I�ul1�,įL���\s4�y�Nr����9���xÝ�S������)5<��;sd�'S	�o�F��e�����DU X�m�Lv�<�*�Nr�������6���9a��MLCιnI딚³-&5�{�s)�_9�P�i7i=z�j��y�'=��<���u��q6W��v�AT  Um��AU��L��uN�5�:#UUUK� {9��A���o���y�w��'�Eo�'��}��'hV�q�:������'Ić�I��q�v�N5 ��u�P�ym��33w3iw[*����5
��\a߯/w6{g����;��{��Xk9i1��'���fh��T����`v���g��_������g�xzUUTۖŶ�xOL+��߯+�d�(u�����g��fi=uq��a��MLC�����LB��Lq��of�g'�%�3<��n}�۠ت�۔ɢ��ZP�r�=Xbq��8��I�
̴���31Ԃ�'yEm&���y��'hV�q�]�c�OU²jf�}���3,��]�ڸ��R����񓬢��xy����1
��\`�y�\�bq�����ffCX�H/:�YsE:�ݤٙgٓ�����oC�UUPlh���r��RyR]�*�5 �ۿw�Ϝ�Sm�ݷ���K�  c�*[����ԩ� �*� ��@U@�    *� +( q��[�B���J���1T���UT+/V�dT�UEP�6�6����ug�W[���D��"�m�x1�8��н]�i��en�y�U�
��T�H�2(�5m��P��y���7��mUw������;��  @U�wIZ]�����p;Zx�,)	īU[V�+��w��y�q�����<B�-&5 ��73;�7i7i5
χ~ׯ8N��L7�Md��=��rO\���i1�:�ڂ����8�B���}���a�i7i<���t8�����,15�sm�f���d�fZN��Y�� ���\�3mϺ�v���e�ft��z���@�89�H��1�ScQs��<���Q��^2{����q5�Y�\� U\m��-P�B�{ ��zM w�Ms5#�o �`v����/: �����V[k�%��@�r�8G:c-�.����I�R^�]`�˚����H�B�X�,X�z� J��V��jrN�*&���/��7�K
�h��kh�[��UzվY�77_4S��ZM�I��z���&N� �6��np����kQ.kmkޤ�x�V�#uHL<t�5��g;Y��-��LD�D����c���5�͟m�����C��{�.9m#�M�GE�UŊȲ��=ssǋeg-u^w�M�Ь��2�oR󑡽��$�$�n#O��eZ�g5%f{�.�3�ٿI�Ǟ���W��g1�x�ܶ�'6m����
�*��*��Ul� �������K�� @- 7"�2`�_oV���9����mm�h15�p�[=<'�޺?D�*����- ��ש<wV��j�?w��u-r�Z֊�,��ؓ�-��2l�1nRX�$�;�]�'���Z��;���̾�$%��m����=?T���ڸ�M��pT��rᔰ��D�$��4"��ֽ��e'���q> ~H���	gm��X>�r�*�@�k�[n�7����_)R����W�3�縊���3W�\D�D�.��m��� *���b%�m�In]c�ې�^;�C�{l�� Uܤ`E8����-t�H��e���s�&��u�ۚ��r_5 Uk�.����}Yfu�A�*�'5֪��.z�fB��o�k�=���UU[&J[i��<��B֡�x���QҰ�|dxG��-���ka�u/��UP��fA��8�b����7 ��=��+�����C���)�+:��8�*D���q�߂O 8�.�56��/=�u�,�y��9��w�પ��[F�l��� P ��*������٧[v�r�° ��ľ��o@�/o��� b��D�C`o�Y,���@H��Y��ꚑ�m� =�Uq2�T@���;_z��jxOj�Z������;�~z�&ú��\UUTµ˒�d� T��<,�K�J�M�V1)� ��`Y9��\���$�dݾUW�\Ժ�/��0��F�Y����!�%�*���]]� z\C�<ڪ�db#e���i��w�Ǡ\��8������u9�@�Z��e�{�<��*�l��f�i:�2NҵJ���Um���6U��+-����J��u��� Ȫ+*�� *�P*�ն�
�   *�
�  
�TTK�� �@��[   
��n*��6�E^��Ų�9�6��݅�+ftj��zл<kl n�IU����v��PZ�kǧ�s�^�����s#�T<'�{{7o~ǚ������6�Ԫ;�Ϡ  U ���ª���:e�+��w�mE0UU��.Y).����^|Ĺ*�４u������
�Nz��YXI�t�yUU~m`�8�A�k[��mFnV�;�T� ��-��I��27\hG6��2��	j�
˚���Ǻ�Jhd��3+��|y!�V��ͩ��Z]�S��H6�N>|�:�z�޸�C��K�(	n��Y�$�{�D�wB�
tI�Z_a��W(��`Y9�Y���!$��{0�
�vyna�oelf��.�L�����kh�6���@  
�e*���VN�X	��u�V<�^ ��-UU[ ><�n�z]3��8��j��Ά>���u��j�*����O$����0�Mfsq�EZ�;��;���%b]�N6ҕ�E�7	 �d�ޛU��e�����k�	����
{Yr�'o�9t��禺{�Z�{R&sZ3�ם7lȊ���$�h�.�I�0ȥp;��[Q�S�_��¥4�N��3��� �R Xሌ��������Z��4��lwtL��B�٭e�-�z{sשqU��E�@�
�T�ڣlUUVug8�j1���Gǯ=��J@=����/x*^�X�<�M�� sYr�&��U�BH>���̒�b{�(q$P�r��3����i��7sE:H�^(�Bw��P8���ZQ��)�|�9�`����jɐ�<Ǡ^���4�����u��~�_�����w�\.d����D�'I��O*6��9��P��Y5=��
�Z;�&t�\���9�����ܴU�Tl��w����"�Vr�
�����$�Fi&�a�K ���c��P����!�<�[j���b�   L��llJ��!��+�6q���zJ�I�UYء�A\MH��=��-~0/�s܏-Q�*q[Θy%�ki�z����Q�5�.W�Z��sv�&W�$�oy� �д����',�Z���L�ᱚ��B����5X�v�{\���jћ�O
��2��k��m�UUdJ��]؁�Xym�Qtv����q�^5�VY�sz�59j�=<XN[|mVbJ�m��fA��=AP�ۼo�4�wZ�U�A͐@�z���Nd\���7v��   U �g@�U����A�����Q��g5U/&�u�5�9��8��y�td$�W����,Ĭ�U�{;�j{T��x�imU@0�����x5��5b%aǽ�T�ј���_���Ja�@����QY�k�c#cf�d��<����{w����;�^$T/w��5u�B��^մUm0�Y�Ap.�X	M��qK�������y��e�(���I�2wb �!r�l59�[^� 3�{K�2������H]��{������c;�g��Q�e����ڳ3�U  *�;\�a��PU=f@ 
�v�]Xp����W��
�� �   TU   
�*�PUU  �@
l��6ɺԬ�ov  * �U8�ʦ� TUJ�Ęez�@[&�Wq��9��
��D�ʪ�/��h5�1�՞V��۬@��اql�EVE	R�2�d\�M��z�*�WGu�� �  R�fU^�Amiwm��`7eS1���7�65P��lr�V�Ǔ��.3���������o5�BL��>׉H��垶�z�A%L��
�\
�'/ldK��^{ �	�����f �ڪ��Y���\�9�.[{�b�G�I���X�*����>aתjFx�C�v�[�l�̶1�V�3�MJa�C��j���Ճ�<��Z�;�ԙoC��G����$q���l�r��}��k\���Yi�q�zl �U�w|�wp�-���#m˥�zm��   U@���r�9q5ڲF-�q(䌪�Z�F��C���u��=}��\����<+��Ƞ{��&���C�V^2�<� �kB	�cV�H��}t�E[���x��W�'"�r	j��*ֵs��ڃ�H�ɋdO ������J��«��M��	ބwQ'=. I}���J���@�>hC]���w�������7+��e�|��x�P3ĝ�E�����BI$��k#�*f��q����MO���/`f�OqLx��6���rl��]�j �B��Ylu�-�B� �Um� *���M�i[��8J�XD�AUT,���[��`w���[�f�� io�x���l��@K��ɰJ���7�q���>@��U��a ?-���`X�Op��ԩU��ݴU�ɋ>�#m!��5�4�eP6q����O�������o1��)������u� zI q�%'#M<�-X?EZ֮`7��-�I@T=w�s J�u��WIי�W*���qj�bK��4��@K�v��DP�y�{����nW�§�'� p$�
^]ջwt @Bp��ӳj��9���3Ժ��ֺ���mqN2	>J�<I�p�h]�O��S����J-�<ތ���#݁C�����Uٹ�:��X�h�U�^�h:}��e�`�G(	j�m���$m�����Eo�$�!#�'S�,��rn2���Wٗ0(�M��UUU����]��. {Zl��I"^@7�z��U ��6mm�R�b)�cX��zI pڜ$�z�+���xO�:܂Z�~���\�x���& �m����cUt��
��P  U*���,�U]hݷ[F��J�U�8�X>T���
Ԅ�p	5��`]]xP���^p4�[k�qN��
"��Njޘ���jH�{�ޅqX/f� ����<Iۭg2�n�QM9b�������u@T�K *nFx�Ş�SZ��_d�S�-��v�u`���ւ�v[}�����K��2ހ�;�^$r���L]� 6��@y��>h�ˈNBs����rp�@������x{0��/=�"|�mU�b�4�#o�(�?�����VEUbQ�AOq�K)gZ��5���   �V��J�r��@�ݫl� �[3�m6F��� Ve *� �P *��
�U�� P ��  m��%@ 0n�ڕ@*���[eB��` *�*� �P ���c�A��4�ة(� �Wb���M6v%fU�pgz8}z�XA�UT����l]jGp6��S�cNl�֙YJ�n�e��w  *�e*��U���&�[{u/��m��{�}5*�U"ʊ�Q����o�jFp���{����Ά�%�x
�\�r	l�D�z̕UV�-+K.VG{
�5-z�/ԑ`_�����S�V��P����5UUTbړ^�$���*]�����nV�;�T� �#K��t[�5n���J�q��|[|�p��ᓾ�%��n�i�����Z����{� dUUEIÂ��8��X��tv��ۼ�S{�/��e��Q��|��
y���U[ �F7WUTT  �ڠ�V��� ��l��NY�/\��*�J���q���׻%�Aݴ@��d#o�J�n2"C�kf��#�%�B������Q�r�S��d������F�ZN8���Z７yێ�6��z�p��{��Y�oP<�Vk�TX�0���f��w�\�v��DmX���87���Qfb�ں��@�jqF����ڪ���2Y�l�^]�
ao�� o8�ҥ�r��J6��
�0�;�����l���Md�p��b��s�=�oY	�m��r�eq��nٍ�u�$�
��bE������,���
H
�"��[�� �*�W��j�g��m��xwW2���w!�A�T��v̉!���̒�n0{$��kƳ��xߎ�kΎӃu��R���>��s�AUU�-s�L3D�t���c���?l�����8��oy�Vm�DHpo��:�m�F�@�P��J�u�)�M~_w���\�mY~�Ds~�+�	F�21燐f�i�=q���W'�� ��,.K����٢�����{��ͷ�{$wD��Q�I1��Ǎ��7`�a��@�u����F�&K��.�qR�^�� �jqFݝԦ���$87�ā���m�o}�T5��M(�l9��Kj[mP�&�lU* 
��
q��{�y�"��Ll�C(T�R���R�u֌��v{s��+�֕=$ӝ̹x
�N�Z�7!!���eq�Zu'��}mګ#i
�/.�$��W�)���iM[�^V���H����hd�ڕ浙��v	_<���`܎9���c,;�aMo�6r{EÐ�#����3�Hpw/��Q9�֕.��ܻ���c�iEP}�ҍ�ޓT}�0Sa�i냖Kd�j�\����VBnb�|�Z0Qz	�P��̅�"��G=%��o����&�p�@Pn��{�g1��G;&�y��eUw��y�l�U�"ѵm����P*��UF�l *�k�����T�:��]y���B��:)�sޝoG�ͫ��ױ��{�0tٸ��I?n���q񬝚ت�U�.A����MtP�o�&�5��j�m�k�xт�[�z��k����ZS�V���ְ&�c�� uUUp�B��Y�ܺh�O{v��^j�|��*�d�I;x
�{܆V��2"y-�^V��P����US�8��I 9 ��j76��v�{u|�q���]u�^���w�1�ͤ���g�N�����f��퓼�q�=����hv���I�q㬈���0y�ێl^:��ﵪML�!6��|��K�*�Z�]r�s�����k�]`�\q�Ğo=�]��:�C����q��ﮱ̻�]غ�z�s�^ c�{�z���v��ל��f��w��6O;�{b<�=$��P�@?/��������KO�� $�x��~�����hp4�~Z B��;:�!	>f@B� 	��8d $:�IFG9`������d�
��o�d�I���������O���O0O�s�5��u����:?d:'�f�z	 $����|<���$>P�R(I�ȓ�$ ���P�������D�O�>���OA�>?�$�~�?D?/��Jp%!>�>�>�`�~P
�} |��e�׽�48$O���>��c�!BB	 	a$�0�$!>Y	!��p���|�a���~��~�� I=Ϙ�:>_A?y�?��0�=��;	����������'�����> �@	'�Ϋ�?~��?����}SN�`P���P~����C�����q�w����}p ��>���"!��������~��!�S�4�@$�P}� ������ |K��(}�)@@�Xtu������0�I�>q��X|���P��aЀP7��&�i8C_�AW���$�p>����>�I���}�'�>s�����;�}A���@����~����?�?9<���@�O�$��'�����@	'�􆟡�������� ����{' ��$@�iQ%���>R��~��a>_t��ÿ�,$� ��?d>���g�}���t~��Ϡ�rIC����D$��!?	����@?���>@�O�>04)��}����O��hi>"""������rE8P���K 