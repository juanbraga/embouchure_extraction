BZh91AY&SY�����_�`p���2� ����b6;�}�$��U=��4JJ�H��Md(�vҢ�F���D�U"��Q�(�*lȢ�Rɠ�Q]�UHUR�QUR�I]� Ԃ@PQJ)
!D�E
*��$"�D�TD�J��U%TUPJ�����ID��  P�R���{��W��ͯ�ݶٴg�^ƏZ���7������ƼlR��䪧�zW�xsj�]+��wE���r�����k���pS��V{��C�B�Ξ���_r.��h�*�Ex�*��P��RK�{��/n�����u���3f�=c�=bJ������v��Uϐ�h���c�{S�j�y���y��<�:K����^<�B;ﶜ︭�8�� �������lִ��;�d�6eHS�
w�q��׾�J��7w��l,�������@�_3ް�N������i�a��x������>��}�w�q �s�P٦�y���7��A�1��{Y�4��ʕE*�T����DA*R���m}ֆ��g�}�t�<���s;`:� 3��RT�z_=��k�;�˻���Ҷ��<����J���}�����ý��nw���|�� =|l�}ޔQE-���e.�[Ty;�B�) ��|�*�7Ғ\3z�}Yy�R�'�\��x��m�Z {�v�}�|���;��$�O�c���&g� =PO���Yl(�:�,5��}��<�P\�\}��`�֑P�>B�H�*�*"RQWĺ�����P�73���4S�koc���P��y�����T;�sǱ���V���Х}}���ۍ�J��ѽ��#�}z��M�7Y�s����o}�-�(�h4�� �}����>�=���O�v�4�&����r��wzk}�w}w���{�Ry�7o��
��^��>��wb�۟}]��=�ݎ����
u���ȩ㽟}������%$��_ �JP�E�$D������{���`k��Oa@��"�����mꇡ�:q�X�7��z�ww�=7�'}�x��|�/t+���v',��z{}��9)�X�����)%V����N���G����¤����n |v��׭�]��=�&��w����{xu}�T��y��kt���}��� ���{��	��{�|��ﻪ��O�|��}�7�B��*��!*U�ʤ� E)�)ﯹ��E��w((� �g���� �M��4�}�K�!��4_t���umW�u�=�n��]��<��ϪQ}��o;_`,�[���^��[b�7^�8mm������ O�	�*� 4F�*�FI*� �d  h T�!MU*��    ��UQ1P� �    �?��RF   @ziT�h�4���a�4{Jzj{��?��������f�#��_�S���VUY7���ƞ���I:N�����I:N���wI't������N����$�'wu����I'I���/t�t�����O�'t����߯��$�'ww�����}�����7���5�|�ߏ����u%�?&��ο`�L����C� �^��>�J#�)� �dt�2�~��]~�]��}�M���:g��^�}���vm��P�e�]������=x#�{J8���v��畑�`V�P*k��wƞF�sq6�T+l7YA=�v�{���Ld�.��̒��W��S��]l�竛�#�K`5�3�w�e���l�X���7K��N8Ջ�R��bTWbOM�{]t����h):�k�u,��ΓF�7ߦ_8k(ʔ"����e���ʺ�_5���q������O)�
V�ȓ�f�=/x�J�H.�B����1�����C�/:�)������A����/�$
R��A���l�;.��O���EMش<1�g�3Ni"Ir�fc��q�I�M��[�o	��1�J��/),���!�H�Y�ty8��D6���N��0�ܢ�J�ʛ�*�E+�y-��b�����]/]�4O�޴�N���*>CI`����m�[�^j�y���5[N�],p�v6�mMZ")��h[�[�iVeV�Fi��Ѕ֥�0��)��4�j�ݣ��,Ĵ���0=[���d��Ⱥ%�I35j��	�����z2i��㣭X@Zl�%�9u��,�l+YYB���]fQ��rџ���Dv�����ɋ��%[��tu��8�mz�A�]����oX�&�O�97��8i�[Zk+I� 3&�tF�Ɗ��¦ԥ���p�h's"rbU7�-�v5�Q��YI��.�R����Je6@��{YY�PYb�R�{�+VR�hx�G�~u�I۩�.�֌f�Y�!���tU��ΐ(�U�Rv�v��� UG��g:�� Rr��bȧ�T~��Qi��s;�)Y�e"0�A�R���5�P�L��Y+�?-����#%�q�u���Q[�F���'{��T�V"j�e��+�7q�v㴑�̔�S�oM�'Yv��2��s(�P�����:�%����;Xr�Z��M	�R��CDna\�G�k0�aދX]<�t�*g)=f�A�{���m��-&%u&��m��b:i��m���f�90Jf�<���[4H�Tn��@��]%�F�h���ifX�y+;�0�D-KMDUŻ�N0��5�3��Nؓ6���y������2�ˬB��5l�a%J[i�[�=@�e�ZI�v�J����Ѡ��i3Q�H-�@�]��O�=�in�0�o.2Ƀuv`��;���K1���YA�x����PۡM0�S��`��Q�`ɸ�Z��IGiJr�I�ZJ�]]�yFg��&5t%=�=XJu�\������m�����z�#e��Ѧ6���yq,��SN��`[u���.U����;��tk��,�U��k��;w�L����J)L���c�Z�n��[J�ߩ�jxظ� cǂ�mխ;L�8BV�z��R�2Ϋ���0;ő~rfZ̽e�t����-�����{�<B�dS�Jvm�m%�M2[v�0L~ 1W��iY�z��[�5�r��iuI�=�j�V�,
�ʖ���K�f22�]�>����}�c�8�g����wA���ס���a��t+5��4�*Z�d4�v�JN1����T�.���!�ʼǺo6�l�r�`�U\�ia:�V���p��A�Qe�N2*X��멤��<틖���A��@�O��>G�������S��\��N��U���ܦS��g<��i�Q�ee�r����\�+(��*�K3(V~�Q��e�P����������>�)��\�v�\��m����6��C��^C%NmY`�j;�ik��ow�* �v�Н�ll+L���F��t3I�ع)7mJ���2�v������+w2� j�au��ذ�3/�7L�n�CV`	;z���952t5���V��2�9nhK�ӅM�?�Qk����*�

��0S��3u�kFP�	?e���G-j	%�)����Yb����U� l��$�2����al;��n~ �fы#d3P��䡴�Ӛ5
r��e�v��wr�^[r�ȓ:��ǈ�/`��M�;jdY�4��ӦЊ!���Qn�IL��nf�i�����OSٚ�lj��&�E��*��o�;���j���v-޷oD�Q�?�J�!n��f�J9���B�Rdt	جe)�+���M�D!b¯�+C�K%�E������K4�ʳ��	z�Gs�m+8�#qҒ�jVJ���ִ��{�qǖ�B-�*��kZ^ܽ�P�e�: ����s1��o,��\���Zc)C�`%����?LAI*���gC̬�۠��`��D�~	��]��e6��%;j�1F�Z�v�J����d�Ua�۬o&ų��,��f��E�N,�v6&��ڴ��0Kx):���2��6S&j1U�45�v�d���ׯu;�Ɣ���x�5��]rîi�S.è\yS����&fT�A1���>��?|C�4YG벀�)�� �L�H}�o�| _r:���_��~n�~�G꬜�h�ǻ�[���5!��No2�XQv��r���m�œ!1�jڇ7X�bGFѦxt�����b�>�˅Ō �9|��X�U��d�P�z;7��!Հd�l��l�E����#sD= ڦK��{�y<n��+�a틫V
����WĈ��8�&(GS�p�Gb�-�yVWEm��Q��R�[5ߺ�KSb�{�że�T���Md�4��꣑~_����S�i�f�hs;1p�˘/FN�\� uV��I6TP�5a�p@(���ХR-&퇍l�b�Q|+�
��e6�9hg�ɻM���u�o3p1�`�t��o�m*L�˿J�E}�V?_��[�U��ڬ!'�4��ojod���
�8pH '��P�}�VںV�Wf��utk8V@�$le��F�.<$sl"Ѥ��R�V��1��Tz�]���z�V�B�����N:�y�s&@m�)R,mԽ�.ż��f6�q6H}��I�Hts��G[���A��
)T.�l�!Rm7sF�zڢ�؃ �-�zRP]�*��9�`��_ne;�N�R�?1��#��D]�������x���X8l�(�)��8�6������k���ͭ"�
�1,�[W��!��5N2����Z�H�J��f�G]ۼ.`��x*��:N藃m�=!��(�<��+@Ʋ�uz���h�Y�V���de�6n���4e\њ�I�G4�ͫ�r��4gc�̬PP�z�!�HC�s7mM�!$%�g��d�.V���1iOuZ���R35��8)]^���t�M�"N�"ď�bYn�r��$	��W�za/���m���	�"�*�j��1m��A��xu^��)ފ$�����|T� �w�V�U}\���I��h���ņ�P�b��M泯K�h�IX�*�D�d��I�	I��L�c�av7�|F7���yIf�v��aUr~�[*~DXU�Ʒ�#Җd���Y�FL��P�k��	�q��Ʉ�i4Ƕ]� �ǲœ�D�wT)u���师��TJ8�X�e�̌ ��TalV��9�S-�����{�MҼN�·h�#l�qU���Sow]���I޽�m^�V��R�[�e�gE�.��Zi�]�U��jtF�:s2���� M�[��ە�N��m��3��K�1,����Jk����#��>��?%�"?�Bv���5Uq�V`�'s��{J	uqؼa/�mE,&�h��Zr��4QШ����o��:�h�Uf��ڂe�B�@��7t֪i;x�k����+b��تǰ~��u���jxD�u��Z-30A2��6�.�E+4K�jGmk�a�C{�m<鴭��cI���(Z�i��DV�{Q�aN�-�y�]�gAB�3�Ǫ2i)�%�9�
����y�^&�D�hoXj� /B�c��5
��7i�V��������d=D,���x��;��):tkcø"FUꮄ=c�;���M�ʴ6�d��I��A�:��c�TT�^%�Í��ׯU'��"������^�U��z�e�۲N�`Y��^J��36TtULu�G�����KT���%b;0��.�y��N5#oҢ+�"vB���u���r�%jl�E�.G��N��,v�p&�=�О4L0�GN���e�p	"�\nP�M�{������q]��js���z����E]��ڃ0AL�7o0�)�y2]�ت�m'I]n�^�9��A>��h�6Y
��״Է��MS��V�/�����(b�@`��)�*գ�c��P�B�1�6u�չ��I���yf��&���� �n����c]h�9��������Qi\(��F]<�M^ѧFSؕiՂ��#���h�Z�kP���˛6�e:RM�e��\F�� ���7�mK��lԒR�u�%�15eIG��c8�gu�Se[���B�L��+q�o*fU֠��f��E ����m��Ab.��o�oa��De��Wk��ɸv�`�V��ɩX(-�i�2l�l�
"[��*X<�L€�WÂ�D�.Z�Ǎ����"35�-\j������,H��ݚ;qd\�ᝆ��Z�n�e̺hb�x�:�[_�ȵ���B�`�����͛�2��/�wq*3�i�����"~��C�����n��;މb'�� m-V$R�ot.ob�+�Z*J�V:�c-���3hjǙV岓��-�Zi�\P�IF@ؤ)>����.�x���3+v+��t��e?aQ�.k���6(��O��3�����
5r��jF�(��`U[�s5ݲ��
}N�8����������@�6�H�²���J�F�Gws���Q%mم�P���J�x�Z���rp��FDF�o���p��]�w3���[U2*�Ր�H��M�x�Y�yI�}�ջ�/�Ӑq�r�1�X,Til�{��Ҁ��;e�ۘ���wN��)ne��q֊C����q��1]w
WD��2�J��Ssz�]9�a��3z̴�:�'[H�v9_/@�칵���{��ռ�r�9o�G��T�X�Wun�;	�"�� 9[���հ���P]'�s��y��f�sS��~�H�E��|��M�3uX�w�ڤ I#ں8�zoj5�{����S���_<��øN.ŏ������IBբ��2��މ�����&�Ƴ�(ŃW�
�B�X�ƽtrf�A��in�efD�n�r��t�b���N]��"����-��y�!�0S�$�vl�oz~��g7��tr�^4�J�
�T�D��,ci �"�L��CPf\ܽ��w�)f��O��۠U��0�Ê�S5���.�[(���*�HN<��
�������ۦ���� a�H�r�7&l����jT؎e�m�*�,���
%����sCz��y���h_Y9�T�Q��:�Ib�:�%E��{�Z��i�{x�%���lQ,��9N�1�3Yu��/�@�S�K�ڛd�J�en�����(�Yz#� ��C�Cf��J��^�y�i5� IC_�&U2�wN[��BM�n�� lI�1,CU�f���q�,�%c��jax�ΗZKn�[I²-�5�k���PkW ��lމ�oq�����t���G��Z�[F=u�j�.���n�(C������K3��F;��mP�XXu"ygvj�.j�to,Ԙ(9��k�sHt���#3�`7x�i^���N��H���y�7h��Tr1J��w����F[{��΅u�fn�@��^�ʚ�إ����s�����TY����V;Vg�]���f�.�!W�*7/Q� $ڐ�%��������lV���A���V���U:<�
C:�'d���-��4
Vh��!����f�Ǵ{uo�(�\6F�wa;9R�n;G\��34�e���m��J;�6,bނP/%�u�Hv���]��U�WE�٧���bam&�T ��JJ��2�
�%�À*F�#��/[�����A���uM�G"Z�&�a��A{�uq�MVM�$sX��M���@�5��رR8��;��
����Of����ԳZ�䡎�z�\�)�,4��Tķu�i�����_�N�%��Vjkz`�pRER��-�r��DZ��+X��N	an�fU��]Ib�$*�ٻ����z���B5���wU�Kj�M�1R�&m[����.�E�n�<MEmѸ^:��3����Q�l���%л"���^A0#Y�֢��4XtOkO�]�`�?f�u+n��s�Z��GO4
)72�VLZ�X�'.F+`+MAe@�L�sP�on3�:+?f։/Ʊ\�t�K�E�y���S��DT+�n,�ј�H	J�D�GS�+�����-]�=�F7W9`�`�k6��o0DܽJ�H�$uݣ�X;�Ø�$�;n�N�[�P���sM�d�6���U'짩!����6�ʹ�h�ݢ�sYz8�i6v��/2�h�ט�p��ڙ�v
��R�����[������n?٢<�:eX=�F�MVX.�������Snf˰�(eZ.fQa���
�Y�01+R�;MT9��n�õ�ݑ�#'�D��mH�ۺ��akn+��օ%7Mٙh�^F��DK�gVk�XSJ��:ǆQU�B����A��p�hQ$7�F���7u��7Vk������Րx��ݻ�-��2��3mVK{l�,��P�9�7�4ՙy��;�Ֆ�W�M��mΦ9�ˎ���-X}���+���*v=�AQ�w��R\Y��w!J,���'��1 �3�R荖@�Kou�,u�C��&խ���t�Sof�V��;9ü�B�u��]_�`���ܼ��jV�����˺O�Ж-2F���ԫJ�UQ��jBjWʓ;+b���M*�UM�����
ꪠ*��
@�모�#UU�U UU\Q�UT�uU*�UUUUUUUUUU@X���R�UPur�)�UUUUUEU�T��UT�uU@UUTUUU*ҭJ�UZ��V��������&F�������V��iV�Z�T�����R�HMT�*�U�UUUJ�UUUK��U��a�k�檒sP�UU�U*�\``�<�9��vף���P�f�$,�Ɣ�m���t���^W�[=F�c>��4+�9t���a�ٳ��"�
\�t8�+��f�������qm�cv�[/��quv5��z�7���0ta�U�s�;F��ӈod〥��.�گG����-���n��dn�;�D�Z�pf3!YCh�I�&���"�f�%3�g^��)7�R�兖ɸdF㫓9q��\l��n�[b��;�����b������S.#e�����Z���-w[�n�x�c�R��7Aַ�����6�l�@N���"ϫG�DE��e�-C`p��&ԍ�1:�+�u��=Ȝd���ӵ�YwMάm�h;3�S�7[C�������뗫Ƅ�m]���q)�Z'�YX�kl+��,��7V�+]J6%̮�[M�*�%�	�ˎŅ�����5��Eu�l s�m��8r�
��5�3ɭx�W��ƚm�F�S+`M��@��5�)���WEGGK�E��l�NK�,��%$�5!����a�u�V8m�b�ѐ.pР���q q6�Z\��'I�-ãZt�g]�p��A���u���0��ia�-�砘�v3r.
���/N����.�Cϟ'; ����h�4Aשc�\i6tfTF�Ml�Q�B�e�����cof��.�ٖV޺Vk�2D5i�-ؗ0�%�5�w�CgΓm4t�=vڐ%S3)��lë+�@t�A���%��6�����	s-���!B�зq�-��p�zrxe8��F�P܁f��u]:.�+���]b�m�yS����n#R�p[�cӌ-����v�,�]3Bk5�ʥ`6�;��gX6�8[<Z�v
9Z�c��;�]�9wNku����n�S�� E]��cu�i/:�E%e����%�Y`ZX�,�F��i]���;^V�3n��
�eۭ<�a����x�-��q�:�F��CZڊ��nc0���1�V��[���}��焂2e���m�,�4TD������I�Rۃ%�]��J;+6vݲvk�0�=�k:k�B�4� 7W���8i��Cp.��<2l��	Q.��Xóv�B']Hӑrv$��E�Mx�;g:�L�ñ���o��q���C�w.	*/N�n�@�<�ꃷF��hu׶u�!h�����6��-K�����Z�!�Wl��<Ĩ���⫱�X�V�t�rC�v�N!��x��DA�i	{u��ĂK���4ح.���i�{K�����&�h[��6��b��bb-��a�p�^+��ٔRؓv���F��)��0�"9����(9�)�Z��f��6rG�%3�+s֣7	rl*�ɕۍ��kMte�6v�#�{D����u��W;�=Ɛeq�٠����`Lb4��F6;vj�L.^�{:N�6�{����;x36#7SW,��&��L�Kmֺuz5kogkǴمz^�7=-�Q��o=�Q�԰�`m���-���uZOA��	9�,fS�/]�]X��F�����F��r��Aú�B6ݳ̒�;�:�u�2��u�-E�6��ْ�)��[\�{4nβi+�X�n,vB��T�tu������/jw!A�][$g6��j�v:|�u�n�[��w8��4c [p"��b�z�d��x��l��/F�]��
ر�Ee�E�k��\L�J1�@��=2Yhj��퀛P��������L�qte=���:#��ش��ݸ�nN�Zu$]X�!�F��e�#.��hˮK+5�XM�X�H՛V�P�����r�m��`�n��ص�%��Ӯ���2�3.��u.�SGB���ʋ�.�H�$D���0Z�0�h��\źm�q���%�MJ���F����Е���۞��/�̂-jE؛XMƶ ��u��"�mric/�"�L�K!�r�V�(T�G�.,�Mo[bE݊iq5r2��}q]��N�
p-s�x(��W�+5��IF�!KU���V��m��QJ�����{��6mH���ɓx!ݚa�w;��n�On��'�f���\0�l��3���v�c�,�̱�̶X����*�k�.N���sd#e���R]G`.ە�n�dЍHv�-[���Ns�a��n��jX��ڮ�Gq#���-���O����X��ٹ;#l&��\��םR]�i��Ye0���G�ܚmub����暷�Rk,vQ��u���js�F��l@���͍����R�:�9,=���4��e6�U,�`䅔��.sƬ�hM�� �`jf�D5Y�Ma�(Rb[T3)Q�kI���_�(e]K��Ym:Ҋ��Y�RK�v������������y���C�j�us�<�v�k%��u�/��	�їj���Q��ք�j۞�H��������)�4��V�ieλ�s`�S��(CB�Yv�8)�X脸��:^МF�l��4���oq��Yc��*�>
MV(	l�ź�a�u!���rB�z��Ϸ-���Y+7dv^�kp{i��;�+�cn��D�a��[�[��95OB���oC��-"�b��u-��BWS�D�|݆�i�.0ݻ\܅��tڐ��U1cv½2�'m�wYwW��0B�^����	mV��@6d��ƅrIvs-�Z�As��8H9�ր�u��AnvްIIJ��Fmv��T#[3��MF�v`�T҅��4*b���,�1��\f���`���� �ǵ:�j��Meb;S1�x!ݚ]�t�{���m�S�3�4��l�nrmֱ�(\ƗrF��:��%�!�sy�:�x�W=�g֡�Cq�Z�� dyve� 7P�e(�q�ٙ�9�����
\r=���6!��ܐ��MV
n�7]�B�O ��VMN� ��6
�IQn��T �)���p��F8�\[�,Ϸ���.�OnB��Jnô/j�^[(O]  �l�(��[��d���#ٹ=��s���NR�G�qo3�6�w3�ppRbt������ϦLr�nj���-]^v�.d֖Y�4�	��i@�Xj͑����h��5��&�Z��/,Ǜ����m�C�r֪]#�$�l�A�i��#n]��e��F�mD0A��`��C�g���9;r�ʚ)sR��
�YR�+�Zlg��v�pn��.SB�j�\-�	vk�Բ����p\^�g�C�<�����G8W
s��A9��훳S�2����Q�z�X�`/66:��L���������0t#�M��趛8����ȝ�;tK��"����GnݵԜn:� �AuşwWv�q[�'��c��h�{qO�tv�
�vӎB+���#o%�ԥ���-��1��fj<�`-�[���
Q�Z��h뭱�����K3omθ�6*Ō���f�4�m�%)K��(E��i�T�@�]6����e]��j�Vj�eH�Xg&�Y(�6�n�n!�@�S�Էqĸ�T����R�ui���x�z3�W��mh�ͳ��8,5�m���M�+&�)o�ƛh�IBin�)s��c����9fWh^2b�W]n6 �˵��Nx�Ƴlõ!��Ve�-�X�l,�[,`J��憸���[8AK���m	�����{!� K������؅M4��F�hn�ڼy��sLsn��z�{N�5���[�8ќ�t;XCL܄
VƼ`:��֫0�i�"뫘�λ���=tq��<d�stQm��f�D�̙��nǬlu�ь�"�Kn�d�F�:)ٻ��)��Ÿ(�0�ۜ���u!m&�`�.��3Mi�n&�U�`��	���-�6����Gvd��e`�̦�쨰fw� ��klx�f!��fꂔѥ5�+�T�K��2d#�B�CC�N`:��Ǉ,�j����͠<�k*�԰[�6����jL��t�����Jck�^\�j��s��Q���������>���l7p�\��b�����v��l�E�t�A����n`9y�p����і�4;���iu=]�m���u�
[c˥,,�����v.�-�nX��`�宰L�n��]����S#s �iw%����b��U(���e*�u�\$d���k�:����rъv���+�1Q�xn�'l�l�v�-�U�#���vj8l]\��;	ǒS�lG]������KNE����m�9:5s�i�jLt�ZK��6H˙���ː����T2`��!�)\$L�չ4���mV�������SM`�Wdt �CR-����.�MksI`�Ҷ9����`30+���k� W$��)b�,A��\����<�-�-�nlk�۔�zUr����\X'lYa�mJ ^:�{��zxp5����n�n��m�=v��hV#�v�)���s�N��M����ų)0�B琺��z�6�l6ݪ
���7OY�2�,�u�:(���Q�u�q�8�`^�S��R�q	ŷZ�ܚ��3��Wa��:;����Fkq�-v%������1�;^���v�k�=�4�Z�E���ne�3H���6R��b���x�������'Gn�Zz�y��,t��4�D!��
jI��Ư���Q�X�10=���vj��L>q������CԶ�CJ� �V�����D�nل��A�XR�8..Kt��Kw8^5�6� ��洘儩��V:ۊ�@	eak5�V�Fۢ�Ŷy0���-kǭ[��ns�������ݭ:*ؑ�u���V�n44/��'N������t�������O;�����I�I�;������I:N��~/��}��ϼ�>�'wI��N�����t���ӧI N����8;���;��t	;�t�'t�Ӥ���:t����~������������TH_�]�'s�����ǫ���mR��mJL2h�pz�S�D.^S��	E�7��9����a� �H�<f�h���b�O�r��=�e��:jN���J�����rU�ok{�ݻ��ϐ:0hq��@d�xm+��t�:��p���Q~�ց��o��Ǟ`�39z���п3O,��"��J�+/����%�s��)FD��T�ćG^��Y��n�)����j��s侠E	ʝ��'l��x�kg#o0�tFX����TI5g��W����^�1��~�	ޤ����[��ռ������]�����CX}�7��T]�x+5t,Ұ�s�ǟs]�[��mZ��fh<���v7��c�,��w�c�G���L�o�w{�ual�JЃPm�S����k3#<�ԩ�J�m��Af*�����կ�,{��S��^�~~�}ko�%����������۳2MǛ^���H���"�6�wv��^a���9�5y���{�UƐj���G=���4��RXY(ժ:� 귊�u���jS���+m�ʱ�a��B���[�936��[Y�;�μK���R��]��q/�⧆J���2�MGBl�T�L2�������adî��H��ͳn�XgSp���z��ugw'�ma�f�k���M?[O𬈒�Zű�����n�YC�0׌4[�ې��*�g�������v��-�:�dś��Dַ/[A��G�=b�
/�h�&���FY�l�鞲ڒ:�nƛ�1H�Ĭ*AJ�#oby��<I�u���t�Z	�.i.�ś	�X���L�ZJI;;�X<יX�5�3�=<3��$~�'��N��ǫ
�����_����=��2����˹/����!0@c�t��W^r��8c�*��M�{����+o3���|%�Җ.F��4e�iX,�[pIMՌ)���nt�RTe��S����o�{���ɞ�S�c�[���2�y��G���|άә,��Q��rv�M�un�z!�v/��qU�:�^�ͼ�W�Eٖ��諵�ר_|�M�����|�!���`�YA����QUP��꛷����W��'���6�\2�KwӾN�׿=e�N]�<�Bv�E8.��ṯ՘��`l�
�tyB�)�n%Rx������x��#��8�p#~ݔ�1اŒ�E��;v�y��}�:��S �߹����M�}�����b�=������gEꗕ*�J�|'�����X�1wq��0�J��n�wf��1��<ͩ�C���P����&��FS��\$��[;l[��WJUX�����;z���<�*]�W�|�Y\�����Vy�$_
:Hp�$-�֓���K���t��N�s��>���X���M��2��d8����^�&'�E�����M@�0�M��]��̗��2Ɗ{�����1�۔K�ZZ#�8K*������Ef��xY��*)*Ro�����0\��ޙ�ٙVt7��v��,R5�׹�;2�{�6�e��f��?�j�^�{�\"
a4*�u��^6dC��Y8�gf�s���z���d��̒�����g<֏�s؟�L���\Z�4s�%[�r���0�p����"�k- �ҝ�x�\�Q����)��^�	�zӒ�N��6�^��ڻ�ܼw͞ǧۜ���x�~èU��IY�9�*�Q��`r��*e�u�������n|�̷���?|�z�l�L�����)�S��u3��6��<�uB)߳3"� ��@�sx�E3O����n��&�9{�^-"n��L]�J��u��sb4t�ll�Y�Â"�̭؋�7fUq���9��k���h�t�qp��O�c��{��Vq�d�ƹ��r���ic�'d	[�$�]�6��ԹNǪT�P��MU�A�QC���雒�F�Ͳ�y�/�����9��p����(��Lf��ײg^d��j��f�h`
;���!Z�t��i��Tn�����3:�x�{w�栦�	l�I���Z�*c� �R�Q�5��)^�&��-��~��;�/��'E=��N�@)�P�����q���3��$� �B������\"� F�ڨ�Z�ӜջX�L_�އ~ˍU��f��C�ϲ��m/��va���u4��[�~�V�B��(� �k��{9m��s5���o\kz�ĭm����<�&7J�"���jЄ����/g���E`�[�&CA����Uͫ4Q��Z=��Su��$%2������b���:���W�	^��p�d�E���\��((�рC|�婏��y�lS�J��6+}q��%��=�;��9��7ŝ�����\�����*H�D^�o�x,�qv�'k��~��:TJ��&��b�3	�
[#3�WC���Ս�/g!=�+����ǽ�k34�,�DfC.Mj��=l'��ܻy��jQS<7y�9*����ˬӣEp����%E<�[f�.���5�����1QOo���	�%=��ϫ������['B����Mky!�����5z�P�z�1�������*�>F��P���F.��#v<w�zM_�b�(�A���o>�	��/2�<�����{�7+���6���Z��&&�ŉ^s:��^�8��lk�ԗD�&x�hJ��ü��׮U�؅wC��'s���s��.�֬79*��f���n��[�%��x���%��&���w� �']�ώ�|��Z�h�C���^ �p�rɗj+��.�0=�WA��$�@A����.�m���o8";�je=[�5Z۝[��R^$�����{�A������*�3�����N<�;���w�N
Y>�"���{�׍�7aTg���8Y���v��ܙ(���VJ�E�Ow��z!=gP1ƬYT�X�=u�z����n��6xX�Y˸�L�U��M,�ښ�c�YŤWS7L� ����]�^����_�U0���#�}��O�?iJq�7?�ͧ�[(�]	Z��gz ���o(^�U�5�j�s�B;�7�fJ6�`^=�kk�u�6Ng
@��ɸb��u�Q3�06`D��I`"���i�:=q3Ɵ��<�o�oQ��a+k �l�z���'7v9zJ�Jqv�\���&�Ŭr��\6,�n�Cԣ�ź��݆����\m��`HN�&�t���p/d�u�q@���S.��Y��1\*]��lr��^h�;�
�����(��7�)�C�^�l�wf��r��i�b�3˭nָ�b.8�,&r���N��m��R��:��X�^�_z�w�"ň�è�{Y��E7čM3��u�4ol����'�Ҟ�)�5�ҭn]����.̙n�����B����\��ήy�`�qq�������C�$�ݤ�)HT�W�m�������u�2V?����$��@�Ƚ���@�I�v{$[��L%��@�-�(�2"y��$owq���?�Ƶ^�<��</y�r�R:{˹/N�A�6d"&�A��l̃��NIt�|�C@�O���?��<�\�E\�AY�stL}1nN9�ű	{��L��4��P"�KXjq.[��9�ݼ�ɐV�ʴ��8�꟯n�����\�9�h!�%���Ts�����BoA}ޠ�1�g#����|h�h*T148�k$����^����`{�������C���f�N*�A�˪+�۬�.Θ��f����48D8,A�4��;B���T\A�jn���џe��^΋L���.���0����^��1�	��j ���)qEAw��*O�s46�쫺xf_
M�"����;�v�d�gP8v"a�`�Rr�"J�Z�x�g��V�4���SsR�)_�Q��uf1O	�?�7u�e�.]-���saX��0Y �!x�]�V㡹�:w8�W�\&���E �lf��v�e��lu��Ҕ�7w�����V��G�ь��p�>��ޣt!H�Hl��7%�P`�i��T�����
�|u��1�y[U�"�� �Ǩ�����G�� JΧ��+�R� ���Ud��t�xJ&v��.𮗤�lw�q�	�K�?DV�gss�_G���^��u�b����,����犫�紩�Pd2�n��7s&��zj����֫P�|��؃��q�$�k�Q����k���j{~���k��"��) �V�`%�!I
EE��P+�n ��mЛ�GM+�޺;Ң���S6
��[Gs��1�6%�¨�"�[N�Rp��(,�֬[7d�����wz
^���Ə�*����������9�G�Dt-�9I�F���[7l�Q�U�AË�A��0��	�܊��g&����'����/3V�񌝕yu��������=1��{[mO�wm.�*$�
�Vܖn���h�l���.�l�@Zk��v
���h0���-�g�������@,^�EuFTj�Z�t��΅��h\q�B�১2s�MB��w
�$�q�G��+�.,����c>uk)
�mm�û�|*p����&{&Ë�+̳��{� ~7@�<���ֈ��� ��	���<{��)����1s^:/�o6��Q��$�^ged��}��S0�e5>چ��fƝ�ۧ�q%�={e��%��ȣK]j�WZ���_�Q�2�2�ξ��^�Ȩwv���$ĉ��m���ծ�zϞ��s���3�,�����V;V
I����t�JewW!�
��y>�h�9W��Nt���Y����M�j�y��ɠ���o�ks���s
|�{�__#�۔*+k�X�>�ˀ6;=�5�9�ۍ����,&RE0�DY�-?Z�M4����q�.�wp��#\)��Z���8p+�	6��Utc���+9y3`�9�K8�{�x�pY��3���H�8d~�{2�n��rޥK��C�{C�|_k����TH$*W.JhߊrG���h��xGN��˺��rkD��W��|��3�ͼeY������f���7�;���GSj�՛K�)#�)w-su���I]z-�_�˯-�S��#h���Fg�e�)�㤝��_yY�x���Q�
	�ʂN_�E�{a9�3�i�SOt�]���V���ԮSu9>q����k���;�6���UqDb5���1ÏYD��H�7v��"ᎂ�6>���E�� �ME�ou�7�-纭�y�a�'у�4����}Ҳ��q;�WR�i6�_2���M=Z�^%� �{�j	�uJnşnB���%�,"��	r<v�Ӈֈ͓Q�.Mv9�J¢�#V�+7b� 들��ɯyT{�S͢?;��ow��t
}��q��.����gSM?K���(���o�\��ٽ���Ze2���T�� ��2?g�^�=��a�d�2����3���N��$�ݻ���=�$�?�k�b�ѱ?�QY�,j߈�н~}5[��N�l��x�]�f�}[��E��<s�^z�S��s�_V��b�%�wf��c����@�ۆq��E���l��_9��w���^(~e�\pcή�5Rս��vԮ���<��m�,M	hY*�
�.L��CXT�o�
���� f;���I�׵�M��oc�~|b����}z�Q�[kGM��`[>���6�.�%�^��GIӔ��4N��]���J$�v�8�BS�hE�lՍ�X�Δ��i�]3)/iB���e���W���]�f`v�HQ�44�u�m�֚��;S�����Aű�.
51a�kupو�H� kpSԪ��ZM�ѓ���9��	b�PG��צ�5{=W�R�3v8�mDve�R����8"��+ٝ��+΁9JI[H�ʌtk�3;̆�k����!��� �ʸy�wF�ii�f`�r�^Uա�&n����VU= U��l�U��W���� �`�{c/4X�WM:��Z�۳�y�d7	�l��p}�ޕ�����~�vv*��6g�ֳW\b6޵юປ�&X��xI�#�u�xp�Xg��F�Ѻ�$ ����\y�kŏ8�q����o��;u��vC����yΙͩ(^WR����A �R�^���@C�{�9�VGxͷ�ٞ#2��ǃ�<��������Jՙ�i���Ь�ì��%X ���9�b�x�����5fL�Ö����/7���l+�v�f�I�$#��7F��s�n�l���,f?Q�tF���"FcH��/���2�</�/��1+ܫ<q�g!e��2���{���Ώ���~s12��,f\D#�we��0,�����C2�7���o^1˥�D�������t�]2|�wv���KC���"鬊��v�=q�`���I8v=�r���H=�+��<�4w��T���� ���!t���#{��o�ȋ���T#f���CaU��{r��+��*�e'öأ>O6{��`3��7�g.�9���ӊ����i��Ȏ^�'2���7�z/#��鋥q�aY��z��ޗ��Ǳ���+c��ݮ �.*U�&efh&�S ��8w�p�0r'OKb���w��g��X���y�.��4٬��6��Պ�-.�A9��x�[���Y���ゞ�Sp���^��I��F%��#b_19_��J��L���hꋇ�訛}&�����75[�)w��v_>�>y���=Me�|�Z��M��ʝd����6*>����"e3�g.Х��3G�+%�F�b�k�nk]-�R�Y{t����P=	]����pܨ��[Vu�M���e��ҏ@[`�:��q�ӭ~���^'�Fc�&j�E�+,÷��������V���~�bi�k�a��GSt�E��r�����P@��:4�w���Y���W�m���@rq"K�
XAc��]`�Ѭ�+�}`�6"��n�~λ�s%ƨ�M��7כq;�i&�*�a�.��A*���� ���+���/':�2e	:hwz�g&��墂ޒ"��Ĵ]C����永�k�u�+�Y��D���٭1D����sŝ�JjT�}� 2�]��;����`^�Wl�,�(�*�EZ�@����j�iV���UZ����U���S���:��-:
��l����G.�oe�y(�υ�amY��]� i���ć
����m�7e�䝷��Ʊ.��z��(v�ۓPM�p���Rc�gm��:�����p�@y�ym=��u��N�6�%��+,cp�L�Q�v�L	�O>�q�6���Q�-���j����*WT�Z���]vI4��h��B���������:�6�3�غa�����
��l�b���]�ۮ��bl'j�6�l8���m�g� #���W�L���oӵ��Ht1��pZ�E�{\�E�.���9��k)��F���lK
�6e�+:������Kѕ!��7h��l��8�g�z���$ N���F�1=�n�q�:\"֝΋�N�rusjmx9L7�щ�m��7���x�Y��W��7��OHn��a ��Rupq�k��Ł����Ƨ���vgӵC�7H�m�Ӓ�L�[�h�+�mWh��4;M�����e^%�9kvɌ:�#�؎���yk�WFۭ��9�E��ݲ�ut]z�9�j�f�n	Z����<t�QѰ�m<����:�VCI�x;q��p��4OV�!��va)iƉ�hWKαf�+c�^�p�0�N�x�c��K�^:���r鋓n`ׁ�j�t��2�b�xuق:��f���d�J�m5�,�w1����8�����&l��&!���koh���v�!�����^�P��l��&�ܽMt����[�Fy^:F�2Wk��C&�iM��0���<Nܚ���8�'�������bd�R�ʹF�C�h����f��t(s�rG� @�[-�H:��ڎubQu�/XB��6@	�q�5�u��F6z9:�*�B'l��u�kXiA+��f���͌�;� �X�)a�l�Ģ�YK��Ϊ�b{j�6�/,��.�%��d$a�$%�����O;��8�rDn���").enX�����%i+"��NZ���,���ޕ?w�`>�_x;�uۨ�ڷ�ި[��]z�ֱW;Z�ɹۆ"���:L���u�jﭺ�����_m��?H�z�i����/j��'��+��]�/>�\�ۗ/����;�s���E��$`^\�!�{�	�#MH���=w��!�u��Z����6�z���}�����{r��H���OiG	�_�y�gw	݅$b.?*��H�����豎ad�S���G/��ss׽/g�G[�����;[{r��m�Nl��ի�����[�=;����2�ɻS��^�=0��$�����#ɫʼ�D�Q���TZ��;/{n#��Wy�Z��c�f.,�
a���3�_�}��,5�i�Vw%�M�[뙥��@),�	�_�\��pX����{�f_7�ֱ�%e���� ��qi�
��G�{6���$}�3�z3,���t��{'.�qM�@l�Y�{�o�G�3|�"����o�&z��s	�Jc�R����w������w�WVFE:��6��ms�l@jY��.
D�Lf��]�DN$A��zOw���P��ɸ�f�ǵ�Z�W��T�!�ծ��i#�c�ߖ�h=���ݬ]4�GSy���ջ����j���1Z*Y��;��b��d�tԹ�Y��ɼ\�f"��-��A��>9�zǕZ�V$� r�騰z�V)���ySk\���L���p��Al���Ł[���U��e�N�P5'��m_5&��Rj}�V�%:l]��T�H�ݥ���ǲ����Ӟ�4�}G=^�J���m��7�k�����(�-Z������^�`T�3�L;���.��ٖ�0_���^�����A�If"Y��#U���J%7u�<��ܺ�n%�ѹ޷��:��ĩ�~>���4���L��.˪sZL/_����w�,G�]�Q�{���������|��+��p:���`n=�`Exp��=I2_�u>�d8m�:�����U��޿G�$�sE}%�rp´�li���v�o<�XR��C�0E����͛y[��m�=����|t�͚)HI9I�#t��ahn[[5�	�3�!��ْA�6K>���v���Z�:L�C����*&����G��븚1����-'"��}j�_��0a��A-�f�h�̐��a���p����y���r|��~h
\y���W0�'w��sߨ�yi����X_��Y�������]#��H6K�Kd���V�訽��i��pHe}������F\��ޜl��w���~%0'U�P�����{��LfU�0��K�2#ҍ-RoS��k1�.�i� �.E��.���я�/�O}�W].=����Z��� sB�����JZ����V
�L����$����~��kw�q�n ��E5A�U���JFNNS�=�:���W�/T��ޝ&�%h�B����✘����/R�H��;E��(�4��<kM�{>�ȡZ�ݞ����0#`�Kh��k�o�z�y����r�4WO��EB�S��/�1��Qg����k�`D���h_�m�%����6��aL9�����'��Ҧ��;�eM��h��L��+�K�5=ݮ��q�V^����<;=t�7�%t/bݺ�WFu� �G�%��Ұ:����L�LK��#xs6���)b���X�T�۝uC����@�<��Zʜ���	����0B�&{=^�Y�w�D�T6�	Wr��%ߥ�;�o)�ӟ�_)���^O`���#����<���'�>�ÄSS��#�:͒��7����d�&N���1�h��9uCGwu���j9�˹�ů��d��.a�m{e
pp����VV��7�,a���}m�;�c�0����[�<�eD�V����0���R�f���w{�7�S�F�����6IG�צ0�*�e�ce�GBî���ް�0K�r��{X��������!��}v�Yt���9S=RG���T��뼅oov���B�֦zvd��n�ͤ	�"��9h��\��__O���K[U�R�;,:�^��&k�4�ݢ�;Ksk0@���燗���lnrWQs�ۅon9 ��T���&���M@,&�U�.���=3�E��\IƷl)��gA����-s��`h��]M��^ɭ�Y�G)�[tjt�^z�Fqh�b�t�kM͌��ڷ.@
�kզ�K,k���d����b���u��ю��L8���_%�P� ��� ���7\��X0a��nY����F�o�IZ]�a���z�mH�r�nT3�sS�Q���P;�=�P�Y�:������m:�$k�x�<O���ɸ��/z|�y�I<��������y_�� ��멻�i�m�L�'h����.V��QKs�(zS';Xܡ���БM;�R�����t{/j�7�OG'9��",&�$��{�ywxe��/PG39�nL�-Iy�͙Qګ��,�.��v�e��Ly����˚�e6҂�ʹ��8�kHBfwBU�D�.ҝ�X�k�[��P�/=��L{�%�^̡��S���&y��оު�}TD��HiSh�8��ꬉ�wa6e�a4��o�Y���+t�j��pÄ\���̭kݳ�j�p����ت�8�����MA�h�cQ˟<��Y��.��oz�ȸ���Y�C{�t.��6�:c�ǴϷw*v-�t?vgMG<�j��=*���"�v��4A;�^��_�w>ғ�ٲ{8�V6�ݚW-����Y�{��d"A�ǉ����땳T+-��o�Y��N�W��)��������=n���f�V�b%.���7�F�X89��Qf^�s_C��у�ܩ2D7���h]�5�����`k1N�� ��K�/�X�B&+�Rk78V3��L̫PcT����`�K.��PغG�+\^��+Uq�bh�=��w1j��e���G�;r�t3�mj��ۜ���hF���@�D!
o�(�q��Cu!G���k7n�:�ul����\�--�FW���o��3qy��wWkߴ�5�"��80
��UЛI%�ӝ�Q޼\~Y�޷�%n�<�cIU�<��
��� ����}�G��Q>�3�٬����b����3]^�K�v��M���F�yKigM�(�g��);��ܷW'�&k�&a ��f�M;n'�MB�	樉����W<�&������	1�h}���7�(�Ga0"e�F�
Z��s^�5��~�Ȱx���{/����[�}�����8����~v���Ϙ��YR��e�m���>rl�	��"[��
s�о�m��oc�j�S �o����*e.����u�թ�:�/�wV�L�J��@U��Q���<tH��Ԏ�<Ɖ��@�so8⡙�'�d"L'2�!���!fc�B�窹�z䎪y��W4}�U�NFk��XSf8yA�{u�^½r�SoDM>�8�i0
����ޞ�M"����ӝ�nL��[Ph缢N�y]�c�Rm黾܄�tR&�mO��S��BIR��ɽkvĘ2Z���K2\8��=u4�:��"*�6�f�0������v5仺�jto|#r�W����[E�`��į\͋ێ��Y{~�u���<QJ7Un�댲�����Z���Q#ƅ�Y�[+(�s��%�7��*�%G��K�	�]��P�<�ڙ,��
ʰHA����e�e�s��܀�,aj���=�3�����q��Y���-K,*�x��K�Z��<𥕗Y�I�MYkD�=K���e�9�3�݀OB-0�N�`w�m^�^���g٠�Q��o&{54�������c�K=�Ƿ��^�ÕИ����󒆻�GƉ�YrMw@���Z�m��l6����y���<g���ƥ[�.����c��==~�{�|�qU�I�9.���N��7�=���U^Q����
��>@�w���+ol=�}u�܋`��p�	7��Y<�fW�v&{rA���c��WSGϖ�aX!`���H�ІM��j6�ήv2unL[�ֶP�\!�B�1���:cA�p�1/>x6�����\\��Py�ɍ�W1�>v�go��%1N_ܭ~�s9�@�5�5�Ha�������짚7��]�-������NC7�K�c��4�1���U��+����P��e��	��ͅj-{�{����K�����"�K�ݾ��CZ����GS#�+\��
ǧ�)��]���Џ�:F��:����f�Ip�gd�z��f�z>xCj�d���Ns,D0cn�^֤��U;,����q@I�
����핇"�B�^)�A�?2��5�H�:�R�w�����ݭ��
�D��ӿ,Z7�e�]х(X�8N�]�ގW���z��7Xn�~���Җ�$�2��D�����;�)����G��v��9�_��Z6K �n�x_�յ����q��+۽��eW�vD��\^Z�/��h_o]��s�@~�~qI�{~��_�����IPK��s2nzr����o2HL P��1L-$E�ɱ��KQ~�6�i)>Y�X��"��z��{��V�ҧg�`�d���^@[X�앗`�6��";};��@$��\E qy��b��LH�Gq�y�z����^ck����`��Vz��g�}��p�@C��GQ�#c���Sjn4� �����/��6F&:u�=��.^�3�$��T볝�ͩ�����V�G�}�9>�[-n�/�B�B8!��\-��\��]����EJ�/����W�L~�EtU�w� j�3���Z]ؚF��6�WX�>��6����j|W�wdԬ�tbN@�
G�Kf.��`�[����<2�t��VS#T=��H�{�ث��8��Q�E�p��a�i�%l��#=X)��yk��s(�xm�Bm���üu��V�ҝ	�gVM�y��?_�@3�r�e ��<b��n8Y������r�?�㫓�h�T�X�:�-JJ̓M��շ6��s��sĊHݔq̈́v# �m���'[W6ٕ����@�U��^ �v.Wj�@�[�-����Y�f2ͻ����]I�e&�]���bC;K��E���=��[\k����c���'b�L`<�$��w(`8��3�JPC-0X�Ah>l�ۮx�0�����^���{t�P�-��o�?���w+�2D�s�%;}ܔ;�{�S(!Y���q�w\���ҷ���L�牡��6�ޮRY�ҽ�v�]�L[cLZ�~�D4���2��+�+� ���.�r(G$��u���>}�_�o�s �TL�f�T<u�,�'F�q����dl��A��HH�a=���{�V�ÒN�g��������9)c>4��2U�Q�����+z���-tm$7Ʀ�]g��A�a��@M�<�e��*�]��r��,oA/W�sw�vB��%��,�Oe���݆�6"�U���{�Q�i3.��h���v5]�$n��

&�q�fǌ���G�J�=��G�>��X�is���9���D�%�ʬ��"�,x�}����|B�����*���m��!�R��d�v,�[����RF�Z)�ZT8���m
թx�z�1�bZ&O�Ձ�l״�/��S��П��!���)�O����sX~Ub��}��5q�{�"�
	��)���`7��3u\��Q]���xS̐vX���.�w�s� ��hʞ̿zm�� ��k�Kq���'� ��h߻u�
d+҅���=d�ђ� ��D��ʯ���a�z��E�8�*v�[Pi�0M���V9^Z�]fQ����.&�'XFd��١�����u����︈m-&�Is���V��;pwϼfl�����/�m����`Ԥ
�`�ؘ���mdY��Ӟ�fu����S���(4�DǤ]�o\���-�5ͺ�{(@2~�7*MxÁ3�Gu{��.�s�ǂF�oUw̨�Ӟ>��ݚ]ἀ\�P�m��G���6�d��9z� �껷�Y4��z���  C
��n���]ي���.�t�)��&t ��쩜����e�A�0��d%d��N�k)Uό��{4��9��N�������]��9o��	�oy_��,��!���/��qp�֪�\�wk�+b9���n9�7Ǆ.��H&��eI��ʋd���޾�W�z������W�;#i���7	��G��<�/�&#%G�onbS���B�B%�(����u��a�%x0�EO��r�y�0�,�;�^_,5�ׄD�y(�Y]���G��kw�'��R�z�׫̺�/Gr��*t�O��q����#qE�l�^*�7�f�.E���Bl
���(L^f_]�y����:�/4�_?����������q�6��v%�,��S!�բ�% �h�� �)���ܺEL[���@>W76o�%;=�g8����<�����y�ѻ�w�%:��J�^�Jr2�S�8���etS�%�$�7]�5���<-U�7r�ÒI���ۖ��Ƴ�@���Q�Y�n�Ӝ�+�>��g�R��XEr	���N�#�Zʬ�}��X����1��s��f0s���tz&IQ�e����{c���3�l�ޜ\o7�=��S��=�+;8�QG�T��;�_�Bx��1���=���;wA
�!�+����<�c�/�:==�\%*,.
��U�B�^�:J���n�)����%�q�F�����Ѳ~)�$������X��]w.U�zu*�U�
/s{��\�`e��Y�Gn�0dw˳��*��
Y�9��k�S�o�D]Z<q*�RL��֝���K)��G��*^i�S�����*�����Q�kjK�������r�KP(l���:����,�΍o"�r�X�Uj]�$!�\�s�RP�T���ܡ�93 r���Q��q]���,�P�7nr��8��q��g�%y��Ii��� &�rV��Rnz�5[�@����$�i�[s��8%_#�d��gw��;�Ȗ8���氏l�f�x���݄͏s�Oۙή�U���Ϫ�׸�}z4���C����rh���{��sc���đ<���W�,ڭ/}��>��k�k:��김b�\I�5ڃ{�uΞS��%!��(�[W=��a��sC^p(
�Ȝb��+��H$w�UB��e��z^��bЩK:����=�W�*s�E#��a��A�!M�ڙԚxyi_id *��ʊw;=��Z��C�Aۙ�8l�_̍(p��#,�5[M��ȂJ��cw����j�؁�\QR=���1J���]��.�c3�]���[���]wG��1֦��K�c�o�j�@�\���3��@�9���A�]�-V���l\�� 1��F�p5�$��(����g\u�u�GP���ց�ojt^r�Iq.`�$�n<X��Y}V/.d�2't����d��q��yp_�fb�p�x$c|�T�{�;��]����)�f,Իt�5@T�}Ck�q��?k�����ɽ
E���m=CW+�_p�?���k֦����e�e����au��ٳ8c%�<��"�r�4�8��:;��w�4�P!YNP�KP�=����'�Iз�A�A�{o Bמ��&�c�Q��Mܾ��̙Ļr��ĭ�ۜ{
�^�)S˔��ų@���4�N�ȍ�-r�Jl�����^�+�:�Uv.I�t&e�YI�Ԛ�$��i��W9G�zRθUs��/F]��\q�hp��Wmos�[���utW�۬��϶�؉�۾�x5Ӷ��ׂ�	�=�r�PQT��Ԃ���Vξ���˓?M�N�ݎ������ ����ƺXk��ёۛ��y���>�8�%ݘ�J����p/d��S�P��1Nd4v�m+��BoT=����K�+H��¡y�;�� �N�u�^4:(>?�
�����d\8�k�T)�ԧ�ߺwDF�=Rf_� �Uq�y���{ۉ^�j�8�<��o�R�O�ǀԉ	a��L�x�2/9&�몔�Tq�����=���ӫ��zo��k7�S�X��7-=��Q*��7�p[�^	�y�#I�{J���]WQ}���N0Bp�Ir1;��#2���95�J{3gqԉB=�,���B�z'O�l��!�R����ʆ��o�|�+��Y>��8'�I���e��5�7�pIKl�d��Q|���|�9�T�ι�pݵ�k�b���xӞ�꧘��$*�m-�,,����;D �k��v�n�Y4��[[�pwOR�v�ݛ��J�8�T4{��6�65�����>�8�h�A)J���>/Nd�Ȟ���{]#_8E�P�^:����,cs38���0�%�7��_q�/s��{�oi���ؿ�������7ا���hǶ� �Lڟ<�:jO �\��{k'��Ke�H��1�S���\�{y�v��Ä�^���Nd�OD���iu\�+������S�ˍn���J!��3Ees����f[~�E�S.�kc���fe`Q��ʜ�wjH�J4�0����d,4%�U�P�kX��>z[μ����e�V��A|��u���I���������7�$�����KfS�����6w:9�-��0��	+�%\������%I��=�	�1m(�Vqt�����vm�ƚ�c 1��H"�g]e��.��="�[Y�	d�0�`�lƛ.�ו� V�s1���&�JB��l��k�n�F��l6
��G\����@
��c������s:ȝ���,�'�r�.�f�\��Ħ�1�͡(��F�덈�a,����QE:���un�	�Q�*���Ƕ�U?����q�0<u:k�M���ͨb�VI�\���*��@��3��l�����bhe��#�e�yVa��gQ��9�L�l�}��F�gں��G+��+k�nz��Y�-xS�)���[f�����I(����"�����/�[�}F�)O���3SejX���p���A�o�����jn��9�80��)pI�G8	xXH����]L4Z�G�1��fxX�B!�ޜ1����b�����=�f�K{�Qվ�������駹����E e9]�(���)�L���_jDb||�UDN�YS6����F��||�ތ.��y�+��De��K!���(jP��K؝�t�ck�v����@�
.6��Uf7�[{ݾZ�0�{{�]��%�5�Mh���������Ǒo9�w5O� U�Pt/��}��~�w����6r���#�85�2�":O���(��a��T�^��~�cQ��(�2|���f`56ƕ��} �1A��|��J�/�3����� W���8i.�����m�ɒ �N;�N�Ҟ��7��M,�Ω�J,Ѐ�>|�}iF�^e��zO�_&^:�8	-��$v��oyuxV�F��X��Ĩ���89^dBvT]ku�Ձj��s�ˬ�y\���kP�-?lv�QpҎQ��Y)W��[:+"�w�$��ݥC�2�zЭ}��T�ã���"�E�J
q��V��:��{��B��r�i�iR�A�4r�)V�]*$ڎvDp�u�@n��Hi�na�	� QE�pX Cɬ�mp:4L!��Ο�{<6iU=wC,yk�r���,��:� ��߲(y�w��}�L�����)��X�S�
�J��&j��|�@�;�v��x���o���'m<_R}p� �\����7�+��J�9���1�tr�Knd���ϟ�Ϊ�;��7�	Y��Ɯ�>�����2�B���yV�]]��|�̆{}�S��`<�Z�LH�YS4�OSLg�&�c&�)<
g�ٲ�7��^�h@q0a��IG����2<�'/���p)�=G$�.��vM�� �:|J�ΝUhT#�j;���f�p@�|| �>0���D��dVA\
0X�[�]wn�`�h�^���wr����;�߶��G-�57 a���ucB��Q���h��ޝ�Y-+�~5|/г�es�Ԝ;�����<ӛ��s}��.�˸� 8k�C%��2���Ma����Y�GΎ@��C��>�|�D��(@���p�F�ۮg��M!�n�h&㌠�d��;��~�;{y�zWK�cT/t_����M�����b���Ϋ��~�3���A��v�<���>󻵂��KhhX�<N���Oa�&k�N�Iz�u$����4���NWc���}Ɖ_���x�wq����9��;�;�&���m$^v\�UF�0�9���{��RN�O��T��/I��";�f�U�6����8��"eoLFve�7lw���]�O��É��3���a��
h������|�1;�)�-����W�6�>z���L�{�*��� ��� ާT�"3���M��Cs�}O}�q���}�o��{��烗����M��ٯ%�}�� �4�,��*�^��y̏l*����4��)V!U�3�M���RKQ�Q�SY�8�os��d<j���� *�K����4�^K���[h���\���V9���`�i8�����0�.;u�;����躟��~�	�<�Ͼ�Φp��}�^ȴ��J+�~ �����DW��ӛ�{}æF�3uu}^���z��q�Oo#�Ȃ�m��dG `�FY�������Q�p�qF���l��x�&ی�Ik�ڵvٚK����;sv뵈����0�މ�����?M��m�6o#�qwY��8�] ���C:-jt�����og�ߦ�Z�����P9J�� '�Q�Y8J�Xe;���F�7
�|��Q ����i;�����ﬆ�'U�3�BG����
�Fq^��[�Ϯ�h���൐�a��p�T`1�vW�;)gwd�'(@ׇǥX��i���rB#��Cq5q�r���}kd}�����hт���u �լ�#2��+8�Y��%���.ǳ6�c�(���Ր�w"eN��{��F����S��.�Rb��e�UEg6LRЂ7G����?>�\9��s�İ������EI�}69�p�!D8ˑ���.�3Tŝ�w}UN��qj�}S3��z��}y�j:����$�T]v���O2(j�^��e;%P�{;���_���F��#�t>J��Ao��I>pEb�י.��W���zWz8���e��J2x��F��=s�f�4k��i!n
Jʹ��{�L���2:���͎��`�����5]��ի�Eׄg�1��֧=��AI�	|J��^���}S�s`I+��[;�=[��j� ��6CDȐ/�hqE�	vŅ�])�Z� e���ꫮ��U�O������+���O��U��d�5%AG=��;-��B�k�tsgs�z{"mu��,$G2�&
y�}�r}��T����D��=�rP ��\z���ʷB����V��L��eﳳ�u��ȍo��89�����5�'��7y�0���V���'����,|���ꫦ�sG���Dq����oo;o쑓f��Kɗ���j�uf�Hid���z���~��^�^���H:8[�������F�R����D����软J��W�7��Z�A!��2Z�OxF����v��{p��CW������o��R�{A�sV�bc)���Kd�}�e	+�:Mu`��L��֝`:E���ef�޴��9ƱLCI
�3E���s�ۄf�&�.4n$IEM!�Ԏr�2�k;s��0���!�ݮb�0VӍ�μ���,3e���Ӯ�=4k ��[4!�,UJ�1ٶ�n&-�m40�B�YE�!�n�?kkp7-�]nƨe�����4����f��\�S��t{�e�N8�չ��8��A��zh���#�U7c�g���Ʈ n�r��ݦ�C㧌�N��~�R��G'����u8F��.�m\�Oi���kШd�:[��β�ʮǼB	��Ap�)��l!j�3ut����>R9�\��ƧL�5�}{nL2��vV��9�I|��3G�q�'oy���`ƍMO �	��k�9���X�o�4&��v�X^�@���L��/����#[�̥{���N!��Ľ]��v���%�������ٶ�ɻf�D������|l�,�P�w�ͳAt�� s����z�v��J5�z�-�m�{�
�Lz���$Ox��\��w.�7c<�Cn ���u	+(KL�λ<��&mѴ�`�.�R;}� ע�]!� B��2)�G,>9��8߼.�h�5��n�}}6t�m;���z�.��!ڤN���+}�^��ABg�em
Hs�y��%��9�R������񴵼���,T�ra��?O|��������l����k�¶���$ķ����c�[���s9��o��$�H��$x%�r�8,�B�7Y�4A��i��C���Y��G�����\鑒=�i|}{x�Q;{�-�N�V?gY~:�ٳ{Y�ʉ���Bâ��52*�'���8���m5�oS�83�v�6��Y&�߽Q�+Qɰ�O�釻9�]D�;1Xb�����=[>��%Z�N϶u��D������.gG�&��d��EDF����J�uj�Wtf]a*��4�֥֫z�Pfa����q����u5�M�������̬�D��V�b{����A'����%
*d��T�H.�y˩�&�� .�9�:(�p>g�����}��c%5��9��`3Z;c�ta.v,�ke��E�,��I�P`�*�����"�|��+�Ţ��V�����S�Ȭ(c?_GٰT�_d_4��Jw��h'ӵy�I_o���"p��b=��{9��u�K��֣�����	����_�V"T���̲sokh�d^7<�\��ɉtt��� L�U޳P�疼�B-Z"hЇ˯�����"S	ۃ戠�fSɤeN��>]fk�C�s��?z��V]�M/I��Q���B_^]4���bS(NN/o��w�ړ��5��(��c��I�_X��a�6�[9�l��e;��#A��a��꬟i魥�q��=V�}*p�V�����sh�,=���8�XҤ�:�{�:�g�����"�A���U(I�uq!��ϑ0]&J�Z�ݾ�E���"Vy�O�gnݸ��u+��Ԑ�dOo��x�x�Co�q绎4��Sob��2gwmx�r��H Tk��Q�����)��EVϾO+���ł��̼�>�tfSu��4�C�c�H�^�T�'�
��s�9bUţlmXk�]�D6�Ϟ�h�ɋ5^��{�*��^���^����r�"�厩߲'�݀tv��e=�[�2ϻ�S���_��	3�_(<�Wl�CV�ѓ:���Jv��W{ƻv���S��3��*j���Q�r;z	�5��Y���_��wyt4a8A�H2���D��4��~ϧ>9����ǌ�����u�Y���ku�K����6
,�.�0x�q8JM�C:�=����X�Z�:*�{�z
a��"b�W��y%��kқ۽ڸ��]�Õ�d�Bo�ަ=�ݵs*�zMs�4
dL��u��"�b�+'{�r-f{\�Ӯ������2�ĩ�ں�t��wX�BA�Ppڤ�!�^yS\fӗ�t͇�3'MdĴ
������C�s�>�Yj�}����4rA�W^�1���%{�[:�ϲ�k_v���T<���6�Y�9��Ck���b���:�"�7����o����{��M��O���؎MO�:���vo���K�K��uz�B�dOeҺ����ɥ
�%=��穕�]X@����1�����,�cT�	U\JGJ������Ȱ�2���c���aE �\S�s֤�!.N^��\vBp&c*D�_2�0'��s6žf{�z��*vO���{}9�s�u�6���뤨^�i�NVZ��E[�Ů9����/1d4{)o;�i�5}���>B(��g�Yؙw�}���Q�% ��R�9*�ٌ�9��?YHF���,�}gI�>y��7�+P�r Q�*$���j�J�J,A�'��_e7u�P���Rh6�ǁ��7x�惜�l��_5��B��&4�5�\+�iK�C79�R���m�V���iu;e��ލ�������+%m�wkX��)XwV� 3ü��$E�G?<�s�Oְ��S�JuNWYMʲ#|�d�JM��UU�1��η�d�V���ڦMܖ����3T'�7x)�Ͱ�,��mܜ6�Z^O��]�t�Zc�G|*�������k|��7�a��\�s*0{��ff��|���f��h����?jt�@@��}&�o��YC��wW�	V( ę��s:�sO�8Ǉ:�향FD�d3]/����)O/:=5>/�<��I�R������*�]�������+oَ�����W=5j�Ͻ�9�aAi�X��72d����o��_�٩��Ϲ��b	��?eW|�pF� �� ��l�|nŷ�یz��4�!3
LGq���G�]�߭�x�M@b2lnN��jf��?�t�86'��?A��ٮ5�)�a�	;�y�f:���wWn��]�����Z%��x4�͗ޗX<�4��F7S�Y�|�+'����� i`�cB�E��kE	r��Ɖ��2�H$b�&�:��w�ss�F���������p�
2��n�o��C_m����#�1�j���J �v����Xy�=[9>0��:"Y�J����q�����łsf���2 l:(�ہo1zr�ZC��{��Lo�,R��D��WU5UvT�L���[,ͣ����Ȱx��մ��ov�Rش�T���n��t�侕�rͱ��0Nt�����g�/��=X[�����4�\?W���{o��������'�����q�1a�_"�2�8���켃���u�ۊ�n�r�V�=ǝ�����cZǳ�q���F+�Ms��a]@��MKu13����+��2�����u���Ez� 2v�0iX����>6���B�$�Mm��#u \�s{,m�h@��t�YB������퇒m��O�����@��L�B ��KK���=	|/c����.
�;HF��P��v�.0R��,����f��R�p�i�2,�B�p�x�.z�<�c�ڭ�V��^*���G�K=+�t?$ڗ)
�J�J�T�˲��<��QЖ��=��B���t��_��ĉ��_v��ף����ڛY��)1���A8G�{8^b��6��r$��]��G=�}͗d��zO	-浽���d3���{q>�"���cTo�p��a墓�<�U��ht���*=(+y{R7�{�\������p�=[Ԩ��W��&��[�.Zz*�7*��P����C%0�M4 �iwg��i9Պ��=�H�V��G�O����<��۲�e��s���o*�b�q��oFa�\Ҩ[�C��X7�ryX�z�`���w��*'�z4G2Xa�D�;����Sn�\ת.�ߥ����z�U��>��T�I|���Uٴ;��?�aҼ�N)�7�HWP���j��<K��wU��Z���{���
F<����nGh���E�	}^���,�c����|�:�C-|m�ƣ��6vHW�=��$,�{t�����*�-%Ȓ�t�y��yG�9��%S�HE�s�f�}z7�Ȅ	�`�ٔb����&Ϧf�o��hw����ߓ��	R4�R���Y�ɳ��/�&�^�[�އ.�j]���_:M�������{[:��6���n��u��]g=G;�k�@jK��Ɉtv�O����C}���X$:���1���h�yô�ZI���˿u9�<֣1��F�Ä�N�o�)M�6��7��7��QU�יr~͗�k2��=�v�ՔT����R��t��EN�݁Z:�g�9�jY�;9+:-����k5�XD�%:j���[;�n��#�;��T�]U�t=�V�Kn��c?+ޘ�1xb(�<Ίasr���MbM6�<8�>���(k?+�*��O/�&����4S�x�u�ǹ����=Ө������,���C��9�f���uOH��j�L�i��$��/����B��Lǻ�T[7Q�_��Z=.���,�5U�2k��w���6�-&7�~��O�5@�v��!�}��h�ͧ�9l*Ķ�OTьUN��WB��a�f�f�
Nt�j��q�C �7,�$n�Z.w�/�8V' 7˺A�
Z0͡9G[��Lb����v�"��\���\��m�<lǃ�]vY�z�л�4����:�[�qʻc�v9y��3��F��\�6;o5�TR���؄�"' �Yhwu�c�y��Y���t!�իuٝ�M��dGg=瓳vY���m�p��ڎ0��<�4A7�҆U�V�rAY�}���>��F⸓��P�6fП��I��{�6�۸���k���r�Z̬�?Y��Ұh˛G����i³�
暝�۸j�Ҕ�y�����%���%Z�Z[SRUU@UNI��ff�%]�,ʴHM����/[����7/\�v�ԎL�=oY��]�.n�c\�r\;��Ò��ݧ��/d���1�tl�i�c�5]x+�-0���x�l�`�[1��8K�8f��B+�^��ٳR�f�4p%fq���n����Wc:�Vch���������c��Q���gp�Pl��u�k�����s��a˶�@u(oR�r	��d��8^�cTZ�Y,�4yh��LEH$Mq u����[��������������&��θ�l��F��#rM�\�q��¨�Mq��9�;�ݢcl�P���3��YN'�U(����N-q��,n�:f'%�[�Bi����[R-��-h")� ��,Z�"���μb�΋45��V�v��F�#n%f�u��Ú�ڮ0�d3�)�dQ���
��v���%�l�9�%��L����(p��H[@�WYx%Pێ�n���͖D�,%�}�)\�x6�v�6�f�۶�3�hٸ�+e�	��.�`Ң���6]�HnDLq��Z�d��%�T+�\�S���̦3�
=E6��Nz^7�U49�қ����!��{=���:1��\.љ:�tvӣH[
x�mgx��8�'3��](٣ Me���j�`a����\$��P�f���:.�Od }��^�U�bkh5���%��Y�۶ݖ�\�:�GD�$l�޷�[f���C�^b+��r5LJ��mX�Ҍ����j:�]x��� ��`��x���Ա턏
��M .ѯnՒc��p=6�ۣ��`*�	���4�ҋJ�Y@�eT�]0�k)Bk�2n��:��j��c���m�>���%��ݞj�0��f�X�7V�e!1V���'z��g�g�N)(/U	���/��s��9��,���6����W$����ۧ�+uu��F�����	2JpZ��d?�V�gn}}�~ ?j��~���u�P����' �&s�O�B�#��բ{�y�VX���g=��.'�$}6�m��(��.�,�npe	:�S�ڰ�+]`�P�.�gU�{](ٻ<@������;�a�|��:����	�E&���z���6.v�e:��R*:8��n׆M�ٷ��.l����K.��ws�Ɩ䗎��VGW}�'u�Yq�gg�h"?�糎t�ӏ�޽LB0Ex�\Ok��10�.$*�f��u��^�᧛0���� @91[~��n��֯(�S�J�{���a|b�=SJT����hA�J�;YS{�*u/+��/�˞�{�*.��~�z�|��:�����u��Q�Ն����wAmG�]�X��!�G������Ys�=ڿG��L�����w,���KG����ʜ��aw�_$�]r�w�ne�w���Jh�	�#ӽfW�:,!�79��-�V��[���Jb���ק�[=�}{
O��������ٗąt���pA�Ǝ�S�lT����|/��<f����U�[��-&�lr���c��R�O{n!U�0�Md���D��點d�A� Ú��`�����^5J.{q",�5�v��Wmq��(I���}�ƨ��Y��W9�X-���V�S�7�sWu���m�9�L�u�P7�V����o>Ҳ�:4s,~Z�R������p�եSm��[ў�A�c�!0�Z%�C9Ԝ*�S�n�x��^Y��{A=��4\N�u�r!e�����wx6�v���PcP�z����u��cDHU�
�;�ޣf�NG����$�L��Wb�$^��;�����zNߎ���ʞ���T"�A@q�F
��<��U;�l��W���"�{m���p��Vf�1�,��KM\�P��!�\�N�u[r2�� �����y�Ǉ{3ixϸ)���s�uQ�³���ـ�c�4A�BM��̊�/���;hU��Y䑴���ܗ�.�ͪ"'�V�$#�y����^U��ڏs�I���l�{�����q������(뺮�T��q<N�)�(����.ږ�1�4�E9͜w8��(p6Ha~�}t �\��)e$� 7:��ADp!E)~�^�߆q��}�p�}]��w��bK@��9�WFGt�7�^��w���o{oh|{�/{�:>�5�OMu�.t�x�"��CC�	wm����c���z8�ut:�Z��M>t`��a�~�{}�}��l�b�ј��
���ٮ�~�*˲aʼ�\� ��%�܂L��j�bw��/u�޻ӆ}И	AA���ymL#�+��7V�/6+���W^�y�W��O}���*�Z����|� ������%]Y=�ACnE�R����!�$?�6�(��N��&���D���8:L���^��d稒��N��<��Q��޹&H��|],���c�9[�Nʺk(��h����s��쮭���Z��r
�5>�T��k,E�[ф�� �:~�4�՞J㨱qd줾�Wz���Η�2�O�x]�Ѵ_^-=�\Θ�����/۹9�0/zD��Tii�^߃;"�(;�y�M��}7%{��z	��z+�������R |�]0}˨���%����u��e�^�����S$t�qpqގM(a��p�}wEՙ��;2��!�M�����,#���*g��>髽sc�'���p����
�f��o�����J��΂�c��mvq��vbL�ѷZ�� ���Ο(y�{���VQUd���x0`�}K�||{kj-	�3���;��nP��e��>%rQ�0=��nvA.z���\80bݕ�o ��P����`��߿v+��>>��#�0$����֪G'��9;��\�7ktĈ���n7XnQ�����%�`�U[��l  C,��'��hEGA{�m)�|Nye�4�e]Mx|�Q�Y�QP��˹M��q}1��oP���7��kE���K6o�Y8}&�z���������lC0�!\^��o�a
���[<�S�����T�M%fV�f���pr3˘@(�3ګo$��>b@��#��!9e�Ŧr;�bs�"�,�yЮ��t�B�$�d!+Q>�4ȯ�V��'_�g��.�W�u��:K�T{�GȜ��uq�{��X����q�����M;����N%��u*�k*m˧8�]MB��Tou"��-�G_x�^ǩ�{�c�UƛM��Y�%	�	2��"S��\�� ����4f
X&�'E�1�ZeN�:'��m���G1�Aqk��l�<�!t�Rj��f�
�Gn���ak�ۅ�7��]�#��,v�qn��#��e�����èA���[�͠�������D�68C�uf��`��k��D����̱f[S&��eDlP�p��C0ˇ�~�w��=�+�~���8�F�6Sw]"��?Si�$���w���$�ɨH&�4�r!���ob�X��W7�G�k�{�ٓ�ӑ�@�������W�cyy�M�U��Fa�윯{�fn9Fy묚��^�-o����K1��/�s���/����,��INv�����YE^^fu{���{���)x���f6PQ'(��ۣ(��|4pc\�Ѵjj�yѵ��V��vp��ϋ~s6j�@���@��)�fi��p�/�/���$����ò� (�ń���n���o���6�6h���!��/����=A�"=k���fo�q��;�����$�{۬,�1Z��Hy�B��;/�F��]��/(����wa �%B�~�`�"q%�yf7��[�-�xwÄ1�`�^15n��;��������?z|i��գ�Cu���)�랎�{���z[��탷�+2�o��%&�8NЛ|��1�ޘ�i�nWu�:��D���V�n� ׃�]��<]olfL�z+��Qӫ(͡��7+��.3��Ԛ�I�97�����o�C�|Y��^S��4p�wJ���=bN�?��Cy�<��L��Ϥ��@"E�62�&Պ��2�-�"�<V�}_zU�uʮ�}]Zr:�[�mdƧlt��3�D�Y�:���$�U�A86R�n��K��SL{>�>��,�e=��Ӗ�^�������)������= ��i���
OY�keG�W�W,,�ԌKu�pj����p�8-6L,���]�Umr�28#6��k�6u�r�c�6i��/3�����{?RZY
����|�R�3�Zi��s���u��:������ǲk®�柺=�r8�RBL	��;Y�맕�r����Uq�]�=T�X��#ޯP��ҳ9������=�7�oxґ/�%[��+�������]��u��lT#�WqL&�e6�`�楅��xhk��[��V��3v��ŠP�FA�;��z����"�![
�\=�r�u�"y�^|+��Y��χ�^��R�3���}wl��c|N�M�Y�����x�;�X��|�SH��iv=\������&����@�1������<��Hھ��E����Y�H��	4P2єϞY<�y�
q��'#@%���{ �ɦ_C��W��������I�.Q�|S�9�#p�#ޱ~>ר�LYB;�u_���x����f��N�VGq����m8I�ʮ��)K��o\��,^g1���N���)q�=~}��`�F�A�Kp�����\N��W���=i���(��a(M���ӳU�	.6�h�0\����%;�����d�J���W��M*�]�6B��]���:��傖�ذ�z�2���痥�u���X^�j�yѻ�^	�u�f8ǆ��n�	��g�Hގ��*I�b
LX�<��v���03+.I� �y���'F߸֌�n����w3�F���C�͒�@9݊�Y��ce��Og+�2�ܿnL���]Qw꽡=�j43!"�ęʠ}�n:a@O:S#�?]k#ގ����4�]�{V��ګ�0� � ����;y�C/���L����3$��D��Iq�Q�XjK�v��Я{�5�-؁A\8l4{�S�ҫ+�(�y�[
ք�?/O���k>�b;0�Ӌ���°�sֵ�Ɖ����#�+����%Վ�A�s!p=�3��{a8I��Q�����J��;��@�O�M�zWD��F�ڶ �r�R�J��}3�xWO{خ������#�\��R�N�}BP�Ee+n��}�<��MX���Z�Ib~M���L���~�Dl������� �[u`�Y��h��a2��L��#t,�WۣV��4V�*K4���~|w����U��<ŗ&!�c�)�.�;���s�����n�x��p}O����8~W ��ɟc���Y$�EH�	z�Ǵ0��]���h�~���5���+��zc�,��}��2���cs���o~��i�d(7�h�ɦ��S뷇� @�47.���ca��(,ڕ�Y��rU6���j�_����(��j��<��X�P[�Ծ�֛��f�ӍR�D��f^S��K�^��C��
�ӫ�ݾV���S��-�Rk�����_w���c����-n�����a�H�'x�<����Uv����Ę���Pu��۬��E'F))��}"��%�#���*����A7����:)�9K�ҁ�#O���8��܆��Ӟ3֭ewMz�}Nq�H*)G��*j{t�sM����W��mh�Z�-��{i�x���=��y+IU�wJ�Fr:��chӻ�B�7D��E�Kz�y��ez���gB�^�l޽�r��#O�Mh�����[F5�ڷW��mzi�<G�����>jT�5]�&���@��9lbس��S%�ۇ��BH�!2��D�R��?ww�����i�p����s9��dy<�P��r�t�|��o	�����^)uk���{UW,����PZ�U6b��gp�c'�wq⏏>%|Lf��}2~�]�H�<0`qu�X�3/�8��Q	�f�r��IF'�Wzk�U�Ű�Ό��w�[���_�A���@����ͼ�������P_	3���RJߔH�.��c>�c��\��ٹ�o�׼�n'�j�J���ǹB6��~gv˘S�W1g���w:8�I�h��kM����uΦo��ͯ��i��fd��y���M�т����]�`��jI�9y�{���w�V��x2"��W��<�63��X�h���w[⤆�C�t�s�)����\����Uj��k�4�@S^�l�!ZWd�L�L�2�Lݫe.��.2ȥ��EͰE��C�X�6&�*��fARmf�҈�.»�����n����u�j.#>1�3�rz��͚�s�̅a�u�Yqt�:�(n�yc(p���u���ͮY���C5����l���#f��B��X��"�L���@�WE�lx�l @I�q�	�K �s����?4G��(����+�R	\���M�Ϛj�>H�!�:��NC���UM�+����&���Y��<>�b,w^d;�d���'�[Αٽ�O�f�w:�[u�g�1P�gw��l�^ލ�m 3���WE�0�x�ל��2��T=k����Gy��(�&/���ۈR�
�<� �E�� 2$-�m�X1�E�ZY������y�LHpQ��Sf�%��7z涌�خ����M_�<�����73٢���qA���)���>-���Yڝ��	����q���g��9I�[�m����מ�_ko=�_)6b���7��5(�+�|=������Wo��p!�	N
ɲoVYVc�o�G����
Ko�]��dӡO��O��'�Ní�N%']�f41�-��][��'>��U k�����=v^�ݓG0��`���9lHӱ�V�_�N_��pMe;F�f�]v���Gy�a)�s��o�ƞ�;s#�חS�Iw��sӯp��Q��Os/r5��8!������>;Mw���}�f�c�i�R��gM\���f$��kc��u'��`d��'�ߗ��>6s��u6�nc��y����ڡ�LJnB3K�ߓѽ:6'K�%7wR-A�v��g7��lmp����������"�5�U	OE=5Ѱ�j�+���H� ��b�Fw�l�Fh��uS��ƭ�B��ׅ�����zl��L/HJ��d0�ո�i�N�d�Bp��&-�7[����U1�J�||f��n��}������oغ���i�K�d���xI�m{��Q�#��e^�Vs�;�)G��[�ν1޼���"~p؂�E�6w�&��OguՅ8���W��j�� ���o���ד���t{�{�մhu�\�vF"�2�p�B�U�ϴ���V���P��.M��t����ML�����\���{���Vʀ��:����g8#����v�Z�U�z����\�e,{�r�;�*E����r=�O���&gخEN�r���nv�yL<	z9�V����A��ﳳ;(�W�+����c7�x�gn
�����'/zs��one��[]N��\;��C3�(���Q��U۽�[N�YfMt�X��[��F�Yu��Q|�\�P~{�(��B��dC��gy�������̿wC(Z$q����ri��+Cw�k�������\���p� �n�>_]�-�b;�]1�8�11�����o{�y����R!����D#�`;���m��+rj{v�I bE$��-��Q����s��|�'�͞@�#�w���B�������믻�E��S�5�^����t��R�}6���e�BK�쫎oMі�Jͷ��8���Ь�{����{��`�c��k�^'J�d�����j��g��_'�E���;�R #��z�o>�9-	��exL�c;<7VNQ�f�yy|��D�C��9+唁F�3��]2G��ɫ!�+���շ�*o`OW|�,�O�� �9��=9��;O��8ր���c�JSc	u5_w��f�֫�U`�Y%����V�����א�t�uy��g%���%�$�9(0������rdo��Ծߔ�+g��2u��7��]���Mmb5�>�Q{Y���X|�h�SW(M���G��he��gdf�h��XTl"���?�C+Hh� _{�̓^s��\���R��v�(�Tz��=���.�|?U��HW��#"'�*�L��wǦM\����ȿP�����Wv����*ȹ�y��%8e��lS����"&���W����>�c-s3����)\�&�7O�&x��U��0齝��qMm�
.	��$�	ś�Umr�44ڬ/���b1!�Fi"ue�ef����7��L��;�K��GZ�^Mq���t� M�TM�4���N�a�j}�x�AYE�c�����ta�-��M�������}� �������8�>��){�pҾR _"�5�S�5�˓N%�K)���~Y����ŝ=�����l?�w����aQ�]<Wh"ͧ.��y%wMZ�u˓Ga����yo0r�2���(�;1:Hɦ���T�+kPw9���8��\ȝ/�tb�cq��]���&e�Be�^�tJp�F��9�șe	���)�Dll��%��g+:T��&S�)`;u��J�Rw��9��pv��7���.w^�f�OY?�&������+OF�|R�R�-�¹ӝ����wJ2�8��W�O��n5��@srQ�����y�IjÆ ۖz����JuW��-�]'p��"�u�c��EE�� ��h�;\$�Ck)���g�R�i۪�f&޽�� n�Y�i�ϨQZ�_��,y�]YZqtC{�c�����}���AN���`t.��xvV�gd��ܑ�r�]1�s2���^N^�����-�Z��X1i�=j�Zj����Ф��؝f�Ӳ�E}�_��H�poN[G@ol��I�R�T+�Q�U'p��<�K%��^��|�A����Xq<�S����Iŗ��Ր
�{�/.Mt빩�˒�L�]n�,!Y���j8��s���紐ג�clU����p;ab��tI��I5��N��Zʐv���<�g\�]�͐'�E�j�$��,Z�}C{FSˠ⢝�E�ν�wv�e���El�і\Y�f	�q�;7`��/�0�wmBkEw��5jo;r��4��^sʰ��#fq���i[Yj���es�g���"�,�e�g1"2�G���)== �{ض_�s��+�f�("�-�w��!���� ~�/���ϷLt�O�-N����
�Os�+%{àr��m�AMܓϕ�v~J���DX�^�wP_t����՚�?\��̂cc�QH�*��KL�	杛q�ݳ~8S��ƭ�����Q�~��$T$�I"���1Ÿ5�.dk���|h�%3�������\p�#�F<���.��vｕP�q��:^F���ɥ&5{��;D��́:{ËH����pR�p#A�v��ŵ�6�'�;�͘�#/�,V_<��г9�6b���j�I��q,V3Z�ȳ:�\Ane~���E����߮��ଟu��L�Պ"��	]����S��:��u?V��É�>�pL_OFR��Y�Tr���R��﹜ ���~�G�����b���Eh���<Q�8"�������i�!�9�7����T��w��ܮ�{޽U�w-���P��@�*�N���0�|~oe�P����	ʷ�cq���j������=>�sȣ!�Otޞ_aʹ�:������5�l߷d�m�5�7Q6�[�U=�Â	�@-�O���ц��O}�E��	�s��G]W`b���=u-=��g�,���$rԨ����-JV�]e���wL�E��F_CgP���Ջus��|�䚀����]]2��9Iyh\j*��1Ik��	��q��l����pm���>5�ꝑ�%l�r褆2M42@�����š����B/n��g�!۶s���<lD� `92���Q�����lw-�1vh*;^^C
�b�:��Į�����qs�F69�Eh�8�6KcY���RbjL��;������i�b���l��N�E���^�8(�vu�+-]�^ٞϭr�^V0�Ne�����<���쑝��.���L'��)���Y�G��m�\��@����Tу������U���>9�s�!�X�8V��B6���37^��q}�u��ɮ̎�^ע(�
*�3΍{������r�'x�^�����ԫ��U�g�=`���J�c�	L7�P�p�Vf�����ǐ�ݸ��Z[q�뵋�o^>Ϟ����3s2��M�Ga94^o�G�΍�{���ݗ����PMww�س��C��7K/s�f�o����(�����S���%�&�ܹ=yţ^,���}^ٲ�8��%`�=G�=�Le���Ox�y㯍o��J>���v��^|m�G���vM�#Dq� �MC 'w#�1��=���GC=L��5_>7p�=wk�1V�NXh�7z��Eq���徐��^��i=b�v�z������>�<��1���Iؑ���������-��gB��~���|=+۶O>q����������M�XhZ�ـ&4����`�u[�2
˦C.���:c�:���)�g��&�p�B���#�55�}�z���r����3tS�$��	=�]V�{�������Q7]�]�J��{��o'��G�O%��=E{RٹW��f�Z΃�47n�6&�&� j����a���������Æ��1����tK�b���i�{ �$�c�����A��R�ia��!>�l3���1����6w��/}��[b��_��cvͱb<�ӎ�"8��ԛ�/<��6�f�jH��B&d#9��Z}�����y$VH��4���렴S��V��x�qT�&���GVz� 'v~��Wt�T�ci�#��kO=��4��7�r�#�3z{9�eԗ �9�(Ǚ��v��ؘ��{;�{1����t�"���u��yӋ|#-��Q#�=|��bṵM���<}N��މ$a�>����~_`���Ȃ�R-�8���.uŋ�{w����h�u���ʏ!0hZ���-�f`�n��Ǡ��i�$��w9A6�cپ>Vv-Ë�}�s̹�Z|��A�ҽP���4'��B�[����^1{�lPƵ�D��g�K�|;R�YE�e���-�͑�='Ǫ,du����=��N�-2�߳��W�u=/Ĺ��]��3�p��8�����}�0S����k��z��f������ٌ�8mg��qk���w�^Lh��{�"s�C�L.�+$�&E퓑�u�M�Y5��]H��W0C�ݿץvڊ�D4����S���@�FH�}6 FX޴&=z�q�d������͢y^Yu��������l�A��&��n>�X���5�i��]d5Np��{:��;!x�O��;��{Ւ�/��U���EsX8"�$#i��R�����7��/O��4�:+ܽ��\VR�KK�n�d�zu�>��ؤwa/|�@~ژ��&υY�9{'z�D��g�1�!R�������sUz�sn���t��+_�m=#�O�c������׍�Yg)ڶ��4�ze����g���y����wm���k����sd\��V�sj�{u!节�P$�$�e���y੢�v�.�x��8�Y���<|JY��R)f:�~wvP�FaD�������}�}I'e�6�>��%C!��E�W��ЛK��2���=��γ}��������Τ��=��2�q>�9�c"d�M�k9�U��zj�*�K0Kb���C��v)߼���r�5T�U�=ݕ�4�}>|Anl8E�
j�f��$U<ʥVjɉf};���m�~u��/����qXtju�Y��lf�W8����TBh��@*!0 PBi'�����\���I?�����Gj��7�[f��{QZ <UŪ���·="t��[���:u�L"�)�Ꞃ�	x�j���j����r�]C�kaG-��ק��=OtVe��f��/yZ+A�V-s���WT�����ʚ�'x�)l0$�F̋�"N&�eU{����t�4�AM%�&���U�Z:_]�:���_v,&�1.j���ok���'X!�x��F���o���.��<=�����-J�\꽂�� �ʞ�2g�}?y�b5-�Ȯ+�8�9N_��cB��(���;���A�sۨΈ��t�n�ң��ڢ�`�l�>�ңNT{}ӑ����g{jԓ�V�D��]L�+����)�;u��{�*�GM�LQ��R~̙�g����z���70|tSV^�6�DJ.{�a� ����(�:�ks �Ŏ���N�>��u�j߼1�@=�A��g�7�{G�T�����{s93�qy<ܓ��wy�ƨ)�6Hp��)Ɋ#5�0<d7����v��!,���{���?'�z��/��y1ٌuOD�>��<�n�ы�uv6�2�o"��	����1�<4�i��<d�*�j��K˦��ɬY1�|绲g�S�K�-{���w��x���W��;2Y�����kR|sŗm0'�߻���>�~�S�cK&�g�-g{Q��4�b΍�ՅP4��7���.R���lqt ����&r��k,mo=�X����S��z�9�A�o�8q%��?A��(xH��s�NU8!9�{r����D�q�≤Nze;�w�RZ�y��
�D:/��k���>��[��ƴN�],�L�������{5�)�;)R��3]�9�����כ:� t\g�e"�a5�9�V�x�����p1+��z��+�4p���6��+t�*{!�W:z�v֛�U�s[{�J�u�ġ�A�M-���,��q�=�,�od6�gW�ΫuFׇrD�v�T�k���J¦skJ��x�l�n�`[�X`��b�!�tL�. \�R��[��fS������S����S���k 飌]6������
0������)�Ż�#0�	T��s���2�Pa����0��J����y��9���2T�T
�np�̦�4�%�7���6���O��m���ͯ}sĹo$�Ϻq꾬�eR����J���J6�w�o�_����͋�lce[g�2)��^v�}j��k�xwC)�i8'
����r��ܼ�e��Ջ��)�1���AE�<F� �. �d��%]��>s�q�CW+����I8d�W=
.������ΰ'�� :+!�}W�w\zYUf��X�ݳ��S�|�G�,�j{������}��i@(�!A.�_�x!^͙�=���nqJ��.�R|�Ь|v�����ü��'�C&g�0s��$�p�&6��S+)f�|�MQ���t�A�A4�Ɛ �%;������?�i�}��!��q3�Q���k7tf�+��-3�|�޷��>�[�CNQJ�Ѡ|[ٰ_�'4g��`�q�$h5����u��Roݒ ��~-�8���3XP�s��,?m�^9P�t1b���K���f�����L�gڎuz9�%���t�������"X��t�f��%�z�M�M��.�p`��k�>�f,�H�Ģ�Mv9����hmor�L�^JgL�hO�/\)���oRg{e�_U��(���S�c���x<���)>�͚�+�wnǙ���^��pe����{�(����|�����v�X��Nx����;G#6�N��M��>��ۺɗuAP#��W8V����ah�mW̯X�Hu�y�sv���n��Ӹ��NjB,A`_��[��rܱТ��,U�vg�ԏ�z��2���gnX:Nb;o:Tqt�k)֣�'�ŏ�{��%�-2�eQ$c"-���'���~)�:J��:nD�NI���>��72&zh����Ɨ��V4y����Y�X�`e$��i�W4JpJ`�����ta�9v��;�����M���+��r����8{��5k��"���O�����h�=^�s����g-�w��^C83�u^�!���!#�4Q�e�"�
p�K&�V�6��w`u�y��d��s;W�h����r�/C����Мעi�OAM�}W���@:�Kl�`$��Z�¼�Ll�S�o��t�c=�Ս-�U�]+Y	���5�29��z�ky�7��z=�R�t��26��}�>����Q/d��;.wف���������[�q6��ٷ�,x��u��~�@�����M��d(��^(V�6�TYA"[��.�����S��p=>{��������8���ه7��5jD<{֯�Y�"9h�@���3xwq~�1��4ie&M\&4r�┴k/]�?+s�bm���;K:��m�8�^n�:oM���X�Vv*m��/����
2X��ٺ筳Z|Gt'�i��-��� ߪS���N��Wt.��h���:���K��|��-���v�J���������}[���GPrߧ϶��|D	��EC�/��ɼ������jo0����3��mu��j��Z'��.�
������J2wu��W?.��]�א}�3YS3�n�c��4���7����1��iVӭ�0w��Ї	�l��۪����]B��1�h=��'�'�?\�u�~�v�{!:ue�F]��罤{o;`j`�m��"�uY
/s�!�����U�Җ7�a��k�&������f�NE����*���J:B�h�s�&6��A���/�l!̈�͋��u���u�蟚�C��d1����N�;��v�$:L�T)n�ZL�Uƃ���	�ێ67t�e��l�%�y
�{"b\n ����dgg6ef��So(�ٕB��L��{����"����<�Gh�O	��_\ޑoo�.lp>������S�N��Xd�bVe�j��G���6����y\,`��}��.�C!c�躄�c�b�Ϲ��n<|����k�I�s�����tD"���ǐ�J������og��ĲX1�m��I̧��9��@�zq'Ii�B�дk��٬�^��Z��jJL�L��'d�Q������:���={��]SKP�%[8U{~�=�x>��d���5>�C�]��[=y^��c���K�h&��ўR,w�5��54՚�B�ʢy�k����w�A���;�;���oE{�$����1nlƊ�پyL�XoR�e���3�~6]<��aZ� J��˲�߁��t�-��閏(=q.��<��P�������d�__v{�f�<b�,F�����5[N�ޣ=&��ڮ�*��Q����;�0�i"ѿ�>Y�3ϵ��|~V����كҞ[7u��Ye8��@�p�)����6z�]��\m��U�X]�Vmod+��UǨw�x�7<�^r1r2j��͛�ԠQ3�G;ِ7H�oZ�>�;^���dt;a���o�K���,@�����*j���#훷�o}�Lb��5�Dot�v}I�g�v�N�[���H���U�Τ�0����mO{;PI�-d>T�G�����%���K�v�	�n�G���������ى�%e���P�$�hG��L{jys��`�3��]Tƾ�����-f&�(i�r�i,�k���=uO��m�����u{��t�x�C�g(L��C���YK����Y�Rc�x�e�)]<��t��Z�Z�hl����U��9��.�z�uh��JҸ��F��i��v�Σ���i��7N5�٢��F�0��q���7�qj�Ѹϣ�[k��<���ض̹p)6��`^�lAv��	x������O��l��d�y�i`;.Ʀ�"#���66����%�&�HX�૫�X9܁P��:S��*��bv eM.�:*�BV\C]f�,
�kt�Bv躷;�,���c�/o�~CU���ܬo�u�6=�C�nc+*�,Ұ`P4+�g�{97�(����$��<��"��7�%�쵨�N�t�zȻ�.�߻�րeF���]�oY���:^5D��՝Ҫ.�㔏��e|�_M١6�LwN�=��54� �
�Br��}�6�������c�*�(qw:�8�Sj?�N"IB�lEA�a�V���ێ��*��Z(�>��I0�A?&�c*�׻Z�DX�t(�I�֨�3�p��gH%T`+�Xї�I���B�c��}�N�4� �I�1��䳔�]���$�$d[/"��o�Z=�0�H�{s�*�`����NDo���\��V�6o!#�Bv�T�΢��G�re��i�S�����GKȟ=�笿�a�����r�`��I�0{*����1��o�tWR��:���V{tN��4�����}�U<vu[S���;�Fa��)v�P���{[v�
�e����r��n�����6�s�C��<fw���=�35B������ܨZ:����Đ�-�9����͝�0��6�!�8R2r}����j�����V��8.X������_ϱi��>���>�Y^xR��)�2�u��Kw\i]��o% �S���0w��.ȫb�5���R���y�N7�Zw,�x]��a�7��d\��b͆�.�iU���9��
���:� ��\k�C�ԫ,�
�(��OuM�V9 �X{�Ge���B"Z7?�����
�6�(Ƴ;-�٩�X*�:9��nֹp�Φ�U�BYf�E"���)��
�`q��ݮ�R�QU���.��*�-�j�����k�˽u6u��m��2��f��.����*K��
8��1s$1ˑWq>�J�!A0���\�WC���wHmn)��[(��mvw�I�J`n�9JӝրX�K���srJ$qVʺ��ź����ΪAHr� sz�7w�f�Un� �Z���x�Sw�j�y5l�����`��s-��L��]�ެq�73&T��L�Ա�V)au&� ��N�Tyǻ���h�Fu���o]Qɉ'J7�6��Y�6p��qhmwP�������F�v��G�Qdc:p:��ۙXܠ+*�
��L4��e�R��J[�=��o hҟ�WtU4���jV�&�����G�R\�ͽͫ�i��6�j^p�O�T;Z7�bÏ��|-���s��[��$�s	�Ș��n�F��0�����=B�;�s�z/9�_�s9�j��V�6�io	��wW(A����I[�M��F���M��N�{du!r�F+���s�8`�C�m�Jl��v8�.�4O��}���l~��]uT�P ��J�UQ�O5R����J�UuJ�#-��)�-��,��Ri��z�u��\):\�(���/X�'�Y�x�d�G>�JJ���]t�B�ɬ���F�,�]J�fڝ���K�ta�Z�g��l���u���j.;n�]�h���8 ��-q��]5In����Jz��;:*��=���͘��,��iR��1�	���p4v�h�zZ:nɩ�����7b\�
�f	Ky�\�bY��%�h3jJb�C;Vb�&rB�G:YK��R�ԛ@�,u�+�Rtb���ֹ�� }S��h���i��L0ґ����-	B	���fc:�=�t,v�n��N�&F�`�<���3mU��Qv�O\L����le�J�׋��4�'[t��u+rQ���c.�v��%wƪ9�qܲgo<���!�n8(qW�B��l�:�3�`]�i�v�u�� ˇ�SK� �ۭ�#+Aȝ�Ie)��Qj�M4ԚiK�s����m��j���heEv��c�\�Y<�a6�$>�D<����x������4���a]Ζ�^#�^�1G'Q���k��7hz8�4'6 �oRxa̸��4���WA����#�v3ktq�8�S��չjw>����#���BB�Y�H����5����Z�pv��玞W��*����hi5ZL���̒��᩠cb��R.K���j��m)�Cl��V*��v���j�E�F6�[�Z�n��U�%;A�����`�5<V:�X��sκ�tlqEɘDª�v�"��M�[�%��^�6ؚQ�U�5�+����G[�m�v���z�1��.��]��J��*�P�A�V�T$��	b,�����n!g�Uiɹ2qtL�d/Wpu��v��
E�6'��xa�K�q��ڮ��!�Ѹ��u)�O�޶E����c��v�i&H(۵�v��'��3���������ZXj�i�y%��0�:��"�mX׭����٪��kM�IZJ�4 �fI�#0�?H��u/M�����J�Q�t}K��D$zL$�tـom����w��Y����>���Z�;��x�I�P4�L4Mڸ���CR�-BcM����A����4��n�U�:��`@#�\�<�ɸ>EZO&��〝G���Lwu����v˚蝡��̲P�6 B/���U�!{}�1a>�zWÓ�~��qE��g�bE�c�B�&�)f���я��E�L�9��ùxؚ�*+۽���N�B`2�"Qn�7_j��ጘW���Ђk0 o-a9Hy���9����se�/ũ�H�s�rp7���0�J�a�����Uی�[�JX��wT6c{^��h�Ғ �笪����w1o�=����C�'�����2|7����vv�xE�,
������}��2���(�"2�ɾ��A1�"a6��i�$GB�W\e��4y�5=�����p��F��Uw��=�h�s�Ӟ�,�
�����GhV��v�~5e����rl:��	���������,o�ߖ�����Η1+>-���=p����|�)���I]� �[�4m�p�ņ9�k;��O0ݎ�\��>�{j�^��7:��L}݊��䋞�s��&x��[�^���fc��:G�Ŏn�VM�C5��k:��q���	����9<^�V�I�V�kU����$����y`e��-E�\��\�{�F{��a��@�p�9a�~����>'���B���U�޵s{���NM��wS�r׽Z��T�{Qg��b�	�9�#��.�|���'�T���7F�d��	І|��8��ˇ�NԬ2�9�6I�s�G���l
�>�l��?�����Q��������]l��wQ�ڰ�����x�՝�W{w������m�UKfvNvϲ7�m�iT��o�p��)���>�/��uo�#��c�D
v�B�W��aqtY��z6*u�T�	~>'V>�K\sż��f�&�qD]V[bL�f�F�T[�Ե\�Uv�<,�!S��x�N���Xǀ~6��}Ɨ����;�l�W��y�ҫo��x�@z�����s�K�I�P9�m�,�γ�/����;����Լy]w"�:��B=E)�nvE����T�̐a)�z�n�ڣy��{\�1A i���~:>�3�ܞ�.ĤoZ�Ǭ׬�����0���b�������V���՛pg7��%��"o�|d������	��e� u昪ae�¸ϋ9��&m��ڇY�����h>E�27�R<�Qո�]Y���T�|8m��L J�L`��js-տ}2򆉆�
w�?Jѓj.�[�٤��
I�l���%g`�Vc*$��W�f�sN���1��>��t~j���2a;�����l��u�u�@ �R����-K�j�Ō�]ݕ�mE�z���t��ɹ�����S�s�	�m��:���+��{v��M)�.�בR����)��W��1��Dg|p��}���~΢�|�aq�7m	�52���7����o�8�E���A�r�NU��꭫�}Cto>�yt�w��i�`���\9V�8!���|�1a�99����V�1�N�G�;��1���8�����<�_�����d��)q���<r\�ׅ�,@�'�;uO'�;��o5/�5m�����,%��K�1I�`�t���e,�$�e �����Y��s��g����xMV��ʖ9�Mn/z��%�A�Ge�;g�\�W)���OL�vM/�x���NB�M@���EIvÿS�E��O���Ǥ�I�g�V	Jz���=���9�]�+5OzM�:&�}���pr�"#��~(�U�[Ø��K��6��c�����*��'�s��S����I�DJ��ˮ�����D��� ����=Qh��깚�F��:�/>��t}<vyU�]���H�򂃂Zh�G�Gh�O3\�~���t>�͕G���F��t��<�فpH�ǲm|�)Cku�W˞��NՍ� �Y/��:Գ��o�ͧ{W�v>�_���u�!(@v�Qp����i�(���I"m
��$�,y��;!�eN��kOcpk���V�X�ہcs��m�8먔���l2٣�-�u�!�&�6�Qj���K����8a�aaK����v�`��Z��4(��V��ؐt͍,�[t�֘�B4�DҊ5H�܄� Mn��k*R�/R��	� b:Z&r�m��a�՝[��`y�D��]���g��r$\����ō��P}��^��tY}�2Fׯ����TLp�*@kc��n؝α��W6[A����1�Ʒ�|G<�!S��99�G�����b�q�1�w�g���
����'or�����[��r0�&��qS�}q+�h�K�M���>NҼr��=9�{[��{%��1���ݼ������q��]�l�֙�7"��=c-�8z]R��l�����J�}���pG�Y9��{aԻ�+�%��o��}�Hׯ��_��G6b��Yw��FL���L�6��l�;��{ީ#`U�T�����~�Ro�f΃��:rTw�����N�ҭ�*������V���K�����c�S��"WP�=��E&Z0ڌ�h�/%�}]˚�?1��8g��PV�����_T\�`p��M�<.�F'Lmgu�무�t:�$,�g�TN���Kw��8�K�4�-� x�o+�����Ոh�J�^�k	3�_��GU{Fz^S9�~�qUכ+�g؟}J3�g)�3����8���3����E�D��+���dQ)g���'��x+�����6�?��a�/��s�.i
��gn1��/|2�0+�K����Ys)5K��>'MfQ/��*�w炆�x���*�ʋp��SKZ����n!H��s��Y��DQ.�����CTP��PG�W�z�gx���^�����G#��G4�d�B��Q�)kxSX��l4q��魗E�����@�KX\ˊ�B�W��K#�aL�S�*=N;�qѩ�do�*S�3�/>�6�Y�M��v���y�xQ�/n�K��$�`ᐂI��Hh�;bF��g|�f<{vʭ;�=��������k�.��c�F�KbC�Y_WU�;G���0>���G�wF���4�;�us�����?`8h6nG�o��B0a~��0��9[��a3�[7�]ޙ�v�`��|5z��
,�XW��]�*�WWߤ����".�]�f����p��QuP�������d���C��{���x�T|ylC�apEv�=ؕ��� �}k?0xUR�oV*Z\��\2{������"՚THM
���2���惦./�4�+�ZN��}G��n��-�z�xW7Pwe�\0F���ٰ8��ڬH�שtZ��浈+�s��ԝ��)h��9\�O�X�d�d���w��'O1��z�߽w��7�(���XmǞg��u������ۢ��%�ez����[g��f�1]�Eg�H>�^��p{��p_��1�]^֬�}���N�����K,Y�s���=e>β��Zm��׶�ɇ�(�6jS�A�V$
^��d2��ݭ���AǮ��:�wO���X�����8���p=f��x�jMU�^�LGm�/E'Փ}<2��h�;x�$m��Gz�oݞ
@�T3;���l����J�f��٪���bX� $R�s�Q�d=~(���罣8CW�Ԑ���1U/���oM��+�'��t}�Y�v�J�.=�߳ىg�:���_�̙�{�/f����aɥy����NG���a@`@��"����y��]�B&BY;�Y~��҃�j���3�c=J6w�I����A@�ޱ"'C7F7���^�-x<��I"MF`Q"�#�{��Gj���7Mi�(�&q2�TLiH+RVS��Z,丿R�iH3t�$��7;�FJ��|���=�f���Q�4w'�|�5��;{b�Ö����TQ_��V�|P��	�X�t��c�>�k�}���K]�p!�j0!F($@�A�cf,&��Y�����w����8n6�����#�;�&�Lz��y�M���ʚ<+�����N��Ʀ�N�ʄu*ޒ0^��}yY�m�F��Ŷ��M����QAX��Hm�[Z0%ǵ��x����(�%��<ϪO.�d�y<:�X��.;;�g�q��֗3���ͥ.	�a���ϡ �]Y�;q��.���V����][S0�t�ܘ�J0s���Ps���(*������Bl�\
LP�a��:�L�v�8C�7>��#���9x�Y�\<ߚ��ؠ~c���o+w��=�.�wT��c�]x���bs��/��!�i��)̄iP�r����x]�_o�����D�Td�G��rx����_\��p�>��;}��q��BM@�ۙ2+tj���J	L���]o���8��e7�o��hdiR���kNG<p���#�v�<_�S�^���?`Cc�u⹅�ЯE��p�ۣ;�Q~d�wk:k���@\&Fc0(]xט��9�ʑ��h��t���|E�F�W�7Wq�q�ZMT5�`	k�GY�	;��r�.;l��!h�[�-H��Z��럹HΑ��ڻ�`��l{�v�{G��F�	�ᜨy��t�ɞ/v�=@}J�%d�iT'ܐ�7#޿e��c�<�U���{��H��&k�w��Q�"�t������d�����9�4� �WvL�5�==��<� �-�w(����OK��;�i������B.x�D��&	�H�Z��S=>�*���Yi��[�Ғ�s� ����s��兆�O,�.�3��i#ABXp ��M?6C�b��1���eQ�벺p�~u]�
�gfb?W{������
T�,I�-\ˣ��st��7Gc�vK@�-��6�����Y���:�3�\�ۦ^�|�S'�2��ي@��Hn/K�����&�N5f�e����4�΃F��M`�=A	*M���n��^��Ec�/����	�a�M0L�J4m�b5��Y�����ksa�>�����m����7,5�ʹ�����s	NiqlK�F���
�Ge�X���]slX[�b�(�bV���e�JćY��͇&.Xb��k��FXA�P��&6dKQ{��VM�G�n+��~��ȁ�O]�oq�<9>�j�r�Լ����DbiDa)1,'8M���c�ē�Q;�J����}�����۟+֓�;�Y�3����:�R��n���i�١����"������VU�u��}=��Q�7@��6�1�[!��Gq��~ͼ��V�su�t<����fs��E@��I�-݁ڲ�6�R�wⵋ�c+FS�e�ksk����p��z�O������3�jW?@����-��®�娰��s�!3�~����s71o5n�R���MT��N*���sO1CF\��ޞ�m����/�m½�fv�LVH���Ɠ����
÷8����E��y�U�!�cz}R���ϓ����a;X�Q~UB����tF��E����u��n:!+���5QSy%���I��Y���c�q��}���7ϩϗ/Z��~v���n����s��\i4�$�Zw�x���_���Z���tױ"��{�z�y�^錉�<���q��fA�p֕v�s��	��!�s0���i$��u����u�X���Qr��3��bW�Q���R�QCI����/7%g^mT���(b���W�n)�%�xx_}�x�r�����Ϙ��:����g�O���0���m�E��]?<Z;�]�%���I�B�սt��uY����	Vw��?O�I�^YUf��3����%�4� |�@[�v(�l���ؙ��i�C��WW����J�E
��ɦa}Eخ���'8��khuìԄ��i&B������fm����O
48<��Қ�b�h��wWu{*��=r��3�F��`5{��6gyĈ���Y�!M�+����f�reP��,���?]�#.�->>��sَ�v�|���9��~�<
Dw��e8��%d�^��3I���B����B�����Np�5u�׽#���b9��˯�w��3ѽ;���u.��6���V���i*]�c����˜w�ܡ�6��I:�w�~���o�C��c�����?�D��٫v��0���fۯq�����E�}4��Et/ܾ�}L�f���C�h*F�EB`0�'^3쿔�1��3��&�����81�g*��,�[}]���Wn�Vh��;5]�n_tP��X2��\�X��ɪuniEuG\��� 4�8e8E�޵�1�ؖz�hp�B|��˴g*���a�Q��H�\nw8��v��5�b�U�p�3-|"-_�ƒ$)5���y[��<F�o���ǫ�����.N\p�oj�wg����Lj�M{�!i]�y�
=��q|(N��B�Z�������O��H`�<��fm�o�S����q���Ѱ��쬛�t@˒0QV<뛷E2�L�G�w����n�j�%AC�q�� l�U�j{�a�;�Ӆ�b]�R�Uc�Z
�=�Nr�d���:�P
��ˡ��z0��9���S'f{&�T�j��B�y�r�K�^�њ;�:�����޵#��C�y/����u>��#�����ٵHM�� 6.hNW��+����e�Z�c%y{M���g�����7TC�o�_�Ӊ��»��k�v�]}Ujޮ�]k�f^[��<�`�h&-�ݻ��`��a(=o���e�x"{��J�x_,CGU=w㹱H��R������z^��q2��P��_ڕtN������yU�r��	�`��;w�rX�F���\*�:/�t�~��R���%!k`pu��p�ks[mt��V�V��o�����$�e��z�7�����ٙղY�k�|}��a�:)<k�nt1�� ���>���[�1�6~IP�v�����^��Uͩ�%d,����w�q���*i��7q@j�;tt�L��s7��YO
�g�9��w�5h�]X��Q��\˯+ў���""e	�4k1`�OV�z�}�z�0�.�f��uʝWL�P�X��I5��Y��\;�J$�<���.u����"��b�u��@]<�VfS����ٔ�Y�'w�4̠�8ZW�WoU��$kh�:�2��i�(�I�pL�qӓ�Q}o�Y�8�G�-$�]��͘����s;
��̧%R��ۛ�FSu5�����̔���ӥ}J�%�n�C*�h��\,� f�4�[%�8�ar����DB�#?Va���%���G�fgsrУ+4��qō�5���W��'��3O姰�T��8��u{X�-d�O)Sb:.�&Ǔ��<�]NV�d˾}d��,T}�6����/U��Q���a=��:��u��Uok�dl�GQ�ӉCsC�6�j�#��;[i�6�ڳ����u����f&Ǜ���Q�"L`�����n+)�v���
�F���W���݉8��%��v@������D3�;q�{u���ɻ�ʑdC���;�W.n+���ۺ�5uײ�u"ee�b�Ԓ� 5� s�r�-��WEc3{����`�n�c�
C@����z^Xu�.=\G]�"J�{H㒮2�b#QEw=z /���Moe���շ:���3^mIN5IEt]r����������l�:-HY#6�EszVK�tX��EY��RR �L��D��"oJ�6�kԑ���ap#7��U-v18�	�A/�8r�.�z��W�e� U1T��|v���z�����*aen�gnjU{�	D�G�:T[y�/�#���#���~�}�(#��ۂ�u(�#*��mO�z�Zڼ���p4'%w��CM�,ڪ�&�h�6L�N ���3y����xv��.@3sfcv'p`<��<�絻q�Fg�I�����UW����	0�>W\g<3�]4Ad���U�5�uB�{~k3igO'���9".Di.���)�=M; �*�W�v+�]��܀w�F)W�z'�A��wT�}w÷�be�����WҞ��=qxw��s��W����Y>1�$e �e�-�/Y�A#l�LY������[�:W���򳻛s�<V��.c��:�Ds�qK�]"{�Z_M�en�����U��~���o���[��M��og���Fd�T��Vc6�ר�����j0����U%��g1Ӯ��$�J��_��ؚ����#BF�R�z{ݪYD�(�pC[�p6����^�8�l���||c���6US�6Lh*u��o�ν�|!\{h�Z�=^/��Y���
͢�@�>ɮ7����I�N��7�Q��Ҫez$��Y�}g�5˔�Z����x�]�d�(�����_<�V]��*�ަ�bX����v^�Mf0�0lq(�9Rq5*���xiG���@0�?0Yhqt�H�H����u�m.���j%�흶�p:؋t�ݷQ���1qupZ9��IS&T��sX����q�X6�<E��ݟ�w�|q�)��Kx�bx$��ٱ�#�*��v4��4�a�ͭ��:��2O=��;������c�<\���$BL-^G�S
Er������+�>�c�˹y�mx�>1	�ܜ�[[قw�{?���+��slg$��R�Ey�q��Jq(�D�N)�$nxO������\6NQ�4�ݿ���z�6�]-|����O�p���O{&N����\�o2�K{m�s��@x z��"�:�G���*˴(7�p�'����c�<�:m0�7۳b��8�����:i��ҾeE�33���u��T����b3st�����Y�6l�{m7k��^��\,�X0���=�t���%]��l�&>���Q�[��&�y�q>��~c=U���Dh���utgM�s�z�Ev�I���.����h�J����~#܍��g2Vw��|A���2��6;~_-�p���Mlq�n
09	��D��e�J<uv-ȱ2��oQ��=���D����k��w����Oh�Yk�_m,'��v�N��,��R��v�i&p�e�qK�\<�I�<�d��S_z/P�|�o����|�Ȍ���(1We�}�{]���;;�~�c��2
�vf�uOO��福��E�G�#�[�)~��tlF���S��x�<����\nLw��ꃕ�<v�v,���8�l���q����eG��绣7gb��0l��lU������u
3�N�wc��B����	�N�p�[�߅�o��fL��MF@�-�����U���;wo�FLl������]7��u<v7g�'���p&�\:��v�,x�.��&��:5�{�1_<$w�ʧGy��`���˺���w����i]qq�N�,
u�w3�l���	p��"��J�SUFg �}�i����:���c6���#0a`>n�^���j,g���V��^����B��m�yB��Ph���=3��ze���S��C�׬*�D�Pkv���e�q[^hc�^�����I|�� ��}bmu���Fx�.$�C.�4:<�DԼۢ.�๸@�p E�U�Isxqd�����_T���k�+���W7�/~히c�x�ɏψL�����G~�/܋��9EQ�5��V9u���(\�pa0QnE�/� �˯Y�.z�S3��� R渟_�E0|ZFN��Qw���_�H�9N^�:5�/�1�|߸����|�3i>�v���� j��`7�OM9�WʥH���k\�R��4��(���9�P���K��H�A�@ch��FN���)�2�����DBX��؇2�4l���>�|�61-�;;r��k-�����)x�{��&�ۧ��n�s6�`"K*�\+�[Y�I���Jĳ��Ti�Gz�XٶkR��?njQ�9][�N&����0��(�vs'������X�$Lc�PmR�g���z&'㾃����g�&�~�ߨ��9�G�J]Vr�Nfy�����5Sۣ��g�j0{ܷN�>s�k8I�E�&����9Gz�F~���#y�f�Z�[~�+�2�d�+k�vj3�ɮb��u�,X�*�ʭ��z|�����m�y�x3 l#+��[�+0׸��I�k�����{�֦����d:9׃��N��s:7��_��������w��E)��
u�;��		E�3���q�+�bmw�l�x�u�Y}e�V���$�o}b����v�P
59Ҷ��)U�A���}��U5a񃏝�}����M��0fy?7{4����44Fұ�< �5�8
*�����1�q�;/d��$%5��(:�ћi�ʘ��	4^}���������yo�{�<���o�
q�%)�|&��{nd�0x�_MQ����t6�@��2`�'�a��?t�}�pt�p~�sK�����gZ��)zP�ױv��6�r���yt|k����R��z��e4�	���8�Ӟ;Z�?�@>
��ZW�.lZ���d�4Xks�w�g\U�5�g �v���Z���VJ?�.VûF������H�ng��.�.�<7vk�xe�W��u��Q[��������.WCn
Y�^�^��I��˾��{�Ԉ8A1A�E|� �Yq�v�q8>�l�w�B6>3y��Y�н#��ž��l����K�����O�Z1P�*�˞�3�:
��ۂS*de������C�5՝�����xg���*4�y�8�&�^®-	����F��`��wp3{/\��8bD���/�*]���CE7	�*ھ�x/��C�{��Z�2AP���ݥO��}�)P0`jRi��';�t-���z��=<t* FR&I m#��n�Ҵ<��6����Ֆ�VqWQ�����8��\�ܭ}ޏ�����;'8�mr�*��L(p
Qst�ZX��B}��ɛkR�mҧ�������7KDOq��4 �c�琴⚼v�]��>7͝9���|d�w��Ǯ�w�A�[��8lX��{Ǧ'wM/s(�IF�:�?A7���6z�n,^�<��>}��e���O�,��#SD+�h����:�֗z6iٜWu�]fiY��QN|~�*:�b�I��WTl�އ�O�Y.9����p�ugv�\�O%۔�w���d�Y���+QJ��C�pDP��x�omcښ���h�[1�{\��hSu�{Y�'�Wo��Il[O'(\E��F��������|I�".�)bխ���aYu�+����uR\��9���0���,v3��:P�G��F��0L��#��sJ�A����C���^�ҢJ��X�61�V5�S�^�nف��.5�J���:�0$E��)�]:�k��b�ۙ���V�f������1��M-�;�F�i�)q)����q߆�s���?�dN����.�FO]?y�Y�ȓ��u۾ʏ`Ñb'	�!�
+Aξf�*�ڭ�#��}n� � 3o�:���oC����%�����
�"U�om�H��
�γ���_N�L���=���%8I'��'м2j]��=��.�8J�1�=,^����>Ǜ|{|���,t���Kh�n��q;\/����^��L�)�E Kp
JM��B�N��Q��`�1c�u��{���e�X�M��O�����P;��n�}[D�w�$
I�^�`a�v/^�<�ؤ�ꮺ���\Y���������7�6���=�� �}����O�h�*��d���-�b�d���/}�������_����L�
;q�9M{�6�1k�.�\���=�}/�^�p��Y͑���p�Df�y;���ޒ�I�P	������P#VԴ��	X���>�U�7Ʀ��J�C�1w�����#�Gl�>>���շⱩ���4���`�ýM�\"z��feح��̀�2Ԑ!t��L�6�z�v��߅��xoų�2�M0��)�����~�)�넬��[1�S~�a��&�� �Y�;W9X7�m��DWHuOk.2��`�����9�sy�x,��.t9��7��`�?$��>W�=�U�E�~�oDE� �j[�_���w2��/��|�{�p٢n���@1��O,3��i=�&ͅ�.�E.�3h[�CI�h �p[�L�����K��tG���^cq3��g���tx�n�u�_.�`�X�{�vf�~�ѫ�M�� �_e�̝~�m���g��n���Cz��'g��
3�>�;p��yNz�K���uڠ�zK��5卭혭�;��l��Aq��|���U�ŵ���V9t���d��<�w�>��a<���=�Dx1�����MW�vI��c��*n��#��V]�������7�M��i�^fI�S��F�.�~�}�����b�Qɐ�X�"�!ߍ��.�S�o�#��dy��KN$�����6_7Ąq'r&���.xw�f�!�ؐ�\{�lk�I�ѭ�.�<�W"�{��U�e������C�<�H�e�˪�]*�A��&���Nks����ȯ�鳧��0�Eb�U+�ǉ�w���4\�ŏ2�J�"��2@Ocu���r�T�\f8�mH!��O���m��6�c����zv�9\�N�>:���is����R����u��lN��d��g�*���Z����_�f�x�`��������yO+�<����i�O;(vLح��6���u�PAO���>�>�{ϲ�n��#Ѩ�rH$�����+ip�K������ك��zGC^���Y�$}�K�^��k~>?���:������
��SL�b]�n^oU�ߗ�o��������i	���V1�x@��/}�ΐ7�錝��eo�Dń�W��/`�"=*�\��A/u���wv��)u���k�Ch�fz���$�2Wl�f�g�%ɰ�d�	�D��[��T���%gWgV\oZ�d�.;m_b��Eʭ5yw�`Q�.��N�
��|.���s*�9��Z��2��Pu��Lൾ��#E�oޙ���7Y��P:g�����}+{�kx�{����A*�K�w��B��t�:+�����<�`w���M�0%F��ێ���ϴSԅ;�â��0�4A�*r���fM�FP6�"�@����Ys�~˽cw߅<���r�gƨe)�����~�-	�~���:��l�Q��S�I�`�Iq�&�:�J�d����%O��-O=Y�f����-�_���u���~a�R�������_/	���6��S�Z��FM����7�~�=�>�H`��a�p����t�8�M݌\ ���Z_k�A]"Y���%��.���*�(�=[��PE'NA�a�U��mgnJUڑ�"�u�?��;\�[̛F�u��b�r��5�G�����u#8��xkg;�,�C#�����m�D����qA@M4[`22��{V2�ʰ���c��T5|��Y�z�w��kTd^�\Lż�J}�Z�)�|<%_o�n�f4q^�s6�O��Vx��% ����uց\pg �+����)��=ش������pBpm��gQ���>��b`�i�f�o3o3��𒼛��nsT��:�쮌��Rh|WȰNf5���>콗�)7~B�������7�~ꪭ��8E��-�$���F��K�Z�6Si�BZ�DܐM�T"0KE���6
�Z�;Y�!$(ޗນ�WB�,�2o�H$;Ӗ��<<$E����qQA82���r��{G��(_�)��Տ��=O'�ƴ���y�����������w�7:����h���s��ԍW�
�2�v��<���|14�c��g�N��A�����]�#�����q�{�1�B��>����pZ?z�"ٗ�����˶
�)�vxߡ�����/Z�k}�7f����<=��l6���Qߚo���Er�~}�CҞ��^y��޹u�g=B�����n����������P�F�6~;*#��GW=Ηu�KU$�o:���q����!�\f!�S#]UN��D��]���.T����n#e�2�]OS�� h�ۮ86�sل��ig���o/��R�ѤBؙ�Dcl�-m�2X+�ű�%Yi�woL���\�bxh����O��l��g�`�w
uځ�l�P���9�B]FSV���4�BZ������c��]%�K	fu�$�⛩`iQ�ssX;��Xk�0K�[q4+ �d6	I��'�~�)c�	%W���w>�T�4�!�jg�{�N$���e:�59<x�|�<��^�c����4�܎-�1<v=o���'4{��Äy#��%�m{�O�n<c/����_tǸiWuN_��v�6:M�l\*QbߗL߼+���H9�=Cv�y�k3O��E6�Q�"�ŕ����mk��0ܙ!���Sch�k�<%-'�ǵ������9V.9�d�c�l�3w��_��ڽ��nn�|��#�J���R�*�N֪����XmM1�h[6��cø��9���Dc��U�1!�)�(0X��d�$_�+�{[<6���z��ߡ�w�ג{�v=�4���A7(1s��k�>�`㼜�����0�����މ���.}�^�8p��F�B��D_R����z�k�?{��U98����gnUo��z��X)�a��{[��];��|)����O�/-�tǊ}6����H��}��W	s��"���2��2&�Z����>���V�����8*L�L����]��p�;��|\��v+[��?k�o=8x,7	��{].�ͻL�UX߾�[50(������T' F^ah5��y���m��H����h�.�����S��u!+�mO�$��уu:������Ļ,�U�cF�
��}ӷw(RTOOX�׬M%�v��w�K����y����EG-ĕB�<v<�`��ƳP&�j���ʳ��r�QJ�Y��s�Ve�Q�xo:\�s��A��K�ݏ�9c"XU��k �U��AH�m;rqf�8�&�8�GV��h�`�.�t%��[���"2):�{,u��y7+�H��[�@��K:o�z�Vv��<��px�e��{�ol��3cə��=v��uG���J��;Ky]�@lbw��9e#ڊ�܂�Y���v9ՙ]�ށZ���m<�W&Ú
ܡ$!�`���YB�2ֹ9ޮl˫��j.V��G1�:G\0t��ų�m�w:�T�x�+� f��=ws����<�Ыc^m�o��[�l��T}��m��}�e'��ZѮ�W*�l8�+%d�3AJ��қҳsd·�S$J�Z���ժS��{��,��e��l�0ov�Nw;+9�w91�X�;X���h��A!���T�?+L�a���71� s� ���i�їXd��x��qf��f����Ӯ�O]0��y�!�6�����럴�+*�P��vB;�[ƻ�H�"r�ZOU�Γ]�<�Qޑ�p�X_(s���Ukm�bYu;��ܗ!J��L���<����(�E�}ǖqL��8X�X��rX�7}v;�ɴVvh���+�j�%JE%5�T��B��UT观k���d�;R�QUT��*�٥j��ET�K�n�y��n#�օKCu��v��u��Ӹ6MY�T!�|Zq՝�t�WY��X��n��Og��C�,;�)�Z۶�9X۠d&��/
�Ua��)�f1�r]�fÞ�:Ǹ#=ٵ԰��Pm�����DY8��:.
���l�v���K�c�.����	�'���:��vNú��s��: ��L��Ճ�;@i�ie�*�ģ�WpݱKn
��QЙɴݥ�(��v���J[omT;F�����GLJ�;B�WVL�9Ԫ��&\N��7;u�$�NGO�V2�3R�r$����S�.���ff�78��e�5����]�v~7c)=ET��,%ۘM�kjR�2�G4�ܝ!V7d�n�NԺ�b+�9�g�q�x{("�x�x��q��qZ|rp:�gG���*�"�1l:]��-�K���GM�ֹ!X�6�Ya#*e�Y��M/V��(YaBȥ!5К�h�؀�cI�^.҃ۧ��5r��\�;�:�Mjm1LC^��f����)����'�R�Ѷ�:Cŝ���q��x�Z#�8��Q�t8�`�n����n�Ʌ�e����l�wm/o2@�ݒ�yݺ^ �BHgvL%�۶�H�j��q�:���U��s��K��� (p%�C"<a�,c��װ8��t[1���D�tn�]�[�5�BP�9��r�:��ׄ
U�H됋LY^�6gl�^S�k0i�q�ϊ��g[�z�d\᝚q�fÆ��Y�����^Cu�l���+�磬Ť!�IX����
�tk*�bLֶ-�Z»�BQ��[H��Z�1���4��<bձa��Z�`�mȼ;!;���تLnf,���t��m-�Mřf���-�mS���3\���4� 0��Q��SƵ3\s��n{���n�cFQceLb���f��vd#s�0�Q�ĉk����ZvFg3pAv�BgCQ��sv��`Zk5,$Æ�.$"�'��?h��k��$�&��v����Sg�r��� �?3���+ڗ����Ƌ9�ݎAв���Z���q�>o2�1&C���K���i�-+�\�i
��Ɂ�I���}���0ȼSa�F� ��חF�X�x��¨�U[If�{z����%������G�s���շ�S�k5�^Y�p�#��Q�y��d��8/{��>�+��{E���_��F�⨞(D�k���
҈��S@4�$��0zzez�G|5iD�ڵ���G^���G��J�T��ˎ�vOm|�
��p\���*��Z�A�[��x���׏�{�s�pԇ�6��H��޵���,e������f��y7�3�~�ˍ.�>������U^��Gі^0N�ٮ�X� Z<.+}t���p���E��0�l6f��q�}����9���_ӟ{�9ۿ���'��u���1!P�ot�:�1iv�h�=�x/�{&����CJ��;3�y�����F�R5��9�Z`�|��90�J9 j����J� �� 0�W]��6���.�E�N�«dBN�/�ր�^����W�*�N켻�S���A�ǫC9<q~��?��r�_M]OkeOWWՃK�.��Z4C r�Hy�ΠՓ���xCy��K0eu�;{6Qkr���t%T��&���Z3%e��V=��Һ�Ut{O)A��A�X�}$�y���>�{)i��|@}(x�}P�� ��Xv��kq��۳貫���A�6bzo��y}M��V��~:�W
�.���~Fh%PI�g;S����rP��ɸH�ѹ䞙��eOO٧��c�U�w�y�|O���I�+�Cx�Y���0U��ʭ�+�f�2y�ka)�D+�hg�ZT9��7;��k9�Òa��ɠw9s��ШK��0vV=\���q��.�uNo��T;��0ܾΨY��l$T$�JH�V����UḼ�f�;�Χ$<�c��up�^�3aV�C����d�3R�{�3��}X�l��i�ϮZ���d�#	��N�m�=��:�橈Y�Ŋ81�o`�U`�ĲD�(���	fdS%E�X5�3v.2JJ	?�����-@H�M~�u��Az	��<U����|��h��}4+990~��4cʢ]�Tї���PKd�Ql&�s��+$�������?������s�:{�m� l���Gb��5XEW���\�i>��;�� *:��W�� �*8l�����:�<�?=��?kث)��լJ��a�)�Z��;+.��)�љuu#ȻP��x��P��)������'A
��T�k���=D������<VҠ�K�G�����W��6����޶�����E��А��WC��ʌ�ɂ�P�l1WC��WR����t��wʰA��6_R�;;�q�.�_$jJ^���bG��{6�=0����o���`�EX�M��WOf��as���*�ʒ.�"��d�1�!=Ww�B�ujJ���������:0X}+��Z�v�\ڜÛ�eU��g�U����a�)q�*}��훫�����h�؆ӓ�	�R��+�ӯ"fZи|��4r��E$X�Q��QmX�](��,M\k`&,uU��	�
�bh7�vn�ȯ���Ü��e�:\�o�n����;y�^����]$Jc��Mv�\7:	/�a�8m5����{�������<���@�v2�_�ȫ�K��+�
����+��sx9{Hn[����W6�J���NK�gLe���4 P�,�̞��=;��<doz�*g��c�Kw�Ӂ��#��3r��W��&�s�|_�����<��~�+˞�i�J�jkA�7���(*2�mV,����f.C0RpA9��8�͘s%N{�)��,f�K���Խ=yb��&*=�Ҝ^F>����89]�+<-],�h3lj�`�����xtk����*s'`�;y�.�z.j=u����:_5�����om����Bh�JI	�4�nt��<�Lrd�x��Y;%��D����#G>�[[��	]Cr=������;����5\���픃L3f,X9
[����Yk�iK�IuJ�k�F'tsv�.^L���\\���@��ӫ�*�y��ɵv��8��l9 k��'�)�n�ܛ�hReˬ�%���h�64�JF��#Y�q8��~��NEO�wz����p_́y�\����5�T�^���;��s�%n�`��&�L�\���<�.�m
O��Z�I切ßiK�齵�pnտ����t�k��WU�(z5�wC�3ܩ�&��w�����-  ��$�QU���S��"wn������}��練S)�� �U��%�p.^jT�6��vH,J�t�VYQ�F�p%�����=��ܦ׏���O�ٜ�� �:�:>�-[_����r�V�Y̯U�m(��1���� 6�!(+ Q�6mu�j_b���[������C
�:�XV/{cg`�k�C��˴E;x������GFr��;T#c}�&!�0Z�gIᙫ*�Ϊ���*�_���ׂ��9�d��/��_,�ǻ䲯��P�pɋn�7�Q�=���7������C�7�	�Ȓ[A���:w��Iu/T׌�A�(0��uܫ������]���>�w���¯3'
����ο�b�����ފ�*	�M+��jǷ|\��p���E��F�x�[^)��d,�Q�;��͊��홾w`!�z��
���BZ�+gw�_��ѝ���{��Gmc���l�F�����H��Z�:y�闖����cGX8w����Y��͇���u�oA�SP"�ɫ�?�s�A��㱐q�ɇ���t�b9=���ABe�&@S��`*=���$ޞQN�W�^��n�.:B]`��&5>JZ@��D~j2���̾����K]@���>QBQ�d%��;����&]N�g��vb���b{���v����k�õq��^����s]4mAy~�a�ڮ��R�>��Q�[��?lT���������ᜬ���Q čƧװ�N�+��͙�W}��b��\���7<
��������ʸ����n
��lW����iZ=�^�c��� ��>��I�G������3�Ӷ;�I�����#��{��r�����@�a�%2��
��Xޮ��G��}�|ww�.�#��'
�aN5ũ��αח�I�*|����j�n��/�n�Q��ʾ���[М6\"���)�������l���=3&�z��a\�:rz�ק��D��P��|j ��ӐՌ���~�)_�z�E�^�Nx�;�{��z5�B��Lz�}TdA:�W7z�D����ǳ�3Z�R	�2�Cn���o]��m%oA���m�(x9�E��}n����r �r�+r|���"_,��5�`�� ?(!�_k.���ڻ�f#Y��;�ٗ)��J>�R�r�6<s)�̺�#�P�"�X�u!�y���6x�J�u>�n�]��t�}3;eM�:
�
���h�c=�v��f/�7<��on�7�=��!v`��#��>K�u�soJ;9v�VK����eR"���c�TkӮ뙺w�I
C$��p�Tr��2������*{w���e�v�8w]�4�k�|�/����y~�����a�2�ng����Z��Nw���i��6E�Gϖ�=˹d��M�=��k4���q�U�&u����"8��C��3���O�ӍGs0�_ٝ������y6����7k����y��t$�� �pL���݋������<Fpf]���ɳ��'�"Z�Gt���Q��o��t,٭���{���q:�o��n��3{�j����B(E �Cp ��t.y�:��MN��ڝ�|�ͺk� ������ܱ�N�jCn�ō<�Ѯ��l�ok&HFw��w{z���O�n�uyԧ�޼���xKF�hz��',�M��wZ�8W3�K��N�������ZfI�	�m�4�!�����^��S;Ƕ��>���w�b����GH낽�x����kS"�e��D�=�
 �[�KxF�}yw+0f� �f�CA�@�]I],qSu�K�h.����q:��{dի��+�uq~t^���I��α��7��bd`M����+:���5�����qR�CC���\v�:6����`�[��
�SJ���̽��<�.����w��a����&4K��3'�~�����eVvQi�OS
7>�)�K��d\����_5����1��o�iu����t�S�k���<�s�=rO����H$H�뫙�7��x�����e������AB��Lp�m���#sj�U��#A����݅?^�u��o�QS�|��9�|���a�z!�T�+�90���zݼZo�?u�JN{��Əi�O��$h0�!���~�\Vǜ�B�����B��<��8~|�|.6&��Z
K��0�_F��/F8��bqx+��7e�#M�"1 �f78/�ͤ��W��1�>\�|j�j�1^�dv���[�8:k���x�@#ݛ����à�\ [�4]�f��ȿN���8QZR���3\a�	�X.ٯo���k�P�3J_n�/d�����`�=��\֮�͔�E�n�GQ�4N;��\N���ϰ}�25s���"�5�{g�?[�{d�#&k��ޜ���)}R8|:���3���A-��!�����Ġ&��/Q�4�w�'lDx���1Z`���/�d�މ|�q�J����U�.�.�K	�x ����]ׇ�ٵ��9&u��p�%]�9��/yRz�蔩RH�X.�ِ�sy����Փ�qq�v�ZNH���a���cT��Y�[�a.WM7#v)�e/�η�Aƺ5E�id|k)��t��Qr�՚wf�
B�Y�� �G�h��2���!ls�0As]�r�r�Z��p����CgTg��6��+v���vC������ i���4�Y�n�/O�qO��j��tJ͌[e��Xǥ�
!�-('���]��N~++�~j�&P�YD�~���U�w�!ʿd����3�I���\�����ʦ<��h��+���;g0�NwWz�e��ɴc,����m�T���C{�s�No�[�����Z��=횋����o$n	
�]ط���ך��{�3�b��ys�ˋ.맦P���T"�LC+�V�6|p��)�<�����z���V�<j���m���7t�:d|�iY��;�%���xI=B}w�p!b\N�v!Oftp�-�����x
РP�ct�g��Q^B�w8�O��K�G�A�W+���ziD��bb-L�He�xG�J��(���:]wH���w���\�X�K`��L��']$#F�w�w]G��׸�"�&6t���M�=�c�t��B9/�O��nU�SӢê_��ޓ�y�#^�J(�X��Fo����GZ�m���5_(�CrLϫ ϊ�9>Ie*1?�Aī�,p�\.���j������o��j�����.�egg�o���-,�n	J�]�%�M����������B0�)%�q�G�[d�}K���~�uLF��b���/�����t"���;36b�A��K�RWu��P�\�%u�&N���5�:�Pc̀~C+}�xyJɱ�E5����ƗJ�L�0䞜�G"�[�e*+�,�oWWM{^�|C*E�`�"ޮ8b��1��p�=������oa�^$P!&2A��E�4t���u�<a��v����mjvVb*+!�����.��;\!_�H]^��.>Ǯ�([���a�x�v��g�Q�S��Uu�u���Y %�C�T瑙�[y[�vn<��mW����C8��5�J=3;����O=�A>U�gUX�ӂ4o<�*o4ݭ�Q���`$ ��ˑ��0<�WW��'�[�#�n"G���o�7�b2P��@gwq�ܐ�\Ͻki_ڢ�0��.W����у��o�̳��ѣb.!�� w�|}I<^�L��%����7(�����{�ʷ����W�s4��{L���[|h!>�{�^�8�R�$��6�oF��0Ҁ����A;T���G���S������<=dd�>9?`]��F��'���pw�2���.7�?i����I�-Sxp���oޛ���p�-62S�(A�R�e�84'i���¢���!H$ �>&	`y�N��Nsxh���}=��M���Z���	R�_t���ׯ�o�% ��Z����������c���u�z�����sC�/emS+X��!���S����:�َk��ֻnb��X���R:��U�I���Xt>�A�ֺ�� �Rq��&z�o��,�h���e��(wG���7۲3m�+�lS�;�O�u�F|yNU����μ�e�Ǟo��'�6��4m�SOmI�|��.�m�l�tv�=2�J��EQ�?E�&�ٓ��u5,7��Og�M�u��ؑvf�)�9�����~:����3=����}��D'���ͯ� ����x�a@��-4%
=�ș��-�U����A��ć�G���s��r������w�{px�cu3�B��^�޺�-��5g{T��:�|{��	4B-��OO�uTyW�5fxc���A��U Wm|�x[�>�A8LfLB{�tE���9�!S/@��?5&��|����l8��v
�U�@��"����goaH�<����~�6�z|=�.�K�b���-�h��^Z&�W}w|V�5p�b�9b7��� ��Ao�Z���Գe�3�)@��v��gϐ�XFFxϸ�"zv�_t�vU��G�;TIPc����ʬԖ��D�j��S{!؜ɔ��$�4���xeh'�˓7�b�_xw�����rW�����ӷ�c�
����1��ݪ��x�-����IU�Z��:��q_|*uit2�X=];�����.��ˢ�����S���K�aui<7�s�%E�:��>ܙj���}:�����_	{�\�=D�?]^�_j�n��ȅGg�e���gԘ�%���� ��j��F����U"Ɗb-ם��R�9K������W����S[�0���p�,'ߍ�>��B0(Mr�_V9�K#E�vU��׺�()�0]�?�q���m!�u3�%�6�e�����2�6a!���n~��u�-	:V^��[�/9aa�۵J^u��a�}��Ѭ�����f���n�5ɥ�T�yA1µ�ت\����]*��r��y�v�>�$Ǝ�&e�r!��Q����E[4f�kk�A�k�w#�BNu�]V�����9���:�n�E�[?98|����#JD�������W8�ٵ��*S�4��&�r�2��l��	w�[
�9�y��|�yh��fλ.��>�nN컐���J����Ygz��Rب���ެV�k��:-�Fh�"�>�#���z��5�e��c�ب�:�M�)�n�\4ə�?I[�y6��i��<�Ř%����`I~�^�7,ܦ��9h��h���Um�T�-���m�)�vL���b����A ��6��Ŭ�
�ޥo_A��7]u���n�����t���fI��_k�j养Ϲ�Θ���[5���sV�Mᗃ�#U��o9�hJ����eJ��;�9��+6�,;s��q�T7��}[K*7����{�W2/�֦F����1��D{̪�MSw�
��ߥ�Co���~~_���P`eI�{6�g=��hb��P׽�$�{�;L���n!���q�����K�>�C�=����LK�gHG��Mף�1��̬ �;�9����9�F5��Ncu��sZ�t��j�DJ�=��h��焾yv�N�`�b9�nD��@����{,�.���^�|_��M*�H����fD����4�:ʏ����$�}���|+���M(%�tI�G�]Y��w\���pU-��:��i�6BQ)(�B~LM�#4v�n�XK.���GWN��N�ɹ$�w~��(��x��(|��f(�oygu7ۦ��$\���]�K���lי��`㻕=��	
2!�oΕ�㒮�j�^3��J8
j�W���Vi�Y=Dx�zhǮ�&�j����7���9�w,���d��X��g�:�c;�Bk�a��	R7�E�=��n_��lĐz���k����/<�l{y`����������� tS7s�%?gٲ�/Y��0Ǚj��u�J��x ZNI��t�����	]e�N�>f�=i�}0��wc���q��5��C/���cݥ�;pwr��qmW^l[3�	,4o\wIa� �/����q�6��r�3�����xedĹ�2JwN���I$�5h���g���\��M��t�kq%luRU0v�.!(@��B8i˥����}��e�[�-�mDn�����8$�,L�Ά��2l]�<�z�zu�7o�`Ũ1uM�X����@���^3{x�lPu�Üm���ӓ\%t@�o�����zw`KC5!K�Ű&�8
.�k\�S��3@��PTݭ&:n��x,L�6�G�߭�������v}���]��p�Wn�ΧT{L�u�Twz4��a$� ��+.��V �*�D�,��f���������z��zW���}k�m*;֮r�g�.S�7�o�QǺ��w��k�>��V�gGwђcF8q��m8)�C�x��|RT��G�\53�`GG,���x��W�Y��8��k���CW.[���{m�a��
:���T{�
o��;a�³-�����3�V�
����0ڑ�kv)���=�+��(̍�ɾ&{����P����U�D��8���.�l�ۃ�%���JE��7�ʍ�_h�_�M��pG�g�uU~�:��'X��ت��4��p�l���4eV�c�D�V��VG����9��s۝ͬ1�M4vgt��*|�ez8^��j��^�����k�T����`���M-��vγ��|�0�⛀��YW��8Â T��ĝ�~�X�uw5K{;&D�(�]:�[x7Q�0�6�O�ى~��^O��xg^�Ț����u�۹�K�~��$='#�4�����,W�=~�5��6�[�E�EӮˋ7.��c��h���MN!��$
�d�l1�����n����v����ҥ+݉,D���i�ky����Y�s`aHpH�����9��.l�S��W�H�WY嘪:N����ͮ�n�ѹy�W�\��Bx��Ę�v$�3��aC�����G"L����+�W{��-`n⬳<��/�*Ng��v����	2�$��]C���y׳��[��~C<����j�4j��bWI��{��M�c:SONb��o�{��ѹ��]�`�'D2RL@0��>;3kuX#�'7,6���]��f<�?��������B:2�!���{ލ���������ӛ�ӓ��u�TQ���龏���3OפvA����{vWz��N���3�;��	������Kƽw'��gOWch�s5���<��QHS&:f�>��^cK�dw���޶.g�#s{�~��0��&%���r�ќ��X~w�2�A.��g׹)Ѯ�j��9c���J�&�/�B�&T]�<��\u��W��O�Y}N��ú޺���L3���<xn���ZU�O��b	�IH��{;������s-�l�<�ڐ�d�ק�=��GH�,pe�zu�So<�!)2�B�ց��̀M�����N����K�F *Q}����}3���ȽdkE1���!��n��E��d4�LdWS�W["��S�z��������]w;�*����^�����}�$]U��ˣ��']T@�����(nd����F�m����>���{�mw&��oG�<؋Ә�Dd�7+�������:��k�}�[0
-�ZD>���T M�����C3#��7�~��k�>��{�{C��:��36�m�~S�������2#�~���&�@���U��=�֡�<䯧Q|�W}zCc��l�s�!/�}���Wt���c��6b}��1֡离�z��⛄Ђ[ ��]ۻ�`s��~�����{����	
]�5�.��;%
�M���\�B�u���8C���H�3{�[�����S=�}�c΂��ײ}ޟz��Ӯ0����\�^��B��A� ӈ��Gy�z�9���g��}c[�޷�k�/MwS��ߔI���Z��w��#�yN9<*(^���'6 �����P�^».��>�
Y^�?��`���g=�ͻ����·v�?�_IF�X�E���h��@�;ە|�/0!LΦ);�	b^��e��;wb-���r�?����빗�=�{������oҟ׋-�~���u=������9�H����p��P�;y���y��G;;����~3	���&.%lå�,k��ǂ���#�Q��=S��*�����	�E���:L䁜��]>���7m�*����T"���KE�}�������þ�硦1�mj&̾6���l��\�vd3��4�����MHu������	_;�«󫬴YLF�J4��� �,�)4��R�r���d��ذ����t3Pf.4�O^��y>q�t�h��c/3�xmY����lOOwVS�������P�2�ۨ�s[�Yb!�I|f*�l��G���)��j�}Y��x���ƌ�=	N�$���L�c��B�A�=��T����<4����I�#�Tz@��|q�A�KϚ��}T��b
����r�6g���,�b�H$疂��+2��9��]�W@�� ���3�@��ו���l�/os.~i�����7W;�X�&�V�rZ+1�*�Y�(޷eMܦ�7K�����8��T��J]��GR������zg�E��S�^���b�ui �����C�82���!�2�h,]`,�̩i�J2�n�#�tt#�MI��>�x&��X�ʚywυ��lp����ѕ7Sϰ �my�ԁ�Ƴ0�͆�ҧ3,�:�e�@7n;gu\"e���sƘ!T��R����͈�^p�(�֋e�hdŷ^{pc���#��]�a��[�����5P�Uv�r�E�\ko$�f�X�1vrF!���wߧT���ߍ\�j���R!����,M�oz��v�[I�؆���^k�m=�s�3�؟ɲ�˖�Oݔ���w?z��V'�s�w��=��l�G�u��zb�;��o�Wfٸ�� 6	�E�MW9�y�Eƃ�{|13���hDj3��$l�X&8�mZ��c�獬a��`z�
�`]�� �<�׬}~���W��+����W�]m�*9���8Ϯ�[����l���wi�[�:Q��#�6�I�����E�^��2��m�ނ�ǉ�6+�wTck���~\G���X�r'����[�7Q?���xS�e�킆�R5|j��MzG�o�~I)6�F[�sC{�9��)�EWz.��^C��2�r�y��+��.{�%{z��b��Ca��_wj��o�qAf�F���������h~�'L������t�z�.ko�ӑz�w����8P�>�3�d޹�7�E��޼�iн���{�KH�
@�(d�DlNyM�?M�e!j���Wl�<�(i��/���f��_�=�=3|�jNlд\��Vǖ��.�; l,v^kZ��#���l�����zN��|r���7S�Vv���V�}�$��x/;;	��N��φ�p�ڷ�uQu�>�%���̜��+;
�w�fF�>�<n�}@���'������˲l]�������=�$p��k����.GP�
����ؒ��*�������Cy��?w�f�x{�����y����ወ���mw4��4�R2���F$��R���4~׊��]�P�4㇟xEy���<�^��K5�`YTW�ig_��E3�*޿��pP��0�"C@���7�3�	����5Upm^Z�9�^��l���:��@!�]�N��Q`3��]�Nʷ�3��E��a4��A��KX��d�	�x ��^ �Qc��ϸ��j�L{i����&}���qc���<=0�q�Ꮉ�1��m������0!���`ui�:aV��a�o�~я�fvY��r���2u�M���b�5K����l�	�'6��ƔѴ�t�=P�wu��|*E"�-�q�:�"�'g:������wj-)ѹ��9�DR��O̤������-�v +3�ݣ�^:�6��V�>m�r_����?W����kA ����+ꊌ�0�}������7��k/�:=�T�?�_:�U���n�����qBupV�����Q�`�) �nua7�c�4	rwE��\:�(�se���G�Y�4z2�-����1T��TZ�w9� +��=��#�ɴ�R��9���sE��
Ͷ/;B��O�G3��y �M�9��K�!0�d��^�	QVYSwCtV�Z d�d��S=��q.����`��:�ޫ+{��-K��������Y�y��"��I��YD1k��9g�Ry����j]o��y��S8=閼-N|{��r�o�+f��Kq��p�a�k雩���H�Vi1 �C$F�+*3Q�����rG/��|~^1l�ٹ�j����O�ݾ9M�և�'Tb�&�i��3ދ�{��c���7�jg��������L@���$1�i�.<�_R��Od"g�h��U��[?F{c�k�<�V��֘�7I�A&�m+�d����ʘ��@���� tf�M�������-���B0�Wt�s�R�nX�����u}y���$��u2�j�����pk�q�W��}��h��z�)�M��=��<��^�=��}Dj�����Y��^W6fsȣ�d�'36�_�����DI�罺�0�:맺�������ԫd�jR�$�8�6��v����{i����͉�����s�q�&L&�*��.(�}Â�wt��kO�Ѥ`��^���dpc0��z�t�����{厸X�����.���f�Q����*���ɯ^z:��^-�2��_���`@�w�t�M9���f�W��p�q'�,u�Ysv�������V>eˢ/��ϹN��1����gwC<�6`&��~;*�5������~�`Fu��Q���D^��c�W��s�`f]��f��c�<�ǝ�^�[���b���G�3=a�{�a��%��w�H^����̒�{���θ޻�yR k@�p�6�����U���%6��ZҌ4���i��J���9��ڻ
�㦷V�Gҍs.��cof��yo�7�d�,h��{LͼW̺�������F������Q>P:�����4�\�G\c�hEE�R���G0�1��E{�.�1�U
8z�z�9�2�����˰+���(�"J�,�����aﲸ�:{��<b�|"Ǉ T�8���8��`1oUq��Qz�F��or�^EY ݞ�֫��Qse7;pv���&�7L�<83Yy.�\G���Py{5�=������1�� *M�W�n�WtKQ�u6��P�4h{\�
��PX�Fħ�Dq��L�JXݼ���'+y�nWQ�����=1]$�$���3��q6w���b��X��e&i�%�[�{���p�i�ݲ�=��s��cI��ڴ�v�yx1O�t��$n��Ќ�B�G�.YR���.�c�y�p֤b��0K���X&�Ty/m��/2��k
� �s{A��z��1�gKxM��Y�Ɛs�q��y���Ӻ�ؕnxάb̲�e�&�v���v�U�}>w�֘�d�&����(��G�[���0|����Oxr�W"��P�$�������U��4����	�p�?S��Mg��y��Z��r���:n����؋u�N&z���j�,z�I�&��>��k�r�$�ΪO����W� V���$��J�����9�+�=�n	</�iA|��KXC$�R�?$K�ӶBR��G˰�5J���p�pI$�	v8�n��ϐ��lD����j�۸�� *3l��U<�q}�O�0�9���ݮ�o��ʽ�{�GЄ�n
-
O�4c�ɂQ+��\���m������j�`�1|��3�y�G����U�P\��"8}� ���I��\>=3�0�;��8`��d�3f/�"��I��|F�*�2<��!ݪ ��ޚF���}���2�Uʾ�>��:~��t�g��C��j��ƺ��x-�
�}�e��wt"��-6�&��K�Z&�T�Z�B���������Fw��=�L���Bv�$x��ˠ���gOH�����ۺ��լ!�O����n��y9X"�B;�Nnq�(G���6���Fa�l��g���	�t���,��}s}s`��$h�?�I\�=��z�*4������Z�>����g�epb7kE��b:*KR�F�\9Zqq���t�0N��֦p�Nhyt��[��gii[Yo8�!]�S��a>W�V
�M��4E��	e����B�(th�zY�Ղ���s��Y�<�ܼE���aS�I�7��H�,V+��h8z���WF:˜���m*A��OM�J[�U���&mZ	�wf�CM�;ք���4��JK,4)[=��!�.=�V@�o�N(j�:�,j��VO*��	��t���ۭ��KO�p�W�V�:�dد�2�v���	d�x��:V��펯&ضk���GNh29]�;��
m]*��|�QgD�&�Tׯ���5��?K�KVw�Bw�)��Mv\�:�evv_i
Z�'e_R٩�3.�WT<QYX��Hyb����ˢl�?��b����)��d��-jF�u@��I�sX���+1�w�3���g3��q7W�����<g�O��
����s�0;홤ض(N�\����ጁIȧ����eRY2�s����^G���C�bG�Y1_D����l�+7bB���k��Y�+��n�b����D�79f l@��Y��)��mڋb;K/z'5\zL��p��gM[]�d����<��E=�S��tn�g6\<�V���@jز��XgU��.��9�r�˥z��jX<U��g�msT�Kf���	��WK}}��x�z��*ˬ�­W$zM{H8�Tu�.d�P̬�(�q�n��J$�M�5`�\:��$�U���UR�-:��b�VT
���� y�m��v��m���Ye�	��inP��]�)z���Z�f�j5�������$mҽ	��x��I��1�j����]{L�hx��g��Ms���cK��aدW`[Ԑ��Z0�n�Ws�Д�DNp�����%F��l]s���F��]k�b�^n���/Y��p�����ΑCltuqG��q�w�n�V�3�[.5z�[�`����SB6lժM\�P��z�D��Vz1�tpk1�彝R"�`�n�q秺�W�t�R�]�:3`���25�T!f5J�"X�Wf)V2��g] ��z�Hv� j�qGsv,�8ܮM�a���A�-�LGR�c��/!�Gc���͋-3�ȗWkd�%ʞ.ݺD���C�p���\�385��Ρ�=���-�1��v*�X5���m�k�)M�&l]��wH�xw	���+����s7c(�S�S\S�8䗶���.�lYy��.�aCPh���n������祸��]Mz�,����e2 pjͺ;\����qɨ�Qw3$Ip�6���&��gl�X�t���V�<q����қva9�Ɗ�.�/'M�@�<���rn1������X�iCk)����k�����c�Ӹmb8�.�۳�xs����p̝p��ci��j[B�q���<C�CF�J5۷;k��{���8�ܝ���̅�Z��S�Чl��r`
Ď�"�/�Mwe�݁� �-�Mt�K��X@!6�\mg�0�&��� Ac��f�� �a��6�1��E�28�u��=&-,ppe�_n�:Oe˳�XlSZl\@��/;��d��pR:����X-\tzxn��ui3&�i�
��3��%v���5�=B���"�9�nm�����9��u��N�8�mV��ͳ�#0�\[��3�ގ�ke�!�d �]�]4�T[ 2�j9����ys_��үgh�����p��ʥ��,y����_TI�4n���A�L���'��G���ov����+�d��d������`<P
�����8�� ��5��k��]��s���j仱^���	�ͮ��#�"����G�wX��=��P�~~Ο�����zmm���	����>Y;�!0e{���R�wR�dj&�D��(��~�bN�/,֐0��\�p�!��U�*�W;�_��'��@� �?Ρ��4.ʻJ��}z`��}���0��O��<~b�� ^!X��?}d<wۡ�DuwΎ��-��rK�?}�@}�0���v����ĬiR.�#�#��>�/��H�f�p����x��ΐ4���S#��@�����k���H,��y�;˙P�B��齬�u��_q����Ä�gk�"��F�c{*	m�c�|0��M�@R���(��>#�G��/P�����B��8j���� ;����F��:IQ{;t#
 1�<G��!q|8G����g�j�p�œ�b4DF�S���GX�z)��8�_���� �!5������Y��w��a�#��#�h0D}���=F������?2�8|�">o�bC�|��Gי}�gw#��C�����X�4�`����ͯ��!����>]�+�H��ux?|ۍ�����N�?B8�#�~@u�]	�l�0�>�:9mu��v`�PI�	��a2�{b��v�X�����+��g1�qpf�ܗWۢr>���lS�� } �h�X�Ѣ@�%!W{�������~{�Ͼ�p������������!~� ���D��k���#�Ց�ӫ��ж^,9�n<�2�ճ��u�|��uA�HűihR�	N�?��Ty\Bx	�����婎��l`���r~��Rd�!A5�Q���|�M.���󽯥I>'���P����A����;Ic���3�}d|��p�y�z���ެ�;�1�u}�G�oK_r�k���#��B?}�,�����\ܔ��>�DH7��ۜ�8��< C��9+�����W:��Y�|T�����~���y� ��˵kﴌ�D}����'}�,}�`}�!�!�#��eI����!�f)�R��Iw�����g_�~�#���@�r���˾��􄘉$2`�����~�CD ����99}��=�>�~Ӊ�~��>?C�ʘB��#}�@�K�����2 �['� Y��P�����ď�@����Ɏm������c��c��c��|����0�a�T ��C���\���`�]�9t#��LQ;�� 3�x~�H��#�<\d�#�>��Z���q����
�����sܮ���dI?}�����9�g� y}�_wϕ_M@_[��dG�x��g�W����(�$-_�����9M��@W���}`}�,�8~D1�><[Het��1HÒBaI�J9�m�ՠ.�u�q�c�3 6 �eA(��@�� ���ޡ��Y�>��{P??������{�����Xe|���!/Py��ؚtW���U`��Y�j�~�c���ɩ�H�{�yb��pQ���)����?p?}G�O�A?w.����������,!��X�#�}Î�O���}A?|=��:��U�g=�y[�{�]Wk��v��?��ձ�#�=�Ogk�Z� �@hQ�G� p����|~U����Q�#R%/�G�~� 8Gվa$9���NU�mt�P�ݲ|�rLt���󺬺���4��Ŷtƚ����m�ŀ��\��]�*��V�����d��+��e0A��H�"G�G���`�����c���@g�#�h��G|8��H}Zs���A��G�@5L,�þ�䞯���@����}".7B��ɘ��z��n���&jb��g��BH�9���@D}��~g�#�������qw��<�W}<�t�ͳ�|(��:���������'�~Hu��}�ӝ�{�m
 l�	�Q�}��8@��sڧ>�y�\F�fB>=�y��V�}�:@�_C��f�ө�G�*�}�>���0��$�*V�E���.�� X??s�Ǜ��4���g�ok���Sb�D@�UۨY
�`~y�����t��gn����_	�r�*_����Y�$�������{��M�zu3Y5��\x�a���5�f:h�B�G@�f\ۋ4���ڵ�evf�u%l�-�9�D�h~���,��!���\�Ο��讵X�b&�:�v�S#��C�¿p�W���s�������uTw����n	>f1	B��~Ӷ�$}Ć�m^J�M�4F��{�+P��C� u����$ ~�<~�"� <F�+ܪ:=/f|��d��ç����hs���������8�� �4�v�j���=H�eF"!���őDr�ơ��h>n�X����|J�~��~���OI"�\<{`" #*�s9�����-!�u���å�.�Ǟ��D#�?��L?�+�#�	푒|��DxG������t�A�;nsw[��,AR4�HY��2-��B��D"����5�
�Fы����p� Q�Sx6,��+��+(�Vt%�^*+(��-���*�Hz���m���ٳ{t���DṘ�d�6��x)�-������UN�j��BG87�;c=�&ְ�9H&�^�f�E�\Hu�Xs7����{q\]��L[���"��]V3h49��K
Sű�.�� ݡ�%��ue��q]��pnS����)���\V����I��Yt���ۤ���g-p�ٰ%��Ii��2�G8ֵ����ֱ#	]bX��c����q����F�t}�@�=���D�����鏈b!�'�}A�������P�ܿS0�/�4pkI4jF�>?}�{N���A>Ő����r����HU/��� �=ދ����i��:c�q}�^r� ���>��Э�מ<�p#��9���h���/���G�Pj�|�g*���&Ԅ6c��������H�k���vTD}�C���iQ��]����.j�̆ە%���P����ޢ;m�ckJ6����߸@��3���?i�3Dt� ]����Q�����#�����U���ɏoӔR �1g��H�y�g��n��X���+��<��Xn20�����|��&8E���|A-l��1�{?>6(�U���«�����i�y�x�+�
?p�G��t����|FG��H�w�B�83�!�P��0]��t�GH9li���gV;��o�>#�l{�:��y{Y���l�z{ܯ���a�Y�?ZH���_��ӽ�����U�2<~��+����a��(!��.�9k����OˋJ��W��@d�=Ē
 }��J7Di�������V�	1B!o"8�~?Z���W� p�?���-׹��A�������x�?`���	��!q_ď�VՔ��//솟p��0	�|��]�R��?F���){�l}�}��(`��{���Y��@R������na0Sg_�?���|����xo8
u��wR�Z��M��'�@���_j5ݛn��C:Ė�`�P�~c�xS�+V<��Gq������41�'��FFx����)�D}c'W�LP�Dg���>�,�ðw�^�]�N�0ɀ8[qĄ8��-���������1u$� RІ����;���ms�i|��_?�Cրd�\��E��R�#�>�g�Xs>�c�E	��D�w�`ܝ���+h#�=��d��.>ݒ~TǦZ�/;��{�а����1��{{�lx��B�>?9�L�e�=�+��#:�j���.�m�~��G� #����^�yL�wsC5�D�A��'����H��������:���!(��1��{��W����~�8�?^�,�<�.��@��w��i:~���h��������{(�&� }����t#S;^#��>-xC QE�?1�G�ds_xeVdm|G�pb4G�����"���=�+��^���ůj�_�?ߘ�+»���U���D�\��R�3������#@��o0S�r�;�.�d��K�3o6����yY	��yA'��&ƈ��)�,�=�)�dL���ۨ�L�s�p����d�Cu�ʻ>�2N�:".��T�Mw�uAH��p���z�D!�:� |�u���@Y�y��I}�_?�~B�v�X�p���5\ド�F����W�|/g�4d���pCo�m����ɨ�_�����`���]	�4�z,��#'W'SĬP��F#����9e��&��5i̦no�q����+3D|n�w�����rX�"��G�[)Zn�y:�j�[�v�ݎ��JLwŲ��}wښ+�{G����o�j�9��I�D2�$�g�>���G�BUw1�G�̓��u�=��c�*�E�^�f&�0�7������uk�ޔ��_
#5|rw���	"�u�����&D���4�1 (�/�@g�/%��e1���1�x.����9h@�;7�ql��C���3��W���@� R��=#��ʞA�_��-��/<F�v��$�ٙʣ�ե�E#�6�D,��`3���l��
���$�;]�=i/��Ϣ�cO�j����q�>�/H1|7�=?	����R#^==<h`�{�r��N����M�]}Cl���nc5��ߴFx׮�Χ��! @���� �`�ћɘ#�}�G�DPΌP��SO�E6�2�e��AV���y�u��S�}R�b���:�Pk���יB���NA���!�Κ�y�|(3]`�=��H���:��wC�cqn9�0�ִ���xv���qG�ۏff���@~m��o��۾]�E5�~�!�}��Ć�#�M�	��{��?@��?��I8������?xJ������84Z�R�z/����d���H�a�YC�58�����+"�de���e(�%a�سOV��b0}��ޙ�"��{��$�G��0,�=
�I`���;��h}�w*n�r�j�ڣې���}6�k��X������n\o5�{���pM�+ E��=u��	��w�q�ukt�af�x1�`l���|��H".faT;�������E�cD>ε�s�j";�jt�40�؋j/�1p����׻�_J��? `Rd�Q�>B���<�x�tL���DɈ�y�x�Q���fś��'-�^����{Y�o�g�:8�h�昌UW&J˼����Ȳ-�.�=CŞ`���b�d&�. ���2��
��+\�5��φ*�F=��[yULE�1��#��Q ��UJ`�����/�����L�N��T��Nd���c�
����{����q�c�9ŧ��yC�syAjX��̆G�XS>��ή�6�c�ɺkq�8�Qz�nw\W/`:�� ��m^3��q�c>}�وc�W5�Tp�ɤ����<��乭�B&�(��!�͚�go޻���I�j�H�����?x�-<��eU_ވp��ÊsEB:|�����0:C�{<�}km���ĎIݬ('�
R���#Ǹ�syN���r��@=��M;�KV�k��`�G�L�C��@/��w���1���t{��~�ްl#Ҍ�����cǧ�9h�k�s5�}������B#0R��}�3�ҩ��B��$��.��ȭ�Ii2 ��pYz]�@K��$^�#�������v͊�q�Z�����L�cq��9�>��v�Ŧ�8���N�Q�U{@�Zf�]�`�gC��^�8�E&8pt_�r��,O�/Y��uF�@L���J�����5N��&n�`yc�GvЗ4� ��MYs�ײb�A�t�׭���5��B\B�J+1]�HJ�8J��sm)���ۦ�.|{X��{X	�n9�;%,����vVǨe�4�)��ՠ4ֲ�B��j�ݻ���c��"��K�^��f.�˸�W.�ji
�n\��0�1��;I�N�:J���ܛ�Bb x�>"���웡�����(���e=����ێ$L��<:E�=���p.�{���o���'F�Wfk������ͪ?"]��zs��b�}�'�;�8{�/���[���E�A�#�?r�%�{����a��-S���*�d��f8�e���n�M�8�׻��;u�C��30��$��'�4�[:S�'���8#k��K����W&�g��;�ͩ��Ч U�u}|�:��~�����}{3��戦�����G+{0�w��yu����ǘ.J�8T�O$t�@����W�(|��^��� 8�W���[ݸt��"�sb>�0�D����U1�8p�@�#��L���$Bl4Q`An�Dݘ�ī��=C��ap�P�!"0D��?'��~����v�V��D.<,X��ݕ�}��>�G��������Ԅ�E��QE矂�����ه�_v�=n"����A?us�m���3S:�+��������J����Yٷ��*�������g��TD\�n�p@�ѐ������kf��߼8~s�ϧ�����r��ۭ��O��Y>���y*�5��̈́V `�G6�ß]��7m��\�<�j�6�����5�b��qG7*���&;7����{G�2���%k%s����l#H0�kr���0{&[��� 2����ӡl�$/]�;d7������M�[���)*�~MW���T��;��{����A&��"��+.��E@�)}�-�;�K�;�il�v��S����o�ֻͲ�VY��j�F	��Ӽ�L�Ѱ0�Q&X��Z��+���[�jAr�o:�uwuc<&���f�Z��[�)}�A��?gw^U�m�!���n>��#SKx��A��C�"
N!v�޾���%�Nܬ~�z{J���аs��9W����,H��펪�q�W�3�I�#U�@7t}.`�[�L0��R��;{�螄��j}^����N�2��1��5Xbu�W[S��3U��v'}����9���Z������u���t�X���FlA.�vw8�����v�z��\"���|ը8���Q��yB`
���a����G��k<A�s���`�$�u�"�R�~/�'�����"Pϛ��R!�9G�C0^D�//�|'���x�r�ڱ�]�?%`����Ÿc����]��X2R+��VZ�\9+���$�"# D��76Y�Q�'W3U���a�'�O� O�G_VH�Q�����3�+7�L�UpV�{�K�2l��n"�ш&UK�Uڠ1��G�T�n��}N����e�Y�o�}�"ۺ�c�=�z�ql��Y�]��p[ɡ����n���m4�j8�Q���F}����<́�6�O��
�rìD���\�%g�b<���[�!��4�H��b����^,qIezg{�n�@�&��o�fu���]�ɉ�<L�`��#�k.�mz�}Ի �oo{�m�!RO���?y:��>�������R>�Gt�*&��!���tT�����{:�uׇ�q�ϻ�����7�eݖ�~Ŏx�/��S{��W��X)�<��|��9(R������H��H�|vfz �K��<�Nݎ�>���\�:����se�}�K���W��
��uS;�FE�oU�sO/ݑ÷a{^�Go���6�'��UY�gJݼ��j��
��@�L ����2v�������ȃ�r8��;[gC��ÛT~|�_O���I>��]��ͯY�sZ�=��r��R��|�u�Br�j��vd/4F�$eB̪c{K}�+{�=�Y�N���遄���U��	;���߷�����-��JH~@���n������G�'��I:N����I'I����Q'/�����w�k����:w3�{����N�$��/�gN��$�t�'IܒwwN�O�	�O���I�;��$��$���������?c��_���>��o���|����߻�>ӿ?����I�ww����������I:N�����I'I���x����d�'�w�?�߿�t�N������?��z��??2X}g���K�I:N��Iӻ����:wN�$��B~���:I'I��O��>�������O�i�t�t��޾��������w�<_��7��~��I�wwz�$������~3��N����}�$�����?����I�ww__�{M�$�'ww�k�����Oh��?��>�f=Y���$�'wq>�����~�?���I:N���?0��|}����_i�I$�;�����I:N����K�`_��c�ٯ��,ts��\�| �>����'�|�-����� ���'������� ���G������~�������)���4����8(�� H ��1&�{�}|�{L�Ҥ)�*DzA%.e2�*Ӝ�L�R���D	)�n۷=1zh�xF{b.�1��m�HQ�i�Ț��F�u�[4��i�T����AcEJ)T%"6�}t}>�tt�QT
           8�=�Au��[j           !�
�  �^IB��    �W��=4S�`Z[�u֦����J��wplQ������J�����mӶ��=��<=��e�����y� 7������jm�v_g�v��o�4���r��H�} �*�ƅ� �!"�R*�=�� ��W%��öV�وNػU xv
Ѧ�����4Z�����PW��i�_5|.P�zn����>�r�جk���❮ڻ���^���͟t;�^�'q�x�{-��$�Ҁ}kF��M��6�ͧ�ך��R�Cji$��I�wB٬����Y)ڼ���ѡR֗�i�K�X=��N݅�M�;k��kl'���|=zgos���������[l���Z��;��}���{�v�Oc$����w�����а)D�$��O��P  ;��z�ҽt��{�����;�+�J�ƣ@th:������]l��uZ+��_N��g}����r-o���gLթCG�.TZ��=�������/w4��Ǽ�\�f����n�	*���Q"W�=٩����XZ�9:tzև���!C����uI�,`e{EԸ.�{�����zu�m����c�iנwT��=}�|7��{�CVQ��2Ul�ZRG׀  <�Z|�۪��Ӹ����$�KgM��^�J��vu:�ݨ82I}���5��Y�Z�����7@*�������k]�v�P����f�������ժ���z�{��Jӻ�u������ww{{k�M�������ͷ�}�t�$�wt�2>��Y�u��R����;�mN����N�o���0��T�]�X�@�@ ���}ءUW�<[IS���[��3�k��Xx/j�`�ɱV�O�����r�]�w1R�gs�H`w_}����I�5Tq;9'(4W�����*�
 �Cg�h9��� (�d��](�cX�S��5�|�rk�n�l1�QTHt��=4/m���
  Z}��}@>����x���l�jB)@�B���  ���7X]��g�:4*��s�
�݊��oh9��f��݃@���A�uqYN��PHo�s����_y��˰����z^��Sw;5�_�S����i�Y�)�Bb�T � ��CJU    ���*�&?T�&��@��P � "���Ȫ��Q4�0d�Jz��S&)�G��M?T�N�����H���C�J��|���ʊ����۩E��%*X���L�2� �|��/�C��8��x}����;��������p wq�wwwq����wq�Ӑ��wq����wq��8�������}������~iK�_����9w\�(�!
n�m�L8b�����&�]���9*Aӷ����W�]2�o*���a�Y�T���ySGvI��fҊKWw��X�E���N��3��m�Bل�7i�5�"YWi��-O�(#�T���%K9��R��\2k��m֦P�#��(LU����J��Z�M` �l�6�x��D��ѰhV�Z�oi�b���dE	���\�k�Ī�>쥓�k\�*t��|	l�d 鉹����*	:���'nur(�fL�-� ����'��&Dr(9��]v��3��Tl��[��w]�{���S	s
C[Ǚ���H�j���
{k��b[�DK�Ɔڕwbź����nZ��E��`(�p�3M��I"�1�ɋj�wX]���T�1�v�P�u��V}��0������7�M1TP�f%Ff����F�d�҅F��nJ3iܧp�N������Ƴq]���lX��k�4���� DR�MnB�t&jx�!����J�2�mc���Աϯ��-c�.����;���#d�?+Fޚ��R�7o@;�+S�l�JՊ����n#Z�}�+`�\f�iS���GPu�c4Z�C�L�M�W�C��	�����S?d�O5��x"��ubN�W	�M&v�[�,@
(U�EM�)An�ӗ�K���,F޲q��KsY���%b�ؽWvİ����HBq^�)�6E3�Fh٘Ee6��+ P��x��u�Ҭ3�����)��[\(�E��v%#z�R|�mio^F#�4kcr��x�)p^l"�=�n���a��	V��[����&�Y�ͫK��̽��;E�z�5� Yw�QT�-�������b��̢�1�:��%K9�[	Be4�Cj�k/!ͣchh3#cͭO�OX����M�C�c�gW��gN�53*��X��4��3$X�T�	��6��.X �G3܃P��������˩?d:U�o��bT�P�v���4��ʺ��X��TzAZ�sp �m��4�R�ib�r��ǃ,۬�U���b��ȱ%k�Šf#!���4CuUiNo3������<T�Ǹ�����t���p�K�utP�VE�^n�(Z���_|��>�0�"an6��?�h���C�m|(5$BU�� ��{9T?%�h�_�Φػ�#�A�˺�CNVKZ��Ȳ=bֲ`$f�^� �d�Ė�n"�Ѱ�e�QZ��2M�1]�M�	U2cOM6�8K؅�2dv���B݇I��sr7��M���s�����&�Y�;6�;u3/n�
'f�hn=[	V7*퍽��2�	�P�c-Z�dw������w[0�A�%(Ш�mj���X�ЌQgH*�e�d�NPyZaڛ&)W��51�*�����Z�%����]E��YL<Hm#.�*G3/"v7ib��hh��a�-�[f��tY��H���F4�Zۄ*x�q]\׺�Cu�i�.ր��8?aW��R[R��L ]���7���4%����'�.������3�Y�͋���.�m�Fh����c�젩���o	�@�aXm���1��s�e6���8�\��<z�ā�*F�la�r`R^�U+i�:u��M�8�cX�{Z�ƪ�r�Ҫ�-�p��.��%��%ꌲ͇�]^����C�8M��Y��C���[4ެ�Aُ4�{Q�E��Ҷu(�	�]6�����'y�p�_&X���da�����y��r� :�(�Б���Կ������'KspV�-���POe;�*��zơ��0���ݭ��HT���_�������e^�͌=�����H�ww#;�0��a��$2�Q�.;�*ڴ�0���ܰm�ݼCkh�)أ1U�4U�pJ2Om��i%ӕ	Ö�9�4�ӳj��xqB�h3Ez쇪�~�(~к~��8�}���ܾ�R\�A��F���[ͩ�Ů1��_K�{��h��K
�M�P��j��]���%���P`8�0۽��B���7���?D|-!�q��><
q�8�����}�)�׎=N�׃�q�8���}������M�o�m)bJ���<�]4)o�spLg3qmo�x��N��-^�k$�N���}D{�����ۣ�|�D�x�x� *�"��l��n�ڕ�ᷟ���l�&�O^�����0��1�\xr���f�&��hAm���6#��.��tuk5`:PZ����$5jL�Jʲ���ڽ�w����zL��*��9��K��rSI��:E�tm;e��ߗ�<��O����
��d��J���6{���~��?W�&��$���6�F��ʻ�e�9dh!eR�}T�5A������	L�a]�	�.�[O <��z�1Om�X�dA�D����{s ���`f����ga�z��2;!�wx`gm-�n4E�y%������Vec{��B��u|�5��Y#f�������V8c�چ:v�2%a;����B#��_a>s��=�K5nIF��GX1_�p�����t@���P�*n��ݴK[�d׀[�n��Be���F�D�1[4����5ZZ�;oO�u�o��>y��~?X�O�ts�x�7S�㏂
����^�׃ǻ�?X��'z��QUO�
(%� �ѓ*&l�����m)5�6��B��L��x��m��7cq�����Jb��9qg��*�Q#��d}D�j�}5}w��H���.6�X.�����n�N�;I�����n�,h�n�D�W�hh*o,�8�=��֯]�k�en�PS]h����A�Y�P�W(-�7aH�q�E:ɶE��O0,.���c�$Iwt�&����KR�D����I���#�`�{*e�cL4��J�Lʅe� `��r�	����К+n�.���US��`t���.�9k,e5�e6���&LT�OFM!�'j���6�\l�����њE��0m�gki�b����Gx��8�Dٍ�,�o+2�XqT�/j?ct��T��퐦q�R�D�� 汚e��պl����l諈�p2�Z�T�C�oe��4�z�!6�PT۬�C�ܵF�5�6�l!]�ԛf�D�z����ђޅiT�Ơ�����B��c��n,�����A����{��ffj)Ckf���A���Úk�&dx���&1���N�Řbq�[E��ݫF�f��B�3�f���!b�l��1GU�֎O�T9D����a�f=�Z����h����V�3�Y�0D�EN��ﮋf�r̐F��*~�L��ו4�3���Ʋ^^��x�8�q�3ߘb�G���H�D3����m^��Q��f�,�s��m�	�׻yy�X9Ym�1ItG��W��'q�ǉ\&�4:�W���U`���6���w�>�z�g�������'}x7��S��'{��}x<N2q���;�x�����ﾶ�#�?"��F��O~חr�KN���&��!�r2�V���=+��L�{�VP̩�!��m��D�s0�n`��\ˤէR���	Q�{�{��U��0K����5f�Vp�y�$f�#Fn;bhH������t����uF�����ˠE̻S�ӱ|ꂢ��s2�FB���Aӣ��̬"%���٩$��ݭ@�gpm���f�j9P�W�[
��sRkoe��UU
��W�^f�VM��s5��a�(��x�=ڷI㲮����Jh֢ì)Mr��Enᡪ�Z� =nXӦU^c�^��)�ԍ���Y9.�-��b����[���j�m7�&�ͬ�M�ٱ��nMەy��H��U�'����i��5n ژ��Q�4늲����B��������6�t�%8�zp![�lX�ؽ2����bd��wṃ�Ee��Ż��D�u�ܒ��v��s"���Z*��ʊ��F̣l#Z�ufƢ6G6�����(d�z̒�XP���p��9�Rf����\32�YUjS��X;��'�u��¬Dn�7+5��s#�s]7C%-��@���V�$A��/]�˫��X�F�צ�]�m���Ȣa�4$v�k�a�6���pYZ�賄j����f�^�Ưn��ME[gZ92#���3@�yP�*R�A�����
��	n�x#x��\��������ߟo}{�¯"</p����:H��Fp�`��z=�ܫ�� <��	¨�"N"�"�"�!�N�������fnM�����MT�V��LJ
D��I�>%�K�xw5l�RD�ķ�Ȟ��j�$Ȗ��ո�`ȭd/��)���F��wj1���Ɠ̔��v�d�T��e����?A_ab.�z�h��5NYh
���Yw5j�S�û2�g�H4�Ae�ce[i��f-o6��m�j
	�ڵe��Q���(n��1-յ�Y���9���t�ZGm2.j�Z�@ǲ�ww����ɂBB䧀8,�x�[OM�)J)����WY�M�:����5�R�{[H'B���ݪ�>�"�F���`�$M�ꚭ��K�Ƃ�w�'<g�{��^QTD?~����n�GmC�N.��	����7X���Ә�ɍ@K�#�G�?i|~ ��*�����9BP�~Ϟ|�y>��*�������'p�w��p�
�x���J|�}�rQ�����E8�5+�f�2��[hk���b6�ښ�5B�䂢��٩��V�Њ���:)n:��v��Ct�
�+��B��{)}ph4uRss�<���G�Q�בl�ej����%ֶ�ꗺ���2����)Z�·�rk�c%�1�ٺ{L�aC\vu�/,{Djl��l�!�f0m�7V�Rz�U�E<�PE���R�ܬ�k�WJc?�Vދ�����A������3r�h{kZ[�q��(`(~�ɹ�M��Pطk��j9/o��4�viW��asE�Z+��^�_)��ڨ՚䧶��ĩ��S��ֲ0,�On�d�̤)�R҄���Y�en�r�
4��"�n�u�Xue�Bf���ED���1+�H0��"-#ZE'7��"��uN����J��t��׭Ѳr2�7g0?�ٌ�ڳ\���.n�+^�9-���R����q��$�+�J�v������^��jꈓ7U+�-AX�"��*����~�����݊-O��R���H���
�L��Dn��زₜT��wGZ"��J��F�R��1GN���tR�Y�e�s��+��v={q\��?��7�X���&�*q�� ̺���S&��sEnmA�[ۢ2��6�6��l%�"q�tm��c��J��X��eE�Ǳ��&���Kh�c�Ḿ��`<��"T-��lmE�+y��EJ� Ŭ굓�yi����z� ���u�T],[��ő����c�@;�����UV
��&U�E���Cpc�R���c�4�R�� ���I��[��c�Z���+F��Ԛ�V�vZLcn��8�x���W��J�m�]��w�S���0KXm՘�B]�9yn�a?ee��ЯW�6ȫ%��0䂶0ejZ.-vw%��wE�lR���fu0o6�w�I���]�wa��Y��V�/J���RT�e�4�u�۟D�*側֭@��2�Ԓ�Ż��qȨ��l%&a;��ȫ��wvR����&��2��@L-Hbpf�.i����;d����պ�.N�n�;[�k��P!Е�m�T�l��b�7JSj�0e�,h�yq�k.�p:N� *+����m�&�^��4�Fh	bz)�5j�]�Լگ���U��fňX�+��"�^�jѮ�5orf~����
�H��Ɍ�Y��B]�a�)��9h��A�;Kj�n�v:�bn�uy@Ae�P��EnX䩎ٻ���^��b�%N�ٲ��2����_k�����^}(��'Œ��;,<1nYn���Q�k�vDe1��u&�ٽY+68��5;k!תV;�w鬏U���iR���n�*ڸփ�f��d8|t�̭9N���MI�%\j��5���S�j��kU �7Uzv�ڨ�p%�7U��)�M�q�n.wm뺧e��+0����+u��e�!d<6
��e2V�W��������od�p�:�I�U��Q��Sˏ*襗���iSă��[���و�Ĥ�L�l�֍�{�J��^�w����l�U*u(�v������J:q����B0(N���mw�ul ����8�n����WHMnr���Ǯ�M���=��k/(bH�0���hq71rf6�Yndv-�ۨX�ؼM5OI��[���ܲ��*
�d��Q���+D׷��&��[1�(fR�1U�{f���ʒ���R�5��(�Yvݱv��<���l�[��n�&�%
2��,�Z�R���]�eG��N�,Q{F�Y��A���!Q�AD��  �   �R�IR@   U@     I5)�T U@  Y�Sm���mͲ�q&֖��l      L��*n��.�n��pq�x��e�gA����o4c�������p�{k8V��ֆՆ��V7n�a8��L]�Fn��8e�$Z�s�l̼	g>���5N��w�}��^< ��|�M���\�ZЭ����cko�@��v�o�k�#��4�d{]������ރp8����j�r�F5d,��QŠ����Q[��M��BS�7Q�Ei�
���3?#7�A؆����ZZv�YÂ�Ζժs���c�e6��:�+
����U���n·*+�I�up����=�x��)
��D�C7xk�v����WD��[��C�m�Fe
�ɒ��T�Fv�h�V�8�:-=�;2���f�p���,s���B��m�`�a-bl�����4p��{�娬VmnVGMA�cSb�@<�j#��ǁãB��^�y����Kø#Z��c�r��l`,ǳ�4��#:#��v^< n!��8ʅ
.�l�[�Y׼�mab��꺁��2�M�_ǳ��Qa�U�F���s��|E�ܻ��H��ݼ{�:���U����I���b�l���Zp�ɜFX�^ ���8_<�"���'G��n\C�r�Xp��4��7��Z9�f���kN��%��Z�����Ĭ�0+��%af���м�&��'M"S�y�kl䢬��娰ҷW#]�����5x��s�2j�/g<�ᇨu�6����@{�Hѳ[�k�����J��S���"�����:�eUe#:�]vHBF�J=K-ޫ��e>�A�D:xtWݠ�۔H�K���_&�Gn��:�"ͱT�oX뮊�������'	�g:��zs�t;e����5�Y����DȕLE1aҵ��UՁw=���t��� O
�7L���)Ju�B����F��ۭ��u����&͌9�%��$���u��0�2�k�ޮ��Cem]��ǉm�gg�fުdtӒ� U.n͡�\Ɋ��^l���2�-�N�������{Vt�Z�=0;OdR��1�w�^�j��6l�kb�sU����*i�˖��'	ܹ�'�I9�3S2=��%�v�fMǎ�
p��R�:w���5Ǆ�)7|�-�q]�f��J�
�^W�Why@7ǐ�Œ��\���s�iǯyU��E��S��齹�jk��/].�N�Ǌ;]�s�r�㔢��-��v�ÛP�*&��u�����qچ�BC�NT�u�|��x�+EQ�%K
;�����T���'��ٻ�I7/$�q�{U�)k;��R���=�]��v<�]�rS�ؽ1�{mr]:��ӂp��t�!c5`嫦�i\�=�D�"��Q��:���d��u�+��	�<ݧ���ub_;=��9<���<z�ʦ���T���'EnG��D1J�r��N��Y�Y���X�bg�œ���N�/�N�������2n�f��@lwF�"�J��q�R�|���y�7LV��DTS�5KM����mЙ�����(��ŴCuYז��7�&���6��ېgi��K��.շ�����k�@�qd�����%���bn_*]�U�9�+�+(����n@h[mg�ur���s^	)R����{�U&���X,d9�fL�׵������M�9�v�ǯZ���`�7�1�ecӏqh��&�n�tr^��nl�v~j�FUS:���W6K,kcB7����V���~��9���^1l�`���f�o��A�{��b����~��`��B�'V�y�R��+�W�귄?Xj^L�W���н��.ueL�깤�$��/j�=���f]�A�e�]N�k��]�qO��o�Nt3M��:����0f�\�;�Yb1���;.Ys`���[M�ӲnŻ�Օ�VfY��SL�"��>��
���J"�\�O��g:�=�\����C�
=q1���)6rSQ�;43�+{�����k:��t��h� ��cCuc�H��9���,Jg�4ƫ�Ջ�>G�UuVY��V�	�B����3�r=��7�9y��**y�˝�|�l�R݆�'+k	�*)É���Ͳ2��x�F�)��;cц���N�)7-���w==�-#�K] Ԩ��8��^@u��"�*uء�"�'o.ӳX�:�L���;���_.��1Y+]XRu"��INIT�%�ȪČ�-]fk�yb��Z�yiW�B61X;Gv��5��_0�<+v������7"v��I;C�W� ��V�̰�ͽ"�P&ƚ:AF�T� �M����%a�}w��[�g�b��ǚ(*�m�:�����멃�7����)����	�_�w����A��EX���>ޣ��F���7g*��9>����;v�)װr:�8�\���\�����N��{S���r����	�>=W��o����a�<�C�J�;��ߜl6����uD���!fܖ�P����H��Em�	*II��
�fա/���۬��̈��Хc6/iJ�XP�
�q�;��=�M] �[��d<��W�U!�����{�o�L�����YͧE�i#���Yr��Bm�#�L6>����N�hȦг��
�T°L'�ʑܥ��W�"����3Hu��5W�AS4۬����(B�ȢiA��n��UQ
��*�������y�/��뢩2x�RN9�U�$Yu�E�T���|��>ii�mܗ�>r���&����!GM��p��![�2ʔ��+*U|���R`B_��2�&#\�!'ɊZ[�W0�D���)v;B�9��i2Ra�/�;j�%���J�V�F"b(�堹�P��}�9JA
[�eB�@�Ql��Y4*��76�$��%f��4�P�׆Qa���>~�/��J�J�c-�V�4Ξo&�!��UXD�i�9�T��HjF� itqM�I�J8����j	UF�D:`�(�	�m݂E��-󐢁%St�b5S�t�28䜫�����!�5e8c�ab$eP(�L��m� q�#��)�!��UB�"�WM�V��!��DP��,u�P�r$�H��/���<&)�s6�f�F����<��p�r���D�B��D�=W�֍�����I*�%Ȝm(��5o�)�4�5�Zf�|�Ĕ�_(�q�j�1kd�R1���U��e:P���T\G)%gW�M ��q$a2]m�&���h[z�l�+w���A��_�l�4iko�2�\I��>/�l���ڠ¦�XR4�N"$����eml�ՒJ���7��I-��elp�f���,���3tmM�Mu��D���o����1�JҺ��a��D����7V(�h��&h{'�F���#�������s� ڑ�҄3$)<:�YM�xL�lY)m�5e���|<��:�Ԑ��[L�X\ˍ��Ϟ��>���>��ѩqtIRL~$�̲���X�5�o�"����[i
;Sm�Ժ�Gi�m%�g4�6� f9����.�k��h������ R)�l֤�R��v��e��K*-6��b�b>k�z˴5�}���5�����l�;k�Z��Vkmq��:k
\���T�2�V��qMi[b�-fn�i[3n���fx�ɲ��j�i:R��4,�K{6�I	�-�:��g,�v�q];��zȶf�2�fM։��5�t,!m�79�y��$�M��5ԭ�7����������R�c�c�bd�$�f��d6Փ��y�O:����m���7��KۢuF�1���<-�i-�-������%�����&�ĵ\B�%�+�O���捜�p����Lb��,֚��;E�6�e��V��l˰\,$�I4�պͶ�bc;72n���f.�Y�����D��5eХ��,f�f�YQ�]%��T�Q�Y-�4n�-ý��Z޾$��[���m#)�������'N���
��hv"��O�A�H�����/>2�FSX�Mr�B�=j���\M%�(���8��Ĳ#[%��Nw���؉�u�U��6Vڷ"l��:�U+�:��,���lP�,�H�֒L���K\�Fg�ltk�M߭��3������Y�GM6j���7[�����,�<�;6Km�/6,�$5�1+�4�$[ql��R�Q�K��I���:Y\���$��=��V�Q즲]d��)6��������
����^��g�|/�i�FfĄW����>xDo��n5�w�b�BE<qI�n����R�I"�ee�LcX]]����)�ٟi������Μ�K�U$5��)9Y����I���dӳ�0iq�&�����R�|�3����m�)�M�s��u6355�Wn�[��m#�#vñ��G.K�$��mmYs-�HƑ�f�#�}�����d��kp�m���b�գ���%Գ�u�X\�un&��oMaj���M�����QH[n-�+��p��Xg/8v���sak'�󘎳�n��Z�9s!�gh�Wn��WL[��B0�fva.a�tl����[�=�g����<4kT��lEt)
;�J�yVH�5�ԦK,����[�j��֕�Q,ډ
��Ɩ1el[uGFK:��h�s�]�5�CDKbȩ�a��d�E�:Z���h�	6��"HM���T$�,�b��Z�a�y��3F���ˤ�����+LY	�7i$v�$�]iu���%�J�N�c[��۠n���IYmк��Ҷ57i��/]u�+IkZ6e�5z��	WVh�Y%l)����me�Z�)m3.-�K.X�v����W]4j/%[)���%���semIԳ�&vr�15����,!h�ٱfta�q.��[pȩ)mɵf�iZ1,e��&T�p���lr�dJ=t�s����sc�Զ�s+������8�]�,�Q#u���7l�KulҰӛrb����Ɔ6��%�M4�`����F������hN��2�K���m�����*h�.���ƒ�[Ηm&٭��ҩ���$^��%�5��*6��K\WB�T�ŊĲ��-h�RH�1���6�uɥ�ͷ����ɵ�..�����=nn/;M�λf�Ѧr٨��4�A�S���'WL�,۵тjV�
��ɭ��bR�L���&��Fj���Eыc�KlmGL�Z�䅔ȕ2K��'9f�;7�k#m.e�s%뭅w9�/%�WF5�l��+\�����m=4����u�gi[k#��D�G�"��m��R6[q�X��Ź���f7Xk��I[����,�\ēh�ӖۇM��*                                                              .d|#��6��a{K{<����3�v�Ҟgk�k�}���\A��%�N�,��*<դw�cCkE��S7v\&�\Z��ǛP�[�=yW�Ы��m�y������4�.�d1V���1dԺ�����K4�����3S#�yJ���X���Z���L�:W$9��T9�V cd�;�aׂ����������]�LT�6k�e3��Z_E/E,b�i�$j���{�T"����'w����s"������Q���"�n�}|nZ�e�˽L���)Y]�wr��ѯ1���z���r�Sk�eμ�k�@�Y��uG��.���Y*"��5��%E���6���Z����if2�mn�[Y�[-��G���@<�ϫ/t������@��V�gU��s"U�u�[T��m�B��+���Ɠ	�m�֘�0u��W����w\�B�ǰr���]�	O����M2Q��`�k*��;C����A\�.n�x�Ks�Z��,�M������]��I��U(�on)�\.�2����p���u}[�W`��q����3bdkGsnP�1δ�[��k�2�*V3���V���*ut�!�&���k�ȭ&���]顃bƖ	�{�r��p}kw/K�X���S2S�*q����[���bx�M�9e'j�������宲�N�;b�U<�E��e�x)�eb�
��`�8*�U�$QyD�_���N��M���,=2<ǟ�ᝤHs������[��·�� n�[�7�%�f�����za$�F�U]v���h�w��%0[V0��d���u�oF5�XE��%u��=�EU4~M���-�A6���D&��ճ.M���#����K@��+�T�Lo>�e33�����ݚ@ӻn�Q�-+7��Zr<쮅>�b`Ѫ����M��w�C�l��z��%��y�>y�{������� ����wwq���'׻�8��q���������x����x;��q��q���;�׀���<N"q�{���	gw{�!��wW����q�$=�#�q���wǸ�����pD�<�;���q���
�ǁ~y�!�ǈ��q^�=�D?~�ߓ�'w?�x>���=N��C�Ǐ�wd�"��N<��?<~C��W��8�^�_>E>����={�l*uL�PU��^?=��z�<�P�w�N=��p|{���w�8�;���?<W�׀>�����{��<��'����^�#�#��q$E���N���t�2��ח��!���w^�D����v�h��;��^<D�r���}N�����/='�����{=ݐ'��
pzת׀������P����;53�G��_���"q߼�q�/x�d�*)¨z�q3���r��� d?'}xt��ya�}O��C�E8��R���`x�y�o�<{������@��O�N7���x���+�={��x�B�G%W�<g�Ű��H���ߞ+�޼��x��ߜ���?N<{�랒�����;�L�G�r�|N���dNϩ�'{����w����tx*~�
"~N(�ӂ=��t���~�O�系ǎ��:<z�S��}����_�>ܝ�,�I�z��'wG�{!��C��D��/��^�<����: vC����w�x���@����ǂ"���z���m ,�|N����*v{��:������z����u@����w���d>'�x��wD��?<q���4�d�
W��G�'ܹ�{��w������ܽ��N�'/pD�"[^�P�N=�����ӯ��;��q��L�w����ǨN�'S���d���{��@����r�{gW��^ �����)�PP��=��8�����y�w�P��{�È�!�������;׫�P����wĢ�ݾN"��P�S�������<O�wz���|x��;� ?'W����6޼�������> }�
�������wq���x�>������wz���jw�����㈇O'P;<z�~x�;����/w~N���8���q��^��������Ï^��t@'���=����P��q���g��;��)�w׈�}Cǎ>'�C��?y8�^�x��������޽�SV�����'}x���w���N��v��qR=��;!�㏯���Ǿ'Eӻ�z�{� ��9{��������w�T=z'�gx+�l��Q���x��㼐�=����� ? ~xS���!�p�)����</)ē�u{��׻����uN�f<���; �<J�_'��={�x<���� �u{�!����9||{!��s��N�̇C<ux���2N�<�^+��;��q��������� ��P����8>y �C�y>'W��{�>'~B���[����uC#����-����޽����C�'w��ǯ}N;����;׃Ǻ>�~�q��ߐ�|�8���<}{�x>��?P�'tx���;꥓�T����NP���}NS���׻׾*�;����^
��C��l�g�Xw��g�D��s����z�N��l��z�z������ߥ�!�R�S��Xy��T;����|�~Ol�|�}OP��}l�x��>�~z=���<x������g��=�����<���^�>!�5gǷ�N��ԏq������d"!񈮞y�9�˩��7�����}п�w�u�9|z�(QN���}yO�_����߼�킔N�N�wǊ�ߨ_fH���ϰ���O�~z��{��wz�M���wvO�@����J����<�;������? 9�r0:՟���m~�_i��M�"��ÏO�Iq�������E��gG��z����|�����?P/������t￡�/ߓ�?|�+ܱ����=ߨ|{ת��8�8�����t��X/� �'/班R���p(�J#TJ�����+e�:�����~�	8><�S�_��v�^�q��?������a�����'��������(x��ς];Ƽw�x�xC�ꞿ=�N��{>�ƠF�W�>=����>X��|���w�������|��	�����p�����G���,���W�$ q�����Er���{��@�F|�<@�_�98���E@��UN����=�'������'}Cǽ{����8��z�C�>IP������ +�~�b�*w�<y�M@��G5ƞ���٨6�耔�N���{;�>�z�����D����@���
|-��g��@h��?^#C�Z���E�N��yO_��t��DR�Z�$�G��􄹄/���z�N��xi��*��*=�������{��?	�o7~C!�~@�����yuN2�?!�h{�ϐ<�?=�,=G����?zN<~�������:��4:���o:I��>| |�;�!���{*����><g��������O9�q�S��{�C��^:5����/������;��;�'S��q���|z!S����D�����ߟ��֕����8��|{���玉����z W�����/��8���#�������� ~x3��_S���Я}x���d;�wD��^��~{�hu��|x���S��iߞ/�i������G�~Bz�/9�~=֯�A�*aa���kUь5ˈ���ۂ�������}}�����}�������]H_����(,Zw)Ε�Hsk;3@r�λ �T��)V��tf�MȆ`QsGfVV-���xu	E
�ᬕ���x-�K���r3�Ch�0(:���:�6v��¹ɚ�R��ڡ��;�:�Y��˗�gu*��׍$<��bAD��;��ܺ��MT� �Uz6<]���J}��U��sz5c�!n�%R�� ;M�d�������0>k�����^�4��'�'����q��ζ��h�Z��d�v�娆<���B��d��K.�F�}���uT�x��n�w@�!���e���[N��cr.��,=E��=|v��b�Ź���!�R�Kw�[e���.��8�;��'p��p ��/����=�~�76�p��h��6�R�nƬ:���َ��������~���?~��wT����=�8�����﷎"Hwx�� ��C��>|�N�^�<�/��<C�S�"vN���<g���㊜~�w�{��z�߇���=N�D���u{��o��{�{����M���ʈ��#��輼�*����)��;����{��=�DQUUQUE�t������xT�''��Ay���/)����?ߔg��(�=�*��+�i��b"�9+UG�H�ӞG���'<�<�"�d:B(����{ʼ/<��Ĝ���?7�d^|b��}�9�痕�DPW�Q�^Nk_��9y["��<���t��@A�%Pyc8y�"���n�üB*��DFsʏ"�ӅW�����}C4t�'{�y���~ ��$�����N=z�^UDM	Ȫ��8�򨹈��1#�>��y�ϛ
�¦��
"

��y����DDE�UFB ���<H����_���D�V
��~�y��/E=��{��!����{w���U^t�<���(����˓�DD���"/$�n�a��]�O�kq��"�zhH��d��>}��g�����}�=��N��<��Я)?R��O��EE{��aE�m{����yTydK�FN'"�*��B(�@�<'B���8��x���NY	�E�p�H�_�=�H*}H�g|x��}g	F""�R#��DC�;�ܩ���b=���a|	0��v{˭��Q�f�*0!�>Kg�N��甫���F"�N�<��_�Qz�x���n�"�殓��s'߿�i��М�B+G��ɋ��*�z؏�EB��c>yj�oO�΄Dy^���,|����F�w�6�����d�]BP�i�m�i!��l����~?�tę�&�w��q���
�d���d�x���+�W���*XC{��7��2��AT�����us���gH)�j,��ξ�m�����27�]��"�g�g�c�*��#������J$�&֙�Ma+�~~�]n���P���"���G5(�mQ������UC'֧�y |��"�JW���#a���;}�����r�C1�JT�E� ���Mw�S�7o�̐��h��_!D��Sب�l�?  F��\�!��p�|�<����U E�$/k2|��DS?Fo�%cÖ�
ln�����'�����\,>@�x!�������m?cd�lѐ._n�
(�RQ��<��·�9D�b�� �޾����	���H���^�6H$R\B�%"�}B�0VD~�v'#?�y�l@O��>��O�4��"�کz�&eYU�h�I!��;�:�4��4��!x��ʊ�XK�a#�������2I�$����(BA9�	vő�X$a�S�آ���]$���4�,�lk;�Y�.Kx�s�R:e�U�"�wA�q�t��6�R�G-��K=��Jw�\i����^��Lқ��}8ܛ=̫�*�a�#�wq�M�q[��s�#wN�O���fH�oQ���I1,��vX�r̛��d��=�n��ڍ��&��1��,k�Q���6��7F�ٵ�Դ��?����1���NoN�Ѯ�v��Y��7C7m�����������T�T�!��4	�}>����l>%;"~R	$*��#᭻��@��!-����hݶH��7ϔ*ֿ���ӆ	�E�G��5H��k���.5|h}�|��mk��"�O�=֟��-E����aC�Z�h�~/,/Z���"?e+��ꓽk?�����&$�Y�>j�1��������|K�B�������#q3�<6.Ɠ;+�>�n�3{Rn�_v/$d��_� �&���(6�U|�,�o�4�� �3���LD�?��u�Ko֫��17M�5R_K�SZ��c'�c���,�S�ۥ�#d+,�Ɨm��y��H|�G���*���h��R$Av� ���~�{�j���
�F+���m~I�R`�h`/u�@^%��V�� e|	]BM !�OZ��2�g�{U㵲�(��c6F��5�
b�w�ri'��Gfu��p���K�{ă��W�^�k�B��W����M�A�
H���Q)��P��ȳZȲ.8�s^8T_���Bt��C��u�.H$1�2�x��7�xR5��i�S�B?"Ƚ�s�39�=X����L��_.�!�`Η0(��MV�����7�g�a�8'T+����f���-~�N��lH_B}(�?$~.�g�~��e4,��8�D��cJ)1ɱƢ(����5%�q+3ֵ�Q4֮v0��w����uK�����h ��x����N��Si�og��z�Z�a��zziƎ�C�!J�A�"J�j����n��W|��iޠ���?"�D/eW����"l��I>o�.�"�}�U�|[h'����.Vզ�4E�m�O�r,�����sY�t+�T2�0��`��-b���E�j7�'X��J-4��j��	p��}�3'��\Y�臆�����X��?</j�G�c��7�U\��+�� ��w-�ͮ8�s8��K4=d]⫓��2�-��u#C�,����֨��ƷEyK�����0�\HT�뗴�P����@-V����7{�߲��S��Vݤk�M��'�x�Gs�T�����/�+�#���a����)��EA��M5����4��{Ŋ�v&�)!H�͂I�0��p�9�޻�T��ʍ8�b8����Wm&idn2��Aߩ�����l|WT�*t�`�BB���V�ڧ��QӾ��+�0[a�s�����hPe&��9�� �^���<�������&.|p�K��>1��īt�t@�RՑ9w�G�,V%(f����'�m�a
\���0�Hy����T�Lx����A���dC� e�0g@���9U|M4�)d~E�d`����?l��܊#`�뮨�4��,��O͘�"����rip�U���L\�#V8^���T��J>,��T����"L$.��pM?�:ʊ�����{���]�m!]c{���1ѹ��D����DސBO^�&�S���s�u$;Ꭲ�z�a���d�BThovW&��Pr{"T��w dv�<�'�����'��#ǋ��LCL�~P�ʬ�!����0�!%52�̗�����Эiֶ�j��3�T��7}VU-��@�XA�|�����L����ɤI��ޛ���!�BW����T��V�*u�N�7�b��˝c��exn�3���e%� )���ֆ����F|�'(�0�10�9W,WɴPک���L���$	�??V�Mm�Y�SCMf-���FRGr��^����K&��1�@�V]��t��H�����ۅE@׋Rf5qo���L^�`��#wG���o��D�]!X}t�X��n�ShQ,��Nذ�<��+m{Ĺ�8eK�Yk 3s*Y�#���[��0���m�î����We�N�Q��Y:�� ��Com���TX���}m�h�@!�=�9�������D��C�u���ؿc����R���F�}���=Vݴ?h/��C? fs;ˉ6K�z�_���8�
�6F4E����(' �"$��>nV�=���6X�s�|�3&���	Y,�ݐYl2��ng�6��v±m�����L0h!j
��#D��U}uC6���E:Y ��yt CVP�릤����&�n��**�X��ؽ��]�R�ܻ����@Ax/�SzNm� �Y2����o�_Ho� �S[������WיWP���׷w���-�@��>��/���&Ѭ�Q5��p�I�U�j�%���E��*��Q����"�r3�"���~�E� ����(�OdN {o���kP��N5�gԹ�k��痳<��C�FQ%|�Ud�)@ I���5�oNR�Q��PN�AL����'.L�A���lZv�s)*F��U3
#�j ,�vw�&14�O�0b$�8L�J{j*}��H�%~-���x�ؐE�ѯ�޸�4�_�Q0I����'�P�L�~�8���4v(��2��Yr�^V��F���4H:oC9�L�ڙ�D�"�U�%}qGw����M��Ev\��s�I�ϓ���"�%�\�>i��b�8=T�2]{S�����z�Z���Lu��HIz{�;ҹo�٫;��~G��Gm��9 ed���)��� KZi�̱DV������=������C/�7+��uA=R����=�݅ߕ�;��Xs+�tB'&���c�	q��������[����Z-�+�aޣٽ�u�#7���C�K������=�����]���뒻]M�.� �w i>���]Cצ�u�^k���%]�u대i��n��1��2͐`�,"Ȉ �OUb���ڭz"��z�,��>|�� t�����gO�^��\K�{	r�wX��Q{��h9�PQSS�kL[��rƶ;��jq�!q��(6ōx�L@�\d% ��=xv�˳(�>���,����A���_.)�>HA.s��Q)E�*B~�5y���yo$[2@����I�o��W]� �&Z>�$��-*nE���''�>�PĀ�T���@#8LB��.T�K�f3�yy�I�0x'b1�jZ,�!��L�OȨ�~\G�x�q�4�e��+��R��s�B'��2�-���=�Ք��nDO]���nZ8~�,dط���t���E��L��X/�L�7lq��� `�N�@CWW�c�^2�GJ�}Հ��Y��!�g��Ûe>�./�<��B��x��E������"G��ݩ4P�x�1���d��iJ7�v���r�X��^��,8#A�e�Zp�	����G{�ΐ��/�����)rUܑ3���A�ǖۃ��}�o[��}3��>v��Js��
&�d*4������V#?��vA	?y��ACu[�v���4�#��Ud��
>�b������C!�q�vUm�z��G��,m�
@���(�BJ�<`pU@����g�NՔ�V22I��_a�u�����*���EzO�W��lNBϾa���lL|I�58#�پ�9����o��7�y=����#�ݿ{~��u{���z�����<���G�����{#�㿓� �N���>���}����l�� ��/NҀ�� >��4~�?d��p=әR�/�� �:ǙF=��ٛ��Fc��j��8�ئ�YS�XܚC����R�%ȢM)B��Ă����6��ι̒G:�U57�3|l�H��Bۮ�Ƶn�M!�Ǘ�3�(����[5�JZ���]f�[*%�v���n֪�2ܒH�{�*y�u�A�S�����r��A ���*�v����.tt�R��M  ����l����b�����d�!}�g�W����]�*a�7.6wP�A=�1$� S��n9Z��Z�5���N�f�:�MVˡ��WN�Xpc#r�Wo:l�> �f%Cn�:6F�r��9�C�%އ�;�v���� ȃ�(_!�w/B`������r7�+۠�����.�.��lRcJ2U�٤Ղx�-���ݼ���;������U�Z�'R�9]UXA�UZ��,���=�y�i�fp�#�x�<S����T;0t��?�����1��V]ѽ��Zc&[�t�Z'�&+-��DL��(�$Bu�Ž��e�74r�K�_�1$(�aA` gT �LQ�`e�˻\������'G�m��K�9�Vf�\�W"ʁ����N�J0i�gEgD�p���(�XX��H��%A��������E��]�jf

tj�GO���)�uW"F����(\�mO��<R23dY��J�	�0�_7n�@��D6�$�:a˷�g�&��.�'��.�����}i<n��Y�|�CJ�S��f����\����H���ɧ"��'��A�m�~wMַ��2���F�WG�:���Q�C���! bT�g���3.�M�3j���e���2(�Q!.�~��z��/d�E��>�"#�!}�}��A��Ǐx������q�=�����<v���=�<>I�����a��N�� �g}��ハ���_��yߓ��m �3� ]R����߽hM_}���"M���G��؏g���y̗&�{��H�^�e��Ȏ��>����-޻�\������powl��m7��ONk9TGr��� ��������U��Y-%�o�r�mR��G�����v��ژ�C�2ܝۮ�b����_F�C�2���0����N��f�����iߊ�C�"�~Xh���~�O�~�k0]l��d��������¢G9��V��W�.�;��ܙ�Ǥʹ�֥{4���&s�V�d��y.�j����ΡZ�ƿ\���S)X4d�f� �����/��
Ȩ�,�bל����<[!4-���͋3doAErۗuU�SN��bܕ�,�3K�dʭ�0~Y��D�թ&�1!�go���c_i�Hbڷ|Q��O�JF\{<��%���iJ���5*"�[w�j��l��bI6�k���w��n $�d4%ޢ(�_�8�{��q�,��\���A1Q�L�ӱ(�4�Az�r#�i�YC�Yu�!����j�:i@��#���C�vr�%ݢSD����ns*�p��Ɋ1�蟿{��t����K�v(䦚�c��G���܃G:YS�n�T��	�[D�zΫ��݋Z Whc� ��S�x�CJ����K��
@�I�3�#�p�/		đ��E"�46�1��J�������E�o�i������陸�z���ř�d���b�!����ʠ��V�H�B����ԭh^�B�lL�����z^T~`Б�Z�ei��[՚u�I���ȫ,@��f(�w/ҏ�qF<||F�G�	��H�ݢws��?~H�Q�׈��S�����~ϩ�}�����TOʍ� k@/0�i�O�T�g�/������+���� �j�<���qҢ�����Cb��Oԁ,�|$-�v�M��վ�J�������e��� �gnf�s'_uN��a�WQqQU#��&�}֯b-@#Y�G��Z�W`~�c��7��x~<��>�I���M�>^$�#���{��;�~��57��<��m��%H>��⍲A��n��d�#ۈՒz�lvr�e9SR��tD��Q��Rj?ln���jZ�=4=����dZ���J�%D��]W����(�(	�VA�:�^ҕL�P*O�:Bhc}���͈[���C<iȚ��;�\�48$����*5�"��k]���X��UU1m�(c���zU�F���W<#��{݉o�q����o.��FG�2�������$uL�-)�A,�ڄ��w����圣�N���lXl�Z�zV���/z��x/=(���(��)���1#��r�����H�����T�H$�Rߠ�j�TH)�^��͂�z�`X߁_�ɗg�:���&�K�B =�%�{U��qE-3i�	�� ���9΃�ŗh󪪔�Q	Wp�
Q���X�,�]eҹ��[����~�e�~�����>��~'��ü�ӡt��n[��sH����_{��N=�^(���(������o�n���G<#�T�����y$[9��ߝu����[C����>�w{�hʔk+��&�F��T�}|��Ct���4\1��lQD�gh\$GH��oyLJ���
��Vzw���J����S�H3p�R]��Ph����L-�a�$<�~�4�*��h	J�����Ă3<�[��
dZ����u�m*���g�X�1���>����p�����T�D[}I�\yr���T�1{�Z��t����~��ThPT���[q_�2�`�I����>�|�,S]�g�޴"Ϟ�A8pw0ʢ�c���+��8�+6z�d+ra�pA^�����%�����V�aL�^��<�\~Op��e�M�v�c=F�[u���� �h]��)#A�m�2�:"���{׮�-��^y�e�hW��0�_��7�� _�׻��|�;��ۛz��ޯJ̧<����){�P_J7)#t�|z���/jg�'���=j�=���8U3Bz��_�T�3m��S�J�Rgk��@�a�Pd"�N4[�2�-�YH��lҖ�T�o�ǅ�d�1K�����x0�]K##�Je۴kH�0=�R���	�Iz�,Wc�^;�v�É����'�^���	~��m�`~�Jz�U�lՍ٢��k1�*��5u�f�Ǆ=�5(��)������l���iSQ3O'T{��\E�;��=k�|�«�Ŗ0Y��/�ܫ�����ة&�j�8���j��nT���i	2�e5�rys��=�T�=׵�M�ܼd[yN�Jw�q��FUf��l*h)rB%mf˖�c%�������~�'�OAO?e��ޙ�7'�:�S�fӜ�j��Ȼ�\�6ܥkެ����TC�泩��^�W�v`�y�<�����b�E��L�������;��yi޼�&@M�E�^ ����c�Yuٛݫ{8���ܾ}'fi�e���>Kh��qv9�kz�.��9�|k�Ю4�k��*���L��
�iߛ؞�do���n���7l3�'�1g�[?>y�#mY�`��ҷM+m�Y
A/]f��,K
i�]�U*Z��#�+��1�fo8�F:s��q����;�f	!���B�M��H�R��Ho�,ި���l�������뎁���UV�|˦z�[�W0+����%՜w��fe�Ҕ��� �0_��{w��^2uS��>E�@�}X�x�i��4�;�e0=w�a�iG���b�d'�Uu�7�	Z7�����|��++	�Ǚl^�P3���dǫ�����4�XW�[J�cKA�F���e���ϓ�۞1h^��NU�@�-��W�ِ�
F�Fc��b��O�*�{0��Q.��J��厹Do��혨�� ���{��p�(#�y)����j�.�;��Yߗ��<|o)�~��c�̈́����/��Rm ���l���M���a@6Izψ/J��
<�^F��$����խ��u:�v����/�zL��Y�v3Ѩ%x	�yε�΅Xv�uVd�[��A�Iy��(�R7WNh��'�DG��6�7�����J�1��J��!�t�UR$;F%��*[/.��$�
��J���n0�4��=��}��5����[�dC�yL$O�0S����h,%�Mz�^��:sA�,>�ꋼ��b���ŽK�6T�n��*G��g�U:����RW�\ܤz���x]\3(\>HRٕ���� �S�ͷh�<IS�n������t;��(�P������I܆�v���i0uTu� 2G_ZO����Q�oZ�18���Įe֟���֒�|��O���u�oYW�<�W�]Z���^w	�v�\'d]E��22gU��a*Y�:��u�������6�v���qδw��׻����X�`�n���
�K�j�55J$`���s4�m�a'GA%i��Nu�Y��j�_W��%֝��.H�������ƨ�2��i���>�a��~�G� 4�g`I27ǽ��;ř|�e��E���=Wv�f5�A0�X�v��ر5O��V���O
�C	G�#��/G.�ݷr�Ke%(���R����X�V� ���b�%��͔gG�u�j�x�B�y�tif%*�UDݿ�Xw}��
�i���[����t�2�����V���Wn�KdҊ����#����يV�#���Y��\G�,�.ï��Ci���\�Ǉ"7�T!���=�n�u��7���e��n��]˃��*��pqv�)����&��%%��x�\m���h�K8Y�iŸ������+0��������9uט�e��t3������,���n
���Zf귪��Qb=v$"�;�	r餲�&2�f`ަ�.s���.U:q�B��mi똺�2�o�kE<�G՜{d�y�l@�X���������0�mF�H�$�4�NI"|��[m�z��g2��ɑ��J��3,���,Ͳf����N��4�3�,&�o���pl+i��ʛb��e�C5�WP�d�Я(^������`� �ƕS�}iaK�uv����NV�u:�(#��̕��Q�gpS_%ї��6��;Cr1�X��صcX]���3{z�;mu�W.��_h�VQە�J�����7� t鰀�a��{1�-A�z�Q'�4p�����%�d����˅�:"�����1�K�?�
���F�*�I*�X��)Z'�@�b1<��s4��ܬ���>>-ku*��Tࡷ˨K�+,d4�C+�%cc�i����|���fNŐ�LW_��,�|-$�O|����吮٫3f�� �Ye�ؗ$Эob&��7h�Į2S]�[3���.�-�j��`�E��a�1�Θ���F�Ɩ��]�.���H鶗Y������ԚL7[�YFBQfbHC-�їJ�0��"c-�JR����%(Xq�`VK�ߚ<�fA(���1�JG�aB�lA[6�[�'W�7\�1i[R˥�-1pi�D˞wH�s$I�! ���ɠ-�)�Hc0�����an[�l�ս$-֦��J�XT�����mҽte%.Ka]2ǳ9�E�q&�-�&�\�X�휵+fq�s$ZV��ڶ[ubE܅�䙩�3g1��g3i)�,���	k�"fؘ�����Ks�u�6� �N�.��k1�kiB&�jWZ�ׯ]��X�ܑ��f�����Gf]J�&���h��U�           �ܾ�"�|��;��i��|N���(�K�w�0�g�v��ƹ/�'sY�le7ҫ.��dQ�*���!r��܍Ԭ�;��V7�=����|���5�̥t�{M���!�T��Mqd���s��cx��0�^ B�C�Y�k��<OS���t������x��{�ݞJ�����/����)>�/E�!�g�#HG�G��C��O�ƿAZ�����k�@�X�����~[;������
�������+݊^9��لh�C�$|�!�K�H)�#4�2By���T���~�VA���_���>�FI5��}�+�C��Q�P�i:���O}�O$*�"g���1��Ǻ$O?C�����{|����﩯�����H�G���y����)�? [;]U�������|��e��>�lF.�i5Aj�Y�?|������O�@�? �*$����)ϓ��z���So��L�!��y�^��N��od����!ۨ ��Ǒ4E�;8����(
Y}��ș�^7����4+eH��<�X��'�#�#�>P�*���3�<_�=���8�/((|H�|b||{���������%(GĊ�(~����l��:E)�~O^=}N��?����}� �(Ofc�"Dp",!n��G�(�ޡndiTU�b��	 Y�rG�G�_"��lk G��gᗾ�i~�|B
@���G�*f	�O^�=�9+m�� ����H��!?���8��S�?�� �)�S�����E'�[�� 2�dY�hYN��3��z��}���D ڧ���g� ,��~��4@B ��#��z(�*���օH�r�
��	���"�����i�"~��������?'�T">N*2g��y��%���_��>����}��b�������υ�=��~�ټ%slz��x ύ�����~����X >I'��o��D��������{��>=�g�_�=J�Nߤӷ���?��*}{���{�L����2|@�w����R6����޲�ȁX�� }":ct����x�/]��
䩓�J�N�C�7�r�=�J������{�E3OS��+ǒt�������d���T����'��2w���
z�8S�|���{�+ʡ��<G��W�?���w��7�(��������~dw��4�~d��,��a~��^z���������_��'�C�g|��������&Fli�28��#0����#��S�>��i:y8��������:=X��S�i|I 2�e�A����#bh����d�%��l4B���n&�3bB�>�~A{�G���Q��<{Ԩx��)�@u�d<����z�Z�׏�������a����^�x��ߧ�=���?�C=߾���O���S�N��ɞ�޵��OG�=O�f13���p����﮾߂��]�Y4�c#�_� �\n�I}m�&Ebvee��Q��wb��p��fU���g8v���jXr�E�)�]�U��VԘ�d�W^��|��>�LH���0o����!��z�^�S���4>'�k���'x���{ϳ�O������:�������|x���|OP� �x������������}�a;׽��W��u�w)���'�������8ـ�P����_�=N�R�a>�N<H��ֱ8�~N�����d��ϟ���<���|N<{��I�����P~��@(�H��#����+������|OPȿ���q�����=R'Ȱ��O�����P�0_����^��{�a��Qz��J�2��Jx��q�N��p�8�NG�~C��>?S'A��~c���d�2a"�Pwt���+�g�6���D`��!����k ����{��)�ާy��~;i1D �L�a���8��߰��?��>���Xg�����{�w��93�����|z<z�~�1��~{������i��~OP�?ٹ��&d�)V9ȍ�c����L�s��=N�S<y=���?�z�{�u}z�`/#��_���������~���ys�,��>���ר���
��W�C�z�)����T��p��ߞ����%�w��"/DY7�]1�[/�_�b�*b���}Z�hq!z�B"���(���A��<{��
���׃�䩄P"�:�U��0�E�"�"�"�"!�
T6}�(~���0#�_|p���7�|G>¿R��y�!��=N����~��E��[��].����QK���>yhz�Nx�#�<�wD��<T삑蟤=O����,<x�����$����T
 Q�}J;g��D�s!����ǟ'���*T���~���O�~N�'_�<E��$y����o<�+�����W��Sn�-�i��y��Li�%�g�~#��ݒ���)��M�9�߯�N�$?���I�|NQ����肋��L��;�R'Tl��x�>{���S�{_)��'q>½�������|���""���ݯ��2���?zT�#~�>dZ��#���y1�0U���g���O�|C��^�������W�Oȧ��x����d�;������?i����O�U��N��?�����|NS5�Tc޵2��߬$A1�D���&�]9�.�eJBn�w���?�Ƿ�S�R$�g�����?��|x�{���QO��oz�{�J���d2x���|�O4�'���D���X�p I���b�(}G��$�|Ǔ"�D3�(��}��uD G�mG�Aj�������~Ę�F��l��B͵��9��[Y�٬�ve<̝�Q��e��`���r�y[Xef�U�ȽC`է����)����+]�o
��ѝ;��t.��%�?���>�~V�불�)�?ӻ��������r��c�����=M )����h(-O�So���d|�.p~#���M��?	����_��S'� _ѓ}�yO��?'���D�/���b"<#�!�����u��Ͽ-����d���T��:���cu/� @���{�)�n�x�.��~ #��� �}d2�d"!�S�"z����~�������i�v����������</)�c����'2Twb��Ї�p��NNVߗ�?����Ꟑ#���g��~�?��|yC�S���R�{���j?ȡ�W��m��'N��8��Ǐ�<L��O^����PD?�yNw�ܖ�O���?Y��B͐����<��"'���������'�*�׵C�rLx����	�/S���wV��x��q�T�c�=]�h$t��C�Fn�-��ۻ���cN�zc��G`�g�h��yT�Ys0V�����T��=�Sb���LS���ca8"������lv�h7��M)��]��������lP5�\��8��$B�7�e�ZpD����\�&��N��i��O��:
1O������Y��Ӆ�t� �-�2����V�66��� �J)z~��t���͞�{����h�l��9�A��� ��($�8���+���|����z�����y;İ��T5np�t��ycQ��oT�n6xgK��WQ���P�Ҡ���a1�=���_�������h��ςG3�d�ų,�"��j$絹˷��;�|���{<fbB��˨�lz]	��SR�ȅv�ǍU��@���$�ɸp�z~�J��Cgt����ף.��k�3��T&�a$ �2�o�^�u�|
��f�,��	wJ����)'����w���ʦ�+�O�Tz��@��X�ޫ�[��2�:]�ri�\��BE��\�L�!/�?�C3Pmh�	h��L��hgm
5|ձ�B����J΋6��7D����z���4�rﲐ��(A��h�.�P���ݤ�ɣ	]KI#ںˤ�WbXk�Y���K�m�-�.w��|��5��U�kgfۨ����e�Q���d��M�A�gc\e���(��D.I$�w�e�f�X�їx�H�
��h�AI�1��^s7i��a��q9�,&0n���|�z����!f��䠰�=��wEz���~8�Q�)�ߎ��e\x�,��SCp�q��Od7�������*b�9�V�|Uz�>[�ʋH���^7�;�ꜰ�GTA8�=�o�Iݕ�!5ٶ�{5�������R��X�'��(S�����U����8�}�B���s�{��8H$J�B 6�%lL��,����z����Ul)��5w��E8�G�� ���r���LH"��pu��g�m��zҘo�ws\�nv�U��8g��%U�������䋊� �7����F�{n��坾ǡ�ĥ��L>~ۨ4{U��'�� R0D�׷R����������نjq���N�0��n��>�qJ�4�)�������w��T����.�
�H��s��ڴj+E��ށߜ�Mۼ8�&�o��j%}*�R��2C�lЫ6A���Z�xx~aB��1Pp?iO8�a���ꊱ��M�peeΞ���9��	�3����)6��ӫO'8W�c9�-ʯI�j��@ô>=%%�5)�n�5sT����&6;�}f7�䷺�=�|`�#=qU �♴l��9��.�!�J����:��ևl~���a�]�zc�bT�*����d=� �g\��;�D�9��=�:Q7?(3�g��C�Z*��wh�i5nsήጺʕ�2s/�W2��,�7e����nP�v����]7����aW5�]QUֆ�/���R�'v�U3�SjŊ��n���S�P���l�=��u1�\L׽Zp>ȫ���gZ��M��f'�ܵ�j��L�tRR��Wʯ&a#����7fT@?l��am����D���' k����
Qo5�C��sXCI�0m��s���vD�t�A"�$������]$�"$��u�]!n��R�k��k>y��46�U{� ��9QC~)�+�{��K��P�.9�]������u�.����N��;�F�'7�ȷPމ�J��-o�8��`�4�u>�m�O�� vs.�;�m�L�P_{#�v>j]Kb���[��)\�e<ˬ�*�qQ�a�rz���b��;]_Y@�ٙ�C���LJ�^)=i��fQU����5��>�"�'o�]u�c��Ei7�&���c8�����z�����	S4�K�4�H*�R����9�F���)z�L֦S���x�}0aOf���>PN��~�����Q���v�S�6��ݨ���;�<g�!=��3P���:�!h���0��	��&��T�b
l��?��J�l��f�P>�s�O�*!�7��{� ���uA"η�*���y+g5����M�
��0�o�����T����>t�3�s� ��{�pk��p-��*�is7U^L��j���`��u����'�������������Y�)��ܠTz�邧��0%��S;��u�b�~~H,�&|�ܶQEv�����UT��Q�$��`M@�����g�x���!Պ++��@31U��a���D������g��|���^L@@�ۜ���o6���)by@�A']*U>j�J7ڙ�N�s�?{rylU���o�y��.N��sed��;�ɪ'w(��"�s"v�k����݌ޝ�hN�V��V�Q��ۙ�*Ķ��\;��4�܏�Z3��251�Y)��^E,	��TB5N�v�ӿ������3�]������X2���X>M�p�m�۬���~�����~E�S� '�Ss9��I�/�YQ�g�x,'��lK[����Vʥn[o�m��L&�$�)#Sյ{=f��Q�F>\
�D��Mzt<���ܳ�(�T��6M�`'[W)%{<1d��k�[L�9��&���P��u4o1<��2{�xw/Ek�m��')ݝt��q4���&����Ï^e˵B�=oj.�I��Z��kj��꧖��(�O��U����U�V���z��%H��Xc�i��9�܈n�4|n�Գ���g�թ��r����`��a��vbOf�C����Ʌ�����^��W6���H�̬��#�Co�q�u���]��;]�BK}Ж���J�˞�۔(Y\��h������Q�pUU��4Hɏ�E]�n�u&|{3-�����	��%;��>7��5�j�8N�S�-��7�$��(����T�R��_�&�q2��j`z�M>�ۓa��>k� �ƲVALb�NԖ�шSB�����>��Xp�(cO���#+�H�W��������:�_ `��,��.QU���k�����z�8=���f�n�v+�ק��L@��ty0|�{v���{��֎�u6�S�VZh�,9������RB�ݧ��"cR��bry2*8��q� �G1s�����Bc[~���� U�Jt
��ә�(�y�Tg����)4�!]%%s7��e�9��f��#�����b�ڸc��s�KN�����E��]w�Y\%: ���;]Ɓ<�v'(�DVbu�k*��42^e(�����������fn�oTf�_FT�u�{,��{�[7�h�~U�_'��0�w�.�L���.�G&��9���uo*��3$
��3C[��W�s&}O�A!U�z�ڧm����X9)vC�̉u���q>��J����Ɩ��l-7ͼ�Q������#N��h��5�:��*�����FgMvA�5}]Њ��
vR�HXZ��9��d����s���^0GaQ�\�c���Ę�a�۽ė�6��u��5�3��ϸ��<�cv�� �E�z�L�w�G�����k���$�wօ�*ӗ����I�n�^�ݚmR��+y��V��{����������W<�8|���)@\"jbm�(=pv:L��F�P�Мn���S�{�8�ۨ�_o�M��?�T܌��W+��"	�e�!��el�e��IA�/:�~	�n��V�o%VQ��c�#~N����y�]�}�C��k�9Yt���v��\l�P�UQ�z�"��9��m��t�V�����~��pMMUP1F��X�������6m����J��ل��]�c�k����`��{��,ն��k���sfeⅼx1A��[)Z��?SY韇l˝E\JN8P)��җ�!]r�.Ut���N>�*	����3;I��<A����>-�ŖS��xJu�;�/�z�T�u�I��U�������?m�~<'x�H�p�C��t�wI�(y��	�Y�'���׀��P�������~�%��5���,��� �ﶾ�v�o���߸g�2<��Y��Z�Uٵ��ɽ��5�v`��,��wztҔ�����L�ېqH����0lۼx��	;b��.���D��DК���ꫵ�e�u�h��n�����i�w���'U*��8���Y��F�E"�4WY��b�R�{<Qχ��ne
ɛ,k��a��H[��u��@DRKr�6�li�����;�5�?��������3u����L�/,�m���}�>�rv2��>3`T����!�uD�$���u^2�k�WS���t­�mˢ����O���,Wnm���Nr�i���^�E���[^J�T���� �R�R��Y�rҟ���0����82����W�O$��O��ͺ�Ξ����]�p3s���mz5��� �{�ʴ@<N�ɍ�Q�L��~n�;�)��[����L��ie�l��9Ux'�g�턁���g[R�\5Ij���q_2Q��6ŸzFLe��LM�����R[*��max��E{����T���'���MMd�&{ԙ����v�I�U�L���ޞ�W�c�-��������1zA�8��7C��ۙ&\CN*
��N��1_\��m�����RR�Coݎ�iy��ɯ.�q�����B���6��Y���0PN84�w�n'��<��ǃ}���	�y�p�L�K�~����M[�Fu�"}�\��vD�P�>�1UYm=���<�9�/��'ʷ9W%�i I�r�}^���ce�T��fe�ߪ{D���}3����
)�9}7`ʫ^�Amf�L���OnZ�*��^�<g���dЈ�v�S͹�~�sJ1?�~�7�_N�?j۫/d�z<��e�v
b����c��?$�C�E��J4���ݯ�z'�GjŶ�9/�ii��.�&����)0ٿeby�5Gu�H=�-yU4;9���bA۴Z��a���*���'�ww1,��1I̩��D�0�}6�<�O|.�_\��� [�=4}j�x$��9�k*/ݽBe�Ʒ��;9S����Jvޘ�]�@�ٱ�t1���mG����9�޻8��*���U���I|���[�u�0C�uEt�#�F�gm��͢��J��gO�z���ʶ����V.C�D�F�^Sk�Ɍ���U1	��V��j���A%� ss�M�9�x��=MV_�ָ�+�������m��d�2�_$
Al C-7J=�m����&�d|�Х&ு��ͤ��4t!>.����ۄ<MC��LQ���Cɫ��y���һ��s�I�:���ZXD*�mᔄ�͎�������W�6����L�MB��`ur��&=Kɭ���*�=�F�����g�EO{��P0��H`��&���p���k��A�*B�z�/����bF�e�s�����X�uZ�L.{%71S}V|���Ss�D�n�dO�^y=�Jʳ�چS>��<PD���u����W�LߍFrx��R]϶��+��e:N�5o�z�8i0���V%邎�쒝#�W�iŲdAB<�C�0��.5wM��Z6J�eu
߳k��aMm;�R��٧19!n�O;�7�|7�[�7�w5;�K�;�U�ro�	l� ��3]���ޮ��*{�i���hl�'{�*i��!�s ��s�"	�)�7�܋��j]UD�]�cUqQ��U��t}�N���*�H�����$�	�6�6o��]\��R������/�x�=�~FG8N��v��%>6�̒�5�Sm^��8&�F�>��U�}�c�c�e����O&��s�)c����p������t�]ˣeX+m̝[&��	��=�����Z����U�7&��/��v�U���ଁؕ�xo�ȶȤ�|��[�8�V�9U���ޏ �n�ά�:�L��P��ghKs�-8sl�Ѓ��F����=W�\N��_tɻ}ϯ���\K%u������f�G��5��z�뼡x���ڴOb��Et�^q'�Ἣt�\��x��"n��N��.Z���˞B�:���k���튠�����fG��m�[B��K�BF�����L,�N�m��('{�!�S�*�y�eƕ�*G(�S�n'G%�y룗���4�7ގ5��n[%Us[)^�ؙF�����>�{77�ܛ�ee���=NJ�V��3�>��9���yY^��̟lr+:�ĶU��mmv����l�'uc��EM;���V�U�[��w���U�<2-�!H1�̓����T��.�1s���Y�[��M,9�u)���:��7��0N&�8�@��M��3|�R(1~��|~��.�G����=�L����7�A�S��M��ګ�Z`��"Ls��}cU��vy����Ĵپr�����b����ל^���s��CW��%�f�ʼ������h��s�W?xK��@C�t���p�6�<&�FկKlW���i*�O���<�����n��,�]d�W6�b
a*���Tr��S�l|qgJs.�խˋ9&gJ_�_ᐚ[Ò��<�t3g�.�XW��m����H���=ل��h�D����hqq���G�2#�P�ג��8�����\N2?)�&} ����AN�yE_� �q���'�"�}Z���{BUV�/�S�
�W�߆�.*�N6}c�n�=p?�'���H GQYj{�w�Q��"S�����zGߖp�)�����<�轭Sm�G��Y]]hT���&�
��Ų�V��T}`�����W.ԃ�uu&_<��a�v�W3���2%�	Tc>#��1�)�����鏵pb�����ھ�y9w��]���W!Q�x���ۙ;�^t�ڭY+Z�[�%K�K]J 2&L�Y�s��{b#��}n��մ���ۤU�+�W%zx�:�P�(�:��V{4&2�54�.k]�zJy۫{ק��`�e������1�)Ki�����8���ut͙�/��zyb�Q��+�#-����������9��euKd��WǮ�����j]{�F9���z��4]�w�NP_;��x;.���̰�h�{�_v1�(�R�:!�I����N���|2��;����˵˅������W7:�GH�����i)8����n����-�܊�۝�۝V4�"�5�T���X���\7+9c8�s(�j��l�<����m �=���V]*�*�h|����b���i|���������e�ݪ����m\$|g^G����9&B���|���=�P�qc ��n�9Vû�ڏ�� �|e�e[�>�\%T�v�M�uʐT��.�̬�46��V��kJC���v�?<�\�f������� _��&�{�u3�S�Y8�P�����I#*�R�Z���pKP[��N�4�Ott�o\���2�7&+؎\��ٰLX�W4�iZޫ����)y�ho�O�����]����/�����Oѭ',ɇm���bk�z%��Z��v!�Ӆ����&_f4���d�vƌWz��wsv����4
�L<nY���jk��a�?2�X��)|M�|ੵo\���R�Ρ�9�f����#[�v8�{�ҟ�Zƺ�M��	w�>�9��$�vӖ;%i��ٽ�:k����]G�u���	�q�Ʀ�NYB2�E�F�}׈�Vɺa��r��ȕ�I��6�g��B��=Yg��AuAK�yw[���^�r�i�)*�G�����dHH�Y�6��g�M;}�n�.��6�A��N����
�o���⋞��
�R߸n~���{H�����f�;����'H�5j�%R�(�Uzᣞ\
>0��(J�%�Ló]{	�7*vT���Ya^��+;q�MC]4��r���l���m�<�>�ü�)ɑǪF/y�SS{��Al2da�(�}0%n9�dӿr"&~����ꭨi�zj2i�l�i�'�fV�*�}��^��lMy�^�5f�͸��J�����+���]�[��9U��^&<窻9^U�7���Gȃ|�a����̳�
�����X*���(��Vj{+��\��}�&�q��x��;p*���d�xU�q�v�̗)�ϣ/tUx��UU���3�N���6&=	�~CW9��ڿ�f��25��U�g�2�U!��]+��8}���9q�tddr�&L���>s�$ �"XٌX2Mq��=9I�~���x�/�U�̂`�S��\�*�����H���+��n��&�	9�k��'������eeo+MW�c^H;>���x�M���meP��q~����f��=��ѱ��Y����9�1t�2L'r���fe��\��čp��V��a#�:*䉨�|ZySx�v�k"��B>����������!/y�۵M�~K�M�H#Nk�ug嘼���,��d�m�3�Z��R<N��_���Ta
Zo��s|��a�N��m�!:yn=v�*;)���i��m���G�x(��1�ݔ���Uq�3���^��#��0α�7�U���bWy�*��/Fn��l�ʄ���Em���f�M�(������VZ���z29���'�}�7B���N���������HZ�gs��v�N]�Ԅ�R�����XsNw}Jͷ%�gXۘIH@��Q��P0C���0�RH����u��i.�F�M&�e[�`J6��/6��t�&�M�kꐶ�?�ygig/�3���!,���&�fg��&�,���mum��j�!I	!Z�4���ZQ&�m��3SomȪ������ ��,��w��C�'w�(��^�ҟB�_F9uw�D�w��J����;��m�3s�L?�`��@����
����(�{|���P�_�f��`_�1aA�sys��價ӳ�`X6�nO����+I�Qap�ǅ�Fg�����b���Q��~�	����ۻ2J D�C���~H�����+j�Z�k���W���X��m��b��kc����+aP�+ljd��%��sd����yu���b�H��F5��uyKq�ء��àV!�IV�>�/f�&��l�s��#��z}��gg} �>��\���z0��#���l�NoV��[X*ܫ�۪�mJ�0�SR��׉˹�������8H���NnTW�/�Ǜ՝Lc��lW�/��Ht�L�N_mN����v�&ӸyU.���p�;��fYWXt{�̩c75Έ"�hy5�j�I)�.kT�w�>�@*��+d���ꞧAOVT���e.!>��ع�bs`�8�hZ��җ���n���̥t0����lQ�+���ʳ�G������k�aUr��$�+f��L��{���K��\$�홥���z/���wS�5��D�޲�%��,��1�����I���b�zpA
qT�*�z&��~eK(]�S�k`v-88�Oǔ\<��6�:�g��Gm��^׮$�K(����^�P�v���c�@fŊԇ����^�Y��nt�ԵW���IŎ�=}.wt6�B�	��\�YIΏQ���A�:&c�U9�|����3�%:����c�mYý Oe�>LwPa�y]��o"���718:�W��ݸ5����@sɴ�o���&oP�Ū��]|Y���Y���Ȑ�W�����m�~�x�l�靱5�a/y��M��`y����J2߷D���Zѐ�y����eyem[�^ꔲUz�_�/^��W��T	�Hm�#�S�I��ۆ�b�����'���<�J�JB{;�(L��׎��8GU�	bh��UKNI�T!�Z+��ݏ�4:���S�����R���`���?-���*Y����VF��' m����(�c0**�4ڰ��<@[Į9;�罫T1�v.��F����P�울w$�;�U׊z)1���<3G~����t0R�	A�i�N��Q�=�m:�o�W5���<��D��v9�\-=S?y���Ю��*W��F=϶���E׮��SC�G'�B]�0���ʤ�_�G]Mi�ބ�����{!��n����3L��&^ri�)���ɫ˹�_�l%n�'.hUj���)MW��E��gzO8P}3�s�w������׭Bz�H ����᷒m�9�īM�����YN��{�Yb����G4o�y6N�V�׺�������&9W4��W$��)�z
�Ϸ�جq>��qM��9G�gޫ�O��%]|��ƌp9-E�8sbWݞR;7>���f�o���h��6�����o��q�kf��뒪8�&9�5�K�4�a}x��9�MYMF��yH&�"@H�`((QHEES �}B����QOƀ� �x�[F��"����W�,9cD�s���d3��3�\�E5�d�#��L�W`����Bq�R["U�צ���`�v�􄍻9��gu�1J.�{�+eśJ������Ƈp��ڶ�����qYD#�LQo4P��r�py�ۈ�L��D9};+�f��xT�I�!��q���t��I�q��
X^�HS��u���?��{"���]�0N��"���{�<ڛ5k]*u��~:'��ǘ��yEU [���CZK2�A5�6٦��F�Cd��_�M�iܝ�E����8SjjT��6\h�<VfU"�^���¬���H��u=D�醫�w��%��5[\;*<����
T�kX�y+p�d�n�D�T�޼��LP�qn�����lci��fҼE��34R�ͻ�Pn���~���1s��k[���|��Q��,�.eA�S�{��PT�=�nFz�O&΃�BfD9��}� ����Pt?w�g���MBW�Ŗ�S�b9�4��'c�'��m@J�J&vk��,���rږ> �?O�̮�S6wz���PX�׏?/K�3���Ll�;d�\������,�ך��}]^�������UG��}�u��ʥW�Q0N�Oo���8o��jc��i��A(�	5A�b[H �*��{��Л?-&Ur��b��-��H���z�������>��z
���Lv����-���Μ�L�w*z�n�8[׸�7&��I�P^�q��Dmj��B���碁B��#>�Ȥ 
Ѝ̘|h���[��׭W/)}ȶ����Wu��J��q��c���hC��?Y�ςEW�+��5k���ݹ�]+��ģ�
Q�O̓A^r�'.��Ky\p�M���w��wd���;I"[o�9�f�cF��m�0��c� n��Mxy��LC\A�F%�{Ѽ��]̡�1�<ކ��T�Q{��"c������.�!{���m��	=�����~������'iv(�P$�����������P��Όf��X�e����
c,.K�w��I��:]h���/-T���4������o����>���c��u�؁|��I�d��vII.�Z���p.b�bʻ���I�׷���
oE5^dR��n�n����E�����n�ϗ��oϭo�p�1{s��	����L�UU9����U,�vv-�ip�V�z癪������L�^nW(��"�A���Ή(�q`ҭesNIV�(!W���< �v��0z�;-�G���,eJM����)��q4ђ$�D����~���5�� �2���J����HU!������ds�ȳ>����m󇊩L>~'�<��+}��֥݇�4GFGC�~t1G�ؚ�X����]��E�u!:fǴS�6ǳ��@0��'����}}B��b���J����.˸c�>K��*�+k�j�B��tY��ı;ҁ5Y�Wߟ�WZ�I�>'�+�kq�TE3~�~4�ޘ���y;�v��iMC�W�I�آ>�~��ڮډDR��nT:y\����
l�[�:7E�Q�Ca�lg�FًK<�Ot�>n�6d<=}��@wy<zD#E��rf$�W:VT�L����������%�ŝ=���	�._��H���@܅��rT�k��ü�jk1f��l�����0ʆ|˷���-˓9Ҿ�N���[/s�Y��&��pw���Lԛ�/2=�8H����������`V٤��0�t��K�KM��o�Y�ˠ����e�ظ��w:kzي�Z��]ja�ze��l\�����t\�c�we�.ꤒ��8m�+���K�$u+l��k�m��B%
��[7�kr�4�f����y� ���.g��H�LֱR5��r{�{���|v��!+�����Sk6�sØq��Ξ5� �����.��!�~�-.�lj�=r����6ڇ7���Xv.OaL�N��oo'��uy?��B/z��ƽ�Q�k(I-��
@�'�t�z�9B�7\�X�.ԥ̤�Ey��*�K�v�(���8U���_���m&V7I^�K5�LI�i����"�^���y�O˴�;�}p�U�fb ڋ3�Ngy�+���P�����i�����_e�p�ށ(���-�`1�/�:��mb��}�Y�B�#o�s�v*n*~�As}�B�A���lU;�a��RDdO�+�;w4�A�a��80��;k�R�]�*��Na��|���)b���W��|�d�P���?x�N_����)X���P��h���9Q@��^�v59#��~�p�o�]l���7��|��(gB˙T� �W�u������@�z�PN�Qw����<��,�^��l�g3�}��Gbs/}��t_��4n�z����|x��>�a'2jk��9z]s	�8d֩��J7�	����b���gՁe��oG����9�E�\;�lr�Z�ޞ��k�0�%qj�f�R��S�F� W�k	��E�um����.~=ș�0F�eA1Wm]d������l��k����^�16��L���78_<QC[�c\�fˠ�mN]�Xݔ1�(��'�J���*M]��\��o���vu�����d���Ǌ�8�E�}�%g���\�bʆ)��B{��PE�� ��$g�o�f%�go��,L��n/w#�.���h
22?<��3A�KV+(��1�Ä���lȟ��J\�Ǖ =C���h��%^�*����;N�+oь[���B����ޓ~�Ԟی
�F�ǈ�dG��6?I�/�j߯륂7	3)��
s������v�O�;���,�����9���}y�z/H���Z����	��E�ι�[����Mw�!%�/O�q*�7�y	�;���م�ﳼ"�g�4� 5��ʅH�Y%q^�Y����	�tĈ���AS�fD\:q^8�n^���PiQFc޿�sf��=�Pd-�m�'�����;b(v+ok=(Z^93�Ǐ���͆()w@�=���{R�S������̪��Fz@(�3��v,����1������jU���"}�Z���wٗ`s�k�Ǵ�6�]�6����c��e�r[�,Kq�_�9v��s��p؍m#݌zV���^���jRu����XŕB�1��~g�1u辊.�n���<<��%�WV�{��NUz �y�Y�a�a�Y��� �/�"���=��-��+|�ʹj5��|�iIU����Q(8,����T=�4Hط"��W�fa��ƈ>��̩�|�f���G�������5���r���*����Y�W�	��OU��6��tz]1C�g9���a*�;����"�n�m�*�2l��p�ݰF_t�}P�S�x���S\&�y�px�����g-S�V�;X2ծDm�;d�`ש��UAw��ǎX�:L��,��d��s��`��kPZH̰��X���I[w�����?��%c�+��ǔ���W�u�ջ��.��VzL2�Eϔ�\�H}��{�ٕdM�R���̹���j��z8i�bdL��=��WwDؑS�6�!o㗶�on����þ�|�<J=��|��~�4aJ>[��\���ʓ�W��s�K[��'����B�u�т�@>��<�>��G��"����.��R�P�ͼ��[ѹr�{~ւ�l9��!ή�aif}�І��3p:�d��;s���Kẇ�V�"v�h�Ѓ� ��)�ie����5�T��(��Q�+�o��ew~���w��UO{@i
�>щ�.Ud�mI��=;�d]�;�B<��m0w����Pc�0��8<�6u��Mw?���l�`�J5���<J3��L�0~����U�*�Z�ۏb�Ϟ��Q/��/�_���C;�_@)�����eT<��]�w%�&�:�˔{��F������5�;��P~#]L�)@1��A�A1��f�{}(F���?x���(���.����v�}PG�/!��c���j��P5��@P�33�.�K�a�cHi��L���#V��yQ!C�w=?�#Ѻǖ�;�J�v�nI��^����nRM-�9<w�L��DS���CKJ�k����6��N�0S�O��zs�_v_����s����z�$��c��=.�ݘ�����9���U�Z�ym�D+�UzF#ˎ�z`ϩ���{��"FgNmt��}Ɵ�aO�C��&9��$"w�X�+=�~N5}�W�F��N��Y?d�#ٜ�I�uװ���~��f���;?y��,K�mX5u0�qګ�3t�&�:,n��[��&���I�����԰UL��(�2M_�2�[��.�`oz����H�dTj�x�B��m�c-�)ڜ���V�?W�o�|���kmS�9��>��C�}��OY��*S�)�M�Fm=�$��syz��C���IG�]J����/�}SXܪU��6#{���O�����b0��KZ]�;��l.���_~���~.zO��(i��Y�`3[M9#�\v��y�`���̕��O�������j��盃d;pr��9��v�s��c � ���`�~Z��Ҏ��Y^��N�1�7%�w�:o�b�DZl"Ȝ9FY�ǯr	�T���QD�^Z�j��'(�>¡�a�u�,b�c����aG��;m�?);�4*����A��[�<�����ߛ�j�;���+��>���g}��c{�ͻz�#f/޳酟H���b�����Э��>-G%��9>P������&(�S��q>��9�
���]1X�q��>X�01L��'�5�.Nw_�&e ϯ-�&��Q]����h����5���Y�}߮�qe"]�0go�k�oi?�Nܷ3�2j8�2�����r�%Cx\B�����ޑ�����{�1�6�m�ƐƤ�i�$F9]1���1��!�I6G[�i�ͦ���Ю�S�ƫ�A�-��̌�հ[���gO	�l.X�f�m/D˭��m�H]�[�,H����1_5��I.ͻm���yuXپ�6Y?�C��LJ�������w�4�G��M��h�/z�`�z�Ǌ��&�߮6�6�Ii�ќ�{l�.���.j��f�)�$XΑrL��8�����U����;�w�M�c>\�O�S��	�(��>�U�ֿ����E}Foc�7���}�|�-��5|�������n�q}g�C�E[P3qwO1B���'���yr�{�eא���O¬-�������ѹ���LqG���ݫ�ZU�<�=@��y�{b�/�q�ϊD�������D,�Ӫ�0UMp/����V*O'�ov�����a<�����`�t�i�nN�8�&7#y�1���Er��/�z�p�,�g�Up3���jm�@�u��:. �n9��)W{�^�[���=Z$xCw g�*%���E���"`,~����d��(�py�B>�U���:9雰k���ƒ�<=���S��g��!3ܠ��q����iV��u'z��Z
:�J�P����<>��sԮ���Y�U%��22av��F�콸�S��]�vA�`�#�����&����<���Ы�׮�K�T�d2b�5�u�n��L��gNC�1���(s]��)8��?�bg	�Ө��6m\Y�pU��f���B���Uw�*313�Ǧ)x�����VF3�:]i�'u��s��ݹ�8����
����kƨ��\�$�{�E;���R[Y�v3Y0���ۛ��ɣ1d]�ܽf7c�u����d����oQ2j;�7��O����m�n���HB�T���-їn�_I���M��^:����Q���7�&��������[�W[ӞmH�~(\�î��Pd`�(P��Tm^��)^:��ouR/�7z�B���ת
S�݄]ޚ�˙�J58����U����.t�+��j7�K)d��ܨ���s���B�5��ӢV�/���9���m�ṍ]����ڞ�o����*���q/ww*�����w!�e�۝')��d���l�&�WQ�4œ��j]:��{�bV�� E!y�w�v
2t2`�0��n�	�fK�)M�W.���n���ԛQ]�m]���X�T�ɶ��td�S ��۹�BԶ��"6��j]el��˫�uq�W�1�;B+!糪�"w6��r�U�&�u��OF(�s�m���zE�'^]C�^�f��ӄW���'0��&�q
�<���V�]C�ٶ�%��+��v�\��d;�pL)�kb�:�M2�YKEj]X�o�z�3�:^:��Y�A���U
G=�EK,
+m(:;Q<�9����t��>�q�s��<w�dW̵��k
uM���e���ʝ�x1��l I(;\����n��r�R�T��4���%��H:·�Umv�4��wqê`I�=tO�R����jd=�ش��YCU�8�&HB��Qo\Ɯ�����uU=]m�29$�H�n6�p�$��ҍ�`��W{���w��n�!��(������zxIzn��Xk�bYV��&fT*�U������grFcM�S�%�\�m�Mi���s*�:���a���N�u�8�iCP(@�v�Ѽi�M�V�Y3z�s�>n�]�Ӽ�}�.�IT�2N�:0��ړ(�,�B2V�۳��5��=ʱξᇢ��}B�<b�J�*'i���՝ꓦ:�\*�W%y�Aϐ�G�3��Y�)�p��4<N���ԁ�Y��&�
���p=p���f]�ƾ�g�v\�j'b��u�^�ؓM�&�o��ؓ��H�ͳ���7��ʳ�FZU��l�Z�H�>V��<��#m�k�ڙ]u��)`i��y|�˿yM*jQ�,�X�/�E���� ���%{<Y�ej4�2��K
���	
�۶l�8���ޖ3aĵ���a4lT�F�%�)4�,���&ǌ��H2�d]��M�ж7&&�Η*�k�7݅�V�$�Y�	����#\�HB�m�H˹��V]��ֶʭ�m0�-�$wH��#I�y#�Y��4��m�jR���ݐљ�B�[mmV陿H�y�ͺ^�.�vh;kp�m�j����F��v�IZmz�Ču�m#krV���)i�F�-biK���	$��-&�Iea2�Kk��[-L6i#�����
2�ޙ^�41&�d��s�me�4%��6gUQ���3\]h�k��lK.d�Mbۍ��M����$��&�ɰ�Y6��Q;���k���l�V�Mf������Y`��iٚE� �K��m�         l���^�6��3��#��1}7��R�'	�YH��"�������p�/�p�ɢ�]ßq�͇υ^U^u4��\�猱Ұ���\*v�=�u���}�8���VC<�ߞ�\��Wl;�/�u,j���9+D�Ho7���&���튻�|��j'�!Vz �0wD��$r��~[���kb�5��Ns{��+�� ���f%�C�Z$�3�5��|�d�LtgB�5�f�p�w���	��|&A��l��i�udH�B�s��ܜ�7\}�;^�F}�61�����-�a�h�)o��!�L��S�8jw�n��Kmn)�9���D�G��6����4.�nX*�U�0g1BĴ��*kT,0[�i��λ'.�b�'���T�Z'w�ۢ�W~>�nU\t�bV���}����ɍS}��a��7n���'z��䣩Զ�\��][)!�o��q���lJ]u��]�<���"<Tܥ�ks>q&�7�ތڨis�oi�g+Ȩ�b'��cs��R�7b�r����H��5C�ӆj��bEw	�(ul��,�����(
���L7P�g��&��\��z4�گ�;��ЙN>����HR�O8N�`��&�ʹ�:�G�����6B�Ҁ�/��(���A9�o�y�p�t��!C�P��B'}�kj����"36���LwH�A�-��~�O�, WtZ����k��>�Snz�K�\.~ذ:�>us��r8\����K-ue.v���Km�p�	^�=}v��b\5�H������a���1�XL����鄊��*h:`e?`%�˿v�k��؜��K>&� �UZ8���L�NTy	�Ձ�]NU�dz��ĭ^lyV�[�-�_&*��N����ٽ;C��7q�p?��q����{�޼��A�tMe{u�t4/D)k����M
!���Dݕg�w)�Q5�7k]�2�gH�~��}Uj�i��m�EV�pť�)�T����W�d��Q�NvA9�',o\���i�[UX�ٵ�>�iF��\����#��k�C�|��L=N��	�˾ۮ��"�>�K�댪��U���<ᑔ2�H�;#�э�ġΎ�7w*F��ˀd8���+'g���:�|7ϔ.ܯ�Sl-)�
�0���]_z))]�K�g홣�JoI�cy��
^_i��I���98��9����ѫ^�b_���q��Tu���3BoĄ
��9�g�i�pU�]ǘ��{q4�K�T�f������ �i��]ր�כfDke�IM>��T�ޫ7I�wY1El��'ϧh�J�jc|��T*8�ޤ����?K~�J6��!���H��C�^�su �Y��^�_{��&('�~�i�i\4g.�&�9�6��/y^��gj�G��ʊ��&~��~�S�Fߜ4��n�5O�Ί�Qn=p8��jrg-�[Yʹꗾ�CS ���2�c5��Ƽub�mW�N��G9R��������;���B����{k�:;ǰ,T�<��p��7�!/���z�v�ݨ��X�t$�{emf;9�XP�d���'�օ������}�"�d��j�-����X���R/�t:}Z�۪�Uu�#O�6T�d���(e�5��GI����n�BXb^���\�AV��wl��$��j��9��\ݍ]W���(�����Sv�Ԑ�v;�!�cm��5*�W tv�; 2.��<A�F�^++������O\ޟ9���!� 33�U��ʶ�\�)��ax�o�J���e1��L�}黓�g�V�];�(}ބ��u~ĸ�4)l����+��"��Y�R.gJ���]Y�_/�SZ�7��bv0���е����������>��9��vOz*kO����$RM˹5��=ib������;����+J�zDm-�<�=���8�T0��`��L�&�'�WYSn=�PkSVzf^Gv�P�z*N���ݩgٙ^��37�u4�y-� �������d�L]))5l�1�1�l��?�o4��kj���LɪWϝN���m'��6a��;�`O����SwkC�M%�����y�	h��ϓ����B^��ᆷv&�g�>�S�Ķ$�(1���W����Dg�^�W[ۜ�WQ5C���.�Ö�ƴ_'pԏ�%���m/��}�|��zl\���� ��z�3֦݃#�N#�#��}�FO��fZg`�=����u�S8-��\f���5ʾ��4��t^zTlW�MǮ�,{?S���ظ�\�ڲ!�����2�M�F��o�Z�`��5M���\��z1�W5O��P����7�3�$z��L�������u����U۵��Mp��k0!����v��K��VȶU��+�
ۨ����F��˸��U��Ox��\:�j!��ʊ��A1ݺ)�����h��}u@���.��<(��[))�,���#H�g3;I�[���[&�+.U�O��Y��"D��R�b9��(�]Wz�ƍ��Q��0��ij��$�8d��FHVqa��R�lȄ�a"�m��6X.6��/ޚ5�?�!���ț��|��^�&�ɹW��t|��Z����ۭ;����N�S"�w� ���2����lh�"��#^�����u�u�Ak6��럠�\M��*�U���l���,,��2�wt[�!�z�ܒ�i���}+��͠h�'�a��mW���O�3ުrD�4�?T>�h���0	��;��^/)xu��P�M'��ȠI�ApB(`���̛�,�����K_��<�Ci����YY}HOfUԺ��Ţo�y>����3�s�)h��!=I{[�s���T�$_G�#\!�ٌ�s}}�U�j����F�?"7+�A�NpF�hdW�ݥ͉���G�	��ذ;g���!u�5��C�k��������y���/K�\w٢VZKv��L[�s��/e{�m��Xq��[<=g,��8��5~�����P�R6��y�~5妾0��[f��������|���2|7�ju�{�#����{�W�|�k�9>=*�I�����3���hÞ9ڮ����Y��'J�{4 ;���"�(ޒ� �^�6��O&�]�(�">�n�5��߯�޳$��LC��s�S��l�[1���d>鮓T�wO;��ރ:��棩;�+)�Q�죒�������fQ��A�:�=���Lʶ2l�s�,X���w����f�2��@�j��4.��sb�ڷp̡�šS���n�FP�X��"��0��}�{��m��Pwpj�%�æ�����޶B�QR���=�J���|ʉԈ"+V��8aN���Fee4}G�j���;��N�/�,!k(i��o6�{��y(TɃ�eҶ�I����1&���|�Ξ-�Nm�/�ڠ�&��������T1�kE�e8M������g��.97�x�w�R��ʑ�)�q�+|�N%�Lm��a��E�zJ�4���p���,]�^�w�W�r=��c���6=�X��h>�=��R�%z�u�~�2dWB�S1N�}5R��@i_��㗻�n빽���]��*rm� �v�.iZsvd��
.y}��Q���M��d��̌���QPn�-l���Gy��8��
T+mF�y�[����_�2#����5OM���^1��@�_�w�1�	{�{bx�V\;��Wa����*�n|�K���Ҡ�r�<"C�01z�Vl����cnvNW|�O�^���z�f�-�_��>C���A���K��u���%���N��s3E`�d�g9:�f8�����e�'��3_�8g�}����}%�2�^��m���)\��b�P1nUmH��tP�>YZž���/�{��[���%%�^�n���LBZ���\8��GAs�/;zf�r*���o�y�K4�c}���p�I���a�"�*�6t-��<l������`uQ�uS�NY���&�7\�-n�6&havՒc�;��+�L��}`K[����ø_v��^�������X�$�EQKfظ��_~6�i�W��Ic�̝�ݹSi�JZ8?�}{��������6;��"��LES���7���	�'_��i��衛���8�>~��-����R`�q��킜��;�Rl@>�NO۠m�'A�F�v��5T��645��fA���@���zVcmCVEwI�Q����s�Nڼ���f�(j|&�x*w�� ������ނl�cf <�����=�}�V���&����%e�>l�N��g���L6*V�$��A
!fa!�At��{x�}Dԗq����b����������0�Q�<?Z�=ǔ�`�C�	LU
��+W�vUs�M�$�s[Ч�c�V�W��A�.�����kQ�up3���;���>��uF��'�'Y�Q��E�W�V���?��ai�^)2z�P�c�#cr��^����-W����obEbdyw�U��?��g��F�$3���g�(�s��ޫ�"�E7��}Xߴul��\6J���cq$�,�G&90�#r	W�����0��zO$F����4 C�?$}woE�쨾>�ҽ�w}cȠ~�f�f�4���k��y���v���ot�[lMX>��m\�U���NQc���]zr��cƻ'���g����ˆT� �]W�GL��@��5��5I� �
K+{�������;����ѳ��)~��Y3j�����ɫ���_�T����u-�\e��x6��n�Z�B]<y�R�*!�H@wV�7�1G�����e��뺷���C�o*ww�F9b�v�����O�yD.�s�U�͹˥�53�;����CT����-Itt."�5X����r6>ER�d�vQ��PN��i��O���Z��r|)r~ٷC)��9Kv�E��\�1�h��eNӠ�Ϧ����Gv9�A���W�%d���6�3B��^VˇЗ�a}�J�/��V��*�{K��f��K�=.��6r�Oa�2��se�I��.���r����2����5S^�֏�a���n���;���Fe��=90�$��|,g��I�YR�%F�/�g�4�	���]םCե��m�Y�0qׂf*֡�wLn���3���ʗ߇�F����k�.�ͯD��]�c��'H~��&���=�߁i���M][^r�=�'�*��U�7R]���W:�9r��H��{���3^���6�N��XYp���'��n��0\���E@�O}+N�s��Nk{ި�������^�:P�xq�٦*�>�Bw]{N�9 �|�Ify<�;���v��׼rU��{��������í��}>��H7b�wH]������_:)�� �����@��[:֚�i����#����6�b�}�)^��[�>���fڽ	Foɚ0㣝̘.�ǻ����^7������FR�퐖���z��N�\�\�t{R|�Xtj�]8�ʉ���S�7���׍���c���D[#t:� � ;Y1����k.,4M$���]��4��A�Q1m �n��Q�
����n�]H%�+[��m2W[xWj�FوF���U���K�f1�-HdbD�ݛl褅���L�ȱɗKv.靤��Z�ΐ����5�j�2CBT���'d�$�A�H����uu�OÅuB��/�Zzښ�,�ۣr����v�$1EuL?eӘ���x�[��% ��u�Ѿ�UQb��^FX	l7	J�$4�!����Ei�'��Q�^�*�<�Ӊ��e���?��vT�נ��v	�(���y=��������aո$O$��r�s!h,�w�>�}��+^�n)� '���<����&��Jɺ|������a3�/z�B�~c��'ʟ��U}�+eLa'	�����w�f��=�ѱ,V�S��[�i��z�pE�E�5aË�o�=ԃ"���+>C^Q�T|�g3W�V��g^�2ci�w�E씓��S�U�tW��������DV�g'G�#=]��yR*7����fg4�P�Th��>�aW�u��ZvJ�4]�����hM����kR�)��྿Q>4�B�����(�:4�w�;�7S	�Ұ�Z����9�2\#��E��k5,�!i�����+�6�b}��)5z�4�
h��7�gJ�6a0=�6�z?$}��\�:nz��Y�r�u���F/f'�й ����6���A�}�Y�\_�+�t�ԇ����[��<�}Il˒�8�,�:�ĭ�������pfv��:�]5�3��+*�2�@�`�ٽn�*E�2rxC)<�4��ck���*���L���v�u��gf5!�V1�����ن7�`ݗ��XV����0��50܌��%��Y��<s{3F�y��Yޔ�f�̎=�A�����?��u�z�)}��:�a�i�pЁ�@�I,ל<M�)3Q�#�6�B��2˄Pp�M����(�~��h� �ھ�"�3~K�q����˟�H�EǗ^�,n���;+�~�yR�
�Zu�=���K'�GU���4�M�Q�iv���T�!݊G�9(
5��qa�A[V�H���,l	BU�+���B~�ToY髽�7uʫ�V(��	��f8d�wޘ5�q��K����C��	����a!���|��`'�w.K��t�R%%��'�M{}�x~����羳)�Y�o�Z��k;Q<�
,c��f<~5ߙj]���.��A�r�#�<"��CnG�u��OE�s�5܌�YO��q�j��<w�1���#
�P��u��]��'������D�b;��#�~f���]Ǌ��>3Iɚ�,��PB�N�<���O[g&��z�4��ǌ����4U�2��9�s`W��)��*�0�m��%�H�d�v����'��2_�9Q�H�e	��4"�b	-�9���~~��v�:[���AN�Z�ΐR1=�*�AI����i�=�^]����v�_�v��8Q�J������y5<x��/i(6�8_㟟@��3��6+�`.��n
��qSA΢��<�ݒ����G���Tl�e���s��u07Ύ�&��GWBu���L��þ���r��^�3��BS?>#_���������3�|��y�\�P@�яma�ݯ������[���~��i��G};seƌ��s������[9� M����3faFO�'ݸ޿:Հ��7�wU�?-u+�}P�m�T*��>_g�\a$��o.�����+6`�����'N�}y�W�Ep~�͡7���UC>ȟ�$��}]<�����W����d)��j;����}�i��jT~���3��� ��~��CG��7���H��e���8��i�������.�e�����wEy�氵C� J4����5ީ�r3���\��a�Y�iǙB=�����ю6vfP��
N��vMbS���V�u�Y����J��qmQ���S�v)�j��$��Hkm0˫k4��@a�3\V�Þ�ҁ<�앑j��g�a�K�_%��ۓ�y���U,�'���@%�K�ly��'���<Vh^٠~��z���2A Y��|["�t����Ȼ���;�*n�h��"�lP�|��r�\�� ����A�'�Tw���z�&T�si_�)q{FU��7	�7�?��V�I؝:^R�I�ܶT��r�u�V@��V���:�R���F��	��n[�r�?��]8�av�s�m�ǦJ�jsA�鲛�AuK�l=�h=���V���2�� � �y�c�㾭��9��Y�A�O��[V+�ف2�ˤ�f�orˆ?-[R�F��OWw*�G 3;�L�Rhm�_
6DT�u)��r���ˌ�`wՒ�hv:�)	Ќ�Ϋ�؋��n�{�19��N�Qs0n����9�Q7+T�/���Fa����I���eÃ�S�FA*E�Y�'�4���&��^m�R����Ѭ��n� �c�ik̸(���F��zo��C&�ϞZԴ��:�UDb����m��з�l�[�E�ӽG^�[����5t����r�㸶Յ��^⼒�b���'|������W��Aё�t��O��XIS�H��9g"�M�Y��B'q��[�0�61bt!m	�m�0e�}��@�o
o���];XK˘�H��M<��i#\��k� ��f��3R���;.1p�6MU]���cx	
�s;V��N���}ok/6�U�f�c��-@��&-w�-����2�Um��s-ꖫA�|%�L��Q#�혳�o'�wwh�P��!���qZo�
C���j�N���N��7@�������p]iP�����ԗ�mf����l�:�I�}�8��K����#K�m*��x�:Z���\�h;��� ���TՕ�c��3�0���.�4{jb��%��3Wtv�ؼ7H�ED�[`�O�m���UMg���G�^~�eW��pj��<qCs��Zz�֢�l2��S��TOac{G0��{��r9�k4��o�׳��`�4���qw(�x@�ts��?Y�Yj_Hq`���D��:���ٍ�Q��������gnc�w��t��B�c��SwhT��yy q<���m����5�ls�Mt�Rδ��Y�ȗ�.i��o4z��=�sǴ%V�]Ӫʵ��j���K"z���lN:���]d���h;��}����eˏ�0�7y)���޾itͧZ�u,i\��7�zp�W,rӭ�&vQ���ﾏ�/&ϱ(Z�)����e�G�r#9��9��q�n0G)]��rtw�`�T�2k���.Rj4��'�7��5�bΎ��z�d}H����#Q��v�J�'�M|-���� 0��:T���Y��K���ꡚ��/~]�5�����ܢ�*�v+�<sΗ�.��d�*,��y7�[�e
�h�p�G���|56���n/S:���ɔj׷�2`��O#ʇ+�\��l
�T
l�xu1߃c�xg��f����r��YB|$���T:V/�e�=��2��t��_q%�f��1��}[����d�>o!�ص+"hĺ��4�-4P��<�y�6�g���Û�S���g�֜���ųQ��x��}}B�P�e���@��ьtg����\3=�E�!�0u�x���f�=��� zG^����dw����{����W�l@��w3��~	Fw�M?�-F	�c��餦�!S��+��p�����M�/�1�ڂ�3�X�_��N�.�^�JQ��[B�W�b4�����_z%z�LD�{30�ǝ>����]JXŽ�ač&�&/�>শ�Y�r�z��R�2pw,��m��	K��I-jW����˦8P��;��u:[ٕ��\�w�9���ԟ�p���<v:]�xS���z
s%ɹ��8-U��Q�!B�(��A1�˵ͳ[(�]qM��6c1Mgd�Hm,iMJ]Kp���qm�CAųX�M�/NY��d-us�dؑ3&^��B٨�M(�Dkq�ٹlF\�m$��lu]�x^u#��5�sƴ����ᾊ�t�V+�J� Y�?H���<׎1��O�� �7�S�B�ʃJ���������I�ꭟҕ��)�F�}��G����o�Оe+#��v�k��t��>��4���>j��vX��c�7v�p�����0BoO�8�V��ȓy��h{=���l2ZgG��F�4�_�_{u��w������D�2��}�H�v7o�3=uV�C�.<`�{��2�u^��>a����de�AԈQ��}ȔF�,A��1�|\��FK��	�3���SUb��Fc�`���Y���9��T��2�]ȃ��b �ʊ*���T���;��љ;U~�s��ڽ��2)�ײ&LT�_Z&*�5�ӹ��Ɵ���3{�z�KC�j>��t�.~����Ԑ)�b+3��*7Q��M]r7�iȽ��"�;'3ڇ���$k(�s�suc^�V���v���$��z�8���^���4@b<)����NȵX�-�k�z�h�F��sZ���;]������aԯӤe��U*��R��C��`#]Y��	���1�Di%![�k�gj��kCajA�N�(Иwꓚ�z(�k���7���/h�&��j����Nv���i
l�z�L��^���V�k�3���K�Qbt{�! A�_T+�x�܈5J����sl������z����,�`��2����u��;�hɁ��t0�t�V�X�}�ݺ*�ԅw\zF�>��/��η�Y��!��жz51؅n���g�n���_��aT��ݛ��l�t�����ea�T�Zɑ�&/j��B�y��&��y�Iʒ�<����E̩y�j:z��EH���M������b�^}J#�۽ʦ8���<���j:2�O�c�v�.]O�/nR2�5�U�G��>O�u��w�⣤qZ7}5RЃ�.0�G-�Ƕ��2aVv!4������/�{�2uO�y�x�������X�P�>�,}�w��׳���ה�����k�f~:�G���g�������aݡ�:U<���*:�ܺ�Y���q��ϝ��x����!��ͻ�0-��A�?-𽡥�mڕC�C��%�?�8"%j�l+�[t7m�,���ֿO��܍����28W�y����/�"M]Z���,�M��7o���Gr��^7� c�c���N
^m�v��hI:�Y{֧c��6�Y���)��,�ա"���/"D�ak�3��;�ib�s\�V��:r&���\�5|x��(�Ճ"J��;� $�鸚�}�졫=��(W��Iq��v�D��f��U�,s������p���:�������`�[TH�ld�Ppi����lS�͇=S/@"�#����l�k���#���Z�\^OZ���CM��㵸Ue(�������A����x�Y�����TeF��XQ���K�^��a��^��z�\��?�Ký��1^��,�^�N^�"�h�#{���Şرc��G��ˣs��[;��3�q��묂_ In����u��[���Vg�������)��Jم=��Ï���f�
,�{[�b��D3���6w�ǯV�SB�	�o�}�q��x�J��`�ťG��a6��
���c���Y�Ar��f^*�F�/���a�r2�1��h�&chD�.����[
�߿.��g�^�wX����%��̆-ZU����&�V�^���2�u;�w��S<HC<�_�S����3b4d7_x�U�V�>9^_f����4~N��d�	7�KO��������!��*��n&6�\��ű �6ݸZTy�(����z=�����Cq���#�f����}���t��U�J<�# ��뛮��e+�7q������2�kJ5�D��/+kik�՛c��c*�l݅=�3���Ү���=R5jj�nG�2ǻ&s���wˢ�:%�9ө�1��G����'t�&ag��rc u�6`7���q5�xɥ�x}hފܼR��;]h�Y��[��YC�Ibr�=�}��\��`K���N�{�c����kMmU�M'�����M����j'�����ّ�{��x�4�����"ޯ�X+�������J�m�h�r	���4���;�**�c�2������Ջ����{����F�텚F���ba1���LOĴ��<�wm�A�~ʸ�7�ף�r/�,�m�
�� g�����#]�omd�Б���u8�����!��˕d���dmgQ�����8�#��>k����)�r&H7�'-�RP7�g��3��W*q5шO���v�B��9EFQ��(ϲ������m���;�����v�J�1�'�kt\'ޅ�R���m�\EU3�n��6(:�r���vz+�L��F�/AN�D�n ��i�W["���	o���L��û�q약S'5�����ܥ`pf�ܬ3�Kv��p˪�E�v9�cq��g(m
B�$�sެ��6
է����2���{��^o�a��e���R��һ*C�d=�kv��H]r4~x��*�D�7l8���:}����#�D�9��2�[]v�+b�Y��tm�%ْ�bh��͍-˒H#�%[f�&V�\D���5�]I�97F3.�M��f�Y�A�yuJW'�ʘ�{�9n/��%Ñ{5���+���ʡ�-��	�]��9�U�����+����>��a i׿��IJM������7�y�H�d?3@c\�2����v���{z\!w=�	?/��:���)F�t�ٟc�KzG>4�d�l3����A2���d�t�l��ĳY���(�M���VH���3�W�&kK�� 侤N�8w��ꝣY�̋};̴�t;U������xB�U~�8;\V[Я�N�)����D/N���f��f�p��$y,�+�)N��<�I�l���	�{��}-E�FŮ9�0c�����<�gw�F���rB�ہV��M���\���.[7��^E��r��ÕཔN#�sݜ���5��r���22w���ց��g�_VTŧ�<+�Lt��^�*�����͜w{�:\�;�����\���Н�{�R�_LC�iϫO��o SB���"Ǽ��dl��dh�7��oV�g�A)�e�·��a�Zqlg	8�K�.׆~�ݾ��h�S��M�~U�EQ�D;f|��+����&��n5ٟ��\7�m�����[�����I8���yV�2J=_.s�b[�������)f�qΩٓWG�������c��g�4?e�p|�^��=IcӠ_��c�{K�(KY�Sh��?,22a@�
q�#+��PV+�7��tɬlT�F��J�5�u�9-�n�Es&*�N��Eδt	���}Fd�k���V�;^�QYZ�=�Bq�{o`�� ���\|�|{�����:�kc�U����B
T����pqױbs�i��,ϬOI�r��S�T���ܠܱOw�f}�j�e�8*����w[�k�і7ڡ*�1�:.��΃g<?���O�|�/~���H���~͆<����/Q0H��wg��0w��;��>��;�j����c���n���i��:���͢U]�jI�77ֻ��b*n�d�;���논�Ũ���܃��N��!��J����=��Э�;�1��ќ��m��Om;�t(����]�,<����xၑ���r�{�_]e!���mT�"�W�
�x7�bu�(�̹2Z�0�w����R����Re���[!�4����M4[,��,���80�'oݩt����kW�Z�:����a����u.�?Pzr��;�vDYa���y�ۻrKX�#2A�yOt���qZk��zr��q�����ՙK��0͇�'ua�	:�B�qOM-����Q�:��xz1���(t�Q�X:+���
cwdn�JSJ=G���=^2�!qS�����_:9.
n�L(́K�n��;���{pFO�Ό�ݹx�`�1Y��UUSb��(�~�n�TF[uJ��w]���E�A����|}�PH��a�8�[����
��j]���{Y^��_�cj����|�~��8���x;�Cr�_n`�v�t�@ľA���b��פ,��l\��kP��P��8����� V��< ��v���Q]�=��5���ǣs�fq�|�|�=�U����\�dq��� ;��L��<f�Q��끾XkW��ǏBuY��\hI1�=
���s���QN��~�=�����I|Q����8}wE��v������ɻ8�m2�l��KSb2�`��&:����OV�sz�1�����q��D��_�T͊��6�ne*�S�gY�Y�>����X��?^w\�F�CT��P$�,��V��M�^^��젙} ;�sZ�n��Y��.�y�gV¸��Ֆk�TF׎�� ��23������6O�������Jz]w;�(��
���ET�t�rowd����ض���Se.����ҡ�k��R���tUus�Z�{���,��{0Ǵ�y�k��ga+��@�����dc+/DQ�OpB���h�V � WnnѨ��9@��2L�m+!Z�����>�N�ӝ�ɧ�y�Uʘj���x����E8��3�|=����={j���[�@{�{~�.%ds�ܮ�n5��
0�t��cc�R�Njz���ԉ;���"�c�7EY�Z��lZ����g7��Xk�ժ(�Id��HA�d-��,���Փ^��=1vʬ���yITJ�=��~���&���^8@S������L���)x�k��i��O*��,��Z9�K��W6�<���0U.�t�p-ğxϐ��+g�r�E]���X��z�/���8�d�@�er�o[�݃
~�ӻk�1����"�{Ɓ��5W��t�4`�"o����E��dc��٭7f֍�O���9�����{Дz�|t�l�{ت.k�<V
v�{9�wO��/�1�*XjN
~�׻��KP�����y>��+)T�&3ƪ�p���|�@lQ۹RU�-{z/EJ��^c�l"yX���蹏�{�Y�9�������"�$�D��/�:��*����]-=��X�����HOh�����c��K�c�נv�=�T(I���m�	��]`ԫ��'E0��r
�z5~x
���2r��nsʱI��T.t��/�D5}U0����-�νt�l+q;/iL�&�4ӫ[q��\Kю�K6�G6���s�J,H�̹��H�2ڲH�ؒ7m{4wG�l�c�4t�bm�	�$�b���mR�<9K�TZ�YC��>�͠D]���
�}�:��O�k�SŦ���sչR4F��~{F���櫹�F� �0h�i�[ꆫ�B�1{z{�z�:���l3���v'�C�2ffo��/}�{V���6�P�����`�R9³C�Qy��
�9!|�.)����B�H��1Ȋ$Di��K��x�G����w��tn�v\��lG�����S%R�s��#Sf&&��x�锯��7�mQ���d��3��x!Z�Y�m��3���O�P�+�=���D�)ɉ��3��!SD�'��{����)v�;�?���߆� ){_�/W�"�]}gd&��g���Y͎;
���mO�G�vv����=�*ߠmǎ\�Ìu�v|����͚�X��@-8db;��b��(����@*��4-m���b�w%\H��� �<e׏��n��uy�\蹾�3��+��S}��۸SS�6����{�L��+�|=Al�W���/����@�{���G������<��ݻ�r
e��2l��t$)̮͋^Im.歙B&'"��f�1������.���mu�Mͼ[w&�v1@��ӫiw�]����,�5��ʵܡ�f���r\�7h��Ю(:4u���dCL6��ཀྵm��;2�Բ�Tw��w���qƶM'$uv�r�����u0���,�u��WNg*>i�Ƿ�����k���*���`��?>ΧA|hj=t5�n3�s,�^����m��Tl�� qYv�)��"J݇�Û;F�@|�'�҇�Q�WsT_W9>�w3e��Ý�yi�3�o�-���փ&n���MhT4�Xʒ�:�$-uN�G
C�m���ja��o;����.<� W%忾��~��B���f�/3�R�ra\��UT�25��ր�+�i���?~�~E�t �F��QN�}���wǃ�<w������|��}�@>Y��Z����A8/+WuԜ��QK��N�ӝ�ƴ٢�n��;�X�B�5��PA�����9)q�G�GX)�4�ʂdP������ԟ���a� ����8~�B�~����~Ó�S��5C��5�y [-3�\��9�YV�1k%���*auB}-��Ji�g����`a�bV�*��F8R��y���4@�j'���]JZ��kg� k�]������}e�͋��$�Zx��㧟�g�'����j@�ޠڀ����"m}�<Hм�\���
䣄庎.�}e�Y��꤮���wMbR�3�jm75g.Q�t�g2��`��&3nEl��!m��D���i*f�{u��غu�ޥ*�F�����-�Q˶,ڗr���LG%��yJc���,��#����������W!%��Z\M	��Fy��H&tP�;����3f)�t�h��Q�Is\��~vW�p�#���H �)$�B@	 � UA���w�K3&y|͒n��*�wX�z$�o^���u�}T�\�p�r^�7�W/���WB���P>�Y�}��y�]���Ջ�$3],gw�f��u[NꨕW0�BCs�����^T�r~����2�ҚQ᫙���r=�֖4��(\����Ӑֲ��9Gjg󮇩\N����l[/��z�u��ͬ�/��o\N���{����s�������1zGpUlн#JR�,{��թ�͍k@A�!]��hb��r��1���U�5��l�:$����6�_��ɴ	�X%��%)b5:[Pҿ��`�W6y+�e�J�W����J��Y�U&��e4�gLG�����'����[�ЅĚ��i����#�$6��	���\���G[����<?'��R�I����ynk+�Z�3��<��:���+"��$���7�(��x&̗,+b�a������P�m!I���LA	t�w�j��;f7�U��Dk��-#:*Z�6ٍ�I�i�J���MX����H�,��8dp�L�����$�ȲaLU�`ζcjհҴ�U�u�s��Md�넬݉��U������V�e�#����2���lqM&��f�Ë�K{]�e%�f�t�[X�Hf�Ru���v�l�9��S����fK��j��ڷ1��[]y�$5�f�ef�0�0�K&���q-HԗRkd�L�UB�CcZ�4�7��H�wk$��3G����5�H�#t+����d5�i4�le\/<Ԗ�dk����&#4F]e���&ԑ��h�bZC��I��eJ���U5QJ            
;gx^�Eq�S��aKi1|�T�����5�-�'��)�N���.2�@�c�T���ݳ�3]���z����8(������rhJ\̍��}�w��p�Ĕ}�|���{����L���B�>��f���㫸�N:�g�~,������]]E�kjxd7/�э���!��cho����nm��R�\"���h�����e!�,���I�y�k��1T��̨�P���x���3�K���`TlYc�y���ޘE��߻��"���E�Y�����Z��츗v=�.��SL!o[�=w�-Q}uc}�$sY���q��f�.��|�򖟂�P鼻5�꾍P=��h\�u#����QR��O�ʼ��BA�9w�� ʄ�E�Wu�*3W��b�ê/�;ȉ�P|�P�n:���̝Ɣ��H'���MA�>�]���6js!z)t\�>��Gb�+l^X�a�c�tG�dz�[��}*�B���������ؽ�;�S�H�Zi��k�����C�={Y��Q��{HZv�^{����g��]_��u>�Ę[^6\c���T��*���@8+Pq1�����5,F'�Ϸ��I�+���s��M �t{e���ķ����嘟�-�ɞ�O��N!z�q�=836f-���R�{��}��ٝ5Š�w�sL�������ka�	�mN��7fӸ3,߬�$��***��\��4dr����L޼wՇc�;o��$�l\�sZ]Nbf��>3+G�׃�8WPsΝ�Iut�q�a�Q�Z_
��4�jdQ�]�����6)���&_1G5n�,;@6̽��>>�c�%�<wr��㏸���__{�E��բbc��.qp79K�b��Bn(���D�W8�z3�{�p���A/�zƽ���	.�ez��RE@�Vy!���M�)�'}��ܕ_Tu�*0��K�7*k��{��W��K���/M��?����i�߽I��Ȫ�:s�h~��{1z�4^��tɻ��du��,��$H��7�K=�q�WQODn��V��XW{�cPphJ7������3݊��B���c~E�m�l�����;7�wv 4�ь����&���d������*���������@��C��.�~�k��^���_���ܝ��Ȩ�� ��B~�/�{D�ѷ�&%g+�rd˘�t���>��R��k!wd{���K�H3n:�l�B�ф{H0$r"=(h�N����o_4�7[�Z���}�xr`�ִ���V�7KR�d�7Wd�U2��'�P��|��zr�ܪZ�����;1�z�&>6�'�z��p���HM̚Ʈ��x�< <_$�j��\��V1b�/��¯�%B���sdʃ�ַ޽�~��u�W��д�>�{�(��Ѣ�k�����~�C���WD���p��5�ӛ0��j��%Y���ۯ�Jw�[��1�qT kCf
������q���wX�;�#��Ŕ��=�pN���-�ؤ�뵵1�͞`�����[�Wv/Y�O�81�v&��z<W���m��B!_�o�R��˵��|��.Tz@�z�~��F�Cɀ��^���|�t�"�eoH���.�>�oW�O�ҭ��4�m$���#�(A�Suhp@�q���!PLNԣU3���-��̀����
��*fl�߮v��+a���xg��jv������n��+g�g:�ѯ��V1��5p�~5�����dq}�&&��b�uJ�W��Z��&`\-�O���^�)r�\ouXG�cv�J�K� =ɬ��`laG:9T�iU�nXjϰ���}tcPɎ��7�D������Ƅ���{C����ΜNV۵�w�h�;�t�-&�%6`����Mtf�׽�H�}�k�f�wq0֪ڒ�N�qu�C�ڝus�{�����k65�o	��
vڥ]}�LlD<1qE�r��h��>����M4�G��.�#�i���y��gd��] �;�q��b:��RX�BhZ�Ջ[���U���i��B�+��U���6]�������ab갏;��XU
*I$��ꐾ{}k�ͯ��ݏ�v �&ͱn8=�\t����<�ǯ��/31������ٻ���Ԍ�z�ùEж>˜���o���q|�;4=����cU6kO��S��蚆��Ȥdi΃~�#ǚ$L��w?xb��~�a���ު7��9;p|v���{�=��\Xh0��&�LV��6TM����x�<�;w>zz��>���d&V��{?	��_+6�,�|�6L��X��h����k�oFQ��r5ߊo��#���LVrjm� �����6g�xTU��iO�Sެ�>\;�2ŵ
;�����{pr�oMlp_u]ݽm�
���'�-Ȼ��΁�=W�ah}�5�&<$�ZbH�S[��j;l�F��'��x>�����_���suDӾ�y�ui�J�J5,[1s��a�m��#��Q..�6�U���ZU�|��h�p��O�\rzG�iuj��9��3�1ɶ��~�����WW��mDؠ"�КdW]oƆ~�ܮ�h:	���m��̾P���m��{o*܋E�ْ1�%��5�wJۛ��K�k�\њmu���(g=�]�������3&A��u}����>����w���%�zp����B���{�ڵy5����6,��;w�p�P�S�{t	G�0$9Q" �Hƚa��s�Ww�����ӫ����9!T�������D��F��h�].��?^��R����[U��9��҆�=�~UH����o��X���k��k� m���
�Mw��P�����y=|�eO��3�*��h� �v'9>�
�-rN�pQ��h�kg��}"�Yu^��X~����a�����V\�ō0�n&k2�}SqV��:�����$�,66r3�����|>�%�ڦ�%�:^���gijOh��&��?P���3��bc�����{�yV?h��B��e�������'����L��Ф����Н�i��2%=`(~F68�t�V��Z��3轛��Z5d��	���0>���2���Mr� �f�H�J`�z�C�����=E|g_,u���+I�(����@�)U�@Tm$X�&��G��ڶ�y!r�0��]|�?_$'�T���[����Q����+�e�ы���ln��e㐲��W�tf��G?n:��
$��º��&4�*T���ޘ��� ���]K���s{��e�>��ͳ��Zx��#�&I��e�ʘ�:�Eq�t�'�W_L��f����/c����P}=z7w�������J8LMz/'��@�%�kW��aw���V7�8GN�s�ʙŕ���B��Y{H~�k.i���W(��fX�2�_���x$� �<Rw�w/5�;cb�hcs������)�ٹ�s?�����5�>?�L��=�*��s#�"ǫ�]�GcH���Dz�JY��"d��:��:�n�_n�-9��c'� �f�# ��Y�w���������A(*��aZ4~��g/���m����iW�~�}Q8Z֏�<�Z��c�U����w���~��21�4�8\�}�0��&9���|�1�x+�=6к%�e�H���c5\۵t���i�������v��iO��{[�����#��<:n�嫵�39��M���>Ú�+|��:Gzؠg��{��ߗ8wlY���q��C�{4R���s�ɣM�չ^ojxnXV�Sts����VmY���X�#h?^��T��#�i�t�؂?^T�0ܖ�L�<͡�x�s�7"y�1��wP��A�/��f=�Y�G3I�9n�r�e��*a�U�߷�du�{ףWTm�g9�c{���C����p�L�r�ƞ�^�m�5��Y����kD�g*ћ����'-���<�a~阛�K���������($��^L��fO�E�y �v����O���;°d�ڃ��YJ4u�/v/�&j���%�2�LzR𜫚�6�87>�����f�]m�%�Rn|������y��Bݫ�u��,q�q{�_rڡ�����ĺ(�z�ԁ�ڹ-5�-n������d�%�M}u��f�����]_�`$�����zD��j�o���~b��q0Go��������l�E�t[����B(Zn�aJ���U�!�q�{�������J���;=ҧu��?
ۇ>�o�/L�*�ǌz�wgq8�.��.o�xS�.Lu~��w?w�@����y�]�����}I_��ķ<�#�E��Ot�쓭�ݓ';Q�d�/��;�+��.�^��EV�C9�jʹ���O`N׶:Eo͸��P�m�u��#�g���7�^!7=[/s�T�T(�!�p���[E�B�U��Zht��W<���8���H�G��w�L'����z1y�b}x����EvH�+9,N������s!���:N��m2�nN<wIf����fŌ�;eޙ�����X6�o�{��L��Bf��*��TM�
�lr�#��R��e#e�åf%���k�d��u��ZR�c�+uu5�&��K	U�fnp��u�N]{hI�V�f盫��Wn��H���m��{�'�-�Q]ۻ�Y[6���5�B�~���遲V?W=>w�w�(��7������Q�C��g���[��K#�p����wG۴�nF�T���dQ�I�7��^����]�r�.��߼��������� t��;�D잜7��P��6?�J�{��
�ƩQ5E��P�[�H�J ����E�=ԘDA��
Ǭ��yΥ���� {��M��*NǺU����8�25�!��=vr�F*/7\�}Q}E��c��&�$=O����ԏ�I��>��>�����׾�9�;�����.���&����w�a�=�Y#����wE #����0fdҕ�ү��G���n�؉m�}�O��2ǽ�M���7�7.�Nu�/?GvNid�ہ����u[k@Ν�b����RzR2�gݾ��+o�ȫ�w��w�k��y�w���� ��`7�BU�9��x�)y��y9��o�G0�>�=I��+��Y>��/�}1���n�)Ϻ�\�Ut�N�:�8���������{+4ai�/��|tcŃ[ě�8^L����у.C��M���v=ɫnة|E�ܵu9��Av�ZI��/�u�E�/�Z�ɻ���yц��uҨX�c�
���TZ�W$s2ˍ�zB̌m���ss�:��T�s��_ӝU�L	$�A6�$�0�6)�,��t�ߞ�Z^���=�b�������+�����i�o�ǒ��F�X7�f��>�2:{4OA�9l^.:O�d��O8���.�\V���.��3џL��a�tXt�g%ԒB��=�f(u�-{5Nq��Nq2E�;�Rg)w	r�Wݮ8k���qKOM�������c3���� #���>� DM�!�F�}������ڃ	i��!�J�l�E��3-������0X��.n��_]$)��t\�^��]A;���ws����FhM�{�h�ث�^��;���6j��i��/�L2{�nƱᾕXw4�˱s��Hs��T�Y�ʞr�mY����ex����p��]K����v�C6h"�������}%m�P�UYp�f
)|H��\,�՘V�_R����:w��Cb��d��em����+��{��b�Z*T:��V�	��x���	=�"oK%F+��M���Q
p';�*�ۥ��R��"=��D�k)&�{�8�ל�ڣ6M��]��8�S��wI���N�4��{�r����nްy�kZ�X�Y�}�$EOJ��+�r'�HbK��T�=j��������z	[�o��]Y���Ǐ���{w���G�_�3$t��Hv�MF�a��ܲ�4����>�Ez�D)龾��ۤ��tbo���|zlF�9�y���Қ�M��^�U�����q�bjoj��.���<�T吺%[��Ry�w�xŞ��r3�z����~bn��w��͆sI��q0zX̨W��Zk
\{�l\�:դ�����YG�W^3bgռ��9~��db��j\���O�9."�7�������ٱ�)�K���C���U�C`1��9�B��Z��Re6�0@B,8%@�&CL��
�sѻ�~*���:������;
k���t��F��=�$�8=�Y\P��[�ڷ\D�����Z��7q�g�N��}<�<Q��=�^���ݪ�:�U�����^��\I��f��=���>���PZ^���/hx��8��ﭪ�x}������$��q8͚��:c�;y�E�+'�z�\�4t�"p�!p�o4J���N7{�I:�e��Vh�>���s�C9�h��F��ۛ���ou�;_d�k��35*�_��5�7�c��F�](B<h��H��2[EZ���L�VF~�_;���e�r�Da��N�$�G5M��4��N����Tc�>����<>�!@�^�J��E"��W�Q����1��N�����h����d��W�e����{�Q��#���LL>��ڷ1lTrr+��TxQ��T��;�0�(�(�7�ʢ���me�\7Y��0��0�,�3i�dH�{*��$�Lޤʽӓ����Y���k���q��0(���q2��jF
�H��TE�Є,׹U���;�dYq��l$7��Dr {)��X���?}��Vo
r���E�c�&s��o��ug@���-����G��})jmJ�r��ǂ�RS�)�u�T/$���UI������	�=VH}}N��]g�6Q��N8�Y�MM&����}*u7���7�{��/��N��|� ?<q^�u�2��4�+��";q��*6p��Z����T"g
+��kF��y�o���<ڍI;h�x�#J	&�?�����̺�w o}�|�� b
�i�د߸1H��b��X7~+H���.� �*���|Ǜeʶ�/2�dC6�|^��.UK�*�wD�
5d����+\����-M����5��2�g2A���ݣ��b�]��Y�mѧ��5��S�Xn3A��r�똄mG[-QZ[��]���JgY(Rz�/-�T�j̰�t��FBwb�ͭ839��T橷g��˓��R��xo�+�ǕC����N�nv\2'OhwD�=��i�pYK-.N!��۴>l�M���I�ڣJ�g&�����o������f�Kڻ��.�׽}�*
lnF�T���szM8[������,���9.e� I[�v�Y[w�T�}J��/��4�Z\��95](��d(^�f��=yE<̛�G������ZD�EM=����3c�/;����g"��[m���O����Y��A<�8�G��3s������eh��V�ЛϺ��C�ŋ��7M���|�m���1s�Lt�e�FV��-��J6�I��򜓜f;jwUk���,��]s��q;N�j*�!q�Ⱥ�J��{RM|���ad�6%f�B�C4�=#c`� >�����y�w�����mm�&��#OT�H��p<���R��3�x֓��b���p������F�GmP����j��AG��Xc�|��w���[c�L,�t��D��3�i�g�j�O����é�;߮����/��C������;ӽӾ�P�W�.d�)��gh�:�ƥ��?޿y��w�.�/�����{��<�>�6�:�g˃|O�:�t2�!���.v�M���9� n�S]��v�})�]�^�d�����Ѷ�G��E�P���YI��M�F%����!�r������^ی>�0�DM�Q�zf�OC�܎��I���	��
�{�T�K�c�?~��V�%/��J���1�d�o��Pߪ�8��#c	��O��>;D�i��LQ����qsg�3g<�p�'��ُVX�K]1�����8�#��>�ɼ���|k�W�_�[Uc9^��U�\v��z�i�YY�ތ��D��9�����T�E�P��.�����"�ys*�J;.f��J���F��\�h�aЏ919�|�!<M�v�LsY������']W+�h[���BE�R�Ũa3��8r`�n�����+:x����BK�C�WΩF�Q��ta12�l�ۢF��l�O��1�g���*�v��YR�Te�VM�2ʪB�lf����%1tl��u��li�b�5��a��*VR�8^����(�@�d_1���t���^�;��G\:���߆n �����Ђ>�͏n�Z�J�=��4X����}�Ϙ�O�j��zwܗTÓ~���"�u�o�?#��!hhn�=�	맛{^�70��OVI��+��$��Sg.)F���Tt�B���k/ԑ�B��\4�C��O�&$a�2����M�͆��ס��26��F�o�W�mʝ���>�c�L�
���L���7:�����F�Z��O!������'���I�9*~�������=]�Յ��X�����B�5�ʍ�u���	�97造���u-g�e�7u��[�6A�c�-&w�zYVp<��W��]��`�A�S��c����i$w��D��]VO�@j&��W�z�c�M���Oݐ�uZ�LW�hA�|&<_73�e�ŖTI��v�A�!���c��5���s[��^}�j���h#��ߦ�g
Nb����I0�ٴ�
������F_�i����I�Ƒ}R|�-' �x�fs�nZg��R�IGz��m�R��yu�UҖ�:�|;�6����@���b\U� S��ov��jf�v�r�\�6H��3$�,�43gI^����J�+�m.��dz;l+��'��#Ӝ1_���#���t�˼,��M��q.(>n@KH�$Pɗ,b'�s���������w �Ǥ�(��W�םGѹ!+�����S�ҳM�O�����yC Q�껤�������� ��N�턓�@��~��U�Y��ޘ�g��(2s#�"�����0�A��W����Y������vש�Ǿ���v:��Q\�<��{3���y���=����jxRu�G�D�q�����ʿ�7(���K�9��Ͻ�e�E�:z.��ʭ�L�x���Wj��k^�w����!�^o�p��ۡ�4��H��y��t�뽠��P�J�S����/�6 ��t�H}�{=�>ʱ����8�̠_��v��P��n�V��A-��O��D�C����y�+�V�#Z�6�"�y#6Ԏ���uݥ,�2i��k*sKeAȘְ���ڝ\Lx���)��EU����G������}��U<{Cs�����lӋ���.�Me6�\�]�8*�s�T�w��J]���5c4Q�N�i+�a�k�ɒik�nu��fC���λ�q�l�"�ѷ����31<�twU
��Z;���[�jm���=��@����W�{[|U��{��퓤t\���ߣ㒾�z`�-ڣ;�l�F��z�fɱ����f�(���
�"�ɍ���ܛz�ڍ1���ԯ}x���87'`�*gw{��$�ɱ�yu���w��9�ןx=�>SOb����eL���܎���@`��I"��*ߺ�Z:>��fJ;ut{�W���P�a5�u��[�im�s�k0M��}S{�/J�q��n^Ʈ�[��9䀙r�|6�q+9*�"�������yN�݂�hG���Y��P>�V]�&)a�{�]>���0�a��q���6Eܧ����ný��%��	�RรfF��{�U|��6���֣s<>�J��� �t�mk��]���wLm������A�xC����B~.�� D������U3��9d0+��eXdڧ�����AR-�i�NT�cӻٹ��Bu��)��]9�8~ϹW���������z�g������3��@�}�`e��*���=s�/�?o� ��ZׂU����s��s���[���W<j���=�ۥ�����;i:�G�i.4fIn�gyX1w�N:vV�~έ��}ݷ�?qȤ]vx2��X]Jh�ާ�maPm�
�%Me�a��C6�-�!hv��2v�n8`�;�-���0*ʾ}օG�a��2k_H�$�q�B����e�[�^����Y���A�fTT��unDǷq�	�쪮;+��H���O�Y3��

_z�ŹT��A��k�o_�w��w<.��>ۙ{?h�N��⽴>�����Uz�Iu��b�>�[�Ϲ��j��²�+ ���P=4cG.�}�z�Qq�i��Pv�R�K(��)�#�E��q��]���(^ㄱCo��u���P:�lN�mX�:�S�^��Vv���h鵟	����9�3(�Y ��:�v-�k}�/K��X�x^���o��2���48R�[!N�$�v��!�O)13�62���73�o��I�37��:9D7��R_*��׉3v!p��y.D��J��#��u�~[�u���/���f��h��X�]^c΋ZQ�t:��ю`�8��׃�M�~�����\�K�����y��m$v$ąsW�fe�
��	r�c�9G�N�R���/���K�F�}i�*(#����RB�ݧ�-��P�Be0�v�೽��v;�f`�N��=Nc2�.���'q�K*�"�B�,B�s���M&s�1A����Q�<�iХ�i�[-�԰�b(��]�������e�C�x����њ-v�fM����mX�dJ:��$�c�X�1[��̠&�Q$ԅL�  t�2�7�N��M�G������"�='�Wdh�Y��"���1�}��/�E�Լ'ن��Z]u���1����3�{�?�׫���:�ʍ�S��*���g1x��'qF0�&��j�b�Y�OVY�p�[t�{˜$І�2s�|R��ʮ��f�Yˋ��o��(��G�k�c5�e�Z���+�7�
u�㦲sMǝ�і\����������n�`Z�k{�ϴ�>!�맗`� ��f���Eg�u����M�fks�Gz�'Ӿ�D���m�"�i�>�c�L�y�u�N��F/fڋ����ړ}�4v����5X2f����F3�531�z�b���;�T�6�0�㽗�X�0���ؠ���V��YHhZ�p�J[������=Y���S#�T�}sls3��N9�_m����3y��L������?��OSfW��O�~���Plq&��]�5Z|��I�yH��~�\@үy:Y�8���l�:����	���O���]b�+>���d��l����}�â�:�Y��sCϺ�>ʬ��ZZ؂�6�b���&�OG9�<�����WW���Z&�(u�sAܼ�O����(㮾�N�.�NZ%	���%���uK{x�{DS^~��m��GA�͍����t�ys�H����9������#���s%`Ԥ�n��ܮ�{�͉Px��";��#/��������}��CTp:^97k�%��x�!�ȝia�o�T*??{�j���X����]$k�bIo��x?��4r���;+Dd˳�)l����������rL�7�.p��Ь��'�z���w��O���~��\>�.�i@���ۣ<�!�_���b��Vr&g|0�j�2Y�qط�"�m����<���g�^`�}����]��~ ,��/L�ӭ��(��ؿZ+^��f��ܤ3�����%��axj�g�5t�� �^~�ԉ_nl-����ф��jz/{���.��ꛋ��&�]h�o�������Q�y)���@����rCq^W�V	c����j���Q@��a�@�$�PQ��	}!$� y؅���5�����h��ޯ#T`(�3���1��{J���j%��$����]�8�@>�XNZ8m�o�'���������TgV&%���5֎Π:7�^+�aѫt۩Wc�r����R��_$��d��a��XX��8P"�⧗������.���L^T}L�@����M|���kU�?V�ؾ���`��z�y��xU;�Ș���P#�$��\r��{�S�NN=�F0�\N�y�)����gcӻQ50��ʝ��$����=��Ɯ,��}�z�ϟ�!b���o���n��Z��Tҕ^���;��!z�Ӎ��z�Ȉ%�;O{���R�u�f	���w���g1���]}o��޻�a���ͮ騼�� ��27A�3o�t��G]�X�����LN��!�ﻁ����΃��mk��"��^�ɩ�B��F����J���QpzǼ ���zgfi'�k�8�e�u�-�oj�M�0��LM��a0�[BJ$�I��&�Gb�j���o;��7�B�y[��X�y�Ew�T=�c{��q��.YX�P���{f�n�i5���z�R1�����1۪r9q��r��U��I����(ǻw�D�ݘ���� ����S�b��k����f�=p+�;��O�F�����ږ�����L�Z+�eD�U��r�=x�zԎ��ڱ�Z�7o�o$S��BJ��C�
}:�v��Ț�u��,�0ɼa�{Av�R���Y���ʇ���$\�^�V�z��f�ܑ����L=&�xͬ$��^��S�����z�"����@�|�U���1��^��2����X<���ze�����:�3c�M�+n�5*gR��k�|-h��|bvcֆ���w=��Ԭ�]�ddéc�+Vk��_G�ԡ�Q�m൧�ip\��Im�X�B���q���U'z�F{��$,�י;��~�����8<����{�����.g	g�����mK����$�G�,���vsY���ҳ<8@pL��}+�:k^�=�r�y�2Cza�Vq#%�E9�ݭ
�d�}���j*LX���Q���)Ç�(
}�ڙ�WO��-�8j6�C��_����QV���yTG;7��?�-�
� �4�e�4�9y�0Z��Kݾ6�aׂ����s�[�źz��w����Vq�(N�iX�1�b<eq��w�J�7�Jn^٪3˔ |;��ٻ����Q?�o
�U�hzC�j�/��VB���fM���a���Uv��޼6p�*�W��R2Sz�h0���X�έ���V3R���n�#��.���;�z�GF���(i'Ŗ�d��&5S4��7ST��]ԝ1J��6�[v�"�6,RXk�v#X��h�I7JΘӭ1��+Yf�F�d��bGJ�[�f�	m���m�Y9��Ҏ���,��rI'���V�y�V��t��Q;����4�]ˍ��v��u�x���! �g#�p�+��yS[�武E��ț��t ��+E���jg��ta�+L�>O�7l�Ш���L"�O2���n�cV#���%W����R0�l\3O�SB�럐��Y�|�<a�� �I$�jR�E�NF:gG08	�19����1!��ѯ޻�e1�����vw}�����}s��X�ֵ����`�� ����wwWctë�πxq�"�C����j�a�ҸS�W�Ё�j�<x����#��'�Yٮ��(��½���V���s�9����@���ǁ���Y�Ш�G���F���Ɂ��-Hj�����)�י�y�W�ѹ�く�o~:.����ꌏ�>Bz�r����}G�.�������Bo��v߉޿B�7���}#`,�o��
;>6�.��B�;Y������3��%��5��~v�
�MR?Uf�֞�{�߰3�Еhl�Ù�(��=X�g��3�!����i��a�!S�L=[M��B*�k�X#Mre(�gI5�B�0>�贆���GP���2�yWВUj��Y�����◝كmU�]�| �9c����#/r?�r�|���w͚���[b3����}|��#b��]�r�lfz`�D�C��C�9t6H��!\�Ҥ�;wQ����#�l��؆�
ɷ�
�݅�f3T�L��3w�H*���EII�O�=��pp��Y�Xf��٣Q�G�ƌ�Ev4�W\Ǘ��/0v�[��٥��um��Z���]���.�T��cjNkO;��ڜM[�:Nj��;K��~������Hz����t�?'����y}������?-� ��Rd�ꈬ��l
w0T���'T:�#�K.���ۮ3���Ŕ������eI�0r�+��hZ(����A�&T��k{��]V�a�*�N���qY2im��v�{���{��̍]e{�^����S���ٌ���Rj꼨�m��+A�tS�QuG{G�����Wr�nmL��Cy��ifk[A]i��l�v��m�.�V�}�̶�;�3F���U�Y�9���f�#ya:Y��#�%���W��TǇ�~����\�Kl�`ս��P��x+ZK���0u��]1�V7]�U��P۽<�*���|1�6bX��dԦT7IT�H8N��5E(?���n#���h�L(l=���k�r\3���ar���=d�1x�a������oF���g~K]łGq�d�x��:oq\�pk*¦�rҡ�X}�dU��P�bo��V�^
%�&Iw#�%���@҅�T��
IUQ2PU  �L�H�w�?�������̛V��#�-��,�um�)�i�����6^�ףj��]B��5�q�`���K�yZ ���냅�ԵdC�(���*�"����2�s:k��6j��7���3�:�˿�����;\�wI��M]��7�o{�ujWvh3z/���,0J�ʱ�#���WE7ȝ���]�C���y�@��y��q�I���{I!s������uG-���uDa�v)Vo�Q����g�57L���͈n��c�GUL�9uY:Um�˸�Ge�Z�?7�I�&�3S��-j�a�!��P�1	0���f�����aէ�,B�i�%���=��6�p�ȖU�&�[-�JL(�D��8��U�ʾm"e���:�V�"��Bdu7%�iKa2�.�d�����M���n�BCu����T��-�I, �l�jci6v��ZF�����:�fZ�wJ�3`f�lS�d�	dh���h��,�e�c�����F"��������g�<.*�Mٔ�myt�szl�;i*�F�]WfM&��)EI�i��xU�:��eؚk)��9!����FD�Y�J9�Ў�ZČ�&�,���#���ml��`���$��7MqX�
J�����Yb":�*M8c#u�d�m�K�H�"E�m�Xݤ����٭���B%�i�d�d�H�:R#M�,[�e��픚�$�{���U���)JAl+\h�\���iz){%Eqq%\�;L�sn3t�`ؗsr����+1&uF9��j��e�%sJ������΋�]$��i����f5���-,�m��m��       ���d�V�uWY���.fv�p�-�mK�UN,�s�E�`kd�1���|�J�{�{.=݂��o<8���x.�:fj����w�q} �~ϞK�����ڡ��^�k�mc�9�y�Oe<�2Pm$�����p�|`���4Lͅ�qާ�g�F\oFH /��>�7y!�K/jml_H[>3Պt�(��cD�M�3*[	��$~���mjO��`�=�L`��UB�n�(V�nFh°p�+S�Eϊ�%��R��سeg�3כ�:�2�<���H;�5(h��춣k%�ؠG�.�qsBEJw^�{�D3�v��f��	� ��rh�k�j1[1a�_����*���ӭ�������'�t�����>����]m�
Fׯ�>nTl-��	�����i���=Y`y����^��ef�8g�Ά�i��?G]zJ��:T����^>5Ѷ���4Q�b�<�M�ۗ��'n��_<�̊��4v4�����K�g�}�ӯ�G�+���9E�@{����F?!o7��mo�(;�"D�S�Jw<�\[�'ԅ��R�Y�~�X�yэ�����}��cf$�ga����L.���+��y���W�T�=�IX�H����3�����i����n����Ul�v���]dɨ��'^y*�z�́)���C��lp��������zQ�ˮ2��&�l�-�eŽS]�d�a����§n.d�wG��"��(����\H�`�Щ��y�7�E�ws�_Z0���g-��=�����A�[�+���Ia{��J�j�?u��R �l�V��oA�Td�D��\U�BjL�X�����D��{���SG��Zc�����t�8}>g��wS9��ǣ^1Zh6
�̚�� �4:a$�?i�MH?lRޛ�}�;��10a�!׫k��
.�΢sc,�~.|��+�~���Lv�R��\�:G��{k�d7��`)zo|�MV���W����5���|�c�ɘW�'��7������(�d���]pavL6�8����p1g�O\�-l�c��Y�Ő��ӏ�����~5���2
����%*U��P��L7(X��h)lNx�h�M����X����v����CA�"����y�k�ɴ��U2�C�߁���d_��4nx~1��Ϯx%�������,~��
��w��5M�Y���QǦ��.��N�8筎��(L�A���Y��M(�T�����C����lras���o���F���;jV�Z�e�[�J�Y2.�u��l7}��vSn���gK��L�˻��WLja��=-9�)��:�Њ�HL]��qb�2��z���1gv�ŉ�o�_~��fz�3�^Y�ҵ{�nmMu�!��G�ڽ�׿p�/��Y����t�?Y����;D{/�^]?�r&��{=cg�*~"���u��FNS~_�aG�3^ϖz'd��G���k�[[��A��ͯwKY[��8���f1�յ�5e��@>�y��t����@s�oz.{�?NP�����t��mɩ:�r|#uǀ�@�$�7]�EeK l���N�[������}=��L�Q��$��r�l����N 1#���&ɯBڭ>������D�����/`��*��w�xo5��_�˼q��)�z��?]F@勽~�ܱOZ.w4n��s=P;���j��v�g�t���ø�j٫f��dsz��E�#V���ywO����_
K��=�-3�����M�L�T+��������kϵ��u�V�b���9/�Mۉǃ���������2���ՙqp��u��wY�3o�A��0��wW�+ײܾ-�+���Y귳CP�?'���y��-��9opl�!ә\���z�	;N�d o�n��(�G�SPٮѶ-���:�j�����B����}���1����i�Y���׮��
���S6Y{�X���O5�똓F�+����:]f�-.]K#)Q�Y%n28d��̺롉;K���& �9�鰪�Kl�S5�ZβMXZim�m��.`�y��S)n�:�#�������E��U��g�%��O�{��y�sE�i^V��0"�)a8��)Z���I���a]v���Փ�����zQ���R�m�F�4��O��og�i��г��C�:�j{�w�R�8�D��i�D��[�8v��F�L�AP����Ii��L�Px�(9�M]v䁤jF�S9��G�o���;��<�	뿶U�ʔ7<�HM��h߇�<z��+Y����ҫC8c��k�<��כ�;#\��si���SSz�\�㣩�ܯ���H��|~��^�TԼ(FOl�},?p��z��2�JWܘqZ[�۵`b���WV##�ΘY��]�]��B��-�ûB.&M��"�Sa�E)�G�=����+gU�4qP�.���ӍHt*��c%Dm�=�|u�2<xO���6#�~�~�������oǤu�x��b��0-�NY^��.*�#`�B�Vgt�]�wCbRqMmeP����[���/��Q_��\����Kv)��ϑ������1��k[_q����ʁ#�PG��Gs���mV��	S�K*��7-lxM���A���C0�'<yK�������� �}(��k*sUhx��Q�qRLs��s �T{?3���(���q_�w�o&�o�-����ܬM��:�Q��(%�#J	Q�L(B�^����)��v���eM�Xs�D�Zro ���u���������U�H�6�	��n�6�6Vl�ޘ�/�E�9S
z�<��ͅ��G/�1/����^�맋D=&��:��V��v���E��rDfeF��w�*#h�����ޣ�voA0k�1�ܪ㑓�uY��N\Hy�Q}*&���i���a9̟g��ռN�Z �db�������#Y}p��\�;�c�\e޲�R�黫a#3�^H�:^�xW��Of|��9���ݠ/eu NeARzF���W�עv}�?l�|[8�1�D�tLz:�H`���Y����<��et�P^D�{9k5+Ћ�(�C�~Z]xd�gr8H�ga���ޫ{���pH���^~�(�_��*$ �E��.|C!��MH[�B��;8����'=�=At�l�V�5��җM��ۥw�C��O�f����z���X�>�`���� ��gpc�uJ,�b|n4輝E�����ѣ�V ,��9g��s6�]4�݌�BF����4p����97nov��qoom[�^�C�My+��;���Fa2	���</F�����
۽є�ECI�P��\K�c�enw���z/�&`)�>;鞵�w'����>q�jf0�gp�n/F#	�2ǁ��/�f��pC�Y�q��]z2},єw���H��������|�l����|"3w ���2}�����ؔw=&;�D�fA�Sr �Je?����_����m9\�4�
w��喪s����+�'N�Զf����y��7�5���5���ͻ��6���R|tP�Wȅ���t�j�����r1q�( tǟ��}2�h�I�|�P�ݘ)0Y��,8N���8���CZ�~��D��CJH$����!M�eݨ�����ņ߼�?}�M�V���Ϸ$�=��%nN�(t�N^����ʐW��{7��aORԳ�?Ӵiu�E�=3�u���\�V	V;�W��z��1]쟰���_o^����.z�熳i��`/O���@�+��9ĭ)W*	��+�}CV�WX���߶�շ���{�D�RW���]U�K֝��ZoZh�!�tX��m>g{J��>�4d�]�-�Q>�n���oz:��'��Q��P��M:�8^X����=���������}��&aKB�h�}�r�r�IT�"&���a�p�O�� w�Z��(oH�a�s���W��x���/;�at���0�t�5��ݠ+�̛�H�=�}b�@����{��OH������g�e=���0oUL�����B�1�+��j���	|�7Sl���}&.��9���H�W���b+Ѝ���?�wx^�a���i��1f�߼�`�0�q�4z�<u����4��I	c�5%�˗�d+:v�|����7��l���gOױ�~��`�R��wL�*���2]�>�P��}����ʳ�;-��Yy�׽�������Б��K�T�8o��Y���W����b�Fzc94�'Ί�!�I�VKߟ��������׵�K��b�#�.߹����U���O��Q�ȧ�wß�-C~��1'�#G�;}߁��l����&�b�נ1*��)����_| ��>����{�7��~�;(ȷP�O@���y���f)��<p��T�C�C\�8B��;�j�c��qᐚ�_T�ڕ�A�Fv������0��g8u"\Ҫ��6H>Us$��x>	<,�65���#�6��Q�Y���v?㯍���|�k���!#eM4�q%�1�m�.[-�nƵ�M�z�q���`ƕ��L],�fëu���R��,�u0�ˣ$�.FYRI$�}ގ��^���}u��J���(�՞4�ձ�꾮�N��^�/���`��i33$���ء~���X��Q�g�s
�<�=��W}�L�ouC~�Uv�v%�:��O��x�Y�eM}>,H����^�r�~gLtfX�;�O��OA��%r��Є%�V��.��j3_�z�I�5�X��xGx�I�=�4'�R�3�~��.X�n��]��=�f8�8v�3�F�&,����y9�yLL�L�^��+j�U�үnj����������U�+ϗ*9������h/��c�T�0�BP�z�H��q���,q�);H�gY�����|/�sF<���vo������aS��$r�3V7b��*"q����|j$�܋ًY׆N��V-�י�^�J��-(�oI�9N(���Tz1n��
P3�N���\'v���̋���g���Bdĩ/����߮h�ˡ���������~�]�#a�u�L��+�u�A�G�1��3+m�N4����7�Q�9ֻ��"R���3����5wVni��_wp����{+*nf��WL�������7�4���=ۭ.9Ǘ���"?{7�^S�'S��laϹ[�����c�9��ن,�c�/n �$mD��o�XᏆ��F2ݘYuv�{z��<��;��fA�7]��yg����q��
����|M�<"�m�~Ƣt�����65n��s*��Wz���C/.R-�k�L7�<�����f�����W�E�3	A2V$��zH�[w���Y�o*2�W���m=�c���||��OG6_e��0r��=JN)}���$��a6���n��^�4�����שc	��\Z���
���q�P�;xb==핝w�~���z)يY�^�
B��fJ��*�N���ʩ�]~Q�n�E�C-z�'�O\d��خ�"|L��=��p{X���	�w��7�#-�}�;�uCz$�cE�B*o���ѕ��6.ݮ�=y1'�"�k�.�(�f;zdz������
�vfm��&���[id;8?u�'W���s5v��KL*3�*waK{<�R%�^���˶�{��O���]n��B�,MMTҸ�Չ7�,$.M�=��n��b3�+���e���\��9M�R�&ؼ����J�A�#�e��Cܙ�)���Y��{�xLv��xwh���k��mN�5�o�����X8�]�m�K��{v��r�>׹��|ԃ3�ʯΚ��gn��Ȼ�TfTFz8A�J�?{��-��˻w��q�B5�$�q�U���٣��������x�n	'<�F����H�2g�G+�+}/�R&CPR��mw^�Q���7r�P);�-�'�\�}79�I���"�FT�^��U���nY�G9�@���K�$,�͊3��МN��V�R�`�yԮ��L^���-�]
�e�p���db�\���k_&�j�/\HW�`��ry�3�i����,��w��	bQԺ\�弰$&)<ꑫ�r��MC%��P��A� ��[�t���U�����y�E��C/Znw�qeLi��9���]�]a�|~���w�/{g7���z�V�t_7��5A�f_��v��d]{cd�;�B�fs������q�֐+e{(�k!������wU�*L����PK��-ċl���{�W�Ο���O�]U]b��d);K�-)f������2.�,���P�1��V�ڶ�1�r{�2�Ua8��r��
��93��OS,�1���RF���ſjۻ�h�3s��n�_&��K�J����os��v�Z�C� ��dJ��5�f���p*ͪ�	{�ő|��:���4�"B�U�aW�Fh������.�`+��	�\����"�H�qˤƞ���pgW}�3\�o�Lr�Ưj�vpj�1��_J*�6	4/����ʱ{\���\)���AU�L��`/#���q��=��u`�'0����
y{���t�|y�m����	�c<���0[�1.w��uЩ���7�����ܹ��P�@@��[5>�Q�q���vUr��4�bb�K��C���PuJ1��HԶ%�>�sw�,��#��fn�
|���je�0��[ӎ,f]�ܥ[��sz�b����4ZZ`�u�	U�G�SF2s
���9���ӈ�juhٽ�����0.�p���pq4xV��uT��.�U�/�1G�-,�'b=]��\�5���ݲ��,ޔ��]c�[n�m�5a*�D�p�Q#�AMĎN��8�Uۢ��GWr�ˮ�-]9���ؑ-� =}�m��eŵf�Fr������_m�|��G)Cf��N��o3�I�:T0e��Ϡ��g�]�*�w��l������C��c��M8��/�cth�1���5>�sw���e��O=9+;fv��=p�uu-���x����K�+8]�����<mwP�y���G��eΝ�V��;N�;Y��,��u�ĵ']k�q��hh�n��\�����I<玗NcZ2�<U�������Ղ��gN��T��t�#�k�"����/�Uh*7�tʺy8jb	׫�%��f�O��j�2%պc�{�6�&��2�,T|�Oڸ��pme�Ti�61hi2)1-%d��̾��oo:w�
�z+w�����N
��]:�[,�����u�df>���v��~��7Q�X������W5��>�Ze�;�Z�{`�~҅�t��듛�}QM�ە��![���%��^��צ�o5��ݓ�͟����])pp8Z�k5�t�鴡�{�:�H�I���I�I��|�a�^N����c7�9��+b���n3jmNr�C�x/���_�Ϲ��޻�Ns`����J(�{���w����V�{�)�s�!�u
_g�wކ��J�vG=��g�2��3�^E����슧GS^���t��5ޱ��<�%�}B9ŝ��e�>��[�d���
��&���j�7��]	�ػ�Y!Tt����P[�`!5~����4\�{v��T��c��0P�_{�}����� Õ�;[��9 |N��V���Vi/H�/�:O���*X]l�%�C,��	��Y΁���.�7?��թ�����'�lFuU�\܊r'�yNh�ar����)�	��Fo�� �!���ګ�x�v��dע;c��f�\�ϟ�oh�+�{��w�џ�����1�+��۩��%�0��[���j���o��ݽ�=;.��9��7G�L�z�WE�źPF2�ì��Ef)��DR�\^���^���bKa�ls���ܽ5�"�۱�2vb��ƍ{��b�d]Q����0[j�����o6`�j�+Ux`q͹��Re�Ś�r/�\�w��Y�ck8��A�Wu	.�[�}]$cV:����6����"��e�5#�"Is���y�.��Q�h3Q$c%�����1a]��<����u��XJk��k.�ڍ�-�Mnk6�n����fש������h+���nƹ��v�nV��D��QāF$MI$�]w���c���h��\���T���l ���&e��Uy�K�KfΜ#В��>�q��/��������'�3b��i�?x��"0���+6wpZ�"�o�s��h3������k�xɁ�_����5�����o�3���a�����[<��=�xlH"�f/HRl�PG0(� /כm��%SD�����j��k@��*f��E�td��tǙ���ã3H���L\
o����Z���-�@ī���FJ��R���8����4ovoU]Ax�.��u�w�	��[+���F+�+������E}�rW[��k����2(����n��G�M+�f�h������_�h�;�dp�c��YR��~0w��k���G�0����4�akQ� S��-����t�	���p�N�b u=��1W��_̋1�{k�*��a�7�_\}
���?j�n���T���JÑ5�Sч��>�*��G)�!��w��[Q��Z���c��Qf�M:�ʃ}��@�*ʨ&$�gj�R&S�|Q|��}RĿ)T�p����+�4�N�V���Ǣ�3X�tg��[1��xE7xU�%u��q����8��*�\F��`�S�'Ձp�w[vpm�3���[��lL+�,�. кj��r�j���o��㞒|I���w��t�l��y�-u�w%�6�!COQ�jC$���E��1��fB\�����`���^g�+�&X�[s��{��]Gs����0��%(M�xC�.���3k7&���<��,��!�Q��랱
�*.3|_�������2<.�(��w�88���(.R���²%�K,LQ�Q�j���[fz����D�=S���Էr�׋�u�>;[2�$|�JR�OuDh��Ęk{�f�:�QR����Ά��^hϷ����nhbɏe��@4�\��|�/�}����RrV.ݐ]��8���Ex_�9��#Ҷj�z�����NdI ŭQ�09�{Tㇸ��yO���|5���|�ӵ��n슘��G?s�FW��=�4K�ʢ�?s�>��%XD���s�G�l���-]��,͊�a�-,��LJZ0�q��8�g��9�'_|[Gpk��;�����x�ǏF��s�H��{8BQM �"@��i ���h��$9~��3����F�WH��5Z���j	Q�2��C�pv6t�VT���U	�(WP;=!����ᰱ�$
��u;�Yi]^@�p�@�{�`k?7!�Υy/7mu.U�RE=����"���s�wO����}��Bt�i�r�xƧa,���U�ϭj�Zѭ�d���i�n��,g���f*�CZ�!a��d{�աrW�,�;�\HL�Zq��u�����B8���+m_�G=�w���h�|6zY������K�s�W��Sk
d��>W̋���-�网.7_]=&dY[��i2v%�z��2g�R���4�-}�:�����)r��W�p��FcÑ�U��81�y�M��fh�4j�����ՙ������sGҦ��'����_9|HC�
��mx��(���ܢ$=��֦�ÇL�k����E��
E�G�n�ρ�C��bv��R�t�hz�Dw/L����w�X^���{��T{�X�c��ٿ�7�������6��½��k��˅i�����:RS&�0Y�r
��	D�F4:�I�0��O��R���I#�2F�Hͺ5��ˤ�P@�`J�[9�H�������_b/�W� f�O׻<��H�:�x� ��fI�Pc�UQ�wV��Bf�����%s��	龀{���6H2���QMy����9�(B1���v�z�N��m�3��u)n��%�*X��:<`�޵n�8]
=.������r��O�1M�G�2�M)ŕcԕ����*�����Q��W&��Kp�n^�7�:\��}bs�_;����%W3���ܭ���՝�cm��	�r�:u�<մ�+���meM�^�����s
%�?|�~�;
6���jj�x/@���V]��ϭ���5;3�G��zaZ�
0MQ�K!��;LG��c�xq�8D�׆Wf�J�tۯ��,˚m�|6��<\���ܯ~�gL���x cݘD��k�/���wQ��0�O�#v���5�-�0jy�u�9g�cŠ2��쫩��Tw ��R��5'�fv�M6W���4��򭲊���Jȩ���i�K`K�jQ�S�=�a�3���(�١���vC]2�+��FAH&���HƎ����Q����|��_o/K���	H��`�&�x�`���j`�	�f�Yى�}S�!8�>^^�Ok���B�V�A~<X��.W�ezIyX�tf4� ~G�+#y���^��|ѹ���Y<�q�4��"=�l�=�,z�K�Wvމ�]V���#�4�$\��f;���-N5oz�����gIYlxa%VT�L���P�]o�#��x�ðjsLM�^�}C�r��Fbyh�p�t�WQ=+��ML��2�:�����p��w'���ؔ,�z6Ϩw|�W�=3�*K�S�NB�-���en�_��·�/Uu����-oR��AI*��wyi|mQ;#q�<,	W�i-��Q�6m�C����k��.�v5��#^:&r?4�i@����nа�kYm�ѥ���R�HXM+.�J��m(�=K��#�3�|���^�Ulw6��lj�Ҳ��X�m-4d4�ױ�j�2,�l����[+:4[L�rI$�}蛗�
��+�au�C_�ksbA/cݙFbRH��*���"j��ኍy���1w�NDu�3	c��֯dqd.a�u&� `�G1�}�7���bF���I뼇	g�5+�RbSђva}=���U^���h��kT�9��g�����߼�� �!Vd7�	��S?9��`�$t!������lE�v���,�Kr���P����
Td���8��&��锗S>�v�h�ˁ�-\��d6��l�����e�e�
�Ku���(���E*�ިv�Z��'�KG{�Eo�z�D�ۊY�b�T�C�������T��1��e��v�>����I+�T߷cm�nƛ�ޕG}~�®ڦj�������Nn��#W:�r�=s5~�z��	�z��/6+����Bl�o�]������GnN��ne��#u�
�8�\���,f��Nև6�T��P��ٵ�2I�IY��R0��}V7�~_�
3Z�<�e��׵[�i0a�(�H�\zt�)�=":Y���T,�1-s��w�aB�HcՋ�,l�2(�)�փ;�ʜ
zE�q߻�߳�����@��[t�U��W��k����D������j�f�I�=c㓏`��wD;�g�e�τk�|�ͫ�6�&����U�c���7;��G8
KfjN��d��aK���{��޼�R��ι��<s����=�0��D,�r�/RV<��L��&�^8�ݰ$�5��`2#\�2M-��K�6�ۦ�����K��G*���	���o�g��C���=,.�N-�)�[��Kdd���scnT鑡y�v��Y�C��2)�4wulSF$^�o��+��)�9��O���z�X�΢�e���N� p~5�q+�<�����x^am���7	E�����E+��ϣ��vˇ��Af�Ǖ�B�
	�̠Y�ٮ��t~��Y�wzл�e�c���Y.έ���-��o13ʎy�c�~���ϔ�V=L8����L�kM\1��- pM��Q�qζ�����B�ދ�,/V]���*`R��"��t�<�ʝ�|T�Y0�����냧!�&�9��s�.d�/�Z��Y\�ޟ�b��\�</�2Y�tp$g���l;Vٗ��~��~��M��C��.Vv�aAGF�*:K�y��]�B�@��3�<��3���z������Ş7oO޾M/��o2����ZBZ�۴0���05�Br��H�~�W��6�FOa�ҼEGÜ����.
�������*�+��V��8sb[��b�R](�ι(�ʲ��E��������G���Q��0��>����WV��vl\��m�z���ӘȗZ�{��ɩ�������v~�%ߙLQ�s��Z������(pK#N���D�p�'�v6*ѱ��S��s�s�x��H�����Myh�EV�����I{�:���l���a�W���6N1#�������/��.�������m�V�i
�漓>��0��m[����28�i�����㏉e}��@����rTSɌ�jc�32���T��h��1�=Y�s&��pU>����d&�:C�}2&��G��Q2�݌Z3��sW�r����? ��*�t7�3(�����塝��$��޾���=�؍-v��ݘJ�w]�&��"NĠ8��N����v�(M?a�>T�\^����}��5 a�G��蕤�:������'�c�U�w+ 7.q��	�)��i?���L�	!��q��5'���]2vJ�+y��uۆ@�%C˅�É����p�\.DoEޅ�^��o��q�A9�������aq�1�e������Tq���Yu�C"CI%�"+:�Fe6F���Y@�_�ֹ�hw�T�+�W7�w�:�X@W�n3F�TuE��{�ck��SWPHP���T7������.�X��K�W�N�i�̓z=Z�nN)�j��lwn��o��\��%\5�{�^=�`Yw5v@�o��o;��4aZ��g�N{W�����r��W/��tG���}��5�>���FS#�}ڑ�@�wz@��_`R��r�
Q�o(ꗂEFNM���R0��3��w����n7�BU�%���p}�YX"k��	�}B���d�p'�����3��F��K�	ȕ����8Cz�Dy�c�(�Ig�����g80�
s������o�^X���VX[�3I3��e�K�����%IG������1p�#�VNG���u�����~xxTöG"�%����SU�W@w�Ĺy&�mv��f�����e;���I���Wy�U�m��&�ץ.X��Y�sV@"�,�r<z�7�Xa$��Ֆ�T!~S��P6��!�O�=1�9ro�b=0�p��p�&��mO9����2,y���QS���S�Q�پ�^z&X������,n� t�b�	��w������#\�LuD�G/h	�f{d��K��v������S�%�B�dm#��5Yf�Bp|��Dي �[��W ��l�[3�N��=kǵY���r���6�e��Z"��ґP�'�>0�%�uߙ�[�Jĉ��|�ҭp;A��ܴ�R�7��\�o3;�y�5�Q��r�jʺއd¯v�=��X��S���RX�ݱF>Y��%��O�lӓ9�U�m��3*�Ji5�D�'r��}�K�u_�����6-쇩+g�Ҝx��*���uv�J��h������uu��М�<�h�5�yfkm�K�
63SsR�jKE��xMڞ]%�Y�F덺�[��Y5p��%v�����hջIס���6�%u�Ik-�j[ �� 9��\Z㪧����kG�)7i��׾��I��<:}g���O���j�e�W\T�r���H(^�oc$���� }�{��Y[qr�(r]����h��-۾sV�x��Hn�E�3��٘�]���`7�Ѓ�77�9����rf���� z��U�]�w�m�;Q�뾌1M�"��E���uc���,��?q�Ή�0����Q�hCP̀�b����T��J��:�fX��.gD=�Y)k��Z+ښ�a�Y�Q��.��;������\|4Ɲh�t�N~&3�[7 |f�L���]��]����di�l����h����/'m���m�Qם��T�"�zRX��c�.zz=f.tK/Z�<�`���ǳ�me�RN�4*s�H�RR!%���L�ET޼��sr_�˨$2���]�<��\��Jr٩iNۼ���E[sqc�$���g]��]əf�;�y~� 6r��A���Cяt���EY]+:�e�a*�]O
�|.�g��	��!����<�p����g1��=�
��� ȇ��A{f�]8����#nB����k�Ԯ�)���5|�R�U42��2=�5+8�Cʳ?�Mܡ��7��"�] `��\�7�I��t��k7r���I{�X��A䊘�uWS�YU�rZ]1M҅�aq#|t���c!�q�7tHI��>��^�3Z�7�U��R��7�=,��p��:&�������<28�p��tq���;$9uwC���wυ1�w��4�`5Lm���:�e�;/m��CP�Y�h��2�n��'+��m���:Q:�usk�m��D͂��*�q�s�IݴvI�^8� �2f7|ouY�����o�m^;4���]�]�e�P�*�n:F���)�Y3����.�ܳ1�f/$q7���.�}���!�c�O������e1hպSf�Y�D������Gws���0H ��G-hT��;:�4M�s	�a���e5[�m8݅�'Y�����2vWA�CC7s�3.�)����,�*��&De��|Y��u�td���ٟ�W���ʽKE�)U���9]q��e�RK�$�@�/V��-)k#,[u�v�em9:8���;�j%K�4:��k���Շ���w������S.,C�-$�H�6-5}XAghV��n�����;���1�&�D�uʔ8���^p��KT�_]�j������<�R��Ž|�28�`��:t�;ɷ�yᖟf�)<���c:Sµ��V��@��3x��ܥ�.���9;��,�R��̖�k!�y%�L0�������1ݵ�i��w��oi�{�\bX;8B(���:���C�x��bxYW��x��+vށ��hl�� II#J8���$����3ێ��ˢ�W:�7Y/7!�cb[�)m�wki����̝]��(�ht罧�z����@���w2q���{�U��h��5��k-@��LAv5�㛷z[��!�ÁL��w"������<��U�#A_����L7}�\�C��wͳ���ھ�G7!�wd���I�:0Y{J�S���X�m��������N��.�Z�BVK�[��H�}�L�vX��ٴ�C���]*����ʧF
��Zu�A�ϩ+��5!YWvi��F8�x�N�%�S�q�m�T*���&�$�"�42���)��h����ZN����v�6��m��0�.���E��6�Ԓ�t���6|�h���|cd_/��i�zᥤ����=�T�Ć�fe��Mv�v6�i*Ka��3�C��,�Mt��Q�t��De���G2j�&�V��X�Q�Z����e��lёk��V�]���_,�|�a֣2ۺ�5\ZE�J�;x�f���&�l�	+ ���c.�ao]��Y�����U�d..�FK�ڻV���Vݶe�Y�K�_���|�mF�݆2�2�i݌�`�ؓX��)��QeU��kիMn�R�%�%�a�^�6Ֆ�5�"mQ��n�)C����,���h��>B��v,���k]3d����i�6sg�%m&����l���M"��6\F�cXR�Q��N�ݮVɶ�$�n�t�]i��%i�T��+��d��%Z�t�f+�[n\/J�b���i.�3^�+��Қ;JԩQ�HI��ɲmQ[HE�B�d��m�          )�˫�6
nJ���Z�����w�{����y�2�W,�v�v�T{J����d�{�6i�;]=�0�l[knC6Ɏ�T}+w��5nݡӺ�,��� *V�������y�꽝�eW`���ӫ�K�@��Խ��3���YŦ�]���$��t�\=�ޘd�4r{�A(���q�ϻ��a�_��Wh�W
���ϖ��D'�&����&|��a� �ˆ�p�iJ�v���>Q����s��¾}��M���k�$��5k���9�1�X�/��L1�;B�w��(f�)�7S���kx���&��&>/-Ъ][�W2j������ȷ)ԡWC�y* �r]���ʖ���y��]ի���\t�<������Gl�D���{�-p��d����z������u���4���U�dmݪ)L�@j6Q	��<�~.L���)�D���5Q"n���;��DH��G��3$N���?v�d%!f�����|/�L�,�M@�Un4#���>���H����C��[��<�|`�h�D�F���:%}�g��K�ay��JM�����5d����τ�7����y�Jq���xڟ���ϵ��v�n{�i�0��T]o:�Sj*��j�n,���g�)���C�N�y�w+���ڸ��%�<�|��hw�~f\Y�fח�>��zNh��"Hts��k�����"2wp}ʄ�$ʯP�+H�c&P��RɆ��܁��j���?j��a�`��ҙM�������:Q�C־��_v.�=��d.��Py�^�	./�7��"K���9���y�[�^����E�z^n���ŗc�::����{�6������v):T����"CU����˧����[a�|;O�~������O�*��Ы��u �������^�h!��M�l:ڃγ~eE���>��=6����&�Z��W��Bur�'w�@mRa�"�B��u�l�e���2��iո���8%�[�Щ����jqpc�a���e�JͨOٳ5S֢�н7q�ޜ�J�p5-��F���P�8G{��B���VӪ�U�[ps�\�RQ.)��U�찫R����Ǣ�ܩ�}~鮖]󇵯�k*�-���w�������I�������z8�7G��������ތ��}�Ol��ҕ'��uA�V)Q��c}���lo�O��UA�e�K�x��u��'�}uy�Е ,5mN�KÌK^�_W�y������ȝ7^��hJdK�n�p�����y�����J	-�aRD�E�.H-� BE��wF���kF�	�I�4o��O��ʲz��7�Q�ڏ�	|���t���������Z<z��n����j	U�6G`.�/�}��j/���>���3j{���hz�����W]r����M[�ח�y�J�3/"��K&�U��ى��"���kFC[�ڕ��O�e5P��Wd�m�'��ꔽ?���)�R�GI���ݒ�W�O�Y{Փ��Z�sM���\:f<�9�u�Zl�Ի��t�aI�-1r=xu�3S]�ӆ��s�Gf�$c\n_����VΝ��g���"��������w[��p�)z�c�r7ՂLdK�=T �Zk�)��{{r�뱼6��Ւ�3>}1�P��$΁�b�o�Y	��+�deg9�/d���:��E�b�{6<��q>���@�˕1чD��4�J�~s0z�b����_�[��.�k
�7��B^�a���U�r/������܌�&���w�>�I1�,�L+T��Q��` r��[^Pwj�k�ґ�i�wk�]j���ua��a��B�4�fM�:����E,d�B�n���bU��x�cQ��)	��i��lt��xnb�2�k+�]��8�dv]���,���sK�"�nG5g:9pץo�)K\%1�\��U�;����Q�"1�ײ5�2�5j׻=<T�=��\]�-G��8'�~G+��$֘��A�eQ�$>���x,������|f�@f|~?��_J>��_��ߪ�	ӻ�N䏦P�+��W�Al���=�rQ4��ma������2�?q�h��j�zQ�ۘ���j��ʽ+��9��⮆N�A�1Ш�qvk�O�H���NW��C{�v��^�W��M����3e:��l�0Ã��B1�Z?z���2�ܭ��.I�����^�8�!	�x�)�jY�&�,qKrrb�K��C�՞�w�.�ʀ����zj�N��Gvv�FZ�˸u)o{`}�Y�2�m��[��jΦ�-�`�gu��BĴ(�լ��^�ۊ�)$��A�R�(��bb<](��QGE��YjK��ӳa��Y�m��&�)y��ɴ�T�̒���Fl�l6����Ivқ[[�h��5��-� ۉ"��(_$���m�{��w�$��"�:?�,�����ju�<�|z�7<��Y	G�i�����Q�8��(P��m9<�#$�KC0��\5 >��F����T�m�z�cg�#p�炀�$��f��ݑ�3� O,���Q�{�OWLetu׹�g)����C�l�Q�U��1�l̂i�{p�yR{���8�4C�%(!
�`$�0T"a�i�!�g��0�H޲2�������ȸZX�6M�bV���-�q��H�J�?N9�[����{"
U��F5C��
��Դ����U�V^9����˥o���Jk�kw��i˛��E�cC-}�*!^jm��[���n���o)��:��(�������~�߬H��3�R.���S��h_�S#�}ߕў}x��x�yz�%Lŕ݊d��� ���=�W�K�]gȥ�+������L/Q�7S���'��J��<g��~�'�� q�y�S�2�s`������'�E��z�6�{l<G+;�MP8�y]K��q��g.c�B��o`O0��c�;�1���4i�ee��-Y��L�d�_s�h=���q����(ɧ�'D-��>�+H�;�XA��z�j���A#5v~35�5av��n�֕�n��ʊ�����pv\�T`Hou<|$�Or�7"Pv��܉���z�Ŧ��"f�ټF��).�\��׾�;
��&*�qo�cI�>���l�]����x��½��s�U����oʢ��#��U��r�1_%����0�uib����Wl�d��r�u.p�s�/�STGH�b�V�n��6�4s���^���h��w((��׻ �;�q�8���딆;���nr�����u�7���%�I���K���X�6��T{e�^4����iO#`�����vE!�T�<������%F����A�}]:`�'���l�f�x��b۸�h�X��,��]��J��)�8�k���1+�m�u�x���=`�������:}G4����]|����V�V��k��2�����J����ͤ���v �u��>T3�
���P7l�w�q:o���u�� �q֌�^ܲ��@���ۡ��j$�֡!щ�K���*�s��:�Mƨh�eC��邾�"��T�9]��н�#���5�B��A���T�*~�n����� ��Q|��H�FGvt�y�������u _���H�ّ��J%HPm@����U�lV1FL-x���	���#%��s/�+L�j��ڷ}Ze�U�j�N���ݍn)��M+�y��'�,oQ%$r�d��圫R�63�V9ϥ�3��.�����x�pc��y~mF���Ώ`ܴ���Z��-t8���'W))��s���n��Q
�y�.���4�e���M�����4�!+��Q�?*�4�6�����AQ7��<����H�p�~[�Q��5��X;w���OYPow��P�����'7w�U�X��`���ʛ�gx���|=bУ��{ ��'[���]�yN ��#W��Lx���ld(%���O_C+AI�hFr*��% ;1��mJ~}�Q'�^*�x���K�y��%6<^�3Wn=�K�����>(;�^ү���x�����ͼ��ø��/l�*�y�IϪ��.�@��d�#A���w��wUU�q䯶���u�o�8Sq�U[�g3���7:�*;�I�R�f�p�A[���e?d������ ;��L;Y��C��p5��߅R��Uʫ�3��"�E�M|�H��%�P�h~`�3O��O�?d�j�o#UFƾ����߲��	m{���y`��а�`����º0x{.7i;��^��-nXc�u��I`I�w�>~��^|o�^�fcB���;'�j��*��q��w��X�){R�{��;�\�UY�#����r�P�3��U�ի�"ԋ������0���	W=�ۆP�Y�HP�89��\�� {
�R�ޘ �t��ֈ��&�*?�����+�,�>���%y,�8X�u�=RX��;����ڒ�[��}��]�|I�k��GvL��yXxn�av]ʒv�=��qC��ǫ&��8�ۃ\���<�MY�a�G��*{�@�S k��ߙ���l$��A���C7����e����et{���H��n�L��UR�>����?�Y�Aۮ�b��.��[���*)eT�n��ۗO��۩thFE<k��.S� P�%c`ʝ�v���ef\dth�qD�G�!�:'��`
S�+���A�JEe9᣷�D� �^p��y���/ڽ+�u����d;Q!pd��0��!��.ی��$���c��[�
�o���cXZZ�0�F!\�>�ؤ|�3ꚙV��A�s���{x����xa�eH�6��ʀ��,�w�j�${��� ��ǧy�r��}V�=��N,�/{�@�P�P٫ʢK��V���u]�)�����@� �LWyE��77>U��y��������	�E�v��1�ɋ΀��'���x�1���Ҍ7
˺�kU?\�l��~7Qg��a0�q�;��;�ʜs�?K����e���º׶nN�����C��J�]��Y[n�@&#�P��)9��u.�����f�2T.��O���k�?���Xc
wՊ�3KAn�|��S����4_=�nHP���c��,�5��ڹ�'"]t����.�L���QQi#׮�s�H�]$1bB:X:dՅ�,W\7mЖh�a��I��1s\��m�3��ٶ���[46��KMd͂FRMu�s)�.���m��Z[�٘�lGMl��L���+m.���k��P"�zxYW��!"t]pS
�؏_.Nۉ���DǼ,���ʤ�����;W�H3v�V�e�_?��	���$V^���:�߮�~���؏�|X��T;���C���������d�y7����'E��X..<�{D/n�r#F��l\�ӯ��W����O��y���eӬ�%-%Μ�C!�#�bv5l�c:�5��{Ha;S�6ꑽ�w�"�+�9�Q&�
u]y8d�Qu.��kT�W��7�x�}��o�ǎPv0F3���3��_�*y�NGFm�.n/�.�º��=�,��w�b��Q[�!�Eb��[<���w�6b��+k~\��i{5u�#�H1Ӭaî�7϶lC�磝z���kk3�fK��~��p�����{w�����w@^o�4�G=W{�<5���n�[d�ر7d�o=�#B�8�7nb��\�����:�~�E��E�>K嬞޿~F;�)3Ғ�c8�ţ�'�Z�t�:���"K��p��C�Z�Yáuz��N${.
��Bf{�a�rMfTɀ�.*j3��Y&
����ʺY;6�5.����Jգ{���_[Tk%=/�dF��t����Ծ�Y��ؑ��zМ��+����w0Q\{_+	�|�� �n=}�WQ+zܴ9[btu�M
��n�����������p�ZЫ�^��R0��=�NA�l?�'j���F�3���L����p��[���ˡ/xQ�T�l�c�D4K�L��(��rs�\�Ny�	I�Z_�Um�� $a:0N�~�f�3Vt(Y���md�]o]��2��w!��-"l��$�Z�yՈ,v��k�ȼqkѻjOnD���^��(�;k�b�b��15+��۬�tl���ޘ��e��YyU��2f����S��,Iv�Ǽ���3�{�2��b�C���q�5�g+rTu$sf��a-hS7Dq�n.�<c�8ݒ���y%�&�)C�E�lm;�6u�j�grS��9a�^ܵ�Mm��o�=���/]�g��LL<Ξ_G�sO_�IfU�dr�JځU����r��(�[�ZFk�j�==��]���q~�4�NW�;M����ڐM����PO{�T��FJ���~|�h��x6R3t;#���->X�T8;5�U�,�s]mK��I@��1�4[�76�dn,�`�}W�	;�*r�!��w+�wnCV-��䗺y����^/�2�{�f3}����<���K��r	C.�5E��Ӱ�F�4?<�,ܣ��*�\����]�ΰr����~��w@�ԗ�7GJ�\wl�]L�i�Vh+�X�k�vv=ވ�Z��k=�Y���c��b��$W[��L�;��rA���Ж���C�xj��Lʹ̫���;�c���f��<б	BZ{�����Mh��gM���Ա/"�j��=�6Gl���n�4�=]Z�^�T�/ �A���I��&�8��-�7Z��u����l#
�����WQ�sB���pUh�ɠ���;n{j�6�<��#��1�;�W�Mwk���P��TXf�:N�({��&�	�h�^��tT�Q���&7Cu��x�9�W���s0��V��O�=�]mV���K�/MnzaE/�RK�ALV�W��4K6���!u�r�o�`���~���˪�8�ĵ>�ℊ�7ss{�RfF#�(ą�Pi4 b|b�P'#���4#�����(!�{jl���dx�%�#��|&ip�zM_5j����^��KG�vw�!/�w�&���;���h0z�<ۦ}1��WR�i>*����p�Z^��9�J�;4v�u���+�c��_�� c./gFƚ46N5u��p���F,ϕ�����W�;1�L�ge�_�ͫ�[����U����<��p��q��֞�� �����k�ֻa�+o5��a�Zy��:��{��U����v�\'Pj�eM��c����;����Ǹ�8㻿����q����q���N�8��;�8�<w���wp��tC��#���q��Owq�po������8㻿����wq����wq�����������۸�8㻾��y�������j�������~������V�_��A4�7`[���X������2и�Jهa�m�w���*��R�y�e���ν�(�v�*j��rL�&͘��9Pb�l��k�z����xZ�y���H�YZUӝ�_R�Vk7m�̣�m���C(v3u�&�9��хP�cgvШ��w)�BKÍ�ه,���"�#ٚ��õY�h=���l�cqb@�d���Q�eJ�M\��Jٌh*�Ո���gv�k7b��e�B��f��+"2�P����):h��1c��'qp�!@b�v�Ǖ2R&��	m^�z)�
�2�Ӫ����+��vv�1�����F���;D*UH�:�_:Ѯ�a1���!��kb�=�KCOAy�q��*���`�#udF��K�1�^��qmhF���ҝ�3�ꈰ����o�[v^?���m�<L=w���\�XK�X+�����mE�ThC��ԭ��
�V-���ZѫabP-bDkX{�(G*+�'(�,0�S�ĺ �6`[�h�cRGQJ�m�Qk�N[�@��'(��Ǫ�@����,�Z��ă{I�L�	&f�����ڻ*�
W�
�3�*��Q�*�2�I3r؆^��Mn\��[�)CJ�N�~-��1S�v��2M� ̎ج��Z�y�mI�7L��f��t�e�4�����+����O&�!3-��,=v��PY	���f�#V~:v�0'4��摮SE����j`J�alem6�3B��Ӡ�ֱT@�l%f�
Z�:�4m���%me޷�Uk��`���ɨ%f��o6j�v	4mU�ے=Z�&�� !�rT;�4ab�-��j�h���E�1��	'6)���T#I�jؔ#.ۺ�2��76A,�e�om÷�IF�$ �p�]lܤ��R�6cD��QB�n��:ϿG�����wq�w���<�wp���!��wrwq��w��������q��<�=��q�����w �ww �������q�����������;��D�}?�����>����������;��q�q�w��P��;���ơ��ww�'��������cw�ww����ww�������8㻿��;�8������_����O�=��q��O��������������#�wq��������(+$�k*F9� ��;0
 ��d��I�|^�}z�)N�4���;��rU!�$]����
"R�v�J̈́� EfI%U"R�ԧ"�AJ�i"�H��*�ƐTRIH�D�
P�		RH�mD���UPD&��T�_l �(���.�B�R�M��$$J�Z<       t# Q�P�l��ćc�#�   � (   �{�(����$
�S�8;8�u���hَ�n�� ҨA�ژ@ m�4��Q� ͍U�o�=��C�h	 ��ڵ�F����m]j4�� :S���)0�6J��htv���)5�RIH��m��5�^�:�m��P�z� :�Pȥ�o`��ǧvȶ+lb�)ӧb��l*��;e�Y�f�U6+mjU$����]�V�-�]ݳ	�ɚ���-5��ҙkmө����H�(*-2ْ�*���r�cvu9�[j��PTͭ0���M��v֩��Z�I�ہ��cjWv�aх��;���Hlխh�Ww]��lT��t�ٮ�j�E��UEh�)D���:n��Ӯ�Z��eT;v�Tv]�f�Ф�m��N&�-n��.�WnY��ؗv�w\�4Hi�쮭��Ge�+gp։p�N�ۻ�UP���bUQV��Uu���f���փ@{%f�����7w��:�C ڢ���m�m�+4H��9��٫�n��-���6�T��\�؈F�igs���D}��w,���T U
F��Uv��lU�e5�s4�a��3����lt�w.�J U����;�����5�vۨ��,�*�lbA�ik.��X�ӺԄ4�$��IU*��©Gj�R��NZ�����P���]�j�V��Nn�v�p�h;�WY�.�nt����:۵��-�Xj��-6�l����n�]V��	62�b@��IH�ѐm�)�t��n�u*�U�`�-�Vmwn�E�-�r��Ե��w7f�n1� ckwiv�p��u��ف�r��m���:\�V��*�T;J�d��v�j�9%C �id2�uӭ�����kj�wr�5X�cJT;��e9��Y#;��kS�-��r�v\��s]�q�TT��Fl]�;A**ET�
lD�k\Ӧ��kiK:uJ4M[;sl�ժ2�n�;���۱�:�����m�n���C8U�h�k�ɻ��֎��T5vt.J��]�EJ���IP�
��*T��d ��a%%*d  &��ԣG�  "�� ��Pd21j��&T�j� �I���O&���Nx���B49&y=��U�jI�\\�i(5"���nk���y���������� I I>󾼹�?�������� HO�$�$��	$	"			�-7����Ѩr�mp�P`��l���B-&c�B�?��/.�x�mѷ��uB���ḳ�!Z���.;�"M޻�Y�ȶ�	:YM����6�νb��Dl�T��x!��K�R��ijC^�O"P�`�� E��`�G��y7�*�@��x��&b�X��h,X!�p�u^�[nB$A�,Ru��XVƽ�b�y+5dyn��S.�O"e��0��Ū���`Zn�X��ʵr�)�������{�]FʄḖ��F�"Q*ْ-n�I�����lɥEv���ido~ ��F�E���{L�T)d[4����'ie,9��땩���+D�E)�m���mY�/"ts.T�`H[V(�d��ܒ��?4Ѥ�7*�
������A�KJ����D�XqRF<�3������J-4�
��n�(4ǻ�j(��Ԣ�V�2P�n}be��2+r�b�<E_��UAV2>?� |1���煃�Y��L{W.�-Ej���TR���u� ©�H�meٱ"��B�1b���zU��ѫ�&
�ǫڵFh0Aa�<hә�t�؟;�X����-�Vպ9CRBlu�^%���x�*B�����lke�����X�hf��U���(%+ɱ)x6ն�gE͐��Z��u`�H֭���o6Ј��;[����N����^��<6ooa&ʫ�֋Ŧ�Q�u$6�J�tVٌ��V�Z�kq"�]^!�i;�/F<vJ�>����ټ2�����RB�� ��91q�/����hKxkm[�����A[�"�t.�`�i��+[��?ӑv��,.��QN�:�x�-�#��]��E��K��%n��׫nh	X�n���W/ �Z1
�zikWBU�3o��w<t�<b x��1b+����U$""�Ab�"(�h Q��(��?YLy�rr,�?@���Q�3
ͺ��!ؠ;�U����o\�Oiּq�6��ꬕw�z�"�4	׵e�i���<:��U]T�(�1�+v�7�O�$taƻ1;�Q4p*-m���{�EU&��k2�ڞF�E,w��*^�w-���u�Rm����I�5������L�,8��Q C���]��G$1�`p*P��'K&;x%�X��7y����71�!>n"�6}��̖E�"�/���B?I?�T3,(����T=X2˪����Ӽ��y�u�ߒ���F"�a�AR傞%O�k<|ּ׉;8I�^�)�"ؓ����HT��F�"���*"�R(�
E�E�)! xŁ%b(���s���k3;����5cp��FC�4�/U�u�tj���i
Oe�r<��p�MћN
�,<iL$�{����b��Ǆ�[ڻ���z̢@�[��u���KR�$u�� W��8^���JZN-�&�����b͂�"ȽZT�.���v�mݺW!m;&���������"�E�	&�wsYw�$��)�Hْ��q�OV(C�Č8�^d��&��MV#c�f��lh�j�6�����h۴N۹�m	�)[��#i���O6[/(f��VL�ì��=9� ��fnk�I����" bE�f��7b�M[��d�?
��������(D��a�ߣS&J�ә��6��5�(��.aD:�FҐ�7�FQ�n<�^@�[N�,�1�v�
�����.�Ȍx�,�̣t޻�Ą#7�4fj�&�����H�iD��W��R�sA��m4V��ǅ<�n�6�e��a: �Lx;,��he�a��Fʧ��eؤ�<�e�A5k��J��0dw+nJ�N�ݧB���[J-�_�,�ڹt�L��q&���N��Ub�F���Me��h�H�f�yoN*��bbi�e	��F'ye�.�r	O��u�OBa��۬��+��K(^�'r)�$K9�J�[.%���t`���w��uq`EB��5�9�y��<;��� 9����{�+b�y'v�l�9z�Gh�>��$y�(ݜi/��e,���ů�cUlȁ�.G0�iGh�F���3c�`�0C3sr�I8K�M	Z�'ר��u��`5���&R���q���u��E[�b��yVu�C+k���*G��{Q�N
ū0�O����а�2��"� �_}�!���cEAVEX�aCi��x�D����V!�e��w�=�O5��~k�V�,�sQ�����/�D`n���hup90ll��Ȗ���wLش\�6�2>h`����]B���{�/-��V�#q⍌Ur�,��fF
��Z���w�*{�li���n�w@(�#TR�����֋o
g#ʑ�(�X[�U �Vn*P��>���fϠ� T��$ے��n1.�/It�2��i
{?�CF��\�6cm-;X+p�\6���N��L�nV�[J����a�ú��+"�,�V!�Q�)a�%�&�^Rܫ׵��Bּ���2���Z��IU�\��V��&4��%]��9Z�Z^A��it"�y��m5���{8@~����Z�LL�7/�ј�e��\z���$�P����͈K�eG'r�Ԟ��V5���b��"�"��qõ�mH �m�(ݩlR�خ3w{�Y�`����X��I�(�F�D��f�.��B��f���e����v���SV��y��*���h�6�����P!���8��4S�V!!J�qP�eԡ�Z�l��k�6��`��Z�>{gm�EX���� Z���"��9�W��E���ݹ��,7r���&b�]��ڈ�
e=��
�l7bX�0eM��3m]i9��13�q7��h�e\4�5`�7 N��V���+KY{��u�ǚr쭍�j���/.c�p��Q(o���	��LR��@���y�b%��¶�8����e�t��.��րu.��Z&HX��ʨ�"+.�,���3�`���c�$�l��eb-�2�R�݆�i e����!�Z2��}
� `��B)H�$���~$~���|��*D.*~�(�Vg.�n�ӏ��f �T��u���5L^'�%�h�#��9i+�ls_�:�M�fMW@Gxvl�n��0Y�͋C�4`n�<��䣴�ۣ3-R��h��B����3+1\ܸ)Y/*}�ʈf�Q��J�/$`��n�*r�f�C�WIj�pX/Cp��#���e	���wdg��d �K�71�����@ ��޸�PW�������*��*ʻ�~ܘ+"���:������y��!3�n�aխ��fEn�bm�HI�0 
AA ��0�Hԋr%wZD�+t0V �&�V�skXղ~��.�&#�R����D*x��z*������v��t�moJȕcE��й�Q�B�z��	x���kLÈCI��F���ޤ��S�R�Q��%.�Md4�s*g�ܕ��킞�׉��T��֤�9�X	9j����PU���_ջz�!im<��6e;��76��*��!�W���b9��!6c��nb�̈́��vm�C���ô0V�̨n�$�PSLi�l-��v�)	��єV1�����ƣ�-�E��(�1����;x�+qۈK�Q&��(1���r��U�U�l����6$3+rٰ��"�\�NL��� ө�=*�~-��n5���&dt+nh�@���adnRǌ%X�4�� �m�х��4�`�V`���iU��dlW���� �ѻ5�5�R�	3�4n�g��j���Xm�"�ܳI��r3��骮�w%�i)�^�;y��]���z����E)yr��e�+U�X��nz���9&��{�f�.�#z��Y�ٔ�W�W�F�kC	���u`T�j�(t��in���7bʍV^��	@F����5=%�z�vSz�EZ��#��J%+"�E����w{cSy��4�2m�OR/Xu5z�V]O(e /E�~y�I�)~�캟C�������#��QT�W�ɘ�ݦ��wD;�ZSkQ˼�BZ1؋ ��X�Q(�)�o�E�-*���V%�ډ����,��E̒��FM�j� d�M+R��RzP��md1�sD*�_�Kn~�t��e��¦[s`KY�"���N�e���k^��;5����B;V�f 3(RD[Y��n���CX¢��9��mRx5��Z����)�[�`Mt��ug���;nӶU=���TUCW��Gl9aͱZ�0�K�]������8������
�X��[�m�4ڨ��0�.1uf���S��{�pۋ�ɖ �7��m�*�^���x���S�	Ʉ �R��Y���DLɳ �YQVp3C@�Fj`Ţ���)��K�[�e�eS�M��؉K"��� h�^\YY����R���yKE,�7QV#`�[���c���$��m���̼;E`�9�&�,���5��F�ܼ>��@�1ԫ�-m��E-��wܩ4��,G�L�� �l�Y�7i;�3i�*FM��{ �4ģ���-l�kv�]�t�#-8V�˴��,]�!�ki�]�D��ȥur����x�b��Y�ǐ�I���b��,9W%Ӻi�2Xu.��+7鵱Jƥ4�kf���0�R
��M��ѤZ�75�I��vR��&Ė�V�%v��+b����2]D�&�
S���c�*۞�"�L-&"B>��A��,UDE��+쫿��7�V�{�����1΋ M��$�� �"��n��g'�d,��E-VZ�a�D�yg������weF��;I�2��&�Շug9dם��M*�B�s~<�N�T���|+5e4^��4�'�@剙kMbˊ����D�栞E�,v��FC��܇XyE&M� �k-��ޣ�-U���r����q��i��\��^�s5S�FY�n0���w�ۘ�[�f�݉��; ��x�`F^�3q���)5h`J{�kf)�,�X�3bB4t�o1�U��nآR��ߘ��@^�(�vʒm���PƱ���&���M_���/r�%a�8Zͺu0��6�nP���v��fc�2e��8X�1	7@	�c�Yb�@�1�5�pn�
P�M�@b��)L�[�y-�6�'`&t8�Z��
D���i�Joi���)8�P1|>zkb�bjr��*��un#k2:6�Fh�YQf9��]�ƯkP�B
fL)��4
td*2YZ�R�û.�8C�mT�wV�P�JQ��T!�3^��1���+M��@�W�X)вZ/�jP�.��Dm2�-g+o!�W���0K�l�٬A�n���1Њ`�+(�x ߚV6�b�{m����B7u�lj�Q���ĩ�zI
�p�˚��YW,��SAS(�w��A\zM,�(-�+7k7�)^���Jͨ��ʆw#}�%Z=23v�{���ڷ��^V<h�
�4�J*��L��
Gm�٩܊�^Ѭ�U��if�C�y��Cj,��	/({30@b�L��o)����h;j�-:E�%Y��4.Z����S*Tb�!ⱐ���ݕq�	���Y�Ֆ����y��R���f�]*@��ߚu��]iy'n�}�B@b�а�b���X,��EJԳ�S0ݹ��8΢r�u���ZdȈ̀+��e6nfZ��$�G4F=58˅�2��M-�:�n�dt����s ��7)��C6��[WR�(�cq��g5�4H$|$��7��OA�;���\��@&�-�,�v�I��,�ǕKd(^S����8�� -�t��G�f�� �T�1�z�)�x�[xn0�m�I)�
�)~���`9Z���u:�R��[�yX ��V㙨<���zNne�st��b�b���4�� ß;U{��z^dl��L�D��U��K-�, ,�&�G_\�oMx6�v�ɍL%=`���d�� j�,4��S�P�ԅlb*^ek%����t��e:�Pj`ն^���2V��v3!U-U��(�E��B��9Kv*Y�c�{Yy>�؂�.�F1��7mQV`Cβ���И�C�$����an��U����tR� 19�����6��C��:+$�ձ+���ۊҸ�9�_�p��nJ)2y+͓K��R�*7[f��au\�o�Vt+��V��uu�FwK�K����$)�[�SgR�o5�K@`�<g-Kk#X�E����{R�$3�_]��7Z�y��[�;�:凭�:$	}�m`�fؾ��S�"�ֻ�V&�I��<�6�$,�	;�q��_ʯΎ
��Ϯ���ה�OG��rK���&��N�5vw"6���G���:Vϸ�&Vw,��+i	�)�t��h	�T��kr>ę��+���2<��F��z����0R��Q���Y��9����R�We�z��[!�q�u�
��i�9j[]��-��V����B�����l��m��tI�nB��n�D�{at�B��̡�G��i*t���A]���2����rq��u&m@��JQf��հ��A��mf�o\U����>�s4q~QJn>�ݵҊ�+���5��T��d�m�NӠ�p^���t��U�oXks;�PL=n!��e1�}��cF񰻦S$^u�bƗ��c�5;�"�i�b�u����*�K�Ҽ������o�A�s��I�R�0;L�2PL�Շ��qg*f�P��0]N��W�u}%%vh�*�{B_v�^ҙ ���k����2�ܹR��z�k@�t����7)�꘠Ӽ���75kj�t�Y�����Ӊ�GR	U��9�ǁ���;-iwI�M#�v�)S�)�lf]�:C���D�=�t�_U��+L�@s�����c�4޻-Tmv��]Ju��Y�A�A�]���.�
vP���-��:��Vr8���y������ �ϻ�]s�GSzb�E�.�>���jwԲQ�a:��ke��k4�۬�V-fvõ$-���4C��S�;`[�񥒬�����'���u5�S�:�elV��� �"�)n��FM�ÊmeO1
�E[����u�AJ�:�7��C9��tҷ��닥e�d]�7њ�
nt��
� 4��cʕu�%�W�@ஷ7��hIoc�n�-�L�1�N�f��˼�Y�w�9��mF���z5�֫�J]��@'u�73��Ԫn�HӠ��EN�Vb��F�t���.�һb_H��vc�R�-t�wr�7���u �XFp���Uuoo4�P�4p\j�c�[�dp��o��EV�F�2A�GKw�Y��q�
��w���&t3�I����V5M�
ҕ�-s��٫+��9�2�,�t1��0ƈ�[�˥�Uz�[�6�KS�e�-�����$G�=�����<%cJb�RtZdna�5k��pI��ډ��]y��'�騴d�6�!K!u���e[��<z���)�d�A���/�hwwspЦ�XA(���v���m�&'�c�}�Ӹ���3|�!���t^�mLv\~�����;Kq�L��P.-	j�[o:[����T������MZI�ӬQ
��)nL����9�@[����ˍ˭W/��h�P8���i �};����8"�V�%�����J�����ѫE-ǍÍX+w���GS;&ԫJ�omNǽ���ΩO_\�d���Mso(v��Xܙ�I�����򕆠]w�6���FΝY�^��ܸr��Ӳn�8�oi\Ӣ�@�Fb(�B�<II����[p^�\�,H�v0�HٍWV�E��SP���t��6Au �xG׳C�wV�xz�r�����E[����a�Ļ6�G��Wg%N{�:}J변�ڝ���%�����Ӓ8�i�70j�v�։�&u�j��x�m*=�TQm���&ξ]��#a=���I��$�:�6VQyD�d���X�25�'e�:p��ckK�-٢���bW76��+(v�c���;9�g	z���N�䀘wc�c��%��h�n+%��0�j�
�n�}�n��N��n��vT٨>gYՙ1��1������Vxw�&�߷K��ޜ���Ku}����n����9r+�b6��n���*<�Q�i�ueX��l�v�D�Y�p����`�˙���)������>o��vc�K��[���U���h^�MYYW�Q7�^�w����jI�94oh��d���x_+�zst�E�1���r���6�b�N}��j��{`{��Հն��н
�r��ݪs���X���6kF�U��2�s�:�����Z<G�+�OT
�H�6���<�v������v�6��]yz+���ݑ>zB;�Cόm&���b��i{���zU��x����N�^�͂����j�[�["*�Cp%�G��qO�.dm�^^�ƹ�[��W(�H.��B�r镎�^�i"�+1��U�7�Ws��u���Ӎd���h��ᳱ����X��X+8V΢���uD�j��
�n�L
L�B�ɉld��Jc,H*i�g2^�Ӫ�R�؎j��k<�Q#�[���w�Ue�h�\���+u��ϸ�3��撳�J��\iY��}�y#������9��`�[�u������e�]{I�x�U��^ܢ����y�u'D�5�q���I�ʥ6����yHwC�l�\�/�>��/.��l��U�<M]C�OV�\��2��t&�ݥ�.龖�K4Htp�,m�����y�m-^P�jߋi^r�k���\Z%�N�n���S����ݗ������L�}���*{����o�B8.�9|U�� �.k�K��Y1Ԡ��Gf�w�����n�I8�X�+�z��e�U�JX�uMsw�^���[g	b�掻�P�D�s4�̲e����W�E{���PO+��
��0n�=)[F��6��d��݁$iie1�Sl֮�cp����oqܲ�]D�u%K��)`�9GR�Pz��p�O#�+U���F7��-c8hvW6t=@n���X2��hj-�;0�>=���gYK�VN�$������b�v�H�����ޱ�.����U��=��Hmk�ݎ�i	��z9� +Wf�p>:�5+�
d�U<�j����̚�U�����t纍�ƍ;�hm>�A7ց���j@N�َeL�;h�bh�eHZ]܂aLwZ!,j���N�x��J�����x/�Ɉ�GG:�׭vݮ��+	��L[Y��&�����l�V����A[AtŉXw�hr�9�������B�hA:�F�����mհQ,�E%w]�Uv�<��]�WB��1�	uݘ���JU�r��|5%[Tʼջ��4B[i�aT��
܅|���x·��h��:����0�IG�-��ʵ�8����ap�(�V �嗒4/���.��i��}0��R�I�cz_0%$4"E-9 �rcGA�:����)k��.�gj���;LF���kĀ�u�yQ\s��MMIBH^d��k��@T�YU�,�D#�AeĀ˕��/-����>�ח\j�^Y�"N�Dr����:���K���v�*�9r���7FV\�"�e���tP�i��X!�3	2�宺u9ī�����!zm��o@�)SN��w�D�͙B��ÍF�[�ȷO�a���-��,{�S��Ѡ��cs[[Y��4,ѻat}_i]pX�ʔ��.��Ck-�[x_c�ps�N�T�ѽ�w��8��l�Xt���<�X8��<�h&%���Y�c6�>��ۡI�Q^�}[Cs�m![{׽|քf�9f�Y¹3 +n�D��Õ-N��$����.��)�׏y����H��m��&m"�����C�5b�53{�Ń�O	�=�g�P���l��71�� ���j�0[��+e�ꀏ^h#^��fV�A�.[w`H������"��s
`��4�~i���h
�����b.�1��ʱ��-&J)�y1��-`qml������b����N��QN��|�2�=��ʝ����2��}��N�c��c�8�������D�/*Ө�e�+�'����|�^�+:,���h=�]>SO
�kE�������zgWC�j!9]�
�:�:&�T�t[u�!�־i�5]��� �]nj����X[�E�����]�W��u}-��8`��w2<���s�#,כHrK���Φ�!HM��.�ҩ����l�z�EŹr�UjH\�$[�æ��ݙx���f�woW��<�r���W;�Ȏ�)�)�S}k��S�/Tif�Rj�t��YZ����"ͭ�j�e�P�)�n�Q|ha�}�Y����>��p^�U9Vut*�X\��qL��J).�4D!~���\��޺��:y�ԥN���ĕװ������Ļ��#,ڝ8ũ��z��i�]��3jHo�Y��)��y�؋��n����Y�1�`8�~,�E�T���+��b���]�Qy�˺�#�qMɹ>Q\���{ �fuK�,Ƥ���fg��V5mu-�dঔX�\�o`�I�5�,^�α��T4��+��띎�����[�{^�b��B#"Y!R������ڼ��N��� /����Vk�����hVc�(�X�B��q�p�,un���=�j�aj3J���l��qRo)D�6��E�㾡շ�'y��W36�谕�>���+�K�������M��ؚN�@�X*����ܥ�ȈE�Хl��"wN�(���=����sm�c�TR�ښ_v�G���b��!�fܧV�CA�.�.L��G��V��1Y�{�뗱Q�jJM=��~�R�/
R���J�H:ȅ�,N�WAjF��m�2H/0v�(�f�6��)��X;�����g�K}�
u)��n]QN�a������+ꮑ<<C�<��%�����
e�u�ʐuEs���lf��]�Pd��=\S]�i��÷X�;-R����6Y�мv�l��o:pO�
�]�z���O��#!�D��P
|�$�l�m��!a�3)x��ȫ� iؾ��������Z�^���ɖ��os(��ͪQ��Fb��XT/2_:�LF�:��A�88�v���z�$�u^|-����(��u�K.��H5������sCug��u�c/m�+����7K���-� >U�y^����%����`r�r2`�k�`]뿏5E�O��hIN]k����/�P���aw�e/�#7����̵.h���f�v�og̗
����"�-��Ef�8&�63lk��iK�>i'Q���Կf�tfIy��{��<�B�����h� ��4����Ð.q��aKl�]����|��J�7�sۑu�K)"W\�)؛���ok|�\�S,I9����8�Yw��C-7�ޥc��Vҹ��UچP}�Su��u��*��mI�D/��ғ9����4��j�:��yr�1�G0q��T:��p���Z��	sΚU��-M ��Q�����Yh���T�p���\��
�*�*���?��e)crb��L�z�!��B�s���1�zV詽��X΃��EM��� �p�nru�v�.!Yޝu��.���aB�{��
c�eEը)�Y�d;2��߬oq�ݼ���{5cuc���Z�ej�LJreyO�d;oQOh��}Wb�k��&�V5qa�22~Zp���1�,z�1e_7��Z(!/;��g���)�3��������ޅ�8�/�Nűm���(ka<���p����Ӳ�m8��X� (�)�V��ClX��=��,�&2c����[��ao@�·��W(>V'7���jD]5��q`U���h�i��k�2L�+M�T$:�I��V��Pz��%+_]�cI�E,׺�TЮ���Q�w��1����%]��$]���-U���N.��k�����,|�%�x��)�슜C,4��V�ۙ�gR#��^�4�GaވT���dB���ջ&�^
vl�ˏ4Ў"*!O7���B��P�7�'�����2�wU��Z�XGp���@ث5��9��wz�F�����,1Z�}f��ձ�_޷}3�w���nc���m��ޔ�i��n�s,b��9"C����˂�n^G��i:�\��wr��S�/Y�-�Gk7Z�dG��1�D�5��ZWz�'G��w�-һ�J�L��ݾYVd#��p�vF�L)�R1un��ʵ׵�R��eEv��9���p���u'@>*N��k'\���D[��EC�
Nw`3i�{���Ӱu6��I0�#I�Ʉ�c��N�ʴ�6��J�w�c�˫[�غ��e>E��3%t��w,��t���sZa]���Ź����S�3��}�3�aR�/�;�s���m�V"wN#c�K3���AR_Y�R����]hICw:CώEG�g6k�w[��Q)[6� 'W
��1�=m����k�#�y`Z�t]�m!s5�tK"�tbo0;�TgnCφ��;mu�v�B
J�t�z��v�"�v^UDxK��En�� ����nm��l0\�u/��T���
0���(�t�e��wzl��c 
QyL�-N��K��ִ�&|��L�VG>����q��\��GZ��MMV�:Y�kڌd�ҹ[����8��f̎Jʬ��՛qMǖ�M\ӎ�r���-˾���ѩԹ�.`��tvvu��{n�0r�#%-�nb�u�����|�gf�k=����&ۘ� ��JvÉ���s��(��o-Yj"x�3�eIv�5��wL���P֜�����K��:�v�s���P�p8�]��3���2�^�E����1#2�(h�����Z��ג�l�n��n	�Ƌ]�k.
۝�.�.��ӕح����jy��m.b"t}�0��ڴt)sn�q�0��Pi%-z}�~��&)�4^tW+�ޮHI�:>Ú��U�q�yF3��` So�I��m\�K�V5f����BO;y�b�5����5Qxfc�iU���*j	��q�-HlC�]=7��f�*`�u\\�eW���HHHRB��>݀@/,$$%d�I�'�@���H�`@�l�	����H�2@�X6�6�I8� 0��I'XBq$RHa!0 �@���a����
�dĆ�Bqzɿi!�H\� i2`c$�Đ�$�`z�*Bb@�I=��$1�1�<f�bC�x�<@4�CH���2bHH,!5�$<BM$40����a8�m&���P6��R��	�����ԝH,<aĐ�Bm!Ԅ� �ꄞ�<HL1!|��d��HN�<HN IR���$Y1���$hI���v�&2Hkt�i	�,�f��!6˫$���8��,$1�6�HM�k(q	�"�4�d���&�IĐ��CI	�$*X�� �� �Lf��`IX<��HV���@�$��@��Ad�IR���񂒰��:����y@��Hm��Ba&��7��Ci�
�����0���I� Xm�<I�@�!@0���k�Oi��R�Vd�%E X6�J�IRY���Ld�	Y$�H]�*�i"�'�&�ǞY$�)	�"ȠI�i��Ԅ�:��m<dwgRE��2�d�`�a�I/(I�I��Qii���'�8�=������ȡ��2s(YCl�Bs�{���HjB,�bL6�0&$Y$׶@1!���1�<v�i� m �`ON z��4�L��!�$P
�q��Y'Yܤ�[ ��:�Hi�:��8�u�I�!�I=a�����!�k)n�y`u	<aXd�Y�PEo(q�P4�d16�l�!4��I�BbCW�	�)<f�d�a�{d+$:��yI:�N0=�`��+򆓨C��f��!��2ԇw� q��0�g,�@[�	P�u��w���@�q�Z�L��َ۫`VJ�}�xԙ�d�l�Y$�+	㌜J�<�8��[���h�j�NyC�Rm�'�m���d�%|��=|a��l�
x�;a�T���5�I��6�r�{�7����Si�ݡ=���x�a��یV��d�I]����0��-��y�2���L�bT����P�����1���09�OyOS�S��&�`�����u �!)���s�R^���:����Xy��S{��e�*#�'����;a�,:�w��%���k�k��/-�ksYZ�"�'��S�g�������z�8YG�B����ix��:��H���[���}+�A��+���`k_a ��C4����mcCɝ���&�B `���E�l�o�(U�4X!0p��u��*�(&�������2
���b�˗�Ο�h��k�ځ�t�P/��Vd�T B�a�R�k�����/�;Бu(:Se�Ĥ�"ra�]j�]pƅ����C�7���Z�<w+6�IA
<pu�:�l��c��IMJ$� �AP;Fi)��ӣ̮��Y�1!�^"#�b����+ש�^`���������	�u����d`��9����y��W���s�!��Fr���6̮�TP�\róJ\P�i���s�t�G.�BS��>$�f�˓���5 )�p��k�NZ�*��R�9�9����FnV}��1.�� �-l=���,U���}bPɩ��	��[�u�m6,^u�"A\&h�WB��\�D7��d�UQ��1A[`�A�KW̮T���d��B�&�1����X����l�wS�Y�!]9��Xb�Y����vHAMQ�����Y�&��j�vz����P:�q�38ݮ*v:�BH���B�i@��w�iq�3f�����N��)�F��΃�*-�6�q�¹�=\k@X�E�e�Ĳ��6U��iꁈ(�ۣH��y��DF����n�-��!�a&���Ӳ���Vwȕ�f,�w��H�Ǌ޳�Tm�*��?
T�֣l��O�������PV*3YpvʔZ@<��	
�cl<i!M�(Ǯ"0����جAչ���u�$�$���=�߼4�{��oȅ#��J�l�̗-]�[C1���ͥ��oP�ְ�WΚ׻w�.<<�gN�;[���D�uc?)���gD����gm�teL[d�YȬ�(�+z���_�G��1��2;fT��V!۲�wJ��X.ܵ�B�Ջb�>�ym���tU�w55ـ�w�Eų����r�+�t��>Ór����Wu3re�}�J��+�m:��/M5�ۄoQpY�.u�v�]�� �)���tXn:d��f�]nT�8f�O׉��g���ơ����ռ|�޸��].Z���J��]�.�g	YA���Z���'1�h~P&�%�Y�C�8�|���j�Gw��]CuQM���}k%�N�֨�Ì�h,�X���k��P=Y�Z���z�W�(��(�� 1�e�����e��t����ьZ�%^B����{Dr�ީ1��ˮ;2�<1��c�3��[�j5荧 ��^����#��ݔ�n�Gڕ;��>�\k�ѻ��5r�>;�,�4�w���8�yАrl��t�.�
�v�������m��>\g!Y�6���}�d���r�E�W@↎�q��u<���^��/��E�L�)ʀf�r)�;�z�Y`��$?bܷ�Futy��\0��	�p���Y��0��s�H�w����:յ��{����^��� Ir�~g=���5t�ޞ��N�VX�d�����0|=ZU���]�V����r��u%���ǅ�ju6v_Ԥilή7��ú��LHB��4�j�m$�I���&2@i%BC� 
�x� �9�LI$�	4��HT�}ޠ@� �
�4�'�	4���n�M C�J�i�T��$/�rI	R�$�0����Bi�����߸���s|��}��7�w��"�DAAm�;B�QE�
�"(
ϒ�DՅ"��[E��N}�DDb	�QTX�I�(z�PTH�TUSIY�0AAV�A{�iEE'֑E"ŋl�ր�b�.��X�5QEb,��b�#1�bX�@U��DX���#Z�jE��+֩1�(���,�(
�� �V�V*�*��X��f[TTuJ
�����A�jlUX�O"�"�G>{���TTEQ�U����AEQd�>Bg�1�Fu*����19J��H�Yc@`�\aLJF �+�� ÍQCt8�"�E�5D��DQb(�Pb�EQYOm�"**Ȫ,`��>4$�H")$��6g��g8��=��o�`!p�j(�X�*�b"1ED�����+\�Eg��PЊ���wo֊*��b�Ɗ�DE�/�U��DE���TPT��QU���~͌�P�P�Q�±AA<���C�i0b�V��I*�X�Em�g�oA�Z�U(�iDTHŌLj�E]Ҩ�}ϳH���w(�Q}lETi�cUA߳^Z��G�F
*��b�eX""}j���a������԰G�Q���
�%g2���v\j�URV�KlQQ?�'�@>��Uˤ���[�	6f����g֢�1DQ(媨,�@��>oF�DT`�"��:�"�#�Q���,]���1V*�h(���/��B���b��Y�[Lʨ��QEX�+�YQJ�gs���;�T}�TA@�z̊�D3)2/mGV��*#=��L�p�{���TNRX����Z�ENw�hڿ%핂(�
���"�QD`�&��4�U�������߹��a�)�����>eTF'��_m}s�{|.�y�]�=�o�x�f���(,byj3�Aq�%D^�4��(�V")�TUX�A���4'�}B���]�
�+(�h)��*�E"���kIƬg�S�*�b��T=�V��(�-�Ȫ��r��>��i)T�Q���QD1*,�C��Qs2
E�������g�"9J,DSm��AR�LQPCMA~���TDF1��V�e�k6����K˝�$���
�QUݠ�)��d�)�
�("c%G��#���mA�LF5b)��{��|�f;q��TcF��QMZ����
�	�fJ"->l��U*S�VLaY^���Eբ1b�*x��A�^o���p)�U����z��d�\ȪG�*��<���7o��~s(�|}���Nv��5rDlfkӳZ��ު��QQE�X�mR6��Q5lX����Ǝ%�*��Q5}¬Dr�X��{�̲Ō-�S�C�Z���جS,��[��c=ʊ������)23�����3v4�m
(�ϼ�㵊'�ED���o�sUDF*��,�EQ2����nr��(�$�A�ս�Ub\{��}w:�f�oz��!��I���   91�EE����3�Q��h��Ȫ��*�heR��N�X��B����̘�L~uEr�F�%pEs�	�WMJyL�D_|�n�z�_�m��l�-A5���i�R���*�rՋ�Y�K��5a�S���N���!>�,��v-�n��	!��F*#�R+�t�o�ǔ���#E��z�"}���,�H����w�5�0�ԛLU�y1�8`(]a�i_Y]'�sVS(�PU��` �h����6��+*����PDXԿR�����g���P�����>�TL�kƣ�x�@$�(bDw�^�����U^���>�(c`�o���zu;o�LV[p�}�Q?'����y�a̳�,q
�,K�pQ|�C�����^淺�+[��orW{�B&��UU�WM��a��r)��("9��*��++Y�Dc�t��7�
�&��PR �!����4;�2�0���Wm��ܾu��B�$���0��{IV!kݕ�8ش%5�D��ɀ��`8�^60��h�&����$v� 7'a�W�Z;C��7�={߲�o��|g!Ʋ�ms�����ܽ��@�L}/ͺ����}]�T��Y�p�-�<��EY�Q1,Ew[����(Z�����UQĨ���]f��Q+�g;�=x,~�/�����7�����DOmue��LJ����a�h��x8��q��T�o^�:x�bQEb"[�����}η}�����׽]��I=O�* "�?I)Yd��h4+f�]�X�.��컼�F�Z�iDT<qG�OYMjsRo+�)Yx�v�ݾ����3%TQ�}ֹJ��\ʹh�=�0�Rc�T���n���/ɤQ1(�n�����<�POw�8�͜�^�K��ʿu�IM4� �	�Lo#������R�ݸ�ՔǸS&O�(ie�4�Ko`@�	1"&����TQ�,�F+l���W-M32R��!y߳��颉i�׬�y��*+~��e�n�>��k摃�K�Q$},%��H28ʜ1_�����ߕ;��c��0*o�c�E��A�
�	���$��ʮ�Gd�DS�]n�ba��Z�,�y�詫�*����h��KO9��n����y���O�v�_��Z�l� [`ɐz߇\�۽cXUG*���^�řĐ8���_`�{�����+.�x��ܬ-���4s�DCV��L5h��B��QQ-��w9�c�,�ES��hٯ�'��0D7s�w��st���6���L�R�E*(_�|�{M�`@�A��;���\_��3ޞ�
�unv�	��a�⁴��(I/�y�J�}�DĢ6��4c�l��yh��>��qSt�3IB�(��fk����MR�5�8�eM7mA��Ճ�n8ŬR��.�v����iFx�Q��3VQ:�������8�^��n�7}.��Zda�#̡�S>�{=�~.�+T�Y~�@�T��6抪��9�����w�0VZTv�<�'���T����ոU�������I�\��v�q�Q�4���[Qw�LUo�}��T:l�4���W�I�,�4}���Q6=����I���z/��Sl�Ot����gfH~4B��� �)U�*���i'u�]$�+ˏ��8��� �h){~g������p�IK��$�R�Lb���㥚�r��j.���6�sЉ- ~"�@Xd�����05M�6ǔ"��l�ݕ۫q��nZ�źt�E�M4T����{_���$5E�F(�I|�KZ#�y��݊��|̋��o��R�cB�n��~�T9����Lk�9t��~
�r3�u�tp��<�Y"�[�SQ���U9�ͧ�mO��_�ڋ�bf%QAo�>��� �AE����|e(C$�FT����@�����R �/����]� �I�Y �[�;���:���}ju̬dҬj�oCO{���n�r���+���U�۷���Ӿ��R����r��d�4�����Nd:+�qE�� ��m.����n�R����6���E[�2��Ç'd72&�yY�Q���<��[�<�S��5Q-Ø�i��,���rG������I.n�Y\@_�D/&iT^Y�`�J���S�̙L�Ҙ[�]4�cl��}�|�T~�1gs�4�鬮��N�/2�'7���ʰ�@���xp93�'�KQ�8�+�v��"	����@3KR�T~�"	��#�S(�$�v&Of�P�^�?Xaq�~Q�\�--K�F?O��Rی\q�[�}����Z�e���2�D�@����v�ԛ������2�>~�T���}w���_/��A)O@�U�r�H�:�yh���}3���0(�J��^���VH��ނ�B�G�U�}E�d2h��]T�D�-�A��!'<�U|��.Znُ��{�9� "�!eDnT6��ە(@���|G�@a_X�sxQ�)�q�mXu���u5ˑ����p�{���7�ٖnA��#�g�C�G/Va�g�Z�ɖ}ճw�_ ��?2T�!��"�lf�$��@JT��I��Y�+ʕ�Nm
o�QA2��ˊ�fP��>K�U_���?F�G��w�v���]��bJVep�{>$h��@@��nk����U��;}ߛ��
�N��Ƹ���I4�-�>T)6�K@^@S].�'�� ~"TLQ���m��q|V��R�q+Lw�Ӈoƙ�X�@�����d�io���T:���%�蹡(��	��_[A������8��X?c�%�0*����F�@(h�i�P�U  �x�Q%A���jYGK��1W�"e�����^��Y���?�����(f��ȲJ�Z�P�7oT�dY\�0����I��evԜ��_����
-��q�ۿ2n=j.��ɿ�!`cHP�ᢞ������2�SN֭7�j����������Q�I ����tĚi�	"����~M)���A�s���x�SC�2^'ڝn�9�^"�4�� .,�+����	��p,=$�U��葮�ʳ��@3�/��^̲2�B�#��q�@S�Vh>A���7:����"��)߰4_��~n=���!�|9�"DRKٹ�ތ�Z�ͦ}u�{�'��]����[�\7a.�F�Yٶ��|L�n���7�/�o�ǳ����q�䬩�Τ�o=�ʚ�����_9_E����IM�ϮW�t�Ֆ�uszp���mW5��	�#k��K�i���X����΍�{.ݎ�z-�{��/Q���T�>A\0I͕ނ�<���ad���?.l"������#$in>_8���W\"�|�/�"��H�K���H�O!'�������Bo�[�Wu��ם�S[�88%eZ�%�w���ّq�Żu�MS1]��7l-(�"�4^���	���vM_�����m��&q-O��w3��n�
>Jl3Mv�r�T��=V��
)� ���'�R�R���?!�D�5�-6����l�J+�)"� ��bA�~a��#a��=V@e$D/�ȑ ��6x��k�s^r֣�A�f�_���KZE��#��:9G�j��iλT�|J�{���R��gmq[�*�y��X��њR!@���S����.�z:"�)���f��Uk~9�����NĪ�ǩV����%�BB�(�l<��*6	��D�,���F!$�qC!�Ҡ��%�A����
|J�}k�7)O	�=+^t9f��wқ(�%d�K���]�I��_���D4���eo��:��G��|h�����*�l��9��̅w�E�����
@x����`�WȴNy.�uxЭ���l�gS��4B��.+?2���L�D�^�w{�� �-Y8����"6�X�%{r����mC)Ӄ͈$oW�h��=����J_����� �C~�}J� �Z�*酇�h�#�X��钾��<Lϫn[�\n��N��6����	��\�T����}�v�Lx��W���É�mdlS^J[?�H�H<�O�h��(�Iԍ/�y�/�&~�vN��K@ϮW��A|EQ��$�H�$䝱�&���j� 5!��y��z�	�0��zNWUQņ@��wK�(�Y��C�)�
�T�KRakF�g<�y�"(5~�Y��^�Cm]���c������}g�H��2Fw^�&w�;
�ٮ_j�''J@�uyb�W�@�v�Ԣ���6�2�q,-y4�A]1��Y�v�4�h��R�u���}E�,T������A������N�h~|�:]�Q���u±�W�9�\jl�Zz�X�7ږB}�y������9�:�e�L��� I mN��A��z�/�4�m#z�^h�0~h"Q�s�#��?,l4�|���u�j>]K�^W ��Y+;)��H0�D�/R�"Hy;�SR��xV?��1!��/���"�l�*Q�-�I%&��c�C�uC��`.k`L%��C+��
�)(�n�F�ȩW^����إ!��haH�$��(��@��x?J��łM�ΚU?���R�&/��9�	s��+d�c;�J�B覂�����A~�~�g�Q�2�j��y7V)ȂCS������tL@�4!�~��(��1p�`_��G�Q�M��U��C��H�T[��O���i7�q�� �M$�����]�̩έ�y����ᥟ�Y!�$��[v��!}ɼ<DUG�le��#�o^o��fzE]�J�
�+�gc��e��VLV��z��yٓ2�o��iNѬ�g/�ܭ����W�:��6~�[��qO�'1Qt���~f��i/��-�����P�C�$B�����Q�0�F�ck�^�[����ء�|s���^������e���#W�U4�4@��YM���-2*��z��nO�����@��(7~�l��!�UŊ�9�x���M6�h�3��%�}�X�#[<p��g�hV��d�Ɣ!> �>=O"<�>H���룞l�QR-��}͒I����a�����x�u|�[P� �Tp������,�-�N/�%�{�6�_����-n���?2�Az�zs���2Y)-���팽8D���GO�І���
�ȒTX�q�+��V��r;/Mx/�<��I8�8ƾ$�{�Et�:x"(��{��[;�Ȁ������/�>�F"P�4��_ (���N�,�ٕn#��X����BQ�����o��j�(�sd/�Z��xv���Ɨ��8�E����C��$�q���߽�$=��-�Ϭ���/�os�$��'�����+�>��l�冼��}������$�0��d��w��s|4@4�{�k�x�*�J�����_RO*���Mt�3e{��?}Dn��`����`��aTmԩ�Mֆ�L�%9-�d�Z���CX��Ћ��eH�7o���'�5o"���=�|�ҏ�﷥�����Z�P~kP@���"DgfJ�p�LHn('п'>��-1&�Ϣ:Ʀ(��7gme�b<^��߯�*�q�)����K���k'���0$H+;jJ%@�!1��/:HP�M��Vi�O���:G���#=1�TQ5�!�}�?�]#��������J{rVSK6�Ң;��{鹹J1ĢPA6��,�Ӛ����*�uH�\��P@���}����������+,���C��$'�� � ��p�-�֘xW]ݟӞ8v�i@���ԫ͐��J��:�y��q�S޶&mq1�A��}y$UͰ�X�1���]��.��D ����v�����(ު�z�������Er��Z'�J:F�n���e#�(��v6wS��b
D����vP%}~�5|8��5�˼����l%����s4����pフZ�.�+�Pu�e���BȌ��b� �+Ņ�������@$�Y��/��΋��CI"(��z(��}v���6�몎z�]�ݵ3�L}XK�k�GE���C�q1m�-��!�R3�G�שRX|E�(2�ny��L��^o�ϥ6'6B?6;����s�4HK���K��m�M}�mU���I�暚�?��f ��QL�`U\hr�8)���2� �c�2�g�4՜�X�_F�jqЬ��$�`^��,�<��Y�uy(i�Qʱ3UM,29<Q��G��w:»�f����Z����U��2*���^����Jښ,���/ȏmxz�&=�n?<��z2n��~C�� �w�{�/��[]��*��db]��e!ޙB�<|T��O��$�<�%&�v`���-�TZ�M��n���f�-0���o �s�*�\J��at����}���!���Hj���!�x`�H[$�N�����n�_qw�� ��Hs����әwb�w���9��n�\i�V�܌-g}*pe�ѰrS��}�| �a{�a�������ר������m*��oe����A�C�)���o��P�������ᎅs�eK3�����s������YE˷��Y�{��t��\ݯ��}�q�z܈����n�Ai���؉,��pA�Uv}�z��	H5pNU l[C����>T��R��y���f�LK+�W�M�ˮZ�b�o,�CIXa��e�LW˘���\_S�Z- �B��Uih����̱,�Y�1@�ûU�L"Sd�i��7~c7z�$U[^�^r�ܡ��ؾ���D3��H�A4�9$U}�V�����㢯�FD2�\����
-���p�~�)�)�P�T��b�T��{a�6�_�p=��E���޷�A� ���'uuCH�E?U:��$���1���e�+�8�CQ/�zUD6�i�p���p�=zǂ����n�5�g��Fk�'B��vD���̉eL�d�� g�j��a�_�P|Ӏ��z�Ȑ�I����E2T4�_"B(�)ʞm���ڥg�<���uvs�0$E%E,���b�s2� �t����T��f�Ǻ8O�hzq �εts�e%r��AN�����\�\���xL��̾��Y/J�n���ʒ�z�f�y��H£��	�N���Z���b)vu�$z+3����TC,�����.����OY���S�.fr4e��#~���H�`����b�v�8�V�v�#RC�NZ$n��"�x>���B�!C{B���K����* �_�T[�� Ⱦ����s�w�2��@=���
3^V���7���TK��[O��6Z��z��U�+(_Ɗ���HZTrB�r�؄�e�P��ܢ`4����x݉�g�Y�B���	wk��@�oL���ע���L�F�&�X�AB��{R?g@���1O�i^�K����ua���a����K&�S�S[g��R���6��������n�߈� |4��Uv<:�0l��x�������zQӲ�e�}�ӽ\�:�]��nt1��w������$^c�`��_��,���l�X5�
�c���F"�d?O]K/�fx�,-
^'�����J���(ֳ���M�d���6��ٌ��z�p�;nm>X~�B��A 򎮻�L&�ѷ�M"���E�>^��P�	ІG���E���r��A���+PMcMd[WaYF�_��88�ނ�{ҡ�ٔ8Ru]X�WS�7'A��Oq��ZTSD��i��"�tlOd�CC�*ƀ�{�t�,�B�U��N�1��fy\}�y��}{�`��AM����R��dA���\K��o��/�?9_4�
�x�p`EƘ��f�wP���Uү]�@B���d�xv�==��Zc��w\�b{�����!��G���v;�b���Ή�F85�Ð�M ��t}�B~e|A$Wg�P�SK9L����U���/�ͭw����1٤��pU�Q�H�=�jȴ�(��!nP�e��I��T(���f��?8���ʇ'H�<�t[������Lq}���,4�Y2'^>��.�,�y7�ݕ�7����-�:�qvu�����8��Vؔ����فP�]\�.��,hcI*�\��G2?PW��;Q�[�-7�Z�[Yu`�m��@����I���&(�5����ar�(�Hq��l��j�'ͤ@`�����(�SU��4��|�6F#�����O+<�|~��,2�X�ha?�?��G�y|AZ��Œ����sz~�ܴ�p�
��a��+Es.e���^�4]�p^q��qbNZ�r���(�k`�ŏj~ �g����T���4mf��+o۷`S�167��+.���/����p3v���u�(�zD�r��s +Ү��d0R�^�a�Z����A�}%��q �F*���'�P"����e���7��Ȑ0�g�R7��$�4A��iE`��7;=k��AuNSjJ����kT�][y��ڼ{�íK��rhZ�q��l�ۢ�MXy���u���9;v�"1q�����B��{�Ur�E�K
�K�ř���Ke4
����5է[�E�z�a�
�n�r�
���BJT2v>���f��㣟��Dx�lYg��U�0LI��F�L��H���3O�eA&n�r�]\���Ϸ��o7�����[J1��N���*���g���I0�g�[�k��ʿS���/�M�˧�+�X���#͛�FRe�C�&0�P۬�L��ʦ���#JI�>��dc{̎-�>��/����L��={ ~s��N.�����R�;�uA�dۀD�뭝�1(�6���}J4�G�MK�~�T6�$�>�!���
��7�u�tl�����Ks=mm�m�x���1kW��&���s[��ug̯qH�]l�0�����	cB�`�P�O�D`ǑmH,��\ C	��͡�n��$=�a�����~eQ"IRP E��L`����L(%W��e��Yڒ�._?�m���nb��n�k⺶�r���g��2�_W0�cQ$p�y�����v+��M%���c��F�ԯ%f4W�d�R)�=Vh��z9��QD�'j}'�B0��Ӣ�5WE�5�0�N4+������ۧ=�^��l��.�?���C�����"i	yb-�a�0��)�����3�F�%�{6�	3�!�ƼEm��hk9������N`�#�����=�YgM4A.�d�G
�!#΁8�B��3��h����P<���������R	[� �Y�t�[M6��s��٩��c�	�LDś�t�	rݔv�CƂ�ȫ���5J� 4<jx�f�I3�E��cO��Ŗ��$\���l�Eq��o0v��fS��*��'\>!@�g��4�4���^; ���D/*�a-#<�e���p��\�3�<��m�˲��gԛi��FR��(�f�X�kfx��0�e9�T�E�Ќ� �Y3qFtV,��`�㋥�Sib��eڋ�k�՜U�R��O�_[�yqq+4���º�oWgu��WQ=E[��Ѕ�}�mt�#.�S�oM��׋�|@��+���pϦK]ʷN��vwRq�"����|�d�dͨ.�z2	'���A�������h��6�Y�|�,i���~}̹���gZ�P��h��:�0{C�TEƁ�P	�0yk�;g��)$�>��o�J�x��G�Ī'^�[�]��w�]W�'g�M�Z<#�ۑsFG�����EQb���o�S+��?z=Ҝ`�iuJ�D��D��u�w�G���wI��!l��V�:����.cޞ��I���]�m���0�B�>,k?���s��0�w@���W��C��W�H�=�`��p��J��>T��;�[�x��{�޾�^�^��C�n<���jr���R6�w���E�t�ML�s� �^0ƹ�Q���l����3%B=�]1��5�}�ڙ�Z�Ȓ�51vN߹�������\��b�XdE�K��8���EF ���|�	Yn�8����Sd6�]�9H6�����[]tH��=������,�=���Xm&���J0�BOT�����c���<]5,�a�5��&�)�.4.葂�
 
�l�w��p�]�tIT�)hYN6\��6a��@B^���y
Ƴ*��9����|`��ثAi�k��R4�hz�(|׈@]G��dk��W7n˺Q��I�d�'�r�Ti�9X$#���T	.uW�`��ζ������(+-���_!m}a���	��8�eWd�c��:1�0�˚�����@�$�Xо4 V�R��+	.�6�O��?(i�uk �ȴ��Y~�z*y�'��߀�e���Fq�4Z�i�7�YO[��?��^�.�Fx��.����t���*��q^0@��� �u��_:���F����G�#�K7����K��E���Έ�fU�C�Z�JT;9䳜���;���7R�d�Lh��3CIf;��ڵ�����hlrn:��R�:gVtq����Y��w\��w<J�,v�)oV)�{��X�e�c,kۑ�ڌc}�/�qS�
�h5���WZmVS��tN��q�F�
y���!���b�����kP}��&�e=�/{���6�����a�]���D�P���n�Yr��ڈ����J�N��{]�-:����7�7X(YO
S�˕{��RR�@<UoB��tH�R�yN�z���
�VsufpndU�3&X3�<�'x�]&�!�[�ݰ������9k/4�Y���;�����X�v�z�"���Un����u��J�o�h#�x�ƷuN�\�0���K�ܠ�w/W[��;Ԣ��{�kZ�ח1R�Y�+Z��]08J��k��
�K��V�ʛ�D}���<q#N r�%�.�µ�.�ݭwl�+p��Rݓ��'{��3�j;����kX��B3-�)��5���om�%=ef�{j.g_)�u��r�>��[ϴ,nv���/`�����΅�o/P�b�u3Ɵ6�:+�i�ڝ�W|]�j\)qt�cΥN�8�icy������2��D��T0[�w��$���P�wee:}�Js�=俇x���y'�;�y���Mmtr}��ZZy'�(u�����X�i��	c����&����ݪ�[�N聭�/8P��"S�����6_pZ��-5 �S�Q������F��v�Q
��0��Co����T����)_W)B�3�[�w�X���-� �*�����1]	�<W-�����g�7Mb�?;�xpe>�"�}���M�ƍ��+k�
T���nf_v\鵠s����Ɛ����;e�Gz��[hv�J�LE�bYΛ��Ki��@���o�nZpc��3yp�z����t�Xޥ/U�8/��J���M�Ι�P�U��^i4-=��T�Z��{J�8�A�d��{yHq73�j�����]�k�wN���1ȃ��⺸�f͔eAfc�YMm̱�Uo[��Ѕ���4�=B�J������0eN)7	r��.��pa��|5��r�cL�D�x���q��mD�weg(��8�;V6��8�8o�pj���L|�+͋C�x�2�<ܡ������mrw�ѻy��s�9��<� *����{Z�_k���m����!ʒ��Y~Kںn����k��rK��<�SJU��ӫ�s�1jI��V9XjFF��J�$�>� ��ꭥOw�W=YN����,�(^�A�� �V]���̵��0{��2)	5�C� 0�Eٳ}����i#n�J��z�ޅ�L�7wo�����ЂC(��>}��F�� �~f&��sO�ڳI�Y�/��K�ܜt�j�=��i=�Φ��l�4��˭wSiOԦ�M~�k�g����gL���}�冹q4�3��9�3f$�iub�
���<���Ԭ�W^~C����+ѵ6;�ֻ��7>���7��t�[1���kOS��Q�����`i:�C�=�1�9p���8ÌZ����l�4`�[�J������DE���3�ti4�� ���h�~���_3�!��!ӡ=�5�S�r�a��?kD��3�m�)�a���7gP�n�㙸�0�y�
s噑�K�玓Sx����kw�g�M�q��g�a�l8�Ң�j�y����?!�ĝ�Y2��5n}��4�f'���CQ��T@'�@�SJ��-��fZN{�
�M&���º�{�m��"��7��V=�:�;�����2C;���7�u���FAE��ԾP�4�a��q����];u�E�\�5�4�ʋ�)�I��Z�����Dy�L�8�yLE:�>���r�%����IF�WT16�~)���M��#���R�M�1e�*�~׿�H=&{3UT��OG�=��O�{ݦ��|a7��9�Ӧm�o��7�(m7��G���bqyN���e1+W�~�\���4�3�=�}���'2�SL����K��u��!�O�u��̱�٭X��@�P�.���g�E}�3���"�3?gW��.R�x3����g��p��+����w�������6���:������ff��Z����)�ۧ�Y�m&'�l�����e��]���w^�S�Fu���Dh2$s�	�G�E�!������~x�E?;a���Ԩ��<Mw��i�ֳY�[��~��8~���.�M ��y3��uw6u��W��������7�37���_i]�B�M��1��1��5f5+5���p�N&e��hM!�̯���14��ݟ4N����Ǝ0��=�{������]�4�՗�s_��3���'�����P�uٖ+�c13}3|�����߿>��<wv��l�HܯѪ�S����#�@�E�~�^����y���B8��4��g�w�}�{�R�橯iSh�o_uw�bj�yE��Zg��8�y�ܤ��G)���ѷ�M&�۳�۰�֐�(���3<�Ɍ���K2�_�us���I+?+C�������;�ÛM{��~#���BG�>��5�
E?3L���!�ٴ8��k��sf���LjWYI�i��s��Jj����ϴpI����D�Z��t���Z��SW3L�~������˫
������6ʋ�������
m���O�yFt]�Kn��{f�0�fm�g�4k�m��*g�����N��N��9�`�䮙����'<�Z�g�sfى*m⪉����~��hT4����f5�M�����w���� �/��2 ���O�i��d�e&�E��Pۦ����渞jǼ�m�g��I\�j�i&��Em.�{\2�CsG;�:6�R��%��*�J�{�:��}��Q����2�6����ĩ �YsudB:�X��lA��������39B5�`Qo6��;����6`�����w�>������g篺&�c�+3ۭP��\�\a�4�{L={ۯߩ�(^�fP���f���5�ϙwc�`��*s)�Y�\��!�z����N�����j��x���阙�/�z�ϰ+4�2�t�<f�M��ݫ�g��[��}�*X�)���ӏP4��-�T*(�h_7�޻a��י���2i��
T-�q�y�:V�a=|N��QDJy��A�(z�*_0�l[�ך�b�d��;�4~����𭰇XQ��bm_���8�R�L���E�jb/���9ϰ�K�7�����L��t�����5C�|���3ve��5��4��l8��no��*<���5G����~gS���g��������?���r�v�`:�&�wG�Ղ�C�tO��*��),U@�g�st5�p������'���įw�Wf�u&�B��{���8�ݦ8�!�<¡�Щ�R�}���q8�
�����}���M0��q��<��+�vg)M�Z��2��ڛ"�
�}���vH��Ϸ�a�s4E |�g�,1���!\CV����ˣ������w&��/s�;ٮY��
�4����q'>��=a�)���������3��S���i*)�>�����۴O J?y���?q�B�D"�4C�?l��!��n���'�9��w/Ҽ��}���E��E�s��~O��ޡ�i#��[�ѝk�Ag\�;��+��&SN��z����a�ɴ��~�)�G��~!���� �dPjb��=�Z����1U<n�3��4�Ģ��bq�m'2���x����l�hO�㻬������G��S�)l6�8�z�5����iЋ1�����r�in;N'�ķ��y�׬�f��!ns[f�S�bO|��7��I~�fR��'�i��Gΐ��@'��?� !�r�@!�g�]V�V}�����L���J����q������4����ߵ���f���i�3W�=�&�_&��q5��6��[l=q2v�m�ִ�f����i󚿽��4��ڝ�b}܆;M�S��\C�g����:��BVd���ZC������|�������Hw�3�잳�%�i(Em��`��|�����>�n�|z�c�Lg亩���˦Ŭ����f/��5���`��4�8�J;f��J�ַ�ˮaS53hiӇ��C�+��֛M���G]}��j��i���~�M��J<��8���7�/��6=Q ޶Rd��Q|�P:���"֠�+
�ڈ�V��#�E���u�4�[�i��?5ײ�c>qh-{�ȼ��}t���A�WS���N}υ����x{�f���9i��C��zFf�[Ѝ9���r���A���me���2��S��@�U
6��v�:8�+ʺ[b��8^'vQB��د�X�݋2�A�+G	˺P�pN=^׊w���i������C���pÊr��;c�]L{+o)_Z�+��9
a��Q"�zŇ��d��~�8Չ.s��m*��C�"yQ��9��ԟ���ٱ�dL��yii_�1H�u� Ea�'A�t���=�ߵuַ5�6��0��v�)�i��p��,���X�>��qluH`��J��#��u��P�Ix�@��ٟ���U~���X׽ �ʥ��$Hb�H�aW����nǰ�x�^�=)�q�ei�D�Cb#�/��_Zq��˝��=�-���{~�Y[Z���HN�w%ftlD��[�4EOƫ�Dƭ�7�F�6�����.�n��Vm+� }�;��%�$g�f�n�G-��uGJ%���=��ǈ�`;>�d���םl�D��R
�p��t)Z�z�:;<���7}��a���|+���^��<�]��7U���r�j�Y���2��
%���
���'8ڥIf��&�]-eH�ܚ�7���Il�=�L3z��) ���W�����?,�0����輌B��1jNU9����fZ�T.���=��i��i���7.��*���8�^Cn�|M����7j�Qd&J�4�KE�"��z�! ������-�4�9"z�A���[$�l�RK�(�˫��Z}+}�R-a���6�s߂t۲.�?�-4��T�%�p2�2!�n�J4�K_.vvݐ��ww7g
prq%�?w��l2[;�,�씺��:	��ˮ��|k�'�i��q�ܝ!uS"�]���^_-�.:�߁!�mm�4 .�iv�nA-��UҠ9����)�������q`|�����Jx�^�ΫįG)|�p�v��f��lD;���2�-&�;[����tJn_>�]#9�_��nX�L��(���]�� ���*�X^�z]��dv�(je�*RD��:�� Y[���z��A�/i�ovv���A*�w66?iF���UClB �A��I�!���3��(�iz>��~�B҈E�r�,��臱��v��=��Ї�\�bt�9�K���w'��	e9�Y+��>�<�R�x7�j���*�l�i�����MN�'�N�掍��,I�Qd�X��Mٯ�¡�8�X����7ؓ�Q��s��6����IkA��F!pn��M�r���y�vT�{�YpI����P�x]ҕ����$�#nM����]V���hil�	D�(��oIC�v����i�6M��(
W�����p���t��ӷ�Z�F��#���hC��_Ex�x��=�"mw���,�W� �u9�4ݘ<�?>j�����b��f{���٫��S�D���ԧ�&F������+�[�U��D���Y?Cs�]ySrn<�����sʽ�����`��̑���]~-
)������h/iF�7��]<&M�*h:trf�gIg׼��\��?7�/���ۭ^��-�ӭ@�>�1�\!���`�N&��ψY!s��x���r��e�$lU�8���j�jFQ��!�3tu]�[�w�g�[M�!&"�����2��-���~��t���$,Gn�]����|CP�2�=B9�w�}�yN?�J.�C��I�S6�����X9|0gD��׼.le�M�;�M�����P񹝱 U���-)m{øq�X��V��q���	��?���I�Sx�;���s �wܿ�#m�*�ۄ�%����9��/V%�]��ouPf��rNG	�=n��.kW�Խԇ)P,1�Lk��[�[.�+�*�ڇE�X,�Eƪ��5��BS��6�g7��8���c9�1��xRg�����9���Q�Xxp4�J9�CĒ���)��ۡ��퟼���D��@՟E���)٪oJ#�LtDR/sn�&�I�	T׎�ܱ��72{m�%ࣧn����P��l�'\v(���[Z���P�F�9Ki����ؕ�Ϗg�_[%���b:����9�R�2���B�6�㰊gȹ)�5a"�'嘺�&�2�*ո
[�څo<�Ǟ�E���EsoG�v���]��x�ƭ""�ݍ�:0&ZK�0K�
�ո�%@tՃ2�fe��Z��0�g��c�L�����
�N��Oҋ�@8ɶ�]x/>0kS_�Q��h�d]���M�̥���F���qq,�6eʲ<B{�B�MrF�����_R�	yP����wJ��ʁ �w/f�,�u��)�~˂Y�)閪�4�} ݸ۞�Խ����P �s�A������M�DW��%n���6ܴ��{ɣ���ĥ�ޫ��j����.�!��z�������W��Q��y��}�s�?Ƈ���)њ��t����n�w���{�ȃŚ��]��5�瞜�L�&Vk���M��z��A��`��X<<HC�|�EB�e�F�TI��H�K�jx���R�,�e�^���oI�/�`ZnW[����lX���N�n�!As �뵎ub=s�**�9�1�H��-Z�iݵ��i��� �2���w��J��}0e�r`%h��w�۹2�F"��&�fIԚ�Oθ
�N 3���ڕflE��r
�}����˱"���t�/��{�Ձ|Vj�����%D�+�0��$ ���/Ab�Q�O�O��2m��'.��W���u��L��mmo����O���04�U�G���!�X�9�������명��i�k�8�\��L��^�������jmƐ36����v���R��dĒ+�9�K������}��v�8߯$c���5N�KH57��oi��
w^iD�r�V�\�3ݭ��M[�~7Xma�뽏����o^R�~%*�ԁ�A��h�V4�R��"!Z`x'�9�g,>iF} =i��!J����gL5<��e��B[�*7h�W~�E Æ����3�}��7�g�k��'u�;ۺW�	�Iy~�E�.��(C$X�)&8��J���||��#�����^�}P��J"	+�eK:B�~nΒ�^�	u ��X�ٷ�&[_��f�~�m�Ӹ[�1	*�g�iidҀ|�^�Yi��l���$�
�֥S�c��6ޜ���p9l5�J�?rlw+����?w�z݋}�5��:���6B8й�0��G�FF��l��ރB�n�^{���c���(�@��G�ѫ�;�pz�oR�^�|�Sf�z-��YdHg�n�����t�|�������큾Vw�ci��[���[H4�k:�+�C��or�j�_OB������J̺P8�w�����&��o]u�A�?���r���7�%�	-]� �j36�d�n�� �#�XUΟ��`���Njej߳��dĶv�̗/V��)P�5�E����=ݸ��o�ה��z���p{X�P�"�p���x^Љ�+�ŋ\�w�K���V��wޒ�].�)�(��W7J�n3x���xǞCo<�=LBv�9JF"����oNC���|�]�����������R���K``Pi���x���v�V�+c&�8�v$jB�'�̢J�_b�c7�ީw|qo�׺�7�ޠ�Ҵ�WU>�2��m_��I.R#T�̰�](t5`�h�s��#�.��̻]+JC����y��K� ��zd��t�4����mWl��f�B�����
��A����ӌjӻը�f��S���>����8�߀��y
�u����9V	�����qn>�,�[�H+yB�,N�C̱��� ����z�Cs.�*�?K���;�c=�kIjf	�@�o�֘����X���Z*.0q�"W��0�+�k��������� S��!	���~�q)���ԣ�d��P��{�$�pU!�_�R�^��rc�����
s-�����<o�<.�a�D�2<�Ydy��ӛ<AX���YO��o|��(f��M����I�]2�)���,weӞ�#1w��\�?o��Z-�h��2	�O@���3�/g����<X�>xҽڣd�o��bo=эY ��*�gV�핱)[��j��AL��v$�Z��72q�$i���C�e��v0Aa�cʣ�f����o�J9f+k�`�R �ݚU�v�g 	�;;j���/*v��:���F���ټj�Ӗ�<MR�����r�ڻ��7{�]�w������o�M��3����N5[������I��s?$V��5r�9�gJx� &�B�LE��}���*��3wss3f�b���Ͻ$�[�{��b�A�Є9���+W�lCd�gv{e�}�ᙷ�*Z�����e7ý��=�_T���A��>#C���;�Ϥ�O�����J#-*�/ׄU�]����k��v��gi�;=jh���}v���1�hW�^�<=��.TpT4d����A^�B����i�sc}Z{Uy&��i�*��G�щ�Z�7.��Y�=���P�SaT�,�$��^����g-<,�<�&!�Bjk©��;`"�5�z]{p����W�4,u�z�K�lR(b���2�s�T��#-�f��A�K�}���{��K�����y���gfo��3-��^[y������Q�ӯ�x�b�Tm�p��ΙF�d�N��VK��J{NtOtMW�/`��ĝ���;1��-T���H{C��v�"���3@���j�� ʏ�G�X`>^�X��܏]�t-�pV��Ms���3�t�̆V�v򰼕¬���Θ�HaJY���WɐI�ώA��/��f4�XT��c�qu��^0�r�������������ǒuqr:�������p���ǒؓ�PÈ�f����BLX�ڙ�5O]��z�g}��鞋��F%�W�´��4��
eF���$�;�1��;fnc!c���x�ƒk S�u���9M�i�Ϯ.Ŵ]c���xW�'.f+��o;j�\�T�,eˢT9���p��E���(����wYG/oK;���H.��.ц-g�k����Y7JKt��T�ۗ\�V9k��w��'���RZ���;�zy��WF��
�̱[�r.�]����V���]~ιh"�Q�t4ń���՗�����6��f�&����d��?<&V�����$|x�S�ׯk/sڝ��^���#��	�!�t�Ѵ�=$�{J�Qt���Z<�#`�ٸ+��3�j���ְ�y9Y��V�J�G����t� �J��j�����WB��#����rHMp<3Ű��D�\q�Y�a���J;��]�/�{ι�9h3��@i�)\X�t�q<C<��:��W�7Cĺ-X'ǂ�}�о�����_���o|gduy/ö�����t�]h�5.ǉ�w�s��lg�NM���Z^�g֑6��|^V���S+��}��Y=O�og�j���Y�.�Ӕ,�lvv�e�!�5dPKG<txzΏܪ�d�@.�囡�r̺��Q��Eb��1�rl�z��~�fd�9/8I��9Kv�O�u#�&&Y|2Y�.ǅr�_W\xv>����ya24�������Y��u��O�(�|��-L-xAUVC~]�QĹ�j���o	Ą+�b�����#�7��)<Ӱ$H��uv�n�톩$��Y�`���p\�㹏9�/�`��
~��+��t�86@��e#SQE���d��ҫs��M������z�m�J鼾�;��:��e�廪���ÁrC+�bO��_����9v�jӮ=Xo��p/� �5qS�����ß�R���$<��'[G�l��jJ�D������nI���A�*;*�m����2P0��S:ͺH����֯��]8���-��r��OB#Eι�X<^H�̡+�ѭ�J=U�����][.B�$t��nu�R�s?N�|z��`tE9�׳x��{�Ğ�n�F���-����2��x��^�fe�ތ���x ���Y��.�չ-�ڷ���yѸ�鞴ǻ˄�F����ǂ4[�yƎ�N����5�j�6�%�L���0{�t��k*���Q���6)�i�L��3�FvF��W��|Hn׼z�"w�u��:7���eO��Rw��t��j.��Z��������v�4���s�]���j�ߴ*�@*�ULm��L����~�P�:��|���{�Y(g��vl��Ş��ԝ�=��2�|�2y^����=��3�0e��m6���Jύ����uI`�{Ń��L�����k�0TM��^�kj�x%�cu��)&$��,��qx}��n�U�wE��}u��##���INQ랞1Ց�F���T�L�6!��+V�ט �C�¤k�ι�b�	��4US��m���.ԯ.�N�v��Y���߽)��\)���-=�U+ ҵ�W��#zm�YӜ��U�]��[�筜�_%�J�'���O��s��Ի���)��=;`�g�S�B�x=�����m<2�j�3��B.IxV��Mr/n�Jr����34􎮖���=ʛ���nh3)�Ӑ���γѢ�NΒ�]Y����GH������1�\3�+���]A�f��7���ۭ��Rov}�_F�]��C90o4gres|����Ǝɋb�{�����K��X�s���Tf��*�{����vwL@��ß7\�h�s��H��4Ƈ�.�쾎�:�*��3&�sJt��4�(��цV�ӋDOo���Z�(t��uSz�a�d�Gr����e���ԙꋤ�z�#d�ܩ��{����!�( �� ��3����n�Źϙ-��rF.��p��c�0�B���������fX�cZ��%�Z&�>O%���t���ߴ��]�эw��j/ۀ���w��d������,�G���4%�U��D��Ժُ]:�5Ua!�V�t2��l)�R�J�q�����i����F� �B��üH�קD�@؅ִ�v��Λrmn�Lf���R$ TWՊ��P���1,l����)�\i��nv�����d$TE����1Wt�(1��U:�$(T�;;��\���;(Ln̰����F�ȯ�ͺ��9�M�G��m���8�-�+�7�0�!�2�c�p';�[����U�m�Iv�_Q��ۙ˪�!��:�&	OF��p�Z�1C7u3D�I�΂�Ⱦs�]�=���>c:�7hS�}|(���bހ6c�õy4��6N�%l�������K
�!�/��6���y�)k�̺��.d������ޣu�5�|�<��$�+����4gox�7f�Yw�51� #��D���)�*���Nu`B��8�Z&ʋn����}6��y��HR��A��r޲�-<��;Q�6��3��J5��I�U��!ٛ
�\�j��saÛ
K0�2�VN&ȫ�:í:���@��z�bcO/5����;p�����wq�w����wB4`ײ��zucOͿ�y'ye�v�YV/h���\�&�-�lu�6��%�M��
�.R�q�]ѻU��4;E%�+�1�3x�J�y^�^��%W�;������T��o�a�WoL[����h=hm�Ӌi��cf�8�ɭ�V�^�U��<͋� ��0e�c�S���N"��]0��{�Vq�y�ݺ)�c�#Yb�Yp�	������T�v�x���<]��{;H�}-e����q��[���u��,s��\.�Y䊹��u�x�� i�L���� ����w[��z�]+�x�Ṡ��[|dZ��KrP�����l ��R�Dg��������l�2�b�������^ս�v��e:�<Nr��ϰ��`��h>[z��\l��w��MSY3e��I�q�-=�ѝ��3�+ni	��"��hW,h]'-*���Z�&��皂��db\wW.�m^�CA,���uf��Ll�+v�÷.GZOt	ǋ�����ᗛ��h�}���>��}�#s*�@؎q��n�i8|�v��=����s|��å6i��L��duvnb���,dq�[[�Vژy��6�����1z���7���z+̂��^}�����;�7#�Ŗ2~��v4��,���G~��=�QW[��@�?�=���fH��+�,#<���\��Y�߬D3<"���?K��8<��Ҝ��ZfI*^�����ˀ�y�=��M�Xnz�;�[[ة���o�ˬ�P��;�D�햌�����d
�X�\o�.	:�y����y�bc�=�����v��*��z��O�M�� s��Fk#fAr�Id���^����s5|���(,,�h��*��16����9�=Iʣ㶮+�_m�g�K��D��n:��w@o���t�/��:�:��� kz���n��G�J��yᴂ�m���>��,CV)�՟rV]u���:�2��ei�)�[���D3���}��ͷ���!��_|��-΄~&��1�Q�����"R�ks-��7�e�t�3;,�_򷵔*߻tC���W��7r.Ϊ)�u�D�I�k����Yg}��l��V���W�-Ź���K�F�}�R��=}��Ƴz���]�z.1M�z{�ݚTo�h��Ƥn��ۋ_T�ͣRG3EISz��!4ڥ��e����e�U��MS`}���b�}}��wgWU�;Z��XИ�9����F�ox4�i��J�O`Bhvr;�T���p4�>���.f��Xo7�˴ݦT��S��zz����[��$W�.��+���P��읳�;�8Mt<^ԔXE�A��{�==;,:[�D���9e��x|����^��f,<�'ٹ׃Ɯa�wݣ�"|��^�P�y�d��K7�;}3�]��;�}�;�2mY�t�r��ӭz�z�/�{�a[�
�{kz��C���f���H�1��z�[wDs��`�ݞ�/Ƨ�����p���<�QH]�ix	𻏛��/63��m�,��������4w
�u�B�oGd.�ó7��K=en�y�0�D��������Ů�҉)09d#=�=C�[�z�(��K�F��a8z�0�,���dy=C�M��ݖ^����.p���u�-�d��ז3s�G2�7����w^�޳M|#閳4��)}��W�[�t�糧j �ӛ�S���y�R��+��'�ӹ4#[��ף�۲��{��)��Y�*��Α�x;������x��Ϧ�l�q �R�aȏ��
�8�c�챞>�������ͼ�����w�!���s��2�d"�q>��9f��ʴ��+��+*7�[�
 �Y�p��h��ل�ZCԝt<�F�����>��%��m�,Y���=�왫�浸��X:�/�Z��_�=��c��Jf�u|�"�z[{���]��A��G�\�{���.�=]�h�o]�+`)�����3"��]�n��wu�J�,b�Zv������<X����Kuq�#p�{r��4���x���ìwY� es���仮H��f�ax����Tw2F`G3��Z�����'}��б���b��l�	�1aݻH�~�A�]�&�:��'���@r���k�Q�f�ܾ0�����ݗ��M+=�?&}V�W�jD��wl�������fQ���{X'N~�t#g�Th���	^�{|&�f�1t�ʝ�~����O�����b��,;��U�E��G��R�t�_��y���u�y��u�c�9����7�ҙ�ks���t�@��� ��xA4�k,.������40�-��oyz��fa�^ʧ�{ꃭ�S��o�othhۯo��KJ�Vx�а/�\��љyÝlOMl�^��z;�u�(������{Uuu���i�H{սy�n_{���|9��'n��� vV����zw0�\M׀��a���Ƶ�:�L�o���=e���$]�.�LB4�f\��6?T����jU�[R�\3�����i���wP���;W�\̘�	���CQ3����	����ϖ��L��a&�O�>	�/[�Qo|�_v��v.mn�.G�����,g�F���u!YP��������I*��rW/��6����������%$�ݻ��u���wY��x[�$$��ݵZ�T���U-�v�.$����,t�л:��~ܯ�{�
�N O��[�ݧ���{rg��p^���her[.绪���q͛���s/��yh�� d�k/��(<��8;�&���0�u��z��[�s�Xr�=�O=���S��w����K(�}����{��m�;׽Y��+~������8�����;s]{�f.]a��i�8z8�J���.��ko_��9���d�V���U�1J�5{m�������''
�����w^�3�)ڣ��!���=��=:���A&y�sT�W��q �sۘ+��7���Ｓ����<��zn{"��7{aړk�GD���{ʞ�(����C��.e�8/����A��׈g��g���cg>��x���l&q=ƥ��BZM��,�M��^aAٞ�8k�o���v��t'X��:�Ii�F��^󨬒�5�µ-y�}���㵋����WP�M�=���A�l�uu@���d�{�G�vTq<ch���h�13u	Bi�OJ��D|9:{G�D������2��n�!3ӟ��z��o4� ?[VS�ϯ�X�b��jb�:U����ɔT����뇞ڱǔ��ڣ˴O�{����o��<׍_�i�o���&���U���-�7ܹا�ϖ^=��3c�*�o/8�f�&���]{�lU�E���r� �T=<kU�s�1,��6��7^tM�cEzԥ��To.ʙkˠ�?̸�ى���J ��@Cͻ�p��'2�j��=؉�{���~��w��.�N�<P+5��\:�? �_e�v{b�(%Պ&^�Ǡ6i�(���ry���_p��ҁg����:��J������^����O�J�/��ԿZ�ry*�}�񔺔�^�;�,n�L/wZ�z�;v_`�<�B�˫�z������7�J���׹��#a�����o>{���/D^+N2����G���w����)�ɏB�֤�<�k� �B���a=�u��nn0|n�ZO �Y7��zR5��_��E��}��TH�7ڢ�|����t7���v�,���(ǩkǓ,h6g@y4�o��O�,��v;y/d�����Q��{w��y���B�5����9c���fd�i��cat����	W�^V�W���y�=���~�=��ΜiF̥+v�s����;9ͮN�����h{E�6�Ngo���F��� a,���� k_[=� V���� ��T[��בbn�����>{��}��p-�_�؆�V1�ݴ8�T���S�p�:}�=ka���ޫ�>�n�����,�&f=�旽�Йpx-�����Mvd޿�u��9W�5D.<�c��!DX���4W�p�t�k��Mޛj�T(;Y��U����|�{$�.+�	an�C�(�0R���wk�����\ʹ�0B����:̮��n�K5�eM�L��yVg�������g���p-7</8QغCϙ�g�c_�B��Q���f��ŶR���U�Q�D8�7����!-�a{��KɅ���F����mȷ~��٥�{��к�\��ÇG�kކW"��壘���Ǿ���m8:Z����7��S�-��/�٭
k���u4�7��k�R3����U.<��j�ȟ<ݕdP!od�\�y���{+�ߨ����elC(X�z���R���DK����f��v�?h���r���i�uЭ�Q��<ҭR�c�bt�pt\M������C�����A��y�^@�S��6�x��1������4�K�^w�Y��y	�I^A�=�D���n+��M�ȾLq]�l��5�]Ѵ���1l�++r�ړ3��X	}�ZӢt�	Nc���������"�t1��ggDe��;ڛ�����`��[���UnJI��X��z:_T�{\����2����g�a������87�0��>�9��^�9��o����M�Z)8C�y9�����[{^�n-���o�q�����J� a�ޏj���Ԣ���.l�w��[��8��Yߝ�m�
*.�g�F�-�1�g�(��oZ�Kޘ�=+��ܬ�v����<�~��t�U���x�יu��p�lpw�C�f�^nw�lÐN�N�νs_�b������U:��>�ԗq�~��Ɔf�������(��"U�x���*���Z:ҧ�|&,����W��r�����.l#^�f��ޮW�(�Cޘ�M�z�=u��� ���{	\�-i��zE�� �wu�猪�y�2*��G�!��}cYӗ�:gV�7�YX���#1J._Ht�'��,�P��>CuP5���J��z��Ku��v9D�S�c�Ƕ�	�Z�C����?c�/6�Ĝ�8�;�y����m�}D�hZә8�zHJ�o�U�����zXhl������dǼt�`��so\y�]d�0:�A+����nq��z:�Y����AJ�U�x��2I��Z,D����O�Q�A��*�Y� ���yc�I��[�Ĉ´����_KN�V���0"�D{Oۋ~�1������)e#.��r莾!���ALqV����Cq��^ϴ+��6l!�	G�_&���&h<6r��w�]��:p��q��h'=O�\�wz�|���.�y�5t*r5���x�;r�)�.�� ��������w;�'��}�V��p�=�ce��;�(�>���j~��Ruxi��2-��I]�W�V`�j��@�Tv��W� �4�;O���e���;^�r�3�jz�z��b�	�pGk�x�<�R�����r��F]��꼆��7^��5�%J�����:�}�=�v,%}$˷3�^���۬^�z~�mwzaGuC�f������jȲU[~�ab^D*����ey��zu��KQ��%�2�t�v��� ��¶zkkc�2����s&R��ol�s��U�=��pd��VhVp��Ǿ��7!)�1��e�]Dw��K�t�u
�=�M5�w�V���{:�yL�W4�k2a�˓�A֠�V]z�s����,Ŧ��y��U�ݙS͗Ț}�SAz�h/T;Me��+���(�&T��
w�)GyِWu���5:x	�[h�	�F�̬+W_n��0�����8��&��祀5��$�,�h3Y��a�y�eօj����p����j��/�����@d@鎆�����j8/ûS.5M��=cru{a��I�KP�<����o^]B�ݏW�m+j�%F��粟�&Ơ����x�	+���2��=�?z:��/YZO��J�ϐ4L��d��ѳ�;J�u�����z͜�!���Tm���\(X#��D2���LM?%&db�'�uO�F����.=̍n���I�ۮ{�1_�t�MP�dR����f�����̈�,a���:6}
�:�}85�zٕ^rg�m<�xè��̛$ E62�c���s��^se�,�o�,''^�$fЋ�[�/���W��s�����GR��}�Ή��2�����[��/ĳ�/����Ղ�����Iߟ�9^4�+�ST��
^��9-�0�{:���=���ї;���}���=俷��qĽ9�B�J�A�ִ�#�{���+���'�0���+,���A������=X���t�lx弽6,o_��b��M�na�uI�6���[��J���5�/�ܶ���S�͟N�]C�N����r�ƃ��Ԩ5��˭
�l43=p~�	��e���#é�m���=Hҷ�;x�3�� M�ZE��ga��a�u�bl�6�KZ��n�c-���e=�_y{�/-bz����˼��ٻ�y�n�uF�x~�����k���p�����w�u��}�}[�:
UC��t��{c�z��>�OU�]M��):�L�T��rֺ �a��7A`�2����.Y9���׵+l�3-�����}��3S��܎-����J�r_>��uo�5l����Ǖo1����܎���U'�EPp%�ݐ]N��<���<>_xQ�#��;޽��3�V�x�yS���[�j�P�Z�[��=9���å���{r:�3����U[�(ܵo/�QWS����[̹�~�T}�]/7*<������Kܹ���Q��<^9ysб�-"�թ�}��Z��3t}�ru]�FD���E�t������_N�R=��K�]//����]3a/i�B���M������$��uj��<����T����e��[�ޔ߲g�����H��G��������vz�ǯh��R �7~�
ą������&yͬ�jׁ_��+���y�[e���k~���V���Y�|�B�WP��S^A���7m\5�Ԑ��|��Y�/R:e�X��0�՜�|ά� �6�F�&�t/�oW�/�Cn��g�r��'8����#�+p^=BK�*�����q[�|�LCa@�VP�k5e�*��K��+Wr̂c���$k�4�X��o��]5`��8�P�W�dGAV�^��-�3w��F.�3��~��U��u����x9����{�<Y�\��_fѼ�P�(�+f���f�q#�ý�;���Α+���`r��x���?:�%'�1i��.h8����Χ��Pyl����;��8�����'w/��:y��w��s��j$/i�W5Cud�[�N���g-�n�_b=Uϲ��/�����व*�&�^�7��U}G�6z�J��)�@Ȕ���59���Y���7}�8�_V�]/[�y��,��oR��)ԩ�D��WLs�9�^op�Dr�,|��-�È���F���:v%�K T���qC�#f�{�;���Uv��A�G:�c��w�Ր=6�+;A����֫̴��|��=���C�y;�
�̾��ht�N�C�����j۔��X�/D܅:ڕ$�7�q�#���<���\��1P[@ͬ�u��7Gp��HI�:5�N[z���F�0+��3�5�T�(��5�AfZ�/�(�rdn��3ݝQ<�ȧ��s����N���'Y�H�>�8RΡ�K�njsxs�����`��f*έS�-���W���K���VfVj�y|5a��/Z�o��,`w�Z�JX̣pn�P,�:�X��c�^�����qY��h���Ty B�B���7uXգ��]WCrY�R�ם�,��a��|MG�v2��>[}�Ɯ�0,�k8�8�櫤���`*�4Ͷut�Kw���5BRw;{I�a=����\ۥS5B����Z����]��u��/��jI�uz�V���-p�yap�~�W�X����Is�Y��X�h� �ʃV�z�V���Բ�q裴�^Dɍj��j�smX�X��G���ސ��n|y�Fc|hf\�+�6����kBpU�n�e^��=�jwEs�� �c��l��Ww���	������nv�3'6���Z�̂�y�ֲ�,І
��d�V���v<��[*pedr�L�U��`7W��^AJ�?�4Y�$���XTl�nZ�j�l!\�R��\�^�X�:��A�Ff��k;��u�+���W�:}Z�V���ޮ�p�!��,1me�ʉ�Xr�g�r�w\��v,c�C���oA����ˋIMِF21�>������+z��Ṓ�i��;�\H��IP�3Z��q;cJ�����;��}���6C�%�B[��۷;l�.�͈���Y�����iv&�ȡ�yn�\aK�
�u)�1����ؑ��cn����@Ǣ<��Glp=V�������X�sͬ�^n�B8��K{�5�R�ܮ�a�B�L��2��������U_US{�z�*��E������$�n��{)�rJ�]/Y#�*�lT�LSs�!%(��*mdfv��U�����gH{=Ү��5�,���ˉ�z��3��4CIy�-Jx�57>#�����F��r��-f�^M{��KUw�wg.�#l.A׷y&�}<SV�i3;|���
��E{��\���)Y��e��;�%>��l~���v�ρ܁>)�:�%z�%�xC4r�fTg�έV�5�l�b��캄Xś��ΙA´�g�]{�l�� �=`\O�j]��]KV��M1��>����L���*x>�G:h��ᔕyYJ������c���]d��sBX�����^��1A�|��Y0'^��AW~Џp\������i1t=bD����yA�\M�ϥǷJ�b�*�G�p�Z�����9|+�J���^Cz��~�4�[�}�oN�
�nvQg%����[M�FTU�gw6�A�N�(S]`��d����/v��yX��|��q������F<��}8�;�>��������l�d����U�Վt��C�����܁Y���x9l����̡��,��8�I�Y9$z\今�]v����Գ��Ϊ6l�H��3oԩx�[R�$�C�^f��'5|ܐl�끅��Xf����.Mj����h�u�v9�,�G2�|�g_Ӊ�������` ²�n�֞Z��5)�W��;!��%6V*��S9�;k{n���Z,��]���"�C\���FG}7�*�W���4/͒��Y��+ �
�m.�����j ��Ǚ��]��D.ׁ�|���6W��{�nS/�H��7�ƹ��ExYc�5�H�Y�`�l���I�����J��������w=&���xUg���������C�����Fdd�ě���n�n*��z�zJ]��K��Yc��Wr�E��d��v�NKG�=� �7WU�B��� ^n,]��W֟}�.�˫1q���a�~�sS�WJt�%�	�W�мO/��U�m^u�u�ێv[��Xv��V^����n6��ʮ�Y�c�z�+��`��S�؎�`�^(-��@�h�����N{®��̴o��˟`Ot�w�t��S�؇�;o}2�;ht)��+}#S1��º��q+&����4+�7����`CK��\�qF֝=g���N�W�v��Tr�N��y���
����tۢ-{�Iݳi�Ⱝ#Au��tF����,�`A�6�\�"�?/r�okJ�k��a*x��Zg�pe�'�l�x����@�!��G3ms-GGzd�y�.�Y1��Q�6����;[�C� ��v�V�y���ޏyÝHg\�nx�s7^�����V�F5�6J�<�v��zsMb�#���[����έ��>GN�@�m:�"u�@vg i�7�qw��K|t@���k���5�_�2�S�}��š���w%���mA湮;��<����u���#�����I��0���ڽ�y����u�K��_��OlY��V)3ƽ�%/om��M?OT,��Gϰa���{��>��֩�i-�!�c�UhvCf�W�g	g��}���Ǜ���� ����}{^���,�HV�4����VS�5��(>c;!Ǟ�R�"m��R��CfTUΕ��{&i�o��x;��i��H@x"�X����,�ཪ׉H�悴5%&��_.�����#+7v�\ �K�94� ��Cala̹�﮽Dy��@�==���fV�-W�`�ѭ+��9��B�Z��y�;�#�|� ���з~μ�q��Q)��4��y�1��"5�^�y���N��÷I�4�����x�|\�udR��^Q漝/ja��(�� �ۯ�,YK�lf�gj�QE��l���X��2��h���V6���6��:s�E�A=�6��jWX�b3
�$����X�)���x���Lu��QFT�iF��Ȏ�˸9�/�X�e�Ry�������G�ϩ� �Z���o{E�Y؏`����J�[Z�:BX�p�<>���]����
z��`��AKx��Ȧ���{J�<��N��r(�\����Y�7+\�Yɟ�{�F�9˫���V�Tw�����a>�W��ʤ�H�: �hs��VϺ��)޼?tC�̈�Q�E�r�=��9O����w���~7��$���r���]�8rr�����U�%���T������o���9�An�$=%x��DNQ�z��S���~w"��<F��٣̣Wyj��Y���E�uK�δا�osYk}x��y�P��G|v�lVVl�;�M��_w$�L���z��i~�'�;sD��G����]�][�d+�~������"����]�ݏ�G��q�wg�Y��J�8���	����X������fx!Ne�TrOrEq��y��;�n.�՜��N��s҆�Yak�a��0Y���Ǯ�ON�έ[�����䙼���E�aV���f��[Y�=D]+!K���:(&�d�co����ٕ�b��0�֪mu�s'7����L���8����<�usm���u��gp��&�5;�e�6.�v�[�oiX���>�%e�޸y�S��^�b:t��-��uf2��q}��K�w��޵c�����$%{��&��-ܙ+߯ӪqN���,����l�ݲ�l��q��Pq"�ˌs���V���w�������r���క�A��s�Ǜ"��M�f)Z��g2��˥�q����˒J|Oh�5�C��b ]�6�l:����Mm��m=p�կ<��b�9k6}�|��Z5M3po{iުT	�;:��ݞ���sN ���\J�z�"�!�]��#�I�Qh6:mh�z8a<c|�����*�9�)Ey�:���9�[��r��-�n��n��V�w����2T�����������yVf���u�`�,�<a_'Hg�4ի�u	�ix��|��˯p��@��K�f��2EE��x�w�U���Cƌݝ�<�^��ع��Tꎒ��mPb��T�Q��}��'7:'����~1:]�'��%\2ԻNc�O��rIo�b�U|�_���1J�-q����Go�R��lS����m�N�9�Q��j,����rZ�։ur;�Ŝ��l|9��](S�+�Δy�l	�F����Hm���C�Qь>7���b���bh�Af�+	4��JK@�:Mp�t� ØهbG�z�FFv=gO�x�]�Z�[� y�u�betc)��k�mfu�;7�[�-`=��
�{��&v�ض=�a�{�Y�o�i�<��cnlV�L��9OYABT^�L.���E�K��[NDs��Ɩx��g��K�zP˂�ko�돴�G�{u.&V�ԋ7��H��E-˫+D2w�"OI��}�ެ[@�#Yɜ�GѾ}2��i���ҡUW����8��:c��U������P�{�V{f%\�u�2}�-�����eQ^p$xI��Dk�W�nP�vg�S�r���_��9S���|�m��hFC�3A�h�Ӟ�ufE5b ܬ�k��wN�L����s���H���p���ҭj������;�/�}��$^�}%�/��ɥ1ʲ�I�n�6�{��{&;9O���"ڳƟ\��2�b�����C�m<S�b�	Ļy=]͵���O���d�d��"7}�z�:�'8v�E�V
אI�v��+iz�̑=(�n^����w+"�<xe�;V0�&�6�.�����m[M�k�I*�g5#9�d4e�f�;����z�7ӂu�v��xt9����wA�Α1�ʕo�d�yI#�CC&/�Җ��]�oTbh;Sh��1O$���ԂUk8	+����÷tVWJHX��X]̮�����],&�d'�и�,���Ś����Ţ:Ǎ�ܼgh*�����-��u�ʹ����ǜ�Ñ����ߤ�it�\����o�EJ���~pV��giFM�"����}P�'W��םv�G��0{ciJ����BU�}�0�U�v#����7x{�E�x_bͮ�p��!��#���Mފ+<�y�/a�c�3��=c,p z��G�{T�R�S�	.���g�ucw�d�}�MsJ��RqW�ߚAz�~��w�S�^������9؈U���P�/�M[̧����]��ϒ��lvs� �7�������#��b�G�{=ׇ5�"v�ܦԀG���F������r�3�S/����A�b��1�3�+��
襹w��md��=+��]u.��Y��;R��J������W�0K��LYt�n^��C�=�8��qΫ�)w=e�����g}-�Ow��m�܉ڒ�ʸWr��/hc����X���N�8n^:pF�_m������ϱLW���9���\���ۮC�ٵ�B�X���÷�4��t�MzԵ�:�ꕳ@oK�����b��K3��Ji���]��T���b���Ǜ�;&#��;��
q̝*@���5&|8|�����7M�(��CUu�0+�K�N̍��Gԓ�QsF�G�ۣ��?u���n���s&����p���iϲ��E��k����{ػ{�3�^U���NG�,:��
K�䱯8��+(��ٍ�^g�\�t7s|�V7�����G�;��O �y����n�Q����	��dz=�ʴ�&e_��uRD��CHC�ۧ;T^f�T���{�Ҝ^Qqa^��Q1΃K�\!�C%��7fo��ze_�ϞN��S�]�6�@����(d��=�q7
� ��r7��۹[�w�+�ρ�_�$~�p�BO
]��07D"�����t*�8�z*�uM:��`��e������eiM�rA���ՆH��'zsʼyK^�7o�sP+�XQ�&�ݔ����LܪK@�}7�Jα=������ҖK����n��v�W���˵��Y�{n�<��ppt=wt�->==�+�Jy�&3�`ɐO�k��m����Ջj�f�6�j���o����$��T���fXݒ�p�jo7Z��r z�N�kR�7�E��M<��v���u������
A9�=�Nz�w,�W�Q�-��?lG]��x��Zᛳf���ս�	�UL�o]�mp�:�f�Dz����Է��O���KY;A�ךq�
*��!6���ǫN���=���n�ɦ�ve���~���r1o��WY~l����l;���lY��J��nU�~�s�l�(0�է� �-��!��N��m�/E�Y̰N�N��l֒}	Itxq�����J�4p�P��&�l	���q�5�{�M!�~)�i�=C�v�: �2��L���y��I�+�C�s�ϒ���W8��m�߹b�5�}�bv�19�_M}�³n�Uo� +<�< ճ�b��W�҄�=�{.~ҧ<�Y����iJ��k/s�[�v����?-��x����^z�܃w޽؃�;������W¸����nv���1`�>�s�ر��-��~5v�yE[4
�_�c��5)�׾}E��P{����f�C/A�[D�&��z�s�W��u�����u�oOec�{/Fy)��Z5����d�m(�;wI���������A�:��ø�N��Bs��β4��,&��__ fM|�G�!ѭ=��b}�]v�2ړ��f����ۻ�0�� ܛ|[ �P���fRW�F�]=�����-⣗������󹒉�}C�-������p��=>����јJ�]fMSG���Kw&=w�1�QoZ��yw5]y'n����1q#.2�y��o@/�m������J>,��d�`�·&ϫ�G��R��㷡YЅ�t�r�|Pr�$ݝ�0��s	��i��g�L�V������{rwn	�㲸�mI���D�@���Q>��rv�]��/:�~y֏����R���Џ]��s���i��=瞤����h~��j�d���=�!�ު)��a|�mŜ�ן1��u�wk����קn��_��
,�|�����y�%]5/��s�!�ڡ9��4-6��߰t�n`�'���f�R�W�mRQ��t�O��c�۪.eOk��D*��;��/�=ۙ�a�{yFߣ�1�$�%=�-���~��S��^%A��櫀;^�z��t�s�75Y{<���[{SǱM䨚��S���=������t��y�'���#KZ`?)�YL�y�鹾����(,����c�ٔ�Q��Y}�ΩG5��[��^���i��Ei�_]7�OW���t���Q�_��U0b��Hq���e{��L+�]�K�@�oF������[6�	����흈�L�+\^qY�`W�g�-���aܖ���Hr�Bٸ�X����m��
���lT���OZл\�ݬ�Q���!ݙ4����h�;���0�7���*���{r*���]�ٛ֠*�rR�Dvj�1���ۊ^���ZE��"���L�?G:T�-�i�R�ބp�Iߵ�S��J]���#V�xvWT���ǡ��r;&l��-B�p*d��V*a��l��M7��p/Fi�n)u�w��Dj������}8fn�I��v����	4yQ����W��D���ʜsY����n��懹>�=[�#�Fҫ+�6,��=܌޴5j���2luX�|C��r=H��ԧ�.�ºw- �v���3�k8�*����/�o��J�%j*�#�+[�S!Ħˮ\{FWf�Ƚe.�}�g�Ɩc�8�7���N���_���WG~�}�&^�m*�_e��اb`:�;�fJ3��g�Y�ę.+r���j:�t�}��r	��1��e�i���k������yr�'Gkj+-�f����e���
ZƎsoP��S�A9Z"]l��qV�ӘM�ek���{�5pS�d�(h�30Qs*��d��홝�����us���T]w,�c��
�^��ԕ�3�k֯/Z�|�VTѯ[b-�Z-A�r#V���]�����tI��=�U��X������Kwy�ޣ�;��u�8�ݎ�7uj�]�Εuk�r>��(283%� C�޹O���f5�!1����R�N�ٽ]̼�G>|��r�"S���24�w�y�1D��mv��2ŏ��� E�:*�f����
9����6��T�X��Gi2����*�<�^ݘ��ޛG,
�L[�:�p�xּ�B��X��7�A��b�j#��]\oR�v�O�������q���R*��}�L+8��˜���9m�"�A�-�Q�ثo�=����ޔ)V�3f���k"Oz�n����"=HV)oK�Gqft���'0���<��t3T}�(�;~�N��2jp;�j@�X�E���qo9�4o�5��tʒ��7Z�:���"5³U�d�K�ݩh�<��E�J�E�P{�z��6��c�hչD�u�̝G3����3���v���?v��5�I[EN�ӣ��c�'[I��j/-'��0�
�YCVwq�X��u���=�7���񨝫�к!Qzr�8٫��+�[���8�tq�Jľ�ou����z���7M�w:�����u.pq���Kq=��-���4�����Z�b�[���=�m�m��P�z��Q�X��xljR(�S��V�����Po�Q�b4�1p���қ5=�9Z����x�^umHa�C`�T#!��@��wP\�{XY�޺|s9.�#A��;H?� ���G%�����>  +	�O�G��ߜk3�ȱ��L����UxLCj��j,c��PQ�Ui�l:�O06��ǚ�K��w\th��.�j��'uС��:�q��j�{�J�V��g�N#��Mܟl�>��`�0�<#�w���k��-\��
�W�X^��&z�Ye:��V��ۗ����v֓��MFG�vyD�D����x���|,.�c�ߠ�ǛE:Ra˜Ss���w���f�3���z揀7�n�U��܃�~"�"!)�ٻ�v�U�.f��(,�BI<�T�Ǟ��䮧�����|Nl��Ή����3��j����Y�G*b�|���w�P}�Z<��6Aj�
t�u�xdN�]��Zs�|d�q��v̼չ����ٷRg��n�(�m=�'���EU��!m�u0��n3����x��5��'`��C��K/zp��F�;����
�[o��{˪��m�s��6�5�J ��>��h�P��e��n�̒��ac��zk��l�t�Lo:�I��b0.������q����������L�y�P�ai�B� �g�����������<�(��Tg|Ƕ�g)B��	��=��.6֝܈|����V��U���A��� S��kv\��+����⋏'3�����y�[_{
 ��7nIA�q|�J����g\�+�,M�c�_]㥓t�� �IJ̃F��kS��r�؇�S8�·fVܡ��RC��u5��W�gmh؅��[X÷�<��
װ!j�������[�����C)������v�|���s��B	2�K�����Lw��c�R+"�tpV5�)��l��GPQ�7D�F[7P@ݢI�윯Kϰ��VZj�B�S��쨲���O|�<5�m�E�M+W=٠��e&F��k���î�*El�e���?����3�B����&��+ZUi���O�%�e����K݃[X�G��w$v�S�#.[�	��M8Fd�j�g�|��)�h��ݵ�t63,K�n�J>
R����\�[����ǅM�!º�`b~�7V�`��?W+So�4p[2Y��WCQ,;f��FuG��/��<&�w��ڧ�3}|#�=U�!��]�A��Oǎʋ�54��כ�V2}�N`�Y"�ȫ2O:#��UPs�nU(��ⷢ�b���YB�&�7���'/=������>�yb��|�KY�����c[���C����UF����'/���صՂoӱ�$�saݫ˷s���Q��X�t�W�:ʝ��JX�U�t_�tN)��&=�^���Ϲ�����;鋹W�Pޤ<S:�v@���4���bdE���Q剑ˢ>�CUm=R*:{r�DfgBC�ԋ��9��؝*�z�hj<�js�KX������`�hM,mq�'�$oC��-4�,��.�='68�[n=��*��w��ݴA�È��=���z�e�r���.�Z�������5h�K!��`�uW�I����8�ڳ\t�>�o��8����|��i�{���=���lU�鄢��Ss4�x�ac��[Ў�/Z�[�J�G'U&5D��h�t5�y&w�P}����K�^%=ŝ���q�(u�\I툝jn&N��{�Ynq`�H9G��q�#�Ls�|9F���zwR̈*���0�/=����}�X6xj�T(��O�NyQ�b���=�������׌���Xr�n��W8J�~���
���%��d��.G�⟥��;�[��X��zs;,/9����s�'s'vkN�ʺ~)�,�Uf�㾕���f��s��ֶ�#�kb->2p�����<��+�^�g��a(�]��q�׳̦.��O�cA�K��g���h�`jӰ�^���+w뮃Mi�/C����L=9��$�P�s�yx��;��zj�{�i��.G�΀Ђ�8�]���wT"�>�{�ў;�=G$ʈ�^aJ�pE���hnU���o��h��Ǵ�D�QP὾�A�}�3�u�~I�>����5�]wV~[��o��P��>�2C{�xÕ���_�MW<xD��3��u�#����_��tLV���A�(�C�lo��ʒs�<34Y�ϻ+c��L�aaU��<P�c1�:��6+����&���wH480�/����J*8�������4;}ո9.�K����h���^w<\���c�\���Bų�+�X�':"�Q����@r�;Z�[�ٴ�H�8u`t*����(���IU�w�\���p��TY�${�>�)"NN�"���5�<J�m���ʨ�Z����	��	ڻ�2�Qʎ�+�>�z� �eq�s��r`�\�1���7Q��S�eP/�Q��${����{{ob��nOM�엥v�����G̭���/;k���Є�ltQ�~/ګI�x>���O OSħ^z�3���|�>�6p�tFle��l���u�#g6v��o��*�;Ȫ"��p��6F��-~Sq57��9}1��ݙ-i���+����`Y菈�ٔ�q�_�Mp��z�R���W��=�b�r ���N�x�GD����v��DgL���\A:���:i��<j�����6m���ͧ��g߄��_�N��؊��\�f�Oplz!�Pa�o9���ES�}��,YX��x��K�Ź�`�.����뜻�9fغ� 5���,zK�=��*`w)j�N��Vi��o��=�7r��x&)
������rF�j�ެ����O�T���C�T�*b��U�U�z���3�0�Q==�u��]p�B��<�=1�Gau�f�=�w)��{�h�Ș��i���һU���NO96|��߭H���=+ʹ:P�9��n�-�ݻ�~%8��?|�9���8���g^p��#�n8��I����F^�h�>X ��f�ǭ�pd����f��I�}�EE#�'9Ϯ<�����Gt��TN�ؕ�"�i��UsY[�05���u�T�u��Ul���n,��3�NPt-.����I�j�J�n����t��$H=j��q�Խ��:;�M�㣮o���yY��(w�!�[�	�Ϸ�ܓ�ɹ����̌��7�)�xZ��g�я�5��A��N�eX����䪠��w�y�>���wƢ4��&@���ґ]~<}�6�*�̘>ROO���wt.�I�]b��n<�|�;"��Я��J����+��u�T���-����q5�N���PM�~щv�*��Gޚ$:}̶.������//B��x�G�<�z��!�oH=7�#�l/AD��
��}Jk����U�{����37�J�%��`n8�-�Dy<���#y�@���g��T���@���{�V�׫l�q�{S��e��s5�.ƍ�����XI�e��eg�/ޣb�F�˨�=h���QJ��(>��O����K�|��5}Z�}��܏?`�qJ}3���6�g� n�W�U��{�j9`��7��{���[7R�\Z����t���q������c���cfqz�'y違� �k�z�ʟH�g���OznE��x\���8�_D߼���-�1*�Xc�����rײ�'s/�Ov���N��I��wX�v���1��Y�7"?I`ŕ1�^Ժ�R:�Sh�s�Q˷�ڢX�GEn�Mm�$�+�'��K�i�: ���n!q,� ��u��n�N�/%�tz_n�݆Y\����.{M��r�������:M�j\�һkO_e���L*�y�"}xM]���?Fod"gbj�G�7'��=�<�8�dj�لϺ�VEn�m��5k)��Wv,��UwOjS0�ñ:�*��S��NLۃ��������^����Ohh}��"��.��>��OJ�������?{|'wbZ�UllD��]+6.�#�����3�+�Z �M��;6�q��Nf�ۋ3���n��؝�����o2,`���鈒ܽ�#;6�����l��{`v��\���;���l_`qzѾ�9�{��w�s������3�OFt����E�\_���\ǲ�����t��Y�9��[[�2�
1�7�P�ؼ�y�w�c��Z�ͻ���]Yxx�.Gb6@�g{O�1n�ꪺ� 0k%���^d]T{��
�Up��Я��Iͨ�B�%Iy��1̖ �e�٦ϗ-��v\%B�3�����$�}�]+e�/�z�mt��*�\�ʽ��rW[�g�3k�W��l؊[�r��� |K� �펿;s��Cir�ӈ�Y*<a��fe"]UyK��A9s9�l��N�)X쭠�L���1}���N�޹�)���X����2��!�lj�Eo'�{A�wf���=I"n��S��l+4S��-֮96��N!����#�uҤL��Rs��u�8���Pfnh�����kK�-�ڴ�۬8.�"% � �N��A��,v�����g�Z4 ��z-�s�鈙�:��Y�~�t"r
�W�w��=�Jr�q]N��e�[6c�㓡vO{�t�d����\518�坃+ƣb�ǳ�V�o��k���l�<k ���҂��8������큁������L���h�y�h��ɶ�;��V�p����ƟLԌ��7��_@ו]��/��}�\_�˴�{ԇ���wby<����+���_���z��W'�(=+��0m�jg]k���@1�~n�K>�ˈ�p�\%Z��h��\��5�l��i��V>������/*D���W�Z< �	~�k�t���o���$���Fw�gMNܹ@��VkK��Yh?]���o؅O������n� ��W�|�����]K���Ի��i�9�H�!����㶷�9q�`s�w)��!��T���̌�g�I�QJ�e����0�?K�`�ړ'����X����dN�m5�f��u��؈f��"��|n�o�}�E�a��K)f����Ԫ��������5�bC�tA�C����^
��F��JYu�Q׿�e�ʖ˅�щ��Am��N��V�sO.��ԡݳ�1VE\+����"��8��gsb�F�QC>b�՗]���.��wPs���9���e�A��R�V������u��r�n�x1-��2S �ݝB�<��L��f����B�Y�.*;ەћk�������w#�}>�'��sp_�4������������j��⟋Y�<��{(G�c<�]/wlf5���(�YO<��t���}'���.ŝ�>3�jxV��$@k��G<�i] �x+<�i���b�U����`��7j�Z�B���2�C�ř�Q'	����^V�s}j�L��,l�/d�2�B�B�T��K������V���OK�د;�	3�Ć��8J�����犎<��~�Y�KU0�+\1��[OW��	��F�:��N'���A���}�g.��'�Y�@������2��7�%""�w4~zu��T{d���L�*"�0e* s#e508C~��1�73��{X��������:���Nʦ��]|u�5��qN뙱 ��Q��<�;�0�߸rJ�}�)`������w;�F�Sl�>�֕�s�gݎ�%Ԯ�į_]h����s�΃��)&��pV�������vkϬy���������Q-Z�s���tl�����2�,5G�r{�Ю���9/�z`�mx���k}�R�d��U�,Y��(Z=1�T�W�����D����Ҵ0_�h`Ȍ��ÝyLp��ќ�]�oQ�-�9%�.���l�+E�3�1�[f��μ<����R3��X+-S��\�*�+�t��ւ0�4@;H��>4�Ǩc�̭i��9r�� +b�:��Z�*�9����	d��WX�i]C��:�L��t.��Ez܊�c.i��I
��[Js
nnj)E��8)�A�m�����Ss�4�Ņd} 3��b��x�Cv�j��N�� 9�{��9u�2���gf{)9�"��sip�c�{Ƭ����h�o��y�~��(9Mo��n�v� !�/2/g����s�M�W�i�w݃ޫ����y�np��:r����r��]�V����s/}�֬ǁ����[����-�ˣW;��q�9�sZ2���82���?Lf}S^R<��������/��S�v���2x���!ƫ��(X^�g�^n*���ҮG![���¯r[�ߕ)aB�]�N�'�� w�㟺?4�=�;c�Y�ޅMxz\v�@�ͼۺ�}���T�Qg��v�vf��.r�z���9$J%tGï��ۚS�7�h���X='����~y�LQ�ȉ֋>/��Y�u�N�Ev�"�nS_@�Y������h+9P��8]�\�����]�K���"�NH�E�{��BS�˔�Y=�Vb�.,�B�'�g����0�������~�M�˥�����^�$p���Uw�ɷF�\u`��D�v���y��k"t�yQ_h���+_Ǹ���K���[�)ϒq�ppȶ �],Y��l꺜�.t����K�J��{��j��<5*��ʊ���s��g��ỽ�/���ɏ��T�L�ۗ/��] �X����Ү��2V�g�"�H���k�sJ⦭ק�_UvT�siʣ@��Ui��1��=�;+��ns����k�����a�^J;��%�Q�����َq�z2��4Nc�i�Ƭ�LJ<v:�j���]�\z�Y���<J;<�d(���H#�OZmm�+1�x/Ѡ}�(���>�:n~;�?��:������ۗ}R{u��z���u����qXt�.���B+F���#f�
ͽx�N���Bn4�d�؎��t�Ss[��Y�=Z��]{��J���oЇ���(ʃk�]���xo�ek�h����3�[_���;�n��S];���wןU�5�|��v�����z��{3ײ�w���0n��G���?D�U�p��VO�
�)����n�l����^Dʋ۬�Y�����ۿ��;E�M8h��ͭ�8���cZgT��܆��y�^ij��kY�=�̥0e�^#�ސ샷�+Lz�SnZ(�%\$�ڬ4G^>yS�����ЬG���״�)H���l/�Z'yiP߯+m���k��ÛL,D�otw����[���k�VU��4�8�tl����2X߻E�x������vѫ��YEn��곚�@qbV(5�h�.���m�h�3XY��0\ㆱ�T��w���α�+������넉˺�Fm��D�H/>#��ͦs.Q��}F�͡���W��&��}Uo�ڕ��}�S�qJj1�k5�d`��EC�p]�c#R�jͫ_|���6���
�b��`y��+'h�֪��o�	+��K�<]�P�m?�����UU<�XR�>�|�ۤ'�^za�{�Ry�u�{�3�����T�+�'wLB���YB�֫�����#X�G�N6�m�ˌ�{7e�ln�h�뺙x�&������<�s�ʈ���~�$�H��`7����{�=S�W�%}�U�_W��a�3��W�T4xtˮӾiߏ�/;��a۫�On�1*�n���"�#H�pU�-m�\���7�N*���ko9x�n��z�@r�!���<�f!�bKe�U���u{ފ�+�C���WD"dU�>��+>~�Z�㰴!�\:�)DY<Jc�o�~�i�ū\�ӈ�����
%�+���]��w�q��9��H�0!-�Xѽ���x�is�zf��g�}��d 4^�[-��Q��-W:`�3Gtv�}�B�H�0a�(� r�U�PNm���yׇ�K�3U�Z�\��Cr�9�f;���6]5�\�d�����!����I�HS����&do�|���R���yt�r;�7�a����H}�X/,�X�ujNڂp�e����Q�8g�s��2�ᄵ.�����K\ʧq'�(��-Z�r�ͻ�*~ )u����*��J�v��kR�/ew8�A9�nn�B�-�p���DX��'o]>a��T�.���y�Y}��S�۩ү���1���/���U���V����+���d[�T!#�(�ژ�}a��Z)rxHt��c�O9�c1X�q��O��PfB8uKq#��k�m�ҭë [S�49a:�!+g2I]���*�g
Ud��)�ܔ� 
��~T+�����_�@��]�<ھ��݊�u���G���9��u���������с�U�R��R����=�"����)��7v��Q�Ȋ9F��m�o�Yj�s\�.D�On�}�+�� �+ȫ��=�����߂~���	�U�g=n��v�)�g[�����[�t��*7s*�Vѕ3XۻP[<y"2v1v�3��%�Д9�����}�!p�x�Ҏ��mf�|x	m�י�*Rt�mG֖���|af��q���W6�D� �y�^q�9X�Z(H΢�B=�����X����;[���w:tzi��}Q�1�]�{1��n���EU־t5��5)t v`��+pV:�
��+��S	�Wv���eĴ��`�u��@�
����d'��](*o�խ(P{ȍkcǷbjv1��I���ݧk[�f���!w
�o���=�fڜwM[��r�J�af��I���9���݁:��&�VS�3&�C�P���keMu�K,��;�x"6����-��%�Q���1�^z0�����q��ST��_���ʼQ:_���5�H-�w��䓭�m��CW��m��u��®�,��N�41k/�l�S4S��K=����{z�����m�ߏ�a�Ae*�����k7:�Iӷ�i�:2c�2��̉�\�P�̕�)�I�ױ�^��$|3`�����;�μ��S��C�\� ��Ln�3o%�#�S�ڼ���W��Ϧ��/o�YE����z

�$=Z��׏��4�~}*b�4ќ.�3Һ�Ϲ����g78��\�/n�D�=��:��Et_~�<1��)���}^p��z�Y���b��'��քb���!�/��6��Y�򞭂|��T�>��۸�>��]�mٮa��n�˭�Kw�F�u�.������m���_W�.8�WDx%�H���/-pK�_
^��iE3�4�'�u�p�R�^�3+�Yb�����m
��˻�&�qA�G_���<������z�P�/�ˎ����S����S����$7�czVw=����S��ι���Ց��a+����2���Y{��}Y|מ�c}@���Y$R�{�>�=�cN��s��s���d5~�l��O�V�E�ҧs�_�!�C4_�{�nK�|)�o�UU<�*B�g���0�������_�Fj��S왉��QdM�����V�c�ju� T��颃�q�Y[]M��&��R����\0S�C����QC�׹����3�ND��-g��j?P�kUL �y��_&��E���ߌҩ�YQ�Iwv��v��k��~�0��#yˡ�~}��z7�"�zk+*&\6�
1�!V}}�I���7�y��F��:�T;_��]������0.]\��JØQ;1�g}`����#�/W���=���&�,r�C���ɯ'%d� _���K����7
�w\]6����2�"9t�����|��Z,hYv��֡s]���I��M��9.$-��E�+�`-q��K�n��7�G���7Z'��<��F���WP��byAO_"T���fk�}_g�/�����S�o@�����x	�yv����w��r��mt_mL�������5�aa��5.7�{������f`RryD���|L�0��(v��V�=>p1B�7�ռ����^��.8,��p��忲��:�#�8^����}�+-(;$Efw�+WZ�7Xж��TZ�#f��������Ew��9��3�]��j��
��og�+�鼁喊�y�'z���f�Qs��>Mw�:��q@���#���0p��n�ς���>K�}[yc3%H(���"�7>=�3�G0X]e*(�<�Elx��g���:�N�x�ʽ~�a��dz}�ϳ(*)]��W�mt:�̡���ٸ�Pv�p���� �Ϙ�>����{W9��V�v7�'(������P���N���x�)'�7��GC�?�Y������rt����|�«jQv����s3�Kh�����2���Q�tQ��~�޷�.�S�^���Y���Ww˻�FW;�����}���]� �ݜ��n~U!q�q3d�J����	Y9�"Vka:�;�,�z���}{�'��H6��wN[S��^��y��V8������[�:��E���JY:�У;6P�\7&��Xj���:)�E9��Fo�mT�z�ٝ/	�/t�φ{�L	X�jj��x<M=��/a�8/<#��h=17�ƽ3���V�7Ǭ����*ړ;#!A�UT�W0__�ẩn����5]��l'�{�{�zG{0R�1J���F�ꕉR��D��3��c�>�ô��0�X�Sj��w��B9�EA(��_;��N7Qy����S{v�2�(7��D{�iuǄ���g�Z⺪K:�o�h�F2(�{���Ga�GT������ڙ�í�I��="36ǈ�n_�j�s+�z �L��5L�Ea?��fdz�f�4D�1�ʚ��d�M�:��p����]eA_�SK�Fs�1,o�̒�����aϓ���ܪ�Y
,%�O�;��4
�t���;�Ao�3ڽ}�Ej;3U�`im��ά�����1����Py���s��}�5���\樀�O�Θ�۠	eW3���͵8�g��G��u���ݡ����m
YiWC�V��ᆛ8.��y-�a�}[��i�2ՙQNMm�a�ܣwy���jB:15��]C3.�t��W�BF�;}�?f��h��{i�o��:��x�,��G(e�vF��L��j�ug1~�n=�Me���̗Q$���n�.�dr~��#5:�1��#���Ӌ���G�'�'c�~���"&����������=�಼�S�ʞ��^�>[�ïb1{yw!>���b1䩬��7�̭�q�C���B�g����G�<���G�<4<��w�j3�В+<E<�[�Cm�l��s
ȗT\b~[X�NT��bC5�UOk�)�e��Zۋꚜ�BhIt"��o��/e�]�`��T��f���\�o9c�����J����L���٭�֐���z�k�����}�<9|g���"1�iѱs1U>�[в����S��N0@�NM��1�����=��N�>׼ܴ��Q�w(Q����Y'�S�߉�E:2㐪��������c���xyZ���1�����=I�]Q�}�{"�K~����u7�b�9d���%�I[~S����6�Xws,4���!�����n����\zx8��2|����J���\���H�yѽ�&��ئ��w`�8=q�hͣ�f�,+ ktX�I�b�˭��y���K�L���b+��v��.����� 圈���7��,�Ht&/�mc#=*8�G�wgϺr�vu�=C}�v�o�d�#D�L����~͙�8��Ӊ�����.@?����N��G+w��_�����K�O+�7BO��Y��݈�Y�DS��;Qy�'������0�/r���
5z)��S��F���u�|ϣ6�}�מû;�?��Qn���Nϸ�#�,!5j~[GqΝ�R�LV �ƪ
u�)����u�S��T��棣1���J�r�಄�{E�X��M]�,τN�yT�4{���2�9�>��<���hV����׈�c}6�tU��#�ɛ�o1ܵq�ȹ[:�� � ��Xd��g���W�z�������5�L=��gC�*!�=�ȝ�Q]$���?s�;��>Ƣ�G�Q�����i���</Eѹ����^IÆ�i������=ؿl+aІ5;'{n��(��h˘#�:��)�*�9���1�߭om�O�!R����k]/:��t�Z�uIA�-�a�)$��i�<�-��F�jˡ��ww�3���h�S��ïUƿg�5�\;%�>(/W�D<~�J��$�9�oJ����\�۾7�JG�|�����R!�E{9P�\;��I��j��AP��e�� �J� w0�$��3k�lQ�P�ClE�|��t4��N��R�]�U%:�$��b5w�����ѡ�iܗ
�᭦�NO�N4r��]��R]��HIjuH{�{����7қ��Yi��RfUx�/ŗ`Ӱ�?�����s�w�'׵�F�@7f�*��\�d6fv��hـ_���&o"�6OY��p���A~u���](�9"c5m����9�W�4ʹ�"o܊������P��X�~��r^�{��z��T�����1���د�7������?]�*0�}��~��8��<i3.�v'M��Q�-�[Q}���oHp���3~���D>`o�mb�A�o�C��3^i:��n%-�o&xNPP��,�Bx�6[y/C0	4�wsn_Z%p"��W�Q�>s/=Z4�r̦-$W���k�x{<�f����;��ozֿJ^����@7��I��,�Jz(Us�Y�Ųƥ�[,�:k���ڮ�>�QqXk��� ��2�٪	��A=.(��/�[t\C�W+Iw�[u���۸�D�f��K�ۗ�g�"�wn��K�=�Jٲ��yw��ܡ7X��z�.��䢢W����c%���iMT��ܱ���b${/%sl8���g[jOB]���:]��'sw�t��-��;u�]+�\��kw+B$P�4o����S���o�=rd�9�m�T1��fn3�V���;f�գu�R����R���\w�g)�/n�)�7L���O�z��b�&M�/$Ï�a�]@vOr�tmς�PI����m�	��b���	��u��Q��Y���������Q1�<2* :L���8��n�	+k���W��X�z��m[�p��wW�5q7��.yq>6�f*�#"���V.��k��sF�xS�-����	�:�:��~�F�܌��
�v�e�*�h�Ɉn���(x��I�<��h������u�{����y9>��CqXA�Rq!���c[��\Y��n���xj���:��8��������i�D���lf���G�LbS�N��0����w�O����d0���:l��a.U��t��O4�����Z]l[���gֶ.j��֟�����s��;���ŉ5��V���Z���EBWO��c�e<m��F�ūe�mV��y}��K��$�s�~[�A�{c2j\�[����Dt�xj�%����xRA�wp�]���VF{y?]�?d��j�s�S��o����)�ȿ~�ڲ���o��,�2(�U�z\Ƕ�����,�"^�?���x��{۔;ִ�	EQAL�� ��'��/Ά-�?b�~����e����������x]��+w5��w��[7� ��oyL�O|4e[Ed���oZ�WPm���!�U3��p%·����K��t-3`_~1+W��M�x"��wq|ե�ج�:pƥ-��u6N���W����W+~a�ˢ�z��;#M9%���݈��B�d��sTr?-�\S$��� ��jycit���}�L���5S��ͼw,[�u�Kyr��m�[��ߠB5#��>�����`�uV�:X}�f3f�����/��	�!ٝ�ݮ�]h�]�o^�oMv��n�WJ��Dy%y[��tg�J�V��S=뜛5Xf�x��ޯ1�^���ٍ������9��8��/����8���W~�4g�ޕ�XU،�Ɖ���͹c-��|��L��RD*�+�o�j�Y����J��k���׬�w�E��K�l^9�İ�f�R.�wt�*���|%	�[Q�&��W��[c%�����왾[<l���N�\�Y�����Cݙ�)Knֈ��q�p	�$)�.��SC��6���J��^�DGǖ%��uJ�+�[�M�T�����p+�{n��}�9��h��\�G�Wq�Y=�� 1��)��6�f9����N{kE�ʦ����α�z�����EK��J�2;�r�2J��9�Z�I��{��H�L
���0��G���� �c���J�x��[����+-��:i���P�)��� !�`p�iNut�#N�.R��;�ʹ�	�o^��wv�ͽ@r�Dj�{f~�0�-K��uP���xej�}ȼ��[�5�����]C�́�[��Tx�{{�{����Y�H̓ׄ�J^��t�n:��qN���]����x����S��7.�c�w6��n3uF��b*vS:�G�W[�a��<bh��}�]��Յ��e���+��^���}_LY;b{S���{WM�(Wf{×_1��O��Cx��}ưs�5���T������͞�x�X����y��D,�wِG���׶���t9������ѯ�K/}�Kk���d��b�l7�9Y+��zY���6���{+?n�ٺ�����l�}�B7��u���|Q���&v[�j�����Rv�����l���\<I%�F��^Ǽ�Ԣљ�S��\�\�lm���2&5�E��4n����j��l���m��(t��7&7%��1��37_���aV�U�i��u�����
��gE|�=�.Ǐ,����2��_o}�iߍZ��lt\��Ҕ������ff��o�F:5�tq�w"Z�͇���|f�|�F o^m�j+�6;*�\�b�V�#���Vv	�C�L'G�PK�nn	���]	����f�^_�υ��&:<�c�+\����u{��R�.GzP�bU#P�R<��-ܽ�
N����(�p칃.����bU�U�=�M��c�A�k���w��A�*vd�����B9C�έ/m�l̦9Է�5���,�R��XnqU*�+�^��,wj��\O&7��)[� '�GH�{��![y�n�(��tX�Ԃ	�{`]�k��w��:�����ݩ�A�&�ֳ6 sO�6	�^.X���JoP\��<j�ݹ��9z����Xș6�ڣ%젬DR%�u�63[g��ӵ>yzؼ�b�O�;b���Ae6�NCGE=�jM�!\r�%���ty�oGA�=

��j*��U��z�o���'��Hz�U�_�~�jJ]����w��~_uFz>�~ހ��C��o������D-�M#��H0N	�"��������7
�U��o��y:��3�j�vuT�R=�4W�ȋݗ�:^Wm��Y�{Q-�܇�����E�Tc/�T�^��f����^)^w�V����=�m`��c��{`�~��}�}_+�5l�s��}s�GM~%��?�ƅ�y�r��Iw���R̹��?��ZQ�/>�ﶍ�uv�2zV��rj�K��.���n{5U�j�����(��1�+Ut
�Q�����u�緼`�8�یـ�;���\��a�+c�]-\6����="A�/�����?6^zd�I��F{:�����4����h�ع����U�ں�#̛�C/Y�[�lc^�_�>5X��K���q�jY3f<���9,�D1J��P��d�ʞ�b��̴�M錔>rdv��U��*J��Q�ռ��3���j�CW�}��*��Nm�Z���L�R�h�����@rv魷U��E��͸�RӜʰ��IX�&�b�(_�����L�v�]R�_��t�.�꯫���.Q�#��2�YQ��˭����ܾ�௛�!�I$�Voʦ��=��ϩӛ�4:�JYɐ�}E�
k���UiA�֊�V�вD6e$�ip��u�wr�Ś��՞���o�+��[U0�@ @ZA�z���XL���<c_��~� �y�lȝ�U��b\�`u}���n����;����=Q����K��u�݇^-�M�ʴ⼡Jgh�r�Z�Y#ڣٹ�C���v�K:W_}�UK]�v�^�Ӯ֎��Ӫ��U���X�n�)C1&F��{:��gF��J\�B4&��N���.���Kx0�`�u̸����hS��9�)-6�bc�3�t�S6�vr��o���j͙��˔ꊥ���P��q�_�`:�Ƞ�V����zm�{�G%H%˺:�O(��R�'+�h�An��f͋uo����2`��VL�P��Ï��g=�ۍo�]�tO�
�U,�	�f���d�� �w��[�YR�#��7ϝo�׃
���dr7I��Z�,]�)�ƪ�+���S'T5��)e��˘�3��c:��Ԭ�68k�cxÜ��*��F��X��	��Y-p�����Я����e�$E]��vi!�]O�ű@㸭��vv.��7@�F���f������ea������eϡ�o���W_z��1R�ZfK?���������������~(�tf��A��@y��{*�\*�ȝ+oF���������;,eE]�q�����ݘ�Tk�G�@�lqk����"!�{�N�W�V�sHGn�ͮB�)��yMe�ܪ�����"Z3�]lQ�]&���S�� 7� uj[r���9�;w��{\�Ї @/n�IZe�_�;�zk'B�ua�����,���_!Ǣ��t��	-�<-![pj`��:�"U@�ʙ��t�0��>�*�� #sܘ��[�]n�{yi��[W��ܝ��cZ��{G����#x���{1j�׮d��&�i�Xێ�������z�7�����</�=�ZP�UMZ��^�ԃc�l6(�ql���܅��۴�p�顱�2U��8!��+�����8s�h��G@���
"�v�mE�d;}1�SK:��m��t8;U�J���S���J���6�m=r�l�n�X��Ւ�T��[�5�^���kʸ[�ޡtq����&���Z�Y�d�;i,ѻ8͕��36�%i
qX�
���Ե*�s�6E��˓������t�X2!�}/���3!!�S�b���eSf��,�����Br�E�C��W�U�IR�~
^��^k�/^�xum��].��g���ۻqq�k��f��R�k]^8#3M�P��@�u]�mH6�wG�dWs$�=�}Q�R潐p�a���u�eO��F���]j+��O\��z3]��G�f�XM'�'~n���.��Z��Wn�"��T�I�Dtz����:󕊛�o�;�ݑF�h����h�l���n�t�EO��1�R-J�����JE�I��h�g��f��^
�YQѮ�GK��4F��M�Fxܿ�Ʊ_��I���.����t�x��ӳq]���D��a����q��et�������^6��w�?N�����塩��l�XK:�N�����¨����x�"����j�ܓ�vM�9xTޤn>�8i�E-X�
�ڿ�4ې�W.���}W�B���<�g�>�8�y�O�<|�����{����ˏ��^a��`4\(���P�F��3vg\	اؓ�`cUͥ�>�$���z��wU�Z�d�1��
��*�1ˤ̻ѳ�񭁾��)@V@J'Mz-�B+y�7_�<�G���ɍ�}�g�'�[Q"6���^�c"}ѽ~j��#���M��ɾ��W�JЭ�<�����,�W@�yn"�ȼD{MIyNi��,���~��I�
����y\���	롙� �k��sYӣ䝼�ht�jt�p/��sz���Uywj����1tn�v�jcB)�;�5j�V��N
�TZ������yՍhZ���zgA��u�����U�m����t)[��:|��QSh ��9�����Y�M?��s�S�5�@<u{��)\�1��ޓ��y��Q��D��Mʁs�ؽ!ӯ^��u�v�u�,qT�r���)��ՑsPs#H��øﳹ6������z�b[q��>�Z�AG�r�Y�N���?����uB�|��v����f/e|G�ЊN���}Ŀ� !Vz�T��홃��w�OW�6�:��y[��5]S���!8F�t�Q�������?�wV��O���yB�U����N�z������l~�L���ٽV���8M��̍�]��Np�n;�{�N��p��k��*�L���h��C��t6
�;y��$R�꾍���G&n-�9u~�jR����)�>d+��"B�o~���i��]^޴�sK�i��gwD#�����@�f�\����J�dǝ���~qӕH�e�w諦�C�3Ȯ�"��D�8`��`��5g�wH;��Vx�"&H.����E�O��x6�[���l���5e{���A���&|�7K�����%�����jf;#	�B��<�b�!��Ĉ=N����Jbfn=̀h�w�h�o�}/GM&�o�f���-H�<��'�ݵ2�9�3�}�se8�q�qU�T�2m��nj��/-80��Qv7ԑsS7eg\����{��0�-j��ofa��f���QKN+�Ap{Z��&�;��q�����f�h�FZ����6wA{l���ܑv�{:�����g-�g�Rr�,�ס��硻][;�+c�\'ù������!�t:PT����1!��H��\=~շ���G?3r�ׯ} ��g��z�N�T�+����e?}g]��՞ho�~�m�-�[����s����!�	�g�a���<l�N�k.�W�M�D��!�J'����o��H�^9�2��oHI��U�C34��~�[4%���{��{D]�Nq��S�]�/=���9<IN�*���8���ji��M����{U��T�Q��)r3%�w1pw�y�ݛN饾���#^�Ȋ'�������%^
f�3�%,�&�Ύ�}�C|��dF��<����F�C�f�p@�O����Q�羞�ܖ����Ƕ�K4���o'3����Q��Z�_AG|#�Dl����>?Rڍ�\(e���Ô/�K�U���͌�r���[�P;oܽ�4`+�o�zR I�w�k�H�9i#�zVD��t����v�JBo����ój-��e�^j�ל��.itFL_+̢�8͛"���0	o��D>�1�X;>���i����P��s���wf�V\P�ͩe&���H��c���	E��1[%"��y.㝍P������o��CP�7hП)�����2�R��h\�ԗ4���8��/�5�&h��J���G^s@���n��=����Rn]1�����bi.��W5��9�3��^"W��.�gcm%��E�����vr�i��]i6�e!@e{�`�N@�k�s������1Z}5�5���@�qN�v37l��I�����d~o3�d����8ߥ���7�_E3�G��9�*����/ݬ���Jq+�o�����aG�M�gD��w�W��֯���ʹ����IΪڭ�v֛�*l�ilb�7|�P9�0�R���z����<|�DS1�s`������QJr:Ŝ�KJSU��骛��Ǻz�<��6Z$J�˾j�����OB�|��򴽓�C�q�w�G"�=����Z�����6�����{��_A��K��Mj}&���~���Ƽl<��:j��2����4��67�y�Nx���y�w:�U�<�e3p�k��������1F��Y�ض�2wiy�1_�����~޸&5�Zb�me�':7B�tB)̋����/��$��{�R�-��|�~?Y�hze����>�&�Q��i['+$msU��cdron�P������o�}=��V|{z�C~��r��aR{>q��a�&�ǳ$��pz;��Z�
��^���u����d�B��9w��U��^1K��u��آ���X�Щ��{+UN�gio��r��&���*�o����am�����7Mw]v�Sv��]K{�n�T�yƀ6��yض����9@�K#��nԜ��XDdo(dlu�b���:*�dgT��ѫ}�k�&��@�ɕ����#����4n����yo2�.�k��4����T��r/P������m��G6kΛ��P�D�9k�F2�Q��s8k����e��[�ղ�ۗA�_7*���}�3����c)y��O�"�ھ�NX�Ϋ���Nի�Q�UU��&ݡ1�L�y�+R	[Pe���;V�>���.(�1��@�Ƙ�w)��9o�(���N��b�+�<L�Æ�n����eǜ⋆d �i�r"XΈ�}5�2O������H���s3��:7���1Z�+��2��r5LD��V��J$�l���ݛn�/-�=�o����Xf�+�P��)w�EE�������AP����[:���sU\!�>�1��>\��cn��
��u:8��{���s��^_w�X�G����r���s�}��f3�Y����͌��w�w�s[�S�����+��bK|k�R���W���Wΐ.E��h�р}%�|5o��O�X������dt[�d���k/΄��>{�)gr�w� �qsh%��\���ݽck��WX��e���)-�r5�UtF.�F6Upmb��];��Ln���ct��9�M���X�lY�vL{.��֛Y����9�e�)�W�Q���J}�{��]{ޚ��vO.��9��0�>*�zzz�0:�}��#W��Y����n*��͟$�nd��Q3>��P' ��=�}�]'�ק��7��>t�<c��-�N���]�����ٟB�k<8�%� ��0��7�K���W�zG�3��غ��A���6�-W����Do�=7���/vU�3�d��T뙏>��Ϣ�橱y��U�+�ʛ�ø��6��N�nAJ[U}���Q���q��b1|Y6��Q-ʕ�R��ɟ��!^���v꧊!u����=7	�H��-�u=��G�:b:�����|~_D��T6���\y�܈���
��=�Fr��]u���LOV�Ow��P��Vj�@�S���aj^�ڨK�߹����Ѧ�+A�u���=y�~3�{uOI��f\&w����}����^��z�71��K����������@��wb��##�Q�0��'$���'�����6�ׇ��j�o[������-�2����#˫|{t�m�n;&�|1Ǥ������uC> ѕ_�5�2�� ��Iή#@���M������-=͚m0��b�PݵQnլ�\\�b���!ΠK,��_*O��!q`l&�\;����O���}�p٤ݞ�e񤲀[�ENV�@T��^�l+�ܹj���M[�i��F��՞�!��U�i���>�uOi9�=��#�"g˦#w�e}����6i)��Roc� ߶9*;�/l]헷���{�]|��w���Vq��>Ү!	��e��m&��?5��s$�� *bW�W�̪�W3wu��S�gg_�w:r�\���UB���/�1��F�_�˼����qW�ez�l�oiܳ�}�V��bsg�E��ﱱ�t>PW��?h�Փ�7�]Ƽ���O��]J͜{a0#�4:c*����佞W��7����{]��5 �ח/q�ȓ>Faޝ���=����=%0K�IqjP����l���M�DI�T&�x]Wv��A��k�K�[���^H ���M��۴˩�"�\��Wǲ}Z��s�����`:#5W�O_3<6ӧ}�w�1f"#e]�R�莨�����N�\k�I�$w�ԟ%��%��v��Y�2����KF`SU�j�Y���<_/ݕ��%W7߉3�V��X�5�L����Μ.��'ʯ����{'�⫫ccS]Y䏢��j���أ�%-J�/h�ϵvK�����J�����i��ee�Su�s�u�9��U�u���;�7Q��WPB�!]�3��E�&edٛ)sݵ�o��[/e��k�����(=�������y�S/V�6�i>���w�qjZ< �1�hB6_m����:�.���R�b�v�+��.<&�/t��']��Cx���oe<�=�`CWvS{W]m�̄�~�
�t�������������24��[��鞮�}�Ǆ���8���2i�7�^��:��/��_*�YQ�%�6�}N�\�ٯ�z_�t��~[|=����o�׷k/萞²���}�k�����ѷ���/'��&֞��{�Q��n ��	K]@3-(
L-����X){}�tTӋT��P��F�^.����y���p���E��w�����A<;B�����r��!��������\�"z8u@��\���+��È�ze�ޟu����Q�Ab�0�e�?���xe��z�FsV<��ۥܲm�DH{9�x��R��ҽ�B��jD�M������/nzcc��J���� �����J��td#�
(�Q~{X���l�7\��h/��������==�v=!�����D�ys�2�X�p׉�ik�=f�5V�p��->�ҵ���bA9��	�ze��{^�w�4��-���\�:Xhws��Z�����k�J�3ݎ�4�wkh�� G�j�W��d��-n{��7غbYN�����mD�h�˷h>���,mqYS��F�Tl�[5v���[O��+�*��u��}�=Qc���/����w��(��B�'����"�5�V�y�
�)yS�.�!��m�Ԉ`��&�&�xs:��[ۥ��+Z�ƊW���m"�� `���y�o��
Ad=��;��)�ώGFe��Ƀ��1S� ��-Z���ޮ��F�⚭��B�d�ܘ�ul6�&^�"��a���t��p��r�S�+�=��֪����]�Ͻ�r���v,2}��e��35]9'�Dl��୧��t�z��mv��I�CHp���:�NV��q�\��  �^J�A�Mz�r�0۷��z����̤��׶��:h�=�vk��ĥ9�'D73[��_b�띞��A\��Ky,�&ʿ��F�+�s�Ժ��C�M����xv���^�YV���4�y+��H�~���ըL�ڀ�F\���mLT\���N0kRH갱7�x��8#S�3Ԫ%��-Es�u�W��DW��$cs�} �,%;f��>Y()>Vx)��g�3;�	G��ZF��#"<�z�������uU���G�I��6|9��M��D�N�or�&O�����95G�o�&���n�s���ҕ�ȱLVm�Mi#6//d��w}�ö�31�,j����ڽɭ�w#5�!�M��a��|g��l>�q����Bg��ꣽ�;��]������^���iKN؏�y��!�j=��;���V'�A]X��N�;���B��,�Y�����&�.o�l��c'D�:3,wvG����)Ų��.ݩPX���=*_�4��Go�P!�-��)V�]��v�����
�*Y�!�ʽ��H,�t��ɏ�?�ĩ��.�4��c��Hb\�o8Κ#�������k/�=3����Z�[�̿N
��&�4�ph�Z��i��Y�U;��ƌ���ݜO������)RU�1�������E�Y����x9w��������������䷵�c��yA�V�{n����+w��f{O�~�G���<��i���Y�;�,���<$��vF_�@&�I�{c��É3�G��3�	 ����iWC<4B�a��~]l,����wt݌A��*n���9�ϓIp/N��N���T� �b~�)�1��5��F�̻:}f'>�U���S����w��`�D��|��~[4E1!M�9�r;r��G'�SO#��[�碱ي�܋����]�{�.4��Y��N�e۩��@'��W���U�0���7�~����5�//���{��%����j��!ê�&gf�z;kg�w�s�֫,�fm��5韗�=�������3w�*��r�[5sQ+����x~w��vaO]@��K�Mwh�xT\��٭�v�f��r�I9c�rc��wj��W6�0�.�]�]o��Gu��Bv\�n�wI6ͧJ�����Zֹ��7RӾ[O�����G��!��(�+��xzc��z�Ma�)á�'��[��������V���f�uԀ��ŋ��c��V��h6\��4�of�qv�-������֌j��Oc��<�r��V���wg+w���eǴ4Tg6��ݴ��}�f���� ����_sO�kU�r�W�U}Kr�-D�����+4bU�j�i�2�����ф�燠���*���j��+��� �����3ة��Ws$z[���=NWtJL�]c��3j���IVi����ʠ}>�����3��}z�Ϊ������7|ȋ0\�������Jb�'3� 3H&u].$1҃&j�N4㬖������pw)�vnl�;v���BNJ���@�1��N�u ��m`�w��<�on����f�~͞DB+C���J��;�!��1�GW��MB�3�t�ͼ͜�u.E[�E=OQ����i\;o;f��6�(��M���q\���b�֣4��ܗO�����R�+��a�][C��mN{�QYy-���}���ݺ]wS����v�I����)���4DU��⵹+k;q��LȻo�3�b���ZH��|;V%�_#aPr6�sJ?mΏ+�	k����b�n��0�����>�N�r�M�xM�yʖ��b�:��ǽō�컕��yl�r*�ڰ5`L-okZgw��$��3xV�Ѹ�έ|����7��V�+�l$N�qu�s�/��$�8B����m�9�NMޤN[:%L}r��Fk����C���Ԇ�Zͱ��`�'����.��z.��2L�mU�t�s�ޛӥ$Gf�����u+������d���'uV۷Iw!��{���Us)��YI=�}{���Kl�����v�ܲ���U�|ԫ�S�Y�]%�jx���	ΗU�+��[5`�)W<�|j㈇��u �N��;�=ܦS�5y ;��0�Dh�M �_`d��E)ܗ���	F¾�{3&�O��ֶ1�����)��jw�7�g�t�T��J�ޛP9C�����_ue\�5=� ��y����'.K���n�ݓ�.��zs�Ļ���GA�*\�N�''Ƴ��چ��:�v����u:���ӕw,�N�՞&mwz=Ӈv�n�F"�wU��<T� m%��y+�0�
WJ��(^��m�ٳS��'�%X��e<�/E%�3��8Np[�}��%H��_A���V�G.�k"3hA1����Y����Ƒ�xGf�S鎗7}���7F�<�w:�3ƍMV- �]�EB����}b��T�rX�U�+vjs��0�x7��\�鄢$�ia%](�r�٢d���B̸yi��],�k����.�W3��e���W�F�	zin���U�Լ!e)�a�s������qB��v9b�N4�Cz�U�|�m�̥y��%[����T���(�c���b�e����c�z�?#xT�5�6������߲%���X��<�7�Pڶ1��N�`��p�Vq�y��h����o�]a=��h#X���9���Lf�X*wmsg���M��b��~��u��t�wR��z�Z��������1��uzk�^ފ�9#@���L���Ml6�;�p�n*,�"uq�X��#�[�=7q�b�)�v��0��8�wd$r����%~['�~�%o��.�wj�Z��|6Eo�dɀt=3ѡ��cz���e�5��ӯTQ��l\;��ʹtR�ش�Τ�X�����F�{��V�ri�N�{�B�RAz�t+}�.�xu��C=�2���N��?T���+�;nl�(�h�����z��b�Wc��j�EcA�܉�F�6���sόP1���r�ڱw���o �>���oǶgv�m�qCbĕz��۪��Yݷs��"��ɴufm:�ʡ	ٟ_M��Q�on�����8a�*���k0��v/7�k�K��<I��_�;�uF��g:�����2����wpy�����.�c0�vv�$��:��]o��<)6wo"}d��~����%Nه'��#�K:�g������f:�L�5~��;��J�֜�.�l�J�U���z�(��)�FZ8ܼ�&K0��b��=z�����u-���%�֛��5qn#uw&B7������6|{�%���#4��.K_���:P�]]���y+���;��K�5J�8�Y �V�q�9�r��3���%]Z�5sqav*�c�s�Z��H��s��<k��ȯԬ�b}w8�q�������F@BS�nȖ�P�ν8͆�ؾ��;�û�������7<$�v�ة��z�����Q�	:�s MS�|N�s�xw�b������:fO*�X�׃wǝ��M�!^d�2g�gp�h�x���I�mM�磃�W�#̳��5���ݣ�{�I�Cˌ�c�)��W�����zcJT����{|�eM�P乇�s����w^]��J��ԫٞ��ɻ�L��'����ّ���|rh��âR$s�}���N��هT��8�VC�Y�����ҟ%��1?��:�2'�s=7+A�RM7�-��ns��"�gM���y*��d�Su��τL�]Ϝ���ЀϺ�ġ�W>9(����ߡ@��߁s��k�������ԍ��,��K/a����1v�]�]�OL�wq������W���?=��6��t-{hVTx{#v7*��?d|<�iT���'��M�xS������F'7EYT���؟fyM��[��+Ҙ޻��b��~�+`��>�YG���:�b)/#~�N�S+Ru;�r7SA������R�l��y��(��IN�l��8%�մ{�tj�՘���ve�v��{��Tn�ǝ�)n�=��	D����Om�=!y1Jxi�$�a�œVn�4��4fޚͮN�+]�`i�LuoZ�AX��Ky��-�2c��s��R�H�%n;m�sOa0���{���VK�:��ا�"���LU.��p/n�Ɠ,EP��IM�3�Զ���/l]yz0X٨�GW�<��vX��.M� �c��u���-�'�C�H�!N��5��z�be^�=�vs����1Y���փ>�4]@~̝� �~�(x/r���ڑÓ]�h�H*N�.G���)�P��[�߇�;)+ůEf�T$` ���f��xY�~q�]��%��w�x\޼���W��n_�T.^���z���\^�Z?�6�e�TH���Q�i�������jM�{|AC�f-S��3G�tw�｛�����p���d�c�u�Ѧ�Q�ʩc�"��k��U�i�� �;r���mA��ús�5����x�t@��p�z��ف����=�|L�z�*�Hz�SAqu��M����}�2�z��v;��k�U�{ty����^wG��-�Șn.p}�]��vL��LS��)�ұ�)��\�i�c�M��w�b6�Os�y�F)TN�fqn����&��#)��2���w�s�Z�%���
�Ղ���!c����j�MWJV���
����b��1r*l�s6,��u�9ͬT��?� ޢ@b��vq����P��������v�RN�_2�h�υ>̓%����7�N,]��fl�h�W. Q�,�-�4����j���IK��S��݉� 37|���ۺPQW�����绲i��fU��P2t+��L���?�6�����H�67In��-=,�fk+�i;>(	�U�cDe���Ĺ�0����]������鳛��G���i���NPen��$����9��zr��j�"��ծ�f!A����,�+�/#�柌��u�f7��:wÏ�H�4&�_'Ĥ>W%��2rg�9Y��ߪ?q��� ɺ�L3�qJ`̘#K^.I1�9^��~�bB2���2�x{�;Aʗ���U��L�!�_�&��ӓ��\�N���� ����Ms�W������U��e��^�2R�s�p���S.ם]���I]����=�5'�Ss���ߘҭ9��X��)N֏�����M�t����ή{'-��4��D/nd"4�qAr��Z��n{H$�Sog�)��$mJǳB��Y������>�S��a�]�u�O���f+�6],���+"A�t*�  Jq�R�ǆ�p���ˆK���SP��ꎯ>�g��O��{��+ԗ�	N��3ya�@~��7�v�x��o,j��W��(.��w�@9|]k�x�*�2Gs��� ����Uŷq�d40��͸5�����	v��b����i���ީ�xQ�\ɯe_o�t_�o��>�a�3��8~���MY�k�H�2����{��>~Fs�vz:�A�����{7f��+���̕�p��O	���� s��U>��[f���gb�]�y6*�uL�����o-Vړ�6<���O����\�XB�@L؝�9����f1�l����-^�ˊ���\����V���w�l�7}\�3GKO���7L�
���k因�v�[��5�i�wz6�n�
ܝ�ǣ�Tu�^k�h?W�]d��|�<v>�Wq��׼ی�>�~9��dk�"��+MOF��~�ٱ�a7R��u+�W�{f�}" ���g�;�i˾u9˾�O���|Z�J�pz|���؋Z��f��w*<�-���a(}�Y������}p�φat��d���3�D8����nL!v<�� �}���gZѕm7��O�e�xo��L�th���I�VS�Y���ī��S�C�5�y��;��[SЭU�%��A���k \:���G~��D�I�Vwd�& 8YO��(�xj��F������q7*^����`����(?l�F�P@8�r�'> s�w�ӡ��s*�}�騎դ�F�|��ue�}6����[N�>z�:����p�w��ζ;7�����>7y�:�re*WZ��Ro��]fX�%>Z+u��˨��;���O��oY����+�s۴���$�kp4P�N�x��{�OM��l�fK�s`�ׁp���yc\���/k\2��ۢ�k0~��ڧ=��zR���-���S�%����yA�:e����}�н��S9$��t�o��o\i�(�����Q��O��������_z��YM�'k�m�_�y��R��N��쒉�g���_� b�v�t�������IcB���S�O�nd��ᶅ*0�^�f�� N���a-��hQ@o�k�j�(6y��e�Y5=oGf���
��%*W3U2�֊�j�8R]·�� �7��*@��DlKg�����̿gl½`^�2qC�8!>}}��.�C?��1����f��ґ;9�AyLnS~4� �BK�<�%?m^��o�,v]�۾��=]N{;�EW{ �L���s@��3���	yה����˘��w\�%zǖ�t57{���b�m�%w � 
%=��:rl,�&�$d�L˷�{Y�YwOx7:-���ڑ��=X���"��1�P�F���%HF�
>�a�:�����Uɹ@j����ݔ�e�����yW��n�`��%��%]jfZ�B����2�vܝ���o��W����F�t6Jp���_FP6�xE.�N����
9'j4:�\�Ws L�v�0(�6V�B�y��۲;���z0��e�-�t�[T��9��e*�����7�zVJ9]�٨��Y*���h0揫;��{e^yy,�m~�9=Vj�/C�M�?x]*�1(x�J������ʹ�a�ލ���!q�t���ą�V��C�~����]	�s�îq&d�n��8#�w
�횭���.��'��4 P�;ۗ~x�e��z�IA^�ə�_s�=��g�B�3�y�Qu1��r=~S#�����\�_`Y�*/v���nv��=��c*I�&���,������?��Mv>����Ha�R�b5�Gfp�w��ly�g:��]�+����. L������e�1�0쑯��4�Kǹ�[����]���WR�M��V�G��n�~��~�߾�oMh�t�H�7�y�:ps ���	݈���#�r	~W��x/+~>�F�G��ˣr�j�q)x����|�����*@B��I�+�����r�دDh�x��*]��d��{��O
\�9M��o�M�=q��S=�1մ�ɂ{�c'�|_�hP���{��`������o0���$�d7'G^�V_�x�A`��(�PV���!M�-��j��������G_a���V�%��gt�Ź(f��$�6��|�n��P�z��&�"��|�c���o�\�#��U̴��Z�C���5��Y�n�V�����I��?�e�tM��r�Ef����Ez�R�I�v/�=ƯJ\v�T��^��I��
�m�˫�{�kz_�9�_)7��v� ��Z�4�Tk����G �ɤ��ꡛ��y0���C�.�-	�ȣ�.4�c�g�f���y���}����߅WK*!��vc�;n������ڨQI���?*Vf,��v�a�n��>�����wr��cF#��^U����G��;_�\�,+�I3��ln�#=�W���k�s�o ������T�xK��yAm�^N�3-%xƱ�G82~���w�|Ua�}y=]V��OW.�ދ�܎�Z���#��'��ɍ�#����U@-̾�eyDw�{{4�^Kn^e�P�U�V]������Rp.��$gg</<�]�łd�.����DjUC͝9@�fu�"�@�}����eWEW9��'p�lZT�ouJ�\���%/#oG'^Έ���I{w�/���3bl_��W�pc5aC���3���SZM�͋����|I��w὚O�w�K!R�Y��O۲�8�����Ui��a�z8�qUoʁ<���[j�͡iSu>�~CS��?�7�W�Z���"X��w&����`k�Q�ZXlVSImvWu�Z�R��$_#Ҥ��yė6a�ޠv=����M��������ս3�Y�n:̭���J�ާ1�\�-�p���j��O�Y�g�4�s7�Jx]pXD��侤TPV�����fp�ߎ�5���w���K�Pՙ.ު���=�;.d��Lo��}�?�]�{ʮ��W3ƺ�dh�� 8.U�2˞���Y��eOJ�{.�Q�tI��چE���޸z����Co���� T"���R�1���н1�҆����~�O8�՝)��,���X����uo���X��)�ā��� �g��kJ�����nݷΝ�C]|lo��sr�#���m�K��v��
�T/�d.�'5,M�@�I�G��U?>�Y�ȩz�R:/`���~ܹCa�-]Ϸ=>ݢq��"�H&�0�%�[�qn��`�˹֡�[F��N���!�]C��M�W=��;d*|(�q��œ��5P]����[K�����)����k�ٝwț5�ܹ���Z����}�M�,��T�]v����^35O^Hr�x�Z>�F�\�n(�����y��F�hS��뚾m`~�V��[��fy�E]��A^?,�D��y_���:+c��ø�'ˣO��B��v�LP�� �:�_v��O���k`�jJ���r��i�R�9���D�+U��z����U��u�����ӝ2�A�������AT�������%�� X娼��Q��]6u��z��^����J��������<��T���7+K6/\���LRGk�����e�;�.�c�<�DEap�Ą���N��&��eS��3����C �^l?F�uX���޸��S��9��[wP!(7jv�-2੭�!���s�>>ܓ^�����R��y�&Ao��|%{��X�Ȃz=���c��3����kC���c�?j�ע�~�G�ՙ�G�D���w�HPɹ��:�Q�=kϢ+oh��Dx�;��͜B��t�ѵ�b�9��~��EІ�ߍA�iY����p�z��=�ݙ3.*�X�nXXP���~���]�z��yC'h{}�%fZNX^$�|��Ƀ]߾Hс]��v��n�l�/D�i��7g�U��l;���'��7� ����)x�7�U��.!�����Z��}�hmb���)4A5�?
$xn'v��K}����)�������1���<_��iȕyT��x��w������C��N����V]M��q����T=��4iF5�������A�����ٵ��y���w�ayϾYu�.���X��ޣpL��7�&g:��o�"��ݾ�<��\�^Ïju+na���Q1�	ql�?p�<���6L���N�W8����sk={�14_�����@� �Up��pW�i��3iMJ=�i8�Y۱�]@1��h�(5u��e&NůF��{m��0��ٺz�T�kf���n�^wX ��'^���;���}�5�q�sn�)���
/vb�+j�27+�q��s{�cH��D��������J����W+��*��[��DA��_o������qL�w��p5��^��R*`�^
X˙J�ܫM��}%a�y�6(ud17Q�@�<�c�]R�֊=۴�E��Pڇ[���K�X�*�So5�!���X��cx�¬�u���Ma��U㊞ފ��v�nC\���Zs�sO̲�QKd��pf��N��D����1.VB�֎[�u��Yj]�B�z����z�K8	Oa7;t�\�!F�}O����#>�="��(p�0�\�C��V�WR�{�]�j�P�*���H=�l��H���i��hκ��,�6��P!��9���dE�Y�.���LK���^f�+��b#u�5B��W��Sec]	#E��ܔ(�={ߛ���O��G{<�;����G�8�^o �%r�vQ���� {/"[s��l\�p��ΥIG��Vj�M^=��'w-���*p��������q��k�PӯLW�� �[x�ԥ7w2�EHN�υ[�q�Zr�N<yZB@`b�+����W��[wrV�N�[Z��R���^9{�ڔe�r 4����Mڡ[�^�=V�u�{���s)��1%�f��uć��}VZf�#��b��rnr�AHWz]�\��y����uթ5L�[����f�2��Rܼ�O��k��}b��N�k�9�o*�c,�����u�V�_�ͭ�U�wR�ڍ�gr���45_|��4��M�4������ê�un5�0�\�wGA{ٯ�r��J��,��݀�ifr���"�8j���T��n5ٖLT�ug;�}+{�'}1:�t$�v�?5�G��$����W�e��K_�[��!%��*�������h�q�V�fu��ʶ�z�[���G^�XK@�2�DMӝֲ�߸؛{~c�/r�5�6� �;8�z�6��6܈��֮q�7���c)u��Ij�{�0/�6G6�+�{�������N2
��E�=V��փ|t��,�>���3���=nWU�q����^�+sXmV����
`��F,.n1Z7n	�ț���3�:X��U�/�;e&+�u흀\���^�B�i�n�����#�υe�e����w�������C.E�P�.W�awt�Bɛ�.���Fa@Yu+u�b�ؐ*E=]U#@a�34�Syd�G��|�6�ʉ�����⛂-��m�Dx��b۽���G�/�7�T���Wgi,\�C��vp�r�6�� ��h�.���]�f��oQ3�r��Q�]K�Dࢥ���\?���ꠡJYͬ�ۋ��3���jUɝ/0
��ͦ��|s�۬x�8��U��Ҙ�'{���اw�J4���M��Mgm��k���]���b�s	��҅\�g'�WB�tE�}?n.�K�ЧvƩ�߰]����{^I@��}��z�;�w�U�����')��`�.(��S����'dV�QS��Y�^�B׍&�C3�**(D��R���D��Ր��w�����|s&V��ȇ^˹�V�KBT:��l��x�qEFE���՘��"�ʏV���v�c�T%V�a�u�E͌�赚w���D̦�jm2 ���f��n�ޟz�i�j�p��o��Dߠ-�+�u��>ܧ�g��ܟ����[�3�ԜQ��rXt�>��P	S��g��W�)�S�ټ}����G]��0|{1��՗q�Y�8%b�З���67�?P�O��w�c�&gNIXy�G'�2����~�+[�M)sY�=K�_�1z;�eڝs�k�;�P�U�5_��%Dϔ���׋�\fW:�[�W��넲�ѽ�~5�^��+�q�lŁ�Q�>C9r��Gޖfd������S\&m�
V�s7c�N��o�����g5�gp��J;N�m�k�^Uj���o��'��H�)B��ڝp�s��B:&�iB�� F�H������*�F�\z�hV�}V��(!Vi�1�u}��h�����XAҨ����{�Er���ƺ�)`��-{��Z�V��tU�����I�n��-�Z���+3�]rɰv!���==�Fa=�y���[��Nz�����e�EN��}M��*�#C8��+�1a��q�g8`�
O=`X������W5����ϼ��O�K�� T�1���h�~��@�g�W�ݓ��|ek~/������WZ�nȾ�����8;ًE�7X������q?e��>�����]_�DtJ�i�z��o,�e�XW�%ßO5F��Ǣ��]�d�-��Sj/I��Mʙ�t�m���C��ݸ^dbɊ=��/-
s`_��Tl��Y7B�Kl?JW2%P�<b���Y*x��xE��DG�1���^�2轅��4���p�)�@��;��V��f)su�;�&��g%Y~[�O�	���9�>4��`�7vVm�͗¯*7��J����ֺ�B�l�댭uB����<w��k��`�\{��b�������M�{��n����r������:���^<�
#\�]�=yn�`)�Y�s�����_M�L�^g0َ��Nx)�D�����a��j�f�W;��
�w@n�Ŀ
�w�d��}?�{f�w�,PN�����6�fa8�T��}έ�u��b�s,%%kC�f��蚙)[���Nf�_
����K��q�I"�o);��۰:n�8��ك��ɮ��"��J�nN�7!� U�p��F���Y��"�2bzCemAO�]Z��Q�R!�굿��V�ߘ"�~wΣ�#��l��}��5
"�*N�⦮n��o��q�Ⱦ9)`��27e�=g=����e�)qz:�fBۏMo�=/b}�I9��#����6Ϳ'��U�7ٌ	���v^EC�Z��g&U�	Q�V�����8a�o��{㚅^}��c#M�S�m4#��"&C�X�����G����Әs�uN�$"8+Yc���nB��;�>�vr��õ8)D=5���"F�=T�	��ޗ^�jYɁ���U���7�:�D��w��g�|G��1>DsP_^N���\�m��r�]w����|V
��h�e�뽨i�p��P/���1ٰ� ���=O��%Fe�;��¹�^h�1{��=�齭t��O-fJ����_���`��Į!=����F��g5)��{�O�Fx���G{�!�A�ۤ���~s@�ܮ���l3���&��H�i����Z�A��`ϛ�����,M��ᢢ�q&��FRj���W������L9��޲��b)Wҥ�"ă�����^�ؑ�g�)��ڵ3��
�,:�\�qU��1�of�}6֔'t��;gvM�u.�F���;
F[K��r�
���w�Dvg7[ף^�Vn��k���^9.�ws�����nbߌ���F�f�خ��]���Z����q^��~}��/�$�#L�G� `�#:�yO=�8���u%�]0aOp9�y�x��������·e�gk����u^
��CH�;�6Tu��O���rPv^�<�b��������x_��}��|/ܖ����[�zκ=�u��=o�*�v>ȍ��'/�m���$��\���`Qb]��*awr/�i��n_����C���̲9�����4&:՛ӟ|���T�{b����t����-!�قo�^x}b��h`9n�`�č��S�R�W(�ߙ���Z1W�~����ʗ��O�Wk���v���hl)�~��:=�{�]I�fxze3�����-M��SdW82=� �uvU�1J��ԇ�pLw��/،��zxW#9�������+�ӟO��3R,^R�b�rþ��\vXq���y�g��{�M�n�e���2��e����N�����~���w�V�k��6IQFǖ~Nk����n�/'�I*�2��o�ѡ���_����n���V�#��,��:�Mj=�D�/�����|&�(��ς��-t܃V$/�k���zq݃A䱥g�o���� r�{;7O��}���&�f�vV��4�;� ���;"�\�v�sm�z���v2�n]!4ME=���H�d�s䴨��}*k=3�}��E�-��o-�������q���K�f�1@���/dz+'���Z��8���I�H3�x;���1���F�^�N��k��	y���TW�!�c,T���f�ʺ���-����2S�X����OF�=YY�vqDv 4eLl��bXwP/p�Ę��G?��������yW\���t}�A�y����7�c��qXIs#̟S��q׭�����P��۷	��,�7��h�R{־յ�.C/�ި{q�����	�̓�v�iZ��y$}	mt��E��w�^.��0x�WH���'���1n;U���HM�N�ܫ�^F&z���2�b~~�^�-QŢ69�L�)s���:L�qѯ���q�c�ؽ`���,���%9�"h=x��]�� %�k�ԇ�6���}��~.�W�R��+��h_9�Fg�c�Q�ݓ��ZA^f���TĈf�;�hϤ
�US�;}^�Y�\��@��+�N_z�L:�튧WCn�8�K)���q����iu�3|`��R������*hS}Tnz}��{r�[��f���=��n�u�.��rgk��A�]}�
�; �!ˉc:3�W=
��Ѩ�p�D�Nk���u�Edk�+A0k!}yeJ\U�i�̂��Z�y��)
[�2U��u� :Mu��;N�u�0}Y�n5�7�����+�C�^zny�[wk/7���W\�>~�VF�	���ڍ6l9fߑ3-c��+!db�W�IQ���0�-{a���kǞ��'��闗��\�w%����K���i_n�OĲ�9�5%(�U�	c�o��'���Q}\���Z��B�Q���G��7�^gf-^:�#�]�-w��Dbه�G�ɸ�<7#��Q!�n^�ޘ���^g/�9畺�^痕���hm�M��i�9�;y�=8�(�ېj��(��l*d(��RG�\��%�Q0�T���>�>��4����rz�~U��/Q^��|��nK�w�],{1���W��ǐ���@w>��veS�"<�خ�uAZ�&��P�i���B'1�Ž���p�������/qQ��*��2!d��A�z���y�j9�$&S�T�Li��B ���+b��D!�OZ��P*|+�ո�0̚�*=3�hO=�u�P��;�f��D����'*kp�9]�W�"��ّ$ަ�c��7��f\D��yfjŘ<���>o�lD��C'�����d ��3/:b\���^��s{�ڲ�Rq[)쳚��Ot�'7�^"�	Xd��Z���:u o�W�t��S��;�]֭Y㥽�R����QGv�'�8��9�d2k�7�,��Mjm�
�U��m��s���֠�f�s���i���&�x[ʸ�EK��ڱ~�cĮ�"�c`q�.��}o�}��|�/'t�z6q�57Ug�Е6`:�_,��}lv�Z��涰�b��G8�o�90r��=׍�&�fNCo��o��зr<�ߛt�Хe;���İ5eSۈ��j��On�~���{{Uw����ȵ�3�2n,�/�7'��,�tFn�~"���;�,������H�#����z�]�܋
	��>w��%p>�~	c����ͳ���W-su|yzq'}��ʍ����,Y��L��]������^���W��l�G���"��j֯J�����u�O%|�x�9�)U�}���顕�o��w��#)��ur�]w�_]��a���L��<S�OEE���ᇺ׮�{��1�}G�Қ�+*�`�L���u2��،��*}�=K��A_-BM�'�*���p�Z�o��:����ֹ�7>^�ϑS3�c5�}��Yo��|�X�=^� {�r��v����	*fح�&�:��,���>K䢲E�ʅ<{X2�g��gc� ���
;Z�
C-��&�RЩ�[7�}/�$��vTor9Fo)l�jU�u}�J��,��54���i5V�M������*3Un��xRʘh����n�@��)��#��}����HY4�r���e���o�19�e7�Mi�2AN8��
�+�>�u�}�v�˛�W3:9P~R�"$����RϽ|uU�]ww[��wV�r`�~4nD�L���1��N~���^f���λθߢ`�Dm��g6�N\^���}�� ��>���>���&�����@"R�3tOO��]����:N�ۚ�K��$�OY��Wޕo�as���Mu�z�:���0x_z�����]`n��&����d����0W����%`=;��^j�I����&K�6I��
<Ufb���Td��Z�훯	3tT�V�rSw&`t��̕l^�GQ��ބ�����w{(j�aT-g6{Wc6����@n(�j6�R�:;ΖQ�[�t��+k�1��/�Z�ۍ�t{?t���n@l��^�feNY�w����d�A�nA�G.-b��%�&��mg�5��+���uw�O1�ۗw��P/&wa�F#
�-߼���Uw��?3��&��?g��,��J徚��#�-�����I�N��,�j�Ra�MqI]�Ȃ֊Ѝ�у�P�=�'�2/�Z7����z�5C�év ���GVG`.���7;�}�P�z"�]#��d�')��N{R4�`������sŋо����e?dS4��l(���)9��*p��R�Yy*�z�<�V'�m��xr�qF�n����^W�AS�q+?D��r&郪��t���i���)��o����Pw���u0��*$�p���PvN��D��i�����,�}��̯���/��)��1J���o�l�T�^+o4h�ʽ��u�} b��#]��e����``�r�6�_�^�Ȯ��n��q�����W�Ն�l��@��S ӠNQ}����5����>�ig'/���f9�|z�h_�s^��ة�(7�glS�y=<}r�]���f O+GC�`���t�r`��ޅ���>��7Y�1�J��d����Ccm�ӂܹ���֛����`���VOq��>����G�{3�^ӝ��AM[ǖ�-]�YK�X��ݐ����*���/w�bp5v�~S���!��Ϲ�'�s7jw!�x�~dl|��y���Y����OV����������U�m9�W�%Qk}3�Ea�-KD�� ���)��SCV�/9�\~~�=����Vɋv��k��-^Bo��_��1�0c��!����	�]`��0�=$ʱ�Ͻ�޾=C$*�އ��o�;ӬQX*Y�)�2�ޥ�Q�_�6]�	�|ݜ��O�W,x7A�/@]w�@Y��:;!�+Em��y|�qP�n��:(uYCw����Ks���C�9�cl]�)wJv�e��){E��NMZK �T�P�u���B�������FhԷ$�^�zv� j�[b�p���w���PDC�Ժ���};^m�߯���y$�f�9���hd���]M|	�\�O{[�q�pӱ��ҿ���s<�@)#��'2��W'�Q>ܼ1����3T������k��������&��}�R&�r�!=6���k6��p%����U+=v{L���J�x�~D�����
4�bbB̋��\���8�МԶS��YHX֦T%+�Z��-Đ����s��>�^y
|G��v��Tu߾K�s*n��[��o�)`���T�����Hs|��\��s��d�1J�㯯|�fځٛ��)�*6[ε�k��7�}mW�F8*F/��0	X!�YSV;G?D�w�x�zL��>�T4T��;���FN�v�/��1g2��E%7�8B��L>���l��f�v,߻I�*n������� ��FzP���Tq�8g��b�y�K{0�,,���?_�z%��rU�n]x�a��a����{ ��La�/K&:˘"'yWmX�.U��y�vgrS��~U�k�طa����P	�z�\��zi�Q	O��6���n�۵�YgyJ<����gp������6����K���YV\}�E�;(�NU����NY�_d�K�
��Ȥ�L%�w�W��Py�f�6�4�p'�QGنZ���I	�,���R�W	�vΒ��������[T�Z�0#��U���6��hw�k��Gݗ�],z,1k�Y�@M��%sn��p�;}��Q
�wj���PѼOa�}���c>���x8!�9S�<h㗻�U��|1=a�!��IFb�\P�B�s���f� ���,�����W]�4Ƹ������E v��!��2e�<}tb�{�]����
�z�� 	���&1R�9�8WgZ�On���m��� �K4\ :Fk+ l���g�7|��'	����f+�e3;o�D�K(å)��er���Uep<{ֶ͇�Kqf��<�{�0Rǵ��㽿��(̃'z����8wr[ݝ(sٿ>X�A���έ�쾜{�9*DF��&q�W}K�[�T�a�e�.�Ut�\+&D���3���Ls;z���AJ��o5�Jf��7��}S��Ք���԰��uw3�id7\GI�BPz���2QX:r�BX���Ni�X�m��JJ��0���9��˒nXb�.�ʺU���t���uӫ���Z�2S��"��%W{��.����pZ�,X�P`}2���;��ڬ�4k��y�jt�*�h�ش+)eVH�`�l��wj�Xd�\T{u����Ǥ����"��������GSYa��ЦV�̷���U��ju8��ni����H�Iu�M˛0�0�rY��_���s���Q��&��Z�� iݎٖ��������,�S^��b�݈Chn��@��P�.��4 B7�$����m�sX$����;0�ܝ�n�\��Һ�E��E�z��N^��SXt��j��`2����9�����X�
��{��qd��S���ЦX��Y�rе��	[����Xg	�����Vc�޳�tt��bBvu�Ck����}�r�%e$����rn�eZ��@O=g�;$�+��Fg-ה���:�aS�fѾ�{C�����\`����Ū�����]zc�suƋ�{��W7\F�v��e�oj{I!��Δp�v8�z�]�N�vLt��uͥMduj��u�Foi��u0`fӊ���A�A����.��b�Shbk���T�13Aƃ�u�����W׳���5m�|�f|�t��r��ɓ�qb���?<�\,mHdsE�ȝ����Gc���I����v#{�+��l�O�.Y2�~��+h)s�;����9B���m�&2.vv�H����K���tH���G�!D�ޗ6�XS~or�*[�$�t�4�y�������"&��v�z*�4��:<u�g79�&q�oL<�������:l��)ؔ�8���d�[2����A�� eUC
W7��	W����gaY�tܗ�X��4tL���p�܍P��*�.P�>8�9;��wZ�	3�Z��ml�c�ds\�N��z���"T;� 7� E]�;'ҝ1��S<2W?S�YHm��C��28�xS�o>�bd�����y��y�S�'5w�|�ۘ�I�^A~�0��d��.�A�'��PIlO�)Mߎ�[
h1�C����Wwyu�Ճz���T�?8��G��[֫gCf��*0(�ՙ�Q��&b�mm8�*6]�j�.ӕCdS��4��<rE;��;{KCP�3}��R�cNc� ��EUz���{0��]D�Q�z�Cm��#$;=���A��ؔ��dg�gm�;���#lN�������T�v����6��k�t��/wꍬ��w����}z\8z�O��ŉ�;[����Ѿ����)�w�/���6�G]����{�dl��j�}���깷W鮜��C�駆daY�/�z�;f�����d��c�>ف�;���[5�d��먫A������m�՗f$��k�R�<���ދB��h�ӳa�i�h������To��	U0�C���C���\���N[��ؿ%�57�3��L�ǝ���8UwU�N��SzNТ#�l����͘���T�{�VZ����JyiR9�8�:�W9�`�JG�c��m�M�D�g\�;�C���7WA�}b^����xN^S5���ƪ�@�1=�yy�1��4����t{�+30󱸼���I<�`������g��t�Q���B��eg�DT���4��3�خ�-YO�tǭ�5�'p�y1ӫ�wh7Tw9t����y��>[�\��3D�[R���<޲B�
L��C���#���d�{��ol�n�;hu/}����y\'�oNX��~8����ڔ�S���}�B�{ru��۫�D~�����M��kbn�݋���Y`ڿ]��F�W�숄o���oꯚ {�tƑ�y��K�(}�UvW]�	��s�ߎ/`�x�.3�DI���KU�R�4<��Ov�t����2_���Z�>�_�q�^kTe���������F�4;��g�e��2Í��~�+G�D��qn�ݸjȥ*e}�"�^e�G�����52����^k[���M~�����$���o����?:�D�Tf��*�Y��3b��%<B�b�VG\?��O{o���uQ�BƼ�6.�:�]�t�-�ĝ���=�4�F�q�QG6����^9ѹ�@�3'v^V��w���G/;r�g�|'d��t*���EEhE����Z�n��_+�7���8��v�kI|^a}����S5e�^��'@22N�-�4�u@�Yɽ[q��;՗��#vC��{X�W(k���F�nS�]�̏:���<�_1.�DX���s�M띂K�:��vD���̎��u�Dy�3Ol�㩍�j�yy�;�Q��Yw�q8�Un@�Z�Pz%C� #4��V���w�f���_�V�Q��
п���0Њ)d̜�z/�S9�*�!Iߋ�&��WyZ�L��+��O�=ÕL,^����T�ʌ��P�LxҤ��3�2�����LXMj��I����=��C���Tmk�&�~�=�̭�S���\аwy�)$�	�o�>yz"	M!R��{U}A�~Ν$��5 o�m(*cY<���^�uLoNl��B��Y}�j��S��=~$�o�V�c���%ȹ�r�'=�k����D�\�7�g]�xu{m�1�d��;��Y\�j!��F8딦x����+�9S��$W��-MW�AyP/5h���#��m{=Ǧ�m�jq�W�f|*�����=-eH�}��>7�/�[tM\^�^[����Rg6p>,����?rA�dE�YWU�#����2��YJȩ��I�'��gM��a�R�k�n��M�d��Qı3Pw����^�솺��B���B=b!�ҩ*��#BEO�v�7�i7+i��4�vr�RI�w"�!��%�wp|)cAU,��M�1٣>�ػe�ze�NO�r��C�*צ�_;x�!]���z�K����6�4ܣ��9Q��/�:���l!#�Hg����"��{kܭ�|����َq��~���흥�u�O�Q}驰�w��zca�T7��ؑ�#��V	=�d�yMx�]�Ώ)�w�D*:ҟmږ{M�Z^����/{"VJZ��~~SV�ǽb�膎�z�]��E6}�����}�7z������te����q4j��<^U6��j�tf���Oo/@rz� ��Eo��!���0�a�D��Z�Dk�Q^}�$.�9D쇢V���'�CwS��8��ǆ����ʞl#�������lK���gR�>ܧ�6W�f������ʟ��ܵ�/.f�����G	�ܸ��o��� <�g{���Nm�ѫf{�ƌ��C��w"��+�%�]���'=2ĸ~�����]��
���Nc��\�G:�,�oW����:+Tv8��a��^�dUf����^����lK����?g���mD�����e���ٰ��k���O��&� �W��(�A�Q������;b��55;�S��ˑJU�����aE!/�ٸo�_jRLz��w�~�R/�g��>:
���B}z}ܤ6�H�'͊Un<4�y7B���T��u��t��jӼ/,Q���"\̨�R�5�H 7�����W2���;��g�x�Z(�AG�M�=��+C��O�]0v��k�&�7igp��9s�oXu4Ǯ���Z����Srwt����n��X߂�A�p^��R!]��~�=�z����'EI����{U,��v��㨮���w��عb#�=��՟-]�ʾ��Y	T�v��%������xe��b���x�*W�zw�:-g�W�K܌V���]��������t�yt<��j�4�WpH|j`#�psL)K���wD�Eh�d\�'���E�	�\�(��W����[&s�/W�y-�ߖo
�N��s�m�ud�0^uL��$��(Q,�7&�n����2������RUL"j*:`\O]�{x��VM�t[�<�d�0
��+q*#�����ޑ��4P?W�M�ex˝�Chս���ju��u;�,�yԨ��h�|��R��~�9�R������}��Ee�R��<wM���申��נ�l����;�#֚��{��]�}]ૺw�CѐC���j��"�{N�r� ����i�����G���cP>4��1�r,��X�Ֆh��*��.�"/%���Y���g�yֿ1K�~��,�Ļ}[_)_qޒ��^ϕ�Ak�����ϝZ����֩k��:��D�3R�%��n����d���Z���[��[��=b� 7�a�R`�<W��=�� ��=L�cU�U��]]g�vA��L��m��]�\)\�;*��?��x�qZ�k�h�`�u^�T�Z����ܶ"2�H3�ӮL�Z�}�:���
/|���X��x�`f�;~7��^�kB���2���U�fC0�y0�ҋ���O���a,�눲�M�4 N�o�ζ�䃇�_�c�>�:r�T��:���kЯ�V��bSN����g0��EA�
q�S�=QՑ7=��Q�ˍsCjMv���1�3y%���B4� ���o�S\Q���M-��4��u������=X�:��=^�J�;���M���>��HY�:Jvz+H�.�^�Q��v��8�'j�ٷSY+k��|�ɰb���B��P�RYu��V�=�v9����\��z<^A������]�ǐw2��ʵ���S��/�U�[����7#'���=�˹�7��7���{Ʌ��=�g��G���}�Xٍn,�S���������;�f՚��*b� $)��R8��i�*��`���b'o���	�����N�ɚ������}OJ�Bz1ywZ {'��'��Ǽ.�y�&������X�ch���ԅ�p�v�=^�^�7��Yb5LI�gh��`�m߅�ڠf���n\)5��t�L�H�7f�f�l�j-�W.�V�u�^�G=�Ȥn�a{��ڔ��GQL�YRRT&fa�E����WK��`�`9���5��
Ύ�1��ӏ~ٷ��K��]Q;;K��7s��z���O)��*�㙲o#�=`
�S����;����u�y������흗S�A�Q�gr,�Q�`t�=�վ�D��r7F/8�7�2��P/�HҼ���>x�K:V���zyxXTz�i��s��T��������)���GFFZ�Jr�$�ES�t��-��y��������0�R���F�xɌ�46�Dl�a(a�LvUuhu.r�e��	·�^�����N �P[��Ѧi�3*�D��"���~��H�l�=B�B�ُU32�91�ڍ�&`/>�	ڝËW�`쫌Ҫ��7Ҵ�_p��/�3C9���0f;�9��K��揰�r�O��5�MJ�Ӈo��p��v&�b+���MW����´��ꚩ`@|m���v�)��[7�4Ĩ��3�[��i5ږ��5W$��JE�gUr�^v;A��g����6-�E��ؕe�W s6����#� +޲�1�s|�.<d���#�h+�:��3��A��R�^���Fb��gu���-_Y�O��<��J�}N�.�P�4+�\�i�g���T���Y�/���n��f�$� .s�{�Էq��,wN�Ұ:t�?GJ��e�Y�ɖ����s�����q6z�3Y�ڵeG�Ą�L�n��wV>�2�������ᛊ��N��lwR]�w�0sn�\m�cn.��y���u���P6����o��.�}�{!��|ߔ�}�K��Hl�LX\��U��(��~��ɣ���#3�������s��<+�4)ԯ+�zn$:�"��+9�<o/�M@��*���t�{듦���&4��A��ɫ��&r�No�Sg=i�'61n������˟X�\w���R�@߃���w�Dj��Ny3���챛3�{�'gu��ۂ�����c�׻+�z �:�6�Ay$*��>ɨl�\HB�ݚ:�0����E7�ɣ C{ћ٣D�Ա�����H�q�nv��1̾���o������W��|ƓV6����z��
�E�i����E�g��E�[`^��_ں��]{1�K��ދ-��%�7�o~�eos]��y��i/� m^G̎�ht���2�M�Sv���}����q�]�zz�\�׹�p�^�[��ҳf�X�0�4(^���W�.�Ez�ܪ/#�t�l��wK��8�f�)-���
-{���ëce%X�n�a}{r(_�L�:���ʃ��y�Zw�ׯ��кȪ7�6����C��/im\�*띲�j�a]J:��;��PųKb���^��Bl[�N�24B
��x��f\���ɪj�:v�$V)�Wڷ����	[�����)�}��ݬ|Y��m��05�M���.mL����
�fa�{�y��2Iڲ�Rꃍ�j�^��h�����:��H�)*�;.�&T��Gȗ�3��Y�XY87���#[��vd �1[��
���!x;�/=��Kd��ٗZr;�GRJv����W*7U�;Ν����
2N{�|�R��a�>����^�|���2�:W������$LS-3����x���:���Mo�?1���z�#���g^B����{�I���E�U���
{��v������qxܖΓ�f��gz�X��:!�����)�'lz{=X�r�&EY*��^ܟ��1m��ǐ��8"���2t��،�Ȏ}���ձS{#:��:�<�ǯj�h�;ZoVr�h�/����u�.�c�ۭw+]2�7y>8��(�n����eiҩAF�ݓ>9�=�'�sʕ_�n�]����N�wlŀ{�tu��Z-_���c\xW���9a�=�Q�Ac��t�?:�8\:�^�O�w��dy�_��<e��:l�=��=a�g�gDK�Js=����"�d�<rzj:�]c����5G�����#+��I�AF�ɯv���Rq4%�9�����z�U�|�p�V�G��vom���������}��zg[�f��誸2��{����bN�غGz9j�v�M_fT��X��Ν����wN�iM�+`�X�[�`��*��u�ӈv���8�rĩ\ޛv:�sȄ�MP��2�ua���
݅���j$�0>;�Jeܼ:E��Ӛ�wʋ�U�z���l�Uv➍D���/Ǽ!�F1������or���l�.���0��7�k��Y�����!(��b��U1��{Y
J�5�t]|�l!e<HQ�S{ޛ�7�.�HQ��ֹ�ȯ2�F%P{�@ʝ	^��n�S��7yxx�O��Wi�*ѱrK�2�>�[��o|��(��wvL�2��lzw����V�n��k'����h���虋���1O}s>��v�sC:v���b�ۚ��^�P�ꑛ��F��z��w����;~poƷ�l�c���i���A��+4��5��+�WY׳mAq��W���b���h��EM��ޝUeED�3]�hǺ�Z�l*6?h��n�(��j�z��Bv.d圽w�z7-)ɼ���`��ӑ���U`}Ss�/��=f=Iܟݛ�w�D)�{E	�]U'��)�q>���=�������k|6'�h�C�ޗ�.��t&��Q�����,�.qWf6��m��~R����ў��.��^�>>�=zP�R��_V�O�@:��z5Z���¸:c������V�9���bfgv��}]A�xoZOi�{�z��3���F����]Z�g�ނS�wQj��|�GR��g=�h���y��e ����X�׽ߙ��{��/�k� I I?�II�����@$�$�II� $�$��$�$��	$	'������/����8����o+e|��lK�X��;.e�!f�`��LQ�`Ҕ�K�,B���2�v��L��5NljV��؂���>w"H����iT͛p�c�r�P�搲�FB��	�M�?xʂ���l��,iU��5sf�hî��
fR[�]��6Xeh���p��j��n���OQ����$ɩVZ���n����ޅrU���
oU��FҺ
A��ueL�4ì򽼆�Ӗ=7Z2��i�cuc��Z�mlG-��#��eƬ��*�J���f��ٛ8�m�O&�:
��)��c�g5�t$�#t.G��,�U��5��m�ˎ#w/E���a���+��n�i95�L�QY�M(��;{��A��@V"4c�P^�e�`�{�
S�FI�Um��bDjpX9NF,R�����ٵ��˃6����j[��Rι�mE�Ɏ��tm�榞^���e�WX
�#m!��w��gBE
�F�\�sT6+�����6�MS,�X+3Z��U�L'
l�B�xK:��VFP��
Pf8:��w-�%��4L�oYh��2�Z
ӰqiHU�WI�Z��w`D2���4�F��:�7I@�ǌS;�0ukÛ�|�R��CFۿ�cnĎ��	��:�Z���˺�f�lb[�	\��B)�v��7[e�al�����2ʊ���_�e��b��<r����+�j��Kǹ��M�ڬ�v��jG��X�jR&�j�@V��ͬ�����̪ ����ɒ���[pK0Š�ܨ���1�M�n�+7d��U'm�L�/t�V��j�.�l�s�]��or�<ٺ%D�e7�n�j��,Tĕeߝ�{��f����3$8ݪܦ�⻉-x'����YL,uf;̌TE�G`e�dJ;�p�H�*)���m����^�����j�q~B�)��H�4 ��6pRɴ�^���3M��CIn9y�b1X�p+ъa�Z�9a�`�˅�f ��5X+]�a�Ȇ|^�le"������l�Y��a��l�Rk?�����HB�$	�2I � 	"�`$�@"@!$I! ��	 $D��������$�$��B�a !$?��� $�$�� $�$��$�$� HO�$�$��	$	'��I I?����HO�1AY&SYZ0�(��߀pP��<�� ���pb��  }>|�b�)RJ
����IU��(�*BA�eQ!RE!J���TI(��JJJ��TJ�QH�REO��  P�U$QP�DA"R)ER)(UHH)R��J�� JJ�$T�B(%$*�*�R(E@�      ��$�):$�U�Zid�El�-2�څP�
�Ѫ5E(�c��ҭ�JH���i@V�kD�����:�)R*%TEB�ھ���X��W6ڻ���Cw�4��zu��T[.��e;�[�Ms��]�������[[�����;1��9͑˪R�n�Xb�U�QEB$P��֔��.UU��H��2��a�%����ø��e'Y���hͺ�9���8�8�٭ v���I�cb7 ��]R��%R�AJ%U$IU���@A�Ω�Nκ�]v��n�A�J˵;�mM�Ðs�n�hUT��gMb��uK;� �G8��$�P�wE6�����Q*!B�� �J���Ж�G]�˸������\�ݻeIE7!g]�ꃮ��5�a�f�T�TkB�[��'j�B�Rέ�E*��;�V�Y�꒑J�IH�*@=�[mQ�:Μ� ����KJ�:�eWr�u���r�  :s��J�)&���i���ڜu7U]���*�	�m(�N�Unlm���foy�($TE**��%N{q����n��EU4��t��U�6�%c������J��b�$��Zj٦�*�֊���:�ql�h]V�;���gQ�-m�R��B��TU%T�$�w`�ww-��N��s�f�5���N�bj��G8��u�1[v��F�cA��.u�v�e�5r��ƪ�c.���n�:��[k7X��sTJ�T��UAB�Hw�6մtgF�Y+:�5�)R�uuuk�ű��뱬��C�n�S.��v�7n�[lvVX�N�;
"�[��T���qU
RB��	*�*J�I�u�5��S���v��@j4��Ի.�֌��+��m�t�e�qO^���\��Z7;�m��Kpَ����==�W�mU=)�:Zչ�]ݏJ�6εѤ�ytth   }OAÑ"��&*T�    4 S��$��Q� ��@4 0I@i������#���S�mM �S�A)RH      "�ѣSj�� �@h�$@%Q@ښ��d��hɣ�2=M��_��ȫJUd��Q�#�333����{B�9��1�v��Lo�����EVk������鉱AU(DQU��Z�����ە?� QU��r��
*���TQEW�b���D_�E*	��n�b-A�@�jT
��Pq��
���������D[���PIQ.  B�
( D�"QB⢅AEAQj 5j"�V���� �B�!QT� ȋ � ����B�"T j()��Q� � j�QB���j"��(��[�)QV��T��AJ�5�A*�
��E*��%�V�7* �Q��*"	QZ�#PZ��P��Q?�K�f�%EAR�TFFD��@*\S�㈩��1��Qn5����K�D�����������t�;13�lNM�~�am�i�r:�����k���P�2�ss9.�M�P��r�F�w���tý�Gb��Y������|�%ΌF��O��&��y�i=�JY�y�h�eݳ����Mm&æU��g@\�����:u��ݷKh�ւwi#����7�gd�zɞI��Y���42ʡ5�n"
�����P��*IFX���$�������Hći�3�K�#������v)ȅA..�ȗ�NX��j)���j)q!��w7 �SqM Ȓg&���b�\D;���2!�%A$C�J��!����j	�&❈v	#�g�8g|�{�W���-�t�7@�KQ�+=[��)�]8 �DTm�4��M�=�K��5X�`�c�n�t�c�1L�'m��1�mk-fN�[�F�Z�uB�^�K��������˄>ra�]�c�K�m�WR�aY�'ZݮƂ�MSS�1�d�'wK�y9�:=���g
�Ϋ;5ʳ�+��e����-g\OZ���ėI��`F�N}��]�j�>�\���R�WIv�z7)��70��(�H&�si<�*ӷ�)��*�[P���6fNU���iu��4�9vv��p���Q�qm$�0� X�r���h��&�VVfS
�d'�C�֌��z�lj���	>n�9J���h�F�
nxV����Z1mLTun�����&Rl��x�T��Z���rL��n�(Gka{țX3�EBf3H��$2��,��eh.�܌ S��^���z_�������]]���i̺4 �Ǡ*��nKj�'���76��J���MC
�i�p��)C+4�P����@���9V�Ҋ�c^å[��pT��%�X��؞�+t�A&fBE��`h��A�@��Gu`��5�3Ko,�L�T�;(K�H�3&�\���
�(PxO�~��rr���m�B�\����tX�W_�Sj��;q�/��n�CE�I!{o�Ȧ�EH��[��G)c:�qZ��+��-:�
��ÚL�KtzY�F��v�B���,f� ��4��Ml��,`L@2���R��~;2�'@�#����bq7�^m�n�&��	tp �]��M���އ��-I�52�b�F�*VKz��G[���f7r�E�u!id�\��'pIN�/��HP�L7b��ol�,՗[$]2�pѶ*()ۂjZ8S��}�]ݘ����;z�*a`$v��j�Vl��S(J��bm�y�����@m٩R�Q�Au5[	Շ2�H�ǅ�^� �ne���w+u{B��2��@�N՚�^�MϬ��@�%�Q�X��U��^�r_�h���
�5QO 3#���%1�Vh�.��h��-�)\L�ڶ�eǴ�@X�m�\�X��Z���*�wfn$c� ��0A�A۩M�V��?�*�u��n,�����Qeǉ���:��4nVJ#]6៞�n��VU&��P͹��-���*��i���������1L]��f(��zEd���WtЭ�[`������n�J�<[�SH�eK2<ɏ.�F�5w�Fɬ�l��ŶeJ2�[�Q����1<���C#o����Q�
��b�rY�bҬ�xc9�V�V�8ݽ�Lӱ�b]�H]�LƬ�C�h0Uf奊�5�@�U���>��M�t�e�R�nT��aJ
9��K��]��ֲ�PŤ<N�VPM�+m٫j���<�9K(f�$Tkh�Z1�Lb�U���#DX�T-�Y��3Pw�J�`ӳX(�[ձX1�b�;�Y��<�v� V����	�}X+ꂴ}Wf�,���n9�Q��mv����.�)�u`��F�<��=`�w�4�GX/�neg\0��T��#1�]�_`�������ۮa��f�1!2��j���jY�M����2v�k2p�i��Vk��E��E^�Xe�=Q�l^~b���%�@n,cl:�M�)��J;y0�X��M�K%+��l66��)��\��ɷ�@55����yIVɨ�,f��J�2��K�:�8�ض�RiX�j��Y6��ak�H��لMZV lY����:�nZ�).�@PE
���4�h��lnV����L�јԣ���/
�D	�B��Y���I��������Ҭ���ng�\x�7�i�[zNޔ�J��W@�R۫v�O&DM�seN�OI	�ɕ���(KGE
�H���o^���W*���@RWp�mdicӢ�"��M�0Q�y����9F�����l"�8��Y��Mٸ�w��XԢw��f^��/���1����*`H�U�c��eǆIbvlِ!Y[�*z�ae�h��3H�x,;�"V���d��^uRv]p���e��b:���f��)O`��Xx#�cr�ٔ���ۓ�W41�l!]2�Svh�]nb��mfc8�Ŵ��3V �QY��<�ZI��.�[ʊ��n6�nC��6��8s2D����ѧ����`EH�(J�.ZJ�V/�2�b'W2��3*���J�9B�ࡈ��Ȥksr�����Z���=�^�AT��%��LH�ۚqҹ��?������d�f�&�Koz�/��t�7��9����&`��T�/�LLJ���PsX���\9�9Չ�Tw��W�Gs�]�O�X�p������q�h��R�{$6���Cޅ������*����i��t&m�$л�=�h���*���|��)��w���t_*'-�U�r�N4�V�1v����+s�LdJ�qb.��XU-*�-e�RU���| GG0P��>K������c�����ͬ��o��ٻ{BJ%c}.G]�ܶ벮�WX]��7�`�n�l����Ν'`��^J����A
��H�z�N�cok���먮�I�p�%� 6�r�dЀ�Faq���^J����gmb)�v9��9ǣu�]]��u�@���F�c�[ec*(�f�"���&X[k7NQ�1b>z��53i�e`L�2��Up�N��t�Vbl��{�]J�(���sU�C���!V�0��d-5��c]fVVb��� �c��'\��a�g��+M�<�AM7�4�b�mYx۷���Cܚڒ�/M
�h��i��E�ݐ3QXF�%���7bܥ�� �� �V�ص��^= K���6�x�%�-�؄���W�.̭�̆�ʳ��r1`��D͍Q�O&�8�P(�*�a���RJx�㙦���'��K.�-Q�̌��R��l����4%��i@X�'���gus��M�Bu�3.�����F�%�0kɺ���0�u6c�3A����v�=���J���U��ǘpV�:N��J��&�������q<�T�;�!#�p�9�+W@V�]�wx�)w�o�ӗ��2K¾I�W�Vi�͈�2�5u�%�5�[��{R_ڄ� ���G1���3��p��5�^�[��!�k���|��x(]u]���eT��䦌8�&���J���ǘ ���^*}e�@
�n)�^<˿ݪ*Q��֖om4�Y�J���aޖ3,Ht���*���;���U�[ъ�.�[��z
��7�-.�m�6�6�[
P�+�wz�^Cz�q���E�n��x��(�y�9�;���͢]�V�h���ȮU���,��x0)������VhӔַ �r^�ܸ�l�Ӧsl���#Ý�{8g\�nbF��RNT�2����xJ����w���n�2~%�e#{,?n̷Y�a���@�-��l�{
�!�4�������I&*�d�U�ƢH�T�^�r�rX1�"�!��~�>����A�j%�{���ۼэboa*�N��SWu�YX�VS[������%�f�vov�Y�
S)Ln�7�X�@���_�}�K}�Ƕ��9i��B3/R�x��ߌ̸�S��4�b��J�IRʖ��^���(�h[X��Tݯ�@*70�b;u�U��v��g���4#��}����#���u�(�̈&�V�[ǌ���S$���twVw��5�"լ� ����P�+]�{�n�6��o/�%Z�����^�m�KX��	gt�/uw�O�ԏN�d��&�w������
������جH��MLq�H�x9RxC��!��b"�.V�I86��q�ZZ�4ݲ(�u��kB^�y�lVfk޷xK��9�
�"c��V�-�(6�'#<Gs��9�o��qAݕ�Ii�G��`e���*P;����᫵m�H@��4�WW���D��K%�poE��ۂ�f�B�����a��$�&����n�Y
4t[�rC����K%+D[2��[���[�R�G���vܷW��@�.� ��*�%Cz�!%���/d2+{M���m�+t��	�m]e=�e�(�q�يD[�z�'N[ubΊ@䁇w�g@�goN��n�/r�ړ-U��Nc����JBfGO[WVi��
m�N��0��d;�7)'�#N��^�f�苵A���� (��������+�ݴmdSk#� ~k.Ji�c
�YK����c6Z������uj�F�A�w
�79�4_H[��Y����(����Ǧ�ͻݡYl[��T�֤*ʐ&W>����>*���,�c�9��u�b�b��@������khJG��@+/ �F�G��XR���/��ׂb�%�1��]�rE3PI@� �3r�UicU����\�6����cn츃�W�^&�f*yB�*�op9F�1.�zEiJMA��X��N�U�u��Q��hG����h���E�cBJ�f"���-�u���Yp;=���49#�n�ᮄ*Ӕ59Q�չiڽK5UиԳ��ӭ���-0���,��]' �U(l��Zt���U�#T�|�spYS�W
��}X�����P�k��q�?u��t8�o��
���#�m��e�f�T�]��{�R�7u�!�RRᛁ�t����me�P��ac�S�d�n�f��S":�d�g�\����),�Ne�n��5�В��ºQ�6�x>����#���=|�E[}�s�*&�]z�S$-8��'p�k!��ʷSW��Ƹ�q=�1]�%k�{$�S=]�͇���[8��o�ǯWGՇ�ɡ<�����t�N)��:�p����ؠ\U�0��֐��3���A>�j�%Jμ�1e5jkmRK��&���yH^~���3����nu�J��:)tU&b][Mr�*����D���j�e7�1奥q�j��j��C��nZF�|�dQP|��Wm<�j�rR�`�&���� u1�GU�q���+{#�{u���l������6�6qU�Em:����d]���މ*�U����B��o�(� �ڥS.ޜ�a��Tt���j�,nj�g�NG$e��n�XI�@���u�c��6(Һ�wm�R����*Wp�$��
�I��u��	[a��,{-�Yej�vrm��I�(:��}���F�-=�]��4`�@1���juvZ���z�@Tk V�A� ����سhG������_����[J�2�"�n��#8&ټ���Cu+��Q� ���n7Zѫ��X��d1�"�̳grX�S���S�L���d�nB4sPb�&���U�R�o��e��jUӬ���Vat-�y4T�1[Z��!0㘐�a7C1�rQY�n����ōRnR�C�n�n� ��b�7���{o��(vՆze-OF���m�udאPF�7F6�mhE�i2l�X�-Q.���a>¢NU��(S��ؙ�T�dP�9n��x�tÀQRQyH�%��ӷ��]�ne�M%{����=vqٳq;��%��e�����ك^ǙN�fmD�U�\ͳ|��|���{na� x���mi�d��eȯ���-�����CV�^�)4�V��܌t�B6��7<�f��WLtʙ{&
X��+bp�eE���_�94�ގ�jZ���42�<L��K�i"��l�u�7 �f�*l�+Ppw­'U{���M���,Ihm�z&m�l}��3P�9�����٭�B��Q���E`;B�ӧH�;]�쌊�e:�ݖ�"��/n�;�R��k������[+�䥖LF�D��2α�/mQj开R��7�e̺���I����T�:*��'����u��{Ę,+��d,:��L�Y��CKh�[�#����a��ۨ�ei���[��f���`7����^Ʊ��wA�
�e9-YL��ۨp:�j�͢��`3m��p���ҶF��ݤ	�ML9���/+MB�z���;�E���nӡ���(D�۳�?	B��]�Y�J3zA�h-SsV+'��c�9���;mm����N�	�/]f`V�Ķ�A�
cF��+KVq<NP�Y>Tg�ow$��ҁL�Z�aw[i����4���*�ŭ���Z�bXЇ#���0y�$Ď:utn�uk�j�ӽyoyd'qrwP��c� .�Z���Dm�}ٳ! IV�ሺ�)f�d�s94wT+cHJ���4!S2슑��R��3Z�d�r�XO���c�?n�^_=r��c#�m�L�� �y�X�4ѳug�G�fr7�m�)m���Z���s�^� �(��̫�@� �Xʮ����դ����V�*��;�iC:�=z��;��ɝ?t�ˏ)�{�������\��]���,�ep�8�]Ǣ&�jEaQ�bU�y�4E
R�I��v���k=������j?����B�_�o�_~�➊>tw5�M�$�)�% �EN|�Uk�]޷���z��L��ﻖ<36\��l���Iѹ#}$�����7�F�H�I#�$�wwI$�����G�H�I�#}$�����7�F�H�I#�$o����7�I:II#}$o������G�H�I�#}$�����7�������I7{���ԁrdKX��]�u��9*X�����F>.ntԹ�]�ͬU��&�[����W!�xj�D�F��&�tr��ʸ���
�r$k��I:Sf�>�/t�99>���N�Ϻ�����]'��T�ܕ-,�Q���K��t��k�N��i�����]9tK�siո�gr-��܆J&n���=����vq��}$o����>��ͽ�SV���F�}#iM�ǻ�j�]�0�r>l����Km�}.��=��#|%%�!<仒N��ڱ�NtmoQ%����M;��w�[�[�m��yۻ��;��e��״qj�4-f��̱�&ɯz�&�Z݌�&L���3�yZ:����Ҽ��`��+ZM�v�����cFNWN�S�ɽ���縐>���z���4G��n�	��r����p$7J!B�MlV��t�(Ϯ����n�aV���7\������L<�4�����쨙���H2�NW]�}Ve衣���Gj=|�����{y�;������1���9��-0e�i�ZS�r.�9M,֬>P��l��v>�_�D�|P��i��w�/:��1#w�ɷyS���c""ʺ�d�Opl�f�e!��!l����3�2�orCY?��]�M���;7^�kέ69e�"���Kr�N�R�����+(�]�.ꬦ1�I��E+�*p)�!��Q��� �q�Xn ��x���/��G���.��l����X�ʈQ���]��ϝ�>�E��V^�F)��p<fϕ�#�U-q\4͚}CvД����MΔ��y�m�g�|5���9��RW2��Z���ud��Ac*�)Z�$��g��ȷ)�{���S���V�c
���c�;{KѨ=� ���z���ؕ�M�ϗS�cՏ/(��2ͽgf�9T]Y��i��*��[3�N�6��|�O;��=,��+v��E`K_-ӻ�˛\�(���6y<� a�%h�vr�𦍬Dm�V�1/�WjN�>������xU�[��j���@�x��v�
f���j "j�YMTV��\����[����)�x��r<�e�m����d�3��k�Q�(ss�'��ee��[�.�gi7yϻ��,���E	NʮkS��3tMq&�,��0ї?f�b�����{N�M��qU��1Q�0��u�6�@���jF�֡����{]i�Lm�o�W�+R�ެE��n�G����`��#��\̙�G��AI��In�+ ��p}8!Y��.�� �J��.\���=ь�y32��;9.�gzC6�7���-��i���d�p�X������9��#]w\�ms�byB=��{����@'�;�ݷڟr-���L���,�Y�z	��Ъ#�u4,k�
]f�!ؿ����vh��AMe�Ō!�u	�Ja��'�H���l�ݗ��j��Z�۔Y.�*��c6���]c���Xq�r�1��Z�v�4�L��y���֔7�oU��)��w�{� l�Bc��y��s�EeǬcg]��r�v��M��S�W&ꁪZ3��Ԃ��_1ba�|{�k�������x�!��C#7��أ�]�������/uculebln �.��"����n�=֯D��V����#��� �\d*�X��2�#U]&�H�J�|��D��֔��WU�ֻ�������	��:_�0��x��ܧ����͢�p+�%��5��3���7u]�Cm��B"��S�C��(�����x2�j,��7�[�9ž�H�p�{��+`��;�H[΂^�tnR�//9�c8�9µ}��i��û��	G�ɼ!�ѭX�<��۲�c/W'+�� �V^�m�r�YRf�74
�5�#��.jZ̛��gj���|۩ԡ]�ЛCP��	��;ړGA����XX©[�4uf�+,�L/B��mX��*Ճ7�comB��ˀ�p�k���+E7t�kF벹h��O��`�1!F���d��7��uJ�0 Ju�nI�nCJ�K���W����R�5�]��H�0�`�8��6n�Juã˛Fa�W�nY�Ki���]���N�%�L�+:D�¹�I����-�x��V���A�g�j�r��O^K�r�WwW:�ہF�1�T�͉�7��GfC�]:׎��v��GFY,�IWmX�$<:ʻ��T�s��.w+��Q�/��(�Æ�����}�_uE�d��f���^�ޭS��R>������G�%����2Y�G(*���;.�wY�V7#Z�x�F8�Rrum��<�]��&rU�Ete��ԟH�<Ց�˜�D��]/���t�!�sD�g�sO�/pf�t�d�vL�@�2��V���ِ@nC��rwR[���L`�Gh�:��hպ�<�;��[Y*��N���X�)Q�(�O^ˣ�U�)��� �����N1s�R+?H��.���Y�����ُs�w֧�Rك9W�g�$�X:�L��I��uśt+��J�<{-���Ma	Ӭ�v�=U�bt[#�otX��v�"�m��Jy{�z��V��c�̙�,sc���P��R�5*WC��3��,K�H{V^NV�T�ߧJ�~%��#2��*h�|����ɔ�կ��I�δ��g�)y	Ǎ��j���b�A�)ۇ�>�ݛ����h6�qpah�9�Q�-w�����]�Ł��=�k!g8Ų�eb6��ݮ�Kr�%���"�9�,��2�*j���t� 5ͫ�e ���Mc��F��y�|5�yC�j��2�E��E���c9����]'�yJM�(p�m�.��¯{����A�Q��u=��+Y[g+�ӻtW\���G �u�Nvw[�q�=��꛶6Z���g,B���~��{��P�E�.�R��̸K�y�m^��z�uk���=��n�Rɂ��v���¶��	������>|]�����e̢�F	p�$�1���7x���W�5eoCK�[��Y\'r�6�u�YfH���!,�P��F���p-�y���Y���I�˟-Ṟ���L�-�Vb�^-s�;]c�A}ۄIa�GB�s��ǩ����֝��2�s�kyG����;�`�x��+i�v�i9һi�*,�(���d@d��M!�[���x�v3�3�!ٝy�F
kS�A|gr��U�(tI�޵C�:Yv�f,V:u�Z�4��<��E͎���*3��fV��r�Wv����f�[�ư�-���;�]*�3�崚Ȇ��ci������W)�L�█��� νk�͕p�5�wl�7I�[;=Ȑ&�T��	�3'C���c85��Kx��t�Ȱ҉Lk%nJ"�n�����uwcF���h+H�W�p&ѵ[Lwu���*�e	G�w/�7�$�J����#�g�d�捒V��72��<�8�H���9���S6GC���((���C�,v���+fh�:�[&�q�-0�[��9B���d
W}�I�Lg�[��f4�-��
�l'�zH������B����q�wj6�2.Ƨve���Z�ײ�j�G�o����ۖ87�R|A�U��`{����.;݂�2U����0ڳH����W`�G�7���v�C6l��ITB�+��WgZ{Ղw>�8l���ӯ5bA�{:ô��(\�Wv��9+q)0ﶪ�͙,Q�Y�*pkd�s��pQG{��v�%�me7�O�Ir^nL�Ҽ:����9�ϖ�5�r�D��`���'d�v�F���ӱ��� uB{iR�KԺ���������%��Q>Ok�V�THd|��G ��ط�P���ƭ��o�t}B�b�pSst�aq뾇y
�.�03���|4V5�tY�����	�d|�Z�O'>��|+j���%��4�1+B�$���Ze�݌�nU��wj�:��"���h6,�����`�5���&�Z.�Vd�x]lu�]�Ci.b�����V�}z�*�2�|Ry:+i_M�1ʽ�����p�!5�3��r51Vv����q�uM]��%<��@֟�7�}�gڑs1�c(QG�7$��ʖ,M�%�[��y#.�]�lrNw���}���V`��
�{+#��s����^U��j7	�,���A���ySZr�,�GL��(*CӢ�<�FC�gN��O��6rnQlb��w�w�Զ飜��p�o/$wʍ���9?,yի*)�"j.�֙��849���Ʊs��n�F(>Dv=�pг'M�ڋ1�������8��&7�|�qC�3g�/��FȻt�w������X�2�4�ac��J���͝����G��
��� ��ic(��
� ���ۥ~��N�zAz��;U�L�Ә��pmm�W���;�v�6�wlKlv+�����5wE9J��G5h�)�l�tm�"��]g~]}��Hh��,Xe,P�
1)ݎ�D�[�߰rMtYo�EH"8��4�����4�9Y�$�Zl�@v�=�)��������%���HmκK�c��e�����j�W�RDbF.��=mf�6�th�;OJ�F��+'K�@uј�*�\��"�n�Mw���;��~�־Ĝ���8Ɲ�,p:o+:�v�GxY����imGP�����G���%�'��ё�@��8u+����}��9���K{�7�`U8�.9��gr�ŋ��'t�9�Z�2�:R�+$jcMe�2�ޣe]��ɫ:U�*ζ�k�;-�4���%4�s���+��i�Q$�Y��ݛQ^6� ���&jZ{�}�sD&��&h���%kA�qV�O^���LCd��;�ee-n�2��D)k�l�<c[\�ܫ��ARN����4����zU����ξ��J&Z7u�Q\���k�ЦN��W�d�`�}�h�u���n����W%Ά���^�����&��z7��	ChQ��Z�n���n�է^��X��
��-wY��,�u�K���ھ�#�"�fEp�f�ۼ����V�_[Ƒ̛[4�h���@#m	�gH�e�G]em1�fX�D�K��}�Ii���&w;{*�\A��&���뙵�5�E�Wb�u�Q���b�s��jջW��E蜻pm�:�Ɔ&=:�s���e��%a�w�`�B��t��.���Y�;;M��+cMRN��+ ��f�c�i��~�b�7�n72b]A������>��[:̠b�gcZ�M�3^QUr,`-��YZ�/��K8^
FޔfNױ��|iЭ�QU����}L��C��w�S��� R�~�����̺����Z���:�`fyVw��v.qX὆@p��"�x��,b�W�����)�Y��ۖ�]���r]z�~TEh����cNAk�e's��������)G��G��EA��n�mL����H�Pp��f�X���ׯ�ͩ7��|e��T��\�u��)c���ݸ�t�cƫ�Ɗ��ܶP�wV����җo]dI�j�{�V;�0�R������$�	K;�����o^@��ai\W��� t�7��n�����kꝼ�ٍ�0�|�GC[CrZ��,��9�D;��)fG۞��
F{0]y�+�ز9t��PkIf��`���HS��Q�V
�{\�';��{Jd�
��:��3z�m�`�Y2U���)�ˡW7�LD�Oeh����3�e��L�\�I7����mY����L��}��ObD�]���	�r����bv�Ƈwm536-]�5��+z.�e�}5c\1U�J4��S��oH�,�е9��/:g
v��g���%��e�Vl�'Bl�۬�%��;"�n���3��m�[����A����V:��Ӹ���F�G�K����\�l[��5?u�κ�G+�tF�����u�e ���R��B:9�MԣN�Zy*��ı�����Xtl����4VVw&��=x�P:]7���8C���Y�W�\u��i���ف�B�f^WAh�9��J��]x��Y�dV���w�AV^�5
 �ԕ@��z;M���Z�j魚<�9�cv6f_+�r�c?aC�k�ߞ��	�0��m���Ƚv��,a�]�@5���rT
��<�z����mc][2�j�A�~m�o��#��˫U|�jǙ��A�h�@��t��s۩��hӸ����K�.�ۖ�w�Ry�L;/�Kʳ�^�sOrb�����۰0����p�3���2��-	wè]��H#���4i��=��L���%�v�H�(��")7Pۃ,6j�"��\N131��ű#ڊU�ũ�(e��:Y��H� ,X��jr��n��p9�c"a��f�j�&3Q��uYr�ӗ����g7�ֲ(��T��E3o/q!:�����Q�Z�*_Sl��b#�7 �^s�E�당ґev��e�k����' hj��OZx��K�*�&/iز�Y��`�_��otwd��=}��%R���U,�fs�����ysj	(Q���s�F�r�\�Ӥ�`�ұ�M*C׬C+��E�{l���k�Q��˛7��%�5�[�kfc��� �FX� ��S*򞊕	��-S��fv]�����K�8�Fl7��������[��zʠ0e8͓d�2-�0�"DpV�]�6rÑwL��L�v���ϥ���|bÖB�{se;�k<�h�Ʌy#�;B�=��9`ݘ]cw~k,faa���y}̤n��{$��U:��A9��ѯFj���
r��}�v��zRt�{��"8�7����޹`���4���ʝ��jG�N=n�T�W��ѻ���r0�!X�����t�[��kkR�9����&L�:Z×�v�o[=�sx�>*��o��tfr�Kkt!����8�Ś��}�f��J�}�@��z�u��t;���R�+5޳5�T{��x�4f��˅�c�o�2V��ΦgyZ�L^�5��ޢ�*���*�߬�@@ȡ4CQ�J�G�����Qj ^)@EI�@dL�*!�U����7Ũ�1Bf8�"fb%�dL�$FB�p���$���3K�b��Pn+���CCBE�V�R����*�E���qj v\�I1pI��b(�WI��D���X2%DL��1d��@�[�8��� �b �$
��aQRWPD���1.$�� ��BD1F��� ���������H�"�Tu��0�@K�-Au.ȭFE@91����� !�Ȉ��	 $I1b��b�]DQ�������G0[�ȡ��Q�	 ��&�r,�����b���(.@n*�";�%��@���@����\L@
���NDq�D��5
������5�P�FA�1B��9b=�E3 $�2
�.�b-��K�K��T��*.b�P�5$�SSP$s�WSqB�7n�W\U+#���NĨ�rD�N�D;��$ơ ��H�pA����PA@�
�QdR��"75�U�A�D���.�����4:�	Dj ��n"�
��d3�����""�$qA����.$��pP�1�qZ"T��(M�q�f��$�ؕ�*
f#��P�G1Q3D�1
��A�F@j)p$�����#pj!Ȇa a�!��@1 ��D�@� �pR���2�@��#"����(rEA�S0S1
�����ɘ�j �"\u.)���&cp@� 1I�T�R����b
\Pu7� 90MACp��K�]��b"��	�+p	�U7�E�7Q5�)7MA �@�j	"�\��"�p1 �J�"&`�](�	�*ESn ��
� ����ED��_�PUO�~���������i����|b���q��fl�F��fo����ގ�I%I�*&�U�l��yM�����ܼdL5λ1�Xӷ�X�(�c���*E(v#�p�L�Q�NT��5[s����L�i��A݉x�-!�6���ݽ�Q��A����R)V-.�VgbT(�K[T���R�o,��
ڕ��A��r��:���]�jk�O��zg���i��f�s=�A�}Ɛ���+��S���ݚ�I��ݝ�]�bzcӏ���P)8{M=��-)���8���;�cXG�eFF��ʺ�S�n	mO� ��Mk���;kp
����eb�b����̎�+��j�����IZ��x��Fb�SF���}���+]u��L��o<:)�G��6�7����9��A�o\���᫳yZ�\٣�\U�)#Yu�ocFS�WN��u���k��a��i�Ц(���f0���M�[.��
;�+����b�������y�W%�l�]�"�j�j:�tE��8�6�~���yc���n��IW~�6s���&�&gFX�3�D�R��4ҍv��eY�ב.���S�HOq=�Li�'�`K��;{K0f�i"@pEy�o;���w�ݶ��eŴS�UF�L#��htW>q�a�Iմf1ul�j��YO��S�e�B`��:�aO�SӮ�j���0�;c�W�`���,����{s%Yn���(��1��7'��F}��Gw7�Wm��К�t�5�/5���NWD�8Z�{.C�I#��B���5ӷw���݈�+��e��ڎ�?�MkjOn|�-��Wk6l�V��εߎ]04��yiĮ##0i���c�{�u~���B�$���ػyʕrm ���t����J��)Vx63<>Б~�ˣ�����3�b��ܥ��qȌ>@[���g{��}�̚�-W{W��K܍�R��M?F�X+��2�qኸ���w�V�=�jo:�<¬�Y��vv���M���S�E��vH|u���Z�|F��_�ě���Թ��L���Ez�a�.Ĩo���=J=��7ԭ.S�����ǊrqmxN��^���Q�[�LG<y�;�pא>�_�Y�m��"�9RJ�;�({���.���aS�=4g�������6�8W�o��Q�� ���d{G2�^X��Y8c]����+�E��׷�Y��p,ǵҌD�|NR!6��g"ŋ�>"ǥm�$Xk,',�>��X��%�+�[hى������sWG+fI`���nq�GW���O���Ky�9\�ʭ�A�V/����I�X�5(�����κ:4��k�	D���Qa�*hYƹ�׳~Z1;֨�ף�����vυ�lή>��Ko�����A������ҬXݍ���x-n���:���[t^װ�/m��'w*Sى]�_S��.���k>U�{��M Y��=�M�I|���[�?{��S�L��%��.˵'k�^�y�ޑ�����+�g6�G�3#u#�>/%�;%-�*�~�JWe9Q�M����c��{�`����<�+�i��}��<7ݻ)���Y݃�鞿t�ý�ڷ1X��	����%�Ѷ����◍��^���K�k����v-M���r�ڇ�ߖ���q陿�)�U�8Q��BU�{�B�Jy��:�K�/ڧz�.Ͳ||P�I���i��{n�V3�|�~T�Otu�o&��߇�}-e&J*ǽ��D�<��ì��Ѡ��x(^իK/�^D���C���w��;�Ǭv�r`��#8�U��f��h./1�ۑ��}x��Џ��+��s��ef��v����1)�<4���+�D	�OQs�P���`�L�s�,���.wr��<"��_n��
x�/�n�E��(C?fX�u��*31!Ő� ���|�g�;<E�p��'����ʇ�Ss�/���j/`gI����� ���#��o��#��7bp7�.,���=���<�n_�fF�s�݇�Y�=hзp��
>�X7Ow�H��\u����v�a��������bU.�3����)nQ����	�(
��g��e�bj��=}��^�����x.�-V1���猙�V�Yu���^�x�r\ֲ�q����=~��8&���������g۱�������L��g� ɍ��������ƾ�(4�==�{��#���x��.�r���]�,��o>���zCiWx���;u�&�6�W�S�*(fߥ�7{�yikǵ�To�o#/6�rˮm�)�	�YY�s�I���R���
쐋�r�W^�d�P�kFy��s�[��q�Ok�ijoy�B��V��e�`�ne(�5�*�X���v8��!p��ؗJk�f��&'�H=�t�F���pZz��I.z'^�&ȩ��"��e] T�d�u��.n�L͢��"IE���4r�vZơ���,̣��(Ĥ��%�K�!���w{vaNo�ss{�S�u{�[�=�z��%6�R��T��q��3Ʉ�;�^���D���^#{��߳\|�9Sg�5p��[���1mo[w�\�
��5b�z��?���ƻ�z`BmG��#:��!hT��q�M���]}����� �u'�>^���^ꓳ��̹$���h:1�������؂�>S�<v�8p���!
o2�Y�׾���h �-�Վ�S�u��}��ű{������"nE�������y[��{ʻ2!"��⎰��7��CG�t3��N�}D�D�x.��Y���c����ꝷ�.���t��u�\�Gπ*���V�����/|u2���A̅�+6�JD'{F'��5im�	Wv{&,�M��΂t)[�^��|����ˌQ<�v���k��w�V�ir�}w�z�M�|k6���if3}�C � ��SE�X�D��m�ٖ2��嬚ku-�F'R�x6޳������y�4��(7 �m=�\iY�l�.̥YX?N)�Nw,n3ͧ ;�wn�P<�e�x`=y�h�o�^n��P�
7b����R9���ys�5|`W\0�F͹nP�@щ{)\u�C{�M�f���dFLx�?tq����<��Z��Y�j��xb�\q���T��"���C&5-��M9qy�{=y.���x����y�,��؏��_ �"�{%^��rٝ��R�B��7-Ԧ}���E]9��ˆU��^�4�T]��3Kۢ��z���b�֒��P<U����]�!�����߅)R�@��n�*�ׇS�%zi~����cS�/J��Li��`�^�:dPLk7A8�򷉍/��_(��-s�~��5�+�M�< ])������(q���gjur�1���Ś�s�^�Ѕ�[��/�����7��G����a�b�T��+���?e�T�\�nݽOM�۴.��^�Av-�L_>8��s|9x2�h��X�Gs��-e,Ŵp-���l��V��Ph��S�R6{{�i�Vp��Nr�Z]��vyNj�j	�֏���X+y8�l@�Ո+�8�8Yسl4����ir���J衍5y�Nsŋ
��[2qW����8���B=�j���l�*�m�t��_�\s�	SS�|v�<�2��]v;z޿�R	��0�����&xi�-�ٻlm4�)2��1�
��ԧ�O����°ߒ�s���٨.�v>Y
�B�W�^Od��Ӓ�+#H���탡׾��<��$�,��{�q�H���+�����YV���ݽ�G��	����J�j�7��K6����Y���vlYG��[!%��*�K�]+>�g/,T�����Ú�0�����L�����5��	/��}u�C�Aܚ������C��k��mt�d���^�>�Q�9*���~�W���!^f�Vj�P��#	u�#��ږ��ӑ~9+ϑ�F�Ҟ$7f�3��f������㈵}�b�y����H����k/�^�^�~��+��,`����^"��k,��;�W�E���ᓣ�^��P{1d�M�=H��EV;VO�E�P�|ԭcy�[���W~�	
�Y�Vrd-���&�gwHˏ��).�{\1���_Ǎ`��u�dx�t��vJ����X�o��ug73�����|ޞ3�-]B�IO���i!6�e�c.W�ڱ�c�}�Ѯ�_p�-�kl���ޱ��|����&Җ�,X�e�M�iˌ�|�\_�=���	���=�y��u�[�9:��
�
����E�Ů���9^�Y�m���k�������
�+�1Vq^A�v�V�^�B��4 w�=R��1�0hYd�kH���t��C��ܲ�����ׇ�vյP��K���üW�35Sgxps�"�Z\?�����먽B����Ǵ	�+s"�f�-���e�3��|��.�8]�:[�3��N��k�e�{���	��=|̼d)%(�?h�K�w����=�k��<|���u��7��j���Np��Ǎf���6��W�T,_��y<�v%�K���{4�îl�m��_����߯y
:����>��]�B�FP�Zq��]�I�3�<�x��VC+8nN����=M���������7Fw�U�V}:>�7��G��*dm#�خ7{�{7�G���<6N][3��KaJ�:R�H�J�b7\���(m�a�RQ�^�ԩn΢��mrMv�{�t��|-�,��RB�U����ƍ� Tv�_;��8��}���}&�b�{�hA���>v��o��YL}=����������؊�w��z؃|,�/:��g��D�ު�:PY��Ҧ^��������w} N����~�Ȼ��lAI
��C$&wtޗ�T����	^8)&�og"wўKcgv7dB�j*�	ܺ�{&N�ڟ%Suu�SK�b���u{|=��(ssۥ{R�(%�?Y�<���:rs�t�LAu����.�o�.+<��/k� ��É���G�}�����^��0��S�����縦�dX�y�C�ؼ�MON
�{�'&��_�nL
�,qg���Q��0��:�k��Z�	�3��\�We��@mh}gu`ޚ��V��^e��֬vrMu�n�8�:W�J���w�5>��?��a@�8\Ek�����޳�؎K4�}ؒ5Ǐ��I�u�fRx�y��qݾ����~�k�+Å|U�h�/R96N���&�؉��*�M��u}��B���y8�ۻ��2΁���:�\!R�ʎ��GU�5��ɥE�I���{�K]�~���І�e��%��Õ�,��ʶ�j�wL䃂ݍ!�l#�&s�q�O����W��B�rfE^~����:m�|*z����#��l�oy���2�]<��΢�T����Β8����oV����"���u�lŊ3���$e�hN�L��̹4�dГ��=u�=ՙ��ٻ��6o:}I�։��y�Ubǽ]d����^���s�^���X{����О�D�I�O{o��w�|��Z��w�0��w[�����Uk��wL* 1��<���Җ*�#��~�k�뽋ۺ�	><���Y�Z���s|��=u�יW����
5��̧^@A��yF����T:;M}-��`]��v�W5X���ad;�����ѻ��D��u`mj`����ͮH{ބOo��2�yJ�h�C���}8R�N�Q����B_������htU\�dcN�wjJ�OC�P�.��c�u�l��أ3ܽ��xj	�N�R�ZWH{�u�T����%3�%A[OV:z�X5��WHt�u���=R�e����u��_X���]�yEW;X070�c����M�� ���w9�x�YeV�y��I+;].@�ۈ&쵛��n��-_�ǝ u��tK{Q��wϱ�4�d�z�d��<ܖ�C��V�c
�u��];Y�W���̧���0�v���[5�>��^��Cx�]O��U�5���a�o�j��@��I���7=�7��<�9��'��&o(��p�4*kԎ����Iy�_+ҹ$�x#^� I�Y��ȧQtq�;�x<�!Tv�3�%����V�N����S��U���*��o���Ȁ��uӫ���p	��{/JI����2�a52�	�`\�WUz�1�
�u�}���S�ަ��_/P��6���|h��=������a�!�\��<i��>��Wo�&:Ė|�:�;��xu5�[�����f��\3��3�-Y�5gmЕ}�i��)=uܗh��������njf.�^�{EO���}�@��!$$$$�I0ϙ95��Wn;^�l~���!��P�H$�gn��D��GOwj�% �KU�'x�$V�#�nR<^�F�i���p��鼯	sA�Hە�q�WV6�XZ�/�麞�c�m�!�r�
�j���M8U����7X,h���d�յ�X�l y�R�M��4��*򰺺�%���u��֕�fU����3|�+6��/)5�0�ٙ��.t#��t6�i<�tSqZ�w�.�����*�*I�P$ɖZ�Ӥ�}�=C"�3C���72�z�{�H�z�gn0���|io~�;M�֣N�m�O(L�'c�uJf'ܻ+95�b�,������Z5�%�=,k���]��ki�t���+pG̎�� �Dy;{�nZ��lE �6������Y�*J�$��O4�Ԗ}�Gp΍YlW
̝j�t�ʖ���ypm��rL�{V�JJ�-��bӹض���#:ݼ����:�Ζ5Dͼ�b���qvV����"�֔��p�!���,
�,�eel쒇6E88ው.�Z�����XH�+�E���������K�hkzrѺ5y'N�)Wm$N�s�]AQ�l=�ݧݛ��ХѠ��j^���t�|�8�R���0��QkK'
M����1�U��O�A�����L�/9CtpM���vQ�Q<��1b[�gn�ԭ�k;.'Z�w_Rz�#W��������SL�B��[�}�k����ՙ�k���Dop�嚮����]0���{ӕf�s��zwwI&6�τwg:�q�줵�h�N�IQ���Z���G۵���vsԷ�-�U��@���)��8)�с
@]��'VE�A�v �J�j��Z������t�c� ��tc�`U����j=���9O-��%�)�-5m�\���w^_�~b�~���K2�e��fh��;�֖^�Q5�s��ٙAO��%iSy#Yv��������<�e��#�m=�f%����G�ݰ ط��ȶ)��.FU��&lV���.p��n��-H�������C/���ܵX�:��V��(��m��;�u��P��uM�]ڈ�,_J��kJ�ݺc:G�ˉ�[��Sy�h<���S;�_4�­�E)np���ǸX������|��.+SWvl��8�㨉�WL�=9,�h�|�)_h���a�6��D#�o� �8={XhhS�f�jX睮tM,y�t�N���j��V6��U��b�]�	#�����m1�H�
t5@��6,Kv&[=�A��v����~l����W*yV�u��t��^�2�Vj�J��&;�F���|2mu��V�ޢ;�w9���5n�)j�p��4ui�J�T�iv���F���޽�hn���G;]��Ue�r�c�÷���B��4eӮt��q`.�K�Yǽ��Dpz4�]�kyv�"V������aH7߻�{ѝ�l�,Mr�e���,�e,!�V3�UW�ST�A����-*�G�� W��m�@]��.9�y��s�e�y�%ϗ�iwO�4%r�Y����|�;�Cv侤NeT���k�&eO�3��U'fϑ�P�u�;|���+�ެ�޹c�^�1�<�V���̯=^9�������u�B���4P�O��à+ݘ�,�}�s/���@59�-ιs�s
��!K7^g��~�*�dW)��t���v���:*-��c6\�ܬ��C�웵�o������\��n���#�
�jD�"mqc^�<W1j���q�����~~�Wo�ʪ5��a���M��(�<��qH�l@��oܗxz�zΏ���hV���Xj3ڧ0���Ͻ�f�5�*Y��N^��~?8ã�:o��]'S���b`��v�]zC�:�mp�<t|���p)Q���;�C����0D�#�zfOQ��%��o\�灚�[z����a]��0ĝ�4/����s/���N|Gg]E��}���q�{�_�V,�;�f�{&�ю�Q�]�*+�C�c~����m%�^͝��0��.��/O)�Vc�:��0�Ƥs�<�������HQ�g�!okؒ8����9B22�:�𫆜O��I�u�$,D'�!6���x��3��� �>��5�0��/Oj�/�1�"�1�k�=Eڭc8�S����V�mLWZte�C�s�;�m.��N)��v�v�C���l��^;��wÔ��U7�y�γ��r��3(��T�z}�R�~�G��j�t�I�1o�f�F����FגGK+�����``o����q���&`��8n��*݀���'����+�v:�6�$����n�%-�]�@nl��.��j��������:��-�R�����Ƚ�&�*�r��3hC�Wx+��&���p�+�])�]>��h��~�l�����f�u7�⫡:�2ga$F��Y�L��j&3�g֏%��*_(0p�du)X}���g����K�:6jx�5�}.d��Wow��Ϛ�лS�\����q�@i�C�b��4�I#��]�����l�A��-U
������O�1|�iv�O�9��;�N�������zp��5�٧2�ǣ)�� -���Jm�����`:,W�..���׃;��+2Ɲ����'�X��{��KWVd�֫��=>Ñ��}j�e���3���Nic�������*��S����O8�Gt7��W��[�x���9�\�; �@9T��q�Bn�;�~����<� b�jT\�Bz夋���c�@�?Eb_DH���(�X~��Ŷ����
25�>���&�ɯ4u��P� ���<R�.��i��ʬ��2u��^Z�k;MoLk��+&�L�XQz
:\������X��K!:����{�f�[ݢ�ͥ��;ٗB�� z��y�_K4;������U}U�N�}Ѭ��7�w�Ƶ�Ip��o�Ⱥ�`}=&��)�%r�إ�jc���J�� �8�+�;�v:�s�@u��j$�S��E*���3߳ZǮ������[�����Q3T8���%�V�G���A�����$�}�q��7�c�N�Z���s�H���P�*}�5�}�c �A7�ao�xS2�)K�v6����{�|G�bo�c�5�n���.�O�	�1_|ay���)���u��ÐK��O���P����kT����GҢb��t�{���^McZ���iA���N���qYz}�]"���ѕ��K��o��b�[F��WD�&c��>s۠ڊ�]R��B/4���	��&fyF��:IG�f�agBP���S0C�B���@��%b�=�]��J�h�[~�
/jY>�lޱn��'���"��F�+����ڣJe¼9��{�f÷�+^VvK@��R[b\/U��݁�i���¡�Sj���Gkx���ܵ�/�Ef�(h�b�
�q���ీXT9f�!�v (Au�~[#�ӗc@<��g�l��U�����̗7&��%�hA��u��"�q�]�q�������i����ȯ,��'
F2lmW_������cszD��ڂ-��׏ �35�Wlޘ��3���͚���k�.���rQ���F���*A�8�����S�I��0	��v�/Q�75g�"D�b��NkD���q^�������5d��e��^E���%�\;SbZe=ΜR��i�2��ָ��(:��G^����8�Y���D��_VТ�rx�Ü;�tn�͓R;��Ʃa�j�y�9C��L7�U�}���ЁK�B��2X����Ct.ڿ-���ʹ��\�u�62�>�dm.�C4_��*�SC�����ԝ8�+�G1A]֮n��.=>��g��×�V�(˿-�_[�s�HU�|h��Ϻ���T��3)�����Ӗ=Π�n��{�eH�_m�G����B���{ ��u;狔X���(��|!CۘՕrD<#�
�=0��8ä�E�)�ݾ�>��j�郝�4P~<3��K�Щ�*U�&�Wͬ@��Eaڵ�����]̛��˳���B�kg���ő��
*��b��pb�V݆t����Z��BF�1��=�Q�4r������y����8מ�!u;�+����;�>Gw5�<'�0wm��;t�ZZ���Y T5�\!k��'��R[䱬�3z��*�a:�w��ں�!]xA����mà(���[�?+�5��k"�b�te7<FP���1�!|q�t�����fgU�W6����z�2�� _��b�%���7��8��:���}��ɘ;y�yW�8����gY�(�n���J�ۨs,@)	V0�A���0����%u�	_!0�Y�v�δ΁j����ց�kJl�V��/Ss�h���Q����y�d=/_)�v=x��\�i��d�U�Awx
�N��#jsn�z��U�qͮ�kնeu�0o��CW�u��t�A������I��	�D�W�s�Nu�����o��I��Ǡb��?�x]����ru� �nm������'#��"�����ԏ{��u.j�)��?i{?qU5S�y9*���Y�ǋ���g-��b4/M3[�����K�1������-��Uph9Y�������-�?�z���;�?ZƳ&�<O�|����k�7������n�ީ��]l�M�V=�#�ňj���t�_����nߨ�‏���F��ތ�u�������Ogt����
���;Q�}�_g���7���w*ibz�S1�=F�mrF�dN�-�5Ti�zⴊ�f��ɋ�<��|���v�>��5���]_Z�]m����;����/K�h�p�r�>����ްP�q,�
u]����gj��t�8}��+xYa�˧���jc5R��%��*0��9�!�S�d{�p��y��|}�q��&7��$5������K��U�cv�sbz�+I)��:�s����H�_:��T&�/�ڵ����k�[~������ٖ�̪��9C��n��L*��S���*��|���J�OmL���viY������Ɩ�j����[�X����`7p����Y��b�ү�]6ދg|0m<��L�#=��O3���qu9)[_^{��YΘ��U��j��~�wDQ�5�2�;]}�x�ck%��]֐�y�������Ǳ׳��c(�,z}�~�1���Qүj���O����������<�h�WnBV=����S���fЪ��b�ϛ�*M��N�E�R����pt�>:�>���9�' �ZF�Ԋ�$���բ.ߒ�1��^���9'׷�w�'ײL�Jeg��tK�'��3ϵ��2��+!�ێiT����ǎb�9�@g�k�����mY�������p�h�t�LkR�!,��>9X�GM�6&[���?�0�G�\���˓[U��(���墫L��$(Uοz����fb}�}<�5��m{��F[N{�m�Ɍsy����!!��{���%��9{����ZKɐx]��[A{-�v�'�����{)iޔz��k��Z|�}{W�C�̇2{Аߜ5�=��1Q���g���+���8����[b�:U�=ü|R�	K��c�]{�Sō97;uٟQ$�w�����_`C/d��{WR{����x���
LM�X����y�.�^vM����w,��o	o��N�L�̷�f��ar��Fo`Ձ�Th+�cɤT����6���]"��L��Zgk��;}:Δ��]9�A��y�H�u+�I��Lz@�(h�r�!��M�6�Ҟ
&]��K�{k��,'�x7�%�	���������q��{Q�_�Z�ұZ2�y�)K�_�>���]4i߽����=��3E<\N���Y����ު%.P��lK#���k*/}�	�f�7���:�U�[Jjz���5�u�d���@�Pt�1l&�)����f����Z�ߢ�x]Fޠ���4�T.��<�S�����:��QJ1̥v���f���mY�y���=R,����^�e�鏻���L7�V{˭ab�����:�q�S0��P�+���9
1�9�b��Y�����1W��wUf?\�	u��k/�Wǅ[���<�<�ƽ�S�����鯆Sj�Av}���� �,�y���]��Ў}ԙ����̲(8^�<�M�P�MŢm���}D�y�^�P���{�-�<X<�(ڏeLg�+�'���s�}�t��c1m
�7!�Hs9~��v���^����k��Jx�2}��Y%��S����F<��e)[W��>"�������[����Y��Y��:�����5P撄R]��	��zN�&,� ����ۻQյxJ�#��]���O%G�k"��YGs}h	�[R�
X�o-�.��g0г:[���:|qb+2(�/w�jq:*^�kޚk6g/���N������$�=�~V����:��2�HGU�~��w�̯e�6��g����s�xůQ�[�o��M`��1�%!}U�i����>�w�+qyUI{6 >C����x�V.�e��o�A26Z��#E����[=���\��p�߶���z�ʂ�''m���M�����js����G,��`o���{=e�m�Rҥ�����'�y�Q���_�����|���B.ݚ�~$�&��������O7�����Ų\2x�ċB���/��>�~÷ �K�C�3�}�5��S1̊��c}"�s��ͬ�Qr���I>`U�qFP�;�|nN��q�h�N�UTʏM��7;�%ufVp�R�CڽQ����(AJ�M��o¸�ol�OY�m<\�CI}ꓷ,
���"��j���R�.m|��U�N<���7O�����̯	��p���cB4i�L)�p�:��O�L�]^H��+�<��ICϰ�k/�E�4����s��J�.��9��U�
�Y&��4"�?*��է��h3sW�k���O.VٮV�E;�3֟X�F*8d������}]+��fkRXLb|����F�w���V�
꺇�-تlc���f�G����d���V!�n�+��z �[w>o޸7�Z��SÓ>���z��x`fy��ܼ��\�,	��f@����s'�1R�D��4��80+��jnS�Ԩ7����Z����_ΚD�8�I��Xj�]��4A��΅m�	���Y�H-�gc`��ʾ��G%NU(�7�V�k�v��e�P@���y�h��(S���[�����Kl^�@��
���ᙔVls+7�"�M]�<�;w�ډp��arh��ϣ=�;fg�緎�u�*� zmw�aJ��3�޼����(��
x6u��fs�7��S�9*��L��tN�f���ĺ��}�ۑ;^-�;:�P��ё~ך2^��+J�To#+f��l��0ƞZO�oMɷ���PD*��59�D�Z4�a��l�yW���aՃ�ng��wE=�I]F�7�)P�|X������XoOsed̼Ӯz���
^��셇�#n�<pX��3�̱.9yr|�Ҹ� '8{r���A�k���.l�A���K3��9ؓ���kk��ijQF�;Oa�o'��
�ٜ3��l�h��Y�r���K���,���QƦ��*�A@����3VPi��ڜ��N^�U#8�gQ'擴�RywX�&ZS��Ͳ1����>�A�i�Q�J���[�
�G�C�ϐ*��;�M0��O!b�hr}�f��r~Y��c�,�c]5.I>��7]��{|����ɹ�av�Wٞ���Yj/� !u6=䋮�����Ê���ʀ�`U���*�r� E\�9�P�T.�L�~X��m�c�L���<T]�U-s}�x�O5�=�4�M�_ ����<��)��]�L\�8%��^f�����d���ov1ّB�H/�����w�ԳΕ�ju���8`�=ϧj��W���-�F�)��(�,�A`�jIH��J����sC�� ��=0�ٳonW�-�����ni��Lnd�E��Y�p�m�I���_��5z�C����zgz�U�ȩ�'�*D2=D��]�s���҃� 77��_��{3n'S�]v�Rp����
D�ɹR=j�z�@q�A�
\U8�w^jLn�z���V�.Y��/'�6T�x>\���S�t+:����?`�>�WrG(^&v��~��qJ��o�����V�n��j��/��Aq:n�KU�MO#�ZB�Cd`�_�e_�z�۽��>S�QMC\�/LOZ6v/��(�?zS|�gs`[݋U\V��u��N��F�V��aS�GΗ⭪���q*�k"?�z�߲��W쓞KN/�&	���*����+��?v�+/u�ᗲ)����&���쾹�OBBO]P?+��-��e���T��催�ǫ���l�_}�諾^��`'���+5u���O��`��)�5���1�����]�ť�9��\���]�(x�7.��nBo���k���F���cFs�V�ԗ����5���}��Z�]N�j�T<���u�i��l��KE
]���E��Ρ�=�J��B��d.�q�3u
��|��}[�lv@�K�н疞~��-*E��mvN�HN��ټ��ĳWF��訝�<h�I�e�:]�0���b�c�D�u8q��ż�Yƥ��9�Ԇko�'":�J�[VZ�wk]�sh�6���,�N�ѲMͮ��Lp�G�o.2������J[\�v�'�,7�U�t"pj܌�.� vZ���(�KMrpi���Q�q�5�,� �iR��ݕs;S��g�TM�;+d�|s�����N7G�r}��4n�^�������9&��Yu:52�� r�Y;X� ��y_
Y��O������-A�����,�G�[�]Q�GE\�\���?��]�']���K��, G'=����fJ�y�|�X�Ы��7�V3�+��.mǺ+��hԡj�9M�3�b�At6���6u�ѫdg���X9���f6+��o���ܿe:=A�),�p9���s:�j�ԇ?ćg���|p"�AA[�dL�Z�,q޷1��ts�Y��	1������Zd�a�ޛ�vwW;�6�rr��z%�X�"g�/s���V��.g>SX���o���W�MZ�kkmKt�����%�z��
�	2�+_�x:��ϓ��Vמzw>���I��Hy��D��,ɔ���$�}�;3d�sCD�8wbA��y����tX͝A++N.�1#�:�sq�S��}1�o�U�z�>�x5�*+W>R���ف�C+�'������P� �l]pe�5��0�we����	��$+%M�Y�;��틳�nl�MG]wg�����U��3;�p����pԿ�Y�����f�啡	\c<�ê��*I�ׂ��5)EY3{ Y�PP<�M�zZ�g]A2S�qM���C�C����˽S�zȡ�\z�DL7�r���[;q�jE �OuA��2��&=�:�B;@:9������*|�-7ܴ�$w',�ʶ�!�ٵ|{�������+�q�=�u��ܾ��;��ޝ��ϩ�I�?�ƽ�;~�m���玞Q-���wxE��'w֝�r6��)��obo;la�J:�����/VR�x��e�f�[Y1f��Y���^��)�<h������-#���x0��I��em�V�,qF⣱vPy���k>�'X S���S�j���q��� ���XmDL�Gr���}S�0*�|J�Vt�r9Oc��ܨT�̌��&�xZ(��݊H�`�_S��}�ە��Nun�w��S'����`�w7ź�%Ǎ�^#Ynz/��Rͽ��yH3:�LV��S���_���<�o�p��"7qb[g�Ǐ�s�
�" 𢅩�˻TXZzJ��^oJ� G�x��@D��q�pL���'����j�o4;@�opj��"�;�q� �"���j���r�#Ԛx�ղM�W�ۥ�g�Y&WTV*�����+�!K�wHgy�~ȨԳ�R�W�*d�BP����V��5v��R=�n��d���}}P�[Ps2�f>Ӿr��*Eϳ�*�E���2
��*�]���y���<�+�/`�jj��1�&$:d�����qi�ڈJ{�#�\����\��wl��#�K����4sZZ����#�����V��p����^�l[�=��sx��u�<��'2�����`�f`�"*�����CN{oz�$���e�*r,�r~�v��*Kk�R}v���=�o/��Z�	=	9����ד3Iq}��k{бҝ
�R�鉼I��F35�-�]�㊆l�»%Z^Mԉ��BN��ik�)r��p��y�cUE�̜�Q7����tl�,X�^OT��]s����:q,��@�EX��Hj�Fq�ކ��g�R��$"@�rYTm{gkD�h��s1=��;Y�;���:@�y4V�&� z=QZꇩ:����tK��(ySZPQ~���K�#��G��K��D ��ح�� E�T��bKar)7W*I{��[f;���s�����Γ�=�<�w-7-4��2��Ou�^�2Թ�>p�0�v�����ht��v	ط�	�N����T�։�QRiodN�v���[%^l��Ç:yPŝZ���c�˝kֻ��s9�/�&^eKT{(H�l�g ��ݙn�썕.�	s�Q5�A}W1+Uud�H��+E+v���7q�;�2Y��nU�_g�z�XGD�����Eo߮,�R�������sHGO�sNm��(ײ}��r�9�[��Ù*���(��+��W\�y�����4.�E��U��������t�ܓ��3��Q:;u��)��D����;�i�M/j�ǘj�8<�o��:���M������gZ3'��ǅ��T;5�i�3�WQ$���I�f�SV���J7�F�gUG����x2��(z�@=M^�u>�sy�U����=��{s��6�7��pO�z�]����O�����Q�.��k%6���9}��B�	�0��IQxU�jqb�B٭�*�����D��a�c��:��բ����WX���g�볗B�:�ށ�..�Sp��:���7�Pn���>��(]Z����+:��^x� �s<��̰:����q6�Uo�|3���J�z�Wu�e�y�R�Q������:�=����Y�Qgr��bQ�EB�H�#�L	��xx�����fD���2�m���#��m� ڟ^�W5ɶ�j��JJ�-�u�p��OY�Z�����2 �}>���j�U]q���� X�'�8d cB������@3mv�
��bd�V贉w��8
Q��Hh�~V����}��X�rQ}�:M��=�������q�.�l�t��I=}\gu�G
דE��f�˖��lrԤD����h|H����5T{QR��WKN�ϫBq�nv��[��KO�Xz�C:�1��]R^�,���C��'��鿵�δ��g����ٚ,q��HC9�U>6|qlUI7�quESU�r����>I�댁^���nV�Sܬ����l�.�'�,��嫤���/~��y�=n����b>�==o���5�jg�%��]}���@�V�[�`{z�^������5;iQY����Df�Im�1c��>f�1��$Nl�5V7ۨ�u:ANś�(E���̍>޺��<�=�Lʣ.щ%ל��d*���Ho7G��ޥHS%��@�!R�]DӧC{Gsp�Ժ�3a�6���?:+2�'zfM�)�?�e�'����6(|U>]�ȸh�]x0-g�������L-ۘ�d�V��k�TV�F5U}�n��=���>l�E�qL�/30A:7뀰{նU��
��'e���m��XruziL��
O{N�b ����U���	���$Z����Mf,���ﷳ&�PkW���.��j����[�ˆ*aqQG�#�
����KZ����>-^��B�d�J��B2���y��1;>��B��i{�.ݶ���(�ȕ4�!J!�t͛��fw^�h�$��u�:�c�j�%�2�V�v ǯգ2��)�K޸Lns�0�mJ�%e���V{k3�y��k��ΥcB�EI]�*�&
���.�7(�kR���h���i�k�]J=�{@�/����0`�e_[�+��B���3��"�Օ���Iwdl��!qZ�鸐v�&���:��%�]5"�+a����K;��	Mu�[ߺΞ2'k����,����I�3�;l��i�7����y�;��L�q�,�N�c'�,K�m�^�02=4�}z��o2`Ɏ�4~^��m�U�꾍�8�d�WH��<1k{�!m!"�0���R��T��X&E���+T�\Ƨ����J�V�g���[Hi��fR'WN �nq(��8Lu�K�6��/*Q�]�kno��Ӥ��m�,�K��Zm(f�÷ݫ��|�U��M�Mo�����^I9	du��`�̞^��
�%m���ѹ�{��1-7�q�:���׺Q�m2#�rb`[�T<lh���:O�s�G߮�\U��Wut�w��{�N:*���uu��>�!�191�bpƲ�1d��k3E;��="�\'¥tf(+m�dp�;��3�áf��ZjӚ�|�N-�dk��.%y�nA��;�U�v�����w�pH��W�ݟ��6]�."6���L����Jv6�kG�=t|Ϸ�3�����";��U�f���
���]�,�B&/��X��~�\1q��I��u��*�ݚ�V��5��I-�a�^�9�ez�`=�k��2СuR�f��DȂ��5e�)oq��Rh����k����\+#�¶Nϛ˺H��
�V�2T���OV�N�FF�J�^�ud�VbŁ�cI�5�D<{Q��ۼ�t�b�r��m�S�KX��QQj�˸N����,�o:z�M5�����}P.�l��3t�Jm��]6���ԑ�ʚ�Y�WC�uCiH'����>�~��I{�U^1�zj���A�+�2�E�z0�ىٽ�6VyZ��R�.T�u���Hþ�g�N��JS���B�O��j���{38�">�w�-mN+��kA����XNC;�*H:�Ϊd�k�:�"�:���Ǡ����#!�
�mKʝ����p�g>��ת��<�y�@��1x�v��n�Oi�.K@E�%d�7�� ��Nd�TYcUƦ47����.��^��Gl"�7ד��s�֪.ͨ�U�r�tޯ>P���tP�f�����7���'�:Tg	ԠA���V�~�U�YՖ;\[:]l�2�#MI����U���9��D��On�8f5�n���!��H#��ʤ�jgݫ�bezSʽuR�߼߱�Uws�(���tV�Ulj>�v͚Z�l�q��-�&v��wܻ�6�����qq�y�v��ܫsKa�����(R=3Քu/uPm�j�x���w8~��y������~���ڶ��+��k��=�������:��ed���sS2���mQ:�'Ѱ�h9�j26�^wK���a�G���a��;�^G;S�t�cV���;ܥ�qo.}�p^<Y6�H�������u+�Z�շ�r5Pʷ8T��M<�VE���A�B�,���;�v�`�LR7J+�um��ӕ1w1�du3��yp+xi�98���s:��UZo}}H=�{UOf�_g=���bWѥ�ذ��/uiw<�XVчt��,]oV?s�rϧ��T�>�zz-|Ь^�B���q�=<4�u?E����	�<�u&���^x����|_������'�Q$/ϕ}gfu�=�qoڭ(�m+��(�����RP�]����#�/�&OE�7)T��"V�%d���P�5��㘸�<gpL»s���b�#�*$7sG�*�ͭ���[Cn�ܤ<��k�c��H��21�|�è�qw,}�.q�<a��x!�-����JW�K�8�VqLz-�>>�s`�X;�#rEg9S =��s<�{I��*�i^����4V"�ǧ�|�w��+�s�:���Ԕ�|P��~��Y��-$��!�dM�IǙ67({�g�Bp|��:���7��L��.��.Y��������ឝ*����.�>��0+������b�Up�\�P���J��TD�P]���<������,�H�����PZ{�-�+g�֩{���i��P�8�+zq�y�΅�|�i}�T�Fz�n��+9
-e���\ ؁>{:�-d����8��}f��ȨR�!]k;1��T����F�V\�����"�J���a�3�V[� ���l�PYZ��5ٽ� O^��˼�̮���a*w@�^�+gsʴ��v^TL��Ǫ8�δ�v1⮍��y����0ڍa�`�@�-"���䝸���S��M
3b�����	�cB��Pj����ٙ!�{�'�,S�.��5:=5�S����T��_o�Ҝ��Ն��4�W<Ε"����DW���P�9v�hS�t����2I��Y�LC�X��Z��{��u�65!`ҷ�z�ƅ�o�;�pL��˨��Ԟ�pCk�}Ժ����@c�|:��͟zj!���\�nEШ;�&�oeHb}�uG������g����+�ڸi�p�����)�ǖ��nQٍ�-!:�C�'r�����@�-J~
E)γ���kjf����\zr�9���[���]	LM�魚�ah�*�=y���_����ˇ޾xQx�lfa�bByv��O�C�wK四3A�6��c7��de�S2$�Q�'��u�='2�궟�=ň�҃5��	�$ED��>$䵆���3)�LF���z(���\�Cp�V�ڼ�"iNOU��������Pӈ���*�gbw
w�3X+��f8v�9z /���t��1����ޏ��`���.��2�SQ��N���ĺR��;��{J*�NɊ�1=љ�[�{�Gͺ�,A�K�H����:�}[��uv�31��'c��K����Z]�۷-��F�B9˸�+0�T���L c��vM�]�4��{�o��+u�vk�Q�w-�6#�JӔ.�ɻP�y~��X�6�S
�AQ�
���=�dtQ��ɿ����P^��%n��^0���N�qoA���o�<#���)����6�,��9�;H�Wt��O�T�`�[F��A���^���*5"0��K{+j��*'f�g�)oӘ�Ut3��x8�.;j����j�~*ǓY��lfjb� �콝ɫ��84T{2+��fX=#��Y�f��v�0�Z�k��(�~wx�D�JhY��W���`���-�I�g#gY�\�K;2��d�L���A���m]{���k"���^���(���ػ��s�cS��u�^��1�%�6���{�#��j�%?��{�w&���Z++�0%��m!$�r'W\ꇤ��3�%CG�˧{�r����8
�^��������9����(��Mޫ�v�a#'T�����d 	1銇{�T���޻��ܲ��nvz�]PlVʟڰ��>G.Q�M�F��FJ"���#���'z���3�X�f%�y�3�҂Mz�2%�@�ٗL��)��'�o��io�O���kO'+LƵ��C5�~��!�3U��q8b���يԫ�4
Q�R��#�nxj��x<U"����!6�WeE����*�� 2�T�!�G�܉�5�]�6����=u���W�&������2��/z�ǚq�en,|�.��|�)v��Qu�Q���y��;�Q�v����qWKb���*.��������9�RZr,�#��ٍ"˛�CYر-�?g�
�g�fgl���h���'T{�Wt��=&���h���5�)�s�o���3|�j?��{�q�Sn��d�0�QG�7����$����6	�j��!4�c� `��+���~���1vy,X��.t`��/(����W�+�1�7���ڃ�u���˿�������LW8`����{]}G�ɑќj��`�ݏ�"s����s3U�har�=�9�"1��%j���*�h�R��z)�z���
�.*�y��#����(2';�L���Ԯ+}�uʬڭ�R�s$(5�s��4�Yq[ٕ�|g���3�'oT&T�yTC�\�G&W�~�W�(�}g%M��`���QR�Q�xk������#(��?e�ܾK.p���cU-�(JHw���!B��^�ꢤPW]D�NCA�,ˣ]}2����Τ�]�=1͹bC�K�6] 9+^]��w��Zw��x��h뾍X���}4+�ȏh��k�M�3ݟe�Nݻ-I�"s X��`��M�:~4�	��fJH�1�>�}[:��}>��
����s����9��g����sJwq�n�Ɇ��$v\K]��o���t��~0��Fj;�Wfѭ>w:�ky9tvT*<�2�W�R�@�Eo�k]���Ԣ�)R���������w-����l��R��%o- �s5�M��A8���;�L��娮�L��<\w};�S���;��q����զ��8��y�C�o
S��)���i���Rrw�����.mF�#���W3�3��>�-�W/<����0\����g{m���2:+f�1_<�Ⱥ�7φ3�A�Ȭ'.�:��ˌ��Z��Gc��l��eLPIg��/v��GEұwz�1�s{Hz5vz)�>�^/���O]N��d�����w���kb���{��s�;9�A�|2ik?f�V��xw'j}�(�wH��\O��t�slq9�J�(������\j��{p�yF�~��,I�6��q��ǚ�����(�W��б��ɟ\���8�f����"d/:;��UJ<˨s�6�ݼ��aJ��GC��w������)��6ݷgd�)��ix��}p�=�9�7W�׉�WN�F�c���fxUH�"k��X=!N7�z�	��2(�yb�e�ħI��J����N˔M9����ۮt�]�g?Xu
ʩ�b��b�넚�9��@�^�Hy���M�h����9����o�2Vg��YؿF\����:#̝�j-`GA*-5Kq��ϥ������K�캳�AsNRJ{�Ï�r_��,��Δ���L*ͫ�	�i�֤w�W�3�;�B���п�@:nZw^W4t����ȸ�N���'�вG�V�Ʈ���W?+�h���'�v��}��}_��ꮈl�[�k�G�
h����:ᶳ�iT�Hv��T��Zl�]+�;��v�[37�d>)a8:J��jh��]��W�9�3�Zg����(�N���x��k�H�>����xC$�F���QML��y��j��}�F�U������铦r�a�60n9�F�Q�8�hy;��R�޴��^о�*��Adӝ�s4R�ߍ�������r lI �쬣�Os8�J���D)W��"���eRoJ!��U�����r`��+�C����y�=.�����G4�W7NMW'JY�A[Qucv��j[SD��f�39�����cM�sI��t�e�����a}lnlWFe�4y��9fo��o��mk��j�"X7 �C_=�qīmu���}[;/""��뼵��X:y�g4g*�ܷ*"�^H�:��;(�Q3lZ�p*Ձ=+�*�畍�݂�}�d췐��[���?m�b1�.�tzU�cJ��ؖ�9�B7R91d�t�i��͕�{zԥT>������0<�d�ʲ+��8A��; ����7�hM}�����S�w�����\���/�/�����zt#��5���8�l ��[7X[�`��U��0�x��x���� ,��!���.2_i�a�7ܑ�)oD[�kKۊ�
�.����f {��� �³�M���U] ��JDf�gd�̛�{q�ň�tM�p�.l&��X����H�}$�{�s�ĕ$w{�s�m�u�p�v�$vk�ֺm�Y����M��ƻ*�R#���X����BY�(��s��r�5����K�+�"duh7��Cskk�̙�W�I%%__1Rb�z��;We��2AuJ�<YJi��T0:��/g-Ս�u��$viڴ$�,%Kz�*M����}��:�k,輶�i)�.k��Yaov9q�,�B�X�������ɘ��^̇ki�畜�\��Z�r�ᾊ����+0+�"3�FvW��w�V�-}t�]�5�p��,�H��=[t.�vof�]ͩ�З�5��ܜ�kv&��.;Wf���bK��NRj�n�pdt���H�`}�Jݨ8s=а��c�V띡zNYA@��wM���qI�flR�������C.0�r�m{),a�aP�t����k��ӋlX�yJA�J��bIofe�^V�G���XP��0���GbI�;H̷�͛�R����sE�d�1��oa(����ĳ���G���J�j#���u��2wˁÝzg.�2��+���k��s�:��$��d�-�>����}.��v2n�ݦ9O3o�twv��vR�u��;C���8r��ə�:�e�2*C��ƪ��+�0��ԟt��`�lq���4s��V�b㵏��]��5�Yt�ݮ��_e�W0���>���L��`n،���-�i�ғ�[a��^6�v���{�>�e0�_����ݹ���U]ŝ�6�]�Dx�~Iq��w�7�+���}�y���2<����"vz��[�͆��"�W�}F�~�M s1��L>��k�4��C�
��~�9&�%�mgeg� @YwWU}��5�D;�O�pߣ�p�IeM����
���h��J����eJ^�;<��pM�WcDԔ6R���F:ZW����P�}�=ܬ�s��MJ�A|��~%誼�
���Ԫ�9T�l�F(�)y���ȏ�JD���ϣ@^*��T���ٝ0M��ɹ�����>m�(b˹�n�����" �kڪ�'�!�䣰z���ۨr��xE�f�R�n����%�Kf)��"7]��.�q�i�����
����#)�(fp�ޅA��P��QwO��a�0c?@S��+��W���̻���:��坒�nfC�퍎Z9]uZN/1�k=���/^[ �W>Ӗ�7��)��3A�t3���b�uX~G2���7�S�L�ףNJ�Qy�ޚN�eK�n�}���A��{b"0��v�iG���<r+�Q�N��.Q�}[F���	p�����W�p��vx4��C2������{����]Bn�prR�z_�j9�^�a��vGz).k0l���o|[�F���S�&A�3�{�ɉ�	 b��N�]= ��Jڔ:S��o̕�_�4�?^_�׶������XL�S(�R�ǝ�ł�\�\(��Јjq7\�\�3�3�I�&e��|hQѾ���z����}Zdg��c�`\��·��p+�5M���վ캐��R���>y�� ,�bs�����/�Q㊟��MɊo���*/\���T:��ު�n�< ���C�!M`�?G<s�n��-R���+Zͧ,M���^��Y�Gn����Fu	[��t��o�Qn��R}�l�On�y��x�x�-��X�s" ���mӬF�b�뺵��nV�eBRJ2�ˡ�޳4��N��Wf�E�ߺ3«�u&��p���Lt�H��=���΢�Xb�:�	���Y�g�Q'����z-S�M�Z#�9�ܫHp{J;�[){HO;��m��(��r�A���2��W<�����w��Q�PM�hҴ<��=ޜ�����њ�?��zf �F1"�iB	���w��(�<�Yd�%��oqD�b �H�!}��U�TXU��q�o�-N�mY>�x�,)D���9���#��\�b�33��[^�.9���kכ��]I!�c�{���|z�݆�uY��f�^5)���+߱���,�9\���	��n��SY��:jiȬվ�
�a�Oj&�Ѧ��0;q��Z8
��|��n#Ӆn;��e�Wr�rN��~o��N�[\/2g�{�r�!5�G_��Q�)�B��J{eaO^��1��u�ʂS�f/p��0�-S�g�u^:v\s�s���$ WX�!��*]=�����W}np4�spM��_1��MV�O�,�����-l��R* �ʳA#��G{Y�t��hm>�����Ņl��S�g��e�D<�n����8.��[X|�=8}���GQJ�T��V�2�aawb%�I[n�z<j�6���+ǆT�W}���w����z��ŏM=h���T��w=����6z�<��,�C��œy�ߌ[�;���)�< ��h'��|�{(�݅��3y�S�!�Q�5��Y$Fw7 �q@U6�9S��\�7=�G�U���xȍ����R�pQ��&ϖ�<:$qVΙr�̂5��\�UM�g�hP�o��ߒ�8b����wA�����7��Q1���ME�����ǽ��}�����ʩG��G	l�.��	L���e���d� �6?b�(��/an��l����y<���F3�	�q^�i��ĳ�vL�����g����|jY�Tq���(�rT�)�׹��7��YSCw5�������]�EL�Ϭb;��OK��Y�py�5�"za{�3��L���z�LsB�ׇ0�~�fhSQ�S�6%'Uͼ�ɩu��.�P�
 ��0"^M����p�7��#�ƺhX��"8�p�w��7�ΈC�7���۾�k��d�F#��{�Ʊr�+���4��̝��q�G����W~�}c��O{�-}��E���Ƿx*b	o�,�M�p:͸�</̈́�L��kU���9��0w[�ؘ��oJJd�3vSt��C���� VCs�����;�U�%]DN��j8��^=�:A�e`��\���=U�^u�����G������c;=�k�"h�\NqI��P� ��9�vq?_5]\����
*!biE*�6;�����gx�C+ϊ�M7��8r�۴o7�!}�' 6h��R,� �tk"���͔�N�~�}��>���>���em�V}��;t�]3;XC�Z+���B��� L{�>"��5����h�}�\t#��LxLg1�ڭ ��	�N
�\��K�j �1��k|G�;�y��vHD�믖�9�K=��.�-W辀V��1S�a�3�^dqS
}e{�.'�{���-��^$ �٠M�_'Cy��j���7��/r׳���v v��9\�H˘��V�E�sxz�-i�q�ze�ULx<�(�Z����b��zINߪ�.�:�eB͸v����r`V����Tw��+F@lp��8�Y��yH�f� S���~Rի�ݒ����${��[Rn��&���ݣ�Ӑ��~�ԍ��[��{1R��T�)���%�uj�����k�*}$������}�HV"O�U����qe�dR��r�Y�d��IO���Q�7&�������O
f&)."��>"��>t��M�+ 1{E�D4��b���_s[E�˨��e18fșt�7��ګ�7ٯ�F��><��Gu�s��w�%\�^��ܯ83k���_2���Z[�j��R�>W�.-�յzv�K��u�J���&c�yY�5��\g���t�[�B@��=޴BP@Qy�s����A�ei�H�P�r�d�94�Ĉ�p��\�<[C.�3d����/%��볋P�G���q�QHS��jtl)������gS�)!�����P�s=yG�f�><�cr���}y�i�Ə#�vr�v̢x��s����O�ν틿A��|�ٕԩ���,��\|�����vf�CL�x��;��o��y�\��ND���,�g1p��G!�U/j_>�)9Q��BMF�s4z�gܵ�0ُ��0Q��)T�.x�]�����e,m���XU>s7;]���&�4��(��:1yxuwv]�i^'��Cay�x���i�ٞ��c<#�|��m� o�߄K��To�`B3Ŭ�A�b�w m�ݨ�`�nj�A!^�}��zEbb��'K2�GY����{#ſ���rQ�(�-�����H��6�O-��讋H�ĩ9�j}W�]g#����7��-�ȳ#��Y�_eN�\�]K���q��}of��t�*�\�p�^���z�'�׸����"��y���6�X'�֝�ͭ� P��=8#���gX�'�h�%K4�'\/p��s���jF�`��}S\x�-)c�J;��[{Iʸ]�@�ؠ�n�j8�v�5��� �c{}ܗq��wWu�G�RǜI'ER\��o>����D��*gb68dً't�mw~R�9�c�X�^�,C��5{.7��_��E���J5�9��w���o��%�簅�{|��˜���,�*ubg(�ˁָi�2�^z֟&�1d�u���I���,�O]TD��5P�z8��58s�3p*o@��_C��>��j�V�k8+�5�ܓ0��]`7Ϣ�De�7�A�v,����	�ӱKmJ��'i�E��]DĜ��*�(���{��,�e-c9�%S"���=ɮ>9u`����+v��ɪ�g�=�k}o�x©�e�P�g=�i�ȎY��jǣ��Y�X���L���%:��"��� ���{[Ȏ�ug?�E���^�w
u���bP�䎎5��f�G���^q��O�]NlAȾ�T���y��|u����U�/�۶c>�ד�H9�͐Nf�^�V7��Sg�o"���z|&y T3�6���͏
�j'�{OUB�b�lZ�"�Z�#�:�(��g���؋�oǸf���fOl��h���f�.R�~���)��NY$M���:�T�3w�{�����w�o��P�{��w��D�0ڍ�Rwsk��%n�P�Cgt-ah��w����$g'}�rDU�k:��+�@T�:n�ڑ��A^�}�((
��pͼ8�Vn	�֋:�]G����sR��'E�1����eK]���GG!�h���3���@�X���0��򻣹SKq��*R����O�v������wսR�X?Q�):L���A?96��Q�xܘ�=�
���YY��2�����w��fi���Vf-;�/���ZF5����'�1x��{��./gzS�L��7qt���fs����܈��Zb����A3���}������LXڴ���"%��0L����*լ�e�]Z�|�~�s���ֲ]���:I	u��[ij�r����K�U�t���AS~Qh���;�/4N,j��<��ba����J>��'��:��k*%ߢ��i���;YPE�x�3"R�UəU̥�<����J2�e01 :5����t���I�3�G��5�b����\e���UUd�%�6Q�b�&�g|�uA�S���#vkKY�/��*��kĞA'��6~օ��9iWt��R!L�1-B�1��/v��y%�e���
��X��� ��K�L�Ve�+�z&8�S�?\�����s�I��1��J�T��ٟoW��4���V��gD ~ܾ�!���m�"�=[�Q��@�*��R��ah�nn���Le������y/Lӽ�o��:�Es#KF��>k*��u�m*�:&�Ԋ�e�9��)U�ru�hu�!��Q8y��%;�0��]�����̺Xk�HW~O3���i�]*׻نmuh���bAK۵��'���V���կ��8�Ř9d,f�2��n�����o�������.��w�+�����ly:��š��o�1���Gm�N�x�B��b��Z�V�~�/��;hBP�����E�\�/�@L�h~׷�'��уs|��{<�����6���'ykzҿi����]{;*���~�]T!m���7�Ǣ��z񊮛4���yJ_�t;/������.P��R|�Ⱥ�Z{#����s�\G�FS�ʮC�zgLx��R�a��8{�z+hʎ��Ə^!cм����(�0��[4�o�-�
'�myn	S#dTx�Uc�V����2�;��O++�ީ�P��0|%� wc����k@d�oM�<;��9s�5��Xo6z
S�j��9�/AL[�F�:f���q�X����x�t������7&���c�%>�<v�^�A<vs��"�j�p'��f�:�vB��Nc�3�ݯ] b�I5ޅ�<��*d�M̨��;@.X�TY�f�̎�) ���]�]��|�)�4N��<�Lh���ȄsM�%��1��k�&H���ʖ-fYZMEǔ!� �|�����ky�m��@2�G@������bx419o�5��ZR�+37��9�V\���B=h͗x���p�����s�uqa:�gQ�w���X��u���~����|�c���U�4n�Ț��օ&#�f᧛��u�Ԕ|�
L�(����y�e�N8V���ܩ�́�b�b��'�i'Zf}\�ױ�x�v[���,(ĉ�r�y����S�K+ې�j��W�w�L�F=� �ȏ%�*����?L�atm�J�N]-�]Gn
Ԉ�X�	*��!m)IV��Pkoz8q0:GO������GuT�M>�8�ob�V��R:+"�xnj�5�0��#��]�Qʶ<9��f9�c���V�Z8���Y�s�O�92�����Ip���i���UL{Y�15	�-_�鑽D��63[r�}15$��TrI�����jtaf�s��D�,�Iк{�Pr&
"�"��-�[,���A`�V�������K"��!��[׽³D�Pq1��aLf��G���a��N�c��v^�c�$ɵ��L������^s�fMT��ީ����ˢ��ي�z�}Tz��MR�%En�;|��I��m�M��u�'�>�dĹk�� ��ɣ!�ɞ�w�����uח�� �e]z�z���<c/g��'`�nht���/~K�B�����<��ಧd�O�e��+� Ԝ�J��[\<���`>��K�w��ľ�/�r�㖅�P��OA�s#E�|ӗB�گ�їJ\�YIX�J��;fL��Im��L%�	'm��y@e>��Jn�C���]��O��Oa�i���;���:�.|5�'2�fWk�缪NH���Ss�Nƹ�_!����qz��o�Q������yS�\���}W�?����̙�[g+����_K���=�so
5ʣ6�(x�-��{w�o7"2���j�y>����u`R��Kۢ1�a�-����/h��#,�9]"ڥ�YҸL���Fqǵ�ɉN_��u��M�zv:�Y�'ȫ~V㡕U	�ђ
�I�٨�U�ݏf�p@�>�������`��+ԡ�.g�5dLv]��*�/@:�p�~��^}aQ`*�]W�t�1���m����Z�`l�k��`GGb�Oct'w�I���{�Q��¹E�=�ߠ0L�=�cz��e�^8%JG�pߍΝۂ��L~�Om�)�9��*�eutuD��N��Ie=�v'��j���njoV*ys�����U�뎼�Ӓ4ݲ<�b{��v����WT�F���p6')�S�]5-n�	9��썟8�M2W���ц�U�)��G�.����~��ew�2��7i먮���?y�?�i�����Sѓ������Z{��UQ/i_dv�ʟM̜oCį��vӆ�^6rCˡ+�5�gԜUG��F��מU���"5#Pnv����B�,�C��Qۭ'P�ݫ�yp���z�z^�R�~�r��Jқ��=��r�J���G�WBJ]MVj���2P�I��ruc��
�}p,��`�ҷG��i��f�U��-��"�/�(�aC3;SWA�}gSUn�C��̵�奌Z�d���d ��/K�#u��YO9����ɋo`e�=J���ˎ�����H���QmG*E\^$��(ص�s"�,
7|�S���i��S�8�`�y""���a0n��]ڛfY�K96�]1����ɋ^1g �'!�u���p?�8�1B ��K�yb��o���c��\Oy֭��VbPT�7��Sv�El����Vb��u��]�]5�Ҹ��7t�x�[=Ԥ�X�W�P]X�jPB���B��k�V99�]amu��S��d|�3������tN�`bciikh�^�Y�KLOV�V�ֻ���]f���u�{��_7d���w�Yya�m���H�{I�g9�0��۹ا��U�E��y�oj�ʅQ/�$v;���j�s/��9N�V�:����ܩ���t�GVu�W�aa���v%(����O>啩Z�ݖ�զ%ԧ�*�k�Uo-h��.�]9���c�����n�]m_�s��T#5}X���$L�;ۣ��D��h��)H-�Cu���|Jt,�9뽩'p�����{;wUg-��U�b�����t�F�R�n�9�!}�§�,{��]�F�GMғ;��K�GW�����<�#m�Mz�*�;"�V�mrTN�1��ɑl�=\[�$;�ړM]dN��{���fM���75WoX'A�eVh�5uh�3�ι]�n=嘊�� �*A��l�V;��tλ��vn2��]-ۅVX�;�ِ@Wj����%��G���х����E��^��,'�ވ6i��^-<���鮕x*���ݹ����W;iGY�&pC�sS���{w�(m��Ȣ��ڕ�+����e[�e��ʮ�)���0�V'��F�,U�~L���i'�h$���>K�Smd۸ҥ��c�'{�r�,��p�KTI�\�:��Q�7������:��`���9r9�6J�������Y,I��f��u��x�Z8.�ֱ�U[Y���6]-�=)R0���N{�C�GZ�VWLu��W�;��5�KA:��M�Sr���E[λ�5q$�.]n��t�5��u���+�K�es7��0�\[�B�SY����x���-��Brs�L�o_�m�:�MEG�b�-t*YN��Ш��J�f�
5cq�\/��L]Fi{��o��i�j���͙N�����l�DHc�9�RQ��If2�`+��x��U��o6�j�V��ү+9�4�_ZKQhf���
�[S/��`��ᮄ��s���6� W� �s�:Q��7XȾ��-�m�o����t��5�=�`������1:��Y��b��Ӑ��i�C�w�����)N������ʺ�
g�ֆ�4� ��op5g�@��]�]]��T(���+K�c>�J��Ɔc9�R��2���)��k���.�z�t5|~��H��e���+�� ?���']��7��Ky|�!�2��UUяF��@iy��B������^��� ��}S+���+�0�>ȗ��������S�k����
���'�G��R�+���:�u����l��_�C�t:�2�8Rt�x�g�K8��t:���E{�nN�|�ͯk�<��T�K9Vi�̟Qں�����m�C.��4@�1���N��8p�sF��"`�V�]�:E"��=M3���+y�޾�[����1ò`�1f�j<=]����#�8��R���S^�w�c��bY�s�.�L���{�Ǫv7T�i�F(X}����4$��ȣ��@�e�u��*.N[���{9g�Ϙ�^��Q��|�Gn�/��"��׋��XٟA��;꽑Z���LT��B�VD��N�1-p�?���J�}�ӎw����5>����7s�;G��[�}��ݖE�D��W-���]S�T! c�?�KVn�~�^����Wn	!;����{3�ij��T���x��R;qm��9�E��bS%笧�(�)��h@�Z�Z��S�̬��ͨFfLSA��->�)�	��x8*Ṭ���9�;�if-�r���9%r�6̇��!�Q�_~땈J��N��t�[��'"��'ͼ����ұ���z�2N�������}�p�b�Y=p��4/�2 ʞF9M��Ȉ���tU6;��у�~ݚԭ������rF��ڪ�83�xda����8�햇������aHz������C���t+�dP(���6�t�j������r�s�}@�m�)�{uѸ�?iuի�0��.i�V�}`6�
�=oB·��/��E��@�|���`�9Y��v8��W����S휣ً�{�ԋ��;�3q&���jǖ��V�����F$V9�N����� �x9r��+"d�֫4l8�˜N}�z�M���?E��^u٫���2�{f�Ƞ�s��Y�E�P9��{nO��4����x��.u*Ɵ���;�f$Եn'\���dO�v�x�	0e򉫑�IL���_QR8��zq+�y7qz�����o@u��x:���R/#��| <5�n��$�S��c��w�n���
�{K�����,
 �{�T�A�*��!�cW��3��pQ�2��T�q���+}r�u�\TQ=��w:�u !T��1b��/��^c�C�z�dol��/7WR���E�3���;��Wh�uQލ�u��b*z�a)��ya ��U�)z`������^�צ18�<*&y�*����Y}sW�1j+Dc��k�`���歝�9MI��*���6�u�����V��+:q�VB���ʉR�o/�2��o��	���[uD0���M�W��o���x�r�ۿE�gD�X��ӥ}��oӒ��0��#��g34`f�	A��C�.���shE��k�G� b9X�}�".����ֆ�n�ʫ�c#�3�W����9�ډJE�I���40���&�3��*F�?��9�v�V������$�l=Y��1������٦'.����gI�t^n�����zu���Le.�X�3zE/S�|����S1��mmo!E�9#m�\]�fx.��,�ḩ��m�D�w.��z]��YW��A睊��o�1�@�H;^���6�n1
7�����%n�	�t���ޫR��|�g}�lx���|���MtPt�XͲ�>�+l��*=�RW(���ڛ�ck�v�۰���g}�1ߊ��^SU�^E�eN�=�ܫ�xU"���Υ����}�۵�j�}޷��˗�� ��V�j�iY��𩭍+�@KQ!Z�[�wqF��i^x��	]m��=Mz`�� ԨD_�9~��A���]�7�g����tN{��x2��&�*w����Y߾��� �W�h��6��ó��\;(����k}����;R�a�")k4��:��ЮF�N+�zpf�:o^�E4_��,�˔��^�a����>X�Ӗ���f�Αmd��=o�՘��W���꧹����1k;Q������5=�>��_f��%=��x��WG��;9�r����}��z/��2�.%�//�[d߶�B�.Ḡ0���4�ս���~�ڈno9� �L�W�C=JC���.�Z�JߌU��}����20�?�Fh��5oA�G^ZC��4�@���L{��}Yu<=�5 5h��X����_}I1rwJ��1u;V٘��Þ�v���9a���`�n���mt/c���6kz�F�T�D�g ��E�3����=EU	��-�[�^����S�83Ww�}�9�uq�D�#Z��:H�h�q�<���GT�8�z�g*f�uY���)P��%�y�ܬX��|�+�^�K�_��j�'���i�f�Rx�w���8��\��)ث��us�h�}�z�����k�.v{EΟ�\�pH�Y����/5&b�97DR�
WL�0^�
�̿c<�w�{V3��)��- Z�F��c�f�D����o0�t���}]ɛ�C�5���W[�ؼ�|ntV���;=.���&���%-�zJ/kS�%��L�۵��d���xv}ѣ��w����x�xm
D�̨4����R�T�oqsq�M���`�V�gd�]���0�HR�{��Q�J*-9���<zA퉜��u��kk��\<8hV��vl�fԒ�e�����������&%�����$rԾ���L9�]�w��;'��X5of���l
��E�?.�I�n��t�/o8|���)A�d\i�>��< ���Ke��k1f����rxۿ�nUŕ^��s�=m	jB�o��s1o��6�3'׼�����W�e�~�p��#�w�Ɩ�/%[G�.�w@���%Ҩg ��u���`�W�z��z���z���S�RN]zn(�?��q���Dυ{�j�Ef߼Sz'��]��wAJ��2��)��b����ү���p/VJ�P�y�� �v1e�5�>�|$ۡy�٪k�����]@��x`����O�I�lN�.�������3���� ��g�7�U.d��6�%��'Gc��ɪz���2/3!�Ms n:OM���:4tx�%;�N���!�[$Mz�O�V�,E�Q�*�`�7�������)�P?7���>wL���dY�5�u�^)�Vr��a�7s(8;�;.@^ϵw{C��}r��`�5��udL�/�z�bb�h2߱T�oo0o�Mx�8��f��wSP�4�����^����{�t4��{��7�a>���i�.���R��e�#�VkD���Ẹ:�U����R��F��>��⯫_?���ȳ���l�&��Dne���2�D�wB2�뾮�yػ��nd�IV�^҂��He]����D�o5Y��X&MqR�V��6<�����C�-��;=oᅊv��g����^����j}/����uKJj��>�{	]4n��e�
�(m񃔤=c����v똾�����sy�cW��Qc���{a���> �d��$�xf��J۠��펻ί
�y�e��}�G���\u�'<+����.ǵ���f��F���hn�{��6�`|xn�\�k����W{�囩[MF��o�mXS�ę��I e��W�au��l.p��7:��.�	��E�ݴB��*�~�x���>^��+R�:�$�b%'z�>��v=���g��vQ[�t"Vus5#ӋQ��%����@����D_-�{B��N�h�#w�2��!��}g���8�W[��ݻ��Ճ�&k�u{ܵp�R"�
���z��ᕪ�ʧ���|���b]ʞ��7�s��Զ$�L�M�EX]g-�-���M�ޓ.���O"�����DxѦfd�����OܼI��aΣ�Պ=1X��Z�]qqح���d�I�W�z���y��E�á=�I&���+�)��QP|�FP �k�j��U̥0�s��7Q8sʡC��3���Ѭ�8���hm��
Ƥ,Mά8��j5�,�$,�L̋!����i@�)�N�F�	���ø��������+���N��U�i���oT%�\���n���w����[B7���u�tp�.{���y���Q�!e���ea�r��,D��}T
����p�F��vh�=�H�)	�JF
��5�I�np�^>�
��Ѫ%w�N0������2�ir�����k-)�7�Ř��c�N�Hً���,�\��s�������θ��ຖs���{�>1�aމ��Z4/�g��ʸ��u5�����O�^�ə囐��I�ζ��O.�6�p>��\��O� t�}O.�����\}m�{���~�Am_=��I�'�=���Tu��u"l�^Y:�Dԯl��>��Oy*+��qBhͽ����M74f6(-m<��]6���n���z\^´���䎘4I��Ao���h�,���=U���>��1��.4{���T�{��23y���U������I��gݔ��e^
�[���a�1��c��{�������
�:B��e��:��Zc2��:�'��+}��lqyn��>�2��o�OC�y������I���3Mr�()�yl�U��#��c�bj�8�Q��.�V�(}��j�VH��<q��s�v蟇�M)챟	�(T����[���h·������ͤ�ߎ 5���Ep��9���f����X�#^�sΡ�VWu��/"�=vt!��$�3�K�WwPrH�]���O�'m ��1N����Y�`"F8#��]�ۺ}�G�<뽻4��_�4؟�g�}n���F����[�8�Ǻ� ���M��q{Ǎz���Q���y��i���� ."�N��,u\��:�|%uz�ͦ��EU�{��&]>��|^����2;��U�5Ҕ|蹏���\���0ś��,ָ���@~��"w3�Tb�=WJ ܜ!VzuL�n߰WƁ�P��(}���q8��_N;"˺�8�<e��}��z�<��=�q#FEϩ���s�t��e��B���	u
�C�Au�>#k�e��hܷU�ۓ	1zwBb�N�y�Ȭ��-��(�Y���%�Y��lI����QL�@�(�9�v��L�|���o�fϮ����P������tO��R#T$��Ye��mk(����[tx梨�U{Yܽib<�uv�ނ�G�q߫$S|m�|y�k�`�i(^�rdƪ��|�58����I���*1`�ok�}k1�e�jT��S�z�2��^�3���š�J�n��YTnf�g8%��Ø}���}$T�<N|�Ɵ�����a�ў��/M�z�k<�q��Μ��u\c -����
Y����)�tQ?Axo-G�Bx��y{zwH��]��o$˛#l�*��:@6��#a���wl���"l؃j��m��H{�n��)���k�ZjZT۠ˎ@���7�
0�}�|���}G����p����k��1��f��-<�u?� ��<tT��E�Y0�1���g�<+D�*�;�F���3��Y��7�ۓbY��}�A<F�Yq*�]�bFb��8~k�&��<xwD�=�>��9h��8�B���;�i�yT4��=v�o�T���/0�1��"]���8�+P�q�����=���61l+��8g�7�;��z��^�P�
%�>+뭭�����Z���7��	�kN:�(�׳���2���ϴ_�ts��#Y|ftC>��n+al)m����s�s���s�8O���ꪘ�"1'Ss�x������bQ��gMX7m]GJ�N�x-�n�>�0tv�l�t��xR�����sU'���įƩP�������y�=R}�]��u��g��l���`�Q�t:��خ����<k>�L{�&6-��~cӲ[�RFy��V^�w^��}��Wޥ���9��#=}sb=c���fWb��eޯkV�u����&�}7:�a�iV�����]TWF�ٌ���u�k~<x��b_�d-Գ!M�O��jجKh�B���������D�T�*Yg�ݱk���ЦTRC�uC>��v��F��&c���v���)��nl�<��p������2#2iV��5�!�'>���9�S�ւ��[�hѬۧS��c2fq�`�N>�,�����x��so�q^��%i,�?VZwJߟ�B�sY�`�'�<�V;wёV�cjI\��eeut9��oB�AW��k8T���{�����}�)$n�}��Fq�DH@<�*vv����V�+�NT����J�$L�\{տAC 7Jo�w}o��5^�w�V�/A�oN*���bh$�Op�7��x�-��}Y'#^�󺭱̏�M�&RA=�]F����	{L,�A�G��N�,�ȾT�_��*�/z܉��Z�����O�T����e�Q���WG,����vq�bu�%��5_+�O��.p�p9�Ch�<��|;�i�
�*+]fd�WT��r̥�yWUN���L�q���@Qޠ�Ypcv[�+�!v�V�LNwW��� c����>y�+qc�f2�q
�vPƓǽ�e����`�`̅X��D�;o8H��)��^'�r|���	��]y	e2���L^e����n�w_až�ǧ��1@�+՞uG���4��M":�TY�V��3��w9�vc�܃���ő���&p wNN�\JZ��
�ח»�ꦴ��t�����҅)�4����%wd.�B5T����U������/�yb�*:��5q��7��1��|�0�7P�7��W_3�x���]��ش9!��fب�#K��T"��#�޾GUYu�;�y4�S��=ʮ��w�G�ss�+|+m՗#]�-�l��V�nH�We����kT����V-N�-��q,"�Yǈɦ�kd�������:���jl+�X9�:n5����&�7�8cX&q�jJ��7O}Ǆk%\p
�v�3Ѕ���ggeꢗ
q��܀ㄘnr�����b���c�JU�
{wʝ�5�́-_c�N:(P��[�=mޟ�5�v+�q;��M_s��&dC\���!�W%nr}���ik�{+�'�W�<��]+Ҵ��+VznV%�2�Qaǽ��sn��)�Qgz;Bε���Nglv��@Tڭ��iTW9u�ᤗe�Zū㴰*B�%\�]�R�$Q�f���3��:�[���٪*B��wS�"Kh��ƥ��C�4��U�Kا�����Ƭ
�{Ћݶ�
���R�Ԗq�M|΄�l�x?:�2�
��H�|hWb�T� �r�6яk5���P��ͫA�L;�b�����9d@D��ݪϹ�������@�$+B���j�H-cmT��oK	�2S绅ۭ@�CB�D��T�mA\�V��gN-��5n	�f`��]�]��̗��<�X�p����-2:�n�!һ�&�p�����	Z��$��gg��W��m( �O_h��ks������nR8�s�&�\�t�6�H�Fr@��'u*Øv�Rw6�J�M;Ϸ�g�*M���a��:�Zڂ�<= �S��:ۂR��Ò�L�P��_"3Z܅���į�6I�O~�z�*����)�T�\�Ұ2�vbh�m1;����2�<��t��wyk�8b�$[vTYOi�gR�o
z��WM�.�x	��%X�Ն��/����1���]Q��IR6;{�;��
�f���F*�����i�*b�n�&R�(�r�n�8�ƻ����Õ7x���'ؾ�x���#q.6�6Ь${���N2��/�`r�*]�d9��ɻ�r	���yf��&J�_2Èݰ��ʍJ�h��Utv���@���!������>Ȫ��`��^9o�X��ó8�+w,N�����P��.��#(a����tS�(���=��&��t��r��K�6���z�� ���I�����Pdհ��;6Rዮ��̓c���Ĵr�.#TGY�@�}e/
e�:K=eNi;��Nɰ%���4^���\��b����Tʽ�SZ6�ԋ����l������ur5�R��N��!�ޱjzo�v���M����*�CC!������u6[��SH+|��'c'T*.����#��IP�*�2�R��ʡ��5��n�Ka�	w�qt�(�o�̰�9ɱ��5�5����wr,�W ̹�s���k���&�p�߿Uyg��o9��ɸ���j���1{�JuN��mi;�]��$X{L"���qo1E�\o�w%�V^NJH ��Ҙ9�s�ǪY�t����>+���Oe9����9��١�a��*.Z�Z#��/'9�鎒�[3��~��0q'���NU/M)��9�ؙh�~&�|�ΟjK����ٯ̚���Y�9�B��g.�I�7Ы����o3�D�}�Qun�>h�f\zq79:��l�g}O#Bg6eY��n�2t�À/V6"�w'##.ޣ^�Z��:�5��?VٹY�#�^�����LRv�P�2��*�H�W1��xϑ�)�Nr%�\�Ӏ#�]��>��E�U�&��R�l'���0�4E���X��%�� !�=e9�9�V �=�#vGt���i���b�z�UO.��E�M*x{�P�_��e{m�6�@#x�����oX�m�y[�X:sw<����A����횐�c�o��ÏVr��M�I��K-�u��ڻ9#U��н�����#s��NN0�oZ�ޏOX�y�J6�7k]W���߂�:h�L��g���*�=�]T-�b`m]���Dh�Y��j���6yǅ�^���)�]��{'7����?u��$��O1=E`Z��V��Vh�亵q����-f�T��{y1����S(�cAlޣ)������t-H(]���u8�j�<��ts��Q��v��Rc\���yP_ubV��Q�=��h�?'e�]�Gfqd���,{=/Ԫ�Uo��O§�عk�f���ڣ2'��Z�^K�3��&\]L�����~N��݋��*vM��UiC�}��
}s#�Sq��ު܀��;�U�c�ݨQrg�,8�JRy;O�1���t%쒽�=��{f��jG� �����E3DL���y��X��c��n�5�*y#��#�s�E�D��׫�N�^��*���E�#{{���jnqMS���F�3�����>��k����WP�j�u3��)��٥��kqfׅ*��`܁K+�� ?Ew�*���m����U�n�\�c�[�-�:�@6r��cGɍ	�S*Go���^��YL���>�y�nU����3�^{g��Wo�sO�=�K��L���
�n/ Ң$x�3������㗦�z/a`���`�WM��n���pw�˱i��ȷkZ��3��o�(�X&U�/�vI��?�	�Xw�������6�
�$V_
˨,��(�7H�������X� X�}�c)�2S�J�VfD�*3�'��vV��H��w�;��S=���3���c ���q՛��)���ʴh�Tm��o'��+ ��d�WaU?)�A,+ �w�ٝ|��7�q�ilT%5�pnV1Z��j��V�nFU�b���v%Ǥ)���\���7���r�"�tc��})t���xm��ׄ܏�q����Q�+��h����&�����,��{�B+ܣ2�gfO.�a|��	�Ԏp�%�s��f�v./�<�5�zG���c��z↔�bB>�#z�o���7U��c	*��i8�1�n��3]gg�b���̱(g����L\t�W���/�o��t)Tz����k��pħ�\��V��o_ޘ�����T5�nK�ԗ0a�:��⸑���_�eN��u�����}��Uv<�fS���g���ﾓSJ�cײ�u݁3Ą���ќ{z��rl��Pb����dȾ]m��ڹ�,D�L��Qս0��v���]ʓ][;��YQ�ڝ�Z:�ϛ��T_�Ư��X��1U���Z=�M!=�N��.|��ɊW�̕pF���s��s�U?z{/}���G�@r�-u����UA��&
���r�A���>����ճ����W� �zTİ8!���:@�co�31:9Ъ��8�VJ�څ����ުT��	ȕ(�t��߇ugԸ��:�I�bf�X�B��o[�W7 �+�ugUos1P`Tj>?Jۘ�#ڲ�P���;!l����sE1.���7�\�Y@�\�s�՟!�[u��7Ȥ��Ǵ,�9��{ۻD�j���?G|V"Wʂ9+��Z��+z2Po��dm�DF���L�5g,)mw;'U���_wR.� 1}�gW'n�]��[����`��?Q�Ɵ��s��ڼ1�e���q^j�����fF{��?�C-]�z���B_c\)s���:�`żǏ�d�x;׆lX�n��;{����.��C�"N	<�&ϱ����f��4��P1SU��cv*���[��I5c�b8������4��U
�F��:>��&�2��ھ9{�V�w__�K���ҭ�r�Ex��_	wƳ9^�d�3�n�yw�ˮ�*J�=�h���s��N��P��^'�Y߇ ���N�)e�#�)7$)؉��7-�����N$8��W6�o���ӽ9�e3H�b���.o�_�4��:c#�߈��t��\�ڀ|D���B3���V��k����$#���Ӱ���X�+�A����)�^�/ݤӎ��Wl�1,�p�}�����#�E4cD�~��F՗�g��vf�C�{^�Ӧ}�r5J(/5���i��Zʉ�x�3
zG5r\t	Mz��qC�N��U���y,��`)�sÚ"MD�%bެ��q�46���1y��,xM{���{.��M�g8�&�ڳN�|���ʃ�,p�훴�7��/��La�v�	�D�d0)WGe[�@`����uF�3'~�]ȬQ�X�3�6;|�ʶ����ua��t���-�lօXk����B�w���o���������,m�\�Ⱦk�N�l�����'�X~	�`B�n����������<���E�jÁ]��Ϻm�O����}Jp<v�t��ݒ��y��V�/T��MK(D�%E2t�i��Pn�3�C��w�QC������&�秙�RP�nqN:��eyQ)�M���s�ǿ^	(T�$v�������(8ܢ�5��&d���S#�8��!Gv��X��{zL�o'G?Tt�z�R�d�p=�ɬ�ĳup�7V~��1���������5׮$v���b<����*a�n�ɟn��t�7�|��n��qL�����t�ߊ|�xv7�<�u�nHP��0�{�,Lx�I�SҷLW�b��7\-�r`�P��[��U�罓�Jn�ڗ{}X���G��T�糲��X,��*�}����F�?�S�+���Uw����3ڜ�Ӝ���8�eTߗ*~���,cH���;�l�Phx>qG�罴�ˡX�BSOF��e�e:��\�E0=\��C1�F��F�ｗޓ�C�����aø������������Ӎ�$��d����ݤ9���]�:�n%V��k�&\1�(�#B���J�%J~	#��DP7��综�.Auٽ6��zѲC��5,4]v�V�܂nD��*: ��t�WD>`Lںƪ�v¯N���펵��D�1�ϬX(#�9Uw{�v�P��!��~zǢ�*=wK����Gr��.V�������d�1,tq>��|��a�R�M�U{�%���3~��^Lpe�x�d/*�ݺ[W�ܹ�3�ʍ�07���?B��W�����0�ʝˬ�bB;��M�*�c:@�zeNW!k�n���\:�7�:�QѮM�]S�|l�Izt+�v+=�b�
	�Ѿ���%��M���B�51�����d��wh�q���1*:���k���zRg�eZϦ���P�3nyc���M��H�![dR����;sB��p��ڪ
R�jg1����صL�|o��M�[Z�������3S0;���!٥�������v<ec�E=��C2^9��ue����(nBP��������{3�b|�������뉫�K�)�@�D��~�o9�]��-�P* �5�)��i����s}���C@�>+��nO�U�6��p�I�[�k���$��0�+LI�����=?bp�)_��9t����`��w+�4���/��`�C���_G�^C��FHSR�7����m���_b��ł�=Ƕ����_q�L�MFӸ�XAc�A[�.�[��n���^]>R�b2�y�Zj�)fXˊ�/���Smҽ�g?��S����Cc��'�So�jեm��ѧy��E)6'�z���r M����7�S��km8��ܩ}3�ٵ~=�F8�8w��Lt>P,qԳL%�woַ�'��Gq��pݕu˞���y���+� F��8ʬ�£���4ϡ*�/���%�گ���XJI���Ã=��9�s�f���E쨗-�����F�b� ���Un6q�<�F�,�f�G�؉����n��a�>��rOS~�{�w�%�dǪTPO:0�����OĀ/Q�������h+رOu�����`�Z�şr�d������;�!цϘ����ٔ
и7��f�R=cV�=Evן&��G"{���k<ǫ|w�O�`�� �|�^h�鋓r�:�5��k��Y���n���/�j�U���w�W�"�F7N�j;4j�R���>J۝�I�zn*�$,�u�JR>�Y7��������=򧘾ѾZ�|}ۂ��DNFM;)/LY��|q�8�	��;I��54-�tM er�{����i��k>9�~$۫W�E�ؽ����0��7�@��{mOE%��������31�C���^�B=����ڶj9^��WyXz/e�Ѷ.��Xo]��8�5�t��۝�j��p�F�%���a�]�l�jq��xޠ�W��ͮJ��0d��Z�9-�_N��Y�9��Z4��}��+<�co�[�Auj��T4J�J�϶ɡ�P��3���\���'��`��E�_��Q��Q��_@V��@E�yʓ�gdL�Խ�nZ�U�9}�^�]�g�(U1W�\6_}֡\';#0Μ�ҽ����VK;C)�fP�m1Ʌ�0k��$���	lwH���j}�����&�:�w)l�&wo���Y;����|�]5p�[���9"o2�w���=��
���������w`�=�Z̙v��O���j4����Rc%w�׶0ʤz�\t�������[��\�{8S��2c��S]굟���}ګn�N�l
�w��Äyki����=n� P�|e�^��"��zWoZ�YQ��=��������Hy
�?��^��'��_lS�w'޼EP����K|��&�#hm]8B.��@��G��-��=%���׆��j&/��e���O4��ZP���� ��4�}�a�vzrOKY�Y�h#U�b��aЮ;ҡ��E�y偰)H^��P���N7�:|{0�Ѹ�~='2q�U��R~+��O�ٮ��᪪�uv�zV��F�dP�,W>:Nm�HuaG�ө-����G�u����웱^��X����s�B��%��V��1�~�f��{¹|_�vm*�m���|�ъ��]fJ7յ�̰q�Q�����.4W/+#���b�wc���	d�_�f�)��[��/��ݖQ�pD��"+U���ɬ����K'K]Dx�\�����pb��w[]:���ቋ�/<n��M}<Ԧ��Kй>+ӌi��{^&h�}�֟�ovT�yu۸>i��k�eɉV��*j���OfѶ�i%����˧��Ԡ��i�K�ek���GśM�@~����q�����6���~Ȥm�k/�uf�U��rjdt�����S�|���4e|_��f����NS<p����!���b"�m�s�ԕ9���!L9��5ls��ˆ���%��=5�R}��w���ʁ.4v��w��z�N����PX�Y�zp��G�o�>c�g�^'Ȟ�����G��}&�}&\��HT1�GҎ��]f�-��`롳lZ�0��"v��v2�^�1�+�3ðL�in%���`W���-�43,�LUm\�o�D���]I�^�l����"���(fx�꺱W��N�:�K)�'̄�ݳ�*�}�����_y�˖G�c*g5�)+T�rq�~�P=41q�њ�}ڽ^���(C�걲D^z����x734���K�=��z�W]�խ��|��G����)V��Dlz���W�n���i���.Y�w���gt���ݹ�c���u}�L̩6d�x8��hwm�]�](� Kz�V�=�@+(�v�ԟP�:��E)��y���6��Λ�,��i�WKC�nwd#b�4VSW��ܩ�ZZp�1�\u�ɿ��
mv>��-�B7cwfط6��s�un�e�c��z��F�y�6�!ժ�R��Jv#<T��j���j���tmMw��݇��{�g����"���	)Q����rp;,�ڄ/����~7����(Й�@Lo�~��f˂"$GEէY��뻇t{_���څ��Vpگ{\l4�-]2��F.�'�e��9D`l�Ժ�u�&���t}�~C��,�'�b��qd��h�^4�/CӮ��oG��w��V�#�����Cr����ldfL���f�a�o,mw�W.K��CQ�뾨
b��>Tn�Yc1&A��#��*�K��V+{�{�_0>=��ү'r�i���Kc _�5X_^�����8��mLV�Nˆ�c:�_T����(�*,Dں�b�f}J{Q�H�x��𰶢d8u)��Q��=��j�;�X��n���k���u����?(�Q��
��<U������A�<�x���VvT��q��;XDI`��8T3���~d�J��Lz��"D�wX�|S�=����"y`�lmw'��g=}O̓����'��'����;A�Gֈ��!b����O	9J��I����p݇����ެ��ʨ�#� �Q7�.�A���Ŧ� -�N���:�4��}�ܝn�T��UG������,
���Q+=j�6U����O�f���Eq����l�O��	nf��6�������Z@M�OoQn<�W)��oZ����+WA	�,�P�U۽Y��/��O4�ݫz����N��4uM�P�Ի��c�:#n���NĢq�mGW�y$�sh��]�H�:����YӨ��'||{�+����ꬔ	O�0d6�W*J[����+g���H��R���7�Ʊ��������Ζ�
�w�%���xdi�Z\�	{��5;hldAm:�]����oF%j}�w1�����zG�5�w��J[ytxlN��������W�
F�y0e%ݑ�M��(�z�������w;�,.���"-u�'⹫u���o�j�j���|�=:��������]�47�J�p����`�D����`U�Ap۽[��V�%lF�(�sU�Շ�WmuGg0�Z���N��i�,��Ș�oon�s�ݚ�ëk3�N.��'��ݗ�S�_U����wR֦��Wr��M�x�}f��z��<�B���ƻn���ݱ���ޮlϚI�O�z�p,[�v0�*�PY��a��u��ͽ�:,�]���פ�'b�ۇ����tO14Q�Ѭֶ���îgZ�qf�AwKL���l�{~
췊<2�e��$�y��ηv�T��G�I��H�s����u��8�H�I�G_4��o��Q�F|G�p�#�$��l�����s�SU�A��.�A1�Ew_@��b9�ЗO9�j�"0�U���ޭ��d;�}u����"`���9�Z(�kfH�4��]p���^��~�*�7���w;s�Kx�
��Z��t��1"n����m���2�Wr�+�e�7��T1f�ˑg�"\�^���Sz5�p���=v��c������#s�t�Ǯ�3���j�З��~�]�-�^n�fLT �v,]t[�JK��PW�/>��\�{7D�
9�+�VQ�����`�(��u*GM_v�2���o�D����b���{E<����T�S{t���������y!��x����: �]+	�:$��ٸ��<����1�s�`Ww�%0�]}!x:�(�ՇH\�fNK\:�IYX���'��Pa�C�F�-Ҭ�������e�9����XU&6N�W������.fA�;��'Mj�z�V(Y\/m=\�{:�Sp�f��xr���������e�.��_6ĺ	<|�jq	�?�n>��VuM�j�u�ЗE.˚0��}.v�m�;�n//%(	߽���;J�X�F�Z�5{�:��=|�r��
U����	����A[�ܶÜ��Yu���m[`����la��	�-�l	��	֬qn����>�{=���9 �F91�)�	�u��"�wQ�T�L�A����ɝ&#E��Ao<L�^��W\�Af��;���^�ۡV�P۰{�T� ˋ>\@s޹De-�r7t�OxH�[�(P����e�(�#�S�a|:b��P���t��7 ��5ۯ���-ڷk̠�_V{���ϡ�xi�>I�b~U�S��}������b��7{�2&rD��O�Z��,>�+`���2�N�oy���H�aR۽���z8{R��ezLl��-�g�����w�C$6G׳v^��i�����/1+>e��Ґu�YQ�Wt �N��Es{!X95��D�th�3�a��՜l��U��$W��=��ڶ�١�����-ej)B	������`�\�υ��=�M��AП�͎>])�u��^o�'��j�9f�h�2D��x�ݍ�d��̻U�/X�h���잭�ҥ�2��
=q�FB���;��ʎ]|�>���:�{�����{ck�O[g�Ш}G�W��/RZ$,½���n����,z���Ǹ��e�|ي~�%a���SC���:�d�G*��2��P��)^i{5\���yǇ�}�Iꋾ���&��ƒ�	����IE��~� ���'ك�rX��2�;���c�>���Y�k8�ռ���AQ�Z��a�<X�a��[�U��of\Y�^nSh�Pc��s9k_$��޷٤�lf���fS<����Q>�7a��\�o{��u���7��ʳN�٥ˑ�*��r^Eq�-����:
�Oyo�pڢۦZ�ۑC���NpN&�vUc?���]�x3٪J��4DRD��
"2����<����-��
կx����Aܡ$�2��^�4ȐU�,{��X�R�Z���}��JڇC�٘9�P6K16��z���lUM
ʄ.�wh�yR(���ٽc��1x�y�A^m���3�{���m�"�&0�X:����tl�lz�b����d7����ʣ+�������T=�{�9�_]��?{)���BL��x��=�F�N��3���z��{�\��\`W�����3�d�����Q�F�54����(���nm�Lth��� JU��K�A�t����}�B�/hۗ]�݉�q��.���r&��41�sʕ�lr�F�}����sƆd�]1��������	I9Q&�i�R��C���c���l�~�{ �>�!���֤�o�g�/6{�/�v�,;���)���+R#}�f����'��Uz��r:����F�᮷ǆ�I��g3�t��֩�a����|S-x�T�0vt�H�#\m,1t����ǲ��@��w�@<e���1�P�����8�<.�Vv�R��Af�@Sq0f��o]g֖� �ü��;��\\(G��E��Gc�dƺF�Q�|����{�%J��u1�.��}6�:&rn�qC$<Z�>�ވS�Sy�Mr=C��>�W��È��W�uL磸x4��K���'��r0.���:���;����Q�a:ߥT�}�SÙ��V�%�R�m�����^������un�\{��ܵ��KP;��ְ�|`�G�s(ѧZ�?��՗C�hn!eKy:}�^��o�����/�-'�FK�5�ب~���޶����x��V���R�0(n�D[�D�ɗ�񑳺/Zv�-3Nq��[9���j%�S5�k���"��Q��ۨݽK6�b�w��m{֨s9��F��)�~�iG�v��..~�K�p7���N�fi.�.�Lb���U�("|���sk�{��p�re�`������e���]v:n��B]c˄���ҎF�O�W	��7�w��=�:rh�5�4��xG��<��b�E+�� ��^�{�;��]�a=�*���v��fY �^��H7���n	�y�D�>,�G{��;Y�!�t�\Cs���x���,g�7��tV�Yh��S�0��zyz�R!��-С����� �˺�3u�=����#��d�gR���y��k�;��r��׳JV-g46��l7�q(H�ju1)��·��W�;�rۭ�a��Xɝ'MpW�=y/PW9糯`�ྫྷYl:n�v�+�ۣ؆T��Օ�WJ4G����7���Fr,ֻ	N+���
&�[����t���9-�J\{]yW���'��MC��yB��O���ѣ�F�Z���_�f��¦ڡ�g����f��lļ�t�Ym�\����'�\�W���@���v`��}[ab�gԣ�<��Ʋ%>/q��ZZ6�^�n-EX�w���_ ��W��`c����j�m��]
c^c ��v�����6�U���j�7}-�C�EFқ��｣�=x�ўҰ�[a�
l����?P4mp����!r�,>���*�#��vX6�I��C˹O����9[n�U9�j�*;J��p�*��P�;1֦m3#p�8�	�̻o;�N��5��/�ꦉ���T�{/�مG�c��}Hy��4��`��;'���d5'���Ro��
�A�����>෼`.Ó�V��'ӧ��c���pJ݌ ���zatg�.0U���c_n�L#f�s�n����L��-���w_٭b'j�0��z"�ɯq���Q�r�Y$����2�QR�c%p��L��	j4Ų3�[�j&��E��7X��p��gJ�������h��?0R9��+'I�lI�W
�B�2��� �f���.�0��1(�����;ib�y������Ĥ�I��WC�p���� ���wy��pi�"ח�(t���5�n����Yxƿ/��x�rʭ�=K����y�0a�[�9OSW��uj@���2�����W��<��q��D�p��� i�x�SѳU6 Y�/����3����X�^��n��39̜҇������:t^��ߪ���ؓ� ��d��L:'�||A������h�N�j|�,Ɍ��7��^@��>�Z��Q�2yè����phZ�:7�Z�cP�G뵅ѩ>��N6�J�
����ճ��lR����#��r{�"�q�}6�*}0�:�0�bL����_��J��+�b�O�^��57�Vj��b*�Pē��u[�>��p��[�j}ٗ켞8j�c��ꑜ���R��h�&��U�r�f����%��7���n�S4/,���6�s)���n���Z��H>7k�*sh�C��6l����=0����]��,�6�G93~��o{ѫ�T��w�Ԟ���j��A�=�ߊ��_e6r�辻Iz�B���}�k�'=�w��|�s�nk9��,�ߊ�V/||R��*��把4������	L�/q�f5�K�S`�Z����ݼ�鎚������ �+j �|5D�Vy8��ecg8�6 �u����k�z7,e��g��/o�x���E�^tj�Tx:Ź����,�;�4��l�ǘ��U+ �f�;1Y�9M靈�_H$�.��w^�1}�j�$D����Z#1��m��#ue�Y���x�=��l括f;�E@�;���H��-%Oo���-��>#�]� J]��F�)�ɚ�,��K���T.ֽ\M����F���J���PZ��(:㺽^�Ed�}�����"��z�o�/��nL����꾃6�_�Y�L��b]�y����u�]���)��E��r�J̛t�ş^�m���Z��U�,%QIF.1۝��`y��9(��c�� ]�̼TP��v���Q��0�o���z��y�-2|�l�ܼZ��ǭ9�}�Y�S�C�Cg��opā�Fg�~�ꮣ~�����!��F�pUy@�<�\��r�D�l Ĺb5w���Pz��[��R\�r��'S�	5V�	dI���2hz�F�Ϊ�C0U�n�$ch8��W�zji��p�uVr׋s}����x�3Pb��{Q#&�uu@�I�h=��DnaSnWx#�퍿n{�r~�=��z�������񿅶�H3��p�ץL3�s;�/Uq�1���8j�k�~���[Wk"���2e��W�}B���91+Z���+�3y�+-
K�'�jB����n����±�䖃Gzފ*K쭗�2��&�܃Cy5��꛼��}�$��魶��f����Z�B�9.xw�wh�G��| �pl@:]W�x�Z��$;}�D�����f��>��x�
���w�tܰKٽW-\ێf}�=R�G�ca�L�&�y�Ι�͛���S��f�8W/L9'��GH~jTh~��ic�Oٓ֠tgV���Z����No2+Л�a��yI�}8_Nsʋ��aOdޘC���������mQh�vw?F�1�v�����=��!1b�qEs4)��f��V���i;{Q���s:y�G�K���������W7�b�ǌn�f	���'a���*�*�5T8G����N�[ۀވ:����j�y���*�����.0_x��f���ZzY�u�u��:�c��*��wݣ��@�P=W�p7�yT(��8�^�v
����"ۺ���%��.5@c�z�ʛ��e�Ą_���s��gg�[W�Z/�����,��&\p�iF��3��}Cee_a�'vaX����Y�Ŝ�y&�X�vj+G��Jm��Yvlf;�/b5� ���}�H]��~�i9s,�u-+�cdw���I������w����scc+��3+����Z�u���n�7�bc!���1~�&�T%��	������P���V^�_h`8��ɶ;���Pӡ���@���2��(�~��o4��v�-������ �κ
�.X��CC��1���,��TTd�}G��C؜�ͭ��#�ǁV|�U�{;W>JI2��;:}_\>��U��SU � O__��8<��:O���V~N�����󍉁���`u
8�֬N.�"���'sZhK�����n�oo�6С���+�0�B<�Z��_�8�GУ"A�϶+��-�.����!�d׽��ӽ��Ө*_f]>|�� 9�8t:��I"��5����j����߻��$W��C�[t�G�S��"�ڕG���G:x��^z�ѡ��eJ�67jҵ�$Ⱦ�W��\[�-�rw}�S�r��O;ι#�y��
�1�(_�+#�8��mS�#���Fǻ�ŞÇ�_����M��n�Ygf�S¨�X������n"�&��Ǣ��&F�d�%)j��u�p@VI����ٛ4�&�����v#��^>�L]%VͣC���Hn=�R@ß;�G��m�'ka�e�:D��Q�CY�Y�$ �`�uV�v��x�K�|}�Ex|z�����������[ft�ýk�_�W�)~��XbX9�n�3^4�8��ﯩ1�Y��A�&o4O^��X)�#�g@�yX��Ґ ��r����آ����"F��՚�4Pù���lt�����5�ˣ>�������:X@���2�_n��H����x�Eo`[���Ź��&��8�wX�U˷�#osJ�5��h��@�Uׂޏ;���3�-U҆s��/G�ݒK����^d�T�x-�צ@��)��B�����{i���;�z���fn����^w�ÆF����t�> z���X-�i����̍����(v^��e�捙��W��E�jgUM������x�^�J��υ#����{w�6}�w+���Q�|i3���գ�<s�.���c�!�.�����k��}B�{�)�J�\��,g`ez���@�2�Lc�t��p�=x*��C>�*��"���t��q�+�ꟍ����n'nj�"�tT�]���Pb����K��l����4��Fc��01�w����Jƣ��y��Z�Grk�Wm-/Iڵ�2\���z0�� ����F�F*�F;���s�{5�]��z������QSb��*^j��z�UPPx������n�@fN%ľ���4�.��E�����@4,�.���o���<�c�q���u�O�����vW���{T[�y��N]���\��P<�b^��
��p�<���ֶ�f Q�g�{�^e�fiP�a5t�ۓ���U'Y��N�po�-��_t�:��:ֈY��y9��A��U�F���kֺ���S9�΋�z��j���j>X�Ăd�O�u؁�}�c��7����w�$��������e�_�mFخfNc��Uk�;D�J��%J�����{~�}���7����*�O���9§4.o5ϡ���5^����".����oNk�a�g�v6%��aet8�'n_o\&1H�սLdd�n`m�T{/=��kZ��^R^٫��{Ҋ^����͑�LO����[<�b^��ث+���x*�| ��Ĝ�I�~U�R����4R���Z��G�3�)i��V�!�S�>*��X�a	�%G�ѽ�;���|U�7ǰ،�E��"�ۻ3��wm񍛎N�Y���8��9ʲ��ѩgO����]u:4u�u�W(��С4���'����.�oվ=UV��5K������ps�>����#׋�����5����9�1�\���\�mW���~�[0��g�ѤXTN��SJ��c��M��v����+��X~d_�p4k��Z̕�&����	E���ue]���"�mNo�7D�&md]J2 �1+�\�DI.�7\s��?_ˤX�i�Q���ˮ�~���V֭��>��(�Y�xԘ6Y���*�]�kzs5�ҧ����e�{ҰY�z�d�ŭ]M��UE�8j�ŕ+̙�>9��S}�S�ޫ]]����I�R�P�3s�k���M,��/���	�g��=�;�:��SW{te���%�tsC����wvM/<"�A�,�`�{��7�9��X|`a���`��S�r���+{6�:�V%�&sJ���g6���}v����F�fj<��#�:���v�G���vI`�Ʋ���<�7�_t���bK��wIo]�{O��k%֓[��$F������c�ZΦv�q�i���x�Ԛ��X���ð@u�\�������K����Wqכ�]Ĵҗ�}�_G�޾�a��#�0L��m�ۭܬ}���Ԣ����S�Rt�9�E�4q�(��v�_Ѓ�+>�N���]Ҧ��J&̏��p�X!R���j��	�J�2����7v�F��԰##�Ҫ���S�a�y�]"���f-̭]{,�v	�Np*n�ө�mN՝��.�4�k��/C&	��z����ڛt]�w�?V.�<�Wqv�F�p�:\�y��.��eq��_r�T��yf��S_m.��l�v�rgf5u�+C5�.$��]v���o7B�)!�f�R�YGO$֦��ʰ[�Y�1�e�}�+��٧�����jrt�X�����U��kC��Y�c�VI���2��Z�ǖ��+U7�v��9�6�o;6l<T1š�{�)qP����5boS{���q���UHr"T�%�Ky�oGO�SQ�1ү�d�\�G�6�m�)�;�Ǝô�TA�e-n��v̀$aq#������܎�D�V��ד6��4��Õ۫����NI���t�Hpj}f�˝�vY 5�mwAֶ@�Ig�R�f�K�Ep�1gՕx$hHL_�u2��G�Fn�X^�Ƿ�5O\5�je[y[�F�#~�n�m�_F���,��BѼ����M���9�)��
�34�79Z�at����Π�*��K���ݶ����Pjq���0V�$u�ͮҮ�5.�˧H��8w�)�l��vV���U·wn�Zm�2~�x��YԗGY���7Mi��d��� e�_2��=z�nq�I��^�7:ļ2��j緢Tsm_�;���F.ږ���x5;�{q�j�u9��v>��}f�˥{��l�{�h�̕��^�<:��Vn�Lb��c��jm�᮹v_\u�����We5	�M����d�H����DS]�o�"�Gzte�-�Ȉ}NW\թW
h�i�Op���N�8;d �H*�ܻ��)ΚE�pو�UH�w��`;�j���mv�����]�#w\?m���2��Mp����2T�f�N
:��{!��9U��-�ѫ�]�}�����L��KK�vV-�o��b�
ں}ѯ�1d�K�a�gOS?*#�9�;\)źT*)]P����&���r�eD��WIu�s�,��{I�W3sT����T"#��Dsk_��gv�ۮ����+��sa�ngN�j������|��\E�j#�;=?��:����s�e��5pO{0|�l�d�5�+������d�3�1]K��_n�F�ݣsz$�8�s�E<��O��Ziƃ�	�r���j�nyc>�/F��͆�_8{��a��1��d���ne_���\��+�������r�0Ts�RkT���}@3�zY������0(����������z�M
��0�e���6��G!W�0�EL�G( ��Y���oCqh�F�.��R.c��°� .6���/F
�x\��`�Uwvrq8�F~��fk�beƴ�zh���US��ڃD.A��y=Q��}oUA�8���d�[81O_��V��U����Hj�������l�v�On�[��yVy�s���q0о7��ŭ'{/�����5�j���	V�D�U�n��z�z��<�/G�VN�򚧲�}{���J���؆��}�Gh	�� �:ϰ�����q��z₆���|0h���ɋ���u�{��E�^G�[�J��E9�)�.(�g]zX�[@B~��	ﭨ�<y��䪔�]�ܟ8��tk����W��u�A����g�%\ �o(]�*e}��i��}�[n�����	��싦�?K��YWs���rR�K���wױ�)7�؍�͍��V��5�˚�<NaLĴ�T;1���f@�E���@�62�v�C���x*^������:f`j��sGJ!Q�wKcx���'Y���醙��� �ڄQ�^�4�m������d���[5Uw ��B�.e�㼞J�K�碮^��f�<��6kw���2�$C����τ��E�ι۰�hx�������V��'�ӈ�XbydqjFz,�1|�j�Σ&�Ujh�w�2̺c��ذf:�K����-n�4�� kOþ�EuC�vqq��a{_ ����x��^��N�d�%��<�deAGX�V�7�����'Z�*0z=�:#�oe�Wc�sc� X����s�s�TpY�(��q�B�&I���Ɩ��3�n�7�Z�o�/4�%&k T~�mt\u`�]�&�݉њ�g��y&c�ŷ0���t���v���N�C���.��O�F�4� .��9ψ���v�7��="��_���U�� ����a�nC�~u~5�GE�%n��lK�T�o�m�CWc�a���� �ӡ��@���oL\��gh��+r������G�=��V*%K9S�X�����"M�t�w{��\��\ ��c�^�xu	���h��$��19��.���W`����b�9]��p�'��鲧��SE�K���/ދ��&M�Z1�%���J�ŭ��R���w]j����
�3�<�Ly]N���j2��i���Kېo<��B��|���N_�s�$���z5ۏeۘ]�Ӽ�y�b�_b�s��]��.l�YI\,���"�Yٱ接k����s�����ee��$��{g��_&�u�J����|<緫"�1�y]�OF}�o����X-����2d��=];��3:�o���V�<}�쇦�b�x�l������Xs\ L���`��xϳ�;e��R	Td`�v돐X=�M���z���*d̷A�t�n�w�����C�w;�Sy~�o�S�hEa51:gO;���ژ������ԋp��B��0s�j*� L]d�y��[2� �0���۾!�5޴�ob�
�)�7�4y���$����c=�@�����5ݮa��h�^��!��C��:�N	��O���r:��x��3S]�g�����f��B��OFR���=o4\ ���a�7��xT�:��{��7�3�I�_31#�>��w�{{�1�u��"<����#��W�{k�ƽ+����,�OǝTi�7�@'�u����©��~V\cc3�5)@�0���W�q]R%���`���S�`�=�~{u�{w��VZ�ԭZ���"�f�7"�3�X���2{�k8�/�1:�A��Nѽ�p7�.�)M�!u�W."hAU��r��Vv�A[M6c�T|�3��.T��A�A��������R.�B�Âb���1p(��خ��G�fԭ[w���\�A!�,����,�}�v�Q!:�p��7�2���z646qe�'g;�-��,'�`�#�c�T���ؖ�^vw8}=y��C2�OkxK���F���]�6l�v���hɆ�7Vm�۫��~��)jI���>�W�|��3�4�|� �z��������ŕ� p��&�7�+[��dV�,�
.�c�hs3jC�Cɥ=`-$&\�]{Y?Wsg�ůz��)�n�Wy��������sHE�E�3?#�������Wl�5�����p�5z/���4� |7��w��+����|���x�;�ԋ�:���_ b�,�mCD)i���V��uem0�u���W�T[�/l�4B��ӣ�x���{����Pk.�4�F�U���zҚ��*�@"�u���56�ہ�f��B1�H���0��Y�NHf'ڮ%��7�K.gMލalk�ݵ@ST�oN�g |0z/�!k�ީ_L��{�'@N�]�C)���`nB�Mx���*~"7}��3��Z��FIf��M�Su+��=�avK�^ü�1�\�>\�r�;����u�t�?Gq���?��������u�?<щ��E'��u��"�q���h�} FiW�R[�d��V���7`��B�OR�_%;R�D��ظѳoB(:vԣYh���`��Zeaͩau�f����3`ɹ�a�pμ�� +�v8�Z]�J���'\ufF@�w�����V̉��e�9�C]�5c������+���a�Y0�K�M��}������x�k䗑�SQJ&���\��ŋ�����[�y[�n&}H9��d�1�-˔dWާY�^{AN�f��4�Wc�ܣ�}|�矯��HzJ��e�Ȕb�L�f⺬к]�'�~�VD-�!T�L^��T�o}�c��`�Mj�l��0��&�w�>�S�O<�����b��l,��ݳv�{��:��~8�j�H�Ԡm�A��H*]��FW���t��i_�v��ރ򋔙r�&�E(���h]EՎ���}aU��.�3�A�[Nn.D�5�DÞ������0��c�Ϋ|���&�r��m�#�U�˹F.�3P/���v����U�>G����J��ڛ�}��PGX�"���&���ov��o\���/ܦ��1eC�PI=�V��B�<u��T S�ʫ9[�T]�����h{�{)��Az�e(]>q����K=�5���d�p������0��=o:`x�֥���[��!1�"yk43ňu�����,�Mkv&)��L��	ӧf=�PA���xl�!wZ��b�N� ����Q�j��t`��ZY�ʚT��������KiG�AYpK����QC�6�;]we���ގ�N,��vs�D�֥�0�&�@za���q�����`�.>��l��⩫��/u�����{\[k�f�|�Io�;��\X
��V�rK������֫�G���νw;%���7:&����L۽�]�YhU�����2��W>���&�Nj9F��/ӞC�aȕ�#o^Ԩ}�7d4n�y�;U�|Gp�"����'��S��}}��e���#�]gS�]��Nз��
9���s�{��N�J��, �t��Y^�5>��������!����d�u�����ϳ���=5^����CA�KJO�ߺ�&��N�5�m�=u�qV��}��Odt�����b\�\�t��w�������/�]u�b%/9|{dȧ_��ًSا��O��.�c���S~O/�5P}&Ɓ�
�K��� h�c�"�/�*�t'����5C�z�Ș�]P�9�<��{��[5kC`q����DcV�S ^�~V���U���
:��5����.D8�j�Q�=�-�]ӳ/#΢���]y�w[

X��p�<5�IU,����8p�"V�ܪ���<}5���D����~����Ixd�G�e�+1�w� �~��A{��W��}w�S�eh6r4���� m�M���\��}8�>9�#��{�"Y����8VwX*�NG:u���UN��Q����}t�"�*�@?��kK��2�.vDr�<�.���f'LN���!��4����3.E����ם,�VK��s}�Β����/�-+۳�[�v1�7�k�\�"���&o�y�Ğԑ��C��ԩK!�@�mNm=�W�3*3yS������P!_���g�4���b(l�r�ˬ�����یɞ}a+�ٸ��J�Ր��*����㴼�utm�H�5|{#j9�F(�h��qxY
aW�������o�j�,�������g���յ]���.v�M?^��^��ʐA��k�/����H������~P�.�v�Y�)���ӊ��1��>nA�hGf*�Ew'�T`���{G-
�f�\�ȇ���]�3��Ȩ�5~�P�r�WQ$����Ѽ*���S>��ѻQ���$F��>�Dt�\{_z6ƣǮ�c~Sy���;P��ӷٷN��%�p�N3y��㕒��~�����=�j�y�#�zc	��;��7�0�Ԅ!�J�
pp�_b�υk����8|s鏙�j�R��{z�b�*�7X�Q�33&vʾ�ze.��0�)=�C�/2�p��k��P(����8҉<k�Ԇ/{w�f�y��r�x�ȋ@ƃ  �\?0�ݙ��kc��6>�m}R��~j�E��P" ����^��"�c�u֘Z��͢��o,;f��S�0X�F1����V���sԩ0b�z�c�v�{l "��V�$��i�����}b�x��׽k.t{��L=Xur�6�D�q�N�[X�B�r�y�x^Jk�I�8dQ2_��s㺚K�#�63�c��q���=ΒQ�-�����샬Y���$��1 V��`S;��	���%Iڊ�D�Q�)J���j��3�t@���ެ�=9)�B��!���t��~�j��;ݧJ�<~C�5Cwl�c�'��F�5�r3��	]�R+������$�����Ӥk�9�"}��>��{����79�K�W�����3��D��r����Ap�ձ��/�u�X�yD��x��[)ы����Ÿ�d�3�T=�^��]]��a�#��Sڌ�Ґz׌ot�"}e��^����w-�ŵ���zژi#ϧȾ����h^H��>�"�ϋǮ@��#�ܭֻ���eEA
�NKp���O.W1��tS���{�_����q¤�R5��1~��u�.��p9A�r�fj��������c3�;*`��&�|=)�c��@���Dj��m���+U\=����>2�]��	1훻���ZV���^d��s.�xFv�sӆ��+�'�V�)k��)<]V)�D��q�z�10��,�p�	�b�z*����;L��Zu<DR����h��Q� b�{��-�t�m�¤:�J�#B�1�����7s-r��W�˸����dz[Wݛ���v�C�J�w��w2i�K��.X�4�ڷ�����Hnv�C$���X�|���-�OAf��c5R�����n)oc��}p_�]������n�ܮ���mK_�|�����}]9��Uk��1��ͪ٩��U�p��s��'��vH�9���M#,I������s�����$��E�	i�V�o!����c%���X�s���F�'_+u{�'��:����,x����G��{VUR7נ�ڶ<O��PD��=���Nu|������Dž��"���u���5�y��y�C0El�1n2fv}�w;v}�]��T���e]����a�EEnG���*��Z��ֻK�Wm|�Y�C�)t�s�y½�,�ۺ�;��Oʉ��3[z�m�W{�{�NѸ#&�~t6�*9C�>��W�ZV+��T�A��qX=���;U5�ʥ��m�f��gլ�Ք!%���A7����n6zɠD\R��:�;w�;��RB���b�O{��I�m}s��&�"2=��1,�1��|������[�+u;�z*� ���-�溾;�ݜ�;^qU{k�j�U)���g�8!o=��~��V�����0��@�980�X"�����K��e�i��
�sYW�p��\�JY[�z�Y�K'7=�
B)S�>�g�v��.���XI��a�<gg`�V �\�Ю�X�<u}��䃥�����1��tQ�9�9�RWx�-�=cd�P�C[��0샐G+�Mu3NU��	�U�yyM�_]|�ċů���ou�?�w�dP\�ˤ�3�0�
'��әy�u�VmG�Γ46֓�ٸo:�zw��m�{7ׯ���[�T �Vnw�K�N�U�y�!P݊ǘ�n7Q�mO.˕�某�K&���>]�䤮<��C@���ٕ_Q�E6&�l���Ux���V3ж�}�W8"�;ݙ��o��E>^���Eà�<UNK�n����2��oS۸����d�	�Ç�z���u�ݛ	nxÃ./��<�/������ι4��>2�N8�C����Ȫ�y�
}�OU������Ar������P�]z�۹w9��Խ��J2Q�|�T�Ъ��"�v�:��'F\R�d�P�N����	�>��C�"z�����W]T0^`<>�u�,ߢ�X�R&���sw>zJ�`�k��V�Ly�'Ŀ	�wr�~�jfF��d�}=�x|��)�9S��5���8�x��h�'���Z.+���/��]7j�����2r�}c�h�`�>�8�w3䂬�p�$�)	�߫��zqi����
������\ス޻]7ﾯ���E!,,���xRˎ��䵶�։X���{Ў/rf����o�A�[�Z��a��ȅa����okQ�V)mǽׯ+ �J�ֱI�jU��5)���Oua�v;�*�\6���]<:b�6��f2��5��\���A,Z�ޥ�]��Ff�8�)]�(�)�I��d�m�`p���T���
�vE��Y�O��f����*^p�Ů ���I������1`�T�}����7S6-�r4�S�q�� ^oepp�E��_��'W/`�$�m>�)�nuua�/:>�&�\2���w�9�{I��f�W;�ҟ���.�^�a,�+�l��9_GW,�m����ton�B��<�\�FF1���f 9v��x͹i^,��t�zHϹˎ�V�9�Zӊ^�+7��yؙ垎���ʷ��:��hp*� 6����.�iwq/�W=�I�J�#2*L��jeT��(�Лj��b���Y��:>�M�i��RH��|��u�&Y�z�W,����2-E�8��W�A�p~�,J���6��,}��{��Ԯg)����è����Le�ɄJ��p�\���wwf��fء˪��B���G��B�VX۾�A�-����ۮ���3���~����`��AN�*G&��wFi]��]�!a��[�ee���u;��n,L���R>���I;�KW7t�I��:1Tm�4z�%ӏY]�w�=��5u]���/y�V.We�gv��9Y��!n�҇�@C^*0�ZP�Nq�J�tM�.�2�r��=3�9�y��5T�].gM��m����w9�}|���� ��|�Sn�R����]u���J9����^����*򱋬�Z���݌*!68���6^�E��{�w9�W�k��n=-»/E�����FRz[��{Ha���Z �K��Mk��o/_��$�eN�S��r"��v�B�g>��h+o'ut$2��%h�ӳ_I�͢�M\J�:�����@B��
ާbR:+w��Ҫ��Pf�Gz���C2�6 ֡8�⦥�r߶M���Vӥ�.�@99���g���0�s�ۜQ}���hT�Y���5Z(���O�u��I�)nv̲�a\2�"�:��V��+,S{՝�K��̣����9:���0r&�1��&�����WV���::m����������M���i�]]�R�� �Yu������u���Ӧ�9,}�H�8Ӑi�w�-�����&ri��47i>�����*�in���3C 1T<��x�c�1C��;qhGw�s\�߱��G��F靾�Q�N����\z�Q��o'n��ג�E#��H��J۫=�ug1�{)ΰ$V���Q�I�*L��]�ڛKs��}Y=�x2�t���������X(��?��'�m�CZ�Q�B�����TYλM]Y2����v����c !��>*ؒ';���T�����޿����7\�Qڌ���5���
���/�)U�ʟ<��q��"n����q��u�A�U�|_fn�9r���T¸��L\J����iY�o.�^��֭�/]�o���{�򊋅�DҞ^�s
l@������vs�,{1����kiO^㉞�[}����屷藗v�#��<>��u�qqu�唩@,"�q�Z���;���ט����;�Os��L�"8DTt�TMv�����2<E{���Z4�,v�/-E��U��jxyD����)L�{*��ۉhU�iA�>�1�]��j:r�=�ϕ,�����R�*�Dh�ix�CB/�N��Xq�ox�MX�2�KcS�b`�T��1���e�ה6'L��tD%2�֬U��c��P<���Xő��|zKl�`s�����Eb����u�������م�U��ʦ'v�78�}}�#1p�L>m�K���K��.��� 0���,fӚ�R��q�+�'-�i�6\��ö�����KJ�f�<����8'��H93F����d=���+���Kxi`���
��㬍��^;�����k���rm�;۷ ������$D�P��ɜ6v&�j�p�@��S*_�����a�][���{�v�Cy��1�����Y�z�ꞃ9\*���&�EM���l�a<&/�-{c<J����t�3-�v���p\��}�.(�dJ:R��r������{��U{+��gǒ�i�P��WV�<gD����aqT����	�>�F�W]m��y7�l�^Do۳�h����>-na�[���W�*vc��1sj��;<e��3���Z�o}�'עp�Z]�1LL.����m#��������g��$��u�/��W���g�dq�9����=���=<eX�Y���]C�Ci��4}�l{K�oמY������oӌ
o�!�zsz�J�g;Kq�X=X��6���Wֻ�⡒=��gcy�#�0�+��0�s���#��1z<'��YV��!��Ò���^[����Ex��-�,�g*�{�lE����y�A�	��t���MN�γg����*��#~*z�Wz(~���8��ui�@s�Oٴ������:�wHEkx!k����y5P��b$(���⽷InJX�z��-���d.0�� /-=U\M�Bf���J$m�9�`0�J:��^`ξ�K�y�:���+�֘ܭ�&Em>Jmh�����h����s��f+&��87$�"�r�[��C'�^��.<��o�+���:д�x���	ɣs?��덆`�l�"a�?�c}�b�|��6W� vY'yU�v�N�3��D�?Bw���FsL�w���펾����m����(���)W��5���=����ł#�X�3늘|U�d1o\5�mM�<��k��a�=u�;�e�t{���o�ln� �\��z�`+M8i}�*6��A^-/,�����n`���}���~�;2��@�NAq�'�^�Vyfj��=��Y� @1c%��8�$TIOnUB5e�'�ǌι��q�>y1I=$���c��)�����/z��:�5�`?di�zĻ#l�/�����gϮ2T���J|��Q��v�f
�w=Ն�0)��Y��!G���!�֎vH��vʢ�6�I:�(��u!��όT$�l���&+����[zB��T�)���6�Md뙿UE.aX�5!}�ݩ��ch�L�7�x�:��
e�f�~
7`7�QH��+M������ܚ+U>�c����2��� ����c����,�
��5<7i%�����Sv��1@i�x�pD:�58����D[��� ��R���Yc��|m|��T�-����o���&@�ggo� U�����;E��˪4�[1�B���D}u˺�u�M=�����	2ƈ��H���lNA�l����>��n,����$�F��z:�Š�vf��0�Z�������K*�Z���{�k��.o�oi�EF�vյ�����74D�G����K������g���������y��`�|^����<!�<m}Νȣ_����)؟�V>�4yT�ط|�I�ێ�z\��9�5\'{ĩ���7��a"b����ں~���#EԉwfA�ҙyO"�m��m�Y��Mlˏw[�Ϯ���ӑ�M�H3�.�e���9.���hF9=���,���E�����^{�*����W���G�{�%��*�����&^\�k��1��ͳ��6�FT��}�@#�Z`����9��0��U��&{^���S_Nɾ��2��:��!d��#�
1#o9�<�q#ˑ~ܻ�э�濯�}Wy�q09m>lTF�LW^���)ʬ��m��Zq�~,H��3����=9
V��%�gf;���0��ytS	p���hC 8B�Nm�(���9]m�,Q�9�6lP qϦ�����!)KC�F�}:񜅵���.��7{,��R�Io-0�F�'۴�I���7���,H�ѳ�7};�8w�����3�,�y4�F�-�6Ї�[هy�w_%���u������Q�$̹}���dZ�{�g �MB}k����˻���/�sn{l�3���
�Ǝ׌�\�#˼b&s��k����c�=��4s��X�l)M鉃)�h��5|��~��_ޖ�C�N�?a�Wa���p�v�K�[��1��N��2�]�r�����\^�.l�����:u�hZ��º���X��J�����,;3�E;�x	���7�ק�{$�=j���9!�b-n��f����
U���
Ŗ��iF{'ҍ,�D�R}���oר�<���v!]����+��sgݘ�\Z��U�wz���rYG����n�f�CO�����>u�X=���2��J��V���V�2���C�����Ğ�]w�&�\No�2e�6H���6</ʪh*g�t�\�����_bkQ⾊�[���}������=�{z:�.�~��x����G�E����Ju��s{j�e�������6d\�F�dE���"y�T"}u�jW3DaN�Q�I���5���Y��ې��,��%VG���E��߯jjx���
����&	�o{z_<���|\�֨�+g^�la�\<G���ǔ�v�|/x�\�>�k�=�0�����U����9�wb����'�iJ5���#�aæzEu"��f�Y��q�E/���*,�G�0�E�W�^c��,S�rv_R;�N�ɱ��ܧ�C�r~�75��&7��]��ĥqc�z�fuJͱ��	E��[0�H����H�K�]��z5i�����tY�M���!�u^�5����_0�$�ǪQ�P�]Dz��b�^�5"}����@B�l�u�/�S�Ԅ>N7��d�~���H��Д����}V���7�����C-�6�������!�V�x p�4w�Fw�SC���f�����o����, ~>1��T��V��M�F��*�xr���G]=�b��d�#^�߼�B�����N�예��0U�׫iq9�G�����������h>��%���s���
@�=�-��V*2�rգ�!�� ����f:�g�ΧbbL���V���V9��t�0�(�t�~�T���{���00֔���x�imo_Ձ*zcY�.�a9ǯ-W
�Wu`E��Ȓʔ���:���D)v��n��q2Ne
�,u�n��|0�[�Ar�]C�f8��c�^��o�-NV޾����ٺ�/A��}�{yQ�%���+����kn�v��3���w�&�%N�M��U���8�Q�����(%)k*ƭ������o�G�>��Y0�����-"K�_���H����D�(�=����Ut��w�H@x���{拏�᭴�3�"3k�3����x¼v����� ���y;�:Ѭ�9��:B�嵷��������Eg�C��q�r՝�J�������/H�Q�w�SY�ϴ�|Wn��2}��ݞ�ׅ2������u��"�~�R��ë-]r�z�k���<'�{�vA��:`�dd�������>k�<�
0���,4,�)5ׁ.�H]�v.b�n�q�[|��x���n�nLdu�@|#5M_��z�z��r[���;��:�� ����t]�`s�K�!���{>�#Lo�Dp��A��teץ�1qY����ErVf��~Y@��ny��W@�9��k��՝e��,�^��NlC��,1�~�'G��_�$F�a+�=�udi���w�����=���vW~���8�!&�eI�d���ҥKʽfV�mT ]��Ë�*Hyr�뺕ݜ��q�j���r��K��ݱ���[wn��Wh�[E-��2�[�o'U�Һΐ��WM���2�KP4��{]��ݍ}�e(xS <o���P�q��N�[دz���ϻ۞�=���~�Y�t�i��z*'�3��ڽ.������S=���|Qۇr��4w_ǼJ�\���W i�{Vx#�C�x�M��jFVz���3\*�ڣ��b���� ֗j�[�|�xA��z8Q쿰�9r#��썇:��4�������]�rڒ�*�˞[_�u���#�3���L�`U��c��C�G׭_ e�뜷j�O#_7�Z���y��s�Ա�������Ւ�?�5��?�������zڐ��ġ^p{<゠%�ˣF<�B|^���9m���3�wr�w�9���Q����5��5K��\��7M}��a����JځSӻ����"�E�;����*	=?Eۏ ��;=����>�iq�Rf���Zi���E��NT��2qq�;��P��TI�} �U�"�����yy�؄�LN�O���8��tҩ��6ϱ�����qn8�={���w�gـ�-U�s��:�1�z �v�֑���5ĬdԵ<�p��C`��}r�W�7Fy4!�K-�]�d�h��-��g���.������0�V�,�$�:�+���Z��;��ս7s/���;����_<�0:z*(��:��IǮ���#u��7'p��S��rXv�#w�]Y�/��ܾ"!.rY�K���[S�t��ܛ� �6����|3���Q�cjX�ݺ��@���'�/a�:�E��Ą4}4a<��	ƻ������kj�꘹��@��ר[��Ɍ?x���;7v͡�v���^���W���W����� �=�)ȉ>��6��#&�y��H�_@f����A�Q����ڌIz��k:h^�;��O*���r�ޘ�CMρ|����زL@*9\���r�ʭ���[�^��ܱ���F�̯��F�(��-��R�\=�L&2�.�b�E�F���37,;v�� ǽr�@�ܲn�if_	���qȸ��P�OԏW��g+��F�eT8�>��1��p�ø��^��S�����O2caH>��ݫ T�^hM.(��2[��^[zl�;�F��v���C����T�0[;H��g(u�՞ㄔ�
b�{k+��Ӈ:�h��^g~��e>��ɼ��{g,��!�%Q��qN/'��S�J��;�v���PǺN�����I�Fu��#r�d<�����++V�Mד�T��S.+rsn��V�@����˫	��fpκ�<ӡ{J��n��C	]P�&D�����v̚"U�U�%-kg3wz��±�ӡ	/Z9��*�dCt��<7�[ �7W�[�} Z�k���7�n\UL,X0�\�g73m�Λ?�M2�x��f�-������u!]�ڧ�����јJ�V9�Y��l[��伤d�<��/\�yK��̡Do�a\�%{�D��|�dV1���h���SS�s���=;Vx��s�h��)���F�]'�ãˠ���2}ҏ���R��T�7��ɻ���_����ުD�ws?:Q���ވ���^�W�s9�37�D\'�!xG��ʜm]�t�o�����sP���"bF�3�U�c�w��^����U|��s�޵�}�yȳ��+�z��1ǆ�mk����80�Y��cv�+4����Q�(E��mykn�](�s�RbȮ��֪	�e\5s�nR��&Mz:6�B[�@��lC�(4�׆�˶7u���ի�h�����*���F�s�4c�o���*��ǣ��%�
��z����:�B���j��X�mE���W'�6�Tk��=7����ҍ�߮�����Ta��[�NϢ�%5�)�D��.V�O.�]����]Əv�:�fOB���ͪ��RG
BՄ�kZ��3��4���fKI��g�I����o1Aku�!3za}{�X�9Rr�Bis��Y�eoܕ��t��Vc�����5�[bV���|Q�4�e��|�wUɇ�LUu�.��u�t�+58^�ՠ�5�M�5]pVy꫱A����K�զ7��X�5`���4euBy"C(:�7�9|ް��odB��b��5Nhu)�{��j�{KrpYC�A٦���e4 /]U�y�%ճ�d'g�[�s)���,/�VU#{G�3u�-�����Gu��鬕3�Gk�]Ҁt�Yٯ��:{�u[@��Q/�ش�ؚ��jt���Mh����2�eW�V�cZJ����𲡋����AӒ�iN��Y��^�{1��p�|Ò�Bh�4���ڰ�sQ���Z"�rF���(p.hI�Nqh���C�iq��XOJ�[|�W��8V�.���M����mr�4]�u�r��0��EK\�g:�t����\��*;�l-� ,U��4��}�N�p�C�ur�'���L]Pg*;��E+�8��<g���dy�V[�eQ�,�5���yt���C!ʆ�:�i=N�:�5;Ds#��{�/d�(��ҞP��j�'����|�l�2e�ue�F�u�V�*�n�ڰ�1X��c��oej�ʥF���uJ�v,�IU�d�ȪS���'��00�$RVb��;/�rw�169Y�U��h�u���7��Zt:o�F��q'�x�B�N�n��{K�����>��T���,T��h]�}����v�=�5��I�>������XB��]H��&I<�-|��}ӻ��6����Jyv`ܓ�k;(���D7h^�&nH�^F+�sM��esV�rKmN*姤���]�а�R4�R�j���uE�o�K�R�wJڗl�zph����K����!�}N���S��v�͌$(
]/�[��:i���\��)�rT :� �T�w{�b���!ot�E��V��f���5׹��*�u���u��D��7�1���L8��[��-���EԌ�v����;�`�bR��Cӗ��R���/���R�����Q6���ig�جu�.��9��"�<�����mP]�1�hm����8{\Y;ZFvz�~R��VVV]��<̥#,#���� �s��5u���!�m��XY-Ko��{�N���r��4����Wrݹ|���c�@\7z�ǴPi�pt)�]]�kjR,���[���[���M�l����w�����-$�e�2����s�.�V�Wu��
ۣjt�ڃ����88Xk����6�s�m�+$=ܯ3����3�%�[��v�5V8�����k]�\���0]�0����6��6h�&n�x��OOW�W��m�2e#�K�-$.�ԣs����e��f� ���
�Ftb��ldb����������S�5�H�����C�3�f�`��=b'�nP<7�ߪ��g��ν�� b|76�r����G����<M�5��w;l[t�A��t���Ȟ�u�Gkm�N�v����e:\��r�^�G��E�b�ҷឳ���>����M)F��7�O.��M��8���4��?�ۑ� t�z���-���j#�ˆh���s���B=��S�3��S�%���3���E��n$��ۛ;�7*2�FE'����W=���{���Q���a렾~arpcVID�2�bq��ﻎzY_.�ũ]��?~�Yם��E���J`TyM�[~�%B�~��/f�x���p(�̝�A;2{�/�ӗz���'���Ƅ?E�?��)��<�0��o�����@��Yeo�E�F�Qv�.S!_�Qu}K�2�{�]�=2{�=�HyS��ɥ�7�G�t�g+�6�^����¢��Y�0�ݕ�}���$O�V��ъ_��T�I��k���vz�xk�j��
��d�eq�ޑ���L����S�VN:~HK<厥G
���}q,�N{�|��`Ky��О����I�%U.3z�f�Ѿ��ہՎ��I�������O�ŷ,
�����h��>�m�{���Z�.����V���Q�Ձ�j�u�n��'v;lv����@��'��(�ɪ
��9��d�\o�\$��^��ڼ��X�'�t�#x+�� gh?��� %�ɾ��V�VS���S��:=����MZ�f�2zX�p3�j�2�wj�Qc;��ȕ�jp��c�p8�h[Zӵ�)նq�.:�w��ҏ~��a|�/3����}��%1ި�F�e��j=��V��P���9?98gS[<�)hʚ��:������ݕ�{������~Y�x���ܛZo�υ,#��l��w'wR~����>K�խ'k��H20�b�n�Q����*�7��H����'�7�_ލۊ�[h���r3�=23�J���"�
2��S��*��c���*�g�8&���+��N�Nm{���?,^6}l��[�'aq�hk�B�j������F]�MvT��󧿾�8�9��s��pr��>�����e����
^�`n[L�k�gz����f޻�_�Qޙ�@FȎ�ƨ�Ҧ2�iP�yC��{����m^���P߫����x[��Z+�ܺiD�b�B�OO�|-N������4,_��ro��V_}���a�����	���I.
�ֆI񯟿vU~�U�~g�!�(�c��D���{��#�W��h5���%�p�G���l�a�=���|�Gs�ڬ��58�k�{a�=j�b3XY����u�0������7���S���.�ȉ�&z����禣��m�р��J���bw��cS��rI������0�HF�.v�N����$���ګ�dft��
�b��g }:�������P�u�R�v鍉�k��+��gP[����FGv�X������;�S�AVuKāp�����`����~B�r�T�Vۘ�xz~[(� c���[�%HNڎ}��9�40��qǯ�k� G����TѰ�N�/��g�WsW�T	����ʋ�s�+��
Y���"�e;7\��F[�G<�Pg\b-�����/L
��3��=�u]����[�oM���O�.�����
YUWx*��������C�9�j��W�+���h5w�/a�kGX^�V&'W��9W@q?	d��vc�W��.�����J���ʗ���C\�,�ջ�����Ƚ��ε�W#U��T]�T5�|V��k?���M5���F�T{�������S����t�.�G��OC0��������b��3�B"�K�,�e�;��A��R���|������CrgCF������3�2�L��M�L��lDӎ���T1�C�a���Q�����1��ş/�ʇ�Ԫ>	��F�ҁ0v�TZ|��:���(�z�:���G�G��;JXz�����mW�|��Ɠ�����χa��ж���tn���!j�3��'�#RV�Աi�@������_i�.+����O���U��J��J�11�z��+Z�p{����r�N;���b�f��(&s�kE�zb|�wX�ͮ��폩l��.~��+��2k�v�����U%�yՁX��pٜͼzjrt����j;�-��׸��rJ�9A��<��!K���fՇ��;�<����h�b���	d���q0#�å�K�\�{K=��r��|��K��y
R��q�q0���^{���ܿx�xܾ*�u��zp�gݽ*�Ő�ŻY�G�~��w�w� (ļ����G���$�����W͇*���0W~��P:X�����u����A�)/�wTL�����-��ޅx���a֛�i���b`�:���B}1S�u�0G�:_��i�;q�&!��͘���
?����҈W>�}m�^~��9@�f�J�ۯ{`�o}�<~�C�p ��R�|�i�t&�#'��]QQ�~���e�ҹV����_�ų��>�I7ɖ�Z/�Tiq>�S=��=P,�@��!\�����l��_�P��N8��
�F��g�LDz*"k��l���_��S��fl�U�a��7��]�k�T�7��z<��3շ��:a��WfɈ��-of���r,�q�3�8x( �����ڟ���T�>I�T�[6�?]OU��4�����1ƨ]_"K5WU;PtDd-�|�;��d�l�a|2��+E����r����P��d)��F��__5W�U:�)��~OҨD�����~d��@�#-��YyV�=��.�\��pj����S9�lQBPI����b���6�oΟ
�{�
����pu� �V���c���8�2d��5+ӆ6Ή_����z�c��ڴqh��o���C6�'����ir��|����]�՛r`��c�!�8K�����ۈ����?f��۸����K�ꔪ������G�7�� ��s���E|FP#���s�`������s�S��{�ˈ��r��z`�>�ǳ.��d����ĵ��ʢ�f���>u�'o���:��$��ݼ9~��UE�d�3y��%�"��I���M$�]�=�( ϵ���Q���q�s;�e8�ܮ;�;U��W*�za���ʡ�����P��:�Oٰ�����ք,1��!ǺbȲ��a�q�W%B�O	��!x����ϥs?��?��o��۱�vm�~��
n��6�������`��4-�3�~�g���r�O~�T��Z~?d��of(.7�Φ�THʆWϦ��"��6w��ݗ�������2cGTk~�%n଼9����lW��g����. #!������qϜ+u��ݟT��G�#��%���#��8o�qK��_T�X�����M���T�}E_��gbp�G�S	|>�wY�ޗ���b��[�o����1�����[L`�<���GV �Z�a�k�\��'��C�>�h�+��9=P�4p�#�j���U�T�R�{,��05}��f�`�v�=P_۵�a��}�p������"�>r��.���*b7�� sGG�p?z	I�̓f�)��'Y݇Y�:�9E`Y[�']�=���K�G4���EJő��"����0�{[V�A��p��\Z��|e�O{����)W>�ّƕ��"i�̛��eu�n�*�o*z2MK�7�/�`�PQ�W~ź���"���1�=N�{_�۞�Ï�NmN7�P��LOa�W�9}v���}Y���b��Y��'�>�oJ׮8ʥuR���z�����"t}gG�^����w�n������߳[؏"/rN}[��s��N�aqL��Ɗ�s/���b���" ����H��*��kF|��]
���+vn��#��P1��E�����V����<窲���"��t�����+�=_e��/�����z��f/�(P��?X�P+�w��QYz��o�Dv��D�(����7d���~sw\?z�o�e6.�O]�)H����u��uԭ���Q��}�Ʈ��N�B���,�@��I��{U�Y$t��^̯Bƕdz�����~���叼K4�#�4}�N��>��R���u�{f���H�jqCDp�~7 �_c���IWU��H�?W}��M|%�¨�E�&���B^�`�)��1��v��!������
=���XU��n�-�Ϋ-?Vň�87��+>���ϴ^ø�ֻ�����s��3$��In�|�h��Շ��!�5�XW�@{DҾ=�-4=��&�����[��ZiW(��s�1�?�Q�1��b�Z�I*��糣w}� g`|U��˛Ԙ���Y��~S�D�]�Q�AD@Ha�Qs'�_E�����Ec�C�g�����NaAZ��b;[�PNj���=�U����O�>��B��ق���U��.�W��T�wc�+�N�~K7GAS�w��c��i���y�Q�-�aj�/����Wp��{�fb�Oi���9�[A��S�&�����]{�-m/�|����8m��ů�L�/;���W�>}w&3��9^��xw��{���^��6�}�p��y��ӱ�؈�pş;��Ӑ�	����W��B,D���U}�#���$��`���g1_�"`���f*����s%�ޓ��6x:k�"}�������B3�_|s��N��O-��p�̇=��oA9��ɐ�u��=�&v���������5��$\�\2ki�C�xJ���|V�����M^O�폈�Q���q�1"=?G[�?x�)�2%CLLb(DH�<as��>�|�
��,_wO_���|�}vP��V�ۀ�:�������K�r�:��&�D��*�]��{�vL�
���,"���`�1^�A?_dxi���Ϙ��t������Cs���\���{|����ʨ���O*���2�Q�䣓�j����n�}a���S�_V�Q��p�>f���٨}4��y顃긂���#��ѷN��mN�Q!�iE�G�DV/�LA�����@�� ����/��P=���0��nw�0�>���2�R� 	F��$|�C�M8����frT4>�r�z�+;��uG�dT����pr���u�W+����	;�!ꦾw뺯K����c7�
��Ӑ����bf{��}����A�a��e��l����;|""k�ԣ,gVH���vG\+v-&�>�,�Ab�O�dg�ȅ:�/�3�b棜u�	��+���w�f�lŋ4�?W�G�J"�;���7���i���w�h92M
����R��.�ę��H�(��2R��DС�3�wI�٥�q���}u��� Fn�.�
7�>we��6�;��hە�n�ˇ(�]��Q����40})�&�A-��eq,	�䩳+�H[�Ҷ���n��C��H�ڒ���p�dԙw�ָQy�2��Y���a�J�ya���[��YOL7��x}�D��q��nDgj���s�a@���7��z��םTs�����:|����7;�g�����i����1�4}��\E�h�������|�3W��u֫��r��.��Ķf;�i;{����a�TX�|������}��������a85�0ك��fh�;a�k!��>�9~���bȐ:#Zl:V��_�}%+e�}y�9�d�ۙ��$o��M�VNR�nc�`1�fYsy�yO�잝�Q󘌙�����46ZH�U�f!gW��w;����U]�y��cq7i�';K~����_ZH�ÿ�1x�:����/�;Q�!�$�}���S�����)Ͼ�㩸t}��I�2A�,�y9;��NCp�#��Os��b3f�Gpν-����>͋CAf���>��á�����h��y^���b�\P�g��悧 `��5cF`bz�n��;.=����^J�O����A'ܹ�3���/��ΐ��sA1c/���W��������8z��\�9��7S�*�>ֲ������:�s��531�P��K���LE!���p#��N��?0����C�����_�~���؈���g�h�_ч��jK #�|�������G���R��nۃQ=��c��6[���|kE8`���d�ߦ�#��H���)ȗ��9����{��k@�Q��S
r�*c�쎟�R]1���T�>��Ws�A�8j�p~�Tu����\7r��^o��vR�c6�#���v�s�y�^|��-�ԨTU��<�#׹K°ggY�,���Ƒ��S�1�v^��]n��H���������C�b�+�&�w��.�
1Jv���׼u�惍���G����7q���o��q��pQ���]}�X۪��d῰8�M��UX�׳Y�L���Ý��p'����~{CϾ�LoҾ�}>�?p�̭[$
p�׉�����թW:T�C蕚�k^�u��>��n��Uؗ5Fy�}��u�Ԝ��f�r�h�����h��}�Vj��VO�T�6Z����#5��C�.#|����g"^��~�����ǫ��߽a��ē��a��q&���}���b���l���E� ���Q*bDp�:������K��������ha5L�����+L�E��Qf#*��Ev�no	��I��B���g��y1t^^@�����������bvw�̕X9e��a�>����1@ D�&/@��t9ڣ�{��L�yဃ�PXH{�M�q�rB3ܡ����`�K�V�~@�>c��D|�w�y�/s�h���i1F����G+l\��N��@���-kZ^���!4�vk!�5��Q�f&2T�hv}�A��q���!�|b)B�O	��]���%|& �:Z��bGbD�{K^���;��}��3�q��,G�E�b�1b"�j���1 ���ܤ�s)�뻭n5��5���������q�X�C�+��FF��fsCS>��h�MI�?K{��Z}@����sc.D�(pĴ�On����^N�7� ��s*��`�f����3X}s��my�l!��H�k@}j6����;��͆'��%�ui=���/�d���ԫ
�a\�r�������+���b�pPGۧy��d@��k�c��{�[qQ�s��Ɖ��Vaøe7EGq��B�y������2�CF��[�b}I��!�j��7*��D�Qy7��}o��W;̣���֮����V����U��;u�Rױ�=�f_��{��Ŏ�m	wX��f�7����n�dװ~�9`1�^L]���rP]P~/_X�ȥ�x�o,�=�
����ݍʔ����Mo���쏥ҩ�U&V��[G���ȓ.�����5��fm'ŏ�p��lL9�NN�=ݻ������r/d���7R��̥_��7�n\S����|�0�Q3�
�K��k��𹇣�֋���F�����FƉy;츔�n���I9��A�C�MZnstr%�7�dd�]��%3��S՞_sQ��̌E����z�������&#.�~��_�����>�dYwFG33�+t�!	��_���a���@��;��~������M��1��ߨ>�k)G3ϰx�sIg��kt���w_�N�>� X�?X��a�}�v��}��՜�W������*8�p�	��{�7 ���٘���S�����o1<E3�k��r�ӜR����:�!�� �#۵�1�����>���|�j���o\蝏`�S�;.9��$.-cf�3u��TD�c���N�sPA�'kp�)XjG��>��w�OD.vcT����ɦ�w����E��U�?c�}�d�3�Ư�ɬk9ٞoz�@7 ��Ư]ݩ�#��Zݡ=Og`l��L�f�@�	zպ��Y�����J�AP�І`f+P��P��@MD�\��!�>�{guó\���z��៬���x��\���{h��}��n�Y��^@�uX �CY��9�}T�z!��wt.�'��� ���}���#����<�>����U��^��I/3~�����������n:��QYVZ��]A+�� ���=	��F���r#�P/j�5.�`����Ӹ� ��.�DE���3���^������yC� k4�����@�c�$ϻ�=��	�pnn �P*��t� �q3n	��N��S1s�E�A�!Py�C*�b}9�{~]�9�9������pw���(j$�`b)��.H�
T����8�p}&.�[�otMb�[���f��&��Zu����JE����5�ύF����)1u�.f�)���6j}i�S0��������_܀�*��?e�?���PT��P�Q�3FES�@�r�e
 !J�PE@D�� Ty��pPA�*���P[�  �_�ue��b���aU@��������s�O����&�����{��ݒ�|� $$��u��QW��RB 
*���G_���P��P���#���In��=&"�Bga�9��3;��rw<�P��/=��)�dBP���)Bp��형�Ĳ����n�P�zvΪ������l���1b��em��1�{R)a�y�1R�Jy3w*i*��F�jBq& Y�Z��
�ڃ6-�*��o0C�ښk\���)��HP�Bj�dX��;����B��+������ֳ�FBY�q�bx��`I]�@��ܫ�p��J�-�`��1 �ӉF�17�z�ԀJc�w�Ob�1�-Z�(,�Eh��<��-[w����*  �T� AU@ "EU@ �U̂ 	JT+ @�AAb�A(A����'��g��		$��(����`���HV͙���BI'�uHF{�<��h���p	����5�(EW?�`}���������
*�� ���ئ����I���
*�W��ʕ2T*��e��fJ7e��A $$�uVT0ҀITdk�TB0.���8$�� $$�u����@e� HI$�n���J��]�.��}���SwL��Ƈ�q�l��?��=�m QU��'�z["���"v���ŉKVgA�;�2���Zl�z:�z�PVI��~lӀ�w� ��� $ ������.�h�MM���PF�%��kQmM}�Ԧ�*��j��T �I[v���QD�b�ڙ���)��v�j%[d�UYY�Ԫ�kE�p� ʫ��RP�-�&m
QRmJʩK@髉��듫���d���!�\WKQ�]n͚i��Rv�u��VڇNۣvӭ+�������)M�ާ�:l��7]�w���ۥ[T��KI�ԩJ=�R�W]:%Riu��l��١������vQv�ݹU(�+D����λJ���QĈJ�	IR
�     ��    ;��[ xS�;��ÍPS����vK
=����m���9��-v��{{hU���V�E���Fl�{���ǳ�rw;�;�-����RR^���԰��@��C��ݪ��B�ͩl���.���#MU��q�OGlw��=��3����=c��+�u��G57��g�z��@ʛ�]U���{n����	U%(
�U@��ݞ��Www���{m�zB��[�s���Ѩ6ݱ�ӝӠ�s���n�M��:����[`��v�9ӭ5ٹ�t��4�����Tj��F�٢���hu�]3V�lMkbtz�Sw
��l;���ih��:Q7��{��h��;��c^T�oK��Vm��pf7`���V�Fק{@�N��=잣4
{�u\󠊂"J
JE�\�{]��Ws8r(5A۽Aw�C�gp���]
�ۇ[{.�u\��Եm�����<+�� ��7��]���aMth#XwnJ�16R�{j!��/�.�hLu�u�a^�@������wm�c�yC���2��4�����t��{�y�)(��ri+v�!����=�wC�d�7rU���;g��U��2��[�f���I���@u��w�zQS{��j;��1cZް�4a��@��9���,(�����m{��=�Q��"�eJ�^؍Á��.e�k0ًk��m��t��7k0=qIᷣ&���=&X�JkF�Ӻ�=��TB�{۞�X'n�^���mv�6ݚv�5;�\�����{!\�Vk��8n�E[lf8PB����RJ�R��N�l`�:t.����`���m�U�g���ú������;��ɶ�'��Sֽ+#g�T�;�Т���ҚŻpRw��/l��Z�m7n���]�Ѿ 
�� j�R � S��$���� 5R	<��'�OS@4�'�S�IJ�   ��
"��� 4  ���%(��4@��}��߹������\cH�=�F��u���o��a=#Kx����Z÷���X�_�*-3�t�B�Av���*LW�R�yJT�QP6¥@�l���u���~�����b$�s,�GX��ksJ4E�&K� ������md��n恍�˺/U�@����;��Y��9���w?Ró{5����X����^�vs"�y�v��p�Tz�=��Ϙ4�@�E�f�C8�iv]��d
�5���[\d��Ԡ��,��o����v���N������J&Q�|1s6O��LgoL��7m[0e�Z��X9�۔�Hu6B�A��j�J���Wu�Ύ���b����8l��"Jgb�_3 Q��x[�iS�RJZJ rٮk4EL\J�#Yj�IZTC,u�9���t�k�(��Pፚ[�S:���@ak�*��V��r�7�����
�7s�X�V��5W�/�X�K)�$�,s�����6��"��-b�u��3zSP�e�b:�8ӭWRf%
�+�ǲ�� ��9U�P�9Ne6B�����c��+��^��-��@���e�Y[��M��021Oݸ:�y���h�#�(�%?�DItƋ6�����p��Wg�ڄ���r7֌Og�u��jY8#�0�2֍��x<{�,�7F��N����o�v�.ۦ�n�w׭�2���Ƅ-�۩DIR�q���;8,�`siPh�lơb�����
����n���Q��N��Y��[t��b�XtR.��CN��fм�ڬ�A�e�
���b��j���_��cӏFk�)WuiѮQ6ء;Dg�T�L(�+mu��@m��7�EiYsE
��n+�,eYH����pu8��e]��ūN�y"���d�a�ԚY@���Rޣ�[	Y���M���{T��`ţ����BT.�1
E�'�LԧP�o1�"�z]����͊F��o%�3q�ZS��\T��.<?aɇ�N�/Z�C�p�"��X)#fĚ�,�EbJ��wb�.�"�oE4Q�P�[�%uJn|�h�@(����u�y_�]2�ɡ�ݜu[���C�f�.��/jK6@�9�2���]�JSz�7�1p��r�n�U�DGut���|�	�p�d֪Q�eq�*�B����wZw2.�0�������#�i��s��1r��!����dr�V��Y�������v�o%g1���
��@�� ��kA�+��ossO����,R%cG2��n��
1�]E��]��kt�b2�'��<���O�PHBuv���Q�}i���He_�ץDK��I�|�.s��Gk&� [�BZ����k�7S+*d9.	E�T=��n�jdCF����7x5����ujooe8�V��V�r�e�Å��:31���-x0q�s�����^Xk�Q^gӭn��+,��36�WO�[в��ٽhC,����~Y߮Uz�A�m�Z���t0�{KdX��n�(�ѹ�'��n��y�����~��ͳXeeYP�}6����o�.�����b���kd�m�pQ�J�o�	�2�X�F���)\&b
������l��do>�p��ʎj݂��2n�u],%:�̑yN`�V��� �bB���i
�6���
2�z+�xH���F�]jEk��sqZ�6r]�u�t��|���r��N#0y��e�Hr��/z���Zf]dT�<�=�e�B��R�����7*�еŚ��2��`�X�m59��T����H���u�#C|�1pκ��;l[�'���^W
�d�0���t�6[vAo.��C��"�q+��f��.�����£ç�.K;/�����=������
ʽ���n�S�]�K�����yk�^%x�4a01\�\��M�|M&��js��Z��T�eaB�w�S�]V:]d˛̛BVN��i�����E�^��eH�A���k8K_=�^���52�g]��6LTvӺl�C,Qk�%9�C@'�r�8�<����y��4oz�ܶZ���Z�C� Y�S9H ��L�,��t�Ӡ�3�����M�4��%h��׊'F�
���f���lb8-�r�Q�n�Jb�	��-�H��e�"/Q�s����-u����\��Tux8��Bh��L��vOS[q�5Q�8�ii�;0�&�3�>�a���g�ح��F���K0R�c��x�в��j�ײՆ���a��7���<���bS%���b�YȆ�˂��Q=��nLv�+b[���Aωq��Pj����=.�ՙS�Ah�yYn�j^){��N��?йeG�չ��C/3^`C%ɦ��`�U4��/�L�uTn,Q�b^ɕ�Ѧ4��m���q��m4��&IQ�X�U�t�+?�`���,{	���Q��1�tM�1E),9�Q�Q���}D�..wW����p�-�äL�mQD��]�P�{	n�c*�sF̢fJ5+�M���t�z0N���[�#���G�+3Q���Z������g��h�Qa�6�u��=!w�r^��e�٥��l L6)8�ۃ*=p�e(sy�o�����=��q����GݏV��������J�@�@4���D4�[��ӷ�p�fұ�r��e�݌�ڍ��l�Ummt	fmkxVY�6ab�PedZOn^#��$��Q��URN��T���ԭ�e�8-��C]�ڹ+2mZ�*��^e����m�f�&
����iC\�c��5{YJ���d�*	.�b���Nm(��S8�I���4�& �8Eu��(�G5s���N mnٕ;*�@/�7����u���(�i�u���]'!��JCMz���bچݪ
b��en�ŉ�3x�N�;
�N.m�(sBe���ǝ�៦�, pf7λl�� ���X E���i֦�v�͚�u\e�³Q�B�а���Ǣ)g<4%z��GQYo�g.�뼊�7�B�^�K9��.4�2��#u����g4��.��VEZB���G�.�E�,� J�!oD�!��W�;9M�Ћҥ�{l�r��	�)���SU�CH�w�z�9G�Z\-jYyIQ��y�;N��̡Z��������˻9�+��\��9��,0�D��2���u��ʡ{��忺���MÊ�6Pʛ�$��`y(m���]�ze��օ@:J�u�𾢎�msk���n9]׃(�8�m�2�$���Ԧs6id^s�-T+���M��t�*f����D,ٻ���Zxi�~L6ﶝ�Ky���۷�k�V��O�Q[��5��oW:�o�Z�.�:�*K��2����9&r��S&4w���p�Zn~]�w7�i��l�P��M�a�����e����2Z� ���N���	�pdO[��K���c��w&Q	&�yn�
���N���9嚱�?.��4��v-�.��ONg�\%���� �톆�Z�.��R�œ�-����^�(EYK9�ޕ(>�w��Ȱ�MWx8��U=��ϫ!�X��ˢ5�.��pv��Z`�ce!�E��N� Ԯ��Z�q�����՝s1
��n������Y�:
fXb�����{$�v��L��f��6T~N�����~�ܻ�.~	�og�&�.���I��b�X�t#]+_uu2��7e2đGl'�mV{��4^����qݱ��r�cT2�"hWJR���ݑL7����0����L~{�/-Vm�O6H�W�b�z���U����s2���������wرet�Quu,;��=�g$� ��|+�$�n�qR����j��[rbq�\%G]�]쭋oY�d5����t�2�
�"Ҝ�j�B�ۑn�6(�6��A�)�B��㋟w��V�|F&��"����C�Hﱦ����ф��<_cv�7��LU��ۂ�p�u.3��8'WO.QY��@��M"�e������5�HT�v^���F.#��9:z���v��CD@w1�s$�M#FM��Dt��5�N�/��;�����j�b�y7�ذ��.2�:3"{u|�cV%J��eech�Os�t4���.5�$(h��:�[ܙ��}�eV�c����=�SǝR��Nԡ+���܂+t�]���<Zf:;����f���]���õ�(�[���#�$,�s:ء��SV���Ѥ@b+�,�n;��{ۢ���J3�U�-��b��n����ۋ�Yľǖ�mڭ�zoU���.�' 2��I��b �6˧���yF��gkCJfA�i��=rf~���9GrS��T�o1ɻF���']͈z�K���%�h�Z�92�ۂKL�t�ػy=��:]k�-�{r�-���Xn��"\��T�,$��-T�"�T�ɦ�p���]!�i��ԐTZN�DE	C�Lɶ��kK`�VS�M[k9��ݘ���X5~X䆆E�0�T�����A�Y��ٛkj*J�=+�n6m~�u��(��"(���[ZRȰm����V<�.�/�iu|H�(p��)�	�u|�hnEO�+�%��}�gc}��j���+	��*��W�s-A@1�&C�F�f����q�7w2\�WnX�Spjw�B�ʃJ�t������kH=�#C8͂.�f\�b��ѫ:��Ta��Y6��#��r`ۍ�74a��
��[�v��z^,�$1�T×� ���V���d����ZJX�,Z5��u'-�q�؂GD�ZvßR���#0{V�7�����JQtZś�gT#�����/�3bU�`��:��0�ij�"����%���ݦ���f�q+k]��f��NS�n4��dduE!��Ui��6.H��M�MlIM����:��.�i3��P9t�rr�n���ֺh=���Zu=ѧG��j�J@����0�,�a��b���y2J֔(�L�n�^�*Y�����u`p��z8� �bT���kb���<���,�<7� �XB�F~ۼ��x��F�S��d�A�!ܳǔY�ˑL��:�ǹj���+E�n�K4�pi07��I��z5�ih]R�5���N�	:9�آ�Ӽ�٧K�9,�T�ؼ6qI���ⵞ�Z��e�-�X��È�}uؠ gT�;֓֕�+��M^`#�Ol�Afw%)n����M���-��p�1�U�A[��l��N�p���h�8���t�!<��W{�<���ŘEV�P�gS��*[r�=���8�ݸ�y�l@�=�j�kz��X�i8DR$1Ѯ*#����j���xݛ�8��쥴%�n���q�W��t�nXL=�Yo/�2��WKN�B�LHIh���P�J]ŭh��PNtib�j�!(Өгj�ܽ�1�Gp�ڡ���q�$�]��:�
�M$�
�5VMƌy�p�N�MH��[�%����a[ר�Y����	9��`�����j��'Q�}��,bЋ��Wӯ�X�ۦ{#�q4�^�����kj��R���=j�"@�YH+aD�Q|��,Ǫ1��\ʛ�M��iC� �෹���e-@,�R@�+	�l�ŝ5m)��cE�r�^)[JJ�wS#ӎ3Csdd0�	d"�d���ul9�g6��
�w�v�p�m;Uk�hQ�+�*:���4[2��%Fi�E���D��A.�5�#2�)V��i+���wZ�X
��Sba��E��x��f�R)2�u��t���'2,j��U�Lf����`��p0k.c���j�NT㼛ݾ���m��_Z�[�Y�%��V�RJ�X�l>�]:��OJŸ�.|�^�쮽�-:Lz�M1�@��RP�`yQ)��+rem�2uʎ�)nbXs2��jZЂΗZP̷Q�ب���̢�i]vv��_+E6Ԍ�Z�'��]�c4n�,Lݭօ���AŅ!z�v�[h$pCN�R�����u��ma�KEZP>5�ZÔi&k[n��|�Qԣŗhf��h��q(�fP�<w���.�?BD��s�1-W�]��;�bKr�p����h�婭/�k�U�
ʾ�>JLh�1���^�wRhJ���7�
0�Jm>�����q
��K.�.�S 0Ul<*�M�3v��10.�r�zJ����%���:s%���H�r��dNvw��VYn��P�M*���d�gN�e4&D����C5�/P�1+���a�V�׻%ʛ�J�a�U�Wә�އjI+؈vrZ,$p4�����2�3<q^�eZ��	��ei�hѰ�л۱t r�P�U�9[�*?�� �&n^�-ê��줮���F%�^YC�r���"Q@�*�d�c)f��G3��x���nu k�n�����4��z�\v(�g[�I=pՓ��U��<ĖLŏ��܂Q�][˹ŋgb�Պޣt/v	r=�S�ˁ50_���M<�&	�l!����S*\дl�p���8�1��K�r�{4�"cXgF������ܲ(��K���vԧ�?F�^��n;B��,X����i~|*�\[�o"�3K��'M*ư�Y[}������7/L��J��s���%;�˔�6� �I& �;�*W@��Ϝ밎��Xwb�
K�ī�}c{i�L��Jyl�}���j��)�EC��n���gnA�I�n"�0��j�.j	<�������lB��LP����L�8u]����I~[���Ӓ�=F� ˃�q��7zEX�O
b7�-&�!��
�7t�<A��n>��6�9��ܤs�<�fS�w8 g%��_~йӰ8�$��^�%��+F��&��kMl��I[�D���A��{ ����aY\�R9��m7���s��kyz)7uoH�NJr����[F��w�v�D$з�a�i�FV+�m�U6Ž�c#��	+��Z7z�C$�VX�j2�/�%����u�(L�4AS\�U�3mb8(o(.!�X�h��i�j)��iR�bE�
��[���:��sowwwM�Xx���$o��m�zZ��|u7ՄnȻ� �/&���k�;��n��sm��#}$o�������d��\m.m�$������0�K�����XY����J�m���ݕ/Y/�I�#}$������s@�����]�bsZ��I�#}$o����>�F�H��#=$o����7�$��F�II#}$o������G�H�I�#}$o��>�F�H�I�#}$�����7Ҥo����7�F�����f{ww;���7R�H��0cq(�	)$��#rWId��(�rW$��i�@s�K)l�O-�K\�H����d��m�e��I���n� �W%��`B���aZ ��JX�$�B��S�D�T�]alR��Sm$�7@��$��#�R[$�[B��]�� @�Hn�h66�TC%�Q$s�����)]BuT�Fa1��6�H�p�l��&���^�"O7m��v���q�+hU�	˪�j�Dݕ�hc�@�*�0�[��@X!�D�+��c�|�$4TO�ٰ*v�TqCQ4Bߵ��{Fh7��o��Y7׎ƈd�^g(&QMk@F�=���䂤�uO���D���ӱW��ǔOM,s����sSW��~q�.ǝD�C�"�,Gq�t�,�;vnP8�<�~K��1���>�xn�ՄG	5�K����cn���Qg�C����5
��9Z�Zr����s&��Z?E��pT���`=�̗xH�j���'����ous�܀"��W�y�l��\"��r��=1Uօ��d�+V5t'If�WV�m�����hW�m	�>sJ6%t��is�jCJ��7��V��pvZ�� �M�dfi?&�{ZV�8�Q��Re�u�kM��d�/�\�Ѱ�f;�%
'5�+9Gn�ʌ[��L�@iŬ��? �e:���[�`i]qK��^�j
�GZ�rBnLΫ:�1K1ժ���{w���uA~*s��dKB�^�c�ط�N@w;S��R�ø�tS�e;=Z�]da�pI��=���v�2�X�V�� ���,!a�*�>�hS�e'\yW\���J�S��͕r���ރ�|��kB�X�д�t]^T�V�F�Y��vT'L���N)+wh���&K��t�m"z�mud;s��IrR�����`�b��]DN��]�k�k�n��U�qӵ�z��^�@��}�1��ō>F�xÊ�H�۹�snܰc"[�W*,p��wxs V�,�bBZK�n�n���e�x���	=W�Ǜ����sa7��K���sU�y�QV�kSr�ަ�q�4�w�#�e��%wO3��H�ܴ�d�!��fV�]���[�S�_����g�cDmn�
�ת�p�ZW�l�[aK�m���Kɯ�g�\u,�:�:&M`s/}z�q���[XQ�ձޢ;��(������%q-cn�3N�7F�wP��0Z�j]�
jm�畨Y�L��Ɉ5�뢭8�ܝ`��;'`8��zY�k�vc�4�3?f83�
��Ί4���x���n1��d�w(ޞ�y�k��̮���F�9��bŦ�q��]���B����ʌ�3�y*��V[�p9����O놣E�ݘ"�.�+�wY�*7x�Exe�ʺ��bAJ<�L��孻���r;��B��+Z9Pf3\�F镒�1t!e5B�QY�,� �"rT���?��_E�k��ҭ�)N:�d/���ӂ:��ҷDJ	��e��]e�n�n�u�"6b=D걧��v�=���1- �ڨn��0��wk3iʨzL|�>H��nZ�t{Lfi��D��x��`��7]����/�ë���&lIM`oj��J�Noھ��ufo^,ˋ��]�`����k�Ovl�/�SF�e�J�R>�}75R�f7�'Kh�"ɴy�c�M#8%�~ǫU]��֮�	fbt�e3cP�V]��ڣ@�n]C]S �*�%�Eu�}L��3Jb��-
��0h�U�̀�ɹ����R�)Ձe��FL�4<���+X�Nw1�ˇz3ih���}r��F�]#��h0g:�n��{��WlMSg��w�����kzm��vEG[�j�6Y��-��đ�Cd�f^�ej8D�K=�����ܰ.�'�MM�ԯC�	ǉ*�pP�,��\ˇ�v��ђ�ֺ���,�?(����Wg)B�b~��C5`U'�lU��S6�\`\3��ޝՙ׷õ�v�m9@�2����l'a�S8���b u�@3E]���\���'7/��wO��dfo.�*���]�`�Djz^�������XEvŠ���e,�c���gcFA�?K	��W
��,�H6�.!�y��Pn]�wĊ)�+&K֋W9s�w��Y�v�ĝg[.�N�|q�1�j�)Y�%p^���f6�䥽84J����Q�S��;F��l�[:�����,!2�������'���t?޸�긇�U�y'��&�2��m��U�� d�Ŭ/5�Z�Ał�0�M-��I��?�C����5��z�x� �]e0�� ;���nl�a�L�u�2�N;%��1L��nMf
���v�yͭ�VΑ�8~�.�n$`{4]�趲+��nJו4/�Z=�Ԧw���ޒ���Ql���2�m6�n�'Dƻ�c�Z�ð��w���R���B�$�Y�.�Bg���mj°Ff��}���!��i�m��(WL�nN���\VJBm� C�S��L��ܣg��	�2�����w;a-y�T��?�8;�=��N� �!=����ِ����em-Y� �g�+ȩ���)w�:n��n��:f�|��.jo���ev��	�&�G� �%���wz�-[Ȃ09Y�4�v�\�\����QY ^�x�j�7r��YJ��=�0S5�ގ۝��a�7"x��K'p쭬5�>A����£��H�[8�o�ǜCl���'�tE:�O2�����a��˯���oJ�w]�� +I@U�H7 ��మ�Af���6	���i�;�ΆseDD)���(ٻ)����ŔHP�4+�Lc
�v�!����g�։�uY�M�h���oJ��z,�9]`˕��S�c�li�U�(+��/Kk�w,�9��b�+�i�q�ZQ�H"���6mZ̵��,�m_w��sٹ��v>�px8��!KFd�*Hٺ̏��)˗���,��/��klQ�M
�b�oq�-6մgF�F���mg^\���]��Aaco����*N����FC}E��m�ZwQ��40�ѝ*��&:g�8a�aȜ�X�l��l@�#+3Hb�~�vfNEPv�͹�����Ÿ�2 1�p��9����k]e�n�tci�(�Ь!ո[���s0�dv+�=�e���&�0�	�E�r"�кU�`��m�묵�lԝAT H��l�S�u�Z��ʝA�%��/�ˇ1�2�A!0��'H��Z�|��� �D>����J�M%;��k����#W�]��N�D	Z���y\$��%h���]�YW�׾�En�(`D��Tv�ͷ�4e۽�Me��x����6��[T�t,
M�-l[.-M==]�N�Ew���U-�(���r�|+c�	i��v?}9�O.&����v�+O��
�/�$؀7�3,m$\�;�{�gb(&�K�.��G���DT�&�V%�h�)�58��eib����N��k��Y�3%��%w%�`��
T�k��u&V��)�bdYϥX���T{Vj:��S۪~�J�W�� H�Ϭ�z�=t���w��ܠ������	��3mV]$U3��եL���5�^���G��w�^��cA��}P����Qɶ��Z��[vN�^KTf���[�,�8�W�FY��G`��H'	7y!m�1V��z�7b0)�GU������5�Yݒ�Z�5�{y�d�"΍R�f
��Y�(�i�U�`��RQ����]�tܺz�6��0\1l�!��Q"j�̼.������G�V`W�;f�����מ!^X�+rӧd��nE���3� �DE��5��x\�\�]\m7(�O�izbyU�p��g}�[j�{��KM�Y;�����	�6�<Z��|h)�j�j��=�K�$	��k�߱A|ʉ�]TA[T���#g-b �ե	<��\;ki��D=`�
�
9f��FBHv��U
�u9��ݒ�AB*n�hr�B��="��>�^z�LQ�[��|�
�����3 ���h�d9]���@�9(�W�S*n�t���h�����g�MFы�hl�-�iV�]d.��Jv占2�.�'ɛ���
&��8��o�^��&�m�he1e����b�xHd��QX�V�&��cƮ���w7��(g���{w���=�M�|����Z��ɤ��l۹�eHS˪�Y5g�� q.Z���H2�u`4��p���0$�m\꺏J�Mdt��"����Z~�2��T
8��ҥR���us2�Z�zM���)�"ioq.�Ǌ0Z)��[}F֪�4I5ّ-9���t��l���h�̫��B�%�O�K�LT����aԦ+���u�0Je�{�]B�=���ˉޗ/Q�q���u�|8{O;��mK��>�I�͸h��hV�+�Xd�x*��G�8�\6[Czw�V��1h��`���kwa;nh9��]Q�<v�V쳃1�̤�J�b;rFH��7or��B�*r�5�$�9)����a3�;#6��ޘ��Ej&�Ώe`J��CO��X1IQҍ�N������k�P4�/�,U����*v�Lr�u�ڢ�/�л�:������ꀓn�%R�P�RҪ.��� �C��0��%iΑ9Ubӱ��`� �*�F��*H�4C}n���ޕu����۠�oK���Y�&��(�v���6��	��D����db�K�Z�$PKh��xJH�"�Wa�20�I�r�-�
$��E#g+������Z먫0�ۤ��<�Iv�j� V
�@qF-KwJ;�b��[Smb��]��GZ��vK�-T��̝��J��K.Ӫ�M�+꧵��a^dR%�uT�"��Nx*��זC)^S��ʊ���+�,�x\{�qӻF�[(���n�(����e�����E��xH� �ف��F	�M���H��K���T?��L�#E�O���~'$���îT0�a�f��n��@U��MK�r�� A���QSf�l4���IM�)����|�e�4�%����D�]�%S?���^\슻��b.f��H�G�1��y�]�Y���p�J1*�tFb�%L�r.ư@Scz.?/��^��1��Sc鸪|�G����Sʴ��`R�� Ğ��F3+���niw`��:�VK���6�Rzכ4�#�[�Y���tRQ�Ο�J�Ф�{j��Y��ͷ��@=e/x8�=\�ج;o$�e+ˤU	Fَ��.Q��sx� �)!�R�C'��ੳ�eN�L�u���+/��l�3��ZnlӘ�f��Ŭ��d�9��V��`�Oi�F'Q,�2Wb�2�t�GOduѤ���+��8��:9Z.�[9F���A�\�b��6��n
V�3�;��Df!}�aDX&��J�,�DHN���i7�ㆉ�&�=�6��q?eg3m�����{�������e�qՠ��W)@��lc��\�Y�y�S����FD:O醍��,P�]*��9e���9+��-��<��/�КB6�>{���Ŗ�m,޵f͵�n^�t`�ghP��aB�5�&����l�E��9Γ�z����[���D5[7YwWݛǙ��U�|�tob���P.�OK�w8��i\TPr�Kr����ۡU�X#�9i\]&���7/�t$����q��"r�tr�m��إF��R�r�G��䷶������t��@��c�p�"P�]���F�	�T:��__Ԏ�Lc��Ii�`��Z(T2�oP]�Ӥ�+h둹�^P��sNp����\�
�C��*tgP�I[b�Tr���,��:��E�a���)�I<y9F�	p�H���%M�XAY3�R˩�	��4�F�d�S��[\���޾w����Tpg�)RpY�վ�+-��gO�ں�u\'f$Pf�⡱��;���{��Oy_ڠ;I��F�|V0��\%����$)#�nd����l �N"�q������6�4� �*Eu�\�f< G�F��|<©H���.�
eʀq�9Y�e1�y��b�+��hVຏ��Y���m�� �V���:JRR� 5WGt�MSeY��zv�x�����R����;˶���o��˝�N�de؁�hT�[�TՄ@hj�V4H-���P��tUEnS��Kѱ�#��� ��Hs�N囷��C�ܩޜ��we��-�ଷ��ȿe�<���Q�Tw՘h�f"m�G%�y�͂F̢)��7R��Զ�n�4�.��k�{�5��R&td��z<�C��61]�=ơ���£N4 æ�m�lE������w[X�igo�����*8'q�fГ`U��=E�H�;�;�.E����1�_��nY�%�ꭓ����q?�jK��[A\���`��U�>�f����f\Ȑ�ǽ�c�ZZ�;��8:+��rZ�[���Ἓt�G�Y��T�e��U��TiQJY�oq��W;`������!��̭��Ԓ���z�P�o�����lۛ�T����$��������8܍�oe�U4s�Rʻj^�Uv�@E()��f�T��hhe05�F�p���_�3�0�ۏ�nfdI�3n�e�7DŴ�+�č7Q���� �3l��.f�E&�}�ku����'z7+��88 �q�%@�L�E�	;�T�L�igE*ˎ6߮�8���6�<��s�N�u��C���\|�}#�o�lOu�*:��pBLrD��܆J;[�[d����]�d�[[V��wE�n5f�H����3I�R�B��2�����*�+r}�,Oj�e�[��tci� ��beR��G a*�H����5���IGA��{a�)6����聳v����9�]wN�I�.ʤ��o
��b��A9�p���
����{O�t;���ڝ{�rQ/��itAb�($�8W`�6,�Sn��m]�E�N8J�M���:�d(7Q�\֖.�^�[I�  ��.(�n�{���[�+1j��&IOx�*%�K���p �!�c"���8�����D�5y$1m'[]�����!��@��Ex�$#����W6V2��x�6�f��*�R+a��R�;tM�����)��~I"�m�x���h	j�j�
��� ��S��8;9��t�Q���պ͔WHx��;Q���.zs&�F���K�_8��l���e�8R�Hc"n�en�P.������Z���j���-D���s2�8���������f�s�K�~����������PG� �4�ܷ��ܑL!o�z��V�#�,E��(��Y�9�EZi�(�*u�XV-�QԻ:!KT�:p��$���d2KD���+U�ըw<�J�i���ܵ��w2���E8Eb�N��}cqq�t����UE*�k��Lq�T����V�j�;����U���sK�AqL��S���kӆ��Gj��$U:��8'�m:�D݊�Fe�`M���}O�!0kӚ����k����Vn�ΆqWm�8s����c�T{<��A��a���iq󙗓��]7Y�on�*m�깼���i���뛍q��� �:��p�Y¶����ai����2'�^E�^��e;޸�3\�Y���AkvC��鸐�ph۷ZŬ�]�GK���i��ێ��s��8'�V1R�n�����ϟ>\��<f�Jpn'
���+eg�A/��z��
�d����[�6�d�.��q׆�Д�y�ծ��K�F����x�y�I�CǞ�k\��ms6MVM�0�w�g��J'	GW\�LMG�1;$�ȘԀ�u��e�k`]w٭��B5e� ��#G;2t�6�;l��
�v�x� �L�|s{c���%��c���s����e]�Íf䭳���o&�����H^Y�_�� �BM��
-��^]�֏>�ӷ������{�ww�|w8�?�=��|
�~^T��K�o���k9�Y��˃�3�]����ul>����;����*@ge�Lx���#�ap�c'��X�=����>뫦�-os���^f:~�5�XA�<;k��מ�0{��+¯�J�Xkq㴻! E�΋��}�I�֞����]��1�eP��@�₹�ve̙���Q�-e�E�{�nn��'r�}��Y�#x}Yշ~����	� �"*�=ԡ�yc��Y���^�KBjy{e�s�%+'�||?��U�5�Z�q�\�gSY��S��Gi݄W��ʵ�;��9H�GcWFZ�MP'�N y$�A%D� D��6�<w�O�皡�"z�(���`�pvD�xQY�o��*ӥxeC^����;���P�Z��[g�/��Ғ'���u��73Dw��T/=��[�$̐W�?=ݓ;2_?��^e5y�� ]��]C?H�E��^;p.t�t�L�E�hksu�;-J�C�X���v�u��_W&"�'D�V���X���<��nNCd9{�U��X�Ы�4�vI:�V�	zR}�Jc�܈\D�� �w��f#�ٔ����Aq㉭�~���A����R'��)��Vh�eysg��2u���yJ����{���~�kՓ��s�&^;�62��WZÙ�ZJ���HK�1����yyb�q�nNՙ^��J��w.�<��cw�J�h�����I���y���n��)�	*WyM��v>Q/7c�T��^���fmp׉pבwvfÑ����|���^ĭ�eə��|�pj��g������c�v�l~]V�>lOW}���5��a����H�'LCċE��;b:h�a�f���\��i���ڙ��c=�}��w��2_[����5�-�^�T�={�݋�5mx���I�5�Vw>uʈ��X�XLf۰p��U�lz�t�Bn�]��o��#:�:��fZ�Խ�
�ut,t|��r�i�F�a�!!~܁��E�y��7����ah�[�n��H��(���P�:�Q�1pW���
�n�{��W!ʲ�w���R�ͨȽ��������kdV
}S3�#M��Er��T��{��As#�k'`\�o�Y,����;��@��q����=Z�J �/����K���y�`�m�wi���#jW���y�t�vb�F��ƶϸ���.:�I�zr�m�p����w�i�X1L�==��:<�C�� C�]V�f�g"����[�*z����cnk�����H(�{�{��w�Y�'�2�g{���B����7�1����Z�@}�f�_��t˫���G�x$}w3ǉhP�8�ů=�{���0?��^-�'-sF�
uh5��f�B�Q+��}eF��ip�<s�#��&�O@ǰ>�Tx�(o*��cwv q`�j��%��qd��5���?2Y��q�\%߶
k���$�C�;x@�B�>
��]L�ߌX�d��<��l��L��z�׷wNf"3��'��7�����g��!'�$��А�3!�x�q��e�)�)�\Fy�r�������o���|qꬉ_XDź��(x`�N-���@h+���G�Ӿ�%�иzb����`L��yR4����銘.wD9��5�������s$���@�"��Ct�a�hk|ǈ��n^+L��wp](����5y�<�w=u2]�I{[��۹����k]
�ٚO�jߟ�<�-�N��`R'C쾎��]��u�����۝�����`�ݏ6��բ�
7I᮫�&<��3��R�jnՏ�:�G�������FBwU{�U���=�tG�}eoHߨj':Nc�~�u=AQ�Ϋ|�+h���E$�9��FuB���f饤\3��q�*�rW,�<"���T4�ą�Z>^���T�ޓu�!DQ��u{=�<�X+�Y����m�9K w�����ڗ�������E�¼y1fW�H�K�J�O<�i��-�۩�+>�j,��׾��1t\�ai���R=��<l�{��k��͢����1rxPw��q^��W�Sk��
��͔����l��1���vt��*��@���+�.+2��y�`��E<���k=�\u�{�A^�����$��H��j�A;�F������g�Y�E��j.��|�q�Qɾ��žG���m��P`�3�|]����1�[����F��VZ�^ac�?wv��:͝��j���(��/M\h��l�E��C�kC��ǯwr$���r�����Yz�"C�>�����3���7t�Dk�R��=C����D�����\XbR~�gi ����p�\
��CY���
�M��e讄�OM��f��j�+������b����BGK+l� "�2z��oǗ,*�+��'�vP+�(k�#��]G�G�xsM���	z���7�F]tL��g����o,䶭��,Pj?�b�j9a(�_��DDO��h�����K(���_m��[j5��}�U��X kYʾ�%��H�b7ƠȐ��dlO��e�����p�.a��J�PT�nk��|X�4�6ψMj��3��Q��c���?�@ouRB�5V3f��͝�Mο-�((��o����}�c��#m8��ӛ����o�OӖk����X�Ì�[��Wo��]⇝l�맲��ר7x��D�����)�wr����%";��`�N�9�Z<5�OC�����ފ�o��Q�Ho�Yٹ����Ï���8�]e!������ ?S�� -���:�p&�b�W�~D~\�\�*���o�>~��DKڷ�W��G�K8�jU�y�G]u<Nױ@�/j��fj��彽�t��d�W�Ǉ��>��:�(ћ���z=T�T�����כ��M���r�$���t�~�������ծ�r{�R�=KG���~��|�*�,DB��'��P����EI���]�w>	��/�3���B R�ȫe�(8��ׂ��+��l{��zj �;sˏ��������ڼ���ǯ��K����� �[���J���.��h]M3G�����*���yL_B&��SLY�=��,/ˤ��+^^Gsjr�w*�荚瑝�׸���K=eLE���D�R�+3�-�]����E�qz[�{;�q���,Ǡ��������r�T9Q���c���������<�EQUds`s:`�o�9
W�ޓ�2�>��s1ו������=K���럮�.���r�g�z8)ݕX�6�h�G�|�d��!�B����/�{�k�A׌�Ql�c�obv�M��Т,�)\�{'��Ad�5h�k�up��m�{��ٝ����ж����������U�~Uc�rQF�E���T���QoD~��go�X4j\�J��K[��mF�)Av��`����q����?N�c���$+���=.Ou�3�6,Z`��#��>�z?V������:E����X�*�=Ȕz^c䠍;08�kMu��>|S̏>�[y�BA��Ǹ9����-�s]q�=��3,a>��*x1��o��7Gn��W��ၘ6?$��=oT~)3�&h5�6����P������r�i�$z�ѿ,��2��{��8�=����kH�U�]>�=��]�����c]�I5�����}�K�j�h ��i�E��'��	�u��xcS���K<���'DZs��))O<��� �̹�v�sCC����`-�A�]�}��>����2Qٵ����L��vB$5�$�ۤ�@qSYr�����`^�^���޹���v_f���i��b��f��[���XǏo��}YB�L+}�[���0��Ɂ3\
(��W���~���8w��6�M�������m_�y���+(GٞfϚ�7���c��kgYb!�N��h>������{I.��"��]k�ጺ���r�>+qei�ƍ�%<����F�'�s�cF�K6ߑ#��!e=���ҋ�Z��\2OҲ�(�?�l[/�5 0ܪ����e��$f�L�1r@��wi�$g�F��)l��k�cD!٫�Yvx>q�E�_��b��������#�Z�/B9�d�{����n$ډ�z�Qc����#�F���f�`�ryW�����+n�=��'�'e��x�y��4o�xJ8W�lxz�7�X�Ԕzf̫��FحvSFٞj`�n�2��k��'nJ�+�W]x�T���.���׫i���A�8�-��C]�~�oh<��;�Ux���W��eO�E
].������Ƌx�򗥑�#����x�F����R�Vj�4��[k��V;�y�+�c�v������|����������҄.�Qv	�ۦ���evn��|v�з�o#���P�GnZ�vd��k�e���w���][�0#�]7, yE{W�oWrv��%I��d���@]�=ۢ��|M�\��m=J������T��򱣅 $1x��>]��O�Ο{�y���&�x/�U���Y����R�d�z�^�N-�'���� S�*|j�����@a���w#m�5������~��Q����;N�L�1\{�B�V��^s�E�н��W�Uwsjx�q�B����h�
�P8�4I:a�غ�X�(2�0WxR�#���`=���҉��S�j��*���p~�Y��N]�h�s���{��#yz�=w�̣�ubѿB��/V�8�Ò�;�
���*�qY���a���\dg�^��ٜ�Ѹ{��胣����WV��f"w���W8D0M0O{�x�k��f�엙�|[�{���5�n�s�B��W=�WC��c�g�/�<}ŭvc�����J��]z�C��#����������FW{:��⨎�G�\���6��{��H�'ۈV^d��U�h�����u�[~��~삄�mt���kxM�o�Bo*>(Wi�Ą�2��)!��1�j=J��/��D1-f�^�[�N����uJ{/2�\��m���4fwL�[���[��wp�]M�]��k�m7c�X�z�l�IcQڝ�U��>�X���ɲP'������U �}Ɂ*Kn�<,B�9Ce�F�
�f�R�����e� �i����h�e�[ڕM�q3k����E���'b#@'+������&�K�\��~�t�Tg�ƃ@�F�3��H\3\T��?o�F��T�簰\u�[��H�N��@�N/x��W���ǌmR0|9mcZ��D��F�L���U��L	�f�%����ObV��T��v�y��v�i�Z���h����l�N�v��m�$�wA�'��پ��y�?�1����_��ڕ��|�r�zfyY��4�����gga֮�%{����2�4}���L��8�a!����s��
��ZQ��K����E��/
xr��w[~�HxAV�w�<ٽ��B�ij��d	���>>�\�l�C��[�-N��r����I�hD1�ix������E�J�6{��dѺ0m�w�G��%�o�*�}W�J�kV�b�@x�Y�JlQ�l��m7�2���,���]�W `p��cnC��f��v
���&��z��0�ګ��^]��̙<CC \�}�7��t�e�2Y٪h
+�SlBȯ��_���"�4�H�9���I��T�9j\��_�)�{��:��sܗ��|�֭��-�Oi~{1�{�������b�9�,����W2f�`UX�D����{�d] σ9k�/H,}�&Y(w6�D��X.%�en�	�eВ��2B�2��Q�gpm��:�K��T�G��p���w|�<�k�iol��y���]9�}v�s�t��6�p��8�g�}�v���H�S�歞�d��W�ұy`D�%]�KvL���>�/-<�oh���376餗:~��+�y�鰳�uh��z!ڏ�fڞ��c��N���к��1�	c+�v��疣8�`{gfw[�X�%���^�\�����A�5��W����x讫�U��m�wوMv�5�{�vu����Y���+�ףؤ��t�BMX�~�~�ߡ���U�y�d.�m�=�>���ьeī�4@N��U�ٛ��z@|W� bAu�p/[�[�o�y�&h�Q[����s�ܞ��	��3B�錫�V)p�s�w3GI-�XBTݶ��T[ކ�./V�y�;av_��F����J9k���Z�
��W�x�y:xi;�*���v�ȭ�Et�4�ڥ�!;�;ⳇb��R&��R�Ӣ��K��{��k�. ]ܼ�47�?{�Ơ�ޯ�d���-�����8^-�ۘr�E�;;7�´*FO~>X�m���'�G��.`���]���h� ���z�����e"9q�'r�v�vŭ�{^ťo?���l(ݽ\5��p�wj޷(�^�B����c8m�h�X�PEQP��[S�>��)E�ޫ��!��[��T�Uuḱ�ٸ���r��T���W�b$r�-���.E��l᪒���#�X�yk�ʝ�Ë�%�"�e:���YLր�jm]Y�Jc�yK1"o���`��~ԤZ�!Ӊ�}jd�ӝ��[yQi���;S]���)��sg]|�9`���ƎL΢�[C4K��Ŕ�OG8�D�,]w��B],ܡY���3�(�<���n���c�3������f2�%�n�`һ�$�/��2ic�ua�[wz�l͛ߺEu3C��tR��ʚ�_Sk�0�-bCwk�	*�죨�G��i�Ypt���U'x���onpT֠��Fk6~��V���h94����R�KOjF7ݏ5
�g0%1��GW%�p�1��k$grU�#�iB3�*�T�,ƨ�pO�e��@��{�q^�)�5�e�r<n:(��TX�*l��ז۾WW%_n�Cǂ�c��z��֘#.��ܹ�e�k�j���Kj��g˚'!\����WAbܒ~���ٿ����_��i:%H������-MJv�ne#Z˸�յe�G���i�ͺ�ư��%n�����Ua6k(�������!���P�j�9n���qT83]�`Ur�[����0_P���Vw{86�8To�f��z���"9�Q,	��/^��nH�F��UH��:�.V���s�٨���܊�_U��\�Q|��G�Ȭ�<�c
�V��j.����+Rk+O�.�h�Ӱ�%vɭ`�aU�y��_�5uh�6�Ջ�7ho �u�3O>U�]��6��dr�gR��׬J� hV��0��� �p�p� t�sX|B�5��cj]F+���MU�����]ƫ������y�*׏T��Pkk��O�6�oq�]�X���0T'Ƭ��cxQ���}a
���4�H�k2w<�����z����­�{.�����k�4*t�:�w��vq�8����GG\�1kL��n�p���8�!�"�gt1W+��$���;b�.�܈S���I�M����/�}:x{�s_��۬�Z7
�k9������U���ɐ���e#�U��ʬ�_�!���,�̋�~��Rg�G444�x��S! YD��<$Y����< �#L�P�y��q5:� j��){�� a�dh�^u�s�Y�O9����W֧~�a^Ë��p���Y���B<G�A����,�Sc�"�\�#����0��i�<��v.r� O��<$_W<&j<�x5���#�8���3�IeX�	ze�gG><��~�,��>C�$Q� �σ�B8	ǜh�8����bn�.Yb�4y�>��9��z^�|r�e�a>� $
 �0��Θ@d� �m @_M�c���K�tY�k�/�TCL0�H9Ӆ�<y��1���޾Q��.qb #�J>!�YF��r?��,�t�"h�Q�<�|x��d@B����qԯ��1B\;c5�w{PGȉn2(��n A�T�4��R���9D29��-�ʤ �G�i��� K<� �����(�F�9h � |yS�Hy�JޮY�?,��A<���	��< ��4 a�ǝ#G˂��0���!�=�bϯ����H �����@� �4���f ,� ����@i�<�P��3� �#rn��US*#��H�><�p��O9~���t���gX�a�!�G���gw*���m�wX��adq��������+ɚ<d�e.Q�"x00��<��G��<�OO'˃彃O %R� 9�,�Y����<���?s�|XE�g�<�EZ��A C�@̥|�j�����k�v=��Gǜ������{��x��#�񇌋><�q�|�!<�(�Q\��*(p��_}8.���$28�\$ҏǙ�C��@�!�CN(�\�<��	�����ϯ��)9������<{��������9ظ(���!b� d"Q����Q� ��	���8ˋ��=|d�x�B7���%�#W��#��Q�S�����^4G�٣ǜ�9���Ge0:D4x�t�H��hB�$Q��>|�-s��Ǔ|�(��� ć<yG�D �'�~��6@I�#�	�"�<� �x�:E0�<��}���y�2̛�fn����)�����uԥ���*�><e ��V�PO�k Bջ�nvAcS���=+���su���J����{�8[b��I��mà�#r�ǏS؜�f�n�?��Z����r�U1!D|@�B� �#��Z>Tx���,�"<��Y���G�x,��2.Q< �s�Rr�sH���!r�0�"0�8��?ydi���� ������>������s�#�x5,#��s垞@-p},Y� �r�#C�@�ԅ�y��� Is��p]��d<y���`����	J��Ň\��G;?��4�\�C��
f$�ØIH�?x��
<x��QG�x!�� �a� K n�!��E��'�.x�"����d�
 yQ2<@�J� <���dryB9Qa��k�;��k���J������� Ev!�x<P�	�������<�8�9��}�O8� i�DsH�����M`g���W��h�C�QR�<F H�=���Ň�!g��������������m]xa��Ds�� $��8�"oX���C1�"��q�q|�.�	@��>#@!�p�@� '�ߐ��Y@��釀|���/��x��|@$��,?)�q�WO�o;��<�:x���|@�^�?P0˷�(�#�GOi�I���8>�h��E<D#�C��_��8yϚ!��F_jv�x	��@Cg���"�sK>#O(�ic3�_�K�e}{�w7����|@��$\��Y���x�(� ��G��r(�	���:t�"B!��}`C�#�{��3DWە��U#E��#��Hg�G�9ͳ�>��7���ݞ��x�񇁐���W�8Eq�\D�sڇH��g��<#����a�G<Q�� �<#�b��!�K<w�,�g��a�\��Ls�\dk���&�����|�¡*k�nn� '��f� o.�#��$��ඇ%]��#J�<��	� id� ��v�,�k�QG������<x���hC��o�Dr#�	���	L�<���{Y���>#�i� d��3���w�q+B���<@��s��j�L ���>2/���C<�H���ψh�x��m�G�`�9�C�<E�C�_	��E@? .�#��2֟��44}V��-��Q|�Ӛ,#�U��|�HM�����7���i$��ӽ[˸�er�ަj{s���w�#[�6៯C���������[B�m���+�8�b4y_�Mt��:�!ucu�l4�{ ��0���s �j k����Gȋד{�GoB *�S�]�F�8�:Pe�.5͆)�����(���U	j���G$��X�~(��Y��WZ5'��fB)/;Le��+$C*��f��l2�NH�,��EWJ�aR� \	�i�H J�Ϝ��|t� /��!�&�����h-V@�>��db=~#��@$WQ#�!C���s�(�#zX�'����O<@G���pB�-�3X�m�}���7;��0��	 ny��0��W��!:l�>o��x ^*C�#���� ��s�"�(�M����rGt� �0�"4���|G�B����(�<yG�@
�<�ˁ�@���_ï����.�ٽ h��S a 9ћ ҏ �x*��H�G�#��S\'�<�ޘ�~#��g��|Y�<x<z@���E�3�#����������AH!��r5��|^�s;{���2S�T
FI ��н�<v�;�p;ɸ�N}]Gϧ�n�Ǎ����y��NBTcrJ�2j�3l���!�ᇆ"&<J�������:.�l�\lQwl�Fg�1��Y>����K^Su���k���ud�z�fK=��c��dEs�%p��`6C�N�dV�QMmf��Ӱ.r���q��O1��p﯃��W����4��xY��	�D���_](��o.�c�nk��dWk�Z��g���Ψ��@tם��=�'��c�d�B�t�v'ۢh�̼���B��GE�Z'��X̟o+�t+�d��
�H5E��DO��EW�S��EJN�e}�v9b]8D�/n[���y���mې�ƙ�)��6Ј{>Z=�Gڢg���9?g>��=쮫��i�7Y���Hb����4=��XP ����73�4��s��`�����b�$J�כY�R�r���xܭ�T��[Kj�tw�0���$�Ŋ�=(�`�8:�mA��P�յ�,�E�ٲ��e�����ԈS*����W�k�țTV���#&5���<2>����\]x8�1���u7�G����{"�����Ѵc���׹�\Xb��bQ$��u���*7�f������W���'���Eқ��s��:"��"Z�ͨ0��Ƙ�����j�PTן�ǿo�W��v.�ّf��_t'I��.�`���������e}w5Y�jTzz6M7�̀@�r�*�{�z����!�ʹ���>1Ys��4�9�_Me %s���N�>��f<���}s�)2���e����y�D=�ק��S��B։�ۭw��kc:y��J�Ż%}M����ZDÅ~�>L�����i6��7S�.'���F'#��PN�Q�v�� ����p{�"1D�ϯ��P_\�ހ�Ɗm��E�������ܹ��Cb]Ĩ���#^��4���J��TMU�ڙ���5�5T���ita�l�S8��'�lL��I'�,��hب0��^����Sl|�����j�܅�6�<�R@�����NP��چF�)�D��]�8�lW:�#�V��=�K�?'��uM�ݞ�.�F�W��H��9��5,�Xq3�i��e�^}�ɬoجfk���p/�̺�����%#5F�9t��r�NW�swe�jA߳�Е���v�ww1�������.��4A@��1�a���Q�]9�U��ʳ��:h']V���%:͌s�0�(��̀�t��������M>����W��٭i �~��r���J(},"`�zbb�Zr�]dx�mu�*���b�8{x<��.ˈ���s��I����m\��`\���ۏ'�͍�Ӏ߬�����Ft0�ZaD��	�9�'w�������a|����=�y�?	U��h<��C��X�����j�j�"���ejq(J��O�;h��=�02ג�LO�D���AV�H���v!��|�v*W�㔐������f�+Ү�"��9��x訝�\�\<��b|I����''���Y��g����WR�lSr}�M�|��Zo��Y����Xn{e�?K��.�*r�~��ϧ)Y�ndl�	�,�삯&k��fLe�^�x��3���˵(9ʴ�Ubkx]϶a��'w��1���;�Ս�w���;��;���9=�xN.��pb��f����0���Y�]X�z�Z~e˯�u��\a>Y�������ɘ�|��9��]e��)�%�ع����ޞˋ�U��PUkS�����}����`D���c��p�#WvڝsVi1U��Z0<��[{�x���J�FS���`r<����w ]��cw#���9y�ؚH�MQhei������VN�â2К:��7�-;�Y��7�w�Η���tVr��<�,�\��y���8q�=��3&Q�A<Ͼ���	s�z����U�%G�0���4�ڙ�/z����9�G\���S���F����.�w�r��G��X|����ӥ7�
<`�"��b�G����>����I'�jS�E��N��x���`��-����_��:�D|��H(h|Wֈ��{;�ʿ�<EtZ�U�B&��$��	kz�����t��Xe__�ڗ�p��d��/h{G�U;���qQQ��䀽zL�-bJA����Wa�1�����\�A���~k�S�^)�{LxR~���ݺ�����/ vr���W�9��#�=dy�I�&��ѵ~��l���]��{('Բ^Q�\r�E�����o��0b[�󬡬�����X��<pyr��O_
��TdFJ�nI�N>s>/}��)k��t"�vK6�xl�>�M���ʺ��>��������$C�P}�΀�s���3�N��뜳�e��=�����N��3�Rs���7:�}�,��<�������=V�]��:k����.��V&v�aZAT�X��9��g]����v'�#��rǹ�gn�S7겪��bjϊ�&&<�g��c.����O1�6\Z���d���r-��u��Ȏ�����5r�\&�o�S��x�[)e����Δ�V�M�5ًe�EQ�o��u�w���t�H��Z���'e=ޮ���nwg㧃�mË�ʎ[`�y~k�h�m��\�r\u$�T$����u�&�G4��9�Y��G|o�BKG��f�4<	�S�\洲;b��Y��E��Op�"��Һ%�۹?uzm^#�܏�<ҍ�j~l ��������k�]{h:첰^�l/9A���Ĵ"lt����^pn53��W�e�-ȝ�5���%a��"��匬jv?�%�<ܬ�B�h�}8�Wt��X�f��.,z=<�72�v���ʩ4�>��z����/�r�{��f�%��|C)��}���u�}Q���c#���x�������U�ϯ��p�ʜ�G�i��n(��C'�G�ч}�hC�����w�Q�j M-��Q]�zvD�
�'b텝��k�{H�v8�<+��Hg�6G{*{�1��s�!ˀ��q�G*�����=�`�W��]հj2(�U�X�V5�H��6����oB�_$�D8�V����lp�������:��3��N=>��~�B����4|�����Ys���nG�R�9�F!N�/&=+�e�W��ǖd�<���W�O�>�$�S�Tv�ׯ0�SV#"t��w�~<������QI�J��܋q�s=�į�q��LU��zx�>�u��.|)�;y�]����h��Rv=1a�A��*������ LwJ��b<�"���%��֦�{�Tg�z�辿�/70e�e��v�����<Gݓ�Zuzu��+t�:��"_\�������J��WJ�r�1�p�O3.TCˌ��"��q'd���F*wpY,��{p��.I���X��y(���I6�YC���ٝJ;;E�53f>ls�fA���կh]��o^C��&��c_�#i��w�Ft��w*kQWp�+���S��������qy���F��3�����zw�K��tX���Дk���������+��ff�a�W�����,���c�p4A��D�i�k�I|8��{�����i��3Rr��s��V����^����ؗ��]��W���&��z���K�r)��j�bw �l��6Lɞ�ӽ����X��'����v�Vk��U
�Q^;�GBxI�F��f�ޙQ�k&%�P�(����Q�-�Y�o���R_g�~��|��(il��l�r��As ��/��أ����-��I��f��A�7���2��L<��b5�����3��1>|�9��֭��Uѳ~Xvr{�y����s������pjSI�.��{���O ��m;��Z����l*M2�����e-��X�� y&e�L�x0��i�"��^Y��gz�jw�:u�ʲQ���Ϲo�k�]Z��Bq��=��M��>�A}���]������Z�?P����x��U�!�IVZ-}��5�>~_u�P�4*��{�H�D�#2��]� ���}7�
��=�ռG������y����߹�&"ɩ�_Q:5J/.�xt�?}�k�\Wb�_H��avn%�#�rz�W���p�s(��K���b�Gs��������jڶ`�ʽ�4.�=S�w;sG@�R=lL�of%\�*]��8�l<�]g���tK�-�U�ev��z�0�l�ӂ�VxMU�]�jE���h�>[�W�M��%�Avnt	G�U3=wc����ȏڮ �B��/P��2��V�v�o��d���TI.��[����Ʉ�i{���۞&O�"���wVe�W��Z>��Rz��}��2���5a mM�F�3 ��?`�u~��d������;|>	{r<a����Vs�T��4ugmA��{>�6K�[~���~��otץ=H�d���ht�}
�;�?��K���P..�%�M\N�[N��n���' �X�UE�+�=Y��%�'�4{t}ye.v.9�����T�՝�s�Lum�=��ޛ�廐J�&���]|?h�G���LL�!�g(u��	�@e�yV��`\�⪅���>܈q��y�Y���u�������
3��~��WK��M�ъW��j�"��%{5}�,U�{��6��i����l*M��m��_LӽMJ�z�Z� �B����&��1׿0Μ�z�d����0�}mZ�}�=�X���hW�P����}�ݽ�\�R(�V�碄#�R]���'��[i��>2-��s1��"��wk=�F���|Q�[k�u<7�3���)�$y,���*���gn�}7��X��`w���P���k]ɮ;J�oy*@�:e�5���ٽ\��gs����ev�pV����}03�k��rՑ_���c��әv��Q��cV�B�����3c��9b���t��H����Z�G�o~���
j�	��3`�!Vζ�m|�MfPvܛ�d�:��\|�{�k�n�3&7�2��N*]�5�4�+Yt��/��j��3���I%�@1$��@���Ib�^��te�K�V|��qU��CY{)�OϜ�07+�O��wY�R��87��m�p��F�{��O^ Щ�Qe�dV��=�y�9y�(3qCA2�#�Ó�:{� ��T'�u��c�)=���:9����r�;�cިq�s�	���8�6���$��uW:a�be�ϓ-�W�L�������X��7�A���xK�~�t���;�co�g��k�h�{�6�U��қ�K�-o�Va�5�;���n-'��_P�4��"�]z�PG:�id#U�(䡇��=^�vg5́�C�6p	��yn��9�z�31t���v��CE͐�88=���*b�NM�ϒ�@�A��_�����ڿVޤ�,�ͫ쯐����!������c�N瀬��/�T�VY���y��i�5;-u@�V&���S����a�^(pX�hxL���������N��	�Ԇ_���W�ƚ����yݸ)�F ��eJ��V�ߊ[oA����*�)_XgB�&��j���c���q:�T�GR���A�Ȝ�!�=}i`4�76����#��}CVT&�%��qh��W{��1���l��5����N�����8�7\�����\ {zx_H��yb���7y#� �6;N�Y4�sU�HQ<5�)r�o�&�]��zI� t"�.�kAo�[�w#��;�莴�B����8�gV���^*�*v���!8
��������a�wvDݽ���p4)N<����R5v�Z��I6ʜ���wR�vŋ����Vی�W$��Z�C.ɋn>e7��ޖ�%Ҙ�@� ˷�r��X�D��:����w��f�3��v�V����:�	G���]����B��۩�[ѱa4ۗ���њ'��!J��Vܛ��T�Jw���]^�I]�k�K�/�Y�ԗ6ٽ8j:2�w_bڑcE���u������{	�K#�Z(�U-���诲)oZ�T3VM��mE�m��K���S%n�P�Vevv�*����y���*xy���:�`U�Oz�k����nq�T}j<D��� �}��墄,�c4�':��j�f<��m3�T�!��0V��A�Y\���X0�-p����η�ͭ4̘¥xwt�5��9��5(i�� ���`��=��g_���(�۲�w�6��v|�b��G}��y7�z�8f�	�[���ww33�s�l����Xm�(�A���dC�O��+`�$�N,)e�l�*�ۮ��F(�R�� "`��W����.?7��(2�c��\j<����9mIhHRGDC�Bm���GkK�[D��M�E송͖s�����{��^PɊC2����&FjlƑ��6�o^�lD9oRm,e�vL�x��t��f�
�[�F�Zt�H��e�$4���q�n��)a��N6�D:�x¨R���K'�w����/v�v��i��=CEJP�\��9eR�k/n�m��wZ�i%�5�o,�k��L�Xv�gq��Ţ�:�j�5َ�
y)a.S�!|dH�˥N�e#mes�$ep|����XIm�Ie=UPM�t��e�h�N�d){ڨ���n����S"��2sK+�B����UՆ��6� �0�G�}t�;k�!g;T�U�vu�58Q�\n5������M�4<�N�Oe�vJ�[z�[<:�n<c�2]�)RSR��c�ĴY؞@P"�H���)�n�RFf��5J�Z}��P�h��gj\9N�X����3�aɒ�)�Ј![��`+ҡ�z]Љ��pDM��Z����B�������1Wqs(�Ղ8Mj�.��l��{�N�c�ֺ��TY�U��Z*�%M�����Z�O�u��۬�0U�
����Wq֬h�oUٽ��1	m$�#��ݑP.Q�FI��N�"�}��+�������!�t#"�˰[i��@Ӈ���ҝ���4Ke�����H��Q���{59���N^��Y-���2�{��k7)ܴ']���]�3 ��a:��C��*��l��9�B������v����`�K�,�-���:�6�!m�Z�WĜř�{���.��k�Kx�2�t��q� ��\^E?)���݈[������qq�[�H�E��k��{������1DV��Sv��pK����(��OmR&"�;W7+U��F������]b\��A]?����j�{j�[��3Z�̣��N.w���g���y��m�#%���vZB&��H>k2f��r��Z��e��s�25Ϗ%k|[I�S��3��S�/�{)�۝[�b&�Z�!WL�#�ȹʷ�XԊ�����T�8�s���1�[c@G����@l梟��ؙF[����^��+ւ�˄�uw��V}�P¨�Iz�[O}g�#Yz~V���X�Ud_om{2g��BHs;,E���Q�>ێ���'��Q�$X�%5� ^�mo��u����O_��ޚ����y��
�^�$l�i�SN<�N�IӠ�œ���[�m[������⹝��ܲ��U&-�ND�̑G���d�K�j�������z�M-��vꬮ ���/kc��P�\�ϕ��f�<��ØV~�.�9,����}�x�+N��{�%l)�Tsa�( )����t�G����$�Co7wL���Lu'�dH۟M�;�=��蘄���3d�7�����A�bf�H򙘃��-e�ݎ��Oѝ�u����*�ߗ��Z�,���';SP5�E��o(�Wԭ c�{>�D�	�yx�m��Pϼ�f|n�}���?�����T�?�l1�j��y�*��o�>�Y ���j�~�2����:GC7��jX�*�������'�l��"/^��;ǣ^qT3�_x�vX}hh�w@k��!&nC�(B�k�VC<-�Ā��K�����#�s��V`*=�o�AN������T���C��(@к�{]�= ��j����n v�F8-�oݍY���BU���&�v�8^��-�rt�N_3ܵ4b!U����xA��K��p��j[�4+lN�5� �I�D�t���.��Rɷ���Ko��K�C��W�%��;j(ʒr'��2Vѽb��τ~4�a����);/��.��fm�W�~�1����9����G�1Vn�Ӈ����c�R����;~��KPv<*.wj~��̬�F���G`��r7yB4{���g�9-y^y%��==�r���yS���e��v��ݶ�~~�Qߚ-9�4�GZ�b���xP��f�s݇��㥮C}"|@��L���n�S�xu>��R&���;�*"Sl��<�GB�f=��v<�n-�ݰ�e�ͳ� �`΢�h���R�0k��Ŕ'�Ǭ����f�}3�=u�2�w����A9��vbrr���w��cօ]OqѪ*�خ�"숢��<�`���r�C�<3]�ox���oE_w��ņ���̪0���6��d���t)�TXt��Z���PTM$�,���/�hw5�~��_`Fj}��g��%U��n����qkWs�񨹝���M-y=ݤ�֨�+��Nu��N�����eK�j�E���:��|�Ι�O�d�B�>m옠<���W��~�Vu�����3��[���`�+o��xS�E��/1O�Nϝp�!s4�i�_kܣ���#>�&����f��D@Χ`�����5�<~�!�#����4���ٛ���Չ��/�;��AW�L�\�����\��9ߴ2W���]U^�5�{��	M�|��\�w^�rZ�+޳2��q9����B�\��u�"�5z�}l�X�0�Y����+Thξ��[�6�m�5ib��u*�z{�~p�Q�WQ��G������ݽo��l:>����V�).Z��ƛP޼��j��l�������M���Ǵl�tj5��^l��Ƭ���)[��ؼ��3��6����+<3ƽ�H��TC!Ujz@O�#����ż�� ���ݳ�����[�Hg�R�8�ߝG��.�9��Ő]:d�+���=;�S���K<ī���~�ho�tu�ũ��lz���)+�w+m��hM9�q��ɷ�-�&/���.�vp��WD�4��M(J�<�sٹ��+�jД	�gsV�4:I�"0{D�t���l�M���"��g�)�[cd�[^�i�Y�����ڟ8]s�4�*�4�q��,���xb�X>�k��"��K�v����[��a�o��(W��-�X��m]�;��p�6� �d��o��R�]]Dn�eu��HO�Ɇ�{|��e^w�aY�62�au����;��>7*Fb�E���Y�.-�CJ>˂��~�xO���=V��	��z2�@�p �V��싴��ぽ��`p`�]�sBH�E@9�zP�}x���x)�������9ު�ܮ>��ʉb���$٫�z��(L�>־Ys�{
+R>*�3��ǧy�F̒�,�H�� tђP���q���|���Z��{��͞[�Sry��>�9�g�������ϫE�.]�(5�-,�yl�Ml.���<Fv�	ZڃV�,u�;��]S1�Z��4���,�%l�$ ��O8"���ɏ4���D*P��w�r�=�L��o��%���6s�W���us1
��|/@��Bq�=�^��.=�ql���e��۞v���Rz��_h�Tȟ`و������O��̫�5�5>_{Z��r@�9��z��uX�~&Oܱm���G4tP�b�)��	�)N�b������	�.�a��>Hz�Y+}���B����g"��������9VNͩ�ثϼ�z�S>��8��>�`�_k@���}�S`)�����z����oGt���ڷ�d}��mӾ�D�Mo�L�v��y�ǷGQ�+��C�%9YD}9��%gـ�b|��^�X;��Ly���Dne���qMG�^O7[����wy��l'��*h�.�]��[�qΟ�^f��R�_����]�n����*~���~��? ��#3�L��Vr���Ϫb�Ҧ������@��9/T�v~�!��.�To���@��s�����Gw-C�.�{�r��Q�┇�t��RL�Ҿ���flq�W�aFígXO�!�>���"U0���������o]��&��[㋆�!���L�j�yu)�{��_����w뱶�7�^�]����Q��c#����D#��X/�6ʝ0#�d]��=R�J���,�/Os3w�C� �[�8�(�.�,���-�m-P�;�}��ވ 7j@��M���0f�s��*�h�T7|��,-L"��.�!��[�[i���W$�5c���Xsj�qGkH�@����u4c�^:�\q��w�eM��X��h���Q���EZ�\�7����Ƙv��X#��AT�@�E*	��-r����2��������
.;)ߴ��|�y�1Q����ϭs�b��G?{��ۏ�:ֶd�����&�����^e���(yg)T�<��  �̑8�0cz�KN�N�n5h�-�$騯Jv���n��ت�\V�i��}q�z���j��F�n"Q�{�"qFM����h)���;���K��?N�6j@�	!_{<Ի��4D������_���F���ٕ��/�:�^>69�f�mm���3Y���0}q�z|�@~.���/�I��&���{��Cl��0m?�N_|�_W�U���u�FH�������7�M?+���%�u��g�F�l-!�3�{��\�W��w�=Q�.�C�#���)�fRfK����mһ�]��S�^�Ͱ�%/U/�<����"^C]e]�;�{���ǼvY�eeB�cέ1�O-46]pFd5�zy���_A�V����]�t��SE��lY,h�?���-tV�d���NL�����-Ë��Y���m�w������t�Ǘn��T�en�£R��X�%NSYW�����Y�s��jY�10������b9t�&)	z�zVz��ϝt���d��p6����C�߶�\���Ԃ�ě���A�닯mnC3�
�k���{R���粭��&��z���5n�6�fs�=i;ڛ7r�U/{�g@$�����ћƣ���1���������<ى�W&�$�: gF�K�����o��˿��M�eW���tF����g�Φ=^��<�_�ZڐOJ(aʶ鼬��
��.�G�����W�͗p�7䟝�8�j2��LD���#��:�y��R��GviM�a;]��_G�C7����O�
�fz,�^�w:��� �E,�z�2����{��e{A�9w������� ˧��~�23�Ee�e��\��e:�����Q��|[�
M��b����K�d����fID���zн�ۺ{�R3�
+�Ǐ��<���.*�_����뱠����k�m��b�0�E���4���|7��;^�E�T\sl�/$�0x߻�קME1@�HR2���O���A��箯˷@��Zg���[o�7��F���T�6�u��E���I�yPR����Q�>���E�UX��2�o�˿z�>q�Au��IVϞUƒ�H��/�͉��[u޸ݿ���}x�\����;��MZ��,s1���Rb��z���;��^}�
��J� ��Ƀ:��o�Ⱦ���Q�p��Ŏ�A������OCZ�]_C���ף&�1^:DJ#�����:cÉ|y!��=X6�yT/�E�;�qL�����CUܟ�̗g��-B읬�s!2g0k� �Ҁ�\���k���Q�^��5�%�1���˰,��gA�)�Շ���+�f��<���=|��=��>�_�}=�ӄ�RQs�G;V>[���`M����WVqw���HRLۧ�S�Bn=�$R�>�=��%=�)��,W��:?e:g�D���\c�=tBֻwTC~�;l�8C<��d���]3=MnY{�7��Ҭx�Ιi*��Ժ�먹���>��t������#S�Uc��1��~I��sP���q�3>�Zg��*������.�=H�p�RTiP
�-aq(S�j�h:R�pMS'�?ww~��vY�roV/xyr��~�5�����55���Ǣ�ƶƆ8,����T�+��Iy͕7��1�}3��#<��E��B������,o2�NS��ڈ��V��~���4�/p�R'�3�ϕO�{����ew_nlz��(t}�Ƕb�^s�����ܻ����**
K�=�2�8_׀GC�s[�Q!���
��y3�U����������w_�꽸��u3Zj���s��157�������#5���^N���F�e=�Z*aTD��������4q�;͊��ج�EǸ�5��7��g�s	\��udM�����|o�^H��3�+iW�Ue����C�
��.��`{���L�t��KM��(�d����g~T`��[�#yp�Ƞڂ�������Jc�-i��l�+�P�OftYJ�wm�Â��nqѴ��5{�B�V���X�Ǫ92V`�ڽ'��lTn�y{�O)�ΓA
�[�/M�7�����Y3��]�D�LoK�zU� ު/=�;{q�M��c��>���ːhw�`������4�ofI_��Z��rL�|@Ǯ �B��2��SmSR��zÞ���Z�=s��oge��Ҝ��-eҼ���&/5Wz�qƞ���Z���m3[��.{��Y]h�P+�-�}-���/%�P�j����r�뽍���T��=YȻ2wӱ%��+u�or������p�||��Ɓ�徿wA�dy�v��� �O'6�F$�"�vM���/F�f���w9:w��=�L_�#wm���P)��F��[�3��{��ɗ�^��nWޞ��C�y�$<p%ϩI3����7y��>�@�9����cW�p{r{��f}q��u��=����۵��s�]�oʡ{v��=;k���y<���{�n=���E>�O��ɀI�t��C�s�^���M�>�׶1Ԉ󏦝�}�n�=��&���Uy�YН���3�4/7������8�ÉU�m�xFk�������c��b��$;�7�%"��/ia��B��K)&�g#��Jx����ŕo���Bt-�ùW;Q�j���rk˔j<���[�|�I�>t�s}�����3�cud�y`y<�M֜��p�q�iC���%�U0^�1��� ��T�a֨J
�M@ O��ʘ�PՄrN�C_���Rˉ���"�S�Hg�_n��=z��o7	8��5?�K��2�V����bh�t$F�(p K�Ptz�פ�a�4����=��������B;L�)�N�?��³�v�ʥ�y���}�tӏk�g����}.��K]	�����W�1�T)}����t��Y���)���Q}]M�U���}��Z)ہT>�K�긛�����S�jO�jg���H���~�Ɩ�kR�U�M"w�%4f_M:Jg�������3���͗��z�v����`���u|}D�s3��L�=5�G�>��*;o]l;9gv�><kwe�Q���|*������SC�y�\}�����Ϛ��@?A�!�*��L��d>)�f�i�����:��dB�a��US}�;?X� WP�O�/Uj��*�}���勓�{�z�1���u�@��G�xAaf'�Lo�a�t�̻6&E>T����_�**ڄ����zt9Qv�fq�r�������
�»^\�Q4A���EZ�����1^��d��g�U��i�[�'3����$���T��x5�AV3�m5t�Yo���#���^ZϮ���xT�R��mW�U��\�8W���h&�9�G��ʣ�M;�\���QJo�/��x&tDz���[wA�oњ(l������J�Ė~w����^C3��Ϙ���۱-�o�"��q[焮q5�Z�g�dQ��
(��y_�n�R��vR���R���
mJ�]v��=,�7g�;�����K��z�p��C�Ĉ�/B6���\�C��ͭ��w$��Te�f��V��9w�x�Vך�G�P'�S������������k3�Aq�/�6�?J�9�Î̛~�WO�B�U@��z��S�������t��gH+�z���u7��}�P�o�����S����cܭ5�|ja���s*�)>�Q2:f:{��l#��Tx�G�#ϯ�lB<�ۧD?�9��N}�^|�g/��B��
S�c��=�0ϕ�8�z������D̩A��l��uW;���=Lj��q󍎛�[�&-��0�b�X*��~Katj��3MHT0Mo���Z���+8��������#��%Sֶ>͛�I��Id/�9ž���˒�7����ǖ����^Q=�]=^���["rϓ�x����L}�p�f���9ӏ�Џ8�>���t7z�S����\w\�7��'�#{�CH��L�ǭ#J����`��|�o�#y׫#Ҙ���^U���즽�������F_����}�0�zyd����z��p? 7��(�>>�j>}�uO�hp�B����d��䋙W���n���Gǹ��[u�����Y��;	�&�^*�[�zP�{4�̍�#����lt,d��v�jbj��d)ʞ�y_l��r�;.�-Z�3��aZ.퓬�:p�����P�|6bsq����Һ�9�j����� ��O ��=@_;��͠�8��\6MG����������>��b�&��W����KJ�kUs(j�>�T�1����p�C�c�.,����Ch][�#J�k(;A\Rq)6�v�0S�0
,�V7�c�XÑ5���&I�`�]5����]&izQ�� ��Ws�4��f���B�7-�Cn�!C�=j]^ҽ��^j�IŇ.k=��$�w��N ��9U�3E�!ʾ�w&J�/�V�J�G���J�s���K4B��w�a��՛9��{��d`Q�*aɢ�T�آ$��I_Nn�VEZ2놪y]A]�N�E��Vٻꊿ�]�{�����;�~���e��t���wmt��ш'q���ݡc��\ᵬsռ�;X���:��!Ӓ�� �Z�O��Ն��M]s̻���[�©��L���zJ��5(l����I+̳Roe��W�!h+A�+YXCͫ��;w��</F��*c;I��,�U�Fͺ��ɹ��ڬp@nQ�����
�h]�R���QJdؐ��X2���6ɭ"�i�;�eN�
�hj�[r�3����醌 7�k�]�.g�ɳ.f#�;Ob�<' �!�|o)�F�����ʔ�Bv����sm�$��$ij$_��z��uc���&���fi7t�h<�F7kx�I�]����٥oh��lqFݚj���J�LrT̤jVWeFL�oi�7K��	���LceDRP�`���m��]�NS����c�3��u�.l�,[����;V��냄�Plc�� ��|�溭��d��u_u滙��p�c,M�r��CT�M�b�c��f�S���R�^ʼ�r�PH\��v�m$�9�:i�U��/+�o�f[Z��b�S����ï�����u�!SL�WB�X']36��;M�c/zu��3�\�\�^.Uׯ��=��x˱̪TkA���"�����&�W�������5U���L���x��r(�C�@N_#q���ְeg=;gn~j��Z�RK�-�/��]����Խ�|�δ��m�*�l�����?��`z�N�TZ���-ʭ޵8;G�:�����ۿ�ì`;�	��%U�{)�6|i��)�n��6���5G�2`/*���;�ӂ�÷md}�i��Whgp���D%��;���ϐ���v��>��Z���:ԁ(L��c̶}��^��131��G�)N������yG��>Kê'Q`�>��H���F�.o6�>ttp\�ʾ��Z���pG�%�[��DT�?��^�����j���}P�E3�[�F�b��]�'��!�B|~��ܺ�l��/�ZRҁ��4}����Ip:6R���ǟl�I(�7+sk����ٶrĪSL^M���$@7��a�(yP�&:=P�rDU�}^Ȟ��
ф�����}����/zA���u��qm�b,W�j���/�VM��Ji:�|y,>��矧�����_k1�h�uX��H�+�^G�N��6��E`��k��>q漂���C��~� �3���3&'*��}��މ��w���5=�R��	�v��0õ��wI�&o��v@f|_^m��*!ڻ�Y�Ur��Pos~�O��w��}1�+��7E�D{ (���������ٓ���O�4�,	��<6�Y�9	��4c4Q�c_��]�-�Լ�,y��'&è»���-�������'k8۾��]��c�֙}����sq�mL=�����^Ya]w��k�M/�¹�J;�
�~o��]�᡹�*�J|��4�𢶻�����焸7��c�/R1V�5 ���u����fv�|Qzg|�_�s��6�Ҍ㢥�}y�z8뫁*`R���H�R���ԧ��S��S�_����r�{�UO��PIW�|ۅ]�0k��k�϶6��P��dW7���ӊ O�V%�l�?Uҽ���'zw<���_g��b&���Y���6&=���t�y�fjLC���c�Ϫn��{7����O�{�`u^�6�����n���ⷅ�dPk;�z�e���΂�ǧ5�dρ:4f>�5��
_r7��{LQ��LVy�2��	<��k�I���r�0}��E/]���1����ھ0��Nz�g����E��
?s�?{�OUy,u�)�ӕ9�~8�+�x^
�S�!s��k�|�^Hb���+��^ʍ�\y�{�=�&s��k�d�k'��Eu2/Fh���?7���)Z��c�ce/�8Q�~�%{o�X������������կ�v��g�}S6g�»Lf@��y�p�ˮ���|���E��g*��a���8�A4���+KTN����ed��g���Z%�j�(X�1��4d�%B�j�^������,�F��*��c��
 �i���۱)��3��$�w+sDw���7t���f��ړ��Xd;"��H�L�g?���
9J86I(��r�(DG���a�Ujǥ�N�)��_2��3$gt���#i �U7&,���+���ť����45�vZ�b���nJ2
��2��%� qA`�>�2�r�/O~pz�<��|4�m���9���M1��>󙫞WƶU�՗�v���E]�x��r�g�\|y�����+$�P:=�����K���	(0���?nL��Ƚ��׻�~å���{�-�v����2�ZpS��5yC��;�:-�o�w9.���	�<�����,y'}��OEG�s��l@����]��nM�7C�*R-G�*�z|��|������"�?[ed�������v=1p� \T}pp87S�.�s�7}c��s���I�K�d��#���ۋ�r���?/ڊ%�������_;�O+h��e9��{��M����X��#�s?xi3�J0YU�j��!���y)�6߯2�����p���1�9�PHx?:�2c����㘑~':�)�1y�Ǟ]���؊?��{�����8��[�5��er�<p_xゆtx(}��id���R[K����eQ�'QVG��yR�H���-�E	T�%x?��wk� �Y~������o�ͱ���d>�q��u����n������G��ov�w���돣�)L}l��n�x�Ǖ\�����i͢���-iN���*]zj���ݖ*8��1�_�3wR���ǷJ� T�����������h� u���J�5�K�ۂpR���ͽ�ς9�1+�g�@IJI�*_a��β��)�vi��4"#��o��\5Ub��+�{��f�b�ݽ{!<�����ss䄽z����ԃ����n���+�Ӽ�����x�V7�����:|c��[�� A�����qa!�^Kg�ks����ψ=S�x������ZH���4�ziC}]�����|�c׃�p)�u��#�{C���1�u�ى���P�"R����-cѬLQi�<]���'�I��X7}�-���$_���[oG+]�9�S�k���nl��o����>�]/��%G�ߺ�n7�L-���?|��c�ExW�~E�'2��D���:N�֣����\"];
�g�����+嚃c�_�o�"�-̜]ѦgCR ]P�թ(�q��<�p��QD[�$!i�ӒA$��FeCx��W�r%�O�H���؟Lg��.�����ߥ �N�x��$�/��7���؅w��ڮ��������Ej���� �2�{�Ӆb��ޫOf����a�~�y"�܋�ov�0c��D��&ct{�t{#��=5={9߼P�����lP=wmo�Y����\�e^1�s�q�X�v��Q-6s����������*��:K���q�b��:h��4o�[9(W�����X�>���ik1�ܜ�/^T[i_TJg%:�_����	��^_�� �8eGG��L�Qn\[!�2�CMD�ދ�%��8m�a��6*#Tz�������n��{��w�;%D�yI'��f}5����&�OH�f��{&��<�bj��]y��Ed����8���"�3��:=I�I�j��8�Te׾���O��u�\Ѭ�هO��us���5lVZ�u��y9BA�:-�Y�QQ�=�Q�sً��nz/���� �ji�e�Ϸri��,F����Dr�VDU��:<z�UX�t���-�d�d8�H^Ip븊Q��^�呔���nH_k���$@�@E��/�G��mފ���e�Tv��V�>}Y��(<w�et����no�d�x��33����8t���<��z=+Ǘ��������A��W���}�<��U��,K�x�X5uo��{|^b���g��M3�1�ߩ��@nκc��>ۢ�Ճ�Ȟ�y��ZNhC����5*��-؟�]| ϟ=���~p� ~c��3
&v*r���齗��VS��}�:z"��8K��-�jq1��z<R����@��_T{���铕�I�O�w���W0ǳ'�?$�}�*QwX�#7)_��w����?fQJ1�˞b��P�t��]m�ҟ3͐���R�a�*�@���,(��U��=��y�6Jk.�����u3�5
{EjKf#���H��`ۜ��d���+�c����1�_�����]z��X�������)��e�''��i�����YhG��'�W���^^ @r
֏�y��&�������~��N����f�fhc����R���Ӆ�s�b�c�]g����{���Q�N}�Ktz�	�Uѿ}cmk�ni���	�C��IC���K�f���9����3��>�#�G�G(�Ts�b�|�=nV�����o��=�2Ua�gcu�R֟nR�w�rj�����v%�Ig�>h(Og�S��� }*���eYd��~����g{:�46���S�O���=_�y�u��iB����}�x��S�t~B��~U�ֺ,�>�_V��W�u���>��D� �W��ꙥ�H\�s�B�g��ʩq��1�mtE�����zȞ��NNg��ꧻձ�p�5}�+�(~�mO�j7}��Nn̍0'�_c��f��^fl�o`���9=F:��<��>�u����dy�����P�{���
ާ�k�לЪ��k���j���E^�U��f8jݦ�q�ٮvr�TԡY�w��ir^��X�����yf�H���۾N*s*B7y"q�\��ӡuQע(ቷ�s�\��}�H�������C��V�D�I���-(e�g.��U{���r`[嚡����o+�<#+��y�]��;K�M�ӌ�j�.<��ݰ�Xӡ\���`'s��G=w���=MF��cp�!���7���3X�X�e�ƺ�ώ�_���6�}�^Tj����
���d���M��m��(�Z�%-� �/�iƼ�^�7���욎��&�8�V��L��y�}>�N�/�j�n�H�̑F�P!�k��|�)�r�:�
3Au�z�ۿL<���X���o�&
��{���N���8}�,J��倿1u�/;�9��e�{�����{W�(���9}C�,� ;���*=����y������5�*�R�&�˺����씅�oʈ����IF��z|"��M�\}�Q�n���s���0n����ڀ�����:+#��Ͼ2?�P�O4�V���묕�����R��!����9U7��G��U�2iMǿDuO�?N��h���	����"���zb�]uv���H���^o�sw݃��T?G��ڻ��ƪ�rg�Tjn��w����%�n�➁]	�WS�Gl�է�hľ��~��p�CT��<s :�ܲ���iא���V�#򠼨{!�!P��y|�)�SO����Ϲ��h�����-Z�Nv_±y��}����ﴸw޽��ѽv�IZ`28R	iJ�a���&� i1}��� K����ie�W�v_��V�^�%ǟ)��z|na�|��� �Kٔ�����L�K̙Y9u�}��TWs��fv��O��z��E���w썗��O+�����~^X�t9��iчkzCU8f�l8���������^���nsRÚ�}���v�'M{\'[�t�aY�7��VF���n�6Mv��+X�Q��e
y�=�	��t�m�0������9�����_x-�E������Y�x)1O���Q췳�hû2�wUG��R��n�y���|>���{��E�Y���`�����7�5[��.��c9QY�f*�:�=2�sq�1�y-`��3����|�Q�)b7u��\~��j߭oZ*p��b	QڟS�K�~N�U�ݿ]oE��?8��f�|ǕGxk�ϝh���~b�����;ޗ�4�T�ͷ��!@��w%q]:���O�����ZV��_��o��v��X�[o�����	Nv]�߶���k��c�w5�z����ŕu�N�=����_yV���']���ɮ޿^X��
�CfU�&$�8$q�c"�P2���l�8d��P@ׁO�|2&^����;'"2z��>�H�x!#]���{> ���}v�}�. �К��oP���xOb��W{ALT�-�>�J|5�+}�֮��}�S��n��/O��YIVv�k؈ˈ{�o}v�x�S��/0�
�v	����3�~n��v��"P9��n﷢��dQ~�J�>��</"�dG�����[.��\{�d�mM[�sF����W���;,o�é��j�kj���5��tqc�dfm�mdn @�h��Y(�ǻ����]7�,-Y뫍v�\K��r�2��>㸹A�R�a.��'p%߭���Oz\b*̄��Q^�{��V�mDS~0�v`c�F����#�Əw��495�J�p�������6���nOR� n� �xeb���1��*�8O�ǥd��OE)W�hkV�Qo���=|%��x��G{�	j���κB�w2G�0��u�=R��lO�QV�X��@G�8G�್$W2�1"̬�z~��M;���kљ���<	���kX6��/���Ywۦ>ϧ���6g���y-�]/��"`Q4��$^R��{X)i��z�#��k�)Tȫj�ȹQ�`���kTj���}�~�Ð̫Yяk}����zy}�Fޛy���ӱ8��	bK�}w��Y�h���]�'��=Q��������~%]�*S�M{R*��vG����Z#��ҐT{+i�l~�"dN�{$�kڶ�������������J�Uy�놱�W���1*|r�Qq��K��ea���fa�{u��W�BÅW���YW{��
���U�y�:�����lW���΢����2i�]��Ë�|\)�����u���n�ƱL�yx��^��4D��iO���b�ˇ��s��G��)K󼥲���W�z��Z�vFtޖR��ًE2�}����U��f��e�y֛�]�"ˠnF���U��u��Y�n���L�0�[9WR+��8�%���C�"��h���7��݊���������7�GJ��\���ˋI���r�/�#�H$��>�p�z�]%�c6�u�E׺1�:hM7*�]Z�{���~��Z�yq4Ὓ��u�Jή�먮w��.��^���c;����:!��gݘp�-[U�T���j$b�qP��8��
��������lmum�v�F�J�g���9ͼ��� ~]���i���h;�������x3L�٪��7>;q$�Z;��>9~1w�����E�8�9��c�*�:����M�~;�ϕ���w�@v�EN$�Ǵk�o9��\�@���y�s��I�T��r���^{R�֜�`�!_�[=P�e*ٮw�~�a׮��
��yT�t<q"|*�M��X1�2�<�%oҍ9�q=
L%����N��B�Չ~�㫢|�爯���V�V�u](n��o�Y�ϜM��w/��M�����=Q����^��7ڹ��A��3��/f�=~�Pn(�"�,��{�<�fA���&N�^�n��Q�V � �'�����Oo�n�JUT��UG_QT�uA~�c��Rw�n5�V�{( =�_��_6Ed������xy�)�L�S���D,�߲"�L6�8��tgk�ӄoU����Үq�sA�8�Uh���G�P��b�X���jw���bGH�\�W4!+��n�p\�"��r�12BR�D��&CʊI�ӡO�sV��Y�5�X���n+��ui�q�Y�����:y�@��Pѻ�V;��dX�*��\�+K�ꋾ�B�f��od��D����}Hڇ�)�q�����VvZ�c]^�bG)��2u��)�V�;y�x�d��ћ���Z�lb���]�����EcQ��m�m@r�3��	g$f��#ٵ9��S�EUؼz��:;�Be"\B�����t�;�,I���e,�Rpγ���G����?om�b�9��z�J`t-�k
ˊN�r����g4�n̐,�v�S�,o/��f�f_Z<���ư����80���ۉܺ�(C��J�t�f��d���5��&���	�@d*fe�[j���
�f��L���m�ת������B��z�;��
 >���Mw������}�f�[��j�b�ʵ�:sgv\�!ՠu^q�;�Im��G��آ@�|�.�;Y{�ݤ�Yn�����um��"���1MAƴ���ƁC�-�Wp��[��b��NӣTRu��S�J}�w;ծ��]CZ��$�n���]ꐞ�R�iBL��L��n����L�g\��nN«�J{�����f]#w,'����;��1ta�X&9����-�n�r���n��۶p��F�M�+/	�u�y�G�6��(��h��D�U,��B�u��v��R��bknZ��?,jX62� Z_(���Y�O`d��l��k��O^�^���e�ę��h�<͏��Z��������чR�����Y��fN
��5�����¤�pS�ۂ��5�I��O"i�3\:�0w1t�r2ʚ-�cYi8�3gh7Փf 0*82��bn:�;����+\*��Z6��	K�c�)kv�
�6�[�)��fu�Ho)�t�x����5V�ط]y �6)��X��z��d��/涆�
�k�L�U��vL��찐�MR�Q��wZ�ui*D qpR��� :EV�?+�M�P��ܦ2�FT�E�.�T�b�:V[��}}+8f�ܥB� �׶���.]�~�&�+ḇ
����LTGFZ���i���`%F�(�?�l� ��v�J|T�p�\�C��L�LDl��(��ػ���!��:�$��<8-"��TX���%�gs/q�I�Η#w�4v�,�mwB�@r�9� CE�M�a���ea�Kz�*"iH��`J�u����M9�w�S�����P�����֑�	�U>����HRuJڱώ>S'ϵ���)&�PN'4�v��iԈ7�n6�l�3n�M��ed-�V%J�
�V���>�Ab�G������)�� 9�V=#'Ԫ�|.�}w{����>k����� �xۨ��!���M����Y�r���6��u�ɬ��	��N�&��#��^��1K�D�5���$L�	�F fE��(a@_)�����Zb���~�k�X̜hR'�6\�̳�����eV�˥m���s�7W9/�l(.[^���n�g\E�z&u�	@�w��R�t�ED�a0_�8�M�H��.�+�&V���g/â���`w�e\mu�PU$�FH�*㭧�Nv�i3;�]��1L~��'�-�BZ�c����K��qن�c31�[h��(�4ֵ����ǖ
��Ҭ�6E�Y�[T|2"k%�q�Bn���D�μ����w���a*�(����!0���[���*�gy[3�f�t�D�LD�aFy!� 3Rg-��u�鸁"�'(���wA�Ё��D�	%�d����?��3氏u�j��G�d�͟�:@���U?|���m���}����a�]VG�Zx�VRێ/f�<�I��_xm�?N&~��զu�2#ߖ?b��XOx���g*H��:��߷�K���m���.�j�I�L��S9�ʽ�A*;G��J�3ۭ��ڧ$A̚�����;z=�L	�FO](�>W��9��r�����5=���)}u�2��$g< C�Uݧޮ��������z����t�2[Ƞⶨ>�jF�9�l����n��^���z�	��[��?jL�kV)[���h�^̚���ld�x���w>����Q�5l��n駣N�?��?+ܩ1~�<�2���yҟQ���V^x\��9][Y�O/�p�������3���S�ijB+q�@�o)i�h�2�K�]d�ҟ+52��'R�+��\�J�]ub����d��B0��&�M�
n��_w��n��W��uoU��=��)w�ޓo�|�c�׆:|��W��m אU�6����>�^�CNY[�H1â|Ue�^�"IR�f�b�b2d}������_@_��L���(��9�V;��@|�m�n�@S��֫fK\����l;{/�Q�4ܨ���=].SUƁ�.��F=M�ۙcG>'��9n�wrj;tm]�ⷕ�����pٹ�R�^iMί���:��;垕>��0Յ�ߛQ2tX� ��u��w�`������0)
��l+kR����{>��w5�v�I�>�y؜!����}	����c�t/{1}��؞��K&Ӫ��~�%���F{&���0bJ��� hx�����>�H�fsJ�@�������פ�teǅcG}�ָO�]a����P�9�Ӛj��ה�m�Wu����p�߅����7P�.¾��n>�Ցq��^^�~��������SwY����%�W,jbat~W7�y��`ϩ����˗B����G'����J	o%��oAq�O��%�7��>/��eP:�&��ut���+2"��:��H}<�m�����E�/'T������X��΋����w)��(�CW��}=�cWR^�2`�+�}2Y��^����)f���,]>�9Oﻬ�����u}�+A��x��M����-3�n���a��y�y{����}/�x��uȈG��9Ti��Ԃ��{n�Е�s���| 	�˷��=���5�$����k���{��s��~��z4׾Gϸ&C��ߕ*5�)՝Ѽh�"��	|$wt���G����9ܯ���5��x�E�*�*r0����#��37�t�(.�q��3Y��J@Q����,2�7 ��,�h��9�����)�icq��I/���x1ݏX�^��=��Zdv�{�~4[~�"#�cj�C������|�Ki����)��\�M��:�ؘ�o3ު�yn�)),ts�<#�\�!Vh[�*�i��(]�h���e�Iw�M)�y��(������y8��j����W��x�������u�΅��sG�Y��Y�%y3�=t|�W�M?��,����Z2ES�i��Ђ@1c�#C�烬��;����'*h��e�ğm)���;sr��:�m��F%�[6�S�eH~C25�Nɋ��r���Ŝ=ֲ����`��W��<E�n��]s5����*^��t�.�Rx��D�%�yX>\`��tnI����n�w�m^W��w)������ۚ^OQ������B�5��{j��}=���~)b�%�3m����Q���_���hD]�hC*����[F�>�����Gs�7��G�I���������H�;���uc�ܱm3���y�:J�yz*Ǻ����O�׵2��0DB�1Ϛ����g��[%��5�c2�*ߴ�Mu1:�_к�6[5�{��+��;�>�x��Ts�T�=�W���X�yb'�S���gT%"�1>�93���LL��iW�q�Q��wwRDڷ��,I���V4���;��T�SOj<��ѷx�g�.�{;1�l�`껜�Iʄ�F������|�n{[#�㏾���1e}��Y2DJ��i��˪!���u��򋽔�p���R�.�.~c�>�u�8������W�="�F,ı�u�c�����wyԘ�ש[>0!;\g�~B�i%ةc�<���Gt�����ܷ�t*�I �~�L�}�X���[�Wn;_]�X��w������,��C'�����@�ȭN3~����B�����idz)g>Z�=u��y�����S2��ݚ�k���[���{�]v�Jʬ|�Տzez�0�讟?�Հ�ޓ�Q��o>��_��θ*x��&^��?�EHx�\Z�����R=[�+zIJB6��EvdR1¦�q������9��|.�C��*�����wU�䓞��%����-�s�� bIb�X�W��w�J�?\�P2m���O�3/,{3��}�&�oUmn��@��=x���ׇ4T��;w/�~J|���3�<�y���/ȹ
FD�kh��M׌�2t��둫���G�*B�V|&?��"��ԁg���ȁ�+ع�s���w5���2�U����f&<T��p�ʉz�U�S�d9��U{�� �h���Wݖѫ�Y�4}u��k��ٽ���� o��7Or����9��R�3����]8Z�S7�eY��8�뜜�;sf��v��D$(T���&b�ϴ��~s�93S�Nr�9{ye�	h�!�V?�� �����W1&���t��/\W��<�p,EAX�b�P�VSad�$𥝦.��WJ�VH��-����/<#,M;%����l4M�`��^>�7%�a��v�k�m腤lg��䒏���d	>1*[9+6���/�n�[�O�y���ϕ�
ϻ�A��v�b�Z��UI�Wxid7�.21�͡�C
����t���y����l��%��5�"%1�J=o{�j����&��9
��:h���դ��\X������Gvvįz���X�Q�}?E����u{��twE��+����O���U�y��O��܄�������2e>�QQ�y��hi�S�h�����}{V�ǌ/{>�.+K�-�ª#��oT��p�>������oR�7�XTn����N��_gi��)J��˱�۝0�'(����Ӫ�OP�5a���b���D��37�>��Mo�t�#���q��Q7����Y�.�qk��.i�c�3�õ�!T$$��EꙏJ����!Ox*3�.�'xt����9pt��J��h*�?]gP�ЏX��L�Є/�ʌ��l%��*��G�=1�.�Ժ�3�����;Y~�ϵA����1���}]��Ӻ�����vi�Jn���}�c�LZ���Ml9�+�L����#�W_:D�~4�@��WV-y�m��<{/C\��4�r��M�u�����p�\ޛ��	�s����U�8���u%dїv��5�@^7����ug`/�<<1�v�G6����5CQY�c��o��vEQ��+��?O��2�<��ǖm�:�v���<�)�-C��Sj9���xn��{� 	ߡU����p�������yK� ��E#a�Rk�>X�3���U]>*��6(���S��f��n�6>�S���~�����.A��a�Sf�a�N���y��V���}n���O鶦�|���G�'ʭGp���?Ng&���Y���p��l�pǨ����m�\gy�ѓ���6;2�T�2)�w&�w����Z���]G�]oc�<���W�Q�h�k�{��>鈎J]�_��|�rY��Ǐ��(���8�
�����h�n��M��Q��X�Ec�������u:BO����d�����w�+m���/7]p���������#� GF�J|'�(W����@	*x����"��t{��h���󍏓�Ô�LӞ�}nG5�=�Y�"6+��Y{1�MV<��jUi��w�|��B{j<��̋����P�{���ܥe���������͇/��*DW���! �~OCѷ�3����nɌ��꺌��9�5���1�5}�x�8"Q�U*�ů�e�vwڟvS d�P�C��}hU���V,��Ć��ICX���\���q��v
Y-)�0�	���u�
�ceZ ��<��{z�Rg*��MR��?�&=�~����B0�^�1ꚦ'\�>��|r�>�viogOmT����S����Fy�{��=�c�G%�<���G��I��;�P�K����B�\x�g�θ�����P�>+�;�0���������2D4.�f�Lǹl�ˋ��_�p�|}!Z�H?���'���s���sm9���20���ND3wt��N�\��!�ws�٫�-�a:�U��G����9|0 �
���q��V�RY� a,�����W��f[�NK�B&�>]R�b�	۞�iQ���О���zm3U��������L�}1���DE۱M��rwD�A�f	�}E�1��s��_:�w0�5̑�g������Z�ە��>�l/�(]}=������F��_:Ny�,
C�^�
���L�][݋�o��w/((���f2f[�y�ߎ�4�N�^��}2���8\jި�D�k�yݻĞ����κ�_
Y���BC�"�أ���2���ݎ�7�q�/�<˷��N#��⎫qv׋�V�N�9
b��񄻧���_*���z�IZ����#>��Y��YS��ʹ�u�v��`a������=9�3��m��9��z�k���}�6.�*����UnQi0����F�M��^�o�p���|���$-�_A$3�v�o���H��{ou��Wi��u�d�s3��G�e�O��.��u�K|0[��xz�=}�vC@?g��W�{m����>��X��_HO��9;�&�{8[�g� �_y����-ch��Z����'�F`�C<�*�nˉ����Lm��g#T.�ۄ�Y����;"Oٻ����r���c�Z�5���9YC�^�V�g�y�|{���-C[ή.6�t/�K��G	�R�x�b�O9�≱��1p�Fo��^C��O���<OO�"��||�Tu�v=e:�s��R�r��K����1}�׶=�ÇSg�^��"��yh��a�ж�z/����To]wV��V��b�k�����o/����Oh����|�Ь]���A{���d������N�N��{4�'����{{v��QlxR����oy�B����������$ٕ3$*�Ҧ17��6����Jx����|��3s�����H34���\�^|��~5ֱ��h��J��:ՙ��9m�-�E`�A�ڱC����M�Y�?w����`���|!��m�����dc�~��ّ�e3m��4#����Cb��f��9.���W_{Z�ؽ�mG�bZњ����kw���>��j��DZ�.�����Q?"���Gm!-@]�_w\Yjd�I�julo3�XY�M[K;�Z�|�
|WF�LM�Ǳ�lv8��rEۥ>�2k,jpn6���N�sY�lM��v5m��NT1G��&��Z�kX��^p��'<lAu+�c�s�wϰ��n���i(UBKJU-LU;&�mQE�:�B,7�(������:�7��[�E�}Ml��U�,`w�2�|�:��F}��	}���AU}�g{�-��q~�R�}QgcC�,�n��9�ب� St�[�:�K��(w��lHթ�}ݸ�^��^d|�K�#�O_��~��^�*�]bf93�� O[�L���'�L����:a��Cqu���L����H^ntOp�x��v�j��#���j�ι�j��ے�Nj��wr�˕��њWE��Z����߻sь���b�;�u�R�Nz�K&ọs�g�{�Ktz)�,y��lXAM1&���ڢ��7c�u�7f��:�>�t)H�f
>n����]�_,��yd��b=�EĪj'�^�]Whv�?]�%�v��f��x=j�`rDB�%��X�qžulW	��[��݊�N�m&; c�����J�Ҏ�b���t��k�-���H۹�;�э{�Uל��
$��u9�wkP�D�K�s��7��(�����CTg��~h|�M�=�3s6��X�~��&�V��%�U_^?T�����-�����h�b`9��K���J���.�KmP��v�a������{���%3I�KqQ�g��j�NfR�v��*imClv2�����y��Ǩ���ݼ�n����<=A21�g�5u����̌��>��Y��t���p���>�D�Aӹ�r�,����)o��n�RB+3ٕB�_9�2}��+�Ё֨ƾ��z9��h�����O�q�D�����D�5�b��tf]�"��\�$���N���g��o�)��F��n�'��ry�9�ߦ���j��v%�@3��4��P]Pߝ��k�Ȫ��^u��#?���P~���u��L?7�<z�E�~�4n��j�]�X���#&[Kj��=������/2�wxx�v ú���|Ǿ���g�5���-��>�Ȫ�ûƎH��<���my�G%-N	�>�'� 7���ئ�������w����W�~��W�n�
Qc쾟K�x�r�r��_n�ob�c��w�Q�g�!vl�s���.#�d��L��;��d�L���]=^ݽޮ�� �~j��N%����ޣN�D����{,^=[�o�Ф:��
z}�������ݘ؄�(�'$X�]hk'�]�����-ׯ�|9�v�?u��=4�e��5�cJ!׽�������b���|l#$	�X���ɮ�=��/!n�{�5\�����;r�%�\U��{�&�{�:�Z��TU�iky��=M�^�}��P�ld3�Ⱥ����;�7��d�Tɒ�:�z�t���/�Cg�Q���а4Q���\�]+S:�|�p�gIF�����V��1�	.2I.�Vn�'�Yݛ�ø\ńQ��~'AiX���Ď7���3�����[j-�����|n�i7B��ll��o�/kf�О�.~ĦM�
��,!�^c�m���Ap��x*�r��LC�r�7��>��o�)�%(�ר�\MoD�}����"Lf�ԃ�z�.=r-o�R8�{�[]�yo�e�C������,�B���T�n��mF�Ք�� L`"��}��6���I$N�-7�SNZ��J34r�#��B���A�b�1�_��,C�W�S��D�/�Ocb�mfc����⯩mΎvV�����Y�i���b����y��i��0���ƢC�v��ɫQm������7h��yVZ�D
�6!��Pk�{JܛR���{C��}:����
V����:�k�]�:��l�uҟR�y�y#��z�z�^�Z���K�Z���u-�\�:�'�8����k]�ۯBb��]�9p��\��M�n��3���mGlԝk/���R�[���Tf)�3�C{���>���G�9�FoUeѫ��Rh����{J���ji���u��ޜZ���Nuѭ�'m�����Ln��f>��o�m,M��+5��sF�g
HY���T�[��Q;&���oR}�ɓwc�7r������'ڼZ�Դ�P��^��<�8p=-j�F:�|+M⻊IX ��EcO&ʧu5A��%]�em@�P�"���*͋�}ZM��]$őd��r4��so�jgK�HM�=�6C�fY��� ��x��fC��I��Z�����.�Y5��Ӕ0��R���Eu7y*f����Z.q0�9�P{���f��\��FC��e��!�WeX��zbƇr���� V��X�뮛w%�wp<ܶ�;��:Kl�[��6����VWj]�.�`�yO;���_.����r}���v�9���Al�y�ܳ�����_}����P��ek�&����M���'{uy��{}ބW֨�^y$+��.�TUU��¾Ɲ�:�Q�1}p4�Wܣc�Ş�W���{�����d���1")mk��4�T8�x��T��8�y�t�@�n�y�+οbu��7u�<�C�ѩ�uy:X>��̯�9�� w�=��̋j�-wܹϧ�oH�׫���u�'k��K��;�ޘ��5����Axw��MɅH��F�m������>�L�=cz*q|kș���)��l��6W���_���-��Kɤ�����S���6���3���.�zeP�W_EOw|�l�ʶ��tL�~W�����g�C8"a{��{�a_QjϽ-r�<B�;߾x�q�h��)u!�3��� �Qa�J���f��qx]���2d��;��^m�tx�o)�uX�O�^��슬Y5g'ݟdچ��&�<���y������	����A_}K���v���f��,������p\:kn��G��W��E�L�a�{B�y�<X����W��g(]���+���S5�'$�]YP �0]���4fd{a-��8�):Aݺ����0�٢{��i��b̌mk����f�EԔ�Rӏ�(�+���y �}��S��v[��3w��.J�J�7�'?_��	S愡��b�L犂�s�������V�٬6'���lq$����4&}�С�(�W�2�I�ë�f����w��T��X����ݒ��z}0�u��d}]���~qJQ=���%$QE �%M0���t�#`H��������T-��	�U�8����F5w��ؤ�����Ӏ����~m�<W��bzka�el�q�ym���z�e9\���u�ԫ��|�~��*��L+�d������ܸ��s�s���@��d�C�޹�,��+s�xR���.^�u�ɍ�������jь�,��r�uV���|�]'��r�nE��k��w⪆��V�1y�4x��3_��5�G������WS{�U�����8�7�^1|�+v~����*\��b�W���N���-~K���}_gA��U��)���̜o�v��w!=��f����G3R�����D�C��=�&#�2��
��Л����}F&R���ޚɘ3y�V�op5�>�ʠ����KӼچ^l����u��V���5���A ĵ�bʡ�����Β	��j`[��f�<�V3hWV�ݣ��6-7������4�1�: E]���T��Z�i�o�ߢo[������8�.,�"�%���l�"��U�6�r[�ӕj@��us+�PMAgn�蠨���Ę��،͛B�(�U�O\��'����ʝL�~�.|���4Ӊ�ي\G+�w
���hh�����˧�����R+�~(�*!m�MM �t#0b����g}oO���l,�}�rb�2�)�ѾoiX1�V����W-{r�@�~FN-������e�����ݫm�U��`��f$ȑ�7��τ^t����Ϊ2Xэ0���S'hs�ۦ.7Ũ���������ƭ��:�=���8m�W}�1�ʦ������6�����H%�ћ�&��u�i�v*=s.��3�;;�MG�]��Nq�ou��F;�fS����O�w�ѫ�U~�Ι)��	���վ� �K���f�E0�]��{جg���/(�[B�<����/���M�]�::2���*���A����u��U5B���F
�y�_��~Y~���P�ώ?p���0�rꇭ?k��I�M���{>C4���*�h5s�o�OgZ�*��_0ؼ'A�l2�2��	jVH(ɒ.4ɐ5�{h.�PY�	��y�$P}V�m�N�d"����VD��\$Q��B��o7j�y����
�Edt{f������H��g�zg�̸��7y���*����׮"z�ՙ�i�Nߌ����7-N���e�����:w���7h!�2�7�&r�=u������S��R�A��;�wX��2��-Io]Ǵ��jŴ�q���]��W
��W:7.�*P�j�☉3*��ֵ�E���D��*�����Q�{=�#����fߏr���ǳ�����^�j��ٍ�͋	@�'+�c��}�J梉Y����YDz"N%�.�/v)Ы{�}~}�m �z�#1tsN�����Zc�Q`���`g$��RlS�����=��;���Wv�|wǼ:�ݹ�׷����3<��4${3j��i=�M�����{y���^&��z�L������1�����6~��~��m,���G�g���'�z�s[�{�\��gѕ�ry&7��#��/u��|���o;�u���^�?0Ev��|db�a K��Q�R��~IՅt����X�nW~��^Z&����^Yi'�{�ȇ����]ͺᙧ%�	�U����-la;��{�Kc{q�*�l� �*�q�۫��C����)�v��L�f�9����e�j�K��'��
�U��v{7��)��Ѳ�词��n|�q���O�{5c.^0jEC���$������[�+�$�뽊Emw��_�w��).�#����`V>YJ!g{�(��6��99��bB�<�D�9���4�њ��L���x���5�F���u]Z�]RuY�`��wS6��[b����R���)�p��<r�MW�MdBY�������u���'����U�:����-߽��M���R���6�����pד�Ԡ]:���l48�u��޹_	��<'SST����}�k�&z��c��6�.+�ǹ�T�7��>����z��m�B��N����윔v2��%�91��<b�c��yqS���g�F:������Õ�Is�����-ݽ���;�?\:5�V��z5���!/0>�$Z5r݂&'AnIB$Qh
Ih�HO�!�ş}@e��ڎ�IϨ%�2=��Cf�|�W�%&\N�\����W��"*9��}y�$=H]�`3�ћ�i���R{�uֱ�Aon����qyW���s�y3SYY��k��G��z''�^�۵+�z��{�Ε�ǹ^�z��"T�[֕���{��Gt��=�=�h ���s�Փ�6�]V�s쾊�R#�[:MY������jye��'9Y�{����oP��囦)��:>�y5��Q���UZ��Ix'���㛫*�u��]���ޟ{��]�K�,�
��Ewˇ\�쿇#2�u~����z����ڔ���~
]�=t��i�+R��M,��g�T��*,�u�Rv6�F�[M�wr�����u����u�}���劲�jſ{l,є���vu� ��o�䋫3�U��_�������~O�q�a�W�Nb}���D�kQ�^��_��]8:��䫐����A�K����%���O
�����;�CN����K����{>Z��|�a�
�.�ԧ	c�̪�z����8BZ�QV�TY	!-NF�'���N|��:��W��*��۪ΥҪ62��r�2�j�3}σ��.l��՘�K򬺽(��8���	q���)@���s�%'`_����������=z4�Us�$���[��ߎ��Ր�<Т�튗��o��ŷ�s����<y��}4�����s=g?Y��cΒ*c���������X����n��@ɬ�9몸�b[^�����������0���mP��ú(��UE�i术<��b���Vc�����Vv�3�w[Y���E~��m~����� V_�F�^V���G+�(�L{?}���7ۇ���U;�{[�2�{��>�����Bd�j�o}�Y��]�	��c�7~ĎP�w�n��ڨ~=73-ݛ۹���9��|28� �}	-��ށ[y�S��a���M�Qx(��^C�L�k�ûC�zn6ng�9,;��9��c�����pd�+��C����´>Y � ����}%�ճG�8�Dx.�`C�5]����gqA�m�PkpH�HHR1C�)m E�b��m+��	L�B�
���Co0L>��F�2��du���>[æ��d_\��N?$	�Eu�zhi�B�O$�u��F;[j���\�STP�mW|t�ON�.؟T,�GO�_nڻ@����#ҞP:����oJk.�z��`�\Xg��f�!�H 	�d����N�G]+O��*	)�L�'5�"�A�O��n�ks<�]����Mmnw[� ����L���~���dw�y�j��R����GG���UR���4�e'��v��az|��T���+��:7�,ܧo��wr��񬿱�[@J��+/�׵���Ո�������r���>ؘ��[Q�n�L��uigT�u~������!�iA��ݕ��[��姾�Chߣ�{B��y�3[ ґ��j��>\����q�/o%�h��/9i��y�����cj2!�k�m���)}����Uo1ғ�֭OL��$�T�$t.�R�iM��u��Q���^�>��u�&A�c���C���9������r�S�~�W�q=�+��ئmb���:�� ��~����4��9Gm�(�7-�h��]�)�Q�2`�7k�`�nFu��]�r<�~D:�9�w1Rl�5'l����J�r��J��^*�pc��7�L�8��^��c�x�}'���C=��%V��2w����B��Om[�y�i�����Qj��M_N]�94��[-����:����yX���/0����{������q����M�ⵊq"r���S�X����-�nV��F��$�¦S��Z��:�F�5z}��c�(�zn�J<���帽F�vw��v)�UJ󟻽��Z���������3v�u��L�VG�,��s�Jt��u��Yp���y	]~3~!*���ڮ:v�鞫�@o��l��/8ML^!�~�*S&vw7��px\�f�]�o<���%k�1�Z���M��$p��j\�6}3��Љ�Tm���e�{s]���z�9��R�rS��~�/5}�3+}Gr�V)s�h�\>wd�a���=ʂ�Wf�w��G�N�\kw�_�t�ԋ��ʌ�u9��ǺO|���m����M��QF������\��� ������(R|Q#L�{�X�ߟJ]���[��R�E�7
���y�k�/Gع�R��<vRv����Kzt��l����v����[|�H��"v���9I�����Ê/��h���Ý*+uj�i�[+��m���E���0'�j|��e1���H�e*�ږ��#�o.=$�g�2��\R8��_,�� ��b�����:a0;�{=�>`c7�����
k\��9�5�uN��V�m��ɭaG�.&9G�7�j�q�E�@ж/o+o���Wo;��克ќk[ؑ��>��6~C�}�W% q���9�H�cv������5�O\_Fg�#�������g���{/>�䂋�r�F�ψ#r��H�fu������ˢb��>�}���+2�}�E�S�Ҥ���,��^�у��}�4��2vzz>:T�"g��s&9���Vn;����>����d����G��X����� �B�:���O㾞o�F�Y$��L�^t[�|�k;�^>���̑}�P��ھqsf	�ج~�Q4xG�$I'&i��z�S~u�1
(���D�����Z����{���Eh����{3(è�Ն�sj"�/��"t.�{��9~����m3�2Rl�VG�CX)]х���lߜ�H���Û�O77�菎�������DfJ��b�+���cnw�1zdE4|��v���V�9Yx��b�^��n,�$��;�n�58Uv*eqWs�j���P��`A}�I��=�Q�^,��c`�74�7R�S�?��x�mX�,����^q{�a�|���`��r��{�C�j����i���/2��p��[1;�V�b9.�b"�𫳚��ݥ+�\�
���qХW�1�t覾5�����:̩�s���֝Պ�cy�r݅�d�B��gwD93O��s���K�S��Gl�=w���2��GK��Q��l��Jo��C|�p�,��0��
I��vZ�ڋ����zz=�G�$�e�-k[AnZ�ټ���}���X�y��Q�}qLM�UӬ����gj�t�.�!����L��Y?�{���Ia����%4���"��L4��5���$�%�?���_}�w��mf.�u������CE��g�U��t	��_���g�WI�{�W>Eg&����.e/-dӫ���o&��q�|� `��R=�]]L1���t�	���zo���{)���ܞ�.�D�V{in.,��f����1����e�g�v�ڥ�"L2��B�͸�:����3G���s�8���O>�)nL3�H���;ϥʴ�f3�~괉��W>����Q2Ǵ��fIH��s���Wx=�58�5���>fvt9sWu\P�W��l����ʽ����	�g�<���U����+;�}w����O�]�WnhݱϾ	z�Nz"�i���^�c�������HE#s�����Y� ��^_��O/ַ}�%m�O�-��bMG���Pc�5R���l)�C�I.�E�, �b��O�p�R����bu�w���0qq
���{��W�GX#���K�X�+��oB��)��`��RL ��E+��a��)��Ы%��Y�.�+���S#�x5��.�3�n�֏����j�G���Ǜ͎�rF���ŀH�*����P�le�c�Qnu���R�}}S�X8��$���e4�����ӏ�?�7����Xd�n�K��%�;e�����Ǫy1p���,�/��Η�,a�J�ę�*��LX�����de�c0;e ]ʸ9��]��L����[��Z4-��X�eTj�Dj��Ol�/�{"���J���S���4�f�J�keƥ_I��甙�0���4��A8GF��嵺*�F�>{���նic5�f�]�(JЌ�K�2�uh|�^p�'p����팧�r*��rw{jn��>2��7���S���V�[I#�`�*C�ۤ�,igv9�k��L�&d����lݛ㭌ax�FP;u� ƒ���
��ju�]�n��.�x��!G�ZW����J�g��+��=��&kN���m���� =!���5��/��1U���y׀�C�J���F��D�ef�(��֎���C�C)�n"����!O��eQ�ڹ뾛ܵ�LE+�.�De�����B�J3���i��;Mm�<{1l�;�,u�'	��P�?%V��;�aŽ�Q��n�d�Ծ��&	�#9�F���w�AG�Ǐ�yz���7[؂�%�X�����,��j���966�s�s0�Ę�`
I�m��A&���S*pu�d(JӖ�m��X[mtR�܅��V�,C���9�I�p�E*g�'ҹiQ��<۳y*l�7)\V�*y�E����F���:�x�޹�oS�0S�F��t��*��Tw�ݤ%�.��W��끂���V1��&�j��.������xv�G��R���Rr�O=�y�4�s���'`	� r��1Hg밼��kr�z��-#��e0���ɳ����V�#\��)o��K�Eb�z1a��ed�m�t��W24�h�'�[�7�.��v���p4�e̤r��~�m����M���'n��vK�X���E��Lj�زF)������e��h�  �%���M$'7M]�ՠP�T9��[i�B�p�|��5=g����yq'F�Ј��EU��y���+�X�����E%n�[j���o��s�[1ִ�q@K�Ep]���XL��������'O���c�I�e��Imt�}���������·~s�2��]�s��uLx�8q��ɮh8��]Y��*�,�����Wt\9��R[�E3�t�:�q�5Tr�ns�M3�>��r'Ƙ�K��;T�gQ�:��-�s�#/��'=�L(6����
��TE-�_k���-	d��"���S�|�5N��އD�]Bs�D���U���uG`��̽p+bqYtBnm�78�S�x�*d����;�=|��]Ul�m�_�o���7'l�ƁX�f�ڊ��W&1jՌ�����L�>�Q��([=��l:.~),�Nk���HZ-��-2ŵY6V�V��)Y��7Ht1�tuj*FI�LQ�m٤#����nY�?2�����+�d@S)B������#v5�d���-�n��r6q��D����#$��WzF���+M�n��[X)%�7pe�ʺ�:Ap�0b�ܰ'x�����<�0�BA5#��ݍ�*'b
�#�]��^��+�x���}�]d`Q�ĸRDm�L���謰U��}8��
�a5������4�o΋���|��"wT݃�N�e�,����۟E:߅�Oev��)���D�by�2�QQ*4l<v�e�mn�,�t�����1�"�>�'b��G�T�!�C���N3<w�����}�w�7�]_*Ni�:���ҟۨ{�5��Ea{��9��;�z}|�a���2Ԙ��e�R�Ԁ�����=h_|T�1-�׏�l5	����^X��d�5=ú,=>:�d듕9+*��/��n�+ǽ�g:��Y;�������܊�-!14��U�,�^�n{=��L�k��L���.�0�C�r���h�;�⛜!u�V�wy�P�Э�z�60�[|��S�&`�F�{Ks�t�-o	��n\�wޒ�]]vW��z������J�����=�_ٙ�湜�%P~3�~��|�2u�e��������<�e+U�4�g1�=�����wg�wҌ�_	���4-��{��X�:izR�C��~NלvU�]���UU����1��уz�����Ilr,\�UӐ��5Z�(j�E�ChQD�h?�;��j��K�5�)���#�N-��#/�ЏNF��vr�X}ԟ�u����iC�D�wS��N�� ��<ex�����.�M��s2]�y����Nr��ۼ�����:6�XZW}Xn녓��	��YW�[����J��MЭs}Liڷ)v-*��x�mY��C8q�p�d�٤I��\�����a�ۺ�4r�W@�r��<ʙ�;,�òm���C����墥̏Q���Y,���e��Y�ݙ�xJ�=uם��E�[fW�a��4���y_%s.!�W�*�����]{t��D>^�k��)�,�5��q<��#<�|���5�o����﮷�.��}H�O�dwSn�:�������%����4��%Vx�1�c:Ϧڊ]ꨟ����!�[���7Cc���Ond/vT�{�]�^��)�^K$�l��+݄;�G;�'��l��S�>=��E�гo 9�So����/�H��[յ5{@����:��!Vw�h&�6��%��b��Be�QH2�}�5�x��\���~]O�GmU�|� ��_oCf}L'�W[����m���ݯ4���Ѡ*�K�Gx&�bC�[6���`�D�<�O�UڵT�g ��w؞�O��52�f�3�?f>^m�
k���=CִA��ň��3�N�*f�2��5���ם;�/V��omL �������NU{�ۉS�G7�7~�e���P��q�Zy\�n���*�[K��f_VT�L�~�]|X�(��VT��
8�:+6v*8�k�pu��O%�E�ڈ4����YI���#V8�>������oV>�e>����=�%=S�I�������0p*�q֧��Ծ���J� x�8��=����qv��.`<뻽�����r�`�[��.�o�UJؽ5��Tf�ɝ���FN�V&͈\D��o_���U�!���
H*#!Ϲ�vm��.�vI���T,���Ʌ1�j��Nˋ6q|uʙ𓆉�On�纶U�ŖR�Nn�/]��;F�A����Ѯr��tuE,�7dL�U�3���9�6yFv@ګ�����۸��,p�r�=�?v��Qu
r&)S�p߯Z�b���-��5^
���OS���̓�ef
�,���>�e������_r��EZO7���wf��:�Mָ�/'vm�͉�����,��z��)S��_$W��,"���Y�q����AH~1�P�����i�1�$Ga�ڭҖ;���mz�2�'"�^l�:7:}Y�ni�e)���U�u(�lz�O���.p��K���d�o�#��ט��Gm]���������Z�]L�C?sϠ��f�ה��%�(QWZ���_@9Qu��w�>*�d�_wh�"��o5nCg:��ڛ|B
�^).��i�0wr��u
E�;�JK3��Rw��IS�7�C0���f�ۋ��iْ�{f�Bo��;���u<�l�)V��+wk��c��J�k�A؛�;��$/Lfd��&�����u��p��P�in�5雅��W����]���Q�?]D�q���- {FӘ����W׹7�����U�SK��A[�ǔ5^��g)�I��JDA����Κ�-#߾������S³"�8�S}���:�t��Z����3#��ןy��9�n,����ii��j&1���bf�/Mx��|��49zv�����i8��l�fu�"����^3���w��HS۵�P���n��̋���a����"��y�q�W�R�ρ��v<��7sv9�u���f��ޝ�)�.��}0/\g��î��
���ռ��y��(>�ӏ�V��϶=��F��,+ʶ{��8�gt��u�^N�k�u�$�j�+s3V^��ӯUc���b���뇝~���\=����a����9�����u�[�i�NS|�ߔ]m��b��R��z#5� ��\2��x��7٣���F��h�e%׻�W��\�k}�u�ǰ���5�!�܁٤O���:��q�G��o��qo���ut�Nt�(s-1�L�*T���]�J��&�B!�C.���N�5����u����W[ֱ�����Ko���7�|���"tu����j���SA�#l��Dw�ه7xa'n�D�<�۩�Mݎ����!Pd�eBD
�b�m(-���jXD#-��(�h���&@�.9���m���~*��F$8�h98��%DJ�ƝRٳ�Э� z5P�?%�o����v�/�,�/�w��mQ�C,��9mm�v��efR����>�y���]��3��w�K7�UOu߲�*^η����\)�};����8��'���j,f�Y8��7ʞ�r5�&�hQ���v_wz�3}���G������s1ݽ�3�̜�>�rq��k ���,��>���ͪ{��X������<��a�{k��±i��pV.3`I�^�=UژX�U�s����[�T3�xWv��z�{�~�?fE�4z����Y�	���|�5{��;�}��x�>�1�S�x���y>���o�%o&]T?vߓ�x��{�.�3^:U��s�iĲ#�0ʟm��Ok��0x��ʮ�"x]nd[�|p�&a�I˩��L�]U�^[��%����%�j��5B�rʊ�3�4s��ϔLhUy��d�>q6.��J�mY!�c%�nQ�iK*��}����2�d{(�R�c3]@�!a�d^�|������ݍA��~�3��Sy�`~��\N&1��֟g^�5�
 ���n��b{Ӟ���װK�	�tn�|�Rح�'�^Q�7���·Jv6�ڔr�)R��6XW'W�^����z�ܘ����'�����1�o#&�LS.Ǥ�L,�Wҡ�9A�WߺV�}*2nz��8���r�_	����N^���p��>��|����31���Bڼ�,�~���<�Mjm�t�/[y�/���>��z�u�}YV}�$�T��eq���4v9�1�y��ʠ���]����u�<Z�B�fz����6Ѿ��̓"3��ܗ�b�8�0O��
���I���~���}GJ�u�Չwj�=�nJ�c/��ْ	�v�O����>��Q�x�����?��p���{����j����!�|��Jnq^*�{�do�V��2Z"������^���ꀻ��
�8l'X�O�^�8��qD��������V�W��,H�p�+��ʗ,6N��2��W��r�w��2�W�?v�u�����\}��n"Tl���6�Y3X3$�`�M�{C��13��U�g8���y��>����6T^��\t�d��]�8�W���g��^���7;�iۦ�D��[�F}�ٝj��oN*j�NU��^ٮ/(��p5��A��f����;ڕ�E��CC��E��^"�SᥭY�xp�Q��n^�˺ӭŜ0��rt�K+kD2�ƸknGՌ�Ρ�^�kb���6f����f�����l��:��H��}��OMqYg�����t���I��_b�׏bD�3��2���[��F���j}���:�U�D����϶�[��|��x��2��B�fC��K}o"�C������s��N�2
ٟtfN��1�7J������l:�Uk�}F��"͑Z+�3�5�ӹϫ�e+r��W���v8��&�=N�cɼ��]ݵ�*�1�.����ځ�� 7"�����g'\�5��Rڅ#��v��cT��G\�gg=]4c׏H�.x�I�Q8�8�u�w��!�R'��Eؽ)����_V�qo�u��g�J��ޭ~�7��DB��r��&�if�u]}����/����ȯ�I�k���]�ʽ��ߟ[�tn��I8�Ϯ�>��/�ߗI͵���G;���0��_0�ߟ�n7іf{������r�uZ�+�5�����=�J��;̾ͨnS��Ҳ��V+��P���<F�/= �6��K�q5Zs:��7QU��,���l`��{iǳ��������B������B�ȹ'��rw�v��B����BewY�+9Ŏ�o&C�t't�-��uu᫦!e�5���r��\�¬�ˆ��<���"s��S�8��<�Zl#��mAZ���	�+3����{e���.3ӧWa��1��.�Lr��^��.τ� �/�W\=��2l,Í��Mt��ˋڦTf�D�ۏm�Zߩ�I'� �Q�*MO��}5��u��v��t�U���k�p�.okش��%�!��5m�)%r���Nخ�����]�{y����j�Q���t�~/������>�N������
�*˫��ڇ��|ʑyꅃ՝X�q���1�$��ȏfW��(���/�e%�V=�~2�2���!�G��0�}p�t��t���]w���]��.m,�sww�~*}��z
�<s����3F�z���KT�z0�7�]��	���nQ���WG�����ٗ�jJ=���jw+���[c��ø՞ݧګwa�>���rP�gܫ�>�B���ڊ�?��T�s_%s~&{��/gv�9Z��@B�����[r���nsI���7S%Z��Ǐ���aV_��~�1**�i��j��Ûތ�q�K&J�6�E�ߴw3ة�TW$I�a�<ƭ�ݛ�i����S!���9��D�5��&t�T����M�i]�#.�vy���@��;�B�Č��b��v�&��C�{�[-<��$N��f���d��wnw�a��,��j�Q�����M�{���M�MjE$X�º�Ln�2�Qt�f��74{���$L�,Cz��uw]wN��D���@єrѕ�Ɗ7��jk�OK�x�d�lW�w�����zf�B<��#W�Z��6&����*�,t��E�_aDo����S�G\����,���C�N��P���{,�6]t���d:�"��N٫��+S��g���)Iߜw�gMB~�3B�uS���Pw�|wN��}u鸻�0���#�&��j~�Տ�(v2�wU�vʽ���dO����;�:*������C�U�q���`Q��zǄ<j��,H�I]��:�}�v��mzz��]�G�>�p�[f��h���eahopd&�䵙�(
ޝ�0�q5-am�t�֝5>���0������%r_}���R;z���8����Q��J��W�A���h�?�ͭ}v�5���i�뭘���|=�c.�:U�~^ꔨe+�A��ж�L����/	%]�y%�}����R���w�r���ٝ�GB���ﲓ�/�!���5��Ha,�unj����X䨤���P�Mr����)��ߓ��^�u�Y�d�~��t.S��ħvy����Yj�A�[�?
��ݴS�����a�Ep#�zt65{-5�����X-J��x�p��ס;fA2��k{�:I��Կ�2W�KxI�����y���9���;Hz|�C�ڒ�iZE�^���������m��i�%�u'w�wZ<����u!�7yڕw�-i��}�9,�Շ�]��H�H^1ٰ��]�b�9H���2Zr�4a� v���k�Qimi��l�42�+����x,͊�c�3��寭ʦ�Cw��_Ntg��9�f�\tWm ߪ�b�|�t����w���rU�b�ػDIH��%9O �;���^��eשm����\�ܭg��G-�g)��/�9=��7���֚.n�_y9���#C��6�ܭ�E%���fW����X����G������v���J�ݵ�v��ת�O���E�ċ���n�w�`{{��<v ����kY؁��郞��M�J�xno�u�;(�E:s~ݿv�m�z���G2�#�(���[���u��Vn�EfvU���n�ߢfM�IH���]�Y����!��qV�QJ��a�x}�8�����ۄ�b��)���ۆeƾ���ӓ
�m��z�!E���ef]^���fp�pt�[�j��B:'�!�diCo/��C�&\o�ρ����\/���Q0�GȬ[~����f�Pw�V-�k]�z���p���|�Lg�εz]=��j�_T@-^&�u���q�潫'ޯe�O��'Ju��k�F��YP[0`K����4p���j_L8����U�|5r;a7�E.��r'��kk8-�g����cf���	�F]-��擂�L1R{�\��Ϗr���پ�)��ͧDl���h��\�ܓemB���j�̬6sW&J!�+{w2;����P3M���n��y�]�u�8����ѭ�tk�uÕB*w�W=y���d8�r���Vն��\�m5���1@�ٷܲ�P9��X���r�V�%�;ۚu+9�Qn�*t��Y� ��"y���fKzΐj�pY��z&.N�j�}űtb�cr3&z���W��z:{�w�����Օ}��r���&'1ߵ��N���X��L��pqw-���<��N���pbh�\�d1�2��1Ge2D;��3���,I�X����!��u�l� 2�_��S`ι��e��t�"����m���G(L��@}��:�u����(;?wml��̹���b���u���;�wJv=]'.Ѡ&�s9º^u�%^�zS���k���Hr�0�ѤƦ2o%~E��f�;I�Udɮ��a��8�H%�}�4�t�Wj��a�s�;EdѪi(P���AŮ�<����oJ5�h#�����7X�Mmv顏�ve�� �}��7T #�<��2��"W%,�39.��M�O�E.C����P5��6K�	Ro�t�\,���l�w��%v�`���[�����\O@c$�4�,��QNyf�[��d*�x��R�!��&��fI}��(p#m)����nc�N)�3"[��N��N�F��6�F�Ӝ�"Jk�<���E��Cw'��S�1IP;f���X���]h4�N�;��D����==����4�!�s$R���k �Wl�]ҕ��A��)g�##-�r��KsFu.o�"ኖ��]	��֪knf1y�F��ɑ�{0�l��0�J�˙�
0�t:w����ѕ�bY]kX��Lc�aU�j� �R��mǱ�8/t�r܀�V�cIɬx�Y,�u.UlB�bb�d)T���05�V�Ƭ#7fӭ�e��=�x���/�'s�^�mWR;�/F��W4$���P��Ma����u�t`��9��ER��3�L"�mX&sՙۅ��Es�ɦАY�P]�7�y��wH�4�q�(mhAe�;����������k"ޛP"����q�2c?��|N�ҽ��}]vDu�?\N�:�<0?L�Fy�&}Ď��y�w:6y�-�ŷ:��2QLqR|������ߐ�c�$�]�.� ��Ǜ1>�	2�fLξ�j�*�gzs�s1"H���8�c5���nef?-W~��ꑆ�������TF���)����e����M�{�3T��Ӓ��9���5*��+�2=$�6[�\�RI�m���mV�o�AF�|W��e%�l�����z��K^�xWN��o+~��8�����z"�Q��6�YY�l���c�wzc��A��=s�~��V��ʙ(�H/g��w�����m�
�L﫝en��Sy3�˪������"T���TL��:�o2�='=���9W,B�2���ܦ���'���Ѿ� �=���U��طH�T.����'��m�zr}�a&�1�w��)�"��;'b�?����%PҞ��oE����2K��3y����>ռ��T7�"}#���ڣ��DWݵ��X^�:��>�Mn/.�����|�΀�Q��=ޡ0��0�pJh�t��˸�j�z"��c�K̇�۬pq�u16���L���]���hց3�0+�KN��ۡ��:M����;�`83����+sY�myT��/˶,lH�L�"���ˋ���U��KK��I���in��7��!Lz�,�uw�s�m�E��.�g���w'䈾�����>�A������|k8k�M�z��lM8�m6%*_%N�|�m��}���������d�����%sbꯩ�]46���	�w��:�2���kA��&��ۯn��zxS�ҳ��aS���ߥ�tD(��(9`ڮ��Ro_xOb���ꊎgK��JU����t�Fb�	T��m��Ut��z=ZS6w�kb��l���G��&��q}.��uM߇�т$�U�v"N�aAvx�lXY3�Ue2zs����d����Oy��o�r�Tk^��n�\���/+1�Z�e@�;��W��c`_���H��[{����loa��ut���jú{J:���JI�j�#�����)��b�+�[�y�n�X.�ԅ�5<�x�1 M]����*W$�k�o꯻3jp��v�)�Y��:�&'��M����u/^�6��Y}��w����}{ �F�o1nL�&$ɗ�J�;��5X��'Nh8(	�A�.�(�����֖,��u����L��.͌�ͦ�d*l2�!BH*�2���봍��c��@��c�8!�`x~k��.T2Ir����ڃ�k;����B�g�Y�5�g��cE�Ȝ-������v�/Y,q�+U�i��eq� ��t �eDځ,����'���7r�v��k\G�љ����� ��`��*H�� ��Nr��}U���[�/C�\� w�qA22�&{ƺ�$8��<�K21V[���g
���gW~��5-Å�'Y����Qo��÷��4���(�)N:���(���~�����ϲ����V��=�6�}�����>���?��S�[��c8���4��)�h�]k���w�>t�>�j�W����=�NCo��[<i�[=���Y�nf���ږ���A�<<���2'
�������]?Ku}���myJU��u����S��o&�x{R�c=γ/=��9w�u����|qF9�|��]��,�n�ڧLpY�|>0bv�Y�^�T�wU[��n|��~�Q���i�������_*��:�J����s%۞�o3���'�͞�w�r�$�_b�-(�4BhBW�3�ݡT͒8�HZ*����S������x�o�ݣ1uc}q���&lG�ּ%���^S-ƞ�1���)9X�R~vys�tjǞwc�
�-�ޡ^r^cH=���:0n*`��¤R��C��U�B��A��î�t*�țOs�׽ɴ:j{���>4�9��|��S\z+�R�X�(W�qt����7��VS*ͽ��%t*�ejjF:��o4�	������c���9��9�w�ܣ��C�hNp���+������E�\��"�^?}W�=S	�����k����Jv}^��P��)"���e��}�.go��jͧ��9�������p��ݵ3~�;�Tږ�:��C�f�J%'�J�S���Z�(����mRW���zײ6�ޗ>��~+ϛ��*�>��uqy=u��͛�$���ڳ�r���\:}褀j�SX.b�����YګĐ�wY��m���l�M��k:�by��;=���+�7�5N�y��,�U��%�T�%�)�N�~h����O�3:k��i�C�B�υ���#��xv��ф�yJߨL�^�����	�ެ�+����b�TQ�s$L�"c|����j������nut�R����[�y�,��z�yWS�d1L���e�ߡ�V`�{V�RC��{�y���c�z7���e�|�q��BWnX�΍'D���>ϓ���}�i��3�������\���@��g~
�Ҥ[�i��<��c�Vq��U��]���B���BN�Xmh�E7�$�+*�:�v��+��X�fs�hD$�uz�]z��. c�[�8�J\6�¯37�s�5ү[��W*��=cz=^��_o�|n �� w/qwM��o�wV�Qݖk21��ȇ����i�/pT�2 _nށ�o�Q{�p�e���&V:i�[�T�T�]��><Ԫ�H��'�����4���}�w��~>gȻ\�|�kk2��\��Mz�z�a�_�U��5�ħK�������Wެ�cao�`�"��aHх�܍H�
��*I�$��}K����E^��FM�	�}s���_o���3���dvyή\))�R{/u�mM���7>�9=c�Zx��У�?Lf�t���ySǶy�_����Tؚy/77U�"Z�ݛ@ʶ���xSsz2wv<_PX�U�g�	2㧼�vf�m��\�m��u\@>b|r�D�;٧c&c�k,��)�{n{���s�����mc͍�N~_e��pǸ�O9>��|�B��rSW�9���o�h'й��D�uc�8)�Ѫ��y����s��ׄ�F|'ِק�y����������/�
%�!�v������'M�ד,<��;Y�y�b;�u8�A���v*�f�:�N�Ӕ�둧�r�_[Kbs.���9��Q�
sF�&�ʊ��d��S�
��*G	!����z�ė�K�}{:�s3Nz{�h�3)�6;���c�R���dH��EQ��mtOc��L��Bݪ�C҄�>�٘R��[27'�L0�ƹ[����=������o��k��z���q�gn���}�<�wQt\!k?9N�`��6Z/�X�v�;��ud��yH����P;M��ʊ�?�ϳ�N�~��NͰ�;w_zV�d���z3E@��Hy5ݾ��mo�`�"����N��^m�&{�'��ǺK�s��MA���	*�"a'y�'�����z~��'v�U��~Ȭ������ʄ7�����_P��ϳ�k1%{�=Ϗ��D��tE�7Q����o�U~�v�*k׹��*f���|&k��5��O:Y���B/�lLW�;r�}D|���E�v�}X�;����U�cu�J�
��1~��H2fw��D�����{Y �W.�o3n�NN\���*��?a��T�aE����KΩ��t��U�j;TE�pJ�뻷��kf�F��g���:����gw8؈��w��;�oכ�B�d`ۺ�[���7�ҷ�P$�-ެ� ��y`<m�#��:�oO�r�M:'�o.��-��nZ)���A�ǂ����
(�J�I�) �U7M�q�-Wy	Z�x��Ff���7�{�{E��TUGX܅��qZ�j��_Y��o�wH'��-6���`.{V�id���b��8��k�Dne홀1�5��y��B�!%�����|�D����ѡ���偠Uk�a�a�ϝ�C�6��V0��}�gcnjO��
�rЏI[�4��a��+]��������[}ջ���DJ�y�u����j�ת=��z���"���UO�����S�7�5_^�
s:Zj��֋�^������z���s����@�=Z�{���1{�m��۶�Ie��5���j���t��H>4Ǖ
�\DQ��sM�����׸�'����y���~�YU��\T1�pwe�ї��x����6�k��4��F�_�+���b�O�I?)������m����5³�2������㝱1��.�~�Q�F�	��0�;.Z���V�]�����+�T��N��ꑎ��,�f����^<J��'��n��y絴���`���ef���v%z����0����1~�@���{@:�T<����	^�WÃO��T�*�G�U�W��H�J��d{��y���x�����H�}F�(�PW�{�.�ϒٸk����F)�A�Y[���>u�Z���v�*�r��Z�I
�mb�; 9{'�e)��OD��(�Q�L�b���)��F��Of�X�g�'.}B�#z�M�0�w��[�Ƹ���@�87�hL쭌^��*)��/î݋�C&�]Ӳud�Zb���!�hz�ja�f�!��sQE�}y#U����wp��yg�佘܀j~o���>�I>��=ή8�No��tO���I=3}����]y�aJ��Q�N���:;n��[ZW9W��p�D�uI���F�%�<2̬����6%j�넧����<j]�����@����1~�b-��dߦLrѽ��:�Mvػkzb��v*�r���J>�ϙyq2��6u7Ƹ�5Gb�L��8� I��/ڣ�Eg��,40;x�]W{b�\�4�H6]ea��m�9��%������tz�eE!!T��nvs6}OTO�ˍ.}gۅ�#L��-2z���ζ�>��ʈ�	t�h~)-~�����}�sX���v3�=9S��i�r�c���y���}�-�b ���|ea�Β�Q��\����b���u�|M��+�����;29^��e,�L�[X��2w'ۗX����W~r�J�P߫���D)���X��a��~��kP��r	�WW�=G�^�sE�$�.8o�7�.e6+�1,�O#�^�gF�n�D�\5�g �K�^�S�����4�3�r�0�uT%�)�J��+��9v������EǍ= (8u�^I�v�In�`ܠ/$�N����Oo��,�\N�S����q5r�M��n��iTҜL{�z����f��'����ŃU�U�n���mMB�N��]�r��r������nVt�IJ��=R����o7��._����{���t���W�N�+�~��3������d�uV6=yݞ��7W����&=;MQ��������s��>}���u&<fp���8�!z�7|\�O�bK��a|ͤ�~r�4��Z9[me�[�=������};�@^�a6ǋ�D�y��Б�_�l߰0X�������S����!�������԰Tlg�RJ�F>=�0�ÃF|!d{/ 2G�����bb�S@H�3��}�b-Ҩ�v�3mP��q�j|�벟w_�ֶ��������㞆�������5����(�G�O>���"M3y����c�xF�A�`���7r|X�ٰC켗�rC�?AҘ���4G{W}��>�o�Q5�8r�sv3�{y���.DoE}CNX�3��0s����� =��	��<pu?�WϠ�M_�l�����h�]u|�>/����df��pp�utW�	wO����vk��7�5����2�vz�g��G�x*���m֢�|D�9��3R��'-͏BT�W�[���J���K�ΛT����Z�μ�����
�Gv�)���+�\��I��`�*N��3���g�BP���\Fi���#��RN����X��g8ǉ��Q�VU�꾑E������^��{K�B�������e_<�2�<��ec�N���8�G�9�qo�q�Ҧb8]̈��}~>x����5���& ���V�����s�}��#J(9*�֣��yb�^�@J�����O���>��
O
Z�!Q������S��Dt��A�A��������E�� �<��rNbG�m�]y����ӷ�wg����k��Cݣ��<u.&���ެ�!K�� [��o�>�%Z`�[��*P^ߋ�X��437"�<?1�?����@)$�y./4���#��
�������oOTG<�}��9�`��γ��f�]N�������C� 7���󎱜g��Yί���ЊM����������b���袩�xUL����L�.{�1戞�A]�D^D^�O�<����[N�;k.�tݪ��=�������f��ry��ڻg�g/�^Q�P�{��lv׵�{J�G9}��FE�Fl����݊�P���֌"x\^���ع(�.��9h����#@��^�������f��n��&�+��9
���������Y�W�!��,b�џ�c�@��>ѳ���=��s�f��7���q�٬Z�ޔӟY�M�Z�{�VʽŔ�cJ���5|�7h�ù�h
wZ'K�rq4���y]�J���V�ݎ���0�8q�j�P�ޛRv[;ߟ�v��EGn˒���ʔ'ad��w��(�^Uw}�p��2�v����n��R;�!u�:\�5vζ���>�;V���[�����A��=�+U��X�^uu�k^i飪��c�=��%=�*W
�*���&�ܕ���I��Kϑ���O� /1���I�Fb���QY�|FU��-�3%복�6�u���B�t$�c��vg�[9�X���u���9����;]0wV����Q=֦��J�,�B�V�\.��p�c�!�WOr����l�h��j�HJ��`c�=[�ȣQ^֬��	��f,+�ܫ���ƞ �^��������̡���r���ip;�'U��Ch�N5�?-�̆Q�;��W��]�ݍ��oP�0�ߝ�YڽƐ�4q��]�(i[w(u>퇴rp��׼t�x�<� sC8����ˠ�[��7+���G�s̨o��iҩKf,�fX�y� +��j���B�vf�W8z�a�PM.��*H�gPx�����Hb��4�t.�$6�sz����h�i,c��뤅J���B���`��뷒�n��"����nG?=�|:���gn�`X�iR��9ʚ���D\ko\�֒����N�W�+�@:�����������1Kds˝}�L8�"�"�VV�Y]��Yۋ�k�j� �YЇ���c �J��x�/��s��s33/wv�H�4Y+��&э"�ݱB�������H���~���&�)-�,bY��b4�ՄQ�IF��)S��״�6؛η��m#A�u|j^h���[*~|OM�@ ��?�C(]1�,@6n�'���� �-��ĄaL��٫x@����;`w��o�1V��������<�W��ǯ/[����&��R���.�+��t�q��Ѿ�ej����m3�M��8�M��.n%�LZVP�dʵ��,��Ce��+)SHh��J���6l�"�P]s2��F95�2T��X��k��ڕ+�t���C�m�v�}�Փ�<�a����V��:H����c��ud�DI�ч�Ъ=f���pa��ʉ����p�9A؆�L o$(&ZRM�����є��M�PAY�{��I�u,�{5�4�E�T��$w�Lf��'�۱��e�wJ��)���a�	ڣ���S	����d�}�[���ξ�)�M ��&e�Bոڌ
Uht������.� �*���ˆ�\��R��|sT�HJ��'/9��C�8�#^�ݳ���$~��ˮ~��P�e�U�UWm��v���1�d��Ù��Q`��E�3N���N,�ԍ���*
�8�d2α�mؔ23�a���p�j�l��L�Z���5��}b��0�t�5A󧈈���E0���r ��i���s��)�h�"g^��⹴sT�~w��8����P��T�P��a�$���!�wAK!6I�{)���w B�?Үڲ2k򢠬M�rh������nF�\h!��D�� x���wb�I�Q��Cm<AiC�^9D�2��y��[d�����Ѱc��J�.pN:U���Q���>F~w�@�XR�!�(�Wa�_n�r���f����VWau|�@��a�x@L>8�b<{P�I��Mv8�K��rLԛ�sc����� I%Q���_�\%�$���ʑn�MkR�μy-~#V���\Џ @D�1*�'	D�Jۮ��d \y6�2ii�׍��L��8G�\��)�KH"�$D�Q�]j0���T��Kc+l����4�2"�zn鸦 ���vJX�{�:*�j�6��_U9��]���:�ኩZt����@�'>L҅.���5_�b�K�ca�Qg��pU�N�~�}��M�{b�G��,κ{���c4}�0�C^0������#�n�(�
�.���$�T�9��pr��c3W�{���@ޣ랢EI���P"6\x2=��'S+U���Xp���߆����W�����n���<>�Y�u�X(;�S�[����4��Dp�U�Dj��O���ٵ���g�5�����ڹ�̹��� {w%x��wE>���r!�g>5�x��,���/g���~�:�/�݇ǴFٻ�7�w�J�������q��@�]<:Fw� �@���	P���p�^���ë���v/W�_�݀6ᕈ�e�i$�!㢻h�yQ�ww���^:
'����U�#pb��a3sT�v`��Gp�n�\hx��_8��0z�
�"�+������	����B��٬i��p�UA�
}*�p���fIFz�ZGr�j}�)Ƈ˛�R�%�����|uR����C�
���2���y|�">Ր�ddK��#��O��{1�=?L<�!yV�+D��|<�>�מ��3_��C7?2��r'�Y5�b�4֝�ߑ}�
$���b��_:A���S8�i4���w;Cc:g- ���k6�N��F�&Y����*���w�B�t�V��Hf��O\�U�����뛓_g����zl|7'�TJ��m���B�C:n#۳^]4͙�6Q�����]��evER�6Wok���ga����]1�~^���z1�󱠇�I��Cx���"�TS�7y��O%�U)v�G����:��yq_��>��~��״�| ��b��j��Ԝ$�(���z�O�r���^�Y������k�M��ά�����eq�N�W�'������qGiB1�74w�i�Kݧ����q<�Ezdho��@�7Nb=�3��}_Jk�!(�&eU-����|@�<�wX�"H���8��? F�]}�Mn���1�^�茐!ď��H�ȟ%��8I�&Y�<��9*��_e�8&��%s�}#�ș<��v�j�囵(uտ�� �b�BQ��!oÞ����9��er��̛����kP!���*���C��t{����J�֠��Fr�g�c���ˊT�_qwy��=D(>^�Y��.��]�^U�̱�>Z/�1����=W*�Ϥ���c�f<S����0}0s�뙙A\N�}�O�&�[3t*���F�c�i���T��?O���ǪXg����,m�[�[�3iuf���z���w19f���ʽ	����wvT\�g�Xd��s6���i�h�֛X�ۈ��W &2��@Wт�u�"w"�1q�E�v5� _72�YoQ�Q���{>�?+t���g�'i�y�G�21؂�Q���v'�Yf#Tz�p�;Ǐ�3���Cy1���2���?`�j���%"T�FWa<��K:�\E����n������S�>���-�2��5P%� �ڜ���P���^�R8F�ٻ�m;Uk�?W���;ʡu�&3����&EH#�xt��@�G�)E->�߫I
?-��p5���K=l@��XS.3�!���bv8�b�Ұ��S>�?,C3N���jD#�|��is���}L8_Ń~����/�i���{�g�r�f�V�rAo�:�E�y&'��Q�uC^����S�nwo�B��"c|�}65r6Ǒ�v'׍]����/�7���7���9�5rb��sU6_Q>w1'pG��7��&iGz�p=S% ���FF�;{ӣ�7�}���AC�;2�$N��@�9L� �&/�1���2��@��w4~t}�fO��܍f����%-�����JC҄�����ʀ7�|�{_e� V�8*a�����F�A�}����@�מ����.K/;S0M��w>���3|d�P�#؜��w�V�c��W$8f}�ڍ��?��E�k����eL�lU����ݵa!w@B��c�۵}boM�sQ��Gڐ�����n�ѕ�q�s<�۫���I��r�J������:E톘�O�A�sd��b��zŞ���h���!�ў\ˡ2P1idM��,9[K�Y�P�m�c5XzaIN�nn�[Z�į\N��j��>\��_y؀x�AՌ׮DG��xs�pzO�Ʉ$QֹE@q9�ej�5�@�B���
��q�C�9(6_{�핟w����F�V��9�����H�d�_�=���)8�Y�@����"O��GU�v���)��>�n)iZ��hi��'��k�{�2gBBw=����~����%�e�'e����{�i'y�tA��/6}qf���ݴqXϨ�?-�/�%3�bU+O��T��4�>s����&M���#ѹ��g�����%'�?ŶQ�q�u|��.p������l>$Y� {z�0�D�Uh2;-����[Z�ϡ�=���MS3�a�MK����o`x_���>N��+(h%B�~�=�^���_K��ݞ���؉�ʻ�_`�bt��\o1F��\]��h��%���>���S8�U<y=�9�$G�� ���Ҽhl���s"b,8���N�	�p�< ׸/�쬅�v}��ْO���!��3�ϭQ?p�����;����j����N�;#-�j�zo�e���}�]CAu�-�ƺغ�Nr�Lgk�^�*�$D��Դ�,v�7\������*����`�".;�7����V�	e*��������ѿ��w#�uc\�w�(��e��f�X�D2������e3r�i	�u�Pu Y�`�x�M{��+�w0 $'�� #9;4����H�]�A��+L	׮���nPlJ.�6K?A7��ur����E�^\�r��m�%ܔ)�E*��,]�M��wʯņ�1WJ�K��|OO	���ʓ��u��gꌝ��!��ބ�2��RwA���כX'���������Uv^��W�d�i��O��?�~V���r�k*.���v���{�U.���w���}뤉̬{=t2;s�A�ǯǀ����4��å�\�LC����ﮚ�t�6��w�K��.ˬ{<�4/X�+�>4ْ�a�ǥ�Q~�0u|T�|&�����r�Z��>�sS�PyXԥ�_IY�};;�M��]���N�M��8?������pV��Q�@y��/k�p����2�_���}�I$�J]ou��WM�T{1#��$ϥǶ<mgc>���/�/?`ܤYe�lR	��,�n2�e��易�&�Fw��ڕ_�W�V�����4r
��NG_�_2�4�9ϲ�����+���k))Uuۻm��s�c(�ǸzLK���U��s�}+yl�h5�yzc��l^��)~
�d��|����`#��ǉ��+UP����ЅG�h�E Q�Q`�/��ó�.w�����m:흏Ρ�<��WΖ�KK�/��~��s6�Kt�A�{�a�+}����t}Q2��`��p}���+���`C�e�G�o+
���5[��v����cd���t��t4�\2��Gh�v�<y�����o��®�T�[Ŵ�H4�2���k�XR�.�+�����6[�E&��j�)��E�cJ�c����Y�=jXטx���n.�ʞ�W�˩x��J��P5�3�����%�I8C�R3�����q�G���מ�>�K�:�{X����&;�d�#�D���p1ş��w�`xצO�>�&��)���*=�i��CS����L�9� ����>��>―E�w���Lm}�ZC��T3~'i�����P�+�LX��R��΁�S�4��7^���|���� Y�b7�C�F�U�v�UU��a@�?Xo��Ԁ���
j�=ޚ���6
�Y�
Tmf�&ts]zâ�}��_:��y�A��\rz����]r��v9�����k�[�/ �^�z.2]|1(5�	�<���]��;n���z���� S�b=Qm"��@B�$�
�����&V�dYQ�ɶ�f���������YƧ��I0 ֯٦�꺘��{/b�����
�K�3.#վ�_�z1,r�G�Ɏ	�?Q�T�?}�}���ŋ�K�䛥Kؼ��M���.�v��~d^��-<n��ϧž�B�+�e�EF�v� N��g�͛��
���_5��G�mf�����TF�V�*W�Yv��>���L�&E�������p�š��1a�JwLs�knY���2�=��jP>Bo����Q�Fּx��}*�{Sq.�u�r���K5z�%
ǯR�{Ъ�C=×}�ް��%�gA��Y�/Ge�5)������Y�x<|n��U�Q2%�$3�����ꋻV��&aF#���}��)�T.�<̏T|$��K/A��F*�p;�&��[��E��P0��C�O/�<�E	�b��:���I������۞�&4I�>�(�I�����V�nɚ >���|����"�i�U���y������]�����;Sp�d(6�ϧ&f�S��1���4t��^�zu4g�e�(s{'��{F*ܠ�'�[9��xWV�y{6�?���|zcF���S���)�M8��>�Iɑ,Z�xA2b�0�m�AJ�RE2����������`���4;���b`����k[ZAco�hT��:�Ȋs����sT������T�����N�&��U��Y�|!ౚB�wG��좃.�.��.8>�}Z�L�GFz��x�i>8�f�a��a�q"'Y�1轙U^>{��)��O4�\�;k�	��:4E��R����{n���p�_����Ťל�B�C:�;��!\%M��~�*Ǣ�(�JO��k�p��褹^�f6���Dgi"BpK��Q�w9s�ߦDN��
�&��P�����Mf�h���Q��s�ur�
�|-<����׉$gա�+B]�z=~�/�iH߽�K�uc�)�T���|�o�#}�����z�?p����j*�,�t�a�qC�g5�1m�8��C/�=�0j��[�P�\f$�J|º쥺����qC���q�,����(�Rj������.��)M�]@������Ż��Q�ʖ�\QS�����N���ᅢ�ђ���v,ր{�e����? �پ*9�/����ƫ��L��.����ƴz�X��`o=�6�۠��|~E
m���9��b���_&��iY��P��X���Vo$�����	�'�J�YPQ�۱���mc���.�>�Y�����|>*�;K(U:��]��F%^B)�C�h�r,�V|=�%u��1^e�m��������a ����۾�NLz�`;)�6d��AH���o]����-�\܏�@JJ���G��'(N5�m畡^��LD�z��+ywq�{3�#��C�����?j���V����a����t�D�fb��J��7M}\tl��(V��q��P��J�r�wg��m����Ow
��g�mhV����P�"#�5���D띏 �0y.9�3����9��(upd��˪?�~���{�z�����qd!s�������ƀ���#�{zWŹ��.��Ʈ�=�3b�����hw8�c�T�>�>ȭkz2 ���Ԟuv~
4��8������~7��?R�<�����P�.�P�H�O�!>�Dm�nM�O����<��BV�{�|Y�Mz��d�]�R��"�y�-Tφ��ӏ]'k4w�ܸ'�%2.mZ���˂̠�Cot�EP#yk;ؔS�u�m��$�+�d�-���"rK�+����$à�rם���iݗ��Vh�F�.�ۼQ��9x��H���Q����2>H"2Q�F�b#4���΃������[�!d�vb:ݍB�!�����fh�t��!P�
�9��3�fcN�>��ǟmJZ�5��T��GL�����-p���S�Z�|̍���@��)Fe��J=�s���gHb�H	�����o�ف��n3�=q�^Ⱦ��נhf�$so7g��)���-Բem�j���U9F��^7"�W�v�G�\��ED�չ���]*����x
�r~/�kճo�g���+$�~ov�օ?����}�A緧������#���������)�H�_Nq̓4h�*�'�@��X"��߅�������@�ΗMҔ�qqQ�o��~��kv�7������>����P~jLW��#��m�CDO�ʩ�`ץ<����$Xc���n�*���y�+��^�+�D����wu�H+�f5�����{���
��T���~���q�e.õ�6"A��z�mwvn_���"Ï"4z%�h蒝!��x{��+=Q&��<Hr}b��;���se����L�hhs���g��>�l:�j��x����r�����u�w����������:�}&�Ղ�-5��v���D�Q�L Y6Ap�Qa��s��ZYd�j`�G6�ݴ?wq�1A��M,ڕj�\M���W�Y�/W�tӧ��5���>�c�4]��� �p>��^D�Z�2*J�U������io��p⿽�W]AYӋ�9WEZ�b]L�H[��Kx�sz2���tۼ/�y?������J�ǍS~ �|��7)^�[�R|4J�i��c󡚷Z޷�O.�\6��Rr֐y�/!��]κ���;?�U���*8OY��¿\e/����}ìs3�}B�/P�w�g�F1���by]����c6���͢v;�y�X���nS�\��;G�&���[^#у{s����=^���g��aȳ,���>�h|�����R&���}7�Ɩ�/1�����v*����mяE�j�܂9j^
�C.`���?��fb2L��j]
?`�� �L8�(Nϟt�����d��')�?~['��׏���t|~�GQ�,����
����E��}9��TgD
&{�1v�7�C���$zE)7���M�TX��g�8�c����b'�:S�����`��pcx������o	��%�l�m6"�`�N����6�M t����~��|�~�6s>�v�zݱJ�zpZ(Z�K&�b�Z[�@��Or���Ug�ɉ�G��Iר��j7��G�$���|��\h�#\=y^g����ۧ;�o��Ya��1�\^��ٹQ0�0`��y0`1$8����G��n#�Ļ��P���rr�:ؒA�񮍉7��%;�y�lc���n�V��@��d��ɝ�	��ϋ�<���	�V���		΋���;��ft�j��O��gq��v�4@�ki�F�"�$\ݵ��ƪ[�z��z��I�z2et�@�[ψ�Q�[y�l�Wq��y�)���/"B�K��P;�%Et�N�}n�<K� _,������'y:����s�뭮�JspMi��]�2��h�������e���v��qiwɇ�0��jWo~��K�ڛ��WU���O:R���M���`=�-Lӝ[�2K���[]�r]��)6�>9�T���r��v��!1��W)J/;S�$|N̦aCI�;�K��4��i�IEō�������uNȽ�G'�a+��2Vs=('�t���t7v�����5�r.-�IV}[kV��ޗ�1;��_����4�-ؿ�hj�1N�u��V�
�E*�n2[;R����r^�2�;7���t�>M��O
4��V�ԯ�}��dj���f��٦#�p�yt�Xwu�`�3uX�����U�,h�1K�j�C�2�����xoxH�c�9B��l)g���Y�����njk��aس�������k݁�L�$0���#��[��w�ֹŚ/������ؕqr��1+�_�n�}F,���Rٜ������[��`BnR�z�]��b2����7OνT�ښg?�a�۶��������!�P��w~/|5~Ivy�v���g:�������ׇ� �}��z�]]��)@��J�i<˩����"� �J��h��w�h���-�폸r�/�>��D�J�$m��N�XK���\&��l�S�$�#�e�d��ܰ��2SO��[(��I�[�%��-��Μ�RW!�%47$=m�<x���.t�b�,u1(]�L�9:�+Z	ʖ�v�"x���];��Ĳ@+TSW\�;+��)h�
�'7��ͳi�P�Y2��&K5čV�\vAjQ�Y��u�0�o�8�9���	X���~�Wfk�u��`vu����Ro0iiU֬16��(�/uj.?�r��-��u�;U�̬=Wvx�'\n��L��Ow&W;��氞���`�9�|8iWo]��v{^ѾLU�����@�f�w�w�0/���l��t��1�۫yǚ퓙��\���$$�6s�a��JʏhcP�nj�}�{"��+�'p\����v�]%�����+��v��$��Ր3m^b�as��R�g;�ׯǳ���6.nr5͟Iȗ�?nw�s3 L,���+�}}^cI4�R}�{��&�|�N�y�<��>��,!��C7:(�/v�e� {3�)���g���	6��&�x���s����n����M�h��dD����)�ˁ���U։�&)"��Ofpx�/�䘥�zθ8�1�H�z�(h��tXY?�o'�[��4}]�e6Qm� .Q���5��(��) �>+U�R����9�������`ă��K�HSܖ�vƓ����i�XȘS5�B|{3���Y)J�J�����
`{f�P��Jr�=+g���s�&�3h9�yӹ"��'K�u����MX��f�w���:�������:�>u�u����1����ӟ�<�
�!�Ձ ��'��W��9�>�(�Z3Vo
~���@{��+��|j�o�կ�X�z=fO�2/KW ^� wz�i�;�ms��b/��f1b�Ed�fR��[�3\NCp?��D�EڇFa��H���&�r�	uިy��.��yC#�22A͞�`�۾Ϋ��i.E�a����M�7N#�	dL�^ن�͐+F���˩n1�"�����퓛�fT�/�)��8,��~f����x�WY��J��o�l,n7�%��kG�?��F�_\)�㔫p��Mcu��7��̜�reb{�xCp�=-|>���� �io�(V��a��π��*�Ö��Pq����~K�����>t#�#���#~^Ӳ�(e�>Ȯ4�����_�#:"�sʘQ���^U����\`)��A�1W(����4p� 5�{5\Z����m�f�����nӟW��;�q|�\Q�Ρ�nL%v�ms����@�����ᗞہ�U���\� �_��{�����&&D����tl�`�Q�R��$xB]徾���y�x�9����s2rFn�ڜ �)2ײv^�s:�swZ�����fy/U@��_s����=E�C��v��}%+��:8���y�h�K^u�=�K���t�-	�F�2X���?k�f�m�u���N���Ɵ(3��ǽO����������1��b2n2��������7���v�s���(d�\y�㇏���>j���.W`/Z�z���.*����.���3S3����d�+T�２��cX�à.�+
�����e6V��wiv��_��_dN�����&�g�0t������t���nog8�X��:���H��v=�;6��CзeX�������6ݺ���]f�e�kS����=R�Jʹ�֚�zL���B[�j�S�F�L�*ICnu�_�u�H�+���9N����bA���x�d&��	�� 5|	�UVGkj�}vP�9��ؙq�-��өA�@�]����ܸ�º�CJ	 �f�).)�i�����&-Qv϶M9yE��.|���U8(�s�>����:�L�"��)�&bڝ��B�r�R/r����Ӎ��i����sNo	#��b�mV����,]�$��\�Y
�����W��o�C=e�z��O���N���}fGߟ43O(���<;dȌ;��WXF|:�`�3�:=b ����R�ѓ��E�|�0�����(W׿R#j`KkDZ˵��������.�;5?Sq�� %��x�(~��ɦ��+8������m|�[wM�L~�}QQɡ�,$�AQո�����DAuy0�&Ffdb�B>��Q5�<�b����<*�9�i�^�]zO�|�g��v���C?����(%��l2�R�7���t����8����	=X�z�nd�Ѹ0��Z�s���U��g����4�|a�emz�ϐ0�����-n���L��4\'o�5�ﳳo�N�3��\+��n~u����p�$��h
�/1P9B�<��{ �ϧ˲�]O���k�t���т��>��
�bM���>��q��#8)\���x�{<�レ}���<r���*�$D%	�9X�kX�)kbn�6�ʅRp4
�dߗՋ�T^	}�d4�Rϝ:� ���Y��G�3뙌S��m���)�2�߮�mz�h�ﯽ����TJ����c,���a}�>r:���^�����KǗ�"ӡC���_et?y�������eq��ޝ���WX݋��wg��t���pZJ�'[�Jx�]&��C�ެy+l��8��s�Ր�[i�w<�ș	T���~�l���w5S�(���l�#�t�����%�����B{����Cܙ�cc'2�/��{砏��T�]^�*��f�H��(@}�ԑ擻y<�{�p�^�Ț�>RG{d�K�|%���믞��>6��1�s�c����c��ٽي#c���ċ9�]q	���$�����(���}8��f��z��=��W&b1���7s���c���x�ŵ~�U˖9��އ�F�槖G������[���U�z���J,�0����k��~���"�U��f=w��)��K�����w�މ<�V}l�6~��L��Dl�"׸7ʨ���w�۰���6�ǽ�ƻ��������ezP�	�ep��8��`�f:��R}��ԟ	7��t".�V%��oS����mRJ�m¦ϋ2��q���Ub��f���Q4x�\|(t�(C����5�;����џdU�������
�"}W��(���%�|kq<���mɏU�K<�(�.��J�s��ί G��-g��Q��rzX~&��O����"����bfm��ZCφ���6�<�|��0���������2z1v�66:|Iާz=���?S�Z:�IB.lDT�6~�G5���&��5!ԯ��mn����}P��:�鑙+�\������*2�_f�ֳ3�M���s���C�'�,����_2�p� b����Qfaq��$�0��k.J4����Ч0�m�
�6�:5������V@U��OT�%���íR����$~���ts،
v��C�Ϟ���ht>��9�=�É��6�&5�X'X�,,����;V����s��>�P}�#�K��\/�G1��.���l���ѨL{=��r����z/�s��f�8b��T̈́Bt������"2}Jx�xS���f����c�A�`���6Pd7cL��@��U�����W�m;��lЭlX^S;�����~�x��h{��W~�=ں��Y�f�e�>��qgz��	�Rp�'Z�;i�Q8�G���%4��"D4d23>$��Z�m�����#�6LI.|�0�v���/Pq���}}P��y�����H��Tvd�����ﶢ���KRQp܄}X*�s>�z��"�#ϯ1w|�ʯ.���7U3�OFݼ~q���,R�l�#����4�}�'���3�ؠ�0�W��cg��ο�ݳ����X~��/�}t��E�Vd�~���ϫ9�R�}�`��xI��%��p��1��}f�骁�۠(�\B���R��3��d~iiOQ����"�F������}$��g�+j�nޓ!���L�('.��<{��#�{��n7�A��rN)��:V<>�1���bQ�`�Is���]��3�Pb՘0����Δ�B�++���	����Cf�Ȑ����s]�,��|v2]&/�WV�QCl��	`=�.�Yӿ��F�ǃ��1J�R�{,uDs�.��� ��v_Z�� *���F�Avww��3�� �Ȯ"�G	vM�$X�c�z��ց�÷�A�깑uW���K�z���Nǵx��vQ��'����b��2̑�<ǣ=��ة����`*����]�v9m�n*��V��>� �\�ț�K{	1�1��09���@�f�yO��]&���M�˿��Q��b��F�!���Y�\әuK�����g� �9��~�=x
�ih�(ĸ��\:w�'s��S]E�&�]���o�����fD�a���ti�v7z��)oL���	������
�nkH���������u|�k���I�{>2{�6��B1C���w�AT=�?�*���T�L!�MG�����r���رs�Zԏ��>J�B�S�6 ��J=�a:^�O%��q=^����,�'�[�/Vh�}1j�h��? �ٻV���}R:���m��%� 1wS/"���R��Q��R��fb��/�t�f�w�-3��4��Gq���'�t��˰`�x�O͡������Hq�W�Sx&f�/Cs�o:P94��hŕ�b{��������h�
޻ �@PiH_� S{�/��7�J���`H��s;��ʻ�9��(0 �E�x*me�ݧ�Fk��� �n3��1�6�2�c,�[,���]�����9�q���R�c=�+�n�{.�j]���ΐ3h�ҬI��$q�`�y�2�]4"Õ���h�L�)l�F�+9Uj���ثq
%Qùi�>�����vYkU�!RUF�]�e�Hh���
\�/�f���K��!�m��7υ��B&�[B_��Kt5s5�0	 �p_M�h��w�c��څ������l,]eB �֠���>�:�y���
�z������ī�+Ta��1U�a�j�r ��s<�6VT>�I�N�=�2��D�ő����X'I�{{�><�-!Q׋o�a<�+��^W�k���!L� �x�=ѹ���7�y�t�{���>�|/�e�D	�߾�	>F�,ߵ�8>�>`��D�*����.l5�;g��a�c>���8_�h����a�d�{2Qe���(�wI�����dz�L�G|=b��I9W]79.�5��LZ�뱡��b�0l)W��᱗5O��L��D�f4] ���٢}�||$��=�gef�>���j�vrbݠ��܈�<G�hB+P/}�	1����hk����Y�/cY��1���+��܎��B����vl?=.D��:d`,$����~�]�";:�4�Vs\vfG�5��J�WP^��{ԓ�vp�P|P�9֦ڮ�s��K��m�ؚ%���ύ�.�Z�{��ze��C-�L��
1;1ݓ^W�I�e�cܗ��Lc��y�7�=h�CWJ�p��!=&\�?��S��|���r�=�k]"L^��!1D� ����^{�Gy�mzʑk��9{��7	�ǠR�;.��;��x�;�m������Υ�hj�m�L,��a�w�����0�T#�������-�/��v5NGm`��n�v�32�!W$�P)�iw��.��C����>?ݠ[����^p�����B+�����yl�w5��iz�ɽ����o�(�{%nf�-�-�������I/ S9�
�ye`�j�A�rӻ��>�v:�r��e�B����7�T]��˽=8���:>(� �W���_])��Jծ�%��QC���_#��YD�~�*��\}+�,�2p|�s�M����>g�C#)��¦��_ٜ�@�_D2Ȟ�E��8#Ξ����1���LvdGDa.
tt��+��Rf���tUw�jt}��LG���U����SFhi�{�ݷ�݁I�D���k��C���U��f�W��e����×��!��r��.������/2.��ʩ�C�4�"I��S������:���˩�`��5\Ey�QX��3j�� �Ϗ���܀|r2��0�25C8N)u��]ϻ�E��7�X�5ڔ�7����voR���3p�dS�R��.c�������B���]�3�fMw��t�˓۫�vTX�d04��LxS�)=/3�9�Pzvr
�� e�G;j$��"b�YN��׉���Q�cǉ���[X�y`����ux��&P�X��0Vm���q�,6ܭ������{��9�Js�u�6F�����ܰlD3U�F���h���>��e�������%�,��X�'k�ffRҬ�06��������X2�J*�ׯ,߈��c��=)Jk���p�De0}'��͜�y&aW����rm+�<���ƙ3�nq��e\4]i?�O�Dl����׭e���"/��7�������j*&�D�O���r N:Y�Q:�E�Ȧ�
�YM!�2S�S�[^��a�9f��ۆ��5��W���[5��������8:Q��B0�;�p;v�w.���=^����/����k��C4���E��M�ؘ�iz	Q���٩�5���;EzDmȆ:E��}u�|�U�b�>ň�4�خוOּh�k�����`)�W޾�N�o�l^���-��H4U2�ӱ7�Av�vO�$�}kn��{m��y���O��yБfэ΢g��.���T�(��d�e*��ևg5��R�����9��L6�1�Ƒ�����DMw��q۶�?h+ot����}9�]Cim�LV{��2|K҅!E�Ifr5�~\���'������N�H�F��G���koٙ旭O�|��4�R��{2�V�W&����/t��<�4dᲗ�^��Y}Y�]�_n|=ZjL�CLi�,}2_kՖ� 4�[�hC�:�X�ͽ�WŪ��N�Y�<��(�n 6U�k}V0�shP
�����&�:h��mFy��{7��;9C(<� ��͎,�[z�6��W�ExTu�1��f� zSA]�k�:;��}W�$�ǓIPF�ò�����Sz{���w�����=�bx����}Mx�m_�� �wr���<��e�7�a?�>�8~���4h�0��1�)eM"WlC �`�F�*aq����|�r�Ͼ.���_Y�/_�ۈ[��F��=�]{�����d���̪I}䧻��ϲ��g���W�N�h$��}�����hh������*�5#�h�?#�Ӈ��잨^=m�N�vu� lWj���՝a��z]��K�[	Wyp�����a���v���v��� ϻ�9��3fۡ�c���h�l'�h�����۸�����ֆV�^�����$T�C0��R������)} ~ WY�O�-��uW�]���nWÂ��-�9��I�&���L��a���7���1e�^a�}{�m��W�ӕ<�!﾿����� ����a�׹��6Q;��������u��v	7Rx]��>�N������}x�u�ǟ���վ�An8�r~�����Kߦ����?���J���Wd0�YD#��2�M����}�J�� 4��a-x�g��T�՚�{T��į�|�n�W���z-?�?n
T*������W�?�u ������U*K,o��Ty|k��@�{�T}�*Om����T����_?/��w?tR�b�0�H������R�m���뢥@�׏��*Tw����*T�e*��L�*[/9�k��zg����@뺥@雦_Mz�T��@���k?��Z\y嚥@�\]yW��P;Ye�J�ˎ?��e5��m`*�� ?�s2}p#\ǝ�Ua�QU����}eQQUm�I"�R�D�F*�JJR������((���R�.�U!F�UT�*��"s2�bR_            t (          @    P      �� 
   6�^�>���yt+�Β�p��E]��ʛ���J��O ����d��*�iOy�{SJַ�(�jv���� {��Qm�jWm&Ǽ����	HR*
�=$$��s��åQ*Hq� a�t�$q�^=�ѠQx�B�{���T(��\x��dU1΀

��ԗ�T)Nl$S���)�<�ڔ(P�J�B
�� z  @  ^
(P�22���B���d���r"W�5E��7%y��
R���� <�JQ^�I�	y5$���AT�ȩ*�h�=�Hz4'�"������� �v�U*"r4�X��*��1"��P���RQO.{���8����zۜ� �E7��o.���U���z$�we��ӗ������8���f7�ݷ��ݹ�Ҝ�"���y�͓�^1��a�+x̺�'�v�E)JS�  �      �̊ɣ��4<�n֓�"S������%��3m�g^�,ؖ� =�׺[miy��vk�Ӻm�Һ��y�G{v)�׶�ڳ��x �U��^�z�Q��ws6�i�U�TV�6ۗ=��-�ػ����{9� 7�v��q�;��n.������U<��m���5�8�{��Sb��o	���.�;��[j���w��d�y�짻6cA(T[j�^   �   
  ��ֶ�����)���;�UkN;v&���qgKM���@��h�J�ڭ�5�e�m{���YJ�a��vVV�K�z��Ҟ���AJ�r�N4P�"�l���K��l���{z�b� � ����е=ۣ��픤=�z�j�������%^�zRm��[m�y����j�x�͖Q+�v�V�̒B�QW �       ]�JV�x�:m���^;�X���m�ҨS�{���� ]\ڰ����@i�{�f��ۅ����m)�-9JX�x {��n��k�U�-{���mi*6ĤF��fӖ]kUF��=��dE� 3;fޛ����)�o=�^m����l��oE�t�{5����Z֤�gW�EV��0��˕�U!�`9)_ 5<������"�`�JT   &�&�54ޡ dh���R��U ��F�S��*�h  �� ��P  ���~��&����<)���G���'��:�ެ����s�w�w=�(U:γ��T����B�<�UJA�IH\�~�����q���q��~W6�[�%6:�r�0�m-?�k��C��������("ơi��S�~
�v����J�)�s:+T2�\SƓ��S�b���4���ă��2�M#́V/x���C�k֗��+
�t���2�8������h,Tf�u�Z���=JdN�Q�5�	E\�nV>7� 2��CP��5[~�nB��7	^�m{Z��kdB�Pת�M���S����\	��j��u�B�5��|:߀�@\/U��fp�8���kd�`^�Zi����t��SK�4ЬS�l0��+Y�y�\-YhN��� �l�Jb��_�~�c��u�2�oN�dǁ��PE!B�-�MP��*XB��m�ˈk�ц@�x&��Kil�wB`�"TÀ�A�� ��9׶�
��!TRVǂ�yQf
�2�ԇU���)R4�S+�m��k� �Y1kD{����6�Y��*3e��ѵ3T ��;��T�[����L�ˆ�[��.�U=�
����2����YzV���2^�K;���P>� �YZ2�jqD����K�r�l�M�ۻ�r�V�{��%�Pi{4 �!-{��=�TqC�ۋ�w�LTY��b����eУ���;JI{�lN�L�x��Q9%t��iT&%)�d��)�%�!���d���N�١Ǘcs��kHt�z6��U�x�Sw(�[k%J�Z�&����_�եU�o1�Z�PAcL�ի&�h��*J���f��B��A�v�2�L�l�ځ���-W,Qn�Z�>��Ѹ�(#���J1�V-�T6���i��b�V��ŪvLGf=D۩�d�IS�BE�-��8ۢeb&����WK+��H�g7R���(�_k�pLp,N$d����MeSSfҪ�j����cU���'u,�M�/e�.�ԍ6!�ʩ��iB���L��9u��h;2�j�m�0����!k�^�/j@�R�LY�Rb��hG�"�1S�:Īn�-�km�F�ZyS�i�9��g�T.�I,+�Z[f:�m+�!�u��P�ō�)��hJ�tuMoN��٭���37uM��,���'M�-4��!��J�cF,[�2i�XVܵ���6�m�n�A�����ZI+:�e��n]@j�P�]���Ŷ�šƅ��a�tik"c��'���X�j�4�Y[��L&�V��n�4�m�@�tr�pk[3_�6��[���o�9z#mM��nYM�2j�</f*m�ԋ�s1�М�pY�&g��K���Zx���i���e_�ɒ-յWC��ԛ����0f�v��Y���[u�յ�%��tZô��:.�����Ӱ�(ʉ��;�ǂ£�C�7V@�(����Ze��{���3��Z��T�Q3A��b���+X��,�J��/Be�9{�o��.�o-�Q�":L��d8�d{���hy�G(���^�MD�
Jlax��T��y��u�e�{Q���ڪ;�F�ov�GQЩ
����S�w�^iP�L�����S�FelH���-AU�'��i��YL�{I�L	�(֓�"�ըH�0֫p�sb�����uiՑŐ��{-V%i��k3�&�!��Λu����re�A*d�*��܄�����T��j�X��d.3L���K�i��!y�H� ��k�(�� T0#]�$	�f^�3>��/��DYU�Ce��Úyz�Q7��rB�L�<����MdzbNLZ�e��ֽWv��L'�� 䀐8����6J������*�,���н4���:).ᚘ�{1VŶ��;�0�)��^�iH�"��I��I����\ݤu+�
]�Ֆ��j�)�c��w
�ifhVE��D��#,Ԯ��x�G/m�+B����[�.��uPҵ'1hf�ؖ?����zd.ۻ������k� nf���Zڪou\��F���Zv��A9�x���A�UVƨ�u�������EȊ�׶�{r���h���9LŶe�hϲ��w�qT�NmD��ei�8�TDق�Y�5Ё���qF�(/'�f[��fX.��9�ݱ"��R��ۥu����S9�������طH����,C13�[*�V��iу�c"�����gA̗Sz&-�4���a�[op�Y�B��Ai;���*��Z��Z�7�	��D���.�-"�x��+�4B�cIf]W�����ݧ��R[ ��i7��u�
+�I^���A��wR��zm���)6gÖT!�o!�p�k�ˉ^�2�7�w�����8fT,ݽ�(��2�r旪��Fc͌4&[�P\X����\n�XV��ZP�wy����^��*` PܖQ@A7hn�lЧ[xf����I��x�ݼ����,���tH�rC&�z7�P�.K���v*O�F���;�i��%��Qg2��2�F&⦪
i�������O5`����R���Y-���J# ���z2�:ӌ�⻡o1պ�r�)[�'5=�5%��3x��p*6���Q8H�&�-ĭÈ�ٚA�i���n;X&�k&^�*,r�]�cF%6H3�v⫢���^J�$�!��&�'�M�ɋ�d"���${IV�a��ǭK@kJ��e��[�Ƴu`���壪]`�)VM���(G�H�L�Z�Y�T<U��ɮ�Wt����V��� ������ȰZRPOZW����P�%�J���ʚ�J�sj^k��������p*@� �I@�1�$��U�i&�h�J����Dc���1�e*pj����,G�+2-��|��%CUXӥ�ʳ1/&;�����s5��ʥ��B� 9oV)Cjd���ڬ{���-��b���[bn�n�T�j��nZ�Q�vT�ґ�J��f��V�K�B�oU�6� [��C+l����MQz}][q���L�Cr��E��xJ�ݝ�X��MZԺ�p�:*������H�somRV/��	W1���hJ���[VE�ҊN�j+���P=8���i�'!x^�̑W�)Є^MZ-�6����\����J�%6�A��ѓ ȭS�k�)¯G[�q��V�t���.�wd��ʰ΢V�Щ��f�c.�5x��F�4&m��d��cϝD�`��;�B,fkzX׺�ű����sNA�n���7q��`Ù���^-(Im*
 ��IR������%�i^���8�kK�!@ͩv�������ڈ\�{Սf��U��dbX
���$i��,P��ZnM�xU�6xku�������X襣+m��l[�*S%����kwh^kZ7/��3,؅@�r�dP�E�&��]T�yr"�b����dL��QV��)U��2a��T1]6tc��	h��E@!���a�%��7�ġ*K��!�^bxڳ��M8�ҕ��UɠRڔ���l6�hn�h��/u�`Դ^��2���`�ED˵(�1���u^}H=�U�v��t��h֢���1s!�ܠdU�r��ݱ�Z1͉GF\Z��x�B!�{c35��8hH�	j
*�;e��3/k��oj��vh=��̷��l�tAx�6��9�2�!���F�t抴��J��ۂ��������^�KW���j��d���I0��3X��c��mђ[�*�2��A,���,'t]"V�.�*�v85S��X�Vӽ�U�e��#�1�+U��%h�M�y�v5���t�L	 ����Tw_c�AӖnڂ��Ƕ ����%ϯ\��� �X2֪8v��S�Y��[c���/!�!�9J�nò�$ސՒr�IT�94U(�.��/-a�3�/)J�m�'��B�TN��Ԅ�xF:ۋF���X�":�R�,����	f!��V��X�Y�Y43+#Ҷ�^ɪ�o�e�&������"�#�|���F���{G!�P�*�*�l�J\����w�����Ђ��D����0	��6]D�nͧ���ul������a(5T�"�*�WF+n�4��f��I��mX�]�*��cF鬒���^[+q�V��a���D����X�IJ���!�aAm惩T ���H%�0��!�k�n��-U5��[dI�V�Q%iR0�Q�0S ��ɔ�������bI#W�aW�Tv�� �N�n `U%���F��j�r^��@��R����h��E4��b�j�̶�w��٫+B{T7�V����ưy�˳<�6�+iiP�	خ�S9�X�7�4I�{�r���*�A�[=HҼͱ�4�DcN�\8/��u'��A��A��BU�1:كK�4M�P�r��1����fneR1�{���x���\���2��>�K�-�`����هJv1Zu��r�����8��E�f�)�����f���J�i��ب�t�S^�`f�Պ�N�,�Xk*��HQ%=��a�y{M�sh`�tȯ4M��h砶���]��G�U�P-�sp̶r�M��TN
��n�p�re���Յ��Gi;xV��KV�I �Z���#�7ͥ�Z�r�bs��Z*�*���"r1�����E���`Z���|��L*0LR�ha:������%�t\-���Oj�ُE����P�c;���1���Ӓ���V���,[�n	M�h�Q0�U�M�x��e���\�ȧ����Cj�[�o&�y0���~�j9>+����F�k�,�op�oE4��fɢ�����u�fl ��G)�%�Ľ���R��ТJ��`�ݹJ���ސ.�Sc%,��l6�Y�����aPAE���a�6�&*f�j�zkN&�E[tF^ip6$�h
ub敥���yL&�S��-A��a*ƫ��mùSY��i5��C�F
�E�nVnJq}��h5���֑X�Ƕ�,0��f�1���[!��2��#�4%�V��l|�W�f#�,la۵J��V�jǘX7�0��ɸ��Pl�9��-jl�-��/2�{�[hޥQ/�07�-uCMh��Յ5���)P�a���x�� �*�a��J��Љj��t�����j�ɱ�E��XA��W���"����<z���8JR���[z��^mm�6�pℑ�s�&}f�MQ��%��k7j]�Da�mE���)�/]����q�/v�w""X(��,��k�W�ʷD����
T�(�TP+/�)��4�Ul�w���R,A� ;��jH��#v��E^�*`�.X��*Axq�Ғ��Z����Z�1��VR��G�͎1oL���Y�%����ZSF��m'�L�0]�f�1k�`�ݙT����T�m���-Q��7�Iϵ�x�NҶ��I��_"��Ȥ�!�3��T"�B�Q���l ��y�1Nျ��'����֜�)��l�m�%(=*��
�'(
kRh�Xse�U31��W��у3E��X�톩]���r�Ԧ���X���J�k�1�DVP��e�[q�Z]�^�/)"�����oU�M�z76#.�ښ6И���
T���,Kʓ$cv�ZX�ڱ�9vK;6+CP��+�{vh�c�n}�cb�Fiķc�4���M�c��e+ �(�M�Ep�k�f�c�1Ԓ�+'���n����V:�;u�M�Ð=X��=8�pߦr̖uE�E���R-�E��N��t��>��y�'!��m��6Y���S%J�o)vkͱR8Un�jbldTL(J��V�$��錕�QNݩZmL��r���vZF�լb�1�Q6K{w��3�-{��ô�=X���K{B�q��Y�,	f�NF�T(��9��ɹ����NZ�R�X��M��oF���(U�tí\6��Ya�+wd�Z��}.A��Z�^s6*m��k/I��V�y/ ��o7GZEU}4�f�V�ʄ��8��9�h��YJiR���uTF�ẘ�f��͘4�@��@ڦ�.jѴM�x�D&�PZ:��Eu�'h%�e��IC0$
�fX;N�D��.$f�h�E�p��o6����UL'.�=V5�^�X7�a�N�XYֳ�sI}�{����(nA�gv��w�h5]\�aa������[xNMlW=3,� �J�Ց*���e��8c��.4�uj3��������V��f�x�/\�q�+��oR)dzi�Ģ����q��z�]k�S��t��ZN4�֔4�.����iCW0߹��k;�E��Wk�%�|���Ф�vi�ރd&-����Wۍ�On*����ɲ�!�L�̓q�Keu�D��h�R���g^Z��<U�{�)Ҫu	��^��)�m2(�2��$�t�����2i��Y�L��/wja����qͺ��Icwi��������*F���`�=���q�;1���{8�؅�u�F���<{0�ܷ��ľ2-�~h�H�X�t�a| ] �)�0h�=�8C���n�ʲ��ʟfG��m��ۉѢp� �Z0�6���]���C��!$��(90�.���̻4��(��k�:��
:M.&@�E�d�vOƅ5�sn���	u����%�4���p��0n��r�c��K:�����2o�t�N;�M��3Ŋ��7Q�>a3�ʦ��� fHYjZj���T�EV޻�q��i���ZǪ�h`�B: �!9���(�]��l����M�A��Y��*H��c�w4�kUir�rE�.�0`(fS֜j��e�Y*�m�n�<�Y����H�ޔ�U\�C��`�Wbaa�.�2�v+VtU].��.��M�1��H
g3��V�m�����EE�e���v"�Z�51\V�l��^Mڛ,k�l��h�6�n�Z!�\QWzݭ�%�Cu��/~�wV]�v��Pȕ����Z��2v���*һ0 ��U%V�T Flà� hj]���ջlQU(�����Q������j��������v�����+�9jU҅P\K�TUΊX��m����Yg��-g��%W)�*U�7k����hխY��� .�ki�G  �]�VU��j�U�U����:��8J]
l��n�K���1�#O��(����}�o#�ݹl�7:�{i�Ӭ�v���}���}�G1��#y�x'd���xϘ��n1��/�ڸ��ȷ���r��ΣB.�Y���C@�X[n�v��xײ<���;n�g���؜G�CŖ�]���^����{)�@)�N�'�8G�S�m�z��ǎ�nt�]�N���I��݇;�.���1�'nN-��]>Nm�uu�L�og��mk����n�p� "�]�Huۆ�λs��nۮ��TO1�>:N5��c�狗ر	�twd맇�b�q�=��x8p�'��.��v��Y9��N�KC����S���[�`�v5nynی����x��8�yY�v��ݮú9�\�coF��Om���mu�7�Wt;ɖ-m��n����v��N�F@�M1�M%�H�(m4OM�Dr�����"n�ٛ$P)��{1��<�R��<k�%a:�ϝr9�;m�.���<Z^�.ݧ��i��Nץ��]���n�Z�uʍ�W��c�^��G��ۆ��-��mpm�Ͷ��g�j�h�u�<��,Y6���9cy�p�ԗr���\�4�������δs�*���r���`����[ckg����6Iŭ��6�ۣ�C�n�3�����78؀�*�v�a}��d��h�o��o�q�ڸ� ,�6�)��puteM���Ο[��"�q�������ݜS��r������Q��g�F3K;��Iv�&�;��X]Z���<�xLͬcik���vw[9F�u�,�ٖ�+��˺L<�vYs���KU\��.�EKgH�����l���sӴ/nQ���c�}�8���q���*b;XNWd͵>6�1���9޳ӵv����{]�rq��S烗�F�E�ޣ[��u��s�n];T��s����[��Ӧ��>-fY͋�g�X0Y�dd��lnQ�T����r�������̷=��ݠ�u�&s������n=S�������;vÝ��m�pL��s�yK1�޹�wY����man�W��J��v�Yӱ]�L)ȕ���ۺ�����bG�M��!��n�n���{�|��F3ClrC����`�3��ZP�<���Ў��8g��ӷ<c��&G۱����\���9Ě.T�;`����Ԟ&�{N�O&�Z�E�Q��u�˨�m�1wkY��z��8�Ӻ��D[��$�*�������Yݜ�ku�K�^��nM����rZj��xH8��m�}e�uWK&��s��;��5NB�Io�v�_V�i��av�p�n�OD	�;��v���8�uְ��]g�s��fLOm�=�kv�������͞|'V����ն8���w>�+�hpy�<����I�[��g����\����g��HR��@BPu8��Tձ8�"��N�!pj�lg���m��pq�N���V�th�l����=��{Y^�{W�v����;f�d�v���qm�&�%:�#�i���b&{m�N��qn��ɒJ�sڦ�v�t;oc�T�8���'��lӝ�Zw��i��PlO=���;n'H��7k��ף�y:l�w���ao;<��,%�V�ۯ�;'[�6�j��s��dҁuH
�Tu% �cE�&�S��6����I��=�˗����"�7j�[a�8�܆,qְ�w<=���u�md�^�Am�?'�W|��n96�w;c�������X6�Ǧ�B��c8�W����t�m�gƜ�纨�+Ì]���e���c%cz�c�Z��p�v9�Ŋ�'����軄��D���Fõ��v��#<�u;x�CVY	磕�~���ؓN"Z��V����1�=��#��Oh�n:5�;\b��=����Q�<����Q���N	��J�݅J�c��s�Q�O�\[r�4�#��n�Q�@u��\W[<��Z��;v�nv�bk.��Sq�5..�{$�4F����ݵ.�ݼcsvUl"BF�r�_9�7�X���р��^��0�T�6��ݺ�_cZC��G�Ey�U^0ZpTx�˥��y1��;<���n��=�v�����8��M��s�^���v��;jw=)�덯.㵛X�ûpP<����=�OP�G=��n�Kt�J��ݶ4gk����\�u�3s6+n��!g'Iu��y�"��g��^���d�g�p�n�노����u�Wk�ċEڏE�h�w^��wg<��󜫼���*rwY!ε��z�vN�nlY0���0�E��֝�m����!j��̠n�<�eǷgj�n���v��ӃXOq�r�;��ۇ��v�3���m��f�l�H�7;�l�<�܃Mֻ����}��>���]1&���u(F�ZN�Z��#�o<�:΄�ܘ�{O�;;q���cH��Wk��
lUn�d�C����F�.�Z"h96�t"�%���.4n��Y�q�v�T�9��3����T�Ɠ�q�v8�NgR�3�-��/5�]�gg�n�ck��S'C����¿H���`MۏΧqb�K �mu� ��V���$�L*(����8n�\Q��W�;�|+��)�Ѱ�7���c�NI읭����I���݇��Lm:�/�kg\4mƬ�:�pd{2h��,ݸps�����M�� ;2yj�9��tS`������Y��Gaق|u���Sqp�K�{��v����[��!�nj0-���>��<s=���t�;:�`}>�p*����jۭ�.�gcy�c}��<�.��s��{uǤ���؃/+���9��V�܂�:�4�;�o��v�/!��v5�az��:�Լ'9���[��d�֘m�X�t���U��2b � �Ǳ�猉�]G���!-�K���Н��$:y�j�ɧ��Ӵmѻ!����;��nw�b�n�u۫5�;�ɡ	�F�d��n3r+nP4��:�9�t�܇d;z�a��=k�avں��\�����u��C���Mb�R=�y��۷i�^9��|k�ST��&����A�1v>>�m���$��lޕ��v�BJo&v�'�;�o��kmz�aw`��ݷ�V�
��v�y�K�9�nyp��rwk���6��N��p::�Jp<�Ʊ�vS����^�\���1�����3��=�cn�QL�M��琤���m���ʷ;`zӝ�k����%�d��Z�p�7)����F�T��I�Ŕ��h^Nb,R!X��nU�0.  ŐBS`��+�+�J� hvHmon���][�xѲO����u+��sղ���=��8��wksm�Me�Iv�t�v%��
p��A�F�t�::牋��2 E��y�ڝ������:^]���l=u�ݓ:�8?_s�w̮���r:ys��2ݹ��F�n|�\�8��2;gb��V�2[-Il���j���Gnɺ�K��ݨ.y��d��Y��9���b{[q��^9�o<�9��p�6�w��v|�s�,�&�X�%��;���ݶ^J���@�/����v�y�v�p��nV}���n^��c
�wRv�ok�c�vn���і��{n5ײ��7Z=�=u�;��ݝ�2Z�pi�̊�3�ub��<�q�����'�ՎMp
��p�POr�Bv�H�t��mNÊ8v�YٷV(n�����ģ$�;���]��m���v7 Uz�^8������V�5ڹ��NS�/+m;=zl�Y1�\v��'m}��#�]5n����]`���d,p��3n/i�N3sVj6�B�n�I=�l�#[�k�}��Lj9�]t�ǉ�쓌\��nǓWu��v^���n���u���Gm\a���s���s�'H�8�ŭ��E�Ōl&�P�֮R_cp����cȃq�f+c[�ź��q���Mvy�t��&���m����˻�-��^��iʞ�jT.�)�ST�����&;6[�U��L<�WI����+��I;h���9¹0�����=e��5�%η�{:L<�q�������<�s�v�M�� ���۴�*�����lX�OF�,gw=�d�r��K��m�Z���\��Z��6뇮%{&��3a�>G/E�a��8�"��a3]����y����ޔ�u����'Vt���l��[�Wf�ףH�-�w=�rQ�s�\���vP|Ξ����.���o��n�ᵈ)�'��ɬD>��l�c]��q{<6vǋck���l���{(K�a��O�ψw۞��L�ƣ�����Nw=\l���(�U���6�NY��Լv�K��u�����bG����pL��k{�v�#cbu�q9���ڠ�{Gil��G��t����G3�:���u�ϾM����+c��'^�Ol;\���"ܣl[&��8����pڍ3��i�m�o`�-�b��}��f��o3VS��y���Ѷ�n�OV;F�S�y���E�Okc�{q�'v�8���J���ys�DS+ۮEf�f�qu�oW<^+0a.���"� 	�=�sq8���� O�&�.�#��j�n7ݱ8�|{r���m�G<�7n8�zv�1�.����� �����q��۝��2u�޹�qE��V��4�RG�%����`������:�xrog��.^`g��S�����^2�}����qN�u�<\�^P�qu�'�Wg^Ӥn�műp)lkŲ�Y^w>ْ`6)�n�;=����.���/%d��.t�V�������c�wo�7"����gs�s��Sm�s���n,��Z7��lt[�:s�y�G����$r�ٶ��9qɷ��x�m��^��]q;��{Z{m����ǮMҤn��\�.y޳������u[�z���a�;��Z�Ѻ��z�o3��N^8�b�h��T�N<���.�,n��nջ�z�������h��m[���$o�����t��ET#҅PaQ^��߫n�Ch�k��2U*�!K��j�*�VtT���YZ�s=�sۚ���d��yӎ����[:��[P��D	c����n�2�V]Q�ۭ�&#�m���n��6�v�6@+uTC�VM9�Кl��`D1O���	����W6Ӱ6�0�k1;n��Wo<���P�m���ٽB�k�(���zz;9�����n�iB�X{#ƀ�t�˓���������8p�w<��[K��yJ�m�<tggm���8;{g3�[��9|�S����]J�rj�Y�������®x�k�q�헣��N�v��l�����0!!�����uN��61��T���h��f7e��8��i�,�*�U��,m�ۓN�i�p�Z�ey��63�9�X���C���'<��MWYޓ3��nC4�Z�3�zػg��c�
��X�b2���aR/k5!
 hsNU]������V8iϞ۞�\�+nG�����'��2�x;q�h�qv�hW�=�;���x���:�
rt �6-8�ҐL��D& ��0iѸ���j�	��ŷj�q�Ŭ�_���lfs�&�'[�#��Kc;�4y#/l�
pi̖q����;݃Ŭ�;��]=�^{��&e�S���۔Mjq�n�ޢt�n�pF3<��E v��=;��>�%ڴm��K��K7�����ۉ;8�!�{u]lm�}V��r�e����Em���^CRY��U˃E�ݼ7�U����ܻ.�Z1�YѺ�<r�q���W�@d'��8�{1׵�4qm�5=3S��d���wf�r��`B9 �8۶��[[<dԸث��p;tZ�km,�D�����m��]�`�8�\I�q�[�h7V��	���]�rgb�^Lj��KvT_a1Us�v���Gm^Y�Kd\�{u�Cp�u���A�1ׄ0i��6-�nݤ	M�깊m�6���s�5ȕ6Q���y�a�sqɶ۳���A�kխc6s�q�ʊ���(����$�ֵ��k[��nn�dt�),E2\cu���n��;2�my'���U��'�|��=��v�vѮ�8�Q�yn����s���=�<6�i��y�L�j	��X^��st����9�
m�|ٸ����wa��eM�nm��ї=ss8{n�3�u%G�7=�o��u�y�ڼ]Mƣv��ݷ ���+`�`����[�Λ��wn�޻�;�a�5M]-i�f�!��C�CH��rv9�o��woa�Å�D$@0DQ�����_�M��Ӝ��+A�E��J��wB:�^�l�F{L<)Cʙ�&s�o{|�*M�0�l�[�%I8�@׬?-�5�N{aU�a���ex��{Jz��@+=��;��Y��}�Z��U��.��X��4��*<�g�"�8ᝁ�S���l��q�iw��n������j�]X'�u^ҽ{Ҝ�q�L�*�R��4B!� �p�
H��_�i�Ko�:X]�H����5`X{�CP��/h��uZn6��ޡ�YR�hAΫ��� ԇ�����!}j	$�ZM�4�������mr�����>���a��f�]�9^*;mu��ѳ��崞V9��|ﳮn�,��4\�4���:��<\c��J֔�6u��<�VցT��+v�$��	#fI2�7�d����ᖼA�}�3Y�?jx�]��oDm
z�.ܯF��H�ߝdG��y��P�1�,�������o�`�9��}��{Ѝ%�vB
��]!��{+���uJɴ*��Q�2�V�r�;E�f����jN�{IF�jv_	b�7�Z�,(���L,�V=�{��-���}�S˖F�<=X#�Dm	���|�b&v���9�a���r���{�7���Zڋ�`��B#Y2���� ��*�s��_��D��?bn�M
>��r
�VB��A�(�W6ҥ��Y���,~�Ay��xQ�q�h��>i�li�iX�$���ٕ�-yg�vxk]U�j�n򐠙���F8�1����n8ag8��*�7�:s����Y'=�a��~��,NCg�槜�Χ�w}7�d:#[X7�;&�e����v�f�x�;�筹9����j��oq���,��dHG#�nI+ê�=��ګ�����OER'=�>��M[D:���ev�۝�nΧ����5��EL9
�*˒�;ʕ{a�۸�=��gy����7k8�g;�_B��5��d]^*�֘��ۗ�^v�羰���L'R-�9Ӌ��%cT�3{�n[�Q3�7�	��l�.�;�ҋ�\��>ܡ��ԓx���c�,:'r^�R��n��2��i,������9[������{0��m�\���:��Ku�Ҫ�E�������N���Aďi��=��wʨ"�ޫ�P���C��fJ\0i��A�E�P�u�ʪWֹ���/z�^�zZ���f2���]�����̓GF
���YcJZ����̖��7-�io_�mh�K�r>(�A�-�_^���]����Dߎ6��	'j�)��D�b��=��{6�m�����lq�fC����1��%8l��7�����Sģ־)�*4��̮��[U���RNq�X�{��VT�ԇ?��h��8����WL�()|�[O��k��}�2sIE�Y�zd�y;ћ�W�e#Ыi�_k�]f�Ɛ%�a$�!�8�Q��H�^��}��Xz�z��u��U�0<�3V߽8��Ux%S�iL=Lc���po���Q�Z,(Sq����(xT��jb�.�&5�s����@R��e�od�=<���G��㺳/�]�~������y3w*�]3��3س3N�.����4$)�g��bь�2�d�����Y��@�v�� ѹ�w�����)ox![[b�0��i�!JCOBD>����`2���Zx!��Wy���0f�Vy����3�7�g/c�R�.��ϊ�ƺ���wa@4L.u�Fuӹ:狱ֳ1�xv1��z�t\�2��1b���-OELrƤ�MIU���~��	��^M�H�w��:wϷ�7�a�/v-╍�t�nd){�j�m�^�xy�J&LF̐�2�Z�=!�Zv<�=�V��~�u�����
x��aC	a�w����3|�_fu��{����L�@�f2�(\���
>}~�]gZV���J����}�x5��#y�����=�ї��N���ӿ7W�ROOy�aq0ܑ #�|�swhG��;�(��[�Eu��J�y�+�n��=��p�-��l(Ԯ��m�'v_?R, �ĂQ 4�f��a��4OT�$���\:��ٵ�;�)��/˱�<I��C�TD7|$�,��{�y-q����\Z��Z+�v��wf�p�O��_=��6���\|{�g�ܽ�+����u�g�H���=4=��یRA�&$:��b�N��6�v�v':�V�d-�u�ێ��3v-��q�,\&z����}gQ��E���[�Ϭ�o�kmk!9]���{n<n�Ѹ���nϧ������cLe�n;h���.���lZ&��G<nZźP*
ʨ�u%P�S1��T@��P�4Skn�'��"`Ku��n*U��h�X��ŮJ1��=�kP�v�ђ�!c�cvռ��=d���v���9ۛ�g�6y�x�2�]����b�k��y��U֍n�s���aJ�^��zSqnC�ފ�r�O_g���ť�5�ѻ�S~0�_����U��)��i�͆�l�Nw�3�T�}���+�B��	�?yH5��FQ�G������;Hc>�?N'y<��
<��oT�,*��l��-��;m��r�;\i>~�=��{�<�4�d��]e�ˌ<7�\o���/�y���f��Np�Q{��[�h6TdE���:iǆ�Ztk��#�O{<���5�J����WO1u�gy=͙��@聫��&!Z" �M!��x�--��t��$_]̅�p����H`2��|�]��u���9N��vݖ����۱Ҽ��P�������klb���8�Eɑ��]g�䌸w>�n8�Շ�!����`N+�!#�/<4��g�*.W���(�dM�[[�O_Foԝ�^���mM<�y<֫Do�Uw���k��	�$~�D�9ez�z�.��i{���s�:l�闛Y�ܫ@�����B�^f�}t�rv��{�(6^���
�w�)�ܭ�4��lے�ۈ�Xf�u":ڛt�dI�K�D�"��3Y�jVsJΗx
sp�iFbh���/#W��<Vg\Ҝg����v�i�a��q+��U�2$W�40�z�.��ұӳ$f*2�q���,Ƚ&�*�����=�֌�I<>����&���𬧽D���B�v��9ָz"-�>\�P�ݪ�'@�>FF�E��}���Z�\X�"��<f7~;�L��ɑ�LWc��Gg����;`��/٘N,���j[�y�Y:[T)]�9S�a���w�޺���1���v���>pZ�n:��oc���j2�NB���uWl���zs�A�k�|_�i����5�˳C·A8���?T>r�ńE{}��%H�l�l����JgOJ��՗}�๦��/{YSU��E;.�p��s)�U���;�N��՛U3r�����Áv9%�1��b/���RD���>O_����w:8U�.y%|1�1�X*G	f�ķ��:v�:��|*j&��؈�v
��bWOuű�w'��%�{'�z�Z�	��{�V�eb���T� �� �Z0�.L�!�+cݾƨ-�n:��mA��,J��\wm*���}�p�Cs���\�ias����v&�*^_V]�8J(@���Y��C����K.��=��BX�%ӽŷ�v����M����.-�)�k�C�F��F����������r��v�+sv�/b탎:�b���*��v�ȕ�(�.�=t���#�u��d�҆�J��]8~����[���}@K�u��^�ʖ;ۂ��|f�	lD
�K)�BҎ�S�U�+�3�#��~��^��*�dK}��^3�wf�Pm?:�Uy����MFa1��jG�޺UK������߬ ̹^���9Õ컒��l���VA���o��2�;jp���äІ(ӄ�ˁ9�p��fO^>�y�^�y�W���ͺI<@1Qe<�k�x�,w�K��u�/xܺ1�5�o5��ŏJ�^�gY��Ȯ��"P�!�Z��z�K4֞���ا>�wVl���s�M����N2�c� 1ns�Nw���t<Y��1ĂA%�H1�:w�1��U�u�Zaiљ�z����.�0@ǅ���Q�ӯA�E����Ґ�u�Q:J�O_�����B�n(ؖ���s��С�]��c���/ j���.��똊Z0DCr(�Z�J��tuwE`.�xX5��]}�5���Z�U��syS'��_����[�R(�Ėp5c�k3}:O,3�e���Mm��+հ�}=�j?�����a�pUP���U*�K.�ܣ���;9�yxQ#��l(����jȳ4��T�.]����A�kQX���1R�w���g�À�2پ�`�����d'�}���(�SF��y$���j�P�F�����y�|�����^<���lk�+�w�f/j�l���l��q��/�O���O�uWn�DT�o8G��r��yފ��`./h�8Ju>z�'v�GV�NqP�]S���(���ˁkp��P�<�0��K��y�Vŝqj�Sm�X.:<년�����ѣo7L��>��ɿ��S�k�nf�M�ڥ�s��.��<<V7]Rh�H �͸���޲!���u�\n�f�ݑ��|�f^��t��v�l:�n-�L���k�?t�������ܩv�n��Ƭ�Fs1f��٣��rq`ù�����[���oG7n�k�6��M����qή�yu�@m�y�gdc5�N<<�^MB�e��籲���ۨ��FS���Ga��nt�3��h��Dq��ƶ�ee��3��z����_�v�?]��6���7<�Q�	�NRۍ��pGg�U�CsZWV�n[������������7zqoxG]0���e�M Z��~�)���9�p�[�����~a|�,�TCE��d�N)���V'�6�{J{��}�h��N)�J��O1l�5xv.��h�^ᵀ�Ըy�ž�l��1�|[�u���걠���	)8�P�T7lV �3g��S`07�_���!�p&���Y���U���-w�>��͇�G��;}�(���*����pBc���C������Ϧe������g=��o�m-<�w=��vxG���Es�7x���]�ڦ�.e�e��/]�_f��"���90�ΨeE�n�#�S��<6���m���
�%�����q������/I	��w[�7��/@�X�#e(�E�t�p=\Z#����˔�Ɇ�UW�#-��m� E��G��pc���"�e�?[�^�d�,�����X�Id�pI�R��T�_iM�	�1Ĕ�HV{�yu�P��'y�����~;N�5:JH�o,f;zgk��x��˝v��Y2у-9�|�>(uFIU[��N\��fS��}�DXi��4���;�����iG�ܮ+�#t^�"5�*��)���H�lɈ���y^����p��ȡ���r3k
[�W:��+=�s��f�����$ʞӵz3�OD�f9"��G	ڎXb�>�
�5Y�w'[��r��-�t���á��w�uK�1�1A�l1�{�빹�Q�2�Ի��4.�LQ�A�r
�����r�K��6Tܦ�Ru��z��7�YTS�^��;;SIץU�]��֗f�C�kϓ�x^��yMDV&F���if7u��nyP4�Js�n�5=�۱m�C�.+W�a���
��P�r�]2n��	��s���B@���㇗lMF��ې�֖\��[<����P�����~'/���[�Dm%��Һ�{�^G��M�V&�.;9�#CaBs���g"��&��{��S�t�4k�馇9g�X�}�$i�ĉ@ӌ_s�sA���<vDlt����CO��%A�:Md��
ȴ ���-�'\�F�1�fB��ۣ�Kr N���Pçhn�N胏K�=[���8*�@�c�C_Ed�U�]�e�c�L{{Uͻ�Ci{%yW6vgq��y^Ru�Mˊ�*��7���&�=|�*d^�f+�}��@ҩ3�O�����
��F6U���8�|�n�z���/opt�uĶt��9���/79KU�>F�����7̉Qx�Iy��D�ތ�{yZs'�&�f���w��+��N�]�s���D��;�l�L1�Es'��ڵ��0]��T�3�3
�0���Ȅ�\b���ْ�D�c��vs|�-����s�z��	�Lևs����9p3�N=m6ȱ�XCA�a݈r�;��7�� 8���-Rn�{�m8N�v����;Q͛�Ƿ*��gmK�{������#7m����طKoK|Ms�ﻺg+$
)u�T����l���}>�\{��f����'��{��6Wg.�x������K�2�ڠE#�cH��7�@��f,ʜr�����7��ؽ׳T��s5(�
�І��h��l�׀�)�7}��`�Z���RK�n[g0�x.>Wֲ幏f�jS��0Wnm萫�嫙�P1ĳ&��tT�r�E�޼��1F�w۵��ee7�r8����X{֫����&�yzR�mhr�]�	gze�R��$(�!ڑu��O_ܥrm�Q���r�`���yiۙ�,�ֆ��ւM����|t�8A$�[�l�4@����4@�g�/�)_G�L�8������L�䯻�D&���E8j�0���>���/9�~9Z t�}��F�����'�����φt��|&��M �#�"U�>�=�i̸�dQ�[ IF����<�t7�H��ܾ�����̆Q3�
����;kdd
��Ӕ�O���ή�-�Y��_O|��A,�39�� ���m�ѣ��/��FDn��8���$.^fb`
c�h����� A���#>��2 ͟|B��>U�__]�[/*����6����{�e*G����������;p��^m�G�ݮtjC�Es�u?�\0JP��K�>7��zs�^�e.}G���+P��mџ"O���BO��&�#�gۆ������H"����g�T���}6���M-�҆�(��r7;�Q�*ۖ�&C�|�Rt�G�Q��O��+\���R���>� ���]nq�΁��}�3��@9Jb�$?S��"��@�
O������ςn�]��U373�}�0'J}5�$]����)Tr��t^:*iJ�^���|����k���z�}���&��g�1>�4Q��r��V>K�Mb ��_tX�+�1�i��d,����M�c��t��n�������~�#�vjJ�S4�i3_
u{f����\�.������|�z�ּ>�[��K�>�.�@g�H�2�	�d��ْh6}d3��`e��y��C1
a+��v����m;;�;I���`�=5�zN���4̙x6�v�f��v`ĺ�1�Fz�����y�8D#�o	 �pN���*i�a�}��Wxc�r8:�j��z�6k��j٥c�T���]��"$���|&W��$��Y��I��X	=?��H�dxn��R#�ָ+� %���wm=�j��kf�OvY�OʽOϺ�@�\��� 0IhD�@	#�+�I��S���E����t��D틓�n������}��o����zχb�@2�n���"{��}�ax3���ح2���G��s}�@f��2��څ�����Q�J��}/6\�Q�ha����!'Ȋ����i�*�Y[�Y�C�s�^�\4���,�uI�	�:��Ev����>���S�7�� Qӧ>�����n�r>#ǍpXiC��6������p�k�M1Z¹�3�MD����D�4E}׺J��U4B�e�ޗN
�4��{Hk�}�'��7j���m�A�>�{��ר��c�O��%�rx:tI��3:: ���RkYߧ��"�6|������/�M�*( �-�g�+�7A�o�zoqa�ia���[h�����}�>b��>P�������|�T�(X�ӟqO��"���,�@teUͶ�t�ӧ�eΟ��aV�RbFZ���j?1P�'Sn&���_F�?q����P�<��f�6Ķ'^ו~5�fׄ��EV��G�b��>�0>�� �2���6k^?|N -�i�u��H�0ٶ�@�I�C����!�LY�Ta�Ud��O-N��:�lQ<꯭��Tլ�8�R�''g�q>6���;��*�*�)�t[Ցh�+��O��2�#ʉS�Q4�m�Ԉ����r��l�n�v�΢|�/i�K�x�u�Z�<v֕���L�Η�x���b8��ґO���.T�CI���f&y��0�k.ƅ5��ێ���1���u������[X���G�/����E�{�nK�].㭎����o:��!ϫ�ܥ@ٻa�bM����+ӆ�b�]���q���oF�h{n�*Of�ʀBZ,)�c��`͂x�Wl��X:���� +f��ι�l�p��{���������� ���/xYJ�>�uB>/�Ȑ8��"�	,��Q�$�6��>��Ȑ"-.�m�V�/@ϭ"NP��D
4|>�Z�NU_O��V� A[?I8l��.��|�44�n���I| �����.VV��>E��j�6`M�C�^s��(ɓ'MDw�2h�#���D|~�>ϐ`�'o"E�,�
(i�R�C
�a�윭T$�τ�T�Q��9[����!����b����H�q�@f.k�"�!ľ�F��q����E�Ð'�|>��$]}�ft�"����t�ܸ㻞9�	;�s�ىX>�ß������s>�ޗ��b��4��S�����ӒƆ��7^�*׮�g-xQ��8��P�;W����+��91�|��H��?|���#H�(���)TY�Z�[�'O�V"Z?�n��,�P��k���>��D������ԽG�D�$�n}�DF$�"R]7j��D(lJ�P_����y��T\����{ߺ�LX.��>�wN�|~-�Fāt��ޟI}���K K�q>&�q���N}�H��h�\ՉW���[�G�4K4|O�^o��)H~�V7�.{4�;&GU+���=�\,�]�˶zJ��àՈl�ָ�ۧn�m��ΉC�o2i_��/����5����N=~������=*iv�%r� d���u\ۨ����~ ��*ؾ}�~6� q�MV׫Ke��7���!�و#g��66�3*<*���w�Y��o��y>Ģ�C.!��:�2�����U#4�ZCQ�uyۡ�K9��z<����&m>[7��ob�Gd�P�����#0f��H��Q�z��B>���D�7�WU;k��q+��%���i�o��ް�4�6����[����6C$��CU�{��ܬ��A������8�{�-I�n�H�����^B>$	������!���ҕ����p����h��׫��e�nr0y�+88�q�|��}�^��V9�0�5��&��?�[��\_����zȣ���|���p�Z%!
E��AY�婚4A�j�3i�&lލ�� }�s�H������I�D3�M��>�� I�$H�R��}�@a��G��p����˼Jn�`ϡ����kT�}k���CO��֦�Ğ0U`��Tv5\��YV��k�a�����;s�D�>:���|5��^�"�y@�m��ww�}�×��| �g��ufD�r�ׅ@��r|2z�ȮCqX$�?��ҏ:����/P��[���M�3�]a�s=�sv�܆����F�n8�Ύ�����DD�i��s�����1
>C>��.�zs2�'��J�g�|"B��#�	>���Hy}��O��d2T8���_�}.=jr_QO����ᆏ���Q
��M՜�x+��>׸�|n�O�3�� �`X6�9f��/�g�)� �R���>��hl��T0ΡdQ3�"HvW�e�2(Z�^��G��M�>����T�g��@���H���qQ �ӆ�����{G����$�w����6�vD21�Kl��Ɓpfg�{WY}77�
�>Y�^&�O\2Hߢ0�>���Uxn����5�><>�Z�wn�:8�mz�uھ<�9e'�����0,��55�E�PH�b�s�q���"{o�]v�:�����W���A/����s]��J����l������d@F� χ�(�8?C�H�EU�+ޗS
i������d��Ƒ���2�U�>jL�����񏏺��RQ7��@G�^��}L��+�u� �1P���!�K����A�$F!�� a���$T���2|��"$�zYץ�}ذ[�<����4�/���/L>}ω7�_��t�_!2���h$�?M^���ydG� am|@5S� ���.�����A>�~��\!���?*��x���꣺:j��M�t޳�-�B�B%�z5j���#��w�I| �Ot�g�Y�ɕ?e��>��<|>��6n����S�G�B5;�O����E�N񌞀�IQ|��u=�",!�
������ݿx�5l�V���m|���6Y�g�q���3��)�a���̂4�A�D;������ttx3����$�@��bC!�GH �V8��p� (��$1J�,R�	_}�j�r����\5������qVqʝ���ݫ�� I� 0z~̉�*�� }TυL����\�o]t��ϕf���"n�h�,��V�>gw;�����s �I��VA#��Ǫ�2~:|1�x3쟣���_U�,�4��6���O�sp	}T�M�To�`(��q�1�.|(����i��m�4��l��ib�!�����՜&d���u�:p�3DP�u���ѣ�cm9����DO���^��n�s��\�Zh�.�Q��I�Xs"FY��d��v��������73���T�p�S8�S�SO�����{��Fk����	l�
�_[ȢڌlDC.5nJ�f(/�O����և�%N��f�&`��2����G��
��A>��"�}��#�58��K���gHFϤ�h�� n (����H�@a����D���
��A%�A1+.���\dwN�7nƬ�p�m��\q�� �m"g����Rs����A�V�Z�
#iXj�4x��؀���m�S�#��6%/��H����,��Ǯ���CJdt���.�&k�φ>@A�7K�k/�2E�|�b�.��Q&�AF��������4E>�F������*d�FM����`�s��'�����G:��>�eu7�H|-{:�Q��T�>�V/`2~��@�&C>u?j�y{���jڮ�jO�,4{���t��u�11���pr����N�,5V�k�.}�..��kb�u(��jL;�K��>׆ӏT��V��(ƪ��x���ë��|`^��}d��H`�Q�����ϣ��T�:��ɥ���a��(A���K���%�|OƉ�{]���� ∛�kz[�)���Cfb��߾�����0���W�g�jJ�+�2��Y���(� :���n��<ڕ�Y3NB_G����R��F����T@{E\	"����Kf�V鮋	Ql\_=�[�}��k�p.��Wn!J�:K����LO�|#�Gl��DJ�g]����8d�!�$	>�Q_GRI��̍>�DY$���x��>G�p��ެ����$s�!���M|k�Vtgr�o��,7�5#z�r��R��csvV-�bt�����﨔t��A���yVv??2�T\0�L�V�m>�	��n8�\p�c�
UQ@N&����EjE��&�:+�v6|�)ݨ㫂���/-������M����N5n���vm�^w��qG[�����>w���۲��C�on<K�C���l�[��v7nۊ��s�]����uʆ�'���eT2b׀��pi���ی��-2�N�Q�g=������2�V1u�g��fwA�7 ��
n�n�َ�Y-uҋ�n]�@��mu`�Z�1�]�2uR�K	-&*|j�b�V�kg���^W��E ��/}5
���(���Ϩ��ߙ�ϳ�IY ����GG�F��E`��9d|}G�>������Z����Hg�~2}9�G�XE���=-�=�:������p���A*w��h���"����Ï��;�K�12O�Af]I���?!&���W��H2��S�g��EY@)�3�d�_D��	���E�?V��,T�p��_ál[4o�|�T���m��b\5�A�'Ú�j�2|>��R4d��YU���?0�A�(,�}������>^�N�.$2�|$�"}1t��}��g)	:|/r<��3���Z�G���*jY$��S��|a��}?|����z�|Dʟ��厌� !u������R@0�,\��$Y���-Q��#���}_]��U����a��� e�I�?i�����Ă�f����),�)z��d�<u]�� �,2�N��-���A�����_q���ԍ$�"�����O�H���Q�}�[8��Y��!x��(���׭���8(*kc�����犚٥�f�޿!C�%9���uϔ�ohF�n�V����k]c�\qۡ+c�ų;bvk�K�g�nQ��]�ؤ@9*"���8�}��k��D�w@F~���}�h�4�H\�sK�MϺ�.�4���}�p����]o�Fs���u�le%���0��	>��J2}���20�F�@~}��+��Fו��T;X�8GlޗN����E�\Mm��c��soؽnsx�Q��#'#�3��6�5B�ɝy��ޛkU���W���P��k�fti�Ы���(�I�J]lT�K^��~0L�o��:$vg��,5���9�_��.5H��)g 	R���G!$}ѕU�C�C��Q9���� �������!G����B~-�1	3��n/XO�ٯƺAQ���}��L�K�XQx[� �9�|?�Y�����^Tp1?N@Y��5N�tb����ix�/W|�z���.o�|0�@�Љ�6`���v��P�P�,%��-������qB�@�F#�F�9YZ�5z?d���Y�>��9�Om�O���?D}�Ƣ~� �6@�s��D�ߙ�Ѱ�����uH��#�0�1}�2b߳�o���쩍�kĩ��9w!��ς>5�0�JGN��#��'>�j>��q=�U}

��<x͵c�w2�y�.��{v0�R�|`��ϕha��r���ʄ$�V�V��?�<�,�D5q�`�=�8�m9�>K�=$�h��V���B��;�c��W-����O	C�^u������b-+C�^���2��I�d`>���$a��>$#� ��h��� W����>���!�h���6EԌ��r>�c�GO^D� �m��"1�[#��(p��N�{j��	�Ͻ1 ؿs��q��]:inviR	wg�R��D%�$�:Q��"���t�2@e�J5�CO��ˉ��? �>54�T#sH�x%� q��hF�����n2���.��T�&Rۙ�� ;SW�)d!�<d�+��e������?;�$�"'�����s�xᔺ�u�:ibq.��{{�w�Qbܭ�R��B^k2�_Y|3��)���u;��҉�X:�ֽ�D�Cٿ��"�bnW��"H%����!"�����DY��6M u�"���^��Y�~�Sߟ���8/<ųV�����dl���f9��i��l�I�.s�r�0;u�L���Αƍ�7��S�=?F���d�
@c���<Q�0�C{*��\��|9�DWO���>��?v�;F�X�Gm޺"}�A����z��+�y�(�uQ��"�xk��AG��������^�����/�z�Xi�%��>����@a�>��CH��~ϝ�	8|9�x3᰼����
�I��n��J�L#�҈lz͹�ێo5�{.�+m�݋���E�Q��8�tl��)m���᯦����>�zP�(�6l���"M�ρ�1�2/�����P���p{��j��;��>f�-���Jy�}JN��}%F7'�8�7�:(�,��N/�{h���?�q�*�9a-���k�x3��@�S]�Q-zȬ�U�}ox�Q[�}hA���:W�oN�IrD�$"� �*%��3�f9���˾����U�I�^�kĈ>�����;�����CP$�t�\�3Ci�!(m�����L� �Z������ˉ��G�@�K*<2��A/�s�#/#�L����ϫ]Dh��:�wY�@��j��v��,�#��xQ��D���|%�g�YB�"��n�:O��XG
�r�ܷ�]��[T�T��%^Ӧ���\���ϰ�7(I%�]�!?=�D?�K }�ыMPhQc�.Ր*�ڑ`��Y�'�FJ�q�}�C��s�#��-�	ۭcEp�Z_,)�Y|o� V�0eq���Ǜ�a�]��16UŗG�B�?����Êӂ���}\�.C�i��#���ր��Ήg��Q�YcDNZ[!��"϶��D4g+X2�a��ɟ
>ϐg5}G���{��+�%�>��}�m�ź�"En�9 ">#�:}��ϲ�>����,���	(���)r5';���WꂡD�.v�#��:9���܇��72x��Y��u�{N�m=����GI�r�e����e��A�ƍ ���%�J|!;�Q���il؃S���4�in?F�/m�����)u|��}O���I��"e|Y�k�]/"9:�#)zϴ�>h�ćT�r�GХPl�RKx��&]��$��"�D/�g�>l�Wm�@���!������ݝ� QDI�@��"�9�d���$ɓ���@!��}z��ۮD�Na&I�>�����O{�(��	"Mv���8(-�Z07m�[�:�wqz[�|� Æ��n�Ș�`�^�;�a��TDFnٯC A$A�N����3Jc�JD�]T z>� |p��L��!��O������5�����G�46o\bC�i��-�J�6/�?5�s��>� ��8�o|e�>�_h�("�������z�;�%�����a֐$ˈ����Ϝ�������Q�r��-��>>���w4F��#�^��[��6�X!�F�e���Z\5����
�Pա�@2|>��F_ѿH�UtC��s��=
�
>�@+��ΐH���Yy�:�(�}��	�~��%�eY�,�7ǭ��x(s��g����5�/�lä�a�R��9��V��K�M�bv�+�o`N�jD�P}�pBh#cFŉ���m��#��kQ8N�b����,s#��:���~v֮g�_�r�H��:m,>7��������\�E���'�/u'I:��ew!|*�+��DÙ�đ�ISv}r��~����[�̈́�6*�ޅ+�:�AV̰�1v}jԠ�>��˹*W��������Kz@��G��_��_�ƭߞ��oO�|�X�8ԗ|w5�;�]i�����m�ujљ��̍�%GS�jf+W������!��w]�C�M�r�ү�3
����^)��Gwo�eH��"�ne�O�\��L8���oQ�:�7��J����h�xf���v��b�����H+�m<�U;��h��ze������ͅ��e��U��=�&7�V9lJ�}�F�����w�Y���V�ݣ�g묤&�Lm�-���\��m�W�JOU�9��;�4�i|�=�j㻃����sk�N�vѽ�q�B��J�`�sy��י���!"aj�T���E�D��Z��Og,��[���1���u��pͳ�`�6�A9'$n-�#��C���9�Ķ����_Cf�p8��u��D�����;�$��Z�Q�E�z��$�Xa5����!߬:U��Df�I��Vu��*/���Q�$����J"$W��;�v��c�����s��Y�JZ��:QxU�#�^�J��_0b��K��z�M���tg8t\���jBUj��Um.�ǃ�;�C���8,͡g�&;U�9���X(�R�m��U��U�C��{ �sue�1�f�xv��s�� �6�2F�9�C�
�/ZY�u���vˁ��
��)�,�s��낥%�x��������a�t9�+w�6�g��^Q.�I��vݺ�s<��c3q�skmt��3���yw�F,67�{OQ����A��mFn��/�� �{\�h���l׵�H`�(�f	�pz�vjuDJ܁�Uݵ�:ƕ�&��`y4o�v��i:��h����NM�����:#�c��0 f���JU����/Q��ulk�/�$��S��n�8�@;�݌���6��I.I�5�IIS��kt���{�:M�ˆq�)�;Z����aM��1���ݷs��֛�8�ֺ1ݖm�<��<;@�;h/n����3I���PQ���M��� ��Q�&"��,@n�l[n\�P�V������Z�,��V�6��=q�3Y�[�u90��x���{h��q����>:�f;D=��¾�Lxv�� ����ǥ5��4"ZF�FSƌ��N�m�'G�$�m^#���玍X6�;Eq��Í��{sǮ���-p����]����:�N7[��<F�g�8vy:p�����Ul��r�cۂ��#�����j:gj�{7!=�ݱ�Ġk66�N7
�\�]�]�.)��]���}���.��O|�\�q��6C��k��������ȍ2QYQ\��o�6����;v��c��tֻkCv�Ss`Ǭ�v7n&�R�x#5Ź���t�f���{]Q�s��s���sv���n9�Kwf�g�l6J�y��l���x�q��u���ҡ+�9���lL!�N�ݍ]��v̑um�\ɸ-����r�r[u���ž�_`�P��k����^�%��`L���Eۋ�k9۲盵[�oQ�g���\w�;n�몮�ڃ�g���sۛ����9��<����	��=%�gx�ݏ ��nr���=p���U[�����wm��a2��m�Nkv��=<�3f�{z{�N;tʫ\����hy��6A���7N�Q����)�����-�im1m�f�A�G��o�� ������F�N�g�!����B5��v��Vt�c�vI3���t�;��XL� }�'���N��� ��6�fݶ���Q�vR��@m�A���#W�Y9m`���,jv�㮺[v�[,����D��/��㦶%�)�s�De��>�"��7�����0�l�,�C�����w���7�>���E(�j���#�>6B>d"8ܬ �$m�����
>�7�M����.a�[Pۆ�6�O���oclg��6ׅ���m��<� b�xϲơGõ �YD���ӳ�"
��|$��5W��T��z�(�	d
2|��n�$|�=��Ga�b�L��/5�?=|��a�߄lnyq�8��!6�Y���	4GG�I�@o*޾�A�MjG���&�F_	�s��O��$�L��S�Bc�U���bsPmf��� �D�ހ*�a+ <���_/a�{(�o[4�����Zۍ�N8f�,��0���3���;(t$@1]|���ߪ='�ٿ�<(�v������r:C4|�|]/a����}$]�"K9�H;>��Pqj�YI���ߐ��S���ջ�\���O�t����h������淏>k��Ӈ�4�HI�%d^}8F��x��2_�D-9���o��+;϶��W�""�����hq&����4rG��x�$�ӷKd6j�s�~�]4��!�4�������}���\c�m��("V���{9�m�N�g���7=��Q�t"10����J]��;\���Tr���]5��a���AS��<�ܘ�(p]y�f���<�T�ɓ_�y�So�D���5�
�~Ϧ)(C:Z�+�&�9EG�wn	Y��*̟a�^��փ��,��>Z�$v�ե,�gE�g��� �mp����7#�j�5��輓Y�,��\P���(��͊�j�1̵�].��*�Eܔ����N�6���=��;��5�w�����u_S�Nu�/b�V������Y�Z�-A�Y���z����L��<i���ę�J��jg���{7ϻ���:�5p�\��h�)Q�^4�*!�3�F�ѷ���%e��J59�ҧ���[���O��ag�`�HQ�н�N:p��	:E��@<~����8p�&�sb�Ę+U�$Y��	"�z|��k�� |l��B��rG�aD��f̚s~cO������qo@.���>�E�	����j)�4�ř��EY��?J|{��R��5����r���D�dO�}�Xdu�>�(��W������������[��*^ri`�!�]*Ͼ<�"�M��)�5�t_���4��3��of����|5T��̌i<ưg�&���a ��GnK�\�FDi�~��_�j��B�D�"���&�6�K�W���d
�����'�I����8/_��������3�Q�%��k���x���Y�9��O�@p��u1�nӏRvͯ�	l�ذҤ�]_����D��ߦI�ߔ�|�H���� ��H�}󡇍�T�z���>�-i�.�ы�����-�5��soA�2ئ��	���"�;h��[E�4��fC0oT>��Uϴ��'����'gU!���P�B���s�)0F�hT/\* }v�H*��} �� d
�g̉{�`Y8�'u�2~�~��������8�2����}z!���FRK;�%�W�\zb1�i�Xa�5��9���$��MH��}�z��v(Q���^�]֎����34����[@�C�x�]XB���zƩ�+g3�C6\y������Z���l�#��ó��k�Z9�|�3U�ouy^�������8߷�ā`�̥$��҂b�z���ٮ	�ϲP��j������8�m�H�H�n\�O4���D�ϳ�th"�򾊒(�>�9��@�D^��3�"��}���E2),:p�#b��P�ޑ����� ��4��Wܓ��t�s�U�=o���J��O�=����')M�+t�׋���m`����ezg�w�r�~Æ��^`�h�����r��τ��&�\�d�?|Gփ/PP�Ps��.�3�(p������b*]����da�Ȩ��^�A��X!�&���#�o����B�k7�yK��9�. �Gj�S�\l�5�݇���8��< ���ga�4��v�D�����P�P�B�'s3�u�ϰ��-9@��G�:,���{V@�" �������!�}�A!ϻ5��L�i���l�����D|D��:h�"RȺ�$e��aI>��OD	�����=]��NW��wӆ�y�s�&E�== #�{��0��t� ��-^��Jc�=٩�w��x;O�TFEh��I�qgя�R���D� 2$���Q��9�܎:�|:�}�џ&B0+�rFZ�(�>����a�e8(��,��8k��k8il��:�,��,>V��1�!� ��&W��_|���U��ȍ��'�ָ�Gո�~��0�h� (�!�;W�g�:A#��ZL��<������~�7壘* �ϛ�����C�Cs���x�L�������[��<&SK���ư\>��݉�G�}� �ʃ�(�>gi��������R]�;#�b����M�sYSR��,�d�t�s:J������.r�����ݕoP�9�1�n�x��{�����%9˛2� <J�����s˸���8���]O©z��͟�c����
�G�+��/����B��
���<٨k/��g�i0|K(��86�쎯�b|�q)���!*�q0��>T��dP���M/ٟ�y��\>����va�W�����w�Kj��C0ఄA�=qs�S�=X���H�v�K;q�)n�m^��v���b�W*��J�r���_���lT���bbٯ�L��4�ƌ��I�Ck6�Y�>�����)G�0K����^������}��d3��jH�ZL�<|���P���Fev)��&J�0�����+qJH��*9l�8.ׇ��f��(�jIQ����k��䕁+{|�#��^�2��uYg�d����f�~"��������� ��

���}��N��mtG�jn B�#꽸�����I���FJ\+��4�I!'�:�e��K��Cm�xf/G\IgH��(���oׂ@㘅�̐��CL���Q�?}ۋ�������]��7����lS�C�I��H�'P���H�	��C;�Q�F5�uM�>�����-�P�~�[?q���^��(,C�&��=q_1V�,Ú���A����G��u"�"$�d��@V�A~Ͻ�غ$�a:��|":~�`�5@�Vp�D�$mi�O�b�UǄ\�|ho��}�H/���[�[�Ì]^m[A��[m�zغ0�o���>�*#���DU?�(a���0}���I�6c�X6�۪��������(a�~�u:Aa��/ݙ�>���A�!���T9yϦ�gqx��j�ȓ�cՆ��o�J&��%�+P���T�)$�L�O`�sH��C�	�K�����	�/�s��*]�ò��ߜI9_h������n4�������u�6�H#�n4��ެN�^���5�7:�m;�NOl��1�خ*w8���o\u����M�==�mY�r2:�a�n�i�	;8jl�q�M'o��َ�3Lۃ�5˱2�tl����.�ە�z絤��r��M��(4�՞��v�vX6�s�ll�=�K�۶��rs���lK�;�����iKg�*wj,�냇o��t�p��c\q�Ǉĕ,Âuf(ܨ�P������l�� ����5�\��=�&(t^F���X�ƻ�����g�Gܠ�P<h�BY�H�K��D��N*(�� w��$Qz���mW��&����R���j�4�:�~�T���]��\�!#�2�k�I���,�	܊n]��#B*~�=�I��}�>��Һ�����9�;Ǯ�?���ˉt����3.��L��4�H��u_}�"ϰ�| �"	!H��!������t��l���Q�޵��-������B�ԅ$���՟ ��As="�@"ε�(�:��r0��6��W��$�d�¨��;�(�tA&J,�]?q���^�eC^�̓?#_�oTY�����g��A}�}ŋ��i'H:� �A��X���r&�1�[�ݠ7PFb
�"�^��DoMA��Ϸ"GY�$I�O��v��D����}kI>-n7�$���Q$Ym��,��Yz�]�'�����Y�uw\�w-:I}�G��M �+:��[U[k��eNK3K��H�*y��g�3�|o�/n. 4���ɏ�*�����~ϬHl_��'O�%�[(9W(Ao�r,�3�aE<�`���Ov�LXw�������kf�ƅ��/)�7;�z�����,��Yv�n�w��{Ny���|�n�u��g��ګ��GUP�V:[l��.�~LE$|M�8�4��%����,At�>��e@�饦'2�����H�g�>P�j6��=P���DXV�j�U���I��$���(9^u���Q(�dB������Ƴ�����	-y��^<Q����s~�P;��s��p���ߡv�ӆ������.}���-�T<Tϸ Җv�t.�U�P=�v;�ax92�
��Ꜷ��²�\I�d�����2�6e�w�i>м^ڬ��`q���n����A�9��a��}1-�5�!��Xk�_}X&��P��j��7�����Dqó[!��y�?]x.��DB+���%�ƙ�a��{sHǆ���y�l8��XQd��ǌ�hT�I诳M{Hʈp�>�Z��B��5:�6�"�>�!�=:iL}��I�<�
�~��K�\5N�Sb�6 x����|��\�R�9jnىS�=���Zp�	�v�/7�/ߧٓ�5�~��b�61���(�M�CPG���-�K�h@�����ڃ�u�}��\����6���Q�7��M}���6l�]b4�F���i{��?q�>
V:��������UI�M�"�!?���^EB�>�|���ﾞ�Y�Od�)%W��f�}^�]��}7��{=^�QA`�0�[��~��nr tL@c٬0�"��Ñy=���R�|Jh���L��b�;�<��⺭�K�Q�=5�݀!�%�^�͍��M�$�ھ�ǎ�=�K:��A��dA�4�j��k�4�)Z@���1���cN�?M�齚�z�@���W�V�$��<U�*I�W�ckl��t��lk"<�|������Ν��>R4�K>�_>�@���<c"0؀�P���n��&��N��E�}����(���j0�?j�����	%+ nud�Y�[���S�o#�!`���|(�Rh{>�2(3kO���� �Kf� ��~�ž�9\<i��}�3��Oھ˸�3�\��֮ l�X~r�*�q�T��PM� ��-��^�M��m����[q>�,��dQA��r<(��gO;ϔ������4����~�P��[X&��V�B�'f�f�,�.���6��U�l#�j�t�D,��MҲ{��U��Y�l�x#� ڹVF���}:�"5:Ћ~٪dx( }���6u��tP�g�=p[1>���>+E-N��eq>�BȲZҕ���ؽ��/���+�Pg�R4�:��4�Ш�o}�#괌}��O$�}�����#����m�m`�w�ű|҈v|ԽI
!�����mwԑ? ����b���X��!�swHǦ ������ϭ!49i�����FQ�@��ښ�����E�iYsn)�G�pHEk�n���)X��|�tU�+W��>�!�� ,z_}�q�ĸ�ߞ�.N
g�2���0�#&��$QqtG*�2���,4����������9F�J���e%��۶�2n*Z�!Z�L�emc��ƭ���:餷3���W�������>�G$��AB#M/�܊>6�3Ú�&o������/~�ߞitK����@�#�Y\��uzf�����4������>��a
�B&����|A$�V@߮����P������~RXݒ�ʇ+޶#��g�*x�"A'�%�� �Jq��@٭#� ��*^R�oc۲�R-���� �)�XaϿN9���{w����Jo[�H�BH��E3K7~�H�Dk���FGg�~y:,�d�C�"�^%У��I��ç��S5�g�-��x�~���.��|-"㹳�@�
������4p�.�׍5�	��|Dq��ߦ�;��q�8Gݯ�ϾX(�?��J��"J$��
�9ˋ>|D�X�֓�&�i���pn}mQ+j��$�%�p`1C����2Ҏ�@�u�ߧ���b(q
� N
1O�6Bߩ���<j�>�
	?$$�B�"��d#��]S�q�Y�L�L�F���E��!>�E��a~���r�hg,[[�h���=ZU��]"�H3�F�fҬ�,�e�z�d�N��9�r�W�� �B3�4U����4>!�d|r�$���ݾܽ@Ylr��:�%��4.	�@�~ �'N�I�Ǎ^��3fx�$�!�bB͑4bo�H��0^۲�b>��w�A���$ĵa�$iz���U�xY��7+$��>�F ���u�*x�L���LKg�o2%���y"ؕ?B��|������-�E���m�:x�$p8�=lr[I���G]V�Y��<%D<��UT�դ*%����x8�<t�`����R�e�D�BB%I}T��)�����(Y>"yx3�p�I��D�� ]�ʙ�3��|&B�H#Ǧ�R둁�4 Y�?q���3��BkE@��`�6�ދ���uO��ZF�rQ�Nix��zP�x�7F}2w���~�8���3�s�]��>L�3���c�~��	F���^�ޫ�T$}gLϳ�CH|��,��.�~�L�H��K̃�|�&=�	 ��=ks��!�{����>D^	�{�g�_j6;*�U��ú�~lG?t�kg<������/믝I�41y�"���)t&�w��O�SGܔΐcH�0�%G�o�~���~�KIQ��~��T��
�f�4�b��CW}Ջ����O}L+���#M��E���H�"�۲[o@^yڍ� #k/�B�Q��#�^?v��h �>�fO�R-2"�H2��}J}ց���(�E��V������ɯah��ܘ,��I��Ҿ�Gs��'⦫5��di�6B&�a|-D�0@���˶ƥQ�]d�r��t�6޿�
3j%#�("8���Q2���4�l� ��H���c����o�3�����6�? �� Xt��Q'�Q���5M|+�>��!��5���L��@3qT�0�Fvx��һ�5v�:��ec�]԰tf�]�-���Bޢ6i�;��t����oz��44�Sw���mY-"��t�F�=���}�^���v��V�ܮ9Ԡ��U��i�+�i���g1��ݝ�k���vmջ<�k��1��F�3Q�v$�nw��d�zr��ثv�$�C���z����b9��;�Y���]e�,K�Q	qٛ�M�;�1Rݸ�
����^q[n�g�<j�z�;m^u�&އ۱�[��L|�qi��]E��q�з���rS���Ma۝��m����9|��:�8�)ً�V뙒��0��b�6�NWm�� _�Y�E�z[?�wu?����7כB�b��'���Ù��������7�DI'���iG��8 ��;G�N�ԙ����'#  D�@�Gн���͌b�5���,=��H�}���*�u�;	l��I�O���,6	>��F	�%�^���$�-H�6��E�1w�A��*cHQ��w�W��������$�Y��Zg�{��pP�XQ ����S[����_u?=^Dw�o����h�Z8�+�p[پ��!C���1�au$��B�L��gE��z�Hj���������^����1|p���N�����,���y���*�#'�Ϫ�ٮ�v�&h�w�)�<@=�ة�o�7F���a��h�(jU���Ō����	PH���[��-���8/�� �@�o�?R�'>�D^�<��%(�8��4|~]_6l7������Yȗ2s�7�!=��� E�U͛0C/z��e���g� �{���6t� �~�� ��{�Yǥ�ϟ^�����;��]�׉�X�0���������_�����0�%�I�(N��k��Ō�I���Ϩ�ݼĐK�IFt���?�Ԥ�aIw��@� f�"mx���#{z��$��k��R��ś9�p��
�� i��"��`�Q��͊G<�m�(�vݸ��:ܱq��]�`�)��6樲;i-���G�O��j٥��=ɫt�i������ظr0�����cؼh����pA��B	ף�J�`��g�N����g���3y�K8gW��d�Ў����������/��!�F4�v��ˍ֭V��%��uD
��,�^�0tQ���d������^�G����+?a���D��F���Gy[W�!��ӿ+�n��W7���MbĢ�vJ�g�]��-j�����h�˿Q�ݭ�b�U;[�ɤv������<ؠ�:,��rb�63|j
*o��������M/g���
��iu�a����8]�"g7�׊W�������L�ͩ����Z�(�F!w�>,���]c
�%{��͊��d��f�������8ٿ�Qnn& X=)?߳���vJ|Q���`�b���4���Go�L���=�h���2!<i2�&���ko�|�Y|9�'P����&�0HG�;+��cv�aZ�ً`.���`z�������S��$���{�3�!vG��<�q}��QR���s"�2��D�P#
2d�ˤ���{�~SD��{$5ݹ��Z!t���������ݦ�"G���4�>��@�N�m~�&W��K,��^9��Lk����}?H�L�~.1_s���8�	�4O��C�ټ�e^{6���@ξbI8��W�Qe�(S���ѐXE�>v(oF4�G���џMqu�D��<5�q��,�[^|�6#�P~�������:�v�[�fv��m��Z�m�mI��<�g�`��i&��r1(�������j�f����-�஀����3bG[;����hO���������Ϸxa�DX-!_T<H����$��Y�>��<7�?�Н���ӭm&g��&�DQ����葆�#�v�]���?�@9����~u��S������^5~i�!o�f�5�>?w7<�?j��¾��7���͜�@��b�u�)�͍��д��K���$>hDދo�ז4A���F�N��x��)h��Ie��[4	���x�r�#R��� �}�=�S�]�qR>����o����I��%r;��_Y$�[��ꊣP?���S��t1)��63Չ�uޫ@�����_KZ+�0��}|]�9u��;0�۔��B�c�ۛ*T��2:�B����B��u���:���O���չ�����EI��m�Y��m�$#���NxfkL��d<���ѵ(Uد��e�H ̑�VW
i`�6�\��[q�
^��Ցu�Jn��+��R�dqH��۝�Qv�/d�7��̊�+;�1�S8Zץ=kT��	%��1"�����:.L�X�C�
6(t-ϒ9�%JeKtͻk����d����>Xvf��e^܈(8KZ&K�1�����'TͧȰ��'���2L�}:���-A����[�]����'b2c��e<�Rh�Gq��us�E�cz)NtcFf
�Ɣ+m��6n�Vǽ��P���U�u����$J�BAU�Z8ζgs�Q�=����޳;y׫���J���s��}�,�Ֆ9u�*�"�b��n���wY���Z����v��v���Tz��ug9��;:z��b�oi����'r���«8N[��a:�5�S�
&�N�W_4���{;�����9��n0��>���W�z��)e���
Mu��[
Zv�,��;���G#�*��-V�4�c�&�m��m�:��I�J��35=;Q'�Y]o��ضb��74^��r�;ʋF��3���\�fXik.�wB&N	��ne{��y��v�F��}�R2�]pZ�L���vӋ�Sm�sE.��Zʀyj��ʵ���JL�|uԺΨ�2�TE��Ԫ�Z���y��%
nRq��U�%g�0�6���o����1fiAj�m�-@�v.�;���S杀���#��Qc�V�e:�ɱWy~lbX���g�ש���0��9$��XL��n!�u��;L_a���^�� ����>�Wt�1g�����T���� ���f�{2E���b�d_B��볶��f����t��Xl�P�$�����<�^Hx����tZm��X�v��Dm�k�̀q��f8�n/��3��OOb����7��AR�B�k�$�����R�Kp&{n��on/@4�jț��$���TK�<+�~�������v���F�om9�KU���y�׺�ڷ�m�V,�Y5k�e��R�ߤ��^3Q&��GE�.Oe����D��3��a�0s�s��s�?t_K�S�d��i�A�I!�:�B~GR"�m�S�5I��VPg�c�s=��f�͞��'�����
�:��\��4.�w��}d�]ٳ7ww�`��
 �8PI:y�2��TNKs��f���\�E���bWzI[|��;	>|*�=J�'�z�ȑi|X�g�z(^ahfo(�MV|�#�ݍ�ۇ
A���qԱQ�BJp�DS�9M���5�ڮg6��5�}Ն����[6���`g���d������$tz�L�縶>�n
�V��)���4;'=��!9'L6.��"ח���.i�`�.{W2ԑ-���u��ȣ�g�_&��椝�2!�,�Tv�^�<��L�$;���-a`�4ۣ#�5�["k��*�m�|g��9�*�u�����Z����$z9w���"��ʦ��'�>'N��������Ǔ[��0y���/��:�#G_t�%x�C!�m9��F�����0̞n�@$�0a3`T��7.��d\�9���˔���<$ q�I�@���[s�<�G�LyՈ����!m9����^���ќDU��[�*P��,��-A-��)6�O��f �1p]�b�v�f���`i�H����E(h\��'pp�]]鍂���X�hZRA��2YT}ނ���U19>�_��z���L?'�=���N�+��DG<�C�f�\=���&���[��=�}z�� O�޻�ؙ����驆�����҇@4�r5w���G�#�+��r��U���>�ء-7���z�{�]n�Vm����s��!h�%cJ���f�>�O�� ���\�N_+���l4��o���y�C.!/=��J́6'o����v=��ڭ|���Su�W��/���E8�_L��D���X2"�B��H\v�����}��,�t�d8�J8ݶ�^j��.&�z�en�n��.�Zm� ۏAs&@�����,to�>7��/ݽc��Y6z�Ѽi�ok��ucp!��k�����*���	�m��⨐���=z�	�����\�F��[[s�>�f.Gb���7Ck�S֧1;m�]��h�JW��\�on"k܎�M�ݟ]m�	�u2sm�Fy:�G/l�[��'aٞa�a�v=���ۭ�ݶ\L�=�^6�AP�w�������S2�\�]�T�Sz�1c7���.SƽքI���ۥ�
��W��jʩ�7�7Y�$f��Ob-Y�Iy���Y,���1�X���/S��{ؕ-]|r�u�����3`�3ި���	rBx�8�&�#;2�"��ǖH�B˞�]uW�OJ6Z�՘F��7�[O��YJ=GZ���\�|z���7����r@�& [U�"��>ݙ�(��Dm%�U����#I���	Ї�k��lo���z~��x�nx`J��	Ɯ��i�Te�}c�X����K�:�"�2�	�|W�dG�Loy��H�t�!b���7�3z\�w6�f��R���fP�UE�u�FJaH��p�kmqg�G��\�v���V�";���_�7AŸ����ee�7F�ȳg���U�/R��k��@���&!���̏���-��z�
"
���gg��Z��]�v��7`�"��:zj�Xc6�`�[��"R܆5�I']c�Bh��*n�r�c׊� |�f����Uߝ/Qgγ�\b���dµn,� Q��d���B��*yg��f���b�!w��[MF#%ȬO�f�H�[���8��k��]�������-�_�ٯLq�piK'E�[9�VAc%�/�Z�ŵ��s�ҏ������+���sr�&H�=p�X�x��a�ֺj��lG}�1#}�^���bj����(�;o�
W�ɋ���[9���^���K��r���:�6��#%6K�n�S�ug֔B�0�/{��(��}���I[�Yg���=osh�~�(Y�^ꡩi6��:u���ؤ'��U�ڿ [�I�"p�!��,)��}�^�.xKC�Q����0��t���h�{O����$���l�|*�Ǚ���^EL��뭺\�Ti�Oǖ�8�VPq���	�*"`#8�Uu��-2 ���d<�ŏ-�)�� 7Hg�s��u��nTt"(��]r��Y+�(<�M��;'�^ml����˫cQ�q]4RDϋ�q�h��֎y�l��s��w8����ٺ݌��*�E��{���J�J�>9�&i:���Ѧ�)1�"��ٟQ�:G	�/ ]>�Z�6����A��u��}>����P��Mд�Q+c)�N6�,ٌ�f��T}D-���H���Ku�-]�KH�H�s˦���2l�!�;O�3�tQ��>���TT�=�+Vu���g��G�����Ȓ�f@ڑ=�L�|�<3�o��*fE&j�4):�����8b˾R#�7{7�Y�gR{�%gw*���=Bjv�[̙���X�]�q�� '6���ͺ��qL'r��P��G�2R�[��Z�E�R~�JD�Z����FJ!����g�6+N��2'sfobZ�wo �|�,��j�t�������s��Y���2��J(Ԏ��*�3Q<�����,� C��uQR�s=���O��>�A��L!'4qj$|�#E��������M#����]#d��c��ɜT�3��%c�Gж?�����
�[l%6���D5�r�.<��˥9��kW�\� �8��6�,�ꗪ�kf�u��tE��-�������8�8���p\���{����/�N1{�U*�1*��=5u�vđO��}DA�l�=�z�N��ğo-����Z��ۻ��͖U��i���!_x�BlH"i�o
m�0]K�e1���F�ݧ�T�vTa���T�Y��>��4���}�I�K�D"z{c����J��a'�/Pä�{p^��@�)GT�RV9%2��=�|J}�b�.U�φJԸ����HA����v�+����阰;�'�|(����uf��@�Ss��m`�BԐ��f	�����Ϩ�֧͛�+·��>��ֺ�^�无�X������r}��(wF�	v?zߝ &��+��x�µ����1"��]`�Y5mv"�{q���(��fH�*�i���ǳh<�sm��O)�H�׻�@aT��:�+?	�r裩D�[w��1�����/����$���@�Ռ����W���3 � (�#;���Cf��װ>�*��Rg�g��՝.����E�!��g��W��'\Lo,����H�����6��OM����;Wol����Pت�
p0PX.�>ㆥ�k^
��T��t�Qg�L+���T�Y�ǯ*�����/#*w�)|�� �Y��Hy�i�d"q �J]D� �R�4�p�$�w��D��A8z��B�[4_�^*x�G�'}�k���}��Ow#�uisoR�������'�����O��λQD�L��ɠg',�@���ED_�N1r@�>���aӕ��s.��H���B����ڝ2�z˳�/��٩���B4
�v��+څ�ڌ>���ꈪ��M'a����x3�ή�_R�����c|�y�T4r^�7G�Kr�7��>W����2�,5��D�!
�`���^wP�f_n�����A숓ޣ��m�08na�mB��&������������W�b��v�9˺!�Ok�;3pĐjCr|%�U�F��w$}`��
���&�:F�Y}U�)9Pg�)�W��XĲ�n�ӊ�իFM��Ы��Is�������M�9��,;K�k������f-��h:��iU����v��ǏS�$��*��"��Ѭ7�������8՛3p<�>[���n�V�!4������ˢ��p�Ÿ��m��s�Y����i�n-.��t�g����y��EW�r�q
-�ss��]�TE
W��� 9�`��M�|�y��zOm	�l�`���79��.j�+8��R\s�:a�pjϜ�v����s9�s�:wn�l�(�\c�W
�9���/�5�F�%���m�:��mۖ=�o��s�^��f��ul���XӮQ���ݛ�ez�aO�ϧ���Β�	d\��rn�,�sE�7�٬Ҏ�ʽ��0!o�^�{Jϴ�=�,�4@�����ЎP�[�U$��?{�b4��^���o2�9$Q<��<8�!6���30ҥ4P@{������Sy��ȧ1�z�ӻ։��ۙ
4�&T���,��-�3��A9J;k�
#]:��E�1����a#1O!I>L��b����0м�Q�+�n�Kkz��9i��<�PR�	�u�l^/�Re�4��f��%8r���}+�V2ޏu�\4����B��o�~�N��7��jr���/��OT�������������=��.��߱�PW3��:�p$j�䶽끖؛Pk��d�J�T��.IP�ڲM�<�����熛l�/�Ɠ�����?���>�4F��c�e�A+]�.К����8����~a��ˑ��0�Yp�{`��re��z������2��s�`[�ny5�D��7n>��r��S��o�JD�A\JHRw�������XiY��������q�v=�}���
kꞫt7�k�F⤄�V�$q(�ϛ�8���m��X�f-u����	���t����&c��כt";�zZ�ii*r97��z6���Z/�[ʄ@��֫n�n�9���{�}:���t��p� ���
�_���B��_�Qa[X~z�����6@�g=yr�:����ݷ�]Ok.�w�Fd/I��3��0`��)'�0�J@�Y�#޽�B�9=28����ƪr��$l�֡�Պ�O.󙎔��|������禤N����ö��q��ؤ�"��y�Ӑ��&#N*Gr���W�ٶ��A{�;��~bo��dz���4�X_t���#df�#�MJ��NMT���Yj��j����+��E�~g�O�r~�㑆�'>!��z��ŏ[�3#m����؜xm�����n�~�>+�~�+ʾ���I��P�f>mX���a
+�
�>x3�8Q��J�G�{g��5/*\<ܻn����V�Wf�Ŏ�F,����iy�T0Wm�첵~{����g�>�س�o��3gK!�>ژ�������hj�!B���N5;Ŭk���_ƴ�/���]e ��f��iuт��~mJ�J+UuS��j"�,��Nm�*�Ԟwg�Z�f�b>��N�f�g$yިg�4� �!�\���^��ʔ[�/Y�E�Hؾ��##q�ۂ4�Ɗu�g��!��g�g���l�/e]{��
:Q��{�~F�.�s�G����:/s�Jf�ث�̠�{Gk)�i�g/�@��#�v���y��A�n_�����L�{=�R�p -P�����n߮�˴R];�f��F�q `b2[�5��J�"���G���C�����Xx�O�  ���U�v����&�Q��s�P�Xck��F�h_�s����\�~�XR����#���K����_�lo��B�0�F��QMQ�H��Xs7U�{/�|�f�Iy1� {j�PJ��!��(��\f�z���c�ټvDO��ʫO?<I��~��s;����-x_n��<�]���z����g�e��s��y�j:��V�����@�j�h9w���)J�3��hhfvgZ�c�%�{(��n_9�y�N��cG�`p�M<� ��f]�5����Y�����%��+�n5����W�f:bES�T�w#\��8 |s�(C%Jݗu�ّ��wF)~�)d����gqf����U�\^�B��q�>�*;}X|���-��#DEp��8��*���:{j$
u�}��vEBq�����b����Ū��`4�C�<�1#����k+�m"mu��~��E%M���B��~�m�Iy��#N���X��:�W]^:��d��g��=n��{�y�G��]�P�w��#bT�êPM�5.���gmY��FJ}�=cuj/���vԶo-�ٲ�+�k,G�7�E�l+ͩ}�&����jU߁�l\�J��b��J4|�i���3��vk۱�ogq_Ks)\��N�@.]	�������>GɡET���`ҝ�wP9��ӳbN�#jP��PdN7��\��i�F�k��rlvϟ�����mX�'�Dݰ��[[I�u�k��ssc��gv�H������g�\#�oD�����[]�Qj@�����.ԏ���#,�=t�sF�9:�ㆍ�Xͫ�@�4Y��?e!V����&�	LB��;V�8SUV������u��7$��]����S�՜i�5�DL!y�U���=iw�*�
�ٯYoO^�(:��Vt�P$�IV2$�)��q!#��ʓ*����W��x�>�n�gZlIf�pЩȳf���j&�vMi�,�aL�l)���g/���t9��29:Y�l�	�#y�ibIMF�R����⵪ծ�N�\�In�ۆ��a��S���#��'fR��n<&����*�Ss�A��2'�����3D�G��3$�r���\��?~,q;F�`���ܮTA*#<���PV��S �S���������"B.5�ݣ+^�D�>�^W0l�ڲ��\	��3������Xy�rY> �y��*�����xzrzZ{8W�<6�X2r�|���c�䮏-(�f�E�p;�D}���OGݽ��S1�0�K��*D���@r���[��I�o]u��,:P�q������ �kq0q��me$iPN��&I�
�E��6���|�Mɿw^�N[�S�����xB5jy®�C�Xof��7I��U�]د.�u}9�d���&ab�.�n�<�R����4f3��z��m*˱֌�5�N����&�x�L��̦y�s����W̼6[h�5c�p�r�a=�ٵ�i�����#�pq��XZluM��L���h������r��sm ���B�Rj.|�����-֭�<7U)v��d��5�Yy.�'jʦsV��)ũt	v]E��4�Kl��©�7A�fϫ)��c��|�<\X����o9�}ΉyE�m��=k7+r��ś��m� �F.�y�R����9��`r̸�r��>�޹��wB|�cE:�Q�����br�.�Bu�YPk�v���ͅ I1w)w.���e��^��.D)�<�E|\��]�#�a��ܹ���ɻ$띲^�:T���,v>�=*���vV���]>��T�j�v]�����Ch[��z���q�)�j�%�801k���N��ݚ�����N��m��*������|���J.�o|��O��޾��@{
K��fiT����[���ɿ�y�d��K"n��0ub�: �M!	/��
�E�-�=��O���p��s+��2�m�vb��B9��EJ�F����΂���N˷�k-r]��W��Sq�pn��6��.��]��f����yvLL��ͷ97�m���n.d�[�ٍ%��8˫�ݠU���,��oR�ll��	㧺���j۴+9��ks�랽�r����/aź�q�t�l�	�l��.٘ڞ�_g�;���m�yn���t���W���;�Lk���\��&
�wch�q�-�}�6�^���6���NO۷띞�"����+���:�jiB�CB
7Tq$���
��&{E�p��vkBk�4����@J�ۇhS���.u�i0��lcP�Z�TR�d{{{<���^�y<m�ʥ]�ݍ�fzn6 ̢h���>뵩v:�[�����m���y�z��r,���\'ێ#���:���1���.'�X	<��
/\���Mڗ`g^�q� �\�� ݝ� v�u7V�v��r��/i��82X��n�tg����[�O.�1��1���b���ͮv�=n����猡���.�޲�e��nLv.5�Y�3�:��ǌ��wf����;צzrv���>��:�̼#�L-u���;η<�#ɶ�r�t��S��1ˑ�X��U�l-<q����p�T��1�؛y�q��[X1�v��')cz�nbդ�]w\,pl��=햋E��l�&��41�Y�ٜvS�&�O:C9sūw2�k<��q�`�7��808�v8}��)�NѮ��� ��{r��Nw8�;vh�v�ݩyK��n`�݇�n2glJ���í��t�u�p�{��A=�3�u�ush3���2��6�.\G����xj���c�0Fsqryμ�ӝ���vu\��0�i�c���v�"sE��N��F���W��+@K�s�Bu��e�S��y-�Y��v��cuiO]U��fwk���wV��=�N������6A����gn78q�m�T�N]J�P�[��;,��u�q	����6y�e��`�y�t�i^
�
SF�չ]p��9{cC����g�j�cpBZM{i�.�mø��3ܰ����9.�w�ol	����E���y��f)l���`M��6��y[�j������+�W���k^Qi�� H���q\����;�8s�[���ܘ�;v$�^z�D���ͺ��O��uZ��hWf�sһd���B���;Wch�ڢY�"$S� Ze�`Q�D�U�1�s�TE��]�Ub��@�'ȣ�3nx��z)ͺ�6�����}Sށ��-�����]��&x�${``=*�0x2ap�p�"����ɂ�z�^U3�ہa@���ؼ�Qbx�����g��UG�b#�36��sD
�^�����!;cH�����|�h��*�(�(�6�iv���YI����5�E�"�?>�A�X$<��W}*C8� �)2Ϟ�9�V�v�:*�{�2Sh�
�sw���{�b�3�}�:�6��;�L��ܟ������*��]P�u��=B
��Z�v�n�W�����q�$����j%�ṾD����"�P%����Ԧ��(��ƪ�������X4��2�	-d��|�3+Ƭ�A��Sc��uO��yױ8w$W��7��c�<����=kTE&�4B���uh���kn��A�ѸN:�\�3�m7d�XT�U]d�;������,��^�R���7�S�e�ay������i�S=����k������\4������]w�_m���,�E�a^`>z��*��G-[[	��?U_��}���x�Kk�q��5�eɛ�����y�m��zk�]Ҁ֞�FA���L��6�en%�6KÛ:�j6%��;��5�s�P�9�.�ʬ�p���Ⱥ
�{��z��!�n��B�#[{�;�j���Q�}Rvn�1�BI�#Go|�U"���j����[э��TF�����-�1tP��{x/'C��y��|���8�$����qY�}����A�	9&��b(�^Mc��}��l�QtB�g���m��q�ܪ1ۤ� ���#�w1/�1$�D��tٍ�ˋ�֩U����J��̿�q0�j�[\@�a���(��z⁜V[�&RJ����������B�,��Ф�k�q@��f1G�uE�o:�B5V��TX��6��\�Ě)8�&룚v�;NF��t����ᑧ�ͻ\1�A���%YI�����!H9#H�Q��ĝ��&E���1
#Jۮ�n�)�̑7PVs�8�9!�˪����I��P��|j�l��V���+yo�!�1�T�4�r�A�=S=~��N��#��e��E�X�F����
�t�o͔`�O��M@��:\z=yu뚾3�Hk�T�]V���iGm>�7�5�K���h�#�ڇ�@���r��VF���j<�!�ՙ��!W�e���:�'��oga��o%��i`��z*K˺w�Sū��O�-A�0ݣN�Q�F�m8�,�1�1��&�ķ�q�a�����ޓ��#�WX�q��?:{3��,{�"�FS8��#�#RѨ'#���p6�&�h#A��d3��W��2ah��a����K=u�6�����}5��M������4���yR��*��b[=��-}R�ezW�[�ȅj�iz�l�?��J��i�pű����-��&A��=Fw�[������\2�䨇'w�緙����ܕ��4�TJ�t����h2���k��n4�х���9���Nms�!�J��,�x>��T҆��}����ABn550��T��`V\����Du�Z�uAlk�Ka��<L�أ$C��B5wj���ڭ�1�$L2J��r�����nH'F�}�B��6{�i/9�a2's�yV+���'z��Ό��B^�>����3�f���t�����h��1�\1،�"���[�N�.x�n[�bY�+/l���[�]��uj��Ӿ�C����\��U���2oNP��hK��dIR(�-m�����g�n��%ּ��tk�h�I��Ҵ'y��P������2B�Wuw%GPV2�t�g��q�=�u��z����޻����|#�̩}|�m;��;��;��fiRes�^�h�[j�+#z��V�����zWAG�󪬴2|�$F��M��Q��y�4}�=�"�5s�ꤏ�z�=�+v��8}�T�Ϛ��>�D��k�Du�DjZ�sÒ�@��3�_�~�4��Z��T�U�+%S�Ƙٻ,�7���Ǝb�"
��䀣q̒���%!,��|H�������ߢꖆ�!�e���ąY$+o��iw�=]ᕌ6�1��2�dد�L�n�i{�]�̯�s��B9��H2��ڌ�]�h,���Fn�.8n!�i7.��x�=y0˷�D��>�A���3�\�ݹcZ��p����J�M<d(��8"n�S����$��3��>æ�����,��΍��MmM��*�3��PIwK�$:��j����'���˅df�8�p(�����{u���^�Eo�	��W^W夅U$ة��l��l���Ϭ�uzۺw[�G�Ɂ��|�_'Wzp��Kzf�qbh��DBƶ��F�)h��E�A����8ĺ��t
�40����2z&�|Z�c|s�+��cY'��^4>�P�B�#O5���Q;�l�j����j�{vzjZ�!:5�pݮ)ܑa8to�3�e�ط��Z2�UU�g/���Q��Sw�hk�w����J�N~}ߙ7���+-��y
'���MZ@��hαn=�Ǯ�Y��9,f�x�[]��UD���֬*s��t�9�68�N���۷g����[�mvŻ������%�<��n��:F�{c7W��9��@p6�V��Ձ���9w�G�Nv^��b�\	c>(���km��J	�;j�1B�؅M�l�T<�ּv�[�zX74�먅����m�85{U�48uQ/����g�ӈ�0t��y-�O#J9ζn�a�9��\�'A�[������������{��5'&�m�񝳐Ϩ����������/�Pf>�D�U��N�d˳�P�4�E}����VEc�T[V�Rev�g�yV��-+U�7u��*�����dl�������(�ș�^�s0�~F8�sʨH댹��-���bY�۔��ӭ���!"&�.C�=A�٣5�1[f�y���P`�1�-���")jI��]�Y>���y2�}<�ԫ�	iU�cJ��RZ�k1�9�6�H6�E6��������U���aU[F`�a�P�2�3�����^��5H��|�o<��:w��ۿ�HVp���@�pbF@��Ju��,�q@�.CTo���Ry�z��6i�S;7v���T1�9]Mhh�W I��@.�bDvFk�(t�Y�9�G�Q�9�q�H��σ�Tܼ�ͲTa�b�J�ݱt����]Y�j�5����Ndt�l�<i�AԨ�"nX�������H8Yܘ��M���U��)�w��SQ
-�z��W�~�У��f����ZV��,r0�Vj�J�p�uIDJ�SnW���ܝ���,me�)<��71�#���9%y�wS�{z���;�zj>��0��iTNҝ4��Md��U���1;v�ևhm�o�^e�Fg����B#A��Lo]X��뗬K�;��Kj�rp�&I<9�H��C���y2u�Hנ�=ZT�"���R��X�6�<ˈ��F�����+GY�uI
5��,����{��iS�M�V�?J�HW�M�"�a��0RM1ȉ�;����Ĭ�,�� g�[=���["=�~ta�u��E�.��(�^���swA���F҂`q8�H{UR
�ח�����*ݫ39��@l`{�69��m���AT/�����"�/,���$�;�7t8�9��>�Cz��e�`?Hˉ�|Z�B��p���^�ˋ��m��-d�y[O�ز�k'a[�x��"<0��K�ש�fӬ kL�Ѭ�{�׆N��!�_/J�`��w#���}%sr�p��A������+hV*�#�q��*��Xt�<g�������}!���n���M.�=��O����3巃�Efӯ[�z&cWod�V"�@��#N,����1�:p�
�oE1>���rv�ٕ�yPTYυ���c��}�0E�t�'K��ή���Цu;u!��6�S��Kzk�q]�<�tB���[XX=Ζgm8���C�v"�k���I�E��_�,o��+���*�7�$�%BBp5$�=(��-}F�B&K��j��[�k���z��!Q<�@��0��xhCھ�K#q�~jL�?�Dr{N�.�m���/�m��CA��� IH�H!�VE=��7�pD[�}����/�ٛv!����3k�Gv��./����v^�_a�ǻ���H���7���cg�8����J
��4a���5�9��	�)+�[�q�թ�7C���Ty����;�z����ɘS�^�sH�ݓ�}�"b��b�e��#��\pd�x����Ȓd,��y�����t;��q������n �%$5Y���y<�Ewy�E�Sg\FY}�h�Nf���:�����;Q��d�a���lFYA.7���ņ�`��fk*�lc��9��n���YBRTYVw�]�?y�m�(Q�1*�7���lp�.Lǻ�,�2ed��8MgD�BH�s�b�V�:"��v[@.��XgD�>�a	�1θ���K%�ݳwoBz}��{�F��pK��V���1���B�O*\�՟=!��c��vy�����᫻��vh�X0�.gL�d-�v��沘�ug6�+��CHXϺ���-Y�X����Zo�V�<G��y~�\����^�(��"nc�ti �T�W3����KV�m�}���_oԪ����R)=~t!Ca?!-,��f�ʏ])̉�$U�͸���f�"��۶�r�^�n�Bё#��Q�Hp�r�h�6��8m��meg��u�c����ay-O�y�X����5j����b��prP�%c���]�}WRQ}4�[���|�#��ңqƕ��Fw���N_߽�8 �����n�U� �^Hm%���^�8IC;��3��0*5Q��庣�U��W<fRY�+�"�d�^��7i�ӵYb�AÏ ��Q!�0d��I�5�n&@���#e��ׇ}�=)�2�4�s����NK��\XkW�]y�W$�C�����r�$�U�َ�g{�m<4�i"q�}��aWAy�S_+���Z��E�\�����{��D�j�9���g*mT� �㧦���/��9�'w�qaK��g"	�g��-vTԤtn�qFZU�:��E�Ǳ��V|�8���qP�S�d�y#1T�#���w�����{�3���;�L��WX(R�Ae�2Xׅ��6]<�=��P�/݋R5hY�� kP�bi�!+8�%�H*�� �}Ϭ�:oV��Wٻ-Wk/pS�y�m��+����'cQ��4VI�=�nۃ�/5DE��q�n������.�1��=7!��^]���7�:ѴC<j�:8��+�zw9t��I��K��mňz�k���gm��P#��u�1�����qg��[�DŬ�Ѩ8�#n�c��6z�2��k�s�3��2��h=��٭��H!�sv�s���y�O6KKq�ür��t;d�y��ΑzY��c�&�N��֢
q�q� ��9#�^�ancK�fڳO���Q5	n�<ԓ��n?6���h%�����������BE�ƕ�M�6j��gVH�]�e�W�$J����Ȣ"D6�i�MG7� ��A�p���˨, E�A;�r�;��x��D�-$I�g*����D�4fԹ�B�z��rW��Q�B=���=ǫ��oM6�~��̕b��^��1#i�Z�Ь�z��p��f`���Qw�m&��1K��Їy�˕�����^�<�Ć���{����)5`����&O �� �.2B�3��S_���;}e	=�aң-h�|.�V�&G���a]e)HL���2�ʝ�'�;o�2��1��2�FeF�8���e��B��աG���2�%+��jH(Y~�m�<���yJ��]
�Ch�Ω/���|���^6�ꆫ�[ĽFe�L'6c;��SAhp�������s6�Bt~�=U%jj�tT7h�y��vp�8s�F�qU�c�[s�S����I�َ� C	&�͐V�o���c��q�M�jYy�JCl���d�%j��ȭ�Z�F7�Nٹg��s7khY�5�}yb��,+)���IREW�wGB��U�Ckfq�xvnT�������\��@h�׽:]�J��+j�n�Z�ɴ%9P��������9���N��J����i���
�g�k�zK��/���[�L���.�{��ﳃ�R��`'���<7&��y���~a+�mӚC"	D"�6ۄ���5���U�ͅ���A5\�b��Ƿ��I[k��ˀ�UC��Į���	�z#u��$�Ԣw��2F�#��������rn�Tg%���wѝ)�tvTN��'��
Wɖ������`��#�B���*���؉�5"/�i�aD&[o)�w)*\�I|�+�6(�ղ�=#V��.aH�^��kӝ��'�����y�4v��Pg���U��#-���_�um���۴�c5�L�T�a�
�q�b�<5��:��'i�`˽u^�vV{9޺
�R�7;̱�-h�ضH�u���%�ښ/��W*z��rg9��h���$��s�f�#2UEѼ̄����[0H�QIqẓE�S̽g}���s��X�<���ql��uZ4��]����~=�r�S��ж�S^���\�;���~q�gs Ȍ-Z���{�+��Tt�=ohl[���}�җ���Y���=6��{��0H��u�YʖT��i��*�BM�s���f��7&��꿤;����R)G�L%b�y�r3K���J��'X��/s"��6����T븗V��@�y�2�yu���v[S�M�I�x���BJ��p��܇-݉Ҷu�2SH<��a#R�N���LL��e�Z�87�s9	��F9�n�6*"�+F�h�}T�z1���
���C�h�H$���t)�6�
Yս��mh����̵�g]#�\p�e���ռ:hTVi���E����w=��f�q��{*��N{�i�4�w����ttr������gP��W2�(�#��[V�MV�h�oOSf��G8+�]���9�BYV�5�x+�]�e&���+L�7��;��F����|E��ݜGp��s��X�����œs� v��+��KJNvu3�#�xS&�C\WV���YF��I7�ϻe���Ȭe�����\�U*N;��'(c�<�D#�r/Q��Qx&l��LTn}�7x��/��d4ۛ����"]㲓�wmi7�7����n�p���cu�7\�����W�#ܴ�n��\s����'�L�
�n���/*��5�T��EY���`!�3r�}�k��p|D��^
x�+]л�S�;w�!��ymϏY�����y��U�o�L79����'�maݩu�JY�^���\��%�����N}�pAa����=����x��D5�U,��;z��yǬZײ��|�`}]���>u[x�-�&D$ �vX2�c��ss2��B��9MP�m�[)���fy%h"�]�1V�J[Ǿ�u�Hv�����#���fl�]�2����B�.8g2��*
E�um�'�ѧb_,��)1J3#1�����fy�i�s��P��H�r��)<a��]��֤�j���ɾ%;��>�W6E�_>xnu����"�ݾ>�5�wГD$�`�u:����:�m�a�sWrC�u�����Z8[u nH�
8rW���){ȫ�<sso�k���0@����]:���!e���ά�q����{sj������A3������� �?ԕ�dn"�mt�^4l��;^�~䯴?}�^z�]"�ø�����k�Jǻ�oi͢�ʮS�/R�D���r�d
���7 E��8d����u2�9{<k�L����f>�q\�:����H���jsi=�Vkȃj�J�/�y�(u�;�ܖ�U��@���F9�BJp�d�h�[ej�@w���s��hԬ"�+c�K�ӈǲ�������HsE�Y�
�_��q�nm��B�;�M�{�=O�����=���-�mC�X�2�׵\NȰUئ���w3"7~_W~�n��f�'/g���)s�7q���v��W��J� ߘ�S�$��H�ԛ�V�)��"��u�ʳR!�ә.��"��"!K|Փ�]���9�rZwy�O�$Ӂ����
�YIuy��.�o�n��Yx�����]l�dІ�=��g�I�p��L��
hf�W�Jo��h5���Lڊhx�ʷ���Y��q����D۳[7��O.��&
�JVM���`��d����j��.����5�w�U��=9Ì�WF��/ݢÛTc�*�=�^��p���̩�K�)wM����La͹6pP��
"�(�E��2�n_����ay^c7Q�gk�.�z|k{�j�Y;��o{Ǻ��N�q{n�+��#Hm9�}0��h�٧&~��;��܍��Aڇ-3��;}�M幷q����&6g��R�[E�,��=����k8���@v?d9���5�-U���4�	��P8��w6
�Z1�?;��v%�ZX۾���\:/3v�nJ��U`4�5y���7�x?!H��2@�wY}�@��wp�S��w*?a؀w��`�q�G���:�CaY��3l�]�8�X{�m�Ȼ��!�:�e���;ϻ��}ϫEUr�;d�-�cY����Q�������]�g�1κ	zSv#E9��+�KoV[6�w�K��7�^�:\"�>ĽUN�[�g��_!\L�nN�;��#s-�S�{�Zn
�����������{;�c ���j��z5��p����`�8��Ѹ�:� Sc �����.a�t�l�N�\g�l�k��=�]�ܝg����8|[���#[/[=�d��b�ո�z�����q�l�s�9���ω-��Z����f�JmѠ��6��dQ$罢4�{��7�o�}�2�I+��]����fMq�&oudlScp��%��لH�79��B)Y�GϏ!�T2&�VL�9�\�؞�O^�N�pw��{1ޮ�|+̏5�1�����m\⡳��D��s˞@��=�lo0z���V��;#(4x$j%9)����#t2���yo�}��U�c�����yFE��6E3�y~��I��O=mR�HZ]KnDd�;V�y���(8n{����p�^ FK��N�}yy���m���^6�;�c3/Z��@�9ޮ����&wW���?*�*j��x7ކa�M&p������>h=�מ��8�������ց�v�J�˥�W*C	˳K�K�y�g���]����=,�ݜ�~)�7LN�]�L�bV=�Y��pd1�3[F�۩p���4���m*fݮM�g�Y��W#pU�(N����d���Ԭ�����X�*@����W��M�X\�����4�&�|c���e���W�{jN�_B�\�=�#��j�0�M�\7XE7-���ݹ*�kLԽ,����|��M$�y��>��t����[��_c#~,̗ǧfc/upduf��Q8l�,�b�}]su���gH�	M�sv�e�ԙ�=T�O�c!����+�K��[�slLwB�a�,j'ыC��6��E�qXz�g�k�`οB��*!e	����������ۘ)�Ӆ�v��?Q{w������QM�q��	�w�qu��_�������Q���|W����2nj.�ݹ��]ᠯud�T�'w��v���vem�O�nJ5k�
ЃG��8�F��]�dj�>r=Io���
���u���1}i�&�Mgua����5yW��=�W��H.��x��W&sdf'F>Nk�z3��{tsøG8:��A�p�wwE�O�k�-���6��O�~'�����զz����D\�@���j;m@��N�;^�b�/W<ZB^���]m��vev��)��5���%>s䄆Fᪿ�<�n��ߕB���3T����q�a#��M�l�sQBm�Q���㙺���o6�ۭ%n��)�J����*8v��,Lcz�	�f�o_�
v�WI�����ZZL��s�U�~s��ҭe�N�&!�&�B�
<��-�*T��c�I*S\y[u�Ήؙ��P�u��_u����wH���zEr��h�0�4	�Iܟ=��\w3RU��4Tj0J��7n7G��2'�x�skR��`Q�0[��{�=��e��1W�-,Oؽ�.����x����l�u�O�I(.��M����sxa��a�p�9U�&�qu�8�<|� ���X�V�>pc�u\_FG�/A�!�*9�Tj!�SԱwd�f��g*{s�m��r�@� ,�=U���Ȇ�s˶Ը���DSZ�q6��[�@s#��BeC;IJPQم���Mx���l]�~ŗ�+R�ޭ�]�� D�[0�H��9I�۫�9mq�����}~�*ZN"�E����D���h���K/�C��{���Y4��:��������DTMn�i<r��q屸��ڝ�x�8��e.�����nUvb&�em��q��d!F�%Gxn�2�I�y��^"dnoG�{ٽS}�]�z8J�KY���vw��¯�%^ˇ�����K�.-�o'6�hgv��	6�i�le��_�w�;�����9�ܨ:�6�r^��d��Nm��*
&x|+ݡEol@�U��cDo@4�����)��+9xi��9���׬;��H�f��=��]�Özq���Z�kQK'�GSb�Fzf���=�Ѕ��D2w{Y��Ҕ7u���蕲"-�LvfJGycy7�E�M�8tT�sٜ����X<�::յ�$wN(�l�yT��X���g��Ť�:�f8�"+����>�g�.�x�8�)�S��Gf�<��~?y�������+���b��nJvB�DQW9�zNe�#Ҽҳ�S$�Гi�x������B�U�r*��2k����E'AA@����!�͚�S~�;�yT#I"��œ4�ߧ�ww�O�&&�tk���t��Ӽ�n�k|�Û��)+<	���$Si��-��f����,P�n��ּ���XfN�� �e�l?n�����xJ��K���6��]E����A\ڲ+��(�!E8�p�a#��?P�fV ͗Gڏ�x)y5`nČ��.��'X��Gx�.�͋���Ψd(.����:�M��F�촎xn�u]�PJ^�Aq�#fH�휵;|�Y�~׳�����������C[��詳�v-Y;fJ��fP�|}u���tK:���ҸO2l�>�5s�\�Z/��34���ǵy���l8a�q���w��扦�_��D��Z��Ә��#�bx�g��h&���y��GX��ۓ��Pއ��#�� h�uظv<gk��RA������Z�Wr�\i��[r%��ɍ�1�oF]v8����{�n�L0Y�oc[s�]Y�K*�-n����3;v���ϷnƗ�Q�N.���6�w<���N���Q�6�J��)"i�h� ����l��śga�v�a(Up-��{�뵶l�m�nx��֜[p��$NͶ�>;n���Qţ�ҁf'j^�Hש*�;��]	�-�=ب�]��^�W}����u�W����o[�����2�,ՠ�{��=OA�r���r�����OU���5�.�p)!Q% P�䍫�\m�����F�5���S���d���#��d�����<:"wdy[��j�I�2VdՃ���y-�Tx�,� ���d n����{��E{B=)6ݓ���ШF써�X�qvy-���{5��/�N����5��S�8��,R�U<<��q@��)�)޺�U���l���J�{d��ق����1������z�x�� �A��`����q�(���[�9��w]�$%bx���[��d2Dс)��֪�K�[��~M�N<1��/WIΝ׹���B7%����P^p˄T�.���ݴ��e�`wZ��-��=��eH����J�<Y3�w)ԯ^q=i�ur�s�zL�F[��������9dk�7y�8zh�����T}�hZ�ű��{BÕ4u���[��C~�J`ʪ�[|�V���S��H@�*Ez��Qw��\�}�r��F�K>�߱�+1oQqP�F|�z�m{�Nwy+~︾"�s��73j�㷩Gq��5�/�I6W+�W�9�-�g�;�E��b�+J��!�/cg�9��ҹ(�׶�x�:���aѸn�� �oV����		��TECM�ۊ��:!��F��zeQ����iU��Ɇ(�w[��cf��9������l�P���ݚ��R#�ߖ%X#)b���;,����C�Y��O(N��#�m�����V.n����bپ�A�U�����ǰns}I�<�l>��0�n�c"r��	q ���e[e]����ɬʍ��vƃzK ��^Pz�a�nL �d|��4k��H�<e�}*}C}�=VN6�;����do�TuG]�ʠy����	��׆�����h�V+�Z���{iyy��`9��Ӗ�j{;:v��/�9^�1㒞&��~��Hv�e�2��+�eoYa����)��͖�^��,]�� �qб��=S<���u���\-�<S��c�5�A��ܞ*/Y�WYz=�:�B�٨���7�)�=y{z���7օ����C0&�>��!��ۢ��_���J�w�񛕘�#��wI5�wm�\�Ӣ��sp�=��(��XK�+��g�o�<jW��{ku<�f>j>�#E��1��"ȣh鯔��E��]�h�s�v0��"�R�y�J��v�����˱b�*N[�����W7��,(�E8���&.��J�Z�r9�G�燼Ĺ�+^J�:�Qb��k^��V{�sV (��1d�O-�*x B<)4m��ʅ���4�7垪�^pX�3���5yeޡ��+GtuŽ���T�D�p���u�v�ď��R�����U��33�9k���W��ɷ���2����>�xj��������eyu`�y�8�eH#�I4iM��}�푻Υ\~�¼��z��^l Y3��ói���|�2�ߗ�'q%SϵDe��>�0&<�	I6v�s
w��FmGx�}�g��+�m>��ۛ�.�|<���`p��~�}��#3Nߵ��fB�10b�F"� MF�j�w��jLf���-Qb�jN��svl\��Z��(s��f'mn+�z���7[6#ʪ�ਜ+Фq@�.Q�DL'$vǟ�`5!��ؐ��¶�L�.x�ɑ'�%U�>H�"����)��g1>yo�+���~�-��av�.�[h1����ר�O֑WGdq�ÁuJ�y��:�4�,=Tqb�}ț����t�;Y��۱[�G�UKbp�,�o~`� n��!Tp��l�yG��85sbY�������`�����8@��<:�`�4>�]��r9�\(
�}�	�~�Yg❺�J�\u�,SM�����ƅؓ8�Nv�+*�9�'�g� �n��S�k��Ś�&���A����d���df瀅g��w]sC-�L�lI�z��vmh��P{�{c����� ��7��C�F��%e�+��� ������ɷζ�N����d��h�I�2��vF����kw�PE��[�Sapv;N�Ӈ����WaBR9Np���)��<v��S�CG]�?)S�'��� ���j���X}S�Mō>��*��rQf�3��	����㉸�ːd�8ó�n�������CE�̻+/���՚�m=���z�d����R멲��ml��"}^����i�Ims~�6�1
���:�s2�P�O^t6'1dӓ4�c��r�/�8�8總J�5׶�(�7@�:s3�΃.re����_p~�Ie#�f��� �γ7������npp�ͥW���H_dT�3|:m�yػ�X�J��h[ھ�i8^�b6!�Vff��٢���F#�i���f��j}�2�hp�O�Yb�h&�;�w��v�[9�%�f��U$3-��8�M��-�����A���	_����0�׻F�++iҫ�;Y��[��$5kޒ�w6�Ȏȵ�T���ʚ��'ȧ�df<1�Ю�2��D�Y%���ٸU�s�uɭ.oM�֠͌��ޤ��S�ocR+�t&#7��\��"�"��:���	�Դ�=��Jvzz&�u�
��|�Km1�Q��uG��+zo2SݛUB��Ȥ.��f��X4�}��{� �*�d���VD�=q#ڹ/�(R��v�x(V�,�iȝ,w��甌��v�\�Ѵ�9���a�gkj��2�� �{*֦4Ѹ�B]N���mV,���ź_�DQ��X���޺;e����� 紋H��e��e��r����enm���/i�qoHq�6�^�yծ�B�5O�3�S)���Z#3�]���h��Ep�$��s'F���
X�༊�w+YS;��O綖�9�x���
�-��3���u�F�./����]uɺ7G��&&��]��T[݆�)D�ӵ�lI/x�X���F�z/5�uHArj���8W�BE�q��9a��-��,��R�m�~%\:./�(1�޳Ǖ�G&5��#��[�ZR���z�����-Pа{������bF����3s�-�S�[6�S��S����!�ԫJ��]�=k��V���㭀lm���i�����^Sp1���!�����0\<���m1�[�obl��h�5�d3n�'Hn;>9�(t��`�']!�m�wc�!�)G���K��6�Jnԝ��WM�m��n��D��z웂�;f����m�M����s��3v��[��.�Wω7�6�vw=Ma�7P�{'�����V��9I�����vФ4c��;�!\��	�8�ń��v���HɎ^z袷e�2ϊ���Q��[v��1�6��sx{0mj�b�j�ܥ׳k��fޝ�1�nG��c�"�l��:W����f;K�-�w4m˵��Q��<�{X��®�+g�=^���7bύs�6�,>��s`��Al�t ��R襵ʁ�Iöϗt\k�ۊ�B���wW�RԻ�!˞����Ah�u=��vdKn�W��f�m�:S�ψ ȧWl���U�ݭ���t�ݸpn�N"E��t�e;*�"=Ep⮷h�.����n�+���C��-c���xۍr�gA�(�v���%�u�秥ܽ�]��5��uێ�s�q؎�m�^v�ڣ���퇡Jg'&s����޲p\�jG=���.y��m���]x�yݺq.����Ƹ�q�m���v3�N�q�>n7�n���y.3��+�:��Œ��ێH��n�Y���^8Zx{sX�����E��N�\<����vdV�ʜ�y3Y^B7Q��ܕ�'@�F91��[Ý��N�8�*�s�DG[ܝ�G<��e��f3��I�8N�l�P�F��s��v�Ó�/e��E��v/G9�=��U�7E�n����B˙�ۜm'n��a�x��Rj(��Y��۫�����z������\Z�pqw<YJ�ب0�Db�"�!�1�ݎ|`�����ګ�o�{%���7���L,)v��ˮ��ƫ�t��n�7 ��
�}�z�s���'l��>L�� � +Uf�2�m]�F]۝n�6����s�����wR\t�8|g�����5c�y�$�;��Y�N��u��vm��u�Z�:vnJ��{m/ts�[u�8˙6�u�\18�U��n^x��ٺ�G���ɴ]���d8�2T��'�S�Pnf�g��>���/�x����a��=�����*��Z�c��;'Cs��@����n�@��;]7����d0#�[h��*۱Y�ط�ݚ�l�W6��-�sНYݪ���P9j(��|zH��v=��fl0L:U�b�U�r�7Y����Γ���k�(��늦B�D��]������HH�|�pB�0���"~�Z��3{egha�i֬����[�I=)ӛT�|֧��n^=/h��#�w�����L��x#v���p�4�"ʑ׶�(�S�-�&�n�=}�+w�T��ז$� ���]ݢ�+�]�^�w�Z$E�ux�x3j�b_]e�aƹ4�i0�-؜*�:��kh�����5��4�y�K+*��`�$:�i�	Ӥ���������-=�������`�0�1��k*����QDm�\)H�ө���#&w���+��gt�{e�Z��c�H�-@��[|�*���~׻�f\��i�� ��K������6"��#LDw'WkX������rl��/!�6g��3ڐ�����������uY+?.��k��,��l:mrٌ�ckC3���Rʦ���m:�l��y����a�{�����A��%�$bEI�ᵕ�2�s^m�Z�Cn�'1W�Pu�XK4#�bޫ{�����־�cz[y7�p�.�Қ�� c�<�hVqu�l��s}xm�R�2I��kxV���ƶ���l�֒��9��y��pU�=��r��%JKv�h}�,����Ѫ�#~ �~�XNv��Ρް�M�x9-�r��1�9�[�����<�Ź�ieh@�4��*�nn����J���H4��c����5�oҭ�\�u��u�p���oX�mF%�Lt���#�L�{xٱRd=�<�0���>�T��6��y������'�=�ڎ*K��Y�X��jmx<&Ի�4�]�0�Ӑ��#�$��{�]�-9�}��<���q��L�%Q:�#Di�;�jD�]��X�,�g���x�;Y-�uey��V�k���vB�R��ʍ3�<����WejS�^�ܜ<hA��񕈕JI�y=�h����=w���Eي`p��1��m좥uY��_��syr�\6�;���N,R��l��{�uHv�Cj�z�H)��kt��Ø��_��)>� �h�	R5c  ����c�*��a����7�殤D#��7�
��׽�}���'o��2��"��C��=m�8��]��u���^�*�ofep�/Y����������Gϵ�c�7�喲?I2��]$z6pp��߾�C -��n-��tl��u탵iiV��)�l�<�T[r�{����EA�}.��1x�ʎ�}���{;ӟ���+�v��+$^�X�B�D܎H�o�HVC7��V�C�����bT�#�x����vSx's�{<�;�`gu��xjZ�����c�L���������3�ۀW0ND�y�L��z�KH�
�yӛ������a�y�n;��������s��҇a��xa�1��,��vrVQ��H7����v}��R��H0�&G*E7$�,=�N�*�;��s��^�|��jm�	�2j����}������>�Hn�1��"��S��6�M�d��t���b��
q�^�A�ק�:��^��p���ȕ��Oh'S�*��v�E��[�3��P$��
�v�>�N�������W��0�]Z�?_��Eՙ'�2#�g����f1�ԕ����	�o_�ڭ��0�t[���Y�}o	�����;w����)=X¥9�v֍�1|����YuQjP�Nԅ�[cTѷ��X""."��:�l㲖���qPZ;�����؉��撽&<�n
E@I�W�܇{3]ӥ�qAj̳��us��4G�9^I���ZE/R�9fzםy��7@_����߾�i)�X�rV#��M�.v��+��Qn:�Gl띧7�lM�8��F��5�<��MgN�5� MzF�v�(	��w7^W�S3U��H�r����),�NgKٓ]U`��Y��}�G`4�p��)r�0����������TZ�M;+Z��\��d&�Z�}"e(^ypOVf{5V�Oi�vU܃�J}IOw����<C���a��j) ��]�]I��T�������#����2����a�XA�k�ԕ,{���m/S6x�{�ݑ�PN���X�\�"%4��P��7WGt�5�]®�5�>r�Zd�.��N��
y�����u[�0�\�\ �:�*�g}�]�f��KA����孋�B	��M��"ܒ��@�ު�WwCw`���9����Lұ�/w��
��(�<�O�E��f��xx�d�Ʈ>�٬U��ޖo�h�ȍ&�uP�<�&�!�z��?պړ9t3*.����6�*�`�mE��=D��-o#��w�3;�~�2I�G�WCv�����Gk�D6�/<s��9����X���[���x'I���'�����F}o8�M�V�n�b��{Uv��h'p�7%u�j��enx8�;.�c����gU=���Wcn��z�[sm� T�m_7����2t,�� �v`>�n^���N�my�-�ƩE;n��6j���Q� 烧�y����X5�ˡ��3ݷ	^{N�t��u�&4kc���V�=g���/���j�:�"v脰�Z���MS'���ն���Qƶ��O�=��C�����Д/#���Ml��-	l r���QuM�
o��X����ak���� �RC����蘻'��/j�w�703�!x-	�Ԡ�=�+����o(�VѮ�3��{��.W��v��=C3���V.��5�M84r��J4�}��n��V*eb�/�-�4���c�>x����x��������OҚ�6�V�y��Ir4E���Dx��ɸ�s����3�S!�.D^�7�s\�R��2�u�rP��е%����jT^�Frz�
>ˍƠ��rH��f�^ʻ���Y�E�f��3�q��u��3tOVXF�.^�V�
ξ�{��ÔP<���z��"��z1�5��u=n<��]���èT묎'�Kv�gU�6�1ʖ�dJ����۟3����R�;�+R�_Xs�jnE.�I�
����52�o��y,
Ϻ���[Z-�O�]c��X27��p)r��g+3��z����g\JW��*��E�ޣԠ��&��/S:ƾ��č*[�U��#�WA��*i/`ɖ���H=�;*E*�'r�ފ��dWAγ�\wkl��O����Ĉ��f;�D��[�sL���A%ς/��$ۉ��3�Ls+g�N\`i���z]�/is��2�?[���v����x�s�GNM���u�{j?(�>yjV$�y�k}�rHl@�JB�u�҃��M�������jU<Ǟ��29 �׭z���<��4��d�����݈(s
{�t�>>��3�j۲oӻ�$cdl$Ą��*&5Z�������X.
��ql�o�>~��K�Ȩ_�{�\��xT��?�Ww�Û�66��F�����طAe�Gud�z�\�l���,��q�i�UtT�
�\���e�;�[H{�i%z�����Y(��hVd���7<���Ǔ���91��zP-�Uνy�!�c(vq^&6�*"�P� t,���-S���Zk/0sk�����j`WZ}����'_�=9�QW��)�	\���A^�Ֆ�mQWcs��X�R�QQ���Q��۠\X����L��){z�N����匙�Eu�l��x���b����X�:5t����]G5[�X���dZ��}���5o^�E��/k�e�>��:l�W�����3jȮ�p׿~��M󽶋�M��8�E%M��M��2��c���'E��aӽB�M�n�Kv�2�8�B�1������Fʖ�~�K�*Yn�P��<�)H�DH�%H{9�5
uTW�įVӵ*Q^Xj �iYg՚ ��d�����;;͚�Z��w^9l���xE�k��r6I��1�YH7�vP�A!`��3�+o#;�u��n��n-�8v��$�G!�%���ԙJxל�۹Z^ZX��x�b�-h��z�?����)���[܉W5�'�'��Yu�)?2�1��Rۇیq�ܨT�.i��}���9^w�{'��H���@�Ɍ[]���L���U�!���a�:4�q���̝���q	95���֬{^b�w/B<��㺐���f�#���>�}9��*f�Fnw��J:j�]^�/E��d�#�*��]Ý�{��Y��wU�x���lW%������w\&���g����z��9�8D�����K�wA�=�z�p��0��p�X���)z��w���z w�h��mv�`v[ů��Ӿ�����^�f8
m&r8Ds|Q���������%����^���3��f���p��}sr������z��u1�>��hy&�[t�PT��l�h����</&3d^�����:�V��@�IHAf"��'�ﭶ�ggy){�-�4���y������x�g�ed�}"�r+"nI*r�sU�>�F�⳯����YlAI�$n8��=�E	�=j��"+�e96u?�j��Et�1�XX�k�YU�	�F�����[�#J�LE!iI�+QNt5���%���q�ҧ�{��4�r��^%�bR��%�Dpӄ�i�<\���繿d�P���;s���2�xNN"�N�oU	oR�@�\{�,�L]�Ȼ�"Af�h$��8�$wW��S�u ��x�.�),,�P��)��D��Ã���h ��Ϳ:�S] =1�6�w�0�U�ˆ��=�3Ҭ�7�@D�۽r	��9[}5[��ߪd��B�gl�B��,�Xo�.o��3I���;(�>�x��J�ĭ�əR��b��P��o�1ÞI)�ٚ ��p!��U��Ep[ϋ�p`�㮽���O[��Gv��]5�N$���������\���i�v�5�k�Gn�S��mdg:�reS���k��r���9�D�.�aV���	�Zq�9�fW����ɷY+9��3u���Ltp���v*(@�Z �`��p����r�z���S��[�eݸ�C��{a��%�ڭ��V0�en���td����|?���d� 4��;qz9{=�Xd6X�dI\�f�V��9�5���c:g���$���ɉ����|�� B��6auՔ5�Vt�2.6̖�v�Mߣw��.c{-�I;��6��D�1Ϛ.!W��?w��C�\����ю̙�1J�1�����q;Re�z��^�(���}mna
y�
�=,����J�i�N#vFt~4_Uj�k�7Z#5wn��ֿkKq�ߡ鎻��� �|� Q�Wym�RHཿg�
1�b0�Q���ҕv��B���θZ�����]%�<q�.�L#F5ʖG��bۣ�%��ɪ2�J�w�E�@�X��s���ߠ�m#��-��y�}i��Z���9�Q�xۮG�kY�]w9�lh]�M�޼&���(��s)P�k�b��L��e�f�� ��1�ن��V)�� �Hy��5&�`��.��ϭ��+؎��������z��bgy���bV��z�v���A����q�5���gG}Z(�~�����*�;�˼7�j�Q E�Љ�w�쁗x�^�5��U�h �S�6��:豎�쾸�hzx�A���r�J��H�G��)msՓ�d����WY8��wXU�ZsUl��W.}'��>�ꔯ�&)�ۯMf
7S�,m�G�{��+.@}��ۿ=���ޙ{s����n�	yCz�!Q�+3iTpϢ����_�3q{G�����粀�6�!�٢�T�����~OҗO/6W�U�$=��2(aA�̉�U����Uh��Ǉ���6��6��;�P�j���%T&�OK�Z����\���}�p:�:h\�4ņ!���,4��C�1Lf��iu��s����C�4ݘ��	K�
a�[Wd��&B�=��1ϏvC��*m�+�Ћ��R&�A=���@�Ƥ/mѶ|+��'X}r��,[c;5�].$�(%�R5�O%�^��fk	誒��/Vm��m��+IW���^���Uؔe^�"�=U$�>b0�c2D���v+��,�瘟,/���뚨״���h.ꇅ[acY�7=�
1�{�a����¼W[~�+��,`i=Q31�����m�b�%��A��wI��X�J�5*�!0�1��R�x����m3���N�,�d�E(�E���������V8�pXƊ���|�Ӈ�|Tܷ�F����.�+9iV$��(56��g�NW��"�~R�_b\�m`����u����e1BE�r���^iA������[R�U��&������X�?o�A�/�9����Z�F�i+s(��تT�mݺ�|�|���/*f��Ba����{�Ao3[Fv�Z+L��P
��A%jC6����]�(i��𳽽�Z]
�gP��Tݴ0#�*����#j!�(X�����/6�=,��6���w�wQ3oli݊]��<�:�: �d�)��wr��Z�p���X�n���e�u.u^�t@�7',��Εe>uj�������v��.{��sǌ��S��k/�����sغ�J%�����kk
]ܷr�;]�Ӗ��%��DP��_.�5��q��|9��٫�v89�Qx�	�G]^j�w"�#P�[�I��P/��,��4���Vr!x�*����Й�Q&�׻*=C�Qݭ��V�l}�ϮNY`��I9���]��֋鯺�#�:� �6�����B�.�g;uU���{#�y�]�o\�ֈ��ɸ�t��VN!�l	��mBYP���i�'L`�h��rL�k�;�-�/p�Lf�tR��3��D<j���R���I�,�OT��;.�l.4�wf����P�I�.hS�'Ty��h3&`��HJx@�z:�p.��K�������k1u_T��CF2�(zD�ܗU�#������)"����r'�{^s��9|�|C ���Juu����c��k}�m]�L��՞Ӳ�(͇�ws&{��H��d,��H�12�fvX�^�1�4��P�#����b�U��hSy�(U9�}r],�A@Aa�7Vy��rU=u��_�2Si9(��(b�9����k�j����9�t�2抱�����L"��*H=椪�����.Њ#M�CS��Δ,qTH���w7�#چQ�;�u��)MC�S2T�o�-�wf���~�j�S��Q�rv.)3��f��YO�Xk/�ɖ32�awiS��ޑ�̩�a�*������4��+<�0ݼ�/����� �%�$;ɤܳ+t������m_%�f��YJ�5x��X��B�@�>��j��t�Bڮ7F�2�ocL�:xF�f)l���H�F�l�}���`�K�P��Ս���S}낓��1ea��G
m�\�+�!a�9�"Eף��p�%-3WV����0x�u�u�!奎��][*b�E�gQ�K�R= �S��R�e��aq岊&�zľ�g+d��{z�<�5�m����KLE8q/��3���q��~O�&
I�k�<��~]�����Si��dY<�&&/�����1ZO.��1�+I��fm�{%��B��BMW��Fn5g����%lȀ�ۭ�fF;m�;��V��d��N�I 孤��Έ=[�M�Թ�{�G�W/]~n�������jC��	��G��WpQ+���҅c{�{�d�' mE#J9
��N�P���5:K׻UewP�������Z�u??]akQB���=❭��|5��]	~=�}��+/Mx0M�\�Fcf$c��-=��imu�Z���|���n�1OH���1�����b�û�
�S�����\�1s���4�� $�$�K�֌b���y޵j�X�'��WO����T*�㑑\�gQZ���k6!��㮄O_>��Y1'�XH�g�2Z%HZR8e��[��eZ�����Jx-W��:�L�^3j��ԑ�.�~���q饀�=�YN���u;�_���ӽNN���6��ǧu�����:�(v-�-�_��4���Ђ�Ӳm�fR�t�e9��;��xQ����5?����dQqFm/%�^YٛW�WVN���Ϸp� �n.�wQʛ]���w�&�u�I⍸ݒ�s��Qk3�ճ�>&z�ܧb�n8�7nr�%���.2�u��V�"c.68��*����[�Ir�G��.�{qۡ�ݼ�e�*��';��qb١�
�e�ְ�Ѝ�>�g����מ:��{�]qO�9gnNnMɥ�G��s[κ�����շ�}�8�x~�I�����wC����rg�cWDp�ڵ�0�-I,���*��KNwo>ϿL���9�_Or��<7��b� f����Sԭs�9�˻��Pxc����f�},��08Ki4�q����Y��h�c��'���4g�;�טeܓ#I�t3���洊ޞ�j�3hjQ�I�y��B�{�E����T2(�]҂��-�d����a�S=�/���º�TǴ�A~�OC�m�T�u�Ç})�M�/q�P��=ZN�H��2-$�-�OHֆ^�����-�w��K_m�����m�š��QȦ�+mG'�Y�gr�kW�B�d��!i9DcJ^V�{��!>�e����&.�flqއ���ٌ�ݾ�����i����m/�l؟�)ڸ����d�3L&���a	
Q��Q����b5<��.�dd8�d����Ɨ��/P*L![�%Hm�.v
�[��A|6�N3.8uv.���!�7��3D�Ւs�c�~�ыD�ru�M�;�ܼ�Z�Z��Qn5$��������4k*��~
ѐ\���o�5fR4��x1_l�:)���ˋW>�W��'V�&7*bx�Qx�����"���:�QgX���^UӠ�@ff��I��+k���������~��o��
	��o�h�3/��z+�"9��)i���¬�<�Zz�q��0�0��h��j��c�Q��r'6	qܨM�:����7O>�}���,�P�����s���Z1�b����X�h'���8ɓג���.�o�S�g����0��ă�DN���<������j�i���M���Q X|�~#��%��o97A%5ׄҽT�f�	�	K�]�Mm���J��*%i5���v���cM"^�ojs4v��D9��tq������m���cOn������u���g��so����6;smv��4�D]�"Ԁ龆�?RҼhY�6��U�[jg!N͋��ͭ=�m�ںx	��τ#���p���]t�\=i6Ҽ�&��қ:�ﷷ��-q�5~���W�kvٽ�"D����֔
̚!�~�[L��}�Yv<Ǆ%{�a�f���/�gN�H�V��;���H^z�_^�3���<�t�gk������,�U�2�+;tй�c/m��rMnu���5�`_��,�֥3d<T��9v��]Oo��C�OCE0�K���ʰ_G��i�8�lH�F M�9A��] ���\~�8� b�����&��+Z3rK~�W.��o�緙ꮭ�P�s��w�tY5i3JP��!9%�
���O=�c�mh�}�^��^x��`U�劯e���b�~ojA~T�p�o<Pe�n�e� �m	�Eh��1+���8�t]�{GiI����n�%�k���m��4�~���d����H&�K��n����{�=̭�p;��䖺j�T���J�uݑ};]��2����Rx	��	�e�
3D\��%^+b�5��5��=�����IIE�+�>���7�&d��O*3-\{N4J#P��3:/$x�e�#Mm�b��uߊ6e�� )'��~`�.�\��f���?b�X��䊑�������n�E
,5U�h�I�X��cQGy$@�w�� d�i�I�]Z��׭���!ԃ~YsČץ��y��0�Rd�wv-؟7��;݇1wZWi�4�x�Z�wدvk�Y}'�
�	�ѭ�QNj��k�1�V�:��iF����w'�y�d��ה��m�V�"dv;i�sl�	��6�P��n��2狖�
�� m\ޝB��P�½��]�U$���M�__�n�uА.$A�����:�W&�[m�f�̷�Κ��ZԵg���Ӳʢ�n�Ol��]�B?�4N"��Z>�m�S����H�ƪ��Md>�]Ӹ�.�kްފ�g̉���n�pd]�v_��̱�����3б�'T+��]�^�Fs���N �2�?y��{����9��E��]e�TH����$~��� OzJn����w��W����A\}���������.����.ۥ��*�-�����/�i6d&���F.���ѣ��\�_^)�+\��O�Xb�:Gvl3.���p|jݒB��y[���oyں�vwp����8��F�q�	�"����c��䲮o��Fj�t���}�;��B�̝��-^�g��6��^:}�Ո��h���e"�^5ֽpyL��?
��3��8�m�X.M�FGu^q[Cc7�˹X��B�R^��q��ݪѭΰw��6��x��eS�6�`�G	�WH�Ge�/9�IXS�>XnMά�I��WQu�3n{q���U�I�n�f9�SZ�U��n���[��G�UQ�LY"r)]zmD!Y,�=Y��ù������y�q�.�:)�݋	��n�Y��^�k=���vM�p&Ӽ��;=^���bs�����ĻXӫ��N�ma��]��6�c��	��8��6ڵ�[l��ϳ��&ݰ���&��=�����y�<ɫH庍�Rt��'��35��2B�*L��G�{�6�;y?n��^{��D�K��t��pTgUmI��H�K�o��\9��P9ۦt\Fc&.f��K|�y�0����]�M�69�8�j���s�q{�C	�bQA�\i�/y��y9Z���ܰ���;X�_������I�Ęj8��:o�c�2޻"��H;�r~[g�z�j��'�@�-����qyu�]f��M��=��*�^�6��iIZ�vWvH����z}e���[�~m׎�����No`m0����xi�,�>����������wjD������rD�fG$�������
�J�駸�O)��*������u�J��8ٻ�5<I3�"�x���Ku��[��dױ!<��=���Ǉ�`��D\縷h9nw)eڵ.�su+W}���z�bnӯA��t��-CקE�e=�N��{ԝ��y�ʝy=
a�z�bJ��W�Q��B������z͏{��n`���Q�m r�)���9퓳Tպ��A�b��hQ��wzp����M֫��I������c�XWW�Q��e�w���������ra�<y�U��7�*��Om�����ꠧ��-���fD�I0�8�� �q.D�o4R��!���.�3J���b����#�pe�J���z��7�������w�VR*3m6�m�
G�>؊��/z&�zb��;�t����u
�Ë��z;��s0*�9��{֨��<�z��0��`�5	2lQ �"�/�G��W��+c�~�@���Ʈ:�1�gb.#���Zs`�����xmX�o�4W�~�3}+�8B�y�c-�r&J+$!!�Y-�G\��q\s�:x�[��,�jR�mӢ�N���M�p������qg�_��(D������<�`Z-nt��;Pr̎�v���r��U��C��G-������b�`tѨ_!�ǝ|E�U��'�kO�ͱ 	�����%a��QɁi}W9�v�G�:�?`�l�I��Z��'�o�
�%M�Eg�W����ʵ�0�y��������Z�9��W�Z�Cj�0��W,��,gw���V����΁��m��)��mfd��s����Ѫ��L{ל��λuhj�+g7�A)�g��0�0�C�o���i�G3ٮN��n���׮�Kg)���7W��+V���ӻ��?b��(��Kۏ�_q��7lU!��F�=C#��`���7���<_��)�� 3��a��z+�	�r��q�Qlzz�bxw�J�3�~'��.��,�iJ�S?Pt��@z�!��lk�B,ra۝�V����\%��x��i:=p�]iI�Ыu0~����6ǥw���GiY���CykA���Oyk�2t�.��h�%A�}�휖���(����P�&��P�m�9s�)�s����px�PCM�x͇�4�3yѥf{.cƲ��2{=5�/���q�z��R�^衰�7�l'�]"
Fd3$��vvV+T�=/N��������ܯ/�r�y��q�k(Ʈj�9L�ɏVyuf�i���ʦ���|E�#h���e�������ݵ�o�Le�燎�o�dB�2�#�|h�ޝi�k�Ӄ�wJ��Wu�P���cq6���
����**�t�W��ٹ��S5ٿvQ�G��Ƹ���)�\G�3w��{�OL��Yq/^��1� �`�$Y��qٳ�ymdNaD4��&���y�t�h]͘;��J'�u9�)���g%�l8�M��뵲{V��c,Ċl$h0�.��*3Օ��v��ۧVԘ�mj2�y�QPͮb�j	a��8�v:���=3E�;�K��ǩfъ�=7���҉T�ړj/i���YIјh�u����z�.���p���邭�1���kM�=५��Dlu��^ٶR����]�)ԉ.�Usd*s�!g2S��{g�'QMD�i|�FC�x[~�,[5~>��޻gq�B�0�̌�4|U(1�όᚕ,��ip� ��Q8#nCK9�(EV��������tg�}<�h��CX�O��:�ڞN4��Iҽ�#V�^�����W4ߔi���q�h��n$�&����)��{����5��ufp�T��G`�����B}6�7X��-�2�ǖ�v�&X���U�S����ǡ�Gt0��B��U̶EN��[�9qYCv��7C���)�־�#)VVr�虨+�
�h���H�Rtޠ�Vnji�Ɣ���v��՗]V��E�6��'�ZR�CsGq�g6��G��VGw�<h��:���tl�/�1Q�}�mg�v��Ie�1���\f։��ˍ]�ŋMontK��{�(��v��ŲF��u��$����}��,����E=����r��l�,54:V_|����:�1�����w��$Q?�w�[�����V�	�id޺�&���1p�5��;���ᢑWz�7� co�\��yۜ��f],]��7�{7hu*6nhݼP⑫X
=8�6� ����c�;Y�s�:��j�%���n��1����'�xf��Wq��u$�ԓ�h���������]���S6��� ɦ����%A�inŅ��;�Wta�S8��d09pR}�lP=ٮi�m���$��ur,����,Nޭ9�[�n�m����q=.�i�����m��5V^gN�B�Pv���ТZB�`:��s ��wH��J��l���#��K�ɑn�I#im�
�}en�J�UXmޝ��}/9v���,�B���gZz���V��Q���y��N�E���6�n��|6�}yOa���0�� Y�q}v>q��YGGY9��6(�P![�ûRc��w]�&�]��EeQ'.�F�P@����C��w㹢�q�Ǚ�ΉW|pq���F.�E�w}(H�ʼ��!��ǈ"yEJ3$r�	t*��dkжi�B��>��:��kj,�2f���Z��x	��ե�'���ݞ5���K�wDv�Lm�曭]���Pa������S�nۗѰpv�2�g�ʥt�L�n����q�Yhz=��n:]�ƭs/Ql&z��F]�]u�l6l�>G�\;��m�=��<���Ÿv�#�%�G���vHb c����Ogq��}\�_i����B���a.��glF��.|n������Z4L���V��EaQQ����y��5ۆ1iG\k��c�lsԆ�9��BҬ���6��j�_l�I�F��OWgqc��z�'9ug�k���z{z��֧��C������j�ݎ�=�v�\����A�;q��x��$w$S�$7C1n}h��-k�(=ʞ���1��-vx؋KH��:,k%���;y�Mq U(����hgn����'���z�m���N�L�.Sq�m�V�k��q�ݒ^P���%]c�&^�Dۮ�r`��+�u����c�cGe���{tV7��5Ni��+Ҹ�*�<�bW���HѭW�e�ySn��u�� �ڹ��X���k��:J@vl�.nr��p\�O'l�Oo������]&���ի�<�bƺ�ܹ��V06IK�`��j}�:���c�ۮ� �'Oם�m�ǜ6\�hup�z��+�X{z�w �8�N�.�l���z�k��ps��t#�z�<gt�2s���bq�	�0iT�μ*v�^�@��ݎ^zN)׃L���Nsc�o]��>�]��8.J�u����^�m����|�c��;���^��r������n��0�"�ŝ�Y�\��`�Ξ%�챾7m�I�kUχk�-���o6��;��>,5����;����[���b�;a�Ǯ6��^up7[��ۮt���m�1��g�������p�y��\ݻ6�ލ�]��3��G��n��;��9��Ԏ�����,!�Hp�M5��ˤ�h���N��;nZW=z쩯dy�<x�F2�������9w�{|�묁�����6q���6�]n��;Y�\(�D�8���}�[shm�9�p�\����&�u�s'��}[=��4U�:����p�a	�]�m��wN���,U��r�-��ۙ��;s���񧝪�ԸNn�tl�������˵�On�=�^U�����\�\\���6n�e���M����J�0ɶ'�.
����׫��t�ee�������矉�x���	�ozCv�3Ogg�\>zp˥���ht�
u��a;ml�K��+ǚQ�#*H.�2�����F�s.D�{��u.�����"���M�//���h�,9���<=�m�W9�6s��sבZ�T)�iEFHI�W!��ѫ�W3i��C]��v��X�gMK���ú�K��`�����w�^�'��=��_�E)�9
���EKО(!#5s(u���iWNкů�H��Sú*�/
���O��B/gs'�%�yud��2#�Oe�TI�E�-ڎ8]w�u$�����:wI,+�9{R�/�̄��3ػ}����2��->r�e���
¦�������u��Ln�Vs��<]�*���W#�m�G[q;�-�[K@3���<�F!��\&����]�^�(5�����!���:ÇWXH�ؙ�SfN���O.U�>��>��G]ݢ|���H�� �]s��1��#��g{�W���Ɗ��\��5�mq�����ө��/]N�κ�pƁ�Q�S���*���:�U�Y�OK��\-�*�;��e����Bf;o��nn��Eq+7�����5"<g��h��YY��D�j|�IĔ�g�j��ʛ�����](em�y����lm���͡�]s�.���A�c{+t(�K�2Kpǿ���x�WJ�vS}����w��ǳ-�O&ߙIx�r�����a�$�c��5��ک`�]�k���<1�O��AD��ԣe��
��P�%-p�"^�]-V3�6���5��2��u(����P_K���Or���ޙ%�:��.�û@�O?�k�/]�6����r���pP
�g�܍/T�;t�Y�Ok��eJA�Z����(-�Y�����Y��u��W��)Wq�>�C�Z�#��a"!�MY�G���ƻ�hKnn
e���ܖ �;	��[��\[�o�ϱ;Hk��1e���2ȉ]�򈪩�f�V�\�.��\����ȸd%r6�i�\(��b�zS��6�Ǽ�>nF�f�~�6W<%mds)��/0�c�<h��̮��J���Z^Zç��_e%�'���#�ǂp5�P]��[��H�mk����UЫ���n�:o�oN�:��MZR�i���pC056�d���K5���5jֹ]@��t8ǎ�u�)��wf���p�+*ȯ��!fG���B�%CP(q{"���rߓ�B�H�T��*���DeTW���q�ۏ�4F6�PP�E^�Чrn�:�ڱ6���m��Tr�ӧi;\��۪��x� ]��7=1e���C,�y;;]�k��_���AZ7^5��4T�S�b��R�p|�zt�T�b��DmÇ�x�R�!�d��9`��PI �n9&//d5;�[���Xrziή���:���V!~�svc��r��~�~Kg��2S~���o	C�-u�⍇#e�%F�8��	��l���׵��|��V1E���w�k6�Ù-�_�'�G�+�d�(ߎ�yƑM:���#m�RD�,WfQ��6'{���:`:l�2,����o�)W�X)�U�mf,DQ��4���>���˒\��=iF�*��Tڰ�"prQ��͝�[z���gT��up�h��Q>`Cx1�(A;,^ʖ�z���I�8Z;|.}�4O�J!)���8�v�f*~/y�Δ�`m�C�5�4퇤/s�>�_����Sɹs|�?h��`���>~=r!���J�D<�Y(��r;�.����������M�C�g���;4u4��<�[�0�6��n�2�T�38���$c��	�WO.zvǵiC�=���qԎ�i=��ᥰ�=�����v��"'
�>>gaI8��`j8o#̧ݎ�Olݵ��qrb��x����#^�(@�<嗵�m&��s�ʺ�e��ԛ}��k��o�!�jF�1���UO�>�'�����Ϯ-�}0�x���]+�m�=��!e�,S1[����U�vU�C|��e�����q<+��w���H<�1���
�i6�+��&�^�=*��+隶!h��Qw���`��D���8�k	�2�0Q�s��^Xϔ����lL������r�t,xo���2��xz�ρ3�s��zK��]g��:Z�<������6.�+]赣���F
,��4h����,]ge�N΁�\���r\k�����됺�T����ue�!٢�M�v�ny�9u�7�\u�yd�6 �#9��s��s��8C���D��k�V�P��l��ɋ=]L���n�<�*�8�c��Gku-pr�l��Y�uc%ͻg���8�C��?�s������œR��;6�^�86ۚ�4�����Q�@��Z��mջv����k=Z�zn���6r�ا��TN�0<��`�n�<����Y.��D{w&ٖ�g�su��w����h��<EqY�p�Gc5đ��l�R[]Y�¬��yᇟ��{�^#���sĈ=z�	���j���f����{��_b�!a6T
5m	XÕ5���G_W�.^ў!�P`�o5V)|iB�'\�+%�.f5�w����i*�m�Xw,s�5~ve�7m¡.�8�-����g�yl�Z1G-��;��5�����w�ٺ��)94����7�]^���B���%B�m�5W7�i�U91�������u�5�j�rb����:Z���D��N�:K|�FN����J_H�=(d�� �8`�r�ici����.K�5��Wx�z��\pc�vz{c�Fq~+��*F��b���B��񒗉�.Ԍ���q�ɝ���"f&�N, �-�p�xz��'q!��Z�՝�E���#�%nB�R��6%%��õ��}�m^e�@��j��on�������\�ݧu�Sܯ��5T�>�;�Y)f[�k"	C�H�8+�kHS6/3y�j�>\�<���Ue�W�tr�Vqk\*��d��9-�[p�uU�+���9��
_%�e`�γ)9�\�֌o�����2����{*7H�W.��^�{�BA'v��ߎx�/�^�)ڧ�[<YB��T5){�f�xBI��|�a�!�Üp�\�P�����
���yw]�B��J,��ͱ|���}�^��)䇱L;t���U�V�]ⱿdHIa��;�1�|'k[0r����/S�$�_��>�uQ�'��zO{�Z�5��Y{�%[����w���؉����FnB��a�I�����IN���dY�Mm-�<�"��r������"��JR�e	��R?5���]lO������=�j�]7��� �J0�̽h�fz潢�l���p����s�ܙ1v��Z{2���7P�mJ�b%��ؿv�gm�3�~˛��M��o_��xNK�P�jg6����ץ��zkڕ\}�13�I�b/?TNy������d����C
��'H��(��C2˽vF�3}�nx��aW�^�qeB�M�}@�4l��y���}�ۻ@TF&�a��*�����ƻ"��.n����J0ޙ�U��9]K-33�	^Vn���bn`䖰o�$��Bs����C#���
Zgjէ{6��݊9g���B:i^ީ����Y�9@�=ʺ�}I�T{q��eD��~��}/Vp���y�ʄ�]9i	i�x)�Zϻ�o�I�{�E���zI���/�-u�0a��^9�:�h��NU`�*n�}�g^j�Q����� B�H�Ch��WU�=�����5J��>cX;dY�w��$��z�|�+M�u��W~֗<�*�8Vi?Q��ۏ_��{r;[��	H�b.������펭#)�oN���1�*L��.��h���D��F�ܮ^{չ����v�h5����J�_w3�W�7q#�r�f�ؔ`͊K�����VX�x��yf�&�@�L&ث�%£M�uv��7		�[����y����w�\o4ŭ�����݃hIkӏ���yK�H�k�*B!nB��]Y�#��Qtn���OzT�u��E��$uU�q�P*<Nl�}(Ȟ��*���T2���Pl"��D��_�yZ�Q���x�����wHp�y���i�J� ���;N���ޛ^5�h�l,�,a�Q�wf��Iv�,�P��6��%>�����9X�����c�6J��j'�����kT3b?*��H{��k�E��ĠRI!I���b�����"t
�{1�EYf����jem`��@�6U�ǨC%�����D���0⫬��r�Q�B0�k� Ӏ�`��.�C�t�mn��º=��[
V�f�q�	�Ap���.��~�oie�����::��u2,P����*��$3����ݛ��W��wh�z�u-���h5��!4�7~��l�Y;��6��VvW���A�R��{����X �ӂ��s��IE;'�x/x��0k٩��(GL�'��(#.'�	�@!����������==��I��%"�9=�p�5�=��>�̇�r�	ORuy�������~�$%��$zw(������A�=�נ���![]����}���^:) �.�]7�3TU�~���~6��j|���6�^��������GJ�φ������T��g(�޴�{���qSq��&yix�ܬN�xY.{9�q�-�݋&2�=W�6�M�(��T�nV2q��`��k��\�ה�3z��hb\c���~���ݜ�Fj���F�rr!l�p�3�r���N�w»@=��n]����YE�򅺛t�7U�{�Y��]n�c��j5�2c�m�g��O��n}��Ƕ:�ˑ����f�v7ɵ�9�����nҟ��}�B<�:�����wl������M�lЀ�.L��'���r�$F榌��x�z�ݶ{>9��wn�w�U6��z9|�[CE��a�WR��.��:��[O¯>H��Ѵ�=��Ѳ��X�]�r��$R0u�]A�N��/د_���G}Ί�z��͘�q���������K���g�[��hb�Y�>5f �)Hl�"����cf8��u��Sb_AF.nCٻ�(���4�V�KQ'��n���_��f^:�r�,3_�a�Rm�nֹ�L�����⩛���7���P���q�8�@�R���]���c���dX~1����©Ie���OLm�#o 2���(I^;qp�ߟ��S����@�w]6d�s��w2�]D-:�]���ƕ��k��$hP�"�}A�L���OZ��P�������y�ƻv��i�O}~��Ϣg���G	5��Cs�7���=D�E���^:�ە�x'�صD��K�3�c��;B01���qLn��sr9ḫ?T\P~��ܓP�u}�J���\��w��Nݼ]�u�2XDZ�g=����E����|�1��nG��[I�����4��ƚW�D�-®T���8��+��8���}O&���G�4�޺ƍ��͎���WT��fbZ�N島�ӫS�b]Q]n����-HS��\�G��Y�ƕ)���O]������)��������H�܃Δ�4߮����igM���8bU��cљ��f��}4w�a�S/��5�v(͢�ǂ��H]��%��.	E�S �?S�ΞQ�c7�I��>����}s��@�������L���j2�G�z�>��<��[-��$��z�5d���̒P��}ޤ5���w�u|��4v��d�T�:g��͎��5�Dו�N�:�2�du�.���˧�ԹI~�q7Mf#�Z�R&�i"�U��(:���8�q�d����u�/A��]�n�[x���phQ��n7�O�ݘm���-���<z��uGZ��2LXٜ;�}(�S�O�_��8bV��w�_N�@��@�ٿ�f6RbB�]�k�Vw���K���Ptod��8�zpI�G\�rU�2&�����BE�fX�f6jx�ߤɱ���pF�0�-�p��@�3��/wT����nn:��,�z�[u<�J#"}n��p\a���X�R��s��ҩ�b�g�zԭꔬ頒��@���-=:~�zs���x��v�p{A�)�+t��i���o���j	7-SWoI#�q�+D�bʝf�]S�zY(R�[��0�.G	r�;;�qH��N�V�%�iV������k���=�~ƞ�PI����TX�_P�s���&�7��e�)���Q�6Z���4�����7y��L�� [;f�[M�`���^6�VswO�n��R��ؔ���uuH�f$T�ZU+��T�n־�+�ݹݷ��4:u4�e�̚ulY�ٺ����{�Ȃ����4��Vg:�����	lfѾ����]��D�l�*�f�C��]>K*h/��
K�X�7/�m��Y=|�n�����S�Ȼf�{�`h۽�]kXe��P�8	h5���� ���.ab�����B��n��g�"���d͒&�rn�$x�j��y�ێ����l+�/�YT�oM�!]���յ:�(Sy��J��V�6q冺ҕ��n�b�փ��,��E�8����r���k�A���ՋU3E�R�'mZἎb�naLKKٚ�>�6�+Xw'jEue�5"M*9�XN�{6���j3khЌ�u朾2�V�bP��/��f�@�"�0L�ìH:�c/e��]ܙ�`�z�D0.2�,=��}j!1����4s��H��im�B��tʒ�b���j+�K�W�8�M�׳Qr�YG�b!s��<��1��r<�e9�^�س�c�F]����]�t��y��T+�ϐ2A"��Z�ݟT�}\�h���:�0}��WmXWB�����V�2i�a2'��T��֥h�W2XW�y�˹�|�Y�+jH�{:8���J�0$�.E��$&����/��QH ,^E�Y�6t��Z���痼=	��.�.2��n����N��Q�߇\>�v`����_F4�b �̡����@�i*g��*p�
Y86��a���9��+��,2�@�AqD$�{�����T�cݮ������(7���w�g�o5�\��V����>]��z�-P�rJYjKs�_��0���f4�@�rVJ!r����j蓎Wvb�n�>Xr��
{Pq��jD�!ii��}���Hl���ݷ�h���S�]ڸ�:�Ǌd6q�I8Ґ��L�"��D�`.��#����m�TDHveYS��U=c�����x���?nW�������f:�j��mk2f	�v�Z8$(�m�ӊ�0�uB����������7�/+)1'�h�IGMrӓ� �1R�׈j��hH[~S7��\ؖUu.Ͻ;�\)�2J�+�7c\���.�aU���>��.ք(u�|�*CH��H��^^��E1g���Bp�����n��ЁH���9���"���&߼'^ֿiAg{v���z�辮��hH��Us�wdQ��"Sʐ��(^^̘�r�"͝��5$����jRs90�]�e��a�z��IΚ`��*d�]�ݶu�]U�y��m�1��W��bjn��eM���7�!v_r����\_/Lt��C�C)�¡K�b�mZ�m��Ww)������K����4Z)QhK^��e�5�N��LsU�~��ǯw7�{{ݡ��mУ��YW|�'���{]��^����w��Q�k���FPH�$n�e�,��}W�������5z�ҍ�w]�9cm�לh��t�ݭ��!\��}W�_�8`K��n�d��iAM�.�
�?y�y��p��!�n.��S�����m�	�g�sR%p��="ڂ���5�]�H��r4S����mX���1 �I��6܇���k�@2:{.� �4_Ȯ�ޮ����\��w��f���X7��ћ�2�>*�ҿ[�t2{Mғ�-CkO840哝q�W��w���v43&�J��4�o��k �To�2���.�f7�:m6u5#h�#�6I'v6����2��zɪ���v��_g��79��c�{wU�>���\۳�;�ey�:�Nz�]�wk8���dێvU��㵇��a�k��d�<�۶�ն�.6^���ܟ{��(�����i;q�M۷���M�`�髥ڭG\�ǫv�x:�C���'c�%����ԡ���a�w\��!��mU�jܝ�rg[�i�k:c��nmf������>uᝥ=&��^��˦ڊK�, �6���z��?�����>P���M��w
H���8��ش����ܫ~���r��H�!3o������p�ͳ�ڻ��"�����G�ـ�m8�
9*��B���e��=Y�'"�9�'[��E�]�΋�\���|��2���u��o���>���s��1�}I_�rc��	F0D� �&��*���ҥ���Ѫ�v(�"��*�l�wL�5Y���Sέ���,��K2J�����[�iPs��������T�n����w����3�����w��H{����%�@����h�f'����W|������#u�)�\U*.���l�&P�H�a(�rc�>�d>�����ؖv�>��u�U7�u�[^���R�{(Omn֯nr�V��u*$� ��5^|�WQUG�-q����=x�3FmV�P���|��v���m[8�[tn{Y��F�	�T&�Rꩠ�vTVZw��:���{I��p�>.��x���|I��NG��B�.�>6�p�L�@���{�u�x�{�>�M%�b��"�9
�h��dT�O	RD�dh�߯��@Zdn`�Gy���q���:ʋ�j����kø`ݢ�x�R�Zu�ُ1�C�V�5�7���Oa�x����Z��^�Zۺ�cͷ'��tzIJ��= �	U:���v�|ݿ�L��	�9��{�Ek�JVh��%�,|&�|�s�7����^��LZ��0�BL�uQ��;\��fu�C���E�2D�B/P���V
dx�V.�噼-A��^�y��S!d��6�:�ya�X9���+D.��M7�S��t���L��(P��Z�'6��X�Y;����#�i��娆{HN�v�ាRY'��R�(W��pB���r���矝�D%��p�cD���Z��Fxx¥�������̅wA���ε�E�1k�l�G��,����[��/*	�	�>+���ㆎ��ٚ��nC3��;��,�X��T�f!��`����DW�QՖ���4�d�P�[)��a>�x�s�6�C �C�I�3}�o�இQW�+[P�-���O.���Ct�n����%Bد�E�J(��**sX_��y�"&��S�4��}��`��_>9�������c䴛�C`�IUe�^M՝�,��kf��b4�́v�Z������3�I�2P�u���a��s�&w%00���^o�bO.1�.c�0ݺ��0�� ��\����<�	��N��+:���(f��W_s����ʞ�=�[�<ls����3:��Y��G��ϵ���p��j�V��G�����6֨7�lM�;0g|��[E���z��􏧘�ezR���ˬ +����J	�UY�&I%��t�Bݺ�I���ks���D�xջmd�YW�q�Z����Nw_��'xr�܈�2����դ";�
�iKx�G7;HyP"�MUk�<��IV���������2��&͜�~Hj&�;�E>��G�&�V�&������k0ӽ�nĹ��2﹉����"�{��M�kg2͊מ��5�U�yࠌq��m���!�f%���*���ˎ�����p-+���<���ps���M�X�̻�sz�����-<�g�����&�0!�M��v��if,c?n�8���ý�Y��z_�a/ܘ�!��sQ��-��������^_�Z�����SEuN��L�U�q8�,�2^���sl�=K�y�(Ⲏf���z��D:��a��fAĮ��Mg��c���/���I�_�9�6�J����r[���L��|g�hO�۷u'�*��h���͹�&�"h��C\|��(�&U��BΩ��������Wo�4�?o�������Y*[&��n#q�<���a�%�0�vh-�YM<�9��r��d0�
	Å�A�}��:��;��	e�u�6�U���`��u*�G��I釿f��ν~��������2(�!�Ifd��f�D>��"oĶK	LD7�cԄ�L��X!��E5���r/8]g��^�{�_�H�M1QOD�_D�R�rn�kB�����+|������ѱ��^m��;q���XJg�#�9-�����bUN���L�h��
��O�">y�*��F�E�loi����d��I��`r��&@� j�
�=�~	��0���'>K;���?+r���w��ؾy��v�p�N���4�_N1��I�}'�_Z?)�(���_��7np��r~=��շ#nh���V�B��&�	�n���D�9���f۲r,$	�4o=�'�?e��/\�b޿����o�9�oU��1A�~��}l�'9`�b�x�c�T�sg#�&F�}��',@lM�S��Z�8�Gî�h��`uӂ��7o��x�؍����V���I������g�i��ϡK�H^������g�Y8�۫��v��XȀ���l���]�^�mv�C��x���t�0v�ջq}�����@;`|�c�7�jUP&��H�42V�ۭے�v&�5ی�����np�ÍԯQ��N���5׸��v�^fgn��:�+<e�ݨ���&�.�����W�p����usF��
�i���N*{���8�l���vmcj��=���,N�OV�.��naǕ�c������n����MD6�������J�������d�}�T��*�n`d#y��)~���A.�=�B;��P��,�[�U㽪٣~�-��N�6��R_6���I�M6�2�a�ug�>돱p�^��¨+z�j�{��d�"v�Y�~���~��f�L�	��x��������������|}�>������o����irB�侇C!���+�ﾏ��~UD![v%)�j���ؿӳ��U�.�.������s`�����=�F�YY*>�v��5߬v�!J�Fݷk��z<ύl�D}�;���Fݾt,�n(�|�U@�~��`��}��V97���\��ܩ���1N|~��~�_R��*g L��v(���l`$�X,�t��z�.\�����{��I�~=�qݔ�Z���fjK�fZn�\wѺ��{��w�[�'	l((���' fr`���ߘ��dہ8�f{wmkaN��=�k���./��\�Fa`,eu��R�J��*�U�����7��8�p�r���	�n	C&s����G'�91�d��*{���Te[���xT/��+J��?�Q�R��3�����` тa�Bm�pŭD_L�}qL���<�7�j_��4��6�P��Ԧŷ(�<�ʳq�}|����u]iS�j���g���̀�|m�fZ�8�]sLy4��t}�nIU��zs����+ّ)��W�^��;�#��=�ȫ/e�ܞ��T�������$����&��@���P~��H��+�"㾜{�7���e��D��gu��u���3���$����3B���Է��7�}��^D�Q�p���m�%�DC�X"�VdT�ﴡ�P�2��y�hZ��~��L{E���r>N��56���&#�I�>�#���<2l!��V�42�I��
Hk���(\n��~�w���Z;�ݨ
�:��k��3��Vr_�c�͙�k�3�>����e��rs+.:jAjt����;�������@��Me
�n��<�@n��v�%�%�9���Q\�mǰ��͑������?�jR�����5����I�g���xh�\��-[n|?/ҁ��u	G4`�����_N�g���26~�}]���J�>%�C�M�wN��}�[̸�o�:nu��Ի?=�ꯑ�rZ��s3���?����u��d[<l�]�vSP��WGź��8g,����{no��7pa��6�i�����}Ӣ��_g�n��FavNӺ�|����hб�3�56�f7L�q��b�3���C:�=Qۧ�7��,:͵oqG�9��Z�X�f�p�|8oVK���m�ݡ}
�@bd�ާ��7?<i��J����To���3��|.��F����աW���JH&a�Ⱥw�3A�K�9v2O��Z]�_�'O�),^���Qw`eߌ��°����O}ϵK��/ܑ��)��X�����Y$�Z�8�Ɍ��{���b���b�+~ϟ}�X�����=����!֎�5)�䇷1]��*�ܘAO�ꈱ�߾۫ssCX�-�c�u��n�s�����u�tv۔����8y^Kh���ah[,,V�5ο���l���o*���>S���NdC��O�U�ф%+~<��EX�oS}W�:��@�k>t~H.�l`���~�-h��ǮvD}oh�X�v�P�?4��ȷy���o!�_v<�K�� L��~�ݹ��N]{V�Wv�:C1ְ����pSp�v���ҿŭ��M����(�T~Wi�i�;��Օ���o�O���2�U�d�[��m����I�Z�}s�Ђ� ��B�)D=Ͼ��O����3Ď>���沧G37O��}��{�g�Z�}K�6�A�8.�c=�A�%�
®�f�f5��͗/�����Lb�F�,�	�碳6�˵���*���VZ��`Ȥ��aw�����܈��i;�������p`Rn>ß���'W�fW��&ᱟh��F�Eoǣ��&A|!�8��ϧ*+)���b;�Tc� ʌxb����ϸ���S�_8�͊q��f���jYnh5		�nV�.��$��Z�"v�{\��^�G���|f�bH�_	�?/�vn�a�ㆈ�.*�����ј�]�����'��'j�2���2P����9�Y(*�҄LCl�j��j� ����2�
��{>`�=�ϙ��fMb�s1��v����7����n< }��~�O���+�h���o�A;���$�&DB��E7�k���.���9_�x[�z+���l�f�3x�g��~�B��o����aW<��MЅ��G��A��Pn'mQ��w+���Gr��m���Ӛ{蝃3��d�"�T`<'`}\tǩ?eK�����C_8@ÀЄq<��%وݯ�foa�䙴p�N�֢��R>+�M���;����sw2Զ����������Pz�*��B�3B�;P��*�څPv�T�A�B�?T*��
��P�ЪU
��B�;P��*��
��B�8�T�*���d�MeYȈ��f�A@��̟\���7S2��I(R� P*�֔V�fb*�� Ԁ�-�BET��ĐP�l��ҥ@P���	U4j�
�$ǀ�U$ P
�H*�@P� H��TJ�$� P�(�R��E
R��R�$�PP$RD�a��(((��R&0T��эe�}�ӭ_u��f�����e��}�_s }�}�.�{�4���e�=�����r�>�.�|�{-bU� �����36�۷�7��  7�}�o}�!�w�s��c4}�}) �w�����zɪ�m�޽�W[4��u����x�v�޻��Ԋ������m[{�{�Xl�7�_p��\v��z�l��{`4�  7��TT�($HUTP*�����e�;�xz�wy�ט����w<�ﷇ+�^}��4��|�)H��j�|���`y�;�v�ϻ�}�s�Wū�^��x>�^��p�v��}�3�=�����a 
k���6z
ж"�N&�J4 ���@p��;=k>ƀ�_K�q��vգ^#vґ��c�i@����А_ tGF�vz/0����
q���垴=��]�
 �xԔ =�T��((�(���qS�{���S��:6Š��;cY'��
ǠT�k�� 2�`�}`�|�
 z"(�gA�
��P
:��rt��aր(��D�� hp�n��xz��ڮ�ym�zʼ}HR�������}x��;j}�:��Ʋ���=L��O�:�Z��Fx���}�oH��ԝ��]L�����itX��:^�lv�  }�T �
R (=��fm���r#�K�c���:��^�)h�}���Ҿ|@w���}����Cr���|a�k���a�nx��홓s���_a�[�������5�<��1Gy�OX�s����S��T���}��^-'K&��;ݼ��v]�{܅��m�}{�����*��y_mko}���v�����}���g{�}{��q��v����F h H�=QIP$���@
PW��kkI�;����v��}�ic�����}�����}ݦ�E���w}��e���u�wQﯾo���o^���b�����oJJ���y�ﻔ���;��vݻ�wwǹ^��P� 4 s@�����Bi}� Z��ȡs�@� 7z���K�����{��ۭ š�·݀G���}�@m��8;�}�����`�0}|���Q�ͥ�;��<��S��کR� ��b%)Tm   �=�&��Ѡ�'�J��   OȨL�H�2 ���� x�����������������
ٷ��+���z�;w�9�K�9��UUT*����� ����UZ
�����UUU
���UUUP���
���T@�UU@UP�9������X����!Uu,�Kri�o]�Q��^m!z,�c���P[X�U45t�հ�4f���Y�Hjh�׊!o#�j!�f�����|E�����x�VVbV��XƮK�aа̕
ɶ�#,�b�a��,�zq�9c��|F�[n��Q�f�Tx�|�#����Z�[��ROӠH5]��U��e��ilʚa<�Սl�i���8�pޔ��.��(F�'38敺���/1H�AgRt6\�ڎ��i��Z�ߢB���(팣q�y�y��T+e�q"�ݼ�GA����L&7���:J&a{̦i]��-�G�5�
�Y�:��y��h�tP�4K׀��"�B�ÐF�en��gs�A=�J���t�)+yEh�z&�w�BM��VV�(M��_�2���s]XL-�m\y���&�rGv�p���"�]0�Պul\�-��SLٶ�.AF<�/NuN�5c ���4j����j�����%��
nI����%�b��R��0�Y�*!�ۃ.�����Z�`i�H@�5*FA��6�teЅ^���̢q�N*�"��.��'�+E�6�SG+f���C�gp9�t*y�q��k������%Լ��v��w�N����D۱�l]�&azL��3+A���j�DHA�����Ū�eVȄVa��]�J5�j�e�m������1���ń-�S�.�(fұ8����n�I��6��D�ۭz�S)�2F�6�`-옋��%Hn8P��i{	�VҷS*�x�޲r�n35l�/[�J�� /Z��<K�(�� ���X�vfdz�f�8%7t�S�d�Ҩ�,�ߎ�Ժ#t�����kT���b\��.�Jj^�E�Y,V�Z���{�n�����*-$��ѷB2�5��� �T�5J��
���&a���  [x�J̠um+Pwa��+F�(�1���%����`�55�X#J���ۗlk�D�7J曛�<��5�H�E�ڑ���Z��/��:�Y��?��z�H1��c���+��B�р�7��b��$�*�V��NcV���(lA۠f
�w�8ŬQw,�;�^�r�V2j��K+V'5()�ENnZ�'y���@�R|���:ٰh�27�黽Z�J��'��F3���c�Hc�����a�Rb�w/S`�6�،lj��옡�*��Ơa�w��&(4ʨ`�c�\Ɏ�����2��S���ی�sbgɵ2�b���Yd�ܩBDU�!��`�Ȝ����{
�l�$�n��#B؆,�;N�����3�oҙ�]X��d� �{2�@��{�;y�z���d��,ʻ.��J&���XXSxF�!�Z�4ɹz[���r�7`^���Cխz���lh{[�A��aV��r�	+?&
�c�F�[787�U��ES!KS4<o�{���ۆ���2;�V���0ʆGUZ��ɣB�R�m�"�qnO���*�'$ �wỐa�v����	Qm��%��ɉ�#R����@�S�:��P��u��5L�,b�l��`YeK�CE4ͽ���M����bG,Y�f@H�p��hG6<�D��Sɉ�F�r�HV1n�Q{B賖�Y�IS %{�e�s���J��)�ӛݷ�Q� ������m�:��q���w(�q���ѫ-3dRt˫�Z�y��g4���`Z��bU��+v��Y��QJ���V�����jI��n#z*��&��˘��#[���)��W�s�C͚Tđ�R�VK��Vi�u"��r漡D�^�T�ͼL�EF1�Ǫ9y�������A}��Lk��&4�6��ʩ�/a�U��d��0X�c^��{{�փ��jB^�tV�t���P�[q8�73vb�XE&-����
/uK�H{6`��9��yu�V槮�i��
�bf[�#;�_::B"U-Ю+�i٦üun���JŹ�!d5Z�І� d#D�W���O��FM -oo�p��f�ǤO�<�4*J�0�8���N�;ͻ��3-3i���H��$Q���T�O4�;w!u�Z9���]�l�K�J��5�KA�6^�A�~OeKJ���m5N��=�m�f��JM��!�+�U*a�muo�A�4w)�ڟed�\JG��YN�>'Lcl	��΃G
yD�7X4m�y�g�IWd�C�7�j]��Bk��"L,]�e�xԂ��F�;*�����)�h�M5�J�^�z]5��w��.f�w�T�9�eP��pZu@tf�]��8�c"�y��ܰ�)iܳ��󱕏B#���P���
j�'*%gE�hZ��lK�)�EP��/M݈jUrp������f���R���gq��;��J��P����Ӿ�ݬ]6����E�T�l^NI�,��U�'4��wl=B���ZhG����t���P�C���lŦ��d8��^Y~d��y(���P��i^��u	Դ�`)}v�2�Z<��Z������y ��/<�#���Q/���S�v����7�p�@��Zi�骾-�oz4&�f��GB���/mc���o�(��iU<b4��.(gr�y�5���iT�#�P�@�̇F���h��DK(#�F��p�	5}��#Z>"��9�q?VLւiqr��_�E�G��5�9u��}q�	�9�w�u��7F��f�8��q�|COF��˖���3N�-'p^���*��nbKw8]\�&k�ǹa��]�{2^U�"��QB�YKu��V�B�m,Lە��1vd��x��˛	j�C���V�P�������^Tb��q�}8�bUK�`U��ʧ{��f����C%Yˡ���H�A�@��&���v�̂X3��w��f�0ȵ]DZ݊���Ò���h'��FI&kj%N���(��Lk	�Ѵ=Kfe�r�^޳ո$U�e^��̪�ݚ@Yf�KF�����)De�ł^	6�i��ܻ����oE�m�1� N�"�B�!U���J��7�l�3r]��Z��Ёm˗��G% �8JU/ �V\�Ŗ��іk1
o�_i�7��Y
,�[��5(G�u��-1�R�
���Dl��.����:����Zd�%�8vm`F6o
�m��V���T��lm�ņ�p/�l���*c�uw`���J����~���A6��fKbU��U�9��hC�u>�k���{��rQ�$�8�8�Ew��'>*��ZgD!��e��e��&pS3l���z�Pm+ W 2KEϚ"�
+2����Y���H��	bPP9�FZ�2��yi�׃�T��-	�.�q��m���Wy�otP"��R�HWfK�i
�/h ;6�A���6����ՒΥ��`���ӑ��m<=�
�m�y�q��zv3�5z,�	d��n��RVF^cX#�U�a�C`ݚ����/Iҋ� ��Ƃ׎�54��5#��k0+�n��t�I��V�Xz��7vQ�ubYv�)f��S��1i�]�)���.�ZO����v�h��b^��
���A3+A/e((�zw4�9mM��ڼץ�2�;a�3Y�j���[4��$i�x�p��r:�-ꗮҺ[�,��J��N\�n��ݘ��(���	t1��+N�b�me�X�NM��9)l��ڹ�!��iـ������w��cHUt��wB�X��$�J�f5m�,V7g���0,��!tUk�zDۄT-��V�������&N� q�Ǯ�"��v�S�	08b&e�-^ޑ�jWJ�5�-�z���R�0.U�f=y*c�����v]�0c�I�5�t�J������M�A#�S/!ڙ.���oZ������Bۙ`����:í`ï��_2�f�U31?j�n}��t�#�J �It�Z�`�r���QbP�jL1�12��w*�[(���f�rh4Ej�e����F���]n�.D�UU���隘�����[�
:3i�)�T��՚�C�f|�݆�n�cUn�r�4��� ה����j�iC��Qa����dȴm[MwP�\�,����W���)��n*��=7LT�e^-K�-����q�B�h8j�#Tȟ`y���U
����ûm�U>uu�$LG)����Nmw�zQGxѰ�oh{�������bx�滭�N�ޣ&�vtm���b��mhZ��V�� h�H3�e3b#�Dy��-�SE�n�Y0ѭ`��l�n�w�K�7\��f�)�aˬ� f�j^^Zؙ�:��U��7nt�2�+T�.�۹:��-G��K��]����2�,���dCPp�f0I�P:�k*'/!�t�0l",�̡t3b��4�c��N 0�b�_1��њE�{���V�yw�Ee�Zwi���a���m%�Ԭ�����r�Y.Υ��Ayld�� ҵ�����8c�f71�J�(D2mCurHe�w��Dp`�pE���=�Y�6��e�f�U�n���*x�x.�
K��#Ux��ӌZ,��,g�3 ��0$��F��ׁ�OU�Bˡ�n<���]�(�صԻ�.�|�������*
���Ա��M��h#d���U7J� �F����)Ӥ�L�+4Em��&iυ!�d�b���=�u,)��W��)2���ۉ��urĐv�4U����U�g�1��o^��l�ۺ���2�2m�b%YF8�c']d��)9����9تm�ܹ�[�a ڬ!S�U4$3.�$VK�p�CXV�).��V�w�[��
G�%e�AY��wIl���^�k�t��&L���Yb�]<���[�Ybꦅm�Y��L-Um4����N���b�l7<*]�0ma`ṃ���bD��l����S#kv�Gs�M�ZȺIm�a<� ׊�A;�'oA��%��m���ʼ�ͷJËMd:��.U�2V�%䢬mą��5:q]�Ѧ�&6�)l��c�s����0Y��n����"���,�������E��e��0BlXV�p	%S�2��(f;F�2u`8t*��E��#uU%ܱE8��2�����I�6Y�ȭ��D�����a�w)���Y��B����I5��-Vé���U�bB��P�G,Ќ�	���UD�N}U:]�?�M�'�'�ҸD7l
��L�d�7���xwsv��܋i+�ѰFX��hv�H�(�����I�Z�lEY��[Z7��)-�8��ڕV�	�U9*�y�6���Q��[��\@e���5�"^�ʼ���[L`U�!����Z��h�kمȽ���R��$Rt.g۫2=�	m�v�3f�ɉ�+U�Q��S
Hދ���"���כ����oٖ(C2�Y
�:�&�����U�TU�%ͨi]I��(%�5�n�[��~A݊V���\�8nʹ���d[��e�ņ���[���wy�e���qާ���ڦ4�52�;�m��y�]��=V>����ْm֐�Z�N\��m�Zw�ZQ��B��c�*=�ք�B�Mȵ�������^�˥t�juzS��j-�A�b��IҎ���t���aZQ%��8�M�Z�s76H��j$.A{+K�1�cF�f��A���P�EYL[4<�ݏK��^�Fy����f:5���O7�E����q�طn� %�Z��lS����P��5�I�hPP�[T��Llhk�Oj�I��:��
ܢs��O�Q�wvƼxFm������Pղ�<��5�V��"E�wl�I�fx��fO��kq��
=F�+#5��j��87
�)��3�)����;��W��� �TC�m��AM�$�vapS�E\��k�Q\,n�X�~-\,l�jV]����9(-u����)Ѵ���Ӗj��ލz��A8w.�40K�աY.�]^�$k�$�#Ϟ���[v�Ҍ��Z���:�d�׭��4'��]Gq���wNZ�n�8��(:��z�H���B�J�$��v���k��w׫&n�Bu�9�� ��"�Wb�S{zH	0� ��F�]An	�)]�t�Ӷ� %6#)�$%����;:4֠qm�)��/q�J6�Nd�H��R)�;�ܦ��qb�b	UB�۔��]�N�ε �g9��k+"�D�m���r�1갚�2l���S��v��'6���h7E�,i�Y��"6,�/�N��E�!��KO�J�U��Z��uwWhkPMsa3D�Sp������&pmeD�--�E�ǰ�'y�Q��@�Ӳ�T�w���`�So>���y�d���E\�̽H@�������Ne�hT���@^�8��uJq=�)GOhfc9{�nZ��yR72��(�4�}SȢI/�6�!cU��hr�×�T�oK�4ɯkfm
a42�FԊ��ܻvT�u@.�)Qn��O(���+1�ge`Z(�ɗB�&N	�ݬs@&۶�Z�0f�Ni.�4���EEJ��L�͢�,�!am�.�6iE�t/qŹ�X��Y����//e����^����zZ6t�ƫŸ�Y�u�F&bv1[@�Xc/2K!����!4K����.�
��cۍ�=j��Q�J���:F!x���j�7UVo�#b��ʖ�\֜��V�sC��"�k
M��d8�I�2��)ǷcM嘄�=���z�+f�Cr̒]2˗��@�PN��7r�����׿�Z���V\���V�Q7U���Ki��E���YUxe�:ҧ.;�LFn��[�M���4Řo�u���F�7d`�f��A�C~6.�B��t>�n� ���Wy�BMk�����p��8r�j3d����,_q��,�4˔&���B8�qa�>~��ŷ�J���9j���ڶ�U��YW+-���V���yn�P*�SS�+*�UUU+,��U*�eX*���Vڶ����mUUJ�U+��-mm�k3*ڭ�"��a�MJ�m��mKAS�V���vR��V)�0�T�[8r������{�b��эe�[���;�k{w�k��1��G�`l���v�8���`T�.޲��n�[k[�L�3ٳS�¾7;��K�(�&��5�S6��c�n"�,f^���ݗ��H�|�>�:.z�14�۰}=v�q�8�eN�ˍBܴ����XVS�k�����Y��Z��U���h:z���2�JƃJ�c�Ԕf�Sn#PJ{{����9��;�cD�L�4�֍٬���֎l����� Yp��p�$�td�,t��`��,I��S����b��ݺ*r�6v�۾o��'��*<v(���{*v�َ���sc^��˃�{pk����یЭ�f-c�������g�g�W\�7WB�
Sʡ�vb��l[[���]�j�Ƹm�/���x�u��5��t��g��g�ƻuQ+���a[�C﫮�k[���ݳ����yX���vy�a,��SSM�\I��A��'�����[<���݃��xNH�V������[{�^��y�������Tua���I��d݄�է��t���>�3���]n���r������oM3��n��z^ht�^N^�5�]�k`�����$Ʒb)!c��0�C]���y7�;yz�u�դV6f��#2!6x�M�����Z��B2$�k���5����'7Y�+�\�l�u�a�h������u��G'c�N�W��Vw#Ƕ�p�L��s�����Vs=l�N�6��PTe���V������Re]I !�	l�{ ��5�ָ�a*��Fc<g�pt��B�ל���+{v�KW,m��T8����'ۭ������y;��n��Z_X5љ��v�=�SV�h�P�AK��3�S��P�cq�$��9��j�`�03y7]�/�ok�`�λ1��R���S�������<���ȼ�[qWHl�m��M�vI(�ל/ջ�۶����_g�P/�w.]��<���]��up� �1�0+�h����b2�R�Ƶ�;��vf�u=ʺB�ݍ���Z�[�����Ɏ�Ϯ��\M�K\!Ko\��W�nNf��Sb�7l'd(�hW:�M�Ba��]%��k�v��ضsM�p��cOq��o������(D�+��09������	=�ֱ���:��{p�I]�0rFy�rG�I[Skv�廎֍��g۝�ۘ%H�#��n{�X�f�Q%^�[KN��V]�q�yk�%-�n�ۜ��m����}�����f+c��Dхn�;s�k�۴vus܉ =��rRu�5��q5�׭�H�����Pӕ��x�n4���BC˧d�p��v�����v�zG��E�Ɖ�;o]5��D1�XV�#!���m�t����Aʢ\��Ktv<�Vz;[�6�r,u�.�l<��ݮn Nz&�Ov4��i��6��K�lJ)��g�{�dtZcv�/��L�������w�[�=u6ѹ�:M�,��K�z��w=8ۡ��x�د-�k��
�}.Q;L����Z����6��L�՛��Y.gF�G3��>��X�c�nNw��m5�t�,^UmA���ff͋1gEծ��#V���H���G��
���=���v���Iֆ��[V��\�7V����v����y�ܽ���Q�v�5]3���܂S�J�m����z��'�l��c[�<z���'V��\�v�ѱ��	�[o#s�m�8�C��Z;B�Ol�*͕���}��X�*�ܲ�2���UT��8��&:G�+f#X���6�ui=:/1���[L��'e�t��
֎r$s1'�wq�����Ο%#�]sv\k��p��xP�]y�)+1AT� ,9�͵��|�n�v����;stޥz�L��; �d�z����In9N{<�g�a�p�ok�[��3�\Mq��/�\/GGj�R9��bym+��&鷃X�d��u�1��:e��@����Z˜�����;S�v���q�8�����=h��.Į=����u�j�\�%��n6NМ����p��uNu��x8מ��U��d\:U��6q�xvɸj�c[]V�D�nŪ34̒��-�mFf�vlS��3��k�[��\>7h!0M�9��Y���ջu��獺��Qd�3��u�ŝ:��RhU&r@����h�����]n�V W��li���"w6��L�qyꝑ��h��j)w5�ukcЂ�p;t=���i�pcd-%�$�c�8����o]/�ʶ�e�+5Z���;�I��8������:b�u�5���m�W���Í3�%7)�:�����P����v|s��:����SZ��k�0֩<c2�L�)�������RsJ�6Wß}c�]���ccR�,�/!���^둽u�7Heiݓ�n��Z�M
@����)��y5�2e���p����㍂m#[rHIf*�l2���H�c�v��s�.�̖��ۣ����<pRJ5���u��\r6�j{)����]6-\0Acqhۇo;�z��x7[P�u��	�),ܘA�cg��A�˪�;�qݗ���͛���:���m�D��:�I��Gk�V�/\Ͷ��7]��+�y�G��3Y�v�ڭ�k��p���]�1�;a��O1׬�8t�aMf����S@��r[t����(������Jn�'O�y�/N��Ip9�������d����\�y͍;hv�2V��4�v�A��%�"����d����E��հ�3M4^4<�%�pe6ۧ��8� -Z��-�-I�,��	'�n'��|���q7pMX�����@�z��B������pv�:]k:�Un�٫����yݠ�����:����q�v\����*��]/cQsu�rsg4m��y�ݸ�I�z��fޜ�g�8f�n���Ul���Rm�+Q�l[�Yo.��G0v�˪�y�q��8L�cX�b�4�X��fv5X�4V�͑\���A&�%��� ��3	M)f�İe �08\7�;I�N��^_c\U�-���s��Lvv䢲v��3Is<Ib��}nГ����>��}�뇫=�����[��!��=�dێ�7S�۪+��֓%�n�Μ��o]k\�j��Eײ+� ��v���ǂx;u&�fKX�Rք�YAfn�Sv�U��m�z.oBb��6r83s�'�2�n��  JXFbl�1�2R�ֻx��W���C�m����ͧt\,b;������v��c�Íbºչ��3pq���OI�ݰdq��z�]�wn�Ȑ�U\X�:�ַ\�t�.�;����X����f�g:�����옎���o#*��j��A6�`٢�X��;`8��Gbd���+��֨�q�W���\j��'@!������7+�Mes3�ᱮ`�g������al-��
6i]���c���p��8n�=g�h��hz����ݲ�qs-�d&�Xt�4��'�Ӊ�u�ᅃ�2�F	\�'��9�'��V��� �o<r1m{vV��e�r�맴�:�Ev֖�D�B�X'���rͱ�\a�i���4��C]���M�gA��q�z����=ۓt��g�Y�;,��M�=���T��U]�V�g)�ܬI����</*�u�ft��e��woo#�LԾ��H%8���.�[�8ĕ+��z��m���w�}Y��9�T��W�0X����L)��j� ��L�����]��s �8;dT*�Ĺ�����l��W/*�.�Ɉ9�n5�r�:�"i�[�퍬ɠ_gn%I:;�^��M9�D�p{S�sv4�Y��KE��w2�k�Vn�K�ۗ+m��s���Kn�݊f�"+�q�tt�������Ρ{�k)�N:�6v���͕0=��\ޜk]�mq.i�4���g۞'.��;A��{kdFf$�@��������޽p�����Xz�rsj�g<�.۵em^�����VȪ�%	mf�C�;r�'�D���l���	��O2z��J�vґs�(��q\f�V:A�7%el��s�m��b�&3��]X�f�S;�b�L��m��e��]Xa��N!m��nn-���V�-�\秱�,�w[c��ۗ��쫸 G�0MMs��	�25w�7����N�#"�ꋦ��@iX)����\��g�Ղ���Jq���y^��*��K{^�v_^������fCvđg��nrs���]mӣ���GPr��\�uYmS=����q��Ur���u��H�0ُ'&�6lg��ym	,qc��Zs]��\7iJ��b�82r��ܝe�V�"��<ua�8{l�2zv���f�h�=mۋ�ng��U��G����NN˗�g��['�>����;e�U�q��h3#v�i�<c,ĸp��D�ϵ��ݹ7!�;�T|v~r}�GH���q�e-��.���v)��nb9�\��c[��$�v������,;��rKv��v��g8���ņ��-۴ v㈧V=�.]	3:jrES\Dx�������}���,�+�E�ב]���<��Z��d�j�y�v.�Ē��S&`������z��p�5���Q��b��l�4U�Z��T!��e��SR0�o<�	�&Χ6�9��ڮ4Hr �R���W+�9�גX���Þ���z���a�u�� Y�[*��lWhy���S[�h:zN92���MaT��Q�x�F瘬�*�k]���<i���:;]��5PP�[��&�vG�K��u��[�8S�q�p*��(�tx�[��LqB�������p�lf��W�[�+5&M�\��yf%��Gsm5u+��"����ݥ:^=Om��퉦TVU-3�j(�dt*��2A��ĠŎcWM�m͛��j�*��
��tW�EUUT*�p*���UQ�T��VsP<n�j(�Q�r�T	m��(T��+k:э6܂n��ێ���.ۮg�K����uǰ�x닣l�:Vjۭ�k���P���j�&bK`�at�u[�枳�w1�K:@9�l��n�붙]����aw�Z�޻L�qP�
8B%h��-��
�e�x�Nwg����gƧ�����gC������Id^ϱ��ִ���'uv�d�����8%�j����qy8�u�c�v�����*��Z6Nf+e6�-$m�];u�4�����9\)��6z;H������-�zn�����qr*aVw-��,�j2�)-,%2B=�X�;Em�Ϟ�y�ً�s���5u��t�x���`�=��k��"��V�뭷�ӭڭ �e�$��I%��Mx�����\f7<u��B�isMJf(�h�A��q�즫���(W���7�D�:�>m��2H�=6.|]F�㞹w����R����pGIԱ�󝞮��X��vv��n5�I{+sj�̴c��:F$ɳ�
��šS��N�b�H�a�rR���6(=P�kj����n'��ϑ���[�n� ^��.2�g��[��������y��/��);Է��Н\.ݒ[�u�N9��]�멻s۳��cvP��;V��b��r�q%Q� V�3�Y�Mc�и�]6ٔ�a�R[%��b5�F��6�x���1�3^��z쉚w9�[�.p�3;F���٤4�f&��B��ѳ9������Bc%������n(�TShVlҔ����%��\FM���cib��ڻ2:�	����p��ږ!����Mn"b�eX�57dq4nr�����W��afVa�3�f�ͥ
��8��4F{Vw��T�e�w��̴rA�Z� lG7��s�,��R�LሎGM=��:;%7��t�ׅ%�gm�ݻ����x�e��\��K틎G�j{n�gB3/�j��fWRQ�##mqcb��1�,��f�S#��e�@U  �3UT((Uj�	�U@j�
�E *��
�H�  P&�P�	� � @�� .�V����m��՚������r)���	nƦ8�3qp{:��c��;��<�Hk�&���id剽s]�:�c&��هX�%8{a;s��:�R�k�GK�ǉ��W�
�uF�A[���������A��Gꓳ�<x��l�d�3MV�ԁfyY��A�v*Ù��^�-�+˔��5ћL;YRČ�f\�q͸�ɺգ�{��h5F����`�xƶ/Z�Vb�-�ƒ�T� ��@����?9.�&KD�\��+j(��N���>��Rۂ+�����ˁ6"o·0���h�������l���*�%���[9���u��x�Z3��Mkr�p[�`]�T���Z���n�d�
K����e%J��M���am5̴]��Q��o���=ƴ�I����wk�/�҃����]Y�',K������Xk��MQn�ǭ�Kڛ�/�uu�f����^޻pg7.����Q����{�RJ�N������72P���Kz�S��W^�@�0JAR�
)���5(��b�g+��-8J����zY���{7x�Y�:$�ly�,:ڧ��>���i�}9ME�)K���ISt�mS���#�*��;n,�6����b� \��3]���91MѢj��B-����i�Rg�]��9fڳPZt_cm�ow���3k�	����1Hcئ���2'�k���%�A"�L�fn\��&��Z�^�/pn�Z\��%�1��c�0��N#�-��J�l���1����0�\t��J�N�mt�qg39Ͳ���q�nW����f]n��^��vƬ�-p<�eoe�	v��3�E�5j�L�{ԍw^�2tj��
��K�-����V���hݎ��_�x�]�Ց��9��ۣ�}�ߴ��L�s3\��ɹ�F"Jwa$�XhR-�SLf��Y�2>�vW��w;��U6L�뺊��ں/_1"�w�U�ؙ����Fi;��!�J_&(Mm �&��I�u��m��7l_X�/g���������GGn^Ұt�zb�� ��O��]G4�ү�&sqt����Zvv�nΣJ���9�*8-`6,0r%=�g�rA�[�5��؇���1��k�q��A� ��//P6�*����jM{-��y��b/L&����Id���tl(NXO��t�n�WM��N���W���fU��.ܖ{���\m�+f�Wr��u�"�~u�bf�J�I鴘�;�t���ٽg? ����a���#���mX���#�����W��	����9����L���*Z]F��S�7l=��t�ûc��F�G�������ka@�^�1f����c�0�4�e�Z-�.��l��.O�o������l�-���m��Ѕ��~�Zj�(A���iq7w�*�ݺ}W葼=&O l���&J2����
/���e��{p���|�yz���Ӵ�G+p:�x������@���Cl:����t5ٷ.�)��g[��l�3�K��RD9n;Fk'b��/<@k�%+�\��`�N�`�U����^�ܔٮ.����#P��X��\�qt;�u^
>��k�=��]ɢ�mhk��
h�Fx'�t�>�g�I(���ʏ�%�rŽE)*(+�d��l��|<U��Xʇ�8����:5�Q���L�%0�gty}:ٸ�A�X)(��!XL��,>Ԛ[=Ѫx���̼�xg��eδ	՜=l����\�H��P:�����{O��]Cb�t���yX�v�V���W:7��|���)���ƶ��pW����a7].�VQ��m1�e����-���צ�U�vCr�Y�F��3w�do�xX��}�Tf$*l�IÔm�&oZ�e�lc��w�g�^�GݧǕE���r!�[�=4y��^���������$��{���o&AJ�Hܟ�ܻ`��v�[�ۊ^��Hx�R�����ծڌ�M�.V�i�q��y���~�՘��G�m�R��
���e�7Y^~t01�jNé�:��ف�m��j̓+(�&��`�k4�z�Z!�;}~��}Ǳ��C���)%=Z �&��w���̠�./8�)G�^��ykp? 8�+(�.�%:���s�K�~���$��~㣸X{��V�^�����bB;�����HG�<��E
Ϛ��Т2�Rc�.����� 3֣�]:���&��ڗ��+K��������"[�ʛ2
�٪�S���h��&KI�:%��#QK-������*�V��S*�M��63+uXĻ������M`��#�H#5]��}�ێd����\-Ãk���f*.��k+�yՒ�>3�'kC0��a���&�)����f���tў���W���p��za^��y^��.x#gs;Ζ�ǎ�7,�Oa=y��U�댏nK̈I��As�:���]�Y�7;�]��8�vĨ��G]lVh�냋%��ڟc-E��g����l�]�.�V2��xs��cDq�s��� ��K��"R�b:Saxֻs��N��7k`��p�6y1m2q]�U�X�ݱ7�|��
؞{gSH����AӜW`�ۍBCm�%�^n�v��;H��j�omziN�Z��s��Q��T��f�bG8Ǉe�v��M�Qmb川&�9,�=�x&#I���@��bX���M�͑�v��|r��{��T5����u�"N��3ά�$ 7�;i�k�B&�U�L6�I��DZ�c����MeG�7ӽh� �����|��k�;�20��hq��~�nӗ�����{��8LJ�'J�m3�n��D$�(Y���6�-��"���Z����LY�	�S��
���[���v�u��ް�"��S�Bm��;���*�Ol��p~��J�Vc�N�0p&uF�\�u�΢�Ùy�t�W�"�_X�ч��<Ͻ��iL�n�*fm���nYMJԚl[�kA�F��ؤl\ۗD�WQ%�@����T���bX�/��}��{�-U���kiT���犾K�m7���}�]�@�{u����d���{��o-�nA�7�y�������j�P^�&�љ��ǜ�&�����(����'F{7�MQ֣*YsXu*���u�A��y�������^k8״�Z��9�"Rn<�❯7c[gD�gN^-i��uN!�5�}Nr�K�<�/���	�*���<}��[X�󓔻9�(�}��!`1"E9q���^��1n���g}0��c�X��Z��^�|�*k^�f�V
�0-�<wɦ�<���b�
�;@��"1
D�tM��F�f���>x"��$)y�b�xo�9N�>f��b볜�/��,� ��1c�x�۴�5=�]�n�S�p���]��ּ�<=GJv�֐ȑÙ^8*�<6㱊w-e�:5�-����V4�;�>ȝ�x��3E�r�ۜ���!/wz�<Ku�ro�J�HѤ�l"�b>�����`wv�*1��y�װ����ֺ��V���;�ƎSX��~u��cAX�{���iAh_�JD�%��m�x ���C6��j���5�yތ�	J�u\���,���{�.��t}�}�+���\h���زJͩ��$�;���j.q)//��yѲ�n$������gV�W,]�I'b��ݦr�{�\,�H���m&w�~}��A����}%1�s��Y��5�����LR�n��
l� 1�*��t��{�Z�d�v9Q�0�B�B	��)�n����	E|=�C���sF,k�A^�t>˳;o+V1��4$��Z5�]��)�S���U��H��F�Q���R�)z��\��fC;��nf��rZ�eƱ%�Ս��-n?n�ߋyk|��Kun��ז�%�az�I�԰���oM�&�kN��j�"�k{/��aA��b5^��
\Y�U"�M�2�2�����:,܈��󠽎��3ݪ�WD�|���m�{4�|˺:/��#+w���ڪp�C� CJ�(��Vg ��[��ӻO����z��S��;g]��y^k����k�<Kx��]��n	m&RP7$[��Z5���K �3+�i�H�Z���O����������MR9��ҏ���]X�����q�;�������@��a�#��"���
��n�Y'׃����oЌ|6�`�*���٘�@%�D���`V�����)�@ 	�E1������{<�]��fl�̾٤�*:$�4嗙��U ��{@fK��m�s�&��H|�{Qk<�:_;�w�i���V�+(�by;F2U�'WVpܬ( ^��Ƶ��%�ix�\�m�Kl���V�DD:༉#J$��.U�m׷g�R�V���������5-��ZF3э�b��Z4]}M
b�"�k1�A*\���\��e�3��^M@���l����ck쭺��smn�����b�>����\�Dӧ@ ��V�[]�lϑ�}l2�J��2vo+��� ף������
J��c��@�� �'T��z�r�'��2>"{bW��G~�� o���.�Xi��6�3�5��7���`�}dAm5�J��mi��.��{�hi��U�����԰k(v�r7��1,i���w�Z
WZ��3�%b�����cU&�����p9;�Lr�yK50�x���7��׻�{��j莻�
���V��J��z��%���n���������"e�i�Շ6��h9*��{��0`ݩ�2l]n������/���t��Y^L�D�n�Kʰ�[�i3c���l#s��\B�7bb9y�뗺tr�9s��wF�[ss9��8B�&������.��ݭ����$��G6��7�i�v5�;�\�3�K(�����z^h0�z��r.o���}�!Ls��<<u�6(m�����*�Rv띦8琷�9[��9��ڶ���gpy˝K]X�:X��65�|{��������չ�p���f�����Y�O��;�~�������MM�}�qb�4����m,<���K��vB�x7�6��J�\�Q�}�a���!�S0�4���ܦ!q���swy5���{O�[&�F�;��i6Z��Ɍ�9{ϖ)X6��2�����-��@�x��ŧC�������2��	�
e&����x���j���%��}*ܲ��'
m��v
3^��9W�/m����ޠSCۯ��e.�a�e�L2K)�a��`���_��r�3~�^�Ɇ{3�;	'��%�V\$��n�	x���gt��X�f�:��ףu�ۛ�����'\�%X�v�y�\<�m�jӅ���;ר�n�m�??�?ci�.XG�Vy������R�������=E{}~�@�����X�4E^#��$��TE0Ln��ۣ#�V:����g��r�����
,�c�D�j�Z���mUަ�]�QK��"���M%�"�g������vV�M7o]��7Co��:Ä��Mu�h&E���}r�U3n���\�3�=Vu����f�re�&�Vl42IM2��Y���w�R�W��ٻP�{�:-a���[�dXU9;���Ht����]��{nY]�Fݔ���ai�\���l[7F�����N����VE:���]KF�b��۷��z�o1�:�l�E��j�E��v����`�G�m��|<o0�x����D�onHħ)ֲ��E�2�rT#���v��t��in���ؚ�F�3N�Q9��8�֣����麳r�mڎ:�6�sm�v$z���O6j.��[����e���:���m��^��Ou�]1��w*l�qTh���YM���W����0�t(��!0)4`� �ޯu���hG��+���s�M@ׇ��!H\8����Ȉ}�.�J��M�@��E3wh� ����f��v+�{T��{
�R��
�v�JӗW�p3X����^��1��v��g5>�$�Y\�|���׵�ڼ�a'�>e�;OV�59}܅�Ucs���Ε�*����a⮵O�(n���eK����c�k�)��:E-a�o�yi7�.8���=�)�J�9zQT��y/�q����w��D�3��1�wVn���ʛ.¾���zEvj8�':����җ��0(e⠨vpl&vQ��c*�kH�+�ʹ�y�+A�1�'M��WH�Hڡ��������ݴ����+~�C+^��a-ǒ7��E���[A],Е�6��6wmK��2��y#^��wӥ)s	�Ԅ���+��pݦJ�J�ۭc3!X�ӗ�)wg��m.�]�0X[��tYV;���:5Vࠖ�]w�-��݃fh�Sz�5c*�wS��h�^�̛����C3�]�|���.�oz�a&�m�V��'�!y��9�����݋��.�����y�mZ:��ʣ��ۇ���`�7@��ͩ˞�6/ms��#���W���$D���4��ڍ�p��w�rB˵H��ͧ*�:�t�en�m�,Cz�O��4&M�|�8���vi���a���On�㝽�5��S�Z�\ۢS�d����0���婜U�Δ���1[ �|��_Gg&6nͭ��+˥Y�w{�W f�lW��^�L[y�d/��?s�ͬ�CGS��͛K3���;�Ѿ͋��N}C��jqQ��.?����a"(�GU�g��s��ue����ƅ����Ļʌ�������BF��<�~޻�lN�����H��m"�,^���}C!�g���qn��XE��u�-��\s�o/�H��GQ�]6�$���|�C.����¶�L�t��~��2��XѶt\����gV�vm�RX�^�����Z7lJ�>H��7�>O�E`��xm;�X�o8��>��q��-m��ٴt�]���<��J�n{L��%8�����t]1c�P+�����*�Ar�z3�
|�������D�Yh{;�vo��P�A���c8d��a�"48{}6�#c�n�t�����8$3�(��8�MV*(�>>�z-	��s1p�Xl���� S�	2��$�q���ݖvͯ �8�V��~o�~b�Ө�a�Z��-y�=���e���	��F?� ��M6[7�^]n��cB��仐!�{mB�z�BV�ż���ou��8>�;7<Y�H��2�#��ݾ�ժX��7b��wV��;�l����ge�o�;�Q���x��<�^�D��0y"t���o_6&/�u�;��3�y4��_{����Z���+�
]�)����e�G>a^<Z-�QU;�}���3�*P�>�xI7�b]?"J��dY���퓕-���jxu��2]����w�[9��n��2� �拶�u�f�vж�#��9 [������$v��{>v���9j��4V�F!�U�0�Z�ۦv�`ʙ�llY���z��/.'g���:! ���S�t���mq�Y0c��������ŭy!���^���b@牘�&x�����JdLV��b�ΤF����Q��w���d�����MH���9��i� g�c����?Z�f�5tݮw�@�

�V�E��jm=�Ŗ3����K������4n]�A	f��7�����(��4�  ީvӬ�r��_��a�������wo;��q9��],�r�w7��r�->aq�n�� ʹk��\'Mt�qGok錩���Tބ��	� %��]����� ��D���Q۠o�^�*��X��fC|+�����-<��I	�C)e�+�����8���烑�2qqk��ʧ:��.6M�*E��h���b[R�t�9V]�wkb|	n�x��h޺M;��ۮh-��^X9�7K�f��8�eѮw4��ݭ����1a�t�Q�n:PM�O��/��N�՝3�K
�l�񘱩��*�.�a	x;(�\���r��zJ�4�v�Ms��s���6�x�:���7]�u\Q�ƺ��n���Ƈ^j/m]7��C��^��m�r��Ǯ�y4�Ɖ���M�5�	�-��*FlJOv�R|�����q�mtf�Q&͎�������!���X�\�Xkv��g���W�k���Z�t��[�+��Qwy�Vlm���m���Z�+��~��R�35�"�u�wH�V3���ͣA�M�ږ���P+�܇���^������322��E�k�� ��:Зc.&rm�(S}c��E�@a��5T�3��?k�]���l���o�&c8,?�=�u�@qn*O��WJ�٭6�n��b�>����`��)
2� �,�h�5.{t�58��j6/��Z�Tv�B�;�e�i�F��NA�CÌ@�
���������nU���o��MR���I��ְkQ��[�|am�K6Ў@����wc;�&��%JR�����;�~�ε=~zs�n��&h��R��G�C8u�i��OwZ�ۂ߽6� ���;�#@�e �Ɇ�m*�,sb2�/�����=�{|�1nS�|~ǚ�c�~�N2��)�ӧ�.��(�{�x��R�u�Z���pBm����ĝ;�ҕ̬���b�J,������y��.�y	^q�iVM��zw4@��/h"�]TQI�%1��KZ�{2ô��+޹��|4��*�J���l�(a[Z�����K��.�r��֕E������'�O�X#ڇ�-"����}.�2l�<�OӶ<y�x�	P�bY���:�Y��y��w�Qw������H �S�i'[�1�e��ߔ�Q�D�/]Xev͠�����]w�]��V�-y�V�/Q��[��Ѧ�l'N�1�]�����3q�d*n]v�v���f�q�۶�ׯ=�˙����o��~l�wy��
.�6���m�鉈��{Oe)�����=����e�{�.Ln*6����av�ttρ���'�=�*�]�Z�wN��ӈ=�mEqW�|�]�.g��aǤ^���'��ө���H�J�5K��kВ*F�>�=�<P�.%ʽ��$G�l�S��lE�fg��+��e��b��
��Kڼ��w��1I?Uo���Z���S5������2X�~�O��T6�>KR���z�VzM�Y¢x���
ekΞ�����gT���,	��*I��om�(���-�򭔽��Y�f��-�SW����X���kAV볭�hۥ:_c���񅤡�H m�TM�M�i�Yn�k6�ygնM"80mPX�RG�+/���Rf��Б�m��w��9�s���e���n�ƓE�D��X�@��⻝�*R���sw��/g��d;G0�8�����a�p�����IO;�=����My �9lj��W�QB���.��Wf�^&���U��A
%�E�m���{�q�U�� z���,�\k�b���g}������B������y8�w/`"�Q?�M�6� %Y���k�~����uIZ1����ג{
�
=,�.�潴�Sxv�>q�fe�~ߗ��I�E�ڣ��;}!�آ�u��^��܈�4
�&@����4��yn9�^y�n�Rߟٝ�=��h�Q���%��-q�#�W*a7�;��x�2B-^c{�"r2�K�4�JOY��*����'w�ݼmާ�:ʴx:� �t 
c2�]����>�i���k����O/� PW&���*����vXp^�)خP��VT}V!|�_�S�74l%��p�q<�V�8ٴ�U����;W1q�����#۱9y�.W]��J�ǰ�:�z��뇧XSQh��s�̝C�2�iWAN�"��U�j�:Lht�h�0:��&�K�Uǒ�j�Y�����Ju�۫uZ(�Z9����q�o#	2}���փ��̱�;�3�lHEӦ�vnb���tf�r���=��A���Ļ�Վ�;�q�ez��L���B��'53�B�K���uE�0�#�S�v�0fΥ�/�
�m�8.�����9�u{Q�Nb�"��:]����
-{����P����I�qZR�@��\��(P�M�xg-~&�}mt�o�h�.ס����y�+�+6��,��qj8�<"�jL�Dd���d����gfguC�sF�y������p��ϔ�syV���I�r��aZ�/�c�!u޷m�Il�����K�cN9��	��$�WMv�����e��8&�����K�ր��U��-P��vzq:��H��\S3@Kv���@4�b&���X��ݜ��u�:�FOkr��!ƍ���v�u���Fu�:�mZt"�7��;F���GKmtYR �ʴ[hc�ny�9�s�%6����e�Z����fXSn���ʮ�<�=7;C�'Wmv�/���G�Ya8uC�aջm�0�Z.m��l�M���۱�"75\�S)�����݌�ƿ:���]�g܌
�W΀���J���]����������c���
(N(��nL7�6�G��{���&{T6�$R [f��9�o�b�IB�]*����W������C�H�:j�h�m�A����K����wxn��
��z_V���j��8t�2��䥍��Ty�ocU����x	򱉄`DƓ�T-�r#]~3ww�Fm/3��ٝo�&����N��A~ʜw�Br]f�
��g�^�ޜR�z��h�J��A$�E�Ω��b���~�k��o.c{&�i���ǚ.5�H6�9��-����.�����*�]@R����}��dq���/���wg{5ӱ����	�G����6��s�v�<�8�A{�����=�����zlr��Qe�ז�6�Ml��P��!�P���ؔ@�Zmq]���x�e�+��$Be��h������-In�WDc��.������r�;�J������U)Q.���*:��r� NޣIɋ�c7:c�8k�P]��C�	or�l�g'CN�J���65٧���A��{Is�`��"��X��]�U��r��`�5��KS(��LUSA2m6�,�3C�ygw|��������s��oA̹
=<�G��S�S�M���C�AT��P���^�Mw�O����s���Xȼf�� �����qQ"wpYOn���m��M֫��*ZT�`�ڣ�J�-��֥��\�h�}n�U�����]������N��������:r�Ƒz]�����`=��-��[
!$�$�X���s5^;fl  wM��]���9-��W<U� 
�L�h��^qG�b�[F�nZ�lwyT�T��*g����'en7ls�ϥ�z��1�"lU&�7M�	n����|��G���o�J����|!�`}k"�$3Wi�M;z��m�)�#���23<�~`���t	� ���Q�ZL˫!$�z���S֗��n�h��[r��C���������.��u��sy�ŵ��]s�Sr_^�'[�` p�u�0|�W���}u�ed��kT���� �ukG��{���>�SW�y�[�#�(�� ��%��mnP�dB'���9�Iv��������%
A�H�>ce��m�\�5���In�N�r��nX�_��7�(��Ϡ�PfEH�[���x����3�2^s^X�%���\Wf^�����Me�д]�j�yj#�Y�$3mi¨�PP�(����g!GMb
���F�.�e�v�<C�l�t����n�]0�-B�d���Oe��.��v��\�.�,m�W�-�5��k�t�뤶�dJ�(�Yv�(����wT�*���D��2S>�knD$Q�]fq���2j״[�{3Ֆka�Ü��0q%���;3*���\��4,Z�ft���ADP@�N20�F&H!�s�nc�aC�n�y�뮕�ڱ0���U�e|�o�N�;�<�-��P�U�$�U2�h2�Pf=iI���u�	h7�B���h�G��]}[��<�O�guk]W���>]�!��{Pެ�tvQ>��'Yr9�7�U�,Y���E����0=���=w��2�p<�p^a\���72�`h:��'{��ea�Ƭ�[A�&�E�2�mՅv�;8L�3t^��e��<q�#���m�W}cz�LwL���W��[�]�;����X���n3I)��2s�n��rk�=�Yu&�h#l�;#`g\�Ġa��.��A�Ɵk Q	�����^>acv�����G#;��M]�AJ�s)�7���B$ˢ�4���p4cN;!��h�'����K�a�nf�p��,���~�$�M���3��Y�p�W&�m<�0!\�I�tz`%`&� )�pf ���ŶB�P�Jm̂�w���p�*�<&]k��<�µvՠD��g����*�ߗӨύ|���[t�-��~�_˼p�K�5,r����u��Nڗk��k����rȃ�{��1_f�&��&W�ޅثܮd���0��HIԽ(,:�kְ���U�;�{=[�Jt|�-HF��^���A3�W7O��#a�+a���J0/���[���޾�QT��eRFԽ�֊|�;��p�:Tv-�ٻs�ӷg��^˼P�ϱ3�l=�+����gut�n����=n�}����� ��e,ʵΎ��ѢeŊth����m�:*���]ƹ�Xx�$����r�X�Z�Jn��u�����Lm�m���<��y�&S��L?SKם�:g��f�Y'_d,Ӈ@�Ca����B{������T��*֡���,~od���0�����woWN�F��n�j�7d}N��4� Aq��Rfӗ9���:��GsMp�m��gM�� ��q|h�J*ꋞұ�C�T,s����v,y�����9�X6$�����W���f�ϻwq��4F�k5j�ĩN�c�;�ՍyW�ɝ����s�Xw �(��Y��\�Q[j$v�:��{*h��ݔ�k��o_i�L�P!I�����G5�k{4]�]��s&f�ݐa���
WТqt����Җ�avlQ �®PY�Qt#m��I���^���j�-w��9c���f�h-\��P�Z��0y8���F�,;s�U���rk���e��W����<2u:T(�����e5m�J��R��rܩ/���p(Yԛ��sDγ���P��J���`pqz�n(��|�3�eAl5�K�w�l��v��ع�l*�f�I��m�5/l>����-9_�k �2��N���K�}w�C�M�����<r0^J�ѻ{|�ѠG3��²���z��d�=�?T�k��r;����dX������]6�l���J�4���ر���V��@�VnsX�0���m�K�&3����թG��l���;�f8l0q�\�O'5NB�3X؜mFƎ�Kk��;n' Y�+������E�1t��X՛��F�����.�0�[�'d=�%O�i�e��L7�N��WmH��ƵI�m2)�E��ҝ���y]G'��qup�/S�4�xeznB�����'T����:䛳-��s)X�Z� 4�iXx��u�m[v�V��=��m,��jK��	��3JJhE&h�(�Y.âP4���������t����+&��n]ۉ6{7s>��p�xu�␍�:gg�G[�\�{z7`�T���m��5Zx��(�3Mm������Z��u��g���w�W�m�\���rt!���=>�z}��̞)�}M��ԝ��������`��\���6�U�T��:��,���T���p�76\��ݨ�ݞqS�B5I-FN��!<��l�����5��n��G+�i�<9��v�������wt[`�B0�+h�6f��Ұ-�1�t@�a�)��!��fVj��݀_P8o�t��ݞ#�}�M���v{NI�75ݳ�V�P�{��]���.�9��i2ט�q˦R݆"��Z霩-�v�=���R�۶��=���,;s�9�w]��B����<��ۺ.N���-�����Q�n,u�w]�Z(��2@�o^���S�E�)Z��o�I���1�S�v�]�8W���lN){rOs�n�=�0Fci�5���V؁����h��Z�\lݒv�7))�t�4I�<2�Vڃ���g�l���!�l��J���n��B�k��Z���6㳸燣��M���hy��S�iHm�X\�0f(.Ͱ�:�73]�Y�l�S�ks⪆֣L��5�K��-Z��Z��c� ���\@�ݤ%�..�ЀA��k-!����t���c���:Wʼ����	b����b��Ҽ��qܜ��ԶĪElY��.N�)v�8h�ɳp]�Wd�6�mg�r��9�����y�6Ƭm֨�4*D�[�:��]�j.7a[CvC�l����;���r|�}���
qښ�g'L���n��61N�Çp�'��r;��tM�ݽ�Rx��օ�v�����L�&25p�n-h��Bk��ǖ�8�Ql��nm�����Ӑg�pDRŹ�I,t�%�ѹ���C��#/\3���Y..� �������3n�z����3p�ENݨ8:�.S2oχ�1�K�绵���/�/B�S�̹���4C��E{��Kŏ�]�ծzᣭW��8[e��M��6,�=��E�G<v�:/[��Z�⾷��⡠�;�z��˹p^h]���>���l(S��� Pi�H%�\�@ b��pk�6=��J�Z�1(=�dB��4�V{�17W���e�A�|���d����_V�k=� ���|Ǻ�ݡ�����pU�Ϳ@��9��r��=#��S{��IPH�H��e��)u�߅��L�Kxx��Eߧ�*׮���}1àiD�޼沇���G�o�A{�|���*a�B�8�q)Q��C\6�x��]{qk�ny�9�ηE2�ɐ�{>w]m͖R):�ǭ��G݋V����h�JJt�fv�b+��4�K�z��[wR�rn;r���x� ��댄Sd�E�[m!Ww��n1^˾;��]��l�Z�Lo�ژ�T�2S�����`R���՝vv��B�V�4�{n�\����W=N�Է�4��Vk�M�h�ץ<��ۻ�, �e�}됱/Z�Ҽc�Ko%kG�G��p��:�t�m��Q,&ǂM%r�l�ɱ����e��1>�U�����ݴ�Z9˽tz5�`:n;��+�+�v%�]��m��i��M}������W��:�k��F(o����c�n{<3;��;� W��S��ZN���ߝ��L�ʦ�L��>�ĩ����Pe���E[��2����W�]�[���O3�㷺vs`20vb�`��S�@cP�Z�"���皕��8�IYۛ��<n��mc6'ugtqC� tE �h II����|3 ��_CSS�m+c},Ƭ��@F���MXw�P�b����o+�KJ�G�±�V֩�E",��m$�cQ:�k�G��툼��^���f�'1;��ǦPX�@�뻶�@���ޥ�>�5����	d�HT�M!Sb+�޻⛻�/�g��G0T/~�c�{w����RՔ���*�Z��(�PQ�)�|k/]�w����5+�k3)�V�]`X�L}u�'�(���o�<;]b�4���9�&����<d��a=={x�L�K��Ht��F��3�D���U)kK;ϼ�٤K���U��n������ڡ�yr	r�/-�P流�;����a�TL`�����(��,�v��Dی��<:"�[I��GVk��FOu�1��Y���7t����GԺ]�W�/I�+p�LӅY_9��M=d��l:4Ri:c-��<�v�Ͷ���Vw�zİ6˧����7>`M���h%q���m�7��d^��齞�X��s��ʭ�92�Ej�/��$�f����P��g=]r�҈�(
`��"�c��lF�2v���6����nRT��}%{]�i`J]�΅v�]$!TmK=7������������
��,�`��:0���i	e���߸��M�O��=G�]��}��ȝ��������pҕ�)���[�u<�RX��SoO��WX�sm��{�t����]Ū��u�1+��p�*�v�u\:��o�F�k�{j�F��c捬�iw	$Ü��R������+aG�����Μ����.�x/Q�zgM��9P�q+-WJG�{�m�%Wg6�qrT$vh�(�����2�e��ݲ��e�x������c�D�~l�&���k.�2��9��*�z>=3%�Iq��Aw��n�ߏ��9�=ĳ�Lp��2�r�yh��g#3Fg6k��h�u��!���(�{��4�"-�n<�s��z��3���1V��/���{]ys�CM�L!������m�H������G�0�F��8t���j�5x>ǯ��o+��W����j^�δ��O���j�+�����y3ʴ����J�
�4D��(�Ѧ[s�'u����i�5�n�U�.]�"�&�i�}��T�.�� �F&�/��7&ꧨ���`Bm#Ծ4��2�9���p=��ջ;\K�~Uk@rk���jc��h�ő���v�{6�����zu��%`�Xq4��M���V�e�-��������^�@rmSy�Qum9��^��Kϡ�����9��Kbom�蕓����Ai[ '�6(Ӿ�v\��6d�/v��%)d�n:�wٽ���Y�9���uΎlfN���؎o�����Iw��݇l�5��4`��E��t5���,v��,���z�샺v�N�î�D0M��\-��<�ܼ���u/1����'���k�Sn�5��y;d�����
Ƹ�����4c��\�2Ǒ��j����u�Y�@���g�A6�v:����zx�ysbnԛn81
1R�B�lF3CrnF���',ruV�h���&�4=\��p\,Ul҄����5T�s*Kj)6�9[f&�F�nX��q���U�O�?���������-�S+ŷ�}�0ժH$��qd�����������N�v(��?twIq �a[Qس�j���߲3���W}�ɚ'P�>�J�+�k�C�e��3�E��O��)�^b��&c�<��,�) E�i��"��~�M���/�=��>�T�#�v�Sj��	*#~NP�g�B�Ru���n<A���v����	0S-�h����Feeh~��n��nf�i�mQ�}p!��V�)�k�����w�Pݼ9�f�n���n<1�.�p�����P�t�b�"+�4`��������c-�XZ=���op��4��/&�z�r.����b�й/��J��
���k7{��"�,��iFJDD�����L1sv�]����S�����>��n��>�0A$���'�G~̄��ɿ%�'��MEQ�3V�^\���\ݎ�Z��s�[�gL	T����)l��At	L�xnK����s�b��pyo�զwE`ɾ�U�i�d���u�����S��(�18���ט.4d׽U����Fn:�sRc�.�9��4e���qT{��t�u[�z����c�n���f��j�XG�,U��y�=[+��*&�m)�[�K�o��K>F�"EJ�A���������}�h�tU׍h��6����`{�ןCW/x���E7��z�b�m�]v��dZ�d*T��[�;q��$W��`��/�æ�y9ߨ��Iu����1\�,k.�� S8o�+}�30y���(A��I�):_hH� ���y�uR���Z4[پN���Q�x�{ҵ�j�Q���}��'=�f��
����GC��,<���m���=v뜗�W��K9R�y�jxՏdd, &5"Q�w���fUːu��#YT�C4��;�ӫ��=�9ܫ�l ד������n��^��6;�m�� �D�1A��iK�I�j��~E�w\쾈�_����a9*Ǵ8�'���(�y�^Y�o��j��^˧�Y^u� �Dj�Yl*��)�o���%~s�`�5��J};�i�{{���QyA�!J	RT�e�x��m@f#W������5	Ma�c�E�w�k`a�CO�wZ=��/μ<�n{uv+�9����6�FUe޻���08�,Kb2���=��޹h�|:��Oq�F��t��Sk$R]����ڄ˻~W��y��H=�y�������R?��[l^x�*���a�	$�Fq]k�bo���Q/t��5*G�_I�&�:�^>}�@V��v�Y����4@Sv�琼D�ugʈ��E��!.J�;h�:w-���D�i��V���~�=oz��Rn���� �-���)P;�o��ʩ��W6�g�A�Z���D�{4[�����	|S-R�cl��egC~���q݋Ygn�6�7�|e��[H�y"��9^%���f�~��Մ�V�$a�H_����e�,��t
u��KN�=ٚm�SJ�m�Z��.f���F��n�S(��R�6�9/-���ɸ���2���ИE��I,�
��f,������,�A�gW�M��t.�ކXK9a��v�d��<�h-��Z��v����m���1�~JW��s}��]�d�p�.B����L�v(�O2q�t�����	�{��]���%��{��ɾ����¨�H] �l �ML�;��L),��%N��M����\9�Ov҃��SVj�3A��v��u�ې
�������kA�.Ro���X�ۉ/33��R�����\����y�p���dk��u͸���Ln�����<
�o�tJ��qɳf0�^��W�F�#1�w��qQW��ѻY��$+*Ǐ/�� �EI0��oN�
�9����{<F{~_v���J��W:�o��,�7K����y{���Ϛ�ʺi�|�.4���9fP��TK%��i��v���Z�{RA����&rbd�L���ei�(B���r�dwW�9���y�� E�:�r�A>�D��ۉG������_�}zv�n?_�`��N蘢���
�2�2��E����
7jϕP�����{�X���j&��6�o�S�71I�a��{I���ŝU۫�iOm�DZ�ǝ_�,���I�-���J�}hZ���{lc5^*�F�Qw	�5��7^�	ڂ���\�;�����kFp+MĞ�����ۤ���۵�Tڹ*�I��MSS5V���,9�����ӹ�6ǁ�ӗ�7M��7T�R��5�+n9:���à��)�f3T�ln���<���o]����q�f�%��k��KYtULZl�JFX\�pH\���΍����Dt�z��;��6����u$�L�s�1[\�;�j�2�Zcs>��N�s��cj���y��˕w;��vH�]W[�Wg�""뫉�(b��.޴�Snι��.��K��2l�k�	�wV+o3hF��ֶ݋�a��a����?�(�~���ﴽeg��z�z(�w�
���v���Ff/l��[<E�"�����9��hJ0A%H����3n��=Q��WU�
M-�<���.�Bb��X�Ѭ���u�;Oh:�����}L:�GȠW�2�T�l�V��h�z��LP�uw�!D��Jk�Þ�r��$�ۥ���+A�k�-o`w�>�a\45%Ȑ��Z�i���Q��:u�pfZ�mgh� J�@���=w�OU�Y�oϛ�2�X0>��o16]D��D�f�y�}���"H�$�G��p�y[�5��bUJ�8��xz7kU'+��f�!wzwm��Y��f}r����u�=>�S%m/9.n�y�n�����n�cY�����nL��z��v�N}q!�D����εT�߯�ьq��c�U-���ڊ_���y1���Y)�u�����R���%g��$��<��F��T�Kn������ϻڇk˯!r}���D$���u���s�W�V�c*X��峒�1P}a�����wtoc�D��::�F^�&jN�%��M�����Pӆ���S�YW��Ц;ʦ�l�b�i^�J�+�w�j�ϒN�F\���ɉ�8�S�����Ef�q��,���Y�5�[��� ��{���v�b�Y�����v$�^��E���d���{ؽ#���Z~*�n���m<�T���r�M^��qzJAy��a�����ompy4�D�8Z�$ ��pE"�ɗ�ɍM���X(��
�b����w�z�K��$������H��UtW�U��ʰu����U���ʖ�P |�h �nK�FYV������.e��۫�Im��]Z��r��Z��J�Eչ���-����g�{ʀO;>ʓ�zz^���OD4+��wJ�)���H��ñɁ$6Տz�8�H�hi���/V�[��o�OR��8R�h��4�=�S ��^����xE��{+�iDz��V�0�|��9Bj�(��#q4��}�0x��|7ϾĎ/�|W�����G�Yd�y�JbS$��7�5L�h2��(D }��ϱ]#��CC֨3�u�{��{U��
��~����������)�|ח�c��;�����K�Z�N�W��1Dx�\�x ��5-�������3%dǳ��V��j��yc����E8�u��h�/��Pܺ.�q�ZVH��5�3f��'��<x˫{C4�w�K:IV;B���������Tv �t<�zZ��y�΂���U�ŽfYw%Ù�oӽ�Jj�M�b9�t�E�&WKn >|���k�R#sp��������V'Y���vw�"^��9Xh�8��|���:ݼ����oT*�ۣ�2<������5S�w6�{zD�;O>���MN���g;b�[��=����~�_�U��BF��m��G����]]F�9ټ�;3�4�m�h���wE���]퐓��i�X<��C �ݲ�-%�D����vE�]�p�d���Fq�R�׮�η�VS탟u�V^��Lv���3d{�����E��Ͱ⩲k�R�(`�8nu,�g!����R�HP֓g{��r	}��%�r�s��{��V1C����0/r!��f1���s�ff<�L�]e�( l�� gc��l�vK�[Wܭw1U�z�7��u��+���m��������B�b�v��å�Ɠ��}��t�{� -��j���޼u΃�ګ�$]�Le>��F5�{��W`���+i%:�t�u��y��(n��qwI����K[�	�B�O>������R�4{����=�{�%�sN�~cG���3O9�pf�8i��*П}���c�h0֐!?���5�;?���W�F��Rە�#����4�9����GmggmX��I$h�ڡ��}+�Ͻ�|A(�"�Ρ��F��=����)i�a��4};��m�Q����S8,��1,��Z�Fd"I$d���ȵ�R�Mmǒ`��c��̞-&B:D�����;�:p�@q���#,]��\=���k"M�!���2܌Yյz����}ŀ=��C$�l�d25��t��?n��40�T.Xˠ�t�F�Ds7�}���i�Jx\1�z��']�����
�Î���&W�y�����c�Y�6tc6i5�j�[��'���Pg>P�#��i���,qp���X4�:�G8�+���OA'8�Z	"+��TW�KLj�>H/�u��jS�;����@z�4�w0ӭ5�'��s��ƒ@�\A��i�R�XD4�!�������!�y.�:�~O�����qPq��7�Y�L�t�k�Cv�?}����p�OQ�b�CkM��pO�J�+F��
�������ftw���T@3���u"u#�$&�mu�vD�I�� B"�>3~X4��4��$p���#"����c ��Z�lt�
�g-���������Ϻ����4��c���[$Y���(hr��;h��	�:Y��c���}�.��.se��{�?3�#�EV#�{�_�sPeM�B�i���v��4Ox��:X��p� �DWpY������
�BmW��ӄ�&�{��P��C"�S+���J/���ᜧ�Ԟ����'��dR�f
ӹU�wu���ff9Y�[��(=�;�3�4e�8GD:�Y��b�U�Y�i�$��4b��G�왈�,�NV���}�[�v��z�OI�Rc�3d巟`�i!�A��f�fd��p�N�)�y{^�wa�A~���G�w���|.��3@!�5Ft�U^�݈��GP@�l�鬾����3�pj�A6h3C���{�g�rT��i������wV^�v9�g��X<�+�z�L���<s�^Ms��?|�q�<�	��-���5���i����hKHȾ-���*��~#MF~��~8>�ڥ*��W�p��txP�����M����_�J�ޱ�� a�|��f�>��e ����,��NЅ�!���Z�"5)���@��.S�K��������R�G��f�ެ�htg_H8��@�l�������;|d�t��L�d�42��l��C^*� ��X}ֺ������X�����!Ф�![�4�|��:t�k�,�������H��I��4$AyW��5�g%,��_s_��o_GH*�3���{��Y�¸X�>~!R,4;�|v>#��z-VmPdp塾��.�)�q8"N�Ӥ|�ĵB�7�_�T��D,���z2���AE3mH�h3_/��ސ4���
*��r���-��AbG	5�o�����_KΌ	��T&c�d|j>=�$��I��")���i�$3�^(����*'�o�vX�ZBj��� ���#_!���=���������[�B��"��I�g�s���9��T J�y��M����S�N����ϯ��>W!j��]~�t�*�9f�'0��_L��w:�ҡ@n�C[ޘy.�1 3N���1��s]b
��ؔ++5�)�3pd9󳵲ˌ�7N�v+\���[�k���%ՀŶƙwZ���K�ȃ�#�p�\Z��N�c��l������ m�h�m�VRѻ5�v6��5�L�Ze-V䙕(���#V;c6�O[b_a);0h`�J����u��	)Jm�����V��g�����j��<����e��ݪ0�4'Yy����pp��o>�N�ɜ��n+rv�Y�h笹���.Ձ�F�6��I'[������Ҝ"�Wb<��a`��JI'��Gƃ!��ZЄYϕ��U���@�����,�9j��Z5��zl3Pf�Dn�,�؈�#����a���Gn{;�s���:X^p�b���!����F���:�@3dY�P�A��E!8�A�㱦�:QE� Y����L���@��۹�-�'������z�5V+H �5����C���Y��ȀFf�5o�+Fut�!Z�26ra������Ui$p���E����1e�=����drPj8[r-��|y��I���mύ�u���A4,��fF����o�Gȟ��Ԗ$ ��0g���xK5LC}@nI�ba��8A<���sa�I43�ߍ�#N��`�3�U���L5e��S��ȏ�D&� �����F�_w���Yc�g����*�v�;�cƸh3L��㡄f*���;��B�<E���0����`^-< VY��G4������#D��ǜу�p���Jĉ?v�0���֒d�2
���q�t8p��9��@dzqϷ��!���VkH���G���qv}�3�⟯x2�*�֞4!kX�L��OMi�!�0��}�k�|��t�)�f�F����f��|+bP�!���;�i����1������G��y����!��dX���V\ݲm�����<""�Iq�­a�}�t4�t�h{��CeQ��o�2���A�VD42*������}�z�����Pt_���Tb�&��"^g����Hߓ�5;&KHL���Ǳ�j��K6&��sß�pu4!��A��@q}{�,@h��_a*j�ă�Nn��Su�C��hŸ5f��TЛzT��b��-�T�ƴ4�=�x�]He(,�y b����:�����2uڻ���ݼߨ�l�6[#��h{�����՛ţ�?��	6�j��$�.�wSǆ���@���4�fW鮖��½�b����)����:���*�����er�ƚ�����I�X,��Ȁ��vG��B i�^g�(i֞ 3Ϗ�Xxy�\����"Ǽ�a���sz�e�����3CN�js�b�V�>6}�a��d#�$�^�.�h]�%4��|����HC��ht�q~0ղ�
�n��_���~KƬ[\��(ЫU9<�)������K�#����1SH���C��@�)d�gǘxow����]��t4й�?;9��Y�ɻ?����}��(�\9CO�_�
��^�ߝ��A������Ux`�o|,:F]�*��l�{l|k�a��d.[�=�f������A=4���}~�݋#�MX#������f�����?M�}��0�R�R$�i��R��M�ʸ��nO=���9�^���ن輭n
GMnMs��9�s������#��|͸p�:GMa� ņ��Y���郤iޡ��Q=��"��t��~vȄ���俴{��8t��S҅&~���5�����Xc����R�� �PϏA��� ����M�cH��k>���U������b�U�f��\+������Hχ������B4>4���yCMx�D��,��?}�AK�!���x�41���:htk=�}�<���)������-��Y]L��ɠi҈��aϒ%Rҽ���:A4���08l�6A����0����!�S��o+���
�r܀���!�Zl�vݜO��^<ߗ>�}�+���,f��v��"�JYr˷�sF����L�op���j�G�O��W���O>�3dbAZ�{��GH$���������iӴ�MY�|k_�H5!�Smz��!TS�{ߞgg4A6��v�u*�58�g�	%���E�V}7��6xhB�� |��8�f����]���ax�.|���_�'d�o�;�^4Mh��H��-�����f�\�;����k$D4�h�$��lk�,~���#�5e�F�so�nm�e{�ч�|�X�E�І���44�c�����x`��
c�֊�`��t`��߶�p���b�Y�D�hgO܇�؄�_KE&��e.ӇdPݨ�m3a�!���|��9G��uנ�:Z5�gh?��=�!��t�^^ϝ���H�Q���ސ0���ec���-L�Mt�GCB?}��Hngg��s9����0,���S���u:U�]�f��H~�}����&ޓ�����;�Rk��ۿD��$�."@��z~�ߝМCj���_��A��5��4]��8��]Ha����K�[��iB,ϵ�f��&D4���f�< #�٦���.P�0���GV��K�(j�z����&;9н^G�$�����ī��:�~o�u�j��Y7��9 �oǝ��I$jӮ>c��~�޵\*qႀ�"?-ㆂw����*�bn�iu5Bz��ɵjILI"������|+EhD%�+��0P��P����b��⮤���G1j��},,���Ciz�i{��v��i`���!T���Z��[��Cty�V
�ա��{��`Bc)���� -�t^'�kh�ź�-�`�vFs����ܱ{o�c��p�?�'���F�p���v��t0���&�����6�6�.��4�y�Xi'q��	�s��4x��"�Y`١k��&���?!�N��^C�P���e������p��:�v�2�~ZD�Qo4X����	��A���ɇ��wlw��+�+��Wl�5�ȱJqě���n�J[��Q�t�a��uv��tF�h�k
��G�:��C> ����P�	��Y��<0�Y����wן,z����VF��~�`�CO"�ԛ��>�=yB�^��j� h�"P���]�j����Y;:^Jp"L�^��O�V���H�l��[�li�
M"�Ç�����E`�kۗn�o�S TF�!s���C�F�P6X,�,���,�|����C��y�f�4����o-��^���t�
=�E����Ӎ!D}=g�_�"Љ�EyZGgcB5d�@?{�	�!�L��4V�5�Bb����c��q���}�B��Ͼ[�����ߝa�rn<�q#��m$��a�3�N�ZF�0��	�H�hn}�u��0�h�Ď�6�>B�dY!/�p:�=�s���U�����H�j��q|CY����g/�M]��h�ݰ���,�����i��6j�Vq�d��<��h��K+�f�}����p��T"�Y&��)}	fiv�k�)��������=?b�3�7����l��!ĉ5'�#�>GOi����V���`t���
#�B� Yd����>#He�!M B�C>ﾖ<k�����LT�%�/`/�B?eN���r`ٖ�iLc��0A�.�2)�$�)�gr�Yɡ�Ӵ�JpI��o�s����/7�N�]��Ɓm#Qط����������v�v�ܷ�PH����9[S�jDA�5.bJC����	��j�����zܛv����Z�S��2(/v;3�y������wI��S�����݉�W}O��w6��Z+K+k�5��[m�nUZ�SluK�-n���0L�N��"��wIH=���.Їk�h.wTa�3���m��8�1������Ŝ\b]��'nK��_Q��$񌬫�����ݹx�7:9��jr�˛���I�D�]��1ib��T���n��P���^�������<Yj��i5�N��3������>����VG��T��Bds��lH�A�"���І�u�M�!�28p�\#pip��~,�#�\�E�	F}�� ��Ͼ=�6kI����Z�s g�9޼�s��X���,�D*FM5���0֑�A�ֺ���{�E���oجsʽ�"?l��YX?}PA[���U�e�%y��h������,�]����=5����G�	�g{.��Vc�4;�~ Y��_s3��$p�N��5��}ϱX#GH����<W��+�	�t,�F��#H�-0�4X���e��K�_o8hO�bA0F�ьmI6�FY�@#��S����(P��T��j����F���j8I�C�� �B5�ϸ�2�T=�����uB�r���z@f��&i����?��@�'��j��i���<k��~%'�k?�l5Z#MA"�^4�4�kH6���D�{� ���:���j��˵��������l��CG��gx�b�3Z��X4P'Eh�_�`�F�wM�b�:����}�#Ǥy!���� �v��}���:��#��x�����]��!���k�Wc�X��=i�&^[\^N\�u������ϲ|xD����	3�ц�J�~:��`t����+�z@�� �dO��%��޺�\�{��j�=� T;ߍ�'�m��������^"F����h����!�������x�m�$%�Ӓ�o����qQh�4{�]�3>كi}����
�U�:R�9vbor��ݾzS��$�w`�i�
��imO��]Ak+b$O�0|-TV��ҥ��&b�f����}�������D]�D�K�_��a���n�(���T����������Y�w"����h�c��!���w��j�� p�Y�,������Wpfm̻mԝ��و�� RW{�[_���!B�����)/MX+��������>�ol��VޱŞ�����ǜ�|�	PF�0���N�üm�@���<�����C�6E�گ����i��M�b���0�@�X��||�؏7�3�7߶����FN:�s�O�h�D�ud���n�D_3�|�Y5�!x���%>_w뱽���xU?.�U�}4�x3�>�R���-WH�6�^���2ҊC�t|�k�_ �Cj���>�|i��Mgq�M���+��~���e�������B���^�����C6}�a7�M��6/W�*���Z���hZ6�4��0��(�N5J9���q�vJ˗q��k�NYtX�8�f%�f�K�X4aeS1�Ӄ��8Q �3�g>Ǡ�	��!�������|�#<�Bf���5.}�daSBȳLl��{��`)xXװ�7t����4A73Ä2,����
4�/��A�_�ä#E>xo���)��n.|GH�� �"�:G����>7C�8��O����A�y>u�dk�+>�4�B�v*�i��I{�>7L�xhC~�'�i �!{�r] O�>���=?�$�'_�_�\�ZVV�q����M��4�h{׿+#��2^0͐�{F�!s�+ﳝ7C�΂5�y�ײ��W�.	{�i���P,5`���Z����;݈)��>wG|��p�S��h���N ���r^Vb�L\�Z9�u���3���J�ɠ+G$~�L����P�ʬ�o�C7~��Zk��K}�cH�_B7�x�,7�GMWiԝ�)*�~?��=���9�оD|��Yfm��N<aF�G��F���	:��VC�PXe�{�L���v4��Mf�"�{����/dF����Ta���<���dK���m��d.��pi���p�|@�sw�ϦV�"}Ն����B0{ܾ_,-���U�"g�jȆA�١=��:F�|���'"f��HF�����<q���< YG
&9/�{Ǯ�����-�(450��e�Z�'��g�7s��.uЕ��q�u�	��9n��OI���I
�\{��%��xF��D}d�a�B���w��:��H<�\���A���8�߆1~���W������Ɠ�+_D3]B�{�f���c�����O%8Vl�?Ou�9!ۇ Ӧ����44���}Μ�#�N|���<wGJ ��"����d	��-rд���~eT*�ϝ���:Q�D��,�e8Iܿ�.������>�Z��I� �5��3L}M���N��S-�K��?rzs�}���u!Ȁz��_>9CH�`\"��F��,i���n�;/����;��
�͉f�Gư��z{��ᠢG����O�^����5W0G� K�#��2'�����K�4�s�<"<)�1ads�Ea{^&�Up'�u^7�H�(� �N�t,�����.����j��Yj���� Ϟ�1�X{߃��4�A\��uv��V�n�#�ύ��+{2� ,"���e_�{��n�~�7��N��C��1%�nH[cTglA��{�g�S�߂����!�bQV�<�n��$8�����ئH����ONzJH�㖳	b����m�;eU� {u�V��9�����w�}���<i�P��6��, Y�z���<$�4N��5��3\��X4��>�Px�Փ#��m�k�o=�Ͽ5�'�m��_q�A�BS,�ח��ص�v��V-ڊ�`�i��P3�g40#f���XLAq���Y��C"�EYF����ZA��Z�qB4b��%���n��td�;<�4,�,��X�����!��I�x@���1,"O�>�c�[ZY �A�w�#t):�����8�����y����D8l՟,�9�ٟp]��q-'Gk�&m,T����a�D�}�������&G����C����T+M~ GH�֭|��60֚h�>���?|t��H�:�{�,T38Ѝ(C0ӑ��#uVl�]9�ȽA4\~����t�0�0�� �]�|�r�#�f��K����j����;��6~�d����H{#�-0��y�67�i�M�8b5�Ȇ�v� ��!�l*ObD Q)����1� r��g�������p��~~�֖t�p�"�Y�衜�W�e��8��1>�1���Օ�����"Ѝ�#t�XB��(/�~������|��Nv�E�P{u�t�4��l�����`���B��;�#L,���8@'�S;���9�GK:8D�Ua�|�ǳ��9]��=Ø@��&H�-3�޶�5������.��δh]#- �B0��_�\4X�(Y����6��f_�Vp;��?�e�D.�q��;{1��-���
c=�����ͪn�d[l}:����Rf���wL�9n'ȬT�LRQ��&���.� �s��Od��5��>畛�w�7���K�+i�ثeE�8N[��ٹ�gRK��u����F{3;^5Z�`���']����;X�#�1�	�I��`yt��OW��W��h ��5/j�ϊ�I[� |��v���}�Ev��-	�`.�����l� {AJ[w~�AxS�G؊��C8(mۘ,?z=W��F����Xz���ej�x=t��´�a�Z]\�@��eu���z2T�?��a�=Q+��eЎ���i�JX*�lM%̢�+j�{��}����1t�+B����)��;w�V������h")A���W���1nhk�іf+=Ƃ�mJ�Op1w���%���[ُ*����G���5{�v�)V:Ӧ��n|��ĥ�o)&(�6S%-���v���8�G݉Fl7
����;��^��
ۤ6�\��M���ά�-�j,�ާ{֦��t���[�^����.u�3{�5���F���78Wx�s�kBu������vA۲dB����th�f�®fҽ��f>�{b�%�u�νLh�q��Kpe+ �MX2Sl9�wސ�Dۂ���Dh֎e�����t}��G_mc�g��-�u��R�A}'5Q�9w���'d^�H+S}�����y;��Ҁ�r�h��]L���;�ӫ����m,�������Um�mj�:7f&֯*�N��������m���m�j��%����e��uR�	r;L��Ѭ��ԅ�9^&9��1�nq�m�oqk��5uЭ���h2�lʖ@����c2\���^*,zJm��L��ĥ��!�^m5��-f��R=���q���0Ù��+61R+Ku�<���]�cV7���{̼N���9h����i �p�o�*�$�0�r�-����h��s�S�oI��9�a�gn�h.��[j�� ٷO�	��[���E���:�^\^M���m�v s�{r=��t�S���l+3�n���^e̴��S����+�r�[��<d.k�����H��q�rݸ�`a�Gm�8�t-��X�5��vNN�`68�נ懳��{��O�;lVI�4燍�Z'&��ÈUI)��76��}�Ie�
tV��V��;f`�[F�7Z����E�gaY�\)Us�7;\ġ�$e�L��f#ݫuΑX3�,��i��9�.zg �u�H��rU���&�g�Dg���m��rh���T�c��� %���m�l�t�a鵖��HT�v�N��\l\�prf��q�+�"��.�V�.)�N%��z�ٸ���&r���lRi�m�.5"V�$�ji�`�ͼ+,e֥:k��NQ݊�,�ۛkک�yb�15v��D�U8��goe���d`̦�d8�ܸ����m>�7d.b۹��k�3�r��Vz�nh˷,�ք�D��0��6�U��,�5�Ϸ6�x���ż"�`�cur��	�8Z�=�$"�c�E�= M�"��ٹg��m5�^�6��嵗Tk��*w�����!T�ʊ��5�������q�-ʶvls[���K�W]iE�gvr�N2�6.��Y7qŬ�F��Sa ���Q(�<:��1�y�W^EzŹ�2��V�wAv�<Xt�����ܡcvwa;;n��j��2�[�#��Ҵ�[���,2�eV�#��6�}��NuA��!�r���Y���5��Sm����W<{F�my�/�]:�	7k����h��i�lT��Q����7��6ݭ]�xٞ[�)��/Q�ڵÖ��hu��*]�.���F��虭�,�s�:A
#�A�ެ����f�V�1���i>cl"n6L��v�R������OlF�Q��ݪ��N�N:벊��F1���
n�(�mƇS�n��n��y��F�v��F-U�� X�|A��N���p�|Z̿�����k� x�U;B��������oH�1Y���,�M�����>��}������ή�0��Y��w�~=m�$WS4�,�D!t��_����|1��i�L�E=�=�R�F�4 �j����FZ��� ���"'�wkkƄQ�FZ�c�ov݀��:Fb�;9pY���X�;� �$}HD"�!�dp��� ��X)sՃ�]��P�'�YhEg>:9�`�MF��H��	$�^���1P�(�����;�|T!�a��!��߾ྐ=9�,���/�n]�w�G�R"ψ�s���M"	��Z{�Ϧ��f���8Y�,�tk�&���"�=�
&5�P��S�&�ʫ>�p�¦�n�P��?�W����[ٽW�\<,�PПz]Ր�:�?���kK4A��A��ζ��|��q/�!���A��n듳��0����g#H8a�I��	���e���HDD�H.�F�Y|!��,��C�^����G�=��D�G�3��J�{����7�s+������Y��R�Ap��7��xG��
 ��D�}�����W�w]5��S�o�%���}���4ʶ=��{N�;�[)dk��OYqۺ�!�A����C��V.i��-v%�܋���^5�,�"��4//>�4�t��dCA�2<�K��/��B/Um��1�[��O���^��=?o��ߍgc�d&�"���C9��8�J��E�0��a�G|W�0��0���ψ#���4�~�G�@���������/ ���6�G{������6�\W)뵝���n�QS-������7�H|��T����`9��ch�e󶮹<y�7��j�ƙ���jp�����\ 3�K���0q[?rC^����\]5��˻va��P��_������:�|/�{�/p����v H&��Xm"���D��#�����gׄ�|���Q�u��>��GL�#H�ڡ��e�3������hm{%�i^~��?�БU�����?[��'��D>�E�o�\�s����]���#uW�|�� ���Ph/��0Z& ۂ�:zxB5f�a-埗asO����0|C����J�����h"$T�����C��mt�6�f�3�+6Y�P�d�Lڌ2
��ڔ�Ͽ>2��W5��ϊ����O�P\T�H��+����)�(N*D�I�}�/P�8D<�>��$��C����܇W}��bh����]|a�{>��YgM/!��+P�>}�p߬?uY�@�f�hB�$�O�M��p��]�B�;Bd3�;��`�tϾ��L��-�Z�ii�7lz��sN<�n�d�x����7@q�˙�)��U��HcQI'�t�F���Y����'��5�LMq����>:��E�h��;�b���LR0�v�g���`K���j||�ad�qiR#���z����;d�G�ΊI�n����\�]0�z�'��	��.z4��ZW�]��\<<"k�}�����=�'~T4M"�Ԣ��$L
�&�=\6hY��}�;��H�y�;(� KXE�����i�o���}C�w1��ʐ!���v{k�BƩ�UV�_�p"�Hg�A�|��#g��uV�xWH�Vp�d�"�^�����ӽA���)���4
��e������Ǐv�ivX��-u����O��J��YI����FӮ�:�Ww���ؘ�I�A�>64���ΕW�{44��"��C��I8a�u�<�}�|0�����0�D��䱭C��aB@�[��⣪�,�,ϵi�W��x�#���;��ß!ӆ��_rS"��y%7x�]i�t �"����9��!�����H)..f�������#���]#�'���t�y�p�"H��~���G�HU�U�u'g��X��$P�C^���w�Ð��A��/�l�Ԋ|�=�hg�d�At>�W���hdX9�'ܳcMq*�%B4�,�w�}٘xi$\����_!���M<���h���$4��ےc��W(�]��:�|4q�b��� Ӂ��k�yph�m�K\M������Y�Oݩ���ӎ�!f�9�t]p��8l��T,�m����t'��;�v�;Yj%N������>߈���>y}���T���9'��ph��%jg�U߸�f�~�4�d�����_���ͪ�;�d8����⡇m#1P�}�E�5�+k������|�$	���	�Y�m�`ϕ�]@D�p�42/���䴁��wz Di ��L���҈�g����ߟӏ�l��2:m��w�#玡nK�����S��>��g�#��n��e��@�{DZD��f���	��.Y�q���jz_�z0�H1hj�+��ŀwMh">#qY�����,8�I j�G��%��\1/�_CrX�B���p��>��">��}b��!�y��ʳ�bdU|B�fe.1�/�}僤x������s��1 �T@q=�Hi���`h;Ť51T0&:x:~��2>���]zJ��ww����[�k^���s��kM)��i�>�-f���֊̻Iu��nN�{{�����:�{Up�H׎�s��Y���� �e��xtO
O�:;혇ih>��,�W�N��$��3�3��`�G��mi��������s�-�Vy��*�.�&����KD�?�Y|Y�Q�6h[��
H+]"�:E�y�����|a>� ��0�IKd��T���e:�r��9���ɍ�o�m�ϴ�D2���T � ���{bb������,�$��s�u1!��,��*�����_H�L�uV�bF�f�DB�`�O���`�K?_$�>ݹ��<�MQ��h	·qP�}�lt�G�q�f��CBrM��W*@�Q�qm"��!}@;SU��M^�c��+D��FZ^^�K�Ȇ�z�"4�;nc���R�-c�?e�1O��Cc�ǅa�\�`a����qX�@��3����v8�^�D�*�Fhp��:z�i\�G$�8^��O�Ӧ��}@Ya��{�`g˄+��D����!Gv_=�����T!>�+�y�O�#��à�8{��������YD2�CSˇ9��.�I�j,�ݰH�^v���V�y)\6Q��;:D�'�d� 뻉��}����h����N
��g�� p�{��!��}�u���H�\�hr�a�oe������q !��ܙ9�;��߇ʄ���􁦐$���Y�N������*?�J��:����F�qB	�da/���k�w����V��3�����q��j��}�s���)�@�Ơ�k��4�uOT�4�@e���/U[@�w��#� �wW�e��P���_b�y�������/[�RtK^J�t��pa���U�C{�F��PDZ��`��k�`b�v7�������Qfة-(�}�W�T�[��e�hkf�)�m���t�[<Wm����A[}/O�xL8�^N����b�V�Y�@�-B��ő�
zn�]��yL��9�yy��xCoDx��G�����=q��ps׳������T���rm�qNq�ܚ��(�\S�B�Mb⺧+[Q%M�V6�f湘rv��8u�p�����:�7X���m�yl�½�A��nz�9ر���&�MO�VTOm�l<�ۙ1 �9�v:��/;�.����������)��Ng�]�#�.�`�h/e����=g�w��f= Y��;D��B���9黳��G��#� ��t�l��妰�3�ҥ�pQ^�vA�}��V�٪m��{�dM�$,�$qI�8|h3A��гC�����5�x:G~�~;:��f�jy6s�t�y�co_e",�(�L�i�k�h�ˆ�2 !:���}�X��PpwM��>�� �ܡ}U�=j��6� ERJ#PH���G_����9�|4u ����FP�<=6C7���G��0]B'�4���]�}z>�Z�����a� 3\8j4;y�����w1T�#���^��e2y\(�Ց��"�{������gW��5�MT_{�Ɇ�P��<#52G�5�1\>��T�}uV�C1�v�O�������B���|>M���Ji�Z`��� 7�8}���3]���}�ōX���H,a�5�!���D!"cy��ˡ�0� |yj��v}~W�ư�r��.;鯋��f����o��_}'����������Cd�у�iᡶ�3^�Ś_���ķ��Yio��l)4�����-�۵]pk��%��nYR{\�����\�-QΏ��VE�,�ϐ�0��׿j��8I.�M��Ͼ��Yf��sEÆ���Vk�CBD��ق�R|�ϳ��f�A��`�,���;A9{���\4;%9��+'I��-m�����6תi����t�C�aGǫ��c��+w����g���ڻd�sq�{����ZF����O淅�f��r��F�(�,�	X[�'�*e>�Lڛ܁�a�Y�-��3��Y>O��4���X�!�@qW|��x�8�q�|�ٲ�$�$h}o��J���.�t{��G}�T(h3�����@��,F����s��(��Ejr��Gx��ӂ���b8q�&���ί2{�9�ZY��2�'��p��h"y���׈��$T����ن�ꯒd	�W���`�83� ���18ۃ�e\AfDw靿������Yu�_>YC� ~�:������1п�8���qP�U�"�����<4��؅���`o�B��5�.��*Ӥ7M� a�����J}k̹P�!I#qe|I��-�W����Di3ٟ+��4�[�	���Wr����N����Upf?�uE� �@�B�p��h����ӧf�kk��"����R8p�ל�ü3�j4� ���L��n��<�����hrPF�eMՍ�w:��O-��8.�<^�v�O�<��/#w�<zl�~����S��C��3Q6B#�V�s�-����֙�9lBH�e��ߺ.��!�46Ր!���`w>�|���|GƸg}�j��\,�k����5��Ihr*�!��o���tpI0@�pB�9CM}��#�L���MMA:y7����2�~����Ϯ���no�5w�8�� CP�U��%\Ϟ�xh3�G��1Q6p�_n`��<t��7������oՇ�ƴD%��~�3`m��a2@v���;?	:;'``:9�uY�W~���3�x������B��:�⾦ ����7���2r����.\ǻ��۵���`�e�J���!{[d!ݫ�����L���.�7�pR
����wn9����Z�O���_�g"��&r4G�X0�5qQ��,c�֑"}����V:�������M��"l9#��< ��"�Y��g��/����C57����׈��Y�����"�^|l4���6h{}X����,J�,Ղ�g����|ou����dE��u�H�*}͕�n�~����û�i$��̢Ӑ_HkH�U�,�E�mK��~64@(7C��C�H�V+���'�$��~ Og���!�(*�ƈ�R�Ӈ� Rk�>Z�{=}44�<`"'Nb@�'�t^�/��5��A�����[�3>�˜��e��E�$a�i8q����J�0�N�^��Ξ��*�J�KG*��K�R���v=�ߪ'�<%��s��	�HV���FYJ;�����Z�%��s����k��!Z�6'�o�����s���VG����0�Oɑx�����}��l�
 }ϯ�຾mM���s��r{⓲c����d}k��WCH�3��x�;H�W�!�N��:�!�B� ��ߎ��hC.1��4/��X�U���G��r"�nz7��w��8�ƾx9�di� ���;�䫆��Si��#P���)���0�ت����#R�����(sx��f��m^�t44�����{:09ԏY�D 2M	���YH{����T�,�ߚ��H���07qXZ� ���@)f�R��qhժ/G��'�J���I�u:��{1\��|1�h��1f������ ?yw�|$�w�����u��|�4r�s�M���*<����u��N�h��8�0'�jS!��7<Q(5�)^!��P���¦���8:�]OT��g��AVD>� �5���:ij�w���qBⅨTe�!��_D	5!��hj��CH�͎�j�G�P�����?k��Ư����.��Z>CEc4G�
`����dѰ�!E�$���k}��^�H��i��!w��x��S�}���������h��AD$j	%��\n:LS<�[nn�u��۱c�=f��ɳ�V䉱	w+������=�b@����I�d���x=#��6���'��}�4�M�	=4�6k�0���9O�?�{v��9��G«��9�E}�G�}�c����ۯ���!3��49`��_Ba8��H���_$,�i��f�}��~���z|x>>~ɜ��A� �CP�~��e| �՚>]�X@%w��� ���;�/��\���.�]��1�� -��$���}��rXMb�9����Zo o���dA�<�p�Y�)�����f���E��x�ݓ�,T>�Vl� ˿/�[4J��k~~Ջ��=4GĞ���X� <4!da�K1P�}��uWz�ł/�Q�4Lՙ{���1l��q���/ǛK�� �j�x>ڂ}�o7O@�U��f󣕤�u&D!�d|j�k������G�x�C���ƀ�=�� xhC݂X��3;:{)C��Ӕc�w�}L|>j�!���f*t}Y�8�ƄN��H�,��g'W&�g������zi�z���<����s6��6Uڼ7L�z�CS��4;���F���|�p� �0�>�Y���$H�wP�}����z��D$������ۿ|���./����V�{�R�3c8U�j5������o{n�-so�dY�Н�������-��k�V,��M��է�ڏ���2ix�V7$\�m��9���܆��M�n0��c������n�nI7r�n�[�
�Օ�WݏF���=�/rl=s�6X3�X������Pu����qq�Y�ծ�@М8��.�����f��9P�h�Pe�785;a���9䧘zm�gf�u�#����t�4&s1!ǅ�	�\U깵��z����Wguq��v=s��a-��Ӆ�VX�ɸ묙}h��2�<=�n�37Bv39�m�]�ٙ�X:뛟�d�=���thIH~����"��}l����Pf�������#M�	��z�~��,��V��	'�{���� !�Ou�H�^��U������:e�]�T<��:S���k���\����L�½=�@Y�}���U��DϾY��9�� _��wSF/� ��� i��
��æ�F޶I�w�{� p��/D�� ��P����T?h�@P��O���՗9CH�q>5�/�hq�
@��iv�^�$􈑕������ts�B/�X�8t�����<�(i�u�t�;�W��t��y�G9����r�8h3A���`e�A�2!X�� <��5��;#Ǥ"�8���@��x�|҅�Kh� ��M���B���ze���3GA��f���s�(gUt�a�_<t,�j��|l?X|�ư�b��ˊ��~�߆��`�9���eQCL'Ǔު=��Vp顖��H��t�#%��C���{�U6Dv{�zOLExы��2�a�)+����A�k�2m�zo�7q{����� _�D)s�Y�f]�a���^COx�M af��j�>�X��I�Ǹ��� 8=�O1�r���L1�ؐ�H�g�n¼�d�[���]���s4�vMM�sWc�'<�a�H2�^��_vسD�7��p���tX�ZE��Nc�5�*�}�� #_�U1�<HU��}�O��U�ip��G�����՛#����!�������i�곘��pՐ�"��~��o�\m���Ͽ4��Y?+t��f�J=�E�gH���p߻7_[-~'����X�/Vꠃ�/Pp{}��nP��O���zt�9�ב��.|4t91�U���;MnS+)�������_7�8'\U��uX���yCJ%c+���1o�����`]���֐�EP�
%D�#���ZG"=�wW>��4z}�}��|P���KM��\��u�g%9-�V_��`}���!��FHa���v��V	^��C��<jjEeͤ>�@��w�<���!���i��F�0��3E���:hm��!5����������ڈ���i�� t�;��_Z�8F*�ދ����L�+4�0������z���<5/�cM-�/�]�Gx�@F͐8���i�v:{�᧟}��	��������6�����QW�n55�>I���	�H�ZD��~ f,?F�x�~�8{p�lT_��
B�$����%He����X��ZF��B�2�!������D�@IBְ!����`��s޺g�f�P�#���ް��[�3>�o8y�!��f�Sj�K���0%��Սs�r�Onv��m�ȷ�F� �퓕"�����p���iS�:-���=TmP�H��S�}���\$������~8ha��;�5X���o���x��>�� �CǏ�Y�>�������"c��?���S��w5t�p���41��0�5��9�J}r�	�>�s��������Cf��|��!_gn�ܜP�49p�Q$I����`o�ή6󒰲�o�h�����X�߈}��y��{�V�+`����6�\D�N9$���NU��#�g�}��W��Bd2���������p���k���ϗ��?{zѿmJvo\��\�CS��t(��7�҅{h��4��xa8dy��0ھ��4;����J(WS;d�s9b���Kxؾ���i�����d4[v�S�
��]����l���J-�o�ζ�e �[Xp��V��a|�6㶆�ն�����5�Dm��̒�,����Ć$���ہ�v���9;��KE�����kf��N����l�s疝�i�c]��1���DqXevv�;��69-�ٜ�h�����q��a��]v�	χf/�	���6�Lӧ��y�zR}^p����R��5p�3+V��w��C�l۷��s:���e��?_[�TV�L����6-��Wn�Mw�Rb�fX�~G�f���_&�����d��H�Zl�i����!�,t�Z��b����S>��Vu�[]:�ݢ��i�8fc�W<X�����w3I���}r���z��v��%���k/�oA�e��\�$����r��ɐ'M�VWj�Cz�5���#}�wʾV�[�2��ܮn��g�&��u�7ug�:1�ܠD��7ڂ�M�PKٸ���s��r�%���h@l%�L7K"��f���}aݻP^����s�6���+�����r�=�n��k»��)}FL�������9���9���u�`���:�U�-ݾ�x<;e�'v֪u:��:m'��z���"�r\y$��v���x�+Ec�m���=z�n�ܲ)��ݑ�������}n��+ߪ��{��_��g��k�ȡCd�E���b����1��Ѐ���$⩿o��&��
1D�X'gJ��8���=ό�`�!����&-?[u���j��?�WQ�^;H����^���s��k����b���SY-�ހ�s�-��tה	�F�䉴{���Z*���u���|}*t����<l���/o��㻎[��K/�d�{׏���y;�ߊ\�֭֌�d���ՎKţnθeW�v%������l
q��+<���!RS��
p-���{>�}=�����퇰�����^琊lK�L���C�O����½��**��6¦�K!�۽ ��j��
��W�8=^��'뜫/�x(���.��^�:�����<���`��^�3�{Gm/h�=G;�v
(.@"�N�m&k���N��7n�j�RCP��]~��N{F'�·�zfG6;˱���ްV=��i�J�՛!U
M��W�5v�2�f͝�V׆2�I��G1�f����M���Da��y���V�V��}�f���5��_fZk�JN���p��b��K�>��f��m�J�����Cta�6�H��4�{��㝫U�i�Dk����)6�e�)��7h�<�귋u��{B�Ǣná�$�7k=������z�L%��E��^�mE<��L�>d�R�ӜT���2���q���di�E�"+����J�+����v���=b5ds�Ŏ�^���BA����Jq�	|s/�r�y~������׃|c�2ȩ��yp���Cp�̤�4��y<AZ<�����ɡ��
2~�K6_�$}�_-l��A��|E��V���&k��l�;<n
�oE`A�y�ȵ�
������+��V-���G�U��ҽMW�W�$�H4�b�����]�/���_Cռ�cōz��w/�*�z��[:O]v	�f�yX)��_�̰�t �-��W�><#��ߤ�xy�ő��f��;����
��D2eOb���2�2��5غP��.���Z\�rk�L�\�V�GQ6TNI��$�j�Q�_��1A1�W
l�Ҽ��W^�m�t�������pW�<���뎗bGD�w)c���k��(c��t�wա�4��uͨ�_S9���M���R�*O]*��0�'j,��;�p�k`�K���{�X��B�B���7���g���z��ng<��U�H������۫�8�)��;�Ι�m\=�;-Z�e�q�r�ۚ�V��T8̝n��w\���{�i��n�s��H�M�H3D+-�&ME3��يE�� �P�J��V��g�[�n٫m��Csv��c>\6v|r���S��T㝌�we�'O ���nX�������qnʐ�CX̻KI��ٖ2�e�q�Q��0�i�E�y�����&qd+�"����ѹ4(���F��t�Ѓ,Ż��m&�x
9����x��C��~j�B^u���x�]g��N>w��/lL��S;z�yfj�=g��5���&i
)4 I��}�����٨���;��c`/t���k�vm	E�'v��m�hb�&��+`���.U�mʕ�7�n�)֬;L�gh�~<ôm�o��<�U�OS��vi��\*�g�q��˳���|K�?S��I�1b��kMX�J	
:]4GƑi773U�#y��k�Gy-��4�F���W��~��m4�}bH��i�;���<�|t���S���?��$�H�-��	:�.��ld�T��h�F�o��=���%��n&gG�z��u֢D����f5IO%)Q��󁡵������MiXlA3j�,ͺ[n�U!�i�����gR(�h��ru�ͧ�u�u�0�BlOrH�KR��w��o�㢘�܅wy�<�yQ̞^�[��@1j���պtiցjԆ�����bl�aM��m���3N��7�v7beYy}(��]ڔp�R+�8���A^�)���\�u�&eك�A��)�:�ĜE��w
�\Ν���Nr%�(s��9�@�!xՖ�_����s�]�ROϽ����f[�=^�8��P�qo�n�؈e�)ā2Ec��N�^��P���Ifc�4��Q���Z8/�Qz�j���k��ƨc��=�4�|�ب���U	�M��l���d���L��ޞ�x8S$��L��c!�>tn���+�R�Dn2��~����[�
���Y�PA!> �IQn�J -/˺ĺά��m���Cb*��JW��u;YI�W��i�X���CM=-������5P�a��ͫEq6	,�cZ:Ym�۩2Tva�1����r���#�-�N+��N���=�����&��Pm��w�+Q���p�U}B�

�	��=�X̝y��spx�Н��'�0Y.��i�8S!}rn�Su��{�q�ˮ>�R����\�Ea>�)�v���-��Yf���fx��M��M�I�xM��4���2=�{��;�V���;����j^�ӳ!X<k�xWP[��X$�[���lZwk�ξ@>������>ia�GCEϸe��4ڹ#-���A��Z|5��f"U뮛8�_?zG*)�q��aF[CgtSt�)��bC�A��ꮛ@����F�`��a~�(�(>�Y�����'�^3��}�/@��Cs$��Q�8z�>t�i0��l!=��H��!t��ُn�;��%7�i��b��=)q��jK�I�9�Y�,ԫ���ۻb�dz�I�����*��D��u���#�'����u$�*�1�1�x��q�N�u��h�z��^"��Ooo�����}�J6������H�0o�{]2e�A�X�jR������DȬُa��%?X�Lb��h"� �m�����^K�mz���H�E�Zt�w����}�Y�[Z�΋�4w��=�D�-1 s��f�M�,��2���)Q����N�2�Mf�������e�B��r�f��	��dT=�o��[�)�_:ݻ���|`>ɳB�-"ئ�n��椼��fEՕ����u�m>�.���9�[��`�B�۝�x��}_S�]\J��)��<}���.�n$��99ՓOk��]��.��<��u��3V��Ϋ�rcd�W$#������q��ݺB�X�	M�t�g10�����<n�1c=�]��>w��Q�כ�f�Z!�G{m��C�ܮ��B�aSq�_�]����tNj?2�anK�e[��Y7���k��h�푯�<b2�h�z,�	M��E�s�<sN���Wo���Z�7��:X[4�6�q�~^��<��Oj�
�_C�WyI_������M�-��[�:�/�'h2m^ݘ:!t[v}�8X��r��s��Z1��Ž�{Qj8����[:��A���6�d��4�I2�d��Y�ՙ�=�����L�OO�UE���	�Cln^vM~=عe��c�+S-�pB|[$�A�E:�s���]5���(g�%5�����k�5����R+Ӧ�xn���V�7�װΞ�ܬ��7��D&���L��*]U��y����T�5.�E۵�`�^ ����K�P�#��ַ��N��^��,����ucг�	���ǜSC�J���Lu����Dx�W`x�a��;^���(���Y̹NR�y��Hj>9��v�)ߴ��?��55���k�ܛ'�]�Ϟ�`�K��[��M�6b�#
J�jP�<q���8ֹ���\��av�8����#��;j��������ra��ݥ�5�Ks&{kdK�{8��4���v�C��;+��K�#����u�ˣ9��j��U����z�&�ƥ�9é���U���j��ˊj�[����i�ח�(�X2죰=t�*��tiq�v��bⴠrv���%�+��^:��T���2n+*�c��$�i7p�uM{/��3W�d[:�坄)�%g��lҿXְɃ���)F�vw_���fWH�$��t�I��r&�tO2֖WJ�O�xC��8͵��_S*y��8��}Y�%ʋz�p�b�f>9{�G&X{}J̉�Tm�N-���	�w�2��]ز���&���/C��`<��_���R�G�{���ظ-��xj
#M��@0�[�#���5��6#nw�]��p�{�uX@��IR�3� ��]� �������������Ey��A�k����pl*�2��Qt�M����רgMyf��̈׃֥����=�,�*�nv{�c
�X�qȐ0��$S��BtU�:�)iq>��t��{h�I��ö�:D���apU�J�j>�^qv��84��t�K��䂵ܦ����ҵ~9�m�F��v���W�0�H�t4	e��<�GArv�L>"�\<�	�y�];@�nĥ��Ờռٲ��%]^ЏK�m) �ޥx�=*S�w�<�y��w�m>1:wF�Uq��1{�b��띴e�z�襜\�YZ�kzN?z��t���ʹZ������a"c���y9Y�1�O7x-_u�!�Z��w[�k*���V�%P1�/����({�P��qR���aJ���2 �[b�-7��Gl�[/���"Ѽ�ؽ�>�8���svܕfs����6�&�o�-�@���k��r��Pۦ����&��]z�o��o���4��ղkF���]ǥ߫U�R]���1���P��W�����齃&4r���T�N��M��=�S��3i�ѯ2\E0��uѢm5����-م���>w�|�p9^�3Ӗ
o*�8m����1�]�.�?$��dv��i%�stގ>�;%�i�&�aX�"���ƪOc�j�z�(x,f�ӯrNc��C'e=� �jo�rZ�g����V�
C�4@��#�;�C�Yxm����E�.I�̚!VVu���{�x�<�C��BC�n�b�K��/�a6���ƭ��v��;X�I[��i�5a�����)<wXRvĨ������,nM�U��o]��3��n�V;Z��H-Z���"OR�vsr}Z(��$�S,�u<f
Cӭ/s:��}gy�Y�����T���n╾��59�G����z*S���@}+.�y�a�XS#B�-3�7ʊ��yh�Ax�]e��x���^c�M8߬��5��Z�oB�[�X�{�]�oʦIEfY��ט�otZN�b)��P���wY0��(ѣ��َMf��	�3�4��hƳ��_26�u����t�,����О2����%t�@��,�{���1s�V=۽���+���;��E�he���+��p�t�MXtP$�c_Zb��o�Y�^�ݽo'Z��ܛ�g�ٝܭ��K�Vx�Uj_M}�(�zs�+r�!��N�xދ���K�.��%0�F*t�m�#!�~�\y5ו^7C�^amI���up�g[���gL��:�Y��rzf�V�M�%"�eͶ��d}�ֱ#I���+#t ��s��/f�^�) �*���U�����vȁ��Vlo�'�k�h�lƉwO���n�}�3*���!lN���d<�WNRܷ�V�[�C�lߙy]���<����^�j��	��D欬�F!�* !��m��6]�x�>O�jk�ܤ�g~|�u�z���.�����RGE�����`�^�[��v]g�V���lKr5cݱ��2�_.`9g�ur��q�5�ۂ�u�l���A���83j�[��ۍ�:?�C�s����Q�9�x��S(x{�� ��trۖ����͂��6�t�F�Q!�M$؂�EZ!�A{'�*.wa�V�/���K�m�(��}�n�]�	�]3����J�����z1m���+��^��-��M����Ʃٻy��k�JsA���싻kg{����'�tۤ����?Q|o�`�<��wi0���1��m�񸤝`�~�:�:����^�{j<���G�����ߩd��w�fP��𱔃�);�Gp��a��M3L��-�,í��4����4������~r�	K;��Ǡ���7�O\���J<��{���>���]s��%iSh�^~�^�
[��%�����_G����V��rcK`3�������y6@9�c��V���.���ɦ��ﻐ9�Z�c�7R��4�a���Տ�	F٫|��eWc�,�+TY���az DZ�6�6U�t��S�*L˭}�x3G��l��S/Z��v�����f�CQܳw�c�*�
��_*�m��:��[�pcs�mib+)đ�2��h�<!��*�@y�k��ϳ7Y���qI��mtr���jEb��ud�Cyp�m�{��Q9��ph�I��YW�;kUC���]wg^i{x��Ǚ�=Lq�.fNaR���I��Զ_n��6�D4Ʀ�M�̵��܋����Xfn�ǡ>��O�[$wx5�8�s��;";N��������+�*���6M�BV�vyY�vwy+���.���ì� 1�*:�¥d�^Wu�F�F4���O����R�1A*�z;\����d�c�����ʗVl��ԯBs��V�q���p���A��;T@�(�X�[}M�=8ʎ��st��g*�>�������O4�Oq۲�
�F]���j�_����`�Cpi��N��tA[:��� �.�a6=���Y�)�#K��*�y5�}���`��am`�l�Q���]��*�����E$q�����ah��ñ�|���4Z�u�Z×/�U�nn������|����^l/v8=�o�bθ6�ڽz,BO�E��H�M#E5I���&�E�`�m���*2�WB#Jղ�[�&�˶�p���4����٠�U/2�p�����e�#�ؚx���^�u��,��q��5���,��兔�؈x��]c���9�W�Fs=�j�:X����-�6���=#��Fy�l<����剣n5�p�;v����|C`.xO�����Bd��V�� ���n�����6�{��v���P��eu����B�u/Bj�S����چ��\���Om��]ډ�5�qع����h�=�}T�M�f��֋{ ����cz�>��n���=�hN��*�kW9=��V��<;f�M�w=r�C0�^�]%V��=�lm7h�8x�mT��t��3�f���.7*DPh�&f�m3*��e!��6��1.�jU��)�#6�&2�ģ��5�Q��4�L�Sj�`�)�+\�&��"2�X��	B4m���oZ:�a�s�.�'�{�΃[��uJ�M�U�U��Z���
�y���i�A\�0��xs&���u:k\P|["��u��^�g����*�ݱ��8Xy�'Up�'W-�;[XG�
�;�mMX�5��[�bH���F����-���Y+�g�8�T����oN��;0k��&�,lj�e�Ѧk U�&�\�Q�˨�&����`���C
ɭkv�h1fe&]�c�ݍg	!��χ*�6T�"���lOQ�Up���7�qJNǨ܂۞��ɸF�,�r]�4�Ob����<Jlㄭ�W4�ĵ[U&�b�t&��=<�]{<:�v91³��n��\�lۯm�<�N���vѮ,���k���\6�ו��]\v��O\N�&B�3N;��X1�q睱jK��\�ۮÍa���>�/n{&��n�\N���;�ї��ȘzvB�O�4]��-וg]XV��iq�N�����^]N�׹���3p�5�ؤ�G��1�[��Һ2`�ID� s1Ֆީ1]���稚Wl�+vr��q <�y)ea�e㶓���]��5�Ǻ��ǷьU9����������<���K������l��p����t�!���L���)����e�!��`�ϓh燼;�<]��c��i���u�@�v�یY�lIn�E���1ȔDg�Ol��b͎�.}I�D�%��4��1��%�tHb��<u�ŋ����;J9�z��]���Z@h������wU��������8�H��Q�n.M�n�w*E��e���JJ����9�}���/9b3k�Q>|9=~	�nu��ť������e�b�n�����usU�9^u�n��yB�f����m�ǹfܵ:���,&a�UǪ�Z.�����Vm��{��aF�ʃl���� 	���%Sf�Le�g��^S�w.�����(�^���(9ssL_�u�dtC뛦��x�7��;u�Z9յ�BK�i$�E���y�</r��w'Vo^f�g�Ksǣ]��v��*��z���F3�m�8ٲ7i���4!mtE�g�,��੶(�ހּ��W�r+������mR���[37Y��5f�S��0��3Pˆ{,ӌa��ܡ+4K�VU��2�����sY�L:���M/`eF������.��������vP�&�ְ��b��������R�尭�)s
G����Q5ϫ$�B��;h1�������µ�|������s���@pTM2���2 �iݘ3�U�㵚ܡ]W��.t�1mb6-h��0�l���K̸�w˺7Vp�A@�}���Ǻ�ٳ������w3y�YvFn*S���F������lڗ:��v��~)���7K���A6�4�6�)��/���ր���Y�s3ͥ1����яY����<�Z�rinJ�ݫ�)�B61W�^��m�t���n�&S�|R6�LP ��^)eݢ6�F��S0�����懼����U���6%vxJwIy����	,&� ��m^6�ݜ5Ay^V�<�e���| Лp��9��H5��	�^U`�9���V��tmg�:fa*Ql�D\��tl�l�(�*�cn�f=�%��qO��0T�!��]ƒ�����m����剉.��b
tv��N�E'[�V��G)>�"N��rAҭ�֡��Am0Q�F�&�[�{�� �:�õ�Q���jF^��4a�	zG��x�X���.dW��y��^�6��b{I�!BB�rI!Ѷ��5��/i�ʡ�"Y���*n��<P�݋g���YZז�ޱٜ����:��|���Z�q\EtWO4��P�7w��N�(I�f�r^�G=P�Ũ�"A���V6�k�z���1���]γb��@�1_�B�_�}M"��x#���$M�-��<qww��W4Zˤ����������Og��u7�e1{ؙ��}��ؗ����(@���6�L�w����+�e]eǳ/9`�"N�٦��쎷��,Vu9��nd>]=� n��Pլ��Rc�*�9ma��!\h՚ Ѵ�nj��i���p9����n�,�"P�-���d.�Y���{���۷�gU��М�m�WHSX���kR�)ﭜ�I�D/�-�9�ݗm=f��co�;��"��K���`�[�^zY��x�u/~>�-z�o����3��m2g���8�}g)�̥���J�z���e���٤	��f�Ӛ��{���|���"%���j^	��c�>w�E�ǳix�n�]3T��]]��)bʺ��C�Pa�%5_MƉYoU빵8���74�E �A��u�.О����z��^�}�~*p�E;����(!'lV�z�d[+w���J�uF�\����U�����^�e�����7������̂���t���ſN���4	�^�Z�z��ۼ����"x�f��v��2^��%���x�2*K�D�����G�j�k)��a]ƣ�5��2�Jnj��l��\�-lƍ�T,�oB�Ys�Qm�6����u��{�+ȷ�@7�K�U���4WR~[����Q�co��7�!Y����Ӷ�Ǳs��)����Rrpi�%3�5M��Ǆ^ʃ��s;�ޛ�|2�#)R���fR,M�$��&,�������-Z�3���#i�զ�����z=��:�:���Tf��l�~��`޴�yk��<�+�1�JnM8@�U̯[	T���.�4e�S7k�{@jq+BZ��"�X������D���s݀"��L����gW���c}�`q᥏0g��\]6<��d���E�Ku]��\��Vaܸ�{��6]���1%�آ����Gi��X�:[�3wݐ�š��a����@�וTZ�L:��Y�鰎�=��맥�ʊYaa��x̮�ϸԻۙuz-2q�8����Ok�P���7V
[�N[m�Z��8A:������d���#�b;g�9g69�u[�� ɐ,ҋ����h�4��˖!���\B�bEnfΖ���vd�܊�2�<�4L���3�����z��|��wc���n)�Tת]�ٺݶ�/;�0�SX��˲U���;<]i��.L��z{=�ph��g�؁���|<;fN�Fz��w+���a-wk�Ȃio]�sp��oT��cA�8;g�f����Y3�:��t1μ<Z�"N���M���W�2��g�m���i�ź�b�[��e*X�p�Jf��0���"7|��7˦����H�Mu ۠����ڵ|�\�Yɇ.�7��"�[���k�v�e�G��.�D�qk���G�\�����Y�Y�y~@�̶�H��E��^�_-��g���+:�o�T�j^��-u�Z��ݙ�o˔��e"��^VM�ǮТ�:�		B>M�E�9�RI��`2��b�Ø�����}�9O��ۙhݮ|���}���Mܘ���O��\�9t��-y'�gZ��*"��Jd�]2Kg�k~�e�#|��v���Kq�W�y�ɹ�ˤF�{�S�Hk��#���׳��ef��/��ךmׇ��y�p�0\L1 <%�U��[X�Bb�띶�W6�V��Fs�����é��X�u)�����Qwӯz���k�F��q��Gh��Ff��ߏ�+��	6� �b��ƯL���v�-dA��TSe'Z�kCכ�vm
��Ng����Χ�mwjW�֟�=\V�=/v�pf��h���+g&)"�W��\�M`$���n��YF���o��]�����X#��=2,��p�4)Z�Ä���]�zd���V����aG��0�'�X�,�P#a��SM��'`�m�/@����o���m4�$��2�����oP/%.�.��p��!~�� �k�Kh�AE���?X�γ��h�GL����N�yB������n���"��=R	�3�LW"�i[^�!Q�8+0uȝu���N�gfJ������{�]	�<��k�x�^6�%և�kzsP�Hc����=x��} �
܉=�Q����H[<����ggl�X9h��	����:u���ep�v���5vb������|��R���d��,���s�e�3�'�^g��h��<���5bYF)��/����'b�PIA%�	�a��UaТb���=W�ﴽ�Y3�(�i��y�WX���>w�0a]�b0�������0H��B�4I`�(��$�����g����VhǓ��k���G���>�O���v<au��YS��;w�U��4�[y���s
��+�}���^�얻s�hM�d�ֈ��s���e�أ�	�q�^\�w���ӳǼ��� /�i�����E��n��;��;î����fo{7Ng����s1q"꤯u�'�a���y(rڂ+�S���������|��"�D"�(2ػ��c����hzSH3�Ě"������V���Ϋ��ʠ�d��˕����B��|�����cn�\��M��x���pE9����ۚ�PI����k=�˴��c$�2�%��l<W19�
�]�9���Gц�vZXC$r�{�S�f�h�{d��a�d��ym26��Jj��
,"i��j	s�����:�*��lK�@��4[�y���8�J��*�-��߉�8�{�p1�m�L�p �cH/��)��e�>�d��4j$WN�4g?W��b����x�{���漏�l��Y@#�X)���t�!A0Cn��sl��å�-��'m��	c��c^������=aO`�8W�N�!v���`=x+ļ�qޥM��u�� u�7�Ǳv*�54�{�bg����e�ώ����S�zƉ&Q�@�ܙ|cÛ��L���T$�QV��h��L+$�*T�w7���M>|Vk���m��l$�QsGW�i��hV�i�N�p�AD9�۷�X���U�_�����9N��.���ŷ(x����2�;��*���ۛOh��.=U���:����q�X���G�6�'2���
Z � ��a��V��M�V:�{na~<V�a)Q�/W�$I.��e2�����g6:�y0k zIƌ}H�^�zU�6`"�{�C�:�	w�����W7m�xow I��)(Ȣ�k�Yj�Mfim�����ö���E$L�@�(j��;����X9��ضBXt2���9u�7���K+������Le���,���C�,Ư}����|b<����Բ�)��Ҝ>si���m^�يc�����3�;�5ʑ��m�i���� ���_y�ٗ���7]�Z���;���)
�*�t�1��VL[������Ppm�J\V=�h�Ͷ�{QV�U��|�Z�z��C��-�ЯF(�d�!��loo��\Aj�-厽?�.�Ǝ�Ky���GV�h��I�.�=F+nlm�Y�&�Ƨ���ݒoZ����>\:�U�2�%������-����6�&���&lC	4��n��L���ڽ���쫰��w����d3���ڭ��<):%�X�s��X�'/.ںg����v���t=�\��2gwg�Sԣ۬�W���s/=(잎D�q�_�p��� nRbCilŨYs� �k0��9�j*��c4+�&��7���ַ7�,�#������u۞̲tn��u8�e�-����`�y-�4���X̒0�^Y֡�q�wm`郘��G!��^�a��봘��=�3`4,a��l`�|��Z�
�(w���+� qL�G�/�z���F{VD;ШӇ�m4��A�#�˲0j(Zm�"6]c-�t'�a�{V��.o��`�'�P[��B��G�zn����՘[��6�$ʹ1CA*d0Kl� �ϴj�?{hd�o��щ�i 7֩�����I=I
��!);�N� %=�]�l5Na�GB���wS�D%J�R�i�Rn���<�'�VݏZ�1gm��4��˙_nm����勐��L��b����/<�2�����b����$�w�y)|�z��
�e�]��+�5��,�rm���$gv�:�:�]V��v�F.�6Pl2�a����m]��B�K7��wD�����}�{��l��O�}g� Etj����<��>E/����2�[N��	aٔ�}���ҽ7r7JΏȃ���7�T6T��}�fփds��a������u�wҲ���K�#��[,Q���5
46����|��jl����G�B����F�pF�$;~�gVS���|�k�E���μ����*�gh�$��E�M�xg�����C=G4(��u߸�{JW�߅�����Ld>�v�3=�'z۱�ڊ�5^;|�����0�A
H�+,V�y�ƅ<����]��շz�ވ�I�,�V��0�;8c�����X����q�Z���e��
��S���Խ��-� �=�O}c�������V�O��t<N�u]�h��Mex��CV(�;��j�W��Og��t-�0]YR��[[[^zx�Yx��h��w<��e��;�g����ew&�rh�]�5����G0V�p��5��ԯ2�.�����xn>��x��-e���������6[F�ƪE��Y�H�>4���n^�_�i�C~�]�qv����
�<��1oM�jI��]3��1�
������y%KƁh$!�hl�4"</d�tQ�A��QȘʯ�Qn1ϥ�����_�u.���L�
( 1�Inm�6u�AiY�]��:��8�9D���W3�:\�È��ֵ�[�c�AP���*�-���f΅#BK�)gL���f��z�m�/s-T�E�G��W5ܱ�f�j�hK�����ͭ9{٦�pṽt띖k.,�VC=S�����-�t���x��g�!E����d���:6E��S�B��t*�cY�1�V���gX��L+�i�V)k��3ln��Y]3��ۻ��	Tm}�!� *X�˭MV9N�>��t.���>,��b����\w6#�æ�4��ixr��z�����fM��n�Qʗ�WY.�����B>|�1��;��5]C/Xz�0�[��[7d�U�v��<i��L�7���Չ�jl���`��Y�5��C��
�_dep8������'X.�N˾��l�a։Bl��~WM=�v����γ���7���0���25˺�����\���d���]wn�޾8p��l�wN��XФ�'sfx����9�wP��C{+k��S	�ݽ駎h�{�-�|�N^r5؛keNwt�V
@i��2G�.���~���.q�ں��{X�88,���o�
gU�'/�9�s��{�]��R�Gy������)[�V�[�u�x�A������N��Wc�p���=v.�h�(h��Z�0�ُ.�,���ž�r����i�C�t��X�f��I֝����
�|/��A��eM㷖�!��ݤ�#���k��~t����ݏ��׼y�$f�fM���ZՔ�a�h��m�-Pt�up讦=^��0"ǣ��G��ͮw%�z=�=�x�2uY�o�ʃÙ�k���껬\�֔�舏�no�DJ@I��i&ϫ{[��n]XU�52��N��l��w��"�OW�\XΆRa׌pZ$��e���N�����|\n��a��a�������x�Ou���ݵ+�]z]+�F��G�0�-6U�N�BSF���{��ye�u,��7��KIT����(�^�n>q�Pt�,:�(�I�]������/�xL�]8�ؼV�S�ebŅ>ō�[��;ڲ��/�P;G;̦�E�)�{�>�\�Q-�B�>?@*�c Qhӫ�ss��^�?5H_>�٨�u��n�޾��ӛ��E����o�#�V��3#`��	\¤�U4�%�2sY�^��H��6���;���}�ǉ^������ď�)�_x��T���4�̉���^'=FZ=�K���V�ı�S�]��R�P;���CH'��;;WU���CA�,ԓ�O3�(�g��م�d���3N8�$�
8��_M�w����*�&k�P�sAä��N4O{_^=��KKQ����ꥉ���u���[J��
�X^�M�Pm*/9����Rp��L���u�6�u��M�{F�fShBĉ2�J7$gd���k�'�Z��-慻�l0�^�aL���I�x�+PoK�䙳�PG)��ooK�wg���q!�����-��DC����O/�o�@f^=��ci���Sʵ�
8��Ś�̙�S:�]�L�`s/��u��|V4�q}^���t�4
I6f�d.���Qy�XD�Y�&K9<�Z�e�t��]�S��6���E�9pм�vй�3_	Ф��M�kv,N��"�L�۝<����GK�/�}���,X$�~�Ǻ
���ƨm�	_�(������Ma�j����k �K 6�c�V6��]�tZ �B�]O"	��t!���{��ʅ�����zQ$OaV*g�=��|
��[S^+��������ߕ�MPڅYVY�pk��Y�έ�m�I�$'/Q�$
�a��e���Z"���/!߭X�FTǆ�z#5���a��TY���M�7nH3͹���I͒䫴�{r8q��t�v�,����Jh��������{���x��x������3s2�I��ё�WZ@L��W���]��V��\]1��%ݮM�P�v��P<m�U���1�u�Ǯ8�r���7���q�=��3MRʙ��^:epW.���<u���<��ʡR]1[vu�`�,j��Y�u���[�rS�S�(�]�=�QH����n�һ��Z¹���ա�������}w���x]��TJۜoIw��M�fL9���]%�@rռ��t3����zХ�ǼZl����06�������:WT�ZZy���e	Һ�k7��[�=�O��c,�-��`�YX�ѣ����e{D;�[��6{Bk��M�I,#5��$�1�5�V#U�sg¨�)�7oVN�J�;s<�1픣�|��ʹ7��� 9Q�<,�A��y����L �5^:e_j�6�SN���!QU�ω�yghL�'�jч�SZ��;�ʝ�Q!�K�E��>���"�� 	�X�8�k% 8������ֽ�skY�x�ycWe4y�`������]<�ͳw��y��2�Z:�Հ�<,̶,5�cWB����ҳ�����8&�à&�,�X�e5��1v$���xk�A��̴W��!#լ��Ӱ.�/lZ�f���փ�W
�U��}�\�F�����I&�9��}�3!��|�[��*+I���=y��R�T��mB��O�7��n�P�#9s�F�[%<��g��f���N���xU���Z�O��^� ��:�t�׼���qڽ���}'J@+�{"Y�%�"��Q���yQ�Y�/�2Z�-���I��K�^�A�E;���U�>�6V˞o�w���]/+;X�Y��r�>�$qh��(�����5�r�w��b�l��/������lHD};+���s7�oc��^&߾"oiדV�;;���W����*�
J�e��crHezfdg��\%	��b�w���@�%�7��/�n��>Rq�>�*+��/K3�|9��f��hK�7��v�-Uu��HǄb;��n��-�p�^.�a��)�u��w���ے֤��$pJ��xo5=������^���:�{�A|sE�ﰿ���~��޹oƌZ�h�V�ym�͂��j����ҽ~�����f�#�����k|�E�A���V簻y�.7TB�mh���&���X���=�O�[B��e^�W��\���3f���>�4�U��4N�ܗ�=v4]�͇�#��ڱ�.����aᘵ/�U�B����zy+[Z�-�����C�v�H�{'y��;݋H�y�C��P*P0\���d_�c/A7�=t�f�z�^�9^���S�]�,0�
���n��B����]�W�XtBi�i���VC{�ý��ı��dd%�C��fP���<S�;V�;����*Ź*�ś�P�ƶ�Q0`�h�����S����nV�M�R��z
��y�g;B���'LF\�H�)�ݜ�q�;=ͱ����=�3Gm�\���Eb�����lD����&j�3rt��UB�#��(Qd��fy�Zܭ�Y�sss��q����Ep�iwk����B/Ɍ���������{��љm�o1<�mP�ER�E��tcw\��F)<�՛˓\;ff�/o޹o������h~��@�qy
�W��s,:[6�{���,�-4� %��a4�����(eJ���ڳ#ip���{��	��U����1���fֺF�+���AgN�v�6.u[�����r`W
0Jv�t˫��'1áVA��r'Ē���uo'�M�W>�m�f�Xx�9���^׸-�a�O����I��)��E�?=�{�ΒDb��Zٷ�s"˹\ ��G>��n�+�7�=wI}��,�>���X��g���C5����m���fQ�&�3��1�.��]4���W��u�]��O9��2�R3���3�<��y�h�|��i��������7u���ߗz�z�{��nʚ�����BJI�H-��k6s"y]�\����^���H�O{�Osn{Obl�o�җ�^�YB���r{Ӏ&#�ǯ�{��(TH��4����^T|{+
��II����;�s���r�A��RC����Z��3�>ܟuab����t��4Ji0�L��Wn
����
޴�4����ح���}�[U�N�ʘvMd�;o�j�سa=[�f�4���ӱ��N=���\$BDR8�=��p�0��<Wi��] �����`m�0��G8mr�qS��E��N��C+�Ԋ�a�y�w;ȭ]�tx[Z;*d.�)u.�%՝��k���JC�*������K5A��D���w��ׇ����̦���ռ������"��@�q�\\�\��ݠ|����WN�.�2٣�����Wh�GJ�ͦ�a/Uљں��Rˠ�ac��vZZ�8���oY�D��89*P"���gb�ܽ�������@h�6�r�`fRZJ����9�W:�j!�9p�u�����#`-���{t����W]n�v;w�U��|��Y&���N��9���2v��0��0�shלj66�;��w�t7��A�*! D�� RE��~k�.X.�������2�@�w8q��B b�x��ۮļ�Ýz8��� ��@�ĊE0j�
i3�k�y�̫��M}��7
+)�#��=X�f;5��a��&P�k����*|W�t]�{,!8p����QT�A�I���]��o%��L4}��/D�X<�V�v���"�)�x��I'x��+�,9v�=W/=�S��h�YB�E1Ӥ�J�4��Tc����
�Y;N�Zy�>��tEk�c<b�G^�۝~n�,���/n�F���"5aivkÂ&�?�Il����� �q^�Z�'�/�	�7,|�5��\">�w$<􆘼��U6���w{~�6���z
	k,�ӭSv�۷o-�w>t��b�s+����]����e�E�(��	�4S^��s�l�ڕ�X�A1�87uP�Q(/��1�]b�=KaLc@�E-�w½�׏�)^b�#8�@�J"��� ����;��|�j�R�.��38cÁhTd�3�f�����j\T"�g-U��;OLnű�����(��1��l5��%���f[��f֞4�o��Y���5���ң�o�(g��aʛ�q��5���>�@��	p���:K<h���U�2�p��R:����n�?���?��+�8u�n�[^fo:�۬�Pt����MS;���çK��w��^r�o�J�E~r���cc}��9i���"~�6���Y(�M���,�;����&@%�j�j}�0�y4q�2�����"��2M����D�#��a�s$\ߍ$��9���d����(���C_�|z��t�BΎ�n� ��`HA6m��Z:�v���eE���Y2�3y���
b�^+���b<�ߒ���gf,�;A�3o���v���i)��Յ#�2d��[��V5[\����������ԚUξ�-��<Ĥ�o�K^�hn��3�w��y��/{�u/:	��#/U?��㈚ay�8��O}���g���z�L83�K|���Ͱ,���V0}6P�n�]��+��X��M�f����D�k`�*�(��)W���rǄ,��<kY�����]��B��9�*�|���y�����f��o��קcC��z�<b�&�PH��-���%��I;*fP܆�.	�گR�c���妽��k��G��;��ݯh���s#��z���w�v4o!e h�`Xt
)4wj���&�]��+E�bh�Cے,����X/�n����y��,Z���9As�f��$��	�Z)�DK(#�N01pc]�� ::3��J�Ƥ�	�7-��GB&�4�L))�S�B�oH�pm�c��J\֪���:��z�2K�0藕��T�M1X�y_�H,��n�.�"��@�V��(,���BB�2C`�� �+�:v�U��6��p���*�G�:���/{�@���T��6�W*~0:V�8�6ƘP���]D�E f<��^��j��;�{;��#;��2����C<}��)~)�G͐�Y�TH��TP�)6�F�j\�G+3�ͱ�px���i�>Zu�%�\�iS<���ّR'ع�Eֵ��爃sҬ��W�e��x��]�J�ܶ�.Qܙ�n+'k-}ٗ�˝X��$�ɶ�ޅm���2��N����3�Z�a�l^n�Ow�� AP�<�5�j{Ƞ�&�͉V�����\�����'��[����{��7z-]ݗ~�3bϾO��,�U��|���Ts ��R���.rv7X笠���)�Ü2�u�&�p��)�HN:Xf�QtM��sT��,�?���Ef�S�e-�ݚ�����y=]װ��מ<����0	Ql>��x�YWe7�! :S �[%6=�QO���Ƽw���`���K��`/��j��!f;���3:���.���z�נ�JwO�y����ȕ����sv��7x2	�q�0���[2�Ot�Ŋ�P}��f��l�A3a:�Ù���@���.j��ok����AG�M0�i�Z�N�Y�oY��E7G!�.lr����ى�7V�wZ}�z{]V됺�:Ҙ�=�ß���f9��:( �!6�A7[�Ժ����ԮZ9�E�
�3icX��Bf�r^t�T/_��I�e��V�b��)�z����k�5�vz�Y[�7Ku�Z���Ui���n��ޗF
T���௯�*�R�����Y�:�����FK㳹A��"�b�ˏ�Ō��n1&�ѽ��;��;�9��k��VJ�{&̀�\�*�<-`B�_J�1I�u��=ʞ*Q^���]M�}Vq凃v �l���t�tZ�&��Փ(�;BPw(��	�`�<�����#j�E�c�!b�:������o�&�E�2n��;U��_�
\��R��b=o��u�\6�}�:���Y�-� Hi�]���#m��\���)��Vejj���ͱ�㲳W9�N�W��8�T����Fq]ر5j�VNF��
�eԚʎr�Z�(��%����ĵ�
��{tmn��5Ǚw�U�c�y+ڠ�e{����Ĳ�_m�[�o�[�N�^o9��'^�,Xk�"��qCV�P���c[�ގ�����[�v�G�9w=g m[5�\�T`*oh u�Y��χ-���R[�G�̡�ne�f����O4�b����~R��[V���+��<ƅ�1C���,�5�������߆��OP�ٟYm9�U�F<��ͣ˞�E��N���n��gSߒ-��ʸC��V�	��N�P}�b�>���ghǈ�Ͱ/k��1VwA�A�������N��un���`�{H3� s�n:,��^J�8hn+��\�}�j�236ol�h3���{ܝu���}[J��Q���L��c'^Axj�:�
j�f���ޒ��47D� ���à8�]C6��yY�pd������m���k`�pꩉ�9ԡT�ϵ�mS�52s㮵FŌ��|�O"�7z�=L]mp�v۲��ó���:1�k-�\m`�ybl%�m�.^+v���Y�)�ra�(6�sWc`���r��Sk�6l��-��[���&jekP�7M"���K�i,9����N�nݚ�[�X�`�b���v3�*ێ#X)�LW2�۬�=�Mj3�V�5�Qf��t2�M6�E:�W�X�/�T�:^uԣ�S� �R��gl�H���l�s	���� �B�HmY�/2�,t9�ɢ�W�ctWW&��g��%��tyjʣc��a�)3��)��|�wf62v'Q]�As`zwa�K�`Bl
�1�vV4ۆ�x�ޱ�rv����@�<㣀�;7<v��/c��j��9|�}��׮/m׳=�%�Gh�8�V�:+[B�R�+0��2���%K�c�mч5q�U�D��xI�x-�q��&p�FS�=S8ON����l��i#`N��Hd��l�s���<T�UՒ��W��Q�^�[pq�[���i�����\����]��Κv��Xx�ay0��q�R�b� �u��7Y�XG:d�8�2���lIT�w`�E����9�$\t��+{ksz��z���w�:�O �֞6�q>��5f�8+�[���lp�7]���
�
��v;t's֠��s��wW�쩚�d�l�!O9M����p'�Ej}�`��^6QKF+��/GP�L��F����]��J뮭��ռ�.l�Kg����D��P큋���[��9���!�����4;�z��}��9zI�)ؒ4G��G5��E#6i6`���4�-ѱ����n3pmk'�c�����Jt�l&mv{\8�v�s:�.&��z�k.,�x�������\$�e��#S5�F8���&�ۇ��m�OS˜է�����
����`�oF����3tvu�ڶs֚d1j"���uփ��槥��c��۟gm��/p�d�{m�]X|*���{&2����ft�R�����i2�����]R�e!w�z���c�n;[��ܝ�=���3�a�Z���ݸ\l$m��D0e��l��+@��6&�VD�ʑ��vr�U�s�H��Z'�y�J25sBK�lZÓUK�)�ͬ�\MW�z��@�v���z��]�P��u�o$k���J�ƻv��}*�ktu��q�]hɏ񶞍�u��!潢��v��o��~zp�q�Ee�ԦM��]��Xm4ӝ�h�A�:�k^'��Ň\[MN��D�7b�z�X��Y�6z�v���Ok���C0�f���>g���l�ۻ�sRG�T�
�S��	��׎��;�c�L����P����PkW�]f�Hץ�c�]㶪Y�=� +պ�o/;ީ�C��:�����o�N�m����ݲ(�KyἨ&��-dG1j����R��Jޓ�{ O����y��Jo�}UeR2�Ҧ���u������$�!�o1Ei�{);���U�vV��_v�.oPe���~���^ɕ�6�QJ
���T]2B��lfmF��g^vyE��n$��]N<�ŷ�M����k<�4z�@�����7�}]�CjK�����zv���������$��l�ǟ+�,l��ڤ,��&z��i��:-خ���݋
)�i�@��#ƞ���|/���$��P!<�)���us�w����A$ѱt�����z�����rCآ��υ{④�M��i��=\��V��H�������D������8��hc�c���z�3z^gTF2/�Z�ƣ��c6
�i.;)ٸ��9B���M��)[ySsl嚀�ܼ�q�1C��n��������=��}�n��}�*(i,��ǝ�r(���"�%-�FA"a���?��&��V��8�d�Y�繮�z��:�jL�Iw�����O=��Ӗ������aE�E�S��$�`����m��m�4�U&\�h����g�%��^{敺�@�ӈGҕ����r��7���~܀��"��F�kqh�E�re��nU-iT��y�Ց�Z�a���o���ga�;��x6B��q{e�Z��č,N�h��3��
)y&B�L&>-�Ha|��Y�4ԩ�)!�B:39�h2�O�n��:���t� #A��):�_e4��؅�gP��rSV�;�E_b+\I�Z��vgM��U�B� SL�[!����E%���E7�9ú0gj��a�a�M��:�s����yKt-�"yߦ^A�m��]HwF7*w,ۥ��/�R �A�m��V	����+�L��%Ѣ�m(M�ý��[�s�t����4�N�$ҫFkʻXc�;	�ϩ��̼�5�i2�� ��^�Xv���4>J���9g�n߅��[=K�#Z(��b�|��8Z�R+X��"m3�]�N���p*��w2����-D@2�ɕ��9z��''y�4wV�R���Β��Zˊ���ޅ���"�T���=���k��fn�(�)^E|v���J�I�-��TKg����}}b�`'%5D�P^l��7/Vx���<$��K�)��K�ϰ�ۖ1�u]�.4���&�msX���IeLBY��2���6��7�c�﮷ٯS��9&�.y0����^-��)��R�m���u C���jվȾUt�!S`�Kl�m.���&�G��Ӊ1�8�1�=ZwE��g��3��Ȑu�+�ݫ�k������R`ٚ7q^�,���i�RR2G0ܐD�4�@%�ᮎ�EI���\���Q�yK��=�R�W>�]�f���N�^�덎{Yjć�A�U�a@���/�9�.�|�h�2����L~8�n�h1J7�����(WJ�Ɂ�=���́�-W�u������v�z9ٗC�`us���{���z���ߴIe�('[���.�F�Ҵ�����k�����7#���}�oF��D�<	h Q@��L"[�c'���nn�ډy!�V0a�:�ש	;^�4�A��R�R�qmԖ̸(���m=&X/���痢��K����;,���	�h.��33��	�f��.͸�M��m*��x��h���A6B���)�(�S����fY�E��N�X��Ck�Z%t�X���ޜ�s�{��&wjy,<�-���n�d[{N ёHoͶ!6��NtϲY�[@]��{.���.�CF<�5��hro����f�_������;�R���d=$���[�F�(% �ʥg�S|O��{�4V�z:�B&G����-������n�Gpɘ��U���{��oA�o���T�#��X<A}	4X���pk�^���ٷ�0(�3L��{\m��OI�}��^���ץޜp�>W�KN��g���І�ֹ��jL&&R�T%��a\��q��_r�g9���owA9�of��p7캔|y��z/a�
dA�+�yR�Q���+����}�k�-y7n�Q�c�AX/7����㨨����YB�0/g ��V7Hq�5��JO��(c4+��T�헗��� '+I�B�z��5Ӄ�I� �^m[P[Z�.�X�<�9��#cVX��p�=f\����npy�޷a��,q��"�����)f�[�����pS��j���;�͌���Z�9۫��x�Uۊl��w%Ƶ��*po��hɹ�5�ڞ#xn0�;T3�8�mvB��ݻ>��^���Z���\ʺm
�3�(��:䄲�Gu%5d�u����kƱ�#��d�КmY���7=GQ�=�0n뷯6j�te���?^�ГFz���?7�O<�l�u��iL��Q���	����x.��:ځ��Q
q�y�;�g���gؽ/q��,�:��eV��ʏ���t�wA�43�<~9�f WVX)t���%�y�%� �$&�d���;���L��Q{�,� �>V�pՆx���EČ�Yӽ�Ӯ�x��������N�3�ӓ"ג, �-��L�ϝ,�Ӻ��e���Wj�KF�sk0n\xh	/+'r�o17�W�7Z	7D�u��R�g(f̉I:x:qe$W�zg�~�K�L Y)����'{��U��)A���ځC]��7�4s�_v�:���鹴%K��Q_��ټ�]f�M(���}1`�u::�HPH"����5��4�^8%tb�j�XGMZi����f[��X�QPl�E&�H;��ӌ{6��̬��ss="�!�t��=k����1�]�J�u}�}V3��Ǚ��'�Q�,��fD�eHL�9�&{�gy�ދ���5/�B=��vf�H9Mn. V�.��\e��rjU� ����כ]}ڇn����Oy�ս;��wue�T�:�k��3;�����
Ly�h\���[��0!�W�?���5�jx�g���LS�(G�<^e\��g�A�h/C�>��mPa�0c�<��|����}��mp�G�h��ꓺl�;8�vq<	v���t7���g���.M�*�I<�����<y�!ч��A&)IH��&'��AȐX1��I���p�6��ut9�q��k4��[RW}Q�
��{�{F��WU�)K�w_��{�r�}��Z|T��&�"�c ��p|��f��dt�1��$tԶP�8�
����g���¾�|�h|��z��o���#���~�7n&�㎲�/�,�o6�g�|��Eж]	+v�Ÿ��Pv��M*Wg�.�n��ƨ�2��"ͬ6�@�0�X���w�������=�>�~��B�* ����w��u}��������w*�G��ey�C�f�^��P��a`ˍ��|�����2ovJ����x.��ȫ�z�%N0w}����Bhū�Ś�F���y����-/s/�0j�h(xfU�<���:��qڑ�%��BϢȬ�=�=έ�@Rx�V���f��C{^��(q��3%�+"�{���l���,za��pcG���\.��#]0�كs's���]�i
�\���ɻ�Ŏ���DQFhOl����D2E사U�B���;����j�r���.���t�q���q�vgG�W�i���w�+0It����{D]�
��Vj~f@�;��$(��d{�E��C�;ڗ�C\�Exi������`h��h&NΠ�(ٜ�x��ټQ����B��<7��fW}����2���s�z�XWӸM�>����P��25���U���c���b���&��Tr�llr�����Nmv����7l��j��ܖ�l}�C����>��������E�K����#9v�N�<�a������F�lUN�+���zM�)����%���m1
6�'�����1ƚ^�l�(`�/�T�n&i4�����=)U��a  ���3������3�ƪךP� o��j��x��
!����,u��C�$%7��OF���C��	�,h��胫2� g����m�:�ȏ/Og�ol�W
E6w{�S��
�g���p_�!�B�Û(#�6���	���K�U.⡇¬}|~����
���j<���'�]m���A�����2z-��;B���1C�پ���8�����I
'��N�H6��6�V;`0��Pn�����=��X�8�t�.����ѯ��ǣpfk�Z1gq�Â�#�&Ke1��W�oġS2��*��+�²��7�=l�����_T���G(��&��>�ES]/P���=}M9are�p�SaX��Q�TJl=p�g�����u�X��"���͈^6��XI�-���,����?<�����jd�+�RA�g9����w����U��r��"k�VWYC��Q咹�2m��&f����$) iý-��>��)�X*{4{d]�~{���h�������¨������=2Y�L�c�WW���*�bM�B�B�ef�''{sM�'x-ʰè������u�(�y��)�p�}�E᭩��ހ�EKnS4�
�|�dz��0D�a7A&���Ɗ�j���a8R�vP��xo=�%A+�bj����-���$��l%�L���0HW+#M��o���~��<_.+��ƩѤJl�H�X5QZB����^_h���<�"�=��ޔ�U��r*��@c�0���!����5M��V=�KZH����*�g� �'I<Gy�b�
~����U�F���ɮޣǮ�߅��=�>תc�V�q$����Y9��KUP��P;jk�ݢ�CW�^@��k���p�sS��Ηg�+�g�>���y�5��<y�J��v���up��I�Ѝ-3��]�@Q�m��t��d�pd��o��y'�$��^�|�ƇV��:�=kn����z8�\���A��۵�6�oc�sc�	�{ld�=p�ח�	8�i;�'
�u�K�/g/�����k�}�x.9���������9�b��m�eo&͂4e֨خ������)5���z�\u��QtA�:�<���hsuκ�Oeڊ�w�
%�)x�"~�WX1���*y=6H#d|@�ý�J�'e�^��wc,/:=��2��w�n�a�ԍ�[0���<A}GL����Ӛ����w����`7M4z%D�i>�~Z���]�3;��Seh���|�T�;�u�H�|$8S,8TR��0j��3�8�m�f�ȫuHN���V������;�m��4D�{8�&{Ƶ]$�Ws �����iE�O�����A�\8M��V-��� qݧ�<Е`�l����	
��g�~����VE���QK�mz-�4ݭ��^�ȍ���C��ظ`�,���C7k+n�|{^{�ہ-E��/]���:A��(������0��4��(��D8�W�k��(ZyY=x4i�D�.�/{���N�C�\��К�JF�Ʋ꠵���=I�S�;o��>�8��]]��S h�R�Lm�>:��tEAU����+��f����o5��M�B����9��<#�!�8��*���sVv!�6�3��I|a!D�-�f��1_�PH���1A�$X#�[N����}E�:�]i%�˧�����7m�P�\��(�K1��$��7u �[y �Ӛk���ʺ����y^հ��m�|�w��p0��؀X�i��T���2¼ |�+�XB�K�{�Y��=�-b�8��4ap�� ��AH2)��^����w���G:���]f�B��N�~�������N��q���i��U4 a�*�[��ϣ�3����:�>�)P��rǂ%��PI"p����Y�����������z����`����H*�K$�׃L����t����6���P�w:�s{+��P}~��$\'�gפz���J^��"H ��9� ��;��_6�)Vo�^�88I�z${� �M��P���
$�y&^�b��g#��ATE��'}݉&�6㳞(�vM5��7�ʹ�Ӄ��v[�,����0.�B;���u��5[�߯�o+�guY����PdQH��!���,p��Wd>_S�݃��d���.<��¡�(�]��'ئ�+�R����8��b@��R*�s9uy�d�t#WZG���au|2�@PG��� �-~�_q=��]1�^��lU�yw�x��x���)�54ް�|�H�6ۃ+M)�L��� ���Jj�}� �� E�����aB������k�H�T���Pǘ4�Ĺ�k)�	����ͽ���]����`\�]ksA�v(�U�|č<�w,�����[[,���tOR!d�{;�O���٣r��ro]�s'�.�#�W}3��a��-1γ0��i{׎!n�͸u�^����o3�R�>�u�3�Rp ��-���a�ξ�JL:��ϰCCis�x��N]��e���L��mj��_&����A���1';ox��݂ U��L�w�y�O���<���{�I��2Xy�V�ٜ�fm7�'ֳ�kj��t����'|�gKF�p���2	�gLX��Ёշf[���f�U��K�&������]��Ƀl���lQI�9m�����&u���L��3X��cpZ��:Ǣ�
٪��N�b֎�X#A��8�B 7��]���g!3#Iu���WS�-�h�j�D�u�d1�Lu�+����7b���ΣH޷�S�9#_Um=�������Y����N�no��h��t�;9ō��0���:b��	r��,��a���2���N���i��1��l�ۥ2f��x���~"�O��0�ڙ~(�'G*�P!���X�fG�4C'e�&͘vb�\�7��k���Ѕ3/N��Ϻ�7�*���Y���˴��ٽZ7�+2�悪.'9T=te��6w��[B=W���p�;���MY�̾՗��þᴳ-�]FV�z����������u�hS�ˎ�v��U565.��v��oh������q`�7�s��#(o�tov�
�s�,M�e������1o��hU��{�
�S��	oed<>�K}��h��C솀�?D�����A�R.E�5Ңb��:oB|w����.=������r���5�����j|��Ek�+j^;�oN�� {�W{���j�=6�MtK����2�p	���˕�D�Q�␒�U��Ȇ�5��h���|���q"ګ �t�d�5�#]�;�3�����G�Ƞ�����3�49rJ�!xuw��@|�X&���ID�Y�M6���n�7o������}���f��	��C	+���Նe�������]d�9��IR3!1"�F����]�A�\�=cr��D�B�7���^x�P��l1j�v��xk�^��gp@�f�Ut��hC����(�N!L���������c\�a	M�(t�]b�&��I �s<y����-���� ��\�/�}Z@<H���U�C��UV�Ѓ�����{�@l��4��N�-��b�����k�kN���>���-��K)v�Q�r����\�6@�:kM]��L�N^�t�5��a<O�^��!l��ȣ�㬲<�I�(=}�t<��^H�4=�x����/kǶ���3\��
kP0�d4�-��>є�%���d�������	��^j�U>S��\ʤ>�z:U�����YhU���+E����@��;ڃ�;X�.%�*0�Ǝwq�ϙ�Z�����^��N�ҩe�7�ڸVR��M��c��� ��ڈ��M��ɭﾭZ⪊��P�*�T 3U6:O�%����� a F�46�h罂���@��	�f�{��\��Lvb�Q�ʿ����p}���tՐ.GT�ՙ�t-� iȅP�!�Ӥ{ע�7_$�,��Es��JSl>��(�Ti�&H��Τ6��R�\�o��4�
qؐ�M%�k+0c�B�8=[-< Y�1��+<�{:�}���'��2,�f���\�+��x��@������]s�^�׏M5�m�Y}���4&*��!���Y�y�,a2�hFe&�gN�!�<�4L0���D�ҹ<�o;��ZE� 2{{�^
���0�;�<�Dif��iS �
�j�l�:kfi���a:hz�\@M�á���#J	��b����zB�$Y���������ÄS5�1����ԇt��'��ot�8|�B��*��*ذ�5Vz��@a7��`#Cv� ��y�Js���}�sꗖ��\\0����_��x��x�x*j�sy�`a ��ڦG�|}0��F�������l@#A�t42����=��B=��\��C��D����d�dG�4�HS5�� ���c���lWH�-@C�X*�b��diha�(|xP����\>�Ъ�f�"��� �xn�`i Y�����ű�W���zF�R g#� !��!Ub���t�{k�W�8��ӵ�P�;�݁�+�c�O;v���a=yz�S�Gtӄ_1�F���N�Ĕe,}�[�Lp�J��%z�3K¨�9�R�eͷ.;xЖ��%ז�p��ܺa�;���Z�ZM�qx���4E���rn�?b��EX���f5e�YFYYXҌ.ґK���m�ԁr�^2��6�E�nW�s�g�j��1��89�ϻT�Nɋ(���q># �p�h����*��M�刈���٘�csB���3�dUp�n�n��|���VݮC�ܮ�S�v.���g�:f��u���x5�U�)��q]����;^3֪3�Z݄�ǃv�L̗ .��flY��3$GH��] �D�9�כ��552:hCj�_�x��I!ևHt N 9v`��y_O<�@{:��(۪�3�V0�Q�2	"^ֺ|�j�����4���8ha"��@u7}� .�D�Ձ=�b�Dt��ↇq�i5Ӥ��`��T"��&ﮙ��>� ��@�/ʀ������`K��WR̝�y��t���k@�L�!L�Ћ�{,:+[nM�P�� �@m��;����3_MYA��5<�ʼ~v�WT����R��o���oć\>�>�?V�{�`B�i 2����Y!d
>�^����%�J����f�#��r��f�,I82�#��U����;��D��y�w�p�������4��#Z@�۬ Y�!���]#A 2�A�*D(�ٞ9A�5�"*b�M�����pG�����5*��5�5������	L&� ԍ]4'<��=$�	��\�h��&Цh0@dS5�����G���ZE#B��gHj����] q
����a w��p��3}�tHHC5؄kHQ�w��罫qvb���/[��� X�J�_�$�M�!ԣ+њ�2�SR569F◣������G���L.Ķ��I��Ĥ��D�=9��`V�l� x��DB ��훠4�u��a�x� N*�7�W�g�=`���ݤ9;BW�E��K���yn�5����`�Rl��m8���]��CE�A��"�ݧZ=�sv�b����̴'�%�W�������|�M֬yI���b���ag������8�j�Yv5�\�|0�3u��K��������VhF�}<�,�h�)�ԩ�@im��+�4��CP�MD"�=~�`x�h��r���;���#Ư8�i��9؂�a#�J)#R�p`�t�3AyUB;�%f��b�m�P� �^!��b���ц�b�E����@}JT7��>�`x��d@gƂ56ݤ 	���a$�L5�V}Y0���_���3&L�7 �4�h-i\�.z\�m�D�<"�*����5�Q�Mj���іF?g��p� r HF�a@���h�5�*�<@[;�!�48w�7C�@&G�"�B,��3���h������EB'�����+��#)�h
��.��]�#܍�oq^�����U��EA�H�5K�w��j�H���p��-��9w������=�(����T`����V�{�8�zU�ї�n��x�%v��x���キ�5Z�0�hsb�q,pS7[��D쟁�hPdv*��Y�)�����PF��d�3�WC���@� t�}Bϻ�t��d#���dt��6F�� {�4�8@�dS#��a�F���-$�~�%��CH���(Y����GG
pE
��֎�G~]��(l}���)���Y<6��+M"O�
 iF��^���:��֨. ���y���9�w�\�IM������@o�9��^$�T
�8�i=�BȳUu�L��npg��i!�&��P��aK�(1Y`�BY
���w��&�*���txە�����m��� r�e�>[=La*[̀�� ��s&�,����G]�w�0E���,ŝ���G;p��b�N�,��M����P�#Mڧf�r�1�{�����8�ni@dS����K�o������=U��f�����u:�QH�F��d�! �壘�S\~"�z��0��� E՜6+�i�|A���6>�7*T�K�=^���ג����zQ 3�#�������l�yE�٣uǓ�8�������ϳ�� e|P��>�	�����5����f��æj���qd_����Mi�� Y��+ss4��4�K m�vhYz��VG��i���5�ܔ��n1�3\��C�_^����Y�8\�֗�^�,[�y؃�Kf��Yr�U����vI�L��x����a�xh2 Z�5R�� {:��~D]��2{P9�T�;#����r��A��������LN�G>�鼘�1&$���>�m�,�sZ� �T�m����|�-�&!�Ƚ��m��U�(Gʅ�3b�d�0�"��U�����,�3+�( �h ��t]�������R�C�0�<EL�֋$�8a��nCtj��+4 ��:id ���9�uXk�gHؙ���C���`%�,��}v���_@�A�|�����n�雌hY�Ϊa;3<lV��@ꡮ�����a��S
"��H�a�4���p���$Q�>��G.w��9�Y}�r�ՑP�~���i v.�
��	�xBW�.���F$� a�h���Gڟ_�̜r^��QQf5� ���[!�ۏ*�p��/������.E�ٮ]Z��`�laB�[ͬ�Ǽ������w�lt��5l���5��+�+Zy�CUv�s��tJr��JLk�{����hi�e�j��Z�^�����n� ��4���vxح�L2+�M���S�Vt߸,i���ІqV��g�$)tߟ�,oZ)F�!J����卜�M�Xj��lG)�*M��u$R��H�Pt�V�퍋���d��3H�ZFw�-hiȤhS�@;~�v7
 Y��&Ml��<��/�Z��׷���� /&!�����o�<Jp���/޺x�E�㈸bQ�t<F����)f͗L�~�q��[�>�����UsZ"��#�o��t3��4Ր=�c�j���Cx��U�|��Urs��}����{�� ���z�bI�w���R���f�D��4�T#÷���e��	ea�d3O�^�b�� �{{Ї4D�+��g�;�l1��k��i^�j�Ixus��顡��H�_�]kQ/���N����aψ�P����U���:t"&�Ep�΋8yw�V烬5f��3�0BW{-*F�ȫ��W$��,;��i�GUE/9�y��v�*���|���!�*K��{��a��$�� MH2�a�BWi�����5x#���P�x��# �\sM��r=ns��&����C��i��lx�&sU�����+�PD=�jz.�&���A� ]�}�<�4��� ��޸&A�]~���f�4@�Ҏ>Ǐ�N��h6;��ז��ɛ�ЉWY�a)_�կ�ss.)�,��sȫ����M[vZԣL䙛�h�kq�ٴ��;L�ּ��C����÷o��x��ۭ��9rvܰ�er��R�-�u���Ɏ�{���R���c�)K �̩���4e9�`��jRb����ʡeh�ƣ�Q����r���{�х.M3+i��U�x#��Iq�n��Џ)�K�q���9&e�BY]�bb����e���dA����Ic�v�u�i�E��;-�m��j�㤂�p��2G�x-�L�nR��(Pmk�]��Qh�Q�p}Cا�xkک����n�)<cրF�P������WmXkE0��U��x_� |��Up�>`.1[;x.��젍Q�	�P�P�4���k��E�p�8@�dU���n�n����E�dҴ����Ό5}>}#qP�Y��x󊀜AqB0���{���\00Դ!��x��1��P�l<�d☼�T�t�|g8�K-���06���d���$�����`Ύf�4:uu0�U�@���P�h �<���}{���.Џ�Y�3��׽��gP.m��a��RXx@2���c�w�c�QE q�$wC1V�4!�y��ݽ�;� 2	� k�7E�0�����N�!{��t�C<"�	�U-��!��!ѡ�1�;�+��@�;I%V��lY Y�1W,�9~;��\	����w<��=f9zII_z���4A������u�V��u
�;�uP��ȫ�ŚF�4=��`��c= B�MWH���6���E"ԇ�X�8{�����2 ��7]���<�V��G�:uTK	���@�X�lxU�H[u��-�b�@m�ܟ�%'���C^��=�uXFs��,�UA]dat���:@�г"�x�7���o��{��'������+H��4W%wxli@g�U2��Y����i��	E7l�V�������A�����]h>?(��w�S+rߕ�m1&ؒ��,�R���ٔ]-[/�zܿ���W^�{�h��q�7��iM��w#�Mv�X����¡��grðN����������h F��C��;ܠ\~��]�یjo�Y��N�?�d�^�t�F��Z�ܚ�@a�3� �dA��ຑP�u��l�VB�Y�<w*��?!�3=��^x&{n{��1�P"�Ѡ�A�B��}��nJ��@�Da�doy�ɑ�¢i��Q�pEi�0���zO>q��AU�N_`�+�*e��c�
���;��@�U� 0՟\b���f�*��P�W|N�m��M���>W�@a!H�"mߥx���E��!���E�kh^�C�ZF�o��Zhi��B(�7��o�3��'/���#0��3��b��!瘨G��N����<��R�("Uԩ��=ַc}�G�zޖ�%�ؒF0�$����>�+�C�Y��:�(����S�^}[�nx��)6�n��A�Y�Q�����<xA�.�^>k ���n�����2�Wgs�7@�OYk��ok��P�^j����%���U���Ǟs����;·�Άv�I��|�?���P���b��1���A�_)H�w�4� af�;<lW��OOb�(G��T���w(K�VEY��|������16��dp����ע��]Q�Z �\.B�7D�"����R6Ew��4��W�dA8��vAm���>�"�C�>�
�R�ڥ�<�8v
s%��Rھ��\�xf��%t�����uhuԡ�����e:�E��z/weM�9�8f���dy�&�ǰP�{o˸P��-*C���0�Ϋ5|�R����\��H�6eApج<<�d ��E�,!���ꮊ׎���n���	�!�;4,�sگ���(2K v*�Ut���T��+�H��F�ە�ϑ$�7\�X4�!7��	�ݾ%���\2�G�@�a��� $n��վ9U���@3Ø�ȿ*K�nxD'G��\S:��xGH�W:���[�����4aUުv�A�d���_R�W2��	��۸)�f�;��w�nIm*h8
nKԱ�(�V'{u=��u�d;Wm�$7Wt��F�y�&n����{�}/16g�sB4}~Ю�&@�P�a��5�n��'�@3O��]����]� ����*�MB��'V4��5M~[�Nʫ"���$x�8hv1Ŋ� Ba8�����|��$9B�w^�O���\�N�p�}URӵX�t�U&���4.$I��$w����23P�i��R��wU�9T[����@�2A�Ԯ�q�_m
I�>�4@�B�PTZ,&�U$.�*�Y�Hz��.���ZB�"~l� .�f��}��b�d�>�z=|H�˾�cVjKvE����}<ls�N�аi�r0H�q�Ha��m�p7����"_xq=�cN /�����Vԑ��f��hxctW���U�e�]�����;��Bb�������z��ګ��.�o�_�=��{wF����
�:�mjŮE������'0��t1lh�rՙJ�aD�i����P˷P���%s�x y�I�	�)��(�����&� tr�U�t��#�ڳGM�7ه'�ύ]�P��o�8�
����{c1>����%,��ngOC�4�A.H5E*� ��A��8�b�7=&e�>��z��`��sηd�l����ι�4P�8�p/6��y�x���{���#h:W��?K @�����21��E����=옩{���*ՐMe��V� �cƤC�������I�cw�O1Ve�����+F����2��x�C��a��.���:_��C�lB:s/4�F��A�KmT�!�P�}���x+��H
̴p���%�Le��m�j�W�#Y^��3s2�.:>�ov��!�>�=J��8��;�,��b��L��II9;ad?��4&�M��������P��y��m<�ةK���b��{QV�oe,��^�o
=��{9ۜ\�6v����z.%�����mWn.�6���ĲYÖ�/�9��'�ŷ���%��|UUU
���*���UW��P���U� ����UH
���U�UUUB���*���UW�UUUB���*���UW��
���U_�UUU
�� UUUP���
���U�*���UR����U`����U UUUP���
���U�UUUB���*���UW�UUU
��@����UZUUU
����e5����P�-� ?�s2}p"����Wkn��*m�gjWv�.-ݝ�.���HC�њ�W,ѻl5R�:���)���]ƶhӮ��j��j6n�h��vO�D@UJ�IR��R�R�UAE"@� ����
DP����T
)D
�)JR�U*S� )E" $%m��}��3��J��ټM�kۅ�����}˶�[�.{���Ԫ�Ϲ�u������ˢ��o5ӛg����}����v�}������Q*|����e^��{�Y�)|l����cYU�[4���پ��{����Ê^zt���P}<�vw����_U��t��}��S������}��홏��IW�o]�W�)Oy>��8���i|r��n�����z��}�޷U�k�W��ָ�[�¹��w�
�(U Q PP*t}7��u޽�gmݻ��Ǿ_5ݰ�ﳠ}�q﷾�sI�ν�(��Z>��0�9Z���!chؾ�C�4��DF��������}Ui��w���u��L�$Eܣ��y�kJ��w��]��_�P}�T�7�_{�|wwZY�G�׆�l=��_}���>�ҁ�<���}������8w����N&T�}羃��p�����c�V�*$ﾨ�J��DR@�$ �҃���>f,�s�}�Jw�>�PWɮ;}h(��>������n۟��/w}���q���w�K,�,�_[f�����}�玕C�뷜z2"�KcY�  >��=��U�
� 8��w��� >� ���c�@zt�>�����c���`�@糠 O`x� N��F Q���P�H
 (�  �� 9� �����r�}�>� �{�  ��Px  	�=������ �`�}�p<@  {�z�*��  H  v {�(�m6��m�}����k��_`�Y�����S_>�{5m�gL֪;ۧ����GWe�/x��{�֞����>����k˻��;w����J�J�Q
��ԉJ
((��QTR"�Uw��5�Ϸ^�kY/yǣ�G�}��N�k����(\��{���U�th������۾C�T������5��>@���kmm����|�����^1�b�Z+[Z��(>@  9��}�  (�w�*�� h ��h q>��� w�7�8�i���7oMW�W/|UW{�O��{�z�5��C����w:��y�`�
����Z�� ����)P  �F$�Rz  h)�14�T� 0�?L��bU  i�T�IQ�F F�4��)���??����_�?������C8���0�g�^������|�w�@P��U��7��(UU
�ڡUB�
��B��UW�(UU
���
UB��P��TU�~>c�cT�n��o��
#N����V�:q[��]d�8|rM=\EYE�p, �����[y#(��EL�#v5��e���U�C(m�0�Y���T,�;�.��'6P[ ��VT� F��z@��%:�,k��!z��ͼvG�P�6)˓rŷ-�N���O4T��v��u�<3C̄�c$D�����9�I�>����%�*諭cI3�th�jj����Te�����y�Y�ުP�/r�N�*���z�Dڌ����9|�I���,Lfc  �f����Zo&��f��S�h71���J���0*��37%	� �̃U	��Љ���,$9��lp�HѼ������m��.�̄�eO�/QKXp�ӵ�q[��̉����K>��hD��S�f���Z�n�NȀ�Mp�1�aF����9W���F��)�C7w"g�1������޽�1�n�Ay��"h�WW�m�N�G6O��b�$Gx�#"b�1e�܎1����+7a����J��1��X�$�[RJl{ �!x���b�7�QS"@i�Ы����U䥤뢬�&�n@l��c�N��.8�7���1�ji�DV赎�&l7Sݟ)�Ud�N�Nd�l�H.�!l��'���o"�r�PMv��}®̧�Z��M��.���#�G��J[uu��a�Gf4Y��'ɉ��	� ��-Xt'���^S)J�����Ee�@+N��nlhJ�8�/rq�R������I���)��0Ś��i�������̲\�����Y��õwx��d܀L��c#70� ����88Cz�z�ڽ��7t��Ep�n3D�.KGa�)b��n�<�4�\�aX�sv���H��GV��7J�����H<��5��\��z%K�@V��[.R���bn�Ã\���^Rx��H9t��*JǞň�ጌ�|XQ��h�#���2D�gԶ����Ytѣ�ثFMZK�ڠ��H%|�@1S����┅Yf�;�N`��<���35����d,w{��I"A�ĸF`�된���:PKA��S%�z�)�ܸ���l2��9#�NƮ>��29ǐj��7�C��ܲ�!/�b�ؼ@�['Y�2`��6	��6c�p
��H�8<���0�,K�"d�sigƈ�Vk�&֯�1wj�H��Р��x�K�d&�R4%UՖ���2�JN\�ma�qU�2VI(
�3Rz�Y���N�Fc��n8S3�*��ѶK��~T`�V�dv�� ܋�]G>�R�Ƒ���~(,�)+�&n�ĵ���[�1��k3�g�鷆�"�=��nx�/f�XҶB��4����]����m8Hw�d]7xʍXd��H�l�۳��J^-A�ͅ�\\��;��7j��ݥXY�g��E�#�:�-�vp��`R4Vk�I%�-�j�ݨ�7�0�+j�I�v򙳺E�P<�M�P���`�ww9�}�L�s��4\N���t/*D2E�1�ƶPt��pRgg�:�ŷYx^��	k㊤6u��h���&6h�L�V���p��M'DX� I��k�3�dwa<)��z9F}����m%Z!�aة�X�|�cDM�e9kR�8wM��zi�'���PA�XQY�=�W$�@5#���ݥGa*��w����[E]�O3��*b�m՜���A�.���t�$v�f���],;M�Z��L�[�G��e�P������+GW��uެ�ޛ��Xh�m�3W�+��r3�X�z�[;H7I[�C��ǣ7
d,�ݥiͼ�D��V�))�5�e��U[���2Š�u�j�ŕf�y`�JH�YZh�Zqgh�̜�U���t�Ad��7��ҍ������$�`V�!�0hM�7�t��Q�P�f�E�m�{�nd5�y�#���8�L'B��"��"F��cx=!���g�k+��5{���J/[��Sa=0�TC5l���L
�s+�J��4BK���*�CU��Ѧ%Y��otJ5ψ6n���XVElp���w��/Fk��sn��vH��!��4s)bU� ��7R7!R��SUq(���,�7e#�#oo5�Y2����$!��U��X��2�գB�@]�%%BfSF��j<.�����Z/%�Oh�`�,k����J
\��T&Gs�#q��J����m��N��C�j���4zjʵ��7bF�f,m�i�An`��"�W\�[L�2ʴ`X/r`�0C8�&ͳ�(f��4����ŔD�X	��1�(��U�8mJN�J(A�R� 	�/k@:��d���+T�]�a������y����@�')�ode�!��L�q�m嵋�.�iêɹ��*�.�e�zA����Ƥ|�ؙ�%��i�����)A��)3�s58]A�\���ܻ�0n��	gjP0Nj�^4E����nZsn����`��񁉗�"�5,4������ phU�@�m�d��OB�N�-���@����ږ�m�NE!Ȟ^}�A*�kP{Z� �;V���Dd�������Q�t�RVA�,�N�'�.�c�v�סe�r
�v-�tհ&�]�<��&i��:�ֲ�4\��',��!�(��]c�@�Ы6�6E[�%�NІ]`�0��X���Y5DdV�m�اGu�73�C��0:��3)1�C� *D�x�׆d� �V�ҫ3M����1<�҉0����{���I��iux�	�)Eݻ�r�7Z�K�j��hɴ����Yl�[�:VEl�w)��5����o/m,�)���r�ښɤu>�t�aI�.����5���Q��̐�������\۰~�6TKC(�{ab��GE�+
7�U��rNiGM� &81S�.���*Q���H�Rfe=6���S�\gq����F�l1�@Npp�Ax%z�#�]�x�0�r,Fi��;)��cLO$����&�j��0I��-ݍ�V4l�˕�bV�LoS�M^aϝ�0Xn���il�W��Y2��XO��#6�Ѹl=��A��nn4X��D2�.伽Xn��+3D)�u;�� (A�G.��z��}�@*����5��z&ռ���d;��E��3V,�B���ƶc�>�mm ݽ�њm
�3>y
�F�Vc5�XWZ��
g�Br��%Ö�T��/D��u�Cs�P������N�pSZ�h\kn
���V��̑�����D��N7���;eD�v�-E�.�PՑ��cqSB��\��ik�J0��>���W�L?ޟȲ�%ĕ|����Y�ئ���a��k7sq�����3L'����Z)��$��S!@�f-�)ּu���5
c(��ܰD�X�:�ƊŸ�v�,P=�C!r�[T�Ǫ�H�)[���TiҸn��%�!����G���<�I��LQ;6 ~�J~�V!�L�(U�Me�����bd�ѷF#	r��d"�׵1�s�f�V�E��l�������Yje7Db��:��A�8���6n�؆�7��$�MCA	��&Qݭ�/&<�f�� J�13ZL�2��7�en��h7tdN@��j��CrʸV6���n�
Y2�F���47rn�yj�. ��.-F�x,�m�L|�2k�^�8��6�'9R�p�;�X�H�����[�q�pѹ��*�����9���#����H.�	q�6:��bj���x�Wr���]:妧zG-.��B+;�v�]�hgu�m�����!V����g>�
<�#�Ţ�՛�2��lF�uk�Ξ�� ��:mQ}`4�;ҹ7��L�w�k-�W����ġ�3��'�B�*z�5�P�� h;��ԛ��
��곧V4�2e�{r�OR/Z���P��n%&��h ��	�cz8��-�%�-n�a�ʂ�*SVĂ���ː�յ܅T���a8�&��A���ᴯ�3s�v���[x�ą3Tb�TUk6�8����t�ڦ�0�L��Z�m:�d��mD��L��⊙
�����;�Hc�Q	C���,�\&�ν�O9��FE�@�p�R�PS��7 L\&����j���v�ڼ�d� X�\ۃcOB�FJ�lE�[�n��yfx��K4�)����>�2�o���-�q�n����0/x#�����/v��X�J���t�SA�\�EX�f�-��]a�*��t���X�5��pЃ4],�d�Tbk3]��1������6�2����zܙ	��6�VJ]�b��u�B�aN��V� �b��M����gj��WL:U�ı�G	�eԼŉ�FE�B��2���N�Z/�G���:��7S3�������1��AO^�SjU�V�ȍ&�#2�)�{(:��R��n�w4U��YF�Cf�<6!���v�fMq��z��]4H؃��nb`f",6\c�t��ĩ˲��(b��r���{f]�6C�Mc�p�ј��[L`�1&e�͓0�ʼ�eP]�F�-��5	.^,�8PB�.DrZ���wx��3�.d\�ҕ\OM9Ve�ؘ;��6sEり؈�3L��
�b̀�-�:���W��џR/A7��1�[3H��7�����M��:t-���6v��:����A�+ulXV7���n��Q���Xʰ�Y�b{ d�1��II�=����K����&K��?�+k�܌޷�̘�zM�E�jD2���;޵�҉,z��S���)
���dӴLH�wm�fXvP܁ۆ[�l&i+ܥADi�8e�t��J�ܲ�Bh�d�2+N���6��+0�.�Rr������ma�p�+l<�
�����4��:O6r��s�1���M�ci*јm^����Gt`M��o�0��a7vL
1WY�G(a�h݋���X�p��/!�z�j�0m�{��Ȯhf��X�Q[4l�r�\T�������ӣ��Rl�wV�!��۠����9vv��@Ĭ0d��nW�D)�OK�d�R�q�Z�+���˰_��BavX�̺D#p���$!vF{�����,e)t7w��e�)t'^�+V�+$�+�Z+wU�K�Xv��H�Aբ�)���1�nٻïsh)%ej@���l�1h��Cj�6�ֱٰ�⵹c $���lY`���dx,Y�`ٹ�#��J���ʅE]��r��{[`)�8c�bS%0%'y��n�Z�G��A�%q �w%&�]s��I��Y���BA���$�����˘
:њq�5�h��{kQ�&^���LM��t�T� �G8w]�+"�ʹÌ���2ȃh�+08!�uw��>2���$I[�p<SZI�#pK��Z��3X{)7��n�B6()��:�̬�#1$�:6@�&��Kǖm�4Him�CZ�ȧ���� n�ע2�٣Dն"�FQo&mL��a�jA����L���:�H�e�Ɗ�W���*�6�b��뷭�Y(���*�R����@⭡�J�ûE�B)��3��#%���;{PЧf��+$�f:��X��Z`�##eK�Y��;��2\��T��1R�V)R��Lb�e� ��v���{�A�y����F�E�n�|�?X2�r��9�����(�;�84�P��k�	�hV��Z�`N�&�$]��/!ueh�5�C �Z�a����VB��*�#$�r��3&�B�SW%�� �4!��;N�,���;��R͑LhW��m!9o�%��# `5�k�ܳ��#��*\�,�(+��(%=5F8m����u ������\���F�kxk0�z�l6������hP��������^�F ����l6�n7p�N�@��=�� ���BL��E��s��(PͬZ��ʷ�x�����/f������]9ꊀ�ebF�3�ٖ
xcYm�b��㼫���xRQ��R��
H9hI�4f^���L��0�<��L!e��=����i�
��!�ҷ+3�d�T���4��7��p@�ĉʗpH�t^���pmdO^��gE�(1+��)����仨;2�o�o;���h�oX��ē�*��ͼ�%
�䆎Q�w�L��5Y��5�� K�;b�5 �A9���ϓ���&��eB�hy4ݣ%Y�T��r�^�H9#�=�*�FD���wMLᬩ��9VV�����kB���N����,*i��m���	`akN�Ǻ޷�&�r]�rJ�|ísa$���6��`-�����y���+b�1G whG:w	ttS5�ީ�@c��
Ŏ���i�m�ä��Y�|8EgN麌kXO0<Z��Hq!��9�+�N�*͊n�(��-���eia��ڷz5�֌`�Mt/,T��c4�j�+e3�E�C@;��7n�K?YntҴ���A�����;
��A��F����S�tD�lb-])���[DB�60�ђdƱ֨���m �@�r���OV�BQ��z�Z/RZS�4e��o(Sr���������Y�o�P�  Ʀ�*D�m��թ��&�e�1mʐp%2r��mkųt�'#���Bf�q:����M���Sn�<�c,v`�[��oj�{��Ю���"�����&V8�+�΁^�hKܰT`[�L���B� �����cKǧ,;&�h�������)[���
;��Rh0́i���Q*�!�h�t�LuZ Bv 2��N�)i����F�=�	�RY��=m��O~3��[�1�p���u*��]�Y[�8�Aj�ճ����b�1��U
VWP`��ն�v�N��0[ `�n�%��l�l��Z����l���*�*���3�z�4��#�ή�ea87-�c�4tj�����W.N���䃕u1�j���V��s����ۑx�%* �8ɳ)����l����'t=��3����t'7[��l;^55�%��:�<J-xK��Qla���ś#q�����,ZE���ą9�m���x�^6�coZfr�Ӗ^]��\l�6�vQ�h�K/=���K����p�s��;�.И�\�;���.}<;L����6�y���I��|�/Z�����8�[G(�<ذv;-s��6�&�a�"����<�<l���W*�t��"#<G;�(f5�[e\ET��XS�n���5�Լ�k�=p�jGJ�Ù��+�kt�3	�x���vq�� ��ǭ$� V�\�W�)r&e��`�4��Rfgɞe{���g���n�u�
�������5om6�Z�4LYc�n��d���� .��
�{Ml�Ռ�tPB�au�;{b<s�+��,&4��zW�͸���B�3Ӧݫ=������J�W�nq�v���;Q�d�/�sjI�e�.��8��@. ��vr�Ȩ����t{ۏnz�k]{JZ5�^2�}����2�lݠ�����U�[	�"���F�6����k�Z`n�SY�����9^ju�^<��|=�EV���i��n����.�K�p��y���[-�)�n3W�*�+���(2 M�݉�YZŔn��e���K;��ېz9�mj2u�Ӑx{MK�B�d�y�q�Byf���v��s��>|o����5�7��X�X�I�W��ֶ���3zBv�ݦ�{iCQ$󘆛ҺVh�t�-�1ր;a�unz��=*��qβ[Yg�7U]�������v�M�U��;h<����f��M�N #�s�e�7X� ]�q�)��4oD�F��p.��u�ya#��G]@qƎM��á}l$������%��s�rr[8�&��5]�LQ�ٷad�Z�`ڞImd��:7G3��.k��T�[���e�!��1�a/2,l�I`��M|�:���A�A%�; ��+z�.5]-"�p��Uw�Fƍ���j�l�W�	m	�s��=v�9�n�#����Ez�qd]������͞ڗs��+�S����g���<$��:5�@�9�G%���&�u�C���K/H8�3gm�۝;�u�M�ytmf8��˴)yN�f�l���s٘����۱�T3(��"�vk!q��$0x�p[p�υW���m3�'�ḣ���cL�5z�HD�m2�FY���uvrׁ���J@��`��n��n���]	ق�lc81c��5�"�4q���.�;;t�'C����r��WY�Ks��}ӱ��vɩ�±��Ռ*��R�ۥu�)���<�Ll�Z]��lv�nn:��tY�r��
��frVٵ#��,��<s[<n�	7)��/mbحɉb�jkh�te,%Ь�&�-WTOj�x�$�J㬝�f��2��'F6��=�u0d mt�Bq�:�4�:�y�j�3���
�n+�,�6��
�J@��:��*�t.�f�T��.f	y�&'���7\���۞��]=Oesn�c���L�/..�/x���q\p�M����:3��ֻmr�;���g�jӝ��\qJ��ѐb}��s9v&�l`Ŧ�J�D�$�M`ѥc�Ɗ�P��pCcjj�>y�K�<� :ˮ���D[��{rK+n�v.��W>�r{`�G�C��ZH]�����'o5�ǋ���̅o;��u<Ʋ㮞�G�H�X$�^]dn!t��	��^� -c/1�o�+�VZ�u�����jԆ����QzIsmSaY�ʻI���{�osC�4��@gی�� �z3<Q���Nv���_,s�YVO[�>�m�v�]��H��V
�u�pnk��ۛr�>C�HnbVU�kdŖ,�,ж�����=�rv,���/os�xq�jQur��v;n�ky����b	��ʙq��B�v9�>1��Ƴr�[�*ygy��� %qbNƶ�	�6�e�p�;:�왭z����p!�';;�:@��(��s��N��;���W,�9\*S(��8�.Vb�ݭ\�cvL�)E�[ծxp��9�9x��@���i�{^��T^�����n#��8��
���G�-6��3�l����3U�E�9�O�h&f�m��g�6o��S���+��N��@k�ێؕ��{�!67<(�1����v�d�r���v�v
�����gm'`S�5<n�L���n�̞�;Ko�(��s<"�f���#��)�F������b��e ��Vh:u��c�ɳeh���c��qn��Ac��\�V��q`h0�̪d� �Rb�3+���`���V}��)�t+U�Z��v.{��!tۦ��]mvr��]�19�j
�	��g1X�ٰ�fv�V�4�Xg��Z�-s�	�!7k�,�+���n�kt��z��&27��78�q�=-����x�N�F�u�0R��$�c��Fj�Vb^���F�h�����>�1{=c��q4ġk��y���K㼳\���d��u5��\ܷ\f�E��+�P����Q��-v�I1��ǫG��� 5��Żv���=7��I�'^n�ݎIz1z�[�Z�4R��v��n2�4qkG����54⽈Vf��Tj%��y`0{W��X�ѷi����1��˷1��r�r�-��û:�#�N��;<�����4�\kn������z�Y��y)���b�a�+(%c�ە!wi�R.�Ϡ�z�ƻN<v乺nG<�4��J�m���ε��%���:������7o��Zm�Շ���q�y;p�+PjG\vS��s�6�bk5�c)e�o;�
�X�{=�}x����ȶ�5�Q]�����l��"U%���x�)"��Vx&s]�Ց�Lhb긂����u��]iL�mѶƼ�78ơ��g�s��t�<���#��k;���nqVɸѐMVq��="�^^��=�s؞�W�:sv�c��=���@]��z�)�ݎ]�oLV�sݬ�"m���[��Р��倾٠ͣ:|&1�y|u;x�s��n�w���]7*�9/X�w=��cײ<X���c<��ܶ�kX��"�P��nA�q5��0#�p�4f5��;�/&�9Iы��5�2>1+¶�I�WZ
w�#4�g�5�`h��s�c��x����n���ti�Mm��Sp��OPDW[��O�a�x�㦔����B]�묃c����x�(�JW7f���yv㭢�;��1K4vF:���!k`#,�/v��8#��a�� N�l��H�3yyK^Hp�/<A�E�u�w%�Ӯ4�qm�y{��Ղm���۲�Av�d��Cns�5��(��4��Tp�Η$�*�]�{Tg�ޤ�+q\[�µst��m��#�f�m���ϭ�k�V\�v���N����(v��.CoO�m.3����y���멸�u�ӎ��H����I���js��L�=@�\E؛nR[-�a�144R�>�]%aFzg�_=�x:� gt%�ϰ������"����j�ݯn�:�zx��s�g]3��p,�n�Z���1m�q��i͒ԭs��}g�!�ᚳ�;0s)j�{�^����h��<� m�Wc�x�`����6��Crs��� zŸ=�v�e�xN�n��T�����#խ�s29�5�(�8%9��f�
al��.�Ʀs��
��h2�e�%(�����$�B��p1�v�GU�SG	�W����Y8��'�q��g������:�����m�.s�F#M�'h����xO7]\�=�f��6x�u�T���/������dh]	c)rH:ݠ:�>m���ۮo\�6횞�ѫzx{O��w]��Z���v3��s��x��n�蘗J���i��1i�:$�FO7g�m�n�]x1v�&�OLl�E7/1�1����ZB�eq0�J�T27r�p�N����;q��r�f��W/;�'Kr�ӏgO;yz��AvN;�K��^ք��L�Qm�o\��\M�G�s�l��t`:B�X�:�i��1퉔��l�](0����H�l"�L��]��I�U�#�JE@IX�[u�itGML)�-"-�=y�t;i��ȗ���Єta�kr�X(�$�YA��P�<a��^ko.n{q�+3<���_n��#��l�m�[{jꨂ�9ٞ:�Lu����������]�Y�����X8(8Σ��=0�i�B�ٮ[n[���'�xlt�{w	nx�`5xݜT+X�ZJ��5��YhM^T���c�Ν���n{V�<��<Kc����5���Z�A��f��i���=��#u�nLW����>��\Ts�g��| V���k�,6���m�sA]�V���9g
�z� �UY�Q�7+������i[����s��.���c��hi$���
�-v̜��k�xjlAO<��ɞumĮ�<܇��9��k����`�$������1�v{Y���[�u���˳\���b�Z�qۋ��8�g+���%�j�{Z��X���c7[f(�*'WF�
u��ɳ�DvU4\���̎��6SX&�:u�=f}q���d���%��m�5K��(���@`{3q��$��V[ڀvݛz�Gm���Lp�9Ͷ��.]<)��pa����;8�>܅���ۛ�n|v|F��s֗��Lt��	"	R�*��Ew��x�>Y����YL,t�������0���R�mm6:�vEe
R���ƧQ�a7&x�p5t�myC��VZ�FҲ�ض[4n�`�4t��}|��l�iKgu��M�Ղ�t��d��(�.A#)R4<�	ᦌf�|S��읲���v�u���V��
7O�����8c��	�DJ��
��TU�
uU@UU_��UP��R*���(&�ZUl��J�V��q\�nݜ��<��́�1vqnx�oDp��n�1�oV��q�)��w��`�B^)�'��l��=�1�u�Z'^�5��c��+��uη��k�]���2֬��I�b�,��Rx�<��Z�7�W��p8���.�䆗2XwVw�ɓF�s�Y�Ӌ$�5�κq�&2�0�\`Q���v�fg68u�n�����r����ha�&�8��{!jz\��r��-�ld ;�\�Y�۶]�x .ǯv���]�5�d,�{5��x�װ';1gO����E#nnNͱaHQ�Uఆ8�ϲ5�Nc�l6������wA��h7F�q�����	��m���"��"�N�8؊��[��^�(����s�Mh����;yk˙l<�CU�C�Wjkҵ��8�RŧWj�7k�q�{
�0/��R�z�ø�q�<�m.TƂde�`���u�T�1�`N�Y�1�C�m�zlT&��66\�̛����y�`��+�n�1�z�^�Y7f��:K/hJ�۶M0�v�Ųm�m�msّa�N˞:z{b8���9��k÷��ϴ��1������A�y�x�&bu����HNYN�N���z8m��vTcZ�&�\��``������0�Uv[���Ѯq�4s-��x�k�;�o]t�2�gl����S%�taaë`q(u�0�,��b��̽U۵�sqۛ3�Ov����-vۛ�����*P�p���u>�\C`��z�p�=�z]]�m�$5@�Ծ{e��!+�df΄Z%jm ��A�&ZL혘�ee6�7©���pϰ3������ZŌ�kD]��e�fn�2��ep�g��ε�4���@��F���aS`x�f��>���/[��8\L���
�k�(��\s�=��Ƌv9�uz��rq�:����Va����<k=���3)���fB��Y�^y��Jwl>�Fm����ͽ�z�S̲�.�`�܊��@P�� &� 
�	�UUDСT5D�� M
�$P�P���H'@�'Kӻ>z�7s1=u�c�;v7\�����\�*R�)�Sh��9�&�������2hE�F	��4�WYJA��%���4۞�x�9M4��i���<vܛ-s6�.`�*�۷&8ۍe�..�S�a����\wlrv܇0���y�f�sb��ؠ��K.mܚ�ʺ���s�n�)Rtp��\nE�f�^�7l�[�iI�G�i�;��{U�v9��#j��ڵ`�R��m+RX(���e�k[bԵ��?��x�i��#�˂<����#R��Ƽ����M�}��L�$����dm�6�����("�%0���!�x��R�Us�s�9�@��� �V�Q�[�R�"���
�w�u�AMÔ�s�s��c�h�r�jSR��� \�Or֜P�#��奪��n䵏�3c��{Oh��vv�>� Io�(�@��-����z�z�j�k�h��h�vl��{�����=�5��8�d�n<A-�
�x�ӡ�A��F���s���lp_"s�h��v]�Mo_8�Ec!�����>����o8��X� �K	�	p��V�<z�v�٦����(�γK�L/a�����Pb�.�!��t��t���;�dy �+��X��ެp}35��T�9�r+{rx]g��E�!p�.jg2ͨ�'Vq�rF�r�2A�a�5��`ڰ��s�=ՉYe�����v��E<�ې����̬� ��e,��X��l9eMn���M��e�8,�Uh�<��?�M�C
,��!�.��\�/o˻�|���\M�z�@&���IU��t�C�?T�~ ًpҢl^`h!�8䷜�>���īw�㱤n���\�z�⺽xX��w�4�v�{ �4R��[<-ُ㦭��ǋ,��0�L���6	zû�U�v)^٨���U��*�(�'><ѯA�%x:
̙C<���(P��6؜�%��n�V�W &�� �I��p9�TI������;8R	eħgK��� �Ve��gاq�R]MB�מ^V��W�l���8ɣ\����nc{f��B�!�m�t����nw���;�ǭq���\�,���Σ�����,�Y��[���ݺ��.�����eFn��4�%v��^�J_�Õ<��wrһivHk�6h�5�͌�h�L6N���e���ofsY��e>�n�#N�d�R,��H�VNMҤ�����Z+��'�� v^!��r�)׶R�7v�'U�@ESD�7��
�V��i{,�4�-z%wt�~~,;�k����g�Zbc�p������Gzƭ�����xgu������|�A�X��h�\F����i��Ǻ���3���gt��:X��Q��O5=���Dtlַ�6�ho.Uھ2a
CE%I�m`�9��������+��+lڳ����1ݤ%w�C����[��)�ל8æ�[�L�uw���$�,�m�S����0Ӽ#�j�Dv�}$y.�m��9��B�ڒl���˳]�bXk.���}���k�5�#�x'�J$�r�,͝(�����j�hX넯!mv�{6��mu�䷞�QɴҬ	�Cv���y燒y�ͳ=�T��!�)H���-�̊�]��t�<�>���l�V��%�]�:�Ok�J&�f�x��"�qdt�e��f۾ٔ6�L�ױ�.)[m�"=�F���jA/-�k�U��(��Y�Y���<r�[b�:j}�&,�so�򡆷y������n)$E �-�����uߺ�t�$�b>�tn�zH���MLGk>^�4�^���t�'�
P����!f�F�:��?-�:?Y5f��4�L��u!"��G5E����WQ��$9P��~�&�E�}t����ď�r_ۯM�le��8-�^0�;Iv.�e���lXsG�TV��4)�^�kh�P]�G�S���A��(���D0���X%��n��In_pE� ԑ��H[�-�i�a��aSwZ+m�+wţǧ��@t�I���7f��C�(	VX�\k�n��
'�f��ӂ�*�������~
��9��GMb��'���v9Z�k`IZ;b�EWR:ֻnp�h���;'��C%(9(�T}�ޔ��b�Ɲߩ�DCG�e�t���݃ioކ���}ޅ����j���9˖G��� ���J�M�s;ϽR���ש�|a�>�f�b�f�@�	b~׮A��Hj�E���G(��)ϼ��}���6�������}��V�X��mu�`�&�dn�}����e��/�&Kn>H�w������5!����@�Y�B�dô�FJz걣�[�g���y8*�ͼ��[�<�� ��[ս)xWwe.}���k�2�S6��;]Y�U�W��Ȅ�����8 �(ړ	{�RO���Vi��_���(��(aS|78T{=R�V�zz�+U�ҙu����QBïй�,�')R���#��]��L�k���p���
]�V&CE�Ⱦ�ܾ�ӹM�M�i�\��+w��4�ʽ����X��rk�Ͼ��&���OV ����b4ƶ9t�����f�ѥ�Z��^���bxp���lBݸ��r��C���x�ru��nv�7�͎��,h���V�R��JѷJ-�4���+�IGi}�\�Wv��@�F�q1B�F�Śd���a��X�:!���z�l���<tq�=�`P�q�H�Nh�OD�ݸ3ggn�<�s̎5�[-vwf���]q{t����]�\0��f��s�k��L���=�\�y�n޶q�t&�gA��!I�SpG�.Y���Ͼ_pw�=�^̖Jj
Ḧ	<����4g��seK𮘳Ƥ4�X�UX�7o �91Wf#�hLq��p��
H2��I�N�?V]<�U`� �����5e6F8k�6���߻��F��J7���1���Y{�:n��u�2�q�\�r(T��(4٠BN�Y |e�l���k�.��to���O)-���ͪ/������^x��(��|�[�i�D[^Τ����L`��-ɕ������Z�z�J��a�?[�
�~Cn�nO)�k��u�P�V
�c7ٴ�-�*���AU�S�{p�Y��_�Y�F����0[I5	N*͎�4��{Ʉ�C��>W�~y(V�=`�,��W��1�޻���}��0�y�w�/�EF�@��I��lD�x�U�^v�M�a7kw9�e],�#b�kFZ鰎�҄�,2���m�W�V�p'�YP�EypN��_9^��Ƈ����n�j�g���h���Q�lxE��%����k����6h�#����!�6e�cW��;�Y��]];$����Y98ky�iў�ffQ�F�)B�Yhmާ�Qf����k]�*4r�n�h1�]�t�Fb)����u�N�m�\�� �gz�×Y�)
�[+W]�4�MS��n�T�=��v�N�U��ǵj��X�0 �Ԭ��i*C�S�y��F�=~��a�{�f��"� R ��U<i
^�q"J�+�j��s�`X(B#�/;4��K���vX�T0�]H��Vl���L=Y�斓eGv�������eFI��n$�Y�f��@�۸om�&����3����]��m潰����#�ͣ�Q���o[��
�,���{�߳����,#N��q�%��5�h�E��v�]zo$W9���{[[�.1��F�]Ab���'cKy��f�Ȅ3�j�I�Ӵ!��	�x�s��Vq��fn}�zjFv�G�~��5����B.�L����Li��-Y�zJ��{�!��2�9*AŐ9��]�!\�\Rʄ-ܔ�A\�,������0�'�ax�*�1YlT�|��,���۽	����{<%;՛�ϯԽ�)���uW�loc�}�VQ߀�������æ�����&�Z��T��5ڍ�u7���F�d�0���S�#����VX6*y��F��i����48��[y; �0��~�7O{�/"`��L�Np�D+�8]�"lͲ
�Rꂵ��k/Q$]Q���+��:)�m��	p���|������Z#N���!�D��B��d�hA���z`F�s}ݰ�yqV,-�s]�H�����|��f�B!����W�x7��a<���m��ѐy`zn6�!DZQ�L�W<�pX!��CY|�^�GH�=�<��	�/Iv�Μ1��]}��X�e>f�6�g�'Qe�98���"��C�n!�H�N�Z�(�+h�O֜�\���ZT{�N8�h���ܐY䇙k�#��p:����_pB�To�rR�����Z��E����xP��#���sx!����f2l&@ϲ�]/	~��!�
NN`���K�bq{��hV��(gfҫ�*u�C	�Ӵ�1!�n�]>����@�4(�{��=��;û�p���D*�#e%n��M�����WA��+���ܱ��� ��wZܦ�1m����f�SE�������f_Z�mlY�ܬ>��a��WX4�uţ��]Ѧ��Xu���I[�iѸ�m95�m�9�KAB�H��հ@���e�cM�v�͸4� >w$ a�X�*�ܲ���/Yx�V#�5��vu�,�K �}�0��؀�g>�z7s�yM��C�x�� �i�$en>!�7=Z��\�νv�;]����<��|]I������m������T�����ԅ�*��Gإ�6�M�纮��:մ��V`�^��:�*����>���nGu5�z��,IO����ov �Ђ3��U��G�2�9hQ�I�n��ۥGVO��B���0b5��Ie�GV����U�dI�B)6[s�>���Q����EQkv��m�%����D�1��xHk޾ʅX+b؎���C���`����
�"\���*}��/ۄ5�ױ�T#H�Uf�S��l����{>��!��f��
��¬iy �5�$>�̷*�hL|�I���$ft��E���Ǳ�ry3�9�U���XR0 �*q+X4n�:��=�G�����識y���wuP�n<��c�&AY���^ZՍ��~�8#qul�J��>�M��s���cQ�wGgN�\���}�f<(���=Iǯ��\U5�r+�ԟ���T�.�%9a/�k�oԫ�Ϟ�[�t�0�(P�Nth4�a����[Q�ˍ>�2�l�����*`�ق�kgqb�s�8����5��x���b�Z����E�Y�&X��v�Ğ62�`�$�H����v�'�����Km!,��v�m*�fk1���s�w<�d�l�b��١l����5�����/=.��P���N۷dOgA�����;��N�J&I1�:s�c���E�ۘ�E ��ݐC�2=��^���#�9R�}uw�ua ix�����޴�5�"Ɂv*�K��X�W�+],-�ണ ���ԄեH�GK\�e����Y�GBy@�j�d�'^����&�V�������ζ�;/�r,��9Y���f�c}gP�I�q�"I&P�h�ɩ�5�}��{���p��U�q��O2��WT[ �&2XHW2C���w\+Y������)�""�I�c���9j�������q^]0)wV�K�ˣ�kn��P�Ԙ��RPx9ouϼ�ab����9/O�_9=�}I[�A��o)�D3���k�����}a��OVG-CP-�xE��޿{ϻ������������2,2�T��h���-
g!�{&��죚�>�@��)��)0�rOg�.Y8�ޠ�B�%��.v3�B5�G.na��ˤ����_4�f�ғ�ɯT�&��Cx��j;뚯��Xz�f�s���y֚	k7[��ɯ����#�بE��=���p5FF�%�/MS �e��Y��vU/l1�Ĩ���E`�R�4:��I��*k;(
��^֬X�л�b��GL��膶,&��5����v�5�ht�7����F�c�}��1X�(���ͿPwV=+<�&�^�?"K��t�������$��Y�Jj��nŁ��4&w���F\�wƔ��b_m���u����� �X���<�&��J�}�!&�	�Y8�L��H04o�	��W���+pwr�2����4-���w�`HF��9���y�P3�xYY�-��_\�r�T�U�c-u$]Jr�i�@�6?Z�{ɦ�wE+����X�����oԼ���B�[���Оi���L��LR��B��8-UF�vazI�os�wX,f�Pz��Sh���O�z͎<3�{%u��.��X۶���<�7��/:뛱����;|���O�Y��k��
����uJ8i�.18P��	�Ic��K���9h	��K�p�/����$10�ʑ�Ø�3���o�?b���ĨE�f:l��8B���>]� Ulw�Y�cN�yn�߃o�u�$�n�̳( $��V����@,oo}�L@��. ӑ����An���TAڛ�챦�߫ 7g��rA���9�|-0IT�SfG��z�@�E�奓P
	^�ܵق+&bo�\��yq�+��oX\��5,�r2���ɃOf�Ais2��ZCqˣ�+�I��6gUe���.S>D�� s!��Xʡ��FYU�|N��Q�B�p����3.�'3^��*�=Z�G��n,��!VXt�l[n
mh��˧/�V�[����%�jܧk^dsz�����:��Wn*}�;�9y�8�@��Y�D!]�X�V͙+*�j���"491Z�/T�����B�Z�Һvö(�!3*�������#����X��܌<�-_�,X�#ɜh��R������x�mc?9��VAde��������õ�R&�}�x90�Ue�1Pro/�WM�`�փ�AηZ��J�xi���{�8Nd�(�&�bQ�S:Ӧ��	�>׆Z�Bɢ�Ӱ,�nd�ă��n���7
Z=k�.��zӨ*�3��T����<"Dn�f��VoW��63ܐ��}.eiqK���J���}.�l8,��z(*��A'Y�[�۸-�Z����Qn�sUk�u5�ݓ�D��l�v�a����"ie=�=�uC��˛�ٽ�j�;�s8=+�%j���cvU�;��(��gb���k6��u��bu���oG���Ё����� ��v���Ѱ����S�/pK�n�O�kX����8Aל{%:CWA|�j�f�!!<;��o�Z�*~�s(����_����J���� t��Y����C��3|�磭ΙD+���g�����5��b�t��^��n?@�{�|6�vW
����Lg@r*h�}��i�13e�	7�w
ԋ� �y��A4���qa�C/!�}L?0�Cj��{?zq���?�c�%$����ŬQ��M�E�5L2��{nJ4*�Q����J����X�{���� 4�,�#o�َgnz�Vh,Ƅ<���Eגc;���X6�WY@�6�M�&6�,�۱��+L��Kn���@��3[������̀]�=���A���z�7�=�F�ʕX���(�a�e_��3f�:c�f2����n�aBNM��������a[�-*�L5�l3��4W�"�W2���MՎ}�7�>���@�hUL�&��D��II(����C�����Mk�J���O� ˌ�6��ې�/84�f��<�/��h6��b�=42��=���Plu P��m�}��*�y/����`|W��F��BER5ߵJ���{�
��ﰉf Y�]�W�Y#G�/y�3(�p=6cs\Q4+Jײ�[ݜ`�R��-��,h���h�X�a�Yn,�U��M�$C1�w+"9��>�U���R��>��n�WT���W��̟��Ԏ�|停�,��!B����D��~��Ɏ���9���A�t�M7��F�K\�s����,&Pf�;�Z5n��w:Of�]�&=J-��i��b��;o+��4l�r�nB�˘3[Lo�ﯿ��*����D"����Wk������>Xj�P���塧��<�.,�j���/s��U�aׄ^�{c9��G-�R�Da���	��}�}W���\��i�X*��:�31Fj��B���Z�a�m�E�A�S���VE�`��{	X�.�$���IS�qE ݯ`�0��l8���@cT�"�����Y�t>P�*>���o��o�"�*������N�b�{4M��
���|��L~e'q��B��i� �[�-�[K����G3�P�ag"3{ ��.��p�t �M*m�b.�2��Y�g�������K.é�ۢ�f�a7E#R `��Ӛ+���u9|��ީ�FK�,���5��n�Q�TY�;'=ֽ"�� ���ܝ�.������ˁ�t�Y���;/�'c����
�g�pr�\v&Aв�lGu(E$)��#r���t�:�fU����i��n]�D� �W��X�<FL&�luJ���sIc�:��	�O+�ݪ�(&�f��4��i�aI��Vn��e�mv�Uz��M�Fε��us���������T�Z.���wF���^�y��n��y�YH�g%�����vy�ٍcI����ټ1�8����G�z2=x9n{\
�������s�`��z{��9-��.�� �h:w;.	�]�mQ�θB}��%��S�δu&��
n_/�{O;b��:�Ӏݸ���[���6;���8 e�{�0o��1e��?_d	����l��v]/0���
Z�Dѹ��zCR���t�4"�("(ԃ�D"�uȕ_q,��P�f��xl�U0n���3)k�7J��X�~��zy����TQ>
��ԣ�1��i�8�d�����nH�l<�gWs�W�q ��ё��j�	{��`B��f����]x�\4�Z�W���K�����%�Ai�-����=�f%�Ͱ�:w���Dd�i����"�!Z�C�>�,��f}����Sȟ�/���z~����SKk�d����l���Ni�T�fV\&�[��>��4�d��T�zJՍ�r�<��e ��ȸ���,����D��Y��-��M2� �hź���j��O^U���Ǎ��y����["��;OC��y۴S�&�nk2���~�u�;���,���E�A�vy���̉��>F:��0N�75tެ����n4Hi{a�V�e��� *6S6����¡�꽺�|߂�>G�7�����i�n�i}"+ ��F��wg*[��֩�`�{���euL��p��v���9��#YQ�=հԝ1��[G���E\�K����"ңo�U��H|��US�:�eA[���
�����|�\zy���3n��hc1Yl�0�t�d�%_'[���ƪ�D�H�H�DR���ޫ��^��OWM��O/�LW�d�L$P"�9A]/���c��l~�kDl�h�t{�b��V1���@�[I�h�ZJW��#��~�Q�0�h,B�w��.n��:gz.g.;�WJ��8�/� �!��%^l	,)nH�B��e��8{1�*�O����2陷Z9ؗ+���wKuЄBK4�5ĻaU�B;������:��6j�B7W�Os[߿�����>frb$�Tv�a���+6�% ����fD6������Vy�&m����6d������&5i��X�u�t�Oc�]���a�aB��E���&���c]G���d�n1\*�
���b�Ҿ�}�2Z$�(  m׳��[uY���Q��Ү_7h�!����Q�B�0f ��PێοE��'�;_+�rr�����0��}���z��	}���G%�=:ƒ�ln��+��S\�v6+8��k�u��v�q�OEY��DP[��̃٧j��X��{o�Vo͏D{6���lHk��s�Eq[��O�u#\кH}�pC�e��b�Tn7L�/�Tָ;$l��1��j8;��5Fbe3'3�H�q��n�:t�ETǀn֩h�^
�*��<N�*ϱa�=�	�2 �6b��o��CS������������Ǒ(���,��A���(�2�>���vȍ�^c��n��(���T�3�ۗU�N�,W�↸��J��I���[�S��a��tsfvm�,!]qM��e3hm,��L3�B���˱:����
�&2��C~����~���V�7K�*�R�Vt�EM�_3ܵ�qUɡFM��v��,y5���+7)."Z�Y)�M��i�>����	�-�8�
�k�=m�(�#��;��V
GȊl�踛6���m��Q��x�5������%&	Gah1�Y��V0P�z1UxP��8�Q���iͥ��88��QP��Cn�f��"�]�r�>�𱁍�=MM�m�@Oa"�<���#[1�vm
�._M�:Y$q�*1N�L[c�#u�\Z{���`�*����K��]���.㕜pyaRm�|���A�Vr/,�3�1h@l���ct��'^i9�	L��ӫx1���cw;!bc�^�O����X�dq�Kq(�)Ȯ�2)o7��)k��F��z?�DM��Ǚt�	yi.1��+k0���zc��l5;eX�1�-,۾h�]k>v�{�D������o�j�����������1���t;�����{n{���@����l0���E�le!A0N�xW<U��Z<,g���a�B�yMNy� �:�S˹|\=�;��d�OO�����<4��PQ�YC{1��?s��G�N��A [,��l������$>[�@Z�"��F���#�Ȝm���>"I�|� |Y�j�y�#j�G�wN�����y\U�֥4%B�1��m�j�M���|�J����P�9p��6��㧗j�8-�;������`|{t��g�� �~�X7�=��#a��1�K	�vA�2��~����c6h;�80M��
X� �+Z�i(�e��&���vI���M�*c9@p�;����4��s+g���P�.	�b�7�&>�B�ї��$�$J4����a���,�Fڝ��b�DW"h~R;�{�/�Ls��#�B5�Iz,��H���g[6�ݢ5�j�Zcl��>Y��љ�Y��kr�d]`��8��B�T����݅�G�߉��ֱ�-�0�Ʊ���-��%���8��8�d���H��ۤ룘p�z�^wL��n"b���Vm�آ13����k]j-bі1X�ݸn7c	�㪺�i�B'n�A��7�`�.�ޅ�,�.B�nTx��͹�9�U�K�9tH\]�ؚمm�zx�m�Z�i��=��uc��vq/nS���|�+b��Ͱ��Dlf��\7A��MZN7Zn�n����;�g���K�[�45�����{���e�D"ȿ�ج�n�?c?N��Af��<$T���{r��Q	���^5�}�f�ˤ�º��Fi��D0��`��{����nG��ωž�w�s�1!��H� }���4��a3�D1{.���۷�^׊5��Ns}��`i��Im�h���l�踘s�����c�)x�Op�흡�9����k�{� �)*�I�C���h�����X
L��6Ϊ��z��7r��o�Dp��9�"�wn�}!��e��ӄ��pWGJ
���[{�Ү�L���a���eI�����p@CjF�f���>�E����� a�)���v�c���=j=+b�a�U�x��?+���/\�WvP��`rD�FP9b�b�kӎ��٦Ѱ�fK��/d���c�xtcnZ�Jq@�ѹ���z*�s�c��W��ME=�������p�C#�?$V�ktOf�93�,�i��".�����
�E9��(��9����)�ԿTm�I�ۜpe��/u ���b��͹�SOo�hs����[4�)���nS(��{�����',`P������*�m7u���&�ٮ�s5[�]4�_qF��$P{��/�/�Π�>S]LX&0rfK�to��uޡ!�mkf'	�@�RF��Q���.� ^IP��셝�L�6G0a������sc�=��|Y�|���x@�T��ܡ��KLh����ILJ�S��n�+[�>Í��S+g��� L�ϧu���>>��������uj�����W(�j����r �/N��M\�
6�q��uP���Yg}�-ƚۧ��o6Z����䣳OE�==������?e�B1#A��!���?[�0�Q�p����sM�h]1d���]a���C4b�Ղ0�@�pee[j4n
��U�*l��ƘaP�)����iA���7r���v�55�5V[�l�ݗQ>C�n{���6iϚ����2l��}O+��|����8��Dn��¬U�::��2E"�N���� �d��r���B���g�y�.t��:˩	C����_��gm.!rk�s��(�(�(��|u�EF��3����`�T�YQ���E%�ʒ�z��1�zɬ �x�C.Ͷ��F�v�2WI�@�J�AeI+`����:���jy�jW�'�|�kfHjN�^̫�p�˪%�e����w�'-T11�C��tAD�Y��e���> ����nE�{~�F/�ȩݪ�_1[�Y��p��зQt�
�tH�g;>m-8�kjў\{��o�u����s�{�(�֭W]&T��L��������Ve<�*Z���`!�Mt�K����cJ�`�3�lK@�ii�O���,�mA�C�^�1[R�Ix�Mr͡[-��S��V�8�g:��<�QԷ��"�6�,��l�v�>�I���!����>{)���wwv�Lw�1H�����[M�o��¬s?+Q������,�SD�(�I��к�����'��+��<;U\n^�6;�r���=�< �Of�}:r��ڰ�טJ�t��@|5�#��2&�\[��ϯ�:h_lǟ\W���)
��5��1��f�Y�(���S�`��A��(
�я�r�<!�M3qv�s{��aD���f6̱D}�J��k���׭�IVwY�2�:�Z���Ϲ[ʙ�#Hh|B���P�C�A�	�ˑ��î���y�5�gU�
��@͂V�*�Ҋ)r��o/X
�4T�p�Y��CJ�	�LҸ]��,0�|V�JP�s��(Կ
j�`n���Վy�+�u��
l��b%#\���G����W�4 �
[a��_xw�2���L4��~�mgu�c�ȀD�i�v3]���)멡T;׃1 ,
T�!�t����n�7rv�H��ؓ�e+��`���m6�S��9"Q�䇵�\�w�O{
{/��kӮ�תU���T���j&����^;b��I�!�b<s��N��j�y%w���Zjet)q���g��=�LtF��������ς3�{�CT����l||���T�4����R���>�L�mm�`�V4꛼l����0j$�D��i:�ǳ��۫ny����iUw���w�t馊��Uq٘}�H��ʆ�
�����B��ʠ��e��!V\Y�L��[M��ŇV��ݖ�޹E�X�N���[ѐS�s��̱e��!G��ᾑ�3�RDN�=yE�xZ��8(�3[�E���`��0!a��JExz_���]�j^U��Go��7��Du�w�ɢj��Ӂn`u�:n��c�E�`�Ў=�wWq��C�(�/�U_�o���brX�0�o�3E]�H����3&e�k�@fm�p�P�c����TZ����r�6�o���c�؊�i�j�����BL�Ib���d�ճJ��v�,�(q��j֝�<��c�H�[�5նz�������a�}��0^�)��\:6����X���m��ͪ6����"/+Kr���n<:2a>"�+�K��Z9���\Zd��W9ٛ5�}o��3��gH1M6�7*5�VuU��j�]x�P㎆��hEF����
�T�#�5��-j�ʴ_G�+`��Y7�!�m��7��q7�9���@f�f�^��qЫ$�)>�GR�����nC��0Y�\�,�&�ގ�Z��
����,�M^�ht�M��(6����|j�|�C�,���Oa��;jq��ssz�0z֪��  �I�*{l̺B��R�zp,T�j�+�w+	0(�ūU���x6�j�eY�RMV����ǭ�V=룥+�l�vt�s�I#���;+�-��,�s��1YT)�C���j�o]��ǀ&)�-lA��������[�v�b�����(�ki�Y�^�B�i��e9K�PM9G7ơ�[*'p�{S��Ez���Yt��h�K�u�1���Q���AO�V�o8LO\���@}����*8�5+���Wn��B<���AQN�����Y-,釸�xqmB�`F�j�G�d+��#�t�}2���J����[�Oh�BM`��f��7|6�K�Ĭ����[���VIَ��
��w�Gـׁ�*�J��a�
���X�?Q�Z�]�T����|���mG����J���h%f�a0�V1�����Ya��V��`"n��7]9�y ҧ�O�]�9��
�)+{	����r��Ab4���@q�q�R� �����krh浶]�!��[f�!Mq��!:3=�zؽ\rur��g�n�պY�X�\חW�j��g����X箛*8^�{� N�Obw �T�&�8%ѴtfJ�@ڧ�����많nN�5�Ogt�����]kN�F�6��rlX9Ԅ�����ɝ�Yy�θ�W,sc�pɼnH��Y8S�`v�ҽ����3���`,X�gBZ����tҔch�f�6K-��e)#[%�鄀ĥ��ݹz-g�ˮ�<��p;CFg%ҵj�*:Wd�y���\oe��9��G/[J=�0�;v9�6�x�wWO]��1��.#�%����c��Al��sv��:D�|��=�D]��r�km��#�v��b�\��DJʻ������/��ՆI�k!qv�Ӷ��^q�G����	�O޻S�f�u6���=e��pM3���Z#��	�ٖ���2�gz�{P��-n�X9�Q�gf��V��E���^m�k��:}K���Ň�<��Y�2K��g��gu8m=��=�WM���`���t��������%���k��{l�=��U�65ܘ3��� �C.��lIy�n2�U9]��7����y������k��-�n�E��MeƸ2�,"��-S�j��"��2�p:>]Z;|�҄�z�n2�&�Wf;B����s�1�׀(��{vv.��y�촚w���X	zs�Lb_'�g��v�^�
��ӯVv{i. ���Aa.�ncamҺ�h-�Z��#rh������nG��ƹf6��fk�N���9�^I�vLOk�ywW%��ͬr[riNb�Ff�ݳ�N�rM�֋�A���L�64X�[s�������cg,9�\<Wۇ��plб�4�iݻ`nd��;�%P��qv��q���n8�Ԝ7=����[Sݪ}��Ϸn�y��%/]�pS��cp�&���ѥ�*��\cxs��`�.���Y�OY��1�s�.^�H��jG�7cB�o`l��u����Nt�n2	�qn�x��c��3*ػuu=���м�j��KB��L�1�l�M\,�-8�P3K�.)
��ۮ-��OhA�)g��.�V������5��y�Z��k\s�.\b���uʹ�m������W�c=����×W"Nz�t�LGp�9�N�LZ��턖Lmt/��lo���2M0���o�1��)�U�y槇��*{��Z�YP�#��0�!���i�ȼ%\^�ۄ�e�$C�4Am"�� �ԫk�H
��J��T^~�$�o�<8���t|��2
�E��
����͌C�%��]�u1b�Rg�N��[ƨT�yH�[&JM6����V�wd�y��tPM��(ix�Z{_��Mi*XɢAb����Yip�o�_l����������ߋp\E��vj]EΞ�^R�ݷX&TU�rڵ����9����į
3J��ܹ�?@{%H(&�h�_ZK�&����\��U��Z�+t�7l����߮�;}~��ņw�?d���ֻL�Y���~j�Օ:�W0h��8�#�#������	�s��FWJa-j��K囥���B��:1&t.��m;� (�8{'�C��R�f��ܬ1[s���|���3B!��=���,�F�}/˙�FW��p&�� ���bؿ�}̋��s��}�t�C�XwM�HI1�ŏ$�R6M�	�O}�%�Ŋ)��^�愨�;�	�L?^k���KQJ�t�htέ���{�Ɋ�v���B��d�&glys���-�u��;qd�L}!aۛ(^�nW���-��;m���[΅�Cg"!r�5�"I�ډ��f�#"�9=��\��|'i̐!DwBڅ
�u(��GTE�0��w����HSO�J�� �NF�9ű �5j�w\'!�_m �H�3	��va�u�Gw�^
��i�/G��F���E2ni�5�����<���1R&�M]{��@)��+ƧqY�Ɋ�*�w����,�x��{^t$�W�	�OG�<f��/�Gˏ�)D�*��i��<����z�=�S]��Mh�t�X�P:�A��v��rz��c��c^',��;��D6�f���p��u �l�]��"���j�y�BR}�>�pS�Ɗ�f�`DQ�r�VP@��n�-�S�`�A�Ʃ���32��{-�n��b�i��|6��/(WN�1X3���w�T߳��CI-�{E��Y��65�ύ>��ƃq-H�2H�rH��+�a��נ��h7U������,f����S=Ce�G6݊a�P�})�`v�?'(��f�[ٳ��%ۄ����Q�`���<�^��k�l�%m0ԁm�ؕ�&ݗꏊ��gZ��!6�}X3U��
j�pIE��p�M7���oU���6�y�B�
�[�#��<�>�ϗ�k����UXtYY�=g �׆���cc_TM�I��4�@��UPѣ	{=)�DW�{/eov������#��5��6���~��m92�0|�w�0F�)�ڗԒ������}[��zϱ�!�J`:4��45��h�&4,��l�'��mؖX�`Ěi�[m��N�-��EH�@�����"��}Mn���RS[�2����f����e�GG�V��R�a^�t��� �ۡD��ɮ
R�%FW�q�`{E�@�r촭ؙ�uY�zP�sޛ�{�r��-�:�<�[�=�X����<���.�LѬu4���E��S1�c�P �+�U�-�x��*q~�o�����1.�'vs��X�[h�6�d$����Oy��b���ڰ�n@h*Mi���x��]��㻫��f���q�o�ea^���8�]�g�Ϲoq�|Sg�o���_����{[�RT���_� �#K���`���N]�{�]m��*��I��g��k����4=鴘�z�!�BHva���#s�����h@�1��<k��C�Tx�j-)pD�z
�.^�k%��S���7��B$Dk��j�͓�k:�Jv��ɞ�T7�T`�> @ƒGyubs����A��2��-��n��a�� �:�	1I�A	��TCm�]fCӓ�o{�cqM�b��ҳ�H���P�||�M-�I��e=�f�D|W����C�{��}I�L%d�$��d�>
&�oY�I����Z��3~�q��KEQr�y�h@e��(ڕ�8u�eౝY���$�vO��c�>ҋ)'��#mŰ^��q�G3�_����"���َ���%��,�lOتU���g�򧜬Q��T��ij�|O�c!�.7i�Ǚ��w��E3Z�������� S�Y�����.����Oz��`�e 8)t�o��H��Zg��(�.F�
� f�1�֤i�4]�i��H���Wlz�׷��;���,U{ގ��՚�iB[:�+<�H'c�p[�>+1�v��usYȄ�t�{��a�H�=���L�Y!j)݉XIwn��tn�d�B���j_������ֶ���V��t����y��r8�.\![���Ýj�y�4�u�,�D��[���V�<Z�����ϊ�kt�]��]�nE���۵�I=��+�l�\���u��Ԃ��;���r�g]e��¥1�K/��B�c�\�<gj������nfs��{D�Z؜����kv���u����Gh�-���][م^�X=v0��w�e{o ��U�W�����/�<�]�)K-��<�H�� �Y�J��y��ɗ:Z�a"4�p��#����tH���{�o�
��LH>�o��7�#��T����S�P�-��8i�:J]h�J�(��*w{Aqm����)�W�&%S�{i<��;c��9K�TX�KE�><���w�ףC�TI�9��̔n���9�y�Mow7Fuf2B�P�$*3�s-�T]��(^(:e�B�����B����;�[���΍H���׀��ֶ.,��t�M�YE:f`��V9H'�3�<n�^����M�k���n�)�؝�c��v�/�Nr.��M:m�0�Q��>��>��j���⪬�\�,�ԫ�܎g	�r��dK��*�k�a�~����ǂsv���D�����m�o.��]�GJ���8T�q�<�˒�hgN��:o]��lnm�=m�:���Dj�w~�-�8����U�� j�:�K+�9�_��$����᥊�_�,J�jH��ʗtG�Η��!� �)�ɢ�	���%H��;�U��Y�L��5zL�*a���g93f�f�n�;�X�m��{��t��{ĩ�#]xᘜ�B�g��
>Ar̗�m*U�8ZXQ]�j���`i�ٿ[��=c��t��!�w�M�+{[��<��,�N���`*���`�T��x��ys�>ĈT�t� ��������O��	��n���OW'�hzn��<$�:1��$F�z72z��%�Dn�W���2���`��o��?B%�<��\@�/�@P� �^�U��Wu@���O��C�L��r(�uc�؀�/b��W�p{ɑl'��Å��W+�P�mu�K�l�������6,���r�-�K��^�ˬ|������֙b��t5	���W�'��k�+�n�cnj�F�Ÿk�>�� M�
u��4i)�LV��xݗ)c��9U���� �V��|4.���-�,T���n�{��0T�/p���(��E��A�D�RlT�M4�;[��,+(�a�=CY��=�{2�]Fl|dǩ͝��W��#8���c+w�M�-�E�@�3�W詬m/k�c+Ufh�v��{־��6��+Kz�����Mf�GR7i�;�u���S��ڜKȄ��X�B��Oh�Rra��g�mRf��;�C��AB+�+v���b]��9D�����N�t-��eh��:����yGBZ�wE�9I�ӻ,i�D7ݽ�2�a�l_<;�>�C��ךM+������ *�,��B�ڻs�?jg�� ���7y�p��68����ow��E�⫣��g�֪5�<���ΓF�s5�2�m���g__Nڜ\
\ڷ5̃��;I�Q��}�K ��b�]۫ՀՀ���;���SnU{��w=��$ ���v[q�\(���W��6Z�C/�xf������IY�$�٨0�	&�*Rm�՞F�i���Z�FK�t����fR��=�J&3LzU۹t�3���B��vT��7f���h�N�h�ʫG)�������e=�%t3Oo�D+gf�����o�lfi�A �_!w$4���Em�p�i��l��i��k+��z�^��~�Lc�t/��ȫm*�M>v���#䃦{ɉ�u�[�����I�Y4Ke��4�,� �k�
6+�dE�(��&���\Z�����K;Eծ�q�ًL��n��B�n��b���ͨ�t�0�I%�e����J#�ǝ[��﷈ڋ������<1�t;�	J�T�!�zU��r�B����	���=�D}����7�pҾ9�s�I3��>:�d��ݦL��+���u�[=�z��Y�u�x�z
c�n����(�L軍�~yG0؞���&�^��Vp�����%�$j�5&ː�J,�L�[d_L�U
��G���w�F���P�钌��>m�5��{�;Zr�>Û�h��l�v�#<��i5Bœs�/Ws�>�3btyx���wB�)���y��*̭��S2�����őYpڇ)�t�H�ILڱK�.���u��γ���r��
1�BV�_e��Wq�gr����ӝ�>"v��KW �*����[']� ��D:	&ةb�z��,j������C*(S�_���{�6��ث����[����c��\kV�����T�JQ��(�����P�V]~��4��Lϳ����,��UUtj���NYJ:����r��Kn�mL6*s�º��$Vͦ�($c"$#���k�a`[��bƻۖn�p��|;`v����O&I����`�T��a�x�v��n�M�0��0�	���qu�I^<�&��Ms��l6�uq��nZڭ,�uۙ�E�6޼vmB�O`�ӷX\��*��Ɯs<�@�[I�l��Bf�\#UlE#,��Xhڒ��l��Օ�m�p39D�mu��-g���5����k�ˍs�9��.-�Y���;�4��u������X2�*8 `�b!���P�^�e���/n����Z��Zz�jd�V>In_#8xvm�F���H!M��"��ծH.쮠�e�h�-�/�}擄��}�m
+9�gp�UN-Ӛ3��nyh���K:a	Y��([ʱ�j+q�{v=똠R
JȢ	l"i��!6߅��>�4���Gެ�3|Ħ���e�G�� z���˽�3goRSJ&��4эV�c��<@��T��f`��$��~�2��aWR��YT�o�՘M%/tl�P�I\�)Uʾ�(�omଲ�_G��^�`���-�P�,zCCe����~]�����^���n�%Y���NW�9}�C��(����DgxV�2i<T�~��H��q��aRkf��#.�V�UT%0�Yta4�1�mlo�6mB�٤ndmt�{PM�xz5I�T�w 7��45O�A���Z��Tq?�8'CV�eS����u���[ta��H/xs@�H�p�At�8��}�4�ף�\}�1\���;t���d�]����'����Ӗ�<����y ����2y�1g%��+y�v������+�0)���S�g�2�2w��H]�8B;9��7|�\����я���̊���X�-Q�Bd�������Q�����R���c��6S��]�/��67F�/�y��醞���zr�%C�ts*��f`�8��s\fD��{����f{�%h�Ɠ	k͉F/��7����I�ۨ��w��~�� Ȋ����ܺB��R{�H	$�E&%=$�y���F�yB��j����x�J^H�.z;�;��vS��n/Uܰs�Э��}3�G�Z��B ˢ�I�a����YbJ;"�v0�c�.��ͳX��(B���Bn'�s�dRؐd��}�tM$��qUfrK�m���2�5�4t�߼3��D�Jc!�=W�v��f��U6� (���b�`N��u�U;��oإ��P|}���I�����9－Y�o�|4���o=[X]a�anK�-�bp�b3JH��葌d}�p���7g¯eN[lBlE>�=���@ӓ�4)����7�|ײ��)Lk��QfĞF�u�q�#�룽�E�ǻ�,n�N"�ZMt�RZ)��HBF���6�7r�q��n��ဲ�;��՗)�ӷ��ݨ���N��>o�o(���ئh��E-kQ^z܂�L״�=w" �g�����v�N+S6^�$ݙ)҈G�6|k���tp-� �(�I��r�l��ѻ��=	i�z^��3i���X�Ma��X2������ �ʾγ��뮫�v�+:�Ҕ��.�K��7f��ep�Дʙ�ym��)^&�����f˾ŐX7ԛ���Ǥ~�'uw7����M�X|���%!),wo�iyM}׺�#�=ɊCº�vq��ةP��n^��XJa�b����ҕ����AB�m.��Z��c/�l��:��8|F
#a���@na�&��)Vˣ@�"�qC1� ��g��Q�������f��Jg_6˥�db�U�)� ��LlL!ưr#��}��.]�f1�P�xo��T�BF�E��-J��Z-�]��/t*4�!�moY��W�F�,r�!��w͋]/�=Ւ!����\�K6�%^g�=�ԁ�[��6�_3��e���N;0�w��[ÂU���[g���r@�NM�x�C�*iic��h��65 e�7�т1=QuN�'ݸ��Hu�O�vd��ۼ8]0l����Xl5$r
�h���?��b��Ǌ�VF�}�{5N�L�R��h�ɠw@����Ь�F�U�C�qLf�l�v�N��������*��Q7��#�ȜhA"���~�aF��Ix�k��mծ����\�H,a&���H�*��q�[X�����k�yL��✙���]��IJR�BH���k�&E�w���'Mޒ8��r���Uf��Vi}&�%��q�}ns�m�d�0'���h��|=㇍��`ŏj3ƣ8`�<�<q��5l4���s0�������J'p7l@`�#�'{��v����\���l;�㞾������]���*o���=�ud,����7�Ԧ�G�����	�B!�����=9޽�n��g�o�Z�y��t�̂��]a����IpK4+�߭���$�^�~��慜�v[�/�I�"�0�fa�=�Sb�a\ؿ��7���\hh�Ǽ�{2��ע2+�D�4k�_�_9t�R�)�(R��%(�I����d�̫�0���>_v.�'k���]�h���
 O_��`U��1ew��:u��ұ;k=
�nQ~7���X�ǌ�+UzaP��!c-��m���]�J=�	~�Q5�.�i�U�I�u+V_�]�he�ňWyK��ai�@�@�o;�����ss�}�9����~Ξ�ώ�x���|7��At���_�:�]��o<ʥ�ôy)��m��_Y��{Hb�h]6�k�J[sg�擙��S�m/a�:�^Ÿ6{g<ܛNA9Q�^�փa�;9�Y�Έ��;�O���5L�c�\�o����dhy{דY�zq�S.MhK���|�;Қ1�L͇d�����6�=*��V�������~ʳڴM�A�J��a�I�k����/���<wG�'/R
n�c/(���M�H�M��G̻Ph����z����~T��v�j��WG������Y�i_,�;A��Տ�"�!�$[199�:x�KC���h�y��C�ѩ��|�sJ���t��$�&]G��o������vR}�}t����ƚE�]*M���l�{]��!�Ԕ{��<_{	�����Ч�=�)#Z{����$�3����U��p{Hc�ӵ���ױ�b���\�\᷷����Ț����p�؋�f�r�*)�1�"�J�K���K��+@]E�	�t��S;xW.�����Ƿ	v�@R��H��6�:���u��^�2W����z��fw���u��Tl2�ӻ3����;]lo:�`�.f�Q-��`�����l���Z؞���������<��>��{X�M����PkbU*����(�]��^r�v�m����i�+iul5f�T#���������]s"go,g]��9�֭���|�v�
�ŷ\��M�]�ԙ��b;�'m�mv��,�=������%v���#����\�,0bHO��_�	$d����
;˻Y����c"/RJu(�O_p��]7��f3}ޕ�z�^� �Y�J�\�m
A��I�S���sG�f�^��[i��;�ڥ*�x�Y^�7H��[I���璥�1L5��Nx���d��-�B��#�f�:�N$9O0u���i�t=sܒ���Xx$�J�%G�*�#����iӧ츝F�� #@&�(�Vs	8�� ��s��\z1��m��E�g7r��&��N~�Ewe�MwN���av�҅��.=��sZͫ�h� I�2E4%��i׫�/>;"�}�U�8&ӗ�58����D�G%�!�j���i{�<q���cT�����������ڶ61L�\[m���gsѰ�mJ�q#6!t�����]R��7��y�	�"�$<����y���
����蜤�{'	��M3�`N�z�C����ZN�,�+��
�n�Ln��}H�=��1M���0RR5����-�=��{��2��+P5JW,�r����{4�C�����)��}���W��bc�w�t�g.!>6���v	� �!Sg�a�.�v�.�w^TY8�&}�ݑs/ێ�B�n+�%���a�� ���a����M��,�U�H�8�X��'��P�'�Gb�)At9u�=G*�F-��[��c^{��R\�Ð��m�����t[4�]2�R/{���!د��C��Rգ�4^r�[�6�f�6aQ�s��U�&�&�.=�47�݃�zn���ЉS�i�I�XpF�� �\��6r��ͻ�9�r����ݡ�c�<����ϰ��I���r��G��	6��k�j�����=z|m��
!���&����G��2Yݝ��h�a{1��X�m�웳hPI�i4&���fh[f]˦$�\]��m|�4�ۜ=��%��r���X�	Ϙ��{�.d�w�۶�kϯ�߷�0#v�&���R���A��8����#;*eNS�z�I�S|ROt;��w��+�#�G�p�pM8g_���k�<��g�H�I��b��#�g�G�Q��z��}'�TN���n�m��{N�;�.�09U��B��S�H��J���95,4M�e�<Q�J�xfG�A:u ���v�2f���t�"J.R�vlA��0�x�����3�ϔ�=��&U�j�H'M���I U�y�VoI��s�r�{��a�����ݏ5�u�W6���e��5�eb�=��g���Z�y������&�:,���I��m硩Z��)�r#�2��/��˞;͝�.LR����`��Y�XV�u�Փ|��r?-z_�~G�C�ڶ����b�,����]MF���.T�F�\�B��)�N܆�uk* �L���!]��;ҷ�������u�F�rB���y���W
�~�YR��E�� nm�p񻃹����Ĕ04�[=6��}#��kf�=ʰJ�0|�S*��oKg�{K�x�j��$�︉~��]�QU��U�W����"��ۦ��ifE�r�\�m���ұq�7���AD�P��}x5��PX�k���V��g� �`6�l:t�L糚a�/O 8{�+����u�R���G�ub=W��%Sd�j�}wre��}~�&S�����: �g8�O�w�7-^{�Gƴ#�������9W��cɍ���B�l�4guY�]Ll�$J�m6sdJ,0�x��k<�Y~�F�	*T�D'@��ۤ�I�Q9%��{�u� �xa��Rյ�r�j�O�]���U(£�9x7�u�2/�ɮ�}������%��iu��C%Ƈ(W������s�S�zmu���N��C5Ή;5�Kg���ЅS\�v��2�~�7�V� SbZa2p�X��5<8��S\�Rю,1������N�9����$UFQ�����in!���^8X%钟#�3��������,��� ����,�{z�z���S�����}�pHb"*0\m���ތ�it�-rL���|e����#����Z���޺uf�>��u4_'X6.zl>$P8,&[�p�C}{8�{6�q�=�YcB7M�=tl�=��wW�X��8�lr;��yO6��4���-�k��T�TۤPI����%�w^��CZ��u�s$��y�p���涳Mz��5�U���='t���S��b�V4� 9��G/��ySڗ���%���HW-w�o"���'Ҝ��^���ދ�����t��ƭ2J|[�f���Н��l�Y`2��~o���W��O=���Nx�fi�6ոG���>:�0�ء�s2�B����In�ׅ8���Ol���6kYpʑ�шcp^u�R��p�۶�t�\l󐹸����|�*�Q��]H�j�9j�uq�F[m�<��j�܈R��@^cu&Xź�ڒ�YڻmN��8�W<K�jާ@gW@/�wn/VN|�9�7[sl��stu�ͻM���Epi��C��k�7E��j�$]���S�8���g��֪��K�C�LqΡ8��.@}d�ٝ�^'���=޴x #�u�S+	ރ˄Im����(�+�U0��0yƷ�n�9t�l��@>�0�U5D�ͽ�$8v)S�'^��^mF�yK�>Ӟ�����ˠ�=�S"�r��r�w��ѧI~�ާ9�|0��n�FF�MóO,���˘9�_J����t͏�(#��ٕ�]�L����i�"uһ�jp�,zw���B�K��v~|�%��<C^����P�]��w<�I�As6��V�K�^H|.fS���_G͟IO�.o��h+�D�,�����~Rq�e���W�!���Y��z�ڎ�K����3��Sz�ک�;��ڳ����e�{w����~���ҭ�mmc�RU%K2A�5Ύڍ��h���c�=u�)��W||��ru�Q$L_~���m5��om��;&���uA{&q�t%ں=�aUY.�4d/�\M�<�]mk:,�t�Ad�LI�
M���*����g�����a�å
���í��U�Ǝ��7Wd�g}M���J�M=�;8�p�%�e�x�ܔ�(�_.�$j��mNjuN���v��hm��Y��=�(M$�E{t����(j$7\��3�]���^[��y��)��i �-�^�q�1(E3ǥ8�C���1����o*^����h��H��'�ͬ#!���d��˭\��a&���x�1�x��fS�#���_C'3�XaYa�s<Y�}��p�{i��� ��x�Vc�	�6�`ăB�d0��e5������q���/v��v�R��e��Gmj;7��W-֌�������K{�m�ڬ`����o��6Z�|�g��nu�c�VB�[Xεa�`�lU�.�Bw\���%6M$Kl�����n1�=�Zg�s ��ʞ}�q�rOfu#�1RM�J������"l���O-�)�j��Bҡ�:`��L^�I��&b�D�eG֍��.��Z�b�m� :�p� ��悷M�Z��;�wp�RHy�����
PS.���I�T���[��W+[cl9Lo]N�__�ߐE�Yg��M,zeK��=|\�e��������t�9\��k;ge g_nǽmf�oMF*�3��Q^>��K]�w�]nV7E.�����A(S��h�ZM�8��&c�w�^?��Y��0�/�+n�C��|$���)_���5�j�JA�n*v)z�N���󺓍t��Q׳�F�@��̄S:$�g��/U�@��6�9�qk[�F�����W����n:L�Hc��Yjyִ�݀o�.��rAW�Q-"i
T�n<vy��\7i�����E�FPs`��0Fmt��tj�(�p�,�!dȤB��b/>�;O<��#Y�-S�P���Y�ĵ]�^�{I����=;�Q[|":4�e�MHn��W�7�͇����W�z�=x��o� ~�~�!�'�HrR��۾�#E-|z� ���>y(��nf���J�~�w�#�6QO��"
)��;�]��~�H#�A��=��Np{-��S���2���yQ�l}��>����9IҢX�U�.�6+��������{�ו�u����}����P���]��s�m��e�8q�:�����DAYQ[�lQYc�7���{f-�N��ɔb�/���E���Q�參�p�V�Ec���:�+.����}�C�^�F'�b��y+J�n�w2�E*�ɀ�!&f�(�֟54E�Z�\�������ڮֳ9�^��bN�0�۷A��w�_�QT��xx���O��@ͳpsO��FY�x��s�cy7�3������"	�Î����:󥞳+0�~�d֨�E�\�_��W8�{��@vb���|�[pOA����sw�}~�މ.��J|�Ͽ��%�;�GZ����)����ږ��J��M7�߶���n:�� l�.m�cٴ�G:�7�Mod���c�a4k X(�[�}����'����%(��&��ͤZJ{*X��-�T���>�LQ�I��@:F���I�`ڳ�P!�Û�-��
����֛��ܩ��}�]�
���&n���j���>�9��;��2؂H�����؛4�)};|s���0�F���l��0������Qwm�{^�<(:α�]Y���r��}BG����U��c[�{
@c	weTQ6��8���]e�����n�ҷ�:��'��]�Y�*������l�f�I�����)��qܗ��u�rP�9TT��ﺶՙB�(�|�L�� A+�r��ܦ:|A�bIݧ��/O�};)=v'�I���iYۏuR�&{��ւh,�`�6��F�ژ�-=��z��f6���g#�p��ZuN��o^�ڳR΋VB��mշ*�;1-�˟���2�+ �d�n��f�.u�S��io,������u��}%�d',�`U�{��>�m-(��冦�v3��3J�J���]�6��a��ݜ����{�"�����!�1�/I����ϒ��;�k��%!���f��JP1��9�&��z�@�7���.��q.�[0{ip�gvl)3ц�m*e]�-�w��C�Z[h� �f�n�R�[P:��S#�!@�N��q�٧I��XWL�v�*\Q�z)�Jk:�U��;_ X�D���IV�:kX��V��k��V^g+0�n�N�,m��J�]�EXYG�]=�x��lW,�9;5�BU�:������֢�ܨ���r}H7�Vլ����[���׼S�-Χ�b(g`�u*o4��;�{��.vw^�%�\�0����.d���9����l�<�>�
m�`�!]��d�au��{]�;6p��:�R}��q�gʟWj���X]JD5C�{ӸW+��a�&�2M̛�SZj6�j�16�m��Sb�[j]�u�t�h��E�i2�4�ٱ���4�0Y�ۘ���Z㹬7Wh-,v޷n�̷�jݥ$�C)�E�&���eX�\��n�^q�5%
p�v{@O=��;;/\��7N��x6�\����͢�͉ure��c���	��2�Z�
���v3]Pf)FU4Cl)j�x��������=)���^ �n��7C�ћ�꣉H�m��� ��ML�am��p:��^���MݸޯE�w=�AÑ�z�Ɂ��������\2���㜌l�Z�7/H���ޱ�D]cESqP�����{]����yލ���]b���
ʫfef���й�qi�6�v:�d{u=[k�w6[vF��Y�i�*�h܏��y����.xfx�.��.�l�ے��{=�cz��uV�[����DV��ۘ:�c����z7��];nh���s�en�Af��m�5����q*���]r�"TlYZ�Y�-3�Q�34�Ε-�l���-���v��l$�&��ag�kq�kp���7m�c��X�ĸ��뵳�e_n]��dJ��Ė�iESiC����t�]�vwT��7=U�����ԗ��d���N��/S�#Jk��cAFK-M�:��R�븥ᰲ���qVCiX�={��ۍ�׷]N�^�c��sŜ^A��Rn��Ox�^�d�vv�`	��@mm�q�w�Qn�kǑ��̐���u��4�;�燫������m�=�b}�u�=�p�Oc�^�[���B�&9�7=����ͼv{.܈ګ��'\�7nl��r^�t��6����um��G����	lXڳ%hf�[)�b����.��*����uTI���H�_YnݓA�d��q�qh�&�7D�+�.Wv.�[g����۫r��Ss��掭�mps�zVH�����e)�ˣ�� ��6�}7��+/Moo͒��n�.�;��"��&�z����.,�SFݙ�Ѓr	T��+rK�Ah�����c]�͸{>w-u��\��k��Įl���q��|�v������w0�����sKV8��Խd�V��Z2pk��׵G�9�j]�%����-vE���ln��-�m�zC9�=7k����Krmɉ�sfBy��Y:���u���j�VQ䠻s��;[t3�z�]v8�\
�X|0��MgG�h��L�z8�օNխ�u�������Xx�u��B5Z�x`ݢ�NcqΪ�!���e.��A��������=��2��uFWV��EZ��뷦[�o�c�3@���G�����1�<�{ΤA�R�A��AR-�We����?[�+��+���룝�#�gi���Wyͽ$WY�2�oc����)c�v��)z�*�$m���=HN}v"�G������W2����ʏP*�ؾ*�ny����+AW����v �hPj�i�,-/���P>U{3�Z{,n�y��|�_��+����I�H����0߽F+is,V�+o�I��t�t�1י�$˿e�=�=>���
�j��F
̚���6L��P���eʛJ�|~M�s�����T��y=F�s�OI��\�-�����Z���Ocu�,nȮ�+/[���v,bh8z$a@ab	���H�����:��W�1���fWgx8@�j������`~�"$�Q�{�N�I&�H��M{<m�<���M]�����A級�����IaJ�ݺN�&.�5���)��r��h���$���能g���u����#���V���B;��ۏʽ�Wy���+2��z�(�ee��5J��\7H��+1l���R~I�I�4[j�lk��o���M�ޱ�c��8� {�11Z���o~�Xݷ������U��F����)��
8o/*��!���w���@��T�=Jؽ��J$���T{n,�'(ޗ�:���Q�`_8ﻗ<�/��nY�΍�80=O}�bX�'.B�ިO��d�쒸�ͤ�D�ue�g�֘�}Q�ܹ��vb��U�Uj�p��{�y}s�M���"K�2�1hSf��KY�>�]uۦ�9]ָ�<.�]j[�18�YqU�ң9�j�s�����9x�#�9k��y�7�??�X�n�����L�!�މA[z�d<��f�[�]�\�jO>�|�T�wU�=�����b�;��1y^}�Y�t�K�uR�
!������YWd^�NM�u���a�I*d0蔅���q���7ػ`��Bl�?R��=������=�@Ċ�
gZ�/
�R�Ə��O�Yƪ�u�r��d�b���t�t4d��`1z�4Ja+��N��]�XQ�lW��5:j6w=9��˗�����i�#@�	�(�R1Q�ߺ�Y�gM׷o��י��w����:�}�8p����	�[�(+;λח��2E���m��E4I,�T�M��p����D�����v��&��؞Yj�����F&G�in��c���u��7��}X{z￳�ڻ2�j:\��k���0ѷ;h2��tU�5�6�s�λnQlkj��4�	����1��_L�I>#K�<&�(�I/��*V,׼6	۵e^2=��աhȏxuX+���i4�j�M{=2|}z�T���l�=�����u� ������V��J����3��ݸ7k�ߙ��$Sl�L��c��l��fK��L��!\g5*��A1k��vO�%�+,����p�/ �4�	�TAn�f�iߝK{�-�S'Z3�R5~=�J�gd�\��%��S�s�H��{�2JZ|�WX�6#���(뻸�Sf�6�����yV���6e2�������A�d%�xP����J������ͩz�Ӷ��C�Ɗ��QD:-��x0�mu���S\���v��[��1�������ڹ$�h�R��0�5V
a.������ �X��g]�]�V�����b17�<#(��]�����2����)nыAƵG�$v�[4��M�.��%��A{,��^����4,w�/�z��-�Rf�I1ō��c�Á��l z��N�w�^gyћ������zs<�A�u�K�;�Ձ���{U�1���5ieJ�Ҙ\2o�Xf�.�2�c���)����k�M3x��8���e?b�}��{:��#ӷ��[��]�j�J��ޜU�A�Z`2�c��$Դ�mn�X����]�Ǯ'}��/�v3c�GA�4���4�]���32\
�K�����t� ���^���]�>�i��u�WVb4/:��ׯJ�%p���YzP��;/.���6����]����+mW��r����
Y}y�>?+V���;�YwD92�we�'\��p��h|r�u�p�X�wONw����2d02R��bM�s98K۝���_5^ �âm�q�Λ\Vy�c'��0�v�J¸KP�,�܁�\��Ӹ�K�����(=����ȸ�̝|H%�X�f"ڛ5u`1���e+cd��S������:����m��Z�w"1���m�9���DD�3h@��16b��r\]�Z���w����ݳ�g[���OW1]vn��ۅ��֎K<uÃ��tm�L;���F�Wh�O-q	ֻ"ew7>��%�u��Ź�+k+�\���\������=y�{|#Zv��D�.������M���o5��B�{e4�(̆Z^�ވ��"n�so�[T�)�N�-�]��gX�{��H׶c�8>/���S���s��Ȝ�@GG�*��R��w��(�ѳ���ȟ{$� CgQ�`��	�)εvy�x^gz�N;�����a�V3i0m�D���g]�-�l<o�t�H&���6������ݲ��V']�Ut�8�)֦����3�L)��Q��f�`>N��0�F f9�d)��8�����Nlv����Xy�	3`��㓮��!��3�纟ޝ�M7	٫�n�t���Y�ro5�6.�o���6��ˮ�gɘ�y�֫u��b���?O���ú�	ʻ�ܻJ�S�ܶ��&��=����X�gB����*���:N�;ʔi��4���H2�3I�tpu>�]�����}D���rf�[pإ�pe�.�*���Рz�*i�w�g��V�;��n�g��欹Z�'��})S�r��2��U�Ez�����k��*�0�7]^���Wj�m;��ODA��y"�e�f�l�Kl1��#3����ƙ���|tW�H�ٱ4���b�Ύ���e��*
��p!����,��Uq/��}uO�;@�Yܧ��k.=u�M���m$_s�kۺ�/M<-�-]u{M�1uwyC�hD��@	�$H� �������7�|���m`	���'���	��J �[��	�';n� �I�BS�v��t-����h�t�meY��z�;a\�A��r�[Ѻ�t?�	��G�Y�n>�kk�ؿ�_��Pl�pDr���N���In(�ң?+�O|����GK�\��x2Ԕa��R,�,�\�s�{�1g�$����B1Sl�a���,XҦ�^�BU�׀řO�O�9�pn�i�%S-$�l�D�=�"w���o�������W^�"�7MB�O���,бw�fm�*`��W�tܹL]��F����"��j�}ڭJ�}�(�X\U"�Y�{+'~ɧץ�n��<o���L@�e�(��z񳞛�r���V_5�{ N��]��go��9���=W=ϗ�5��\ꝇLpn��\�,�L��.�i�|�Irټm����n�z���vt��t���(o����'���&�>|
�� �$�e%(���H���=k�y����FK�pŖ�3�jM�ՠS �q-St�a탆�O^J{��T��}p�����fgሀ��y=`��p���i�[�<�.����!���C����#�'��{�T���IO��X��	x=�.y��wmt����3����-Ů���SM�6�4�a�/	���Ơ�3�bOF}�:����u�y����Ũvzǒq��{�#TCI�@L���y��&\��zg+Sh�C����,�y'P��x<=ʊe����7�O`���8����I5����H��6;�jTr����	Yg�頎�v;�{�E,����{q⬛�q��Q Ђ����9�j���"�I�W$�0SD%I��i�?S�}���i��8G�3�Acȃ����6��^�dJ����u�+��]�����&H�4��=��.X=����k ���q�P��i%�;s�^�u;�'&������.��$�s����5���]��O�U�;<��S���ie:c}Ͳ�:.�n�L4�^z�ܖ[�7��� {�E>ab4�Kӵ���&^��x�ղ������\7�$��<��2�B`M&d&�VkǁP�y_&�t���}ǟ��� }{�ѠM���"a?{n��ukJ��>�%m1�7%8�k�kO��y��v�1%�ɝ���9��{�U$_r�Y�F�zX���X�.�����Lhڝi�ǀ��2�J*C�3���=�:neD��]��'5����N��6��$��y�tn�ԯ2��z)X+8-�>��iF��l�;�MT*�hK��c�H�4+��#��:�℧�$�,ms����*�]�����^'O�94�ۮ�^{qvt�Z+��-�X�\=���v���Zw0���S�볨�MӞ�\	���t�a��F�3u���lM�+��B�ox:9�m�]��pW/Y�����gqGMkP��8Mfl�R�v�����w2]��C&�Ȏz���g=<���K��m����ZJ���M�t��
]���vZKx����H���F6ģ'���v���sZ��n.ӌ��TB흳�{$dm�%v��Yݭנ�L	�
&�:��t���2ߠ"�wx̡����w=��������.d*P��,:�.��f����T�T�h�H��a�����d��~��ZT�ka�?y\g��Xw'L^Gb�C��+��c�vV�B	�;0������΀̠A˴JL�3/T�4A�Bed���:�����r9W�.�;S#�=�������=[��+XOÊ��v}od��}j �Sr��҄=Z*Xf��P�^8�ǏgU�t��ya�:�d��1�{������C�V-�ܦ��$2A�[�}
�n��V|u�L��9���z埡 �Z��@���3��lD}���_��}m��=���j�P-�YE`��j��F�Y��^:C���Ѭ�·`��y�jU$�E�n��'D�|73�Ÿ�2����+8�k����Q��V�؂�@m�'c��z���C ��hP�S�7�6�y�
w!YQ���-H���P��(P��P�7Qj��g�YSN����l�}�]�/.�ztbL����w%�ܰ�V��8�}���V_
2'YV�Ig�`���h�2�7�ޙX�j�h�q�/��I;��5f������g��~�gR.�E �j��>��k$����	��{�)E�s�g*��W�/;�=��x��2
h%�N��$��q��D�O��/�+���r�!ʲK��z̭��
(�꙽�v���0�h�!N�[�Z(�c{}����fZ�X�tJ8
�T�ېjEz8F��i����n5K}��V��uL�yR�6~���* l��5��)Y/-�����{6��K �b(LQ��c�<4�8}g=1��\�4����]�wU<�`8*ـ�L�����W�)^~^�q�/��G�÷���|�:E��K���@o���e�,��k҄�e������$����k�V-���7�c3wu����W�v�i.�y޺��V�0\�v�rw��Ǣ�Cf�(&|��i����I�hk(���u-�*�?i�tG�T�)�uc�*H3�g#N�M�=B�ko~#�Z�c�� �*t<�i(9�2��r�:�3��BQ�+{D�:+��4є��O�=�j��y������{;�j��|+�;��u���	t���v���o䫴���GiM��[#�N⥁�6	�&:��ׯ�4�<��Y���6 �x5Bt�H1�>��<�:�f�*�b̭��X�Eqwә=���,���w�GB�=�kV�F��v�՚����N-�%��mC�?f�V�[��)*G"LȞ�{�J��P�Z�w%�:�ġ��T������7�:��f��;��f��;q��\�G�]�	EKuh(�*�n�NyV�?N�&�W]�9k��eѹ٠R��/�]u3ua���h.��;i��rve��x�1��.�����*�;֩�v���E�ɀ��d�٫�Ou��DQY�8K�����$i���ܚ�לB3��ǇZ�4�]t�n��G9��Ʃw&����@�tep�۠�`�������K��t/��P�j��]ϴ�)sm�N�.��S����$n	r���ժ��Ly���q�L���N�@VlIuM�k�Jǫe���6�FROK�����s�]�@�;�v.KW4�z]��i*�1@L�`�HiK5{Iǖ*oh@쪌�����R�A��j�>�/����'��?
I	�
W����L�g[�����b�.˝N�`,�`����01{�w���j��%�k]�����`Ԛ��y9��o6m��)E����ԍ���u��!*t�M������x��>��6-yD��=�L��B��ۿ+�|`Yf��Y�D?{Xg��4���@q�F�痻o/<�2>��x`d4��C1Pf�B���6kaE!�'"���� ��@��\6@ÿo:�p���8hY����ͽ��~�=����@��CV~0Ѕv����.wu�f��'9�0<4�ڮ���f�=���w5<�~���q�ާY�͍�\�S={:��y�C��\n�)�kS�\�e�8,�tN�須�{j�8@�?}|ᾚ��>�VT	Ǥe���t�F�hZxO�ƚ��>7���|�ɟ�i=�{OH[U�� ͚�畁�t�e��(a���T/�˩?�Q�p��CڸG��1�*o�Mm�o�n�����>���M��x�MF�|	?d���q�N�0��t�VD#�7�`|t���݀a�ZoˉU���b�p�ϼ�[���(x�f�A���ς"��m���<#�Cf�ᬈY��G�M��G�3A5ZD#�5r�<�{�y�F��Շ���D��Hلg9�`y��F��� ���~fY�\������h]�c�F�m�nG�U�[ҡ�B͎}>��I�p��\��t@��ϕa��w�DB
����WCN����g�����`\43	����l�}ҵ�h�iKm_�s�qd��ۇ��#�Q��J�!��}a
�8���K����4gt�R��&c�w6vW�"zM���ե�=w�kI���˪��в�CC�tu�u$�ʒEh���.՚h"=��Ol�]-p� x�UGӺ�/�������p���,׈�&>@cy�u�{��ha��P��G�}�X�t�5�TȆ��b5�q˿|���i�XO�3P�-�s`k�����Wd�A]s�(qF��h�K�\������H�qt}�] a�<F:Y8G��<�뾋�G�UY��c��Yo�ӕ�::��P@�>�����f�/7ln.i��ߐ�H�#�\����ڇA�I<:S�,�O�z�ߙM���&n�`鮫/���Z��3�x@$1�/�l���/Gh�0��n�'�8n���3^�hCB}~�`z��XQ���hY��_0X���lг]�{R����t��ﯩ�%�얍p�<�����g�/E�;�ϻ�V���!��F�B�}���tx�5�o�3������h�D4͐!���)�+�����A�ZG�P��.<�G#l9��V����
%��>�N���!���X�4�b�6E�����y�B�J�=�x�h��8jb����3}�l����Xf���flI�ǌ�$?�|R�ٷl�Y�]��p颐بC�@m�@~�lv:Yl@�THT�a�u�h���X�_��A�\HCA�X}����oUlb�����k��2�􁦬�Z���%߫��8��E4�ʳD)���7��n�R����W3���L��F�I�J�u��ƥu^3:L���XtK� �W�Gߧ�|���,R[,�8�t���]6�VSs<c�=�L�Vű�{o)���Mb<1J�c��R�	pm+jF�9���5eE �v�>p�F"qf-�`�h{�5�7'N�7P�q>�x0{�{1��nM1l"K0X%�r��p�r�F�`-�M�/�2�UYfL�fx��A�4��{i.����^��l�GR�m��'X^�=��/f�$0���5��m�B)�ݓ�l+�[f��j�SkZ��0JH�`��-A�HT�l�>��LM}8h,[��0������G=��ޡ�P�^0�5dF��y��}�,�5g�4s��e!z7�s\�7���A�����\�J wy�CM��ΐ0�����$N@�	�XF��F��<'��WC7�K���	lw=߈����A��#9��X��}(a� "��f�k�M}x�Y���hw��*�C2Ǭ?u�O;ށ\)4�
��*!�bhm��K����<'�!��RJ}�,]4��#��4����`p킾�*P�s�鋯�mp��`�͗�UFtЇ���d#����:,Y�51Pe��v�F������"�2���2�4|D9��{9��9n�<�H���~�8t�j�?�t�	�{�x�>����f���[��X_�qPF� H%���-ƨfM��><�vT4���NޖD5��~-��6B���K�#do���/}�i�kN�f���[���t���r�9�+��t,�ĈQ0�:�9�w��㧥�j��P����,-U�*��t��0��c��~���ƿ�C����{�-��5����Ŧl��%6ϭ��)O�Z"֯Xn
�sp8�<��*���5�,Π,Րg�>6y">P�Gx����*+7�t��!�>@w�[�h�=��\�|��@]^9�ƴ���s��f���%��@�A��oˈ}l8�b-ô8k�Bh���D{��zJc3�+ݣ��
�r��O[3�KM��V�� S��ڝ��؋�׳w>��ս*1ˊ��������v����p�����tCy��!��ދ��\!��-5�����XZk�Y�p���Ɗ�9���`W�N�D7!��/I)ҝ?i���.L[�mU���O�����Z���ր$	�~˜���p�����C��8k{����CY;���c�w���t���=��i��g z*�\���!���49 ������c��!�)����Ӻ��At��c,/s�F��i������Y˔,�]��W]"Ow�CH�dA���� �7HTQ\���>��C�>���`��*ᡲ���l��CqP�7�d��[Gi�Oc����hI��9��w�t8C�>���#H�Ȳ9�8=����x��XI���g�g��_��]���V���5�Ziy�9f�i��W������
�g[_B��ٰ�B�k*��yݹ���x��Tt������;]r!&܏����3��վ�߇���a^��{�����wU�5i��Є?�����e�Pd>-�@���A�}���xw��:M�$�8�����+*����0�4�������A#M�`-Ŵ3�|x~8h+Z�!���g>�p��;��w�o���7�t!�yy�cƾ��VA5�B��/-Xy�B��f���>Y�+	��H�ߴ�w�`���!����Y��e�Cy|���R�Ȑ!�P�!�p��`i����Gٮ�гA�Ko�,���D5�w>G���q/�͊I�$^M���*����N�JIJZ���ס��@AQ�S�w�]�E�%ٸ��.d���̦�Xr��ր|n�C����ŝ i�Ѩ:@Ŏ�y�o�ho�� !�����E��20����4������=�z #�w-]>:j�������+��J��&�/o�>��^8<���awI�!��k��
}ދ�!�C���C�8�C��ѓ�9M7C#�c�0��ZE��g�������XhCL��o�z�k�K�r��~$p��B��g"F��n���?f�M{��F��o8m���І��.������qUO�����]q]��vmq���y%�n�E=����s����Og���-�Ӌ�0�Ϙ�4�0��X�Q9�k�oE�,�����z�#O��N�K�߸2�}��$���f�֨Xr�����|:'L����������pw��'���`t���yߐ?.YL��p� �[B��`Y�'s�t0���a�#vv�ZhY���[�����*��S<�_��a��}�ƸF� B���[�A�o���<����S��>cݡ���!�Z��'�� �-��9CH�H��E�G�YF��o�t4�"�NJ|@��|n��4�5~��W������+�c���Ǔ�'K5gN�36hg���b��t�=n�#"�x��[L�*F�Y�Ƒ���!���t�w�txi�}�v�~�85V�z]#mV/��t=|`t�.���KZz��͎���Zp�T��U��?�֝�?
�-�<�T=�5n�]ލF�l�*û�t��[l*@p�1_vtp������������7�;�F���U�ߝp����ӆ��T9��ܳ1�ܒ�2H2�x�B�Q�Y�k��ˡ�����V�==�\^���n}'�w��t'Up�i��ΐ/�Y�a�����h}>�:i�"�F�o�l��_]����hr�t1�t���=�L�}\J��n&����;9K	m֖��K�ɿ��/�c�W��7���~���CCmPg��$F����#��5tp���������o��C�EVY��]�̱v�Y�졆��Yk{1���#�������'��O�<'��)��@�O��WC��|S��M��=�F�#�R���{��a��v�f� t�߲�z�І� 0yY_|�t�<4 &�<�����H�t������m��j6�Ƭ��&� 5�{��W#@�4��*^�J���C������������!F����`��h2qCA�s�cƴ��T�|�5� ���x1DA�NA�y�~�fq����2��/�t8GuT4.��L$�h�w��&V��!�����x�֑güu]�U�ގ5RX��yLU�
��"�(2><�Y���
��2��E$�(a��؂6E��a�������43�g��V��o�f�x�8���g]R5!f�4Hw/��>4� CA�}��a��!ݪh#C�5}��o���9ɷ��7�����kH�̓i�nbz�zaSqb�֘(�N��"R���7��!r&��n���4rh ��!=�c�>߳�����:��K�U��g$o6�9;Ol�t�\76A2��:8��t]z^w\��;���� ���ݎ۶�9t�,�m��4��������6n&W-���*6�JGS�[IQ���rV�i�#c{!�lɦU�%D�j��L ��u�*��9�.5-W�S���p�c�^��d���{d\����[l���s=�_c��.��=t��Z��Ef�.s�e�LX�\�Ү���	��y��5�{r��.����ˮ�5֥����sR\��D|bI����0�F�����@�GN$��*���[�t*��hY�f�g�����C
5��@BH�����\4c�����������'ܒ�\,�C-Y��������ѷ����2N:羖,"	�!���"ύ"�7�`D����@Mz��g��򱶫M��Oo��r��3_f�����7k����|;�`t�z%'�]���#�hq��������Ư8�Y�}�U�#pa�f�&��m���xЇe��p���u�̍��, CXA��f�#���N8p]�w�;ZI�/6���NO�@��鯉���������4,b��<5�L����4�f�8����X�Α��#�/�[dz?q^�C�Ϻ,gz�k�z�6P�L�k�1Ϸ���J�*&�pe�VbhC�@B߷�u�h3AG�w9�{�>��߳�B�h#��W:�����5dC���¯3�*�Fg��=�\47Hփ�Y�0�����7�/�>M�����I�˒X�0F�tͶ��rp��9�ڕ㭛��W�.�쳧n�h���3RB�=�Gw��>�8ǝY�¾�s��CK"�I�*_{�CO��!�hY�M��&���·}ћk�hi�W���_�M���X�XhlT��h���g���uM�Ą#$�(p�!��F���`�G���R}["Ţ�;u���><�l=�n��xQ�d��i�uږV���[Uu��Ʀ��G
zn%:�=A�xnvٖ���H��Hd-ü��;5�a��p���5j�F����oU�֑5<��@�/�4�#��|/W�Â���:)������GC|��~���Lf�a�4�Ak��/��.�{�L�V"�� ��:U��j������ޚo���?;�����4�@E��=\"jd��N�e߈�oBm�؂C��pԈA���9��=���ߗ��?+k��4����Bs���#�N*k�h3�Xo��,����g��[�n��	������ᡞ�HGM|��A|l6Q�
�!j(�WCa�,�@��߾V:G�*���f��ZF�V=�J�w��t4ш3V�Ś~ |~��49�@�A}3�t>�,�ڡ��N�>��m:�� k����	vD�2�o]��u#˞1qqկ6�q���ʶXb�������k��bhC� !��z�Xf��uU����Ρ��y�x�d3B�:l؋��~�>V|6{�;�P���"h|�|��f�ЄY�p��kH�����$�R9NΟ��,Ѐ���3�6/��9����z�D��Tѹ���#9��,���Gơ��9�o��z�B��� qU�43�s��<@a��_>�m��Z+�����]�]��0JE��F�W\#��� Y'Y��WC�hw���,�j�ӜM�P��z뜕����]�<�rX�����~�u5#ְ�Y�x,�D3��!�����L�t�9����v��a͉�Ӛ^�).�S��K�����P}FҨ���a����Z�(����l���a[�11c�0���a8D4!Y3�����@� �����T�	~7�u�u]�'B��B�i����)�����1�ʪ�T{��;���<�z��#���qV�j�5��5�w���3��dG�� �s����1�i�}����t4�f�EL�E��/�l��9��.�G=�B�l��#^��p�I�ç﵁��}�M�{������.k��Y�5aW�u����7!l�P3����h5(\s��b�Ӆ^�,;=GE��fښ�ы���c,�������^���5��}��A<#�T5�9�xՑv�!�:n�5v��:��Ǆl���r_>����q�|8�L}D|Gg�X�����ӆ�h8���3XB�
>?p��I���[�hi�?hB�@���_��i��g2�>��}$3Cs�xՑī웢�a��x�h3d	���;k��0��$LVh+�}��F�H7V�yC��hN݆�	e�q��Et0�ք(���@�*�}��a�hf�_*���Ea<yc��.ny���T��^e��\"��@Y��_�,k5P��kHf���k��(�i�q��4�C?!>鯏���ϯ8>:~47��o��9��2��C�OF�1�3��V��~�0�����|�퀧���sW0������Hg>A�����x��DV����)��^�\��Zv�wf[�F������z��46�:�K"�Y��~w_��~�I�c�@�B�Y��{`�@���|��I��E�v�����,�������!�hr*�g"<|q��̀�����A��Śf /�tX��4��m鱽*�~ |7X�Uޡ��>��Ͼ��G�ɗw
a��@Rpx��q�����-��b�VyȃK={[��tvճ�ì����sa���߇����= CAz_���EBfd�E�ޒ�{��u���D|E����8C8}�w�[��������\5�4�qf�4�zm4MEA��5��P���\m��EH(�-Ŕ0�����t�	�}��a���s޴.;�|g��	#'�hx{��t0�E���>�w�ώx~~��8���x�T�g�|u�a���}숾P��{�Y�AϺ�; JF�� NA�4�F�C0�d{��f�G��~�Zh{�l�dt߹�@�{ۡg���[�"��z���Bw�|6��a_<�d��_���H���٭"���#�0&\&ʑh��_Uw�ƚ~�!ų}��v�;Vt�Ӝ=���b�5��p�>?3��p��a���^#�/�o>XǦ�2�zw+�4o�C�~��6+�b����g�!f�3맄��m�	p$�:kMi��V@�>����iEP�5f�#�t~�[�{
=�L���*� �?
�~{�w&�4R��a����.�X�����B]��(s���������/�(�GEf�(֏ԍ��,8=ڹ9�t���Ѻ�/���.����D�ڸ�i�8�ۮ56�M��@�ffǎA+Vfp�D�ﶵ�@��;�f�$�	�X�͆��`��:ޣ��IY�����_Ax�^$���9Y�v2�v��u��ϰ�]�S�,]c��ė�!N�!�0m+����3�D�^J��֥��v��`/�ތ�J��h-���ԐD�2p���\�%[2�-}o(��ׯ�2e��B�������t���NYڃj���B<�HWGl��Qu����k#��ku��n�㎺���+�����sjh�I_rk��J�OΕ�eDJRtoA"��7[���%�赳.�c"�\u�C��o	�;[YCv���7R��d�o7W�u`La �vynA�A��j�>��p�	7r����*��:�t�z���ԠN#:-s�����[n��]}�W������N,l1�Wp(T�=1�ZF�ɮ�������V%��X!��X&=�&-
�:��+3'
��h��4R%���֪4�:(bp����Q�@�un����TPS�V���݅{D8ɱ=�2r�b���ݣ���m��-��slf��'�:�n ���ŧ��F��0�dCC���&82�)��yw�b璯s�;�=i�=��]�L��ʜh���q�ը.��#G_0N��T�җu��(AAQ[װ��S�,�����As��O-�k9X ���Ed"�vv�@z��#��;���s2�eZ�NG<����G�em��3ƍ��KV�ezp�z���vȷ��8��N
u�d�������\�ڎ�v�)�b�gud�v۸���qGSc���[uyXH��Ŗ���f�۝sX������[�m�J*Xw'gW��Ã.1N�j�-�]�Q�	�t�b�H0�v��v��Y�/!t�mvlYv,t�`c�m�y�ܼ�+vƚp5�D���;5��v!���lܥy1Y���ι��fX�p> Ƭ���C5c��6�*iCGf5�.+.,���c*ݫE����`��Sh�է��7�\\mͣ�v}v�K-�Ķ�-`�n�C UX��TusF��h�os�n����������h{�s+s��d�\
������L`�.}�\�	
9D�H4˦��uk���j��7DS�r�`����N׭[�q��Ŭ�����$nX0g ��-����Gc�,��َ��0U����W���4&S�۶æ�oC�����EH�D:�2�byw�s�!��7�̀�ݯ�-��E�^��CU����{i��-��Luu��h�6�c�G-�\���;�^�n�(��F�Ź덷s1��ln�Tq���j\s�����<w6�=]�q�������Q���^�7g����j�e�ڕ}����WX�ݫS!��v{p���k��x��q"s�UF٫>�za<˶.��ٙ�v#	�%dΚ�]	���ێ�.xCy�Yb�fyԝ�xCS��Z�m�1�^��ǲ.�yٻ�$�`�ـ�h�z��ke�R;m��V�pk�e�աc�v{v��[p��61;O*K΀P�e%�-��[/�¬#m�K��u�������@�*�-jKi�T.7���;�u��v�Ѻ^e�s`��S�'��f����뀪�\��$-��J�f��]�n�\:���Aë� ��מ�����nű6�F��<	%f�r��yٮ^w(���^Y�������FMI��f�D�q�6ږ��;u��N��77����Y۵`2��;��D+��'����s/Q�m���]˛���l�_ob�Wf�Z��]�{2=SD�;��׵�q�Π	ކ��qc��n�������:5lMq�b�ky:解�Ok�\�n�c=7 O!��kt�`���,�ړ��q�ܪs�x�y���;y'�o	v��Ϣ�Ӌ��hnֶ
l��2���&u��dݛ9��CgLM�؎�Y�nĶ�OlΎ.��kg�ăɠ�ap�$?P���_�\ߘ⮔V��;���:@���ׂ�{U	�s�a�
�����u�z<ml#�;����hn�!�; t�lⱹ�\?yWN�P~�D��<���R�q�G5n�Ξ����gx���拡�1������!�֚	c��f��^x��t�!����{��:����D�a",�۟|�@�;8���=ٌL��^��:{���sxs�|�N�$�-��@<T��g�u�f����t;��48�C�?��WB�k�jZ���8�;�4>�M#߹�᠊,�4��E������>4}�r����CA�ؾ�":�#��\5�!�6`��W[�#C���"��!Dt�b�d`��o>WCMj�Y���X��^Y�,�׷���}ސ<y����i��T����-��Ͱ�0��F�i�E�xp��p�㹜�� ��L�h",�|2i{�?v���.�⠚�jÆ��g��FP�A����D�L��6�>��n!�ȳ@������u����uV7N����nݸ,����e��X/Tn�l\tܧWt����1TnX;bY����=����3X` B���z/�ho��f��7^"j�h�]6hY�6�����l���~��T>;h�s�f���;��H���4H�T-���8P28o�5|�c<��4���~��.��"<��x8;��Æ{��y"��QQ7�x[�7�%�ܴ()��Cr���`T����)�۫��04���v�՗���4�����;<�i>~ |h2��}����:�-b� Y� Ϸ����6s�2�����zl.�������ސ:B4������}���P鬈CBd�{��Ff���@�0�o��t9��5|��Kh?C.�i��i�4]4��ɯ49�{��,֐�z׏ư՟��G6.>"8�e(1��,��Z�A���#�=�����B��p^�4��B��6�{��ׯ���E�4,�ws����.�oJ��^����3�h_%���4V@���}]�j�a+5�,�ǝ=���<&;�/�V@��{xn��x�-�i#��?/�}�ns��?a�f��CBA"�w�c�0E���B�5��o��#�Ȅ�b�-5�����3p���g�6���뇬�N՝xq��r�4�ɻ��(퓞�Y�cN.%�kiFV����SCb��@#�ϰ`f���:�T4N�P�0����t8�C��͐��_wy�<�s�|`���/w��,�Z�Xl����aj�5=�,���z�aE1	R��S�b�5�2'�K��&����x�:>��¾|h���f���Eڣ����᠍h"����cxA��!Q]W ������V��;���>�5ޡwt�;L �&DXh���ZC4� !i�}�t4��G�*���U�q]j��wݾ<ٿ��g3�$�^�R��x����q�N�<tg6IЮ�pU޶zf�.��گM���t�V\�C��A�L㞩��/�k��j�f_�u�{�!����8k��<lC_qP�n��#M8�Ng������2D�CMzA�+-͊JB�7��]Pl�yZ����~���B�{�@ľ=5f�Y�*Ggٚl|�hC���p���t�T�Z��h>�{���4>��#ӟ{�Iu�d��܈� �:_U/��Br0	�f�r�ſAÆ�s]G9/w��U�o���G�iG�C�_}�pX6ۡ�@Y�^�=49>Ϻ0"O�pІ�j���5��0�8�"x=����	��y�݅������qe�tR1E�f"-n�tci��ma6��������$��C�T�P��O���Xt��:�B�"	�ٿ`�nܠ�x����?_�D4�ڕK���l�y����,}���~5�U骴���_�X�[<4.'-г��V����
��!5^�;�����;�|�~�CHw��<=�T5�O*��Y�훡�*��Gث���C��/��j��:��3�c䫄;��Ɨ$��������|``��8�bGQ#OA�}�K�@@������CL� �r�H����^�:a�N����7����Ƕ�!����xh3���,гA��a�4�125�Y�=�|�*�pBZmÀ3���zG�h���mT��	���h�Gy�VhO��H�C>�p���׈f�<V��%��`t��ԍ��Hݶfr�X��5�`�6}׆���gX�5�Y0I}�q�`�׼��wVC�c8%�T��۳�c܇�������C�GBf�4�l��(��p�[� �����$������!�E������i{��# �,:xD�>U���t<�3Z/�Y���v�V��A"�5%����pX������0|kH�@�|���i�>�'
R'H�B���6�yv��T�Z�s���=n۪�A�ֻ8ͭ7`ѻmR�H��Jt�H�>�۞����_�C@�2k��5��/�(rw����D�Og��ߧ�/����i��1�49{�y`��f�5�����a�P(���pe�khY�5g�k�\�Gfw����ok�p�A���U��t0���_a�ΐ;=�;�xh3Ǭh@hw>��0+U�������gvNP�D2<k��0N�&��`�������tb��kO�0�Ծ��=�Ct4��d~�t,��tp縮�E��Դ߬��|h38�S7]���x�a�@B��we��C�5şN1���:s�2QV�$�܍)"� i��pC�36�#�<[�E�ʝ�����#�!g�t,�B�O��`x�*�F�:E���\�'˦�E��M^ 8�X:>쵏��k�syΛj�h�5dx�� 3��X�a>ӄ�	��#� p�f��~@Y����u�i�Ȩg�;u�i=�[��+�s�`#��8��c0���t�g`L� om٠��cMi����CZC436��5�')wy.1�1��7���t���}H���kiqj���6'F��B�n�B�L�d�J[�7���"C��]�f�`��:������sF�y�g[]W-U�v�8���흠Y�m�!v�牤,*�S4��s!R�w;m��]tF�`b�<;�⫦��ɬ��3���|��|�M��F��,��P�oa�E�u`�E�b��y맳�KF�;�Y�<��\�:��R����#eq6�ctK1e�XC1E�/4Z�c��Sڛt2�v;)�P;��0��y���^�]���X�v,���Э��k`�rf��ud(�E����&Q3Ք9���|�,�ކ>�CM@��sE�kx��~���;��^y���sq:�!��E� B	���z�f���щ�׈����/w�3C��c�t֚�d@��w�H�
@ԉ�-�t0�����g���:�� .#����;�D�%s��P�*��W��ݿ���\4=#�,Ї��/�.�zzhB���xA5���v'ʴпdμ�������p��9���Si9J�)ŔlB<l����������G5p�4,�D8���|��zA�_G��^�A�6j.{��v�І;`",�$�@��ߍ�ڭ��@m�4ȄC[~G�&��!	l�AR���X����gVd�#yދ5�!ٜ���E�}�.�#�������D�9���߾VEt�g�D�/��w�����k�z���4���I�\|A�SM8���+�p���� Y�@Y<��K��a4���!g>O�x�nsք����p�g�5al�T,�"}�p֑
��@_>�To�wCګ�j�۸0����y�_��7��&G	9v��]�Y�g���vu�5�:�c@��	J��fF����J99C��4<��d	���t4�����B"��Gs�.|n�uY�C��\L�����}�`w+>�ſt}|��|�2- BL"�U��]4���ư� ��[=�����P&aH�XǦ�s�a�f�C }k��1��;5�ǿ*��<B��	ǗR��)�N2����Yzf5On�RU�Db��"1���Y5[Z*Tإ��N�c)�zXЎ����*������>!��g`/�,KMY�0�_|�����4;؆�_Z��m4�|��89! �ޡ�������Q�'���vO	?C>w|pt�i���"��}%���h�Z��yӽh#�o�������^4,��`wt�4.}λ2��hB!�k��h}�}�`-�$!R�Xy��߂hw�x}��c�t�@�ջ��ih� C��h�x�5k�3C����3ִ��ψ�|�W��>�4ٮ�C_3]�j�׈�T!�C47�;��Wk��mV����w���+<: H�Yӟ}������t���#wA�߹5�+��㾚�ުk�hCA��v4�w�Ɔ������ˆ����f��ȫ�CS�=�����}�����*��1%tXƫ��wX��1�m��rj\)���h�isf��]���4��.��"�ߑ��p�@�f�#�K=ϝ��>#�Uf�ڡqyB7>廭#��!��n�n�{�`O8>�nt�k��4�ÜC�a���῏mW��C^�Z<��@CrH�q��]">0��!�o�^���/}��y�f���B�WH�[U3��c�NqгA�f�����xhr*�mP�}���n*��i癿�"=���0�R�/���M���PD���D�i�ȳP�#aW��t:zk��B	��`��G�U�N�{������b�OE�kp=h�W�A�� F�Z��� �UѸ7��;d
���*!B�w*�8ܳ��&V�&�꾕dm���TW*��Ua�X:]RL!��f�a��Pg�1�������!aG!$Zrm�!��������ON��H����v�a�� ^��v@�}�9��WC�*�l!v�Y�{ �s���Κz��;�7�����x}�AM�v`�U�A(�#^!��ٕ�0�b99t4�> �B 2֒��W�H���F�T!�!��w�����&��Q{�`���ր���`a��o�4!�����4�405A�`�GƧg~{I����/���hl�eeL�&�sj�UQ�*�v�OX���Y4�f�응9���I
���RG��8k��YN�6�#���~7�#�<lІ�(�ҿ��t ��CBڠ�H�߶���l�j48z@g�^�M2/���5��>��7 ��U�hg3�k!�҄l�Q@d�hp���hY��Y�|��"���b���=��&�L:k���W9%� D#Uf�;�H���C�$Vh_o�#Vhw�x'"3~��j�>I��?< �3�%�d��[��!�koO �C�W������]4�� :1a�ߍо*��m���mA�p��OyJ�>�</m �g���-|�%�i�"5_ы4s�#)�r�q�,|kH�>����������4[�����Nq�"��hwt�|X4���n��]i���>���2X-5dY������߾�3y�~׆2�&n>��tb�.[Ox��c����'�u��ƥ��QG�[�|�ώ��*Bmx��'�]�
�*<���(�p�k�3A{���L�!L6��hq�	���}��n�$�hk��4�#��1��n�G3�e�ˡ��<~#
"�Zc43�_�X���� {U��H���	�t��*��
$ա�8���W&��è��(54O�\ۨ`��Z�[��ڧ��54uv$�-n�i�2��l������߇G� ��G����#�*���̔,��K����񀍚�D١~Lһ���#���︰w����謇�a�a�j�}�t8h���b� ��~yq���ArK㦃4?|őd����Ų��������W:xzhx�Ds�a���D_i�GY�#=>�9� #!�C��lm����"��zl�@��,�����
k�BeC����C4ѨF��|�������w4���n�{<n�sò�FLs��4y�řlf�����k"�@���<��<4�A�#�!���.��5��!�Q)�Y�φ����b�/�a'Z�勡�,
���hy��wB��B���5ds��+��uг� r_ÉL���<�W�C5�����bP�Lψڽ��0�R8]&��ǀ{���4�\9b�������ae��B�F��Zߧz��>t�|G8��}�hCC3/�(i��D#�Vhr{�2�� Y1Pf���>qw���3���n5�8O�:F��YsR�CD͙�֞�O��.���͡���h���u2�ز�(�8W+o����{v.m�KshM�g�h|7gt��uZ;ux��e��X展α����D��SsUf��Te���KW��eܵ���q�=������\:7I;��/k��p�0HLF<���[٫ktm�6f�t�D1�Z�1)M2�t���,�}Wg.+���r���\�4�\f�&9�vo�l�Q3�1�qQ�f�t��mu҇G �yܚ:m�e�Eі��V���e�D�4�>͸�����s�q�;Mnڒ�0q5���l	�QD�\hW�'Zگ���rx3|��	~�~6�5��,І�#����>w�]"�H�g}}�`s���z�xyh4!���i�x�p��K�F͐!�"��q��	HHH@�"Gx�D#��i�����$ٚ���x �<�������T!�w�ߖP��xY�!�|�㹿uXW&�dkO�5���X�!�<j�}Ω���ur�EP�h.��At">�4���c�+�8i�q�� }������p�4>\�A�b	{�wC�p:��3��ύ�æ�>5��������g�`Y�f���|�CZh�A��^�Hd-��b�n+��p�4,����߯@�>"n>��r�p�q�49j�#��{�h��`>6F�VG���0���@�������n�a��3H�k�r��܈�j$���juh?�����k��x.��hv!�x�}�d�'��-7���m��5g� Y����XOCMP�G��k�+M�o��<u��#�xvP�W��<����,Y�<�-Q�d�t�Mq60����g8e��ɮN�{uU��u�c:@�T`2%�;Cs���g�݀2&������������dwC��A�:a�P����܈����oY���^0�9��{���V��vi�f������r4j 䀳[C����#�����0����D���&G�[��&�i�z��ʂ�;��k7ßjj�<�i�=m�/�k��Bn�����4�zֽ7+E\H3���4�d]��y��Mgl��#B�{�h��h"hO{����%{�,��P�\h]$�s��P6e �
&p��_8lЄ3�B�,���`t���VhCdQ�Du����6�T�p�D�o�a�%���櫬7�4,�e�G��43>�]��i��T���h_�lkq��&�%$�k|�֨Y�~�|��2��@d��oE�\��op��Cw]Fڬ�O+��Uh#A}��/=4>�@B=��zyo������},2,��U�шCP�����\�Ja���gMaи�2�{���3Ī���E�陧�����W�'����Ƅ6D�hC��U������3�B5fko���>8&!��BύCs~cNuW:��V���������x��]��]jbh��iAm(шg-ռ�ss�b����v�W��$I$���8j�HY�"�_�3dG�L8G�͝#��4�i��F}��t*���@�a���ٰ>�).o���~ C�P@��gH���kMEB⯈���ϵ���	�Rr<��VC t�A��嫞�%���gݏ�_+���\"���w9�v	�ȇ��=]N�}������= e��MXW'��}�0�ʅ�=�|H߾��<h#A�8A�5P�-9.�!꯾Cg�N���<��j�iՐM�0�:G��,<�~r����y잵���v؋�����u��p
�T�+6�ʗ��8vtN۶���,Fm��t(���Sʄ8�W:�trX�~�{[L�l��2��ƻ=�c�7�Z���*�7��xI:m���CE�1���L�z��}��˳x4}�ۂ��$�r����$;�w�Z�2��`�Y䯬����2v��87������aI�\;�����MbޜѹEk���7���I�	�n5. �ֳS�q�5B�T��7������7;%�,�Ku��`H��I����j���7v+2��&�~��J��϶�w�&�#�4�\�0q�Ns�[)YS���FȬ�d�;��n��}Q�\^'����(���b`�W�-oh�*�2]�Z3^�*(]p�+�z�	�iK��pix�|h��^�+�H�M�8fW��z���p�v������O:Y���}��
'v�G�8��ЏgE$9��Q��8�0�=U���(Ǡ�&�FB%��^�)�� ?����=�j�}Ds��x���XtszC��m��)�.#E�v��M�d��[��ל�97�֭��J�SE�Z:!������[gJxrX�Ђl�@��1�$�$z�j��B)ۍug$#R2v�^wr�$����P!9�}ٜ/�K�pG�2>Իy.�j�ؽ�j�K~�`Z�'�{!�1�o��	�&V�i�u6�1�T,,���4y+1��ǲ��_2�E�'B���{HJ���e�ݖ[���3צ������i�0�Ӧ������ZB3��@Y+ь#Mw��x��mBC�� )�t�'ƷP�Cm1����O��y��P���Λt!,1��}ώPބ8jD3��}�e��A���_w���ϲg�����c�V�>=��@Y���/y}��ò]��������)쒒\����i�B!�g+e"_��W3����*�����ϐ="�ل���`X8t��#M������ڬr*�BYS�0�4��*D}�8sr���p�?=�,���LGDKt��찢֖�Y�����[Rݣ.�f��2�73�͐�8k��<�	���c�e���}dݳ?�����ME@=-W�z۠^M�V��O�Ofk���AR��l�@6����ף�z���=�3x]��3a�y���b��x�o]o��BА��[�VL�@{O	���@� $3	!��5��k�'�b����P���]������x��`�:�\/��$�����`� YP)D#�I�s��޸��~�}�1b�ԋ�#��W�Q�s׾�U�͎qΟi�ˬ�qM<���h��_+�M��y�qM���E	�;iή��Ýӭ�3Gc�1a��23)�(��P;������d�X���(�E��!�ذ4�=��Z�k\^���+ҧ�����w������{Ղ_cH��h�q/���O��Qsz��Q�n�M��C���n3���N��w#k�R�Pl���O<�|�qk����9��I2�{��D"p���HH��,���g�]�c̫P�y��f�~��"*�d��)A4��:;��٩�J�Ct�j����Pʎmx"�F�
>~� s��=�Ǫ֭~��P��h�X�)��v/W�Υ{wת�0&��
�6t�;=�وv��5v�,zy��WB	ٜ1Y����$Mt�4Bi�`9����Ǖ����?_i�jB�캿�Y���N '��g�����[�M�ٞ壣*Q8�1��Q�x@��d�g����Cޔң�j����؎�Y}��^�&g�������v>���n{�����cP|v�(ZsXE�	k�!�����R�}%c�����-7��6�Oz(��=��r�,��\Q��OnLm�!�F/^�w��h���v��A��֋��D�+�c��e��Z�ݮ�z��U���Up��@���हW����5����s���u̬�V�15�+,"��n��2^�v�]��H��f�132�Zm�;�ۜ-�Y��U��v��Q��:���o��WbN�Rx�q��vC���v Ϸ=M�9�o^�E���%�[*$E�LGܺ��[�zz5�e
-�#'m���rՄf�������m��J�����4ȣ�e���Z\a��%G
H>�����}�{5#�Ϗ��L9��0#yry{l��PX��h-�W��؜oE��7B�a�I�Ld��h:>�㚅�����b1���e��Z��]��f�����o���yL�sƷ���-U�a��Ma')_�l����4�;9��g�8��e�ɨI/Q�jm�Y!�*y�s��x�4��L2�e�4�o�n����^�(T���Wl��|�~˵�� ?,d���� �v�8];]������w��y6�0Re��Ld�!mwK���Ǝ�Y��?Z������h�Nȱ-o����$ǋ0:�N8����u���u����m�{t��m�q'9�mz�v��k��G��̶V�u}D�<����=�=�'�G�{�NwB��oC�>Ӊ3}�6�<<Z4y+9����\�a�0*i$um������s�^�K^���=�"˼{v �-����b��t��{��h�H��8�ѩ�qQ�}�IX�u���w��X)ô[ɢ.���:]z�L�jV/�'�����,Ã�ʛ>�/2�ٰ��m'��aZ]x�ASt�)����2x�V.[��}�A�c��7>���g];:q%������3�T)0�H�E��x�g�O�.4w�<�ͫV�"����%��|�yݓ"l!�_�}�6�Q�O��g�� U��w����l�d���q,���o�q���Z1��rM�ܔ�3�/G�=�u�m�=8J�M���v����'|�h%c�)Nx��Po=d������.k�㛞�a�j�����)V�qu�����J�����2TH���l��u�z�GU�{;�g��N��Ot{��],Yc��ZM��.�j��KMJ��{f��sChe���w���_��)�s�jm�{T�����Kڮ�2���<�⏙	P`�E$�p�I���x���U�k�}�=AX�{v�$i\.��r�&��D�(F�f����wDmrB��;y�E�O�������&�����N��,�f������VG��v�[�N>~�NV��=Y��E���MK���`��3���4287x�
{���1��my�nS��#Qu���7�ʓՈ����O�SU۶���W�x	�M�S�9�뫼��M�����!�j���t�&)���ue�g��-��_aݿf��ӎ�8h/��� U�]�;���������*�ǚ��f��/gB�6\d��L�4d�TRI�u��a\���(A�����r��gxx�EA�WzF����d6��[�j�-*4U:-��-:��sd�>����4����%�-�#���e^v�JrL�Ľ����dv�
�T�l�b�i�S�������J�Y���fb%��Jɘf�g�˥�3ζ*�8�c��u���g�o�J�4t	���F��g��1x#�wd�m����� �X��
�4ߊ\�ihL�P�e�nޞ&�V_�~�H�r����%-g^���7#�B���*-��]
Z����͕��S.�kԥk��=�wu\�����wa�4I���M�i��*&�w������/�C��W�Q�]M���Ww�1ӹ��d�o�%/y�oObTWP@6�幗�j϶��n����g��Ҷz��v ��^.���s�s�#ܹ��7OicW}�ߟ���)��W��^�'K�$��3�ף��G��u�9z1ޖ�0���9�Qj�4 i�`(��pr�}6�n�X�߳C��Ąp�'�$X���Ѻ�ʕ��>���]�{�RA.��s����@Q@�'	��ÈF�*jBޒ����u�S؁o���y���W�g���\z�$RF�	�$�}��h�<���ɮ�ka
������μO0��� �][�}�u���˥:RGa�3�(M��N
�F���d܇f$����oz��r+zz��3�Ɏ�ǟY/�^" ���+� �rSX�P8�5GެZVa�i����u�3]�)pxe�N+�<z��xٶN�����AZn�l��{X��> �W�svi`©lJ�T4ܾu���۟<�m�/V�{twE�%��:��,R\�;Y-ɜ$�In/0[�3�A��n��Yu����ω����kt�s6�΀����a:��-�Q͢�a-�Krv0�u��r
W=�+7���&�w������5nn��{Z�Փ�r�Ci��c��c�,�h1��׀ �=��K��ћ���G1�av����차�bR�o,b���Kk�Bk[�vnx�v̳ct�N�{u��'D_�Z�,��s�8&�ǀ����O'��`�z
��9�
��g�
���0�����i$��z�m��������O�4nv�����@����*���W���z�~�%Z\m�9��g$��l�M�1,hrz��Ύ��z��v �bf�ɞ�$�ۂ�<��c*\���Q��D��pdӻ�Op�֏9�>�7J���{��]z-Ǔ�*��b{gW�z���g��[�43�'��h��c��#
�Q���h�I�~��{E։z��bT��7k���������|��G���^ܼ�<3�B=:x�d�;cQ�,l5�ف�4�.����I��E������W��U�Lː�w��[����3��jr�c��y�2���׊���ֻ���iY��	:��鷫#Ֆ� �Z��z�h���8v1}`na,]��L�B�t��tν�Q�xzj���J�E�c�j�u�e���>��.�S�&��+�(�&���[��7�˥|����{9ۺ��K��K$d���*m�'Eٷ�x�G{���$�KВ���|v;��yg�h�NׁbĞ��O,�CU�"�K�(P
�MT%�~�g�f�s�W������5gΧ+�Y�K�sp�̄f�b�"��y6��>����[�YN����/��7ڐ�tZ�����Xoi]��~l�z������z!s���n�J����K�N01l�=���lfQ(ح�O�OF����B���*8���:�b�a�
��9I�Qɓޑ\���`Z�r!F}���%��י���}�Kwբ�dG؞��-\�h�E:uM�4��W$�5�U�^�����x�\��[S���roj���]�_
Qi���s��D�o׷=i�Gn���7A�6پ����pX�%�8�ssDJ�P���]�|�:ھq�gC,�K&�/j���p�u��GtU�ΣV���}���`��E <0�]�O[Hɨ��Z0;&���"=+o+Zb���W�8z�K^�ݞ�H�Qv,��k�Ý F�wϩ�2z�O{=<5�K7³�O&�S>SGL@�T==�`Q����ez�y����4���l��m|��l{�j���Lq����z�l��y*H������[�t^-vRM+����M�i����n{k�"i ���xy��-�sW!�s�qd$[E��B���$�m�{���/g�7�H��}��\�n�'~��
�l�	�?g�6�W8W��.�:�^�9E9z�G��=�3Y�bˇ���\�k���)�/}�-��by˽)9�x��:-隘:�����X�:7`�a$�h��e�n�5�U��n�	���5��ҥ,"�uݘ���pf5�>.�3}��A��5�pޱC�Qu�&b!�X�W���}A�<���}�=Y��紋�DZuO=;�)1���_�¼F*�;�73{;�"G�[�����ɬ���t^Ğ!{����d����]a%����jRG4�������X�N�o��X�����ugW+N���ɕ@��(�1�9
uϽ�җ��4�3U˫k�s;����哫/�u�&A��}�=�Ϻ3ȏj���ƌe�d�R����]��b�4�����c.z����u=��{]\�	��M�7����u�jӷ�-=�Ɲ�륻�cW�!�h�LƎ�U˙�]��T��y�h4Z- ���^�6�F�e�{͏)�3V�w�/��:8�=���l��&m���>��=��rg,�չR��j�)��C�]&����o�=���W��hy����
����>9jN�2+NTt��V[؝sm�D�`��B�	��e'��;�|yn`�9�x������r{�RLD]������V�g/_V��ކ��>H4RH�����.�w?]:J�=9:GE�p�.�vl��+����	��u�g�uUP�x2�7(�(\�6g�$� ]� (K%�(��]3&��� 'F@�����ZUe�pFd�u���i+A�����B2�=}�b�2�gr��M�Q�-�a߲Z,��;g`@m��_vB��\gl���7i;@�Aa�Y��[�*,P,f��}�i����C;HT� R�+�S
�$��(r��l	r��2lޝ�k{��3���x���p�/K�d�w��kYZ6[��j���-�%;�0њ��;��h>��Z�)k��#�%ū)t�����ս�Iu�]H�d^"����l��׻����4�@�c�c]7���I��� O9iH�1y�{�d@9�jрkc��e�t��������{gR,��n�ń!��p�X)�o��!��M��u̫ΰJ
��<4qi�57'cGW$�3.��6�f��桔g#&��-���:��hr�y����COAX��&$�t�5�*�����N�Y�ɽ�ݕ��9"��9dIAM,�>���--P�;�&<{����]��Lɵ{4�-��_�|9k�A�a�D���f�5�eQ�lv��3�C:�,'8��%����$`�6�qC���V�G���N�^ �׃&���۹���������aMv��_f�G�yWPd��ԗV��!�e%WDE�B��{p�$������F�h�f��R�����+Bb7���x��c�hd�7c6a6��>�V÷��c����h4S�H-6~!�H%���A�a�l���1���n���Y��ӈ��XWv���T"u��[�4,�-q����8���n�;u.����^c:N�.\g��o-�Y^M�R7EX�6Ū����0���i���S.��"0�ia�Ê8HGF�aлg��:��M3���9�q�}T��L.���V7	c�[S����kn������q�r3�<���Z}@��re�Sv�dVp��\1\X�9�Ir����3�r��O;�O����]g0�͘r`U'{i�k��v\BH�[��˒�����g\�� ��q��y�|FwQ��P�҇t��dqj�<��Z����AᎥr��ÂoJ�ūy�k�����u1<�zݼ&���z��m�#ü�y1u�Y���+�ʺ���9T�2��e���
��|��xX�#s�yݢ�c>C�����i$��f�8��6�;;����^��;;5���.�p<�]�%���#�Fe�e����N-�k.T�z�a�3��6�z�cF�ַ`�:�h��\%�ύQs���K�W"M�χ�8;RϭF+�h��P4w]e��-*y.�&;n{5x�t�޶�ZðZG�vt�y�v�i%�%]p��
ha5c4[-�:%95�mHԄc����@1�.�
��ۭ�����:��y�k>zZ�c�,Iie��n#��2�ld�i��Dgb%��t=�7n���̊�c�����V�K���;s���h�[�:͹"S%!ŕ�-k]m�:r.u�9<�Yr�Q�p����ʨ�l�ui^�Vr;аr��B�y�ȼ�|Ҹ��m���vѶ��g�%�r;��TJ�ݍ,-El����4��ݫ���{d�;
n��Ǜ�ɹ�=�82,��6ں��ޗ�s�8Ձ��է�1�%2�A���"��B�f�q۵�d�e��-ę���%vC�s�5VXń�s6���f�3m�Z��4���fq-bʳYs��sLV=]�_.�<v��y� w4���a%�19����{��ke��n-ңś]��[�qk����m��ٍ
Zc��t֬03(���^0s��cv���t;�hΠu9b�&u����|���چ��&bצ�.��,6��V�W'��%X5��t��b,�\�,E]��\6���{pp�؁y�h�,,�@��c<��>q�:���4ֻh�1���u�m����X��^�l8���G-q]��vӛ�`p왆�>��mI��'�x@u���v�	r�??'�R{�����|efn���y��~h��D]K!Y:ta�uþ�*�v���2��tm׽֘z������Ov�d��ժ{�w��L����6{�Pfu�'ʺ��^�t��Y�2�k͌�O�m�z���\!(Ti��8r7ӻ�s��.��v����}�0!���ݎͯN뮛��5����Y
TC����p����yp��9u�{����oO�5�e��9�v#Ꭾ
�x��V3��>2�6��w��$�
�N����1��\�k^��=�!�1�NB��e�zʯP��e���2u���N���zŎ�<�f�*~<ҧ�|�O'�3na5��l�c3L\�L�YB=tmʼS0���L�m�����]f��:�q$$�o:�#��OeOy]&�.�Yy�¢pR��޴��\K��P���~nJ�5յ��i�m�E�����Wr�w�OV!��Y͞ӵ�e ���^�`�"�����V���f�������֫t��-��z��N|����u(;#��@v1�7H��5���)����q�N�ܬ���Ggu�Q�*�]zbr�<	K���4.�1�Rc�J��gQ��gԯ.p��~�7��{r��ū�ւV
g�o��')'�����@�d6�ZH��==����V�w��{�W3ή �{0��k�L[�C���C�Aۓ~�ۖ7;|j�C�)Ӣ�MJ�$�&or�o��	t}��5ґ�w[�Ӷ���$B��=/�
ӪU���i=�__S���F6�x���xI[��^:t����nq�9l��s>�*��V�y�z�[�i:�$��=��b��̲�.�W`���|7��U?z(K����]Z�%���u��_2 TE�.�N���DW�sO�ͮ^�o�sX���l�BL��x=�gOgY�o2�@hny��2M$�i2�b�ʋ�{us���:�]t=^�m)^=��<֒=}�rZ��f��]�F��jI{9��C3���JI-xm8hY�~
3�$�6��[&pVM�Bfk|�a�ٺ2m��G%��v`��kWx�[� ��)��p�s�+^���X���^z�{�0��_P �� 鯓A��7�>{�珝�tz�t�۹�'V�I�]��e���4���R�v��<&o��9�fuぢ�A!	Ro�į���|������;��]k���ީ1�o?��9�<��>&�+���>�����'�e���)̭��@�-�=t-;�oG'f�K��Kr\������N*o���j��r�T���ݭ���5Vb��tVmnC�8�-q\�(���$i�٠_��SY�'��4��h�R�ᾩ\kz��s޹U�֒�|<��"ϻś��ݡ��{x��y�x�C���#-Hh�&�u�;���:�ɔ0�����]/�¦u�[���I��ן��oD2D��� ���Il0i4ۭ�����j�{n38��%���}֜�F,z��=����{�����F�jy[��`��j��-�Uҧk45��;�f�>Q����I+NB�}����,�Qn�����iJ��ޮ׎�>F��ĺ�9Y�������L�N�(��⼎*��	��t��
����h�Bo���M���,R�Sڧ6f�5v:�G�Q]�ub����:�*�sjl뜷d���ّy���N�=�uU\z*�v4�����F�$���`���'w̃0ݩx7/��'��㫇�����s}[W�K&�3�)���{779�0�M�@���:"���o�c[��-H���#&��7m�l���q�z�/=�	�ϑ�;��j��\������k�a�I�m2�i�ˤ�������-�,�>*�3��g1I��\������Vm��p��2�D�`��H�Rj�6�-���O��z,���Ly-��3���/pL^�*iWMX`@,�O�y�;F�|a�}��,��&	���k�vN��ۯ<�8�Œ��W���u7��3�+�$u��������J�ſ5I��yY7j��9l�ڼ�ۭ&�� T^q�W��`���d�w�WZ�޾_e�eu�c�r��OrS�C�5+X]�dq]�'0Y%�<5)rdσd�>�x9�I"]�E�s��x5�v�fzy�PM��]���nJ�U��f�*3U	Q�ӹ��x���{I���Դ��r�ͳ�Nv���[v�jQ.wnڊ�mh����϶��:u�=�P���emQ�����B��=N2��Sf.��ME��-�5�7b�k�oh^��kt���;8{5v
.ί>�{����6����3ύWD�O[A�IIݶ�f�1u��S��l�Xm/�|����WK���������*|�<��p	OK'wz`]\��W˗�f��MMڶ��uΕz��M�h۬���s}��=�^luq�zH��.$�م�L�^۔����՛\��{�"�B�L�i����#zFn��ȥZ�{ȹ��)fVW�ܔ|�xs����}/�ԫ�Nw�$��M�!H����w���[y�!�To�.�}�5�h�e / ��;�-A�%���~5�Վ�gL�J
�zR�Y�2A�!�р�	8�R�bu�W��;
�w�J��
��r��L�/�v�M&;�s�tG��B��e�0���Uv�E�R5t�,sm�b�r�;uR�i�	�ɖ�+��P�G9fz��8�����ާ���>^c�N��j�F��pX�z�@/m�S��m��Y�&L��I��XR	�à�?2��m�����Ŋ�V]�q��oZ7n�p�J�>����P��U-���WirL�� �N�Z��w[��塕�ݮ2���\齆I���o�����b����w��9T\�Z���z
��{-P�~�m�G����Vz���b"L!���&2y03��qޔkZ�d�}ݕ+(Uh����~�z���]ٝ���e��sǤ�01�PB��{�(�$�(��A�����#���9>u�kc�:���@�A-�S��&�(|��ܾ�u��lq珙�~U����L�p�o�=�P �� �7���*al�s�;m|� �Ѵ}��Ψ&�[S7'�#K^v(�Rh��7�|.Yv�N���ܶT�L�;G����"�_52/��띞-��k��3���B�����.�k�4L�ڮ������|ǽ��� Fg�㾁�3�&��nu����S�Y�>DU����Vī����B��� "�[6F�D�Pt��G쇧����sʋy�C��`K�,�?o��'K�B���)�CN���^�z�N,��,6�D8��3ˇ��
 ���IK}[v�����*�2�i,��rU�n���泀�|޾�71���I+���Z�:>d��t����Sa-��LS�����!�d�(Xdup��n�x�qL�!�oy�oy���t��ל���h"��M^$�t�囥�aݩ�R��ثhu�ݕ�y����y��^�nnU��BϞOf�|7�OW#Ym���-\8M�P���Ȝ63-�5q���rWHf��3�$������M��3I�d���}Ժ����Q��b�j�x"�{���e1H�"���;�:��N�U�My64S��kS�����Ze0�)�E:I:�2�y�_q���^L�����
����{�>eض=,f�����U�Z�8WQ�@�7@��օ`!�8�_�l�o��Hr�,�.��iµ�����|5�������Oc��{Sg�t��k}�^"�i�!�n�����[wַ�$��^h��~��{gt���W�wU9:��3	i�۽�C`��I�vf:��z�e�o����uy���Y;�{{ԡ��*n�1I�FT�e!KD�|52��� �q{^���[�Vr���$��-D�7�ִ�LרE8&� Z'_b�%���GJ ���:	u��&��9��~/ơ�}޻���zY1�)����������29O��E��K����]��������*a�oe��r^K}���Q�(���j�1ܭ� �� EQ-`y������˔�]�h��kz��霮�)t��r�2@�.I$�
b$�缜[��c�39�2�	N�J�����>�����GO=��G{��W\���t�ָ��{�\�N���#,D"��#RŴ�$�_3,f�*ˇը�q���/w)[����>���y6��z�q9Zg���K����������2T������/)���]eҤ�	����L���a�+�'ۤ��Y���p4�&)������B�ƶ�P�f�+�
)�SR�^4{�>�f�C���R���X��u�t�,����e���m
�\��>��=~^�V�[T�vט$�(�RFۆ��d=bn�;�)��v`�I[�@�ه=3�a?Q
�!�:�}���J\��(�s��2?U�iM�z�X���خ���s�<`�2�� qe<V�h��DR�X_�v����W��fgΙ眷��|ֱ��yc�s������,5�,R.���&�Vŕ`:6�'F:M\er+s��<	�NP���S[g�]rJ8�.�t�����`P�p���m���̻�L��\�k3[LT�z Y���$�
�:�'R�,zh�0	n��ee�4��,b��W]1�1��	_#+4UM�k$�Y�"�����v��kp�m�/�.ʓv	��'9��ɤ˘3��2�L����îv���^,^g7�P�fVۥ�x�O��:Y�9�BM�QX:�67,p�lKe���h1A��e:�֒}�|����X����������Q������p֝{[}=P;�"�~����a���㵀��o�i�)�h�j�e1y��r�Q��G����-�'%��]��sݹ]�٤=>�!���������H�o}xH��ɀl̿*Ԋ8�(��/	��ě�8/f�ݐ�.?zi	��SQ�=L�L���;/ϥmK%�Z�}J_��Wi����,ͦ��A�M"�Nb�&�ך�b��@E6����т��U��>H��Q��ظ_HP�KE*L_������s�
L҇GX΍��$rEu���G�}x2gvK����w�������)qJ��\j��瘱�ؗ�S����W���Ց ��>���Jp�dQ�P��.��<�ȍ�C
s]Z���y����;R���v 9Δ�O�������,o�uk��Nμ�WI���o����Nx�z5���݁qb����!�g�/=&�]��T���@�um8������!���k����k�9;e�W��1�h�pu%�p��e�n�pw�`�f�,j�s�N�f�6�q�ac7;�B잫�/�D����Pַo�d����U�hh�C�����z��_2��w/��T��!��V��)�J����5x)����< Ǥq ,��Q5�p�{�/�_9�\�y�cE4��u�U�z� ��ޮj�81G��8�|�\XQ3X�Q}�W���h3L��4�=�l�؀���$��@�N(����~�DR5�s�a���n�����ޯtv�G��������Z�gmUY���&>7��x����tW3�j��� �CH�S I���?r[$�$m�Evd_�% i4:@�~�u[i��Y 3;;L�����:�ˬ:@}@#T��|�Y�:j�B���^�H�x��CM3P��>�.��{q�yA�QI��d�6�y���:	xy���^�n&�w��9�����;=NrfB�N>�b7̀a����"^ ]�X���4֑X@F�N��WP�]���a��ȡ�au�ɚn�{�����w�ǣU�8D4���dVe�w[h m��^�@���t�FB�M�
rXd���MPFK`"����E�`�w���xOQ�MV����@G��`sU ȑ@�4=�
�w�u�j��H��)��E��K��M�w7H|���t�S5C�{Lh��@�!#v+��D4�x�-
�}�;�@�5�5B*���b����A��5H.��U�}�d��h�m�� G�Q[�x��x/�U���N,
Vl���N���"�x����Q[�.�tb�1�]��i���cԉ�ڋL[�q�GB��Z6Q�B��1�����ڭD�Lff���\T�\u+� �СZ2��N�'7A���m�`1�f�ܒ$���yP�#Ԯ��p�}y[�t���h���5�Cw��0h��<|&Ή���#�s�7��K��-�.�%h]aW)P�s�m��9!��!ܘlkż���5��Dp�ɨ�����=-�t$� �.��F��ݘ0�r�[�_P/��կ�y�3�������U�JS�e�݃l�����.��gv���ь��r�R��5F�)y:�G���֌���1U�����c�I�X�Ţ�b�.3�E��=3�f}|҃/l�2��^��9͂�����+�s%]�[�~��ҢΥ�h��+E^�w���ዡ����5�I�hۦklek&���l�E��,��Ű��%��ѝ��r{+/Z�� \�l0:<�Sjx��a_��P-��ỏy�X�1^X�B0�]J��yZ�]�/�R���;X��i:�����9�F9q�y@�����"����ۄ �p��͕~2��̧��ҍ5#�Ӂ�6��|t;�m������/�vnb������|	��坎��Z�(j�f��,H�IJ~�W5гIPvV�՝b�2��&W=kwKxU��S�Ss��E��Ү*E,=��4#�� ��aڜAMc���]<�g�x� ��EI��̠���TH������R����U�2%'�n;�7�~��ٜ�5�Ik����(t�d�A�o8�c�{|�紀���_�p�LгZ:�����U���	�!�hU�[�uXEa�T2�֮��P�CMW�@x�x@^�� �{=�^�M
[��<�Ut�htІ�j�Ր(d����.S;Z۳�NI=�xN��'��0���ڪ=��.��B��B�ШER"���Xz6����t+�� ȩ�� @�y(�|�"��\45�@d@Y�4)�ߍ�]�lUt��(#T�� �j�٫��s����ؒ�8�h`��/�Xʏ>˸���q��!�%$uV]�j�]\���m�A�DrOP5�@�*����@�C�w�V!4�x� a��U��F���; V���5z��B�� s��+ 7j�v�黜 Y GA��E^�0�5C3ٲ�YX5Q"��PdR j��N��Ϊ�"O SZ��i�P��ULB��B! a�
����`�D������ "��Ua�Xl���;9�����@B ��o�f�hdN�N�� {7��)@t�)�(#L��V@�C�s��Y0��9�/���� i�C�@��@�����f�JP��c��p� i 3UA�ZES5@N��/H�@��+X �H�T WGE�� @����Ej���,`�@�UXzQ5^�Λ�H�,�Zh
�UtІ�;��!��|�f��B� Un"'tk~�C���&GP��B�MP�P�T,���:�[�8E�5睊���5@"(�L�/�
=��C� �� f���"��P�Y�*��#US���,�j� P�	��@q�P	�+�(z�6�[~���ǚn[^�>�e��D�����RU�W2�.w�u�l��B�w}�ۺaT#�<�1�=��&���Pߜ6��Rus��]U1+�5��4(a�,�8��Сa��="ӌ�m�
���� 2 �j�
��w��"��"�2*��EB �Nnyz�y��
f���UX@�H��@�5B�}���& +��GrӪȪ���Г׮��#�T4D�)>F��?Mǲ�o���͑E�L� �*�^!�֭����#m�sÞ�[�FrZ玱Ӹ�Y�m�+������?M��1߽g� i��s�^���@p��<j� Y<����B�DV������(	㯄UY p�L���H�
����wB�;���3{7�t4+���@�d
f��4!�{��` 3ZEx��@EUCU�!T!�T��G2@c�э7�CH�UVj x�i�5T ����b�P�y�����U�@���Q"��L�8�o����{�� 5B�)�Wp�]T5Z@�T @DU�{��3��T�:A ξ��ھ����!C�UB�Y��>i��#�6�)Hp � 4�$�� � ;UT!��⡋����� p� 3P��T#��A��8@ԍ4+q��R5Vxj���z����xi T�UW~޻��b�� |F�45U
�Ϋ�B��C���!��P�@CB���ΒC@��0"ar=�C��h@��咰�(x�DU^ {��CM�@	"�m !xF�T��wUD�qtС �!!� w��Ph@&��(Ua�f��tΞv�{�t������c�����T g�D�a:ba't���������6��CMP8�S"�f��4�}b�U�s�r�񡦸@� p���"���w��k,�LS�����uX�=Gƨj�F��>�t()�k�� t�骦D!�X�VzF���l"44	E ���@C5N�nD;�Ӏ�w/iv�W���VC�ؕ�پ�%�z�ꋺ��5X,�ӤZ;B o)�V�ȵ���
��L9ZW9�}�����{|��gs�����
*"$5m�����9�b�q��IK�Ŧ�{y�gk�n�69�b�p��Bv#��]=��Gi���eɳ�5��c!���>S�|�9p9-i��Y������v�,�w;y�ǇF:$7��������]8�S��K�$l�l�rl�4���XDH����=��htKu�/���2�I�[ 0�l�8toV�̼:�k�3綋���v��Y��+�7gF1�F���.��.ɮ�5�E7MM���.깮��\sQ����w��;܂�R"�k�s�f�p�� ! B"���*3��t+��d<j�@B 9�wVhs�y���v菈��(aȄ�!OY��s�,U��#H}��гUD�8�a "fg��!�"�C!-H�Ӥ���"��Ȫf�hp����b���c��7 ��%CH�@oPs=�uU�GӤ�(i�k�H���wT8F��p�$hV��X@}��;�Ui�]��<G���
h�MU�4/������-I�p�$t�f��� ���>�S����W���H�!&��x���H��w��E@��f-��y@i���+��ܘ�a��GuUh����;��^�8E��
�hP~9{Mf��\g.ǝ'�c�1ӱ!�쳷ޒ[�EV��Fo�	�N��a���Cx����8@�(q��, 0�E,�qUf )��������VЭ5HФ@��-my��� �C��s�V�T0�]�B����
��s�/2b�"6��H֮6Ei�f���Ei��peCT0�qP���DY�k���@�V��`��p��s|� f="�"�7�UbD���j�����5f��j�4=�_���<"�@�D4)�9���W=����/Ɍ�\��AD�-#�$	<����`��e���K�Ke�MUT3�!)���&���j�H�UdY����#ة_����!�z����#T5���Zj�4EQ3B�=�|/;���Y��?#Fxk�44օ�s�ڢhk�qX�(a "Ƞ�ڨj9�{���(�H�rG�@�S5A7���uC���K�������s4/gi���<Ik;m�عX�Ӻ�J��ow�	#..w��6ڷ�JO
gv�\l�e.�ﾻ���>�<��4�3���� dU����%���0�!�jZz1�a�X@�����+N��\�H�{�ws��x��<;��1N	'�g���[\[k��I��[XD"��(j���w<lV28�p�F�L�:�n=�qjȨB46�A�o��y��3z�ކ�A�Tz7�8@�M�YF��(9�;��i���U���"�QM|�HT��a��iõ]4�z�����:ߕ��Mpך��qv�,�1a��C���ЄW�s���h2���P�f*�>�] �p�=���U��>��z:"�7�"����B!�}�x&Ԓ&،E#� �4h+B��uZhe��� �-�"�@C7�����g\�t�/:l��5���A��{r����V���T,��vЭ����V�5��R�45O{����!1ԈGpM�T]��w\�GDv2Es;c�ru!���t+�Rζ5v�iI�b�j3��� ���:�;O=�n�F��hhx�%W|uYj�����^:5f��@IF�}.�����^8�u����c���B͑B]�8��T8kM�L�`�=^����n����r�j�q{�U�|F�5/����:�`X7��C��P�]����wC:x�G�Da�7��`�i�0��ha�>��_W-|%1P�Ϋ«6Z�91�5�T����Fh�,��MH�I8r�p��"�mB*ҡҳ=�=��k�:hi�j��xؠ�� G�˻E;���cS��c��AO�q�V)'�)}ؗ��ԙ�^r�sJ��z]!�^�ْr	lÌ��	Ӏ�������}h�զ�������Xp�wf��������t�5�誹h2MU�h;��T�)RN A5��۫ ݝ"��>;�o�5�^�g���'�"H��Y�@�z�ng��4��x�N�8��WUÇ��� Y�UE�������h#��۵j���)��L�c��� n4�Ah~�Â$���ZzTB���u���n�P�P��j?{;�$��]W���Af�� 0�|�U�*�B��j�;�9�5L�mS#��h p�O�O�O�?�x���^8C�z�v�l�����8�a*D��x�.R�B�7��nAڞB�"�6@f��w��`t�p* ��Uv���A�M�B5��V5ҹ������{u�v�dF�`a������C�a�A�������IE��-���O�G0W�&[�9HU`��hc]���:�:������} �7��{Һ�e3Ϳp*�ƫ���A���u�a�h�_�{Ǡ(��R<��CEF�Y6��H�3Q90i��P��e]�M����C{n���>;h	�xn�ǣ�oo���[n�����8Ge���AN�P��K�X�u�������'�:$�i �I��	�n����+�vv�~�\b����t#A��3F 9�獁����:6l�M����c�MF��W;s4�>˶�)Oj'��3u�s<�	U��S�ND���z0�mF��d��������%2�L�h�-�a1���s!����e*1���U�E$͎�9��Cͷ��t��P��1�!�xE�V@��T�����B�	f�k?U&yp~�wYB���d�}��~	�dx�ٳ�ōU�F��'���Gݕ�X��P���Ɩk�>a��D[�=b�l�5D�*h�3����'<ۓX�ێ|�˛<���떸��a�IGm]�8t��3LÅ����GZ�w���2�7l��,�d_�����x�����VE"ט.�WTu��U�����к!vc���}�闥%R�T�W��j�vݩ��Y�c}��#	4ΐȦ�es�����,�!��񴾩F���[�g4��ʽ��B
',"�v:�3#aMb��~�l���!�Qi�y�rŎ���sL/>!�"��Lv1��D|�l���!m����b$`F8�P��O��*<b4����7I��ڬ�6_{���D"4��z削Ȅg-Ԉv�}��}9ׄ�)�ś�pU�w�4P �1,�j7��r��-6C����a���)���(����Sl�w�t�=_s����V�`���E�2;�����E���o*�3���@��V)�	$oWn�uc#��eeB�;����۪4��׍�hω����]%�v�Ot�&��yG�qv�����A��G@��:
<v�|�!�������_G��`�a4%r!���l7\XK�ݸ�9�"��r�m��Wh7�2I�o�]�:��qs����Ҍ������Q��F�ܜ(�#è�썸1�v�����Cj-���r*[��3\�7@���w��5Ǒ��k�=P&�vv]Ӣ���ŉ���]b��n��z��V���q]�T�)����cj.�0��1̹�֝L�.�Bh��r�h.7k�9��=��]��W�y��8�3Ym(
f��A䤕s@��-֚���w����U'�ߕFׯmҝ2�=��K�a���_��s���<�^K'S��Q���v�]V
����8Ҁ��O��@cr#M���Q�Q�����TGf�?N��U�<b���3}�0�ҋ��)��2�U;��a���4���M�Gv	�:��а����`6�L�a����:Ub���I���}I�\M/E�zi��L|lVT�G+g���(��bϳ
�L�r�V�C,�Y�x�N@ԍ@��U���v)�}��uX�	2��t���^�e
k�93(���Z����Z�� �����8PB�3vN���ZC;��qr�i�J�l������#�����y]�+
3��Z�^�c��Y��4����_4b@������t@��2�����H=a��Gϼ���1�`�M�J�f��Sdxں�+�"�:·۞[�h�t��lœ
�'�yj�4�2$S����3��3�X��$dA���u��s���!9�a���{R�ʘYzo;|-�m�s���8�~�����&��H����>�}
��R�sj^�S��+���ɀ�'�`+Z�t��K7pTɵ�57-K)�V���7\&f�m@,��\t����!�c�t
y�SC�y�A�5��9�7�Ğ�ׯ󝴍;��4��4�2O�0&l�}����]B��@2�X�nN��Q��Qz��[,`t0U1}��r�ӓ���ًl�w����[5&�%�g�����Iz
p���a��a#Yd����N��Wob�z�w���d��͗*��83�>�qu?\�5~�Vzxփ��H>�jA��1t�M!H}A	�jナ��5E��a�I��k���)^"ǙN�*>h�Z��2�mԳ\�3��^�]Υ�q�b�ה��܉a�ݳ]���}�B�i
Y�Fܻ� �`�Mp�)5�Q��k�œ.��,	�-.��K�Q6����>�����	����U� �K�Z��;�m�yT@��ڭWҟiߩyܗ�x�b��{�%�z�%��BÎi�L��S��b��K�U�҇�<�9���n���/�"�oV�L���t0�t����*�kE�D��3k�\}���`�H:HP,����a��5�6���̜�Ϣ=�P�_���J�ޯZo�3���M�ٻ	, �s���2hWU��vj�xn.8N*#R�y(��-v�;u���K�F�a��K�ytI��^{���a�b�i����r���p'��x$	��Be��#��ռ*	�z��9��/l�p&�+��}��>�|�9
�!�Mu�rq�Ҍ0*c�N��<��K�4���ˠ�����m���l�^���Р� ��6��f�����WWv�u�AQ���|��hc�����$�h�� �FϞH�֟�Y�\k<z��h2q��l�r]c���A�F4j۩5j*n�+�6��V��	�Y�E��-��I��֥D��8����[���Qa���p}>��^>�Km�w>�=�[<�I*$齾)WK�3����)�B8�དྷؾ!V�/W�@�W�T�c4�����&7CMQ��w�U@�~�n�c՝�۷��]�
�Vs�*�#�t��ZE5}�:���7�F��]���)���n�~�\�����׻�)|�׺�8��E��yp�'���k��N�E�Y	6Bm���q�*wv.�|3$�=���,��(������LQ�)�۞��g�x��T�_`0�s��L��f@.S&��KldFU��AmaF�(�;�ؤ��yb�Ms��ni-8#�f�h��Ξ�F�:�Z���,>��t��K���P��E��J�-�u��W6����x�E���q弼�ћ���I��@ۏ軔��G�wv6�8��U�c��f�{+jԣIO���q83;�"t�q��]%8u�٦܁�y��I�Iƺ۞@�U�Ϥ�5?�]�:���2孺��� �eN6ȻK)R\(=���>B�}e�.�n7���U��넓��q�4�H5N;�qIA��x��&���W= �B�y����$e�Q��͏�}�'^��%O��R���>�=}�=���[ƛ\��7Г��xp��f�Dk��9ʟW����Vy���1���xo�Q�c��^t�\!�����
� ��Yt�k2�PE*O�=�i�x<Իj�:������'It�>G'��[C8�4�5�C�ܩ����e�����:�0��Qi��;ne�����0�HĔ�'^!MwnR�q�Gb�"���Yg-Ǒy��ۑ�B��UW�P*��U�P*��U��UP��@P��U�P*��U~�
��U_�@P��U�P*��U~?�B��UW�P*��U�B��UW�@P��U�B��UR�(UU
��@P��U�P*��U
��U_�B��UW�@P��U�P*��U~�
��U[@P��U��PVI��e!@�Ė` �������F���%l�ն�(�)$)��IT+mE*�E�� P�	R
�(�R*���D�Jm*��hʕB�KmEIO}EDU�@QUJ 
UR	T (R��T ���T}�RED*�*� �	T� ����
$�ɠ�J)@�PRD�3@>��[����lk�ޒ���;���>�8|��z�lf�ʐ��l�{d�7����[{�⽛*�w|��{h��z�<ڮ��Q{�a��yn�i({5��P�@��$�3�ci,�뺼ʖ���Ρ����x���*�;׶�jk��̦�f�����f|J�|�l��4�KH���f��G��zm<���#Z��Ao� $��TP�@("D��{[ml=����̋��AyV��w�Cejyt�j^����I��^�u�2���ӥ����;٨l�����6ձޔD7��(���^�m�w�/l�R)JT�ƶ�{r�k��kw��W�m��
;���������{Zoz��)m)�x���U�y���l�4��[z;l�O;���mVۗN�k-Zۈ�*vlQ�-�E�<�I*� HIU$�	J����7������i���==5U{�����{׃׶	e��Ry�F�78�����5^��=2m6o=�Q{[+ky���-�5��nћ5�nw*��%U*�H�Z�=�J�Xj��w�m�����w�{fM���^Z�/{�z��-^��
��#ɮT4���Qw�&�S�{�{l�ZqK��[ye�Mak�a�i�5Y)�<=I � �J�!T.{С�{r^�LZw���3\A�-fk�U֔Օ�DP���j�^�t�1u���iw���J��w�u=�J����W��(wo�є���b��*�),��h��=�$��z���z#s:�}��%��tU}g��u"�=��z_;�u[`+Cy����O���R�vt<��(��o@w�� >}�����C�Ѿ���"	/>zjAQ�PUR�P ,/��

]�|�t�T��hU��҅N�����t�}�J�H{��Q�ϭiJ��i�ﻇ� h�1��_uå$y�:��y���)�W�>|�%|�)Z#�^��G��(P�: _UU@�G� >�s� I|��=��� ���>���*�tm��̓糩%)=�����۽��|��)/��'�]��ZU�{�B%y���}�������w��)}�r���Y�����U��~�R� 0�JR�  )� �T� � �2�R�  '�T�OM�  OH5Jj d�O���~������3�~u_Q���O_Wǃ������;\�r�{�G��_����!DGRr��"!(�QP�B��!H���!DG���J"D~�	DB��B�P�D/�W�?&����_�՗vu�:-ӽ�Z�M{�M&��h�6*ė"7�`Bȶ��v7���jw���e��@�7�m���o��0�+|���ʱ�?*ђ���x�`�e�f����w�X�nh[�Qћqfʒ��y�ee��){�9�E��aX��b�GpљM-���z����Y�h�7lȷvԄ��#!�c*&���2a4�m0��X��z��j��T�сL6�P�J̀���`4�)�:9Zw]���<ʈZiw���x��A�NQx�͔n��W�|L���<xoBj��6Ud�4˛M^����^��:�Gn�ge�U���T�[����h0��&�
��Jd���1�M�p��%U�;�	�z)��+�ة��� �En\�9��,��^H��^�h�ya<����h(�G���mD�dm����h(��`�)L)��$Մ7K�N�ɺ����
@ՙH,���0���F�MZ(��e|�,�J��pb�e�}�lm�"P_"������֕Z�3&̣����I��F]ni�6�c-�mZ'r�j�:��ZH,��,~j�b�Rn�.7�@��&M���o
u4JJ���m�%1ݠ�F�{-�U�*��ٷ�-�w%:��d"�Sc�	�G �Fa��1+�t��{0X�񶡬w��Mf˅"t�Gf�Z�D`�͘�,*�]EA��9+v:�j=�񽩰�� T�OT��|����1]�Νϗ�P*�+v��k�S��P�-�WN#�V۷-��"/udPC�j��En��m���.�[�I�\�V\{-M%�m���/D�Ke�������p�b�	��B���3~(���f�4����3X,�YMU9���FC�+i��=����l�[f�f�X+V{�7K�A�1�8�ɘ�b��\L����3�)��V`cX#u�wl�������I��7�@\���Qt��kl#���K8N�G�nC�Xql�e�R�Вn��D[92^�dKTkX4�je�����DM&h�M]B�cGmK稹&��f;OKȒ#���/�Z<����0��>�V2�V�mf�wj��vV^�zΑ��]��J�u��D#�^��D���tMt�����d��[P�=`�w����f��X�<�B��[�v�3G�hYi����ڽ���A����]���Z����[[H����l��)]۬6^��  W���r:��򶋌f�{�O�Qd��P'J�V)S2a&��%1��cx4h�D���B^�� �� ��`b��2�:X�� ���d�&��C!3j�ܹ�֝��EZ�k!sNf�ܼ������7L� קwl�50��i��Z�M\���s�6��pl-�E|w&MX�MJ��taW�S[�7�Y���bҀ���N�b��Y�:
e$���Y�ǥD��-ٓ#���0^Y��Z�  /sv��,byRiDjG��wBgl��{�mZ����4�6��深d�M �uf؋�]�L�ն�ɘ�R�֍�:!�d9y�����L㠴�x�6��S�^i��+�0�5���ñ�MZln�J�Ri��Mܬ[crS�K,d�%�si���*�ͫ�O^��LjH�!^*��^-���8jThi66���vֽ�!��D�ے��o��].�8��Իa��J4�hAMĔ�8(�i,b�))Y��
��F�i�0&��1f����-�R f��1�1�֝Gv�IOI$�,�DӍȦ����K�
41,�A`�����ܥ^�����xR�{���\n��j���N�]94ͣ�pK*�pV�J�j�e1�C{�m�#RҎ�M6rѽ�[CgV���QeŹ�4����=�-d�m���Oq�0�ϳN;z`vZ9.��z"�n��!�d������+RǆƼ6��D��d-�8��3G���>�H�T ��/B�r͵������[Qh�Dm��4��k�@QP�IV=�Q����sS~ɩy�Z��w
���*�$�m���*�{@Ȧ���5��(846�$6 NfɃ2�{nosDm��C���7���[A#���s^c��:rU݇�u<�l�q�ճj��ڲ�n)�Ջ��w*Ȭi��n@%Ƴ(&ë�(hzfK��(�+P�jR�{W��K0T�b6�b�����J,6��wٻ���[�Da��\3.�3Lޕ)T����4�ۮ�1�Ŭ�X�C�-D�5��d\��ǭ!�hTԝj{corؔ^�Y>m�z!���h1�ְ2��)
�1�h��+�
,iژ(Sm\`�ޘ�u�e�:���� 5$�2���7k)�9!I��^�֭:� 35�x���
�"&j�VlX�� �[ha��͗WS��r�"�`�lծ�o���M�%QVf��9�����O�ו2���M��t��(�c`_)�.��;Y(̩����ur�v[��S���޳-Х��4��5������*���ѧ.�7u�GjՉ�`�����i�Im,ג�����7��;2�.ФV�V�/e+)4�zi2 ��u��M1�P�|�5�҅�a�%#�f�y���A�qL����K4���L����P�U�XA�&S����껸.n[f��	�m�[ �:+^�G���*-�u,A9q�,�Hn}�#����0@[t"N���QW*m�å�.�/��W�[�H���
x�y����0�����]�`m9{��Y:$*�D�	@P6�ة�]�Ě٤�:a���wD������
�(fAl��@���l_t*kw�.]��e̹�v�'D�L�Qe��L��;x�n�.i J�b�l[�����ϐ����M��WYZ.L�F�)�y.'&jecY�;ҩ`�f<�׊�; n�:a� ,�u:#*���,:N�Z��u()ұHe8����Aڷ�������4�$)�gb���ؙ��X�VP�5mr�WCjeE��wGm��Uh�7��s+E�h4(�B1Vf��v�N��Gw&�;1�%�!@F��ii��V�f�1e͙	��n��6�pӽU⛧vC�SgЛ776��Ҝ�a���0+�SE��B�͎*tA95�� ket�M����Xv'"]RV���^�o���f�4X-�/#۴ޭ�5X#���Ch�Z��:qh�2h�)^V��e�\�p��T71F�����2i�)�;����[qLt2��u��"���5)����Z6��S�Zi˫{zT��4��8e�a//a���nKۑ�Zsa�x��H�F=M���哊�G��͝�v���(sY	���a�G/r��h^7N�2
�
�fS�x�10`W��P<�uxvE˺Yy3 �4�7-p�,%��⎚�U$�Ŧ��gN즓�dSU����eH��Gk.�{��������SCi�!6Dvf�nY�XUx�X��`�,�ɿ��VC-��շ�Ǘ�Rʇo�ّgd���b��!�JҖ(���Uk�a��[�Eb��h�"����)d8�ݚӷz5��5��.��Snæ�o�.Ƌ���x��T��[�t�p:���a��4�y�B�*��^��ţ�^����u)�.�	m�V-���[�Z���J��� 5g
��޻3/e);�h��DVJ�T,'�X�58� �+5vt�Z$�[�{ f��slޫ�pD����W7*��3w!�7S��	��eF6dH��c6��[R�J�s\-��o�K�yС�Y�#w�&U��.�K�$�yMS�v�z������:��8�+��-���4G��f�4`�u3
��	�N�[�
zG/1,Ot�]����MsMǮ�YH!h�������MB����-k�ݩ��V���T������F���G&
h��M��N�+��]�k!hIG�y�wf�gl�µ.=u�$N6����V���J 3Yj4D�Q�!ŵk	Mrk�o%���ʺL��l��mmś4�]6�hGr�[x$�~D��i�e��5B��h�xvۅ�vŦ���ZȬ��\�1��Ш��z.mj��lX��v��5�W~�YnpR� ٽ��Y��%��*���9��B<�T���k�3��c/s�z���Y�>��0�3e��|�.G��w���#8Nf�����ެ����%Xiѕ�.+�:��f!gF�َ�-����	v�{�T��Z���	��q�Ϩ�eB��Qi�e(:f��h��@,K�]�����φ�I;F\ ޳ �KI�Z�BA�\�m�1yM�jEZ�|�u3
_'E��X�;��S�a�ۻFƽ�J���S�s2���t�
�o(0f��n�r��N�]*�����m�%�d���-e췪��Kt�#B
�w�;3{z�9�fJ��;�h�+4&@�K˧E�Ք�c�������xZcz�V�&]6Ϥ�]�C������j8J��9���,��F2m=�t�Ñؼ�L�9w�+4��7j�����G���#VX�	��1n]dp��\�b^řI�+�J���V��Q�keQ��N�S�M7[0@�S1��Mj���
��ddʳ6��*K5�Le�JrLڑta$��-5�[/A0�V�����3���u}�w���f�St��t҉75�T�4PӴėuwY�2��Mf����\�(�D�2��r�
Cb�A"gNd�mn�t撷���[�,��p�nb0����b��є+%4n�t5�*3/F
ѓaK�6��`Y{a��Սu5���˽��3NN�A7��&�Ċg��
�T����k�b`5gqs8j%t��K\�.���
��]�ؙ�Sp��zEj�4H�i �,:U�f���O����̄�eQ�U>��A�nS�>��֓D}R�5�4�Y/
��iŚ�����VViL9 ��+���ҌҀ;�,�v�'�|�������X$��f�̰hn��Ltpcx�@�����d5�t,қhi{���)Q@��fi�.:ݛ{w����X1�Y�Δ�0T��9
Ŭ[����f-�V!9v�6�a�E��w�D �r�v�Ʌ<�S(����gj�YY�]M!AI�;N�.Dj\"�+ke(D��`�X���*A�婡���[[	��n��qR�ҟ���n��W�&�l��+����2��씖`w$cb�(��M��r]{��Ƕ�
5X���uآ�Z9��rn�]����{�� �{���c�7D�:�ӄAh�\@�N���6��R13�Pq&.���s`c7��pty*�y�7(6Aڿ�82���d5O6�`W�-�Cz�;.�<R�"++]nd�]*f���U*�e�&�9�r�U.�[�;#@b�N%�#7�u��v��ŧA��F�9Q�*��3܇*�c2�Tw4�Mj������mui�e;��S���L�Y��Qtr��d�w�4�u������I�Jy�V0�L��B�aQ�:(f��*�ۀ��Ҥ�����5�B{%��*3c�D0���
��ۃ7�ӑb0X:���'Vf�6p�1����%;���[KjM��g��w�1n��=̨� ����������{+]o^Rjh�L�L�#w-���z������ǔt�w(#�^�q�uTɴsE5-76��;Zu���VԱ2)�B"�,�FKL�trܡ��'p��	�&����OI���~DF|�����R��j�am���6whct�n��.J"P�)Y�(U�A��$72i�#��ۿ]�U�`��j� ��1�$9��See�mT m�)ea���HiV�����YY�RZ��a	�t~�M^,E���e{�&;�x���\hZb��`�#Zk_׬��y���v�µ j=	�P�	̚)U�9x]�QB�%�@ŉ#���8��FQvpMb̳�~ݎT$cO�Jm屆���b�\2��U�D�	%n��cl��)�9�w��h�z4�*��U�rg-4+�*�i�{i�M%W��p*�b$і& -^���ٌJ2\ ���Q&B�o��h]	b����KP�@�/S�~�ˌVe�61G$�t.!����-b��,ͻi"md�����^�ܚ
����ͫ���
�i��3)ʙZ���n5Of��,�Qa�$!H�ۨ7oe ^鿖���w���2��г롺������/��9��3@ólՆljԤ�IjȎ�b]�{/(E�W݊��`SN�L�X�4*@u���K]B۫���;�&�����N�]����(��o�����Įܑ��-PVZ�Ld�SW�k�x�kh��7X�l�[�+w0c�2�������	,T8�)gF����u��C\�e%t�Cnl&k��-7����n��l#�7ʊ�n`/+�vf	qd�a�0�74-��%��az 5�sH�.�5���J��P ��7��.@��[܈�����'0S��BK���c�{Z��0՜F�$:�L,J�|^�:��X��؅������5�6�(�$���j�njV��u��ALє\f�bW��Tu�Am�Z��]�9�r�s�p��6�,d�6J����۽�Ush��(j����f'*'a�2Xz7oK��b	EV��h�#76��/f*�@��tx�sF0�N��E�-\ųh-��*��ȵV�� {VS��ƅ�=����d�B\َ)�MhHJ�K���w&em���~���56%��9�h�q*Ѱ���n�6w��`�M�4��%��մ��Y�fA��ڭ.S��8��%����m죨ڤooAD�� ��[�q�@kյ���g�WE{"7�7�F����
���YQ�g�haP���>F��?f"4e[�P��j�x�� 2ѵ��$G���:X��6����慀J[�aKI;*�9_1��[;��Ô6ai��������$���k=vQ����k'�wojy]�n�t�q�*��ܻm��y�5ώbլ�	�R
7�H"�8Gu���lt�yl�5q�������:�h�5�u��������i`��z�Q��t�`e���z����������;2��MX6WE���@%�f
�ۮyg��2@�g�o�[oNz������R%�è��[�z��e����n�k�\[�t�mkQ��л֏�T��)TU��a�3�����S�G��4�'<�pd�n�p��rv빮XQ�QD���P�Ct��cϋ]�n/�&F�X�&�-��n�3�/Tr��̽��Vx78�ݛ<p�&t낵1D����W4��p��Х	f�ˇX2L���6JC����n�.�][��c+��fu�
$��-v��]l��4t٪5����@%%�s�[.Q��kG9���]�b���`nL*�eu���u����׉�-B�w O�����gDq���x�R<����i�ұ�H2�-��a�^�K��S^&��{'7�q�P���Mλ8�`.@�"3�`�������m�z�o`-��Q��T�<r/[�Zy��cm�xz�x,�,,�T�q�l��A��㌤U��tX�:&��s��=SnLk�1�%�&V�9�Il"B5�X��8��{ ��n��s����/d@���X4��p�{H��z���ۃj��\�E�L��h��e�I�������s�x�t���Z.`��Q%!�Kz�y�s	�4�����^p�gL�֭�p����sV$�m�疦�5E̡�'bϺ�f3h��&��k-�yn(��&��<�:Sy��j��&t��O+��j���،1�޵sݸe��s�t��[q��/����ټ��G'&���u}6����I�q��X�v��v8�ɱ���ڒd���Q�q9�U:����F�5s��ѳ�����Ġf�M-�K�J��2d�QūlZ�����bi��n,dK1�G�i�`E�z����»�E�%�뗍Lk�ˣ�a�xϣ�0�����s�����9�=����c�v�ŗ�%�uM�����7������fEq��k�ˇy㡎��c6�9'��7!pmy�{x'�+�w�	y�^�'����cF�K��<^����u�&&,��5�"�P�S.�iۓ���n���o�k��:���#9�ZGMx�������%��U���Y;Iϒ��v��X5���j�h�369��� ���&�n�N�.NŖ�m�<�oy��wcD�qZ��ǚ,�[���/o5[O[�w�M��,�Y�M�W�r/gj\؁X���&2�ͣz�VVZ�-�R֕lKuX��JBfk�a�Ffj���Dŵ5HA��S+�JvW<��۲�{�튴qm҆d5���.�N7XwV"��ʰ�����1�x��''&듉���Qs��0��U��Q�5n�X���ٸPN�H.�� ;����v�уY<N�;N�1�O�䤞�v���N����c�A���#:xJD>���u=pmf�ԋ�܉lͷL�*U��rZ�W�Z�5&��U\��X��&��p�\�+���<�*�<i6^ܽ=.D�m������^wc<E�:˷my�]�ƙ�
�I _��Ҏu=��;3���+�D��&S��#�x�V����tŷ7[�+exx�ܡ=S�Y��izx���{]]nݮ�ԕ�ƺ1p��ƹs=�Ns̛�h[y3���lQ�p{4qe���M��yl;2�1]Z�)�n��]���c�6�����^Ϡ6*֎��	�e�m�Mf^�q��[p\u�`����1��(�:m��c�>����/&��&7i�*�͞n�����v�|aBBY����.�Qn�j��M��Vg\ה�\J$P֥�&ؘ�L�Bwn��f�{rqE��s�k1�(��T��G�,��؂G-a��5���R�v;Ol�rV�(�:Fۗ������qT�[<�c�3QA���;'u�|}|3=�dy;\.S���	ivb#��
޸yæ&�c��r�, �2�Quڂ틝�\�NzƷG[�{���e�g'��}q��{uX�\� [T�ٶ�7i�[�,Q��t���A)�u�R��eZ���M��IHa���C�������Ȼ�"a)9t������sͬ�t��Ì����=u�uP���s״N�[��K���K�IcY�+�(����yͭw.�\�6����>3���وk,1��.�b,�����8����1�m[19�}�$��`�㫓g����N8y#��ñ�YY�Ͱ�m--uV��eR�۪r�K��z��A:x�d���aB�f�5d���&�-n���㮪�u�	�QVd�j�U�[���f,W`٘�Li�K3.�1qڻ7SE��vE[�=�v�I;�$��9�U��$�vnS��N�B���Ҩ�bҠt�-�v����t�6q�pu��)�-(��h���66!%��1�Ę�)�sR�HK�sYn]4u��Z����n�
��Ƒ�xV�;X�\=1��҆9s�]̆���L���r�5�@_�ȧ4R�է���֪�z�Ts��CY|]��x@`�'��'WIf�
�@v��1ֹ�x��J�ۗ�x�״og����ж%f�3k]^����:cɺ�u\s�<ًcɔ�s���`��:�yh�u��J6]��'�h�lb�5�܎˔nav�Љ+�h#0�K�2L�I����m�uWF^� ӷI�涳�����WF��F(۪.�����mm�\.�n�X�;9�ئ79w�/Z!�1��5�_��RX���50KPSn���d���IJ�BF�R�uf[�L�Ɉ�������f�v�_;MY��V�^��*.X	��a���������'j�tE)b5.��9Ĝhx��(I�v�n0N�!�����cV�u�ak�����\l�a��: �s�<�hM�W+�wf��<���u�����h���U�r܀u���l�-+1���� 2ԕ��=Gm��q��s���(E6-�,ΰ4�Qx,��Ϝ%���y�F�V�����_[���Q��I���p���t�+�	�4ϣ��M��k����	��Q@��3�(�ڑ{'�^v<k�\��ݢ��F<+Ҧ3�<�Ɓ�[Uh탛�a�d���i��8����7����0����<�5����bEe��ֲ���U����)��a�8#-3k�B͔C�ҬMn���m,�)!��3�k�N0O�楇C͆.;uu�zF8�4ց;a�����:�C�F�Q�n�q�(�"-<d�s���gU���BҚ�,h��f��{y�n��UWI�LHh��e���km��q�۹��1�$0<V6k�v"ެ%�m�b*,�џ��l���<��n4�ר+�Daж�#v��R��
:!	�٥6A5�Si�e��E�*0	��,�N�l�n޺�q��˜�u��A�#����ˎ&�
�t�V�.��>���u/m1�;X�98�%B,L%c�-�5���e҉�I��۶ڧs`m>�˸n%Ӯ������7S)�R/\�m����+\������H^��C���kncC�K��c[bḕڌcOA�&箫���݄��㗝��O=�v�����������Ά�%�:֟\g���*�aS'f�`� �16�w<j�nu�L&E��V�99�>]ַ�`^� Z��\��ܮ	vf��R�5�R�W����/@�����Yse�5��J���U�4�'{p���<Kľ��݁�#ƷAnN�9�,���<q�p�V�l�ZG�v��ܼbTS\m϶�7$�Ŵ�����`���H%�b;!�7d"�t'u�/��W�v[��p�tqٹ9�u�Fy�kpZ�Ɣ�f�3�M.+j�F�Ӻ@קiwN��ۨ�A��Ic�	Ů:���;���m�,d�Ms�����9fa{B˚�.e�ke%$�d��Li�WU��rԉtP��dҹ%i�;��_7����blo FP�k�;��-�ݨ�fV�w[��r�r1������L�5b����ͣ���1�t���3�����+,$f�"��f�e��e�Rٷ�����'��m�c��x��Hu��=���(�n�r�anW`�ܸ�'�;���n�Rv�N4�:�r�d��&�VW���u^�%HX��k��A!�t876�GX��<�lr�S���ˌ�JG5<��ĩtP��s�3�3��#{!�v���;ѻN��y�>@��QN�-���S8Bm�Զ�J�]d��'l���9����=��n�guӸ��1�
��������@b��赌��I�Sj+��;X�6�@�\���9����ݑNz�i�]�89�sty�)����lGf�؂(z��j6N��c�|�^px�N�����X�� U��n�l[���z]F�;��YS���ٹ��mc��\���n�8��wl�������ck�
��Rkt#Մλ���κ竈8�v��5#�6`Ų�GJMV�3��T����v�NC��tF��B���0ɱ�.#��?O� �#�B��u�yУ+E(2�g;BST �_m�� z1Z�H��QF�s2b)��,&,qQͷ:-WG���a��ӷ��	�q͸9�}��h��cH�a���CS��p�C�M��p#���(<�O���}�\��h�����K[�E.!0B��{���� �6���f-�ݺ���&�7
�l.g%��U+��P�m�c���; ��e��W�	��<�g[��: [Z1t[)�j��ؙ��w8�r�dU�8ܭ�{i��g#�փں ���\L`cJ���M6ȅ2g�2v8�-����q�P�����hE�7;��\t[��3ـ��t�/&����v�]����8��l#�w{sҏ���e6�˞'�4��a2�
U5?�B�P�D/�(U�Q	(��"!(�Q(Q1	G0FԷ2-��N�h {j�-�W<k�S݃��{qF���ccGgXLg���u�"7-��B����c%�%�����Mlk5�5taɷ"���N�.����\Yz�"�'Q��x�cn���=�Ů�8L@#{]g�nG�.}�a�wX'q{.�et�Oq"�L�˸!PѠ�m��[��x[�=�ei5:5��f��B�e��X۔@�2��˅B�ή[x��9��wY�{3�Zj�%-
� ̹���sj��r/gB]Vզ�	XJ�9�ی�E!]���b��u����>�[9����=���&#Gc�<�s��s'�`F��k{gg������w����]k�`2ʹ+-f�Ha��Z�kGh�֠��j���>y��+������=��3WBT�,̶ѸrhL��&�W�m�f�;im�l^x�XT�Q�WF�٦��g���z�<�n1{u��	q�W3-i�@�n�3jl��m��K16Z�c��j74���.Χ�|��;6J(Z��a,�R!p���,vٱsֵ�.bL5�CSj�E��#WV�%82�FY��ˡ5I��3H�2�mɥ."& X̱�Fڕ�F4�ݴC$e]�v�F�=��e��V�:x�uY�$�6����ҕ��W0ڥ�B��9�v{<�;sz^�[N{;��<�nrx]i�q�u����J�u�Չ�7�������2���e��]جX(��&;ll���4v�N�P`��^���k���un�x%�7N�<s;B�s��k]����IqyT����7<�X�t�q�Ol�R�Taӑ��.�P��y�+@m�ŹN���@Зm^S���s
�ɹ.�6����e��Q�0`�c���K����ؑ֎��5�q�b�R��=���r�ĝ�x���'Cҙ�]t�cI�X�;E�qļ���m�n�r�Ť؄�K.[.��Vˌ�.�h6�3R����Y�
��:�=t^�Rgv�3XbX91G�ӧwt���wwB���I@BP�I(��$�BQ �"!@%���B� J@(���%	B�
�� �(Q!DBQ"% �D(�P�J�*jL�x9c��ڀyۦ�ֹi� �!�7��F��F��L�lѭb[]W���X6�`�85</c��8�qK������׎,/&3�3��c����^�m���޸s����ؔ�;ԑ%ګcbca�J�쐼���[�)kۓWX�͎���'9Z����7�g\&;k����B�0ֵU{���})�1�z��k����w>YC�=rJD����'���m?�~U�ùF�w�F�e8i�Wa����@���� �m����}�p�Q�
.�Cp�cM�w��y�UC^ �	�l���ɱ�x���T�H�އ�
M�q��n|왲:��N52�l"�(�#2H��b��ٞ����Wu9T�|�}6#gyx�7�P!cg�75���Lro�a�����-ȅ�Hs롬l�(`54JRd�`EM.z�`�@Q*��(�j:�;&�&�7�չZ�~�\z�������IB��Kֱ�J:D�S�d{S�A��
��<N߻�~)����/Mz�(�:�ÿT�4��~�ߎr7��[�!Hm׷
rK���q�t'c��X6�S�Ã��[t��'!�2�kVԋ���t�������u,x5�xe�)�<�&Rr�K
���ek�uc�~�}���9���3YA�q�'��|u이�X���V �Ս�vT���w�MCW��
њKD�vx9�r�,h�R��DF5d��xF��^A�1�:]G���H��&�4��9ܘ�4��j]Z�ˢ�h+��Q���(J���@�2&�V�q�l
_i�Q�[���}M^K��;�^��D��r\�&�K�ǩ�����dC�@A��m@ �;xvVv���h���u��al`%�Z���o��ZSN��½���X,V�:�͋PQ�6Z�RH�MB���įfN�}�u��f,OG�-U��yL�+wP�N��~�wG�6f�O�kNPM��p,>>���|/���Zℇ�h��+������SI`7fQ�%HPlU�w=K� �kS�ln�� 2&࿥=����3��X���g��'��S��H���X�ˏH�?3N�҅Jy��oZl�%!��+�D��ΧV��B�<c���3vg$u�n�����~�wA��[�sb��S�Eb�Aۢ�6ڌ}�����,���72z����u��[�ޏ
��cM��a�A)�����n���W/���¹�3#��т��]AC� �u���<�RU	$�[C��5n`~�����1�$�~>y�Y��Ą)L(������Ǻw6��$�{��3n@���ݽèL�:��NU^�U���S��CB�t��
wb��@����y�\z@��&�l�~jAC���HF��3Ճ�s9nf���C��ê.���@^�}2�wi\_$�����F�-��I䖲��A����kM�-u�	p�����rڸS+*p�	���n� f�-F��:بز]�;�	fr���*�#����}��v�F�=:��HЀ�=�,鋮�4E@ ��rO��tǻ�T�S]
`�M�Xtq+w��Ο_JȠ���y&�;�í�.=��8	uy���ԣc�	�L	�r|�"2����'�/��R�Z|v(.�P�+#�~M�C9��zL��q#6�e��ES�9UT:��EJ��h��9��h�Y4�v�q�|:���0|�1۵T��ү2��S�kǏN�j��V�"w6%z�V�:I�F���T��;�r��镠����Ktv�hAG}��M�Ս�ǟ�m����_��p�Ҹ�)ȯ��ӽ.��=��]�����s�Uw���\�C�=듗�:�mw��c綁U 7+j�F�∤҂6��|nyv7I�/bxY�,�8�/3iq�ot��N5��y�-H�l�����g��OϾ��w� ���/i,����j !���ܱ^i�W�v=�

h����B�m��2J�v]
�j-.2���4�J��Z���9�>�*��N�,>�W<u{�7;��Ѽ��-��Fۂmf��ݲVci�8\���ˤ�Z�>n�_�E�Ma��%U���gmg��=ŭ�X�xjz��>��Y�>���Y��a���F8�R!mA��n=��\����z��Q����}�����<,#&L^�g!0���Ԯ>�"���C*���)ry��1�bb0dN9x5�*�G5w*}I�[o~�|�`�٢�d�_��*qr�F�LͰwه|���
l4�yj�v���n�(%��g����0��i��$6/����������I��"����!)�f�����I�����ї56�Y���bkjT���P6���ݜ*��yM��n�90iMa�wa`ѵp�B�tJ�.�l�j=�s�Hvh�c�@h�]�]���be6��y]Y�/�c���G��<%�/[M
���p����ό�l�^�����̘c�7]=�T�֦ ί;�e�vf����{<�ȫ�wU����,���]j�����nP'�.��y�F�����7a�Z:,[���/g�^��3Y�:�2�jL�0�:!�:	*���qF� �[�6�:8.��9��g�g�gE�N�ʊ�C7���7c�m�V�x�!�PKu="��ʼ���#ޡ~;���i�
;{,�~lx¦��^�;k��䴾�Of�Y�z�������vڦ����R�DP�=Ho:p�^�v��k����**W�҉��΄;��W��X�
��R8YOB1��>�I7��M��{O��E �~��t_Do1��R
"��h�e>�N�|v߆e湚솮��Mm!����Y����r	p�-�nݚ_A4ڱq��\/��`��h�6��O]�טj+z:f��u���{�9�e��}�~ynޣ���e�,Ź�R�/8��'6&�-�V��ݰB���w#d�*�қ!6��+C��q�H��yN���k�	]K���ͿE��j�,eF0�S���nő�2��/A1��%�H�[� kJ�G���M���E/iX��s6����b�.�{�ş%�=�<�����6�B̎�Y ��u��#Y��v�+�T1|0`�~��k>s¦�4;OrH^�J?"� ��Wr�z�a?s3#Ώr�����'��o�([�bƜ�bG9�L��WW{އ��p�O����WG'7N�n��p��G���<�Bkӥ����)�%�*"f3	8&r)Տs��/gS���ܻZ�� �4C0�R�|�D�*<U�A�4�l���$t{jy+`�O���F0�-&8/i���\U\�r��]���={���SA
���т�!
CN���]bϨ>.)X�pt'�^�6����!���l��6���v��|)a��-,nl{'(�j�v��p󹖍c�7��E!I��L����䣸�&4)��s��|e�P@�� ���^Y�:��.҉� D�L��k�	���f��̷HVG ��}z{��MR�:�/�[زt�2]�X�7i�����������l��|6��E����i�#/�P4�#��q�]�7��W{yC�Cۜ�����m�K7n����Rj���ĭ1\i���DF�2M�ؐ�M����߫o-��6{�j�]��`=N�*���!|����浆{��=1����i��	1�Bb�jj�u��&�����7���?o7��lNrL���,�'�o� ��֊'6���Hw.j]��֘��T�u*�۪9ƦvA�Kc�n̞,��B,���Bv�k{�l�:�K�ܲd��߽���*IE�3�RO{O`p���|�P��>� QI�vU���l�A�t�=�������ᛂ�X�Ѷ�ńJ�c	�c2@k��]b��(�cv�����%%�������AQn�d�c�8d�WB�p�	6�.28�e7I@�7v�g�+�z���i��'p�X'��늖B��_1K (��v*�QD�o��`��>�v��e����P��2@�Zh:L�H��4ڡ�ѷ-����^X���׷$P*G{{�mg@qձKv%�X[]����>�I�}��}�g�L �Ϙ_����K.$��ͻY��ZL���{�p_��Y/�3w���]�7vˮ��G�M��ZhP��y��Lm J��⎝ɢ4_f���FV��V�Y�)���)h��0G� �&��2�7����t\h�i
r���ܞ�	���(�(�V| f6�^e�j!����e�L��;��ge$"���.��œ�(<�]�(��)P&�v�k��U
	�8f{+l�te�`���[����k�GT�63[aKb�p۞���}JLr5�')c��)l�FH�4�M�%�\J��OM���Ã��'N־�m�N��Hڛ��,W7�˩��Q����"��ٔ��%T;U�Yk.Ns�ཀ�NU�i�,S�!a��ѱ>M(Kp�X�Ww���;�x,m�^e�-V�+ͳ�W/i� �)v��ҩ^���\�m,�h� �&�9`���ES���[W��2��B���N����J4�z*lJ7xzl����S��/J#�}��)Hg]�1E���Dl��?Os�,�����o�!l��M���h������������7��=��A�t�Q�~�3n�R�Y˘��&ҫ�8�Qѷt�7P�w�0�R����%^ZpJ~˻︥<�,�Z��6�IP5�eN�y��}Y�Z�	�������<���lxF�6w=�ې�ԪE��h[na�E���hĳ2��'�0vEܒE���d,ں�k-��-C0��	\\��E���yf���i�:��GR.��4r0\��VR��H�gEG�zض1�%]���wUmtf���˹��&ӈi��@�uф��p�����l�Y�M�U��t��e�����e����n&қKëؚ1����1,eV�mE��jR�*A����Y�z�Bhc������7���y����@���S#�6����Q���^m�'�?�F�{�Sf4$-�/�d�:�՚<�*{�¶�,9*��@��77��9Iw�蘍��b�r�З;2�̠;B���}cI����@��R�jD���_Ic�ovp�A=|��3k^�>1&U-*XU���,Ri�
��;�7j)��&'#�k�F(��	�=U��f�Y��ǲ	�����vM��O|�_���i�X[���������=�r����/jF��^g��x���+ڭ< ��9�/3=�=.)�L*�$x���q���3R;�H�mA"��»���n��ݬiM�%�-J���Olsh�b�`�LI(�q��0S�x�s��g��T��u�{���f�������L0���*�#DnV�V�1 fT�ϴ��i���yv���m艹�1�l�/�~V�����7�]56^�껝b�B�.��0]=Ei�+Q�]
�'N�&;����6>�ǅ�bK�:r<PK9���K�([BfHZV�d�Lg����h/]\ܝ7cQ�����LSm�XXm�LSٻˏ����;���r��a���D����r��2h���ϻr�u�Ne������-�l5H�
l�Q5�jc *Л��
��i,�G�U�A��v٥�Kv��|�>��֥�ǳ�:N��)�L��&
���cc=+-{�V�2G����� /�\d!���c��:jQ���m��d�m;mɋ�%\���P}���ϐ�k���0f)L�.X�; A��v��� u�8֙��|���չ����zj�>L��qlG�{�҄΂��ƝZn[������µ��S�=x�~��W�����B9]�����R�Vϲ��R�=��]�c�c��s�k�i�
�􆋺����*��6`^�#>�@�S�K�EjLn{�q�����MXzK���$��h>�օ�ɤ��RTk:����۸��Z\S��8�� s2���L��r�J����a���'5�W���Y憢�Э��"S�rb�M�>!'��a�5��c���\%6�Wv��;Ȍ|���R�1���j�+zZ���{{g�Yޘ��x��J�Cz���9.'܀T��Z�B�V�ΐe�}+�u�)ŕ�׮`���֬@2�6A��_�&)j���|�%�3W3LM�"+r�Z7�n����}��l�w	�h���VҖ�|z?��-K���p�*!Ԇh��PwCG{�/.,=�xȻl,m�,;�d�ʇUEA�(��ce�V̭ɪs�}W���F��{Nx\����G�dШpB�|���{z�E�:�q�&ɖ��h7��^�ٜι�t�p:���FP�=\��6^��2��k��;f9��+U�*�����e�L�זd����֎a8ti�d��]���7�6�a8.i�:�n�|�9�!����7[Y�i�z�ˮ���7f}s��w��]��j���W����b*�p��DW|�l��tA�O%��[x�S��Zq�3*����Z��)����׵�غТ�C-����X'v�9ӻ����Buv*�e�U����ӟ<�۩Y��iB����X[b��7�D��%�xi�]�e���^uK�lp�y;��R�G�㸤�o��9����X}q��f��\%Kе"���Ν�3yَ��qf4�;ʜ�����m�4� ��,���P���G�q'w�xv�k��O��y��,���e�.����=�.{�Qn`���%�)�r�Ւe�oN��{騏g��SUF�\��t��G��m<d�$!��)Ȩ`�Ay=�'!m`~��h�=���:8\5��£��{yݵN�X.֞�s��L�fnWz?��H�>w̭�y�ߣ��E�lD��`�[��h�l�u����e�I^�ۯ64�	���Cm�~AV8��lj]�qF6��]2��V��)�:	�,�d��#�������=�3 �h�-�}�޳P0��wV�Lٛ�+nz�>z@�J�����*G(�^*s�l�I`߫k�EǋQ݃`���^�w[b%�H�*A������]��=Kե�n�$�V�[N�F����jg���X��W ��$��"��+�ad�I�w��ΨF���U�[�t(�ڑ�X��ף�Ea���VɕM��Tݳ%��x�����5����1�¨b kCz��eV�:�tNPy�0ݸ��J�#����3�hF���옠�]j�Y2�I�5�h�I�P)j�Crペ�L��k���1���?_h�޳��Tt��y���e� �.'D
�%_L_ZV�����w���سա����X,ɮ���g�݀�c�;y��VD����4�r�
���DF��̑��+)�m�z���d�|p��`�OZ�y�LM�L�rQ��s�;��!��������"1��D���rپ��ᴫ{\빫.Q���ZLhh6�T^�뵱�۷Db���F���{�u�}�����Х Q�#�9�+I�%��Ŗ���=V�}\V[��)���^����<�'>�o��I���5������8�!�!x��������D��ׯ0�����Iݧ����w9y"���cxj�!o �r�h��B�'P"�!��Ղ�Єx�(���Gw���Α?	��F��pm��z�`�!����ˤ"��(�[�sm������.�X#�־�Ԡ�}[�+H�%�]���7�P����Z�2v�u�Y����|61���s�j�LMZ�̏R����i��(A&��Nۧ�ۤb�瞜^4���0.�tsB=NN������PF�{Kڱf��\m`����Q��R��Ǝ^@x`���w ��G�l�gD�u�qT��3�2M�cX6�ZM&�B���ˢ��c\��.V�V]���e��5.�s����s+�ؒ�	q��v��Oc\)V-���x��l��eN�Y��[�N.�L�ñَy��-�㠽�c�\S�}���n',���i�3�[=�a�۞6�t��%��Uw����=;��4�������\Ƃ�'�L�pe �|�{��,�3S��jvH��9�+e�J�7;	ʚ4ʧ�D��{�'[c=�,*���|�l�"�t�
u盪�ƒ�D��=úB{o�;l�����la�\l����H�4
`0�F��ä��O�Q\���{8�<]6Gt����~7�'܊O)�����=G���iW+��S͂C�:<%�.<m2��z}�]^�^�	w��k+��ܞ4m��x���1���0ˬ�@��>a�� ��1$d�F�I�l��)����uQ�7��L.S��e�T��gk�[ä�O(��-����*���McW�j�&,"+^����ߞ��u)�Yv�&(1��mћ���V��[��Hk.�y�7qq�������K�)�b}���PQ�.Gօ���3.���U��8`����{�^�aٗv�:�,]��Y��Wq�ߍ�k��8�:�R�ʺ�9�P���2b��|m����-���]�m=��v_Y|]_r�7m�;��5�K-v�V�og0)<Er�{��K~��sV���*�QOE?:}�[vf�D��$)Y\�D_��S�l���I8!f�14x�7jςҬHJMH`�ņ�������#(Q�/kb�9�j�����R�N����N��]�/ֺ�!��5��O�#2Ya�L���kn��p]�QD�+�!J�Z���T���?�}�ʬ�.�o��6=��61 �D��&8�Η�BS�kd�CG�J�B!�}ިF(���{v��$�Ԉ��Ay���L���"ozɗ6n�廡�Kh'�4ZTID�P���w���R�3�K�gK�\ ͪav�jTh�,+����e�S׿�y���|��޼�{���%{�Tx3r*�q���ex'l���e^ӱu� �,z{�6x��ķ�l���d��b�Q�n���"��up��m��C�^I��HP�c�� �r��v��zbV�5���j�]�so͂@����
�.D���tI]ߘ����M�mrPR��hs��E���v�ey�v1��v��G#F�Έ7���o,����Z���G����j�e��7�ޚ��;v�!�۞����K��Fl�{I��P# 1)�Tr�]iY2�Ǹ���^���Y�:�|ov�M*�=�bWn���!�8l�z��E#�kF6�$2\��%���(�}�xr��7KOt����+l/[����ލ��\�ʇ�y2���d��c��P}&8>����=���{�l-l�%&�����En��B\������R�K��f�!0��)MORKB[I�מ��lq;�_�;�3�~��5

��j\0��2�"n��9fa�+tID�,��)CI=L�����{{wefb��-Il���ny��%/�rWmq�q�,"���ji�y1:�`�yи�� �p�LJؕ`�9:J0�PS�V��zc���L/��3��ӣ��d�W�ې�6�fo/Y�>0���:\�5H�§L4ф����`5�:)����xi�����~�p{<��^��g�6���emZ}F*�q��8����m�W(v�Z6��8���4�)��š������n��f����8J�ҳ+h����~�R�wK��X"�ȱU4Q�x6E3l����i~K�C�*L3�r�:��e�t�l<7GY�=����jHtJV+���gg�O���aF����m�d�uK�K�}G�[n,�U�b�;��7�-5��GMR�X̦�fb����@Vz�����XNuV~�*�$����T�v��!��t����˱)�Q��b���B�9���"Lq�JEXQ�P��\�ޢ���nq�<(b�On���W�(�gٛ�oV|w�u�:r�=��b���,m?0$�|�1�	
Iu�/CɊF���ܲ�!����0����l�Y|Ǌ���2V��祿k�I����dq_|�2�L��b�ڨa���[$�d^��g~��l�_�jݘg�Ӽ�*_Nɒ�%2g�9�^C5�������P8���q�T,�I��C�:�Y�� I/*"�_fd���sU��*�/�'�}b��'D�Xm�DSKqiͫ!�fY��:I�ݳui�P%��ʕ4���
���Ї�{��G[}��h���SWD�/�e�`wT�OE�!��[]��r�^�+�
��٨�=j�4�9�b���(b�8ћdP��ҕ����9Gby��Ɏ��n�<��C7��۳`��t\�;;4g����mq۷Xg������$�-�U�0j+�).�#�Z��9ܖm��y[���u�׃j�&�����X��C�,ک���\�:�d7�aRz�kl]1�']�o�d�PLG�s�<��5r�18'�6d�;���<���ԭ��.wm�/<�9��a8:��kn�����YlsѸ����w��^����)�$�A�r��r�'�r�߄ry|��;F�����M�N�K��T;�cN�L�E�L6�ݿ6���<�*n6(�4�fm���HA��y[�%��iޞ�E`l%o��pҋ��zC��p���>�$m��	�k3�����������#�A~;��`�5�5J�F�x>���;�E�6t��V���=��%���j��w��TQ�h�L7���]���J(ֵS�n�ж�1��Ǿ�>� '|2�o`�!r>ƗX3����1�R|ʌ�'t����8R.�>a�M5��#���ԽˌX'E�=���Y�o�ư�4��O3!��R��[�藊�S2Aۊ]�VOn$��@�*-�h�q�aHJf�6��ͫ���RmR��,��m2GCk�������<��������'h�o��-wy���}���N�m��VJb�ɤ�Z+ƍ�ٷ�F	�!�5�cZ���і�2�y5��ژ�>4q�V5���B"�J�3�R��7!�y���)۵��޼���1�n�4u��!j��%�.yU��=�.grɉ��|��fyΆ�Lm�/i���J�˒����~���~���3�
[�H$�FPP�vS��̤���:s7�Iѭ�,F��χ+	f����E�bRez�#o�J&Tr6N;�e���&wN�� ��!�ܦy;ns��ǪU��E��ޮ���Qa��J�{��Jiz/�+��ʑ(�a������54��a���Tk'�G��b���V]�� ��O���g�{~�ڕ��F�	�W<kâ�)Ss��~��_��y%?j���o*Xoj�ty��۵�Ϥ�&���\5�sq����� -��
2ӄ��`�!�R�b�:��}D`k�u�+J�6��^�,��$���>�}�˙ª�qu�-�`�!NH��8n�m��+��_������ո��z�"���ߪ\
/���}��)��Q��ѓå���Pkq�Դ`ދý���h&�AQ%�[�i5)="����_�+�*���)[����{��9����]���2���!Ŏ��cPeڊ(aN]5WAt�"�M��B��x�\��e.�3f[��{��������E.������z�~������Q�#�ɞLzmPy�&���φ��crB�����1��z�^��Ǽ�⹟p��(^L�G�5eQ8kJx�;����ESr��ey�P2H���l;/7��K	Qc��`��E�z�V-��)��߬���J�������� T��E_U��� ���%�$�]�ʊ�v�]���]�`*-{D��<��7$HϢi'�*�U�����|��=Jͱ��5�Hϴ�U�v���:Q���Ց�/;(�<�7I-��>ȴ ���t��OϜT&2�]u�`����[_p������s�h6���M�^^�����0���S:(�>��򝷷pq���ϚM:H:,�Mv)D7�ni�k,��(�H�}Ԣ{��������5v�d��̾��#��^�P< Q4Ӂ�\pnxk"�C_np$'��_# Q;��-[Ba���/���)�E�'_mHc�X,؏>��%���$
��T���%�,j�v(�n�b1�"�}�Ĉެ�t���=��ɣ�u6汚�,��������
b�I2�."$�v��J#a	��>>Q /�>f��r��=`շ������n�4� ��dY$�E�-�TA#I�Rkηm�	5�y�D�p�g�{˓��jx��6�sq�":���$��L\���_f��w�v�}�Xk���T�[�F&����^�U����v��s���ad,*�,���Fg�H�B�rI��Z�Y\k��bv�Ȗg�ח���8�4{�]���z��i���00v��8�h�U�<z�V�":
�1�w�k�R�l�섻ϓ �^��
��4q�y�3c����v!�^2�Rμ����#A�l��Da�$d������ޖWJ�{�~TQ��%:nG*U
��T����8��'�u��uEVd�b�q˵�x�h�:�p��	&ڸ7.l����ڿ��e�`:����WKo�٢]�!�̪��	�S�<���q��Z������>���sX;��ʼ��d�SWv$����H��c���n���&�w��r���l�8��P��K�4�W�s^mof���mԬ��Ivx8-�ˤl�K��7���魡+޷�F��]j+Y!����*��{vH\�K]r���<6X���3�h�{�x�
��U�(���u�=J�.F���·��{;"8+��j�	CEq���$�&L�4�������M��Ht��W\�Y f�ܶ5WiS�d�!�&���)�6c��O��*���d�5�mL;Kb2^S�Ib?m��C��.��0�`��VBL;�z%t���͏v��j��Q�}��w~Ooev���B��]�ԪS��{�E�:FN�]`�Z[r+��+�t�=�JV%K}uûulT,�x'9�gk��%<�>Z�L��� 5կhC���6��z�ɕ�t�Q��hӨ�CI��x/p{kIn��b����U�ݬ�l�������ŵ5��L��R,+jK�³��r1�}ѳn�S��f3����
��T�^vE%�qXk#ܲT�R
]�_e��"�rY8�l������T���\u�ŭ��4��i��մkd�0_���67��F�ۖI	ڇ�(A3nrѻ흏Q��9,��|��(C�2.�I�uS#�J��T�:�p+�Sֳ��I;�--�k/���W2��8/�X�s8ԅgq�9�֎l��$bX�|l��ppG�[]�lдE���^�aJ,�c���x͊�4�[,	�LA=h؍��g�뤨���ا�Ѥ��[�a0�=n�Q2<>�ۻ9��L�v뛞8����ua1Z�ƺE���`@�a�y귵ö�!X隂��ΰu�.7�cs�����`���r�3(>�y^�?����o���w6؟`ԙ�l�9ȽJ:�#�n�Vs�<`6�`fi�j�sư)�ܴ�Z����,!L�h�;0�vo ��mGQ�j
+B����k�<u�9'K[� ��VhKF��M��q��=�����������ܨ2x^x�s��/JY�0vK���f��N{f��t�d̼���i���
�@�J����E��iuZƱ�(l��J0�]pVFn�x�g�\�4u�<p􁎍0��NC�9z�m�BbfW&�ȋ��e�i��ds���`�W���1�§�u���+�\�s`s�(��k'7�+��C�Yc �՗����5�j�$�=�F����4�[�z�e�]��u�HBu�f�����4���e�m)�퇒��<���0�L�C6g+j��@fe�q��4V�N�j���AA]�Ҩ�B\k����׈[�f�0n��ȼ�C���n�z�^�䍺�踔�jyy��f��$u)v˩ZX�o
uà��g=�#�B������{'c$;K�X��v��7k�mKt�3�v#.8��&78K��(����h�ea� ݲʦ���8��v��94.p7^����h۞��@y�4 ^&aWP���ˍP�n��+�2���^���a�����"�	5H�:���[����㠂�c��՞\�3Ntz�0t:U7:�pg�ٱ�f�=��P�w9W�`�������:�r�ٌ���	����u��I��5��[�β��x2r]�����;�v�eMi�:�(t���,�����#���8�p�4]͉2��b���6in2.��K�.眕I��������9,��*��j;W��wl�J�/.�6���YC���B����){e��%\�	n�	���XQƖ������abE�.v�e�����Vй�m2F.���t�m=	n^N^{F�R���\I4��;q�Ń���2��\ZCy|��|2ָ��&�MF�$nz�5 =L��MV���l룻J������u{�]�iۘό��ڻc�ht]Q�g1$
Jl�%L��6F5!�]CqY���c�����M�\�B֞��*q�[��D�'czYe�3��$fl��a=����.��Zo_%Z��2�2z�P�K���Ɨ���+.7T���M6��.���w���z�
���1�~�+����w#�kP��@�9�[�@������d�Y��2K���wcǶ��{(��/�G���֔�D�Z�&�N,��㘯-��6�����cmOq�)T����!�\��ЏkS+(�̜��w��J�h�T5>dm�|/�r⸗�����J$��^I���T��y���QY��&�>�8ey'�^����cӑ'E�{�Wê�p���h%�(�
B�b)Q;$�x5X}-t��#Β<^����Br�ut��+��5�C�O���˱�����3՚��$J�(��f0q�t��bAu`J�Mtģ�Y��bh:	��?�%��`���qz�8�"�������s�ɞ�!��ң��cARgP��ٝ}���X�n��}`݈D��������B}��2i��}�p���j��~�T�/���Bf�MuM�B[z�nDHԯ6-�d�;'+ј�@۝"1f.T�� vg@�>�z�7eG��6Ib4�D"cq5eʏ�I}��MӀ]t�[����^w�S���V�lo�(!p4�%�`�M5v(*GMo��M>��!�����,���G��޸�^��M<o��
��{�˿��:������ X6"�<Uy>k��j�'M����~�#&�<3��>�%1�^�2��fF�����Bʕ�M�p���d-�XP�E��\��cޥvm�nmL��ƍ��/�#=�Z(AL�C�K�M�y�x�6�v
�'>�Q�p��K lT�Rd�d@��g���M��{X�:� Tfo;�>6��x�n6� ���-Ö�G������s��"gP{PGC(�d�Ƙ�`y�۩eWKQ�l��:��Z�85b"j `%�#���d��|�ەg��,����=/q��o���λ�:#�;v���V�"2637�o����n��RA��F�+�$��ӑڛEwl���kl+�{.1~��uЛ����j�͡���}ί-ǗD�G�sD��n�;�ҜX����;�vw��E[�W����6�����ۘl'��
PP���3�x�x�"�F"��٘�A��F�L�����P���{������l''��C�c���^�Du4h���k�J������vCa�U�G��� �ܔ��a�&Rl
���3a�ub�X�����>�^]3�Ƃ�PcB�u�-�41���r�9F@��=���F�a�����32�����A��$��j����:<�`벓("��F��r,��4&%���%����G`^��Z��B�,��v��6^�T����^[�sU��:��&f]�ѥ+�H"5(D���r,Y��[�� ����U^�ɞ����QF�fwsw��6˔Ü��\�MYܣU�3^kֆ"t0lia��l"�Gwc�:
���c��^N���7������Fwe�����G �4^K��,$HX�s��v�`��FL2BA�G<V�?7V�����7b5'�՟�9�#փ���}|�s�uD�C,sx;����
�s~GD�HVք�F��~���\��0Qw8o^f����(��o�z�6�fu�����n����	�ɣ����o3؀h2(���(NGH�	�kA9ъ��dլ:�m��#�u����j����:��['z);/&��n0%z'��K����IȤ	B�a�,6�+���Un�b��&�a�Qs� �c]��2������2僑g#���<�ɓ�j�E�<	�h�:�v�}���w��R�j+yr� �O_7ʹ����l���[�5��]ڳ��U�T��޼W��-�����[�a��՗�?z�ZA���0�d�T�L�h ��x9sŒ/ ��1zA��$U{�]���M��Gz���.����]�7s �جR���$Z3J8Z������x0%(����/�}%�T�N�=VS��t��[�SD��K6$�E���y␍f3-�Me{�_����{�i�O9Wf:��y��㭬����Y��Opg���H�ik��Y��,���7h�d��l�Gɩ�M
����
�L'wү�s�q������8he�Z��&��X��р��(e*�x���?(��6)]r�sӣ8,��Ц�&n�Įqq01m�]�d�'\��-��E��:�Ώ95�狒�3��b4,W�1�-��&��c\u��S�9�&�m�̖MN<XgZ�&C8�Ε��R;<�tfX�:h�-;�ɮ�SB+�S:��
�H�p��n���S��c4<uD��:�\e��&�3���Nہ�Ggn%l�z�����#M�@1֡��D�Ȏ��}���$�T<l��|�NyW�fP�AG�w��/<���o���#I��PP������\Ot�zKЃ8
���JΗ��I���vR�"���"�n1n�1��:}�3�`��k�Wu��R�A�F_�mP,c��9Z������}�/X���j�o]����ٛ���OY��Zf�e��gZ~紅Z��t���w:ȱ�>k0A�3q�}*��2���f]#ڇm��D��JTI�:��-�6����$���0�#V�;���]� 2(��1�Bl��5n���<n�z���ˀ���x�VO8 iƘ�)X��}�.�\a4��:^�kُ�;�M��U����s�1ޒ�|��V54�f��"�ȭz�ͤGġGGx�vc��bMd�4nerg��xpA���œr%DD$rI�B�\��:ݛ]��Ol݌:������;W}���h���^{�P���7�|�����ut	�U],Z~Ł8raϤh�"���ęvn�;=<�����D�gE��q�ўÚ��`U�7x�t<z�	T�����楎�d�k�FK�a9N��iӻO~�+����n�]kxz��B���&��:ϑ�ccj˗�LjՅ�^S;S~n"Xiωn;ʬ�	f*�o�i�]�*��X]y�ݦ�2+ͧ}G�Z���k�{�9^��5Z�a5 �T5������$`pK�Tߤh��s�Y��y��/���yK���$b`CKK�@a��J	f�!~ڱ���L�~ܷ�4\c(�+ %}aƒ-�&e��0C~lx��vy�>X��z]�Q��iB�:������8�S%��h�ܟ��ԌFS/�@�yp�Cn���C:��1�j��X�F���Ľ1�.;9��w����X"'06\����2fѕ��W��e;��u��3�q\��i��ιd��ҳqJɥ��~=��H��S8Ga*�Add!R;�s*��q��������n�
�]<;+�[/Vp�p롻Ƹs����A2��燊'n��*[�Ĥ��B�9H{�y,���I���v���$�y��N�A�]�|Z�>�5K�#a��:{�mCƐ3FW\�N����u�hb�.��x�AVv�3;;�a�"r+�dD���+�R�͵�����=Rq>�^�DGSmwvY�ɵ�r�*�Z��� �$��I�=�e��ZA��S����6Zg�5��Ll�T�vv��b!|c������v��,<�"�Zz�]ZI�L�%nNû:��ݏFڸU�����|J��g�ҥ�A8Ð�����}dΛ��wj�=��R4��Ţ��5��G���`��B����/H96����>�I��iVI��7�Jck�ݦ�"��W���>��=W�}�7+k��L�|ba/FS1�+=~�!u$4�%��7|��,"�;��Zک;y{7�2�BM�}Z�I�H���+f����6H�}��������U�I�_�TI�~����*�9�:-���<w�7༩��M���ঝ��0QR�7%�WFG��dpo�����I�^�,�my;��s�t�KllFꆒ����&�m��xT�ʫ�-�!m(`lD\���x��ypU����kx�8|���~	N�c�D���p�V�f
��F� ?1��/�0�e,�#�>I��Nj�����u�Kܫ��O���d軓XS�uG�t�R�Ա�ʚ/ �	L���a�-{�^�)���n�Uo,5A�Jl�Q�H�m>S
����9��x��FM�)���������7=�5��`�(���g[�0ޮ�T��5H��=u�o�\(G#a�,�e�Ŷ�M8qۊ�=ny�[�ބ��f+2�x�'HZa&A��nHbnL��]�.��~<���0.�7�@ibek||o��Z�i
�ۓ|ʜB?��8wlշWU^���Ȅ`�0��}�Q��R���}�F]i��t�W�7@��Ѥ��-(e��j��,{���\�k0�G�ݾ�'լy�(q6B[�ډ�cnGy��k��8\v��'c��5�/}�6j/�F
��f�;��w�(p�o1�90�˹�鷘}(я��r󈍣����(�C��R��7ݮ�u�7�E�0�oKzm�Gguq�<��I�Z�#��K�����_�k�F��4UY;��u��1D� \ �to`��&-���!��䊚�* �޽�+�u=�	��Z�6�:{�:��D">u�;��מbܕ*!�VO���}��l����Q7\�<��-u����e�<�o$�ֹ�̫5|�E��(
w�[��>�cQ�w++e��<�H��2�B�@&w"����I~�,�r�<��Je�R�J� XV�!;g)�=��=����[p*��nx.p����C<��	C��c))����&��6�l��t��۩n�G��M϶�2I[u�{n��1�G8���`�X�Gh�h�6sqf#fL����cF����@Bh@����L.K��ͶR-؂��p]�e��f��E��7;:e�6��n�w2��	�Z��h�l��}w��q�(�.��n{V
�˩�ݓ<��]U���M�~&���X��mT~Kw�j}]Q�>I�n����h6�].��cl��/Ԋ=*u�����W��09@�o	 �M�0�=�BYɎܰ�?	�[��.�g-m!}���wWj��*��Y��P\5u]�|���e��})^�>��D���Q�11�B4��(����B�2����2�B�f����E�ה\�&���!^�Ò���T�]u	�zF��,/o����~�P12'Q*���)�wг�{G�^�Vz�@��ާ�aG�M��	�9��~��U�n��
�`ȣ���D�j�/fs�U�؞T[����Ґ�9*=��65\-�"N����W���hgyk�M
�+}ԪV�_�?z�l���(0��QyS������l��>�1ӺN9Ƥ�Ny��e��bk˺:�p,r���N�V���+�E5�$�/.k��؏��zv�_w�Uw�~ES��x�����$`���ū-�O�𙾵��v׭xOn���ta�k���dV�ئiN�;�;,f�56�FU<s���K��7�h�͎c�L^�¸'��gC�̂>�ߔɻ���=��I��}��o�'�JCa�{\���֎��%)��&R���PB���A��38�'\f_�����Ss���Ї(��jN���C"��Y͙��j��a�{�t�^vV�~�>D1i�ܒ0�qF�6n�֫W��� �� �m|Q�a���$,ۮ
{6m�Ͱ�r�tMøc7�.�K;W�К�Cn��A��[���&�-��Z6.c�ȧ�f���u
�Y(��x�����S�>��(o���3�^$����[�'l�Qc9�^�G�#G���/�#Q�˝���Qzx|v��,�E�l�͎�#���b0�J8IRH����<�~>t@��=Y{�9r$Ԓ���)Z�����!O����c��gQw՗�������#HD܆�$p��:�WZ7{�^��gm�5e\Y6yn��a�m�{�@�����+н��7�ۨ}j�����\v
�rE�"��Eʬ4)S�ݑ�����.ۭ�㔩��V�y�������$A�����D"P��10A�[g���7N�W���v�ut�L��m�B�_@��}b[[8p한������5��y������z$�G��ۺj*q\�\��E�xp���oX�P�;�R�7� �]�=�[����gN�vfn"K��9��뮝���(ۏ�D�&eA�Tɯ���b_�w|�j����l�OJږЊH�ّ%A��WF�M&�(��v9(�6��F����h�8-�H�7{���w����܉�-AC���/6�nZ������0:0'�[,kZ���yb27%C�|+5\�Ѹ�n�'��v�������ݡc�]����"��۔Ef��|rC�恬�P���U������וY΋۹���{�c�ئ>�R.��g;�Ɲ\�.��5x��`83*��;�ͨ�R�1d���rK�� �����ggvfM�FVJ}�WLF\.˔�zyn����A�����M�y=��������Ѣ��� {��N�i���aݧـA�g��E��sO�ў蹜*���um<�+�f�yR���D�k�[6��{�揍L�㬫�L�S���fQ��\kIeou﴾�i��k)��R� ���>/zl��Wb���;o�B�gZm3٫k 'Xr<�t�Ȫ��o;��=�]u0]�"����Hsu�uc5���Wu<�B�(eߔN��ǘ@��p����t�����=(\u:�s���E�9]iGHwu�hNʅn��������(�u��`��X�/̨�]�D&]�j�q+/䖾�#	4ێ?n�K|Z�}�و�6��'Lo#�[?P=W�B�dh��~�n��Oo�)�p�����٘+��L�>��ڧ"6#%� ��Wkث\��xz���� w�K���q�CJ��M��E_�t�j��ޛ����1iدCxeږ�u�^���_-���]�T1�c"�7l&��&I1�BbfZ�9�i�vzJ�p;[��E�6DMH�:����j�+d9AP`��F�=�_x$�лqYP��m���v�)�뮴�-ݽ_(r<���V;syhJ����n\F8���oi���Rwy���tgh7���@��[��뼀 F)�w��fd��^�x䵳˞��h�M���
?�FDb0$��z!����ʙ��A�o�z��5�k3ӕ�twF�V�G�rg��#��lY:��enxe�Wp�)��Uǿs爗��}��cׯ��V�ڷ������0�f_��l>9�~�^���[@�È#��O��dY-z)���(�[�̨Ė�%�N���0�m,=\�Q��>x̬9�}MҎND�T�mШW����EW�\E��峜ū0��DL̀�E�	(S����m@WSd��|r�0w"e��M�E짠�Kв��?x�����:�OW��_^��罰�)h-"���;p/���wL#���m��[�L�����l^c[C��g`'����]_o���o���\�����NG0m��Kwγ�Λ!�F��$��{�-БWI� �?�`X�p/ $n���TȦy�=r������>��ֽ��.~<�����~ٻΐ9�4P���M�#+��:Ŕ��ԅ����.��x���o˹U�n;�����wJ��>� J�AUmc���.4��8����n��{�43͘�NQqI ����e��η{��NN�	߭`��Eԭ����)ݎ�`a��޻��ݼ�u�`h?l]�΅�7��Ҟn�ݲ��:���ER��n�M�����[le���U���k����w�.Ɂ鎼㺙�햧N�-�#��C*�'��4GA��҄�#�O�pQ�N��\f�e0'���v�K8&�|�S�a��W�4��J�T%e��PO'+��
���w�sߣy�d���0����m˥k����s�6ƙ�V�\�1��7Jˑ�g�k[�>��<��v�')4��vYiw:�E��TmoFh�6�\q��y{K����{r�C�;="�y0^��ܵ�����`%�=�����U��w��F��l�:n0(�f��S�gr-�ciWY��\=N�'�=�=q�:ml�r��6�bba���p�G6�z�hqk���c�goᏑ����t�L|�f���"=�3>v��ݮ�VM՚8	�/��90?������;Μ�Yq���	��ڍ�a����ڃ������$�ub�T������q�҂I"�M�ߺ�H��/�X��;�)���A²��S�Pv�7���6��%.^�`�'�%'/�n�y��P��G�oW� �l3!P ��h���4i�v�I�^Aӽޭ���w]lЭnT�^4!X�zm��S�K'���_rb&��CR���-�Xz��oyN.���'�ps["��Ѝ�|�x�`�Vn� �חKy�a�ޭ�{����E]
 ��(5���t/��-4!��,�Y!N{�q4뻋�^w��Q]<�D���5����O	�/��b]�Ѣ���rs��#AW�?~/������eR�C��n��z�{lK��ᵻs�Ƅ���[xn�"���\y�ݕ�x����0��a�UP�BJ����r�G�n��g����|՗'pf�O�B�Nǅ[��>%Ĥ�l��5f�7%��j̀0z���OT�i�ў�ja���
H&�B�j�1��}7C��q �� ���KjS�O[=f�۝C����{�$���aI��
#�8��q�f���Ͻ����Ś3��~^ӗ��0�m@�e�Wy܄u]���������J�vǤ�O��M�k�Y�r�YI
 ��᛫ܲI�7�=��G:d0�t�H��ot���#(u{�C.�kC�T��<��PG*���;A��ƕ��S:Cu��ET?�|���/����wf�$P��Q3u�1YJ�ƻ!����]�W���ʙ~-���v 7jwuμդQ��'й���rZ\���]�`�JY=c���X2�����@���+t��S���f����n�t�D�#�[���
N��fȵ�[���ϔ�C7C���<���5��6B+�N�.��0t�t�����v檼�	p�P2"9�6�`՗����6j_\��j)o��3���{�� �.k��#6z�.����Y�W��|K��D(RkYA5#� �q��v�e�/��t�%�Z���r�9h[����բ�nZ<�����K����Oa8�k	��]�ݺw���%�SW:z�oc�2��ҏ0��Z
V���,t5lpi�����W�w�:��(#l�lbG�!)����o���Po]	���z��7�P���U���Q��%4�U�J��w[�X7ʆ�T��;sO��A3��$6�NF滳��ƶ�4H&���wG3�*Aӱ���1� �k�wz����>/^�����(��.��F����\j�Ř��m(tgϲ�?X�n�.Yv; Uw&�џ;#��y�u;/����-ZM���#�,4C -e�]���}��S����t��8ǦT�-�;��|y�(�ﯗNH�겁d=�QWy��˦oooǄi�&	RG�}�HFʩ��]����ͯ
n���~U��_-t�	$Cj��o��ڦ�\�Iqi���%�C������c�n4���l�tޱo+��7��{�UL]�2<���so=��=��w�Op��Z��v�Տ���'c���c~�s����5 ��qԞ�u�]T����{��d�(=�ɛ�yw�:7��u黯ݧ��g���ܐ�[*�Xy�;H��
^��3xh��f��ͷGy��`́�-`����8�w��Z��{�;��R����6�bu�sk#n�=u홡	�����v�ybL&Qt�4]_����XZ�Ä�O�pNK�1��Y�0P��m:�&������0f|-Oy7�-�7����͹�z�|bi.�l�h�Ie�F�XG������Ȯ���y	둂�\�%X��Pqv�nRi��u��&�r����	��?8NJ���5�k�����2.�a�+���v��b��oE�M��o��H&!'$��J�{��w{»�n�f�!J����B�X��}���+[��W��mӔG\	�z<T|"�6Jp�P�ᵸ��]�7ڍ��/!�A4<�R��8��_t&�v��F_��
	Z7
�����[��u����;S������*�)�����o�c��Jk�Hs z��������*5�;���E�a�~�mn��[�x��f�r@�v�F����S���\n�X4N4���kOۗ|����hnY�JީL����?vi�|0����zN&��4��w�:D��꜏]�6�>�0Ǜ}�7z��Ƚ�EJke^��i15:�Ƞۼ�k��n�7\�";�IF���5��&����f�G"l͎Ŝ���"���́)1��q)��%�����(F�i��ݡ��ϔf�rp�T[L"Oe�';ig���@(��d���m؅��hL�䲇F����b�3�RP��$��UP�L��1��1��m+l�5냓p��0�^2���1��;
�M�gYA!+v�ػp\7&Ϟ|GWM'~��s��Tt�f�Ƅ�Ù`1�6]7)jY�e�8��1��vY�,c���ܤټ���ͮ��g��zek��X�)�U�S����<}�>�����_�Q8�p{k�̡l_����F|��')ӸL>#}��7�c��@ҧ�N�D��<$�"Fԁ^�l�u~9垇~��h��9�v�R@z�^����'x]5��r��,�iyM��L���[����Nc�����JQ�nI���H��+�1d��r�G\��/�j�`#M�;�ӭ�G7w�,�Xe�
�u;�x�kQ]�0�(6>t�)��5��L~��vYg�����<��o�HI�K2��۶13:��D��ⰏU�(�c��:�̗�3ƩeAO
[XU�!q�Z�9��\3��������z�Z��,NxOE���Ѕ78�V����;��ǶuF׽oW�y��j}�~�����e%+�I/lR�i���ݲA�0zm5��΋{l�9 ��q`�����M��A�i�Bj&����P��/q�D\�Q�鐣�xɡG`dR��Û���7�[�%V{hx���3�}������z��j����7�^�ȥ������BWVe�n��K�Ǝ��
�1�1LNJ�{%��jh�t��֡���3����FN�)-���^����NAj�e�T���^q'��E��+�R?]��f���:��+�V��{f_��� ��PM�����:<�2��cX�d;V��|�{ҹom+����:|��[���!�٣�%Kɕ�0���./�A��P�bj�D�Y�\�oE��u�w\�MLwy^���dtb�VF�P^�c�z�����z��ٜ���\�N�!.coteuʷ�:;H&SH�D����~�a�I����]�c�Fjw�z#�J����h������%�o��1�T	_���o�����[�ht���_@���咁��l��[�6�ɱ�6q%�#�;h:	�m�a�V��i���	�����R23�MJ/��ɯv���u��E3�'ӯ����{R��n���ʟ1^����gRnc������mF!�E$�cW�&�y�������N��h�Q�G�%WKw�R�t�(Խ�=���ܦ%4ί6��wn*~��!�n �v�ACO�q�ְ�J:HO��&�3��FaK��/����9{��"$�盾�w&�������۽mEK$�P���J���Ѯ}�#z�O�Ԯ�h&Az={�.,�&�f��),�l2�%`�f*����O<�JS5�j���h6R�Ё)iÖBUT�"{�AG<̻4m}~����c�3�0F��{���w{g��^�l,s�*��ir��@�]�c�e{ĬN�t�#*7��8�Om��]<����ͺE������N\}���DOI�;�ƈ�J+��{�Ļ>�������%2!IZ�Q
4���G����$Z`���LgU�3j� w�kl���v�u�b��I!.#�'q3���}*��չ������믒*���'���~�Cd8z���)���K�U���q��U�����)�RJ��%U1��WY�<2����[�Ѫ�䃣�n���ڌ�xD��Vg�Ǯ����N�h��KW���Y�Y�6�3!PȠe'���t��ȼmY&�,�����a'<ά5p{�ڜ�"��5�LW^J�ڳ���3@��09y�)0��[f8�+#��o�{��xg|�u߯%��
q]��-��a��>W��g#��)�^G c���������̝�As��-t��� aj� r�W>l�䪕f�Z,�0GsPf�t9��X��:.ak����h�\�����ʟIҫ}��=��?0G�|<�)x�R.���7�u-�)Կo���lU3�5t��B��~>��7��b��wfX���
��j���A�wU�+���ʴ0�6[���X��c��Z�S@{ckc�1=����ŗ��������֙�w�(:�ҩj��>=�������ٜ�&��F��k�}Yb,7���VQJ�k�c&����U�^_��k� ���uy����7�߉����񒽵�Už�w�������w����uЇE�F��U��te��v��f�B��uM���j6JP@Ӓ+�,��Q/w��K�m���Y��jM���6�#ʽ�~��-w��gXS^���U�B�V���"hf	*�����o�.<�6�I�yeoC�c�y�-�Dܬ��_yWh}=:�k}���~,?tu��n3�D�6�!�W�/q���:O%j��e0�`�ʽ��S�ҏc�u���v����έǆ��%PA��[�q'Ef�靊����g|>�B���9���ɫ����}�v�Իy�ɺNus����ž�5d�}}�T�/��s�0��ٔx��>�X��7��ۘLQ\>�]Vd�{��HW�*p)H�X�YO�[�V<yM�����Uc(��:Ƨ������0^��z�6a��-��
7��r�t5�W�g�E̪ϙy3	�.�:�9�|^���>x�_�8�g����� uԵo+ߓ���skp־Lunm.�V;�;�kuR:.o%�^���؅�10V���%�	I=݅�m�0��8'h�^ij<)��xnl�Z����D����'�NO��/GǇ;}:ڬ����Xk7I��'��0��s��z�*���+4r�v+ѻ�En���.��b ��s*����Kr�Ǘ��x�6��ੱ��	x�8s(����R��T.%��n���m]*��.64ڡ�բ�3���1K����צ�ʩ�)24��%�-3��k��NC�ҷ��W|F�[q�T�!æ䌗���㽩.	dC���w�v����F�Ú���Pe�ڶl}p�1�;P��9�:�	�=���Y�7��z
�{i%��|M�%�mn��}prLQR���r[���r�6�,��D�{����6������멏�=dۺ��Fh7�&�z�iE�*�%=Ǜ*��N�Bעu��
����&�[���W��C�_>����Q��c �_@��Z�t�Av�4eZN���"��0��d�հ�T-둽{6��^�*hv]�;��il�Q����"�F�h�#�b.Ԍ١���� GJ��I�::ګ{W���3��F\���ps�x��@q/-K��ctB����v�Xጻ]�	q�9:#�z�'�b;\f�FU�����L97[.]���s.��b1ĺ`��NmѺ2f޼Z)V�h"���:l���j͊�q�Z˦��p�a(����-C-ˌ�B��tݫf�$�޴Y��mҮmU�C\��n5\���#�[������|�����r��Y0m�<�5vuļ=��܄^r� �2Jˋ��sb����ژ΋�����[�Y\���&K��tϘF�s�ݥG��m��]F�CDĮcJ̖�MF��\���0������m�q1�ڮ{B9wX0YF��l�A��.����F�be�ban�G�WHM�Y����&tIn"W�1�ܥr�
J]mF]t�f�FǗ���r!\v�<u�tuq�`c�v�
���y;o;��oBt���cl��n��yw�&5��&8��<9{��G;���݆�ޢ2ŏ>���q�ݎ�"����"\�Q>q�m�Jl6뛦|Nͱ�v��6�F=�N�����M�]�ǲ��vo^]�=����Mg����/-.nIΜ��������n�J)ܗf{H���n7ceN��Y�s�1R6��k	m�1s�gMez�s�fj5�J��s3
�K�z|�gcR��t�4�j��PcpC)w�>��%�m5a)�����&9w[H&d;b���x�G���K5.� Ѭ3afo4�Ғ��%�$n�ћc8�Cp��}��
q���೺��pu�]���N�
�JY(�.��f�.�K&f�v�Ȧ��f��l0� ��έ.k�V����r�s�b��t.N��<���v�M0[33b�ԋ�ŧ
<��SKe"^'k��8�<Z׸�.ۉ���F��+�鋴c]��B��=mhX�! �"�g3g7C�[4c�So%�������U����{r�C;6�^�o8��&�9;\����uWLܳe�eэ��#5��ıS�;G=���{{��ے�m#.T�^ҁdЩm���c)���,�7�s��r��*��EɢY74.ҪL�M1�Ec,�Ucl��6�E2n�-#;TU�`��lA�He�����y�@C��F��R؁�q(궰
ݸ��)��p�glJ�`����v���:�ۋf�щR9��i(t�]�nq��1�ʖ6m�f�ı'$����WEy��ՅQ�R��dK�\���N��h/Q���Z���<�c�w�Mqvh�F#�U:��"KdSjFR��6�E�Ur����z�k�}���P`C�ޫ
����	^��ֽ�vy�v鯬�Z�S"�`Cq.�|Л�@��#��lߤ�9/�^<��K��	ZM��v.Ǫ���{ܳ��)�y^� ���=�<�(��}�]�-8�A�ۊ�\v;xn��ud��%���EMVQ�{�H�,��sou�}Ƈ�@>�=�6g.�"�G>��fe-%!���@af(�q�}��TR�.��X�����OI�Skt�����$]Wv�W����J�~�ڰ4 v��,�}��Zx߽�}�;����TP˛rmi�4o�EY�-`�l��ݍS6zn�4'`KMU:t�6�Uܑx�¢�l���b��O\�W�.c�n��mҧ�T}���ǜ����tR�v���(K��`Ut������(@��#�;��m6�Uo,���6=*�������m�xi�������;3��ði�띢*��V�wF��-�+��u�.��pmdleԡ�kT���u���}�}ޡ�4<�'U|S�W�z�wm���W��k�@��+l��Ǩ�[���L���EE"���:w���u}᙭B���U�.�3���wk"�ܛ㜆Og���>7͝�Bq����h&K��fO!W�v�Ta��D������D�]=���)Bv���in����Ʌ0��ү��ܽ}h��"':i�P�y�W��Z�^Ã44����&v(�24�@�
LϬ�P6)����M��_���˗=ט0��^�/w���t�w^��* � �Y����=3����*a��{���7���f/L��͕t�i�8�rF�u;s�;Z��"N�gwk���$[��y�vE�Ko�wu�A�/f���H�)� �U�X�pZ�GW�_lW�J�C���p9��~�(�4��?�󌲑�'�N�}+c�m�����+���0�[}��̫R#�8��G��7M�y��R5�i=�L�H��4y���k6[`�"�@�`Q��(��U���͹�r�p�M�v��#������0I�펲z�{�\2P��`�Z�Gb>�k6��0�8lr��\uurF7^�1� �9��IP���T�_#��:�l��9yb�('�狰�0�`��-j����AR��t�wv��_k���>�xĦ���;ş@�i��S�!�>��)|xE�G(\��^�N�ef��E/J�R��� H�L�6��دE4���ל������k�
w��ׄ��B�~��QH���G��y^�$s:�ߥ|�ϵ̀B�(
�Q�6����7m�;�9	^7�ql�[v�4������r �wv�A�����'%V�4E`]��,��֜u��6��z�4|6��SU���L�E`�-��t|v |��V�����)/Ś��~��1S����T;/t�XTD󸼳�c�U��|��+�p3�2e�0z�:v�b����^Ҵ���L�|�R�q@����*"�2gx)u�;m�A�����Qg�Ѽd�[���_�ў�e=�(���S�Ny�X��x�B�ם����~,S��[��($پ�j���\U���T:!2ܮ��-R�H JM�@�ຜ�W�ʓ;η���}%��rH���B���n �e
��	a�(�4�"�L-6]�r4h.�w���ך� ;��@.���C'���$eˎVnv���z&w_	j�0/�rw*�L�||�:k�w�Y�V��[��*�;�)�D�O`J�~�����0kz�.�}�VqaU�h�!#���9�s�R�� ,�ǒ ��7)p�n�i�E��<��lr���v��n.6�=ӡ|�OJ�9v�mP]���Mm��z�l���>�x�T��n��han!������yw\jH�M���"���
���������=��ԍ�<��_P"�̊	�U�Go5Z�)���b��t2ܱ��D�6N\�{�y�"/��D@ې߼#��w+.�8+�.�5ޛ�nL��~?j���YM�.m�xV%��ep�8��߸U�^�Ap�ۄ��NOY��(���`�%�����Ϊ���f��Ǟ%�4�o�ݐ���U'�q:�����[���3HS��ݤ�ϐ!�dD؎��i?osx%��Z�E�&spר�J��6�g[��<o�yI���)�{p�vO��^O}�8VЪW���3�z
�܏]����T���O���Zv��aL��g�����mLu,z`wΉ��<��`[
��u9��Ycʔ����I���A1!t�B�6G�bO����a뒩�Hmj�;+cO�#\W��gsL��w���\;O<J�muvb�1�6��g�=t�Z�̲v�{sݮ_@\���!��:���!���w[`�MY6X�w^��9
\3)����oA�m8�n�6��qt��on6���U1�\��d�޻C�[��!�"Q���3fbR]3(s�Ӯs����g9�n�ؽm�x���v]��&5�V.�r�fj�խ�1�K�Li�2�g]31�p�b�@'qRL�w��y�4�ڮ�嗦��E8��w����+�Vz��*�?T(���K%�N�4��>��2?Hd��c,k�2�X��c�e�D��H��03x��`[\�tܩr�1	���y�[�^�ʧ5�=�����Ȋ\h�#�=�!�%C���¼�Ӵ��wf:���g�C� aHP<)�bΕݻ�G��e�+6�o1�RE�H���fˈ�Z���a�{�4U�ߦ�,���s�N�3���W�P���ӷ7�������Z�1�9�(�E�!
G����Y,"d��cR�d=%�3��j��)t���`ʭ�?s]B�N��Ǡ#�����ϧ�.�������.X�
U�jC[�4�V4�uj�#5L�`"�*1r8��i�'������ˣ���,ujit����@�Ol�yw���Yٶzj���#�
/��d���o�WrKRo�.��Ȕ%#�FrX�L���^�3���Go�$����g.���}{[��q��� ���J.�5Q[jөV�<-���Dl�xg
�I�if#SP�@٭��Fp�.wV��tq��Fi���ӟ���T0su�+��S�5~!-K
[��j���a";�P$C��p��B���;��9+��2�������&�����q�էv�{�[F�5v���EM������>�W��w�����X$�}E��W��޴+	�>�5oݡk�r.T�}k����0�-+��R�5���+�[�|�GU������$7�a��k4q(��#���u�J�������rN3�� 컕�=�C^��I*�P�����!������NX��k���l������I4�MuuLc[�j�Ij�5���-h�.l;F��:��+P��I8��9(aD;{~���!v�
H�՟U�k6V�R��*���	��]����Ԕ��*������3%���)H"n�b;�M��2��rS t�Uo��(�}ϙ���F�cd�]�q�ɋϘ�	���п3y�pA�ӱ��M�ފ���}ןF�&A���N/&o�{�7(��і�I��]��{%u�e+8E�B��ZZ�a�b�{��r�*]$uOd��� ]�B��:J2ҳV١0Q��E��7���[յ�F\���i��B�xc�>��.9��5���ˋ�NQ��2�BI���d@���Ew�����ީA؉^>ߩ����\}T&�|-�!^B����]X
+
��+�z������>�XF�=75)+��L@�fC#9+誊�o�1f7�P8!�^��h�Vn��T�~�(w��\r�M7�[�)�I�g wUT�ޜ��޼g�^�YF�m� �V:8j��F}����n�F*s��h��3�s*�jE��Y #e�f��VZ���
��m\$n�o�d�����(�R�3���mMyxڣ�Z����D��	��B܍��1FT��C�	P{z��,� +#>z�+��¾�B�,�����b*1��t�f�8�������z:K-tl0 n8�Õy⻝���ɯYnjBe��)^��[���-^a�W^���*[`ţ/�ˮ,�������unﲚ�d���ڌ�T�\��O���}<���q�`�\�z��R5V�%�F���7���U����Bl���s�9�EM�}}݌�*�r̚kzW��[6��1wh�9��;v4i��,���qve�:��_�YF�V���߳pZ��c�$�e��0y��'|�/$�Z��-Pr��x�l��!���ЬA�� ���N׻_SsIu�|3��΍�Bi�D k�=O�&8�m��B�6�ş1Ƥg{#�&�\�YF7c	r�Y~��_?k=_~p���xNͿD�א|�ə�)�ar>��>���:G*|'�no��Ec�k9g����h��m@�*I)�}��ʚ��
�t��ӎ�z����-�=^wpqf*��ms�((�rtm
�J�}��?L�c��݆n#���*1=	���Bc"I%ߗ̹�M����<\�f�T��m�!�W���􎳧��ea��υ�xo͏vV5Ǹ�6qt��$L")��/m]֌������V������@@۰`��(����'��y�&ȦG�^^~��nӭ����i�k؄�_>y��2�!��N_ y�ܟ�/Y�x�Q[]�ʸ����ψzŽ��^��q��ecs}�9ૅ*^����r��u�W]�;|��l�t�<��w7�^����4�wh\�������l�4
����X�Vڡ�]��zfu���nc}��7bs*\��0)	�h�͗���7ײ�^��;�B�s��۷I0�q�M�.t���Z��5B���GK�i�^�;���s��с8��)��:�� <S��W����M�<j8p��'j�y}:#��]����Zz.d��4��a���:Fv��d��Ƭ]"l�s��»��nMۂ�i�v��nR8���7��}��;m���c��w+��%H������ �;���]���k!��	�"�A��m���k}$�
��;*O��r��kޤ����Eڪ�K�@���z^=�����V�ӠY�KU�~�B�Gq�\�qX�e4��T���9�e�W��c��՗�T�V���˟y�L+��u�=�3���3kn�6}�Wh[�]%{� wȖ�QD1�nn�],VS�}CU_z=�N�����n����x���zJ��[�b�P�v�)苧��+�mk����n�A�SN�L��������７�ZW�.���AM?x��� �2wu�����}0od���.��v2n}<�i�Am��e0>��[��g���x���jV|���=�hLTz�u�-��<]�p����{��{��^q�<�������>#���?�l�u3j놗��Ɓ�-ۖp�w+�]��w5����m�V�3�p�^m|��<B��>�&y˒��� �X���?]���a��1����Y�es��y��͏X�W��Z��E��<�d��)�،V�	A�2I����bW3 �B�=�=F�Ҽ���<�d��������N�(��m�)�;�]j���5� �t�pޝ�����źV���G��DL^5���f�s�yE���mǱ�W���q��|_(�����Zy��""KqH����,�j��%D�,�0(�jC�!�^Wu�S^:���J����Ы��j:�.���lh9�>���%�- �-�q����re��-���sű�%-`�oN�Ig&�^^�=k�<�+���xY��U){����$E>:B���m�!D�}���ǳ�DAZ/lr(���v��eHnzpޘ�ӯ��W�w���FϜ5���d�����>�~�f�ۏ�\����H(�	M�hEz���C�q�&�7dm؝�a*m\m-�D�JI%N�x�e�y]{ǧ]�kF���5���u3�h��D��p�I��n���4(}�ѳ��_�p�]pň�>B�!G$6%��*ERo�U�֤���7�AD_,+'����>Y�8r��c*B=[�5e�L��ߎ���0��K*�v��l�	 ZDB�u�w�qlG���X!ȪC�w��3����wP�!�;�D���t�}F��qy��QzgN8b{�R�
��Y�%�;k%B�("Nhӗb�Ȫ}�Ld홠Z�:�F��pY��]����a�z����r���m_Ի��r���qFm%5fZ�SAuo���\��ü�2��Z�2�mnb��*Ϋ��V^�����գw+oY{���n,���
m��\yjWu׀�]psNaˋG�G
�!���x�"S�7g$4q����Ɂ$s�7wY��"tO�*�h.�oJuk'v�'X��@�\ś�8�C���Y�wM�Dhf7Cxśu�hD�M�����6��a0�=&�� �6�o �ːn�=��Fm2oU�XwH�(�"xx�E	��&�ŕ�:�z\ a$�᳧n��T�E+��ܢ^c6�5K7��`�[x�ԧ��l���H����qZ�FibL��CwB���7k�-ЏV5��������C�w(�m����S��yGl�Y�t��-,�A��#M��u��S8�.r��{��Q�zv?�E*�:3em��/&J��VJ���]���ZJ��/@����T� O����5�8��7{�4�Cg�F�pi���蛸�A�X�U�'��-6��92�/�+3b!a�"P���s([�O��s	��hd�2W�����Q(hn��T�E	r����(Z�!Yv��B�X�(>P�ʏ�[�����:#�կ�{�Ղ�&���n�صz	ļ�5�@�^:�s:.�{|7`[�[�N�.���Yؘ�b�b⢮��*���ܩh�yo*W���kߖ�(�m��ch����c�VQ �+7���ܻ���Lz���!�#E�	���l/w�G*9c}��ט3�/�VN#�?^�']�qôs���VP�#��Ӷ�ͨ%hE]���M�t3շCs�78z�ch�
B�,�_x�u��o����)�&��X:���vA6nx�\<%?Ed��u��s�n#c��x]�;��ח]�+&���<�Ǆ����8;x���*9Krgs����r��=��<���Z��X2ʗ@#�bJI5��⮫&f����)W��o�^�G7<W��aȂY������ѽ���쪴Q;�sۂD$� ���a�`�Ex<qz��&g��&���h�׀L�����i�d��:3<�w*��1Y4��>/�k��q��g=�C�]N�c#𦟂p6��d�卲(�%�N��^��x
K�&آ��WҊ .5�1��,��Ru�ADD&e	�Z��3R�G/:-E�u^����\wo/�-�N\�V=LV��W�w=��j%�d��x�Y�"�e��T�m�s�A���G1h�%Z�J�X�L�e� #9���u�����=�Zw����8I{1�	}�S<��7u���z� �Q�\K��QCN�� �C^��3��8��V]�Bn� ��G�KV*�7o��-�0fU���59n�F:�C��gJ�Jl.��4�"[0JB[ �a5��21�6b@�sV�u1١s�D���O�m`��.�pW�!V���#�6����e<����ľ�\�����~.՜O����S�J�������܌)�ɸ;Ov�>��ԛ��o8,$�}0z�maX�Z/zxn��&����%��Ć5��x��.�F��HJIH��eQ�n��zK�O+�X�߱��g�oj«`U�}nC-�����39�![��y>�B"�|�}>��xR{���t�LUmw&���FK����:}��4��kqяO&Cr�]��I[�M��� D�9	�.eNa���r?K�m�#(ܦ!nV8�N�Iu�&omLa�gE�
/�^cν�<!��˥p���ca�﮴&A��o��Cn�/2�ITM�4�`�����
ٹ�eG��N��[;�M<7���*i֟'n��ɒa��U��B{�;O����Zoy�5��Z!�lˢ���F����m�V*s��;p�헺E-��6�NM�Yx�Lg<�NsY{-�z�;(v�g��#J���r�Ÿ{b�d���q�;B��-�9���8�-�v4i��Y���g$fWMeP�^����lGmxlh�!�V�H���{f��8Z��)ͳ�LgS��ҽVs������5N!88�Լ�/�;ew��M5u�K�4Tlg`�`�����R��M�	k3(���,���%'����>}��m�2ȷT����+y/:�^zBk���n���˫h�X�?z	l�7�u)P,����NsL�ـ��n���OJ�N�̩�3Ҕ�=�7��p���AG��θ��>�;*�vX�Z����r�����Up%J��	 �r��P��|��`j#�!�}7L��nh[��eK���B�h(��g��s��0�㳏�}���u�P=1�I$ MO��DM�iZ�Z�ؼ<��uwFT\��9X��+��.������27k�[�g{=wW��8{(�W��bD��W�f��x1!D���rdJk�%P���Ša��3��(Z��.�o�T�o/�z��� ��]�Y"u�eЅZ�@���R����FAnR���a�cK���0n������r8ni2��fAF�]��*�p��	î�ȸ3�z�EE�Eܯó���į��wf�g>�h7~�>���T�l0V�C�CQ�e��M�Y�P�xu��L�/O�,�Fo��jƇ.���wd�;h�rP���u������!9S�	� �H��	������klN1�S�Uko�&��B�GA�A�Z��������^��R����G��i��J�.�{>>8Ca�����;�����$�[~e��쨪3�(��UM��˖J�͜@�'��4�4
/ޮ�p����4
m{4C{q2�zyzk=�{�՛�4��j�=���r{v�v�x`�q�&�'Kn��#�9���N���߱�l]����D �J���uw~������p�x#��0+B��������77:xO�}IЛ����1:_�[���t�%M���3VOw�]L�,�m%!���Cq���W2���w65�w!v�6�i��M�7L�DbV�r��sA��yZ�������:)�w�G{V�q�ƻ�<��W��0���=�l05,��W?!y��5�}�G�D&��e�����ùxS[�}�+ܷC�<(ڕ�������Y)#F��Hv��W: ��s����-43;�΍ƪ#�����2�M��E$~�H��33�{8>#.t�Qxtu�	A?b�*��5�@vs1J̝5S��R����.��0:T'@_p��ܫӓt��k-q�]�G�Yd��/�iɋH��Trd��Hf�ނ��Hf��Ļ�%�,:%Ģ�+!��\k޲�\�N2�
F�1X�u��+�������#���L����h\7�� ̳[�9g�)��>��y�=YjK���*���X�<�[Bj9$���!��'�˅��-�Weճ-���c�o��!51C.��������/W����l0W�`L#;�0�h]mIO�[�3u.�1�r���>	�t{�����dӒ��؇6xx���6;�~7ݾ|i����*����*<�)��v����ql�\GCb�#��#��w�^�W�Ԑ�U^�4?�|i��I0Rq=�D��wf�=��˲���캀�Y,[F�K�u�[�a��
(��8�^�5���n,@W^�ڻ�����<�� b03W/v=7C=0�{�X!V1ēW@���=U��;6�CoN���Z�ߪe����e��Ff&����$FaHDL�u�0�`��`�.�`}=����8
Y]�:�[	��nt���Ih��43�#�L�β�ˏr\��KSV������v-�u.�1�$?_n단�a9�\9̪�&p?I���4rd����9W����Z�qn	�Y$�IB��������O]�W�4�F��-wv�/�k6��_�9�5�KJ���YT*0��Qlz w�D�Q-��&MF6�2*�6�*T.�C����p茥�%�VpN$rۋ|Mmת�ɣ���κ�Z���Ы�A;#]t��2�+̣$�`��~w�7���k�]�g��IY��F4�0g�ϵ�"3B����-�݌,Nq̢��0S|o�y�������S}m�J��b(��}h�	}�%L,�>�")�*jF�dBJ� �󾜮��~�M�3��Y�IK^��&�ܻhV�(p��
r_T;����XYg�R���{�]`���Z��Ir;)�X�6���������ێ��]%{(Z�x��A���e[hn�Qmmɂ�f��>'�Xb����b��G>(2�H)�)�`�ۖ�壕�4��2}�K7�{��m��t�GI�"�:�O�!��M���+�J/�z����n��{\�1>��˺t*��ڽ�����%�v	6�T�:O]�*a(:�[���ۻ�B�X���c�5���}���w�T,��@�L#�.�W8��+�7n�.����8�<0/Uǂn��#��ena�,o\l#���4f�l$�u9Y�,]	�%��`��	J�]1mI.��o#[�h�+N�5���,��i- iCv5Ƶ�U��<�j��]enn� Ҳ�Z�٠<�Kn��N��M���+g�^�����\&���n3���b�8}��9{	��׳kj6;h@9�yB[�6�K�.��Mk�bcsJ�D+��i4ecl3|���>�|)y��K���ez����w���*���}Z��S�`��a�/I�%L�V���/*������&�D�:/}^T�er��x{I��Q�v�::v=`Y�.�:�9�)xoM1l*�u�/0��;��������2�x����N1h�${����jciv7��� 4e��Cܦ���d�Y�[8�� u��؉5���+w�
�9A�f��4�U��	!���8�4��[�����y�q�[�۾0j�'+Wc���v��S���v<��%%`��o#"6)�Ŧ�O ���E{cd��b!��  �f��3��5F)\���Uޭ�ɘ$���We����'K�X�Ln�z�񻅇��S��pos��d�]�����Z�ȼ�n挽y4��鲼���[�r��<C���5����h�Ut���'���(ҡ��<��Xy�i�yn������]=Q]ӏ������>F��픕�ѱ�ɥ�h|�#��(��L�{t�aU���i��-��ʐ`������~W�#xM�0n�x�g�8�p-9oEx��d�������sΥ�	$k^���	�~�j��>��`��~Wc�R�3� �S��JV9xێV{�ֆ}�|/���F��N݉'g=��:�,7A6\�6腽èz�8��%G3;Ҟ�d���Xtɞ�/(n]Zkܽ|�c���\�gO�)
RE	qAg��WY�^meyb7V�#-��v��.Y�[�ܾ��0֗s��C��
��9�3�^Ckv̏|����v�[8ST$!�a@�J:�2�����].xŉf�o�L��,̛�Ŏ£>�1'K\�7��^�����i� ���ْ�z�E�LL}nx��m�] )�[���_<�ɢ2��]�ɍT-���ae�-WPS:����|�넮5FW��2�8l�Su�ς�^n5��݂+��r:i7��\r)*Ӓ_��ʔ`�B�Eq,��L�"�E$w�!�����,�<Ξ�vN�*��L���YDs-U�M��U��/��k��qmܵ�
+|���m�S���^B��aEEѸ�ML��{�梜�{��e]N�`ު�_�n4�i��f�G5	��Lg�ne�Y�����}�N|o;@˫�2�K�Зf�d�2�����DA�è���*1�T�\�z[A^{��KF+�`{���߰�e4���]�(B@�M�,2]�]N�48)��ǧ�f����L���8�*���L�S��m�cŬ ^�3b���6U�~D)4f��d$_ ���)��ф׺��*�a��QCק}�V.J�^��lX7�O<�#�0ш*�]��wYVh���ۢw/M�{��=d�<`��j4!���m�0O6��x��b�����HF��V JlO�R>�J��ˮ�/��{u�v3^̛�]���a��|��%3v��.)��r����⓮S{i��
���&�����!�G�Vc�=������Z���d��W�g۩�t&���m9�y�3��콮� ]_/z��^�k��j?=g��<��a��ѢE�i�L���V�S~^.ƭ=���D"H)Wt5of�O�״<=K��B���]7o]��Wo��gFpM�H�a��I*M7��D��.��W_�4x��''��;������Ԍ!ה�p�y=�{������Sx��d_w6��k���K�&�JQ��?E��m_k��y�4�e�\.�u.��i�t8�v�s/wq�;;Ɂ�Jw=N$�MHp���֔���[��Й�6N���)z������Ne�M2�/m��͋���S�Qk��&v��:�^��׭��,��A�ܦ��&�3��1��uvsyG���nRQ<��YyܶQ�.2�*��4#a��A*2���F�t���BU8�K�R`H�Hҋ��f�a�=f��o�.T��>����@���a�р�/g\F���k�WT����Q��I{��"��=n��<j6ҧ�򡝀hG�A���;�����)
B�f@A%$����˄�o�u���ۨ����/5!�*+�fb9���n��P�s/����<��E���YP�޸ܒ�\����`�Oi}�7�{8������#��+�8K�'�ճ:w�l�!���ݮٚG)�+9N�d����)jP6R��M�8�����[A�Z���+�����$����x�Aa�9`�ƣ�������/�����{��4iآ�fp�������.�#*S�_)���״sqob�8���Tv�"	�����_nt�)G�G}e�m�1�ֈٝWJ�]Ε��WeaK�k9(gat����14�g8Ouu�w���61-�(}�>2��(õ���wJ��=͜�vuY��*(7�*�W8F��y�a�Y�q�e�[)�ً�����*u�IM�;sWt��\��E�B�2��F����YW+�Ei1$��;\��U���{)yN2�ֻ@�H�����*am,8/Tj��S��e��-n
t�ܸ�ɾҀ)�:��V�G/�������w|�V��!N�F��w[`EVsQ[Gr�tz���s�k5�;I���oX�J�߮�
���	cgMA|�֎����i;*��X��٢�|N���3�;b[�z���n\�9�Y�D
�ƽ�׺����Nwv�������2�_�����6�)\������͑�T�V�.��::��� պU+&�_ْIH�p4�co �m+ٺl��8K�l�n7�ʪ�1�)եĭ���u���]������)5�`�F-I��Us]+W�C�`��������v�n���j"6_TY�����
����$��Œ��N�ۯ
���M�X��	����7n���w���ϖZKM6b�f�%*Jq:Ђ���N�z}�v�+4����D��%��>#l��e�v�"Y�b�(aw�����ϳkp]og;�ۮ���*n�jGh������F'k�{p*�k �������`��I�h�;�R�7��t��{���<�7kw��0a��B�:4�?L������;��2���kd��$6����h������r��s���;U�qh�L���ծ�d��Y-�Nq*���g�M5҂��뽷KW�7��.�\�p�x�3<4&B75n�5hK61(s!��a�Mfe!&N�¶�*�O;�8j�n6E���3���uP^:�5�d�f�+�V�Lj�PL����]1��Q͗g�o.�x냫���Gi�rZf���rj�-���r�vRۄݷ&�> Ls=� /-v�8ќ�6n��<��ût�;x�:���ua`�e[��n�c�;L��)K�e�8��UݕC����>z�A����;3��:��n�ςB@f�����Uq�8��y;5�]u�	G��\9��<�)�]�'�I63�W="�3s���mȸH�j��Җh�ꃶ���7A���Y�%����%��;��8�L6�wlC�����wT2�MU�Џ����5n��%�y�GV<�T���ݝ�ռ^�^#����ʁk���v�� n��랖�Wn����zk��8���8�l�������ٖ���׏V+m�M�^�k][38�x,��c�V`����;�Ms�ttn.�\��I]�x{��8q��^���Oi�-��wf陹h�[[�ݠ�u"����٬�,tLncK�t#-�N滞��;9ܻ��^	\�7;{��ə6��V��۶�%A6���-	� E�'lt���x��Jd JR��R3'\<�;��f�]��ϙ$89���(:c�ɰr�v��DG<�6ޝq��n���D�f�B9��8�z�Km�q5�k������Bls�"��%���� 9e4���t�ޚ�z�]�q�RV.�㦠��7nz[�݀�v2��L�F�k��N�&�+�r��q\�f�a�u���܍0ƶ++LL�G�g�5l����$��C�^l�Fgi��A��&�mb�l��&G��m<s*^��qY��<.�e��S<��&E�@�7r��Y�G��wN.�5X�GdR6���` d��j �6V2T�3�2!	�S�`���=������v��y�B�)��Gh�&�m�I.ж�y�,�{�c�;a�6}k�������n��3
َhVh���oF�m�i�a�c%dr�L.��^����^v�[�]�w���B�݃r�]�;n�r����϶�E�6糎�����v"�˳�+�;uM�L��˘-�t������ޏK��|<ҕ�EZ5��gA�'�j��E{kηsݕ�<��{,�y�R���lz�5H{N[mp��L�Hd�xi\H�����L��Լ]�tK{ O/��p��*cK��K��zL]ʪ1��}~�:K~񧯗j�s�/I��2�-�!r;�+��{w�>YJ3v��A��16�-�=��ޞ�1}�m��;ő!/Hm�S�8�|YE6�N4�qb>A<�~�t�0�~u��,9�wD9�����TV� ܛ���]6���C�f��ⰷ���մ/�.i蓐1b'!N3Y��W��av�K��i<���m W�nnO]�VO,F����f �t|���0����M��+�1��x߰�`��M��9�[֣����he�Mn*Q�6(��1�3��$�S��$6!$����m�ׯ�'�;�ԥ�-��o��m^�|���ym؇ȓ������1o�q�ٍ������t�%��&�Q(�5$��a}&֮�'O{��ܥ�jx����r/X�=X0���&��Ne�p��fnu�<Ou%>,d��Nd
�;8�����r���6�kT�i&����tX>�=�j"��[�1]�/$��n�ζ��ڲ�9ӻ��
��ڥ~��(�A�-�M6K`]��ɸ
﯆I�;إ�P�sz	��;<&�W+;q��U�L���t�N_��cS��4��V�d
�E�����j��|X��֡����7��`���i�L�\�V}�w���u(���q�c�)�~ǅ^�΂O�jT��\rU�i�= m�J�h{��]7��{��}I.3 �`a{���;�<�3�&[�9�5�#t��x�:^%\,i��#���M�������)`�c��E`2�� ¦�ЁF\�'"�!%��K�T_u�ճ�*�)?
kM�/F�۲7*gx��|N2��7w
s��U	�����LD�f��%��f��V�qɞ;N)��U����f���򉄄�$�)�\9��u��==��^I����/�K�<�|�(1�"�.�� A7��U�W'Xi��^����)D�/$�7{H;b��ͺ��9C&V�ϵ�m�V�s����X��T��(�����ܾ"��3x�X�R^��^��w�V�������O%q>�H��N�_pa�!�D'褝�$��`�����������ޖ�zw�{*�q}�����;���D��f�zա�z��Owj�h���d��pD��n�u����TM�ҫ}��{%�>���'@\˚�y�B��������kE�T]�]�P^�������c�a	��KQ��a	
ң��m�Aq� �H��ڊl���*G��µȣ�=�ڪr�MF�N�wz�3y�
��yw2�g0�I���ڏ��6���<d�fHm��V�qa���s�o��|�b�*�|�Kgq�\����(/{ܩ*Z���J�-Sz�`=E��㻭�I\ɓm&i���a0[^��J�/��ڹ��\���Z�c9��`XI[0^t*��-�\w���41?����c"�=�
6�H�&�m0d̂T�M<�G�//z7��7uY����h����5S�^�Ծ[�a�^}7���:akF�9�y�h�R�0�P �b���؟4/�],����r��5�R����79��9�f�후��z^�ڤUi�_]vI��y� ��x��T;yS�"&H�I� �/���V��W�����5�d�ҭ�${���Բ���Rߞ=.�������\0f������=�zr_�oך֚�n"������Q����:�c:�1]��f�03A�4bU$2E��ۏ�#$�ɚC��o����'͆k&w��b񶬥�}Y��o�v�L�
ϧ�V�E�	�(��9�QEk�������g������YH��g,1�|^e����ciN������ ��J��y��V~��}��%A���o=R��Ar1D�j�N%"�dK[)=�~���uN���YX׭S˛�91��q�J��B��J�{�PX���O���x�D�v߸1a(	�($e�W�C�C��-�
n�R��C���,R}�]��fǓ�����J�6����<v;��W����nX��T&-�($�h�Ф�N��I�oi��C����"i�X�Z5���X�
@�)֠l���u�����j�e�m���mc��Zu�z�6�����9r\�^��/+>{��9��p^�Ș�T�WJ��*���m.�L#�w�|�����\�����i��b�}�7�^�l���ނ�p���ƀ�Й��cf�us�ӑqork����`U�n�����@lH9*��n��L�bɕ����ۊ��]�cT�գI�cAX��֛\ql�痉����'��v��u��.��g�b��W=z�E�nv��o�����3���v¥�34ҋ��]a��M.�<�Զ�i[�J׮�ʥ�Y\A�Qҕ��z�ۋ))Fsj.�r:�.^VC(ܠx�/�Ē::�Z�0�k�4;�Rl�����1�!$����͵������{;Ew���y�X������du�aPA�@�Ŝ��l�e����^���"�!1A�H��QiL���`���7�!�ؘ�����8�X�Z^�~@ɼ�]�{Ҷ�
�T�����27iA�B�m6Ct	�dn'5�=�ʒ�V�NI������^��xw1�0���i_z	����a/)��F>hb�9C����h��m���Z�uv�{mg���ni^I�__d�7�(�s�SƦ�+�mp״�ϵg^�P��|ɠ��v���,��̅����L%����+��:�7'�b�V3jOX9���<�)�"sٶ�7��Áfy?Q�$�{O&?a�����kf"��%Yi�8��� \�#.{�HW,�s��\��Js�^�Ik�5�1̄����28p�t�ܛ��t�|�к������Jv�F��uj���h�t�׼67A��u?]�X(ϙR"�N/[��r����dw=}�"����~�g��>�Z���#
�|V�g�e��ˮ���݀����»#_i�t���a�`�:9���v��ә�<fj�Xd�͍�^�}�����y�;��v�G��A�xU@��wxX��y�v��J���<�jX�1䄈�EI#P�	���.f�O�g�B)}�zqJ�)\H�v��ϱٽ�iש���_�Ԭ���0�n?Y���v��������}�}n���d�t���Z�,ɓ}�5�t�"�P��DT�Z/���8�Z[�l#os/#�)�<��v�F�NI�4�w��Ao�LN��f�����&
���:�,j�z#�I�����r��PN�~1E���3�M��>��*��� [�,3Z�Rh�@�bV��`����fF���f�G��b�-B�1���]̾������Oz?^ȴn@����s��\7�97G)�{���Y�m�۫���aV��T]0b_���������mXn� �۽���A��Z���M�{
�e1�홷�`���x`O���3�������!�-9,��2��ɮ�}eS*n��a����ц�u! �����ӻC�iȂ���7��r4^֐��C�����h����t��o0�_R��N�voS�'_6�s�rvXr���`]�Q�ǯ.T��n�i�4�,ϒ�B26(nk1���L���;W^D���Kg��o�X,��I�~�T�����W��i�접$���{I<HJ �q�pAx���މݯ)F=�h��Z��X}@漰{�Ȏ�Je���lG;93}�:`�Ul��2�?q����nD���'�d�h�Ճ,��)]�.2��}l��XypnɌO�ɻM|fpe^�ق�Y��V�9.6�ߌ��5{ץ;�}:����35H���V} �g}�B|3M�Yr�ǲ��b��H�,�	3�8��!��� C^���e֏����On��/���-��_�p��댘\%os�'M�@�5z������n��ې�B�98'�C~��qp�_z3̦�v�g��R��V�>���P@��doHf:`�����ۼ;w�My����� �(��MYڋ�ܧb���w�7ln�Ss����{��G�e)����Q=/��vھa	�儋=���HG���\f��גƉA�ۘ$n�ͭ���p��K�cGZ�Y��]����s�fЮ�L�]�*@H(�-�����up���(�%�C��2x/��BІB[���Tm�'�zP��l7��ӥmq����}ww�5W�_��"�E���i���ӺC�Xp��-���a�2�ť��]���`���	��reG�.Ǵ+l��l��'2eI��^��|���xЧ�O��n���	p{Ƨ�L�D��s��>&�_��[&�GȽ��!��mp8I�Ѡ[dO�Qȳ%��j�����<�g��ˇ����_z��xxO&|�i�s��$�8����a��r{��}̤v�ځ�a�&�n��2��^<��W����P�<q�6�Qt�0����N������e��9^Y�V����t~l��BH���Zf���wC��&���ޜ�F��?[��ʍػ�}t��E9j(����&1��2g��V/�����i��N6dA�" �$��RN�ל�X����<�T��ۗG\T�����7�A6�u�.���F��~p]��D*��*����(.�j�a�й��� �y�X��B�����m�R��ø
�i(�E�͡Pk��Et�·p�7�/�w��Xx�;��� ˭�̽[���A.:� uM�r���	��+���͹�suSl��1�qm��۷k�C�$����kmo9rK�9i��f��sH��Ҷ3�]<��vv�|f9΃��h��[K�̭�s�xS;%7j�0ml�1�ۇx��V�]l��RSXJ�$0gh]��x
8�6kXu���c����NL U��M��@vn;�;ɲd�����#�]��&(���u��h�����Z�����l�m����и�@��H��I��R#����o�?�-<����?�xbL���[�W�_�I���'F����5ЕV�$��1wtS�!ci�>`��p�R߹��Q���p7�k�k�vӞ��B��2w��a����D����=��P�~���Y��<�u�j#մx���|X�E
(�lg��6�!�.h�O�tp���G��=u ��wC������0`�㙗����[�Dj�/���D5$0�ue}��SWZ�ok�ٕ��0`8ԉh�8�k�N�J�nd6��с�>z���J�D�x��������MYZ��<�Ȋ�Ɍ�"^�k��볖��<�@�8��ʞG���ޞ�'W�{`����:�'�v١�P����f���%E��p6�IK�g�����{:ц�k������a�r�҄`Mi��nA2޽-�S��2�ut�\�V��^m��%v�+Gs%��~�֛u�ך�����W����C.�`$G4�9�����+���7FxVgE	Rh�kfqbGhgs�԰E���lm���f�%vYoz��;8��M
�Lh�7�jf�erg�g^��t�F^_gK�|v��U��t�9��879���S���������h����3DoǛ��
E&%#��R�ƞo8���V�66���l�{7��M��d�u/>��ՕӺn.�h�e�B_
0K��$($s2��/��2�����c���,��A�Fu
�ʯS�a]�s�����,�{�Ow'�nҽu����p\d)N{�^�h]�~S`uw�#�/wN�^�gF�+�q6�&X�h�9�m�ٟ6*{.�Z�Dz4��IdV�pŔ��"sݤ�7�y�n��I���Hu3M^������&�7����$h,(g�2�����F,�U�*�k�Z����:�Z��^]絬��{f^?sqj������e�3��)0�_ľs-&"qD\����ztU]R7f�����=uݶ�[�(A��>�M�]M�����^ޔ�o=�^�x1M\JW����Ђd���iH�7Z��8_�?2m�[�2��Z���;r��u`��U���Mm散�:x.���}[&���۟M�����5��ܡ,��ow�]�x� �{!9�u� �[�|l���;�3��A��
�Gi���\gP�{91BE�:� 9Vn��C�wu�F����t�ʳkL�00J����:�rQ9J�9�׻b`MDӴ�n-#`�[�񑬹���_˝�O�ӊC�n��������@��|������J1�ٵ�!Tp^��{j�v�x)�W��m��I���%�*̄4�K!�O9�Y�/y�
좝[,�Ὕ�Ч�`�aؤ闷7O:�j��{[��9�����C��3Y���nQ�)vP���G�8�[����7l&Ns�=�8�IsO)�GW�7����3�m���Zq�x{���wk������PL`t�N��4:a3.�1����xY�!^��ǂ��%Ƿ}r��E���K�8:��:	���rm/2CtwS�@ݤҲ�r(/�9`PZGp�O�dJ�����ۑ�W�q�26F�u.V�9��th=��0���Q��_h���.@`B�a�2�
�n��t��7�����qʔ�k}��֝٤W���(�����98n���2X]G�#���V�z��W�nݶy�}���P��s��\k(��Zfg��J
�m�2�D��Ԫ׊�G�Q�ln����޺�Γ�IcuM�S��\�mڜ�����&��qr�*u�Mߢ\:�Csz�5hwn���.�9��!1�o&;�c$���TV7�+��:���kq{�^����3��Ӿ�c+��ܫ��#)�F�I&�E1� ��Y8Vs��s�y�����7(�U���߆���O���պ��f�ա�V�r�l3�������w�
�	�����������]���������V�5]��D.���P���$�Û]���fS�Gc�{�z���R ���ʳ[���1�ae��y<��
n��7X�s�-�x�5;f`�*���)\)��Z��3?K���?;up�[��Y
ŤH��=�+]#�}0��h��+$K���q%eQ���f��{����b �$��~���VpL���}��I
s�I)�J�Nf��4���p�e�L�Ͻ�V���"V}���j��}�|G���±a�o��{\x���V@x��|��
�X��xCG	e7ZJA�i�T}���j���j]���>������_ܲ�X�����[�h�0�=�=�z��-�l��۞�	pL�TB�d��W+�qs���/��f��2��gܩ�]��!i�H�ץ��%����kr���حt��w�<Y���mYD����T�j\AN\��.�xX�6�W�>��v�/��X%g̽�nİ�"^$H�\���i|h��#�֬L�!���괟n�����*��ݟ����?h-�_�m��������n:���id���
�f�#D�,āQQ�����YlL��vK�T�Y!U���r��/���PܗVQ�5K�4�)�'��^G����2�t�����:.�D)�%�}y�|BӀ'̛�,��v�_�߅T�#�]���^�,]jHTy6�W�f�ظ�B
0ek�&s}�M�~q��%$)�w.G�]/�U�s-bq�]���ƛ�����X�\����h�[	�Z|�,��(CK�����Ow�����?gg ZX��|���X���TB�*"D�P������I�(t!I�f�����n��;��������@Y�E*	-�����Xp�S���EH��],d��B���NjJSR꨸Zn�x�����p�/J{w�������s��Q	�]����b��ݩ��d�;���
τ��㴶����5)H�;���~�xZ��c�'ӎ��y�������:���������-�.��..ѷD����"I��"�����n>:�[� �
s�fr�8��t�\P��{ֹ<���.�S��|�%��ϯ8_���mtT@v�*�&vޣ�\������ׅ�}مV�1����7ئ�MKnfi��d-!3�Ң���z�Ig�|G��S\�w���#��!_�=E����s���K�)sŋUr�{��W�6{4B�ᴤV�.���������oeL�ayy_ؾ�kFgo��i�F4�.jsӨ�
�BT^l�2>ɞ{ן,KPq����aF8RI�V��_����w�z�#��L�G��(�G�߈���n	t���[��^�D}y���9��]\�丑Kp���I=��;wzU���݄�G��[&hXW|x7�UH�(�-x6����,��V����&�hZ�}��Y����vjx���gk����U�$N05�q*��p�A��YRe(�b�XJҗD�mF�,\$��㫎�`f]��4k)�M�DE�њM9�2u�Q�<��iZ�ƣ�c���6@ �V�]��gr�2͋hA"M���;�f���PB1C�6,r,�\���%4���1M-��#��b82�g��
nm��ph4n ��8�ӱN5�i�cgt�4ݘ��-|ZuLu�X��c`�nL��e��yٚ���P�I�]=���vv��j�eS����#�}xe ���]	X�u���#�B�1P��}��!s�.BrҐ=�.���<�[�;���I	���ۤ|Y��w���Zk��O/Bϗ��;��f�1H+�H_dX��%Z}no��W��M��{�0�]�͉X����>㴸W�ڣ�4];֍p�b]���ғV��j���t�{�7�a(J���s�6�@��lܭ!��h��>)�
�U;�#����i³-�~Ʌ9�ɶ*$�^5&ۄ� 2x1G{�Я������#�ᅅ�J[�H[���o�e>�������6�F�
8sﮗ1�G`XB�s�4��L�UD�J�|%� )#'k���W9���pK��w�wbb5�"E��,U�Z3��0{}=��>e�*(�ȱX���w������XpTE	�w�����9�W��U�փ�8�	_&c-�m�y����R�JS4'"�#��kb�$A4b$2% 0{�w��kẀ'"�d@Q��ܔ������^����=P���$-�+��+s̫K�/���gnid|_��\.�:_D����Υ&YKE8Y\�>~M��{�.����%�e5݉j�n��BѤ���l�.��/U��G�ܐ:6lp\��<�GR��9-z�.��r�R5畞��Z,Z��֑B�2��=Y� ,JN�(�u�Gᯯ?+){��7(/ٸ�;�&q�Dx��V���U��8*�t}]�X�/�߾���a�`�O#�v���"��*+�ʸ�h�w�_��P��,���վ۵6���
�]�aD�J�U.�ѽ��J�"v���|�Y���8�W��{��/����0�W���ﴏ���҈���wӍ|1�|tVtYѠ�,g�ť��Q�l
#H�^?BO����'�H�����Y�_�X���%��f���oD�8dp6�nK�x�i3�gg�Z�H��o�����H���_qѤ=��qgyu�H���o�«���HD>X�Ssyٵ�hZTtK�lJ�b���Z����%X�H"��i������f��F���W��U@�)_��G����8���*�4?�H�B1* wMSb,l]���k�E)�>��R`���)��S_s�^��s�_��
�d�(�B��J8~8���ZB�ާ�;�sT��:��ij�8'�7��f�ůf�K�w��*�i�$d:p��Y-�惡��y�د��6����*��G��0���V��g�.�qԥ�i|���G��^���* �rĨ�܅E�wن��*�8/����H��z��͝����nsa��Tkm֣�J<c����[[]eK�f�܋�O����_c@	X"Z]���Ti�1�1+��@![W��?�\W�H{�\#]�Rܢb?�w����(`��*��v�ZQ|���0Js�ٵߚgH�Noy`��J:�D�]����:�)M2]'US��௏1��\��ƺ,(XA���lYGN�������=s�i�G��_,���q�t�"ZH��H�׿;�- C������s=�|ŜtE����y�ϥ�8G2�}�$S=��Mq>���T�J���h�_D)"�J��{<Z�i�+y1�^<��@Y##�{��;ƨ@_v�͑t�7߳S��׌NǴoS4"k��Q}�_Av�j�X�t]J�G�դ��m_|m$օ�k�m��b��u��2w��ϗ�-2_�;�f��Й|%C�]�_}��k�q�t������ο�/7�D���Da��������k�F����"��(�2w~~��;1�&�}g�}�a����Se"u}�I$����p�����Z�5/Mu�f�a��{����r��X�{��|�����#5��l�
`��Ds��_�S�%2�'*����J��ӂ�D���v�,��v���DL�
HW�"�lyl�z�z�^_�W�0��+z��Ċ�Ra@�8��j����ְ��i|Q��{��|غ.K�i�Ed{�=K�k��+�zo�H�W��J�K�.�t裤�ͳ��[Z�<p��{�h��0���,J@e͌�#4S�����O�!w�TF�A��\,־���#��Ϲ����oV, �.oj��T,.�^s�M�M�{��s��#Uސ���#�ȑU�9V�n8B1
hs�u�I��U���v�hȊT���6<Q�Lt�%�:1=l��ɘ9�����H��BǢ��~����#Oómυ#uRwK�m��!����p���[��^��e�|D�Q2Mg��>�\!����j<O/����qb�/���v�4�E*�3Td.�4�Gf�,�F��rN�/���؆@��*MP� ��}V�A�P�߸Z���ϿK��i	�߄�9�i{Tn4����������?5�b-Е
�$d.j�Mbi���8Kr`�C����'�f�f~���1��q�Dz�G�����\Y
��r��ݘs��p�M�TG���c�c�%w9�r%�)E��\���g����b�}�+*=�q�B�N���1��[�ӎ�N�eG�s66����V���!� 4
!�Sz������2�һ�?,���i��c��k�>مD"z�����L���{|�X:+,�>��z�^'�\�:-��-�>6Ќ̿�����y��Q���W� �)�̢�p���}��Kq¤q}ʮ���e�9�R�����o��~��*�ò����̳�ퟮ\���ٯl�6;x����I^{�78+a即�ݎ|�g��.���P�*��o�/���
ψe4����;��w�1$�M8�\D}s쪸𴎊������K�>�zr|o}7�D��6)�o%�i�Ϻ�o�s�e6&E	�˲��f~|��p}és�%�7���e���
J#��J�OU{k�p�[K�H�}_�]{;j}����I�#e�a��'/7f��/W&(Xt_���֘���U+���(���:��x�ª�~i�ӷ�es�D�W�b���5bR]���n��"T�+(/���t����
�1�p#��W�kl�z�6Y�ߦW�i�f@�������|�����l��DH��Ɨ������fS����q�j��}Y��M!�TGM��~�A���r�P��j����j��&j4��VE�����ki�.�+ܻ��Z/[�!}%�*<�_�u\x�8�am��[VC
�K����rzC��0,�$�鷝y��C_YʗW��.#�s>��|$W�g��$hO���/�
�-�QY���{��!���t��������}�1Q�����Es皾��~�=��G��_�!p�tTG��V�Ro7ih��}ڸ_H�)4��]�^���a�O��^�h�L�=MI���X~�����-���'������͚T�C⥉	Z���gbĸ����RΟ��ok�%�T����Vs�|��o7�]س)���-s>����_H�	tD6�6�b��;l
���h�ؔ%��+i4�� :Y�un+,D 	s	��P�C/>�۩۶�ݥ�3˦З���S�	���Y,��`\킔&���l5���j�ng2!n�_;� ��np�F��'�;��W۴��g'q���]���!{\r؇��n�E^!e���� lii-��dɻ8��b=�'+-��^��iJH��.��;e��v��s�ՕL�k��uD��ĩ�M�U*aT6��^"�RBb����K������}Ư|�0�ϴ%p��sbɿeU�{��%gEv�w-)$�a�� {U���Y]�ۦyG%� (����Oy�-v\N���q'n9��-�|�2�)m��.�j�Ck�I�C�@���d�D"v��J���/}D)��G�MJ����*8B�=-��[=������.q>���1��z�EH�o��Z�f�A8>|�����`�#�<+!N#A=�U"t9r杩a
HL�{)�Ƒ���� 4�9p��S>,�|/3nn(]���6Z�*����hd�:B���P�}(<kJ�F	s���^�rr�Q̚���B�(mwLs�
J��"���%�������$h�~?�ӡ���1��]Guĩ��u��w�_���m�]h�Qrae�y��S�.����BL-�Jn��N,i>@�d)�#��rm�^yM{Hg�<�y]�`�֩��$�*���',�0��SN��T�p��O=4���=�D`������q������g�~���M�^�ߢ�������8��0�J˦@_gيҴ��	;�H�h<Nn�(@��o�H�i�׊��!_��\�zNUZ������"�#5������.�vYLJ���˻�7d����jՌ@�V."���l�>��8T1 _o�;�U�pTH�b���&X��ɬmw�ߕ����Q'�X���F~_�}-�
�U6R�f�ח��>n�(VJ(_k�,�9��V��7�P �ɧ�J���c4b�{�ʞ*�uN�'J�&�mN8�e��Xp�O[K�ϻ�2(�DD/�Zk��};���.���:�.KDX��e	E"��Q�:�eD�W8��橯�/V�KTܘiڂ��������Yǩ�Mɣ;��.�A���߈�ݔ0�5���m�Z~���yk�����9�ӈ��]���@xE�L_y��҂��%���>�_m�]���:@��7�%�S瀞sB���
uK <{�mZ>ƕi�B~��Z�0U�]i��ݘE��ϳ���;�g/�(�a:�eJ�~x��W���J���,<)|.���o8�h�h�,�J�;�9�}�a���QJd�]4�կ�|�+q �<^�c���@�Sy7p��e���)�|��z�*9Ɨ�ދ�j�|=cJ���Y�=|��J�m*�0#9�\ռ)�糙�V`���ڒ)���>����9�0)I5U7�� �\�I�����znk\��k�Ԇ���e�W����@�c^ߕOQ����0��c��$�mV���i³�K)�4��7߹��8.�{ ie��X��%�4�T����E2 ������-�y���8k>6<��Ꝟ��6�ݱ���J>v�˩�2�L��\�|�����Ք 5e��3陸U�WM}1$�+$�*�����&� E8���/~��"�w��__�V�G�ƤZ4%]��.�϶�f8d&%$�+"+�uX8@�0@��H,|�#�t�a�5�QJt�U�t�x��l_v��Ï�����vk�Y޸����!��관�)=���%�i#� g���Y.}����'�9	����X���M��.�.���K����.8��v�<�w���ş��Nʺd"�?�|�W⾩�O�t��~q�{���G����Xtf�<`0ؙܣ�SWl��GS�ĩ��E�4V��Wbt=�ma֫�.�N�'�)LV��V�[~�����k7���;u��O_�Ƙ�X=!z�xZ����#��_a����USsH�JJ*j��n�<�&;����:�����	�wW~��-���H�K"���V)�Lz��Z��ʆEM��Ȣ	��L��B������Qb]Þ�`�+��r�	�	J��DX�b�,�^��%]3T:e)�Ub�9�ǭ5-�"A[J����OUj��8,����Z�4Y�0V,�����޺����ϰ����Dp�"��D*�C���iM?q���:*«�s���t�Wr�E�Z4�#�s����AV;��HRjw�F	;D.vW.�)�[���Z[��f�fT ��\K
��Ơ1Ց������]!2߄������|Z�8x~��1�4e�8ⳗ>��[�~�$I�� 2�E�����{�W?ۯ�E\���GNߥ�z��	}�E�O~����[�����6��G����/
�ԒʥM��y
�Rh�O��Sb��ϽW��ω�}^��*�]��ѫ]k�ݹ+�I��>~��»h�u�)s�\W)u	�aG+'�z|$O��1f5ÄY&�ׇ;-�ʙ��|�M�D4"��k\�L�K�J���ԙÂ��yJHXv߸� ��=�sՐ�.�)8a�fA2�!������p�Dn���|̬}���q�zt�����q� ���BAEc�r'}��."4���6�0[O�QeU!d�P��)�R�:��Z5ǮgL!b���^�>�]�,J��ڬ�\`�\*6�*(߹1�����.�2$��I�TxJ�g���x��Ks��S�,���S���*O�ƚ�|[!4��Cׯ:&������祡�\�L$.�=�f@,,Ӯ#�|��[��5���8_l
U���~e��]�A��P����v�b����m��&�,��<�,VB�~vNܑ���vn��j@e?�RLĞ�g�n�J�$�~��Y	�<l��
f���$B�T�-/��=��EW�ެ\Du�T���5'�L�$�^��z\��Ȱ�Z�fO�HHщ�s��"v#`Cb�[۬����C�d��j�\�9�&��2�(AR.� �����Q�0>iX�B�������>��u�
 �p��H7���>��Y�~���'<�0+Ӽ(Pbe�}iL�߲V��E��6FeZ����o�������˧�O)������%A�V-#�|k��t����)$��M*��VY�59�:x�U�.���s����4W��X&u>)����H��dX����խ��Ӧ ��˓}Ɩ��^�qv�}�Eޒ���?����	/�	 ���_���m�Ta��0���?2.���i|���ww�
GrҎ��Z�����;�Ǯ��w��4,c+�N�/����H}����k��@����a�<!����|E��Z.s���TD����%���F�(����sI�����9sJ��zQ�����]|f�1q~z_�u[~�w��e��DX������z�����j��X.F�N��g}��A�Y�Q��Q�pK��py�L��t8G���}J׈޵�ܘSm��Q���쩚T�R�,��#��y";��??@�1J���ӞPߗ�M0�&KR+�n�Y� ����|����=0I���w��ih�H]	;��	����!�/u��2��%�_����.U|������
��q~˄:�B8�锲���cs�n��]��{nIy�3�L�}|�+nʨ�Բ!��{z��h���z&��u�@�.�b������cU|��r���:қ��b�=�P|F�:��Q��ʕ��"ֻ݋.�@��o@�V��v&��=�����]�s-��܄hҜ[���ʙo��\}]�W
V��k��7�����>��N��8N��֞�ȗת�pl�j6���	%i��D``eΛ�F�x&�6�Nf��}�X%��}�xV�p���\y#��ꕮ��8��-�7j)'K΂�np�H.�o��u��𩽀a��V)��:�3[��=���K�w�)��[�r��%A�Cv;�\�P`�U���q����H&�����k����Q���ҎV,�B�v
��/�۸��5�|(�!+�q��(�f@\^�b�� &�V�^�f�4C�a�$gr#q�V���0�{� \ba�FnQtop�:HPW�p���	�3w3�͆9�YS��Ѭ-����]q���ea��f�giܫ<��[\cT�p\D�����,��2�wC�����r��f�٣.cw����9�:
���6�"nu�:2��h�&k�L"��.7YZ�Eݹc n^P���^�:[a*�Ɨ���]gB ;J�>�mR磧.���&��Uh���|�.���B_����7OLۨn]��q�{*���d�sMI����S�&�m�d;�2��Ŧ�E�5ݪ��>y�[l�F�cH�=��xu����;^b1=��;۾V�Ū"+���5&K?�6(E�n���K�u"�&��c��lm�e`@����m��<�r{XЏk�n�N��vg��6`Fڢ���nd�:�t�ڲ�I��ܦ�n\ȍ��$D�ϐ�c�2݌��8��S�"rc���-��ܽFČV�r1��u���8�����vc��p=7��M�b`�+�B kV5+��u��/�[7�4ںa�l�<��ӎ��-�KS�%.J8��n^��Ke㎒��-v�o6,��˛ǃ���8'Q�s��=q�V<y�m�\��=�� �\�ؗK.�6��1%��5.����O=cv��Ů�=�h��XM4�@HdWQ�	m��fL37D�ՅM�6��Z�ʱevk�8�\p�t�j*EL=Pv{���x��^�j�M��t�s8�u�6�ENz��'u�LC�=uh㶮9 "��G-a싋P�V�O%�-�9����b}��Cl�n�b�b9W*KCD�B=�ea�m����b�B�X�>ޠL�`v��F5�l��p�b��v��P���a�M�8E�ml�s�q�V8;�]j��^�ny�g�5ׄ����UǑ�^ݯ(��Ot�GH�;i�.si�l\Y����k�F睞\I;c��aV^�-m6�AJM��a����B+.I��t�ͱ�lmۓi�Ѻy|�Hs��덎x]�.��P�=�5PF�m��Gqk&�4Y�e�L達f|�3"�N.��93�ז�G�
Ax�͓4�����ji��7R\���	�,b�7M<ݽ��/���˱� �����w�yyv�x��C��Jf�%
�����;a�q�lg�4I��]p3d����#3,�cZ�|�� �5U�l�`T�� 	o�%khQ�=���k��o���3�X�\�=�����\��Vگ+4D0)v��P��{;��sl�EF��%�3/'SOC��;�n[{E(��i�F�K�	)��G���S��y�e���������9G�g@��i�t�}6��zW���! �n�f���b�,�TKc�YV�ݧos\���/��.�+V�GB����Yy�q5��ն�!5z����;8������73v�v�m���;��'�����^+����[�!�,(���z��mn)�Y�+��s��{c�x6\��=�a�N�	�?�/���]>̅=�����g5c�o9��<:6ۍ�]�f�RI9��W��͔��-I؉�� ��k�ڻhL���n�>8����
���j�6�;'6GbI]�']/)��?��>_���5����Qx����XF����T�P�n.��j�BM�)�)!I6Few}��o��3d��w��	aDi���|�g0��ĉQ�^,L���t=_��I��U6S�<����6�������d�{��![6C{��+�.�@ �qL*V��ti~߯��B=�p�4Y�,VN��8�����>"���
�9�h���_�o�z�}{��߽o/�'����|uXe,�ZE\�t�z�����{�v/��H�D��龠8Ç3n�]��]��K��瞼]w�y����オj���Z�{��:,6��b ���م7����q<k�|"�k��ӇEb�\1W'�_q9�SRS*j�8.�5dX��<�"�U�O��8?m7��߿;��<W�wۆB�Z��Ԑ�y|���rc��`�B��L�	�����:���){��w�tl������Q��*�9�[���;徘���Cu$�ML�gƌ\"N�D����Yo	$�|��צ��<�64կ��O�I#���!��g��鑢��
�ʵ)��<F���ɵ�������$]M5Dk�ݪ�]q��aEݽ8E��S��s�Т�I��֜��Om������k��]X��CE�E�36lB6�mعO�=��/�.���,�\abT����.6���M���Ĩ[_J��^��#�<.�����`fO�f��`ϯ�oS��5�pK���b��vv�Å�|ڵ9d�[�,"EEK2���<)g���b&�D�S�\#z��c�Ե�I*�'k��n����k82K�u�UEiW�Ҡ��u{V��K�ʦ�n�cRg���m���꺝�VS7�oti�����j6�K���8�܄�t{=�a;����GcK�Hʾ󾭅w��#؜{�6{\�H��t~��w;��=��g�� �� (�g����#�2+��r��%b�2|���d_�1���K�X��]�޾Y8Q!߽J���i��J�wj�@,Ϧń/f�)$LO�=ɸ_?r�h�������؞�r�~��x~^�a��3+�Hѷf��Y;��*� �ZZr�>x�!?���ɝR��RF0Ӓ��C�x�A�j�v5kߚN���,���9׈$x��b��!��Ȋ?+��鐶�i�G~��RY��R�s�,	k�­w�$�?3��k`�U�������덩�Ej���k�ҒpXǏȧS5Q3SU6�B�$R+"�wW7��G|���Y�J_
�-�ٙ˧5鳛/�ms���iE���h��L����0��#���υ��8a��vmr�c���)p��Ҙ��p\��w|�?��~���!���	q�W��Ss,��"�Vf��d�Vn�a[rՀT�r��+��M:�n�}"�
K~��H�x�"������Zp;�@,���Y
�=�Vt�|��� :�VF�%fS�����+��/���{|�g4��𳖀�_ x���s�+Wׂ��Y�M">>�JeZ�=JոUg�8T��KT�j�8Y#�����kY�w�|-�o��T}��'y�;��&I�W*/9��`Y���Kͼ,Y�"�s���PRXp��>�����^_�վ��8[A=�p�����w��/���,���L�1�h�0��ն�ݬ)K���+���N.��'W۸�,=N���o3�D��u�C��<����7U~�s`3y���ẼN��c]_J�}\;H���0�4ڗR���[�%�[�'Ml(�;Z=*��r~�ۓ���@?Ww��@#���H�O�����y�M��8| ]��h*;7(!Z�߸�+и�͇q'�u}'��6���v�-�i�����
t�55C&��;_{���f���QD�]�c�8��J4��g�V��~������t5S���:�<~�����G��?yД`I�d�&���_.�b�,����z��~t�iNĳ�)i��a���5�'68���Xw���B���"��٫|w2PTp�RBb���4ؔ��Z����
�*_��l�,e�ٞ3�vU��1�Fi�#�X�)�ٴ�kL���'+�t��������Ytу�ь�T�'��L�P�E�뤮�\��7�M���"D��St��=p�mzmj ;�(Yd|�E��t>8f���is�zx��*�̈>_#Ռ jVE�����t0�|I���*��r�_F27�3�S3bH܎����!��]��Rdf9;��M����b��_z�y*H�|y=�y�it��WH�MK#o�R�繓kH
���H������ٰ�A>?��w7
p�]�7���Yu�ê� p�A'�َG�0��Ȥ9��$�/�}>-,��x�|��F�RE!�g�9�p��;����%>�4B�_;ZE���H��"LJ�:�/�{�k<�80"ys
��X����r�rQRK�u��B�4qy�!Q>�U�O��p@����}͜�b�&{�:%�}�T{9��� }��,#ƛnD��*�ܬ�p�*/���U�pë����R���|�ӥ�1,��;�]�r&�>�YC�1�V�8�w��FEz2��F���&+�̧lwM�r�u0���u.�tzFPYl��8���ڭo��$x�wf2��"A<���遜B*T�!KsS�]��������n�ȧ�rm.Q��^5Dw�7l;@�!�b�����+:�_3Z�Qㄣ�c�\��p�.�O	M>����mfeM�op�����a����W�",�y��������
_����nA˟6��1X��{5hxɍ�iأzM���jw)���Fl,�?O��|м�Q�R����n��)`��1-��&E��q=�}�!Z�$���P�-��{3�N$��S�����$�`�D�˽n������DN���?{���4�6�j]T��q_5dX�gUʑX�T
��W�'������_���R���B� ���_j�~t0���3�UMҲĨY�;���}}o����#��]�?` i���C���D��6�VX���������ʢU)�5KU�-Q�|q`���_ޛ���E����E��]��Wÿs~�L�>}��\����U����Q����0,���߿oh�DsC#<�m|���+d����PJ 1��i��ώL��J�N��|��}���~�����"��U���>ʀ�D��U ^n;��99��g
���8C��iw���k=]�U=�Ĳ�k=���H��7��U0�Q�ケ|Ei�=�(����sUY ���L��Z!����NF�'��I
�$H��}ߦ��}����]���p��$���L��B��6�A�6@:w-)��pv�ª�W��\#I�aM��LTx�?ɮ�_��_���h
�7�n����[��F��\t�r+^;X������mr4zg�(��Eۭ��c�7��q�y|0>S}��ʘh��K,P����k��ik�I���z��5�T��G<��#keb�Y6������vƟH����,n2�=�2�x9���n.v�fW��ԑ爅뭎�vrzŞ{%��M����`�����V�H��b��	o]Ζ�J�LQtt$ؕ��c��X���?o�P˝c�\ݸ[-�'$u^p�ύ�u�7�*��,�#]��%�b����Y��9��;;�qD�cF��5���f��1��,��x���^�m����#�P�K�+���~,4��b�c�,�˿z��-�2
��ǅ$q�0�����P�ٳ4
�Vq�� ��i}nȠ�r{ɿ�^��t�������%�O(����|�=�H�T���:pO\?6�kߩX�L\���j$yr6a��������>4����Z���_�P����(��F�z�hse�W�N:2(���t����}?��F���������~��{�A-�
M�����J�"�T�����.J����|��bY�[�z���qBL�[�F�d3?{��?k�,�Yr�����y~������"O{��q�;$����V�*Iɡ|/w��q��\�
J4�j�W�|���_(�[uTƨ���\#k'�d<}g�뵼 ]p��|�dQ�[]���L���ӑ,����#}2�1m�HA�:�����zVg�X�i��-�3^�W���+H������|<p����# �|.�[�Ki����3U5YH�w���&{�x�ʥg�o��xX�����#�o��~�9m�X#Fz׼8��\�������Y��kw�~���>'ڟ���%dԃxa&�W~���B���c�X\_z7"�Ȣ�?>���r�j0��%��κ�+�[���b0�ؖ��X���6�Bh�0P�l����ٱ�Qv�0�?3�}ǭfSa+rO�~�@x�U6*!zӅ$sZ���U���TGTA��	�����n��G,�xw��m�� g���"8��}�|pɟ!��Y�{���z�l�>���Ha�vh�jCL�-}��������f~~��uk�D+U�0vd�5��FoU���ɌaDWv;�jk��v��PTҦ�K�# WqD=x�8$�8�]=äS�^V�~x׾c��-C��K� sޚ_7E4 S���lX�N̐FKE8N��R�!����o��+)*���e<zi}��,�b�W���{�����&14?��������7�5�����^�ﻏ[Z��*m�±X���ޜXi�<j`�:���KC[>k�*
�۸����U_v�y1{�Mz��Ɠ>&>�9�#��hT�p0�����`�y���"W��h ���h {3,-�)b`[��ssR�K������&O���c���<4[�΀Ac���|Z����Q�U
BfY>lYU���jl�%ؕ
��ߪhMٞ��#�RQ� n@�V����٤-�k�w� ֦X/��O�e���0F4����*��.��IsOu��q�`�JJX0(`����\���b��Z~lXY~�V�5�I���C���O����,Ġo�����k�b����{���2�a(-��*�Lo��VA��qd`&D��	kM���{������>/�n)5tD ;%�T��F�m���N��<�7+�9V{9ڳ�\��Z!���ux�|A���Gҋ"o���`�Z��0!������yQ]���0@�#�@H�c(�"�Ĉ>�g�V)��esS5�*i@a>�@ 5P@���ݛ�Y����Í��G�|ѣ�	9���/Ϥ��	6����X�>>
n�& �! Kd���Q��,��}�?3����;�d�H&�0��1��da�:�f!I�Ռ`Q�Du�7����D9lc����%�?}���}�>m|�:j�A��t�������Ȍ|�H���)�9��o�6 �y�Ee�3�N׋[�<9jq�%[���eVU�H�n`י�� G>��IZ,�}��hjS�C�1��3r�Z�a���썺0�cu{e����D�(�%M��xk�5۵g�u�Y�P���^k�����gr������W���]�9�=��iM�˽�rxD�m��1�J�k�@n}�ͳ.�_
��%��r��E<�B���ڧ���[�s3PQ.��R�+Ƹ�9*q���rL���^�� -?�g��_���a�#'-����W'�hRD�R&�g�>�{&��Y��>rtm&Qx�#m}�K�����VW>�HI'ޯb�=(|jI�4-�D	��fQ�U!I���u4�!f�ه6#�Q� ;���E�rW��Ûo�k�s�l}��A�o�~̹C�$r �.�"�ȣ-�Ͼ�U�A�w]!�k�1%��x�^*;�{&�7��V4 D� #-�ڟ��f;����~�:�r���b��k�wE�#�����M��>�OJ�y-+5WKsƎ�Z�~�����MS��E%�_zs��;��h �r�6 �	u�{Ȱ\䯎c��q��X����������g�r"ld�c�I��>�&�҅$�����Į6� ��I؟!䃴	���6�⛀��P'#���|H�0�E <����j�{�"�V��+�GH�f�!@��ߝ1�������P�
,˻�?��Ve�gDȡ�z'¨0���/Vfͫ�ZpHE{��_*�����a- �T�{��U*���e**h��i��D�H[c�vw�y���-�B���^#���7ʸ�=��dXc�����5�UN�6�f�:@�'�a��3�!�
Nk�l__=��[,�s��)���G`ud�#�0Tw�aB}Y��̎�*b��S,)�<��w�Q�+s1�?9�Ĭ^���ݫ��9֬���YN$E���z��\ 
�j�!�b�R�GreP�~��k�����K:{����~YJ�~ѾSK#�+���h���V���iM�:EId���Ue�������jβ2�����eml�h�뽼�ƴRu�VF 4`F�uMM,Գm�����mw�����+�%�W�,�,0��*�)�����@�!��"�(��ˇ����s�����`4W�f�-����h�F
q���^Vz�.����O�Yfh)a�s����h@��Ӳ�4i��b�<{x�� <�y�b��`�L���s�Wؐ���h�G�p�G�).SDJVrTqu.�
��OdK��1�n��^���N��u^[��q֎��X�ِ+���x@>9)���B%�w?	��*�GVMI�Je}C߭�Dh��D�	i3�~�'#I8&.q���%�	H~.�V�~66n$�NH�NN	���ЄXĤ`��e��M��GqY��\�����p��ui2�Nw{�İ�Rp]u(!e��cO/����/��eD��?�`�\c�������1G��
��<������r�N��)T�d�U5UU΁AmQB�[})[���[�<ʴ�:֔`�w�v��֯΂[w�������iyx�����<]w�&{Ǐ��Vv�j�l���Y>i�'MΒ��y��ri7O/۵���R��� �٠�<Y���1��{{�����E�4�"�Ä|�*�dQ?p|�T���m��y�w;�@?b���D�;���!Z��g}_c��[\q��LU"� �*���;6�)��0�l��->���	�N!"���b7�Pr�aQf�E��p����4?K��U	�j�ਗU�RE�0궕�|?]^,��eӏZe�ީ<���b����%��U �L�����ks��҆�r�ҙ@KU�A
ړ㦔6�h���o��)�]B�Ba�4��y������l��6�e;
R�/+7�N(�oH�¸�� ;�6��X�N{�L�ۇ\��$8�:,�﮴�5.̡�Ba}nw	*pa�z�pR�>-�an����t�c=�V�9L,	���8v2����]�0�b�f��L��!��#GK�v�wosu�� ۴��1�on�r�k���[9ǭ��͉���,c�u�Z��8� {]-v-�V:<4�k`(-l�7l�ٺc�j^�;
� cKq�M;7>X�<&�,�8���-c3�*X�J��5�.��s��H*�C��ˍ�^�����qh��Ÿ�0ԇ]���H�r@Y�?�(��r��ȡH���f~m�� �a�+J��#|QL���q������%C�̯\��lw�x��5��K�������b�{֭|-8Cӑ*#m����{92�)Q32¨t�j�ap�U��+Ƥ��+/��8��g<�����\;�= ���Y��ź��-��z�ߗ�q��F�$)i0�����q�tT��L	s1�X�YD��άH����D����z�\q>jȢ�ź�M�(�tɒ����)p�2�`�(�o�O2�zut�7E
�U����U-Q5���#H��f�+e{�"4�Aֆ��w}9� ����-��$�NPbL%�3��Š��� �������
SM����1Rc�ꥲ���ՠ��L���P꾾�lUC'��!G�!wޱv@�F�h#�j�Q�`�z��9%Vm�6���0,V}-,�{��,|lBmL.J/�׾	����b��7��$������2x�m?�e6+������}�Y��-5ՙ�l�׫%����*;毭fԩ�u�ߝ�CgI�ƙ{6)����k�u���s�̵�}�J%�#�J&����V`��J/£��bb�iJ�=�_�\���\Ȁ�>�̱���TC�|���7�~O*��h�P��4K�Hu���#y,���ԫˣ���rd2��9vF�,lS*H%R�n��>�:��L�n�� c}𜹿�X4�1 ���[  �k�������R� "F�Њ,�o���?o����{��4�~ٕǂR��@�6lV!��M�a�oxd�	~�؄���C� ��"�rT�hm�/���>g��\�@�R��jϯ��ň��[�t�b�)�_���))l����Q�{�b2�ʖ�r쥖���|$%���[�������n:�|m�C|�h�>�^H��@��L��}=�9M)ALn��rn0 #�	�"D�H���^B��}̟?�]|�>� F8�~�?�� 3mm7���'�ԁ���")�݋�}��+��h�M;����.��0V�S�U�l���9����4 �,�����ߗp! �$�K1��u`��>o��N���l��緜w�u2.	�� R�)�5&�W�ܿ=��1V�)����e���a�6��~�߃��u�X�7�ZC��$kd-�Cm1 ������M�^�)T�#~�",L��"% ~����$�"��1!�~4���wl���N��N_sx�c��4�Ʈ\  (�Jd4 m�f}�2}M�өR���:㤖=E��tA��#�v}���k�	:L�Jc �p�RD���_�Q��� ��o�$���j��$bbr٥�`[�.�>糫#[���m@ٟ�����L�JO�=��;*P.�c�ɍ���$�%� �_��{����VY\��Js#�S�[��4b@z�ί<i�lm945Ts���ݜZ�-���(؎i��~� �����׃6�������8zX�����@��@��WHi� �R�_9�^�>n	���&�VоMf5ptf�3ڙlG���ł��]�����1�D�6�"d^�N`� ֙� ��O�v��o��6�(UR�(����l0J��XdY$���Z8��#:���U� �ze�s>��@� �� =��KOR�U��w��������_ `Џ�,�$g5�Y���S�������Wm:m�!)Cj�מ��Y ���=>9^�)P��>CCm�I�{��ʪ�UT�%7To���	�`�`2[7����=�N`  �i֥V�A�׵� .W|�kI�w�� W�M@$72��乾�h�{�_*���0����_����F�%���ѳr�&��ú����P��2ֽwR���V�X�I,��y��柕n�X$����c�0�Ϗ�܈��ʭ]�ѧǰ�<��t��� �X�V����-���L�!f�P�I:�5�c-A���(��j�����;�_>�ζ|J<�j��g^M�ٳ�B�*M�U�x5�p*s����RX(shd�7E��v�SB!�o(�;v;Zop
��aC�V;30��>�lEѝĶȈ�]B(���9��>�v��s���]Ӗ���������d�F�3�M��C�J�7�GW�}L�ϝ���5.�$�0;�J�чf�)cyҡ֢,�s�g��-⫆�_I���t�\�^V��f&�7R����d��{sh'c��:i�Ű�cDVS��幫M���M�ťj��J�8M�[u�z�UĔ�Pm����W�׹W��e<�qn����H�
T�Zc�Օ��z�wX.e��a`7����F7�(v����{�f,|Wi����v�6�{y�\2�j%z��hhi�
��Ʒ3I�.{�7sV���q�w3g`$�-n�$����ҧ)3��nf�.��������	/���K���"rݫX��%�1I�;����
�=�H*��5�e�'��[�d�Gw<�2���uܐuC�i�Äf�^���!u���f�tr�3���󷺨�Mq���ҮyA]����ں66��a��I&��ү>�*����x�ͱN\����nƘ����� ,Ҩ�����7k[)���[�`ch��9�1�e=`�}�����]>|_~���F�n�J�>OV�>�e�6_s��>��*�� 1�
��ŀ�����Zk��Y, �V�!��j���Mm���m @���n��`Ri�����L�����R��r�&����� �_�N`o�-8rYZ�4����!�@��3t��3U5S-��� ���K��& ����TR�{�x���f6�<��#Z�hD�yߛhuz��O���B�"y/�Ic
m!|4��D�����z���X��}n�@�-��`m1m[`C�9�pM�ƕT6�Xi��l@ ���z��r��!�W7���b�f�E�û�u�J8B�k�;s,є�Gl���:�V_�%�-�� ����cT��{�ʱ}��Y� ��L R���ٺMM+j��*Ji�^�F 81)i�ne6�m��F�~�n��Ş���!����$A �� �]��!=��^r�msmH EWs [`��G��
��D�f�^$ �%� S�u��2�؄��Y�1$QX
3����߲�$��<��$�P�*���T��iP}��2:�Ϫ�@�-� H%�/	��Ԁ'{�W�[�D�K2� %m��j�1�LP�G��j�Z&(����'�J��i>�2>nHz�B_\��*rL�R�AT
�f�bQ�D�����]����D��"�%$Bd�%%��뛅ӂ�$/���3z�z���DY�G;���lƐ�	����;�f+䴖�Z؃��������A���	��|�F����ǳ��1��� m�]ݛIpK�RD&$��/�V�V(U{*8a
�UӘ���j�t�	H����h]��3(�΂����ռ�o�����sMkw#�,��U#՝q:r��^#8EB�_c2f(�=/^�Ǧ�+������=8
?���� a�*���B]"D�r�f�|��̪������J��v�XB���
��;������ |�R���)=�y�}�2{W7$)0�S�D.�mE�Җ	}�*ݨ�NH!&*Z*
,������*#u�,"�Wx��_n~���#���n��n���̸�e�q�6Em�(��mx�WA�r�5���k�FU�*3�@�|BM$��RBl�J����`�Z���@BLQ"]��������_I3�[WN�C��Ӫ;�5���@�� _��P���
"HI�X�3�� �\��~M�ҙ�N�S�敥��,�B�}�IX�VBT��ό�U߰~"�^_V����-٘J��*MA����Ɛ�b�BJ�dT����1Z��H�u�l�/6�I���O��yCM��&�9��XE�)!&)"D�~��q-���_#"�ҳ���qK%|Dj�yf�<��P��",����|s>.�Ji�"H�ʪR$�\��Ҫ�J�4���
(Q��k�����1ShU���;�����F�7���e��Kx!�UG\>��W�*��Y�����+]�P�g�;�36B"��.|��D��E����E޸]�"�gHJ�y��_���;���g*�0�@ۈ@�D���Pۜ���.�T�uJ��!H�J�������+�X�
�ħ/��)�y�;��4�Q"R(�Drk�J��	H��A���>��܅�J�%-�����ۏ�$���Q���}��\�tn˛Z&�R��p���y@�<�="�]���ʎjG1�V�[�D!��%i�R��gf��n�`�@!Ж���0���d�lذ�.pL7P�{	�ce���^&�.��-U�
Zۡ�]n!Hmz��;1�ldT��M����.��#�v�kGTm��C2ݓ���	�����y�Y�a�h��&wh��A���-�"�cQT��a��Zd�J����F;"�P��ZD�sM5҃pΔa������P>~���؀ې�̅v%zך�G^2v7g����˰�3�����_��.76�
�f�]�e,e�m�?��]�&(�,�n�ȉ"}�[�����,K��q �H&�鸌D&B���Ӆ���

s�>�;��V��-�b)�(����`C�IwW���!ϻ��<G7$���V$�~zK���
f��(A�-$�Sn"HQ��후,׼{��Omɱ-'�x����]���H���M+!*��b���*�s�����T��G� ��G��t $��mj���vy��İJ�R"�L��9�qJ���jh�T�V�-��&B��S-$]�Ԯ#S��!s�BT~�	�U��÷�Cde�)��-�s�(\��"�I��P���0"�Q"��W�ߪ�j8B�
��dT��H�m��JQ���3�'�>�X��j�}W������L����\8VX��}v%%b��߮n�$��2��Q�B����Az�y����mV`����]`�@^{�*����~������=��7���R!�	���[��j�j��P��K��n�FDDӃ���Z#r����}��]�~��ڥUf5$+��XY&	.w�j�YO�8]#D��7�!_RW��3|�.�ho���C?|;%l�=��s�̥}��Ƙ�}t�	�C��2�a�QP�S]�&���F�t�(&n�L��f�:9��V�b�2I� -ʠ(���̪ Y�UN�����IN)�{?b��	Z�HZ�D]eT}߶�¹����7b�����Zrc�U�}7B�!H�qȡQ�%s�h�6�s�����؎���
	1+�h��U�7����9��[��S�B�Q1���Mܙ�
�uN�e��\����co^�Ғ�sK�H姲���7��*�E^VD2&+";�n���Bb����ED%���M�EZ��Ϫ��9T�R%�k{]|�?|}�Kn��y���a�T.�\O �D�u(m�E��Z�U|~v��w*�k�~��t��F��=�9W�m͟D�L��UƛU��`�����;72�8-�ܹ��i�Fg�j����Q��IP����Z/⨙NGQT$���~ 	����%��}��	F{���0�g��$�-�>e�_ut�mF�n!�	�m%���W�H�ev~��'3����qo���w�( x��Ȅ3�����21�\d���j���#��(���B���ʸ�"b�&l#�~��mM�Tkb������_&���.�`F����A��{�|#���Ra
յBAo�d�)n�)�(O��jt�7�Q���R�Yj�Q�\1h�h����Aun1���a��ˎ�$;0�gV[s��32+������T�ߵZ���.gn��(���x���#��/����U����9O��ί�$���B�Ȍ����K�"C�j��B���գи$
8[�%M,�KD�֩HS.~��p�������;�$~!�m\�ݗ�n5�(�B� �s߶mh�H�jB0��ؾ�� V��1���]�-"J�⩤Sxq}©�r��NI��|!p����
EB]���k~p����҆&��:��ӑ֔�r�g9�˼�� �T�U�8�Io�m8*���l�_eq}qg+oPw0Mz�O��+ak�z�
�[D<���l�՗�u�� Y����/����d
!���I|�>-%�16�4�i%]�����
����O;Ց���'�����n�3����8��Q�&Pj(_"G��m^�|�J�)�DP�B��Y������@�%�kp�i@�ێ�s�G�H�?s�GNE$��Rs-)T�U��"hrl�	f�����ң�4
(�,�����Z���U������D+�>4�?|E��Sn��$f�T7
�K�&#>ݫ]�� ��G�I"���=�E�bB0G�Q�]�������&�
\�a��u�F�kvG��f���i�q�l+��e�g}��H�q�VF����|�4��])*��:wk�#���B5�5�(���y��������vF����	�e�Ds�݋��ΐ������j��>ßL�S���,�TZRG�ǂϞ�����un��7���B�sTwA��
!)4���u����J�찋	�f��L;/���GŐ�9{��5oɟ��|���=X�/��F�G��<M�NBC�T�T���ͮ�X��	P��ݛ[\�VD��nȷ����_2	��wyO��$����B���-Kq�C�,��j�&(d���݉i"���"�ִ]�5V�}��&�$���ӏ<H?}��?}w?v�u�A5z!z=\}�� �%K�@�
?{�_�ơ�z� ��)�*�;��%�U�0}PM�n|��z�����l��s�	�\;@�EV��%^;�Qܹ�+��s48�z����*��QL�ܫ�	�)i��2�HgwC�be��%�\ږ(T%º�,H��	fA �$;�a��$
?$�/F0z�*Y�H�Q����b��+ga<���Ec�"L��&.������"?'Bj�w�VKXB�t&w�	���>z5���Co+����m���� �2ι��ʮ�ڱ�yS����ps�փ�ш.��r{�}>~gB��~�l���U���
?~���4uGϪ��G5�m�ŁL���ժ��	�V��}ܹ�0���dhKk�s�4� ���"a�"��@WP��1�х�̱H|���lTb������l�^ߢʔ֏�_b�|��C=}T(�eN��	�_ȏ�c�1;����:��bP}O��Ϣ5z`��� �jvH ����$*^	(҉�ԑزkΈ�}*���+�
ih���M%'>����ig�g;��d(\����@��J�@S�b�1l׻:��<��lQ�3��L�"Sr!��^?P?	�
��K{�� Y�w�U�#�E�����7�]�{��F��,"[ N�Ҷ��?@V�j�eo{'=�90Ĳ�e�$���D��d2�4�� *�d��������J��ULsN�a�U+n���[A��ۿ;�b�D�x��j}�<D��x5�*��_�������+�ߩU蔚)B�l�#����o/j8($KL�0��|���]z���+_�����U��&�� ܥ\�ǂmp�W�&�ޭ{mJf�T�St��:�v;I4N��m뻤W3�)E�w������ƛB��U�k�Q1VT��M�[��c��z��먘��o�e]�k�΄2g��m:.p\8��S�6��ZpU�rd��ӣ��k�s�޻�(�+����BF��A�7��:��6��*����4��M��[.l���.����x�9�e���j�q�n�5u�j���[R��'*��s8��W8���`c:��%ൻ"�J����t���b.#�،����[��ZUn���Zy����U-���7)�d�4k���$�XW+!4�#�Ut�kвk��K=?�߿K�1DE�2/��|�w��W± ��E8Ɯ��`g{E��4xx6Q#�ʰD����"0[)��Wg/����h8\i6c�X���b������l5�^�U}�ԫ��D�ZO����"�{�K+���z��"�}�b��C6E��P
�Ћ�����?L{��#��{�5��9Az�=�o��\�	f�2�Ԟ���1ވKڂ��5dEi�!��˥�A{$����ˎ�ꬡ�O�Ͳ?\������
��F�e�'�d}x�k1�Gᕧ˵ ���)�������/y�<��(_=Y*[��1��5W��V����(�) cL�����GM|��P��mZ�f�^�Vza�q�ѕp	��}5 ����b�Q5'�/Zt���i�}��a��G���+�����L���}>,�s�5�YQ �#���UX�������HOz1�g:>ď/쉄�E�QQ�	{*��oFۙnpv�)w>��YH�U&�Dn�cB]�SLi'����>�7��,P�i�AI�!���N����E��?C	&��_k�+/7�=v/å ,����?���n����r/�ҋ;�<�%x5	l9�n�Ɵ��&���Vt��R��q�R@�D|���Z�ٝ��z���}m(<���;������:�3H�\���s#���z��G��P7�G�Ѧx|�u�B�̓.8|F���:�"@�Z�ow�|���T[�f��W�<{#v�˅O�-ēL� �?BK.&�v�,���VB2
޹v+[��hk<��}<r��.�D��L�޾2��'�Cz�ay����{65r�U4r3���}I�2Ϡ�� K��� 5��F0��w� /���EN�Nua�}{�Y��������U���Wz��
kE�֨W�!�B�UHh�������bK�/vh�=)ġ�9���!��ۢ^^;�|��^
�u�����*�2(�
 �k@��~�S`�J_vQӫ��;���H=��!ec��u�ؚ�D�0�,W�+:ܻ��ͶY$۰hGq�J�-��+j�基{1z}1�U�*�:����#N����ad^���ee������^ӧ�o#������&����b�b)P�9���� �NE0�E8o&^���/!"���Q8����� ��cҠPr��h����El�s3�#�?	3΍}V~#O�٢M5����=\�\���H\ăv��V5Pl5�'��٬��� ^��;��ǐN�o|e��Kf���I$�]�(`�4(|w�Bto�)�t �ݠ4�X��k����,u$n�x�9p��&]�K�ll�#܍!���Î�l��,�����ni� ���`�~��BC���H��y�ͰIQ�u{�b�-�o�p�����ʚ��,�a|LG�=�����ļ[��E�toz�����깚�0R�"�*%�]�]�\a�h���H�U�	���W���G'IAom�Dw�f��-��ƒi����[����-�>���Fnn�R��A(����(�3y4
M�t5��U3�ƗJ֡�Z֖�sz��bC"I.@PD����$�*n�S���J\)���{�PC�>�lS�S����J�}f�8M�]z,�Ķ���Fs��:{7�:��2ͣ"g��ou��d��ٷ����i��xx�)3ٽ#�>>�D����B{�.�?n�P��o4���1���AҬ% JN8��;�������Q�J�%�I��2��G�t��6,�wz���� b�8b��N�HI�����m�2�0p�a,#���JH.�H,���Q��=g3�a1�!+|�g���|U��[^v7��T��J��)��)Hs S1j�Oĺ����,b�󖭶���C{�.r��;�}�;H��np�)Z3i�����{f�)���=����r��(���D��K�-hTy��.xV�j���+��G��7\�cg �h0�p�s�/��/���X�c7HEh;<�������O;��m�qᖺƇW(�z<�|c\`�v�M�q�A��$u�L����ه^_z�`���z���I�Y����r��\
�hZ�b��󦝒uA�{f{Y�/dw���u␣�1-�cqص�<��gX��T��L�eD̜z�L�7��}K9�ZV�:誺�~�:��{��� K�gɸQ�Ed�͓�k;�D��������< ��W�9d{���D��ϯ�HQ�H��٢���
��@��XM��Lmԯ����gi3&	�첕@�]t�>�Csi�1w1]J�A�s<�X%����b$���Q�kgs��#*�n֌s�u�����f^X��ɷ/9\9�,J�DBQ�#�""���D%
"?�"!(�Q�"���DBQ�#���J"D�DBQ�#�1	DB��DBQ�#��D%
"?�"!(�Q�DD%
">��J"D8���!DF(���!DG��D(��b"���DBQ�#���J"D1	DB���DBQ�#b"���b��L����2��� � ���fO� �t�ǽ�H � �@ i�YPW�4
 J� �
  (ڪ� P ـ �P
P���_ �        
    (        �z        �� $       D T�"�d�^A�c�H@�eJ^,4��gOC"�4q:q�,d�x:�S�{�/n�V������%@�ףOZ&�/3Ez� �JUU�u:<ڎ�=4�J��
\P��U)�    �     ����{ed�� �;�kV}���]ڑ|y�z�;��󼽽��������S�� n������U��w��<@�ϻ�����|�v����[@" ���Ǡ      �C{�o����rz�ӳyz�뵩C���}2��������� ,�/a����M��f�������/�|��<��$];�@�zR�w��/�};���>�J�H�JSo��1������=��Q�� �Wۯ���|�����U�>m׶��כu��}�A]����ﻀ� ��}
ݛ�4�m���s�ק��|�q6>�x����=h���@((�}��@     ������h������OG_>��N����<��������E}o��W| x=+��}�}�zzK�����RB�w_}�2�wc�{h>���7���C��ON-��]kˢ�gp
�@;���w�v���^���� ��4O���w�5m��x��إ٣y��ݝ�����=���`�� }����v�y��+{m�_|Ͻ_wWw)�}�}>�M�u�绁�)�T *�  }    P@{�m������H�/�y����f�y�y�+/c�>{땦/ ��zϮ۽��S�L���/>�wm�����;�5wy�S�v�G� ��OS�8�����y��{t*����wk�ҝ*���x��n�� /{�mݣ^{{lG�ݮ�;�<:��|���ъ徽�5L� ��w:]��}���.�o�xI�;��yv�u�=Ԯ���jTT�-�   �     w������{ϩ���m��w����;�v븥�c�g&��� s�����69���n��y������n�[k���}�}��M�� �^�_[ww��!�#v׍�ـ�D  B���n�QEU�S���ztD��V��(��IU��G�k��6ʽۑ)#�TT<�(*��̫���Jk�X� �)WFH�'1����mJŪB���a%^1���t��(�T�!2�J@ h"�ф�����@a1��2h  ��R*���@=��I�Ԩ   JzD	)A@�2)��/��?3�S��U|��k76��z��aL���sF�wE>�َ{��j�(�����PUU�PUUQTj�
(���UW�� ���B�*���?��������32jG��2O��fQ�H���ܗ c����Eͷ�m�p������'Y�'��P��jx�'r���(VB�d��t'7Z�T���WN�4p��a�r^���%lŚ�t�������`4���;��0��]ҥnR`��&�Y���k��Wj���ۻĘCjeܒ"섅���{<��M��70Z�Y��*��n����K��s=@�L"�8)����[��X4C���袦��"f�V�J����7c)�HxN����֛��<L+͌�nƚY��R���R�^B�����*_Z�Es*�i�{�ݗ�]��n,��[L:�s"Ͱʻ����]ӏ!h�N[u�]���m�[Qc8oi0��kV-�e�b�ܺ�8�a�P�/ie�n�:,"7{i�v��ٗa�څ�'��2��Ҷ�h@H$��j�fZ�\��mfBIr�M��J
Ypf��B+���9V�n�����f
hz��L���W�DV+{%�BSGs6:X�[y[�ʃe:*^����ݥ�J$е�j�c�`_�"c��$����EI.��M	z�)QV�bӏv���	yV��3�r�zBܘj2��$��~�z�$�х�j�9C+--j�N`X�Z�`dnI �;�Yc/�ih��[�2-ʻ�x˔��(��RW#�D�R���͢�|I�Ⱥ���j����rG����̻3QR��Ĕ�ȳ�Gg�F��U�6�Ǚ��2��@D��>ѧ�����f�����1m�d`�e���1��f��רB�5�^�D�	6�c)�/r��k�[Q���2f���@��e�dg@�jR��(4��1uͯ\�X�8���V�=�CH{�	�d��w�����@W�½�>~�̘K��q�>��q���$��U��8R+�旕�5T�RS��9IYʉ�k) ���)T3#ւ$�x���tR��ǕU0�ZW��i�m'Gv�n���/f��A[�6�;ufn6D�u�d^n���Y�sЗ̩
gx�O^��õz/�y�+V�-��ѹ�WFܸ,�G1^�v���#[�1l�>�5ca�Z��뱀�%%�o0�9q|oSw
�*ƣQI`�˨W�*��pۢb�m��ŚM9��1jv-�����[lmM1^�X�֞�ca�Ъ�@j��Mj�j�֤rV
K,nZ;�*:���.���Db���:v�f�yt� ��ad�V����6@��3L�uӭ�mz�P�%f-�trK֋�@n��B�Y����xTeʶ������з��. �J���֬QI��)"��,&C�5i�n�J��F}�z�#1��zw.�ћJc����d�b�����AKt\8m�Ǚ5`'��3�67��J"���yo/r�B�� c[@TB����lCF�̘^Y���+ɉ���\���Gt�#J�)���[�6��R��h"�1te� yv�*�kiU�b���eѼr��f�w��%X�4�FE�ƭV{�����ٙj	pQ��Wjގ,��\�����[4
\]�Xr�Ǚwh�y��bE�7$�)��9-�����Q/S��>�1eEF`��8��։�L^W� R�� MW�j;A7U��d�xA��E�5��Avn��b�܁�^Dy��-��%n�Y��I��@��Yi�q��-˗�eM����/)"���P���%�pLғ�:�0F�c
H��[KM�0�*��)-�TrC�� �"���YPI�h{e�T��`A~��<��Ĥ�Q7U�s�j��s0f󉪙�Y�@ ���W�m)4v� ��n&vkDY�feE	 ��Bc/w��49Use�i0ާDtc������-�n�ի�����4�ܐԳ��/*a���6�ܻ��LP\��S%!X�4����7��eŻ���Z�%�l뼣LR�������4E%��ٙz�$��1�9���m�U��yB�h3^��JXܕ^FJ絔[�m��3Օ���:~H9�2<tl�ĜTf�v�י�D�����byw���嚛!l"�j�݅FbҪ����E��W�.���m*���ۻ9o#��Vv��ʋ��g=E�5��|�<�����Ǿ��q|�f� E�BrYů+��E0c�f,[�gL����a�nf�q��Nb݁�ٴ���@�N�kt1�S�#ڼV���<uOZ�H��jL�5K�x�6+��y�y!J�=�.��ڔkNk/J�0�E������c+8��C��������[��<���)����7໔�6�m5,\Y��n�C.�����`��A/��^S�S:ѺcR{�Xs���
��ĩ��p�p�n]��Pn:"��rQ�W�ʼŃx�X��G�(�vw�C!:�j����l��%'�y�tw%�i�\�f��� -�e�aoe驻k���v;Z����m��mʳK���`���J���)�m�ں�$cQ3�%��b,[N�D�|h���3GݔIB��Q�[�iQxJ��L�����6.�<�����o�B|���Zb���f�2�b��Ũ�2)yw�S9kB���4���Y�	�۷ ����j�Mݧ��.��5d�J!�ХQ�,��D;{��JO,���*���jh?��a2���>&wr�؅�GV�`
�N�@i�a<L�o1V="a�T**Ri�)���/e+wn#�s[���dݠ��7�Vͫ�M]`���Bm�Ŭ�y�5�/2��5\M�viU�B U��LZ���慖�mb��a�i����3] o�ؐ?cJ�\���wrމ�U�/M�hbXąѐ�n�,���J����t�&h��F�m��Y��B��N��؆�b�*t좲V�h��	��f�Aǣ�,[%`�ƨ�K�B��U���^c�3�+VQD��4s]�Mn����)��,��]dj[�9=H{����Q�A��A����t��᧮�+�jV��Ę�cs0�*�k����F��T�&��a�U��1ݙ.�+��]Zv�;nj�4m)+L�(��:N�j��.`�e�
�n�����E��d�������������і�A����!�n��w�dq\S>z���aҒ�/Oٳ����5h������00�G�y�ęQ�[���J�ݪ�w�Zz�	�.bU��e�S:�Ҏ��kh�+K� 
��צ�W4�x��6�:�S"�?@�n{ؖ��˂�ʍ&E/�z�U�*�EkfhXѳ�{J�;d@l�Q���9�ǮG���i����ք��k-gl!+CY�<f�ö`�ǘaㆣ5+u�|��ߴUkBY�04���uY��#��[u����V���	2�w��i��q����͡0��E�#3(532QR�����f
7{J�$ͺ�r�����3�f<����,: &q�[�/5�@�ͤ㨢w,��[���8���f�YqwyQV0(�V�J[1�Ɣ��}p��m]Z[v�ɦ���Tf/��[ߞ2t��h�	�o2�B~��ٮ���z��-'z'��'��Uy/V�=w$k0�C%^k�[��[ז�m�w��[y�#�/&��mTe�"�U��Rn^l�c='��WWt䧥nY��0)��`����n��n���l�LH:x�����6�պ*��u���CD�j���R�)���9[�[Pa;Mъ'j�4+�Yf�YԚ�z�����6�)�Ѧ�l�m�����QҌ�h#m`)4��"�U��T�1�{)�RS1��ygH	��h�ʸ�ŇY��1�{[��i,m�KY�Uz#�����G��ʋe��yZ�Z�VR�s2�Ą�wmM�fb��Y%1 �M������2�&�=g���&Y�l�D�j�6đd�u�B�ԑ�C��;�a5*[5,Ԋ����lyV>���ϼ�ۼ�$��6�	b0K���[��B]�ck&�Le�ͦ�³b�T"ϼ�Ur��"��TQ�z����6��Fa��t%n���dӱt�
��O�Îe�/-��1��))v�Adb�L�+�{��)����8S��[pK��{X����.+e-m��E��5e�V�{W�ڽ�o-3�[p���]�n�^ܲ��TWc�fބ�R%Dl=
�g��^�Y�YP����y4i�oJT��ړ�M�4��P��ٽ����m�����I���	���W���'��7��n���G���;�����t��6dGi�C�0D~@Y�U�f�Ȯ�9��e �X��$�݂�/i]3DA3QR�F�ᚁuwv���h��v���5�j�V^j����(��
]�M�!30�+%@F�{����(�K2��M�[1�j1��u+`�Uf�d���'�4ثY�0��c/e�P���9����^�n�NG,\]Qʉ�r�U�f�50fJ��n�koL�lj[�3�l��ޱ7
��lPZk22#�g��e����JVU��CU��ԏُ]�ڳn�!���W�����4�B��{a�k.C34�[�[w��
���P
3�4��(Z��iGw2T~0`�.�^:p�h`6��L�n�[;�/�%Js�h�4nٟ��q���{{X�`	y��j�`�M�Yy�Bf���kQ���	n�[�GOX���c�ҭ�N�7Z���$�X������5$wnP� ��ܭ��kwf���SDf�;1ɪ�,�̴lj[����b�.���j]���y�e��ܿ�X�⺊��n�gU9��ni�,Xw��6�]���Ki\!��rdp춵F"��-�l��[�w�^�qa��3N�>�yN��/S���P��Q��⼡��9{��^/-�6�!��⶝Ml������ĸ��T0^]����kRݱ3&���9�;�v�4`̷ʷ=�����U}.eo�4S��8�K�t�7��wPٺk5b����m����ұ�zgan�'�Zؓh�EJ�K�Cw�~`�38͸�QD���!��u<�b�v�"
���k/�i����9e �{X(IlMܲ]#yY#YD�]����RfǍ� �H+��CQ��V(����un�¬�it�j�)<�j�h	-P�&BP�.`̽-�G%<�bg��uag�R��b����cL��d#l\�;Z�N��(��@ͣf��*�5�j��&'�x�#�K�L��`y��&;���!��̽Ȳ�1i�^�NB�@�T�K�NYS�Ҩ쌱Fj�i]hf��M$��ڋ,�5�J�[a��,ۑ�̦5�64"�f���K�
����GF�[�\��	JRm�B��/2�1�\q�5t)#mf���fVA��,wYxNY��W�@;3"Y�%�eǖ�����1t�íe�� 4�"�XF� M���w*�M�]q��- ����JZ�pٺU0Sw.�Ai����sv�Y��l�\��P�FQ�PZ@QY�BF�C"�v^@]m^FJ�0�2��53UY9W2]֨��&~;c=t��̱Yy��B�
�U�v�T�*oMn�SN9�x��PÆVl��t*��T@d�M˼6�qʻf6r�e�c�+Tw�^�Y�µ�nfn��rU�KTё;��c(�//ױc�,k�ɮ�V�\b�/u�e�*8r�����In�
���F�$�q�fRɷH�V0�h-%J����5L�lU������G.�F��fm� �
��X�g��>�Hr	`�KY/)��i�F�*Z`��ֺvl�WyL�.j�[ˤ2�.�!R�\t�Q�y�Z��"�XL-��.���i�K�X�5���ͼ{C1ۗ��N}��Rf*�&C�\z/^ B�4�b7[.�&]��/-�7�%忦,T���n��й��4ΉP4����+.��Z�Wv�Eq����֎7+t�X�DYX)�
��lb��UyV�ˎ@l���H�lR��<��2�]3FLyi�H7lw�E��E�\L�����Yt�(iY�{��Ƞ�jN�[��ם�*�����x�<Ĭf�7�D_̡���[�vndD^\������j�"�!��3�ׂ[�jxh�����D/��6�Ub�}�� v�@��h����AGh����I��?�����a<�/��7~�t�,l�9�[f��3o#�\R�2�7�uk�k1a�.^��ܻ��d]���dPI��V̀���PkD��*����*]w�����p)t��2t�!:�BVIf�j���*�Q��Q�b��**����1֜x1�����k� &b͌&�\ߑ�j]�0޳���:�F��Y6U闙��n�*��Fll��]�X�"i���elIp�F��6���b�Ҁ��ɏ�b�mL	��W�ʇd��S	��䭗�u=�q�,x��t�Rf��Ι��� �7�R6B`9�s"�6/-fP:�41����P����Z��/s& mZ����� ������Y�\��|�gQLjT��$5Ev(V�y�� Z��R�����7xĶl�65a�tVl�p���r,wXp�7�m���J5��[
��IP��,.�d��d��YJ��(��y����[~�Ÿ���j��VT����3oze��=܂)�c� |53�� ��ƣ��F�qZ:�0�aƢ�ݨFH��ղȺ�!D'B��q\�CH,��`�|2���"��W��A� ��#�f�Ԩ�����+D4�#E�[��7�� ���,Y.�:_SMZ�ll?4ǟ�9�>X`��wN�捱��+��V����ã���n���,ݬSA�dÍ��f�6�-噔(����!��������R��*���~�_�u�����������\�f��̓��MN� l�ۛ%������nZ�Uj����~�/<�=�A+���MI嫕V	P A�F�@�A���4GAag�yy�O*�e�ʯ�a�\�/U�tv:�;u�u�9:��up�"����$�[<�g���cv�:�!�kq��M�o�`��}˻uUu�v}�Q��������sA��n�xݝ<,u�{��N:��x:��=���t2��`On^n�#���`TqۖCj�9+@��/�1��c�s��q��j����n%&A�0X�j�y2J��^����8��vg�<ȬM7=n�s�����W�Q��c�k�ܼw;�Ƕ�tq��%mr��A�nݹH��7R�Ů�-ɺ�����^�cs ��z����mc���(��݀��?Q��v/�8�6F����Nm��/��f���hr���:�wac	+b\���rt�<>�]�0��+�.mذ��!�؛n#A�x���g���&�N��:dB�vgf/dx�]<��Ӛ�h��KX}k-����O!=/u�v�-�^Da��P^���xͼxǅ���t"��9.z��%�[�Tc����9�VNw2�9�=�%�����q�gv�U�;	�k��f�n۲�u����(�"�%���p[�.z��\rz.�5�1�6��Icd2
�{]��L��܏[q[���׳�#p��C�[kw�筹����n;]��'����LZئ�]�t-Լ�X6�d�S['��w n[�W`��������q��D9�z�8���z�Z�����-X����[�����)�lV;s�n=ۧ�/g�b�c��)L�u�Tӝp��L&�7�e7��kL�v��C��p���ӷ=����']g�<:v��[��$�<�(\p�ķ*Y²��^�l��7li7
$j3S];-Y^�J��Uـrû݅�1��S�O+�9�Tck��;�b�sۗp�ʰ��D�0�ү0T��ɛ����c�uq�O�\e}\)�/sz��g{N2tb��@j��v�U�7�����pVmыgQ�s�Y�8�:x�U�=���냲Yl�[��*cc-ګ �يSO)�ζͮ^9�=��MGl��s;�ex3ݞ|Fp�o��T���VӮ�x����1B��{Oi�{������nv���ګ<�Z��C.뱞8��g����SY����v�<��{&h�ݱ��k�������%��Z8�\�-�jį67��ss6�Oa����֭`8�v�O=���ۣ;��Ctq�
���Ol��a�[68ˮ�;t1�[!���h�ѹh�k��M��1�ݫpdx�k!���ɀ�m��g�t�s���s[�U��͹4���9ћ���..����wm��Ӛ�ف��da�.n[�	&�Q�=�#qp��x]��ú�ؙ�ݠݹ�nW�ݶ8��W��Y��o9m�y�N�������n|�a��;"�]j�����:{v�]�9�q��X]ٖnvM��6��gf՝Ǯ�l���0�m�8���\TU.�3.��;eHt[v=E��Kv<T����7kvщ�N�<1�����\W��yw�6��z6ض���m�S��k�E�[�;9�ڮꎰZ�s�K5[�r�=p�*��6�ní3Tn.�6�=;�l§Z��85u�ø<X��jrۂ
tp�pX�]��<b7�S�g�N5[�GA�fĚSy��7Z��m��*����F�ڰ��E��\qۮs���8㎯7;\^z��K��ǩy���g��=���⹍�n�SP��U���k�j5��;�7.(y�I�U������ka��s�{n^w��l]�*�.86�m�w^7`��Qά��뗞�d�p�&鵵���7l���7��B���n��ne�2)�\��L�g�7f{Og���� �;f�t�n7Z��ܥrԽ%��d�kgn�dMn�8+nU�b烘b����e�)�nwK��8�2\���pGf)[
���8�q�偢�i5 FVD��h���W��#*��C2�ݮ2]�;ˬ�3��ǭ��9���xx}n�.����y�!��|�uq;�뎂}����ܿ)�<$>r[&P݋���i�x�:��[��N�����=�7R�cM��gq�ۇ��&^�9���Q�t�gqX�Ǩ��H�q�H���Y69�擮��{��o.sx��:�g��/:�#v��W�9�ew��1cL˖�uq�R��.ݱ1�36�:��h�gj���m��պY��̑��v��8z״b�5��S`ty�'�czM�74��ms7[^�QX��a�/�R��ۜa7�7kk�J��<�n֒�s�N{pY��y�k��۳�U�n�Wd�[��VKw!�9�����OmzwC��\d{=�w��0ב r�j���s��������p<-��f4�����N�k��)�`���^v��ګ��GO�ldd�+w�;��h�vǻJ>zwI�s��1m���i�e��k�g;����J۵m��!zj�\baz�j6�Q����[����^]��&�����&�whV��2g�vi�z����g��uE�x3=6V^-��'ní=ո��S��\h7+q�6�g���)�7Tt#����V�i�x��n+�F�u�S��u/I:f�n۞���s]��tn$m��u���qǎ�#��5�N;p�ƹS����k��(; t�W3v-�z�u�]go���ŢYb���m�2J��]�v�F}l���oV�`��ӹ���h\:���;\����z=�{;�I��(s�Fe�Ӻ3��[W��99Vl��]�:Nݎ)���e�n�	�׋���2r\V�/��cWn�ۗĖ���^���j�#S�����Ce2���z��s���v��]n�=h.�CGۊ�Cjrup��^n���ػ{;����\nz�8��9k�ç����Y�ź8�ށ�maq����ضzn����V�%����vl��#��W.u��&�\f:�<���\"Fо�K���ۡ3�j5�Nu��X�Ϸg�mi�f�k>:�v������S�&���s�v�w��y|�g=�=�<7�ׇn]��B�V.s�Ht�i��=�w;���K���`wb���ZN���������g������DwnMe'���m��Kxګ���=P8c�8�:�u�gnš����+������zݑԘ|������b��{k�˔�ܧi6nx�s�\�v��t{m���k��.����J:�U՝;���GgݸwAS�I��3����]m��mO����&�A�ڇ�upx�]v��A�\c�N9vm�mc���p�x��R$RY�\�h���X�M��W�x٬������Y;l=u���Kv�Xn6�۱���c3x�y����͖a�m�CƱ�������c��vy}n8E<��˶�c*��n}�g���'���ݵ��q�9�SQ7bą�����`��۝�sխ�n�-�ݓ�E�$�λmgrlM�[��.m����;mn����[�#�e:u������ə���v+i��g�]z-t=��d���N�>�qL3����r�X�xE��`��ca���\�ษ�'>'���Ļb9:�6�l����1�L��nz�O #�x�d=���s�ެl��knw8��vk�n\\1�v7k�N�vC��l��t�ܝ���yƺ�td���5�!����X�S:)�%�nk�jѱ�vV��kk���Ƒz�ME�AN.�y|�:�q�i��<,=����)nV�읝��׮^x�`]s˯;<�X�����n��Р`�ݸ;܆Đ�nmY���R�7���9�;X:�4+l�c��I��=;����p�@�u�1���dzHM�Bt�j�c��px��x�u�T�M�
�E��^tj��f�NӻY���Eۊ�{����Me8w]��R�O<��o�i�b���Ywx�7e�\!,@k\��:1���T�g��:����;j�65{h�ș��<�����r��ҶC��v6r��r<l��v�]���W���[��E�Knl�^�;�QîR�Q 긯v^���Þ,�p�3�F{t�tc�����v��Ů���P����;����F�����|��nk��8LN���n*�92�f��Jp{���ۮí��L�����EI���.�k��gt�w��i��{u����jJg�Tm�ACm��j,�F�{�v0ryJ��8x�)��Ζ�n�<�q΋�w��c�v��R��m�m�]F2S�������� D�X�l�648�'�6y{T��0�מ���x���I��2�j��@Nø(+���.2y'�;kL��x�����v�B1a��6Wr��ǣ�n%Y�e�Þ⣑�[ssڍ�0u������r&ci��u2Q"�v��Ou�\��ɺ71�-�6ćj�h�Wc��lq�3��uf�����nE�m�+9�����03F�Wb3����F9@��x���۷u����X�B]�y��X��6��ױ��z��0�ƺ۳)���Ƹ�n9*�sێz���rr�bW=m��\�nz�nx�3��۵�c��]�g=v��ۭ��-�;�u'6c�cm����7�{_?7�>�v3��{f�(g�Cqʷ<��sg'����sx�w2���v��c:|�+g[u�v�GU�a�����q��s���N����mY�Q�q<�5ih�C�OU���\�23��`q �b�ô��q�9,C����O��������yh�In6����k�,�Me�v&2�Kn�,�i̻����	>VÇl�b�n�N݊Ύ���ݶ��ʝ$��;�lӝ	��m]Y�����HW�mQ��/:�h�]��w_����B�uO�:��s'6��a���q�^$^i	�Kø���m�]�q��>���>A�:�l.ƷP�q���cKv��y�K���g�rqW ��p�=xx�O6�'�wc&1Л^T���ʔ�O>��`aܮ#0�]8ݸ,<��y�q��n�f��� ݸ7&v�<�J�=5�O[��u+�ίj����M�RF#un^·�3�J��q��˸{>���V��UUUG�+tUPUW������j��TUf��Ȏ]�	��r�,��1Yݎ�A�y��\��{pg�4��te���k�z�a�79�py\�\�s8��V�8��U��s�Y�A[`���>;N��UЖ��sn���.��dήՇn]�S�dk�m�q��f�]���u�qn�wf@�m��f��W]�0��ns�D�:�[�����<]��gן!��[q��&n�\]l��^5�m�A�l!pa6v2��8�ϓ���]�f'V7m�'��Z�\�9p]�5&	ۧ�N��p7�vN��<��	8wh=m�]�8��wb�n'�79��Ie=Y��pqΗŞ7k:3��.�O�nN�Ω�Z��eC��:I,x�e�xvx�bn�:4��rgH�|񵍝hy��V;[��;=IvMqւ��s��n<�����;E���i{q�}��u�m��s��p�>�d6�{v�2�w�չ�/K�2\rʼ��!O�:���#r뇬=9�'c��t'�X���9�U�Ź�E�fۋm���gh�� ;�Dq�xwF9�S���-��j��T����!p���y��Z��^7�c�V9���i��y��5k���9��tm��z4r��.��c�_W�m۶˲C2�#�E1ۭ��.�5���듄�=�s���+��v�D뵕�m��gV՟Z'�c'Gٸ�f��]v؃�;��͹�������mfc�m�Tz���v[ۚx�x�ȻmN��������k�l�mq�F$I�p9:͎5�H�^�� ����`ٲgcq�G�:�g��
���q����8��;mhB�6:=+�%�NݺNglίnsHp�8��F�����K�;�>��q��'̽�Ñ���s�[��б+Olku�7���"{n������O��9���0Ss�G��l���ۺ���-bF���\<�pq��f*㝇�ml�y;���ۂ4�V�ծTG����+�2���"�=�.bо�@�m85G	��7c���L��Ȅ�c�QAA�D ����(����B��h*�*���zw0�7y��Yn��:�Ù�����Ht�r�ȣ�P�q�vpk�vX{rSrs�g�cc<�_pk�c��Cӎ�p�.T�aǵ�ۇ�2&m���sru[b�֗�	�#�l%�Yָ \���c�+�۶=%	�T�qu3�9F�j�\��8���gX�Kr�i,�z�u���Ӝs�:�ܷ6�o&�a�6�jMu9����aEFԗ��b�7d���.�=��v��w&�M��e2��l�_��h�֊4��I����(-\k�������^��
�%y��z�'��]$�8��b�g���e�;�hq�\�j���bu>w�̸d�K����rq�j��Z��s��m�T@e]:ƫsf��MQ���ǚ�<B��|͑����^��]{@q�*��J�J�ɭ�m�i�7����wz�ْ�'1Z��[63;V�l�9�/�kHs���W��4���'$kdn��z��G�|��%W�p���E�\6_w��s�J�LA��
ҥZNr��<�]�{3Dj%w�tbTh�o[֡*���9l �?���J�s[�[f����X߽��5�͵֪��+�����O��,�� f���w�9��p�f�����տk�ܡ��G��'��@��>�5���tq���p�2�V���щV����8��z��F8骴#��Ӿ#w�1��P�*W�~4��!x%m/$B��~�9�^�x��-�Q�R*��� �W�u] ;J�P�z�6�gq5��u���B�,2ea�]��jag����$GE[����$zwlw�V\�#��-r���(u8��N u�^�곲��m&�msp�i$�8�z�{�ǩC%b�F�Z�[�����C��Vns����[4{��Mlj%zJحV���ݹ1�r�[&^^�F�� ��;�D��(�b;V������6�B� ���Z�1r���c���yp�5�Ͻ0[���5���z휰�u�	�j�� M[��(��ѾJ��4T�*����{xV���kmGodw)M'}���u���o_g�w�-���b6]zM,��)!$��Kmm�^�zi���LC����t�V�5lBN�V����ϙ�Y��2=R���V���k|��buģ�hֲ�CRV\<��U������/�tN\��a1f93׍�@5Ut��0�u��XͯT��m!�#RnP�#���m��b7��o!c�E }1�c��x�?66aֽK�b�٣Wւ��Oʽtha �����Öi�&�}x���I	����y^C�o�5�1�jQ����s|��ZZ�s�V&�/;����܅tN4|�o�M�d�ףF��1�4܅u��1����Yr��rQ�H�z��k���g/��w���i����F�3!��pE��Nݹ���N��.���S���n���\:q+i����)m���V��n{%v�q�ivÏ�5&<��q�W[LH�#��"*����x��O��l�/F�%/�$3۞4=K廓��|���t���V�$�K�k�KUl@����� �?Co7>uMӛrڟx٢(����w=�y߯�F�7�'�H�k����@���J6���;�֛��4~`׶���
�P��u�'!�V�W�~��va�y��m?&5]���4��������ҫ��v٧HmS�o����Z3�aR��s���Q���yy�����f�O'%pU��Y����Sf��m��9 ��#���4��췍^�+{tX��ca]��i�w_K����u���
�ԆPK�w,P����5w������t�_9��\&�]�喷�2^%i��,n8b;�����o/��{�v�h/w�4Й(�ү��W��m�R5>��7��wU*;�W�V���-�)�t����쿥�n�
#�mɈ-w���&[2�Q&f#Uyv}��V}�ʎ���^�1+i�� � �Qګ���_=��X~���t�:L=v<B���U��sŝM���Q�d�9�����d���Z[]�����g7�zZc�%p��W@�e�O�a�7c�5Ûs{uӸi9�n*�3�=��͞،u�29/2}�䠏��Pq;7�6���Ʊ5ܲ��;�ߓ�{�m�2>��UC�(óࢽ�g�TH��+I��->Nv{!y:{��˻�U�mD��9��/�x]7�.�30�N�;��u]q�]}��Q���޴��+�χ���}~�[kmU�o�Lr����毳�op<�����h�~�S�i��nh�f�Y��y�괋Q�N�7f����8fK��xӝ����xB���z��; d#��D-_*K��~�����gz��yZw��6�j��M5]|�-�y|Nr��OjQ�����Ld��[���q�je�#U���v#�?t�Ǩ�]˩�E[`D|4��z�k�Z&��R���y��/��Ʊ!i��tߪ��ٳ�sd_X3R�	�vc�s�.��j���'La�r�YKtsk��J	b��G���� ��]k�o�4O�Q�޲��J��2Wks�bcqV`��+LGҶ��h1+�;����1��51��	�
�ߛ�ħ~�6�N�kH;���y�F&��\B�k��^�k}ۮ�1/+�y+�mm�rɨS��>777�H9ȏa@����6����y�+3�]�sgy� ���l��Qq��K�::�>4��#�oӉ�旗t�d��N��mVO� _����w��k�R��'��M
�;	�¯���U˪W��U���%�k�f4]vl�B7�	1%��bq��\h�%c�M_������k��ԕV�skHz�����!"�{��}� 3� Y �N�`<_�=�'�C?Z�V~o:���G�བ�r�����,KS�Op��W�0(�q�a�#�YpǺ���Y�i�kP����h��{���|��V<L�ﾽ��˝�����6�3��$C�گ����o���u��l�^!�K���Z����֦�hR��
�B/�����A��Y��'��x���?:�!�
�F,�'�FQB��C�) ��l��4�����!Fd�R� �ԍ��պ�h�����g^$M��t���]�w~���s���{kMU�bz�$B�ꧤaĀkʩ}d3�Lz\7K{N2$��_3FC�#�b�V�V���J:�k"��_����ƫ#k%��������m�M���a�rY�(p����`����M֓Ϭ�M����;�.@6�C�}jic����%���r����qf��)���4��G@cW���nQ�A�U�69�u�x8�qXqI��:{m��m�gŔ�C��F����������i��Z��^9�����i��d*[N*Sv��y�����H7��/���t��F�mƱ��ݶ�i2Ƭ>м��㓛�?�ɻq��g;�+�vjF�m��[/F�<�n8�Tv�G��N��.���nϓ�۔+V�������9kuZ���+]�NE;.�di��N�S�^4c��~�c�q����v���j�5o=:�/��m?k�;Yﲢ����?a��~��X���w��z��$"}�~C�i��6�k��"�h�Ь�����X�{sWeQ0t@��X=���Ƃ'R��̥�;v���Nw��r���A���cE�٣Te­�4-G]��W���>O!�,J�ן:�3��dǿ]�s�|7[J�f�7�|��n��M�K�J�W�m������tP���և̏�S�>yo�.��*�u�_��mV��f5��sU��ܚz���J�J�q��Β�<k��+�b藗��c&���oR����w~�җ����<����e�+i�i:�����M�i�o~�Q�6��˞j���&����Dz�h�-�I�e�簶<�(l��B�V����:c�">t4P�cO1K�Ƹ�x֓�1�4���"N�j�~G����SomY�!ksyIǭ�-�h{z5E�Q�B5mF�����t�|�i�Hn��p�����`��|���2�n�3*�lp�ɸ���N:ĥ��9�����:��nܽb맴{Gn���E
����k�ZHko�&�p1�&繕Zj�:�)��4k��u0���<|~�d
����e
cF�Y]��z�C;���\�5�E�i^��jћ���v����+���±��G�C;��	3�+�a��G2��]�kwT9�5Cx�A�X�p[���-:��8��on�-�ޗ�a*������޹�mD���n���՛�y-��Z��Shm�D�F����4k�]B�"�-��氭�k�������oO�ƫj�>�Gp�bH��f:�;C�rc�V��;A����Yg���a v/��\�`a������泝q�v�'ʴ��5�Q��ᶼE0��Y���.uqѬ�i�>h��&��ԛ<]�Yyh[���C�?^))�D��[�����%u:�o�ڦ���&���q3%y�}V��" {a��n�0�T!-�j�p����kþg;���Tk�ߗ7�>�]Uu��ŗE�VB���M��m���a�������
�r��HD���J�{�?Q15�@y��k�Tm<�ng9�7��-:�Ľ@�MOr��N�{��t���N�L��Ljʼ�p�~��j����m@Ia@�Ev��Ɲ���n��{ǃ���¶�H]�7V�M�]h-��a%�V��v.=��W��ᢌ}p1�B���wZ�_ɶ��д118ѡ�\��k7��]�[�(;r�>�y�&7\h�P�i�~ʹ��˶Ԙ[3�q#F&���^�����G�o��f�t���QЯ��:�6� YH�>�F��e˩�A�g�V�6��n�&�̚�k�v���̗�K;������|��q�\�Z�32�����^^U���q�%�ry(W���QƻsI��{,�c��Y˄|mG�/,z���V�Y�O�}^�6�M'�-;��f���-Q�W��JҸ�"�v�\�m�9�:>���9��J���5��f\�4"y�>�g��m������u���
]>�+�+���7��m{p���/͹p�Xֵ*���Ɠ�!��	�$jAxl�@��0��5HW�j��R�#�^l�t��G$<�d߷�j����h1�U��~ճ��"�?v�#���wgk���9����@�[^z����O:����7&3feѷ�F�d���{F��c\N���z=S�z�M�p�egӟJ-�ehh]:q�9�{F�=x�b�8�_'��۩�N���5{�I�m�Qն��'������Y���m�q�XrN_o
@p�\S�N^��$����S���U�aˍ��uB�zC�jt�_Y\t��]W�i���Z��p��ӏÍ#�0���~���͎R��6ג��O5~���s��/�+Ms�]k����&�U��&*� B�א;W'�F��3���}��o9ۋ˜�m*'���SS5+�шNn�j��or�����IGɏ�։ɧ���l����%w@�Y�o7�������U�9��s�ʗ�ۙy4��16�!�'�z-�Q���͵�J�[q�>a���];�����q�ncy�7��쿏;���LCY��+M%��e�H�M�^
6���~k�G�#-|(�&�cxaq&,��m�ky+�i�}�����n�4/����i����!�q��z�u��h���啦��kR�1�p�RE<�
'���_
 ^-�O{
�~�/LZCʔ�S�Z׳��h��0���j�U�o��iq�ĬR�T \Yj��|�h�:�̊�y�#ZF�� c���R����C�1<յ�<ܶ �ߤ9p��QfH�ۼ7�GZę4�lcv@�q��1Qc��h�]YX��ׇ����{�a��'Zƻ�Zh��\��֕�\��:J����tq�D���4L��<����i��5b�k)+ν��/<snn	�	&9�x�cu�;�'m-ˑz�<���۱�G66w��te^[�p��[y�<����}�cF�I���p�[~~b[�m�ӭ�����'�ud(>�i�+X~[@nl�����{����>Ѧ�v�9zAO��i��w�'p�'ZM�}+����a�32�Ye���A��Z�_]������;)�G�Ds��Wy�,ӆ�Gġ��L�n�ƻ߹�TI6ґ����B�cĉ;�����ԭ�v�r�M��ֹ�UN4w/�g��5�l�\h��w�/��(7@���H�=�m�WI�8�y��&����4z�~�m�n(�s[}3�/���:эw�o�(�\Ko���N�웇�w3y��ԭ��9�F��Kh�}��ccx3	��5F�5}���M��{3Ҵ�+�9(�l��Y�Y��۟��IG�kW+�s�uG�(��ֲQ�K�ܙX�__�%u��F0��%c�ӷw�/��g��_��H��w�ݨ�=ˢ��U�!����'g��E� >�m�B�}%|�_j#��sN��������q�rF��ùv�̺�����v�4��Qn1�ch-��f���4mn{%-OM*u���3]�V�(r�BڈĨ�~&]��^C�M�p�:%��e�ñLǛ>�1�����L穿4ج��]�Ñ�IW/�N�B�ȷ��dc0c�{ft�v(�Quw�(-�������Qo'=n�s�{fC=�S��lv^+x.��[��ݜ��\���\u���Dvۭ��\����[�ss�@\ޭD�]\V텧b��]�j�Q�䭟]oZ���&qmm��q]�Oh�y�-���w�`y`�W ��+�ݎ��\=�����<��[���`�6����vͶ��+�8�sM���n� rRӹt�:�e-����.ݭe��`���]<<�9�]�4�h�=��rZ���[\����kn���*Lr����������F�����oұƋ�#Ϳ�ݾ�Yތ�0����4�C�{n�������$�Di@�ʭc��N�:6��Z�!Ʊ�vܣF������ĉs����kԀ�M��<��en�=��-�w���&�m�j�3����k�y�M�sI�w�t�}J���Mh@o,?�vЊ8@�ڌ�>�V�����qƷ�44kT�vv�ј��IxkY���Z�,���.���ݟAyV�'�%�F�Qb|׳Y��jf�|}p��줳�!X!b�Q���	#����y8�z�m˼h�w�5FnWɭN��_uܖY�	v����CA$�lZP>[cmW����ʎ�d.ڸ�.������MտL���g�.���,R<�.�:hnQou~�&y�j��o�n�Z��$ި�ˤO1W#����Gn۴>�[���4y��/��.\ȸ�s/2l��C2�B����eu6EA?�|[�����%o*�g��@��e�4D�ve��l��eʎ�5���s~�k�ޮ�km[FԽ_]��ѽG*n�̑�.�ķ-s/��\,4K�E�\K>��v�<����[!!��t�~�Q�l>��O�@w���:�u+2�)my3ڼ��y�2H��C��6��Es����4��F�Z����^G]�_	[N;m��JR��Zs�Fa&ٖL/&��[Ak��y$�X�&�=��}r��|���v��q+�mZ�M?L�6U��m�ɥ\�1�vkՍ�pl���ޢ��Z��zK�i�Z�E,n1��pg����:�p��S�x���$.����s�n������/%�ޜ�-�wW֍�}p�B�P��{�8҂�zv�==�wS�r$�k9>�H�.r�,��2]�K��m�Ԛ��֝s��o�ޥ%�|�������ߺj�ݑ����W�UI��I�Q����[ZN�כ�Ƹъ�k[�a-�^��J�G*�������-"}��;K�=�C�wu��i�q��� �#A�_']��X��{گ��x��)K|�Lc1�f���I�5�����:��y����{�j�4z]���Ҙѻ���0��w��	�^ae�������((���($��H���<���2��0a�E�+�U!�ۧ����Sҍk��3a=:э��� �z�����'͂N/���|*��NwP����A�z�����L�Ln]�♖)nf.��iF��c���v���TzS���y���J��p�e�c��y#�ƌ~�bi��5M��a���a|@���_����@g����N��8�?
��U.LH����N{Y��J�w�tf�S��m�hc^�ƍk*r��eܼl��e�]J�Ľ0P��s=5F�^����ǵt.��aƉ��(y�F�j����-�}��h6��V�ՄCN�:�ؘ>_Yd6�[wXf6ퟑ�<C<R[Y��r��2��D�o3Q�7�cF'���/W�}��k��cG�x�Ģ&�ݱc�� ;y��
��=�������v��3p;��͸3�)���<(6��@�e��L'sMs�����A�uVv�Ǌ�L�	��2�k�&\�'&�����ʢc:���%h���I�l�"�D�es��_;��`��ѢE-��-���I�}��'F��GZXl��W,���a5����}���4 o����b	SF��B^��V#���/�c��޽��ۍSx����
�Y�3o|o1�#lB������U���x��Ҝt�<��-�6G���Z�Z�׊4Pw�=�Q�z���YQ��%%��f�l�v���� ]rOjz�Y�=����z-�I�a\[��&*��6����0k{;���ͫ�t�#��]s��ۣ8���m#���h��Ϛ:�orR�d�F�K��ʯ-N��s8���E�š�
ʅ:h2a.%B��QVm_����⡙,�QZ�[�!f�<��h�V=��������,��n�I�7����;]���s�`��a����q�)�^A�X�c�r����+�0E�,hZͥ؜[.�*�t@�i�us���e=6�aΠ�o5��<�A�_I���"0Ն�r��4:�*�/dRL���gLc��^�+�Ҩ�~�����g"�-��ĳ\��|�o��ע�mÂM��y��\������+N�*�Z�It�����*b3}r�P��Tow�W83�PQ�(J���T�1�g/�]yؼ�*�Hs-֘��CD~�4�mVӷ��<������$>
P�
P�~C.-�-�%���4P�
*&f�J7%h�B�)X!�����m"P�
Q�
�4D�R �(� �$h-�B�)F}��]�J�J��)B�)B��2rB�(Z�U�HP�
bJ��n�B�)B�)F��g�����/!��]��J1*%
Q�(�DJ�M\J�HQr)B�)FIT��-��㺉B�I
��)B�}��h��tcX�vo_�H�)B�)Gd��#Zj�P�
Q� D�J�f�p�J�(R���h#��"P�Y��)B���եj���u�B�(^�(R�HP�G戔)F�(R�(R�(�w
��J�J/5�׽�)B�)z偉D��J�)F�(��
P�
Q�)B�(�����3�5̓���([h#U��P�����+�D�J��)B�)B�܅o!B�)B�)F�(Z1�'�(R�H*%
P�
Q�:��˩yr.f6Y2^a����҅��V%
Q$(R��{"P���@čh�B�\�KJP��D�J2@�TJ�h��-��3|�^��C�Q(R��P�
P�
Q�)B�-|�G��~��J�J��P�o����w�smVډB�w�����%
P�
Q�
�J�J2B���4o��҅ƃ�
�JH��r�g�V�)B�)GپitP�
P�I R��P�
P�
Q��9�,�J�J7!B�ܔZP�y"Q�%D�J�J7�}�7�6�(P�TM�D��(Z�ʫJ�C�p�J�h�B�d�E�D��)F��F��)BյY���=r�9���}�-�[\Ȳ��K�]�\Fz�lM�{n��)��8㗇[n����ҟK!l��q�w�/�B�)B�)G�
�h1�B�d�
P�
P�%VnU�
i%
Q$(R�(Z,h�G}���B�)B�-W��5Q(R�(ԅ
P�
P��e�4D�J�$(ZH�F4F�����{])B�J�FIU����(�DJ��J��(��?J-(R��P�
P�m"Q$�m�%
P��{��P�
P���}y{J5!B�)B��"J�(Z4��(�)B�(�wz6�rB�(R�(R�3�h�*!�15X��)B�B�nCh(R�(R�HP�
g��4�
Q�%D�j�Q(R���ϧ�d�.�c3p�J�J��)B�F%
Qr)B�)B�\�[ԫJ��-$J7 }��J�h�(�?wK��*!�(R�HP�,�{��^�7�\�U��.��(�)B�)B��Pw!B�)B�)F�(Z�5V�J���oe
P����5W�]�P�
P�
��o!F�(Z%��ġJ9%W�F��D�J�!ˁ�Th>bP�
P��3E
P�
n��vB�(\h"P�!h̲�(R�ƃ.Uk�V�)GyvH�jB��(�J����7��(P�TJ��)B�)B��js�Z�(R�(R�(܅
P�
P� y*%
P�
Q����'L���KYd���B�)B�@�Tk�
�h2�
Qr)B�)B�\�V�J�J��ݔ)B�-�˪����t�@q��4Pc@��ɬ76�U�T(Vڠ�|ʪ����5UTq�(*4f������=A]J�6��}*��mUU���J�U_�:�X�o�����R�����
�����M����+�UV����4|���U�R�q���X�~{y�/�ܵ�� J�U?�bX�Z F�Q�g�_�fk�槀��5G�*vUV�_}�l�Q֊�E4��A���j��J�7��������R�
����- ���6�
�_ߺh�T��(:�hnQ@��ڪ���U[j��4f�k���Վ�uxV�:侕x$��i�4�w	�����P���֙��E����y��-2�ݭ. m�s�	�A�{/�/;�ς���U_u���K,�"��B���i�R��
�C���q�;2�Ze���y���6�Z6�\�]m(4��{����R�G�ߥUnw��h
����~�F��������b�G��x��Ibi�����y���c��0E�)��1�J~5G5x��q[��qp�H=����V�%��[����va��b	h����Ƿ,\ӻ�r'cBS�`��������vE��Ԛ�k�3��+���4Y	0���1�R� �[�s�j����Y���]7gl�`���!D��2�A�2B�	D��f�U+����`��Y��OY��sP���BF����G��;4�[؆v5ldV4��da
�x�!�϶j�V:�C���zʄ��zf��̞�-��
� 	��#�<�b�?V�Ck�3���S�"�aD�˷էoT'��e�k�+�A�l��O����F��*8ہGp����^>[�~��yO^�k6�P�� �Y�]��������SX�����|�Z[��i�w�Q
^8Az�)�e*�ӻX�cQ����[��]ʀ�Ǘ�)���;���C%�m�ǫ/T'�y�(h1��R��^����WZkb�.S�jh7Y��xئh]�G���a����7k:;nxw+v����F���y6�q�T�:���wTe�i�m���s���8⣓z$ύڸ{8Wh��W\�x{6s;V�ps��k�Nݝr6#c�������m����v�{ �G$�k��q�I���w>�P���b�V?Ϙ�8O�6�5��ǨZ��;8�m�m�wI��۴�ц.�,���d}��cv*(���p#>�Y`.�ǫ9ۀ�S�7yP�z���n�{���o��{����5�Ӎ��{s�V1������b��O�/��E'�����h��"��Θ ��L�N5�9j�0c@♐*����êe��HJǷ�f1�98E����Fԡ��1� L4���N��P���}��e��)���,�pSS�0�F)N��d׳��sM�vR	n�I��]�M���73k&I��L=�0	\!��Mu�	nkǻr������y�}\W������p��C��ZZKz蓎��4����3L���vJNj$�p�牺��v�wL.��}��/��*��q�K�S76�2�.��
�y�S�M����{�_�,խݗm���92c��h7m�h盍l�a���6lr	#�Y�J������ՙm��
�-%�]�lnv�ij�;�㵼ݬ��A��P>��<=�$%%�_�S���k̀������&b��j�7���<p����t��9؛���F�N��k×y��G$2��}�c�ր�/\���[��h�]��8kE�ܸ�P�X{*,uZV.p4
����Y�[yкH鹅�3o˵��y��W�[\��z��mLs������mrр�jG���7����Qt�[<_QF����f�-Mk��aH���as_6<j�3\�9k�$ ��M8u���=����[v�bPCN��d��^��5��s�y���X��pj�k��=���9ړ*q���F��Ñ��E83^XE���;*�:5�t���R7f��a��5o�hz���7~��_���֬�n�O�Z3W�vd̡S��~��������]�d�7:�ɶ���b8l��8ۣ
�w㣬[r��&�k����tJ��k;�;���%ho<.i�y\�}�I��R�*�@L1ؓ�}�`���/�S;��U�2��Q�M-̛M5����p�-��z��&g�t����[Q�r�3;��Z���{���ӗ8�/iL3[�ĺ~-���~X}hPl$�GŹ��H�Onr�k�[��HZ�열"�r-�~�0�k��]i�]hԖV�ئ����	��+U�ѡ�w�4﷝�XJ�²T�J�$[Y�앦��A����/��6n�.���U��}1z����	������q�۔����Z�dE���
��xs\�|X�ZH�>֦E�hw�b�;�ב&[4�v�v�޹���s��{���}SM�6VZPq����L�ɘ�����P�'j�>�)b��:2;��Aq۰p]p�ul��y/�mm�&?���{4���B�X� &�ג�|O�H�b�m��x����V�#��X�>��¨�m��R��l(��U%WA���m�NyN��|DU�x�p!�{}��a/��rt
gY{DH�y�O]w{~C���!W/�q�D�%�BͽM�6+."��`���W��J�����n�����x�V�О�n-������ޝ�nҮ�lH�M�&@�b�L�N�����;�=��ws��Y&�<�1Qru���'��mw_�k���+lS�*�&�V�$���%I�6��i��t�z����Ư�+vv��.�R��Y�mt�z�(���#������6#��R(�1�C��m�1\\n�*�Y��8�v��`�M6;]k�1�K�m�+�����/یC�o.�u��P�\�p���1ld9x�4��N�ѵP��ҎmXgy��	��w\�g)����m��x�ۻ:��5O'vu�q��6���T:�;xN���H]���I3����Z^z78�P8{v�J݂aR�aqOl�t\�k�]��D�2��#öNS��J�X�Oo3��;��x�J(ư��Y�t�w����:(os���R�K+(.w:h���c�#��G>-hl�o�z�T&���}�*���2ū���p��{�#׮�;ۂ����"���X[�������;E�i��]n�<>�3R�tUX5w1A�CW�x�Z��S}dĔ���܂�|����F��z����t����e$���ͪ�Rr.��6�,X���Β��`�W]�e�� ��d��o��Q;���ˉ�$XF|Y��a-����J�usM@͜�;L4!ot�c�u���a��N�-8-��
eu0��A���U%V3~���n�Z:��k�f̓��V�aMԊ��c���Ю��u��0��#\:u��l��z��78K�����/���C)�;�߾��x{9���!l��p�v��y{F��):�|�oHG�WBfǢ
u����]���t�A�q�[��u�mg�i�Cv��ݠ��pGv�m�o7q�md
������ڦ����km�!�ΐ��9��=[Q�7_����_�Rtj�������tq� �/'u�欳l�ikZ��V��ؖ˅s�Vg��Mʖ�g���>+�$��Zn0=8�Ux�X��ݵ��m�5k\��q��}{7��D�p.�-Ks�ϟ�b�^�e^�k/�nUH�V���L� �:�y��or7w~�����DL�w��-w��
��+!wX��mV_��r4��gN�:|\�y�.�*-׶�e��FK�w��,#��s���Ѹ=O�X��$�)��q8,xy��
w��w��u="���t-���YuW:�\���X��s�ܻ�H��kUU�9�A$P0`	1FH3�e���k�"�%u���_�f���D���6����[�&�f�U�a�/Vu6qTm�:w���@ϯ�g�󜱋0vKIE6�A0˒��!����/��.�#�a�h���JjnL�"t=]_3L�e3О��z��^�űY���`�<Be0�G>&�y�z��L���<�xζ��'8�u��h\�D<���+�8	ȋdR������|�<��ng+M֦Q�9,���y���g�{$��6����]:�I��҄4I�8���]kc������YZ�^��R�R1��nJ���b�F�)��jI���W��E�
9�����kU�S�9�v�0��䝳8j��C���Y�&{:{/c��K��"��@t���������<�x���}�&X'���"��NA&u�%*%w6v��+g���.4����R��H7��<�=�[:0�U]�,{�۹��,�q(%�1����m��}}+u��ö��rj*�vI&U���i�[O�ui��m�M�m�<�ܦ�g�Ӓ�^A��)J"W5зi� ��84�D��3q ��x�9Ʌ:vR��ސ�xdTӶBsrk�`��N�5�.����G���j(*nWqm��L��ۆ�ǟ6�玓�![gԘl��ڴ��vK,DaQg7j�Y�&y��N�Z�LhP��:l�'S���GC�����z�,y�"GZMyj`�h��%�b�����W]�:��jv��7u�kO5{vf^�E����2�&H>~�,u<ٻC+h��S����`�'��&2Y�E�QD�I���^�b3��j�o,���y�R��,Ɨk�=�q��%Et8G��`Ҿ��=�b�{<iGZ��Ve�Ʊ���ʌ<;e=�'�Q̄�W�L��}�OH��Ն��.���za%��*��6�������Cn��ZⓉK����.߃O��Ǳ~�����x�|ۇ~�O]�{��T���VxS	�b���1��q)f(xT�`�V�3��yy�v����2JF�<N���%����&�.����Lc��4����G�R��:*�c��w�];X��Y�z�:ذ���6���퓭��j�"�b��Ir�3�,�]�Ϧ���ݼn�vBB*�i�e^��m(�u����ۤ5l��c.��^||�k9�V��L�k�綊��>q@`N�0��T����ɍ�����)��*5z|/����+\(�܌�md�+�!���x'7�a���p�&�6Nĸ���{
�ma�RB8i�Ȳ8.������z5y*1`}=�v��[�~�Hם�ɽ%ʡ	��p�CN
/ޟL]C���je༵~���F���9
��+ř��~�7=ɑ$s�J��ԉ"���nq
Tr��_��R���T�s��#gG<�V:��\�9L��\XD�`�����l��UZ�z�`�V�yB�ۖ�p}�,�w��X���z�O[�^6�IU��}�O��֮�)9�9U3A��*x	�S��2��
��-�®���c��X�=�頫�6
�v�P�Ќ(R$ָǧs�[��bU��Y[$p�v:r��[v�<{�Z���D!UYhM7�-�w�5��N��|���7�=ϴ4ڹ��k��e�B>�Z�=ʓD��	2����*�҄k�LGl���s����5Gد���k�7�)�m���L*�k)�Q2����vF�������w�Q@U ��V��-wY��wy�����o���wR;��ȳ%�9�o���Ӟ�5�N�;�yC�\�P!&vf�����w_TW��Ȓ]����e]�]�	�+:��z�c�� ��%�L�S�'&/�܊��ys���a����x]�/�Sn�	DrJÑHF$J�R�YAL�{�8z?�nY�:{q۠M�͡�w�f�Ҥ����tP�ǈ/�E?g���,6r�$�N���cr���[e�D)���N�n�)^�Z��;l��ݹ���fᔲ�ɷW��䅎�2)a�iY�j�¹�C����0� ]�V�Iԕ�;�3�o.�K�]'M��$NƄo����sg[�l�.	��HYwN$�Yˢ$��تh�]Y�B�z1������tJ���.d�e飻7�����\��JU�d}y����A{��1�َ��qJ����8\%�9rx���XLjo�/	�|��lh�#�����;.@���!��&����%N��Q��r�갣�:�]�����ڼ�C�)oF����l�f����[4��r��fgu�g-�.���s8��5gb�6���H���S9�&\.�����1�e�����RU�6��&Ͷ���ۦ�*���]]�
@�Y=��l��En�xn�8fRK8a������o}5}W�a\,�7B��r��|��8x:��/t�_�eQ4<������P�SI�nK#v���,�*�؞�خ+��C�%��cӼ�c�������k�p�,�A�U���[񟙙BSZv8�@GA�:䪔�b���j�r��څe��7yX���{��=r�jth�oVL���NVa��E�g]�8�q��ȥ� ��e������4���]VJ��Y8�J�vΉӂ��+D�r��H�(1�=����s&Z��+�=��5��&���7�t��4���S�����������
�j�d�إ}��wH&�%��v���;�{Q_��U�ye{ҏ��b	&\#�N�m����ۊ���kɌ����l޷�Б�1�%�nc��>�<�>#��=���و�m��Ba��Hٖ��6峏�p�OHFM���Xv-t���l�v�u��m�??vT�(y���v���x��:U��=�n�֝�/k��M���W/m���S];����n��㮑�Bny��듎݉ _l��y��N7i's�g��v|�N�eq׶�q��i�����n�[/6ȉ��qqѝ��/v�Gpv�4�x��u��¼�]nx8��:��cM.8������NN��v=�սaa�s�=��8\��Z�nDvm���� <\
k��;n��`�����6����9N�v��q�hga�U�3Ru��mٶ�#�yv��h��8WW(���>9���W4ۮ�眙�bH�L멫�ۧ�7X�r���ȓs�j��Sֹ�p7����[��usA���O�Z�Y7�q������z�`V���3�ͯf����]����8lv6xцf��/�s<��qϖ㍳v���>9�9���[Ü�]�]��
n�s���XnK%�Y+��6���s��92�:���m��v�'��4�*�i��Q�*<��ݍ����%ڳ�YN���AV��
�Ѷ�����]>��Ϻ�ʗ[u��`�G5���l��c�:���4���vݺ��v��Wd��19�<�*jsH��yg��,���y�� �f��[c���L�e:��t].�vݦ�<s��S��V��n����s�\kc:lO���
1�q�9A�L['[�8��E�Kbx�u��Z=���u���^��:�pctvᄮ�"[�㣱�m��.s��ϵ[�g��ܘ㍊XL�qZu=�v�qk�w;��gccT�:<�sV�<,�7x�;��O;`�l���L�cm�q�:�jE�Y��m���v}O!;�ݬDj��V�9�ym�-��v��?>>�l�6�&"d�q����+3=�m��s��eήъ9a9�v�f��k<�t�������u�T�:R�I:[��G�i5�Gh�P}��"t�6���;1�rOZS؜�M�÷oh:p`��,8(`ٺP�g�)����ˬ�fɵ]�H1ӻ[>�Y<*n��n��>�VȖ��q��l�ٕ��m&�Qȷb�
������ݷN���z8��lYvx�^6�Y����Yt���f�N[-�7ifv������;vLX ��3�:��ؔ��G�*7nSxջq���/��!Ce�$��'n���^�� �&�'�*!RL~c���%����K�/sC9p�V�S�<�s8;�a�qY����:�jG}��.
���P�V]m��6��AjG�����.o�a�t7;�+���9� X:���͠�SH˝IyAI�e�]�zu]j[��^5��<f�On;g�#��-�Vq�r����	��Xn�r~[&;��+F��r�F���Q���5��zGٗU�[�����=�8�P�T��Џ4w{��y	�)̥�x*�ӹ�v�z��,�)�:=��yi�����̶��S����{�*ؓ�R��1
$��c�ȍ�eUWe��?b�|�!��tW'��\�zjg{�����h�4���#M^��	��!X[}�W`�{�i��a����T��2��8�/j�����{A�;{]x��mc��78Q3��,P��c�!(L�s�Z��ǽ��b�'^�~�t���s�Z_���m��=�+����	�Ǭ�s�udF�w��Л"ʀ����+$���������Q�}���[F珰.����S:���lT�
g3X�g��w%ό9q��Kc|.uo�ːi���j��t�9X��NM̝�V$2��Ƚ���O���#8�5(Y��g����l6��مz	DWV@���P�՜��]L�|\�pAM�b�����w����f�N�vd�fm�����-9]A7�4џ6ɂ���k�`na��8)���ܩ ���0EQO��UCv��"2GC��n|���x`*�4gw_k�އ�k���9{�M�
JR@�]��V�zp8�Ω˵Ҧ8�Ԋ��p�V�������2u%DV�dK8v���Յe��	�˂�v��w݉V>�Z6>h�C(5{��n{>ݺe���v�	�w�)ӧl=u�x��nt�; �Q��L��=UTd���^3�[��ה����:z"��Gt�}�n�o���;7�c
��*�����łt��xvUaac��XRF{�S�\E�O��R��W=J����f<��S�DB9a\>��7��[R,;��z��V֋!`��9�@�xlx�-��0���!�b���t�&�o�iC�7��,�¸R:'n�ֲ�Q2�U�G��`Y�CI�v�H��:tJ�����c��s|�瘚�6p�V�jќ�m���=�K.e���Pb���Rf�DjG"��XL�Mls����{V
�&��^7��DJ�L�v���6�'�@�j�Z��J����ض�ki��0���`�B�i�ኰߚ�?F2�f`8�R�>�0���wxϚ%خ��β��{҃���B]y�J�R�5}+��׹|��i�s��2r,��Լr�ŻnF�	���V.�!*�����!�#*m��3�HM��b@�I!��K�4j�+ƌn=7zX�mU���u�����gFZ&�3�g��]㩸E�xJ�L���ooJy9S*��);�nf8<�N�劃2��r�u��E;n$�O ��U՟kC�][�/�i�#��3�ჭ�_���Szj�����D��(�Y@�޳��m�V���s�#�|�Ϻ��#i�hٶ�4�"��9}!"�zQ9�W��5wtw���oAJ&�Q�^���&ܞL�e�e��9��ދ���D�у�V�	l��nP��`-l���\!Uɵ�穎��}/6�P�RW�m,��Q���U��T1�2�RO����w��l�H���w�+{YiYw��+�6ȁ�qr?�F5`�c'�GE*�")]�h��:7���ϥF���Ttmg+�~�ѝOƍ�U���b�C�ܥ��P��T��r�6���N*�M�'k�n���)�n���=�xwF�#׋`���ǐ�r�F|p�I�m����#զ��½��{�C2j�Of�n;��E՜�Ӿks��mI���̸�h�{���ds�������m��2_N����������uhp9�xx2���!R�t��ş���5�&�$E�zǹ�jsԋ�!dw���뾞I`�kJXb����^7�O=�<���O=Ix��z����w�T_��v�\��Epc��Q������Ez�p���
^���"�Ж�aI�'�_�����u��,�f��<4qƁ�|
T<,)�2C�|&G|t���wO�ʒ�S#���4�P��or��O3-t0���Ŵ�, Lqo���=~��^�O�7Y�O3�.�r������&�FtyxY/qx����w`�{���v�.��-<�;^:��I	�3&W���b�m�=�ӓ���U�@H����e�j��Y�R�>�(����ŮL�v�r�s�3$S��il����ۃ��un�i�rf�ϖƳO��X&��E]P���s�۶3b�g�[�U����؊�=ٝE��N�c�v�^3�[�<��΅v�Y�g�P���[� �J���,��q׵�5���^2Jh�z�n׶uo����}�58)39� #�GbjᲽ0
I�vyݻ"�@v6@n�5D�McV9v}�ٻ8�[�'����F�U�x�ݻ6�n���J&�ٰ[lq汷�:�;v�R�h7�B�6� _~��e�W韞��*%��{�<wxw�Z��{(�n�nϮ�W���vzp ��;����
#K�j��h���M��� �8a�����uy]O<x��C<����x�����H�a��y�r��eNON���ޛ<���bDu�I<[y�����-)���B�h^k���nM0�F���)�͡���T34�t'�4���K%m�r,����QG~����i�O��e���e0đ$��cD�B�;9���V�!��y�� �}ܽ��|�u�kϧ�OH��W�<B2��3%�P��/kA}���UD����bn(��8�ȳۛKE��^U�vk�H0�ŧ5j��Q8x���������ʳ��,&��|Uի���L[U�%�������f���&��sH��--�&�t��f� 7�5�*�ni���;�Ȥ�I���~�XG�*�\IＬZ:�co�XDU��a����{�h�~gU��Kn��*�·O.��Ds!7�<ϒ�֢��AM�e�e�XWv6<�FJ�Εk�L7,pB�4(��5v-C�V8��°���.	��)Z&�|�Ƽmv�h��Ȇ�u�y�U͂�ʶ����6���j	�}�V�V_�.�=���b�Y���͂�:�'1���{^����Q�"�&�-��kֺ>�"JfJ�':��!I���zy1��sʋb�н��`ڦZٴ<n�y�JM�@yCP�#�V�{(]���{��z ���o�����OP�`�Ji�E�o��m����+p�҄�-��R�cM�[���;w���\v�3������w��m_>�(��B����D�2-@�mU��zx������7��Hi�k�޽>��fɽW{e�����^�����lys���jѕvɹ�0�,��s�R�9�Փ��H��Q�W]��'��y�1�u��3-g���mo\���g���x�6�JFݮ@ױv�yH]��4~.ʜ��	�*.e�p�K�S�G��Xa(��X�Y�T൮�ٸ}�k�q�>8j��<�ɗ��^9d����˖�x�{��������ŃY+�u�������mx�<
���Uⱘ�9	��1�{�����<��3{ݺ �1T�� AځȈe��R%����^���~��\7D�ù�u��<A�Ԁ@�<�c4OE<Q�_N��v��6�W-���%gm{쳯}���t�h�`P0�=��}W���i�t����ɸ-�̷��ܺ��Y~9�(e��'�wC���%� ��r9�É����Kv��:Ȟ�-z�<�"�iN;8Ր��3�rY��l�	'�$�e�ܻ�v��K�DeFd�Ӹ� �,O�)�c�,���E�}��n�vEZ���I�Tg�9���_i�?F��%��a�"�	:�5Y�3}eH�P�s������Ǭc��H9
�b$	 ��=4. �v��8��Nv�2�ĉ�ޱ�zn��ѢXO�'��m�@Is�ۮ�0j�ܺ�}��ң��"'Uƫ����ʬ\�H�;���3ݹxs��c=�<^i��g5�H���qS�`�}y�K��MM)��1ynM�\����?{Ȗ1p�^�8|D=X��}��^]�w��t��Ȣ��=�D���P��A�ũ�-�O���AB��fz�g�4�jz�E7f���|NP^9!O_�&��,�"N���͙����Nn�Y�;̕e^)TTOo �����*2RN*bI�����N�X���G$]�[��;sbbn�y�D3�%eay*�.�R$U�)7Pi=�z��z��-�ݖX�1^ּ-��s,S����a�b[�+{e�g��h<��W�	��̜�!�`�Y6��CV��p�.	��5�lr"��]D��I;oG$o�u�M����=ﯕ�*�zT݈�j�ʴt�{r��K�(����9;�]�L��G�"��k�y���5}tMB�/�'��lg?#ȬL9��v����4N�/07mڌ����{w�G���v"�� �R�� [KN�lU���nb.��pqZ|���ӪY��3	�׋�rw����id�a�(�2��B�S]�x�7N�5�(ok�Z���rF�X<v������I�bK0jD��h@{�qi:J�&����:��U*!&��n��HԼ�Ʉ��OzyW�{���W�QI�V�Hn+���2^^�<Q��^�������	ƃ#)zД�	>�.�����R�ND� _T�V��+��˭O� �w[����qoڠ��ûz\�q�I0�n*�Z��Pz�n<t3��k����`���D����_o�'�����&�4��mm���W�: �H�[�._�[��r��D׵���Y�l���'a!iK#��f���{E��fA	;[�b���eh6,�r�V���t�U��*����0�E�� t�u�!>j�c<����-�>�����3���zt�tݣt�8�wz�O��4��L-v=�=+z�}�	H�|o`��r:G6�q����J���8=��2ov��룙i��r1s#�4䚸oO����F�36�#wd�ZΨECm�����@ָٍ�����ƺ��,d�\+u����e�5��v�cd\����mŹz��̐�Y.##�MG=:��Mn�������q����w����Z;k���pv�k^��ۮ�m����͎2]�+u�/v2����Ѵ��@��4�U���v�u�A���v\sl���']��=�1�kS�<O�zMȕ]���N�8�C���u׎9������o����]���n�!���3D�u������6D�7/l�|50��;�V�bT�o��^�"����g	p��E�\d�䬼��I8��.�'F�燺�W�Q~֙^��X��
��w\'�zCnI��V_ɗ��ݙ�8�ɾ�{��vu�FQ1�Ou�8�k�$�VSv��2ojs;f�n���`=טh]�Q�E�6s��M�yE�@ �lKޮW]u�{���'���>vʃ^0�D6��T�r��1�}*���e�R���3V�C�ҕ�o&��eE�������j�J�94��a�T��q�.+M̟q�NV��¬�@���R���P�8���a�[��u�\��'����D�m�����l��Q���ٌ�Q�Ȩ�5�:��1��PC����c����٥u�,s;ڻCt�it(#������E{=˽������<�^�w5�����a��*��䙋�'�7}�kmw���Ⱦ˶*7�������Cz?\� ��I�
]���qq�}ӄ���/ w�<���_T4������8EU8g���AH��>S��V0����Sr�Փ��Ζgj�����&�g���	Y-�ٮ�k���,�C�SY�����km@.�Xt�������ᖺ���)OS���e�z?O����yh�=y޿r��:*��~(�vq~`ٱ���w3vy��<�8/.F6�*B`�xe�[j�A���L68��&���UҠ?X�:b%�Grf��K�Յ�HT�v޿�zz�L_ՊiMg�O��۞����"��s{޽���#�L��*ޫE��c������k���	j�W_�a4�g=cڻ#Qvq����+�!�ILέ#���E���)���E$������E瘳fz�R�["�,[�tT/c����v�����^(�|<�՜}hD4����1�`��(�k֪��LJ�w-?=�9�
�o��c`�,V�@���p!w;b�w@gR�dwsd��O���-�.�Fb�F8�q�5]�Rv?f������p(4�5]8�����d!Y��7Z�ڋ&�����rdV��S��Ye6l�뼙p�|��H�}c����H�������.��R��.��&]Y��Bցg7*#��~��S�=���_f�י�'$���0�-�"��X���
6w����Jw����27�pr7#qв=�B�c]�ҞGܼ�z��׆��a�X�k􃦪��+P΃9m�_8΄�a�!�ie��6�f�q�s�c%�;��EC�n �Ҁ�����U��Z���̗f��
��V�!dN������[�[9W��*h�ַQV6��h44eM4��	;�p��9�N^S�ߎ�ںB8F�5'���&ohu�b���.]�s��+��r_Z]3]��N�W]HoWY�De���K�Wp#�<kM�\�r����M��k)w7��L�fu,3�����2�nD9��o���ub/i�u�ovJx��Z�s����w[��t��l̬�0���-��.��fH�:�FH1`������	c��+2�)�e��=�ӱ��'/sy��է�2�V]es�k�dZ�w߁���j8��g2:��T�R�c���a:���D��ew;5ٔ�B��\�"�=N��X��5�:y�z�3���>m�wr�31�(HY޷�d��U��z�ѭ��l�y�$�������٣cX�-}�~�i�L3kP[ኔ2���M�[{�x*1ʴ^˖��dz�=������SS�u�z��̚]\+g���XJ���GU7�p���X���f欲]3��xz���F��hx6�N��3��s�<���y[y��>I=S����<5�OI�ո��^��3[����{��l���:�8ma��9�ێ��STwD
��#*k~�r�fԽa&w�����P�H^�s���^i�]ߦ��h�5�UKf������BP�3)e�dU�}Ҭ�T!DS"KQH�,���*�e�ȯ==��9-{!�-��-j�>�YtH7���cu�?R��;*������Ѐ��aɹr���x��|���� �Ĝ���=Z�$�ɒG3.�e����
b�B�6}�컻 V[�Ƶ�;'��d�(���f:΂UR�q�]�y@N)�:C�*�a�0�R���f����X!����ߓܒ��Q>j��[}I���x��ts�3�:��Z�D.���u/;�x
۠�� ���jO�j�U�u�����|��f��g����_rƏv1DѢ�W}+�����|��k�B=���׋�,���ˍ�ۑ�>���f9-\��S�O�x� �GU�*����ʧ;����}H9��GЍ {T�a��\���\�KG/[��
������K���gu���̞}G��[�S|&�����D8I�$�C;�����@�^yU��cB�Y�<q�i�po���8a�z��syR������{�����yƳݬ��oz��m�yم�$���]�����9"G���YSss �2��C�;#.g�sж�j�t_ʵ,�{<�'^5�"�#�Ō�W�<�-�q��:�T%��2^S݃�%�AP�n.˽�
�@\�WЕ\fjU��^��A��VW�p��~D�j/o��`�<nb�F���2=�Q�须o-Ř���/gr�s���[ʿy�����Tdƛ֣�}���y����3R�}.���F��SR��?*'j���q�q_6��y�6�o����9�O�a׫�M��۔7<T�	k���X�t�u8��u��9�u�I��*P�?��>P=}���#Ԃ�~�c��"��ӗ�l*�+�68h��ݞ$1����H.��G�쯷�|���%�Ú�L�sX��k�ԏ|�(՗�-
#): )s(��fzo�!��^���s���隚�]�\��������gs��}���֑���J��iG��J4}l�����@>d �,�ē1�Z}-<�q��|�7wt�q�5L�V|_g,(%�~�� �Ň�hG7ʅ�����#��F�%��y�Tl�4�������&�5�&r�W���[s�@��;�b���=q���������>�s����Z|���/�y�U2�����2�Ϭ-v����ҍ.ذl�[��5<��aaS�E�'g�`�F[Q�$��,Ϭ`��T�o���f[*��:V�}�{z*xE�UEzӒ]My�#%Gйf9��Ũd�0]ܥ�4z%n�V�2�t��P�-Z�-dH����
�#��x�]��e6^3s�	�	�졙�d�+�3}*�mV�kj�I|P,�����s�Z�s4�Vv_O�6����q�=�\���]�\v���<��s:�������]L�H�<�8�c��۬�ޠ��8����E��͍�����vNsN.q���3� ��Te�,!Fu]n+(��<G =D���ݒ۱�s۫��Mct�Q��6\��r�it'��^��'X��.R-�ަ܎u5���w��]\s�[f�K��[�n2���n�(ZsؗHq9��S�M"V�������|;z�{�'?/Τ������X%f; 6b+�G$�x�U35X��w�k-x�C?��Bff�ы�}HQ�Q�!(�
Q�䱜W���`��J��|�mgݎ�������"�:�FǼ���uLߝ�{��A�EDlP;����屺W�(�7�n�'T��3&�p��ad�w#��c��EߺEW0!�y�ʾ¾'���K�}�/���{qC����~�Q�9���1bt���'��00z�8��\_2{���5��[%����[,�͵��YŋTs��&E�^vNؾw�Z�麗G��J�=��b��Z{�r	�W.|$x�?BN0ep굘p�����!�um^�3>~Vs�Ze�0�e���ۮSG�����-�>�83�Q��?u�Nث�����K�Br�Ɔ���<j��U�Ɛ(y�R��k�t��8�k���~����I���S�L�[;U3ݝ]e�Px�����vֱ��d�-����2����ȟ�w2����T3G���w)��N#�����g�d�:k�Ӥs��(bv�X����:�����VK�~A���V��TBh@̐��_>֡��r�u�*� q~�}Z��=C/" ]Y��xk�y垵�˰e���I�t%��j�8RH*�W�oóX�F�g=w�r��.Q�T��:r5�=��f�Ty�Kj�\�(�va�p�Sk��ͿN0��5�l�\&[�x�-���9����c�hH��{��% ����N��{�W�Z��װ��9�˳�� �%1}�*�M�K�7�
6Yf!��Ib�����@��C�7=��Y��:\�s�+FQ�bg�]����/@�}5���R�Y����Ơ�͞���))�M�V��s�7�d-p�Fgw:��U��O�cK=ӹ�S^b����M����b���]q9`g�K�T��������4	y�������������oUiH�0�L(��w���Ec�^�ʏ.�U��?XM0�	�Ӄ� �ð<�s�YTnw�xl��Ɲ��ԋ��qGkn���HF
���J��//����m!�H�W\9W{���v���j��yuC!�^�ֶ��lo^zo�I����]������K����mg����d��7�klK�aK�0^bÕ��2���`�@�#����_n: sXa�:;s�#�D,��Q�\�r��8������&���$ߦV��Z�Xǀ~���$<�&E�˗��㦮J8�.�s�����,��Ri��M��gdx�خ���~�sKX��3S>;�a��X�K�����YY�7K�U���ۘ�n���?��-um��jZ\8�ҁ�D�ۦ.k��|(�p\
��ߍ,�氌�9UKU�9X�wٿDp�N�X���M��������R�i��5�gЊڡd�(��v~�|�Ax�W9qK&�ni$ϡv�)�d��18��5� ryz�7G]�m��Z��c��<�)k*�R�J-�`�O�@6���8�`�ԃ���?FRi���b�'=�^��}��7���������y�g� �j���_����)bvbm>����������wb-���o;��W%�ԡ8�srO�9nI���ls��G^�l ���������	�>C��ҏ/W�
���Q�� 6>�A��`%��O����[�]�l�����V�W@��3�\������βn��X�J�+��)h�i����tY�]cΔ�ƽ�c�	�#L'�ׯƨ�����?-Am���e��"�Uv(yLKI�����Z�y9{v%֫ff�L�����F���D���k_�#)
�-N�ڷ���eҋ�h�Ҽ�ή���W��[eaCeeB~���Xy}	 [��Af���0�F9}��E.�5�-z�Q��2��ig�<ԺܔWҝ���;�a+Jr�>��K甠��f62�eE�zp��x�?Y��#�a���9�bp�!
+�Lc^zv
t͛�֚�앸'�&Q�Y���8�%]L$�z�w ,������t`vBEi�͈�rG j4�r��@~���j[OlвBX�DO̩Cq�ھ������08��[Nг�+� �a�$~yLU#ޣ쪈=x�[Z�WJL�Ș2���Ʊb��yG��-������m
7G�Ȯ�Z6�_"��'�H�.�v���o[ K��(��i��#�𜆛"�d����vY��DƲ�Y�Z�{�F�_�,�C�J%U��&a@�ޫ;�?��w���vv/���.�!=VRL/Y�[&c�W!�~�޻uĬW�Ϝ��!4K����^�g{��L��/��4��a��A:���?5e��$_����q����~N��X��fތ>O�Y�&�ޗ��rRB �Ť�Z�i�Y5Ί�R��˕��$�H��W�vg޳~��K�}��C��0�]���D��d?\����ٟ�q;o�"����۫Ж`M��Q�����Ujab�s�ycOY����f:���%y�ι��vQd��.uY�~��p/�\W�z���
��!��0(Sm����u��2���22,�emv,��S3lo�-��x��頼�dF���V9\{W�Fp�O��$�$�z�(�&E��%m߫���]x��J��%���'����"�R��cy]n�*num��
rr[��}����b�Y�O)��wpi���qa�Z����{�n��V\����Id�������i�k��7A.����m��34pv��<�ٞ˗v{]	�y�Q�6s��m�:8���/Ll�	���kpm�6�N�����HN���\���g6��ý��z�hobv��IwYݻ��{u���]�NY���eq�u��/��E ��m�[Bm;p�&!�GNy�t�ț�ٞ�k���3nl�'<��Z��I��v�էt�W��xm�7y���;���t��S����|���+#s!��y�'�3�w���������$"(��}Dg;�T���V�Q�0���c���'o��ڇ�x�[�^Uּ�#�Yi���o���ט�Y��������ƱR}�.�hY�����n�ʁ�G���G��tȖ�g�4Y�W��_�UZ
LL@�0ryv9W���2y(E�t�B�G�ϑ����Բ�ҡ��-�|��.�{��eN�9�z)+�L�4��y�A7T_�~V�a�GA�0� t�́����k�m��'η�T*�\~/��ȣdZ#��AB�Ja2���CmQyPׂ<}���H)��4��W7���"�Umqˡ�b��Y�:>����^_�ar�M�X5�Y�A�Vr1���j�a���b���\2Ȣ��|}֜��̈́��8�6nb73d��X�r��令��{kG$��9e}O�>�S�Ʌ�,�ΘJ��Bd�T�g������NO�+T�"���N�X��b{Y�nЗ�m�]�$�����ڙq�:5�s���6!Ӆ���e,5~Q~���X�a��}^�����*��p@@����tbw�њ�"Y���
w"%��]U~;��jR/���G]>�X�'5��_Bߝ�{z�o}�,{��.��gQ%�S'����Y�=�M��I]��ʴ��B�e�(=�*�"+c�)t̗�LKw\�"T6��2M�y����������y(熫FT��C;ο��%�A5|ݭ#;w֬a;B2��B�/Pt��a��zPr�A�De��WDa��oc�z�Z��h2��j��}iJ]����>���Go3�gc
x��tivc����2�U��F	�K�|�o�����a@e��Wo$�{�	CTu@��I{��U%L�W���i\}�7�g�C;x=o�e�����[�`aG�K!��UT]ܳs71X�(��"�o4Śe�Gz��2N]mηs��=�������I�(��z�������7�?[V~�4��i�f�3O1C���|�!�Wl&��畞����M�uYކ����wךn�G���#LH��_/�L=s?3�"+>��J� �������M�mz����7��qp���Űs�a�b�=sm"�$=ㄦ̄B\�s�����6h�6P�if���!Ca@��E����fn䉃(�:��u���3t����)�WP��5�{��4*p��o��2dt!�>ȾR�mn9�W�b�ʶ{:emq�`�:���o?)���l#=4��.f�Jq�U�����[I���c��t�Q��'5iC~�<B'G_K��:�@�.X�97^�i�]���1������_EqA��*���M�*��qs"�����X^*-���I1Z�J٭�o��Wh��x��A�"�oC��6�����lt�9�<���؞���M�s�:�LA)���ŭ;M���~����*�]�2N���bL�`��x�ɶ�i�L�M��?3^��~��F���@��4��79z�3�N�������]�^��ߴ�鈌+����vQr��v��hY�4;��P�DY���>"9I8`a'���ԢN��vt������%E�L\�BK���e*�eF����}Zt_X����p��sw�3���Õ��d{e������|1�� �u�9�E�y�mݫw�T<�Ei7�jݷ�^�����ˁ�.ax]7��r]�~�>�~y�W��_o�M� U��uX����ҕ��f�ձQ�u���|�fM��롏���*w���iK��1g��!{w�qh��A�LI�<��u��3�CU{\o�J������1�4Hq�|m܉;k2�eP�P7B�03����X�k�M�����b�� =�d���w�]�^IO��e��/%�5e@m� ڄ]mk�C�!+����]�(�|�{tn/.������OfU*��a|�,��ޮ4,V(a߻Li{ٚ>|�����&��rE�졐-�����U6l�/4�m���?� *��W�#�����u�c���,��������9�r���;����%|��ҷc�ʺ̔�ꏘ���eؼ��4��\���ڋ5��u����{d�}�\N�&��lK�[w9u�Y��:�%޷4w'��t�Њ�9˾Sw��8��S�HP�[|�,�d�p���R�H�J�d�/��;��$f I�kާ�2�=Ucx�!t�����qP���[��S"@�͊�@��6r,x� C L$���N��d�W���h1|��X��n|���:oX�+nơȱn�����!��șV�,Y���fd�{�]Bn��$ڜ�z�U�}���L4�ξ�a� �c�_Qӱ�:㧼s2v��>���}[s7Ԫ����L2�)ѧ��E�r�J� ��N�pZ���
=۴t�xw�}�>Ɛ�(ɧ15�6Vv�����^�5�X�Ԏ5�kܫ=Ұ��'�z
4o���w���@;Ӷ}�f]7@F��r�dca�A�&Sn���}t��X��=�B����E�ծDm��m顦ߩ@ug\�9mɓ��V	�����0�/��B���O����t,�G�X`K�ݯo�#RC�6�NC��=a�]�����֥G~�QՓ{]G�i���E�p�G���3ו�@���_�X�Ϡ�{3l:����%�gm�V�͚0�����ۻ���ɖ�s%�^�lT����.����{g�E"|f'_�/g&.ԕ���|b�>TQR��7/P���C!3׎��CH4�ͻ��z���d^�I3+q�EMm�}ْ���!m�骒W�����O���CL����}.0>�:�1n��!�r���Yۡ�CE��9;2J���홒of5��U��ԣ��fE��mV�:���ʬ+zTnh���[��u�������Y{R+���S���{�iKu��q.� �A%Y�}g�fV�{t�:��xV�z%��b�'�o�����"�{���Wf<4ͯÚ]�?(��;�4�	٘\|Q�|r�+��\�-.�����+v���6��vn7�v�W;W
gT
�� �ȞO���Vi�];Ⱬ��g���Kc����/���J��m����G+ivg��x��1��K1�#����˓���"�d�VV��/v�+L�j޼�+{H��k��)e�L��*>�m.PK0��흘^�iv^)6GZhW��z�<bCW�6e5/�{��G^վ5�c�N�ZA��J�i-�5�(�(X�!m��Q��h�7r��@����JI�6t1@Ͳ���N�H�v�_�d���n� �2��A8 ]�����ٝ����y��ϙ�vKڢ�(Mw�0^�7&���5��	�W�ݞ�ɉ�:��V��{ÐI��ݣ���թ��79���)��F����A�]��цe����tT��no�>�i���W���nz��f��o-.tX/>�D��ˊ*�h\+���=�*՝��AF����o;k\�gN��1���f���U.=�����^m/�ͫN���E�ۙ*t3p �����ltu����b�����ūn�	)���v�vv]�8kY�8]vդ����h�c��w7D�܏Xn�u�g��''O���#ڹ�3��6��K;�r�؆�u�ǯIn�X�ŗ���]��6��v��z�{9;����.���{�XvQ�wN�<y�a�c���ϨXz���Lo$��	KR�mr&�nZ�;��)݃+d�ʛv#�-�rr�s�"v�����n94�9��G]�-�^-��p&�̈́�y�<h�ĸ�;����'6�N�\W9��H��:n����:W�nv���LH��%�*9��0�����F�wlnq�e��댈�Çf�=�����9�g����ڹ����;���+c��/K�l�a7�F	"wX_g���-�d�Ǭo,�n���v�z�p�kܖ������$�vbw<W�
�++/$�;��%�N��u�<7=��#�&�&&��\t�vA�s����:,m�k��1Z3�yM��*��M��ɝۺ�z��l��%�u�[���˳!v�s۷;�X�%�s��!�ku���c���q.��\�tt�BoE��1�nwU$��uF��m=gC��c^ۦY���`���<�nw;����0@�s���k�lpf�nu�c�)�P��l����u�+:;�&�F�F؆6v�8�t�xۮڽtl�p�Y޴�����mu��E��P9ѳ��]Qq\kљ�����ȝ���	���9�\��rnΞ��z�z �kv�����8�#���v��nˇ�ۻ �z�,�۱�F����6:�۞�x�4<����O�x��Gq5+���`��v�s����nݺ�*����-&0D�ݸ��$U��&{`uԓ�{��Ɔ�+�F1���1�����eO.��nۥ�2��yϧH�Kɢ7�u��K���Z�[ pf�ծ�x��S] j�7	Ŷ��[j-P;Bj�mry�QE�I=v3GGۮ�pv�cq%p�y������7e[Nm\nOb玶�3Lz1��P��
P����m���&�k˲�����h;n��xp=��k�xðhsi蹺-����^�NOC][��k��T�����;����j�kiZ73��!h��7'8��H�;�nh�fevn�2�n,џM��@iC�ps��3q��=�mvp��v�[n,uo`�;h��-�[��U��l�'������؝<w8��k��[h�X'�K�g\��>
�X�Q,�p
�[ߪ��Ј}vh",���"�UV��GC0�~�iC�!����Q�o3غ?�.�d�)�ZE�Omm�f:5�} �����C����<�00�p2ڒC�=~�^�#�����L]������~�P$#Ƴʲ�9W[R1��1_.�Ϩ5�g�aJDB���!�4�O�`�;1���+dE���-b+��IA�#�$�b�PV�Uگ�2����^S`'jW�1dmz��!�V�5J�jt:�;�[��1%���Q�a��5��ٍo&W�d�.��}����V9��,I#��L��=������U{�z#GQ~����,��{���F��3�z�;��\�_��x��Cj��O�A>[�@�[·��PB/�I�����Ж�I9#JCWv�����?\����u>n.#�a�Z6iƈ��&����[�-}�e�b���I̥t7���k�I��S��^C��p?R��2^���:*yۨ���m8FIKɍ-�#nB�#�6^*�F��X[F�7�$�묣g��d� ��v!V���I	���*�[)��dA����?)ة;�=w�L������^�%˙%x���[R��]e�M���w��x��N7�}̒�w���[v�ŕ����׷f��rb~�����;���\�rj8S�^w� ��aCyi�R(b�IX����x�Bv�Y�W�<Zu��ϛ�V��C+*�%K.<J���䧥T�ʈ��J?K���e1�ri����
�O�����#��+W�4��>����z����1�,�݌FJ�2Z<Zspk�,zMfEM�n=�^�Si6���Ɓ阢��п_����D�ؖ�
��l	шI����8\�O��-c䶾���w�U�dr(�4�~���r�ke�$�{�k^���ج�#�� C�m�~�jδv���%�6l]}�PHo�t�ū�i��V�J�����H�p��}~o�B!�=u(��y��ϡ_K����+'k�E�c��P��*I��v|,��}����oB��=S�Gi#���|ma���,1Ĉ0�bn^��N�Om���K`^���F��z���[ny2Q8�F�VK����h�)P$]{�J��|�t ���݊�����ժԯYo`4��e37ށu3``�^�p���R(��n���"��0��%�$��gKj]��?��{��t�׈�u�A���7�a���&��~�Q���������Hz��Ԯ�n���O3zl��3��^�>!�I$
�'Abӛ����;u�ϋkULi@��]����u��%x�gws��}�e�0��p��`��6�uf�J��=��C�V�g1	��1�ra��#xvL�^��5h�*M���$�;���Sx򷔮��R�h��6�S*���>'����]�~������H�cd�Xl�^y�[������n��3���zp^Xb�eFϼ��u�	S́qvp�(��>��6U����^J֊��g��v�/�l`2�T��A�i�(�tݪ:jWzJ����@��G6�;�.Y��Y;�-}�_2�1HuU�PQ�D�>>��H�dz�O�*�{|}�L׆���`�� �Q��5q��	yV\8R���s�N���|:X�Ʊ�U��L���!-�Zq��������J{;�	�e����Y�]���e+��k�Z�߽^��a���\H�������C�r��pV�1&�8�n
�������q}�ʾG��\��*�K���]Q���E��.�R��%X�v�Vp������c�nj��t' ʞ�z	;xe���T�v2��$���T��~��2�o�9�Hg��~9N�-��;��:g<�ݡ},��F��"�{�5ߴVeA�������M�{��{{b��_��b���ͽ�]��d���4Ĺ�o8�V+�U@aR��L^?BA��
��EMtG2�����ז�����U{1LGP�f���o^�we=�E�*	<�鬋,�
�O;oO܇=�;3"R�c��:Ӵs��tsav
[~6���9+�����[��q�';�4r�mc��ɮ?-�54D�"9��ϩ?v����qGT����9�}�yZ��}DB��"Uo*�2�g�C.�z5V~��q�:4�}@�Jg`NM��b�l��K��q�gz��C�%>-�Da�V�Yeل��G̼���;x�)�B��"Z�7�{ �x��q�I�~�[�hҝ�����7��de�3�ġd�>��qW���,�X)~��X��wܢ�2�#,N⾺���<�R�*M
!�b�8lȥ��P#qq��F�b��>�3�'o�a�[��+D@x�[�d��^�7������:7##TN�i9�<-HjvK5��X7�x�~TB��E�5��5g��t��{_�|�N�*#�*�a�}�� 5�~�� \[�G�O��h@��Т�D���W�95�k|A�wf�������U��/�Ѧ�Pwr�*"�/u�&�$��*;F�gor����V*�R]�)
e-���F��\f8k�7�{&�C�o�Bۭ�����-�!�D�ߥ;vx�Ւb�\��DH��ޙ��d�� vWd<��a�o�8UZ��;�f�r𼛼�_4�d��F��Z�=�=��X	b�,ea��"��L�������Nō奛̂46�������S|�-�j��Id��8<l=����n���>*���Pm2�u��Sżt����˷Bh�ܰks�7$��F�p�����s�۳p)a�x�\�Vx�Ŏ>��۱���7[ooF�'��9j�J��7pzW��֋#�� �g��l��8�;=�ŧj9@�Zy��v7Ŧ#x�ػ{i�9�1�n�^�x��8����v2�Z�6�j���>����<��1��u�,�ë�F��u�5���ڞgET�"b�2�fV궽��0�S#�qh�������i��g���CJ�̌!�Α���[9=���qݍ�VN1Ӻ�ǰe��l5����Y+�@�A�*9
����I�dUu��p��ڲ:X4�ў�|�Z������#�X~(�����]����Vx�:&{w����0��e+j.���@�)��28T���/%�T���7ǋ�׳�m��ʭ���J��ƤV��k'.>����B����m7�/��	�����e�ܷG��3>�}���>
����K)?s����uW`T�λ�˴8$o4m0����̈B���#�C+��9��.ɠ��P%����U��L�����O^�ܾ��?-�4�aCl+��޹����<C���t��T]!zh�9�a�Oҡ?j+�(wֻ݇,�I|ۢ�B; h5��B�<���U��R����:�����r��	�i1p���o7�{��o�[��S�0�RA~iw�q���<�)^k���X��χ�'�Q����w�0E	-�]����*;
��1�H~k�S���ҁ_�7���w=�� �h�����k��:0XVH�Cs�X�����ȺXr�RU�z�q�71_��YH��97���{���Xi0!�2<~���;�~�@�D,�d�z�;5e�0*Z����Sia���uwjaw�yw�C�u>��OJ3ҷ:����訜�5\�^2a��|�}�l}	5�6�S/����(CE_%���q�s&<x�L��y廒��h�� �1�h�lP�EL.���gm��lx�����Vuvx�gt����ׂ�
�}�>���+/�s�L{ɷ�1<�'lڱ5�]�C��4G��}F3$T3�EP�O���L�9Y� x��h�+-ax�t~�n�+`hR�L⏼%��Z���}��t�D��* W�F-�}�}j�E��4�L��D�.��.8^TD�yj��'��Ί<�A�a�j�mF�3U2I�޽ ��񚑴����{���҇?�Vs��'Ȍ0��D��n�~��w~�|��2�~����L�ehh�
�,`0�)Dc���g�"yD����mN�u��hn���G+3ڬ	x��eFl4+�yP��@H��ޔ\�"����dK�۸�f�2��ɋ&D�m���Z�9v�<���=st�ƳT���|���FMn1ѕ���1ZZ��v�J�s]�Ҿ�W�����M/����'�������{�S�m�51�����#�n1�ssIO+���Jvʉ`�]u����E�<==��Z��cM�6Db|�l��h��j�LO���>��Ʋ�=������B��a�r�Y:
8��U*7/��]�,���~f"�"�ۤpY�:����7=���#h�!�_;���8�*"�@`Jg^.6�aw��<0���Lp��z�O.���=��*�G�mحyJ�eR�s���Qh�E���̷t-���X8���~�#���[��Y��%��hK�w�4�f|�٪q���[���i.�խ��,��5��)ޥ��&[ �X��iG����(�ޤ�E���#ai��ݡ��G�����,���m���o�Gz�b��'F3�c�Un*:&��&����$A&�������8�\&:zr&	3F�/]��א#�ak�b�v8i�sz�9�+{bL��w�f��pY��KhOY�V�S붤hU \��l�y1���E;{X���'n�9����
oh3�wyR7�6��f�`��.�`���=g��*���� w	�!gʹ� �Ge"���1
(��O]vOtW��-�/e�g�ba����V��K?zvO���e�D/��t��P�e�m��I�S][�Qjd�a�G�eK2�s�yf�f��ѓ���}/_v�ifS���e�{Gk���eڶ/ƱN�V�x�i�s-<Ɖ�9-�
J� ���YUY��{1�{2�RU��y�kI���ɫPُ5}t�˺����\�YEG�w;��� ��������xoi�3�/ ��)����Ѷ�f�ù�5u����a��F�2�[��^}�F"b Dۇ�ʦ4~w��Y��20�	���6�*�v�m��Axv� �?=� ��t�X@�Ϩ�]ʝZ8Ex�1"_I�2�I��� ��y*+�=e��*��S��O�����r�c�۷�0���A;Ρp��A_m��3�s���F�
����[zr�@�`�Zp���$Hr#p�>�"�����~��f
E}e��1��r����y	�M�_��n�/GR���ˉ�R��;���0@�1��VNX3�;��eޥ�� ��~��}��T]q观2Umˬ�ſ�Uc�ϙ�X~�/�����^U�:V�0����,y���!�N?.��&�yw��-˒�'s��;���u�|�b�j=�P#[�7W
�ܮ��������:J��}ňS�s^x� ���
�G�F׃�v��qs�sm=d��V{��}�i��;"bŴ�m"�Fu�f�a��S�{1���vL��P�G[�\˛��랮�\ʎ�ˎ�X6��)I0Z��571��B�ڤ���w���m����K��g�<g�Fs����q���ƺ�r�k�9MI�:��!�;{�d�=�G= v�`ɮŗ�o2HD2֯B�ɘF�ͭ�竁��{8㬭��v ���Y:8`��Ż>ƤL� ��̆�<iᲾ��kmu���b�c��Nݔ^�g�=�����ng]K:���6M�T�lƕ=��]��뛗�� ������d���Qs�P��;kbz����gn��;W���UV��6׳-�;��s���9�uiQ�z�fV��VYA��#�>�`��[�������h��H���;��}��7�'5����mZ��H�K�w#�v��4o3�<�)S���}=�2�/M�;Q׊�=Ҩ�yȬ�*Vr�fd�M��b��8�Y�nu�pH~��u�����d����bB�28.2Z�a ��4���
�+��[���tͫ����i�L�>�a�6�P3�Q�С9��G
5�A˩^��Z�
`���Y�ÄO_���s�?]�-���XQ�������W+�暯�!i���
C��#c�PH�_�u�UCQ7m�>]6�/�{�R�;-�7�N������X�s�P��ѭ5���ם��I�ޣ�G�j
6CQW_{��p��d��������3�\���a����h6d$"�B�TBk9�����y�t�����0㗶�(�uߘ���
j����P���T9�����n�*v��{�Q"��;X���+K��w�kާ�`��3=�!��7VC!{a<�pN�&�u�	�� �Ҥ���t��W{��P��wK�gX�wD���O��qe�[��jaW��
�Q+���X�WM�p)
F�չ��� �vգ����|�e�����H9�����a��8g���z�)�C��E��05�n�8�F����s78��g�u�a`��B�'n��]�-��cAFI<��B�ޱHf$�{�T+}=�O�6�����E���]y[S�R�Lb��q'��j�iF�<pb����,��M��D=�����OzV�{�O&C���r�wu��n�t�U�/�#k]��#}�{�����b�AA�>e��p_x����7���:�1| L������,�囹�R@�G�J�������l��y�����ꛥ*��[Hk�[�	�P�4C_�"@����Ů�eZ��u�/\���d�K��n�n��d�"(ɒ7#��I����NjB�Ʉ@�̣1�)ݥ(���R����Y�:�<��r;�
Y=N�NI��w�G�����6�	�����c��8E�γ���v���"���VvT�<�B�m(��+�p��ӈ/S]&�9���Y���׽C�!1{�h�֙��"��ؤr�kLwqQ�?]<�'.Z
�SH��0���Y�ޏf\�E�T�2�x��q�f��A`���.w	�ª��ׅ�-��y��e6����M�)��-�o���Q7W2����..��g`���bW������4��hx���R�T�%��x2KNo��\�:&��5[�F^�3������wLi)��tr%0
��v�`��h��+o�R����T�g353ؖ�c<�2�o-'q�.�Z[�l�}�H�F�T���ð|��TT�p�F�vn����Y�/�Ѽ��o�5�8�i���مl
Pܳ�Ǽ�\��J�9{t0	3%m�?�m���7���ł⡼m\���6�V�
f�;�//��t?$7*+V���/W�\�=K0nUZ�iS�ٸ֌NJ�==�7�l��9��VT�=�)ռ�i1��n���@�A6�#8,�ۻ����1"��VS����QLGLv���a���C�d��s,]o��(���U��nh���]>FB<�mLg�%����Wq'�<��iU��}d��'��͚Џ����W�P��m}aڇ�^5��Q��2�5��f��ǭV���r�����WJ��:��٬4D*��hs���ý��R��;����yl�6��b��&G��_f�4��l�񛔲vGA�C���>�u�*��kl��ݭk{��9wg.{vr����r�f�c����+OZT��2�N��te����_� wC+;M�귈�q 2��r]����l�hN�4�ș:n8hp�w]ZSk���k�t=�XMj�r��N���[cn�X�8��t;�1GC3�6۪��� ��ΰ� 1�&$��T�����w�ι���E�<�_:�v�v3c	�O����]�=�-m(.N�w-���o,�|47}��c?s�׻�֠� B�  �ᱱ�p'|�o�� �|��3���{+&8�F	Xe_K̜yC��lm����f{�LW�{�l�cv�X�ɠd4ˍ��Y��{F��k��nՈ���jlq���� ��y���⌔$f6����;�pu��'�v��j����$�qOu�<}��Y����ݜP4��!��^d^s+���K~Z0��Ɏ��4$r7�'$�Z�^��.��U~5��/���t.e�hCN�����U�	�}Pر<7�B��EXU&�"���f}ˎ3CD��9�y�u�y����p�e�1����0�8t6��nd���=l�ta��ݑ���Q�o�����,��u���]t�^�uY3�邬��YweF�>��W(�q4r?���{�Bq4|/a޲Avz��ÍvHÕ�3;�7_V��:lz�r�̹�(�MK7S��T��������=ٙR��.�7C�ԖK̠i��MҮ尲+�����:�:�b;se����f������V苧|��#q��S7%:6M�ɖ�$ㆷvЮnJŦ��=��{k�A��o*r�т/;Ύ�ʖ���s7w��g�����rr�v0�{r	��D��9��4:�]��$�v���e�٭���&�v�;s��ø�|�.[�n^'�7	���>��B6ˊ)���~E��,��_����#uꌍ�ˠ,���5���Ϩ��Y�hxv�WOt�J����9���h���<�/��Ϯ��ns�#���0@�pߧ�ۦ��7��,�VQ�oA�oi���N8�0f��[�c`���Ia^�f����f�6q�c��Ǝ-�{^�+��L��i��K<X�����)�s�[�=��o�}����ufr��z8�1]:z��]���t*���l��.���l�w��Mx9{$8e�=�V�2W"��ii�����H��~�z+<]vu"lpl\���1�nAqw��y�`�L��Y��^Wt����w�	,Dہ��՗x���\N[����l2&�m�o��^*���K
���""������Q�u0'N���gH��k�.�7�� rz�;1�w���э�{���x:
ۻ�r<6݄Z;7ޏ%��\*������Yc�2��9r��/;6R+�H�A8��s�O3۳��num��g���[��6�0n8�����`������m@K���6�T0�^;"�ҧO1;��#�'F���Uc���;:ͷa+�i^��W�6ݥ�QX:F�^�G�l�+��uͫg�����x��S�Q��g��-�c��ypCf����[��;{c����8"9�'g��"��J�[[n���Ik��W�)��8ͮ�]x��h}�y��/�0�:������ېH8a��m�^c��=Ƿ;6�U��J:�*3�|n�������{aH�x����xvt��`$TC�;N�a�3^��ow$��҅�:��R�F���d��t�Q�Vz���4��l�<��{oE�fI��L�bBwv
�2��`���~��c#,_�~�.�~��U����S	눙l��rK�;#�u��	�mԵ�Q��2���=7
*�F�4�9�������c������x/g�6�����9^����kh�(�f��p�*	�1�H��>�-6Gc�����Y�'pƫu܂��"fJ�����W��� �>�l�iэ�Ξ�����f9�ۍ8��OW9[���s{j�T�B��|\v��֓�p����ɹ�fj#�i%�=)�x}����
��/�A�gAy�6��.޼71OT�v�G��N'��^�5`&Ϯ&�X�i8-�����[�s�+nv�}�v�Ri*�L��r�B̼����$o1��-�$�e%������X�Pp�x�Ѭѷu>�+z���#��X�Q�#���E�������V���&A����� �����h�[y����n�O �����W&X�]IK]ht�dw�}���[�쐹b����2L��wq�mI]wt��/��}uB���c�k
XnD:ST���y�V�g���]�?$ �{,I�J�}�.d�Q&��X%?14�2�M�����8�73Wc�T����e':�\��\���d�r=>�3<���gL����#u��
�Fn"�i�Ӑ�x�n��W���Rf�����Z���%�m?g*5�xB��t�6�ڍb��'Yڱ����^'��~���8��Luݵy�L��q�2�~�1����`�w��Z�F
���,{��;�2:3|m��%��V�ߓ~���A1�U.\���{����N�)�2#� )���Tsm�X�Ɔ���{4�5pZ�X����d���+��p�<C+v�7������n|PNdQ�q�iR6��Z�xJ;mykq�We�^�R�k�*V]�<DEގ�;h��go�u���Ƒ#����� 7FȬ��o���2��P���k�ځ/���0�t�x֟?$�-��A����Pެ�}��T�W�w�G���7u������=M2�K��P)9f�~^�yhN����Ϛ�\y4Z��Z�c�i�]{r֧�Z5�(�IƯl�������I����*�`����0&�<w$���M�8�m�ՍU�T�Ƭ������M4ue�[��n�� X2r�۵7���]��J�I����iǙ�=^�=�K��OB{�jU�B4��vt��d��LK{��aw4�����)ɵ�E�歪��~�QBȟ> �y2���$�DK�l�[��Y]k(�G�m�tC� �v�f�!q=h�6��a��V	����Jsr��p��]P�4 �/�	����9zs�[Tf4�v:)��in��+v�;oF}H"(BB-2d�uW_\��ݼ��nx��VK6
�n&�v��X(���ǝ/^�ܺh��P�H�"�Җ[|�2}c��Q}��QXO�,�������"�1�.Y�u�R��z��R�p��Ȋ��2�$�E����U��5��d�K*x�eO�>�׋������Gmc�2$�yK0���{6T"�
hL��cus���^���Xa[�2r�;g���W4<�Qy���>��>��آ��r�r�� .���X"���{�|SF����;l:L�R�c�_3�a��ʯ���Or��[�h_�G,6xlf0�)��J�3��pF�V���+1���l8oMpU��J۟L�k�e�F�|�l{�aӀVB7�O�o��yǓ�oO�� ����"��N���R��tڈ�S��p�<vȹ�Ƚ�1�%�5n([#TA��+�O`ԭ�6�^���;}��<k��e�u�e;H�/G\�V�m=7F�=���S��kv7nn^f(�%��s/O1-�2����my�}3��x��b�f�H���6"͝
�x����W*^���[���G����j��a1���I�\*�*��{��k�n�,�Z�=�CM��ez�6H۶�X];���':L���u�_v>~".ƍe�}I?�`$��R_�;CзF�ߵfk�x�m����/��κ��Ղ�}Nl���VJ��m�N��)����?=w����/,���)`� 6���A��J��ӝ|�{�$��`�Uf��8�B��+�A����7P�Q6Q��ԥME��|�,�����$ܬ�8�^L�M0�9F���J�X�W]����iTl��I{j*K{瞙7�����n5�%��1ÙX~��y;V�Ы�Y����'�!e�zS}�ΗeL:��#��*b�x����Rɻ����L}����fJ��J2G6���5a��;�%n�j��4�RL<��b�G,n�K��q�^KIwKevݴ&^�=�x6�۷��^t�-����mr.N�܇^�&$��jw��v�����n9=��]m��v�2��D%���}��L6�b#ks6�u;Ֆ����v�j��)v(������k:pwV��V<K�0t8��n��x�������T#��2F����n��E\�K����6��N.�9����un$lu��9ֲ���[Mӱۭ>r����%�جqB�+J���C�|�5��d����C��TR�{����pQ*q�S�����+��Z�7��Ȥ��5ݽ;�zR���x��$���	�#H�A���F}1�xSʧ��V)E���~�!�'���?O�"�,�Xs�ӯ��X=�Vwh�ι7����Y�9������yyn"�3����+R

(Re`�^WS�7,>��Nj�l��k���f[��w=����N�R.I�3�v:����,���j�8X�ۉFCL����];���>���	}z��~��y�5'2܁��(n�x"l�Q^�x�X��\N�<Tn�熹�Oa�V�u�C0�l�	0�����쭛|f-���W����{���\�@�^��ژౘM�~�IK�-T8�<��r�إ�^����윻{\��
m'!���nM�ָwM�㳣\^]n�\qyuTj�S�岪d�Cl��>v��P�7�&v]�o^�[>:A��" �6\6Ӗ��Af�r�zn�;��o}� �7��g{^��IUb�8�m��L�{<'�~0�[=٦���z�n3C*%P�[�{��4�ٍ�됉�M41�҇*�,{P�T0���Q�}�;�|���{�a���O�E]9'Z���H��N���"��f)��j@d��/3���*79��K�y1�S�z�!�}-3�.^�M2�}ca�lV�Ϳ�Ҹ��cL�)�Th� ������{Z
]�FmeYd��S�쵛嬦�S:�o32��)���L�UJ�H��M/y �c42�]��lo�1oz�I|��8Y�9D����#==d��Ǯ��Z}<WhX�-8
&n�d ��
2�r�C#�^l2�ʳg���^��v@~��{Ij�̈́����e+޼9����g�$���-��ֵ+ĸ�"c��p�Q��k�ƴN���lݜm�{�Y��)�"�S��ݺ������H!�������@�6��v�I{�JPAҡ�8Гڶ�����תM�TF5� [��s��L�4h���"Dlk;�wp�YkQ�<Փe� 0H}��H�����g�����O�����u��7i��d�J9<l٘�$����zs�{��=�qb�C���78�W���6����YMr6­�m��/#7~ ���9*M�Wҝ����W��C�<��<e�7��[����9�\�s�Cp���YOn>�c�}f3F:8!Λ�{�E�Їbb�
��(����fb�۝�H����w�܆u�M��N[}/=��1��O��jŘ}�˞i���r/��+�r,}C6o��jE��Q�P&��.���<����ŧ6B=�lܬc9��G1&�r��3��9���Q*R�&��)�o�����c�g������6��ݸ�5nZ��/=�T�ۓ��W%ۏ�9►�>v8ب�b�n�+h���
�p��Q�Sjz9�;}D���Ba:����	�.f�.�Km�J9S>�1Z<�.��D�l�*�u��S���d�!���kعwWU��ڬQ��*��[�����eu��-�B9�w�W���
@��M��[׸��!�ë����o��(����2�f6�M�;0�f�:�_�+�tވS����I�����{Ƃ��7�� F"�N5d���L͔,>��"6��'v1'4���sj��������{�{*����]�H�~)�7.��8c(g�٦�P�y.Oq��}ґ��z�;��+UE��[T|�����h7
՘�e������1�ٙ����7�}�V�9��WFn��aN���=��:�Z�s�n��B�P�AAo�ؽ��g��׫��S�f5K���j8;wv�nuھ��,��u8��$u�N����y^~�m��ѷ�J�P6�r�.@Y����jT����v�#�ݼ�6��0f�W[��u8����"X���;�=���H�#��Sק=ݜ��0g�W�/'O&mv`��iA⠙�q�yخ��V-���.+%jer��f"�R$=��T	2ۯ%����y?N���hޭ�kٳS�
ձ�4��]�e�N����Q@��k5�՞�2�SĞ*�$�1�'�<rA��&����n�q{�)��v<��./��`J���䎎U��Ȭ��^�ц�K��Y$�Db+-DE���E��x�-��>�d��V���K��՚�8ϻ� WQ�3t��*G7+%��Y�1�]o��ڭ���۠zjI&��1��pǷ��u{o!�I�1籛�m߈;B%a�o=���~��n�aQ�)٬~����	IH&<�N�Cb�r!Ą�����|v ;o2Z����T'f+�����T�A,�d�R�|+f�n�yW�ܢ�l���_��.Yю��O����x*��s3��>�t�ݐ�u�;,�d�7��V'0��ch�g�rF�����lZ���7ۀK�:��2G{rjDt�x�U�P�vc��L���S�v��!�}��x;o���H�m0�"/�a7��<�ع�prݎη\W_%[*٬�a����5.k��]$`����X�[KWUm�;���L�r�Ϊ%G.���Ql��������b������4�)��f\y��u�v�V"q �ᦸv�=����V4޴��f�;]��6k�Vx�Õ�v��Vꕀ�ۮ��'7��襖Λ�#��s5��f�	�0��Ƕ����$�(���|ԁ�̛ܝj���ʯ�NR턀�E�Cc@���vl�<��P9�f�f[��ɧ3evZ��W4fL�f�C�0L2�˹�,m�"�.�\��黴&��]�,'5�)j�Ƒ��k:�;w��z2��-�͊���	9Ç[��P_uu�l�v��Ρ�mV�FIG����/�w���ʹ���e�V��d��T��)ef���,��d�ӕ�m�g��]������*ӳ}�@zRg��֨j���@�ķ�b\���7���%e�f�������GA��P�p�Ӷ@����!�d�ԍ��f���F�66�n���zA���ga�nF��Y�9;��y�f�W�@X�GB��D=���jW 
yW����Gy]���ڷuƦ`{�?��v������ݱr`;`�ݳo��h6.���=)�g�{�X<�ˍ���+��J�����X�j��v:���w�]vݫ�F��e����z��a�'���Ƿ-���:�gN}���5յ�
���!m�or��<8v\�;\Gl�6ݝd�L���r��SsX�{v����6�#:on|��g�m;on}v6OE�A��4�l��Y[kqt�rCU��M��<�Ә֨ɞ�U.�<UlA��=nx�1�x{�l��9v!ې�ʞݲ�o�gw]g���h��x9�y�pm���t������;�[�<ռ㓧�&���.8��ce�bat䔗i-$�a��"�t�Nٺ=���9+�[��nug�7o6]��q���J���5�bԽ������t��^z]��I��X���OjGg+���1�ܼ�z�&��9|q��nێ����7N��r�g�"���q"��Խ���ٷDq���ms�=�j�)����|���9������cpq�J���cױ�ӻy⪷n%y�.��ܼt�m����Ԏ1A��g����m��՛�疎�ѵ�v7fSf�3��	�h��K����M1����;u�7o[�x�k��f����N8B|�8ղ��s[n��+�s�+�%��r�X��;vi���m7^�9�0��n�pnb��ݱvŅ\�7cglsΞwp;ź��vZ�@�c�l�Ʈq�F���elk�7�)�b�Q��.ݞ�$ϋU��;!Ɠ�]r�����<�������V8sȀ&bg�t��Fmڞn���&���n ��a�y�x$�^�$oE��;dF��y��:Q���>�(��Xz�tqS�6�w<�ڋX���7gV�l��9m��\�,Qn�ahݗ�e�o;��v�n8`�'��uyq�:涹3�n�a���r���s�&�up㵻s���VNx��m�k S�/>�Z��9�ۇ���X��۵���5{Y��ZWQdh��l�d������U���7<4����r����0[�7lg������n�ѻ��mζ��^�-�ō�p�n8��7:+mG=c��4�َY��p˦�ı��݄N��k8����4��:�ۮ�qۻ[<�Uǋ��C���8&2�ӄN���m[�(��sa�����t<�x�E�vωh��퇴n�zu�;</\���U�5tO^]�7�].�7r��=]mϷn�;�臱ϩ�6�R3�E�w���ᮩ;>����Ơ�ݶ������c�|��碚����{��N0Vu`��sƈ8�^ҷ�낗��I	N�=��l���b��m!3'�Y���G�v�2�@�%Z���ܞ���ѻ綬�_u:K%����KIg�[�oY�A[+4�f/g{����)�g���z�b����HI�Aqo����sB��+��X(�G�OKJ��V7j׻�5V��A�1;RdX�%y���և�1��ᣁ���"d*m�3�X�Q8ӭ�S�8�&�gD(���I1��;�\�L�� �LU�!�=�]�r��׋�^����gK�&�N�*4�4�$!����i^��	�{"��cC�j1�B�C�r�R[��ǻ�=�|˕�t���u�9�溷[H3�~�u�x��]�v�m�7vK\����1��$�
՝�Wg=�ËZ���'ɬ����ݭ�k��Qn�:��%H��e�R*s���Y4��ʡ�iGn�ꌘ��-��TV,g֔���Eʇs�0�� ϶�w-�[�&�ͥ�F��m��*�S&Y��l���u����4�YzNV����d�۫D�j-:e���s��
�F�ܮg@���|f��O	�+0�W��K�X�j����	��+u�v�Y�Ԣ}��J+����B�L�gp��P�ԑ��{��-W0)���}Ö�&:H��r��f���α�J��̪����U�v����K�K���p&�r3�6T������w�@߬�ry
N�k�9u�{���?v*�d�d���7C������旓�~��.5=�N�e��YGq�M����}�<g�Q8zP�U���
מ�U�����ޏ��yȧ�.�׍����N�{�f�1�׶U�5M*b@�e���d�{^����n��oc�m�M�^�n������V(H4�	X�?O��]�z_���q�]9R��hBU�ʡ;�˔^�Ҫ����p��C�$�6���E�$��8�*H
�M���䶾�������������o�'3�ӃاQ7�Y�/��adK�v��~7��=ڋ>�UK�X7�ތ���] M��(@܊��(�@���ƃ��3o�Po�;��3p�=x/n�t���ѵ-4��oqૌղ�+�g|�+�*^�l��m�/ՎO�gm�4q���t BmT����o���]t��Q����ws���׫ʅ[����ǃH]����eo�-�l�ۂ�&�{,�$��$�R�[���B-r��˫�YYەz/�;�3b�ð�y��h��.��a��2&`�Ɠ������}W���z��y@�L�
=��륫N�̄\���r�үKw]�뙄{�L�){U��7���֝c�EC�ZrP�nx�8F�ݵ�7���4v�v���9^�'h�D��TH&��Ē�j�@�ն���WZ����Q�U	�E3�+jzV*�_*���[O�&2��ԏ</\�	�݃s%��1��ͧL��ƺ�Z�����[Ä�Oe o��]co�C�V��e�U�S�`����]L_�޽��y�a�����PN˞]����z�l�2%s�������^zb�	n]3�o&�wp�e�K�#i� a�@c�z���2���)wg��y5�1C�A3��ȨC/����*��F_��F�.����[ͼ�#�+u`u"��Ӣ�ݝ�;^��q��U-��g�H��ˊ�]�{�-�f�ǡ��ۡc�ڽ~*΍k�r��gw5������t���WiJ�ٺ8��H���ur��7��]��D�y#��GxU��i���/ui�������D��)em�^-�**�u�>��y������$�r[ldn����������>59��\�7N�/(�U�;/R��z���7�Zv��92�j��<�ں�����u6�b�BB�*wU���x��J�������Q������A,*f�u���z��Q�����ݺ=*��5m��a��;��d�����q�6�D?��,�;����z��UU+,�Y�����2����;�{�j	����m{�����Y{�#U`�%���{�T���{�$���Â(�V�߮�/�}�s/��oMOi��n����c�t�Ԧ��Yf`C��B���{��5ɗ�i�ћ闳���i��ғ�^�p�G�"��N�-��]��]A�:���<=��ѣ��
����$�^ӯ��95"�����'�X<Iv�d܉v!�ڐ����dki캽�g�!���ֻ=���&�;�r��f��&ng���i"�_:�n�i+^��?_��{�on���R�ŏ��Wn���9������n�����o͋��m����ȅ���t�(�i��خ:�f�l�&�.�@�v�v�^���{k�z�*+��\����.ًA�\��-[n�6��ev�-�1)�;8{1�7�-��bn��ɇ�v�m��L�y������׭���6���q;�R�O+�����v(�-�J���E��"���z=�Q�er���8(�f��j��^F��[�1Q7���Duޅ^����+�(�M�^l/xˑ֯r��'�ly����^(������Y(����݋��L��Y��Y�D��Bd& �ݸ��z�*;wQ�O̦UZ���(��>�\�G��^v%�/LW�j��[[�Ȗ!Y����+u�\�b���k7��E�w�� ��D(��Z�	zʿdv�n�����1��4�����dTz���q��L�f5,BD)8�z>�W�v7�a�}��:w&��1f�[�/n�����OfY��Z^_9.�O?:�d�W|��!Q��R�~�X/\��k"�����;j�Op��j���1�eE�V.N{JůoM3�������#�|��xՄ�!Qi`�z��1mL.7l�����72$���vzΫ������Bs��v��8�	�q�N-������H�L�
V��-t���j^X�,�)W9�<�״TG�h���k�c�ll���ψgc�7' �p���Ȳ�FX�e*��;V�2���$�iA�4���>��j�ɻ^Xa�ZW!V��9���V᥶
z��?p6�����K.��)E_o(k�ph���V�R��ͤp��~oמ����y��ۣ���"P����"�He��J���^���������)ꣷ�%n��h��l��jw0�����z5w��=�)彾�q#�9D�//�M�o�b��9u�,�̎���4̀FXZΥ$N��ֲ+Q�y�fU7dw��.�	���j�,8��F�f`K*����}[R�5��#$R�3��;�;/0N����.�,�'�aos]�0�C,]�8���'�NoG<��2��[lK�2��o���)6r=]�6{k�x�s�x��-n׷�gZ7]0�r�O{�Ҹ�(՘��s�G�S<� ->�bl+����]ю6+��u8N>�(���zd��B犽0�|)��a��>&F�~�O�(<�`�,r�Ul^�`�׌�<[J�r��܍�Ѳf$aD����ԑS���=3��Nd�5��v��$�X��K�j,�V�g�#�h��+��X� ��}YF;$��o��=~e��" ݁�O��V!m�1Z]*wda�o��b�H��s~T�ʱ� >��]�7;���QTT�JW5��o�	��u �6߆�X��E����=�U���	�R;�D�c���X ��Ѧ��l���`�;Ǒ�%[��vyU9rL`�������b����q�o/;��n���/<p�W�,۞�Ȼ1����1V��(�Y�	��A\+�/or<���M����]GG]�n�t�۴x7F�q���{u��u�+;������5S`K$�J�g�@%p�\�IwԱ���b(9)Cae)��ø[)�����Χ�G�.����c�e�;�]���s���&P{z��=2�5����y{8�;�]i�y�)�s;V,'>7W��dt5���
���s�0��C6\dG1�:�Z��쾮��KacNA.��f���d�'��,S�Y��ѝN�w~��5�k�݉�"Y@! �z���z̩57������� �]ii�=�X�g�V.#ƣr�gU�2ԝ�>��1ѩv;)�����+�2|N�u�	�{�cl�ʊ�kv�X�U*�j
ӨE�Tx�FZ<뱼zs�7@W;�0Q��b��|��n���\7�	�w��Dh�oowv�Ƭ��Tn.hO#c��ĸN��3�u��X ���=�o�������-z� �p�Kx�Ν��c����u�("�M�gYpv�{t�*m�23��w�ƹ[��Xu���J"�)�u�b���}x30�ͩ+���ZÉ�U�j�҅�����ڿ;Ƕ�`N�$垙@Н�J����DĐ���7���S�t��3�1�� S����Y �	]���ј2g�0�u�̬�Wf���J�,�Mݨ��"ؐ���^%<��8{;v�iWR3�hC��]�Jݏmռ!��;1S��XJ����2��s�]�HF2�D��^A���|�=��<�sL[wN�Q�ZW q<5��
�p6����wg�g'��-�G�| ���ZN�`~��K�(a��ˋh�e�T�ƹ-�:[ܙy^���E���O_K�b����*��p��N�t�F{�7tqv
$�~�RM& ���pݻ΋��KJ)����sM]ca������$p��������F���9�����۽a�J�K�����N�ސ�v7b�v7lچ�1OL�T���幍��Og�۵���S�z-��'V<��"vu�޴^�㵛nܓ����q���bNį���|�Ё���z�o6m\�7n��#���][vN{G`0:��K���ބ��d�y��c{9�v�{2��\pݕ���sv��ev�m�y�ʶ��ᨍ�Q��)����$V�g�q�.[�ֳĜ֓�n�u�n��S�+J���Q}Oq�(e�<�o{&��9��z-E�~�Uݚ���xZ-d�\�<�9S%���B;Jx����=��w�����b�5�
m��"Ӂ)9Q��3����W�]u'�����e��EJ�,_:Q}���\ʌ+:i��-/:Fzv�cj����3q��Q��{�ck�|���`Cr!W��P�y}���.
-k.3��v*�پ8c�k��²��F4�}�*ٱ]���'�@���J��+1��u���kh4�s�c�v':7;o��G�iul*z�3i]?V�51�K�-e����Χ7[��t���!E�2�*�:���F=�v;>M�0�ǘ�r�ӵ9��ⰻ�`����*.?a廼�Mu{g�G6 �q��V�ѢWKi�%�;c�爛�Y�ػqn�n�6�f��{%��׸��f`��=Ks^Y�Rՙ�	��������"ȺY��*��JT�W��+"��kx�]�d�$�Q$'ZuN�"��{�sQ]wkq���N�t�wp���+IN���yI�"��C��Ol�6k�YG"ۛfi��.�V���)��
�fs��y����W�eSO!�X�v�6yb�[����Z ��8"�%���]�m�M�Q���
�ˡs��:���q�"\��A�}*�到�i��6��y��;��w���Ҟ����[Ĵ��Q"�P(d�#���u��ڗ���Tr�((��>�S	-�ҝc�SO����V.�ZCT[v��Q+3�j�8M�N�o#`����$�U1�[мx���jkf"��n5uμ!����<h$��@V:( �6�c�^�PSٞ���nR��γ�2D��Ɓ�#�v�om9��Wlz�v�7�k��D=��*:���rRY����Y�#Y����B!�uU{��^��W��E.�i���W�o9�u2>�h�ST�;f�Ņ��"�J}9�X�W�<�zi?>�ŝ�z-h��Z$VzL&s�]v?d�Y�b��x��)Y�n鏭81��s@�a�b���mT�5-��Č[�R��L+�L�oՊ+�=�V_-�Tv���m�S�#s+u�k���`Z��A^G�oW��1/�ʔڹYso�Ҋ7�j\�;��:����6gE5�wY�>�9�E�흕��/iE�S���]lԷ�Ut�����R}�{���S���-I9��ŉ��>G�t�ϼ̩�C+�U�cN!�<v;�k2�'j±`��qۮΑi���ч�d������lNK][5�1�Bwk(�ˊ�R�8�����SqMT�5IǢM�10KV��V%
(^�`�9��b�uj�o!����E�o���Նӫ�ەU������*}�ڊ;�CQ׉��Oz�Ս�Y~�kɧ�a��b�Z	�J�Z�.�ʬ����.X:��[��m�zSt"fK�~fEb7B�@E[�gq�uҴ�fk��JJ����7+]�=٨�11s}ܴd�����F!yX��?�l����lj:�9��>�}�x�_S�&��Wze���*Q,��������r�vҒٴ��Ͱ����Y���m��6N�e3��#Ȼ���+7]6�V+�#C022��?h�� �Kn1U��@�\7�6�f�۷���'��1r�&�[~
��R�籰�z��{tHU묬�L�%�����J}����m�hk���'d*�
�좯\���G�i��[ѼV�0<�5��z]a�|	��,
󑍆��N������\*x��1g�: }ʘ��$7l�^{���%)t�FM�t�ܚn.}��S�r����f%��ޒ}2��b�.�E����b�ͼ��X��3�ɇc��fz�ͳ�^';8�v%"��Q�̣*@S)�0fɮ\2�a��l;�-���ej��$U�y�s2��γ�,l�2$k���w<2Qw#��'�<��P�qO?X�WK\�P9��\W5�����_��:��*�N��G��,)��t%Ҽ�`Y�/�ZW�����f�!��I)BB)��Q�]��+`����#b]��3����&9���&z�a���b ���2V���=J���Kf-E�8yfq�m3Q�'�r�X[k�E۝<2ۊZ���U�Al�`��q��b��WN�1��c}�dǕ+`fPL�[*����)K��ˀ�l�wb��ҳƵf^��V��Z�1,�!�ϫjA���}��b6%����!�C��>�>���� U�ּ�����)qe9;sx`^)�����l��4
!�hUgtt��������蒶�z���G�&׷h������a/+�L��}�:��m9���n�,j��vV�n��ξ��y��f�nd�4P�{��v1�ެCsHZW�i����nVӆ�R�
W�h��\a�p� ^j�T�n�獼\��9x�3�em��VJ
���yqV{W_(i�Y2���2`˱غ�ѻ���x�E��AA�u�n�L[λ/Y�&�Z^}��'93��k���~�lL��-U�{��#�J���p�u\W���Q��z{h���?�Q�#\9U{/f�eߪ��h�7�~�����)I��ay�d徛��u�QЍ ��HF�dUwc,e�+K���X=�ԕ�dW�T�.�����,:�36-Ʉ�����i�rcǑuoVb�q�֡���~�`�xg��,�7�D�#�rc�^�U7�L�ᆀ� ��8����
&)qq�C2v�z{珓Yۙ�����'w��#^'�ΈVӵz�*�2�t�חw^�[�t(O���yD����>����	�'%���N�/��f��C/jnN����[N�-�{r�\u�����D3"�u���S�[�ش.�Lq��&�[{j��n�U�`ٜi�e�������_�:1Ywb�-�����P[��k�ȓG˷{�bɃxs��
�7-i��:���N1����۱�^N��f�����8�6y���[��v��P,!ƞ�:s�`c�w��B5����^R�񗭗{]W>6��� :�!��eT�.�/�l��"��w[R��l[`����s�,@�����p�ש̎��8�����C&vi݊ծ���x��`6#��moVۊ8(g���V�*��e�<\���ɱ���ke<zm����6��Ʃ�ܲ�+��O2���GM�ݴ0�*��Ä~Kw�웩у��Og��b���cwso^6l�S/�$=�+6�;����d��چ�<����L�rK�՘�b/��}�XU��R��<.�|�jjg����kZ�=�ݥ���Xۮ��[iرur��gz4TlH;-���_0���7w2����K²��ޘ��}c�X�6�kkF���Ҹ��n�e��t`H�j�q8��)��EV��:�F@�U�h{���4��9�G{���l�}�ύ��y}��l����p"��^IX��r��^U�8(��"Ɉ�N!�F�-���6C7�ٹѺ7DS'e�$�Ӷ{jj��;��[��F��צ�]�L��(�p41�DP0ȈQ���!�۝t&��ٮثM�H5�����)�g�N@����e����kW�Z���ŷi��+?yXơ�+��Ȯզzb�Z��4t�9��;w��S������2Rf�6��3�������kL��٧}�H	������D��;����{^��q1k���+�J;�VK[�M���#��2�zK��W	zGpZ�{�Z;*����X�v���H�O"p�wT��^)NjW.�xW�t��t�����m'�w�9,�E�cm	r&�r3��]nP���o��]T�S��ZD���T��ņ�n���c�� pBi�nг}+"٤�cJ��V*H��,�f�*3q�t����G����i߻�ۿd��37ڻ۠�vl�)p�e�+˂���\�As��JR=�q���P	1���a�a=���u8���Y�Zmj�]���in�U�\[c%e]�Z�z$�L��i��3�~��8���nVv:�ڹ����8lǎ98�G+u��cn��2�v��v喒;cH&5�i\2dM {���z(�B;CF����F��'�{�K��G[5�[�`F�]�z�ϋ�E,������s�;](�=��o�4�i41���!�R���ٳȤ�{�]�֩�A�/�ߗ%��h�4�nVt�^�+�ߑ�ߨ�/̕����k�M��0ȗa�q���T9L�u�-'XX��ܣ��ظ˄Cw�E83+�ү��<ql��R���ҡD��7Rù�\�H��^!��W�W��Ù=����#�y*�|����%�4��ռ��F����]�����N���f�8�h�{'hR#[X���8$��M�rj�z��z�*��Ep���Y�%���o��x���q�8n�x^�s�Z�|K�{x�=��r�:�ꬹj��Ԛ��WH�!Ϟ����iݷw%�[�,�����#���c}\lt�]]���F���'�N��|�K٬�mA#���썑u.��n��ڣ�n��?U�Er�[��E�g����J�\�tɷ�U��ލ�@�R$��̕��E��S9�y���4�+�mN��H�pL�Ո*2K�(��G\r�;r�w��'o7�3��-�"��=�v<�=��w#��fK�����Y�1y��7|��,�S�9�u����f��vx.Z���{��1ʠ��(��PIF�Q̛��a3:�:��	�P8�Z�掭�	��t탫3)�W*���;L'b��U�*�my~S�� ���!A/��Z'�u�\��p]Ɨ#v-�y78�^�ʍe�d�������Z>��̧��ģ�M���ڑ��l$��&Ñ�(Y�+;*����V�k4�
ߴ�s�*�;���Ӱ��Om��5MT3K��u��w�A4=�S/2Vf绮���K���*i��t��D$�)��]�퇑9�n��p�ũ�ؖݎ���Ev{�\-�.7V�(�U[s�:��9��/Cr�5�n�'-ش���+�g��;����mEQy*��C��=���+C�z�3�%�n<U�T&�x^P��}<�*�U������q~��C�p�(Ӿ�xv���jH�j�R9�ɟ*�;_n����������WZx<�6RBG�ۏ�N��͊1�t]�U�-�0��j��Ͳ�nD�
@AR?cݩL17�^�?w��z�`ǒU�M�4��LW�5f���	�߽���Ѩ��X��<Hp�DF��Τ���(j�'�����7��2���L�*<� ���~��,��D�~��Q�����;��kL��#%;]D]�l��i��b��N��Q�i���.XhZ�� ����W�MP�9���5l��0��
'/aIp.�i��c�0W�n�3��n�х^�s��x�'d�ݹ��	��q�i�#P�������\�j� �0:\j�\g�mE�θĆ3VݔW�ϳu���-�wV��1]q�OU�={5իrhp<�i��g����4c�\�.�m�۵�t�gT:Ѹc���{u�O5��;��;u�q���]m�;K�Śx9��p�磵��c��2�7Z%��u�2�v:�yT��8�`(E��6P}������,�\5Zz�%��
�+vmRn5 .-��"^xphu��{�<E���n�>N�(<��Aa�Q7!ٻ����or���ޡ�]\��O��d]FK�;�,d�/*~Х�QVy�tj�i���C^s��-�DԂ	C6��rk=���FeEHy�+�A+-�5/��C�]9�^�RÜ�m�����X� ���]w�.��HI"4�N]�{ެ4o9�ܹ�]�"�4J�������M�
����e���L\���e+I�m2�j<R�D
-�JH��ǐ�>�[����%���,`;�e�w�xT�4����[=	Z6�ݒ����1�<����neC,(���"Jn�O1v۱�umU��=Ҹ��	�X����g�(���5�"�1%=��2op���0��kt��U��K�í���WOQ\0[hj �ή���]|�'����f@\*7"��?&d�����.�9�z�Q&�Z�7����Q�8S�|\�C���暇��gc�)҃���Q���\����˧igm`͹��Ҫ@Pi���N���Q�d����s�Y�u�x��6�TU[��*�ǎ�$@V��y�3عt��w���݅]*w��������''VnM�o�{MT �mQ���יt^���J���B|2�k-M��!������o��67��w�J�oHo�.���A�AF� �g��͞�vqIJ�޼f�"J��X y��j�=�����J�c�٧���������*~�rM�Nf�9�Q��ɲ(��������n��2�o-%���cv�#y�W!�2v�/k�dڱ��w^����[����v�8�d�$�l̥
�ٶsTNa�R6L��,��
�J,�Ӟp�u�E	Gw�a�)�ST-�ed�2�J���6a�ˎ�M�ݧU�ַ�qzd���wPzr�MPǻ��Z*��::X�.�?wݻ��Jf_�zX7?�d$��&8�&I&cޣ*�=��]�<U:+}��U�e������'���ۜ�ذ`���w��j�,w6�oQ��d�r�wA�a��M"�Љ��Tv���p����GC�Ǻq]xX��WQ��v�2f��5�/:/��Vﳦg��+n�e�������
B`��#x#��6Gc�0��R�{s�x/��[g�=�4���ڗ�4�3>���̅��ѣ��u^���h*���ͼ�ӋsB���6Z��P�N�ڧ}�l�vR�-�y�Y���cEe��;3=؍6��\Y����jBZE�ϚM���cj�xy3rm˹��/o]�z��X�}�o��b��+�(*�<���G=�g��r^Li�hq�r��׻�K-�U�D`�;T2�3hv���b���u�M��ۜ��bJ�FY��e�}uSw�&>��r����BC��{&���Ň�/ҽ�2��&�o�2�'��-���S{�ur�X�X�z��ǤQ[|)��W1��S��<o�O��+:\d �<�7������Bq.׾�G�m��ؤ�E�fiD��� �T)��t�K����IF�FK}��\��̿i�è�O'��Hvߨ�3�.�zv�nt��a��]�ע�8r�pf�=ʥ�q��܀�;�}�vK��G�r;=�[KtJ|�o���J�ƳQJ��_Z��|���>�R�j.����D���
ij��)-s��}�*9��m���5�
��/c%;;w���׺�j�hԁtdޱe�?kN5\v�=���ktn�]��6��MW[���j*�Pq�oX3� �S��DR)��={�tm�b����Y8���o�:n$p����DY�V3PVq�/�g�C�e`�y;��*Bʂ$�N�Tݮ��B:��/n!��oJ�W�=Բ�6�&	�X�]k,c~�4?Ov��t�fx���qs⌎�*D�!�D�U��J{G�P=�eQ~"U�TZ�/P��mK;�Ԯ��$��p��a�e)lNKht��q8�<<�Yԇ]�`��7�w�
w���<&QY��#��wN��/�^8v�Kp#��G��;�ՙ�3|�J)��O)�0����鴟?d����)�^�X�6����x�ky�]^/-'7��L\[�mϾ٠1��F[xٲ�T�sƔv�U3n�zz�vf�D�x|��숁��)Dn�ù�&\���.�j�zH�kYƺ���1:Vsh��]��Ѷ�����@��D�(^�R�a�h���%olw�t�Iu8X�Jv�tP��G�Rv�Hǣ��}��ز5��=^H���oK�^�R�d�>v2�����d�~��6�L�J��!�iY�={��Q"u3h�a�=[�;�m4ũ��X[Y��y6�cR�F^�lb�+�X�b�ù3iOVX6���U���K]D�ޢ�nN7R����Q�3Vf7�Q���%��nx�}�X+z�~���Z߷�]xyr]������{�ו�@�d�N�X,�v�'[�ض%B���K��Յ���nuug�^�`z�f�����;�A�/ZO����������Q�B1V&�es��{W� 3R4����lY�7-��A�ٍ�Y*��ҷ;T-��83�i������%]��Z��tb��1�ԋz7��u�*=�D KԻq�n��y���)���ط�.bOw�I�0�XU.���k�CJ��$C#�q�{kb;7p4�v���6�AW٢b���A���ͬ�Y��|O]��͡q��9Ũ8/s]� y6,��#ULM;���b�F���s7�s����&��!�0��3�5�C�����ܱ�ɫז.i�N��b7�ض���S�Y5���� ��p˿Yw~7�J�;��C���y��u�k�m�|G��w�&Tjw�Px�B�!x�uP~��M��bLA7��sW�㚀E>��QT�(�eV���;��ا��y9Cq6�:��2}��b8M�i饻d�A���;�0�a���>�	��\�۹8�u�=���yz+Ց�3Oc�P��P�u��;q����F6x�3�N�a�:N6W�9�]�v3<�(�j�I����j}�@j�ؼ��m��G����1�x*�N��81 �������l{��瘎�NB�x���n � ph�ո뜑�Es�5���p+���G��^���5�Ë����qs#и��AO�Nu�/;�3Ţm�i{�Gjݖ<@��6�^��26�����=�[��9�v�u���:�S�!j��rv�=f�'0����3���!E]�g۷59�a
Fr��GMq���0��܇`�Yb����y�b}����?}�!�r6܎��4[��[[T���nת�v.κe��:ūnx�v�m۶Ú<���ԁ��ơ�;7[��9�i��@/<�;�Ű`4wۏ���FM��u�u��QSѲb��˖�ق�.Kc��5��u��\1�o�������*�鷍���i��� �X�h��'\�-]T�-��n��vx�t���Ӷ�A�2����e�q�_���7�h����8�9u�{=��z��#�,��#����s��<Ӳ`؂�슉h��p�i���*n{[�{MY��s��Wu�����^���M4n�n�K���>y�v!�^$���xٛ3u���z����-��u���7�׎x�ݭ�]��ۨOsܞ��7c����v�s8#z�f�A;q��ڧ҃�C�]c�m��n=�/p��[f�v�ۜ���n�\
Dl<<��֎l�s����n�-���qܸ��v����ֳ��ʱ���h����;J9��6n��۞����g��ug��Q�Z�\[����!ֹ����v[l��ye�pc3ȉ��c���l�0u�W`S]X��<�l》S���mvnM��ɛnN��8���b{F4��mH}�v�gs^Q�m��:�}� *�y�`�R���ϮD���u���{]�]#4���ٌ�T��C�������u��SY7]�v8�;#����[��\�l���v�r���g��'1�Ɏz�I��n:�!�FU۸�M��ۦ0�����M�u`�Z�闫�<�)�gH!v�e�8�4�]ۊۮ{]���y(�p���{<�.�J�׷��b��9-q����Wm����F�9{y�$Wuf'g^S�yN�ci���i����������S�*�0>~��,�6��-��>��J;y~��L�){�8�8^�Q�*�,p���|\ 
9Tיw,#cY���B����Id�٭��ܻ���ݖt�r��������`��f��^/��cHA-���wR.%�>���M���=��{���&������ǜ�y$�y��:�U�<+�ꦪp<R��r$���͵^�N!��Mxs��y�\��;��$�W����p��=�|�/�8��$f�Vѻ�\s,�0ѯ�Щ��llN�K(���{�qy�؉����h-Ât�s���[�}nK�n����K^N�*iyq�O9����b�&Ij���e�x��c��톯o<�Qs)'Hݹ7?�q'aTD�)X)��u�I��MP�׺�u�'}����#vݭۄ�S���5w��{�E���'��7w��S~���x��R4��(��8*�7�^��Tx=3ǲ#���v}��OpϞ���w�0~����x={��k��T�� �Pv�Sl��\��Y�N�z�Y8��sz��	ڼo*
<�X�m^ى���L��5���"�Q��bO���C 1s�Ծ<C��ٶ���ӬpM������ڷp��s(����Υ�m;y�m�grH�'�*�bI�Q�欜m���7��D0�	�m\�+���B�g�N�>j��٩q/=��N�ǐI���+��W6��5��T������X��
�|�&F䊯���QW��S�LX9�ˠ����X{��
r�BJ�x\�Vޞ*wmXDj�"k��V��||�(���vn'�����C�݇��>9۬q��d��Y\��J)����C0�{��=,�ݽ�"��rxBƼ��Y�5�&ߥ�[f=�'{F*������2*R�#F��EJ�:��%&k/o|�2��큱n�b�z4�f셝J�-1hۘv�S��W�����6jЉ�E�h�d]WO�^O�p#*	@=��묦��f�4v��Mj<�}��j52�r�Z�NN��N�/���\�]�W��G��6,�.�DpwowZs6�J��%%ʳ�k2!��ʞ�^�dmK}ag��[Z�+kx�t���r�C��Պ2�mw�J�(BiD�N3���j?G�
5��`����e ��B5钴�[�A���"��N���}� ���6��M[��!r�A��H�*(��](<��X�/{}Ϯ�Oo\��(���~����.Fk�{0�7s�y᳣ʜ����r�.�v۝���}�s�ѳ��_e.�}*緓�6�#p���y� �k��E͞8wY(�����k�o��t����;����t�@������'[�+b��3�S�gxy�d|�W<�PDR��L�� Y���L���}�$U8�F��k��@�u������1��dK��W��;h`�FKi��E�rر���*���u/N��W�n�`M����%7��m�ξ+[k4d�F75�M�6��;ѩ��E�H�
.k��N�nǺ.ܮŰ���$��S$��`1���|�U`�*��p-����rP�����5�廸��l+v�Q�G�mh|x�6���A%ݳKv�X'	��_]�<T]��!u҆���*�w�ݣ1{%��g���-��ى{}�^��ƛ�틂{C��y�ư(��3ne��3�~�\� �i�g�#Ei�{{l{�r�����$��c�����:�۱��=`&v�Oj�����kaގ&��6]Ǩ5���.�s�	���������SEm�/�9*�[������MfCl��Άaټ�}K����cݙ�Ƃ1B�m�AI�w
�eR�*]����jQDo�&�r��z��TvKDl����r'����u"J��Z�%��ՙU�z�vf�:X�ܰ+$�����-�n�GN��}���V3�Y�yhR[����	H�7�z�fof�y%�T���
���FTQ��W�1���=�ݦ�;��|"��k�w����fd�E3�N����h���׫h�*U��_6v��pfYP玫�!-D��A$���v�`5w�����o��� v'ƍ�C�5�=4�0�����O�'y�V�ǻ|I| ���� ����.��ڑv�,V��Y*��T�;�B�z��Պ֭5���r6�@�Zkc�f/ym{U�k���y��/d�9d��^\.�6b�ʜ�Ѭ	�j�ζv���2�r𕷫��m�h�k1l�j���� >����q�ٵ���f�iݸ�3݈�s�k�������׌u���qpMxuW���{+�w�l�����ƅ.6�m;����k��4��ع.n�5u�G�3��5��b,�y��5��J�c����z�2[���=�i�㮤�����R��tll<[.[ۆ�Nפ�n�(Z7;��tmr�p�+v�����m����A�9=	^�ǻ�eNӗ��� �+�PMxѷ����XB��mew�R���H�(�����%5�h]��q�뷣<��9�6Hx=�����o?�ׇЌ?r�Λ(;�R��s�w2�f���4)/{�0��;/V{tq�����h珪�^ͱد��tU�)d�]�I������f�2��F�B��#��ޯ��#/�������1��i2`)p)�KbU2�li
*�xD�\�oX��G�I^������^fnx.�� �|3a�O&�L�Tф��E��7z�B��c���{	1f SZupb���e�(�TD>�k�E�7�o��������@���9.;m9��u�z�v�]���F�L�k�2
�7WG�]\��v+������w����8s&�C7�M*1�w�q
a�(�]{�o�*��௕۞�tʱê�.��"
7#q�yN�ji���Vk,�zvy����&���B|<�FZ7��[O+�c�*��u��Ν�MC�Y=:��J��x�V�Ս��#z���!=X3�R�A����ۗ͋��M�k9��B������]��֮�bSЮ���3�G��Y>C�~b�Vр{�q�{3?�{{�YD���T)�������s�5)�Iv)G���O<�7�[6��Er��&D��	���U��;nw�XdmU��G�T�;�a坴v�9}�{kv���:t���f>�X�ӧ�8�o��'sϋ�Qаt���XcQ�}��u'E�ʪ�ʒ�d�C�6B����ӻ&-�ˍ���|�1pf�߶�����yh%}�ɝ\Q1�g��!g�^c'X��<���.w6:k�O'c�U�іF*r��H�(-9�}��s|��j��S��7z�7�t�����8-��������֥�]���hx#|�qH\�����2G��]S�x}���:�7%�J��]��Q�=���k���^�%��R^� ��\�6{sw4Ue�N�&�H2�"��
���cr�^��^^�F�t�)�Q���$Nf���gQnv�D3�$�4a%�\���
�A��#^ۛ�̽҉H�����X���xV`��9�]�UV�y
�s��w�����31٭-p�9y��oޝ��(�`R�{+�1�m�`M�Uv��M�r��*��q���50�ځ�l�q��H���Ƽ0+�ۮ�][�������;���R�n://�+����~�&�ʬx�l�q1�jC3�n4�0a(�H���@ߦ���-�į�I8�]��:+N��/���`"	!$A;oZ��Š���
��Gx�P�q�8�nݍ�q��%��$T�
�9���s!�c���H��Qn��e���w��Uu��o$�i��ͼ���z�X�����5 ,VQo7��ry�m�U뼛�in7������3��r9�=Ԏe[	�a�	�'�y�����ge����ۻ���Ϟ�I2����.��h�z+���$k< ԕ12�ݲZ��49S�R/r4�6j�j-�p�{
��-e#twZ5^��Tqh۽��p+��<ܛWN�0jY{�L�Ǫ�`�7�'���Ԟ�-��sw[���3CzA-��F���vL�Z&tt�]��h�q��f���C��Y*�|:�7u@z,��g��.R��%�_���k�_1e�@�&R*�/�b�%��������*���	��:.��J�{d�5����KF��]�V��~�ȌdʻT�^H�1�p�=[��/�[��Pc;A��NC��{���K��nE��l���3٫�5�KP>|{�ik��t�����v��8+�nөA���o���~X/�^����W��G.r�"\�������fy�S���;�g��Y��K4 5\�ZY�GK�}��N�]f�C�_�{D�`qHC���&����;�zЋ+]�n�'��P�Ml�}5PlY'a����ݘ�h�|��e�)��7®H����[�d-6��g��w�4�6�d����ݸq{,���dte�5I�|� ;}N���	)�rq�xȢ/*�{r
�쵕�I�.edl6d(0�m�j�|�۔�ԇ٩��Ԫ_.�O��s334I�N��)�9�l�U�J��x��Tr��vkd���Y�5�6r0P�X��*s-j埋{|�2���8,r�13��mOn	��ɳ��o}x��SH��Ĳ��Ż��X_�L�v}j�z���J7�g��e9�mǫst�g*y�1�a�Wdp6��q�ŝ�=~B||�Ɖ�Jf��ڻ(����[]kv���st�Ǣ���!8�OOVl��sհ�䗢j��������:m-���v���[�����v��m�����f�y�'q�dΔ���n;����q��(ѸN��c��9:����Kq�&,8��s��$l���z�pi툑C�6�utk\�=�U��)ߥO4Ix@�����o����=�&��ظ64V�赒/&5m�/�^;��\ӽ��7��d�xR�2BD�� ��|ȫ����+KO�qyf���bOu��/$;FV]�p�V$�u$ZW9�_(i�WZ��B��{�H&�R�F�X^��"����6�'�^��������mY=����w*�Jp&��(u|�o�C��<ޞL�87�
9^���y���sdr�o��v�@S��yҐ�K}��u�d�)�<wu�9]2������k{=7�5�q��e`!5ɞO��f�3�����Q�
O0�L	�s���,]vS�Q=���r�mUv��E�#�!�Oӕe�L�HG5�sU�.��le���=�����y�&vm[ƈs�͵J��V��P��+�=�i��H��IgS�G|+�E1�f�)��v����Wq���d0sNkHX�������(�$��έ���7�]i��5����:]�ٷU<���4��fba�b{��Mb9�^U��-R�1��KG>�)���^jƣ�������{�߸��^TlX^9}��{�*��l=��W`� ��N�5Ċ�U/=q�NiX�hO�"�$�d$@ ����Zd_T䡂1��4�V��k0�݇�tʁsуc��3��T�`���)�����v�λ%�6��XWpf8Z1H0�5b���MT/]W|O�=�[�J�o�ǝt~|��b*� �&�y+4�!���n&�]x%Y)9CL�˼����Y6Ye�U�z:��H�C	��*^�����q^)�L�����q�,�3���o��{��A
{�ݠYW��ZV���S���q��Sחv�fqy!��кZ�FM��GCu;�v^.w������$����m�/���)��uYr����+��Y,ÄgM5:�\���{�,�Y�y��I}�����;L���ՖWh�iBH��H.�C`��x�nŋ����l�ry_���+V�\.����-��.S��©�x�y<*u�I[�u"�3sS�ż�7����o���� Ԕ���	�B�V��a�iշi	|���\��m�������%��z�d�T.��(�����UC`ǽ@���ZO<���b`ޣ�6KKy�e,,]:�n���2�p9�8�,Ϸ�w"j�f�(�w.��G^�f���/{U\�ȝz���e�پg9��A��Ծ2�$ut���F����R�r�Z'f׶��
��[���ٔ���^[�ڠ��Ta(�x��X:m�B<�cvb�Z�P6^J��@�P��J�5*��H���]��<�ҏ!A��ٖ��50��x.��&�t����~�a�7/cˣX��;�lE�|�ޏG��p��d����:9>�J>m��:A�8���{��PCj?'��pe�y�h��P�y����-�HA�eܷ��f,�-rm<��[�,},��y.L��s��C6�y�u��8�Y��/�������}0�r ��\�3�z��Z��k��g��u�|N%�q�q�I����-tts�0q�]F�,�����G����F����Wp;�������z�h�jV��G��m^c�+C�us��[Ѧ˕y�s�yǢ6�e�oN�Qb���B�δL|^X
����aI�+oc�0�Deoc�\��M�����|tj�z%	��e;�(���g}�WӨ��n1t9�3:����o�2�LߎZ�El��AJ=� �b��5�-5v�,����oS
�V�v^�^��S����F�3��W����O&��sl)R�h:����2�h���pQNB3��I��:�95.��i`9RE��xVo6ѡR�b��f�Û�/�<6=�]^y�!��+)B��u�^aȺAa��ˁ'$
D�D��9��dр����2��y�X�o��(��i�y��o���ֱ��U�?o��ܓ��.�]'�*]���=j��Y5�/�ya���b�ȓa$f���hֱ�g1�o�tU��(�u���Z(�,ƖBb��)UB�xJW�󝥱B��_�����vG__�����g����������DTZ'R��jd�����'Kt�<K�࢛�x�Q��v�x��v�v������⢖a�7:^�$6%�K��,��xf�g��EKs/������}��/���}�eW�,GL��J��|�y
k����Z��5����X��\(�lN���3�/��y����S�p�?c���`(��y��2�v�O���ƶ�N����῝R����(H1#�7���y�3�/q���j񔦥�_[F�i�e����qԜ`���L�w�V����4�dγ�9��?;6��߯ �(�M���N/��^����C��?P_�XZ�_��f����f��Ex�m2AQm����sTm�r��q�b}������o��L,�/!	w���=���#U?~��L{��~��
���X����vy�u��J�o�(��/�1/��V�I�mS@��"�L���Y�Ͽf͍q"��t�[�5�p���4�����"ӑn̓W��Pƻ���ƩP+�<�w����!��ʎ�;-u����|�S,����ՙ�7�w�rqKײ����l�=ɫiw��9{���k��͵�T�����v�`�F]��Í'dW�}�{�Ev�{�����~�*����s�{�t��G�Xp�#�<ף33$_ِг����rDm��]�In|��9��{����^M���=��	���I#Z���?�C�zEq>�7��v��wF4�q�?)���s��?rr׳Z�n���L���cwe��m���v��O57�v�g�r]K\�&F^��=_.��"o�Ð"�E0��n+�k~���E�L�,,�J��E!�s�o�C�"A�m&���k���h���ή��4�u�7ڸ���.��!��;��D:��`�����;H#k���B�>R��}���Kl��s��q�ƙ�r+NI�\j<�v��{Wr���
��6<=Fg��]^�mÿp�}Q<4����:���wDƦ�q���=$`��~��SӨc�~q>��܃��>�׮���y|��c��g)�|�=j�	���՝�|�˹y�.G/&��_z;�܃J�s챤��o�k}7�i���3��=�Z�n]r����F�g�3�<R�����{T��E~��{	�҈�YZ��#>�,�y|����gAm�qـ���{N�'��E:C��4љ �=�;W�L�L��1�n��ѧ���� �N�~��	k���n�G�H��>���yV'�]'���~�M����J��c��μpG}��ٽ����|�鶠��$���aW�y�ߒh�~�j���E���D�}K��~wX��K2Ha.cx\�9�8��~��n��D��_�p����KH�~$����^1�_������߇��b� iEn�J�D�w)u����6q_By<D4u.#A<��-�G�ߴU��7��k�>x�pF��?iW�)�G�WW���\��N�n�#%�㣎�ް+�:Mt�9��})�O�-��Vm�v�����y+&��g�3:mw�nB���[ݙyle�h�m��p�fR�&U����n�� ��uu�*�s�sݐ�=��o/*��y�N��L�����59�˞_���ݾ�;�:���Q��m�s�����v�'ziۄ�=��@utlܫ�z�p\n������Hn�w4ۑ�<��/qd�<=���.�ܜ�q���tʡ��Ђ�'klU�{xH:'o�8�(�����<�����7`��d�c�ֺ��Q
�/=�s�N�s]���f�f�������x�'��H�w_��h5�q#X���߄��p㋢b�������n�Q2TVЩ!�����a��]����|�] �w,�N�^�T�5%ɩW���>�6�Ўi��և��,u8������w�e��"�/3fӏX���u�	��c��DĽ߽�3�V�~��O�#$��^"�M��[�{�u�w�F8#�f�GLW�}�΃C���]*9"���f�ۈ����n�o��~��G���ָ�����{�Ծ�p�D���<{��m2��������ܨ��ڙ+���Κ�R<�Џ~��?nkY���q��J1�Qo]���jMÈ�	���_��X�'�I�"H����5ٶ�߿s�\x�H�y?:E��{d䷍A�o�߯�����r�eˇ#O�|����? ,���tfq����p��v;ψ����H�0 �*c���<Y&������q'�Hxߕ-�8��~@]���~��0I-�-h�F��{�~�����»O(��~����J��ں�4��W�7*'�����d$̳&L��a�;:��y�i���M����\��������$t��Wgc~R
�Џ~{�Ϋ�=��]�{����6�;�b;��k�����]���Y�Ci
H�K�����74oL�5��s��?o��Y%;k߽����)~՗t�	kG���f2��e��[�4\یB��F�x�a��f��mr{m�C�R߉]��R{�/ܑ�g%A8�o(�j1����w]x����T��h��5"�O޿�4~�ϳJ��RH��Ig!��Ȟ����$��}�R쇭.���2�Iɦ�G���7�^��5��ʉ��^���6��9�k������f��u�����nu��|�w�WdʗR��~�G�u�B��
�6k�,*�9��M8EdiB�{��\6�}�e�]I�,�ej��[KC���Z4]7A���Kx,9����p@����?jUs�����?j��a�d�O�a��*h������q������:�mW��HD�����u،���ص��4�w}��d=�������s�������H�TJ�(�7��ml�iܟ(Dt�=�?��@3�<h�@��_!#�?e�Pg�k(�,��W�\���~��I�n7����x���z�Z�Aq!�Vx��~��D���3ݒ��2.в0�+,�^qF���)��>!%�!f�ͯ׻��v^x�t��s��=���I9����Ѷд�*o��:���r�����m���m�V��Ɉ��^�?~���������ZP��oMP+�v���$���ޗ��	>4C!(�i�S*�<��s��~b 6؋����6�q�u6�O�u������aܾ��?^���A�{;�⬿x�+���
�<�h���k��E�3��~���_s#��t�B��_?9�Q/�������0�G�g!d
>����i=(�ɻ�I�b�W�#Qb�I�o32�N 	���(ݎ����="��4�R��(J�8��^���������1i��{����VF�O!ʓ�$-��~2�:�4�	D���Y��ܴ�y�w���;z����v����~~�S5{��S����6���oW�����8Ѯ~'/��R��2��a�����Q���/1��`5����N������U���u�V�#��G��{�_�'�o���*�ge��mb��j����u\{��q6���~^L���!�P����(f�diO~��k�B���;��m"Af��8=\�ܗ���%��}دee�4K�B����{�k��������kt����X����s��|@c9�N��_�ۇ����"#�������?Ⰴ|g��i�v��<�	�:�\&T��Y�\lt���5Ά���q�A#O
5�,�
�Q���@~��������
�����Q�Q���iy��m���cwx�7���7������&�&/�'r����{�x�'�>s���wG^'Rd�/�����[��ɐ�{�*��lj~����,�,Ǟ�Q�����z�4M���[���3�ž�ie� ��V#_o����0ú��vm4ۋ��?OR����^�(���s~��(������Q���#g�KOH�]Zbno���]>�Wu�����Oz��m�19������P�]mǭ�3Wj�gomi5���kh��_�E1ƴ�#Z�����b�O��?2��0���wQ�����Qu�Ց�7��ct�g:��̙%K�̱��˴��x�q��2�}]�8|P=[�S߳V����:���i-�sMںϿo5F�����>T����??n����Dv�|}��g߿Y�8��FR��#^,���X*�kH���ʺ�Zi'&zt�O���_L�Z�]�&EV@äw�D��@a������?d�0�<C����n^{�?u���'�:��ɑ߫�U�$O�_U�0��2bD?R�H#7*�~#J�ܨ��W�P֨S��b��}^�X_x�ڲ7����L���[G�{��u3 �^o�������G���/��`a����/NF�rD�My����w���_�g6�#����)}��Ƅs�6,�j����{��q����ѽJ-��i:��������D�9��mf���:�������,�2���!Ƣb�]sUn�����sf���ge��׷iOΒj���	�Y��O��F.�_����kZ��C"ϵ
�0��:&ݺk�g���`4-���z��"<˓�h�-�)����HJ	V��E��7�jͣY9gPw��&�=|u�$�n�]���yƽ�G��-�&'�����;�G��]�4[\bv$Ӧ~��<��h�ibE���6�X8~�H#m|;m�!��vy�H�:�~T��W~��%w�~�8��)ףm{��V��:�?�i?6��V~�0�(א�|/�
����hW{����������#&p���Sj�ֳ6Ɔ�u�:�:� ��\��:�v-b^7��2�	���~O?����,�)�����w/���V��'�9���V[\O�{�u�=�{#���M˼v�!�����O�X��8A�\!7���G�&�n��ۗ��ô<M��1�G�X����|�@�A����8�'2�c�!��&�:�i����	�号�Y��|!�����@q����V��"Ȯ^�&/�D'M�5�� 2j��:k��\�5���#�_W�y��j�D
 q�BH�Xe���P�pW��h�,�f��� ��΂��诇jB4D?�g9
+�{���&<�_<�s�zu�3��Kfe���3�^��t��M��f�����ډ���M��'�&��Ƽ\1������#p�L5H$ZR��^��]��z��v�\i~���Yg��b��~�V�ԏ�CC�-5r�����=�n�M5��1榧G�ޙ�@W�ڃ7�a~���Q�G�~��v�o�u���@�ۢ�7�@�����xҏ���}wKY�_F��ߐ;m��$
"]��_a��<�� R�wˡ�r��`�fk��V��rq��b~�i���|(���~�+E����!z�x�OM������ۛ�܉֏�Q���O�D��ٝ�q:����u��i[{-\u3C9��^�jؚ��`�j�[=���$|V�w� ��t{�#s��PǼ��M�V��s�2]�����$̖K�-e�.��jH�]�ѐ6�v3��d����a�x�&��>�g/�Ӡ�n�����e�賺L9�i{ZfV6�:��u�F��}�(}U��db�mn�'P<1��ێ�,h��F��c��i�g��:z�I�#GN�6l�q�n���[z�7n��<s�v
�O@��\�J�z��Ӈ�9��\�]lm�Ռ�g��ȼ\Ǔsme�<dj�[=mے2fǎi��1q�C�n�v��7BT6^�v�)�]t� 1��L��?OBy�
��4i�ƹ�w�V�Y�z�~F��x���Q���D��!�Bd�����٠o<k��G�*��x�!�H־�,8~����5֣׷��T��jᚁ矸�P͘� ���q>Cڟ��B5��}?w�� iS������?����?@�_���u��q��F���hc���ע$�����?jW^O_7���7)Ck7�|"*���4��9�#O��><�.}N7��f��rj&8�$Is'߻�a��i�!�3�_��X����]93�~���1ʻ����,�]�zk�(r�Dl�"��w��|�x+�0��i$]N�~1}��amq�חC�2D�.@ӉH�Wd�
Q)o��K��#]��t<�E�7ߦ���<�䭴gY�1?5����?4���I����?�b�9HC"�ج�?aF�^-�o!�_z�l#����E����~T����h�oF�
ݶ3�Ԍ�2�h4�4�'�i��kJ����Ts��͵��/sڔ�L��~2��#���E��F5;�k!�?s����u��m}�oZ3y��G��X�Z���J���7��׿~K����ٯ�GvHq�X6R���#��d�Ds�{g�7��s��3�Y�k��%����6�/�׻(ƈ���?8��N�_�W���W��a�L"8��z�{�l	i~���g��?C�2=���@V�;����~�7�G�s[A��d_���߼hy3���5�R�M���O������6-��e̼5GZ�[;��|� ~���*�D���n'T��HF�����Q��r�Ϯ.�����n�du�<h�ZruZG�����lS(Պ�!��aEo{w9}Cur~�?���n��q�v^����W��Mm�{�mm4�����l-�q~������_8kl�q8�K;��wo>ܪ:B%b,Y�?>O���ւ�ʊ6�^�^g���%�&�m�k��g]]����U���M_Q�ں�_�c��_g�г���Oߐ'���wJ�)��7���=������(��2�D������4ci����p�i��͖�z�����ٴd
�r�ם����L�u�&�~���r���{��'T1W�>�
�x�F�/�u6�5��g��g2����ͽ`~���?iV� B� 3�`c�a����{���G���f����`Ɩ�R��Z�?}ٓ�BBf*1�d�Á!h�9�g�5F����m-7�hi�3;���ܯ���t��������_h�4~}�(
��~��1G��_#�k����E䮾CM�\�Ƈ���3ֿ���v�Tp��Cm˫�t���$/-�F
Ĵ�\�b�d^�`;	A�Ú�]���/��,��(���~]�ex�	�8֚-�Kx�!�w߳T_��=M;k��A����%
�F��i����H���ͤ�/[5��<m��n�̣��bx~�9q0�*\�r�&���1�?��!dY~��<�ᕌz�_<�o~�[��ן�"5����7G�\�}4b|��_�j��'��i�&;B�~�Һ�t�_9|ߥvc�~;|��4L�>���r[-d��w����Υ��xѷh[�����k݅��i���֓�د���?eQY��gCe�˯=O˭�m.,ߝN���:��d]�1��9pt��o{X{fP�V/^P�{h�E�m���I�~����m�3݂�$����܇�(���vi�{۟�Yo��!���M��������\�"[��~'����|(�g�_��v���M��z^�ύ�E�hy��15���Y��b������<N�g�0����ӷ��`m~l����:>4h�?���}e��8��3f�k�%|���;~CM�����2�ۅ���7G��n;k��N��8�Wr��Qm���|��w섵תe�٪3���kmwP�F<~����tXK�������w�G7��5�N��kW��G�l�֏n}�r�~,n�fJ��H���e��.��s��u���ʘ�q��
e��i��;�����w(ާ�]t���ׯ^�~i��g��Vէ>�Ѥ��w��ᮦ�[�қk�B�,�=��[�~�������x�?s�]bq�5�rhSN��8ϐ�J��Nϖܚ�v�P��J���� �8G�(�c$����^a� a��V~��"��XU�a�C�̏־����n��z��٭��i�&}����u��7+������;��j�rQ�p}9��9xd��:�k���m��)>29d˻�yx�>~k���N�5��r��{n��gVE��#O�~�!~���_
�?�6E�_,����~���d3f���6d<����ro�Dk�y���j�h���p�v��d����9G#D{����]W�fȄi����Pe�����i�X���_^�59O<ԭ>cE�����@H�y|(�����}�n��Ѻ��g�k:�ۊM���;�q��Z ��&&��^��5���W�	ǹ�&l�D���&^v�;�2Gy�9Oz�Z���:舼h����h紎��r�Lff.[y�a��.�O��ԈbD��w��Zk�d>�]�g~<X��_���N� 	��3����*�
yx��l�P@����������.֓�Ư�u��\�����֩ޝ�.�;X�3���]Wk/+�!��A6=W۷��\�2k|:F�HJ��ZJ��_�ȍO�?� B{���da���n�d�0�j�G�����l��T�;�,I|�>��:���x��� 0�Ə���:�Y�n�|,��3f��_�!m�؊Fi�S�>?~�!���nv�����okE�Ӊ��PK�_B���V:����+��5����o{�Qƈ���@�H�33�,i��rF�{�r�hJ���['�4B��"A�&�	v�㗅�3��:�4Z'�s|t|�S�՞cF�正Y�n���F&����͟��K�Fj��s�P׍�(�@n�s&߷+�ٓ���K�ƣ�o��l��0Iu������q�x���� �}���-�^DQ��oc����}��|%�pk��>�͐>q�&4k&���形���Τ x1�j�J����4M{�t\���^|�ܼ����B;��}t�Θ�K�N,���C͹sMi�M�>�_sTm;%[�"L�n"���G��@Q�|.���7��p�Hֵ��'�}�%�XD���V��3R��PUW��EU����
����������PQUVUW�
�*��� QEU�(
(���UW���(����UW�j�(����PUW�@QEU@�(���U@QU_��*��U QEU��
(���TEU���(����PQU\
�*��1AY&SY��sJ �_�pP��  � 7'�`a� �Z�3�����{��gN�n�����zU�����̃N���N�:hz�]:
$�[����st��S����q���%�����    P�oa* t� ��G���w&�Kam��ml"I5�յQTdkld*���d֤���ۊk=՟K  ��/j�� 4 ��#{��o$��w���y���.�U��m>כ�wV�z{�u%�{;ݯh��2���ͷv��w�]7�m����te��)����(�D� �ٵy3� <��          R�    : ѥ�@��"��vk���[ P���(��={{ w�ؠPs����P4S����   � r�g�� ���^h

;�� ��r��/�y��]�� ld=��h�6� ��9g������ކ�=��O�����:���Һ���Y���woZ�Ҝ�;�4맽�w����Ssg=����zv��m��� �.�8  ���s�h�ζ�,��yy���z�5�{��{oRU;7��۳������k��� ��t���JAX��AN�ӛ=4��ƍ DU^�:s>��m�)���zze��=8�g��o&�9�E��[���P�� w�������wk/oo^�Uڴ��Um͘z��y��M�:�� z�� �N��7^��w)���A�]
6�S��f�7UV���!��L�w��:�ϻ�i�%^A�ug��<�{�9 =�x�@6��p���+�����C�!�[JR�i:��O6v������M�^�xt	�;ܸ���^�u����/]��)]��p�
��� ��=� �>�osξ� M+����g/C�=���t���x۹����{7h<�^���ON���x;���açV��=��^Aҹ�.�K���mJ�Xv�� �m�(
��]�#�L���w{�XS��c��OO;ކ�����6wg����J����9�}�^��]9h��ѕF������\y������l;�筠<�;+)ˠ,rtw^�{�Z����;�w3I.�ltgt�Z����:�� ����	�2`@�{FRU@   j���� �  ��H$��L�� @�~�*�    i�!)Dɥ4�M=O����?�����φY���'i�4��踩�hp�Y# "�
j4�w�*�@��\"�
�(
���p�G��B�W��P�UXUB�Uڪ�
����
��Q�TUU��
�(
��EB����UU����?�����u��E�d�g����%��6n�_�3�u�����0���G1	���E քѕ�^1�9E��`d����B�¸q1��:�S6�^��0^�{���k��/ ��]n&���X)�N�����N\���ӛ �O�oC7dB.m[e���Y��E]�h�2;��I�6�-l� �g���B�C�*�?6���܂e���r�0kY�)N�c��ۖ�ΖuB�rH�8֛)�Uɺ5x�(V��S1n��f	�������r�ٙc�FNx�V�������q�1�oSA9aӒ.��<�7���N�b�����L�J�wY��d>�pA���{"�iX;�c`�Ze��'AG�7��Q�[To.��馱�-^�J1�u�s�����1�rWZ��(�4�@��1P�@��2%�=j{�D��M*W�6�k�o^���B�m􂯬1|��]Gna��$k�E��N��aӿ�w1��ΐ���c��r���2u��1a$�=R]`��Kq�.���.m��S@��������ƳpԻ�LZc��X��5/va��M_T�}���1V}�-Y5J.�I�a*��Z}8��9���
 7�5��d�uz�"�fa�`�̄�ډ��D�.;�ͳ�};�����Zo�ͨ�WM܍G�ؕ}�����o�U3��raz��&X��w�8h�>!����:X���Y[ha91��fy�Dy�����ά��e�\J�d��+�Cb�ܓk.`� �<���
νn�R�Ӥn�S������.���Z� ��	B"V	I

��`Ԯ��)�ܲ�`��CJڸ97"6�r���e,�r�S��R�+.^"�Z6F�;woUkv@Ll &�b�ՊB���ʄ�tYP�A�'�wT�KW�nf+r��:�$�v���}6ҹ-c͛��Q�E���A��9�X�0��>���LG(�� �[K#]3
�91<Ҧ�`lц�J�ff�E���M�jJ�ӳ�eb�J+���Yt���H�{+PD������(��]e�7��r`�v�F^��t�}�]i�{l
[2+x��/�� �:tBԷwg�I�Ӧ_	�~Me�����Z��,Ԭb���J�#6u.���Wv3RJV4P��J4�)tІ"n5$�q��Z�D��!Ia(r�:2Gŭ7��HL�y�ˢ��L���k$��]�/.�X�(�r�	�[��â�ӔR�ߋi]Y�,!^��KU�KX˽Y��$ktܑb�զ�'��րUsN�k0\�)��"	��[�����kK�F���+.��KÆ���]�u(܏�+�O�%�Fܹ�n&�r��p��۵�C��������e���^�t�r�8�=��{�d:�8.�����(�u���Y"��p����im; ��@ZE�Y���G�P�������V0�N�/fZd�.���4�o�D�ݭ�J"�^]Ò����Mn��QZ�
���˺��V��azlT�"z�E+NCY��i4l됬��ɒF��m
.��21�.���xͼ����Y��2Ao��w9������|9cɰ�JW�t��wL��,!�KM��3I�<Aʗ�ܘ����E�V��͙�VsE{��{����^]�88������M��x��m^��^�x����tC[�)���%�H���0,Ia��֬wk4�ע�1����V�x�����dd2H� w�D��q�=ԚE�*�R�o�%Z���i��&�(���yL�ݫzѼY��3�iY��4)`1�U�jŬ�#hjr�".ùIEP�.�#hP�;)�.fަ��zf\۵��,[y��ܷ.��V�7�����v��X�c*Dn{4Ԭp�Ў��{g>�y-��+`�e��B��F��aX����i�2�9F�|�X��c�9iݕ*�B�ě��+ Enݬ�Q�J��[#y��ڜc�D�ۛ���9�����(Zb�-�Q����TT�4e;xv"��*�-�w��vu���I�q�.�0'Ȳ�3d�V"�&��?�
#A
��(�����];S�70�� ��XZ��q�c�yw3.�뢇P6��eiua��t��:Q����WE�w^�N��g�� �P��,���UUo]3\�X�W݋$v˗3��:l]EEٵ����l<�Ps�t��:��\����}��8>���qy�EW��ш<^��9v+��qA2r$��U��T$Z�ѣ��Z�+۔�Y��tV�����β��ok]���V��i�t6�')5�Tk�ib� `F2�;����\3���N�o0]�l�8�[f�ͬI����`���<��Tm
��P���%n3�v�͎�:SlW��p�,�a ѺM�A�jf�[�D�\���*5��om"/�/Vn�܂�Q<�����8A�\E
�Ý���j�f�[Һl�������%q�=��j%�9�reX��nȏ�Y��m��\D�4����6���ɳjڔe�k,U�r�K�孰��#�9q�y������]��\�;|"�x�O*�om�d�z�M��b��g*N��!�Yx�Y��ɂ�����`��ΆZ4��!Uj��X��FG�S7J(�p�h#��6f��K73�8�čؼL�Y�ō���p�����%N�c�%��;`�弭�/^IST�ûz�2f����&2;�C3T����h�#��cf)0�&(�!ysp�v/ki ��iHM\�^�7u:st���f?���ݓ�εQd����L�
�G�$�5Ayi���BL���zM�}�/��u�W�dZ�G�۲r�xQZ1��f'H�7{��R"b�j;���˨��ˬ
Z2�CQ� ��ʉ-��ҹ�M�n�nNL<\��ʂ��8����p��8�����.ŚdnL5Č�.̭&��b:uݝbaݓ'vZ4��h!�%�HCG^�ц�`.�ݩ2kl傐9�L�����,�8\�۔��h�5.<ATw��e�V-C�L;ùn�b�L1�r�G [̣��ݩy���Q!b��iB�3F�����
���+��W]�k��E�ŷ��ih�rw�Z9m�h9�����[ZsM3�5f�cn�B��y U�/��"�Ƌ �����"�U����L����WK-�1�-�͖\ͻ��d��C�氘���Ȳ��͸�*l����r�}x���[`AG	�M�b�X62�v�&�8��"]]�6�ȡ��Z��f��Nq���S)�FI���myk���c@5�	q:�Ѻ��2h����J��)���;�y+SLY�rȲ�^�F�
�b�7����x���nh���\U�.�3��S �Z9����li^�8om�/���cx�j̛nuAC�5���Y4T��L^�k�")�����)͹pY}�Dٶ������`7V��)�l��n�eu2�[��'[z�����$2���J���{5���Zm]�K%�4��QZ��N.�ʝ|v���:̥����}D��[+i�� ���I��x��Ŧ�J@�ޱ��nf��J�h�m���ԡ�-���vm�]�]Ȩ\����^cB%��#�J�!�v�J�����>-��"��^��m9VލPR�O�X�<�.b���*����;���V	Z`{n�5��`���h��K���!��*��oj�c�iPʴ�޻�Y�ڴw詈�f��귳�r��^{<�
@�Z�2ś7�=�jd����r���8��"ƞ�kkN��K��X�e�x)޻���ܬ�ƒB��~���g�>�Z$�t��H�Ѱ^�ʴ(㫽un)_L�)k�o�yʆ�<7	�/,f�=p�/�����V�edoI�v�kF���x�ܾ���o��P�5��:�]h�B.����h��6&Pv[��{�Z锎-�9r��o���`9��R���j���a>�f���*�F����PE
�@#@P�*�f��H�@�TMA�
�:h
E
4(B���"���T�ut�8EP
�����9�L@nv6�-\�T?ZT����He�=�hʦh4l�ޘG�!y4$�Y1�a�&첚�;C��ge�U<�G���cy� ���W#�����l�H��	3��i�R��.Êڋvh�U1Mr�K�+N>^͸U�Yh-����iט�y��H-�f�Xc�ѻ�R3RN�4V��Z.�`�̢)�0ѫ�����nʆef�
ͷ*[��i ��
j���[u�(�T�f�uq���TU�!{�^��b�b�F�`�5ML����j"ͩc�C,Pvi�@W���aZ����{���9�M&Jyc5Ewk���Ы�N���)X�ݼ�r\r�!2���imӃ%���W��e�80C�A2؜:��|���m&vF�_�^�I�9ӌ��P�����-sC��yB�ԡ��Q�Wr�G��U��O�j�[�3)nYf�pЖ�۰�,N'�]�hAЇ��{e�"�u�5��yNu���E����qUǀ�QZs��W��N�.��c㪋�yi���e�[�H����82�^%5 �qP�h��Nf�b��|8i�p�*�`���A��4�zA�Dl��*WF����l:��$E����;�"�����)1U׌/����H��é���{S+��鉨�JVh!u�����0��hHF�V�V���6ivEP�*U%�ɻ�g,ŕ �FI�*Uk��fäQЌW��()���!�6���8�P2R�8��7�r��6�neKx�7b����lܼS6�e`g	��2mMǼ�Ή-�h]+��f۹(\f^Y�&��EN�Ue�)]Y�Mv�7S&i������Ʈ2�G©&�d��� w����o#��xF6��(��)0��.]�������<��+޻*oW(�Y�T��:7Xd��"���!�h32�wb�iE帛�c��1�Oc�(�-�-��hܙ�m���*Kn��^5R����å+�M�uJ�dH��ߝÍO5*���܊�ɹa��E�~d�@q!�#zM�Y�QB�K0}�*�M�J�L�utS0[8����l�gC#'��ˏ>�t,�x�,��w9��=��ŷ�*�$���aW"付��sDv»yĂ-iESK
ӻ��P&�:n��a��ڻ�h��(5�ͼ͙	�'vï+�d2+��o0ԴP�KL�e�&�3�s���,Ú�< `x,@�T��sU������Q�;�W���
Ų�tiL�#6ԖrP̙���ç��gV��St��Ze�wm�h�B�qѫ��,�D6q�k)7wR��V����+DL�;�.�X�LҦ]J�w�<�ʧ�9U��i��iS�ܜ�<�95��9�o���D�< �
4�(�@� DbD�I�
6�0)VB�6
8`"���	n���X �D�"���7J�SzA�PBY�2�m�x��/5I��+Ad�ɮ�i����jfY܃�m��{V�YM��d1{��	�J՚|9��˰S�7�M��X�!�e�rn���^k3xd��pb��v��0Ta:�>��ٝ��E|�30_�Z�V�sfQ՛��R#��:�LƄCtՋ�o�v�npd浼s9��Q|ˠ�\�o
��ha�|�!zP7�� @2�@%d���jA`¡0��0���.A��(����P|�(�8Ռ|���6X����zC�03:�iz�ڽXk�F��\ ^$��JpR M(OUܯnrXN9D� �EA ��N�.�� �n��۫����ĝ9�ı��ZT w�U'��i<�6�i:��P�B݃j=�s
!*]�ڎ�c��"�7{�I��Ѝ<ܯ����q�T������`�l�.d�ҫ�0�hD�n��7#ǻ�h�]�:Li=̴Ժ�J5�*�h�s%C����e���k ��p�:d��đʕ`݉`���`�'z�7�	�J�iE㫖J��-��;��x��/��m���x�һ���4T�8Z���ݹNGJ�LM'���L݂奀�,��f\�nB��G��Y�B�p^ �MM[�9H�zًv\���`f*��3�cCCfUޙ����4�n@�k��WׯeG1^��55
́�F�Kn�U���6��AŜ���-U���d71�69�;g,��m�nDsp]m���v����N�m��ڗ�nK�n���.4��[�+5�5�M�f:#v*ӡn)"1"�m��1[��J���+aɗ"ۦ4���4�%`������7�ڜ��.�l�\yA1�k��#f�;���,���Ed��;��m�o`\a�j���r�L�5]oi���g��E�1	W���qZ���VK.�NYT�>V�ƽo]�k6�!0�_F�]1+�ݼ����V[�Aua�*Cj��\����u���:T�L�W����z�!�+ͼ�]懀�݂��k�/�VFF=�����F�)#Ț���CF�Yʎl�z��%�.�0�Z����vzl�ך)���.�#}�%�Ǧ�#�eDm�dP�[h  VA�)$$�@V� �d �G ��p��	 �����@�(��$$�dnR9[h�%�8�h	D��PH
;d��(F 4� ت%uY �rm� � ���ݶ� tȩ,�Wi+U٩QKm�q��A0(                                                                                                     ���                               �0                                                                                                                      
ʊ��Y`P,�a	cb$I,z�v~���fbk
���>�(�)�jf-��tG1�d���7�e��R,���k2�B���ib�Ud}��m�Uw`\���W�X��(��޹Y.�(�R�]v�ޥ� *Ť7�mo;s��xDܤglFl;�f�%+��r�QI]��V�L�Va�\��.�,^��T��0Y�/m[�7"�yG�"߳9_HiT'<�{oGj��u��Ħ`�F�, \C\�*h�b�9�(��ا9zw':�����󞢗]��M��w}�q�uh�'�o�w�0����WW{�6�e_b����"�w���el�h�9�nQ��vzt��-�%4s�@�>��w�b�+.���^M�AS1��U�d�op6�[��ji3�7wSm��ŮvI��0�]m��V.�f�\Bo1b7��r���w/ �z�0�6�kYp������8�	y���D�cp��f���h%��v�5vՆ����B쭭ܾ�V�\�3����
us]�t�������̦a�l��=\gNѺ��e]�w7�Oumr�_,�^e��n�iVul�k5�r+�P���-��a�J�p0W����E8�I�|rv�1(�^�G"���x�@�]��ܹIM���U�η�긐�mu7�:^V�K�����\N�ĉ��'�^�A{�7h;v���i�M�tu���#�.i�`�P`C���7�L��2�ܙ /^��G1k&��<�Į��Wىp4��L����)��iR���
C�A��nH�r�=��P�wn�dXo��XjQǫ��Sç�R�]r)w: Nvu��a���}҉Y2ʑ�F�2l�i;J�T��RN�)ENX����d<[��HƜd��ۋ&rn�fL�[O.�>'�r�s2,Y}%-Ev�mp5��O>+�9i%�h�b����{��X�Da��/h:��k�W^�6{j����챋�[�0������n�vX��]4e�[.�� p*�^���]g;�2��+N���U��������.t-u�VMo:�wG�'&1���w��U�^�S��=}��>GMD�2�WWI���<rƬ�i>�����=��#L��o&�SҠ?���D��%���xVX/��)���Z��%�>���v��:��{��޵rZ�.�)gن�ޤ��PҒ��*�%S�%�P���$�W<>c@�u	�O&�7���6�wPx;U9�Wvi- W��o�՘�Ί0j�jAu.��1��Τ�c�ɖ�կ���e��
��33w������e�<�5�ْ��ـ>{\�[S+�p�<F ��8�m~��u��l��u>�:�l�-W}y�pY}��O$c��Jx�T�}���|w�;WN�<;u�(}�Y�����s�nM��"R�e��gn^m�38�[gh�icKEãCo��ZȓX'HWv��B�o׿gˇcy6��&��E��b��Aw~u�5�������-!�6�G����4b�"wui�[��e�(��u��swU�ʉ�qq��M��O�W��[Vu�6�@V`[������]ݽ�.=�(d�m^ �'WM���n���,�/���t���#��٠��D���c�i�_"�f�F��8�ڹ�ZGe���u;�&�r�����Xw���]s��5
Eb�7S���,Y�i����q���-<��8���T�	z��^�����q��v��ɪ�|�K-�hu-����V��gM%*fn���Ɣ��̖��ޅr��垹h�y�b����;��lp=vK$��[N�c��Y\ �q�ܐ���n����05,ld�}�{��� �~4jop��Z�_���#�ݵwa���m��F��X܉��Ս�B�^��.m�f]rQs���q�s��b�I�C��S�ɥ|���ە2:�w ����m��oj�5+x����$�n_�ÌMjJ�Zr�Y����[WWvihl�D�ؖ[�b��9�rT���2�����W+<�x�[w��]܋=z�
���1|d��S3���o���Qzb�������:�bM�>�j�����ʝ:�C�4B�B�ku�Ķǘ�M_L�G48sC����6k�d.eo��TBDˎq�ռ&�Xt���9� &feLdV־�M��7[��)c��]�̫��]"N��$�pL�6�kh(�\�� �}�H�	:6�y���ΦCj�7���}�Wv��V*�Ц7��B-�6&�]�c��N�ϟi�Tr��O�����޲×D2@xg.�(�nEn��&(؜ݾ�g:p��HJpB�C��=��5�ѝ�f�H�	��R ntĦ���p�����;}��R=��`Z9��{ץ6x�
��=���*=�fU�ػ�5�ğM�E$%MB�3���Y��u����Q��F���ݧ�f�l.L�ߌ��н��{���eR����wc�ł3��z��ʛ��a�����" NN�h3lni�#(4�y�������}��C6p�k��j�\�R\]�%̳J�	"љw�� du��Ѩ�c���i�HFumΛz�16Z����
=�=:�A��%�^�|�̮*�
��wN���T�#A/3���<o�^����0��.�mB5���;�q���������s���8�r�7HΣ��i�p8�- bVC����n@R+J�����7�+N�p3K���p���[�{s��@�C�&��$�N��sp���ݷ��]u�GE-Q�Lǖ��d"��"�h�;s�O�5�E��3{����$C�u�y��NF�.79�1�)��-�#0�����h�)S��3������P{�x�3rU%�W��x6$��c�ܢ��*(�H��xB>i�,z�T�j�DJ�h�ȍ�B����=
���{�� jGŘ�	�PR�H!Y�V8X��xA�	�95�Ҷ�VKbvR6������	��FhcVf	����J	�����M��.�<Ʊ1Ű� ����SOʅ�D�����������%|ڄ�ɤnf�������<�9��&�X�H(���N��d�%	�.������[�@�
�� 2&A$
�=�/�o�0�.@�sڍb6�� �\P�Dհ��BAQ���%�E��FA���E�E�kA�b�ɼ@���EH��`�P�eNǶ䤒µ�x8�)�i����v�n1��R��b@�s9^��E�LW$��i�NL����*��R_N���
m"�`��6�Tm �2���x�QÐ��l���z�}���r���z��o���łP ƫ*����]�W ��rȖ)�Dɂ��M )�s�Y�B�EkUͻ�d�&�%�$ĭ+	Y���I�379Wjұ��;wkټ[�(���պ	F頠UR�h�lj��
3Q	�N @6Q*."�.��Ҍs���v˩\Q^�ENL�,$Pn2�-�Vm�݂k:[5��uGkV.!������)*��W�t���4�1B��7�W5�!�������rj�C,Q�VU�k��1�p(D7��P�9s/M��m���YZڨU\�F�U�n��0"�ˁ�/�0��<�Dw���d�}~��t$Ȉ�r�kcT�B�\W�g�r�IݸZ �a��]�,7tKj�=�z�����=陏)$p"vJ)83^jX�a�Oh��q��p�K��u%��wx��V�����&�Q5a�Btu��872���)��*�8�����	�ن���k)���X��cr9b��G_oM�mIk�>uԗsx�3H��@��0��3h��KT�lR��S���vg�5����VH����w��b�e{�tv�X2=]̚�7���D���������f�Y��,���vZ�Si���t�����L�ꃱ�q����`�^�TPV0�a*��,�q)�%+Q���[GrH䑻2�`��0��"��2��X���]����c���
���+�()$�B���Mc��%�4�JԬ�u��x��$�ұ�t��R��k]]&-�2�94+j%mT�V��7����&���#L+���l�Z�n'�� i^�a9����\&K �N�e�.9	#t�����f�7�|���d�-K���*�Á�O��$�}����`��l�5����e�A��g�{;Zv��+Tj��؋�f,Ӳ&�[m�B^G��wei�
j����m��r��߽��ǊM��G\��9��M'.T!��9�����2e+�O�����DSyM�[��߷L��4�v�)���7g9�a�r�Xꊙܯk{c�DDݖ�5.`����\NH��2�G;����Z�
��X��͹�B�ݷ��wl��d���'�jq���-u�7�s��58��GѢQ�0���VZ������*�
� B*��w�o��k���p�U-�n �+ �.:��D�*� �CHO�ge�߱���K/�b %p���>Ӄk�lF��Y�S����!ȓ�u{��>��)-J)B��OnfI1�k[�ي秳��7'\�l��WR^���z�i�^�`�N��H��+SO%�&�5�tX)�m�MKYff��_9�j ���N:c�1h� ሐ��.�<��b�������I�]�W���r	1������Ogv��7�\46����է�
a2-L���$�C���*� @Rg	�g7n��	"T����]�(M (N..���Qh��&��w�m�R)l���,�b�S�1��!�A�R>L[�%�YA��uzڜ玬z|뉫zT"�5a᭣�`�ʥ�sʎ�m&��Y���㒔)�L�����Ƙ&4�cN�0kJީ
J؝X,x�ݍڝn婎L�dt����ܶ�۪�QQ7�ֲ����ԍ��c��!�C�x�|�c%�>UD2S�
$`�)�-���6���Q�r4�&$�az��E���:Z�6#z:�јx���)B��ڰ��xo�s7m�D��nɌ�m��9�w����TcoZ�C�L�B��N�:7��9kE�q��IIh{8�4m8�CR�K�KՁ�qH��ҩ(���OU\�VQJ��=��N��B8�vۥΑn�opd���dlMB����m)�.���/XhhD���x���	B-���]<�.��,DT\�1ݬBHZj���x��B�s0[�B*Fǝ~�/Y]Lt
{�1=�����v����;������*m�JlP9�Ƶ�n�FD�����fꭦpͬ��liݐU����2��{��(�!#��<�^5���p�kj1D2@�)���ZlH�*���26��ҭ��gci	�&wӮ�;��z��6A6hݲI6B�_b�F����jB�
N[|����A
��홙�(X�����[	٠���@2NYǜ���l���Z�-`$��p*D���e��%Ooo���mi^�PB��	��*��O�y��cz-�څKM՗	L��I����=�{�������X�A�e``�!�JĮ�&�Z
e}�s��9�y"!
29���4�;�am�q�*W���	
Ԝ��N�`U7��л��B�5cCN]6.���Y���%���o/���ʺ��W�r��VFCtys�s�reSS2�#sh�yi#���&��p[�sY5ܰ��Q��r��0��7n!3&w�6�:�Ʒ��Ӌ9ቃR>XU)����	���^�4�E���S%�85�1"�p�ї��*��[#'P6�#�T!!�4h�SR�+L���-�jB/f3�����ё�Ӵ�:+j�n�C�!R��\se��=qۍV�᭣5"�:�n�䶻i]+TX�L%j*��VZQ5X����!"M�k�%��(��q[T�{pdǩ#���$M!�Ef�p�$��i��!0��{ d�Li��5��aalzq7e��T�%�����\���d4���R(�u*���a#�B�$"�陽����Q�:�lt=cyS�>u6�����aeUHi�XRv;\.��֚��D�ThV(G%�X��ERʜM귧Uj�6��-+���\�EB����HTUUd*UB�����
�j�@PUO�X�� UP#˞��l-�����hnB�\�X�:� [hX5��                   �    m�                      
�?��h~`���r��ٛ���1'�d䭅�;�������96bb7ٗ33����-�E���dQ-��7�Q	;�kS��y=�w}�:��.�s9�U�N[}��B����m:� ���aG�䝞��cK�-l��p��k:J�%<w/�����Sݮ��Z)6+�H���]潍
j�U��975c��st���z���fb=�o9���q��d�1��8��3(3%�l����%��(��/�y(
�z��Ue2:�h�M��
�o-�D��2�s���UN}@��J�*cITS^RӖpr�-2����*�o����vh��}����eU�SqV��[dpB�r͊4s��+����ǎ��{��,C7,\���B{��a�m������EN�)n]����ʲc`�*�J)^����`��cW�Xgn���v��1lM��T�]��"'6��];-s���e���C�75��S���<![zh��d���+�����7�s*x+e�GScA��]��kcr�[U�\��Ӵ��m7�;����$d`�����g66@�PV+u]�G4Ǒ9M0rڸ�.#Tm�&A��+a���	I���ozb �<��;'���vm�d��%TjJY�
F�,���z�a;$Y�-����U[Ʋ�R?:'�i��9#�Bmx������v9V��K�6����W©�Ĥ��	��UfZT�*Z�e���dX�VɊA��
� �L����Yk�D�Dws2�D�P�
�A�m�5["۰k�wk����[2����ѻ�;u��9�`�Ec�"LF���D�)!\�^DG{�x���/d�����n�˪���ő��Y�Ƣ�� ܮ�c�40�$�v��h+U84�l
�R����p�H�j��.auje�ƆN�E��2GY@J��RIh8���UP��4(B��UB���JKZҋIu�r�R�P    -�   H"K,��O��<~�$>%�"�fY�څ�m�E3'��&��d`�,l��R���[R<�Ƈ=.9ǫl��ԩ��5a-Q6�:K�NA����yX�J
��)�u�n�1z�M�܈�6�LE��xn��J0ۧk RЊ��m:Kn��b�DB-��5g��Jdc�9uK�b��:A�oe-�e�M���=�V�asV5�L��(��h�q�F��;�M<k�%~�]��r����^�;s��0��`�$��5*^͵Q����C�t��za�]�7��nX��\�G����"MN�Ϲ��b&Sz(r;/rvݝ�s�A�gOx������rR\#�q�V�Z�.d�4�0�L	;��}xQ��ꯤ͔v����
����%?U�Wxg�s�S^||���{��m����w�5Dw��l!0�	���O�o��\�vz�7���7��)�Ӄ�u��y�,��{�̳�"xp�U����|�f5����݋�@ۓ#S��d�"��낃dt�F7
i�h�L��@���he���0�|�ց;�R��1����%Ζʸ`��2�O���%��{�v�gT8�0Ajr�9"Sk�F�h&v�������ts�zGx��akf�!�܋M�;�*���Z9Q�׃a��
0��l�h I4-��g/Z}hXfY����_#��ѽ|�륄�R����Z�&U�i\������H�l���x�~�!(��T�xcj@R*a���J>O���<���e>7g� ��{��1�[�V�����2�s&��;�笳�
Hx�<�ĎtV�jG];jveB����3�(���ҩ�P�q���0�/1+�W�.�9�����y/��vD����<���|��J�~͛ճ+m���6��t��=�{�����`��� f[�BX��w����2�VՕ$�' �׫lVX��`�,��9�*;RyYr��l��^ߺ��pn��
�ݻ��+{fRh-�B���+���	5J05d������,����ބ)C����YI��חI���LdHծ¡��4�������h7����x`�;əUU~�0Yi��upsδ=x�boS��x���۸!�>ˁ��^���3��_Z�}�s�"�U"B�T�uta�TH��IG�y��2�nK��ul�owv�%3U��<�=g*Xஆ�߯�>�5�JJ�>��}�-x}�.����_K�~Tжy0��xw��	mF�=�.��W��o�w�o�=]��Zv�F�'���<B�7d��<��wg��)j��#1��xh��<Lw���5A����i��#��c��[j\jP-!���IV�,�Q��mN�Ly����s־�ʶ��a��Sw��M=m��M�0 1V��O��y��&��R�,�J<��R�Bo_tz�ͽZ����sAC�f%*m�7x �و��3;c�Bhʕ��,��b��yL-���RB*+x���P"rz�Z�glJ�em
�A�-#R�t��D�3���q��T����̏�Nl�����gm<ܒ��������Zp\�F*z���o}���C�I�e2��I5gw;�y��b����%��o��oIw�{nWcj����������-������__�*�7�wٍ�-FT�K�;w��v2�&�}�w)�*��k*.-�k���S��9vfL�vt�κ P!�~K�u@W�� �鋤��h8�:h������Ӓ�CAidpM�~���C�{,C�6�ܡ�>�k���!��2;ۼ�m��&R��mb+q�%	�pgVm�v`�p䛺�� 8𧳘^��>Z��ª�7cuH���lf==��Ӽm�Яxu�~��x����y�j�׸���Ip#Hg5��>��ŠT#�&vY�x��Zx�W^�ν97��b(�Ob7��4{�O��dS���A��/xE�6j�7^� 	�7�^��y�b�@��y�v%�G.�q}�qn���q�{��2��r�;���i��&kr6q�̼�F���z1��Vg\U�lQ�<�����HjI�&;]��,ߵ����ID[�ӮڙtܑWi���)it��˼��fMJ)�+Q\��Zi�̝����W`         H��T�U����
Nod�^R��i`^���P�� ����,�}��I�n2���@J!2�QF��Q �ORm�k��s��뭄�i�e,���l���5bcv���D��v*̲W]M��|��u5��3��dq��!"1�*9(XFU6[����,��x�<uF�k1��Dʅ"N���
����{�O�3ݐۛ��Y�'oAYYUf|=s���z�e-Sq�P�#/�����Mw_��n8�B�x��^Zcefڳ��u<�|���f��U-%���:	��u�y��w��<@���/���6�ͅ�6�A�L.�
�c���p��s������;|�l-�z߷�ʊ".Y�Bw�辋̼��j�&�մ�����
�[u۲��~ӌ���1��o�}X��xu�W�Q���Z�㋌�F`��헏��a�JWMci�b椥<ʹnWoW��z`�,m��x�o7�m�ug�r	UUW���$3]��'ub*8�FKm�rAH��H�(�שܱ0>��Ԍ��[��\��(ȅ�l��p�.j���ٺ�)�Ѱ���!��W���R�F�L��Cn�po�g�AG�..��=�婂y�YYj�%Y ���A����&�����.^��.۪ � �A!�E��D �A2��7
�gA�7w�n.��ޭ��89���e�����G�Da�RT��S;EewyJ��ˋ1��.���Xz{� ��FF�8U�[�A,ћ Ƙ�Q�ЁP��W�hiw�@�۳�ޱ�dj�C=���co�<=lxd�Do��:,��p���]`M�� ����5�U�{M�Y�K�Ѓ�齼]{�x��}P�1����ʋ�WD�Nw&�ur����Wl	�;�<5��u�#�DE�*�e�l(H������L��IǎZF�"��uA+UӨd�;X&�Iq?I�[�Tb���Wze��cu婷���49�@j8���ǻuK�D8���eE7v�8��
�歽�b>'*༫���Gk����� ��J�<C��׏�����P\�������/��6�+�����5��v0�#��'�:�ǽ�Zf�j���6QØ�H�T��7����jcw���u�ꐼ�fgqc��B�W-�@j���U������e����9�a�pQ`ku�o~gwQ��W��]m����ù���KT��ET 	�罫]�YLy�6�=[c/4	���������˜��4��C�Y��,H�z�!@z���Y@��_�3�?bC�65D
��K(�k����}V�yjL�P���^eD-ݟ0��c��,f5���@E�ήxxe�Ja.�#iI�����E��me�`�J�u@��Eq1WJ�������ϖ��٬XLN>�)ר,𑹺���Ma��Se-�^��M���w-����O�����}m5�A�X]SN|�U���y�IO�8��X�m�h��~�c��u�F�trQ#��:�  ����7�
c�b���äz���ټn���[��|���,]Qkt\���mY�i��ܕ�M5�=������������Vm�#�ox��`�|#�R�Eݴ+\�8�K�"a,��\�����u�@�)1d�BU�� ��*�kܬO7�'�d�6��Ծ4_S��=�3y!W]�SFf�e������)X��b�9ُ�{���x;s�l��Ӻ�1�
N@��U�4j"�&õW3�w��ۜk�K������(�$n&�BA2�UhE�hY#;b�4����fD��:3X�ڸ��snc$�\�X�ʠQ5���Vth�h�\j޾d-$�\eJ����5A�}Gjg�^���0/r�"..����#�z窂E8�͝�����w~"�>C��v�0Nm;�4ь�=�kB5���WdDY�{D?o!��
�s�b��y+�ܡ.S�Ms�, \D����e9�����>=cj�eo�@KeN�^�a��=�ӕ��%��ym���׎wٵ��K�I;��!�Uk׮I}�͝�[��c�[�pf�;���d'�p���}�̷}���~���	\w�(5��ݬ�E��$�@�3�Wy�\[	�코�v>���W�"�Z�[v��vm�{(�(��;��XB,8z�;�+.�DP޵��g��10ۦ�:5UIX�K��0�P�@  �     U{�:qvx=����/�zWf\����S{�}�1�K�U�y�m�e���xZ��ڪ!4"�$�nW\L����+lr"Z�*#VQꃭUFӰ�IjeewN��V	�]�p�5�|1�5r,��;$������P��X��-���H��'7'm�N��xGj!Z4��-�8�Nۖ,�#Q��OϽ�r��;~=}T��{�2	�s������}��<�K�cQK2~�[�
Ifo^�݇~爘���P n����^�W=�e@�O16�}���"�3m�ga�nN�<o��^�bEB��NC�����7��m-�.�H>� @
G�O)���X�%��'�{u�~{p6�ڹ�`nm��-�S��X
��$�2rJ�����nw�=������JL��@�"�$.]0;/��q�0�3ݎ���.����x�w����F�0&I�>Ŷ�^�Ux\%s��>�LށU�Z|Ѡ *���{xV%���M��3�^<},h���|JvHø����,q��䣍� B*�pm(C"V@�R��`3�p�=���Ro%l��OM�Xb(��7�i ������ޮ��*�4��]h��.��?�/'Z3'��=	8Y����u[e1z�P̌����@t�&�3<���v��� ��lD���{�՞�z!:?z��r������ʧ���*{Eˎ\+s0�MK����(�P���؇z�:��=�뫗̼��k�p�=#�t�J@��u=aS;9/��/��Λk�N+.��˔�GD�N�n� PTZ&�i|�ј1�����!H�ko-�6�����ǋ�2f�A����K�hO����9����޾f�ꂾ	���yQt*�2���{�a��b��qrf�1�l?h���t�\]�`����yl��M."=K�Ax���Pw3f�*).��`(�"͹^+w�KdI���!([[���dNX����ƙ���itc�&귤uda����=k}��"O�O���n��<��.LG��x1�,�di]eP��}+�����Q<{������`��T=�Z�T/�)c�{k>�.Z���g�ܿ�y�����Xp$��#��EZe��r�c��m^���B�́.�L^�q�]�ޞ6�{����Z���ގ�f��I�ݔ��r��/,ؙ�2�9�ܬ��o&�г��Xw>'�_ r�}$��,,C�-�'���}�o}�:��?]�2����$����A����q����3�	=��X�{$V��ml�:us&�.�Vݫ���G�X,�cG#۲�BU��;�θL
�y7G� ֜����+TT��9ӝ�v[�aR�v�\��nʱ�]�wDɍm4)�e�mX�t9�x��}p�>K-;b��ޡ܌Zq�ēD]X��x9 ���G!�2��fcbc�D)=����S���;��B�A'�rRu�R�Xo��n�[�c�X�B�z�c(�;=�]�Y�k<�������4\ԝ�Wjk�� �iʕa�j���KXU
��y�7���9щx��1����]�ƫ����g��uWt*��U̵��M�Ҿ���#{̺R�쫻bB]C1��sl�x��������������Ļ�4u
&��F���Q=a�Xlvլx�x��P����J�26�}�{��.�;[�*��"�"���^j�:�.˼�:��S��
[�1w�����g���k�aQV�T\<���R�LԸx;��@�Q4��O2�D�QUD(5�R�NFy�p��� �Y$iݢo����:�SF��P'���A=���i���"�;�	'����v 8�So%�M�U%]�l
�t���k2��[w���y�"�Tֱ�����{�#0�:8���{��8��7����.=���׽��s��F�5�Z:�ģ��l�%M`J�{v��ֻ�a7�ͳ�i�q�U�6I�k��Q;旚�"H�]���h�Zp%\ė��]Gq�p=����`��ee���u���%�=Z��h�yk!e�HpQ_nr��ë�A�]��{�sU�X����@2΢9|�`���nt��*>�R�x�-�g�5ƻ��ĎS�_j� �ڸ5�aV�9&������|j ś�QJώv�]�B�lL]ۉI���j�S��D1�#�q���)u�����?v��d�K
�#�R�f�l��'�y�b�s�uX���ܾ
���(�~���CZ-)�X�OȅQ���Ud0���U��P����MĆ�Y�Y�$�1E�E{T�(RA�ʃ�i�{�0 ��z����;�Λ�~�*����';3�.�j9�/I�9�w�*�$ok��j`:D�\��O�b��GچE�QZ�]Lc��J���a5T�s�V�P�w��7O��?��Ȏ�����߰��:wT{��=T�F�(�@��Y�XD�˧�!�ɼ�lY#ꁬ�٨ZL1E'&ھ�+Je�l�^�6�N��O��y°�RL��T3�w�Y�j^m���l�m�;��*���ڠ*%���?b����DHh��)��l�/��״�	��؆���x�J�f���O���i�@&��3dz|� 4�ة�c���Cp�f��<�媤�|�Udx�ț��(� �^�^>�}@
���Vy�	�zi��I�t�g�f�[��5��ϟW�;����)r���?b%bQO-�G�,���F�q��B�8C>8k5ߗ}}����f��LB<z@f���������k�wݾ�hia�%T(r��'G9�ݽ�|�Fe1�)dN�L�����V���XE���q����x&��L�Pf�iS{����s�!��:�3Փu�1u���>�>#kh� i���Yr:C:B4	�x�{����I��'�bMB�;�B0��v�H�EEE@���		�5T		� x�=�8j�	��Ej��(4�L�
;��$<}����U@xЪ��ƪ���K5Z@�  �S�� LTB�2H�@MXj�m*+��ʨg�
���� ������WH�����t�]�� T_E1��9n�+ՍJܢ(�Vp��V�Y����(+�j�"��lP&�"�	�-�EE� EEk� F�SJ�	�("(+���Ej�48�E�'T				1!^4��uD��гC"�"�5@�@�A� D#Cj� (�@��M|��H�H��jqUEEE@�S"�"�4!@�,�m
�:DU��3H٠����4�E(��2((A����B!"��De������ �		DP&��&�hHP$P$P'��F�EE@��5@�@�@��H�H�/�A@�Y������EEj�"�4(��R�m
���M ��A@�@�M H�M�44(�EE���G���("�	�!@��@�#@:�52)���<B5@�@�B$((T@!@�@��H�M��3T=��v((((T	�)���xg,�9UP$P$Pԅh")@��T�f�DP&�(($�h	��@�C�U	ߤ t�Ej�"�5H��M|EEE@�)@�ƨCA��#T1*�DP$P&�5H�EhQ	����)j�"�!Z r!@�&���H�H�H<��M��EEEj�"�HH�ha���H�~�b�"}ѹ`((q*�ԅEEj� w������c�Y|�k�P$P$P&�(jUE*F�	 ((( &�		�ޓ��D!��EEEj�"�"�5�UL�Q���� #T				�6��H�H�H�����m
���窐�E��P'ƀDP&��	!@�d �� DP$Q & 5@���@�]t4(Uf�����)РMP$Ps�A@��H�H�䪺i@��O� ��H�iV�"�43��ϸ�^����Q�!DP$P$P&��a�&!@�C
"�"�"�L��			 EH
$P$P&�((bB�"�5@�4hP&�($��Ej�"�"�"�4�T�+�@�W�0�j�~lP&�5H���@���B�4�R5@� ��H�H� �@���D������2|�0ðb�@�@�@��MT5�
��N8EEj�"�"�"�= r �u=�h�h
��3���((T		����5@�@�� �P$P&�(U��$P&��g ������H�K45@�@�@�@��H�H��	�!F�((j�`h�@�>44�T�"(jU@�@�@�V@F�$�DP$ �F��
dP$P�PF�4&*��((5H�&�"�"�"���qUEEEj�"�"�4�"("�B�	���j����H�H �ڴ<�Mz4��P$P$P$P&�\l �2*���R 2)A$(Vj�������MP�B�C"�"�$�$((((T		�F�(�U|���6����@�@�E"(u!@��H�M �"�5B$((C�� !�H�H�MP$P&�)
���hMT� x��S 	�DE@�R U�(_Z�dP$P&�((T		� CqU3H��EEEE���>�G
 
���MW�P�H��o5݊���	"U@�f�EE@$SHP%A��B(�		�F�����V�E#�@#T�"(T>��E@�T��MR4R	�����ݒ�((T-!@�@�@��j�"�4���MP�W�U�pP$W<�2(((Ej�"�"� v� �0�		�5H�Eh|h":@�E$(T			�m_������{����}�t���f޻Q����xj4���& ��(��H"��g�Q��P���        }ˮ��l�f��c���t�_����WY`v�R��z����=e͸���ҕ���ĊQAF�ꎏU��JF%]����*�di�d�`!;i��-wS�b���S� �2����+m���B&I,�:0���B�]I.�\T`�	�� ��P�^F�|ˏ$�cei��'k"��������.�ʊ	�d#T		 j��			�՚�� ��H�MP& �5ƨ��H�H�H�A	 ��j��4*���R 0�EEj�5L�P$P&�᠍E"(4�dR5@�@�@��`������"� �F�jB�4�"�4!���ê�H���5@���tҠ!F���3��@�H �(X RU@��:��@q�(�@�@��H�A�R"�"�5@�A�jN�H�H����C>�v� ȠA	����	*��B�"�"�h"(EEEJ����HP&�(B�EL�(�M+q�			1 (�J5@�@�(((T	�  �B�5@���� �:@���H�H�H�Mt�s=<\�"di,ʠH�ąj�"��T4	�>H��1*Ej�4	�H�A�DEEEE��E"((CH��a����HPąj!��:�9U��((j� !@�@�C�UEEj�"�E�CT�P&���褪��"�48E"(U�S �T			�@"(b@U�(CMj�"�P$P&�((D�]lQ4(�Ej��EP��(P�"�C@"�J�(((0�A9 �MP$P$Pi"+�L��4� B"��M MW"((KGT	����M#T�P$P$-Ş�K{=>k�G�Q��}�3f�\�N�BA�@�F�i;�҄���� jBg��@%g]H�*�i�d_JЬ�⮘@"Hɂa�c&)n�������Ƀ8j�>!g-@:o�4�E���%UU44�ƃ�Ήd+A�~�P����[i��9�t��q6Tms��TZ}A�b_�B���c�b�x��b�B���=��ӝT��xE+CNr��V z�"�E�Y�5f�/���3U[���#K�V}|sݿ��wް8B=�Lol�
��(�.!��λ:�k��;,?!��d��#��
&Q���M�w���/�=����Y��!�cU�0;4fs�>��s�� �D|Q�B7j��@�%��L%�2�ɹ�0L7uVKn`��j�a�+�	��(j�"�E����w�*7�H��Je�k)���ղ;-b�&�B'D*� SN�Df�->" t$'�2����{쁑���ܳ@��00UC!��uƃ#��%�h3XV�$�I�|p��R9`*�WI�G��0���9�:Tg�5|@#�aMYA�>/�ﺉi��(����(�v�I��kX����kx�2{�����U�G=/&?��m2m�q��s���d�jv����9��8�[¨H��H��XP܌�F]�`l��ؙ���}���V��x��{��*_��C��g�B<q��- ���B4,�k�'ڬt���@|B/�Y��Y
��Ӯ�E�$�;�_�	��V�m0G�"��������*+h|Q�B̖��С����B��Bh?���L�H��d�k�2���!�K5s8�����)�fB��i=�36�|�h4:P4M��4�Ǆx��t�����E^�u�3���cy�AB�u���͟�X��2���kz���6��IM}�:���Z�o�٤k(j�
t��>!�h�@�|�����ܲD�@��!<�-	�ɆcCڪ~>1�w�����^O�ш�z����z"˪������Ȗ:ƣ���e
,8�WCڀá�`�Q �F�Ht�3��dY3r�_-t�d]�(P��?Ҵs���<s~Li��<"��z7�Z� ��x�#v�e�:��j ~��1�Q���"�{���u�{�o'0��� >���
��!��czbb�����$nQ�Z��#�^'ͷez_��|�ج%EVD�/ؘ�(�E�!�q5��!i���J������t��"��ä��ݺ }����R�=�#�����h��xЇqWb ���
1	�͛8ibea������F�l�zB5����H�Ξ�}�0��-�1��9)z��}��c�`��L9�X/�?;���Q労:���ėkk�>`�$�@ԫ���@&@$%%y�ho8���l�o�xxCeܼol�K[�v����Xt��$I0J��Dj���#�\L�@�+�P�f�>��0,ւ4DT��x�5�#Aر�Y��Ǫ&�6�/k��T��g��u�$[f5}$�+s��IR�,T>�B��V�M�ɱ�m�!��x������s6�*��`R:�wD'-ޯ��tq�i���BM�4�4C^�*��h�U4�-i׌4�]�
����x�!��G�xC~nA�$C�@�f�#Ϯ��"׏�<�p[�,@y��	>zI1
&����dfz/�=6zt��Å��GH��פ�f*f����|Y���y��3��/WEU��U#xBa�Ad{HE=�� �yb�W�Xi�"�l^4Y�L�f�**E�V���H�Ks��η���`&�a�4���C;W[k��.�Ԥ����d�y�"Z�"�凩a�3@!I�k�U-�9B�z� �ӗɤ|m/�Q$��8�� �,�t��@'`����㰄CF;X�mFU �d�k�&׷<ѹ��E�CX�(�!� ,���$@%�P�i|���AF���ǡ�������XڊY� ��Ч�S�ֳk3���fw��a��S5��cF�@������� �Ė�Rr&��}�P��.��1�@F��O5D�~\��7�e��}�[��p�i���h��ښ��Y�f�����Ȣg�18� 3H��k����56+��/���a�8��h� u)��� ��M|o��s�v06՘�s"O�6"0ѳrU X4��
���C��H�Bv�!7Q0����� j>�Q֠�����l�F������x��jy|a��W�t�A|�GƔU��#�TϏ�2C���Q]�x���H`M�h4�Xa�E�����C���Nܞ`x��-1�%�R�  ��$
$Q��f�&�H��/!��0�޷��!Ü���H�!dB(ў� �VEI�_Z����9�w>S,��%���n����\f(w�˚��V-l�%�T�G���k���J������*PS(")hP�B�(���x9S�x�{�0�]w]i;�U�f���n$xv<!�
-����Y�b�z#�!��~8rc��T���1�"����z��a+ 4�U"�$C��͚�G�TK5��%�l�����`�}�{�e�?�Qq�!�P]L�g��	����:n�b����/ܖjI"�Dt�7�&�"��|ܼ���,�D�*A�sE���4[�-tM�# NF��j{��,uae"6����k#�.����"��#@���j�)��\HKD�	�L׌,ys�Cϸ�C�믭p@�5��֛4M��7S$Yx~��<^�P���j��q�<#�H�GO8��Z~�f�.���Gq�5A3������F��\8в	D���5��������uO�n#�@�Ȍ6� �;����J*���k�B�"U {�(b�!�C�{>i\�����ƆzzL�Tmjrp_y�zj��Pb��6��ђ#F��>�@��Xq/�4�E��F�Q�HD4�ڦxa�^GW��PքU��oKO��}�YX�0Ґ����co�`e�������Ԏ5�*/���D6֪�]|l֔�Y�'���������<��Օ��4M��qK��}��!Ab�8��}H���DݠȳH᩻�0ՔcC���GK�t�(33>�"�#��.Ƽ��s>͎��L��o���t�� q��$	�����lY�F�����h�5��l�f���V��L?eg��;F�Q�4��dp���<G�ճ8����0�©���8i��:�?-�dkA���6I� �Q�+@"6�*~��-����=:,�|[��#O;m��;p1v�+�wYڍ�S�;OJkN����v��� 0�H@E(*�Ӵ�AZ         ������)�ZBMSt�S������9Lʓ.��>=��*DhPJ�T���Bu}n�[��,�&�%{yu�D��J�ng�n5%j���e�j���'UjWiP������qj�Kt@���U5QV��R8��#>��"�R�5���X�j:��Ƞ�@"�ŖRw)�(�n�����b�uJ���E) ��q!�"�_w{8�n5��3��V������xh#^X��*uWŖNV���P�����+��Y��a�	�*¬]]F¼�Ư7��`u��p�y���P���`Y��Gґ,�'� n\�~��&:Ё����ZK&���5��%z/C8�9�LC�C ��Ƴ��.޺ma�񤖎t00��x��e"XP"�(��
b��Ϯ��Kئ&��,��gU@eD��HCf����D���x�j"a�1�q\�$
b���/�L��P��F���cʑ����� W��f����t�� ".�!���\��8�%��B7�'��ύ��ݾ@:k�kƛ�.�6{�d�4�2�H�8�g<����Z
���<hY$#���Uܴʔ%���jd�a,�N��Y�=wx�x�4�T���MDI��u�C���g�b��M#�q�|t�C�lCk~LB=�΄8|X�Au�~����b��#���4b��B���Pf� ���Ȣu��ުɖID M��_Z�D�HGH�i�>U
h9�K_u�T(wv��:tw�di�6k��#��N�gA��C�@����kT�-h{�Y�Z�%~m*U
!s�m���c�Q8q�F�qMR7AYt�}���Eq2	����#S�f1䣬����p���a
 ,��F�,���Aq:�@��`4O~@2!�3��Um���T�>��f;��7Y">�ud�y�p�����7ͪ���\ 8t�~4�a�����b�g	#Ŝ:i���({�B	�:KgB2�WX@&�S@x�B�G�?�Ā���J�}�͋y����BK�$��r����o��������Ft����#����8���U��]��j���qҮr�	� ��{�Nٱqn�r󝹲W��y����,�?*Sx���>"�@��,4!�-^� z*�V{����>�f��GHQ2ꆺQ���c�����lv�z\��r�4E��{����� "#Zh�V�t��=,�&�����"�}�t��kㆯfKu�3��>�B�Q��ϐ�r��N�,����!�e�N (!T ���	|d�"�i�tԵ�~4؇b���?�>�!�RKY�D��O6I�}C���]����������C<��dv �x��8l�s�8F�a`�Q�Hguk؃0�h�G����!�̫& ynY�������Q�CY�ox�k />����� cB�(@t��p�m�h�#]�dY�K0�u1�"f�Viyt�U�o��߾�v��#m"5�A	�4	���W��@"!�A�E !5Aw�	@�!�q}��	��*��=u�&D5�J��>}}�������Q��&1<znev�W]DE�v�L�Im��CmB�Gƨ�!*�,�QЇ�Ʀ��=@YdB:Y��>L�*�?*C;�B�a���k�Y��C������寈<CMG�]�gܻ���0�GmLT�/�z�!�V�p�`�j�� gLiDQ<�L45*��vi��aW�����Q�5��7�hs
������"����u�=0�D�E�a�o��z? Y��xk��Ӥi�B��]�ř�bI�xH;�v�s��X|F�T��� }�!�Ŧ�m� �>A�4�t�H �I�DQ�h�k�Z��m�в8A:]�@���iZ�7Y��	 �^��߽���9���
I�<�c�Z:�VJ-������)+��=�J(�IU*G9�u�[��yV�s�z"{
y�x�n�a�Ía#ƙD{J�Eڠ��([di��:�V*O���d�B�E�	�t>�c����#� 8F��T�E�^�9�P�쌭�}�3]��0DC �4�h@ �AsTA�� M� ��>!F��H�W���da�F�8�kx�e�Z9�Y>�dv1{Rt��5��e�6��y�'*B�j�F���a�4��_+"Z$-D�T�T?���A�DƆ8�U @F�n��|e�`)��Q]�Xk��BZ���$",��a�#��D����l(��5#>�0L5����N��}�m�?����g�m j��$�و۫7\ʦ��r�V����-���x�ƽؼF�ل>�����<Y#��t�n7	B4��Qi�"(�|�`{ �}�8h �` 4	��v���� ��8�C�<p">�=��^�5[�ԍ2�3�Hb���i���>�?�p�W���:�s��� �Q�Ϙ�>(Z\�$a���Ŕ����6���yw1�M��SD4��}hC@�y�P� X����3�wh,�Ҍ��ب?*C�]��Fb��I^w����PGs�5җ
)!�9��@�~5-@o�h���Q;���Q��h������B4>0�j���jZ�1݈�6�ùׅ�A�[�e�>��Q=�U�|/�Q5Ӆ����ӤYæ�/X��52>�p՚]_+� ��*4��t��ο����=⯺#�C?�}�G�Y�' \6Y�qadtb����!���?6#�2�pK�B�^E��k�����v�+���$���td�@�H���LѼ�xPП�ζ6�#�K�ޮ���h�!#MUPdbpD�m1A�c��� C
,����͡ٽll��6�u���|���sy��kN^����E��WCO#V]��!�k�k��NOY;�B*��Lj���G�14	���I�5Z5�f�QD��h��o�����y<��������Z�AiD,��"�&I���A".u�Y�qV4�t�І��:(R��	���g"Qt�[��� #�	B���:X�@�5TV�ݴ��6�8؅������ҽ�F1��ȖXj(���"�"��	r��@�+�LY���j��e�O��u;B�U2��*��Dŋ���l�ha�B#�q� [��@kB��`�EbC>(Y��%��
_6�!�(����{8j�z��t�4Ȟ�2D4	�G�
~{�6�G����!�>���T�#8���z�i n� �ա�iZdQfs�aҮ���G.R��z\B޲�{����>-!�����@�]8��1�I���:@$i
*�\4cDY}��P�$;�ά��;��f,5�����G���D@~!�=X�?w��\8BCƝ�`3�20��N  .�� �\��d�ea�@"*��4��i|���b�f���^H3P��?(5}g�}�=���h�ީf�B� MT~Xza���ϖ�-����414�P�P4yi��>�`B0�Ȳ�Yg�9'mny`W�Vx.���& !���#`���VAj}�a@���S��0"Ҽx�>�p�I*�,EW���w�gz��H���N���UB5aa����p�r���p��"�=!��l������G�ثꆉ���He��#U����Zx�	冈�%���0�R� ���PCb�6�rxx��_+󁨣���3F0���U�����.��Rŋ�$X�lc����ٺO=���2�Jw���e�W�GS]���E՛��޻S�}�FOX|t��cV�sdh�2C�!�9g�s������Su����軝��83W{� ���ٸ |l�.Y|M��&����K���w��J���ו��r'w�����׎��]�9Y	���H��vOs�۸�y�kOqX-�m��Ө��e�Ҫ9�뵡���#A葏�UȺ�at7��+V]��ح�3��6��k~)�y��f����QE7x��胔f�pˣ+LR���>�|]�QPz��.��;e=I#���iݔ���*��Spu�+�X�5o&�h\g{f�]m���]Yy�V������]>�?�d�6���z����Y���F+��h,˻��[v�Z1�D�ێ��~������mfde���mI�1������5�zU8�N8����o�^�֦K8Y�����>��w0%��w�M�.v'�� �݇�C�S���W&N[�-�ɯ1I%�5#���Ss�*�Ɲu��a���I|Z{u[C�
$
��b h���͒�K�Z���5-�ê���܈P/�a'���h��	��x��Q����U��/%���bb!�%�&��X�1Ҡv��V�r�l��6�|�8�y��T����ݕ���bq6�	-��Km  JW�E
                                                  �P$s�����Ҧu�.f�un^9�p�z���n��Wy�m텺wH	��7N��[;i��*/r�����(Q�Xn쵬Sa���6��l�E\k:�[ƽ���w^;�=ơ�h3%�e�%�B	�`:�EZ&jW>�WE�u����0z{�N���i��1�!t4���23,�d�I���A
��EC$h���sf�;��X�̉��闎�t��V��hV=J�J��K�["wjT]·v1$jqX�5�[+�����i��d,<����g����.@��
*�'W�ʰ�����<�\u�U��,q��"�˷�ܛJ���(�����\��!VL����a�����
4IW�c�EUѱ&�\2\r�;x�=�狿\B�Fԍj�{9^dU���:K�T��^ꕫ[p���=���m��I5TX�#�B7��3N4��Q:�P����6�N6UZ�ڨ�i�5m�vK�DԒ}����p�=1���mQI��1�Z��v�Z���߆;6[�6��j��ypzwq��}&Lq��WS�J�`,m?����_�2��X�e,���W�3UB�b؉�\���ʪm���0�F�)��GX+�KR�#`=�̖���E�ٗh�#�w�N�����������z�Ad��f\
��v�k\����F>��5�;��8��g�Q�J��r�*b�6�@);�����Sy��$�N�D腈�U��΋�:�}�*�p�	�&0,4$Z��(]Q�d5%����3�0�\MF�R��/���8��Le\LT$���1D!�8d��w5�1��&*m@ۥ.�L����aj��q8U�$d�(�,v82E���2+b �$��EY�����pqJ���$�B�,h�#nT� X�l�I�B��:�A9J��	$yrKSN�        'r�I���.ߺ��ꜝ�Úi��Q����*�c��Խ(�;�e��US<�d21�ʉ �L�U,i���hBVʂ&ܶK�#4�d`�ں�J[�+��ޠWE�s')"���Q
Б؜T�2�+AV�RƉ�)U��2P v���7Ef�ky|���B�V[Y:���X"�I�����ӆ~�� }�:�K�>�:��)}��dB"�c��#���V_� ��lY�h4���X�߶P�ܾx�(����@F�����_�;C)��>�5կ�|D�D#=��}/ј�L6��D�=,E�5ϸ�ݝ!�nO0v�͠�׷���u�zX���4��g}��t�4�T�3mX}j�*-0��P�Ul����qP-&���&���`���}�Q5�2_�8����K��}D�%�}�f�٤Rc��Q��"$-/�Qj�qGo���8Y�|m�4��P��Pe�_C[f.*P(���d��c˫THf��y2���HF�F��4J��xt��k�(��o�"x�E�tG�����âT��"M#��F�G�æ���Ohϑ��Qe�b�dhu�H�(��N��� �/*�dC�A�%��/���0vVD��"�ŵT�x1Cލ�S@g ��_��\�5⎐H�f��h��M<�����ZHI�t�+��6G�5�:���+(�/�c��Q4CC����'����-sF�1nax}7sۏD/ �G�4���p�>��<��H��W}����|\ZhP� ��Ԉ_%)=a��d}4֍�m �W\�Ő�șe�=A�'�@�N;F����0�^zǨ�b����X~J�lbUf�jB�� ��,�3�9���:i�HG���H���-�Q�ke���[��������ވ��8᫶�:�j��f !F��Q�F}�H� � �������p�#���q�T�ƺ{���(�L�Y�sS�p�5�����Ω�9��8M��Q~�FdrD�����4�j+T�6�
��Ph豽�!֚A�9��M��A�QD�8�zi6�h�� }C뭪���>f:�����9�!e��qR�e��5�a9�`XS,�H_+ �⩚�!�O"�Q���F%<����~C��,�$�F��2,�Cª�b���tٛ��<G���"4����6��1.C^<"}��쐒:,��dv��jZ���;�g1�F���e�o�]��xh���XG��Ϡ�<!pj���N�,Uޅ�z��s'H���Y!���}�:E4�t�&����g�ݨ�	J�hgzɦk�A۷��5�;�<��4��)��P�k���K4Nb��W#xw����4��I�#Mk@):��#衮�G�"��V�7�u�?M��h�6i��BHi�C���a$3j�:J�ؑ���,5��X#��NrW�1���D5ֱ�5lJ�_�_��<�[��nsn�Cu��5���J�LP�<D���⠏MB�u٭�uL��T�h�_�;4�"KN�@",�v���`^�i>A���i�3J�-�2�UX,P�J�MV>�e�<����ZrAB �k���c��R�b����(��\틡�˾o��È�"�3DD<i�ϐ�d|9�D�A�hQf�I���C���
�X~0��Y�|W��o��P�֡���l�@�T��Z��4�do	�=(�_��!ptT@ǵ�/P�D!U�Q͌z*��i���'�W�uG�<�&�'�B�S�@F�D,�D�*dx
�"�Aޱ�mMXe�'�3d#d@��T�])J���T��dVz�碘ZDb�{�i�G�7���?��Z,�R5��eDU�F��+~'\¨"(~*�P����г��;�B�rλ=:Y�;�m �ͭF���=A��ֳnn�&Mٽ4qn��]�������>���[,���=��5��<���7�s�ߧ��'� Y�ߛ�� Y %uz�B�)})����ൊ��B>j��h��H׊!|~�5.��`Xtd���ZV����ͅ�Xo6QX�0�_<,(�� $��|��7��E"��q�cXh3DE�@N� 3XE�TH�@ �ß*�{�#� |Y�gm��k�49z\Hp�S�� ��(b�!�@�
!��Cg��hQ5ؼ`��F�
4N�|i���:&4��W-z�GT=#�>�-%(��D�(�'����ePiB	�����af�%�DufD���ϘF���Hw�y.�a!��HI�dY����V5-�e�WTx���L���c2[`w����$ߞ��ҎTK 2"���P5�B4> �1S0�9�s���Ӳ,�_�1x�����@v�!D�HC��<�׹�?��y�ͺX�a�:�2	CI����~��Ϧ�I���]��Z�dC�M*�(P��Cd�p0���%_�4���l�PHj�G��lQ�I�u��;�M��_�L�q��zX4�r�2���(!]V~#���)BZ�$�Q�@S;�e2�����8C"qK�����g�WH����,�jo�+��-;��� š�4���@�p��!����|���2�QΠM#��bK�鋚��h�G�sQ��5���B�0L#~BuB/��ޮ���hMT�Ǧ�*@�=��4�z�mv�Vl�nʳ}�Wό�af��^��h����ɡ�/}�= P�_MjW����T#�UքK%.��P0�F|�#M�8C6i�,�51Sq��Օ�0!~�͍0�!��wt�x(�6<�"�Ys��2?:��ʻy�zkyu���n�L*�D/funn�P�t���B��]�%w�Z��!X�����7������
�*�g���ƈ�"�h/&e���zc9a�M8w�^�u��)�-�~�{�3���( 򧎷Gb�cv��h����x�D2�#�k���7��t�e�ƢິB�"ee������O1bC��pB���LjT:P-"SU�EH���˕�(�4JhR�f�â�C�G��'D��S��Y*����u*��{�l�t����1�5O��/�q�[�і	h�Q��C>�@���7���:L��Ǖ�Ƕ���#M�[��
|sx���r�K��(��è�t(�أ�T[�^�t��T��6�ԞxE��{��q��Ǝ�!���(������HL�ukj
�&G��qzF�K�4���5�F����PڴZ4��Fs�D��I��}#��<�0���z�{
^�/���w�UǛ��bY��-YX_C;��};��2aVm�p��a>���n�F��cv��(���ns';|�y��n����B�X 1�Z��6�����T���5,����j�yeM�$eW<uVo�~z=�g��F��mn�аLiiym�v��e^�i�8�sL���o��&-��c��yϗC�>l8��Y�V���5c�HN����)�?�d�۞8��]�áB鲚a�Q*l�(hJ�" I
h$�ti�jn�m���        ,ݵ>(��r_gm��-xy⬧Q۫�++�s��xw{{/N��W��-Ǚ�媨�Y&W8���H�f�җ(�u���C�7tH�ى�Tq�qI�]�9+g	�54d��I5I\�Vk�02�}4�����#�m��V¸�s�ԍh��b�h���zmUT�j֫dh�)!h ��U
�V���:4� �ѶKD�Z	Bۛ��R�H���G��:�����"��0z-��8��%�V��<�g�"Ĝ�̬�e�ӆf8d�j@����F�8����w�*��=�b��3ж���k\�xKr!���u�n:Nvn־�y!^�1=.4����%�6�f�D��2��:��;�R��tSU�\��d�;gy,�n#��]�a���bS�䧊� 0/��v�ؖs�-�r, �=��\���%'�ȉ�{٥��mµG�2<��߳�g?C����A�ϐ�;�@�������4������m�z�E�b�)��"N�C���[j�<���5�z�M��fx3Z��nDz2���Y��������X�v��U�"�Jd�\���z���~T�;^"�cUU{�Y���Ǳ��d�i�P�/^C��GQ׻V��MX���27�Õ�����J��+ѷ�X�91��\N:���ȇeIбژ�R2�e�!V��}��~O4�[��{C�w�ߪ/f�����SrY�@���f����^�+��mn@�ꔍ4��ie��0���A��;�qI��1�Ä��w3��\�g�Y$k.¯(�h؍pHY�玶�v�.�����S�^;�Hg�r��NFQ��S������H�D�h��Ϯ�g$��W^Sk����w!���	ۍj�w9�<�<��>������r��m�3�,��a�*$[xzv��5��`��:T�d������lLt����u�캝���Y�$�m0��s��b��3�{�R��)�����Q�<Vu&n�e܃�6��݇�#�j$�r E�C�� .�h9Ϧz.u3��]��mz˧NY˂�mHPb�m��[Ҹ�QC0��a,��Z�����	�/�8#���.'�hr��%�b���ڢ �`�/+�h�A�����\c�Q�O��IJ�7sDR��=a�)W����niv�,4�pDW���~\r̙�i4�0�۲��*q���o�mp��?=a��婼͊������ݢ�-ߺ�g�6&oZ�R����Y�QAL%r�և)JYj��E(X���I���llOJ-?q;?}��{s�sA0U�ܫx��zA�}��͊��>����jmӺj�M��h�A������c"
��'�����K|�@�Q��J�q#�&�+���>Z����&k��]N��8c�1c��4�o���c�K�Q�wG���řX�a���5k�Wc����û�6!��z��b��$T^�<ֶ�`����F��E�e��=��Å厢~=�_�x�i��	�������om�=��j��o7��;9x�l��%���j�T��N��7���f�m2%5���l�����Q�{z�p�t'z�0������'
D�;#����c�&J����ϔ�x��']��rk��H�hD�5@j������d���;��E����+<+.0(��u��8ϩ;_G0K��*&,V>�։i4ɣl���>���lP���R�ʎ���W�9�����i�f���Sݿ��}�xF^��h�#7hF�ƈ�zc3g���}����{;�Ȼ����- '���B"++�ɧfE��ʅjh�Wdc,t+��n��}����YW�h���v��K��O�4�"�����4#z��(DZw���+f`�ڇe4;5nEr���g����c��dG�b���`	o6���P�U��s�z���Ъ��٥�l�u�pc�w$9�Q���++�����OZ��U;x��X�-<�������[�^5@d��%�PuR��^5PJ/�����#&�6��UAOk�0�%xzTܽ]����� �H `uE��'1Of5W@&���C$tݧ)��
5MeixٛU��L�Vd��y%H'��2Y]kę��~ҝ�՛�CΦ��d|y�u{� /�YB�!�'�r��TS!)���z���ìf��Mħ�{�*H����T�oULB����:�Tג�;c��**�����Q��f1��4���f�XA���Kt���LhDg���J�1��,y��G_g�[O�{�0��y��D°d�aMs�'vs��1@%��/���>8��	ό'r@�� ���jHԕ7d�Dc�Y2�n�䐠�t���Y�a��%�(1��*��RN�Vμ�u�czBU3�MMd3IO^����0�B��ֽǏĠ�t��z����cbcӤU)t���s�d�ػ3��8a��#jp��E�����8@��G[.WO�	?wf��ψ�V��S��'�7�{`ᦘKd �p� �D��?��i��[�z�&5�N[02I�24�7�D�'v>"����we���?�v����j�]�R�-�\Ze�)�qN���L��O���j���>�y��E#)�/���3)�`+�;qG��٨�����8��k��ScN��ci��~6\׫���/|{�a�GYx.Q��|����UFN1.��5d%2��>ۻ���\ߟ� +t(P���a�pa!�P�x�mF�g���1�(��v���xMc�$.�$4bю�N�ƺ��J�9t��NPB�NT�j˧�Aݹ�5��ǲ��=T+��_U���ZoZ��}J2�	�@        �9%��7����<w�=�Ӯ&�U|,q�GL�7:�ǋ�T��nV��)1K��TA
W��$��Ul������Zj�GukR&宻%�T�1 �ʊ��Y+��ɧ&��g��%�S,��_;�I2dm�5 ���]r���,d��TU�p�b��Q=�5d�ӑby-�82�K☢�A;���Hep�v����͵�N0��j�# ��;D�j�8�~.Z�̸�o>�����jH�9��يj�'I�U�Plv�O��;0�lcKL�/�v���g3���x�5���鵗dt�5���O-Cj�]��E8X𞏺6ȿ�qC���
�[���"�S��ˆg������vM�x�UT�6��naRb����5�]�(h��"/�4J�=ۡ����x���B-�U�g!�+8�x�ky�(sM�f���D�tZ�#��w�qm��
Z�ĩ���L%�xO�&hΉ;x��^O���;=�ykƌ�d=���RU����R#Y����౥$�dKU��.���2��[�n�옸c��ݾ}֞����M/!nR�R����Vg���9SqP�0/�̤y/�Z3�{��m��T>��8 �d&�y���]ݯ&+)j�lR��YDh�*�S�dc+b�����R%(��y����e%,\���a8��/��3�݅ޙzxo�B�o˗Ɠ�9I��n�f��r��l���p.ED����,b�':ꋸ�9��-L.h�zz�}n&6Ruki{�"~Պ�m_	1C�H�VT�No�l
�UWT@EL����$�Q,�FA�Mk�Ą`4�P�P1�H*b�F��ސrf�O��jyݞ=�K-��K\�j�O%�38d����x������'�����Z�A哕���3�$���S�MMF�%S�Rw/�]�r���U#"y ��_�y�9��;��1�\^��<R��2�@�����N>U���l�J����25?�
	j��[�yMK���T-��܃����ǝ�U�]�K�$�|�ݔ��h��y�¥0�Z��|�M�cZ��y��|;���:yh��HF�q�.+���=tWQT/T/x"(��Q=�4�Ep�=�^5K�v"��t�ɀ^�N#HQ���e8����*��gq׳Ү��"�s���k1>IG`WJ݇"��,B��X�en���@�qB4����b�?��h��	��0��Y4N=�@� [�_;1���3Ħ{b���2�_��&�9ȗ ��T:�i5��r�Z��TKT�9�Y?@7$�3W�]*�(i��,��n���d aeOG>�4�~/x�`,?<���I�kQ�49���0m-u�m~� yB#����>V���ZӷD6F:r˃�(:j�77�m+#E6ھ�s��N�-k�''(���P��
��:�2��w��H/w��7�k�J��x�:���`�� V��cV7���"�]E]���Jn�����&��W��p�9��� �7�]���j�U��p�(�Վ,&t�[�y�|��/�!�t�;�]���kn�.��f◥W��t�D���J�)�
�p=�4e2�MRak㴡2�u��7x��(�b��2��m:�Z��]:҇!x{RB�Շ�:�V�t��u���v80�-�X�-sv��
�3ln�7��I�c"�D^Mح��j��+�|V)�se�}%�]�l�	�*�=�STF��o�H�vhY.'Ywm�X���������n�Jn���çP�;/��V;�v��轝.�ب�
��a�=u�r�$oZ�3"�g)P�σ�[H)�K�w���|޾��%�^,:-\�Gf�"��̀�-ؐ|n����b�|y��}�#c{�6��C]#���-�҅�D�zVf�8.����Y���H糊�A�T\ӵ��i�Xq+a�OȮ��M��2����AM��ݨ����f���J��n
�77ѐ»H�2R86�a��b6d�s�]c��Qh�����;���/R�0	(t'�Uq>,��,��-I�#L̇cH�ذ�6��\��\+B��M<��k����A�l�HZ�U//b����i{D��Ϥ�]`�;6�B��JT���+��V��#�SL��.�%��A��*)�I�)_F.�r�\xwhӚ����J;uf����e�9
Kr���6ݳm[�+Q�y��r���)��������m���&G�<��Z9�θ�,ʇ.�1��侕}����[
�ws�a��늬�=s�B�2��
�ˡ�U�4�9iw:��Z����,V٭`VR5���W�;/�Y�˰X��l���Nf�`�(�opn;�ͺbRw�w����v�*;��v�k��{�8>i0���9��r14�hh�*{�xy�{m˘;e�v��L��\[vZ酂%�u�8N�:tX�}6�n�Œ'��x�r-�q����v���9�)�!�MCa���	Ӗ��˞~� 5@�#��� (Vϛ��]kf�qz1
��q_}�%�LȘ����#9(�¡dk�7&@��U������=����xriO�R���d5ґ{��_@���3���5�|��m��4<bbV��U)�ˤ�cz�le��ט;�*���3�YU|<�^|�՗��2^:���c��ɢ��H2���Ɯb�g�mۼJ����h0��2�0b��&������9��2�0o=̆�3���^7�
�k��l&�$�骝��r�|w��l84ܾ�����&Ӷ�{c-�4��� !٧���p�u39��¯���`�Q������Omr�TU�i�OeWj��w��RA��m���'N�z캱�T��wta�΢g`��1,V7�E;7��C���9�r�W��뷽Y��֔�����L�W��:��Ơ�F����Ɲ�M�<�E���?�wG�����j�oF�����y֞ǘ8�Or;�	;{!�Za���9\�`E:��PDi������.f�R����h������P9��cg���޶��a���l��r)�HxC�;^ֺ��[��y��ʭ��Q�8�(m�ۗ�}��d����սI*�na���~������r��#U��>k�<�������B�rr\.얪��[iE(��86X��p�QHG����aA9:c��a�&Bs�T%���9�8O��4N�c�w#��M��yN�m�����cNo4����9��]W��Ʀ)�'z����N��P+���V[B�i? P�{�����r��PЕiS$L]�5�:{3O@z����~�L����i�!�%y�����i��^^��N�Y^�݆�1MM��u�5�?U5��n�yo, Ufc�lƤ1�V��*q%���դ�[�\�;�"�8�7�^�i�?E�~��7��ɮ�S	�����ފ���%���E���m��k��oNuO�<�z_5�{n"R�*Lu�E�{�Qp�ܜ2w	�G&�K]I��~��*�����Ӯw�ڥ���u��'�W&]�j6����Q�y�-O�� <D4T�OV���aZ����Ю�Y�me���@j.��8�K�u��˳璱p��&��� ��uǤ����Kn녒��         �,�ە�
��`�z	Ys'ՙ]Yz�F��������!�ӊ�bP�|�	�{m�
�r�����F��1Ě[ep%t٬�d�I�u���Ӳ�D�W�S��� D���N�i�H�U�mb��D]�g�A[ۋ;&i�������w�'��&R��X�ݣǒ�u[�Ȉ襮��@/K���T�+�!��+2j�V�2;��! �27���j���_���qg�?lst��|!��!����ĭ�'�}�1T�����mG�{�#ǧ1�`�EE�>1ͤA�h����b����*i�<�X���܈\IV�gB��뤜�ל[ �Z�i�\��c����gwt׭<�B�8�X{>?|>����UH�_B�M����P�49>����:(�G*��$4�f��4�o=�r
���Y��W�1���C2��qa��wڜ�`Ν15��_��<[�N
��*���K[1ב9�����憧������ �R�;
��c��'1���p�^O��WRu��T��GD���*�8c������� ��B;R�(��[A�-�OJ����qT7t��_/�]��a��W���Y9h�W���cڃE��q�pi�
A�nѷ$�q������'�,b��n�I��^e�Mx��<1����gK�A{���h�����J)O��\��ե�ƹ�'�|M�R�Xd�X�XR��� �7D�>V2�ã6�6��a��/3'��Kn��ƪ�v�q]���gg'@�Hw�S4	M�CR�PWZl�M5��ղ4��곞�Y�nڧ)D��E
ز��U���ގ�a+��y߄��d�����ξ��,��cy��(n�.���3���y��n��b	!��nd=��yG𶞥s)�1n�=/#��ｐ�5��YQ��t���,�f9D01��\b:+��ل���n�����S�5{��d�_bJ�����Y��fd�~#��j��O����|�17�$Od��p�̬�'l�İ)n �����O����䳾H��c,w��(]5�-e:�1�B�=w�|՜��z��,A$�=5�!�5e�gnx�??��&�+�d���1~yf�d��G
����H���"��@gwd����ᯬ\�mlHw��;S�vms�L�a<��L=�ƾ�\΃y�.���3��V('�;o�_2HӃ�o��$z|OԸE�HY���n��}��d(�m��;5��rˢ	�k�ի�t�߽%:���t�ю�� �̖ �</M��Q-D�ڨ������2�!�h�zt����o<M5]�fj[�4�(L׹y��ɫe^M�#;��o�6�-�J�$֗R� ��B�!S(�x��N�r�=�gb�O�|;	He��Nn��G�)ߨ�s�c�i
!y�х�|���=��D�@A��ۣ�^�k̻�������w{ÛL�m��)��*]�a�B�5,��cِ���[f]��ܼ���k�5\�|��� �������	��:@ �԰At�,�O
�n5qsӧp�l1�.�Pf�!TJ���ݝ��<P�;�>=�z�D�r~ '�m���V�k![�m�X�E!�V��+ L�DB(l${A`��^r���uG�t�ٗ�T�)���U�F�EL1��AI^��o��zN�H���xolw���n];�50n�E�]��B�Kg�Z���}Їs�u�J���s;s_���\�46��d��c{�U�����}}�ƿ��pl�SJg?ge!�muSHi�b��"�Lt�7� N�z��̎���"�'���{#s�\�䜲LJ�N���u<�7=�nuV�z�io+���u���=�'.�57=t�sa�no{�>x	���
��(@y�ڐْ*�	��b��u��ԝ�8Tub_"2�d��^}�XT  ���IMQ4Xn-�]S�w��}��c�]��ú�$☒]�T���=S�-W�
�e�@�����䕊f[nR�OE
�~��)��b�!����qO��v�0��q�Tc�T��sd�2��D�g/&+�Y�du�ԱSBb�ƭʲ�tZ)U��JԳ��>��	�]�;g"\�%@|:x�it(�U˜��A��,�#¡�"	V+fEe?[#2�G�|����`Ԡ.� �T�٘�����#$��i��a�Э��__���7�S�q�TC�r��V�N
��Y�D�,GF�4II�z|ԫw�6�YML��sT�n�h�d�;����˾�q�=,2p}=v{7~̩e={�߰��BYBO/�}*�8w���{�>Um�����<Z�S��gXej%K���q�9�Y�t�Q�뎶��UV;yK�dړ����_�(^�D�FN��Ḟ�Oǧ���~�0�<6��% �w[�9�[�0�g:,EI�t_{9U5յ��n�#�0�3��Q�C�z4�h�'t;�㓦F,����7;y�/�|��5�A	P Řm��d�0rPp�        `���1ѓg�o���̲A��Qmz���ylQ��K�2�i��VMa��4ʻ���30@����XH�(�,"&�N��jx�2�G�^��{���=9�(�L�6���cP�S�}�dR�����G�*&��j!#p� u[��nX��*2�Z`��f�I^K��uӒX�ٷ�%��t>�R롱���B�S��8�z�1-=����ox	�ϒ׼@L�Ɯ�6�X�kdx�����w-�	�wP�0*��q=��FȆ�l��S��v�=n�H��w�T���	��!���_O�X�l�� @��η,EJvϽ���?{#xJ�%F��qe�Ѭ�a.E�t\WA����	�{�t/�۰-�+uQ�	�:���[6�����ˣa�(13�d!�*ۢV׋���*�k��T׷[!PZO+p!���	`��zD�@f~�=ڟw27�r��=W�uIR�%š�j��l��R/%�����|��;�6;c�h2,�s��Oi6x0��y�_�C��ܱB�����	u�sr�ݤUY[�۶=W�U�YJ�h�g>���`'4�(V�(�(ɖ[f���}������Yҕ��h��	�I�������.`KF�AJ�:�Խ�n}h�;݇A��Fg7?V�&G�˴��'�zvL�p�hbvɻ�GB$`5E:N�v�qYxZ�׷���:�z�ڶ�n弬!j,;^��Ts�%�wPƐ���`�Hg�k�������HD86�n�C~��I"2(�W>!�{��T��XNkv,b�������7�b�^ ~*��;%���{���nL�y2D�OB;P�#�i����$�I�w��=v2g:*û���4�HxĔjf��١���nh3��{P=2����A����bN�����Fk�+��vi�<��> l��Tn<u6���⤽Ơ�}�fU�ͺ�w<�� _7'����������K[�V۶78��m��d�t�V)����m3NX�؅X��@��kH��i~Ō#���kc�Za��@M��Sչo/,��� 1VAy�$Ce*�9]gγ�����2[�B,�d3��6�4\�{�}�Y���g��a2N��^�xt&�Q��9Ki��[��i�]�����������8
�N�Kͮ��vv�~�ޜ0�-nzᨋ�a��/Y׍��Ϡ6��$i�9�o��G`�Xb�c�&:��30�|2�9���4�#i�����|K���l�x�yx�`�q����Y�t%��] cȎۮl�xyV  ��J�&s �>��V����,p��&]CRgn/�X�c���x0�Ƌw��Wy��wk�&tGi�y��y��W<�.��Ӱ9���<��FZ��	Ժp�Cu�͸������9��:�Փ���5�d��K$����#��W\���~oP{�c�gj{d��u���=��f���݀T8��694Y=��YW���&�U��d��; V7%t#?<+��k��0	�=������DBnp�'��3/�͉���l��͹�c����@P�oDQ�����r~Ĳtj6?0��B����3�=�j�ր�L��\�g�߫6�m�G��E<���xb�ڱ�_M��:�Q�d��OB3'�s���3�c��$�h�2�$�s�Neޘ,T�9b�nd'��Ӧ0nr�7r�0ݴ-���3�(�~�T Nn�X0^7[=�K�J�c�uN��2�E��ʇ�Xu�%��se��]�
��x8��o���M`�Y��L�yb�`5A��M �S S! j�e���c��b��%�軙]QُDdԽ�C(���e�!A�j;�.u���mJ������8�&g�G���S��G��}wBX���0ԍ�;H�j��/�cxQ�*C뉸ȵsM�4;��/��\^��gh �p�1I§�ˈz��땊�c4D�f��Դ������%��d��{��W�=y�����Ǥ�][];*O4@Z��/ ^�� �}OѦp��u�9�ý4uy�r�\����	yO�o�j}Y�вA��f�FWD�9��u�xg�C�xŭ;x�B�}5�G[e��c�w1�oC΅nB�ϊ,�u��K��ƒc�@�n���/�AZ[JTa�ly��H��dðhaZB�݃�R��lu�7�"B���]���'��͜�b��]g+Վ���S<��t���G�K� ^� \�|��@���
w.��D���z�wS��
IG�BsA���}���W�v�3��׳i��O�B�L4�BHȲ�D]�;��Ǔ���n�L�j�x��-�H��#�Hq��̛�8n�'��z��7����)v=mY�`�{���65�6ugY���P��^^�ǆ��!�&�mB��p��]ᷯ��Y��j�f���s7�Ժn�-�+�6
���q(����@��*˳|�Z�sF��&��^�kv�V�Y��N�����m����Oar�6�u����N�����!���7�b��ӶH�\8��.�y���,ڐ��`�?]1?��I��G���Y}�����wٰ�;$N��u�6u���qdPfi�H�D˷L7�z�Ûtjk�J�Ds{������V3�X޷9��V�\aX�I��J�D-V��4��@�ĺ<��P�M�7�fZ��k�]�o�]�m�װ��Ҵ��B9���r\�L�L�嗒���q���:`+oN�Mt�x��
!h$�kE�2�х`�2sl���6��`�m��z$�F�M#ʹ	҉4H&��5qX�Y%7|m}�k6�s�m��宭��][���n0u�F�gC7��fƴ�+1���(�3��VWQR&���݆��rm�q����Y UD���N�e�48ۻ�P�5U�Uٻ���D�#\g�E����ګ/�XM�����аP��Zv�/o�Ĉ�0i�K�9���lufv9mlG�3�~O������� 	%�	$l�Wl�$�R�Iij�B@���                                                  �X2GH�s�f�^�9�vAWT���2H�籃����bͳ��$�L���K����$:Z;�Lk����[8t����R��	��T��:I�̙ڟ=���&�ث��Y5[�R���	���,:��)���twݜ�Y��"!]�"�0;�*M�W\m�^��G��7��6���kA�S6Zn��5f�7`nv�m�$wVk�kG��_5�4�l]�٪��W{�'R�{�;ų:���j��
����T6١�ɹ��6,L\�nF�YA'|y�WY�{a�1#6�A��T��X�jwDEh�Sl&���J3)��L���U�Yk��heɁ�I�M�m�l8Ia7tn��H��a$~�4c,Ds�o2mV�ȱ���n\J��V�FW4���X�.��]�ԒǱɦW�4I�.YZ�0X�f �{�i���g�SW��ݣܱd�U�K#���"{6�M�m)��X%��岇& s��p�!FF�ȮNͺ;7=��N3[�Q��M1Tʘ�j��ɔp3�\���� �q�F��7����@턑#B�,�AF@;�防�eOWA�[�1�r��NW�V�0�v5��uJH0��M9�gl��[�"���(��;����.�}.8��6�m��V�E�½�SR>`��2����BE�l14Y$�I#�T�~�M�(� Ed��}1��#	�����K�3��mk�D�oM�Җ�D7n�pk&9.�U>�U�L�{���4%��ƙ��["��2�0��A0�k��cS3/n&��dU�h�ti����q�ۻ���	3`�=��������Rљm�ܵM�N�vI/6c���W��^�R5�e�f�1��
'�cN�+@��R�T+u
I�]�+(�HH�D�%�6�r��hE%�

U�Q��[�]��zc��B��Q�ZWa@��         �s���Y�W
���e�|�����M��w��EU�[�*�evu˚jc�TK��#R���D�W*H�1�UE����P�&��9*�n��m[d��xǙ,�v��yIn�7@Y�
����˷+x���@Q����Nр�m�]sr�"�"o1����c���L�,�n(@J�si�eP�6"0rV'X�UxYrdtSr��MJ���1�a���ͭ��*�ǜ��A�W'���8�ջ֗�L��.�їWф@x1��ƅ�w�X\��;�L�.r:Ї���r�f#8r�YB�_π��h��r�4j�ݛ�S�	�Z� ��UH ~�؃��2%D�w{��pX���kOA�
��疘���w�-�����Z��1�:b��0B+�Jؚ�6������S �����o�!�^�g�ê�~ɐ�@��s�j�C��=�{	o}r&1�	�\k��F�=�l�_�px{��6\@Z7��͎�¤��e�A�� �ڙ��v�=�~-=�i�:�晚����u�j��&_�wy2�&J�+7eQP��	m�����n�!F��7w'��ɡic!g8��N�2��2�6ܝl�"k.3��Qe�l±$s!���;���}��=EL]0՗s�_��o֭��=�g�=��R�	��!���t��A�����u���ɑ=���\} ���0+�д�� ��'���n�fnl����i�٠�v;{n��O��0k8���1���3�
�%Um�ޑYX��'�I5i��q�6_+�����N�6;�F�츂50i��2N	����(u�>��P�Q+j��(���t�K�q�c�2�ΊoS[܈[&���
r-�ِ�Y$��"���5FL\�����*vs�`l>P,��$�<�fo�ғUFឃ�#p2 gb���j���Y;Lᘳ���"2;!��!�H!gZ�f��e�b����o�q2�_L�u���ڽ��^��#���K�i^�}��ݑ��rIBz�e����e�`jZ.\Œ�+��Q
̨�`��@�|έ��j^X��l�N�'=gg�#P�	�n�P^�O=�0:����i�^�1��V\e�%���ib�Ӷl��HqD�|�E��*��1ZD��e��Ŀgׄzg�+)I�*�w��xM#�yU*���K���^C�w�o���V���5�^���kR�2dķ�J;����̩�O1H?�6�E��v�K�"��Rwzp�H73��RՀZ�1�i��wVF��$n6[T�&�ERi��Gg{�^��]	ַHU���כ/�}"��<�5�Ņf����!;���6¥�YS�q]챋pZ=Ci���؀�H�,��k�)/��314V�ϵ��N.�@��2\c��5~���#X}e�lFӐ\!��}�:Q)�_.��5`���w�M̀�%�l�]d=��JM�
�w&��U�sb]Éݫ��e*]��9�~���&�ySTMJ�p� �^�Ӌ��c�,�׿�����^[�����!�%�|g�3�D(�鞲Y?nMƬ�t=)��(3h��AƑ͏���Ç��ܪ�l�5�S\Cc竳�8�v��/
x��S�������ѡFk
���}����"��*���M3\��a��ue�&O��@�%�XQj�dH%n�`��Q2J�}��)홥��n��o7�� v���zk��D�j�c����ަ�]��7v�'(����J3*8z���]yΆ�cBv�3��С�z��H2��jvW���F�	�8ˉ_�cE;F��v���R��&�"�%$�U@RF�G/y��ޞi��w��δ�fZTA��au忥��I�ޟ#c���'$�J�@k�~����!R{&4�s1|� �W�����ێ�^�j�ȁ#�����{���[�F�~�ȟ@6O`	���$�تɊ���hj���p`�LUJ=B���$D��>��tis�2lm��i��t;�|�}:"�}�(�r3�� �����iةw��	��J{�|Kc,�pȸg!���"�n��^�~�O2r-�_2S�y��k�mv�t��޲vه=?^����x5r��-�q���{L6b��0|4��$k�!��k����<�����K�yϱ�'��sxd��Z�͔L��M]L(d�i޻0�3�[;�%���B_2�_{��f��3�B�zgh��h�P�	td�1��q��rs!���y�\��m�8�ܽ�q�B� ����ߣ�:������f��R{˞aH��m�q�;���u�f�o��dK���O;Q=-nӹUIŋ�uk\ J"�t3�k�ْ�	��$�.OGn�i�5K��Cj�U�kZҺi7�Q�svG�V��         D]��YrnLs�ה���$R���ȄL1�f���F`�m6)�W���S&\X�r�d�9#�x��M�U[��M���#���Ei��X�Ђ�G��C�vkm��4(�dMU$t-M�Z��%h+j�Rvu�̭'�u�(�q�%�V*�U�(�h�2�6�v����GUP��
��`��|C�'׊����* �	�n��6g-&S���kkJF�K���_�T�+�n�����.�G�V��Y�,4��n����M(��F6�"|"����z��"�=�uH(,Qը���g#��ɫa�d�6v/�䓳h70��1�68u=m�	+�,������+�iQ�j|�HӢ�v/��ops�Q�cJvI�d�&qB��!�lm;�6�)��n�9P��L�	ۺo������d���}\h��x��2������WX�EC�L{{�x)I�Y��|�5 ��6��$�\�5����ˇԽ8�yv�\�,0���.u��vs�y��ܝ �;󕧛*eN6[�J�#�4ꐱ2��%�I���g=ah��1��`�D9���#��Ӿ(~�P+�w.��F���1���!�F�,874cݵ�Q���ںx$uJ�"��P�(P���3q��-צk8�"�r޳�l})���x�%�z��cW
�
<�Yc��X�`P#ZNl(B)��9����aY��q�`��W)cP������BPZg�3���W�]��3��K�?�|w&��QhU�"���~~E��*a3Cܽ����}������ȣ��o0��~��w�f�Mw~p������]ٹ����/�:�k͘�UP>͕Mp�Q�U��gcA����+��)��C	�3ύ ��~oK�^7����Go.W��ǶsږCi�X��'�3�L)-�,�%�e��b�jh�;�[�˜��m�5~ή���<�ȡ!�B�0��P�/�C6ʗ4Nۻ����>�sZ]���Ʉ��W-�*q"D�-��M��&+j����2�F���+���3��Y���Tǈ�A�b�[V~\jw��ڰ����˼E���ad�dtt��5
<LDK4n<�	d�r�T�b���p��]�mj!�W0�nx�yb�{�z�����w#@���xss�<j��._h�9���Z�<���s�XJBLG>�ѝ��A�rS�mH�p0�9�!��񇳿<�5��c��U��C��X/�S��{g���{@�$$
KQ�u���L�c��3�s�|����S�`N�1�Z6�<�u{�+���>�!��o��8��m�uO�W��Ϥ�N`��z��,��ԙ��]
��y�sLj�ǣnո���`<Û�a���g��f\1C��tOi�,����l�uI���p�a�'	Że}��y�ԛ��툭2]4��O;m�>` oýu>��[6�M���]}���Ii��L�t�H�4���6`m�-�cYטm��T�������rZj^���" ��>�F܋���=惂h�C��_e@�3��Ǐ=�5�kٻ�z!�'dd3�?-<��&�ͩ��JZ��	hd���.�sŊ���i6���[�֝�V�ů�"=�
��.^��tG��Y5��3��c��]�fs�9�4-"I���3B�F �{w]��g���%�����QFܴ�Έ����G׍�XPD�[<�4)��*o{]ORKa��S(��OMLx�F�{��xoؤ?-��<��N�;��v��_����.i�u�Z뱦���X�c"�WYpE]�2�@I�0f ���+�^B�S����7u��[���L��K5EWyҮ�c�dRY����+(Ǝ0SjCkV}��@?_���k��٦�iЏFwL̼�6f��dW� L`度��Aw6�sT�������2 �nۮ'"�Ҳ�hPtz�tTV��A�Ɯ��h���H7�v`=��C�0�1.� T�-����m.t�;�MK��S7)t�*�b������Y�ʼ�1����B�`PL��(V�=qL�x6�w�wP��Q�� MԀg�����<�0j�]$4��@�x����������5�0��G�v��A�t��*�pHj��%���&�0űA�D��{d� ������{��s��İG_�_A�ͼ�Q��f���n���A��,��;Z�KK����s3��	χϑJ���>�=ѵ�Yܟf�W١��.T�Ŕ��3��E��Z_7�#9�-�j��K��`��4���W�ɋ"��(�����n����
�l40�gI���u��-���Sֽ��P�~aT��}B�a��t����ܑ@�B4EIUSkM�knr݀@%!lN�         K$%*2���Hgt��T�X����O��uҐ��O.�����H�$D���.�1��iB�N9}V�`�YkQP���YS�d�ݮ�.�-{1$�ˍ����c�cV���&3�ksm��E(�V#�cݭm�Kq��n��QK+��Fi�rP`8�dL�v��j 㕎�̘��ẞH4J�Mn�%�ng!-�m��3���pJ�W8����g���N�������4��f���s���� d�
*V�ݥ�c�ȩ	2�P���FZ2�LV.砹݊��:��Q"v����/y�a�y�W��On˅�#[�.�����'��1��P�̯9�pҎG�t�ݍ�Ԑ�n4,��U����?:�J��,�'鶈L� d����e�t�B��WW$m�a�H�sb�qT�׼��&�q��"j&�a��x�~ԡ�{de�����bzlb3n���RO�����Q��0�#�#R�8��tG��;
��4or���հ6���TX�Fd�����X=�cäJ9��%�@r�f��
f���+m��U��-�f�<!k��p�V[hW%R�BG���ty,O#�������9 ��2�ͱ�����#��ܻquOk��=�=�c��4�
�ij8���F^Ff��b`li��gn�<�a��Dq��靣Ѭä�0��G�}�'C�Gv"h�K�9-�ϊ��w�c�zb޼2��ڑ*Kc�B���ݪ�O�͂^���_l��^.�Xq�ص����4��{�����{�^���bP����Zb�fO�'a5[J�I�������������"_�#�z��g!9�-J�7v_�M'އ5������e�8��,��@5'�����9o"C�xz��_t�Α��ģ��e��/l��lI����� ��E��6�us'�v���@��kñ�o����W�^;�>��.�^�d�	�̜�g;���q
�V���c�R��3���M��C0v-���mh��^l��i�n��l�b����^t�Tr/�Wn E,��<Vj��VQ
�\�C����Lm%w��5�����s[7��B>/v`<�ں��ڎs�▭>{��M똞e�Zu�]Bq�
�0uz� �U�ܲ�nKIt�&����R5ϧ;�R꤇�n�<UM���O�7��.�$�}��dj��C���;��.}w���@,R$��C�����/g��i��g��1��'f�ױ�b��G�!�S+|}S/2M[��0A/��N,��i�M���5�t-�h���3�O�	ɛC�go(����ݵ��B_d�#n�*�0�7,�:лl��.�Y�ܬ	e򝼯X�f��M��(�sQ&��7�vB#��r�B�
0#JA���@m�mY��H�#�M��J�8Usto���6�[�1��7X)<�ڠ�xw�;ًg��v�;������0��,8�G:XI���օ1�яQ��C�lj^gJ�U�ļ�����l�ަ�a��j�5$��}N�v��@�oi�>,��q��ʏe']�u�^�s%��s�1�/o(��3���{��R
޶!��l�*�z��%A^T�R�+�X��q:�i<���C�	��}�֮��fn��>v�!�:T�f��Zۺύr�9��/'Z�&���Zڗ�*�u�g�9�f���+��gl��n�>-��$ѩ�F�V^�7�Z���A����7�F�|�o�
5�S��Ŋ{V�j>���� ���Csj&�m께(�	$r$.�A(�`(6ʝ����K�]�d��w���ͯ{����xNf��1���Ȳ�镛\�{�af��t�k�Y#w�p����՜���{���b�T���ҜF���7{�Axs�u�a�gO/PyTD��őHX ��1��8�jBb�(B0)��.ś�IA�m�8�]�9��̇1��PU����Á+�8e�Mp�Gl[��wWBv���K�V�B�"��v@'t����d��@���G�9���k�~7o�r����7vѲ��v����{�s-�[,�R��B��G�ngP�a.�nDzs����ElѸ��X�m����,�=s�FuE r_e����2��W}�kM�"z��:d7�*.5�s��e]5��������V��D����ǃtV�)��λ5��0����	JU/�;*��QguΫ)p��o]�
]�6��ٙ�P��Ύޚ4�m����0�|\�UٲF�<����͆���t����S/�F�j���{v&�n�W# �@d�����7чwr��y�N�vS�d�3�+a��"5�}=ewCj��!��_H���� ��0%
��h�oe��_`]�JJ�B��+�Zǜ�Ҝ�rY�U���R��%y�	�7u�5�%+8(l3GC�AN��PC��ťJ�Mc�s����+����g�Ģ�"���kd���O����`��ϼ]?�v࠷����Ų���sM�\��j4Ya<�p+���rL�y�X�o��L��l_<8�y��O	������N-��N����k���<��FP���:y�'�;���$��̅\Ce[<�F����[�qL5�O4�c�|-<S`PG�(i�;~]�-�t����y��ݢi����q��~�SY�?�V�����-T�ڼ�~��GQ��WTle/5Ӻ����S�T0���ަ��Om�P���Y/n�*��qE�å6�D~��YX�<���ל����~F�i�SQ�O[�Eq�N��(x50�t*�g�k�Q1��Q�QV�dhm�q��W{�+�K�V�J���AQ!V1d�!n�w{��o�wxz�uw�˂*yi�����"v��*7/�5����P1o�0�9�
{��R�R���=J+3���~�b��k�7\÷r�y`#��90�q(��^���9��@����B	rە8���i�՘ꈠ�f���A���Ŷ��]��7��3���<-E��^n�'��랿I�0u��є�P뗱m��	U�z82q���|�	�C�O�^�@tm����nd`W�V6����oͭ���x�¾��-��*f*�C
mG��
h���(,�xb���ǧ�G�8�
�^��H�	D�i���zh��7J���c/���2�pe
�s�4��Z�q��t\�������Z�"J������3���<�]&�������x+D���aS�pɝ�9��?8h�zf[qw�R����p�Ӥ��tE���ީ--J���4iw$��������E0�Sn�q��76��8�Ϝa���O�����d�0�j�Ut7�J!s(U�����Cr��5x,�Oú;��3y\Ҫ� ���t����zvUroxWGkNI@        U�\���μ�r�d�qg_r=�ܙ�Ww1���*�-Mch�6�!��U��j�)-j7鉶ő�tլ����e$��i�]Zd@I(ʅ"CDFI�JGSн!��%��%9�feOD�ۖ'ǽ�n`�I�H��V�V]�Q�l �;e �!W2E�H�lJX��� ��J\�$��o^+�)&M�CE0G��ei���'˚�d�- ,h��l3�w��w�S�2����TQ��*}~�Й3����d�2ɒF]�n�˞�n�|����e�δ���C<2 A9�w�2�[��mw��8tt��Kk�lf�.:��[�4�>(�\���t�b�t`dl8<أ�\M�}��7Y(��`��q���N(��@�.9|Gd{�����Lϝ=�� i�LQ/��5/��Œڋ����R��Y��z���c*�j3K��� �1l�����y�}t�����l���d<�8r]�\��bL�G�/!���[0Z�Ls3���9�-�\n=�4��¢+��cP���L��A��Ã؈7�]���^�ق� �,D�9C����[�����hn�	�����ތ�Ӊ��-�܁����A{�6���5셀>^2���G�C�r�(X0���72���J�p��bc�]��徙\�W65s͠S-~P��54*S�הmM��uXĻmˎ^^�gs6��w���(� t�L�@1�c`��h(��W[O6�b_T�Ac&���p��2q�`d�U�3gD�;��c\^���OiW���L���;�ϊʡ3�/E��C�vH%� bZbЈD����z���]5'��oËD�^�p_^lp��Df� p4񒣡�pb�G��K�Br�I� 7�ݻ�#:�*��x��N����/E����ǳ����q�u{*Y�1rXC��[5�B֕[YM��1+�u��� Ʋ���࿉P��>,�<L�2�t;8�6c��|�m����f.\fs�MOf��/�f*�L Q���_�̹yZT�X��� T���:"��m9U���V�BɄ�/�~�/��,^�U Ó�0��=��иj�/F���X���6�#���|l���}�nL�gp^�4���J���4G�.q�����;x]��I�I��]���=���T�r�Csv�!�p��w��`|���p\�u;�+���Lĕ���Ȅ���W�q�����8���ww��<��ze��ǩn�r�{g��u3�a"�!�H5Th����`����zέ�Y�A�h�ƃp��1a���<͞«�w���NW�s��7��n+2�za�(fz����c��K�ˌ���o~�-�I�c�>���laXx.D�훆w�e~_]�=�2ͦcy�"d���IwwJ5ܻ<F�q���鍭�s��DZ�j�oo�>�����<x�(�-g���sN��߼>�:5�nI!���mm�m�m1��$�����1�eB�Զ�R�n&{�Ǯr��o�����Pg$!�x�Qb��}���#{qB��o=�l�m@Ww=t�T �%��Qt��,�hT$L�'+9��z��nym�;�ŧ}%ZG���9��"��m�g\R�;zr�ȫ޸���G�R�˖�GVgэ�:���u�
��x�=G	�g�i�7BΛY-��E���3�_��6,bGq�!֞�d場��֦F*�bT�M�Ù�"/u�):,u0궡��[71��k}Gl�	I��c¨@͉��fH��vͥ`��԰�zvP9�F��d��385�S�r+�阩 `a"
�{�{�7}a�������=��$�"�2�e��L�ǻ�TJ�}{�;^�̗�")O� ������� h2���u#�z��־�uU�%NӞz�+'b-��8�r^q�c[e��L�r6�t�yi�a����09^1��{�YnD��qH�5����G) �������dJ�ᙁ*���+�T��V�XA� �o7�$V�8�kN[�4&J�hI���^p����\�P%�h�I����$�{�t��'1 ζu8��s(���k}y��ݽ  ��ff��(�e�w�Uw��Z�Z�hG�QD�9mZ���s�*��4���g����ZH��O����)/Lu�����j��*�vLn�?D��ںZ��B�uJ�Mgs��]ph!O��Zj��L Q�QU�ޯtt�m��J�k�q�Q��<���{f)f�ܡ��Ņ��⩅��e��'0vz4�ڧ @���Jt;�y9�'}�ܼ�w�֘�����3�&����gqG]?:� ��	��a�n<�Ċ�������Ź;ܢb��Cc��
�a�׻&=�Z�_[?]�ӽ��ݾY�L���o8D}�D�ES�� �t�kM�;5M(����+q䑖�        )G#����3���u ���e�0����꯯e�2wb��MI���SpV1�@C�Y�^�$\UM�w+U�;�<����l��x�r���/X�dQ]c�,�Ԋ�@��,�Q�$�KU�Ա�#�\�MFUSX�&�N����on��:��V�´en�����13(�2���W,�<�Ve�eR
�Q&�m�Y����[�)3�9���pB�z"����r��1�!w���ȹ1���=!�/�7ޙ��W&rgaa�x����%Й�r�P��~�ۈ~���H��y�I;�:�|k`�X�&o)U���N��L�@m��4:����5Ïxg����N����Y>]� 򖹧Υ���ŉ
�a�s����2h,y)�d���[==6a͠��6:{�,h��߀�&����	xj��XiaA�i��0Y��s%J/�ˈ����րL?��j.�s����L�{fa��1B�kw;3B	�j�Cmˁ�� ��K�F���l�Mi!��?�5P�p�*��Brx��5w�!�wk���kyj{p��u[&��IR#B�R�O�c���A����d#�QJ�٘�������'%�?J�i @_�>o���m_����Ih��I�m���;FЬz�:�VD`�zb��|���>��(�K�wx��u;�~S%�C����L��%��WL̡	�|��ѹR�t���|��;t�*ٺ�ڕ>�P,-���HI a�A���
�a�L�/{�+�$i���fE��$��B�y��z�N]y���>�)Xk0T�<��:[`!Zݵ.����L;�"m�B�8#�dn�l&Y:tS17�O�R-Е����Tc�/<}�Bڀ�@�sl��-���z����B��曦��:̻BK���V2y�O<�g���,biZĦ��ձ)�xM�����T��^���g/�Px�]��>��h��ysc*,˝
����[d-��	`J�{��j�����n۶���>��@�Y��|���DP٨�#�Jr���A�}4�5&��Oɳ7,�l	eo�X�ʢX�*E��Q�0x��UՕ�cmKk�hU�/�V�3�����.'�n嬉f�L�B����e	}�b2ovry�܀��	�����KE�X4/�;8�c��q���;��r/veV|o}��}y��zY7����븪<�4
�ɀx���*E
��{�Q���f]�`�i���b��4�td8��0��H��W���
�!��CT��)Jx{��L���/p�	J����:�ҥ���ҫ r��TV]F�������C4pe}�D[R��\W8*i\�ڞi�8L�����g����79���#�<K��dbV�S?�=��J<��脚@l�?;Xb f<�(��k���s�=�Y3����*�z%;�!�}Goz\�T�<ne��>�p��1���WK/�7͔b4���v�e���n�d���j��xQ��06�vFWg%&^0H�ځ82e�<�+�v���Xd3 =�4�\��-�`��n�4�Gk-$RKSWEeVq��!�$�![�{0-��{�d�����p�Ξ���`{�x��/M[)�i�4�
�_uPz���E5Bte�+�����|)B�{�'��Ol9l o0󉍑�nl��6L��^PqZ�(�nØ�!�E�����2j?X�=��܀�
C�98����ũc�os!^�2�����V�N���hǀ+��I���u�d�s�x:�p�,���t`�S��g\�ec6��v�o����%u-�xQMM=��X vc=�̝L�_T�(f`��+[]����^86�]�S�1Qz��k
�������q��:��w��"A�ۖ2�ALn��J-2Bl�AEܼyDw�C�z�9կ�MM&�9�u;�uu�����c�IȨtѮ�q�4ix.��vP	' �݅o��E�3�w�Y��D��	��{��!8�%�ˮ�ò�H����~��Ǵ���Z�V�!zA�Ż�w"���;4�(�i��+j)�2�)�@J �"{���˟No���#;H�����5�yƼ,��w�2���Vtǁ���R,WQ��)��`mعv(@�A�ăV�\�dn�Xt񇫅hm��3^6�1l��I�lt�~iij��z< ����TN0$3�����0��K �_1�T�i�5�͘�7B#��5�����fq�wyd)���v+�g�	,�8D��>�mas��f�S9}s�`��#,��r�YUsLy�9�����0�63&�(s�Q��'x���J�����.�L��Og*�Pw���j��束Epd���or���b�vV{gݧA{#�i�=h:�
����EY�hB<�4n�Gn��|��w��� ��c_�a뛖��.�Pb�:�	�ʗ1��
IRs;U��2.s4ЮS@n#�3�yk,���`�owϝ�a&��l9���ʳ�
��u�&dBt�"�b��d�x�����Kb�+Ү, ��w/8���1�`ń⽹e��5U��7S3\iQ:�u�)�����@�q�ԥ)�h8��V�v����̧�p�6r�����pTx���P�=����F'��v�o�y��Mm_;��y�M�m�3�,����[�g��;��u�W/&��}�9�[u��g7���n�e��}K�ִ+�K��B�a�ȓ���c���b�39��A�wU�4��m�90�#���T�+1��#V�s���^�� ��mtW9m.�v��J�ra'-��8W ���X�h��Z��:Ҷ�i��,�����a����5y:wD�����,#�@��Lmޗ��Fr�Ŕ�E���o;�8�ӓ������X�v]�9Q�GuwT������0K)���"#-0��B�:�"C��� �
Am�FMi�`��Vv!�U^P�F�F��#60�!f��LӮ��`�H�DK+�9҅��|��fܭX6�ҘNgh���o��Ͳ��B@Υ}�Y����[d���ev���-�-�����	�Y
�7"�:�                                                 SV����{<�����!�N]Sj\ôj�Hkc�X��+�f������M�����ŏ�v�RGz�+8�c�Eq2=42T볦���v�k]Bb�o��
�˥;{@(]�;>-m���yzլl�2�;Mb�ٳ4�FQ����'jd:҆w1�rs�R�i�!�ޮ#d#�c�{2��}R����r'w�.K�05�Ճ�9�;z�]���Z��`�ٸ2�N�Ef�X$R(��V�]Z�P+��NթSՅ	�J	"iY۰X����g��1�Y�����w1T"�̻��[ӬW۵���Zѻ��P,���{��,.�����j�[�;u�q�RLS\"�̊�*,dʴ@ɢ�
�<R���鋓�K��ᵞ��O�oaEkD_)%C2s�FKE�V�r�Suw�	*U�N<�^���!TW�W+�=D*�R
�c,��ޮ��h�ӕ;#���"(���e�H����P��{f�MݔD]���Ʈ���jU�6��by��n��7���b�V�K�r'��[�ZR Dv��:��^Ԥ�VY"�)[+Q��V��WtM�X�떡IA�(�l�����nɝq��I6�-��9r�v�Y��mI"x�6�U� �		�R�"i�22���`�h��ʮc¥	�4.F��E��������%lQ� �u�n^�������`�ٚ�� j�4;O�VB�
U��c���R���g�LΔ,�U�MA�J�5}5�SZ��e53ٌsp�&��,-mF�������i��rT����cljz��}Vp�}��(��\�J�-r�,PD��P���9�o�.-�Q��]��c{�uE��\��Y�[�,���7�gy�\�ܳB$T�a�ۦIl�U�Kd�#WL��%���[!t�(�!)k$i�DV*Ս�%�jT��ӑKXGJ;���         ���#�sk�'���j�M���H�&T��e��\�[Y(V�!)NRR�Ös^�%��50��fE3��[a�ר�յ��h*`�,��EQ:�A��j4G�Y[r��F�z�d�[
ԱR�Л�M
6	ƈ�����4��Hث��(�)IdLh� NJ�}ڍu�.�n�*N��[k�FS�o!����c���I��0�O�%�O��ӏ���g�;* F���EWS�}IZZ�zJ��!��3{6s����>��A�{��N^d�)�}����C��H��'@�~U.��V��m�a˫Q9��]Mo���-�F��ǎ�'�fӎ?y�D��gۍ�|Y{� : ��^�|�`��%U}�w�"�RN�Z�JI�L�e����E�3�\��4 Ϋ�)�/[�u��o�Hh8�G3�IR��m��{(c{$z@_��(���P�`I��Q�S�m���P<Q�T���J��9<�@)��*�B������8�`�//���:Do>����8��vA�y̵�a�go�D�)��Y&_'���z�r˰��Fb�^��t���Jآ�D�!!I����e�Æf/��N���#�
��έ�Ìҥ�r������4��w���S +�!SH�9�O'>%����qò�huD,#����.A�\M*�n�)u��F��@u]p$%d�Ww;,�S�9 T"	��&C�oVP�|�
̸���fVd\��5��ꏇM�B��qV���յM���F��Q�M�,;�_�B�_�8>l��d���Z�[��x᤻�`w�2O�[�/�$�wyi'I�5f��6wF�%ۧ��k�8� �U�
�AF#~/�C�Ҿ��응1A��
�󒮸X�9"W9��O`�\�a\�׋�����kCu]'eOB�[0>gq�[��F�;�{\���.�.���P�X������@�Zɍ�T���T�^\=��Y/��/8�A�$r�Y��yߥ��P����IHZn)d�ש
�ɗF4©IT�S���Jʭ���xӶ�i'��ų�*aAzDP���3�_'	3�~�u��M�&̌��G7�w�XX<-���>��os�*7���I�س'�����%���T͜e6�|v�c҇^j���������L�N��5�w��!y�w�y�5k�'� ��b;��C���`(�	�Oe��!ܖ�Siw�E;[���ddײ���o]���*�� ��T#IH��j��*�B�쀹����u�w��95�;<TX�+��h4�\6�K����
��T���=�L
v`ƨt���F��T6�{K�t\r�)��~{�_0 0���1���]44��O}�bg�e�'��d��L�ݵe��/lg2��>�Rۆ�D>�e�p۶�?��]��C�]u�h�����N���9 �P3�z>
�Ow�.��ݷ�����e(�V�FT�+��X��L��H���3j�,$\�h�|��d�����;����Cp��w���k������m֘/��C ��DA����$>BS0�1*��7Ey�����:�1�.K��<c��.�j�)�='(� ��t��[�O�X ��0��@�YmN�%e�
wv+�k�C�9$>���Jx���c�㸶T,O-�oy㋣y���m�-GuW����{Z���៓�?�q��1�i�@�IЫ`3ˋ��j:�GF�w�g\�ohO�3s���1P��Ғ�I�632Wy�Y�f��r�ފ��iV�m�Cpi��թ֯�%"���+���z|��jfu�WӉX7{��ڲ�NI�\��͋�V��a�c�J�rb��mh�DXq�ЉO>ف��Ѩd��o%˧�\�o�k����K�5��A~��LE�cu8��u�{z�1iZ�,�zݝ�wq��NZ�q��u��ܐ��[ޘ' ८�p)K`��}y0)ޮ�xU\���D<��5V���̀m�P�p�(�;*9��u�Q�hТrtK=���
&3�7�ퟗ��x����ӄ���A��4GK����j�xZ�qX����d��'W-f	��;��z���B7I��*˖]�<���^!�]�!|F������f�>Y������$����BE��ҙ�p�k�s�˃
���"RM��=��NS'g�J	h���f����W�z[� �N
�-��*�[���j�Kk��77��8�ڴ~�	�U��@��N[��%��-���F�}�:T~�%��n�V0kky�x��jI�5��	9���ݛ��ųN0w�z�n&�W<�+Ӱ)A	s�b|�pj�F�';������͔QMA�}�2�Z2� (         8Ez�f�fڳ��g<��o��[�w0q�/�c;8��I��0-8a%G`��ʰ�M�6j�D$�&|�r���+(�8:�(I'2�6,�E-�$*��lLjHꌱJ5`�	lr�U�
A�m��q؜B�*��Sy�"�qL�������e�1����A�!hny�i�U۫%�ń��t�i�Z��,cp���LFR���3<f�+%�}ny��PyA�S��������{�^�K,��<�^�ˁA\�vt�ϛ�Y�C��?��G�<��b���/�����a�TS����g�7��z~��7��ts��P�v�^,�A�;�/U1W6�L�nT�����K\4��c�>񖆝�;�A���-Ev'����{�/ٵ�\��GD^�Yq2�A��lI��}��2��TN����3�i�a�v!��#��f*��}�z�	E�&�.���� ��V��꼟4���us���=���1-&=�׳ׄgqdc�%��}wG˜��[�-0v�r���O̫r7�adm�Z��'�7`ȣ$�Rn�s��l���a��uG�P�]:P��pp���A���p�W]�R�;T�i��wW'0�r��*��͈[3�8N�3xv��V��ꦤjc���:��e�byvd�����dRe��LO4�����(�+-]a�Ur�jGq4A� &�TR%�L�UF� H J_L��8mJ���u��N�s�
7��].Tr�7��*=���U��36H���i;=0ȶ��͢t��"[&kKla]yd�2���$\�v,��ɮ�^caa�Z�k̾�@��x����8l1�%N&%��|Ғ8��9���aN�$��N�M�P��Xm��<71��"-�n'��� ��׼�
��%�:�X�N��;�TuЊ�S�T3u�YE�.�TvD�B�H��N���&֍6�Ue���Q�Nxōt#(���Ck�=6P�RJ�f�33�n�y~��%{� 5#4�Lr%V,��# 9Q�g6��G-���b�姯=���i���1~ܧK�ԇ����]8�!v�x��E$�(�N:�������"�"�.p�/�;SR-��"�s�!�G�Kh��"/��V��ڢU㰙����έ�w�����0*�\	ٛ��Z�U��-��թ�=D�I=�UW?z�'�6-u�dD��=�b��Xz�T�r�;=C��t�E�v���� *[-b����_8@�{��a���2����\c�5�"�T�y�J:N��egf���!�y�HgY5��̰@LU�FPBu�
�ե>��x:  ��z}Ngw "Y���>��ks�\??^���(��1\m�ΐ��x閨�[T�F���ɛR���ɂچ�qa"2��zPf_�v�#�1#���I��B��q/Y�׾f�wKе��ec5]�1��}Ջ������|���$�VB�Q�(����B[*�Ar�ˌ�E�BZ��˾�������D�o7��nK��ב�_8���g�N�K�\���$�o>���iJ�gh�GX�{1O�u��� �	F��V�P��NQ/=�=yĭ��c���hcL�.�v��|������=k9�'���(n�zC0y�2���D3���qQ.���0Y��wN	c�` �{bk�b"(�ۆ�n杛Ӧ�F��<�py� [�˻�LS�)]TN��i��\��&��7$�z�]?x���-�� t�ϸ���zt��M��?u��x�8Nc����\O3kyZ����C�ҖMFĽ��HJ(�@Sp��MS@����UE�
�Q����C��-����W���0m�����֨���Ul�����bu�vA-L1��2��F�)~���Q�4
�Ɩ�,�E%]�QѨ+k,�o7��Λ�Z�������<�g�����$�/��W��e�8���UQ~s1Őv�A	!����W�]|褿���-w2ó O�C��:�;eHMI� ���1s�{𴺦#��t�y���1E4"e0�qW���yM�*=�&s��X��8�����(Ӓ�fl�:f�z;�a� ��0�d�bo��h�r}Į�D�q��r��}\��tq�h43i�wf�lk4'�+�ֻL���8�s���W3w٘J�)AS���Sd�/ZZ�;IM��@xv��O�!�.�v*3�gL��~P���+�=�Z���%ֵǝ]Y��&i�Ћ��2�|2�j�H3_o䘘�������1�m=��i��YA�1otṑ��1Lл����:#nS����'kN�7���Գ��'������4cBk��-�'X�M�7�AX�,lC�M�����-�q�          E��ww���w�OqK��޿_e�3n�RX�H=Fk���� �qB)-����؇`������8�U빓0���GSN�HW$�6K4��։ �)+�A�J�*��PJAI�u� ���
ǬF�,�j�ѴP���ƅ>ˍ݄nV"�@e��~��(ֈf�C�
8���ª��Yez���e��^��%��5� ދ�p���A�Ѭ��/��c����,���#3�W��ԙ7i�vaE��Z��K�0B��Eۮs&4���5���6E_������Tc�ȸ�́���8LL�7W5�f+eU�tD���V7e�k'��i�($�V���[�C��3�k<���ȅ�P���^�.�n��m��F�u�}ǵ�-��%�qV�̙��p2�&����똖}�\���O7# �E��c#\�7��G�Z�_[�͛X�o(˖���;�$�u�Ge�8�=��P�Q��n��u&���Q�v�v�i^��`<<yݜ5�x�onq1����b����w+��\�j,U��-b�q[m����h`��%(��gp^n���-�܅y)�����Y�<�l���#�RW&{^�#�z�?1���ө[�����&�gp�$GOا�3 �gAߞ�vl�H{JB��JA���]j�Vfྥ`�t�Դ��r�D�s���ؼ3��j���6m]��JjQh�<��td�M0��aH��ʕ����wZ[�Tp���4`�a�$CR2�ڭ{���DD�5Y�8Z�C9d�X��f��LoR8����ݗ
Ϣ���"5A�tD�s=���N��W������a�<02��0�"~FY�������.d�f]���P�v̀�N��z݌��.ѓ�z��y����b|Թ�w@�w��.�Ы~�f޼��Z��ɍ�0#�C�kK;;�5/�g�1��.�¦�0�j�c��ŕ���s�D#�\NK�v���+��P@��&��[Q��Q�e@�Gk���rV�ӌ�e����"v��W�#T?�%�\�fc����߳T��:�����s6N����,�eܻ��V#��=�1�]w������zZ{k�b�[)9mZ�o�͘����f<Mχ\��5��AR�'�]^�{��5�應*���cM�e��44�;��F�z��#�����]�i��������븷���wi�z�u�X�� ��j�7�����	�S�xk+j�n��敓�^R�t�s8�\�����2��ؤ)����:�Z����F#���v,�{Y�j�.�;�71��J^B)M����W�;�]Z�\��w	c�L����N����Ytƒx��i|�;2���/��-��2`܉;m�OH+��%6s�HV��0�޾�V��9]�Y�1�+:�gUf[�Jt��N7]R2��:�m�]��>�n�m�S�cZS�ZK��la�O��u�c���������<��p�ޫǻq�?U��Oe����l J�]����K�j��)خ��_[tlS�r���Ε���a��:��9>_-�Vb�U��&vG+T��/6����@�:�'V���AV
�:K���gwd�r�zuwOHYI�D'���HN��R$4�J,U!o�^�g�����ř-8n4��{d5Kk^a\���p��Y�F+��ீ5����qڸSW4�ڕ��?]�e��Bj�ErA���˴lק�cL�\u�b #H��$�A�JaO���iX��҈��X�I�W��G����w�w��8�Xyw0 HTl"-Mv�.�,���%Ț�Re"�F`"���&�H����/9��iŚ��¸�a%֞�y`��X�̽ݣl�m���켲��f}�r�Qu�9M�3h��)wE�-e�_!-�Z��sPRHY3)�7�ow������m�8v^VaN�U�|�|ym,J��Q�Ð�Wf�N���\����.�y6n!d' �MP[]�ς[j�N��'��7)��B�}�` ޿��6��=b��fn'e.���V��(�;�r�2�J�2�)ڬW3y\E� �B]�F=��oY��k�S-2a�f�Y�(Cj������p��E�Fq����|�d}�MŅ�W;���P��3��Ԧ�j�����&�8�V.�;�p�&t�T�ȵ���q��p��цgּOD!�{�����Ɓ >�[r�h���� �~�n�p��݇qp��2[�����a�@��s���u�"�.w��Xkm48z���b�@U�;�p��1M8MHZ����H�S�VMU�Q�\�T# �Dz��6\��̠�D�m}f�vQGi�ӌ�Ǟ�t�a5�{&���3��U��*���}j����ﾗs��^������s0�B�.�^�"���.��%�en��q�yC�+�'"f�B���t�;�:��f�iu�<�<�UK7V�vX�a��8b�1*��xPNa��S60t���hVU��PʧE���t{[WI��)�ݒl���xv�����XK2��/s�r��k�{0�[z&�t����znh�)�gȋ�O�n=ߖ��u��|PV��5�͌N�M.�0�� �'53�Z�oZ���̗Vh�	
T Eka�sD׻ww�|���99���n�e��oo�ňs�e~�KN�莜�� H�59��ߍj=Z�l�X}��t�JD��J�ں���ۏ?.����_��D��k6����)KGl�+�R��p�"s�mW��A�%r}� �v" �=�����4}��P�9l��^'���u
y>^H���r���}j��j�욡B��= �Aà������=`'W�xzze�fw�1��qv�m�]^�J\L�*e�;��T�b²ӂ�w9�b�)af�Y��ò=��_�o>�x�Ɨ�����L8�W�B�;�Hn��ʃIu3w�Q})��0�C���xBp�CW��"�a��2��8��)��M���1�P�݇�|����!���>�c2׈�*f(�r�\��ul2&��3��LY_B�X3c��|	.+��C��J���{�)���~���P�q7�=jr�"�F�h9���ۓR~8 ?��n;4�[�hem������{��]�}3h�RE*�:���P�F�A�
�'�����NY@         NX��^�����Z\3v��}�[�C�y��m��}}/Q%�qY/ox���ɔ�F��*��U6oO*�,�TK+�dadH*�MȄi����:�-��:�Y�(��Bc�)P�n�F�RR�#Q�`����)r�������Gk���#��X�WA=YF�Uh||7��,��1������w(�O1�B��&̳�b��?N'���*��5�a�^$]�S�^�(��{8f&;�A�����>�a�q��΅�ɊVb!AE^̈�⩘pw���ڬ��Y�m������*=���v:�z��H{�I�xs8&h���� ��C�{\o3�.Rc��Od̘���b~��ȡ{n�ʖGy]L�#����#*dҎmeE�G=�z-��n���M��Y�t�I{�-z!%Μ�:��[wv�9��K�%Y�]�N�uWc�WU�����OM����2ɼz��bL�2bP�vg!᪣c�/���b�{nws��L�S�t���t�YvՋ�ߊar�;��2n�O%1�[�L{�<������C��lMƜ�m����c,tu͑3�u0���&Ӫ�NRl8��>�"��H��<�O�jbq�|��y�I�����#~�+l��A93���cU�w�f��r����)�����qo?�r�,'/=��a����s�̫� �F�+q�oƍ��a��D�$p��c�	Y�cs�B[� ��[Zt�|ꠥ��[٬S�����.�˝�Y�-G%0M1,�m#a^�rV�,�mz5;��hO)����2����o]o�����l�~����T6� Ƴȭ�=	byJ��7]�[/�rw�.����6L����[�Se)������0T�i�T�tRZZZ�`�GZ.�-�]�t��5��k9LAn�ff�ᱞ�sy9Hv�� "-��AO����E�������)eþ'�R��jG�'B�X2����Q��}�;�\�4h��.>u�t�ߵ�*�᭨�W��lܙ[���yL���A�P!�6V�N:&Em��
&-�
�s�t�1ޚ��{�#N+��CAD�nme���c��xV@�x�{¥���StWGO��S:T�X@�w�/�ʉ��KB������o���L�3"��������E{�ڲq�H� ��2��e��P�8>�9e�",�մ�}�t}Jx�d@���u���%q+B�c�XO9��ŭTc��Y��AQ"(�0� ��(�A�Da.<bcoo;Ӹ��u'��6q}�ـ
�dv��6�cʗ|��W�90�+���s����G���B�hm��,#��w�pVt�s�w�/�Q��n���4Xe^�]{(�Xku�	� ����^�k%̛Qd>�~��� ��dz^G��cW�煓�u�=S�¹�ꪚ�`)e����ȅ���]�MO��mC8ٛ�~{%N�ҝ�.�����n���壕JV6���>���_�2k��|O���@g@}���Z�U�kp�) ����M��s�)U�2Z�l.7)�0Z��D�ʺ�)�pŕ�7��8�s5�;>�"ڰE@�	��پ�gp����e�s.���q�gd�b����Qp�M�i��9\������X�ÇI"�X�g�b����L�c�r�6r�����r^ (F�X�l鼧T���!��W	�Z]=�^���L(l��!;�_^߫s���
$f��R�xC�v��G6w,�7�W]���}��\)S�Cw�m2|�]�ɤ�B�WҢ�����I� �{ ��D5*���Is�snu���7�y����HM�Vph��-vodE���յ�����K��P����9�0��q,ُ!��z�
R2�`8U�/w�0�� ̓��M6�.K=s�{�.w+}�� US�.Wq´*²�����R��&�et�&r��鲴W(x���zNTh��J�fh�����Ц�v�MB X�SU�=IdZ^�n;���u-N�.9�'N]ؗJ��1�R�jL�UgB�wʓ0ʯ[��4�XR7�;��� D��Dx�.<-V�˟�m� >F1��hm����S�L��(��W�㖓�ty��Kt4h�������+�	L��sm�ӏʲ�9S��51�}�zϾ��jU�E�gXe�xʪP�It��}��a!����\&i�YnˑGB=ִD�%N�_��a�O��|°`����y�,e�L�X��n#;�-[��E]��Q�m��p�x�6��E9��pa��Y����h�r^�U��06f�y:�&|a#��Bv�s��<ӻq�����qrZw{��"�)�Q;6�rj�w]�        �g)�*�ܼ Ծ6���,>ɕֱvY�+9��z1��8Q�H^UKS;�30h�@� K�QJ�����ɷ�5@��P�+j��䃶�'0m�W+�(��V�R��aKM;[�eˎQ-h�4&�u�A1�H�D�l�$$�(䪚u8j���4�d�������I`�j��_[�&�RN��!�wH��@@8���,}��tzN�/L�M�+��7FN`M�KX6R9\_3��uݱ�̃�d�Ȥ���w�)Os� rJ���ny��B�ݝ�c�Q�t+��:������}�Ib��qu#;��8�v,��a��,|��xc���;�B�@h+�p�F�%�P,G8�ݓ13��>��1PL�V�"����E�t�
һ��f���Kspy�V�2�+���A�㴦M�}�j[<%�a㩀M��&��Vu�%
�;�)=�O馽E]�����4���t�Ǻ��AUg�B�h����/7b9-��g<��s��^��� �+��
W,V�m�M:�,@P$9e�1��n)-[~��5ە��b�S���qUѯ	:�v�((<��-�=]1��/�ڵL�q�Y��`�K�vv��n�,�_~���Qm�]�`IFu�F4�&u��cc/b�&���^��ξ`�јHoT����,�h�@C��H&2�@��	-E \&�;��2�oo�k��!���24[O�waf�{��W�V�Sım� ���q�F���x�;�&��v�KpobU3�9&N3��g�G�q�m˟wp|���g�\�yBc��p����7�����wS9��y�i�ٻ^�,���)�C
'!�g��旻{�}��b67��t���k�������51\l�WS�7��y�F�jKH��Zr�s�w$>�[i�L3C�o�}��'������)k�Z�	�a٩і�nT��9S��s�|���o�$'�\@�`�PV�$��ZTIj"��8��)b@�p�H_B��5� UZ�����SlgO�_d�,�l�K�HE6@++vu{�M����/y��z�Z�P��ddu��K6��zs޹Ȇ�i!:ִ}�d�m�59	uܛ7g�̞���;���fQ{�����L4�2R#z=`H�Cs��_Z>աR�f�qc>s4��4�e���*��F�&d�{��T�U�d��y5�i��8
���):���tzaնM�Y����E�=|.�C���&�ԓ�.�w|_�ʗ8{p�������)4���-: n;��Y��#9�T��P��=��Ъ4EN7�e�����q=����11΢PƬ�g���܅H�ܞGo��\�D�+��+ݟ��«�+�zgl�o�^ZX�)��޷�UA�q�ԃ�yf��r�$�=��o>[��n �/3,�5�FXGj�&�;�
�W�MGj$�er���-�:5�㡍�0Gtc:��}�W2!�ˬ�A¥��{��ݴo3x������H�'eGI�F�F�ˎM�����Ւ�msӼH�C�z�3I�u8��B�&�-A���F���1��d��8���-)��,�����%@��d�-��N�Y��{���$�P)tNu7���i�
�1�!6��u� O�N�G��fD�gYBy����6 娑w��=�����D����5w����j�*�~���4M���e���^��f6��c������fZ#�.��2v��C���'M�!� �_���������$]X�[1�`��?��i7q�K����
/����F"���Л��]���P{Y#]�(��8�7��&���`��?��j���Z�R�D��{g7N��|���HQ]v��zFJ6
%̈́��+jr�T�5���˩DTHD�r/P�S���z�5/7<g�V]Ϊy{��������}��\���Éb�F5pK�wdȾ��t��8���Ͻ�i2��[���Cz��t���I��TH��P¶F9�m��[��nxp~?S9�����������&�W� '@;�pqzq�xMN	�sT��D��<����]�<��^r�$ɒ)�bX�L��S�`k�����ٙ����S5��f�o
��Y�zi�K���UTe8�O��}=L�~L�2I�l�mƸ~�����جX����}��3�L�����Cgt�lCV�%dt��C���{��Aܼ5b���ؖR������Rͭ��e���7+�W%v���z�nK�N�v�,ټ�����+2^K'�OP�[��C��������ծ��r����[���u�cP޾Z-rE/s3^Z�E�$�Y"���ȴ��hq���]Qetڷ�N�Ɏi�r�f�/��yI݂�����f���!X�����;p��v>�ɤh�3/�̶�N8����o�'>�mY5;M̜9�+�P���Zkl���z�f��Ƿ��L�t��7�+�bj^�]����+&�����쮮U/{
�]�o7uN����Xe[�V7�s���_d5��̇Q�8ܼ��L6y�6��Ir12�d�2��
����IF���W�����fK 1����f<՗��Y���#�[��_u2�����-.Z�ٳW[�q��fX�����@ޛ+�
��Y,��M��;:�Ӈ3^@8I'����N��#iV�"q�|�&&�����
t�'cci���
)B<�K/��'��F�jh��ΆI=v��K�juk d��_n*YK/��әd���fNY@H5�����"��cMAQ����j�(ZVP�@V(RKeݙ!u9�o�+�Ѯ�x�g" J@Аy7l���\;��o3�ק��Xe���v�Y�+q8䄊I]�WY(�d�JB�"�WI!@                                                 P5X��$�ͷ���� ���U��v�3�l���3^����㼳o]��G�-ł�ݲ���o����)��Q�� d�϶�>V���no�D�K��B�c�b�}��ki�[On�mr�0>ܭ���f��m�̼�/�I[����Y���*�n5�Z���ӻ�qt��Q�T���CM�>�}�WK/\y�eA֎w[����k���x3s\�W�e�n���:���vu0\�ih��YX|�{�Xc7�D�K�p���ߑMFy�F�hܛ��z��6����M|w�C��w>��ږ� j�ȂEV�\�����,s�o�B�y(m+ }�²ޣO�&[�p"n�e\&�B0�VKǌs�^��H�PtuN�&[�e��Mu�*YS�LS�6\�����n�Ŏ���3Oo�:�Z*�7�u7G
:�@���.E�7K�Ȳ�ӈԩ�QS�]9%��8��v
'$c���%zcu��T�S�G�������:\k']�ȅ �Em��9��!S#�n����U#u8��"�&m96���A�!��NjG�Q�i���ܬ�����9��Ʉ�u�7F���V[wl-���rHY(�TK"�mn ͋1���0���|fcnU�pMv	��D�� �M*-Z7'1��Q�� ��a�8b���
+l1�`GQ��;GU��C#���0-M<��(x�j��IF�%qA�`�`��N��㚑�CU:�/�=2�����$%UTQf،Y��%��	)�T�Su�u[C��wM�^Je�:֘��̙TȜ,(o���-��{Y��.�;��lh��.Țr�Y,��qMbB\���dk�vBD�#�����Q�[
�F�dNV��)c%���;�6�g�M�=�J8�uܳ!sQ:jSE�#�Q�4�}�3%�m�ʇ̔Q�A7.[Sh��l$�p���HP�         (ϧ�m���q�8���>��ЁV�g��g�ub+c$��1��TEDڰt���r����"�b��u,y�Yhu�Q�j��B�,c�K�]���U�ܕC�9\5Y[�5�!%��?8�[,�X�t`�,>͐���y<��.�tC����ԑ8Z�4VIH��� �^U�sY�lԩ�[C+R	�+ZpD�u8�c�"�SLԿ�v|�;q��n�ը<[J�6�y�ݥ��gn~@z���2���)����j��o�7�Y�)�C�$"j��7j�h�ַO����z��DG4���V�J�����l�Y��������zy��"K�	��C���;Nh���q~���c�y�eDU���E0��Y��7n���Ve-��Fe�T�5Cf{ݪ�wOvA}/eS��$o�������}���"S�cI��I�=�g7gL7-Ә�6=��%�3��嶡kk�/"���5��ɨ<s-1��Id�]z��>@��iw�w*��l��l��1m߀����5.�Y։wVa*���:���=�`j�
���8haEl?�\Yg��W��O�D~d�fַ�J�k��m��p��7b��0(�6����<��$�;%F���L�Q��;o!��^��4[�e~��Փ�,��6�z���v!T�΋۝�V3� ��AM	$(�M��[d�Q�&�*�_
M<�z�&��w�6�*�}�ﯴ�i��e�G,�2:r],���{7��|��ޘ�+�c�]����$ ,�ɱ�d��} ��2���%sl�L>�m79�5B�OW�F��`%q\n�7�w����.�
��C1����k�8�b433��T��4���p�5uP]� _=ӥ�|�j�a X��糕�[�oZo�"�
3E����y��f��=�J4��I�\j�ν������k����2H.^�+�n2�o{�M��e���3�%'GH��~n��m��F���t��2C�l$Dl9��,��ʠ��B��%(��y|\���~}1�v-�Ӊ-�Ft�^���i��.����}ha�x���P�]�ˉa���}
n	Y�!����z��`����5�&Ve�R�c��p^�W;��7S�{h��G���GB�w����B���ڊk�G$�C��-��7-;�V��)��_M���̦Ͳ�-�f.�I�q��੶Kͳ���ϳ�u/�`����Xw���i��n�d����vyd҂=ޥo0g}k`��n��!�����%;,CuC��c�Pa���b7�;]\�F��
:Dy9`�!47�e�F������M����6��4��|��֪����b�H��|��oHDN���ww_^��/k@َO+Fo2S�#���Td��}9N�_3�_�ݵ��fݎ�4L:5�| �b�[����#0��R�j�ڋ]���J�Rm�32�V�Y�Nu�����k��i�S��K���]�Z���o�#/:qP�{��x�"����;�Y���ِw�-U�]�ds���%t;��@�F���#�o,��#��^�L��G��[F:��*�v�a��%&b�؊�c�����3Ӳ�=ݐ���{9[�e�ؖ��S(̞2e�L8��������	���]��y2t;�����Y�9/mQ�B�%��xoSj� xs�mL���@����h�)� ۽}j��P=w@��u8�E&�W՜�U����rD)Q&�7(JL2Gn�����ooD��o-�Ž#��[SWjl��q�Ҵ��]30=_��B�]�	�*��N�$]"1�M�9�.`��<0qy3Z�� tz'�y�2k��P�xV�J��)�5d�-9�3����`GZ����n�oj��� Y,EF�n�H�Ylt��PE��2���it�M&v� kkg�s�Y0�d�}b�+ꓖ���nv����ϱ'D���Ĺᄧc�(�ar[�-���#��hU���r��6]�	o�_�Ź��i��B��mi���.����(X{47��C	:d���Ū_bQ
u���Q&s��`�Ų+XX�)�ƶ�1�>�T�BX� o���os��2�g�T��eU^깕�nᰍs�P��n��Ź�\�7K��{&��k<@FY֟w<EL� �#����#%��AE'd�udd�OƖ�Pc��*Mz�s>f�o0��C�L]��",\��+�9��,ĩ�H�?���xa^�J��{�O�9pR�[�a��U�v���AOE0�F��Wv̭G(         J�?����9p�U\'\:�aYDẶf�.8Tu���)��Do��.WA2�,$<�ړ[�Z�0�̪��-+s��ɒ��K�a[�� �Z��/~��V�!0��Ѯ�-��)wo��MUqZ9d�V��?��M�0�Z��q��$&�:�V����� [�1�m�.��6!6�[d*��8���Ie���#e�����ŕ��#�����Z��'�6q����v�WCd�)��-sr���n��zc��lN���*spE7!,ό 
��D�<1�nj��3%@�e�9�<�.����:w)�!TJT���X�9W~�8N"s�TEt�H<_�CP��$�x5��m�I�h�= ��y,�E+hoz�o�����-Ņ����ӻ9�m��zT0�ǽUB�ત)�'מ�c2vyȓȎ釦=1s<t�)dU<zzj����A�b� Qf�����oM}"�i^4�3�{��&�&�x rc�q��G)f�h��s��S�l�K�ND�#UY#���e|�|�\�"��R!E%� rڨ1�T��n��Vb(6R�[�mϭ�m/���"4��wd�saCv�4�톤2|9pvy1��R��*�VE�m�0)(2r�<�aw���Y֭����_N=5��F��g�1D��|X^����c��hq"z�@�	
���p�Z2��P5�tQ)V'S�,�93����F��Laf�J����)�vlt�N<��q7���A���K�_Y�D9a�C�H!+uk����Y�ǡ^� �#��bҸ�l�e]��o�V�X�;�{��P>u��6|\1�J���1�6����EC��9<����U,������VϘ.�.�K�C2x�1å����!�G��ȓb"��gY"��9)e��ee��J�"��l\P2�\��b��㳼kY�����/���T&�g��Shq�9VY~ #�QR�U����M�D��S%Q��U"��m�#������p����\��V}�GG/�ϋ�xĄ�z:���Fw%�Njf�;�)`B�c��d�
�8�Vi��uuUR�K�ٮ�W
�.i ��qܣ��s#e:��4��D���ۺ����{^�"V~ ���(b�?��N�#�����D��o[5ݭ3rĊ�k��it�a�̱Oz��p	���W|�W}��}��Q�$�,�-U�r�!#Q��D �4�A�x�Z�����z��)ؾ��7S(�F���7�ޤ�u����2x��v��U{߸��Y��9dӕ]j�����Z��de���M��gNc�.�Or�6Y�u�S�!�	����R���zC;�w�݋�8sc����<�]n�d�Vđ9m�e�ʠ�s �gY$�.��]l�
Z���}�&~)_���pO64]�Bd�(ت�Ycx���؋Z���Q�LY�έ���C�9��pYoIH���h�wj�ȣȏx(n}liI�E\��/�`�z/Fq�)�Zb���E�U�d6��4k'�4�@��/����R��ZkÑ��]�EpW��4�>��Utz����#�ՠ�i���e�,5����{���6�~�S�R^J�\�w��6CͲ��$�de�sŐ��C�	Dԍ̇�{º���_�2��Ts�|NQ�΢�ͮ�멦G�6kM7(G���0n�Z�jNL!����R��y��[��*t�_�B�U��0��$#@�@��L��y3�{9�<j�u��E��y:���],�.������$h WL�L$S�"B�F���޽OU+qȮ4�Ћe��^��T�\��z��
|���ļN�52��)}�]���r�`1'%@
Z� ?b*�ex)"���J((�"��'?��f]r�����+La�D�jCI³P�ԃ]wD��qŋ5��L�d��2��=���z�r~��� fO�}QO��eJ���P�zm�����r�֔X��e�q���&�&�h�у��r,Ff۸�8�<�6��[��N�\��"��Vªlq��ѹ��qܠ�Q�R(��yK��CxǼ�YOPk�TE����;a���*2Z�|�o���-]#��2�������"����s�02��f[�5L�~��X<�t�ز�������5(�]H��YK�A����U{�\�WΛ���Իk��3>j��y��m�����^����3l�����uA���a�v�Y,�Qx@q�"/F$�I���=�        �ݳsr���A�If��D�.Y��UKXw8�̧�UH�-��Q�+o�ڝ�Y*q)d+Պ�;q�kCUj=�iX��MH� 	q��}B8����8I"^:S޹$��GQ5xV�*��eU�	ԅv���do^�o!`�-�$F��FԀ�L- $��d�R[��P�9-��'	$���r�3)8�%Ӥ��˨ ���r#�C�9y���l*�G"Ƞ=�]����s+�9��+���+&y��j�*I:w���0�5w�jbf��7T9C��b��4���Θ���{���ߢ�T�b�2'��F��[�Ϊ↮�w�YU�Iߟ�^ZX�i�Yk� �h�5������0��d��f�^��0�]�l?a�<>��b��up��b�Z�.śJ�8�|�*1�ڏ�8 e�sZ�B�ǡ��Q�	�D���M�$��Fa��c}��ۗ~eZ�.�����l�q�7����y�K��5L�����H}R���H�q5��b�ЂFܱ�7`���	4V"Q�dtT�H�'``����$@\ϳ��}D�t8OkzК^]��G(����4pv!�QP������q2	;�b����Pͻ��C~2Ӷ���-��^�_9�l� �/&^C�6N'o���U��	�.�o����wIdDn�bP*�ҭi*3x�̢�ȫ61��b�K���>�ù�vs��Y&b��Y�,�+z��%��f܈=8��|	Qj��xN_9�}�{(�+�7�-�;�a2	�
�yt�U���*����CQ�-��
j:.�;R�c���\*��8�z؍�]˻\\�P���*�wG>��x��{I�Y���R�[ۢ9�\�w�&-�ڰ��Y\�oL�i�@�Zے����0��Nh,��ܓ��1�\b��m��w����7qs �{q�g`g"��1r�6�c)�M�7
� ʉ+Y~�L�H�wD���J�#U�Kb�VN��һfr��la���w�^�Px��=�/Þ��DUvɽ�ϥϲ.���r#mm�ݛ�K�vv,sG�����t�B]��u3a������'�k=Oa����|��N7�5n-)�������ت�o��qr�	��4;��� ��ը���m�؇Q�hH[53z,��5�N��}�{@�Tz����빝q�'5u�V�;s�N�waw��,ucQ�3���gv�Kx�v���x
���r���tZa�g{�Ҟ������oH'G�w�	/�u�R�H�8�6�r��Y��a������7ۘ���Qo
܆�Ǝuի"�_`,@3m)�����Χ�Y��_m�j��gu�E�Ҷ����n;�%�8���{h�9�:�ۺ|HW�xf#�����&Ÿ$n�`�gr�n�˸�k��ۣ��/�[j/2Wa��Zw�Gfo^.Xk���c�r������dށ�%�˺:���#*e���{�B��'q�����3i�7���h���������������t�
w�ﯗ�Vj׵�0���*e���{��Y-�j\3NH����ז�8۳:.�	ͱ���(�m�0,�z�[��Ҝ�[��� �l�`�F^��0 F�L4h���h���&�጗���m��si�]*�c�q�	��L�����`�.	�k�����"�3U���$\�*쒢�/���"8t����+}\��;���WMB ����`m�x/vf�-�ѪVY�\5A  ��d I��@�F<M��N�9M�bF�i�{-�C�&��_u������
�P�4ZF ��ff
�m�y-�G��qΧ�p��v�s�q��ھsp�R8��k(`�7��?��v�L���%����}i=�M\IP��cv:;I�m*�sMb�A_iD�R���i�r�GҒԱ�6w;;�D���*m��0�� �k0ej��6���/�f��<�ʵ�N�,����N9���9E���oj���s6���Z���n�rTy"����&t��Ignj��R�'�mh�N	��}X��X�7��M�n�(V�.�.{��=6�<����5��z ;0	�_
��Qr���w��~f4��n�I%�஖b�8�*�j�	'|a\f�v]��C[WZ�}�]��$�l�+��k%��\Z���ٽ��^3ۓ�)Go'�z��'�MT�Ao
XD&��t{����j2��u��s��DO��p���緘D��a�Ԍ��]0ͥ�`��f�y�=��]�zȳ�DOo�JZ�p���v��O.�F�T�B����\��ū|o5Fi����y�E�������ǽ�wj��J�wNX[klu7-��b���j��H���`��"w��,HEll��n�(�q�h�KZL��z��F����/�'" �Cwr��8/����7�����.�P�l[�P�c9vӨE�c��Y���1M&��^�{m�wN���Ѭ)�3�.윣�"��T��@�S�>n��\h6���؎�ȗm4����	=H�<�씞yS>u;b/FQ/!E	;�s�ŵ��.��:e]c;�ص5��<�)Y�n�>rF��w�m�����v��b�]������5z%xr<6�
�V-`����͵F�a
�c$Z�2�T�(4��h:A�!CW�΋΂�|��$k��ۇ;#c�Dl��fp\�إ9-Ut����*�HDζ�j�����'�j��aK��4 �v�D�� �ПLT]�\����F-��r{}��� �f0v�	�ʛ�5>�5G�8���(�c$��p��`�q�q����-n��s��5�g���t(�v ���H�S��WK��-��I$(;�r���q
*E�y>�ۇ�W�~P1Z�T+�9d��$��ʿ,g��@{7�U��B��nfl�	-Jc�b�݃<������2�c⊈�R3����Vr5�#�F���m_t��\�q_z�����P�WfEP�z�~��*/�j��̻�Ȧ ɍ3�I������p`���3��4x�3;��/5�
���?W���p���,#�j�+�t���&�W�����q�;�Y��R�Uu�Qe�ԥ.*�GH^��\��sv�~!�\v+��ڵ��7[S���cAj||�����T:j�j��Z�s�q�m��         v�nV����M�g2�|�g�����JrN�h+�x^1ͺ�lU�S.����fmd�W��x�b��yw�3X��[̳(v��]�7URF�j��֤�J�O�����"���5�x��9�A��e��84�������D��l�F&����]MCb��VX�K@RT�=S�(�ә�:�)��Zm�7�:�:��}\�.id}��DN1{3#�珖��t;6�,̱�����%
.�a��v�K��^e5�sC�Og�c�/#��FU<΍N�S��k<�;pLE�5�b��ɻ3���R1H\���G��a�p}��#��׏l2���;p6�*�x��eiz����a��4z�yN_�:q�o}�5�F���'K�x��Ԇ��)�l�ڭ�f�j�q�x�ְd2�1���/��{��U]cO7\sa�<��)ܻ�c��<Vq6�^z�f"��vS�Q70Y�n{�ެ�m��}�z��יx4��7Xc����1�cQ\ԑ��T������F,PjB�����d�sB+�}V�/'8�{��R6i>�wME�5�SS���1s�ncZg4�i��!����+ ��W����e��gQ��%EB�}��j*��P��W-IKŎ���:	Yu;:�sn�`H�8�aPm���.���[xQ�}Pp�=RN��ǻZiӟj����&g�x
E�,�dsf_c���|�|���?�k�>�<qH䌕"��"Ι�9s<1����C��KK�P:Q��pӮ�6��ɰvس��IݑN荒���"π�.��U;fN [�еεkx�pNE�-�s�O�a����h�;:(��F�:)�ݓ!p�h��閶��s��ȵJFT�-�Z��>�����*���^�(nZ׍�����梒�R
���-�HX��=�%Nbؘ�ln����	�(VB�w�@��_�n\'-duo=6��1�Zz'oq�G��	]w��I*@�k#�L�ୗ\�;cg5��z{vV0tl*j��_Y45R�j�9�vFݨ|f�ˊ�ۻ�Q��n��˙�8�n�����B6�3����|e�41��ع�f\��v� ���w����+�W��w:m�#MT�dd�*�a�w�sY�|]��n�odM������n94��c�ୃ����-�f�vZ�%��vM�r�x�L<ҧ�h�6�zol��C�-�{��b�7tF>�O�l�	���N��%= ��|~����"^����駤�Qo%��;7�=M�h�vĲ������Z� �gpj����<'<�۠����s� Op��b�&��TT�++G�	� �uI+�&@%A.���X\�W9�Ok��{Ʋ�C;+�R(�,hU3�1�����ݦds���8r�v�p�9�^�C9}܈f�ͻy��V�B�h=��<�v�H�~�K{��}LOѼTDL���Kb��2ř��e�;���Յt�n�ų�\�]�C���ES���eEՏ-u��[�������8����;n��~��]��T]�вFa��)�NH݅���Zy�fm!��<7&5\�/.����[��mvh�ۥCC���D,�a��Y��
D@�� �$�	D(� �@���:�Y�o3z�|]-vy���3yk��'yoR��N�ּ�~�F�qn�;�Y<�q��SL������
C�$!V�B���t�a5�J�Y3D8�X��|m�q� EC� m�!�*�8*GK��7s*�Ajq�j)T����Q
�/�j���: ;�FV�W9/���C���1���j�I�����]�E�N�&��%��Ya��1YhUC�z��s^��(;jV,i���;DSc ��z�k�TC�[����{����t����#�e���<�����yY��4���qS�K:�F%�/,Y�+��=��X�]�����?����o'�φ��f`$�.��L,B+o��M�L�4׏�ݑ���Ӎ�ɧ��K�ا�8���-q)��ܝ�!�f�46rVFH0���1���$t��x"�[�~3Y׳�VtE~u~�.�q[�L�t��0N�U������M���J�`�;�J�ĉ� �'[IiR�$Q !�|�t"d��I�         ,�m������v��"�)mV]CB[N{��Xؒ>pr�m���ɩB��!��E��&-`�5����a$Ix��g�Q���u+i��S���xۑfG�>�۽7��n/Lř)]P���J�c���(;;�T�"G��ʄ<M6*�RWQ m۴mF�9ǁ�r;kU��,*%�B6Q�j��3Iqv�|~�s�d6��s��5��L�������4�&�:I�[m�4��JQ�G�����vn��(���97k��ڋ8�	��s�������[�4�Ɛa�޽�
_3�k��G�1�4��3{�pb5�Qm����TAI���x��g�嶡&��<���:CW�ȉƑg#[4зL���]�f @~z����:�^u�T��Er�y	WJ����P��1�*�����NZ�ɴ(�&��f�4��_z�Q������t �Y���O#�i�_�Nm�5�Ix��1Gw�Y�J�@ a��6)��ᘕN2Q�7,v�Wt!�QA��,�v���͠�1z�e�\�e�YK&�98��T��mW[ONjRB3� 	!nؖ=1S�dF(�V7&��.mh�|�I@�ҭ�B��f`�j^�Ëv�qI��\�"ZխӬ)�#C��|�P��s�=��[��l ��˗==���iB��T�p�9B����վ�q�N�TӉ��0����Kr�n����s<�69�oD�&��=&Of9G�B�lf�;c���woÑ�@��Gw��y���Q��H �0y���h@���:��S���;�f���v�oxVjA��P��J�+o6����#e享W��r?��&/�Z���"����߮(�:DDs}��7�"���4Ը�|�߳{v�����l�Ys$��9���%�s2cV7bjж�,�e���UXX�R�*��������8-��e�qZ��=�{�8�v�['%�xjӓ��0&��������ђ�Sh�L�,d{��jz���a�3�ԾɞA��\�.��M�t�������wpQ��&.��(�{=�R��
Q�a{����_9��`����4�@f�=��X�݊y=�!������E�0�vڻ�<lp�B�7s��4p������@(�Q6�V��4􆐀:�s�����_9�fH�^5J"�1]�U2x�l�9�(8n�9��:��J�Ͻ�hW���AY�hxotm���K2���+�v�g�(����¯��#������9D��5Y_9.v��[������f�dfU�]u�3�]�.�
s2���C��͗�~�r��1�z����v�7�����S��i/�|-� d5������;Tq(F�!eb�T�0�i�TA�q۷�&��+�������%��-b����6kD�6^'x��P9Kt��cn�p7�Lr%|��+�V�EƆ��75�Wb��LB׽5s�Â	wU;[��������Q��k��+[[�(�	g�!�$r�ݟlL[WPjJ R���[A�)�~ !��]̱��g���e�t�n2E@d��#^e\�M�-e��&��w\��zL��ﾮ�ܤ��k9a>Kl5���p[�����>��!y�1gVpo:#V��I�;��X���bw���v�*�ARԙ�J��mN�Gpn�n�<�{U:�qG��>.'N��iQ�ݝ��_غ�[ݏJX��=�"d�Sd^��v*R�v�M>oZ�@��~[��m�}Ń]�������Y��:G7��<��s�$D6�F��p����b���N�qȡ*heH�	�E��T�A�:.�b`l`�n]�b,<=7��tF�y%�����b33]���,X�I*�ծl����EHJ"ذ�أ)II���Z��r�-�<���K`� �w�%l)�n�:.t���hT!-������7J���z(�VL�`�H�!�8��Fu�!����*%O/��&���B/��7f�ѰFm<��^��*t���)�GMA��^�y��<�A��'UK/H��7�ݓ�h��[�Wf�8՚�>�@�z���f�&��5f삯ۄ���W��w����*��*���P�(
������@UP�� �_�B��U_�T*�P�	 @���UT,��� �hP ����*�"�
 	���T(
����P�(
����B��*��������j�@PU_ߦ�������c��B��*����P_��UT(����*�@UUr����IT(
���������UU}��U@UUr�PUW��TUU���
�(
����������b	T(
�����PUWξ_�� ������B��*���ׁ�O�����T(
���?�����=T(
���	�@PUY�~��1AY&SY�5EDm�ـ`P��3'� a���ٓW]�ʂ���d��
�����Ѧ�6�4qE��
U]����7a���Yvh�����C�(��:Ӯ٠r���ګ�� �'���(�J
��KcH���)UEQB�U	D��EQT*��Q%T��
*��%	K��ze!"��*���2!"��uT��j��kk5'�]���l��uٯn�����m��6���m��Kv�u��k^޼�mk]�89N��Fw)UR�JJp� �P� :+nQs9���׵��r:ڙ���]7��΍�=ƫn��N{�mԩv6�{؞���{z�8�v�Z�]����T�@"�y�4��C�;wz�b�{�y��{��^�N�-��^��K������;b���l^�磽��wK�ZV�.`RRJ�
�-z{���z��i{j6��{�[�p���{��(7���^����0^x����0 �7#ۃ����^��4�RB��U7n�ûl�=(��;�V���X�������q�����{r�AG�y��:d鱝ٶ��y�N�Qֽ�攣�J�<V@Z�jIR��@w�����:�mҴh�ÏC^���= uי�=�4�z���hg��mN�����=4Uz����!ћ�  fv"B�A�]�]�{�^�u�q<9�u7T=�w�4��\ܸ�:��w=�7gJ���=Q�����=:��2��@ot�t�I��� �j!"QTU\��{�������{@ ^��iwr���׳���y�z(���炤����5��Ѯ��s�%)��G= j����	�ʕ)Q*����u݁l�<��ݚʏpίe�<޺�ރ���y�ۋ���yp(Uw�Uޅ��v�㝶�O{���w<Э 5�����)�{�ۻ#Þw��S{�r����N���k���X����=�+w��׶�r-GnX
��k���޽���rg�"��JU!���E?!�)IQ� ���T���  E?5)J����@5JT d 	4�$�)�  ��������|��2�9`�oM!�?M�by��˙�{��[����BI;�G�� �$��@����0�@�O��I?АH�BBC�;�����s�k��?���b���i��-�Ў�D6�nX�- �L�nȾim�ͽ�Y�	p�,�,����J�de��ʊ=G����gK�a�Rm��5M *]�f�^+�n�ۭ���aA�B�O���T�-��*݂2�`mݫ!�����ǆ�������	��i�%m�4�fͦ�Q�Z��v�ޅe�{50�[�b��� q�ȓM��>�H�pf�jڣDGz6;�X����r6$����5�x,�^0�h���8�Uq �>
1����X"ӛ����y��w���	nt�v�ǟ#�"Z9j��r`b���ۡ�=f��YwXx�u��+.�i�T�a*��� Am�T藔M];�K��EA�1�-f�Y[وi��F4�lS��m�k�*����*���*�5��w-��xM�v�9Y�T�tY��-X���]��g��3ٻ�k���7AI���^�m�N��{���k�N�L���nO;ǴN*�%�t74�Y(F�S����Li��4`R���?n�V)�A�F4E���Cy�ݚ���`����j�ۺ-�f#��ۇV'E �׹@��*��SPг]�^��Թ	�j`Ք��n�XeBoY��E7,�ou��ĥ�5M��a[w�p�UXfm���5Wj�驉nIb�h�Y/,�{c"�7�n,&�)�E��7] �m�E 
�F��2��:zuLcSR���eZW��FV}��3�[w��RŢ���/%�#�(��Da��+i�Q��� ���̫",ct J���YG�gV�kھ�`��ggtB̩��CSd��,��:��i�[g� 0��[��,Ū)���p� �x��1�G��ʒZ�DV��,�U�,�B��nJÏT�y�{C⴫fr
�ⰦLo(4n�Rf=z��;YQaȓ�R�㤎3�7���=�5̚���]���1��2�m�.��	��V]�9�J��H򞵗emH�9��o �t����!Z�h�0��T_�7Wgn��G(�CW۹�YT$��(��r���u�U�b� ��F3P6�`"���c�Ybee CWwS)7%��_;: �Op��4l�Ő��/)QB�4Q�^d�mbme^�0�B�#v�%B�1�8�g�h�x,*��eԊ�iL$/T*�^�K�D&�����š����HU���)�iW۾4�ΜXw��T���j�S369{��t��f�rc^kZ[O{K-V�n���Iz.�T-fb��S���˱��;4p�
��+�SjZUtDD֜.j�/���|�o^����n:�"/�jf�gxo����bэPӈ2��F���XS_,���Q�h��hx�p���B܂��ʻ��j��K!�n��Jf���ٺ�o,��k�z)Y�Uf,H�v���Z׶�pf�\0Ou��U}j�;��];�ar��n�1�ҜCˑ��NL���*�k�mޒ�l\G5F�xV�#�scBP�V#a*7)�^]�i�v@;V����&�Hn؄����)V���S���Y�hb�:��1Цp��2�k*�;�e�gwn���KCzV]=)Cb̭���"��v�����(n*-�܋�M��0�[Œ�-��&Mރ��U��)�V�
{��,�h��� �-���}����t`�!��@oդ�.��&���&�Ė<�B%�͠(V��|g��u�7z!��L5��Q.s0�E��<��痗@��=a'�~�^��h�M[(Ƙzx�z�3��jAꘝ�h�$slA[�*j`2�U��[4Oqw|;gWj)jA�j�ִ�^�rP�3ኰm��Ƭ�c�����s[�y�X"�(��"(���M�ۭ�D�}��X(��u�)�o^�˷�RMB�v��G4�X����]!�I��W��%7���2U�.�m̪��;�Q++Md |>O5�,n��v�\͚�|Q��g����٠��������1�>�PL�yupʵ��t�<���ۛGq����!x2Ɣ5��v+N���Ϣw�����G-�l�VN�-S:�n�K	y�2�o�hӨ�Kn��Z.�{��@�,G��&p6��rfU�Kl���ZdȠ��[x���G�f �Q7��:Ǹ'.���wrJoj�UVkJ�f���YCw]m�����[�q�Hf�s�)S�#�v0�o2�pO�I@]7ٔh?���l�^8��o����UDn{�3��ɜ�6|�`�ta�&_̋x�(:��/2�I���;�4K	ԩ��y�i�t������'(��ɿ-�O{{Xc[_A��?����6Y(^�1�B���i�o��c�S=�on�R�m���]oz�;�5�i^o6YM�c.kq6�Mu�Mg��S3kh
n����u[5
�(�#1ad��ƶ�8\�fF������&5��Q̬�ۤ��c뷸%9N2�����Ǯ�".�����Ջc"��F+;��
��Y�S)��b8�[XΚ7�㚯e�.Ht�$)��l�b[MU��nbtee7r�D4w��LP��z�T�yx���V�۾c7����cv�w�Z�c�R�G�4�:��XX��ZKf��ed*jn7ZZu�VX��u�A�jY���{��f٪8X�ѻJ�	WpJ��h�*��\��+F�Bm�Na�94�^mk�hYf�ӫ��ذmq
,nl�3س:^�K�œ5#�7^�N��ģD��t9�7:'��ۼ`�GN��8�(��""�(��2��.��ֻ����X�z�q�0�n�|��a�E������/MɬX��k*�V��y��̢����j�[���hH�M͞��:������Aw�8�R�DFDG���;�"Ol�2���:�iL㲳pi��4�]=�Fj	�8��8"+�m[3���In�t�Q:�4����X�PT�:���Q"���{;�c��;��1n�����gT�I�C�/BB�)�o~��� �^S�;����)�� э�g�k�;�t*݉��U�6�m�4��'r��lSaV�Y��[�߈N�����0�z���p|f�V�O᎞d�o�N����%VB��T6��l�jmE��ܢR��4�0!LR���q��ْ�h���h��b�nS��vt�QM��4�VT�*C+JW6���{���7�hk*�:�+�bn�È�)6]L����˻�i�H��1��<2h~�T��71���^Pl���L5�G�7G��k�(���:��k��s5uVv�T��1e�Y�Q��>���-�=���%��(���5�k��_�2�� Ճ��|I��v��e�Ha�D��L��U

<JTw�/�v0U ��Z�7�G������U<��8)a��߮�%GB��Llw70�� ��y1,WCU�J��wF�h�sBa���O>�^)Y����}%Fd�c�+��h�y`<pڶ !֣A�+`��0�N�*�������Z������
��U`�յ�)�[����t�S�:�7gh��*�4R=}�4�2U�\i�x�7y�F��ˁhx��+l�֞VX�N��n����W0��:o�����B� (���(���((����(��
(����(���
(�� ����(#���k���f��ֹ�Мj
6�9��s�7�/��n���AG3��ŉ��Eb(���4�J`��{7��Xv������n�#
E�
¤�)���pa�mdqM�A�	���si�w�J��A�˖ %Hx9��P��K��fo�}(�"�"1�aL8���:w��f��:`�)K��^�w�ۛ�u��j����S7���78 �tp�v�!�ӥ�U&��CA�fk�@2��uY�uwc1;��}oi������Z��.�٫�eE�yb�-T�.���f�̛�f��`�R
��h�{ί=�������� �\��s3�u�3/r���w3���dODDE�VT�Øݐ�H`ӈ��uR�e����j�N�C/�^Kg�Q��@���f��(h`(�#5X���3T=wJG�3���on���4cC�L�T�����A�{��ו���I�[q�YM,/QB�*��@F#"1ə�"8%їg4�7�R�"�^��ѽ(d�tP��HՋt��;H2��k]\��b�&�b`��'t)��IM��9ZMCbM5�Eh��`�����E�:������e�FɽxܪF���OhP�+��z5#���i3�i��*�#J�_��R�m1"4o)J���z1(i��׼7�k���G�a�̵c�i�Xf�TT}��R�ޑJ^�۹��\$���[2/ ,�	����Y��q��$�.�Y����X�i�k۱g8W�^p��׎�5
vw��)�o\�*��ߚ{3fU��֚T�p:��Σüӫ�q��k�܇��)DEDy�Z�c��5���}�k��l�þ۸h�����Na��4�RH�*��u�)m�W+ި&��<�Kw`� Р����i,U�Ʒc����S=�~K���lP" �4"R��7�o�׍���2�4��cs�	���1���V�ԩZĥǜzk�3��L߶�P�Ⱥ5���hͣ���-*�q���r�H�M]�p�-��&Ԋ��{��b�1�!�{&����d0Cݭb�ˠ�кd�ݭ*��V����2���Z�۸b���Rҗ5�B^sZ'<��5��s��zS3�Η������W�{�v�5Y@#!�KF�,WWXI1�R铡P���2������c[�A��6�@H>($щ9��,���N�P�֐��j�5��]�dc1��$^��mk��i5� ��QŭފT��)�"����=�����Ӷ�+��w8�Ԑ)��VڡT(|"�����Y�oඣ��t42����G�|*ˬ��\Kv�&3��;Z>�л8h���ΥN��)Hc����vl�y|��^pԙ��љ��e�Έ�X2,���j�m켧Z��`��µPᢝ���N�w]���-j*�eR<�M�V蛮�#m=uQ���X�۩Gd՛[��ba!��[z{���Z���,��,�y*�� �deXnKm;��aʫ�opMq"vQ�𜼍�&Ӏъ��r���$�t=[����A5�b�[y���S6�nK��z��Ċ��E (��a`�+�,�i˥�����Xf�wQ��I���֭FdL�]�;aX�x`���w�Mzy%`(l�ݠQ����y��j:��~b��1U�Z�ĩ�B�e��w�M����Ø�0�Y���Kʺ��f&52��k��;���R�ʻ�k*a���%К�|��赸���K8V�*��GjVS�Ɨ�ޣJ&�-��ѥg~��i���3I-�B��%̪5�(�����RdW��2ʥM���w��}�+E�
���bq�ZJ2���Y�ҭL�l�ҹxsL�։n��H���w�+T^�-��f'���{z��v9��E�s~��	���
{��T��h�� ���`�R"ż�c��e�Y��z��[� ��+;�@G@�2;Dm@5}j�S�\��l#{���q9�f�v`�K��R��D�ǖ�������\5�X���o>j���cت\��6ؐB	�f�v�W�z21&�f6��*��˪6�u[�b ��A��Nᙬ ���=Ch�Y��q�Qb�B�`Z�O]R����!hD��X�|,Z1�q�׎יNs��Kx�f�DQ'u� 9j�6���7%�4�6Ӧ,�5e�ˠ�0[�I��!d����z��uO�n0��X��x��M�k3�v�7S`�ь�A��IMl�H5w.���,{j'B�WOr��R��YJ��O�6%`��=�OjY��Z�״m�B3,��Ν.�C1;�w�[@V0 T�h˵�0���)f���$"�)%�!�,\�m3���C�n�"S{n������v@j��SÎ�p#�7dm�Wk6�Zr��zդL�nMݤ�R�q��i�Wڎ65�Y`3�#���1�LfƗ�dgrKU
,�b<t�+�Fh�"����x�]���j���J��������U�6�� xu���M�Sd�Ǎ>/Yn���̓�)\�@i���A}�!ud��R�LZ�iOc�k��Hִ�t��+i�E2s;�cU���w�� �IJx�᳻4}�+������'���ˣ���$_Q�W���`�֝�eaK37C��&��L+V˖'\X>cp�M����ssp�G3�b�)�J�.�Ү�n�V੆���B�*$l�,F,���k>Ϳ�me�XR������BTk�,z�Q�( �j 񁚵>8�E���ݬfԹS��a�2.�࡬�D��cg�����g,饠� ����� Yӑ0BKhٻ9�,U����sn;|9��;p�������1m��t�nPIl�q|�������/M�I��D�כ�U�� ��r�@�C��^6�}`��n��̭�7n����`�Yz����cL)�Q^�A�õx�۱��Y�6ۡ�(Ѓ���ٽi���Y������{ϕ��|����27���FPH�9;&W�8�&��%���&ۻ哷��X�{Z���bSyl��l["ɻ5��9gn�k�o-�d�����z��زE�,�'v�KJ�t>��}���<�N6�%�s|�H�IH�D��$�̙�w+��ַ{R�۝�f[��(�w��-k�m%rr�Ks:ZW��Vb��ۄ�����K��\.��me+9�9�ɰ��[��}$��������˓:﹓�t�l[|���$�aRn�b�:
��0�Ȟμ�Ǫj@��çvv�Irý,�8Λ�B��m�Lwq�L���r�2��(�=ޓ3#�3��y�t�\���n�������e��;7�%H�{�yn��G��3or݊lI�Rr���v��,Wٙ�(З-��';�v��ջ����ݝ�F�H�I�u����[��-ޛ���ZYo��3I͕۠9��Ny2�#���f�7Ğ�sR%��������3�vDr�e�o7f�e�8v�-�Fq����ù�(�8��D�r�mӎ�o7�0=��Y��L�N�dj����-�\W3]r�Vn�x�;���u͵�^�ؒ���.q'�e�k]�+pu|��E?�3,������2�o=w�)v��w�� �jV�)3!�ŌG*J�ո"Z+j�A���b^����(u�f�I'�A��{�½岁�nq�̳ij���秣Wr[43)4�i��Xmܖ��K�әU�K�j�i�Ov����V\�b�'�Of�1�u�0dG�,TQ;{6��Ĥ�ۣtN�o�V������Ռr7Yu�&a��d�oq��p���]^�T��C7P����v{V$�pn�e�<(V��ݽ�'�X�`R	�{0ƫ���qi�s���,��i��n��	�,���r3-�`L-�O*Ҕ��Ωɽ�4_n��^2��Kݝ��u9s���$�v��nҶ1藵6Z�0�q�9�R��N�W���+�\!Q����6Pjh7��{]�ΐ��syS��Y�&Q�Ί��lkɻ�Gw"rp�su6fJMָ�J'wh�f��-p���͙�Vh�,v����d"�W5��5�uٱa���+x����P�8k��&-ե�dmnR�@�O�%n�s������^�ۉ��{r�9�:�%��$[X�ˍ��s[�ͷ4��#\�ە����.�\�F�i�8�P�q:��^4��-ޒ��~'u���F���ѶgB3n��� dEdY�w#��7n�ޓ�@&�ww����������n_{�8�Im���ָ�fhy;&<s���]�f_vˊ��v�1��!�8��-�I��-٥�c}qvmhXxњ̨�^$��&C�V��Bfl�ŋu�f�u������䵤���&n�̓�u��,b��Ss��Ot��V�ܓ2�0_�ۺӒN�$�X�y��Y��ǯ{`��G����ڽ��9��i���McToyK�N���T������ֽ�C����j2�ɹ )m��97�wn��ې+��N�ckt�	�%�k��
�ܨ�8��L{�v�k2+If-�9%��q�m��&��mW8�ղ��˙6ɓn�F�P�-n���X�W�:Lɼ�n%ٙ���n��mۗ�s�KԖK�&j��v��3H������H4Q�JW^�l������r'y���|�̱ܲ�Z�W4G�.�� �\�ou�щrw/�!������w&�e�S��OY�ڵ���Zz�l��g�
w�{fn��k�V�7r��n��w�(u�b�Ɏ�E|�݃+�ǣ�G��R�sImə�[�۾�����VC��CVfv��m$0�خ��.�prd�sn�x+kUӵ5I�JDv�;uY�����.�g^���Z�B�a�yIC��+ϲ�*��g5z*.ѶL�}+S�,�r�֕�_t�e�{��K���c�)-�2�T�Uw�KS�9\����@�R�j��5ͧ���Ղ���֢�����_7�V��i�H���Nf��k�䨭%:��{"F�
�꼲VR�K*tC�5ϊ�,�y�GU�w�7$=J7ڣ�Չ㴬C�VM�i�q���hn�WC���]��ve���a!�Vqd�Nnf{2��+r����O�9�&	$J��`�!��}��ǽ&�L���w�=����uUݞSO���ǖ�!O��F��1إ�}&
	�ve�\3����/���C:�[ 5�*a�gtp�ֺ[��CXzj�IgQ�}�0�Ce��LT�Zp|%d��8�/
���r������n��5�&�^�a��>K7X�lye�n�s��:�8v�����ĖfN˛W�6`����_�B�ݼ���J�u�C۝��{1J:h�jVp�R�k�b�E���g53D-�7r�6�\%qY�huZ2��ҁ�˵��-������GcYք��toc=0n���5�p�d���Zqx�p�X/j��E^;H압���܂��׫g=��U���1)E��y����5�N�%5
��n���!v�l�a�5��ݒ ���M�F�e&�	.��gFG��o���f��1˵���Űk�����N��~��B�z�e��q׏��3Z�}y�r�O~�{{X�wO������R�Kv��m��Z��-Y,��>yZ���L8-�SA7Fi��
A�v[ڲ�m�s7��y\aM��p���i����}j3��28��jԚ¥
���:�4�ӧJy �fu�<�	��fW1an;:�k��RA�:G���K���5F���|���>6��TсY��U���)��+wJ#h�6���OS&*�eJ��<y.�Ȝ����7�@�vӝtKPKl���.�q�L:�f��s�]m�RɉN�u�C`)>�Q�|����uwk{�Vb�N�ީݢ��sE>����.7Wr�H\+->�TX)�K"`�}����G���շ�q�z{�e��L��9@�|�1�Ve�����3uܧ���ӎL3q]�V��a�n��;d�ԯ7����X��jl5w-�}Y��W�kmWs�'�<yUي�vKMXBB�;��3���'XJj5���7"�c�%�;{2�ڲˁ2K?rw�w�!��ǀd�e�L�y&W8�E�����0��)�0�V�"��i<�s��pN�w�m�Z�����P'���l��[�Υ|����t���}]+o]n��ݧ:��[PC�DVb��'$�������X�/\.2���F�].كN���+r�LTVR��*k��%Y}l�;F�R�c�*a{y&逌5�-��|�62*��Z�[�њJ�^��q[��w�6(h���������ۮ���K�YK����v����J7*�ңV����4��³���SE�I>/5V���]��9��V�u9x�N���A)��U�u��N�r�ojEy�IW\�X��uf�.޻r�]<�2�K����9�_Z{�R�¨�-wN.�U��b���f�iޙ]� ���Y�;�h�R>]1��gh�o�t+�V�V���7H���%�'8��6��[D]�u�V:]��DSj�W�<�e�ƩI�b�s���������U�,�齱�����b5�Q��§ns�G�n�.+mn /)��������ϷE�/�i�)�[Zb��M�B{���ǲ�Z�F)�Ai���c~�,�}bo,$n�jMԩ+(����-&<X�rֺ��n�U;Qk�U�H��u"�+q�
�$�	��Ba��5�%����S;5���[ �	�SjlC�J�Z�x�՗/Zܔ��:���:Zy՜��N��-&�6�C9t�׆RI�����,�,��d��#�FS�w���ųx.�/�՜�cW{z�ٻ�o`k��]
&,�<η�A�����f� �ow�g��#�r�C�R��e��#����^��A��65�eu�<j�5�`�P���r=yn j]��|{+-�"�;�-���[{��̏�&�f��{��n͸ֽ�j��ٴ�^��@Q�b2�Х)f���n�A�7��Aطr�`ի��'n`	ƶWn�w�c��v�g��F����h t�&pa�fh�:� N}�j�,IΘ�x������`���SWO$B޴����oR���v�O
��n>DL1�}H��7ywC�� �T�-����R�eoA�q��Z��Z/�oZ�-��]��#X��xL�mGj������&@�ՙ�ϋ`f.�t��4E�wq�I;�Yړ'�p�l���PbG6,6�dg^g�N�/-��_J4P+�9E�Lnof�*�v�.ͅ3`����Hlj��u��n6���Ctb֥�{34gHMo^��KU�u��jƭ�N��P�Q�� �!�4��0`���1��d���X4�����ڼ\�+�fZ˹�Wm�t�ٖ�5�НWE�;n�+�n���֧N��h���t��;�̥rk�	���ު�ÚhM���r� 46��鱛:���p�7��ʰo"�P��o�=]ӥ�Y�Ա`�gy�Jj�;;jq<oOvCE�ti�l������J굻�N���m����m]��u��Rї�wS��G�uK��Ϟ�J�7o
� ���K��]n]����NtrD��/s��p
� n5{�@fm�޻jJ�Lۚ�7��9kzFpT�f.��en�%[2��R��"��|+Q�V��:�Ѝ�w��¤��a������U�
<����X[��� �Q%�z�%b�C@���YE�rs���c�]��R���u��ռX��hp�y{�޶�r�IdV�[}��7n�7ꭅq���L�Qw��p��ӕ�w]|�E�>�Y���ʾ�*0���.5�� ٸ�vw"�^Ӈ=�y����=Wn���`Э��Q��Ƹ*�WٸܣY[�ރ��y�/�
u5��d�h=:խ�Q�c�,a�P��N_o
h�������0��a\;J��c2[�y�<��*����1
�
�%q�n��E�L�p�N>��g�ت\*�َ�ŝ� y5�3Rr	kL���C���DmtX�Z�K��[���*��;��Ѻ-%��fn��.��h�`v;M�8�uE	u���˸�X$�ɛ���F_wKk���5�����KU�+.�˦���t�vJ� 㨵]N:/�$���q�1䮍���_�O��T�[��o�u��H��aKx�s.^نD�e�-�f�*tz����/_rvKxY�����%��U���ն]u���'6�'�H����Xޭ�I�Y[�W��S"W�i�&$���Hgp��v�ľ��j,d+R;Y���gT���שN���q�E�bdz�+;c��֦��x���1���D � q�ϔ�8�V��V���7 o[��&�jAjΛ{�IڳV����!ؽe�S�+1VV�EcT9FU��o^9���n��temC���j�cem�K6��� �lbNQ�騘�*p+"�sc�q��.�4�b4­��/)���K�S�P�uj	�6��[�r��j��f�v����L ���N=�)fdS5��P�����!"��Nj�琩�2�m�J��i��+�Q=�W��Z(��1MN̳��DA��|��f���
���Z5Ʃ3��&��H!ة�O�)�����p�F#�;8�L����C)��A�ԃ�j���u(�đ��|aw+eÒeWH�T��Q/����1�[L4���1'�xHO���	��ݹϖҹ�`�,Z���S�,ge:R�T0�li�V^�*�xO̜�:F�������kg]�)����]F^<;[o$|3.��R�v�7�е��b�"�Ǉ	�s�{���h��1:+9�=��m���+ �x٩n�lU|��:��Y��=��Қ��k�֥ڝI�t��^�8�+���pL[v�c�(�SR8�3;k�J��J��-��r�6y�ѣ�9Y�"�gS���=����k㪺�'�]>�T�Uhop�[آ��mұ3�٭��z�"�p�J@��]�[hX��r��yN� ��i�_m�ҀO�;O���[u��'.���7U�Gz6�Q�ed�Aӣ��_t�$�!�GJ����C3b���+�7�7.����43����¥�C����>CSM'�,�Y4;�"0��v���`^6eB�Z��[+�r���N`V�f Zκ�oj��إs8���z�1V&�y�&���9F^�b�R�/%��ȉ�9YM�f�̓+e�m=�sr �f�L�$m8&k;�m<ek��8�b
�,2�5�G�@��3��5�3 �a����&z�k^��d6p]:J�z�3~��ݥ�o��wn��W6�˝4�3�d��S<6�4 [Pi��^��scq�n��K��ԶTŽ]z3Uf�K�L�%�ޗ<�M�Z��Z5�m,Y8E2���+�����^̈Y�V ؐ�f_��{�G�,jIt���Ӗ�H�^����J�{����-�]�YѲ"���oE.��.*BZ���3}�C�m+�� N�������b�:�X��y].�f����:�Js��� ��>�v���R�%�q�=��Z�M�J��e��'�k�guj��8�#l��M'���u��ϴp����U��ot����D���S��;�U݌I��++�ٽ���7�۶zJR���b�~� 	2 <�!Sx��ڻ�t�jh�4����)WثW�e��Gm���#'oH��ӽo�%ujɄm"�����4ٝ{Pn�4ac�D�4�Ĳq޾ҬFf��fͰlI;b�7�QdIR�9_]s��Z�ݔ��#�+t��5u���'3�Os�	i��;�Z;i!�7k4ٝ����b˹�jh�V�P���X���.���J���ݺէv��á����K�k$�z�AJ��B�Y���@�E�����<���F�����y�!]Z��<E����_V�Sm�[��u�n�k"�Ij%	՛oo+]H��	��e�Z���y��`9�T])��d	n@��	����ݝ|~2�ٻ�(��϶!ӎcX��է9K2��թ��w��Y�ֵ[�\��1�\�3�:��0��Y�9^oW\r����*S{�wn�ykݭ������Lh�E\\�\�Gr)�n5\��y��#]_� ��$��I?�	$a����÷��y���m�ٛm�N�۹�J���Fq������.�Q��`�%މW�n���IVa� 8��y{j͑�h)V����ӕ��r�8��:�g� [���c]�ZLm+���rkOXkM���k�-�G����$��٦X]��4<x!
���s��l��x�����#q�aH�A��9���e�	=�kvvt�ET���+{in=A�]�^��$��*{n���tv�����[F�'Y8���������l��r�AVu.d�����ܭw^_(Tz�&;Դ�z��+M�۝�Ɏ.%8�5N�9(��a���X�73b@�����i���=�
�{z'b,
�."]�C)Z�{P�Hm�6'HIY ��Wբ�L�����J1��-QU��_ï��ژeYT&C׻V�֑�w�Q�E~�37{2=��tWO��B6�]��e����M��QRL�z0r'(��#[���M��e������� ppKҳ��%a�*!���k���p����n�c�uա��B����;i#�RK���
��Ɉ�M�0wԯ"��RCe��j=�`��'/��]6�<�0��x_Tkr��ߑ�jK��r�x�P��a6nJ�C`�ج&�1��6���H�WH!�4j�kS2L;A=
#�3�D:�<au��Q1��bEON��q�i*Ύ���a�K!�YRjY˥�!�1��+O#�S�tn.�������fg�r��w�Ŷ�=d!vQ�+
�1�53i30��t��ٷ�j=��$�	�.�<]���q[�_n�Lfeю/�9!+������L�&�ȳ�"]�`���D�p��4c�Ͳk0҄�Js�f�� ���:�ﾡ:4����K�V,�S��Ki�[EW�<�*
�bY(�EP�,��ĺ�>�7ɛ��W���EtYMnA�K���K�<v���v�j�@jBP޾0�d��4�!��� ��w�O6��直�Sl����`�(��g,[DTRf�k���!���!]8l6�B%V�@sZ3�;��Pv���*O�ӎ&;
�	{�.�jm[�t�FW���=�
�i�\����1�0`b	B��)��g&���ᮗ�����Zr%H\`��q�2G`���7/>�o�� �(p��(uZc�K��hW�U|y�V��}u��|J0b
"E �BE�TE������ ��H����X�>�tb�-�[�^]��N���h�]F�׼�=�ǲt��Cܰ�U��+�8Yd(�(�86�����Dv��h��KNI�K3m�ة�N��A�B��gS�"{M=�<�\�!G��[�7�N�U����Oݴ`C��wg. ���w-�0�����Uq��d����F8�i!L`������d^c�2+Q�լ�)Έ�}2Gjt�|0�.��1b��Q�h�4A�Y%�<SE
�4w���\2��,�/p*/��MΖ��z�ִ����-�I��S�޵rWT���q
᷷�\�PSfF3���9[�ұ��3t��Ffa�+$�;/��VT�U��:�p#��ap�4�)��Mj�۝"�����: w+��rv�5��r���h���Q�v��%G�t�|	�\ �,�Nt|q�R�W��i�;g_�T����K<�j�v�W��]Gg���Q_��'y"Im���Y�g-�m�V�,�d
�i�1 ��J�,�(�`�V,��Y��D�g������L9�W�g+yVh�场��l��(�yD�2�ʄvnZa�1켙���J�5wbfro�<w:C��r�d͝,N�ny�
��HXi5	�8(/s��h&pڢ�H�O��3�����o��磌귕o���y��s��H<y6ԙ(H��Ykg*Պn�ٟd4���øe>f	CGtH=��7_�2v�*+4�o�����F-�����$�t�%��	��q�$>�%�;F�w�;��.0��p�Wv,�Q��q�J�we�ݰ=������|�Q��p�4Q�g����N\a�uM�E�6P&�#����|�W�RMSo ��K��J���O7.�i[�k����84-eՏCb�R�acұ�ԭ��LA�殑��m!0�*�sZ0C�+�!TGM���Aπ��G/�V�u���R|�3ٽ^�-U!}W]q��5qf�-�K�m%F�iB�6vpAuu�B�Aէ����Ҟ]��GJ37d����P�
ha�+�0��C8*�c�va2FEf��vեN��3�XX������WZ��:�fʋ�b�����>��O`�U(J	�3n�j�(�����yV�@8U-XHM١�P.����]|*|z������x{�z�������,�����"�5��P�N��*�\ k{��n�6�5��Fì�$��Ȕ1�#����^�
���#�{ێp���P{Q5څ�gn"��x#&����V�Ɣ�ӂV�
��G;+����ܡ���4��?{��hcc�Am䣧A�ؠi����X����@�xsb��Q�b�v��,EɆ���W��]�8	 ��P�
^�W�(���#~п�[���}��n����ݪ�v�@y��l_j��_X��m��]�0�Ruh'8N{���~�]�_���"� �;��<%�����o���y�ZP��u;��e!Rҋ0�%S-�ץk ʲ�8�_J������z��N��!�uv�m˦��b#���)��b��]�]x\��-a\Vgv�Z_
V���9�Ҹ� [���@��U�EZFDF����\Ѣ�������1�cn�x;��M!�����U�7#Y\�WU2��1�{��H� �n�(�b��$l�x|���(_8v�����o��&��y.�vƊ�ps&�.$�?o6�qҢ<�CT�tl���UW�t\�v���ȆYP�&�m��_��+�8Å�3ڭ!�@iq�U���t��0��Sw\�Y�J��t�tu'G���U�x�^�A�9sD�˒ں���n��Ԣ;$q�qu�9���~%ڃ��.���;{[��2Р��(�!�v�S���<�V3�n�+b` `�{�������Ew�� tWV)fn���8!4�һ�����N�u8tn��de�ul)�ޅs���!p�6.�=�ǀ��yQ����`#,��Ȃʣ+eD��)H��H�TF6�K"# ,��e�JK��A�P�/�g����ͮk����/�	B��k*��4���S��f�:{5=ܴ{��Dn*Y+*Ct�;U�u%ٵ����w�+�2μ&>�ɮ�\��q�h�ٷ��ĸm�{o�o"[����B��˻5ˬ��D��LS�v�4Or:��R��ު���+gm�tO`R���ˁY�w�/�qkh_S�L`m*�c5�u���1N��-�{��LW�ﾪ�^����_����c��K/qNG�`ۥ�n�t�Z�lĪ#,���_i,F_u覔��N�\�M�����~���I�N���Ϧ�EB��H�0U���n�{kUf��Ʃ
}| �6�A�
�0F�����~���E�Q����흚����zepb��Ye)w��5JW.�++�u��Fq8WZe���ʺSh^j����K����{�o��9�<��,���ᛖ�	R�%!�$�oj'c�o��=����|]��7�d�ӻ[�08��`�TP�]2KmiC�{E;���Qw=��S����/*p��ApF�NUs�V܋&.�[8��ָ,���f`�ˋ�c�gRp7m��_T4���S���+����!�!rg�t�:Wb"�Xע�Ȟ����PEe����Q�F�|��z��k�,�U}J�	�yݹQX�}��}G���6�C[����Νj���.�A�[k��]�U�+��q��0[$�t\J� �lq�W���  �1�x,`/:,>� �/
�SI�4t&뮸��yd81���(�Z3Wn�i���ǒû�9U6�� ��+����Uu�PD+�9�3�,���4�q�`�+1T�Ubr����{�8XB���_`�[�i4T�k��+B9ْ����{�b�����M���A��B�;:�f^k���]�80E��h�����K1��2V 7�]=|�kY������E0��ꯪ����j��6�qƩ��Յ;yD�l� ���FdR`�E������4@R��ݚ��tNd�mh���W���%�.���r��s�fE���ecƥwJ.����Gua�V��A��f����q�MA�c��q����V���pE�� V�����ޜ:�YF߽��V՗M�C;ǢP)qгN�����J��q;���ü2��(�E&GI�Y܂e!��tq�yS��Ӷv ����'wz`�|Qъ��!�#]M�G;��fp�L$;n�Z�Mg�tl�Pd�f�`s��o���{0&Wl7^G�I��sm�Z��"ˤ+C���~����Dl�"�K���,Xʪ�����y�*E��s�A�]9����:I�3ƀ��<U�ANd��7�|�@pcP��0QR�֌%3p[e%�(�����������95�byA�z�<<W�sP�[�� =*'nt�.,R���5p��-��M1 ��|n� 齡�_n�'/��)O������Q�g�[��� �LIU+!Y����}z��2���"�z򞙷���s5nH�u3��d�԰����R��堑�Bʜ��Hy[��u�u#O��v�N�[<��q� �T��1J�%t��[�(L��'r�퐾����S�
Q���qq�c���w���ezWoWv�t�S"X������-j���_fcE}�2j\�Y�d��c+2�̭��Ǳ�{�������kSJ��0p�$9��w,�*��D�����
0us]NEAO��r���,u�$Q��tWN�ˠ�C�J��8��m�������(s�3%��X�sZJ��u����QE���,�:ڤ�T"������_p����m륛�$ǀ��RXl��K�.F�O����ԫ�۹P�ʘ�o`[:;�/�1��Er�nDgGU�"�ԅ�^
%����$1�
�b۞է���Ğ�s���i2������-?x�d�}�n�� "
��R�����w�ky�6���ݑ)�|�(��{�*�!�<4�쁙ف�p���`7�,3���ٮ��{G[���k)�3���4@����W�(�У�p����:*4�,c� 6,x	��p�F�������Ĥ�N�4����j[�NZ �;:�3�i���(V���,Z�L(�ЦϢ�T��� ��� g�x�s�g�����pXr\��?I�6��>���"����Z���H��)W�|��Ѱ��=�e�K���؝
����llS�UUzb��Nl��ݜ��N���#2bC]@��1�{z�ޡ��>^癅���X��&>�ϋ��v���!-�~�g���3_���P��m����Vf��b�"����X��%����
���֜9Wt��i�-��#�f5vf��{�z3�\2;DY x{��E[���6�XQ'�d[6BY}Cc�S�=���c���Ð�c�ʛ:�6M!��N4�'Y^�����g����?K��_���5�����{؂�θ%Tf����G/��`Y7`櫴�w����
��G�m>u��(:�d���42�P�ܞ�]F�i��Mm���=�����~�$7v�j#"��-�X�t��W��óZ���ϵ�4�sLu���.�t��uĩ��W0S9�2;�Ћ�!�?������~jCA��0;�Tŗ�m�+mD����V��+ɞ���0�Y�a#Q���^7f��!�sZ̥絣�,������7`�y2R�6�*�^|B)�I��Z�OZ.1e(���zP慃B�MՄH�}A�b�I�P��F�B���gnR9ds�moijT��u�ח�U浚�t�Z�(������ý�����A�.�s�̣�듉]�Me.g�����g7��ǆp�&�������w�2���|� �$H�� ��21����""Ti-){�4.��+Q��`Qf�2��QW�΋'�f���(u����k۱�]h�J���5�
?&'K���\�P�rS�yr�v��ܷ�Mۮv�{�9UAHa�Z5b"*K����N\�y�Os�i�x�*zMp�j�Q�)	����/5�͖I����eٞ�z�c�e��P�O\3;Mx�w�����qs�ѯI>x�{�[��Jڦ�G��m���GV�s4����,�AR�v��]j�=�`�HY��P�P���*��J���<x�/FyA�
*�;G��)�5�z鳧��ڡ�J��IRNߺ��gޖb��i$���na��w'3�H��-IE�7 {�	�ۛ��\�u�k櫓L#�	X^VVZ�۽����u#n�xH�ͼ�}����˩��No����t���s��L�
�(]�QJ�Ƒ��<�4���|�Ź��ޚ�G[� ׁ�*n�&0��;��[� RCj�t6z���5�Q�,���ʶ]��ٽ{�寎�tf�̨�a��i�\����������5	��V�0��jD��}l�"�����[�s,�%�Ml����w��Z1�N>��wEs���mu�[�z�0�k{�LN��9�Z/��O�F%iu�dS��m,8q��k����VN��7��;y��q��c��f���=��n葡���+v�9!9�B-��WH����e7nR�2�Ư,���� �
~����C���k������ӡ�նS�z�w��N�X�p��۵���/on65��TP�H���.������T�P8�QP��n�C��(������nJ������j.=�Q��y��%����/f�Ȟ�&w�võ��vs��#1�6ټ��;�+9�yp���ڛP�"oU����tr\�i����� p]Qp鯟*�g7�$�\�����w�Z����E2��r��M�B�[�ݮ�+r�M�>�p"��G2\����no,�`�� �У|Dy%=���	����r���Y�����,�f.sB�CvYjX����I�c��@S�ux�qr�z�j���0�b��˛���N��ɷ,�ɲ����3^l��M�w�_��R~JÞ�M�|����ퟒs,�~����T?rͦ���
ɴ������
��+��L.��n��M&������V~g��k\��ؙ�{x!K��:@'��szQ�%&� �H�����@�Ο�T���t�0�5��1����!��Ю�~q�0��t�f2T_�p�W��l !'�`�/{����O�0��qgP��!�P]q�$Ӵ
�=�+4�2T��6�@�ߵ����
������~ְ3��|��ɧL��@�Si1���	��=�w_��߻�?�$��h(�O�RT�?3޺t���*k�'��׳��S�*M}f3䗔}��B�é�Cΐ��3��=eO�W�V,���?k���{���C�1�I~�c��S�i��S�4�L�+Ҙ�0�1��<�0?[�5���6��3�X|���*x�b*�$R!�DE�$X��H
,�"�"�b�F" �	"">���5�?�c�4�V���k^�����=�F�L|�Y:�2����>Vm��`�|�j
?3��]0�
��G�m�I���Θ?4�T�L��a�+0�t�i|ς Mt�>���V�ҍ0�1?3�cZE>�ɴ���f>@���
��O�$�*V
|��^��K�LLf�~!�����h?�1���d��M�a�����<_}����C��;�'�X|�P��P��>C�T֞d�P+�¥|�Rs�c�11�?1q0�?>gާ�8�$�gn?����v�����o:�R�N���|H�TB>@}'���q�Mg�L��&�_�VM����$�~f��@Ǩҿ�T��=�,�1�q1&e�����ֆ}ׅ��j���}�<Ͳ�{�������?%C�Wo�l�(w�d1L���ߴqMd�~!�1j
|�H|�3������%E��I���w��ത��A$�$��#i��������tEa�P�+t� X쑉Z�e��i�Ia�x��iN������ۋf���]��s��t"�8������ǵ���B�N��3�Вm���r�5�P����Y���I8�ow�'�����y%@ݤ�ȿ�O�﷐�T
�O�\a������*e{Z�����zb m8���O0�&0ǌug� ���d�N�Hq9�!��N{XI�O3���3I?0�i��~s�5|i�̝J�XVc
����V~@�LO�+*�v�}CL1
��@��q�?0���Èm?2VlP<���O���+��| �f��"�F (��1�$�C�bO�Ri'���u�B�v��ݡ{|�g䕟��i5�:��M0?��쐗Y�J��*(|��NT�2E�Y��^����]���<4����0�- �߾���˟�߯�߯�ME�!����Qף>�b����FkB*b�k��a`��AӨ�W���,QFa�d�ŻZuf���6A�P`s[F&;:�����)Dp�� 9[��Jkt�L���O�����u)1�}�E�eG/�0���5e�v��w"8�
 �Se�B�b���GUU�Տ��cފ���{��J�^�r=p,�gF�[�P:/}�f�^�4|
+(��c�Rʲ[,d���!,- �U#�*TH?jgKW1�ɺfa�V�v*-��s�m5�lƹ9[��㘻���F1�K�/x��^c�qeњ�1�x7x��Z%tQ[z:�xX�y2�nH�]��aUq7�gO$�~����x'���xR��q�=�_|'1t����3q!�>|�K�2��U|��(
�7�yo�\ۉp#2�s�Ua��Ξ(��Bx����}����9 o�3������T�$R�~�2]��k��@Vh5z~�:FD��ꯪ"�.�n�ڕ���v�Es��A���H�\Y���jy����͵}�,*e�Q�>�+�������Gƀt&��5��W�^'�`
�-ѝ���B%p����gS�
-_�y��˖u;�<4�� [�؍ǹ* �18�����6��I��j��s��D�Ӕ�<<=�X6��ʏd���5z�'
ځC)\ۨ8APT�ѱM#�v��r��9��3�8�(�%��ĭc�� ��]���������S���+𘬑�EG見�B�/�����w#`�����	^J�"%��m�.��,��Y����2S���N��K�}VM9�vN�����j�\�B����d��Tu�
��@���Z3N�I�����r������P��'e��z�b�;��ȍ���z.��ѭ2ZkG��k	B%�+svB�u����@	���K8}�����˹���UZ��q��X�8�62$��F��������D���A���۔hY+MP޵�+xn*��[PK4�9L����S���)g*�mf�5�:�������X�M���r�Ã�����f�x�Ţ�<:T��)Đ�ו�Jٹ-���P�Xm��\+��9ꪯ���xY��EJ {��M9�u�QWb��	f̀�P�g ����a��	�]��ys��r���f�t�trr��K�SO�����u��k:p�t��UWܢ��ޙÉԶJ>a�t�J��5�6e)L��,�K ������$X#r����}���}76�*�j��,7Ǫ��G��n��D.�����`u�rΑL���:�+!0wZ���cV^��[�9����1�����0)�=�K�����������e;����ۯWA����B�Wz�������{ؓ�c����vDlow�[r´�G�w�}�U}�X���r�[H�D/;runt��g���5��rt�y��}���y]�.Ws����2�xx	���Y��۔J�MG\���R��{�2��z�d�ԃ�鰝����)��=��$>���}�}����JX�Y�&��0�JmC���J
�X�����5��fi�ü�'k�$Q��v	7������OYY͕r�7���j�N��l��m��0�A�f���7��Μ�.�都v�),E[��_~�Ȫ1PV
"@AU�( �,TdQ"� �g)�ڷ�~�kp�Vٛ�!��������%#�Eq�b�#TX,�(#3)���#2&�N�fZ�o��̭߻���b=b�-�>*�ۺi![��s:��7�h�ktF�緵���;�wp��ݬ9��*��A��S�ɲj1���َOd�xo+������������tjԇ��&0�MRy��f�w{'U�� 9d�lΤ�Z$���&��f����z��9�z�����BYy��W�CZ�	�SG����(�tk\:}�=�ew�?,�b���J����"|�P���/����̦�u�)��ݾ�i��M�|J��*Y�'͙��v�غ��۬��&s��F��T�{�~���ʞJ��W��&��Nh)������<�+�m^�<l�Y�ea�#��b�~�(��ǚ�Q؋��Λ������c�]���O���.��K����.�����w�m�fDH�*[j*���ҵCI3�����|�>�C����N�J�{@0��#kw@�Hό�w3��ۄq��G1@��WY3�8pc3v���H�5����'��g���<��%q�\�gt�35.�Ӱ)��<S��
�
������p���gz���E�M���˺˼cv�N�?R��{��k#��voW-���Fu.�U��O`{�J��0N�Y���V$�%�qn�� �Bv���N;:�`r��q��L-��G�_}T �n�M��m����e��n,��W�Պ�GeG�T�����t]tǀ�� 6cds��t�	]�<Op�7�=����Z��j	󕤽��zm=]����$��ȝGk=��k�����X��y*�o��M����yP�8\�'���%g%kBm�2��}�*��(�@��]�h��r]�m9M;��Do7n�F�Tn!BGi�Nc�]�6�gnY�ҳ/L��n#YlE!�j��q\��sxIٵ�;Y���e*}�W�ꪯ��a]�T�[����k��|2ַۤj��1��S��u2�y������vc�����F��OL��K6�.���`���d籵�V?y����<fܯIY՜㻎o�u��jl)_pC����/��w��;�����s�u�	��5t����l�$ӏ�^9dز�]Q,x 'f�/x�U3��A����j�+d�!S&I
�
�� a�������6���qJp��*�;s�UWЖ�j���<OS�8��=�}9;��ֹ\��d��ۗNtҫ���̀�)߹�vsϷ��T�`1��_�̺�5��|9�7��82H��}DUT�JA�K���Z�����8�`;z���֫�(˨�3�]�d8��u�`��@�1O���Mś�ot��/����2��⼓���u�W�q��Ϻp�dR�SX�ƋϪ����'�*7$D��8  �����O���_^�����ă�}��)���t$ĝ[��HK�_X^��﮾�����\�<|�^Źs�I����y'n�=N��v��>j`�
�o-�=]7t��3N�^x{��������mX�7i�|��9WCzU��P���/C��R���e>���/"�s�a	&�,>h}�ā�E,�F�}u���>�ݿ��o���6l��mt�����\�L�Wzx�(��'UUf,<�kE��u�%��DD?���Mf�a��G$�j�� �'K�"B���Y�]�IM�79y��^ws�ߥÇ�dJ4�fR�bR�GQHX��q����d*�X�U+F�H��%a1�2�c M�!a��Ƞ�$ ��%)��0a!F 0�� ��h�+U+�j �%�L�R�MaAL��ff�ݸ�l��;
��I1S��z�bdZ��GiLJ�{�d�X�2�镎@�cy-w]K=5}� �Syʵ���Rތ��]�$�v�jc� d@��ړ��(�C|��q}ܡ�v�����{3M�]�kg}�y屩l�=�}�ǽ�?zK����~�v�nnK��8.�>�0ˊ8��S�/smP�y;N.�O7��leǴz��xy�y�B��y>�*��C��+�/�vJ�	�+w�M��\��_}�O��<�}��މ�"^������1��g�u�%OU�7�:AV +�
|�:����5�&� �a/9=vOގ_����� �G���C���뾆I�N�d��h����O]�6����[�x o*�W���xL݊��[�J�5JvY��q9��}��{���f�:����^�ݴ�����-|6mFj�l���;��G��񺅒6�L����A
(�+���WY�V�ˡ��mh����(��z�[2���VƔ�~�o8kE򙇤��77�ݦp��h3)l�4��46i���H\������( )�zM3\�Ղ�J�֥k�|��o���*���V��U���ե��wR����IH�bл��9w�o:;�}^����b�m�{��Y.�w5��w�����,+YE�w�ͣ�f�}��ue��N��(J[SZ��ʇv��DS��_��c��̧Ǻa�s���U�lR���*�ٮ��o��z�pϾ����	��TBH���`�5e-��(�P�/{��sf��R'[��z�@:^d�d���	Xv�P������8�y5�}֎"����j�	�{F}M�*#�M��:lTY	��Ѣ_y��겯g�:5pY�aw��|��J��Ǽ��޺���o�Ѳy�"�1�ϻ�4is��M��u�m����Wr��f5�e���*����w�gn�eY&딄�GqC^ O�4i�#U���!V.�r�i�����H�`�k�N4��1�#x�g6^N� �޲���j\
뎋�P���!wWZ~T>|*�P�lD�|:�Dv*�+��C�E]�pG�3�fA��]zG�m���3g3�i���
��*�jc�4i�A����9��}�����h�-ڭ�t���C��#��=7%�ƵcIJ��I9���$i4�կ��E�����i�徼&��x�Mrm�#�5/h.2�oĈe,[]�-Yۻi�q[�7*�!��ڻ���7�r��F_Ki�زvR�ኣ\�><�`���ΓO�O4]��;�7�j�==�S�^�v��m��Ֆ���ރ�E���ڛڇɛ�\��٪����X�����
ׂ��;P����G�|�l6\pCS�Z���w�7~ѻ�;ާ]R�G�B�<�:��e�y8���={�5-	A�i���=������XپY�f���b7v�Exz+n�"��U�nIKu"�f|���ot�܇��\�,���wmd{S�9ʙ�lJ|��I /;�y�]��E��K��_J�ŗ�<�ӡVh�JEq<�v�󏬴���wP"�T��kM�������N�#}�=X����d�.A��v��.�c]��yKW�z`��_f}y6`Qc�9֤Ȱ\W�dv�d5��m��j��+K�s��Ʒh��2�Ő��u�s��կ��0�:��6%VA{�w.��RYKK~G�y4.��N���)��KwWNp�Ms�!l���t��ܭ��L;��ɦJ[VF%7������a�)�(�5��-Bd"q�<�X�����9د�_Ρf�X�Z���אqz���I����A9.�5z-&���QL�H���;�@u�Ǆ�:���&c�,��M��̤H��qT��rk�Y��i�^����X�lBu�K皬Z
�;�y2ܗδê�on�����.��� �7�sC�u��'�Vu;�4I�Vi�.?G��ZBs$�}��B�Grz���=�ZOV��u;��]��,ߣ��4���꽚J���;�4u�?{�O�������xٚc��p�s����UݓB����T2ojxq�d-���qt_����@�,\���n'x���f�7 �]�'�G��y`/zHU��3/�VL_|�#r.tH���������n�A�u�]��?�\��Ś���qe�������ɾ�X�
������<C�տ}R�{�I�R���r��Cў<ԋ�\7��2�۸mnm�u�'��a�v�jM�8���C���M�j����[��6��+1
�10��K����X�*UH`�Eu���Um�ň�b3Q���DRk���������QE[j�"�i��4�e3z�ڋ�sL�8�F����c��\�Iy�5t��M���t�[X%�.=�;�ᴲ���6�z�Y�+*S��]k���wX�9�	E��7&N\9FӔ��e�g'r�{���
�L	���^��H�}���O^;�V��gEo��v^d�+{�+����ۮsV�7�GUd�K	�7_��������F��	�5{S�>=�}(�����:�����1wD�w&�����u�q������������l�鞩��L�D�A���vku:`a��z�q�����;$Ur�oY�TZZ:���� $c���
A$����z�awSN{w59����_s���Y�2:0C��XRL�gN�C�f�8�V����dq�y�8�}_}Y�i��e�^�B��XWE��|�M=�c���i%} ��#lT����}�.g�v{I���<pZ,m�b*R�kJ��17�k��{��;��J{ �4��ĳ1���l&��ء}�VI}[|���}U&{ꯩw����2;vqU��CQ��6j�ɜ^?�g���yBd�[��V��Q�����y��Q��b�)&��/�>���]@�����������띯�U*�7��12�7��_UUQ�A�Ǽ�o��֊��j0�8RS����|��N��gӹX�Mڼ���=��?�<<���4C�G���}6���/�,�I�"�:)&�X��y���Gd���@�uaΗ&�!O-;سS�"!i���`+wT����g��:�Nogb&A�����6b�蹽+�wQ�_Wպ
Rf�I�WV*�K��_3�^d�tr�ڎ��ˎ���q;���E-���D�Ȧ�ILs *J2�.\dDӤ�b��K0��0nJ��8�^��|��teA����>J�i�ul�Ń\�g^N�.P�`��̽�� �}�n�&��V�C���'��=}��;�&��mʇ3zdKy�	Gh�u�{���������Tnɹ�Knkz��(\��5�o���;����߂AeJ��v���k
�D}�E��V {�{��
������%K�Yr(�I0˗���b��Uv~N�1�!�ᒼA���o*~������!�[�.sB�X�����{}u������=/�X�-����}f'�U���< q���u�,i�I����'���޶2㜺.�{���uk�R䯾���ګ��BUURw��yy؛��w��6-��.M�2�;��$�&�p3��������H����_�s)�=���r�)l�j%�H�	
1eRH6Y����VFTKYKVR�)b*�*E�°(�T���A(�	d�DEU`)`ƴm)�7)h
�
w�ӒY�Z�z��{�!��!co�R���[SG"k.P 怑F56p�*3gU���#�V�..��Éf�B���X�R{�#�ˏK�2�zM����s��{��q��C�W&�;n�}_UK��Ӌk�m�ok��Y:˔��E�/�qV\Uyڒ�|����o3��e�����Α�tWx~��;���B��.i�]۩1�]䲕.�f9+:W���*Ai�f�lِ�Q/U|���>='�z���t�[����Ey�v����>�eڢ'��3� ��/UUTϫy_�b�~�lz��{:2��T!+��@;�ů����)�0n�Fn����\��:r'�W�{��{�����(�������PW��ьYɚ�3Ϭ�2�Ҡ����b�0kJ±rY�"��}��ӯ�[��W���k�m�@�]����<QsJ�\c8A�:j�f��,@��z(���|����s6���N�f�Kы*!7eL������U��5��ϧ�g�ݎc�p�'MRW.[(\�;d���{�p�Ub}��"o]���sg~�=f�B}�3z�tn;v룒���W��5.��s)?� ��\ݓ�s}�����k����Q����Ez��z������`ud852[)���t.s������nb���_v��=�cQ��W\Ǉ��xNo9������w���:ĸ��$���S������*^^ۺ�ގ\�]LF4�K��t�����vS�����+�=��꠻0��:�N��:��v�S';�;s�^�\�����M��3PG� �؛����b�c��uF=K�s����(���C���Wș��V�Nlܶ��i��$���{��f..(޵����K4Sɨ>�j�6�6d5�uR��N�x.�L��dG�a�!E�3�\�Q�9;k_S���1��vf�$����/w}��;�gٯ�
(+ ��� �,�TE�� I ��Qv����0f���Z�éu�ǣ5��7���͆3�rf�;L�4/�Z/�w���ʧ5Z�1s9�����Y�H�oW^Κ%<��:�KYSĦ
��,Ύ�P��Γ%C����&)�E��}�u�O>�נc�U�p�_(P.�����2䘷�%L��y���[X7۽}=��r,o�j`yx|����w*U�o���zzop��T�E,��]e���}����L�q9|潪��Ys�˵]�i��r������I
������a��vY��|��/���/9����"�"�*:��ǀ7٪[~)1�G+mLg��?s��Vˇ%��UZ��J�x)Mp|cC(S�oA�v_L�L�F�oV#W�Z�2ԧ�g��ECm��$W�������wl�Y�܋T��mMx5vmj�2��z�ӷ��d��ل�VB�)fg,�Y����D
�Q�����}AE�Qt�P��C�t˥s�v�]�Y��|_j//�!�4e�uZS*(�OJ��T+�� 8�������mu�u����fZ���쭇:�Ͷ�65y�s�R��mŚ��ᓞT��[y�>��7e�{�w!d�f:�b�3r>��_k�ٮ����z�I�z_.q�՗6'5v7g/8jW��U�ȹ.Cߺ�y��;��ݮ����x��[��ݟ=��-f��!��UU=W��}=�v4��\,�	;��f.$ԥ�Fg������>�ǡ�Z��DU�&���䣓���S%6Sk�fb��5W��=6[<� \��kOu�=u7Z�4{�m�ݽ��������7�Z,�c�|�β�f�$Z��ײ*4�;� ��{��y�!�������3rY��S;�J9X���&ٙV��}}ϭք�*��ae)�U�W���V�v�����:�N�.R�ts6l5,�A;�w12J�bs��];���8��Ͻ�����0��RB,I��c����<]��t�Z�z��7���X��u�ޓcc��v�{���܊~ w��+s�Y�ø��	�x1�gQ���sm�h.j�].�IW�egN��x�����Y������BM��wq�WKs[�Ns�vʖ���NRѓ�q��2vLXxi�ހD3z�MȾњ� }��=܌yuz�c�Ȁ P�ZF��i(�UZZ�cdR�1�c-�*%�V#!��Db[	D�VJ	`(�k,0��%��(��������_�}��@dsʢ������d�/TGoM=�n��re�T,a��H�
�fY�H_p����ι�P�$�N��S��o�O����8zd�v���|�rב�D����~�� �
 |'�|M[/aơa�Ӝydp.y7\����2H�mf�k���O+�zL�H������=mC��z��S�����@��}q�O5т��rԽy�3���'bh�up�:ol\�E��V���0{�4��FۮD	�B�&v�D�^X�Ev�Q�ᮥop}�tPH9�S��j����}^ �`�����[�#66��ƨ��:దdk�5;�Qa�of�z���r��]ܾ!ApHOG ��� P�  ��.�?A|ެm)�����6�]Ss�0�����i����^��L��7�]qg�`*9�jէ��$i�ؾ�H������U;����ªR��Ln��W��7Ƶ<�cqw�Mw�������*�z邛�@PV�hWR|��y% f|�44�����|�a����eݻ
�&X�DOf`����n���c���n	�md��V�K�*�FVs�٨)���M#Ӛu����:շC��DUN� 
�]���խ������n�u�c�D��5b��G[yxk'Z��{��$�I��D�딂Φ��>�}�vk��:Ƈ(Q`��W�sn��t�ʒ��w@�t0�R�-S��4���I ��֛U�s͞��Y@9yM�\�N|>���@���W41O����J����s���Z@@nS��4���h���s�=�ڈw:sFCl���5����⏳��}ܕw�oV�£��ᵉVe  P4.����#w�Q��&�C{�_S�*�+#���-Oi����i�/OVS�jGġ�UT��-���<N$뛫(����Y���Z8UV�!�F��P���̳I�L�[�Ӗ����4�Cv��1�7�'�3��\��/P���Qn�7#�Rˋ��|EI��q܎��:(�Я6��}�3�r��[��Z�9fH�:�Vڥ?�J��_[��{rº�{\l�lc͐h�Z"M�E^2��Cٮ^�M�N�=8���[(��m���-����3��pY��y�C�vk�}f2�s/w�U=�S0�LE��"�=VF�@y8���݂s١K�������$/q�xJ�o�@=���W�ek�j�y��H7�|���S��Vt]=c2:�V�*��z	���l��f�G��_$����>��ٌ��m��q����/m�1�:�t� Kd�l^�ۑ�:��w��QXɫ���I
�Kd8�r.����e��K�;k*s';��(r��h�\~;����/��)�7	 ���^��R[�G�����V�-X��E:Nr���a��#-Ib��H�F��
�f$�*��fC.tyGx\��ǽ�&N��p�;U7�s���m\�\��}�t���r���-�[�o�7�É��ќ���wD�e묏/��-��q�,ԕ���e�������Kxnq��h���\�:��aYc{o�>�Å��1}�fս�y��ڒ�>3^��pP�Ǯ��� Yrt�S�ٝ{�q_M���"E�ǒݳ�v�����Z����te���Xn�|���yz�k��t����mWeCh;]�jWZN��)�QZ�(�w�������]ݡO"��Ƙ��+[rk��v�ڳAAգ�iԡh@�X]�i�� ^LG���S�{�}��zVNN�T�\���n9���`�7n��]�ԓ��ʋ��{����N�� ���� �q	��N��詷e�j꛳zլ��EB���(�W:���`z$�8n�6�.�_g��[^�����|!}���Ƥ��V��3{�۝F����W�x��b������QD�no	q�k/�y}_WX���.�W�O-�N>#��; 盂h��8ɦ�Fus�|$���#wjRd���d.}����RVrF��%/77�|3�eG;6i�q��o��T�,"ys��OY�b{�7���Xx��ǀ����Y#wٰխ�l�a�K�&���h� }@}T�����-h�1 �"��fR�Vkf�\xN&�5�a��i\I1d�_p��BA�y\���,��h9h�Wc�����f8�������S�XNTrc���ΗQi㜎^��$�_z�g`���	��G1�jm��>��s*��Yj�L���m	�;�w�j�d�o�Jo�>�u4����S���[���}U~�~�S�+잸�	o��;qjkpj�QJS��/�꯾�����gE�A����=s�����et��R���	�ъ��k�tTpE�����0��纺_s�4�'R7��L�I��m��O�/�V ��"Ē��턞�]4�3�`����n�������U�u�A���,xC>��'**��Fީ��������z�N޾��s�V=U�V�O:=�$��so���?  � #E��E7���t�������HB�"��������2_L�s�^H�\$�$�h^5��{������'u5\t'��B�CX8W/�%���J��
�o}���,�S:G�z)awa���a��ӤY��n-��/����3�
P��Yɝ���8:?�课�.�=��^R�]��Ļ53�@�<�d��w�M��)ǒJQ2(�_A���w�_Q�ػ����!Txd�	+�!Y��Yn�5�}n�9Xp��;�C��T�t����U}�m�w�M�ƹ��7h�V�s�<k����g�s|�G:�����P�����w��Aֱhvԋ؈���E�׉�ꯪ~����ݢ ���5:8C����oMG%��w�ʛ��.f.�..��)^D��"
o��fY���	'�cB+ ��Η�w�����?8�o���J�-C��OAZ��������jq0a��>l�x����%B� XDB���bC)`�+-l�V�&��r��^��O�]�]s��M���H��i�4�K��S�ٹ[�K�S��;��zZ�D����O7�[I�7ж�U���PN�y<��Z9菢Ge��fg�E\�I���0�K56�I��/:j�y��s3�i
�I<�)a�.�����ǵ�q}Y�.��^�}SԽ��Š�Q�ڨ�@W^�e0���W>�����=�p��g����9������N[탬����;U[����j���a���8Սf�����%� w��\��~�O���=�s����/���a�4��649��a���Ͼ�����8O�iG���Kز�q����:���Q�2S�pT�6,+)Mj4Զ�ھ���%��7�/#S��sE����$�����L `��s����j�{�����(�;{�T�����Il��;̻j��2��e�13ll�%<.,'x�"�֜ٸz�:�f��I���""��#��l�>�_I�E�=����:�(�3���G�ʘ�e�p�	�d"�&2��E�K �na���Q��-QTh�R�2Z%Ɓ�L�&�0�fkY������5�L�<�@�*rO*m>���m��R�t�]�uBՁD���]����"D(7[Ҵq�ޠ�}��wP]$�%���H�H�GW%���C���l�΋�Ƅڐ<��w;!b�ƭg�"<xqD�c��Ԓ ��(�.b�{4c���H�'�/yocȰm�G���9��)�qS��u%��7�}��_��xw���g�cz%I�S8^�r�>��hPj9��, U-#ϯ�W�)�/o���ˌ����2�ٞ�,�Z�������c��`{�}8n0e7ɉh��p�]"9�,oa�|iˮ�Q\�<\�#X(��s�D��ݫ��&-qLE����G����_z�na��+�s�,�'R��u�w<�j�j�NU�a��eRh��|$�0���yp�� �P��/7�%^���U���za I=c(�{4�{:�|p��E���-ľ�X��c~ҳ�6��\��֨�E����U������ {_�O�����h �J�"��"�(� ��}T}��N�aѿ,S�g5��Q���[N)���x`���w����ɯ�Y8�ۃ�l��A�E�N
�f���F�ItVl�U	}M��m�IZ�ܛ�ܾ���j%�jgm�`�<��R{tص�OF'`fH�0���'S1<NS��3L�Ft-7B�&�1՛M���DW�W��'g��}�5���,l���p��| `8�St��%�Ә��6�yeuh=w١�Zw=�C(H�N��"^�h���^`�xL���%&��Ƕ����)��^4%���Ȋς5���EV���P�u�oWNWdg�������uew����`�H,��,�����]�R���\O�����e1,��$�3�oCA��R�5��ӕ^����
Ea�)��%7�͍����Twhk�E/}xe����b�I���wՠwp4���.@Bj�8R���O*��ꤾU��C{��Rk�t�z�!�:s<�Heo�@{n���S]}�.#��5��Q��Αl)�1�|�	M�U8��r$ J �	%;��p�I&BP�m�Z2]x�83�c]��Ť��V���w�e�[X���Op�씮ؚ�7h�ïmb�,�܄�{�n����Ngc�Ʋ�L��I���}�_;��lX���RA�وy�_W�v^>�F<�KRwB�'�*Yi²�	C�VOYθ�qIu� ��,���n�ʫ�-��b���T�""���I�@�(
�G�����s���	!�t{�)��]y)P.��t�sf�r�N�U��D�Z�X���?���KtEO~��z�
��3���!Q]�M�Փ&��=��ea����[�]���p���.fJ/w�}����[���7�Բu�'6)IN��\�g�����3S�8m��	m�PY�P��hV#��T� �B}D}�\����[˿M?��<'\���S[;un�j��ȽGB�D�C��F��8�-f�t+[�Z�Cs$"W�ܑ�M���>���i���f��r����|����F�b��,b�wr��r��>~S�\f��ev��� �E��0`w���_wW,��3�k��������*p�p�1M��*��C��o���knI�S30��(s�6_,���V:k�)Ј���n.�s��1���0��[�>��>��:�p��5R�H�]��`f�휗�l�&�Vސ�g,�������C6�9;oM���׸��}��b(H�,�a�/�����������6貄q�q���
���A���(�q���u������Y��Q����n��B��G��>��l����hH�%;ͪ�)�
�T�ꫧ)2f�(�\�j��I��q7/s/��ESw���y�*�,�t���������}#\�e��g�UNЩ����^s��Xd�,�l�С�P����zS7qW�R\��c��T�dB`�4�]�Ƕ2[&�`�}���Ut��X�<��z�.x���̎W/��L�v8���������·Bx���T����0��"q�e.SkJ���e�K̴���$YPĔ�kU�
R�T��0~����o��7EA��M�Ć�]���F㸅��A���&��-�JE��]�N�C��Z�o�o�XhKׇ/^�M���-6�:g%��DDf}�y�3���6sp��$Ui�Ry[U:�S��[�t�����y�eB
^iI��K���=&s~��+��>��g�����.%���'�R��o��V-Q�J������B�&�=���'��ڸx�����ӿDF���=^��f_�#>��]�!�O^Ss�&Fp���h��r��a�⺩�T��[\m�������s�er'zr1��H�D�
���G���gyD�z��T���97O^E췛:�/���vq�I���z��76����9\�o,���K[��d����o;�s^���c4~3*LοVMl��^���}�W6n��3����98�2݂5P}k,���)�F.8R%S������ʍ��~�Q�R�KC}������-�.�r��^`�3����}���|�����# � �2��IP�ui�8=��k��{nة\Ejy����1��Z`ܛe�!��#�c���)���ЖL;�;�-}cwS��-���`�ZZ\�Z�N\�6�#��Yn�z��Ӗ���_?������������^v�o�}��ry��惤����|h}���RAu�M��Cc*�-��w��_;�����{YJ�m�a���b"6c�3J%K�q�	�:���>��]�+v�S��^��6�t�n��	M��B��t3��gȈ�פΞHp�a���v.��,�{����{�lz�׬z����5\{�v	���mv�RS��^���0�D��5���J8p�酳F$��F�=���hz"3
<��$�'�d���:��F�u��C����_Z:z�΃&��sJ��3����3\]gU�.I}W��WG�}p�?�K�;}{��(��*��I��p�;(��S/��A.�OJm�_2ù�IL*��[F6�f��dc�Q�M/}����8�zQ���?E�%_|�͊�͡�]��a���2���
q��ԑ�kj΋\��>I�α����k(U�F����Σ������
��qRK]�6x��NƊ��WMa�s4�}��J��%],�L��-�c��hПd�߳�:�Qm�ƛb(��A튈6>��P��B�XNk�j��<��b���DC�Z}��h�R�}�M7T�z�{p���κ��4�J������d^�/�R���]h���bV�]����GK�b/���V ��(\�2O��� ��E�޸;-Me�E�,uJ�}�or�y�S�}lw��R滽틣�!&F ��`�S\��IdX�5h֌A`,�.�X"%�V1N��P�dQH��7� ��;�}�߷�桱*@����1�c8������mz�� k�~�m@A�ަ:�;��m��"��O�[����H)7U �-��Q�j$w��5��w�8�zͦ��q;�󯷯s}rv�b�r���f���e �KQͤ�a\/"��.�a��B;�R�#�״�V�����_v�/�U� FRz�r5��
�WY��Xj�Nj�2�z��ۧQ��n��7l���-������\�3:J2�[ڨ+*E ����{^����6ކ��I�~��wr��x^��ݧ+��5�PK�.T���򲊮OKV��@-c{} {��/�
͘��s��,%
�:U��i2{��b��V:<`P�#ɭNƷs�0�-�������$��+Hutv[�-N���d�z��#E�x�*}	�F�R�K�XD�]m�j�����w�:�#tAp�9{A������ �N����R����n��V-j"m�35�3��W\���i mr�kjK��J���*ꒁjY�nd����������C���l��ã9�b�-��G	�l�0��
E�<-t�Q����:Uj�=ݛ}�s'E*�ȯ8�fe�
IQq'�`3��3,�bԔv��wp:o%vC޻2%i{Lb�C�����-�S�Wڞ�����Z5��e͉I�$}{!�L����u�{�r���f���U�Y*�v�Y��Ѐ�=/8�-&��K
�dn"�f�.8ށ�{��Y���E�]J�clj�u0��n��h@}v��.���Vڸ'9N�5Y6vݥF�;�uuZ�S��4�P�me�P^�t�Z%�n�`&��֯e�)$r���]��p���ٽ,�i���L��N��Y3�֛�v�m�R�!�%hY����{MnG)F*��s%�ZÀmc->��c��y*\f^�7��pI�t�&Vm�՝��*ox\�����ad�ړ�xun�+�ڨ�aG9�D�ᡛ뱼@%Y�!+�*)YC*X���nU�Ҳ��e�#�NOty����F=zx���������L�:KѽS}9��7J����:�B1J�?}��k��	~ ��V�UL�"E֑/�Uu=�B�L4Ƨ�%7Y�\�;�zt7��Og�����NF"����k�����ϡ��E� ������^�н�;�|ƍ��Ŗ+%rN����ޭ�A�3�-�}3ւd{��4��`�>�k*�F��菼\}��@o����������E1�!��S�`�2�6�E!��gq%쩮�D�ng�nݏ?ግ"���9uS_C�������xe��>��2}X��)G[�%�-K9vvW _yu��K�rU���-���r����^�8T�Gސ㴟�?D�3�($R""O�g}��y�?������Y���L]�M6�C���Y<C������N�Q-l�2V;,4��_C�����¡X,%
Xw�}��{�x�m�Nܭ���[԰�j��p��x�36]I!�ī������Ep3�؁��,�۸5��Ɂ
2��tn^�Y�|�m� W�#�P�|*��8��·�QR:n8�>:�J%FO�����l�҅�=�_�>��VO7Ǵ\ubbI1���r^�NOG��C�-�I��xO�����፹˭�dps��	'��9T�L�)�0��X�8%kn��-9�O̇�R����� �3��x�uo���I�	Q0���D�FqN�CgtOZuy��罳��bX*$Xq=(c�'yR"Q�z��>���}�W1�=>O��Fmw����R�A�;�	9� ��6��N����װc����De�W��
d��#�l���tnk��p)I�5Y`��T�\�fUP���b�T��/��2�4 �S;΢�
m�2@�=W=��}wu�zN�/�-��O1ﾍ�ڿ6=��B�\4~@����������bJ��IX[@� ,�`! �O��F7�Ler阣@ّ�r{��F���U��JՏ�;B���ε]u[��(UypE�ʡ"|{�f��!.}7,�-�
X�Wm>�W�t�l�<������<�N��ݸ�H�KoV��	��-���eW���sz��އ^��̹��W��V�<�#r�h������NQ)�Jv�J�5��-Gq�빬��dY��6�G�Rd���>V���o��|-~�.f�ԧ��~ԏ��F�U:c:�p��^[�ncC���e��Pz=lE�6)FU�,n*�K����K��V:�\M�Oz>���|�&;#z�G�ۨz���'�L�z%�c��|���3���9٢��Զb)I�WX��z�����g.��{��}w���2)� �?IW�)X~WQ��75jR󨥢�XPh���=\�ht��.Ii�:�td'TU��˒����-Y�uC�Ս�H�cˋ\� j���qł~LZIfV�<�Bg(��<�N&��Ѻ�U�0��v[�&k`ȌZ¥���-�ق���9>�����Ý��jA]҉̸���$!H2A�H2A	"U�A��&e��%���k�3��3�U�B�2G�L7^�m�[:��p��WҬ���jlˮ��Z��է�tAsY���wر�X�֫��|�廸�i�۽CՇR��yL���$�:�.@C�	bp�E#y��q�gV{��t�n(�3��s^p-��>��'��Hx��������%n���v���ǹ9�f/v�]�qf���踑���.��;*������<���"5[�BҺ����7��������{��3����`^�,�*$xtP��i��ڛ��\wF�x1�WO'�Sq��-�k� L5+D�"9?����ݥx@�A�O�����X�yMp{&�<��_������;š����	�UK��x&���s덂o����$w�K_g{G=C�"M�Qm�v�ˇk���Ӛ.]����+˥z�r�HLX�B��G�aD��2-Yl7J���}{�c�g[��Ν��.nt��p+�&�a3�'L��Ψʥ���Ntul����ɻm��e�l��Ȳ@Ȓ
 �˳	S X�(T���[wu�ꎅ�m���;{YR�īos8j�%�6˴�hy�N.v�fH�:�}r�]�YA�c�(�2���+6Ac�d�ʯ1R�=�+�M��g�$��p���Y!��	Rg�����ڿ\���<�ȗt�����V�Ų�b=5�I'X`hҾBgF���]Q:����tٳ�d+�Ϊ(-�R}�|wb�[��(�?����Vk#��vY��=��k�.�����Ay{3�^�ײ*�C�.�z/�@�|/�v;z�<̰�_�{��`���D��s���i�����~��	���d�ǰѡ�Ͷ���zp���\�R9c�+v(^Γo2�xG�w�G� �.~��A�l��f�Й[ ������SeI�1 �vS��:�p�UoWŉE�ne�D��W��׈~�c�*��~X�_��/{��dRc���Q���(���XsR�j���r�$��"�M��u�c�at�eVM��T�����\�|�z�`���=G��1�m�0P��
�+�	T�B���X$Ƙ��v؂Q�(�)%�n��+��٪��(op�"�B��
�>Wce��rm���&Y\۰�M�2�:�Ǳr�.�x({=���v��%��U'����f�74�˩�6���9��$rS�+��J�����#�?A��z�xu����f3歃�k���@���;Bi�[�e�@�,�(���?��/�qO���G�l��4�F�۾�����8��A=+��
%��8����\�4�#�<Cc��������2�7�FF���qt��?gXl��4��2�Ŏ�
�	 q���ĻWޭ��_�����A���M�g��+��b)B=>��?G�G�����>�g��z^�
�iy7m��]�T!6rev+L;���3o"H�^�;�Ǝ��v�i)tDl*���G�/�	��
�����.���X��:*�&g�Օ��W;�Z�l�{Hz�K�����x7�9�O��犉*9�q�������������Dƌ�lF�S��_>Û�>��!�K����7>�0U�k��(;¸�a\ق2MXчkf��O���dӂ���7դ^SOS[+��>�<���p�/��t�2S2B��aG��V���=�����xvɺ/T�XK�mto�/U��BE*{_~x�<<H�$ r����Q�[߯�������U��9����L���z�-�&Jd�@z��m�g\��3b�K�n��W�Q�\�Τ�]Ͼ�_G���wU�ɓ��ԵS�W.��xC�@����)%XGi��ʓ�ۋ��ʘ[}��n7C-��v6�Ȭ����4����s��y��Z!���C�b�c���٩��#�*r�u��#KK��9��˽U)���H�� �O_3�b��Ι��)z �>x���;5>�g�=�8�v%v�R�x�Y���q�/���.fL*����Z����舏Gє����zȞ}�Ҫh����p`����Y��9��ƥ�]׃#�>>��/#���Qm���
����N���Y�W����W9���狒{���lb�\��2�����L��jT���ވ,��}��������uF7"���)q,�b�1&�=��>����O��ȉ+�+��<Ƭ�`z4[�
���<��|���(�Pԫ���s��׾�����,��S��W&�lI�r�ϣ�<0����0��qY�
�t�梇-�}���bi�4�q����4�(	�B�z��,9-nt'�"���V�g#����N��X���a�s�-i���fS�=���u�v��2�a�����l�`'����ɔ˛�H@��w����E	��(P�Dp��LM������m�g\gI�6{&�W���a/�nԏZU��Eqv��3U�����:��j�Ǣ"�y F}�9ڽ�{�y�������h&N�j�碌*S¬�z5M�w�S'1��f�K��;lNʳ��������_��`�$R"������n������g�[��r@X�m�)�
F�`2,!@VB��T�("d�1�(2"2F(�0��Vؖ�߾����Y�S�o����ٗ��p��fE�(qͭ�1��Gb�ofc���m��WR�Y]W�L�Q� �ζ�Ź����� j�1��i�v!k��	�͡} �+6��w���=�x��s�SxLF�iOE�l9�����}�t}\ǥ�۪�����c#7���(��R��dA8�;x��=1�a��P���\^��72t��������`_�@�k��Gߥn� ��f�:<�
�����R*�h�z�ZZ�H,qG.�ʮNA��Y���}��^�菣�Y�[�](�⽴�����)���^�$Ë��Rzԅ��V��O����r�Bf�@�!�+F'ԢL�~��q�����(9Ć|z����s9��<[��E�s��F^a_����A��r�;�Q�	��D�/�[�o�@�q^�L۽�bœ���Ȝmw!�_�oH��Z�Oy����I�h��j���g7�|sIF���
=����U��IiH�.^��i������GG_I#{�>ILg�6f&�Τط !*�7��C��D�S=�"�>���YN^����Ob\kn1J���ˢ��|R�9+��E��tFp�G����}�R!G9}���Y@i� (�ܒ�z7S��^�o�3��A|*#菣^� J�u7�К�k��MMG���-4I3�<����� .��̛��&v<��g$7�y�����ž55z����p�1"}�[�t����X ��ٶ��!�s҆�\e�h\�]���y�ev�O1�P��Q;yR/)`g%��|�6���T��-�G�G�ᬻ۲���1�M@�hO���=W����i{�!��q2[�s\��i��[�uE��� {�(US�����k�����?�,'����os����2lW��r��L)�	A��䡡_}UU���:�;��ǎ?��~����w���x�����pǞ�Pg.�=�.)A�ƗE��ʁ��eVh�>/OT&� ���̫rU]|ξ69m�j#��]
F%(X����>���y�K�sR����P b��"Y�I���r�bF��|A���3-��d����
���Y�|+h.�i�u�P4h� �[m%�qތ�k�qcp�V�"%y�9�i��q�4Su)mm����8���j�՗��T�����J���[�+H�|�]��[֊��nS��pFq����X>�D]	�ok*��ʣM��" �Xb�e�c�*o<�_}��n��"[�\.M]Nsx^����x��Zr� �sT�,����sW3Z.Mi�Z��������ΥKep��iE��QU�Y��uȉ��40�2�3��jb����0�朩��1;�f��rce$X��L��N����p�>͗_r����3�I�mp�� Y.�J���ί�NN9I�xe�]q��ܩln��]͢�a٫��tE@��(e>;o�T��o���W%�:��Z�麗[���?rk�jnX�:�������}��ô���d��c.Am޴�U�9�d��߄�giP���p4�Gi"'�ǲ�Vq\si	��hPV���wB�qS���n-¯�96f����ݷr�bRhA�9��K7V��zm.��ȷj�����:�;:�ҨMA�>\�������S�ɨ�R��[��N=ݎ|]�����V�m�Nw�P���ɳr��K��/�ē����v�w �n��g�x����ڄ۹x1��=�_I�n>�\�ٱ2~	�c�:
�'��R�W��wG����D��΃��[�vru�D�Z�M]�KQf#ӱ�L��ѫ�����_5h�᠜oW<����9�d�yC�%�����:��-RQq@s�vgB�ѳo�]�}LKR�eu휻���(��Q��v���ZlQ�k�*����5��ǒ�t�wch��%v�ʴ��[���t,�g1�����W��%5��Z�Ӝ�h�9��	���<44���}/���W
N��O���*�Q�X͙�:U����y�n��.���F=\xf�Gjoj��)K/���:s��`�cs2�����R�u*N����T�5��]Q����F��W��'�i���B�p�4��e��B��M�]�S��Sva��.Iv={�W]B��1Ńx�|�Ѡ��u	�[�hnj;Y]�:��Á�LwFs�g�a�}�Fw9��m	�MqK(�;��.q,�n��G��s���Ŏ1؋[��l책[�/Y����Y�
i:�:-;�b,���;טM�a���V9�j�W���*.F!+���N_Z�TO
�Z<��GPޛw2��eJ��c(0�)Dm^ݪۉ��iM�����A��@>V�m���J ~�yF�<ڤ{_��
�̏���A$��v�Oﾸs��HW�^>/���"a��0Ks!�(w��A�7Xl�Sv�.��j;"ᣋq��ƨLN9$M𘔞�D��棉V;�׾��z7�G4S�s�W\�����K9NT�: `���}2���\.ף������w,���D��:-Y�3 �`dD|��{�sRS� D>99s���B`9�ɞ'f`�ͪ��ԩA:r�j�vq
��\%3$Z����)�(�ݫ*l��䝔�ш��6��}e�cU�>���
&��ױ*��3�>��L���T��k}��a�m�xm�`u u�_	�ϣb+{�ߣ|�GV
v&�ٞ����\���u)�x�3������]���7�-�'|=�iC���� ��҆.נ�����qG�V�N�=�T\O(�D�X�m���(�.cL�~�I�nţ�K]�Y�����N�y�{EQA��f�b��ol&��޴������<���Y�f�دZ�r�V��\z�Ǐ�WN�T�w![�ќJ� �g'��7�a����vQ/)�bf����a�vu�v��l��+r�h؎��=���<(:�/�]�{_Gʎ�e7YaK(\��Qt�o^�b���i�E��V2�e[�����;6c���l�B/(ODuz"��z]�[��9�u��zX���7������9y~��"P�R)�����
U��r9wsL2-���ⶫMkL�y���ﾯ����ԛ� <?:*�����o��\�� �m:��K9f�׊q�LF��3�n�p#l9q7(31�y�}�o��FZ��{=:hu�S.��r�8祐/y�Y�@�� ;FkC�zm��Rr��V�oF쌕�ia�Fݨ�[��ﾓ~�UxA�c(�ǂw��M����څf��1�Ԉƻ/�)�|�G>S��XP�Ϙhq�"�A\�d�E X��LRQ/��׻+z�4�P��D�����m��,�c1����ȯQ����,΂�ws)J�g�8eu���G��G�8<���:���Q�����5�s�z����u9�ʠ�ζ�MBzՙ���U�U�s"Ί����{���(K&Tf���V���u�V�sYP�d�'N�7���q*9}	�wTr�'*���f�n�og�����Ar�'�1��PJ��J����D��j�V���rG��E�>��V>�)���8���EL۩/nqL)�[]6	���0�v��C��yݹ���QJ�X���Nf��r���J�9]G�D�g�G����9v��1�n���WP��\�����x:�Nn2��Ӳ�S����9��|���a�5��v�0;�cX��=��і\X���zC#P�J�+�2:�T�i��{kG"�Da�!��Z�Ym^8�����D�˲+��ֺ�-��_?�T�A��x?�R@9��4���~<��-�"#�Z$�Wa�mP�1��1B� �h�@PLI��[0��H�E$pe(�2�
��*[3�Y"��f�?Q���J9�Օ�yoz�4�{+_c�/�^��:�6���}��b��f�ى�(�t��c{VaN�\:Z���W6�vҵ2����nH�ӏ�f����>�<���먆L��w� S:�z~��Q��ѽq2�3�>��w�;�^;$8T�%,T����FȺ�+K}�nW	y������2Ulu��=�8{n�KF(�O�G��ؕ+Ş��+�'��1<��r@��(���k�$�T61���b��2���
��jM��L��q;��W��o�W��4�ٸ�����v)Qާ�0��u��'A�I	N�]O���R��^��8����eO0ܗW�z"$���t禉-a���}��e�(Z��qR�oӦ��URg�B�q���F��Ũ�ꯈ����Ce*&t_�>�m�)#����a2��N'R�Zq�.n[��+����a;�Ї��{���v��z�O��f����"&D�1փZ��X""�2"ŐD�Z����>���������^��z���g#嫔g�d,s�i�+�u��q������#����q�<r���ۤ2��.5(�K�]CX�+`C����Y;U���8�^ڇ��n���ƭ��tt=WY����2�h�
���~�(�
(T�^�}�5�^����JK��r��mF�ef�ඏP��F��$�Qͷ/�:�wpB�e�s�<jU�T�U�5���*�w&�E�e3�;1�\���m-K^��Y�s|J<�9.�U�0��p�K��sp�$�� g�X��s�!5I��S������RWp?���0��E���������Y�\s��o3�7]U�P�(����]S�ؤ�d����ٶ���ON�ɷ�={�6i��L23���%33(p�GAE
Eb-D��ڼ�M��{|=7xҖԗɚ����{Q&���q�����(^���g�V�5�Ļ�.�dO[+C���+WPB��1m�@���9�wO�Ȍ����E���,�����X:%n�!7+-��8�Ζ�wt�������į!lG�����*��63�B�7��YL@GE�)�7w�ܓ�_�̑X��{��ksdfi-��rۿ��O�3D}�=��~1��d��}��k]��U��e6�f0�n��ޚ�1۩ۚN{s.Zf{M*!�*-��z9��Uع<Nu=��}zfc���u�ߴj��X�d��XY�x�|3׮�p�B�q�D�̻� ��N�Ƌ�[ĭ4h�ھ����Y�^�D�ۭ�>���}�s@j���-�1�4ǅk��֘��+oZ�Q�B=���w�۝����9�l�����K璼�ӯN�jXÔe��2�Ӿ`�h�
�.Nn���`h4�~9����z��X��8d�<B��f�2��Gֿ}K�˟]�}�X�<���W�Y�vT�'��Zd�G�dIe��SҤƜ��Hj�=��E(4���J�C4HK��>���R����?f����{\u��$uJ�B�d#$Y�dO�*H�+`93Fi`��k[����9�~2�Mt޻�w����d������c���S	T��)�T��"�xަ�S���*^����:z�����#�4��Y���[/)訶���\kf��<r�����Q����:d��ꎮ��r�{�``ze ����K�NӋx�G�V,#�\���������}W:�ݢ["��v@�#ﮬ�Mk�N1��Z�>��5�El����n1e�[s�[�|���� ��W"���i;�쎕,�S������/O\+3�Gw����S�}�|���U���$��`�0��'��Y��B�SN�`$�m�sE�{���s�=n2�(�,q�O{i�;��u��\�ʚӀ��/EH��[H'U��q.���u<��qt�F�`���D�	���=Ml�}��qs�L?w�3�}LL}�^�~���fizw9&e�9~��߃��t}]r���ĎYjf6`e�:J���J��m��;y���"��h�LW��$���Tr%�&V�[��F8R[^�����[���uK��/~�y�<<%�R�oXVˊ��Q�7}����$ì�݁����rmF�;\�-� �l���o�YĻpU���:>��E-(w��
�����Z�˝L��OM�Ğ�n��I�v޸0�x�:Q�!�N"rJ�{�e ��"�������6�z��i�S�
���|/���h�h�r1��p�"���5-�/���Noa��+%��f:qi��8���0}G�5�=��r��`i��W�g=�؉�囉��'���泂%rinxK�pطJ\Ũ7��a)�$�U���#��zz}���	O�tVs�����_uLS�.ے^���o��jZ��]�kL�r���:���0�n����Pe:.]�_�*_��ɟ?]=j'�0hY�*���]Nvv��u���ҝ�d�,Р��T�%\n&����P�Np�ҽ'^�!�j|��)6M)'��R��l؉ɋ�"ȁ Th�)ie
(�VDID�
��`0F�V3���U�k;=K�U�lV<,��O*j�u㱟��z�]r'�&z���էE�C��K.CZi�T�{P[��s4�P��R*�Ǜ�8�~�P���_x�s�A�Sd�n$w3E�g>���_���v�5����Ԍ�G������t�7�oL�X�rH=�\�C5�>�C~��'"��OC�κ�E�-u䝴�hs����.���gk�ܡ^�Rs��=�l��u�챰�*���R���p�=��s�*UL*%�5DDae���݃\�Y��=�*���{3H���l��=�?U1$zg��u/��=pWTU_�j!ю�kVM����<|��{ّ���UU�v�Rw��7�/����G��'��YW�<�'S��$wn�B.�����Y����k��d�eӇ]��ݩ0+L�ަ����:T�����@mֽ�N��^�22{�\2l)������B����Χ� �zSS}Qz��`ul�q�"�@o7=
����~�9�/߿�����oa�6ֲVV)�-a�Ծ�hR&��y����eky��ZW�k��re�v���@�m\�-U�k�RyF˼r�K���O�m�om����2SJ_*˰��6�H8�d���QN��ٜ��uD.9)㸑�n�eґ�Eh]fwk�m�`V��;�%2܋d��3�#�g LL���ϲ�ɉ�	P�.��]�OK����\R@�k�	p���CB$�"�l�v���.���K�Hh9{}��>�{�e��u�S��� �1�ű����e���bo��W��"�k��:�3)q�N3e$�<p$ ��k���i�fN�z��=rb�fY���yn�_^ћH΂��Q�1W�M73�j�K�J��q�8nF5[##
�X�3j��]�5舶?*��~0=�q~:�\�V�T��ZǇ�������\�5��L%^Ng���=3��0�B��.�YS֫����}���(9���uz��t�s!)��&J��;C�Y�w�K������\�J�̗OgG��>�U=�@��$ȝp��u��U!ޑ�x@P��T�P��Ŕ퐑�6��l�Q)��ԃh��Z���~bP/>0e�d��wX�*j��6�m��E�$Am�N�'݉�s�n���!&Z�aV5!EjR�F��5�Af����6s�ܴ�bf��w�H�:L�+`�q��+���ID-��ѡ�b*�)��Zֳj�gN�Nz�r:q�(%�ѡ,�Q�ݼ�{Q�54o��=w�\�)Y`֪�u��gy_��@N��j	��ɜu�e�*�]�����^f�d��)�I�Г|��)���@��,,J�..ƎKޚ�hJh�4eh�M_%�j�;�x��\~/��8�"�[q
��B`���-��0%4!�o3M��2�}w��0�[�E�;8A@�ra	XB���^�M�l�ݹ���R�9LЋ;�࢓)[l���`����O�}~�g���������8؂����z�r��y�^g5f����"͛G`[D�j����RR�r�������dfUUi7��!�^+@J�gO��B��n��{�o�$s�-�	{u�;�L�We̤`�csʫ�"��O����%L�..u�f���x �V�����b�ڒQ��n�9��X��urZņ0H棙�D���x2aP�;��l���{�� ��M�DwD왹0�}#�:��K�`�����孖&^h��qxV�Y�9�ᤗ\�U��Z����Ě�:�t
�y[��ʒ�A�Us�6���e;D���e'3��2]�۫�']�������tn]��"b�w{���u���:��ļmB�u'+�
"v�_I�ESV
V�&�J4ej<>�X�.t3��GJ�@�l��v�[�Cw|1[{�s�O����9N�]Z�,T�ׇ�I��,�Φ�U��ˌ(,QM�gK����	ʢ<��D�p��j��n���P IVbb���*&�Y�즹"oZ�2�"��h3{+2Ȱ��t�V��k�ev@�|�m�
��{�3��uz�w]}���e_x�Ӝ�ۣ3��������+\b��2_C�+�S��y�S8
f�
���t7�r�K�́�]v`s��I�+F�뷚e�R�v�xyۮ��٤mte�EgL��f�u�i�܋�b�/^XUx�zuä��V$�9�/I�ۮ��J�ք(�',Q�b�7/lk�ltt2�WY�C��X]3ِ���z�L��Zq���&��f^�nm�;H����cB��@v-٣��2���2�e������Z =������%a<ku�t�2�~�'������������XE�'q#w��� ��N�*)6�Z!��١�=�RwG�٘�p� �v	6�I��vЮ��Q�u����9Y�7]�O#<U��Ә���F�Q&]L�k��ܵd��Q9�1��N�U#U�z��xǵ����ʜ�E�q&o:.�Ev>l]^�{.��S`8�P��GZy�d*q�jm23v�yΤ�b)㧁nE���C�R��3�dO`ȖȪ�:�<��j-CU�<��m�R{2)�3Y��DX�lJ���j��P��僖|�{��8�x^�=���]�����z�H����9����瘱�l.�9�&ĳ�ȞMNh�6���X�޾8�L�����|���&���	^P/�d�5�C�3"���f�s��G3�̘��u��,��e˕K�ŗ+����YBp�4O{�Hz~�f���Z[3̀������Z��*`�'�]�
����&nk���n��{�$�U���U� '3�L���(K�&_�G�\ݹӮ���v�jbb&&g�j�8��b�P����߶��ި^�o�]^�S��2�����S��ͯ_�l��]���je�\�e��g2�̡.�]�����)���8��K^g1;��jw�W>�ڟ����>��H��'h�FÊ1�gN׀��qu.ﮖN̯�򭒰xً���D��A���lX��Y����ܧ��<9+�.�{f7�Z(q���5�ro������ ��wV������(Oմ�5dٻ2Y�;s���]W����=٩�j�Nv_Y3iI᰺��0!�T��E�x��sc׏)[�`}}�t����W ��[����U�TG�/a�DOrT��P?��7��)����A��������"7�`umm�'@���}#�m|GLv
�6��3&��v��#5�=�4:�T����[��ɚ�p�v�s���f���6�&2]o'	��B%���!�����5�l��aR&k�t�9�Kh�㮘u���]{�����U��T��X ��b�C�3Yu�R1QT��ʬ�\�Tb�e	���b*D�IE-��Fbb!�_%@�9�5����Km����8-uN���="����7fHV��b�ٺv���-xdKoU������a��c�0�*5g�\=�]^;�@�ӯ�)�@�l�P֧���>�!'�̫���(n�#(� Xٙ�8Yz>��>�D��sf��Ɍ����ﲵ+̯8�$�s��k-��N�S*����A�Ko&J�n�8�}�z%�ػ��h����W���S��uUP�G��Ը��"]y�n��jp�{��D�k-fĄ�6�հ���7�.�q<�Bv޹����.�vm )7�������2���������,�=���f�'i���y��%�u%]�����l�w�Ve�2����?L-�WH>�}?�,��ju�^�A��ur�Bʾdv�T)���y��7�j�:d��`qb�]/�j�/��->�>�腵H�xﾏ�O_�_���{R�᥾&QwP�;�)U�����gň�)[%`�PQe�� �7tj�v��MS�	Y��'l�U�p����;��9��	tFcX���cf�t�^N�c%jVn����TsN���5��k'r�ޥ���z����u�WQ-�5ȶͺ�o����fp��Q^�N*y�M�jlȝ1ՑP[\�3G���?!ǆr��f;��Ýk���\_e�:���\{�Ͼ>��@�yByʬ���s�:p��8�6���}�A�;|�i��x�d8�-b�1a*قw��6�:Z'��Z!�Gޘ����5�ӑ��D���Ʋ���g��#�gӵ��|�~O@az�Jy~��dT�H|�c��<b	�O�E�Z����G���)�ޏn�R�jrs���x�+�Л9�!�<�p �GJ�.�䭦y�bK��XL5���y}.P��x�D}�G��=��7�m.�fu��o�%��1a�d8
��諥��ys͞�)���p�__]7�+6r��uXj_�s�  d��j�>ɱ�7;K�,���	�$z���Çx��c��vn]"��r�N�����m�������.Ɏ��5�j��op�lk�f)���qr��|w�!������2��@9[��ܞ�	�蚖���;���E�+Y؈ݲ��W2�Z��;���C~�������I�����l/�ֺ5Q����p�M���<w��q��̈q�q�m�fTWd�C6v���>�����n^gxuo�F�T�:�5iq5nL��X�:/�!S�WCB�p;���"{vӌ��h:G2�lO;C�Ku.���ȝ)ס��H
9��׼�p��z��tX����1Q��-�P�n�]ƥy��U��=M2��/y�n��7Ik;�g&���>�&.��< �'�UT��Ĝ^vj�zmAvsRz�'�fv`¦�7��F�o&`�⍧B�ww�X�ӳ�Y�8���1���N���&��+e�u�����w������w�[�˦Ghۮ닚H�h�������F(�/-0�����*�VQ��m��6Z0UUS2"�-j�Qb�����%x�P)"|*3��
Gq"��l�:ƺ�l�݉-�*s��~ưٳ89[-J�)ۛn�eϬm�n����kT��k΃�u�l�Ox�x���݀�[e3�e�G��a�t�J�y���2�%P5�:���n}�}�`鮙���7�dv�*�E�R#;y��ɪ_�TG�DuC�k}�6J���Z ���L��(8!�;$���R���V�;�+byاv(��l�eL��.z:e���o�Y~U��;Δ��q�����+�
����9r=<�{���h��k�C�S�z�^f�U�&7�W����g��z'�ʆ7Ī4�UG�]fh
龺Q�U9�Ud��	�܊/��0.���qu�UU�U��Y���Y�.�>��G�Dd��P[�0;��tp�.g��h�+������G�Z$��}eS;�xW���E��e6�_{3����+�W��I	l�W�P�\,�R�(ɨg�-2�Y�ͫ�5�}�g�� d$b@D�d�	~�f?n��q7O��i����tr��lH�ca����.���Ý,損��(6L�]��]4\�)mVʢl�E(�HK5.��	D���r��a�u���4�̧7��
)��%�t���%��^�%I{9���(�Be)n����p��2�N��=��{��o"�FDt*��ئ��^�<7�{�鬢��m�w"@)��זDr�E�f�H�&L�+�)[���!�s�mk�i�Mgu���ÉHl�N(�=Q��}�����S�C�z������ښqN�v5����|�J7�ǁ @���w<��g�]�� `�G�Υ��*��^��1pHvtXg1��� =(%Н$v���j7�4��l_ c�t�H�4��n6�S�=3	�b������w���n��m$.���ޫZ�U@6�U��r�sQ���h����\��힩����v�i}�2�z7^���#�5�]��'�l��u�J�����)�`�ie�m�J���*E�X�	��a�0$�.Z,�Ȃ #X�¨[F����*j�fI����缼�%Ծ�<H�L�)jF���]�7:�Vo�Pe�ke��wJ�+5�̋�Z�{����q?I'mn��f�E0����S����b�����-��l
���2��sR���	]�[��}�������vL���;^b�Xs* S��?m��P�fJ�7�/mL�ӧ�s�%q��yg���`lN�u?�`򭪱?㙨�{�u*2���=]� [f8x�2��s�rk���l9'L���!�p��ՕؚpwL��3�.y���mI�R ����{Ω�v=κx3�/�6h\9� r��3,-�bۗ�\̱��+h��c�p�n�{{w����LB4>�����(������_��Ǩxk�6�">�T	��K����,W4Bb�Z:xx>�'z�\0��]\�������i�Lө��px't@"��s��Fٕc�ӂG�L튍��'�zuvqq`��!s�uJ�X�5��^��UU�La
������"1d@��0a%j�PFDd��MC�W��{������t�9�KPD)Y�A*!�'[��^򊞍p�9��"��ö����V2rZ�]J�7��u"&uO[*�D�����V�Ln��4ٌ<���G/}^����]�kxd��v���P,	L��OWl��Qy��g������[R��ץ𔶅�� ��lG�6�;��v�A~����G1 BSu�=�vN�Z�w��˄���s���'3�M��/h��L���2�e�h��\e��l}�DG:�pIW�=8���W���)�Mg9A)��k9���2���196V=�Ƈ�����
����vVUt��斷^}Q���l=�����)|�
����)�=*g��	Х�뭨](�E��	Q�=t�Q5�ap߾�z�S�z��U�N=2S���q���Ng�GzL!��U[:��7�ն���9à��ҜjtA�N���9��6^S�"Q�!QK�f""�2i�4�w<�O�}E��Ӭ�G��������"��A����㎛�e��+�%��f�����[ ���!�^" �n�L����6�]-\��޳d���ev�9���T��t]���:;��k�:����:%�4�g-C���_q���v�;�ɽ��ۅbH��'��$z�G�}�{��������ɏz�X"u�cs��;$J�wT*�愌i]�����S���+n]��k����he������V�у�"e��ל=3�q���.�va�s�ʐ��SCi��/��ғ�/�{wٷ�.�� {0%cH����g'�>���T����z�f��׍�	bIp�݆�(po�(�*�l2Ea���+��P����u��B��W�6��Bu3��0_���Ҁ������?<�N�t��Y8���dB�����1@0jG&U�KvBA�/��-\	�����ވZavǡ�#ͭ���OIa�e���>!�.�rU���Ϙ�*V"�����L֎�d9�Ģ"/�ܞ��l]U~w*u�a+ʹ��<��f�oT׮����g�֙7쩋�m�ÌM�c�jC]��T���):n��t2�Y�)�W�@�6����\��%��8����R�U�Mpc�R�*U��b��Ʀ����������p��ӎ0�(�e��u��1z�[�����r�y�y�op�KcV��[��G1\����<8[ADZ-��)w)��(-;�q�t�U��+X�P���F�ˆޚ#� ೲ���B�c3�2�я9�h��^f���X����ǎ"�Oqٚ���&��	�N�z��1y�p���N���M���WZi�U���iE�i�\Ad��4\)i#n��{ ��E�q���b�d�e�k=��L�a���,b������Z	�]kI��S��x�Nh�֭�fwP�
�7g����-�}��s<��.\��._�h�8(m2�;�F�4ػپ�����gȧ8���ͺ.���-���#�gmF#Md������3r�H�J�@`�7y�n��{�vE��橛�B�t2,Q�֮���֔ʢُr��;�U���&A����%}y���2�ޙ���n<�lNqH+�-Kr�>�U�Kx��n�j݊�M���h�q�xMc���%�#32�����
FV����ٻ�J둗�3�R3�tyLrw�shge�<��;X9XC��+^�1���"Ș7fg.��d[U��J�u�ܺ�$4���&fn�nl=SK�_]Y���ݝ ܃wě���#��:�����9���a^�l�9�����Is�"F�ݵ��D��/�P�d�3T�Ĩc�)m�Hyyw�C*J|m�nc�s�g%^���s��Rn�(N�یER��f��'0k�&�Ǵ2�}��U���z�`�����R���C.�n�ڈ���s+ُzy�U�ST7��eH.�r�L�^],'u�I�d�zU�8�7��6�y�Vf�nE|p7���5�
�4���IN��ΰ�A�G3wv�5.��=9�u�w3c���:��ڽ����6ٙL� ��cU����ư4-j�� �|�����Av�u+ߋ�N��L�ҽ���B$�z���37Oq�H ��Wz�s����wr�=Tv�:�Q�Q�ξN�_\y)Ы�F`"d�GQ)}����.�A����%�z��c9xc��/t��eօ;C�M�����,��ad��z�jT��3�rD1�eV������t�Ofk�U�J�Yj�|5�6�}{�GSx�S5;_�M�u�r��T5��g�	�Us�k���DL�e̜e�XF��b�ĴM���RN�uv����]n�Ic5p7���7�+�i�N���{�7N�0������[�D����/՝[$2�@N�-Sa����hN8+�1S�;�]���'�jE�(�`���Rr��N}�~4�����WO�T���S&����Fn�l��ܑ��`�q���>�6Bahs6���U���-Yv����Afc菾�1�����*s�ڬ��+����4�K���cboS��h(�EbBg,ُE�kl�'��e}��en:k[��Ƴ�z"#�������`�������b���vJ�o3N+ȁ���f�K����UR{��b�8w<w.�����D�|�yzS�٢�A�GO 7w��ؙB�.ÒR�2�M�<�t���ټ�9�1u�荊K�ɌB����lsV�Ck���S���uҫ��l�� u���"��k�\��Er�;�p(z����(,� g�߿9�0�ww����,�t�"����'I�զ� �UC�?�r7,d
K��v"'3��y]��28��J�����w,8�:踑�[���Ф=����<}������ �'����v7��'�D�=��<�k:�l��� ��&�j���u��'�����Q�΄nE�W�ﾪ�7B��[(��L�=ǀ&J1�O鿠��W��}/�aV�vR���I�]Y���|2y�f���P��-��_+OP���+�K�'��V��3���ӵ6�J��KŘ�Ğ}qt\�|J5)����;A���v��^��R%�_D}�������u�1�Q`2Z�V�50ȩզ�p�d��{��c��f�.)�R�#���'B�Ʈ �%��9�}��+��ӓ3���:Z��٭�z/��8HC�JFJ�h`�L��b�]��������MC�*�s�Z��,ɵx���=2?<*G��`3�8���9Ń���wt�|�
RԡI)
���YҁTա#)@�FF �� �0���() @HV��P�J�"���
�<�d���m���{Z���w�6o�P�jq�P��Rh���z�K�v�,�Z"��܏4����[��S�e���kd��t�,��4��a�S5q�<���G6��X�xN��6N�>]�ܷ�v?8,u}�g�>��ze]Ӈ=׮M��;./�Q��S;�}����vc�����><��끹��S��d�N�t��*TP�Q|
_��}�z�|>���#�<������y=��r�0�4��Zva`�ěc���#�r<�J}�Ifr�ғ1�����l�l�Y���Q�w�0ǚ�\	]6ՠ�BFe�	�hn*sfa8��ʓ̹�ks
�T�!\�՜[���T��B�t����b\�W��jnt�K��c
}kF_�]�N�nw,eip2�0�Zw��b�#�>��R�J�v���ﾻ9i+k�R�֥�f�Q��"#������[���ɓ���0���6�D�w%���q-���ʄ������6�1��*si� ���\>��Ȁ�@z��5='lӡ9��7��FD.V���Ѣh�a`a��vK/7j�Ө�@�@:w9z�^*�td̻���,t��/�����kӿ��1e��t��;�՗���T�.�2VY��ý��/T��t�O�˃*Ύ��j:c� Y%Ļ�LHh/G��f+�n�.Ӄ��z��[�s��-��lv�au�bâ�Oz\�9�/�X8��ѯ�+��F���f�]V
�s������"f_�=+���>������گ �'�׹���Pp������C��6Y� �U{�W^;���{vhc���>�Y���y��Tj7Q螡�	��������𤨃�
�A)V��w.��΅B��Գ�3W��e(-���EG�_�,��I�X���x��m�, $���C.�[B�����(N����g^9w�5¹_K�φ����W�~���|N�(Wa����䎮�+�O/q�+Z�%��	"�q	b��.J���nFjW.��x����9�r�]�|fF4ʬ�����׷t����Y;#4.;��ce��=�|�FwX�U�0��r��^	��:r�R�M�|�	�pT;ܖ�x�)���DG�:ԙ�^��DI�~s����la�{�c:.'�a�|j"�s��9��J��=�sX_=��<���jŮ�`���&��{��G�O�3:\�� �2�pNz2�xؽ�%�q�:{�#�}��,�:���(>|�@#{�kZ����}\;��ZVB99-ǲ�juDU�z�X.q�V�OYy;znjz��a;�D�`'���%���6d��G��|<=�G��և�a����j>�Vkǐ�j��n��u������[�O,Y�����&x�wn�9n���"���E��G��G��N�E��}�zq�4��YJ�h1��az���]U��,�;v�8��wy��<d6��VK�������G�G�[t|�k��޾~��9ݝ�M�(�MFA�DHE�P.�ӢkWZ}��q�{�����b�F��ȓC�t|iv�y�H�֧%ٱ�VM��L-�Fb鯲��o������VɘMjge�d>�ʋzH7ۏ���P�`xU��,WYDʯS�8��D�:�F���Z�ҥ� D�DxP��P�t�WU�5�T���Ʃ�2��皬��ݕ���i^�Gb5%f!��rK'y��Y�6s�j}kS�Қ�}�߾�s>�V�]��;#�� g3�P�u
�O5���/�����p�5jX�דg�Q;�N���a��w�	���{�%����C1��U����N�"T�"�=�`�%p9�F�xWuk��h7h�vt(a��+a�H&��:=5�dD����Z��z[Z�+5k�f�K�,��L�Rˇۋ�n5�y�*�0���g��L��3 �w��C舌>�.0:���`U.�����[�V�m��9oNI4��-ٙ���{s��2u�mD��%+�f�yx�W�[*�*BJ��ZU�������ɗ�N���yY���4:���]�۬����uΈ`+�XfE:��ck�:*�����Iz`l`ѳU�7�������'3�RzZfwf����Ot�-2b;6���'Լ�v�����|^UN�n]��ƛ��sX���D�H�	���,ú�7:vD�y���D}v�VXj�A�<%ne�
{���;�Ĝ`�<��E;-�<cw�����g�离�d<8������C`[T�l�U�}��舝~������T{۫o�|�S�@�W�i�=�<
뺥ߌ>�e�V��e����tz������.r[�[}�LW�}��><}�dtJ��ǂ�$�'�ѽ�tێ�;1+�(�$[dݏ�FXH�ѡ�Y�(mUs;���ͼ��/CUҍn����WX`$w��3�T�,�� ֯f�c�Y���MTj=3;�4:�ZgY�6��N��-5W�K'%]o)������	�����זϬ��^#j[���"ǻRy��BÓY�}���UH�B�`VE���#Kb�Q-(�m����PB���X(�#b1%J",����xр%}�JOB��&_d�U�X����]3�EN�W׸i�Q�º�s���]Y�����A)���ځ���kE`+m���Iμ�|G���#V�#I\��A�yQ�ؓo*�X���U_4��ʚi��n�~_�3�ݷ��6��q�Jn�A�E������ڍ)���Z��[.f���=-���MSLΫ="����	�5/A���^{�2;L�;��ȧ�f���;��ƅ��Ɏ����~�����*^t�ؙ�{:��LwS�E�
C���h7�(m�f���+Y+x��:���ʩj�ӝ�\N[��J�����t�|b���9��Ǽ �����e��A��t�3�Ѕ���u3i�0g~�y�����ޓ�g̫<9�G#� 5ڢ���(T믰�VVu��県(g�M�=���S�M�l�8��l�WJҞ��u�7LR�7���L�i��g����?���x{��o�p6!�� 儔e@(�`\�����j���Ǚ�xK�[���	.ι�)r�Zh�#�	h#\�5��:��SM�ћU��f s�%���z(d�Zzq�}5�r�n��M�,�X��S6�T��{"�1{L�������S��]r'�WL��r#���U�G��]8��L�T��k��=_U|_�.t��0;��<���f��qBG����1l*rԣѣ�sջ��/�Y#xÿO���S���J�Q�k��,/3�Dn�v�`��8��^Gc�d\�J��QR�L;Q�V
h�WR�3���'Vz2�FC�R�����t�,��.�,��T�����5u��"љ�{�^25�{�l$�"z �U{����e��a�%Lܩ��vV*l:-
�7��\4S�ј���C9:3o���ַt���^��i#���@��:TDEO�)��+�r����6�������EYuZٓa�+�9�4gB�7��+��>��D���[����)9��0�iɌY�h7�a���k��9X�Iܦ.
tl_D��b]S���Xy��ln�IuWVc�P+Z�8f���� �U�HޛS.d���N����Sn����R�^I�q3]G�e�Y|8¬%�]*���n�P�ȆJ�c���1�w��r5����2]��Κn8i�ڪ��ܚ�O�8�?O��cX��|N���jvѳ��<*h[�ܶ@��I��
���Y���';E	Ak}qHq���E�,n�-x��빹���#E��1��'H��VY
��r�VTZ�l�\�K�W�f�v289��R�ƎzL�}����;����ïh���?���,xX�uՈM�>��\5Ő�!1-N�5;3)�c���ȇr�`OT�^���4ŝ�p��/�.\XR}<\�Jsg��۲c���#@���w8��2��;����T��~�!N��v(X:_N��%B�x
D���_W�|�s�GC��������\��BX�w�C�쵗�mH8��+���y�xԍ�%��>�{�U\;(�N� ���G˅	��.��H@q���*�7CU^\��S����Q��v���j�]@@|,����t`��`vIg����ۙ2�6:ú�
�%y�
�]���z��,��[JZ�1�(~�S����Y�����@���#iD�}f���*��mA7i�*Qӕ��s*��}���s[�P����:u�΍&�ȳ-<᝷!%��ʱ��G��Q
��B��!,*�əWK���
 `��@��hT4��1�>4��n��s�Tw��ލ��-)ē�X��K�iɆw���N���!�m��z���:^�H����%j�A/;�;O^���C�ek��CL�О's>^n�{�v:�obW�
��M��i�eJ�~���5A]Q�aZ0q��,��w��0��c5̝*��C�8OqIJ�	@}�Я�*ђ�|�jt}b�*�M��):��5��@��;)JtD2�p��o�Ӊm����oh���T����������'%6�vTܷ�$ڿ��Uw��_��H��GSg�)<�]?��#�W���So���gsV����VfwWT�%vv(���M�k�@�jA����=o�&�+ML˫���E��`GmI�bHR������X�ʘ��&�t܏��N'e+O@�\4��E�Xn���!�&�g�\�70�RპN�n�G^܍qܙw�*	d��3�K|��#���S��;�{5ͳb�oeٱ�z֛�-SV*w	C���N��;��&z����v/������,���/a�t��qa�Y�o[wrEQ[�5�n��oH��ٌ�����ov�h�!��S1D�Zٵ)�XV�o>���-`R�l�ޅ�p�t��]��&��ZA�����[��K�ma�����6�V���@K����bt��B�=�����)��˲��e[�@Xǒ�O/����շ�6}��&�=1�e'd����3�qxV^������݊glKm�$:�K7��mmv`W��tH�4#��\vn��RJ�$��Rж���6�����}vԲ�����xe
ΰBW�ʖV�����Kr���=�;V�N�F���)@��Td��T������+�sb�/�V@ѝ��ۑ�Z��&P8�%o��|��l�\�%ڋ�#4E���'�F�(�X���RӎƼY.�G34tA�Q��wDk_I.��ʈ.���%)پ;v��"�������QE��v�ߊ�֓�/x�N��,-us�[�L�P�3D��oq��	p�����}Ml��G|+�:,��)�3\n��s*Nu��Ѷ'��\�r�C���5�ٺ(Ǝ����Gr�vU��O:���u�#R�����}&ԙX�|�#
SR�s������=9}[��[�鳅1�9�l����:�	Ra� n��k&]�ѕ�
�5r��Kt�/�]f-q��e����M]J�Y/f���vſR����}'_�nJ����0T����ykK�'Y�G�ܳ6��.��vPjX����A��_��}�ȬF�����=���a�V��`��UuR�������p��v�	�"7uat�>���џ�>�w���;��P��x�!�����R>����p۴���ԙ����N�?����]K3�8���FX���R���#d�k�0z�F�F�کA����d'wB"!���{�µ�V�Ǭ��E�w�{���HM�W���ݮ�K�M'\q][����������}7�e�n���m��`�Y4rv(PD�Uö}�����~o���.$�2��¢�2�+E��jZň� �����j��ȱFY����k��l�X�m1dɖ�$T[J�FH�̥b:�ӖB����;��9�y߆Y�&&]��]l�ebɭ�Ѣ�K����}]݂퀙�F ����xU��;"x�N]d��Z�_"c�Hvѭ��n�rh�N����g�*��|dJ3Ȃ�)����/{vm��T�����űn����zv�""����{�.���Z��]�s,`Ψ�Y]�����k�3Od��L�z�Ͼ�.�
�糽�=���p��AP��y}�t�ӓ�=���[Q�Iܖv��X��8�v炚@!Q�h�5���PO��rz� �J}3�sɞ�ݐ�M���Ʃ��Q���As֏O�]x>�ӑ(c���2g	9(���ܫ��c3[bx�Ex�;
�P� ���Ҙ*��s�b>�#�����ۦ=�e$���y<�5�����Z����Y
'4$v�@{X�ҼxtN�c0�-�����#}?{YiO�3:K��ѩu�P8�w2Q/��IvC%[�?y�~��qVIPEQ`_�eP�
�G����{w���M�髝��6��ʌ��r�ꐤ���ŧ�v�p$��
cs�M�����;H�B��EO1�69�=.,����������S#�X��/菴�4�'8+�5"�R��zM���|�����K�H��J��������"zE�vY:��=�tW���y�ll�x��ç��Ml���6H#G�0yz��oK�-���;�kfS������o(u��S34�D㏢ً~,�S7�J�R����4��m��Q��1�ٚS��e5�Č�u���ӹ�JMh��*y\=�~��Yz�Gu�{�~�@��-����=�t�;�zP*�����OI) ��|�a=9BK���S�в�9+����y�u�j���El>t�y��ʚ��op%&S���z�]�/�ٳnkSJ�yu	��>���z�3���8�t������*M�T��Tb
sW�l���ke���7��m_Z�V��l���])pgF륷	/�N;���NK���@��G���F[v���ȫ뙁�0��C+'q�,�w���.��z��{���,kP��!�/>����cEn�q?�ܲ��ds����7���7$�6��r�����@���c.�MVVZ�t�=�s=~&B����_G�!�6��e_���&��#��|K�vQѡ_'x��Z�]9	(�Jd:�z\�]b�uڤ�8e�s���h���< �W�D}�E��Sh�`�&����v&�Ye�b�aN���rm�芜�[J�C���]	fL6Q�! ޝ��p��DB�5��k�j�<R>=������P���d�:E��I�t��	����{�F�Hx��UW5�m�}9�R>���m/	��]�_���bq���[���ӝ�O�^[Y_���>���(wN��\����K�N���y������A��!EE�V1��[eS�y��n~�n���[�����kM���z�`��(�+8�))�Z�a+���7��=9m��;r��}F	��h��a�9v��4dݼ��$-d�zhlm����zn�g<�]1��3��j�Wk���ɮG��sDk���]}3l��1خ�%�����#<���R���:*M��G��B���tC�z���{�@�pZ�[Uj����<���@n�m:|.��7Q	��j=��*VJ+Fp
��i�mB�b^��B����������Ht�gtm"�2�}�6U�o$Q�M�(��]H�"��]��l�Fq2�V⭜��-����oq����t&x}�Tq�k[����H^4�K����yY��ۃ�R�}�s�x{�z���Z�g��᫞�b�L��i�h`�xo�q�MA�����/ �.SE���*��̫�a�7.��DE\:E�]���̨�:��]Ȏ��*]�3*
��7��ӄ�k��7f�$�A�e/�#�9[����z�[1W=�w����|֓�6��ܛA
t1���+���εp���qm;���.>�B�g*;�S{(p�.}�R��i��;�K�z���C������|��q�f���즪��bW]7�|�'0���v�+�0A�����w�ed��T�S7�*���ɘ�N�l)H��v�ʋT��(xyN'	p��}3I�I�^�g#�;���׻R�:j��&h���nN�8Y8���M-iq�'��{������o�e�Ӷ�8��W��>1�Vz�m�>��دdX��9�ċ�P� �$hlL���O:���V˨��h���JFtڰ�ns/�+��q��	�fa��2��g��M�'ǥ1�
6���/��qT�=P1@tfg���҄�vx����Q�\G�	�^�˭�h�zg�PtZ��&iH��r��(v�����q�	�!�#���:�UMKE;�:���c%S'�+~��g��|}�_����u��+��Mk%�n[�!F1�,`���#&-"8[@EX�A�EZĂ��(�D�qF�c$L2�"d�T%ˑ���)V1Ffi1�y����m�N��G7�/�A�*�1�Z7v]�W�!�Q�R�t]���q	�>a+/�7�)��O�ͻS��c�Zb��$i����g��'z#Q�HF���DP���0_��ϯ6�����n�йy��U�ˏ;�}�ѵ�q���S<��d��V��3���m�c�S���X륈�u֗&%�\>�P:���S��&�oQ�r���3�P�֟Q�=3�hN�>��}����s��,ҫg$�=b�I�5b�Rt<�8*z�27�X�ö������[���x��>��#/��C,�Zc�� ���N���u*m���d6jp�V��T7 X�ё��7A G�G�N{�s�w��ToT�j:��B���wY<��̎ᓖ�Z4�|
����B$�&�F�D�f���\�����__���՛�p��0f��}�,��6Vhk�M0�	��
����+-!v1��I��G�"�V��IȁbJ0
@�D 2[aTI�./��)�H�#TA�ϯzg��|Vd9�KGA�\�7����k����m���ׂD���5�gu���2�j=�����!N�]C�{���0M��+OChF+�/��)������)�e%�� �[d�AaVt��7�:�э��mvl����p�}�l��w�� 3���Cw�E��-��$����x���C�6xr�hMl��xɞfwC����1߈5}>�����T�<�;�m�;����U�֩��;���.��t�a$F'��.��|�d�ٱ�o?��=�>�Ԧ=�����΃x���qq�ܫCUܥ�:��XY�+1ҵ;w��_��|��`���8^��'Z�荚��4{NTy��8ܬ�g{����n鼞��y
�8zp�|5E�{u	i����� F*��z�j��(is1�v�����Z|�ʧ\ӕ�M���X�d��G� ��u ���{����|�1r�H.�xk��KQ��O`�3.�z�u����I
Wu�狨�4n�����=¸����3wjܩO��2}C��î����
�P�xy��&�F�'���ȏ�"��*��ݞ��Wj��6qQF� ��,
��u@Z�%I��M��=t�u�Q��9;<i5zW2��fSR�h  �(n*/˖�}e�'\)S�uКe��n�r��,���l
fd�{�uM�(M�=l(��j��R�l��1�L���g*1���D>9<X$>ν�SV����όF�[�-_����ݔ���JD��n]L�㠀�eь/���h� �aC~�����C7�/�P��°X\Tɕ�/��m]8FV({�`H�%mWpw{A����t��6�넛�V��  �vh�0��M���Q;�X�ΫCPZ5q2�Y��]V�}qtު��r�y�[&�2�`��b�������5��~��l��"��r@L�"��H���T
�0
0�.��	�������:�+���KL7]�m*o�kJ�GN�ڵ��4��љ�0��={�\�^T�œ�u�ϠLT��Wv�]d�N�\�.�ő�
���<D��/EI<sQ�!����C����AS8Srg�m�ջ����\����W��D���vM��H�^H���u+�w�;�"����@9���Mb�4���-Y���J˙�ﾣ�Ǟ����\G��1A|=���~��l	�G���Gʅ4�"7t�{Ig;�p94�Z��ZZΨ�:L�J��|N$`t^bKh�������;��G�FՕ�}���y��9�u�UP2ul���f��U���9�fxE�A���U���+'OJΒm�p3��m��ä�0�f8����\M�a)T�s4rz(
��j�3{qQ�[���J��4��>��)��ľ8Y��:Wa
8�{���t�oY�(�]�(^H�L^įJ����>�y�wBz���<��y</��r�5��k.���竫hVY����U�R��|�{��4��֊�n��jͺ��53��`�}���{G(��O[Q��3k,�ެB��d�iQ���S��l�}�|wY�g�As}���0x�R�*�[h����W�e7�D�{Y3�r�.l�b�P�`�)MՐdl������Lv�jje�F*�4�G�Yh��݃ڡ�߸���02��y[C=e˽������q�D�$9Th�nl�X������˂&��g���a�C�*����$�f��֒P��u֘h�u��Wy��`Z��ʁn�I��{k��^8.�7�nT壕�]w{`:_p����>��"@P��R��
�H��+i5�E�D�u���)�E�#%T�̢��H,5l���Q��\#��R�����\/-r��)~�M�Z+�X��-9���ݼ�ְΤ3��Ŗ.�����Uc{�^{Y�8�Q�L0)�
��ӭy<i�i=���J���(|p���� �.�)�O�Zx]]�od
�k��J���V���?a�W�11��O����{�+j�ܾ����hXTT)���B���3iA.�r�V������Į�3�Jn���:���6H�$8u훂+}w}.w`n�s5K˰��g8�BM�;rcE��&i�ҝ�1�d��@v�G7�7Cn�����`u,���A��Y5��X��[��|'q3��8��,�O�K�Si���4e��,Ys�(�9	���,!}1��藲U�ܭK��0�Jw
�6�wP�O*�۝3�y���QMyr�&�
���	���<��xp;��wbkGF������*�-�G�B�0&H�kq"]5��\�1Y�d�]ui#ep8��5ن�����w�j>�*�=z�t���x�-L�:)A$���}oj�I�au�j�U.�Tb�5P8����
���G��#��%]V�:&Z���ѽwW�����0�x"��k��8;h^^��ᣁ� Vs_ *��-|�4�F �W>��
ŝ�~I6!u�'��i�a��u�H"�����"V�o:�ގ>���w+~�B�V [ �j�A�)�-:�9Ԧ��ݗZ�����Ho9@�V��c
=[�ʆ�ۛYV��Q�=��<�P�"�w�Q���c�dW��a�L-�/�W�>�et1c��PPZ�_gǷ���셭V�����A��v�V�l�ܒ�n�F��76*��k����Q��l�)�]C��t��; �H�zuw�ͅ��B�E�0�;�z�V�i�n����J��y�E��G��o�z7ז�r����N��z�-����4v��ަ襺��ҷp���N,[zc��trGQq!��er/7�V;��VPGnjg�S�I����R=�BW2  a�{�����_����}#����qJv>�����;z2P�����vbC4��ّ��t�s�h�g[�p����.��e5#�X�4�y�"0(��g��W���W���O�v�'�,̍!u&� Ƣ�r����3�9�i����<��<�����U�s��P�0�17
9^w�C���xy@�Bz�D]��֟nν�����uV�ǀ ~�g��������z�bg������ Y�7��hE���۫.xy�Ξ�r� ���t��6]�k����G�s'�>�tZf/6��n�*�;Ev)tB��Ź�5`�z�2c���g�<lpt�ރQk;3mR`��T�e�:�No-UA�l�9�.vWH%�%�i�"�,T�Hꃍds(0R �3-�ز ��&[ ���%�YFT�]j��[f��EfWٗv/Dk}6hkH{�yN�;h�)�����䵛͡�)+ُA�δν{n�G�*�+eol��0��K�W���^�W��Jtz�I�_��OxҙA�:u�QW*퍕�P�t;;�*uR�׫���1�2V��Y)��t�\��Cl�ᅯ�'R�9�t�ڎ"OF���3������ƎI���Bko<��0_]_?.��ڑ���i	�M�/"a@�ضS��P�i��X�	���<��Z��9'8�䉔'Ww�L��ܠ�p�w7��N�m���ZT�C]u�ġ��C�Nu��Գ�a�Fe��b���}�gGS�����᜛LIS�\Y��$���fo��X��^5"&O#��]o-H���/{uSn4��������s�����k�ċ�ę����}�'�CEӓ�4z��-��v���N���uUP]���t�C��A�F�/[[�|9j����o����B|$�0� "�RH�3r��Fğ�ղfs��JYJ�Ŝ [&�yu�b���(VR�/a��K2���76SW=w���]l��r��l�o[�c�"ΐ��!��G>�O�r���2�Ւ�3@��WQ���9�xD�9�og=q/'p��90�����v�q#h�Ⲩ-�C�g� �x�r^;8�����XY�[��C�or�煠�T���M�1o�023]�t-�R��a�t �v\چ��������}�\�='���i���k�$��p�1
RÇi�s��%���\3Zۨ*�!�bb"�Aw(�t���ճ{�*��#�^菩�P�A=HW�<=�0#Sw�ye>�Z��5�F]�f��b�ŧ�Z�G�.�y���+�1%�2�>%�uf7��ޫ��{Jv2w8��-i��Za��]��S�S�֒p�<}#a&:��#�l9�J�ؕXgQ���%��������*��+�=�\�/^\�u��r���)���Y��_7w���d� *��R,�@b��HhЇ��(r����k^���n�R�3d�	w�d�5c��U�َ]tVNh�*V���_Cmi���d�n!3pڵyW�4@ӡ�:�;�x�ԺD뻀"Z�=&BLS0� ��ޭ��<�Tq�Nr�Xyw�(���u�Oy9P���H�Fi3����wX�	XF7�y���	۔f��:_�Ɣ���F�iʢצ���V��Q�P�2��{ێ*�i�ΓNm�7/�'��\������@v�M�^s��)�Z�+_	i+���+.�|1��MN?A�^����N�������n󐳭�R��;mnc+���Ȫ�9��NЙ{e���:2�їX�7KG���}v��n��a�'�(nuBcH�a���YR�3�[;�ܫy��ݱ���p�5��B��Z�T��S/�N��(�q>�V��x�<�e��d^S��yVkPR0Nbv��Ys�B2ƹ!��$���ZW}����l&�4P��X�̋�Mv�5��^�xiH A��d�^DC�:Q�ٚwb:biZ�Q|�&9wg=�OEu=���ݖHQU�)�t��1[z�}V���:���gz�73"�Vܒ6���f�wv%f��s���d�2�S�68�\�Ǭ�XM�,¦h�{���C��x��4c���5�x݌�uW+9e�&Pzn����G�����OT�"Ұ� Ӽ��YBV�r,T}3�r+mU��I_E��:���e�M��/�P�����(=Y�xg6�s����p�^$a(B�̰Ie�/����.V��̽U�K���>��j�h�
{�͹F:�)�6AD�ͣ!�!�T:�zY`쬱��Wr^|X��()�K��	�4�� u
6L�yu9��wh��#8��r�S�j�[j�c�q4��V7"AޣQ�tkc�X�z��&���nڥЌww��u�r�E�3�����W.��e��
`w	�D4��2��@��u�y���"���MyP4���IY+**���� ��� I�0�OT�T��H�M��y�F��1:�Օ�jDf�i�X��=�U��Ko���˶{��ܧQ>Pn" B��p�.�)1�%n��K>���L�OS.*�//�ܜ�ߊYw.�gr��5uE��eʤv�kˬ�욵'�\�g1��y2Y"2��p����w��r@�uO�b�lZdU���4�kX��l������	E�|�"l+�MwB�{MX����1�k��N���>3j;���U]E��̷���$�"��ҿ@���G�����+�5CqZ��;:��t�-y�,�1���g�a��w�y�Ꮐ�Ş�,�� Ȝ0g	���t�D�F��:���}�Bi���^���aй<7%�S���d�N̠�L�>�����s��{��5�߬�~<���o�Q�a�"Ϩ�ML�W��E�x{��c9�h�"�ZxR����9.__BN�C����a_3;L��+�?X�J!�(�,Ll P�"0�*���$��I"�E&5@q����:~�X.һ֮�ƍ7��Fr��N���Վ�gb�&�1����!�to[�0�we^��s����u�r�� ���|����+u�<�-Vv�=:��!|5�E����{.m_�j���M�+=���3���``�k}��Ρ�7yS��lʌc5��e9&eT��&Zd8��Z�7nb5�^%�Ǻscq�5N[��,hzY+d�6{͎�<��gC�uVH��х0�m�Z�}�kKu�D�K��[
%s��E�0`�e�Tڿ_��I������@j��|2⋝ah�JiX���X�L�Ry*���~�� w�ۙ�t^Fs��d�� �|K��L��sz���l��;�����Zp�	�i�1w�{+�	��i��'�'�:�tV뮒�?FZܫ}oLM�7��mY3�z)D��8��{�W4�5��5̵<^�\d��R�Q��c�w;��M�&��Ǵ���pR��8Ny̛j� !x�D���R��#
}�(���J�Ĺ�M-��������͝����];r���n�>DWc'Y�Ƙ�t��]�K��]�6)�l����g׏ɉ	FγW4]F�4�%�)a�ȍP��^7�T�<�׬�7s]N�uq,eN'�}�D}��r�A��8\��DDt.��U73j� GP�eHon�Q�Kq_O-9���6��Y����E̫;R8���s����2'��N�`x^�Yn��2����^��	��!�;\h��e��0��|��|��Q��;���]�%�`Lk6e�� 9��9N����fq��f�����|�x0�a�v5�S�`s73�)���z��3f���syE�}�Gޘ����_��{ެ����wc�
��d�2�t�� %|���g��n�ƌOT)}M�m�|+����1vј��ȍ�����vF�Ej�[�{�/�M�\�c�	�u5��rv�C��71���N�+���i�M��zPO9�+?$%b�2b#�ĔRm����`LYE�6;�V�c�lE���on��Qڐ%%�����K�Q������{Cϥk|{v⏟B�.���v��z�f�m�uT�\�V���J`^*s�z�B��;��8��}�w��|�r1�KQ� ��v� / ��u87,n�@�-���:���5���+�W��-��~�:R.�l�̖��'w$��H����pki����)Y���h`p�?�;�n��l�6��O�F-9.N_8�6j�H����Қ�HL��3��^�"�R�.���Y��xbz9���^�6rԃ���x�.ny����=��]J�~C��f��a)wz�]�Zw�z8��p�9�C��S����ĉL��N�f�8O�--�J���F��|��=����I:}���B.�9�D�f��j#SZ�s�`��h�6��X z��]��r�i(��UZ�_���`l���d"2� !�ď I>I=�X�M���t+�3�;%��]�|v�X����?@�f�SW�}dی.���M7̜��U�W<ٸ����w�7�85���^��ņ+ �wx�p�L�zd�k>�����=��"o�w�4;�콤)w]���.���zaP��~>��##� ���j4��(��L��-�y4�F�	�ா������}�֣�٩��Z��B��{�.�V���~ѷ�j̞6W�.ƅ��l�x`�,�=�;cﾈ�D��!06�C~�Osy�S6\^5Ma�M��9|v�%ꔍKw����_Z�,��%�/&���6���zK��1t�KK�Pf�m�=��ƥ�)t\�L�Aub�]˴�{NC���Ǹ���WN􈈋��!�t���b�fnw��n_c��({7�&�r�њ{����Ŗ�&�����ؕv��BP�͗Yhs��L7��I?�	$�Ą��Ia �$��H	$�R@ I'�a �$��	$�� $��� $���@�O�BB�HHH��X@ I'@ I'�I?�I���@�O�$�� $���I:H	$���
�2�ɭ���b�����y�>������>��A��ƌǾ���T�B���x�ծ��g\C��,�
(S���o�}eA���gN�]���.$o�oXօ=�r�Y��78{��U��<q���`�kky�V��#�    h ��24Ʉd b0 � D�T��� 2     �� �U=& 0   &�0���J�M0      ��ADd�    %hHe124dFFQ������M��tNV��*�5>aڢ�5P�w��A@Q��������/ 2�#K"(����P�B�To��ފ�%�S�tQ�v���O�A�k�a�~Ka悠W���C��_��8|_:=ֲ��O�צ5��G/JkE7�b��K���u1�ZK����]Շ����MѭM�	���7B�$�^ �U��r')eV��D؇h��-^`pPoMDu2�%���z˘��Y��@ۼ�$:��Mj�q� ��n�ja���IF�c*�ww�b$�J��ݭ��)��˩�n�f̙q[cr����۩�ű^�OEx���\!U45h�w���ׇ`m�c"{]��d�Zl����
��e+WƲ�f�h��\���ƅn����h��Tr�b�������j����<K�.�*&d�0`M7��d�VQ�H���k�\���t�,ԪNX��wHnH�1F]=��Ik�Vˠؒ��~�템�Ն�=$�gC��X�uh-��Jǔ@�F�D�F+-��Mܫ%]��mM@���G5j�n�+PF�b�ދ�~|��ooL�Mݸk)��/q�e�a�	n�J8��b �r5l�����z�����jbl�i���RL7)��\��Q RXͶ1��Jm	%���v�Z�>�E�3#��8�r�	*4�Զ��/�d;Z�[�/t�y���A�5[�=c�����*�W{�S�x�h�9�qa഻z����}�u��d{(��@��&�_I�5UW3��$<�T�PH[���@P�Q��ȁ��z�/qSYuQ��m��m(�J6ҍ��m�iF�Q��m�m(�J6ҍ��m�iF�Q��m�m(�J6ҍ��m��iF�Q��m�mF�J6ҍ��m��iF�_��J7�_6ڝ��UfGʡ�5�|�70�D��1t�fsu����\�'k[l��e�e�쵸�#����y]��C�cΛ�!T�D�56�|ޕ����+���{K�����]�ʁ��_Y�yWu*%��D]�{m���"3b�TΛ[��'R�\
0;��^��@��������q9�e���Ke��e�6���a�/;�E��d�V{�[2�bG7+)�t-��b�ˑ��gz��.Hl�@oiN::K�Ɩn���"��9g����c��A9���z%-�f��B5;Z������0���8����f���AnUm��o3(��[qa�n��&-=/��7��-��U��(V�ie��̍\��CH�fE����di}o sYLP���QL����u�=A���:�_V��L�g7%X ����(-��&'��9y\Wm6kރ6�;܋)gE3��(���wCî�@�̩p��
ˑ�Z �����$�0��/���I^\��_7l6ژ2hȆ���B��(qU�d�g3Q=�����Q����#WQ�\I��2_7:J�r�	p:ݖ�2�`���jq�3a�`��d�}���6 y Ȇ&����0arq�ӓ+A��;���EA�`��g����%�-��٘7����!L��63��h(�CT����<5��}˝�6TQHF@�F�@lRP�A��5>K��I6���IF�Ŷ�(s���Ve�)��ܷUl�|�a�;/UJ�����	�d�$�WER9Ah����\Y�� D��{w1ۍ���3D����M'9[U�T�nz�9��K&�˰AeϏx�j����,(�B|�ܒo��[����(L@� xI�1�RF��z^\aj�*���ψYOПxx�����M�w3F�&:3G�]JkK�� b�Ǧb�ee+����+���2������{k�<~�󲨀�<.��_�]Aӝ�I�XDߕ�U3x�,J��P�+���NV{����sw��M��_���w��[3�� �=.�����&��ll�r��ۼYX���-�>:�@�?��TKp�h@���T���r2f�dS��ն�hY�X���}
�w4	�����������C=[I,�z��n���vw%.`W���u�P`��?��{���$�� Ow��
*���;�e;���z���}�����}'7?{�6W_]��O{�j��_ٓ| 	M�~�(B*x{Ǟm�����Ϣ��P "�x3q(�Kh���fYP�m�|u�a�L����."�
�p�i��X��ƚFٙ)7�"s��9��`i��w��Ղ�%���f٩*�؍ad[�:��X��-r���Z"]�ҎƟ��P�����̻���˼��Zm���JGmS� Τ�@M�f�{K/��u��y��k���3���0���-=E��/��B���������or}o9>���f* @� �4�}:����#c)�� �H(P! T���*��@ �Wv"+®��q؈�7�vv��7:�r#�,M�W�"��"l�]R�%�v�V ��:��M %"-�Z �
�F(��E7ҫx
���	X�� l�&�B�p��@A@�T1� �*:DM�������R"Z��@� ��@��\4��3]�Ko�k�w��ƛf
$�%b����MkE /�B@
�)4� J�@��@�q���(�\�3eT�@�C�w�gD	���⚙uZD� QQ��vװ��έw�����,x�Ьf"Q p֫���L��#�L�TĶ���wD1B�Z��R��/��z]�<���7�.5���'Y� �N�
�붋T�E��*��a��R#�U��UvCɫ��*��Y��M�V����5Q�ZV��*Qp�=�� �:�s�炮z��� �h�4KG����xRZ&��X�o4X�W8����+Zf�mF�WE�G�� uҧR�U�y8��Ru�p@܊ש�-=��CQ=t��&��B�@p��E��w4���דe��V%�#Fڊ�~��iJ2��z���~XcUƺ�C�h
TO5q��[Tc��B -*n�M8���ֺқ�GhBڭ�!�K�cޜnިw���$����2�֭+\�i^�x�Ct V6׍���'.(d���ZH���T{���ӏ&��B��Ŀ"щ\����e�D˖d1��4�7��o�X.y�Y�\�@	H�N �>��=@�����!�r���@U�F�\E�V��rQ4�y��8�@�
��v���b�y����|��C��#��bG�ư0��[X�{�uל����"
h<ߖLj�@Ƶ��u 
W��hi3��y6�kR�4ׯ��i6���5�2J<jIE�p��k�oMD�V�p	<v���C�%{���#�������qd)+�
*ضV6���)%T����%�Zy����j����t�"� �F"A3������B��Yp��gn�IFے6ڊ���]ќ:)Kw:�T�w:��ҕ��j3pĺk�b��s�U�+�ut#U��N�F��`�ق��ֳ�K�H{b{�!�����"
"�z (G!�:�D�16�­�� @=����1�V�q���[U�݊���cU;:U�mZ�IZj��Р�O\hP�����m�]�TW�B��@%	$A(G��膭�S�����u�q���h�Q�7�3��(�J��ZL�U��U���ܺ6���iW�m��T�h� �s���S��F5���M���5��Zq@��((�
�|8Td�6�`uP@#� q�IL�X��pi}o���V��o�!�8w&%i1�@�mM�J����<ܢ�[MO����i���khZV���Q�Y׀�[tF��.?�j�v��=�6c1��8�P���Յ�)�;�3r��xxg�֞�����8y	�B}a�}�	W�E�G��㕏����yr���j����_0 졆|��9�xϹ�W���M+Ǎ��V�F��fUk.�����;Uo�^�9��_��1�l�xG�y,�H �5i��f�ii6�ԭ<��I�ŵ�՛^�r�Ycj�<0|-�tޡ̮!57:}�B>�ϵ���U�=�/�{;��1�q�;[Pd��g+7,�X۰��{�K�d����*%�]tP{�7}mA�%蚫��Uk���dE<�� �hk�V~T�}�#q��쨅��Wu�����DN�~�^����Um9����y�V�]���(��,��Z�F�I�za�a�r�eЀ�pL;���@Q��&��_U�
����%��5ļL�	��h��*�ܕ^r}����I(�'��^���p���N� ���2�,���;�w�I>�S�Y��qj�d��*n>X�&�N��ͮ�U�*����>���b�뀈�/>U��%A�T+[%j���c��� �'.�]2' �ߥ��#��[=Uc�ផ[rW���n��L���<�%�5M�ɵ|��h�@*!�jf%[���[V!t����L�f� ��իu7D]�yNM�ު�gC%V|L?wXòѸz t����
�5-m�x�QMU�b��;D���:\{������;'{��_��+��[�S74*�3��$��-i�.��yIZ�ukl̽�]{�L�ϪX#�ql�n��rh[@ꊹŧ�^����o�O�+N�I�q�j{�]��Ž��3`�{,s�W����W�[��G����2˼�s&_=��~�=o��bY���*�U��;��Wӻ.�"SnM����� �H�+�:JT�1��Ԇ��^�(4ڽ�а�	�q�[Ǌ�L��.Ɯ���dB\��ic$Qm�|�����s�n/�I(ڎ�dW%#+���S �K�q Y�L�\�w	���'g)R\�n͠�t��R�] sr��YU�ջTܲ䘻l��N���u�2b�$���:��h ̓�W7�n廞�Ķ�/�y�4�N�yѫ{�ɩr!�����љ���_YoM�(��Ox'w�%����O���}�$�U6��2:���vs���梬pjB/��5>��\ο�r�k'Rn�@u@ �玥Ԟ���(ż���$�}��Н(> ^;kT�{-o<]�R:��Y���x�������m�! �f�R])׼<yl�7:��vI���E��Ci��v�,u5˦	������������ل���%�<ʂ�`���g�u]�69��U�W�����[<w�'�sN��ު�-
t��v�)�׶ß0=�eC����C��8~yU��o���KPɌ�����Uv�і� ��H��}s>��?}�mC��[�]K��^#�EW;��RI��
����ftD�7�;ha>��ʜ�х�S��?�G��m�	}�8Zxpڅ"s~w�H�,`��:i��RI���1$F�FA����Za��w�����Vz��oһ/KM��IF�m_k�=�2lJ����Ƴ�vN9y���WOY�xu�F��\)=#%�y����Y�nଃl(^<���+qeVްU��p_�yu;������%���;�)�+ڡ�#����0R����)l����I�W�0�{��}����5L���1�#݁��b4�ՍSZQ�e}<Qژ'1�=̷��f����˫�D��+%�wfl��K:ݧ� "��&�9{�JE�&��� 	�( ��	*�;��u�����@��"]��v����^�����2��[����h����j����*���;kz2Uuė�x�i\��7{�����v
F�R���	&�hM�ק-n�G�z����]�	7X,z� -xy]��\�9���]�\\��϶e�j�۞�Z�P�yB��>Q��
��B~�CS����9}7#$�VU*�coۨ(�c����4���*0�X�>#�Ե���wݵ�z�Rdn�Q���KmQ٦�=��-7�8��E'���UN�]�ga�'���R^jlsk)�VJ����Ч��2�:�iG]S~{�\��An�_���&٫�K�d�×�a�7v�=YB�':h�$��nH�i%4k���>����#�י'��C���J5:�ݘ��L��f찅����+re�M	\�f��U����v�,�$�4�a�ۊz�<*�3�5弣�]ػ\�Г|�&IÞ��w�xu��9L�uQ;�M8@�S�����{�x��� z��\�x#1ɹ��bn�qJ�O4i�,�l�ېa�Y}�@wI(F��^��s*�.�YӪ�&�����M��UΞ慻��7�>Qi� >�mWWs���W6�Ց_H�ݳd^ï��omfCYj�dO�鶙E��^<��|�vvs�3o�r��H��P���hq������ �3��DZE���y���4�ݎ���]��/J�S�ˡ��d��B-=ɪ~�r�x� � <T�9�f��6�rΝ�Mj�8�k�ٓ%;��q~�ºwu�Û�z{ޭ�v�`�:����*�ed��L�P��R>�w���i-����uP�*L�z�L����z!7.��
(��Ww&��4xçU�a��[ʖ�IX��Y'I���)���5�f����1
��H&��7f�zY+�.b^�+"�2������*�j�rF�m$�I��9sl��b.�kq��:��YS����fn.���w���C:,jK"7���D�4�(�L[�S�`x_+s����:��n�]�J�.LӒ�[��BTȽ��������<���~��ׂ��k�-���6{�2�ҹvӛ��Tw�ݝ��g�7�J&u8��$��:�ߟ�K�XY"�້ֆ��26��ue��#����А�X���:��q<�Im�ljldj��8�˽n���'D 5L�.��5 �a,�����65#[��rӱ��۾S����cy�|@�lh#�(YcF��^�e�w��]�t$�����J0ݏ�TT���%��_|7� �r�^u�3�a�۷��(�f۵~��,����� ���V�wB��LC�1׽�"���xP��  Xf,�1�4$���\c�W�M!Ԣ�wM���+�u�RN]KM�;jD (��wbf���Ut���({�$���U�O#;����֌ʃ7=���1�(�䎯�tssN�>��su�N�{�&+<wSˊ@�`Z�׼�i�dp:�?y�G��|t�&�*,Lj1�З̙W,d[�m�܆-�K�-�E�c�E�����d.�a$n&l��D�M6�J6ܑ��,+F��Xg�p��	R�nt1ګ\���B�bS*�)c��z-�8���f��Nrk-l�ب�j�.�q�/�7v���5LV@\��⸎�"t8�J�Q��_T��5�.n��^�53��5(��(�B"H ����ӺS3����E��<ͻ��
4E���2ǽ� �X��^��;k�c:��2�\��f�\;��$�����j2	�9��*�"dp��u��+� �Jmr�O���1�R�;F�\�*rIױ� �t�P�B�F�a�A�#�Y���w�>�r��C]�p�N䝰�H�>	��q�û1�Yiƕ�ǔ�䴤����Q�� t1�i;ϓ��*,��.&�����O�iy��t<���nR�H�-Y9�u.��6|�Ĉd��Pex ���u��}1$�(����kO#Ѳ6�8Σ�h�ƌý�p@I�8��l�`�4�F��EգyW^����j�5�1
/#����r�X��Q=�h)��b��@�sX�;����׬*Y�"�� 
um����k.U��6��Ցj\#u�m���W�&^��8.CR�A5rAʽ�7R�u�%���ՐI&d�nf
ݬ��Ykj����#I(ڍ���K<�ln�0f �ܺ��Z��>Ǚ4�{�}�{5#�LJ��Ћ��iڔ����%�K7�ؚ,rM�>��_����l{��CMB�6��9Ʒ_;�n�~+-�]�'w�r��C x#�:�i���ͧe�<����LW��"��A��[Q�˩����9C��䚜����q���_�gE;�m����]:ё�{�ݹʛ�G�0��<.��{��(�Nܬ'^�P�GuҠ��_c�B3��� ��Q�Rхd��p��I����t��Ƈ#�x�={��κ��c�Q�W����t��GLk���F�Ώc�a�+4��\��b ���r�	�`C�l��e8Xi�Y<g).�e���Y�n;Ѷ���b�K����Ք�-���+������i������<���qY�����I�5��ʵ�"=�'W�e�C�K}�W��P��[&gNX�����Wwmsj�*֗G���3��[�Im�2�����,�໅�Y׋�f�XY"��a�{�l��n�����Y��Ԏ����fvy��[���~���F���$�I$H(�2��
(�pN(zA��_pn��SX�i�J�\Da��@"J�X%k(^�njZ�a!QF�h���D`h�
��b����c[~���;�H%x��/X�ߨ�<���+�� Խ�"�L d�ږ�
��@;]��?G��j�(�#�@������F��!�A� P��?c��9���(�9�SĀ���F �)u
*�W�����ýF���f�ߜp{�� 8�͎��7Y$������?�o�Uh�QIZ�(�젉�j��0����Z�ٸx��=F��QDv8^N���W������1��@�݅�`�� ��p�?HX r<�G�P����@?P���Qm���>�èN������<��Fϣ��w�Dwx�><P��y��t����C�` pE�{G�{߈�*7}�v��Z	@���S�UO �*"��1hR�`&�UE
WF�8��B�6�U��2�71OU�n�9.=^�w�E��N�S��p ��_����N�~\�U<zRt���=J=�5}"�"(�� �*�� �DQ#�6<|��ud�����.����"��D
+Ǫ ��<��/�T���m��N"UDy�7 챧xpYM��� �
xi����@�Q�^rG�`��T� kΪ������#�������\f`'�B��! �b	�B��]��BB����