BZh91AY&SY3��n�_�pp��"� ����aw��                  ;�                                            9          ����@   ��@@   @@�
1�����` 6V#T,m��� T��T��Z���Ucj�Wp          uT��j�V6� ��� 4��MP�5U�UJ� h�X�R�����ԪU�5J� j�V3T��j�V3T�bj*� ���P�ԪU��T��*�           f�UbX�UXکUb�� 6�Ue�Q1�%YQX�B�  Z�%U��J��*�P� �f��0�6��E\  Ƌ#UU�X�N�           �����,mU-X�Ы� 
2��+�UciT�  ���ڡch�cjK-J�X �J�,��cjX�R��  �R��*���ULmT�cj�`          U*�a�U��U1�R���` �R��*�cT��T` 4��Ҫ��U�UL  �E�Edh��j��X b��TS1uѫ���<  ����UJ�� 0   A�~�*�4�!��h�   �   ��mUJFҪh�b�@ 4��� L�h���4�@�G���zA'�T#*&@4   6$m��D�8'L�9MZ�j��j�Vyi�9o�! ���Ȅ$�$B'H8��Z(}$H+��X��Ҥ�Є$��tH:�Wݾ�W��U%��d�E�R�Uf�"E�c
j��ZM�;��΄ܵ�@�P�:l��ۛ�F�4Q�f��[�%��h�� Ի�n�4�m�j-�D-�I�\�I�-r��S4IB�R-$��6�L��k��$gPUӚܷ1ڹh��X��*R�Tʔ���E��N���-�Q�1iRfX�-�h�Z4Q�c[�����E�1�T��E�ѴZ-�Z-�F��\��]]�D�k�F�ķ1љe��-r�Lܮ�5F��h�F1%�E��TZ-�I��Z-�I��Z-Z��Z�Ԗ�ELM����0H���	Q[hU�R�m���L�d!kX	6*���F�fK[2�ʙ���#E�ѓEAc�f�RŢ�]r�f��DՆZQ�E��h،�6��RQ���!h�b�Qk��h��F�l���h��2�6d�l4���E��6$�Z53Qh�Z-0�l�CZ�A"1mm�X��s��բ�b�We�%w]&(��R�m\�ZKE��h�Z-���Wa�E��h�Z-�Ih�Z-�E��h���E��h�Z-�Ih�Z-�E��h���F�nZ6��E��h���E��h�q5�E��Z-�E��h�Z-%��h�Z-���$�Z-�E�ѻ�\�Z5w]h�Z-�E��h�ZKE��h�Z-��Z-��sn\�Z-�I�W-��rѩ��h���Z-%��h�Z-�E��Z-�E��h�Z-%��h�7-�E��i-�F�nZ-�U�E��Z5���h�Z-��h�Z-�E��i-�]�mQUH�Z�h�Z-��ܴXŤŋAQ�E��h���E��h�Z�Z-%��h�Z-���i-�E��h�Z-��h�Z-�r�h�\���(�]+���h����9snZ-%��h�W5�E��h���E��h�Z-����h�Z-�E��h���E�rܴZ-�E��Z-�)�*J��h�%�m�UʪM�EQZ-���&�E�Z�܋�1h#F�pŝۮSe�n�m���H�bH��B�i$0Ț�4X�Q�m����v�E��Z-�E��h�Z-%�v�Z.�u��i-�E��h�Z-��h�Z-��i-�E��h�Z-��h�k���h�n���h�Z-%��h�Z-�E��Z6�κ����h�5�]٨�%�U�E���nZ-��h�Z1b�h�Z-%��h�Z-�E��Z-�E��h����q���٩��ܴZ-�Ih�Z-�w�Ţ�h�Z-�Ih�Z-�E��h�I�r��k��E��h�ZKE��h�Z-�E��Z;�\��1˰ܴn[��E��Z-�E��h�ZKE��h�Z-�E��Z-�\۩ۑ�����E�Z�h�m˙4Z-�E��Z-�E��k��E���s���h�Z-�k��Z-���K�M;��sSM���h�t��\�Z��wZ�E�E��-r�i-�E��h�Z-��h�����h��֋\��\�Z-r�h��փHZ-�E��h��֋E��h�Z4Q����h�Z-�E��k���E��h�Z-��s�-�E��h��֋E��h�Z-�]�h�Z-��5�E���E��h�Z-�Ih�Z-�E���R����jŪ�Tm�d��Uͫ�(��Q�۬	MnlV��j�جnl�mr�b��i��q�ҴV��Ԗ�*,mnUN�2�J�۶�j��\ܫ�W6-��֨�X�m�j��j-�����ۛ��[�l��髳J4U%������ֺs�u��4��][.��Lқ�\w.����p�].���m���*�ܲmr�͆�m��
�Zwj�s&��b��i7.u�h�K�w��b����!��KF�k��\�ֺ�EMΎ�'m�L���\��E�l�6��r��k��ӻwv��jw]�`Ɋ�ۊ�nZ+���K�]����ѴZ*�̹�6�͖m�7]wwj墮��[�wm�2˕ҹ��IbW6�u�!ȧwM�h�[���F�'-�ˣ\��*�wj�$�t�k�E��-�\�Z-r�6�Ep\���Q�}�s38?��YْI$iG$�I*��RR�#� ���k(U��#b�{��Z���W���Ywt+׭[v�x���	� �ø��              m�. ���@�؜�  ����o�l�]��.k��� � U    �U�����
�       ��     {lp�͠��n�n�@ ��燁�1��( w �����eS��z�\mn�  ' c ��ꀜ����ez�k��e�N ����	��8@x x8  '�k�  �W�ͻ�9���ݣ�of�ɽ^`|U��xs�Pw^�{�ʨ' `n���x�t�{i^νU[c�r�  '=���V�����u�P�1�T�=���	���vh  N ����	��8@x x8 � ������1�p��T
�P	�Y�y�  ' c��P �͞PƜ�� < < �6�p����	��8C�  C�   x ���y�N ���x8�a�yN�C�V�  ' c ����<m�����c��pSc �8� ��.���/������.-�\�Yuj+2��	�� A��` < Op�a�s���	��8@x �0-t  ' c ��� ' c ����` < y����4�`�s� <x8�l���c �T< ��v�;��з���0��I�* 8	��z��k��7N��Lbv���eu <<r��������ov�]�s� ��woط���]vʀ[h`    �P�ЪU� ��T��� �� �m�  =�>����� ���ۉ������
� z��	��8@yTܪ;�Ǵ��\��|��^b�P8E^�o��~��U��S�y�  
� uiwl�   � 9� �:�ۘ�0��l 7�U��s   T  fQYB� [  �ٷ���� �            x �v��T�i����  �p�� Pj� �|���u*;3�sp0VM��� �m� =T ��׺��M���6��U�XZ����*gǳ���+؎�k��ꡌ���A�zN<���
{��e�gb�    �b��@ù�     *T�    @    T      �    *n� ;v�@ wTٶ�Lwq��      e�    
�
�;���  
�  k`� 
� �    � Nm�      Up �p�'U   m�
�Tl�n   *���7Vչ�  zd     T� �*����l  
�T    @    �    f�t{ �P m�  �� ���ߠ     V��UuYj����o6�I�[�gNh��]�^�ӕ�T @  +(  y[��� u+�{�R�����Å���s�^���� ��n����s�*�*����W=��u7��٬���<w �  J� ػ�T��[�M�o3��֩��    Z�V��m��wWt��t���۟���9�i�lT�X ��OM�q���ڥ]ޭ�������>��/sSc�֊����l�����n   ` � ���(� 	��m�^�ou��Ta�����eܫm�1�p���ո�    +�P    ` m�   �V� �   ��  �zT  &�  Ӹ�m�n�                               �wu���S�TU          }�    �  �                                                   ` P            �й�                         @U��       �   *�       �             @      m�T  ��  *�  U  �  U                                 �       ��   6�   *�     @                        *�                      m� � 
� UT                            
�         ��             *�P  �TT     � ڨ        U                P
�         ?A�      U             �           � �U    U 3l1���  ��
�U �UUEU�                 � n�                       �                  �   ;�                �}    @   � 5P    �         P                            
�e��T      �>�     ;�                      �^`���                     �mmWD @      �>�                           ;��      U6� �@                   [              +�*�f@    �*�         *�                 ��    �`                T�                   *�U                         �                            T*�                         @�o�~�               �     *l��  6�  *�   U*T               o �  P�   @PP�    ?A�                  [9kmm� @ P   lb���      �     �          �}�_G� ��uP              PP     5H@T���p����N�r� � ���U�ҍ�  �            
�       Q� � lomm��{�wۊʧ  ��1��  < �܉��8@x x8{���N � @    ������1�p��*��:�  tӤN�5��� guT����! ٺА��.��'��7b$�>x�cwg�ᅜ8tޯ{q�-���-lb���x�׳{�G��`  >u '<ۻ� �@  �f���o��<�a8֞��	��jwy�3�w����X�w`����1�p�����Q89�8Ow
� �
<� N �����*�{q��N� Nx�' c ������1�N�<O<�F۽��
��;@�;�lU��9Y� ����{Gquf�� \[5mmER��d  ���Vdy���W-U�5��²�M��� *��  �U��^�
�تm�V� Ude�  *��  PU Vuw��l
�5W��:�r5^�G�<v/(9��s�uh���{ut{��+:��z�l��` U�UN�:�z>�	���z�p5��cw�      *�` U�T         �  -�         U    � ;�      U UEP          QT     @T  
���    T P   �   ��T{�   p    ;�  �   P  @       ��P`   �    UP �     @T   @ بU     P�  P        
�          �  
�*��
�  d  *��   ,� � <   �U    V�mV�f@ @
���@c 7� xm��e�  �6��ϟ?����7���2���w:�/l�گ���0T˕�U��La��]�v�v��b��Њ�l\kr�{�.y�*T�eP�Sm֭��&��z�ws���>(�� ��  *�@P   �;��*���TGp[j�I� �j�@�  � T 
�����˘�m�{�ϝ�v��m��m �$��i"SI���Z����mUz����T�I0K �m�O?�s&?����f?y�����?}�^���z{~=���ϕ�����}^�YL����A�2�	9$I6�9��O�%�G#����B�mB��Æx�Ob6�~�/}���h�e��nH�	G*��'7.[�y�y�����KH~����pr3-�Km� e���P����8im�rjE<>��2��Nue���a��x?Q��NHۍ$�A����)>7���O�%�G#���B�mT��цx�H�����r\&8�"4���������=܀`�V��m�PU^��R��K(�E���}��ܽ�yHf��	�O����?P�p�j������I��፸�nE$!�CO�W"��mC�y��e<4�S ^�p�x}x3�e#����d�ܒF�n2)����e3�R:|or9K"�xK�
G<?y��0ک�Äjq�m�H,3���:a6�f�0�z}���)�Ρ�8�"�4�����B�Ý��˄��G$�$@���奘)��:k�إ�P���YO#�����p�xnU�׶��޽���q��`�JΧ-<�PT;���UWu ����Z�0TNI	m�#1��{Ŗ�2)����e<�)>7���O�,�x`j��nIMHܒBK�
a���\3ƚGM�n8mC���{���<��R)�N�m1�
��!-��`����p��ȁ�O�K0R!��tב�K6��=/x��G�����Q�ܒF�"�
�8E<>��2��Ox�/��i��oS�T���{��Y���&]eD�$�q�����O�t1L6�~�.�M#�nFmX~���{���<��[�EQ�*�v��hj��ٳU� a�^�U�R����z+�g�#q)#m0��pӄte����4�)�if
D4�Κ�6)f�:E|5���	�#q"Tm���xi>�>@�\?S��ѝc)4��-�dS<#�-��y�R:sȡr9��[��r9K"��/`X)4���C�H�?S<i�t�m��"�¯�aQ�!1��m�$�C4���R<p��eƚF;r i�x��(�R��B;Xhcm�ے6�IȠ����U���8}L|�S�x��2���ze������+�D�	Jw��=ɶS�l�܀;��*�t �6¨*��[R���r�QT7��)�t��ds�������y�d>>"\SƚGO�W���m��J[��G�m�#�C4�������(~4�0�ۑL#ǆ粑!aƠnI#n(�C4��%r()gǄu��e<4�S T�8{��e#���T8�!#����mAL><#��S�H����#Ǉ�2��pӄx���M� �K�I$�|[9O#�AnFi�x����<�3O�x�8|p�2��M#i\8D�$f5!d�#_��O���x{�y�
��q��ǎ�p�� �ٞ�l�wo��p�+&ֺި�6�z�-�^�� 2�
�
���w;�=�N�z|n����edT    U �   <�  w*���w�*��B�cl Pp
�P�*�� 
��EJ��T��w@��l�/N��wm{�I�wN�-���������PT<U��
mT��wY�^���dd�bI:a�ˣT�3O�W"��|xG_�VS�Hᦉ�%8G��Vd�#I�$�F1��ze���у׋)�t��dső���	{R8i�^7LE��Q9$%�L2)�ǄO�x�H�[��G�m�#�C7�ļ�������J6�qH�rZ����\�a<>�K��<3���
p����Ur�~��D�$�q��
�ㇾ���R8i��dS����Ŕ��GO��G<Y<5�[{�����{m���l�9�M��v��w W��@w T� �ܽ��̓H�JI$�D#�`�pӇ�:�P�`��� �#>�a�����)�ުg�TNIM��6�"�4���ʅ#�;VF8E<>�HpR!��ˑ����<!�����H���p�8}L|�z��)���α��s�-�dS<�y���<� �Q0��D�mƊr:�z�9!���O���P�`��x�H�[��P�)���m�~Q��F�M���=�����N�x_��R8s�d`ӄS�o+
D4�����jH!~%;¶��m�V��� m�lUU� *��ePU�mOw;�.N�2�PRͨt�;�,�����c��O�Y�2��Nue���a��xz��[䍸ے6�A����)>7���O�%�G#����1L6�H�V)�M#�\%��Q�ܒI$�G#>�a�����)�ޡ�8�"�4�C�#�;VF8E<>�IU�
m��JF�,�CO��PRϪ#���)�p����C�S��u�a�:�{>u��F�6p�L4����e3�R:|or9]��G�����,�岣�Ze��1�12�q#RT�š|^� ��U^�b��AYK]nn�p�D#���m�Cm^��:D�f�0�z}��G��i�P�b�Np���eB��֯I*SIC#�GR0i�)ᷙ`�)�����j#���)�p���'�"���Lo�rHKm�1��pӜYo#"�i��*��<���܎Rȧ���#���OVݎ)I��I
�)��:F���4����"��r���!�{�<'�S��!OZo�rHKm��,e3�R8s�d`ӄS�o1�0R!���q�)g���{Ŕ��8D%������E^U��U�n��Vٮ�H ��
�R��
�S�]ڛ�F�6ܑ�j"�^��H�:��FE0��:=�xr����܎Rȧ��%�TNIM��9"8)4��,a�a�
F���4����"��r���!�{�e�D�H�JI$�؄S��"���eB�Ý�#�"�e�`�a���q�)f�:E�(U�d�ӍĉH���xi6�1=P���U�c)���n6G�>>#��2�q
GN/���6�q��nG<Y�z-�G#���a�}�<E1Oi�dg�C���>'�$������yM����?��6:����ٹ <7���n�k���n)Rl���5���ت����AU� p�����1�w�v���:�͞6�-�      w �   �  ��� ��lwl  m�� �  @�
� }�`� 
�P+=m���n��c�<��
ڻU���k�Pl;�U]�PUj�
����=�]�禣�Bcm�$Q����=�LcH����ʅ#�;VF8~����
Fza���x�q)$m��#�!�:�x��~�����-Y�2���V�dx����22ˉ�Km�$��R��#���#�,�����p���,!|ϼ����)�M?x%)�#m�J� �S�C�鯗�e?S�!�1�E8|p���T)9ڲ0i��N�d-���$���qL�4��.5>G�C�u��e<4�k�'j#ǆZ��e?S8��kM��!��J#�"�n9��<�� *�q���l�m�(+)n�Y��2�)F�q�ڐ�	0����m�R��#���#�,����#���O��>�"�a�$ID��I>m�����F}�0����G��Oz���@�{<%����Ĵ��9$�$؎	�����z�淚{����o�c���-}=L�ّ�ҒI$��#���~���6�Yo|�r?)��xѷ��Lt�Z�����d�!��Qs�������Io9|.rs��b���)�a�8�ۻeV��;6�jN�j�m�p{)TpJ�T��NKڶTLe�[��3��~�Bz�淚{����B��*'$�&ۍ����o����~���6�Yo|�r?)�}�b�6�p��H�r#o/'��?{=G�^�������~�}V�=_~���ַ߽[��_W��������[}k~~u��>�����w�<����w�><y������շ����m������m���[}��ߍ��߯_�/Z�Vߊ����ϟz����޶�m�����z���y��#���>��|>�:��`-�Kq����׆��[�m�[}��׋η�ζ����ߪ޾��^�^���o�?���篾<�|kzV���������ַ�o����k{k}������y�%;���
�Owk7� ��V��
�l*��z�<�{{��`JF�ID�r<�~3�a�xn�sַ߽���ַꯟ��K������>v��������֯���7߾����ϝm�}�?}������IIq�$m���m�[}k~z�o�/���o���ߍ����׍����[�ζ�m���z��z�[�[��ϟz����ζ�m�6�����ϗ�^<x�x��Ǐ>|�x���lk{��߿����Ͽ��6�k|��ϋη羶�����oַϿ��~=Z�Ʒ�C�����ﰀ>����rG��u�ǟ[o�o�m��[{_|����ǭy~��~lG7P���a�C�.��\�dS𫪛-��rH�m��yN!�<h���9/��^j��a��c.���g��	�g�GSe���1\B2ҎF�-�&e=8�o7��*�qUW�ز�ՔG7+7;w�d��n6�RI$�f�8E"͎|O��ղ�q�O��c�[�<GN]Y�R�]���8�nI#m���H�H��v�q9м'O�S|%g��ʂۅ��K��g�ڹW��x��ۍ��$6����no�+!p�5���q�]���H�]8�/U�p���Q(�q�$c4��خ���p�|nn9�6����rK _n1;V�
GJ�7R�|�rHKm������y�##�&�����t��7�Vo���h���<ϵ$��(�����j7n�:��K�@�	�����UT��6�˫۽���T|�md |<Wf�<�r�mݠp[j�:���sܻ�ѭ�wZz�om�y�@ U   
� `   <  �  ��PU�VP �`�  6(� �  @�P *����נU���s�v֖��c�-Z��wmV��3��ku�A}��g׀+ٙ@w T�*��u�U]�b���߯�����~�#"��1nǖ��):;���)�W��`�)�Tרġ9$p��HYo���b�Z���o/�lb�οo5�w�^�J6ےH܆���7T�Oo�fܫ��ʲ���Ge�V�rH�m�܌��y{�v%n]3]�!n�k�/��msF��$��7�I"�����_{��8Ň�{S﷗�61m�g��Am��B�N7;�W{�yAk�l�`�ª�UATm��*��k��\�h6��v����u+y�p�oU�U���y�:�³���`��Z������G ��K�Fr<�>���G7P����>��ʴnr2)���c�U8�#ƾ�ێI	��$�(��)�W��`�)4�".�yo�q��6�uL�C�S�E֒m�F�m�iǟj�W�ݹ%�w*���F��ҭ..�ϳf
FA�-\�\i�nI9�����:~ʛ�+=��T�-<�|ͫ�h��dS�l*�r2���{gs<�^��T�N<��wUz-���UQl�[e���qm������N!H����Nb����H�Q�u{�p�|3�e a�t��B[P7$���n9��p�|o9���6��zW�"����V�=��ѽW�V�q��!$�=-��mIr`�a�?��)9м'O�S|%g��ʂۅ��G��3j�So�
��H��Ldi��[�窜B���r<�q_S͂`�8iD<]^�"��Y@��F�m�����>v�=P���sy3�m[���"����V�=�����dĒ��T��b�J���PU6ø�J̡�R���mn��[�L�RI$a�#/��f
FC���\NGt/	��T�	Y�&��h�Ѽ��k�rHKm���>f�έ���t��-���N!H����Nb����H�?��m%��"��B�WдX�^J�&,�y~�X.<vcʶ(�z:���\`�N��2��rH�m�܍��Wz���w�<�"�������Sị\VGt/	��T��á��%��Ĥ�F�Ȏn���F�;�)�q��T��Ի�M����r��V.3=�CeT�R�%;��:�yU5��s ��*��� PU�m�^k��h6�Jj���Z�����q���ݷ]t�}~�f\�������)f(�-�ђ/fg�xǹyy��:����c�^�l^��t嬂`i�"I�)�����@��o�z�๋�:ǽc���8.$dqF�m�a7#>�����;�}�^S1�r�rC�g�U�g�2̅6�m��.IO�w����=یwח���O<��Y�~���~��
h��o%]i�lf�-�qգ��ǎ�}�}꯷� �ٞ��m�����֠N.a��ԽnC���T�@nj�VPWsn��b�<����,��u�����      �   <  �*��Tp6�Tw � �� T� 
��  � �T� �__| ;�Am�Cv���ޝ/+x��tʀz�*�z�P����^��������;�Ͳ�K��M���M����u�r;s��F�{�R�^\b����K���m�$�I�G���7��Gj��w��J��/*r��Ѣ����iG�Wm��q�ڒC$s=cǎ��V�q����\`�]璫�sV�ӗVy�E<�������$I$��#���ł���F��#�!��O*n4\ii�銆�\v�����ۍ��$6�
xG���f�L^/��Ũ���*�,���⚵t��3y�l��m��0��<m66Ֆ��X 6ø{��-EJ���I��!H�IC#��b���4��[�W�:��[��o���X��1=V�i+��Lh�B[l�$�b�qY}���/Rn�����짚F��h�Ȏ]]"���-{"�4�I��(��3u{˃s�#�vv���\1x�~ʛP./#��c��,���To��HKm��x4�+WH��̕lLXO4�&��ǎǹV�q펛���#��/����F�7$R1|�6����
�����.جb�M��O1Z�F��#�#H��9� �أ�έS�;���U��;Հ)��UwUATm��w[e�].�ڨ܁�˫�S�w���0�[����ŋ���M�b����6�\^GW������I$���R)�G��bb�����U�1a������x���*��s����NFbIF�MŃ�b�y*���X_8��j���v���7q`��/���u��H�%�a7#�#H��&�#�xG��nJC6��1A�H��۱��H�R�hM0�n91��(�x<����`�#&�į��
���bb���U_�#ǥSy���o�$q��|䈶�r��uM�ǈ�⭷�ٺ[j�
�3��/w�6�Q6�m��3HGup�7�X<x+��U�b����V/p�c�*:Av�22ˉ�Km�$�Gb�Z.��SlLX>T�[�h�6��ddt�8CѦ�-���B���qBb���*m@�^G�,t�1X��\J��<,g%[]l�&H1��H�q�!��x���y3HG\aʞ�ȼ`�^o%Wt11a�U�XG�1m�I$z�q(ڒ���C�u&�=u��S��~R�y��]]پ�����u���z����7��*�*������*
�v��y�A�cRI$�6����۱���<u�ʛP/��'���,�+�^ǈ�'H�$�H�m�L�F3H�8z�<��
��Osܫb��Õ=ˑx�a��դi3b%&��iI$�*iUJ�b�>�i��.��ůq�h�����<�ł�K��:i�$���$8fi22:tX-���o�P��u�ʛP/��'��#����޶��H�F�!+���^����eu�k�ƞ�V�q�*{�+��z_�m�������>����><y�������t��|� x   y�Wګ�l��v�� �� Um�����x���v�m�� �3qQ�����y�۶�6�{�^��{�����O[.؃����[��p�������'k�u < ��v��0^ݯZ�נ	�S8x8 s���< �6���x8i�x���67���kP�Ͽ~����VکT�-����1����΁T6�� Ը�Y@e�   \��[�Y�N �C�˻\��U�T��������    � ' �T���� � V� /T��:쀪 ���*���
� ���w�܀dͬ�םh��Ż�����p���n�� p�n�=��3�[�wx��W���n䱜 ;��;��N�pm��8      6ʕ   �           U       ��       -� �                  �>���             m�          � T�(U ;�   w    �        U �
�       z�  �    `    *       ;�@      
�eP �@        @   �    
�    �     �      �  ��  �    �U�@ 
�  �P   TVn�om@     ��^P��m��k� � ��m�)_����˷`6�s��-�*���F��z�ԇps�YX8@~�������G�/WwmJ��LR;�UvѱSJ�a�s ;�����ޮ��l\�w�ׯl��9�t �   �  � �P <�  �   �� ���S�@ � m�ت @ U   P� �E����|����*;�7����U1��P�ª��*�� U]�ٔ��{�A��7#ls��H�G��α���-y�4�1u&�-xˏE��ؘ��+�@�⑸��I$0��4����%*����UԋNiy���&/or<��ۚ�/YQ9$I6�nA$��O�į��-7������)���)���f����e@𶵑l��m��E<#�xĵoP�:k�J�b�.<�%;LV1O�Z�=�x���H%�9$I�)8�H�8w*yJ-�Z.4�M]1X�?F'yR/#�>�v<�S�i+Ow�7S�rη������ǯP ��U^�el�Ք-��m����<�R�V���2;�c�V��bm\J�{�h��̕lLXs�����`���n�4�m��nH˒f����U}�dS�0�璫�a1i�U�U���|�i��B�%�.HۍF�a��L�
{mͱ1aܩ�Am��q��;�);���7���#�l�鑖\M�$�I1��uN!�x��E<�����M��\S��Z,n/%[�TJ�Hۍ$�pI�F������ǎR�.E�b���N�Ɖ�Nx3�`�)�]N�2Ii�"m��h��w��1w��� ��{2�C��AU�s_;��
���}��w�z��ůq�h�m��&,*yP_��tɤ3����a����m2��x�`��Φ��	��[ܩ��y�1�Zb���\J�xX'-?Ai(drH�F3H�8tK�r��x����د�P�<r��r/+��J�ta����|TNI	m��`�<g��R!�vq`�^#�-�՚~������F�sp4۬(�I��9	�>'ǆ�#��>��=��R<w��G�x���l�4�E�W1\%�!.�׻���]���c���ª�UATm��*���G+֘�I�/��a�f��@�C���F��᛼ϰ���	w�������I�#rI��$c=��R8wy�c �x�o��F�Gp[�<yH�{��0�� ��rH�IF�H�R8G��w+�;����H�bP��S}т�xx�)�<����j$�2F�RI$R$��Ä�\�%ǅb��nU�+9O���a=>�����ɩ��NFbIF�M�dx����'j�#������x�"�-�/��t��u�rn�|�],�״���s��@�wUz.j�mYAT[;�������uWu#m7#�@���Dr��<xwI�>&�N�̌�� -6�yj����A1�ˊI	��$�G#�<y�g���ixM��\S�o�ܫbVr�9w±x��"�l���q�$m�ܙ�6��w������N��<G��0���<D> ��:Z(țd�ےH�r׉��O���	Y�!�&�X/>pr}���:@軚aI�#n2T,�#�W�x���� ��Vx]�#j�W���[�p��a	�32�̭껠VP��i�k�6)�U��V@	�n�M������]��Y�5[� ��c�Kc]@]E �p���Ɲ"n�M�Ck^.�󺀪@    *��   @ �    UQ�����PU 6�T m� 
�   P��@�C�w ����[�ٛy��x<��kdEV��z���J̪�*Tiܜ��S&5rIl$�摄S�s��L��WO���dx����'j�#����E�K}���m��j0b�H��7v�eG�����|%Gy�7�a<>�'�ک{V�!-�$�@��G�M�Z�E#�G7�X�b��:�\,8M��\S�ؚ*�����l�C4�¨�����w ��ۚ��xlc�=�g�(�4(q&��IpHǔ�b�����{����g���繷L}(!m�La2�n0�D�[*�k���ª�Tm��n�9$l�Tq�Km�$;y�ɯ�t۱ۖ�G7��%�9�m�@�`���[��"��BZ���m�Cr��[��wٻ�[��]�G�j�b����$�nI���y7T�Sñ{��cޞY�wos]�h��.)�I$�C1����-У��k�6�v����/I�50]d(��$�q�!�M��4J������+=վܽ�]��n�Sy��J��r45�n��m@�{���J�qUW��[-�eKmwUK��U+yU�J����f;��C�=r�z�N�r�Q譖�qW���P#}$B��$���z�/�/	���梇M�S<�>�cwRݷ�.���$m�ܑ����{���d׏j��e�[������z8�bub�%��EI���{�w����z����b圣�[-~��6�Q��A���{��׫r��/���C]����3�<+E"�e��a�}�ue�*��� ���J�P� 
���w�.�j�9�����y���r���.Z1;���YyۈTJO$���jH�jY�vz�u[ݡ�x�\�<c��c���Nug��Β�Q�$��Z�C���7x�S8����6���T���0\`�"☬nG�㍸�Ic<4�w�m����,{�l�q�����,�c�1L�O��F���ID��I$�e�Z;:��,\i��6�'8�K�
xi���'��p����[�so+7��t��^���
 6øUW���w*�U w6������uQ���xE9�n ��Op[ł��M{nm�1a�q�W��)��fbu�i5#rH�������<t�ELo*m����cܩ�H�݇��U^�ç�K�o�RI	m��	g#���¶Xţ��Ͳ�ƞ�ySl�^"����O<#�4���16ܒF�0���äp����xE<�tTq���ȵ�dq�o\S$b���Q��D�m��H�i���Xf�Cp�N�)xg*cySm�^9c�Y��Sެ�n����3	�C:�:���R�����<wuSl�����؜�:�ۭ@;@����؏���UE���sn�<�s��o�ޕ�Ul���w���m�      �   �  ;� �U<PU�*��6�  l   @ P @ �@6�� Ke��UV�l��/��,��n��=۽�w�@P�U�-���VS�}��k�������ؒI�I9��Ǉ�� �3�gnj��Z;:��,\i��6�#q��c�D�NII(�@�Â�zE�q��i>��2�Nu[�:D4���`�qS�=���cCm�[���mf�X��E=&ق�iŔ�Cp�UMR��4T��ی�9�2"'aJ���������5���<�)�,�y
W�Z,�l��F��]�g�`��m��q�$m��y�3��䳕��,f��^�{	�Nz�ҭ��:�Ŧ#�4X���ӌ���xᱺ���W�cֺT;�*�J��R�*�ç0��T�j-2���K����*{P_8Z&ilqe1P�k�feP�c4^S��)5$m�J���y���<h���4�n�瞩-1`��R���h���iät�\�$/���$���je԰L���*m�F�}��mЙ�4O�d��C�LZs�~�l�2�=�<(�	ꑸ�nF���OO�n�`�8���K����*{P_8Z&h�8����ꜼȌF�jI$�����OJ�ʛn+!1x���7a��R�LX3��)�p�Y�!��31TU�s��V�[�R� ��U^ɲ�x @ʹ��켁UU�UT+e�ZS�m��3�cܩ�)�zr��e��6�%W��b�9ň�4 q&drH�F3OӝV���g�7�i���/
^��H�gx+{]C�i�8�D���B[m&�T[�}�ʡp�h���ۊȿ�kZ�j���^����__�������������p��2�-��&4��F�H`��[�h���+e�ZWuþp�L���*m����!�3{��8t�=�l�D�m�"��2��P�:r��1�xF��ᔘ�c=i��L���xR��2F+���?{����]-��t��Kךލ�P�j���Uj�
���Tx��J8���#�I$�˨t�=;���b����ʡp�h�����d-#Ǝo��O�Ϋ���z�qI$I$�f���M�,��
W�Z,��V����u|�`���T����+�6�ߣm��m�H<�Diç�m�Wt=�Ŧs��f	��˭�&+ʧw��b�C�k�@��#5$f$��"b�#��Of/�-4x�YLT7�yT.�p�T�8����j[��Hۍ�#l&��<#O:��=�Ń0}��p����8��l��N�]C�iӟ24�ƞ�	�F	$��d���p@P� ��T��T��-�Kj�NݹT.���w�������,c�Y*���&-3��%[0L͎ñͦ+��NuR���������
f��2�^�qL����Sً�D�'SƸ�^U�3EV�#,��nI$�c���8���V?d[0L͇�3�6��f���ht�{B�<�ät��w����q�ڒDT�8X&x�or-��}���,c�Y*���&-3�_�[0L܋���i.5�H�i7#��N�<��/
^��H�f��ҋ�D��M#��S��$�Ɣj7"JF���QQ�W��p�Ŧ������8�����{����8@r����2��`�w �]5wp�Vc:qU�ٵ�lw [      ]�   <  p   �x`��� �w   � � ��*� �   
�� � �֪�y�T����S��l�����l;�U{(
�lF���z�vkyT�U�t�Й�4U�yS|���쩶H���z��b��>�R�w��zi?	�cID��I$R1�xt��f�u�u�ʛb���B�o*���VJ�V�#��u��	��B[l��f�	����,��c4�ȴ���u=%8i{L���P�xs7m�ޒ�MHܑ�R�4�i�V̈́�t���yS|M��i���6�0|�iM�p���1�ӊI$JF�m!�O�"���f-S�p�Lg+{�|,8Ρ�.�F�:t��5t6�!)>n"����W*���z� 
��*�t[*�l*������j^����w����\,=ڭʶ`��Y����i^9�Zf����N��B��ED�H�m�ۅ�]C�i��ta�g��NtZv�f��o*o�VBb��}�W����^��-	G$n%$���l<E���B�ø�E�q�*ك�����1�or�ؤn7����"�b�j��&ۍ�dDiû�^"��j�!�p�ڳ�e<?s��PR!���-�����P��P8��l��m"��,�v��J/�-4�pYLV7�[�\1�"S����CH����I���^��iEU7m�� C��J�P� 
��w-�K^�C�`�U*ff���&f���QI��a�)��Z,��V���5�	��T��o�6�n4�nG�C;��B��DF�,b|�%Wt=�Ŧs���f	��}���0��R֞��M(�-��H��˸n�/\S$b��S�Q|�h����b�������yO=
�j�n4����yuN!�x�o�idi�S瞥6��fx)\;��h��/%[0�7.i��Lj�I$.<�����T����+yP&X�'ʲUw-�GM����i�\�R�%���������U�ع�� *�Gp{(
�p m�U/u�w��2�U����M�+�Zo"�2�^�qL����OiE�f���)��q�+9���iԒI'�<$i���%;��.��L^;_���"f�6�Ԫ�����;�u���q!�I$���l��[0bӺ��8X&3�T[�ǽ���,c�Y*���&--I�=
�$K29$a�#��i�Qy���N�i��Lˆ�xR��2F+�{J��#ON�ޑ"-�B[l�"�4�7��V�f��o*m������*m�&n�瞥6��f��6ffI�����xn�U*��w��l *���U�EQ�ARQ���kS350�2����qy*ك����X����T[�ǅʝ��8�t�OQ�ܒ$�nI����i7z3e_.7"�d;LV3N��E�e�@�*��H��Ǹ
T���d��"9�G��׀ᔌ>���<i��O��.�w�7�W�ݜL[N)*�"""�j���x��}�{��S��O�-��r=[�^�cm+�m�[���;����ɹ]ͼ窶W_e���n��&�k�z���$D��q(�-��r<��u=��' lPC������Svm��$�]�ùƪ��`�^��r�����ˀ�������U��O�<�z� 6�T     �  ��     ^� m����m�  �   m� 
�     7��}�߿@�v�0�ҽ���"��[{�:�ٷ߿{�ߴ U�Vz�J�� E�Ӻ����d��ͶQI�����' ����^����S�z�n�{�w׃�nH�RF�m�i�W��w���m�/K��އ���~�~w���\22�)"[m�rG�w�C܊嵩�^��W8���Ք�p۷��s���Tmƣm�q��^UU���^x}��2���Ӕ�HG�4���$��nI$�c���i7��G��8ݎ瞥i�X�ȕ�p�W�%^�#�m�Ii&�!1�$i��v�s���lڶ� ��Y@� `�%!�($%F�q���%2��S���ʛb���r�u��8\�d��C�L�����f��:����q�ܒF�q1E�+�xo"�+!�^�qL�����f��S�Ƹ�,Z��ģm�x��ç�Jwyn��L^;_���"f�>y�Si�`�B�Lպ�H�|Cdƒ�I$�H�c4��G����1�or�ؤn7йSʁ2�1>U���a1i��b&e�PLʩ�U*قe�_vC-1X�=i��L���xYM����*{P_8Z'��~}�}�&��+�*^Y�<��%W���m������[cl
���m���MHbI��0�0摇uw˃y�"��W�M����v�eM�D�շy�#�O�P���RI	m���+L���h��^J�`ţ�\�`�η�SlR7�\��@�c�ݹ�����nI#rD$c.��#��Fy�f	��}���c4���-2���N�T�Α�vq2�*'$�&ۍ���D�9�,�+�q��T��3E\7�6�VBb����6�7b}��5	C$n%$�H̒�H���.��/Sp�Y��m�1i�i�8X&3�nU^�����Xd��-��#6�m~�}��*V^�:y@P� ��T���AU����ޗf�m�W����������~5Y*��������*قe�_vC-1X�=i��L���x]����t*��Kr6Rk4��a���S.���`�M1X�k�O2���`��M����]���]�Ӓn4S��,�{�wy�Si�2�N���<��m�1h�[.���>���d�m�rF�M��F�}�<�>��yS�^�{	�s�:�i��V{x�������ZԡiEґ��3��<C��Ҏ�ۛSQ|�Y��C)���\e*�ŋ��{!	��q4P��d��F&��[*�^�T�V�<Y@�
�m ;����#�ƒP�܏.��4�y������M�|�8R�K��Z,�ǚxt��ʳHQ�"��$�H.���O��ǚC;��B����4��5�귨i���Y��S�[t/��6�m�"��pi�OO����L���4��G>W�E��{��+�qYط�F5$�I�o�<#i��y��gݏn���q��z��g̱��+�8����N%�I$���l��4��zZu�q��u6�#q��ʞTQ�"�Mbz��~�}���ڎԒF�;��\�ۻ��@� ��eKon��:�	�  �=��ۉ͝`Z�0�[h< ������u����o��ǧ���%z < �����[hx8أ������ 1�p^����<�=Ľ��.h���E� ��1��	��p ''�8@`�����yl������T ��ud�Qn쪁T����l�UOV�s5� � �Ul�  *믝J�m��Wn���ܹͥk��H9h�5e�m]׀*�   
��M��TT @   l�YU�ClU *��ʪ �� �  .ʳ|�w� �����:����l�p{n�l�N�0�m��kd�/,-���3-��J����=��Z<���p�Aӓ�¶@�      �
�   �U             @    `�    
�@ U6ʠ                    U@             
�    
�  @ �  �l� �w    �    p   ;��    ��
�T     @ l    �    x�      � �    �  6�           
�        *�          �     
�T  q ���   Y@ U     M�  �`:�d�d    Aυ�U ����   -�m�s:ۙ���)�a{7���U=J��V�cw-�S2�b7��kh���bm[Le��p�f�P.clU[j��.�u�ǎ���L2�^����       � 
��T �   d*����@Q� �� � �  *� �*�C� U� <m�A깛 0|��͢���g'�t *�ت��*��l*����m����Yw��UMUT��U*ق��/�!���4�&�-qYм)z�1Q�T���q��s��"�Q9$%�̌sHú������g'�ySm�d3�ǷS|H�ݎo=�?i��X��JbF�R(�q�����s�ɶ`ŧ��\���v:�`guw�Q7�}4�����NIM�$��˫�Z~��:�i��W��zq�3ORo"���St��jW�H��9�H�e�܈���4���4�Cq�1]�K�3E\7�6�VC��qf�{����l��Aq��L0�j��;�ެp��R��R�J�P� 
��w.�{�i���(_�>��V۝�c/]�/}/2:��W�1���6�-���aٽ�1�pooe��b圞�*l���-�\���4[9$H����������������s=o����A�6�m��I#r$W/9}s�9����zs��=�㮋�zW��ȋq��m�$�G#�����O)2�16�%V�=���r��`�}Yo��xU����KmHKJD� ���z�l^�m���w W��� 6ªV�z��L�ʫz��9����x⸓�g���󏙇<E�³j�\�AN�="[�$HQ6ܒI$0�#�T��׽�3K#Oz���xp�B.�Pڦ1���:n����cM��JD�.�4�ټ�yHf��B�O+�X�/2�UoC�K
�C��fNug����Q�$���q�����Zed7	\�Wp��T���p�L��Xf��ݽ$�Ɔ��n6�o�ߛǳ�wR��~��]S�����T�<l]�?????���T`�WtSi]�
�uڽn�P�U� UaT*�����I��IC#�I"�����E����[۩p�k�O*��M��[ob39�T@%F䐖؎	�<#Nuh���Fi�M�Zed7�)�1Y�T��^�#ONlG���%MHܒA0���}��H�c4U�ySm�d&/��Sl�36'��6��f���PڊI!-"�4�-�:G.����Hһ�ͷ�x�ؤn=�\��@�çH��_a�##��$�����]�LZs�J�`��˱ͦ+㹬y�u���F�Ѩ��mqG�E�z6�k��Ej�����P
��U+ԪU�R�*�y�'7\�m���bH&]C�i�0�#��p\�dR)���G��q
G����4�4��.V5��7�I#��$#�a��<]V�H��1�#�}7N]C�i��YHf��+3�7���NFbm�����4^e\��C�\-9�M��ؾ]�m1X��;�Zf\7�\�;�[��Sg4�=�f�2�#H��a�FWj��FE"��m�y��x��A�2�RHLIIrL҈ӝ[t��L����<lV�H�̕j��̾p�LZ�ԥ��)����n�-�yEG��MU��N���yV�S���wb�m���6��p�5ݷB��Բ�[ku�
�۳���qb�˻2������.� �   �
���   �  �   @U ����`� w � m� 
� *�T U����%]Z����m��w]Q����m�nn�nZ�h ��
�P w � �^�$rF�m�e98C6�y��&&1y�r�އ��Zs�M��/b��k��a;���q6�m��E:�̸n���J��s�������!�v�\�dR)�����7IB�n,�]����&iDi÷Nv	��s�|�#ƛP�gj�1��}�T��l$�I��C�{2�Y�3�݄�s��ʹU��/=V�لi����w��n6�R(���p���L��^�R��Y�qn��bx5C)����{�4��F��IR:V��sRǮUUM����Q�*dW�6�q���6�j% Q�#H��;���M���?e[ L��/iU�g��uZ�!���J�$�F�m�dR5j���w�	����_
N���5O*��'ʮUo��.��2�b)�29$a�#�<#NuQ�͘4�#�����+!�^SR�³��n����25LoK@�B[l�"�4�|y՞��xC��/�>��&iDi�ۧ;��8FN�e����Ԋ7$B��������<,u¯t+�}u�I�v&�LLbt�%L����ֻ��˨m��{mz�PT;��z�J��T�*�ۙo��$�$����q{���sc��^ܽzwqk�����B�SZb�H�2F攊j�<޽稡�_W����xn�\U��.�z��^&]m8��$�Q�!�	����U����!e�L���a�����)�ޭ�'�4���d�oy�e��y���;��Y�h����sk�g��y����sd'"d�"rH�) `�>#��f�e�:F��S����E���ʛQP�.ۭ|�M��[�F�rH��Z*5����]T m�p{( ;�*�@���ڒ3��rF�nG�YF�3�L#�Ǉo�RͨR0v��p�:n\bz��S�]H�ނ�m�Km�#q�2�'���ʁ2�1y�����\,=���<#Nn-8)i�E����R(�m�X4ú�Hɡ��p��Ŝ�h�����b��辷R.�w^�#,��nI$�c�旈R:}˼�4�4��ӝ�`�p��iRͨR3���xi6����cM��J�\+4�Ǖ��^M�@�c���'��
G���Y��i�n��m�L+�Wf�+t���z� �b���Tm�PUY�֩��]��̥LMR���³�)��Ze��]5>���Sڋ�D�9�,�+8΋����V��J6�-�di���%;��4������*m�&h�����0�
Y�
G\$P�\i&��I$2D2�GL���a�����)�ޡ�ȈӇN��N1<w�R8Vm'c`��F�lG�f����&pR0�Ӹ5�Ze��]5>���Sڋ�D�37i��(�IȤ���4�i�V[u"��W!��f\.��ySl�3�h��
G<*���$���'��R���ϝ��� ؠ*�pg��m��n)ƻ�Sw�w�N�@���.��ܷ��*TVٳ��6�U����o;����ݚ�W��*�    6  @x  p   ��@le ��
�� m�*T m� 
�   �<V�nwhf�Tcwn]o^S�sM��.{� M�n��^׬����l�U*�
�U��t�;��L��4����w8�S�H���#�=��Q|)8݅��T	�1���v��%$��$������B���<�i�e��Ȓ�
�4v�ȴ����a��p�Ť����"I��r$Y\-4k��*8΋�u"��W!�i�!H��.�<����,�k���4��IH
G<6���P�gM�!���:e���C�����YHf��Y�l���D�J6����Y*�<������U��)��%��h�7�i�7Em�
&fr����z�7vի��wke�Ϟ��Uj�+�J�;�*�@�mw^�6�櫺�{�_p�|��E�f���i�������];��oj�l��e����q�S�sy�y���A[nt��/�B���S���В>Hۍ�#l����I��/&�L��^ed���sW�V�,��Ԗ�Vq�>�j�,��d�ےH�q`��#&�㦋e=��p�L�����+8΋]n����'��)8�n2T,�#�/��ySl�3Gʞҋ�a��P��j�gM�!���:n�j	%��rA�������c;=r *�ت�� UaTU+��:��n^P�&�4�Ǖ���7�&X�/2�Uxy,=�_�[0L��	��3�q�ڑ7!g)i���X4ú�+���8Xk)�E�4�\S�r�����I$o����OH����7-=���$$�h�)�E���h!
Y�Rx'B9$IF�&"O#�[�OU�S��r�,�3O{ɼ)2�1>U�����`�m����I(drHÂF3Oӆn�Fx�4�v�ȴ���S�,5����q�g�pj=	2`�8�	B�&6d�ȥf޻��λ� 6ø���R���U�m��$���$���2"�#<��sT1�*Ἡ�M�Og<��H���O�,�xf�u��nF�R(ܑ12F�h��y
هJ�U�b�OfvT_
N7ay7�e�b��jf&�TF�$�m�Sc)��p���1�xF�������;\�-17ET����v^�IH"27���h7&]C�3kU�1X��K�ԋ�3E\7�6�C�p�n�<���.�L�eD�$�q�	rE��p��i"��nq=�}�^�e�+�9��Ǯ�%6�1��~�n�J�v�ko[�w˶@�w W��@w [�Gv��ݻ���k��_����v���}��j�)ۦ�G���7p�w{��3YB'$�&ۍ���/��*�={lu.z������xn�\Wv���3"N6䍴܏V�|K�E�������nq/�C��{U�d�M��m�$qIW���3sw�^1��y�<���܉������Aq��j6�T�C���5���*ʯ<o^'R�WK��th�$�HҎF�B8�R(^jz����r���y�U/l��؍�Z���V��={��ᶻ�l��ø��{���<�PV���W��]ޞx���:�ʺ�y]�=�    U   ��   �  r�   w�*��*� �` U 6� 
�m� 
� @*�@��@U� x�*��黭��u�l�Ͷ]��k��� m�lUU� *���
������n�j�9#�o}�r=W�<�Ѷ^��<��A�eB��C[�`Q��i%Q
����Ȫ���2嶇�z{��Q�b叶|^ƣj(܍�$#��������n�m��{ɹ�=tE��t�u��Q��M������wٯ�Խ�p��-xVx��<G��t�B)���I$��x|GL��B<x{��YH�='n�E8i�z�� �t�{� hM��`�&����R�M��-<�PT;���U� U��:'u���Am�Ȫ�_.�B��3Ǝ�<�\.
[S�<,�Om��ݩ�S.����RI$AG��G�����OH�wy&���_<��H�^d�-xVx����N)$��L���iD�e<4��n!)��R8i��;�ᦑ��I(m�$nC����³����Ŕڲ���4�7���i"n�㦑�vq2�D�$�q��,�8E<7F�D4�,����4T���b�i��6�WWL[����8E^���2����齕�Ҡa�*��J��*����m����I'�8�R8i��$!K>#�NeC)�t�q	H�x��=x���OMxP:5��rH�I��2")�OH�N1<p����:�S�)øta��3�)��Z���+��
bfBf��#�h�سH�����4�4Һ�H�3�1���X�Zt�!	�00ӒnH˒<�ȧ��eӂ����ARψ���P�xi2�BR!<=Ϩ�"�$n%$��S�)4���܈�p�H�3�O#�a��:�S�)û�B���É��O`��c�w�ݝl�{R� �ت� [-��
���ڞ��޷n5]�R��E�(�`��>��S����ś�W���?;4��M�cRF�i%��OԎK��<Y=3�]�H�OO��
Y��<=����ҮW��S1��H�,&��G���,�p�<N�{z{{^��<^}��������������>|�K[H�6�m��pG���N�w��?ah}4���/bϰ� 8���a���Y��Y�F�aG���)�6ϸZz��M�"񧔼v��(��C���������`�5đ��fIJ���R�^� �<*��[��d��aIb�G$���l��C�xi2��y����翟����{^���;������������3Ge4�\�����#	��6��g�M�Z�G�)Íʻb����
���H�m��%�)���g�4��}Z�?<}��4�<zg������V[��i(�Q�I����W����W��y�a�x��>����<�^�bAF�$�M��e_�����ɿg�[�����O������y߿�κ�As��w1W���W��ueU1��^p���n ���F��7��K��7
����v�p=P� �Z�U�k�λ��S�w�n6�nV޻���  T� w    �  �  A�U �� *�`U  ;�� m� 
� *�T U��m8U�@x�[z��"�lݫ`�[\�V�[ �wJ�R��QR��7O���B��܊�w�E��U����G}ο]����&]eD�$�q��sgy��j��څ�Wۨo�ݻ������3��d�&fS&���9��˲W��{}ɻ7��*�A���$LH;.�܋{/����g/W�l�����nH�RF�m�i�<@�]w#�O�֧���5o��l�(��*��i���2j���u�S�7U�yUH��`l;�U]�PUj�
���ڎֽ�.�WuU$�G�:j��Dt����x�O�"�3�g�t�>8v���`�6ۍF�,�3�~�{h|4�z-�Y�Ӈ֬P���p����Ū6Yq��I!�I2��G˼�<@�]w#�O�֧���4wۨf� {�U�$��n4���ϙ<;�x��ws1���Oۡ�?t�o��1� 3�~'�R(܍��<G�N�3�~�����mȮw/����	6�`�H#fEK�*��om|�T U⪯E������[f# �1��n6�n%#�������p�������)����j|��#�B+�Z��I �H�i�{n��H���y�����ȴ�O��sZ}��;A66J��#I6#�F3�wa�Z&x¸o/�8V.mN�K�T[��p6�z�)&�nI!1E�x�R-����׆/G|��K���>=*z�&4
��!-��N5�A�`���
قQ��U�^4w�"����v�1��������B��� �G^�m�U��6���Z�@�w W��@wlYJ�v�K��J٦Q��<p����2��&�:F�N�3�|FwC���r���D�$�rIrE�G��ۣ��l������c�:G��ܻ����,�Z�)#q)$�8Cp���>��<F���2����c<D#����0>{�0���H�IF�&c#����s��}�3�g���R�3�����s)�2�%��Q���o��E�G�������:uB��G��1xZy�-�U^tJ���k���m�M��o��w
�����6Ք*���>6{�r���s%$�G#��1t~��,G"���􎑺njO��n��"��pQ�"�$m�ܑ�s ���v�1����n9Ӌ�z{�������}�����_^�����/>&�-��m�|�H�=�>����;˺'��{��߭�&7$mƒP���k�wS]��>�sjf7w��p��=,&&�N�6ˎ1ݝ���zs�n�`��w5��Eg���U����&��C�[wn�n�>8�,2  f���T�]{@ Zv@Pcwl6��ٶ� U�q��8@x x=�7���qy*��{��V;=e|���wX�8@x x8l���<�� <��������c ��V��@����	��8@x�S�������v0����#�{����lR���-�Gl*	�]X��n*�uT����k�� .` 8@ ���v�l�P�{h;�U{�U�Y7�x�A=z�;���UP     ��n=w  *����P
���ت5��d���  T�%UAT Z�Yno.�*�y��6U�o=��tr�=j�n�wv�{{+77nM���f�os��g@�8Cqݎ����m	�	��;��      �r    U             
�      EP        m�               T                  �  T           *�� Q�   �    �   ;��    �@        ��  P    �@    �@      pT      k��       <                        +��   
� �  @
��    �P      d     ��b�[�     UV�����
�d  �8J�k���ۥ`oj�l�dr��9�ݖ��xb���WH�< ���S�gmnw�c��לw ����$�Wm�� \�J��6m���Jm�Sr���t����K�|  *�     �   �  N U  � 6�VP �;�T  m���m� 
�  
� �Wt ��J�����sn�W����;a�V�G;J��My��T;��Ql�m��U]Vb���Q6�m��Nx<GH�n�|�H�=h}#��R]Ô�Ӈ��J~����Y�B�jI$�����8CӺ�:E#��w��G�;�N
D4�]Q��=#�{F�q-bI$IF�&"H��wq��Zi��_q���ˑi��?'�<p����i���)&drHÂF0zo�~_^ok�������z������ǵ�t;�e#�t����"-�rHKm�%U��4�T,�R��b�i��8�"F�`M|�oa�6�������ͷ���b 6ø���C�̂���.�����sj�I��r}n��9��~M�̧�x|N�9����n�z�K��D�m�����a�ѝc��F�<F�F���w�}O��OgͤdrG���!��=<6�ɧ�i�[#�H��u�t�GO��#���{�����nIM�d�
FG�������(ۚ�R)�]�c<D#��r����}W%�IĤ���ff2:xF|7�x�#|�^ͫ>��7�&p�&�/�4V.�ߛw�W�y�%;�f��ʪN��y`�ª�UATm��*��\��y�)���$JH�r�O�C܋4����wL��:\Ȱb�O�b�i���|�I$m�ܑ����G�<�аR��sj�W�{м&���|.>�n�_���J��vC$m�[m�$I�?S.<�܋�
��O&�<������U�?3����i��X8�n6䍖[�>g�C�YC�?^�r,�C�x��ՓO�ʬ����<C���Le�m�$�C�4�!H��.�<���}�
G"����y�w8�R)��k-7���&�wr���zEm�k��z�J���U^�b��VPUܬ��;�UK�F�q����<|w�������m�q���,]��kŸ\,=�_�Z���AJR7$��#�<�F���>g�C�WC�?^�r,�C�x��w&���^`&��6�m��g0�#�>��)օ#�ܻ��#����p�<.�'���x�!"��Ȓ�I$�	$C)���1��G���<~��]&��<#�b}2��8V_ZD�$�F�lG�`��7�^8N�w����tZ}�z\�C�x��'z�#������-֪�:ج��m ?�l�� �fe�R���qַZ��k'���w����?����^׏�Ͼ<�{�k������>=\��n�8<G�/n������i'j���h�o2�^>�n���V/e׈!�}ˌ��>�݁6�Q��7!�5��<F�Fk0��n���|F�w�!�+�􎟽\�TNIM�$�(�_!�<x`��H庴��/
|74�B���*m@����S1�����I Q�px��Tb�!�mfE�^>�n���V/eׄ�����~�}�kk["��i�pC�U؀�T8�N�T��@p���m����VW����;��Ue
�׀.v�퐸6*�2���k���w��;���Q�����Wu        `   <  �   l�PU�U �6�T  6���T �  @ *�U  UT*��� �Sw�����N���v�T��vn�`�ª��*�� U^�˦����m���z>��߾�X�W���Y�Ⱦ�V}&�6����F���>g�C�W�i�F�nF�He"����|�H���M?Sz�5�8G��5l�x�<��0~�ȁ�$&$��(�f`�u��Z���n�qZn��{��o8Hԓ9#n6䍰��K���ϲ��F�{��W�V��M�ګ\,4���$HQ6�m�h7|�|����<~�^�gj#ǧ.��~�U'�i0��]�@���#�F�EE�^���q� C����lY[j�
ɽ�J2HM�~�F��(X.f�q
GO�w�ϏW7����߷z�/������^w��}{_o�s�e"����1&�p7$�I�1��G���2x�㘇E��2<xFh��n!�8{�Fy���<ﵒgTm��jDی�a�l���}�8E�?����;P�=8.���<���")�cRI<�<a!��J�)>��G���
FG�����y�	ik�IQ��	R)�]�c;�0��d���b�����E���n!�8��w��k���:+;���m�^���5R����+(�
����xt%$McrH�H�aûsY�H�H�7q`�P�(~#�a�~ʳ��OJ�v$������d�"�"f�ם12����+�p�Z{9�M�<=ۡ`�p�=U��6��5"��
�a��tgR).���C~�ns'���C��w��#D��u�29$%��l$2�b�Q�<�aûsY�H�Hzwq`�P���!~��6T�H�7�&s����LTq�^t��
|s��B���]�x��n"oZ�A
)�|[Tv
�����l;�U]�PU` �
���ٽ{(6�J�����Ì=�.U&P�&+\�d_p��o%[p�L�ٖ��q�%���IXB��di���7G~��f�H��g��#L3���p�m0Rͨp�8q��	����q���8iVyO2���c)s�Sv�ם12���<w��B����$7�m���$r<��������
G<>���4��LV��B�,�i\�J��X���#�΃!�6�m7$�'2��u{�Q7ݹ0f	�����1i~q~�l�2�^^h�4�:zP��܁'��GP�$��ݞ�@7��� C��}���l�-��
�ٶ����[�e�T*��7���~�����O����ۅ�f��.0a�[�̼�F�t�=^�",���US2IU1m��&/��Sl�3v<���Û��I�p�&,\�d[,b��"ޓ!m&�%Bی<�C�i��;b����r��0f	�����1t�,��<#Nug���.5rH�-M)��c4���-2���d�<1�R��m���%{������9nB�0}�6�I�m����o��Rո���7n���q�S��|�5R�;�~�������V�#��^��©��{�Q�p��pw1�ꠜ��F��۽۲��m/r�^����j���P77�PV�YTx�E��;���Gwob�Wl��_9��    
��   � 8  *��*��@ U6��  w���l  U T*�T U��*�ᶀ�m��p�\z�uu���wvw�C�Ww��P ��
�fe�
�"�ʹ�u�6̀<����������ۅ��z�b����r��>�Nh���CO�3Ĵ��$�F�m�TUJ�`����Ʀ�>f���E�+#��g�1Q��9-�Z}��53?L��&�nH�2�D;��\�ɧ�i���+��gc۩��ƥぷ~��_�Q9$%��N%s����ql�=�r���}V۶�_*~ۛ��1�Q12TU7�7$A�w3v���r��û�����o���]\ĐJ$�C$q��79��U]��kՀ�w
��UQ�U*����m-O���ڨɻ���ܯt8N�{u�n{����cک���=�/di@�Ĥ�I�����Q�4�x��Bt�[�=��fSv��Ud0]eD�$�q��ɘ���шz������n���*����Ûm�+�
x"�d&j�H�ӭP���z��u	�on�m�{>Lw:o��|U
T��PTDUT�UR��j��Cx󛊔�onq�ǻ]����y���ϐ���u�|�Ϊ�Sn�� 
��UU�n�ڲ��l�˥w{k%J�_6?>�~~��ʟ������{���z�ҝ��󲩻}>�Oe�l��rI�-y����[�6o��Br�;�[n��G[(�������Q47x߻_�����=����3�\�L���1b�
�c��4�J'rI$��Y��H��Ve�b����r��0f	�����i>ތ���iέ�#RH�6�m���EUMZb��z�y�Y���<1��R��m��3J\�T�Cq�9n=[�k[zE�^���gw-�v*����� ��
�*l�pJ����r|\�jI$�(����(�D�sP�:n�eM�D���֢���W*�*��B� �Z�rIm��H�iåiLw*+�	��9^[�,��.T��"f�>Y
}�����2�J�""�����**�[0L����U�+��7�i���/
^����t�_8Z&x��lI6
��!-�Hr!�D;��\��be�W!�]����쩶H��W�st�F=7)ǭ���R)32R�V�W��s̅l��Jc�Q]И��.]�H�{йS�܉�3n��"��E5��QGQ�]��*��mª��*�� �
�wK^���(�$���I����]������-�&^�z�����֛ȴ��n���ӧH�6i�6S�F�6�?4�/�-4�qp����\e�S(f����p��v�eM�D���{:&)�$I6�m���ç��b3�LX��B�Xť1ܨ�t&&x�˗�C;��[7��e���%��ƃ��&X�����Bb��U�U���o^�Zb��z�y�Y�xNt��6ĒI%F�G4��0��n��4ҹ�¦+����&P�y���G�7}H�%(�%�"�CWRov=C� 6ǝ�k���N��;v4�z�)��{1v���Tq�Kwr�Y� �e  ��*��_+m"���z��w�jl_6�        `   <*� w   �Cl `+( m���  w  ��` �    
��*���Ԩ��m��㽅�|�],�z�ӽݞ���T��� VWqUW��[j�
��U5��<)�U��_���{�D�����8t��ՌA�b��������-)��E{�13Ö��ųRF�%�ܒD���3���(���#O`�̅>�y	�O=W�V�/a�{S��ON�l0��n6䍰�q`�Y���<1��WM��D��r����\e�S(f�;����I��M�#m�dk7T�G�����F��{��E�+�7*�*�LX��ȶY�:v��%��m��J\ae�:F�yr�F�}�?mș�0^fB�t<�ŧ����f	����J����U3��+�n����v��Tl;�+ԪU�
�S������P�6���c4�ݹ�˨����+5]n���OL�D�Cj鷤q$��M�M��o0�a��O�KT"���^�M�"�v<��V��e��\�L���|Bƒ�I$�	$C4��:f�r��&.4�˗lR7.R�.E�p�����4�3>�$�I$F&ÕR��./c��զ+�&�ͦ]G�+��i�a�w��p�xw7i��%MHܑ��f����ri�N���������ە7ċ���Zdp���x� �$��&8�Q�$�&ڕ�N��w�P��U@
�l E��t!�i��U��{�9�~���z׹�+e�ZSʊ���.]�H�t���ȧ�����e��G5B�a_8�1a\��U���vv:��ç��7x�g,�>��Pc`���$�nI Q�}yy�"�ye�^�a�-�{���{ղ�kQ!�&��I��#�N��4�T�F]����;��	��;2������S�*'$�&ۍ�L�F�<#�d)�E�LZy�J�`�{���LVi���,g�!i�:�i9>B2���-���I�=fހ*T;���.fՔ-�m�����s�Wu��;�ߜ���D�-s�SƸ��-0����e����㯚�?y���	�)$�Gi�{��/t,G��"�L���1b�y
�c��r��д�>9ut���6�nH�.9�C;�ޅʟ��L��/3!O�Bb��U�U���y���c4�X�QETL�[m��bC�Kź�H{��Ӥa�ɺ���/�\*b���}���F��|��5-�\9���4�;��b�25W�Qi�.n*U&U�t.���i>���e��a�� ���o�b��^�=�!Tm�pz�J���*��.;ͬ�� ������H���9HF�ޡ�/���xF�q�+�)>��0a�/~������n4����84�:A��/�t�z]"��Q�T:E=9ub�F��\��4Č27$��#�#L#�?t�W&/��Sj�dj�6��\�T�4�V�H|�N%�Iq��d�$C4�#���aOy"���)ڹ�<%�q�O�=N ��x�#��������29$p�#0�g�͇��H>�t����K�R!�w*9�H�����}�7��wm�����ʋe/j�Px���;�R��g��-��]�z�1�p�e�Y�����ݞ7����T -:���wd�3��*�5u�w���     P�   �  ;�   ��
��
� F�@ � U�g� 
� 6�@ C� @=V� f�w��;�t��ٶ�*�i�� 6øUW���6�l��m=i�����7�������3y?����e�����{��x�{t,G�º���f&�R7$r$���b����C4�#��V񅞨t�|ns�#j�P���E<#��Њ���HKm��He��!�i|��*Ջ���oj�1X�)�sk���<C�.�:F��|�)�#p����/�-4���LT7�/��̡�*�;+�1�>����6�7a�BoP*'$�&ۍ���f��t��Ռ@ʸn.w���1iLo)M�>g��ǹ����L�$�-��
8�,��r�ttR�^��w� T�m�����[-�e���6�M&i2�1�Kq��fc�o=��{�����N�ck;*�b��z�y4�-�<F��5��bI$�)��+<���#��LV7�/���C4U�vWtc����<��Sm��mFr<���ޯ	{�`�8t����Re\7	�;�V���7������Ҿ<���d�ۍ���!��6*~ۑ3`�̅>�y	�K���f	��޽�-1X�:�\�(����6�ŃL��C�=�t��0�*Ʀ���3��LV7�:剔3�����z��zE�[�Ʀƻ+ll� U�
�*�C� *���m�x��q��F�0n��#��}��&nǕ=pZb��sqr�y��872i�H����&�#mƒP�܁�?t�b��ͫ�C�_ug�xt��i�)�C�LZ_�_�[0L����:$&� nHҒ�4�:z}�t����C�K�X�+5]6�4��/�\*b���WO�=$�ۉ&�If�<"S�k�1�b����6�7c�v���fuci��P�+��,D��I$�
�U���7�����3�^\�b���B�O�r&`�����!1i~~��w{��W���[��YU[:y۬Y@6øUW�l�� P�ii�m�$�F�m�$�ӄiέ��\84�:t���L���h��,c������4����&r4�RI$p��#q���&P�xvS��	��k�T�,�=��#�O�]���qI$&ff"&��Ze\7������-)��)�p�L�ח.ؤn7йS�܉�3�%�v�qF�R(܄B�˫�CJ��;�+e���޽�-1X�=i��/�!�KӧHû9\1����"I��D�	˨p�>9ubHú�����3^��1�b����6�7a��_��W��-�ע���P���� �cmWt[6Ѷ��d��uTa�Ą�ȓI�$���ç��b*�LX��B�[�cwJy�?u�Kp�;d�`��qF�J6�{�1�7�Ӊ{�����Н:�~��n���c���=��GTB(�-ČGf΅��۽�˪Bt���6����}m�4#ީQ�&��"&f`*j����=�Cx󛊔湷��d'O%�����?s�BS3u35UU�*i�y��?m�Ǟe��;omyנl���f�ws{ ����NH�rF��ݷ�d  ���U 
���P��rY��nn�˄������l���v��Ӌ]zuC��L�ob�p}�8@z� �l0��    ����U	��osml=��1�p�� �p}� ���q�� �ǳ��8����=��7������v�� j��*��mW���l���s֋b�vs ؎ˮ�  U*�  �Y�� �P[��:�m��0x =;�G{�*�*�eT   �T��6z  T *��`dVPfASd�� �  ���T Tp3MWs uS˻�n�^ݹ7��q� {����u:�'��wF��緶���* ��7�z�u ���~� � �wݹ      Ve   �         P          �       Tp         � P �@                  �*�*�           w  @VM�T �   Um�   �   P     �         �   U    ʠ   �       
�      }� �e� *�   �      �          P    �   ���`  �U      � UT    
�6�  ��E��{(:�     W *��{�c��T��`<����}s�������;y�� x|�+=ULc�S�pw1��,Ȝ��77vݻ�k�����J�W���޶���*UT �6�������W�oo�{x��l�v�:�n� P    P�   < 
�x   k�m���Y@��� ��� 6�}�} � 
�P
�گAT
�Tw
��=K{v�iu��������nɶ�j�U�
�*�C� *����C�j��nIj.��d_��!�?O��4��0�=棜�h���v*b��~��u�(f�|�L%�#n2T,�suw�H��r<��f�yS֢ذf�\�L���5|Y���6��"NrI$�Ƥ�g8�3N��v�#q��ʟ�-3`�̅=�����~�l�3r/���̭���m�#�Git���9����2�+5Oc��Ɖ�_8�T�cq�N^}����$��0����=V8b����6�7cʻZ�b��sq`Ә�V�˼\�"�!2I!mD���K(�w
��J��l 6���r�w3y*UU������{�p�R��&x�˗lR7�\��b�0f��Sť�m��������j���UP��&^�z�h�+��6Rd�7/S�L���R��|�D��h�D���!-�H��D;��\��iC0U��O�1x��eU�D����i:x`wYo[�H�jF�D��Wǅ���+e�ZS�S|��yr�F�}�?lZf�Ey�T��)$���I��]]��:p]�!�p�7�޽�V�c4���L��q��?�4�4?.6�)l���(�MHeglo. 
��*��[*�mYAl�����p6JP�ܒF�?�9ut�=8.ة���\g[�����}��n���F��]Π�Tq��m��	��ذf�\�L���<�V���7����	�:������9�yl�B�I%��xCɋ�<#�x��[�ť���V�/a�cT[�Ҽ6R��n����
�i���$J����61Y�/�h��s��LV7�:�0���pͫ�����q��6ۉIU3*&j��"f�yWk�ذf�r�2��,\�![,bҘ�R�n0L�_�������^��ʥ�YEU��� �R�U]� UW��[ݾw��Il��q��s4�wW��}Ձ�3�B�t[�--yߡ[,L������#���]���q�$m�[84���E��S,b�T�p[q�f��.iwV�>]�K:p��`�#�a��j��*�n3a��k�T�$Lݏ*�p[Û��I�p�1b�"�c���69qD�h7 y��F��c�Ҥn=�\��b�0f	��>�yZZ�!�p�9՞�?l,���$�D����֛)2n9Ƌ��S,b�T�p[q�f��.1X�k�W�ffR���p����B�`��m����*��� yT3;�{��J�UDEZe�W��p���*m�&nǕv�Ń0���Re\s�.�� ���RI��"�8t���a�&n�!�ve˶)�z8)�b�0f	��>��ZGJ�<	i�9$�$�bI�8C/c�9�V�C0���L���E�~)�1Y�^8-��3J�jfbGAPA3UUU*iT+b����:�&P�h����v�eM�D���b��Es�|ӊIm���1�L�ux��8��1h��:U|���:����ǽ��u`�ç�-��l���Y.A��8C3ݧ�xn4�w�����V���S�c�w71���]�Qr�@�/Of��s���  ��*��;�2��nO,�{.��k׶ʷ�vy�T@    s   �  � *��l �\��w�*�;��m���B�  Tl�� �`g��Nz��*����)u�Vۺ�@2��t *V�UU�EQ����ٝ֨�i{V�JaF܅������87�yӄiΫ9tC�D#`��K�꺯j5���ca#�D�m�ؑ�v���г�緛����vS�=����d	��ݿ)���H�JI$��G)#�KLe�8b��2�8X67��یUԼ�3j���`�eD�$�q��Ɋ�,O���p���~�e���՜�9�B0�L�V����i�FAl��IFpCH����sut�"���,��c�I��)��O��8^-�Q3�{����J쳣l�ov�Ѐ`� �R�U]� US��Ow��`��D�m�����^{��#�a��p�2��,\�dZ���cyJo�aE�p��!bm�ے$�e!�W})�b�,O���p���~�e����˿L�!vyiI�f7���I6����n��^��"x˦f��\�T*b��;ю�&&`���'
��ۍF�,�sj�U#��}ɚQ{���/������Re\7X��B�G��"F�*�I!�9���4��R�'t{К��M�u}O�������?�߰�[n��UZ����y��m�@6ø�� �� ;��HM�#m��mH�s�fp1�)�sG��D>�b9��F��0ڻW7>�ؔR7$�H"�4�<!Ӹe�c����d	���[�(�
�wC�����('�$���m��R����)�q�b뺗|);�}	�~���i�6��Y��Ӟ�14�)$̎IH�N�:�.����񂗊��<��!�D����4�Y�k�rHKm�"�f����.n1H�|7�W��r�fiDi��7�,�w������U�W��z���������� �b���*��eQl��wSm��14���#�(�3��
�����y˫�"��g�^�&��4�0��
7�N)$��m!��:��۾Y�ӝW�~s�D9��)x�_y^�!��q�%��m�$���9����v��a����q�E8C�e�_t���3J#Ox�s������$�n7 rDs�"��X�����;�g�#��w�<�_R,�ΐ�z���|c��n%$m�!���ȶ �*����L����ϙ�4��/���;���mm]}�֪ݫ�o��'ymq� C��T��T�]�]�am8��$J����Ԇ}�o�m_R.��a����q�~�,>�^���O�x.�$F�RH�	�0)�/xe؎}����X����_`�������-_R5=����m�[m�$I���ћ	�ܥ����M�_��)o���be꼻�2!���k[m�ܑ�-����*<*7��A|��)�
�>���.1H�|�V�Q6�l6�rHa����W�>���҈��+Fo�Y�}�AL���D�
|Gߎ��6�l^���A3�+�Az�hqܝ��0���b��uW�ln������[ܻ{76�窀 �eP���3���i�{�󻼺����w�m@*� �   ` 
��  wU   W�*�����Q�   ` �Cl �ʾ� �R� �d7��z���W{��{[k�;�T׷{n[l.�oM{�� l;�U{( ;�*�@��|�[i�IFn@���߈�#��!�yw�h���a؃�VU���p�9՞�tB�J5rH�-O�|ȇ�M�
^+W�W�|D=�]������a����7�$�=M�m�X4�,S��^�{i��ul�3r;��R���}�AL�j��;�jD�JI$�0����p��������\�s�3�.����L"�|�\���P�$�F�m�$�l�ɾЊpQ�)�t������F��ڭc�F\($�7!aĢL�U#����T6�U]�TUj�
���R6�i��F$�RI$�����[=���}��=����o�2�#�a���_4�HKi��X4�-��(4����v���"������CD���O˭XM�\n)nCC9�_p��Y��3��ߜ��Rw�R�z���|`��}w����rH�m�܂I���4�v*}G��n�&&}�ǅ���Vi�Ox�^j6��F�RI$�!�_g���&U�pŉ�¤Ϭ|w:O.��Y��|����i���%$�a��S�o�g��
��YN�PT;�+ԪUWu 6����W{����UF�T�������|��{�]�[����|�x�}L���	#p�d�J3�����u�&.v�}G��n�&&}v�[��<k��q0��D�mƊrf����ћ�R8FZ���b�iLX���L���s�7�0L\���L܍�����g��˝CD�n#O�b����ik��-�2�)�PW
�go���"�m�[m�$E�0i\[��Y�1Q������4L\�T*��z3�ݺL~]�&�-�Q�S�H�1&�n�Svؽw�ۻd[h�e p+-�� B�-�q��e�����W���ﲭ�3r;�����Y��sI�p�1b�1A��;�ҌmĠnI$�c��8�1u]K����T۴�ϟT)��:G��4���Ћ���m��jD��R+6��i�q��zR��77K4��G�������ϵ527$�H**�����������U���ʷ�g��}��p�H��I�
F�Q��a5���wyS�R=6=�C>=#C���p�q�H�^.�\���2�
�EV�޷��t *�ت��*��l*�������Ӛ�ݶP���d�)�)�w�20���i�q��zR�£ک�V��Ʉl�B[l��C4�>=2����S�vE������U���ʞ�_����j���)(�nI!�F0i�OH��8��cySl�p�N��
O&n�S�'�uca���I���G�exv���q�6�LR+2����w���~w]>���(�n7!����P՝����ܬ[����{�M�N^�wy��wB��۰��s^��'\z7q���x��G�6��ll�m����뺶��m w�����@��P��;q^�ws<��ݺ����z�/�ݹ �    
� ;�   � ܪ �]��Q�� �� 
�� m��T m����
� m�`� p� y�UTn��]Z��E�z9X�J�N�N�e �]ҩ^�R�wU �
���k�n�کG���̿���V2�
�*qI����gԏM�r�Ϗz�7�Zq�ɒ6Kq�t�j��&X�W
|S�az;ql�3N�M1Yb�(<�Zf��a�ܔ"rH�IF�l���C�	�n��4��"H�����dR)���,�C�t�OF�0�m���6�MɚQp�����`�}��Re��>��\Rg�����yup��j��p�q�!1��$��C>=�'7s�#Nt��j���w5f�#OL�~SO�
婕��Yn;���u��ls�l���km�l;�+�@� j��m��j�5M�a�X4�ڼ~�{>!�tM�3ut�=`�&����Y��>8Eﲒ�L�a�ےH�qg���۽ɔ�)��{��;j� ����h���ߟ�;��IB�q��\?I�r�ύ�MV7.(]���T�Ӌe�������\j�6�S�~WO�c���W���`��3��n������0����Q)jg���m�"���S�kM�_���۫�������t9Vz۬�Jiq�|�nF�m��MCsEY�۪�*�1UWt �6¨*��Z�дAA��JI# ��];�}��5�^�:4Nn�E�P~3W�W����$�F�m�$�f�"��e���¸��Lú<}�����MҶ�O�I�KL��(�JI$�8"�a��Vz�O���-�����{�)DS�i�؎x�!����惊I!-��qF0S����MU�g��1���ta��S�|)<f��sw>�6���m(�n)nCp����/:ql�q�w1E3�da����Ϫ������}F�S|-�Q�zލ�Y�[��:�Lt�(P�*��U*��(PUn�w���ڪ6�rA�WO���Bi|y��^9���;E�Y�8�@��re(�p�7���H�JI$�r�?w�tANU?bj�<,9��M�F/M9w�l{������D�m���3�L#���8�-t��b�J�1E3�db<�Zg����$p�h%���>!����_8����S�3����x�o.�Y�8�@��4�F�I�䌹&R���M�<~�肜>���h̃O��wyz���XQ)�Zm�2"�A��u�=m���ݷ��l;�+�@�V� m��^�n�T�U䣙HgǽZL��|)�z�A��/'N�Y��S�.��i�a�դ�E��m�$0�������{�!��ڳ`˫���=�O\W����K�#�����n/<���ܔ��y����zۃFf�.٥��q(ܒI$0�#��|����ⱻ���oV�ս�j��b�m�x�n6�R6��4��O�c����x����<St��i�8qLVx�����W:�i��{��=b�0��ݧvW�6:��xw�*���㝰�;p��c�:n��eP8t-�wgp�d�Ku�����m���{t��k�w9��ͭ��p�      �     �   �m�q� 6��UPuPP�  *���� ��C� �P�����N�=�Mː|�QYV�r�V��o\��m����Q�ATwZ���*�^տ^��_�~?ȿ��/7�V�x�Z�u�_?�T�����('�9#q(�d�ϼF�w��|�~�����&r�2;�P}2��'_�,�AI(drH�2E��m�4���qi�{Г�������P��F�D䐖�&ER0�݋}���v�E�Y-}���C�\�9����oTn4���$�
a��h�}�0��ב缇�n����M�>$w�Gɽm���e�̑6���u���@P�*�©T;��m��Ԇ6N)$���I��t�/�����b�b����qi�{Г������%�bm�$��D1�3j�f�Vi��t��_/{��VG�[�V�x�ޕ2���D�m��.H�}���x��PQ$��a�缇�N����/K��rD��7�6���sơ�Y+=���mH�n���%�d'IbH�H�$���t�z4MٗP��R����Y��}��Y��_��M���ʶ�j��빳f�Ҫ 6ø��������v���]ӑ�r`$x���>�Gv�<a�V��n�t�>��G�ˇ�]Ǡ�n9$&6ܒD��B>9�4Nn�����鸇O�vʰB<x}���4����Z�m��m��nG�K>���f�}��F�՞������)|y��^H~�_y��e���$�H�qg�1��ܘ	1�����7z����������ｷ���ם��=���L%D���-��ï���O��>ds��>�x@|>�X0���[��ߩ��x�2�n+�s{f���@U�U^�Q�AUfwV���2cP7$�&�#4��A�������뻵�����0�ki��,�{ ��m��mH�kЍ�n���n�'��^_}��}��׵��}�y�=?_�����x��RI$�0�}�0�;��:p�:�\�����9`�Ο �a� �t�q�$i&ÆH�a<7w~�GǇ۱���4����ƤI�+n��˧ͪ�"&&D�JI$�8$c4�>˒:p�WvE���^o.��ŏ�����*=>;w�v���������IwLu�u�PT;���*�� *�gt��������f ��NU��� ��0�7�6�0�zi˾�3a5X����m3u��Q(�R(�b5��!��٪�b�N�Ԕ��������;�xQ���ʾ�$��Q9$I6�m��9Ɵ/u��������x�o.��@��re(�p��/[R)�I$�C�@�x���)�j������a�o*m����.�Rx͏u�J%�9$I6�o3��CL"�P~;���v��3O���O���>��,�Ҟ�}ֱ�@�����|�9��ܲH�!��IЪ�"C+X�FjH�%�!|�""��iO�$H��*�5����g�o��c���=4���ky|��ٔ�����n���r$t�! �v���O7Y�{�z����ӧ�wSw����el��V޽�D�$J$D�BB%�$)�qQ+��y)�f�$��6��Ӟ�2z����! ����<��t�:���_�l�	�q��Zݚ�8�Q$�t��u)m�$;Z5_$)�>չ��|�{?a�[��SH�pV���� BA�ۜ�k4�[oɝ8��Z@���ٯ�@���oUnъ���[z���Y�K�џ}3ݔ�	Y�iңn�w�ݷs^��tH�qg�k��)W�ѷ�O]�o��d�Mf.124��~�A@����@��}����                        ��           P       (                        \�        h  �&�bj�6�e�V��cV0�X�U15T� T��]jq�^�]�T�-rݢ�S� �U�ה�8�J��ڔ
cR� ��R�A�)c4�)��)u�4�+�          :R���R��N��������� j�ZP�T��V6�UX wmiW-J�Ynڔ�6�J�f�U` Ԫ�ڕCR�VZ�J�ʪ�  �%Ys���R�VYU]�T��          j�U��V6UUcj�LmJ�` �E15J�U]8�T���UX 5R�T����U��Rcj�` ��q�R��u�+����m(� dX�*�j��&���T�         t wU*��UKUU1�USUT� UUYj�XڥUc5]5rԪV  ڕS-UKUJ�©V6�v�� �U1�R��j��f�T��R� ҩ��U1�*����V3J�  : �      u*��j�V6�J�Ԫ�6�ڪ�5UX�UF6�Ue�Qc�� 
F�����5*��U+U*` T��l���WZU�U*��UV  ڪ��UUcj�V-Jcj�� �~A6U*�`L�  !?�$�*�S�2 4��B�F��#&#F� T�ڪ�#iT�р  �����UJi�h�a J�2�%?A4@Q�6S�'Oo��~c�~��z��߾}������}�w~"����*��?QTA@�""
��"
_�_�����rD��O�M R}��q&��q��s�ےx�9��3��&��8���C��!�u� �B�@��2�ЧI@*�-`]*�� 4hD�"�q �� 2&� $U��Qx��Т	��E���t
�@�Q9�9�8�T�4.����J*����: x� �:`PCN�  q @ ��@�dN$y�
��Ƞ<lЈ<H+��(0��H��8��Ec�Et(����.�}�>^�l[[���4h���+j�*�AMDS5URI�Q[��(�U3#BP�@R�P�j(J'm&�����(J�"&���a��"�ֶ�SMSL�2�M"P�%	H�%
P�%	H��R��P�%��H�%"P�%)BP�%"PBR��BP��T+JP��N�	T4 �ҳ4�H�"�@�	@	BP��	HBP�SH�%	H�%	@�	BP��Д% 
R% DД%� P�
P	E"P�IH�-����Д% �)Bb5�M:t�R&�@��*���R��4b*�mkLF�16�����"��jJd��� ������H��f ��(�*�(���AE�-mEE54$�--E%4DUlb��%&��墢)i)	� ����*��*(���#[X�[gM;i������������"����*b�#m1E-R��.э%`�AT�PPS��$���
��P�4�SD�Ƣb�b(�CA��h#��LRLM�S@ES1%V3��E�U:*�,Fh����&���j"���h��$���
��5���������gSE-�4;cV4�U��EScbf�g�[DLDV��:4V�֋j5�m���@�4��%."%"ր�t:GN�Q� рЛH����2�P � �P�$BP�%	BP�%	BP�	BhJBhM	BP��%	BP�BP�%	�%	BP�%	BP�$BP�%	BP�%	BP�	BP�%	BP�%	BD%	BP�%	BP�%	�%	BP�BP�BD%�BP�%	BP�%	���(M	�(J��"��(J��Ѡ5�5�"tѡ4&��)���&�N��-�N�	C��V�hJĺ�M:���(�6͝	BP�%	�%	BP�%	BP�$BP�%	BP�BP�&�J��(JCl%	BP�	BP�hm��(M$N�ք�4�.��(J��ӡ"��(J��(J��J��4�J��B�b�(t�R�Z��!��%��t�E`��Д%	BP���%	BP���4%��BhM	�(M	�4&�J�КBP�BP�	�4��4&�Д%]��&��4&�К�И��Q�BR��4%	BhJN���!4ihJD�-��6�P�&�Е�4%8����$6�N�К&��PhKb$��К�К�����&�К��E��1%T�D�E���(JGKH�P�JJ��4Ŷ�X�"+m������˭#���Д�1��KV�[!�ѭ%[Dh��h	*��,j(�6�HZ,�ƬŶ�cN�ITZ�Lb�46�m���Hh�mA[E���MAI�6�Qf(���b�ŉ�N�4h����kIM��F����)(��hJV��
��4�i�
)�І�)�BP�$BP�%	BP�%	BP�	BP�U���"��(J��(M	�"BhJ�К
��P�a4&��%	�(JBD&��(v�p�&��S�	�(JBhKa)IA�(J��4%	�J�,I2��)��Mb�`6ɝa5Aki+��j�!(J���)!4&��%	�)��M	�(JBhJ��D`�E��%"R%	BL���4%	HHl��(J��(J!(J��(J��(H�C�(J��(J��"��(J��(J��JBh�AD�(J!(JM��(J��(H�A�(��J��(���F���Ѡ�cM66����mZ�E����mQKR�Ŧ�րѥ��Кht&�]	B[	BPL�H�BhM	��4�Hb�iM!�4%	�"��(JJQC���(��	�(JM�.����4J�	BPi4%	�(M�D:]d�К)hJ��4%	BD&�ւ6�hJBb�Д%	BhJ�И����	�4%	�(J!(Jt:BhJ4&�Лa(JBj�КD�4���&��4%	�(J@���P�%	�4%	�)M	BP�&��(M	�-�КbM	�)��(J��	BP�%	�4%	�(H��4&��(J�
j+j�"��H.��*�D
Dŧ@�X�hA�V��)Ѷ��.��C@�B1Z#�-WT�!H�(�%#�)Ih�	��b֊&f�m�M1���Q�-*ҍ!�T%�j�jZ(A�KE8��u�����b�:�F�Z5@�9�gkcF�`��49��m�Z,ؘ���TE�� �)����DUBU:�-UEU1D�3����DD�BE�k#�iH��h���S�� �j
�5�h���dĥP�ecg�E�i�
V!4��H��Q�4��B������kIZt3-SI��4!�4EU�1�ES�F��h���(-�IV1����IF���+k�E:�hƍ�t�Q i�H��LUDM�ŋ1T;P��5���5�5f��D�Ƙ�j�Nm�+glFpSV�&'cit��$�""�4ƈڋ[gNH�I���t(�	��ӡЖ53���b���CBh���Jq���4U��h�&��hh4�fa6h1�)"*��0Sl%�����E;�т��&J����"�����F��&���"�i�S��Nb�FI�_�^_�����&Ad�$�����_F)v�|+����U����u�5�Zx߂Ƹ^wu��n������,��W�V�O�4�G����A�TBN%{��{[;c��   aN�^�aRʪ     <  n%���;w��ҫ� �'      N    �    �  N ��  �8    1�p���p �   '     ����    �  N �   �'     �T�8@ � aTU ��� ���VĆU8@�*z�'
�` <U< ����� 0 ���   � �     p �?~@x x8    `�    x    �x��     8    ����1�   N  8@x  '    =��1�      �     �Uc �*� <���uAª�*����    ����� 0��⨜i� ����\� *���@�� �T �A�d=��6��{wwmwgvӄ�lٲ��J�*��u��[��s{��:ݨ�{�e*�:��5�p�+tP�U�{��@�;{!�/f�{>�<����q^�U�х�-ݍ�!�����ͱ�7�t@��P�]��zֺ���&���y��z�����S-l*wN]�Vz�����9r{m-�eE��ޣnm����g���q�ʙ��r���y�b���ݙYewk)z�1�݈    P  n b��Koj�� 
��Wf���� l�^�V��w��1t�W���1����[� I�*����	ù���*�Z�`!�  /��U���Y�� mض� )��Z�5������GwWn���v��*��硶.��+]TU-���y��J��g]����xα�k��Y�w��A����&�WLkqSױ��}��vޯ-J�\����8@ �	��������1�p�^ 3�3�W�m����]5� ��R�/l�z�'Z`*��< �w �p2���K&��(�V�TU���;�녥]�9L�m� c ���p0���ko=z<�Y�խon{F=�V��k˺�z����[��l���vy�j�S�J����)���Q�u��m;ỻ�7u�[eeof�T�{����6�ݻ�Z�u�ol�Y��fѱ9Tཌྷ���n���m7����;w�T��Km��Z�M�Yz�P�   ���j���^�s��ڗ7k�5�or�kغ{d������6��
�x�
�ʠ �wVy��  ��VҀ V�Y��eTR�M��;�)[[�V� [-�k��T����Q[����Q^����
�������Y�ݺ�n����[[=R݅ݴ�۸ o;�y��lz�[[�v�T3t`qVT��-�.j���T�=�}{����+�x[�ˬ�^�goV���]Jf��2���m����fԮ�mwoL����޳�[PΜ*�Wv��[*�T.[&g.�R�]e[j�ŵ���ݬ��@*�;���=�˴۷b�ww��;�� lQ�6���U�lڜ%U�gi��@���Wsf���iWw+kmw6�f�%�j�b��9&���op̮��ܪ��w���*�r�-v�tҶ�swo�ڲ�wj�m�ί�����w��_w�'nk��2o=��U�[�VѴ�k���gvWm��w�oo7��N���7�UV�ղn��j�V�n\oE�v����sΥ��1vh��ܽmE��{I�w@T���t[ �l�z��@WRݸ3-;j�AY����u�׼�m�維�c�kn�Ge[^�Wn�9f��ۮ��}�޻�R�6�Ż�ؑ�^p6(*�2]�ݽ���u5��{�ǻ���N����Vn���3*�=��l�X�W��o��8��
�m��nn�]��i}�ڪ��kw*sm�U箸�z�Ư2�˯s���<xٹu���{w^�N�U斮[7���g�Օ�w^c+\^�y���n�{m�����7Z���sݳ�g窶�եA�l��w`�*�n����5�=�����2�ZY���Nm�ݻ�x:�pZ�z{�ͽ�m��E7M��zݺ����Sm�m]g�պ&��P�u �(�t�Ев��=��{e�ݫs�J���8&�JU�]նr����sLm@  �Nw�hǺ�ǭ�����6�z;�k;����9ӹ{�n޽׷rW]����                                                  �~                                                                             �?                   �                              �
�U *     T� �B�*��  �X�m�A��   U cl  \�                                      �    ��   �*�   m�*�� *�      P                  �  @  � m��    
�w�� �          
�                                     �  ~�   �             +    �       *� TT  p �        U  6�l�<@N �R�  P�?
� ��        
� U    ���P@ @ 
� @ R��i�ݭ��-��
� � -�@R���|6�w*�-�:vu�59�                    x�                               �               T�         *�@     A�     ;��     ����*� *���  <[       �p   x      �                 �l��  x  c   �߀     �                       6�                           
ʪ 8       �W��        
� �     P�m������h�e@U U ��~ P     �M��     
��U�               ^��6 P    EP -� �T  
�    P�T*��     �?     �U                  6��           
�    *�        �   �  �           �          �              �   U                          Pp��              Pm�  �   *�          �z                r� �      ��� VW��U  �~                     m��U
� � UU� �   �J�  �S�]�     P.�   U   
���Tl���,�e     �e���BuP���m<wxW�G]ܖ��.� �T 
�U  ���@@6�W^���N)���� U[ *�slM�J� U �  U     �m�mTPm��N�y��ƭ�]��wwog�=T��J�  ��caݺ�p��Z���j���Um�+�� �JH�n;�ԴD9M1��j�g� U>�A���z�r��?A@����Q<{�y��u|��?{�������`� #�o;z< �  p��  N �P <xTU@ N  8@ ND�` �� 0 ��   U��W�� Ur�   m��SkIS��W��ovڭ�R�6�^km���A��f�sw��̖��� � ����Q8��=�6ʕUl����^�����˻�m�YE��TN �m�*��J�� �
{�� <wn�+]�w\��{���my��s�T6�fչwbQ�m '{��s��t�Pb���K�-��U���B��2Ͳj���w{�T[{E�R�k�=�e����2ʨ�k�ȝUsmG��}����i�u޵�oq�����;t���m����ղwV�i3w<w��su�[�s�t�i����uv;�9�w��mn�*��׺���Wq��;��Y��Ϸ���ս�����<         T              T            *���6�*��       � �  U     U��P          �   �   p P�U  *�6�P ؠ �w����        w   �    ���� 8     @ @*�         � U   ws�Ъ -�P   �T      T       @P              �  
�  �  �  
�@   UP *�� � B�@ U�W� �AU]�ڀ��  jڥ�� i����מm�[�����+�I%���$�HI$ �$t�qT 8@ g�Rݺ���0sL�f�nzm�0�U<�����K(mN�׫�v�V��ݲ���Ӻ�A;�v��ݻ�Ʌ�붭3i� U  P �� 
� w  �;�*��w'�*��[*� S` Q��� �  *� U ��6��Om��odn��~*H���� 6:t��i��b�0@ @$ �L  � � ���"��co"6G��H��-L��I�2C3�͸{G�f�R�"m�$m�A�dyg�3)�k׆�1�K�0�s}�X�ح��yΝm� F�
i8M��s(�η/�y�g�'���Py��S[����Q_U7 @�F�����=�o}����k����^�l����ɘn7N��� pa!�i�S�[��>�є��^�m�����m�;y�=?d͒I$�H6��viR����t�Έ��Uk� *��TU+�YW��[�y:���Q�g��p�}��++r��m�Y��Y�,������N���r 1���g7/����]�<{���h���~�l���d�]	:E2  B@ɻ�^��6�{�ܺ����YO�5��g��˥��꒯T@ M���{/w҅��ۋ~�l>�����yx��Y��O5��~m�7$�H�V�}��m9�w��l��lߖ�ݽǿF��/7g�J�I$� ol�z��دm�n�O]� U�P� *�m�ծ�{z���U���=�f�fLϦm�^o�o���,�J���1;�8Icc�$�)+���X������m�|_�뮚}D��ׯl��_���Im�����zZ��y6W;�~�޽��WkO�tR�S*F�$�2J�ykoMu�׻��3>��{�e=������$���H� �R)�V��[��n�{z����׻�z�ſ\6���I$��n�L���U��m�㹽���� a�^� �� �wn���}ʛ
��z���]�Z燱������M�~�����7ᔚ�$��4����{�}�v�;A�4ۺ���_<�n��E� $L#��<��="��|�=��w�z����^��g���֑"E$�5 J$6��*�ܼ��un�jf�u��_-�z���z� ��0�>����׷����>+בf�Yw�wc�0��$�I$m�$�B����wj��={�� ��U@
�pUQm�e ���g�� �C{��\���x����e�c�2��V�7{~i6��A����{qo�{�Vn<�j�V��醺��>�#����(  ��כ��o����/^]��6���Ȳf�Yw��4)'i  q�<���\�|���/v�����/�v�^kߤCcrI*E,��m�����ܺw\�Q9O���l���Gn��,����� p0P�nvjj{���a�n�Ӎ꼶���e&����wz��l�[{]�N����n�U�V�d���h�j&T�J�`e����s�`       �;�   � �U���
��;�UU ]X�   W�   �*�P A�?
��xn��[a}V�w���uov�o�l�z�v��Ymy@T;���U@�T��*�u��i%�#nJ�t���sי��y��.ƻ;u{�z��_�N��+J�RlnI$��e�{��T͸c�}��;�>X'�J�ُ7ҁSr�$�67G+�۶��������[��tu�W�//�o=)�@��-�����y��l�v߭�]y���^�ׯ���?��A�I#lH6B����;A�4ۺ����M7��g�v�����]m��ZUo;ײTy�ۭh m�p{( ;�*Tswm�7�PD��I�2J{�o�[�ͷx���������y���߮f�`:�I`D4�S/-l�Z�mL��l�>�k���{v��;�9K��8A )�=����J��Z����k��+&}W��k�~y��J�?TA$��:L���Ҹ'�z�Ay�U�R��{7}9���N��  @B	���NP}���e���:����Λw���UNU�������u�w��O*� 6��*�t �wPUW[�[w�(	 H��h��������J����lu�z��̛��);` Tܐ׻�Q����y`����m��:�#�ۏk7o����L���%]]֡}���];���r���:^6un����m��L�M��J @�m��{��^��]��֞=��?Xھ�}��;�h�o���� I!��f�57u}^�����׍cT<�gus��pU��Ϸ�<���f�n�� C���̪ � *�ηs�v�U  hc߽����C�g��p�kה����[7V��O5�6�6��$�V��w�a�:n����K���Zx�S��.}��MR�A$� ����wU���|�����.�{����z�����"Cc�$�u�F��k���xcz�/��~˧t�}�(Po:�z���!$�  �[�mL�-��>�l7f�Ű`��׷��Q���I$�^��ȫ��o;������0 ��{( ;�*l�8���2����fI &��K�S3a[w�w`d�ܫ���a��c�=�<�i�DI"P*�sǅ�T}ֳ�5�����ܾ���p��֌xQ�� ��	�
�y��e���:���軮v�qwK�K�}��@�I$�d{{�=V�n��,�h;e�u^�{���v���) n���P�(a!���5���{koB�#_n����&�����Ğ6�I$�I u`  �� c
qU�V�����}�m�l��w+�Z9�G������r�Bxt�l�����N�ҫ=)�wJ]μrw{����ګ���U���yT       U<   
�  � �<��pm�lP N� *���:UM�m� 
� P ?꠪[u���*�/Wv��@ .�Z<���Nɵ�:�f�������Uw��cU;���A[�����/tt"P�$:r紡]���wun�L��l��k4͏v��֒�c�T�Ϭ�m{�x��hS~�m�!�/����}37�~T�H���#uM_o�F����b��x��t��ߛk7u�H&�� 80��}��߮6�<P������mf�v����b��QIA$�IZ��x����/#����ǥ�B�����ާ�l�$�D���
pGy�{Ou��2��w]�*��T;���BjS�0I�8O��Mۛ~�~ˮ^����?k��:F����zܒI#C��n�*ߕ��=~���Z�VX���'��(�F�T)Z�F���#��*�y=�d�Uf�W��j>$H�2~�oL4��Kbh�U��A����crI$	%^���CwTG���õ��z��ײ����ߥ]j�-V���
p	$HIEUPC��#�m���#x���t���3�u��,��3Yb�����߮���ov8]ǣ��G+t�^�.a�^� �
� \��v����r8������3Ku��,��6nʘ��+�&��x�5ޯ-U�ž)�cL	"PIIGE��_+Os�
�UkR!��#�Ϗ�����C#ǋܺ�#�巶l�����I#$��UkNӪ<l�<Cfؾ,��I��I �)���;�����o>����������%��b��4�}Sxr��67�x��I`#�9*+KD���{ݘrʜ0	7�70_�G��L9W�}�C�fR�"�#�V�u��Dn�%��yr�~|�����<�CfJFI�W�w�.^����	����U���۶�^կn� m�pݺ�UATm���Kn��DL�F�"$�<���һ����t��Q8�(����d�D"?<�au��U�~���H H:	y�!FT�m�ϸ�#�&B"D5S��<�*�W��4���~��f�0~`H@�)JK�U����7�U����m
�$C�i	�K�~e�UX�@y�⍐ 7I�.�5[�V/߿w���� '�<@�ǳw�'�{��G���|\��WĎ��}p�=w�y�]_�
��h��萜p	$l����<y��x(�S�*��V8�?72`e59�B����ڶ��I$� �%2��[�e��v�w�� �wV��l��
���:܄@ @���Z��2��aGڥ�D3���Я��~���ԯ���]�xQ�+ܞ`8������ĩ! ]~����ֿj�ԥg=��
�#�z��W�{��<#�Q�+�G���q��d�/�^�}B�=��r��1�G�_>�=y�8=[�7 @ b���/�������ߍ���W�!x��+�G�˿~w�%z�нq��w�ǁ}����(�w�
�#�z��Z���;��*?6��� B��~���>�|��λ�}���+ԏP��w�Q�!�<H�׬��z�ߎ%z��(����8G�^�����#㾻��Ѹ��D�H��~�ֿ~���~j�~ݚ�>�y��(�9��W��X_r��߯<��r��_2=�ѻ���^�������}�w�����׻����C� 	�    P<���ww��m��V�V߷YP�mmOn����x��@����{o���s��Z�f��|��K�q������չ�n�����       
��     � P�z�*���  m�� z�  aT U    *W����x ���R����u�y1�Nyۭ�nҼ�wYݮ��޺l�m���� �R���]U׸+ʭ���=#ԯ������y���G�Q�W�{�x���^<a}�����ߝ�G�^�t/\uѻ�����|���7{�
�U�( S'-ܷ}ǝnkG�{�7l}g�k�J{�-%�wE)I F!���{Ϸ:Z�07���nɫws�}�f_�J�!$� �Q���7<��Qr7�t�N_Sr����˲�j]�
�Ȥ��I"d�J���Sm6�f�Z�cG�{�7l}g�}��������yݽ��{����kw�]�@l;�Uz���� �*��oc��I#lH"N7��Q�ݕ�����!�[yUc���<-����@�I_&�s�RA �B^6�����jw��`����K4yKYS�os�%���Z�n�Ix��xO���ɋ�R)$�@J�#��Q��+/�g�$�]���۳VT���7�6�z�yO�v7���W[���ǥ:��#!-chlm`�z���5~P>S��*�N���T�`����s%�Z��{�l@���U  #t����֦�	�}�5~P<��=[?Tf!𚸲�4yKYS�ws�%�^P-�����@+ng}�<��zmm;r�y�����W�� �+&b�[�m�� @����6�4�5�{˳�{ �5ee���Xh��P��祥4C���P#�|��̲}28���HQ��-M+Mkx����Y�%eL�^�Q����w�U��{:{�0�5e{yH*@��+KV�6�ʾ�OykcM���SW��|����Q�p��Z�|�-m[ckSY3ZI��j����g_�P�ީ/�	��A����Օ�v'�(��P��5eOX��S1�#3S0 7!+��X����x�Z�V�����o}Uf)+*`�W��L5~P>S��*�y�<&/~VoUUUUUU$��+���8�z��� 6ø�J�pJ���ݶ�Yn���	"B�䕶����`�X��>m%�n�f���xN{쩫��>^�O���.M/�Z�>��)�"�� ����Z�l�-eL�oXY�<�(|�{�R^)b'��{�0
STly��QZX��x����}?8�E$���j���9iM�&���/�l���f��WV���l�L����z���0��@����,�4K3UT���U@S)�&,߷���3&MZSv�J	k����9��)�A�9ﲦ�Tl��잨J�Z��I$h����ɥ�ַ��8N/lɋJh����f�(c�T�n�I)b'˺w����dե���ꪡ8�uڪ�q��[�t��V@�w
��UT� �
���Ww{$m�6�(�������|�Z�|�}�t�~�.�a+ZŊb�㯵�U�N/�f����6��;�/�|���*�dq�t}��Ϭ��;���>?m���/*�_-���	$�"$������.��F�8v�'T,��8��ۘ�~�3`�TU��o���%I �9�;�k�i��6TU��/�f�L�#
oj�~ㅷ�V8�<x���g΂D �$��"�V�W�|g��-?al��28�W�v�ix��˪#����y��n���   �  N ��Uyխ�x��o]�ܤ��{����k����1���e���6^��<�ӫ7S��n��-���띹�=ӽn�ۻ��/sݻŶ        �  �@  �@ �n��*��VG l   ��  T  U T 
�P['�U[�<�w[�o�K� nro���y޳d<�m{ �wJ�����s�p���Ȋ��P?8�  ��?�^U��0�˯�����eM�����Q:���Z���nb�����h�e	��$������QƩ����T�*j�˻�Y�b���٫�h���t�J�����ng6���P 2�=�D�5|��VSf�+�|'�~�0��@�;�b�T�5LY�lO9�bַ�}��t�h��$�! +\ڶ����0��M�t=�3z�j����~��4LSW^�f�R�T���~�I� �?yk6���V�T��X�����}S����.�OTQf�����f�)�b��Y�8
����m�y������` ��
��@T�.[w]J�����-SS2�UL7����Gdݚ%���{Vj����{o��W��1��S��1o����1SUUU�T�UU1����2Q�%��W��0��M�t=�3z�j����}+�Z��k[�e�#J*A��TT�L٪R�	��vyy@�B�z���,MS��w{�0SW]�:TV������o|QKΈ9$� 	�fs_����+~�m/�)��Gdݚ%���{�M��.��������Iy���|P�$��T��)�j�����c0SW�7nd��Z�@����A��'��ʚ�m%����YZ��%I%F ��&�ӛ�g�s���� ;��UTب�Tm�B����ݎz�@�P���_뿝����O34j���'g8ݞ^P>P�ީ/T�5O�����1M_6w>*�"�nI$���*+Z�,��=�f�)jz���/�S����쀥<�]�{*��%uH��j��$��I��������1��R�Z���ٌ�1ؗW�w\��.�^�9��� >P��:@H���������nN�|Fajyme�&h�Rl������
�uIz�����|$�1.7$�r�!�$��7�ǜ����-uC������3	�vwD�_(�˽���jy|��]UUUUUCm8�sM�q���y�w- C���w�s��b�.�w�5�R�i ���ST����Y����1��R�Z���H����m�Q���7I-Ͷ k����� ��<�) |'C��ި�,�y��3����OC�f�+�@u���o��6���t�$ ㈑���i h�/����0	Sˋ/�����T{���@'_t�򁭯���4�$|�	� ��=�I+����Յ��.����0���b��1U�@�����N�f�c7��� �@q��V�&�z� ۙ+8��P�S?3�y�6�<�Zk�B�W�o,�BI%F�u�+ӕ��b���݊p m�p;�Y@w*��&�z�۳�+�������O�����HD�}���9�J�\Y}��~Xh���=�]�^RZjouʔ�@$� 
R2~Wͤ��/wd�� X�_.�Ք��J����/�)��Z��1~���|�T�nI$�$u�$�����z6b��J�@�����)/��s��P5LY�蟪3��ړ��
( 7 t�k[C{R]���g���^�j�HD�}�|��yqe���r�$[��^cf�j69�+��U�����~���j#�c���:��9I]R�/f���y"N�}�  >|b�E_c����mnZ:�q 
��ww  � ' c �    0 �<  :�
���   p�p    � ?�� � 0�Z`=T���p����TmG,n�a��շ4�n����{^�\��6����[wcy{8�س3� �Z��U�.�u���x
�;�YUS�m�B�rW�.o��ׯ=�vw{6�X8x*��� �;vO7<i�V�ȡ�S]{����-��������m���.�wu`nnי���c�P'PUm���6��;m��{p��ݼ]/7����׹�m�oe@��F�og�s�u�2檷;�eUTVU[�)T<vg{m���ײ;���������wS��w���{�[]̺�f����YKm������{���dmٞ�]���T�˻v��������m�K�f.��ַn�x=L��&3˻7w��<{����家��Wos�;�V[=�                                   
�T  T� `        � @    ���^�           U      U   *� �  qP�e�iK�񋭴   
�    w   �     x ���U       VP�      U     *�   @�l�U�P     
�T�_�� +*� �  l�    �              w   [   �  �  �P    �� Wp � � U [��*�������M���ͳ�7��ieG�me��P������������� ��0 ���U�{oj���]u��US�8;ժ��p���������G�Zڔl�[��w6��Ͷ�5�Lv�9���lg���a�M���ֻ�qs׫@         
��P  x *�컡�@��@ �  ��  m� 
� *� PU/T 6/@W�R�z��s���=��ww�m�W^��� w�UZ�*�� UWv/jnmPm��
b~� �{���&3 �<�)ѷ1A�R�@����_��>z{�m%��l��JR�ܒHRn��3���K�4yJ_)�V�Y���{���R�$��_}󘒯6��7�pק�I`H�(��a�Z��av{fye�0I���T�w��n��5uoN���m�k��-c��� ��>�_�S��*�y�4LY��=1�)��s%�k���㕎��릕����V�OĒI`�ꁪbϣz~����M\Y�:f�R�WXN�r������%�զ���o+�� �I��1I<����պ�i78ޮ���;��{+eT��Ke#�m�4��9 ��?y%�ַ�����,4L]P�n�^SD0I���T��;&�XB��շ��R�Ƞ	 �I�Z�כ�τ�V��&�w�Wt�"&,߶y��-M_���f(4K_(��m�ok� �@����޺i`����ꁪbϣ^�c0���Ş��h�)uM�������y��1�m�Q�I$�0�W��M-L�}����ŗ�OUa�b��cvj�̬!�Ow�s�73����� 8�p����5��w�5L]_��V��&�(�H�C��F�؜#Ο96����y��v�ݵ^�9/;˂�p m� +Ԭ�;�*TN�mo���FQUt.�E�G[��q��x�'�c!��6%m��AְӂU�(��}%
�F �i2Ҭ^U�]7z��j��	=�8�O�K��Ȣ�,LV���Oy���I|鍊Br��Z�˃�l�#��d�dk�"|xSٔG"�v��SU��V�٠�󡠒T�����0�XdY�=|�`㧈��$�,g��8y¶��#��~AHR&�RT9H��V�u�W���36��q2Om��
|�K��<AL�.�<-��פ]�{���]�n�7\���WV�'U` �-���^�אI 
Tˮ^X�*s��wʫ�k;��dq�|��a�¹̢8��J`P�$�baW�*�V�k�R���c���{�t��$����ww����H�m���U�U��ކ��<x�]���Y��d�۫��~gk�+� F�H���_/�,��e��
6~Q�`�/��8���S��b��;�R�	$�@ ��(�:@��!l���aV��1���g�z��t�#�'�����Ն�nվ5�����u۷� C�����UGp�
����]����wQW�Z�@��fV��#H�9_�x�ܲG� Jn]g#���<�KD+Wwq� ��V��v��]b�,T���f"�Q騲0��[,�(wa5Hh�7�$�Z����b�^@F�P�p��<\��8�[V8�>4fm�o�j0 #`K�^X����g,�eM��F��
�J������
�\��ږ�H�H^+U�x�'�`l��Ի��i��l3�O���_*������$���I$�{   c*U�֕���� 8@U�{�[�p��䟻��[oY������ܺ{m7j��;k�w.��m���t��
?6��n�6�P-��@       �U\�   x  w� ��M��
�lP��
� �  6¨ �P �
�m��6Ǫ�;�q[l� �uvjW�^۹}k��w 0� �R�+��~J����L�v�n��UV��dY��'��ϰ���\�Q��)��-�#�aV��/�[h�v.�Һ�j����g��0q��x�'�g,�qV��#�9_�x���V��(J-*��U��B�Z�U��������:�X8�<Aw�a����I  rDG|��vs���f&_f��%v�j�w�e�i1E}t*��I(:��r}�2�>�����˨�^Z��t���H�m��4�jz�n{u���l� 6��J��S� ALI'$?FےI��_v���r믻�I�]E���s���Ek��G#��יo��ӫ���2�u̼����3�n������HB8ꄾ�1�]���~�z����I=��)
��A�7$�H�q}ז���fwk�}��z3>��=��J�� m� (J$���ޏ{;|����=���Kz�^�}�{$�I	$��1��9��z�w�:�u^�@T;��]ʩ�
�n �J���6�@:Qr��o�����ߺ����-�V�x�󽠄Ο�2I`6)#��]�ǝg^��M�j�t~�&];o�(r�+��� $6���3�rv�|������#�^��}�{�� ��Q��$�D�Z���)���b���2=�n���:�\l����~��jy祰T�<vX��]�ڵ�ۃݯl �����ݲ�^��c�w��n� -��g�T��T޽���9A �H	��w�������2��Mu�����[3���T�Ґ 9Fջ������CObx��X�_�������j ���
��$���k!Y��sVt��:Oj�t�C�6"�Y��i�s�Qj�3[��`  i*�ψ�&�c8Y<$���Hg�U���y���a�Y�r�%�S7$�|��W˶>��V�YilՐ�,��4�,�gHM��l��0������	�y[�w[x�nl����U� m�p�����{�T����w�ƂIP��*�8�W˻���Qb����g�t�Ռ�`�+�U��ծ/xt���� I"�UkTS�c�,���m�3����{n�!�O�������w͛�F��HJ� 
���jgH\�R�C���p���۬dQg�p��`gK:D�IЀ�D$�hc��kUZy�8���Z�d�,��c��3���x�8Y~;�PrH$��8�G|��U��JVȲ�3�c�,���m�3���������^[W+���I$�I$�I *�@  ' cU�S����j�uP<��{���W���D�)���Ӯ�S�VW��{���|r�Z�J\�׍]�d������]}�����+9�       *��   x  p ��T��ATw @ �m�  +�TU �� ` lP� m�򨽺�s�%Jר��ݽ]<�V�;^��l�-��V�-�S�T�_��ڶ��o/MQM�v�w{��?j�Y��匆�#㶞�,�4���7�a�Ƿ���I`.Q%��^Z���5Z�VU�s#��b��=�j�Ζ|G^��_3!3U#%�f�c�9�,�Hg
�JVȲ�3�c�,���z�֪�v��S7NI$�� awX�!�X�X�di�Nj�D4��V���dx��[�a�x�2�� �7BA�-^��S~�r�H]�l�A��g:�fE�CeɊ��UkV�����I$��I*Cu;ob��Z� ���R�� AU#m�1o�j0 #`G������x�8YW�
�X�D:T�ԭ�������%Z�>_*��py� $U��3X�#Ǆ��!�����;���*M"�0Ȇ���m�K#�9�t�PI@�It�{έW,Siw�X�����2��N��k�/L�N�Nu|�W/���I@ @�;TpB0�����!��p�0�	yc�x�t�<��#:ԶI�E�A���L����/�m�z��Z���N՝���UI^�x>*��c��s�*����I$�$�@��% 
Ulw��������U�F� *�\�aR�"d�� �#��媯��%�C�`�j�E�g�WX�"!Ï�{\�/��4�=<�"JzVJ�I!_/*�x����ʭj՗��t���x�8Y���S�=��͝�/� H܀�|���>}�r���y&جf�_��>�>�q����hzn��H�U9^�XZ�s4(Ɛ68������9׈X�jFyu�{�!��3ڲz��!�1�DC��z�������IPH���<�Uy<ߎ*�yV��wZ�b��{Ձ��Q!��p�7W��� [G�]�e�^ݷU�\��s �m����sU¨*[j�kٽU���A�2��_*��w��FZ���rY!�a�$��� ��ewg���p�[=��*�F�(�]]����Δ�c�P������2,����!�C�g�d"����Un��$��� �L�����/�>����F���.;�qq�1Q��ά��;�y��uj����PM��D� ��V�j��'.1��:��y;�M#13MM9,��0���z�d5�B<w�ڥO����@?0��yV��3������Δ�c���Bs=t2�}���=μ��'}�I$�J��)k�y��2��իq� 
������ K���U���m�����M����y��:h�kj��F���!��.5&*6!Yf�"RH Gu��G:�[;�5Z�^�4�X�D4�t�5J�FZf��rY#W._*ͮ�U)I�p	$��$��V ���'j�t�b�T�z�`dm&t�<��jhi�C!���,蒈��IȔ��:�X����;�S�Q��m�DC�B�mC�֠�ҳ��2U��l��*�Eq� H�֪���|\Ձ��Q8^K6�F�0T��s��r�w���UsPc���Ɂ@X� p0��N5^�U�x���
��L8]�������d"�}�n��{m��g<u�9���"��^�;��=�#�/�������ݪ@       �  �  � @m�"� w �PT�     P` x@ U   ��J�-��G]�V�7��܏�[=;6��{y��;� m�p�o�T� ���}|uUi]UR%V�!��y&جf�G�I�u��/.W�^F�t�5�5yS7���AR��!$�HGW�֪�(�^�0�ac'�c"�3�C��h�qr�Oy��G�j�+ɽ"J�IP0!_+U��r�Us��y�l^5��g#uS�k�g�D:U�~��D��$��Uq��>�d�a��vI�+�A���NՐ�/����Z��W�o|SEQ�A$� �08�j!�,pV��#<�佈i��Oj�E�f��r���l� ]*S�Y�������v��k@�m���EQTw
���yjk7r�ݠID(��u�������Z��Ƥ�*�#,�9�E�Q!��qj�y�ݍ�|�d�6�$�1�U�δ�t��El���L�SNK$3>>/d���k�x�;n�!��%�Bm]�I$��!N�UZ�����Vk�s�*X�j�i�3�<��"X��XȽZ��obFB7$� ��ˍW+]>��v\+da^~�C��M�k�#,�?j���X�C
��ꉪ�����3�����gX�D4�wUl���3�ji�d�a��<�lV3X�#������� <T�����]ܾx֝� 
�� x/T � 
����b��l�I"P2B�
��ɝ��20��I�X桨����r,����Os�U˔�t�� jO�#�E�f��r���a	��CZ�#J�u�p���,�q�T��I�N8	q��o?�αQ��5����S�g�"+ Q\#-3MM7�*�˗ʦk��H��I���^�e�._m�CD8�T�^B�24��I�X桨����r,��������I#m��V��-��нUq�>u�ܴD8a�.�T9"�!�s�hd^U��|��$�B��mD�J:!�^kܶŴ m�p{%@�� �&��F  q�1]r�Z�Ynj���Sb�h�F�2�Xξ�X��'Wr�����x)�CI�%�&�	��<�lV3X�#Ǥ��h���+�^F�t���5�1��*��  ��EW�֪��m�؆/'��i��-�DC�B�~9_#εW��썢���I"*��d:C��I���FY�sV�D8�s���ϵ��Y�eu��C�C�ψ��R��T IB�Uv�>�?@�a��K�=b�Mb����!�^/�ϝK�U�˅��$�I$m��
�Fm�wy����^� �b���*�`P�bC
p��C�����ƢB�+h,�#|��zE�<$��d^�h�4���"S��T~Wj�H� 1�W�U��<�U��מWڱ�/$Ճ��<GS�|p�y���eG @#rI$��U��ʙ¹�|E��E�YtGY��m�ƨ[�w}pכ�-u���H� ��]]����D�c��Kw��2c|$��/Zγ�$p\�������8C�~P;�-��1sՏ۷��������m@ 8@z��x8@ �+({�����=e�R�t�xolpۮ�V���
�[إ�{�J�S��^�u�y��h���N�n������i��@       0      ;�Tz��A^�le  `  ꂨ �  � T�� U =e��? <
���ͷ���n�{7n��N�e� 
�l���T �p�USӆ�u��m��U�?��ٿ��7��/��|���x7�2�4ߥ��
T��9C^o��=+��tO#���1�ι�ۘ�*UHԃi@�8G��ܣz=������jf��fo���|��m�1P\��n�U��������[����!�*�M[#-q��Ӳafx�beR��"�I0$��
�W�;��/P�5����c#K8T�E�r���&9Z�C������� ILCn�L�)RI!��k��X�� ;���� �� ���� I 9#sت*�����WN�G�w�#K4Ӊyǋ�q�#��|aϋ۵b:d�U�&�n8�,��9�����22獳�����WP�D<D9�����Fb񦳚P%�J�  &ZU�˗ʶ��(�E��_.���!�^*��X��,�Ri9��u�L�bt|�#qID�)!_+ZFyu�{�!����d#-3^\�H�,�}�<_�i&�ު�jfI '$!W�ʳ�#�إr�Z�e�y�qx�C�w<m�,��^���C�C�.�_¨��������֣˻]� �b��E��=s���Xݭ�ҐH�H��U]�Gϼ��U�|C����j�di�'j�t����K�U�˷�N�*uH� Sa^5�9Z�C���Q佈a��{n�����.&ܴD8a�:�eJD� I$	q_#εW��{ʯ���Rb�b��g��X'/�q��j�����v*�ƥ0$��
�D<D:TҢ�FZf����0���m��kdx�d:C��dBP�D�)$�	Z��W���Y���i�!���.�/bD0��ڲ�z������$�I*0(CLP��W�WN���� 
������U�AQ�D�A�ӑ�$m��\�\j�Z��ڇ!�A��s�J���PL����=�j����AH��AU\�+�kU{���
��+�+�s�Y��ji�d�:GI6�c5�3�r�H7E$�I �A�H^�Vk�3��
����wr��r��Q8��p�/�'t�������i�@$F*A�/S5�8[���Yd/59j�o��ő�_.��Tq��������3$�$��Gu��F��G{���W��r��z!��6*6��L�SNK'�Y������?����;�5�ۭ;��t�޻k� a�Y@�
�l;͝�S� IE�-֯�����
��NW�^~g
���P�CHX୾V�T����m�S�	 ���V~�/e�22�5�8[���Yd/59��_��9��Y��&��^pI�J ���W�&���k��l嶺L��O��臏�fA)\#13MKq�N��n	(Z_�j���J/Qn���Ob�t�k�T�����¤�,{�F���n���H  ���|�j�K؆�O	������m�G�,��*��~�>"�\�^�}�v��u��
e��     �p0     `U^�^ N �    �   	� N �  x   `����� c �U
��P*�[��:����weeSm����"��Իm�6[���;{������PWt �,*�Wu]5������ 1�y�eV���wQg]=�<!uϫ���� ���U��P�PN N�8�� ���ۧl��[Ұ��
�zސR�Tz�B�@�{|7{ȩ\�U��f�YZɕs�
����8�گG{�U���wR���j�Mݱ�����ީ����w-�����ol*�jb֭uݬm����x��v�y�z�&@m��{�d���s�r��U���;0�g,�,�&�]w��=wn��ٮ�l���U�ý�s�v�{M�ݻ|��oD�n[�ֶ�f��޽ލ�                                   m� T�Te;�          �     P    �       �     < @   *�  
�  �  n�6@� ��ص�   
�    w   �@     *l�    �  a�       
�           
�*�  P  �  
� �   �   d P          T�     =�    �  �  �  �    J� U x   ��
���kKm�q���� m݂��+(-3B� 6��Υ:�U��߻�wm��~ 	�  �� m���Cbg�޴�ڢ�0������6/UW-=�;��c�6�@Nz�B��E��V�;��YEVݻ��]�y�'+Ou�m       ��   �  w  ��<PU�PTm�  �T �  @ U �UU�<�U:����
��t �]j򢷲��l�1��� �J���S�T-��Ǻ��ݟm��I!}��׈��)\�jՓ{���<i��;��p�7y��3���I벩D�I$���]�Gϧ�T�P��t����&~�'�c:G5�J���~�i��Rq�@��pWY��Mi�YFyG��,4C7�������SyO�j�_f�L<�1�H� �P�q_#�W�3Nu|�Vk�mu���,�5`�i�!��p�7UdH㮤�D��I(l�_��U��������MM9�a��<�lV3X�=]��u�7��:�$�(h��Q�HU�����l�ݷ�= ��
�UwJ��
�W��x��Ub=����sM��+���[y��X{�N떫>u��� �t��t�k���=W2����y�ɻTz��|�s���ޯ��7d�F��$�&]����{}��ޱl��j����ݹF9{>mR��ې#rH0�o7�枔O�����)�d�{M���f��C���$��#���0p�,C�B�mC�֯��~�C!�[��:�̟���ݮ�I$�JbJ]�i��u�m�n��un� l;��� ��W�t�Y[Y{S~���Ƣ���|p���S�g��*ܢ-��x�{�}9rk�ʳk�m�"!���]j-�y}]�s�^U��Og:���0�£���3M o��X�jDo��%�� I�Is���]�;�/U�!�ܿ����[P�5�3����^U��w������m���uVx��sV�D�����7UF�P�w�%\���!NUw�o;��2���U"Uq�<�ɗM[~�;.�.i�Je������ϻ����I$�I%�9��V���M=�w^�w`
�b���Tw
����l�����;�k�:�7�����1̑�3؝cZ�[��Hz,Pō���ޟ�R�$�FrB|��y�8L��~��=�j����x�8Y��}���u�^V^�:*n��A$تY;��rY!�a�d�u�����;n�#��T��24��9�MzUF�I 
o�����=!���(�^�0�a�5M8��L�g�5/{�U�˕im��QJM�$�(ҵg!�A��s�J��q�1Q�:C=�y`qx�C���XG��T��o <���{��w��Z�g]��m�� 
��T۹+2�r�
���n]9��$m�I���|��)�:����9M8��gH�olVq�C�(9ې���O�BnI$���%X�H����5D!��:q/[w�!�\�XȽ\k�8�ڻ��I A�eƫ�r�S�v�^�αW�����t��PL���8��E���Q ���T��	 `;��U�>��U���p(����)���-�B��|�z�(
�BI�i��B�qiT��qF�9�j!X�X,�����CHdx������� � �� 
�cnwkp�غU��EZmu;���wj����Z��ޞN���=��ku�]�㹭�n��<�owz�����%�n�;m-���[f�y�      *�p 
�U<  p  <
���� !R� �  �AT� 6� P @  T.`��r�s�m�yp��_k�;�^�sgnۜ��n@�w W��� 6ªw��D�#rH�A�*�z��e[���C](q��8�+��V}���:��W*�X�7��?�AP ��8�j!�K��Ŝ#1V��C=��2*6��\k�ӎ��t�|��jS�6�)���t�\�W�=|��y�TįX�F�!��G�����+P8,��s�H�
TJ�W�!�-�SNi��y-�DB!�.�8�j��y�_/*�x�y�~k� �@rU����#L�R`qx�C�˂�<E�ब�C�BȨ�#1q�W�=.�]B�j��\����ۖ[k��
�lV��^T�-��T�ow��ܱU�n���H��ج�X����܇HqiTįX�a�d�(sP�B�m	y��I$�7%�E���彞��+�2(`~Ş"�q�!�h�D0����G�b�,5�1`$6�!$��Uu��.5&*6!G��/�q4Ї܆�b����Sn��I IB�Uv����ؕj�^U��ج
��|��� S
m���yU���qJ(D�������>u�
���zWv*�C�=�a�#uS�Իz5\��*6oIRI$�� 93�Sl���z�����UR��SLU�p U9��N�A��eg>X���T�1����[��2z�v]���?rN97$�c!���z�JU��c���re�5ݾ�e�Nt��A�H�m�)�)�{<�f��s�N��ɇ��!�<0?j�"�^}x�z	��P�q��q��S輡��F:TC!�AA.��#�{��o0��X���M5UT��U@��:x��]��D<D:S�Ԯx��0�d�a��<�lVhq[�M�uv�c�M^�s��awͻۀl;��_e p[hT����f7$�So:Ok�J.�r�j�;P�h2����g�+C-K����a HR�Gx�y���1�DC�B�mC�bF9�C!�[ΟW@����b��K�x�]*�XAD<E�����N��C�C�M���3\�,��0��beR*���I 8H]8�y}]��|��.��a`�4�ң��4A���c��"�oک�T��J�IM���!�cD��d^��xD�DC�B�Ct��b�O��s�^U��WrI$�I�c��������e���zѻu ���*�� U�*��Z�ٽ�.�UAa]VF>3Ձ�C�\�^0�����D<D:S�4nx��~������@ @�r�����.�u���9�Y. S�b�24��8En���L���o�R7 �I��Z�3ɼU�!�x`~Ռ�����D8a�.�T8!�a�n�B�Y����B���o:u��%j�X�u�y�8��x��k�#5T�:���mi�4m� I$% _*�t���tH3>!�b�+C�����d4C���JwX���jQ6���	$�I$�   A 궲\�ں�J�@U]"Tj��5学�ŕ���D'n��i�y���vm�u-ꯛ��{���WW}�        �  �P  � =T�op*��
�  6� Y@*�[` �  J� U+�M��V���� 5���T�9�{p����PT;��p� wP��{A���PwU[W߼�
mX�,g#<��X��g��XȽAj�1�DC�C�R����܁��"�v�ZgU����]U�F<f9��(�����a�^��ob�Hp� �A�_���\t��ѸFb��%���M�Xu������^U��N|P:���I(i�S��^X��r��]a�
��G�����*Ɔ�5�C�,d^��{w��	$m�I.S�5\�r�S涡��#
�J�2!��]U�FX���>u�WޒI$�BDq��U��;���t�� m�p{(S�5Ҡ	�k��g���*�߿�~�#uTju�"+$4n�za������s��^l☛I��D�V�82{���4�k9���^G�z��j�/T�� 8~t�"��xG-a���qT�Q�q �Ua�����ERC�������>u�.X�uW��Y臈�J��f!�¦�,��*���S5&�� IEӏ��Ր� X�6��#O+�9�z�S���V�U������I$�P��V���Vۜ�}ڋ� ��*����AUR�nl7n����W6z,"0Oj�E�P����[P�X��+�*P�t��D����I��+�V�|���>*:����r�y�D:T*����#�dPrI$�&U�/._*�������4�G5d:PRA�Jh�T�+Bܔ�yb�}���t�꩛����  M�Dw��*����ڭZ����;d^����!F����qS�bk��1��$�)!_+U���P�q��1�XAE�*a�x��S��s�W/.����$�H2�J��D�l�n˸{[�{���*��U x AS8R��I* '��]�~s"��0���6�����欇H��=�ޔ�W�/..�җ)�lr8Q���JC�U�+V3���&�V40�Y�:�dn���!�#��Z�A#�
0S�8����W�L��ä8�RT<D<xɳNQ"����{ϧ��e
4��$�Jcr�=��Sb�p��)�K$3>!�b�+C��'��]d4Dh9zMa��� �d�*����f����G�̞���m��]o���gݝ$�I5��U9�[k���n�k�>[w l;�/YJ�;�Y* ������Sbꪄ5�i�^=(M�a�J�:j�DR��Λ���w��\��T��F�#�ً�W�\�ӒRwg���ryܙb����t�"���L$9�Բ��Jn��s-�m��wׯ�_<n�Rc��H�$ I$Iԋn�������=(M�a�J�&9UBYFt��U[�H�=���Kv]�s�w����"΋���}����^�T�I$� ��  x� eS�ڷMV�˫j�wv�z��n�����Z�@�������v�x��NݝY�����-��W�m�^��{���n׳ӝ��        �  U �P  w   w^�B�*��  k��  ,ڠU�U  *� U �UU�yT*�ͩ}V彻��8�e^��w]��w-���m�^@�6�m�@
�UU6��ۖ�-�*�PUWu^��sn��
e�M�1�Ͷ��<l�隩7�� 
=;������f��*d����a�J�"�/���H$�r�Wm��;ϭ���N��f���g�w������7ɮ)  #��}�;�g��뇹
��-)>�q�,�8=���iC^arj	YY$�(T!z�b���m��U�W�[�w�^����)a��#���<� J�y�ll��V'�N�{ �wA�T� UT�m�w���F�#Q��!W�ʻ�:�QX��,SՂD6 ����a�7UNS�!D6��t�T���$�H+�Wn������C"zvجG��ͺ�h�-��r�z�/.���d�F�
���\B�8+V3���M�E��>�N23P�<#���0�X��(PF@�GA�WV�Z}�s��j�A	DP�!��c��H�#�U�^0���obt�2 �F�*��E�\t����/e�(��0�&I�+�ʼ���B�
��gQ���I$b4�ƥz�V�QC5��@l;�m�@w U��Nn�owk���w�6�F�t�ȡ�C!W1Z��7�/&�V�0�Y��q����=hT�E]����U���l��,���'��#�X��j,�H�!�(q��&�8$B��Z�[�A &�ⵊ��v��|F�$���ͱ�	(��L0��l��*�^_d�)�($�H� �H�wY"�S#�9���L'�����7��C>k+�!:�U� �h�+�W�^U�v�j�Z�ʞj�#�½ҥ�H�(�D<x������w1on�ٮ��w=�^���� 6��J��� *���
��Wwz�Y�ʏ� n�w:�_*'Q��>#|�����"+�j�k��GY�S�~�~  p�U������t��,e���i����h!�:�3U�U=��M~1QQ�@ Q��V�>�MXȽ@xG-�Y�ڇ �"g#����Sy4��  2,�=K�S��H����׋<F�rx_�U�j���]��|���wb��4�*���U��t��9�+ �4�t�XΛ-�]=�Y�Et�XmC�v��ػ�N6�PD��S�tҿѴ��iO ��vU@��
�m����ЪU�*[��dg��2�x���z����~�kV�y��+����biQ\��$%�ڻ����AAU�0�����tk:F������6[�B�$Ъ��mUA���?|�V*ɚS��+��k!�@�*ngƊ��$�A
��]��7w�	�(����&���g�I�8�������}I�D��T���7$���q�u�[�q�]o�m����z�n���-�� �I$�H@ ���`!T �w*έ�V�c��;�we۰���ݎ�/:���5��w���nۇ���f�w\����n�����{�w)�����     @ �� 
� x  � U ��
���  6�  
�  �  � �   *����bTN뇷L�]n���U6m��;�[ݮ@�� �����@�m���W2� ��&�ty&Vn�����}~��绵�A��$�F�)�����n7�s����I1����R���UZWwUU���)��R��d�{�}�f�tG$�@@��׮f�;��ٵ�/���+ｻ���	RH�$����U�K��W��Օ����サd8~��ʿ��<X���U ��t[���s͎c���ª׺�cU;��*����ww���#R����Uz�;�U�������,�ҥg� �hx�||o�DD�r %�*�T�kW�Y����V(�f����*�����[%�($ �I a%]Wʼ��{��~ū��wc�i�pX�サc8~�^�R%� �#��b���;�/�K���8���qb����J�1�������ȣ�@ 
�y|�[}޺�Uj�r�����}�Y��%I$�H�C�+�&���7��m�ۙ@T;��]@� ��  ��(n � B��o0uC~�0����?q�30x�>8S.�UX�Lt�6�7$�HԔGz�~�G*��8�I�>�Β���G��ŏ���Qwk���F����~������fɸ!F�N��\��K�^U���T��6��	$�/�#�#�<~�wB�#�i�9����it�u�/����JcIQI* V�2!Gj�p�fG*�C,�jϨ�:L�2�gK?0�ڪ��Th�Tp�����ݶ������ݔ �[ <���^�{�*a]Y)Z�G�¤u�~d��!��&��24�p֘~í�]Q@��ww#l�!|�ʵZy�9�*�mn�W�<~�wB�#�i�ͺ�\���.�(�$�T��}�����U��N��8�FG*��#���Ϭ�;�t���Z$��ےK�.]��yUok���Wʭ7ҥ�����8�t��pB!Eqi˒UL�-Tȥ�DQ��o��<X��"<Xn�Y�����.K ��~�瓇]���g���n�;]� a�*���T�VPU���zίRI$m�I$��U�R�m.�y�b�,@�(��8�!Ij�?CeG*��#���.(H ��TU���Wb������G�Nu(`A�E!�*�61o����	u��2+�� _kOi�{���|γ�EР��F�HT���޸f�Kz>�}Y������ǿ.���	( �>�ޘ$�^�
t�D3�	�eL|A8S�R��/����-t�H�[Nժ7a�0:��T   N      `     ��Pxx�	��    �  �8��1�   ;�` �	� �����ٗuT���ў�2�Uvק�Sk����8^�1�{����vݦ�r;�zZ�!^���WvݷԀ�T��T�R�EY�X�M���ݼ۶ͱ���   NU�;v�ꢯUY��\�q�0Q�mm���L�n\A��nm����o6�n���UUT ]7]��ݵ�\)Yq�p��ŲEr��NS�k�m\2�ۻ����Wf�E�S9z��uem������J���y]Z�����mwB�w����Z�����{gf:��ۻ��2��m�]R�^�Xڞ��y�ն�������ӱwM��c�������r��]�۽źז�#-�%�o�v�-�˘����ӻ֮�]Ӯ�                             P       P*�e U`      T *�       
�uP                T� d *�� 
���*�U�-۩vް   �    � �  �
� �  p��TV� < �   
�  T                �e�  @ `  
� P�    �            �    U      x      �   �*�E�     P@��.`  � �Lݯ7Z� ��UJ��
�  ^���۵��o�;��`' c   < �
	�\��&���{ �M�s[m�zz�����Us����%�um׭���T)Ui���)H�j��k�es�x�       [h   �  p � ;��T 6�UU  m� x  � 6� P `P 
�����m��I5�x/Tͽ��vwn��޼�oY�����dl�qUoes�
�q�*�qG�� �"���Z�%əE��i�׈�V�����q�󸜪�b;��Hu$9$��v�b�4��X�q|#��aD�\Ń�Պ�s�ұV*�]ӽ"Br0#p7v*�ql�$ʾ"���`�q�Da�1��#���>�J`�8�)�B!RHnI$��(��*�K5Q_*�򭙶�F�\�x�5柫<F��8����L�D� L��˫�J�\�]nP��4�G5`�8������~����V������ӷ�N�U���� a���@��Q��.�B�
5M�9カ�U��T����\E�&U�G3�����<#ٔYk�^�Y����F����.�#
�J�0'[a�m�C�3��x�{k5fe�Z�Ϝ�@"�)��n�V(9*�G$�G�(�RP��5}]��uj�W�U'��0$��
t�Z��i��Q��qB�
՜Geβb��.�ۘ�U)l��Pl7$�.�X���wk��V�ZgV#�<ȡ�������4���'��i���o�@�u�@l;�Uz�����` ��^����hQ�M��X���}��W�b��x�E��C(���:ܡb�iq�
��8�	#�
aլIWe-�j�ya�>��!�) �Y�qX�/9#)�o��� F���x�*Q��{2��a��0bC�½��X0�YZ�_*��5���N� G��CH�f�G�µ�����t�=WʅKWp�|�V*�5p4:o� ��I+�!�i��j��q�s��i�)G) �!Ij�#��R� �|ܛ��c+k^K��mR�;��{+dU�Ue-��W[{)vڂN��έV,]~����z�=�*Ťa5�0bC�½ҥG��i�5)ȣ  UwZ��*�n�,u�+���0�i�f�<G)�U�(�ʾ���T�I !E�իʾU��T���4�G5`�<D�\��qx��U	X�c�T�m*��)���$�B";�8��Tʾ�0�<fn_dZK�yDr�U��]u�Uk�x)yS�������0�k�*ǈg�v�,#�B�k�x�+Oc�hx�:_ճ�wwwwNnwj��*�^y�n�Z��6���
�*��*i��VǮ�-��U]�Wu���5/���G��8�[�,D���9��'�����E&�U�U$�� uu����Q��y�*�ufI�oP�ff��A�4>הG#g[mw�� G#� �R�GX����J0� �(����|�`�9!��f��_*��ۧ�_���$��SL��C�qҤڸE�A#��zܡ`�X�����;�U�����J�I$d�G��1����"���c#��$ʾ�0�<f�_DR��J&��        �-{�nWW�vn���۰�8��28�lguw�:�M��h�{����%⭴�N����=�uԖʭ{������u������h���v�      �m�   � �w *��l��*��  Q�   ��  �P@UP@ ��P���m�z^��r���ݫ�յ�v�˱��X wp��UPU` �
�w{ �rI$m�C�.�\���f�<��F��0��TX,��2�x�x�m���X�yS�\�w��	 `�X����d�#�����(�J��dq��J\�{�:\�$H��% $�"�_O�;xI(�Y��Rh�^�R;�_^e�7�ڡ�ㄐ�5�ػ}�enI1A]�a^�*V#�+�ѱ�a�����R�	���b����Nf���i�y��J��p�#���r�QV*�.ޒJ�I$��Q�"1I޵�c��=��d U⺷�V�q�d�2� 8S!t��*���{���N�G��=%P��9!�T�w��T]���~	� ��C��f��A���הG#��u��?��*��b��t��  ��v���<D�1`�9!�.f�G�´�<~C�qҦJ�E�yT�/��wVj�UU����di-ʱF��G���#O+��8�Hx�2m�N�I$�IDw��T]�d�:�\x�ܾ"����=yf|F�rj����߻�|�� ��p�\�{y��w���@l;�+���pJ������B���$�G%.�V㧆�#�w�h:C�'��G��U����ʵy^��EJ�$� A|������du�AXQ#O�sVU��e-�j�yb�k�i����&@���֎�Q;��U���{�O40�������+X���yD3�a����$m�WPu�+G��!��A7j�q|C�x�y��"���]�����(��� �e�1�3�\Q\#-����du�AX��*���{���}��֩ВI$�) w�w��[L��N��^�l;�Uz��������wi���W^�G�9"�����B���
պΖF�s��bD0�ܘȽAj��-��F�h�v*���ʞw�+��*�8�+�������0�|͎j�~_�o��y��$m�@M��k{UsR��!�L*+de��A�_�ه���jc�aݫd3��S4�T�Z�t�,��#O2���c�
!V�j���'&��C�s�?( � nK�]>~Y]���!t�3X�#J�b��p�#��W*��T��$�I$� ���s�ٻҼ��ݻ�y�@P��������T@�I8�8�p 80������F8��Mq�Y��g��D<D:T���z�}[g*�.U�����20	.��U�X�j�v��Hqx�������+��,tZe��r�g"�w����������וrŷ��^�}hp��D:a����r�diy������z�4��8�m�G#>=�j���SMq�����z��8����B�i�k9���P$��v�W�gu��#�j����,gH�T{B����]%c����~�w~��^��   ��p ªl���H�OqT��*��k���p)�^�m�n+�Ų����s��Vڜ3]Ԩ�:+��j}�b�=�ۻ�L7%��c       Wt   *� �  ��@�
��UZ` m� ��?ʿ~ �  *� � J��V;���E�wm� u�'n�on�7]Z^��m�����R�����E�@�JJ��RJ'ܭr���?mU�CO����L���o�(���T�y�E���f�*I%t��]ѳ����(؇�Y�sVkƚEM�0�7z/A����Ƒ�)]��$�daW��=Gϫl��Z�Vt�
��A��{.��7��s)UV!*`I* A��m���=�Owm��6G�rV5�fߦV<�XH�b��9E�n�ͣ�Lߟ.��7�������۝E}�I$�Im�* ��o&��λwwZ� ��U^���6�*��pI*NH��H$��$%{��鲨K����&�K���o��i�s��u�+j	�E$�H�(F�}[��¬�ʒ-pV�s3d{U�6K`��w�W�x~���$�@!�2]���ε˜ק9��[�Q�T��[���'V�Z�69 `�m�������y_p�d�rK�;�Ar���x�EB)Y5Wwi*���.���4�+p\z���r�ȟWǍ����۽�wm��� I$�NOm�������]�j��� d;��{+eT��QU��u۽�B�U�{c�x���~�Sf��C����J���ӷ�T��	 �@a��wT���-�`�=4�QtӃ�IrW1��; ��pd)훿ewe���k�S�F�.�һ�UQ�JB���Mi��w�֪��j��Y* ��I$�.�z!�C��;�����m�e�t��r�V6j,����H  jA]r�Z�Y{�w[��Q"���#uK�NC�C�9���oV����"�I$��F�7	t́竻's�l;�+ԪU�
�$h`:U�PrI$���U�._*�ɔ���<$�Y��x�������(7*���L�!�m��5Wv����n���p�3��oZ�|m�ʘ��Lחo�(�tä(�C���3���U�X���ۍ� �p�����x��F�#,�9���T��T�\adn��w�W�?��^W����R�$�  @��Lה*�a&PWƢ�v��Hqx�������*�%J�	��	"�]o;G:�N��:�VY��6��"`�Ld^�}k���W/.^T�k�Ҥ�I$�ȓM!w^��bR�l� wp��UPU` �
��v���U]�;��:��#J�+���Rb��,�������*����U{ϧ�zSAخ��"��z!�!ҲJB���j���0�ɔ�+�28蓵d:C��z�^�P��H� �:L�]j�-^NE��Y��"���1����fҷ�\��+�^��U<�2ҭ��$ܪ�nY���,��{q���cH��l�2(�\jLUb��=�j��x�C�ޟ~j�@ 29����^�3�A��x�{JR��2�4�*�b����s�U�[M��rI!�I&0 �  0�᷻��=��T��y��{��TN�Fz�{�wS�$��eFٝnw�wF�j�L�mۭ�q�n�ݛ���Ջu����9�      *��� � �  w
�PSc�#l `*�� 6� �{eP�~U6� P  U  T�V����wG�� 6��Ծδ�x�͊v�.� m��U]�-�S�TE����v棛j��PUV���'��?��`digJ�RXe���V�y�,��7�J����� M:�Ƥ�	 �d�U�=G�p�;�]4Ì� �ҹ���ʷ�#��W*��T�m/ϫ� tU�/�q4�Y��g��D<D:T�T.��v�yP�l�n�Hk�H 
d�<�U|��=��qx�������)Ȩ���P�w�y�굪��y���Jdm����x�x�Ҳd#u3^\M�L�!���i�!�A��s�J����f��݃��ܧm��m��;�kם�R�� 6ø�J���Vڨ*;�V�s��n�*���7����αQ�F.,����t�i�S%P�Fb�F��-��� #lR.�j�Wʲ��s��4��m�3Ds^)�=�#K8d�����
�Q�x7����rI �Q����(5�"Θ�eLdm�h�4�eΖt��r!�������U\�FrB|��5�;��ʢի/{�5�G���׋<F�lg��ҤU��6��$�r��WoP��C6Ydpǔ���i�~۬f��S��]j�-N�J��H���$�"7*�ն�v;���up�Z 6øUomTF� *UU݊��oPUm��߽��Q4G���X�FyA�M��t���E�f�OfQ�gH�Ą�P"��@r4
+�*�V��9��Y��;�p���{Ճ��y<>}��������6��%{}���u�ǵ���.��o؞xs^+hdJ���rI$�R���U壴opT��h\���V���dg�ٴ��D<^��2<�<�������6����b�:a�M0�5���UsR�"r�N���Z�e�y�g?�G�����@A	$� ?(�E&�R� �'Bc�
��U��eT򲂨�[s���qܫ���GY��7Uq��'!�!�U1J�L�PL�D6a�1�)_h2<yߨ**U0�I#n F�g?��]���digJ�Q:,2�?V9Z�3���S{Û�U�޷O�'�����FZf��~�DC�!G���F���(d:C��I��NY��*�N�p��;���9�*;���Hݕ|k�d���:U�>�Fbf\�*���L���?�d 
w��֡������y�p.j8Y�DX�Zi��Y%j�d_�=��7wwwv,�Z]v���Ṯݎ9n�P ���*�_�~ UO:�ݫ�w8�U�wKcC�C�!ܫd].5�x_y�Α�~����24��QG5�AyQ�H jJ.�U�U�z��ڟ��Bzk��3iz�>C�3�\��v�lw׼�P���I$u�\��*�[���D��<$�X0�kJ�\а24�˹T��ǫ��X%�� Wb�c!�~S&ҽ�!�xN�+�</��|Α�G4Ð�&~ң(��F����$�DwV�5���)Z����5�Mq����8��[�Mg�#���߿������n��1��1�  *�8����Ƽ�T*���YV�p�OuU��ﶶ��tn��bl���3����a��Q�n��֗ۻ�{���u���_K[6`       *��   \�  � U .a�p GpdTm�  �P*���W�  P@*�*�z��8^� 7<���@�<
�K�m�������m�� ��
��S� @/-A���U�_�����y~?_����(+�-3��	;V"���2�������U#���Ic����Y�#Ee�Ed��c!�~Q���|�~g�0w-�X�֡�}��t�#��S?��$ E|�u����G5�]n��F#��k��<�g�MMj�y��|�~)8HI� �E��:T�T.��v�yP�l��A_�2<xIڲ!���x֛
����ej�����H�L�*7�'�?,pV�g#<�zz�z/��oVTȫ�_��gI$RBII��&��-��n���� �wV�E�T�UKmwS �*)N� V����w�u�\����&9�ú�!�,�9��ƹ��l��?�#rI`�+�kU{κ/A����t�=H["�3M@�ن�e|j ���Bj�v�%wwUJ��!��3�F�t��a�f���V���dg��=u��O��}���"@)��E�G�%o�(�tä.�a�k���m��t���D�UkV������ 8*�X:/�q4�Y��g���x�t���\#13MG���0�f��݃�ݫ�Z������ۖ��˺ 
��
�R�T;��*s2�n���x n��z:�_,��B�
��ɰg�,��ΗR*���QBȲ�E�����[$T0m��;�v��o��|Fb�Z����Q�=�Nx��kdi\�R�C�8�㛵K�*�UV) �H�uʭj�e�)[�����w�˓#uW��臈�Jsԅ�/.�t�G� $��R_�Qr�V_X�#�j<$�Y���L�G#K3�;����h���55\#�(�ܒI���NFyM��Y���r�B6�>�8[�Y�:�:B�9Zg�(`rUUX��Ʃ���ծ�����;r�ۻ��@��U�PN� Uz��=���CtaH������x�s�D�UkV���+��-���F�5:�r"7X�>���ܒI Q�_*��}m�D6a�vL�|j ���;n�!��]����^Z����P7�H�%@ JCE��B�j�p�3�l���D4�x�;�2����&ߦQ�H��*�Jm�H���r(��n�W����d:C��I���FY�p�qi�����9r�^��wd�~�$��	%�g�"+�.����ʄCfCα�]j��wg�|�Y�墉{� �;���w]-���[iU�� U튫]5Q�*��[;��no=������*�,����*���B8+V21�ɷ[ζv�K��{����#$��$��r��w�m�\��o�(Ls�;Td���.b�Հ�3RWuE*V������6{&�=HJ���\���~�&���I#lHR%���<�
={�-I8+S�{/�����c�n�v� FĜ'A�>�2��.a�+竟�P��v�ν5JꝐqw�jP��A$T&��7mt          �   8@  �{mTp��=��  �	��� �0  �k�  ��;v�1�p��G���USdr��f�m���g�ڹ��^f�V�n;ܶ��6���y��Z��_�� +w�^z<6�h�T��>�+Ԫe�ﶱ��w��tn��7vL`!^���~{~߿���WmS�zp<v�*!�FdjBh����ief���ۺ����[[�bМ��S��v��5��)uUn U*�k���l���MY9�[Kd�� ����v�y�7��[�p˻�Rok��Z�uV���[:3�5�'[��EU��Z���5����Kmoom�m�t���ٯmҺ�۹��P�1,�L��@�����"Z��{~�{���.n���wt�����6����6����{v����mם�2�'y�[T�9���z�ǭ                                      ��
�Wp          �U  ��   �
�             �@      ��T   U@ ]�
�P�ݵ���   T    �   w  T ���@�      � *�U          m�T *����� �`��߫�� ��� TU  p          �  x `        �@    � T  � ٹ�     � *�@ �T���l������ �;��U�  �)�T1��ݭ���/w{���,`  ��  -�A�S����f3�d�����p[�L����{�'I�`����.���ku��S�/8��[��=l���vX�Ow����      S�      �p �U��TGp
�c l   �   m���𬢨 
�P
��x
���og9r$���5v���<�wqz��` U�
�*� 
����/�q�H �0Y_c��G�����9Ydn��=��Nz��E�f��**�r�S5�;� F�6�;�y�v��A/���q���)�T,tZj(B�+P�p�3�36�Q��U�]  iBB���\�M^���\z��*oݔD:a��a�k#J�u�p��n�~�R ��U�_,��+��-x���p�dn��S�=��J�(�ʮޣ]����� G	u�.>!��W�Zdx�d:GE☋�G�-^O��Y�#�*ҽޒI$R�#�i;�n�y�wzٳw���ª���� � y휯Y�ڪ����k���(6O,�XD>6��Lde�k�p��C�!t�CX�Tjq��M��$�F�#��j��#�ا&;L��p���^#�x�8Y��g���ԫ�������1�AI �Wʮޚ�%�l�y2��<$�Y���Oiwާz��W������6�� ]ٺ�C�E�,pV�g#<��<�r�!��w*c#-3^\M�E�0����TdrI t�E{�y������1Q�FY�p�qi��k'|�+Z��g��I$�I �@�B	,��ۗl��v�;�܀
��*�tm����*[oUP۩z��T��{��߿�^"+$�.�����b0�L�x�z��ݞw�ʷ��I��DH�*���Wac#K:d����,�B�j�p�3�l���E�C��ܩ����|�ץp� � Z.[����ʞM0�5���s�J�Rq3Ys�F�e�)Y���*��^qp$�6�WH�9F�jug���X�p��˲��b0�L�|j&G��RG"N@�#�
a����{K��;�^Zt�BÊ�EX�X�FyA�yg��W/��{�%I$�IR9 a��n�c�v�oh U��w�T � 
��R� ��Ĝp  !8K�W��-�,�HS6̴�ҳ�D2U���蜪֭S�5O�� ��
����^!��p�7Ux�A����J�(��f&]��X��0�n�_RI�P @z�=U����/��b�L�Yң�E����Z�U�U;�|4� p 8~a���q�w*c#-3^C��E�0�
a��9��y�_+U��\��T�1S�#nF!^��W�/yJ�~�9��'b�p�7Ux�A���C�MR��2�i4������v���S����pWu c�
�P w c6�Y��[ H5'��\�U��9�窾YRv��Hqx�����,�N)BÊ�s�L��p����rI �Q굪��Y�z+"6��L�e�kˉ��C0��⴪��(�oL��L�UI �|�V��w[�j�Z�e�)Y�M#���8x��^k�g���U�E"67$�H���W�vΕ�-L�ǔ��#O�~Ռ�׊`�h�F�V���t���J�  ����h>"8=[XΖFyK;!�!�1�ʙ\z���wZ��yU����PI! ݈ 0 
	�+k'���<U6(�r��� c�أ�s�U��ªS:�'e�M��6�V{��i��iҌ"R�!�SDR�r��       ]�     �  T:kCl `*�� 6�  @ �� ��U  �  U�<Sr�ͰU�6�K�^�c*[e����jێJ�l��� U�Uk���;�yAV�ul�m��{�S 6!�L_�U����U���x�Wx��*���R���*��yIy�~PH(�$�E	^�����ݛa��#��+��4�7��}�9��|�2$�"�I$�R���^U�p�WE��"8=[X0��	'�x���]u⫏��|C��F�V��x�	�f���U��X��q�1T�V��9J�_�����7 H#l+�������3�Hdn�[#1x�{6V�ժ�m�|��)Y��$�I%F�T��*��֫�S�T;����x Ag[�v��P���uw��9�)�=�8�>8\�DX��dLpV�x����<l�D��QPAcc�r0N�UǈZ���u��Y	�f���U��X��q�pU�0�_f�LU�!Q��7�
�9��u=7����O63�Hdn��Fb�6V�ժ���p'� ��Ƹ�Sی�֔��ќF�fI3��j����WV�T��[�5�*PI$�S	�Z�Uڮz��1�]F�;�_o�ڋ��^O��y+ܤ��IN�m*�jj�kw:ֹ�z� ����P w � �����
V�X�Y�\��)�z�M�>#1W��X�/*�H�MUv�B�u�U�$�H�!������|��:G5�S��x�ʢ��J�v���m���h7 �
�����ww���^U���\��7��6a5{C8BvY�4|F٠��J�����#�V�5�7��"���kM#��lY���˥�yV���?ͪc�P `A��ƌ�C���z�)^�?a�헌�9�+b}���j�ܷ�I$�I$m��O�����rZ�wu�n 
��*�tUF�l��ѱ(�9�����$�uu����[��`��/S�,������#-|������j�w�T��d�F���l�4~��%E�������|�M�+�~B���R����~a) A�$��~�I��S\~B̅b�\G�������#���y-�*�]�� �D�9%_�T-�z�W��홥����S�w{�_����Q	�?!9���R�7$ �E˺��U���_���ӬG�x�eW�~��͍妏�=S�< ��q�ݛz��w��nӽ췺 +�
��U]�T
����Uw�y��($��_�H�ǼU��b��E1U��d+�x�<���O�n�kn@�� $�J��i�O�U���[��0��)��q�I'����#�(��)ө$�('�P!rE�?Q��?^=���t�k�HU|*�w|���|@  �����~B��lس�f*�\�g�̂���f-4{��*Ŋ�*6�����P @!}���e�iNʞ��a\n��氋��qԭ_*�}��ɸRI$�I% P��   ' �M�ս���j�S]G�������n�k���Z���*���z�c����[jm�Gn�ɮ�u]���ާ%m��h�͵        ` *��  {�  *�N!TGqU M� @𪪪 *� ?��    ��b�T��mg����C	�ؘ�EB�ЪEL��w W�@� `�6�犥@��Cؿr��R��x�y�����V(��X�����]�[������)�� q��/Wg)_k��Z����yt��?2
i�|FZ�F��RHx@ j]j�^U�ls�_�{3�-�t�^*�S�g�E��k��:�6��F�:����n��Df�B2׍Md��q��<,�"���#$�A�r������+~����W$/����y���I#��$6�Wٖo\kgy�;�Uܯg� T�����-�QYAV��ݨ��������F8y��,�����|u<��_�T,�y?�t6I"@ۧ]g;B�.j�?V'��Y��"3wS>�Zh�*l�U�ʾ#y��P��
+�G�2=�X��׍HU}Di���U�k�<�E�G}�0�0$� �R%_�ʵR3ES��Y�%b�_�2y�c��~�_�]�:�������$�h�Wv3�iy�J�E��:f��X��o���_��j��p����N�$�A�]���JWtn[=u�7=� P���T � `l�]Uw1mlS�wZ�W��+Z3Mk~ߟjy��
n����}�ےH���ຢ��>�����t/륦�u��#��2yH���7o
J�7$���]��8��eg�c#H�$�V:,0nq��/:��b��Ջ�r�<p�D��p*v� FĜ%����;��!�����aWΚ�~�ˉS"�|����{�t�@��D�Y��^#��g����c'/4����^2���Z�W��b�	$���؊(���W{���� a�_e�;�Tm��q~@PI �i���_.��o��ҝ�6�q��V:,4Y:��\���o
�)$"P @IU�8C"<WS>�]�Ȃ�L�~.�7��/�y9�|�W��x�y���� ��͊�B#O��08��x���b��i�h�ժ�K7GS��`<KT���I.��]^�2�v��dh28��w�]�O��dirR9���u���L� hc��Z�y�w}(���38��������02�Yf��q�W�� 6[>�ʫ��4W�{N� �m��u�Q�*����Y��&���HlnI$�!��[���r8�!��,,�#��س�f*�>�j�*�Y����UHD 0�U|���,2d;sn�4Xɻ�����i�K�^U�m����%q��Dj��"M^�bE�rOX�C"sWSi�!+n`d3�J�n����D� M��5֪�{8�^U����5��o���{ݏMuߩ��u
�� E$2�E&j��Vɘ�������ھ���~�<�v��H�I$� 8J�P   ]H]�gw��ޝf�9���Z��-��<�����μpsT���Q�;�W����ۻ[&��SM뫭x绵�nU��tv��{�vަ��      �p     ]�  �9۱
��;�V�  �     -��T *���J�  7 �kfˎ��P7]����˷yݴ�gO^�z 
�¨�Ue� AT��f9{Sa#l�d����w��:�g?y�������"�9'�Vx���˩���M�+Z|�Ĉ F��]��\�S���!��<�����
�CGE��qg?|����6:mHI$m�@+��U�>�G���j��ESUKy�*��d2��sn�5e���2��*�ܒL%��ן3j�aW���E۽DX�U�~�!bE�rOX����#4v�	"P��Uq5�3�C8Bs9�Yg�*ܯ-�t����ؙ��j�U3��I%1	Sl�)�M�=�W-On�l;�+�(� `ܩ�n�Rت��S~���<����=b���|3Y��ݔճWc�ͷ?V,U���&���($�@H_k��Um��^-f��u��J�~zH���U�?=��Y�tR���@��pa%����SW�	�d�1���3E�t��#�x�F�_��UPI$n"���V�3����G�,���[�����uΈ�����3Ki/$ F��w��yW��u�h��ܼ��-Rʞ�ޮn*���d�]W�I#��$~n� m��ݮݳ{� 
��UU� *�
��Uk�ˠ(�Sq�*I"�����N�g-�*�Q+$χ!s�f�+��8�I1�F�
D�w��}�ܙ��b�]"��h����ş�*��k5�:~���R���UUUT�I�]���+�q�<�۬�Y���~�é�Y�:��z�P���)�'H��$ۅuC�V��\~q��Y��=b�x��N�*c"�6��F�&|8���r�
8r8"8���������o+p*��Ί}E�V|~Ʇg��[��%I$�HR�2�7�QD5M2��L��Pl�PxVP 
��a�P	$m�I(a_���i�*��1w+5��8�nm�F��ɹy��<���ҪA���$�F�rz�Pg5�5�����X�BȽNI��8~��8��W닺�4�d�($�+/3���\�9�,�\���t�r�V�U���,�<����A�wUWBp�NQj���{ѫ�yW�3ESU^.�f�⿇����]d�� 9D�B�6�n@��A�d�^U�<��i�J�5��,y��g��b�bE�rOX��Z�P���$�H�6�8J��N�m����q��m]�}��� �m��F�*B��HE @Nڪ��\O�{�>l��(s���ܭY�=�y\��_�S��Ц�)   �;�E�V|~Ʇg��U���x��:!��lz�7����u\�@��7/��ڠ�=C�Nj;����ȳ�`�]?18� 	(���8��n�2�&WG<��[X0���(�/��@ 8Ɲ��=ޅ׹��_/�O_�Eҭ��H玟�SM[#-w+2������   @ � VP�rεٶw����ԇs���<݄z�͝՞�uv���l�[�+w�8m�Wq��]ۢ����Y�ݻ7���h�\��k�^���       -�� U  x  p��
�q` �B�� �   �P*�T� T ?��  �
���T� m�r�w>�2����͕�۔ U�Uk�Q�*��+Т�i�0Hq�	���g��欳�/&��$o��T¤����j߼�_/כ�Iz   ���Qo$���?��_t�h�hcx>�$p�z���n����I"��E[��M�L�O��X5� E2��.�k{���_�ټJT��$� 
�U����x�}%�x��z<����XT���_���i���n9H�r��������&ۯ]g���ӫ�KM�w��5_{�d�$�I�5)�H���J��g@TxUw�P�@U,�`8�!	$��۔آ�B�\gTX,��������X5�ma'���y<�i7�$�$�$ ���~�΍��q{��7���5��Y�����*���>��HI$m�@DNH3�rb�r�V@�4���+���Vx��#I�?�q;ǥ�I$ܐU��N�C�j���6S���f��V��|���ӑ�$��ۑ�_�U}�K��#�\�����f��x�}%�NV~��w���V�ʪ���zl����{^� l-��%P��m �ڷj:@�� �K�U��gZ}ү���LX�[���,�����~�Y�0������48�$J B�!z�u��%�P�(��(s�������Y�oS+W�^�t��p 80����Z�<D�����B�⹚���b����Fm�~��w��M/˧�P @!wk#VC(�2n��7�ڪ�NX���6��>k�Vx�v
�X��f'�)�*�����J/�U[��&*��u�פ�~D�q|�NV*��`��ۻ�����gG��o��s��k�{j m�lUU� *��TVm�5^�֞�ª��s�7K�zl�R^�����-L����`��q�����ݝyc��U�㍨5�{�ZB
5]wIRRI$Pc�6����,������;���75��)*Pd���HF}��7����{�M���m����51�Ҩ�C�R�I$rQ!��Vq�fn�÷wz�LY��:�};E_v��$�I"��{��g�j��_7��� +(w6�� w PT�za�۶�Ҫ��c�2�y�呫r=�[1�S[yrF���'�^��1�9�8�Lڧ+T�vz�	Ǣ�E�{]�뒝�(#ʤ$��$��I=��6�>��K�ü�˨鷓n�����4R�7v�$�F���v���nϳ}8]����(�_b�v���M���6�.�XC/3;H�r���c��Ks=\zW]y<u����>x���O�" �~ ������p������Ȩ��<"!�R�C�$
�����NeC�Ȁ�ǌ���Ex� �-"
"_�ŏ��EP)P�������z~�?�>��QP;z;!����}~�A��������������!�}���* ���,
�*�2����	�$EC�c�����(�����}ρ��ǵA@��|�~}?����|�PDG�?���( DA@�����"����x��oЌ�b�x?����\��AP/�~=�"
��?3��G��~��|8P<���栈(�����K��~�������A@��A��<��9?s������>�����
 ����)���Ć�iOo�(,����������0*��     �      >���q���P��;��(���t�@�r:(��(�`Wl�����ЭswU��jUVCT+ ��(U�2�X�R���U)s��T� 9p֕��R��ҩW�J�۩U+�h.�UY�)[�*�����r��@    �4�&C 0L  
����@���  h    ��mUJ�  4   4 *����*R�      ��5P�Ri�      I�H) �	0�<��@ 1����O���̷�$g� @�X@�	'����@	'	�s���N*�� $��;$`H��@�Ad$I����U=�� $@���19��?��=���<g�)���db��I(J�X"����I���-���11��V0U�DTRET[P�+���TQ`�Qb"+0QX2,Q@DUR (�ATET���J����-�`���
[TDcX�), ��I	mdVD�DTR����4�ƖZ�DY%�,��AUE��Fb���Q����mT�TY��(�TX�dUkDD�H
E"�X(�(�b�*֬AQD�c`DA��T�� �,,�d��l����"�U����T�b����`����(ȱb"ȰDQdQARTI
ж��E��PY�"��+EEUR�TPUdH���@�UU�Q`,�E �E�T*�Q@Hł��Y
�U��+m
�
���J�(`P�B��HV+(�P*E�Z�V(*J�T�RT�RB�B��P�������XT�j(���ְT�X�+�T-�J�i�+*V�-�KiP
�QedR��
"	J6�B��Q�m
D��J��*�$+hJ�d�E�*�T��([IAJ�QKl���(��"� ŭ@PAQDdPY""�R���� *��T�)F�"�
�dE���?}����f�>!��~�݇�O����Ӿoy��p�(�U�P� [���T  VT������m��� +km��̥����k����}}��fո����%�,2
����mn�[;���@ 
�P  T   �0��j�
]m���  ;�AUf�������\�P�ud�T�]J�P EQlT��Z�V�<���E�1�*�P    *�s U  ��m�֏w�e-���ҹ݀��m��۠lP�le
��uT��l�U ���UP��]ٷ{�@*��R� UM�Z겁T�    *�P�� 
�d    ���   R�P �  �P[%P ��~���PU Ee   UPU �U  U   P     TP    *�@ @   R��*��l�
�        QT ����̠ �R���07J���   �Um��Fd����AU���+)R�f��ATAY*� 6y��*�Z���.eP T� *�� m� +( Y���  ��V� U ��cb� ��S��l�Y�Uz��UU
��o%�m�`[  
�}>�l� 
���U      Z�] U
��k��{�ٲ��{��LG[��� *�j�cJaWS�z��Sq5���Qӕ�kT�����Ͳ�6�9��ݨU����������Zӹf�{���Ue`nAk��$ɵ\�����;�n[[������R�2��.k{�����m���]�i�����Qn�d1m@�V) ��Vك&�Ҷ]
�Gmj�
E4�[�l�l�
ٌ�0�j�p	L� �iȐ2L!Lm]�   �U*�s <ٶ� �
�ޭ�m�� ���  ʭ�P�=n�d  ��@   �݀ }�}���-� ���VR��ĵ�58]$��\���*f��s3����N�xI�i	N�	>d�zp����0���d_�&�O�>L��A=���fw����9kmUN�+�s �mme  .�`U )��
��W�J�VW��=�YV�ޛh�� U eU  U *��TP     P � *��@�6@[!UY,��QT*T V6 �v�wR�� �N��ck�yu�e��F�-í��]v �e��S$ �,�jg�s��u��n��*u����`����շwԜ�=81�EP)Dpf�ʶѶ  � ++�UC�wo��x�x;ѐ��3)nfffU����g��ߥ��b��fY�o][��<����c6�ɲ����W��7~��>^wd�R,=�1���s1و��N�Y�C�Y���Wb(.2Y�3l��gL�=�5�CY����t�f Wͦ��,��̠u՝ V{�N�Y����v�=&0Y�����Ɉz�����:�SY��i�9|���fU�]A%١Y�峫�)$)̤��k��'հ�\`��2g=�˗LC����)551��⹜a�V)�7i�-�s2읦�3m�պ�[�a|�����˴�`�*[��d��ot59�MMLg�9��מ]a�X�:��Ma�u���VMMa�a�����NΙ�&sp��&�k�0Éܤ�lY��|�|���]�����+w\�Ox�ݜ���{]'�q���&�C�u�.�&�ܤ���W��� �l�&0�s66g�?	����q3��'�`*��U\m�x ���m�T�b��wn^uR�kaI���5Wl��d���'I11 �e&y���ŝ fR
q'��3.'s�u&3��Ncs��T15&�0]�s32�Ś�؜���ݗoK�b�j���u'��t�l1�X,ĩ���Y7ΰ�9���naٜ|�W��l7�Tǉ7w޺��y�I���m��\a�g2�eB���Ӧ�>6u�9�~�-ʪpm-v[�f�NӤ
�n���)�7y�:bM�'i���a�\�<�Θ,�+�K��w���ܹ��8��_6��ʘ���fP:�0��w����*���4�T�{���ג�bW�K��z���`q:꓉���n��{�͕8���M@�̤����N����c�0Y�^2s��7.����6u�9Ս��=�t�*�jd-f���O~�j�"��B���e�;MLf�u�1+�v�]�޻¡�P��)8���ns3a�}]a���03)�q�o�Oz�jjc6�b�~c�lh6�EmH�#��� P�h3Wm�uڀ�7p�ZJ� 9v�m�X��ι�+�'3p�{���ޫ�N���]a��S�y�@�̤���Ͷ���s�q+�O3p�u��_;�33��8��_v��b�{˻�!	X�J�I<�Y!g�s�����36��1+�%�p�=罭����551����=�쩨ff7)<��̸�'հ�\`��O��g��u \P��Ĵܳ�o9�&� T�oFfq�;��03)�;�+�4����m��$B�e �+�VN2�!iR
AM@��R�[� ���R
AN|w�jAd�T��R��Ă�P�`N��I:Bkczg>.�"�|��;Hy`J�e�'�9�qNI��rN�/ǁ�����K�ܛ��!���C�Y0&�'-��0Ԙ�#�m�́5�+	�I%��LI'����	�Y$���y��x���+	�К�&�X�&0���nm���`Ld T&�NyBq�5���7�}<�Ξ?s��x�c�3UUV!9�_��	8��8�p%`La>9��f:I'}��B`O��I9�	�����] N0�!1 E�1�+	�I%�rĐ>~��L	�vI'����@�'{Bj@��u{��`N0��I$�,	�B`N���_~m��m]w..n�����@ ���'�����z��wV��wq�iWz +ᶺ<	�v��Z@��jX���ύ�����̭���Cw�W��<P�jF��{�m��q)��  UY��L���7wO9G���{�>'Y�a����ޮ㳤��xη�T>:���Y9���N��ݺ�|��';��:3�:����f�C�Y�A�`gg�����½0Y�W����P�59�[��p��+��a��SW�.,�uN�>Ov��jcp�3a�`���f�P���sC��MML@�h�O_��:��X�dmZu��n�P*s)<���̝'հ�\`��2w��㙥Cިjs��ML@��^f[��ʘ�dݦ��&'��9�|'I��a���f%q���;����R�M�Pe�=�慓��:蓉�����1���r������rܓ�Rk
̴��M���̢�{I�I眷�P�r�}���%���k���"��d�e��T@ V��T]���[��[���=���2
����h��u5��rx�fZN����� �d�(�ͤ�x���'HV�q�:������N��m'V{ǅ��8Ԃ���QC���i�]���h:s����^Iָÿ=���q�0�ԇv�}�r��r�cR�O=�љ��}Rn�j���usX{�'51!{�k�0ηuUV&Z�=^B��s]g%�z�^;'�QC��ݤ�+=��3I�WoV�d��;]����ɈV9I�0�'��o��q-��N)9��u�yUWm.��qiC�ˌ=����}���Ć�OXVe��-�3H.�w�P��o���f�	���\a�v���p��N$<�N�����ζ�s7m���ԺV��5 ��u�P�^��LB�/W>���6�d�ć-'��33!�yI�$��g��sEz��N6B�O���s��Γ��
����պAk�ۚ��VWz�T*�Umߡ���}����n��Tn%ۊ� �Ǖ ������T� d@ T[ *��T    @ � ��Sd
�֡YVڥeb�U}*����m�*s*���sm�P���z���W��{�ֳ�-�Sj�&��I��E��]q/uOu�C��Uw��U1W5VʹW"�Rݡ���ϣ�sy�h"��\�Hb�*�  �
������.��7`Hֺ���M���U[V�S#6ޯ'��Xbq�/����=B�-&5 �>�f2w�(n�n�j�z��I׷�Ն&�jb��rO9I�+2�c^N��=�ʪ��c]��-�yΰ(y������fu�`^\a��ɹ��sMHe�x�f[�a�<�7^���E������'HV�s������C ��6$��?c�{e���S��Z��Q��vɸ���"&���ē' Wl��� ��Y���y�� :�&�|������2��ڛ��C ��ҹJ�m}��k��0~z)�=}�㛾�A_1>�]���oס�H�B�X���z� J��VQT5.��m��[�{`�&ܱ��d�m�J�hbD�K��{J�5U���������f푹�;�OZÞ�$��@���犴/Vo5�6�>Ăf;o4#���ύ�ᶽ���x	�5�z	D��e�R�[N���[>.�����Q��]'��b��z���$�\X��*.;��rx�l���k�z���S:�`����bZ�ho��DU��eM�Ei���Zf�{��+��m��53�7�@�&����ڗ'6m����
�*��*��Ul� ��,��i�`J��v��0� q���B��m��C�o.6����p6l�?H�c����+X���M�'���Lt�=�GIs����V���ȓ�.�/� L�0[��6�#�8@�_}su�v�����̿ �ȹߞ�1.�� ��/���,���om��#rᔰ���,��H|h�浽���	�[s�N'�^�C�>BY�m�����YEWP;�U�SmУx���T���������v��ȧK���ZX���$�"t��;�k(*�
��+�2�NⲞ�v���[<^;ʇv��	� IH��4y݉m�4���7�S*�՜���b]j�߱>� I����jX�wՖg_4� ��K�����6�
b2�]LW >�ܶ�ꪪ�2R�M�C�K�-j���Wv6�Ro���Bf�6�v�XUl3�I$�ĉfB������y/�Yj�w��n{ت�����
�ToD���bqꂤI-��ox$�2 ��S�X����1K_@1Ԁ���ow�Ciw��UU[m��j6V� T �J������p��ӭ��1��n�����,�K g��+�?�/�<��&��{��c�	>��~ީ�>"��� W.%D����ް��<�ԩ����XsK])7��V6����ʮ*��aZ��l�o�W�;*e�Ku*h���1)� ����}�f��9�$��r�
���.l�O�uxZ'�a�s\����Fq!/P�T|~]��b��;��!����F �6Y�����g��VV�<�R����9��wd�7m���x�
�Ȫ�ɵޑ�嶷����TAUT��=W�l���V[m�͔
��l@ -�TVUPd U 
�Um�m@@   U @  B��*�1�l�S��@  EP�UU�ml��M�dJs8mm]��V��3SK�Skt+m ,lp��]zn�=��mڎ�|�iӷ���p;�n�\�� U	�������^Wo�W��A���Qݶ|  P *�� <UUlHR!���,&�tKj)�*��69r�Ix���Of��$�`Y7��F����1���'ޅd�ܬ$�:K<����� ��BH<��vfU��t��]���4Pl$�w�x#���UU@�-[Ysl@���t��8.Ky2��aZjC�K���Rlj���
gY������������AU�!Pg%Ix� �s�EL�H7�ؘL�!Li-/�0����� ;̬'���=wp�W:6�
b2j�'��J�g�/3Y� ���khlڻ���   *���
�qY;�`'�os�sυ)]� ;�02�pS⸿U(<���E/��k���R��/s�׳Rv@��O�������^�w�3�=H�HM��[dv��f��~�aoN*�Y2��Ր�BiE��:���K_@1Ԅ�yʴ��	�3��;m~��fDUUF�%�I|T��Ìv����]�6 b~ǻ��INëFӪz�c�� թ ,p�FB�rxJ�m���YA�-tUA�;�ʬbN�.m�����WYhT[1d*�� N�m�6� �������sg���=y�l�R y��U�V�	 ��Q"g��N�W��i^sT��\$�ȟ�n䠦!�%
c�T��{�.[Of�y4��9�� �A3�.�<�ާMH�ϊiϻ��
������#����֮:T�.y�,nF����������o�*���$�H�btK�t�j)#� ��&�g}]q 5ï/
B��Q�ux��� ~�Rs�r�WmQ�FE�fK
q�T�m����٨���N�e�*�
�GO�('{B�H�m��F��1T   �gu�6%MĠ�6���I�j;�G
��*��5�C���#<S����z�V���;V�x��Q�U�,Ԗ�6���� _
��9?	F@ߡ2�ן����֙O,�����
d$|�Ұ,�Y���U@-��g��R��}��@~��۹,)���qr��mȔ���*�~�mપ�"W���/,@��5uQ(�usף�o��v��T��s��l�ղzx��[|qVbJ�%+dpyļ���	�&���e��J^sSʟY$�f ���Nd\���7v��   U �g@�U,���[����ܪ�ZA ��acm#���R�V���B@w���̪
�֕Om�i�/gvڞ�C¿>�[@UP0 *����M�6��a���RQp�	��ʧ�]�m�JYk��{�[Ȣ�-��񱑱���w���uP:{� ��
�9*�E iw|^Sn�(Y[�ڶ�*���1�^
�
��� LN iY��N�Q ?�e�J
!篮��3� @��Z�>�O
��ֿ¯������q��l�	�u�����_�����`��Ql��\�`�Vfu*� V�k�l4���
��� T݋�t�[*��AU]�  �    *��  TP �
�� B�M�7��7Z��m�� �@ �*��T�  *��{-�U��m��nb����1-s�Rݶ�kv�ĕ���GE�m��`� <�;�dw����v�{�es���3�YWZ�;��P  
�K2���ֻYm�vh]�.H:2��R65P��lr�V�������io1M�]��;���%�T���-Jc\�I�`Om" ��v�Ύx�
c֢D���K_@&�����̖� 
�[]
�=y�L ���ʇ�������R����'��ɪl��x�dힶ�l�̶1�"�h]�u�JYk�'�R��U4�X����j�3�eV���"I�E��
6Y>�7���n�I�βӾq�l�1S~�ԣ��غ�tR8�{r�{^�w;���   UPmd��k��VYV�(۵���
�Z�F����sn�잾�.[|��<+��@���&�y�9Y~e�y�ք"ƶ�H�*�mq��C,9۶��Z<�' �.�MsUv���[�<�D0���4;���G8�o4^)W5:��0 9�s��	/��\ 5Uq��'�B֐���j�32 uӂۺ�~�ў�N��'6�}���v�UKq��8��q����W�l�N}`�������Rݮ�M��P�N�oxZ�!�lVA[[�mP�  �F�l 
���nV��Q`�\CeU]�FL��;�@��eV �2s^~)K��l��-�i�`=�h���8 j�e���dg��O���*s��HWPm�,*Ħ��D��*"�C8�	������1g��i �{_������y�J|�x��3y����>�~����g@�n�@����)=i݉r��T�5W`݇$��% �6���z�J�9��*�@nfxەUUV8�rD�%��4	ӽ ''���`�H�p�3%���mI�8l���z 0���n� ��N�[ Zvm[��;ܹ�z�Ruz�V���-���Iq�����j|��}M@1?K�[!iE�,&��*��v� ��U\B�`����G"�4U	b��Kh*����̪�' �d��I��[l�<�m���5�/:([}� >�j>�Q�?@�[G�[(��������+6K������?c�7�ތ���h�D��VN��~��ޜ�l@���:�mRS�3m�`�6I x�p������M�$��΁��R.\=����������TU���0Le�E\Kdm� �  *�UUJ�P*��e��-��V��b�~
� ��˅jBn|���.��@s�9��JF��� KHzG∡s�� ���ڒh�̬
�Tݖ��oc��L�j�t���z�'��lm�GT�L���$g�pY�e7o@�
ۚ�������:�,V=z�ۺ@�e��>UT0-r\���X��J���.�,e:�@m�����H��_�. I>�����ad�pdC}�h�sϰ�8sC@%��ȟ�J��āz�����s�mUdUV%�}ƥ,��j��W߿x  �Z�m*����cv��  �l���[@/TY� � �@ �d*�V�  @ 
�P ����  \���jU ��*m�
ʹ� �@ d� U;D���dcL�Ģ�P#D���*���m��ܝwj¬)-�a6�7c����UJ���6�֤w�\��wn]:�͹�m�VV-�ul���� P ��PJ������on���m���_� �U"ʊ�b×���dg�4���<]���u�P(��Rq{�K�N���UUiҴ��dy����s�I@*	��OX	Ky�:�B�֤�?6*���ŵ&�\@��k��TT�~�;3%��M�e�I���-��3I/��w�*����@@�g�O�'�~.f܎ҋ�Y���uO@���ּ9<ү|�������<�Ķ���t:�n�{��eU���\}f\	�6���ro ���񶻌�Q�w�  �  SmPT�HH �A�I�	0��	I(� 9&Y#a��]�R�Hw�Tm��Gܣ0mt�m\wRUIg���ʯ�	�o�ڟ(�Z�Zrw�(zݩ8��%S�Գ�V�I��U�Cp�"#7}������J�|��$�X�0�����y�s��n�Du+hj����.�T����x����t�zz�*����%�V�e���)����~�wU(w7�*���} s#"$<7y��W�W��T�e�j����&�ն��޻�T}���o��)��ͬ�%WT�պu$���7m"��8��1���L����R,� *��@� ;��U�,��m��cCX�;Rm���I��+nUT��Js9o�;�+���r��L�;j���m�G��C�<7H�bAw�R$�k����Z�L�f��t��-բC�x��=�*��u� V_�j����m=��0���o���Vܤl$UߺW���x�o�����_l�6��0��lwBF�Q�����y�����_��ڽ� "�%�b���T7""&�b��m��$u�~w({$��R��m��2u��o8ao W�[|ij* �&L� �;��Aܓo��K$#vg%9;u�)�����|�����M��sj��=�ȣ�v� ]�W*Ͷ�*�T U@�+�T-��,�^�m��6@�lU T.C*�]�H�段՘�IU$9%S�wW^Q��;���)���9��{��vOY����VF�1"_�*�wou�ɻjx`�}=���{	�~��9}�nz�s���$���UT0nG�`]�c,;�aM��q'*����>%9w�Sr����uR�ϭ��j�8��U /s��B6���N�DHxm�6�r���Jj�fd�
�']�S�r2""�: *�	im�k�jٲUwcyk��ux)�>A�<����2+��\�s$�n���P�I-~�cɐ�Ue�L���-B�[j��m� @��M�]�*���6y��0*��&��5u��7��!ԭ����؎������GN����Y��zN����8���lh�n\�)mY ��C����a��խ���ddD���9�]Y�*J���M�w�wp&��zL��UU����b���dD�u�z��9�*�T�\����MG���ۥ�Fd�	����s~��6]���*���$�J7M���ۨ�s��ub�:���'}�{@�v�;�u��:�z�����'y��|u���hv���'Iǎ�#���q�Ϗ�ؼu�,��ǈ��s�{���T�s+
�7;	��[yˬk�=2{��Ļ��:��Ǐ]Rq8��z��s.����]u�Y9˯1�>=^�i9�N�u���X,�n�_�d��Ƕ#Ψq��MMu�I�~J������ I-?� BV �ߴ�~0?�~��L��#L0�w��p�@�,�g�g H�� �$ '�t�I!�B�x�f�A��za���'&�O��� ���'���o\�s��q>	O����3��&x��L'G�w�i����>q'A��z I?�N������I�I��| $�@��I��}�������}���LD�S�}?�����>�!�~�@I���4�3��!��Y!����_��N�����.��_2}g�g����a��?���>��!�$�P���@Y	!?$����B����~�Nϕ���N�<�����p���>�:/���I���_��x}���������� ����G�� �}�m|'�'���'���~A�}&���}?��>����N���@��������| $�C�?�����g�>��;��!�Έ��! O��� 	'�g���'�y?�?:R����	��<<�C�2C�H�@	&>���ad�ПP$I`�d�%�qe�f�tN��뢟�D?��s<,�� $��~_��'�O� �a���H���P|�?��������?9���%T�-�������� �'�������@I�O����'� I>��}��@��O�ϑ�O�C�p�W2~��C���C����~r��(o�w�� �}�|��Ϝ�|O����|ϲa�	�>�I�?T�'d>�@I��@�s'�����}?a 	'�?hS��᾽O�������'��w��]��BB1���