BZh91AY&SY#שؖ߀`p���2� ����bF������%J�"���5:ε Pj�ю�j�Ȁ�E*)���lK&E]aBv�H �Em����(��a� h}oe4�Z @Hl��� t( :
h�� (�Ҁtv� ����@�9 �7� � P���  �(�գm�Jv�  =�Z�u 
      � �:�   � �N  
�F���� .Ί�(հwv7 m�SGU@����V�HV��
r���n��E���4ꅰ�j3�����wm6��Cmö�]��v�g�� �Z�4�QѺ��ӻ
��Z���Pv�WI�$�DR����0ʄI��F:s�֪k&�clm�j-�)PE�A��b ƭ��
��l��ɶ5�	j
�V�Z5�L���r@��;i�l�Lc[[�!�M�&�URV�̣-�5��`1ӹk4�cm��-��m�KXf�kJ�AF�a�J�"�@��ՙMm��j��j��6Ӷ`;� �� 4*��0�hŁd�)IR�ێ�l����e��JZ�5� Z�-	k(ͦe�m�ݷd�*�%��J��64�w
W*�1��@�wأU�p;�[�ܡ#[5��m[CZ����Re�t7(V�@���X
�g]vD"ژ�i�l������V��������&�*��v�
D"4:4h�lv�镶.�Y]�N�LQ�EU)E�ZYA��ֶ�P�Un��f�l�����fҥV���F,4Xm�E6j�-R*�I�v�jAD*��6����\�6���t��֩���a�jY��52�5�,�wv��m6Sm�`��٭�vq�r�&�VQ�լ���,ʦ�Ct!	��a�F�4.�6R�m�ZWp,γiP`�Y[i��T�H��*ʐ!l�����[�3l�@�[lʅk0-6eMwuȵ1��������Ѫ��4�  ;f��A݂�wg1l�j�]vΓ����6�6(V�Tmu؅�a�uU�V�jի�KM[��ل�7kSl����qu�FD ���� [.�H�h���,ֳ���m lִ�S(�+ERQ�֖3�#��l�-�l�T�t&f�L��V0w����il�7eJ����ُ� �~ ���T0 &    EO�0�U% M    )*h�DɅ=&��CM14ѽF��S�@��PdM d hi���h*oSQ�Hɉ������Hт4= $��&d��� &�~���<�,�!GBY��!JE^�0�V�[^%�c���tr�	B�
D}��=��ڄQ^�UU�DE~ ����0DDV�yb""+���H(����n�_�g�Y|G�'��3 �$�u��w3TJSBU%4�-f`D��*m���~��q��]~��I���p �L�c���Q�IH��T���r�p�(@��m�$$,�!fM�X���6��vmVn���arL371�ӈs���0�ֱس�^Y��d�D�G��ԭ&շ���t�%���OuM]#�Ɲ��n�F��z��Z����v�j��������! �A
���g��Yd@	*캮�w^�M�R�z1���]��� ���U�Q�bd�sj`Y�n�JXQ�p���y;4[�b���eUaH'Wn=�j%$��J�̋u#1�j˘�nd��6(�@݈7t�lge��
ۺm�$�e��zf��N���{�TD)! D2��B@��Cq\�^����b 1��1���wGʻ���{��]H8�i�r��.�ɲM9�i�9�&m��XJ�������.�Њ�8�ay�YZn�u4�dZ���/U�������sH�����4K`�{�.�n�3��ǫ��=�ْٞD섗s���y�n�Wu6[��Y����\��:x�k6�$͞�i�W11Bbq�{Zu FC pGN�p~e�����h[4�!,�wQ�ݱP1u	��'B�'m�Y�p�,X�t۹W�ȝFY�2QU*7K�7�?fS;�]��P��e
�H��!B�$ �!!�h��B��#��	Q�N 6�B��Ir�ۧ&Q}}{��W3&̲ę	��泧vѽ$�d,oe��ն��*7E�uvc�l��E�t����39LX��oYIWf��Dˣ+Y׻5v�� i66Tr��T�f���n�rF�Z�� ��'/����h��V�Жʵ�xr(���V��+M�Ρ�����b&n��u=&��%಄3&��Ibv���0PZUee�M�3
�Qtq5n2�Q�
圾�Յm��2D�f]ec���-�j��J���Y�*8�9Yf"��Ne%G5��+��m�nT�L��f��[k4c۳-�[܍�5w����f�M�O��Ru�̘���ɋ6k
�elי�J�m2�Z�4[�=d�1�p��ј
�q4���˧b
�N^���,9�b�k���zo�"Y<<�SY�x��L��:�S����ԈS���@A�h��Fbvݫ��]��ɱ]��^Kn��Y��ͬJ��ε/7F;u�u2�
 ;Efhe�EHN�N�k�ӷ�X���*)Vh��0a�lމksF�Z]]����9$��ձn��K^�jL��X6�Cc�oN�=�)KܷZ�nhYX��Ŗ��I\ֺ�����f�_:6�m�LD�
�6�����A�G%�(��ͫ��.�Gfuv-GS�ɬ���.��u�21;�ou��:*�e=�F��`D,*���#M�*N�Ǽf2��k�{����w5���rY���oa�F��n�M�ʶZ��z7Qt�ʼ��jE[Y�ĝoK5W)��.!*���ʎ�%�BTD)!.,I���G8�G�[��;�R���7	܇������)�H4��
�J"2X�Cչ�\��Ɩ��S�?l����f��K�mb.��Ĳ�%X�y{�TJ1�T����u!a)Aj��	 ��-�o-^����+u&J��&)��
:h�}}��n�-:w����ܹ���ӯ�i^E��7�+ls*n�q�V�J��B���.�/��v��Z�d��:u}�8��s[��v�I<�]UV8��x2u�#������S��j�ɕ�����J��	�M���;@i����ua���)�C8�O^��&��&����J+FD;f�F`��wU�3UK����e�x�j)��	��6em����,~1c���9/1A6���]i��a�ԡ���vc��w�M
w�,��m���.�VAqV��v����]Se]ū+(�� ;�������w�/�1�GI����o�ҝ(L#�ifT¼.����ͨ-�1�
��U�,8�TYY��+ov�;�����YB̎�����ٗ��%Z�� ʲ �ӇD�¥C46�
�H���*�)�ꭱ`�W�?�l'j�&��ZX_��sr^��W,�|j���|M&
��S'���˼/2��I�ɹ�9���-6q���k�񓕢�6ӷ8_]^�-OXo�+.Î�髰Y��a�-��b�kb��A\����gE�c�����ʜ��S;;�YUΧ�H��joLq�@!�!$�!Cl1�!�SFNKKT���2BP!	H�1B`�IbL�Ę��C	�HDwI9}%v�W;��u��i����+`�+[���/!��;�	�4P��&h�F�d�� u��c³j�藱b��M���h�C5�,R��Q�+ZOvRyo1�Y9eFIwe#Si([��$��K&j�v��D茋U������h�.NP�h�%�+	�rڹ��̒fi�t�f�6Q�Q�]�R��t�p�b�A٧f`�-�v��lCR�V�%�f�y�R҆�3 ����� �/K�ZxE��R�Mڥ]gutق�6�x^J̚��lX�'E�mݵwr���C���\�jeq����ft��j\�UV�.�BI��Jm7f����T���Lۂ��j�I9382����5��4�l�a7�`���W����jK���z�XԷ�%�
�H�g�t�7&��Z0�����0���l����d����4*{#�{����3�uu�e��U;oS�<fY�y+��r�wZ3\җNs/iNai��B��i�b��"F��b����6"m�W�[/0�A��c갲��Ԅ��#�T.~E���6�U�9��dJ�x��Yz(�[��/0[8�̱�0-�
����!	"��Y�75@�bW�SS]�r�D[*be�W��-�7p��m�V�Da%�הl:o-
˭�'Gp�t켬+����ə�&Tes(�xf�,ki�u���h�)��xpU�S�Iv��5?�ޚx��[Ai%�Tg[f�e�n���T-�W�䞤o4�;҉T�����G�զә��{�����e>uZV�:�]ܕˑ|��5��7�n���A\�]N�S4طr�d��*���9����X�Qi:V���͕�n ��JP�&1%�%�JN�K6�w,��ɻy�e`�Q
�Y	H����5�u,�	���A6E��v�E��-����t�zRbVn-6�;3�
�p�����2�g-^*�'Ky��V-�^
R�U�3Lt�)��`&f�;G���]�hSfa�{nː��J��v+)vq4��j����;J׵"��u�nayp��,[ʴ�s.R��*�69Y��e#i����cR1X�
�T�oN�LVB�B\D�ۄ�)"

�)����6�8�����-hBƙ	����B�(LP��B�.$�B�i)���+UU3:����%GUvٛ���� а�6�v�(vU`A�4��ֈupJS���w#z+s�[�3/ynX�`��
��	1D4!Y��*�I�M���f�gPf��x�8�Ƥ�*����Sd��LG0nK�0mS�f�H��̺R���ok4�����Q���1���r0�њE�Z�2��7A��˻���*P�	Y�� �����J��$��R,�+r<wk�5$��ݭ��dJ4k����1��h��sPY�a�/i��؉�m�MR�ٖUn˛�K^�K��s��uJ�+�)��M����+�&�^RӴ5������e��أ)���Z���[;r��X6)���+d)E@�\^:*������P�G*�Ř�<�E�>���}�uY6X@�S�dһX�m�+V����x�J��sF޲u�T2�82����f[���YeJіt��j=�7��)��xn���B�r�%�0�ݞ\�so�ы9Xg*����}���
�.z���b�ܸ�ǙX�ڠ�B;�/+,h�թ�����"��-�%]"1IR��5Paa9��A�-<�K�+"[�P�db�I���he^]�j�X��ejY�0��Jˌ�%�o���^d���˩�V9�eѮWb�y�\���oVӽ�Wk̵4#�b]��n7eUeݘ#Bv� ��T�d�� ���"�8�Iux.V��`�����k-��6���f�wE,&��7`�q7P�R�]arѲ$��լ���+F���4�3�\�/;�AOVn��Jѱ���֦^�)��Al��7Mb�.^^�ˇt�"Q(&n�H@a�MH%��*�B�P�0e*�A�V�H�s��s�9x7Z�Y�}q��i������7$,��P��r�+.�#��oH;�̖�����xÒM5e=�+)8�t$��Q� /v�.�Y��uJ�r��J!$
"2V�F�(!Ԡd%!K$D!@�B�W�Xr���5p��"G��+h����L������R�2�(����&-z�Z��\��G���m�+7�ì]8�4��U�;æZol� ����X)E\]��I��[�e��<�]b�;����VK��z��*���zh�yS���D�3";"F�Z�v�����)��3j��ŻY�.��j�2�Ct�{��B�ʣ1u:������4R��3��ٌ!,i&��$B)U껪��4��!�Ȇ��)�o7�X7�8D5���p���-�2U�M[۷��l�˴�awB	�!U/dX�����c�uWr��]2nЉ������Id�Ιuw�3�����cg)��E�OV��vg.����Y3t�
۹i<�6���q�y.͒��F��2�Z�y5��a6��d,�V[����t��ڍ���z�e��,��$�+2��U�7Cn��R��;ˬ��)չmroE����Z�U2�c��ʕ;�,����� ��c�B��֤�u���4r�62���.�:��~��ܶ��i �-F�	���Z��n9X,��:��^8�䖝���-�:@h;.�6wpK���\��H�v�)���[�a�r��ʍ��sY��.��X����)��p�FR��CU'? t���/&iK��g.�dS�	�t(ێ�@��Q&[�����Lb�t�ǍȎ
�j��Q�eܫr𽙗M�åmy�)b8�1p�"<)N���R9�ZU����4j�&��&���zƤ�h�OoY{y�^�+2Qܼ�de�.s��1p�Ҥ_>��.���{N�P�h�:�6�f�m���d��GuM��cT�[j��ڕ�m��n�J�pm�Yr3�3?LU�Ar\��s!�r�&�Aӽ���F\�R�+�-��[v����2k��z��������$_	2��eڨÛ�4��5w�S� %��R�[�nsm`,��[56����ݎɭع:$�<�]�uf�έ"��/6�UK�dC�v+QV�oFI�-��a����.�]�Ս[� ]Q,M��)c)bA♺8�����c��N�Y�eI"V(�"A�*�9�W�o�s	WQD)](Y���Y�W3��%M<��|d쓜��Ɗދb�7r���y�s�y���B�W*��&1�4[���%\n�N�,7�b[$����<_��K�E;�\`ܵ0����e^�U6�aB��҇������B�����G4�2��td{�Y�=ӎ�� �D��l��'LCF�/YM�3cn�քM����̽B�hʝ�2���ju��t5h�$XsV2�*P���SR�8wPt� p̵� �W��B+i���2��#�$\N���p`�E8$�l�r/(�D*�\® ���D-�]u��*�4�5/q�Z֩��X��w�by*�V��t`cMu5ڭu�+obV�eqbowfX�t��SI�vU�uvr���n�z�@�sA��Q���W��.MX��{gEj�r�4�+p@P�W�S��K6��}:��<�t�k�[�ە��;!O�14r�2.�n�j�،����5��TQ�5]W��.�Rq�8�,����A	F^�1+s]�v�ܰ��Y	�C��,NIb2�W���$Ʈ�]�oHW
ٺȌ�&f�I{B�mh%��E.�n�k��YY��jV�4BH���(M�)��0�j@9
�Y%2�Vmlf:Pę��krZ��K�{[�T$�fg�8�p�O�0(:���4���_}9%Mo��ۃvQ� ���h��Y���i�1�i{]S�¨�q�����T;3SW�����W�ג�lTsp���R�?�1╶�	��DV1d5�<1���+F�z,��,��Ȓ��M��VU�Ԍ�e�(��ۗ_���.@���x����d��SG�tّ��"�3MU�&�R���� R���3�L�3o���-�]G�,�z��{��,�a�����;)�)�n�-.�]ѕ'=n���ow����^{5Y�9�͊x�f���zZ�t;%	�n��±d�ȯ[�ཽ�dQ�]�Q&N٦��r��Y�3�����I�,M�p�G8q�N�8,��2�}� �Ie��Ѝ������v��V�p[s �ނ��]WS"G����G4�v֫�3/B��]+�+�,_N7�ŢFXޠ�+L����6BY�v��ڑ1j�;��y��e�Go�gL��E��&�Z²r�j��+j_�^��&'��!��:��o&���+FF�A�ΌGk��Y�`��ͼp�Y9���+]���w�+,bth,���`��%oWI̜���)�`EM7��$D�ɵ_(ְ��m�S1���h�J�v�f�W}�[�6U��Ԕ�ٗ� ���(�1�E���2�e�+���`�;�٩��z���Yw�33�&��t��X&q�Y�]�zِS��1�~��f�u�i�Ƶ)�3	J�g2䘳-���劇���맴NӍ
���Ty���X��������]\�e̵<-�MU��Ҏ0���R�;y)ț}��3���m�v�,�[�d`��.^"2����ĥ�.O-��j�Υ�co���8���/h�P��Z����+�d�rm�x�E��˝�2�v^��P�'j�V����'�*���;�DT����PS�=`���H,�z�3EӴ.u
X2���P�6�'*D+)�{�3��N�z���k�"S�ݰ�<�0��V+)d�(����j[�o-Q�8��-Uɕ���2c*�q�XR	k4�]9{�$��l�A��-w)u�Z=��+!��:Q��M��&Է�p>�C�����ã���(��<5]3���'p��H�+����9��`�LlJWei*-���/K�%ދ�� ^fΰ��DjV����Jp\d[����z��uj�&lR���f�!:�e�җ�ca޽��_oMp@�1����$��]ӯ�a1[���������u��Dy{q����	}����ɪY��c�$K��8�<	�\#�Q}Ո�W/%��53�������[}��ra�W\��4�.#"ѻx�|�r���r֢U3e���1'�ƪ�J�Nl�*�MT9Ի��������Ew;
tai[�h�/<~5{�&r�]3�QR�qƱ�B�E�W&v^��C)E;e����HʊSp~���]�]М
j�t�r�Zr!����j�f<=R��<yq��n)\�����%[��ӄ�|�%�gQ�1���8r���eNy�a�� �@�¹ǋ�ɑ4C/n����V����M�J�o��W����`��4M��t�6+f՛��}�9�@��G-�6o;��Z{�Z�ۍ:Xwy���i�S������ujG*ӥYy
���D�hᙵ�c���<�׵���:Dڶ/�.n��E�K9uF��]-�ޛ(�P��h桢��>Gnn�.���ȕ���(�����s������$�b�E�*�F�����6V�m�H���6+W�3��4����U�;�7�;�/3L}�M�WA�4�����(V��x9��Ƃ����[��d7[]s�U�F�0q�B�.tv+mw�)���	�ԋ�g4�<�Wu�sJ�M�Ѻ�,J�����������}C%�������n�N��m��luAs�Y��v��<��\��������:�ф�\������{ztF��cniD��V�M�6^_U�2���M|1B�a���, 
����>+k+.���)���J��wmZ���e�����?�˔3s�$��Tyix��9���������I#�8̎ȲQY6�e����բ��L-��jT`���
��r��"��V�r�a�T�l�R�G��7[:��ݹ���P��iO,���/N��;����ˣ�q����uvngP�Ӷ�
6x�5u�6�M�ujo7�<�7i� �p�ES�B�L�!�}{Yc �19.��ດ����e��K�2�Ġ�X{�r�~ٽ"�I��J�#��G�o-�gt��|z�����\��=�x1�8�԰*��er�W���'-
�i�/?e��6g�.��� c�-�*]��V.+���d�,���g)wS3��O6�S��6�=ޱ���1����ڽ<��k�����Y =2/E(��w!QRД�R#t�V��������z��Vm"F�]\Op4��3:�*���S�A�$�s5�p�M�.�,{���M��[ѱ�0dK�X��G�c5�Z�* �>�"u܁���|�����s��o:�ƦbV���{y�3p�ej%ɇ+h��kR�3*�&l��'^�Q
r��z]�Y꛳�L���-�q̀So����p]d��̵E�+ǖ���q��w�ˡ�z,A�VԔ�-{��fe	08��R�<2R̬��I���X��3�X�mM��	�Nr���!:Q[uwSXL-��N̬��xٝ��dޮV��D�S����lo���*�#���j��z��^N�J��U0�^�3Gn�Ό��v�3A�p��X�Y�8��D
�L��g�W���=�$�:��Rͨw*�Xi'*N"�&��%Ixd}Z&j�/�m�gW%�*ƻ���)D��ܚ�ހ��uL �cx���5�PZ���ǽ�*��k�_�7{C�B�KN#zp��嵻3X�}l��6+:�qX��`T+� �$����h�4�l\�߀5��,$b,�U4��W]sa,B����s=�1��[Ҕ�3V8hgd��g2�;�w�eLB��gf
�7�]�˶�1�j�t_ %]lŸr�em����͔Ɂ�1��w	���m�0p�̀(�F�I�~u��7�[��v� �w{��z짃��Tx�&�H�E0�Q]]�eo��2h�&�ڶ�ųq_b��9��
�yw�S5�Ж�D^F%v�Pjݤ�p� ��˛S��oRz!%�t�6��$�q�N����m�Q���\��sW]]�׃YJ�y(SD�n]��ԳQ(��
��� �Z(G���]汜�tu?l�q�����C�e�lU�m��/ájQ�uk���LL���L�A�e���ΎU�777qj|�HjN^���Z��"����)Ǘ:Cx���"d��[��<�,��I��&z���?e�N�7���}PdT+B�q��fP��d'FV�Yn�����(Vv��\!�M�O���h�z3+UL��~��\c���^eu�\��H����圳4s��b�gt�`�S��[U��N4⨜����vͬڗ�q��
�25:�˽f����Jc"]Hթ�*��jh�r{�չo����F�\w+1�T�u�6�Z���-#k��׺=�U��i1ʚڷ��*b�E_X�jP}���2�U@zfX-Pl�g/��W��U����Tc�Y��<�w����x�i�(jԎ%6w�.�aO{k7M���N���[j�������-ݗӾ'7�R��l˕�.���:��#[�&~�nث瀽�x[|�b*}�m)2<��⃓yY�̫�����ʧ-OF�њ�fV �-�+v�P�.oƹ�ڗ�ԇ:�TjjBwVb;�]���Xt\���.�g%��I���p۩���\���]���W<єT6)7.p���ީ�Y3��Ut�ݽ&�Qc7:j����Xi���Zٸ�}���t�f2�z�כI��u���ų]2ll�.~٬(@�ݛ�m��[:�����)�T�����S9f��L5Վ�N�<o�f�6�����S��V��Q��\���R�ٸ�I��'_*ܬ���^Y*�U�w�W�uEp����M�8������u�d�ϔ/2�����S��q�a�ʡ�`���A���V���>�V�F���+�]i�Ճ��;˺�g���j�7j��hL�ݏV�h�,L�������\�g]Բn Ym��pɓ�E�]iaV$�z[U՝�e���4jX�/q$��0�8%�-7:eh�����w����֋Ѵu<Γ�
�'h��N�u+�⎞�E����c����g������}$��p�ǒ�T�_�ڍ�ƆeY�2�T�u �w���ã�/�������3?3Fe��h�0e4$ځ����p��Y��/\6au��ewt9ܐ�7)֮8��ƻq�l�Z���3#S�v���En4�'(L��.�J�qm,�{����/7����1"8����,~�㼹�9�XGB�Y�LM7}jD=�c��y��L�)��HMb~�V�v�*2��[-i�t����I_u# |��y��v�j[�+�t]�4�7�-����Q�[�}G����$�̣tm�y�]�)nV1ONŪd�QUw�b�%�Q��0���;G9QTC�7'5w��S��J�����@v`$��WPRM�@���6��nj��	Ӱ��^�%V�k�d���o*M���#��oT�э����]9���f[�D�NT�=��do]^*{���%H�	��T�x.u��0�;�����Or���7y%%�re<\������yk�V#�4CG;k���p��s��$��/Wv��:f5�鷻��E(���:�ɚb�7�]���2��h���}�����=�a��0�ޙS2�s|�I=;]��`/v�Xq�kZ=����;A�N�k{�҂CT�z����;����b�rS�W\�V�z33�r�%�ζ��3�le�]wBRtã�㧍n���;r��,(B�G9�֮��$����C7�9��� �8�Hͥ��Z�u]������R.GkY8kT��hd{�H��2rz7Tꭑ�N���CTS�ՓU�@�j�s��u�S�d�y��b��	���;^��Ί �j2}��g�m�S��g�Z�<�[�5h�F+x�w������f�K�ac���v��8��][��M�ɸ���y�Q]ꣽ�Pfh6�	��%ci�s�����P��9�����ӘQ�[1�͔qebo:��-�����+-�ǋH��V�ά\��N�-��#?5��|:��t�RI�;�U���D�3��=un��E�fE�8�����Eͻ9Ϭ�ۜ3��f̉�vغ�f�뫒��3k�e>0
8�G�a�e��ȧl�z��u��٦{a��tG�7��NC8]���Ԫ��*�<釨b��i��3�d嫞ݙ�V���W��j��Y�u�A��M�s����v���QX�B,V텛Q�yu8d�ɓb�l]F�8���vwOu���F���
4yb�;��7�[6��o�M�Tc�wm�v��e^r�U┴FK�����{���=�9��(��2��!�rl��v2�u+�N��@�<���Q˫�����?��iW�V;Œ�,�C� Qu��+;sP�ܞ .��Bޫ�������s�|�Y�Y|d����=S𑗸�W��+x�@�[;8飥�-κ��u6�_�I�yT�b��p,A�����®�62�WX��j�+K�a��V5�s���k��T�a0'���D������	у1���xFn2���D!��R����۾qu�$�>�:ٰ-�Jv�m�9O���FfT�(Y����[B-ʻۜcmӼ�p|:�lP�{6ƽq���U�ő��ϼ���s%��4��\���q��Q�5����ahG�y�ft��m����y?(nB��W���fvl��.a�w&��Cl5հ���r`9{�w8Wxa;:fU͊.f��[��Ty�eh=��5�Z�	W;M���՗
ZΗ��'�Q�u�yug���)�t��Z6cwk���+��nL��Ɠ���F�l^v๔���t9���)�}�X��!�M�m�
��騖IQ"�����#ݓc��eA���� [7_>���`rƝ���[���,��oq����X�H�*�&�F���Y@W�e��"�5��p��p
��.TХA�#Y��yAdR�9�zh����m�9�#��7�Z�$�f&�5Xbf��B� �"������N��8�M�#sgvը_NI�s�֙�	�]�X?�	S&��a)�Lr���8����ԛ��v��Z��J��Of`Ժh�U�{�\.qq/��=9b��Aw��<�c/.�2�P_c�=��0K';�7zBx=A�@�<���I։L#�B�r����ؔ&�������X&5��9S;k�����u�r47n��+R�13Kd�+)@`@(/b��a�z�� R�^��G%�oΆ�T�S�N�:�5�	j��ջ��-@����2f��O;9���vH�Z|�$2���I9J�f�f���ٳ�pVG�3SM:���*�|3��s�n֍���D�Ȧ`�)Fa����Q��mA���*+*_U�9����s�ob �fV�\���ݑ�3����4�L�X`���ᴺ�g8�E}Y��8�1*��a�k6�F�p��S@��}|4p�\��S�v�k5*Izfp�0ݼv�8������@hՆ�f�ֻ��9e�L��Ԇr�Ī�y�rk��m �!�K;��V��st��7D������j�{V��m^��9�R�u�����.`ū��҆n�8K|�M�;�m���8�|�M�VW�=�Cp���]�TTn\���3i���ٺ��Jю��]t���o����k��DB0n���~�©n=�rI:_u�'e3�+32ó�wg���FX�YiM��t-\���O,g7W���%x%ߺ�-��H[Y\�����0���ɳ�9���rS���.�}����Ѽ�]r�;#Mu���YD�9��?9����݅]z�x�͇:�ڽú��{���p,'����U��i����'E���ۅ6%�h��AH:�4U��D+(^�+x�H��kR�1>(�Vl���fEӤ8�O7g6�v�����(/1�Pi�u�b�f-�^kI^��k�6q��fa�R��D(P�W�ǿJ*"+�� Ҋ
�����T�TC�
 �=޷�� �7"��*{e^$D2�@9�Cp*w
�@<H d�@	��U� �J� &J9"/P�� 
R �/�kX��!��!��A8�L�<���;��r(����
���S�z�hC��T5*ws�M@w"d��(B�!��G�C S���"�����D�y�y(�X�*��3�G�e7ܻ�PP�B�(��T�(�A����M񊚞�� А(A	;j	e������H����y �P�└���0^<�\�r��X��5)�RQ�����x�p�@.@�'r�B��3x>@��O!��0@�P��x)�x��s�@�{��E��nD:��M��=�<�'Rd���.O��P�@n�ԉ��J���; �uI��P�*yu ���B�8���G�qrrP�W}`/p)Ġn 2D� � M�+��A�8�P	@�� B�';�$�L�܇RK�%�J��� ��Ӆ�25	��%b: N����\�{�P��y�$sև!7)@�9�ΰ:��:���Ru�S%]@����x�h����)�$z��u�^%ԁJI�|�!̇Pn@:���>f��':�7(���j���Լ½I�fJd��ԣ�C�2�%n����X��7�Jy�jD�@2;� �.+󄨊mB[�(�4�I^�b\B�H�Iۄ��­q
�"!Z�8�M�;�7 nr��j@��SP�#�]��du)�^�$8��b�C���h������Ժ�u��@�p���;�����<ț��`.����T�^�7�C�� ��#!3<�3̇�q�@��Y�A	%�BRB�E�&(Wm,!,?5
q��-#-�
D��ģHS���P�/�s&����S�P�����*!Kp��r�I^4��Kp�DD���BZ%׽J��ov��y�u�d�f*wǘ�(�E���	p���I	h���*�U
 ����ǐ�&@R�r/2BR��)S
� <����!��i	i�$�P���LQDF�ʑ,[P����p���"i�b�F
0�4�B@�V%��B�0Q�Id%"RFd(���`���h�Q�r�4�e4�P�>ii.�F
�[J-
I��$\ �D�nt���bb@yL�D�	C	ܹ�&�A2D�����J�<,��7\!&B�um �4�0A$)(�K�(�E�6�O4ĕ-j$�TBʩ��B�(�R-L����z*,
��"0P���J���-T�%bTC!M8�l�!Ta<��H�H�P����vT�&(�Do5$`�U�#q��`���ҕsI���i��{j��֊�ǅ�����p�dȕ
=#�dX�+$�	5�	iJvb)%"����q@a)О>!'U1g�$Gc^��k�8g�L���h��s)W��E	�\��ɩeVV����V��~�m���P��-5ۙay7BY���^	ގ����zmN����>o-�+�&Y��[�>6}1��+9\��i_=�fr�6�&6ݪ�N��LJ��Onǥ��ӄ���{3
�S�sj��M,ɹ^�S�H�s�@Y/1gRڙ��uuX��=ڶ�	8`�0��!X��&�Hk�m2���P3�2��gIj�K��׵�Q(�w��&��#V��^�M�́!��X�:\��<˼��&����Y����J�:�#�W.t��vMoK�&�]]�
���ۀ*`)7�+9_@�bT�kUnV����4�]�x�d�ح�kzHq��&�4�����e�W�c#.o��x旗k-	b~����-9@ki��R����F5��z��W��J����(�K�Uv�h���k�ū�	΂
���W���o6,�J�\r~���(�ɦ���Q�:��#�i��PT��>J��a����m����6t�J��[Σ���YX��sV�d���j^$��Ss7�7eC�S�������R�;��3E~������r�`P��[��0�	�pf�6T��HBR*��d�ܕz����E5�9�{���:ݺ����Rt9Z��^�QۦfmeM�\�
�:�g"Ď�UD�`�X�aݭӜ�^�a>[|��	e+��X���m\KI]7�%L]���e)��E����&1�������ev'/2гy)��m��-&ЬI F�z#^�3Gtmֺ��@%&
M˭)�c[h�5jm�)�!��k�T�B��T���'��֧b��ʊd��a���S��̥���T�uV�VI�pRJ�f,�z���˖ڛ�xQ�^���8mR�W���.��@��5YD��+�e�^�m�ڪX�yj��X�eZ�T/�8 o�����T��Yُdp8���h���_��PDE~N_���_�}ϗ���k߬����Q>����ms��0��(]`ν�'��U��V&ԡ@K�G]�r�T���V�Y)�]����o#u�k?^A\(�}�2g*� 'C�.ː:�j������+��.^�xa��w,em�武��h�7�(H	�͜v�t�[eJژ��f�Ε��r�&ѱ���t�Y���[��Q_' ���I[(�v�ڝ?���x{�+:����Bլ{:��|li[M��f�*x���k���z��CM��ڑ�j��]�FY��ŪP�p�ø�鬑�f����e�|:F�[���Z[�����[��;
1�{q�+�k���.��H�ҊyY��������]�6J��J��[����)��D���������Mb��2*�9�����Y�a��N���eB�[[6��/zE+a�痃U�Hs����B�WC��V�:���*_T�uCP��䘳���[W�*ɵ�/�rU�2xq��TM���q�+/hؾ�b��^���$瘶��s�$Rj?����H��BF��k�S,��	�k)��8mͲ0��^��8E�E,'��$g��gX��V�]%�f�Ҭǡ>@dr���3y[yF�R�ɫ2�f�[�c_�D����4�m�|����P� �<r�~��;
�1�u-r�W��*�Y�z�X!����ea�t��:�����/;�#�c��rǮ��&��$.��-�Ź2�E��7U�i巴�cN�\ϯ,�(��Q�j����������1ܣ9��Ձ�֪mҧ����x���^�v�31�O�,@Nb��R��5��GN��,����^�|zn���tu����\�<״PG��7����P�AN���z�ܠ��r�ܨj���k�:�#܀����W�0T�_$W����8�9� �Q���N�P��[�������_�Gt����� �&��bh
�����$!���)��z���(�@! �8jƐ� @ @   �B 8`	  ��T¨A�i�I 
C�! "$L�4>��P�B! �PB"   B!Zaxh�i�@	H�8D @$$@� � �B���@!�@�
z=���؀@�A D$^"��:0Ɔ
�Z��� !�  B@eJQ(��! � �p$ D AM�B!@���� I�	��B�� @�""  H@B�&a �	
  ��/! H �H�4��2y�
}�~N�;w����l�fW���@�� �B@$ ����̈́ ���$�B  B  IG�2q50�$ !!@ �4 ��$ Dsj+���!!	 B@� &؀��0@�� �!  D`� @�D��T�bP�
B@�" ���S"� �1@		_�!�h !͡		Am®��f��#  B  7 ��q[֘��BM�!@;e���}��.�h}�g����O� $ 	 �cU-
��(�HD'�p @� �ڑH�$$$@ D#��A�p���_� �� 9�#콥`B$+ @�"YҪ! �n�i� �#F�7�1BA.q"#�#��ڡ2G	  Am)$H\'B��� B>�J@�g���p�ͦ��H ![�}�y�NmνN�f��O���]�� A6�B��� O)�T B�! @&&��$��G�KE��@B��#>�T��!/Iӂ��BA���a0���!�"�pJ��`�  �m� zS� AÄ@   D�z��!\&46�`�_6|C H�����[h�UW����uW�r�1OɈE��pĈ@	�̺�h��0D@�j��X�@��́�J`�4�m �|0^���K`��SM ���!���I��KbC�� A͈��j�m��>j�n��d �#Zh��l�� #�7L�M ��_=�s��Ww�]8���(@�@ �pЀP6�a�� H�&n�4@#�& HH7ޕ@� �K�`_{�T0@�B�g�P�[�D��#�<����*ъH��~Ɋ)�i" �+ꆈ"Ę���ߗe���Zh �0 ��XKf��B}7��ygQ��@� G, 7���1+n��1&W>� �Dg�5ְJ����O�iL����@��� !�%/K���@�yyL�b@ �	��@��+��� V;�œ�+�݁���=�p|z���M!_	��Ċ}=v��+ �G���Ђ �@AcP|CP�A�e��B�m�-8[:ib B������j�uJ���HDw0���`ԉ�@D���L�,��J��p�EW�΢����W�ga}x���ǎ!��f���3=2C/�J  K�G����q�d4@  H��D�!��d�=nF� ��#*b SKi����J�!�
\&t��|&|�+�]v@�E("b0M�b��+m�G;Um�m*!e�	[�5�Z���q��P��i푣 �����2�����HgN���7���)�T+�0����wq���$<���!Ȍ���	�~^J���0̰On������'�/�1[U®�eZ�#n��ϲ�{>�V&A�rG=��
�	�&�L�j�@! '������>��[6�B�Of��,M1�o)���!�t� �\�x"R�c\\�B�'ys��� �U�(��5Y}T}��_/}FSA0��p�vҤ$�8b$_z��qL@/�Б�0>y�#�Cf�)!��<1F��E:�L&@A�<�� ,�dGK��[<�d! D �l���
u�%H@���=峟}/����k��}�P��(L��:�4p&� �1��}S !
��(b�Z�HJl��`"4��*���5�4@�Z=iy�s�� �:�D��j?�x9ߥ`��R�@����V��|��c�t�^���^T]4�D�4K�Ty�����V�����Z�!d�+.A��Hn��ԥ��X�_ӓ�@ �F�q+�d�8[dJ�p�&y���}+j�~����J�~:p~�	G!��#g�L�#F �)������&SK�`���J��'6AՎ��@��7=[5�JX4�8��VZ����@��5^��|ՊE��ub��E��M� �s�_9�Uk-�tO�z�n�0��b��EC5���1���Á��_Jp��S�Wb=���W��^�� Ɠ�ɅED I�=8*Bo�iZ4y�=�H �_Ā��ݕ��s���U�<�3fe ����#D@"4�z�K>��-MG���4v�q�&��_���r� �����<�^8<�A�Z1�� +�B��ғ��L�C!���1�JK���=k'՛���>�Uy��&��4��JR�Lم��9��b�m�1q}\%BX!H�e�|2Y�^� 6�D�Z+����jo�+_6,mH�R<�!X���b؅k2o�W������2n�z���� B��A	��D�g��L@τ�{
�8_K����!B3�ۢ�1H%�l�)` �����}Ҥ;��]5�4H V�E�gս~��GW�����z�k����">p���4#�	�>i|��% @��8)�f"������`/6��� �
<����[LH<;�Z�D|;v)O�U�{WΖ@�K�T��x�iM/��n�muuw��B����HU�n6�"Y}����F���#�Nq:֓�-H�3gK�(��zT�*���,�7�H�uEb�*�v�g��ΤX�p�r����*L���к;[CX��_*Y�����?m ���C��:�\�h�nd�{8��;�=LB7�j�$@�A�2�H�/��X�_5b"7,Ad7=4@-	��S� ϚRͽ���E�D5�8�5uĄR��~�wbX�4f��W��}��ozr=(�!G�_:�L�"�
[(�����ϯ׊ʙ'�9�����R���v�8�����J�������H�����
ke��{{uo��fv��c�^�n;����L{�W�zA��S�ԟ�N~���Eԩ�!� `�������C��˔" @K�]�>lbS);��J�M�N�Wėl�$_5]x)些��}�<��S,A6�B�Z4P�g\�)��*�pЃ�Z���T�i�tQ_>!?�A���oJ���2�1�WUE녈Dxњ�K��}�f�7n�A�B$̤Ȓ|��#�@�Zk� /��7�!�]��9!����_]PH���f�|�/���ガ.x�`����}�����?��'ٗ�Ьa�6U�	=��������Q�PB�%���!$��F	3˽:+�`"h~+Gm�����OJy�n�S���O�A�v�U��O�ABNΫm��@%���mX�\��d ��g}�HB �Ғ��3�]F�]G��[5ʕ\8��1��@	Bڽ;w�	j1���T�j�ʟ��\z=�ȋk��^l-�6+#��y�.�MJX��ϑ���5t�j�rf�բD�����'35����:��lp�~�KXa[���[�/�E_ت�_9��N4L�$��*���R��u,���[�N���"� ���Myʴ�m V�{:�<�e�n�����R�&:k����%O���S�HB����&�;m-U�T�|�'�L�Rn>#1�,�)}-y�8�|E�~,��,�ֽ�{#+�U��s������c�Ѧ�+�08ν��V�۱�L�w S;��.�,��Z�Z�*�frJNV9���-a��6���f+���*���Z8S������H3��N�.���;��㵍��Y�eY��� ]��<�tG x_�5)=���S�:]ٚ?��I�N�4�fOe=�dK��,3!m�̫�p����g�{:���$P�<|TW�(Ut�Ղ#G	Uo��Z�dv��v�|�������ʩK�4�q�emE/C�4�%U=W7A��_�?�9��ʹ�fW��.\�{��a�ͮ���]�B�y�/���djP���ܑ�ڡ��`(��#b�����\�H�͘��_���K)45.�bRҶ��
}�^,�Orj�dd�/���Z��eGv�z(t���r���U�6����ŵ[��c ��U AM���s �}��U��{�P���\%���$\���VH�l��ʿ��4��	�;,nhT9H������=��_8��&|ӻ߭X�5�����Q�NB�*Y�X�1�Ĳ)	�
�hD��'T2F�G=O՞ϯ��k�J��u}��6�YK�J�]�m6�M
����bPs[�=+j������5f=��^Sg�r%���%�C�^'.�7O�ꝼ��õ�}~%}�(}��B����_m;#��F����sV��1��@M����쩙�\L��!
�h���g�!�U�+������1�>����L�^�ڇ��\��u"j\?}T�B ���M
EZ�J����h� ��s^�d�E���=mtQ�j�5YC6�z�ǯ��$d�޹�Ks�EuT_��'�/L�,���
��R���E�,�c�aq��ß�N�t��B LR����fw���~���;��F
�-Y]Ց�m��U� ����->��N�4$��z�  ת�(@n�+*{�.:\t@,y�*� ��U�ʡa�h@N+}�&Z�d�l����ޯV��[b��%Nx�x��.e�(v��\��7y��7&pza@!�[
n�'X�%�1�):�=�1���*�P���*M�	�����6������*k���X����L�Hμ�dy���-������>�:6�qRgl���W�Q�!a��/�@�G�$��4[S\��j����]�����L�=L�̫�y�'S�rV��t�^�m�Ĥ	}ĿM/Y���qP#� E�R���˖���!��J�)8>��Z̕��2wZ}ke\���</� N��{�ޕ"��澖��*<(ī�W�M3���>÷���xu�@�?,��F�gj}j�Ϯ}�CO&�ޔJ����h���j�+ʷ�s1[����v��k�l�B2IuK��߲���2MT��Ճ��^jX3�HlĠ4_K�ȁ��ŋ�`/l]W�g�F?��O����&��Uׇ��ʖ��,W2��F3^���ӫk���x�PF�B�"��7��'�j�
����������Ҡ���|-��tG�%��b�k�Dq$n�ScKDWvV{FR����$,���)T��u�X�u֝7�+>n�uO�ֵR`�b+�Pfj��`#A=H{Z��Ҟ˞˪�9墯<�`��j�Ɗ7m].p���P�?NS��|�8r1"_ۖ�(b!��}u�D5��VK�h�D�S�B��r;[����43:������!Sk�{����e���T|t��h�� �@Y�k/�g�;
M0�M+���Q��^5z��uָ8��9�������H�c�{�`S�+���
r��k���6V�m�ˏ��+�,���C���A����S�=l���-��S�
���=�9ߗڽ�L� �2�*�!syӖԊ{�0��Ε*��Թ.ϵ=_c�!k�]�ie-�ܰ%��NE!s`�������ul�d+����E��菢��9̕w�Z�GR�*s�N�6�p�!G�}�BdC"|(�K�$
"!M������O�
$�(���W9G?Iآ"HP��Dm��"�b4�'�XDv�U^�(��G�D(ߗ��(��Tj�ooZ�%J�C�K�]@�M��%�J����Js
V(�,!-Db��J~\�n���ٹ���p{��$�^�Ի��_B��v�z7p�9�Is/M���jBs6m���.���c�Sepq.�jW�<1%�,��JN`�k*�i��]���N=1dƧ�r&'-�����[}����Y�)
�.�������Iq_�^�~-9 ct�_54ԌUS�`��g���?Z���#���P�Ը$�"��ڕi��8��6��m,W�}A�7gx��G��4[dS�=�v�_Q`��Ԧ9s� o0$��dY$٘�]�V��^��xH	9j`���q��-}���/���+O���h����S�I�zI�����ҟ�ET�-�SmS0X�#���QM�30�x���`d}G�0��Vň_d�zl��`6��}�J�������'��ȼf�z�M�ߟs�B|��*W�>M:�)u1{�
�0��n���+�O��]��+���S+�i�����j��2Z�"�D�֑�?L�e��S��J'[�Wǉ��<ҵ�k3�Z�"���Kq��]���쇹�޾�v��+|�}4?�0����-P�KB��G׈ �j���ۯ��b�kǋ<�+Ι�~:�gaLݥ��1J�-����� ��jQ<���2O��^�iz�j	��N�8��4������Hx*�7
c����J�|�e���Wi1*s�_]Y5�|d�ھ����xڍ"O&л�2�R�Q1'kY��)��f�)���\j��	Ovk�'��ցvr�����kշ�n����sv��W�>M@�Ǹ�hI���'��l'?@lE/���T^�P�!x�oyJ��pH ��fF�+�*8��;�wǺ�ϻ-�9�~aB��!$��7�4��G��ԡ(_��Mʸ�v4�����˷�����Ώ���
%�#H���M�?�9~�zn�J8���Q�R�jS�2�y��ۮ�}��(�JHJ��Q$���9�Bg�Yޫ�і(�
Ȉ|�e,�y�*�7#��r'��z�K]�(����W��'7�e��[��gk8�S�2��h��6�x���F����5�N��u���`o ��N��	�=s���dF���CaZ�DUW��5Mz�A�*h�鼿���rB<� >z����C���Qr~��׸�4Ts\�;�v��gt��2��ʢ<������}t�>.�W,��壘����%Ri��*��j{j�˹�ۂB����������Z�򙉊͈{*r� �EO?L�ʐ ���zROV��tx&����s�,^w�� �:���g��^�I�6;;��W��O8ڧ1��kE ��9`3M[v�A�J�-��a�O�J'��8nVߎח0)On�[j�y �O}S��A�!��3�����1�H�,i��p��<�šשPC�����W+q:M�2v���]��;յ�ߚ"��vԉ��>�*��F��<��:�����GR��eK�"���a6Z�LY�UY8W�5.h�s��\?F�DU�H����C>o�}�Z$R5��b36TH�>����-��0}m�ݐ�x�)V��		�)�EY�[SǇòq��~P��b�A�`(��P%o��>K�/6E�I�~�<1O�*�/V�m�(+ُ"��Ǻ�0�3�.8�H}�:���sk��>ߺ{!��� 7��f<�T��U�X�8��D�^��p�g�pV��0TzZ�>Se���b�\-3n|�k�y��[S�ez�s�d��(ð�l��Lp�>=�-Ab&hi�)_J�������^�.�nVhE�W���ܞ]����u����H!,	�F�|�L_LKĊ�MN9�}Q�(���<ҔLDa��*���s�_{r����O���>xt��O��x~j!Eq_9씥��ݕ���t����֒U�]|B��J>���;���α�\U�_�%�3���]}��C��3���]т�:��vݷ��Co
�y������n���U�ʒ�&�j�Y���m��N��9��YiM{MSwS��S����L>��>�d���VV:V|�y�|\�(ȧ�};E��o�Eˀ�!6 p��]�qA^t[��zU������M?����!y��]ҝ���X"
���IB�d��dH�J�;�jf)�ɽ5��%BB"S|��/^�d�UӉ\G���&%�m{����}6�3>�3�on)���^����<QdP����^4�����!@ ��X�P�5XÎk��ؒ>]{X�U����`�CE}k��1��ۑ|S����yB�#0�����M�d`"F}�Q��(]�*��ү��]�כZ��ǣ�m�g08���E?�^��~�]/\�E����;ۂ/�X���S?T��Sٵ�W�#�K��jQ�y.��o1D�8n�Q��C�N�)��A1���-^�A�n�f+�J�L� ��2͗y�Q"�i�';�Q����廙�8�+s�0�2�C��-�	ۄ�7}w�G�eZ��ȜJ�O����mi��l��VMK���k���nf��Pn�J����n��S�JX/Uor�9�/��Oҵ
��Ƿ�&�������hZE���W�/�S���!B��Ҥ�/
o�I�|�%�,��dY{w�;�d�ݨ�i��e$e��v�o�o.��zL�O��0Si��Z㯭/�vT�t��!t�ｘc��������H����&��KT�i{�MSm�ļ�[��<g�0wn/C �>�j~�T�{�S�����9D�6�ޯ*��v,�q�NJ������o�'�v0�{�|�n*ZUn��H >�c� BhN��O�DR�)��8y�����^*���;�C௯;:��n�]}����v��k��N܉���p!� >��*W�m-Ŗ��=4$�v#3T/p�U� ��<�^Y۩�&��Hݮ��	������vև���]߄*V[����������]�L�|�,�	�ߦ��mZ5�g��b'���e�=%�Q�����pu��j��f�%�#�+���n���"
��ԮnT��j�T(��r����͙�ي�)rw(���+�&��~=k�a1Yc�V�O�&+�I�������:�s�c��
'�1b5�+���^ey[�]�Ձ�4�����7��=)��a\��~�r��H�˥�嬿����M^���[��ӊ~�o5��A�za��	9����Pa9�Ԧf~r��1����\T�������߈��v�~8�=�V��O�r�+�]���/���HT+E�h_L���z�����ԛ�8�Y��r����2}�	"��0|X�Qj�Фd���TMv��cm�N�|'IĠ�nR�Q{H����J{ܟ�|�4�{����_��#�{p�/�B�}���h�k����D��4��f���Җ���|'��T�/~r�]�i��][�����<_S��㞪agBaXH�"��UP.���,BHyUKT�s�S��U�N{.�|�=�����W:pp�-�^��}�Q��p쟽��0R1xS9�G�t�P�/�����Jz^SA~p�Ǧ��i}�J����)��S����ՓF�kM��fO�׿ZkEo{����a�ʻ���b���7-�]-zzSn�SS����&'_/�̼N:5��J�&�oTR#�&�(&a2Bg����y�]9���1Qݫɔ]���sâ]<f����I��X�q
�~,=Le�ht�WIL�n�d�5����N�\�
���E[*�M2_N�����rˡ�u��-E(�m�<��ںDښ�A8,Lk{�y��z��n̡H��B�A3�9V� q���Z�$��~�D �R�b���"��f[�~s!VF�r�k3��7�hW @7��ڽ}y^n5k�gϳ�*Xp������իD�;,��h��,������Ȝ��W�[{5og90�^I�ySv�̈́U��aǷ�wz����>*NY�Ц��v�ET�z���·&���@��_t���=�]�<��� ���#oO5��v�^)'�'*fo~T�����>s�7�-�;&b�#��f-}1�*H�$���*QO55��f.<g�&սB)qe��^�u`��oΗ/5bы;�����"WmK����D.���c|1�ېu�)V�R���\vj؞}�P�צ�yt�∽tv.%�e}No�5� R*�5	1�J��ӻ� ���ǉ�Ja�觔&��!n6S���
$|�(r"b:���a��c�d��.(5�����0R��ν� ���ݠi���9a��)�׬�wu�rf�}Q%��W*�;}*�Ɓh�N��IپWpk�~g�3��c�6����Lh��10>,�����*"}��=kEw��H�Y�Lm�1�f��RNH����Xd��h��	gX��/�-���f��m��������H���W�2�1�׎��E3E���&�ި<*֨^�U횑`��_'��$�5�߅ʟ�~��\Tix��9�uS�,8��䟫����c�pIB3��v��mpsV#�X2���0t}]�15���Ū��ν1f^\(J}wڲ��)�T��8X�����vq8�U���� 6e�.���̼ĭ�lV�U��sL�:8�f[��{l�6�i���.������)����Zxo	�l��m�q�(�的��ui9�Č� ��	�/�l��f��Q7CfEw�-%�dC�;Wh/����42��b��}-��Y��Z�V�h��ܙ�rƃ��iX���?\ZJ{��J�^�՗��j���F��=�r
=}�EҺ��7����c��wv���<�ö�͈�e��1�����\T��WS��\&���7�DRY}����]]oI����"�Hp-V� ]�Z��Ԛ����������՜[[����+)�R��%o.,:�8��)��/�#�J�N��{]�-:����뛬,���)�eʀ���7)l�*��Q�s�����v$����̥{+�CUfpndU�3&X3�<�'x�mf�̾w����\<G�x/���<�����kOq@�Vo<yR��T�p2 o-��Xס���u0x�Ƥ�{�vmm�1�m\9[5D�2fLV���{�g%;N6��E�.�8�5R�/^�͐b�`�1����̀��&�ۥ���U�q�fDjդp�ȱc,��зccZ�*�_Xk�^��Afu�[u/S�Z8dC9U�ꛫ&�^%y��f� Y�I1Su$4,)tpC�fu�X��8�ziN��|!J�1�j�^g, ���u)��(�N�sFQIICgg^�k����x�(��6��x��+��I��p�Mҡ,�N�	5��] U���#^�Ճ���b��vNo4�̈́�;�X�q5�^�2tO��4z��(�y�%_=�z?#��ٙ��\�&�ݮ��m3"�}��vE#�+��j�����o�`�R<:.����*h�1��⇇VL�`�u��e�R�;�o��B�:�V��Q-�����&9ع+e� �ĳ:$��= �bgQ0و��2o-9rj����%��׎��Ą�
b�,��0��f`��O��̥����ݎ���՘��"�������&]u��S�A�6ti��n��Mf7nKv�����;��w%��b{Bh�:�d8Y�\�i����W��Ź/�0v�N",�Jb͈e����/�%��T�p�]c�,8q-$�1ŁJ�x��6nXz�~�kk�v��鳹�3;e\��t���[��;�,�k'rM�ё)N��u6��j��Nv��r�f\yږ�7[%{=�h�D%
\��|�O[tM3^�]�'�]?�K|ojgqe���;.��o�KkV���­�uj��@J�O����S+b�_TQ�u�Xg�¡w2> ��)�^#��B��-"6TyA�=J����wa�^�!���芃E�&x��y�]B0E��e,g��o�V/@��s+!nٝ��sIzrs�I^�!��>�0��ڟ�y�@��0�(��n&R��F;���	q2ը2�$�_Lj�������z�����UI��jtu��q��q<}6��|�M�rn��ο:�!O�
 ��k�7.���wi��&�^(����+*#$�c����j�dOf{��r���E��b�4���+�ئ��<S�De������z�yw��t�x�t.`�1��q?J�e��@���b�\^[�~�����R��4(mMY�b� ��*r���	�O��x����.�#>����=��ۯ�9���xX�Z���Y+�S��W�͚�����m��N~�i�z�ː~�q�jP��<3�kUEJ>�t�sn��\v�YPӉh(�̺�_T����*���^������@��>:���ę�
2>���TG�ܯ��*�t��ry#ބ�i���pܙ1�$���[�m�E{�n�!z�o%��Q�b�>����R ׻*�GLjd��	��! Ho��?��N��w)�}r�P��j�!/��2X5�����9�����lt�T�0�$�E��oo<v,�FF���Ǉw'�D�;k�Kj�����}E�SJ�f���ua�qUf5��t�U��SY8��{��Nc����w�]������C��Q�>��&,g0gL�P���-��T.ɚQ�}�q��#���������g����(�jP���nUQ��^Y�MQ� �6��%;��8�ýR�l�J�ں('���s�B��xvZ�b]E�+y`�eX�)������-�m�9��Z��E��-��v�p�5SPk+c�5x�{��&5{�0ә���\p|7#1�9Y�6.6g��1�Tt�Тe�bfJ0&.B��(=7�Ϸ��E;�=o�޺�B�ۘa�1�<ØȓB��H�$��P�ڙ\:S����|v��r�@�)�^��M.����u�7�Y�7Hs8����
~}%Tx�[p�0����i־"a�3�D��4N�x����V��L�-c|N@��w����&<x,�nl\�3BP,�)u,�&Ox�.���[��|Yljc���H�Y��I�"ĭ�"���g�BR���.���G6�(�'�����񅼚۵X�*��k����ԩ�Ϧ��5B��mG#A����0�)@�{;�0}Ĥ-�jzo�K���d۷Yj�tw����0�U��Wh�z�A�nne��Y��T����A���f���s�v��LTH�[!�s=2/�D_ZNI�8˨�-(����̪�z)]}ȪZE)�^�K��I{R�1���`yJ�X�*����0�H�R�[�Q\,ʻ�N^���8��|�y�&aLi��s�Y3�Ͼ�у�^T(�(���
�e�� I����휫� �?9��Rq�L�ѐJY�n/z��={K@����T-|o�I��H�E�?x�Q�OЧ��,��f<�d�ko�))>q��ͳ[n�&�m&*`U����-qm�)ݎ7�I�A��~+y6��V|
G.ʛ�����Z	�3��0��T��&*���h
"~�	1�g%%P�b���f�]U/�{Nk��*�o�b��ԱJ�k!n��oy��Ů���sv��]��ٺ�/:h��f���9i��D�X`�-Ω3��l�?�Ʀ���&��|��Aa��o"��݀�٨XV}`���i##3v�;PQ�틪]kU�s�:�����/�i+O�!�5��'��9a8�'�I7��##�J��������R~�_�iص"Hv"Æ����9 F�Ǚ��Y괺��-K�r	[Yx�E	�q3�1T�/�!�0���*���y/��4�+��JjX��+�"�fE���2��B�*����2��@�Z�?&��~�����,EU��r��0���at����238�r����fGŲf����F���\K��W�80GpO�5N&�T�����&b�+���=�8�ɉ �	=���4�[�mg��ٝ�X)�־�rab���*�����b/��`�t/!E�,�� @�a�G�Mo���gާH
a�{n*��| <���*�J=�v���QM;��4��3�(�1�yt�^�f��ćK|����_,͒!r�H`�9K7�*�&{<��E@�IR�#5m�VPK�%<��{>T���$7ó�����3^ܯ*Q�;81Ao���GlĈ�v�e�\H��➬��?n|�!��D|� .p,N��XG+L7H�{��0;���Z:����%��D�NB���.Ni��##�ѥ�牭R%�Jhm�qu@!�y�s�g=�v~�V�j���������U�̋:�8@�V��^�f3�m�VM]u9��R���y�8������� F�"�#ģ���N`ή��J&�g��ӻև���l��.� �m��\���ۚb9�V�V�!^�{��������D��[OE����ʢ���̮��l���+�2�nd��^yM{:i̿x��:�����#��6m`��H�p�����[�֭��o\g�TY�6W�
�i�T����B��_9��SQ����6���K��=62�\�7����Z5q����\��IT�We�C2�5s�)�{,�̜oKm�f!�w�b['z��2�e "x��Ųl�s����}#{p�Wv��"�=�yq���S�16�s��Ń۹��$h��\="oUeq���߼;�с�����b(�����`���n��b;�^)-L%�T��N���S/e��`��{	���\]r͔�;ݦ���p��dɖ�{<�}o�Q]�W����+��.U������-��9�\�]�/�6����)�£g��Ê3�]�U@�أO%�Y���*w�wM�*Nt�d�������/�%yJ?u0DM�X�74��;�2���,��^4:�w��OB ���`�̭Jd0bY>�5-�q�Q��g��3���T�0x� l���{�샑���d#D����R���Y�>�I���L�qB�+>�exb��K�Kj�W����/y����'�)�t�SR������)�}�ƃ���5�'�yGuVԈ*F:b��QВ&#�ra[�g�ʡ�ܱ�QP��P�W*�M\(�N��g��j��O�Ekm�0����dO�j>U>䔉�)i0e�Rbw�*u�����x@Q�2��D��o��C���S�m��M.�����;��ޝ�<�;\Ϥ����M��DC�����B�wp�f ]wʲ��<�3u����BEw��r(=�k�7ح]�&���wA��b���.f��Ӊ�� :�ֈ�����Hx5 ��	.�	ݳ�@���{,�R�aS����[ݷ6�X^R�r�&13jK��U*;��3n�In�ܷ?	�)֍��u���[�Fw]e��6�_���]�B뽍#v��G�rX�/��2��M��j�gyzvI�ʗ�p7�_^[jw����NV���:��ǅ��7
��]bqQ��}�A�69�������&�FuR1E��7V�	d��h�Qk:�z}��bU|�H��(4ܦ>��R���[�=��I��]�cY��p kG�(=�Tg�ٺ��Q����פn/`���3�{�rfaX�/!�N�ѓQ��P�PS�%�����`��U �����m��)m�~���0eL�lЏˈ�[�|�	�9�PJP�Z��݌��Fχ�ڷ"R�l��Ys��Y�ۇ�+��é`���kG�1"�����ty���uF�(ʌr��[�}#�6��
ʣVnɄ�W��H�TH�H�H����鯻�,�����S���}�;j$�D�YUdpJ^�ݒ  �3�&ҽ��/��;7BD٫�S=�Tm�䨐��V��1�^����g���7lh� ��~L�Ж�.���G����1��##�UѠ"��l�Q�HF�a0��'�8�����T{��UO7Xמ�h|C�S��8�{��Vb=���M����gx;�&:q �u�nF�1��U8�/�	B�Kv.e�%��dO��k���a�����^����ILA`Ǉ��b��(O���"g���fba:K���ۦ��:=�����229/�<�A�6�,+��~��+h���w�}ʉ�ˌ�7�!/�qn��|�.V䏔o��ic�R�S޵��|�;�~4m#�Lb�_���8I���7�l����r|�ٵ���.��@}0�o��@�"c�1�aPP#Ҏ�U���˹�;�"��}q�{�Ξ=��I��w��G�2R�z����փӻ�Mrj����ӵ����b�@;[� ٙ�����t�	�,b��WV��UM��b�W+x�	Y����z��h�{��&�c�D���\��n��I�wL�v8��\�ۛ�f`]BT7��4!��	��O_lX�+�ʩ���((o�萊[)pVb��\�h!"([4��O�<��EH����c�#��m�.:F%�����l�K��k�wĴ�Kޮ7B��'�_r���){�f�!ϔHw�_E�(�Q.�_��W�L�[:1	�e���
j�߰LդD�t��wA��g噭K�=&�zj_�$5�?+�Fb�b����!̫Nri	<���q]�՚ٔ���#����s��"�<���V�P'�N�aUi$�u�Y��i��Z�>�Q�`L��>�`[[R�nQ���[E�$z a��e-�"����T�u˝A�9���oB��K��W���4o��2I�c�pHVU�R5פl��0�";�)�HՀdo�!|��o�Um�e���=?>	/������}��  �$��e
��0V�1�*��u@U�7Q�~����!c���(l�en{�ҡ`Cq�痷U���b%J��	��J*�vrϜھ�Q��@�} {��C�V�72���Q0�R[��_M*nI�Q|�za�Z�f��vx�$��}k��4�H1��D�;���a�<�X�M�LJ���ib7Ԥ�P�����1��W�%y��w6^1]�]:�be�p;P(A&��i�S�捻Lt-�j�P�SAYy�s���v�#��d%� ����g�3��� ,���Y��.��1�&s*R�c�7�7+Lyy�H)��W�����A��@�����p��蘽f+�gm`��"NW��l��U��ą���j0	y����aߦQ"-���+)Pڂ���}H�\�f��T۱����:�S���X4�beTO��v%¶���ۉ�y�Ί��Pb�$�c(�vE��eZ��>��»b�(�4.��g���o9��ǽ�=�,B��n����-���r�<�� Y�I�	]|���[T�+���� ��(UG�nW�c%*nT<��cǭ߭�^���$ܗd��g���[<�� �F�̚<a{�)��^ؕ;!L�x`�P�*V��,A�p��|z�]-�jsKv��|s˗��̕#���ե��w�jf��z�����"ߡ��+摽e9ȝ�y}�D'$���\�#m{=�,��;h��AgY�6��7�I�ӕW�>��y�R>��[�b	��R"�BQ=A�$���B2�b|D:y��7����E�]��>GoqX����b�
�Y���r�z�г��l��QF��mg���]X߲�������sG���S���߇�B�i��X�f�.K±ź7V����+�M�I�����p��x�e��b��EI�S<��~4���,�Gxf%�B6~ԟ┘Jɉ)T{��L�����|y��2<a��Eᨥ�<�\2�/�Q�*��� �3�0�&��L�c�|j���\Μ]��%j��J���s���Q�n�D��T��Q�QQ-�d�� =��)�����4����`! @m��C�|̞u�q���{�c3��Q�M�)��V��<�V?U#A}�^!�l��C^;�a��I3��+�4���xm�"� ��g��QMY?!�':5򫧶��̬s�����MS�Q'{0 n�����{�~���WLv��i\Y���7IR]ˣQ�/*RpB)VE�UFU�Hʎ��vs7ϩ�¨� �;7�]�r�'���V���t:@Z��X�o6q[�pH�M��/2��+&�6hl�K�,G��
�,�V$�yl�bfl�(-z�'GJ�����hs ��E�nn��k�@��3Y������v����o�<��v��}�	���\\ڷyt���2���K%у�i6�fN��ua2=b�$r�ˬ�{@Ώ��	����V)�j��O�a=k\j�'�C��o�v�J�b7>�n��#<�����}[�� ���59��ݙ9w~�.J�	d�h+`g�{��^d�}�V&&��d�8Wu�P&�����^:�����)�T}�L��*.��ъ=�z��J��Ajnޟwml�]lȚSMC��A�K@�[���	���'�N���XJ�r#Ƕig^�R�d�[�6�����u9����f-��t�~ڨ��u�H�ja�T+�ck��8���2:����6�&s�,�s��/=�������Bjɝp_��B��C��r8��J4�T̜�^�5C�ILl��a�P^!c\z!gY�����Û�OB��Fy�*�}���R+���Z���1����S)W�.I���� ��{�>��K"��g���R>ؾQ����W��8Qu��J29u���r�i��^PТO�	�`����сu��/Ի���f�V���,�ށ��6��ϯ��nxD�d�
�1��\�LU yn��k�:v���WZ�;)m�ze���{�suX�Eֽ��CJ���_��0�1�Q�G���ƩUP�TFG���5s9��G��7Ʀ�.C��S�}�����_pw豕��_�\rnLkF��U�bV0c��f��^��g3o�4�Lڧ���S8�r��Y����z�QzC�s,_8CW]���*�����{�u�sUJm)7T�;*U�z�kc��)v�Z��|8v,˳#��>��/�i��·d˝F�W3�:�j�5b���Ai�.����%���W"A1�f����Q��^UL�<��@A7�3�zy/T�a���<��	,�4��Ej��4k2c���P�E9���@A������he��'����-��M�(,�Y�vs;pz��ue'�m"��"��G�
�`[_zsoև��DL��]bo��_
4[^T�J2�QT�@�ؚw�3��Қ�g�F=�R�j�Eu���?b�R3.���P-ӯʬ�{���X���jx���-ıb5k�v�}ѳG�ʍ�P�Y��"�R3�W�*h.n(a����+�QB&����J��+�j��o.U�r_�s��k��i;oLeay�8�yA}<�'�ʫ����Nhu�]Ⴧ�2�{���?��l k��LЀ�4�y�&�s�↸.�֗5�ނ'��ymG7�t\�S����(��M��g �w���$^��~��Ina׊�G8��g�%.}��VC�/z�<�7낇fԫ�&h�3��`�M�]0&���"�(��ؔ-"��4aeb��{�����-F"�0�E��3���A��ȣ�>�P�E��qW�hL����e|�-�߯ל�n�t���y~��+Mp��\�'�F��8�"��0��Σ�漙0���Lj����"�'��C���n�`M�r�\��b�4k�������J��Na{,���0��^
�Ni�a�l�}���}��*�����~��9�x֌y�c�[Fu*�a*ԕ7��f���x�+��sqW.gu�k�pÒ��o1�?+�-��2k<ս�-(���KUn6�ڰ�K�H���u�yAw�S�L����{n۠�A���`��7O�Kt�a�E}���V\�?vڸaB�vVh���__vx�4��'\j@B|���p%���u�q0<��ON�{[����l�
OU�^S�o䶽��Fa.��,���շ��y�����`�P�/�F�}u������$�]�Z��b���#nm]b6��T��&�&ip�5[l�u��h���	����������䍃L10�;�[��!��.�ZtV� �7ꬑ�=��ࢣ�w![�G���b��H�jf��M�}N·=�w���ь��8y��
��|!i@�o��(�.0��B�=a#�3�$��t�1�=�����zP1�	��$�s����e,����WO�H\ӘG���Y�Hux�]i�~���NTޛ�iz���Z�����֢�/�O�<ķ F��T<v��Q�N�A���3�C�[�sS��|'j<��z�����;>�`�-�S��,�=�~�[>Ƿ<_�Sq3c�
��d�a����b��u��*��&ZqC�2Pu�!�!���	W�ۑ?����������ZI|*����P(��q���WR:�=y=��gJxlנ�ۼ'7&�}�L�e9���WYٜ��C��Fme��yi��2%��.o��=xIrw��nc������܋�"�kn��tJK ]���aT8ʶ��X����u ks5�]-Q[�Q��왡��q,5�c䀗�e��#,p�à����B��!5���S�Mx�������!�N�e� �]���:�;E-�z'������vk�1���u�ǥ�x8;s �O�h-��ܮ͎3ݹ�qY6��Cwn��.�HPܝX�C6�-��������
S�pW$�z��N�!�����N�l��b�כ��w;�!��"�](v^ۙ���JNx�:�ow
����;c�8��t��i�qq�T�;���éQ6-;Ƹ�y��y˾��ӠyJsB b8�3S)Ԗ��jj���zQ�YF�9�X0�QLܲ��5a!{u|Mv=O��"�2�
���.�tF�}k����|;�mu�C�e4l����CX��� �<��BfL�^�e���N�}ދ��T��R�{�H��Z��*IC#g#v�X Pn��ֺE+re)�57l�[�{�eL�fB=��
K��[ӉB�YL���3j�@3s5���gf���ql[-�����$Z#n�-#��4%�U��D��Ժُ]:�5Ua!�V�t2��l)�R�J�q�����i��([M�k��B��üH�קD�@؅ִ�v����&����j[y5"A�A�}X��5�[�#�l����,u**5ƘX���n�8t	mo"sLU�4�`|�A��.4��RL��']r�7�e���W�"��P��s�d�m��*�I��������_�uu2/�ɭ>��ޓ7!�$\���ӑ0w��
B[!����M4gP��m�BV�X�����6I�<�%B�p��mƶWS�8rw6�шvE�q��T�	�$q��-`��0�:sQ2�س�t�꾺m�wN,�z�V���ع�^���ù���E���W&ʰ��2jӉ9�y*��;.NB�� ���V�0���MKEڧ-�)�U�J�D/��ڈ�m���:��iv[�n������I��̦d���
B��Vfꐋ���:�sU��| NR�����!| 띨�Kd1��k�vc�}��q����t��3�^n��+Y�z��7����\�j���Hk+��5�5.��Yԩ%��m^J���̻�
u���ͪbf���ז�����P��mndQ�=���k�8+���;wrwAS�yFʄ�lV��#ISӺ�z/&��Y��w�b@����h���W@�6��Z�,�+9'�kY�&K�q�L��jsTJ�Yi�Jr�s�*m���7P�۽���S��W���vɬ�����0��+����t�p��3j�̬MsǨ똅l�QN�ow�5%��0m:\z��CR��0R����-��ڕ�N�ɈD9c	x���5X��e�ĺ�ԗ\�*=�����L΋��]��?���ޖ�TG7�Gi%�Å:���Ъ��Fb�C��O���U�%+7�J��q���I%|�����|��Wy8!3��4�	7�-�)����������qw>�0u3V*6i2
fY�E�V �O�̛�������I����V��̺�)(�n��n�Cc�Fl-����ob'"4�[�U~��gEs�NQ�8D���/��<��n�m����e���9�5�Z�O;�+�DTdZ�ˆ:���z�Ɏ�r#�ӕ�s�$��.�v_���7���M,1��v��Qy1LD�,ٻ��<.}]��u�}����M�Q)ײ�����y	&)e_İм�0�Mc/P������6}鶅hE��^�������Ru���Y_x�`��dsϼ�s�N��h�̽ŵZ� �> uo�#d�)��:�a����Z]�ڸ�e��䀀e�ݩbj�ᜡ �[܃�Nt9lsӾ��{��'o�����РL�{n�苵�Vp�颹Ay��ݑ�(�LK�s�tuLnyD��H��M�X엧k�<���3���C��c���I�i��fc�n���Lz]�b}lg#�dUA��Pfz� U�n2[���b^����!����[պ[�a��̜��t;ǥ?i���<!)��G�Az��m�xb�,�
W]R'ǧ&؊P`��G���]WRNG�ż��^r/cބ'�RyT\w޷���T��⨒m��6F^�6���7���iGz.�Q��݂.p����~[3�˱,�Ý�V�h������4n��z#tS)�B�d���]�π���	�9�C. Fy|���Ί���ε-��X�1pa�9�d\B!A��꛽ӓ�:��`�t�7Z���Ŏ��V̓6�IH�e�m�ɡ%ꎯ�6w	Ԏ��h�t�d�iܽ5�,�.ֵR��;����b�e��x�]f��5X�HYv��r�*x��\,��(j�~��8b�������[�sN���"�CqO�~���������2�xy�jg�
�г��3���cd2�L�A����8���L��ʧs!D����y�y_ܞ?N�y��i���t�T�E4�����ɘ��Hd<�|�L�]�I��2��A}���E�?����o^qWB��Q�w�t�;p���$��ʍ��\B��f�rh�u���)�����93V6�J)Y��WzpJy"�L�.d�:�W{���/=���>�ih�Dt��ٍ�f{s-̌��Wƙ�v���A�
\U��+�|��Y�=�wtI�xV~K�jm��(���6T���t�,L�sO�-P���	��<�2�t���fLbdz @>�:��u�z<�$�\�x/�g,^��dM(ay�����5����Z��s��X0/	!���۞Y�9�D�mP�<KE."9s�Br�6l�g��ۮ0�+��b������O�Qn�,({��phO(������]ӵ�v�%q����n�\z����I;C�%%�/�Fi �ᶟ�8�;W7�BJ����ܸqSf��'�,�la�:W�뭼KV����_�6�H����^x�9J�yc��7�]�{��.��ϱ8��t�E>��ݱPJ�j+=�U�
�s+χ}ji5^P����oM�����AuL62*w:�Xsq�Y�&i�~3�� ��g>�nQ#u ��pJ�TkD4�[�3q��J�bZ�gnt�"��?c�'�yP yC\�ɜtZ����5��:�m��md��M�nc�ݘ�X�S��}�NފG�~�\Ϋ}Nn�e���9�Vu���&4@����TLQ���+��C��4���xĭsMy{o�u��]'���C'��)y�^q>�t#<��p���
<f+3�}�a`mr�>7�x���՘=q�1L�Ω0��D��͎��T���ˇ�,q�)��M�F �hfs8z:E��"�y�Q���y���QD�4kS���~a�[{��:�n�~���0utF9�V���#ЕH9J�@�H��k�_������2=c�dRr+طo��dŏW�It�A.3S�-4��Lp9߻�&���,;��N�b�bx#�<�"Z�O�M��R�rg(���%|�h��=&�.TB�/�}:�7j���͓JE�U)�ˣo�y(�<cكEt���R�n]4.t\�4#�����ȳqw�1��3u�_�`m�&L߳�".w�%��cek����4i�e�@�;<�-lu�wtӓ�+3241G��==eA\�mG��� ���G�;�OZ�ޢ� ��7[e��h��v���ږ�^���C��^�}P�5J>L�UF�Ns���= ��5���l��51�ʆ�r�\9��c'�#���ޫ} 1��bG���c�j�\�����_؅z�K�89�L��:�ҋ�a3h��I7(��)���!���ݧ�8��ܥX��Z��@.-˚̬�BM/��J���m�t1%��c���ؠtu� c�
�R�αz�J��9P.U�����B�&�����#�'���s��3�EUۛ����_������d�U�B���+˰�ZLA���{T����7,���*U����V.�|�L;:�b}t��|}o���Jpl�Z�@����9�ܨY�H�p��'�<�.�WkQ�"�ǱY{�(6�8��Xo���q'�N}���ث�h���qz�N\yE s^u�P�^��̐ԭ�0�[q�`	E@�15[>֎Fi��a�H���H�,��^�o!8(�=�x�(_�s�u�)��S�����5����`
/}>\�4"�� �Udۢ"��{nRH��PcS�h1-�gFE�����J�'p���#)�C3}��yj��'����E?ޥ{�>�ě͵�G@f��Oij~��U�%�StJ��Q�T���f��P4�����ad1�'��b0z��Z�T�7躥7�$� ČF�U�xO��+�A4G�O�1`n�T��j��&�z��]����@��,LixT$F͋�WDۧ�8�wW�������5�����vU�5?br'0����[5��! ��W>v�����;������ 4w1B�J�"c��M2�pF�ܱ�̟z�e���H��)-h�UOED�^ΪL��3��B0���9���NBB�G1��8e���f�&:'O"�;Lܬ|��q�y����]G$��Ğ��r���r�nCEWqƎi����ꅒ�ضJǹ�zHh��`u����� ����h�D�j��y�E�,49���nA�7w�V$w,0N�2�0��Q����0���$�M�^���')�`~������0���;���M5+�Сhgw�҉sUQ	T\�x�n_�T��G�ע��,����3v3�`v��'�T'�I�X/\Mm��5�Gݏ����S�}t���`����f�W�]]h����1����\}/5gwŸ^��e�s�^ё�v���ߠOzŻ��R���G��W����Wk$>?K3T����_�:E���܌��닚L?sM��9d�8]�KC��%K��	�p]Tu�ً*J��q�?]�S����=��3r�Ҷ@&.`�����CP������Qۂ)b<|aᒔ{����m�@֕����uy��7��W��"M[�E�!�tW�
���͕�X6��VǮb pz{�h��򁸼�nVN"��yZ�W�=N�F��J�����6q�(���6��+7��x��Ϥ�o(V�aK_NE�q��p�>o7����<���W���Z7Hm��"��^V�VE����BOiW�77�*w
�̥>*
�=J]r�_��ګ����z�r���{&����M�xu������i��L���+J�U#�~��'ϜR�����|�5sb�?�n�5^
��uQ��"��l��I��S{�%�p��*7�}Q�u�03���^�� {.��S����2Г������t�`��ok���)G0�㵏o��:Yi�?�1���a4��~9{.eȒ���&� ��jb̫�κœ�M�9��5���%��9��+j���~�r�V�B�-�	��ܗK�U�ڏ����}hd�<M�{�W~z���/�v�B��KL.�pn=V��]++o�H��u�<��yhl�������4���i��I���p�!���A{jV�#��"�G�J�F��ΥG��)W��-@�[��dR�E���qS'ya���((PrT羨k˵yX���8&)hOn���#@)�����;f�/��c����'��Q[��ƛ���{�{� Q�D�U�CUl���I��6-l�w�{�|-�Q;aL�����Fҵ�M����.�F�#v��MW�a�0{j�m������m:�k*�S�������aF���M��MN�fyT�U�kfv��3�Ԏ[^\Z]�������W�q;q��5of��궧(s���� Lm'&qvgV�x|C�7&��=3�Z�~�����k�Vf/��Y~Ҟ�+��jb���Y���e&��9�=i7b��Ř'*)�G���3.˪���k�1��r�J�pek'�����~�5�Ez��yx��|�Ӌ�J�}b�R }�'e/]Q
�ӣ&S��c��F�����N��r�\'��	���f��\�dϟ��Mޣu��g��Cc����l���,�T�/Lx/�Ұ�ʋߜ_��iE�<~q���g�|��mG����3�'�����Tu���vSp�ݤ���C�h�jC��]�Ɏ+�d=O4J'C��EY����Sg ����Ӡ�oD���i�ݱ�x��9�so*�D���k��j�2��7�s_,��_D�����������V%f>�{ȓ���nl#+� #�?@��P���;�F6�f�r)���_kKg���}��kLWݷ����N(��Ht�̛����zp(��$=]�G�\��ݿ(3�Hf�ɤ>ڤ�k1��|����هY6jl^v{0���D�{]TP�<���TW���dU��g.xE�1٘����5�|����Y��Uv�w�2�y�1��'��}*�!gz����h�n����S��9\ƔW�g^1��n�o=7<���酲�x��8.��g��w{*;4 g�}�9���ݓ��"7ڳ�;g��!Qp�(c���n�]�����Ε�s��Stʁ=pEǞ�ӆ���=������F@�-��#��Y,�+#��ƣ�{�5�d��B��^�?��t}�21/騺�`>�Zn��"�\Iګ�deA��D��S��3��+�.�:n���~�%�y[��=��SS��n&���j`r":N2�>�P>0�E���`��I��ڃ'}a�X&���V���ӑ5���4w��9 }Z�0�ق�=̖��?r����$�_5�խW��wtƑή}�� X�Uʴ�Њ��|.�O��F,�΃� u��l¼�øZ,��;��+J1�Jbk�m�H[i�� �,�mU�
�د]�K'8�O�%?1䠜�S%C�c��Ig-�Œ����ن��J$^V��ɜ^�4.�*"AkEWXB�Xgc2�f�S#{s�M5*΂�㧚.��ϻ��O�Oύ�v>����9��"�sT;s��AU��AOQ��h����&33�<+���v��%�O\�QY���M�=��V�W(�C�7<oش_]������F�>ͪ�#=�l�O�T�}�T�s��'�d��]�z��~�N#fߕ�5���O
w�eq�;<��&*=�[8��n��;��zV	�u�����,�r�:��8���F'�%�WYZ���k�V4^��G��T�|{S�H紨[)xH�}�x\�v�er�4�y�NO�����3������ZU�y���ͬ�|�%��z=�U��\��xQ�w�����yݘk�����9�� �c�t�Ƞz�Ӫё�,����|<����/���J���Fr��'�+�����+�ks"�����?e�)�v�1�}(d��+Vv���P=��=�%{b��E~c"(~���w�Jc�{5q��t�Vַ�Uf��?���fS�R[��=�.���5���aC.qɇU��n+�������y�q.�tS`��]5FFy�������0+=�Z>��}3$��{'n���bS���O�y������H�hm1��k��T�R9�}p/sB��~�$	�l�%��-^"��GZ����0��;�la鸧s�c2AH�V.f<n���͝XS�7�J;ȱ��	�w�hs��L"�EPOv�=lI�oE#�,�<���۹�iȇT��3j�7/y�]��̆^��[N�2(m�;(�:�y�2�����6���Y[1�`��ӊ�^Qή%��/�yHK��%P�j��>V�MF:�מ����I��.�j�J]��]l���f{�_R�k�a 5臙Нv�6���үx/���=*Y_,t��V�|�������5Ё22d真
v�u��R��4����_�����qa��d��ʼ�^�A�2̽�#{s�j��,�v��Yۉ�������D�]� Tp^0��*�C@�N��4�$�����&���+д�U�cT~��p��u�e4"65��s�X����T{��yt��.2��09�W\��bQr��x�
�뾑��Bn.����@
`[�1֗��;]�׮�_�o�/��^�ۤr�}J�j��=G���b0��yé2�+�9�L��S�P��O���}�{��W�}��A�·�:Q�0�Et8R%�~��Ί4bB��p�k���:��L�׎����$��<X ��yy}>����X��|�p��E`����5~���MݵH��q�:7�g�:����Nn5�����wo�������k��?f�^�"tH�B_��z<���]A^S%��&˻�*��͸���yF�^�V	���)��i�j���*N�\�nV�56�Wikw����h=H���sT���y�Գnί��g��]�C�铮�%��_t>��eգU�ʃR��'pݭ��+F�72ؾ�Ֆ�5Q�Yr`躖�fF���&�Z��ۑ Fl��;t�#V�f��:U
�,�~""=Ƴ�Δ�K|��|>�Sw-��>�d��vm>��^I
�GTU�FFF�Հ��'��Z
�ݕ@�����Y*-o֪Z��[�)�0�t�X䜇�f��m?et�ս�u���{P�X3��Y��Ò��L��F�=�#'���1ٕ7=��ӏ=p���6��y������^Bv:�@�3�A����4��)�v����=�Myש{Z6�k*��7D�&�l�M]Y��S�<��_@���)ԹEq2�g#�0�u�NK[�nA��t��yB�Pޠ̼5�u.�i@l(9Φ��%^�§Q]�^��4GT0��P�`�Gr��#٦w��պ�]�8K8X��mU��fn�P���N��O�]/�oyr���sz�Ղ�>�{X����D����뛙���s��t:�n��2Z���(���,�=>O�_A��%'f������tu��\��+^G���5�,��w�E��*��b�!��A����V�<'ϓ�j��o���S�ӹ�%w'�]`��t_���f{l�毺�t	2����ˤ���9! �8���vK�`���@�{X�����8;���F]/��L����&Q9;��{-C�|�2j��I��UY㕔�Q4��߬�%u��u7��7I��.�fNd��[��v�[4#�;�����{�e�}\o��Ɏ)�:�ٚ�k(���g0��//��n
9�y�I�����/a@�C��s��X��L3�ѭ�tvi~㙖c0�{�,��C�9�gК�@"��F$.�5�X�vul�ǥ.�]\{��w(�KU��y���y����nZv�{t2��n`�#A���.���٘iVe������堕�fsTx�{a��r��:�����wE��ƭ]��i~�Vч�r��%pҰ����j��`�gV.�q<��T��+Sy}�{����:��]�"�t�]6����K�ɹ�_�b���t�ؙ�%iD��*ΈxL��]\#(��mN37��7���[s}[ֵ��D����s�q���w��b��D�O/,�w����uj�b���}�>wWѺ�R���j�)koW5v����}����9U�����*�"�)�(Pܥ�:����l�W�+۱�r�)V9X�Z�C�Z�{���v��=Wպ0��n��Q}�ޥ۶S�*	"aq��9��7�
�	�9^�oe�!�SƞЫ�7��IB����| �ef�<8�6k4���v�s�Z��]t;.�{�`zm�VjX�7�b�]�'�N�F��KU�f2^�\�V��3)X��L� 8��]2#O��2�M�Qs��RHsyG�:��C���k%͟����mg���_^� �x�L'�)�:����j�T&�ܦ�O�VC䧣R;K���Ƚ1j�L�rT'!/(V�����Z����,��Q2V��@K�������H�)uΝ����Kt:��p�Pޖ3f0��<U�!��ס������$!Ϝ;/��\�i���ͱ(U�ՐX*�l���C,{��yw�N�,�����1�{�yZ�D�jVU���_h|53v0�۽]�/��J�e��K��H��%���7{��wX;r��#y�z���p�I�ҏ�b��)��)�S-��}�4���_<x�Т�	��f ��s��!{C�>��7���֙B5������?&0h�!��YZ��Sp�������΋�ڪ]t���n;��j�f�{�iwY[W�ӯq�x�OG�ۢ�A���K�I�]v�#
�n��r���q �-Y��dn��	��D��9*fcf���9��Wv�E�s�<�'AĩlW{����ٳ�M�ٙ�;���M����"��Y�U�Q�z��8t��b5J���D-�\;y�c}iݎh��^�Z����Ĭ�ı�ʔDѺk:7�i�k�8��P�3.."�\s6���韥��n�����}��v@zo����>Y5���{�;h����	��W��;Q������ݮ;ԓ)�}����Y�]\�����Z3PE]�]��Є�P+$�'>Dq0'c�TaYƍ?��G����Ң��;Ī��1o��|I�~�nj�uz]WNމ�M�V�ݹ9�0��̼m�̢dŰ�v�~�9��a_jTs��e��I `�N�:��W��vSY#:ڏ	�+�s<�ňwk��<��/m�v�e鸼�8�D��r��Ld�+�kv��ztz���c��IJ7aCQH'"^Ho	__�'��Lc4�p�um���>�J̍�i��Ki�Gb�s��#��h��!����d����6Y��=��x�k��ҎF�b��S�%�fr>;
 �W(]�����5��i*A��X��b��/��<jK��"����m�e�9�u/<U����f���H1�0�N~�`뱓�Y+X��k4k��GB^˳~>+ᚒ�Q~Q����x��c��^�F��\��̰�WJ�#㣙�{�H���i��T��\c��X�X�uAS0��ɥw�]Z�Nyy��v�qŪ ��� ���~>	ܞ���e��Un��O%G�x�s�}(|���w�X3czI��3ݪ�2�r%&�A��ڜ�w�|מvf��� u�G���2<sQ�T��(�sV)�Q�]����c�D��m�ͨD�^uz�����իW�'���%~�i#D�~�&��f�1��ρ��[�H�K x�+�1q)z�ѯ���3�<5tU�r���jƳ�7��{ <`g)�IY��{�B���@�͝V	�|�i��T�@��y�+����&Vfә�N ���Ȇ�	WCC�u�ޛ\f��] �̌�P�Pn�iƫ�f��	����/i�w��+:q�Y�_t�S��������1�i�룄T��jz��ћ��q�aI�q>��i��ڈzC�U���������g�͑�Ά`gm��J����9���)⨯BLO±����]�����g�����5�=�'&���D��6��ڄ���!�t*}���J2Zw��?	�+�lgyHq�0u@!�#��bULL���Q���N�EW��×\z�Y���z���{bz��FF�P�μ�h��ڮ�zF���C:::y�;�X甬�9��'1 �au��⇒^���}h�X�9��O���x���;~��
mG���o�$���$'�с<>ChhI�+���*۞�Tz�u���s|LF�m�q7g�ډ�����/x^�އ��a򊉻�&���7w&/К,E_\� ��#<m��L�{Ǯ��5�(�^�����9�j:�\ݸ]�p��*<h^#1ｐ���	���J�m�{���皦����X�b��{aJ	��N��E緭Q��W|'qb���4�.����?-5Y���C��zvX�i�->�'>;J�Y}��uz�b�����]�}`+Ó�KZu+G���<���[jƬ���їJ���ԝ�6��Yť4Z��Dkm�=�5z��KȷNh\쭶����0;�)��릷9�op���ӫw���1�דTВ��x��Ck:�{�t%���`hf����KI�[ѥ��^h+����eTsn���1�M8����7�0+�qdΜQrnҊŅE��mS���{�_8�^�AM%��f��Ί�&�ӯ1��q6Lmt�}�ʿ�]����O�]�[	Cޮ�'��B^�����|Qq�{خ�ʯrYY��t��zx�_8Q���+�SmK?<�	l�4\�m`��.��[�w��(n_���Ş���_3�CΥ�����[�gw�0�XJ��������Q֑�S�s���xd�ÿ���;'.w�u%�hb6�x����N�w���\o�ZN���Y<��C�a�[*`�T��Ծ'����a��m5B\xs��or��Э��н�k�ٰ��\��KS�.)�ͿG[������S~��/5�T�0� ����e�=���x^)��6xf�#&:�|$�W����-��*�x�'>�26>{�԰��$K�izV']���Ã��rD�q�Yछ���p�9�>�eZ�W��(�I�"\d<��솟M�is�N��U�o���s�]-��slI��n�J�J�����=s����z�$淠w���5�4NF�.���T&�B��7+�n_��y��s"*���o�CɆ(ygV�Q�]=f��h֛Q9,qd�[�$Uʳ���R��e�wse��1���_<�c4�8���|z�K�J�s�3m�7]���������~Ղ�^�Wm����b]ZB=�uH���p�{vx�����v,Vvt���<Iߍ�;� �x�[��6�6q�˴�Kz��YP5�v����l��0i��m�»�.E I�-0c�s��-����펜��.�������U�{C~�;7���ɫk�g�����ܵ�z�%د��jh�:B�|��/G!@��D-@�희���\��I�R��6��ħj�g��V��w>��3x=���W(N#;��I�C�d}��'}�0��=)� �Ɵyyz�Ǭ��y�Q�b�ve\ޭ���=J��u.���� ��o�"�(h�򢏹���w^s�;��o��ވ��R�q��Z������X�r�p��R��D�}�y���J�{3&x��w��k;�n��5W��uEX�,��]�!������,jw
���J%֩>j�׹=��c�yP�4�i&D�C7�V7��p�uI�CS+'�2Q7�}�Y�$Do�t`�زA�*���>��J�!y��x��N���z�o���a��3��G����%=յ僵�S}6�)��^^�kU��5��gm�-z��=6+���.�Z':}=��P@Ke̹��R�Tc���0ј7}r�>m�<�&äs<\��k4��(�Y4�z^a1S�����Ǔ��pԽK�M���ut��>�/��m737�#�^��Mѧ�(��|��ȑ���mEfҥ��G8X��Nd}{�w8*�ڣ �f���Z��x���F��a�vג��fPk2��P��d� .�����5.o��K�?e�s��'Ӄg
�y��R�71q3yV�)^Y[��Л�P��wg�H�� �kN$��.�հ2{��G��.M.g�y��;��VVׄ���U.�����nIV��
z�um��=V8�'M���1���Z�ёt{Pq�������� �|^���v3��sv��lę��ݹ|=y4hӘ��u��r���z	������ي�T/=�3�v�cnWI|�h�Zx��B6&��R�KXWi� �'�=�UĞ��qX*����]��kk�X7��M�矖�'�_�0��Rs��jK�\��;��c�8f'�'#Ex�I�O�u\�S�*|W�p�vP� t�&���n��R"�����t`�1ᲆMq�xģ�P} gU�o(o�M�JK5E�Q�G�шF�* �A"3wF�v����zb��u)�8L��Y��f='m��\}������>8҆׳����n~^��=[����W��匆�O+0cҝ�MmqC�2�ݼ�Y�M�	�� �Yy��6���S���38��[��s���������*CeVx�g�u���O�hƋdH�k�"�� �yIh�M}Q8'u��mڰ,�k�}�����;)��M�K�N���Ú�u�"�<,w?җLٮ�Yw���k��+����*�Qn˕Ơ%��'5v��A�-�y�q�1�`�mե�3��n����&�j�?�.����:�^��瞩7�ǶE���C]�WX<�Ê�!x�W���#Wo���ܹ�pͺ��>l�ƗHqU��"�J��X$��o�-HǾ�A]��wu����4x8�W\%d{' k�F�g�F��Nϒ������L+�N�<c���3�kC0=�׼22�Vά���<'�pAx�vӪC��*5&/ʎ�H��)����Q��+�ax�[�|��q�6w����w�����Ղ:Ȭ^>jfU���!| �w�&�K����M��9���>9��#B�z�ƭUޛ�aW������e��ݴj:Ǘ�c���/�Vo7n���\oִ_��
5������X����b]#��@�U�/�����4=g���^�.�1������F(-t��&�`ctDK����m��8�����@-�wh��|�	�A�|�/d�! 婠v�|.�^_a�t�%GDyn`��2}��|c�zol����%<�i'=|��ޱ^�:wy�����3�-@ς��Zɖ!1��(a��}d=BgY��@@���:l��u�t�Y�m,�)���&��1TƜg,Έ&���v̷
Ds�%%uz]j��)v�H�G�W�O^��[��"�*ﺉ��w(�mPHIH�'v[ ]�Tw`=��=Z��o��$흚Q��X٫�9�������݇k
B�I[�xFy#����3s�6�@�h���{�C7�]��Z_ʅ���m���/1Bv?y�z���E�8�#��pq��9<�b��k�߼�p�3���O���ޘ�1`�ʿa鉛~['��B�.��q�ut<�����dvԓ4/ateH;P�g_���L*�v+B��x����ɨ��!=i�>Xsx ��'�,���=��av���F����l�ծ�"�>�EX����U�o�ѓ��"����oMx�E�7k����۞��.�V�]U���K��Έ�Ʊ��zE4w�q9p��C������ܡP|����/Zqz�W��%s����G��}P�(R�["ga���J힎"�1�ls@����6Jw۲w��5�^�ӗs��c����r�6	�o\����V�	p� ��W�yz�\b�_���ԁ��\�deeugo������Z�ݎ�j�&5�Z��c���׻�*_U����C|WWV�����]rbn�E�w�<[q�f��1 �^��;\���4W>1\<T�f����d骊S��Nr-xf;��۝ {3��*�	خ<�=�V�}v���Š�	;ʉ�`�-�­x۬=y���-���0���]�V�cl�oll��z�h��R�֍�|]�N.�R�%�f�y���׬�RA����*&Z0���bP �_:b��y,��G3;�_l�-
:�͐��Tz%$�ӗd?I�V�f��cT�6�ѹ�3$&/��XR:kR��\��x�R�uG�p��kY�Boё�.(i�Uƽ�ۮ<��\�u�F��e�I�rF�e�y��)���\��p���uM�Yj�~ݒc#��/\õ�o"�����H&�1KQ�*��t/:�#�H{n6r�(	Gz\#[�9�Ǐz��mݕ�i��TZý�n�@��d8)�J|���z��'���]"�.�vN\�"�|�LJ������ո��F�����f�7��r�Is�N =�/�N(���0Tzp��A쉼}��;�g�t:yg`���s�Rs���޵J`Wzm������O�'}�����&�f_�1���\�גF�Qrf���4i�ԭ����(��}֮%��M��k�Gg�ɟm(�3R�f���G��%�~�91z���j��LcJn����E@~��7�|f�)��(�Z��{"����9��{54�Hܖ��|��U0�"�*�[8����ҳ��q��\J'�7`�頑^�ռ����iJ�9��wԍ��D^�P°�99ۜ��MK�Ô�x��*�ݝ0+p;�a�˺���*����������e꺌�H���UФ��ۢ�k�Y��Ҟ�	��2d�My�����Wǰ��师[��h::�:�;�T��'X�ǈ�4�D�yB�6��K�*R�Vc��*Y}�Ӑ��,��i�57�U�z�{��]\@M�6�z���Z��0�,l��� I��ȿW���	Ɋ
�T$T&����释{.F�4�1�}>�
ǫi����!l�Y�z�&͒fqqS���~�~v{ᷱ�Y������Z�_'0�3�Û�=�n�����ݺte)t2X�7��K٭�6�Y�u�FA!Z靍��y��#յ�Z�`T�	�K\2(��,�����]T�����_�j�#{�d�3��@�����A�1��c>��YG{#��_X��v��N�1��O�R��:=��r�3���`ZӚiw�v{S�f3/����^�����J}��uMR�6[���#��[]=WkV[s��~���=^��%,�{MP�6���TI?W+�#W��ö1H�zP#�����(>��#�ǽ�(�P�p�ʅ�X�-��'��.��[E��53Wy1H��^�TK�J_R!?zJ�mw���2�A/S��-cB�/��w������B�������L�4������uL��˽��5�5GQ�5�@�#L�ɉqG�sW�X:=��J>��O����TXp���oq��V_�[�F+�S9�1�|�����B+k���I��,U��lee����f��Z4E��i�R�({��ٻ�ͧN���-�9�j;�����՛�3�ᐽ�5�]؟^�h����"����!3��j&>TQ�G�1��s�T�?yd���Nc��,�e	�&��Q��~�Ӎ�'V�VYTe�����w�=L�Fb��H�y�UEm��R����2�<����hhg}����ʻ�|���*�,Lr�e�z�ʴ|�s���^Q�!	�Q������(�#4k�kd �r��w��ɤK�|�PTZ�/_J�w��ܕ@��������9�i���8��Y&&�����t�d�{c���x,՜�e��[������d |ڑ��@��dd��i�U�],�=8K��H�ٮ��"�\��Sa��jG2Lz֘��Ey�m�)�:���8�)�.�(e}�tFv�N��3uql ���~~�=t����C^�u�|<�=9��!m�Ha��	5K�Ǣ�n+a��_�!j7Cn��w�&�u�oP�����`����%ĸ~�f �}��0r�Q����i�X��Ֆ�����NX�=��9��]B�U��E�ꌋ��z��\5�M>R���]Og=��ۯ�1+���m�,�-ۍӋ�7}�_vy����?PxML9�/D_՛��rD��)(�1�P}��y��.u%h��mF�乪 �l� �j�Ulnҙ�_<��4�\�,��u�f�5:�;{ �z����bțyv��۽Yw_�m�(`��f��r�?��]8*v����Nu�"J3�Ohl'�
k���C�v�D-�Z5��k�d�v�8�!��|0 �۸Vj[�_iG����3%
�1��ن�/wz*���obE����W�#;���|��ՙ�pu\.��g&^L����I�Fb��cb�)�@�r�if�#����s���*1��8��^u�՛&:�b���E'���/�z�ٓKOq��{.�+EEb��T�4h�Ξ�JM�t:����y��h�^�.�w����-����v&*|cجn��o���e<ZܛbT�j��e/n�/�%�e�HT�;�yb�����r��ƫp_n�{�78��ᄱ|�\Ď��ܹo�
���s�6�]�¢a�BJ�M��fs��N�wtT��G��(����a�ι�������u	-�]Fҫ��Cb��;����d��J�n}F����첉e����7u(��a];��Y$�59�\�Y��*5,�
Ծ�2�n�ᩧ�v�|ͅ�Z�Ⱥ�%6]r��2�4�E�)u���?�Y���������T/^�tw�[�2��6�,��Ze=9��M�������9ZPR���������_RR�����t�Ȭ�fX�[�*U�K�Q0��a�֣�����q���u�w��(k9ͽC�򧎂r�I��+�Bm�[�`T��8���V��-�ݝӷE�&�"�N����u�LN}/	�xc֫/*@�&朾�uß>S�s5
/���U>q$���Qm��,�aۣ�\Iq���V�R�鲑5o�]mAc�.f,x�
�n-Kn�ޓC>%�JŔp,�<n�q#a����}�GCF�-�'f�pҨ�y����03E,�6�z���Bl�&�8Y����=MM%R�W�fN��޲j�f;2:Z- ��T
'��[�5@\=-v����[.�t��U�Զ3"Ҙ���802<E��Ԓ܉8(�2��f��}�7ӵd{�eՕs	��M+�`+%��x�A��h{kvT{Mw�Ge	4',�g��rW�+��^��^q(Æ���x�o�|�[�ԧBd��P���/�T	�8\{�"h���k��~#gR���Jv�K�x��楴�&�3u��:l�b���c�@_M�Qb�y�e�����Q:��-/�L��X�A��wj'+��i*���a�
S���i�r=���nN�Ve(5n�	���c��Md8)� �t�8�ā��J��kw�1�� �VW ��˽2�F��C�֜��n�2�	ıx��D�p$܊����x�!��wE��+��M�%]���P ���X̾��ޣ�����I�����w&m�6H�%.PnEZi&�+�R���&2�Tq7#�]b�Ԋ��\ضt0'i��˙jd�f+C��߲�BIB+�ճާ)�3O�s)|*C@��������U���宥f]��{�w�[��kfd���Ad\�K��b�ow��D������t�◊f�}x)O�i��44o3�G�V�e�VL�]�s�྅F�D.���v���oP�ʣ=3P��B�:��v:l�ڳPP�Ұ*ZFƛ�L�j}*$w�;�ǎ��1h��y&��5hY����;��d���m=�ڼ��>;�~�#�V]���/����a�b�K���SYˁo�#;�B7��HIP50}�"�} z)X~��/k,;��b<��LQ���FkӞ�B��ɵ���jp��w��q⍟���)�.��O�y� �e���cx���b�>�]~��V��ٔ�U,��̚/�_��y��xU���LE).=R���k�r�c�e�Q�`�X���u_���WøLt@���P����8�?_JT���Q�!��9�;ٕ��8�د��W����^��y�+���L0��u�7�:fV�F78`v�UQ>��uá�
{3����Lb2�to���*:+=b�(���k��΋�b�ؿ�������N�~��{���̢�=ȩ��"n*�8�I2�����9A��J��Q%�T�[Wq\#��VZ�Gú���7؍ѕ *�`!?�f����ih"��W��B9�WdX��b�P����dݠWX��%+2�����U���֭��X�M2'
�b�S
�K�*K���ާ�Qmٜ�N<�P�HX�B�f�Q�Ѥ����+�Z�-���ܐ�O��+�2�w#"��(aU������Wds��/ڦ7�� %=�y46fP�r�v�8����{;�B|��;y���X�b�zh�΄��W�5=K�q��ˉ��#�I��N����2̜�f��y��(��{�4{�s���C�Md�RՒ`O)�|��>�U�����(�U�|���1u��U�9G��=��\�~B�*N�$[ EX�(����&��з��)U~��O�s��Ga],ot�"b`�;˥��ypj*1�Sјjo>��3E%�1�N<�%��q��6���4��(ɇ�b�բA>[񌝶�V��xT�C� ^��B�����y���`̞�N��־���Z|X�T��_s����)�b��M�ZnR����5�"+:|`���'أ�����~g#dӮW�5y�͵�c���G/qPH�DE�4��Ⱥo2��h]�D�U79�r"�d�.{f�w$�,I��S3i��e�j�]� ;���C��l������սZy�ʩ��Q�!@���$�ꦶ�k�e���y#� 	��n܈{S�u�����E 4��2F�>
l�>��}�ۼ��/�`��?�$��-(vgB�Y�����$%s87`�����S�[�66c��:���R�V7�ut�n�_
�ܡ�uhr�n�^��8gk����^:&r�[8v�[�����0�F`�����pwvR���@��,Y�n�dۮ�U}]�:��t�\�	��kN%\[٥=��k�6�4{}:].<����4!r("G��D���1��Q[7����f�i�lv�"F��
�x#Ϫ$aM����N��*7i@e��n𘩬Q���Yԇ�r�ͯu�
�x�pR�S���2/<Y�qkTt�j��,4�ύ��Ǆ3(�R���Jɑ����h��a��\�VZ��>��T/Χ�
����L�y�]w�K�W{�s>Fػȡ�Q:M@i�<�y�ب�UJ7�9ޏB-���lH�K�|hY��y��#�e)aUɯ3����>�3��t���ϙ�p&�C���ѼV�;4=�N_n!ݨס��[
�#1�~y���V�M�(�U�x��Z��tuMlSfy�ܲ"}���3ח�������УXM]qxk�8q6oU�c��y^�m�`(��7sCbW��,Q�~Dc�2᳛~
޿l��R��k]��	�jȵ��/ށ��l1GTe�Z:�i�_oX��+Y<�"s�3�/�z/���NZ!0ʙ[�8ׯNWL�Ů
dP�W�s���(H�"&+1��3ݴ��@�����A]�6���A?�7oKal�~�15�f)��C/7�J�4et��p��X�������1k��Ջ��1�x�ssԊr�0�eK|5�i��S��F;2n&sOp��(	x�2�0�f�ٕ���4����`K�(���{*f�s�YI)����r4F�^���Η�F��Y7eƊ��x�p�z1 3�Usc����*|T�b<�$}�'�^Ji\�u��"��������=�y�z�8���{��W�3z�&3ҵ�ƅtHضf�(�eМrg��޵�^��3��aۋQ���R.]eBⳊ��,�`��n|�u�+`��zR?m�y	˷�'�J��Qw�'�	A��$n��Šs����>�����-��Z�1A��,ud׳�D
�V"w=�9�
�4~�Α��;�_Wf��1p���rU��"M�y��$;����|�$��ǳ贅���걁������Q���{�� ��@8��1�A�<�B�Ѱ~�>�����x�R}���6u�P����|��]�c*��K�%8��v0R۞�*��f:�1�ĤL�>�%#tyE9>��C�Sj���՜9<�iG���B�a{�(�W-�K1Կg�yO�!z�#�����4'-���e@��N@�Ó1�-��W�Y6�z���:+�ӭ�K���J6�NL,[��1��V�#�1C�=S$�!�ۿ	�9��	ܖ�6T��&NVw�r�Z���Ȟ�'˗s�l� n�J4�T��5��В�v����V��ѓ�zS���l�w�_W�I��Z�#׆(Z;����K�ͫ��'�^f��-)�r�)���������2�j��2�9�3-8#�����r���<E��7@:���;��ԏ`L�\_���[h��W�Sv���4�u�lM.�M�uj���L.�R��^�y�ȗ���
��8C~4����a���Y1Ӝ����3�룵�ڀ�UΊ֣��S����8��������m���d
��E��~q����h�xItȞ�3�L՘+n\+��|�@�i�E{%�/�zu���3���G�Y8!uA�Ax�;�%8�A<p��;���>�mG���O�=���A��S�2���flِ�L�
�t6���d-�ݼ�uzg�-\�2��3�N�J0x���k�<�بQcZ�Z����Cw�W���L1�A��v}N��'C�-�N�����O`E�0�����0���[&ﳉ���=�f6�(��sbI��޳*�u�!%��]o�&vGيw�b�z��r�G��#�mx����l��N���)�R�3�,���==�o�Su7�CW)��0��<��sg��8�=��I�.��^�]�]�V�\�T�#�Kv���:���o�ѵu��������9��=���M�V����,/=���{U�W��i�ؽrkS�X�r'���q*��Ux������^LڰS1i�\��M.ܫewh���F��A�)�z����'/��boz){v������i;�Me��S��/�&��sX���w�L?�2���h�� �������q�|~��h��_>�����zj�;̯B���̥�/��Q����|�׋'��=�^�B�z�#yxG�-�0� o���n���=���dϥm���I��g��{�,=⒛����#9\�wz�6�y�9՘���Q�G�	��I�x���q�d�S����a<�;|sN��##>�ST˭�H�W��5��è`n/a�ު�M��Z��d�^��"��x�uln��Bw?*�~�GGa�W�>�f��痝��~���h�u��Գg=��ad���B�����?{3����6��� ��i��۹�1�2f��u�Q��5pIE.�%KG�e�ا�F�'^g��kQ�n
�=шNE�ج��u���@���q�ۼ�`��q�=�s���s��9:�Mo�ӭ�������
�"U7��tl���������ێ���A6]%��o�c׾ܝ�_�c�GM�P��}j߁9��YY��
��vr����ꉍ�/s����|��ՌM�s�r��ݸ&U��|z8���؞5���ͺW�N`���T��x=������p#�c����N.��d��"k��U��iX�a�"����M]g��;X8r��G@y���rY�� ����+�>@S�x'sP�� A�f����ɖTw�,�ݎ7a�gr�y����"��\���˚q	�v�H��-�Up��2O��'50C;���әC�ܾ��
<�J����nwz��'ʁ�@�k`�9%�9F����� .��ڽg$����E��o�>���K_�M-]뎨��<ș�G$3�����u6i�	��9qc�{U���ٙT� ųSY�+�j{�}�Tt��C5ի�tW�3�1<��1C��c������e�� T���d��
j<���sW�9A��{��8��ˑX�gDσS�O�)�.㒎�1ݶv��?x��Iy*ۭ�8rKc��8b��N��cNC�b��鲘�̽�K����p;)�D!"=}��q��r����c�RGR�|���:�y9���}47�N�➄;T"�Bޏy�^Q�m��v�r���X�G�eJ�+G4���a��;:N��뇈ܠ��LK����E�pL"��fOO�b�k�����X���Q�������d�%�kϺ�k�[�V˯t�+�ޜ�X��ïr�i���ϰU��J��|kFL�>�fiJ�&��Wg��]ޮط.+���ge��Gү�r��0��.5�H�쥖���ԟ�ό�լ��=�b�ݛ�&�R��t��J��ă�/P9�sL\
ꃐnMzy`�~]�egݽvw��QdX�0���\9WwF�	;�C�]���)����T���0���zw6-do�3�V��rV��7L�y�-�	m
�C���BN�Y��
Y.�Kq��"5̭t��0D�	�A��32}{v�t^���&�+�qX���v�D�jf�BϷ(�^��c��\A���ͼ�[�ۇ�}��}�f��o8�/\��~��;�&*�j�q��j�Gu��sj�p��#��(���Bc��*��-�9fa�7�d�b=�"���h���^�����_��{i9�qd��Og�do�o��~�^��}l�Ϫ\>.�# �~�Lè�sK�(��i��G�\>"�F�����.$�{<�W4��S7�����0��m��#;������=�s�F.w=b�EfIyֲ���#D����}�Zؼɔ}f�9]�ĲIF2n�V��d�U:μ�&���x"P��f{�I� ��9#p�}-�yc������n�����7w�_�>pD*�ԍ�_�r�c�v�����xfG|�v-��Q�A������j+���ԕqJ�Q�Wӗ@D����MY�+�lLzp�[���������ޏ2wrbS��+����|���k�x����q4�)�r�]��0�2�<
��.�w#^�+�h_)J���~����W�}��!낛4�����vR��s��i���¯�·�Z��6A�77J��i�/ׯO�w��up��l��P�]����o)U��#�h��g,�^�@�y�8m�=���A��]E���z�TꝪ�w��.'6N�ӊ���BD�i���B]�̈́�@Zز9��)Tb��Ü��=�]$�{{0a��s���ͻ�"�B�{�6`�E$Dk���9��V�����n�8�LO�h'[�^�� Ix���ޥ�`�˽�j?�\��#��w�W�}�fd�V�~v����)����r�hJ�d	s_I�Sş}KՌ����eB�Zg�\73�����ݟLs}����yJ��46�zh����}� 葯^0�e1�D��Tꗔ�C�7��r��c�_\n$޼�,({�����P��sz�k�s���G<��YI����ٯW��n���	�O0�`���t���{���_e�����6����lG�&�U�N��%8GneeG\u���w�5�6槟-~*g1l�B��≊�v:�]gUܮ�RT�*J�s`{��R0��|�wq �L>�����ge�L�� 򍯩K�zCZ7��e�Od���%�"������z�R�(ݐpd��I�T�>Wj�n�3KG5�^cx�Y6s%D�ڰ"FZVe�;z���0�k�Y]qәp��3��gY���}Q1������ͥT9O� Č���ͮ�}���S0�8��v���;X6�s$�]f���v
�6��߷�8��"�h�S�:tԭu�$��c%�����m��n��7g�c-L4Ӛ�����(HP��oc��UΧ{��ct�{�����c,����\����h���z�ߜ�k�[gtQ����--�¬=�qI�T�يJ
�0\[�(X��hjH���w��/�[,Ù
�3x��V�P��%�΍�.�ǭ`�}3�p���7_��]�N)�]z��V�e4oI�N�	BY6�d)��U�� �WLt����=Y{� j��vj�4
������7�c#X]Pwx�AsA�롞
� f�KK��l37�\�rQ���P��S�nz��(���C��q�=J�r���"�*O�I�#�]q�%'��d�{Z�ο!w^+g�sY�v�Ps&��"��z{'z�+�w<=FL;T��yZ�ܡ��YYx��ݠ��ݺ��y�u�5�����(R���
m4+\�c.��\J�{�D�_�t)����1����se?z���&-I�~:��#�P�,Բ��������}{e���D˂ߖ\�3W��5=��KI�1�$�~�}Eւ�m��_n{;2
2#7)�E�Q��գ��)ݵ0�(A�-۩��:ю���o�AF^.4B1�gU^�V�	�
d��y)Dǲ[~/5�^%���V=(�jfǊ����NI��ol�UW"��]��܄��>�U�|}�4zq�^{���3"E\c\d��0��7r����9�fɍ.汉W�����m�Us\_�3��{�Y�L^;Z����ո�MJ5
r�N�5i�rH�1��lLE��ef�sr�]���0��/�C5��%���U�}uW��	ۂ�(���m��� ]�ʓ��ul͐�J�IG���[m%
�;6����/C���\DE��Nx�]�_Vn����mO��IXWn^zڰ��=l�=�ϢB\�gd�bImX��w+�^��qZJ#HJ<B�u���^���$�\"�'��+��6�h��9��\\`�osq�i���ڗ~�N{�U���4�q�!y�ʝ��gJ�쫥[Jy��#��[�,����D���L%��DY	B�u޾[�ל���^�k�����2�t��/�,N�l�Ҿu�U�������fϺ�P�beh��n�r6Q���gz��v5��ŉBL�s���?[�q������>3Y��Bw�k���$�8K��733[x^����)Aewu6���3gz���KhS����uuI\�ک�t�AE�$�l�$���+!/ռ`�}��˽����<%D(�G8��(�"",�V�������PȂZ���.����{��*svR����˥(B[�pU�X��"�#�����ӶnC&��������]t����u�b�1ե2��kY�gh8{+�&�#e�E;3޼W�����(�U�>�+裊2U3-削fEy
�%{�	v���f��/��w	�N��L}v��gbx�7k�8�M+%]�^�ܹ)�0�#��v��.��)���'eH�ep����)e�Wl�&��1��x����[È�멡$����r}Qt�����<����ZE�)��5�3�,(���R�^�]N��l��^/����:}�:�S�p�E�׵�q��m8���]��,��=���Bӎ��1��~[�I�+���d�mUUg\��SF�!a��r3S���R�ʭ�ke�h���-	�?\�1�"�(����l(�ĶM�7[�ܙ���k�,��a��7�n;���R��]�Z��9-��Y�@�5� �G&
̝FS�2���!"�2��f�mlM�JmՊnL]��g�(�BqZ��
ft��Փg����ά�۝��g6�����`ɘùzd���V�E�n������ս�c�7����k��{���g���c��;���N<M�%���
q��g{R�Jѣh��o�.���u �l�f���WU�M���%����&��ժnSK���_7���ݹ�#�S��B�M�����yv�!�v�&C� �j̫���79��W"(p�mH����)f�9w�&��m�X�T���""���Q��uu�����A�p��,�u��f�>o��fd����=�gj�a�l�Pv,wu.���;R�ݕ��7��iV�̀q0���A9,j���*f�k<qnw\[@��7�nݥ�.�l�K���+�ۉ���ݥ�����B�JQ���klr¯��k9�S
u�7�IV���,�	}o�e�v������X�;+e��t&���H
B#W��:q1W!�!��vS��	
ї�a��.��z�Ӊ��6,j�Ѹﻓ͐cԲm���U����	0m����>���۹�]�g�vl-�^ �.���c�^6�/�K^j����0�[���p�_L
���m:w�	��:����~�՛.L<M ����;��{;N�V�U��h9�Zk�k�{�Z��ǪN�*C�87+ns՝ !ٗ��*��T�enK2���UD���4��&J����iCc9�}���G��D���^��;mR��늩�~�������A�#�T��M7/P=�u@]WFɶl���YU3>�WS^���B
=/6}UWW�Y����n��\"�TT�{L^����ܪ�`L.���K��ו2��@�n�kd{�_V�V���eb�=~�A@y6���L�7ںF����Y��fe:^�?
�n���K�;�����P<(����7t%�'�7ld�5$:�Y���:����Ľ+Ӑ��U�K����jN��Ɨ�����7x4��ϔG����{l��m�N��b⃅'v�4��A𲣅ϩ��#,B`����(��K}#Lԍ��nm[��V@~�̶J~}6����ũ�$���[�'/p��dm+�_3k|(Pb������9������h{S��r7����+g��-9�`� VGLzq�
�]$��3q��#��G���"9�����,f�����c�r���͝5��
�b`*��:h����hV�S}c{BF�_��/b�+��]�:i�ݼnL���1��͞���'������^�W���M�z{q���#$�ӏ{�t��2g"�R.󔤄�C�иg7�(��U0����#�Ny7k��3>cj��{>�ʽȻ���G��l靉a�-�`���=��>��n�،�ћ������=V�/^+4Dp�%�i���K��ꍈ7� �;E޻�*;�ܣ{/zf�}��N�**���=J\����^{��*[��@�m��]Ѱ(�N�G�1P7&W��W���˗�ݚ� <$t����%W{&�6ţ�)�h�v/���:*�N�$��z,W��eu(Ѹ�Nh���X��G���F�0�>��[��#�^�r��p���\>�X�Fb��+�����;1�hU���3�R��鑛����v-t.:�Gn�>�	gn�.�N�X��l�9�ht�.�?Q��쯾`�ҏ���F�!�,�����3t�s��o���G:3���B5JG/H�)��`-�ީ��י��9���ʬ�h�Cc�����e���6��}	�!�˸�5+��i6b��l�D�^�;9SN_Q� (����=�b��L�c���l;��}��N�8�~C�����w�w{�dr�[��Z&X�:�K�D]�v����T�ܙz:�:��]3F��V�O7���L��/{���� ���n�s�.蝾b`y�
ox�_��3���#��S0�J�]h�Y�\%_<�C/�{$��u��Y��Z6���k�p��ɡ՛`�ڶ� �^�{Z�q^�w��F�Ɲ�E���@�`�"qe���l{�C�Q��E^5�;�s�}�A����N�|��5},�ѽ�P\���'��a��le�M���zM�b�*Tk\3,��c2�	�ی4����'=Ҥ%޵���]�;�"�*X�2�x<��6<@[jhP���2��x=t�1��^/f��_��a�����ݾ���yzDd���ny�AB�BbL#7Ȳ<����ԟwEBi5f�����]�(���g8*ɗ��l��*gՊ������aV�e�m8��޽�I�W{���33n^Y�A^f�w.ڕ��S���0c��t�̌It�/�Ѻ�'L��zM̀��t\n�F]M�Y�-�=��o�8=XN��8�=��ƧL��5�޳m�v���G��f�ϒ]}�� �P|[�joAZ��O�_X�����
<���pZ�u��Ҍ)��q~;�u���k��>,ˉ�dU��3�1w�"ť�������Ir6aO��ǘ3��(���19�<��Ɔ-�Ln�r����*)���O�k�i��Jobs�I�Kk<R��8����<��0Яk��Xq8D.ʷb��wpQTjL����Y��b�޶T�bu��M�Z�s^T��R�R�u�� &܂��	oS7��l�Pfu���9�q�{;���K�ы8��\m�:����a�+�7����Ǎ$��d�P�4x}��1zyHY�L�������i�P.�tq�޾�@�Lt����l{�}�w�*��/�"rj3ᒃ{��`�y?�@=��\=��Y��J��p߽S���T���t��MB��;�`���Q��Q�PA���%�>��JV�#ٍPCs�!Y�o)��s�ɛ�>�D��~���{�[})��3����i:50�>�#^�03ҽ��Eūw�ړ�Y����h[�N��K~�R槲��`C~�W+�:$d��h�A�r�pW�-@j�y7�{�'諭��*�oў� ,�^��Rk��{.2��f�8VO�M_���p��v]
Ž�nb�F���q<pU��W`PTD�B� f���G�6�
�qGi���
P�Y�WWu��<��r�Ɇ�ue���Y�;*��<�K+N�&8GN�H�f�s'������$�.�A@�RY�5ڕ\�f��#&z�T2��L>�~ÓYi>g�	��3~5���������3�y��/_�/�˱�ti�t��cS�j<r����O����rDN�=
]l^Y�ih�?u��h�s�o�[��n�������aǵ�Do4��;��,{CL�]��^��V:y��wNӖԬ��c7�%���uK*��Ф7�h<�4ުko����[Z�:��JB�WZY�J���s�Z��*id8��.�uL�q��;���Ov��ϔy:��=u���eGf*�r����V�����ݜnes��&mO�;�&1����2�>ߏz��@���F�\qj����<=�*�FǕ��d�`�]E\?S��k���cyGC]�\d�.��_��7c/�<C�f��b�A��w�eƉ�z�h��?O��{�uҟN�'�YǏ��0g��E@Y���A�g_I^LI�QU��U�!T!�Nj;y���W����#{Bђ�r��b��R5v�דǦ�
�p4�9Q�IG'�nR�n��	��#���g��l�%T�u�����]�����ډ{=&wؒ{��ݼOZY~ٹ*��K4R��`j(ZۀIe�ݣ�Jն�MǊ���J�{X+80�4d��?Tp�n�(_�MyV���K�%���0YL�����1 ����Y���!@��$s�Y�Ms�������a0PPg�����ZA�&��L�	��%����p��#��؊�3\�M%r2��Ds�Ԣ`�F�Ύ��5m�����X+�يmt��ז��U����b�a��;����i�ʑn���Z�ؿt{�ζ1r�#Y���g��&Ns�h�ڽ]������H�;�RJ�u:���h��٤;��e�M5�!�i8�����\g((�v�#]ҹmBi�v�RF��r<�G��<2��,f	�6r��,����l��Y���RNeGP+��t�2L�]Ҭ|nP���/�D�����f9B�ʌ���O�1�q1���;����!L�zR��f.���}����-�҃�n)���G�)���[�`(<7h�+��i
����%|e������N�=���ק/LR�qu�x �!/!	�?z����e�s�2TUO���QF6��j�>u�k�V��w��a�^�������u��d�F������6|`;�n��h�tm93^���^��㍁Ug�ELq�^�V�W�哑�����}f�Q;�a���5�BNE�{qh�8[�M}�����������#I�k8͉H����b�Oj+n��\�i��"cH]�H�����@��c����O�8�\�t��My*��+���>��,Y��f����W!�;��=��Y��+[ 6�v/�>�v��}�#c�}�enuKn
/-�Gdj�w�S�����i��H��
[�u0.�d�J[��;6w43jY�u��z4�8֏&���e�0T�nR&+����YK�,ʇ�I��J���"6�J<�\O4C�juV�Uy*�Em�R��H$D��xI��:��$��/���lk���p\�����u�smU�W:��gh�x�_$,>X��a��>�u��ֺAÊ�G���qd]v���Y���ȴ����
��±+)d8yW�.�^X��6s���8?L1���0���mT��56s��{ك�6}$�?]��s�Z�Z݀<6���i�X��˺UՔ���;�߲���w�$�^����C*`��>=Q�,5��C��{�*p�Z{�^qQU1�w���Wa���$�QsQ��f�������}w��p�^��t���+<�z��E��I��\ �.�¯Hr�?C�� `����]z��*	����V�-�t�����]_X^�AK�Q$r!�%�Z��@��%�/�s��
'�5Z�p�3���0̼�yj�]�2l�Q�h�lMF�Յ��E@�����vا���ݿ2���c�Y�q�ߎ{�DrQ�j�ߤ��O'Z=��T��)��ۊ�XX��a㫧�2�7�Nщ��JzqñϽ�mz ��H(�Ձ�M!xc��8�t8�]z/o��_n]Zu7��R���Ռ�T�7~^��l܎�^�wؼ�U94�d2���ڈ�FѸ�o�wy EⅤI>�F
�f+D���c��|�e�6^�ѹˑ�.��oxP{����rD�CvY������Ë��|�a=�*�f����%��:�Q�p���
�(��;B'�V�L��r�������,7�"7),Șd�W��2ƕM���陧rͪ
.yKD���r��h��Jj���	�[�����Q�6h���rXY����x	�P�|�[DX����ȫ� �!���
��%�b�n)���BU�ȬAo��_}t��4]�\����#�+�Wy�[���
�ߨ�n�S,]�
5lve��<
�Z��1���х�̬멝���z��/��2S������)���y0�k8d&�n�U�/��P���#N���s�L�^q��R|#�X�Į��^1�H�SD��~BA�+<�5��q�9W���m��/\�lvI��Kw~�{�@�"R�q�/Έ�y�o�㻵9	ˢ�kw}������Y��M���?�+!�r18��_\L�mj��
��/�t�٩ pR�-��&'z���V�����~���{j������VVؐ���.�'m�΀�#�lT10s%<^6��,^,�۱6н�'i�	h!�N�:M���v�aQ��Mk����Oy����T�(O7.p�"�3c�a͆x�ŭ���zX�J�Q��N����Z��0v�B��u�~�Uޖ�8Uu�{p�|��޸�mN�n<��v�7	�/ڑ�����v��mZS��B��S��K���?��H�~�1.]d��^4� ���o^����� ��2�����ϊ�r�̻B��j��3O89֋��h��n���v�SF��S��:$��kAu���v�Rmw1����T���6�]څnrԗl�p���������C��.���T��X�ū\ �F�¹�r���H���������;���-�{y�'�{�.����Ta�߮�,��]�����2Ϭ����Ik��1w*��F;8�N�~oȀ�q����;/�/��Dz<&�3����y��M���K՟l!E���<�+��>�.��F���q�q���1Ǥ/	��?vw�qVc+Dc��T���}.ћ���Ӽ��a�8F�Hp���:\��x��j�ӕk�Ջ���`1 �xB���o-*#;�dP�m�'�#|�ړ�l��^��O�<�< �
�FG6 ?U�)�S�/@�<O*F�GOE ZZ�=�}FJ7�bQ�ƺ�z��{<n�(�t0�X�X3�\J��z���Uh�bSS�=Y��^�y�����Ǹ�UU�^�>0D��S%���+����<}�E8��n}}Iɣ�L^�(%&c���`����o���z�ϱ��ǎyP�֨d,�N��BV��ǝm�1D�V������D�,N�֏��J�1,���321�[7�y��2�q
��l��-j��0B�46}�h��O$u�2s��;�U���޿=�^C¼AQ5#�.M�����n���!3���[}ի[;�);ky.��J���B�k/1r�YW�Ծ0C��;�@�)mf���^Xu���5�� ��C��Xo[���j�)�;�_L���{;g@:�X�Һ�W���oWn��PQ'�C���'H=EV~����ŵ{�4aS��fZ׿R!GG5�6����[ur�d���&|z�z��ŝ�h_
��F���@fVĭ"w-��B�w��^\ׇD˼�PBjD�!����Cڟ3h��0[����3�D���Vn1�cH��4@�`�uSS��(R�8���B��0z�=r.v��Jm�8/®���0�/�o�P�ݝ��zo�c�O�$GR�����-Ѩ�z��T,���Y3ΐ�^9,;:~x��;Edq錉�ǨN�K��T�hW��m�03'�JQp��5P�A��{X3��uxw�`���Q�5a�D�q��$'���t^�Y��L�M�#;��ҾDm�U��U7��\u����zԻ��3gfZ���s\�㎥�?�6s�៿�
�
�b�_SQ���4�^W0l%1����Z���M�N�|�²����Bc����=�5M�=����qQ88����=Sܱt��Q=��f�_�î��%ݦ�@�ï���u�D�Af���7�}�yyud�&�q��I��7z�=IZ��u>cb7;�O�q@ur��(���*��.BB[{�
��W��A�Զ5\$
�b�7���s�Mfj�Im`��QQ�a�B �N��n[z4��@��΀�[�2^�s����o(��d�3?q�[������t��U���B����Q��f�/C�̬�|���q�f!Y��ST��v{�]z�6�hDDD^���\�%��O��+�t�����kd�*�kn���!D�	\�+^˜���U�^�_RS��E�X!Td���Hu;b�e�`�N�+����) E�>�R�>ꜛ�ɪ�9؅D(�����~s�<���2)�U�N��$MJ�:&b�Y�)V�P����\@�}���&�]Wӣ�eӵNM���z����KzA������jI�(��j�)V��g��O*ԠQ	%V�to��N�[Z#��^5�B��<+�h��}N��T(u�����Q�����ʶ��UiA���4u^`�[x]fj�����p4�Z�n<�/6�9ʛ����J�N��uUU�*��WfV'��4�c����6�f��,�8-
q�ZS]~ܺ���7%DN�-�]`u}�[�##�n���󷵸:��_c�����}6��[;�z��}r�8�(Spo�_��/1VI��]��U*���=�{�Nk2��0�	qG�yŜ.!aǛ�|X���3�d�&*���YVЀ��+�-��ź����H��sU{>8�4
Ƹ��eݓ��[�w������U�VNń&�q79�ˡV^��Vf�Tn3ԭ������b��
��WKʗw4���/�vH0��]E�0h�/�S�Q��9p�B�^����� ���E���������6Ḷ̌��$��M�s�Sۅ.�r�4j�Y%��PW	�}�! �Q�L��y����9�F��F��ќ�5dKw:5^|�J�_i�����\̐�(G^SFA�U��(�߬؛'&�R�-Q����Yd�A�s��
�˺�"��N��3}w-��k��7��r����s�3q9�X2�X�Ir+C�%���&��؂g������zF֑F�
R�*ɳ�&65�,+ݑ�4�����k�;��kL�)Pb�4�u�w���Mk�b�����8Zyk�^��t4��Ҧ���`�7+��m��	0ڴC]�f�1S�T��@��XB1�f]���2˻���	�Das0)�!��+*��2��kk;23a���=d,�<:�0qӛ�������ϪBBz�����s�I!ޛ�35�v���`�0��6&bN�Ԗ�Z�+�Ӊ�vvK��ήM���I\�0*V;�����fwp�YKK��pG`������Z��̳;�/xYٻǤ�K�n˶o�:w�1=�G;y �]C4�Ε�?�GG�:�g����3ī��	��f2��� QjӰ�$�6�A�]#T]`��.�ɻ�Z�~��!�ӹp�S�V��L]	��&p���GHY�x�C��왈�m>��x7�;Vw@���K�yg:���7+����x�(�s��*�P��돆eL���ri�V�]ֳRJ/�:YyՄ^�.=ѽ[�q~�<��-���ө��u�QʫөXWY� q|/��Z�~�:�r3C��p姨�W�+��ޖq�@�!=x/��Օ�Y�* e��W6�K��Z�������D���Lh�&�grۅ���ۤ1D�@���R`Ҭ�W=�K'r�/���a������E��Ntɕ.PW:�7rY믤�w|b"ΑyK�|�K7}� [�
3�+�{�x���~Q�7Ce|/�@sG4�S��ض�l�6�U�Fd�}�L�޻�)���vƩ����m���{32/f Ю'�r<o��%X�%r����9����I���7����,�_��N}\��Mo�V��a�?K���A�:3b��ܣ�2���f=ν��3`�W�0��W��j�Y;/;��`A�ͳ7��nٖ�7���"��!e�!��!N-�go�ؼ�v���<%F*gxc$��T���6�U��2�=V�@f�ǹ��mG�G�b�}�����`���#�&(��� _�����7�v���Z�;�D�gwJӉo��Ƿ4G#Yc:<��G6<�TRvc�Eϗ,^�$�U�������T(�ΨE���s@�Vǎ�~T�Ka��9(�V�k����h�\e������&4���-(����UqQ}o'~��|� mq�b�X�9�`�u[u-gnk�i��q���'o2���1�����iB���(�I�~u�x�g=WY�po>ޡy�:��tl��TN^��*L۵�����ZEq�b�W^��r��-���X�[��bz^��&S��9�Y��J���z���3Y��#� �zR�_��g�eCÎ���0zt�P�
�+��	ɍJU�]
ߨ�z'��Ӳ��9�����~ꚶSQ��N���Ɂ\vf�M�ͮ�wt��6�o���g��WsU+�>2C
k��ò�Tk?[�;9�X�%2���ю�Fb�������}��!����g�bt/C��uZ��9��FO�ĉj���h����A��kË��u��h_L}���[r�]
�S���c�[��y�2��o>��R��w��v��aW-΁`Nu:�g�'��ub��G�!��^o����3`}j������+OZ�v4�vf&��^�Y��ғVt�{9��C�l}��$ٰ�E~o���ԗ�o��=�����^C;���E��
'�/z��g͞�a_| 1|���n�j3By[�j���E�N���3�'�N-���+&��'�f^�`K����	�_�E9cÈ�(`�2T�N�mk�� �aF?�s�>����AQ�i����3�E�Ga���yKu�#yвOir���}�zʙ�7Q8]�sI��l��|�,R3Jh<�,ա-��z{sCj�lp֛�y��qm����6]D1-�4ɀp����M�q�9�
�1K�ݲ�]������xA�]��q��7����O�nV~+ZaWٗ��n���}/�({�Q�g��'o2���*�L�^��h��g��9��������-(�sOndt���O���]��b��s
C�ۊ�������iy۾�����ΌR�rz|+�OXoA�C��y+0���p���Bzdm��@��F��&%���UġÀqF)��������(A^ݬ69Y�} �l�T�%x�Q�|���MG�6�p�x�;#q]+.y^���(p�2���Y;0lj�_1йWD�Ӥ�r4 ��8D���4pW��~C/�՞��dn�&�G=���ȵ���ԩ�ZOo��.1��r.*�U�Q�SJ-j���!�ne����;�GE��.;����P@�r\�s|�� ����LLj[���'7�>'{k�ȣZ�z3R�G�g��Dz)�Bh^���U�y�8qj�����=��9��S�#���~�v����
�jv������z(ݸ��M>�3G�~�Z�Et$�9�34�ZR�܋��6�;\HYQr�]�[��P�y�����nvFu# � o�23. ˘n�}
�5.:�v��6��K����y�.�}j�\ͅ1K���)K�9S't�FvZqr�N�'�1ی����P�ͩvRk���@���s�ͺ��/����b��=���1S��Ţ�j�u����!��q���V��`��ؔj��1ݽ���W��S�QD�:�����R��'�f�kbc��^�~%t��4��jp�v�a:�Kָ��X�V�/x�R�R��>�s1Y:m�b��67h�� ��A�Yn�o��	'	�e7�&����-h�/.F����F�ӂ��y�mH��_k���l�F�U�Z�/<��QC��J�7�-�93�
jQ���FF1��sݗ
oJ�ʒ�zWHO@�ΧJ˿E~���V,��ć�l����7'u�Ի��i�/X|w��m����&�כ�/5���V˭��r�����6s�w3lw(ֳ�&���C!Pwn��F���컜*]�!�74T�7�h��Λ)�=����u����>�ng�t3%ҭ��*}�"cٚY=E[��������O�t]]tC�W�$BZ�I;_:).��p���Y��L�Y:���q*����?]Ei7p}��������;;c)a���)�,��b�J,`�K9��`E҅��Tyws��*v�DXp.F�a�2@:��$�v;}�pǱӌ
����_X��q��2f���\�L�kc8ƯL�kؽ���}d}Q���9�:9��v��UI��uT������+���ⱺ[I��N3Eh
~�� �tb�Ò��;�5�7�Ooe��҆�+�']�+xS/"�S0tY�Y�{���_��t�6��2��R�Ɋ���3啥1\jM��`e2ܴk�n'BTC��<T#��!��@�.N�If	s}��#�f:_w�:W}�,���^����6���hk{�R���;(�q��L�/8߇u�Rs���k�B�G����thu\� +H�ݗ��Ŝ/m����;�}\�8ol[ʝ}��ϖ�!O�Qos6�kxS��2�9Uu�;:}�a$�������]Kr���W>�Q�� ���8&��Wq��L��=aJ�Sl�|�S]`�׶k���w(q�.q��ѽ�öey)��##� �ƻ�Ց^�f�2�{�6<�Z�x}���軘v������a��Ϥ�b:�[Qr�'���`�י�>� ���t�� 9���T��3x��1G�c|�fW�0�o�=Q�yQ��(�ú�&��	�L��1�����ǆ@�[�nI�p6��3��
��Lʚ㽓�b��]�ԴD��;�?ln�d�H㋯m��d��ʝxl�y>��÷B&c���6}B�:��[���� s�9�13��V������0�V��%T��MBؼc��֥l8�iפ\�D!�I�kr�|�=M�:��P&(^4��N�F����>�	�y\%��k9U��c���f�&m��a��/qt��K�ߝ�C��EC�A�ז!|��㱜�T< �����{�c)uĴ̢�n��'�o�w"�;c^j}o�M��I%�k^�V\U �n�E���I'��s�=⾿,���7�oƨ�v���ܵI�gٰ��Ry���|�SN��n䉅�J㢏C��ԣд{�Ѻ�[%��H�?U�]�s5�;��g
��*B�"����V z�_@Ǌ��ԅ]dҍ��q#`���W��G�b����?{��3�Ztgѭ�y/�7
wu���gv�����n�r���w�ʄ��ژ�{^�ϑ���k.�d�k+���gù�oB��^�ۇt?X*<2�y�i��^�r`$C�Q���=^�ȤǯP��_��ٞ�+M��'�#�=�g~Q��1�#��$�
�:@���pt�.�A��3(�dw�m�l�S_�K�I	�d�];��_��ȏh�"���2�d�4Nv��͗�Zn��7�Jo��]��3�QV~���3B+��sb�Dǂ�#I��/�=0"c�M�A��ӹ��^	�=̽��j���4�L�T;g��/����9�}k��wOŸ���r��l��W[����ϥf�q��Oލ�w�nH�b�x�)����z�2=��>9���W}ܯ�-���LNJ�x8ymo��$%~�=�X�4�s%��	�[E�̭�X�:dh�9i'�j�o6�m��!��
�iy[��+�5oa궲�W-�A���_�ʼ\/�ԑ�Es��N!�j̣2��7 �YM�R�-���̼i�:%�p؎6��"�e��7/u/�����x���w���{��1�w����}�hdvB&W�'4����P5#���y�OL!� b8�"7j��8ߝ�k��~ZPC�Dй�«oT�{�2W����G��������c������_'��w���.���}:� ը�P��Zy��t֍�0��%YgqyP���*��c�8����|Lׯ�bF���U�L�"U-���Ɍ���R�蚀��Ƙ�|�C��a�E�\�����=w���q�~���y�"�#L<�r�(��\O;��N���Q�v<�yH ��p�#&�<����3:J�2�8c�)�v2��Q�Y(�0�V�vܬ|E��6"���� 4���VW_���5N[������阺��Κ���uh���R����-�l
�97uʯ�%����Q��c�j����7�G���ɉO!���gl�`�+v���rP�'J֭}�qn�8��a��oI��qdf;2~��:�A�VfDok���G����ƫ8�bB���=<F��`U����;Ѩ+^�x:�a䑄`VE��T��R��"�~ޭN�(�o��@Ϋ���+�T|��t^�`�����D�}]A
8�-tG���"�1OWMw����xO���9(��W��ro7/;�qx6��m�46�d�]+8�NW�]�����5�;ʒ�U,�h�n���sBw)�i��xe�vb�&$��jh{
s�A�!-�OP��������+�dr��1�y�7��n�'J�[����}��V�� �����z�Tx�U��vf���D�I�˚���A?�b~"�;��**;Փl[Ⱦ1��I���=3�xxa���_�Ce�9����6�m�g}4}.z�/T���7ܕ��e����XA��Y��L^>����P��(*���$%��뜚�y��B��g��k�Z/�l��TNv���ʄ����VFEQ���]�2�l�^���ZOZ;p >x�H�ͻ��e	-��8�����!k ?J�"�5���z�V���=ciԫ�ͻK��s�D�d���<��	�m������˱�L��檕�������B�W�@���
uB�etM�1J��ِ���4�_��M�9#�C8�n:rs��ќq���x�U7�tl�Kٴm��s�P'g�Ǡ\��	x@V����fTvr�����Sfժ~������Be��B��F,>��?P�z^)��Ly0ӑV��5��:�T��U�4:�`���U,�\te�Bbx9|�]��������]�:�YO��H�J�c��HER��$U�m��1�ve�)X�\}*؀enuk��蔯�g4�9ٖ��*m��խ�gW_u��{u��Ĳn���t¸k���<�Eluڬ�9H%��f ��^ũ*v�=�"��B=o*:{��E�y��W`��E�X~!�-�2�C�Hy�c䳦��i�9u���Q��!�b�v�g����JP��͑G���_����@��a\>�p��TFk�13ѵ9<WD�˸����Y�|�5�����X�*��Θ��nB1��<fNa)hou'e�!�y��z�^n���M��WK�ڵ��<�k$f�~��`ϲE=�s��޿���9�*�!Y���Nk��>xU"���HY=���' �FD.��~��j�d��M��C����pX ���VWG,�4rֱs�9�yn�c/��E�< a3פB�]!��:~ފ���mw�.�Ѿ; ,$�3#�AF6k��S>�<Xvf=��P�M�e�X{�lM��Qn���p{$.
N�;F:�����A(��}Gr�D��Q��L�͖�"�Q�uƢZ��mN�^�����a�҆wo�������c�*4-�u��8�ˣW�Kc�|>�kl��s�RS73��&�A�FL�aqZq��5����Mh��o+2ue�z1�rv��εBoaٽ��y8Q�b@�+ں��V�:\yW�����l'�Xb'rs7V��p��&��j'��X9�hA��jФ:tt�\j����]q�����I�F���,;���u�n������Ɖv 0�w�����9�J~����|�O�m��8�����E���q~���Bc����!ᘮ�q̏�4ñ���˥��J�nT�z"�!R��]}t��3[=�@�xjK��Bk7�,ݶ�SB���/qW�$n��Ͻ|�ڼlbtl�$���o1v�D��dj�ϯi�Ԏ�'�,�%��ߌ*��s�ص�
 )�s�i��Js��U�1b��@���i�lz���~��d����%�1��y���0���gS��V��T��Uu9��9���G��F�F���ȹP22��@L������w��v~�������xO��S��Ĺ\��7�����]o��!_<�VG}�/gvFř�~^�^�v=lu�i����%��7�^EV���^yh����FO�4�/�ػ��l��6��60bR�X�@�O��3�<\�q��(��g�#�Fc��F(�>�?\P�T�P>�����'r5c���+if w�p���ŧ%P�9Sf6�D�N��AvcT5�9cȞO)��������|�IC��կV���5���:�gU^WeK�ʡ��7��۶æ��yπ]9[���T����]<�]�"�0�ZgIN���LtVoxu�깺zF-ތ��d儦�(��S׮�V�>Y���%�����.0�Ӻ���E�)��C���H�8�g�.�k��镼�^�����<D��#^-,&��:�c�N:S�vE�e%��܉Nܤ�D0U�|g1�m���. T/���1����o���0�V;��̊�r�����h�%j�W.��}���.h�<�]X�������f�l7�bôX6����F~U.c��sqK\��:�� �S�0"|���S����oT]Q��N��Vd�+a�AӼ�
����!��]�X�;ww��{U��H��vU~��6�/A�l���]�)�Y6�T>����%�⡊�*�6�%WOo4�:��LK#Q�Qj`�t�5=�2E�$�aRL����{:�1b]����~`��H�j�7M+�z�#��-�����o�o�4�N�J��
�y�(DU����Ҷ��$� �� ��� Y��NS��+M#Q3H)E�OP��[O��Z��Fv���̇	�+��iwp��Vk�V��JX��An���������f��]�W�>�.���_}�a ,e�b�;"q����E��éK��m�E����3<���j��I�sQ�������A�䯎.�n���u)&v�U���Wj�3�s.����v����-��^��*��N�z�:�_*�3��É���"���/b�^�(X�����D\�VU&�NV�AL�p�"*��̝յ����c������b����*�E��l��I�y̝*����S�2q�$�y�왲`�ܫ�j���\"���]*��A-n�����]�Y�e�+%gq��&Lc�e�wt��q�݁��ɘ�.�P�ȨK�sw��Ġ"3��L.R�ƍ�`���Uu�D{����u����������w�����j�il���M�V�Ƌɒ�)C�Xcd�t�&�Q�G	*��C5�2����[n����Jcm���:I�v�@DR�X�֯xS.$F�ƮMP4 �Ȱ���WԢy�O0��W���F�k���jn�M"EC�,^%g�˳
~�'�`_��V���G��| ��s��������'n�ע_RN��M���b����4V��1��Vc��;Yww|��X�R��mޙ��=;F��������V����ՏNu.y�z��Cl�]mE�v��v3O�b����7� ���Z�t"jU[+w)Bİ7FJ�`�&:�ƍ��r+�xQ���j��j.�lq�O�4b0̰�_^\O��nV��)bf��ۅ-p�pƄj�f⮃2�kCe<uA�Jy �YsŀAwQ�1j��[���՚+bp�Ke��5f��!o�h�ێ��V%����9�mp�l��������N$d�2#���Ywj���UwN���[�!�'N�T#��s�t[k$ג�J|p<��0ò�X���9�^���t=֬���N�O�ו&�C��)_(��B�V�D��LMg�菣�'د۞��q����8�[<��wC�2��`�=9�(ns��G<Q�u�vk/Q����CN*���ۇC��9�#����5av��(~y-�������W�ya{��Q�;�f�+�-{	���]F+�N ���eҳe�7���Hh��,��ꨔ	X��Lzw�`������=3
��BB�q��黍�9CY�+��fd��k|+���|=�~�̒wD�:�6�ڕB���5�-�G�k���(Q�ھO�QN��;�x��w�/{(Q�i�?�
(<�4l��~�p=F��K40� ޤ���� :np8�.�h+nV��Q�a˜�ϰmƛ᧚�7�
�e^?rQ��Jg�.J���C�{y��]�Y���'�{r{+l�=i�r*:;�,G=���¯�{�y�|�
�z���?`�U���1�9%�u�qֳ��?@�5�=*E��i��:XZ5��?�I�l�q�29Lp�r�'��o�//ЗU��"c-`�X\����n��-J���L��rL'}�b��<2����!��+��O=���ԙaňƩ�p���b<q_[F��o=�h���D���9�_�E�����\����}���f�ؔ�8�~�3�1K��N��V?�W��l	�&�ҖW��+ݤ����zhe��k�%����L,����!�cWN{�L#g��@I�-5Vv����̬oo�v=n�T�g8cw��ȤάRc�o��8�C|���X�<ݱ�d��u���*���Qp���������v�q����aOg����KEY�Tߩ����{2l�����>u=�ËZclLp����s"/�_�b:��p�n��;}~�qP�]�6�����y�d��ڬ,�WS���Y++"	Tٽ��k2��5���u_Lp���b�=gx{K�%k�a}>��qt�W�a���Cn#��	ʺ(J��_o�1��#5�d��c�VmU��k�,��z5� �_Ӣ	��ח����Bw'�aX#�����5q��LP�����v���ﭻsNZk�~�6��:��}��1��)H�z�f��lh.����Ny��ͩ���Uҷ5F��F&�ѵ����<Z���g��Mʎ�k�={s-~�#�p�i��rvب�5ې��+F��ˬ�O<��1Ռt���'"�}��f�)��І���8>w���Ǻv+Ӟ����1EĿ֖F��z`���(�+<�X����+���y��n�67�:8��f����-ʐ}�Μ!�2p:o�kZY,� A�lՅ�jD���G��t���e(����xu�T��E���,^7� �xY��Ì,	2���y����͋�aw��h��]Ѣ:��X�=GhU�1��8Gy;����_7u�
\2փA���k�8ٴƕ7��S2�"�M��<ə&hXFnmt}�N�J^X�pu����P�T0�E�Z�cjE���wy%%��ƆB��{��k|�ň��W��ƪzk�:��f����iY1B�L��rǻo��s��"��^���B��%�b����r�@ђ��Mz:U1~)��٦��X�wP�����P1��\��|U�ø�[隭�λ�;��Q��J���a���F��K� ��R齛�WH�fN����fp��V�ov�j�6��#±n��A�FIpIy:�za�n{��|�]��#�E,�n{;G�R
��|�x
oN�G/�i�=(""�fh4��Y�� u��E]j����Q"�4Z9�;�n$}�>LW����k�}�R�eb�r��w��w��V&f�R����2v|{��G�k$]�j�xT��BC��>������]1?&�u��`u��x���Ԑo�g�z��a{ς�
��>��w3u���Lw>Up!e�үGwA����TK��%��U��.����&3#�9%��J@>���aɨ����e&ѽ*��:���n,b�PQ�ޭ����A�������rڲ�(��۾[��2�Mb��	��=�R?^#���ܚ�e�;��ͭ��R��<���ry�l
�Rd��Ñ̫w��b$5J�=�:A�I��3v�˕�z�t��S�B�ī��A[��՛'^�l�I^s
���u��+-�����F �7}X���Ld��P�ot&20����*�	ࣴ?���O�Y��n\�P�����E$�w���c�Av�7J[ef���P��1�H*�������@���J��NV��=)Y��3���N�Q�[э��^Y�p�|0鈞V�eOu���F�B�U{r���ItMԐ��f�����Ge�9)��܊jU^���2�kc=u��4�s)Y��-	)-�e_�I��".&�Z+�|˵q�vr��}�#��yw@�x���Q�w&c{��D%������a���]�U��IS��֜8N��/(�Ul��~t�-��cgޥ�.3�����`U��c��+gn+!hK;<#�Ve��;�n�^h�Fc��)��v�bxS��dly}�lyA#NT$H��n"�Ac�o���,�ɯR���j9cy�vL cX��Q[8�QlW�mKdÂ��]�kӊtP�`z���.4�ʯ��=A�w]+J�����+���z��x��s�"���s�y,�^�/�jO4����~j����<*gA�@�"Խ�pr��|�F�����������T=��.���_�1�o���V6���j���Ꙑ�ⷋ�W������gK�:���sG,OE`��9��.�x��M�j�u��;�[6-�q��^�
��;j1B��I��^o �s���v;�a��WMA,�.`u./N��4�!�u��c�˩�+�L���s=s`��:W[��N���^q���8�����S�ў�^�26�P��w>��=���s64p)xw���L��@q�te>�v��*{n&�\��i��q;p���x��z�ɯd�>����9�V���S��]0F�r��>
���;��PS�{fs�ݟq97>!��P4�u(v�e�w%�s�7}��n.Bs1��&PWQ��Oo&dn�9�a,�|sZa�e=,̈ ��XiT6�Kr��7����(���W@[��jH�i����d��h��������s��x�'�MA���^�I�[Q|"���]1�ri���S��	�s(f�i���8����}�Vcp���"z�#R���U:�Zk=C�>y�l�\�m���j���x��Qך�h�e�}M��P�{��\�q���9��[~>�;�ҍ���Y��BN�`6�����՟?wu�̉����k��vb�v<�-M��Zc�;'���>���T�(-�`�=�8�vF\�K�n�H�ʭ�Ȋ;�D�"��H���jw�WC8�:���L��*�q��l!�J&���"o �X�R['s��:�7����Xm�d�o��3nM;�ϗA���'.n���Bk�ޅ����|і��`��Xb�Zgf
r�0�b_4�`&�����*���"z�w�5)�� ����U��r1AT�f�u���/�To���Ơ���y3���|L͗=�����ເ�,y8�1A���&�=)®+f;C�}*cR�J�9Z~�<�M�WWy˽��.Px��}mҕ�>��3K�0=�MȌ$��f;�2{�$�cO�6)� 1�.�p�'���f(w�33	�=�	̜�Yq�]�����T ��{�<�þ��Pur��Ҵ��'o��5�B�L�����f74��ġz'�&Ş�^��J�(yn���b�T�ǃ��Ư�)u�72H	i\�E���1��ݓ	�t�Y�q���c�8�TP�w��̎�E�r{�d�o����r��v,]����~��P�_/�\t�5s��|=|
2Nz� ^U�i��嫙CLʟYAi��Z5��R+O��V���ݵ�;f��WC͞�7����vT�!;�r�s�d�f���zcnp.�$ϝ�[A���`��K0�Q��	�
O��&7f�xO��]އ�4�n�����7,X�S�K�Z=�s���Y��@\��i͠��c;��>F��8ڎj3<3\w�_��};���	��[�z@Q�Y����S-�'[ٖ��,tt^U�p[��e���v���3-N!tv�Q:�($Y��q�WQ�c���w~ژ���H[:�v�n�74�i���;w�B8pK����Xq�s��\����'LD�7[q�{�p������&�j�՛���F,�8�	v+%����2�����i�/2� �{�Y.����t�w�:.���h�Lp~���%�����go�R[�=F��s���[�T9��~m]������Պ�hB&��J���P��Oh}�>�fF�3�x�`�؁T�:��x���g�:<�=���Z��}:���D,��+`���3:�B���٬r]S��U.ɾ&��΍�c���_{�����7���H��i����8P~�}�W�z�X��5J�zy;�cف���Py78�jf9�]_h���~a�I�������q�C��먨���]ʠ^�J՗��v�7�WEoF����v���cY5Z$Âb�\gJ\�ƥe�L�a	Sq�.5�m��u����rb�4��4,ddd�[ss�4Y{JW�7�Z�����N��[w.<�b9�v  ��[.?U��g�zjF��8
�^�\��]�uz�Y�N�p��n�>��G�ߜ���wk�g>���= ��O=	n"S���]f��X��|)�`���� ��ɰ�}��wO&Ub����d�����K��Ϋԗ)�W��՝����gYR��Y��)I2W*���~��{h�k�Zے���p�^��*v�-�i�^����}��	�U��Tz�.��쾊Q�N+�u��Ε�p�P�ʧI��M��Ġ��YyoŹ7���LÃ�i�� �W��uL7Ȅ�y�
h�R�q���]�{B%B��oU��ufz�{�C{:as,i��N����_]���(ܭ�]C�^m�,���c�HkW�|�_Tw���*�G �d�HZ���B'
��^� D���Μ.��q�x_]a>��G��=�����}J���]�1/gf��3ݓ�=�P��u��o)Ln��{\R����!�#K7�6��� ��0o��|���)X��[r�u窺4D�z�,z�I�����L{��f�x�Go��beC�ȕq)&)����Ϯ��L�)V�{.%/B�<�såjމ}>b�-�=�l%I-�B�����Ԏ��cV��MH��Ys��"�����ڒ�Y�C�o!@������[�}}�Y���E��yX]=���R����(_y��m:������=���x�s" ��*�&zG	�Ψ\�Jf/���"gʦ�{��)U����\�s�2�g���ܓc�f�.���Q�_ni����\Q��}|������v�]��i��}s9�v18�1���LR�	WWe��5v�9eixi3\N�r �i-����e��)i�E�=*L@�Kw�۬�X�d�1���W(�0�����SZtK��u��wR+�j������=͌]��s����gt�;��+��O��.m]����� L�v��@ŬG���6���f��eF�Po9�&=X��DT�g-Exam��>p�V_R��9<��1�h$�s��F�WLg�b܊J�y��k|␳����0�b<|Bz�nB�ҍ�12��rĢgޡ�nET.��ͨ���ـ�=N���ZY�=�]<�r4j�atA��"�2]�{#�i�<6�י�SJ�P���@�Z�p�eF�A����M�6Gx�u�͜vf��+M�sިJ��O�f>SX��t�f�P��{��{���,���q���R�������= � �z�n}�R�v�ŉQ^��Rἃb��7�"��q�jӝq\���6�$��-ߍ���I/Rq%F�p>�T����E�&�u�?(qK܋�HP�Y�o3!�3��6��o�[8����lM����� L���Ӟ�,��%�>aP�*;�q/�/�7�(�o}����U3��4E|ԣ1m���Ω���*4��5^P]�i��ʙ�/� �E7ݹ�,�۲���xV��i�Jٌ�4��s�(j*�!Hs.1��q����a᫶ٕ���}W4��	̬Ŕ���6��m�W�gn�3˦�����k���lM9��f�c��E�����q}���賴�B�;�H��|���][`�\]M�KQ�^"\&�6�{��<6��O�xM����-]�_�����uFWvS�C�8�oT�1��(��o7�F��9�J{`�����_x}+nJ�h0�mG��P����ڵo���9��U�Р�bZ?c>�&���\�odD�����whǎ� q ���id�\��UܣM��T���H��= ��*M�h�=0��t	�\\t5�l]E�'t^�8~�>���	�SFš㪅�g@'0B�D��f�lO�8�)A�l�](�jI�;���e��γ4�#�G�e�k��v\ږ��;�U�GwA���j��=XX����}<c#fT��z���:���ת�$M��ۗ�l�jVT\z-��w��\i��qS��3�����p"�Ξ�H�Z^y=�&�B��U��e��|}i�h<�_w ��YΥ���t�P���+�t��}	ג6r/�渜�.ܿb t�E�b2@�ea�~;�۶-�*}�}�\���/u�\yМ��K��������&�x��:�T�ф�T���
��K��G�P���{��zj�W㴵��cEM;B��D�ﶼ����i�r(�X��G����	n��� ��h�0�eQ׋x7ݙ�T�y�)��w$c�4_�bd`�+�̴��X���Z;�ܾ�1)��ɢ�k����C4m�ZZ�����`:̘��(���Db� S��/f���{m��&���V����֒�� D;����͙ɥf>���_���/�!eqU��lY��gO>�O>ޠj��K�i9��)��iN�����;��{9Q8�g ����ucF0�2rH/a�v���aN����uf�b ��RD*0�8 �Y��P���h�/5Ⱥ�l>O.��Mɂ��25ŬL�WVJTK�=O�d�3��AY�H�uqG\� z�P����ek������9u-���l��I�8�mv���k����.�
�������.#(�e^ �]��Wm��+�i�΁'K�����v���i��+*���Zq����dR�ݬ��u&���K>$��Sbb���x���Ueѽa�x��¬�;�+iV(�J�r:���^q�v�nC\���[G9w4���ǵe^��X�9�H�;;h���`0�Zf]���/�ܽ=C���xv���r���ۊ�mMÕf!Y']�<�e�([N�'��W�u.V�N(��,zE�5�*P�׹�z�"Ƚt�,�:�j��t�J���6AU�f�A��g��rNO{���0]�\��f�67pC��7���F3�mK���S���י���F3NСswp��yH޸��0��� �i�q�����z9G��G��KE�|�\��`O����ɔʺ��$�5@�h:���V��}7��m�q�e��CV�����\�R��{�V����15L��B��|��&��q�X�S����
�Ѩ��W��[3��R�Vʺ�w'-�K�ƛۗR�ͫv�p���[�H�S�8
צ�Ohv�o1���V7�/�4AE3��R���tYӨ���(չ�����m
�U���4Wl��zW�!�:cF��fb�trVsHs�ܴ�s1~����)z�@s�#L��M�[B
��7��o\DO�+�����>�vY��,�:.o��y�ۘ�m���n������X�C���z��pf�&Z4^"�����7��8[eOm�1���\
�;a���M��Y� *I=J��Ϋ��W���Y�:Ⱦ+6\����gm!1u�4��|?,E�y�n�̭�Ԏ��{��G��� ��U�G���dB��.���y�^�Vz�]_	#�6N�9����n�I�;v:��w�O���`{�8�q;u>�"��Y>�>�#�C䇇�����eϓ�S.�`#�:;���3f����k����kk�&(pP�B�3Ew�*��7���Bj;w�R�[nw;������Ir]����1 WA��������3�>�J��Ęx)e�0�H��+5dP��<ɦ%4˪�N�UI�����u�]��1�ݠ'F����.%��y��$�f��v��b�c$B�qURE�WJ���Mc\�.�	WvXܭ�S4Q6���N,9N����/5��,b��{D�5
�+d�O�P��ߎ9�����q��:`c�����!d������yg'KG��)�km�����N��z;2lc.�T_��p��ܦY�WB�ɼ��:I8ԗI(�sN\]`*s���x�i,��^1�'��܄h̞�C6=��~����W��	C��(�O|�}��+�݊L�]��G���;y�7w�&���[g/�jZ���|�%���)�u3���*�Ɋq�^�撑o|9yWb�jd �y�ag;z.�+mc����~P0�f���|&������[�/. X�醢�ﴤ�Y�c�/v۫m^v�ڿ��c�R�u-�������1S�'�EN�����6�;,p[�vAx��Ţ���\[:w,U�uM�����ޣ��T�C�2�����w�<�}U��`�S��>9�lÅ�!b��߲�,�J�7�:=M8v���7P�%T+����z"����+5����AQgyl�Ň�5�4;��\ikux=wO3��a�^��H�<+)gBx.��J��q8��b��J��VZB�Tj� Nv�W���S�c5Kf�5��;�������q�j� S���ط@�*���yX�r ʿ\�&L�f����#�a�cƄ��ōW�N~�8�PwJ�2�vj��j��	&-�4��C�8��U3h�Cb�o���#Ԭx����8�~έ�b�pV#�߸���';��D4��a���*�A�:'xjyA*���Ŧ�~*(,���4���y�äɘ�e�]��*�,��軨�6;��>� R�����ˇ."A7��sr�w��G���s�*U)��<�ľ�q0��FպΗ�pdH���v�#�0ؘٮ��:�ˡ26`P~ccj.��JX�����j����Ƙ���Ղl�ЯA��j%`�N ��~�'��y��V�tၙ'o��+�NÍ�1�h�/=���s �2 ��6�'�B�x��m�OmS�L�nԪŜ��>(����y��{Ʒ��$X,���=}>�Jl��"�[~7��O�}y���{<���N�a�3��Mp�l��l_�<$ .�����0��^!�Wq�j;dV5���G+��ٛ��ְ@��0�'��w�Zp�f�Uʴ�-nw��>w��{О(���w]���¶�b4炻�9G 2�6V0�&lt����5Om��b�jd�uFٺp���Md8��Fm��b��k�/����PY�[$��T�f�Kڑ0(>��w�{ta�| uU�*�9M���4��
����CEZbw��%�S*�=}MÛ����VC{=#�ΡE�2����󯾊��"~+�Wv�%g�T�[YtA�G���CWy��غ�
�����nX��S��dyT�?mq��8���tX��>6/�sHv	13�U�k	��"��ۃWi_Dه�3���n�{\���$�W�籂%�N��t��碄1ލW������xv���?�f~G0��|�]6��q�V�$٘�W��z;MK+"Ю�f��3<Fp�Q{��k�G�Z�8xe%U���C(oq�&�NƏ$����p�[�5D-���9Wb+ܾw�YR����pI��s�\�yb��~���]9��Vz������6a�SK;�o�ű�Za�i�j[����P� �ޡw�o���I[��Do�|�2�~��/EQ�ښ�-����q��'#��3؈�鍋�͑��˵K=�[����դ�:~-�o@�GC���G���q�~�k��+>�y��.�_͛���ч�)]�%��������Գe���]K�i�����i�6���c���i�X�q�tdL�P��<���X7~uC��hPoO	u�u�@B����a��OtȪ�
���F�K*�]��]9o���%vX�)��-�t�%L�#��r�I3�M�8Tᔚɵ���5���U��}�}*��]�(��C��wæ�3Gi�b���B�:��W�Au��)g'����
.Ri��v�>̿Tߒ8��;�0
�C���K.�X�+?b�sV�����~��޼������q�S���.{4iD�$��˵�������>NH�߰�g�=.�\�|2^�iY�Ļ��S�Av�����t:�r�Ҽ���z��x��c����{�l��x�B�ޞ5�3��ެ��?Z@�5��;�̢.;���@��zW��P�&�o]Z8�"�wJF_�_�t$U�����dI鮌�1��S��S�ط��h��Y��]Nl��OWG��x�����g<�}�ѻ�1�c��U@����3�I�?�[�47�$u
E>�~q�M��@���^�y��]����u��d�r� s�%_LL�@�ݸnԟ�}P����gCƵ�� -���u���*Q�@���p1:�Y/ ��ƛ�[&� nq��Ǚk�M7�gYW� Z᝵�B����e��Lb��-��ݒ��7s)�퇵H]ؗ�k�[�6�wm1��MN�zͮk��yZ�Y�U\�f���S��5�vٛIu���w�n}���͞����ʮ��G>)�7<bٞd����]�f3aS�	y��<��U��w��%a��K��u�f�F�����lR0b�f&�E�*�K�R[� �*�5��1��5�����%�u�ůG���"L��b�$xX�o�vߩ|�ea��p識�3!�!�u���m4R�fBб�J�l�&�e)%s����7��;=��s����Y�}%�d�~o�%�.����A�� �r6�{L	�m"�a�1��] �휤Ur�}�>'����>��S�B�����r��R|�so�1�1e��7z��9��[ڎE�WO� ���Y88s;M:���vY�=5w���d	V�e@�[X�|(m��O"��ؠ�������J�Hp'�x�4����s��vfy��d�z=�4�z�_��r��T���:;	������Q�=�h�o��C��-|6+HN�zM娬�m@=��vs�l�l\<,\#b��.��,qrV�.�a[Ϸ��l�"�s�o�/W�iKc�*�r�U�UϽ�}�)���;u7���)[oxbvf����t�1�z� ���0��܅�rD��e��g��C9֡�˨A��Br��g�/��9��FgX����Lʝ����,�fu	ɻ����۝[B&^�n�$�K��~��={^���<3��<}�%�g�z��Z�T�Rڞ�&�G��3�m�WCxQ4n�Jz\���!/|B���	C
*��`�85 B��*d���y�Y���:�1��mxwk�����Mpb^��Y�TR��_X��2���5�7a{GY��Ӽ���g%�ȳy7&&P�n�B�|���]iK+9}�q�t;X�?Z��F,�Ne`~��m�J�����n�%b0������.+;��j�z���N� �"�:[fͫ3��N;Y z�'g[�,ƍ�zxx{�9������u���]����0�wn�R�q/�|{�S$�GЕf�e� 	��/F��˅^�1;�:�%X}��oo���c�
��*�x�u�y��3:ٻ���E,=MZ&n�C.��:޷�|�Nlsj�9�f����h	L�oDp�м�L�����Y����V�3QK�(��CV�̑e�1���W��)'���mv�8�Ս���S�\�⯶��ZWz#K/�"� c3ΞA�3���0r��>���W��f�Ev�k ���&�$�y(�z�*��*���X�������߽���f�'fO�d��:x���鹨+2�g_��Kb��j�x��1P��M���8��������>�囫�̧����X�͂C�={��v����u��[��{�S���='%e�WU��rP���')7�D��560Q�v*��B-ҨCLG�n|jI����y] �%��$�x�i=g�n��G�j¾��}���nA�}�������1"�`w,��-c�NNN�w�=0vu�z֢�Y���E~����7�j��b�%j�X��f�f2�$d�.^j-u�����������҆>�<�6R�E�2:��3�Y</����"�?7}
2C��nj�l�6��ƉnJ'���n��f���c��;v'gZ��ڻ%����|�5�W)��6#9u1&��Sɬ������+B�5}P%gxs��J7C@���.��S:�o埅�/�$�;���4;�VY\Yb(�>��wv�6$Xy�[ӵ̬֓�&�\y*�ͻ���3�z��x���L[8�9��Z��\�'r7U^SuR3�u['�]�����8�g���C|F��t��dx��B��"ہ9����<�;n�?r�>�vK�O�����(����_��"�NǷl�\��r�{��w���*�ђ��J�� Q�xWhܨ8(9�U�/�8̘�<�3�����ɀU�&{۴�#t.��O�x+�W�T�nsw�W���K�mt��j���׭�������R�/�~��C�ބ�׬s�K�s�Vzb��m�3�H~��G�b�Ϯ9Ϻ0�첐`*�/ۖi��$��Zzg¶�z@w%��k�:<�����3Uq�.<@頯n4��
�(����/��k��b��źˉ�cg��¯�wJ-��u�p��Z�cg~J_�`��̌xhY�Ng�q���PՄI"3w�'�]=�۷�U�S#�n����?����K�SP�~p��
�_���X�W�S�ϲ���}�b���S�{{kV޷}ě�n_7��uK��Ǵ�N�� �
lE��<ū�pc{��Cuil���jI��|�>`hDTYΆ�����3�.�۲��a)�ٙN�#�YX��7��n���_f�I�:�؉Rȼ�6���b��JV�|����u�-�ض�`��O���D�q��D��z���Ƌ9"Ll��*�>�~���0��}u�������1��.�����'1ؿ]Z=���������(s�>��mwV���d�]��0c�$uu����wd�x�A��3�]-����i�+��PzmL,�22^6E��x<���C�\E:̟O7/���q����=�!�'Tl6S�ތ��ά�g��Y|�ٱ*�2�=��<c]Q�fRڤ��q��'���?y+π�x���>���9q���8�.;3��@�x��b�Σ���3~�@�{�]�Go���˷�ʻu�ډ��j^����J���ձP~'��׫��@��")�<�GB������M#
k#/	.��(7,����텢>�����Ʀ��a����2���MR��<T7ި��]x,��Jy�1��_���=����s�C�y5�$�{�W˷-T�:�sBKYy��G�w�ɂ=��y�t鏯4;M���r�b�k�4.�h��P��F,���Sd'3�؜��p�~�7h��R���9��i;�eeEw�xFk�;edWCv)f����sU�@�%
��ʔ-������J/0b������娻V^�`��k��t��&ۙ�U��;?�\T��"�D�%%§�<7������<w��X���5�G��X�R�9ރ�a��,�C���:Yec�)��z�����M��^|�����&�
�l٧����{OI�靥��|/��%VL��j��٪G�oهceB���fy�j��S������C�G�]�{6�[�^�&��~~��C�Wobs�s��)}�����S�6^��s���ڏ�!���� ��p�5v��%��hY��J7�]n�ؚ���P/����Y�'4���y���d�3�M��l'7dQ	����=+�qm������sY��Ur�!`�E�h�!
���!/gt��{i��U֣��ӳ�eS1���n�(�d^�{z��b�G��
������˥�]��hz��#5סU�D���M\t�B�Շ�J�NѴo7I�hԠ��� �DX�;	�I����m,���vrճi�`�u d��n�[��ܮ'���%ź��cd�J���-�ƴ�[��qZT�ي�cx��d{�8Y&� F6�T�����-n��:~���mM�"���c�%{�ך�k��7�=Y��w�V26l�/������9c�Ė�NB^�����!���@v;�hs@��h������q���g`В��FCwYK������PU�;�	�Wa>�ibsРN:}�m�r�ܽ��h����Wuf���ؼ<Mez���'�K�r��Z/�W7��劒d{!*� �<N�,^��u���(С�X7�7bm��(2��(U�5׋��c*앣���y��Q��Sr-Wґ�J��r�x*�XKᡐ�cC͕�W]��i�[��e�f�%��x,���>2:�<�WJ0{�l��pƳ��.�V���� �	yȘk�E;B� 3�e�AZ�1�hM� l��En̝��p�q�j��O
�u��5w±T�}�Vn��:)ջ�B�I
�6{�wȐ;'�k����N����| ��YK����3�6���|8���Ż�aV�͇�Kqf��<�{�0R{)����	��q�����ĎݴT��wj��܁̘>齃�%+-h�����s$�xG<��}�Z,- i ��W�2�d��*f��	����Y*�Q���"nq��ssS*�6��ȥkqk+V+�5pK���K
N�ɪ�q(�S8�j�_=������q'愠�K��d���o�{7���n��
G���ͳD#W��Vi̽�R�QYo�]�8IF���՗o2��U⩴Σ�g(֝�3-�j��!'S�kj��=o;;.A�ҹ�W��\���e�D$�x5�AZ�x̦9�]��oT�ъ�_WY��Y�!�-���e�ܬas2��\��au�Rs�92�&��&�8å6��+.hD���)}�)��������6pX��̇*��]m�ːp͇���0�W{�R�e��u�����w����g/𵙆ʱ��.�"�1�J����C���WJ��&TԖb�N�́�p��ޮ��t��"s�K����_k�·_r���{V-G�k;!��y�!���nE@K���X+	�2qH�8��<�ۢ3s]�:׳��e{G*�������(kK�|.�'��s��*�2[�&�����wFEc+���n�y��mӜo{1<�S��e���g&YB#)�{ʆ�:���IN1�1����u�=������0���R�79�V7��m�7���Zj,'a���픯^��v�v{�R}8��aŉ��G�o��v���QЂM]�sí��}Y�+O�t�[W���v�;z�n��"U�]�3�pLի�Ώ���73�"�������l��\u�z���ߋ�ӗ5�1m��L�4����3�p����,�l�k;��[��u3��̓Y 8bh�4ǻjd�4�������3;�*Lm���4_i�X�kr�᫹d�� �V�n�n뼫��f�e���!O]{ٹ�v�Eֳ[#�]��0γ�nEJJ�+��+ֺ(CP�U��o~;O�}C�0�A�����M�-�L�}_Pg�۳Ŏ���Z�Pa�#��%.��=���x߈7AG`�{��0b�<ҸΩ��o���d�[�#/=;O�Yן>������`O��ao��1efE�G|aW�P.���Eǰ(A�^�x�	ٽ�S]�r/�
٤�g-<�p���YX�N�v��ڦ Q�������=�_�� 6�j���/�z��Wㆨ��y֡x�7�g�Oz�L����\�=��?�I�p�[{��kk�_�˥GqV��Z�w��gϼ_�����GӺ��>+�R���s�Y1V�)����>��#��$uth).`5��<�$[v�c��Ac=�wf�U!%l�w��W��/�#9����u6;zf���9B~�F�<*�0����gT暍�};11O{��T�-r���I�3(��1]��h^f�d�rL7����2�4�ͭ��{�\/f�FH~�wsf%�dU-��-Ֆ����������:sJ�]ήoM��}�t��cw�V�D���F ��ORNl���Ȯ{�\yVPf˝]�+V�=����UӺ�N�l�Y���Z[�Ϯ�4�q^�κY���,�%?<�]���ܡ����}q�����=Ȫ*�0zv�v{��&%�t��Ex�+=�B>��N����u��9o�~����\����潔��~����W���q�d����~7��)�9�f5eF?���۽�0�N���g����72Ԍg�~Ӻ)ܞ{t30�z|�5��(w��sؼq�L��v>v��ƚ�|�\�p�׵�׽�>�Jȗ�y���d�0ng�G9E�(�PG-J
e��st�������ފ�B���+���'�_q3%-�sJ���Z���(cMY���*�Gp����*�3ձ�*�.CвMY�1��+�@|�x�v(8���5�n��z��o��}�,#2�X[���RS]�Y�{���W�u#Gȥ*kǪ2s��5�����j��1�[M�CM�V�'���p5{B�{��F��Sg)p����L�K-�;�2�v���v�8��un�������҄`�3J.�O��Q�X9d��ֲ]�f�=�i!y�;�*nㄻ��nS{�A����Q�ʹ��2�^�]���K�q[��L޻���Oh3c�lx�<�3�w�WeH.�l�o��lI�N�;���=^xegL7����`��}u��<�>�zD;x��\�qĐ����u��u.y��c��0�X�/'�,E��{���ܼ��e��ʴ�.��U�S���
��ً}ޭ5�3�U�
�U���%9�L5��E)��.,se�n�dǥ�T��;]];5�l��(K��K�м�tա�;�L,(w>����$��a�6~Z�}mC��7��U�1�;�\����k��ڶҎ�I��}��f��	�K�L�FUV��=]�����]F�Ln��3V�= �~
�c���o�>��۾�,�U���]ׄT���}(}N��_`;�xЕ&�S~�c���{"�z$��5���Y�p�s�<��/_c��0�ў�_�{pSb5�]c�G��#��33�[<�,��@�;`��^�������'�'^!�Uz���]v��U�8��8��]�Z��y#�ۻ��+<���Ƅ�l���i*Ĕ�s����e��\_35��( q�I`����`�*���@�'�kN�3�]�Uu�q ^�]��Tܩ��-m���N��r.��mC|�w�]A+r�����Wp𪉍�8��/�=7�Ʃ��ߟ����?\d�)0�FjF9<|�����F��lb�!���$-Cc�;���.Q�':��U�yi��+L�}X����ݫ��::�&X����7�ʷ;���n�����%S�'�53G��GE���y��Q�����W�6���o�~���}f���1�O��9�L.WWP`Ά+�ڼ����2�
)`����"Ж�o��g;3"�|a��{�O�����]�M��-?SAՖ����{҈�:S���{���^&�HB��^�c�O�����ԥ%�#������z�P�9���Ϸ�Q}��Hx�M��k-����BQ)��ǖVe��f�&F��9��OLfMAO�Z](]��/� h霣�8�T%�0޸�o���1�O��j��aFjl�:�I�y�W+��HZhvr�J��s���f%���_ 6����x�f�9����2�M�4UXWS2Buz%ӻ��-��)?:��=`�Ħ�R����{��n��2-��*�+w:�.��z�=��jz��3)rZ�}Kz;��ӻai�g�?��=�X��7�F�v7���]3��FF�2�ۨzi� �6ɏW�/�����0Wf�k&zm��}�=j�tTy^�1�|_��4�Q[�\�0}i�k�W�9�&��O����Z�F,!�^��:p���T;ܟB��!³\j���ԝb右ܼ#@F��Jr��6�z2'
��н�Ǻ(O���'=�A���y���j
w&������nt��!'�����tQ���S�u�©'\�0g`�Wt���Cyj=��p�˧��口�f�3�'�Z^��$V��\vz�S�a�BT6�IÏV&:\O)���:�`����z���/���M����z��Pn٣���{b��������k��-��b��������"	=���VB�q�o�ۘ����>��P7oϞ����?���4D����_\λ��gYswq���uK��{
�9�����uc����1�؆�S6.}2��eU�9ڗ�}�L:�]�S�`ŋ��^���k�
�ci�#������9k��3��ƃa z�y�v�=ol�t��,y���x�	3��6�F�U,���o��q�F��Y�Pg�Ny��bne�������3�s�^�(��xT�tn^}y�|����P5M�%n��l���QP�S���� 5��Y�*3���rdi��5�y1���;�ӝU���b��QW�[�%-r�7y�~�u�2ԓ-ؾTs��2z��G�^�޸��eЬy� Q4a]Z-���{c����#���D,��ۭEm�ԩ�Au=�n�6���$�O�����U��Q3Ӥ���'�F�[9=[8.яJ�w���/�Ʊ;uG%�:0ښ�P���Ix(;�)�C�}��n�I�-��?	��+��!�H�vC̘�9�^tE���63�v�ӿ�����`��}Q?�K�A�b����,�G7q�*_i�|Y믶^g���}�R����^'�v�Ȝ�-�o�É?M����L���Ȯ�5�W1����C'[K�$�Z�Ic.җ>�y(��[6��{V���ef�y�R��"�+�R/�(J\8s��,�����^���h�p�Ұu��{v���uԽ���j�Ko��Ω��[g] ���.u����f�u��S�u� �2�:�g�����ޡ��r��s8���y����~����g@��XJL�o�c��w�
�/5���ӾV���0w-F=Qo�*��ٌ�Q8�J��E.�9=���άA�2� �=�}P���T'
b}���*#N�*�[^�u��KZLz��t6kV��#�kDyW���[��Ŝ+w(�6����(v��	�3�bW�h��'��8=Y�]!�f����;1��,~%Y���i�������7A��Á��o�.`�k��굾��ۛ|Wa�p)1Hl;��E�a�I	��>�{k+�0��R���1E�#7���@�6���^�2���Pī�u\@W>�>fyg�_��XXL�_d�2GD�׳�u�.+�g�T0L���>�T���B<ߚ�{�~^n�,Z=.*�I�����~���vIi}�ֺ�;��=�/Lc`��u�B���l�G��{��߉���͚ù�6g��,����`��u��M3wo��=� _w]=�b�{q�.���Ӳ�OD�P���W�8�-*�VL�&�_Zp���(�g[�w^���S��jdN�o��L�S�꾛��.�Y4�Ps��Euf�9A�J�ng"�5d�$�[�S�'.9����>��:P��ָbn�p�40U���1�zzB��ײ�ɳ���"��bG{�f,�S���^���~+lo�g������u%�F�'7ݣ�'��,Mz�n��^�6�t�Ƌ��U�N�N�)�/gg��x6ZƷ����c�wen#�����rz�%�^��Y�;[&�j��6��V�N
B�y<79��yy�'a!�:���ǝ\+Ԯ�/�ϡW�ִG�G'��)m��oq����}ϕѠ���{�syhd	�[����W\�ks��t�g�� f�~���6�d�|*�bNfϣæv�=�x��٥���E�A���k�����F8������G��UY�����%�ۥ�Q�K'�I�K�����o���C�H��#&�vV�n�ꁠx-u.恘�ɕ�o�6�+�s{�o~`@2�v)�и���鉱�����5�k�/b��F�T+z��1؅I��ͶUup��uiu�#P�v�$~�%9���z�����:��_N,b��}[������7ôqhWtyu.�]3K�V{7r�v��9��6�m�wS0������nu����r���W.��,��=���~��ּ���%��\ym�3����ZB����߇�^RPN�b�,�W�b�LL�e��õ�d��̖,y���	5r-��w�p���X:�V,�h���E��|"4:x����It�ٕeþ���79oِ�����Z5g�0GՕ�Sr�V}]Y=�q{���ޟ\��_j踨�>���}F�0�4π�I���x��xy#d��?s��{\֛wS�����>^��咣+r��Li�1n���� `]�Fd�ڄ��볋�`,X��qj�	��oh/�4���m���L-b�t�¼�� G���P�ɚ0�K��VIQe�/R8���.�W�E��뢳pwy�Eu�B%����;5ɠO��#$�[��킏b��1xz��¼����F-�v�r[�:�^u��\�X4��g%�mU_�۹��r�ORޱ�_d�\��>��w��(=���kxta]7p�I`�-j�=2�d�[�B<�v����+R��]#��u�J&����w�T#�;SW��\0
��n�̘s�J��ڗ˜8��N�vu#�~xR�8���yX�C?m�m%=���R�Wu;��O��x��Ľ9��%�FV�㛰�I�kG���F_?B�q)V�����vh��ȵ�r���C�ګ
w��fֿ>�3k���:�Q8&�X�b��7i��j�y?z���q9yџI��b�	=�	yҞ��ѷBڮ4�n�L��`WC���t=0DG������u�nz��ˡ��c|�N�}��o����[u��g�@��#-J�:�?G]@|s��un/��ԏ�`YFr�[-/�%
���~��^��{u���6�)\���.V��M��7ϒ7o�b�z�w:Er)GM�Yy��g���{�8���|b�AafE�-��z��� �Ϗ^�w^o) }���4]o�[��{�0@5�/v��;����'�uc�Δ�ª��ӝ�n�lgT[���~v����|'�i��(�����L��+ܼ�Z�#ƺ�^ՃTʷۻ|U���9H�5�.K�d��+�YuQc(f�I~�Mfb<о��ad/��t��k=Ϡ4�K7Q�(Gֹ}B� [Pp�R�ƸQ��Oe�Kڗ����KLNf�w��e�/һh�2kw���<�E�΀��͇��so���1}[2;���nL�.����A��.�O��>�> ���~
������f��
(�<h�9��
 �ɠ2EDԪ�������?L"(#�G����������/~~���|��>���?���R""+������`""+������}����q���?�����_����ւ%�<�@�������I�g�J�j�^��(�%or�ۖ��:證��|�p�¹��V7a�f�Pm��ґ����SP`,ʔ-f-�BJ�f���2��a�h��R�S�-�EÅ3-���|jb�����0$�8�9|DP��N�-��CE�eͫڱ�/If��;,fЪ��0k���[ �5�j��ݦ�����ֆ7rk�P�p���Y���k9�YթXۢ��D��*V0+%-Q���U`�AQ����Ҍ[�.g7ϧy��b�'����G
C#���t�ǲ�U=F���� I�R������;�ZuY��^"ibW�bΜ�Bg,����n��/:Lu}u��*N8�LȲ�SL��7�6�0کL#SY�3`�ә��2�m(T7w{���7fl���|�ݚ��[	����3(����2�²̅���;�&��p
84�4�f���֛"��zwX��T�ǘ�#B�r�^Cx*Z-ȶ�il�O\�p-CKb*Ѵ�c�)b�w5XIF�)F	��Ay�h��vǇKN&�v.�s&��*nCg�ƻf�F�f��kP��4)f��d{�Z,��
s�����8���=��Ʊ[Ss���X0��XQ[5f<ǆ%x��Z{OV�{=�ӓ8�O[T�uj�O\J�%9/�P���e�"�˫�W �ԓ���,H6V���U�^-J�`t/#�kf�:^���Mb0�(x�T��Li�6�6���) P����(��jӘ̫r��9��mX�țgT[�n�I�jV٤ڎ��"j�ZI��f��#MfCn��^�"*����Ϊ�6�I4�;�aM[MɚM�%Z�d#I�����)�[���s���W���76̻ݏ���Ef���5wI�gE��*���V���*ʹY9qMv��XM?�J�rԤM�Մ��7!�YD[�2�9�y�@Y�P��2S?e��Z�v���t�י���$9�]��)MX�7;7�S3�_Sʰ״��X��+J���2�˺:mô1������Bc;�����T��e����l
3X�L�rm3!����K�i��8�@/V���c�RCL^ ��Ya�]�LK���$��M��Y��-Q.]�{��aC�0^�u���W|r��wK-�@��P�:���̔O*�����M�UT�8��U�A�B\�P&V�Z!��r��L�MN(��ȹ1P��#1��gr�Y�j�֪x�M�2�tbr�uN��\���ޚ�e��+��Qz�ˠ]XbH�M��	YIm�U����˗�j�;C8h \��l�bk���ô�6�Q���+̄��7�u�{~�j* #�*��*�H 2���$"�������(�
�(�# �H �(��?�~J��}/G�}>]g���q���DDE|����kO�����~~������_>!�����Ϡ�DDEy=������?q
""���rlQ��k����M��í_����a�ٰDDV=������DDW�~�B�����<G˓x����������Q�qY�C�������'g_|g^�""��� ����Z�L�z������|O������|""�|�g���g���
�2��q3���� ���9 ��>�x�{��m�M��u�vj��Zm��@ sJ� �a�D(m��[�W"�ƺE1��[�w4�a����l����P i�R�EZJ%T�
e�"T6�ʹ�����QT�`�T���6���@
PJ	)*%
�R��6¡B��Ap          �붪]��*�;6      (���� �T]bIK�P��� � ��pPHPV��� ��t�� :��vw�AӡFۣ]�8�:�vgA���M e]���wvƍ��R�]��f`^�à� (4 ��x@ ��� ����[K���2�����r�ek��������W`�Yx���n��v���5��;�Ս�������>�o����K�:���W;3;gu���׽ķn��W�F�֙9�¨h�"��ƾQ�x������ˑz�Օ�9���r�+�}ܯ���d�����ʛ[���w�d��{�Z��G�n��뺙S�WVM[��wo<<���]-S�_}�^�:�.��_o�a���k��*PM`U>;��u��]����޻F6���9-ܶ�s�����c�]��{�=��Gn�s���n;=������a������ݽ��u7��:������v^�zy�٫����i��U�����l��w}t���׫��\�i͵��]�w�>��o|��뛹���>��|v����ޤ��ݍ�5s^\�9w�����4�.黜շ�x�Y�)�c�m: �F���3٭�����q�'�Q9�:嶛{�n��O|���5���=��F�n���k�07�����;[��Ϲﵬ���t��=ON�ݲ}�[ܻ��I�������WY#[XiE"�>�N������:�����lݵ��ӝ���Wm���s�Y龾�K�}�ou�}�Er��|�W���Zes�|����s�ӻ�N��y��w��u$����p�*Tv�JUQT�<�|Z�ު�J��]��[ݞ���[ݎ����yc޻V{�׷oa�yj�Z��ɚ����']���v���y�]k6���W��wk������n�[4�hЭel�]���:����w�۹�n{�}}��h�u�׏:�m�s���x��}�����f&�|�y}:��7���Z�â�h�%�h�����-��խ�ﻮ�㪀N�QZ�YO�|�]K]ھ{Nd+^��{�'���wk��7=�ػ���e2��z�W+m�n���vMfv�}���f>�.T�וW��{���mt����eT��ʷ CSh���� )�IIT� h S�M4U!M?TG�� ��RU@ � �@OUU  h &�����i�Mb|�>�?e��g���7k�e���bm�����r��i�]w�[n���N>_� HI;���@��nI$ C���$$��H@��X���O��!BI���!$�@��̿�Ώ��?��s�,�����X]��hO�6���ɍ\y��T�	���RjF�^�<7�R���zC�i+�T�*�	p�h���z7^^�؎�Fj��0-�a�UEYH�m���4���i��r��l�T�P-j������P���d:�/k%m�I,�n�B�a�LG�e�Z��7��#E��
��Zãw9	�G�gwzku2�9�s4
�7C�f�}�CX˴�>�%�SL1"1��A[��p��ر5�W��Tt�k5BHi:_����Q��F%�|ܭ������T�i�!$]Ja��Ma������4[�ݨ�7��G�t�.�F�]��*"��eb$�%%�`xRN�p���
���h�.��h�r�Al[��LrP�tf�V�ֈw���Q���_��PX΋	�VH[Wb���)�nIFe�~h4i<�Ϭ�m^UBOPrR�S�`
��iMc2�m]�6s�A8h��xE���J�-Y	 `pi��wME�1�0�r��Z*Ҕ+�s�y�׹��e���������O>�#��%@�C��{5��/3�̖켺�{r<���6'�)��c	�DZ�Dn��.�0Vn⤂�q$�m��n͙6�I2i-ãE4%l7�A�M�+F0�iL��e�馍9.��)#v'��
ǆ��LˍQ�����ʅ���4�Ѳ�<v�^V]"�8��y;wZױ��ߡ�l���7*���V�ĥy !)x6���U	h�E�
/]8,�`lk��ǥ�E�j�i�)�K:�w�ŋ�r��ʭ���Ï��M�U{��OYU���N�4��bPG7ķ5����c�m]��[�ӗ�.ْ�o�)C���7�c��4���T1�VC̘=�(�@$�|�L�-�Ys/�B���m�T7�V]�eڪ�6��#�"Qp�B�P�x*D�Ecr���?3.t���˘�:�NXγ%e^=�3�GO,���]m�K��*V���s@Jn�h�a�t�Kq�sb������675�;$ũ�2��>��D:�q&��')F,b�PTGOU�i� �`���X��(��A�G����Xd��!�k59���s5�����ُn��z��F1T�� ݃v��,P��^f�n�ř���� b�(���@Q�^�n�9<׸e��n�6�*�Ř�~�#��PiJ���SrVΚ.��Ybn6�5B0 ��\4��ۨ�[����lx��f�ڞTm�R��/]�@��Y7 �8cd��M��aZ;��٬S���2�z�ͥ�D7Mb	.��#�k�yYT���J,����-�Ì��,Ia�'��0����j(��!���.ގ>������{H�w5��c�V
Cl� �no|�>��kWt�e���نJ�{�[&�{��>6HiZlE�eIY+:��@��̍!b~�OA�2jMZ�M9�߷�ߎ3I�wٚ��w!��@ǌ<����4QeDQZ�]RTհ*VN�q��C�1I�E'I$82m�C��P�C�
�R�ިi���ac�AHq�&�0�4��C�06�� ����9����dՔ�i��<��C�!P�-,a��r���
$�`i!Ԃ��C����O Wic
�T�YRc�1�Hi�{M0OAM$6�:�+w��X!}Hu�ąHV��Y!Ԇ}H|��C䇙�1!��Hs�C�
����u=��Y�w��5ϻ����0X(�7oL��gl�v"5:�Oh�j#���v���0ГvYM]���+&S�5��F�P�Q��^eqEr���=ǵr�� �:�L�!ZmԠ�˰ⶢ���8ULS\�ZY��oB/&T*��h,�����,9�!u���H-�f�Xc�ѻ�R3RN�4V��Z.�`�̢)�0ѫ�����nʆef�
ͷ*[��i ��
j���[u�(�T�f�uq���TU�!{�^��b�b�F�`�5MN�2TOC�DQ�#�wh]
��2p�I�k#ʮ��q�7g5����f�Jyc5Ewk���Ы�N���)X�ݼ�r\r�!2���imӃ%����L�1� �bj	t�ӈ⧵�6�I���u��x�6I�7�l���L��ij���ה���d�a#Bv5�h�n�.�e��.��u�%���,҆��	e����bi;En��������;��D��2�7/+Ptoj�&�TB�ʂ��cH-��+v�ghB�9 ����ӊ�Fk+V\2���>�s~��W�M@<�T��������������ʅ�_i��X��,�]���*�JJ�e(�F�T8��"�4p��mȦ$�n�D��Z�؁�ᙆZTi`b0woje`נ8�15�iA��.�TV��x�	�Jيі���.ȳV��7o3D�7X�l�n����ֻp)PVl:E�y���p�Ǐ4�ה&��6�P2R�6��'��9��q����Gw��w�`��4�h��YN���^����I���;Adk�p�����J9�70���V#��På+�1ɮ�&�d�4��1:קs�j� 蒈�l��j��z.��a�����uBwkDc :A���	If��r�b.�%*p��y��QZ�͠[yf�S�`4��a�3H�""h�T 6ΌH]n]�k+T80�6�^�XQ�[�[A�.ѹ3H�k5�T��O��j�ooS�JW������wKY�w�a�/4����˸���q���%�~d�@q!�#zM�Y�QB�K0}�*�M�J�L�utS0[8����l�gC#'��ˏ>�t,�x�:����|�e]�n�t}��ȁ9.�94�����^Cq �ZQT�´��m�	����b7�d����(1��Wy.Z�Pf�;���GV�8�)1�P�̎G�["��û�.�f�D|0��Ŋ�������r]�"
:sj���N攰P�m�p�駡7�!0%sq���+Nf��N��\;m͸̍�XB�����ϖm�8�5����k`+n��ʎ˕�&uޝ�͗R�W�iS.�J�؞leSׁ�����4��B�l�ܚ-XwJl�u���Y[	hXb.5�#��m���
��ES���򎋩��nƼt$߸=�S��J9���؋�\D�aEܲj`�Ι�Gu�43��s}���9���Ω3�H+�6c�Ϛ�)�iK�9r�T���p*�W�iE����C�]��y�������m�iZ��I��Mcr�]7�z��( m$�����-�;K4Ф۽���B���Xr;ͅ�BE[�ح<j�R,Q�Q���yiݚ�4����T.���<il1�J�d�k5����n��>�4��$",8�~35�o��{�&1Ao5�VE�j!�n�H��E���2�ρG+*]��$��֨[ڱ�c
�G�L���C�RUiQ��a���� V�Xe�4)&���z�׵��QԢ,�DQ�۞ �n�uU��j� �O_�0� s41�cT%��� �V�8N%y��y)fcXN:0�e
xdHPy��BT]f��G�-�hEl$j�0�1�	[�"Zgq���F��RFH��?-�:˥GN�f�{0��<A.�d�T�Bd�U6���Uqܧ���]oT�imdQ�5u��̦������nA ԐӰ[B�ݬ?\ի�K,�4�.䪱>cRܼ͹h�BnF(�3j:[`�˕w);"�D@�2�N�a��(c���*�8S.m�A:1a"V���Z	�я`9NŢ�H"�ȺRg���[�"���m�R�K&�Q��c/7H&�����5��ฬY���w���^\��v��I��I�~i�Ùdǖ
L7�}��ե�.ޚ
�c�G�nh��S7^��ڌ��7,#*�VZ�ɫ ��@䱴+fA6��\��P�*���g0�˽%YŚ�����fn�9pIjô�]eĝ�C%FL�ذ��h��<jDhm�H=�f��@zI��iQy�		�b�\uz0L�^Ը�ї�GWL5&,Z�8.e64�7Z$;�6�FS!l��h�o�4�A�% Nё���������9���f��)k,�e��t+Rě�N���o&�wt��2Kf�I"��WB�%bSf���NmUK� !D�~��`�H�e7Z�65e3�o��m��.��kv�u*�SNQ��n�WK�U�R]��J�Q�xɗR,�X���f�Gll*��Z
���:~G±�d�i�
M��/r��-46�h&VǹcYxZF��� a�p�0j����#%�Ce��u�l��]ؖU;�s ��or=�/�Xv����R��C`��Q�j�^Sz��7�*�N6�wP:z��L�u����KtwH+nJ����v��0#kJ�e��-������Gp����Cbjvp����bvVͧ���!�;��[��*�DD�$�&��jPᎯn�5�:�e��x�}���gę��쬋f�4�Yr��F�[�f��/okX �KGlޣ��ʽ��ұl��)]\6�E��f����n=�$�e���F�J{�"T���(Ԧ��&
�b�swNkw6:[��x��� ke1��,`:��t��H��2M���m8���IV�Ҷ�X��V����f�p*�fjR�2k
�{����:�n<fI0�n��!̅A`�bC�<�+x�(!iDY�aąc�_Y��}�Q�s�:[�h�f��)Jrt�s۷�Ă�C�]8�CBő���e C�!�s]i�op�i[2����Bכ(�K"G�mf�l��5���eBݢѦK�F��ɍSB��#��y���m&�@E")u��^wu�
���o+Wz2�dɭ9P^C�T��D����.�t�ZD���K-���&��t� D zD�M��3n���B����Y�v�Z&`����V���[z���J�Bd�+q՝m �mH�P�i�yh� ��q�ö�w�K��*;[�f�I���Ȑ8�i���+�Xt���Œ��g�n��Z/Qj��f����ը�`^��T�F�C#Y��GD���f"��z��=��K�aQ]�t����l�4�<ǲ:j�j[{)ҿ�݌��������2(T���O]4.��m �ݿ��7^�����.�8� �&�	��>w���Ք��GssJ���VR�������A�4�e�/":���fԙe����6�p�.�L=��Je�O����Ѫ?��x���ا U��vJ�Ǩ��mfJtm��G :TSvfKȀ�����E�)�0����Q����V�V4�ڒU�k����*
�1��*HLS�"nR��Ͷr�㬤�Sj<pP��*��h`ƭ[T�Z���P�%�ճKת��+e-g+p\9j�nM�b�{-� 
�V����e�LzVR����ՠ69-&(�{m���X!��טf��K�WCH��V�E���`nV�N��j���1^�Q��(n�>0U�Ph�{�� �n�
o*e+Ҕ�tn��~���C;��:�[28����@��vp��:n��f�ܶ"�u 5�]�Nj��he�WMj7f�r��nx��@՘e�fJF�l�&�qk9N�2��o#�(,H^���%R�طyZ�U	i���e�u�2F4.Y��{fPT�Ź�;A�ۗ����jV� d\�՗�2>��B�H,)B[�W7*�RŪ��1B~lR��ڎ�����6�z27J�� �ܵxk��l�Xƛ�YJ�O�ч s)p�p�����ǥ"��D-ؖ%��������|�mQh��4�Fd8+�i%���)�n�bf(��P�����r,�e*]�F�Gi˻� �~"�\rl�ee F�F�8>ͣj�2�����!*��u�C�C�`���)Y�j�cڬ٩딫�FĩکT��z�-�Qx�.�dz�*�E
"�r�t�V��%H��e�ɍ��oY�����ٚ�&Pȱ<j̎�i�{�C̨�	�O0<p���Vdz`Y������Lx��Bn���B��i� �KYl#��.�k)V�QuU�HYW��H��0� ��A��y�u��&a�M˂'�lf�^VF�������L�[,�)V�_b�3aYUoQY��^�/~߁�n��E��Y@H�piF� �O �[�]�{�n����E&鐨5n,����l�A���#���Cۭvp�1�������ZӔ��[�6�J�Q�Y�V�iEV�=�!1��� 1P�&᳕w(����Z���Q[$Wq��Gm��ۚ�ˉ�����FZ����F�II#}$o������G�H�I�#}$o����7�F�H�I#�$o������7�H�I�#}$o����>�F�H�I�#}$�����7�F�II#}$o������I<+������sG.�{E"M�q��ʹeVin=�SǇ��9�N4��Zn��gPe*�]�5n3%+s:H�]g�	��v���>=�	�n �w8���BQg�8�(>4#��Mʊ� �:�i�诲�VT���0��tV�N�4K��3s#��7$P��Ӹ0����N��GzvKUt�kHf��9�4���uݩl-Q�R�X�g8N�UJq�˅p}3�̅1�=���2��v���]ȋ4%_u^Ü�,I�,^#�����	�Ի�������a�f\ڦh�]�`��V3�{��sA�`0voQ� ���e�, 0�,ݡ!Ȇ�����7]FF0V���B�~�]�L�����B��n��U� ؾ�4A��q&��5N��d��v�U���9R,���.��_m[*��o�����M��N� �#��a����|��}�'�_]ei24	��ޜ��Ovn�WQaG�)1�!�='��<QT�r��'��$�s��um�)[aN�N0�"����*�ד��77�%������9ڔ?w<��%pwz*c�S�tFn��Y3�Ԕ`�e�O��;���7i�q-��P<�9Q�CG:Y�Q
P�����0s\�Y���7p�=Cq�5��؍�m��u���'֯�Y��f��Y��Qf���W�m�5���C���s�L5��'�F��u�c�;L����}�	2¶r�j��T�󥇝�˫zNo�!��M{3,�}�s�;U�4��{�W��N��0��|e���J���r5+��L��ر1�΀�h<�8����`K����3���0GNh.�b����iu��]�څ��u�y�(����X5��j'�RF0�W������Ϸ�9If��tb�ʻ�d���Wcx�h2��L+r��v{#3�{\�7�;b�P�_'����SwF��.���k�p��}��7��yǣ����go)Vk΍d;	\t�]ì�]x$�J�ʼ��ϕ��ᨈ�CH�����)om�?`Y�������}����d�uv{o�u�!��2�4�n��RORX'&u���k5�NN��S���*��-,�0h2[�܇&�V.�L����UW�v��eoH26���g5b����68A�����:#|��rc�X��6�Ð�le^<Ĕɡ���24y[�y�=���{�R�73��"�_H]�r]�>׌�T{�����1K�&a��v����}҇C\1�����0wdt+���k/��[y�Ǎ��L:�N��/�vd��Gq��-��3�8V'Y�z�R0�����R�cJ�ݧ���[�Ɠ��hӞ�u��ѐ�ch��@�*6��nt�d՚��Q��nPΫZ�-iz4�;1+1\���]!Y-Y��;��q�6H��zك7/h�)�,�H��a�r	{ĳ����T���,^�{�>����o��;(A�f������F7��tYg�[��QY*�w@G8Ǻ����I4���� �F!K�����V6A"�[?h=W&>53QWK���y����a�.���y�KK�7�H`���e���kו"ĉ�u�X/8���m�Y�V��o�dtEv�_)������<�.'3)u���d�8Ď���ˌN�������ʵa�N�����}�w^؛���hů����3���%��u����2Ig8����㔺��!S)e��>M�Ա�Ml���؞�2�6oiN^E�Ԥܳh��T'��m���t[{�W�y��v_����l��z�WZz���ݙ[Ida7Ԭ:�w)��S�n��_ʛ��7���\U��U�cl�r���]]�ƕDWt.�K˛���c�
oo]����jΌ���P\��#́\r'��1m�F��9�3%^�����.�"�d��}�Y���'�Ħ��o:���o�rIb�����NB�M��Z^���e�J�]"�yR���e�b���N1��u�+xF@a7������p�$����b@�IMGAV�2�\��PɂZʺ�Bm��Ԉfl�]w- 
��i*kp���t��/jslUI[jw]#���O���o�f���.̲(��	/!���,PT��A.��Q��n=
n9��V��=���5\�[�;ker�r�d5�ab�cy�Lhc�~x��g;؈�Z��NL�)ϻ���sM&{z�}qV���}�xu�Y<�N>�k<��%va_q��g��fgv��ϗ|��y
�Z��>߳��ҨN*y�ގՔ��դ~z��K��}[���i��X@����T�]V�b�"�w>�
�|��ř>"_^㘺��TL��M��Z�d�Y�!g�٢�*N�o�W:�r��I �=��`騫��/f��T�\{��8���5_<W5��7IB�[�o�=��-&_۸4�z�p��qU����&}�v4�Ecv�r:�$t�;�a;�l7���+f�� �R�Ł��jQ���]�X�i|l�s4<��rܷ 짘�XY��PUd�B����Ւ�掻swu���׵s%�T�gYAީҁ�e��
�\�3{�4*ܖ�SI���V.��e'֢1ZwW[�(쓉�Pòl�E��g����]��+	� W�v�#{�/��w���ui�yn�n{��l�T�MC!*e��d�h���Ex	�����K�8��y�A�f�H1�r�⫔�*�x��C�'&�QҰ��f�ڰ�\�9A����L��$��f�b�!gM�������椪�$͠��XY��<M�yg����]a��Ls���S�Ǜ/z�W]l��9�n�
n����W�)W��g�۾�GU�[+��j���T+����0u]ג&s�:����)�ہ`�7ik���3�K���{�N�F%[8�F�9�ɡ-�qӧ}$�,�P��K�;��w�fܡ	�8vk=o	�e�.�Z~Ź���58��n�])�����]�T�GfI� \�����x�:@}Y�V�Qx�l��/����(�bi�ts���b�)� yd�dyX>��w��y�E�_*�M���V5r*�Z��uy���r���[�U�J���0�t�#Sy���/B:A�ne����"t�ɪ��\�V�µ�A�Y���
�0v�z*�<Yv��{�ȡH����<��w��f'YgrE�z8K�S6o\�64T�W@\�]΂��xE���[�z��s�\����#mR3=�W��l�vdٲ�d$+2t3&��A��(9���z����t���6��I���c����S��6.,];:-tˇrB���ɚ��p��,9͛{u�[;i��7SE���&ʃ�\4�u�l��#��ib��s[�n�F0��HG]����`�Fʻ��_�ui�h[����!���WF�MӇ6�L��:{o�z����e;�˝SK/�e�xpv~䍭睗"�h�"�D���]4e�[.�� p*�^������Rw�������>oW��,�$���[:1R���3��ڬ��u�NM2�`&��oP�������um�Mӫ���O��=}��>GMD�2�WWI���<rƬ�i>�����=��#L��o&�SҠ?@b��s��{Kw���x_%���t��������mh콮d�D�4z��������^�K��X+�H)������>��{�f���g,���.ς�L�k3(캂�O���m;o8�7Зe��Z߫=���ƻ2����4�N���3�!P�ۆ3ja�����UwqU��(2�^����n��yJ��_i�yV�wgE5E��zH�ޝv�k�b-��d��%���l�Zխ�ye��t6-��7��2��'�o,����i�`���W�9�%��Fq��Z�d�S�o)P9o���Qtkt�t,vh��I�Y�w�����ؾ�ǆ�y��3&":gF;A�4���M���y�36�R��D�욺vi�h�Ȉk1�܎�'0J��%
��f��H��Gk6$֖)�}S���PVn'm�-Q�3V�'F(�
��O@�����y�lRJov@�.��������.N��|�������@�Aap��f��ga{�7�Y�J����<�=�ÛCaYh��ZkV�2�Y�X���u�k�0�/���.5��=�/���f�W��6�@V`[���Ewm�,� ��B�n!C��� Ro+A�¾�Kw����s�5���׈u2���tf�pݫ.��:L]��}�orW�\���{W1�H젦Ժkt�\�K�&�$;��b���Q��
�o�����OnVe$���`9�k�Ƭ>"��Y�������}P�#-ҽף�Sc�1Fǀvє؆_5l��G�r�(��Ӵ:���j�Y�Q6S��vf�Fg5�L�X�|��ͽ��F�Er���׷�U�΁��$�&���6�a�Nt��A����	�] �| ��W���n�1Y�B� ��62N��3XȠ�w���}�����cwdC|v�����	)��Ơ�lf��A+i����'�gg:�KD=$�
R����7�(��V\�1�sh����t��Tej��(�
�AZ��k�mX쬩����q��h�,txY�[/���H&y�+}�GX7��m�u�R�9�G{s7����Y�/�I�,��t�t�[�g�kCnX{q����͚���۳y�+0�k���P�	i�'�����w@:�0 �D|{.WL��:Œ��Tel�!�v�vt��@��x�<�u�l���"����al��.���/sv�(Bf�jf�	ɣ��)#�㽫�X�t��vEɅX�څb�}�z(�]fX�fA64`E��V�7�_qe^`�uC>e��=�wI�(f%Iɥ�,�.�m�]�B�&V����Ǚ�'�a����f�_"�N�����i;�j�'��1R�e��\U{P�yg�0����<�^k��^��`���ӫ���[�^�̕4�st-�5RB�%��ttWvwDa�8��j���zR�;�	[F��;o\\��;:]��.�g_�r=�pG���-
�<���e���\ggL�=��QĂ�U�RoG��Bޞ���Y˘��(�*��<W*4�ԡ,��[E�#c�S�W�Zϝ������`���x���FL�f���;/u^e�6��5��	fw@��M�ew	�m�Y��2N�ŉu�y�81��;"��gis"������xKު{^�fɋ��4��sd]t9QN�!���I�mo@����&AwF��S���O����^��w9�Q�g6��#gTM�^��H^�)k�$("�_h������-�Jy:n(+kAF�\�s�c�e+o��X&�KV|��ww5y�.7�b0�Ĺ��F�&�tgS��k�fD�ھ���;��Gmj
[m�|Ag���ԓr!�\J�&��S�ӷl�I*F���\�OJ9��V�ل�v�r���Y�h�[<�̷P�/0�"�s|5L����ǳi���)�t`�i��3v��Ve^d��7�%�'\���t�ݓe�K�}O�,�,1���D2�hT�Q�M��H6�/;5#d0mC�N�T��"j�6��K����t��r�-)������Ί_/����e�{-��5Ò�w}(n��<�Y8��|�����4��jo2-���qj�_��3�`"*�L�r��f`�+�7���r���5���E�О��5:L��=t�BC(g��ǫvػVu�sr>�\'Ae�:q�*�;k�������t���_%�f����h��=��'L�J>ʌ��$D)nM��
C���5���:�d���϶ݗ��v1�nq%Q_������F��hl\s���]HxI���L�ge՛Ay����@�7��Z(^bꖦ�3��n�W{h�Ku�j�W��s�ˊ��ft�y�t\���ã}|�ṉ��<7�x�P��U{��Hy�
r;��HW�fF��uD7�UM!��iK/���(��t���n�(�!��/����;���νg����fa�Əˠ���"�Ky��0�+��g�t��|�ŏ(�pE���{�g��-1ЮW�:�����82��{p��{��ZzuDJ�8��7�v-�u�/�V������vt�#O��[��q]!�| С������eh�ƶ79��!M*��<	Tʮ�S:�`%>��$o��Q�wZk�b�a2��2s����Ek�t��q��u�}�waݬ�rӾ�ҵZ�9ɍ�T�W����"XCn����)�Z�Y�f���t��Ns��8�u�Zk���vЮ6�<BwK�p���r<��"�R5���s�ܴ�0�V�枰�Et�WG��L��OZ��.��Xj�V�ZVD�kGOՖ;^W݃�A��v�2�󃋷��!���iJ�����!U��v�=����-�-%H�'M��sTt��e�q*o=�Y}��Y\I=e�%,T%*�I�Èkz������OM%}�l��+L=�&����ar�z�]�nV�^K�jV�l��i9��u��K2_f���b����W�(�����ں����Q�J�"2�Vmǘ�[�r�Ճ��<�($��*!*�q3&e�RVkk@�u#��R����i�o�m����άk����|�U����O6���v�5��nH-Wi��G�1��pB���7I�������(�ln������Ǔ��˼�3�����=Ա�O�ݑ�T"U������;f'H��z,R�����[�-��*g>����	y�ƙ*���I*���%�K��f!��8��~{�;1��|Ñ*�
^�3wB��y,����
��֛��j�f�anul�WvAN5���6��ISZ4]e����w�o��Þٽ��ܯ?�$ HI?�HO��2B@� �r�Hy���I 0���$1���$��d��H�	$��$6�HM��I��1$�a&�Ym�!�R+ �c��X�����|�8����i�%BN2L@P�	�B}��Y4��1�`i4�IHM0P�I!�k�+ �P20��6��	!�*�@��!�Bu��M<Ia'�&�!ĜIԁ�ľ�YY	Y ,Ām�,�q�$���ϐ4�oRԆ�I�@+$8�8$Xs�,�!���6�4�Ch�M3�$���^��@$4��� �8�Y!XT1l Xm�c�aX����6� �,Y�|��$!�ʕ��R(�H+!aXi��IZ|��=��$:�ݒI�&��xq�I�N!�a	�H��@��d�M!�O;eH�HC���4S̒�w�bk� �a$=���abpO�����a�H@�fV�R� ,4�b2>M&�	\��L����H��J�@�2�Z�I$�����'X��@ݵ$��b���3��L g�	'��>d ����'R��]���%a|���=�ߩ��O!��!8�8�	��#4�N3}��c����_2SHm�$&���+�b�f	$�h��>�O ��֡ ��V@4�)$3T$�XV<Ԭ��HT�HM�Q�E�I6�W�儛�25�>HLd&]MnZ��β���CN�I�R=C��v�|�N�VI�ႀy��c�H{t���Uް��@�qЙ����HN&$g����jB{�_j�_S?eϬ�;�	�ܒfPFHV@�i2�I��3��o���&[!��F��k	3.���}B����K��/P����o��5���c	��ך�}�a�{�8I��E���k,����&�Y�2�	��n@�ם�MHr��)�D�����	Wt!g��B]'���}�	�c�F�����k����~��#�U��[��c@��6��+����@��֩*k��i���9�@yHc�`�����e�h�y'9����`{V���'�oz~��3���g3�\�l�˦�0�ZYL�f��I�=�w!r��k�����3x`/{d9�����/,2빢r�����Y�Y�^��}�9�§y,>ݓ��z��W�zִ>������d�!��ޠ��>z w�<���}��wƧmٽ\��h���������C��Ls03y����b�����t���/l��{��_�a��~�����١���8�y��9�y57�g�]�q�$�L̎M�����d�{�w@wN8�N�ْ�h�尿P�k$�� ���:�G}�=���d�g�jL�>�{���!�������~�2a��o6f@i������hu�X1���̴����@�'>��;�}����!�����j�fi��o��:sxIq,-Q)
�Ino5���:���>tA׾����o�	NRc���8j�eˁ�k���|w�oz��:�_}��)g���5���Y��1�2�z��d�2�yߵ�Ht����p5l��\���hd�#�d�Lހ���3vB�ތ^ӽCF�!�5Od�޽ͅ�C2���yϵ�i�C-��:�r�0�ԛ����R<l#��G&a9�絰�ֵ�M��tC���%ߵ��ޟ?jw��ԙ�����g���!���a;�$�dô�d7�2{��I�Hf�˩4^�d�R}�7���k!����f��L��w;��hw��\3!�<��緩�w�������k9��F� �V��S����n�I�R���X�|��`�-�ff�6Ò�%�>��v L��]ίMp�iR�#�);�����$���k8F�Ƣ	rB_&��U�Hf��PF��u�^��70wQ���U�\Ne�(��������b��VSqڼ��]�:�4��2^�Ȇt\,�M���\)[�|(�v��Vz���dCM�D��J*�c)U���;�gS�!O����%� _�w�����#����L��%dcB�sGa���}o&��f�o)���͛�os�w0N���Q�8�9��+H�-�w��������%�G�\w�<�C������\l��j�����:��S2>�*�v�˷LH�M�ê�Nb9`�ۀ).�F{,L�-�Ӵ��֤��IE����i��,U�}B�5�#s��^��ü�=�h�ֺ؉��?�2A�
ٝ��X3yН�Q���v1�$ms�W�8�6��!v^��bH�a���$��J��h�]c�$.�Yf����%����i�����W]��� ��8�yxA}��u�$�k�ч���yw���7lk�2��F)V�7QL�Ƕso7�T͘�UK8�\��&��߷4b����L�[�v���d���0�z$�Z�\0�����^pt4���X����Xc0S̸���,��;Vve���I��v!��A"�{��ymҲhs�W/��K��X�2pj���$6����ݭ�ۏ>�K֡Y��[w����J*,�DBjX١\�S�
ʏ�o'Ի��oj��e���Y��
3J&�4m�p��$�����uշ���ܻ7�8��qt�H�)���w5+�HA�+�]ɀ�Z�����;�\����ii|�7�>uՌ�ѽ\MQ�a�(�nt}:"�'�ߡ�ƌ�U6�#�,z��1�l��H����S��^�����Bt��9��[��2}�&�!][j�Č|о�Z#�}O,�ݨmE�f��ȥB'��s���Yn���\g��Aw9Ll��������s��;�k���\�y$�� 7�&�&�:����"��$��!���@�$6����a1���,�ޤ��4�
�}� �@�m `c	�&2X��`E H {��~�ޭ�)�ÏĂAiTv�`�*�VAb�2�Ȩ�E=iD�E# ���b��@�&$U�Lj���X��D���EB*���\b���`�1`!�����?Z(�3M�5�Y1�s��TUu�c"�c(�F",
o}�����EUV2(���A��[DAAG��$X*���h��`�"��a�<���b�֊���NYA��E�j ��?B~��M�\��
�q���a`�QEEF�D@В��0ES,�F?�0��T��'s��}�z_����qUX�P�ET�Jc*�h(�s\��ս�*�ƣ-(�����
�?���J*�Y/�dƢ"
���Ň����"��Xʢ����O}���"�IU#�QUr��m7�Eb�سT�
���;��(őUF��1UE�*�eo��hA!Q"?��e?4c�.�~qP��%�ATX�?������>���}�8h���QTQ(��C3Ϯ��(�Q>�M���"��B�EUE��(���R�#"��}�H�5E��������r���+�&|�Mv�E�d�F}��
j��C[�ғv|�U�3��~����
��
�#�,6��y�_�(��)��}ىh]�z5>eDO�L^�������g>�?|~E��veDb�+,D�?_�����E`���*(u�P���������a������?:q�*"(�K椭CGh\��(4eTko��F�������?\qh,e����l)EQc�(�&��ǻ��E�Tq*�Z#��'�߾���ߵ��~ޮ��6ܳi��Q^�`��`����\aW,�����^z�"~����]�>j*<�f��GT�*,�*3��F!���m�#�RQ��4j.�R��Ab�}u5*���3�,�"���}lȏ�B�J��ǝ�ϻ�s/zbTw�ɤ�4�(����TDjUV.��Q�UF%��3R�UVrӗ0�T[h���0�`_YY���f�����[b�Ս
���tET�7�����wTݦ%*�%���h�Ѷju�v�9s�]�h�j�q/�J�2TH��=�2hA��*�ݦ��*�j�)~u��������?aD%���d�� �I�o�A��=���**�m9J�f8*�׷76��GT���u�4�U��X =,����Z�6�z�"/�� ����W*�a�(��I<�+�Zօ1
}g��۹�޵8�
(���w��A��
?f+�عV�-޳4�1�%��<Պ�빆�o�=�݊'���\ǡ��?}z	C�:;���I���vǎ1$DSg�S$�X?\xh�$@��w3Y�����a�7�W��h�r�pEph���л�t�MEM5�$�ibG{��T��I>ګ�5�5�}�:�<���no���V_a���sĐX
�O������w�y�H���=���}2�UU/
��[$wf�]�N�a�M;v���a㾘�n�����7ݴ�U]��yB'�-��\�w],fe�; �3�@��i��Iǘ��S��k������(��3�kB#�0���ːPƥ�Z֭�\��3���T}lb���\y��mGT��c��ZsZ6oI���Tq�|⇙�L����vi)�b
��������s��z��]��*��+S�j�+�bi�&��u����iaFc�K��
_���&{1��-��SW�aT����w9�Wg즙�fU-,�5&?�Ŀ{0]R�f\��$����Z��v=�II��$i
��,YG��Z(ܲ�z�Em�@!��5B��]**�6���8���y���ִ\�M����oJ;s�ణ�uq���8���s�����Ϸ�>�o���hE<Za�U�R)PS�j��^ځ�.�Vq�(�Q�X~��uee�Y���O��!i3���LDJ?,���<�OP��ǹ6�+�4�
?�>�G"d������b�輥Dv�#m~��5�Rh��l��x���/Z�.�b�/�d��kumTZ���ϩ���`!W�΋�ۻ�����	L��K6C/O�d�T��R��@��"5ڠ z�`�AEQc���+��Z�hT�����i��b���v��a��%��G9���o�O���9W�w2R���"��//�12��}�QqC�`܂@Ho\������ty�U�~�1���)�����M�e�������(�R;ֳB�����;����g�E�@x�E��!��ŏ�����Ǐ5�ɏ�Xdf�~�i������7rbW�?f��t���ם�	hj�5|�m�R O�+r�=���[SuqL���uk�-�(6- (��t�EoB���D�RH�B-���DY�'FN��B�ߩuO��Ǟ�/�ʕ�v�tH;M�	 ��0�mF���w��Kv�Ѵ������f��1��y��-���q����.Ĵˊ1c��wX��J���ڵ9i�U�6�:�k/S0��平a����n|}�_��߷��Ţ]f�@�Ύ�i�o:��ъ�n���Y�ZCVa�5L��I��)i�N�\Wv��t��C�oFԆ<ݚ_bFv��p�:�ns�Y�y��ş6�&`��^'�f��ۧv�ײ;��l�wWWXz�o����yO٬�����V?�e�S*��$"��!�GMK�}w��<�|�;����u� ����:(@^�K��?SW�@ϩ3h��̮�Y}���I�9�ĉ�bо�X�[��OM][��2Q�s5��z����ay�N�el�UB"=p�%,�B|��,d�w]K����p�����֕���p沩����2����"+�A�P�A |�����-��aG&�D!$Ƶe	�BrNU�ㅈ��˧<n�{�}Ï�7�ͼ��"6K��%�|��a���q#�TZ���z�$`H�-L�ba�`��,� ͟�w���Y�xR>]����@�p�4y7D$f(	����o�|�x����ƤAEx����{�qb�l�`4U�>�N`_ 	�Z��Ӳ�:����͐4�	$����8~e �ʎ[	��?^\�g�ߞ�K8����f�߳5,G�c�X'wmkS8�`�&+�l�:lR�ۜ=p1fQ\G�2Jƙ����SH���p�5��E�@�#�ڻ�i�nJJ��
D����AO��o֎z�18c���P�����Yi�j��w_fޡ�]�~���?2�(����ccuY;>cZ�1���h�ޟ�� �7UwL�U�����o5+��	���jR�!��4�����(}$�P�Ȏ0���6A��DI/s���T�'�9��꬐D�>��;�P�q��.�0h�|�"朙�L0�J��JH!��[$F�%��(~� ��{6�c*י_,TD-ɡ�����C�<ǳ��W��VS̅�T�OG1��5uoA��Ҍ�����<�.Ѵ�u3�]:�Zt�QG1%wp�w�z�u��mV��9;8WZ�R.6UF���;�E��f}������ۆS)e+BRH����O��T~� y65���I�z�uX �ʴ�)#|��W1R2��u:⮅+i`�x�l�G"��|�,��B"�$���H�g/���m,A�[�&PiD�)x�5M�n�W���[ B�3������CΣv��}��[�c_B3q��0I`�h���-!�$`����eJ$��/-LP)����ý�G�B4&�)+�|�ן��{
&��� j+�����wŏ[��Edƈ�L$k����Ӽ�k��r��sFR�\y�0��3�m����_Ԑ=�}����J����������m��|A��A����ű
!tb��P��4~Ŋ$��\נ��$N�������s�m�1�s��(���W��t��]���Q�f�5jd����M�mo�����q��ٳn�`����$C!q��6M���f9M���%Żkz��@wBTc����,L�ԅ ��I'�$/�C)
۸�D�%0�[�"x/�L�=���m�O3.��S�0�	�t\���/�z~�϶^[�^ki����֯N�U�K���Ca�y?�Q5z�\����p¸� ��d��)���D�|*��A}��<a��u�c��i9�D��F!$jFPM�.�`,��ݖT�lb0�mV3�O�$쐩?szn�׿��[ǻ��,�政i&��i��K�5�ܮ�~����9l����o�|�Tf,�����s�=��ΎR}ĥ9�	�w��q������>�Ovy�򐲠w�O�b6��{��{iq�ժg;�gQ\�k�Z���t�cxǁc}u�٥%�l��z]Ҙ��j��b��9k� �Q�6�q[�����OM��� �*�dy�.�4a%��cR~V�`��[ޤk���P�k�,�[��y����N��T	�g&�1�x:�6�����ώJ�tz��p�B�'�|���1}y�.{xǟB�>I$|�q:1]�u�����Bl���Y��
p���[�3eϾ���i�-�B�L7���U��Ͱ+B�6�g���WW��,�"|���ڛ��gt*�d,�UR<��19qm�n5�}s���n�S��i�L���0�={�c�^�����/��ju��9�A�{}y�7���Eq���j��"�=��Z��[g��~���g����=���g�GǪ	u6�A]K�$̚]�c4�X�Zd5�?rtJ+��2��p�0�ǵ&�g�T��x.��p��=�$>�<��C�@6��Y'���b��g4�>�"�l��c�U-�o�����{�
5]t�:W����i�2y���$n&}�8ׇ��~c� :�9��x_��MZ7W�绱�5���q����;�}�������>D����?(�e��)7�N��K¬��:l��&!��K�kz���<7E�r˟��ݧW�������������ʬ3l�3�y�i�n��H$�0�����.�&V�F"ۃ%}2���9�+ɇ�Cؙ��4��N|��~�{��f�����w���Oz�t����r������!�a� [C��,� RR@�.��"�E1c��� �B��tw�@�]���!�V{]9߱�}��l�B�q>���g�=S����ޞ��׹5Hܡ
�;U�svr�+��(����V*�����oUoI���T�WLN��+�Ϟ��W�q�0���jeO����-���&c��R����v�1|���M{��'�1m޶�)��{���e�4�/y|`tڳl0֬w��D�:.$AC�c�U�=�T��������B��ã�B)�������[�n��*����7͍H�f�RO��ĵQ�`���S��Ҝr3�&j���6����T9!Q��G�<sB�6.׊� C;�@t�?|:�JG�]G�\����uL��/�+,"�D�c{��A��qt����3�e��g� �!U/t�P�D�7����!�����~�uW�^su[*�M)b�# �8�	�#�1Aj;�e�ځ{/_�꼙�"��0��=�Ȑ��� m^�YӒE99ۡ?I��1�s0�6
D(
��`���"e�i��7f��kR���R�c�v��a�䡑J�P���Q?qЛв�Rm|��!�uA����{W3U�$(|j�V�f���e:&�C֓^W<h�T�ܬ�YN�Z~�MQ�G��`H��lZ=Z�f�,�fT����gS�+��Ѭy�֑5Gϻ��c!���W�V�&���O���05Zӎfܭ����i~��t.�uw����;,ڷ�xc�}X~���<�k�U3M��ް�8��Ӳ.�q)t�L�C���j�WJ ���1f�jWJ+-��y�b�v-WzLֵ��!ߞ	]�~@�C�����H�=�5cDd��K�y$�� i�~���~�����}��~�����W!e�c���-�T�
��h�u�B�Me]���5� ��ӽ���������'��Ԛ�@_wY����:�?u�K{�%��%v�ƣ������v�q�N�܂�^��L���S����IM���f�K�0�Z��z�O�m��2<a>�q��,^��Y�9�2��bl
!�ӵ]������ݕKD��v�b[�c4�!D[���ݨp���
�.�>٘��Ê��|	�tr*#rH/@��g�D<Vm�>�2������nRܯ3n
���flά���+7��u[$S �a�����Փ�T�i��G����\i����b�����¿{7���s��Ӟ㯹}ـ�6�n�(���c����[o���	tG���s-����2ɫzDUD�]a��?��r\�-�a]��7�Wk�u"L�����|*m3^ǗC`��g{u�}޽�wU@����!'��ξ����7�f����{4��=�&�H�'1���n��H�^cL��Däd��uk��N��`��hP��6�:q��F�&�԰̉�U���N_�^t�5M���z��I��y�d��:�L6��'�/5d��'�u+���(Y��ͳשN+t3�]u��P�(_����B�K�3���=���B�"jXj�)u(/�HB�5ƴ�x�x��4�o.��
���h�g8DrI�OH;������u��/�3�;�C�^�P��$���B��x�]�7��5����3��~��tQÛ����@������!�BS>��Q�n�bƚ�ɄdG3���{��s��|�ʴ�i�kė,���w�_��Kއ�)�c��[�|���v���@{�f��8��;��(�ӧ%��7|h����{�f�B�Uҝ%ܜ�\^7���7e��􉿦/R'�m��$a��y��ƟmUU���W�?*ekD��^�C�> _uT�u����O��ż��-�5�^ZV�$�D=��Փ+ʡ��;���DeW���䪂4+i��c��(��!w�iiz��(�n���h��~ޙ���R�����o;������4z�\.��c�z��cʶԑ��8ʙ5Ҹ�a#p,����4MֱV#�߮�0�,	�\8C/�L#�]%�ל��k��tͽ��ZeP~+�,.�i�R�B���,�[���3�t���1��i�|ΰlT���>gh�K���xc�*9Z�7��0yמ�/ �7B�'�0P��S��ۆ��\�!�Y'/�GӲ��7�G�n�L|�ʯ��֋����s�c5y��� �5Ү���,,3|���p��i:O���Im,��j���[����6w�"
i_Wa-F�i�`K�E֕�=�!�7M���z���0W�HC�5����w�͹5m^x�g�ސ�!>�f���5���n;9t��jo�kYݸ��y����C��g�j�Q�܋��{On�)��>(#��K*ˤ���5�$%h��>��({ı�Z��dB�C�8:=v�� %��n�����Yw�����k�پ���o���� k�̙l����k��������o���9IK�k��(D�˷�����#'xKl�	�QL�pS[�³pp)C!�u�jlV9�,�`8y�/��+/O3�]6��*�B��d���ٱ�T��BJ���=Uk��]}��Pʘ�"y�!��{<�~��]�!�z�Q`�Ϻ<�a�̓�[vuЊn��bB���tc��մ�"*l��/����U�c`����YKH���/��j�B�#o�)�ȵ(Gx�W�	��*�q�0[���6r�SA@��<�&��1r%�k�����f�~L�����o<l�_e��wH��I��$������szЩ������)����BYe��3�}�>>�<�W��<a���}�Q����dL�<rA��8.�t]dXG���hs�y���N��^0����^�h�� �)ԙO��k�j�▄�$x./90|�w}!���Vj�pd;���;q��j�bm�|l��nFPC1�b���,5���	J��M�A�a���`r�P`�J˽3fY����N�$7!��V9��w�_�yW���m�%�:Nqc��Tdꖜ���ٰ�:���sТ��!~~��X�ͻ�`��f7�zi�n2	"����;�4�w��`����޾�hiӓ���׈^w<�����{\)^|Y����=� �<�2.o�rA��a��ԇ��z�*-;(�{'���7�O��Es�Wϝ~�
�M��������8��R��O�_[�G�.�ۡ�|�o���DV�8��B���i�V����r�ڇ�1�nۣ���	�J�,��b�G�7�����W��y:K�3	�f��p���6���ԉs�ݫ�z�oW��&rIg$>�5��˾�,� [�vՊ��M|�:�cPx�ϩ��zpk�<�CA��gtư���w�$KC6�ELߠ��u\G���z��A�NR8H���)�v��pP�����cx~��������n+���y�����2�6�Go$��Muu�����v�lB�x��O�H�����t	�~�ϼ�Q"��7�'�0�&���NCɣ��{����Cq�l.��d��يv����5��7��rW�����3��]�7�x��֪	����$>���K��V�#��:{����k�W�����l�4�W��.u#H3ϨO�������������
oY�	&��W;�����8����M/ �S���M$P�@���џ!���1��6�ȉ<��6��vK˘}R�_�k�cZ+o��G�ת�Ǌ�b-���?>׺6�-k��BIςkfM�ȵ�>�����d�h���a�8շV�"F\�V�
�R>yyF�A�ɤ#�;P�D����}���6m�[��&���+�勭Bm��3�/.L� x�@�7d�F��aL�Ҍ(8:"�1|��X+�Z���w2����ڣ�F�q�pt�o�6�/U�Ӧ���s<�U["O-Z���]�yػ@R�WM����&,���p�P���UjP�@�����4:[gNg1�/�.F>�|{y�#1d�P�4�����т�B�~�Өqi�D��4�-�^�)���&:� )���i�l��F��v������	5Ʒ[���3���E��<	m�'�h�[�8�K�\տy�i�f�|$��X�a�jJ�Yw�p�R���w\�Wё������o�wZ陣Ac���{N��e��X8���%��k
,��?���
S6z֬��*/����v&B�O�Ĵ��������u3*խ���p�(�5��_5�ܬD�:�f��wԨ]�<�o)��e��)��w]�5���O[���j]�Nz�a�z쯲�3w�e)1zj����8��:wA �OWЛ���C�S3�I=�1>̇�.m�2�Q��a�.�K��#��y`I#.�_\��K��Т[��9��=/�2�:��f�N6:��$��ؾ��ˬ�i�4c�z��q����P-��M �\K:]bf^>�;Z��u�yKM�M�WgP��rҠg<�w&#g�Nq�/�������e�N[��������6kz�:p�6��h��d�r	բN�2���,�U���0k���+��5uE��f��������Nz�K�:,��4k��:��P�S��:ʦ����{�G�����F��^K5�[lв���곛��_6ϸ��ۯh���C*uU�]�0R|��v��2�G��YYmq�֊ނw4���H��qwv��7�3I�W;Y\�Hڥt>۹���VO�s�<�H}�ǥ�$�+�,u�4���u=5O����iS��H���y8�j�B��W�~�ѵzg"��j��mt﷋��kw'�D�5�b�ˋ�hX�٤��=PH�N���4i�kqwj2c�Sf��v��C��}qDt�S*pM���|��Pq�6���*QZ�+�Yw��'+2ӥ���wV���n���ɰ�m3�-K�FHIǝZ�Ѣ ���'�R��5��� �t�{W�;���skN ΆV���r���)c[�7�����f�t���\�n�̪�\]q��&U�Y�s����YY2}g�8�U;/<;\n��`ë�A�X;櫱��V�b�*ؤ��gQ�ͫ�շ�o���2����ڗ�(��ھ3x$k�w-Éژ�|]� O
�S:�b�'f�� �
�^T���&�t�S_3�;�4õٺV:;{v��'M�6���ǜ�ܣ�o%������%��X:ɔ�U�SH���[�EQ$v�/k�[�� �;1��� ;�-M��i�yi������Z�;�g�q��3��΅c��춚r��Re��A�*�h7�]	�]·;��B��;JsT��.>�����T��!�Xu'���5k/*�X�8/�g�i1��*�1����	��'S��Pٟgc*9�a�����I��O��2!��8���!��r����r����\ٷ11I9z��߷�O���*u���R~v�1!ߝ�C��!�Iv}߷�&�3�ש6����i�I^%a�<X����Vg�4ɤ�T����q���������3L�������>�c�>�^vܩ�͎X�vҍ����q�t�O�'yJ�CL�߿jy�=}�>��?��E?�bm�J��+:�@��M��XV��4��\CW��M��N����m�N1˂¼/��M�;d�R���!�Sxy����N�[+���־���x%`�i����1���Z�ϓn���R�]e�c����L@ճ�3�d�6�p���?���*n�>?RT�,1��;��h�_�����_$�Y�Jw��e�����7��?u�P�ba�Z�*�C�p�8�N0֩6��ɉ�CZ�����D��^�m�����ѶVJ�u��>g)4��G,wM3Hi:��l?�~޴�I")"*E����SMg���|��*���`=M�d�26_jUs]:���&��f�pt���';��a�Tia�<������ұ��>݇�v'PP�������$����hT?�LC�~ށdį\Ci��֍$��Xbv����;�oԬ1���!�̔V�9�!�"��X��1���%�f80�R��eOb.�fٌ����/穟�P�I�Q�����f3���x���d��'�X_�lSn�� cs'�����2�!Y����a����+�����'������Ns��y�k{��/��1
�߬�ݒ:��8�a��?��s��|�7M�a[��:;�8�)�i+�4�[+�4��Nj��5�����0�uG�*V?�{B��uXW����PD�&~"F?5�ɗ��#re��_��d���m�~{��Y���>v�V����I�����m8�鎝I$J�,�Mr��yI��P+��\�˦bbc&[�9�bO��������?������`bҔ %�c������q�� h� ���=���Ǭ8��ȵ�����?�s��@q
�����:��6�����x��G�h������`����̆��Q�ϳ��C��C��9���n��Xbu��	;���U��?�[����}������*2����C�mnqZq#c���f�FHr�c0]�(�����v����n�Q���$��e;���z宏��ٲ�s�\}כ;��ȯ������Ρ�W�	���	���B@M򃔙�L�k�Ă�CI�����aĕ��9o��b=����P�J��>��+�����٤�?&�IgyM!��
����5�x@��5��Ԅ׏}������E��|�O�m��ȧS�N��<�?�$�R:�K��4�d*T��~M�~�_ְ�߰H)�Xc'�ŋ�X�`H���Lg�gl�?;�/��}�|k_so�/�bf&�i��k��Vy'�8٦N�18�g�?�xͣ�kAXq�d굕�i42�3����6�X�M�7�&�,cd~�O�8o�����B 8�#8PS8׹�>�����4��݌��b��bkT��a&\`���>@�6!��>�C��:�e4�[n�yI��Q��&��*<���m1��r��	!�x{��Z�e�{Y~ˀni��vj\U�^� G��0(0�HO��80��j�O��b��Rq�8���P�aԾoY�fĕ?'��`zӆX6�9f�Y4�6��?f�ݐ��6��Ͻ�Mr�5�����?~ϡ�-�������3�m�.��r��>��m����51�Lq����2}���b�0�&� ��LN�jq�+<�=B�H#0I^%���� ��x���`����ya��kx����)נWw�3O篙�,�}n	4��c8���h^$u?�@�뎓i�Tܸ
d��wHu��a�+������ź���~����7�M��B��P��AC���߬�{�9�g�����:�u10C�6�M���d�q8�?����d��q��%a��4��Ca�mY��3����
���M�Y�侤��L*y�����Ѐ�Q9��m6�AO���r<�at�,C��m�n����B��; ��~0��N?'��Xu�ۼ����/}f�'�I�]��~�m�����?��1��;a�����:j��~ea���y�	���d��?�0���[g�S��<���f���}��� 0�|�^�����v���=��q����0I̳L���������I���߿~�9�SC�,Y��CHmS������͌������i�'?��e�n�X��T�{5O�����4!i��>���8�'xi���x�\������`�E!
�Q$�w��}��o3���Z�ý^^n��G �WJT�-�PV��,t̠��՘���:�	4R��������{�,���X��Wم�T�i��3x���Vr5z��ʯ������G�w�l�>g�� �?��d�Av��
�l�L�Lq����$����d��k���C���Z���3h���LC�4�'��bi')�nOfL��La^"���t>�}�~���7�|t�6�q�?'�C椎�̚@Ef��c
�\�g�����5���'=��M;Lg���
�'�7Mo'�s�L��+�K�f������l�YRT��][�g��T���^i<����`��o� ����u�T��i��/�횁Z��*}`����=	���q�4s��ۤ6��'o����oe�ĜnP] k. s�wt�w��2�=џ8̋�ڼu-v��igor�du��g'����Z�]^�1�3?�l���+�����h6ͤ }~��I�YS��.�X�k3W3�
�|p�r�=�ǁ�0DBB������W/{���'�5S�N��1MAܥ�ٷ}uhO="-k�1��T)��tK���=T�!�	�u�-|���m�������7�Uֲc&�DC�����i�G�k� xj��0�/J᳚8M�-z� ��(7���"�ˍ+�Sa���32r&p�+����p��Ӓ�C��e�ꮑ<�����(�[���t���1DG���n�[f?>L0��B��C��}7�O""sS�Z�(2*������ݹ�S?0��B�������e�l�\���ᷮr���c�T�~`��G�%�pe�i�<_��)tu�c��ve�˻��*楥����)�>�%r�&$��s»٫�C�,����g�?Xd~ۂj���;�������v|�|lZ�R��	P���:��f��</��*5i���l���wN�e�%fa!�|�z0�#��Ĩ��Qr�����8-�UܟN�w+4��]Ky�����\�V~��-�G9��O�|������B#��Ҡ��f'�ԏz�Tt��8�q�j�Z��K[�N�:ݧR��J8�����f��Lc����E=���̥Tߧ�)q12 *ο<���[+t�⭃�G�u,��q������G������FY��N��M�LK��RT�{��w~#P(y40�^V�煨��v :T�sV��`�7�]���DB�������({�	��{�a�3Q/!˱�B+Me�7����)qĬ�������˙nE�U�o�v]2mU9�m�@�j�mؼ}��ɴ��C=����a"=���-���ݐ%cS]�$�B���E�]�3olW+���{����4���� �m���*S��UGF��Jv��u"��YL�0e^���$�4e�]c<X�FrU�wpX).�&V9-z�
(�-�7+s�f�j�}ծ0��߼=��� ԼawM�5u��8���g��,8���ᶧ��I��,aZHVzH?�a
��oٓwW"y�J�k�"��#�&'�d��ig���ǧz����r'f��<,�^ۈެ��YX�c�����f�}A�ձ}����=9O��0����wȹ�UP3������ӏ������E��]��WX��������?T>��޺��gU}�_�(�c���2�1��Ј?k�J���]�U�OW압4U�}?	���(r�������l\���BƖ��.��n�>��yg3��
*������n����T�s)&f�V7���n�.IB�Q����S��d���¶�9�ESX�)w;��8�5)]$뱱�{8������������'�{�T����=� ��N☒�ϭ-�m[i�nN)^]b�����T�I@��-�U8�q	��ry�;g�n����F�Q�t���,�T��{�f�,l��MF;�}|l�/m9���Fj{ꓯ�Vr�>b��W��2u���c��)�i�B��z�_�on���������2*�
������lc�r��|��TZ�U��Eɉ�S��N�'��Uu(�	��*�K<�<3�vg	b�P�8��.��^m�'tk�M����s3e׎��<�u7��n*�CӐf�5.�*��)���V1�?(�[hJ���E<�K9E��shQ �^��n���[e~ݙU=��Ƌ�3ɮo�b�B>���-��'�߾�Wx��W~DK��9�
	��!����o6uٽ�x�jW$��0�ӥ��K�]0G������,V�Tn��o�a�p�t�k�+���m�X�6��mrP�c'�v�ᴨ����跆/$wl���.$�7�<�S\>�/���mFW�!#�"_'�/��`G��҂��˶m���{���v�=$��/���~�ջ��ak�M���(�y�Kc�ΗT61�>w�\�g�]�JM��U��iMEAE��H �Ed�񨩪�w����vc��2aC�L9�1��;	F3��4!Q��Cԧ�|^�o���^���5Ik,Gy��_k<c>Y#��0�YtLiRU`�Gf=����o_?jg��9�Φ�.=ܗq;��^���16��N}m^�&2ڳ�D��ǡcm��jb]�P�^٫]v ��� �ďǆH2�u��l�k�+���}����c%���܋P����M�O�'��Z���a��J��X�o��mȕ<����=� #��#2&�t�r�f�l0��ƾ≉���ޅ��_��.Fe��Sd��jf�#^�~���Nl;OřY�)Nc����BN)��~���ƚ6{���ғa�~�=i!럾�i��|;e�!<�)ێ ꃰ�~�a��DA�ݲ��"sfe��s�ܟj��fƲ��A���'�7)��o��Z��&Re���ڒ�%!�/k���{�
���`֮ݸȭNdh:g���t~�ַ�� ��נC�_�̢�S�>C�V��e��}m��˝�t�y#7��c��0%�b�;�%q����ԡY�L��_^����r��.��s
��J$��>}�5t>?�5��m����n���L��9Dk�o_��&���=�t���\Ϝ�㒙ض�%�j(-�=M�I�1!�C��/�yW���������
Y}��}��"K�ـI3�r��R}�K/>��u�%�kc�����sfX�jD���T���{h�x #� 긒��WHrOs9*z�~�:�u��֋$J)nґц#�q_���7A~��^��Y�w]+1�(�:ɕ��ѧSKR����"�r���n�!�}J������#�~�,X��g���ֺ��#q��m�=��ﲆ��A#F�����1�뢈�%Ϟ���裈.ʫ�
�R��ˎ`/�˶�9ج=��3�M�"l��;��.vk�=(,����S�vN�j���f��+ޖ��(@b�r�܃�ȉ�$�(.U_�{�@�b�Q~oN�I��\��A�<Ҏ�
�q�K�R,���t�{!�j���iG�'�j1��u�-n�th��e�����뼓t�?k��'=���MFDr#=]���j�}:/]O��L���&����w��M�ꇭ�����6���\q�'�*���2ݶ4:�E3l�G����S�[ŭ��o�Dӕ�ʈ.�UH�>���}{2H��u�`		U����U�Qg_l��[�N��N����F�^�߻'��f<܎/��M0mY� �-�epy|m&�]Ҩcg����e*^T�5*�.��Yن�c�{;ZlBb�{��]�r�W�d�$R�7S<��^�Ch�J�.N�Q��"a"GQI���ի6��[S����N�(L��a>��4/�P�����]��'�4�(�5�%��L�E�c�s������dm���,\�{:�Q)Jܩ��{5P�C .�]m�AU��mZ�ү)L��f���8���z����H�{Hӎ *�xD�ެ����?9<�D\����tf~(5LdƁ��w��8Ԭp� s|�}�*���y���"�T9�����쑓9������>mP�����З{,��%�y���XA\Ƴ��ڳ
�>U��.�)�2�5O��b9�'��u�
�wu��{ku��;�-�yy�w��|��ێ��e�/t�V�t���\;����Sn]�ٓH�|.�Su�g�,�P�q��d�z�b�P�?k�)����{���:��Jힲ��4�����c�,��t<9=Ϻ^�};��o��.U�I�L0�gp��E�d�P��q��'<<I)ߤL1O�K�G;��J���B��wt�Hf^���*��%�߽�IéU�߄�Ԙv��9�c������)CH�M3�&�n���T1s9E������WZ�4���^�k���n�!H�׻�s��:�ws%O��[Wb3��\�z�9�ʼ��@�&�ub��);v'�)�+��5��]M��k	�gu��
aqĠ�7hU&�����G��~���OUm7ů��7���r���g#C�#�g���z�2�nlsy�����7�u�a�e"��jsX��?���Vݢ��d���#�s�?YB�e��p��˒�"�x�)�bJx�Z��(�I�mjrI� ��)�� ��:��0 u��#.��mprr$!�0�&ju�TɃ�
g*\�"�"�A���C��C�ݓ�C��vE�{��w��7����մʐ�#�r���n\�c�Ǖ�֕�_���7.jl~��Z��S���/�/��i��#�����}�䍕]�2�v�xn
�&M���~|vsPs�L��{=/)t$�(:Tʰ��&��Ҭ��,���U�'��s��D:?U~�/�� �A�����ޥw.5c��Zx�R
?>��A�����^-�$���e0�Q�3�����g��k�}�e��}�p;�h���w=�t(*�Q�:>޲�QA�|�A��!�>0�8T�u���-L3k�ܨ����V#z'Y��U��(0�يdu���|�d�5�C�b#lky��ß:�Yݑ�o��o>Ю�{���p١/��y1uwz3�ކI����R]ͥ[:}�T�R���� nig�ʞ�Sv���D���u=�{��0Fc�%�0ga�ч����d�M�O��W�y�>Ho���E��~����Y��p35��r��OZ�a��4�7PP����~�D�k$&%wr)�C�i����y��_����fR�}_p����}8����3Z4H��"�Ik��d�ZEU�����p��zA� ��@�'��Cv��duQ�'�d��M����t�6D0-��X|�L������̠��
@o�I}�5]����1������r3�D^��!<�d��Sz��u���c�~���8K�.\*���A�� �0�ZA�1ۉ���PWm�P# l�����U߿_�L��G��r�ʡ�V�P�Q�CK�n��;�͔%�[{mvz�Pa��X0��zPn_x{בT��2rʝ�v���ݢv�^f�h���AQ�}��P9�Ǩ���&KU��kϪ$)����������.[S�`��<-����]{l%&d@,S��C�]4*(�t2)U���~�1�)B0�_��$浏zWj�<��!.��&3�WHL1�~�jR�����á�$���J�?k�sҊՙ��N�;Ȕ�W�궴c����(�֟;����w�	o^o�տ]���rm�/�ĵ�E����V�p�j���Ք SX����VZf\��)PA���{7v�ƛ�e���|J�ʦ,4�/�N}�s�0�e����b�ϕ�[��˴Mq����VΦ�K���\��:�Lǰd}Ё�ۇ��ﾯ�����`�o�櫫�}Q�>���O�3;���pc��R����׊�u��
�\�7n�dVIٍ�� �5�,L�*�� �vVP�KT$bn[�"��$~�Z�7�_�T���%�������>�g�kkyr4^Qx�Q�B%�b�%��Z��I��{��{�bH��̍���|���i���_l��U����\��ī3'��`�]����g���ܺ���"sfS�-���}�
^=j��X������hZ�6��G/Q2�s9��V�MR^-�?Fӎ�ҏ�dȸ��!^qO���5��]k�,��~1ӳ˪�p�6y��詼�h����SjE���Ե�p\�&���������ڊ���&$I��M����U��/6�U�/M-��׮q=��^Q��#���Q�����:ڱ��M���Ȏ���RC����N��F�P���VGWg5\`ƻdJD[��`�������G�-5����[���
I}E��>ߺU�Zʒ�d�zg�}X�R(.�T"�ڀ��w�5��1"m�KM�%��C��WZa~H�D�en|�3=Dd�[����=#Q
i��M��mIb�@�T�����U���PG+��oI���wz@9n����e1ޟ��^���%zc�"�R`����3I�H٧){.ho���P� ��b�֫j��嵯�+�����V��C:95���Q�q�4�
a��>#UT:9Վ;H+Z���dw�6Ƚ;�t��=NTb��oϷ�.�T\O�Қ:A��צ��uwV��%��G.��uyS��T4�9<^�D�b��?���ܤ���ֹZ��^��oI3��h�y.xs.�#�hk��|�������cy��7�^eY���ӓ)A>�}�Nޗ\X4����DN��l��DD'�n�+Rw��Z��Y�4H��c@����m֍�t�bW3g�$�4ֶ�	ʘ�u��ˮ���N���
g���Ҳ�@pü��0^u��ќ" ��L�����s)R��rL_q�$����֝pl}�aCZ����6}�oׯۓ���!Y�P��q��Yoηw}�㶽����ۼ:S���@]��d�	!�AH���8��X�b��7P�X*�ph�%�݆)Sz��\�h�p
B��e��?��	Ѕ��O�g���Gpz��:��kǷ�m�~�WU*Z-&x�	M	�	T�պ�8�Ց����Q�e��պ�L4wd�">�<��f��4B���y ��Wtkz�QRw-��$�/��0��E�:��U��o��<+l�B26ٽ��dd�"ֺLP��L�=�!��
�"�Q�Tus.Bڊ.��y��KdA���Cm$��腒�Aԙ�sl�;�{r*=�۲P��N�E�b�&n���Ҵ�Of��ѿ��쏺6ߤ�����=�Ϲ�;�8�oc��]N0((���=�+��e��T�]z������VM�NB{Y���}�C�s,�c�@ԋ�(]���jsV"�����ÿ����m�'+��{-u�u�ønq���S[e֒�[D�DZ�������
=��.���l�[����˙{9D1����NL�{�>�[]����=�w�1�D�|�e�Ԃ�.��HZ���R+o�.w��V�[�z� S�3wu�_D�5��;�ڡ�ֵ��K ��C]�b�m��3U���қ�uз���:�Y�'�)�Z�x��Pq�z�&.H�uҡ�-��Ubr֐�Ct�ǩ�����r�4&e�`�][��q{ڎ���DK��A]*\Y��c?�����{� ;�`��eǎu�=�z�±I���^Ж ��aS,:ୡ8�2��Wqذ�ę�=��y{�H��+f�o'm>�&�$��V+�w�U����-nͽ-33NTgV+�����tNqf{��9���/�Tvn�oC�f&��v��K���b������l$�9P�Gw��)A�Ƀ���b��]�A-n�{���n�hvp{���J�'ҳ`��V���#@�7���p����Ƭ)A\>;m�V%��C��Ϸbl�V�4�2�g�+[�V�ݛ���89Ƿ�Ae��GE	�Ǻ���q��� z6�������q���o���oV��]���<|��WV�����.-���/6k� �s�nL�\���i:�,����H�+"ol�u���u��Q��?@��u�2��O� 
�0��(�\Uӭ����'P�ɩ=͓�
y����ߞ��
�Jn1��~��~U��� �;���4��ȉ�����}4�>��'ݔ�h�;�7J���baJHU'�^��܍Н*���0 ��[h�M�D}hŃ�\�`-�i�o/*{$��b>�.�X�;��^jP��2�9�f�7�wm���.�NU���Ҁ�P�o?J��?uO��Sx�v�f�����W�$�8�3]T}'��َ:N����Ɗ� ؗ�y�x�A5��F��m�!���藑>�m��$��R��[g�Wo�srq��N����Z�0s��3��
WO�h���2��jz��h6�y�<��΢��ǡ�թ�5�OV�@�*�r�2�׌M6aJf)z�P���Wwĵ���㒋�e��>Y�����Q2�1�d�Y����bV{)�X��7�Ϯk[�	�M@����r�o;M�g�U{?~�U�/���	jy7�e�w�mm �,h��jsUW�T~>�e_\��"��L<��v��Q˓9��b�ۖ��$g�w*�o)@//�(BGcܧ� ��<��?zEE6���X�S��Oyi��6φS�a�1C�4"4E���jl�.��*�����UD�[l,=�����p�ٔ��r��\���u =�}{9��L�YV�0.��wI���	u�4�k����[1����aYЉ4k+�TCw���˴�$��q��N���HC_��ۣ|����� �(q�A��ߑ��"r����9�0u
Lx�����z����+�^��Ff�T�ʙ8{���p� �*�t�KOT�f�5�8�b�y�IL?�+�-�^��щG+T��<f�	�O�<cCʕx.�~��|�XܞE����Ϧls�=`�}�]NY������%����z�� &3�%׶�V|��QS��/.F��������@��w���a�����<5ꯄ�,�mɻx�w��wP��?�ԫ�y��݂=��(��V�t�u���>�%���
 L�l�'�ܛ&d���NS��)�l�K�z�4Dѐ�6n!�f�
A2��k��)2�X�.��,�Y0�{o�8���lM�K��Í�J,���<��ͧ�~���7�ҍ,oN1QU�$2�%$�ʺ��j�b�A��^�vj�+�r�3��q�B��2}S�$aB�ʩH��~Q7�
�A��f�f�m�p�,��z�%��+&Q��2�7 �6����D�ޑ2����1NsD*���yM,^>�z����i-3��kftU+�� p=%�9��vv����9BjO.Am�l���T���|�&�0s��v!�eR̅�u&\��m��m���N�}�Iyh��5V�+�N�	�E/� =5k�r��'Dd�#�/m��&�tŢ>}ց=K:�f�)�1��v�f�}1�O.�weu��	�g�j4�K�}m��yP�U�Ѕ�;^��^~�s�& [b�_� �_�'�ȿ~��ۢ�Tz%�.=vi4�������8js���A�5�$y�]��.�\Ct�.!:ρ�<\��B���I\;�TFJH�~5F.�}�}}�y��sL5� +Ҩi�!���P��`���p�H�Yх�%���J��'�/~����{l�=,��u�(���b��L۫~�B���~'��ǝ������tN���YOD1����]+l
�����#}�d���WO��bZ�6��1��$E d�[^&.!C�D��O���D��My�B6����]��.��'���e��I$LM�ݖ=5w��^O���;�a�tˍ8�DWB�x}q��]1����4�o�_u�Js���(?함#�!n5�(7���+��j�N����^Ψʞ9��,;��1I㩶j=�7�OaQ\Q��B4�6�ls� ;�	a�"��M5.Ӥ���R]\m�+Ű`��h0s.���Crk���v������s��Z21�&���K�v�N���Jd-�O�����(�s�$����{^�k�R�	E�xi��]� |�LBb�w����6��@�]�B���Z`u�*l�f/q�W{�����̳���graN� ��O�8�����c��f���r��`�J�6���Quq�L=�'g�6�og��*�2f�f��_L:������ڇp�C������޷u��l���ze�l@�3�~,�=�%ї�x�����1�F
�� ���[ܭY���Y��	�q�e���w���~D��?�"����ձ�js�)F/ R�n��RVaO�^�6��8x�-�R��f��3��w���0:#,i:���2��L-�m]�u�{�us
�G��hL{��^Fڨ�9G�<�ܰ��P�����~�n��A*��0�sx�̓�>2$VjZ�d_:T}g+�Vx2�SW]�=1�Q�v{(�����q��bx�~OQ������>�,u׬���.�E�'r�5|I~�y�?�}ya@���&mBk-1�Qug�boL���>})�6숤���z�'���o�5��*���424�Q�S�������ͻ,9�̝�@�cyܞ������8��/s���	�>Di�b+����Ute���\CJ�: �9�H���s��u�=|ܼ���y�� D�J^�Qm,�=��5����Z���pC���z��N?Z��
��NF88��UHSN�.~�|������x[}�I ���^�|�R�)%6�.���tr�@1@W�{v�l|�QmU��0�h/����r�50�1�B�Yd*�  [I�և���v���ߌ��|`�<r�bF����K���)VY�Zs���L��2���o�θ+��b�|/�Y[W�3�2=}n���7�����e'���|�2��y2P��Ѥ2+��W��!���{3,��>��������ȱ�FHpe�	/�b�m�~d���TM��%pɨ��1���3H\4E;��e��}��r����ZZ;[��{��L����]���i
=2��C�<@G��Ӑ��m<ѓ��S��|�ϫȴ!��h�ۘ[x�[���L�+�x'\@��{�C���:i�X�EnD��;���L��I� ������.���9ZW(h����"�??M�ͣ��*�I���3�=�����$_�W�z��X��MV.��T����Us�)���6M62�ht�W$��ݱ���cT�zk��ٹΝ��S�S��W��̃���E�f#�1��Α��
�nXڐ~�m�1�n�I�.����L�H�<\T����cs+i:c;�Z�Lw�=Lm6:7�O�-�Y+�ɦ�%��tK�p�޾|�����2r.4`=��ӒE4��SA��@������v��'�z���V�Z�,U
�R
�F���E��z��i-c�+r�w�[��F\xZ�&�����a�V�S���@,6��u����@:G��r�����G|V������ng.2a�<p;y�[r����w+�_*��!՝�|�,�^��\�ֵu;��S\Wz��:�]��k���]�˱�MV����!�C �j \}���c�q�Ӷ'Sys0REe5;�����k�./����v��x\f��y0͒�q	Z��;������\��J��X?5�j� 2��>A�ן�����s��f��L�>�I�����E>K=	q��8�HƏ�B�8���E8B=Hx���qFq��,��۴=��V���
��92�ٱ��S����2���̟���W����@`��WC���8A��D��h�eKD"��F����L���˰�GV��5L�L���/��,.� �h�$X*�~���y֛����� '����9��>�u�{���o�u�n~љֶ,?Q���OyK�H}{��X2��W�х�?\�Iչ��Z�S��2�b�,����s����VH��P_z�B�V��r�Z�P�FNF6["��Yyn��=q����쵋H�����"�s��do�.�pBNr<���ĪQ�p&�<-�����Ø���1N��z��O>�*�x� r�R��RъC�Q:S�)�8J�1��:�W"��7{�������Nh٠�y����7J�u�^��*��2�3��v�R�:�*�y��[��$�� �u;�5٭�&1γ���d�c�>�{8>6��߬ MF4Mj�F�X���g��4��K�7\+�r(�0����h�9�����wڿ"�R�ie��,�#�?��X?�Z݉��OO�5�d�����!��%3�i�i�ń���"�b�,�Q}�����*)$�����M$��}�]l�:'��36�'J3�Q�����B [9�G��kX�:�����\���(��dy6{�B�����ڵ5
bop�i��kFF�m���{q�)���Q;�$jtEH�p��,��i�����h�9����U�kk|�s���g�&S6�Z4����|�����"�F&V������ÔAS�V�,��1�tN�@s�X2��Ț�	�wk���V퉤e0'�5q�7[iJ!�d�[��C*��L�)��@=>U�]Hw����H�Q��0/X	���>tm�E��Ixz�멾�a�3�"|�r��j��EU@�����$<6T��;��xȇ��6�'��F�O����n(.��n�}�����+��ٖ��1&��W����C:���HzOׯ�k`�X%��e^@Ԗ���җ�;���d�^��+��:r��\�E[{-���4�J#C(Ѧ�'��ѡ���e���!��!|X#`ChS��c�}{a��q��sY	T�ou[�9�A)k�l�R�x*kj�tU�h��vvc�������ٗ�$�z�E�p��P}X2��\�+j��v��Zx�V��*�K�|j;N�z��G\r�y��S~n@�[�tn듉Y�zp9.�xVӝg��l�6@�U�
�x��ГL�o��lu>�D��y�F��}�w	M�`�NР-t�v]�lB&�U�ߡ;�u����<�^���Ŀ�^̃w�{�W���Ջ&����z$�Y�'y�7��ݯ7߇�/�����w�[}&��[QWUa�0uH���V�����Y]Y��F�)�ǈۙ�Zlߝ��v(��j��>�"<�N��'�v-�͋� =x�e��x�5*�o���Td�Z�\z!E��>M7Էl�I.d_��ڨ��f]Ũ~͕�����@W}5w�^�4���:�y��>�56O�V�t�6 ���V�d�����a�!9�F:&��1y��{�;1��u�y~�Q3N��){�1��ya�>Y�R0o�����y���5z��oH	�J�P��U�zZ���Q�7h�r��'{0����f	�L�X�9����.���3�����;5��f��w#���2Z�Y���;�I�4̠����u|s:[����}�Y̘��I��3&fE�}�o�5�����Ʈx�~{�]�0�����Mr�}۔q�	vy���㵍����Ӛn&�\���&�IS�B�~�9a�w�^W��q�J 1�"2D���!�无n����p���m��=d]>�W��9NK3*��v�⥋� ^��,�t3��p�&f�Pځ�-\�Ċ�w�1}��k��)z܏����R�A�B����U���R���N��o�b�����7���/���j~�ܜ*�([�?&�uunT�#�����m}�ja��&c�e����;�J�2�U��z���-�n2�/���?��sj���|�wR��ws�>K_�1ɀ���#B^^,�k�TH�K6��Y��}���#��V�H��*�~��&���ſ��Qՙn�~�6bM�i�@���[��8Z��x&��P�k�P챢�Y��m߿zq���֮�g*��~��t?��r�8ݽʓ��Xˋ�����RT)~�s�s��rt6�;.�1�i��C����2�n6��o�*>����mي���#M�Ҫ%,%ك��`-zžY"��,��TT�1�qW$�F�	�7�,c]�J���܎"Ι��<!TƹS[���Sm���Gqͧ�"�h�QI2���M�X.�����o�����.oO����+���
џ70�E2�@�X���������m��.n2P4���=����.�My�<X�nvun0`�c��Q�;�Y��K����1+o�)[c8)Ӆp��^ FU�2�s{��u�\�ŧvw2mr��\�퉫�մ.9n�G�]{�����j���Ŕr��	T�u*����w����k�g�_��{�ys���PDU#�:�}��fj�[����^2����~�7Ǧ�,u��ʚM��ӳz��A'B	"k�����L'�.~���7;`�]����t���wCR�:^EdPO��	�<c��Rt�Ф*$O��FGsnc���o�>���wz�S����~~�T��nc#�����%Y	�����1s�Y>�&����d��}�o���@���,�����]r���ɑ+yX^����<�8Z魽�6aB͟]*y;�K��-K����agu8����6.^�lP�n'��ke�޽	�����{�6/u���3>��g>�����Lz
�WA��6����n�Q����&�+F�Z�@���OM�i��en��8&�����c�n]bڹڐT9�Wd��Ҹ��=�I�@��Z�3Rws��Jh{ׇ�p"!4��Q�����wlo]u' ����Ԋ[g���7|29���?�P;�>	f�Ð�[�
K;3&
^U��[�8]�x�>/)��YR�jp�sx����L��Y�-l���)�f�p��#��P���ʻ�-��VƆ�_+�X��by����^^k3�ّb�B�����岐,k��z�ㄥ�gm#Pj���TڑJ��v:1t�;?q��4���'���қ�j�ywǘ�k�\V�r�'Gc�6�__�2�!-\�(`�Q�4���n�Hlb��ý���W���RX&�0��
�bac�Qv���b��v����������2�A���q0[30�{��79�}�����Ys�ϧDb�P䚹�!0йN�`��^���H#�ɢ�S�}6���B2F%6�kOv���3a�b�q+�R��*���7FC*�P�.|����hݣFI�,X���x�����3�{����w���ߦ��>��'�z�ח[y�r��'S�nm��l�q��;OoXkx�JeAD�A�3%��!���b �Q�`]�l�څ`A�"�i��Y��5ZJ��U8�S�[�����i\vf��&����5�:��+2�e>�Zy4�K��ە�e��S�wnl���g��5u�*�|���'n6�qA6i��1n�s�z�j�uY�;������=���u����g�w�J*I��Ն*`��^��w'�cl�ZV%�U�t�������X8v��aM�P���G�o��iW�kf�e���WOD �ż��*����d�}�/�<�N[̤gQ}xM�jS�Y�N𗧕r7������j����L�7+��x~�qg9NJ���N^��m�{��0M��P^�E����R�]X�Z���6�:zuZv1�lV˺��6{����3)��B*���(,oj�1�N��)K-���.cT���2��+�F
=[]!��Oz�]�X0dp��j����Tm���o)�'���mI�Ǥn�C�s���Sfi�B<�˅m]��{��5���|G6#�&2�뽢;�X]y��CC���P����d�#5̵��*���(�q�]A^hEf�u���Ȥ�)��O�u���Ge��7��3jN�8fM�{�O�9���+.�IVus����(��S��wm�Oh姫�_&�ٺ�t(�Vw��n,��j���������luu��3*�����U) �;�U�lK�aЁҢ�x�e�����>"��9�;i�ՙ��om�n�=�bV��g,[�#�Tky�L�,�X�j�&�52�3��2��$�pn;�ͺbRw���-[�g�,[�B��37���=W���ʋ�����Z�\q[�au��S����8�f[���QY>�_Y(\{:�4o6���M%(�Q񗢎��ǀqv��]�6��kv����[U�ʫH�}�Ʊ	y�����ܢ˔�@�Oj��Z��T@�(Is�x7W9�g�c��٤df!�r����Q�ۻUق݆Ȋ��hG~��<�[H���;��3n�����{_X�*J�@w^�%Q�{��w��S�6%�3
��;��e�;2t�{�r����e�cϽ�N�;�!�=� 2���?�1~��s����|��L�NDY�*�״���뚪�]��y��[#���+����"���N�Q�ٔ��M�kְ�VJ+m�a$��C�҂K�|�'0���w�s���<?d���?0�֩*���Oc�$f�E.*�Oӌ֗���'w�^@9;�����ȳ=-d����k��	$R�l��y���v�A���Mo=X�M�xTB�>_��Xc�n�.?��FU|ROc"F�̺}y��zb��0�ܻ���#&��T�m`�=P "�hg�Ɓ�r>M��I����G�P�_7=[G�퓗�Mx	��Op��V]	�G���R2�Y�wOK�7G�[=w,�;-$m�����oS�4N��o�zS��r����ױ�Gc����?�˧��5G[9��=�z�+��V��s���cR�ܬ-�<F��D����IPXd���������"F���J�S$!��f�k?��7$3�L-]
�k�kc��hhY�k�+7z���VS���uR�9�n {.��¢h���ۙf,�sc��՚-5�d�}�1u���B�]�V�2H��u�8V1l�Ga�c��L:y���F�y�O�0���r^�12*�dP�'�K)�9�HD��۩d$��H�Έ��(Wn߅;��8<w������D��J�>���)���w�oA{����O��$��.8�S1|O���V����y��O\�&M���c/�����w��rM�HYwgډ�,H�O�5�amC�Ď䶬�ʫ]g��3�o���@��¿��� �����]A�����*g�b��L��.KwN��0?�-!�"�b~׏�i��p׏��(���D�q]]��a͇�p,7ǻ� �Y#kϳ�������|����Jj���ۛ�oM0�Z�Ky�^�Xw '�S�x�B��q!Z[����Ad��z/&�����9x�PM���fE�U0�fび^����^�ͯx@\&� �^0ۧ���b�~ڎ���s���by`jy_�TV�<Z�{���撘Qng{=·(j�Z(�zsȓ+d��ޜ�{N0�K2�0��b������MS���Ӵ��	ͥ��C!�;4��5r��c ����)�����U}BX�gwj@����n�-o]�=�g3�a��cά�1;;���K���o@/J7/8�n�1%�껋gp�B�Ä�m���Z��V��O=���.=��f��5�X"�+NJ��_C������@W�����^Y^&��N%H	�L����}�DM'��/N�pV��u�Ԫ����e��/ZX��E0Mۧ\���|���Y����(C���Q��A���:�3����ܦ~�qy@^2������^T1^-w?9��k�(3b����*3����x�3xS�;�U<#`���Hj�[�4-`�����v��A�Z�OЇ�M�|���U��e4��)�y��p�ZW1"=����+��[��U= �#�ۏ���7f��~W�U����}Ѷ��su�.iM�Yo��[�=.�G��w�(c���5�Kx��C����5�B�&�c� ݭk��]�;��7��6i֣7�UR!Tr�,�����-�4<H�bV~�RXM����@��D}��t�c�)L����(���u��f �@�r��?D{ͪ�M�Tb�Fp���&'�|2U�$�%7 ���oF ���peo�Ns���wx�%��� 3
��~��j3�4����[}���y��L`�X�54����&��\� �j��5s�9�����]����\�թ��q8�ٖ�O8��7��f�-�vka˾�\A���O�py���v��T���֩[��K��{v�L�6x_=��(���^�ѕ�#�	y昳��G ��&ȏ��k��x�]��µ�s'+�f�S� ��*sL�����B�yj��Kf�"��^�ÔD'�L��*߬`�UL��L��vq� j�]���a8�,}�%�Ud�B�ײ��-�Ϳ���9�#�q��s�K����V���y@D�[�X���T\<��>^(�'g���f�� S�����p�Q��AV��iMġ���+��t����&f~���SO��*U�&�����>%�c``սB_lM�2=�^�k6���ٸH>�荺�$�A���g����oԺ�u;�gζ�p�byO�!3�Z�,Y��
�`vzg�v<�j,�.qr�>�҂B�s!ږ��z��r���1���k�l�jz�ߠ���+����2^%�"�#�@��ܷ�T�V�^X�֩`˛w	�`��HS�u׭]�5A:�Uyxl���LO�y���<�f7[��&''�6�U̹��#��U�7
�4P3��V�pd�7'oH� �{L��b��ΆNu`!a��<�Ӯ�~�|o�ܽrjf�5�2P)A9�}�t{���f�א�Y�`.��Ô�.�Q9%����Қ����ja�K,�}�X�2�ְL�+�6���m���C.����z־[z��jnN���3���>d{&T�+߉�c�nt
lS�'D�j:��b�wI�5L��=�`)�H�s,��K�t�0�����0�k��vNh�*pUKVm�������=�Y�>�uw�ڱ�����C|���@o{rAW��=�:��DC@/}�MSU�Ҫ6�b�$>�HM���EOM�iC_��)���#�t������C���u#:�W�ۦ{S�#�8�'_�5��a�	��Ŷ/-����g�F�k�������7+��O�GV��oy`F9iw��6�,�A�,���%4�H��WI�극��9&�X�uwMS�g^������ ^��.�m��X}h���ǽ��OS���YTCSf_u��|=˴l��"6"�#xn��)���A�Z����y9�M��{�=8O������]�[(b�,��< z96Ͼ����A�^��f��:���ݻ��QC���!���#��H:߬�(�j[�(��^�h�9��!80��?Eǽ�y�V d[�bf�aS��F���?�~5�8�׉��>ߞL���/��`(���H�a+�}�g��t!�/]�2�kNLU�;�-�������-V	(��h�w!#2�ga��a��n Or!��S�
�5dxr�븓��ް��(����T���	���i��J�f0�Z�����<�GH,N��Y��?�*�S�8������_Y��~��q7S�F�dPyߐd�kvWeE`�"���6��_�O�(���1;a���h�SW<�\GF�/��ke)mY�7]�b-x��Lq�0t��;�Ҟ1~<+��d?g�\|�g�zJ�c�l�O'#K�z�uFܺ`!�b3��k=�}���K��gdg�{�ˊ�x� �7E�D=k�ӄ���ě_�\�W;jmIU�e�mYQNY�����؞"$�˭�����<���ܫ�P=�+VPO�5*q���/K=5�v����C��/y�k+���VK����O���q�㫾�\�G���V]�n���"��5z1�ew�sC9���Խ�N��$<�Lviv���WhN���5�����{
���c��Os�ne���q�@!���,�h���MW����; 3�b�|`�
^*�۰�x��@2�ųw<K$��(`�kʀ�͜�<�9EU1�GX_Vxu޿�^[n[e�2�w�$�].�H"��@�uM;[�2��s��|�_Hܗ9Dj�;�N^.9��ttՕ�r�%d�� 哔��v��yq��ðzݟ1}~�O�6:���Fǩ�a�����61����������G��=�D"�C�>����5B���Ց����"��龗,�.Q����/7���w�s<v�)�9�k���d	��q, ̓Y�"�M����V �LL�Ql�_�v�02�T�>]GQ4'��]3[�#�it?^�<����P�΃�ۧ5G��k�+�%�����aC��x�A~Ș-�m!����
�5����a�������w��-��/t��Y{�.C��t�T"%�)ݘO�ak��PyK9{���H��/}�	~�Y�qο�}��#�Ύ���܃Z�Li��fa�V�8c&�IēC�Fwj�3��R�ɔ:&\Ès�؜�P.�_�RĎ�|���	��/ߕ�D��i�2޽�������H�k��Y�dC�f�q�I����ϵ���������{�~�D܀�} kQ٦�8rj����9��k�F�|�����I"a�Ĥ�f� ���cO�ls�c�]��2L�f!��?fC�+lQ�SB��O�"@���Og�a~�ƴ�J��02��&�.���N{|r����n�/o���f..u�x"�Bd�*V���'I���g���D���T�	۔/l�|Rج����bFr��C9�;5ue�|c�ߪH4�"��vGu������QVG9�+i�J}������܇�԰�FBQ�����ɛm,�enMl:W����:9̮�i��vjeu��-��+���@)ݪ8n~Bȟ���/�hޅ��� ��1�N n6>��	?|�(I��/���s���X��b�OV�&-b�x���.�ݍJ7�1M6J�;Q
܌��T�Ȉ�)����!0�R��y�vDvi����u���T6���|WI�R�65�����Q�l<t7Ժ�~��{*��^�l��ۥ�h'������K�z�#�qVsIH11���$~܅��?}dk����A��Y����_��*��7V0�d=O���U�3�}W���7�r̚��}T=��{P�8�M��0,5�Z��!b̚Ck�:z�U��vL�|��Hh��_=���4�A2}�r��z�9{�Li�"�&����˶��+1�]ܠ��gq��pF+����^��ԫ���v�Hg����3\o_:Nꥶ
fe�R�ȅRsZ�}�絭��������9z�>���Lɛ�S\�L͌ �n���fZ̩X�b�����𠓃I�:X���0���?-	h��X1�GH��];;c�����*�-W�w�UD��(���K(p���;�e�ZP�c������%Ձ��v�L�Eޛ�2ۅ�;c���^�4�52C�O*b`���=^�ԝ�GX��"n4s�]�T�A�x��.�p��*X�R4�@M�r�ts��_�oR?{��o����F�l���Q�M����>��sk�� �&k�m��1�͚ ��÷|-c�g
�[鴃x˖GR~؈�U�m���c�0�7�S[���f�s���8W'���Cd����;+��o��\�XK1��]sw�B�j�=��W��5�Tzx|�R��3]���y��v�D�pv�Gf��� PR��ިt�_��]{�1oozz2��x9w�3��d׻i������hf̓����X܈~���2����lQ3�;zڽ���Q������S��O"�pHF�8��c6�P�iU�f�ߞ��;tB5X=J�n�#R�*6}S�ƌnL�9r�䘄��B}3�cm��	�=滛�ΓguU�N=�85�k���
��������͝{�Tt�Q˳�.�WTQ����q��,j�Ӷ�;�O�v/���.��z6�XG�q����]�����ꚉ�Ic G��\�ʫ��}m�7�:��c��#[���%O^��z*ͩCe�]H�a����-��R&�C$��)�Ya�G��#��U�}pc�0� 7Ik�렶Y�"v�Jz���L�Lq�����i�<H�%��v��i���&�T�9��;o�:��/
�>p�d���s�YT��+�i�]�Y����㪋���FE�y��7�V����y`z?tvY�/�dwۢ����7ql�gv���'Ses�n�e�ءٚE�;���̠ܩ�,�Ԑ`�3�?�Pg;��T��/��þ�*{V�OWX���7Y���?�X�N]L7ƥjZ@�r���z��2nxk����/��y�4zګ)(鵍�ه�e��ű[*�5��/kj���#�;�JŤ5���G��WD�Z+��W���1p�-M��t�u:�y��S��vz�|��ː�#+v�&�ҹґ]6^M��;c9mX%�Z��N[�[�pJ�kD����qū9����n��R�WU���S�lT��[[���"�c@w7��Xl��&�`�q������n:�ƥȢh����X�,�`;|�=Αު]�2:fX9�ծ8#j��]v����۹!e�����S5�����t�8ri�������O�90�Sw�u�D�=�6h����6�
Ve$#��c��m^J��a��/����f��Z4�*�������&$��O��j�mYO�4��9E����yY�|{.Q�e��x�`WE��[9�n\H��o-���]+��nն)����Y��mZH
�kֱ��2�$r��~���7�o���k�]���d���g���0��q՞a���^�~4y���`	%�6��~���p=�����]��}���ru��̜s�[�a�}��G��@o�a���vF�"�+�,KOP<�J����W�'<�Z�Q�рjy�F<�C���G���[�<�@����LQ_]�����T�f�|�{fr�^�y{�J������q��ER�=#:Y��ƴu�|���빅�op1�VQ�⯖[��t�o!�ޡ�I�	�[I'{��r�b��gw#B�n��E`}1)��Ҭ[�?�.�'?H�}#��h<ʐ�e9�غuv����.ޠ�_kt-q�ua��� Ӽb�i|/.�$����j������!-^��feZ�У%�����،�A&�o(�&ej��Ի�lݒ�y�U��Pmo1a�]��bFVo��n��ż��L��]�yc�� Y��Ό�����n�qvǯ����-����͔ٚ�T�:c35��l�_ȍKR�:cew"�C�=f1XpXu$���=V�L]�	���к����E�VZ}M��:v�N~�����ǝ�Y��i���m+�]����+� �id��i���ԙ�n�ɽ��b������_c��G��mE�B�y���:�Tgfՠ�H��僕�K3ZT�o����ݩ	:yH�]�R2�
��O��L �+5�l��Ҝ�Sga�������X�x't΃�����2p��j�z
Gz���*����[�"�:�P����ۘ�E:�s�oH��b����څ���y.V��`��#�{vr4�$jf*�9�m̳�ě2���S�^���T��9����\n^ڭR��odށn�y�M��_��i��n�Q�Nk�Yz��݁K��Rx~����v)��)c�d���!^ZuM����!a<�\�Xc�N7�o�'��v͚��� q|���%�e7)�K
_Gj��@�C7s�����3��WŊ��1�ʼ�x{�����J��*mV��u��W�3|�r	�wU;��t���SP��T���c\8E*ݱM�*E'f�;�A&���ݮ+�V�Uf:T�X�=�w���:���5���u����0+Z�ci��s�*5&"�	�PLO/UR9�h��U�E�yV�%�Ju�Q�jV@��)�:+}]����Q�%)��jG<[c�?�͗=F��Ff�i��A��4����sY �<w�7��;*-����xWq�˲s{8��UU��N�'����Vk�#�	g�b�����y��N�|ox
���¦]Α0+�e~��o�ԥ�w�Nz��rQ۷؇n�����,Е]"��`��+9�5z��8��&dy� �}�o�%��u��[�xM����,�f�_dh������kn�a>����%&�v�n[7V�-��^�h����g�ֱ�i�}��o7��ơN��O�5�*��K�NVF�C!�)5�5�J�\�2Y���;	7v?z��!��2��>�����궮mݎ�â�7l�R�#�f��z������Kr�^)�D9�%Y���x�9�t�����n��W:���,��ӭ�rSo�����9������L�l 酅����@���%��{��ދ�9�C uQ��>� ��~Z�va^}�E���Zـ~������5�d�4Ah�O�1޺�Wr��������.)��<�;
������u�yfɹS�@G՟D5���Qd�9�q�!�T�P=�̇�]��u����!U��?�~����7��:6h ���9��P����:�s������������1�1�p>]��WU�,����X'b��1E���Z���CfC֩��ﾱ�v���'���i�C6(bK��c�W+�y��|K��z;���S)���M��E��R�&�^�=�Lm��OeoU�>y�s�l�mW@ng./��ڂ}p��mWoj/8�fV�&B�+�5���՛3Mާ�J�f�� ^����4��"�׼	�B찲�To�\60�#�xq�-�3�V�J��E�&'%р0@��(M��c�f
�$��}��mݸf����C(�c��۰;�r��m��t�Y⣖�t�}ݔ1��ã�w.��2�E�̄�+�Ը�̀vG�(�oWv�w3�s����4���H�2�3'M+�S��,��Z�2y���a������5�'��t�ڕ\��I)zo����ur��_�����m.�u~���S�á*�p�e�dW�-�q��i���7͐��P���
�����,ه��x�a_���#4�s�{læ��!ZUw��.ܹ*1i�/��X���C4�U���m�LZ)��<��SD��exBn��3�����oZ�h��Ƌ������SA�o�ɻ�xXN=�BT���\��ً�mY�[/-���y���yз��Q3�����	B�c
��s3�Wq	�ߝ?�*�X8[�Q���	�YH���3���R�0�+
��g�ߛ�����a!�$K��L�7`�9�r���P�Qi��n^8����k������R��Qn��b�8'Ld��>�(|�p���=��ɕ��	L��k-����|�_v�>���J���� ��u�{�ީm�Gv9e�us��ӂ��ӵ	O3��
	nN�3���7�����G{�5 V����k�mb�v!�@�rve�n�Ú7�v۹2��ސ\�#���Wb/!�>��.��i7Ox%��@C[߯�rD%�V�Sѝ��Rf~����xN��<T����.L�� ��㿥���u}s]��~�%�{˪�F��@ؗ��S(åѷ�$|=��Y�v�V�]�M�}(��[{^�}���X�8n��Ӻ�0UBX`��Q�K����a�����p9J����/S4�~ozW�����ql�׵�`}ʲ�6*�^B(W�a'���g��ml������ڿo���'�g��c�{qY1
{��J���߆��/�?�]r�4��N|2����-�ߢm�ܛ�[�{����Puw[[�^V��~4pw���`_~���������(I78�'���p[
Ԣ��l?MV[t4s�UY�� 5'����8ó��xOC�UD�q��`�ovEkY-ʞ1��ס��b�/��˞57���>��	zR̙��s\(�=������ґ�e@��S2�L�ՒC"T	Y>u�}�����7�c��o��.ы�o���Q3���Z�E�7xf�GG����b��C�����'hY����t=�����Ya�t]x�{9���ѫ�yq��~����}��h�\Y����_B�N�rT<sS^���i�\��v&�Ω�R���{�kj���snF]��X�,�d|y��[ �zp��5m9��5tu�h�~͆�%�3��4'$G��>�6�/Vn��q���5�sP�V�d��y�ѝ����#=�"�����>?�n~s�$r�ʄ@m؛dS��(��we�g��,�xoB_�ǹ��#���B���=�o���_~5�����,�.�����BM\�W��d����:y�n�U�U7ON׊�sck`I{w����K9��Z�Of0�"�yeS��D��C�q��N��ׅ��,~�ٔ��*P]����؏�]���2����g3���P����Я?hSP�}��Io#��롴;.��A�U�K��0mr��x�1<-(�����1����i&o����{\��^�9ۿS��7;�*�0u돨�}N��ۖ��W>�rwh�}'3�N�5^�J������N��n]�6���˒��+��63�Fkջh�BMU� n=��˕ܳ��e���rJ�ef�+h��~�����v4ښ��c��U;(�8�#�8�񢞘���q�t�d�j���߷���.n�S��:v�f��[�s�u;�e�Q�XI��lE�g�q��o8�iz�4Ҩ�����)�����y�E��'/�b�7�9�
��!Bo���G��KmR�1������63�p]�_�}�O\�Zx�l�έ���(������>H�6 �xn�]���b�p�1� �xz���������f͓&�gAGr��3�\�1��#�ܫ��_⟱�<˝ʗ�D�75q�o��h�\ѧ��S-�|�����(�Z�y\���L9
jv|��W�ݻN4Mtd"��~ۭ���R�w�}�U�}��a�YV��٭8�zR�%n4zU�ó��`�ȥ�`E�׾�[3���}tJr� TC�O:|[ա�+��������:
\o����/�������V;]���X�Ld��mK��'���D�N(���w���m�꿿L�ηE��Q�c2�?�]���S�9Q}�0����IE9�S��BM�S�d�I��7���vC�������vCF�C`����v�o���%�����R��]�ɦBj>[6GP��w�f�K��UMޠ �9H�ʴ�"�@KxZr���&�;;w����8�i�*m���Y"�thw�ޠ�ez��UU�-7��Mz�X���k�_V�S����Q֍��_s�\H��[��J�Z�f���I���8a�}`�o�;�n����*��Lx�!F�Ό������Z���^7kk���ɻ[�˒r�/Gm�����9<��:�D��7 U�cr������nb�A��%g>���Fuϝ��δ��VCٍ{��-XCF�P8�}�>��B#+O�����c�?���vm!�6�ng5!��]l��kl��C1�(Zb�tz�����<#�gU���m����ҫ1,�p�S�/�-�e��Bq	�ٟ=��dւo�Jה�;��е�+1�`�U{��rf��w�pѕ�#�ogU����x0a�b>3j�8ҳ����k��L#ٗP����g;m�!�e���۠���Yu�E�ı�2ι?�m���~�2�ͼպ,����D�X�'�4����b���CKM���y�\�wԶ�XɞU�4��cn�Z5ɋ�l�!4��W����mvnDE]�=#p�̓�@��8yme������S'��z�W��W�����)��;�T��ՁQ��q������p�s��g�.����J�v� 	��/'*�]�B C�Zwn�Ҙ� .����3�6#c�w�ĉ�\��bڼ�r`��۴��N�N���
������2�H�Y}S%�6_��hw*�ĵ�{":�]_s���nw�f�7���8h�nT:5�¨;��	>�K��.��(0��oX�X"G�Ϙ��r�f��0���hO���]�.����]݄Gh�zNmn�+����>�� ��`�bDT`�H�����|A˧I�U��W<�S��D����ʓ �Ҥ�Ĩ�Em�PPR��
9��oi�\m����ow,NQ���q򹻑Yi�v8/I��r��B�Zk�L\��D^�b�vH�C�4w��Ha��{tiVϢ�]��������B�+�#	�բ���>���Z(�K�a�-�^�oHt��7�U���{��*9g�ں�J�j�!���޽ٺ5�ҹ����(Kp
�%!&A� ]�������� {�s��tbv���n8�4����FQ����cB�ܫ�9��'�P��qʿ<�n��-���{V�v��s��`A�b��#-��Yk�!F�!@�]�P=럡�ER�	���ՍhY�h�U ̓�)����\�����˾���c����euh�L?zۮ̞�5�UyYt¸�4=W5��jq�ͨ>�AZ�����+܉C=9 V���5]�Z~B��;���\�U}ttގx�˘��y'�U�D����/;ݼ�=�^הrY1�_�P�n�^����1��.1MR�d�5���ic��+rg,0�L��q6��@�M@���˰�6'}[����Y�-O�MfMoF�P_%�6j�1tՌپږA�AC^�ۂǵ��^Nx�+݂��&���T⮔Ν��^����˗Yw����X�1E� +7�U��2ۓ�-�G{$q�W�'�b�.�l��s�̚,�����gmS��h�\�i�d�w���ͬ^S�L�a{=]�W��5*%���,wB;���qiE��o��P��G�Kގ�m߮~��;�v1�KÓ��屾q��ЭqRܸ�E�i�C��ᷝldo�|Õ�2;oؼwx�w~��v���L��S(Yּ��;�{���$��n�(a�Z�qB��~�e�_P�3'����ci{u>��|u��o��]���R�BRE�X�K�y,�U��W����ٯ1~�ﮪ�[�
�Ӕ��t[�*7ޓ�i�S&����kj_`y�Sm� �ad�X(�S&Q��g��^�?��d��	:'75�s�ֿ�ƐC��7un�T'�F���Zi]:�����+�9E+*�֞�U�1"�a.�j����!e-�_2
��w*�c2IΊ��>�b�k7�݅��fl/;c�T�X�AL�K\�ڼ���R�p���=�+]��!X�˥���n��ZǉBΆ��Z�dαK{UL��Xnu�ְx>��=���������ֵ�k->]�(�U˜`�wf]f�"VWa�.�R�$ﰆ�����#����w�9��Nư�aй��x�=��>��i��|(�yپwW�z�	4���ξ��C:��s7MC\������z�s^<u�s��������f�Hi�q���� C��%@����轢�������j;���v�-x���ƍ	`�I_]m���kwF���뗅���ESڴ�a�����3��a�wNG �u ڗD9�N��c�{�-���j�C�*�܋,��Y�ɗ�LͲ0<w0��Ps�[RO�Ztk#P�0�3\s�*�;����ύ}�����_o��H���a����5̦�L��:�"ϝ��^L��&Цc�;њ�t����H<F�,!B�0�e�Male1��g�� �4��+8�#�d�|��B19�Ɩk0�&w9�w����^a��u�s};�k��d��%�d���@�'X�~�{�M�<n��t����y�x�7cnGö�2��Kh�$"{]�m�v oW%yh2���&���D©g���t���s4�x�{�h6geT�J�t���+�!�%�d+�s��h�ךqv�)���
;nγ��ݱr{z)�\�ed����F�P�ļ�i��L(��T|w��yV+��_�b{;�I#m�G�;�{������D�up���R����nO��:�{ 1�[�os�X+ �纉5�a#c���8T�fB8u'�Wo^[����}fp�LE�ÒuR�;.f�a�ڤ��nTܟP�|n�\�xozk�nr�pȕu�&�h�˜�Z��w8�jN�̓+0��:�n�p"1z�-a7p�7��A,2$d��ǃ���_<�{G;��3��n�:#��}�V�ؙ=d�<ޝ]���ydT�8޴��NLc���Y]����yHe��g&�����om#5s�of���B��:�[�0e�`%Ѽp.��wn�	�KW;�o���3��$��g l����GO]�-�ϳ/{ ���G�r�L���]�ت�S{��v�g9�T+���]��>ʗM�Գt�Q:v�#�:�>�wx2
�U��4�)t���b����|�d�Y�}�C6����*Ù����.��o\W$�\���j��T�U���HU���w1Wf�R�}GyҁJ�dȁ�pOV�I���U�t�C;��4+fa�WnH�hdeWMP�(�|f���[����J��3��n�I�2��j�K%�xN;!w	G�O����B:�ˤ-�Cv3�����J�n�˼&�D�u�����mh�t$􋙻�v�P�t��6��G2�v5޽�޳1]����{��j�liw�\6�Ę�9S�IV�.�Eu���|�&/I��:�j�_u�`�J����;_{˥��(�f��h�OvS��\�q��R��͎����~��Nm�1�*��T���bMw�a��X�ڪ�K7����v��L?�Cz���˔cv=��$�c�kpDT�+����/�q>��ˁ��Ź,����ˣ�K<~����߾�����ͱ����
�����z�l�B*E�t�u�_SZ���<��7�+��<����$�����u*��x�q��.���atr�����>�V1C�_A�鱙'��s}ێ(��r7T�͞Ow����`��\˚�Pt�;�LdC��o���ujX�z��_0�%?z���*��4i�Ǣ��b)v�:�]�Q��+\st�tCUS���)�� ����wxxW[��s NpÒ��4�l��
|Φ�u�Z秲bښ	Ѡ�qy��NVbil�h,[��/�<iSnps������{m���Tv�ͯ߉�?m��k�h�2|H_SIB�B�O{a.��E�^=4��v�3�8pb[9b�����`͝�-�[+�[{��lCJ)�ؔխ
��a�Mq�E����+��ҟ���9��5��GM#m�=�ō�⠅��~l���ǵ[S�v�˻{��Ό\����w�,�btQT����NW�ݎ���t
�V)�往|}��+6D��k ���C����]�hV[ٗ1����!��L��Ǉ�n��o����9@�~��� ����å�3�1�r�%��V(�}���CE=6�6ne�k	Э��XQS(c������ޗ���T�x�Ɣ
��]bi�5z�@�������Y��V��&�� �΁���!�njq1V^�VH�;n�h��S�ީ��DgL�?M�(�;Y�+��-e$��g2S�zfc�Ϟ^5�ŉ	��+sg<l��p�\�̢`d?v��tn�tA��œ^@-X�t�Lԭte�=�x-�Uv7v6��v1����ݰ^�	J�醴WuOo��<��/	N�����3�5}Yi+�[h��W]+j"�d˃2A�}������Μ�19MV"�pe�C0�f��B��,dMܱ��`�]�z+sK��3�F�(�8
��"ձ;8qT7#�8���Nᱴ��솕*4�"����S�m.W�^�a��S}�q6P��v���T�e7+���%Z�$~��.YG-�\�l)t�'<,Q�1�r��ov�]9�
����{x|�9��rDU9�����/�����0+U�����ww9����SO(xEF������oW �FtpY�H�hk�
YQZ�y�km =,=�5F��l����r�:��Ԥ/���7�_�`�ڝb���y�9d�s@���ڗ��e��cn�rj�/�e��^Ҹ	�/Lc���b�Ev������1����I��x_�����e:iį��m����jI�+9x{�~^�c�y�@����å��$vCd̛ݡ���MT�|ܫ���OǤ��~x�7�4l�P�n����s����.ȅ�x�w=��F����NE�u`//�6
y~�x���GY�e-9%ս��/���y���D�i����C.��\�YY���Y�S��߷�_K-"��o3pg���W�h�<�%�yi�Rɢ�ʛ��q�u���:�S� ��%(��	%��y�xye�boCܟm4�*�;'1��A������l�dEbh6Ū�,��j��*P�2����=�����}����^s#��j�F_Ĝ�����ީ�Z�tH�ǓV�e����n�!�-d6�@0�_�����ҡ�2~��K(���%-��=ۛ;"�^MlwGf������>��]��?c�U�ְS���n=��+%+� �|���B�&�1�lx��+!�^����Oq��`���c7�}X��x�aB����$~[�Q�2*&�h��;��[�Rو���f��KrN�:z�Uid���y�Uʩ��|�w�/�Q��cC�θܣN�W��Q���0�4�n�el9�9�Nü)�㸟'u���N�{)��z�<!V����eeFK��>��o��G�?ADSƲ�����vP�~��$ ~�=������3�(��5i����k�#��2L-s*`��I
����ۼ�ط�ƵU� 7BWf2��Y�}V�Ϥb�M�ݍ�y6��% m��8�=Υ�]�M×�iu���ѽ��o^_t�/���,/C~���?\���#[���I�g�|Ӎ�~zEِ��V���т�S��l�]B�yٔ7x_eJ��8���q�T��q߶-�Bb��~��m�G�t~�1����x<C��1"�tn�X~u�Fí�B�v�C�h��Y3Ъt�f�!1�{_K�8�egmj6�nd���v����*��͞�4�c\U:��K  ;u�7��ܹ�E�M��a��������5�E���Tݦǽ���ɈJc�9�(X�������97������ť��������һy�'21���<��Ī�r �ߧ����!�#�*{~Mz؜z:�WY["�����8��%�`�!D�;�klcU�����qA�O�p��u�0�v��(ɡY�O��ѹh�7+B�&y�=²�)�_MͶu���MޝYc~+�cA�1�2�Y��唾@$Њ�tyB�'H$1隅��ns}5�뵜,kKκ#@����n��:�ƞ�S��!������5+�՜����0Բ���M<�YE�9s��k��G�#��7ui���G�|��� �����M���8�\վ��Yj9�s���+���~��� ����P2�'�RKjy��iTzq������u��`��7V�� :*K` �~�������k��Q�$;��ݙ��t'm��Ì\D�TL&{;�#��_אor���R��?�l�hl[�,�9���#B3�	�z��[[+]�+9>g����߫���0� ����n>j��y�?d�}N��;�4��rWS���ox���r��R����tha:T����K+vƝءճri�/��G9T���N�c�X�3q��*��V�f������k��e50�����:���`���C��e�Z�)0�4NU1X��B���\���^�2�Jֱ������*sm)��O-3��3y��KmFs���m�~���x�ܽ��A��uIJ��z�������ɑQ"������T���Q���w|�}�������o��nT�����t���@*�%�����q�/����RWƱ��Bm�j"��^�ז���&v�2��Α�9�4���\�K$/	�p a�o�(?�8#|{v��ۦ���]�N<�xy��l�M�cll��eJ�B��=O�������An:�w�?��J�_3�e���������n��u](�E@Z:YG���_[���w��4�}�h.��S��l�q=�y�Zp���v��t�D>WC&w��:rr�1fW׭w9��D����-�u���Р�������bO4Fk@&��-�"�������V#�4E�)j�1hK���{��3����뤚��Y��ڻ�ߐ60+�}��f�ɯ}�+J�q])]�����2V�/i~����ߏԹ8ؕ�|�˷�8;���fk��X[d�n똫9�s�Йt2Bq"s�#�m�U��6�7��h�`�+*���L'�b�<;�6������~�������"�N2�B��@�E(̔�뇶�I���ϸ��be�!G�2�[X@�(�/����3�^�ͺ�W��ʱ�j�����x�vEzU�w��e��-I.�+kq|�h��l	��*��bW]�̜nd���
���8c[��!���z"Ve�%�W�W�r��V�0P�C�}y	��D��>=�_{C�~�ɨ����*��S/��Dlٜ#�����%׮9+g� "���|1�gi���]�����n��y�}��Sz͒��.u���q�Oi�ɷi��g��ٯL�0u?W���}�_;���W���'���Gǎ�E^n�[����?�N�B6���^�ʩ?F�1	!�d��6[��湯��W���3J��g�u�U�+����Sӻ�X�n �5?
�H��=���U��j������䫦��3s
�ͻa����yTq��O����Fm7�J���h�3���p��nHY��a7��K^mA6H�dqr����+�*�W�����7�8�#RU�U�C����]N��k}�K8���^�wc�1���aO,���z6;w�Y�юk�T�:w���L=$RkZ�pK�h˒�+bi����i�\�;�>90�v�9�U�*��VT.���Y�g�ׄ��Gw"*`��$�鵒𝴟<�M۲����)��l��6�_X�f���e���;3z֖��C,��u	֕��X�8(����G���3|����ׇ��q��� ��|x�Q�:���Y�w��\�}t�ч��N��Y�BR�K��ǽ��}�p�F�+lD�էb3|��Ɏd��
�M��NJع�tv)������c��L���J�f��鮪�o �ܹ�w��w ���mƶk2F��{�w��� ��TU\����X���ֿ�sX��6�v��p,���aV��UD.\�}�
�����Q��`�{�;�!�)���5p�#���;�¡�x.-{{i��1�azf~�Ay]_��d�>jL߇�c6�p
Ծ�vN�ʔzW>�^	ӕz_���HU��`����z5L���Y�ʅ͖��ۻ�}���u"��WL�d9��|��L��pv�����f`���q�1���TE�Һ\�]\�t�-&9��v��D�;�Fx�"E$�iU�v���*i{����FFu��j5����t��1�^�vɓ�Ti7ke�PJЎd�v�cÙ��v5����P�ۗ�u}/���:��
&�J�Y���sl�yݮ�&|���7W���ʐ���R�ŉd�N\�z�%��滜��-p'�ݨ�_�=�=o�g]޲�xי��W	+�'l��s��Y���T�����]��݄�ţ��/�oE:�o�Y'n���_�g�'�r`1�����ɑU;u}p>���6*:mY���zN��hk�F��]�^)):�[�8����P v���b��U{�_�vn��S����gkUI��6�V�~�z�ŗ5����.�O��&M�޹�Ʋ�~���qb��R���K��2*G9�(�ͫm8�2��<��1Nu�e��+<�i0U��؆�:�E�[g�{��z!�qc��O:Uێ�.�
t�#�����*.�VVK�Np9<�ݴH��{ٹR�V����7%���g������0�։�+&�g|�?6^t�2�E:�2�u���gB�J�9W�rpbE�E���[���@T�r�xo�:4K���e���l�۶i�DK�����fe�"��\���Io\�:^�k��V���D�����ɨ3:���j�CmU}����Ym���}rm����9�w�6��=a�P��Q�[��|�ث������ӄ��i�v��6孬Y9,��W�e�{��e&��㸲��<�C�V�P3�o���6�o{��m��yv�ؤ�ں��;��R�@}�0��P��m;�h@��X@�8�P�� `d���q-q�9��m�Mi�!휊}S���;*C��� .�݄t;�(�9d����J��r�����M@�x2}���N ����y�9;E7�d�ޱM�:|;��w|�K�gt�cYm��
֝�Ø(o>�!�G� � �
w34'r�;�xo\���S�l�!�Z�
�&ӝ�b^7!�k+4¬jB�ԥ��whk2�l�#M�#
@�&
~i
H��� ��m�P��@�
"P¸'8�H������@���>���(��}ʶ�����_��́��Bp�8hgw��W���[A#���l8�0Q�Y-��+�BD^^�*`�Xe"nE���`9���٬{)q�SFp�ct��dX��A��|��uR��Xb�YYjҩ�	���8fde�B��Rp`%�e�wt
��fp��C��'L�O��j��1e��jj�9٣�1m�a �_1�f����Y���9$��$����K��v�{�r��Ox�ކ�b�T�I�3���2��Hr'�J�{qr�G���c�Zq}]*�	^����z��лֹ<8��Ή\v��a��0#�V�;,g*��ې,$�z]`�	��ۆ<�XB�5+��
ʑwO �F�1�q�C�<�.V�qB.��l\{��w��fK%�؀˵q�j'"��]ue�H�D�{����F�7��U�Π�#����on��×Pu�����7��Wm�*��j�if��>͜���)�ӗ��j�]V���E��K����b�xZ2ޡKZ�^�\��R�Gtdѹ�������W���U�΋��x��\j
[D��ͧ�S(���/bZ������	��\_�62��G�J��{a�]Nj'J�~pkq^H�R��J�l���Mos�9��ᓎ�˴N,�$6�Ene���`�s��wW�J��N�w�2>
��խ4�:̏30��J](����w��^�g�{�h&͎�e�'�הz�.��v�� �ܮ*���gr�iL��	�xl}�};:����'N�9�7]�7����l�}���*��Xpc�P���`���:�1���a�4��d8e�lM�٢���������Iۏ-����Ѩ�DU�f�3n\�@���e��4RZk1k� Ń�ww蚋j��{n� �"�K�ˊ�(���o���Q�s�Υ�����`��T���t?=���5�J|�mmu�
��r$��uϲS��u�vU媮�cx�p�I��N�}���͸��$�I���<�^	�寧V�Z�#�M�іxf��D�w�pV胯�k2�snb��Fڍ��P��=�H
[�i�2��7[w�}l%�қ�0.S�� �}��U�ۂL�dχy��0��)����/`�^��@����L��l��_����O��>�e���}�C��ۜ������L���V���hk�<W�Pj�{m
�VJ�!�[��-�C{._!\⥞��x�U���,���˹����?�Ƨ0EF�aoy�:�u9���4�m���l����$ڽXn�9v���pQ�pJk�&>�^i2�U��u����ځkv{z���<s{͏:�+��d��ʽ�z�1����NH�ֳL,����u�0�NL��������U{�s�Q�����ͮ$�߀��-o��n�7���'Z��*�����fK�o]}��.��ئcd�����K%��$p71��1���/-eY��׫��7���g�G.��%�ç.J$�-=}ڵr�\76�S�̧�vt����F��)t���3���5�u�'�~�u�I�[�^_��`쯣ﾇf�0�!�:C����[RaE���5P�&A9�UUgb��	ԟ�``gg\�p3j�+��};����L�Ta͖��wUBl�y���E��\LC1!�@����>Ӻ��3�����{-����J;�eHI�����ZѶ�Z��ޒox��^U0�݀���>NcsQJ�}���mc̈́��1�55nnSI�Kuh��X�;�g����#F�;K�[���olEB7S#��@�1��,e����ܺ��Q�UBc�np1
E�ƈ��zx��s�\���,�t]`�������j��G�Q��{���Ͱ���O�k<�=M���=Wx�lF\oZ��秆��2�ǫ������i�Z��ϫ/����[h�O��܄���f),d��}�y�ީ�@d������+[E�V1�=��Y�'�=ܔAC����vی����u��FN@���n����$E�S��ucYRM{A��uW`H��c�;��js�
�Sw+�`1R�`��]�7�ξ�6�vm_VfӅ7��'0��z�5jzWf-�y���Զ�)�|�R�}w���`/�>ùKح�x�loi3[٭-5�J���ל3̱�3K���v��O��v�]�93�t#�i��n���q@ޚ�OaK±�[E���x4:˶SM1���	T�/��8���f���!w�¦7/f�ק�h��������Wl+���-��~����y�$�������tOW����}�q�q��o���,c�by�C�a�JׄVwt6�q_��  �Q}�w��DYVh���p�"�=��8`����=-�}��x���t�����2�Ӫ�� ͛���~t7G@⇧�mu���S4���[S��qȫ����A��:9���Dh3�ln� �Rfe{�囱z����k�b��5�Wbl�G��S^���PȀ#7��}ۤ��e�7s���r��p>}���E�E�v�3vbߴX��5�S�܃&�zCMS�Uy$.����8S�%��oT诸�/�Xr�"���b�Ѳp�����8��Ḟ3e�miW,��B� NԴdsX|O�*B>��{Q��^k�����S��-��+^���:2�ܭXM���ѓ�j��6�m�Ƹ��z�3�̫��2���&0xm���j���(���ҿh-�?��밻�[�#�����0v����C���9=!
`��4�[�0o �a�d+�2���]��5D���QaT*-H�����k��J;~�U��w�/M�F̴R�:G���K����ܣ3J�n�����j�]�^>�D�WZ}��X�b t����7dA��%�o*'�w�cF�F�����)Q��tms�kԪ�0#�N�&�DzU/���/4n|/K��I��t���MT�
��#6&fm��&�@���}�K�!���.���puj�(����q�2����v�.9��/�a|�2Uu�����2�2]�QьiV�}����8�W��6p)\��vu-4�\(l߃Ef''�~�ݖ���Ǻ�S�GJ=͜x��Y-<��c�p
.w����+mV7#��+��gqOgOԵ�^��z4��(��۱�oz?�����=a�2���k�dwQ{��e۬bdI�ҧ�k��+A���e?f��sVo|��D��>���9�o㦚1�N���>޾��tyoѰXw�y�8jW(D�w��a[�M��͓�����Em��5LF�p��4���_��Gm꡸KF��'__�C�ߨ^�b��H�>_��]�[5䌇3��3�N�eg"�E?d�c���5@ R#���鍷l��Twp�����l�v02���l)����AS����-�i��f�8��A�!����ٱ��7�&���~+������M��-���V�7��ˣ7h;��u�#тc��V�c�ߝ��W�Z��j��,�)̍Xk���+����3O�w�z���[�;7'N�� -�,-����jر
�Q�@�>�YZ���u���c��}�զ.h�{e�R�n�U��2)��v'e,��u����T����ٽ�CY)�0�b���D�����*hb����n���y�u�ﳉ5�#���,jn���]�yf�rw�(%��ܹ��I�d�W~n���?^�;�ll�م��^��5�1����;�ɉ֊�'woqF�q�Tƽ�bWv���`�rG��F��"b+$��;�]�Q�/k�q
Xvz��^�͘�j�w���7J���t��՛��{%L �{�(1v�8��y<���}��븕~�~�X�^�����Ich����Uzc�[���~�刯$|D�2��ݛk8dJ̎���Vsk�/�	���=(��DM0 ~�s_]�������D������/��܊Pf�@8Z,Ì��;V�UT�NŹraދ�ő�]�H5t�`T4�D�cn�
o�zG���*�ʿ��\�<��x�*�R���~y�Qv&Y6ْ}�ҙ�7+u��r���Uͨ�_���|f]UI�!�:�
[�˯�2і��(*�E�@�]���x/t�,�3�n�͐-�]�Q�'Cݗ����r���A��F}���͖��\���C�c�z��ԫ�u�g����5T��]<O;� �v-�����|rX�U��^B�f�>��/��� ��W���|6��!�3]eyV�_&���ׅ���E�^��똜:<h�V��Y/ug�g�K���h�!ݺB>{�����<�$Gq�J��&VB�z�U�߼��;�q���Ǭ����]�+F���k��)���M(�RH���z�S-�Øy����U���������[���6~�#{��[�{�|����Au"$�X�� �~,���3�u����[����sIk���>�?���2b6��tE���K׌Y�Q���=k��B���RQy�0��U�S�]�t�i�¤3U��v�Qy��ӊ�-b���8��s�eƖ�C���T��ć���X�ܝ���~��.�q�CV|N~mV�}p����ݚ�[����T���񭘱���L�p���l����Д�#*j�j5e	���K�`���(!RKjҖGX�s��oo3]��[��z��t�f�"�!m^6xS�
�c������R"v��{^pSN���Z��Y܇}pr��]y��㥇�>����ks����3���e�wwsC�R��	Wz��Y[��f�������Lm,��th��dmH�4�#*�p�1�����0w9[)��?����ߧ��[ޜ�T�zl��,en��{wGS�GO\$՗�����1�ʇ�`�뙘}����ԋ�h���fxU=��t�Q��U�U�U.�WS3�じ�|�UQ�eBe���^��E�%���5�3�@Gø\P��AM�4��^|U�W��Ƌa��3�3r���ѹ!�������~��{�y�|���zq Se�S��ט.�aa���=��VĂ[�qٻ�`��8�zW���6��i*�hʌ����lhS��C$nc��`M����o��8;3��CF����\'��"��hjzoP}Ir
�Ud�ժ�wMdp�v���q�g�F�CA�!��j9�v��\校wL	�z��H������n�3��[�i��H����te���I$U���r���ݽ��L�j�$�M��ku��s�e�U���R�s��&a��:���9�Ǫ:�j�����)�d<{�&�\u��������S[zx��.��@�B8�g -cYk�{��a��\�D�5NmF��
�=Su ������<��$o���:��5�#���}>�φ8��㙨^���e��Ԏ�>����I�_h�N�v[5؅p��i[���v3fưX�4�7E,�0ӲVڑ��ugD����x�� ��p� &1~{~̶c���*=^˯"� �0��u�gL���_P��9�ܠ/ȧ��^-���.�vX^�ܨ�6���������ﮦ��D:h��߁��3:�h���wg<��I�Sӡ�W�q�L��5�J&����/��>
,g`�;�}Z��[�[��l����� �I��|�ݭ���¿�z=1�Ut�f,�K�N�R������P���ч�ߣ��+�鶣6�~5����7���B]���yJ�Wp�Vr�v
��j.1���K����禼)��.��w��D�ҡ[��np��bd`���OD'p�̼v{މtfX��5���^��ǲ]�[�1�(��0�Ʈ����#	V-�؄�W�Zn4�o��|���%N,Ź�f+�\{�D���C��V�ݰd!���P9��Ty�vY�)����^��a;zB���$$�����g���������͢���2��;��η��Ż�'�c����4�O3|lԝ�ܓ=�"¢�n�����xy���ۯ0}Ւ���I�_U��v-���lF۩.�<E���ҫ�~�����{�����:���+Z��[���v~p��b���Y�.�ě�ߑoů�P�{���]�P�Z��q���Z����k��~� ��+���o��wO�ƿ����P�ù^�N��TL�Ƶۭ���s+�g�"G�ۊ�Ӥ�K��k�����G�嶲��~�޾�+��PQr��{�ۯ����#mکysF�U���t:���y�r-��z��/#d�Mh��p,+��2��Z�{�1���Å�#�DCnء�Z?�����l�8�wG��Mr�I9c�s���c�Nq�ݫ]�6�j�m�L1Sw��2���M��5�ޭ��1ʨ�3G]�yWɑ��9���� ���ne��SQU�΢*�i7!�@�W}���R�)�7u}�]�ݳ�no4k� ��� 8�Nm7,�87�I{E��Xb��n��-.�v�����q⒨iq\C{�e<o�2��_,#3�yQ�iʬH���ʐ��h���;�� �p�hMm��᝭V	�q��;�� Cl	ۏ/5��}>�+�k��=��w��V��p��uOV��;^=�81��k�٣��5��[�f��ty��qX*��m.�6���	������vq
蟛T!:*Ba!:��q ��!��k�q�֒h�̌���Lh�mh�k�U��(�v�լ���pW�Ս
�Qp��8�y0���=y�gY%?�\�]��{(��0��ڤh��`Ƙ-����aZYZ�P���]YѦ��0�q>pw��7�t�n��W��7�2.{���}�����.��G4O��i�A-6?[��s�l���%Q�ڳ�R��� �;�.7�����x��l#�ѷU�i��G����S�X:�
R�e�Q����'1w:S{��ZT��6��xM�yʖ����M�X�S�5>�˹PN��_9�Vd`L0+keM�rb�=�tY�d�RY���7&�˧Y·��n��s���ob�v.� \�GGO("�M��BZ��轡9��y�Fn���ʊ�i����D�nU�pM�'t��m�ےee���2�L�Hp&�Y'�����9-���s�]�Gr��
����/B�mN�/�6��#Ne��Uʚ�^�F��S*1��1����d����O�>FU��b�,^�u�ɞA�5}Ƕ�6�n�!��y�H5�h#��M�ޝu���X��H��'�C�q�'�KU�Y�FZ��׍R�R6�&�ə�/s���k�F�E1�5Z�u�{����X\|�p�_F�k���"�hW�QMڅ�}O��@����	a2WZ�n�{�f�D�A��M���d:0a�\+��fSiR6v�V�?�>u�@��ŋ�]y�Z�N\ ך9N�HrպB�G
���}��9T.j{�s�'�ݕ��R�NPEո�։ǙOa�N�]�҃��J].�����;�7a�A��'p�G�y�����T�5�)M�Cu�wb�� ����|���C�\1i7o&ʂmd0*l�4�͹uj�d�\Ar[@^q�Owj��tcm�HY����W�_LUg�N��Y[������J�w��Zf�N�M��%��hu�d��v��nAy\E� ��:���}���)��k�S-2e=4D�M�;MZ����A6�=ȍ�98EƦ����2��Eg2���鳧rr�숧k�y6q���F�P�i!.Vs#Tw��ۮ
�6۵��<<s��u�i�f-Od��±�w�u�Þ�Ξ�|���! �ާ>���J�}3AV5��VM�r�"lշ�2�2�o�C egi�S؜!C���ؕ���b�h���yk�)Z;��Gv+���u����~6q���J����~,R��`�[��;[!�����y���o F�q���$�(6i;�G;�����[7�5h��	$ܑ��!o��oRyHo����In�\�q3F���Z�1��0�6B6!��U9[�-��9LL���OGCB�<�V�p]ٻ,� w4];݋���G�5�x

��>Ms*Z����z�1b�\���Тƫ�s��s�\�՗�s׳]��w#I;C ��}��O(�(vr�l�Yͪ[�rj/ې��{o�D��c�L,mF�^�'��x��Tӽݕ|�:9\����z���[�گv����M��N���MCg��v؄���ab�_���k�[疫��7-T~�܇�g�>�\K#?8����F�=�h�IH��}��ﾻ���}^�xS�vޙt�gur���oF��a����0A���L]�����N�}38]j��!��úK�ɱ��wPY8X�Tn��Lc*^\�����w�} �	 ���,�����ub��w\�vt���N����1O@F�lѹĄo/��DwŝI�È��:9=�-ӽ�9�6ΝO{����J�kQl�vX9r�*8��D�62ᡏ^�IU����K�Le���6iǞ`ߖr�$�~�.{�[��K�B��2��Ȝ��fݴ�=���׸@�~1X/o�͝WQ1U��IL;�P���k�%X?��a�v��^���?}7'v*;U5�6�x;]�<X����Q��ڭ.M�#U�֠���� ?8�G�L�����gS;E�=F��J�s#=E������� ��Cl�A�=a�ܨQ������@���F�z�nn��m��i�b�ɮ��y�v�`W$-w::t�  *����}'�ŗ�:�<���sρ^�;�$,n�l��9ԶCq��}x.�M�����)���I�P�+����5+0�
��AaX G�O����jK���m�C��vnb6j��|�b��E,We���,����WS���NdC�F2�6Y�1��\����n�2�#Sw'l����jS�;���ݵc{��1Q��;C>��ҽwOܐ�+b���n.�~H�Q������B�X�x�+X.hs�s6?mnun��c%_�yulok�TL������@�٥�+;#��\�L������9$����������hrBE��ΊX��f�s��I�S�Ԩ��L��Pz98�/���ߖ��Ϡ�[��d�.#�������]�W�#m~��8��}V>����U&F50�%M�G�g랝�M�v��]����0YVP�c�n��[�12:��N��wE'"��d��+�YB{Y��޴߻��w�R9l�sO4�>�ɚ����vQ]X�^�S��^
w�+/(C�1�ߕb<��?G�{}�ꬺ�AY�=d���#����� � �v�{i*%�Ȼ߆]�l�鿆���!mꬆV_
�5�AbaAN�8��U���%�CdG4���S�}h.��]26��J1���SJ��{����r��y]��~�W2�u�y�u^ԝ�I��k]��L��Do*���Mcg]k�[���'��Wi���GU���#$ffh&l�LH�R�9�K��8{C�W�`��T��5��T��K-�.�bZ#HL`�T��Ū3�vRzݸ���{$~���La�2yF����~v���{ݑ�9���0�e�+���Gq�MOS:�o0�E�	�ֻ{��R�p�՛Ѵb�q6����-��2���j��>��_�	�w�:��\���_E��f���AtFe�¡ؐ���D*��1٦��|����԰ pun��Eܝ��O"!�${E�{�%ʔxay�X�=����y�N�㬗�u��r�?�?k�Ԗ+��~��|��1�bݔFP�������]�@��;�."�mzf"�"b�7�������ax&��t_��9æ�9����'�B�5��#�O����9g�}9&�l���7�k�b���MŰz���=�.
�U��~�s���W�����.��;�Q��:�d�nt��7-H%��1�8�@�9�]^w��������*����W/*=v%�j�ÖJ�+5����uwF�Ж����˩*���˜�qb���y�ݘ �VG`2�v0�(�_o`3t+�1f����r"w��4���K©0��E�7��@��.�}����R̬[Npg+FqP�Tӡ�fܘ�Q^�=Wy����ᲥS]��)�Ҥ�O^?���}�u<�z��
~;�*�ܾ��9���SY('�����f�\��^�k��>G8m:󑞄�����O�QfOu��h��E񚏖�V���ƫǫ�y��:m`z����/����D�4�V�u����߯��:���H0aI����ߔ����&޾�dE�\�\w�)N�P�.�j@k�F{6�ը�;K�\�pjK��D�v־|µ�N8�[�ż1��ȾT�n�I �ȓ�����^��_D�+6w ]!I��zlм��~��51;yE�U�^Ke��4C_/��;�.��^c�{��b��o�VN6NGBZ]��])|��mu�� 5r /5je�ZB���kwi�����7E�ww�+{g0^ٛ�)$B������uK�X����8���\�GXr3o��ԕ�@�7��q:��z�1�;mvodE�3B�n�Lev`��`�M��r�4�ՄV�Ё��ntc�:O��^Q�����UE�9���5��~����8\*�+n'O^�����2Mt���欎�G`�%ӆW�S���OΝ����]
}��)���P(���#'mv�G�3�����G�7A>Q��:��OxW���R�*YWu:��bmH��6�
yX�8��x������I����B�f��wuK&c�C󌌓xi��X�	�
�M�	nU6W�i��k�K:K��/�M�h�,���>�C:��Cq�%��9���[��Y�f.�f�����j���5�V,�y��+�U_�{_N;�w#ʹmȊ|`�����}����o����=8�݉��V�����ep�Z|\��G�O�r-�P|�i�~7����������z�:���7(]�k�J�$��4�D��1Ͻ�׿k������o{��/��T�7[72��L�.��Z�)��v���9��1�1/��C�+�Z5X�G�C��û��P�|�-��t���A�{�S�_fFsb*��� ���*� ל;�\+�ؓ�*����w�D��B%�^oƵ�v�툌����Y5��s��t�+y������=CGڬ0.�n���*�c�ڨ�"��x�=>q�&E���X9Ӷ�.��C͌������U؃M���`7���މV�<�2���Ol]�-տ<�y@��.�%��r�*^�_��2|vz��=u�N�.��S�cDV�h8�T2������,P7k��E�(�r���� ��w����e��ޡ�*>G�B+<��˗�^>�?gx�~x�.N�j.̦u4�r�{M;�X&|.^��u~�]��֜��`����{۶lU�%���c=u��OΗ�M�9M��t�I��v׫Kt�I�8m
�Б����D���k��o�{���Iʼ��f�浏��[~x�M��L��~�]��b��u�����
¬�J�i\k�5�Ѹ? _�I�
.��DCZ�`�U@X
,`�F|�7ƚ����}���9~�[���
�S��T� �]:��rg��Pa�&^T�4���sn�˹�ّsc�8M�>;k[|�gv���pw_q�y;5��忼&��wv�<y���y�~C�~��@ت���w:��6I�Щc�����!v�-���ާ��:+<��K�W�<�{�sA��3�wbS�,�o=�]�K���iܗ��zꍲ�?	��q����vI��>��u���|o�w�_��r�-��\�^i�}�n��vU�m��dk":��#n�6���F�$;#)7�Y�br�y�Z��s*�ō��=�]t��d��n��9��������o�CYt���~�L~(k��{7��'u�,��%�VFT�V��N����&�8�ݞ˫�T�{��U�L�+��H�N�»�ꕆ�^[�����b�������ަ�	�qS��N;�׭���g�F{�o��Y�յ�1�O,*����i͏a�o+7�W�0���d��_�&��������n�}�q�/n��G4�Er3Ky߾�]�φ�2&em�I*t��w�%c;�,�khhe�7�Sr>�F*�lg*�U�]ګb[�e���S:��N����'|.��(.-����w�ਚr�t���l�E�eCiIj�����sX�.��Gp�C[G�2�!�n�ke͌�R�:�-u�:��F!?%���=���g�~|}��z)��}�peK�`p}�r3=�05�0U��}Э�t�:�@��Tȡ�U%N�Z�5�(|��v[��u/FN�2���H������v���m.�F�T	k��cj�F�
�y"��y����4_4�q*�w�������]hU�����ݣ���Cw��9;��@�"o��3�*����T���{;&���y��Z����5�����N���)+���F���wYo��%;(+WLE!�&k��ֲ1�[Y_.�aW\ F�7`ߠv}�C��E&�R�bL'[������ʉy����'��c��;����.{;����g*����/%�r�f�;����p��}��y��~�o7��{�ɾ��\�����U ���]�������AT��i�1g����g�=O9��v���q[�;��3��I��1�9�5�`�� �rj`�7/��v��Fs�9%��h�S�y�!�lU�x+(Fxp���V^������lBp~�0ڙ�}}�O�b1�wTe�u>�4o�\�ҷ��~��#���//+��W6C������Q�>�)�C��ivٶ�E6�gw�K��<&�kP�^s�(��ۦN���+�6��p��p�1��vsM+��p� #ٞ�^��ʌ�Ѓ��ވ}�k�:������K�'B�lɽݝ�{.�x�2��lZh�v*y�m��O��ױ9Z�M��H���m+?l�͈����o�`�grg�K��?���\��߿og��T��ib�F�dz�Z�Z��B}~s̛̬r�Q���xF�l>�y�]����Ox� S��9q#���������T>��^&��'I��� >����s��{�dj�˹��o��S���uGx�ul��|
Y�Cꩺ,�Y�My)�F��\S��ܪ9}�d+'t=�ڒ�dV�:x֥�i�J�Ԟc6n��U(Dĝr���D��gmvs&f^.�i֮"��[�dc{��y�ic�����������A����g�4v�*���&��B���k������ڴp��#/2��nY��݁V��*�s]�Au�Ku�܍2�}�k�.ڌ��;cS�kܮ��a��X�m����jB��G��F�c"��m|r�����g�VT����Ldn8�yy������Y��S�'za5�w~�6��s���_fL:�z�Hj�DH�b/�@�z�H�
t�'cci���
)B=x�]��H����ባsE�a�����!Y�b_3S�X&�vr�qR�X�}���b�{G��k�q�*3�=�-�W�:�)c5���4�k �wr�}�aj]�Tm�n潭M���x~��i�Sۅ�Uփ�|�@ai3Cā
1@���\ҍ5B���8���Gob J ��v��b�=�.`�w�
��j��|�<�������u�gE��a���QC��5�}�mxzeGQ���b��k��I1sT�x.���#c˲^�\Y��)�hՁ*d�����w��#�l��Nr�wЭ�1�ӛ����58sw�|2]N�r�/���_Q��,E�Wғ���Fӽ�;1b�A�S��Y��"/*��f��F�����I��b{��JT[�����%��Y�@O��y�3)��O0�ܼ�r=7���1B*o/�����e���G�U�6�ݑ���M�ۜ��9}��_r��}���X�Hs�mAל�-+��Vۡ0֕fb�a��*��wc
b3u��N_*��A�@�ӇTeX�Bf
���Wo׮�	$Lm�yd;R��z�hz����O{�K[����êT�n\;�jG"�fڬ�v��򶸊h�S�WMy�GLqf˾����f����L��\ͻ�V���@�Y����d$�]B� v��6l�nW
��D^th�I�IB��|� bz1�%M��(ޓ8���]%G���ӻ�̹Z���g
T�n[����ˏa�k��/o,�>t�D�w��k����ʉ�:wE(w�	*FF*xwyP�y����/l�S6;}���i��h�y�rca�]�Z&����#R:F��tD�+X��Q�'y�Ny��f�%�im�nT���ֻ�i�uҔ��+q��kw�%��K�u�vv wb1v��$��)��ne�jl�Zkh�u|�M�:V� �e]J��i¬�Ћ,rW�����o;���s{Uڀv�z��if%�_5s18º�����R�t�W[amv9i:֍���YF�]��$�efG��Ѹ+#t��8�;+v�>]�y�q���TL���c�\٣��w����'N"=���'�|  &Թ袘+z?R�73�]��d�.�J�e65���MgC>5N(8��G8uL!����Z�g>n�F?��B�f��3��wr��ed��A�y��Q.�֔�k)�3�KH�Dv4�=�L^vr��C<h�����ȷ6���D��A��������j�"���G�eۙ��̜�j��L�B
$T�E�HB�봀xs��*�O�����ou:�/�q%�t:�S���I���R8�:GD���wnfT��wiL��a�;�x����x��n��xf~��Hkց0�y݊�ʭ����Y	��ܷZǆ:�'L�$O���>�=>�$Z�v�r�M���}�?;kǅ�6�d��{i��lM'ѮF����n�.�L�=n�&�_xz��E?���W�E`J�����[��4>�}�lOuSP��Q�h��o�8�}�� 5���#������BJ���ӚJ�;"�[��g��C�Ma|�c�p�׹��g3޿�r.��0�ӉyC���1[���/ �(�S����Υ��n�3�r  �2�]�WU���f���,QT�պ���Q\��1E��X#l
*����w�k(��4�C��v;]*�vw��)�N�͏_7��
/Q��;�n�d�r��w�#��Q�j��v;��:)�j�\q��NY�d*t�.��ԻgQ��]�^��}��.�2�iE�O�1���AJ�/7+v����<i����0ԙ���o�׎cF�ޒWr5?j��uN��܄e��S��]=�C�7T���\*٦��Z��t��a������?ˍ�C�].=C�G]t���mz�<16Xʰ�VO���f�~��a�����ڰ�cĔb��A�A��U��mk�`E���f��}G��S��&q*j�L�3�e�(x�qLk�צ�R�����g���6z��z>�%��&�b���
l(B�T�����	ɴ�Y��/�d�`V�\w�Z���w�Be4�hlBh'[�Z��v�'���ঈ�5&p{���֮�y�xЦ��ݗ�G��Xr��%Y�:�� ^�Aܳ��v�ĺ�9̤�J���d�U=.�*�	\8P�{�I���C�X+˖=��	7hWT�����鞟����^wa�;�$l��@˧��3�Ԓ��s��ȑ���'3�����{�>�uό�8�e鹆dbB�l�f�~gX���<f�ٙ��O5l�E__<蝪ݻ��:�2"�:j�k�&�j�ǂp�}4e�){�;��J�HP���!�C��x��I�Mwe�9��e]Q;��~X��j�P�d``!�4�5��nWS<�l�qSɇ�ԟ���@���q��
�v��[��k��^�N*�u޿�{�� =�QV����?��ekǠ���= /fX�i0]�N᱌C,t��qb[1O*I�sT�"I�V�\���	�,�.�� Є5�8w˙Y�����
|�V�U�#R�v���@}�/4z���k9�=Jϧ��M�n���7�-���[�j��<'i�F���꘣�=R�Mq37(G&z3'8BS,$]�dS6ֆ��_���}�;=��@���6�yS7��XN?H]k����<����'ܝZx�{dl�p>�5.��7m/:5HrLC�y�;Q�#T�N������� �>1ޜE�{!�Ǩ[���\�U�����#k�p�nju��)t�R횽�;؆@'��n>,s{�����=oj����#��7�m��sp��D�`.�)�3(�
Yz)�DW�+-{0��m�k�B�t�޽�2�Y�捴4�;�^]�բC7�<��6Rru�t'�w�
Y�gH[bb�ь}1q�,df��um"�Sg����"�f����r��ۃP[k�Ar�l���4g�p������5pX(��[�6�u��Gz�r6���`��:�^ٍ�|g-q����8��V�:��3J&���H��m��q�f<�>��=a��a���}W6��;�Oo�!:�O
�G�e�WM��y@z�G�]^0��W�`��q2�vUS$v��u�15����wo�<=����4M�Z��[�z�ė���d햏��� XӭP���:H�)��A�F��]�ݫ���Ƹ����:�N��$�정EM:IU�0��Zb��7��(�ȹb�[�܉�[�Bj&�b��-�ƭ�*�	Ŗkn~�hɇ֍��sי������ ���+�9�
�+�r�B�R��~�"|+���=p���7dI]ѩ]�Ts����Ž�G��w �:
p�Zk3Z�&({�����B�dJc�=ۥ��c�z�FքDT��<l�˧�F_�P0Z��o.JW7i�Im�����]0�]1�Bs&)��ӹp﷛���g�E�J�J�2`>>>��|�`㋳n�:Uވ�.{�h��K:0bSe�N�7,;�0�ɚt�����K���*��^j������1���Y�y �5��9�N��N���S�ݘs�xp���Q��ם�K�P(��k�z�a��qY�7N�
�_K�8�\��&��������1ao����f4�d�X��A�2!	�wN�g+��ui�y�di3:�Ȍ�����S���,��4)v%q}C4������eI���Q*l��T�^/ػ��z�g:q��s-˄X�V�x�|}�E�7Z�2H�#����x�^t_/����o�/���v��-Z����Ky��/�*�Z�NOc�v����!��+����[.�(!&��\�}�y6c
�Tڵ�B��o5��i@��L;����jD<��i&2~����f�߷���o���sO�r���B��o�iO'�f�I��c��}��U`��ʹ����|}��=�K&�yh����Hp�^�K���.��I�\,Tڨ:��ux�k�Rۈ�Պ�KU���	��_q::^ �J1��|`�3��8��mUÒ|M��Z�ٟ�*�MU�Q-sױ�3a5�iH!|YM�УY|��6�(E���{ab�>B�`�ܥ���
�	�WÜ)Y�5���������SX��ٽ��Ydr�(�JC��ˆivჴQKЭ����j�����w�7�
?�8i/:��^׆�qKE�]��v7i�E�y<,sݻ��C��Cp�A䩗��u�m����:{����VWV��ζ�fh�(�+����������%$L0�}�xce�'G�x�Z�����fx��y}�r�>��jf�W�љ	��g�xy��N������{=[w� 騄�N�/��g>e��BY��.#�ʻ'������9^����qwZ�~�>w�gi0��~c4s�f����o�r�:�px�qD��%Mu�%d���.z�����k�]�a���˙G��l;y#;*wZ��3��eL�n`�b�t�8xxNZe�����z�ls/ia�l�n�WX��c�*h�^��}����^��u��Ŕ��g��P�l�^͐^8�N����3�~x׺Z�wU�:�	-���i����_]��O�5�f<ռ�s�s�����]WD���N�������oE�c6�T�Ly���U�	rI��(��6zөT�k�J�\�F1Ŷx�&��G�J6��&,9n*�r��/�;Wv�w��t��}�:�bN6��f�K@�F�O.��*�8����.
)��<�*Br��N�yN>�;v�Y��<���??��i2�˚3���TSA6�=Bn���çc2Q�b.*$�3���+��:m��H���~��	.a��+��=���7
;3��-�@uX��a�χ�ܱ�T�e�lx��Eq�.���~�l���zp�d��rc�2�n"uk�~v��^W�����<� E��֏ki�+��������`z�+�-���k/"���=]:l҄n�>��΂hV�u�+�LV�������@�[>��	�m�4�9�/sk=��Έf���Yx�0���`g,/�4r ���p;&�ec;Y�|8��I�D�l���XW��p��p��x�wC��32��],����˧�r�ϟ���9�(��(�Hc��.���]�p<��:kf&��	����=yh�3ؙ��*�^K6����p��q���.er�ټ*�i�냆k�g�K��/��jcoaJ{��M]���X\]�`�<1q����>-��\t�tW"���W���w��ֵ�mJ`�W5��πX(�a +�&ʦ�ܶ�����K���l���rۧ�R���&�����G⼜[W\�R��,����_;"Μ����l�
�v維���Z��ރ]�a���+5��:ne��ۓi���z5I���<�ذ
s.��u�'.囤2�n�=���_�D���k(��Ӟ-Y)O���X��o�xoF���T�KOn^��'��E�W��v�][�`�A|�1����i��Sv����R�k���ƍya$>���F*�Y.���V��n�`��V+�_���=^��-�;����9�:���R�1���&�I߭Y����E���ߋ;��^�^yn��~]�o�b�,�o��[�}KQ���^]�B�J�����D�p�d��4��]v��>��]��E���d�
��������AR�k��Tq�c��x5;��ȁ��;���V�̩�ۑ�QXG��[�x)���熧vS�,ḭ�}u�o�U37�-�UJ*dfa�c�.I��X��Զ�h}��1ܞ��)��ʅ���A��v�sQG&��?�Z=����i>[�;�P�Z0���Ts�e�S�r�n)������Źض�l������Z=��v�����u��k6%�¸N3.��	�OG�j��.ޚ��<Z��[O����>b�"<	�Է����c0�5Yh8�%����_���Hr�blm�==�E�1S�q:ʏ���_jC��FaXB�[���7�w��/��οt����
����LI�(��5�<�R�m��;���l�FDЉ~k��_��l(�,HH�be7�g�?�B��թ�ӧ�D���,��վC���vhC�&�uy+5�F��CS��ѪTF���tZ�Fl����/ x�@[r<t�D����⎍���L6̆�,X@g�PM��c����מw��WL�~}79�)}�{J��f��z�n�C�ǆuv�9�
��
S��0͵���9�䈈�
�b�q�����R�+td~�{ee���l��~��|����&��^W��s�zz�%e{�_�Y�2�=0���@�)�U
����)��Ȱn^��|w��$!�]���zq�����(p��|&=���\�˦�w�bDx\��:͗�U�@��AHDKrGְ�1$��Lg{���0K�#��v�X#)���\���t|kg= Ne��˻�T��&��ղ��nݗ��m��P�L;�D�G�vϱd��f(���z"�R���s�
^�����j��b�X�7��������1P�?߱��-���g�5��V}���kV3�\`�}[�i�	�A,�d���$T-���e1V,g�|�2��;��-*	bk=y^�.�O3��7KX�w͊#�Ѭ�#`])�c�#Ц�<<��<��!��LьHQ7'/ݟi���}"�hl��Ȱi�k0G�-y�5����G�߯�Huw��\�'	��>�'ܨ����,=/�T�E���ǲFyz�~v��*��5}z��:<@�s#G�����c*��~}��'��+�{Ī�v���׫yB��r�E�?<7t�^�q�YJ
�̧�Q��?Xt�� =6u�ӼR�Ȳ+^bwY�f�l&=P<��mlҖ��@�s��D��mG�3�U_���&�;Ҽޝ��+�G{��QU���w[��R���^�`��NuNG�:Ұ�fl�X�U(Rh�u1a��g�c[3�R�K&�\�E'2�ջ]��,��������oY �,PJ��se���5)��&���H�ɫ�CYD ����h�}YPX�}R���oq,�.>�"�|-X]ٰ1kD�=��H��c���K�º����)#����U:���!�^�Cl1�	��Q�ٕ��]u�*�,}-cfv@`�X8��{k:�0�&J�㠮����v�ӨMJƋ�i���t-�ЇC۹��$E��eb9�c�����x.��}:�5����7;x������k���G"�R�s���PA6b5jn^�rr���뭌�ƌ�ٵT�_��X�T���&u�d,e�_�,'i)f�@h���
&��}�\(��\2�7�m�cKn�
���c%���CCv���gWJ���D��^˺��;3���&)���fMb�b껾����]�TQ󾽛�ч��۪���:�v#π���@Ս�_�fR��>��\��fed�q��!PTa��DĢ���n�7;��<B�	JT��nf�Z�"�Y�|ٺ���5��].a�5���)X�|��ktEs�2SN�9��lYw�:A��
��0RF �F^[��iS;�J���i�o+���,��oQiÔ1c��Y��Cgwc�Ū]+�t���o\&+���-��'n�f���z�a[l��]�dۆ��ɗ`b�K�2�,Ogmݔ�!�{�W��a�B�}�z@qt�z���bЬd��Y"�X)�jE��)���2T�xT{u����Ǥ�˦�ڵv�l��W5vq��ˢ�ç١L7��3.�%�o�}#m��j	��gq�w�C�Cǜ/7�n��Tvf���b�s�� .��-b\a7g�^����A�Nw͗��v]��рh���7%1���`4>�wݸ2#%VT�����M]3W3BA�ur�Ff�9�
_΍
=��-a���x�3.��l�;�i4VoP�-v��&�u�޳W������h;4"7�-cڅӛ�]0V��6N�3�D�R�1g
xVIA����A��ؔbTpr�m���s��"�c8w[{�E9`t�s��P����ѷ�d�ӛϴ)��n��{ۤ�cM�o*ۏ�!�v�M���h��|j�e��z4� �tL��U��NN7�]5t��c5����=��FU�X��.��7�eGˤ8_t;�d����W�E({)��l��Ko[�k��=��X�.ݫ٩Q�֭�z��*Ka�����ּl�������uR���Ww�Flk��)���'����� ֠�䙽�L,��n_!��ƑZ�	�ɽhS.m��x�^�>ǯ.��Զ<�u�֦���ݙv�Q�0����׏�u��'Ve�GF��ưEvɪIz�߸��¤�u�+��w��~f4��n�I%�஖bbj�U���P�����Lg1�E��*�;f���c�6P�j8�����V���V�ٸ��h�٨���\D*�����������vS�kxήu�]��� <<�Y�d������)�9a�n��6­2�p�b�qH�L����[<�9׊��X7�G�a����-���]�r�(�4-)��F���x���Q��Ca���	�4�u>��T�F?�8��K�O�u�/���י�"=�y�:0K�(�ދ�?X�6m`���:Ҫ]�E����Q�E��v��C�
g��� �u�m��t��Y�}��c��ٱ�d���]���E�M;x�<�OX��V����V��n��!\���h���,���&|&�N�X���~��
�X�~ӯ�kAޤ�.��"�Hw	��G^\����w`�=������Z�Gc�Q�{�u=4Έw�S�=�U#��zc�&6�p��N��5�2ŷ`x[v����Ʈ�$�x����U���c0��T�d-w.��o�^��v���b��a;�R��sRẓ��n<k8�xi�l����̵�v��=�D�oϮ����e��°U��31���Z��?K��rA����?M<�����6�ҭ*
V�XD�DM����M}��M)^��e��}0�ړ;��Z���k��ɤ���uLne�f����1�BB�!D��"sz�u�ߏ�?��Ӭc�*���R=9��ofڼ���u�Y�[�A�g���=�n��jVX}�ך�6>�����=�*$�7��PN�R�d'I�pnr�
�)����g�S�LȻP�6�H��QШ�
��S�k�|��g*~{U8=P��'�\Y<E�alj�b�)k]�X��O��君������`i��L#�إ��'�\7'���[AmxW���wY���Mv��@V���Ag��d+�F�9*{-%�e9ixrۇ����LF�������t�Q����le�?XR���[�9�oY~j�6"�*�:_C>;��{��Zܹ�O2N�Nm.a�l��F�V�R-�)�6%��zs&�+�PK75,���9N��s�Xo���(�%��-fs�忱�L��I�b���dQU�%��0��M�f��^i�65��;��e����˔�f�}�9|@��;+�MX�iͪ�� T�����a(��:����?�c����q����^�һ��1�W3vzbW���Uc��dPgb��5m&)���#��ڝ��(:O�6��Ѫ:]�2�{�~a�߸o���$��6��]}��a��O5T���t����]����3�=��:V��8eH*�[��s��6=�]�8XYwí �c)C�d�\�o.�|��1����.��,�=��wk|{nI�0Ģ�}]
�c�ea��h�;���ޣ'R"һ�8|�-�n�ż��}��%��(R�,_@ŝ�6�d#Ǉ̞��\_�\��/5��=���TcO^1]O���e@�4���ۥD������bvwk�A:�M�wQ�$��i=&͜��G�B�l#�#u�s�3=L;�ɴF������O;����Y�k6�h���ם��L
*��I��Wu��=�+i��r�wo�)��c�;9�nr�R��\3;.�V�}x���8��VN�/L�4l
E���i�u��E����#bA}ݮ����_U��W�Y�5u�X��;؟���~�9{v=@}D�/�%�b��Ay$v�h�?�����^�M��F�s>(֩hC�~���L��G6]_�|-!��a/������#�
�)�./��OD���i������F��"��S�����5g�lC(.S���^ێ��Q��J�r����+.��2�o����\��16	*���_�o��շD��C���̦�^�Յi۩|�z;V�:@���V5�ͣu�$b�����#T����e�����S�1�)NGmv�v�Q���7keiS	��a2 ��s��i������8i�!�����6OF.�ӐRU�2�2�Q�
��oZ��A�׻����0�ʨ��]Һ����N:S7�CM�F�:ۺU����n�+�I����q��)�}!�D���n��+}�oQWxyz���]w!�ۊ-c�3ޒ-��bċ�u��V�;M5!W[W�V���11A��ޱ�N�e�����e�8zy�QO�)js���sJ_5������F��-���� �1b˧2����:����]	��)�͈�q÷|�����[��͖i	;h8(��r!���\�����\ф&��3��`x��!�G7y&�r�O�ܐǰ��0�	����ֽpS�Q�ˌ�7�g��4���i��S"2�㑊���i�0�r�KT=�M�e�� ��Ud�mQu1��rvoYlB���(�N0U6��8E�� 9�_M7����ZM�����{\�"�as�!��2��������\�u��;�{[�e��X�uה]m�hL�c�r�T~�+z�a�3�Ntj�=��1]'�
l�;1�Z��6ds����!��뀮 3M�uͬX��\a)vX�|7�8�����~��#��K�Y��-9Az�~k�`a���k�x䥵w�+*������7$�������&,w��~m�Q��!���iN�4�o�&��l��{Eb6�Y.��y{��<D��	P�ڳD�$��DG��"$�����EEiP� b78 gp،�sِ��S�v`��ޱ�)���7Y���~N��7�qkW�O�z)D��q�~�����T�`�x}0�9��ފ�}d=����^�rv�sT'?��452bܦ��+K�Y�U3�A���A(cQ�u��UX�Wf���3�1�x7	�f������C3^���ٙ�q}s6�gq옫,1�K�\'V�KM���z�)\���w�z�1��TfZ�!zʩ��^u�k��Y�K�Tn�8x7�a���T������\����+����j~C���>
�x�q��.z��ՓbX��糝��]Պ����?Aw�:`�ݲA�����{����d�"�7�� x�m��b��N�DX��e�M����n�;�թ��k���=��9y��]f}ϗU�0T䝻�}L������>���� ���{ۢv��(�0K���ߟZ�x��G�!z�#�_:FŢoPo�ck�8'�v�a��Jz�h3��(iVƐ�3�{��L�eЇ�7�z:��8hy�l~�Z}�z�̨� ��ͥ�:�f�F����a�����SD�A�(����W�����/<���U���4 :Wn�w~�0�E�n��f\(ǁ�!�=�kq-mR٭�L��v�o���P+&o#kP��>��F̴.r�l���m���p������%���"�y�D���*O��� 5J���ixr�s���Mܩ�ܘ蒁@�(;q�=�1
�5}�s�<.�󼖂�ڳ0���[2��"���{��*��h�Xף��`��@�w;�S�d���i��Ѹ] �W�akҶ��k��3�p�gsDI�d���8���4�nC��ǉ%͖ E��tf��~���"���cε�Zo��C�[-i�}��y��}ao���"�d���K�����|j?=�v-�p,��K�v$����eY�z�_룻��	�/s-�2�4H� A���CDg�ŝ��5)\�0,m�Ƌ	��{���9�x1���h>*ڄ'�#cq\�+4�e�q�6�^�Wsi��Y�gQb��q��gr���
M�e�Ƚ��y��|/үu]x�!��O��@ַI)��X�tC6��sx�P�-�Bj�r���1����
7�*(W$D�@V�郘h����L�u�f9���r�ô�
��S�����M0��00&�k�2T8�Zr���5���Fۦa�z�)�D2G}s��U=��t�w|;*H`]IH�N����^vq��G���3AC7rz)GB�b�p������D;2mr���߶��U���~�]��o������LGTF�I�ʒ��&���H����}(���}I�0�g4�{����ȩD�߹�#s�9� 2�2Z��0�:�TIE�'����ň��V��XC��F����~��I��f��<�罱IOn4nF�-����]8��h�ۨ��Uxfk�%��c�|t!�0��si��ʩ���.��1/�Z�n��]/�+T!˜R��.���,C
������CѸ���D�T�e��D���7!���^;[���/�M��yl���jՔihS5ەݎJ��o��V=R3�k;H����J
�3lvp5��$�t�f��4�G�q�wr��T�'(q�}d�Ůp���Y�7�ڬƢ<�q@ye��M/� D��e��,�:�%=���h��쑻�mI�a�!��M�A�8˞l��\��+-��*�fg���eO|ƃ�)rbâ���4�`�LFr�5q�ޞ�i|g��b��j�ʸ���g��)��m����T#����[��K==���\�͂KX[���^��i�B�x����KV�����ue!���ZMj������q�9��{ӑ��1wu�j��hc�<y j�(�?t��>ƈ����_Zt�3}�,]��J���:R�z��.,���v��qY�[����� �zeg�!��m=v���d����ړ��y�&z\�ꉭ�M�P��|Oh̸�xc�z9�vG��N��_����ǖƖj[�Μ�{�n�?,�̊2��2�Bj'�h��zbj��ɩv�hg��C�c 5�l�L�r0��>��"�@߅!����4M����Cq�ms
�A����ی��B<5�̠c˭<@*�Q�"@� ��B#!���v��;���/{��O�y���3�Nek@t�o�4����ǆ3�^��}1h}�nZ<�39�kq�o��)��V�-��;e]�9X�]���v�:vC&Ed,����3{Mo&*�v�(Ql�c��oA=,�Tn��+m�A�3X��;N���
�����]��6F6Y6��0�~F+�ċ��1��T���\7=�!�;�Yh���ԃͺb�a]С�eB���Y��[?�qL�:K�W<�җk�9+�%u�2�y�iYmj┦�CǕ�7-��ng��2��)L2�ۭ5��y���%<+`^H���-�ޯ��`)�V��c�?T�\�N�h��)�t\�xyl���謏/a����A�%���/��=X�y]���'����7��/e�p��ݻћ=�K4���6����:ϽK�*.�^��x\*�;��d���֫'.4�0��m0��f\A]{��~�F����S���(��I=���'޳:�����0��g����_���,Eɪ>^&a��Q����^��}x�f�+ݸ��z���<�vk��6��ʺ��jM� K�����h�5Sz�}t��[�)"�帕rY* ^z��}�<�즽}�:�9��u�z U�Ҏ�� ��W7��i^�>����μ��w��iW�����f1�����M:u��^*7:ڤ�<r���Cj�(Z�}G�T���Y�fņz����m� !xL��VC�v�30�c�8����p�È!���ͪy�#,���$e��v3A�"[8��p��q>SK_QYQ�^5���5>�n~}j�u���� �~�L���";L���܅���m>ď��� fa1�$Y�rkz;�
N��瑣�$�C>;s�fȭHS�̴5/T�����w��̠�+��r*��g�l���B�,�r&Q������&u�>翩�g��]T��˯{�ט5�[<	u��+|�M���}�ϑ�z!+��a���@�53��-z^�I�)�_PD]�~��?Q䟞�M𞥯۬�[�d�5'�"��s���< ��N��;��M���é�㘧���Os5�����NsC{�c��J��`�ֆ�Wto��ב/���"%��Kv`�l��=+3���_�cwM�IN[+�jA {����wp+GnVV{)��E��P8�����i�n�gN#���܎��(�.�}|c�,����\Ȧ�R�[�Ȼ���4%�O_9馠�Иqe��ªQE˃7>k,!G��W�xE��Ͻ�|7������}ߛ����O��$$����@ ��	! ����		ђ Bh` ��HE ��H@�+�(H���I �5����B�����@��o���		'����?��?�ax{������?��!����?�����~�
"ٱ���[��Y_:�p[�&���k-R�(�'�wX4�$R�K�"�̻ݢ�S!jMS���7F� �p-ϝȒ;�=4ZU3f�9X�ު&����z��=�i}�H�<UW�^�1KH'�����M�۽LS2�ݲ�1��+Fǟ�>#U��ky�f�	�j��È��ł<{f%E�
bYvf�ƍ�H�^�;gU\�����l���1b��ibyH�������J7�-^��ٌ�4SƎ���̺�U;܌��ʭ8�rcyW��G\�f���,R�����ٵ��˃6����QR�V�VQ�XPL������9�54��Lԣ(�ʸ��Uำ4F^4M�-�E��GB�vV�AMWQw@md��Yt�Vf�(!Y�*�N4�.���u�����A��o5]T���;w�)%i���SY&�ei,���X5�.ܲ��l�.ȼ�!Ų���e5fi,�z�uzn�����wX`�ׇ7J�ڥ1ɗ.-_m��VN�#��&i�y���=�Y�//t��n�tMb�f-6Ye�al�����2ʊ���_�e��b��<r����+�j��Kǹ��M�ڬ�v��i����1���RØ�hb�4��f�T�U����(�fټoJ�1��J6���J������ᶦ��"op��m3����U�'lU��*6��4��7�
��A�(+Gi�ׇ,�n�1+"�c�x��٣X��Ea&��f"oq[I�B�-T���$vCT�oU�Oo!9�S�D)��.�R��P-É��M�m�7�e��Yu�TN�$��4�H����)����\6��%���M��c���;F)��kŚVF���F��Hl�F�h<�]gئٙ�y�jZ5b.��Z���m�F���-��ZF�VEͲr�qC������ "HH ��D#!!�d�K$ $$"@`HFB ��� � @�d$��?����B����?����MB$$��'�������aM�o���		'�O���!BI��5��		'�/����~�sf�B$$���B���'�����!BI�XB������?�������d!BI�����O��O~@���j�!=��}���
�2��gX�b� ���9�>���<����-�T%XU[V-��T�c64���h�V�e&M�0�Pm��E2()��R�U+6R�&��B�D�6X�=d��(A@U(���TJ"BR�)TDT�*!�AD�P*�eUP*B�HH$]�R�"[h=ۊ� ���"�qZ�w1����)�:wkgJ�WN۶ɲᎪ��]����Wl쬺���j%�Z.�[�wS{��]��N��
)@m��b�D�P���B� ��    0�vųMۊ�jmݻ[���=��-���b�[wq̻b�k���^�=5���[$�x�����[ -dª����E�[d�;�={��T==(�y�oozju�y�ҏ^�+�{���z�t�z=՞��t�0�7���+R�HjA��H)n���ݼ�t+�`�vK;=����7H�T�l�-*���O\Ov��m�7�-�Jr�K�xh��J�@�J�ޥ���[�]�A�g�뗚R��g���6`���n�7��nw�x&�5�y�{gV�)MV�����5�i��y뵴=����P�b�RJ$���e՛׽y�P�=�Avkm���%JW���kGft��)�y9�-�מ����{��D�=��[�  ^�EJPD��ڂCzޙԲ���V�{ޯ<��������m��x��\�����Uh<��[��/z[Z��N�m��a 
L!{5)
�*=�]����`<�G����AU���Km%/;�yAy�y:S'��Wvѻ��z�� /y�<ҁm�@%^�UEUH�/+��^a�eI]ޞP=����2�+�Y��"�Ź��[/�sʔ���褩{{{��Vκx�NxJ�7=�( J�B������[k���=�%K����i�=�.�Ey��
�#���I<�OySb���{�#�G���+6�/w��ke	�O 2��@�"m*JR @OLL�=   �~jR�  Od�UM4�a&���=@ i��^�y��V`�d��� "Ed�����(���>o{�w�}~���I'h��@$�RBH��I'��$�� H�!	!�=���'����9��wf���PB��Yb�������.��,v��l�Z�d_4�������;�i��u�����v{륪����k�Э���Q�8,���eiwO37x���w�{�]G�m�6�g����i�j��a�n�L06�Ր�|���	���S���R�h�u����K��y�#�F�G2�+��U�Gݣ{}y�V��"�Z8z8u�M7�n�ۻ���88r�VЦ���ʰ���7/J��Ԋ���\_v�=��N�+9�k�r�j��*��(�b�1`�No[�s]�;��gw���.�Qoֵe�ݘia��:�
b���ۡ�=f��YwXx���N�j��U�3mh̡L��2�^S�^Q5t�	/!,] ǀ����0-�x,��mg��@���'���,����J�{�갊²�j|��X��W���gW^+䀧[h�i�U܍%z��-+�1��+�e�^a��9ެ��u�R�˸X]�ٺ0�~��T(�ŝ��f�Vq��֭�yԕ�?gg.�|)um�M�]� h�.Ϸ�l�]��{�Q˥��Ć���.�W���30�[[j����-�K(%�GV���:UvE��ڪWE񾳼���:���/���h��J���,�.�S����a���Ro��ٜ���-b�g�;F���gw�㣥�8{�='�����>M�h>Ρ��y��րB\�]����@5�ŀVQ�A�Г�\8��j�t��`j�XN1���P񩡾9�D�d��<��sh�;��^��j=G.��e.�L�5��j�� .eR=H�Ǣ�`'(qF��G�F�Ł��I6z��x�	vS��v��(�՞�K����eH�:�8(}�y�z޷ac���{��l� ��޽���@����m�m�]n�3k�5�7�o�և���l��yoe_2�]��Ϟ��DeX-�\�p[L��J��Z���w�ҫ��:�O_Z��f���үm{Z{hX�:`fu����.�ζ���w0��4�z�mށ�v�}���v���s,%A%�ZSuvv�>�r���]��G(wwS
�f�hT��k�n�m�ط���"wl^u�/R]�t�7Uγw��ϵ*�m��F�+>=��YD21p�G��}ymbme^�0�B�#v�%B�1�8��{��f�Y��6sz���o8��H��hY;]DMY��'�XycBf����
k��`��|P������!��*o�v�c�����Mq��Vn�k����@6�YXM�OǺ� �6u�W"�����u��P�H�F�چ�����g�ү�ǚ9л�h:(9�Twu1.w<���]i�����&�<�wv8�wǘ��PHVI��9Z������Kl`�$�mu��4,�H|hݛu��<s�u�g���;�������g9��lk����ZO���f�b�".�/V����h�I$�B�ܬ^5���ႯZ�}F�je ��՚����rgmн�'$Z!V��'K��t�\�Q9��I�g���]�<@�Zr�*3�2i�w�@H��.Mr�%EӬy�gRƑZN
k�eme��d֑�n�rk�<�J��]���>��X뎌� F�ɇj��q�	a�շH
��B���q�ʵ��7`�լ�b���9�Uej�G,\��ǟ4�ѧv����Z4�@_hguZ�I����ͺ7�����>�{���~�_l���Ei'V�ղ|w�����֓7z!��L5��Q.s0ދ��Z�X=<z�2��51���㇝�<yI���w�V�s�X�4S�.��V뫯4;b���Ul�=���D�]����Z�v1wP����c�xv�V���J�U�F��(�ܫ���QEDQO	��m�[ΉN�R������η�U4�����;VyE�T�u�	|)� ���m+��f��"鋺��Uh;�=��ꕲ�>�µ��_��[t=c�Ѧ���f�xܾ(�N����k9�
q�f��=M���b��ʮ®�ѡ��.=K-4�9�/t��n�]{�z��`L4,�sNe���վec]a��ۥ�� %��z���Z�uު����j�=ȊT�pIP��*��H�wUcr�����uj��gN+���p�j�S�ZE�}V����v����+M�b�z��j�y^$�3��Z&��mo"h�����em_w*�@��q=�C�M�Zǫ��L2;�/C��y#v�|q!h��2��Ђ�m�O��C/!�����tg���9����:��|o^琼[avj�Ru�n�Zx
<���c���ʧM���7�RZ�����WW��W�md�}��)h����CG���܅/��_e��i�[��+k�F�&�-`v8U3�6��U*����.��u���Q�y��e7���	��]�=���Ӿ��H>�,U�%V��D8�0Y��z��H��6/u����icU�GJTZ{[��F��h��b�I�he���Ò{z��:��Y4/] �>,������U�x�6=[��g-�j�C���s�;�m�J��m Pk��P幹I��J�y�z��ڡ�,m������B�^�.�6��1V�4��E�|�on0/�m{�f����\�:t���ìu�h:�;�$���|>9�nu�ڳ��dSB�{�Cq�x����<w�U
��3	�V�1ۧb��6�����Ù�b���K��L���'u{x�#����|��(�s��O�����ms\뛵�o/ |H�}ˋ�C����y��y��WOy����_qQEDEQ�neE�]sI�w{������;4a����;pÂ�.scޗ\�n���\�Vq�ч�����k93(���s����)l.�:�sg��΢.;�yPD]�<f����;�����<�G�=��{w4�G�ee�Y��m�*N��v��|�l4��q9���r)�%�9��9���9�f&���y����sxᨑDDc�����q��n�8tӧG;�b��J��Ĭ]^
�(
��YN�z�f�)��q�������֗���M�&��`��}��8o�؛,������<��t����Yv3WV,����|���1EqB���>f�v�+ת��!w��]wæv�̯�J"�;3�뾼�7x�Y�U�: ���h�[�n���ܕ:�K��|������M\�r���3Z�}���t(��߻u�p��Zl:�N>Ļ��1�H=C9�Z;Y��Я�v����n��s]`�Z6o�T��$DP�d�40���k�����s�h{��z����wԝ��QR����՜{}�3yL�j��um�Z�^�}t�5�SGXmFAn����/.�Gϼ��3]7�nm���]f��p�$�F�b�2�V$㝘x=t�:ݡT(gk���N�|�*�j�Z�W�ZG:ۭZkn���N��m:�eu�CV�WJ��b�z6���mwZ즹��v����օc����Qm��v��%�k���{w�Y�v^:�ַ��}{�z���l�bh�(���;{� �=f���oU��t3.ҷA�(!�n�j�:�@�yux3�1m+���Ubݺ[��4�u�[���`|�`�J���:/��5cHҺָe�{�����{{���Z�N�o-�Ys�k�.�n��\���DQEDDQEQAEQEPQEQEPQEPDQA�/u����{]��{5Ԧ����PQ���׳��q}Mkt�o��8a��N,MD�+�G����jS��{ٽ�z÷��p�3wPj(�`V$QH-L��<ٯw���q���+&���&�R3X��𓕼h��`oل5��aos
��s�����DA��F#L)�Q��ҭ��i;�kiP��4u ����*��g��������e,=��#�1E]��`��z��_m�����O^��4��UO��IӺ�����>���eeN�;���]2�ɼ�q�C�F�{�|�M�BC0E)|{4g��W����SH�D@F�D.f���ú����v]{�;��f��'�"""���6�5u��H&��ij���ŞWY��eR��h���-?B�:��ʱ���T��"3U�1H��5C�K�B�g��/��u[Yu~� =@�H�A��=�*��+gC�uz�b�[V��{y�sW��v$D���FDb3�3DpK�.<�k�n@��Q�o��p�8*��
�5�i��f��-vg4yV6s���Z����)���vk�$���Ӯ��o�2-m�"뮻[�ٯٝ�8�yU�i��+��+K�����ރ�����z".����5#���i3�i��e*"�}�9��<Sg_{����9̻����`��o�^��ͯG3��te�+2ՎXe�Ma�QQ��h���=��Z]x¶�����������B�
w)iyw�c����]��`��vz��� h�b�3M3^݈�9¸��5=֬��غ�K��QOi�j�"��=���ȢiWm�i:0b��H���_\ֻ��q�A���DQDG�5���;��[M�7�f��x�͜;���߽���q��N��.��`�c�Yt{,�:������K}�^,�����9�p�=��Mn�':�{���g83<ؠ.DAhD�/�(o��';�q�tk��;���S�uz��oy�i����Z�+X���M{�swI���W����ӽ]{��V�PD�}�K襕گ2�9�g{�V�oP�=���{��b�1�!�{&����d0Cݽ㮣�`�(��xn���Պ���XkH୷զ�� �>�-)sZ4%�5�s��Xq꺢��T+1�*
߷�I�[�H`DR@r��F�]�*���4�<T��Oo�ZM��X�:��o.��6{�jY�[}�@P�*I�i9��,���N�P�֐��j�5��[w����wD�o�/z�ɫ��G�z)SO�D�`;�@�_�WW]f��]�55H�[v_]q#WUu~�^��N�߆]v����^:D|�h�8מ,@ ��k]~��b����hq4���toU��K���!�V��S��z�t��h��Z;�=��]�̋�{|З;�f����p�w�SVx:�E;y�v�h���twk�����뽬�U��j��������7ώ�w�kJ�ok<H�pls��F���|�����m���廚���] k4b�ɒ:k@�ֈ�Ŭ���a��.�g���hem����|��6Q�ZiWf�mE�S�ה{3�]�H;����;vumn�V��up��Q�uòm��hSK��A�oEj�}i�8Z�2�r�C��[����bζ�u�Z�m�|�������v��ŗC��7�Mg:5ɍ&��
�)���W�]л�ѝ̷���Y���Kʺ��f&52��k��6�򺬪N$
Yzs�����ʇX;��kK�֝^J��GFq�6ss�[K�J�&��qv]_�F���Sf�,c��$��g3=��<%nk^��󝪙�u}�k/��us<�{ަ��h�@�:SIW n�֎<���1�q�g�nX嫃����p�{�E�b���fb{�m�����c��s�������f�]�.�����a�&�m~4HAk�A�h�G�ڼU�[��,��F�l��V�UM]s�����cv���`��kҟV;P�t://�g+8ֱxJ�ya����h�YLh�v��]:�����U��W3\��kGp�	\�t��C(]�+�a����k]��<���oA��E�#t�s�gS�fk5��6���E;�ӽ���\pS�2��x�_��>�K)�\f����Z�C@���F���@=ZE]]��]ז�n��-��m�}o��@�k6�"��������vI�M�p���˘�"�3ʬ�յ��WV��Z�vX�OR�X�!֬�2�;���+]��M�<�ѴsV�Wǘx��vm
@�*�u��u^��e: >m+u�aq�k�Y���ڦx��tV����tXF͝Uc@o5^%c��� s��Y�uލ�Jn��`W&ض/l��X��xq�+L��b������۠�|�m�����T���lM�-^�X�sY��ކ�^��'���}{��
BӮ!�v��=��Q�ƾ�,~x{u��K�+�oP���ưX;[�L�Ҷ��+b���9���׋SF�.m���[�@����m�Ɗ63����W']Z,����TB�ү.�K-=zG����m���o��+=i]Y�^�� ��E���[�������n�r=c+�A�yVk�%�Z���D���i:��fWr��^u���X��b�#p]��(]"~*��o�:�.�E�g
�N�P9�up�8�ww��SZ��s+4�9z<ye�ɝ�+�n��2��-P(� �ڱMѥD�|�W^���a�N�>�>`a���.���}��8*Uվ����%���w_.�y��� ��=�N�to�ջ�(h�c�'���N�K���Y˫������Ǥ*���i\�������Tm��Ю��S&�����h #e�h#3.�)�:)oez��:�[���S����YGCǘ�-��w[�Û�]�Ϟ3�W�Ōo8f�~�
|��:�	�]��m�=lvk���������:�E�����V;���%�K��e�S9�M�-^���;5)�z�����]%{��lQi����`o.���}��wz������ކF9QA"���̬W�����6�ݼ�ḃ\�{���9���K�y����l��|������ϡ�ξ����˗B��l�g[�'H���S���a�t�Ji#	�ĢQ�I%��$�}ۯuwmjw�GG�q;��B�qm��S�l�y�D�n���xNl��t�"Z��9�����g�e��H��b	���$�{�mF�H��L����JM%�����,�2�M�jBN���Tf��wYM�:��3w5q|M�e;��D�t'2�����l���s�{�\$�X��{�{������Q������c�0�;�I*�}�F����u��@��q�M���tΐ�2���-Ù��9���Bcn���.[(;��-Z�˽»Ows���m�iG����Dy���=��M�܉�Z�t�[���v�3,�k�4G��U���Wn�['�ur�û�=��͑���Z���ڸ���^vWC���m���K%���'�$�5�%��:�����JkE��r�MğL�`C���E,���5u[���y�ZH�&&J��^#�$	�m���;�vP��$�9�{���N�ռzV5��q8M�V�m�Y��b�#�%r�;2�]p��"�2�q�6s:�70X}j�+�w�e��Vs��V#�v����$S��:ݺS�-s))���e�iX��6����6e1'#�MVYo5.�Z���W���[}von��>�+3N�ͧ81)8������oU��m)"�uc� ��3[�޻hE��b�Ob�r�2�r���m7W���T;V	�IF@)j9��5�8*�E%�ћ!Ыh�TW=�K�xIWd�;<N�775�wU�ћS��ən�al��]�*��Q���Wϸ%\��f tI�]�o.��=���>����o:�<0��I�I�����kk�n���\R����fǶ�G�X*�j�z�;�0��ju���q�x:�pW�_sB��i�!\���ݨ�6hI+��̕(�:(�&[r����X�Ё)b=�>"�b�Ԧ#����Ja<yn8�g����!������xXi5�r s^�ެ{i#��ċϦ�l���y6!nR�׍��̼��(�1�I��h�X��yS[&F^��/�)I�KY��9�� �B�n�z� ��w<�M��m��p�+���˻3���5��9����}�fgd�/�%��p�G�>��v�MW �[;T�M޵�j���M
��	���˷y��i9�T��`�vH�b̻|�J4�3{���A�+v���%1kz�\oe[��N�嵼�q���Wv�O"O"Nؠvc��w(�'U�ŠS�����J�#쎱'���f���;��r6�g,�'z�	w����ԺI4q]���H⵻nmܖd����|��K�y�}��{�ۮr23¹u�s�U�,��гǵ��`���i���d����k��z0��U�i�:Oʒm�u��ML�)�����;��'t�'	%��^���dQ�۔�fE�VOC"�y7U���#cw��}�������1�JK2n��Zݹ}�;d�Id��z�+���ӱ7d�v]l�%ɶ���Z�l��.:��T��D�#������Y�6kQJ�������-�^�Kh+9�7�{$��/n���E��[к�C���2\��e��\6�󕓰@rU�"�#1��WIK"��v�ڗv)��a��竮akDL�ۈ����Kw�#q&��V�#�Ԝ�����N$�$ރ9�ƹ��FY�Jkӏ�	[uդi�G8�E""�7s���ی8���9���b� ��2���B_V;���i,��}���[O�n;�WS��C9��;gy�v���9#vw.܉����4�-��r��Өk3�\�:�:�!4�n �W��i�.�5VK���7sl$N�2��;��b�Sv��7�
�H2Y$�5i{�]3��0��͒2;�gn�)�`ܤ��6nZ�|����;DD��[��# u�u��C��w�:�"�j�v�����v��ٕ`�d�K�3�W��Ήe,H�uv)���u�N��n苞�ĝv�Óy�9�`�|6�	q�LSQ�7}�����^�^n�Ts�Џ~ɋ)nh*z�%��4;��8��z0�t-��P��}o�{n���m���7ԪG�,F� ̂㙋�@�Z���AŔ����z!F��kl-�;f���]|�@��<}Ks�&j(!5�c+���T�Z��p@��y
ua�FJ��G�ހ��\-��{��y���9�=<2��3z�H/V�Z�`\�H^�1%������͘�i+���qЭ7oK΂�\p�T�s�nt,8��d䠅����y9E��b85��u��&�h����Z��˄��)9浶3r2�M�v{v����{18up���u�:2��OL�m�x�f2�0b0V�D^5�0Vڳ�$	JW�hD�)��,oE�0su�հ�t�w�lM�ǜ]p�V���%�U��Fx�G���G5�ɖ����݉ݒ ���M�F�e&�	.��gFG��o���f��1˵���Űi����]p���ݭ[*��p^��-P�7��ҙ��a���'NV�2��Y:�G��̠N�{�ޫf�:�)C��=�*{5֧ǹ��a��MњCW�V�`�K0��פ��Z�m���z@����R�q�o�����K�	��Ύ�����Rk
��U��6��%ٳd��v����2���N�[\HN���hְ�X�$S�y��NHɺ�(��;,���m�Gi��%�˲��ψ��8C��<��Ȳ�=L���-�*�02`@<ٸ�gm9�D����r��w�î�i�':U�څ,���g[�6R��Ț�>Ot���K��7{I�ěe�����e'NN�/=VA��af0ef<H��0�k�2a�sRȅ�8�kĠ�oQ�{G)�m�����=@.��q6w��ʱqC���B�<U���їQ��,t��]����w<V��a�n��;d�ԯ7�!�g�:���s��+1�ҥk�3n�!K��������*�1^n©i�HFkF�Tk�E�ne��gx��6h�k;���,�7�;�` ��`[ =s�Ws�7��۽p�]lpv@�[ډ�XE�Z6�#zH��%e��D��q�`ㄭo�uez퍈`��gs�7V��tL�l��[�Υ|����t������ʻ� �Rs.��S�$�u�U�y@m�Me_n�x!�6���.��' mU��7�8�m+=�q�	�y �5�ṢϴmB�fS�"�54.�o�;��2��(�b�)�x��o��'H������7�E$��P]���BZ�-�l8JJ�w��m�e�X�a\��t]��ق��+y�����I������P��*\o�owWo�	�r=��]�n�q�qէ��� �$5����g\��GN��l��-�TO�����}x,ũ��Xr��h(%S0���v��0�v��w�՚e�唙�j���S8!�\:=����gFQC;�h�R>]1��8�t�X�pRz_e��7y�{���� ��U�Tg�,[/�9�kz�-�F�|ޗw�F�K
�G��i��w���4��t�t����q(���e�m���7â�4��3���y��%�m:��>+kLRS	�Or��8�]�XH�3  +����ν�դ��wmhϝ<1�Y�Q�ojZ(Lx�0�uWh�.���y^+���h��R�<N[�"``� -����Jw	�Vy�G��(��| �|r��؇,�����Y�.^��)�u��q�t����{�N��-&�6�Pn��"�T�J{�w�62"��T�M��4��f`y�5�ĭ^f�]�Z��P�rB��"O3���d�A�)٫`Kݻ�7�����q��R�A�\�0�FnH�r,s�L�Lا�Ba@�ѻ�"�;�-���[{��̏�&�f��i7��]7�;�9b�����e�z�!�
�.���K���.�{��t�<gN�;v즏:���rüo�Cc��h�1Y�:�@&�nL��j���u�4@�
���D:X�A�\2���X%ӫ���:!oZQ�Yr��|T�r;w�'�+]�:#���X�F�����m�a��In^u׭	�����%����yV	��-Q��X���ak�Ou�vri� ݖx�̊۲q�R�֞
�����
�1�G`MK��I��䳘
�Gm)/�|O�GLi��w9�2�0�P�3m��T\�Á���Q1�r��_nQZU>�-�VP�����/\�z�6tή�O��|�xsZ�:���;� r�H[	o��XHx8u�Mnɏ9�ͫ��R�e�����hA���T��N����k1>) 3�{t�Ֆ,wW�ݬ�v�ɮ`&��ۢ���AI��״�����p�M��׽6.���t���fF2�s��Ս�8�K�p����G5�X;�A�$�(%
WI�#�`��T=��],=��ɾ�����79q={�̔��-q�/!B��Y�Cv���˖m�5;�u�vev��%�6�)a�뭁V�w9��bB�[ےT��tZ�dq��r\/e�.n��j�6�䬁�8��zqҗ\D� �\�����y��m�x�¬1��R�-nG��y*AV"�Kh��Jź��9wՎ�����X�AY��(�9w*�7�غ��)__sw��ܻ�RY�P;�%m����1�k�0< �55�<Ӿ軚\6��*dM۶e�1����Y9�5h�+l�\��{pr��Ái>Y�c�n-�\���i��B�Fƫu�P���S���ݔiհU�d�&�R�V�r{t��ԍ����D��ϛTuZ�W����t�:��3R�E��f¬&�m�;\���޼���2)�7N1z�+A��4���첚���i���4�B�fꠎ�]�n&휂5���.�U���:�a��2���{D���zZ7E��V����2�-,V�����Q�)�����#7stV	k�n�^b����)mu�2#��0�R�D�RK�A�q�u�v5S7��
J�)���ΎcJ��;�
S'��/5g�0����кԵsU�;�6�]�z ��/,�os4�S��/^�ĴjR�$�mwQQ����2�wkN�vS//�O�R@M�ζV�j#Ov����ӫ�Iܺ�ي󬋹��\ѻy���xe��'ؑ�B�`��t��x��`�C�r{z�K�.gt5��iSk_4�g�|���6�+�iW ށ����`BV,�^]�ɸ�⃏%���V�6x�}�� ��X����F��N����<�*�EcT9FU��'��+���5�A��)T�T�ewF>�XVu7���J���vG��N�^�,��|���o[ʢ0R�h2)Y����`�q��\@�=�"�e��oڶx���e���0��ʘ]�V�vda�6S���f�
м��Ԧ�L��rsW|D2k��|�Z織�������(��;�+���1���l�K7����DA�7N�M18�Р�ژ��8���Mj�9R�l�3�o6]�Ev��;˔������5L]���֦_�+��CfU:��7ee��|;k�1��Tl��q�kP
m.[�5:�'(v�n�Z� j�Y%���re�)!�;�X�OwQN9:�u�:]M�W�4�+/k�Z�&� ��N���!,c`����r��9u�x,v��H�f]\u*Wv3}�[(�V)�!}xp�'I�� ]]���� +-S��]]��2��pP:�i�%��0�f����(�饮�t2�Z���4��0�q3���j���4�B¡� Ԃ��grW6J�čU���S�w��ЭM�y��*e�Fl�	��r�=u��B	����kf2�"Jt4��%��wf�]Wnܪ U���zm*dZ��죃�������TwXUg�,���mb�;%*�.��xe�oju�v���
L�N�1���wH[��*�9o�6wlZ�Y�t��ǔ$�Ȭ�*���
�⏃n��l7�ń(9����S9N�yχ5�vf��gMn¥�N�KH���{�ʳY4;�"0��v���`^7#q�E­��rt��)�9v-���;2���Kҩ��c��.��[�_	.�a<컷�
y7X����e$��7c�ջ�u.�7����k�ޠIS�����$V�yvLn��ʳ��b����c�ٝ�A�ٙ���R���r��r=�mfS�������4�m��\5�����Z�ℾ�h۳��ѳ=q+�Z������S�d8�>VVQR�� �����F.	�{��e�3�ņ�걬K�aVNQ`�o�H��s�b�g�0
���i�~	;8�G�ē�Hc������&��Ju�R�x�/���֭͐��}-m�ιp�e`�(�iQ�i_�A��W�X��q1x��},	�]�U��|���/�]���Ӯ�5#����d�tP�/��a��rՒS���1~�~�1���C+�yP��V����]yZ��\�Rþ����;N�"ޫ
�9�w,���*�mVW[�ʵH3.�S'B��l���~�wvJ�C��c�ՙ�8+���L�U�H�fu.�pe�Kg���;h�4e�x���k2�:�E�\L7Lv��c����]vrή�m�Fȭ�u��'�p��}؆V2�s���z,�$їp�ʋ+�E��I	m�T�⤳��SR�yf��%��H�Uh�h���łf�3�wR�@Yw5�D,MZ��1��Ӑ�����]ݪ��݄˗|�e��[�Eڳ3/%����Y�\��V�g7��:ɹZ�����6�9*���!s��^ʺ���L_�;c��ó��34b��L�es���KW{�Cرf��\K=�{,��2Ź-�]�7rV�����^�՗@���3q�������p�^�ە�]��;K
�ŹI*zwj�Vm����M˂��;{	�����S�lԭԥ���:_uu!�kX�9)_\b��م�LZl���j53_y���}�BBHx@$���#ވ�{��� |´�q��۱��ۧ�wq��cޣ���hi�p�'%�e�{;oX@�p�J��un�*J��Ǹ����Vl��AJ��/�ؾ����k���=�])״zn�*r[�'�s���Jmr*��p�E�ɝ�f��x��I�2��)���[IZ���>S��d�)�#G,�Tw�Ϯ���'5���c@���Ԝ��AX�7�4_ff�*�)v���2=���/�xۇm�9�L��'�Zt�j��Р�k�� �Ib������c���Φ�J�x����y�!��gb\zK�����4�C�r]�c�8h�@k[0ƣ������v_#�ΝӦ�:zhf��n7q����.Չ�DR����Z���K�v�A�Sc�:��S`q���o�d�V�ٓo׫���d���A��*��,�-�"�fKtY���-A�M\�8�h�'���Q�q�����3_EI2�l10��o�2���b����5�֡W�@:�/V�t���2b�^f���P^3�;m���u������kj}�M�TF�ͥq �P�h� l�G���>ȩô���d��4��勵�14+	��N{B�fG�SD�m*}���5�+|��#s4kt�c.�cԮ�(F�^��H����4��A�����,�ǳ��䀗u�V�P���_+l�4�N��H�I�qV�r�ތ�m� @���1�u�/V�
�`��W[���Ҫ�ު��������fy�M;���[�(�WV�<�.�{�̸k�����sl�cyf�-�Y�[�q�	Lfeю/�ow2��IR�5���$�m}�PX�ֵ��W�]ֺJ��+tQ�AR͡�i̗*�Ώ+AM���z��č��V�%�
�})�7՗XšH��G�t��AAbXlK%,k&Ա~���P��ԭ
v�s��,WX2��|�ʋF2,�����ؖG(���D��|�aj�y� �^�ml��]H5�;�^�Ue�͑7�)X�YΫ��:�ԷtP�9N� $r�尠'\���u 5� ��b��աdT�SN8��\̹���eFzN����U^�b��`�\�2y	;�_k
,h�ƉB��+y+�
{���s���*����-B��\b�j�G����Tk��r��G�P�L|d����Çq�U��]��s��껾��o�%1"�M2@�H����0�H�J2ZT��̦"�{�{�w�o���鳭,�zP�V�
��i�z�@u�&��a�j��� �h��Å�X��51��G;U��[ݥ�d���d��T〝Z��
�]��@L(S��kr�9�Cޡ�t�ҭ�OS�n���+�?m��:�k��� m
X�0�;W�UW��"b'�^ZB?���;w�u�By{��x|���Z1�a�Vr=�|�� <c��Yk���,Uy�=Mz���9W*#�W-�k���1��=���P�y�Y�z���ᷢz��ʢ�>G�I�����1vr8�S�H;��yh����S'"�J�>�.�땪\��@2���#�-�:�Y��4�)��Mj���۝"�Ȭ��t Q��6tc�tV��w}+�����'$Z�N�ǻ��Aݠ-ݑ0��a�N�9
�x�;]�rW��K<�iұUyi":�ϫﾬO�O"yL��4�w�q��GD�@�&& B�1���Y!�@��"T�d�D� �*�dn�&�&�t��@h+�b������U�&�S�{n��Ħ˚%yH��)P��,��D�]��Gt�)���m�\�5�8�N\��UG:㏶Y��r]H!$,5�@k��e���s��uEqlʔ�M%�y.���k�UW��#Y"9�-h�"yυdY�������նfme�Qǐ�P��[q��{�S�zCtT��P��X݇L�BDk�Dz<9T';Q�0&S�K��L��r.R<�Kbv�����, ���>6���N��˩y��R#�%�W���ވ�9�O�ބgm�Ne�h���n^i�ţ@��К}�p��rC�PG�{�e�S���$U7W
y�wLsJ���}U�b�Υ��qB��ii��-�ݕ����殑��mT���XvyD�E4U}u�u���T{%a~��C4<����3vk%�u�_t��ڲ�*΢V�Z�u�\_�80d����p�g���������B��;�he݌��n���E��@hU�.��w��͓]�E^=]�5ή�S:0���㹃l��a7!��NY� ������^���b��(Q�>�6�F�R��ޏ���{(\��pU�S$`�(K^�;�������ޣ�����?� ���2;��&�>ׂ��t$P�PP�h��BsqѬ5� 5<�饪)<�\Ii��	$j'�*�$�{��x�D���w^�{�}��O�E�ofF(�N��W#�8	g��u���J��ӑ72U��}p﯃ni�H���y�UUy���D���:oM�\>�FNFF�UKJ��i��i�5�c�DF��Ɏ_'�t�W����s��9�	Х�|A
H�0g������i���,�Oi���[ŧ�=�wm��K1UH���rx.��^���ˁ:�p��yny�����\^k_����� �;�"a#�7�n��r]��"U�Zb�%}x�Χr�̲-(�S�rU0
��!a�@ԑ�/B��a͘0
yÆͻrڦ� k��
��8�[0*N�Y$���'��n���'�X���G;�W U`���@��(
cDl��:$`�sB�q�{�,ss'{�w��gs���M!�� C\�9:�E`�5Z�\�x2R��Ba>]�y����e�}�b��y��6br�Ȅ�s���$�w��Z��"F	���p���x�J����(�I�G��~����&�au�h`�z�*�A�~��Gε
"IC%;a����s��.�4F��n)C��	�!����S��N��A�Rrԛp�"����U��';�Բ���j���~%ڃ�tZh�V'i���;s-
-�� wa�8��<�V3��}2!�G�����v���m!��@]Ʋ��YB[9����Ɋ�~naX
�1$Mڽ�2�XJd��AF.Of�g��.=��xǞ̴��D�~aLdd�2J�+eD��)H��H�TF6�K"# ,��e�JK��A�P�/�g���w6��T�E��X�Y.�]�|�/Y9n��F����N/w0�,a4�<�PV�I�9ƚ�0��j�٥ײ:��7�� �'KY�T#N�,@3V3mͬ9��Р%k'zr}�`�$������5@+�W�Uϱ�=]���
,'�{�W��Q���T�zg��HWL��|���1����3-SF��kH]��g8,�ݳ5^AU�W�U4�,٘
	Z�]ϭ���ڶk���ܵ��f^�&�R���J�f(-���^Y�K�Kܜ�P��N����
�z�<d��.�:Có�srY���,z��YӪ��oG�-��A�ٶX"T� sz���C��_{���j��oQyݭr�"�w�4s9,51�P�w@YXu��Fbb͇49�$��*��f�y��]OG���k�=�BC]{����~��̼��������(��$�obq�81V�9�����:��Uz��H��m�l%Tn�.�,]�p����H�ֲ.�n�̋�,�*�U��eР�\��hl,Y�����j��r`B��1k��pY[������	$��YV�:;��#F#x��������n���#��DU��TY)�͛/ 2��ht�:5Q:��ˮu��� �_
��Vpw0���ҳ:��W����u�F��h@�Al޵]�p*����mƮ�-亖fM��@[�Ng}ou�����^���? 9�	sh{:,/� K«���& ��S*N���M�޳'��a�2����YJɘ�\[qn��e�V*��z�/_���.�B6��'Fy�>�׶�l8b�y�;
�U3�X�=�)
8XB���{���p(�\*Rj�)T��jݧ�z=��z��=�(1�S�+R�3J��wh��W��"��a�vL����[@#�t�9v�=�����N���ԭ���VIͼ���W�G>��-���*�h��0��t#�� ���B��%I�YR��2
 4h�(
��٩Y��D����V8R��dX۷�WZwUv1��CK�[�b.m�5��r��m�Sf���:!`�{�ZG��*m,kL˽o�][��Ջ;����j����[��'Q�`X��픫QSѠ�~��z
�:+�a���2%�4�U�#J��>���Zl#/���A�b��0N�ѿ1�"}�q�{ފ�2#q��N:+��B��X�]ܔ q4eu7� �$6h�t���4���C cH@�]0�{����Uo�b�����.42 S&$j,L��;�n��ҕ�-}O��|M))�*'�ɾ4,dDz<�m���U1p{2�{����F?z=�� ��o� ��,w��k�7R���0^X�%�4� �(;�g��W�'�uwI똽^��LNO��0(2��W�^���D{%:���ّ�a�3ݕÂ"|�jT4���Vw``�ѼD��'ra -W2sK��G��rVO1�UUUJ�LynfB�VE1%T��dE`�)2���_Nz�S)^El�6��E9y��m�2:�"��W� 6^�ȯhW7G��;{��5)�/U3O"[YAZ�q6�v<;
�ʖ�$�tp2r������owm�i��0q���'�t��uĂ��bi�<9?G��ZY��C20}G��\�Rr�%��B�1���yC8׼'?��Ɲ�׼|L��,�@A H�뻈��k� d�@��zÿ����]㲿����G$�5.��Uu��r�:' �T����ax��o9oe���(�R�(0���{���E��0�����0iXD$ϟuf��q>z������Q�0w�d��<d�#j���S���^��Q��#�K���W��d�����L"��!җ�-N�َ�ʗ�L�(��7v,�".L�=�ؠ�k��iq4�fՁ�磌ܼExWmUG[~��s_NK/�]���U0�%Z�8�6;�7d���H@��*�aJP_s_���[ύk*{��Ȕ��|�w��E9����V2>�w�{�8]�.!��Զ�<7lthL��~h�.�wY��A��nh�[W�(���{�抖��!�z���T�.:\��E�z#����y3�B�v�л�����U���8{:}+P���:K|Ao�i�f�ٜ<?G���>��`�vUh��{��#��ާ܌��v3�"��M�+�:9�%�c��A\�MGp�2��Ύ݅���"�9�G��l{�t e���y��^Mz+1�&J̼
�UŕOs���Э0#����[c'cB�lH�{Ƌ�z=X'й%�L�[*�R�z+a�<��%أy�xAF�k�6��{��e���O��k��l�DN�D〝��0M�U{�^��{�]D1����d	/^g;��~�=�}��5]򋡉��gSɌ~��Ut�_�&><ƱJ�d�r���l�8(�OVW��G�ׇ��._��:�c�ꋸ�i��Kf;uM
�O�Ki���l���7*Y��.�I�)l|���i�С�9��v�s��U]ϹS�@��1��y˻s�=���;��{���B��g��C�{|���S��׸��u��E�=�5��ۊ;5WLR�c���t�On�������7Z�9�U;���Y���QN9��2`.6��9p�wl˘#4aW(��V���TETT+G+�����0�Y�a#Q���^7f��!�@��F�su�G�A�sM7n�v��|a^�|ոh�%r�U�f�B!R�-���\b�Q����n>�;h��kFܵ�0u6���<+����k(��T��G,�pͭ� �"�
-�#Z��k5�隵�Q;^_sIɇ{���Ӵ:�]r��F/�'�LSF�]��?���k�)eX��I�kk��y�/�o��@D�, ��#��""%F�җ��B�)R��[�j�+M�~��plVh�Ir�^�=�+�ֽ�Q=�І�$��s[��bt�8i��u%>w�+�o΍�y$ݺ�o7�s�T�5�P""����w���H�L�B�'l����|'UB�	H0Nxm��R�?}�x0^eٞ�z�c�e��P�O\3;Mx��U�8����[��b4Q�L!C�I�L�6%^�nɹn|�4if(�s�\X+�zh�q�pe�;!�-�$�VӕW��gF���o?�C!K��Mmp��=qTt��-U[`a��w$�y�t%�'8L��$�I�=�76��׊�N<g$�1FZ���n@�^"W�7+��:�|�ri�a�!+�t�ʻJ�0�=p^Q���/�Im�;Y���TW�ӛ��2�k]9C܆I��	G��e�.���]cH����7tZ��:{cX-��!��$ѻZo,i5�%Jƞ�9�| /�1\�SM���٤Yە6��㓦�t��c|�a�O,���y��q�yX�N��U��/�Y��e���Z�~/e�En�s��C����^�ۍF�0ƚx�S�&Ŧ>}wK��kh�,�v�O���=�2�W��:)�����[�e����{���0�Ss3T���iaf�	湑��C�`��ި�#��{Wb�#]�M�:�+�}��K���Gw�YH�����R�R�2�Ʀ��y�P�����o+us�H�f}R�T�\�]������+w`�8b��Չb��*�K1�<ɠn��we�����l�pU�����-� �ۆ��[�L�1��k��M�M�����t��.nl<.��ܻ�v�� u��L�V�M����G5�����^ F�=�������4ák����5�ʈ��{�b���v��eۋ^��0�ȝ^f�s���{$��$�$���9π�F��=ՉV�U�`w���y� �����ooBo���>/�IOu�-�d�+�\��yVm��p�(�'���Р�)�h�=4����o�����f�y@���CͬS�ͺꗱd��v8λ=#3���v�t��+J�4�f^��d�t/�_a����>O���'2��돐*y?����1�x��%E�+ۖ�P�a]��au`,��S�&�LV=
ϨP��y�!鎪�l�yu��6w��V{~�U�$1��C��M��A�O�*~���]?�>MjèLx�a�Hu�a�+���g�;��6�f2T]^��?3�B�M3N1Dx>J1���*@8��c�$F��"?e4�栺��$Ӵ
�>���'�J��#l}�YO=a�P�,���N�e�1'���~M:g�+�M��I�&������{��w?}�^~�!&�Qb��P�����I��H5�'���s�B�T��f3䗔}��B�é�Cΐ��3��=eO�^!X�.���k���}���!��m����>�c��S���Z��c2�X�JbLtì�k���`}n���N��'\�ea�+?$��ሪ�
�@bQcI ���"ȲH�X����(�H����6��a��'�c
����\��j{��?H���p��1"�)�Y�����AB��|�˦�AB߰���h��LO�~t���Ҡ/g߰��Xg�Nc�z��U=�<|�c��EGH�����C��O��m4�������+5�¸��3�vىX)�@_o�K�LLg���4��8���3���'
m�w�ܼ�^/��g���Xם��X|�P��P��>C�T֞d�P+�¥|�Rs�c�11�?1q0�?>gS�6ͤ�g.?���
�ӛ�{���������z�b��̬4��4��¸ɦ���&~�����$����������(��W�6��Zʞ�y���^���2��Y��4��!�+B���Z�4�Dp��z's8=	
�a��0S�T:�v�����"��Y@�>f}��@�X�O����5��%f3�_'��(RTY�ԘɍY!߃�ғ�R�LBK�"0���~�ݾ��3U�keB<�㔐N���H V��ƴ!ek:=�V����O]v4,]�������*E�gu�y��_"C��=��I��9����@ �`?��S��<�M$��g��&�q���O�o����J��I�fE��|�}�����T�|������f �C��C���������iHO<a+6�uf�1���Ϙ��m��:�!��,�S�9��$�'��$!�f��~a�m���﮿���u��P�
�aRq>j��I��%eC���L4�I�P+8�b��:퀦g�q��J��5�,?����!��?�c������l��<�� V��k!�z��ğ~��O��$�4�@�!�o�������&�B�P��`(�=a�B{7�d�?�������!���M�l=�N�ڼ��o�W��?�Y��/����O3�l�}�ɦ~IP?~����'�M0��_=��S�<ʓ����i�C����I�ľ�ɤ[�w��_�~�߹u���Vv�O��6��o2m�js�LeAJ���I�|�I�k!�*|�_j���l���u�!�m���,Ě���Ͽ����o�{�~&0��@�S�u4�1%@��E����H$�T+R~���`i�IRs긇�T�����f��%�>�I��P�S��c�
���	7�w�n��9���1�8�d�ѿ�MI �i?&�Hr��L�q�t���1���Y�T�m�Ϸa��O��~��+��9��k���1��f����	�6.����馰��Lz�2c�V��N��f�hbq�����f3op��8��o��O��>���6°Ϭ��>t���lD$!����}�w���?���:�a���o�'ɦy��*~a�hN��"��
��"�x���`�3��9K0]٨@�R�����@*U���c$��A	ah@ՆZ��P����!�H���u1�o{{k��z�Eڦ�&<Fu�n
���}@�yP.�K9��5�y��5��+o�
����e��JVx�Z���b@`V;��{8��4��� ?jC9�O���;�8��O^�yH�+�c�dT�2kb��Y=ʯ�,
�M����d���9�1:�hќ9E����U�U��ذ8ā�D^�mĢ�m��
�dmp�اu�ĵ'YwEX�C�㑑:���ꈾ�cvŘ��f�3��U}^/��,Ӛ�f5���Uf?;�j�d�Sn�� ��o���m����2������t���iQ�j@Q��YQ�_���0��U�����>��O�jB�V艏w$�7��7LN 1709�P&B�r�j���SW}�z��Խ�*� ��rǼ_�ކ�8	�ÂF�R�� �APK�F�4h����u���s5v�+aQ
I�0�dWH~����#x�B��
��9��W�1Y'`�Q���&R�
��*l�p�6	���J�b}K���MZQ*!�8;Wvz���!�k�B'��Z2V n���PLh��k*��H4GO%�FsO(#�^�77����1�͵]������R�UՒ���e�#=9.r�KAgph뭺���^��&���A9�Pa3�f;2� `L�"����2��.u]ܙ�+h+��>B�;}Ćuu�#�Y�9����!;4Q�����*�ɆΏ
}�[^j�M�UDqy�1ܥ�t<l ź�`C��5s��c�͝Egx�wMqq�yz5��;MLT�>��!�(]�(U�	l�,���Sԇ�Aj�%8�Z�l2�nK�k0� }���{���yܙ���_� ;�C�NQ�z=��*��9�3�F��'OOWG	A�b�2*�i�Ӄ4�M�}(�sR��F��+uu�I>�mV?DG�SZG8����m�E8����aM9�8e�N�2����e-nwi��V��Eg5B��T�G��WU`P��ds����{y�����;���U�,�55�Wx��뫖^���VSFڼ�^��<�u��F�4�/�'���C��אw'i�BV�k��(h��\jb�{ޏS���������T� 	�zaYŷF��9}��n��=��ã�+��/:�ӫhT����o���'�	�,��_}^���� 4j��x	���%��!�jv������|}���e��)#�mՆ,Tf�Y���N�<Of^�~��I	��	�qWR=�DY��b��5�Lt���(^^�4`�bYG�h��}�^�Iݫ1�G#�b�%�j'���9�+������G�;�g��"�N	٨��-�%�+�۷N��1}�L_u�rb��CZ9��jy��
r#	(����������\�:��g}�Y�d�Us#�\ѓ�U���	�h �GO�b�-�$�t�xAÆ���Z������_��u����AdU�
�b�1U�( �,TdQ"�G��Ϗ�O�������W��:�}�k�w̡��2��(*,	��R1�DWF,�0AE�̲�1C2�	R�4(|����"����D패& ����X�/E�Mvf_����_:pg�$ڳtB�����-l;%]�4�[�l���-ciMo��՛����S�`�@X%�D��V�2#_��_��D+��z��]u��K���{M����n�&m����z*��\�l��ua�MACs[Ь�M���d�~��<H�1�Ƃ{��ޯP)E����^Z������<��pz��]�f_���n�Y��0	A�`	)�����>�ޯz���ڰً��
���}�
�F��l>q���L���1`Z{"݋7Uޏ\Dz?u���⩌G:dt�]	���!Dz=p!�f�>�N����X%����T�QLǃ�m���n������e+!�zޮr�s��?z#�^�@��C-����ULV��7M���DP�R�у�V]��q�7]R���j֤��a�^����=�p{f��dD�����) `�E��X��:Vn
��Q�T����զ��U����%�\1ಽ���l�-�י6�Z�ُƞ ��ѷ�>�v�43yV�|�̤͘��sx�(�8p(�z�O�^
�A�ޑ֣�f�N��M�Dq')�5h��Xlǽn"=1a(�(U�f���t�{÷,�=������R~F��@ys��z�5Q}U�Qޗu�Uzʝk�z��^^z�7O��$%�|��$����fЀ5�&��$�.��n���3](�����!�}��Hd4�1��D;z��k��@r�/}U�R�:��r��5cxߎ�}�²��TdJ$��M��p&1���@� ��g%ic
��q7���ڋ��g�W�T~�{�U7#�s���Q(x�5|3_��tWmVv�KDؼ U!�~�'��V��W��@=H�e��ƇUGv�z#���)��Q��]�֎����Gؕ�8"@Y�ɴ�)���.��绝v�qА�� ��9X��=��l���k�<FhN|�o}�wvU�P�`�"�	�.Y���D�����f�1���19Ӱ���p�5�+W����l���{������D
¬��V��%��4]�Rш�hdtق�ve��%�$L/b�#8�	���	B���}�l�g�����tο{<�A �����o�EA���`�u4�"���&.湥}Kؕ�/X�ϬT,�UJ���7�0�y��F�񮵜�T����G�fz �ͩ��TT�B,00�80��2T(A27@f��WL��� �p�<���횤,(Hh�)����{����:|6�T�־�S\E��y����v{��Đ���Rc�����>���\e��@8	eA��EH�(`�\4C�Dz[-���
����3�dj���H�(T���:�B�jM�F�u��R���f�]�[.>�u����I>T�`1��_����f��<�zSÂ91�\�H x���@��*� IH:`)z�`QKR6�<�9tl"WJ�M
CCܭ��1���ld8o�qp� R0�M����qغG�nhD3��Wv��)&s[1j;�!��:��"B�[�Y5A#B��(0X�b�vo����ҩ5�.Ʒ6�F���G�B�S��S��̇�G,���Tf���=��A�<��{�ȩ|V���j�D��\��Ãq{�������q)^�QyM����񭳌��r����ٮ�4�2@�&�Ի/ڈ�#ǻ7^��1�1�xA�̶��:8����UN=��7]0#fF@--��3<�T�T��:��YGv84p�������@fܔ�WV���ͮq�JE���v�|����C�"<�< �+��	��Nq�v๳�L��N4�P��I����!�K�G��nހ���U\��Ǜ���X6 N�������]����Yʹ�����@�ZB�:GH��`�
βjy����\�J� ���V��U�^f�T����:ȔiJ̥�ĥȎ$��
%
��,��Jѳ-�	XLaL���DuHXj 2(0�53	F
d(HQ�*0H,r�#J�J��4�h�2���XPS#����9������8��F>�y$�,C�R��ĉ�J��9,Ŗ���u��͘㥲�W=��
�Y�rl�f�'����.b��]�����#�
�"=�E]Iޣ�n�#²}��Q!�H���6�]��{7��J���Մ�B&D��E
B���#ъ߽��2^�r��=Cs�,}J�xu�Ɯ?q��r�K����W]g�J�&T�b!wEcb�dA�2 t{�Dy؀tã6�f׽@Y)W���7��jǾ�����`W��c U��$x�U{ޡ�RP���6&/��We`q��D�rs�Ń"��7�X�ԛ�V%[�7bAFFw��%lB-��T�*J�x�;',�$(\�FQ~�{��z"#Q����֥���,��ˣ��L�����t5���d��V9�*�c�W�I����>�Z\���0q�۵!.��^��O�+�RZ5X�u�i!{;!nZ�lڌS�]i�g*�,��"@Jԩ��n���,P`��*#yu*}���L�Z�-!د�"�`V`u3=�cJQ�k7�5��L��No���n�9Lph:"�B��o�
���ǝ�W*�P V��Mi���0��t"6���}��ؙJ�[t�e�K]�]�S���Zb�v�]����E�39���v�j�XrH�`���dA�A��K��C�����f���
�.���;���������򻫔z�#V�e	.֌4]
"�&+�\f7�I"|{�y�;��\��*^<r�]����߷������ЛID$����SVR�["��	r���g6l��u"u�=Ϸ����HVOZn0��m����Ɏ��s���[�w�h�,o=�f�𞧴g����R?4�J���E���@��%���n�*��q؃�W�f~���N$�/{ə��1�j��'�ڲ,�c,���A`6�9�d�N��&���w�I]��֥�Ҧ�'�tk���s�R P���]_-���)�#U���!V.�r�i�����B�T�k�N4��1�#x�g6^Nݭ����w�tk>��l�빃��f�ك
�>[#����7��{��bQWj\�}���`)W]��+t�[�{���ԟ_m�e���h�R�
FŇ��a)�}�E�^�B���I=�Q:��6�i�#;�n,:Iu,޶�[�m�C�(qӦ�G.m �<�ׄ�ܶ�ɮB��dJ��������Ҷ�����-�;;�
�-��Ҭ;�UJ�K��cv2�hSGl�<{2�AS��馌'TTu���Jmf潺��a-Ɏ~���4��{��t���r\�`%�;��dΎ��/q�S{P�3w��۩�U���<��(�3��eL7Y������6��S��+r�(��`�U���Ry����{���{�=٫��R���tV:�D=��J$��;��Q����\�����u>AK�wұ�yo!���	��V:u�dB�\�H��a�ρ�B��o�[	��K�/���{^�K���{*d��A>NS05��Ƣ�~��IX�t}�Vu��Cn98Э���Q̡���-'g���Ej���v�Z�Q�;�3�wb��L�ՠd�\|s�s�tu��c$���������/�M�n< ��"�o�| Foe�-��v�Ka kK�s��+2�7ܚ��sw��s\j�u8'<e�J�����o�W�����"��r�h�c�Z5�� �oQ�C�����>�b�q�JXZ�٤c�着�z���G���#���Ѓ��,���\Ӣ#Y�9�`6-�MT[ V�X�B�ӓO{jmՍ�V�����^�����d!,4l��#�xJ*���$,���]����U��Р�'�T@d1�X��2��:E�����乾*���v��Ӗ��/v��.���Y�g�����gX1�]��mq1�덻���7��F>�3l�R���޾;Í����D{#�J���������}S��Vc���FҟwO�#dO�Uz�\U�{��^�������ު�o�ީ�~_A������-S�?z�a�Q��n�������hո�LÛ�B�K��FR�)�ǋ���F)�A��ӓ�W ��1f0�5�� ��I
�G�	���Z���|�i6b�-�^��񯾔���3{0��[�Sѭ�YY����j��J�V+Q�Q�DDs��<!�^�z�|$�[�ti��Y�A�i���}�^��+���ũ�qeb�CMAڕ�7�qǣ���tx%x��HJ�ى'��mb6V*bbaK�1U��"�)Pb�C�(c��tZ��m,F��U�"�X��U\em�Ud��*�TQSZ�V���)���X%��fi��6Ikv�n�Ӽ׏, �����J�;"�ۭVη�z�l�;0�dK���>5�Wp�*�5W��.��b�|��6�o��p˅�SQu���r�;��;e�׆��������Tl�I��v�\�{X�}��qFj�w&:鴜�P��Σ%��r#��g��5�TG@��}�z����~�R�����^�VqVLa�\߂���Hr���.r7�FQ��Ӛ-u��#Ћ�Dy;��Vަw8ؒ@wu��5ܹҀ�3Mt�Z�����T��ԛ4u�30v*��_U?]�݂0�1�X@XEX�u����0$?�6��ɫ�����ųGLgP��Yy#2���Q��!��=�ۚ��0�{�`z��Ur�|�k�S_R���1�g�͔����6�M�)���b�Q����������O�
#��e����+*QY���eMJ��M�8�aĸ��%����6�+��}b�h��{��[k�"��b�,)��[���v����M�ޯz����GѶ�`�Yo��9D��1�,�Y�)X�<��v�ط��b��^��aZ���}U^��=�*��AJ=����].R�0g�;�}�	�}g�������T#GW���#�G�#[�k���%����k]�vU��N��+1�²\3 Q�r��H+�ԯ�ꎛ/���(���t��2"�I�-����L��ˁ��x[s$�	3�M�{v���Rz��Rڇ��"۱-ŉ�L��ު�W�|$IK�\Z��`|{�X���=Թ���Fsgv��=6K�;n�Uz�H���djfuu�mw���N1�E=�v7co�[�w%v,���fLj	F����@D�Ȧ��s *J2�.\d�M��h�T��
�3�	a#�e���YT;�V�����R|��7�,ћ��K\\e��O�r:�vu��͞Y��M0)��n�uA�	&��NQ٭�SJ:�����F��ov�����~��; �a=6��-uC��n��-�O.�m��E[����v����O~��o��� ؕ��d�����z-�=M���������Ì7#����\��e��{q�o���}����#o��T�⧌/���w��e�J-wbޱ�!^���EQٵ2���G�L��\�´�7�k�輕Y�� ������Ew��Z�(���N��q�fY����EoŘ�7UU�ys�2R��^�[�a���-6��J��ܯ*�Z�+�!��%[ۭ)9|�V�	�KU�g����>�q�ߵ��2�S� (�-2��V�Z0QH6��bʤ�l�-JA@-��������"R2�UTT��`QP�,-b�Q������62�R ��h�
R1dnR���}�$�д4%��^!9�+{����5^n�qJkh ���r(쑓^J�R�h�A{�D|���Bs7�XK���6���u��5��i��S�x�S$�0/E��:�������]w���]�i63��MX:�n��T��2 ����:r'�I�΃g9�u�{�j�L'uҽU^��{�DHN(&�F�ź�ַ���wZ#p��S�����_gr�$U����2����ޅ���e}L��u�o�;8<���^��g|��V��	%�Ĕ?W��﫸{���Y_Sn����M�-��]ƮV�p8ݼ\�nl7�t�1�ϏQٗ�:����Q��z<��e ��#�[���vn\�z6�;b]�m����=��[��V,�`֕�b�2E/~���7������W���k�m�l����jKЭ��</�Z�*��ǲj���u#:
�9N5q�;RP����[}�2�z�����뢽^s�����_Va�ў�إ[�p�'MRW.[(\�qʒ]d����UUi�QY�"�=�����s�{�(s��&O.��ۭ�ϓ�ff9�42���e�ۮ�H��{_�ޞ��|��E��TDV%��Cs��_U��CdY��3H�[����c	��[X��S�NY|�S%���Tμ�����z�=�z�9�������lVێ�.�J�IW���|��E�l�G��.EZey�>�պ��w��@~�x^S��eB{cO��{ِ�t�A:	v.8�/����7!�a��:8yd+O.�X謬#p5.��QϽ�Χv���J��`.�<O�DF�Ee���^��=�2dC`�=��BuIL��۩ST�v�r�n�&2��q���g�ܭ�uU�n�����U̻ùnk"V��-�=��G0�4mI�ԥ"�ח�CMZ�ۺ�P}Ϸ�wn��{=�kY��
(+#$A@X�����	�n�p4W��D�R�	�W^�R��z��Zq��f=��E�^�}^�z�w���-�/���Z���'8��.k�o=XOS�&�ʸ`�VU��%@���.��/��S��W��C��E�{�3_(�[�MR��8q�'�:e��3���.g4��ڬ'�41D"�<}�=�ljk2���)m��K�!��I�Ã����e���.�PS�]��.��ŝh2���`U!������������_D*e�-4�speJP��l�V����I�76��޺w��|������i1�G+mj_����Dq��YT�! G��;:���*͞[9r'���:���B�����J΁��Ҳ�a�h�yk8���Rr�ܨeq��b����bF.��TN��QV���+ ��=�PٓpG�!%��MJ}^����_W���U�~��N���r�A�o	z��铢=�M�<�xo�nf��n��g6ܼۂQ�{�[��z�o��Ϻ���k��;��ql�����KgL�^o2i�U��*o���Z�A�x8��.�k�#��G����T�L..&>�x��Ħ/k��K_��C];%2�v^5�r�Ug�:�Ë���{�0D�s�<���ǩ�a����N6�3's�+'ϗ�w�*33��	���9�z����}OVU��[r>����H�@Ё��{������=�!�`1X����D�P��<�rs�u�d��a�s,̛[�t��gW�k����#vwK=\��T^X�
�2�ƈ�����>�X��17��]x7vQȃٍ�:�N�<�qs�(ml%�u}�'D�l:UI��z�K��Æ��+d��m��7S/Ȑ��%"�!�]Jmcm�%��UU��z��ӛe^�2�g���)}׷��L}�K[w�\{O)��մ��������a��X�9�u�?�{�"�Q�+��#�zX�(��.+�8�5d�e9�f�싹��Y�z����z��k/T
w"�gO�@Q��AV;�/Q$�������Ivv>�L��C�}˧:k��.�l�P�D�z�H��{w�F�L�xzi�0ۃ��p= �;�.]������V�?�U_L_n|�����=�Z�q00�cH�Ym2U���6E*�
�1��B�Xb0bJDF%��HU`Ġ��Ʋ�2�3F�w7�9���5v�5�'����@K�d`!]�5�b��rh��dC��>�l�md&�K�i;T�l�:���%������Z�E�}<�J,D�8dS��@��J[�����`�EbK��T�OE�~�t�.U��a��źUm��V�ڜ�1ۚ4�&1Q�ޡw�k���+p�"%z;���/�.��P�.;(/y@�]�>s_<�.w8�r1o=�+`T�^�˞^���ŭ����
��y��ddy����h���༭��l��Z7h���^�-5�{ޏ)N"#��֜N>Ӹ/��d6�ݨ�e�e���&����˙�ǋ�Z�J�O8`���r ����x�  �9�4�{;��B�VWZ)��X�m��O<b]�5�ݮ\y�}S�{��3
7w����uş,e����8�\j��k��i!_B*����$@�eaU)ZW�7Ys��M���Z�c����s&������c�ͅ�m=t�M�����h���7�����{䀫Ṃb
��6�]UԬ4�V�9�tem�[�� �W���u��Y�P�ɡu�ਣ;l]Ya-+F��*�FVw�٨)���M#ӌ4֫�V����Tq:` *Av6�V�2�³9�u�;KF��{B��LK������\h�h#�K=��|��&\WΓ
�R:�"��9�}�M�7ۖ��k�E��_}ͺ�Ӿ�*J��Q���K�N_h�#ts$P73Zl	W-�36{��e ��7ir�9����p_O]\��M>�i*6����r9i�N�o|Ӷ�;�=�����0�Kj!�����0��w�W�uo
I�u�˳�i�-o{�դ��]�8E|v�⑻�(�aM!�ʯV�]U���k:���]Kn��z�(���u�̺��(F1�U.f�x����:�������C��nc=V��]Y~�O[F���[�6���UU�Bn,�Ş���D�c1t����p���k��7�>9г�܋�k�x3�tG���� �k+-����of�jqݟ����?!�k�(���;�>,^��"��j�FL(��=�����n���0�o��9�w����n��YON %��7��u�5K`d"�D�������H
1�C����-Y����w+��]v�mZ7. ���@1�u�S:�*�r�A�Z��0=��םЈ3�����e�kѦb��]���y��|#&�e��+�׀�Ө5��q}}�`T���!݋N�%9P��üg\�Ƅ�hޝ�g�h[W���y�Y��o,q��Loe�Z6olmr���B��z[��ښ33��a��w*�W*��*�s{ qJ�Z�6��ܠ�zR���iEˣ�" ���E��,�J�Q�l:�ջ�#�Ӥ���X�V(���o��%K"91��݌���b�5�:^;���� ���ei�]���9S�ˮ�.�*9�2�e��:ď\��|�Hb���o���5�v�6��u�vM�)Z�9�u���N��b�M �vzG���/��uϛw�;Zle��]�6F�4��>�]���_am���z��c���]�r2�^���z'�#�⾚.+ɕ�D��"h}D7}o�tq����Xn��_k����<�6�_K��<�<ʆ�v�Ԯ��S4�4jG�P�N�v=�����/�f�B�EQ���Ö��2��J���3��Ꮠzvu����?��F�C}M���/��l���=\�h�^ڏ&v�r�f��q{���G��=~��>�y�v��ߧAQ���OY�W��i��c?�PKhc]�h�q(�k*=�]_^L� �Ύ��^J�8�
U�7h��y��G��\G���H�Z��Y���Z���4^*�[���ΖK^2@��_i��y�ЅIQ�/{y�Ɠù�^�����1W*�N�ϱ�]�CJj����E�	/�=�R��3j��X�	鈈��	wA[+�����[h��8G�}�ow[�"��9˓5A(T
QR��隌��m+��F�Q�ژ���Z�B�Ǣ6��{�l��9pp���y��~���^���Ղ����F�1kE��YP�32�P�s�� è���8�*����"w��־��PS���v��w�t��+.ŷ�.��Β�ا*qk	ʎLێ��0C�s`!Lԭ��K2�Mيʷ��O��c��G�5�]��ܣ	�m�2����I��Nts�n�NrO���+x����+�W��}U����k�>�h�h��&��O�vu��M�<a]�]�w����}�ꕑL�D������N#�~�{���\�q�%��'�fn��aQ�樭H�)�q�$W�ӎ��V�$
�y�{��Jh�(}�����i�9�p�cF8��z]�����!�r�	�!!8�{uǢX�i�2��ۻv͙�ήZJ��3�ѵ��er�	�ج�+Wq�%;=�{�o�ｯ|泙�@�0�b �M�����yO�m$P�"��������3�������z�|�(	7�I(Z�o��T,ܸW;Z�f���7㯍�{#�\i�J�[y�G*��S~XK(ዤ������QZy�L仵=+����=��W� �dw���TUz�ޥ�z/��_d�͘�0���բg1k�.�B	�T�:�$�ܨ�5�; �`ۈ�:Ėe�gL�����&{p��(d��w��k���N�ԗk���B�lD^F�+\�K���ݢv��V��Z)�j�>���I�����lum1I����ِ�nµ{�cdV{��q�R�'����M�Ef["��4��8�J76�5��k������.�B��Ӝ�
Y�P���"(��������JI��[�Og� P �f�|����:[��TR`�_���U]]�	$��R�RLHe,�e����5���3
�Loϻ{ϵ}s��er͙Qa줷Î��� v�z'U\���wtm��k�^Ñؗ!��pN�(ॽ-����e����-眸�x��G�m�N,>��Ǭouu!�������8T��R�6�E��*����ZPɅ���{��Wa_{ԛ�A��O+2��v^��-}���I�4%`� �w���z�R�G��UM���^�P����2���FZ�M�H�9U�l�+�)�$�3���Klδd���]fv��duF��D�~=\5�͊���OI)��<5�;��]�����t�i��؉�gj��5!3d?Q���BE��b�����/3�F��Ӿ����o�:��mTq��#�Ir��O>�;�UC��d��)����8R��#��IoHn�7���ƻ{ߧ�d|�S��� ��A5�!e0�1�X�*,�Y �sd&2�T`�j���FB�0ɒ�.44d��|�4��I�jo}fܰ��nif�pὥ��5a��/QAۭ���E�M�v���H=�;���|�rS���0��ǐH*�w*�_�6V�'jL���Fgg��u��η i��k�ꪠ���R}t��vx�O��+���)�;�q���i�����;�7���IfK���=j�v�;B}.��L��|��<b��V����Rt��!�6[�v5�&G$�=b�C��:�G��RA�EB��[����	�PB��)�]s��ɃꪗY�f�b�ÒQ]�X8�_��@Vַ�ܱ?�)�O:E�(l�ޒ�٣e�)#�J�L4�M����� �y�oH���J�����U>��.��k��K�Μ��zQ39�W
��t�¹������(h�mH���_{ޝ%(6ꮩ�F "��"�(�+�]�кqֲ���{���=�Qt)vwWS��gB�km\j�5�<l�se������[kg_1���w}���d=��5o"NtI:&tI�u�f�h����y0�9
��/F12��*�O�ՠ"�3%d��̽r^�L�o�z�����Q���C���!�j<#2�ٍݥw�L9&9�Ɇ�w�^�Uo�N��v�r���ު�>בgۦJ�m�ѳ!�rb��8���`�=�.���Et��#s���g纙�N��-�����=�=�@`E�A`��ߜ���<�ܧ�wx��]1�Jݬ&1���j�\q�Ҍ�n�� ���9���pr*7l��?G��jm��7�-V�ݵR�0�虫\!!���� �WjNC�;jῪ�UIE���U]Γ���Tb��t����Oa�9'�C-eh� (U"J��OFk :5��<���W^4b�i�.�wI��]i��)�&�ŏz1fH3&u.ȫ�m�ͺ1p��F��L"��@2r@.�p�﫹nZ��=��샶�ީ���sv��t�dz#�U�j2KA�S��&����f�]8m͵��z�����("�5H#��{�W�UYM�g����0�[�.��gp��q1����ɍ)4��n��3׳]NZ�L\��/�=�R$se�Ͼ\�fV�x�Q�v��Q�vv��4�-d��!(Q��b��oތ��7����Y��q�|���d9{�K�El�0��.ӵ�}��% z�8�~��"9S�>��;�+��U4B�{c��R��J��{�;�3���]��t���@%8,�u���$��v�������R�H�,b�y����S����f�	K�Wn	Jp��Ns�Z^�9��ۨ�r��v��*z@*u����E��ΦE᛬Ծ�]$q`�j��1py��\�ԭ�e5r�A��pߤ�P�ު���2��+2��S���6*);��\���
WiW6PМ�#�Rs��=?	$PE����_w�����ϼ�؜/0��y=��8�\��e��v�s9�KШ^�8�n����}���z:�����vT�T�P������k�9 ���D놦[.1st�kv�{�p�n{��DgA���O��W���3�42>7��d����)���R��^ ^s�j�R�����C�z�A���^Ɗ�%oz����{چ�Ÿ�2�R�����	_x�>;�b&߬��cmiUQ%�r��s-$�l�IT1%1EZ�h�AU-2�s������e��2]%(M&��T��F5��|���c��|�+���@�eɦބz�A�	ٻ��=X�/Yj���합.�K.=苷�CR��b���g8�m2������ǧ������Q
A�������x�ٕ��}5��dO�>�߀Yj*t^��<�n��޶8s/�ذw����������s�a�IلBUU�E��X3�#X)Lӿ�#Oy�Wԧ {5�I����{]�p��h5"�LT�:�3�V��"��5����g�zokn�����Ys�"�]Őz�U}�*_��1���Ҥ���:�A����=z͇�u&b��e�쌦�Ѧ*�xU&�fP��|�߂c���{�n�=��ze�|��_>���YsD�~
H_� h'�x�d'���\\�U��Q�v�$����ty�(�����4�U9~�{�ܨt�������fGN�i�q�/vk6xn�u$�ظ{ǼM���;�x��W
�
�b�-�ĕ	�V��
��'�gX����n�NOOl5�n��˺z{�z��b�h�� v��708G&E�S/����LGOm�NH%Y�Ɉ���pw���Z�xc��4_��yv��9�?w3n�H������4�V�3U��{��%X̞������\�B{���T��"à.��۾ٵ]&wS��X���K�J�m�gl�ф���Ͻ�F��@B��I��D��'z#�W+�T���k���"\�K1��ݙն���3��i�wR琣z����P3ވ��{��&��������~�����휢�ʵ��3zrw�X����l���&�eB�}�8=�b�|�T���kѹ�Mfab��e��e��������Jg��s/����ݗ�"�{�z���&ʃxOU��Tiu�yCq�d���be�}3��?����igo�C�2r;U1��	ӳB�{
���hZਸ਼�q0�<���P�S�wzE���+�)}�z���|���}��/���f��hf�E}�Xt��L�G�5|n�o��$S�Ճ�(�]_�phr����N�"h��2�(ح���V2�:����U
v4T7t��k��s0��5�5�P��З���tE
��}o��lV���A^:{v|�_^�(,m.��1�:�WW
�˙�`�G)�QB�iϳI��X-J��ri��[�[ۆ�_�:����+��VCY�E{��K�>-�ڱՌ�y�$; ���Y���}�]�*�^�B�1�}��iUR/>���h�k,�(�Ac�U��k{�P̀��k�c�\
�5��l]�	0�0K����n*H+"�a�F�bg�vR�-
��wF�r��"�G]�pi��v�������5�1R��Ɏ���wg��0�k�6�]K��j��1�9�?co�teiuBx��ޮ u^:AI��X�zS�Fu����L��}�l���6�㚙��ξ޽���۽���,2*!���B�`��f^u�ќ�>����VFyS��*\��3���_���a>��(U� �ou�5;j
�J��紆�d���6�΍��w#�-*�>[݁dQ�ȗw>�P����<{���Vp�wݹ�s[�/��Iu����I}����Mh\�ϧ�7˥Y2��E`]�kh�pGK������ͷ����Znj!�t��(Н�ͤ��.�p��c���0̃a;�U�#��î�rs�3|��R��v�,Ћ�.�H�s�-w�Dh���O�0��{ݒ���ް����XSS;Yr�K�,�r�b��P��j�j�B�C��]����.��Q\ږ�4]�ŀ>����U�����Ǵ�3��Y[/��OqZU�X"��؊�;�[n�F[��D��/p���Ϋ4$N��<���P��0[�A���Y.�x�dQ�7�k:�x#cvJ��3�2ɥ��$��]��6]o#Æ�d�-�w�4�;���$j�N��1�m%µP&q�N����|4���o���G�0�;e��
��x��QԦ���j��X�l�[��f�|,��%�EF&̴Ì"-�"�v�B�pfܛ�t䩹�YU%J�cn�s�ɫ�U�eӾ��@R[(��>�$�ӆ�^V*���胻(��U�Wm,��اM1yv9�w��v�sFޡF�i6b���<�p��s%2�x��+W�8j�ܔİ9�޾�ґ�&}�}���m�R�!�%1�;���Nu#�Ӣ��= ���
��2�����Q��f�9Ѯ\M.�/rN}5J�Jt��{ok{q�ӝ�K��@'ޕ�,��6
C�Q���\#�Ga�!Q"�hf���p	V`Hmc��c�Uj��5�\�!�X���f�@>��]��3�]AU��*�A�c�s���P	�!D����B�"�H�EA������Y�����?��̃k��jH��")���,.�0�r[Ze>��z�)r�EbU�{w�]KZ�ޖ��3=��Dz �z=��FI�?��XN����������8#}>�r5���z�H�r_H¸�s`�>�Jk��W��T{���.o����Z�]�ņ����;��=�h5���Ju�IV�Pcaoܩw2�-��2��41��
�;��pw;#`���=�ퟧ>n+:ݱ.���.�Q������u:����i��dO&�h���;����|߯���́���#�< @���:�����s�J�1�OJغij�p�;ıY��h��%s��և@	X�Yi���8���@��XJ������������ս��dr^HoR�0U��p���9v'u:�ꄫ��s[�TS��Ƽզwec���@;WA�L��yƸ�d|�v,�]��P��¨}����=W���^\�Ory��T`s`s�z1��.�(KEp��8yK%�A�~n��G�6g5���%�S��6��H�~��>#��D��&6�N�"��Q'����D�"��� ix���>�ͧ4Kh03%�6zz~��DG��#$�u��@jߎ�l�~fxEr��^��gJw��#���GO2Ck��n�8��e���u#�J���苏�޺�r������GJS�v�W|�1$da$����� ^��q��ٴ�����U�����l�%Α�,��Ut{��Dc�`G�?�;�]��9:^�=����n��P*wb �;\��W���(����G���w[yw]�\������?<���Pq�T�����]Pn��j�'H
bJ��IX[@� ,k
`�ι�w���ӝ��6�]u��m��xR	ER�
�P���S����5��	P(0��*vL���ȸ$�*d���ܳ��)b�]��^�ӱ�@�}DK{q-�p�S[��M`m��j��Y�%�]��*���No_����PO]���]�!��3��儮���2��/��.�.�:6��J{Tھ���[�%�^|դ	'f��W/�F��� .��>����R��{�rʩlj��P,��ՏI����w��h�贚F��4��0����0���K�Ht��g2���zw�'�:�d��$������T�JO�Ok��N��b����**IY7�hb���4�T�q{����� ��؏��� �� �_s����������w��/��֛��J�p�;]It76Q'�jʪL�fd:��.�#3F�cm�;VtZC,8������Eg��>�>. û΄�����y\>+�d)&?Y���:Si�j��_�� 8���AO���
g�z5ְu�@�D��P ����� Ȃ$ ���*� �j���n����*���3�;5/��������;����b�=}+gwUʇ]an'�>yVl7�1�F��bV/y�y���K���sCs�U�Z8�p_ڭ���(�≪���`����s9�3}$�G��LB$���՚�n�>�h�n�����&d K=�1����w�ǐ��"e��V6�q�FV�Y���O���NNDM��z"=c5VL�wn�ėQ���/W��ވ��ژ��޶�������Y�KF�
|���,̩Z��(/nh���6;Hgc)	ö��'��+n�w�)� =3D&G�����l���Gц�}��f0�ʰ�m �bn<.��;�9g�T�s�!�����*�1q�Qu�Oj�S�輌�Jw���y���Mn;�7u�Uܛ�a\�2�̃�c���z��C��{�AC=O�z�7p�xdT��{ޏ}��̤.��q�g������N{��s�
y��Z��Z��n�S[2��0��z6DT�@'���0�� �,�0�1��*�����?
�}Qп-����ok&:ɽr�u��/��-����r�,�;��Z�q���B�d�yt{���n�U�:�'T��S��T��|wo�~���9���浯�����E&�OĂi��crC�x7��lV*��1�Y��i�V�08���%3pc�s<�ő�771��b󤢖��G��#�0�g�t��~$��@�Ds�GU���v�Zxj�����G�m�*P�J�BCU@Ѿ��wK����߿� �
��(DI��;��_{�C�'[���F�H
��'V��y"w��D>��5R{��L����s�]S��������G��{���`di�Qc��(��>�.�Y����Z�,8'�[|���3�r˪�Iu5�<F����G�U�Lz�������g~�}yv9P���˺q]���4U�E��輾��,�
�lcgj���O��jF�G��Wf�W��\��>�6c�?0P�!
�+�)kw��9�﹬���lA(퀓�٪���^���gG�T6���4ZJ�<[̾��#}�/���.D`̆�%�jL�Ŏ�1�~j�RQalIl��ڔ���B�2�Pvho;������Y\��p.�!�����������s�뿉��v���x�vU·'A��[�pl��7@vG���R |>dE�"-�A�����Y�8{��C�hn�_�To���s
[#|	u���F��G`0�d�v�c��X�q㭜�2��zd��ߪ�@���ߕ)_{�^�؊����j3�(�}C8+� N�+ܓ�����'��ɀ��ԫ�].��,ŨS��{'��;��+I���o�����o_4�� �b�̻sTa�8�Lu���9��q����Q���6�ӳҾ�ނ�����x�����×LdGS=C�fÛ=��.*ݑ*t�V����@MTGM��/s����׽_������Z�,#)Ad$� �"!4�1�+��k͑Õe�>��!�K����7(YpK�EoY@DE.��Ƕ��nm]5w�ͽ��l��tc����+e�w]Q�E᝱S�}
n�~�|�c����t�R�
�FԠ�H�:��<��W$�tu9�j�{wK!�+�&v`5^a��묧�~'�"�"�Po��߷c"b��Z���%�ݘν��t(%%�%=�r���4V;������錣Q�pxb��]�����왆�r^e~�T�y�]z2~��Oǵw����Y�gj�=�*���AS��������_�vv[���C�k;�Q{ޯ��h������.�v^Q���d���ҽ�
����|s領�6L�r]�y59|����ջ�kn�C����P�Ӄ9�l��]:��z"ži��b��\�&R�"X��E?�/{����K�2:��=9\GĊd-��)���UYZ��XДe�����ZɃ�It=舿�)����>�*���=&���%(s"��̋�7N{��c0��x���C���x�~#�C�ѕ���**Ы��y�9=�J�5��t�Ŭ�gA�����z�t��2KO�l�΍�Ji�����87��[�A�~$��U��.��R*K��Z5q�����}�xシ&~<3"��}t��[V�tP;nx��N��U)wh��T �8M����a��ޏ6�\����`����L����H�=���@B�k�0��8�p�D��ר�bc�>��|�� 8 ���2;�Aؓ�X������DG��wނ�9�,Cp�c�ĭ�k��r�{�I�ߝT9U�N�4�N\k%�W{��89VD��S���ۭʯ���P�_�7�O�0sﾫXv���Npd�П��g�J��aDKA��۶�O(֐�ET����N��}/^���U6�UB��a%b}^�\���{�^�޹��r_�y�Z
��0�KݹÝ��ofX�}�@���6S���{���0C���W�_
 W��>p�'��:%9 .�"}�<#�m�HA#�0�	 +�!id�*H�2��P	#IE�H+lK{�����Y�k8�dս�{�q����^�.)��4S��w��G}��aӁ�Y��[R��A��!ք{��ط4u=ӷ��UY�m�1[0��*#�0
�8u��/c����}k��z#�
���I�m3� ��&�@?{�O?�4�S������4,W)��#jq;%�P�Tfב��7) 6�  }��Y���3��y6;���:�M,�r/����l��d��>�uC�S-F��\)cKN�B[=rs<�g=|l�Q���p��a�fy]�E���M�u�{_¾�G��s�������<b�SX3h���"J8�����zn~�rˉ�+gOPp�<���㯥@�M��ޏy�XR �?O�T&c�	q=,��J�����%�B8��#g���o4+�=@P�=<���$� om6�z��o�A�q_h{X��<x=?v�տh(�{�}R�VX��|�Wj���>Τ�s���[�9���Q�&eVJ4%�>�Y���O91�ה��$��F�&|���Y�s2`��� �@h%[�ܱi�I��(������䕴�q}CrE(��Em� �����C�C��C��1o����U��ԫV��إ������#(�$�Q�g�N�劺j�V�zk����W�Еn���B�蓿�~�_��:�5i�H~�{�_k�v���.�-����K��y�u�Iw��yҜFi��&D}k*�R�?��U,��y�3Nl���CE���.���,�d�*�c�U�L'7!\�K����1�0�z�[6���/�sj-I{��(f���{���8�˷b�>*��Ɍ@��A�?|���12���X��;�U��{���G3�Q�U���yv��~�(H
���J��?��2��u��>�K&3��^�%vM����0H�w���J�BQ��a��|U}���-_.{Lr��{��E�&%|k��������ģ^$����󩫔��g���X�o�#U��O��DK�� �7gm`u����!��{ ��q�9}�xq;�x��K�g�h�j�}���^��^���(  �P@�,�$�xUY�X.�<������(�[�wuڢ���U�f��:�o����0��f�h��ۣ��"'y����*։Nw��}U-��]T�Z8��[DG-ɐPx�LMT�������o)��oV\KAK�&�:-V%Yv~Š���+����;n��HU�NS�5�ƪ��}p�=J���UsѕF�aTD"�ņ��m���}�����uĉ����W�WS��������0������=�5�,������֋�Fpփ"*.������y��R�\5tQF�Az�U{�e��r"k.�ẹ��Z������3y�*o7LN������I%f�'�w���*r�6��e�ܯa�>���dΞv������"���* ���>�b�DT�Ep�ɕ�۪� qQ�tr�L##�5x�R��pQ�>}��3y�����=�.���X�J�Wp��W�o��<=f�]���Ҿ�M�7��U�s2n����z��W0楒GS~^m��C�p]������g˱N��z�3O,g
����n�PG�Щ���7�V�(R[�rn��� �o��M��t��<5���̴���YÔ���;.dkTi�N�jZ���]���_�eG�ł�N!���l졽q�P��v���l�LHql'_>�gH��i��i%W^s�;k�����rv��רY��8b�%m�������:�k��dr֜�׋�P�XK�,鄚�Ć=̡8FSzwV[���ΓvBBO�;6���d�!%��)���|�e�/:�ĝc���j�Ct���^Mu�S�:���	�ʋO!�P�V�����۷�ߙ'7,��B:q9x�%���ؠVo�Lp��g E�*�C�ri�u�EY�����t��*�$Z�MNs]+-�m%T�U�RΖs^!�E�����K���c��6�؜�\֊kD���fы�t���!F�����P��6�V^����uq��ܡ2^u	�aU�A��Sr*Е��0&trvީ)�����t����Y]Vi�2�D�� �*�Q����Ț
�6�yGn(w��n+�X0���f��AG%5�a�4���ʕx���ֆ�e��l٤
+4���R{VfY�GV�ܓ"9�l�d�"�J�ܹ�hj����غbm�ꀝ��(2!���=ǘ���2�f��i���5����Ŭ����0,��GsU;���}���+������^
H��C6�mVN�)�\��*�H����;}�8���ҥ�1��A�%B͋۵Cnf���u�v�]�[sڬ�2b��(���� ��<�bOm1;�VJx<r8��@m*���ȡ>�F��v�S���\�΀� 7U�f�w��ɝ^"���"Y���S�q���T'M�� j�B.X��g��}��M?�ė9�����J��1-�ٴ0�N��� �
��EK"AA�vi�;�^(�����ɹ��v�@�7d�9�t�}꠲fS�5%uԃ�;�]�:�{Cdp�o��Яz�Eræ�R�R7T��M���r�����"�j�؜���Dz5����Ǳ�^���������M ��3����*W8$kW�n^������7u�6��-�c���?V�<���g������^���w�;�DI_��Z��ݦb&�Z�w���s)�M������\Gl�=����f�����׽�n�ÿ��w�6>��Kf�.5B�i X�"2O��C�Y�}�'q#�j{o�9Ef�F�r;�Y�w@y�eg���p)Ǐ��T��/y�l��ɨ3��,6y����çWbwC��-ɘ�<7�hqY�U0��Gv��5ǩ��t�\�aa��u�V)� ��% �U�pf���}�Dv��8���4C�G��y[��ʄ�`O�򪳣�ӴXp܃���G8v��ƴ��\�>�Q�$mý"�*uE�芡��U����F?�Y,��pv�G(v��K9�z<ܙ�e�.������(�VT�
讦&ئX�@���q[U�]��R��G����z ����`G�櫕���v���{	��sr���5��cQ�9=��&�Cq"5m&i��{������#-}��O�;ԭ ��\99ƺ�%��jd� ��0@�u!�[r1f$�l��\��t-�T�ۥ�Wm���	�U|d������韴���t�Q��PtNjZmR	�ց.H��|Jo,
t����TV8��`Ɍ(� �e2�*�Ž��߷����/)��<�Gp]d�6f�z��Nܾ|�pugt&���bK�:e���tNC\n9o\�q�-�5�d�����f��R��b��*��#�m�s��_�q�X�UÁ�CR�����+o.X�*b뽼}V���#��#�eC���؋���Mc�.�2Z b��= z]���s-����g*Vv|2vV�iʢ�8�4��UqZL"�$��S"�S7��s���D��(�߽c��y�>����N'\�Bqĉxxv��u����MB[뾮��=9�@�eܥc��\�9)2j���?zm�����$۹�9B�M�m�A�
���UqڙL\c�Ld��B�)�w �:��V�G%�f*}X�p�f�������G���u?}25�2`��$V��)�̯]�ޯvZ^80��C�B8T�4�.X �T�o�x���^�V��l�G:#����p����l����^�{3�����ȑ�u�  
Af�ڡhcfb��AJ������aK���H��Q�e�2���6T�g��E�T��,ݦ}���VV���L�쭻����r�5��3BÖ譧a9�x��x����3u����V;��2��@���[�gc�'�Zo��whvL �G(sv �ሎ:���J��:m�d�TP�{�;w��@	[��3׳���>�_O	-�b���T*��X�GId�{3yש��Ay�w��0�=�=��wN��z#���Aag�Or��K$�!��B!���v�����Xցn+�l�&<��3O3Y��%�E *JW�L�ߢ"q��������!�v����*���<�  �mR�t��I@��VYrWTZn�S-���'����$o\�̶&w}�DL�޷N��3c��/&G��/�����L��L����'���� ��b�R������k��/\	��S��M-�o���RS��c<�����m����qս�_�
͠�Ų��PJ�h�Fڦ �΀�֓�����ѢPbZkȈ���ȱd"�����j�Ҝ�KU�es�W�(Z3����K�؊�ЗZ�N���!ȱ�ɛ� �{����G�V�ee-Ǉ� �c]H��r;mF��i�ң�sA��6a��ň:��FC����)=w �ƥ�ط �?#m>�]�Xrr{f�a�UQ�?x�Z��ӗB�G���f���lFwtc2	Pٓ�_���O	��f���R:d�	�a��T��v\��M��
�:��}쿾*jS�7��2.��H�E���6���E��@��R���*�8壮�`i�a�9�}��1<λQ��Y.S&Fʏ�~��މ�A�~�6������x2;�5˗s��tg��z�n(t8���YS�V�)�K��msO:^ν�oh����AL"5�(����S��,�q�0�b�z[W��6j_Z�����I��.��h�D��������w�HʵŬ���rC�9�XX|���J(6O9�%IA�"�>���� x�  D A o1Y�VϬ��fk�.�oz�{�St��&�'{i��Q]Ļ����c�6v��g8�P������VS�!��wu�$�~l�X�S���u=j�R[]f�n���=�Ϙ�fLX�s3>�Ga�1K�j��2��,��n�����2�S2Uȳ,4�3<��'.� ��n�\���y2'���{���/�����T��:��VX��84�^�� 8ʭΗu�o�Q�Y;��z$��[:VQӘb���+L)�{���v�U�����7<#�[w�J�=CO��^��:��޼�4O-�΁���[��y �0��h��M�7%f	Tp}������eT���L��H`k�ʌr"��З��v��i�᨞3�Ӝ���묻g�jcp�u2K�3�H�2���Q�Ծ,1��^��K��˯ho[:�c�A�ˉ5�[�(awr<��dn�}$�phv�֍�&�OJiWE+K$�����Y��Ҧ�+��>^� @�GT��HJ�$d�"�,��
�(��XLњX=���;Щԯ
�X�Փ�kv�[��i��9s�
G%u�xLl>Ւ^zqO\���cߩB�e?m�>���ɻ�mNh�bq3<�b��Д���3��{��q�҃Ǩ1r�\+we�*�3�s��W�Ӈ?w����O/H���,��c����:�U�	ȪB+�s�0�=�L�\>�4�3�^K����/\�ۗ���A�ӛ�/��c^�r8)j�����JR��1;;�擲�
3'(����*���.ԧ��DdDw}�t>GP�G��^�_^�kE�z��w2�3�j�
�x#�/���S�׆��Q=#�om��w.r/;͌�W�y#3�_����d�c�o�L�k{V
�=�-�U��O�X�e����d'i���׉U�"+/bU'�R�tO<۲�\� >^�=��|��'�V�}9]+�Nx;��H��'sց������\�І̮�˶�i��hX�p�D� ,�h��$�$9+20H	�����J�L�$�1��������U�s�u;����8��a�R�)|��#2�j�Eѐss��g��������8��v�:;��L��F����5�*���{z�b�K'�Ϫ��,��� <|��e �x_]��i�vP�.N�z:aa����Qps ��D��G�I��z'{�s��(?KJ���٦�E�rr�HR+m@üÂ��Vǌ#���^�+:	�4�:Z�ǳ�8�<e}Y����d?E���
69��p��o�ɜS���FQݘv
e@�D�z���7��`8db��6�RU�Eo�ޗ�1���P߈M։����R:������`>�A�N�l���ҽ&y%��q�l	�G���mH����te�d����&êi�-4������x^�Wu�b�����X���<�&�	�\b�����s^�Lc��Q_D�i�b�)\~$���`�t���Q����;�����`1F�dbI)KK(QDR�"J%`Vm��6���g��W\����5ݜ��t�����m>/���Ky�.?�{�����b�5��K���e`�rY�[+��1�Fz�K~���x�f�j������s�C�5�ä�m�,k BuἮ�FM���=?x��za��_&�)	�'P�1޷z�Ďpr��Z���|YKսg��w"�n��g[�^�B�x�-���k���@�n]���]��W7�U���К�����Gnƅ�	��8;�v�
� L��7m̪d������2���n7��޹��r�w3�����ڹpߪ��?��~nE���ZG�1d4:�ZȖ|�>ͻ�Y�=�_�� .�U\����"�<�����Ơh|��z?@��e���/�������U��zV�l��sГ [��,&Ck���t|-P����Y��yM��{�qE���<s�ʢi��M�ŢY�<0왔S4�ֿ3�~�mvR}�׎;\t�;�6��s@@)�<e���k9�ư?�Ӿ��+Y
��"4E�%�dm�L���oA�.��u�1�B�J��z�nL��ӫ*����ʬҳbf򮔹�s�Qf'�������Ʋ�.��ݲM����Lz�$�m���*��L:!���?Ģ w.�&U��Mwk�qk��;�&��ٶX*e mL��2=��Gӄ�m��>�SQJ�HoS���U�j����N.��h���ԙ���c�\���#�V\�PLh{�ף���Ns���Ū-N"ٰ*\�������W`��t;��y�9��1�P��e�GD<�`�����0O4�e9�=��b�>;�S�����w�פդjΦ!�k;:�Z���-y�9-X�=2V:_>b�]�+�>����f��T�w��-6V�P��κ�/rp�\dq�f1��� 4�c�͝V��L{g����t�嫡�Ճ�\Dz#������
\Y�3����i��(-���ڤ�D�J�#;1�aw�,^�}���A��N4�>�)�O/jĻ5���A�s�Ѻ�=w}����k� |��`�	�sJ�jA�kh�CQ�1(�2�Ӳn�;�C�5D�F���Ӣ� ��.�*oº�vv���̛�y���4�����o8���7�[��h�F�˳i󉑥l�6�x��	(���thdX��Jg0ֵ�Ś�Yӆ������k�	l�hK-ATb�7o-��w�M����]��<�VX5���h���W�g���ڂt��gkYl���~�켷W���,kJe�ot$�=�
k���#$���ˋ��������0�Z$ASW�tڵ��%^91W��o"�.-��B�1��'~�Kw��	Mc���E���̵�]�u.V�f�P.ܘBV�<�;צ�l=�nkruT�S4"��(��V�&s1X#��iS��_�����b�n-��e��N6 �cq�޳��}�m�Yx�d�t��Ea�tI{������ˣu���}��+❻]Z�uU\LT�!�^+@J�gO��B��n��{�o�$s�-�	{u�;�L�We�X2��4ҫ]��ѣ�}B��әv/۵TY�����^Km��{�W9�{,��fG'KH�{����Z�	*�0:Om�����&�]ޱ��\��HH+M��,�}�����>ף�O�㩫�D�l��^^Z�be�n��nX����0.��d�U��Z��;m��{K�������wVWj,��{3�:m��5/h���U��;urd�6S�v�W�,ܺ/��D������^�!q�8�Z����.�Rq�+1�/fmf�V
V�����(�W*β�`�cB#��sBӤ�Q3N�n��%�yYW1�;3�{��ດ¾��{�ԮV��0;P�.#�S�2�`uu�����ҷ:%�e��Ԉd��U��a�cEpN��sh�^��2�#@�՗&�r�$�F�d�8�C4�J�ow�`�d�B�F0��`��Z��9��r���t��Om��]%�j��4�v.�@J=�B����]ڎ�.ѡmooe��#Z'�V<����U��]��j�\�n���ќ�h�k'<G��V[�I�Η3�Jß4��E�b=z�ݫ�B�}�p�K�V&�HնH���׵����Z6��УY�t�r6U�{=}�Ɲ�F�	�H�]�T��`(1Vg5�zdg:�W ��p	>�-��xR�2��yk���=�[꺹f^#��ħ_,��[��p3��i�Z�<��0ӛ�kwl%�=XN�9-1�uKA;Ip7°��N�G�e_)v!�F��2EZ1\�,�||ԝќ�Ǌp�"�.�]��)�ʲǻ>�O	,L��n�>CXzk-[����<�L��n�+���w�����#%�WMR���w�1���k�U��c:f/:��W��VW'S-�2��2�ˮH�>m�)j��o��p�c�s:Y�#�c�Mu��hc���,��U�R�vHL}�5P�L�sH��3~��r��q�9tZ^�Q����غ6X)�\z5H�ʪq`�=Jk��z�1�z/Z}��;]p7S���!��0=�;��$�Ǣ�2uP�U�[�a6C��rhf�g[��V��k3���������FY������9��ф!�p�
�5/PjJ�==J��iiWd�^���s�؝Jxz��N�I|�8o}�<�����8V���#:I�8����pR��w�#�3�hr-���d�c+Gsj�m]�DF�\t��
`��uS��˓(��4�4���s�׺뷗��T(�$ $1D��@P���߹����;�������G�v��yi��_��^��8QȮK���X��c]/Q̶s(&��vN�b�.W9�&rZ�&���:oh��l��<�%i� f���I/H�t��5<:�ވ�J̹w���{���i���ϥ��\웩�\�=�u�"�`t�v����ҧ\�h�/!r��������_w_�=o��p�5���A�������%i��0�Y��%�Zv�.��e-�Ǻ.��A����N��\^�L)�K�dT�����)��<�n�����T�:������L>�X��#R�@�D񐚝Y-����^%u�ꦔ������	�^ߑ��d����	A�J��.2����P�6/�^����̎B|jXj�@w.�ڠ�y=ˀ��DG�*f������H8������|<�`pK���9���"��M)����s�J{
x�:?Doκw�$w�4̕iD�� �H�T��P�3f��X�b��iE�YP����\�H�T�#(��Z
����fL�����5����Km�����k�u�{v˷{�s�-�`�8�9�����G�;q���-q�*]�{��0�oToFZ8':��2�lQՙc�]\n�U��������&�f+UGv����{&9��P8\�T�#�	�OI;/c���{є�4>�&1g|n4��X��+�ffVRz8�&1uN�!
f{E�`r&�����{ޫg�scc�۝o�:��uUR-"K�)MK�i#<���J�������hS;�5:��5;:�����S&.x�drսs�'\�n�xm )7�������1���գ�_UY����&76(�ޭ���B��=%���~oĪ�6��� ��ٛxjR�W3���� C�Q���}�No#S5bP̃��s�SG�xOfE0ƗY&�<�=خ�p����0et�jy�@X�j��_G�U9��ǽ�:�+�^�}B��ղ�I9R;�*ju��.�X�#b�j��� ��G��J��,���)�DXd���4�6N
�M�y`��!=�V��G]u������!�3^��6�f�K/ew�b�7��ÑH����O�ĮVd��@�3�5�9i�P��V��u�� [g��ѓ���.��{�}�k!ˎ�AIY����h�3P=�0X�r��Փn��7�2y[�9KWKYwOl�&g��~��+��������jSή���V���y�B��R1h��	�P�`@�\�i�˘e*�Rw�Q�i�Zl�k���u����(f~
 _H��S�7�ޗ��1'έ��kk-���`��Hz�㌓&�fo���������'=��r�oGۧ� �Ѹm��ѥ��!ڦ �D� !�eSTfO-��ʉ��B�[�Q�.��;ٸ�JGgﾑ�����߂���f��6�MsC�]5�V��#@�Yvܡ���!4�x[����,aY�(q33��I�y6�*���DDGTV��8�[Y��������fm,d�G��??x��g�FPKyV�wz���{C����XpV���6a�l5�����t�n�.�b�;1H�](��gY)
�2���7F��˜&���q _-�烨[F!�єخ��8�6�{�ڎ[�j2�,�F�=~��������g ��98	�ʸ�S�	�juR��a��nc"s2a�Wp�.��߭s7���cb��z=����>;]�|e}�U�!�e��r��R�0]K�������:&dD�g�fOg�B#�/n��SӴx	r�9 Rb����}r�"F�~��櫎^�z�Mbu,���l�F�t�%�0������7����ņ�em�Lƻ�te�;���v[$�{�:~�
����\W��?Zt?G���_�6u���Sk�ǣ�y#)���ʅ�dpP:��ʵw�P��/ggZ��`.�T�x�>�{��x8N���_���\�q����8$=��a�eK�$��Z�t��Tg%�(���Z(@��(�/-0�����а��%��)ll�`��
�d*EdZ�"��QQ����"��>�@��}�����f*�u�u�^��1����H����8R�sn��Ƒ]��Fʮ�Β�ٻ6��4r���ܣ1�:�Y�������	�[27��ޞuk�H m4^d��A�|냌��y�2��\���� �\��� Pũ��M*_A�Dz"~�p�����oZOw�
���z2�-��u����20{�K�U7�L3����� �����@3��_x�ݵ��U�俎U�E�6��Z�=�0������9��yT6�Љ\Fe�dT����ޏb�2T:R�H�ї�=�%7�i��T?)����CB'�K��"�������8��dnb��oܔ�-F��xk��Ub����8%�wU{��D{�2��������`ctY�Z�e�h�,�X��S�z2�3�v;�.
��V�*Q� -7_zL�{6��b�~���_��EQ����^R���������ޱ�����vI�,��H����/�L�����7f�{�wF�q{. ��E�K۫< sն��9�qB��F���gnN��P����r�Z�n�.�k�
��$��[�6Zs���8xY�9��1ѷ��rA�^shy��C����5�%A�U'N��!	�}+@�D�ژOV�L���%PUr;��f	��su�����ߋ���UTTDD�W��J4sF�P�2����4��s�D��j=��9]�`v����������ǀ�DDt�n���v�@G�s�Ƨ;6�[�����-<藻�!���@� ��<�@䶐�yeT��/�!��Cxΐc��ս�˗���Ϋ�4�0 ���O
<$���Sj7$?R�P�Č�5�麆�G	:��q�3��Xڮ�ձ��^HgN0e�s�I����֗m��UTp4�5]P1�8�_V�ғ�*�9gt�q*��M��g0�<�ޒ@����=��϶e{x�ҥ`�*fJc+dDdF(�1+�3fd�aF1b�0`&b@-�0��\�h�#"��b�
�mh��L��A���Wɔ<7ptK�}hx���R�.�|!��<雽HVQ�o�LrwZnh���}�`f���⹾v������xQ��sF�[���M��x4�ѡ;x�_�	T{h�4��%n��V�w)������%{�fP��t��Տ���NN��J��ݨ&.~�%|�{]Xd�o Rv�c�{	z��.�F�xNӑ����:�����#㼳6!��j�J�>�z;h~�?7�HUS�r�ewO�lol�suw���P`p���d'�.�9.d?�()��U�&z�t�����FG������}��.~��h��#���j����Rˆ��([DXN��V�+;;1�0�<n�"B�@GN@�2�EM1N")¿�v�����J���Tg���f�����u	ڱ�d��%V��W;xh PBe�xa��w����{"�
͒����`�rq!De�;(|4���wF�G�	���]�4�{N�R�}A��v�`V2U Okc����c̙�"1dHAT�$�B�
Ȍ��jh�j�-w�O�Á���7�j���E���w8��(5��7#�.�Eܹ��M����˔\�V�+ *����
�D���}.gC���h'�*����9�z~�B�N~��N���Y]s'�x�$��E��g������Y����|\mJFWL�{-����� #"=�P�wkRd�����2.f*��3�tG�;��ڿQ��gj�/u�O���V Sˬ�v��5��)gu�5m=�>�DG:�>-'{�_e�^#;�u��=��5��cn*܅v�qu��懃�RZ������=����;��7^}���Q�b>�S�z���iӗ�e�2�҃e]m08��T���.�cT�a��Ͻ�Z��%սQ���:�ӓ#���� Ǣ=����🃙��EUhճ��ٌ���W���V��ujFdoǖz��<eg��S������U)o�DI�����v2�&kO��3�����?P鏲��)U%�$���Z<��� A�>$��ګe�׷]��!~�a�d�dp]��y�+�miY2��ȭ%�4�X2Ld�Z��;ޝF�X8�'4uj�m��\d��qN�|���<�h�A��d�=���p�,L���v=�G��|����~9�A���,�,��
�7�`
"ԭ�Z� �K�x9�r�U7�Z���YZ�,�d�^����}�|a�y|O���s��wq`�����+fBN�#��Bv��[��e�^���-��Ѐ6"�Q�2�V��u����Bt�>�W��Y�u��e,�M����0��P�k`�����޺#�����{��1!{����#Q�5J�@x�@@��fG!�R79��O�-O.�:�&���u�|�r���XvE�Kn7��i�;yn)���OooK�|-���fo�쏛UTlk%���Ո:L(��s��~(_���ó�˼o�9~H==B-H�磌߿n?ê���IyXJ�m(8�37�����5뫯v���u�M�*b�[xp�{խH�AMV
�F��Y�x������Y@V�R�@�+2�e�ɣn�Ԙ//A��R�U�Mpc�R�*U��b��ƧtDs�|����M��U�2󛔄eM=��n����Z�EX�J'3'�sg6��[,j�Qpa��W3;�sO�Q�h�J]�\UZee�t�:"�ʱ�%b��b�
�{��p��Du v]��{��#�їU�y��Go5��4V���~��<qR{����f�5�hL�w{�&�����ÅEw%0�5�m��Lr�,��J,L��� �VX��KIu�{���-[����[&�s.��Y��Zf��oAc��^oZ�H�H��ZM������rs@=n�m�3��8TA�=�6nYn{��S���ü���\/>%�Ѿ,P�$:5����4ػپ�����gȧ8���ͺ.���-���#�gmF#Md���Ev2ff�`�ڕ���xn��cW�v0j!AI���;tFV*iQ�h�N:2b�3FP�Q��V�|��S�,woZʔ�n���V[�ƺ=�ӑ�Z�e��n�x��QL�M]��ū��aH������q��|%�W�c%�#32�����
FV����ٻ�J둗�3�R3�tyLrw�shge�<���c��9ڲ��#p�j
B,��vfr6A��̋j��iV���yS��M�RM��w;=����'AI�5{�>J�u��d �uv����ͨ�ƞ�>�½���2N�l�[�tٙ;��u��Q�eh��e�G�����TO����Ewëu6�6Ϋ�W��f�	5]mo@&�ۥڣh
8d�]�J�e'fX�I����(�ڵ��)�(i��r�.�X��;ո9��VЦ� n�a+�z���~Ͼ�M���?��#Jv�'V����y��n]�q�.�+�������a�|�]����NTly��j$�����!�GE�Nm򭻒e<��m��=ۢm*��k4pӡ(T�H�\hU�o�T5`�ak�@#fQX��'U�z��{(�PB�EzP���wm� 4�a�tz��9k���V+F���5b��p���J�:�d=�hn��7'�cZ�U�j����a��j�r�@��6D����z��YOAxL�Ni���!��n�u�4�ײВ��'U����r�V>&���ZƶoUr�o;2��K��g�̭{9OZ��G"�׫��[��'(�Wr����̡z�=3 ͳ��;�NK0	�bU���w]$sQ����[�Ik�x�qV���Bw\1;���;"�xӬ�7�<4 q�I�t8���]�[B�;{�������ˁ>;��L��E�d�Z����P]l���t�&�SV���d��)�mh�VW���xM�����w�-��򻙹�'�K�\���іr����*6+��GTB���=������1�_���#=յ�r��{ۓ�N�f�㣰�����=�U�+Wh�%wCՉJ�����@#¡�|�`:r]�8�����G�k[�K��ٮ�������b��������o�_�p��P��Y*�=�&O=��,[��(�f�C�d���_��{;���W���rk���h�Y�c	��8��΅o6@��R�	H�����\t�{nsS,]:��3�:(�C�A�/'����8����ᢟ��Х�9Ȭ�eM"c(b(YP:2�E5&�$]J� y�=��" ���
�Z�)S[g [y�k,�t��Z���f6�p� ;�U�uL>�����v��C3�6�mH�Z�ݽ�n�!D�l�I,�CC�
m�F6ݶ�ze�cޏ��=�6�f�Nɠ�%}����?%��o#5�xy�t��/rR)ǅ�s� 8���cE���\�e�Pu�*tb]_{~��/��p)���'ޑ�r;hkA�w�#��=�	4������{C�q�WǸ_qpD6�p�ej��׾Am�^S�#ߪ��ǟ��^G�^7:�c����]M�]�Ձt�kݩ�s�מ�3�S���T���#�Ã�̺���S�+'kޏx}Է�[���-�+��Qd�mҭ�40:6+Y�\Y���񮎖��澰� �6Oq(�R"����h�3��9����[�^��FM���t��]��
�q��FL���T�R����@�LS�:�eq��z��z=�z ���tr�&�����v����T~�]G���-�3����׭�}�k�ٞ{ӿ3���
Id,��YҁTա#)@�FF �� �0���() @HV��P�J�"���
�<�d���m���{Z���w�֮�����Õ��+&���s���Z�3E.^��5+\k��O-]oF�\1�qu�e�9��p���vG�6��,&�8�.xƨ�B�Iͤ
�v����T^�X�FA|2s�{��aR�E�Um�S���3d�5��}/sQ�M�WO�y���#�ɹ�4Q:V(��� tG��W��v>>�������PB���d	��f�4�l���H� 2։�\�L�OQqs������v�2��y]z'��ON	��ip��p���5R��,rw+;L*sæņ�B��m
P��[Ш�,��J��i�4��g&��б����_�������P̅�ܲ]-�bq�̨������֎;uڛ�;�y#s
e�����=i�-�t̊%G�=���?3���t1�2'Oè���Z'��;��	�iOT���ls��Rm��k���ٝuN�qrt�\�!�""#�������[�v����H�L�,R��Ý���fP��|�V.\�4�֦��[�L)ݹ1�\)�o�=Ԑ�o.:;ב��Zܴ̩.�����Y�>!Wt�{��=(\�*ǦY��t��5�����k<o��ד�0�	p�v-�x�"��vV���Y�)�/z��5�E����P�O�:�1���((�����zJ�5��3ܴ<���#�~����$a<�9���C��G����N��11���h���U����, kMR���F{�z"�o1E�ս��R���l:���{\���~��ٺٌ�p6~�$����>����E18gpȐ�H-�/gC��bvE��@�w�*�&�k0�;Q��E������Qe
n~FY��9�l�:�e�rmԹ��0`�����M2��S�z�h{�+����|Vz3����Ӷ�U�0����Mz�"B13���r����F�7�>�H��Ǐ��t��R�)3���˩��ǽtwcӞ-��G�dcA,����gWX�"I�u����5�B�7���}��8L,��i-�m�G�<�w6ܩ���c)�A�����:�.��k��>��G���4%�f�i��@���וֹqY���ٗI2���s���˖-�d�fC�8�1���O^tORn����'�4~��k�����@ą�u�&~�!!a�h'�u�,��`ݼ��׎��XfB�Ռ�$۰��ET �Ol����E�a�5G�Qھ��9QX-��BW�&u��R�q��oJ'0�Nv�9��pY+�Z�`��������U�-�(��_i]s�:�srv�d��X{���~^0B��p �'�u54T�H�3%˕%���z���96.�zO��D{:-�
D�z"=�!���4ש[Xa>�FP�[�}�sNy�W|.����0lƵ�P�L�r�4��d�si݌G��M{ޏG��Wk���O���g2�b
3H"H���
�tMj�O�g;{~��׫����d_A�%�Q�x-�.vɃ��ä7�YlX���
u4O`�ͨ�I�;��LKhS����l�M�^��/f���T��<Jf�ǦS���{%��YLk�[OQ���4
�IDj����:����:����ϧ1��=%���Jo=�Q-�%j�P�:g�8��a0��r�\�9�s�Os8����LG����0>�Z2�O�����D���"������oy��C�nWWa�\��s���c��:e���� ���@z=�������OY���巙��Wr"�IC5˖��H9L��b�%N~Km�1���qpA�r[�;�3��u�m��7)�+��w�Gud��,L��Ȯ�h��8��l�0n�1�U'��{j���
�z�@�x9�	��ğG�쟠���atJ��S�о/vWt�����[��-���*�=r[t1�ء̜�"��'��~���5�羖2��[*�*BJ��ZU��������ﹿ������f��J�����\��Y����:!�k>�IC����n��$�xa`���^�8�͵;�yh���sO%]Z��d��$�m����k����і{�k'F;���e ��ڇ�)�����
�k��%����T��Ǻ��������J=�ws��mc��Rب)�e��Y$rє��Q����K�d���4�$R�b
q���
����l���'d̲iU9+C��z?����n��b�U<΋����oY��`��[,�v|�C\���1yJ�^D��Ⱦ���x�$�v7a��y[�鋏{�~�J���� �$.Q���O;�y\����_��֊��N封��4HD��Dƺ:"�7�6��Gc�U���]��Rֲ)�z�s���L�x�9JΫ:�>1��J���5v'[���P�9V{��؀oY��Lc�� +%��Z$G��2p��Y�@�u�*�`�:l�j�'�Kh�=���� ��12��Q!��R4�)U҈��*J�HE!�*L`U��b6#T�"�Z[)���/��ϼ���-���P&��F]��c�Z<6��ɵ�+�n����>��	�
�6�f��v�����u�0�dx%�ݼ�;��z50+�y$6f[��.I�y�|�s+�y��E���Z(�zs��}w:�*Ce��7��D��gb�.���%]�h��2�okv&kCmV]��۪�i��H�@�蛮�#��\g���}_'���@)m̊xVa��'Y\M$��Q��)�X�p�}�^��D�yӈSl��O_]�J���_��+(l�I����6��'�T�ù��3�C��Ы9��N�һ�H��܊���飮墶N`�C�\�%{Y�D|=��zXh�9##��TG��";\���-1\�������kFΕd�7%�KgD�xb6�*��\�6�:��;�m(_)�`�/�w�1�1Y#l��� ����ũR�M+^Xo�U�Y�@%4܀��Sj~��1���:k#C�I������������x!��E�^�����K�3��Y[|��MEX*'+6�yr�����h)�����L�5y��V�@]uz��Ͳ���{��][��� >R�K�A������˵0K��*x��Qk|�,3q!!�`橉�^\G����O ����˩�e{�8���_b����@g@�U��@�;.A���l��V��[�9�/x�#��߇���`�쟾��f�0(�m��ﾝ`��\���\L�r�اY5o�V#���v��V�ž愫�����&~���ѐ��RΗ\��)Xy}�A��-E͊ݤ�x�@�Vә�[5��:���QM�3�x�Z�����L{F�W�S'�ۓ���Ia3Y�x�r�괽s0�(m����]���b�g:0��}�e����C���>�_�u�b����>��#�7��+��ō��r�����aE�Ү�l��A/mܤt����6��0���G_iɌY�j����2�~��kT-�^�	�uv��8�q�ԝ�r��VfέvM�&UFէ���#�ѹp*�e%مY�qZ�;�����{2ek�/�:E�5G�~ԅ�?�ǔ�V���V���u�����6T� �%y1���E<d:3M��6��.��	��N�n8���UQ_D}�P>q�Uo��H�[8���:i�7]��)r.yӨ�,
��ӆ���f�)�K���&$��BG���z=EK1�x�㝍�b�P�z�ɹDk�vU2e��(]I���V42!͠�vr�a`���4҂�<H�<�����{�G��f��������,���_����j��dQ��h��Yx�@hs�P�܀����s݁,��6���Z����Ւ3Х~��Źb�
~�D���kZ��V�t�4��ej<������Ĭ�W�*�|) q{��N��aJ��� ��uUUT�s~�ȫV˔��̢�ِ"��3%r����^��CNZU��e<�jF��}�h�ڪ��h'H UK{#��vIs� 8�NUΕW���.Wԩ��xCO(��;y}K5R�� �>APY�0]ð;$�u�SpK�|�*�5Z�U 8���c����?�֧w���MI�o\_s�Ó����SL�l`��]L�6�Y�L�M.\L娈�Q+]Y�ب��j�[PM�i
�t�e'ʽn�sV����Ĩf��o�:��8>π�����;�m�mwonQ���`���`�_�|d̫���H��e���SB���	�!�̀�u��J�����n�iiN$�����:]hCNL3���t�h61�l�5�׷w����F���+U	y���1�x����ϺC+^�`��;���w����}�{(��5�V�t��
h|�L�*T��̪�
j�s�_N�e��/�8�H�+�d�W�J��{�JW�J��]
�U���o8��:=&8s��s\w��:a�5sǞ}��YմG�%��\��I"����1����0�3��m�67㨾��� bv�՚ݝ��w��껖�_y^iAx��l�`%'������yY�]��1���a�ǻ�^�K�m�)�a'0s,�!�ܷ$Z�)�%��@��t��F�f�6�I:2�_0�����0V#���]��s�]���I���#5���>x�y�Xu�A��5�ɴ�^r��-s*W}C�d��#r�R���/\��H24LY`)�TF�޽��ٱ{5����^��C�i��U��j����CCD�3�-�&r�]}���f�Vb0��(+�ku�j�;��\�F{y�[EL��\��*K�b���w����ڽOy���jV���bx��c1�j�F�`I΅��(n��7��6㙼x���ɻ��f]/+�yVi�bWO�h�x�Gk 85�[f�I�mm:�J�M�Y;�����48i����3v^��湹}H��� p�ffI���N;Y�q�m��(l�]L�y6<�c��%6�@�4�S&��[@YB�ܾ�����$Ջ� �{�V�Qv7�2ɾ��s�W�Ն��rY���k�x�5P���##7��:Ε��.�^�y4�r�%ʎP��l���A�u�'ܯ�Dy�r�w��JY� �3�{d\��㏍��u�� �X1��cɝ�rP�yӐ�x�#��fh(#\[!�p�k�K��2��ې��	N��۵��G$�z�.�[���Vf��1{ǰ�u�i`�k�����e�b��$w{{��XJ���ԙ}Ml��G|-�t�0��͈NN�ؚM�n*�u�[�r	�WP�����Qn�Z�6��:� �����z�V���WW1+jã��.@��o�����B&��R�R\@�7m��zz>�O���Մ�I����T��{�b}Q���������s2���Oe���NS~R�o\����^����&l�gf��M-�o�1��5�+b9W[p����<ב���s��ߧ�ɔ�O���Od���8�q�HB���|�Z��3���_��T���̸Ƃ[ㆦ��D�V���VդP�˯�Η�Ռ�X����*v��`�L�H����T�R5S1�t |�w �2Ӓ������Z��Cq�nӅX�]qрdDl�����ޅ��r ����?PpZ�|N��+Lx���5!�J��I��A���D�eC�s����}�_��`��w'�v�E'�o0+�I�Ǉ�юk�f�����~����zһ��Y��tZRx�<
�L�7�J͊�?G���*�_u��+A���%Tb(�1DV�-�Ե�TA3+�ժ%�-U�b��)%m��*
*-H�J���,b�1�,	DH������J�A��G�4*������yY�o;��5d��Ӿ�(�w����M��s�ak�F=3���l�z1�X�b�����}׻˥�@���`�A�:@븃��\���F
���;��]���A����t�t���h��ph>]Յ��(E,��٧}wR���ogoޏyO�3�����7���?�R�c.@jzyTҝD��WJ��R�� ������}G�༽{;�%�q����r�8w�~��쿎W�W��Ѻ[Q�'b���=�'=���)	V�b�H�%�*�be�k�Mi�n��p�;��֞N�����&��uO�^�z=�#�&�����?�twU��j��j�1|UJ��wa2�%9�hm9�kU�	\K�1�<��N�>�{��MC�����vc�8�)�	�P�&�;2����[u�q�Κ/^�^��1Ǩ	�$+l�¸L`)/-�":���Z=&;��KH|2�����r���K�B�:�1fS�0��=_o�u�|߿_�8���PEQeQ�J�|P�\�y�����	:�X���5%H'eZ�aU�����ݳ:c<:�Q��xpD�
t7$�I.�nP��M�n���k��`�i��xi��A������# �\΄�C=�{ލߓ�Iଗ=�`��@�ޙ�y���Ɉ����Z�0G��WG\���B�B�@۵r�u��~�tW���I�SgE�O5(�څ�1�7��p9�����̇N-݈������!#�YÙN�}舏V��Z�,̬@��"�%�~�7�̬�k�@ZJKn&��F�=�݇5���\k�8"�5(��14JهH-�����BrB�_}��_m�]ty��$A��6��/Q�ٚ�~��E��i�����In�q^#Χt�Ĝs,��|�e�C_���(-<�>�{�f|�]G_��+�n���E+�p&W��U$	bQ�5nz�g8�CRK�24\���p�&�������v����0�"OR�Uԇѕ�y���b*
�b��*19��.�����^P;����{jX@�vv�����)�imb���{���Tg1t9�J�����n#��ϡ7���ܿf���RuJ�&H��3BįϹ��L���0�
~�U�d�|e��f�9TcElQNxu~��k�q�3��r���a����Kx���o�}s�S)��0(M��7v��z��T�p��ڗ�{��u-�Ҡ�˾���VHR�4�`w��'�VA�;3`G%�]��4����/�PUBd΀̓[����j�]�ncӧI���h�����XI�����@S�d�įb��Yr�3���lqӵ;�M>{2��ۭ[Z�<�`*!H�MJ�CX�l�	���J:�|�g�9�j�N����y}j�\J@43����Zp3�A�(�k�g
{=���G���%�Vr���$�hVW��^q�$�h>�~�<!8ߚ���[��SA>}ym^n~����O�2�酀�?Q�8�J,�\O9�q^q��H1�HҨ����! � ���~fI��D��sV3�i�C��N�TCr�&J�+�H��*�S¸|��7wj��ΚʵԠ�WaV���<kzaVb\C�I����ݮ�G����F6�	˙��$G|�(z�Ga�cR�Y<-2�Dw��t�����J�A�O���>2��Ͼ��|t�&���Q&�ga�tr`�:˭��LN���&A�T��e];���mLz�в�u��0B�*�)��TS������6�B��:I�d�(��NΞi�5;�	�c��W�'0�:5�zud�%�_lmszH{@ʼ5Bh{E�*ҥ2�/8u�,�Ǥ=�����G��U���,��<a��los+�3���=�7G��n�?DG���������k�tb���Ϟ!�뵳!t���]b˚9����B��焸ܦ�Fہ�S2ce�9N�8��"L��y��2qڗ�7�=-��R�
-��!��������Y�DJ{d>)�.�-=����b�P�  '��x'+sP�>�Zkf*糮�+.b��uZE�����:��y�h������D���s���=�^:ShV��@G�n^�ߴ�4�nj�Is��O�ߌƥ�Fex�H�������C���E��M}�@D�gml����(���w���_BA��u<�T�Lyp��UoF�|�%ڡS��æ�ǋ�;���uUUTe��%֯{Ln���^���B�K�>w�OeU݊ݖ0;S����p+٬��,l� g�#�p9j^�6ߕ�f�v�㹇3��>��}Y��r��7��=%�`w+}8�k�2�E�UH�QsVk�����D�b`��2�;��oV,]��c~�W�~����W����G���G>���{��p$92A�������6b �\+�4\�������k_ܟE5�}�;�q4���Kr�<�-N���"4G�r�Vy��E���tb�k�J�t5�!i�wWQ�hٞ��|�ڪW������3��qS��z'�A�Mk%�n[� ��`���#&-"8[@EX�A�EZĂ��(�D�qF�c$L2�"d�T%ˑ���)V0
$�'Y烫g��e;˩ߺ�
k�YPQ����yA�����r�K4�A�X��U�w �o��,���jd�v�t7x)o&Y�c�\�N��jy��v:�jn�tA����lA��������`��sUSaκh�V�.>���{ލ�����;�a�9=��������zM��@:�DF���ҫI/!<t�2��d�E�7蕿y�[���]�y�s��h}[#O�!l���� 9�����"�U�g;ϻ��|%���wkNi�������8uDr�9] !��G���S��� [L�w3�u-��Y�X�I�Ԫ�s�p�#z�/T���i*�t�42a��j��6�踈�}�.�~�f��xg�+9�m8��
����(��z�'��0���jǫ��o�S;�xa������[@ln$e�*&��T�_ǫ��6��#5Wev��ȍ�2�
ec�x���,ڗ�ٻ8�g����1ނ=��r X���0���:�����4��3Ψj@[|]��WqL��bҠ5��t×ϣ����MPuK%G��<��EK3U���U��B�^aT�rw��0�J�
����<�9v��H�<zz��b��(_����J�1�t��%9�� h9�]��;ȧrzu9�^�����u�rk����4��d��ڇ��$s�NX��L�]
*4�8�O�x¨�F���ӌsZ�E�̎; n��������W���/��Gjm̎dn�ʷq�۵
�|��7Γ� � ���p[Jo�.LAZ�PcGl{U�佭,�n�#+8����"�bVV�d��`f�.]�0	���G��g`�*m�^����W�?������^�3���8��0M��|~���r0��Gmh�/f�<��l�!������wU���J�l>֞�n��
�&�U�6�~]j��y�N]2J�@E��.UO"��wZ�>���]��5��g�<4�KkX����{����|�1r�XNN.U���R�v�3y��re�S"w�h�	NH�{'�u��wc�3���#��#l4�f �Y59R��?}���ИJ�.�TL��P01��F2�f���ü{�-�{�f��_���>�sa�Hd�#h]��Ld�*]��Qx/Ca���Z��nҖ�}�gk�H �UU�ËĈ����d8w��Qx���J;�K/�\������`_C�� #��25\��s�u���2�G�2����\�V�ގ��,(yQ,��"Y%�֭�bky+µ5#���s����I����@BX��( ���ܢԜy��}E2������&�<����dW����`	C�g����-�����V;�� �I"Й�bb6�X�D%}#hh��d�w��DFj�������x�V��i+�9�Ú&�t;"Ǟ�P�	�)��9��Y��z�u�\�7�?~�q�&���of�� �2+��b�AS(H�mR) ,����+�1�ir�w�:�A�E�}ϥ��ˎKiS{�ܺ���Ct�r��|�u"��˗z��|0KL2oz���3Eu��Ie^��y���1�e?�fѭ�Bߍ���P���Qק!0���4��}9 -�k.����B�f��6�����?�&��V�	���U�O�/��~��|�I0�P0[�yݤh�^T&�<�U;R��"�暢���x־t��N�gx*r3A��4��?9c흯֐����y��?w�U*�G#˸�V�0jEè�r���(�jd����OM:�V�|�u��.��Ա��]��(�GΣj����3+tN�p#+|R�݃�j�8l)�sSYX�T6܆b�GV-��zc�3tB7Cg���f��5�ڍz8ԛm@������< ^�n��VM�ؒ���h�v>�tN��::OB�dU5x"Syi��t0�΃� ��I���1m� =��}HL,�S|Np/��Qv��-3(2W�����u�j��u�x�(\Gy��n��+��pN�^�v5@�w����y߶�m+���)��n���L���)}��\�
�hWEiҵ�poV!HE�s4���^�C)���E�D�i�ˎ����f�y��,D�sn��]Sv�%�%f[D+fr��r�4R�QL��`��`�)MU�dl���潭Lv�jjeƼ�x���C��k-�`;�{T"�� |��R �/+hg���w���ußX�u�-;k�.�����鉚4�4:2���k���9�v�
��{!2	8ٮ�u���,y�u���o|��ev����[��c�^��b�׎���[�9h�sW]����/.�j#�񆈐#���`CB���(���Me�r�ea10�f�@F(�U1�(�9��[,d6�`�����3Ԩ`�}��\�z�J_���tV���%��Nk-1wo���_�cɳ�lYb���\Z�V.�#���ʤ��ASR�4��(3��k��[���r���w&�sZt�їi���m��j4�'�b�<.��7��׮�7��4;���{BA�3�0��tLb��粹�6���ڮw/�&x���
|���vЪ�+L�@�K���բ��0>��gs%�̉r�tu�M%I4<�v�Y�"��w��v�(3T��+�]=�� 8�]!�#2o���M�n�;|,�.��ZQdkou�:�
A͆� �{���C �YQ�������q�N��'wdU�6�1BtrŐ�;���A��dr�繗y[�o9��:���F��",}�t�S5�ˤ��mZHl��D�n�}Gt��վ����E��r7��'B�[�+R��u5ـN��e]l8NB$�Z�Y��S����9fC3Pf��x	��h
�
1nvkV�̄u�(���.�>�[Ԍ=5i���[Ų�d���n*�#Ji#h��3�1q�J�����9���|*瞟[�;߈�7M�dp|��SkQ�tm��6*��/����p��Xp�5��uIC�ڣZ�W>��
�m[i-˔�f��JȮ-[*0���l��p�LZ�u6�q�$�u�[җ����T�sr��(&�%C�U�.u�Z��>P��T/�en�T6���m�Q�=����
�oz��۾۫��"���V���bؙ�hw�����af�՞+V��d�zk��]��$l�V��̴�[Ǫo7��y;)0g1���S�J��ECU�y�t�¦4ͬ���`ct��]����`�</��$���m�x���D�zs睷�đ:�]S7)�:�4{�aD�[����q>��ٞ�ڵ���(��vA��9�J߰E�9q�F��2����$t��S�#��B.�Eq9I�h��wk��9J���s���~��X�Z?�o��\R�z=�ڃ�C���#����� WT'��g�"��sk/\�wz�n+�F��&9���z4�l�H��vm'�M��c!}˂�<���,[ّ�H6�S�TF�:�dO��ͧ��_8���TسeI�5�K����]�.�dUh��q����:�a��S�����]�ϧ�n�mUW��8�z">��ClW��ԧ�(L �����w+ ��{�M�B�&e
�ڋ���
[3&A�,pw*�Y# ��2����j��Oz=��e���-�gF����˱,�>�1j.�"&0�¨I)=�7��Ϯ�VGV��䬽�gଧ�#;qB`ϖWťHb�t�[r[f� 1��Ab��@�(8��G2�S"1�2�-�"��e�
��R[�eI֮ �Q��hSu�i �v����nYos�����s���ܩ/O�Jƭ�D�b��9e�4���v5;�lTn�eol��1�����5ց䜼�r�������0���)�u�ܫ
����XS��[�n�H[���CW���a�0j�ZaVQ���� -}X1���Ķ*ߙ_����)w*���1�բ�:ǲY�؏{�T�^'�*�d�#,(LS�1�ΰouX�⸪.��eQ��[��u;f�Ș� !����e� '6`��ÕL�\����?{��&Eor\�k% �Ы�G�Kyc&LR��'��Re�SV�i�Kܜ� P�i�*������0Z�`?a#�����E��d���X6��Qn,����7����2HUH&��C�@պ�Eܾ�:�ˑ6B9ho��G���\-�1֗���:��H��*�gB�������b'�ꗂ͊��4t�D��5<:rV�q{�w���E �}j/7�߳n��w��߽�}��r��ehk8 ��L��ve#�P#b��r�Мբ�m�����ngXw|3j�3�bKQ�7(�l��l���|���\�LZl{��D	��1y(M�>���.i��;5�t���6�J�0a�reda����"�[��]�������S���'q���w&���ݗ��'wli�4.��/k&����oM��:���Cb�(�39j���\�1Dz"}2��SL�k�}Z�`K'W�fx��'t��F����~B���c�&��r6�#���B���N������+3!��{�J���WZ5���L��N3B����Z�����챎h��5�{=b���g�aݝ�.6�Kۙ�U�͓"0Zy��"�jv�W��z$3��ql��*�lT[�Gh�����![i�m�=�����u:�G�xX���G�H�,丈��G�3�"""�=�6����+��gQ�y|��MZ�H�_T�*@�H���,��C��i�R,".�c�0`3r��8.��lT�^�h:�v1F3��*�rK���j]��"7��6Wp	�����7 
u
 [yL��є1�!dvvq�2+�*۶�X��#�k�Vd�ht� ���)�^11�q�����r���p#ގ3�Ǎ���<P\�@B߻,�Bd��}K����S�>����_9���HUq�,�6��V��*����"kQIr�&������7�N1����t3
���0-+���T��M�^xw�q�
۞�}ȴ��|*�{�z>8�g�lc�'�ϩ��G �\���^�_��sa��d�n���G�g��KH��' �e�8
���������]��tbV],�ng�c����u ��h�rr����?]�_u��YW�s�y5LOv'��*
����eݠ@r	ma��\7��7����G�B��f�^�˼��:�b.�H�.��/m�Q��-.k[S�6�S��wJ���&#@�n��S	��k3���f_�����y�FRCI�����3�~ך��k[����F0����h����5Yͷ��R7�c,k�[� �B��-��/i����G����u�+��{
IV߹,�W��E+蟆�����!�CQl���a�3��)gS��D;�DȢC�[A�Ubb#���N�=\��28�87:�. �e��Kx � (��Oxg��iYf	i��O,�/�l׽s�d�Y��%}G������E��<�쿅B/K�&1<�*z�Ӝ�>y)�}+��;	�I2���٪Ǻc��JJ��z�w�w��?WժZkO�|/�&8Ģ�8ԛ�<��3���w}L�Q��SN�`��,:�%7Y�m�{��rg�Z��#{n�]�mq1�Q�]-l�]���m����i��ks`@]bO\�w���|@ԙ���5�Hu9��9M/���&�h{5��F(}i��R�($�z��b�mI6��bt}8u�L��P���h���IR�	B��A@����:�?~�z�}ޯ��Uo#��h�qȝUꬠs���s��k�p;꘵�G�Ud�K<�D�mZ�iNv*Β.��<3o�)�I���w�=ܚ?y��?1��Y���a؋���7lʬ׈�ҳ��Ν��U�)�X����4ˣ�
y��eeP@D����m�N��zt��YuO��Cl�1�0��iF�\��]��'�Vls�%R+>��P4�w���80���[�;et��<bO�� _<c7ޭ���D�*.�y��@����<	f�X����cA�����Z���ӻt����Y�0�L�D��b�:����&��2�W�H�U3G	�2��=:�G��D&�YeP{؆)�F�q�<>����|B(�=��/��[�����5n���}q��	c#>�J3FU�f�"�;����Z��c�kK�L{��s���Mb�R]��M����pȉG��B+�Q�0�c`�Y�V@�$�2I ��-|������ɵ�f�K1*��]�pRL�ߐp���zѡ��n=
5�:+���V|x��$�m� 0�we^��s����u�r���t�0�P�g)g��~�.��0Ӥ�N���!љ��b!}�e �.���V-�6z4�hj���(]\�S�B��q�ڍ;r�
�����+��.������!�t<���yt.��d��&�r�G��ʮr]�� )���2�gh�F��d����N�t��1z�Gs�g��P�VY%]���,�^�ˮ���I���
�3�(�Ƣu�|r�X�V���+4�lk5��&�&Չ�q�w
i-��v7gS��T�F�tDF@g'�H�y�/��GD,��#��.����Q1�p�++�%2Wm8I�
R�K;��43�n.�ǫXZ��Ӆ����mG(bcv�;����e{\��i�i�rv���&�
L�zّ��{\��&���(O�B$�n�`5��Rą)T^��o�7��muy߼,��U_�R���y:�x���w���z66�Ι�6H7��4�V5���s��(�>���8�R���X���4&Nb�;��7��hLS�X0'���,�:�N��e��j�,�r�'�>�z=����D����&F�@_�=���
��n 
��N��8�X-��KUڮ�p�\%�8�^��]+S��0'B�p 6��9jk}�G�ب�n�Ix�@���VN����T�ˇsXо��o:аz���̩�\ˢ��H&}革˛y�?T5�W��4��R 	�� 7���-Jp�u���ő�@�R��iɘ9���=�`..u4��~��$�Ɵ����>�^��}�g�y��-�T�b�HcP�|b�2Q$+��'*����K�<�+���wV5��"���� _ty�w'l�z�q�DDN���W��#]��N��eM��k^.�&�fƴ�����18L�x�~B��X� ��B��m��Ϸ@�/� ���FNA�H+2U��Е���o`(�b�Zj)�Y�*�͓Q{�I�ϦX]�Ӱ!�\��j(�N�s���Q��b9XpIHc���������n�Ȟ�IsA���[���*��Rg�9�;�������x|J#Z��V	Ɲ��Ѽ��Nю�{�����}��p�4�Ih��g�@
u<����]�E[�JP�S�F�e
'�^��2:���G�7��<P�c��V�W<���82b����g%�5n��;��V���Ϝ5E
/0ɧԡJ��d�}��oF�dDz#��G)8ʕ��<��;[Q�G�b�r�БXG<�8Gj�3�ze+�Ɩ�òXQGe=��A=�>�-�r��b]ԝ��
p�׷�!��['�� �`�th-.��*CrΦo��S�����*�o\���d��7������sMs��A��P_0������"��>��[÷�~�������Ęȍb4J���-��=C��>o3��ͼ}S�ٽPi����|i���p���b�w$�!�pU��b$bɌm�l��eT	�S�kl�>�����)�+>�)�C��oOT�b�d�t��n���+�8��Ӈv�\+%6:W,�#���e9�hw��jn�e�܈���h7���;Z��f�=�����!j��P�PO�瞌8|�;�Z�N�rڻ'�U��X
d�ǋcޏD��%2v�#�����ր�li/T���q�=�zTG�6��]�8��G�U�p�2.��K�eu�-��{ޗt�[S�j�G��r��Lv=��98�QeNV�T�Tc��v�J���u-����ʥ�I�D]��]�MAIw(�{��d9��/�`��W��C��|�[�	e�+&�`��2U=~�����l�������w� �	$��@$��0@$���	 �K �	$�h�I'��$I?� �	$�h�I'��H��@$�� $�� �	$� �	$�	 �N@	 �O� �	$�h�I'��$I?� I��$�� I��I'��PVI��{t�:�X��� �� $ ����o��!H�0 ����)�*���4R��i	
�)U#l��(�)6�Tf�(�� "�D"��%*��  %QIT�"I%"���R)U"�(ET*)T��Hm ����	�t�UE*TUAQْ��ЉDF�T�Ѷ���Za��"�:D�A�J�ЗA�N�-Pa�f��U+ZtNE�C*ւٴ�kP�Q%$OcVڊ"UHvz�m����w��w��p� �j��`���6w]D�]*k��u27N�ݝڴfS�B�	L+"��2b��.�v똛Q�v�MXr!R*�U
E	*��<+B�)I���HT���Թ:���j���WZI(��Whѭ m��A����LF�w�w[�����J6(���3kb��J�����R�@�J)zPv����0��t:S��hf��$)���\�wg[���L��P�����j�M���n�Tc@Utj��(���5]݅V���Ww%B5�"UP�%UMܝ:.�jƖ�R�Chm�Ut�A�i���t��SWc�v��g]+@U�m4rt֕̃�\��v%]�̀�4���:I �JR)"�T����He����ݰ;k��ug4`j�jv�îr��Rn�h3��]wEX�kU��wJ�]�Zՠ��n�v6m-��E���N�[���T"R(R=(v��9����;�@�:�tk�:�� �u����U�n�79���cMuvۜJʛZiGn�˻���mC]erV]��7%�u�v�[*�iU	BID)$T�6�f���uWh6��۔L�dkM�Uvv�ewcY)�5��ݺ�n�dGwF�l�i�t�v����t�sm�m�qE݃]�u���ծQ�-�;Q�]۫�R*ER���(Tk��.�u�í�Z��U�t�Wi���+�FNحۺp��U��:�ۺ�su���1ڵ;�wS�k9λ��ֹ�뫷]�D�n�m�nj���TBT�$��D��Usv��t�u��k�2����]X�ۺ覰u#mVݻk�Jn��]�mK�Xt� t������   X�  F�lV       �{&���U   T��	%)T0 ��M0���
��d �EO�A%J��C2i�
�S��@   � 	I	Oj��4ѦO$�7[4r���hDj��bC}�5�@ 	dl ��2�DUk�p��;�	� �3ff5�����3ff�� ��}٘`��߆0ffd���f���S�333��0ffl 0�����_<�}�Ʀ>�d�5`р?3.._i�d5%���٭$X"92S0CI��5�qD9�0��Y��8`$fh��0���QJ�4��Tw{�g_%�s�����I�1v͝م
)��K�eݳ����Mm&æU��g@\�����:u��ݷKh��27Wq7���s(]+�4���z�΄�E�%p{�1e�t���`D��N�6j�=�!��.��tv�*�J��M%,�h�IH�Z�R hk3\I#L�Հ�h�b�ڔ�*��@�3%�����k�%��u&Aek:ÖEm�ӏBմo[��:1����N��ߔ2�yo�T2���#S��O/��Ƿm9u2�gh�΍��}ڕ��vθҽ�qG�M;T�ڳ����"�$�Y�����0r�a�`$���Y� 60� ��(�C,�K�0%��2��L���:[��Tn�����Vz�;�S�p\.����ik�z{4�]�j��0�n�>����;�1L�'m廷���e���+wh���P�VK�Iv��؁ҺݙYp��L2��RLw#�um���]�+:���@۵��]i�ju�8�<����{jı[˼�閃+w:���*��P~}�f�R���pY=hdjvn�]&b�m�;9v
y�,��
�Weȥ�����nS�n`#MQ��L
7J��y�U�onS�	�U(*�����6fNU���iu��4�9vv��p���Q�qm$�0� X�r���h��&�bۭ�A���r����aL�qv�Ƭ���s��Y{���a� �ᗅh��G��jb��w7H��!2��gUnS�ڥ4�g�I�0c˭�����ud#g"m`ι	��#oX<��Dc4m����r0N�zf�U���R���uv�7��2�� B3����-�4�V�c���O1*��M�m�*�i�p��)C+4�P����@����J�EZ��/aҭ�Ÿ(�,��bǣbx.<��M��	�P%��Cј֛7�i���9*�GL���t˵H3����t��2nU�V�׎D(<'�׋�~k99v��ޠ E�p�ZD��aSsWt"`���o7B���I�����LdSt"�kqU���R�����席j��j��U�c�a�&B���	=,�d�[�c҃`Ё�2�!K�4��"��E-�h(�%Vʵn�Z'�z���p�:���Nn�5�{q-����8%���HEwWx57Sw#z‵&XP��i�P~�^T����Ԏ�Q%���*�\�R�N���QX�w���hT�
�v(�F��b�Yu��E�C)7b����&����<=��� ����;z�*a`$v��j��"��S(J��bm�y�����@m�F���]�Tf-��W��V�� �܁�m̴#t1��n������m�Z�`�ՈS�K������.j��Ǉr���j���kD5�XT���y�T݁(��*�F��t��F�Iou!J�dշ{.=�� ���or�2��%Bռ�)U�3q ��`����Jm��P�	���Wm,ۭ�M�qf��8\ڋ.<N3Vm���{-Rڅ�ff����S�ՕI��YʷgY�)+�B�670P.�P�x����A�b��,�1GX[�(г ���%����m��lv��%Ct�W)��ʚE�*Y��Lyv�4�X�=d�bmmMǨ��{�ֶ�Zơ���xh�6�Á-9��q�,�%��-*̷�3��j�j���ٴ�;v%�4��t�j��L��`��N��2��Sd�ZM
1��g
���l8�a�˸�g��5vֲ�PŤ<N�VPM�+m�@���<�9K(f�$T��c6���ю�cҨD��!�� WD`��35y4�F �;5����.�@��Vv�N<�� +�P̈́0�Y$�,*��V��D��p�e\��h��ƚ)GZ-R���邋ֵ�ٶ0���4��ۙY�4��Q�r��U��ZK QA�cj[2$���$��FbBe������Գ��K+K�d(���d�@�
��IV�j�Z�a���Fݱy��n;��iլ,��A��^m#%��5���ki]�#a���M�:�F&�� ���e��.򒭓Q�?,f��J�2���5�qñl;��ұ�խҲm*�lB�R���41����@*س[�� ��j���mA*G� �աշK�m#E���4-��Le� Ml���!��1����dL�C[�˺Mf�~!Uǌ�pYƛP�����NԨX�pT�-��wn$�dD�6Tw��oI	�ɕ��o�%���x^$`JՋ7�s`̫�b��uE +1#c���F�&=:(�)�ޓ��d��y�EP:�%�̾���i�����vl��Su�;�3j6j����ӽP�oP��+R���^�:�)f\ji5v��f́
�ܑS��@[.�DT�E��a�I��5k&��X�C�����m&�[��<�� x�Jx�����;��̦Џnܘ`p]���9�Ka��X��⛳D��s��l[k3Ǯ-�v9�� $�����3Z�&�f�lB��9Q�Ym���@�I=�ZD�f���`EH�(J�.ZJ�V/�2�b'W2��3*���J�9B�ࡈ��Ȥksr�����Z���=�^�AT��%��LH�ۚqҹ��?������d�f�Y��������ꅘF�Y��C,���a
2Z� 2����9�3Lӆ@4�Ds5��02-1���r�Ub}Ï{�T;�Ǳ���HR���ރ5z�e�
V��h���@:ݤV�MЙ�D�B����^lZh@�ghS%�/x�7��r�5�|���QV-��z`�S��f0E�}�["P��w�b©iP�Yk-*������le�B��.�O�s�Y�[��w%5աp��5�U�W�0�{�nG]�3Fer�RX�n�{�.��y2���zkks�I�.񗒢�1~H!P	�Bw)��m�u4]u�	9�D���C�,���.?ʮ�f�l�����[X�g]�j�q�ŝy�Wm`wP�%���X�V�Xʗ��; ��P7����mf��3��!��@��B����S6�fVʓ)n5W��_��gNب�"�U9Dvȋ����i
��!�d��!h�2�o]fVVb��� �c��1��ؙ�a�g��+M�<�AM�	�)�Ŗڲ�o/^��4;�%(^�#hѧ��熋o� f����ݨ"�7bܥ�� �� �V�ص��^= K���6�x�%�-��BZ�F�Ի2�o2s*�Ʃ�Ń[�i65Ge<�0�@�Z�Ň�yI)�Îf�7l3���e,���F322a��H2.�XZü Дc{E� 5c��ѝ�ί�6�	�̻�N�J;u��P��&�_��q�ُX�s�H�u	�l��T��,&Ү��.6ú��ۆ�Aan�e���L�E<�T�����8X����s���I=@i
Q7�~;�SV,�d�+���X���I�r��9�a�,SͻC^][���ཀྵ/��-"`fQ�i�!��n�\)�j��ī8�m�L��t^
]Wek9��U.�9)�1����ݻ�k1\I����9��y[�l̻X�S0�y��TT�SA�,��i��D4���ý,fX�2�K\U+��w]?(����n]�*�9n�'oZ]ۊ&m�0mB� �W�������Z�a��6���k6��Q�6��8*"sBwi]1�D�¯Kn�8�.�F����o�1�qH�lm��~�)Y�NSZ���{[r��#N�ͲG�LG�:= �pι�^�č����Ve�+3�X�w1X��!Z��d�%�e#{,?HZ�n�*����oȷ�&�1a!![�u����f�I1W[&�N5D2�+�K���t��1�Ѭ� ��RY���i,�}�Dwk�"��6�Q��Y��:��4�Z4�-����ڛ:CĲ��^�����d���p����Uk�
[�=�(���MLtw&��[��nV�32��N���Y�d��j�%H[*ZBzjKt���m`FbO+ug�wGt�4�x"���%�䲇�	K�hG����s��Gk7�dԴ���J�[!o2ƛ�L8��.�P���usL�c����1�זt�
r��ױJ��n�6��XrU��Lݕ���h^JX�ǏK;��{��"x>��zp�+%�0˼�T�Q�s�6���جH��MLq�H�x9RxC��!��b"�.V�I86��=˨5Y�n�h��F��/v<�6X��>4Aá����7FC�җl��A*���������f[긜Zt�{]��/:�s20	C��MJt�Bb7�5v�� �����(5d��(Q�Z+3K�.�@��l���m�f�	%��363[��B���I��ۂΥ���-�t��qG�ޭ�3î<�.�ZV҅+7��ʻ���GPެ�IEkktK����ą�^��7v�+b���b�[
Yt�3F淪�nf-&H�P�Df�9 a����1Y���|�����\���cF�*ɀ7�3��f�a v�6���T&�<�5����aoz�w�nROJ,F��?�^�f��Eڠ���H
=o��5-�*���e�pZ��J;a��䦘V0��唿Yl63t]Dr$���#�T�5z��Vٹ�ࡼIow�dv_�$Nܣ���k��6�v�e�n�h-SSZ��*@�]zm��id�d*)��a���nD"v�[ԁ?�����khJG��@+/ ��;��XR���/��ׂb�%���y`�QL�P" 4ܳZX��D��v�W#B͠0E�w�mݗ|�45��f*yB�*�op9F�1.�zEiJMA��X��N�U�u��Q��h̨�����h���۱��%A1��T[��Q���W,���RW��2���U�(jr���rӵz�j��q�g%��[*e4 Z`	��!�Y�κN ;X�P�1�����U�#T�bXT�O,�\i,����'��2 �x��e���ia�-H�w�F���Q��N�6�dn��3w�p��m=��
V��Ԕ�f�F�]"�u��M��xC���9;�K��fm��2#�6OFuɡ-��b����\��#]�-	*�l+�So7��a�\��<�c�ϔP�ݷ9R�iׯ52BӋ2wV�����Rf�-����%� ���I�z�8z�/�an��f����X������9Y4'���kY�J��|�
�+_�]���[.�i�s8l��S醭RT���3SV���$�Nk�������Ѫ��9oi�1�^�{d�^���ERf%մ�,���N�p�DO��֪vQ#y�Y�g���Tb̾��k0w���.q�]EA�Bu]������JM�BJ�-�i� �ct��(�i�?+{#�{u���l���a��T�8��"��V�IS�.���
�D��*��H=�/zMЭ�,������a�b*:D�B
�}�75e3�J'#��2�D�����	;P.��sf�WW��WJQ�"��\�J�C�� ��S�5�n�q�+l;���e�Bd�t��M��ę�-���4qi�z��Xуi �F������jC#a�[���{,�Vr�"F���*\���_����[J�2�"�*�M�:���	��vY
�=��r�F@K��X�n��V3�"��7n�cpE��f�䱺 ����S�L���d�nB4sPb�&���U�R�o��e��jUӬ���Vat-�y4T����_��L8�$)A���v��Rz�7�o�e՜cj��[��fT���p�Xa���{��m���ڰ�L����Xݍ�ά��j�&��ѭ���&M����%�޼�'�8TBiʻ�e
bR�{=j�̊�[W�kE���0�T�^R#	sp����k�Az��c�I^�o�%�]�vl�N�e�i��im:q6�`ׇ3���3j$2����m�����;ե�D8B�K:֜FL.�f\��M�q�,��5o�ғOn-��I�#on3p���no�q��L����բn�hX3�*,5��2����i���%h��X�2j���$(�z�$T[Cm�N�&�Lݗ�C-��K%���ZN��/���M���,Ihm�z&m�l~��tЙ�f�� *��kpи�hTeo<�QXа4���V��}��P�C\[��UDP������u*B#t�vbw�{x���kb�v��Ɉ���Y�3%�-\��
Y�F�L�y�P�2i!�Ҕ�J�.ۭo{H�l7Qj�W�\ʂ±��vBêi�ȵ�k4���R;�j����-���V����Mnc����5�ۣ�b��cX�J����[2�����El�*�ڷ3h�6X�Gj�j�#/��V��t���7����66�e�i�R-���j6Y�"[���z�w��N�;S�*QJe�
e���7�F��75b�q,�z�:Q��h����m�x0D��˽�����fn,�b�N��ƍ�I�V���x����~��E7$��ҁL�Z�aw[i����4���*�ŭ���Z�bXЇ#���0y�$Ď:utn�uk�j�~Y0�4P@ +0�5�V<m���?l�ڻ��F����R�U�ko!���NVvR��Ŗ�	X���Ż�� ���-�ӭUo2T���Ȏ�~�D% ,M��,U㻼�
z�wv��vV� )�yD˦t^#2�V躳��?F�#�6d"d	*ټ1Z�,���}��uA���4��]#B3.ȩ�/G�c�Y��� �^�	�<S{����M�K��_�dy͢2陜� |�x�hٺ�ƣ�u39ζ����7���v���W�v+�dR�c����*�zԱ�]uG%�In%8j�F��X�Z��:e�T����}�^)&t�y�n�������Ў��鸤�%8��H�ϝs*�wZJn���/�8]ww~�Ǭ
=x�6�/T��7�H�I�#}$o����>�I'wt�H�I�$}$�����7�H�I�#}$o����>�F�H�I}$�����7�F�H�I�$}$�����7�H�I�#I�<ߤ��w��.=H&D�%�I%�'Z{c����|�Ki�c�(���MK�uѹQ��Z�Rm5�P)��5rg����N�o��i�G+�����i�`�"F�����6is���M����;�t�����ʸ��}��Ia=�R�ɕ��$�-�J������j�K�ӗA��W6�[���w"�iLm�d�f��������owg:7�F�H�I#��\���5h9��iG�6��<{�F�;1%ܓ�#��n-�$���������ܒ7�R[��K�$���=����F��5\�K���Ӿ��y�����7����C��m�Y��{G��$�pyfXޓd׽AS�n�R���&u�yw�ټ�N
n��ci^EV�@�����;@F@�1��+�z)�d��x{��H^�H�[��#�����hظ��zz��P�1(�FP�G�F�>uuŁlH�]����.t;[1N�湆S�%r�h�>OG��Y���krf�eK.�JX�4u�e�Z���M����<{��+%�U��H��L�!/�>@�i�u{3Cy�c�WL�Uop��؅�D"H/��pŌ��W&�v2�M4I�՛Vs��j<�:O
!�]cdv�1
����;��ܺO*�v���OWU���b/x���!65��ξKr�sj�7�YoX��������[,^j�jڄ�[�,x���]�ޕ��.�5��n!O�*:��a=y�;{�L��b%L��a�ɗ�5l��r�%^u_1o$n��6�*wp�K�,�V傮�Y!G̚;�`�i��̤?>�V��̃:3,��%CY?��]�T�ɛ�|�������к�kOueG[x�U,�늻�V����>=l *�c�y/u��J劜
sHw{�ko�R�r�p;�e��xt���G�;Nb�M͍A�nM�vv�wAD�G�U�+aV�g�ϝ�>�E��V^�F)��p<����b�
��+�ƙ�[�rZ��[�79Jv<˶�3Ѿ�mwA�a�+�]Y�H��!i� ��Ac*�)Z�$��g���mV���D4yNޚ�[��*��Q����/C��a&������g ���	�9��u�z����ޢ�Y���¿g*���WU��U%¶gl�4m���&
���F��`E��[�6N���]�	9��+�(r�<�0�g���gi���wb6�����ǌK�Uړ�Mx.������~�H�KT�����NS�xT.f��=DiRee5�R��*�Wזr�8ѐ��)�x��r<�e�i��z�+W�D�ѵܨ�9�Γ�粲�wd�h+a��s�ći�050�BS����	��h5Ę/�ԳxnY!�^����,MO�<w�t�PT5�N:��f*:*&Or�"�;X��w}�=�w(�v\r�#/j�'i1�OO�W�+R�穃v�{C��۔���0n�S��H.fL�#�]B�4��If�+ ��p}8!S2�-� �R��˗)�4tc-^L���I�A�tS;�����qp�-U����٪���F�o9�YT�R\2���[kM9��j���c����%�ހO��}7m��������e���Q`��gu�&sB����б���Y��v/�>���{)�����>U��7�L Z�������͘;��mW]�[I�(�]VU��m5��a*�A��3G%�=Z�v�4�L��y���֔7�oU��)��w�{� l�Bc��x��-"���1���|+���ǣ7�$Mɺ�j���e+R
�U|Ō�r���b�v𷗜�t/�?:�423{�\��Y����^c�Սձ�����̺樊zV=�$�Ou��)iU��m� ��<$�݆�2N,U�Ir<�)5���ɍ�L=�iI�����SQ(�}�K��巷�~�����Թ�u�ߖ^�r�U�p+�%��5��+W ��۰�b�~콇n��oD]�[;����eS�u�p��=3Χx>�]`��6l���:��
w�e��t=��6;�H �ºvFwX�u���Q�����)d��h֬uʞ[���d�����g�;��4mY{�y�U�����{n
���� �楬ɾ��v�>��ͺ���}�j�)b�8/Gw�&��.������i��R��HJ]Jb�f�mX��*Ֆ�G��Çv.՛n~�v��%�z7����cF벹h��O��`�1!F���d��7��uJ�0.�RN3;��iW@ivWj��`;�`^ѩͫ� ]iU�l�9�t�S�؆���&����J�̼\r��%��VkiS4��l3�OlAf'C;eH���:�ə�+FV����8���J�`�'�%�w+�������q͘ށ*of����wԣ�3!�.���WN�;Wd#�,�U����q%�����k�^L9�]/��a}��D_D����R0�ꋆ����:�nZ5{�z�NOT��Au;0����o��8&L�fQ��YA�w���w�� :ea3p�5����Z1�Z���n�Q�|��.�3�U�Ese��ԟH�<Ց�˜�D��]/���t�!�sF�ճ�����xh�*R}�A�3��T�2�7v̂r�'�����֎Bc �r;Di��{F�ՠ��8����jmd��e;���V+
Tg�
+�ײ��{�nns@"m_�,���\����;���/@���� �����;�����-�;mW�g�$�X:�L��I��uśt+��J�<{-���Ma	Ӭ�v�=U�bt[#�otX�c����laÆܼA�H�Y������,sc���P��R�5*WC�[�=V7q/�!�O�os���8w�ҡ_��<a�3*>����kY�\,�Nm���gZF�3���N�gݫP'F:՛��J���Z���z��a
��1���5�᥮���8��m7��xr��5����b�O2���ln�a%�o��[�`��VWFk��V�)JL��esj�V��7r���������\���̻��2�E��GwfWc��`�M�'�N��0��M�8��V'
��r��iz�A[f�ݬV��>�Wk�v���0&��.�l�q�&+�Q�疯���X�b��Q���/��{^�h����*X�Y�	|;ͫ�X�Vέw�g��M��Y0[:�޲x�V�Ր!;�Q��ŷvt�c���c��˙D-���3���_bC��3}����C�[���V�/�W	ܬͮz�Y�>E�s�K7$�Ш.�y�ݼ�?�9�^׳��X����Ra&f�+�S�L��'�R�Vo�� �K�0���S���ݭ;ðe.��Z�Q�����\���`yʡr�g8�K�m�|�i�*,�(��<g.ُ��2�
��7��i�g@gR�<�����W/y�|gr��6!�4�v:$��Z�ǝZ&��V
�ಞ;˵BB"��^8����E�n����%��ݦ���������N�)�r�P幜�-��D70��M,$\��Zy+�)�L�█��86!ٱc۾�W�\yj�lj�9�1�D�6��u�{ə��g��Oq�3�YZķ�hvd�S8�a�/q��к��E|gӡuw,"�^��j�ܙA����t����;�k(��yBB�eܾ4@�d�E*���܌#u�钷�6Hy[4�US�����@�� �fZ�Z��Q�B�'J
8u�(q�6���׸�ْ�ι��F�薇Z����p�Z��)fv.&�1�l>�͘�4�W` 񭳁9w��Ŷ���t�A���ú`{0ag9���\}�<c��b���K7{�3nX���N ԁ*�k0=�`�7zjI�CZ���i7�[i㖶5)����������Y�'��SƩ%Q���wq\3����.�5�w��8l���ӯ5bA�yN�Q׵{�#�P#׹�Qff��ꄉ�z_d�@T�(�I8�9���(�;���7[��me7�O�K�K�ɜ�W�\��՘�@�dv*m��D��`��b�A���5>��=���[�HgTK��-��m;��om���1d����x�V�THd|��G ��؎��R�	\���Y�Vظ䰧l+{s��J���T���'X\z�:�48+<����;�qf�_-�f�3h�a5�'2t�j<�{{�(�Ԧ��5�>��7���^ag�J�k
�����K7��d���U!�:�9�ך6,�����`�5�� �U
�P�2n<.�:�ġ��1R�wyb+n>�
��d�Q�)<�����1ʽ�����p�!5�3��r53)�����u��a� LJ�*���i�Q��}���H���D�L��$�r��yIWun��M䌻v5�y�y�n�꽨��$�������d�smL� �7l�n�Y3��9�0	��2�Y���x��1�jQ�P�b�<ʰ��$����O��6rnQm滨�x.�:���4s����HbG|��z{#��ǝZ��S�(dM�s��H�I���VJ�J�K�ъ
@{&�hY����f:�3�9u��㪣��z�c}wχ8#6q�P�/aP,���s��� ׃.ܬ���e�i���k`��ӝ�;/vK��C���94ös�,9X�;{¹ 0l���_�=Ӫ^�^��q��oS:��=�{��QX�)�{}Ǻ��m��|�ۥ�z&��)S���R�6C�jݤ��*|0~�]�2v�;E�%X�b�)a�Dq�¶��*�=�(�w���k��}rR�rcIYXi�j�ŒL-6A�;q���΍��!|�����k�f\G���X��qj�o5u��b�z#�����z-���%��Y�xg�k���i�*���16Uv2�K�E��W�}�3�N��g��/j=�N@�p�1�x��ά]�P04����)�o�,p82qQ��D{	s	�ftdi>mJ��ǰģ��R��W�O{����
��D8�>I��u��2E�C�m;�i���9HQ:�־u��5��Ս*�PYVu��^��:8B5( �gSNn`�A��Et�u�9�$�k<��;EEx�h�P>Ot����R����{x[ʔ�����%k���-���=T%_�LCd��;�ee!��E�<ȅ �b��El�u��Z�#�j
�uwv�YM�@FSrI/�wy�u��Wt�i2Ѹ+���:⩵%�g��()t�K&|mqĆ��U�]���Z�D�HB�.t7��d����ȹ5o���ۂP�'ֵۭ��񛫵i׽���s|�KEwY��,�u�K���ھ�#�"�b�&�W�n��Z(q�l����i�МSf�� �6nց ��BbY�9lYe��Y[���fX�D�M>-Gۀ�Ԗ�����3�����\A�� ڽ��3kH-��fG��b
�[��d؇&�+Z�n��Yo�,��PGoh�����f�g�U�+��5(~.���P�r�x�4��4]$Kn��vv�5�Vƚ��C�V�����7�����X�ik�̘�P��s,70�֕+gY��[�kU�+-�tU\�yG�� �_��K8^
FޔfNױ��|iЭ�QU����}I�ψu�n��b�u�
X�뉭(��-f]GN��`XF�ְ3<�;��8�p�� 8C|
Y�{���U�_+=���)�Y��ۖ�iةJ�%ש��DV����4�k�e's�#G�9tR�8:�e��Wݓ�L���p`�d�us�X����z�
EV��:E,_q�U
�{���r��m�W�伾<:Cvk:�+�F���ܶP�wV����җo]dI�j�{��R��D���Ң=r�Yջ�h�ow'������:�-=�)c\WotZJ®����D����uF�8{$�x��GC[CrZ�� #u����z��F%���[�ʾ\��"��k�+�^ܼ�hպ�K0���1!L4�sM/���6�w�,��V�n�я@��fW#�������4[.�\�1�=����r�Z�޽ԅ�;���&��tr��ÞtΌ��ъY�s��%��C���:2�}��C+,�s��I�,
�]�*ދ�Yp�MY���Q�Y�f��v�vٖD�Z�{,1v�5��m	ΟHKM�˔8��.N���7Y�L�vEh�_B�m^e�S�Ԭ�r�W�mV
�2��Nc�p��R\~�;���p����E9�T�`9{��b�Z*ec���B���N�전� ]�]��GG0麔i��O%\���8�=]��/R����++;�VG�T�.�xk��(�B�Z�"��x��M#5�\�̺#8�a�y]�H�,S�*��u�x{�g�7��C5X?3,Lw7P��IT\
_@��Dn.�U��(Np��݃5�C�uf��+�sΡ���l��C���nM����h;�%�4 �YZ�W%@�MS͗�!�;[��5ճ(��w���q\�8,�C�9�Ğ�A�h�@��t��v�D�PСZ��$/Î�e.D��n]�ߺ�c��{xpL��
�w���$Z{�忎�.�]�xԿ���/�������B]��m�R��Ma�c��;+G"oIwݹR i�#�E&�pe��^$Rʗ�,:��}j���w.�z��B>:3���Gu�b�ol�1�˖�1����p9�c"a��K�҂ʶ0����r��҅�ԩ�(s|�k"�,�O��S6����Κ�m�΃
�m�{�Dz����q¨���qw:R,��L�t�pTu���QZ�i�KO�wEX���4�����f��r�Fr4{3��l�����b�U�w]h��oc�`b��u�v�J��٥��4Q)� �@r�YM*C׬C+��E�{l���k�Q��˛7�p'��89��M�{yӬ����'T�U�=*5=XZ�5gv�4��G��6��8�Fl*V����n�E���w��\�S��N
�| ��H�
�+���Xr.ਫ਼"ɂ�Cn�1����xb�Xr�]`COnl�wmcG��{6�2u�j������B�r�'�ƍ٣��0�0ffo�����`�`���f����&�� ���F�D����$䍷�\tw@���GO����M*�6GN<�̏u`��n^2&�]��$�];]��b�Z�;�:�R~y:�^�m�,��%H��c�kI��@X�mΥ|�C׺4	3]�r/փ��ZC��=������]R��f:�J�iw"�;�����.*Q��]j���;x����7+Tf�I��5G3q޷���G�t\���u�j����\�u�i�q��� �/UNfӬQ=X-�C|��l���qb�{�w�J'i��;���be1�=|/��'u'����6ʌ����u�,�*�ڟ�A�+���{�v��}E��u��_��F&�du�\�#K!Lr��jdU�8L�帯v�v�pW;�gy��C�2��|rٳ��*6�Svm�C��-����עP�{NNk�@@��!�h8/���H�ˬ{2�*�t�C���<�]�MsM�B�
)�1g�`{Zu��.�g��
��V�W	�kNpv�E^�<�+��6H���9V�f^�.ʄ1��$���wc�r��`Sܘ����̒��\l��lM�LΌ��gf�Υ:i���ʳs�"]s5�jt�	�'�I������N��	���ZSz�D����'�ۯ�NˑnG��G%��Q�;S��Ϝc�u�um�][/�!�VS�eP�:<�v��y�ލh�Y�=]U��&(��0`�70�}�e����^��jh��n�.�	��4��b�:Rs��N�Mq�o�c�$q�d|t��Vp|F�v��9��V���;�K ,��ӝ���[�Ԯ�l�=��C"�����q�����<�������Ye{�[�h+e����o����*��@=��v��9��%{��<�
�hH��:+Ee��|����/ hg�u�25��_�"����������ۙyCz/(��$�U�q8���\���3�U��:��J��+b��7�daVN,�{�y�I{^���Y[G�(���Z��]�S���|����H(oeѪAڼy��"�R��bT7�֯y�x�ލ�C��yOC�S��{)�ŵ�3�+�܀~\3 �T�b�9m;�-r��v���(������%P��=�~[�{�Ǵ&9�B��n=�:�Y�8ף��Z��$@�P�3��f�=oge^S<�w?^��g)j><�"��z�7���@�7���
Q�r-,]Y��=+o"��Ya9fQ�&��?�Д���	m�ѳ[s51k(�:.�R<��3��k�H�V�l[i��������H�9\�ʭ���ub�������3R���M�<��J�8۵k�	L�ۮo(��4��\��]��cU:<g@���1<Fdz�{�3 ��~��1Pn2��G�7J�85���o��P�����F��������^�ݶ��Ц�����pѕ��ހ��*��c�k��Y�Ob�W�8���!vЛ����w���K�/L]!o��p��9(t�����c�c�Z�`�%wf%�̐�8r�� ����+����&�[�}�k��<{Fsք�.�ȸ]�Rt�n@���[vrÙ��}��;iX5+�M�P� �ph؇���r��1^��X]�/��N*�{�97��R;�0yO�dqx�=37�eq5�#��t:��u�C}�O:�G_	vE�R���m������L�֛9���.�r�P������q��\�.�i�\�I����.�w�+g���ơ6�|�<�p�#_���]Rs�������v�r`��#8ӥG�
p������nG8����LkB<�W��W�f�z��E>-)�<4���\�qp���	��ȁ��P��`�L�s�,C	� K�ܲ;O����"�
^,hs����[m��;7�@�ú�d��x���o���g��.�h<8-����ܛ��o�ھ�64@#��v��y��^��G��/�~x�N��ݼ���x����9������Iw���,yr���>XQ�����~� i�Ԇ$q�}nе3�r��LW1	��sω^M�l�ZhV��YBu�(3ٞ���щ�;�8_=�w�K%��\I�����^���p���y`�1�&/�����r֋�~]O�����;k�K���n��z���h:1����=�5��m�?a�'��=�f[��u�rζ.��l�VޟJ0����wԣ{�y!d����v芍̀,��b���E[�R��Gvc�o�g����j�77z���.�K+�'�eg9���*J�G�+�B/4I˝]{ݒl}C�	��]��go	�O+�����R��;�,�7���F��Q�&k�Tv����0a�5�s�S\�5&��1<�A��J4t�ΡZ$O��1��pB��*up�K�q�t`Si��U���x����3Sh���wI�����Gk��YX]������{e�˝��qv`��T�?W�{�nie�ۋ{���n{|$�7�Jhޫ�~P��������R�}�+о�V,�ǹ�Õ5��ȲZYY�i�u��)��¦��X�^��N
����~�LM��%�b�5������5��b����tR
���X�޾�.��A����P~�{i{���2Ӓ��	���s�Ք��ݳj�9��y�g��{K��/E����:�w{��^���|���Ȣ��L9�_�R�;��|������َ蝉{ʽ��W\�GX~��֒>�V���j�� ӥ=�􎙇�T�df�/��r��3`�s���t��u�\�Gπ*���V5������S/�=�ِ�ecTmb��*N�o�i��۰:��
옲{R��ǜ�6�צ�=��wuvp8sY���.��}�*�gT;is��W�E��I����K ����|A���$���ݺ�m�, 9�=o$�����h���h�В��T���s������ܿ��6@�(7�j6��4�ͶwfR�����;��7�Ӏ軷C+�k.C���J
n�(��rvL�8E[��^Ь�O��׫˟����v���E�w�m��])��!zֻM�v���dFLx�?tq����<��[��)�����o-�o��/3��}�_J/���?k�m�9yx-~S��Wg{�ͩd<�;��wHe=�(υ�!�Ȼin>���5��n�3��2*��hzr|��¢��Q��۩]��g�<`>�j�;3���/{��^�c��|��a�J��o!4+(���(&����U�c3`�K��(�}�9H=��Op�v����n�p��o_���~���^�\�l��5�L2�f������2r��G�N�T=��H�ݝ~�Y�'?;E��_E����w��{�0��u:�����H�eə;(v���5�6��u�s�+���Sj42�j���8�q�8&�/ne�r�TM�7БԎN��B#�H$��/�w^_)�f�=�մ�+8�o'9y��.�D���5m5�kG��`,��w� s���P��"{b$�����y�/���ي�[�GCf��,+Gel��]+ES�@��z�e�1��mX��ܭ�G�:�#t��_�\s�OE�o���F~����cl�o�R	��0�����&xi�-�ٻlm4�)2��1�
��ԧ�O����(m�-�?Ko�[�X�~YP�d-�r^O'�vIli�\+V�#}C�Y�~�G��I���h����K��N�~\�5@��w78�=�JSׯ� 8����g�K6����Y���vlYG��[!%��U8}�FϜ���*{xG�t\v;�3`t��7�֙G�Ϳcc�x]�*냭N�է�F��~�OR�Iv��D���^�>�Q�9*���������W��mЩ����K�t�3�>�T���xz.5m{�������Y�{y�߲Y�#qt���eɵ����X[���R�ݮ�|�;�t�����2��'���u�X�yf�E�W�E�����o(���c;��z\:LFj�j�U%G�۰�{�I
�Y�Vrd-���&�gwHˏ��).�{\1���_Ǎ`��u�dx�t��vJ��P��fԮ�K�r's:8/8���=<gNZ��X��We��Bm�2���\�;o�c��ꃗe��v�|`��u�4�w���k甯E��v�.X�e�M�iˌ�|�\^��wG��&������߲��=o���f�oS�twm��݂u�א�5�u���y,�.�F�8��՜]_�r[�=�.y2N ��W=�d�W�\�T�"��,��#|��Ϊ#��gG�\AU���+���,C�Z� ��n���~[6;&1u��57U����;k��=-p��of�:�@��u;��Ѻ2}Q���Pj��+óQ�^�uK��n������cy�rk�2�He��������.�߷�Հ���kۓ�������/e��^� �kS�1΃����K<��p�ʅ��.�'��Ĵ�sظ{���gS��w6�����٩�=�[���U����2��ӏ�v]'��盡����e?\w3k�o$���.�*�!:��*i �G��*dm#��\n��6៮�i����h/4�4V��|k/R;ұ��� ��Jy�d�IG!�7R��~n�A������U�=>>�ցVi!l*�pn�<h�x�GPk�6�Ӧ��V<\Lm�����7�����;��Ż����-f�S�N�Wӽ��3���`tIyׇ�8Z&���+��`��ߵ�MM_�4�?o_�s��w�<V3K��w�l�b��!����qp~�J�]��Y3�L���_N���ã�wIbU��:l�E�o�&rˣ�m��I�o����n{t�jZ����5e���<��O��	��9���u��z�U{|��qX���){^ s�Ma���c��]��z�z ��c�1������Mf��k�o=Lz02=5=8*��x����w_�m̵y���{���;v�,�_���]y5������.�z��
�]n`��6Ί��o��Κ��V��^e��j�g��t������8|�=^�*Sw���q���^�
y��+]%֧6����(V��<�Ç�($��
l=����5��j��R�V!�@��F�z�ɲu]M�4��HF�PƊm�����.�(`�<*-Id�hK��M�5�Y�n��_*8���$N�����8��i<[[�q�k����o�6̼��Y ]��OS�+:Y�7�m�Վ��EY���&s�q�]����W5^֯՞�v�̊���[(z���?�R�ia��k��ٶ��m[��"�jS��碡�s.��a�=����^�E�kB�2a�LX�=�z��FY���tˡ�k�oMA�����]Q�9�n��P}Sf�ԚMh���\��K��Ļʎ�۬���b�f�6�j��N��և4�������GyG������(a��w[�����Uk��wL* 1�ۿ~�Y�c�e�Cd_���`�Z���I2��|yQ����]5����g=��K�!W�Gl?x*�>���z������m��ީ
޷��������o4\���C~��"��ƣ���&=�w��ѻ��D�1��]���M��f�$=羞� �_o!*4GeuR��A�e��Ht8R�������{���-�A�F4���=�Fu��u>�H��W�2���~s5b��z���V�J�u�4�&lYslֈ�u+f=��9X��T�Nw[�_#�.�Z��a|G]��u����wa�1\�`_<���uܸM�*n�	l|#��s�r�*�՛���M�}6���[2�Q�j����vNZ�	�Z]^<Y��E�MV��F�T��*�7����
{r[�^�yZ%�L*��jut�gi^
�2�������{!��{�}X��x�C��y~�|i�ī���c���
�`v5*]��D�Z��ʫsټ���Wk�黐�⮅>�H�>��!f���3:�zW$�O(�	;Ɣ6x�B�E�.
l<=_�wH����{�nbx�G��Ru:��1[�sb���]6��3ך�[d���+�����\�N�"҇8����<{��@����
���{V�,i?d5��ؼ��a��[z�\�}��l�w��g�B�G�z߳�@�,�yW�s�e�N�3�T�?
��J7���M�orcꏭ��pz�Y��<��.��KGD��}�N�A��K[�/w���]+�ud�s������:=�٢�x�2gꢿ]��W�aՐ���������j��(P��(��:�{d<�ʐI�����=2����8JA8��4N�6H�8?#�nR<^�#y��WX8A���W����6�ͺv�m��8�kw�<�o]qS��WKU���i¬����,�_,ݩ%歬���`��rmt��(!W����I/������v���2�-LAאڤ�_t�W�ƨ�fg8?>\��AUĥf��5�x�НY`��d�2�&Vf�Q�� ��N��������^kt��=�%�hfi#1����f�w��4�=9������0I��]Bҙ��.�]y|�v�m���)��8\��w�R��sãQaVL�6�R�`]��|��n���5�ȏ'ov-�[�������#`7õ�c8�4�I[c��#I�Z��o���ѫ-��Y���v��ڝ�k˃n��[�fkڶRT�hl��E`�V���\�1V� �ֺ��aj&m�+/`&�������!imA�-�8�"�����y@�el쒇6E88ው.�Z������u�]���������%؇�5�9h����M���'W�䃅i��y���M�}ٸQl-
]��F���,wK7˳� ��(�	�	�5���p�����p�hfe^�Ts 䌧\uwG���8���z�(�(�oA�-�N��WjVε���k;��)=A\ۻ9��^�r��+�B��[�.ٸ�>Z����2l���'��h��r�% X3N�5��:�;�L��7������$��|g>ݜ��Ƴ���]�]:I%F�[�Ak���9n�yz�vsԷ�-�U��@��xs����[��b=:B��A+\`���d<���4g,��)��|I�
�y)�%]��˚��6��ZǺ1��*�e��������C%<��8�QF�u�M$�;�}�w^_�~b�~���X�+i��s3@�]9�����=��K��^P�2����JҦ�F����]}V�i����0n�E��r���p_��+���3)$���X�1�� ŶF�8��]�.t���O\�iT��aH�t6 vif���^��J�et�u�&;J0Ed�c+�c+�v�_N����Q �~�х����/B��wk޾��>�nek�B��3:�8S;�_4�­�M^9�gW�b���ʖ�[���M]ٳ���:�"y��Ŷz�*��w�2����L�F:m'9����h���a��w�3uS,K'k�Km�<�ӱyh0�W	��m�ګHrAk�儑����u���I�N���dر-ؕ�ok�坨�%�)m��ʞU�]o����
����ڳW�J��&;�F����+i����1�=�pob|N�V�B��ч�f_T�*��b��S�;m���w�w���)���l4�̦��v����J�eիKmmV�m:}�X���Vq�q�ȎF���MNΛw��d�x[�w�v�V��� �~�I��+r>����苈��+�Ә��`���җPO���h��v�vu�
���h]Ev����&�w��󅻸�|��S1L{�Nv���9$x:���*�4�z�]��z�������~�ܒ�wq�1ok��ì������{~���,��c@���:�ُ�e}����V}-�Z���ִ�c�'�K�;A��W��u��VTI��#+#��p_���N�r�i�ZW��ߣ���B��R��e��,��]*�2�2z�(0]<v$=�~b����
sg9�ъ�@F�.�"�y��)=���
E�b��[�%�Jꪽ�����ۢ�m���.+oP��=䇏���H�pe�>�nu�����Ӵ5���mf�[�A�:#nݫ�Hs�Y��<�1�)FEk���AJ�;�� T��ǰ�9�H���_A��}��VK�r��0�T����yiUA-�^�Ӌ��k��
��j������=�3_x��6Fث�
�]���z���juf��N����V+;�ݥ�^��]�����WP��<>�yw!~v2e�5�[��7�;q������
�^���Q�=�`<�h�W�t�j�<	i��.�L�s(��E@֬�j4z�h�WVz�t�|͘WZ��N��S����X��W�?f�R�	:>޽�\��Mۭ:2�!ƹ�Xն��3x��5�]ڭ��em[K�׃N�v���*]�U�y�γ��qu5��io��WR}zhDZ}��\�H�EF/pX�u<ܸDa�3v8P=�DoFԐ�����S�^�򹊎���k�Oss����ԗ���:b�7%u~u��l�ؓ�YV��Lo�sT�b[#ѿySDu�/�\,�*��>v�zrr����S�;@%Ie}��!�r�{F}.��x^�/|�p�0Z5:Z�ۓj���P��}�?���V
?{ZVq���-�W�<�w�ff��[�
5���2ch/E�f/��,93���&P�'fl���b:k��>2Mp�K�&����;3潴.�����߆d��;�0�{�W�Ɵi$t�}k����E=������ث��h%�e��?6qY^3���Nu��g��݌�t�?1cvi׌�X�f�'�h-�ب���U�<��OHs�~Q��_���u�5��,i��xK|qu��'�ɡ���vOxY㘬N�h��?S��2Ϛ\,g�9���|Ν]~�����ޞs ��#)e�8�E��.7�h�?k���d�i4A�.��oXz��ř������ܳ|��CbL/Br�J25�>���&�ɯ4u��P� ���<R�.��i��ʬ��2u��^Z�k;MoLeud�鑋
/�k-3��=����d'R�3����ow�6�
<e��̡CH:s*n�y,4��fRKiU�V�.������[Ĺ��n^T�j#H<M��0�,A�3�D	-)���G6�L�$5����=��rs )0��Y�#$Y����:�T(ң&�.�U�n� �̋	H4e���v-�����l�׆oQ!�������iC2,�!�dCq���dF����"���$�!�W{��B��5qG$�<�k�i<�Y�i iaz��QC#���%��ɀ%�����Y��4�И�4�N�#`�Qa�4�2 �秲�2��>��X9Cq�9w��**�����ۀ��T�6GT�(^x
��n�$j�>4-Te�Sڪɴr���v�C6_�x�ژ��<��[渝�Գ��QEL��Q�%���x���`���R�5!ＳWk���A�y��^L���2�����GE멟���� [޺"o�Lrg�:�i�)Tp�/��م�{���/+�	R2�����fС�8��eq��eg�f�G�wv��=��S��;>&�s$�V��#�g ��i�}����kf�֝���0|"�}�&��9�%���Ka�v�<��.nMŲJ=���+��k��6�m|-�w�_��G�c�ξ�L��{���W&S懋ϲ<C�\}���/|D>���@�9���m������F�,�$��]�7�X\��Z�������#b�� �u�<4M�36]i@Dj˻/@Z�� `Yz�!�@��?9&�F�sZ%�G[���F�.WϦa Y.u�d)ד���.���-����7��)�t▎�Hɔ��ð�dJ�8Qצ�諎?Öf>=�>�մ(�ܞ00�����^:��y'���y�f���:�w��o�R��G��쎌lk�⇼޼��Ohaƛ����)r]
��:s�2��}���2G�y����-}/}��h��s�"��s�����]�έ�Q�~[ƾ��<�^��Fٕ��S�Gզ������A_�{���f�UE�STX�_�mw!�~��;��F~��p�]��ڝ�Ok���_v�DO�|)S�d����~|F�+>.���v���X����=~�Փ���yW�����W|=�߷�[ \X�A3�bϛ�5��:��W�[B8'S*�S����m/!�h��]Tǅ.M�(//aЫq|� �l�z	�D����	$F�;ʇ*��ClM�>0�a��n�t>�^v-����Wo����!�z��'ƼEve>�z��_��L�Qp*���z��%\:�mBߒ�����y�꾄*������$\�b��s�gq��糲�c7كD��H��������!FM���y��]���a����]�՞6���I�dl̆~ôSTv�տf�w�˔����!��7&`��u��Ӛ����gY�(�n���J��D6����aJ�� öa�i΋��벴M�P�|��eg!�:�{:��O/GZ�ww��V�g��VVo�d6��MO$|�6!�1�^�Mɉ���J���'v�1�e��K���f��{����xg+�3�\�h�W�W5CW�u�������z&a���<R�?zo�f�G\[گNS�&��lO;n�>G��|nй�ؕ�EQ8��Q����)H1^P�4�^�sw+�7v��'���.��W辇��H��ǋ���f7��z���t/��]�^�B�C�K)�E}R!8�7����c�l���k����w� '����6e��x�uXY7�<h��f�^�ئ��^�菪A��Z˘�÷( �d��^���'<�N��f!�>�'5w�z�H��b;ݙ���6������C�+C�����P|���Nǻƣ@̩Ԓx��F�o�H��C<�E^?%Y{ݵ<Z��p�:�3FEedӁ���P�y�S]$��"�ܭ�<��_�G}� 3�|%7{��;o�GED��2�M?p]w]T8TS�"�9�<!��-�u|ڕ�Ph�w�zU��E�rIqb��T���ͺcݣk�NJ_�nP��zw�gUvXݹ\���
�Jrz����ǅco�g��󬱚FU���mZ���z��-�?oi�أ�Iڗ�K����5s��d�_�ŕDg�9L��W����-rV�{je�\�G4���Xgca�Kz��Y[v歁�?�/z�~lӉG�nXc���&⪫�t=��}z��_�����KY~|�h�E{o[�D�ս{���^�h_:���~�	<4u�C�O��z���o	���w�st�|�۹''cl{,R�Y���O�pt����A����=�X�\IT�㕦����S�u%��YW U�t2���zs4�[.}*����^�O�烺�향���c��@���lg��fx��NA[�1'��ږ���ҳ&��\�n�sVj1� ώj��,U=��Ҹ�Z��q�wU
�;��nOuOnլ��x����/�G��Tdr�[>�\�Κ~v�������~Ѳ��Zo����=��w��;�������%`Aģ��v?MQ�_�3'��7���gf �������<�'7��:��C�Ҙ��u�o�6ed㕞G��;Mr9;�����݈=����8�nL[��. o%u�d�y�!(��#YȞ��q@���y��d� RA�	�����n�7:*�r��A�:�4���8CgPںs=ü|R�	K�����]Og��{�w��(��F;��z^p/� ����s�8R{����x���
LM�X�����*�T��]:��mxu��V��m�gVe��6����o�M|��kn�.@X�2jF�����X�o{X�gev�\��珺ҵ�k};�:��q�L�y�.�BR�E�
8��L�FpWG�ww$B|�؏���e��p�a�G�-���~��q.ftk�k؆뿡��>{Q�_�9�b8�.e���*R���ǅ����"�o7}�1���S�>�����έx��~��gI�	!��eT�.��B��;ݐj̃�I�g$����{(�i����#4^�_0���nfMz�
��j���ƻ)2���g���Ho�.f��$���o��\��7�$���8��B1gi"s+&<�z�3.��	A���{O޹�:<�1{��ea��g�7��{����	�q^���{r�Wa��3�X�qU)A(�����VT��߯��zz�x�l�n���d�|i�P��7���8K�[�}�9zn"�����z�������p��ζm{<���-Q�γ�ȋ�T����Y@��ϴ�e��_�"m�������[�S�z�zVh�{�����|�*�������Ry��F��/�kє��n	�۩�+|�d����p�_r�ƽ�������\�t.JV{s6��_ �R8��L~"�������[����Y��Y��:�����7(� ˊK��A4�I�D���\ݷ�.���w���9���1;���T|&�/_5�w1�ր�n[r�
X�#̞���g0г:[��[35q�Iu�Z�w��ވV��O{���u���߫%ݷ�O`�^D��6���Y=K�Hj7}@^��Nx��>�Q{/���5�F`�|�Hq���j�e	cB�k�kv��o��?��]�3a]�U�/�2<g�鿏9��*�~趚�^������͝�)�%5�������$�H>�^�
����k�@��Z�94�M�e�G
�5r�SŻ�Փ=�Һx;7���{y~�ò�_�|��k�|z\�ȍ��5Nd�O��T�����CӼG��{]FuAS�k�b���[%�=�"E�zV~��f�aۋ�$����R�/-����3"y�{-�EC���~�g��� R��&�������λ��;�a�y��Q�^�ֹ#�g����g�:ҟ���^�WC1�>SL�h���w����u�^S�I�ۇ�CGw�U�b��`ڵ��	��9�ׇ�O��@��9_�[�g�>�h�zw[�:��OO��X���p������]���J�]ag��[c�`B�?Bz����jGݤ&qF^(݊�cf��G�8X�Z�2��q��F���f�6��9�����{�S˕�k���N����0�ʎ9o:���3W� f�[��b���nÁ�jWp:�M�a� ���z�-Ȫlc��sa�.\���d�c
�8-څu6�DKr���w��:E>&wΒY*=~�����Q���X��k;wbTs��|7S�Gf��(��0�u&�e��O8���\�3}nbX221Z]�LGw�-�o��R�>�,P�3�~�����w����۳V2�u]@��L�`�
��1��F��L	�-��w��}��wD���<���t�hI�����1�^gz`W��.N�z+����]����i�3o��y�㿺�_*� ��yߑ�����;�c�.�{��2xT�$�fn�&���+�f;~���l:^�Z��W>�G�=����pO^��Ӟ���*�Ԣ�{'z�vo�c<0�>�^+NO'�#�<�9ϕ�f���zx�n��4�bϓ�K�����˼j�~чl�6�s��Q]�����7~6�قQӾ����~��Ŋ��(�۽ި}Y*��R�X��@Pw��n�Z�3ϋ4�i��^�;h��OuH� �ψ��ߟT������~]7yB::���zͦ�)=�J�o�`M�D����4�(*_>9f��J�56�U:
�Ω���N����n�Mє��]�D��'iT���nI�]�b�n�G&ŋ�q�����sv�&��4_������w�
�e����ab�9b��u����w%��dom����s�#��߱�_�o���_��f�'$�ζ��n��v}�%:R�̳�Px}��Ȩ?�!��0��S/�͂;�k.f�I|��q1t����ɛ��s�G�-�:���g�E�m&g�x#���hV7�CY���C|��+V�M� *+��δ$�I��]����ȋ���=��7�À����ʛ�'��Ȅ����o�	 �7���=��|��QU���9Ǹ�|9b�"v�_�-��_�Ay��w��j�T|~գc=|��"���LR3|jH���E?�v
|o9��Z��oh��,�ʼ@�1�p�d�G�{}7v��~�^B�R���Q�Q9Yz�+2{Y*4]��t����0����|�O>�#��Vu	���~",2�	_TV�uIwԥU	��opT��ykO�Q���~�F��`܉���N���՞�\��$3�M��۟���9�g�9^Ff�8O�'�`����<���K�>n�g+v0��<��˩Z�K����7R��c��ׁ�6�O��	z#��_Ϗ�3gk�m|�[����uA� ��9��W��G��Yb�eާ1�Y�J��{=�~��^	T����2�	��@ҳW[�*���P��VE$Ѣ(������s(�P�_YL�,7u���p�0�`�R�--��t�pΰb�x9C�(�����'��呪���Xќ�U�u%��ld���_pnV�WS���U��Ph�Wnh�OE-�f�_#)�T��wV�P���ɥ[x!J�Vo�=*�u�R�J��ְyi��н疞~��-*E��mvN�HN��ټ��ĳWF��訝�<h�I�e�:]�0���b�c�D�u8q��ż�Yƥ��9�Ԇko�'"95mYjuݭv�ͣ��FRl��:R� #+�ހ�X:�vp4$�*��BR��s�a8.a�����P��`5�wp��}�8�@�RZk��g�t��s\�RF�..i��W3�8{�py�D��S��N��;HO�l��txg'�=��F�|�ᨨX/xH�#�:Beon^���B��H�_-:���r|��n~�8�2�Pe�Ư(�X�G�[�]Q�GE\�\���?�E.�[�m�}�Ňh����a+9���y�|�X�Ы��7�V3�+�D�w�W�rQ�R����6��͋���L��3F�����`涋�خO��wr����ؤ�U��.���꽫;R\���/m�������P3Mjd��z��j=��%gL$ý�s�ux��@Ol�GT�8�>��\�����x^�w�2����K�娼�p��ϔ�)�}[��f9�V��G?2��.nPN�j��l�.�+�J���5L����޹�my�s��}$��$����Omb̙IIM"N���ٛ${�%�û^��f.��6�x�]ý32x��o�wr#��\3.@Kӧ&5&�X��SJ���,��E�����PZ��ʐ�GϨف�C+�k��S�`�{ �a���l�Mݴ2�_@m�aYבH2B�T�e� C�m�ػ1��Lp�&������F:�����Ui�Y�=��j��E�R�4��d)Q_S����?hBW�5�uWc|��I2�#[+MJQG�L޼��n��y�7��j�g]A2S�qM���C�C�ݮ2�yw�t���Cn�"�b��n;�6�<J�=縍ܵ%)�{�5�nI1�!�"���WO��YP��ai��F�i#[��Ke[Y6�z~ͫ�ݎ�J��y`�8�kc�N�u��ܾ��;��ޝ��?S �Q�8W�O���:k4�A�s!��֤ŬG/5.���`;�������e#Q��y��J뛔euk���9�ګ1wd�p̓%2��O���`���:��9�E=��w�֑��M�Wt��N�E��9���s���6�U��m���@E1Y��?n�"��he�H"�{(VQ+�ܡ)m�T�[[wH?�c���c��{�V�B�&fY��*w�Mi�� NŠs����gGv�c���[)����#Y'k�Y�`�w7ź�w�i׸�W��ro:�M�bի�'��N��.4k��/���#.�Qai�*7�y�� k�X��@D��q�jd�Z�S�����a�K|�wqy�8��d_�NV�-��h��Ŏ1���z�U�-��3M9V �v�/E�����>`b�fϳ0^�Qu틎'}⪬#�Z���0y�J�yN�EE
Uޑ����h!������`6:������ޤ@�N/o�n$s!��� <.�Q*�4<��?W��^Q�c��W@E]�/mL���9u�nC���D	%=���z�V�.N���L�Ǯ˪��̜V7��.(_>��!��꯬g�C���X�����s`B瑇<����W�}E�~4�캉Iܺ
�1vLI�*�Ѥ�9�ex�nz�<�2�h�I\��2��}3������o#��ޝ+�\�]$ϒ�]���Q~ԕ��>������v���i��,�jC�jNd��*�Ɇ�eG�����l����C��nK^~aҎ)���}�ex�N5Z�@oU��i_]X����g5;Q37\�ϛ��*�F����>����<���z��i�����ي��� Z�Sn�r��"/��Y> c�%	�hK�ۋ�Ԣ�!g!�
~^�j���J�|��'W1�>��M���(ySZPH���t!cd���z<�Щ�mҘ�]�i��r&2�6�w�Ş��&��{��W��|��.w�n�<o-���d��/��֧[�{G:%D�n��O�^�2Թ�>p�0�v�����hup
�w��&:Z�SGZ']EKs'3�A����[%^l��Ç:yB��剳�j�c��Μ�5xy�Ә�[��sF�Eet$g6m��`�n̷HvFͩu�$t9Υ��xm����t��N�Z�MԺ�%!��h��v�*rDz%�,j��(h'ݵ[T�I�v�"�҂���E�0Ox�|wr[��j�ﳐ�Y�na�:�GuӨ���\�����Zv���WQ*ʛ��H�ҫM�v�Yb�wr�C�}��@�ϯa&y����y����w�[�,L+io�����[���������w�*�*M��n����G)�f���y����^��"No��X c���	�y;���{�ǹ 04iOW}wZOT���k��@�7C�O=��{�xQ�|��\�
�Ʋ��}�7g��`LMDw��vM�L�����G��Jڢ��Qi��{tW�٥ԫ�f/cCf���W�'^�?��������r������5�>yT;�-�NfeύA�w��t^�U,s��7����0EC�tW�(���2ϛ�Wj����lN*�5�-=��/�Z̿<��O����S*I
�[k3��b���-[�+�w�-��B�}J��p��{�-+�u�=Bw`�Έ�C���!bʥD�9 G�l	+�?�~_���{�#����fD�9���^�	 ]j��q�GQ��Fp�N��h�^Oi��k�o�0$ו篌t�7��ɭ���a:�Q�������5L��s�zpTt���{�P��f�mX�<�}[2-�6��X�N9(��&�tV����z�U�Ηg�c:mg
����3��#�kɢ�³H��tl�<�)�M�؇(�gu�'M�b��5V��T�4U�Өs�Мu۝�������վ�a����n�+�K�e����(r����M�k����9ḽ ��ƽ�)�뻚F�/U�'>��~��.�ޕ�}�lI��I�iʙ�s��b<}u�{3G��ye@3V�N��-]%ڡ�(*^����$��N������|���[S<�,6e~�s����q�<n<B�]�.9It�Nک�%EgD7KU��%��nZ���bhG�
�$����Ds��%t`ŀ��=��/��Ou���>����H�U�*�\7l ���D��n��sv�|HQ&� �#�Ċ<T"�#.w_FW�㡛a��Tx����B�h��7�,�>�X�M������Hء�Th�v�'mUx�-����|υ�ڔ{2�1�������Dq���{2���N���{Y�����
B)kP=�=}�*^���U�.�Q5D���*	�l��߭�@u,=J�o7��FO�,�nud&�a����ِ�[�p+����GX�5V�,�"3S�ή����!�k� ~�ca��x�]Pft��[h�]z�����B�H_!K�j�[����4q�JT���� �2�*#R�T�8Q��N�+��}�*��̞@|;zl��_�i�%ݔ��|�JZqKe�X[��*�^����n�������XХ@V�u����>���>�ܢ��-K��v�+�6�+O{\��Q���|�o>у)rՆ����yx2ioEN�r��G(]T�K�g��!q_�L�ķY5<����(h���)��W���Ts����|N.�kg�L���n���0��w��'d�:��v�������\�uB���QB��wF��%V�UF��Q;WQ�ΫС� !��ϝ#ވ�UXr�8yc���I��uށ#7T$��SFy��(���������H3������!�z>����rx᩠��1}fx.�nٚ�ŭ�����%Y��)A��K����_\G~�1�_{7�si�K�M��ޗ_��W}ۗ�w���d����W���[^���?�+ϡ=�<��� ]n�}�x���\�{�0Nѹ���M��1-7�q�t3~�{^�_,�"��ҥw�ƜZ���#�#D�٘�/2�̼��ʹF�9�s1x�`�v�dH�.T-P�B�B�Lr�]#���-����X�[F���KWr��Z���_�g�ٚ|x.>��E���ry-g�Q~�f(
�����[����j����,�~P>��U��Zz2�|~�)����R��]$r��n�{M�V�h�gpp�JU��i�=�7�����8�<��I��naFiri˓�T�׻ �GY/�͋]*������i�|�5���^�i����Du��~��Y��(���=��dBr��?b�w����A#OB��L=�ؖ��Z\٭��v~o.�#ot*�[X�S�ki=Z-;�Fi(w`}{�Ր,�ŋ�m'4�i��*�L�6;'��ն.��+v��W`2�(��TZ�r�%�S������dǵ���b馟7�ছe��@s�ZSo78Z����m�5^���áD�>���`���s��m����鯡�^4EEG���$���BX!pY�B�(#����p���u�YX�hhQkC�Q(��rp��7$�^]d��G�;}���o/c�Sx�;�_F>B�G������*Ü����~�8��P̛�l!�zNM�-Ղ3����b��y��׷[�br%��K_%C�ȏuZwv�Ox�@U��E�q�lo_�b��u�����z�<��맪Y����:�=�o�'٤�n/�T]�Q��j�n�L�Xx���J^X��b���{�kҩY>�8�*qى��Y�}��-�x����v8��3��KaFQ���~7ѱfU�]>�b}������o��E�V�Ew*��+��D�h�ztTeJF�;��dm.}��<W�L{3.���6߽f�����c<���T��&�ͻ�i��+��YX�.�%�ܧT�îף�\�J8U���Aݬ�r-ɂ��;�O�ܶ����,��������}�d��Lto�D��=G?z��S۴~��x��D�^N/	��z3���^�!Ò7�����˹bv2=^����)cv|/˩����a��;�^G;S�`��<�]8 �
w�Kz��\�0�Ĳm\�ima���'*�V9J�O�O}J�nH����Ip��T�k��ȲVh2��^����{����1H�(��!շ�M�Mʼ]�{G�]L��3/t�&�v}�^gV�ʫMﯣ��j��s"��l��_D�b�B^`q�X��t��O�7��T�����n&�N�Opq���rs���*�ʎQ��o�Nirt�ݶ�y/�D�� i��#�8���%��d?n����Ihb�*�vo=��:����]Qr���7z5LE��"}���N����pd�^jb]�T� �I���pDQ��ct�^�픠�Rr6�wSsN�BLE��H�?*2�c��B��=Þ���9꩹���T�}��e���@1�z�����1�x��+ނ�S���.\ϥ�D�&��c{�)Н��Nh.�p��Bo]"�D�wS���gYј�]U�]�̴�O{�	sS�^����w&���;'���}��Q׉O���������vК��n�he��1�*~WF@�P��y����eĎ
�\`
s�.3���U��Tkx|ឝ? ���r�>����:�D��^a�i���$lVN'w+{Q1R�tؕ2�����<�=33��1F����b��~J�P��yYħ��f�\���&����1�7���*��y�	d�u}�Z��k< �_��|Zt����P���P�)�B��}���*F�2���|�.Lur�a�v\�|^��0�ҫ-�7i+�p�x����
�;���o�롆D�,������;|-��h�w�]��ت�
C�د(�R��z���u�#�Y�to�M�O�x27}\a�"����y��뽼�s���XH�`�C�v߅/��$��:�*SA��Δ�d�$+,Fу@Xj�^��z��_N������t�^��8�2�W��V�rɒ����Cu�iw���%6����Ȏ����:A�J�-�jئ�a,~�X���Cs�w�6<�ɜB^��Iw%�L��h��w�*���)�R�
��ë.�ɽ|������n�tci�0]F��F��b�}�m@����V����:����}��
���P>���������-�+W��n#�G����*ud�v:ٺ(O�����PZ����}i\^G&M��ޚ]9;��>�n�p�g6�&�w�*�Q�jJCi��*�:�J�uz�PW��o���6�X��uA��̆w���?^^L���/cQy�W�C:T��a�/��_rhn�w�k�b�'#��
�Rs��	��ex���w8�$jɩ�b-�N��F#Am�2@x��z�6�v}V���}�}�>Y"$T�����}��"{��B
7Ƹ�s�����Lq�OG��uț�d�s��yB�<�Z�u&��
���R�ƭ��yJG���<���璳~e٬ժ�����ty�S�b�E�^"E7L�t/y�c���&����o	%�(ɉ�+�0͍c7���s�qVVa�::|gq� ��o��|x���9��~��r[yz��Fܶ�؏�+Me�2n�=�m�)��.�)L*�GXT+��\�u�qL����?��;w6�)P1�j�+%s�]p�WH��D����ѲaU2Ta�&'is�&��.��{�l�N�>{$��r=��A��e���F8�:	�����=7'19'�{�����{�\�V|[���O��",�0ly5�{��aB��Ot��b�
���ػ�{�K^y�SW�ƟHdiJ��Q}���}w��4"���V�$�SC�`�zڸ���PUJ�n����'�{� /&��%���-j���r��̪[8�+�������V��*!���\G��n<�byQ�̔k쵻�M��-,}����hG��ք �6��/8A�1�����6���ey�_�=��xs��D��QJ/�Ͻ��=���yb�uȰ�/����$�&<�⣃sF�Pq�ِ��;d*�2�^�#.���"�qѿV��̲�o�p�*�����/�R�K����炼�P�8sxg����^yinE�m��@�ٗL��-�''&8|5������O�����Ҫ�G����k�����-��}U��{��<��f��p���W��1:�~�����e`���/��k�T�=��/�A�v���2�%-�Rv'Yb�,8�G�XOu������2��/z�ǚq�en,~[*l��tO�u���cu�Q���y��;�Q�v����qWKb���5�\�L�g/��of��,n�kX�{�����,��C
�8O�<k(�h	�����/}�jfa_p���g�uY�\)Ȱ�m�߄��Q�J4:���|��u��]}���u��e`�_L�*��x��Ϟ� ��Bz�:�R<�
�6l;����<�}�	���n|ӰY�m-�w/�R��3�'�B��bSP�}��>�P��z�~���rd������{>��k��*A�]!]o�EJ�³��f��tx<^S��$�=�������瀈ǂp�2��以R�3ʳ�>};��T��pj�t�X�#'�����"o�ҕ���1ٽ������n}���ɺ&�a��{��N�CD�]�`�+���5]U�=q^|k<+M)ɬw�K�`Ϣ|�y�1�e�h��>S���z����b�?Wۚ�Xn��B$�����Hv���a���ae�O�_N�����h/����U�֨=��F|^���G�ڡQ4ѳ�K�Ý^�5\��}�X�V*v�jZ��\�LG���k�M�}��+s[gi2lJ�8F<���W��]�h%�u��*_yۦ`V�Y;�鸪��K�U�{��>lr�]�qY]�Y��2}R!K��Qn�̱�N�q��>�����uU���o>��Q�B��S-�}�,���żjnt��J��J���'����l�X�d�m͡f�d)��법K�uk�-f[�xQ{nog`��Z&҇����w};�S���;��q����զ�m����L�8�7�j�ή��A�f�� ���g9.mF��{ ��2 |j��1T��<��J��#��*s���Pz$�>��6���+�#�ך�[���6�M���W���cv�zW"=��S���ڋ�N�f��܊dK�����Fue�Y�p{��qb^i�l뷱c-h�����-�/�������|�.��C���[�3N�Ϋ3�v����}�.p9l��$�˒@�p�w}}È�L}s��Ws"�)�>_
�:�p�!�SM�צ��q�ߝ���w����ڔ-�=^�|���F�S��拵?`��N# ����x�C�wF�̛�^;�^JFG`@�M����{}��^�'�*�BӾU���şH�q��R���[�{��_�ـ�\�����]H��v�sv��J��/$5%mS�q3V�L���.C�?'�j�?0M�B�u_l�z��ӗ��'��%�ձn�^��{��>q�2�˩bk�yG�@̇�GEGa�g/�Q�ތ�Q!R��Z(v�r�QL�@��B���lm�3Y9BO\��d�8�]qIź'�"��Z�ۡ�}���0U��"E+�I*����ԵW�|����rx����+�ᙁ7�=^{�>U�̅�C�B�y�vö�����P�&��Q=��mtx��I1�*����k]�>ঊ�{������:�C��[��w���f�iT�Hv��T��̏�+�;��v�[37�d>)a9|FV.%Ú� 1�a%��NvL÷֙�4���="�����<���FR=�ۼ�ljI���Ö�Z�E4e2x�����TD��4
��}��lս���39��q�5��e��9z�q�#�X֝��z��^}H��!��)Xo��@�CCXv�6$�
�r�S�cJ�V�i�:j�=p��C�"���eRoJ!��U�����r`��+�C����y�=.�����G4�W7NMW'JY�A[Qu�"�j�V�hu�6�n����v4�w4��G@V[��Xx������tfP)SA���#�f�}v�[�RJE��w�,�r����8�U�����6w�i�[���$�J�6��t83�mn[�G/$Y�tV���1��@Ů��XҸ@®�yXݩձO�읖��o�R�'��F=���N�]�n٤rҲ��dlڳ�D�/]��	��k�4�t冲��#��_E��l� Y1r����N~���+�:F��Y�����({/�"�sNܾ\`����e�Ќb��*N���ʉl�aohY�WqVK�Í�5��]#�@YY�B!��\d]�zp�rG��lnM�/n*l,*���?5+�������d�6��]k�s��fU��/���3S#�w��&����gd�̛�{q�ň�tY�=$�Ы���#�o�����t�y�����r�uͺn������z��M� �5�[��z��e]*D`���Y�R|5ĔS������l�w��ї�eR)ƣ풅i�w"��lVv<LșZ�/�M;���9�Wr$uG�7__1Rb�z���vZ��$T�Sŕ�cDT�>r���&=�d�J�	��pJYd��	NޥJ�c�u��^s�3xS�#!���^쾱 �c�2��.ŋα:K��^�����z�:u��*]}�+�;+V�Z�7�U�{ WCEfa�X����Z��y�9sF�򬳝�Eq<+7�8�R�gs�lQ ���V�]ͩ�З�5��ܜ�kv&��.;Wr���U���\�U�wX�D�x�e���$�}}����Hsה��RX
Yi���4�c�q�o,��/�/z�=�r��H¸!�/FׯC{>�p*���>�-p�zqm���f$��%v�$��+y#�Rs�(��]����L��zv�yo��7��Eq�z���-\�SA�mi��*u�Rf��^��:�c�ei�6���{����=tF��.���α��(���M���O<��ؓ�ՒȶX�f�B�u����xf�ݺc�36��B@�wk�e_ds�Ǚ��׽�8AÔG]�L�Ճ,�y�Rw�5T�X-������6�]�c�ř���C�}��v��� Ee�v��Q}��\��V�e2�u��b3;c��y�c��|�m5V]!݅붯iv������ė\w{�x����y'�o1t4FG�ׅ����̓[��sB�̙���N�Q����t�T�=����>8i~C������R�T�e��T/�0"Ϫ�'Ϧ&����C˴�9[t�֚}��/KW��ߧ��lF+��31�T�|����5�#t�@�;����A�GƜL�ۦ(�	�dl ����}W"E2gr�t�����.��~�FͬƘL5���cb���t�O��H9L���{d���Vצ?���yvd��v��5kH����q���%4�&\y��-����ۮ���A��>
���U�O�]T�D�ub���dmA|"�p� I����t����pnig��_���O�z1��蒶:��ѯp6��f������רЛ�IK��g'K���Tg:�x��>�ʝ��t�nJ���캛�jHj,e�Ջ�6�$������/z`q�x3�'b6e�2���b��wW^�)�z�p(+�ǬJ���/y:�a�p�=�����\Y�z-f� (	��C�p���BF�b��X�	�Uޕ}�}(/���޼�~��k;MA�=�YC�՜+�.dgcЫer��]���]WxU8#&���ޥf�܎AdҘ��$�Ye�ڃ���.K���>���k%W���m%Os�v�1��1]�Gyg�mݻM�Z�wU��cΈ	mb�D.Y.sphD5:A]���6��,���MX4L�ֺ�|h[b�t��x7�tv-��K7����a[�wV8ٚ����M��˩ܵ-�N���r^N(s3}G［q�Z�:s����Ug�a W��(1��ʺ�ِ��"��0U��סϝ��N��o�0nL��B��1��/�Cⵦ��o�*�}ѳ~���"}�k��}��T�n��R}�l�[s�4���⧖�~�{΄G��O���>�=�w}U>�j<;!I� �W��ah.�Z!���#��g�k#ƣ�e�js�\S�4�r���]�f��^ʑ���"�މ��7`z�	�Hߠ�_*I�釳yf�D������Έ9z^E�	�W޲�����&�8I>�
��L]ad�6��W�8՟# P�"��Q�ɿ-��;?1�o����:�����K�/��ҩ���	�'j�gi�B�S"I��E�{��P�z�����Q�;]��3���A�~C�N�k9���=�QoƧf(����v���1�+u��鉪�M3� ������K~]]b�^5t�� �%{�o$j�:�W%/��x�1Qܟ�X�^�ଫ�Ud�݂�[�eL�F�(�4>�?.���uvr�+#/˦ײƺ�к�=�Rǘ|w���S'q���hR���:�;%`�֭�h�O�o֔�����u��G���KS��-\!�n�ځ����N�K�r�}��u$"�Z�Ed뢫b���Oܲ��ʹ��p4�spM��_m������m��p�{ծT��uH��?*��v��f%ڹ^�)[ԕE�6����p�kU�(�r!�<�w���A��)��W8�ߛCH%jg*#n���>o|��z���k��|�)���О���U<Ớ�SJ g`dޝ<�6̅�*�%�%��y���J�����o�r3C~U;�g�oF���"�}[(fO0O(�r����K�`�|�[�)�U^i��b�#Ⱥ����PA�Ir�%��զ=w�𞻌��񼭡1�N�:��ܪ�	󩇗�>��5c>1��u3V��º�3����X�7���t,�æ3P8��	˩�n�H��k0�Ğ��kԱ�I�9oVLX���x-��[d�6�tp��R�c�x��ɿm��6�'�)���Ø�E
=�K�[�s�)+��^��o�[�4���R��/З:����1}�r�w��r4������=�*Q��ץm�v���{j�f���P��{�$��gy��~Yq�������@uޣԨJj��3k$
���C�.�h�)Osl�]�
]{�;��[q_ͽoU��.�*ƌ�=>BUj�� �5[�
~��-����T�n`fm0w���m�)�)M������]e��Z���q���y���A��N��8�C��4��G�^c��Qո�,�?NHǷx*b	o�,�M�p:͸�</̈́�L��kU���9��;���ue�LrGj�V��ڵ�5��x�%˻I��l�i�󐍉u3�m
ۑ��Z.����]�`���~t��;̑���׎�cgj�O�+'R���O|�f�w����X&�U�s�5�Sn���J���u�2��ɹ����7�.z�W�enf�Pw��c�U����~E�U
�;=�]�$M��(���|��@]��/�,��J��k�E�x�z;.�n&�r��y��G�g��W4�	��<��]R��lt��?@?Km�o�9�v֯@=��	x0��F�'s�\J���
Zk6�-�]�P��/Z2k|G�;�y��vA�#:��w��(��o�q'3'4O]�q��G�d�֝�r�ǧc���c �W�c�P����!��^��B�d[���Pt�Q�wǴk[9{}��>ٻ�ϸ�S���V�{I*�hw���uH�HA�S�-���k��3�}p�n�+�ZN��~����C�i��P�w3�PW��6}�����p;��5����W�}�����Ou�B��ř��
~g�����2 �w2���"�����Խ���Z��;w[�"���oҏ��/@��p��g�v�Wu�T	�y U���[���$�X�
és�z~�2[x�0zh�	���1>xcԱ>�Q�qފ��$S����#S���4Fyh�_�geb˯�����we���
�u����"e�lh�+Wj��h�f�q��\��&��yϳi�t�q%9�9�aJ�7�˦����ܘVU��֮��E(��{��#o:�Y{S�Z��bW?L����{������?4��Y������g����yO����rǂ�[0��bM��0zY����B��x��rS���9�"����-jZ��y���|En�I�E�2�|�z���� �_����PA��u�|�G��,�qxV�zn2�7#-��ڒ�M��.��y���2kN{F����NM�g�t]�;�nb7OV]�w��gPxy<��o���	�O=������S�{�F������#}g�_�Y����뫷4�={r��#=�Xy�D,��G��C�^����2�E*�E�j���F��ؑ=T|�x᳠�:Y\��5�Z��ꥄB�n�N�K���l��P���X�-g)��;�<��ޚ���u{��0���^c��&LQ��U��w����N�������cU�ZE�������x��G�������5އ�w���a~0����{t�{��.z}/l�O����t�����c�}�^gi\u�s��\{2��R:k�u,�O�����H�q�k� ~q���o��P�۟:_Gr�sV�O[X>[OO�]�~����S;�R����O<�~]W�]`�F�+�x�=�Ɣ��yhmD�ƛ{�^�z�1��9A
wì�ޣ4���aW���JNU�
����q.[��*[��-���C0M���w%�{1���@���/ay�ԒtU,�JН+V/�1W7�C�_[0���%[]ߔ�!�]�\�����;�掍�y,���;VgF�҃����^��9����HT-��>��g�q9��Я5lg��/~���v���A��X^�3����/��oiaYl��UEO�U���uv�h��:�"mgOs$�8�l�O���Q�j�E@.��F��^��(��{#8��m)4�H�+��s4s�9Y���^��Z'Kl���F!��Q����glίm���N@7BsD�T��sḡ�G��K/s�@B퀶@��R��g< ڍ�C�U�86����ᥑ,�w�:i\�eb>p*n���/��O�xܞ� 11��a��������������_��+�b��.9�f'^G���Ώk�����3y�+�#��U�U�<:����0]"�u����(L&w̃��fE"u'N��y�������k}��%��e����ah�s���V~��������f˖ٲK���B�?����^L���wȵ˳۩��o�.DK�:�H}��ِ�Jz	ॎ"`͕��0ݫt3=�]�s�G�0_��;$����3������=���#�wr��l{�)ޣ1���u���wnXW���7/�t�5N����o��+�O��_�W�Qf*M��dG���є�&�OwǷ/S��Z�N�����Q�/������Ld\���'v��S�G,|�Y�PV�]�ܩ��&�1R��-R�;�L���D>�~���`��AGz��>�8z�U�^CT�)gY�'ocS�q��ɑ��]]�uF����f\�s�D��LY�Y5�v��=��ETcM�P��=�Z��8}�D}���f��#.b[ջxc�ޟ<܁b�M������n�+�R�~���٨'��2
\��x8H��Ң������˙9�Z� ����^��W���-z���J�=�=[�69څ;/;��x8c�x����v���Ũ���WLf�op{���C��B�l0{|�{FQ�)k��W�=��	@�q����b���ᠠ۠N��d�WY1�gl`��f\u0�E��/4�vT�:�8&�,��G`��'p=ψ��nfg]�^��t%K��c��~�T�7�u���gn��Ϟz'�q��UlT���R��đ�0]�H�Q�0Rm���|�W���%�Ԗ�fz��G�vC�78�K�٩��`��k�F�qު,dx&9&gw�q=�j6�Aηz��kطPR�L��]���}<��8� 3���Wp#�8�o�¯��\sgѕ�!��O�;huyyS�;��L]@,SG���>��o��}r�RH�d��)u�@X[�\�ҫ��1�i�ݢr�* �F)U�ru�hu�J��TY�S3����/����+���`��*^�#;�y��ΫM��V���3k�D(o��
^�
���kln�k��N&1`�/Q��ԕ=|�(�ۼж���"����t�rW7�t����LW���<=!�˸9.=V]j�Ǎ�b�daVr�R9���)
J��}Yn��uf�C��ɺK9�\��ƸP"�vlz8��o�c[2���Y���l��|({/��KV2���ͳ1�=C��f���������ªϥ�l���T�t�j�r�O��Е����W(�l�X�8CfE���cc/��)'�{�h�E �A�s�����t�4�L�l�ȒƓ*�9B�}�^pU���^�
��}���ww�o�,(n�\;y���߱�ֳ��@��q:��L�ܗؗ}V��=�q?�66�1���ѝ��%mu��}��^c��m�B��'wFk�!�����ݝ7�PH�=��,ݘ(�]g\Ə{ӷ.}N�Ӄ�D��j�t�<8��Js�K8�C7%��V�S�x.�u�,ȋ� [�Is�������v	������1w�i:`\u�i[��֥>�.�.�����ͨ鉧uV)��������[��7(}�q�;�q��^��u�1�����r��=;^"k������[���zҔ�Y�����j��oB�˖�I���],l�������	�l�:�>Wd_}�gzl�i=�`��Q����٬t�v�����Y[ٚФ�{ۓ �X����3��<��)B������ؕ�\x1����mʛL��+!ssq�Eաt_W�S������n.�,*���5�̩������O�ۿ_�H�~�H�k�M5�4{��@]�f~��*o��pj�=Ȼ�'j��@U�fr��M�.���=���u
%�K�uV1nLL0�z��]9򕦟=F��XT����|;x��;"~�J*]\���7tzd�0�@��H�O�3����g��,�9⦹��'���ҷLu�w�+�]Y���Y�~~󀟫�ّ�P����n]v�|���f�
$����Wn&rN�^��N��W9u�w���#%U���z�ɖ����@�;�]���P��ۘ&��Ks�;��#����������	HK*����qb������{P�%�m�z^��׋����X<ܓ"5�!��Ub���Qw�d�1`:��*6`��B�T�,i��'tw�I���Muˋ��2�f��5�"�O"c3a�*ڜG%��s�f��5���6���t7fo�J�`��Q���̔�%-�u��Z}��s����U�x>�A��'�޵Con��(b�VR��ݜ",-�vؚ�:��t�����>�L:�]_�G=}�М�Þ) �I_�Glɒ�)-�����!$�|�(��1)M�b��Xk�����tI�w.lC��{���G�:�.޹�����M�흔Of�f�.�'�z��c\ү�Ès���=O�e�2������yS�\�`�x�?��Φ�)��Fk�&-ݵ菱'�;ު��NK�8�xX=X�P����qe�D���W���Ϧ���9���O�?܇ȳv|�����g'�jjE�t����}2k3�&`/:��o0w��9~�'�X�[���⟞{�{ok4�C��:�T��f�y\L��z�m�E\��oo���6�O�m|�)��ۡ^�Ȭ�QG��Op�:�E��Y�{ӑ���mOx{,^��??�yyhl��j��Ҧa�8@{Ur�����lɭxZ7��܆�TZY֧��L�B�݃�7F�ڃ��� ��������Wϼ����E�Jy!Nc�Z�ā��ʄ�e�	���-�BuC�*�T�90�8ߋ7��*:u��N��QՓ�W#SBw�!����Wꞿ\��-Hp�,�}Bo�����컊Fv啕g|�K�c���y�߰Z�eq*��iȿF�ʪ_�ߗ�~���g��-�T�s�����ùR�S&�F�Χ�')'I�7�����jvCO�p�{	��VSY;��5�Wp]����磖����[�%]��ug�Y��y��[��������C>.I �,1/Q{D>m�5r.��o^��ʵ*ߝ]	)u5Y��^���I��ruc��
�}p,��`�ҷG��i��f�U��-��"��֯qP`f0S3�5t�q�5T��}]�Z����ɝ	,�D�\Ȱ��kP9R7X��󚉮�̘��\�Ԫ�����Z�]�m=��rQr�U���Np��Z70�*��w��:a��F���9c�f
G�"*{�+Ͱ�Yɩa��}�n!����;�b&-xŜ�М�T�������h8E�'Z�Z��K��~��c��\Oy֭��VbPT�7��Sv�El����Vb��u��]�]5�Ҹ�����(��{�I����"����Ԡ��;'\�R�:rs̺���o8��x���jg�5˖�9�,�f�������̼	�������d���j��{�:�m]:���n�A�\����:ە��������s�a���s�N�⫎���oj�ʅQ/�$v:�U�waFś�EY��TMn��H�%�;��:��p¿a���\���JQUwi��}�+R���-e�LK�OT3\ז��Z���]��sN�'ٹ�����ڿ�B�wb�C���*Z �3X�n��]�ţC� �iֲ�1�1)аV,����ÌzF��9���U�8�w�s�W������%��:�=��K�b�NUۮ��D���
���5�X�;�uط��1vP�s�	�~�~���G�&�S�b�P+xֶ�*'W�gc�dȶv�-ƒ��I���'KO=��N��mC\��F먾�GG:��L�א���ˎ��SF)��3D!����]��MΜ1�j<lu�S�n�h�Oi(�tλm�Md��_h��.�=g��6
�F�]5hr���-���(�E��f�jM���t�q�^�nu+A:ݾ3k*���\�Io&��k�jQ�wn�6{+�����	�4�BKN�Ԯ�]VHu��*�#,]UtpiNi�o��W#f�*�Nk�TȨ�I=�A%�h�1�@1.)M��n�;J��}���-�E�سo���i-Q'As��PYF�`�Rb��;@���1Cx]D7s_kݡE��ܠ�#����JjD�u��x�Z8 �gV<Tʫb�g�J:�\�t�p𕊖�r���Lq�j}Y]0��y_$���ւuU�� ��V�ٺ�[λ�5q$�.]k���y�JRA��m�Z;&�d
��"���B����/0��`;�U�{�x=���Ȧ���޿�<��uD���\ŢZ�2T��׽�QK�[!�{tjP-b���.�L]Fn)��M�BW3OSPn���l�t,�`��M��tT�c��Y���ڀ���J#J�{� 7)�j�}*򳙳J���� �l/��u(��}���Vk?>x��&� 
� �}�J4�����Dy���yt.�)9�pu�"����tS��S����s��T)��޴5a�λГ��j�b�������D
��i�t�.}DRIT�Z-��s:�V�۫wt�&��^���WCW��k�sGח�ui\]�3��|N
�Q��o[��^��O���BW�w������h~>�������$m���p�#�|�ʘ<bҖG8��1\U��h��o'�|�W�7��	�¤��z��=:�u����l��_�C�p6(
��j,�k9�hk#��#:.�������޿u,��Pˊ6H'Y���;sO)<�C�B��mT���[�p�l s�e˔�x��o��{�}ɉ�����P�ާ'+z����p�wd�]���Õ��� -��x>���^���d�����s²g�S�i�4�Fg�W��z�{��z��у�y�H�j�fm
<�"
ێ����WV��_�<�M=�`��k�E�>)E{�Ӝ8���kWýy�o���Q���7���yX4N;��	S��X���z.��}���1����ݾ�ه�:=з�\�*����5-��YtK��Dx+S��:D�� �6�{���=q1G9����o6w�(�o+��Cm]��ڏL���v��S��o"��0D�}�S��U�]A�ЁT��qP�)�YyD�P�̘6��Y�Z}�S���p::T,���s]���GwL�p�\j�X�QΕ�$�2B`��G�}w]r�	\�VTtn��u}d�T���l6�d�f�J�^F��:�mY%I����G���q��I�1]A���h[�cG��dLLg��-=әU-ݟX��>�}F�� {�β`{)Ҏ�����r}1���햇������aHz��gj�GUA���鋸!yg���7���rZ^���ZN^e�ZB[��v^'�{Ӌ��.��|�:���s���߬�A^$�z�
߄o����k��������fD�c�sY�P���[a�>�\��O�ӓ�(�ěX6����f��T�����7B5�t^D�5U��>\���HV�ޞ��L���)��eދ#k�V'M�����>�����a�.}GZӓT�m�|щ�ѩ�穎ͅ5�4�����2\���4�h���ˬ7�S����^��٦������&�l¼S��4"��Oh�v
�����q]j���GԆΛ� >Ɍ��ޥ,*�lѰ #��2���/p
S�c1�h6��o6�L&	�H��`͏&��s������yj�2?������.�lܱ)���3�ʙ����tz'�g���Y�E���#>�W��W�;b�ۅY�����R�a��l}�!�� �b��TA��'��O�
Y��zc��¢g���������1E{��QZ#�\�_�J1���ބqYǵ�ۂUk����]G'n�������JΜt��C>�&�\	2�){|��H̬��83�ە&߫�~��q��TX���|�tX��G����U<�I��9���F��Vhw���rv������Z<L�|x��_l�����6�|�_�n���h��>��^t���}�=TaO f�YW�b��f��ga���=����߈��]E�]��;�-��5����[��h�ˎ8��am�j}�"���=o���f���q�>�w�c��*k>�Տ��?�F���,���"w����p��q'=��C��M��VX��7�j|7�W�}�axv=A��߁w1o�(�}�;&;j`�e�v�o�NVkZE]4�F��^��C��Fn��j���ǫ*��V�]o�'E����娪�1%r�^я|}���1V6�[�j��X�N��:51�^cbL�|ᅲ�޸��^��]���?�����s�����eY�o�N޲˞ưH�>/;͔�>�ص}��'EK	;�M�UAG��B�:D�����~	q~ل=8`�>�*ݛ��ȅ&ǇU?�(5C��G��L��NDQ��/�׸%>��f}> �W�63M���p����)�����ns9sC�ԣC�r"��Ok��n�
�lD�ק}���H��E4�R���Z��˔��^�cynů7�ض�j�bY�'mc���\ ��������
���/U=��\S��s�|�{-�[�g�7ٰn�E�Ha�~%K�t:��'�d`�=��z1�F�4����� ��=��Q��9
��t+t	�Ǐ?5.�����s܄�u|(OR����2��}Ez��]�\�I��O��Eo����n8�Ȏ��e�l�r�(��[@���k��t4Ԁ��=�b� ��2��J��r��n(�8i�0E�z���r�̏`>z.�Np1��5���Mg�{j��k�l���-A�=�����0I1����-��o����}R��]�W�:m���s���t~�~�Q,���� 	M?]�v�n8�s�K�7�-G��qvt��0m_�W���kPM��R}�v�
s���Y�"r�r���ܭx�׊�DY�w`Os�h_n*��"�t�x�uݏ���C'���������s�MI�<Ƭ��,ق��/'�!p׷v��O�i]��U�ÎJX�p�z��.�1��p�,��>K]��.��_�wTz;_�����sT3ac"EX=U�R�&����i�
�@��y+��?��$L}}F���f������1/O��H�-Ѹy�Ty\T�)�*sU7���֦���gb�{�k��F����P$)@�d���h�$����%���9WF�َ�&�Wn�xp��#��G���g���\YB�~c��Ǥ^�A��2bY�0�i-L�.KD��]�ZP��"I�z�[٪���F��b�.�Z[�N�̵Vx�s��u�lفr��~�����@�pԽ��w���;5�~/��nY���'Y캾����?	~�
��Tk�A��Xr7}�ȶ��{� ���sU����p��G��=�-�^J����k`[��֙�QS���6az��}X��Y�r�ܮ�?��S�RN]zn(�?���w�_4�=��a9�v�#J�>�U]�csBE�4##�V]�M��:��{��Rz1F�e$�E��8(�ѧr$_�N򜡕s���f&;T�3-KiLɍ��'gm��$�D��N�/�����ٙs�_F	��azN����)'�7=a��2�^�h�uc��XS��[�3�W_'�r51���GҍdU�h��8vHCLz��q�Ui/b��;U���O"LW���J�4j�ϴׅ(����A�����u-tZ����J};Rr���g-f{�h�Y���e���;��.��6\��B�Q�w�(z�A�f�LLF��ko�|������uCW�
�7FL<ɭ~fׅ����뉠�&eoRܑ~�1�~�L��dlOz�8��S5Al{��U���$h�]�aR7������Jǹ����۝�_V����ȳ���l�fl"76�WY��/@0Q�5�Sf���t�<�����F����!��ʻGk���<��&4������ՠ�'�7�o-����'P����)�^Ş�[��z��~y��UH��.F�(�.����[R��S���iK�ev�^Vn�[���1��N�t"���#���/�zX���`m(:_�_���QbQM��	"^ߦ��vZ=�4;�O�3]�mF�e���=c!��w�h�S���~��������ھ�����j:ǽ������[.A��8:�r��T2�,1ө�:�wimZP hL Y7|��\�y�omOAu���蜏VT�<>MFeyM[�Z��|�õům껄6f��D��[G�.ǡ������􊹂�[*�֎!�D��	%
�16�p��Dn��<���^����j�G���\TH�};O�ǥl��_��~��v�u��[�|vm�"o(D�wx��kE��F�5�Y}�x������V��î��_z�B]k��[��(�=��*쬥η�^w���EN�eFTa�>K<��J�Oo�O/�;
8՛�(�*�����*�"�2���C��vO_]tW�ɇb}�<�D��˂���6�N�
�� �G<Y�8M�wA6�*j�u8���OrS5n��v^Kq\v���ݳ�Xԅ�����{��N�,���g{[���&��wm�8�zy�Imv6o^0l�]P���v�@:��Nٜ�0�a|��&0g[�9%�m��H�3�]mދW���#,��{½�۴��O=��g��(�+GE#�t�wM8�boٵ����x-߻��?|����v��r�Zٜ_Gk�����ߧWOD�<|��1�����j�ˑ�Ϡ�_���z�Ve�}���ys��r�i���$Ys�:��;up-�</�*${N�Իj뷊����s���'����<g|���Gt��P�����_��յǵ$����<�6����?�� �_��
��eR���NOT>b�U�v�x��g�xqM�E���Ӿ�Z���f���tdM-h�^!ywS���'���.��\�MEʴϝw��_ %�,��>֟A��l��|�>�x5b�]�2I��j�5
� c0*�q���Vu{��B{i�O.�GV��lq�Y<�1�{�1�9��I���ڍ�L,�j���Sɞ�W6�+��E��k+��t�{��׺��,�����,��{�n�V̼��fc{7!��rwN�E�}P��]�=�����Yl��훦�X��o;!h�uԭ���d��$��N}��(��8LOo<c��ӵu�C�|�����Xτ�*Q��]���d��e�#�z�.�m3��i&����6H� r�'5��,�ն�5�"��	q͢��[��;���K�;e�t��9)Y�A��������U��ݛ͞�����֮��=�n�}���W�Y>�[t�8�?��1�}	����?��u?��^��8w��>���S溇��1�yJ�d��õ)��5׾.s�w����E@�Sj�o���Ѝ�I�f|����틼�8BWNx��LW���P��T�d'��e�J�=@���^��6w���>$MzI<K�]7 ��'yf<(�G�p{�[e��k�ICf��#vc���=�+/f����EdΗ��g{�Sz���k��H�pW�r�y�uB���'p�}�*v2�$S��{r]��U-�]]rF[����Q���]�����[��TS�f$��m��v�����ġ1���yM�q���+����k{�Z���6;��Q-�gp�b������տ8^��Ds�x�mm�lC�'o��\qvO�i>z����-�#!kF���F�>�#�VH�#���5�ub������F��ю��Ajկ�P!�ZF���#s0��w�Lq����T�m�}�����C��=��棷yF�ʮ�/�@��=�~"��i�XP��`�ն=�;�3д|)������6:��Ǻ�Ӊ1y�ﾈ�^�/��0�'�$ �Z����)]�����&�;��{*�I�6F��T#��q7r�~'v�m���m~�f�+64��q��ݧ�ms�q�iͮii�iP�K�����m�n$aj�.�"A�6���Ɓ�u2r\&��<Z�uD��Ž�Ն�1�o*bc,?������|�"!^ڈD���j�OhE��6].w�������#�&������4�������[ �,	�ֺ�p�����O��^���yH�7����b6�l��:�=��5�m���O�������%�?!_3��uҺ{\|~��{w=>#���u`h�9�:u<��н� �d��2�L"#'k�]��5U2/��Bq�w����Ɛ��b�O��d���k��{�KpV���S�gy��ŏ.��;Ry�ڹC(�m�s{�jy����J��/^�s���b�_�����09�T.<�կz6~��4R~U+X�}�I�5�,�rg�bN�l����)⻡쭡F�'<.�;�k�b��'U���7v�^]��`�����z���t��s1�>��4����U�_P���28F��f#'�����0w�����ns�{�k�g�C�Ӳ��r?�w[C���?/�SF�}^ycw5���M��nu�@�K�m{���/���W]w���K��n�,(�TF�s�4Ad{�b�J�A�J�B�Ut���R[E5SǕ�&Ek8~��]hÄ�3:�U�ɢ%q�t�֖f���(ZW��sR��y�ٛut��<��nU��T���Z<1^��]��u���st�)�Z�WB�k{5�t�r<�fL�7� b�)���nL�S��J�xm��
�B�1�Mֺ>��c�"9�7��4%jj�9/�ѱy#�{T
"�<�`[mOR�P"}�5	6ʽsj�|�rhOC&=��y�{�8	��O�S�9�J�34���ˮ��W��w�f`��T����p%A�S�����2��P�w�R[/k�!׈7x�2P���V�Z����ZD��GiR)_)�c�y/|����}�-m�P�����L�3�v�{���d�p�����E�K�������o~��5�~�pJ5Y�#=4h��l��>{�oHE�9cpV�һ�~c�R��B��q�˓�ꮱ�NJC�^�؄��~ܕ���T��wcJ���]w�n������d�t$������0�sXҡP"�uӘ^ڑ���g1�~�����@Հ��}��y,���r����sW�|������V�t}gF5q+�{ER�o�pO�G�'��y�.��N�Fn�Z�:ɣX`Ğv/z�?{%��`���v6o輊f8�k&F\R���\^v#�n(�˅��T�!���r&[U�B��C�QǑ�A�.7ϖD��������@!J��5��.�"�n�� X)�a�x�{��6�`�H��+���<T�M��N��lZ��`3lT�����Wm�{7�L�6�ޮ�Z�V���g��)&��]�ű���
�
є&n���o-���
iZu�#�]�b�7��֩͇]J����۵Z2�N#&����NW�'s���[I���;��������&�7�8cX&q�jJ��7O~��5��.8`�s�B�ړ�>je�S�oN�$�s�̱c�֬
��|�J��On�S���Y�%��b��É�Ej�kq������pWa爣�ݾ�j��o3"�~���ڹ+s��O^;K_+�_�=�!����^���!Z��r�.Q�ҋ=�t`	F[΢��v��k�����_;�]�kU�;M*��.�|4��kX�|v�HA�䫕��J[��0LӺ�w%�f-έV�4wvj�����)��H��=9U�wo�V���QwN��)�:�u��^6q�[�H�z�g���O&˗���*���ڷƅp+UH��+cm���J����4��3j�u��غ.��)�F�uY%+�j��0AB`@]_V�"�v��hUq��\I�`ͪ����6%�����)ُ,��v"e�w���u+v�3�����d��v�6��WP�R�G	�.%)�y���J�U���Zdu6�:C�wef���r	]�e�Ln����������Z�����W�K�p��5-nr�t��B��}:Io�}#9 q���a�;E);�m%\���ۈv3�&�Ys0�`}�mAB��H)�n��}�rդܺ4��/7tZ�%Xa��d����ci^������w��<W��$է�J=rӏnrKx<��r��p�GJ�ˊر��Ni�;����.�<��t���k^���[�o=��2�Խ��OQ��q����;�O.�*�^�5�Q|x0�[��]+��Ù+v�na��~Z���ι�D������xʘ���e�v��S�;�VX�s�S�}�}���=��O�~�x���W}$ŚDWg�.�ڱ��=�~�w���Z���80sx���͹��P<��AN�%]*�F�0�>TjTD�Ҩ������X��W��#����>e�4��j�Ʊ[�շ�&!|1���i:}9 �Ɲ
p��}�1�b�'��7�ZQ�����P�ʃ�ۨ 7n�&k���6�pËA�2�A�{[J���Y�f�\1uٰ֛lrw]X�Rۜ���!����1+��f�9��)�n��,��9��n!'K�Z�ݢ-�d#.G��f�P�t񪂙W��kF��P/��s�^��X�k.g:�5�R��N��!������)�:R�6�z6+D���fc�S�W)��nsyM ���ԝ��[..����#��IP�*�2�R��ʡ��5��n�Ka�	w�qt�(�o�̰�9ɱ��5�5����S'i���w�o��$sy�]pT����ؔ�S�u�kIݺ�ӷ{9�-0��Z�ż�Eq���T�IYy9(	.Z&`�r��������h��L�|�#�e�]^���7Y�xtx��b���y>��ծ�4C@�ed��fl�� >��.l�l�L8|��
���b�#3�u�|Ip	!|�/A���-@�{�{}���rAmh�#�j��o�Og����o�޸6q�FCYo�ݙQ�z�n"pQ�w1�8���:�r�t��苧��W�t(�\~�4�W7����x���Z�D'����m_R�|��7�77w�TK��+�E�*t�^(}~���2��M-Fz�s/������zt��GS�Ϫ�%(tb�����d������n�b��d�b�.AU�XGLЊ|�Kj���+}~�D��&{�t�X;�$��wVz~T���k:��Te����y�=7N�:~d{�N�_�J��y�ڽ|[P�������c��c����zή�TP��Q�z�޷y�`�l���}ꜭ����+s���u%�#6�q1��>�d�Z����\�7/�mW�W�4\&k���e�L�?cJ�ߥ��OP���O��*���P;�ц�3�&�7��+��Z�{b���<ڹ���$��O1=E`Z��V��Vh�亵q����-f�T��{y1����S(�cAlޣ)������t-J���,i���{��ʄ<��#��n2����[̑�k��B]����qt)��h�����1���8Q��t�3��H|O_u�yh�8*����ܟ�ʻ�kǇTҭ�'�:�� �2�lr�]=o|��+>n���[;���#m-���f�t*v�����o8�lI�xv��6gju���|7��W�7:z�I^�_��I^���{f��jG� �����ޢ��2�Y��cgv���݆Z���O�����ٌ�B�Ng_��]Ւ+����ZpE	S�M�ì�*eZŶ�EY^,w�RPY������M2%�j�Q���39LIa���F0���ٿ+��u]sf�{W��U�.�o�x�����VT���OX\Y��S/OFԑ�z�5ĤT��ƈ����@V�%���o�s6����o��?V���w�r\���et˛1�Doi�&ĩ��.LЈ2�z���̞�=z3ˣ�Q1VΑ+�&���S؏(�!Ej���E��"C���>�K�Ͻ�ھ���N���k���>��uH�ٙ2E֑+�@y_,�^T�"�
��yv�h	�c������"렛�v`�`�KD�Q�xi	����髱�_S�VY�Y��5VwiRSukѕh�����N�zVAY4�ܮª~��Xx��u�/���r��\p�\�ܠ���b��h�����TgF).���;݉q�
p�w6p�7�{�<,8+�AK���f�R�]yJ��}��	�IR�%ԯfI�CÑ�j7WI���;�q.�����-{�w��cq�#��n{z����j�1>�!Ot���<]څ$z�����yOP��`�^��g�+��9�PB2��e^�z�·2���ا�~3�U0�5a�Y���R�>/��}�G]ܯ���Q�o�Z�[+2���[�p]�;Wګ�]I��>Dx��P�$6����ul��g�_b����L��7��ڹ^��5;�_�tק�5잔��_��Zݮ�m�j��.R��JT��w�SԳ*��==�W�P^�j$t��rCb��B�+�����_��쾝B�^W̚y��9'X���\�ڕw����h9�Пw���5�^33�Z��:	�&㏧X�yo�^j�1�:�����������ÐA���u�|g8+T���Q��&�{4��¸݇u�=ap,�FOgn��[Ew�)w�B�rM)����͑��
K���J�W�\K�^0,O��p޸��\u�ٻ�]~�nw²�%��L�,j�ud��BW2�Ɍ��py�Nu�,� �*�ys�w��@�$��B���:��ŗ �>v55VvB�^1�_!89u�U���,G��¼�ʾ���?�mTU��fg.e^"��55���n����m�������J��PG%w;ʙ{2�N:�\썠]�X�k&-.�Z�n����*���/��q�*2)f��96�=�M�ak%V���wȽ�5<��;Z���>\G����~�~2���v4Dɷ*(C��L��o8ß>�~�.l���[=к��l��S��(���;RE��h����k�gt��9Rei�肕��r�)�{���Y�7r"��s~���E�����P��Ld�2�������Y�n�̈��*��ۭ��4g8r�7:޾�Yg�
���Y��H�V��Z���ٹ|/W�3�;G/���wP#T�߈4���3��[_�yy|J���:C��N
�����)e�#�I�fY�t}�k���1|@���H�/^�_����T� ߥv�9�)Vo��l4��8���8ZJ_j(a�yV ��2J�}����gz��Nr��f7t�r�Z)Ni�ރ׭�6��|���ϫ�e��(�H��1�kVMD�[E!Ϝ�nr����!l;b�����\LS������Â�l�{Yf.O���ز.��(u����5.�A�J��q��3��ZtV^�8��)w�S�dA���F^��&�申�ް�:�z��Jw�lX�>��~ā�U��a�|x�nm_JB���R����ͫ���[Gu�S]
��p�m�D&����]G�1;$X?�E�Ǻ�^h9��eC2w��܊���#0�3c��<�m���;i^�v:T�ޖ�6kB����Z`�L�&n���N��]�Қ�X=�٫�GV|�Ƨ��3�=��������ԝ�.���T2�Տ*�66�π��Z���3��ƕ_o_\�^�����W܄�67r�Ʈ���s����U�
�$��GO?xf݆�ʁ��<$:�37[��T���Y��v�mC��,�v���#W�WYv���{�٠ea�%�϶��Lt�z�vا�DU��$!{��T��i���"�vH��G�к#5t�P��]QG�L��>W棴�|FT�g�f�����g��rQ���u
_I��|�\�ǩ����EES����������W��r�\@B��Y���㖵���҇�(�z=S4�؄� 9QM6,�H��K ��p��zW����B���>���+:o9o��7�J�'��_�׺��3�u2G����%�M"�NY�\q�n�V�Mh>»�GV%�v�}C�O�.<5��j$l�k�k<[�[mPv���:�z-��vPW/~�k:�����~�%��3(��6�ɺ��#��uuF��iňK��呚�1�s��= ��j+#!��ȁ);;�D�u�Ӎ�$��d����ݤ9���]�:�n%V��k�&\1��ૠ��&����?��i�(Q�����;j�!�\OM��^�l��g�q\[�E��*�[�Mȝ��@�D ]<����Ut^�̎�ztƦ�lu��Z&��%�V��uNI�~����P��!��z5�>�^9���U��(��h�]8��>'�}�l�TC��NV^OϠhj4�=s�븭n5���"ύK���Sڲ.=��j=Wt�������ڞW�j�5�V>��{Yo��x��V3u���tʹ��k����L１[l�~̩���jU�
s�Xq��{�m��O�V�+���|'N�#\��^c��&&��a��/��k�������S�Z�aį]TZ��	����_�j�.� �����6v"2���^T��Rr�M�-S�}�T@����dĶ��r�����b�?��$�z��r��c*Y�����ޱ5��/�i<�Ng#T�+c�~�w����㾛�L9+.�&��p3ނbj����&��=G����}M��h����y�3����>dL*��[�o�����xh\2��x�ϯ���һav0oY�fl��L�f?v�a����F����ԳϤ�ٔo����1|=M�<W�m������l���x;`s��l�ٱ�Q���hn!T}n�ܨ�7|i�V�˨�#;��CfmcX�Wd���_q�L�MFӸ�XAcγc"���킷{1
ν�d�8Ps9ܶ�e#}�i�+ܾ��f�M�J���VQ��l�B�'�So�jեm��ѧy��E&��'+�qr�S/v�'�z���m>3�9��~?L��սDD�+G{Έ�R♉�6j
>��w����H���N�>љ>�������zE���3z�n�~��}?]]�)Y���և��j���٢���c�(��k@M-<������Tq����jG4Ӭ�p|�z����hx����yl6"x�A����`�����g�v_J�{��~\j"b�ָ�g��lP���&di���`&w�s�,�R�6�)�v?G�Xep�կ�#O�o�Xɣ�jP�{���Yܸ������7��5����=^]]�S����L�K"K��=��Ǆ�]r���j�=�ϓK���M,l�z�c�.�@�Tϴ =C.Q��+M�N���g�{Y��cʱâh����d�'�r�i����(I�ڍ�T�Ӌ�1`��^9å��q�N֪|M�{ԡyR�")����<���u]t߬��4��tl��
�c���¾&{ʯZT$ı���˅��/�M���s��Pz}���o�T{��)���)œ��|�>��sD.����>�<]s�[�g0X��הvf*S홡�e��
V�S�9�ޗ�\7HP+��f�� ��j2Z��Sc�h���K���@n1y��՗7;5�J���2	�	bs�o3tg}:�f���Yt�l��WO�m���V��Ձ�>�h0�>���m�C�՞r�nsyA@M��O�p]�r���:��U��;j�i�Ur�*E�w��ۊr�����+�s9�K���\�ݨ��,.{$�<' ��jq]��oX{�C޳r�e��#�ѩf���ȹqU
�n��5���}�Յ���/��q�k��q�#�|s,,�Q=�ٗ[a.�.��)�me*X�� .C���_�t�׶ t\���sd�W}����ǯ��%k����-��F	1l����;'T�95��c�F�q��/�9���}Bŵ�WB��ׁص�o�Umԉ����MNZ�y�!������Ej$�g��Q�t__s����W��[1������W��W�d!�j8��-���~�Q��Y~`��*k�ƪ�J6e�랼�HeѮ�;��5�z�������r��(�t�rM\�F������Z�r:�׏¹��=1/O[�7D�w�ْt���T�ͱ�����V��D�R}�`������Fp��]v�����:�ß_a�S2>��6A^�ެ
����g�_C�����So�%=�H=���"̦�M����=���mq�^��;0��f��>�E1�\<^u~�T����l�!�F��r�_�;6�F6�4�_$tb���WY�ҍ�mDİ�,�mTv�IK���y�Ԋt�c�7�I��5�a���L�c�9 .��_p��K�B�8㳘���#OU�����q�c�ad�	a먏�k�^�rrnh;ݳ�~����(�C}yn���:(Ѯf��Y�o�!�#�[ޛ��(J����>��}�rZ���v�ϵ�2�ķ��5�xwo��2�p����J��k�>؃��CV�6ɮ���c"�<A�O�_L��h^�!�������ő�o�W�qި7wo���˹�7�K�ڂ���{?����Y�v.�<���o~�#͎򱁘��[k�p�
���&A5J�D��u|�rH��^Jj�mx�ɖt�r=[jD;Q���ޑ�Rj湟H4+�:�{ Þ7	�tϞ;�f�Ȟ�7�j3�0���-�ڹ@��cΏ�7v�{���(�����c�9O:��1FS�׻�ȋ_w����C��?W�dk���:�$(=\��H��[z���%��C���V׬HF��=�R�ۼV����Nc]b���KZ
�̥���[��m��S�y�r���,����l�v�w�l�Up���}��~G~���^.�;/���Egm���Ϗn�!-ާ�zP!$���[�g���ŏz�v�v�M�ѳ�=>���Y����NK��r V��v�L����Ҙ�����x��Rl���p83��8��۾
���P#  ���������0Ut�Տ�f��GQJ}��m���ӭ).ֲ�.�)��'lK��6��ƭ]:��O7j:=�s b��Z�d��	�6�`��;�]�ݑZ�l�<��J,��u.�`Ȃ��8��|�NP?�R5��T�����~8�e���{F+���=��`'I��ˬ������r"4��<TN�0b��
�Aٮ]u�am4&s��x���+��.����>rm�;�#n����H�|wr�d��7�uGE�<^�@l��3����N1:��pi����Ț��,��uw��=�-����a�Uhdb<"�'����rz<_����Z��2�`ۮ���s�Q�"{0ϣ�ɘJ'.�m0��z��|j\�����1%E�E��;sv�!��h]>r3yd�J�U�����Q�bw c��)�+��}<#f1d���)5|��x�mOJ�9�o���$��n�]�ϟ���ӝ���G�Һ��}{�s]Y�Y�^ �T��@o�'�_��E��'��q[=�zj�VϞ��,�����)-��4FU��1B�i�a[�9a��^3���Z��qU؉����%=>=��,�a�k��4��p��|<�g.;ڲ�c�i!��=m��oM������RT>�"�o���h%�s�2;OY0����3לEET�v#�N����Z��AYw��Mp [��==�uniU����:��+@����uIYWu:ty�֮ce[k1�T�&l���W�
���4��p��l�k�=/��+U������ur�����:����,Uyf�d�Wݕ�u9cA]v�k��[�4���t�ǡ��od↾��\���t,��v%��j:�[�%��DƂ�@E9�G���ZΝD�;��o�w.Q\�L�%>4�}��2�=uw�up�V2v�9)�j\;���X�5Cv��Q[@��a����\��d�����=KA��/vƧm��-�P˾����ô�9�5db����v�]`����]�9:��-��U�`���޼3j�n:��Gx�FCխ�̎�-3��qap7&�	k��?����G���-��%�����V�+#�v(�tP�+9�JK���%��ff]�V��wn�n�eXc����#L�R��:WQ��2l.f�4Vm�`e�D�+{z(�b���mGn�������rx���{��:��ZZ�Wu-ji�w+Y�ش�sy�&̔@�\��5�tOvf퍭�.�sf~i'E>Q����oA���1Afb���e�?�G�{�:,�X�w�<r��ƜZ+���<��A��7%r��bi|����Yy�G4�-\�n��f��w�.w�����⌾C�)��o5L�U����]�>�N�Fۘ��gk�ݩ��D�M�:��O%|MÂ<���u�g
�S���	)nV#�9����9v1~x���\��\��J�Lz]��;9�؎at%��s��H�+�p��>�������ھ����B*���#��ѓm�jvr��15�����P�]fumީG��׮�cV���=]/!�K	�rrG%�o�(7� ���X�a�̾wѦ���DQf�Cv�����X�[/v��k��5�z홪�'K�9PF�(�)y�]�gs����/�>�ܻR[���t�ɹEK�nv�V��HI���yW���S�eU�%���gy��׷c�#-"��'+�Ǣ��81iR;[��
�5@�K9����b���{E<����T�S{t�=�������y!���.G�qPD+�a=�D��[7 �ڃ�R�;ns���gh�Î�u���A��x���5V��V�MʤTR�r�N��cK�8�o2�*˝6�c\V>�,��2�Bv�y�������*򚃛��c�й�D�5b%�w�]
�+���OgY
n��c8oQt֡5$������9b�Du��.�O�X���������gT�V�7[	tR칣 ��7��a�;V�������R����N��Պtn嬩A��!�=|�r��
U����	���W�/�[�������n��w�h^��B�\� �%֋��ڻ���;8]�jr����mU).P~#g�3��=T��d-o7׽;`U��V/tj˹Gv��Q���wI���Ud�񫒐e�Ψ8�ܴGb����o��lA�^�&���Q�8�
]�GE��<=ڭ���4��a|����V�p���z�9��ٯX��I�?F0�s�{��R����p=y�7ypu7k��d� �Q�k-E¿5r']�Ŵ(��,�����2f^>�7�ϊ��3O
�����̎��̷K��#�Los��7�Uf�;Xg_��j�g]d�����</�|�n����5{׷יs3=>ϝeg������U���"����>��X����o6����Կ'�OB�t}]>���Z��_V��f��&-�����G���;��7I�,ˎ:
g�G����s�u���*�s/�	��xGp���+�v��b���C�|8W�w�4M��G=�`:��;�dMdv�2�Ңb��]՜��l���3*���39�Z�O����CIp������'R�\�EF0U;]�(-���g���E_�}��0���T��"C�3r�����\��UHu��yC�������ki-И콽���Ǵ~� �����׹,Aʙx\=�h�ܟ\ъ���R��hj�o�S� �9}���@�,]M9�s��owU��of\Y�^ne��u:�g3���A8�]�}�Nv�k9��fe3�:�n->���:λʛ��\/j^�];|XE�C�s��B�-���ʩ=1*���N���8a({)�O�&!�.A�\�P[�F%/��r#] ���{�?n��Y��ߠ�)=���8/��������H-��e'GnhZ��[�O}K��h���w�u׷��E���O��v�;E�`��X�9Sv�oc�!���gۊ�`�;�7�>��~�W:�+YnΜO;��f�vʯ$Z$��'��{W���};46��蜛�-�@�y��@�l"Ϗ1�;^��6��kǚؚ������ꊚqsb���s�=�*F� ���j5��`�\]t{I�A�q`�}m��%L�R�uvb�۟X�#*E�7�ӌ3Vb�&�b�˧�2=���x��K��wE�y�����f'�Ur;�U���Ӓ�F���,���q&�<(۞hϹ��7�����^Z��վ˩��9�y$�7�,�7����2SGCv������@����𽘭�����s�����|5[��^��M�"{�aA�Z�Я�z"��we�8�-�d_�z���zy�k*Uo�(�韢}���j��:�7���0R׏ULcgN���5����J����,{.�$�K4a+Iۨ�v�7Eh#i�ȱ4\��%����u�om�+K��͆���6U���l��dwv99�kVo�k�|�|(t�+F;�uzz��a���H�U�)U�Ug��� !9�zc�}P��hù��^��O�HJ�"����+U�~�."�>�N�5��uN�V��YHo����4����������X��*�����%��+UyB�[�?z��:�.�lu~��Aw�O���iA�M�|����ꬣ�Lq�Z�Ľ����t(���3q���t�}��G�B՝��A���]�[-A=)�����g��B����T?f����[\ȃJ�}�p������B�y	��.��C'0V?X���1gX���UK��3ܓ�@@��z����"�t��Tym��3+=�����WF!�-��7��P�gq�a7������E�QS��^%a�F�ڟGkRwH�\(�mr1�	�1-J�:�TR�������#��OkS^����ȷ�\]�f�̪�9>.Q�Е�dY���ʛ�ڝ��a��?n��l�7��~2�X�v<R\���4�����δ{�-��~;��� ��_j�i����!VVHj�H��􁚡^��՘��:��ء�F���2bux���2%��F���Ѝ�L�#�*4�h]q;\��1C��a%�N]��؂�.�|��$�v�V�{#��d�gR���y��k�;��r��׳JV-g46��l6�ġ"���Ħ�1Vf��q꼡ҧ-�6�|�H�7)d'�N��y&��z�>^���~|��u��x����t���x�E@���F�I����5ur�`��n����F.��	NV��kr��~ݪ��(z��|`�U�2�}����`�T�ϟX�s�fD
mx~Vm���y]��x�{AYF�1��*�������u�Á���~����;0��yD���7L�]/DHY�q�,��_.�3�"ؽ�i��OOI���I����hApE�&�/0OXzp��2�ـy�;�.�>������*���v��oɯ'�U���;�����Յ������`a§�zҞ��i��M =..��$@�[>^�{�ځ�&�Q�G^o�5�����NƯ�Sc��e\�M��ۇ��2F�%U�n���EѦ Dg�a1U�q��&��'�Vv�s�n�;=���q�`�`����G8`Mf�3"xl��|q�@�=�EU`�h<���5N�7�~�te�m	c8_���7�炢�W*�e�#��l��Fx
��qi��7*�{�D@�r���:���o�VA��ߑ��ۢ}�3w�^w��a�=|%��95�p5E�5�����+���r.T�s�q�놢�c9 Ԙ���2�I��~�oY�*�W��b���<��H�����&ٰ1'\(~Y	%�hh�Ơ`f���!Õ�[�9W�lk|B͝��b��]�`�l�Rt���t=G	���p	�qmN�w���
i�"ז���]/e�?�u4�g>���0K!��v����a�;��mdSoV�x����d:� N��B���_��n���s#�d���s��bg�,N��������ww|as����!(��������S|�g�ϣ5|�:t^��߸��`�W�Qo��C��O	��A���^�-�.ita��ʢ*�|b�M�N�d?Y�}N}&���uqva�d��m���7�+�xs�Κ��E*���cԼ�@�&�l��_Qΰ�����|�>�`�=�
�
{��>�L���酋c�%���-wH��W���,<����U�֗y��X�+5��:��ai�m���*�=�y�X���<�O(;���>ӝ����a6�"�!��w��S>�Q�{��s�n�~x��sN����ŋ�˲�h ª��n��g�THZO�?zo
�#Æ9T���8���jׂ�����pLf��^�_h�n�.��z��5�#0����Y����Y�r���w�kfp�? l��r8=�X��0���L�/�{z�}�:l�7�r���bov�
���m��T(�z��R�T����7���o7�c�����s7q  �ڈ1����
�'z��l�wF��.�[�Sιۙ��e�sg)����~����Mu���:5g�
�b���um
�y}�7&ȥ�ö�V!bS�]x�����Ń�2�N�w^�1}Ү�%Pc���cv�8�R�i�{qx=��ݺ��zڼm�����8Ve{��dp���GA$S���i��|�>���Z͉��K��"��#=��x��ϭ�k.���`��H���0��l�j��>�> ꊧ�J&�g!1n=��߽���Y()��'�Y���h��c�b]%%��uK=��=�x'�]�
��+�/����0�	j��k+Eq���z/9Ge�|���E���<ڇO����V�я���]�FB����c�����é�ʯv��V��s���4Q��(����o-D���E����`U�X��b�~�V��������]u}df���$�W}��P�5�Ծ�����l����[ΞW��Ag?a��J�H�׫��^'J42x?fJ������xC�����^<��ugz�k/�s.��~���ٱ;�|��Uen�!ss�<x��|Ŀ�m��ųY>�N�t����r��y>��7��{���~�x�H2�����\���){�Z�l	����H=���"`Q��[eL�pļ���Ie�rbV"�'�{]o��W�M第�).���
OS�3��i�퇅c[�-�R.j��>T���ܠ�s�*�r�ssz��%5_qI`��3�A݄޺�J}��sý��]��vV-O��(K���D�]��}����
�FM��������2���r�*�2O��⣋*���Pk�l4�S��
��:g6o�7�*'w�s�ꁣP��0�ˋQF:v��ygqS~�V�P�/c���X�Cj'��h�5�EQx3p�֊k]m�zb��g2�0��_�I���iB����y{��k�V,�l���Z�!+��`�b��OyR.B~�D?c���2:�'3��Up�Dnӵ�L�U��8�,�љ�k}M`� Z��L��1q9�՚UO�0��9C�-��{H��!M��������>9�.'�^;3�|��.������{^d<\V^K�|nj�"k�faD�89W�`��Ǡ��2b��1e>tV-+��������g��P�^�r��`р�xiğ�4�9��v}��~����"�C��줥�c+ދA�5L3�� �,�"�KwSE;�������kJ��n;  _��eR0pk��M��p�JM<�x�]a,�r�����w�5��J�`�j�k�����W=%�n���U�Y=~�٠���F�u��t1��n����+-�{R�=7b��fɺ�	a#Bd�4�E�9�+�����g	ͻq�`w3E���B;���-je[�QV9_ֳ��|���������9-p�t��uCC��3qH�C���	}����9擈,�׻Dv8�*���_ns��XM=]�WÚf����qc6�OWW�Nۅ޷�93��i�[=��-����JLPq���5ΒSnP{��x\��u9���kg����5����ALD�Usz{yMW�`x���^�/�!�ە�.��z������TdI�5��.-�&�|�/� r!Lp�}la̱t�낥���=y`��M�?�8� �ߣ���:�P��)发k�����=��j�Sy�\�
��yѯ�ZD�<ǟ"���\�:u�RF��u�g��S�]�w�\�j�U��Ao���>��+ݵN�t����0X9U�l�Ep�/ڬp4D3����M��rJ���k��M��{����)��~�މ��G�d�<u��s
�L� is��9,A�#�s���~��o�Y��"�#}c_�t�Q X��W�x�vTr��*�.��Q.�M�W쳤b��ڑ$@���7�=k�ѱL{k��?c�]n��Gg#ч�P�8@��>�~GY�ض-]_q��;|:	��C�V�J~�g�A.�����0 �Y�)�gK�;�d�\D����
=����_���nE��ᆡ�t{�b$h�]Y�3E;�թ:�o�'}a_[�7i��ή?��*+�t�����wGKyÛ��\a
���\��<y�v#G��m�Mm7g.��t�5$�5�s5%E�{4e�N*��oD�4��j��=�Ԟ�4Y��|>WX'�;N��ם�}Gf@��g���q��7��y�ꀲ���V�.�C<-��ˇ����>2���=G��[3�����Uz"P����Z����ދ<��O=�KJBz�?L����m���֙��!���b6��a�I�w���T�3�����u;���j��R�{���ʘ�p8~kB	օ��J��qw�H���k����=����ɾ�-oؾ�7����x��z�&<5�|j�Sur5�yu�=�]�~�n��=Q_T�W˱^Y�6��ק1�rf���3%�I�	���1]���z�����4(�;�n~���=�H���P3�<�u]t��|�{������IƉ�f v�g~���5��=��^���]�z�R�l
���0n���}a�3B��x�_� �@;L���ʱ�9x��~s� @��#��lH��]��vd�vz�}�&I�����5���G�gi���>�O]�r5���(<ޡ��ϥ^���ҷ������fc쫛F���OX����M��5���|���fY�T#�M]3v��`����Ru���m�u׻�rJ����ug�u����.�sa�*�)���x.oRul׭upQ���*���\���U��Ap��3Q��V$%�}���c���ٻ���>������*uvK�a_t?�c/���+j6�	#z�>xO���6�/O�`��v�E/���w��^��
q��R��ErsV���^*�|D �����}e����7��5�S�}UʮJ�e\����%ҥ���m�q���;Q��gu�����s��;ʽ�����;�MR������[f�g6��V�@�z!n�S�]�n ɰ�WB�}�x�zs��0Q^�p�6������}q#���� ��o�},v%�����J�ѣ���9-��3]�/yu�q袛6�W�UR�����5羽 ��W�OZ�0�9�t�Ɨ��������DH���4O�I 6G�D��ݱ��8��'��C�o~�s󙶭�Hܿe�	�����VGc�l�9����Y�!������Vw?-}�����@C�u26�}�U��G��k��>��Я���+W�����1�C�����z�zU�07�b�E5�#����vK��<4�ݷx���&k�d�23Jǡ�����Jw��ރa�� p�&�ݱ����WZ�M�=+��6��\(��^��L,��p�cV�C�Ϊ��Y�8i/ix���,�y��Q`��xh�E��%�%�*/O'4�Җus��} �s�>�5�\���J�ufM�Gd�a��sӁ��H�5w�FZ��r]7G4?��z�wdђ��-����a����u��;��kcx��$�T��7��Nr�	��ĺd�i^�S,���׷nH���f$�ξ�P�}�k( ���Iq�����e+�Ty�o��:����Ww�s�����=��G5��kI��ؒ#[���EE1�-gS;b���4��
ӼXjMys,[���� :�B�N���ݗ�U��0��6��׉��q-4��_u��������r�`��@�9��b=ڑ����MQ��a��+�ltJN��"Y(�F�7e��������9ke�*kOd�l���w��(��&�+0���S)JX1
Cqgo�oJ�K128m*�+��e>v����+(�b�\��ײ�G`���	z��;z����Yۀ��SA����2`��8�g^^��^��6@�5��v��:���6c��Y�����Yw��+��wg�EuMh�n~����l�v�rgf5u�+C5�.$��]v�̪}�F��v\��U�j��w�S[beX�娛�/_4���uȁ�٧����X59:n,\oa}C��|5��b��1�+$��r�Bo-v��o�����;{w�Ն�z���6*�%��&�K��&��:�Q��j�gh�6*wc�2B�ܬ�'�=5T�" �H�Z7�Vw���}ү�d�\�G�6�m�)�;�Ǝô�TA�Md�Y;�@H��Ga;}u9�Z�r�кC̏M���붒�ɨ��[�3/-� 	.�Ѩ��M;���$W[��Yfv�ل��m��Z�=%�jK��u/��,lş�*�	i���u���<���i�/kc�⚧�ᬛS*����26#�.~sv�J[ˁ�YFU�h�*���vPX�e����Zg3.��{+{��Kat�����POj�Rީ��mm�S�&��7RX���b_�K��2��#��ٱ�Uf���G���)�q����h̟���.�i�u%�M�9��!V�����jP�m*]�	�=z�nq�W�X��8Z��u*g@��oD��W��=<�u7z1.�6����]૜�YW�Y�a���
���1�7a����"�/��lә�Ũ���Z���"e�[|mV�k�`��W"���B��ꬢ%Ǖ�MBoSt�b3����`q�s���h�YŽ!p��:3���L��z����R��Q���u�V5n���Oc�d�7M.��z��S�a7F"!U /�fՀ�+q�&�tC������op_wi�i��2��Mp����2T�f�N
:��{!��9U��-�ѫ�]�}�����L��KK�vV-�okP�6�X�O��n�;m�ܴ�h�/T����Dr�7Gck�!��J�E+���mb��3-%�ʶ�P�p�Q�>�s^fwiͺ��k5sy W=�sa�ngN�j_WnK��U��Uq��G�v>z�u��0��fN�l�L|��+���5�+������d��jݗ^7�` ��ȁ���cOv�YBb�>�?./ {��A��+ߏ��w;s�:y�K����M8/E�CP���[	y>�+�}g>',T��O��[��;�V�;<�G=:�1G��^.���hO�y��G��'��w��u�+�ZhW]���;�6^,'5�3 ߼��ťw����g�P�g]��6㏜	�<T⇏=7�U����i}u]k�|5&g���$�{���-�1�׺�
+z��hTu����EY�_X[�qP�s,c���w:��,���sT"4�&ͅ�����R��Α�<�;3����t�:��P��>�z?N�������mu�q5��ݸ����L�k4[�6��T|*��)<�5�a��:�K���~�w?�5Np��q���tD��*���f6���j�'�u�갸W���<�MP�Ɯ���f��"�����~y�lUr�w/ޔ|W���Q6FU��'����8@�=+Dy����[[���'Ҥe�%-��m�+�{�b��#�e��_{�p0&����s�}6��}�*5P��&���f?���5��MD~��b�Cuχ��K-.�/�Z�ױx�ڼ��-��[|��x0Ej\�]|���C�������ٌ-f���^`TV�ڍh������=�z*>����30E����:Q
�c�[���N�Srs��r��jG�x�u�.����+���ʙ<��2$�f�q*�s5��%������e��_ǥ�ۢ�u���Uvr�:�x7���}�M7s�S^sWb�/}���^4l�v����Q�X�V�	t���g��*UNx矖�lL�,��������ke��W���9�2w�׏����B8�/��<�>>j�cȔY��e*?�x���$Ow��%x�	�ڭ�*
:ƺ����9���^�FV�'�qIi�G8=Qa���&Ͻ&UUzTl����X���mC='���f���=��/5
��e^�{Ҥ�	��V�Q�%��Vn\�Fu�Uy��\���;�\I�T$�zA�p�)H���D�=5��5��s�7h�mPY]҃A��{��<Z����`>}P��̏NÅZ�9�=Ⴅ%�¬�D��>#=}�ؼ�0�U�����:���qViS�nv����P��D|��QP}�6�w��3��t�P�[J�
Ȟю��.��m�}��q�'{_�(�b��o��ܑ��ͧrlZzM�[�Oe���1of�L��:x���^s���#��=X�zir����緉�dV�e	v7v��qkhChԠ�]�Z�5�3�<�Ly]N���j2��Y���V1-�7�Z�!^�����S��L)��Ҝzd��n�{(������Ц��c÷{@�C������h׽���U�����T��r��gN�\�l���� ����ὴ[�/�����u{|J�L��k��O��dn�ߎdk���?fΰ=�ӄG�ՙ$�p�s�tn���>�w���ŧ�}����zQG^Sᤦ��{���޵x�JoK���P���YK����x�5�T�-����/���#�'�3�-��d=J"��
�P���K��v��^{|�uncB���S�pu�1O����x��{��C.�����~뢸s�b�[����;+��|@�
�������/��a�v=��}��Қ��~OD�\/?p���\P�R����y�O�
�VyV�ȅ�n+����5;���\����dYi�_�S"���$b�~YyS�[n{�&}�[Ӑf�E�h���r������՛YyP�j&�H��zH)��n�ee�-^7ڜۧ��Cc�iN���5���=yt��O�p�8�����$dU�zت� 9����tY�9�hHLFǻbX|T��|
��>�3�R��Cp���R������۬��FK��|�sc�Æˡ�"�bYv��3�t��>�S`נ���}
����)����h���)D����ꥊ*��?_�&�+i���v
��PFq�v�7�q���Ԏ�=����l�uz���4�v5p(��ح�/�f����%�n��s ��oen�f��v�Q!�]�ӭ�sbe�q�@8��Y`	���;�g*�	ǽF�$A�wn��F��ɾ�Tt?-��L�����z%����Z����>WWL�ᒾ���a����S}7c~�Y�I���m(��.�3����rvŋ��u6ݟ������_�VD��*3�G~�V��ɚ�m
�����z������� ����8�Ɨǻ��K�������j',�d�QC��U���{���#d\���mG�h^���f��i�x_��D�D�;S=S^������ ��N���Qs�ϣ>]��j�8늟��u�w���u|�Ч�~�d�����՞�헶��b}�챔���9y���΁�<�p.�/xk�>7��}��q�0P�,D�ޓ�~����9�z�l�p�t�/꓍ ��|���YQ�{i�ո���{я��$���^��l/;a�4�U؛�u��~>[���kM\�����=s���aF�XH�KxT�#��/+��%ʋ��?�]�oB;�'Rʟs��Ϧ<!����v�s�v���.��k����^������&3d/ۼ����B+`ti�
�����~|���Q(
�J]��9��c��oOj�GѶ��hn��ʅ^��v�%;R�D��ظѳoB(:vԣYh���Q�r�ͥ�au�f��G��LQgY�u�N�x� +�Lp)´�J���'\ufF@�w�����V̉�؆����\Ù!|���Wm�4k���º�`���V�y�=r��ct0���Ymڇqfec�Tm:��ӥ�KG,ló���Lu��zL�Ȭ�ۇ$h�ʁJU��䮓�
�{K�}]��^�c7�-�⦴�
��݄DfS ���b��nS���0{�I���ίvw��_������-���9�7����[۟>Mw?�Ոw��*�y����5��z���6�3���a#5."������+{� �[�_MQ�i6Eox&q	:+��&����e�ˌ��q�u�Y�$t���/��U�n%���qK<�l�Y��`�9�̜�9�rS���)����!��9[�s�DޯI،�Ƙtm����W���J��ڏ���tǴc#�ؒ'��we���x潄o�{ޚS�Z����{����
v�V�b�8\ )��3o�#�z����ϽI���Y����}5� B��YgԵE�,� ����0�Q�=3����[0�}��q;̦�� {�Z�n},v�)�_�[\�� �V�{�4=��{{y(=�Q�4�ƌ�xl�!wZ�U�EoI���}����{é
h�a�t>6�������Z�}�����r��ݜ��\��w!�ga}�{���]���:5�s.I����X;�v�wbY��먗V�G{�X��6b�qT���������(���>��u�zR�tw����Z���yz�^$e�w}�}1g+&1˯M."`�"#���Ӭ��g���j����5x����$��@R�#�s4��}�WX��`�������&�]6�����_{.�o��>C��sf�O�黉k�,���J�\����yz9��u���+�[��1$o�Ϡ�l�M�.�A&;�����4譍��C/%�:>�hb��gA��&h�U��>����&�4W�'�F��Ч�wP���o�z c��&���V����Z�Nu�
W\t��)&�>2:G�>�л%���oY�0�#O��wQe��&I�����<?v�����]�>��0��m�
T!�w=ᮐ��nbzc�?�LW�W�7�B�%T?
��CD�����<wZ��^�^/<[�����#�����I�D�i�U�x��ӆ�65|^�[�����C���:o��:ְw����i���|�}�&!D��ɼ�UVa�j���+\��8GD���3�خ����V�M	 �},џ}���#|*N+x����FH>Aޮ��b��i�^
;z,�w�eذ7T���p�x�����';���S�~�H�u��dK0[cc4��
����[�l�Y�,5T�E�.��M�+"�$����˾ݧ6��n!,�$,e�����s����#І�w���Ɣ�+�/�=~y`�Ί�G�h�{3� �ۺ[��2�;\_*ZV�T�!ۍev�����h�7Ofo�C��VV�+1����zN��j9��1��Es�܃�j�C�#ղ�۸|G�^Z+�.���k���z����%��9��E�/S7�&;U�1�u���ݶ̇�O��X��}���"�8�MLx�[���%��yV͘��Q�kFm�s���I��
]f׳gT^�k���"״|���KV�2�SyB78�2�q�N������r��Cx��$ݣ0�o:f��Nj>�];�n*,Tl��5��˫/hn:�pΙ��f⩳vr���B���(+��xU���\x��#��֞t}5�Y��g�0��L�N���W������+�yUQ��~������yVCVn}�j��~�����Dxȍ��5 �+�Z*�X�6���*��{-�:����WA|i�q�;�U������2.�xm���N��_�g���h �������7}ǌ�G��Q���w���h���T,��[>h�A�~vgOw�3�#�!&��qG�T�t��b�` K��[�;�mly�R}���Ta�6���y I+rs�X�8������u����h�����٬b��� C�l�{n�R�c�nu�z�&]q/@۬cr.w�7@59�|z9Ji��η��8����׽ih��q���S;)z���V����d)�Z���!me�p�~��n	}Uyb`��3�]ɩ�uTv{ ET��Y&6�)�
w��͎�{){ƶ��
���K�:u�]^��Ś�Aʺ��X���rgI�}T(�1���O��֠��6	"L���1Pn`j��^�>�'sM(8���>�z~�KϨaO��^��C��N��:��{�I��i��w�:U��Y� �����W��nw�;j��֣�og����n�k~
�v��em\]֯=�֌�3|o=[��My�x�,��P<��K�w���š������n�����`;:w(`�>�"8NZ��O�� ��=��u�x��۵˯I���?{?��o��U���W!;x���,T�ُ�c���F+����f�u/>p��{�9�{���Dowa��6�"����쩆����2�ë�T�]m�w�3:e�/MI�s��fa}b�>q�;?�2�C=���jE�(�׉ᾒ���C)��	=�Z���R�����I��7���J���ע��.��i�++���|��������燮�?w�T������ߖ�r���q�/�&�H�4;��^�XB��FZx������-֣�@Ŵ�ArZ)t��l�ɅHu֕2F��c,3�e��n�Z�?s��C�qQW�����3��;m&�H%j�9�Vo�7�+�w2i�@4�1.\�_r��j�NFW5�Hs7�4T��Z����5[ۣ�r�\^�;y))I_N0o�8d���r��K���}t���V�]�{7�n��<�u����x�%�/�����K��R�hA��P�|�,�<���.�:Z��q��	�G�Σq(q���!�MW9�T��a{~ڄ2W���	�zy�2w���s%��Y%���<��6�O�N��@:���T{�;0痓����z#c�L��V��ɮ��'f\�t�+�дuO��;�k�ʺ��s�&)�<����@� �D��^��>�?m���d���N%�pV����P ķ�#�;��X^� �ؽT�f�k�[�W�FN���~��!�j7,r�������jc.���%���g��jϷ=��v�%Q��$r����.���Gϼ�e!�~�LG��L�<.U���T�s���į�[�5��[� s���P��af��jV���׏�@rb|���nwt\G��%�_]%�o���%�jʔ�<>~9�[�W�|,�꽵{��go+�������c~38)�\ˍ��ܻ2�]�D�"z{�w��˞�:~�Yۍ�5\�h>�� *\�]�_�6r���k�i��Z��f���^��3Bh���V����<�,Y5�k��n}R	�v]���F;�+N��cޡG��ch�80;�vL5��a�qBrY9���)�N���������-�C:K�C��0_+wwed��]	 �����g� �V+���`f��`3�Y�}�w8�����oi�'2���!RhD	�����Vu�*��?n�\�˰w��,�0�WV�Rok��ջ<��2b*�e�!H�}���J���`���>�&�su-L���0�W=��;I@Ȫ�xSv�}���/�c��6�3�x2)�>�O��/����Y.�4t~��!߲�c}u��+�zt���L���E������c�.?���۱�N�-����M������2�/֞�rK"�:	� �V�!�������m�����*��#��f��X�"��`<k�F�w�+(�x�WdfKQu�2]	�4b���p0p����.ߚ���̚��e^��.��̛O�#3��}��@�PKO�nV>�j�י����y��9�E^�aE����#�<Igу��Fj��9�]����.g�D^��1qu�H�,�1K's6�����9y#c(�
���WH���g���;f�8�a��O�#wCݾ���o6�)�&������n�|��N�ݼ���AFm�1Q�v1�c!�A��7����wI�=�3��WBM�{��R5 �S�����5%EB[S��AXz.(������7��S�x���ӑoU�gV�k>���+�R�����<J�j�"O���i�"uY�Vp��a ��an�Y���(VF�$.t�!����@�#:�C8,���xV4v��䵶�։X���{Ў/rf����o�A�[�Z��a��ȅa����okQ�V)mǽׯ+ �J�ֱI�jU��5)���Oua�v;�*�\6���]<:b�6��f2��5��\���A,Z�ޥ�]��Ff�/hᮘ����u�m�֐QNw�F��T���
�vE��Y�O��f����*^p�Ů ���I������x�1`�T�}�TEV���޹u+x���/7��88R��k/�م�
����n¶�H:�����Y:�_B����|�}�Ү��6��-{S�V0�Z�YΜ�����W6����:7��b�}F�d��#��{?L�.�ѷ��-+Ř4�x ����x�f�i�/`���V��;3�ߟ��V�C���V3X����2��:44��ҕ���]vȳ4�Ty�Rgw�l3S*���Gf��T༫ηB̼���mN�B�F�S�`���2ȏ-��d���Q�L�q�t�.�8���X�/#!<m�>����{��Ԯg)����è�x!n�m&2�d�%k���q�Chu;�&���fء˪��B���#�k�D+,m�k����CWf��H�n�_R�?^���0G@���|�#�Tox*h��X�gkN�j�yV�r���۩�� BÕ·���I��9��:�jG�6�I'wIj��	=�F*����Z$�q�+�n�'�4&���u�=�`'����5fH��T7����)v�qU%��M�i�9g�_�yr�ܥ�e��j��V] �c�2�r�̲�w;A���P�w3���6���i;��tLcp.6B{�{s��Æ�Gb��묜��Qͦ�U�u������C�7��J�	��E��DѲ�p�_���$;���s];p��n�{t-�ǂ��<�9#)<e�����Ah��d�5|f��x,0b8�o7w��:�N�]�X��U�u
��^���{��C+uR�t�avk�69�]�3��/��+{�B��
ާbR:+w��Ҫ��Pf�Gz��8P̄�͈&��;mqS��G;�~뾼��+i��W���s鏳���ՋL`�{y����ネ�t��w��o�����ŃJ�����r;��R�A��P�ݶ�Q$SN�lU��J���gr��"s(�(�(b������X9Z��n�DMN4�+Eulͮ㣦��*�O���a����n����C��WA�*[Y�k>�U��d8�)rx���b�����u�q� �J�-�����&ri��47i>�����*�in���h�`�`ʼ]1䘡�@��#���\����	£�Q�t��~n�v���ǡ�U���v��y*TR<�D�<�B�ug����0�e9�,C�NV�����I�������@I����b{6ޔ5�E�/So��TYλH�VL��&���Gg����X�t:s5d���f���	��D=/�~h��z};�]�+�
�cko�	2��E�)�R7�sn�[�;�=Q��bVq<�b�����Z������{��|��A���(�E��/���E�ߞ�K���5K�{ʄ�a㿻ރ�䏧��s�#�C��F�s�,x"=S�}�m)����>=
��}t�i�vznC�1��{��O�>�{yl�V^�6hx�:�/:s?O{w���
�#�g^H��wBg)�U�bOa����	��^^ޗ���1C�z2�T`��骗���C��$Q�2��� �2�#��[R��]��j:r�=�ϕ/�ϕ��HO��+h����D!d*Ӈ�3���Q��r{&����L��<�^��*1���:��T؞3����R8o˯o�,�5��myɡ]ul-�ڏ09̓�a^/X�^�W���yd���Tm��=Lt,[5�t��\Ǫ)�[W�^�"AA�#����)Z�I����m9�5,�W���rr��f�e�L��;j�/,�Դ�Fm����S�{Qo��%��\�ȅ��7o�'�b̝pZ[D��u��܎:���e����̾"Uqk``f��j���vDK����ܙٛ;5�ک�5�SEc�:�6^��^��v���Z#z<|}S�I��s��Ex��NRػsplpD�jo\k���
el�����_��z����}�uѻ�����u��]糑c^�#�n���"����d�v�*�9<��2b�׸�T��yyJ<J�ũ�I`���	׍G��6r��l���ɽg���B�W�����8'��(��C=�ߜ]��Gƾ���B?�;|��}���g�W�|�=�gxߝ�r|ޝ�����s�]}Ƌ�)��?]GVu��3���R����9�璘u��K�S.��՛s���nh����g��Syo��0��'�֌�o�ov[i���S[S7Q^�5�[��g��(��Z2���&�ˤc;;��, �z�����q����vUů�o��\�
ޝ2]8�r�."�"tj4�|�߫�Jpq=��_���x���AQ}әn����)L\�	���܃�|k7��:ᙑm����]���+ޱ����hC���dWg����r�T4#�H���Ȼ:��e4^MT%5X��
?����m�Q��b^�Z��N�л��^ٱ�"��U���&m^mԢFܓ�w#$M5���{��6��1w��9ʕ�U�ݧ�L��|2��!k^1:�<�z:���m7ć8�`���ٖv�"���o��s��I�h��m��xe�N��YK���W��Y�R�N�<�S-�VF܂�&�\ٺkMh���j�����u�K;Ī�)g��ɧnh�E^_�rME�!�]gn6�TWo^/���j�z
��ދǤ�y�l~��WTd��1���5w�1�ߞyV��3*Kux��-�#�7жwU*����Wk���I"=|��"�����BOU�O`���-]{w���ƿ\x357������윾��(-66�����8>���)t���� �kGG�W�|S}�k��yiV�Y�g���MW��`~Su���/��ŝAD~����̿8N��c��~����o׸#�=��Gi�:�c����A�j���f�.|>�c�����W1mZ�Q�v](�Rc O��Hj���܉v���3%L��q������(��N0�|tp5���' ��k~�]|�v5Hn�����.%��f@},Oɪ�I9 �r�`l*���y�0D�K�%첬� �u�fed�A-c�C�j��,wU���P��`]W�LupW]E��\�9Af����$���5�XO���'�eX���O,.>�{�^8�J{�f�J6;�ےq��WiZ0��[���hӥ1PW���B�u�K}�92 ��;8k�̑��M��p~L��US�:.s��M��6�f��꼹�A~��0}|wP,��������+`���Y���˝�%}c�I/tc:�:�Ex3�1���To�p"fo�0����Ӈ��n��b�k@�S\|�ͨe>���Ծ���;xE�G����H.�,M�fr��k��<�|���cHDް:r��{+8yp� �﹗R\<^�$�a���Q��F���/{�JO�����w�y�����l����Z,fS j��U~P���]�o�.�JL�4zS8c6.~�}s\�M�?L�<�G��*��U�i��O��u�J
���??z�ljZ��J�ULl����f�tN�ɝy�̊+�}�G�w�]���e~OO�}@��!�m�V�Gй
^�5h�ҧ^_)�^q�����Ar�oc��̬��AE�TÕ��:�-+ 3�~�E<�}��Yj}���K��1��{�t{��<�3��ɘ��7��(������ď.����h΍|�E��O{�@��(�G���W����]�?~xǂӏ��qb@m����eܴ�q��R�F,�;1�ǜE.����WE0��]nv�2�*d�٢�=�c���@^����aj�[�( 8��c��1uqMr��:�nGӯ�[Ys��3�[�$�G�uv���We�ٶ���eg9sR�[��%};�8w������J�I��U� )߇M?zd�;�j��,����}u�v��Fؐ>�U=�/�[���Z�Z%�D���^��H�I�p��9�߽��lE���`R��]�s����#���]���}���R���Ll�\�k�*�xcq����D��k�b�X��g���:����R�w+y�rZ���T?������kr����g%���é�}��PK'����w'ǫ�Jg�ǒ��u�_/����3�C1�e�!Α��d��E:��UO��GP3z��3���}f��U�$;��E���#C.}�T&�6h���� ڂ�#|��B~Z����UV��}���N?�����`���i�V�/��dzyt���԰o���žN�F3;v���ډ����m�B���NvE��Nϼ�L}rr]jO���I��(lO
y/�>�Y��m��[��L��7�=���y\n�T0	���������^-Z�����,�U��Z��U����P��1ܝ(��]��:o�-B�f�q�Z
��D�X�G'JL�o)�-�9�,���a��DD�T�D�u�jW3DaN�Q�I��q-��-�`��p��ӌ��a�#�R�"�i��׵5k��#���T�/��0L<A��Y|�ZO)�r�Z����fC��#�n���|;{<���vތ����^�ub��s��PX/��r��
B������Y�߾�����/SnȨ��=��S�C3~q%��CAU���ivwS�Z�����t�!訟c�;�b���q�:ʗ�Z8IcΒ{bd��i&Q	�����=M+��<��]�u�d�qǧ}4}1�{���ϝw,����*���F3��y�rg@e�M���!�u^�5�>�n�����':0�q�sZ%q�j�#�`��CH� �B/)Z���UOYs����P�L��/�"W���I_+��Zk٨Ƌ�����[�8l?���ǵ��ۂu5�pɺ�Ĺ�9~���T|����d�_�b��)�!�Ԉ����C������=B��U+j�TX(c��l���N��b�q��ۯ��q�<��ˡ�s4�=�ѻ�(�e���f�Q�'��[�)ܮ4�8��>��Ch�FFJ�<6&���~ʸ�7l�5��BbR�Wz��^�3��d��{���q�>��`�K��؇ E������ը#��Kkx`j�.�	S�̙t�	�=yj�Vʻ�-<��D�T�.�Y�_wr�K�$�pts��NY�i��,u��CXᇺ�:����n���c�^��o�q�����̽d.����#sF���7����N�Wb9*6@{��;����}�P�^SᢓWQO>k�=%�{����0��Rʓ<=�������^�)��Ϗ�v���R��ȳ�P���*�T��HGgl޳����yv=H�{ӽ�	�j�c��V1����"*�7h�nɧ���$/C�t�2��:2�}��V��s�_@����n����ƴy��Xl=���/�,��D�Ӊw�꼾�Ƽ(��׸�Ѭ�ׯ'7A|�fr���]{�߳2z3�5�j-�̬�;�����[�Aѽ�uC+��5���˺�rTsU�"���w�L����Ɩ�;��]}1��
�q�$���(�&�N�̺̞y o�e��.�k�~�CwG��O��}C���K�U�Ʈ��F˅�~��v%��I�jғ�){�����ͽнڵ�UOO�M�CG!̈,�"��x��8w+�͉�S�}��q6��O:ӗ }ʧ�N���+�{����������3 �J ���5{~�:�E(���쌑��$��t�I�-9��m���n�]3��S�o�+�[�fW�2��2PTq�F�t��N�ѴuPPw����*Hyr�뺕ݜ��q�j�N���]�%~���:����ܷZgYOF��)l�)��`��u[-+���(�tںos?v2�e�Im�����ƾ�2�<)���X����g[y���ھ��w����j~�������Xjf^a͛��u��O*��Hu��Ǎ^����&�ù~��>�+L59��Z�m{���i�v|���^����qN��ߔ�r�+�O��-��k�a%��=�����o�.�F��}���z$U Ѝ�#��8D��#"������O-�n3+]E$�Ƕ�[������W��Cȥ�����=ÿ�-�3�bgY-!��z۠}X�'ٝ��W�����3�'m�(��f��Y.���[o�H�/�T�{;���������)͇�p��M@��de!���4�4�}�z��>�����f9�Y�Q�.�ؿ���ʜ{c��\��7M}ۃr'���Yf�;7wW�Uݛz2*�|��	��� {q%j�����	<���h����SU�>8� �e��>��ɓm&g*7�gey������"���{�E�^1u����2|����jǂ��ͨ$�Uml��S�{EC�;$���QeSU)ᘵ�q�:*|�6<0'o+n����#6�͠-QN��vȓ5.�����|�Zu��3P�b���w�f��4WB�uۄ
���BQA�J�]<k+nwg�r���ڭ@�يk�ޛ��wt<[�t�9rNe\y�`t�T�Qku�`��]���F�/tnNቮ����ݛ���P"�u"�84��1.pK��gC���V�î�&��`;���'���{d��WW�����R&���:���|���f�ԉ.z�+7����Κ�e��\���%�I��BDѣ�����^���{�
d�֒&�ٴ>}�0�{���{ū9k�\��O۬���}:���D���K٫�U��]`:_�3��Э`ya�x���ʙ��ۧ����x��y~q�Ue	TuG7~q�<-$2O؆���͞�v��TCZ�����5�"�s���'�n�Ǖ���װ��3���demy���\$�͆fF1`������Y�6:�2xj6��G��C"�Ϫ�ɕ.��9��h�=T d\�n#�V�ɬ���u���պ*�g�Q���-"�Nv�s��?~}�����98�Mש�M"]i��n�#��J~�����iF�������\{|��[��ԓ�)5��V׹�f�X,NꊌZ�S��Oh��n�<Z�|�i>����oF(�=�w�Wr��-��5��%� ��&��}�U>�\˷��eU��ne��W��(^�'l�7��\V��]�,g2jr�h�	��fpκ�<ӫR�Z5���������U�"SYق�v>�B���5�j����a�?��wu�c��B^�sr��.�V�k���*���-�Cf9�} Z�M���ThٙE�Z�`�+��OqV�Y�>�!�����f�-���yG��w1���p!c���j	�zj�޳^����GGY1��W�yz��=n_<�]%vf�C��d���}�WX�5n��G{��������g��s�z�����5��=��5�.�
����+~9ϔS�K��R�ޟ�89��ﾗ�?;J�ުt���5S��/jMG�Y��rS�}���4�97�I�`���ꖊ��v�v��tS�mEv��3 �Sp�.T)٪��]��n�̧3�s�څK��AL��3�����mdW��������C��=�˘
{��2��xC��,O��$���x\�w��(U��<T��+�j�����*�ծ�)f?�+�'6��_�g�v��)��t�Q�=�/���v��j�%b�~�M�72�̫�߸�LvC���}J�M�����@T��9ۙx���W$��;[���c�U/e[��಍M���]{ҬW.���g	�w�]Sş��EM����׽G��V3���#��!�Y����/�*)Z�󈿽�E��y�}��9o��o��M�a��(Q&�������z0/)L�x�fI�`�������Oݘ��*��j�x��܆��bJӝ�/�"2�7�}��.��ra�F�e���u��u�f�ݺ��I�ƫ�
�=Uv(�ƞ�d�]Nnb���fI¥M��O$HeV��C����齑s8�b��5Nhu)�{��j�{KrpYC�A٦���e4 /]U�y�%ճ�d'g�[�s)���,/�VU#{G�3u�-�����Gu��鬕3����Wt�)Vvk�|��Ĺi]V�--�����D���^<�S:��r�S�J��*�LkI]Wx��T��'w�Z���Jp�������Sي��S�p�h����G9�gV�Նk����z���5�wqC�sBNRs�ͣ�+iͥ�^�a=(]m�a^�T�X;\��,6���	���ާX�+�_DT�ʦs��O�ΘΫ%���r��!v��K��^^3J�'ٔ�g	�0� GW!�[yK���r��p˴R�m㈫���z���F�֜�@�^>�/rmbխV:�r�C��8t+��z�ru�S+�jv��GS`�;^
ɐQ3s�<*�����Oe;f-���l�2e�ue�F�u�I�U��q�a�b�YZ�u����E�J�I�^�6�X9j�<���ۑT6OS���'����G՘�����ݹ;�x��������4o:���+����t��cB�N;.�Ju:����H�lkut�5^S�.t��ԓ%��e�VR�*Yu�_.Ԧ�{�k�$��}#m�!����u�����L�y�Z��:��wwtm��Հ��
���'�*vQH!Y�.�a���9rfY�sr���&`}%�R���O+)p�֭��ڜU�OI}��}-e#O+�����M�Q�b�씻�®Q���52j[�K��?%Æn�m�r,Ԫ�Jε8%X/5=���\����j7�z��yt�tl,���x� ~�b���b�C��![�-Aqt���Y���r����W��L�
�r��q_�[���T�&Pq��싖�ow��FX;�v`{���E��)[e!�����|'_MDvn̋��.�t���M�� �)�Y�6+pK�9�o6���0*E���Tf���#h����qgv��v���8���%J�YWYtR�x�s2�r(ض�� �s��4.��Wa�Km���q��m�0ou��y.T�ܪ l3�_�]�b+�����rmݮ�d{E����ś�$P��mYd�բ��%�B�ފm�d����ڻ��w��rF�C�U;Y���P]�5�S���J�ѫ��+��7���\�A���8`���{&)f�k��n�Y!��y�54�ѝ٘���x�v�5V8�t�5Cbֻrf�g""���{Ruv�rk�4s�7[�gi'����+��N��ə2����Yk3-(��G�ӄ�hѬ[�^Y�o�	@�TgF/P��F*J� :Z�����Z�pF��sv�N���M+�ĞN-0�(*���z�`�l���U��:8�0�gJ�}�Wu��dOw�ܣ���+j�KI�ێ����J���VĨ��!@������;&�����	��A��Sxѳ��FzoC�Ki�b)p6<b������P5=��˭�����xC1~.�⾹�tm�P'Z��C��O�cF5:�$�����{z��z�`ء8�F��#C����u����^�{~�?N{jK54�t)��Q�g��+��ρ:��ݩ��f�Z��}n��2�My������	=�r5�By�l
</q��������P8�ӯ�Q���e�a�O��F��<�w�T"4ur����D03���Ez�E�̈�h����'<���u_\1h�t �Q�G�mq+��8�K�����.h�-wNF��֭���ï�'��ر"[���?ݺH��V�ث�{4��'����T�(���/#����uYV������s��/���lLi�B�<��R����˵�X�T�k��j�1,����bp/2�����u�f?�Uu�a�]׾�{��D������w���2vx�V<�yް�1s����v�g�M��m2���f���o;��dÝ����|6Fg��(wC�}�_U�e[2�>f3u]ɳ�� �V6egƥ�x�2���%'ۜ�jO^��F�W\ �8���d@Km�}K2�N�<�d���S�n>�p9�2�О&�H3k=,n��vڰ��]ڄ��X���R�2_9�\JgX�LS�-��i���޲(��d,��hУ�뻷���NО�ن���x\u�Fl��܍����Oo�����g�͇��d�Fb�Ժ�fP��B�H$�9�m�����/��3uӂ���G�ý��K��ܳ���7�zNx�Fg��=:���t쩣9�9��++�u�>b`yK,y�蝸����)�AF��O�A��Y��e7��.n�*�S��������'wM�=3�Rތ�5Zt�������;G�j�r��],rT�\'�5uysgrn��6z��{�IҰ^�� ߩdIק���%�N�.�����ٯ6�{v�4~3|�m�m���S4Y�N{����6�G+po�x��elj��.���3(~�W��a��/�7��M{�VaOO�Jm�ؑ����z�><]�A�����<m���nO��w�"$���%8zV*hϞٯFh�׺�c3�hs�6p�,�#Μ�O��r1��8���d���J_(o�^�uC�x�7pDIQ0��{�M���i�DuS�u��?�� ��[5�y�,A �KE�@�`�H{��Ț2D�a{LϨ"�����*�ݰ�}��RM9_�S��rI���e�p��{�#�;B�zzvkCB���UӲ3:hp�L�pU�h}:�������P��rڏ�n�ٽO���ɵ��X�:��w�D�b28�۴r�TQ�Xxi睊�)� �:��VCY�{���(U�u3u~B�r����sW��d�8�/g���+��=�OQ]�M��-c��o� ���;��&�����*���G�JU����3�#	�K'�c6�<�̍*s�䩣�a����x��θ�[]�뻯N� ߶����tF�T��e�
��u܏}�����D.�%W+ %��O�~���!�F6':����5+�����R	�3�gk�R!r�v3Z�>U�ar�,�FM��#�_.���Aбp���8ۄ��u_�3��m[���P$�Q�o[ϝΪ��\�V*B���P���Xm�?>>�������7b�륳��p����L��vT"�x��+��M|&?彁{��Y���B�ՙ���WCP��x���%K��������귧�j��F�Kl�>K���'�&�{�d{�'2��¡�?	̩�i��ʯ^l��=��<n;S4���x���D.��-�x�썃7�_{��Z�;�����s�������ް����9!����#j�EnD�x�!�vo��H�s��,����w�w���;;i8$���T[w�P�p͏Vc҅C/\���dk�SŃB����c�{}�f���������j�$ټ<�J	���y-ޘ�!��+�k�g{c�[/lK���
�1�L�Z���9k{m�Wb׸�+�q��&��#�5�|��WgW@�Q�Š�lǜ���Ko ���2#��P�..;�VVl�x�������l�.�~g������uT�ٖY�&��ҷ"�L�d���޽;��d�>q�(?f@��a25�r�Ďx��*�Ԥ�1讟�6U���3�Q�����hApN	�����ЕW÷߉?�
�ϛ+�}+���D��X\���9�[x}����L�n���H���=�z#��{�r��D��td�VN{�DV��s�m=0��<��Y�!�wP�51�o1�_�E��n�N`�?ni)�q�����Oo����
�#�P'�&dCI�"��~�#f�@�2����3�侔�臽}��{�	�Wrt���s�~���ʅ�M��	y����\�MO�U����)P�ٻt���uuK�����q\>�H��H�T����n �ָzP�Vh<v#����w�נ����E#�怔ɞ����]0�����������DRYJsI��� C
�s�?T�1�����H=ۻ�~�k'�g��|��}C��K�	�B���,�d]����{:���ƞ"% ����ݶ�h������?\	Uѽ�D�j��Hgz�\m�����G���N	��Kn���L�������C1co�v:��K�V�l���b��LeH-�*Yˣj��t�T��`Wfh�Ek���j��od�fR�{���Pu�Q��x[l���@�]����G�'õ3ţ����ƺ.~CetO��������	o���qB�F�rJL6pwX�u�M�B{��!�8?9�Ð��,}sR�Fzy싘��t�S�mq�B����yI�GA���.V��v_fow�aA���7\4�p��M�Ȃz��f_��;Cz]�PYM��a�
<P~�9O�@���95�*~vt]�Y=��M��Rv\�0k�X����1D�Y��}�:>��C8=�T�A��%{�G�D���+w�����?�_%A:���U��g��C�.��O҆aW�~pSY��^����Z5aҵ�?��������ur���>�{ ��/7M����f�1�z� 9iN���e|=]�Ji���S��@�_�&�@�$畳�oTLГ�!h�#�Q��vV�\��h�nKm��Ǚ��)C��u��k�F�{����9Y��p��=-� -����8��5 e�����Z�x�����RPK��<`��:�ѕXM����U��b�8�����Ӱ��^ �Rش�[�<��N��	��K=<}DG)���ٟB�p1�]3�k�X��k톥���,�i\6�	��u?��d-�Py|`��v��ʄ���T���%s� /��%�A9��Dk�-�@j��<i�W���	#9����0����K��@�P�w��w�Rs3`ٲJo;	�wa�hN��E�XV�DI�dOg �R��AQ�)�r��R�dr�$U�5���kjҨ=�r��K���|�h3���c��8
UϵvdFq�ijȚs+2��:�8/8�ɼ���a5.��.Ⱦċb��=�Uߕ����5YaG�wբ���n�k0�"iN�/�+yD��W��qjbu��6c��������E��FZ��ޡ��9J��t)z{���A���,5��ń�K����J�H|S޸�wnC��7�������W��_S��if3ݷ��"'U�2�=6�n/���#f f�3�k*��ʎ���X�V;x��V�l�2�$�y5��q�Ѕ*�z������1>�ڛ\�M��$)4刬��m��6u}<E���/C9ᅚ9`k����b�"�y��hz�݄���"�W^H���ϴ�4�ޮ1��m�hFE�y�u6E;��$f�H��*o{: ?�l{��f%�NE)|f~�[��]N���k[�{K�n��|�^8ҍ���-�B�D��1֤�i�Џ �D�.\�� 3��nSQi@�=����L�J�f/�sco�)�H}o��Q�F"P S�7��a�a���w�q��K���I��,<�
�h�b"FYz�]�\.3"�S��=�ZΗn*},�=#a���YV�@''B�L�IAZ�.ֲH�Ô7�M�"VS����kA�k�Z��=��9�x�a��jk�$�����\��CP��/o�n�(ay�B�\@� x'm�T���b�jH��y�񞫾���K��e�H�<��8=���0�#=�`N{ �]=�s=.�B:XM�@.0rO�Ց�Bm�x�U���v���OO5W�̺�1^$MR݌��-;Y�,��qO]�Os�$hY��>{�J�+^�G���q�Y�n�X�K�&�=� �]����]$�{}�K/��m7�N����)e���%u�$��T�g���I#g�)�3{r�-�Q���k!�kqn�:�1`n�j�z F.[L#��0�, :�!�rt�*�]"K���KX^����9=w��\(��)�6��`��!�W�`i��3��q�w��\Y�Ô[Д���R�)�v�{[q�qmT�9��M�d�{Y�&����w������T�� �7��6�aaŴ�l2��y��oE�n�,ӑ@bk�.D����y>�8LMU]��5{�:�"�(KA�R;�(������9DA���� ud	>�wA�H��ޡ�ЅܾO���+�.�y;%k�݆��+7<%ݺ�h�/ g�Yg+�$xB ��J���M"-�C�ȅ|F�+$�!&X��FC����u>|�.�![c�Ȍ1�n�9Znc׎6�G-��A�\xg�PA�!��4�S��}M����(���@Us�����ߋ��W���-��飤
��<³�{�s�Y��0��Z�œKƀ�v��d�#�(�(����{���.�E{0��HG9X���p,m4�%���� %q��ƥ�q��9 ���8Q��K�"����!��C�^-$I�D��88�U��Q�w�z��=䣢}W�G+�&��(���G<ᰊ�g�<ZME,�g����Иwސ���Z��`עy�m��l�$47?*>��q��X9� Pd���+'(7�c<�M�+.=C�@�P���λ�!ǭ՛$�������\��*ؔRJ�V?Q�A �1��C{�gn�˥�&s�R!�))����
���oD@��ǫ�6���Z+rf���ٜ6�Yo���y��lԱ�Ю�r��׹�+B�,`� ����&11��%�/"R�̮ 3Wm:�{�f	o���H�kyn���nA=J˿߭h�?s�d�iH>@\�\[d4��7�$�Kq���[ހJg����Ko����;�e��=D�n֞��/Z��d�zv@w�鬆s����[1l,��-�D�z��W��㜭��s�"�,�G:�V2�Z�ER��{Q��
��gc%��v^��q�5^P���9�Kq�!L�W��B�@�Kxɡ�k�9R�2G�C���:�!3�O��x��������V.�|�Q��D���&�K>�C4�pq3f�9��D�nP�a��v����ޖG��fdܩǋ�d�v�D܈!�!)t[v[�XYL�9���)`�W��,���CǋR�>$�b�ڠV!ۙ��uVN�$��o�f������Fhn���-8��a÷gdP%�Aa��L ���-dMqvH�:����sq�����j ��\[&
�o����\��u�C��t�Ke2k�8Z=l�""�� �v�L6��-�p=*[
�l�;�d>�$FL�U�hl�֎�{��H=������Q���=+�rK��@�� �z�@��M<7��KQn�G���L�:S6 8��x��}-�%�7�FT�y7��Ņ�4y0y��H�5;q��/�U(AbH�vy^!8D�C�����Aq��b���ᜊ-`�8\�M�U��<t�<J����0wy�-�ږC= ��m0�@���qT ^��S"�}8C{hqj���jy�KK�Pʋ�g��%0�Oc��6���x����sԵ�3u�J݌�����/����8��S�[W�P��=bx�G�s�YJ��`�γ���9��n4�Ӳ�;&��Г��=z�p>���:�v,��nv�
DȗU��;z����w���mh3Q�|�&tJ���Za��qf^����i-���*f���ཀ�|m����8d�M\ [Q���x��MѾ����y2-�6��j��O�.�>L�z�鈲�338-���:r�`�,��-E��� ��H�e�ZX9�	�ii�yͦ� x�� �-ơ�]��=B�PW�88Ge�G���普@���{}c���Y�[�G.��p;Scq� �0���i�D��>.T;2��ų��h(@�q/"H��(��fε����d�6E ֻ"�-��~S��Qm(t���E�\QطspQ��6�E{�Ǽe�à��@N�i5 VL����{�:v'\�J8y|"-e]^Ġ �� �����#�o$=��m,���� �� �����qh`��ϒ��4��Lת�3�K���.dZ*F�=9�/s�w	��-�
V�H�E���p�ن� {]��*�f���(�����!��������>�@]�k*y��t��2��=s�3����	�u�	0�Ȱ� �� �=L�z\!�o`{&�z�����H�@�@��v���o�'��,	%0wo/�����uQ|0��w�s�U �F�l71�NPdcC�a#Ʌd7���DA� ��QrÈ��%�B 2��íPv�͇d� `l�[A�٧¾���̹=1V_��p�[�$��s� H�.o���`A��,��ٗ\� �bIs�Ԝ#HXI� ��D���`e�Q㮅��qn��A�Lz�"����29��gv\X��s�|8� ;Oh;5ah"�[�oJ�CnS�O-�K�(�[��&5 qE��R,	�͆�j󷈠XC1�rX43C���G��i�3*��M��_1k��ߌ=�f_��{��Ŏ�o,�r��ފ�n�+/)�5�^�� ��y1wG��AuA��9}c���%dɬ����vl�c1k��{��R�S����]����L�Sh�L.�|�%���=��u%�ы�ܓ�.�C��2.���Aa�H,�p��Qj��f�O�-3�C'�0�vr�k`x�|L04Y��
� �L��a�H��@�?� ��w�3�8�l�m�x��,%-�0m, ��
�9ha��K1>!��%�&:��Ô��[H�� (�q�(Ө-�żr�&6,����Hï@SO�����9����L�A�6��a�Q�逢�-n��H%S���XD�D��K2s� g��)�����!����P���r
>��@%�a��s�^F�C�N3��|�:�0��UT� � ���" ��C8��%�i7R�[��a�f�[!��r@*�L&Jn�l-P�	$,�H`�mwf��Im�������N^�=��f�a���r �ŀdZ��Hr̲Jd&�����D	,(Q��i�@�A�XGB��b��-��L(��7ɇΘ��D�n��M1�pO�af���ϣ=���j)���\\H�3�w����/;��$r�U� y6� X.Z�`�$-L ��ڌ(vd@� �����!J�$�2#ZA�- �(�^��,<�lq��Mb�\�f	�����,�ɀ��` )���#�n%:p8�^ lU� ,J��XH
!�m0�A��EH@9 L��Xx���g,#]�6c�Ӟ)Z��.�%���J*g���0��Y�H�3�ٙ�5�f�,L "����	�\,�30�h�6���� 9� �5�0�L�@Xe�n�����)v�I���獈�,�, �L�C0�݈KP,��a�L� �A Q� �� �]��`9�	,��e0��	,�	�6!���ɀ��>�a���Y���c9"N��=w&�Y����d,��af�@�A�"H39���L;� h�aV���+1���*�F�w��_v��f�����3ff�� 30 ��0���d `�e�`�@���t �2 `��, ff`	��`�  �`�0fh��: ���� 0�����`�3ff��|o��p`��������������331������0�����O 0����G���� ����G`���7���3W
�L`��� �����`�3ff��C�`�33}�w�g"�D`�3ff��`���v����0ffoك ���������Z�权 ���ğ������f���	0ffj�����e5�f!I��� ?�r 	 r}�"'�7�V@�jjM��Vc�X-�,[Z�jT��я����U�"�*+h,$�*E[32�٥��[Z��C)�h����i�[Z,(�v�UU;�(l��6�*�M��V��b�mbfm��;��ͷf6j����6��m�mMgN:��ګ����N�n��4��u8��-�F��b���eu�KZ���-�D�i����t��kRTt4)%�
U]���A�T{2��[0�:u�B4�)j�n����T(�M+�gA-UIR��t    m� B� �z�T����O������mT�>�^�f����vy�ٍʹ�ם��Nι���v��u[d��{}�甼��{٭b�R�>���nJ�f�]���m:�%J!ೢ�w7l�mh)�����h�M�����_b�;�[��uw����ӻ7�W��UWy�����F��ξ����"����<��(sM��ouZ���{G����9a��{i^��s��f�}�n�r��;�&㶶�{�G<PK�J�J�U�z>�޶�Uc������f��}�{ׯ�m��Op:o���y�7�p�g����{��_G��P|��=+|;�<��;����-�tۙ52�r�����m��SfسB��ۍ:��5P��;u�u���N���{�e�nj=�{�I�'��R֗�^^Ͼ���ΔL�E{�{�}�����T{��f0y^���wS�������&�{ x:=�5�r����6ױ��� ����C��J���u>���k�-���oj�Z�sz���/1�w_\x��}�}���[�蛷�\M��{��V�|��WS��>Ҿ�]�혫�c�[�k��}�]��N���;J���"��fH�ܵ�&�n��[�"���{�;K�h��{���Q����J�we[��u=��ί��Ӿ�o�f^��x�:F������{���H���*�[��羨<=}�+o�������n!W��f��
5�s�}��J����U!�^����E>��޺;�h���m�Żn����do/��УM��
��f�h����ܺʯmw��6.�{k��[�wv�ګ������J�m���Ӛm�L�^��� ��͜}���6����\s�Z�ݎ{i�g-�}uXmm����x��_V�-{�&�v�����k���M��ټ��w�W��O\���"��෽m�WӢ�j�e5�O��ޛ�d(*Aٕ)m�7����E�U蓉�m�o�m�y>���{��ׯ����o[�wm���{ѽ����wn�۞�{V������O�Y��ԣ�#-�6�U۫��󽴺��&�t�+Ջs�w�n���MW� �M�U   ?h�IJ�   "�ɡ6��  � T�R� @ ��%
J� @ 0�IP��Ԙ@i�O�����#�����ث9�?��Hӱ�2��.����O����~�`������2�� P�����
 ���TP*���
 UUW� *��Q�"��UU��@
��f�� *���4 �UU���O����ޟ�<��"Iw�\w�sx�x�����u��`b�TUw���ح��1���wE�(������w|�?\'5R�.��Xvobf��6��+�8���ݜȹ�}ݣ�d�)�Gfn�s��(��Ոg��.ˢz :�!Z���K`댖{z��E���J�4ݳ?cS�p���҉�z_\�'�r�&3��wg���2�-WC�[�wxj�u�ݵ��ʼ`=���B(+g���Pb�I�=p�W�D�ίE��ه(�r<-����)%- �9l�5�"�.%O��]$�*!�:����:P5�Y�(p��-�)�cXA 0��ʕ{Z�EŹ �e��BS��p��v�B]��ݬV��ےq	9��sq�\Q�n�͖�^
��Y��Ɣ"�`�O�δ�^\��7�����q�r� l�Uz���S�!K�GC�u��,ͻ�Z�-��	
��2�*{viZǹY��d�4�Tb��pu������G�Q�J�����6�����p��Wg�ڄ���v�F'��:�f�,��\kF��
�=�o��qw'u��o�7ֻ�i���
y�ͫ36���1��f��v�Ԃ��L��C�f�9��4D�{���P��1��}��օ�FNuَ���Q��O4�aɱcvʺ7�K�[�^Y��&PYi��VH Ҳ鋈SNC1yo5R�I�ٸ��4�њ�
U�Ztk�M�(N��ݥݩ�
9
�CD^rz��q��o��Ҳ�/���V#Xʲ�b=���y8��e��K���E���H�ѩ4���楽G���E87�#s�S[�����V�=	Pt�4�)���3R�B���P�1�;��ޝ�N@��(n��	Y��=\0�����G���f���Med>ӌ�#�~`��sz���ǝ݊��X��M��G�C1n���a)�y�Ѣ� �J�v��e���t�W&��vq�oN�A��Ի����,� s���"�AwY)M���h�Mö�W�m��eW<�i�b����Q P���d�+Q�eS�^z��o�6����^�a�1	y�n�i
�|h��܈o�q��U±�E��-������a���U_����-#����Z�}�\ś{��x� t�WAb�+9���p�gM�Q�gr�/���`�+[�+��<f��엔��x�:�B����g
���Mv��C*��*"]e�L#�qs�V�;Y7����t0� n�]a��YS!�pJ.�PT�Se��5��vHNj(���fm����lu�����i[y[�1��9��w`T���S�T�m���9��?���ya��Ex]�N��NL��"L\�&f:l5Ү�:��eV3�zІYs|��~���3/1o�=�l����_�["��uqF���)=�t$�Η�/N��vnm��+*ʅ;��#��}��1l����A��
j���o�	�2�X�F���)\&b
������l��do>�p��ʎj݂��2n�u],%:�̑yN`�V��� �bB���i
�6���
2�z+�xH���F�]jEk��sqZ�6r]�u�t��|���r��Onj2�$�P�Vz��6�L|:D6��̺ȩ�y|{��\�o����$-kܫ�B�jk�ˮ�y�1`7����;�SG�K	#��#�ר��a�9�:�GSh�ox��P]x\+�')�g�ř���{���Rȋ�ީ�T�;I���Js���
���,�w��vl��4Z�B�,+*�����O�v�/�F듽�qx���ф�`�s,rf6��4�����Λ�j��RI��m��ީNUuX�u�.o2m	Y;3���_�O�{[�4!�#���q-|�Ql>A��g3:��`⣶��gJ��^{-�+4a�T���\j��j�(��{�.�e�g��!ڄ5�4��v���'ϓ � ��68�8��s�pbs�)i�Z?gu�ѭ��޺���m�C� �W�6��)LR��fV2���͓E�j?*��p�7-�����0���*��6�MWsi��N��kn5&�5�m-0�fXz�ak�0���vO���y]���$n�-ĳ-�0Y���,�y���{ �XjKifۣx^����H� E2[}!�Φ.e��`,�,(�z�j'�3mɎ�ХlA�x6�9�/��+*h܍���.[�4��1�f[�*Z��@��*ӻwO�.YQ�n�ykӡ�fn��l�8�L��g�E�4���Ŋ6lK�2���4ƚݭ��;�7R���0D�*5+%�r����:W�8ܼǳ��XG�v�V��:&�ژ�����(̨�zr΄�3n�>��+l^�Z�+R���gH�3:(]����u��k��ݲ&J5+�M���t�z0N���[�#���G�+3Q���Z������g��h�Qa�6�u��=!w�r_����KzZ�@�lRq��d���tnM����I�t.VJ�;h����C�1Cv=Z
ZR�w�+B��&�i���iҷa�n��ͥc��Y��S���8�������𬳎l�Ţ��ȴ��:�C
dr��m�t<�Wi<��s/SW�[��@8p[�#t�
���rVd�(�JU�Qʼ��;���
ۆ�LLl�҆�`��a�j���A�ѓ��$�يO�8]���]L��&?�4ӎ��@�׋L����R��8��fT�Oa �����#U��U4Ez��_���ɓPǮn,-�mڠ�v*jVV�\Yo��%�w!�T�qsm�C�.�D^<�h���7Aa�1�u�emp%��J�-=��N�5c�.l�C��ȫ..������D%�=�K9�)+�hժ8:��| �8yp��_]�U�X�z���Y�x�q�ı�Vq^]? ;�Op�+�a��wx�E���dY���"�G�f�!w�����W�;9M�Ћҥ�{l�r��	�)���SU�CH�w�z�9G�Z\-jYyIQ��y�;N��̡Z����ͬ7Rӗvs".*WӸ���r	ۣl0�D��2���u��ʡ{��忺���MÊ�6Pʛ�$��`̔6��Uqͮ�2���B���H:�x_QGS�6����^�������.$�AX�n`��wD�"���ȼ,�$*Z�WQ'&����T��,;��f��=i�:I�0��m;f��t��o���ᆟ@��CVky.�.�u��J��]�u�T
���2����9&r��S&4w���)�6���pԍ>4槶�u�7c0&���F���2�U�f��-f� ���N���	�pdO[��c���c��w&Q	&�yn�
���N���9嚱�?.��4��v-�.��ONg�\%���� �톆�Z�.��R�œ�-����^��"����oJ�n;�cdX���jժ��P�Ր�,Ky��ؗxn�;i�0S1��Т�H'@�jWwWS�l-T��sn�{Rjι��N˷Q\��s�c��R	���,1Q\�zr��w;|k&M�	�Cw�*?'RAnN�~�ܻ�.~	�og�&�.���I��b�X�t#]+_uu2��7e2đGl'�mV{��4^����qݱ��r�cT2�"hWJR���ݑL7����0����L~{�YN-�pN����)��vS�w�s2���������wرet�Quu,;��=�g$� ��|+�$�n���jj�{5Jh��18�q����.䭋oY�d5����t�2�
�"�J��2����"��lYVq��Sօk��>�����R��Mm�E���G���o2|6�$+@i�P���h��5_g�«�S4|�	�CƲY[�H�i �E��k�3��Z�B�G�w�
��H�jfi�x� 3�S���"ۮ�vJ�l����h��"�)�C�S��v���c m@��^M�k6,*��K��N�Ȟ�_'�XՉR�{YYX�����Ƹ>�6ˍk�
9�Φ��&gD��uYU���g7E:��c���T�|�ӵ(J�e �67 ��+}'*����)y:�����s6�0�u
��������<�ζ(g�պ�gti��K � [���F�^��E='����z�}pس���mb�6��7q/��q6�V�=7���S�C��
�V`I��b ޶˷���j�N��_�?�7�nl�[���pB3ZN��w!��rnѭ����sb�R�F��In�:�L�����#&v.�Ox��CK�w�OnX���W6���DC-@��.�MR�OY��K�/uJܚmG
�.���:�IE���DP��=4̛h�A��ue<dն�����ņ��x2����j�$42,�2�>��u�dZ��fm���*���N�f�A�
x�J�(U�c�D&���(��E]��I���e�JT�w�7%�r���b�r���+��3Lʘ��57AW�xN�/@�œb�5��r�$�=*нѺ��3W�IK�r�T+NH���8��A#�f-;
�ϫM;;�v�j�&�3c�`iJ9S-Zj�w�����q��H]9j��`��ɍ��d���9藋�\��ݦ���f�q+k]��f��NS�n4��da�&$ݙF��hȴ�M�MlD����Q�E�à?�B���JN]�-�]�#����B�ؼ`/�9�8���b��r�8���՘M��0�Z�uX�u�6K�(y�ݬO��I�T��-[�������q&�ĩ]����9��.y����e�Hm���;]���[v��@�=b���f����+n5{V�Ʈ&�F�ή�#@���L�o0�˺�P���i�s�|9�ile��9��u�Or	;;�ز��Մ!ӏzvX	��"�uxl�u=��k=x�	���[�2!W�mã�r�0�մ��w�.«�Ěj� ��x�e���D���TC�U4;U��Բ�ECX�G���$�I�-��=gn�0��Z�b�d7��֏U�����P~�cY�򁷊�܅)�eh{�=wn��}�*�f�Z��ަ2�dN�v����S0WBU^5`K�)��d�?;t؅S��e-�/u��3�ҽ�nC��r�a蟪�y}pѕo �n:�5����	Net��eѼ}�S.Y�1���.4v�6p��{�cv��;�C5!F�I��[�u��P�I�j����Vᄝf����҅��?X#')�4hv�;"s���-�̙���r��(�-QYg��9�=�1���r�Dұ{�hj9y�Y)S���@�C�THv) �l(��/�����8�M�d&�&�Fv�G);�P�@*x-�p>Unɵ�[ j���mbΚ��ը�dl>
l�/8A��i#�l���Csdd0� =�J�������[���̊���{;,����c��
�sD��JȂ��%����;��ۉ���h�Ď�w�-6#%�{I^�t��F`j�M��j������
�{R)2�u��t�	�D��]0�:c7��ܳ/Ӂ�4i{i�$[V�r��������mG���b��+�##6��\Fܵ���8��6yÝ��T�ιD-f�`֢i��d���ʉO�=��Iuzr��J[���̻B橙����^&Ύݧ�X�<z6/�|cw�g+E6Ԍ�Z�'��]�c4n�0�n��"�j\׌�j]���m�	Ӽ`ԃC#��Y�ptMdz����x���i�6�ZJbX�E.;��h)�pVJˇ[w��*;���R��g�H���}f%�������qlInA��CrZxܵ5��r�ԥ�;�G�C�9�C��F31 �K��.�M	Y�?���F�M��'�N��n��/V4��.�S 0�qK����5��������eʑ�+[Ҙw���n�XL�̖��"�ʛ�e�9��6mYd!���ѹ��[5����:F��Л��D�9�)<���Į��[��^�*n�*(-�X-��Kohnڕ�nh��oP��	<��)���cf�X�l2f�5)p�F��z�b03�3;0e�7�0��o�`��bWd�&�M�Uq��I]mތK���� �a�.D���U��J�R�O"4�g���OWZjAZNZ6s�7�ehe;����{J�]'0��hbW,6����m����%�9���JZ�z/Z��9a���#��
c�ap&���I�M<�&	�l!������U�Y�^�6c(��ܚ��R*����Z竰�xq���tA�-�"�<�:�m<Y�4��;7\mn���߳Z�c�3�B/|�N��<�t�Ws+%K�=����a#J떬��V�7Z6�.nmq�uiX��G#7� ;"�xM���xL���V��1�Ӹ���d2����w8������ɣ�ג�&'ap�'��d�C�+���$;R����g����r;!�\w^媇N�*�mMwj��մ�<���ĥ��n�p,@��w\x���Ҍ+�=�N5B�;e*B���T�0�F�M���U���I���F:J�逞'Gf����*ݎ�rc=��tV$'+Xo0�˦���c��h�J�'I�y�rYeZN�� N*�
/o���Z�`zmᆖ�����*q%tД��mb��+xL�on��f�i�9��@y����x�Hv�P#Xq�q[��D�l��_�5��D5�%��� ��BNB�����_	�1�Jތp9:�ޭW�u-5&#E���+[��aI��|D�T�.�9/��3*��	61��nvQ��
�0kM��or���{�K29��g<X�),,]�i�Z����X��p2¶��Y��5���`����@p��,O7�L�sJ�c:/(VZ�'��k��6�wwt�5�ߟ����m��K@P/���z���q e���pc-t'v�Ԓ.m��$o���������l��k��Ͷ䑾��7��f�)ww�6�K5>0��ISm��x;���%��#}$o����;=xh������Nk]I#}$o������G�H�I$g����>�F��H�I#�$o������7�H�I�#}$o���G�H�I�#}$o����7�F�T���>�F�H�T���M߻����ۣ�!��8�7����A�,(��7!et�A���)%rIV�?YKd�~�I-r I"�Kc��Km��GY$R�ku�d,�\�ց�
��L	h tv�)c���
K-N9`IP[mu��J���I$n�m�I%�Gd��:I$�����Sv@�$�
ݶ�lm�`"��K,�H�����rR��$�$��c$m�$�������MiמּD�n�n����s�V�(���U��?���+��Z�5xUhaT�f#��C�W�ǔ�<H*h���ɰ*ye�8���!o�����4�����VM��cD2d/g(&QMk@F�{;��ΐT�������7��N�\�v*���?Q=4�A�J�'jj����p���⸃��5$^XF�9�݅�ǳK]���䫵�F�^���@�ɼXDp�YT�Q)Oo|��&��4b�5�=q�Z�Ƚ'!vck]�NWtr���ɾ�*~�TxํR����6fi"�+�g�=�y'^����7��r �F��dS�l��.��ī�s�DX�L|]�X�+�l�O}�	�ˡm��7��~�:5��G���s��5�Ǭn�m%��b�ڃb��h�@s:=1g]�w�=��34���u��+UA��^)2غ�5���r2H®L��b�撅��v����X�F-�l�j 4��yៀ��U���[�`i]qK��^�j
�GZ�vQ�Z�W��u�X�����r�%�E�u����dW45�,M�{y�b�{99 Y��MN�J��]�N����;��]da�pI��=���v�2�Ywբ��y�>�8�XxJ��O�Z�YI�^U�%--R�-��w[�*��	K�7��(օ\�	�i�.躼���"�ڳK��ʛ�-����J��$�i��iX�x:�>h6�<��HГ$�����p	$�Fű����M9:����[�sU`�t�e�Dm��(2_iLr6qcO���0��%v�e\�[�,Ȅ���ʋ?e�����<����䛩[����j�}w6G�M;ʞ��2��N��7~"`v����0��b���Z��6�7�Ía�)�ta���ޑb���bfsPi�������;a����˻��a�p�`������h���aQ��A����J�-��l)t������iy5��L�]K����V'Dɬbe�/�]�;X�k
=C��!�\;���+�:^�����J��Ԕ�	|�y��q�v�)����V�g53҃& ���Zq��q����v���W��V�w�`��gv�e�0�=��A��Dq�ǳ˵�$�&E�xs��ծs�ҏ`ݿd���w��Mt##F�x}��U4ԗQ�8fr�%_a�Β�2�s�+ޞ;�F�g�0D;�۠_t��7K���4�[�g*�m��veo"��k����oV������XU�h�h�A��p`<��VJ|`�Ѕ��
�Ef\�@��%m��q�}��ZF&�^�Ji��!}��ڧu���n��ӏ�{�p��L�*���Dl�z��cOeq��@�˸bZ(3�T7q�`^�e]0�a�9UI����-˥@&���Λ��m\�h=Dge�M��?��Xuv8���͉)��_��X���R��8Y�׋2��)�b��Q��=Ѵ�	��\�9�M+NE�{���8��C.�6�K(�"��u�c�K���s^��]����5�Xl+S�qޫTh��������],Y4WXw����t�d�)�(�*���s1_�z�gn��"-o*�An�(���/�����ؽ��(�N�a�m�Lofõ���֮N��&��:m�s�F��w�����U�8��;6�S.n��{)~��E	�Z�B��kVJ3���*n�l�+(Ց��M���,_ �W[��B2���^�N�3��"X�ٮ4�9���j�Z�s.�۔#�FK�Z뷛7k2O׸�;��ڟ����1�j��A��b��"���'	7��}�ԗ8�M�^e�њL�xz�A��	�x��1}�Eq<-%�}V��f�,�%m��׻�"hR�OU�=�!�4M��WL&f<�vJ� ��9MK���4�ޞ���C��K�k�)`�� �\Җ���/\VO��~"�(`*.m�!/I���9��( �.�|H��b�\����vܗ#�n�7�c��u�m���[�g�p�:V��,�В�Y� ��ىX��[Nq|�Q��oa��{�]fΤ&���p��[A�U����{Γ�O�8ӡ���ķU�?`Z�0��?.y5�anKgQV[\��4 �S�v�p�h��l˒���H����P�oD�-�G&m%����}u�,�#8���Ǖ�͐l60hw2U��I�P#�Ҕ�̣-ɨ��e�g.����������;'ҥ�MČc$��;���aGؿ_�݅�_w��{��x��R�?\E�b�G��gm6�n�'Dƻ�&1���ð�6�D��M��B�$�a��2�B�M���e��
��3�|e�p��!��i�m��(WL�nN��v�Rl�{��eL�ʝ��=<"ne�Q>�2p��b��=�ɬV�T�9^�cL'��fП= �hf���M��ʗC+hj�YR3ϕ�_�鳮9w�1�SD�ȫ\����6��7yHz��[�4R��5��3D�m-��M1GA޶a@���x#����饊^ؐ��+T+s�ʤ�IN�;�2�S�4um��R�؛�<IP���vV��t� �c��:EG)�¶r��\���+9�+��!���E��CA' �eՁ:�e׋�t��7�d;���Q�2�O�"k�غ��@�"e �p`Hn���p�gz�5Y?s�F>}̇r���<@���0�v5�aY�\��@Ԗx^��~t���mV� ��]g�cÕ�/�	~�Φ���,LVqv!�P��KH��{q,WV��k4��ZQ�H"���6mZ̵��,�h�溠�Y�c�#���4B��&^l�.� ��9̖k4XG�S%�
�elۮ��'q�w;<Y3`�]f{�^M�4&9����2P�wF�e�P�]�n�d�?�s���jɼ����BH��-���
;d��5�ƏlN\�B��聰F�Xg�?���sm�	w�۝=����Ÿ��@z �5t�Ghxfm>���5�`-=%`:�:�y����S�Y�}���5<�-N�8j9W(�謃����B�W=��{6��ל�˨��8�����SݯD[�*�9�!�o��D��&L�0nC���ua!4���'���|׾]�6����=�����EB�ɤ��M{xE_�F��\,��n��H�+[ 5��+�d�p]X���]��v�׳}��u��b��jb��wޞR�n�3V�]�C��iy��u{wo���0���e�ɧ�Ĺ�ta����6F�㗆�9��5�9ƋܢE�+!��n�)!62a���|�$2�YnC`7�3,V�EͲ7:��84�
 T��_Z��6Ni�f�7!/D��7��&�>=��d��se�Hm{��9fl�7�]�홍��B
���0w*�0b��f&A��U�H;��G�f���w��w)�y*�1^$FLB $ymz�e�8֊XPh;_���]����}��Au��%Ŕ�c	���C�@TB<�"Į6t�
���ސ�l��9�v=nE#��xN�K�G8f	pZ.�����aP�m��/7�8^SQ�%�l�	�Nf6J�U�qޭ�݈��	UV����N�Ҭ��p�L�ʽ��]g�َm�3M��帇����M̹⤣e׃���R�۸��.���T\1t��������SO�gZ�h҇�k���5\��ʄ]����l�V��C����N�O:���)�%B�8� �dm�4F�=�We�^�S7Żm�:�H�O�fw9��7V��X�+6{�á!��u�z�c��H1zE��m�r�i;n�$y��,e_�l\�"��Jv��I��P�.%�VN>��=�H���'bg�^z��$=ln+�t˕���oP2�v�T� ��Ѕv*q*Y�+b�&(��Y<9��9�W���-n�l6C2�gn�k�q���P(��4'�YL���p��g�MFы�H-���M��[t쥳rK�k!�7�ՋPE�rcQ7�Y���<��y�	���I����;h�[�i"e#�7x[�&��cƮ���w7��*rF�s.��m@��aJj@r=�mE�?kvܗk���:,D�U.���wt�X��o$��Z��'�-å�l+j�U��X	�,���Ć���ds��+�]@�C���*U,�J����7H��M�������y'�X�FCe4C1ko���P#F��#�2%�2�QΔ�����h�̖��;.�u3t��8�p�k�0+Ό0�S�f�Z:�%2�=�b����y�t����w�u�%�|q� �ɲ|E'nۍ��Ӽ5���<�ҤX"�*���!H��2��7�Ha[�Lţg���hW/���Bv8��s�;g��ƞ2V<,��d�-/ �=��䌑��m�Y�e�nY��WI!�9pl�w��!��mﷸ���4
#�Yt{+TN�(�����H�.[�������xn���eT�9��r�o9D�-G\��(����c��@3�z�n�ޕ6�T���j��g/�NaR$8�fW��a�0�h�CX�H$���c��.��-W�?j�A�f���z�qI��Y�&��(�v��*���Bj��&� ABL�7��{3+l�"PLh��z�e�r���20�I�r�-�
$��E$�=|a#��A��+@��cO^ur�
ղ@$����Z��W(ǫ��T��YT�H�j9���I9��jD�	���:�T�B���1�¼Ȥ2KFꩊE�徾5��鸌M�rV�`5}��-BPe�q�i�o1��ER��n�(����+�"�5���Z`]6���ޡ�7����a#��.7��b��E��A>�s���~���P�ل=������M�ݙ���*M5�!w�̶w����5�g��wcЕ㎦�g3Y�S,ɧ2Z��.�(#ǧs�U3��?u��ȫ���"�`J��T��c��9�;Uw�g�Yě#H����IS2\�������t�.����JC�]:�AQ�IR�N�)�ZD�0)LܐbOZ�#���XoI}k��M4v���O�7Ly��'�y�I2=u�ՙ:)���S�ׁ��Cq��:X�W��8鶒��G����ޓ��W��E�]�
�)r��^+�3�II�z�|��sm�8�??ҭ%%t����+/��l�3������{\Qad�y-�{���u�<iI^�.���N�Y�J���me������d�<O�^������q̑����W1��zw�����8ep��� �6)r�B��V	�5R��6QH�'�]�/�e�,v�=�6��q?:Cl8�^��
}�i���P���,���uh-�.�gI�k�<��e�W��9J���p��Mu�X�+ �U!pr�Me�n�@��}�*�iP�/v��v���pMp:��u��O�� �N
Aь:�?åO����s5R��1�]i������I����K؍䓟&_������]�a�D��=�의����ѽ��
�Ӊ�wn�n%1QBZ��B�)�1�+�B�.�FEH�l��
�!4���X�I���`3�)��w���/vBA�f��*����[�F��P�S縓U��[6�pR�dJb<z���HB5L�0y�ȫ=�;ͮ�!�l\��p�(Y�u�T2�ol�.�'E��u��ǯ�w�����(�e��^u���0+��,lcj��Ś�}^[�#5��}��RR),��
��a� �]�AE���|�y-˜���ӌ�r&O�z�#a`��8s}�=�p#fJX�I�k�7�}�V[=�J~����W	ى�D�8�lj�\5�v`n���`;I��D���"��Ez�/7�� ���72P� ��h��XRܵ}�asK�ۢ��CBkf�sA���ǮF���R�*�� ?M�h���.Ń5�����fYP�ʺi�ˊ�� Vi��E�-�&�V�)IJ`up�uy2U��?a�o5���DMqy0� kF�,Da��C���"C{l=�+.�ҝ(C3��=8)Е��]h�Z8/�#��W��0�ܧ٬��]�'�Չ��@Q#S;�tFĢ/����ށ�6޳#WLZ��x�����o������n��+h��q�_,�s`��.�Khʛ�`Vj!U2\����h�aY���R�W7{!��ܣ�ѯ~��Eb�£N49;�C;&��ZH��������̧X��lh�X
�]ޢ�����4����`�b�_�� g�V���8�-�9%5��R
N��Cn���}
�3/�իn�kv6��<��@͹�n+C�k8o&�?��g3R��zΦ����z�%��P�ܶdnp7��c�˾��l�Z�R�s�W�@��:�lTe�z�X&��"�}�i��ޮ4{v���񛔰���'��;>�qhe06������>B�1��f�1��W�32$��n2���b�l��bF���v
[gC��l��2G�v*�W�������'�;o�b�P����(P�UUtA���P�T(UUU
� �UU?��@ *����{�������7�O{��v�7z84���o�}#m��[��,neb�%U�e�
�nK\�v� ��Ka-��F�d�����ݜ'K
8�i��k㬝�ܢ����ٕ�6n�h��Jܟw�ڡ�y��1]�s��VJE��L�%]�"�����]�(�8z�l9�&�A�S{]6b�rv���L_����y4�.�$H�/��k �z	�k�-�i{#������u�c6�^朔I}x��������0��Ճ�ra��])+���	�BY6p�Y,u��V�u5�ia(Q�Y�0XkS1�E�fL�����YD��7۶7_=�d^݉�\�ٶ��*!�n�.��1;(W#�cD�S�ʢ%҇S$��Hb�N��#V˾�ݮ��U���r,֑!�H�:���L�]x�7M&mS�*�()���ɣ��]P&O���d�䟒H��r�^ܗ8�Z�^�b��Ґ2Z7v%�����2O��e�$Iq݆%��������`�1��vAy䧥�e�Ñ�k�L��`��i�L���2�^M,|�����Yn-5 N"#����iƾ�?ӄi8�Ƭ�ӉϽ-��YF��!,m�*:1�|m�ۏu#�"�Yf�����-���zEW�4��5ϛ�%�ۯ�2��Z��y��J ͝vR�n!�Z'd/�~�W�V����(_t��֋��		J��XI����-���77"�LN5cjUZ�-��约G�vP�en�����L_�T���F����wۼ�{�Gf��L��N�4�;�UEm�wJR&Ĥ���ИMX�*N#5�����m��|���j��]�gvާ��n>C���j����E��g���G�f^����_-��P�M�~����l԰��<ss\��OȻ{�O�:|*�[��M�i����l��`��o,�H^R�v]j޸�3\�CIɱ�/C9��;]�5�Bw�žp�1�W�*����|*������@UUP����xP������8�Jpn'
��������IF�ӓ>a�Q�K�L6��E]"���.�?gs�B#��tZƭ��*����Dڢ�bn�*j��̵�W�����5M��S?�5(�$	��eQ���'d��`�Hq��`7:��/}}��NlE�[�pP�!f�a%a�{#�*��Y��AB	�������/yi��h�L�s����e]@KZ4��5�M��Yſ9����R�b��@xY�~�E�Ж�
�x	v�Z<�cNߐ<"'�x,s����?>�=ǯ�Yo�����W���'·���b��c�+������������Ww�R͍�R;-	�V+`�7�7�ԲJ�fe�K�F�a8�����Ei{���:�1���鯲����]6`ּ���8!�N��^��5��;K�Z��鋻}�I�CW��pW/[}���$^]�
��rCV��xV�-���{	��N���&�X�y��~/�K޵��裕C1V)�{��W��'�b�Y�Rs��y��l���Y��\�[�MW�օ�Bn2ː,�k 4�jur��;���9V��u�')Ԉ�j]+J�\�0_9.��Ia�o8�YM�������г娞���!�T �Lny1^-'���}fmӎ_��kϭ��;�wW;:�ੵ�2!�czWzRD�W�"W-�ZL���򭘼��~��I� �V~rB_;�J��T��n'�� ]��]C?H�E��^;p.T��B� no��8�	1Wc�<�mnc޴��ꉇȰ��;U��w�.�;	*�9���qW��}b�]9Z�Wv��N��r���tQ(xU�gr!q��_9�æ����fR���Ǌ�VͿw�=����|�)�����͈�|B��3�G��KX���3�<p]5�c�{�x,�\*��n*�j.�Jl/C���Fcv�~o/,Q�kI�+�qW�iQ�n���B� �n�	\����y~��<Ѿ#�2pWJ��+gD_{T�-W�=�3���T��^���g�<bx���5�k���ʝ:.�==F��[��˽݊W������P��f�����5x����*}�*)��u�0��U��%����!�2*�t�UQ�k��MDA���{�jm_:����֦�X�{ϲ���"�A��v�\�f��t,�]V_�����<9{�n  ��gs�\���E�3 h:i+��kpƅvZU�ME�E!�z.x�=w:���Y�HX�U����]S��|R��~�-�b��}��V�\�6^Ϙ��N��lp4�A/}Бiys�G��1�^e�q�6߷�Ԗ�5�z�+�y���.H�(�,pCb�u��eH����'��K��R��h��f%E�^�A�#�k'`\�o�Y,����צs�������	Vz�@�v_~/h�T�8k�0h.�ݧ[�d�iە��C��y]���� h��>�@j'|��M&-�}�ͷ�=¶��s|�����.����ٙ���D;�.(
�<Q���a�zކp��Kk�Vg'�<9X��]��ޗC�� �����
c��c��z����v;|?�e�Vι1O���YN�@}�f�_��t˫���G�x$}w3ǉhP�8�ů=�{���0?��^-�'-sF�
��V�P�����@��C#�_Yk�ףe�\h�
�G?DM���`} ��xP�U{��� �����&K��"(����^��	��Ϙ�����.��PC]�G��[!˝�� S�C�WO��[����Q}���^v{_�b��zI-�EgZB�?m�oj��<Ϸ�BO~I)�!�fC������N�M�f���x/[˱Ŋ�ab���Y����u��Uz�̦w&^�U��1^�ox�jP��y� /�J��
���}����Лx�1S��;��G�������s$��^tI�l��ku�� �+�W����<Y�s�w^q�}sy�C�R|�۷��Qe#u��lZ��]��eЮ����y�xs��GV�Q*��r��6�!կ)�ܽ˾p+�أC�nv�b�7ɂ�v<ڌngU�!Gd����ՙ9��_b@yMڱ���/[Q	L�Dd'uW��_y^���@�B��ޛ~��$]�����"��z��yu�[cqx`� ���ׇm�3�}�ػ0Me��U�&a_�rW,�?{l�D�*���[K���=5A ���W��*7/_�W�4�X�����Qui�f�L�-.s�W����w/�
��ř^� �/�+<\󱧆�Da�����"�i�Y���;��P.5�}*G�P�g�!���q��vWス�Q�=^b���u�����N�&�?L���=ԏ2S��E��\�G�U���iʇ�a'{0� �踬����ႊy�u�g2v��{�Q�i�q���~�iy�8��#MPH'x����xe��P�����H�|��Bn_��y׭h���V�n
��;��R�^�X:e7��Y;��u`��Ĭ�ȟ��_v�f��yɵM�Y2ў��A7q��ɳ�	r�q]��O��t-ȓ�����'#ЖD�t�!��W������o�xb�>�\:h�Z�K�UG�sۻ����v���JO׌� =vw�nˁT�F�/se0���B����i�͜�݃����ϟ�g{�P4A�Ij�) ]BGK+l�*k=�'�O���#/a��(��wK�!��\�ٝ�м����l&K�3��%V�,��[h>��c�����-�F�jK����\�ڎA�J<W�:�"'疭q�p�ev��1�1��ǎwm*�`�af)u4l�����/�f���H���R���	��G�~9#h����!��5��Ӆ��p�X
�׏���X<*i�m��՛�gh�]�ם�~z��꤅jj�f�Y�:=��~[RPG/W��Y��=����q���7	uxt�&���X2�p��È�[��J��,���짽��v� �Q�
��F��T�{۽�k�H����'*t��yh��=O��_/z(<xwA�_��G�!�!d�Ѿ��|8��ɜ��YHx�6�<4A�*�o9m��Π�����U��k�۩�Pz��Ξ�<DKڷ�W��G�K8�jU�y��*>W�ə��3yvN�9V`�d�W�Ǉ��>����D=��xpR�_3���mz�B[ݼ�o��<������Y��ם$�(ծ�r{�R�=	h���o� O�c�_��
���C�W�y'��Y; �4�׳���B R�dVF7Q|�N��s�΂#n�,�r�ޚ�1��r�鹂?-�y�n�v�$=�6��$J>��d`W��g�d���r�\z׏�N��
@â�^EW�d�(޹��z����)�l�ח��ڜ���ʺ�#f��gAl��>u�fĖ<���l3��c1����M5ڈ���TR�-ɽ��������ܖc��f:*b�Rm�P�V���4���q�E>`�<��TU&���t>�Nߨr�g�'�e�}���fױT=�9�7��ϳ�~�N�j�I��=�ʬyv�`#�Y�[�S���~�A�uӗ��5� ��p(�����i�Yǯ�J��p��HW[�]l��^j�ss��u��[���ӛ���Uklz�լtǭ�x��r�k���c����u�*����������h
Թ�+����w�ڍ�	uvE�T0��� �6w�������·M>�e]��YE<s7}Q�V0@A�vҦ�DW��xμ5ﳉW���^� �� �|�x��R�6�����	D�����֪BJ @�%"`�>㛧]w{��;r�^WGg�9�HV
��/ԫ�ծ���6�r��^��k^%
����	���,�Q���P��;�����%�f^�M�~YI�dR{��8�=����kH�B�u��y�9�U�����2�� ի����}�K�j�h ��i�E��'��@o�J�C<���
���W��T��Z4.��8RRx�����&\Hj`d�hh�Wrb��۬�Ǵg�p��7���>:����E���!�y%f�'J����N�r�wU�z�z��&r=�w����/�OV�4��1QճWs-��Q�k�Ϡ�k(W���o�+w��z;&p4(��s^�0���G($�ý��6�ͬ������ml����OiP��<�-��Ą�����A1�� �D\����r߂Z�n��l��J��\8b2�t�=m�bN�V�|h��S����+^o�,
�`@P��4�m�:�bP��=�}(�U�<�� ��+.R��� jJ�Q�I�ܿ�l��X:�w�h���̤ۣ�!��(g�iX�.R���#�Ȅ;5~p�.��:����Y^����R����Du�U��G-\���D�jc�*L��(bՎ�ٹ�#�F��U��n�b��W�v���xT�u�;̀N'�LN��N�~��h�n�p�(����oұ�-@���<`�SU���g�Mm᭽n����]��?^|�x�I��	�5W�Ww�e׫k�*\�Ȉ�m��<
�R�!���.��f�+�.cAx�����h�K�ߗ�9=���oR��?q�9Oh�QԽȧ��W�4.<=X���uv��Nx.����Ʈ��4s��.���@Jw�=�XE�1G9�u��9�����"�/'3;�;W�����SN�y6.��f+�,�\7J�[����3�.�vR�ܝ]٪�WF��5�Ǩ�!=͑珮�g�A�6���z�zwx�Vl�X��X�]}��O�Ο{�y���&��x���bϕ���Lҗ� �;���@a�Ю��+Ũ�5]4���UVU(H'�KI�%� aF�t����~��Q����;N�L�1\{�dH���9���^��٪��9�5<x�򝩜� {"�� ��&�Ɖ"�Ac�6�b�b����]�V�x�f��>�V�L���jj�h����wN%����ш�	����Ξ�C2��Ո/F�
>н[�|a��T���P+"��<�Y댎��~��f���MWD�绷;�X�l�^�GЀ2���(M0O{�x�j�h+��<��2o�u�`��}漭�ns�W���*�x�y��%�8珯���	'w���{���c�}q�"�{W��sw����]�Æ�U�XH����Zo���9"$x�n!Yy��%W5���(�G���[���4��	����S��J��7"�0���u�si	Pe"�RCo�c��z
���.t��k$l�R !���T���-u�O6ۼL=�d4Ȝ��Y��=�;SqX;��R�m�5U`6�RX�v�}p�b���Kg�ݓU�װۚ�2��TR�N�|w �u? ��ḏW{�n������ͷ��֭���}όZ�ƕM�����Ɗ��E��VNZ�h�� 赅G�a5�_������Tm�c(����ܽa��Kb�.��I�]A*C��\(D������N��@�N,��Q]hf�O�����K`4����I��g;7*>��%�T���=�X�:�-^���2`;���/&KxʯC�9",AC�ܑ�$�v��'��ͳ�/7���3H�ޥ�]ݩ^�n��x=3<��y@[HPѳ����WX���gu���>��`�&B
��
R���C��9���A���v���g���c=��3��߸�U��]��ms��ZR��v�]�wD�c����8��X*5�h�=�i��ғ�4sB y�{H s�~^� =6�,x��������������񀔜�
�>���b�"��(7�%8E�;��{7s��7@��w<�F<ʳ-K�ۈ��x�����+.��4&3��j�x�uP�2W�9�M�~�Ʊ������A��}f�(�nYYoj���k��ZT��?�y���U&�I'37҉8*��-K�=������囘���-q�,�[����Վ�K����
j�\ �yL5�e\ɞ���������-���
�^4�����ECWD�X�6���	��ĲL���0�^��FMN����v�w6λ��:R�s�ES�z��;{H\�wˣ�ƺV���=���I��Ӑή����(S��]<4,���ཞ��1��v"L~;�o}^Z�~�J���w�-�2�׽�0�ޒ�;@��������鶗:~��+�y�鰳�uh��z!ڏ�f��"�)��ލ
"�NY��L*��,�y����Z���Xřه���a>K�뒿CYz�7&��b����8K�U�*�����o�^��7g[>m��Y���+��@6צf��m��j���Hs��ߑ��2yV��Mٕ)���K�s�x���\J��A�"=ަ��{����_���ֽ��o�n���P���:+|����� �u���ޝ�9ݦkNVTYV�*ZR�B'I-�)
J����?��{⓳u�g�%�Vkκ<�Ʈ�h��H/&�Q�^.w*�<�"�v��"F�N�N�G{��g3�B��L0,�GZ�w=�����/S�B�H�����3(��a���@��y¯qx�?{�M*��˼��%�,��祻ד�FàQn���w�hT���|��M�utD���pe��1�ڪ�0��(c��8�����@���۝ݟE��������:�'ޕ�ɵ��2s��0Z�S1���+��hVT��"5#�g�����!��kjs��%�2�v8r���-�x\*I����X����sFm9|��Nī�19v��u�"�{6p�I]Ewߎ�ìkMgh��\�.����)՞w��`.��#�)Rf��o0ڪ�U��Oڔ�UD#q7O�L���s�Q4�o*-<r��gjk���E=ݮl�O�18����.-K�aDӢ�h�9�-S�)n�2�pވ!�X��[���Y�B��Rgp"Q�y?�2�o(��g[c����e�K�P��$��wI�6_v	td��j�����ݭz����+��N�����T����]����k�\�IWgeF�=sAt;�����=T��ޮ役�SZ��ܔ���7ϳ�|�����k9U��V��o����ǆ�u]��Si�����t{��1Pܳ�]�>ݗ��7��;)�{�8��ֱ�����T@�Z�,��ھۣ�D:mpC3X��C�d�qf}�>�귋Z`����r�u�)����a-��ٜ/.h��rSK�]�rI���f�ljz~�M��"�:����5)�L5���Uk.��VՕie��b͚�)����Zm��r3ҐJU[�w�ջ7&���dv!pL3����e^n�O)<���HȈ��� ���m�}.��u^���:�����.���ٺU�������`O4��z�_�rG�6�B�D��r�������DA��u],�e�ؤyq܊�J�ʶ0�ui�������oa�b�E&�O�.�h�Ӱ�%vɭ`�aU�x���M�k*�6m!�V
n�4�J�Rboejw�M�9���Ԧ�$u��c��8'.>�%�4��%!����`���D���o]�]���xK��G��j�TJ��[�aʏ�Yʠ��1
��m� ��2�+��{��`�O�Y�[���ؼ���Zm�@u�Y��搕gWW[��(�1�qK�h8�J�����wk�� 뽴���9�ͷw�����a�[D�+i�XH�v\���;s=>y����.K��)��^Om�a���χrZ߇��c������!G�6�f��X2q���`����d�ܿ�����a�ElUCOﱀ.�5�W�_m�@|����Z��U� �#���	�B�Sʀ� �]����Қ i��6hf��ڪ��k�˦���Wiq̝��5٘��o\�}a4&�4��#��dP�j��Sb�FM�L�D{��?ƙ��a誰� 	�
f��A�&r%B �
�kM���DG~����������
�k�3�P��u"�4	�A�·��P$�P�fH�?��bnͪ��l�a�����#@����!����i?l �_� B,׌ 2G �D M�s=�;�3���E�1|D B�a� �hl��x�d�Wo�i����:����4	G��"��!�C�j��_�x�UD5�!f��G�A� ��ƶ !f���ϱG>�تS�5��5}w{5��h�N�NQn A�T���/ڏ�����٘ث� �G�q���� K5\>A���C��(�8Y�@a #�> a��b}��'�ޔ�&�3����4'�h@�_�x�� �4�#��C�>�c��W� @dT�CC��@��j����6hG�G��Y�?~�c,�i ~(�����+�TG��@�(�jED��gߋ2� �3{��l"�h#A�^�nӽ��8��^�adS!�U�F�2Mm��*�w�`i8j�ib��W��Oʇ�ރ��4�h@O�Y��C�k?!L�5Zhg��aF��mB/��	D L�Y����?N����ט>��G�U���VZ	�����f|e��~0�#ơ�~_HMS(��5��R��Dҿߥ�V|��	�A*$�ƷB���a��jt�fZ�f�~�!�@�h/kF��w��Tm�=�/�ƅCO� �XhB>�z* �@鮅�>!j� d"Q���Uf�
4O�Y���U�U"MD��u��I|�k"\k��EY���@ Fگ��0p�����U�T#��!���"4��D�@����a�Vh~�ξ6C%��k�S�b�@��@jB�5f��@'HO��X�8@I�#��Wđe� ���<E�4�4+�����|�2l:噻��V�4���g-�e�CR�r�����Y���:������YAhf����"�Wc��n���2wko�cݳ�y�������v<²��Y�#ۧ~���^�g| �Ug�؆���@�BEU���Y�ha���CU�08��,՚If�*��hj��%Y #U�~͹K�P�;���DidS"���a�#��5J��i��埛�ﻦ��~5m �W�8��C��(x��+�@-P�X�T"�ШЮ k�C5A� ��"�b��0�����eO�=�T��%2�$��)a�G�@j㔪2&)�L���$��i�ƾ#�!f��骲�Y��H�?0� K v��C���4HȚ�"���!�ο�!d M\B�4%��q��dT�B*��3�S_���������d��������F��hh@" '����fM5�R5\Q��8�3B8�DW�O�~~s��ɽ����Hߍ�hCL�(~�H�0��#�Ϯ�z-5��4,�u��N����hF�ӯ/ᦀ$"�X%_L�'y����(�(,�"��_���D� w���0�����45]�5XE�&�<a�?$(��L�z���H1���aMR+2�S�������78vx����a�ta��/,�F�4�Hg�%|@gK5C�6G� Fd��{�)����񳦫�C�2)�낽kJ4	�`@C��ʬ�:j���j�u��T5ڢ�K�,2�4;y�j�b���
(Ԋ�5\�Ex���h�j�P�
Ȅ�����b� "��Q#|�5�Ƙ����5�U>����fȿݷ����6g
�P$�ő�ý���R��N������ك��c�)��H�T��*D��W܇��C"8����?���0�"�(�ʀd�"��C�B�,���A�?�Cꯈ�V�{�L��U|<�f��|sw��	S��ۯ�D�	�y A� #@܀x��d@F���
�e�2؍+�kM MBO�����+x�(���&�d�Ea���Фs�*F�'�ݘ�Dq���Vnyw�c�6ap��1ݪ �b�+�!H��,�>(��H��S4�W� ���~2/�@@��1C�q�t����4���P�~��b���5Z�$ |hiQ �@=TMR:hn��p�*6�'LY�СPbcg6.�%���T$&���|k���ȴ�F��·iޭ�7����Wz�����Eހ,�v��}x�G5�x��DT��,7l�H�^s���F�����H
�.�n����0�� 0��u8�A�R�DVi�%�C
��(	փxL@U��4��Pu���k�r��ҀB�TE�`������wR0S%���I�^�X�(��Y��WZ5'�;Z}��S�s�qW��F]��'�7��Ћe���c�9#���EW��aZ� \	�a� F�%���Ǎ���B�Y�~U����(h�L�G��*�B +ȑ��CE�K�� ���F���,P&���@����B?Z�5���_Zc������wզ �oΪ$5���� 2 'm����e �3U�!^"��C� �����B4�!����H�Ҡ0�"�G��:F��#d#��,��>5f��&k�ʃ$���g�ǋ΋\�Z���tDEJ��Y:t�i +�zA�4 a�y� Ek�)��_��M�f�J"����WƇ��h3A�B��"�����!�Y;�v����V�l	����o��Ԟ��"���M����2�}t���W�o]*��.����%6ɗ��Y{0�y�/�{L�̨�f߶�a�F0 �Rذ|7ov:{��/�r���fg�$iU��e���j�D��E7^���B&1�ʺ�٬<�|7CS��61@O��#�3��;&&�+�6h/�(������u�����\}9��j7�;����|l.|ny�+�
8��I��&�����6����,r�9���y�]��duR��z����Z=A��2QD�csi��ۢ(�̼u�-����rOߗZ�ژu}�f�$��w��l,M�H�s6����;_�,�S)V,����,'�
~!m��My+>���m�����(F�Uo6̣=���v�hy����z��a����2��F��2,2yV� ��nM�D0,"�����'�-���O�~��<�y�g:��w��lee-+a-����K�Ŵ��W@�qc[�M\8�S�ҊvÃ���\E=��)2�f�l�u�m�'+��B��Tݥ�r��1�䍪+l��㑓�g�������筪�����%�s�W*�Q�oE�x#f�3� ��]?m9�st���!X,���I0	�\�H��Ұ@�3k"�c��L�5�����=5q�,9�2�J���r��k�{¯�v���1&(�j�oo����*4�Am6`Yq�X���P9���Ml�JA�x���Uf-���غK��p@�ʰ�v�OFa't%������M��.a�H����謩 ��ƚ��;�����gp�.��\N�5�U0bN��kL����ޭ�g�j9}&�\p=����m�=U^b��ΎK5�h,��3�KO;8���!���QiDC#�P�&�lUFb�7����|
��c,0Ì3`�Q\�	)�A��0�;u���vYI_��`ֈeO���WI�>�F
S�2d<�n��=%�9'�M�=
K�v��Y
���?c�j'"����̅]9ÖŻR�����j���I��"v\�5+5�Q��G��u,[����b����,�P@h)M��e�i��y9����]�8�lW:�#�V��=�K�>��i{�����pV���Q!=}�+�%�K$VL��~2ɯ=^�9Uڰn�؉=��gz�wwcbiy%<F�hr:��1p���j���4ԃ�g/1P憇�wp+���hfe�/�ȸ{_-����d8�KE3�4�8�ʳ��:h']V���%:͌s�0�(��� �o��������M>����W��٭i �~��[�&�M*@c�&�3]pd�Yi�[���6�\53e5������eCq/A�e�9�0n���cLE�!z�?%z.�{������������}O�x�/!�hI�������X_9l����ͣݹ����t�.1�����Ϧ�}��C\>��8�����O��]��],1�'��v<8˖������Q<�]AXB��슺;�ȇ��ʏa�~#)A36�d�c����މ�	�
�GP����E<h7�X:��ҝc���ěShT�z�,�l�᥆hRԯ��ܟG��y_00��Vmc4vÖ��n�����
�����s��Y^��8f��3�4�I��W�g-�l��l_;l��W1 �gMiɚ�����᛫o�Z���ڮ�E��<�i�z��w��߽� �Ώ�V,�@k+V�b�	�z�N��b��0���<i��Bݿ��1,ѣ=/�V}�8���IO"@���xp��/�ss��3��k
g�Vj��;�&1�����ׯ%��)�L��wm�j��R�W_����`2�ޫ��bU�0��n'��/�ֻ���9�Q�ȇ���E���GG[�yY:��˳����6�|��Lp��cO���]�;[Wt��e�y�ȥ�\�Ǜ[N��@�;x�j�R;������|_W���6�3����:�w�o�I�M�A�Õ	�>��}on�w��M�ʌY�-<w[�ҩ�u��\���#�r>�X�>�l��H��掅>�ZN���+˗0���$�Z�/��h��G���ACC⾴@��V��� ����+��׊�B5�\�p>��`��~��N��k���U�oQ�Y/�R��ha3Q�)��2��oZdՠF�qkT�XCE_ml����]w���3���l;�_���9-������v�s� �qd�a���z������[�u�>�ڶ��l�+I�=(�[��7l*��4D��О	��{{�ŚZ����Honj藾���ծ��i���>*N3F�5��1OѪ�"�2�؛�ɚv|gֲ���=�3�9�_t�0$:̗-�� ����E��e�3�9gd�A�{����s��+�3�d�ɺ<���ٛf5<��}{'Do@J��V�Uymr���.��휼�,�t���&��sI�λ�_݊�O��vEn�=��5d�^R��~�yQH�%%�'��u����NG!�S��y��`ձ�hn��6C�[�
�)M��ڷ���)�i�<t-���t��gJZ+s&�D�Ų�"��7��к��޳a���8�|�*�vT��@kw$���6�?!�_]�Tr���溳-Ͱ�˂ڮK��d��}0�Q#7��QJ�M�@��w��r�X�2m��N��Q��l���0>u�֖GclVZ�=��(�U���Qs���{��'��W���0*���=dֿlߘ˙ko6����K�����wM�^�hc��
��j����ַG�c�d�
�ƦuTW�D�c����z�O�:�W�CPz�����¹�#�l�a������!U1�;��6�nغ�o�t/�b��������N�=�_n��?��`K�6��3nO}���u�}Q���c#���x�n�u1��ʼ�k�!�x��;?��ie=�j�*��I��B�O*2�*�����ݲX�zbv�=s�bӮ��p��b	׻Bs�;�t�4��O�	�έ!�i�g��
=�`�e�^��~<h�P���͡qم�Aus�b���]��l�Y刅cX��?Cj�(~�f��I0b!<b�l��NS~!�����~>�R9��'�NU�E�xM}V�0lɰZ�QQ����`�s��ƦP��޸(��k�0�Jd>+�	k�߽��h1�3c�j�7_���|xҮ�[�U��٩�:��<ʁ3w��I�R�Z)
�F��i������e��<*���a����ʠ�<��i�'�c��&�J	F<���P��J�������T*�IH���0l�򓲁��Yo�>_z�8ݵ������<ؾ=����T��	��]�~�2J�8��Hx]pW��<�qs4/D�[^=>�-��4K*e�N��P���5�_�����O����%�8�n��i1}=l�׋����I��T{�|ߩGagh�Ʀl�ַ��='�^л��B޼�F��Wlk��m7�n�Λ�N�Mj#��euc�x�w��y����>�8/���mp ��%�Vw��@�vT\�XY3R�z�U^T���
s�^0��|Unn���pN�K��:�DVR2��s���r,�˂\� �]��.
*��ە�M��ʰ����#���Tڮ����w�X�"�e!�b����Fok��fq��i�h��}މ�۵�ErqҪ/�h�y�tr�d�;����~yXI�F�YF�ޘ��5���-(����Q�-�Y�o���R����?�������»�5ʯ�̂���q�{:l��=U*:"�G�ټ�q�ם�]dF�7ka�`�!�	sۧ4-���뉮}�i�s��kΓ�� Y�����j[�n(��N�y��S�L6ӿ]���-��R��M}gkwײ��άTߐ<�h��eA"�^��ëz��N�ж�g�yY1;����q�f���^�(�6��f�tzOg'S}�O��_c�8+��x�@��mς����7�ߕ�{�O�gX�ؽ�VZ-}��5�>~_u�P�4*�pr��g�
��_���L������Z�uq�Q�<�烍�)��^nݬC�i���^��F]�N�LY�>=�����|ˊ�Z�uB�.�ķ�xNO[#��޿���e���v�LU�vC�G�:�ow��n��\�N����q�x: ����be�{1*�IVs��x���eu���]n����X�W>�OV��Pm��ӂ��<&���3��ۻ�l��;�Q�KkM.$��Of�J?W�3�v:;0x������@�4^��>�$9̳�����\�<a�ܚ���g���	��������^�K��W.�-�(MPAY"�����Gt
e�z�=�ii�&v��
o�c�qm/#p�����}�oV��y���4���Sg:�B��AwVvӛv����]s��������M4Jْ�X�Qx�L���=�?��%�m�V����\N�[N��n�����j��Q{J�OVl�	r���^C�KM=J��E�Ͱݚ:-(hz�����{�>�n�����ޓ8�_� {�����1���~�>�/ c�;�=�j�����3O}Yڡ���&p�J&<.�~���:�fa������\*��p+$�C�L�]f�	��`�/Y�G~��}��~�U�P�>���0ͅI��6�m��iަ�h=_-k n�rl��KZB��ߘgN{=\�P����I�u):�x6�`d~y�6=�
���X�����t����=6$z(q).�C��ci��TQ�6:\י3%]�ժk���D�cq9�mL��[��L��Ҁ�H|A#�eovYWfU�}";�v��n�L]�XF�����λ}�N��� Z2��;�f�s��`;�xWLރ)v�b��>��z�t�ݭ�ǟwua��n[��ɂ�n�5���ۭJ��3c��9b��Sg��\_ Q8���~F��@J��c<#�Ї/��Hy��J_'��M˪*6�pZ�[�^9�W1��F�J0k$0}��
0D��5��%�)�E�R��0f+���K���L�"4] �P�� 2H�L�f�f��|�Xg�Y"�篌���V��k�Eݣ^R��87��m�p��F�{��O^ �4h����+lr��c��"$#n�U��e,G7�'^:4t�jA-ܨO���L?I3+z��2���ֹ8���6G�"������|������K����1M]*yv��X���_QZ>���y�
�}�eN�=�g�۱�%	�%btʗ�3���5�`��=˛z�����M��f|J��e6��W����߮v/�CG/�\��{�����uka�fs�1� �g�M�v#4RR8�G ��ݗ��чt�^�S�W�Lw��!�(=����3H[�t��4·)�'7�_"Z��]D�T��Ňz�HL�Gi�Xtx��l8R��3
IC&�+���ת#ZnTa���S���X���;�����k�ǡ�#�xK������C�MV�Q���)l޸��|"���+��v৶'��t*��XoG~)m�G�w\8����}a�
P�*Ѫ�W���f-���R�JS�o�Pξ�i�n%�8]�*����̈l����Z\EX�pM��J]�j;-]����s�Z�4S���r"f�:ۻ�br���r�';�)p��!��}"[��v�<��H��;�dҝ�W�m!D��d P��վ؛�W��ht�3�ܢ�Ш/��V��#��;�莴�B����8�gV���^*�*v���!8
��������a�wvDݽ���p4)N<����R5v�Z��I6ʜ���wR�s�K����Vی�W$��Z�C.ɋn>e7��ޖ�%Ҙ�@� ˶�jm��,�IhS�@���x�n �vi�iuo Hn�#�1`�yl�u�TW�*�'��G���W��E{��Fh��D8�*�a[ro[=S�(]��>�A��:�w�Vu={�+u�kb:�+]B-s�}a�E��rR��֊+�Kp.��:+�[ǖ�UՓ@���[Qob%���[���+��\��466Ff�;�슞ot�N��z�޴Z��w|ۜ{#Z�9����7�F��j�h�=X�-�Σ���8��L��.�bKJ4՚�f],�l�u�k���F��q��S�2�����N����=<5:w���J{Q$���'oV	- 2�r�Wn��݆��[��;����.�~��iX�g�A��/��w�̧�}���C�n�e�;�����G����ǃowo.�i�%�,�v��m2��HD�P�� �����,�b��)X�&
~��
������.����!����Q�?V��r�
�k����[�<�w�RC�^`�{J���C�,�[�󉆱n����e��o�L��ٍ#u�m>޽؈rޤ�X��j왉yNف�/d���h=�����3��e�$4��jmKp�9)a��N6�F�����*�*�`>�~|o��/vئz
�/��C@�]PP��:�<L��S:#[��ǵ�كWm$�F�M��y¿!S)�Ŵ�w��T�m���f8g�)䥄���þ6h�*��x��x��ϯ��FW���7�,��i��m6��Gd�j��������gm-#-mrd]׌�JJ%�l��0:�`���V��O`m�f�=F�C:DSQ���G��"�"�����!@�������Z�N�Oe���b�l�"GK[j�a,�7���v �IMHNWA���gbxU@�"�R �ZIC4�n�wd!�T�Ϫ�1f�j�`���~i�>B?O!�����Xrd�
E6�t"V�,|���z\�M���Q��v!�H�Ja�5}����S�_|]����kU�x�U��k�jxՎ�XbFu@����u�	�&^������z�v�6�q� A� ��s1?7�u1��9ۚ&�1��u�z����!S�.i�gZċ��ѱd?Fv�\Ÿ�����C�#b�n`-����Ӈ�}a�O���[,��&G��4���7<��NNw����yKi&c���o;T����ɈO<>���f��yC�$���U]��S(s�
��o�~��(�����V6&91�R5$��Ǔw�;9}�{����`X�ōwWP܌��:�cʳR��|b��3k��R�j��e̱c����p;�i���J���|��۾-`,QA��$ڤL&�����\�)�R��G��r]���[\�3�Q��'��< v��OJ5l:J�AH�SJ����r'q�~�O����V�FK<��vZB&��BG�L���`܀��֥��n�dk�?J�����N�7�O�"_<�Sx%H�~~�<pl�dlfA|du�H�I HԵ�݉��Η/��v�m����VY���~o�be�Ӥ^�}�i��9�F���܋T�`�f���k�G��0u�k/O���|�Z۽��u�����y�4>-���g0�}�����3(��|��!���S\�&�U�����ޣ9��^���J�Ϋ�=�3ph�a�
6�#�Z6A�t1�gEC�͞�،�e�M�&��vڨ/j1�>��X�l��{6����BX�v�L���֮ݚ��� ��<�:�{=� =�u1w^�^�:hړc�YQ�qx�曨}��&�\9=�}��z�{���x�TǕMK�|��s5�u{�y����NE�Jޕ͙<��+OM��6�������kX'4�3].�5����b� �01�u�:g��'�e����C�gs&S8e�
�I�
[Z*��~���T]�[���{�R�!q&+.Lr�_����;��J����a^��u/�þ {�b�}���(}�@טg�(D"���M��chd�N��s���>����K�-�ϫ8����q��?48^<�9�հ�;a�(B�k�ˏ���[�m�{{�[�{���埍;��#���R��ޯ�bf��� �������,������܉�5�#��7�Ɔ��I͡*��|��v�8^��-�rt�N_3ܵ4b"��mm���L%�ݸQ��-��'S*���1f�:R%맼�s/�!|�x;o�������;[2�K�������w����ѽb��<#�����QI�}]�tF�3h$����[-���Q�͎̚ˍwM�-���K쁹J�V{2�S=#l0��ݨ�^�ef�6����w.�pcK�M�r���b���R��C�2 ��k*�2cM;38؁�{r���@??@����/՚C?\�!W���]j���-r�P:�j�뼖�,�o�,Y��f�)���f�r��LK��=�������	f\DZ,^�8�1�bA�O}K�L����e	ƻm1�'/ne�ۀ/�}g��&Uc.��^��'8��ᱢ2���w�,�\����:6^��z�n�z)�ef稱�U�FUˠ=��j�)o�p���W��T^�{E�>��痛��ݾļێ$WUw�c���B�$R�d�K?t~����uO��W��Z�n����E	Uu�����WRߟ�'O{r���O�w7ڸ_����T^�q�]���|/�fT�@��i�r�$u�:��1y!3�4$\?�[6,��^N�t�c�+B����n8��4n�wV@6��pk~ʆ����O�����H\�1�k���(��Hϯ	���ә�v��3�X"r���*�V:���(�-�τT�c7b/J��^�O|���h0�mr]���ƞR�jƇq܋e�uU{��E�s%7���hqs!�z�<n�,W�fe�$�r]u���F�W\�5�@U�4i��abhýf�{��H�9���۝�3�{11��{9�4�ޥY�Ov��*4*�=(��K��ٛ�z�=�E��H���y�p�Hgz�0N���:g�1���G��2�:w34]�ϟU�o�|�
���D;��db��"�[�$�6xcl�B/h1���)�*J�l�X��"�O�a��r����Vz �b��1ƌ���{�r�3��\YӦLB�jz���R���RY�%\����C|k�������L^���K8W���  W�A�k�^�UNr)4�؞��W��X9���iBW}a���w���+�&�	@��{wǫx;Q�Ј���qi�ICI6P&�i�_s���̭��v��w4н������E��C��c/*��sOV�Q��P�=8v�H�x52��z+��Kn^�9����C`���P�gp�;�B�b� v^b�r�6��Q�ɮj��og���}�쮵M�%wY.��k&�7�����W8U5`�k�X.:��7�����a�21�C�?nA�:��p0�|^&���k��s�d/D��pA��j��2��:�;3�=�r��{�愑F��s+��׋p�'��V��`
4�5S��qn�ؗ�.��>C�y�*�߮P�~}�|6���ji���H:Xôo-�T\��&g1�5��r<l�(B��O8��b�~m�}�3-	���E4���д��X�n��|y��ϫE�.]�(5�-,�yl�N��F�c4��$��.���ٳEݻqh��͝��xgN�e�(�eI 	�ý��k�������i��e����T|��9ʲ@U��۶L���]���_<;}��MSw�5��Z�<�@�D��M�0�f���HXxU�2���H6�of5���x�
D�<f`�}l��0����YqP���:��@B#9���s��?���{,[K}4,s8QB!��S�)�!�* i#)�_��ᐚrcxC�W�Ĵ�j�Dζ��
W��g8�0�D�	�����r��Gx�p�������w����~�j4St;>�*���K ^�N����Z���f*�M��#����+�Hh��������
v�F��k�xMXz�zĹ��k��K_$gX;���
1)�N!�IJ�[C�e�[q�1O�~�%Z笘��Wy�ŉM��b�T���O�y�,�y1/����G]�n�Н�\�]��a���D,�řO#<}2�ܹ���O}��H_ݒ<���R��ϱ�En��ƶ6��*s��ڵOOw/!��M�MK< \�®�5��5�0��	�57�ԳWY���*�����F!�b\>S%[	b��E]�����ݘ=�� ���[|<mQ��н��j�yz�ƽ�@/��}^;���O���v�H������ݱ����Y�ӄ�X/�6ʝsY��{tT���Qޫ�J_t2Wr���yY�bź&�h6IrB�RE je�p��� nԁ�\\b��̗4T� �������:w|��,.L"b���e"��u�I[i��BK
O���]E�;-@3�(�b�(�Y?����9��ys���c*h�������Dz���/o��M���"�WtBn�X�ѻL�*cv��`�NWo�}r}�b&�%,���X�y-���~�V�wc�)�P/O�`�c��=m��k�*cݱ��/�ɤ�ch��F�C���܊�0��Vڲ��@�I �́�r�X�R�t�Փ�ᾦ�e��r��Řu�/>�W�2|;ޏz=�����mV��U��d���݁.���|r͡1U�yw7"z
���(kE@^fEy���u�������J�3t���	�v��v����ި�(p�����ɵ�w�c���<�wG�����鷅Zq�f@���t��$vfK܆��I��F_y���V�smW ���Y�i���JSM�1���RU��1��hN����`��\Y���w����r��R��5�Rn�#�27k1Qx�k���n��)E��&&DhV�A�h�Ywx�r�R���B-،�4>�Y��B���p�Ë"��j���=*ם]�t��SE��lY,k��\�l���E����앫!�

�s�bܜ���S�6jlܛЦ:pvTD�l]G��1��'�����Ү���^�Ҏ�[y�]��h�{��[�8^i(�������.�90&Z�3��j{�,���)�����tC?kCX���[҅�t�6�0L�L�\6�1ml��^9�㭧�Vv=���������}ٗ]�Nx$����,�����g@$�����ћ�:�ys�]/��7x���^%]y-�n�+��{@��^]w�z��ߗ<3��ۦ�;������孜;��*�jj��!3Ꝩ��v�m%69�M��ls"� �k��mxj��/į+�S��v�~T��t��hߗ��ui6Ñ�������e&ך;as�?��n(�m�d�vY7�=��Z����EN2vjw���	�o�m"�M��l��mOc��k��y=��'��n���їIݏa��5]P�}Mؔk76<f)q��roӊ��iJ_ x��i�o�c��W�<��e��]���
Asw���9+���W����MR�J�(����\s���ܣ�m�+��ߒE�Ir[����*�8����-M���)�Y���e?���%����!7!���}|�g�&�Lи�����>����.�3�GZ�V}�Ļc&��Ʊт��֭���Ŵ"�֨|l.���R�P���
RhNk/����h5�w��F�����ܟ�����J�g���3�O&-�u�C��Vz�l˶°Zm���l��%�*wsD��p��Ŏ�A���� �׉�[6���j��"�!Lt��v��ZꙎ���_�Hxn�-V��U+���D|qL�����CUܟ�̀D]�Cn��K*έ]�W^Cr��\��
a\�B�#�0%�M�Z�\�sZΈvs�d<�V������`��齼���=YӳG
�W�:��{{Y����F^�j~�a�9a�x�����<ҙ�!����Ly���ϳO|��Ox�~��ŮΏ�N�TWI,��O�]":�v]�ks��?����^̛ߒ��@��������wҬx�Ιi*�����J�ϯ�(�M��n�ڵ�B��X3E�e���l�Ө+��}S���f}��_:U��|/W��]z���T�PiQ�@*h��2J���WJP���=/�v�����gu��MD\�G��<�,�8*��T���C��`�c���q�����:�Oy�Y��lT�|L��vN��"ͳ�nK.u�J/1�f^��Y�R�|�bg��L�!fig���]@�������C}t����uӏ"�����e�|�R/�pՊ���޷i||v�h�p5��@\3��'���~�rC�NX
ط�Om���Ջ��r9����{n�aTA�������3<nL��1�ў�:w͞��j�¨;"���ܶq�f��|7���:��Rq�:��
��׬pE�q�4���7��#&�L�&��x�����?<�W�=����U��Yj�E�úF ��D§wˬ��龧�(�2z�c�ƃ�2� �jy��F��27���PV��8wptV��)�쵦�u�\�X:�ٝR��`�ࡰ��4���w�����o�
��e����vgp��G)��۫�gV5у�EB�h+M�K��w�5���[��}�U�G9z��٢���on*�ґ���=��:�_ճ���fC"+v����z2J�?kLQ�TШ���왚�c^��͙�j�.G9�Q��YB��V�;\nwU�&�2�cISR�*oS�1�(^֫��G��F:��Z8[Ak�0���nʒ��Q�5�.�@���ÝP��J��D_.�����A#�����{7�:�}��.�}/���<;��lC\;_N��s�|vRn�OL���[�ɜj�I�T1Oiģ"TN�N��cڸ�Oѝ�Xϻ0^��vъ�l�?L}w�Zj(b��ݷ��&=7�{
�\x_����Bհ�$"�%ϭ���ѳx�S��@|;Ÿ�����k�{~w�4����؏3\�����6���X[V�Sd��ޫÎ�,�]V䵼��ܗ��|����dJ��EUm�GX��m��HU�6�F\zu�	�����_:��d	�Dх��W�`ב�|��-hf����s�7�~�c��&�gm��X|��T�7b�څ������%"��/ia��B��K)&�g#��Jx����ŕo���Bt!�3�N캇fdZ��[���v,+���!W�E�����YT� �l�,�F�:ma���_�� 5�wvW�����Ƶ�wƊ跥!��~�+��SL�0-��o�*c)#&X#"׏C��j�-��>tE���iC���sJ$Bl��f�zW�ĥ��̄kA�������ؚ<��=�����b��#���y��#�=F��H�X���B&fSa4�n��o�u�i�ig���m�J�g� UҔ��Q�tf9��v�k��O<?mv9�_�4И��E��ϽJ<��s5�֌��'S]M�U���k���g�R��R��a+J넾�{K����~%?��W���I�w(�J�FdɵU�)�%�i�rۣ'b(�t���]��Un�c��{> 4��ׁ�uL�S�I�:�g�76����Y�_��V����wm������V���xK
�Ie�r)e\�;ȵ���2�i�yr��c�(�[$>�zp�L�;���Y�������(��鹇hkoy���'��6�ҥ2ǶvK7V�����Ĺ0z��+�x�hn;/�ׂ�Qݏ:��8[Ӥveٱ2)�\��p�
��ň�u�����F�L�ڪ����A��u5���w0�a{,�3��
��B&���T0�D3�Hz�|���Z}�IY-����?�9��b��T��~Ơ��ߛM]5�7�'��e�]�Z�i`�5�^5�>��{Q.$ߍ�)�gy�l&ͭgba�F��Zi��.lE�I�.fbނ|ڭ��cZWA>oD��]we�Z+�Y�Y�ޖO�{-��o�x�ժ�ܭ�=�P����8��-i�˲(�zZ@<�Q��
�ŝk�a�׌)�+�N���S����0Nk��v��Z9�uN�Sc��bDm���R�2hw_qt�{盾{J�8>����,��U���[�`�?�����ߗ�D�]��kX Ω�����c�lLE3�����N8��5#o�PB�]�B����#�����X*c�Vn��u��jq�ζ&��P/�U^c�0Q��;a���#�+�����o(��J^����2��� s�ά�n�2����H.���J�}�xġc�F�*`��f|��3���o��r�\4�ī�2h��i�E�J�V�����o�Ud�1�K#	$Ptqc���H��y�6j8��嫦S��_�����`��LK�-HNC���T�'�A|R��~�l|[��T$V,O��,,�J�l �Q ߅W8��֫*������Ta)�kh�h>���55{I�zt��t������ƺ:����Z�1����eXG�Q{rU�����������UޥT�EI�M8��u�sx�㠰w��[:�-^�Mb�2ji�K�2",�,��{��x)�~�/o"��?�|b�32�'��יf�n�!�յ�q�:r�]^-T�p&�7�oA�-[/oV�g��}��P����r��)Jzq� �D;'���e����_|��!K0Wgc�8D���]�K}oJ�f����\�{����-��Ō�M�Db��C�κm��*{0=�}�Ca� 컣�&mh��1��Z��ֻ��\6k7N�f'7)*m]N_P]�;����D�A��ls.�j�ӕ{���޲�j=�(���ld�͕��_�4�b����ZU�@�Z��CP��:�`a�l�GW˅�X�xX/�ipel���B�ܑW�YA�rⓉI������ɀQfb���j������2N�*鬼��r�3Kҍ�w,ʻ�	�.�+�T�kq�l�v)��i�ER��%�5�V x�Fh���3]XE-��p��A�f�D;�P� n���|��:V
=�v��V�3��W�Y�"G�����χ+�7�K#��@ލ�Qk!؝�"K�������d�j�x�G��y���!�|;?��[P�rݡ�w�]?_�Wptb	�w;2F�ϝ�����v�����:��!Ӓ�� �Z�O�K�&��R&���]��s-��T�����_�vN&���W�������(��~YJc%��$�ea6�����I^8o�Le�h�֬:��&4%��f�dC�Z��o�X��ܣ4Z)�7*�}YP�[��Y�2�7��;��6ɭ"KG\���� �m3�.[��):�M.���C8.�]���u�6�W�[�[�����=I��8��Fb��R���gw]^�\5t�ےI��H��H�=w��-���緖M1ۼ��n:�v�y0�n��ē"�#�ñ���r��(۳MU�Z��䩙HԬ�ʌ.�F�Ӳn>�^]%���������]�D�S���bnp,=�q��W����j�ނ���Z��{���A�M��l ���.k����JX�U�^k�����P3aA�3���S{�؀��dYV��-CI�һ*�-�"ӻ��9�G����ۧ}�*㙜-!��5:R����߅�g��,�M2�]��`�t���HD�7ъޝa��.��+&T]�H�ʏ���}�2�Kwr�X�5܏$�{vN�V FnyE/�Ao,��`�C�@NpEn^���"�f�����7?5GI�|�%ݖ�ۗ�ҹ�e�������Gd+����[�\���������J�靎2�E\��Uw{"��5���}���>�Q�F>��'�UL�ga���\I3K�T�T�)�;���>d8�����3�jS��;v��b��UfP��o����D������*d�ܯ-�2fbtV�Z�(��D�7�C��t�m�����m�Cs����WYV�Y�:�E��,:�6JH�hY>�g����f�J�A??�F��R<�#3\���J[ƈ>�Z�25g�44]HM�* a�������֫l�BKEP�%qo�˭����.�s��L�<��G��Q�-.�╽���s�t�xzr�s�ꂧ=�aG�Ñ<j+;#Xl��ď!��CՇ]M��r���j��7y9����H5���R�T�Ӻ����䲟 �� l�Je��8x����Ã�~��t
�E��*�^[I�x�B5����u
oA�u}��ٳa�1m,�K��O��(��x%�ߣ�S�I;zm;:cU�	�v���kr풝6�	��f������� :¦^,�+y8Wv�b� )��6ٌ�έ�!��r�]11�`r�8K����ЕO�����u�1�!`N�Aᷲ��N�y���s��R�5u-`<Y�a�a]٭͖�la�l����=x�"q�}�ܻ��1�/'*1�����Y�S�����	f�o�I��&���Z_���y;6�>�O�Y�l1yl�B}O�a��[[c��:����L��'5XZ���iT�*dP���(!�O��H�3�I�ι�m�K�Fq�ES�?M�}f����V�uG���P�9T��������#���~�?�������栒����
�W�av~y�>=��&�����t&Mђ�!�VL��)G��ojd�0w�q��9����w?Xx�^#��5o�5�)�T�Caъ&�[�Ά�mw*NdOÝ\��Z�Q��PO�����i��`h�*'u��[���@@��wb�N^OJ�T&���	�	ѣv��C�Y�_r���ڎ57P�J��ꛔvqQU"���#�y-�:��S��,n��CW;����e�YC�v������S>k���(���U���ݽ�:o��ק���:��99�~8�T�+�V��q���Yj{���d/X��5;>�b_YP�<�۩���Dgi�k���d�;J��d0^�ܾ���ϵ�j�^�����J#CK������b�Rޫ�!����]JM��{{{1��/"�'n�$L�q�n�s��{�愸�R�����3�yŰ�][לK �J�|�g��h��	Ws�9p|2�c��Q�1��4dՖ�ѲQWV��h����i���lV>[&��"Vkl������Tr�ܝB�1ҷ�N�!�䊡�ړ��Xd8��&~��u3�;��+�QȪQ��IF7#���k�a�Ujǥ�N�)��_e��3$g�[㫑��R���Du����"ҐL�Q6�<���g�6�]�P�2@v�Ge�8������&�l�28��n�{�G�G͵[�x'��5����f�y_�yV�V^y�V��Uw�Ī�9��1�����X+��":����e�_�m��y�|��1_�_�R��SU�E�4��X[aҁ�C�Ҽ��[�5I��OFiे��v%Ȳ��.�R�)�{3>��V�y+�z8a���9��6 |r�W.�Vw�&����)��y=>c�a�X,o�/�k�+��ZZikb�Ţ�A��y22n~ɭj�7���dϑ9�^���O|�]��8|:��fߐѱW)?(��1����'ŕ����"|�J7X���{T若x5N&���܏�i0����(�5Y�]���ټ�L�i�2������%�;0.����Bd0L�K�?WU6�~B�9�b,���7����T2YRY��U��u�ލ6'�{m�<�-�x=�v{�x(}��id���R��m�*��T}��L�j�:�s$u�G�h���D$ئ�}��ϕ*b�/2���J�sk��;4�4���d>�{�h�_��u�.�Z�]���vTd�����KS����?�9V�;.�WNͲХE�$3���*��b*4U{�-�b����o�^�_�3wR���ǷJ� T�����䓺��k*ZWw����e�F�/ݸ3��P��a���qv%v�͓w{I>7�T��OC�eG�SR�8�U&��u�m�r+�����,V��W[FAZ�o�������GH���ᄁJ��}Z�4M�`�u*����|������n}��X������b�*��N� ���v�s�N�i��s�!cD5 �Bvx���>�x[���h�2e%��W:v��K��^����}v�7�*k��ݶ��b��_�������̝��&e��Ө3��D@{�T�y��s��9�ؿ~����~d��L�Wx)���NZ�yTɮ���{�`����Kc]O��"]��u �����]�����z[�0�$W�x�����2��D���:N��S�o"�������#]u`2��hC�m)&��d1J ��N:�pQUA�V�X�VeǷ��O�N,��Xr"܁!M���	 ?���C�P�Ϊ�<&�f˩:��B[#�U�w�o ���� �N�'�����<�FȮa䦻%Y}}�'�o&vb��s�6J��=��±Aދ�B���M����2S��j��@�s��b��s�;Z�h�.΃`�#��1����7[l(��:�,�[S����*��+t�{� �2TKM���c��|}�����<�=Ҿt�
�?���յ�u�r������X�>���ik1�ܜ�/^T[i_TJg%,���Q��C��엗��M�ڱJ��s��X��*��Ce�0����jK�/xp��y��˹ƭ;�y���.�ڦw���[�Z�:#�r �5�4�9��ZJuAQ��
cMވ���v�j�ؗ���+�qp;U��,�Gh���w!����<�D?	�Μs��AUls;!ԭ���<ɾ4�lV\۪j3�iJ������Ac�����ǵ��h�q�l�ϳ�\�
b��/�.�Ȥ$�P}]ŝ��h~�ɲ�yH�n��4.ݫt���=MP�K��$�vdͩRn����ʢeHB��7$/����%�D��3 ���1O�u��{1slJ#�r��-ܭ�|�6�,xz�ײ�ڦȞ:�[/[M���&�֞f.�a<��?��;2��Ɵ[����O�P�n��4�ek�6�ژ�%���B����!n,Z�,����-�^d�KFǭ��F��<0��73H���Lx!�ag�l#�p��^n�xK�'�c�4\���wR~�u��>|��P~��Fx���ƨ�>�;a�&x�/���o�����&l�k!vq��6S��`�fc�����ʟS�+��\L��\����� �Má���8��y��G��Ќ9J��[����� kfQ�|�\r�C5R6ګnѕ�<�������O�
�t���N�WS0�29�<�)��v�o;]��s�tV$�r8)�/D�l^��\�&�N�	�Һ�<��J1c��1ɚ�\�Xfʰ�l�Gv�jv;+]���j�G�!C��'F�{�N�
 �Z���C��	g-���j���g�Oʲ�w*�fl�I��c'.���\�MUw&��l[ϖ|�6VES2��O�s�Jiw�P�5]_�Xص�;4���"���6������ak��Jӎ���0�,,�G���t��?-%뇪�T�얔��^�a��c7,��������:[r��^���.�,�,���PQ�0�R��F������
���[MGb��������6�zy�86��v����"b15��n��npT�VM>�<}�׎{]˩ɺ?!IM?*��]t_/���W�n����m��<1b ��-�Q	y�>\�*ЯC���UK�uя�j{��8O��m�sYͽ����1ꥻկ�x�س�;�Q�uT�*���{K��7^"4��r��G����؎��y\ؠ��n�ˈ��n�i��'�i�Y,�7jE����꣯oc����}x3ݪ��l8�y��ɽ�-c��d����̊�b�����w���^�g�o�z���菖�t��]�9G2�U��5�\�Eҡu�;z8^-j���N4�:y�O�S'lق���Z{8�2���и@*�p���L|�T;Y9 1C��bۧ�+�r�+o���]Zl��fsPh�c(]/�U�:�bT°��X���ͭ�=MF�릫pػ��^����]b�Gd!a�c^>�UxnW�.��� ����e*+�����4��(;@6���Y'DQ�e��R��P
2��H�5��Y�N�jj8"�rl��i�1�e��3���a�-L/z�������j� ���ʼ)��"'
�-�1�a`�����[��>	��ɛv���p��b��g��B
ν墛w2r��k�Qٮ��l>Ĺ�Z���c�J�B��������k�����NX��5�+���J��M{��C���U4��V�ڶ��k�C�o�q�����7ut�9\f�M�b�1|��ܱ`3��+��������M���=���2��W�s�cF���8hwO�x�c*��4���@�z�n�;�CV}s��l�`���#����R=���c�ѳ���3YN�]�80zt��9��ğf��hV�7�&c��u~�/i���zE��V��}1E���0 �_]n��\�_���)�	���}ul���p{��(m*_�4<�O o�e?*i���v��4���b�ӾZ�Ҝ쿅b�/k�諗����?z���
?F��$�:7�ĎF
8��t��g�h�b�&���g��Ǐn�&g=I���q�� �����S�|��1Xe��*�!;h/Ħ���n�'MK��#t��.���k��ܘ�fv��.䳛Ʒ��d<���x�	�#E,�;�k����s��?ٲ�;x�TP^��:�.DwZ��y����;�6h�NSs��ۇ9�rla-�x��T�Wh�8;�E|WYWP%Y��i���5ھ<�c�D��B��|�w`�*])�}���F��7�`�+{��R[���a�۫����`�B�?��;ⴶ�W`�Z�ꩊ0-]ߛ���vA���Xr}DT�Bwá����Zεw����/��ۛ�]��\��w �)�8���<�<Yl�A7-4(��U;��ǚ]*����h�x>wU�0�QI��e&f�n�e�N-�~s;-�V:�Q$o�k�:��"�&����4��ϓ�y�p~3Ӛ�޾�S�(����-�H1�hwrX����<qySw�1	���\9V���St�FL��I=��}�:\��sP+�}���`�Mt�u��ہd��J��e��N �}�eݞS<�u�Ɗ�s<�|���en�XU���Ѭt�Р����l.,�w��?��@���˻�}iP��)Q���d�j�`��l>� 	J�Mw����
?w}��y�2v޲e��
�sS�0�N�N��dN�����낎^:V���-6���e��-lX��N�{o[/�XИa��(^a�&d���X�y?������y;�"�^fvj=��n�<b��4xf�w�v;P�]n��W�ݘ�E��U��;2[����̲�^�9�-o6
�j�`�9,Z���5��tqc�dfm�mdn @Y*Zjr�mA�ҫ�}�je������l����1�;��!k&�⻉�	w�|�6Sޗ��!+"p�s��;��MI1t���5E���
xx׼��,��֡?w>���N�s;t���ذ �S06�f��o���,�+V��M��C�c�%.��\������8�\tst�e�h�,Y�B�^�L??�G�WS�=&kV ��&��Ӳ��0�ʮ?�V�t���L𜢶6$XǱT-���� ډ���������ϕ=��ܺ7ex�Q�.bu[���WS���88D��<i��Hf�\4i6H������a��7�@��Pw�X�������CWlv�a�F&��-�l����x���L�ޛY�k1��!������3F�Ω1���Ã-��b����ξ���+VER̠QL8�j5]�/~�������N"���
�Sem>���7L�ۣ�d��jҚs8^*����aƆ'q��5�5y���qvW�%"������w���-�Xzf�;�b�ۚ:M~�υ�e}뛿���v��>U����n�X��Rrm�끠q���P��{�V\E.z��맾w���ah:��aM�WɈ���Qv�g�CǙ8�
f<��קi��B�Z����0�^T�&Ќ/�|�Q����}�i3��6b�L��rΘ8������9y֛�]�"ˠnF���T9V�\ț�VX�Nh�P!��e:�|*vnb�W��C�"��h���7��݊����N��S��{Y�kn�,��3 ���#��|���r(nLC���؋w�����웜���|�H�x1t�qlz�I&{c�,��-��Zm�q׶��a�Tɮ��[K��[��ﮰf���Cw�V"��MY� <�l��R�GZu��=)��\�b ���(7[�Ľד��}���YPr���?B�s�YG_������Ŏc9�P檺�-���k��{:m�'x��&
8��0Z!�T�=~�;��4�Ծ�'��;57qӨE�|w�6���z&�x�M�IGWxy�{�����즱,�35~��5\.�������Kg�8�ޖ)!+"&�zaw�R�y�k�A9���rآ���
8�>S����7��L��KmJ�T���5T��R�=r�-�bPm�xc6Cu!]S�*�ی���=6��[�'�*��t�E���}���vc��Zd[��d.Yq�Ŗ�M-M�.m�2^Jh��+*1>�p"�1�'4=�D�«��|�V � �'�����Ou�䴆���^��Q�;�+9]S�\h����8��A�gw~���dKk�Ȣ���!�"u:���G+g=���5/1��*��3��i�7���Rk�W8�9��H*�Jem#�(J]�h��K�k5;�n�aK�#�S�Y+����]M	]u��ۑ_S�r��!)@"fr�[:��f���5�zc���S[+��zC�i��c�զ�yfގ�X�����P9<�8wn��9�����nX��+K�ꋾ�B�f��od��D����}Hڇ�)�q�����VvZ�c]^�bG)��2u��)�V�3��q��s{�6_B�j��Y !���j0-�m�@�fr�c1�`0�d�2�o�<sRV��Зߙ ���V�ۥ)��bMc(9e�'��[7{.������ �Ý��T�B�������+��1��'0��Y���9<��Vzqf��{�6�5���m����NN�N��aB��rW<��7�C$�vS�$���hLB!P�3,BثWw4��������t�칄����v����]\��qPz�*j�X��Va;���F*<�Y�+5�r�v��Ȱi�_Uݱ}��Z��D�:��]�nv����AͼZN�����R����7´���ƁC�-�Wp��[��b��NӣTRu��S��K�z��EZ���5�-BN�F�>��Q w<5�$�J^1��n&�.���k�u�|S;;�J����]Gyʴۢ��§�P:���
;��>헓���[��0(�j���@d����k�n���yI7@�
C&=m}���d�,9�/E�y�YW�U,��B�u��v���)ie������FC��eL�`�MO�q-���2^��6P�.j�'O�ӛFS�v,�M�L�i���Y(�Vʭj&�[t����Ր���TX٪����*�Ky�{�e��6�8��);�i�BN0Ϋ��ۧ������*h���e���͝��A��Bѱ7G��D�h���m�Sz��%81 &9b��n���W�u9�ԧk|���`+w)�t�:y��V��н ��
����]����c�Q�n�Q�� ����[+��Q�~Κ8�����7/5W9\N@6��T����T�*~���z4�+��xq�mOu��)���
/D�w��+��d����Vpͣ�J� E��%�/���>]�M"VřbO�������s��6���+�ȎMv?�H���=�}�2�/^�t�MJ��������fb#�����5/y_D�ִ��(��)R$��kH�ދ�ł�M�E�2� ,bo!������Y����X&�H��t4,C���p�bv
���d�?x�����k"iH��`��7]T�����."���:�2?	�I>w�t��\&iT�n[�V2):�n���fP﵅��)&�PN'4�}�)��֊J��%�jG�w�����+榛-�V%�U!Sjؽ�]���,S�z`O�77�O<$�<CD�\˦lYq��fD�[ŏ�+���U8���Q�Cz+O��%��HEg���פ�DBx�w��`A��@�r-�4L�dÞ�٭S1f�^��	m`ڇSu�[t�y �� �(�9�W���:�S.{�4�Ɓ�"pkCeױO%�k�ʭc����8�Nh���*_��P]lU1��y�:�-e��~���&�ƽ�N꯳D7�s�����OD:���4ɫk��u2U��\N��M��~�#,�F:bՊNJכNv�i3;�^�j�5$%�EI P4�<Q�a�~N`D�j��fcp���N3
R'W�&��5E.���X%֢+(`M+V�n'Φ{V��̈��i)\�r���D�μ�a����5�%UE�Oov�L>k�+r�_"��q�C��ƳQ:�"lO3EA؋�!������5E�"J�����QX*�p�M�#v��B�!��G�z�[�lwm[�mj|'�?�b6��$y������"�����a��!�\�V�9S��VŻ��&��|�n����d��]S�uG0�W��\UN���7�v�T�C�u��߻ھ���9�w�����f���u����TP%o-]Z r���}���,6�j��2*�缮^<����ĸ�$du�iv������V�7�ܸg�̕��"��G
l����5�I���.�Wz��Ʈj؊�9w��t�0R�A=mP\�sB�h�l�׭��AG�td�e�Ck/�Ï$�Ϛ�k��-w�[�hdl��K�r�|W+\��4��D�������c�ݲ"�"Q��<Y�&b��^��ΛS��0��ֶz9߻^����8vk9f��kS;2�h�FPb�TV�f]AB������FU��O���>�R|�\��6O�oX�$v�+�
�$��������-�^��O������B�'��v��w�r��a��l���eЮ�"6�hNQ�[��˷�2��F�L,[QՕQ��b����_vh����wٰP��a<髏�Lj�����Gl�f�9G��ɷOR��w���q��������u�ْ�-i�hFz�Y`�K̕;���nW
�CJ�R1��x�v��� x�}�ٸum�qᓱC�<m�����6nGj��j�Yx>��Y�(���l�xe�5< �O�������I�U�a�5/����_U��>������>�V�N~ֻQ�MD�ُIѲ�d�M��9�9Q�#��z�^��Vj�5d��Ϯ�|z1�ٴ�T{N�����ws=M��)� �c����*��Ģ�\Y�y�\ҳ��4��F���흑��_��mا�TpD	��c�;=_�ÏwmN�&ya�w���&�m��f?G��S����Y��F�=�SD���l
(�M��W�1�,�^���-%������5�Û���d���s���nctK���0�=����%���U����7Ȝ�޽���"g�R���N]��1�Ȋ*:��N��S m��?�? ��[���s��W��ԕ�z��ڧr���t5{8<�qg ֵ�#  є�}Q�&���c�#Ȣ�g��[���M��ɘ�����YL֎�bck���(�ں�Z���ƽ5��^�ei/��7��Dhɤ#���)��l_Ú��or��}��7O��yv�9�M|�E3�b�]b�\�f-�}<�A����ːe�T�ݐ���Q�IN���B͜��@޲u*�-R@_ٹӧܯ���5������P��ثz�ʄw�n+���M��0��\t���gm��޾hH�ʤ���JV=�����uD��P�[z�J����U[٪~��ݪ���d ���'ƊA퟈wc��v8����+��Z!�҅ohQ2oc��'笨�F�;V�<�Vo-9nz���O<g��]��fv���[���!�����,�2�Fw(K���E�|��ڕ�`V�zLsÝE�;�s�Iվ�(�W��R�;elK�n�|>�)��d܈-��e	����n���Xl�4<V��=̿۟���Q�k�D�Tq%�����J�
-ri�.������gt���b���7m��FL�Vū�Z�P!�>t*�jpضG,�utĵ6���4�`��e4.z!�{m��Om�6۽(����-Te�k�"w�N�/EB�sͣ�p���Uۯ��7�ή��(󪹣ق}:-(�i[%��V�����uD0�j�Г�{"K/w�ޝ9�r�ܾ��M�3�!�V���~�ߐ2�ex�YS��7�=��n��8��n=]USԘ��Ґ�q��QY��W(޴��(��+�l���1��_�LК��2�a��u�����ƻ�n�SK�XEu�}u	��j+��Sw-�g��_}�_�nQ��Yj�}����*��T+,D�JU��ꄤ\�`�����;	v`&�UË�z��$���=E�bH�Ł�����������u��ˉ<9���U�|�l�`�z�w��Rv�`��a潩���]�]��O�M6l�r�V����B�����u��򋽔�p���R�.�.~���zr��������ۧyT�D��u�c�����7w�]I��z�����~��,@V�]���;8��Ҡɣ�:��Kȭ�~ǀ��	iܛ�#*�fUeNZ���Օ�{�y�v���3��<m���u����~񼱴�,<������U�o�מ��1P�=���k��=1��5$��[�ޓ+�����\Ǘcm#<�}��]�^澇0��)j���z�n�5`>KIǧ��F�M����
�$񉗂%=��QR1O?�v�>�`�x���R��7I�u�*Z���TVn.V��;{o<6�Fdsbz��j۠wU��+����/�Q�V�@7wfǊ�$8�.6�I���*�;X�V���n���Wm���޲kku{`�`C^+��i��S�#n�`��0�+,Q�\�C���d*d);$I��;�R�1T��^��Av����	vhZcp�	
�0x~�V�!��mY�������6�w9���g�� b&L�"뇶��%����)>�A����4<��:"��".=b^���(��u�;7�>��]`�����U����7��%*fh���s.�-`)��2�y�z�\y����f���t�HP%@,�,7e	���Ɖ��A�^��v�-n.�oۓ�ԣAbU�2�7�	 ���$D��ź���`�Z1����[|q_&���������OSad�$�R�)����ҪDm�L�L"T�,��!eS`�nY�(b0�`ru�|�y~~~�^���j������ǖ��-c`��BN?�&4BM�Jt��k��e�٤_l���e�K�Zν�;͖�X�񫷫'�u9�4U#Uf�&z�O���\���4Ta���5L�H9$-�G(6u��W��3%1�����c֪��켥KF�cJ��K*�{&���h��Qv�Y�x���;^%���P�����as�\��x�n�t��Hw�������uw���1
c�3D|�M?c�#�IK�Sӳ2��ХI2��ܓ�ͤ떽��^B���"ĩ�֨���0��7x�ͺ7뮞~\|V�%/�~�_�Vz�J�\4�Ԭ_gi��)J��˱�۝
�H������<�<9囜yG�˯�kr�S~#���Mo�t�#���q�9 SeƖ=VZ��윝Tf�ӽ�;���7T7�g<��(y��y� E�&����w�:[�]�˃���T��DU��~���ЏX��L��@��M#5JP�<a-�A_8�\-�m%��.���r~P��܋\��;�s,tQ|}�ڬT�e_Wv;�tn��q�W��>������=�?�bԮ�ka��Z+�B�F�2��[T����ii�֊8�[9Μ�9}{��Hok��5���|8LG�JБ�7���=r����i�U��}|�ެ�grn�'����r$�X����b�Q���a�9E�i;��:�m� ��TiOes��r�;�+����YfףS h����g�s_Hz��mG3<�/ݝ�'�B�V��p������뼥�~�"����w�Y0�k��H��W�����r�6qn)��9KHt�п	*�T������3���FWxa�Sf�a�N���y��W=�]��Z܂�֦*'����j���=��vpi�;��J_*��;�O���`n�Q}���5<cyѐ���ٔ���"��rj$��K��0jxή��y�X�	�^9u5y����{�p�������ۧGj��^c˞S��H�_��/6s�>�S\9M���U�焖��Ю9���m�愭����!'r@Im&�oŌ��fQ��fW�z�y��<�����~�Ǉ��T΄1���X���c�i��ov:���Sإ���VO�,A.{N{s�kq����ە�q�^��j+a�ɪś\�3W(��m�|��q�.��|�6��e�Ks�!F.Mj�;�G�4�]�������tŕ�,$˂X�iZ����9�����/� F�]WO�'2ƫ�\a�"��;�����!F�.�Z��Q�g}��e0IE�?�@�օ[�~�uu�;�	L���ߚ7��ׯ�޼?�D���۝s ��]���ceZ ��<��{z�Y�R��<d���G»��y
����{�U��j��#&���|r��|���gG>� Б��&7_�#�Rc�W��Qͨu���`i���-d냯�dJ��Qx�d^Bv;��q��r/��e�SC�y����L��U͏`�g���0ꄴ2��']�1��ez�,fu+�,�\����L�כ�7��k���n��|��F1�c���s��=q�X�GJ�0�7W�S�4��>���P>�yw}p�.�-q8�#���K7�I��2 �u�7��~+W����𪞵�᛭�/�����^ɾ��(�z�c�������A@�9�ٵ�l��j�%~Ñ�#�:.L�e�9����p�9zл3���'ܷ��Oyy/�(|W��#�D�{E�㇮���2�t��X��^x�s-?���������ku� ��C�����R��5'��ȸ��]�L��*0�w,��!1J��������$�3�Uw��z�����p��L���z���O
� ��ޞ�s���\v����m���=S׎s�/����Fn�JR�q��3��L������>�s����/-$��%�\p#�s���u���˚/ie�#�zs�7�|P˘��䲚p,��x�a^M�F�Ƿ"�r�8�k����@��hډ�����nz؏�wV���94��.��3kwu�LJ�Vb��;����MQ���%O�G�e�O��.��GX-G�����"#��ht@MzE�M^�[kw�VD7OY.��ġ���� 0'gw��d��=�`���HZ�\ի3�'w��,+Lt��&X�Մ�A��jv��DJ����W؛��5Z��sz���Ct�����xw�|����1_՞�q��Apι�������y���g{�������EÁ*��u_j6�󌛪��}��"`oW��>x���1M�~
,G���u�����;���{j�*�N�j�H��M�k�b	�49�b�/J�Չ�W��:_��>���f��t�����7�z��E�"���/qҨ>Wk-/;��k��En���V�}���"X���M��霻�N��ا�_�����U���:-5%���ȅ+���Ǉ���I�*fHU��Lbo�����O�Z�f�E��ٴ�q��g��G�����<I��Qd�n9|6�MM!<�g3qft��)n=c2+�v}4DoN���_y�*��s��Ir�8�ɩC��1� �ᆝ��,86�f���hG]]c:�=��Eck��Εw�]�W<�\G(wY�%�2� �mn�Qw'����S�r�>N����ΆYd(�膫 �L��E7D�:Wf*����L����7�b�,dbg�e��(;C���Q|WF�LM��c�lv8��C�+Y��2k,jz7R�s�	k��׶&ۂL����m�QJ�(㟾�i>�Q-kի�VՓ�6 ���1���]���U�ߖ��T��G]R��TZ�T�! �z��r��w�.��+1h�z�:�8��R���Syy��|��U�oM" S��T�	S��٫{�{��v���qfWS��Т�ˍ�c���� �+)�gT!5���]�pA�\4�Qm�wn5W�����Y&������ش�\�SkM7]d��(�p����c��xh&ݒ�:^�ϩ�|�O�}L��Z��L���x��\:�����vν�TI�cZ9��{Kvw����,x�����jQi��:��CS:���C�]H�tAX��d�u��lfq�	'ߪ
&�+}s�c"��gt5*��0��kؑ1H>��-�mQ	{3j�q���ָݚsn��w8�:����s%���;���j�`=ʊ�nf4�3r~w��1�QQ롺���İn�pdc�s{�A�	2;G���m��4y����<��R��{#v+<�����I����� ,
N����*J8\���ǳ�ӻTH���]��T���wlN۸�����
Mo
����y��k�|��w�e��e9��k�������<��2��{�Vnf��|g��Z���YiZ��w�Ю����aŷqН}Cm��C�8�bӗ���O��*�h�y,`�]�m0�N�+��{���%3I�K^�@�Q���cV�s2��.�SKjc��&_0��4�^aǏ������gss7B��~�`�%ŭ�zj�#ew%���w!�6'�5��~���H�:o\�P�q+�'?�R&�����V:g�.Ŷ>�g��0���;�����~R�ܽ��4�F'��M�9.L����u^/ϙv�J�pLuț�WV.{a�v�����j77v�b%�D�T�l��7��I�rh�י�Z��)�{��{Z����������-y1�_Wv�����I���Z��yª�d�sY�0z�#Im/]��}�ډOM(�t�3��s2�l������v�T4=�{��[��@��y&I�K�Ǽ\��?��>�\��7��rP�wK@�� $�	ʩ�׬QJ)7mV���]w~_�"��Z��h�Ղ^j���hL�-��WVo�
X��,5%*���d<B��r��A
�s'&tC�4�U����>A(�Rc�n+On�Ｙ�������,v�l���$����
��Ӽc5靡݋p�x��y����vF������p����c7�d=��}���,��shm�z���o{�jֆ��(%�]doPZi'(�-��R�j
��{�Pd���,CYS��p�n��@=��Q��@~���Zʜ�Q�u�w��wom2o�+Θr�m-o1��)�����P�팆uZ�Y[�x��2l�\ʙ2Q�V�_n���}E�al��1^��4�Zk�˥}�w*gSO�����(�[��/�Jٙf3A%�I%֪M�Ƞ���7�p������N��"�i��:$o?.�gw5c�&��[]�i�����n�n����� %n�0[��Fo����k�MlY��6]�K��[|��kX�{9J}����{&��b������d	J ��4�[�$�f�xȓ �Y�*u �޺ˏC�F[�T�N:���u^[�YEtg+mK�X�v��]�M�$����Ij�F�&0jc��jp
g�Hw�F��ԩ�-pc%mh̾/9��|��Mw��Y��<y��Ur��7��ö�ūq�����WԆ��G9R�:��-��]z�k�Y��΋Xķ��ݐa=ɞ+�D�d��œV��O�1_�nѐ7(�w���0��%T�^ҷ&Ԥ����+_N�jE��X�X�N2�_!SK�D���"�v�u[�����e>�U����G���N�<4V�ͮ�\�Zͼ9r5��~�_v�;����=��Oe,(a�����>}��s9�K��)�iv!-$.��[ړ�e�avT�,�'$U��FxL�0����m���E;��ÕYtj�DԚ:��<�ҫ�z���}�*+�u}7��b��tkx��ib� �s�������+=\��ѽ$�̠��t��Y���T�[��Q;&���oR|̙7p40<�w+��U�ڸ��R�s�D�������8��]�:�|+M⻊IX ��EcO&ʧu5n+tM%+6�}�EX��!P~xCy�̭}u�+���,�C\.F�q1�b�s4A��~2���:�/n���Q�l M�R�e�̆!Y��XJS��_t�8���Ӕ0��R���Eub{Z�w�ܰi�����WRX�wg ���Ut73l1^�`�j�9����@e�>���뮛�A-��Xwh�ő�g&����CY]�vdW2��r�vqɼE��(ۋ''�:;'i	��4�7Q˻ͨ�_�2�KZH���mᲷ����2rT6�O%Y��3ۖ6�E����_,�⟳2�|��ZRx�a�b�y�Pj7��ƛ�^�}|-�c=T�{L��w�<ߴb ﲏ�9����s6i9sk5����-�MKޣ�E[�g�]B��Q�γw��6�z)���בd8�����������̋j�-wܗ\}��W���O�j��J�>/���y�x���<Z]�5yYcS�n����������������a�Z��f6|i����V&"^HVB�A���|�rN�5�=��nfNJ��T�sY�L�dcgCݵ�DM���wrn�ue[Z �:&z?+��}�t3��3&�»�u���Kӏ����6}��Eĳ=�ƨ�]5u,�����h�v����P��
�8_���w8�f��;�e"�͎hn��OW�U��Vr��.���j�n�3.�(F�
�=l� y$�Լ�^�k�Ovmqb��4L�E�\8ގ���P�Yk;�����X�T.W��:����e__���tz��kد;��L�����}ue@<���x�pỰ��,`�����4�4F3F��a�}��m�׃�u��N�u͉��p;��2�Ŝ�E��7�����-�9��m�~y���z�4@ʚ��[�;�kk��T"����2��>]=l�c���/�=�k�u�~>=@I����:�L{�#��۶�׫�SE��l��޵�Q�X���53D=�yO&�U\fRx%�ɠd�~�@ �h����Ґ�֤VV��w�r�Hs��8��W{�94��{��o9���/gZ�Ъ�c&�*B�}&W#+312K]d�oqx�t[+\��~�9���dC�2�r���x�e�*��_+_��zLaҘYѦ�߼��u�y6G,>����|!8&�7g��b�8���S��
�E�,�_vI5>����M�ZoN�,����lֱ٢���yd*����.�=�~��nV�j��z'yмk41R����LWoPx�G������WS{�U��Tފ�8�6�,`_��;��(&�"$�]��V�ݍ��ݳ]��§�ϰvX�s�E�{+21,QIZ�{���']����R1r�YJ9��q&���{�+�@PH��4~��}����`�����RJWK3>�zL��ݥ�zߖ!W�>�۰��%ĥ�{�,��La���Pref��3\YZ�w��Qeԝ��u�$Z�lCA��V1���:���j�яlp�����aG/�ҿMP�U� [k�L���M�M��T�:�'q;��qL&\X%&�-B�l�%}:�>���t�&�i{"�.��N�UڢD�,�߉�
��y6Ę���Z6��Q��d��[|��_E2��N��?w�p���4�Mo&)q�A�*J���I�3M�6����,���}{5�ö�(�i�)$��,N��$�ޝ�L�;^s��v��8&édbH2�i��<��Ղ�����,z�um�>k!Q�W9ّ�5Xr�r��7ԭ�qۅ�uβ/�0 .X=�D��_>�vF��0���z�>��l��SSbl���膧�d�<�gA��jom/K��Οs�'ԑ���W�2ӛ',6Z}@D1b]�m�{`��λ*Rf�0�)��ڞ��Q��3\�9%3�P����f�W��Jvzz/o̩6fc�Yf��j��V@+�FF�㵬�� �]��c���l%����rs^��ſ�<j��
J�}�c�}�xWrΆΌ��iU�w��=g�W�M���L6L�*1cT��$4h3e6�é��1��+��n^ӱ�M�6"�7*����
��W�˹���Qu%{cװ���;�F���=!�@�ˆ��#�-B���2EM2d1���Q�*�ؚuIzo~��A�H�q�u�Ԃ|y2����ǉ|y���t����ݼ}8�R�l��Lx�G�lu�X�Ɖh�&	OR��{��^L���[��y�=���u���w�V����ff�W��g�o7`·u�</p':b8P��N��ά�v�p��s	b���E��q�,��:�}��.��+��¸qѹw�R�����;����RZ�����"I)^Q}d�QrX	��Z�Ψ���zcv�흽�^;)������y�be�,pHڋ��Ȧ��kH2$�c&t{].��5�E�9�M������5�d�=1v���B4�&:Y�e+�b��>�p��D��z&�!Ky�v�HsL&�큻�wa[O�����ۏ����,���~6ZT����h��'�RF����JݡI���_w)ڻ� �����nQF��/��i����=�V��[�y�!O����m_�y�qRFO7��u(Q�ޒ�;���fxG��EGf�1+}����e"���FQ?�R��CI��C._�w276�p���/ml����/,������t_wݎ�Up�Ӌ&\H4o���*yԆ����X[�����i^��f�zՍ���Z�ɉd��^���������6�����{��8��|
?v�4W��OJ�����UH��C��e��aۙ��;J��5f-�X��+++�Q���*��w�Hm����������~R]�GؗU��:7_c�s��/�e�#T99��bB�<�D�9���,�њ��KK �w����#V�ՁM]N�xQ5�(N�2�'��V4�m�>xS��m�y6���J�V;�̽�H��D]55�'����2���z#n$��eEV��dRyt/^�ȴw�iX:��ҫ�<ͮ�q�y�[Ӻ��m^�DY^^���	��G9'�O6'w������v-�i��1�I���߾��4���Y[�[wT�X�/�j�_oq�"J�컃�t�q��q��W�Sc\I�e:-�r	4Y�Cl�R7v����X��uF���'f}C^^:&C�0>�$Dj�E I��Q�ᄔ"E������𰈂��Y��X��\��&b�]S������0��\��m�Ox���j}��8(��Q��_ܵ}g�d	�f��)��{|�ξ�ep�fZ$N��q�-7e_W��{]'�P������;�3wL�q��NLvB���D�N�$f,fW3�X��6�v�UHx��i5����JT�v�6�ew"D�/���g#m8����P�W<���y)
�&���ˌ�&���/�4��ͷ��D�m�=�=c�p̓���N�|d�4F�3�K���7�2���=�b}������?�w���-t��9®sQB���y��������ؽ#{�������p3�Ớz�s��V�58�YI,�+(�M�Q`���L���Q�Z�y�ܲ��+/��v�U���u�}���励6�[��6�Ue�6�Vn!P��fPo5�S�������*�
�Q����c�侬���X&��'cZ���g���j����|�vL��I�D�׋sz(�GK��~7;//
����P��x��K��K����[��������]�N2�{Y�X��j��KYJ*�TY	UG�'�~�%3�U����a7e-���\Uϧqm|N�*1d��9�wH�T�R���v��o/=J�c�\(� ��{�]�ˆ�jI�V��b�"_���s���iv���I9��uu�͋�y���Т�ΨZح4/d��t���tM�E*}�7Uu�5�#�b��
̷CoIO'��i�i��AkL���V&(��i;ϘϾ?�����P�se�&��d'X�Z�^����Ok��ʜ���,p��7�ު�ܯo{�Dn]��|��
�;}���fm����e���u�c�eO+G؅�n�ml�F��y$(Q��ێBٝ�������[��+����0��D��p��FǴn���7�F����+�������HS��:��]]��D��%8��~��F��`wާ����躋>{,�(����Bs���v�-�ۂ'h�K��{���k����9���+C��	y��x�X͝�����J>��f@Ƿ܈�3�P{�݅7����jTƅ�]GK:}Ë}�]��j��'��P��mֻ��cf�o4�p�L�wa��.��E��1��c�u��0�-	�Eu�zhi�@Te'E!�#e	")
Uŕꀪ�M�
��Am���r����S%���u�,ݚ&:�(28����O�M�Iְn�U~p2�ETn�4IE��c����}>���/�v�T��������/t*�ҭ��A��GI��	=�����k�(f�� e��k�~�9����cC��o�*yn�(\��ᕝ�����M���sJ�>T��ѻm�aZYm���g�u�*�Q�4�=�U�82���n�ҫ/�׵�c|3kV!�^���W|�ҿ�>�_kCk����QYj���5����t�?ob1i/��N�]�C����1�~�������졨వ����Q���Ӫ��aG�p*��/y{^�~�l�k�*������ڙ��>���]��z���O�*C�/'�8�RxQ�E{!vG�6W�\X�S�j��ܨ���:�z�� d-��}�U1�óF�Ɇ��jgo*�0�O�����\����
�c��'�n(�Q�#n�e��4����<Q��ME�����g��r�xh#kn{Jc!U���6lʊ��`����L���Ki/f�����xo1��y8�n�l��:��Ab^,H�T�;�Hb}�go��b틤OVu��-�oL������ܣ�H|e��l,y���ONޣ1"m�uE\�5��v��;�%g\��C֊�)ĉ˧ˬO�b�w;Hn��Yi���'��j��ܨ�F2�v]�Xs�~��*�������g5)�iy^������Q�ETK(�soL������Y�����zD6�#EdD�M�i��gI�\Ƈ���x��%��׳2�+�(�E��s�G�|v���к.�α�T<��`B���m�-yibLk����dE�s�������d�F�sK�Hc"G�LnaERE�4Z���j�z"�{q]��EϺ�y�6�S�'��T\%&��� �>Qܦ�<��4g���-8j�ö�aY�bz3�Li�t���ֲ5qy�Cb�Ⱦ<����Ӳ�e�ga�	���ߨ�;"<�e]�_%�&��"v� '��?��b���<�"���.���^��j�"s�܍�p��C��9����I]��"�R1��@oMiJC`PZ����}훊k��LT �m��)�,|ݼ9/m͊Nn�B��&}����f��I�?�҅��R$^TM��w��nm��Ї��W���޿���n�ܭ�T��%��_���M�}�-j��zT��0+����ɕ��;���9="���^���s�k@�f�9U����fn1��*�<�I��ǂ�ABؽ��]]�du������ږ�T݇0T�Ǜۺ���D���J �ǚswo:�,q�;����v��s�5;����J�iFd���������A��r��>W��Z.x�-JO=s�L���3~~[�U9�mщ}��4��l�T�#�+��Te\1Ք2������fiE����=?W��	�І8�jy�R'{��������D�=�}�<��s�z����ΐ]��.�L���u���ꮒ�� y�+��*�����zb�������wIc?P�\I4h��!
 B
�9&����}��ʳ!���Gb<a��V(~=�K�����\mp
54wݙ�o�k��o�+�~��[4Ov֭�x�f��6A��#Q!��Y1`�wLN�9�.Ǖ��?�8���9x��}�?W�HhG�p�0N�]�잣>X͔��q�<�������1������D���Sv�v�w�:�,`����k���)������������Ks 2�[�]�r��=Wr�E�2����nK��ۻ��trޒ�H�)P�Y��Oו�����-�O˥SM�k��mnt��i�Z�Ve�xS��cvަ���x����,����^׭��*���qХW�1�t覾5�����e%Z�|{�����)�_fH�m�:��e~Y��\�"��ب{I��%r���#�s��Ꮶ��g���:�ܥ9�.꒼ͷ����@ө9,6|ɍ4<���!�ޱ��?��xV�+~��N���qڝiɬ��\3�KS�U�s�	O���`����w�=�����)�}�?bh��
�ǟ�;2�2IZ��ZGFOȩ�J쑡�s����w��\%��{6�v����[���ǈ�Κ{F�,�/q�_���g�WI�O}N��^y5��z�K�K�Y?\��G�)�}�����5q��9KF��ז���9y�`wBa2��E�Y픥�wGF�wPYw]�#��
&��O��Aǌ��b2�wKH�J勇bL�w�����zh\#���ʫ_[rbI'����V���1�U��b��f�:�gM�L�NN6=�Q Q���a��S�7K�!��QH�D^����=���e8V	���gG���o2�yX��|@>1}�y�{�Ӏ@\{���3��WvcF�nN���z�u�ck�ۚ7lD��F^��1=j��l�_1��M�\������fKX��or3��>^æ3�C���\̹v�S��y��]�uL������H4��S�B;��M$t��|L\B�����;���V麸��<����й��}�D�F���	9z���D�C4����B��s�'(Հ8<�[����u�]�f!��Y����"�AWُ7�j�U�ݓ�WR��p��m� ��9+�R�Y���vkb�D����X���9�֚�q�0���v���M�#�����`��9��_��\�5ƱX˙2h� �s? Q�J�ę�*��LX�����de�c0;e ]ʸ9��]��L����[�6'[,�sr�LU�F��"��g�l/*�3Ʋ��峒����=�:"Y�������s/hv�(�]��#��4?J]\��#�Mm�=���R\�b��M�wϷ�z+�͆�PP��/��et$>���
��N�3c�O�UM���.���Mr|d%�oIe���wq�mm$0�]���3n��������x�*��͎ax�FP;u� ƒ���
��ju�]�n��.��n>ˡƖb����V#��i�a_pyZ�=���e�ͪ����#]���aA�[�x
�!�?Cv�@Ģj��JGu �Gw"o���e=��V���)��L�=;W=w�{��i��p��������9���fa�,U�i��;Mm�<{1l�;�B���\uCF̮��R'u��vm�աkZ����L����t��Xzu���1]o.l�u���I��AG�Ǐ�yz���7[؂�%�X�����,��j���966�H�Fس���mIX��$�K$��S*pu�d(JӖ�m��X[mtR�܅��V�,C���sb�"᪊TϤN-�rңE(~�ɿJ�#��B��J�g�H��ynTj*��g�)4.ǔ%@M-$l���J����X5G{M�BPZb��cs ��i���ث��S5caYRT��}�;u���JYׂ�3J�]����r]��YD�?�V5�5e~ ߍ���)�[��x�w.����Dl��^�-�{ZGX�rܥ�ו,0��p6�b�����+��1�b�d4j�����'�[�7�R鏟h�+�pt'6�CZ�����'����9�#	�2��_fb.�6h]w3+I+v�Xk�}ch�]��g��I�:����]M$'4T�S; e	ԑ�[Y��]�n���5=g�l�n<��N�?���Tj#�4�w�¥k]M��A�i& ��41�;)22i��;暎%*A���zx�M
62��$�K7�".��VYA9%��O�Eh�e�yl>b���&x���^J��B���QU�^ܚ��K�3���q[$�G/�����~j��窂r
KPC>��x��F��@<���s\�O����D��S����*���ǉં�G>�2��;ۤo��M��}DR�*�_���%�3�D~�1��{�_�5N��އ�m���y�E�7��Ζ�I-���_�9�$�>�������T�'L���Ƃ�U�ٷ�E1��[����-���nc�i�T��a�q�íX Ì���%{UO[!p��-�������P�����I9�왥��I"�K��}8H���Hb��9�{n<F�kڦ�]4P�i;�h�u�G���
/?ܳ�?�W�رB�)��0���	�پ��G0s���-s��^�/ufb�.�[,"2���X�]`8]���-�Ԇ��� C�M|����DK��k�c���}۞�:��M�Ce�Pc%����AZ�v+�a��� �{\޺��g�{�]d�Rp��ؐ�`��X��VX*�tA�čօY��5����.�j�ɿ�
��q�_9����p�=�-�e?V��n�)���Oev��)���D�b~���Ȅu�ϻ7%��%܈�*��L���A����Ka�qĊk�����v�xŎ�����w��z��RsL�j݂:����։~N�[Z�
��|�1���k��z��.�5�	�I���5v ��2�`���[��x6r��aH�ԪE�q�g6�'�!���w=����gQ��&�؉��wJ��ɖ<��3�����I�iJ����TH�s�M���'F�o%�Ż&w�צ���?hn���>�����Y1q�;�_P&v���zt�(V�<����_x���������v>{$:��E��
���wi_;;t6U���k����`�{�p���}�/؏������[a[��FmO]u>���C�s7J�bM ��+<|�5��n�`��oَ��Q��Y�5c�C��ak��j
TΪ���i����`:l��\��{+��󡧽�
��ƒm�QbU4���V�)+�G
Q���a��Nح#n�D��s�l���"�%�}㽑���d��^���ڇh��󮓹���]q_ u罇�>��|���=�M4��o����gqW����/��Q�t�mJ��
��.�%]h	����9e^eoG�/�(O]0F����n��ZU���V�4�1��p���`�,l�٤I��\����M���M�I]���\�*f�6��o0�E�'M�$r�bhًbCFD��a�����y���/wfT���e��^{�8)μn������V���C&�Z3��eK9���R3'�;q3ݲ2z�����",LybZ*�t��s#k^�>ga�Ow�Wo���VZ�ܺ���{f��^�hϽ
z���q��>�t�C�	N�3��(A��#��J��J���e��e<1����J��2Ռ9:�H��MG^5n�ԋ=uD��2�z�� w*&f���_k��!�]i=�an�(eǲ���ݜ��ܣ��N��YQ���,�/u���V..	��3g��&l�H���ˮm]QZ#N���R�a�_m΢@�Sa��~���?�+��V�x
y����n��h;s�7X݋�l,}~�Y�.�n�`�ҝ
~`$E�ɑ�V�!\��ixar��h(ॊ�6j��דUp3�k�j�;S���}�%��4�<G�篳JU�������^�<:<��֟���`�ff�]mn���
z:["D���}ѽ�WW�ݵ�4�T�gYv��ߡYk�u�%��\k�W.[�~�
��Q�8��D�s�~�]|X�(�������S�!Pz�����J7@
&Y�A�ٳ8]IJ�.'�#V8�>������oV>�)�X�	¦��z�>���~9�~ېV|����[��s�j_y	��{xh��+Y�m\�oV�$p2�������Mn��+3]x�Ņ�/*��wHoj�xz�ϲ#c��φ�^��l8�v�z�Z�*�����E�;,�<����΁��hKw��6VzØ~�׋Y>���l���(����U�fk��eM�[��bg.�;����Ö��$4J1��T�*�Q�����F��$��n�)c��z�O;���l��yZ-�.�l�< ����=�^�_��_���"Є.K�U�Mz��&�6��W��k�uQ�+S�x�4�}����I�}J!����v�� �<nM�w�� 2��폤՗����݋Vs^*;Zu�vOX6A��l�S%��r��~��pk�|����b�i��U��ħ����mV��n0�ͦ�|��Ǧ���7.�q4-0y{�O��ʸN�-�/_�����}�u	����=ܮ���l�]�)=:�1�=����5H���:�ڣ2���e]���=B��� �E�_�������.�\.���239������W��Iv^+L��ph����3XJ�����;Gv������l�9��Gv����vd�ٮ���n���%�O9�G�\�#{��~�&GV�����X���ePPgwH=��@�''��Y>w����-A�L����y��Y�t#�ڍW;cc�l�l����Uڙ�S�(w�^�z�"�x�[����p���bK:H�3���ڶ&CHBR"�ъ�	���|(ݻW�׍����b�iFM)�w�.��ۚj31�(�2�N8��{�,_��<�C��F�&�8Q�Y�`�n�:ks�\�:����㌷���9γw{0P��|�Q��i��G��ؔYǸ}�f���ǥ���O��{��N>���T��1��Ǒc�9y�lswc#d�|��'��o�Ůƛ��:�od�W&*���Z E�t�ӕ��^�v�n#^ɢb*ڈ�>w��o4H�f�2o��μ�d�W؝�͜������R�n/C���u��Wy^�>N��g�$�}���r��I��%������ɩ�h�Kć1�︱�	3n���o Qt��4u�m��<:Iv{��7��k��7Ի1����~��� E/,=����=n��C<m�[��B�[�!|�*���X��ݦ3 ��%J�\+�L��:����`Da%S��n��t�]r��t���d��
�,s������\�n� �C��~&��1G-�:J�����7h�O�,D����E9s���x%Ѣe[��[W89=l����ח���.#xR�'8�Z��B)7`q�91Z�q���4�F�և!#���d���L(:M���mr�UƑ$����׻��/�B��vj*1QѢM�&��4HA��6A��نo�^�}�Ř�S�O��﫼�Y���)}���Z�Ԯ{�@�1����2*�W[�kJ�w�����N��g���S�^Fw;�ݱ��@�C=�s��>"'�[O~�	�)C��v�$g�#�lR3�S���8zٜ�{�N�۝��B�/u�U<����6y�s�������b��w��9�� 2��
I����'��W�]�c���`_T�E�Eڍ�"�t����}9��]���E�|�x�.I��X���5��T�����O����<	��z9�����	K����g��tW��wœq���.yǫV]��I�HǱx�~�TQ��#�M]V?=��-��T��h����F��rZw+�� I+S�ʃTj7���2|:n����S�y�}#)�c
��.�ͬS�![R7cc�� ���z&Z1:I���\�FtV��Yg��w��I�[�d�g=��`E]�j����9�g{k��8��)�%Yyu�������	p!�lZ��(G':�}c�{��@���r�:N�
�C���{�M�:n��ҝ�����ÊT�J�@:1���Pb����T��L��U<�8�H�%���yq5�b�p�= �
ae
���q����I[��a�p��Z溹�X���9��w<�)r�ͨ�����h\���]]l'R)M^���\M�W;��������+3�gtW��-�ս��z�	����k�VI����bxgb�%�^c]����g[,�nWCaآ����a�s]N���voѿC�_������Ý�؆7�Ni����U�nymݥ�OŶ�&��.��*�n�U�`ۃ/�e�!ɀI�T����
_��(�zU��׺|<���s��*�ek���ɳ!�|��Jnq^*�{�do�a�C%�u�{�k�A{�r���Jp�	�W
-��.Pz�	,���N��PfL�rVK�����v��Mq����L��_��8����ދX�e�O�72lu��t�ie�<[�t��x��c��M�YTvw��7S����,��f�9���{5�؟^o'J�� .�O�<弢�sf�;�tG9�P���ok�<v�5S]�Az
�}�دq߸�4r0�Ӵ>���qYF��g;c9ig�s^UM��mJ�"�Zg��܋��"�L�r��qs-�Bq0w,���˺ӭŜ0��rt�m��CE� �k��6�{X���5톰f,<�Z�y�gFj����лt }�G{�U�5ڲd��V~G��e_��w]^!���߸"�kw�����6u�x׆���ٛ�6�:���~�����+}��o�.etF�&�2c`����Ʌ$sQ�ݽ�[�ΐ����K����|���7/��j�o���)������]���������`�͂��}�a^y#Ȋ ��v/VE���v�e�M ���ݗ�NqCQP<��_������cE:`j��ڢ���!���������x��i���ٕ7/$�Un���,�m@�^u�.��1ٛ�1][4�������J�qY��[�&=�J2;نN�J���خ������)�Օ�������yf�bo�As2�{�4�Eֻ��N��T�Z.`����N���mm5}(�t%�����B^�&���|�7��i��|J�����=�3h�E_R�ׁn�n�o�[)���ҖS5�qz�4�.:qv#H����8muX�z�*��u3q�z��%��yJ0rZ{'�y�:Wo_h'�Kt����'�T��"����3S;�9��?4���]�a�J�qc�ɐ�]	�%f��]xj�A��t�hW40�$r�ķ2*yz��"s��S�8��<�Zl#��mAZ�=�l8��%����m����3Ӻ��^3|�~L��IFr��P	�D]S��_�׺p-�����6z����r�T� ����4�ԓA'��X���5�kE;���-r���++�E�5��jnc�ī#g$�$Clt��lqI+���_�:-���3"��0=����wniѹ�V:�Z�LW�﮾�<I��ب��g��55�W�RR�;��`V2y�՝Y9"N&� d���[3�^xWr����}�FĢ���&0��w=�B%�y��y�㸜k��`yQ�V�3׶�}��p�[T0����7�a���ː�>���b(��9���y��ա[\P���V�KH��,��]w�dy�f]��l���d�nN�guT][��n���*H.`è�� В���~Wh[�^����=O��|0cm�L�(g#��Ci�uc�<��_���Nڂ�����G�zg�V]R�Y����������W�
���ZK^��+'�֓K���y���}�ߚ���#?M��"w7v-�J�����5)f;���9V2��j�B38ke/�a�_x*���X��뷝��8��H& ��l�p񷟲_D�r	�תr�Ed��$N��fy}��	�ߵ�[��%��G;{��oQT�6wv2��&�"�,[	�����;] ��8/{������
��!{Z���Uw/���I�� ��O;�$�r������� #��L0�8T�J�tkysj7�i���EU���־�6&����U�X4���&��Q��=N�:�NU���&�{MI䔤WOo7�<�N*��Qڇ-�kr�Y���+S��g��CI���cMyL�f,y�UQ��=%�xB}���{,�T���g�{����ca�E��l��Ջ�(v#8;��p�q-�<6>9�ߎ��17GEbQ�fMQ�V/��������~�Vc&�[?�*�]�v��JZ:��n�D�^a����-&�ɿi��g�f��$���RP���!�u�koӦ��������0�j��R��a�ii���Tv�=��ԯ}�{�I���f�}�r��u"h��ұ�[[�Ҹ62w�T�#�iȷٻ8�E��1�r�on�xI(��#�.��7�}Ht�fA��r7���ʝ[o��xq4���.S�/��!�Gk��q���9�Si�'��寝��S���t��ٮ��1��T{���)ma0�rA!H�M�%�	RR0Q~!�,�"����X{��� ?hА�˕>�CXw��;Xb�c�W�]|��@�e������ɼ~��$��Կ�2W�KxI����^�� ѹ�9���;Hz|�C�ڒ�iZE�^���������m��i�%�u'w�wZ<����u!�7yڕw�-i��}�;v�%��{t���|�o2Wm��� �;֨V�6brƴx� ;^��T�]��KkN�t�fᡖ���$P[���œ���Qs�W�xKy�_Fs�g*Q�Ŭ��޸�Z��뵖8��;m�F�Ε�ڶo�b�i '.@v��{5v�f�R�1;����瞚��,�,[֧��u�m�$�s�~����h�&�ݥ>�O}<�V���=��v�aX�>�Q�_o��]b�j�[f�.�!Ƒ`��v��홻n��]�<{�f�K�e�Jd�-��+��p1m�Z�c�kŬ�5g]�v�C�a>9�����6o�gwr�Vdӽ*Qm�lX�6�m�����+q��iz�\�.�8n�}w�7��^���=��O�{�N�mF������G�d�6D:��j5t�"y�?(�!����U�$�R��c'�-��:0�Winr�҂���N��	-d�=�17�A��Ӽ��7�<���SO���%�^ːl��.�(��ٺ�W~�|����}��ʉ�j8>E`㙝s4���d�E�1�y���{�8/�5K��Է�g����]3�2	��1�;@������u��#�Yb��*�M��j��NS�����ri����{R�a�Ξ7Ү�᫑�	�((M�D�U"-mg�,�\9�lд�9˥�{���p_�&*Owk���<���WqW;7�%2Y��㈍��b�/�}�6V�+X�Q��\��g5q�at�B��s#�����4�1=Α������ۇ^C�9�n)-�7F��\9T"��{sך��C�ا)��Mm[h��:K��Y/]s)ݑw,��c9&a�\�5��w����wg8J-��N�=���8 8O6.�fL|�n��ÅoxMU<u�1�WE�n�̚pN��c�Tq������յ��ڲ��s�]9�$��!c;��[I�v���a�	���.��v(��{8W&��uϦCC)��V
���k;�󫠀gn^nЬ��u�l� 2�_��S`ι��e��t�"����m���G(L��@}� u��oaM�P$v~���ù�s%-��g9�~��oo\Zk�.��`f���)�9�
�^Q!����F��ɼ4��OVJ���Zx;�a��8�H��g,�p��)B���t����)�2x{Ϗ��=��W˘ޔk��G}0n�����Cd���FA���n4(8�@G�y����
�Y��(`-�g2n:2Vk�v�\�)�	���T�kC�l������<�Xk_r�D+1ԗ�����[�����\O	YMYC8;s�efq�`r��鸲�y`��XL���-�Jd�]���j�h��H����t�Ι�DJe0r�䛘�S�s�Ȗ��ӻ�G$�������͢�4�3����O��g(��OC*�<b��v�5h�1c����iv��v+�=(�[{
>z{ei�i�Bh���,����b
��+���)0R��FF[0����*\�dE�-!�Ӛ�=j���c��o{܍�هkd.�8�ҭ��e��9����k�oFWi�et}�cw�1��*�6�Z��W5͸�>G��[�� �|pq;9�3Cw/f%W}�E���̢�U���]���bخc�2�ms/�]3٢��6�ae�$�q��e�U�ކ[��CEܰ�&͜f���vSP\��wy���"��W��&o���6��G�v~軈�o�<R�?�cIV �'\r�ZYq��\How��q孄^8/M�|IN��\X�ۿ/����Y�u�u��T���a�V���Ll���r!���y���62q�]1�mz�������
l�M��[�UnU����h�d�b:�i:kt���mZ�deo��.Hu$D`��aɍu|�1ˇ�ou���j��a�z'z�4ˊw՗��RǝU��n��N#���f*�Zr'S��^�N����C֡ ���]�`�U�Q
���6�z�jW�{�%�l��EǢ��w��;ݘ��M7��L�u4�v��n�.V�6���Vf�0���^���/Ev�n/�q��4��;��gy@�3l�מm�#Z�VV���ޓ	t.��w|k�h|�fnI�z�9,ǭvU�Te\ ��A�2�f���,�ήݟZ��p��Zޫ��dT�9X̥ޚ��V�K=H�{�aS���ڲ먑XbJ���`�g�؆��= ���i���� Z
Vj����t�JC[��@Ż��������ݵ��N�ʁ��[�YoB��Q�+^�ќ�F��Q��=ޡ0��0�pJh�tƬi��;,�}\�^uǽF�gAǝ����ʠ[�%������6Wcw4k@���%��KP���~�#}�鋐7b�ε��Ӿ�����Ϫ{^Ƽb�H�Tue��2ޫ�̅2Θ�B�������r�}f,�7���me��=�U^imy�sͻ43�Rv�z���fO�x� c�C������LLsм�����j�R��:��)�p�`�%��0\R�^�1�JU�<O62�:�%�ǥI�q:y�lu��<֡d����7If�q.��pk9uO*��T�48�w�o]f�:7��e{�{�KW0�|�������t��تbo/-ֽ:2�J�&}���-t�����
�,�
ԅ(��y�Ə9@E����ûo @A�U4��L�u�0��.�%��NLc�UYH����{�6�T����q��gn�Ϛ�g�>�
I�T���M�uÛ��D���}_J�Ā=?���铗S;{�Q�nHoa�]��m`yo֧�:�6j�4'���NJ�x�z�j0���Z��ۛ�o8`� ��B�U�ofh���q��򛂸P"�]P�k���wo���^,�gr�4[1�L/�L���i������$W���'z~>���'��gk1��U����v�sk6�@��8�9����Уsb v���v�FS���Df�
��'�{�_���+].�ʈ2���봍��c��@��c�\𱓾2�?�}����\��o^�ڃn0��Y�R�d~ӓB�g�H��v��1}��4^#�D��]mA���0^�X'���h�Zj6�\qH$7?,�Q蘤Ji�4�MP�ח.�U��+�iƯޛc	��p�쒗�T*�Up �w����������&;Dd�k�ˈ�.;-s�z=�a:)w���:�q�ld�P���Xvwwe#g2��m竄�m\�3�p��NuA��`&ݓ����|�slh�9�a[wj^�;u6P�g3�$[*��Ϊ���PY�����[���܎;��Uxj��nuև��톐���Lxu_b�=�:*�v�X�]�f�N��9-�Y�����KO�u�fnN6�w7ƨ��w���i��v��(��k�[��#���"��۾�y8��-�W�Ӆ\���W������,�Ͻ����<�cY���� �w1n�}�4J�bLԟMcFy*���6�<>�{^W��1oՊ5W[i��k�����.��SP�<盓m�O7��י��ӇS��>�֥�3��`��']ґ�cV�r�	_��͑J R
�eL��`�����+��l,��j��͙lK�����E���c����2
�b�{��/=��)f��p��s2�>�װ7B�T��n�u�;��>�p����С�l��r�g�U�B��A��î�t*�� �k�������7��9�x����ښ��^җ���H��ǧqwop7��HY���Z�Vm���+�T�+SR0y�U�I!�rNe���B�r삆�G2��^ۨ�~ ���STw�$(W�#��/R���\�����g�eYc���׫�c��*�St���i1µ�-m�ڛ^���YɼX�ј�96E�s��$	;�D� �)MO���z�WW �������6-�x�W쫂�6���s/r{��2�nw==��.H6��x�8l�H������:�B6l
 ���]��+�gAv�q���H�͵���ۥR����Ԑ.��P�*1*}�|QMq�rߩ�fJ��v9��2�����'AY巴t�vF��V�j+(��ń0
�ce>���<�"�3��s�CWȍt^�m{Z�v�m��8C3��_zx�iRr��WԽ�[\mo�ۑ" ��ɦ�.��[bi3�e�c�����9Զ��x0b�t�N���Þ�ZWTx�_��q�q��Vh��U����������y��W(�!��y���ȉ>ܻ�{y*�B�n�g�-M�Sx\�T¼�RɅ��Ӿ��@�%���g~
�Ҥ[�i��<�Z��S�ʫ��+���?���*���|�o�I�VU�u�L�+z��wkL�c 1m��.�\���S�x��+;iǲ�-җ���vfoN���ap����XT�iU�;�{���gVNf&��OtY��Gui�t�����������O���S�Phuݩ"�vzӮ�Eob�&��Q�%��J�m>�|×�V����U��)bɛ�����۪�}y�/.6�ſ�O���*<\fQx�H�~��?�T�y{ �\�Tٳ�h��)��y�{���y�����Ocaw��pc��&��X2E���(A�m�$I����v�F�������dQ�ǜ$u=���M���T�#qrݖ��e=<*f,T�����b�ۧ.h����6֞=�*Ep��;�'˱���-�<��S==[(���nn��"�݋����Ԯ��!�7�#w\��9:*����0���8����u��n�;��n����rd�u{�dC�7,��)�{np��s����Gk��s��/egٜ�n�S�S�ǳ�N���ݒ�ϰ����7∴�\�w�B}xY� �6n�w�ܦҎv<��0�шb���=�}�s�f���|���Zb����y��oN��o�qm����@O8,G|��G�(3�Z��\��+�#��i�܄�W�V�؜˄����NB���MY�Ӿ�l;��H��0T�CQ���P�%�s{���t��ܻD21)�!ݪ'u2]4n�0 󸛺7���=�/*�߻�{�~� �v�u��1K��H��ٻa��W��Ut.�n�j�Wk5��i�J}��<0r��������H뚄u��J9���. CA �(ҧ�Tg]�H�GgN��Y�z����O���Vs���cn�L�<��Wﮤ��	��u��jS;|}Z�w��3P TPzo��S�Ѓ��#��.�8Jӹy��(�+G^HźJ��׫�k�Y:U����
���mlT�WB��{�j�c�E��pX�D����H�L.��
'�f�̙��Xܸ�r"��u���ӹ������v�}�w{�0���A� ��� �Q��YY�� ,�-~�bb��ې��� �{�"�o��n�еNY��J�6f�����|�R1ڷ���i�[Y ��YW���Z�:��s�>��=�l;�L���]�5T�9�Ova����s����l�+�癋i�`ԍ�}�݌�~�T.l����\bAݛ�y6� f�svH��� ���߯m�9�F�����&�$�g]�5���x��4
Gs�u��*4�L�E.�U;"��3"�֕�6΁]�����e���|m�'���F��+s��v��U��BV�&eD35�Ws"2��XM��f*+u��K���Al�Pe+}g�oՁ�<�	�F޴�c���4��j��-,�#�*�1Ŝ�]b#s/l��a����6B����o��%%���������H����� �ǒæa�P��<J4LڎQX����vv6�J���@�6Z���M��:�
�������s��[}ջ������:��~�i���S����o�qu�eT��nm�0�S}p�U�U�K�&�t��qw��>�3����*������EG����|�G��汞�o$�n��E%��gU�:�x�͈�I�1V'K��N�F�g)5/s�����&6u{[�� �pV���y��5�;�Ԑr��аf���nw}V����h宊�>�O�yx�z9sn�jw�\+<Zq�ͭUo�Ї�j�m8�S%��ԃw�R���Z�����9�@��;�M�vM@��w�wf*ĕE�"R�`�+L�^J�닢3�k.�����`���g7V�Wi��t["v���,T䉁X��n.���QX%/�P�<V�-R����V�^�rA9d�C�,8e�;΂��}=ۿeܸ
���U(��Ets��>0��KQoy)�D�����ku����Wz�=�^<J�1ʳ�r0D:����:rN�
�A��"�]OD��(�Q�L�b���)�=��T��ڱ��9*N\�
��F�j:���Q��-�[�Ƹ���@�87�hL쭔�ޮ�A�JN����݋�C8��%��(���=u�0��3G��Ȋ'�_H�y��>_w���u���o*�L�7uƠ��PH��;��nup�9WQ��lv�PX���ks��>�]2Vjo���r�m߰s��WE��Xv��� -�*:�v�lO��9O�q���~�ʝ=~�"�y��J���7�r���1Lј���jo��Q�;A�W6WN��Um�b�N�;�8

��ܷn�5.ܹr+-��Va'e.*�@w���ʑ"\��{��jt���~X��jtH�40+X�n��^�\\�O��q;�ڵ�q��c�>�����f���<��@��ۂ՛��4�9y]��Qu}��j��A���&����ζ� 2"��3�$�r�p���á�aw_=��*7eMl�dNΧ����s7��r��2�����*
���/�-߲�9����b���u�|M�63��K��錄)�ި�}��\���>�gL�D�^�u���9O%m�o����^�B�c��اqp�(>�#�oH�ɭB����V�=e�-"��I�9Y�9�Y7�!�۳=���W�qP��=U)�p�U��/��{�N��J��ҨΝ�P,�i�]O5T��?A]N8�˷�&�]gf����t�}2#FH
p��`���[�7(�e;�zJٺk.�=�m�����j��7
r.�DT����1+6��#�į
sc�	���5]<��@��)F	�O�c�q�r�[��k�{s J�QU{�n��{�rH�$j�M�Ue[��t.#T��O<�Ŕ��{�[�ߧ�n-s��7&{s{�,�˹^W1��<��vnk��Y���ǻ�+��YҨ��iU��D�c���?��K����J������T|ߴ��Z9[me	Um�����^+�:��B��Q~Yڶ�&�T���X�K�u����8�Ք����ݽ���fR����p���5�'��	��\*��@���.�x�-��j.Me��m�����%ne�����۝�Z_{{Fu�U0�MmݔuQ����;��I�l�i���l�v�MK���E싸���-Q��ҽ�0�Qmpi��D9ݫ��e�6S�k�Õ{�֖l�Kt}<Z����nǋ�ק���l�,��0k�>1R�D��nE���rd�]_a]몼K5��T��֕�SKC]v?i��	�i	8Ŵ�Zn#;���j�
�ۭ��Q�؛ɪ�J��.�޶��7u���[��eepހs*�X1]I�k��69�yA�.���JSx��av������4����eI��]	��<,՘�,G;�k��~ѻ:o`߻���5�4���ʰ}O�QA�ꥶ�C��V�/d�{y�z��*�f����l�޿ZN���+9����.{0MWD���l����eVy�����輹��_��b�
QA����t_����Tҍ��������L���	^���9V���8a�,�1o�LX��ьA�Y��J��_E��#~����&o�+W�`}@��������s!����(������5w���.��>nCY����ݚm���g\F��8F���"L�#�Y��z��`�q�����D޾b���.ٝ[����������}Ϡ�蘣Ɏ��~�\��;�7l�fR�b�ֳ /}c�U��3Q->�y��5C�+���(T7ݵ����gJ{R��nr��M��n�L��(���y���'ﯴ��k�g-r��(ynu.�h��3�@C���]=�>l=��Oj�CPN^Z�U����ɡ�ze��}̵T�D�ʇ���PnkCdܐ56a���'@�N�e�����r���b.zc1�y�%�Q�����N63jT�~�!�5AlMh�sx4u5�Kcտ})�=gi7Ej�燻�t��Z�iB{9ZF��F�Xw9�N�C$�y�N&�S#k��V_�J�;���f'<MRj���w����~1�őQ۲�fv����Y �f���;�]ǟ~2��̩]��}�[��nK��4�o�w{�7^��:���<�fP银�,b���5N7��=�+U��X�^uu�k^i飪��c�=���c�5�Ƙ�5I{R�BZb��I~F�4˾�ˬ���$%�ݕۮ�Isf⨬�>#*����t�5	Oowz���^wmY0��YH
�>st2oh(����۬m���z���v��Z�Z�D�Z�#�8z��#x��r��t�A���%X��S���V�-�MVMUi�X��tg�z�kl:v��);��z�K�97*�r�����?�v� 6��ufP�{�9dh�[�����W��z�
������ح�R���|����n7��9T4��ΆS��{G'
n*�{�I�W}��'�����]
�=Y��\�z<S�*�:�jv^U�թIZ&�H��@�'�r�oS�D��3 ��z�a�PM.��*H�gPx����l�`ͧ�3��ص�����ғi����#��*�/�B������n.��W�=1�����WVsl���m*RU�9ST�Yh�k�m듺�Tt\�ъ�r�]A�r*Q����X�V6woR�^���8F�(>�F.;�ȠZ<O�����q#�[k7ۋ�k�j� �YЇ���c�����:�5Ӻ>��m���u�jѦ��g�����kv�
+PN:6�Y"�V��g3�줶H��gҩ�@p��VG�%�`�NJ�^�h�bo:ߗ�m#A溾a̶����k���IfE��"� 
�7]��@h�EA ��o��$#
`���[�n \��;�P��|	���h�H=e��Ĺ��P��=yz��)54
�qnŴ����h]:����F�WXPAnq��ͣ`z�u�jf
;r�kIoS��;�J1so�V]�`��t��M!�Tn�*��B0���T��c�R4�ٙ*]n,Uc�.�$�Timq�'U���Q,�n�w�M��WAg0ǗR�,��$+)��3G
U����o�
��D1��H97���e�Nl��*���ȋ�8z���Z�DԡH���E��)��a7�i<�۱w%HѰ�$K[�  ��eg��%�"���S��.$w_)���0��ڃ#��v:��J�����a����88��a6�|�S��~�GL+��=��Ķ�e�"n�61c�%������^x9��*}Y�XR�r���Gg�l��5AmT�d�C�w���8�#^���ŗ
Б���K�x�R*0�qWYU\�o<�<��ף�L�Иs:8�!��i���9e��l���'�������/)�r�yc���?w�?�0>�Ovr�r��Δב!�3�.�h�v�CF.Y�J��r�=���O~���c�S�n��D�y{�k�ͣ�O7�Ε�o�j��[�7��s�햁�.C��9�r�I(��]�����Շ��#��:a;#\�%�P_��00n;1	LV�i�Ƃ�?d@�2Oʮ���\�9�b�C�<A�C@�4�n�X�BJr-�Ňj�)�u�(+�p>}�W/�y.}%���rpv|�W�楿}䧔'�J�E /3)b�iq�%�)��[)���}�۶�~G��{�������^P,�I*����\�\BO*�,��]��SCD���7�KT��v��e��x')�"b(�Ail�����f���u�d�ּ����}L�4*��l��v�?SP��E�H�죒��a]��T��Kc+l����4�2"�5^��Z�g�c�R�ݖ8x����i������S��'�uo�*�i�X���&\������d��❡p�Vx}�X����۰zd��q��)�˼KB1���q|{��=���\�M<[�P��� e�hk���2I�f9?�{ѩVon��h����/F�c��>��O81�ٯ����*�**��u���gu�ox�[5�</�����=Zx}D��떰Pw�"�ʷ㵭S/S�_����L�f�E���<�q�]ko�WZ����3�� �r%��t. ���t[��KMȖ4:-B%��D60�/��1��h4{���swؼ�:��Mvp)���C�j������C �@p�i4�������4ǥ��=c��*��fXB�E#(괒LCO����T��3_}���
O"�x��Y!=D>2���v�����;Cp��hXauƌ4��^�qj�R�a��
�"�.�h,_ �p��Z!S���HR2�����H�!�K<�FB
�Ux��㢻.1V)�h�c��t�S���R���`�=�g�d��y��ֺ��T85ϼ�V�|xO�<@�i�TgFݔ���,\�H^T7q�b�������6A���v����� �x���+�8������Q'�̃����w��S8�i4���w;Cc:g- ���k�m uG�+�Cj��W�oyev�X{�R5k���C���f�&�z�]˫Y�y{�b�x�������+䊟8"YH΋wmئ��F�p��2����3>�V9�`���z�A�K0U��F�;F=2�N삟�T�.��N� �,��+��z٧��n�3��,�-v��̵\��\>��~�W	���z&�{ 5���NT�Aq4*��HHwzn�����Uͱ�r��-�9dkh��s}�������=�ie�I���UsMYa\0~����v�ò���ͲrQޭ����&�u=�T��Z��"��rzٙ�	�v������*sD˹��W��t��5<{���f�Bp)����Aj}�f_��ӫry� O���|X��vXM��,2[�#��ƞ�$- ���&.���'��9%���aT������S�9ԍ�B�9���nS���ׄ#.n�|>8V�@����^�Zhq3��v!��>A-���ΐ��H������zV�s��f�^�@���h�W�r�(�ϫϲ2ǐ�h�x��J���\���Gf]��0��Oe�ʭ�K `����k~��IA�>����6�tr��g\Q��gz�G{4���vfV��9���,r�S�����n	n8ͤI՚j�3�	���T9�U�m��������c=*�$���Ҭ����H��m8-f�fv�� &2��@W�W}S�a�KH�zn;��	3���y���T���'y5&}M�#��1/y�:�c�/2��ׂi�HD����Ժ�,��]��cő3�r�;:�������o���9b�!�B�E�D��K	c�ת���N��z&\�6e����Ǿ8�����]효. �����4+��u"!���q��w�ԫ���驘�4}��vJ���#�y��"�h�Ǡ �+1��H���8����sE������QO��˙�Q0���T(��`�q*I���5pd{q@y;Ŗ	@����J�h0�3�P�;��0��n�����.���l�G('7�^l����C�e=9B/�l��AEj ϡY��˕c�c��9�f%��ľ�v7:�j������x���~Y_\H�,�I��7��&iG<��z��s�L��������x�h){��T���Z������͛�\f]��,�S��v ��%Q�)�I�ڬ�~�ܼL��QMm�f\�*���{/�B�>�]}�F�A�w[�>�Wf��Y�r[��]lC̳A��6�-�j5��9�;d��-�2��;�Z�W*���������-c^vn�*d+`�}�n��	��`/�n���-��F��jB~R�~����D��3����n��nŖ��W�^t�l�L#�^�i�Uԅ�%�t���(��=PV��@LAh�
��Ν���
�Kd�1�X�:|�SYb/s{]]�F����ܝn��Q�X&l�|����� �l���U��Q﭅�9����(u�M�rv;KW���d!�W�c!Y"*e�c�(�PL(>g��?g��}��Z�P��>u ��5I�|�F��p2aַ*E�c�PA�L��,��[��Ff:o�,U��������V����G� w�����L��
���Qfu��Q��y�s�yޅ�of���;���=��ѾrE��x,J�i�~��Q���|��MKD��2gm)�!�sQ��&V�p�¶� �H�Da��~��z����>8n�B ��`ީE��ww2��:l��7ގ����J�Wɘ��`]�rn��ٲ�$#�Y�2-���5 ]:��^x{��#W����Ǽ����k�}����$�qF�9��^��ߐ!�X���▨Q�_ۇ��c(���.�h�-�4$K�9��������d*~�D^P�p _k���<�}2�bI��I+����b��K�1Ȭ)��qTS�E�C� gQ��'����oMo�=�qݯ�i�Y.�%�x�B;^)�Q�yp�Rwoj�����.�Uv�fT�#}Ǹ���)u�����7���G�<1�B���FYJ��$������Z7���2S�kF9�2�+n���aV(g�I?0tv�++듁��M��|�`���٦Bh��AT��A&�/N��?�f�袏ť�3���A��+L	��A��(6%���g�&�Ƈ0�]vN��#O�/����1u�@�6Mb	����9����%�*	�� ���(N}���'X=��Pv8J����li��`_F�T<S�H�-e��u5j����-F��moj��ױw�����
#OG�6��-SA��X�T]s�f��꓌��:���1��S$�V-����}*��v�6Oa�4�ʂY�]�qj��qs�LC��$�Lb������s�u�c��k"��!�$aK�n�B�`{�o��N[�4�4��@W�g�|N�s��Ш<�t�x��lg5�����v��*����S������Lk��1��6���Q�Ɉc9��[�bI$�A�[�eM�e��3��,�c�u���gǳa}�X��ʒ�)���}y���s��N>��m����%�{3)xu{��U��"b��eP �?_����]�|)CE�����~S fi8S^���{+�i�Lp�R^fTτ�W�U�`�+D�-=�-/�y�|s���߇0��yS�<"����n��vx��BV6��U�H-	�
���V���?����<m<{U񧮭-m��/��F<eǵ敵�^�ث�dyF2q�h��9۽<�d���{`Ԩ�<Dŉ@��Z0{+�[� f_��D:�Q t|&�}�t0�|��!����cd���t��t4�\2��Gh�v�<y�����o��®n�(�V�N��%���1�{+
@���csW�����wI�r��Ju�l�Ҭ����� �q��`g^d㶠�I�#�﮽4�)�cY��a����v�Q7c�����~�h�䗨�#���
�M?fך�l��\���bd<P�sfY�g]8��|bq^ݻc�`F��c�-��'Ɣ�� �����1-F��KG�)�w,�5n�w���@�w#4E���3�w���&]W��������q/j�Ŝ\ѧ��F
�}�� <�Ɯ��XV��[���on�¾��w,_lwb$��_a�r3^�q`FZ��2�ǽ�D�f�F�hd{4)Q��ts]z�C��W_�����1!m�y�9[�8����M��!�ϻ�|�c%��C_����殼	x�Dَ
ײ:�8�J���X@��/b6@"��Kf�%�T5M�B7j�$
d��-8K߁$���~v�%���?-|Vq��=��!-_���(���������O~�
V{�fz�V*��өh�ɉf��f\]@ ����ڡ������i%(a�P|��<)lt�K���<C�G*}�)�����
�L�Ct���>���<�A[�ڧ�e��%u^G!�ֆk5�=&��jw��k8��=��s�c�$�4F칅�^�[lE�+��c!�[+G;F�F�.��s��H��!6�d�G�tكȍ�x��U����\7�뙥`��%��a��
�שk��UH�`˾ټ�X���ch:T&f���<C6!��[�:;,�@��ڇ����	c��*fshuE�l���\}�Ԥ�Н�5�S|��o��i���W.�l���}�!>?A�NǍ63~�b�z26�O�.�
�\z��W	����Y���Ԛ}�'�x�R���LHܘ4^�O1��l��/����<
A�]Mmm�X2�[@��i�NB�h��=^���Ң�:&�lA]���.��聠=&�/D��Οe��V��;�tab���W�}<
<%�L
r��e�Ⱥ��ֲ�O���y��.���a?Ǜ�C�V�\r�ՙ�\���L�h'�p�:u�P��h�}�vO����5l���&>�SO�x(x��.� ��b/L_������N��t�����1> o̋����=�_etYwq�>
����ih���e=u~��CA�����,72L썙>�C8>o�
U�,����:�7�)���yf��hG����l_IҞ{���`d�U��<�E�t���m�|lS��k=v ����P.�q���M�)��Yz�<�3�{�i ��4Q�'!�|��L$.ϫ�&���| ^4�WX��Ă.�k5G�-?(r�}���K�lU<Ѿ��[��v��̘e������U�٢������%�}�B����x91M��<���Ύۘz���2�Ҕ��K*�<���J�;#��^�7<S�$6�q�K�ē�n��vR�v]jvr���	S�����Bs˽
-���^����.��)M�]@�=7���Ż�Uܨ���o�Oᳵ�E���Z*}��m"�Y� ��e[[��"�q�G#��{�֠����]w�ٚ�����=�0t*���X\~E
gZ��9�����|+@c���Z�h쮱�)j��I1 �����OЙF�����c�/�HZP6�9�r��{��8|U+p��0ǫ��W�cL� ����#+�ߗ�g���WP{Ns�_6�O��]�� g���;3�O�cM�|<��1��+�IT\�ve}��kd��X���gk�=ޒ�T���֠��!q=��B��-�6���^�#(;o,�u���\���7Oדkou�:�$�:}�=o�fE�8�%�F�R�B�9���Ll����3���s�賮>|�?L��-&�1���k᯲�b��
N�]��P��M���������ݥPz����9��C�ϻw;�����i�+�!0���MUwe��U�H7�R���Jk&�c&�]�>]yP)fcz�����m��5���Cc֩��L"1�J���.7�_H�ӊ�T����aglMS̳e;��ܼ��e_b�y��-�)��X̖�n�}u�t��=�"��{vc·��@oM���-l����7P�hiN��8��v�Gq�]˂y�S"�ի��:l�,���ٸ��F��w�(� ��{���k���͒yn㰞7aT1�'�2É�\/��};�$x_	�\�n�H��b=��=⿗3R�蛂����p�U�G����7U4�l���扚���[sD,��f#���+Bh�(��3G��?�C�8+��c�ϛ3�vQ�{<��PH\z��7U�^���NBӹ'�Ŝ�\��(Q
H��vY���K��_�R�>C�ىg��َ�8Fط��p�������B�ϼ���ɓ������eL�U�g���!�zE6{��Z��l�
!��+���[@�ا��C $T��M ro33]�c�CY�lN���96�/��GA�N�bd��-q�e��_��C�w�q�U-��X�;��0ѝ���Q�B�5��"�6���Q�!���)��Zn�IS���|��m�Z�mn�f�(1���il��MɔQ�ؗ�TW���R"v��b��ZLC�F[�yfw��u����q�B���ϲ���?����;�|S���;v��;�m�j���\[p���ô�n�&���=��L���N�N��o��t��;O�+k��!�;�-�zu��)��,�`̹Y�������)о1]�h�/5���_gM�#H��C�&�ņt@Q�ƞ�z޿��Zk�Vݚe[2E:��b!��.Qa��?W��-�E�(G8s{�s�Ae��^nc��Ü�/7��7B/�K=i�Kw�j,8C:��.�E��p�;�M.D�_,���	��<і�s��/ض���R�ǎ����4r����ĺ��������<�9�Fݜ�7�'Z�;768������o�2�8��W[�����ZnwX��f�ַ��˸��*������^?�r��d��?�U���*8g	�6+/�^��v�xh�:߅|�d���5hk����v���������8Qg����L@�vͩ:��2���Z��1�S���Vm�Y�hi�ݵ�r[��^�=kV7@l�{0�c(���!��٨\�ɠ
P�{�ӗA|�����
��u�.Y�W{>h][:�����O:*�k�f�k�,�y���L�&\�R�qs< �ݪQ�0��9B���-�ڌS:{zi��­ִA��N:4ö���0��(^$Z�:����D6��Z5���b�q���ٚ`���ǘqw���/fB)���C,�A�e��N������v2Ѫ챺4�lu�;�������܉������{S'��Z�gߧ>�	�~�����]8--OK&�N/,�����͍���O}�?�v��mϮ���V;� ��6��j�XM|�0<��W�(�C��� ���+�be<�3���	i:�%ҵ	����k���1t�ཱྀ6-p��a]�D���<�5!�8�>5Ϗ!����Wټ5Fqh�j��§Ύt�>9ɞ�	�ߋ�~m{�٤�������%��M���M��ŔuVoA�Dz���Ѡ��X�OT�6�Xy"���5R������x����M�ѓ�+�j�'o&�-��ԶV���_u<ڔ�م헑!X��j�撢�]�P��u%�/������	���}�Vc9�u��t�9�&��g.ՙ}j4U����sʥh<��v��qiwɇ�0��a����t.Cjn�	]W�CE<�J�C�6wY��[��3Nuop�/k�mmvU�v{ ��x��[�R�gPYʺ!�'��z�\�(��O��;2��&��u.g��HW��Y%7���r�o���ݕNȽ�G'�a+��l��j�Y�)��m��(Agn+v��\[<��*��֭���/Xbwef���w�%ji�[����(b�2땈��ҽcPJ�{[���Ԯ{G��ܗ�L����;!}��:�csS"4��u+�_@h���e���6i���m1�]&��e�6L�@-�����p�&���~��$z1���LH���������칩�� a�b��/��o���ͬ7v�l:����MS�ƭl�wm��6�#�TOX]M�W7*[���u��'�bͬ��u-��܏n�O��5���&�+���e��Onm<vgB��pf����{k9��;�y#S�pg�WY�d"�bK�g�g����U�.���}W{��g����{Vr�L����uv�{t�E�����7-$lj�9��-��p�B����k�%���Ś �@�z;f��~��<���]��$��H�}$�ݻ���gfF�	�<�.T�	5�Yo���ܰ��2SO��[(��I�[�%�יB4f\�H�_
���N<Gu�:P'�X�bP$�ȓ�:�+Zr�]�ݭȞ;����WN�"q,�
���%N���JZ2B�	��c�l�u6�L�}ɒ�q#U�y���H-J6k8tt������'>�zQ�Py�x�i?m+�5��ʰ;:�uk�7�4���V�R��x�����Js����c�	ڮ�)���<l�7H�ߦ\��'��+��u�XOpGv��B�l��U�$��g��8F[�{fc(�C��&r�.�TI���@r��ZΌ�����\����2.��0�-Ѯ� �-k�׽�ov��ӓ�.TF��l�3��7��S�s�L��IX���ȩ��S/���33��U�;_n�,\\c�-\{s�{�� �zBs���9�V�p؁c���	��Jn�˜��y�6}�w�<*L����#<�k�������#��N�$�'!���<�i���zKg1SD�f�ږ hz9�D���?.�#�)��3iSO���Ч�~$�8��,\�~\���cB����P�Q��8O�������w�WE���GM�[l�r���dǣleu�P����2��
q̮�^+8X�"����w�n��roJ��>1��#��c�Ow��YT�Y�\����X�x�RCf��?�z|�=���9��F�i��ꊴ�|q�/Qɏ]'ƹ7(ӷ���d%�I���A�"{u�P�yWN�q3��\�k�&`�� X�ւ
�<ߤ�o��Ų���]y���k3]�>ꘘ�~��2�bk�j���.}�Q�ge,yzTۀ6[���`�NjVy^	�b/��f1b�Ed�fR���7E@E��|'*�Y�����w�ޕ�ƓV���UsS�y=>�@��D<���\ �M��<�]{�~�צ�l�tYx��RwG""&��M5܀�����Է�du��nrv����n����z�7������u�	]fv�4�R��0S ������gD+�?��F�_\)�㔫p��Mb�J7��kw���`�xW���ϩ.@���l�K}�!B��s������e��Fnx f�%�10mk�w�h�Sf*���ʞ	���P'6����ln3)�fT�=ϯ"f�&s�mߞ�ec��R�*�@�j�6ȇD Ӕ���,��������2c�b�؂�ڏy3;�5l��M�!�K1��=Q5ل�jd����z�۩x{��SN�C�\[tX[���;�Ix���r=���[(�L�Q�<�4�_9��̼G�8ǚ4��^�d6ܯH���S��j4���ˎ�Δ�E��Ժ�(���7;��f��n%��#|C��f�A��4
m��=��5�]zꂆ�S�ȗq�����:	��iZ��k<��<=cKK���^�jLZ�m9�hjB�1s֢�	�yN��Ȝ�-�q��1�eb�n�D�S���!�Ž?#CJ���pp�k�mvTɤc����q��Q��vF�u{��뵡��z��:T�a]|~����ʷ|�ݤ=�)���ϭ�UEy`M�CK�Q{G��t��J������k`��Ʉ�jd�b�v66.}l�D�����O�·�z�|x���7W���=2s/��*VU͖����f�:��Uz��$ɑ�I#�~-��E�[��a��7�ZI�,��S�f�m2O��N@j�	㪫#��5�_�.ʑ�9��ͯ~�&e�)����oeb9��F�u8\h���G �bK5x)Iq�� oD�Y!ڐ1���\Ȇ�~�w�,+��p�	�չ�������g��D%QZ S�&Lŵ;F�+�$�^�-~�8ͬ�i���.���$}��,Z-�Z��dVH���R��5r=d+�!�}���f�ƺ�
T)m'�����s��[���91�9H�=.�!�|E0�*��$��Q�k3�Tyλ����'g��k;��~@/q�x}���Q�t�&�Az��lOe'~�������p�N�5����=KD.�x@t���xYR���@��̋��l���/�)#��};~��|��� }���I���:n�-zK�f3WI�U0�iϐ���TN�
w�=���y��������H*�x#��I)7�k��:�Ed���g���Fn�p(�����!'�^*�&S:����G�����Cb���ό�^�*P��·ؼ(1ʶ}�C�����U�h��g��o��� �W
�X���_}����IAxخ�6�&nCu��6b��E`��~]f	����:9�ݣ�(�}u4~��eZ�r�@kgίM��
W(�����y��X�/7���܊������J���5�N���7}��eB�9���@_}��%�B:B�QP���g�{���եX�dVL_}��:�ܷ4hcMGN�Z��>��z]��ɛxA��
�-o�>ۆP:���,$���ǆznBb�
9�	9�#�{�]�3��h��8��8o�ӏG�7\�v.�ݞ�����i*��+6u҉��:-�ǒ��̣���K�Δ�Z󉥶�d��!*�x�݂��P�t��f��F0<��>�}�vl����A������r"�}|������Q��(�
^��m�6�Z�!?�궥w���hr���l�����&+)��T��W.nJ����@`�^�:n�Ǹzna�������n;��H����6������3FM��l�b��x�'�1v�������ѭ ��ǷM
���+6m��t�����L�p��F�vvފ�mu�8i�j<�nZ]��-n._���#�v3Tvk���c�l���P�U���ov�щ*ρ�]��5 ���w��_��J:�3��.[�]5@gG����u���FԬ[�-�-��IW��*m ��N�z����I��X��j��R}�\�RxI�[����Uȶ�q�����ъڤ�$ E��lD��?}[�V*��.ӜQ�<ǇLO�����������e;Д>��m�N]Р��'�|�r�qr-�91�����P]��B=]H�_T4�>�hs�ce����}Q�ӯ��pz>�o�2\ή�s8�X=C�F��xM�8�j=0"�����m���s�ԸB2��ϓ�豯��N�+�����Ԯ�GSd����j���>�g�3����� �d�mn���먹}�|��	�uH;�#O��Ò����M}�4�Z���7"m�wdJ�y��x�&�YWȯ�_����������o������6�����9��mPU����ѭ�G�d�Cu����\Kh���R���H��,�7���V�g�c���q55���{��80�ʉ 4w��5V��ըv�����s��,�ӝ3':�w����k��=4���31��S��Z6D;ch���l.��ݸ�;��8^���bxR�����	�~�Vqӱ��μ
GM=>�s���X�!ұ�N�ɤ��r�k�Һ<{��9�Z�W����J��s�F��*��Mצ��=u��'��P/=[�a��N]����Ru;`�����>�4�¦H�Ca����k�n$�+��>�Ʉί�JC���,�C�6��}<�_�=�	_LU��=�[�Lz�۾ڋ��E-K����)��F�{�-ښ��Uv6�x�{[&�Ҫ�ʥ�g`��&N��,T�i-f���p��3�E�ڶ�4�9}��1w���^._��ze.4��E�_z,�������-K+��U�| ˋ�pkXe�2xT�}�X.���o�W[C�t="��.!]�y_)E3>���$E�S�c>.�@z0������j]
�k������m�r����P��}JS2�wo.�Pl7/��*\:�Q���mY����x0��ꇉ�}WCs����0ឲ������0�T�t�
ܬ�^8P&�3O��on����ֻ2Y����d�L_b��P���0�ܢ�E�;� ڴj�\x39�����_Q���u��ik_r����c�_a _�n����"� gL�[���3=%�U`�D��0\����)�����>*BF�:OKD]�s��a\y�X�6vN6�vv��OV0TC�<ZИgg��v[&�5a��O������.ֻ������#<i�n�D���Y�e�._�}�C�S������I�x�R��7m4ޙa��N�~�2���:W�s$n�mVf�m�.�QUMB�n,t�0gԎ01����r�[��a|�������뫣��̢5�n�;�\�w;�kB�e���W��6����]�dA��N�3���Q�<�]g`^�U_m�|�Ҟ����8���[�d�A�|T�෧e�+&�eC�ă�ڗ�m��
,6�k���K�C�^�^���41�� Tⱙ'{�|�|h<�+��X� �Ӆ�T�zf��'�����g�kO��,�J�Ԛ ��фû�SSH~��f�U%�P���\޶e�{e���([��v&Kɹ�8�%��s�YHwH��Y�BOams��H�!v�f�8ˎ�6���6��T�Oi���k�+~�
RyZS9�0��%@�Q,9�۬�a
�h_Sf�,B8�Eū�G�"}�/�����oF��>' �)֐oc=���"��	U�9,	�ngvu�Iw=��k��,��Sk.v�<x�=o�۳������ъSS:���X��	��L��I\D,�w�>��
�K�'?p��&��4-�wh،���4��;$�e6[����Y��a��f���8L�R�\��VuU��ߛ�V��D��8y�� ����%��e�V��I`Cb���h���w��f�Њ<e��Ad�i���E��8D��k��4�n�.f��`A~y��ƍ���چ�Z��<0J��X�l�hA�jkZ����}��e���qn��̩���Ӳ�uڐj��27�q���
}o��D��)X�KG�;=��RUT�����Ӟ��c$��9�u�������+{�a����Ϧ����Y�u�8����I�"��>����=��bT(�nBo1i)5��k-��ڗ��[���_lu�LJ��r���W�y�}��ה�ཻ�����i�5�*��K��b�)��Hb3��Gn��ԉxsC�6ze*#��t�L����X����ߩ3y�Wx�jZE�1�17�lQa���OQ<��5�P�оe ��V]�6�wѬX@7�Զ��o(����sK7
d�� �&0�wB�t�BcL��f�%)cew�Ѯ�Hc�F�Ϭ�;ޫy�UD=��{g�\�l]wf�e�'�iܝ0�/�BQ���4(����5*�4���ٻp��șk>��w4A�TΕ�
��jm�ʧ 6�D��I��j��,� NQ������w��n�ozgƞ�*40���؝��-�w�T�(@)3�����8��R�k79L���6��biS:��y���n��H�ӆ�o� 6�2�/([o%S{�s�-��L�(�AW�K\�q@��z.�S�"�\���NAG�QQ��(�]�]Vˠa�]��a](
�9�.�L��M�Jˣ��ԟt��w�����;�#���J�WӴF�f]"J4o��6�=h~�n��^��C����x�ꤍ��3�T��qwY��e�MwA��\K��~J�;7KI�z9+`��n��!�a*��1W��X�S ���<
|r��"D��Vj�|:�Վ��'��I���2��:���`���=;���3��9�^�9�0TĆ����#���ҘǪ��[݆!�IB�>f�tǈ�kv2 ڮ[1nk�6��`Wd�9��M�����~�:��>#�_ٜ�J��C�=���9b8I�KdpuA�������?cc�>�>>^��H��\��e�ߨ�Nw��`��g��$Q44�^�{o��M�Ȧ�X=�=Û�ik1�cFf��	ٽŊ����{<�3����a�+~�x���	ܢ▌�I~2��M:�$�z�U��se�Һ�?�������{J�}v�斃z�'���.�Ť�q��X�)�*�:���tp��U�z��=�1��p��,��YB_�%�IM^�`Β��s8>��]Z����j�{X�/t50�h���K2�QȔ<9��'�c�^�SaP�[�]1�N���.���r�V����l�Q�}V��bZI���J}����}��_T;��kD��ђ\4�G�+ߤ����2���E	��+o��ۍ`���E��o����h��P���u�w��F{.��5�m!Z/i)+�غ��[�5Y������%��,��< �bx�&��4+U�0��;��������.�˯,߈�zC�̿
IM#z�\��ܧq3��D٨/|v8�zT��2|�䖶�x�V�u��I�ALXPUi?v���}XO��^���T =��lo�8k+1vX<L�ܙ�1�"S�&tH;2�ˮ˓�sӖ#fځK�h���&��Pd��/��˪G,�ԭ�I��SJc����]H�6�ii�p�z-�$>W:�8��-���6� H�m{�g�t���e ���7�Җ�YC�6�bb&]ܙ~���� 5%��f�V����w`w*k��-G��\\�#n*�_Y�6}�>�L�tn�J~���Һ�q�:������]	O њ�<����C+U=��a�s�}�e�$8$�����G�C�FV*� �I�����%ݪg� ���d�2��D6�����n��7�g}AX@���y�̥SvJ��Ck'ۜ<�g,�mM��I���b�:�[��o#Ǭ:%�����I���~\���'���x�\F�<����F���,�Cz���j^����V�W&����F����Ƈ	�]%�{��;�Xf"/x	����J7K�i�1���K�z�ݠ ��Kw��t���W��o�tˠ]��E�V�� 6U�k}V0�sP8*��wc�M:t2���.�c}���c�Y�r��yr�a�:F�]��~�v�b�=��pN:� �2n���6}�|���C�g�C^�dJ,��3��¾ʛ�m�����r�d��+�KH�[/���/}{�r[�Q���ſ���ة�h�BO&ٍ�Bʚ$��m�`��.;��k�X74��Y]��b�\���]�J����f돍���;��1�Ea0�C}��U��{�xN,�S]�z���$��D�L���r�toIw�,�Ѓ�T�`j���v~F}�i��g���Y����A>t_lW5Y�L}�����%�-�����G����)?��{3;(���H�+s^ҋ�{�Μ�5�����0D/��┼ڽ���oe�wS�J<�l8���\b�O�^-G�-*�H��vK*�e��2����(���;�{�J?��z�b��Wnj��`�*R��-ʒ����%�SLK�D��b��R8�v�R��[a2��LjN��kɁ:)2OJ��Ŀ`�u��,�\�qN�Y�b��&�`��甸�M�^eM�}�7�#�-�V���~Q�p:�n4:Th �(0��T���Β�	�ڊ�ҟ}��3��*W�����J9Jq��Ɩ�{'�+����ga��k��4 �UU� P�����H���J�UUP��F���(P��TPB� P UEP P�O�� *��g�ߨ@
����� (
 
@P��� �UU~�_��+���� �UUw���������c��
�( H �*�
� P��MPUT ����� �UUu����@
 UUW�#������ *���/�B��UUu (UU_�� *����(UU_�_��}5؂P�UU�z� ���ο/�_�@
 UUW�(@
�������u��q��UT�� ����@
����D (UUY��?�1AY&SY��% Y�pP��3'� b6[�:aLڊ�e.��H��U ����.�R�� �B��R��RR�TU;4��Z��`�e��vʝw1!mha��
�"D�E((��������U���Q*(R�l�TEJ*�H@!�% E%$P"*J��J��VƐ*����
JT�	l�EM��m����|�����i_|秶}:��]Т�.!�W�K�(�^ћg��<�{�uJswL*n�ܯZמ��=6ȫs*��we}�t�Y�� � 1  :뾠D��� q4q P{��{ �` R��� [�EP3�  b{  y�  ng� 6��@��
Ҵj��ER�RJ�U
�I�I�  ��   �` ��  <��� �.x���  �`w�  =� �� �4  �ء�� @ >{�*��� �� �F�ӻf�H��p���+yܧ�:c�^�U��}̧K<��VŦ�NY#���rt����z�fOMMd3q�P�K���w�o���b���mM�.m+�l��:}:��   �ϥU(�� *D��R��{KFm���gJ��E�n�֍��ݠQ������C<>��)�m��b�zӥ���tS�E����٨U���(�=���ןw\�'���k���M��EE�@[�������[��X�j�z!�֊�ks�$u��=�i��0=�������[CP�RH��{mao{�{�&��(������m���>z�I@R����6׏�T��J�D
��S��挧�w��`9�*��r:�{���U�U�
P9ה��n��}n��|sE�[�+�a�Hzx�յ}t�y���RC�H:�m����yJ�A�@hT�&.�/=�֛X0� �\��km��Ê���m�7f�R\Cu�mj���m��e-�x���{��F��@JnsN����n����[sr�
I
 r)���*EU$H��R��9��T[��U�ֽ�w������ׇ�}���7m��O��D\�
=��o_h��iw��f�lkl�ev�ٶZ���yI��=[���[bS޽��M  ��Mk{�*G�5޽��m��9�TQ�)�5�;׆+F��n�M-�޽���cb�\�0P��=H���Nwq���޷{j����fU��y=R@O�*U@ "��Ȕ�L� 5S�2���F ��U*)P  �*T
�F ��D�5OP x���}?U�u�~�>c������O���/�$T#��e�iO�9�� �9΀��^s���s�����p�9�� �9�ߜ�� s����pp 9�p�p�89��������I�N�~����0�hn�j94��Y�@��@��\�\_e��Ŵ�U�t,֊`�.�k��{���e8�����R���kP
�7�x~�W�`�}n�7�{@��f���!�	Z����9x��s��XTӦ�X,�`��%�&�6��F�+��8������w�zZ@�PЏLa�X�,n-� d#����Ŵjn}I��Fm�J� ~C�Y�1�9/e%�Pת�����i�rX���A�՛�_8z����4�2�' �@c_U���Ǚ➃�x�Ҡ�@����N���y��ے�MN�S�C'�~آ/lֵ�Ƽ��Z8t㽪A�0��)VA�P����X!�{��"�oV�iF��PE!B�-�|0��cT��55�hV�6��@�)i��:���A�L��˅3E���������i��Ԁ�j���dg2��>��Z~���Ʌ�-C�&/\4Ex|����x���CjՑ�<�6X��S5Bf�����EM���h�)�B���%�k*��x���c���{�OY�OA�B=��($����K�ب��ի�����Qau�˿��k �L܋u뻹r�Yz��dĞ��S٤�c	h��t�*��.�\��y4�@�*�4��6]@u�I/D;1��;���7(�yVM)�.+	P�Y4�q�~2ac-��?f�߆��:>g��/NҶ�^;�&�b��*T��P��l-}��c<�sVUĬkS!�Ψ/sp@�����T��-�ߥ($Uk�1JGL���j6K4�\l�E��j��&��AvbQ�:�m
��p�F�OP,+�U@ء��iBdv��J�M�&�fUݡ"��im�2�J�i�+����H�g7R���(�\׸���&�f�yt@)Sm� oAv܍|H�B"�9�%F���c/,�!�X0�V\��MXn\l��'H]m��11#�.�F�f�#&�U�-|�/jB�VS�A�B�f�1�r��!���S)�Z̪n⬖�*�h�x���i��r�"VX\�,ᆪ����'�� C�Yz�Zn�ۨ���1�ѕ��nMoV��٭��4��6�YW�D�7X�Ҕ�P�")*[�b4��[s��1�yZV��˨��F�=�����UQ�v���,7�AB�vӻo�c������9���v*�)�@͘\���h�:�n�܁+����u������
�t�^l�l�#�3t9���ơzc$-v7Zv�j�V��,�)k0hU���*�N�R��� ��LlKm<a�-���' �7sj��"�Rl
�f���Oqf2�Um�;+V��2�k�b8躚�c�W��h#aHP���t2����"�D)��5�M��`~��2	<r>Aj�q�&h6�R��"���.e��/&�c/q�-�u�����U��rb��Z�P�uX��,LFŖ�x�!�/i@`����X�ܦ�� �3�^м�ڍ�+u�X�V�Q�Z4�{��:�pf�HW(;͵>WbK�'x��f����� V���nYZ�CT4σ8�B������LR�J3�L�-��Hޛ�V帳.lˌ��]����V�Sx�f޹(�j{L�dP����n�Ţ������T�U5�	;a^(�����Qa��'B�Ҳ�ị9$�0^T�J�n(�%:�
<�*��If(/M(>�/���v#0Um��kzq�^��cZ�$Xi,I`��ƕ�L� ��"���^���Si�z�dl�$ϳ	���[G;%]�N�̕��[�[Gݢ��L�gV�%�Sq�O`�ٛx��Ѥ,&�#!I��Y!9j&��ڐc���&� f\ݬ[�{�gtF�!�e��m�cm�%)SQa'�eօQ"+uHe,��o�t���x��ѕ�4��7�l����$������	A���5��VɠH)$f�fe�Є�{�U�^e*WNL�pAeD�K��6�f�5�ʔ�ޛWL��Nn��ZnT �)��̸�́�p����U,ӛQ;�ZA�4U6`��h�G�D��q��2<��؟"�����v����1�lY�F�4�{u�Q����1�����æ`�m�$%L 7�c;���U�5���-�'r�Ҁ�P���F`y�r�Y{3m�T�iӕ��7��4��ee-M��ٚ�՝�LҁD��)�TF�6�VA��-�t72�3�,G��ɻOM�2Vf�F�����ƪ92��Ve쌛t[n�V�^�c662M���*#�m+iAE2����e�d]�]�j*�f�N�7oCz
+6��A�sSܡrSD62��oeCs@�Ӎ�8n�ѕ�x����qۨa�^�YD��-b�a�0��we6�ӭ�p�d���IT��n������Q��&��M:�n�R��\�)Qb�T���7t���P�[4E�ʨd�V8-�175PSLTh8��$���U��ˬ"������[���e�˒ ��Xt���W�l��yMt.�d\rϥ��
����U�I��� �eeܻ��l6J�p\bl��x��ێ���/v\509r�ƳgH̛$#��U��[���5�a�@��rD&��ōJ�F�k�=��ؔB��q��xN��մ-7h8�.��&��56���v+2���	� ���H��y��5�W�5�M�w���6_Vʷ�#-�5��n�0:����sB!�'��Gl��ͤ�E�jX�x7_Fg��D�J��,Ò��¬�����<�3RT&�b��-fƎ"��ukY��ܭ���LǢP6ۣ��X�ʳ�S�*�:b4^L4wEh*�q��7o*��p��h������47�yA��q��m�o,f��ԭ��@^����ɷe��;Y#��{`�F [5[�/A
Q�W������YF���F��g���Z�sM{&�x�Qɫ������ÇZ��/73��w�S��u}W]�g&|���Ve�]5Wa�NǮ��5��n;��Y`����Α0��c����1B�ָ3��h]��t!�V�cc���3^]�0�N��T��So��6�Z2d Y�bۦ9+X{\�&�^��35SÎ�	��[�%�B����̼�F�P�[qM�Ⱥ�/t��{���:��@�ݭ�b6@��3�u������樫o^d�%�twUK����pm�O���Ȯs++mxe�Y�ɓH��0
��?!YV�a�\8u˽e7��f=��k[����[Df����$i��,P��ZnM�xU�6xsu���q��0:Y�Em�6�6�,��m�M�2�n��N�����ՕaP4V	V4YR��y�Y�!e��s.�Lj�Җ^?�d��)���j���Ո���5��A�zV�js.˭v�(vm�%x,�$;�V��t�đX-˰�c`��v�R�a��`*�7��w3M���*J��:� 6]�qDX��87������5X�j��I\ƍj!I�>F.d ��(�2��S ݲ5<Q͙�җ3r6 �B�
=u$��m�ʼ��+AEV'al���e�p���SU����5-�tmn:E0�l87s�ܡ���F�t抴��J��ۂ��������^�KW�K&"�1�����3�ʃY��{vۥ$�V��5��0c����t�Zd�̪����OpV1b)[N�-W����T���(l�VD.xl���6�w���N]��0$�2��Q�esB��p^��WنS����>Y�c@��/7)��>�YYm��Z$؋��x,�*��x�zCVI�5%R`��Y���.��,^5�,VJ�m���4�5���/-�	4��u����Q��(�F:�1��ۺ�s ��[ci�	I�mY�������\��/p��QL�֚�m��{HDF�D�P�me�tVJ4��p�U�*�{y����:�N��ģv��%�ՙ�	'�Tv��n<v.���a(5T�"�*�WF+n�4��SvS���d���Vj'b,�fD���5�W)5W���yU���h2�Q!-Cr�D.�6�R�-(1m�GF�[sJ�ʈ��чR)b�d$�8u�z��݅���ZKl� ���*$�!�F�4�
dwY2��^1�B���I"yz�Ybr��;FIj��*�,ML�T��M�{p�]�ܬ��q�ȻP�n	n��r3Dm7(�բf�{Tt������J��!ۗj8bխ��uk*Z��\�q
D:Bobh���2�n)��U`�t�46{��,��T����w. l�mm'��A��A��BU�1:كK�4M�P�r��1����fneR1�{���x���\���2��9t�
ܷE����{b�umm\{t�U�m]QŌ,[6�M�����Fj9[4�o�ݚ���F@j��$i���Z�N���a����S؍�����G6�'L��D�)Ǝzk�8a��W`(4�=NPH�~����W�$��!�[�vӉ�["�ڳ���mc�mmL���H��nJ35
Ů72�Z�r�bs��Z*�*���"dd&cY��L
��76���'$�dJK���u"�1�h\�I�ݽ��4��ݘ�[xj�&3��Kmx�54+sf�,��2���U���̨\97u��җ�GV�t&O��E�+s gi����%�����X5���k&�0Ab��&�F�DQ�۬&������X�u�Z�a��ΎS�K�i�{[(��SB�*B���v�e=ɪޢn��dJ��Q�2�m��hǕ4*n霣�&R�ɲ�M���f�֭�䣍�C�2��cQ�fH�G�Ө�75f�Pk����g��ޤ­��h�kC��^kW��h�ԫc�b&E��52LnP�)��i�Ҫ'`�t�63^b��Ƿ�,��e�f�1���[!��eѬGthK.�'	�_I�	���Z�bT�2���6��o(a�q��ٸse�Z��'-L�fF,�$�z >�(�����kEnƬ(����7J�+��/R6�I����R�����j��,�p���譽�hk%������n<XU��XķtٙoCDʔ��9%��Y�P�f5��
ssYU��2�wu2�v�s��1L,�O2-�*�J�a��+B�B�u��YZ���N^�;��@���"�*V�{�tṊ,+n�,:�+�F�nƨÙ��2C�҇/&�T�n����[�#�ok�W�J��7,��,��A��$���I��L� �&���d6)U�����
�Q�v��A>�"vBw0Ԥ>�o1����N�)�3y�2M�ݩU����T�m���-Q��7�I�kv���=Hx�h�1���,�mT�QyL�k�R��X��fc6S�y�N�;�>D怭�x�±mX�d�&� YGlbՉ�s*�� �� �6X�uS3�5y��34Y��^ش3L�%�@�ƬRQU�7G�ڵx2k���hQ��ӛq��N�^���ōH�f���M+�:6b�so&��0d���%K�ӣe�b�3�d^`h�:GQUw��Z����A�u�ŘpMH��s��*R��f�b�f*͙7Ş꽕�J�\�H��ń�UZ�Z��Ԓ��K���ۇ�Y��x+-�!8�N���H�j㠌rr�p�gTP)TZ}0m�H�V�w%:�u��$�t-�lbB+ӯf�X�D���y��[c�El�6�H�����YBL��K�$k�f\��s{&�X5�ыU������ Ҷ`��f^ۻ'[�8�n;��/p�tAaVJ����sCbm��0kI�^�E��Wsmًfѱ��
aP��@T�Mf���"�BӇ1a����-yq^m^�a�+wd�Z��r\�M�����ٔ���/5��K���K�I�54��������[��*�H�L� �x�/��.�II`F����-��hl�;TVM�*�P���j��M�z��u�&��N�IqN�,���uNR�0��̪���;wR\ܭ���8WȘf�b�*�p���N��ւ/X,��nӬVu�,�kn�L��o�頬V�Z��ݨvn�*���!2�?�뿳l$&�k�8��AR�=u�bI]~���g.��ظ�0un)��ss_һ76]n���C�
����oY�}-��)��z�1 \ޠ4��Hm����8AE�x	<H
�<�F����V�#u�*�9��/2���+�ӒLݚ�oJ�q� r	W������K�[M�� �����ĝImaW[I�k,��e)In!vuᱵ�ʃ�Xw���J��'hkL-{��Mi�Fa�N�Jٹ�����c��R�L�li���s`�ݨA�\�9�V�jL��2�1$�Լ["ݒ�xhǟ]�����V�}z�l����v�
k�녳ri^���97-���:B�.�<h�H�Z���:x e�,*�X
 7P�H� �\8�3��3upU*�����f�nM���$�O��EM^Zۡwד,�"�j(��`V�^ax�T����@p�����g�S�~�<:t^3�Y*]��B��9�B��	u����%�5,	,���W���ƣ)-na�+�ɼ��
q�"l�Q�,V@@Ԃ��#�tr<Jt���0� � �j���ƪ�PӶB���]_7F��W40N!Y����{���@j�rM�A��Y��*H��c�w4�kUir�rE�]�^mv�F��(�ŋ�Ь�SD�:�<��M�OhC0n*io�^SFnѭ4F�{� smj��a+/r�m�ֲe����Ҙ1d׻����
tuĪ�qP,	i(�E�n5r_Շ԰̂M��W����ʲU+��u�:7*ԋ\[��Һ�젅�oh-��O ]����^���O��rA'�[� Z�h �1�V���b�WhuPl�Wm�Ř˪VUc��a���ժ��R򥶺��l�u����m�j���l�WePklp:��P�)W�E�T�j��٩H�mڮKRڄ��N�Yg��Z���T\u��J��8�m*�"��u�H픶ګ`�;<��Utm�6�ʵUl��T�*��m����{n�y���!N��S�+��P����T�G=0�ױL��>�/������9.6'�ؚؒ7��w�nnO�vz�V�r8��r�a�Os;v9�^����D͚w��]�ە*s��:ks1�������Y�rC��l�`�8H�/y���t�4Mo>������Ol�f��Rf�v�Om���f�v���l���M�*(R����=���є���ư�iwh6�WO�� ���g�x~�3�|>�6��mr�ӧp[Kێl	��y�:�}g���{]�n�r�Ѭ�;���l���\'��i��E��]�zN��=f�t�f�'��S����67q�9�9+��A�T�suZ.�x1��N�3;���	ys��/n�1u�ۏU�d�A�D:�5�lqām�:I�IS.����Q�[N�Z���K�Mi鸭nv����&���:7í[.	�oW��vR��:9�\��gu�|�1-q vw
v9�YƮ���q���==.����SU�t7g���W1�^.���z.G=���N]v^X�`!��<�g�j��Jul�q��q /�nn��d��NL�)�n۷;q�a���z�[c��`��s�eWzkք]ә�cz��.M���}هI�p��l1��۬���H�{uufL�[ʭ�y�5��s�OC�e�3����&(�b�m��s�������surO��`Q�j7��{�ku&�O@Z����kS��òa��N�N�;�랱h��qvs��;��1bZ�4p�.c�G��F�\�/OQ���r���vt��k�L�"֩a'9U�6:�ul7V.zB��.`�ڹ��0��a�]��Ʃ�z������9��Mq�/G��q�e�!���.woI�O�^�rf3�m�&:a�Ts���B�.\�r���ͻe�\�$��FϴC,�;�!Np����N6]��x<�7���C�q��L�s��Kt0�k����'>�;�ӫ�d���
�"su��v�/#�yt6"�۲�;�/'Wg��_��tJ�k���@�CW�eܳ���$��l�^�47�7f�9�m�ۛv�;=��]�A�U�5�7:�6�>fۉ�nj%ش�F��Y�y��eԚ�y	&��j�<J5�K�f�Ůۜ]<����X��h�k�]���k��-d�Ģ��c]�"B�����:�h�����ƪrsŷ����^��W:���,�	� �v�n�kln|���+��,=�8�ob�1�ܤ�M]�����d��t��C�6��:�k�iN<��S�����6$�+!�c;�tFz^����nƞy㦎;,jv4�K�V:,]y����n�7`}<'>-�:�&��w��vl=BC��b�w�jf�:9��p!�r\m�b�{k����z{.�6�]��X +�آO�����c&|X����7żb�����q�r��K 5��8�znݠ��IQ9��n�Zg�:wM�v�.�çW9`*j�9C���m#تW�{�<���m�4rrr[]];��sp\��:4��nxշg�y��e���s��^�p��;Fu�Fz�:�7���96]�u��&�/G=ury�3���>.<�Ľn�nx�Qz>��Nk�.����`�cF��+�Wd��.p(bt��g.��IМ��:�Y{����&i�¬�k<>�{Yx�3�R�h�;�&�V��+1wm�=W0��9�
s�F=m���4@i�<���=��\g�����k��ۜ���@��p���Д����P�����s%�ۖ�42E5�⃞�sAcug�l�!�O�nݓq�7#��]�7l�>�ݪ��[���I6�{x�귍ۣnzڰt�����bz���K�-�Kk��j��:������R��b��f���P�]Ӯ'/C����lpR���c�j�g3����"��'���E��nz뗢6��#c��8�|b'o�{�W�꫱�I�[ۅ%��<�zp+c����w�L]��`wnL������ms���y���S������1�d��<��ۍ�=�=Y��[��Z�x�ݸ8eҜqذ�����@hr�BL���&5qm�eq�wa����9�`�t�E�pr<;'<>����݈�l�����Ӣ�i�Մ+z��l�z�8�痳Ȋ���>�R;�n�'wg��x�0�A�ƳC� T�8��D����q;EqGe���3�p�Qan�\-��hQ3�K+u{=�Kܝ��Yp�����s�'72�
�uj�-�$D0
�AA��EGh�'$B�kiiӈ��{@��V<��s�L��t��oOh9�Ю�iq[n.p��vh��Ç���b+ ��t[:�zCa�͞[�ͪw&N+����8�
�"WF%���3SSbwۃ�۩��Z�dS�'k���.�8�CǊ�wY7��}�Ӷ���q�|�F��5ά���`>ݎ㓻Q�`��Y�Й��s�b�؎f�Q8
}�r��"�娹���\O�"3:]7������-�ŮY�]�5��C�tu�e�G�qkq�f�b�!�u��c�� ���ďm��ޮW�k@��-=���������7k��)���h=�֎G{YkssV6X;9���3�5��y��W���/-T�s�-[`����'��>��]`��I;��N������Ô���N��qpn:ZI�p[s!�a�ZZ�^X�	�V�н�(z���
����wDَ��ۧ�������ػ�q>��2aݳ�5ӝ���p���w�m��خhy���!m�:���[øۉ����k������f]d���I��nr�˶'O���G��z��%�ٴ�Ǘcs̶h⺝��4�C�컍��r��Y0�6���^W���n0����ө�q���nܾ�q���6���t\N���oj���x�fu'I:|�t���n7!tte8ۮ����Yܜ<��4컒R�ۦ�'���oM��X��7/m�p�O-�<�y8g�N��E�26H��n���ָ!ۚ�����yڝ×l�΀�nnU�;g�D������+Eܙ�����2E�
�z��ݡp�3������yN��s�u�g�� �8�������Cƕ��u�ã&��n��u���u+��^��Y��va�Wrc����I1ZD�Px�u�ug�-<�e��C�p��{=��Yô�	2��x���mڟb=���� �n͸�6���}�Z�S�W��I�n�qȽ:Ĺ���s�v'�g !�9��G[�jt<�gv�{kqÎ�΍F��ⶹ��@��zyw1�ɋ1si�>cv��˜z藬7;���zON���K��g[���s�u��/4�rl���sW-Ź�<��]���9Y��4����q��[�����z�zw�vc�kD�^�ׅY�m��t[č�.{w;�8N6[�$ng+�d|���躬�[��bu͍��ܭGb�sx�u�Dfx�n�/ͨ�)��d)!:�Y�sx�[ֲ��.gKG%R������(��Ź�Uz�^�g[����[j��\W6�9ܻ����A��	�8�]�2];j����p_y���]5	<\�ѵ����e��1��I:L75X=�)�'O�ݜ���>9̛���nz.�C�����1�L�o8���'[p�k]T[�u�V��jj�h�x\��a�Wn�ti��L0O=4[�"�F�k��S��s�0�e��=��A�1�:�˻suv�|F��I���( �9�;�88s�]��<۟i�p t��М��q�<�f�v��n[���g�];�U�6���zZ�ӧ�;�۱�Hވ��&�="a�3�\���	8�2&*������y�猇k��W�<�Ʒ5K-���+�8w��5�;��8��7U(��:t^�W$��9�]��J����3|�^��3n7.�:�����E�{w����%���x�Q�t�ںz��;6�����7�^�9�-М��%άE�Us��g̓ù;Ge6O}���G\�b5�<��D�ֳ�5�:cz;^ۦ7�.�x�q<R���ok�K�c�]���dzz���z:�v��뮦y�����<؆��R��g]7GF�0�&�ӞN�f�2^�muZ��Ixݤa���V�-����$�[�n�޹%���YP��x�F/}'��l�+�ͤ�<�=<���˘42�=��:��n�V&A{��x��e�J;�=�n{�}o7^8���g�A���ډ	���mj��G��7+v�`�n�Wn�P�ܣ��G9�����k/��I^�8[kk��\��X�I�9.�<���r��w�i����	��d)�v6z9w=�^���P6��*��v�#�y�P<��+x�&��v�C��ptu�"=�B㤎%��wG<�M�z�~9/��t[6�c�W�z�Kb^��'[�ج@��=r	��ۨ'��wk\u��0/*�3��Q'���j���^%{4q�Γky�Fݢ$3/3WY�Wn.u�C��=۟Jm��<���I'�����]]e���Oe�:�'>��;��5'-����9yv��t&w�W	x�su�;@�Zp&�aĸގ��eA�,��b��㭻l��]�ӵ�yա����$�Q\J�yi��j�9��y��s��ϏNM�O�d��*��'����Xl=�y���m�z	zu�b��P�Ig����]�ۣv�'9��"x y|��z�+�p<����MǱsI���3�m��l�'i��KYR�c�7��̐oH���7�N�R]����Y�v[WYn(���x�z�N�p�L�x �6;>Ӧ����w{�9����9�ps���pp 9�p�s��s�{�~�����i�V�#dgU*�Nֺ[X��V�L���T�%�]/*�V���3ݗ�:۞7�x��ĻmthxY1=Z�X��A�Z�Ѹ������
U���ݦs� �������%]���\3��7��yC�tp�ze�zdeNy�&�k��4a��5�ŝ�P�����7(O40[�5yP�r��7]v��{�Cs�s]m�G�EFxsض�]%�I�\�zz�vcu��)���8��K˫��Ϟ� �=���Z,c�+�v�y�ۧ^ݥ����8�츻'Z=y�<t�r�B������M�nv��x� �˥�/�l��F;m��D�mRNC'Gg�d����i���]��we�vx�;vfE+͇p�#���r8z�b��۶���Bzq�g�ۦ�#u�����%�݁���+#n%�د;q�.����F�(�w�p=Dc��۳�B:93ض�vi<�r���6}ik����[O�Ⱥ^��vŮ�t�ez��۹��\뜽]w;��ѹƇ�v�98.'�y��g��Qk;�n�q\n�m^G����C�g��LDv:��:�����d.��SV\B/7\`���	l���7m�\�w
�L��U���GNq��:T�i&�#��ܹ�/��U\����>��t\.`���3�a��v؛:���v��n�g��U�`��gO�ܧe��q��隰{s])����M��Sb�/q�޽Q��������cpBX��{rٻ��m�r����!�)qm׈�����t��I�BU��û�p�q��.zU���g�֓j�p����Q���v⣵�8���p��E�<��C�fMڣ����3[����Gk�y�+�f�ns�3��+:�q^����P)�i@u��e����nL�nV��_�=��7*=��\۰bt�:��QP4c����vn8����u\ژ瘻����9�0���v^z��nz@"{�v�mp����D� ps���3���@���{����{��Տ���M.�g�v1���0\�-�Y�:L�
Nv�:�\�m����wX�2ir��u�3�����o��{InG�����^�y��/�s�6c�I���-ȧ\�:�p��:�R�z���XQ�j��L����am���&�ktt�lW��݊��ポ�h�k��(a:�v<�l�=p���7Fi�Dg���{{��n0��瑸��<$��)�a��<7��`��Q �������VW�N§���y������O�Kh9J�7��k��]@�u�HҞ�򧹕�չ9��[��/,-41�FRN%q�a�=�|��k.�;f�h�s�4<&M2_��u�XX������g��{&��X�Jd;O��ݫ�]gS)�)D�����=n5�����nI7��!��r�ś���i�g�����,��E�x,�2����b�P�[�	 _���{ ��	g�r?gS�Mz'��;W�"���_v���_1Jw��n�Y|8�gkwht�Pk}�R~(���PI ��E���j$��xE���껍�3��������%�@��r��И邱[�~���n^$�ׁ������
vA��)R��Y��o�y�=fv^d���	rg�����]y��l�۫�*���W����~��׽��J�+Pq�Z���X�քB�y��ӭ�.[3و��"S~-�Itg�)�R���
���aRޞ�8;]�AA��W�.���^ ��w��2�/f�X�k�L~��� ��^��-G@3��ܲ��g�86��v�%+��p�2�(����tg�nR��t{{�x;Tw�HQ�w8�^�7��{O���.Ü�[瞡�.�8��A �[
�L*��G����I�ή��a#W�Z1��d)WV�0�~݈<��a~ݞ�j�_���!��ed,� ��r+��FX�pC8�h`~'>�o<��kƙ�/��|���Y�n���2��`q}��~c&�^�H�~�$�C�v�jȠ�Z(��RR�Jv`������r�����׾&��L	v�"��.�+�$��8ⰹ���	��j�x+�ǿ��y5�q�73�Nj��ݸ����s[��<T���ۗ��4��Em�Mn-�r���۹��2쪗�0�]�o��m�n$�v��9R�6����ٞ���L�r���{�v���h7�࢕��(�I ��T˒T��"�ｅ���k��Z^�R��Ʉ�I��,k�]a�@��P���&m�mlr�ʾ,�=���0G@i0S�)����~�w䮱Q�����o���I�]�먾*���	QX�~�p/ ��x��+�9�JX�z�ɒ߼�у�=�R�f���H-�^��2�Ͻ�\7��m��0���9g;So\��<=N����tQ) [:x�\�o����?wۜ��:č�+�r����LW2��2+���)A�Y��D��ț;�,{-�!��(٢�����\����[�Wx6�A��M��y��~�cm�q7��nmNע>X�!ݲ׽��x�����~��߹��~Mȳ���w^���Z@pk����܏u0&�[�a�6�Ծ����ț�D��k��x�u�3�,%��|����;s�΢^����n���^9
��{����m�CZ���M��M
k�5�W�V@���e�} ����5���Wm˞n����D�9���0j���p\���/u��D�� 	�)2�c�MW�y������G�i�3��4x���=<;�_��+���f�Tqy���@Jd��D*,�^���@�VC҅�t�w �qY�w:�ln���	4��R�O���w �]to����Ӎ�P�u�=��J4
�3<=�yT�&s�@V��IjP�K��w[�Y�N�1�d��Vv��ft�3;`�x���6v�/3��]0�(�U��U�㘋��n��*+�k5q�-�����̼ܵ|#+�o��H%�7�1�f����M����,*����HJ�]#����m��a��k����-ѨhJ���fw/�nsv�;�v�Oz�<2�YKI!����+}]Ey�&+�3aJ��@�]��^rq�� л*�r���ɐ����m)��'$n���왡.���k��|�:��O{A�����ǟ��I�kdo��9��ܤb��# �t�A��/�ͧ�R1'^�ȅ	��zJڱ�:�{��W���:}�a�	q�2�Kץ�����6��Di&U$�4�hdƸ����ye����&8�;�����Ӡ;�v(��xPDa��T0�}��k%ݙ��
�L�Y�J�m�wʹ?M�@��B��Ek���<�(��m`���{8<����*�>f�"��W�Q@Ǻ���������iЎQ�d��ޅF[�u���|�|�ky[��,��p0+\���p\{!��N�S�����0���K�sjEh��D�i:m2�%�u��0!�KɳQE�;c��t�򋽌��E���Wch�gkmZ�BV:�j=�}[<{.���\]ps����d秱p>��c��1�M��;p[��a�;=��E����G7=��-9��,]7��ߚ�ﵵtpu���Z�����O\�::5N�*��E��l�]�\j�Rsv��[Y���Xuu�;Y�u͎
=�g��g��n:��o��7�{S^� Z�l�O�'�972�iR�[n�n�`���r=--N߇���㌔��wE�����vw���"�v��yn�r�5��m��Y��v|�م��52f���rެ�|s0�"N�i�.�y#��r$�#��-=��>��"�ۊ?G*mùw��e�W9$(-�IY$�6b7�׀��9�kk��c�ِ�D�7B�x�o:[���9㯦�$��XL���YЉ"����E ����1`�vTc:��s�r]x�������ދ��δ+��ټ^�d�x�ly�ի'��mb!��QF�NE��%^�m��L�.��[��2��/u��Å�4�{7�vط���������L����A�-��Y�%�p�0:�.�&�9([��Nyܛ���l�R�,8Z�N�+�f��YY:A~51;�g�Z>fĮ�O�ZЩ[��_�+E�m/4��je"+�fM�.�E0�U� 4��z:if�^�=��Mu���X�2�3om���q�fnDD��Xn�
�S�d�/��:�V^�D����zb��ce9Z+FM[�Mk;6�Ȭ,뵊Ӻv�tBׇ3�Ȁ<����v&48`ַJ�-jv
�4Y�6��.��
m��j��/s��ۖg� ��أ��P�y��k�9v5^r��\�d�w/[
�p�n��7Ve�-P,ذQ�]	�[If3�@s�̭"y������8R�A��Oz��;�(竵OIε���-{9�ȵ��w?��4�A���U6y\G]�|E(�`n��+��Ly]�.�ď%텞!m�s\�� ��܈QK/�ߟ��\�j�7d�����u>=�\2��Du��A���.����T7:ʶ��r����1r]��^��3Ҹ�q��>��O���ӵG��;��,wmtc��utEM��tAt��iS�I[�WX�~�����ӵk��s'LZ��7������wy�l�a���� �_{�5-��Ͷ|�u������$)��-#{��[굎H߲�N��K��Y3r��hܼpI�:H5z�0veF�˧k@pxz�8>���E��vf*��e��l̺`�M������8^%o�+W׎qf��v�=���__�c��G@�B��Rue"v\4Jݾ(�����F�/L:�v�k�M�����g|L�
�rz�ܝ�g�P��.� �=3�9���`:N�$��f&.F=d���N\�gy�E�vɗ�g���[�a�����ˁ��c�����SP���>�Wz�]!Dq��Sr5u�^5������w:��T@�E=f�թuًGf�4m��_h���ደ�,��P{B~:��ėп3��v��,E��ͽ0c��	���x�8�f�r�g���%�0M�z`E���u�!%�j 7�J�u����ݴ��E�p=y�R�Y���(�]"�x����[��s����EoWb��/��{ �w��^=
��b�(wqz3+˝�����<�h��T
W��/n�
S�J��=�vǷ/�/wE�j��bV�!�>�\��U
��;lu��s��+�F��䳆�M�if��9L�Պu�cZ5#(�H�֖�F�qT�O5t���9�Ż�d�4vl��:�je�����雷����aƁ�$	%eH1	<p�j<����׌� }C���N�pa���������N�JwC2���Em���A�]>�����*uF���D��L3�K�G';��l�*�pv6�k��l��=k�����i�a�8����Ud�q��U�]�4�sX�>��~Kv�cў�T5�]��6��A�	Sa�ۓ̠��Γ�ႎ1�uzǛ�����lN�vv���h���&�+��Y]3y���Z��s��gh]��w�{�Q#C�H��	3�Ea�+ݖ�鏣��w���e��m��L�����
���<Ӷ=I������ٍ��+��� �N�M��|�ɳƪx��w�V����L�Wx{]��/��������Ðfݰ��.��&vx�0�7w���.�#A� �3(]�]?}�^v�m;�g�^���#�j��^���m��
9Yv����ng�V���x���xhk\�q�7�zP�C�
_k���tz��GZa
�v�hѷ��P��Y��'��v�;ɳ��$`���r-��?c��.wW����-sֱ��	�ؙO.V��ٓ�Vܝ�f�9����2��]!7����n���=��|�����j`�u�e���P��s6���[����`��IkQ�B�=�C���f���DW8�ے�{�]ك��s��%��_7[��6k�kP{h�B���l��l��B��kq�-lݝ$�2�SsI�2	��kh�6�����O���-�v��q�����x�����vy�xg���6nM��͕zMj�ӢT�	8��$��hw��_��1�C���V�,��x�ڸ:."�[t��z�;`*l~�Ʊ�9��17���� �Q��{�t"�	�4/et��^���}�y)nk��J�2Y33z�/���盩/ŋ)ɵ5u�h_o{�da�W��R����*Ƃ�CjRNBԁ�{�haf)��}��,����^�
�qLu�D���(޻��oy^����݃Q|={ގ�+�������I�E
�5��@-
8ί�SC�W��$Q��\_�sl�����?�����Y�I�ɞ�����ܚ.;*�W�-��h0Kf��[m���/'����n�"�f�o�ɿW1��{�v`�.�? ��W���Mc&�<D����oF9��m��]�$͠xX�#e(��i���g��5�{U�ǫ��\�0eWV�u��BU�H�!0�4��y�:���x �j0�Z�KG�G�9;���;9�{3rY�T-&�>���m[!�Im����q+u��.K��O�v�r��~��f-8%f!��(�S��s��5�s�ӝ�(��J�־&�]����*�Y��;9�i������$L:�����˻�1�Z���{���wu���
���F � � U� ��V`��f*��ͭ����C�!�%���r�v:��z䭳���1�^�%�����J����6�h�e���r��y�yD���u�y�.�	�=}�����zwT������Q��gV�<ד'�'��ƶ�d���.�i�("���o�m�з|�����5B�S3�x�8��:�0��7�7u��9,T�Z�M.ͺ="�jX��Ǽ�R0b!�91��lw\�ny]�:�w&su�p���8��g��QTR�@��
��)��zA�g�ף�ײGt��I��xx�E�4��Ni^��Y�M=�v�msq�wu���_!�"}"<PI5$��K�����w�"�K_����?.�yd]j(���{�����mY�JdW���&����dvvĳ�a �H1"P4���;�;�.-9�͑u�g�i���֏�b5g�C�ذ�)�j�����֭���U�: E��m����
��Ov�2������ ������z�,��T�����<��ٌ��2�x�hP���L�~"�$E��#L۷�;��l�ѦĹ�;+�R��;{�*���C)�zJ�.��v���YR�>[�㒉�9��;*���y����k0�3�OoA��k��:V�j��ʕ��2������x.�����[Ȁ�0�I��1
&�7�u����mE]�:�v���Y.7���͛������"�V�Ph祟�e]��!���f01�����k2��~��%<ĺ3͗S�s0��&����y�m�Y�^�}3���Z�g.��v�^�
/'�Հ����q��-wq��J�u��=e0=��C|�={�3V�:�f:�M��zot�aU��7ow���l۬���%\�w��e�M96���I��w��h�z�rhݻ�b7ӄ.��'�Ƚ��+��١`'�������$B^є��)ō#4v�_�#�m	1u̧Y��b�s�l��ٹ;��72=�[{B�#����ԧ9Va�m���5}cL�M4�d��:-�����/��p=��s' ���a�BVޙYИ��5��s0)U�.�N͚-,NiV����271�n�wZ�)��#�|�e�^WU�M��b�fkb8"؅������.b%�YR���ԭ�Va��d����.�I �ܡ�����wA%����|zF �@~��<G��]#M�:p�<���З�� Y��<ͽQ�<K=�@�Qr&D�X"�\��O��;�!���@�/��z͎�ΐ�r��j �<�ߕpU�yV�(��t����uΝԎDy"��DQ;K{�~�;�EF��΂Z_0�L��EG��ٝ�Zβ�)�ɂG$94��͙�h�d,�_��r�&����	�/���G����F���@C���� H^TE遐{�f�Eg�3� �呾��4#B<��<] 3ō�yD?�e��v��V�u+I�@(�`'mI*��"g�^���<
�[��M���y�y��ܖ);j��f�q���fM,
:t�n��^}%pt���v�g���Ⱦ����Y�"���!G�a��oO߻��y�&�����u��BH��#�%7�;Z����0�>=��m'��˅�I8�pa�FC�]<���}�z�
��)v1��A��!]��Q�b�}������Q�
<R����_\��4l�@����e{>�,3�<
�̚������Y��خ�4��H�:Ta2�h�"p_�ӤC��z��!�:�~5�#H&��.QZ��|����f0��h�Ւ��GV��z�*��_zMCϋ�<�0�����66(�@�Qn�<&a̣��ɦ��.8"p�y����o��t#�x�W�w�!��,�����r�Ϥ�i416�,���#�����h���<�����~�*�@�2�WB�-�v���J믩��غkYz����6uA��Y�Ӷ�oMŰ���(Z���&���=�B<��4A<�Z��!�=*"x�ٵ�p����*"�E����̫R<���O=J�ϔ�ȣ�W�,�U.}�(�(a��R��ф��8;�`�×hA��K�T#��D��$����x��+<�g����Oz��{I�t7����~n���;��[l�plJ�N<л���lỳt�Ӵ9���-���GIp�L���==�կ�D�%��8E{Ϙy��pC���呂��͜�,�~���ψ�9~߻`m�ߺ�-D����o���yS��+��j!��F����Fgs~�cc�6�3�W;�a���C i�{(��zH"�Ӟ�y��ydK~��ݟ,���ژ��X��B�g�P����il��&�Y���[�=Ha��AC��0ת�t���:ׇ��t�Y��9!�8D�(�Q���D���}���ӧ1Yx:�':�Y�����"}��G�y�������꾋<��7�����@���~�K!p�(����0.a��S�x!�HO�g�\4�)�05��[v�v5��ܑD<���l�����!��9!�><#��5����Hg���`|��Α��|��0���뼘ه���>���~8y�bPOP�7���Q�8�l(L$������jj�`3�|�j�6�B�����}��0��}�M��w}�{�y�L|�>"��V�T�ŧ��7ٱ�:�ʕ\}���ӆ�"����6~4������ׇ;� ��a�^�IT���['֌�190bʅ�=*��L�C[
���Q�b�9�m/�Ɨ�ۣ2�
����,�BI&�d3L��+xp3�����`��\��ݳs��{JC���<)��=rK���ۻ�nv�{S��k�r���T�ɧ��;5�:Գ�{��<���L�n�m�=��sd[xݎv��-8g�Ì�#ɞk���c=�M�]^:wݨ�<��1r��ѻq���r�.�m������J��2����)�a���&,�oX�5���;�\����3��"<l�
X]rp\p�(� =l//�v��%�{<Mr��{���{�tw��>��<S�4��.C�+�B��]�i��3�Z���DQ�g��,�jYT��˲"��>�h�t﯁�Y͞��*��y�� |UuvY�d����Fq,�<((i�L���Q�<��xO��N�}�6p{������=v�ָ++g>Y�F�M�6l�]�����7� :@u��C�Ri�6���ֽhi_-<���G�x+.�+.�ו���W4�w���jaڈ8�T��㎀�]�����8�0Ѳ��Η�}%QG��'�x>���2�|���^|��߲hS#\7}���T��eou���s˄�yF�?�e}�|#M���K��O'��|~S���A�N|�/3���,�F��<b�����f��;O�H���"�v������,�޼1c�j���׏ޢb?�s>`a��Z./&;��y�'o��B��iφ!��Y�D
>}ߴ��%��78��8,��<��]w_*$B0��ϩ3�U�uWF������LC~?.�]���w��#O>��{� \��+����6{]��@f�x���^
����1��G�DL6xO¦���ѷ�q�F��j��<4� ��T�kh��<v]+�y@zus�Z�Mf���7$�8,���q*�K �	��҇��O)�G���(������<�Џ����j�@>��Ī�;ëliɎ�i<�"|Yi
0G�G�k<l�'j��$;e{���8L`��t8y�l�����o�����I\�����{ɞ���1�����oq��YX��!y���K�V;t�;�Z���6S���ٳFRn����΂nf��E6Nn�1�6�FF�F���װ�x'�0�Eg�⼻t=���<E����/�q�����7H$�O���/�t�D��pZ����!�����8�л����RlRL�jI/�O=�.��	��Tz��l��|غL\Ͻ���t_~��w�y�\�so��Y��XsG��ܨ> ���w�=��U!��T|�H�ʈ��=����� K��"�>��7����xX1�i7r+�G�><]Pٲ�,Y���g��aΎ��|�}�(B<t锾!
 2ȇ�AX�u�!Ǥ
<(���]��*�@\�~��8��5Ϸ3�̾�O�������>��~#��Z>�5�U��!�z��Љ���/�O:C=<�G���㮿eoΆ��(���=w�!�l�s��o=�}��_��x�xO��/
#)V.<��ԣ����п!��x� �3�Ŋ<V���˯��뭦�9�HJ�6݅�j�Aۛ����Vϭ�ݬQ�ݺ��$�7	�]�5kZ8Zr94}�z��
"3Ϛ^��[��%pa	f]r���#�zУʧ�*���8(�N@�E5���_�yQ�UmOYS�����y�|]���]e���h��<x\���6h�/�Gq�eH������$�=$�h�ԫP 2��{���<+j��h�xM5����*
x�x�!0.��αd|yd���u��<�"�ϧ�PG��uY ���o�����l��ǟG���V7�7���EN9#ѧ��(�����ayYY��>Z�v�Nb�c��ߛ�0�y�U�w�#ʋ�oG���W�t�"��<+�"z��͆��nm()4P�k^�-xQ�V�e������q��G���R������>,�Y����+˧�� 3�?"�=_fZ�>:p���HC���>���8�ᐃQ���ur��G���[�z��pt��#����|oT���W�>���:�>�5��@��. ��\��D<g���K��҈�[;iiܼ�!�O���bn0�4C�;x� i��.Qv�h�ABp�%�
����ߵ�"���՛=�+�����ǚn�����C�I�y��+��|�ҍ��R�K��4�W�T������BK6@7W�@��^��t��� �Ow�e/�4;谺m��(-OOfd���s�j�Lu�z�AŔ	,�Aa�+�(k]��-�sΪ��~�~�OV�rwJ�pc'�3�y�߹�8}_us�Z<��W��L�.*B�8GK��Ҩ�[�E�J�yDiD|y���<D��d�0!ҏz��r����t�3�H�&!n�Y����M��k��H!x�����_ #�/�޶��dt�3������w��<��!�j�}��*�(Q��>AZ��|F�3�ud߾�BYH3� ���f�;�x�Di���^yD��Ze8��ă�uqgX��p�Wۮ�0�j�F>Ϯ���&�B_����K�㇊���Ǯ�'�,�?j�G����*����yG�ma��۳��4~=<-�Cͯ����^d0������䎸,��:�}va����ਬ��pb���-_B��Is"�H�}�s���Αڼ�\�j�"����|*��3�VK垝<��
�c����^R`����"����u+��v\�x�7PR�o%X�P������H:��J�S��aV��D!w���q��g'e�-��~��f:�a>�O��Q�}&0ņ�qˍF[�Wb�^zzG�\zG���oo�\x�M�0�E��4Ն��D�b�O0�Hg�>��x�Péa�KS�P�p��Ͼ���,���L�t���K�ԉ<��>A%�de?���%�Mq1�6D���v�쀜�<��g/ i��^�Cu��rl�6�����8����3F͟V��<���W:Fl����] ��U���4�e��CO�4dy��D�#y�i�vq��I �9k��se4Fx���.��(�p�n6�R*y�t�@�՜#L6G�w��e*��9���.�U�}� �4��p�p���>��9�H|1s|�x7��+����B<�"K���.i~����j*>>���4�٫ %6�p&Ji�_=!��!a� 	�J2������(��=�Q�ˊ�6{��/oƅ,\k�4|;�/J/�Ş�> Uc�^�{�|���zz!��Z����ӳ�����w~|G��p3����to����iK)F��_gV�🍓ﳾ�|�xO�Su�1_��Cǋ
d3f��!���tMV��#�<���#�Q^B��R�f<��f�ր8~=�
���M�{1pN�a��Èi$]/H�/F>�d	�(��IM'r*��1(y�Q�"����ߕ��7(� e��hwP�����3>Ci�Ҹ�.��!�8����_a�d2%"@�!$����(��0���#�D.	K��!�)�������O��(:[��1r��mnNF�1��O:�-��4J{cB���I��a�+�¡7�^sJ���[�Sތ��/	+�-�R��N'!h�L�,m{ȣF�s�.直n�.�uÈ�n��������A�2�]���Oq��Wmu���y`-�/�v�xW���j��z����8�=�tuW��@���"�q¼���<sί7c��'[���8��WC\�)��s��]�g]v�\UJ�$q�����$��@vM�����ur煶�.x}F�[H�n�]F5�i��[g3'[7m��nݗ�]nQ-].Q�r��ۛ#��lf��x�E��u�h.�[��������Y�!�,�������}k��pTB�/�)\�d��<ߊyD@�9�����m�j~������4��_=��y��"x�h�]��iD��:b!���"�8Z�G|y� C��H#gH�ϔ�g�G����ë�X+����I�#�ܺ5��Y������|��i�a��yWt�q��`>��� ���� N\d`�����\�t��g��Yxo��=E�!&HT)��G*(�z-�������P٣���x;a�maן*�����"��9��5��#N���S7q�t>�
<��鸑���{�+�zx7��!�ȇ��z���ą��8�q��柍����<~��w��$S��|�Y���X��N}���4��k�Rϝ"x�,�VyG��F_ٟ}%�~>#��u�X�;(���N0��V��6y�>��͵̦���O+f_}��!�*D�r>�i,�y�K�
#�@����C���Y�<�>���3�g�����Y>�J��5����g��o�n��C8C"YU<���yg��|.x����������w�~���mIG�^��F�.ݎ��ܜ�`)��\z1˙�UZZ{rnb)��x��3�D��=��p��}z����tu�Q�Wq�xM��+֫��!�#�B�,��Ɛ��٭����}y�M���O}��!鲍]_uW!xs�N
<��KǤ����p"(��05$���u���<Fa���[�B�,�2]��D��XF���i٣bc��f5�-#34e�@eT�*9��p���-:���p��1(�bU/�봳�k�<���D#͞���_K��!�r�<~y���Oĥ�@�}�Z�hQ5Ƿw�,}h|t��\�w�{���0U���ǃ�����ښ�2[M��B<�b���:A�4�!Di�Ͼ��_:@��M �z.|ϝB����.+: ��Y1�!C�P�.���\6@�L��i:���2��pi�a��'��g>�x=��K����S��!�:l�z}������[�n��ӧoo�����P�y)Oj�h:x��r�w# Q�X�#��,��pۯ� M� 3���d�������������_z�a��J���mx��W�_&5
&ܑP�k��C�x�_�Xt�E�����ࣦ��Q?�w�{�T��@��`��0��jЦ�,��O*�t�Q�yv���<��J�ߕ�ڌi���]ASB��=}�K�vn���5DN ��tܼ)�q"+�,�qy�V��LZM���Vu[�j��{<^�F�f/������83�.K깟M�\Z�8��\��J�$�0}v�<���	�Z�b���P�K/�����"l���8E�ԍM�C��H��b� ���rP?.��h�ɂFԒ�g,�p�y�����~��΀&��aV�Le:x-����7�� �}��ņ�~b��⍞i_���GM�!��T�Qy!��_ێ���אt����;��H��%�`x���E���"BM��8p�0�*N��)w*��Zb���T i��G�e�d[}��w__=�
8E>�u��~�sL��γ]l-U���[׷�|�z�Y�Sfn�N�I�6�!�g�0M/B��:k�e]�J&�{���r�QDN�}(i� Y���(� �x=��Ƃ>#�A�=Z�h}rf���QА� )��q�>(��{������d.�;y���U`F�4��:�s�:GZ�<T�D3��+�C)X�`"���f����~�\����W�@)�Giu�MO�4�!�� |����\����!~"��:V�|����)p��H��H'�C<�!��S��n��{�Ϣ�/f��T�>����l>�5��k��=��=��G��h�U�|�#� �fF��Υ���0����,�У����<k����x,�)����%����%���s���mW+ʻ�n΂�ٜ���g���L�m~�=�<��kĞaΔ,��<t����"��O��BW?�u�g��}w���?T�l��?���[�'������>��~ Y��J?�d�϶X���3f���j��Xdÿ]"��4cSr�7�g�G����D�,�_��0����SG�;⍻�H�g� Ct�﫲�I#�$@�TB!
A�Z�b�<���%�<��N�,@XyD{�gM
��C<�߾?n�y�|0��<�n2~&�D��[rE} Bڻ��'� �]]<��;k�{��>�� w�m��<&|�es�nk����F�o��m�3ψ=D��̽�@}k�\����t��o.iD	��t.�P,<f�ԃ�.z�����e��nӉ�����HC��!�e�7HG���<n���C�C���OZ�_���_�uT }��WM�X�Y/��b����`<�z@�AJ�[=��^��t�6�#�i�;Q'AD�WUq�>����|�����\�8�=4r���vw�<fl��E?�T���)��M^�p��ٮQ�]��������|F��!gH���4X,'!��+��<�|Ő0٭��&����F�,�~C�DY�~@���n��9U�\x�h��wuw�Z$_{ܔ�x����񇧟���,a��������Q���*��Q�����y�e4�@A��QHB ��lt��N���v1�ڍ��K�sΚ���t(�su���va��#�3�G�ǝK]�U�-
�"͟uf�'�w��g���B��2͟(�k���k=s���?Ȫ_yd��k��)~46�0�Q�f��.֜�G��a���d6����t�e�	��!�.�k�����=�k2Jlgz��!�{<gH��Ww�ڢ�E�
+�x�����{Z"z|㔀���(�:�_��D��F
�o�����E{�g��`�F�=��Y	�1LiI,�up�mp]#��	����^}�� 4�B���|؇|kt�N
K{�_Ն�� )��<�\6����$@,�`?�(��'��#���{�T@��qx��A��l��k7q�[��#%ډ9%��#���!3��/��C�7���4y�/�6oɐ����0!�E��ϖ��J1 �~��H�] Q��b5/~����C�WH	h�K*wҤ�Gǘ�6Wz��4�Q��\�����G��S�A�ʒ�y�
<�.h7�g֬o�<R�d=ϟ~��۶��W��\<��W�Y��u ���] ��O�ka"�ݞ���^'�|��,<��<}�}��x8����|r����7�{Yw2l]��Ղ�Llf��vU%�Ɨj�μޔ��.�d?o\1*8��ك�-'�n69�R1{/7	j�7�ֶFWq��Ź�W�Y8��+��[�엶�Ztz�q��ʑ����p��E#�^X��~x�`m�l�����)�c��2�X��&��v}r�s�~��]"7i7+�8�6j�ޜ��:�V�e�fep���Qz_o .�{.D>��o������}�02���k���n��v�� �_N��^$�^�7/z�;�B��lGm�����g4v#�Kq�U ����l��)���w�a�؄[7�_qA@�dU͟�X�2����zk2���BUfC鲅�e�z�z����D�2]ެ��"�3^�U�;��؅�t�kaR
�O0V.�h��*�_^��v�{:�U����Ј�GWc�;�v�m�X�3K:���8b7����m�nn�7otM�8hV�1��KΒ�x˖�����y�uY���/?��^�ow3�_�V��6�t��o�[���n��!E,�e�-��y���j9�Dn��rC�a�K�����=�p�u��@>��G[>�
����@V�Ä��nf󑃏����!-�l�7oUu�d0�g;/�u��"L�H�s��X��i(�Qp����%��M�2@�\{�ſYu�/ B���y�d� �?.��� ��5��E6oF��g�2<�N˱�P�D��G{f��H$����,�^鵲=9��Y(�H����]�t��k*�d�b�1�[%5;J�S�[���m���/q�.c=WsˋX�k���!�����#m+�vy����*�ʻwj猶v�l�PH�Zݛ�:�z�vp1hgX5��Y
����GG;-��`ٛ�ڻa��⅞nL+%�T�Pnq����?gxkY�wQ��u��<Ɍ'��K�Zkj�������A-gO%��5An�6��@��v�u���M�z��i-���+����_vV�(��gx�.0u�8���q��q�y�ƞ���iv#�q�w:{	����t�<�'v��;�n�ܹ�{e�G��jN��=��g��½�;m�-�ؗU�#����'�dܚ��Kv�Rl�<l�u�	v��!��i�/N���k�N�Iw��<cA�q��fLP�G�"��mb`�2'<\���ݶy�ln�浃��'<!-s�k�&͸�S�n��s�pr�xT��}>�63Yʘ����Ev�ٟh��>����˨����	뷂�,�05��nI�[Qpܺ�SYd��ɀ9ꄦ�sמ��g�������g���,���ɽ. ��,�D�ݬS��d�l� cOg۝=��kuWog��(�,��Wa������n1�6�8q��S]�qظѭ�����tpA�X�g��dwNY�Z�o*��=r�7�ٴ���xL���+t�P���ħm�R�,!��Njwn�eٚ��������\a]���kû�w�J$a	^��[`݃>u'����0�H|��Ŧ�%A푬70o���8�۶�]4\f�]M�loB�q�i����Xk�s��lv��GM�x�]V��Q ��Ǒ��s�ݹ�twp>��U��p/t{v<z��WJ��z�� fQ����YK������v���Tz��ųX���u�n�j���+a��{u��k#�?_}���R�����m����nx�d���7gq���!y��������㷮��vs�pp:꫎b���cu�[��嵳b&�lݓ]$�s==��N0�����n'E.���t>�֢�mm�S����z��C)<�7�R4q�m��ӆ�w^�^x��U�V��̣&n����L�';��'R���yqͷM-�ܷn%���nIxf�y!��ʤv��,��99��K�K��m�Z��e�qL��!���<�rWe��L�6.zlgƗ\��:F�U�ǬX�8��vx`�An��\��:]���nI���m���n[��n���WN�6�w_��xW������ Q�W��,����@$2]}�säY��R��h�}�f��8���|~�ͻO��.�G�|p�yDx�- ���w>W<Y��g1<�;�}�Z��]
ez��9#��%t�o}�i�iv�Hd�'k=J���Dc�~�B����0�!��3Ƭ�L�_��C+�N�G���>�Ϋ��3�upY��	�4y��1��S�&����WU�syd.�|����	w���A	�b&�RJy�s�F�>"��H�V������o�Q�Q �!|)����P��YM^}u�O�w�ysu;��[�@Cx��o�`n ,���6��A|���.Y�}w�MQ�I4�j��0��di�;�:k�_e�C�"w��#�[�C�>��fń}�z�;��AdCg���Z�"��}�u�#1qaߐ@/��/iB<V7�Hj����OH����"�$��"����L{e�H�CrK��S��]*�#ƏN�@�E�+^o��GH�\���Q�� ��w�3������{��[���>x1���CĜܟ_� ��G��|G�?y��͞E��@�bx!�y	0�.�o|j��~��X1��Fy8m��xY ����<�vT뇎vM��:���'f�k��,:��u�g��㿇=�Q�i|C"x�>�CHg�U�q��:��Cӎ�<�>5��a�B;�Q���z�t ���/O>';eg�{�d��D�+>w��4�e.Q��\����|��m�BF�NGZE��`"���A!���'~��oZ�{kO	}�9�g��y�O���d�.���M�s�4!�ci<*T�c/����crT[w���j����;�Z�T3w�jy�s:��Ǔ��f��.����J�~�MDȭ���I=\dC���G������:<��<y�
�;HϷ�`�$�A�M=�d�5b:JVm�T�������T)-	��n2���g���x!��>�&L���pY#L<��օ�Yk����X��+��(���0|~�-�x�ӥ���C�K+��|��?N�Df�3�.���㇟b�Q�r�4xOr��$�1m�#�J�H�͖�8:{�����=�}�w::	��}��g�yE��<>��@�B�ᯪ��8��e!�Z�(����n{�<�b��e����}A}���uд��_�`C3f�4�_|z�,N��ӎ��iQ���B�����p��C��uO!Ħ�B��W�E�!��:Q��X<U^�P:x=!���:Ff}�$�E-"�\���:�jDZB�<"�����fu�~�D�&�m3s��.���]�����&�6=>�۴%Xl�۵�2�#I8	r/Q�"ȣ��4��}]��t��C�ߩ�Q쓈U�ʨ�msH�A�C�Z�g��K|s}u�u_��x�� L6@��Da����Bΐ�G�T�Z�<M2�,�{�BK��A ��E"�YGH�� 2!g
~��]�4���:��t���<bc�Y�Ĉ����p-@gUG}�A��j�fKTR�4P)x0!�a�"���8���������N�I-w�"�dx�5>̺���D��-ǽ�LBR� ��	Q��7��Ҁç|�D�<h����>[���Şu����9#���Re�Õ��l��m��üU�A���u����)
����ʚ�2V]"�#�0�=��!�{��gu`�dCr��н��A��^t�}��W�p����cڐ#��!���EB!���ʅ�a�	�sq}HU����0�M��$�sON�y�7[c7���@8�!�,ɗ�"������
6A�Ͼw���1��6y�XD"�!���4H�ϾVG��WW(���B?��c~%�=�GO3����1,"��8���>����B�	@�!�r*G%F"B�������hg����8G��,�!��<����)g�߅*�������}�C:�k�D����U����k�~�>"�$
3>��&�#O�|�4�AG��D�Ng�j��D
��$��z�w�����U�����ܕ�=p�g��ՠαSʳF����?}�=����	�O!����^!d�������#�At��G�y����;��C<��y�6��c��vP$!����>U2)3�;D|L�>(�)q4G�R^y:�#��Gm#G�zEy
�����ؤ���#�KӇ����a�6}^`6�7s�v�@�;]��]�TYϚ�t�@��|{��C�t��Ӑ�aD_E0O�<<{>�@�\�(���5�����2P��#A��1��=�Bc=��#��f�"�=]�F)Da��w:ɳ�GO�:H�w>�P�ň-e��t[�*��|��A�ƭ�U���x4��ǉ�~�`9�zF���Ȳ!�=��{�k�4��1 ����
HY)3�����r<�a{�0�Qz(nt����#�����X�嵥���<H|]!Da���z�M�!�Xg��<҈��=����o�ρ��g֗�������1����ϲ��@�Ro�*��Fpt�'u�ձ�_)�;�wn_t�tVuͥV��7U���f��˔XW�e� =%]t��������<$���o�8.�,a��v�bH{�D��ӄ��VI�D}��$Zd0G���X�m��U�2u
�c�Z��Q;�t$qfa���\=����Ô�%o�t��+L��
$�x����W�U�g�C?!Ⱦ,��p�������o����뎆K�.��]�m�e���!�V�Z8�t!��:���[n�ƞ�f��E��^��|F5�(�H#~��y����qZ�x�)
��'���:呧��a]A�1F�4��o�x�O[�_s�gY�!���Dv �l���]���/��U�$=%��4h�g�u��0�l ��#�8Fŧ��CdYp��D���5_}�\5�+BY;�V���?h�^��}�V���O�pT�V�����ŉ��!�+��R<����(Ë�<�u�������v�4�I.�ֈ�K��X���H���(�?_V� D����G�����:0�e�I�� g[��f��u" #���<F��&���D+�b�ĕ���'>]�	u��xQ���A�={>t,�p�|��l�U�=u�:R摠�� BH��|Y'��	#��>�I5�
�-|�Ax�0�WX�����Q�D|�9S��f��$E�> ����}޺呤Y��\,,G��|�#�o��
b��+oG}�f����K����y��˔Y}��ywd�#GRBS����G|�4�a]���1[�� %m�ϵ��è#�|Y�e<"�0���^��=˺�cGO��y�!�>~`h8t�(���	�_j�L�?A���$@�r�>w	"�x�^��dB(��������R&�tL��P��u]VI!H�@��B�c�)۩Z:$�5v������al���w�31���M]B�s��@�D�l j�e�;v�OnD6Ɩ`q�6�즬vã+\Ls/6�)ѹ"Ɓ�F��pT.I[�Iɺ���t-����8�����y�y��3pdbi��b��Lշ�I;���Ƿ)��ۮ2a�|F����(i��mp'KN�(r���'�ۺ��[.�[C�9��=\6P2�Ҷ]W<x'{\x;jn�;���*/�N�l�.��Rp�/]�h=��P{v��滞bɹ��7KvuK6M���&�y�����~nYa��G�L
HY���v�C:GA� B
PR
��P�g���,������p�z�?j��d�u��Z��~�Ӟ�D�g�/Y刺��#׾�Aμ#�A�`<F#�!�O�k:��i����0���*!E�a;��T�^A�t"��
�P�gH������yR����1�?x~ �v<���2��F�#�c�cO4���Vwθ0�Hg��d<H�y���Bj�z�O<�Y����>o����E���݋BGl��2$�� ��YU�"{4��/��P��(�\�\��	�7J�>��΀����4Q��,������.��N.w۴k�vu���ZxL�H@ǁ�}��C�!�OHK~BRg&�:x4]��D8 .D�2Kq۴��AZ�ZB�߾m��l����CǘE��G���P��d��:��I<1wd�
"�qu$�#��z��������������y��ä�Y��nzP�.��Gǟ}���)��G�FĄH�0�`M�\��"�jȇ�;Q�L4@��G鲆I���g�i�m�yxln�s����@3�ߟ�|L\�P���E�}r�j�zF�g�d�Eb-�f����y���IS���GǄW�GC�-�c����l-�2��ĜY�.m�O3ՙ�툆�*�3cv����ڇ]r\�Xԏ� iD�_x@� ��y&�M
�;����#ǤY�7m��U��[�k�Vϝ>Xy�Y���Q2k�f����#����Yw�)iD�E�GZ�R�%���$$�,yG��x><�0�K��9r*�Ξ�P$�	f3Y��w�-��B�h�7�=��6ܴ��|f}����T\���I՘8�tn�U�����;��.`�5��+(Xꝛo��z�C�خ��;$w��NN�����g�=w�:�Z�O6��e!�Y̶,ѩ�t�O:If�ǔyG��7�ע��hi��8��G6�Ǟ>(�6ye��w���8ۄJ7$Z�:�>(�H�Ev��G��n*�6N!��(�	�C��D�J��>��H�lx�y����B��E�]@B�#���6v֞	kH�h�D��D�#�},9O�y��!�!f�%R��&"|��R�t?b�5�����љd���]d��սt.� �Y&� 0�<d��`� `(Hg�D0�ҍ��#ٞ��7U�x�H��8�٪9��4����Vl�F�&�� ����}�]����P6ą�$��M�>�@��G����dY����}��[\'�"����/}�y��ޑ^��P���@�.v��|��Y<�VXa�Dh�߳�+�N��$ҳ�&��y_^�y��O���X�#�0�6��G1;�����={WTt�A���A������M�s;{u�ʭ]������Yd
�F�˿,!��k��J����%��Z �D�DAD������:f�BMf�)r�t�M9��򱄛+�u��e����h�I�Rާ�C��}��������k��˥���3υ�!���i�xB#Nbm1g��4��c����v�"6��?ut������;���,�[�{��\�h�Qdߠ��d���#���`��.�t�ť�E,�$��]�B��3��jR��ֿ����s]w��|y��D��Z~N8DR&���BKO�b���N��,�t�d�.�aE��,� �W�|Gqa����P�PD�%1��ɿ/cwC������w� 3����d�b�n+8�fL�k�њ߃�.�#��s�T��9(� ��f^����~ ^��0��J�ujDu=�<]�Q���I'�����ad3�G�\�,�$��d)F�+�9��r:�0�&!9Ib�K1f�k�J�2�E�{#��}�C��A����C���#�ċ�_-O��0�I�ǯ�h��+j�
$����Y���Q�ֹi"zZ������o�ZD��/��C�,�A�E�Rw8."	��R�
?HY|(�N��H�Q�A �J@�D�=:A��nS����1��}�G1��;X+���_�����Q�HwL"�$R����UdK�.2�<!��"����=6ԉ���E��W�1+`"is���~��Z?y�'�O�~� ��v.:at���Î�-lp;Qs8l±�z�PD�v��M:9�X@d��<˝#�Oy�#���N[�!�k��g�&�S��ǆ�,�;��U"�0P$���!��F���������t�����ac�R��!8�m�=ߥ���I'��28t�� �<_R��bpĜȯ�A���h#�><f@���*^i� �j�����WH�� ����2u��|CHF=0�����v���$��̑��Z��$��(��͡g����*8	7�)�����F2!=z� _r�.ģQ��b	#��t���(�y�BТ*����Hҍ��QdĈ�ٕ��,�غI��~�gI#.v*@��B��`-5�^�7���8�Ə=��߼�Y����_|�QD���㕙(W��$P+P
 0�������� �Hۆ��p�J!�O݇ު	t������ث�W�1j(x�
�E�	��ϋ8B��9/��O3Bd��WP���3�9�h�l̩w/�#5 �9�	$�Du�{�������#n
Q?@sk�� ����[�x�ͭ\R��yɋZ�+̏DU�R������(�]q�gΗĂHW��E�(��v!�cG�mBJ!R�O�;nh$�L`P"�y��B���A"R���><u��9&W�L�b��"��i�iԆ�gra�����:w��x��<ԍ�gֽ�>4�cR�9<��\OP��`������$.��:��.����/@����_oVtn�A,��v�bv�Nya7]��qէ��sP5���u��I'Y杹뮻F�����;�CԨ�K:|Y��?}�견ظ�$b$*"�.��i#V�g=�����+˂#��&���_fg��7�}�5���D��,��56�<�	f��������!B���HK�{q���BB�i4�rC�<d\\�6E�a�}Tw�z�Y����ߪW����ߔ<��$�Em{%a�0L(����ح�y���߷�c�O/�	*����8��H��� �^�l�`��:xA�b��Fc�}���󧈂��|�!�A���(���w��R �e�O,�W�i�5>��X���~!����R��,�����c�&M ���iJ}ߥ}���r}��t�I#J8�����24o�
(�&*,��}��A�}pW��>���<Px7�-"��rI$���p�:���	<6�<����tx��pv��~V:'O:p��C�!�eZ�j�_Z�{8�|E�tbÇx>߲��i������0�h=�Q}�gԾ�g�１�U]�e�#�(���$������l�(�p"�;I���x��X�$xiG�ʿ�]�Hac5��N��>�}��|>+'�k���c��\��G�� `�7%�'�Q�-��0�y>"|_��^��MҮ&KI ���`�C#;�${t����+��.R��!�呅�kvO��C��|���������.�'>����^�U6��X%�e�~��o��%���8�t]�6鸼<��mĽr�qʛ��gz��ZW�i��g��g����+�ݰ<ܽs���͌ݻ�76�5�{Nu��������b�!��ջ��h��^˻�ź���/3+�Wn���[�q�'&mR�v:���=ur�;�$0ɶ����x
�]i��>8Ʋ��m� �4����mkF�d�%��{U��{n�s���A�4d9�A��n޷n_ N�y7"�\�s3�+�eֈ�p�N)'߄<yY�*��϶�#�~-<d�;��O�h��h��#�4v��0��NMϻ3��y�"�<��Gݴ�e�`ϫ���z��Z����Iz��QD
Y|#�~�VQDi2,�J����,�ǾՏS�N"���p��~�]�i�I昐d�Q����UNs@h��G�V���Ҭ3�7�~�b�T�E�^�*�t->8~�@
�,�b�U���p�~"� �K�
c�韄����z~"���������~�&�]"��8E�,�����0�j38ۓ8<���gH�,�\��2;_w�CI#J%y�a�|�cD|p��p(A�������s��*��pQ �����Xy�#!Q;�p�K$��ȇ���uݛ<X��_���g�C�_����ȃe�Kj9(Y]A�D�"� ������>�;�3�ϝQ��4��[�� �੏��TQ�G��ύ/>�/�6W�|R��D6�0%<�Vt�����Z�f����H�^+އĒGg����A6t�H&�ݚ$�ms������>Z�X� e��*$���/�F�4a�!I�C?{'ƹe �%�
�Z@���<���JS�ނNgْ�d�{�B	t�=6GJ,���?���iZG�"�~���Q����:y�	'p��*�$Q��(����$O���$��$�KtH��M\v�]X�{Sex8��#��`�k�(�Ը�vD� 1�d�Iy�ˋs���j��F�D��^�W,�8�<�A-AEs�Ҳ:x}b���A�B����)h�>0��_ά�!���CY���3����h�����H�ս�b�#�<l� ���@A��b��bQ	���rI$� ^.a��������.#D?n��U��xخFy���<��LeL�������v+j�VlT��~M�-YszklI�ٔ���Ʈ��O7&�j�WWf�����VbA�>�K�~��xKO�^H�I�;���s�7�2�!��2�>+A���u�D�W5"I"��!k��RЅ�]e�����bG�#U�Z�bw���|��.y6,����+o��$HK&&�&H�%�ԾB�A@�jG���E/��X7���I&2�@�/z��zp���p�~+�O'F���\��<t��Y�x\'�2}r�`�b}D��
����U"��<���P�>(�3�u�m"l��P��A=�IR	�9#�d���5i�d��N̋��s�q9��Ȝ��̦>��� ��]��tM4��>8���q4H�4�F�0�K1�{��U�:F�C5�y���a��4��w��������k�����qp3̚�,��y�-	P��@t�!�%�F��@	x�(��z�ޕ�G� �
 z"xNR_o}���{r�x7�bq%i�_!d
�R�عg��Uf�Qi��$�.AA�{�|��R<%}o��s�̤<aҺ���7��@�L�ᄿ�˺��w�G<΂D:�TR�Ղ�Oby��ƃ�i�.�:�6�˛~w~x��|~(JH��hC-i�O����Ԏ�\>8C'�.��pl�24���3��<�$/�sR �i�d�=���ʾ����~�//g~�kF�,�?�4EXN�L�Ά����Fb0�"yQ�$����.�� Q��&�����A �����;���K�L����FsGR#�Y{."�}���oUn�7�B:l��Rd�dQ�L�=��j�4�Y$��<?*,���|�mVBI�CD:_w��n���zx�1����9�,v,�_{�]���� C6@�QD���ϾUz�C͇=0�KH�����ʷ[3�M�����l}��q���W��H#�FJ�Z!Z��4�/�Rt�ۯzE����bR+�63+��ޫ@��yf�LmgJ4����;�=�xB)Ni۔���2��m͕*M�eG�N���@nғk�1�S��%^�{��V1�*��7��d��sm�1"y_@f�Ԏ!Dꙶ^"�+ӱ�z�,��(��
��K`H�e��O0�x�qT��El������{��pL��Y�O[�Ԃ�e�yf*#N���/d��̣�p|e�F��(w�FS x����랏� =���Ȫo��t��q0k*TN0�L~S���,���M[��]g;��U��xK�7r��X��*�e��0K��5��}ږ�O�3�;K�Wo) �}:��V�����nr���
�A�1H����ڥ1B��Z�WW:t�,�L��Hx��C̋6�9�f�
���L�%�r��ҼE{q���d�|�R��S�a�vV+����w�N�u��cGs/�Z��q��ivG\9�WV�cy��(��V^�Ȟ]l'��oygۑ�7�C�(|�NU�h�����;��Ԉ���F�OVd�]]�4�zA���������z�6c>�ߥB�cW�f
�G���f���p45^_�Z�˴����AY�9�Nɠ�,("���	Y�yC���� �6\��^ë6��H��y"���Z^�ql�[
�},w+f��]u�m��-���{I�̀Yy�ӱ;�G��al����t�����y]NոL5���Shi��Ƕ���M�O���f�ѓ\}yWܒ����>F�������U�\���H���"���0����H�<D�����ȻoNi$�=��Ȓ�7)7!��b���y"���SY����N�Ƒ�+V�eه��,�{��Fm�Q��b�2<��*��@��G�1�V@��D��:|h�Zh��;5�A��ͳv���5	����gɗ�8�(�RH�,&an\p��NY������u]��r���;巼�	g:a���~}��q,��V���f6s>�n�$*���Jno����Y^]퓦ЄB�d�i$�.5��@y�zΈ�n�L�[Eq���Ӂs\ncl̘f72E�:x�}���T0���o&�ѳ�v�URN�N�z�ʍ���,gv����Y!�2f��+l�U��L3��
�%/�m Ke�w�M;{x��^VƯ���u[����m�t�ߥ���Σ3�	 �%�~˖���S�T��;�+�����3�s���������^N�(�m�d�����#���~��M�(�������}�'i��h[0wujE�}�<�S���O^:�)O%�[K�����ffc�����Y�6�]>V�� P��)F�|
���=U���W@������|��(y����c��z�W5y���d}ި�&�>#Ht�Wu��[�CI�I^V�He=�d���>ꇲm8��cY��psy.Z�/�����q��sf�'�����ӎ9����_/FY���y�nOJv7�,�	p׎�<*7���O&E��X@Y������4�<6��.F`��)��_v�*�|w1��.�s0���b��cU���lͧ��1G��\l��K��%޹�%b�.�U��a妲ۚ�uԹ!���h��>t-?����/����o���:��L�==��@:���?K�'�C�+���-��n�����jT?��;[n}[�Y�/�Uvt�h�fK0@�&r���<��ܱb�Xhgb�y��r���(q��D�˪�T6-bY�>�㾛ӈ�:�/��,�aϪ]k2�i}�����w�E����!,-�hy(xL2�a���2-��u˴�`Q����`�fxjUޏV����/��V���� �WU�K�O����QK��V�a0P�����}��֏���?�������p�g��j~�w�A�����i.~�uײ��z�`��7�v?{D��4���T˺���ϕ�.50�F�<Fv�����I�<Ƅ���k���%�&�9��U���>�ء-9���>go�7�yؗ��q�k>,|n�T6ER"�w>��|�4qL��M9���7�g�P�lU����:���E�0����6q%�����p{Zc㹚x��A��*��}�����h�Sh�1d�{�{�(kXJ�&�N�@5@�QI�Ϧ�ڲ�N�)/<mL'X��v�LV�+p��v:��mc�"�}��I*5����Y��?'����C˗v�WE�bHoM��mluHS�#�Ε^4�v�f;<�Uiڎ�i�=bz�gv���ͪ��)㠃���u���CGX������R6��=q�N��[�ԯ<^z�ju׎.�ӭ���|��c��@d��gs�����n�l��n�G�����L��x��tn���38��[�� �)o���W0�q�0U���Y�q?Clh�j����vPD(L�Ǽr�y���l�Xy�j_�|�W�%��;�3�'繛�4�i�-2)$�e�'���?�������`��'���w֒��D�_��� �Ey,�do9y!u)b�w�ڼ��ש�Z<o4u.3Y�afH#�Ƣ᱄�x�q�w[�l����@fTv�U��l?�xۜ���]��%��e�N�U����UX��w��5w�g����^m��"�,"�NIx4�0;]Du��9B��V���t&��"���|���.��T�턅���i�>i���Ŕ/������,�][��W�����s@E�-�	1{��RG�{�3�_�r�1���c"��V]��3.8�>��WJǷܲ������^u�^�M�X�D�6�~���Cݳ�H��QQd�,���%�..��ܺ՞�I��Q�rl-��V�u�vZ$Y)��}���V �:T����\o�ef/�W�ثg��OZ3�>���3�_�V���dx	�7��H�\�~��sI���O��l[�T�
ny�$h!lM��7B��BH�����������n,O=׺�U�x��~ɳ^��b���ق�7�qpYw�OL,�s6�=Nu���3�7<+�=xG��2b�e6�����O9C�a�i�,�$P��%P�$+_�.�K��{��Ψ���{��/g��<.�>���oE�ݴqK��M S�I�ݱYs�/1&������:���H���E4�0j���v˞gf�ѿ�,S�s�5-!ݘGgo���n�!<�j��j��o�&Ď�19�1��3��ᣪ3]���g��*��d�Cw��,Xx"Geul�x.��AP�Գ]�#�̾�ȿOA@�� �z/��2L�g34aJ*"x���69��!��;%.����p�^�Aֵbb�?I��!]��W"*�Dþ;�|um.:\gӄ糨1����g��b�s�4�P�@��4�&B��!��l��:mv�v�5��a�p7Gu��n��q6����ϓL0�s�u�/�ڳr[,#D
���O�hWҺ��V[��V�m�8��C�c�=��_�8<s%A�R�d�D���H\N6�0�{k�#����]�/}4P�$����e/2]"�H^�ǥ��.�0r�I�5To�ޮW��^�u����_��m�_%�39Aԇ���G���t�-�
bex>VgT����
D�2[����y�^�5���U;�_-����ˊ�w�.� K��!�>禥ͳx��!��!�@����<��6���b�t7]́-e�nuD_��^�J�Sc8V�3>�f��m����4��kԟ�S=�9{U����e�_13Tf��wo
��O@D�l$�ϑ�^]^c
"��l=X�Om�2������*��S���w����|�@q�(��벩e�v���r�g���)�G{�Ɣ]H��"4d�����ޚF�Ue޳VC!y��W�y���dʵ-�瘼*@�Dc�L�ӱS�+����煩1�+p�H�D��.���^kW�\� ��(�A8A���T�W ў�Ѻqֵ��-�ܶ;V�Pn�6m��Hy8#e(���d{K���=��*�a�D	�=5u��!��yd3|5���ߦ����o���d}������*�Ĵ���!_|
Dӈ��#�U����SQ���ӯwi�ʗ�yuz�F�Z�4�$߼��[")v�dB'��:�D�r尓ŗ�a�Y6Q�����T���5-"$8�0�=�`������q�	�jp��|QZ�G��דw ��4'�eWx���U��~�yxo"D�VS�v�W��jH[P3e62�.���Z�1�5�М�'�������������r�����oR�ٟk�=�+�f���7��k�l[�K�>��я�E��e�ɖ�ք==J]����0E��0U�e
��@okקԬ��srE�=T{V�T��W)7*m�Ux���* ��i�/��Ex�WG�x�����0�a��xn��Ȋ�y�B#��H^����h=<d^q�����W�:B�Ҿɯ0a})� ��	�&Z $�`
�y��Vq=1�����l��ɪK����\���-�Rj�=��7HMC�pSW��U��z��<�Z��v�Ur��~��U.?yF�Z����^�<8�P�G*�5�k��	V(���1ð��(�L��I�]D��A8{U�B�[4_9x�y����^KU��q_d4�#��59����N{�Z���"�砳�t��ni��N�{Uëj�٠�y���u�ED_�N8ۆ@��9w�3�HD�o1�e�a����wX+�/���&.3�0��Ӎr��?v��V�j��폌?i�Y��>����w�d�ZdPN�6����c戚z��γ�>�{S�]��(���]+��%�9`���g�{e�@hq�� b�F�S�j�{2����3���"O}G!�4ڌ������ �"j�]}�t�V�V$�*�5S+���N�
!gϼ�͓�(\���K�����G�D�"�������j_���z��K,_��}3�!A+�C��y�����|���Β\�}ľ%S��I_Dl8�fr�;Fl�M6�m\;E���^th4�W'u�Žؙ$F�Pɒ��)�qb3zJN6tKn�3v�(>[�76��b,�4�AnN������s�ʇmۺ��zR9�E��
��t�������Z+V%zN�=��`�n}&E�k��E���*�S��|�R�<V�[�D�,�3< �s�;;���櫅d�{w�<�M�$�ء�7\���<�dE$<7ոz�}�����t�%�޺�*�G���|sAb����=��^Fc�[x���Z���痸HU�㞠����F$�so�e�Q�����g�c<�ҬVߥd;0�z#!c{��ozQ�;���5J�`Şa�~ې����{�gE��ӄ�bNqf�w�x(��ێ�w�6����'����A��#���
�'8Ow�����7Sc��4�[�#7����d
 ���V� J]�ڿ���#A�A�E L$ٹ�H�QOR��ث�����0Va|bO��x*��[\d�B�eF�NM��N����eeq�����n�A��n��I�v�i���CH�N�!m�q��3��}Ide�]��+.���<�J�����MuJJ����*������y<��//c����&�lvxȕ^�oCI��B��+�S �P�?M��7p������A`)��/#��¦��V�����7S�~d>��#�[2��H&��(ܡ�ô|����<a��ˑ'�B�r�xwIZ�l��nר�e�[s�mY���y�涢4���,�#�M^�ߤ�,�<d.�\L`޼{��竀t��%�Nm)��tIV<�Hh��}(Z?G�ԯq�(��a4�ᄲ� �I��M��ۃl���a�wإ[�ugm���g�)xi�iHsz�s��^�/{��Xl�"��7����,�]�xe*�M��y[t�ɺ����~��_"�oz�����19��7�u�|v�����ؾ��
�3�-��������;X���r�P\��~��ЋpXr���GR�!�yH��iP�ת��=1T.���Fl�5�׆�{�"�MWU�A7�Ϸ}T^Ǖ�>��GWk������Ip���뉧!H�b4�dw�<��^ͷ�5���ޭ_���,���|F�V�͏o6F�@ay=��e��6{�l�n	�T�҅�i�3�O����A��a�`IǂψdtĞ��X��b�31�6�-=~���lM���}���W�^U�x�H����v���ڱ��,!�(�`+�q���p��PzT*8�e�X��љ��֠8Yu��N�X��\��]Zm�6Wc� ٠�e&��·X^���u`��c�݉�C��2�S+׼�����(Y�)U�����ϫ���V}¥9:}w����������
C�����sqDuv�����}��8HC�u�I>�ڱ���i�Mvi^߻&��Mq*�
�~.��$D�P)��v����k�@�ዕ�� �Z&�>�ԅ�\p����$V4S�S<�^"��{Vs���@�XB�w������*�ʗ�ytTQ� r��I�����Ml��	�=��3fn����f�����^��A��6=[�.#�U�s-����br4huy������u���v]X}�m&9	�,֫=*��4��i��S�*�+����5�A�F�O�w|&�s����V<�q����þ�.�g��sG|�ʆ,n�F�=.�^���.r"Cn'W��=8(�d
f
�/W8
0}M�⡘3=�*ڵ��w� �P���(Y��w����S�����=
��MW�hLV)��h���� ��۠	��ȋ�2��Z�_wH��tx�e�^8�x{9�������'�En�n3`��o�8�ݼ�u\=��g�	�	=���n�wؙ��p��������c�qѵ֝mu��]Yŗ����`���ͥ�R� �.� &	t�Lϭ�8�?=J�]�����w|�`]J��ܨ�^nǗ�l���7k�?�U�Jtw�í�� K��ߺ�=�u�7HŴg�R�yz|����u��#DEp��0�^�ym�t�*�������V�f-�,���je`�"���n��*a�����@, ڇ��.Ƥ<=	P�HI��W��
/UA+o�Z5��O%7��p��!%(
=k�qn<����U ��!�鮵|�Z�ֳ�z�ʻ�,1w�3����(����W�u�F�v�S�%>�Y���k.�KjŶ6l�Ń7�f>z��M��Xڗ���＜s��'�s�OʻR��J�I��7N�O!�o����z�������0\JX(�ٸ���e��]��f�\����Y�VE\�gM�,��6�+�D�W��vv�'S��N[�������Z��kO&����	�����x�����2q)�%Z?���J���w��1�Ƭ6{�k�~�!��j�S�g��[���Z�ލ�[Z���F��f�٠n�,�v��Z�]���
b��Bh4ڳf��Q�Տ]炞_n�x+}�ǻ~VPB�5��yS�\�]1(�y�����>����MKǂ��ގ�H��uggN��Fq��2S@�H4ɦ�7�F�M���v3��?%7�Ny�.>P��-�t���Ww���X>�d��ev������s�눙4�\k��2��Tx���Ē�l!i�{��kU�]읭;J�k¤�yۂW޺D+qA�u�m�o۶�xw� <�&{g�yVW[!�;I
�c����W�����U�"�/Q�ix)
N�*7�<���`���r����B��YK��:�gl��R�m��wmz��R��O�EF�p��T���U>����ժ�st�ӵ`]�ix�E��˔�o�u���J�� ��βb2�kJ���²���=,J���Fhj�M���R0��WS���{r��Q�2�K��ebX�t���\Ɩ��>�뮥��e�Yb�6�����h�Px��B�eu�3��ϴ�x�l.�/_=�ro�׷�$-���i|2r��1��8��i;Vh�Z"�ݻWr�|Gt7@�����#YDA Lކ3�p�F��R�b}ŪP5�z���x�Z.�^)rk;����ܓq�r��f�Ms�ܮَv|l�vI���C����h��rr�;]L��j�i��g5Y�+�8���Mɯ�腬幣o	�i��+n����8񧭸"�sF�{}[�v��R[�:�L���.�k)���8̜�Hc���pW�I��uk��Q�3���v�Z�ɇ�V���A��؁��-��c�c�t�<N�ڨ�����]��y[x�&��f�0��=ˣ�QN�Eẽ����1��y�c�v�㛑G�Z���:$�cf�\.�D�����|�+���S;�5���_uAcn�o���F,`1٪L�&�wr���1�Y{�q�.y|��l���8�vuÃ w�S���#�ġj����]>��T2�%��y3MnЭ�en���/A�R°��>*Q7��{�v-��qQ�/KD��q���a�8�֗�e�}�|xV��s�|��v�*�� �d�-B�3҈V�A�G|�j��@\��H�4����mժ4�m�����|���mm��]�[��s���-�O7G%n�E��)K�`�mvly�����J�X����ڹ�w
8��K��t��'=���C�8۝YB�
�j��הu���W�D�9OV���en��[�m�<)\��Z�
��A�vҨp!Q6�{t�B�b<�WO���뮼��`Zǭ�4tv��/K���pn��g��'7c�v�9#�z|t���Wc��擻8���a=�ڧ����փ����Y��<ƺz|��9N�����x�{s�n"t�����G>.8#k��s�]v�b�w�
��h1�7������v�`�<]1wN�ëi2�pc�KWj[��2<<��!z��{򮫺��[���Ťy+��>눥�v�[�����W�.�t��ż�����9�=h��m��>�#��{�:�e]>��M]�"ɤ�j�om�|E�9�m�p*�%X�x�N���5�r��7cD��{���2r��O)����Ⱜ��Gy;s��cz�Ku ��vJ��IwF��\s�Ʊwl�d{u�n·pם����鲯[G;�3{ϧ)l��v�e��l��<�	�y�si���'H&7R^�Y�r�NѤ�uA���ݺv:�ǭ�e�!�b8�v�Y1�$���!ۧ�ˣ��͢��W]�e�l�v��kE�L\�'��:�L����G�v�r�&!{E̶q5�\�v�>AG���Qaøy�6�B��&��e;:�]�'mɋ�᭚���R��Lk�m�g�nÄ*�W7d��k���^�f��=�zY�x���c۶�H�ƥ%�ɹ�(s�Du��j���o6����y�c�B�,7	W<��u3�mm͏Y�<g�i�����vUmp��;��U�y�L�F�q���W9�mv���n����ӹ6ۄ\�t��yŲ�q��D��Us�����yw\=�Y����b��l�vm-E��f���l!��ɍLs����E)^����xRx�[�v��3�>�l��eY�6��JM+�Tkv˩��(�1u�v��	�nL�e�p[n���I���hz��:����wVn:T:�݌�����Mv��O����̱&����i1���ޜUͺ�n���U{=����a
vӶk�ΝܧZ����Y�*�#Gi�v���l���q�t�=qZ|�s`�:�ٻ۟F�[E� �������費3s��q�5f�.H�I��i�s�+�{�2�]h�zɪ�c̠��Q�ܯ�SMb<��[��&\�w���k���غ=st�17�,T����x�u P���T0�^0���*w�2�꺭򝾣�hu�x}��
��>�5I�u�z��������/m�,UM<#�l�Y���Q���G_Q�9"-7	*�NJ˘ly��=y[%��;�=�n{p�Ţ�d�>�h�t�cL�|U�^g�P�V�0�P�ɠ�<���֎ЧE\p�c��Jm�!@�NFJ�1ERt���̝���l�ğZ���e��_q���IA�*��q��Y,�0�w*n���頇.��Ɉ�o���$J��ǌ��	�Kvs2�Vg2��'l��#��lA�6A#�i�Z"�_5�i��@�'�r-�;�vǲ�;-�|��61s�m��Z�)7i������s�E�!�I���vL��ۨu�9�ݛ�:J^��FD\mF$�{�h�^"��;La�N��Vx�u�%��NO�
cy�ڳ����y<	�{h�Z�S�FU�|����Y��¼�|�9�%p4�,��A���/K�a>#���ڂo=��l5����]�zk�.�@kOe�Q�em��;�Cu��f�:�7f\�٣E�Y`��^�*�u�Mj�j�ye�i�v�K�$�7Kc�W|�AP}��ʺ��T�`nػ��C¬w�\2�V�ʙ��(�h=��8E���j�t�x;��i"m�A�b{��8Ex!�ɰP��߮�C�V]��:�ۋ��3s�0�=������A�	8�%����+���<Z�h�E_
�
[θ�^V3}�+-c^����8J�Wt=BQ�6O��,��μ�֩U�e.	+o�;�_�I8�s�B�����,��m����خ����i�BI���]��(<}�� !���-��;A���b�4R�/vj�Et������6��]dbM�F#$�Ɖ��[�<��kM���8�6:vmt�r:�����p�p5 �=#H�Q����w�he*lom]xՊ�w/���@���T��ҕj��CL�w̑i��R����a�Uj�EoV�Q��	��M���)�5��_w��&�G���״��/v�q�0�Fk�,��/>��,AWRU{�ҿM��z�ʞ�A���������&q�z�`&Sh��i�c���@�	��^�+#�C��X��|%;4�#|9c���\�H���5��G$,�Tm��!h�V5��=����|����P�,��"�0C���8T9ƴs�k`�[7�W��}'N�<�����ց<t�gH�,zm1
2����$�\i���u�w�`��/9]�}h<g��澜��7�))�or��}Dr�_W�؛n-��|r�ah�',ū�(��`���
t�MO�l�C��[�2������:��h�W�g�r�nECڑK���u�H(5�^���~��OU����2]!*a�_�D��� 6	{�:���׊vz����M�ӡ�bo2�����n�{5N��.K[T\Y��|����~��3���|�ڃ"�R1��]���\�yU=�q����zf����Ǘ�\�p�.��R{�r�����FmJ>c�H�d�	8��օ��w$�����Sxj�0w]hz�����M�f�W�C�O(�h�^� �"~��L�YbN����7u.(8 �m�	�i�@���:�f���sV��2����=�;k�BVu�߶�[����ދ�o���f�]xU����q@ep4b.H�m)8Ϣ�}�%ּ����֏A}�Y��j���Wxt�]�ٕ��%?E!n獾//-w���g����Z�{@*L5HpGxs`�}|�(���y(�w��;��@j�qV��_Wma�Hu��@o`>�q˪��s��d��c�8�ցM"i�
(�2�V99ՋnN�*š3�́.�(��0���8��T�<?\�y}�S��\tkQѢ�58}뭞U5`�w���VGL4O+A���1��gH&��,�7��ɞ��j��'6ٓ�gK˫�V�V�������ժ��1��;�T�@׶s2��S`��*'����&���o#F�ܽ�X�iKi�a�1�!qR'����R��'�A����ͤ!=bG���n�w�w�S�6Э[����u�a<�1`wky]W���} ���8O3���GZ̢�kG>�P(�@�M�N�I�z_)�� ��EJ�g���Bc�|)��Wg��oȁ{s;o��oN�#�V�B[�v*�t�J�6�k���I�e���Kg��(����x8�w�{�̴7��8BQ�^ώ��'uzۺw[�G�҅�ٟ;7�w�����;�gW
��v$|��*�2�)h��E�A����:b]���W�����,S�T����X�� �׺�ON7�%��>�s���L5�DV��ꓥ��k�����j�}M�`�q�[r��~s�0�$ଣHxmn�.Nڌn��Y�"�G:����-Xv/����]d���:������J�3�p����,��Y��է���qDo#XH���]�qvy��ц�=�����UZgr�Y��j�`���n�'��w/r�p�h��C�\�U�0\8�m�5�<�`ta���	�ӛ���������ݳ�I�Q��M��O=0ޅ)�+�6q�r���<W��:�um%�pڲ��Y\u��k��;n�;�4��471F1�1=��uk,cf湁��⮹��*�x5�q�t�C�f^��n�	����D�������N%#RC��J9���A��07��銷38M����@���b�l�e�;�S�V�/|��>T;�X�@g!�x�"v�V����1�\�臈w�a�(ѽ���=��ew�+�����A#�ޏ,S����g����Eg�u��vg�¢�5E'G�
 \��:��l�	�.C�z�M�Fkb6�ͮ����(0x1�2w=4�v�ED��3/p�l�Q�R)���0'rz�=�Ӷ3$�@]%z/:Cl�l��M_w���9);����ҷ}�Yr6�^%Y�whc�_��`��o���ly�]�n���w�ُ}F^�7�ˡ�Qة	]�xc�" ��	� ���
Ơ����myպs�ffOjd�A��e�\]/Ew����^�f��x%�y��!^���RZմ�c�^G� T�]�*#pjs8���CF*u�Z�[O;��z�N2Z䐲%NB�,$�NA��EЊ��P:a�E]��fCLUp��R�y�n<(�P$�kg	n��)�2�`�� ���e-쿡��Vꏥl��ȸ�������I�xH�A!6�oj��6��A+U�W���R�cs���Wk��6���xF�n�����H�f石A�x%<++�s�S�w����D�J�}' �4m�X�+��*��ʔ�#��`Y(w=t�)��B��E����#��)���¢SX����G����n���[R�w�J�)��Oop���GoT:�!��b׹Trs�� U!�/���M�L��i�X-�*��+N财�Ȋ��tj�-�
x�)AU1̝��,
/�7M%ǯ��ȿ0nˎ�M8�=`)����	�:d�08���T�QV=��
,�W�e]؉{+v�@Z���N�O�q��[99veR+�bQ��u�R�9�`�]�=�~�؀���PV�ŗ���K�H�g��Z7h�ݞ�e�
k�������O9�'�ɜU����ջU�Ɠl�������ߚ=�SW�B�"�vp/V�>�������qΛ��>����t�~���{��A��������ab���qƂ�A�[ML�U����.��e�����m�����i.���yf�g�ו�Y�eN���̠Ѷ�{҅�,<�{��[�����ޏ1~,+m�d�' t�	����[���Շ�)V5��!3r���_m��
L��{.��so�NA��Ԋٴ7=���b�]�;Tcy�9�;Mm��u�v�g�M�|�Z�=����\$RB]�|2�*�1DW[��*�7�&Y*�� ���
,}n��&��ߗ7jKP	њ��记Q�jh��*$�޼����B����[���z�./mߨ�so�F3�šB1!"@��^.�!�VFs�L����.{t�6�j{�/"��T�	��k}OL��%��
��P�	�����i(�w�QXA#�*�d:9���Q����(t��岧�c.�ʃGNM̹�N�D�D��2J|����ߥ9����^o9��,b�Iw�=��2��f�>��W���f�AV*(�nNef��^ZrǽWc�^��pn��q�����m�3�e2�9�W��ĳ(�,𭖽���oz��K85�W�o9��t�HCP>�W�0u��(�c�zp�ӓ}^�K��AT:��Εl �I��A��4�{�y�;�X���S�y%
c{����T���2���^�uo�]z��,4�J���˫H�����	��h�F����a R��q�늰KrY���^���N�0��#/���*3�q���͊��Qh�����;Z��'Y˗���GM��*\��ju�!|�z� }nZZC�:�������#�5�Y�6e�Mo��z\4�."�v%��'�p�}�*�t)4Q�-Ѥ�2�L����y��j������mt2{C���[��)��IQ>���������s�.��oC���#��ߞ���{�z���2���\d�ȣa�'0�:�c8����=\�[��s��AF8��0����'�z�,^[��4�)����8�CV >v����ϓ��JΖ��{gR����K0[Mwn�{��朞�t��2(�Ĥ�fm� y)�ON������w.���ꝛk|���-p3��ܷ�9�S_� ���$��*�h"�N�ح7�7�a��`�ٗ�qI�_/�������N��@�M�|^�^��82F킺���=�uw��<�;<�3<�#�	��Cͧ�I6��'�4ʅ�Ju�<r�����,���M��9|������v���m��@p���X5��z��z)���<��Bb��>�]�&�N�&)lf[�+�v��}���7��p�����)mL�O��挭��h����Aw�A-�����МU2�v�L8���bAE��cclZ]�y�%�f	PИ�cw
+a�1!�ğHh�EjQ;�}iZ���[ү�켮֞�Oxf���S���s��6G���ݕ=�^�]m������G�n�G�OZ�c����������sk�n��<��h��Q�z����GQc�5���+s ��ܭ	X�q	��-�oi9��C��GR�d����`s�!�#�b�.�d���݇�]h�,l�%�`�y�Ζ^����\�t��^����)X[�pǷ#�mru�k<��i䜽,��7]�:øw���� *�s�9뫺��[�t�:↞�L�qD�M�L����RLsgY����D[h%�w{6����	ݱ6y����7������Y�؆���綁�b����nt�ys5@I&�-�CЊ�M	o�ו�b�nsK�ԖwЄV�3��R���:Z��+|}�BW�/��u�=9��|=˲W�=���B���*�C��@b0FӅ&�9Y'��Rj�د���y.ܙ�ٵ�	�s�����@�^�����;��-m]��͝�� �mz��\��''A�")�5M~��z&X�=�T�^
���ՙ�z���{Ύ_����������7�hns�5zh��[���{ֶ��s�#2T��Y{w偕 �B��p5$,�G6̞u~V���}Cr7���Roc��zX��O�j?>u�?V$y�
����z��;M1��߷���u>Vw�c���Pmy6�\&`�.{'�vؚ�-X�H����s��xm�:���j�������믑�޻��I�Ż?����~�<G,P!5K�����-
�r��� �R��j�S�X�X4(�@�32�Z�+�:��u䜴��'}^ϥ��[H�b�HU*���K�k+���MJ������T-�()�����w%c���:�ɿ1�=ޝ���˫X��7t��/�Uhf���ۯu?=����X��R��x�NJ��N�nd�o�HxU���%�e��i�w��Ghj۝.�<���˧�nv1*�o��M�uמ���$�=4�ڔ��,'>~7]��%�R�d5�_, ��I*�*��*�\�*�um�j���ى�z
r�3+i���6[��I���,��(�m�w�/�Tq��.���@Y��$�����̬�߄��T+�L�Oe]���k�2�O�@��{�(��>�zKy�yƽ�+�0|��l����2�4y�BJ-�� ��E�5�!ёl�)��Wf���;�^]jMU6���A$�4��ˆ9:K����3M+6H�u�O�e
c-	��?7�0g����{�n�ʾ, EN�֩6�:�1�ifc�K�����4���� �]<��i�[�Oc�����M�r�;�����z�\ˀ}�Zt�_���v�z��z�gvz"��V�5��3{P��" E�Zn�}���*�%:~���N�m̩���Y��+���c9�P�v���6�E)�9��ai<5uYM�z�pJ��K[\�3GU�"��[��$�G��H�0;�#U����bU���"���rl��� �.6�xw�O?{+ʸr�� ��y8��i �e"q�2WCbX�"���[:�)�4�ؑ�]��,�0iL\D}CFA�W�f��ZJ9ko-M��0�#������^�O{r֛3�V�E�G*E$�!J�"�0?On�sʼka�g#�i^.�Sf�� �ձ�xtШ*�d�s{LT�+M�����c�ߍ�GE>�k�[�V���[�t�n���rN��V�����e�B��C#!����6�[��m]�'�������
�1W=�B wEd�>�86���UwC�-�m���Lr��K�/eּ�\w���Æ�v*�ܽB���lS��M��]�>�v4�:�U��2���*n�GQ�,fc{���_om�1z]{��ɫ�C+�j��aNV(k�4A�0=�2�&jx'z4m��pʉ�lF��R��#c�|T��{sb�e�7w��n`Ų6�ʛĮ��Z�n�*�jT�Y�b���j>��e��u7_�C���=[�v�aTj�g&X���31&�2���Yh�k����T��mhU0ݮ��%��S��YZ�w@�]�۽��8�{zżYϗZ���
��Wf�pU��ܾȦ��.���K�QJ�jT�z��˩��fe��syT�>�!]B��������)Yʾ�ׯE�Ľѵ��\��׀�Ԧl-� �h���$��~4�#%z�U�ևF�4�wz�Gq|so.�MHj�Fi~,�I4�*�-���AjX�3�P�W�����3D!_O<��|Dq���f���UA�캗X���=쨬�S�z΁��-�|}}��KA�@����fr�^��͝��ꎷfG�39���V�UX���o�a9�K�	��i�^[p�~�z�o�E�ݾ�y�Y�BLDA8���+h�gSFG�ܶ;�]β&��sv�=�Mb� ��IrD�F8����D��K�@�A�<|4�_}bͦ�G0�PU׉�q���z�P�q����/{F����s�]��śFYg��5�p��\I��p������y{k��/���Ny��X7��_����%��]lF���(z��ٝ�uO��m�	�"J�c��$��t�I�fX����.�i��0z��[	�[	��9=�r���y^��|�o0�S��]\־w��)�1�3w%�}�(ja�I	)Ȩ�ؿ,p]�齉�pO�(���w��@E�:��9]<B��Ζt��y�:<HsE�Y�
�_��q�nm��B���'�����`������m�f��2/�8���2���?M�����fť��]�~}\ N��f�ESI��n�ۤ���T/�OE��7�#����կJf∩k�~�ԈA�4{���r߈�c|��<���B��]���ɨx�p'	�.q��$s�;7�6�� �Wg��y۲�,;q&e�n�\ʧM$�t�uͬ��g���K���(�_B��ɥ�]����V�����wuw\������pq�Z* mه���vwe�ES`�@��`Zі�Z,K�7��]����7������V\ߔs3(C��z�m����=�{^�f�,d���Qâ���&��d��eKYH��ܝIn���o#%N�7�}~|���z����=��tU��幸�Q���Z*��s��}��9�*��Q
r����JD�E0lؙA%K}�ߵX����ۧ�(a�=��|�57
�.{�8+�qP��ݧ{ �K�皁D�IZ����z��
q�)"���U�����k�n�"�0�w��~�Ii��[4.7YSFeY/���]����}F~癊}`�ƹ���^��X���&�T~f海)��iF���[b�9�!B�"o��z]F��1�;��];�+`4[޻�=ܺ�@��f�fp�z���Ս��$Yr?�٫D�p�z�nK���qƱjF&M]��{V�qc]�zwG�l���z5J�϶SK�T�h��̓/��,�u�t����s,�����f��	�*H8��y�s�#�9�a��aalɸ�v�g���켆0�d���fr���N�w(�]�@!g���ZM��o\2s�m��X9���Q� ��z��g1��E���6ɹ�݆�n;�X&�E�[�u�NF]��]�nx�+c����!`�C\C��`>�M�;�_"��̓�}8{��9¯�kݷ�ۭ��[�P��z�-��Ն�!��?k�� 0�e5{��w9��t�_��PCާ�����
�'�7��32��l�^���u��N�E��q��J`��uo:od���<�]H�M�Sf�A&Sy3)�+'�oq���;�k&P�h���hn�X�&zB�գMo�X��x`'�Vu��"k	c&�Jc�����7�	�T�UJ�C{�fk��#sĘ�����k���ݞzL^ɻ��oo�a�HX��A�N�Gh�z�r��Yc����{G��*�*j��|�p��D�Jsg�3�*�]=�~{Z*r8<�7Y��%���P����TE��d�n�u�k��7s�b��9����/b�aq����؝�-"W�H���H�În�X��S>m�Z{=v�[sG8�3ɡ���g��I"ZZ逋b{��w��w��s[2�����ܛ����O-�ᚺ%x_(��炍��6�W�=����������y(�!�d&h��I���n23#����C�����I�-")���װY�!yL
���:]`A��9�#M>�5�]8lu�7RV�2���Z�,��s[�{��e!�<<���!�v���պ�4�����`{�]{�=�Qw#�黯VV�>^;N��u�!!�J9qXz�g�5���K�h�qg�_\y�3����}� �u߯K�W��η,^�鉒�Nr�tZiҦ��Ƿ��b_����%�J/.hW�vЉ���w��� ^j}�<.�n�K��n�j��wxu^�#�c��Q�F��(Y+�
��������Z�[�Uڢ��pZ:Ɨ@�=g0@����ې9�d��0��%O��;[�gsi,��y��<����x�i��Nf!{r�/n������&����R�gn��v�f�?��w�I�G�����^5Yt�Qܜ#V�j�y�Etzр�[fy�N�r�)�=m���U�h��� �̗�M��bK���RP�n��R�:m���Li��ؔ� ��)vw�u�^hovz����^Q3rƼ�dx�ׅB�14�G��E��l�CD���(x�z�^�Cf�]{�C������t�|��5ϥ^n�S �3�e��#�4�^kq�0�T�+�D�u\ױl�K��aa�<�7Z�lO�BN�p~�d����y����^d�	�Iܜ{6�w3RU��4Tj0Aly�Ʒk�.�D�ټ3��8�x�s��PYi�j�e����ϵ�F�<9�D����7�L�{{���KԤf�>ٞ쀾�4Pj�E��>��7�q|����NxB=wҥ���F<��>w� ��e��^�|�_]5׋9y|�����0{ضX��γ����Xǯ��{�f��p$ ��{/f�q��X�� �4���֦����m��⭷3���V���	@���o��|���c_g{8z��[׸C�Y�/���ey��03���=>�<����ï��Jt�D:l�ٝ۰V��ý�;>�^5»W���D��Ƶ�3s�8H]��TR�{�f�uj#�ײn{�l�!�A��w-+i�ӈ7N3!
4TQC=[�)���)�wJ"V�~����7�W���2��/Zםϸw��
�]%q�/J���=kc���3��}.��>��m��	��b2߰s��,+��*���{��V-�؁l��Rv]�HֽG��X*�(m}S��U�jU��kث��O��V�q��� �hvx꧖9�G׬��u��8�4�D8!�k���^�g�O%�)7Y���W����q��r ���	��EJ
��O9����e0k��������tfVK��^G�F�b쓯��;�Wt�Y����ۄ2i�M~JTs]�$=�fy�L�#r����۵�g�VWj�͉ܔ(��"�JE�{z�f����<d5�ߎ�������j�.f��7fh���Nː�D�Xc�Kt8�s��9B���~����N��6�D̴Hl-Bƾ\�y��mcm���)�&�=y��n�u�{ǔ0}����U�gx����r����9�;��{�M��`��m��+Il>V������;��AA:Q��I�������
�P��+�|ؾJ�ݟ��r��K^'�E	
)���a#���i�0��>U��?���AR�wf�S(-��c����4�(��:�/We���w���^�w&쎜=�PM�A�tSc�2�i��㐯��ޞ�>�,x��p�׎Iޅ��Y�2�^��}�:�jV������6��5��U��g�ܿ5�N��w8K��M�"��ul��cz'|)��\m[�,c���V4�Wz�fQ'�=�u"�'�a����ŪIp�
�̲	HRE+����n��Y택��VoY6.M5�U3��ù��A�p�ֶ.����m�E�]��M�u�>�M����8nD8���F��Y���NF�X�m=���J�en��t�3!�ډ�۟q�|mZ[�̡���A��Z-Of��t�ʉn�c��琎��Wf���x͡��xۮ��j�5��YN�aj���\@0�j�������̈�s��k�[���rh89��6���ZL�q:�rq]
�6[�?���w��|�hgn�]^�?J�Jⷭ�m�ܿm�RX����(!�!@yO_�{ޭu�11}uv)2��[��l�C�4I�G��x�G��}JwWw���9�f�����߽�md��n��n�ҫ�<Ȕ9W��8>�~���^ynP����P���#/ώ���w�C;*]݆��}�v��ݕ����a#G��iv��XSv��/���N��=�m��B-]+�2<�)"R�S�9΍c{��f+[��$�ml�x�h�%.��2^*�<��E5b���Sf�tȂ�h��yv[��Q�n����Q�a�Q�n�fْ��s��N䗊k�,��i�=�k;7��f1G�.J��G<��.];���k;!öao�i�nHz��RT�0�H-��pݍ��q%�w&`�{y��M�W-��zzt�an!|AUg�IQ%#���n�c���"��t�y���g�W�;�pdgQ��e7/|��2g��F�<�kz�l��tM6 �o����Ks�{'1��Ѩ��϶7�w�f-��Û�v峳2s���.���n�e�����6����̎���:��M��|��O6x� �u����VYo��n�h�g�γ�N@C}ݎpf��U֬����������k(#Xt���M��>�&+%2��x��֗|o2�����/w�"ٚ(g���~�{�.�t,'��v&�-�$�h��d̤CR Qi�
i���@ڝ)��e��o?`��B�(��/�vC,h�QM�{�6o�Qor�x���������`e�^}�[o{���5˂��ݍ�J�JūE	+ H}nn=�{ӕ�����U-�S[ޝ1p�ҵk�p���y�����������w�?�e�Y�Z�q�ok�N��"҈�$���k$�l��ŗ>��<^�uao7P[�F-i����|��iQ�I�E3�cc�"]�8���dR}#5˷�p�r�V���^���ij��=�j�o��j�v�"�����ZV6j�a�a��]cL>�8�'51k�!#�S�~�\u��]tE��}��r��^�{&[>ďG�oTXi��*����5fo�
!f����C�H%z0�Oz�����M7�2�]�|&C�y}]�嘅nwb�ѵ�[O�"��m�0���cC�/n�ST72�8��n�-G�#�F<N�C;��TG���o�t�g}vB���Һ��	7	w��.�(9z�Ŕ��|�B��doO�Շ�8�ja�!Qh&�J�p��&�Ҭ�A��(��^�<}�e��Zĭ�6�w���,<��KnTә¼}-�W�3��4��,�~єB�E�l���:N���9��S�:��e���G��']+�`����B�T����{s�x��U������&�6�p�1�
L�]���<��T���n{��f���@��0#�fW��(T�*8�eHq�&�)��o�`ݱ^������V���L�}��wr�ٴ�^뾼�yK,�g�N�1��ۭ0xOf�"%�(�R��A�gz+"�� �k��.��U>=���}�B����Ss��¯_�����̹�4�i���B�10b�Gh�e����{�r\�۵3�Նë�(�����jȧ�V�����aM��$��^ܸ�!�6��g6��ez�]��Q�DL'$vǟ�`5!ރ�*��!�mD�8���av�Z�gUYE4�	k�����`/d�}]�3c����V�v�U��{�f0ּŗKdq��2�ͷ�y��:�6�Y��.}����ܩ�	uz���k���%�c<6o������&�+/��1�2���^�v�>�~��]�w���ĵb�4�[R���|�j �u���n���s<7���>���7FR��*$�۳��Ht��n9]��7<�|�#m�WF,RP]p.�tKt��SO�@N��#��><�8~T>k�/��c���y�P[����{K�]�߆mg�M�^�����͛R�A:�t�!�@h&�m1(	d!^�r�bc�mz���N
�9��ܸ*9��g������z�&�ƳxT؏ x��rׇ�P:����R��f����瓙镛���%:}it�c_Et�H���>���e�Cr���e����� z�*(.��`&Ym-�J1\���{�;��B�]mg��d|�X��eܿb~�=|� �SEg��p���^d���z	WPH�Հnq>J�$ңH� �͝�d��D��w7S�>���f�쇌����T���9�g�q�Wf`�t|�9'w;�N{{}y��_����A`G�퐒�ֵ7��Y��8��ͬ����CNJ�[�<'�雮C��r��>yDmܳ��TZ�N�C��Z�,^����5Kv�R9�T��5�<+�X��L��xþ+y��ݼ�h��7*��o\&�:���֬��U�e
Ee�O��݄�z�iP+i�U����om&�=*��I	�mnd?��h�S2�^���[�K�ұQmجŁ�H��`qߥ(��	��óB��L��杗7��א���a��сuM�BA���wٍ�U�V��J������r����4p,.�^����C,M�w�(�XP��y��_W\�Y����4Yv�e=�2d��t��w(K_
{�a�K.�A[*,s(
l���'{t]�#o|̓F��d�NLu��+��V(��
^�<V��ś��g����>�H��y�ΪW2��2�v��yC��)�[����F�Qc�b	���twf��#��+E,�]@,���Ow�`�%0���m�2}�/i��oH�rmn^�Y��g�݉�0LCUD
5���Ef�M4�Ժ�^T=Q�_I/M�5��ܲ����ѕx�t�*�R<߽-�?��f�C�����r�f��͇�u�f�w�=h{f��wLS��y�]Ǣi)�Y��	0�K*��Oh� �%1K�լF��^k�ꐂ�8�rS`�\�4^i�ZR̝�m �a�G��]ŋ��n~C'�f#p{CװK�p��5��h��6�	z��ut�z�^��j�U.6�G�I$���lRUU6�;ԫJʛ�)h�z#@�5�	�s���4p�)�{����+�9l�:��K�sm�޸����&O]l`����.�1�DLXt��8�<��9���%/j�̯�ç�iK�G0ڛ�ܤ����������j�VP5��4ε��Ĝ�z�p5]�l�@:q�S����+�◢8�e��ϴ�ך�Add�(vN٠�=�Gnhۚ�nݹu��n��x3Nm����u���I����c�=:��/=u�Q�gڸr���A���0�
9��`��4:*�r�޼6x�q�c������GY�f^�n'�Y�s�m��P4	wlb���TWI����<�4���:��+'/&�\�uf�$�l�v����v��pc����n��b��V����:��tR��9���7E�Xk��wYs��
��Lv����qs�	���@:t\�n��X:ۅT�\*nS���t�m���x��D�<��5]Xuнv��;t��s���v�x����%����������8�^�zzS��.:��lF�N��׮lݶ�ƷGy^*�sl��.�Gs����]=mˏbywT(�P6a�]�l]E���ve۝��<L���M�r��M�e�X�q$.�#+ێM���]��c�\c���u�N�:�N1�m����۝h�����J��-<���a�N\g�s$i9щ�<�]s�p���O
�q�p�WK��Nݣ�b��-=����y�v4`y���3��&:xM��7Ln(��Y�!�����=�
����g���������qKnSvw�D`w��s>7U�N���Gi�f�90N㧣a��rN]����{����'�۲��к����nݱ��&}n�.w.���Ń�N-�E�A�+�`zU ��:���U<�Q�(��G=ˇ��h�����ȗ W��fn��ڴ�H]��q�˭ۂ�nR�t��^���uy�l��O�eI|t�-ɄS��\
d�$�m�]�%j�*�2˂���N9#��2A�nm�#���j7�z��Spe���y�ӻ[�\pC�%��[��>�H:.�O7:��x	{v�w0v9y(��+ѹ�͝Sl`�ܽ�=�.B�	�W\g�ֻ���\	�p��Ӽu>5ls1�{Z���KȾ���ɫr7I��OauT�l\��s[�u�z�ީ����;�v�=l���]7��f'&�Qf�pd��Glj���E��]m�ڻ���;�N*;n]sD��k�^�m���vxX�
�?8'L��,5kB��~u�Ο�k�X��2���q���_.�w�j ]þw�B�0���"~ɨV�L��}�u�؞ɨ�rڥ:ѻ��0�̨�L~����{K�}�A߼��������<z̠��t�* �T����	"�}�Q�ޢ��h�c�M:QV;�Y�H�����wx<�f����C����7&��|��^��!hE�� �W`�]�K�=���Q�8
�h��<�5L��������:四�1m�w/���ۄ�=C*z�G����۰}�8�Q�l��nEt�h���ɝ��`/
�=B�bl>��{٫��d�&h�h�~��C
E��{�~G=6ඞ�өv
Z�|=a�Eb ���Ć::˨:BLs\�1R���<S�����m�u��'E&GW�;sB�Z��;l�ؽ�W=�y�%y?h�c|[�QM����Q�>�|�]���X��¦��RE$ػ���=[�=���GL�lߘ��1V��,c�b�p�@M�|��gw��q�X�>�h���X���x�������N{�N�6ҳ�7�ό�%
��t���@����<ث���l�י�&�Q����NL�ec{͆�J(�n
�+"�|�=�^��˔�r�ӂ�g�
^o��io�˺���$�������KͿ�n��ץ��]�qhg�� nEȫ=��Ǚ��&�D4���]�{{�_�-���k&Ӿ\�]kF���{+�^'��o�]z#̓x`ʸ�}��\B"ˠ7M̬���bc�~��t�B�O�;���x�r�mL��F�˸g6& b���Vn�1�;�b�0�Wp��B7�w�,��4U�AB�as�x8w��'J��t\�г�C�b7Z��iJH�t��lRi����5G0HV��nqg'<���K�J��¼sW:X�q��<�0��V>�~��}�z�me��Eي`p��1��m좖v;��Pټ-\p�F��������~�<��i�����b�m�\�6�!mz{�N�*mj�m����j�� �l��i$�$�����%+�CM�}�yl��.��9�³(+ӽ�[="�x|��Xe0��K.E���]�fFr��粶��@���&KKT���=7�سq�u���/>��C=�/��;�u�A�Heme�K�i� -�#MŻ��!�w�:\�j�Q�L�vͽ��"N���<sv�ϐ�ا�Y�"̎�}��t�����t�W2����d���R��&�NH�o�J�V���dB�!��Y���ْ��_��n�>Ų�w;����@#tu�����~nz'D�4S%$B*��r�P^�3$�Tm��-&� L�z�E�s{j��4���%�;�[1�+ͩ{�&vRmRV#�ܸX��ZZU��E�yu8Âz�͐8�:�+YS�c��h�kR	(̎&d��E���W1y_�������!�����}睥��R܂����>�qݤ�]g
L�wƷk�{�ԳF�{}�gL���r� �4�M��bwc����T��{��0mߛB��u����<W��~#��!޻J՝��b�[18�3K�o�ˮ�R�G\ۢ���i�L�l0�Q�Q�wA�g�NG���x�j_�6�mH)��Zy*Y�`�Ooz��.�R.�V��s�JK�lL��0�Ȯ!jul
�X�ݭ,b����U����(v�u!t���4m÷�������5�5�v�5����VV��`��8�^_�c�>d��͆�$D�W���Jy���zu�2_`���R���{X�.Z
X�e^�NߕW�;Zҳ����/���W�}b'Ryl-Σ[��z�D8Ʈ���QV�K���2�E�Rjq:�t���M���u��8bQ�����d�7\���R��w�{\"��(j�|���z�H3.�Co�O����)@�AHːfba>�!<����0V�4��a뵍��ʗA7�;YҤ%����x�����E��י(,�e�	}�/����+a��T�E(���.����F����Tҗ��F|����ᰖmPcT�Cv����2P����˖ttht{ȷuوN�MrX�P�Br��@dI��rz��#t=u�o&�=c��HKm���ʰ�b3�e���xy��?`�y���<��|�#��^�[�|����3��6h�Rm2�M��JT�]�d��[���t�pccxzXF�z��gc�/)%�gn�}�N��ʙ'=O20m���U��d���[�;���&�!1V6�����	U�:/s5����jA��AS:�L��6���@�W�aq"��[�8��(n�<�Ev2Om��P�&pr�u����w͂�'�ܖx8F/v�nsv�+\G�I;��ѧ���s#��v�{Rj܌k��⫈,������utQ�uj�\��Zx�x{m�q�gA渍��ݫl���uQ����C��m�����]����g�U5�����n�'tX/<�	ةɭXۃ�15�~~���Fո�۞̜ۤ�ۖ.�V�-�q�,�pvusĐ�;{R]s�X�v�_�C�n������5K��uxFJk�߻�n����{���z��X�Ϳ����moQ��.sT�7�E���~�Ih_�5W�:�ڻl����������#F3"qU�[(s�Ϸ�IL�<��{W待�*�	LB,�꘼^�ew���o�������^{�x��ev���׽���%U���� �8t�SmfG�{|�nŶ�ʷ�O�Hݒ։{flk�F=�3y�g�̄N��W��Lp^�=�q�2I#.F�q�"��u���2��Ӵ��j��#���xf�3\)�0G�)�C]��|I���ѽ�W�g��m}���h�d�I��3�i��^r�W,�PA�	�,�/8��	�����s2�����r�;@��o���kK�ŗK7da�{��D64������p��c�Q��;{svJ���M��l�	��i�=S��e��������Ϙ��'�1��I�c���J���ߍor�뛍=����,�9k�A�q����I��7	`��b&#�+zN���g��
�3N�A���P��fu�@T�)�e�N�KPTb��޳��8rGVE+{cn���L�,Nbՙd�����{��7��,\;�Fvu��et�"����'�F;M)TD���� ���g<\8��~wF�Iu�!GjFΤΉ1;�zb�2�:�[��d�����������~��%yOs�KP�G!ܺ{Ѯ5 ��,��������m��TKa4�m�u�6�{�_�_�S(G"�Y�=+:S�M#�vzQ���HSJZ��~��=+��ԁ�t{��{����'�շdߧ{ބ�cdl$Ą��*#ZhK��{k*��)̦Ѳp[���I*�Kns}�JC�;��'X}��Ww�Û�66��c{�]��O��3V8�mg��rP��tkg�C+]��I�]j�6�����ݿ�������Z��-��7]�R���i�RK�4x�L�N����geN���X\w�{¶�1�gJ��1�Q�p�#�fz3����OM�ͼ�J�G
X<|FMb�@r�W�
~9�%������pң�/�X<.OA�9=���l�*t�8�)H(�8o����Ŋ{ʵ�T������x�_N)�d���m�ڻ޴\Ы+@я'�Y�0tJnt�2� �i��e���yq�3Z4����Z7��V�8i�s�#�}} �FN��7����Y�1�gY��N��������̵o�Ʒ9l&m��d���V{2�}7��tf;���E�]AR�V�:��'�٧�H9�+�=����s�)���Ki�)�M [���cj) =v���xa�S9��&�o��e���ރ�j�e�NhA�:w��{��S�+�!�f��4�U�y~��ߴ�q�vli��\Խ�g5��sk�.<;�����f���i�nnT��1,���z�	|''c}�^vD�;�g9���BByT����u��ir���/�$R�zĿE/-�V؄M�W�� ��I1��Z5n�Q��y��ݜ��`=�g����cνS�f�iR��M����rN�!تp�걷�E;¹�@��!0)�߭L��{f�zɞ0yD�M����w��{x�NLZ��(X7Y��T�� om���e��4�@"�g��ى͑��_Lݗ�<MqV�j�3��#Tvv?��W�cf���9�Ԙ���z��N3�9b}��S��Q�y��K��I��3��U�+%�+t�kg<zIw�x����	o]����mξ��7'����K1�Si0܊H��}*:oF����蹙�* ܚ��d�^���/��w/\�D��d��tBE�55}���_w�n��}��޲b琐3�Ўۚ�ī��w&^ў0����|��"�FFt,@�}�2H�]�ч7I����C�HE���g5o��~�_J�<A�M��=��w�>����so�E��lAI����{P���Um�<�#^[k���[#]>Wш���+g�m۽`�j7Fϲ�F��#J�L �H7.9WW\�y$�qn��,�*�vv���V�`-��u���kW� �ė<u�gfx�;7諎h��)�N�4�L���*�;�5x�gs�L�o���֭��G�X�h��.���n�sͨ�����'�7�S�"(�!��pw6O��JtB�(�u��K��5����v">N�MY�ȯ�J>K���K%�{�r���3o���r�˿T1L+�*M)���53u��
������*X.������ f�)����ز �>��,�q�$�&�6uk<ꮞi�\z�P��a��ogs������W���;=���4�7����t�qe�CF^&=��g�1Ok�,�&�ۍ�U>*ݑ�nn&_&Gc���R鲭:����s�N�k���8:B$;�!�S���:3��A9�r�<�>{WF�,��\욓Wg1����qغ�857n�O=�7v�9�1�a[���f:ï��v7�>�n�3���OJv�n^=�h�Ε��m��kdy�/K"�q�P�OUOϤ��[�Û~�y�KKt�x{ w��l���S��[��uh$��|�CÍo@l�7w{��l$�d�"�m�#Z�T�+q�5!������A:�gd���}�碘l[����ñi?e����t�R��-��d��%2�b�Vk\ [Bcלָ�]ۻ�y<��y���.���?tW5��'79��vܒ2���4 d0)�E�S�%Z��b���s�������=u��^A��Dl�;+��m��2�	�o�{w�d�%V��kg�w ]0a�E2�bɞ�/|2z�u�ة��/c��\=A�t�[G�*S��v�a~Uet�u��U�W�8�����T+@[�5;�F�x{�K;ynj}�fF��zݑ����V��x��^լ�V���w�p����s���vN��h�q�r�M���w���/�y)���v�^���ޯj(��:!6�2��ٸ����z�N�0l�4L��<�KC牐�n��y���B��ɵ�3��&7�'�d�����Q]]	�ٔ7u����nV�ٻ���gc�=��+7��׷^��4G�n�����,����\���x���=��	���=7��A#�Cz�!Q�+3iTp�J�~��o�ў��ŴY��?=�H�o�����1h,P�}�4�Nv濺MY!�S��(1�8���"�FUYq	^��96��2�������Ի�&::U�rV�Y����ڱWe��U�t`�x r8��)�}�[U��=�i�K�z
���fq�	Ъ:~�g0x�Kx�S����܇g�T��W�Ћ��R&Bi��P{uҽc�˼�/5���ϮR�4h �z���m�`�	6�g6,~S'K�{��Q{Wp>��ᕘ�V�����<ݎ!�ܞ�̨D9���^�'��V]0F-I��خ^ೞw�������+���xP�<Q��ږ�G:��>�E��}�t��1rw����k����B��J��0�-��2�?YHz:ءw�¦�*w�9bạE�<[}�E��U�ml[�z�A���	Eɋ�lv�u�s:^�n0���/�	x���/C^�ֲ��8fE��E����9L�8�\�=t�~	�} �rR�Ed�V��s6PpS4d�����>q\�+~�����J9�K�Z��ؙ�o�C��h���3eiûP-F�	��_U��&����}OH��4�T�իs�n�=����iNٹ��Kٵ	�n�d��#n���S��2�XMoooV�F�m��3ueC��M:��;*V�q��}2�VaB"ʾ�V�.���/�yiq�S��K�FMz�ou����a���T��Yd�R�ܥssK6P&;��졛7r��}ǝK�W��D�F��u򅎔�8�lJ#z�8��m�q�:��0�{�;��7j��Ϳd�-ʙ&��ؐP���wf�[\/�f�i���Y\
��o^n��=X�>�!�j˼rۮ��h�
]�zq�
^�7��Wu<�����r�A��m�)��ܮ��YL���C�[��;2�TN��Q���Gw��[a��}rv*�J�sqi��gr[���k��
=Z	��',��9F�g_4;w*�*��ǲ>NiM��k���XF��.�u^�w
�L��DK�Qf��x�8%�2�9��q� �h'	v{4���o@V�y`g=U���|%�߲Ccڡo'���L��<.�l�*���ˠn��X~�r��>��uF4;�,�r�]��U��wQ��\�����z�;/6���)�����<��(Y�u;��V'ۉ��2�Sb��L�)��m��<����^�ݰzT�/��< �=�zS���ՙn�,��ޕ����[c���̶�t�����-�¢�a�r�aAn��zQ��w�����WVW�}Pdu���}�SK}�鵛s�-1����;�ʑ�nE�<�U��H�� ����\�gu����t`Cٶ��76kT�Sj��`PQ	�"S�[u܋rq�Ds��x'Z�A^���]��U�6�d��o�{�GۄR�[ڵ���&��k�Ԕ�	���6�����"���$QE.��
�����z��#��N�����J�K}���˯a�>
��L��+4��+<�0ݼ�/����� �%�"��@%;Y�M�!�ܽb�wl��S(VXǖ�x�j����Y{���M0���|2�a�ޭ���;Z�A @M����k#*��/kr��en�3�����b[���rxu�˭���8��V��E�t�Y.x�ctX�?�&�kبhĦ��`�D���%յ�d�o��[�۹��62+��$[>�-M{=��`�B��͛3����ﭝ�w{�N����3�a��N��ÞMkr���<�J�gh���:o��3`�؆M��{Iu��{-a��u��뙭K��6�ʕ�+��ᗗO䷆��y}���<���g`��ރ�����g��ٹ5�aĤ��R�����>zZa�l>�7os;f�/+Ë����]���'S��V�1�y&����h�bJ�)|�[)�l�W^��#��L��I6f��c�c�Z�����TwQ1����q��ZN�����y���^���������s����ne�N�@[a�� �2��:;��d��A}R^	⧐�;�ī�{4A���?�'�g�-��k�y(cm�̼ʜ��q(R�$�P���V��L�%������q��=���C��w
7������A���e��V/�������EJ�$E�t���m0ﰾG�{EXr���x��謫3h��obE zߤ?n�E�qK�]��T��'�fKG��}�X7��n�ާ'U�uCͳsCպ�����vE�6�^"ȾGwviY��6v��z���0;x:��C��|L�i� �{f��Z(�v\��1/:����f+��TlOn�nR��nl����;��^횐�rݶ�G3�8��:w�`�p�Ϟ`z�C=-@�Zg�g�{�����;��:Ѯ«u��Nq�0n��mW���\������:�IǞ�Ik�v��8p[1sVx�ь7]��6��!7({z�=p.�nv�3�Z�Z�t�F�=�Hs�k#G��ڌ�Z����ö����pN�qW3���>�w=%�l�vs٧�$ҍvw+'-b�tW$ؼ�?Oܠ���w��2�U�2��j��A$|�s��Ψ&٦yl�՝Yo(7���^��e��,��08Ki4܍���r,�w�,Ř�f��ag�'����KM�� (Qʜxl��ϧ	����� dY�6}G�I�u��H�lR��i�su�>�PH �p���c�(`�%�}��/C��)�'����c��\�t��C�1�y��uzE���i��-�OH�k��/���Io>���Do�t��dY=��i}ᔄɯVm�rq]���u�EV�R��l�#aIjH� �.�z��$V�G�ݭ�Y}$���ίU�6�^���Fl?'���/�ٳ�d��R�)>r�˪�Wy���y���:sל\9'�vf�3�cp뛹�%�K���+��vw��-t�[���xK[�ίkѲ��u���GR#��m'a]I` 1��L���~�������~ ��E�@��-��^�LO.�u2X�������xn�Bj:ɹ,����L�c_��ns�ܱ{Ru�4�r��2�&O�d�'ݖa���ֳz]�Rb��$*��s=9L5�؋��x��W1��Ŝ�R�Q�'���nϧ�u=W���1��Q٥a�}'m=Q8�rHÐ��sq�@�H].л��vc�<-�
��˩�M������$֭^���vF�b�W�=�~�쮓~=���@�		�$xM�DY��ZO�:�ޔ����3=*A��E`�IM+]I����s6Um��_��]�e�AR�
�L�I�N��J9a$��٤�Ϋ@���T�Dơ�{�Wx���W ��C���*j�ػ�9Qs�ޯu�JɹYa{��3=�KL6dI�h�K7���<�z�!�F��=�V�n^��p0\M�X��̲���C������S��a�l���� ��v*���8O=��/�*˰���,�@B;��������n�t��<�	 Y!$R�7�cks/}���jx���]�����~�T��Hy�2t��J����Sk]OD:G�����WS �X�=dB���8�nCW6oe1!�u��g��׳�ƽ����P�{�;`w��o{Jʘ�;ׄS]-:Ȥu��ks��6�l��$��.u̫a�2��m��Sj� s[��uӖ��
[��̫֙��9�L4[MQJ�!BW�y
8�������.?z��q�Z�f���d����03}�����6{&�X�cD{z�@K%]�+�	]�n�;Wc���T�!e�B�{k�"������oҺP�f:��|��.KѺ�1SLJK8A".�c��3÷�=FN{�m����ָ���K��Z�.�t�K�]���=7߯�p���U�=u����MＧ��ݬUݶ'�g���.ؘ+�@���,�Xm^�F2u�=!�|�2���ERtSbX����:G�*^��k�s��㾛+2JO��4{��X"+�K�*ݽ�X�ӱ��ފ������B$IT�8�P#�Ϭ[��竩5X�Ie�i�o,��n��/��u���W+כ�AVů��w�����fM�D�38M��-� Fa�z[cf6\�>���ʷ�^���S�H�o���';��cK�=T�a@s��>�K۱�Ž��יw�2j��i��N�=ٮ��e�N��
�	�ѭ�QN�4tZ��Aʶ�n,�U��J�����g�.�ٌn�t:
n�T�l��v��E?�E5Ɵ�ҰT��&V-9z�Iz�.�ͥS68��Wm�gT�J{X�������Q�	�"@�)�ۛ���k�t�*�굺�[���3�Z+�(zn(18��D�rٝ����zR���k$Gˌ�^S7�5z4�шF]O[mG���:~�v�V�>TR�K�1�̉�$.&�e�..�ݗ��s,h����?7��r>|�����c)�Q6���7h桇$t�9��=��٨�$�l7l���*$K`�S����~�ʻ�2h�w��ޘ;Q�Z�����|�=�N��:gm�o��\�<7I~^�T�v��l�L@�`Q�/��uOV��T�y9gg���}�N[�f��:Ż6(.�*��0#p��ݤ�t��q���烷:�v�B�}��t����&��d�����[v�h��ִm< H}9w^�ߍ���O�z�S��-W�{r[�-^�yfd��]��6TqP74N˭Vj��@ry��i���Kɸ���j�m�\���8�2��7����r�V�����k��JI�OLۚ|]��-�]�d��g��WE�Ӱ�ׯVY�����n��磆c�;��U�ӭv"��Cn[SDB�GY�Ӯ4r+����}\���ϗ�8�Z�ϱ^c�}7E��v��]�Z�F̋�N^6�y��SnY�nv�Wl����]�rBz��Û��2<$��:�	��p�N�l�ۋ���J@Tz֩t��cKϞ�/P�Qv���|6��v�X�ng\�i3�5�8H�ס����\���)���n���4mW��v�9Z�H��߬�_�:n~���.�a�o?\�p�@�p�x�� �l���dp��cX������a/*�J��=�ca@IF�*��j�9Ef\~�^_o��JW��ݷJ�����zڥW�����V���ۖrM�Khf��y�=M�$�N�%QI�����uA�U�w{a�Ƣ��e���=��*�2�i<X/ׂ�g5�d�p����+>7��y�H��
h�l坡�7q�f?o��w;�1зV�ۯ-{Lk ���[�N{��5�T�h���ݜ*Ԁ�:����ލ�F�<Z�a��e6�-���
������x�Ee��i<��Stew��w���(��O׼����j�ܳ�[�o�J�m�IF�]r����;�l�����l�u��ֵ�Y�[s�rr�P���8$m�MO�qU٫ǵ](:�OE���Q5~ś��3��,<�u���qhQ{�J�haBy�ND��]24i��x0��n������췘P��8}[�{d�77rj4^+7�sIڏ2:<hkh��.�B79n���J��A��U�gʠ�Y�X�U��nex��C�/!�U�<J�K�������c+=#C�>�Ͼ���d�$�)�i�Y��֣�)P=�X&]�Lќ|z�K6����iM��+�}^�Vl�2r�!}5}�?�2q���t)�M�G�^�#�}ӔYW�aF�o}�uj��L��P�"�h����75U�|��m�Ǉ�`�E�Uh�`U6�[A�}��A��V�<�"&�(;7P���V�����	�ʶ�}�J^���;Vd��{#��;�(�w4�FG16��F�eG72��n�\�[�v�4��#�Gi+-��L,�:H�hQL[m�WcQQj�Å�=�|����,�}���T�k�1��{L�WT=bZ��p���D�p!,��l�u����=������m諴gL�1�^}�Ŭęo�[�b=^������5>��ʻ�c�=V��i��m����-or���M��g�_�r��r����,�*��F��YGFy*���G�l��zJ!��N�uf�w!So�.�#�ǝ-��;0����	�{�2�s:T�nT�iC��X�N����^ny���+�E,q��m"WΛ�N�I�3���e�0���*wF����$(���_+ޝ�۞����Fﹴ�����'�=�;������C��hz �G#
���x����"�T�LR�0�;�pG�'b�WȽ��)aL��wk��V��8H[۾}�М�W�i��K��!��2�\u�n�nx�\��d���˖��uι�i����v�tK��e[���F��Z�s�����{��k�|�%G��*T\���v�g.¨7�o]���iU�=�E� S%6g�p��y6�t�|�2��<���"�S[��gx^�9��T��Z�}�'x��&xwpWUxL�����m���)���m������U�#�ѭ輰U�G�G�糚�;̟3�����9.�����g��<,aYM�u��:����a$
E�j^cS|���^��]tb\���
o�	��4�b�>T�oN�x��紸+����7s�Ƨ�*{�{
TH�Ν�L'rib��d�7{b����*�k�L�RU�~�J�f�9+:��L���{X}S/w��n茓���l����q���,�z�8�نz�;�)����o�+���z��A��VL~D�Q 5����كU�	��Sݻ['�xb�f$S`�#A�q��.�P����q�A.18"��<�V�������!R�4RE+)_o�0�6��l����u�m�q�:g��h R)���d�<���K��������	���$���ѯ9Lf�	�t��a�x�"��,��s��g��.0��{x��ʁ��u�(ۛ�ԏ��^L��;i�SH�I��d�z�.�F�wV��X��j�t�=��X��6�g�^��>��τ�`�'�B�N���t�N�Lׂ��JfY"34z�2�f�O8F�g]/.�)z����1vT�8���x���)Zuvo�û��|�\Z+�ǭ��h�HSE�%�K=lEC�ef��g���N��Ժ�\�}�b��-�5�>o&�w|���=���X���J��,�.�	��ki,j3u���Lf�%{�V�X0��@+�#��d�FK��5���+ʓ��Ɔ�Ǐo�U�eZ��۸.���Y��6��K�04����c=f��L{n�"6�^�
;��0e^�?L�[B30�v,��6��M>�Uw ���{GL�N��٤o�\͒2��f�^T��|��Ɵ &`����M=�on�:Kf�e�T���}�Z/��aQ����w��8�ə�m!y-�;�sĬ����J��L��U�>�ku)c��Yw�1X�K;}��ol���Ń�X3�4�&���=YJ��;�2!�ī����pU���.�u�"4��t�V{3{$�n�#ȇ��1�m.��6Gr����%>��)�Ǧ��Wd��q�m�v��w��-���s.-���B!���ف8uGewFY܃�۫V��)��zm�ʾ�m�l�IM����ȴ3��Y��Z��9��n�m�����o�]�
�껡�UմK�с�j��:
!�.����ZB8̃��
;�n�G]��"�'�(�� [X�c8󱲦@cd�^���X��S�Z{�ʭ��z��t�ViA�a5�m�G��4�TZ�=OE��Vc����>�Ob�H��|Jk��Zz���㭙B����)�J�!�[�E�RɲX�ҳ�V��2)��1�eJ4-}���/~��Y]����t̮���q��l�8���gA�\��`��iv���՝�,��+9���Lu����t�,�AZi�0Y�������u��ە�]�b����t��ַ�m�\�v6���6�7
��G/<h|R9S���[��d���V��e]]&\&�E���[���B�z�7��)�1E͖n���vdz�9rP�`��f4`{O��v���繸ϔ�
0_8�\���o��j�sgg�v1zQ�;��Z��q^5��e�Yb]ˣ�xgp\�dfΈw^N6�s��'����GO��^x���vrB���ŷ�j�ɺ����'s�]�m��,��M�t�#Þ��ؓ]����vk�����R��.��\���g��n�S�u;r)��)�Z��ݷd��8�QSI�N������Ӟt��v�Δ�,��2L���8ioT���a1�h�{�KNt�C�,�s�I<��\ɹʵiy�>|]5������O�Ĺ���Bq����j);s��uQu�v�:^]���v݇�u����.$P���:����g���q2x�Q�.75H��Ƌ+�n�V�me�n]b�U�:�Hr���]r�����RC��U�q�\�e���V�C�V�h�˺��w�O����j�]8�勳�W0��N.v�Qδ�m�lN�vAx�ce���W���>^;wn:Y���:��y��CaGr�ۛ]�zyR���NvwI�Rv��`[�b��v�.��;P�f.�t\���D��,:ۅt������&�S�;u\�4�8����O;F�ױ��XyC۲�ݾ�3���Ť��T��G3��@��r^�-]s�VC��h��W��\v��0)9ݱ�:�x�^����rOlgG|-����t�4UϲX�^ty�헡9�s���#���C-�A��1����#���`��ѱ�Ӻ*��u<��ێMs�{r��Lg���b��a��掋v����v�(�q�1�z�Uqۡ�q��=����"}�3ŶS������9+�z�u���gn�;vK8�%���,/ce�wVzۃ���p�/�Sƹ��e�$����m_On�/Q�<}&�ؕ	q�,C�6��!٣@�ؘ�ۚh�n!��vo�:�lse�{d�5�n�2���23�]K��z�j�Mx\qДa����^�s��F�=���m��X�Ft�u�z��by
�)L�Λ��!]�i�v�e�e�v�v	�
���fx�yW!.�O@M�l,�v�����3i�[��{ZV�ٜ�Ħgj��7L]��kX4A�N�0����Er�1wj_���c��G�N����̼t�f3]+h����AzOY쪩O�_�Q�̅6���zp�y�
T��[�����w�YF?^���ZŨZ��8-����o�[~ܸ/Ҝ��]����g�A��v+�M�l�� E-�(�[��b�U�-R�f����@W����}���}�ܻ-s�f�;�9Nזl7�<�/���G�P-��M��a�{E��D�y!�w��q@?ku�]�1g���j�Xp�����"��v��Q;y��3������g��!��D$�M0�7y�ox�b;�TW�RV��dz����$4��S�=�3��,QK�����=�Eл�����$� C>1�MHSt^^5���'Xێv�)TM�]n�������q��̈�N2SB�q�;���|w2�l���Z(��f,�)���;����D�z��f5Q�x��
���ޕP����]�rH�� �]u����Z:�a_ew*���U�Pk]9��y��R���oyu>��z�tNs��Z"���
vg
���โg���W��/���'�Gr�p�∌ԋ�8L^>��$z�������M�,�&{\@ �P �幗�ʛ��/�z�[`߼�Jr��v�Y�ݼ�������n����{�^�&���@\��,2�-��&�%�w����)�����ٮ���Q���Nۡr�W��~=�H����37�xc��v�AD��j- ��H'E�IaDq1����Q���U������Cy3�龌糡�f�b�̋�tp��_��6�����͝�g����J��u���p��`��^�M�	6���Xy���I���M�:bE������R��H�o2^ o�M?%C�f��@[�;2��ؕ]���n��3���I�ڼ,���{���B�Q� ��e�:cwN�����M	:>��m׏��u���
Zc��P�y��]���A�b&���tVp!�08YV��	��M��i��00we_�,�u��x�̽�!����ces	[B8)�<�	�=����d
�̓2���Z��gY9}�K�t���Σ�ǂtͩO*��O��n��
g}�eO:s7˫��uer�={r�����M�l�S�����qW'Ö6�M��bYv��e�>�(�A�-�m'7!��Ƿۘ�*ȯ��!fG����l��]I�{����'���vj[l���C�>��1�1Wc����ޗ-��4��.u�P�ܓ}7ү��{@*�|< �+�s�I	˷>�㭺ynwe$��]�⎏.��:�B�y�!pqa������0F+�\|���r��]�*ae|��4w\������B�i���8��TMo��I��
h��&�]��o=�G���$��o �t�4�n�}���_F��7q��ط���M�u�3g��RS>��:��ev�9���M��M�)"�~f��l�ۯk��7,�����ς�d�ף�%���9��ٛN7���8�)��h�6�pD���������;�~�)�[h�`L���s�j"��j ��]�K��p�kpԑfq"�yy%��L�I�6��u�7�[H�.J_v���#��0�����:�<컨���Ď��L|��
12,Y�!��oWn{��Q�rt���h�Bar��l�Gw{���~�l%��G�X�~jv�U�<Z;�^����Xl`�N}�9��Pm���`����,R8�,1!N3*t�-�-�n����p�ئ�k�����嘶չ�qCj��	�Bm��n�0G�x�3�x
��O�`:������d�����J��%�Q#�Ctz���>��f$��<||�p0c���<�}�:н�v��}[[��v3ez0`��7]1��:�U�X�{|��l�q�+Df�����͵�x�ᐄ�a�P�#�|�x��<��Ka�Qf���Yα��C�������Ҏ�Pul+������ܒ���1z���TKt @�M�!�~[���/rC�⍎���e<wy�)��<6b;:ם�����9���^zE/!U��S�Y���Ā�m:E3��Ά�L��.�0��So;�K���t��~�x��"�)=;��z�͝���Xo���yS���J.0ؽ�� zǐ�[oT�<eL�*{.:tÏNp�n�׎֓�\����#(���ֱ�+9�a���̗�9�q:o�8\�Ns��r�֡3�c�{Ml烫N���)6���]kK�k��^<��r���ʭ�v�w 8��S�ǋn�+ER���g��Z��� ��΄�u&8n��O��n�b���f�q���&I�a�X�i6����9�Vc��N{�ɫ)�X�p+��vhz���0ތ��L�v���W���7K�����Ji���.'q]�9��ոK�E�vsv9�B��	��Z�������(ӵ��Qm�
	SH�Z}6f�Fe����Ss��Vx��ܜ!����t��L�ܖ$?A5y��R�@�
�I�5�8e�rO�ϫlG؜)������Q?7 ��Gs�&�ɽ���	^nUׂ�j��κ���L4%M������-�!�Ǣ�7�z����s|�9w�O�}e�t�=�z��)��u��)�
l�!$�i�o��p-y��m{ï��m�^G ��]��綆�La[�^� ��yړ:���72d{��t�a&�)��C-���[���u6M�����{����e�]��������W �욇�&ku�Z�~j�'����"��kK���l#A&�f�f2�(�;CQ7n%�1Ύt�sfU�:�6��]Z�G=�)4�:)%����.��>�n����e�Rb���L1NޗB��{�~����3�V�]^�n���[�����A�B��*�(�;z�1�<�#α�h�9��zzl�f����N�sB>L�h�5������u��rIR��n��6:Ԭs���f֐�,�nn��7J֛�Q��1I��OxL�)?z��\3��Yz�uY��V*>|B��UJ{;������W���JB�c4`�4�X���Ya�Z�Stu����+�}(���� ��B�f�쨕�
^���kVˡ����;�!>�
�����~�	�kf��߸G��A{�z�t�K}���w�sF��z�l���_��}�����0����i�H�[m]��c{vN���էjmx,s���z�mgSi�F��%d�����l~y�g�^em��.ݙ����%\��7�Ѷ�ʷ�z-��ٺ�Z�G
ݳ�����1�H�4�+\7[q�ƃ��xi;�t�iIQ��\�e�'�޿y���-�Kg�p�\���^�L��KT�)v"���Q�C@�a�m�@U�oxc�G7$��蠽rxv�l�ã�>�ya��l�\iJ�=�r����DX�)mr���!{�4�I�@T��G��Wo����G2����I�;����G��l
�:ɻ7F%[$�\ �V�u����+��\	.�#��r^42�75oV�7Ib#:n�Tt�b��a[p^l���b{˰��f�q�2�
��?��Xw�~�1,[�*玁L�6H�*��}��9���虎��-�'	!����;��Tl��=y���� ���]	:�n����L��=�р�� I�d���7�����={��-ӏ;@,֚��Ԅ�W;�E&�+=3�^A.��/@;�&���F\.�bK�~��v����!��d��E0����s-���͎ۺ�#���mS���v�6Ӯ�$&(!O�D�r8��ѵ�P����{Ԑݬ�J+����e@�n�9]����=S*�[��B*��$�j���f�1�O�����D
a@���L�/����鈚���z��v^gȍP�*{��6�Px�bx�I*�1r�z��,��$���%HQ�9	�ys�xiy��>m�tD�ޕ<8���������o�L*�|�}�9����Ȭnr5*Í��o3}3k��+���+���N��[�G���ۺ'��6R5��#���}�/<&`�ZTr���#b�G���F0p4��(i�{Y$��xZ�x8f��@3;�����:�ʳ7se-��u�]�D�����L:M��%��a��e�I�*��w�焃�����̇oգ���X�T���Ƙn�����ad��2�l�+ v�4�;���n5�ٹ�mwVkҔ��t&*[ůj�Y�L�R�20]]e��?_�;"��/l�9 F��Nv����$Ӵi���M��S� ���j�j��z7w��Jtt���yF��.�Dآ�J�������ص�m_"�9^��=	����3׸��K�����NXo��;���T'g��X�ye�b�.����P)"U��B����8����]�!�fd�Je9=�����{T��<N>sg:%�K̛`���D����nCW�P���/����{���r(��E^��|�W��^�>H����"R�i��د;�	���mQ]K���4Q*T�m�,q��u0������|��o��Ew�
������͓x�aƮb�<�����|]��`w��W�S�H�.��y'���ܳ���+�}2��A��@��U����5�r�;Xv]9���x�{I	����D��U�"��OL�.!�KڊxN�GU�A�����D�������:��na�Tt�:\��]F7Cc�W�x��t�m�W�2u�v�������qCqq�Â�۞��c����O��[������P����\�n)���ϝ�\+��s���.��<�X榰�j{[��� ��sgt�k��'����&���pט�Z	��WR�f�KQ�-�3��ʼ�6u��u�mg��,k�F:�יNsq�[�T�.c.�@��x���r����ycw)ͫ��1��m;��o:89����}��y�Ӯ�;u���3�+>����	��1"���[
��'=}�eG��d��3MX�u�EC<2��,��.�/]5v!�._יJp�t*BPE5M2�m�v��T�@G�t_0�T��\U��*�����/%��(��C���I�|޻,��*��<�[��0�n�}���n�
O+�V^^�m�~5k(__K�<y[��[Y��������ZT�2z�����"n��ʅ�ԑi �#a%�>�ߠ	�X�nN&T�T����k��Jb����J* {��E���ָ��q%[��[�S���_���u-[A$��Cl���*Ӯ�r�g���A�����z���k'k\=ni�	���m��m��>���5w��:�2�ќ]��/u�k�c;�k7��	�v����
ž��⮃��T�&�E�S�ǗKǻ^P���m�4Q��H���\N4=�_f\�ؤ2}�ݷ���כ���ۭ琋f�8����V<�{�m@4b]�Wk�Ì!�h���4u3�Xl���#�1�7"����&pݾh��ւ�߯����'�%$�pH���W~"zP���6揩�3+��X����ր���0����G�*����@��;7���@"� �6� [eL)o_U�w:e�ӹ�Uݯ��s����蜥�x�@v;�+bXE��X�|'����1͘J��v�o<d��M_��)I��r���ކ��]�w��?.,���ޏ� �����%{u�wo�;��Дqj�TG=�{ҵWW�F�;�R��}��\����^S��X���'6����wb�c��m�\C�؇:U�ц�>�uf�{��|�CT��U��fp�ɽU+Ԥ��L�]GK���ԸF�
X��,���Ez��r'���(�M��uuf���<�xʾ�{�#��Һv3j�Wp��}D+#\��lH��{˄�?"A���u�xVU�w�d�L�U`C��B&E��ݭ_JN�.y��N_�����Vn�U�n�7�b�ܺ�>�F��KZ^��;e��h?T���e�.�YNs7\�\q��[�0;�� Q�\e�p�	V��J0v��뾜䲵X̸���/h�K���,�ѫwdv德�z��4^S˷���kGC6@�p�{b_�����!��Vl��U���r�r��wj����˕��L�em�Q�Z���]G�ү{{��4�B�N�/j��*�	Ν���ݔM��}�^�����K������Vu�vlnƛ�S����66�қy�M�e,�2�lJ�����ٜ�0�O땀��N6.���c�}a��{���4�%�Ų����-���AY��չ�_ױf��`(L9C[MVunP�.w��5�͍^+�n1;룚���\ᯰ��Y�:}�*mY�Tt�62U�c��`�#��۵c��݈h3��FR�뒈�^�U�Z�)K�b,<�/�w͖���8Ё_Py�Vq��3��Uu�fS�MIW]�m����}`^8���Gn6ör�����YO����r�ݽͩ���M��:W7�j�2��]�W^d�7�u�o]iC������N�D5���;�i`}�Z�1�a<���� Dl�h(���Q�_�鳃��Ƈ�l�u^$�0VZ�޺@�>v����{=x�>�63�
ݦ0�6���U�$���zi*�]�N���JKR�zW!R�Zz��{e�x���� ��*C��GI�ב�r�0��2hU�yo߯f�r�Z�ŝS=Wۘ��墦��k�A6�{�~�lp�0�=$#�2�m�Ϻ#%.�Bf|h6��'d$_�K}\��Ľao+g���\�K�iY�|.��`[�:T��nջ�jC�G9g�0<���xױ{bˢ}��G�ǡ(���p"�t�J   ?��l_ׯ�ȒA�� FΛ�=y8s*<�(��ܯ5������k�Gs����`����c������ooэ$FX�'�P,��L����l�^/����[�����<a�KqA0Z�ۭ��W�v��5�/�v팱���?�'O7����z h>� ��]x3�0�䘧�kK}:����q�ʆ�7i�sj�_p$4)��!�,��Ʃ_M��X��w�v�]���t���m�
=q�,�.k�������9Xg�ə�:���|1C^T�sT�u�x+u��+]n,.���IMؠCL��x�<��=�����7{�/�X�<O�n�B�^�V6�I�F��r����t��Q��!��Y��gt�g�!4�U��C�	
5l�⼥HҒ�9^�ژ!�l��V}���PWY�,8I]/�i3�"<���s���x�=E*)qsک�O̜���w=�#��K*ж�p��j�<ږ3P�"�-Q��z|L4fH��^�X�ؽ�:�qz{��q%���h��5t�Ƅ
FcA��E �#K��aQ���<鱶���4l�owD�}��=�ξҶ�Ҭ4Ǯ��Q�� ��Ш^�"q�{lf�a�����xp�wtIj�_�߂<R��g]q`[�!��nn�ѭ��z�G��]6hu�V����s�4
�C�&�J��
ǒ?/����=E��х���Y��먁���*��˯Y�ly*���w�؈8s��עIT�;^����T]��I�e!!.F��9
<�=۠�~OE�վ��W��T�����\�N��M��K&yS�TG�v����3�����ᳳ�;�q����m�#�����zY�t�������Q��K�_h#wfU���]b58�˓���7�k<����y�S�!�ʝ~r3��dQD�1��+l��}�"�t.�= "w&����5/�����C��F��j>�����v?��W	���݂�y�QG�)�4�4�7���uw�E�-�H����B�X��
��m�EȢ*����l�Z��߇��x�еN�؎�/o%��2ثF�8)�_�ں".{M�I�3M�"���,�i������e�>�xJ��"�(1�78����*�I3lP0vj�������~��gR�i�ݘt�8�S#�Y��[�⪩�ǮJ�t��=l<����s{����m۹��{�W=\�X�Qy|aN�Y�!�AT,4�0�u�{]�'����ヷ%���az������g�vy���x�ܽ!�%�7]����j�B��\���qX��Sm����i�n��^��bn�X��;w^a�'33�6�[s��Od@�	q>b7�M��A�C��'C��y�+�8�ׯ�yE&
��5l��W+D�3.F��_|W�d��}���Ӓ:�t{yOfרXi�O�4/�8�	����[�E��8�"��mf�n�[��sH�"�y���Fp!m��4Zn}0�Ѯ�?�$�f]K�A��*yXc��5�r(E�>���Nh�W���Q����cM�zD�/��Bn�o����/�mV��lQP�M2�^ 
Xj�ɞ�vL?`�ը.��ʰ4R벮�������W9��r��jjIEP��R���^e4+P� ��K	�B-�p!.�pȏ;��ն�uZ��jU�����+�R��|�~�J�ECߌgu�o���ܺ���3텰�1��t�=� B@Y&�B�ED���N��G~��u�	��{�;YfT��ԏ��o=YBܼK0S�{F�j��U�V��.�D�d��~�׏c���b<�z�yr�pz��ܡb]Ք���)t�G��W&ƌd�c�!���lgv곆��J��ƐC\�sr�������WI�L3ޓ��&�o��4	���_%֖=ޚC� ��e��"�4{/u���!��Q���1H`H*�Q��o��(���?Of9�:m����$��� �ϱo3W�hj��.�L�]�/�f��(wi;�Y*]�S���E����5�w��zxAŵ-Xz��O\ B�U��P}k����o�z�3�Y��[��ql�u���b�Q@�Dn�2[ffr�s��&P�k��[XR�,��=�&���<�P��w����Y�|4����]��g��~� ZO���q�����O}GœN�f�ʈW/��岉��/�:�x�[P��A&K����������[GN�6���/�����{�t�诅�hA	,p���كұ��9�Fed����wp��({�n_c���	��q�%,�>��1;9S
z��c���3N��Ul *E�l6>���Z�u������]�ݱH��H��]n^��cs#�4�i6�ӵ�J��2ݥ���~0�HS][]c������)���Uq�N���Řz���U3"u|�NR
͙f�E�ФQJc��`WK�Ϸ^��H���P�b1k�v#��1ǔ���Fs�Y�g_h�����X̓�M�j�>c�"p�Ie���w5�r��.M�-��}�|5����&��|=��b�vb�C�m�k*j� 3#�qn��!6��<���ӄE�㣾�<v`ghQ$���h[��ݍ�Iџ:݀�����}��X���� ����m��4 h��2Gޣ�<�	��N�ע�'��J%P>�9���s+5�����+��*����Sj<��{H\k}\G}��[t!&L_x�u'��F��;��I��C:P�S/�2�߈���=�gkfV���+�+(���BiT����`�~��B���I�$qۇH�����ɶY���G���²�v��ڈ	!�~YZ���-ɅA5I�ӫ�Iwr�W~d��N.�.�{}�)���=^��q8�<�k��	���a��ȶU̝2eX�G/k/��/����j�߁y�O�Cto/����^�s���DV+};��C��`�Z��E�Z�*�D�(#(6�m��z7�(��Z��uu֥���I�����Ӎ��d���+��ے�v9+no?{���BYy��$���Y���p5#�>�B[����;�y������@6��yĬ�6��G��:=�:9���=�
�R�=F�����v.gM)�2I@�"��u��/�bki�gع�h�傐�k:�&m�)�uYk�=�u,Ť�X�c>�^ў׼]d�׈a�M��0	I����ōZg#>�SC^���p��
�nI-�^�,�(�ٯ5ϧ��c���,��w:��Y��t�����N؅�p̍�Tl�n���\�$g���3[.9�Rk������ɫ-k�uқ���S�y���ǯ�����'/v��]KYە���3=+�m��9�.?u֍*@���6�I�C1%�ҳA'�^�Np�	�"�T�AԿ`�t��]�Q^��hM�n��~�����ml-QY����{��f��*��峲���ߧXwv֭H�? %��n6�E�¤QtKhF7]f��u�NT��j��>b����|ԧ�.���{VU�^��9���r8$�|���,�J�&�V���PTͫV�V(��ov�����)��hK1sR�v�ޮ/+�Җ�W�V�!�@����G���^��;9f�.�g=WՂ�G [N�gh�t�&���mf�x�l��W�-�M��f�����g��~]l��M��՗�5��rړž4b�n���!l����z��*�nea��)R�����Ă��������>=w�7.�q�O�����dԴ�KU�i���yh�D��j�8Y�{u�3�.��Yz�rخ���b�v��W`��E8I����'m�v��M���K����N6��-�;�k�+�B�AoM�ԧ�������k���9�Jaٮ;	�[���%���V���'O��{^���c��^fd��<']Z���l�u��Fv�����۝{0�/g�M��[&a�vtl�ظ:���k�ŉ�b�w�p����=���T�ãa�ls��:�>V��`�ݗ3�K7Y�{D@����>��� Hda��[xǷ�r��q�2o�:#�)�`�
���6����;�J���x����Hwb�k|�E�mʄ�e�Cl[9�l�8��}����q��St"�q����6�� nN�8ʳ�RDP~Ux�����z������,�@�
ZN���M�G�6�$��t1���C�I���ﺅH��������:x�!���)���uSP�|&�ʙ�fa�We�C�3Y��$t�D�˿����Iwcv0����*�Z0zqUk�u(B���9�.󼧴�"�}�*�s�^3�ӯ݉_Y�!�LR&ب�ńSm:%E��
�����rW>��Hb���AݬΊ,��;��Z�<.T��߄A{*��lP ���cfit9�o{#�kPm�HSI0������qt�I��v�V�"�e�ӫ2]Os0�n	�A��z�8j|�r�G�)
�x����创�y�RobVb�nn?L�(��+�y=���Ҹ��q�tJi�@'H"[gk�7�gZ����k Z��$�ؼ� ���P�z�l͹Kb�]��&����]}���y�Ea���ԝGo�t�U�=l�;L-����GqĲ���N�\ �&�����EL��WW�S�[��љ�Ӻq��p@7D�p�3�I��!���K�H�eA2Fޔ}�e���t�{ğ�l�	�~�(���H^�=s�`�BoWo  ���V��w��f׎zV�{���W�~h�$������:CbUʿ|��V��;�ة��Cܮ�R"���.sp]����R�����^����e�!nZ���m&K*�IW��ѷ��[���ߦ�e��@���z��bF�Gܼ���=K�{1��#��23���hfՀ/�V��O�Z{����M�u7<qu�S���'t���Cx�sZ��o,s{A�������~q'|1](��>����m�o���կ��$��>�M;De�7 ��#K�O}�`�g����S#����E)���7҉�5 ˷��y������rq�|�q�}��]#�j��Y�4_��Ѫ�����ZN���Ӹvb�?xb������i�M��[������ʗj�-�܋��矲��uIw��cf��MY�v�T�ds��(��k�;t�f�_f�[�z2>Qϟܭf�MYx��j����2��U�Ԇ�D���$I�ã��+�b�^���#]���+�r8�g�U�
� �E�i�m��+z9I�q����in��MU�h�]0��.½X��"�s�<,+)�ۓ�^<�X
y���u�R��M�N�@��d�Bl�3�o��-�鯧V����{�*e���A�]05u�ܽ&%���c���n��l�g�,R��An�
�23��q�s��f����\��[���uy���g��N{]*�u%��I�a������������l�L�3����z~����TT����a�[t�S=��C���Krw�K�w��˻�|�]�!+�&rB���~�����;�~������Y]���96g�ME7�*�i'���~�,��߿9KO�'����պ��0��}}�B�]��&�Hd&eH��ԫ�G��w��գG_�1!�U��M�f�j�<ڱ�I/�}ګ�o�����H��I��A�{ս�Y!�l��/�ц�%��`���I�^���xH�\fW��]����.�3Q{�Ԟ�n���e�Ꟶ\�n��v���h�����s�`,
�����{u�NXw'��^	7&+ęQ��q�s�@m����w�>ʕ���xe�1J���t���z?g����g��D�;����>g�FX0�"{�7�v��g�*��e�U8��uT7��o�W!߾??�(�"�pJx����]��)|�j�O~����9$,���\�ߕ�F~�X�\�W^M�1�0��ܚ��1���e6W3�VW��6f���ں�mvk�}�v�R����ϮY�y��5���d.�ޚ�׈2)�$0�m����uOv)?W~������;���u/X�l����o�z�{	A_�I��j$5}Z���v�5K���e�}�}�@d���R��פ���ײ���$v~��9B��|�Y��M�ͤ�����_z�_��^����M{}�(�{:�����MB�IɊ�kĀ���w~�o>OF���H}>�t-��5��g-�3+\#x��k������1{i��زǪP~Z�w蓳�[�>V0A�(#�1$�׷^E����=���u-������ ��~�����ݎ��/��W�'��Ԟ��]b����t�?w���P�:�ߺ"�4\b Њ6ZsL��<��wwyt2�n��O�>T�.���V!z�̻�HoU�F�n�w�����9�� �9���88 �9��9�� �9���88 �8�� 9�\� ��?�s���s�ߜ�� s����pp 9�s��� 9��9�� �9���88 �9�� s��9�� �9��pp 9�r�9�� �9���� s����pp 9�s��88 �9�� s���� 9�~�� 9�g9�� �9��1AY&SY>�k�(ـpP��3'� b2�����&lTUB����B�f٢�V�*9����c*5��L��km6j�ƒ�%KL�4�� ���h�m�ZhRl��[��                                     @       n��m���ޫۙv���t����㷱{n��o'��E��� vz���[y5ޖjsx��v��=��|��v"����K��a� 6��m�O�+j�wz`�i�%�͐�{������hw� �{e2����Ϊ������*�_.C��^;��e'�� ��{�˝=:�S�n���r�y+��m�sݵ�D=h��� ��         ���\�{�;i��y�U׹��g���-�-ם뼲繎� .ֶ���c�3�;�����/7�������v�fn�� �^Λc^s9zim��w��9R�UT�]�j��)R=��=��PP��� ��RJP��kޝ� V��j�ic4��x��.�)�j�����G ���z2(^0k�c��@�_��e 8�PPS�n���ЕH<zt5����         �o��A����*���k@x�
R�:!-O��P*�#� ��	
鹆�y�"@��)�h
������:�T1� �([���&�.3@���E	X��3精�.����m{Nx �{�s.���^��<MtK7�7�w��g;v��v޵���� -v�:�7��z�]���ǖ�y��K��.׍�Z5j�� ( 9�        �u���\N��oWlݶ��w����h��{��m�� f��sǻ�f;���G���]����Kݶ�ۯ���m[�� ��V׷���✇��ݲ:�  �wn_.�e��1x���Uۯ {����ˮ��q���^��ּy�i^��y5�S%�� ��fVټ���������=�v�[^=��iz����Mw:�&�J
��}|         >�ǫ�5�n��^����[����ownӲ�[�{mm� =�m��^^P��ګg�o�Λ�^6���;W������u�� �oVӪ�㛽�ݗ1ӯ�%}�}(z5@k@^㯮X�W֫}�os�|}�:�h�� �+����7�:$(x�tQ��2�ňힷgw��g�\M�� T���O�����S�
>���������J�h�i|<����	�R� 0�L��*   ���%J)��` D�2�SAJ�  ��A5J�h#@OH���� h�O������~����;6-����C)���������v�^M���dC���~�$�J""��Ve�$�IDDlBI$�DB�(I$����8I$�����$�J" Q�DDD/��B��D/���D��__�dȿV�T<e���+k~?c4Z��e�,j6aˑѲ�R�̨Aܱ�t��,-��9I����
2�{KN[���<[)�]^x	��+�����*��xc���a*�W�U��Q�Ǻ�����P�,�H�iUsC��N�4%뒞-T+qnLe��QK�gA�u�B��͆�Q�Q2�Ϳ��U9�S�.\ۀ���A��ٗ4\Ы�Y�8��I�����FLU��a˻�n���e��+	���+i��{��*d�b"�l	��'��4�lJWK](�K�n4�.��2�	���7@�I`�3k������h8�zhD�[�5F����ՙPL��X�6+hQܶB�9t(���A�Y����Ae�8!.�/���ȦU	7���r�a!��5�g0l�¥��SZ�[��,���j�M�*�\����#5�Z���T�o�Zf�5��)%C��X����yWVL�V.#�'�lWu(�v�h�H|d	lO2��'x�]h;���a���tc1*ߕ�C^��j^3q5�k��v���3&g���u�6�0��*����,��+]l��,���S�
�!q�P-$��f:7�bD�5u���be^��ISs$�3p�n����I�R�E��Xd�s^�l�)�Ee ��Œ�������	�<U2�FFI{�Y�6*��]�\4�2^��uV@ktګ��r��a���Z���]��I:X�FU�^P�Y�L��l	���S��Ij"T�N��CTa�^�R�E�N��]�pI�e٤
ߎ` ).e`$U�ʴ+s+P���
im��jyo6P���k��@�/7S�&%��M�X��֖�3N�ub�l��>�Ր��ǮR�wp��k鳴���C���cj���,-En�t��e"鶘�eƞ��E��.X��re+wQe^�qÂ�;zh�;��y�I�����q'CwkKC\8���d�Q�`�y�K7��nn�r�K^������Ѣ����Q�.eN�If�B4�-��-p=�2�ꢆA�`*ne�6�(�c�@�7&��n7�Aۧq����a��D[�E�crQ��F�[���JO\Y�Wf��P�)�Z0�f@o�M�ɹc9�Y�l 6ؐ�-i�y���p��W��x�����W����]��H�i��ܽ�n�C�Ly��B�ct�V�c��91Xc`����r�Hp�p�Ǧ�m�*�-�Of�k6M2kmd�eZÅ�M�91K��?9@�-Kݥl���? f�_�Bʳ�a�;�lt�A�������9�dug ����,2ݲ����ki0J��4,L{y�֓eԧ30�p��v�Y�Ǒ�@���Iy��ZY[R�%�/vF�I�^�4��E�#Nb{�CʢmT6����*m6E�(8��ݶmE�G0.�d�2f�2�s\��3X@�&R��
VU�m3ǂ��hSu �ٖ�F���H����7CLګ�\t�͘�Y��X$$�ֲ�ʑh�]�B,�*�=��V��F�kU	�޺�r�b��2�[T�c-I�"�j�M0eQ���±$�nliĖ�PҧP��AԒ]3z�Q���3�V$���У �P�f�Mޣ��Jݠ����G�e�s2�b
����P'�z�
�l�T�D^ArPg&���T�w�2�e���u��.5
Xbm2��	e���d�� ��ovme�Ŕh���OfIG ���9��+U@�H.�f%��r�n�p�:�yVE8X
@<.�3pۈ
Yy,Y���R��¾�\���ݸ武V\��-�vw0}`�i��CX�,�fi�҄W)DN�+*���ak�CF@�#F^R�q���X;a�(�h�qX��]�7Hr���#0BbÒ�;F�x�`TB³R��.2�*�	��l��s~)�k��4����DL��n�B�����4V� �z���nf�Q�zp����w��F�Wi��ˤ���#R3����j�Kݐ?�,;֓z[�k�ƪܟ%�,�' �֔Up%��(2��b]�ϰfc�"K"]�z����z��*�7��BK�^Zn���a5�GX�m,1D��n���T�ض�f�G�yOS�Xf�6�
�Bƺ�["ur���*���P��,�F�BȬ������7����]�W����2��t$���t0˧��"�VAT6�Q-e�"ʉo�NqY� ������P�÷#k"��K��(b��']��v�5]u�Z��FVT���y���-i��/WȚ�d�ܩ֢H]#HU9=�ӢK���E
��Ξ��b�j�O�/�V+q5/��7�I��ZY�3���[�(!�t���U�{|�v^S�ʪ�]��HW#���r�/�dğQ�V�؎����B�(\#H�:D_=�o	�H!V���v�#*aF�Y�j�7Y�8�G�>�N�X;��;���:;JK�7K7{�VظT(bX��jՙóH	ǂb�gD�,����ˎ�T�h����:ng�O�y{q�3���լ��خ���Zo�-,�C��4n��PE]{�i�B��6K&ܩ8�捜��beCQ@zM�0-��ݗ@(�))
�7�t��	�A'.�R�ҫ�s�m7`�f�Ku��X^�a-MۅL��n�fc+�J�Ȣ�9�-f+ٕ�Y(0s2T���Ax��j,�(?�L�l�G+�H`iE�[��sN10C�/)T4\��I��X$4ܚ�X�U�\9�9��ns,Q�n�Q`j�H�L��xl*Ż����(�ٷb��vA�Wj����n�-ֹPR��ʥ5�&����@�c%�v�H��R���aiJ׌#�e���c���fа�zo#Չ,��SB�D:԰0\À'U��a]�)�ং@����^�%2�CI��r��0�6Ku��l.�3/ F+2m��]�R}��)���^�&���h�b���A1d�hb��C(�)�LP݊�8b[�Ά--�U�b8u��Eݙ�m�4�4��6�YPjɌ۳A��P��M/���I{:�H����J#I��^m1�����sU;v��_n�w��Fu�$�j�;��l�+?%�n�]��@d��уFV����n@: �L����٬^�U+\L��ն�3>���x��#]<�@��N�i��9LRuovmjx���<2��C����C�5p�;I��XΈf���B{�A�jxP�DzLc�2��V�x,G(�bn-�u�#�����d��ը�h;t�ڼ&�U{�N�6�KB �a3PV��f�gF+�#A4Ċe�YD��nSt�.Q��4��\,�rӚ ��Ê;�Օ(e�B+�v�u�Mvn����)�vݥ-���<�0�ޚ&,��f֣*�n[8��[�D4^�A�d�Hf鉇$R��XB��l�ae�[z��zn�b��V�Ͳ�jh3�k�I"�K��㶅L�����LǓq,
H�C�4k0jV��˕(�r��Q֪鴱h�S���P�\{����vorA��u��)q�����ʚ��'H�2���$&����s	l�|��htv�I4�W"?,h�G�s-�E��kH�XEa�V�<J *���OEZQ/��3�/l$�ow^౅%��),��t��8V����6a��悩��<H@RVJ96^V^�,;�*�̒��;�-�Eͷr��L3446��2�� �ș��RkkP�Ab��d/e��Y�IOE��IKEY�7577��9�k��d��1ң�.۹e�����Kh�L��Z�*m'�n��U�]A9h�^��Dü�Y_-�f��b�D��_�jm�y���I� �*رd<F��MB7�v�E�B�)�z�ڄU����[;��{�u%j�-�v��Q�v�Y�ڔ�ɪ��
�YQQq��D�[Z%���ˤ��Q����5{��(F�iP����^�ض1��f�3.h�÷*E�C�b4����}Ȍ�v`x��c������R�Y��4R�]�S&UB/4[��K|�f��i��6S��f'���r�������Em�y�*c��7�<�R�I����50��8��.1�z2^���ȃ��J��*���B\A�2�Ϫ�IU&c��LÅ2��16f�O�Oqöu�y��՛���p�4Av����D�)�K�Px��N��s~��naf
6c�Ʃ��	����.�@�
ŅkV�嚴#�h�H�cBe9qm��5��W��R�%���	J������`4�l7�S��n�.�#�����oHs[��Y���#̌b��:�D���� ӭ+YJ�Sl� В�f�L��&\r����/6��Y���i�#�-��Bx�B���@�Q���0��z�4�Ê�O�T�FGJ��7a�km��d9�S�ذ�U`#4��2�X�P��B)���P�e��o/Djhy��	_hW�^��A(Ф/SC�7�-�%�Q Y��f�`�3$h�%��cF��f�V�m�2��S2�3.�ş
cN^C�GSr�d����0�o0�3wd��V�MjГ��T���[�)2��L\��V�CAD�"���ۺ���Xwl��91۸V� �)U���g2�&���h=�nLٲe��n�n��r��pJJ��,ud��F�7����P�\+)�jG�Rob7��Wh�� �M�(��+^m�*��-���l�:\q�Պ�ݕ��wVJ�=�.���+��KGH3\ā_=�T?�+V6�$�����XE̕m�6����ԭ	3Jĩ)4uc��%c؅��ؖ�UCf;Q�,�S`��J�f�T�-�t�7�^뙡ekR�w6�T�fm�"M�b�Tƕ`���\��-�4�B�(w>w-L��*J:��{��fζ],w�e��7xE}d^���wh!4,;gp$�%�R�&^V�d��8v��-������`��U���-�C�+0�Wyl}%��}d��a��K.{��� a`۱�I!�r�֛CY�wm(v���l���L�42ˋ�{�ec.����ϰc��Ts[ߴ8蠶R[���5RePz����E�-*a���kU�kBS��Z��,ވ���x�m)>ӴSsZ�cZ*Z��v���|��W���dk�fUB��[a��W��fڑ{ ��X�
�n��Q{�h�{����r�u^)�Gdb�cm��;6�4-�n7�K{#�M� �0V3􈗳%3N�Bw{R���u�(��ye�V�>쁼!a
�e�8���KcrС�/ˤ�RJq�V�B�L#&�k"�/���U��j�UM�%�Ĕ$�����Y1�k �o2aH��M�Vd!E���`B<���̊h7gd���f���W���M�ZU=VT��5F�U�Ġ�&�>��{,����Hz�M����v59Zw�ZY����4�	�{	���+p�6�ZY����q�X7DZ2Z�a��:+om�>i#���YQ�em���Y�!*�:��Lq��K����6*�w4��7W�P8�hR���e4@��E{R"�-.�����y���d�
�F��[#wEǓ+,�^��x�#J5&��J%�%
.�M	���v�at�f�t+#�]m#�cei�L5^p�|}�B��&�	�b5X���b��{glk�5�Lk�:�eG��D�M!r�ݷj��f٫²�Z�_���
� ���b�w�ղj:T���X���^��d]Z���ú�͆���R��8I��)=j�Su�B鉴#�K�5�݉�E5��L��r����D�0۬��m�h�E9���M�Kn`f�ѳX�4ö��b�-�z&VZ�e����>������oRjS�p�/T�e��lݲє��ı����]*��T����J���!Ńz�n�N�਩()+��K�t���+�R�"̛ʟc6H�]n2�7�����@7��+ZPFn���Z�iM�ө� 7���A�6�fn�-h�u��J��pfb��K.	��/6]�S.k;�L���mۺ�wh:j����fT[�P=����ʭhf�$�h$�R�y���b�p��]�Q�Ud!C�I��Ħ��]`
�"0i���"eh�eKr��
�B�F��|�i�[���H�V�q
��@�b��1	�"�m���v�ȋ0+���<q]�D^6�#�\�LK�͍2�E]�|�r��*�@�x�Y�8����v��I��M�!1Yr=A��T�`�;�2X�nn�o%M�wp�ݏm19�]f+-=f����|"�$�k�񥖆ԕ�n:Ó0
��fb��2�r���2�6��7n��M���a0Ԍ�����!You�q��=u�`w��#Nc,D���	R( ���/i��L�Q�v���vh�O�&���b�$�[I�BkCF�
���溔�g��/`V������ �RM1�t�u�b�S6��2�	�:i�.;B�������(1�aY�r��C.���N��ѱ�i�A��E��SY�P�/ĕ�1H�{�ߓ�kZ���4u�×{j�jj�;{Wm��B �7�]��Z�����fT�9mS��lgq�#j���Cw��-�Z3�-U^c�KC�2�"�ݳ�X�|,���F26�`�.� ʏe����ie�����&;iq��'��z��iHq��*����*-��E��5J6P;�e������`�S��]㴞8�9)�T(�� L��kM"��i�����QX�(]T��*���%bkJ��Z�y1�쮕.$O.㷛�M"��ke���4����G�G$UG�v�������V�|Z(�X�WE�y��FE���_ڷ��n�$ds+X�v�T���l<�5M�@����a:�q�Iʩ�!�9*������,4R�u($��$	i:U����T�5NմҭU*ʸ�Yl켲�=���tR��Ub���YV����Ye���V�*�UUVڶն��8��j��U��X�kkm;Y�P��l�8=��jU�mm�jZ
���U�������M�i�Z����,mɴ-J���m�A�<���|||���0H��;�kcYZ���Z�����������h��mP6\H��ĸ�Vq��pvڌ&�$�t���{��sҵҶ�v�b�a��5;�(�/u���s;�h�E��;��.Km�=�gq���d���E�w���[�O�|g�kt<��bf�.������S�e;c.5n�<�Ns�����@k�[�m�nZ��U��������v�nl�Z�00�tx��s�^�p%=����㝖�������5�0[K��n�dMծ&Y9�ku���v�� y�7l8���on�:�t����y�mbNvҘ�];cg�}������T��⳶�|���M�Ob��G���S/��i���M㆗����0q/nvn#9���f�s��Z�)ܧk 6E��૥��'\,Yr�]p�Gl)O*�t�؛�:��ĭ�۳�Z�57�k�� �,L��x�Ng.0�#u��<���B��s�f3۫B��w�;���!���|���\T��{u��COn�
��l<�ԦK�Ч<I����Ջ��D�:���;O���ݍ�9��:#AZ.�Óƫ�@n��W�v�a8<�>0���QGB��M�z2�9ui��COm�_7a����gx��t�������x����m	�CuS���C���r�I���m)�����Mm݉`�cc�`{Z��7�n3<M�fN�^�3D��g��m�;u�\lvz*��tgvvݭ{v�M�5�ɰ�sZ�n_nz�su�r�u����An�w[����zܽj݇[N+rv;pN�W��Vw#Ƕ�p�L��s�����Vs=l�N��S`��kt��8���=�VN����l q��㗓=�\M�k\^0�v{#��3ɸ�;�r>��7�9[۶�Z�cmo�ŝ�n�8�^�v��N�sr�x�<��c�kp-/�q���ol��6�����u۱�=q���3�S��P�cq�$�j֭T��ۍ���{�]�/�ok�`�λ1��R���S�������<������ձGEt��6����Wd���y���[�-�i����z���r�ڡݵ\���]��uq��1�z��n�n:9i�nN)r�Z�� �;3n���]!p����[�q��Kbjtd�l��R�.&�%����Y�+�7'��f�)�m��b;!G<�B��Њm��@r�-�;]k��^^ų�m�ۇ��{�����d}�C�E�=�5�n7n,a����Oru�n������:�Wv��m\��V��ݺyn㵣D����Y�v�s6�	R6��?[����o�/	�v�?W=�����w4G�疰An2R�v���X�߯�~7���:�vb�8�MV듷:v��-�GgW=Ȑ�`�%']X��\�zݴ��knlnE9YM����J�Z�$1<�q�OWk�`zܝaH9ga��qݞ��Y�h�Q����[����×p'n�;m�l�����s��Q.F�%�;]�=��ڛm9:˗h6^���7 '=^'�[g��s�v
P�냶%�s�ܽ�y2:-1�i���k&Tnxuu��g;�-瞺�h��&ĖEn%�=u��;���m��{<a�W���[�^>�(��x�v�-\{v�qq&z�͋�`z��3�s#��G�Wk�[��ڷ';�t<e$1��q��]�l�466	�ug����]��R�F�ǧ�8�כ��KV��zu��=c+$8��	����	:�Ln�Ɂ�x�IՌ�{u�Σ��j�g�特�ƕ�ە雔�k�O��qƷx�qu�N�t5n����cӪl��F���qB�+6�v�.�ٚU�+[���0|��m���:��I�N�lr��'=�����Y��0)qͫZON��j��xֺ�Z;�(��6�Mk�n�<���|���nt��(�Z뛲�\ۇP�����z㓝���6�| <z�Y���|�n�v����;stޥz�L��; �d�z����In9N{<�g�a�p�ok�[��3�\Mq��/�\/GGj�R9��bym+��&鷃X�d��u�1��:e��@����Z˜�����;S�v���q�8�����=h��.Į=����u�j�\�%��n6NМ�n����K�2s�N烀�y�y���`9�s���Z�D���p��6ƶ��)�n0��Ʋ�O�)7[�aՊx4Fu��u�ѵ����Z�r�U�hv�G�c�6�]E��z�;�pW����u��<��ͨݚ�}��`�w�l�����k�)��\^jvM�;�7��l7�'�r���;�ۡ�xg��`��\rN1ϜI.����!�u��;;�Ů1��<d2{0�9&��`����/\�����l��n69.3��n]�y]�ٓ�G�s�;���z1�w:��M�qˀ᷷kX�q�觳س��1�뭞�;�{ﯢv�{v��8cQ�J:��uh��:��c۫s���:������׈ɗvw��3=�q���F�䐘b��t�x�l�a�T�]u2G������m���R�u���ہ�m���SˬO]]6-\0Acqh�ۀz��.�˱�I���1f���>��IlN��we�x37e��{ѭ��ۧ]X�쩮yS��3m�n��o&ĜK�h��Xo ���W�����E�^gu=�W08�̽�y��f����8���)�b��,���>i^��s���ہ8kI��<��� �7Ip9����������ۖ�Gy�i�C��1��h��Hi��Ʀ���rvΓ�����MNx��u�g�5�}����n���q�xS.p�l�ˎ�s�gq������y��;�f��8s����@�z��B������pv�;j�Y��{5s��/;���;'A�77�8.Ɍ��pqʀ�ᮗ����۹
�8�gx���Ǻ�Ǟp�vmӹ�����5�7�l9t^���u���f���y����ƣX�gU��;]�cX�b�]�l(�����l����w�Q�!�+�w`ͧ��%����8�����ΰ�^_c\U�-���< A=��gnJ+'k:��4�3Ė,
g����uW�}��xﶽp�g��pt4�KfC���m�n;l�NOn��+��ZL��Q�C��nF��]fC�^ȯr�9ړ[��ۨ!7�wX]؍�S��m��� ��2����썶蹽	��M�����̶��� 0��z:��v�<X8�ѭv6�k֯Ge\���O���wE��v ���]��N�����,h�ۇK�v����j*7�s�ln1��oۄ��r$=W-�����'9�ˮ������6���$���Ϊ�ny99;&#���ʽ�ں��l�u �c[v��#T���a�+��U�K��=������\��4��6vw7<q�������c=�n5Žj�k����x^�q�����M���ݘ�npݜz�*�a�6��;��d'2��[��M���iG�N99Ob�m��ۮ��v7�%����NGv	�Aպ8z 7��[^ݕ�4��Yn܄n:��7N��]��M��a���Ӷ<�cD�:�`ӱ�#�i��+�2��΃n��2m�=�z63�&�g�8�0��vY���.{NuP���v��q��e���ٶݎ�3�n�r��v���:CF2�X������^&j_Iz�=��s�U����Ս��n�W�n��_}�}�՞+ ��Ml�zc 占���d�����d�"�-���D�]��s �8;dT*�Ĺ�����l��W/*�mK�k.4^��y4�v.���v��d�/����ɯa妜�n�8=�)˹�W=>����l�-�mt�v����v���a<\୻�ۡwb�����\r�)7<pn!j3�^���f��͝�kt3eLmd7��F���\F��z�%�t�Y����5��n)^��1��v��u�Z�/�5�͹�z�	�;�ư���<����y�]�j�ڽ��=gc���>���!����v��O$�k��3=�8r+ƞd:��Yԕ��"�	�����g�n�q���9�pm�=lX$�u�K���vv-Gn�y쥻C��ey���#v6;8T��,u���ǷZĶ�ps���R<���lq��n^z��x7���ml�X�׶T��|om�]����8���J�M�l�z�$ok<v��pκS�6W��k��wN�WWX������g6(ܾ��c2�$�<��s���n��n�j:��.���Ȼhz��� p��s�����<\8��N�G	��y96�c=�ԛ�n;��ƣ���OM�z�3\��n1n9{l�nN�2�WN�:��=�x=;v�
k�b��M�����73Ìy*�z��Ick''e�ڳ�C���\�On��ت�b6���c5k%1�ݽ�s�����Y��cq��&�2�vꏎ��O�h�W=c�6�����1�.�2��G �u�����lk|����|ĝ�к9�����r�nIn����<���Z��\E�v�$�q�Ǡ��ˢ�&gMNH�k��\<cv1�av��^��%����:}���<kF�;G.۰���<���]��%͞�L�Ys�������k�{q�F67���PE�\;ql�ٝ����ܼ6ؓ���6�����>�[UƉ@
Y}[��v�:��K^`��s�=���V���[�t�#v��\���hy���S[�h:zN92���MaT��Q�x�F�m����we�t	��K�}��ښ�`�<S�s��@N��)x;n�X�p�
q�2�S��:n��q��(O���~�)1�ц�'��~~���;���6q�y�玶Mz��&�����
q�E˻Jt�z��+m��L�w;v�k$�;wk�h^�g�G!�n��-Ҫ"�*���
��h��IB���J-B��ID(�Q�I$�"Q
I,��?k���m5�<�j��CZP�c�V�u�����bwA���S�n�Ӯg��^ny��pL�`����\{�q�Gc�7 �XmEv�m�3.^C�����n�s�d�:�&���v��=gp�c��t�W�fy�'i۱8��dv����aw�Z�޻L�qP�0vLf�e��[;se��9ݞRNӽ��n&�7�<z��%�{1˄���5�/>�c��]�v�>-�3u�	nڦ�n+^N-�hݎu��r�{Sx�6�h�9���8�C ���=t��mb��z��؛=	��@�F��w�D�7]t�pv�8�0�;�l��st����'ml��8�k�gh��#��Џ3�1tnw[8Ʈ�Qb����xǳmv��[�JԽu���u�U����i$�c����1�c3���玸�=)ۛ$�n�u]�������j�n��+�������<���q�̗n��k�6�Ĝ�˸��x��F���u,q.vz�0���������K��bzz9v�k���+W�����f�vsH귞JZ��9��mS<�=�S�X�����n�˷g/`��b�;��s9�x��y��_=�Rw�o;=�9�A%��76�E8婅�]u7n{vv��n�"�Wjs���mmۮ���9�܀�\qطl6۫v�Ok��;v�UnE��lq��痗��r�-�bm��\!��c�f�����4�s6�n\��fv�f71��H<i�\�b�d��=k(��ت�Bc%������n\8خ���<���Up=4C�ۮ�=���vMN�ݧp[���^g��#�.5�f�c�	��ݻbK� @��vmm����ӽiۇ��{tmy����
��8��4F{Vw���A�ݯmŹE�d�8�K��3��}�-oF���X�n�94��x���z�ӷ^��\-�[v�zr>Hy㭗S�s�/�.95��¼]k��m��gf��w[i93��v�)���e�Ӏm)���SMĕj"�	/�DD(@�D �IBQ��
 $�(��B���$	$� ���H�J!$�Fs�T��i�ڥ4�՚�hh9#�[���S���m��$L�\κ4E�N��C���!� ����&��v�ꅌ�<^�8wfb ����Ϸ�NS\2�x����Y����e)�z����o2�N����3խ����,��v���y�wC��v*Ù��^�-�+�l^�&��ѩ�c�>�mj8��
�q�d�j�۽�[O
�v3��]���n�{o��n�n;eǲs@��,��%!5���RU�������E����[�T�������C'�+qJ'*�k�0�^�����H�X4�`4Pd�̰��s�kf�J+Ƴ�TM@�� �zp�$�L]^�^8~�]����4��b/�!l�#m�2��q6��W-Q��cf\��υ@�e+OUõ�T�������z�O^jV�MU}F_˵H�A�n2�+/m }��z�<N������!���p���K#�V�")+��a��$�0���@�b�̸у��'��J����(�f�-b��qp��.;W]=ޯK.�c;ٻk�
��ѱּ����}f�m�O8�Ȼ4�H�	:I�ԝv�X��h@�W���s�X�m��-�Σ�G�b
0az����Ư���:�7P�ɱ�'NbIR��3A�3k�	�2�U#4�N�H��O��-P�N����D�k��]H(�������Z����X����n�V�[!J��cG�v�f�þ��F�.*��w���L�f��lw&*ߘ��+$&E;�(^е�1�zBp^K�:ł�'��[8�[�g��X�[ Y��U��?&H�H [�o��̷�=Zе����nA���Uz^o\�}<D��W5+J�87��]�"Sӭ�i8�-H�q�g)tY�/'Z�5��㻒U�?>on]��:р�q���߽�x�jђ�b0i�ـa9=��q����_$0q�Q.���גsw;o�k�>�@���b���w��� F�ۭ/q�h�ް��e��J�x���'�H�Nl(�E3����ݝF����>�G�ņD��l<Ӓ�N�@��
D8��&V8���3�������H���n�,�;���kυ�+����)oo��e�@3L��2�M�$�9��}Y��G�N�<��]�H!F�+����%�����t^��#�{���􉽭�����`�m&6wnSg�_l޺8��H4�����c��#�r��!F�����E�j��2������-��N Un��Y {%�s���l:�6l��f���,D�̤{���H�߻�Y�e�m�[��|�M��-k0m)%�Ӳ�]�)��͒>��K�3.�&����I�=�A��h4yח��RZ�`��*u]�$)�۹�@�C�t�(�ܗ&;q�t3\�Mu��xvd���$���!���6L�����&���&�Q�j�T|w��(�]���Q�#�E���;��.�ڒ!�q�3Y;uIy�]�y)_]
�tA:׮�x[�n�;����ȅ�]]�&�!����WI\e�ή�Q}�R��	~Va_%z�8&����)�z��Q���p/F��$�@��~*�wM����t�Ytl�A����/5��@ֲ���-w	�̒�i����I��f�N����o��L"�������I�%��?rZ��ݵ�X�y=�-4Q.���|��w�̴r"�6�rE#�-�Y8� 9�r���_[��X�|�Q{��c��'V)��X�O�a��jf1ˬms��:ֺ�����]��2"��܎������.���P.�n���l�����嬆����.������ZAB�͗	8�g���雎ߵd�Q��}�m�jfx�1b_V^�+��#3��l��[^n�@�Z.��I<��L���a��d��#r����<<�۷��;V�P�KV$<Z�x�6�,�T��	�\J6c�<�pG�I>T?z�݇��=���ry]�43fUS���ݖHcޭ��}q�3��K�޶�ט�h�r��%R7`j�)�z<�Ճ���3ص��bO0�,(�oM�s�t�$C�;�ݽq�O�ד"1;����'z�u��|�"\IBp�t܆K~��A�˰������wI����Z�W�+���1�3�3��h�ޗ3"�痾H�Y�TR��CN�u�q�|އy0!��X�S��I!9����*ߚF��x�y�����VKtYs2�U�sX�dVݸ[=��Ҹ�X5�	5��2�����L�F������ݱ|�z���/�[��FX�΅�Ij�R�=�F% ����N���2��U���������zx�/r��Dq�O^��?[�y���]�}�P�Y"fl��oV�c�~?��l���S���=��{z��qֻd�V3������pcgs;Ζ�ǎ�&���'�7\J�=q���y�	7�.v�P����;f�b֋���n4���G]lV���o[6��t�	z\���l�]�.�th��Ý��;#��.轑���n���6c\��p�9�s��N��7k`��p�6y1m2q]�U�X�ݱ7�|��
���UH����AӜv����W���Ub������$NӲ�@-�G��&n�BQSO뼟��1���rG�^��{ՒjK+�&x���Q��T����š��=$ʎ�nC�p͢8(#I���@��1��IGOfv�vd�v�׾��b+9�Ǯ�U虷S��YE���̋D��7o a��e7��񥂼s��!(ӂH#q��O<=��^*�"�U�'=��4���kav��5��7{{��^�Dњ�N��&8`Y~�D�d����U�t�+�#����@�܇+���NʆW7NA���{w��$�Q�� �I;ͧO��z�A;N=�~;�e�>��})bEb 0م ��Ϫ��x�+mw<��������):��\[<�P&rY� �L7]�Go����p&��:D������<˗m��A�	R�m�uXKp�ےC']B�n���9�v�N���]�Q�T�0�#��ꑺ�욱n�-{�ڷ��a���XA�`y#k��8��''�-K�}I��N/yVK�݅o��������!6�ԛ�ye�r��ؙ9ftnNu}���Y��#m�%�__k�6��d�v�;S���`��맵���Xp�۫�Z���5�w�6'{w��Dg/������\�����e-Kڻׇs��	&�Ĳ_�Z��hƛ(��	8�X��|es�B�?J�ݭ���J	�(�y~��1j�4����Q�{y�"4��H�ND�w,7u���Y�
��ϖ��s�n�dm�����U�c��C��gK��>�K��q�K[��[�
�l/�CB�-���%�pݷ��|u"��&���6��W����G�=���ұ�w��y���[���Hw�j{v+�1m�
y�<�˷<:א�z��غ�8s+�\瀣��c$�Z�r�ʱ����mr�6��Ǭ�D9Ⱥ���噙�-�ķZQ���l�A� ��ප�+OJ�����=b��ؕwE=�X��^꭛V���7QۏzzWn��qf�n4.��t��%��m�x=VhE=�=}G=S.x���o��
ݫ�Q�:��}E��nL�o��G�(#�.�Қ����oMF�`�ȉ��Nک��	�j-Ԥ�h�K��^�6ߠ�����ͬ�Z���ww5M�;%�L�ywxJVY�"�j�E��C���gIo�veAٷ�B;�F�2���*M���QuiZ��UUom��VF^�ܰ�Y����|m�Le����e�wD�pt�'f�f��k�R��_=�趞\"y?{,#���+=4�r���a�����I�-�
�_�q��vR������s�d3��v�m�ї%>:���H)	��	4��{��:��W�Ou�q?=�L}�<�]N�=�xXm6��;Ʃb*����naAesb5Z/8�aI�@`H�g�W�]��!���Z�~�y�G���4���7}n��>3�toO��]�䗪�7CɄo$�]+͝P��S��NF��y��s׏L�@�ço:��Vh=F�ڶSgե�-D���y<�뫄��CtU8T%��J�3K6�lt�!���0�ik-ÿ?v?�W�z��A��^��/��S��6a�p�T�:����ו6�����F>�|Go]��������|�r�5Z����N�X�)#��ܢW�2�uNW`��&�^�¿B�N#T�&"�-8m�i���<��6V��ū�Ϣ�{YWx�Vf� Io��'���=]~بn*C��gԥ��e� ���!$- ��yܙ:'��c%P��<��r��z^�ג��M��{]:*��?������.�3"KU8ҵ�]�V���w_%ַ9��.��#��-�k�Xf���H��:F����[��2/��A���p�J�4�����w�\��6�]�J>�X����~�V!��P���(�B		 $� ������ǳ�gQ�:���O��;�{� �h���GO7��\p]�	s]m:�iѧ0�p�&�5w�b\�e��ܻSsv�"�7�DQJ�x,4����,�e�q����7j�ʉ��'%�ag��$�k.�;��8���:�ev̽���/�����ͿmV��*��(o�hHk���u��3��0�nR��!wrЋ�ցי�{��i��vC��[m.�4���0��Ni0WT�;
z^����MDBv�)t�:p�lm��J�����\��pjx̛[�og��`������)�;�kwc�7f���n:��]��=�]��E�x�ڊq��,�v&#��޹{��@�G.)�9s��F�[u�9�|�]���d��E�0z˯/6��m�:v�� ��N��q�����s`�u,�s��7;��y�����ȹ�;�]��1����l���ء�[��,�L��WjBn�s����+v �g+q	ڶ���gpy�ZEӃtk��/��E&��߷X������o��'y0�CmZ���}êw识?�޹�%bg��zڅ�Z!1�q������a�^�|�W��r̲���2�߉�O֛�zp�+��J����.��͘�C����[15 �5%6&[��8���͌���j��m$��F�1���~�+���x���kϯ�(�E	��wGc��b7������'ʴ�����joy�S1�۾�4��,�������ŝ�e(�n��f��q�S���卙�p�Sd�=��j"�(��a����[��^����Ӳ`k���=g7^��7nnz����J�b���ظy��Zէe�!Vw�P*݌����v�H$�p�ȏ2��n-�=��mԧ"�E�&b^
�T��
u���3pL��x�f8p�M"]*���7w]s��]�k+2� ӇUZ�qu�
W���R���N8���W�j���D�n��Ih�7d��*�75�����6n�X��E6+8��	(jﱹVl�9����!rz�r���/�j�Qu�fA���y�j{��(b�1�J1$�qH�؍��][��X�d2'DmzU��jXM��f� �:���p�:i$���d��b,���$��LG"�T�Kf�ֳ��e���.�F��[���L����g�W^�Ԛ��Y -�Ȯ��j�E��VI��d��
��x��5vsګ]6��=��]����b�֗������<ʻ�A�ܲPV|�C��n@�5Q�wj����Ů�!�;Nt�Y�l6�mGn�t9�ѻ=j㇘^lվ�>�Ic}��ho�������N�ǫI�H���᪦Or�f�S�-�)w�<6�EшZ�B/䋄���P([�=�Ѩ=~Z�0a�mʾBc��u��v��&���(�sB��VJ�����q�"a'�8��U=F��V�i����ey-�������*��Zm?X�/U_X�c�v�Y���R�]c�UڎV�4��n�=nt2�',6�3X�k��A:Co�V �o������� �듩��7~��.�w�[&!ҶX�a}f�X���y���d�:�%p\�O�/3�,�x���n^���s���g�}�����C��q�R�:��+�Y���r���RN�)��F9@�>�7f�n�0=Ѩ�#�j�v����eʷ*H�D��q����τCOZ'u8�p���V�����8�9��:[�u��K�R�����A���ݵ��u�4ql�/2	r���LG���>���z��̋���iWm��%�a�Dj����vjb��}�� �pjbbS�yr=ꗝ��F�r�6\��4))�;2RS�:Eoq�̣A��b;k#�ƞʕ6�T%÷���䔜�h���y^Y&�j	��l�o���B���w2�Uq����X'7.b��\=��|�٥h��v�Ns6��M��+�#�k�ɒ�o�4��`2�`4K�Ӊjy!f�K��o0��I�[�ʮ����u�� �tUN����݊e�3�Z��U�i�����DV�H3On��}��n��cp��tj�\�/����:��-<�-V_e2�:Ų������2U�sw6����j�:�c�3�1��q��iN%���;���NѠ�m_&4uJ[w�����Q���+�q�C��P�R��dVJ�d�K�އ	�Bκ�S������ɉ>W��*.u]��Į�
��w��n��7w�
�C��Κ7w]��߳��[�,��d�S���'��K|jX�G�w1�������u{����/�6�ף��z��U�=���c���k`-6`��
p!~ic1[��BΝkK�wJ���H�k�ϗ�۬,�y'�=���e(k"���)���B��d�8�<6��,uŷ�b냟\�8�+[yz�m"�n�mȒH1��M �ē�>���\�f	�s0a����M�ݿ7iSN�/���4_�:oe{�Z����dU������w2!�"�1�A�4�VL?��=^"�c#���F�?)����9��1F���J䀔Z�kz��[�)�a��R�;T��²a	��N�N��*q���ݖvͯ �8�V��~o�~b�ӣs/@6�|K\�����(2��9AmtQr#�H��K�3+�Ѿ���o��`U�jaЧ^U���Ǽ��7`۫�;x�m�È��%T�gzH��k׈fٽ�|o���8�TTi8����W$�ȳ5���ς��̌����t"�e|N ���nYT�_$+�-��j������Nk�����$Fڀ�
q�FߚT����ևOR#��S�C�g� ��j��Z�-�vp^Ȓ��٣Vmn�n�\K[WW�9
. Z��$�37;f9$�;v�u���ݴ�^$u\�v�o:|�W��v�ٲ(%bg1�H�/���Gׯ�q���S/��~s5h��BLpn�˸ �{�#�,�s���,�(h@��[���)��hM�W^^u.V�˛���1�P���;�2�ۑ߷$]�ļÎx��j��:^`��x�����vQ���S� �)��V\K���]���Ƴ9e��M`=JX��/Dy+ֽ~�9��]�]o%�à�a"��I56��q����2�W�N�����CF�\��"9�^�
�,Qk������(�]Cj�M���RD 1��{+=w�q9��<[�et�R��޽w��<i�3<�Y�_&}'�0�4�iGEf�ܸ^n%�aWVoa2��d� f��w+yN �u2m]&���b��Q:9Ȍ�q�z��R�k���1au>:A0T�ݩ���Wa�܈�<�Q�n�=��t\��Ů˗*�����7q�v��v�N+�W�K��eرgv�'��������ӹ�������n"ss�9���{j��\昹�kh�-��CXw]!���Cq҂m�|U���|�ۣ�xpvy�n���WnvciM��ձ�ͱ�z�������3ݸA\�vB���š�� N��n��cΫ�4�V[�ûz�7<�4:�Q{j��m����Slk�^x�=Q*@�ax�`�}$ڿr#�T�X�t��7fS
�W��e��L����V��L�U�����^mBQ-&��jG�w%ڋ�Gb�\`����[� �F%��a�5c٠�<��z�k��jz�}N���lc�;8
;�rh?��tH�hSa6�����W���|s`�烫GC�W���|qK.v�v�R-6#�=�'B�]�����	D��"[��k{��Q�u3P[Z{h���{�Ijo���v4�Z�[�.��F�����f��|=)����������KqDJHl��������c�%m�YK�NOVD��#֚�Ӭ��.f,��Ì@�;�Cf���	�p�y�%f�n�M���t�%ͭ`֣���<�8�؝�q��<�s��oE�n:{G�Q\f4ڏ���y�a��YI�|.��cr]и"�꽃zC��{�^���AἘ��c�r�R&�8d�FŠh��_�x���r2��>��:"G���p�!�W��yw��&�&��ɾ���a[��iqx��`Ǒj���;_6ە{Yʢۧo���p�@��%W�l��غ^��
}m�{�Lӹ����%x�p�)�(��RE1�9��ZfAd�t��}��;���W�����Y�W&YZ�^I^�t=0w;4�=�ۣZU@��4`�Au�s�{X�嶘���+�q�j<�<糷%�ټ�3(aʻ��[�³��<��^��!/���� 
�,IX���,�o\��<eh��ʐ��j��bƳM�V�[��BןiJ��f�[����qFa:th9�����m�零�!Sr뵳�h�6c��ݵ��y�Ƃe����o���m�\�'=��:h㧙���F�x��	O�?u<�.���x$p�\7�}���؂ق�q�??�P�[ׁ�VFI�a�-iY{l�Sqr�g��Y�+�o����o��Y�n��p���Z����R�N[%��~��Wm2WE�g�J�)���(�m���s]gA� ��]���w^��M#I��M�K�r���[E��	_�� ���4#��/��˼C��Ϋ�����O%��{����p���z�W._	�zV\�oVI2s� ��O�Ф�4S$�gў`��`�+�!�?kX�<����n���\�hz�|��ִaQn�:�捺S��1ʻn�\�\�\d�$D�H܍S�Ԥ���o,�å�Hy-��U�/���Rf�8<�Cn lK��N�کA�����FԐ��A�nV �#��^w4�Hc[;���*����[=��b���p'n-��kj�Zh��a���	W>��V�Q�rK�u��D���V뾅J���2���_ 4��`�
A$���8��yV
g�I�8�a��#t ٗ����])q:mzqb�Hr{I���sA~��Xe�"�Qϛr8pV�l^��}�ܖR�����^�jgx�҆����e�HmVf���Sxv�>q�fe�~ߕo�'A�j�,�Μ�[#n��3~~][���T��1y~f�5O-�6�#��*�_Ͻ�^��mj����%�Y1��ҙ틎�k+,�����W6�0�����Z���l��.2�al��%�N�fԞ�}*S��bp/��*���a�
p��o����uٿ�$t�k$b�{sS�V{Q�I�J#�>u������Z1��y�e+���+>)�Y!�qF�X�'��n3��g�N��$N��\C���#.7���N^c���`�j
%���Xe�zs�=~t�V�����o���
��yiX)\�V��P��)ܺ��P5��PA0��.Hj��Uyz���!\�O:��Y��y�02��Z9��\1M�a!�O������s�iVe���3�qH,$T0��u���������{l�X4K�(N&-=W+y�ɓB����������]y�g�)7	�H+A�\���l9b�:�40.6*�H=0*/T�w�V�:+N�DY�u�zo�fv���3.�-(TF�A'$1�IO�@���us}r �PH�Yw~y5 �z�V��1�+9%և�yߎ��
ͼ^|��tǬ��Ep�����xs2�\�����w�Xo6�ox1*씖hvzs��Q�Z��e8I�u�����7H_��Ny�m�KdH����s���ib�k��ֱ��'k��t�������m�n��u�\�l4�=h��\n�1���}��g��;7gja-��;W�k���;m�n۶�m���r�f茝���Gm�h�^H�h�ۡ���]F��:[��f���;9I�\��ۜq��:�dʹ1�i�<�����u��gd��-`[��۳�)�Nz��Wh۞����]y:�k���0���K!��! 鞻��lY�J�sl�<�dzn��l���"75@��)�k����FAֿ�.���`k��V��U����}]~�{<�>݂��_Nt<Z�H)N(��e�5�0d˚<{�=2t�N�H�D����dh�3�A\3(_5�N_5�з����u]�O4E6�TN���'�/c��fIܙ���hA�n�:�����=3c �ڄ�J�p��-䆕D: 4J�M�d}���̴=�v�ŝY�:�M'˲��=����8︄��^���h��3�8���U#�l�J�B�I2�M�SA�ž2�
˴���gd��&�n��~*7/BȻ�6�9��-����.����X*�W���Zo�rK����	�H�������f�x7B\�k�g��(:x��t���G#l��.8c����z��*����%!�Ƃ-<5�׾5v��XY��Q�֔��÷���o�Ѳ��T�M�	!2�l抴Swdwl�
�]u�ӏ}NwWISQ�X�:�ԉ|�|*��*es������ �uk4�e�6�<��c���cvz��a޾r��ɻ�jNQ��ni�!��}��ᛄ߷�<8n�0�b�q,�r�Z;�y�z����Da�"���~�1�4<�)���O���&�꽾q�g�mn�=�ȳ��h^���-��rL:�Ƙ,8$R#{F4e�jֶ���x�r��ȼf�� ����k-9wBӛv���=�!�|�l<�� ���U�o��/w�[�i��f��a�u��/z���������y1aL��<�U�Z�y��IK��_��y�Qv�U�x9�ݠ� ���S��' nn�۞�)��r[�Ԯx�"z�j�����yv/:�4�rԛc�ʧ��o��ZbM�p˒�~��M�p�9@&�l6��Us޵}�m�s�s�7=S���[՜4�g�׹,�<sN�j�&��9�����uu�a��3	��I������Vmܷ�ġJ�D���U���j��2����,�#���Z��/\��T��]8�m���)@6x��,��j�=�r��tq��V���Ũ��+a~v��On��|E����Kڛ���Sl��p�Y-
U�F��r�S�]{N���IiIvŸ�oz6���#�i"�x�����s]�;��̦�_V|`�̂|PfDKpf/���ֽ��ud��Z��%w�q]#� ë���Yl�-�������%l����X�&c��BjHL��ъ"YWO`�v�p���7V�&�q�x�N�Y��e����ˌ�cpe+.բ��jZ�z��dlFu�S�Ƕ�������<:�y�D(��
v��:��=���Ki3� �LFb)���m�m6�n�z�o�������x�� �p�E�6 X��d�[Y��`VH�*�F,Rλ�e�$E�"��%�"��~7�s6�;���\~��^��s _=�A�Y_,�sW%�2���m���-��I�7�H�1'���-�K	^^������k�d����:�Z�G���NY�>[���-�3�g*�DYN��ܫY�,���<���3xq����[5�[�I��l3�'|N�
쎮f}ͻY�#g.fmV�\/���
��WCQ��Ѥ��!?��ua]���)Ln�����׃�ڍ��ٛ�^��7����\g:�6EO��3��g����=�K%��Rt��L���y\]���sI�Z�7����.1(�}�@�I��~��O�����N�c�:Z�Q�"�+k\����n�N_�� �f9��𕽝j�$F$I��P"6��8�hƜtib�����jJ:�.�&d!���Se�����'�m�om!�z���e�49��J��y���u,:;f]�Bh�M�
u�iH��V�CB��rx;���~2�z�GY{��>�b즊=��<�ՕWӌ�I5/q�	pHKr�	kR����k�.��T~76�v��s�<I�D$-E����\����g�H�^Ù��]xk��2�z�L"�a���,(#n�L<[:�G��x��̰Q��ν�����k�˝��q����,8�P,<�L��X����Խ��k�:��(�l��h�eΎ��#X��:^D	PR�ө�6����n9�z�W)+7��ٜ�o\���y;\��b��>�B$b�2�)�h��U�:E�3A�Hg �bYJ�o�؂w�m����FBb0��ii0m��3���M�w��SLC,�P`Ų������vph�zl�	��5�\�ͼ6t�
&S�Z�����m����u!�{�[�9�7RC��AT�}�����5*,y���v#̻M���fvp㣷��l*d��k`0�MվgZcW�����W&���д)�'?_[�{W�7ԯ��cq��!����f#3�_ݻ�Z2J͆�T�VT�3s��!��}��ל�;����:�Q��`��V�&���ʛf��]�S/g+��yv��c��8R{�f�Wj��+2�qȡ,��F��y�S]��lt���۽��{��@��������̠0�S^�OP�ז�v��Ǳ^�w+��뱡1�F	���xs+ALo�s�\٨�L��rꂊ��2K|![����LG�Ù�)ТC/7ec�ǎ���n��YJ�1�۬�ϋs�,:ܖ/6�e�7���l�d��<2���h"��L���.d���A��xw��o�(3����Aըk��V�F�j���J���r�'`d���[Y�;��]S����ٹXee�[�.f@e�!�"���9�GC��¯���=�1G݈�ǳa���v��.Gw�l�n���yby���#.{L�l�mn�)��V� h1Am��cm2�[j�U�ӭ��nG:��t�zu�����ݞ�=Z�7i
l��.��s�1��6��{t���R��j�;���\n.�7+�7H;n'��غ��Q�:�h�mn��]�&wgn����d����u�,����7BvC�QPrT��;M/�Zx���}��;�����)cb5��{Jv���u�O.���N^:��i����܅��3��N�ks�u�7[���ۓ���vq����]Xx��u�m[v�V��=��Tx۾��6��7Y��:ɫ	��w4k��u�f���~^~�M���`��S��wn$�����hGuêl-��ˊB7\非�nr���݃�R:��\�=i�6����5��$v�.w(uj�=�J����q�I_1��r�n���І�s�p����gd[�2x���6��Rt�z�S�l3{e���v�ɮ���ؤiv��r����T�7��3g�9�#�Q��*y�C�1����#��m�Q�6[�:}������nÔ�6� �=�ǝͻa$;qǜ�}���W;�}��`+�m�Kf��`z�pV�x�_P<�:t�-���>����n{=�$�����+k�R��&훶7[�q�1�qn]�7H�g����Ѹ�v��]klr���{H8�^{v�8G�y�E�nx�:�x�R�q����w@����;�E�\����9�Ŏ�.��K��E�H �r���Ӵ�;�z踥+\|��!c�6��F;jx���އ
�Bq����/nI�y���&�m<�w-�����B�D^�]Q��u���'ir���OcD�s�.�m�1�ol�y�Ξn�ϛ��:v���{�;:�]�g���ڶ����6N{�����O�
��G;�ݰkq�ڲ��u�nf�t����t�l��ö�K��av�]<5�rլ��}�<r��u��5�s�m��8��ܧ�^�n��[lr�WgJ�W�ngv�����wky�;ͻ7���=KlJ�VŚW�����<]����-�a�.Ø�&ޭ��Q�r�9��4m�u�o\uD��.�ǋ���U�s��1��֢��p&�7d:���ظ�#���'�Oo�B�v����e3[��ݍXբ,9,�w���:�r��	��87`7Z<!�ӓ�NN�3ܘ�����.M���ֳ�˲{gllϨ���n��^��9{Gv��6�����	�
f�Y׶�sڸ�^�g��+��\]lA���7�;s�f��o	78f�D�l���$`��N2���w#��7v����e�%�Rj`�ٗ<]Zf�a�t�h�r)x���ڵ���>htdSk�O�ND�.Akzm=��y�dO��68F�0�T̿N�&�J�~X�u���FJ�~j�'wܥ.���ˌ*)��s�
5	��@��� ��5����Vb�'D��5S#+@ɶ������������]O����1��5�=1�
�<�n^uN�bV>ž�VL��N�ZE ���av�a�pގ�}�{�#�Sy�P�*	�R 2�m-E��~
��z�3vчN��Dj���2�fgk�>�ɮ/ܟe��p�iS[��*�yU=��>����"�J}��
�m���ƺ���<���gK��L�Grd8��o[�.���PA+�"q�ai��,�fs��	)'䝧�U���B��΢gfYדv�5˹7����wh���w��%0ۀ�$l��	T6�e�-�=�'���Y��������ډ9��3�Ҁ6�l��|�����[8�cp��}����nĳ(}5�'[ۏ�Ӯ�W��Io(�c��倽�H�f Ky��7a�$����D�)L,MW��F�g�Cs�1�,&�f�_�����������Wg)���T���̧(dj���	�!�&	:W/U�9)=o���"�/�!$i�[���]V,�+�O�-}(��6�%F��=4I�m��A�}؝ǲ�zw-G�o��B&SeSE�BmźN�R}�u9nc)��t'GL��8<2����r<�VA~7�V���ms��:1f��؅���ơp���{^y�V��ӭ������,v�3bq�VwG0<& tE �h II����|3G�}O'�޷�=����@G-�T֬;�׉v*Ծ2�#���ţ��D
5*��".&M�e�i&S2��c]�Ȧ���P�ݞ��bI`e���=2����]���y�=�]��0z��%I��@F̉�����W�AM�r/�od��v�?}TC��y��:�����]�3F.�:P�A�9��ƭlYq\��'�3[\�]�EG�o N��U�s���9�٫��v��*h5��|lֽ��������1��W��|a�0�ƠT���c(�;t��R)����Q˧��b4�`%eCA?�糵C�(���|���C��[�*�� �yqa���6�y�J��[D��F�Dی��:pE@4r�'��s������V0�5;E�6M�>�o"�p�K��W�/I�>ƥ�M��Xh�����=a��n��Yb�����`{!F�V�omu�`m�O����n|��=y�;��3����2��
�v����d|�֔�]���*O+�2�@8"Lh�8׀��nμ-X�pE�$�
[���j��˱#���g�3|�`/5�WA�u�6=7e�z���Wn��BFԳ�}���<��æ�!$xn��m"B���[X���i	e���߸��A��DuP^��=��e|��k��K�u��]"��,��&9l"�42�!��(7�!®�L�ۡ��������ȼ�y�^�x�j�c2S	b�X�{���o�1�SF]A�e;�	7�33,�5VUٗW���i�K[qN�֯��t��R
V�X{/�mm�7&6�u�SN���quy��		l�my!Wo�d�E� &Zl�-����2��SU~�v̹��W�ht����C�u*��C��<��ɵ���ظI����*�[I�H���G-�r�r�{d��Z��&�M�it�%rn�X$9��nt�8��4�-��o���:��z��3�{	�="��Aq���]j Ϯ���0���X9�-j$-k������h?�i�qjo~�=�\o���
����Dp�nԟ{O]-�ØO,>��gq_�U�g��n�O������%�ڦ1pE
��BF�R�ު�3<�_j��,{�HzZ�{Ȼ�(uI�b�c�U����4bo��Srn�z���*�^ ��R�{������ut��ι��Κ�/�2����bZ�_�4s�da,�����)./M���䙧E�wn_�n]\Z3[�M�;��/�(��6s|�J��ٟp��K��}l���*s�T�<���p�k�F{�������cj ��j.Ґ��׸!���Y�Kx�8�JE.��P���M[��|��f�9����m��N�徴�R'&��"1�
�Y�]�x�en,v�N�.�^��� �����,���z�샺v�N�î�D0M��\-��<�ܼ���u/1����'���k�Sn�5��S�d�����ˍq�`;5���]�Xg�wv緻;F3�pn:�,�N  �\�V3� �i;Y{x�=<l<��7I�{A n�	��Gn��ܛ��z{kt���U�8�"�-ɹ�W:�qg1����!�$��G�;es�WA�q�/GQ���b��q�Ή�ڠҒ�������~.�OT�����5h�H1)��Wg����f8&��s���q����)1@
M�JD«��@�N��Հׇ���Wd��XwRP��_�^��
����Ѣ��qM+ܛ5Hl#�C�sD�%�N�p��PM(��H�of��{�ڿ[���$o�Zô̼��).�u"�̭����|/�n��_C��S��\�z�yi�Q��Hܮj5X4z�I��X��c}�N�j���8�kܽT%N����Vo���.e��Ywi��� �$�R�YQ& ��dzo۽�V9�r�:�۳&���83�TǷ/T^F�y��R�T����&vj�H�΄�)�a9v�gO8ގ��u�v���=OW�G��8��ѺS�P�t۶��⸛?��1w��� 7���o�^p����A��e�Z;,#,�7�6�t������<q:'�p�l����e{�A�ID�t	Vz�d�bMW�~��l�.�V"��]��{��l� ���*wv��U�N�/
8�ꅱ��6sZ�C�wF�5�;���{Q^�Ok:ͺɹ6���ԧ�>��s����+{}z�n�@K#���'u����7��e)�[�K�s;qZ[�4�%] �J�XX��(=���+F����tMʛ�S��0=�k��5r����"����^s�T��=T̮�WiD[�$��v��5���{���`�@Z�p��7~�y����mv���+��ōe�1#�
g�燎`���X6`b���M��E71H�%,��R��5ִ8��N���sz��	�P�e�Ҹ�����w��D�e}���ݽ���!��V���"��ڌ�	�ă�u�z�s���a�T�@^aZ�5c�������l���33�v�u���dk*���XWM����}!�[pa�ʵ�Z�^�Y��<[>��L����8*���LEq��U"�wc�~��c���)8����j���$���,�>�o^�^nNE�<���n���[���1�QH-�����i���y�]HZT|��OK/C?e&����F����y�Nخ+5:�U�&fr�	髏	q�ևǳ�i=���Y����>z�M�&{���SVp7���P��+�vݘ��08�,[��n������-/��umz{��[BÐN��[�c"@���<cm�{�{5y�?	�� ��R���o��}��2���`jI^��ē9\��$�Fu]y�rb˲�o>h��L^��c��@�Ӳ	����ę<�u���������	���,BB��՟*#�g�!.J�;h�:w-�Xɋ��Ӣ�E肚��}q<�ڞ���rD'�w�#\�*4N��e��G��z�c��LW/٢㾱�
��QF_ȧ�JOJs�K8֍�9n��Y�Gj'9�7���y"��98���^��ء1V&�$C��z������N2`)��O5ղ�w,�/)=)��� �iz��\�=�EI�36E6^>�@�Ǆ�/)�[�R7��֤��v��-	%�R!~K��v����z%�h2ίvŵ�bݳX)�<gY���-6�]�=XƊ]qp����P{v�e֫��˩|�<8o_I�J��5L�1f���-����q�t�N������J��v��������9�7$�P$0�1mf����S���[�v/�zwݣ�;p�)=�J'�MY�l��<i�{K[��k�P�ԭE�_��h��]�/�	c���@K���f��pgqî�:�(=��[��8��#\l�u͸��Pݍ�*1!�����p����R�W�6c �U���yTo+�3j�{�/���ܷF���MRA�v<��ظ,����&c����d����os���м�o7X<Z�I﷤0����3۽�/w�c�45��t���\io�3lqW������8��h�����f^��8��ͷ������1P��b�d�d�^k����5�O������pϏPЦ�e$�i�W��ݮ���~M��ۭ���n���݄��B�U��炛�;ޞ!��zsu�i��+۩����]�Ɛ�`$�D�w���x����w��^`)k'����=Ƣy��3,�h��8�����-��3:,U��m5��˽˫�-!���1a8�e��v*J� N�
�o����pr��Z/�zV74�t���Xm��/6彴�aV�ۍD�1�/h�[S!�����۞Sm�8}9xSt�nCu@�.���sZ��.yxtA�%;��j�͍��ug���뵠��T<�<�ڎ�`���m�R���ۑ��t�9mʷu�<�V��q���Y�N��I�֎u�"kk��v�S�Z�Lng�P�I�.{�mX�݂5ۙr��x}.���x����@�]uq6�u�v�kSnι��.��J�)�M�׭s�;.��m竎˟n��Z/0q���M�˽y�+=?n�g}��QA��x[8j_4��}L+��[��-�J�dM��"�b��9���b� ����o��ͥ�Bfg����G2z8�[�d�n`V*tL2;�pe��}^�`0i�-E�f�`��j-i��$���B�O
#���2����8���d(��IMi��/�rJK˦��`��E�,���K��^��-���iJ0Z&8l޺�U��֝�̋�����t��^��۵x��������CVv�=�6�@�����Ś���UA��3�ĂRHdq� ��j#1�Pl~�Wm���%c�J�VK�s2�N��ww�r=�7��.�YS΁q�@�˦���W�GlZOK�b�\m����j ���Y����܍�nL��z��v�N}q!�D�����i��l�V��s?qj��x��F	~�wy���X2]d�U��z�Y˸Ԭm�&�v��zC�h�h�Ph�nA�5�A���r�>�8�j���b0#T�����:��t�J��*�C{����`��[�aI��kz��3����c�y��؀���f�����y�oAN����/o���ϭ��T6��9I�72��Wa3�A�q�3ȿ�f\P��{��R]N���&
y��e��ٝ��F'Q��>n]7�s|�Ƅ#����0\�!Fz{��cl'���6�P�!��]ZGt�̳���m=�)Y������Կ��d�r����B�aVC��9=����Ʃ^�w*Ɋ@�^�m1|D�Rnn�r�������x���Kb�����
�y�t���E�t�m�s_m�,�D�N5Q�E~�P.~��Q� J^m�}ߟ��~�?�� yt�k-a�v睗G#������d��Ť��Ů�[q�I]v��aΐ%����h%b7u�2+�/?�n���ط�Gf��44���S�#*zj���kk�~�:٤�LX;����k,������?H�����v�2�x��h��4�=�S ��Q�7׬���9���١`��D�����ꕜ��H�"�:F]�}��U4J 'E0R��d�+Z^~�����W�d=���r��P���K_]��ó��I�&�b(�sD���%�N����Ĥ|�v�Ǯ�=�x�K�����K��R�x��8��΢*c[�Ոdg���`��x/D}rĴ[����?�9}�sӆK��6��*+7+�KB\J��^���0�S����3M���g�^��C�8T�9{��]J��[ߎ��6%){<Qn����ׄ�W�֜�R��"2d4����:B"���9�DƄ���Lס:�hEI��OA��1�[Kd�����$�B��J������n�g��+n�H>�W���E���6-�U�iÇ.]K��&����J/�)��x1CZ>�a;�>,���
�eK�׼}}w��|6��z*Ŷ@L�F9�_KQ�cYF���Y
�/N��m�0�$�nl)����`w��{����O�{6V��huu;pt�Wuj����pP���ɺ;��r`�3�5	��s6p�F2�����yQ(�FvğB���s�퉘1w@g���+�A�xT۾�TS���-��Z�[	;_7�Cζ�:~a8\2��� Him s�,��6�Kc��M�P��tj�oҒ�h�W>����ou�j��M
�mC�!.垴s�7g}��Mf8�^�+5G���WJd�N�^f>ǂS���h�v��eX:���69��y���׫�狸��G��$"b��bi,z����n��Z�d��Mb���m)[�p�'��	0kk�9B��#�	Y�����S���.���M�P�C��R2��D�-��2D�O��WB�L��L�P���d���nZ���ц��Sٌ�++��Y�{�s��X�3���ä�=�k���Д�$���l����L�-�#n����G
��>�����b�3E_s\��E޵�fR[������ִ��B�ySrժ#�I"��mJ�\��7�s�<Jw�LR �!H�[/�}�n�C��5º=k.ƙ��iB�������s���,��Z2����r�pa�Pugezǝ̼��f;�Z�ۨ'��:��旘���_S�&|�^��.|_ح.q��sݝ��D���]��;]:��&��i��읥���_��_gnˆ��˗{��k�Y�*��#�`�!������R�4��]*#�߶�ր�1c�M<Eܹj�uE���0TB�D�RBk�~��g!�v&_�~
�?'�����lK8�M4!s�}�μ�+�N:.[�*.�^?��.����f�4�XY��$.Q�qZ������_��Y�]�|3W��<�}��ȰDA9#���	iT�C��*�?���Hຈ�}p��S�~��Zľ3-���3t�h����;��4t�����C󌞉t�ʮAYtҾ:!r��M� 4�Bh~�:�ʧ7� �rFqD';CL �(��~����^���X�ƾ��>X�@w��.a�d"�U�b�0�(�
q�YB�Q�}ټ"�#��(R+�x�˳�M�߶�h������K`�'K>X�2�J��[ �5=�LoʷԄ���{սQbo=���4K�o4Z8f&bg�N�_&�z�H�*�$�Bb�~��ad��v9/�A:�L�2j�B��t�R*�J�X����ߵXC8)|jzi$��{�4��y�ݹ�jx�X��}V_۸��#/�V	i�%{^�Af�q���ٴ�n�"�f.4��.#
4L���y���+��D�vԈp�>�=��ߞB]�("�c�Zd���IG;�/f��<�XX<�+�z�L���<s����Q������<�6@�k�u�W�gH� T���ʧ�2ꦽ��P�����h�'o�:돬�qZ��y��x��
�KJ���3y�k���]M��ֽ�bXG�j�G鿳Ha���F�_�Oΐ��LT��K,Q�����ت��h;��X����@�-��H/����i迭�᝞�ƴ�*(8a�^���k���AQ�`�7R�B��}���p����ͧ��Y!Z����V�~�mRd�4�\�O!t]4TG³�Th�}Ş!�<�
eГ(�T��9���g*,�sg�=��tS�]8aD}���/�E�cº�Y�e�T�������\8$Ϋq�-p�k}��}T�8�ϢN
�x��1)|!-�Y�����G V}��z�$Ä'N��-��t��RG�ﾛ�-#����:p��������fx1)+�L'y�o��h������fLxV/��/�uo���=Bj��ךӠ)9��4K��J�8~��k�9q�̦ �����
�{w'V2���t��>�XF�£¾&�L�+%����$��8B��㥋@,x%h2��aB�zX�u\²�_ @����wb��j�3���S��Y��M��o$��#��}�*(UI�z*I��y����! CQK��y𙲭���IN����������e۵�ˌ�v��|v:�\�9yy���n�D��u`1m��e�j�N�.�"<����qj��:q�*ɳ��5�Ͼ@�v� ۜ6���vk�"�m��]�u��l �lu��gv5c�3n��_a-vn�Au�5؃b���D7e�>N(�03<�����T'm�a���p-�.,n�Q���:���_/+����y��v.L��q[����78��\�s�j��N��{�q�N+����G`Y�N��n����#�M�uUU�~�)��Oe���~�w����k��(�$�2�IC��G�'zZZV�$PŻR��i�]/�︯Eg���r�_�92�Q
<G��6B��E4�k���f�}!^8�,V}�a�*?��E!8�A�㡄��4K~�"ĳ]N|������s�{�N�{:���=���F"J��S��9�.g²>SI��f�Z�(ξ����!H�9\�p_s��m8��h>�/�(:Э�g����E�:���L�(5,7"φ��y��I�BD�����l�?_iQ$+H��->���q��-�{0�:��C��w��Z5�\�t!d�4�]'����)��n�Z�i�H�s3���ӄJ�d�R&9���_1]7��L���ƓC�����?�䮇�g�S�8��]�+��^#��E7�=�n��'�M�ek�E�_
�	�	��-+ǧ�vH��!���7}�)�� o�Ջ�S8%��*q�>�L�}���'@j"��|4�hm���@d.z�5��~�J�y�"��Q*���_mfw���fs�!R�
�Ӆ�����
]��V�N�����E�U]�0X/�w�q��n��R�Q"�S�ew{g����~�c[BI�^C�@�I��<v7��:��@룃\˼�oliȕcnp]�w6j�T�/	�*4V&�%�ڢ������i)!{�0����ߵdX�\)�*!e8^����Gv�}M�{3�G��~�ab�H����W��=��p���6$O��\��1"�>�Im&X���1i#���!Y�&�hJi�|�V���*��9��H?����to7ct=���j#0��s%��k(p� h���d�Sp6XN���QkM�D��E�̹|�o]�sjg�A���+�"R�y��:q^j�n���=P���*�0Sm�"˯}7��+>�i�|݋K$߃y��u��Z.���o���x>��tp6�[\����ҶT�9�������0�!� a�]�Չh
��%ß��aÜq�O>.E�Z��#���޹̿�o����$-4�9g6դ�=��޹R.53"eX/�e�W}ʅdxRG���b4��T-�(�����]#:�E��_n���7sɟ7�$c̾�X�R�E	��a����	h�E�j&���J�SwZ%��%rҟ��p��L�
�߾����J�D�G3��!V�{�ΙQ�,���8s����?�'�`����*nLZG���}ᇪsO�|�ߩ���g��n?��T6X��Q�+;��w��Ջ�A�:*!U:�Q_���b�Zo&��e4�ٽ������sL.��I���J8%�hSnr�/p����q����9�^���ٌݧ��	�S47SO��>#�P��>��iO3n��.��`�x@P�R]�}�b�޵҅�S��H��Ea��NV�7 ����_�v�3mb_Y�*@^�"�|�����]�
I:vʘR+��4��ώ���� �*F�m�G�����?"3?~r����m��\8!{�z���^;>�U.��}9H�NE���
Ͼ�)P���|X�&pVD��/�;!l����i�'~���8����C$�݈���[a��E�ܖ�(���%g�J�7m���F�!�Hľu)q,,G~9ό�tO�P�c��B߿M���H*A�r�� ���{֧�|N�"�j�|���۩����bн����B}��	��S�ܬU$t2��K �k�W��~��~�^��b�2�.	�%�N�3�穚 F�s��1:P����QmI�h"�xn�r�J\�"FH�p��i~f������M8o���;��� G޸�� M����<���-�,�
��v�f����~ǟ`�JC�`�k�����|i���Ut�{�p���V�- !2�`�A`�r��0Bq�"j"�P�F�F�W"�Qv"���mK��J���t�",�$�o9�򹭵V?}/�ns굄مE���Bҹ��;{��mx1��4Xw�q��S�B\�?��t���	0�L�l�>������'-���2a��FR�8vA37k��6r �.��듔x:�]z��^�6v��������ͺ=�J�4�<��M�Ä1H�=���o�R<��7	� ��E�(�J}�+I��:��7����~������f���*��n��<�V�Y��ȡY��'�����w>p�i.G%���@d.0J������nq��_W��U�VB���>櫅9��F���������p�V&I_l�dY�r*"j}��b_#�����#�#���y��z9��s(��~�������=�Ϲ��[o~g���7:0��,�}3�)Q���Ș��q]	n��%F���[n�]:F9���}6�-��Bfۀ�ix����i�n0)��Z䯇��7�(�QƤ�?��P��"��c�i�j�A����!�9����Di�ӎ�"\Ʀ�1�E����.=`x��{~
��ay��: Ťa`�
�7xfg���n�������v�	�m�nXa9��tdr� =�te�֞ѧouݨ:�"/��[bq�QlU�69����㟿�.���:,#�tV4%���φ7:ۖ�U)��q�4��r��xC,7%*�+���W����B(�����弛�>����nn�_Dqש2�q��3��.�$��z�@][ �XD��Y�-U�Й��T��>����4���u?|����~s�Nw�\곂\�۶�&��m�Y�-��(�j#p�������x�g�sN�T�x^GHD&Bb��v���!h�5�2F���L�,�ړ��y�ķ���z�Ţg�d�!a��u�����O̔+�����|ÂL�*De���\��s�,-�R@&a`+��=��-�$�&�U9Y�;3���CPAڇ���8Ssd~�JT��
�
�&��3��{�ⅽk�J$�$J��!�{�z-3]��9>T�I.W�9���u}�g\�eXv���������V&G>��g�%�l��ƇSS���ڕbdXkJ�>�ڭ`���>��w�pg��mp��JTYϾ�B|����y��|5�K���g9[����6x�[XJ,J�!W�}�b�q�ӈXt�	��"�_�G�i�EF$pe	im��X�V	���S+�{����I���I7��$C�X'Hd~?8����o��M�Uxz��戃�I�T ��$��{�h���L�hX<\��bG�����YS�;$,���V/�0��5���0!_}���TM�NI�����4��[谡P߱���g��Õ�z ��1M6Uq�	X���j�ؚZN����ۊ��>�_cVH��%�Z���I-����*W���k�tK�e}��8�,�guk>cսۦNm����Sypy�K�Y�جi�M#�]�.�654vԤo4G�v����3��}Ҳ��s9Ovb胻�hj]���>_�x�d�������]�v�ܷ�P4R�q��V��ڑ{̍��{.ݰn�[*�c;#�rmگ�/k�L&�Ƞ�m�����X�\�@����������kɁyt�w6��Z+K�]m�gv�Tsm��n0�8���8a6sr�Ǡ8Ÿ���(y�t��ۍI��v�pւ�uF�<n�!v؉�+�oKc7 tu�qg�n��ے�>w���$񌬫�����ݹx�77k��<���7T�J��E��i��8_K�����p�\�qD.[��j��"8O�V�+8/+"���J�#E]��V�3������=o����,^>ㆋ!Q.wsKJ�k�%��F�������g�G�LҢ�*��*h���qi41�Y�$P�-:c�ڮ�E�Ζ"V{>��e�F�_�������s�w��S��+H��,��B%�{�X�/E��we�'���-�!��ס�CQ�Pqj���~x��p����i.hFA�*G4�pV2;���@�}�O���X�6w[��X2/���b�b����i�����X�����>�hS����o�ܟ���z�0��Xrw\X�_7���_r�,�p��)$����!��i���,8ڒd:~��"�D�������A�`ܣ��CC�#\� �t�,��n�[V&G�f�&ԊK���@%uЙ_r���XtJK����/�缟��%��s^&F�$A�d_&�*:C"�tc�m��e��E"�ѡh��o��I�N�����q`��O��0��E�Yk�o��o#�s�����>mcL�洳x�i�rF�o&�����]a�5B�r"�z�X+F���k��<G��oT a���~��������`�o�݇Kχ%	p�ٹ���0%�-�ZG%ɗ�����;�����R�L���^4Lߚ��Y�Qn�ƿ�Z]8.�ם�tJ�ĤF�}ϹW/��aws��-���.l���C=ûnk�H䐸;�\!�B�Y�t�Z@'��,�M����|u͢�p�	b4���Mj�*0�5�6��.l�����3�XF��F���X�׎�1��w����f�=�^vN�N��\�VRH�`u���
mok���l`AK�ђ�[�{�1�����/��b�p�U�����vma��&�'֤�j�u�R�7�w9�LX��n�
ę4�/��Z��£E$z�W{�y1N� i�Y�(���ѭ�"�"n 䒀��Y��#i L {�����#Ege�M��j�w��Ы���_ՅG�!L{�� |+oX������Q�9��kL��w�1����f@V/w��p���ٸ�ac�b�L����Fbi��B�qP��:Fy?��y+쯏:��:��e.��\-�"��{�Jc�}��h��b��M�+�{�#���{�^�Z�S�|���';Y����K=}�k�7�/���q�U���Tz=�%��%S�]Hꍏ_?��_)i[.,�O����X/�C���V��MU�֗�~?�W���z^B}�����{�a
���?v��A���k!��}T�߱���ü=<)뎋5��q}ۥ�+e��7�Jut&M*]�3����tGv��;$mg���\�ݏ<ݷnևv��=���nC��.n���w��p��q�Y�d�0N\}Mo+~��pO��B��!¡YB��k�5s�*Eb��V+"P�
�K�>�-+�Q��#�>�_)b�p�H�ϫ�V�T2�d�?c�0�����3��@����sO��訟5$2J4_KO�k���E��\��2��������3�����.(p�N�H���6��ϋ�>4�!��s��@9��7zW��P��4�M�	��H�D~����ġl���*u4e	iGK!PŢd+��~v�.���,L�bkE�	�Q��Η�������U�����mII0��٤���G��ޭy���0����tS�WSѧ��� �{[Y�	+5,�t�-}���LqcPVܬ��m����d->:E�0I��7~��4��MCy1�vV�H���뉆�Ia)gE���E&��x�����u�?��|��yem�� `����d*ǅS?r�p@k��4�S�k�*F}��8����������\�v�}*��oE'E\���� �Z�
ń�d���̿�)aE0��54\-#��8*!H�v癹�#`]{�^^�¡g�������{Z�(U��	a*(B>,�Y���k�ڹ�8X)e9#m�j�����'g��g2pJ�`�BR�ü����M!����0��e�Z�'ƍ.���`:�J�]yٸʙ�w=F*����?G�����箎����[���q�������� �n'D�����ŤՒ�_n�oDa���>C����<D�7!tr�����p���~�B6��E��%�7��_\�%��RA-U5(���ab�	Em�`a����Fδ0T�	H��s�F�����׍�ã)!�J8����r%Z�r�-�r�3���P���m|�F%��gEd�3L/r��X.���n��ݳw�1����9�9�[
�)�T2h	�7����+��Cb�yҷ񿖋��V- ���Z`��>������p�}مGm�y�����i���P�#��W��im��>KdP�^�s��>����q�%��	���x�g���L��2��T\`&pTt�,�O���NԼ����΀�X���G�~��0�WZ�E�ﺮ_T��n7�X��!e���,H��g��F��x`�R"�kߌ�����׵��7�7�m [����t.���um��N�-�V��ήN��	����	��^C�`��>�.x��B�7|Z�c��SW*��v~��`�0گ_�|ߓ��F8ꪟ!t��D�]2�VS���ۿ=�ݎU*����Շ�]��U�k�Cм�k�O*8)�'��J��^�ő� ���si�d��.)�I���<Z/�}RЎ�8�
`��f��ﾞz_,?������m�{�ln��!u��tv-vݺ�XP��ܼn�t���[ڵ�.���ι�=�������x���E(�۲0d.��+�ƥ	��
�еc��|���iq��DH���zS!X*|!�����f��UQwނ�x��Um;k�P��k��\�$JHRp�x5���|�i�(�Ժ����*0�,�Fq���+��k�1�]�Z��x�:��t�aG���~w
�ن)�"����^#+~ٸ���τ�T�	�iӏ}Ot��i
�H��D��5��]��
���h�hF�!�i�䆾�f �X��x�W�9iS���ߦ����&QD	2Dof�}6�m��"J"���ɯ�?qd�^�4�;vZ]��Ax�3m�c�{�J��斷��-/�8S"�?\C-:B]_+?�a|��D�D�X�����"L���W��wN�����}>�&�I4L�X��!z������]�M@jP�#G�l]�<~��!96�b�[U3�4Xfu��0N��|_��_܎��_�zQ?��|�^c�~T�4@�?Z9!'4
n8��#
$�i�$�N$�W>^�|\�����*��\a
�<���k��Gy��%}�V��_>�fJ"�>�E�/���vY��e�bG���a�y���	�*�K	2�$�����I�/l�����FE�Ca���~�V�"�I]��Tg'�rVhי{Gh�7ݖ���2�Ԭ�y�s(�k�v1�Yf}Ӫ������H0���vn=5w��A6%��r�Q�3�s�t�+,;�m�j�]YU�K]�Y�qְ 8538�v���Z%V#�Ir�$�>� �~���7�\���ͣE<��v���Q�V�>��X}����㢻S㉌�,�X+b��®�^�L-�s�K�X�{A�MY��[ʕ}��M��}{V�*��q�T���fԸM�1��f�'%]r5P�h�����`N�0Sw˲�"�+oDs)���.9%=��wE�h;��owZ��+㏳����"�\pv�p��:d�6oh4��bj��Gjv�%C+Q��Q�ea�4iO+�=���9�{�1v�ʷ��u��t�G��W��3��N�V�4O};o�U�o(w.���B����q�|3�.�c�u���&�գ�;�ϖ��
�Lm �9;5n<�}W|f�����pܝ����Jk�H��߄�h�����U�˝�@��
��ڏi�R��7Q53��]#e�����ތJ4���Yk/i��+.�-��so&Q;�Z�Ё��{�t,����ec�VS�V��u�M_e��F;�lf�;�ٲ[���Z���rv�υ�Y����]��;�k�::ȪbZ�i"��
�'n6���8��s;(�8c�8�;y�Ey�sR�J�U�=����aea�ю�X.��ƃo�Gl�R��5��ʬ�f�+�f9��j[ic��Ҧ��m�6���_�g]���^��fv*pu`�u�ol��lZ䎍���'#���9}�Y;F�tvB�ޮ�n��׭�j�\��)o!���[a�c�l�<�{T%�x�EL�,zJm��u���d��k��WM���.��n����''U9�ƷQ��u�Ȳ��^� �nCX�U���,���/��z��Z-gn���H6�;/�A�m�;���v��ɲ����h��s�S�oI��9�a�gn�h.��[j�� ٷO�	��[���E���:�^\^M���m�v s�{r=��t�S���^ְf�㬛�����{*t\���r�S�{�ǌ���v��y�۩=�9[�>H�n���z��洷N��ی�����q�/vy��m��=b���+D��S�q
�%7<s���ٝ/��8Q���.��V��;fb���5���&�vհ��u/8U�gi�C�H�+��g����mvۍњ�t����p\\���U���q�.!�(J�gY�u��p�c����v �E���&�톇MsН�[���+�8痌\�prf��q�+�"�� �Uob⌧�u=`��y��Փ��6��EI�I�l��`×��gEa�e�v箵)�\�br��W1dN��^�Mc�3!������@� >���v�8�{.N����u�x��=��o0�6Y��8}�n�\ŷsy��f��x��n�їnY��1���ۏo�03�
�;�ss�ͧ�=u�iqo�6��\�7�h���g	����GF�wOHn��{�nY�u�Mx㗣ō�箹me��xlʝƥ9x#vۜp�u���ݸ�u�U@�u�7N5���V�͎kt�t <�a���(� l��Y��[f���k&�"س�v�9�c�p)��m&nxu�=(cl���0����s�e9������x���% /+s��B����vvݣ��!�8e�6�<G;ƹ��<��ƹ��B��Ȼ�l�dwC�����[n�CZAp;#��#�<ku�r�۞%����x��n8��n ^'v�uBn�mE]>�s��Vة�V��q��n1S�cnݪ��mO7g�,�F�V�rӮ����e]�W+��7\<�F�޹��g<s��;$����s��OOcns=�ݻWF4���{aq�d�+�u◟n�8]toj{b6�����V�4�\t�N�(�^$c�Px�wM(�mƇS�n��n��y��n�i�4b����������#���]0�iX���%�_�����%��m�������މ_�J�,���V$/��϶n0�����Y����W�Qr��_D�K�dj�w��vfx�\��$T*$��"�}|�(�|�E�(&p��;�ҐG���F��;��t���ɺϏ��ܮ����_QϹ���X�����t���D*�P�^x��1,81����
�e
Ea��q^ �����Ի�GQ��H�Y
��po�q�>R4$�G�A$�_mcB�2�F%��Ͼ��
��QQI����|�⾉z��V%�|���sWd�����b��Y�s���!�9i�x�4��OH�)��w���N�Hέ����y|�
��;��9[ :�`�9�1+4�gF��p����?������~!Q�]��Ä��!Wޫ��H͗�y��Z#I EKR���2����<��ĊH��jO����+����B����+�E�^>�dX�h!l�d�ԁ�Cj�������<�*����TI���������i�9�ڀL\��?i�nr�;ί���p����D��� �f�ٛ�it�4�)�AE�N}��qj�q�p�wf�����9+��}��.6�V����:,�l���t�qۺ�!�A����C��V.i��-v�5O�A���
ȡQ��Qd+�Ϫֈ4G�ED&���n��M�
�¢宋%²g'�OW��+�p�O���Y�	�c�d&���zM Q��n�d����-�`#�V0������!.
@��V|%�p�5�kR�Z��Bۿ�n
�� �ƯJ��-�y�t�9�K5�6'}���7c,���ܷ��*��ق_�k���v�2�R@�4���S�����^��8_'[�+��+�W���)(\땘�"&���TG�o��H�ŗn�-&Y�������c�p�WϽ۫�.�~��U�*��މg��"��H7$v?F�$�˔q���w�ʡ!�/��U���T�!���P��쵅}��ip5�u�c��=����֥�ĈVr`~ܫ�xA!�8*<��v�ٜj��˟w'N�*��0���`��j%_�4�Q��XS���j�:pL�!9M�:N����A҈fK�+�+ZN_.h
!Y	���M��NB��j1���4"�@����$�(RUlĖ�T�}��R�w�����U�2�j#�U��i�j����a��9ShR�i���D���(��b�#�C�{M���.�T���r�}�O���Z����ww����VI�?5�*���+Va~�>�TH��h�*Z�D��4�����XEcT,������)p��"���M�	T04�f�:����s�vc%���8��Ѻ�n\�M�Z��R���N��кBd.K��eˎ��_;RF"P�9.8*,�|{����y�ԉ`�������S�_�őE���������ad��@@Z_",M�·��8Cq���?�Y"\Ul�o�V������������;.�n�H���ﺮ8p�����}�����A���k����@����u��%uﾛK�}!��}�c	U��W>�mR�!\��5v�}su��<�H�"������[*���nh�"|�T. ����<�b��8_�q�Ex>����2b�P���l���tgV~`�����
�_�Ϸ���˴�1o�'�=<"9�֠]ӏ2L��K)�룲�wq�&|��S��3��ϕ9.�����gag᧐lB-;�iQ�P�ާ���&8)[��+�D>>	{�+����yV�][T�K�(j�7*�4�W�Q$���<W�������uq�뛅Æ|�L"ů�TH�_o*�f�u�ia���/��+3�)�g�7�-Z!���$�~iX��3�ަ��;����l��8~�a�1ؾ<e5?D����ꔷ5V�pR�tҒ�T�LR��d��}xe x��<F���)�k��ߚ}�p�)\/�q�ő�Y)��.Wܲֈ8�):��(Z.H��}�k0�����������C)����m~��.Q��F�Վ:�\�ev�3���8�1^�O i��r5�<�5ni[�G]����߇ͯs#>�M��H[�~��Ã2Z�Da�p�Ss1��x�pمDi~��r'��~��
�h�~ړ1�B_y��+��z٢�8s�o��|X\���Ʌ��{T�Q�\�3��0���L��Zn�d`�8��d�p��kE��V���Ց��?L�Y��W����&p�"
�7��k|��vb���ఌO�.ry�����'wz�1}Ƽ#_�}E��_�#��y��ٹ��������?�C� !��߾!�m|�q"�\#I5'u���xi`� ]�����h�vm��Em)'2�T�V}�8��g��I���^,#�)츠w�yǉwH�Y
E���_����ċw�m}wA�~������,� �7|4������g������@�����e#����Ʈ�(V3�U`����2�W���� �JF�4�p%4�=2D�>ⴵǢVE�S��h����������p��i/WlIw.��qjt��#�g����7��:ڷD-I����h;͜F��K�9�.���;o;A���9y����N���p�Raw>������];R4	�iSuN֖-$_�1�����H��+�� �Z|�ғXD�H��{闦_o�G{����g;ߪ(ZP��Aw�ǅ��~�X*���,Xx�(dYd+���hi至
i��.��F���M���#`���qu�<��c���yj�۬����/mӚ+����]6���A.���T�=�T�D_O{j���zHݒ��~3�;�ƴR)(�Jtp�Y߹��W���¥�"� $�@�n� U���B�?V����S�L�Є��. :@M�u��}�Z��.�.NL+"�j�Uʭ��&]C
�2�F%Y�(�B��1Q�~��>��1E_|Ŗߟ�M�@*#�لȑv��7{مb��ma}S+����F��T -�2R���4�s�;]$\��Y&n���6�??a r��0�CK�h�/�3i\�G%Z\'\_+�Zii=iX���u��ϖ���!?n;xꐄY���/�;�
��ݑ�ӛ�|H��IBWý�_&7�O�Ʌc���TEy��w�Uǀ�<U��.�P+#�l�'J�S%)%��H��L�ϱ�If.������G���6���|�f�s�ϯ�%��vV��>
����u\tS��h��u�!r��D���Z@���Ե !���˛����w�󅕜ٽ�+	�dP�����~��EA(�$h�#N��6;��X��/�'_ժ���ַ�8V��C�Q��^�z�t�w��xS�J��h����k�0��쥜���.�"WN4��j���E|}�'��}椎��c�f�!��g���ysU��w�jd?�Al��3�u=���ӳ��gkd�I�7��kj��Bxi;�栰����mW�;��+�c�4��u�hYC�4�r�ݺ�Pq/\� wۃSL�z[��+��w`� ��>���n�&O/'F'Yݶ #�9��q��B��ő�
zn�]��yL��9�yy�<���x��G��ֺ<�2��^���r.�{Xl��n��s�.��^�FZພ��g��N<�.1�*�eCu�a��{t��La��V\�����cXr��峮�
���i��-�v,e�'Ƀ�:�S[��/c�ֶgm̘�u��q]m�r�f���*�}�s�P�V.
J3>��h���!?e���z�I���Y���VB�&�7S��*O�����ez��Ng0_|�>><*0���=����gDļo��i�$K��Y�������&8�RG��?~��~�����i�<G�Q�9<���~��g�0��8Z�7�]�m� $�$A,=�V$|�B���B���p���r�ϱ���OHO�>�}��#܅}q�z�-�lO)7tȥT�jm&a�J�>�s�i3�t�:�ӇK�ƙ
�ds�
��0��	/Fo{^����� ��}p�]�II0���y���Ĥҩ�D��#����l2��'iGO��4�A��-�u(�z~7�������9qO�yXQ�f����R3�\��`�A�}���t��R�ᅘi�ֈ=ϯ�p�B�y�>1	k�ϗ�s�/�w�}�Fs���i�:|M-�R~�!�G����|�E��0Ԃ����
��WlBT.
�g>��p�,"D�8�Ռ����멨�&��-�|>�����n56ؕ����W��L��I��K�[��n���i�ۅ$z�U�G~��1�n�~0�L��	�Ȁ��Gd�q�mڋ�{8��a.�;rʓ��5�s�sè�eRn���/"�bVQϚ�`����]���*o���O}{IY$1Z�9�����,�
�UM2>f+I�|�ϳ�__d��|�J"�/)ʹ�2�ۋ��~���ޑ��D�T�Ŵ�24�QUSp��ʧ��q&���5�`�_���C��#���O����H�͖�f��&�=�^@xckJ�7M����r'F���6��J�w�vV]N�p����`t�F!�Ծ�/�����;���I]rեG5�)��XB�\��?}ɴ�	Y�5%�0����n[����{�I��K�v���p�V���Rq�l�MHs�"��ad"�9LC#ڟ�E|����@Y�;� �$����W����8�N[�g9��zl0�v� �vd��[��M�E��%T�ߞ��م��7"U��N�(�;V@��q4m����m�c���_�(���~����>�r�~�����!}Ə�sw�be�T�u�
����{�[����&�g�gťÄ4)8��j�Ż)oҨo���g>�-ƚ [�Ήa|Ջ�:��_I4����ꪦi�|����V4-B�lK=�� ZK�b\�M�d`�\���'��͵��R���`+Zp�EDC��PE~�բŴ/�w^8D�6���de#���:�p�&���j�e���1jK?{wOזS��h(�!i�P�!J����u%���c�}��G�G�؎�6��瞺��n�?G�3�?O�#�!���^"X���s�s�=�����ș˕@*[���U�����d-�bT$����i_җ�^��p����k��|$RG���#u��j�\�ۅ�\>O��e�U)�5Lѐ���2�^"J�ܠ�֙����ե���U���yfƐ���1Q��{sx�����H�B�ߦ$�}8����B���,��nb��q�����:��Y?Wѧ��qSUmh�bxo�C��%H."Α
*�@Y'E̟k�ݿ��4^!z��ֲa�j�Lw�p��)0
��\]�����=�ŗ7rAp�D����&��)��n�J�]��iS/tNݭ��O5f͉�&��m�a�;��$	)�7\ݫ^�ӻ������5�*�ޱ���W*X���K��-�����+Y4Lh��Wrb�0�]t`��I���f���2!QFÒ;�H���L(�G�s�y{)�v�/$V�{�>#�ٙ�!g�cb�3�s���)#�!{}7.9�����J�$�C����/����ϹάQB�{��<�q���mFu���K_.�m���*	sT��ZF�-�e��b�k[�����r�VB�p�W����˼�w�{��V����> f���М��HdS����3��_HZyNJLR���*���5|}HQ���~8�׬L#�����F>�u����l��f��3k�5+<�]3��賧�vʸE����ʹ�6�j���Tv�樓�)�	��;p5�VX�������j���N���.��/�X'nZ}���ҟ�߫�s������ Q��>r+���/�V�B���@�ƽ�X1/���%̽�H�BD���{"ȇ��t@�[�����W��y�͆/"/�H�,M
N�wU�0��L��T)$G�ۿ���
����1+���V�N9� �{��v"���޿�?{����߅��E&�!��M^O�w�*�|��XIY��xs�>�ńp�v�Y=[I�b��.�>y�ɉGK"���\�'�Z{�0���:��p޶t�!���UﯜybZ%�s%R"��[*Ήg��}b}	)�`n$�?R�A~t	�i��߾o���ѝDf�;K5�g\Ɖ_�ܸ�/�5��֫���"Ƚkq²ħ�}�� Tok󲕐?/�z�`2d�$�P��qvw�:��s94�|o��a�I�B�~&qK�o��lYm[�G���:��O#%d��vVvV^E�G��x���
B��tH���ruCֹ�{��?I#�D�H���ag�}M�`�	[Z��B�{�з�¢�����O�t����{���Ĭ���,�gO�X>l�_>�+-M�0�-pW�ë�ߝ�pJ@��O�O��&�O��1~���e���6be�lD�O����\n;X[��U����]�
�0���jY��:iH�T!MD���/��]M�$����z��M�����Ym�&U�	�q�o���۠:D�d}�V`��F�>�,�
ύ�8�ɵ���%ç�]�����p}Ϻ�q��k�)��G�g��g	X~(��d	��A#���?~HX����+!���;���]���/�O�����2+�E���B�ʗiQA��.*�=ʩ��қ���=?hU��YN,-��Ȼ���e����"��[ӿ`�Ea��+G���
���kb�!�$A�;R�!d9�8���"s���K�ƍڮ	����������U� ��"Hߧ�����fux�C<K��󵢥��+(Z*-%���6���_�x����)�$YW�3���i�T�&�4�-:y�T��!����x�إ_{��ө}�}ϳy���l��T)"E�.";~Ϧ�8׈4�)"��ZW����8&��0,� "RDY�����V.��z���\�u\,!}.�Q��f8YW�?J�EAhDெ�D8�g-
7<�Y�$�{�M�N�"�=J�12��}��*�����ݻ��D^�*"��!Q����X�=���=/�ҳ��zB���Ŋ�i����_��j�@X� ��5w�E+��b��-��������P����͐�ڽy����R����s�ÚIp��u>�2q��N�J��Aw�o��;i��&��"��N����U�g=:۳t��y7���!)���nut8ۥےMܴ�rV�·�e{U�wcѻ=��t�ܛG��͖�%���w8�msrl�\a�q�J������X�9Gb��G�dö���������S�=6ͳ�m�ϑ���h:l�
�9�����ݮ*�\ڏp�=t�n
\�+����ڻ���l%���8^ue�ی����gֈ�(�=�n�37Bv39�d0'"LD�������'O��	�	YHJD��/�O Tp]߫�V�^�
HS�n|d'��K��H����괪y�^��2�zs���B�q�B�;Hp�F?N7_���
�f����恥��?`�N��QI$5�4�%e�w救�>����-��U�|�;K9��J�Ɋ�Z,M�y�v%�x^��~|4���~�|��\!񢟉c�aG�y�V��:^V��߳^]r��Ƭ�*��ַB@�-��,H�w��E�C�/�7�LQdb��Z�p�L"��k��sUB�K�����۽3�
U8����>����������[b>r*4��/7���n��mp^:%��dM8�氀w����z!�B�%�K�h���&����X���,~6]f�P���w��Y�g�*(�>��V,����KO�O)x�()�LJI�
~��xd|r�2*w�j�&&aŅ�_o9�s�{�b�4����f���`�t�F��6R�U1��琗E҄ۀ�e>"$�q�y����\!1u������/�L��?qv>�3�� �@���
�
�^;_��-�l%mi�L�XIR*"�>���8.�,K���%4��W�{瑩���h*$W�(v���7a^s'b�t�j�u����ɩ���j�rAv9僸����~���*�e��QFKW��U�#EdP��1�P�O}�������Ve��61*;S�K>�۴�|sI�}���{�uċ�ɘ���+��Qd��k뙍#:��l����I*u�k�	��I&W�$��#�r$e��sVY7S�j���S3�}���}���8�bp�B�\��m:*:���ϳn�2���Ӥ`�+���,�h�7�;]�v�i����CcK6>���_s�U!���d޻_�|�裣����}����3ɀ]���i]�����N(���(^��XF����OR�:~��� �kT0�D?:��41A�RB�Uʞ5F#�}6�-ƻ|�b�XB�u�b����JF��p���3Ƴ[.�m1�1U�g?)R���5��Km|, �%/��3U�Ϣ��e/�?2^ O���F҉�[Q3U������a�����g��y��p����u� ��$eҌ½�Z���|/-kI�%i	���˵j��>	2��K鯴�ͮ���iϾ����V��Ӎ3�e��R'N==�XE���&޲�BD�7}�LA�G����B�`��)�Ջ�u��9.E����+���w�[v���G�wڭ/�7�Ƌ�t5n$E��B�}߾�Z*o�M�%�D)!}~�����ğ	fj��X�~�����c_�O��;ԙL�Di8� �՘�9qA�,[+��;d����;��]�n-����m�'�[����~q�sU�$��|�u��U�h�\�]�%"u��}��������g*|a���s d>��i��<�|�������i����!i��E-�h�w�c�}$������,K@��TB�g�Y}f}M��W� �{/a����{�TY
��ξ�;�v��q\P���q�*-M�l��v����s���9ʌ$K	n7�Z�:+�����߁뵡�l�D?�����j"�Ӛ���_�+�BV;ybp�Ӿ���ƤRQ
��H�
�����Ţ�ﲨ�aP��ޙ���P������_��ϲ7�o�ɳ�/b�-e5�;F��[Bu���Q.�_;|�:���(.���X�������"b���b�������ni9X��o��3����b=�6B�
��p���t�"���"��L�wu6^X��)'a��<��@��1*ė�;gcG��C����AJ�׵�� �S�_�Ym�v��Zq�o\}fg���w¢8�9]}��u�oo@P�Jz�,h�i���g[�1�8u����F�i�|̹}�n���|�����~�/J>b�@IX�����t��Jm����p.��u!%��&�~�Q��mm�n�:��:�n
wve\���{���q�8�B��ou�Y�(��W}��D`��z�N�w]E����m������fb��VF�.6��f��(������E���EY�wg,Z��y��Y0�؈�F�u��7�ۯ�Ĝ<!�b���c7��ʌ6�]v��I��w�q��:��t��-N��wF�t���y��p���d���ע�;��XL.���]��AlQ�x�������@���v3,�=���(j4\s��D�-��p;���mt�_����\ɉ��Җq�ke��%�B�9�	),^8����(��	fU� lY��C�F�uu��X��ġ;�렕g*$�r�nnCsAϺ�iM��q���ͧf�Üz�EK���D��<�h�V��.����F��Eo3)�S�S��^]yn�8�������d>�+�_k�V�����N��TE
�~�m_�p�̞N�*F�<�(�Ѹ���2���˨�����Ĩ1�tk��"�O}9�5�f|W�-�с:jw�V�c���3X�`"�P��qZX�sj�- ��R�n�"~�|�pU��uc�wԴU�:n{�%p�����ԓ�~mx�g;����}.t2ar�xT/�}o|�%Ӥ�MJ�R斥��N:+���(R?k�g����`�D��~t�a�-���=���k�_�J#���#X�Q�9;����v���);��,X"f���_٪��~~ � _k������x�X�џ��dF6�ve71�v�m���%�ѷ%�=�^�ؗG������}�VA]ۢ�|ȑ��
x��6V����/�;�Wu�s���:*^�*��,-�>wD�e)(���!���V~VD�~�	�Z���`�Ew��c�2Z|�
���HX�(�!�۽ ��j��[�+=���<�c��s�e��sX�����'W���p^5�2�\}q<�ϱ$v+7�Q
����/�j0���o-*��w���t�"7��lk���_�R�̯h�}t^��r�u��s$�	/_�QV|Y�],���^r(�B����r8��/7�<Q�>�����z��Ν�ջ#�>i��s���,剛�w����l�q�%J�V���i��ŷ�գ{��U��,���rwm�(,R�)��)V�a�h�h-Wcz��9ڵ]16�4@V�\ ϊ��h�[)�f�U<��ǻ&� �S��,{ޙif̓�;u͖MdVL�^�=��Դ��=��aY+�m�Ӟ�H)�̼�~��A�����8�;�c�n�,F��+���9n�]�{g�F��t ��̳�T�aA����Jq�	|s/�r�y~�&=Ycw���Ɏ�Y�(y�͑.�Y+�U�r��}���b�a�^j��6
Aȗ�%r)�
�����n+���k��Ԩέ�ˉY/%�v��c�Kc�~sy�嗈*J.O�?B��R;{�4g[]��6����#I�A&�b9$��Iq�\��z}b����]V��o%X�c^�h�=�l�x��뻡l�h9=u�&��i�`�wpg��h'A�E��f1�i2�����JWZ�[sX�C6��i�Ǡ��ЉQ��ݣ���|'m��P}=�rӞɕ㚣�����n|�� �#eD���&Pcf���xkl�L�������\;'����;te�Е��#�WN���SR0-c"�℣7�A��v����Գ�U�}���fP��[�����nVjWI⸚�I����Dk���,��G��1����jՉ5}�a�	=��Z��)q�u�"�ñp������s�Ȣ���c��L靖��۳�ծ�f4]kc����'n��X�w7���������O8��vV�&;u�cۮAܯ��u�6�z�J�=�C�s�U����v��5m�3�nn���gˆ�ώU��jq9j�s������Bv2Cm��<]\�<�-�R0�ۭ���J���=m����OlZ�i�E�y�����&qd+�b���F�Lg����k��nz�ٺE��Q�(����n��C�uy��s�!~��%�Y%�4U_��&�E���z�}~�6�<���3"�;�dd"#q�[�Ig�He�JC�h���3�X��Q��\?y�
��a��j�3lxcCq7��[϶9r�{j�Jp��I�j4	AH"�E Tt�*@�Ko��<�U�OS��vi��\*�g�q��;���ĸ�;.9��*ݶ�Վ��J-�,�h��"�nn.C�Ww4��q}��ѹoK`�:/��}�Ɋ�+�zSn��蹅��}y��b7��k�*%���v���l�#R;��:�>��{ ʯ��TCV�/j�~ܤ�y�k"�$�\���A��Q]�{��me�AR~E�.�j�k�U������q�GqG���=e�V睎;]2k��:N���1� �s�.m<�u�u�1!��mi�}Cn�*3'�Vn_%ݶ՞Ձfy�md߼O��d��+�{�wF֍F�6[��|@Ul2�0����aPf���oz��V^_z��C�$򍗯1��l4��2�ޮ�·QA#.�8;�#���(oom�ư��t�:���M�&,69�C��!i\��V[�~��N��:SA�!-����f;�sj�����Z&�<R�kj��dE���ā2ECG���{�aU�GK�K3-��пe�^e�$z�/�\�h�]�خ�^.�5C�Q�x��cm���zr#&9$n���Pu�ښ�L�V�{vX�P�iv@�le.u�*����^��O7"u|*V׎g�΃/�$z�fׁm�����R��T��Vs�
4,E��t؊��R�＝N�RD���HM�����i�lu��|�S��p�n�vz��h��ݜ���۩7JfC;m���*X�8����n����R�����&��Pm��w�+Q���p�O��0��׶K�/<�nb<&:Z�W�2�B�£k�
d#o�M�jn�r��{�6yu���y�s%s��+	��ԖU�+6�E���y���]���l� &Jk���\ݑ<�˞�׮�Va����ݩ{�!�5�<+�-�Ǭj���oP&0wl�3�0'U�E!����*:#3>�h	W��͜Q1�<D8�u��^݆3d�㮛!>�MکP'N��F��&��\��&���r&�KЈ�&̌)���T�N�l�IE�x�}���I��T�B�!�~�ök��!���v#A
����#���\~<8�RIpHBiH�xF�&��.�}�1��'sy�����>�l^X� N2�-Isi1g7�5Y�	� C}$Ѿg�����;����Q���nN�c�q��||}��q�Dv���`hƻq��q�N�u��h�z��^"
�D��������yE@�{�繭�j�`.N��켴Z�&ԥ\=|�>=X��2+K۹���i9�kz�Q�H�R\R5y�:{�U�Z��Xx|^#�����t�~�^+���fmhO�:/P��r���شĂYԳf�M��\�ýx�Xb�AE
q�wG7d��7a�4�5'\�˭�fu=���ݗ�q�27@���K������F������6ZD!�M��c��G���ȥ`�h�S�2`�=�t$�+�3�!��US��2�K�<>w�Ruv=3��$n�{��ck��u^i흗rZ�nGl��r�.��^CIç.,�F�;J�z�%Ox6����h�e�rہ��Щ!��������Z�����S��3���Np��p��Y�i�=�u�r�S.y�6]aF�L݊��M/&�U�2阊���h_����7;��YV����̤����:{dk�1���3�bLHQ�����KMG��j�X�T�vo��y=8�\<rS��CS�.`���.{ކ?w��T4�,�Y���^6-|��d$Sq� �8�8�E���h�թ�*2H�� pAI��F�������͙YQY޺�]�ί�X�(%��+�!ފc���I�LAD$����kճ������ m��# ��c#�=���.GBf;�J��b\��.�`�tL��;miw�MGq�9�M��S4ѕ}U�E����Ʃ��X�7F��+s���gt�;��g�7~F�@�-:*�1��Y7׸m^K"C��B�]cs.uc]�V������Xs�)}���|��`��qwT_$���>�lvIF����ʥrP���a�w�g(]��u�U\@��-[ufՑ�5����O#�.1l �s�ҭG�b��WE\�T�0W��l9!�(	eBC�S@���ɲy5۬�<�<�V�^�v2����b��g�:��9ϤB��Gc�q�s)�ֹ;n��7nqo0G/�v����3�M���g�h�izy-�n��^�'��+��v�C����a���r>�U��h7�Fs��W��F3U����L=t�K�s�]D�.۶�b���5���Iۍ��'�J���ٞ75����k �ѩ����g���i@��l	�v/Fq�[r�7�l��p&�nA�)g��[6���3Ƶ�%��I�����c�B�+mb��ز��}!��d�������%�I,��&n�D�\���̧�+�ui���h���jhk�경�����ᯮʥ����=�֊�����������7AC"m�A��o6��	���U����gu&��8~Tc+5Dos��i��g\�w4.�J�՜��*G�Ì�ar8�����xB�e�x�#-��H��J�L��𔨺�m��yf `>�ܰ����`=����,3�T�J,��9�Mpl*�2��R�ˤ�,�O�z�q�זl>�ȍx=jX+��ѻJ*�1��_vP��y?qȐ>�]�����	�S����A�:g�c=�u��N�[bK-"�|�L.
��S��}�����4j>p,5���j�l+0V����n��׌ె2�z�1�c�[`��l�$4
QH��:���۾�M�qW��*���wĆ����1�,Z���d�|�ҁ7b�V�H��VTWG.��-���8�����\����r�U�E�b��/!)��Y�P����[���v����\�h�׿,��>6�$B�p�j��3���mہ����\!�'������U�}v�6hA�W�Y�z8�(��u*ɷ�
S�这�B-�W���c�|��7�	�Xܽa�Hذ�_�F/�ݖ؅����6̣��@[�)`�����7}�,��9TM��2�����Ci=-WZ�`�Dd�������)��q�ĽZ���<VTe>��蚳�oÛy��i���rќ�~��c���d�n�� 3�59��8��z����6�����`�]<��ճ�f��H�9:su��F��/���It�L�zý�U��c�d9��δ;y���B�n�ѯ�]�a��~I� $���&1�ժv!���K�t��y7���Ò�N�{LA&��R�47��#��^�6�`h��7��Ou{/�M��n���.IVv�U�~w^xe�Rԡ��0��X�Qx�3��*q�������"��u�Ya67(�Ӫ�a-�Kp+˃
W.�j�	��N�#co77R���J����Dz�'_CIRմ{ΧaZi|\�7=>=@���e��n���HO>^�u�쭭�>;&9us�ȯR���4��y���|��f#�l�w�)�ۃ� 2��HQ������
mQ�z��G<��9<N�Z;�Xb1���t��ry�a�w��}�h�/�OU�U�Z_����L��J;T2���n} h�!C�z�����p�F�O^�v'�w��V땷]�;�*�%�3L6�c����d��t�Ç����~3A/����K�=��Bk����'���y�}�G{G��p�7��w�7�Y���&`L��1Ó���{O�m{V��6׷:)��}<߽�Ӽ|��\hby�o=_R{�������BpS��U�p��V�PzIL2Hd0�m�ٳZ����15u��f�A����v:�h���[a�t��l�k���2�|�\�wg��3f���iSd�[L��5;۝�5���Ѯ�S�""���si�V����LyVГsh'*#�C���m���	Ƕh�ܸɊ�oY��7;NC����!��gc�;�Z����ӯ_=�s�[��2뱋��ϡ������3�xN�JmAu�5s`����f)!~���Ɵa󔡧fn||W${j�v��8�z�6�������i�@���U��Ԍy욎Aވ���k����k����8u�8�Y�%�]b��%��e�2�q=��3נ�X�>e7�p�g���-/]Y�AZf]sS+�ݧ)��t���}�ndf�M嚁��A�N4�BcnA@Χ���m���-s�z���v�r]�l�E�^��Z� �Ӌ�8)B/�������T:��OkW��^�<��n��.� �Z�L��]b)cc{6�w�a�<c���l}�dt�w�=�n� ��H��[�4��2N}��|�HPf[,4�
��Y�����`�X}|2�}R�
I�;pt�Y@��;��f�X��S��]�����Ĥ.2��2;�(8b���F�RMwk$}i�*Z����4TFn��B0�L,�\A�:nٱ��6�^8�3�4��9����-e�[�:M��G9^.ɸ���|�s��b�C{��nI7��������uY@as(om�Uʯ4�v���Vg�������(��:#;X�*S�W9B�e�:��׎�v
'с����%�:Y��^ef]���Ǆ4{m�\��b��9:�/��J���#ȱ��+���`�$������&|�d�1�a�]Lm�9tJQ���@LK;�y�>ͼ���a��ݐLy�R��d�F�ly�
�}�yt�-a��p�)�D�q`Ѷ���]C�����*�u�3U�?q�nd�(b˼�=��t��;�Oqv�|���`CPk��mm�z8ͼ}�|��^뻚꾷:�BGq��}/���v6��!��!�NWG�9٨v��ł
cGe''!�X��VmP�GH3�gqj�'R�,�ι���xsEYy(w9��^`j�n3Y���V���wut̺Ą���Qh홙&����:��{wX�G]�kC��c׹�f�u�/n�1h�׌���	=]RU�7�Y ����#;�\��.V".:��zI��Fh�G��뎳���k�M[�-1�4��HܔA{�[�y�z�G��M�����*_#L��:W/6T����@���b�CwG9�ܓ�K��V7Z�l�ᎎ�ѯ����۫�F>*������.�橛� �Dp$Kzl>L�c�q=��R����'����w��6�x�	SO�U{pAI*I��m�����e�҃lJ��0w6��v�uU8-��ͤ�n�ds���U2�q�l'\<m6��͎#cJ��m�ӷ��x�m�����N�5�5�U<\&{q/��.�n�ͣo;���=�I�l=Dۇ���c�[q����9�ϸ8rnɫ�M�9��۵x\Ζ*rsǬ���;�\��m��\����剣n5�p�;v����|C`.xO�����Bd��V�� ���n�����6�{��v���P��e�^-n
�.� �񛀷R�&�u9ήm�m��=4��m����]���j�8֌cۧ�N�Va���K�h�� P���l�7���>6�<�C�&��ܡ��6�s��un]�ök��Gs�)t3�����UoISۆ��v�Ç��݉�H얳��O:;p����8�Zź��[���'��\�b9�vp�Ϋc����WX�hݘ��{�{3�t�D�	�n�v�]�-�nG��}�/�&�E��9���pC�ѧ��J���1�V�{s
�y���7n��&�j6��;���X��`|-Z�C������ n^|�ݱ��m��\q�I��i�������x��wnޞB�8��vn���DI�n��ۥql�'j�����5��gfs�ݥ��-Y̶�7Y��Du9�q�-��V7Y�q��s\Fۺ\枎��2�.�1�nƳ���s�Õr�*N\n{�'���*�|�k�`��'c�nAm�XM��#[�x�.�q'�X���k��%6q�V�.�H��.��q���n7I�;�O/^����Lp��7[���=�6��x)�%���ps�ݴk�-�$��&��W�;u�k#�W�8��	���ӎ�=�n\G9�lEڒ���:���Xe��O�yK۞ɫm۵��$+�te��&���7S�V���u�w{<u���OY�������{�[�׎��ۨN�;A��7i�3Is���;�Ɏ� ��N�z��v�.���i]���ˆwQ�l ���8���X���i:=v.��Ź�X�{�1T{x��q�S�!��h�=�����y{d��:�=l��ۗ�Xx�K��[D�/]���z��^��	ngɷ��[�8�]���i䍺� vI�y�Ƅg�qC�-�h�cs�f9���i���Y��e�/�2H�'!]�����n�w<�v8��kt��47,n�7P�(��s=v���i��]��N꣙���!�W���q�v�n�\����T���:.�ف�(�g[�'�ߋpǉ�W	޷c��\���ï5�&-������s�����*��"�d�����X[��+ҭ(���[%I�L���R��>W�)i.o:���¬�.7�+(_���fKلmgL��lۭG� .y�� �j'"��G�?u:W�T�˽O��(#�n���V�j�}����Ƚ-�Uf^��2��qѦЄ�2�I��u�朡Gya�X�����~9��L�쏷���ˇ}�V�gE��5\�Z�u_�v" ��5=�����Ӏ�$(�T�w�/��Z��}�R�P�:}0{}u��ꇟ^�޵S�yebl�C.���ǲ�T�犙T��(!7���u���\Imֺ��t���z;p����.�E7�Dt��C��n:�s���¡j~ཡ��}y�m��-��~�D�N���a8�;hA�Հl&ώ�N�wד��C�'��{��'�"eYڶς��L�)�t+i�vB���
;e�v��(�@�զ]�y���v�H�'A`�N�?�vq�K׹�{^q�����W�JY�E��{��F��ˑ�Nٵ.u7��K\�S�c�3fn�]�&�F���7|�t����=K<��f`ٴ�8[�v�n������d.5,��O�3ܨ��9Њ�ya��	%@�) �맦��l���6A��|�R˻Dm�����a��3qɯ�y9�gՀ��V�G��ߢ=����"	�Wv�>�<��5�<�N�<�F��`M�9�Y�H59�<n����}�}x���9hӞ@'T�Zt�)��.kv̺6n�c�z��0t��O�Nj8��F�4�fb��������o��F�{�e���]3�î��h̆�n�)����
���jҰ�
�mט��@f�K¯� �p&�(�#q�s�m?y���R|;X���l�9/[8��x�� �K�<e��B��l�s"��{��6��`��Į�Cƣ�
e�$�+U׬������C��dã��hVm�~e[ACm49��W[���C����+{Lub1s�v�S�c��+����W]
wy���Ōˀkv�o��x���MW*��R�+�I�}%��T�ԭ9)��I��U��Ĭ��@��~M#���L���"f(v�[��ww{*usE��L\�>QZ�K�9��Q�j�9��i?bU�������|���IwVB���|����M̤�]3*�.=�y�+s�I��4Ԕ�z'��ei�ry^2�����UQ޳��ƚ����R��O���Q�D#�gn��J3gn�E����p9����n�,�"P����<�U�����ŧ��ڑ&3h/���#x���d�d8�"������͈�Ҝ�n˶���~lA���dꦚқ�|�1��Wu.]�y�Tmx�2�ڰ��y�9}�����3��m>P�v��uG�r��XvZ��ꞅ��g��߉F9�2�r8�`��ԫ�b�uJP���ګ��@e��w��;���cٴ�A/Ø���������J)NǗ���@ѻn��|�9X�;u���b��Gh �FO��lW���+��2�����ͼ^�7)�C^�4�u+6.�#�r�{���+�U�gg�
�'w��-l8:ִ:��[E^�8�Q��a���T\�f<>^|�țm�rA�cDU&��E;����#<�EY��`9�/�;�b�ͺ�Vb�Dޞ��a*�$�v�>{Ksau�,RTn2���C��cx�'g�c�ny�r�۲e�p=���ō���wnvұ���/���q�r3�{~��d֏��ʇg6<*R�	��׳���*�N�A�t����@��� ����Z)94bJg^j��/)���eD�w��7��e,FR���̤X�|I~Iɫ;A*�7�����ن���6i�om�EWU�o+$W{9�,.��4[�p����ZvGf��Vg�����>��+D��=�[��N(���ƍ��B�ڜJЖ��Ȯ�c�jw5��=5s[���bxK`��6�#~�6��$�F�V2�|���;څ������&II �[t�U�nw\���V1�]���?{_�IB��&��=^�p+2���<̞��YP�X�T�A��Y%GΧV
�<�0�#�w9��Ŋ�j�ZyV�7��o�5�j�T�'	�p�9Nz{nIi�����'��{�Hڌ(��RS�牄��������qH����NY����noX�%�z�����ۇ�ۂ��۰R�;G���f7=Z��]h�V�J�m��g��옐����fw=����t�!��du�.�l�n�Q���z��[u��*�y���.�� ՗&n}==��4r��l@���>�'s��rk;���̰�����A4��͹�z�U5�S�Ʊ�t��]��lX4h��=�t�:��k��]*�d�8h8�m������6h7����R8�����1���Ӿ��^+�t6yq"��]��߱���T	�=\�R�-�	�j����]no�5�E�/7�\���ޥ��Gi{"��(�^|�F{�Bj�d��� ��<�s ��lH�EFڐo�?��)Eκ��	䲼1��uxı���w.��5���A�2�L�/+&���hQU�Hn"�"�RA���C�qf�vEylR[�em���{/q�mqՓ��1�x9K�,���[+k3_L�Z\d[#��}���)y!��1"׎�1��Y��E�i���5���2c
��˷�vϟ8;=�a�Vk��gS_z�9/�A]��z��.j�� ���:jv�\�T9Z���wO�1��`e������ʾ�Sg��[y��ps����_r��}q�};LrWc&��X�����H&
��u�J	q����1�����{3�B�_S-@qvN��mwkk���5�{�{꽱zM��K�a�o-�4�j#x�K��v������2a9��0��[�;��4�s��۪yw�$t�.V��ː������еkO�~¬��t@´��C�g�F2�Q���9	t\���=�0��
!�:<��i�q&`u ѕE���pۼB���yԍ�>�@Jdjht>�lH"R5)��^�F��K����E�`Ә����(��(�e��ۧ��x�kݥh�&�<-�̬�W�)�EIã;2�ԫ�x�X��pR��w�ݼ����6�M��L�t��;X�0�<|���1J�6������}�U�H�"�)� �Y�a����[��p�v���5vb������A���@����&Hv%�jxˢ�ۛ��ۓ�{(��=n�66�T�#o�K��*B��Q��Ĕ-�A�Ba�n�i�t)�e���EZ/\��%��1u�2�g$5؆���|w�qKc���#_/�j�{�����B��Q�a���sP�;������m=��;���CCլ}8���{+�4�(w��.*Y��x`�֎�M��W@�l�]�u��^F�o^'�}�C6�%��c�t��ב�n@���k�}4b�����kw�zE�� X��AF�RG���̷w�>��b!g�M�f����4���Z�4���z���f��^ڼ�9mA��^J@T��b��`��ܑ�ԉ1��m�<�G�x��jUQ�KUF׽~��V06*�K}g<&��WCZ�yD�ՁAÑ�C���R%�$q�"N�ۉI:��tX��sՃ�5h��W75��{[�i5T�):�Il�ŌCNgB��w/��O}�Io��(A�̙Y��*TY�iޛiV�����L��}3�)a�j�q�b:�}:�~>�+�R#GZ^����Z7x�d�p/�m�Y�@gIᕦ��r�]e︶������BFS������{��ʹ��2�Y���X���pI<B��q/��Ѯ�^�s�u���zn�GQ`�ҏ�I���.d���Ifu�PYӊJu���k��5�yJ~9<�㗚��O`�8o\Bso�5������z�����w�8ly�����^�C5){��Tw�G5������M�46ȷ�(kөB<${>;��{(Y���H�A�p�Ix0�~����
m>|V��y��-�$�>]sM��q�r�>�.�C�:em��<��՟�����β���O���|[r��oIO� ����*���ۛOh��.=U���/I$�9��\O���waj�L����.��hP)h�dޝ�{oqZv�6sFP2G�]ji����-��ѫh�{
%$�������+΃�/�� zI���dz�߻iv����~���:�	���30��'��sj)�'wB����}L��j(�N;�RMV铝�3s6u?5j�mm뺯^:u��f��!�4��`�T%q�;{^NM0KA��k�_D�f"ێ�+կ ���kQܵ��v�q���׻�o�$q�[/~�]�5ߵ�� �{ĦoѢ{o�w{+�U���������I��E������Tl�	���6�Tr�_Fdi�C1Y0�Ҫa+&-����n���K�Ƿ�-S�w������޴֤:;�+���,����n�rV��DLޅ�X3TN^A�O��o�8��[އsy�'z��~�[j�n�]�uq�ۛuў�n�2�b��n�7������A����nv
Cr���'g��C��B�.���u��둃g�]T�z�B�^���vU�z���(`;\���V�OL���K����7��{��j�Lv�!ڵ��A���r�b�ɝݞ�OR�n�i\:��M̼��s�z9Eƍ��C�Ӫ܁�c���^���n;n������6ݮ�-&����g�>����\k���m��'���tqxu�v�,�9� �$)���81�/\uN��3�oO�Y�c�T��̂e+Gc���f8�v;,t�Ɯ6qt�
��6&�5t�]�!@�.9���]T���,�=�Nl/<��������4���nE�y��a��y�ү���-CU)��r�`�$7]R�3�}���o}�s|t��?
�܅:<k�w���������i �UɊ	SF#$B"��p���X5���(.v]��c��0�ګ�m��86�~7�� o=���ʴ-�p�.�p>�4�\�4�e7 xz�Гݷ�FUh9B)�}���Vm��se/��mʍ���?XM��.����"[��}��`wj�fa�`e�<邢��A�)��ZX��rrm���%��I��Պ�\�#.���SC��?L�z�`�@ i�}-��o/dڐR�P澃r�\G����Thy�ׯ{��_.�G�K���K�1b2�p:�[��`��[�6��;�y%4tx+�&NH5%��(�ȸ}z�z
#���O��إ��\]�yJ02����DyB��6V�k�X�w�0��=5�ԫ�4�"1��B��ݴ��ܕq�*/��һeX`˽�Zɞ�4߸�&�O���q�a�$��x\�Q�n��hZA(�[~��,�/iJ��:CP�)����ݦg��{jJ>��n���V.�`���$NtFWK���p�����}�/���γ2�v�8Ԙ/�8q�荜�]�|bL�wl�Y�uq@Pr6�T�좹9N=��L�̪J�{C��}�i�n{"�sd�{'�lR�~кB����}1B����;Y���)}��(��L�\h4Xl�+�5秎u���N̝�h�e��;�g����.6�)���ѱ޿N²%@�2�,��>���5�~w�u�p��M�����D����L$86>�5l��N�l0i5�z]�׮��Y�/��5f	�M?(��3\���M���������{�Co5 �^WZ�M�.u�ܩx� k$!�hl�4"</d�tQ�A��QȘʯ�vEh��i/MCJ;:�&�P���rt۫�s�vwi/�ג�Dp�2��{��X��!�-U��WF*�;-+�Ae�^g�����a+ݷ�:�]CL�%g�*`L����-���������6��M[��oyT���$v��*DC՜�u',� :s{��p�s�Hx�.W{��+�ֶ�X�p�V���l�ᑝ�1g�=���;����x���&^�	HN��}������n�ӛ���tl�G�+���5bBw_\����ӌ�n�Y�U�k"��n�vj���Ѕ��zG�2�oQj��Nܼۮ��*�n�k����$,ppﰏ�1�'f�۸�:��	�.�M�u��*�֝�S��P�ʅ������l;�\����&9�4;��յא��� ��!9���`�x�m�b�b����(f�+�Ts~�����W�ZX7�uh:�^��� �Fɚ�,R�Y9��0r����l��mn��f�����.
�7[I�D�k�$��VlW����-꡽u��.yd�R�٧��뛬=ޜ�s2���rGf���U�.�@a�s��F���H����� �|��*��v�[W����+��C�S&�,�go��{�>�m^VT,�0o;�j2�������V�`�ໞ���v|+�[6`�9Q�H$�F!CBV�y� ��]�Júm�x�׳Z�W+Wz�-찜����XV4�mv�π-�q�X9sܧ:��.� H�&ճ�;�ϴ%)�J�i�K��<q��6�Z_�7�i��H�~�탺tV��ZR���xCm�Q�R
�p��VCz����<}/��9�{˄�{/o���W�p���q �n���:z��|�����F3��y��x2L2ٍ���I���A.X5aV��?i;���ۊ��苍=^�p]c:I���8-�ׂ˃�un�z�8�f	P��rH��:{]F�<�8W����t�ڕܮ�.��#v]pZ&X"��D�v'�uqcG�������yD#ͻ�l�^xo%�l릋S
�-�}z��N��������H��1�W�r��'�&�^�%�\nj�j�s�V aO��aVLB�v(���{S+�lNE�v8Lr�:W�vBRf�ɖ�iH�!)
,��)G>������!�g�T������s*��(茴�_��p7��Q��"���m]�?r�-�T���iH++�y���4Q�V��к�gr��o���+����'����V�����Q�	L����j����ng��g� �� r�=C��Q2������
q���4�{aGp�õ�%��$X���[r�K���[FOK/%�̑vq�#�4B�+��շ.����g�'����	��bԆT��	{rz�f�'[�:�Br����E~ɯ��H�)5��&ӎ�P9^�9����Rp��Lѫ��']�lg\��t�7�lvn��t=;]���;���t��^x�����Yփ�H#\���~P� H]��o�5��i�<�(���wW��Y��X�Zg�>0Rua_�˫�]�L�<����_&N�!��P�l�@����P�7�۴S96����{pe��._W�p|�#M�M����-�.�^{��$`�2Y��:�[-[��=z�b���+P"����?0ݠ� �|7޲LR2�B���39ۂ����j�.t���}ԏ���ݓf�n��m]Ý
�x�h�3��s¢��^�k=���l����{�0,��D�m�;Eca5z��i��xs�t�HuX�A��ީ9
���^C�oJ$��"cV:wURY��`ii���^`<�s
�t��SZ�+C*������?u�k��PԈ�	��p��j{�U�m��M�E[�w�NvS���H�����`γݛ��lM���3͹��礀�� ]k��{r8q��t�v�,����Jh��������{���x��x�������h�zܛ'��7ӥ849�WZ��uۓ!��C���"]���Q��-@�u��S��q�c]x��+���o2Ɓ�:���kd}n���<�ɪ���m��<].;v6x�;ɤ0y3����Z����k�gb�+8.�[;��{.J{Jv�n���r�E�G�{u���9M���v�'!tl���՟��Z^��
��J�Cu���m�<y%��c���/z�������s�dd=LWq�2��9�$�Y_z5�S���ؔ����F)�-7�w�q��Ao�b�9}�y�۪V5I�_��ݟ/=A�b�`Mj-Ěp�X&H��[r�;ݐ�D�m�=��~�/��E�&�k�3��'���F{Yu-�*�ܤ3�̲ 7�a�@��A��y��9j)�:���x���Oj�����9��QR�t]d}�a�9�5������z1q��mT��f�$��P��nE�y$��zj�'��]C�T���h�g��+�f��]���-4=|�+��s�oV�4et�b�U�H帚EH�06TbG�����m���g��2qv���v�W��u�\���R&�#.߭�Q�έ�dS��G���f=[V�:��е�׮J����r~#�����:���`�E$�l�q�̆���c��*��Y�ǨW�|[�u8�ma��s��.����B�����V�2���_��F9:\�*0]��Ү�^.�=��ڍ>w�T����G���by�6IO�~�tU�<�H��m��Z6�S׷�b��W��J2��E��*�Ǩ����D)��u�b���vp�ł_���L�6.�;,Uԓlʀ��P߀��AH�MF�
��G�����1��>���y�萕�|��\���Nr��g��C�x����.iqK�Ǹiɝ���g��atP@�L2�M��$2�323�aC�o.��w1Z��t�� H����Yν�i]q]øx���y55E]U��f�p�,@�*��v��ȸ�N,��fw�m#��:�5��`��aA�D�1Q�A��#mN�	WY͔�y�Ы���޿r}J�wQW�!�Y.�{ ���=j�o�A&J(�1�oMה/�8�@��ʐ��_��=����	�y�9��}��HuA�*>vt�Pj&��z
�z)ȂD���7!�K��=�#"��~	����<��^�6GS�����w��8s|#y!�Q�W�z�:e��,xR��d�����Ve�&��A=7Le���&���,���ޏ�����.�g���!��V�ڬU�t���2�z��WN��k����y�;�㒯f�O�H��]*4��u|�A��9m9�\��!A�E�LkV3�}[�!�ȸ��}`=�#!,��s2�w�Cx"`���Y[�=�6'έ��tk5��*�
+��ۮ��Y�-n��e�f�r�bnr����P�s�[9��X����=K������lA�OY�zq�@�_g��4/;#��b�[��GRu��!a��/D����WU=�ʙjF��0TI�g����zm�N�}�x�8��(��,��f0]�r�F��[��^5~{ި�O-�2۬���O:���DL	H�ͺ	1��^�#���\���37�y��ۗ@��U����L2 ��v��3n2酯o�veg5�QI�F��Wv�Z���v��U��4i�P��R��+��.��A���B�//��O^ʗLׅo�Fh;��Q8�:��ֆ��`�Xk&��|;-R��3���Z ��o�I¡�mR��q4\쮝X�]p�����g��r�n�C�j�4��8̑8��k=6g�g��0�6�`;"�ֳ)��
 �`C�e�=�c�H�ƍLg�i�\�,j�3D�����M���6�q�$i�\���nsOkm�$���ݺ��0�n�Le⽗���F��N'^����E���U�`�=�V_< �����-S$*<��ސ��|�e7�y=>B��
��|X' ��y��
����>��$��ߣn��'�I�-���+���W���:�B���r{Ӏ&#�Ïf��{�σ�4�k�"0{�$��k�ѥf{��˽te��ٜ��p.\�%�86}P��]L��ˮ�E(Bbf�v��##($�p��[^�#���"�sIV=���t77��C�f��ǡO��M�Y��MbA׺��ά�;A���[�I�_mU�s�6�""�����L�Za����O؇J��ZH^���1�V��to�>|��`���K������îQ�!��]�>�O��J	\C.�b���x2�&�-EJ������!� �ntAM�3{*�G�Y���N�|aI5$b03d읹^g<ŝ����6c����v�j��:�X���燵mºu�w8q���޶Z�E�{�γ��F��v�S���M��q��#nշcVȬQqu]�ư���J�r��;��L���[=Y���2nz��lT��S��[۱�l��s�6��s��=�ᎰRݵ ��`8�gv�9q��6���`�v��U��|��Y&���N�1tq�X��P��3���Põͭvƣaci3�	�ˡ�^bY�h�q�B�Q��$����~j(VĿB���[���#��xFeЄ@�8�v�-�y�a���e��eR��i�b#qe�Զ�����vvl��z�*��2�T�%%�<z�.��%���u�Ã�nc���,o��������u�9F׫�Ȳ�����'<7l xx�l�0�JƟw�E�I+�zo��s�rU�u�96u{��F��e
%�N��+��'�'p��A�i�}R�'/�}�^��k|��>TH�C�9�Y�~%dv��tQWǕ
��!�-�H�)����Kg6ׇ&����������	�{$�b����S|1�a��Ǧ�
�d�>h=�Z����u�EN�R�.�P$�j)#�D� ����w>t��p�z�q�S�1cq��Zy�(s�`\��9&{��>��LxH�,�5���T:TJ K��wX�R�S��E4�VJ����>�ٴS�2�I�ڑX�2���EwU������p�v�?M�R��٣Զ�5�uJ��Ŏ�;P�?>����`��5Yb�Fv������#�L�H
|�]�7R�T:�Q*������|b�1����0�۞E;~R�nh��'��ܹx�W��)�	h�'��Y֋=���m�Ҳ��ʤu�����~0	��ߏ�LL^Ѳ7�z�Pb��!ho��V�&�)��\_>�/G`����N]��À�|����]�ot�9%V�\j�,ex9�OQ��3��Q���O�� ."R�!E�^�֮��&���:���,�m��s�+�.�l�ߐ�%����a~�*�/IY��?
)e��6h�D11R@A��吳��۫ �sA��g�����:�v���-��
���+3}vh���Y*!�旉u�����)�J��vb�S��5��/�al�8SL��
.��V���-�=#[\7z��F��j�0$ܵ������!Vb�}Inw�pHq�ٹ�8�w�t7�ʺ���r������8��)�4���m���l��KVֺl��O��
Ux�̗�W<�����On��\JG&���koE��M\0�Y���M���^��.#S�B��.�1-Tvj�i7ה����ueq��'�̋m�������ڌ{a~��[Ц�[RHԑmuCIx:�u�̡�(\��^�����1؍5���=�h[�昻��qx��{�n�wcF�i�h��QCM7�v�g�݂��\�:��4���]h�^va;��?x���]+���2l��:��Z1�%q��}s �`b�ƻC�`�:���D�����5�=�8���,	����߿�sw�{��<�l>��śP�z_T9������$Zq�����#�\����E��]g��)ptJ��,�P�\H�!M�!�mn��G����8��l��nؕ�z(��Z��pe��ҥT�!��`�����S���(a�
�t��(�-�4ڸ΅���>�މ{{��#=ՇqH,R46t�ۜ����|� �E�5D�n!u��t(&ڤB�N?s�3>��\��ϊ�:���o�.<��e�bVmDǲ߯mR�q��E�=���oXF��SH��]��;v�t����2��_X�6{a��X�������Fۙ��;S%���N��a�:�]�oD;��9�2E��O'Y���u�]�	p�$!��T|�6�N�Y�7-7�	��
�)�n�[�ݩOT�}��c�ʒ��U���#�z�3�NN����65�6h�ʅ׬�q�n��Y!8�cut2mv+aγ���������c7L;{s�6*�W��%��{b��>�V���MSM1��;�n�)�u! *S �[%6=�QO���Ƽw���`���K�`��'�N�<�
K~�>���A���⧚�	�����*,A��M�
 ���3*��B�]��!�0�K.<�}�[�9n��;ZνQC-�Q��u��$��1=]�j�����$�τ�h2i��M�Ի���Yr��X��v�>v➧/��ÁI���8}%�s��R���\:�����<%��];��XAf\�&\�<�?V�g�����aM����X�-y�����˧ز�z��bO�N^��S�z>�E��{�z�����{Hb�#���[����r��k)��˹�}2P��D@vu�)�/����1堕����/n�Yf��&돢Or����F�oc�2:��^n^ GM��)x'a��+9�ݪ)�75�܆�Y}ỳxe�9ZjGT���]r\z/T�p�� ���[�����񣑲�\�z�f}2GY����A]��C�~W�=��׏XF�=�h��z溔jrt�l���kC&�ʍ�i��89v����X�q�����rA(�2��'t��z��F���b-Bm��3*?�0b�e��Z������ݧE�9��[�ik��R���U����Ή��1E���p�g[ܧ��@V�ق�Ity�zNdؗ�'Ey^ׁ��pz.�81�v��޲��*
��uF	�g��G�ٔ���b�vP,r���\{���ݓ�����ͽ�owM����j�6�i��^oh r��V_Þ��e%����Ɍ�Omӄ��Q�º�qi�q�T�=4T��=����Ƥ�5�[K�������뺙�ك�s�D��d�0d��Dj�g<�!/��{G�M��g7�ܻ-�͝���_Tߛ2rͺXDF�)leϙ;�Bw$(��M(�������82�_vT'l7��>�*�j�Ur��*'���P�%�.�����`��U�lT+���ޕG�D�:6ԫ|��ئ�9\��{'V�S5<���\t;�	�x���vabӮwc���:����[F7)�hu�5���|�ak^�}\��c������.��+;����R��S�uT���P�yg�ඩښ�d�;'��m6�[�&��_B0v��6q�Sqg�K3�1u��z�e3�f#�����N���&u�<�X�&,&�<\�Zy����B]=�L=�l{!��3��ݎ��Յ�jq��Yk6ɟL�wnîɒIm�����v�s����'<s��Ѭ�#�ݻ4��6���:��=Y�N�p�e[q�k5I��^�u�����Z�l���&�wH��s��+�6:�W�X�/�T�:^uԣ�S� �R�b3�6۶8����pq��t\x��N  8kn��w[v޶p=�=�ɢ�W�ctWW&��g��s+�v������)�\���{��̾d;�;�������=;��%Ͱ!6W��ӻ+m�f<L�X͹;d�EM�^�q��q\���;{受��g�PC��
u>�h����ٞĒţ�]Ϝ��m�����C�ѵ�Ŷ^�3�o6�!�ێ��=V���n���5�Ӵ�j��T��!#�gr�tX�����+{n#u��<T��m�\��ڞ�>$���OX�ۭ��J�\u���Ӱ�؇���Û�����G�gOɷ޳=�;Z��k[���Q��p��f.N��1����OM����7�;\���w�:�O �֞6�q>��5f�8+�FĽ���`�����Pr�s�@�;�;�����\�=�S5�ɞ٢B�r�i;U��On���J��S��l<Gn�Z������O|�onl��H����ګ�m[͑R�1��0NK��{-δA�u��\�պރ��[���x�^��C�������qlS���❉#Go�8ۻY�n�c�VN��:���(M��۸�Z���E�Z����l�v7R�%�	�]��3��\εK������ˋ!�:�i�b',��]�=�N㳋;�ݍ���M���ۢ���9�N#��ǃH�˹�2�vލ{=�f��뭵l�4�b�E'cz�);�OK3��3Y�>�۫�^"�r����t���U����Le۫�@�ɬe�t�ڷm��n�.x���ꕋ)���͖k�x�n{[rw]���3�a�Z���ݸ\lc�ܩ� �y���8�v{(]���d�M�K�vr=r�۝�Y2���=��g[͎�w��gr^�O!\MW�z��@�v���z��]�P��u�o$k���J�ƻv��}*�ktu��q�]hɏ񶞍�u��!��E���O��|�����<v۔��&��cm�u�s�m�2gW�g�j���E�m5;��y`��n�����z��5L矠]Ғ��~�(��vͫhLJP����{X�wr�Amu�B�(@Б��n���]tu�X�^�^MI��Yr����r�P�6�����^ӱ>��� �V����gC;ss�w΀a'>.$��|����F��^���X�K�����1Z�w���2z>`f�]|�������ǳ��aV�p���bFJJA.A�=S׺�I�C�C{��%Y��a<d�Y��R.���o�?]'��M�y����$y����$��PD�G!���	]9Κ���vbV�����5�g�H�Rܧ��#��&4x���[��)����A^o�����a�&!�M4���Ys�����K3=S����	���v1΋v+�9���astjk���7����Mo-���n��"qmuǦ����ۂ�V��MKŷ�y�-∼��^��~�#�M��0�$�G��9[}�I؛���ǃ@<r��ہƪ�x�[4.pC�`��e���]�c9\�=��%ot�*�m�ܨ��t��;5v�MIu�z��X r���m_��m�PP�NV>[��"��tB�Ի!lýՃ+�e��q�m�Q��bXH�	J�A#���O���W�s���D7^_F�����\=�"���YX��6��R�{�T�z�ޡ(/���)(�@���chmjrl�{��v������b��޿G�o
�^�+��q�զ����>iGwܦu��j[����1��q�=*u=++"��J�l`��꼔ת�8����3��=��p&�UT+:-~��M���]}Mz�.���8���CB�ړb+;n���qq������g�Zx��ۧ�N��b2$$�""M����z9�p�u�Wa�yU�g�x���V�J>��7ZV��q������DUj_!�@��H�%�V,���9��ٿ-��t`:"���� Â���u��1��E�tcu��˾*{V��kp�g ჺ1���Y�Ki��4�%�m[mh"�t�7��n��M�J���ں��ĕ=�y�-��\���HW-�B��E�ϯ���P����!�oIʵ��S�h�gi����sh�����y=�hb��|J^<���z�A�l�%�9#NBA�d�+Y(��]����s*I:����D.������e;��,��E�48j���ntw5f��[?ձ2��� �g�m S����H��+w�YwJ�
�T43N�>�I���.��)����s8�ɔ/v��Q6Tӛ8k����<B/����1�nݗ��t����X���Vk���s�{c��m�����9��`����s�.�N�����]�[�lש��q�X5X�^?;}Y��M|U񔛖�R��!ۺ50B���E򨓥D*l�d�T���&�6^�Ͷ!Kkc�ѵ;ex��x̷.�p;�ZTŵM�W�M^����r>��e̬�ipO�@_�H�%#!$�O3U���U��l-���k`��0C�zB��kѠ�����f#DuR�s�-���qe]�Pn�'��0Ŵ/���>�|������m{$��v���E�aC�Azo���c=�Wo��,k9W
�H�XҚ:#��vX����ћ��[���Ľ�a&a���;���F��n�Sx���f�pQ��7?^+��`�h�K�ٔKA��a����lDk���6��]��ʹg�TU*��M���J��X�l,���%�B����<N�v[�۞^�G��/3���1u�ę��jfz�8��]�=��s�j�m��]v{N�<�k^�'�5�4����Ø"�I��Y���;>�y�ӯ�f
��x�>��!���k|=�ڟ���!Z���9�Y����2)Yw��&�!���u�p��	�wǶ�Ln��]�=;^��M��'�E�o����H�*��9�����y�+Ai�ѧ
	H;0�kљ9/j�{F��kf׆6i�K���	捯.�pZ���:��3q>���m:�r��}��k�^���.$�b�Nr�}Xz�u��E�E�t��sG���C����	��Уު�s��]y>�))x��vl}6�c�c\h�C�I�O��ңs]�=�����&XՌ�l��w�Fv@�!�����ښ��:)ӷ����ꥥ���q^���-��)�ɘ(Yy^��5�}��.z��h+�:����,���o>���%l��E�������B����X	=ۊՊ4 v��U����8�u�t��LY�W�V�k^s������:8�lb�����g�˔:��x��=[��=�E�=��Vݳ8�}�E,��+trp�u�@�}�-[%=�(�c<�V��n�g�8y��v�8��ܗ��J�����rnp�j������(���N-�]���wnϡ��r{#V���͹���ڷD�lan��֛K-=��:;�)�&؋�g�j}��v��5��u;�^7�nz���v{cw\�����De��2P�z3BM��������E(i��w����cc.Fpd����;A��}L���5}'�7�|�c��=��ܼU48~~�eڽ,/_���\����w���EJ�.�>�����1����,���]���l��<x1��^����!�0g��ċΫ��]vr[�Ct\�
Xj�6�g��͚I ��Z��}t���n�o�.�}�u,C�T�#놀����刼̶ݪ�.�r���@���P͙�t�t�>�m?���Ư�J|�00�N=��S����(x>�I����1:N�u��S���I�+*�-?8`��������:�m�7��ruc�~�Cdm���ύu�cӱ�Fh9�wK�s�k�%�]$u�[=��@p6�A*|Rj0��tx�b�N���PTPRd��'�v:C<�y4jV]cۏv'�O	Yî��T���	�,�Lț-HK�7X��t3{s��QΉ!��:=���!0a�=���fT���&�XK,����e�r��;t��]M���ӹ�K��<*�ˮor�v��z���O>���ָkub��3��0�B�T�N\w�L���x˺��=A�I$�x�sb	!�!0(䱜�g�3Ҭ��f�4�6C#�h�)u%�(��~�'n�C�Oh�b�~`�t������|�#�Z������3CVu�(���@��|��|�����6^`3��7�������t,^�Ub
�v�*��`���-��p�IƗ����_U�)�w/l�n�i��G���	��rԒ{�Q���hge(ƚt��[�]�4}�k��r���k�.4�>j]�z:�dn������n�rfxܫ�Z�ٴ@�ŉ���?FnW����Ө\G](�v���r�vx��fⱻ;;r��q�u<Q��v��ӥ�
a�B�6�&�hO{_N��[�* ���;��;�]>ŵ����ve���R�|dBs�3*��A�#R��<'�DL{ݔo�F�wn���h�e@�}��Թx�ES��#oň �+�"��mj���+t;%���,ϨY�=}h0pC-�[jG �͑=�Dkɓ���$`2@I[��lVn��7�+�/��q�1��n��U�٭��*���݄���ޘ.3ڨ�$�\3VFʁ҇��tCwz���.��[��,�&=�ͺ��B�]|��?F��wN�k���=%*v�1U����;hi��6���5gN��*< ��ϳ%����!M��F�cϻ��,�`��x��mҫ�#�lQ�x����;K������[�.��N��1F@�m8�L6���t�����ޢ��-�MK�z���;��}����|ٹ��V��+��w=���\A&���1;�U��G�������y�.;���lkb�)��ۂ���Nmv����7l��v�:Z'-�2��Bז�cܻ���/���^T^Z
WG�K���j�Us&�Ы���8l�B�lwN�c��x�x�(��U�9�m�0�i�wӟ.b�4Ÿ�K���0Ᏻm�ʴ*�ݱ?Ei�r��t6�|m�m���߬s�{.�L���b���t���A:⻖׳q67!�x���Ą��p:���.!Wv�8�A���7P�/��r�j����k�>���k��R�iȷ{���*!��5u�" H@�Q�{D5�6�{�OB�]�^]y!Vt�H|����f`����7@X;s=�ú�W!㽆��^j�^�]�뼨(v�Wd;e��]+���6�oh�W��O5����f��n�����M����w�
����U�<���T��b�"��ռ."��Ď%"p�o)5&G]��	��B�Xv���:ǯ�BE����<X�4XC��1�
(��]-�绦Oܠ�]e�5g��C������YM��l�ר�\�݄Rb�zٱ��["��	a&��`v���*����G����YyPH;=�M�
.�I��&���2�k������f��WK�0z��T�M7ٹ�Oeϙ!IN�l"�G��/�#���w?k���Q����+3I����TM���=2Y�L�c�WW���!����&9#F�q;�Ҿ���}B�F�	�|z��z
\rM�5ҽ�L5�kjv�7�8QR۔�i��������`�0�l$�6[c�S���7a���:�g��3;�H��3)n��Y�og%U>�a���Wm�S&�]di�m����o�=g��ìiL�Qi9-�e=A�(�ՙ���50֘�T>��9���WJ�>�L>"AN��F#��bCc��IckI��#�XL���:I��;�:,XX��5�e������f�5�<�]��T��wa�O/���Tai{���3R�KCU�����K_�_���W<�=�c�qsS�����wl�N�W��g���= bF��v�<v�Q.�ٛ���	6�1�Kv5����v�[!����K�KJv�;��g�{�K�uݽ�ѵn^#�v�	[�ι�n���$pLs�W��Kn�<ڍ����z�1n�&�\"u����N+ZN��³�bR�ǇK����,m,�l��ng�);qz��7�Ѻ+U����Fƀ7Wd�˱��N�콽����L�p��[mD�S�.��7\�Oe�C"��!(�W�~�(Y���8�'���l���w��Wd콋�}M�ۡ�ʓ�����ߝ#�(ݤh$Kg)��:g.����@��<u��y�'z�f8�Se-uZ\�7�Z�����ka�2X���A�틞������D�
e�
�Cg���_>�f[��6��D�r^��5j���;�m��4D�{8��3�5�t�o�d�:�N�$�+���Rp�"�-0,g`5b�?Nr�z��	W⳽*��6�G��g�~���«"܆�ب��es[�"�c���X~F�V�CV��ڡ]D�(����"��#�G����'�*y%�C(J�KLQ2`�Xuw�MlsM��,�C���{&���<��ŕ�ūD��l(W
���=A�;��[L�:G���ogs;��ZQ�Mڞy����}���t�ӯ=�ے�]��n:�~xO�n�H�Sw���5��/YW��vn1�T�/y��K#��b���*�Z�ns^ �ki�-�+�r��t�N�lߴ��Vq�	��a�-�E�<�e�\�����q�ݘ)����%<3ʜ�;�{l�kg!��,%��3�SP��Eo����o�æ�dVQ�%��}����Cl�}4 5H>,U>ht�
��%���}.	�k�.I�m+QZ٬��i�ϐo~@���ۆ�u����n[Y�>٫�٨W�I�~
��������O�8y�߮��Ɂ�h: �'�:�d_r>�̿���1����Hy�HW�Q�]H�ݡ$?($�8m礆^+��W��)k�K�>U��^:l�Qv�e�A�vv0�n)+�{mb�;:~��������:��	_r��R\�����;m��>\!HD�A�l$q��α_]��G��CO�=���̝zs/tU�a$Or�����=��/q1W��������H&P��AK"[����!<�G`��h8ٯf��iW4�pz���r%�۸���b�A�h��d�&4ݺ9���ݞ4-���
|���4����g����;�d���\,QS����JU�a��{�Cp@�W�Ϭ����RCAZ@��B	/��s�U���J���V��wj�����M�i}
�b �}~�����{�X'�Tn�]��E���0�,��S0b,a��.D�L��ff�F���bһ�FO�F���=���*���\��S�ʘ�Э}��M���P6K�sG#��2��}�I�L쳫 3k���q��ɜatn�t�i;p���$z�<�﷣k�ؕ�0�Y=}������ѷXo���,�Nn3�Q�la�K���!]18:Uݜύ����V4��W
d&���ɘ&���W04�K�00������R�]��e8%#��X�Ci����&�u�/�]M�������'�0v�k��	�ռ{T���-\�p���z���xx�1�1��3Xsf�7;�M���>{Rsrw̍5��p���u�8����c�N���������¤c�"8�.�h��s�I��7>c�����E��C�4�/��ʣ�gY8jWT����t���]����[à���U˚��p$j��+Dzd1� oZ[wR`�o	����;��]S�=ɚMv�૭�A��ͷu�R��}+#`��2Y�:��o2�]mM��f5om�΃or�xA��r��ˡ��q���f8U��� ����(�/4�(�f��T�	���B�gx�e�:T(����U���Єd� ^W�����鬾(ݹF�P�Co��'w���Ùօԧf�)�ۆY�j6��s��&JӱR��\#7�)Z���l/_>ӕǯz�oSh�Ez�|M�<��xI����L�dַe*-�诮�H�]���;�}�iݩ!���ܛ
�t�Fj�%l���K�Y�YY���y�*⫷��G��Ԯ�n�<ߔ�싡�;�N���<�����鋄�2H��T���s�[٪ק����w��$a
N|�*��8+繪���M
?LD��ʫ]���"	�r-��b��5�=u���.<ܭ5�^��o�����9���z�)�"���2����O�p��%��җ8p��B���U�@3d2�P	�
~�[�U��m@j��w����$wc�\��(=��+�a��A��d	.h?r/��w����t'���BO�����7� ˪���9Vp��q^q�l�aO�I�!��&�Q���(����}����N��VѰF9�S�繞;��rn��{���O�RP[w�ÿ_��޸�Z�y�[��
��B�/Z]�sťz�TʕHXE����y��p�Vw$l�7:㤭MP���O2�|�7HQ�vOgs<��!���ԃ~6���kW�!�/]���<n��Z��e�(K�\���� �����EZ��4 ���}Y5�Mp��b���/i1��/��{�*y�f�����J!gi_��&�!���Ho��}�B͑b�W{8D�����EB�*&��s�Cf�"w�L���#Ŀ@�4RS��V��["H]�:A��vc��R4C?m�v�@�Z���Hn��FPc�rV��6=fP�����.e�o&U�YW��=�l�f}�A���C���� f����v��S�u�?!��Y#����c�6�$C�khu�r�M�#�马.���w�F����]t���F-ӐQ.n�k��G�g�ÿLj#�P�J��C��X�6"���pP���j����ou��a8��@&g���ۇ׋�GyW�����}�i�b��UU�2J��-�P�TE
H�D��^��ݞ(�,�/P���;ǃ�=��!�A�s��ՌaWCG�Hm��q��w��ֶ��݀�������]�G�V���~_g�w|}�Y1����G_*�n�lUA���
h��,Qdzkq�V�&;ưI�"TD��]�^+K��e�{c�HX/	v�*�_1Z�*ƗU����(�*�=N�UAR�II��j�4J���ӝq�Em{U�B��8����$��X��R#����ķ��#LM%DwZ^��F1i$��#�Evoť�`�]#k4W�'��`�tK��E�J��R-�b4�p��>�>���m
 �Du�b��	p��R�#��Sy�V�:�JP
��s�~����]�+U�
�O�Rǂ��cRDiB��{U�İ���(-��đFs������NZ���-Y,�����8��# �w�} ��U��@��jEr�\�k������#����Idߵ�[M&D�.�VBܽg�9��ٜ�̆i%�R"�R*_'-z�)�**��M+��24�i*"&�W'���t\	f��8�J�Ǯ�q�ye>����F�"{���%z�Q�ĨQ't ��|@Y C��)�#�����q�ci*#��G�v����{%.�o7�Q?���E :����J�۵�1*6Z�z�B;�M���='�x%�,/�K���x�����{y�,�xW�hI��F�I�	A�9Ws�%�[�p�^XQ��t����˺�T!kEn�q�E^;q��e��nM�g�U��:A�Ƭ�������M�ŮN�g�c���p6�'�KvE��<����\��9�fps��j����0lA6Gu�O��<�k;�;s�)�ʸ7Q���6Ϸ���E�v�y4���\.[�[���$��U�k��w+���]��i4�⎙��`]r�����V �ϵ�v*N����L�ַc
���:�a�]�Y��f��w���"O�< �.k��~-Gu���et�E�ey�k�}wc��P4 °g��?Nz�[�pK�줖�˘���]�	��`h���^]�@�EDC�G�j]��p��a"^�=��Xu��ׁ;��hx����ֆ���&�p���, �X��?U��:r��\��	pW�	Q*#���ҫ��G[\̮���:W}ݾO�j$IQ*�^��m��nHo�.?�� ��*���S��+K3g�X��,�����n���*�+Շ�0b��;26N.����,�w��C#D��%�q���6�J{/L��FUͷd'�(����qP�tR�P��nid)�U�As�����['x	^��\I^�x�KG-C#D��1�V`�&G����	)&raL�N�fx�SB�P�!c�r�{�mQ��ue�Ւ�\[K
#�Q)����U&�"�I�R5@ao1g����$"����ж�HR��D��������g<��
�&�aeʏg}j�F8W=�\F	.w��.���M�$�J�$v��z%uu��|��<�y�bǰ�D�e� �K��w�{�`��s�e7f���X��GQ����l�w��ƽ,��������������2#�8�n��Q�{' K����.
�`W�ͪ_ �'gP�h�h e�|����|��_�MRCg����f��aKHJ����zw�0�II�"�̯dL��虒TҙsOZG|�2aa�W�:���R��W��#^����'�&=ke_��Kns�*�ܺp�_Ao�T�f���^��ǦU�Xi��ʼ|��ս[��<��P���'&�}��!&*��"u{������E��Q	p�k�9�i^��1P���T(�����%�$�~�G��kt����/90������Z�H��9#S�>g�3	��w�,n�~�.�̑D!G�'�~�p���[֣�^��q��p����E�w���],J���	����JHvvh�@�!M�� ח"��#�Db2��H@��k������"Y�ES�owťZ�j*ZRB�罫,�+���\	r���CD.o�U�3g��P���{樛���:\,J��x�4�T+}W���HHm�r��!B'�m|]_��P��Jm��e�cJ�u]�{�z�f{�r�iT�I	�$C�w��k�	*#�Ҙ��g�{qb\�޻K�� "�w*�>v�Ҳ��D�Ы������w�;[�\p�*�h�̷Od<k���^(hix�n�V��f.=Gm�װ��"�3G���y[P�]��h���{V�z�),JDĤIo/�w���%޸V��
��:��t�B@�B͟*R������8�/r�K�"���*G��ݾ���MϔD��p_����B�#©q�tY�z�F�2�%nO����z�="(XDpX+N3�����
'�Cё�z�Z|�\!Y��e�Z������ ����s�%7�?!�jU���}��@�
c��Rj��բ��p���:����z��#E�N0��qBL�5ٟM��R7T+Ƥ��^�ғ�`GM��n���s��k�I�r{@�P�ebϞ�P7Oz'El6FN�yg�[:�؝El@B�1[�RT�-L�y|s� /smP'F�BRP�s*+���aZ]����T����V8�n�E$C��_��Vz)�q)��}�ξ���N��k��@�R�Y(�#�P���U��\�O�D �u�b�w_��>�Q�i��PE��9�?���ަ��xh?nm_�}>��0��_#؄��y;��+�K�I�M�()!)!3�.>ns��#�{i��4Es��^��d�v��w��!a"(�"i��r��-*4�+����x�x(���1h��$Knɲ�oZVE��Vj���=8�of���n1�3\��C�_^��yhݧ�����ӥ�u�4q�"�ɫ�f���7�"�r�x�0��@i
D�ƨ�����*w�y�wo��`�xk�v9,[����T��D,���:��H���~f! )J��Bn4X�}�+Ia��j��a`y�=��V5��~��Z����uP�8W|ͧq"]�JL�_Z�"į�����̎ph.�(5`�l �_U���a?QS�(adqK���K��c5r���vB���]!�ē��Ms��0�:E
(�NE��r�A
�Kj����mH�t��Yޥ��xewfS�2*��K��BMJkM���H�R��#�&G�}d[Bs�E1�P���?�� 7=D{ě8�����:	�����}��IQ(�M��û$�O�j,d*��	��W�"E��҄����u��9x���x���׎�9�6�ݐ��#VK�d�wh��F��w-�3'^�T���.ƌ�Ae�#%�_6��滞��>��ni.�p��$�	������Q"*[uT�F	X��p	H�����U����%��e�E��~O�:l.\斕�V��I2p��׋Q��T�0���dV<�3���֑�0!�����y9�/��t=���i|B�͹�%8Y�9ơ���0k���`qՎ!֓�a�rr�A���٨���{�pN�I�&"Z�(W}��d-H����.߮����VB�aB�{T�{ҟ�k���U��?X`+�c�1U�C��0��� 
�m�pģ��F �lb��^L�� Ww���=g%y���e�,V,�
���p��2-"Ľ��+�\�W�W��1U��2L��(��NOG�_2����¡%ު�s<cd�iM:�p�RI
M��P��y>v�-�
�X���}��-�JH�w��j��#�.	Ug�M�\�XG����b�y�"U^��%b�T�RG�j/�>���4���T���F	Y�U8^!�m��;�51V�)p����.�`���0�>������*�뤦*.��}K���%�i��P��s�w��wy�ģ7�n��>>"�C�G���i���J�@ɐ' ��G�h@~�N��r�����T#ď�-z�@*!��5WPnGx��H#o�����H�:m���k�n8B��E*k��Ϋ�����)�@%aO
���J__R�3�E��g��"�W�RDǪ��K�=�J�&�Ͻ-����v{���q&��k��S�˫y{��L\|��K�ܬZ)]���նq�u�ɥf�nQ�(W:���ۥ��\F..�-����$�^3p�u�X�.Nۖl�S��P�Ż�w�y1�/`5��W7Gwhy�p6ع�=ru�V�3��C��;[գ���@e"�\�}��9ɸF���)[t;6�1�].0m�z�:�w.1�f�[�883��6����ݓn	�uVܯh�`ݮ۰�9��v�u�inqvNN9[��s����I�jC'v5�u�9����AZ��ͺ�8���9��/c��8G�ĉ2��t\,�9*�TD.{����z�l�#E@D�%&g=�.;ஏ+�=֒訊wR�k���}��&D�$żt&5�h�y4�t�S&���1F%��,��^�ߋ�a`�p2aXS[׵<,�^<�FZ�
�^�Ɛ��O
Īrav��V�kH�@�g�HB>������y�Xw�sT���D��B�#�sݕ�L�3Q"�P9�Z�� �B��~-%Y���Q�.x���?4~�˥?����3����M�B�>ԇ�- 3ۺk��8G�� 	]m�`�W��W�ÂF[�%��lY��1�'�(��8�W��}��;ݺ���sޢ �B�K��>�ŉQ0�	os<\%�-�ଋ�����+�x�1L�MAU���N���@6��}	'�}�`T UޱE}������q"�����_�fU��%"AS��p��M̨�i�����1.���PW�_J��b
�+�v��2!�B���Wn�X%�TM8A�P[��i`����$%=�����~?_��ͿW;��G�u�˛��Uoaj�x;&:�r���	��o��eƽ��ݻb�34uB�b蔉`����5U;e�`������*q	�LeJ}��p��(�jʣ�x���;�O�W��C:�V�?#������ʨN���):ڎ�%��~�r��L�mFQM��-�a��w1x��)��}�-h������؏b���9�ۺ7��<:!|H�
=���S�!W-�6�3��ܓ7�!����{c���邭�^���XD�J�{-M��&%#ʕ[�_�X�@�e�I	X�R%���ڟ8�#��/w.r|�fi"�~���%y���vR\�)����Q$I�ǔ�X���⸪p�Wf0I�\��'n3'<nDy�� ��A�nqa>���
���;�b�J�$�P��ݾ��۹�",���2>dg��+� �Q4�N(�6#�1�	Ox^���z�g<xJ���j0^H��)*#�E�w�p�w�I��;�g��C����p�D"\-"ov緪���#<�x���dC��߮<�J�E��!���0��Q�Ph|���}�.���$�*[�wܹ�Vp�*�喯�*����%]qwحD�$
s�J{�`�n����N�	8D8&&��O�}��wZ]�Pɧ�Z �J��"'��	WQ�}�G`��g����.,5�����V䗮	�*�.2���~�{��wǨd/_qϝ����6@G�K�g��W�Rd)DH��S��x�ԯ�4��o�^���!Q�%�'�W����G�+�"�}��*���%QN�UN��x4��c�G��^s�.(F���gw��/������X+�V>���Ӽ�ӆX�L��Q[~�<�qr��XE��#�>�u�KA��w��K7$p��O'H�4Wv�MT�&��&����b�H�X���x�HI���HU!@a?9����X��C�=�p�j^[T������X���62����O�y4ےT�9А��w�U����]1�ƉB��+$�8E��`�ܮn�z��(\�o�q6��
��$�k��'}�+J��K�vE
y��0J��%�'�D2���h}��ٷ?%]:��/_s�T �y�� �䠄�P�&�VDs�~-pZ(R%�D�N.J�H%ᯮ 0�dPm�}]hn1=�}~��UU�q�vR�	�J��K}���jBp@ʐE5g�@�Y�tҪq
{���^"'�)0�(U��d����BkH���T�
}��!�ً�E���݀��!ӄ�
@NH�����Ӑ@�@d	�>]{d;���p�5h Di �p܍�,F1�)Ռu��b�m���w	��]"&����؀nj[���;�)���BTA����z��2�5�EH�7<Zd>�9���8=����`��Ƣ��:�J��6��k��LE
*����Lj� �	��H"�66������
�^�q��5�����\#dD���ɬ�h��d�!X	�{>�R,M>t�P	N��n�h̘dF0�����3�D}`��VdXY:!B�p��g���V���!ٹ���a�V+�a*{��~Ȏ%��5�����H�����YN�D�t�>��hgrx��e�	�=���d��ܑ�����$���:�U1��4�6��~�9r��t�M4x��q�q"^n�y|k��:� ^�I�~��p���+s@������z+�L����g
�Pr�"�]����5��ih�JEJE�˳����N�R����8��� ��w���q�p��N���J�=3]E���
�����Z�*c�"��j�x�o�[.��y�F?B>d�5���dA��ޮ�Ui�@�K�1�䣷��V�9�~l�v��9"qnŬ��f]��h��v�<�vL&ϟ[oL��q�&r���������Q�jL�H�B4�+?U��.>�����}xEu�+���ZK���gJ�� ��w�m�"�������I�B���/�/�.��8,�z\&Wg̃cQx�>��[^���|+!z��x����4I1;Lne�.C�A{g%;�஧��C}�F ����T�h&��'�O�_>�,���]نG^�[��B���u�*�wX��,����� �'d,��:A���M�!\�6�L���9�\[`�vRF�q���鷭mk�#ޓr�֯T�Y������BRRh9�]�/%Ծ�����M�.S/����9��l܋*��)Ҷ�|  ��}��$�J"#��$�IDD�$�IDD8I$����a$�J"#���I(�����I(���I$�"?�I$�"?�$�IDD�$�IDD�I%�I$���p�I%�I$�"?xI$����a$�J"#���I(���I$�"?�I$����BI$�DF�I$�DG�����)���A\�0���8(���1?�ӫ��n�U
b0JCEUۡS`��Ȣ�rYjb��mۭ�٭n�{nz(��]ں�Ҵ �Tb��t4�ZP�wwV��tw��        �            P           
�l    @ � .|_m�/=�!�v�:�t�{�}������w������ݐ�� 7���{�����GݹW�ż�۫-���#�����u��g��}�;� \�>ܺ�{�=ݯ|��޷��/{�^��Рm��]+���l�ݯ�y�>�T> ����۵���oqݽ�w���o��|m�����x|���z� ���^O���3���>������/���)�J�yn�}�w����-�ݢ+ 5�   z 
    =�}���|�^��۵���޾��V�-ة�s�vi��u[��>���7���V�c����7v��s��w� �&� \u�x���+�ç��ZڳFض@{�{�����p� &P�������%�8^����}�W����	x :z�my��<s:md����Z����۷��v`�kP         p�����e&�{i�7J^oU겶��w�`Q�� ���v����_{����F��wB��N����QE� =�ӶM����������+5�҇N�{�x
<6�B�� ��� n0�s�` �;���tP��B�_C�z � �� (��}������ t&��Oo��  ��/� ���         ����pw�nС� ��tϰ�����  y�� �C�
s�c� ^gAG����7�7�P���� ����5�= � }(P�J���� ����>�{iٻ1� 6�w�����%�x��Z\mR��x�^�Wx ���i�<�)��z���o����5w�Ҕ�{
Z�P�h{�        �����cԽon���oi�w�����o7���� {�{����r���]���֕S\��5�Cn {�+OG���}ޫ����{�
xz��� +k^���@ �� �A��� �� >�BE�{�S�s��x�w������1�f�}�ۧ� �zN���������,�����N�v<]���{�����*D� OdbJT�� "��$��U 0  D�*��   jx�4MJ�d ѠD%Q�� �F�O��������(�FU\o�IUu�8-��o��y{�|Qܟ� I!%��Y�?�HIh$! I�$��� �$���HI4$! I�=?��W���cX,։�nfm�>r���N\���-�ohh�p=f��l�y��g۰��ïd��d&Eot�G�k]��l�DMOFS��WE]kI��'F��f��;�oeF_gֳ��q�!+ʮ��[3k_���W��\(�Q��Pؿ� o�)7V��,�d `��v���Z"�M�֠�����f���5k7wtk�.x��vT[����5P���Ȇ$����Rm�wS��`5��8#;o1�xn]����H&P��`KWsy;�Tc�0f�8C2&�zM�٪��#
wGp;B'o
���0�%dXK��0D}�3�#�*�E���D����Zܧ��܈Y��6��#j����U��N��"�t�CExat<�j2���y5�&�̬r�ن�,���Z����n�=�U�t���J��Ũ�&�ڒU�q9w0�Gc�$X���Mͨf����rҢa�{�Bʼ���tU��ѭ��ฌu)��e���1Z�1�M;�����d́d��/�z<ĕ�7�f�_RMPv])���=T�4�)�svQ|(ڻ���H�u��M��.����fRnj�Ý��1E��]tb��"�,�q`��UǴpL��h�á<�� 07B��JTm���X�+.��I"��X�����Y�u_�@	��W�K�j�b-��x�i?TY<�s���L-t�Ւ�r���Ef�Oc8, �`	x�u�c��E��Y)(���T7�9����َ�wJ[0�Q��f�4I������!F�i�E!N�+C�����G�d:�D�*�F�/����X��L��ةhN�@.����Y��\�J�SC/޶	n�KV|���J�*b��yd
��7��{�aF21��
���E�{Rڊՙ�h�j��<�u���g>��,�� X�N��C�{�Re�t�%8a����Fڠ�iSn���F��)$H2x��=s@zSU��ԃ�ҦK"�j*S�q-[V�d7�uL��Q �1�Wq���y��ў���+,�5� �l�:E�AZQ9)�=Zߛ��6e5�|���2r������i��f�6j�k���t��DC�5�kWʘ��[$wv�Pr�c�N%�m2Y����Dir�bJ��D������FK2����^�i���v�����R�_2�j�r�P��6�sV�ʌ͑���%U�p]���T�(1�E`F�"4ߊ(JJ鉁���-C``e�e&E�����D�m�ȼ�۝[���`�^��Z��l�CPi+[̻�Kv��3-X���F��k3 ;�K�#�vu��KÅ�`h5����˂˔�`Gr�#�Y�5۴�+7�^Ȳ�z��Y��.��� jF��Dn��6%�06(�唍C��:��o�O��͝�,��:oℷ�����s�d�f���n	��t،��ۡyR!�,i�uf5����\;��;>!���-�����= K_U!��e[G�ݱ1�D�f:���/h���>����%�G�[iȀ�G54�wt���ff���8Eh�]�kb��`?Z��!�>�u����Äد�%f,��S��
��/�s�)^$� jG�%�ݻJ��U�>�P�����gU�T�4۫9��ƃ,]I	*�eعU��{�Ib�㥹��6v-gj�2<��,"�̌�m9X�:�����d&��]H2�GH�nњ�Q]����*��Ԫ��A��J���]�=�S!dV�+H&m��
$�0*�aHAHՉ���-�z�`�Y�&at^z*����R���"զ�VVkç�NfNC���w�f��U���niF�hh�E�n�t0+sA�4���ͺzU����D3qK���ӽ���H&����R��h��6\�6���BF<߅�p0��u�tUu(�n��M���)Qճ�/ l0*��0��*��	.�"���-mʎ�M�&�b�x\ywW�d���9��r�3�!v���#a@f]D/l�E��dRb 
�{o�#6�qa�����X��+p�&X��P^!�s/B�c��=*�0j�1��@���	�MpVը�!�h}/%�z�)juyW[1^mb��0b��--U	����:�����k�C1��oP���7^�����nn�*'JK ���Ā�0�a�G����L[����vD�&}��b�Y��@��a�YrMz����w��=�a�.M&\pQ唺�5�!'O���voqZ�*�c��&�s%�����4��KJfO,`r2��	K&l8�j���Ŏn�4��d���u�C2ڽ �A�|�R>Zv�:�;k2�8�LW��C/6��KZ֐�j��� ��b��
��Koa�pc�WkU��P����fS��f����4��m���Ѣ��l�yH��N?f`�5�'7�$�}���n`gS��SnoHR��Rܑ���Ȥ9�ϳh%X`-jkRdAgj�Y��(��u�V��s�7���Z2��0MT/Sy���u�ӽ!!%�v��pRЮ�4*�F]3gVRwh�Z˄�s+(���Ȇ�֥u�`gB�ڼ�5nė�;Bu�X8X����{7$Ѩ��-��X�܌������6��Y2%��Zr�
 �dV��N�.�w��),f�iش���'���s,�aU��k.̏^=�h
Qwn�ܶMֺ�隽�ò�2m+n3A�['�Ε�A�:�]�g3�l!�7[��K.Jh�b����E�iA�&�\��7��$��'j*	����eS�6��3@G;B;�~�6TKC(�{g^����:ʸ�g�7������ U�)�j8�n!�	0F}wNn�ݐ�I��p�r��m
�GBJa?�9��$�tr���56�YW-����lRf�qe#��2!���7��Y�kl9�<��ɰ��#����b����DJ#bV�LoS�M^aϝ�0Xn���il�W��Y2��XO��#6��j���ܱD�	��*v̘�9�,��&�2/x�pվ�u;�� (A�G.��z��}�@*����5��z&ռ���d;��E��3V,�B���ƶc�>�mm ݽ�њm
�3>y
�F�Vc5�XWZ��
g�Br��%Ö�T��/D��u�Cs�U����bcf��hf�M�7g��੺�M[7ŷ}�M^'exP��+qӱr_�g#�[�o��s(��ݧd����)V)�axnY�d���tKr_�i9��{&�����Y+pr�c�����T�S$U�4q&��1��X��mg�1n�K�U�Ǯ�sV�ё�ݫ�fm�k&���4U;��ۥf�=qAm�I���g(fi�v�
�O̨�M�r�ž���FC�=�fx��逥&�!����G���<�I��LQ=: v��L�rSXw�b;�)��;
����c�z�C
��)��{QS��1,Fka:�_n�v�/�KoY�}���StFP��y/mX���;��{�m�*x�Mho)n4I������%qI�6�_�9[��IKE/|kI��U�����c2-�mTHnYW
�Q�ś�g Wr]i�+����i	�+F��� b��U�Wz,"�j�k�^�8��6�'9R�p�;�X����m�;�/�ʾ�3�TrK��22���/g�u���%mHK]a1�u+�R���p�xc5�n�щ���N���qos�q=�Q0�`��s+z�u���X���>�
</-d��*fS����.��=h{�e�W�]c5F�5�G�f"5<~��v�x	1�J�z��4[�����+��_,)�w���0!�Y+o3w�LF;":9��	~2�[�=�m���-[�˨W�kcݶS��pn6qسq/eBj�QfP�=��VE��[�'R��g����%�&F�Ե�
�qb��q�M��*��{a�K�%y0}.�0�JA���te��k1��.YXߞ���I�j�V6V��q�U/L�:����cVX�M�HY�m����i�8���BP�4|�G��kNcoo�1e��vZ�L˨PS��7 L\&��"��e�Aw�Q�lF���;�u�T\ֵbЕ�q���Z�*�m$o)ϠL�y�	�.F4-�p��0-�𩩍��n���N�:� swe�y��.- �̈́j�nXk���F�4Ap.�(�b'\4 �K%��U���w�Lc!++C����n�o�h��ޅ�&Bp; ��Յ�R�nذ+i�XS��4U�3 o�aS`���KŎ��4R�[^������)J)�ˬ�J�Ap��6�Ĳ��\�2��9�MӕU�wy�qrrm����3�����ԘX�&�B:Dssw���"�&U�"�#�ȥS�^�A���;)��2csV�P�X��HS��Ͳ~�2��R¦N��w,ZX��������%N ��F*��(T�.��y=mX^3d:��:��F�-Vl(wVA�\���Y(�6j�� �V��[ې@t��aͽ���0Z��U����JG�5�K���yg�/	�9�FV�6sEり؈�3L��
�b̀�-�:���W��џR/A7��1�[3H��7�����M��:t-���6���(cp��^:̙�Wj�¶LR���B�6贻�M�z�Wҭ�2I$�9��g��.좿��6 )��{�߶멛k���'�$;W�{�ږ�3^��ŧ�b���'���7$��V�y�
1�bF�m�2ò���2�Ca3I^�*�#Hf��,[ͭH�F���t�]	T]Ѿ�U�v��+0�.�Rr������ma�p��[�����N�l�KRhǭ�k��]�_�Z#t�g.�m�e�4wF(�ޙS�{�h�d]]]��U�V`�	�d��Q;���S;J0Xz�h��؅7��#��^^�M�x����l�A�����)VD�[�;�U��
�F��R�^S_�`)�o��"���sɨW�y˙-F��d�R�q�Z�+���˰_��Ba���ثF��S�-��#=���Vx�2����׎����C��Z�Y����GN鷵����z7oU��Qƃ�E2RAMf<E��G(�j�4}N��W���L�Ywpє=����[����b� $���lp]�p�80\�˘�����;<r2� +�i�L��7���#�;�%2SRw�����aůdz���;� ������!� `O�F\����Vm��đ��� Q֌ӈܩ�,��41�r��:7�H)pK˕ulJ�X�E�gɩ0z+Ȯ�m0�$,�L� �,
�i]]�eO��;u	V��֒x���fV�5��M�q%Y�����Y�m�E��wwqc����	�bR�1�m�[yPֻn2)�&%'@�5茸vh�5m��є[ɛS48�wڐcm�)�ৎ��5�`�1����{J��ذjz��mVJ?-8
���-cr�8�hb҆/���x��n ��D���a-�S*��@ђhKp%�p1 �����u�ƹHb��N�	&�˅�%I� @�+eb�(��-�6Q9���n�q�BIG,c����� QGd[��2������j��#�Q�wzpi
���U�R��P�vU�;�%���A�3�p^��dk]�l3WwJ�(Tp�@���32��RBcǶբA�D��,۽��[j!�����N��M'F���3G�>����h�[q����%��؆��.��fF�˔��YFstL	K9F>�|ο{+n��ћ��H�qn���'+���nE�aM�j'�[���"�{ձ�f�9��&b�̝01���̳z�8���$��n�]L��Ѣ�;�RP�#t3�(��9%E�?n^�-�&]�Vl�5w���"���0j�q��[a�4�8�*�ktũ�i�-ܠ�7O��lN ����ݩ����7)�d,���PPPVm1�Ty�d:V�f|̖
��f�B���nؑ9R�	n��3\.���u��v,fڹE\3$���j�M��A�����-G6�FP.$�WmHY`˼�ͱz5�2��u]��5p�7kh��5�n���e����k,;R�}����%���S4Gh�x����5�tj��Ϊ7����lu��n#7t��S8k*n�NU��$B�G�0��Шr�S�l��(�w
1\٩��#̂�ؘb��Q6�Jb
�k7~�f|��l��@[t��'��d�1?z��xM�ufV�b�@�Ўt���kU�R�4 96��f!�9��hf4�JA�o��>���
�0�f�VS�$1PA�4�p�ݥY�M�`�Ub�����,<x��V�F��#Zь���劖�lf�-Pl�s��hz�`T�>t��F�:�n�-x�{qJ�:TB�q�(��K�$�cj�Lܖ�"q��F�� �5���GgVh���q�(PP^K�g����g-��;�aٵ2eMfvE�y:�]RI��4'K������w�R_5�k�a4k/\��CnT�(Y4��^�Px�i�5aQa�Og�*/	�w�T��@�2�vq��`���J�e�{@��*̪�Cb��1�	HE��9a�L�8��Ex
�u|�r��R�r�

�xA&Q�k.�yv�{"`�HQ�ʝ�����)[���
;��Vª�����N,�bLj�GLq�ې��/����sn�'yHZ�ה�e�ÏGT�3JuS�ws�&Um�7�fM�m�WyG��W�ݧx�<�CW����/0�,����(��䗂X���|��F`(f�lؕ����&Q����)P�ꬣ���y�����*E��$�$H��a��R�c���p�>D�����@$�d�J� kn���nʻR��lmU@@�WF�h6��U��KX C`��(�h r��*�*˱vq$��4�퇮<X����x��v��[n�7
����.�W��p�;pu�]�tOF:�YWwOX͎�{g����x�fۨ4^J�"�Ǟ{n0[x�3��80`x�q��H��_��/G5$m�ӮoQ*�u�)"r)cD̊�����	��]���F����zۊ�oN{l��ݝ�@�����#m'+K�z{'��A�8�j���r�=�}";��yg�ѱ�g�7Vƚ��=so���}χ����],�Q��'l.��p
�m�m�pQl�ڞ3z�ɧR��#)x�M�	ň��:[�������qِ�v�I�n�'�ڍ��k�l�ܦ���GU�]�k�];�]����w7!��v�G��`״t=��H����^��8�@Wnѻ`Nwl2�]��]/!��7�ь��!�dx5���j�Z3�L��7<v�v�����Z6g��⇊���W�#�k�G&2q�猃�:5�}��7w���n�&���Mm�䫈S�+��2��u�<n�9�(��.���{
��c�{ퟱ֝aha��v^:�yH��v0�a�n5p�z���S��^�9!�R@/o=�g�d{%��^nX�{]gݠ�=snl�v~�������3��;Y����ڮu§�i�6�ض����^�\��89�c&xNQ�P�b/<�,����VН#���jP۷a�F��M�m����k6���}���{SV��on���8ܯJl�ɞ�Ǚ�7�i�l<�V�<�][W%�� 7m�y��=E���uGQ�\��ʪ�rC���!gE\k��ol7=�C�nqӢ�����Q�.�4ܤ���6�[�9���jш�e<��r�㦱ΰ��nۣ�R1�E�-�n2�V���v�[�e"�6_k�Kr�d�6ByQ��vOya5;l8��z��`�Y� ��v��"5���mp�BKe�z8��1��S���'�s�'��4��ݐ�N^Ztmͷ�X�)�[>ׂSu�ֻ������cv`&��B����8/c��<ۘ�b�n��<��{;:����6�H�Y�ܗXrn��lZ�:{#�<[��NLv��
s�.&yxWucg��<����{n�h�ճ�s�nu��Y	��3�^��k����m���\rI�m�X���]������̸��9�n��@]���<3`�E�\���S�s�����5�ݻx�m���[{�Aٵϲ��9�bdIݮSpXgn�V��l'���m�δ.�u�=d��J���l��+��N�1lm�:��[�8���;���c��{=��(Mn�oWV�{]�p�H��=�5��ơz��]����ϺC]��z{'!�C��1웶�V�7;�4��S[m=�Ec咺
5;f����9-F�˄��GDd^��	�9�nh�X��r�O�x#A��[� �;J�k���s��ݒk�g�E]V�+���{Nۭ�Wn�u��f��=�NkIc���v�m�kf.��;�&蹤m��n��`(�	�:ɕ�v�ݬ"`+���t��o^�L�܀f�ɞ�;�2`�g���t�Og<��۵�I���p�֚��xTc���v��^S]p��mY;E�b�P=��������JWr�'�,=��H���k=����;6�v;r\ȕ���v8>�����<n��F�Ç'��ӷ��X�kc��k�����w��'����֏{muݞ9����Sxvٌ��ϥ9��-ᬖ��'YBku�X��{c��g�]���y:�W]=��B����v���cr	��p۳s��`J�ƶ�-^l.ojrj���ů)�{(�v�����Z7F�`����ʡ8�7�&��H�g>�ٟ�;���=a�խ��K�"���_-��Vw��>:���n&�XG[��vVڬ�v�4e �9�Ws�omN�lF�� ��Y�]]��vݲq�9�;������{;�76)r����v�v�q�:��<�WQ�;I��SYt	��'����Cr���ڧ�O6��m�[k�i�b6��L��^�f�cq�.�Æ�խ�m�v�ܹ݋p�-Ӷ��\�;s�]%��:svݜ�U�$ƅ2Wm�R�v�;v�QY�v㷎"����̺����d�=����xm̝w]�x�m����>{s�h9yd���zrn�n]]6�dzOf�q��G�	�ŰF�Ŵ��A��&=�7���9�V����Hp�ۃJ�C��u���lU�i�q$8���6o-��Q���9=\QJ.�e���=��p��8�g{�L���j�;㶸$g�����6�n'==�w=��O'=��o��?p�۶��5�IZ\��uÁ�kUl�{�	v���7Os�QW��le�ok����6.M����eI�3�7�Y�ܻ���+U�E��\�tnv�c������Q`{�����cptG��n^�8:+����h��D\	Wn�ƫv��x�;�\��c�7ӗ�f^�z�0��f��n��zX�͋g��y���&���i�g�;��ݵ�OH����s��qG����ٟR���wk���s��W�����x7��zgR�
�Msr�v`=k��Ȼ+c��[�������8�8�v�wn��Lf��۬q�M�z�q�y�1��K�5��\MjY{[��0v�[�E��k��SI���Vf���b�=ې�v�c�z��[7]U�����dP��g�/W����L�$:r%�uЃɦ]�R��5+�Te�ѹ73h�v%W�w��Tێ����d㎳�+�7�5�d�j=m�>���6�s�n���4b�}2:� #s��H�P�
�wn�i��O�3q��KmDǘ�=:�cjݹw��jا&��dSp����a��x���&��[��d�[�\?����9��e��݋���øGhy�}[:�*�L��ݭN���\j��!+�N�%����v��n���u�.w,u�1yc��g=ag	��ۮLt��k�r`��MQ�;�Tf;X��v��¼�t�B<i벾�7��+g�9y-���^��O)�����=D�q��y�q����777g`�;e�5�ń�gǯ/�R�\��[�OS��픛�N����i�sŷM3o^{Fwo6�緪�9c����5�n�`�f6�5�yͳ��gF݋���z͗<����.�ƽ�ա�39�4�ekg�V���%���j!��,[��N#��[!�-r*��l����S�ѶSV�f�=�#�����7a�<�[Z���ۧ����m��n�]����咳�u����r�۬�k�V�W7g��yC�Aj�n��8�z�qvG���vS��m�q�����a7mnn�\fGf�i8�x�ֳa���/:�Gd:���b�gu�Nu�$�v����u�(�`GO8Y3���n��ev#����x��Q���7`1a𒎓�^��Ǎڬ=��;�7Jݫ�8{+W7I�+5�<����`܇[�@1y�
*�9{@���FNՐ��k���u�=>8%0�L��w<ڼ\]q7nN�t�uq9��z�=��T=i��f��k�ն�W�r����X���pja�%Ө˙�v_=��7m��g\��8��e��k#�<���i���86�G����N���SWl���8������`R	tR��U�3��;�Y�Bn|lQ�Nr�j��/]�f��j�m�+�ô=�l����i�O%�nw=t�y��mz4v�:A�$�{;�^1��EN�6g<���1ш��0c��om��v�}��ì��p݊dz&N���=��-�pp��4����ZM�ٷ��fn��&��g��힮,���v䎰�s�:��7�м�u�Ɇ.ض��#�ͬLv��{m��j�w���V�u�`{�5�<ľ���^�Wvn���cwbZ티����=p��7�O1����b�Og���u�1�Iod�$0�����٪���<�[���"�`���G��q�������,	�7^�^ ��l=6���;vm��\���wd��-؎ѷ!rmN^1��Ǻz��^�8�f�خݗ��wKr�z�'���z�u�k�v�4�k��]�6��N�$�H|ÛM��n=$AZ�ћ�l[{<�v;y��b���Ɨ���������R[�Ս��F�(�M� 
ۋlgpcrq<(���]�k���X�^y�d	'�s�3C��v���jj;7"�G���c33���nx��tw��>��mq��[���ݻA�x+��m�nA�����5�\b�^��7`.���i�f�ѷm[v�+ݽ6rۢE�R��X<��������x�Ύ{N�^�	�۠�l��;�÷O�( �ۧ�WE��]<m�og�C�րO<v��@���p��N�uu��v�ݷ��#�������y˹�<Z��:�c�j����d|;��l�ny��Ѷ��� �۶ʂ}��V�;NTDkj�Ua�筹d��=q����3��.;VT0�#p�]��s�A�!���J۶�m��E��t�m�WN����N�yy04�V�aw�z����Ďm�s�vw\t�{Htxm�vGK!�8���pp�,ȻGlį�ނ��Xx�= f�;\�y݌�g�%㡬�b�n�lu���=��tj�
�uu�l�����yk[��Ř�q�#��v�c=�1�H�C>�&�S��D'ug�ܸ��v�3u콸1�m�䆶��ݸ��w>���Vݐ<1딷G8u6�Q7���(��^��v�dY�L�ۄ�O�v�q-1��ru�nk9۞�M%B�7J�󱻍����z8�c�M
Hv晽�Q��D8��
�;=����n�s�n6݊8J�ڶ�Okр�;�$C^^uv���le��)�WJ�^p���u��p�����=��g�cnn����~�=�}�݉u��sns���6����3�;��V9��cq��"����mm�QD6hNK�R�ü<���e�Ś�b��6\�=������nͻmVܳ$�2��$! I�R�I$	/�!kZ�ִ��������Ls�����)mj��I����k�l�l�cn:����G7Vm�֛��H˸�'\tj�A�[�O%�;zm���%�Z<;ppK���<fݑ�]��ך^E�QM7G� ;nw9�nG������tl��w\���f�Y4u	۹6�p�,��ht�!��7L��o6s���睕�:��fF7d�8�\t�<�"+��!�Ddݻ8�ݹy݊��Oi�����з;��rk�v��8�ʓ��m�7�q=k���w=��pѶ:<5mv�<�5ה��BOz�Zѭ�kj��м�����f݊�Ú7;�y�y�[�z�_I�u�G!l�:��cͫq�ۼc�W^��s�6���4��n��F^�[��X��J���:kv-�+��&�ۏ-�c[�e��ܦ6��6��)��Ds���W�n#%*n3ƍ��v���}��J:z��;rv�V�`5�ƌs�1���xqؓ`Lv�p�lo4�v��meۅL�X��6듮�0sю۝���m٥6�8;:�lX�e^����k�����d�C�m��q�h�sarٻ;��=<ݮlv�h{b�C���[|L�1��v�<>kgg��'��ᵱ�v�A3��[h��Yw��3�n��0e;p�laZ�˴�u�<��m��^w��e���n��:�ɧ�E�s-����������뮛�*4\��tg��E���z����oV�T�X���*z�z��.�n�s���"����9�\0��J��g����C���5��۷=ݚs��JW�:�VϢ������!{����n\dM]���v��*8�P3���W��l�U���a3>6d��.�1�e88��9D�
�P���m��v��<�����u��t8ݳ���8Wn,v3�g��3N��KWmƥ��bf�m��l{��=���[�@�*nM猻��G�˝�O�k�;��u��N�Vj��n�{hhx�.�e�wF����v�c�������Ϭ�:�!�����=�y�Q��Դ}ܐ���4 C`$� 6�6�bHHI$؄$	!��i7���KZ������*	4��1�mäbx�۬��u���c�i9�y�̚5ۃ��Ƶ�5�Y�;��۱��'k�Ǜ�N���p�4�r��q�np-s1�Q���{q�n�؅��
k�cu!Fnj�q�۸7;���4�rn��p5��fNx�8x6ws�-�N琮��]�`�%�;��b�	LZɷ���	&���ë��\�ě��^�x_vCsۗy۶�M��xT�*gx݅ț������5tݖZ�������s�^,s�9�G��>da��^,?5Y���Ξꢾ^� H��.�����bG���AI)��C�q��]�W��nnc9�5��j�6  �j:K}�X�P��^SL�"��Ô��t0R��V���=�`��_�[�̸?\�K˙�:fN+Q<R�}�Qy��s%��ގ�7g���������4-"�A��l�A�L����S<s��2���r��Tá�ٕ|BN�O3ܹ��9߻$�〈��H��.Yz�'�<��%�QYO���F��ᤣ~���^�I�^SA�R��DJv��>�ڊ��c���7F�2�T�8��ᦃ=�[��!���n��zܳ�lWv�d�"-����Dnv1*�$%E
���1�IO6����8�d�$И�����?
��{�o���!i��i!�m$�xR������<�l�`;;6�;���-��dg��/�]cO��ڻ�
���b�^f`%���R��,����5	��:A췇�J�'�_'�ɲ�aE�D!� t�G.��� P���M�s��r/��b�O��rd�s�]�����ŵk�bp��n+�T�V��~��yJ�TE�A{Yk���|�˾,wY��6q�������˄��&�O��S���D�F��
��F�zû�U�Yuח ��Ī�ٽu-F����n�\b�4>��O:4ǳ7TC���5��+p�@ �3@�!&�=k�D�=�z,
�> �Y/.����w[�v�?2{�m`��{f���UPf� ���k����^2a��K��r�MŔñ�g��<�m��������v���0,�`ե�le`Ёؘ�/c��N������=�.@3O�]�ƥ����owm[���'�S*,碤���&���`$ق�"��n��krc��C)�4�Y���y�t*����7b��w��v{�쿰`v�ܾ�E�^�J��ђv��F쨲!�y� {9�T��!�B6����s�����A��}n�s�d40t�h�b;�5lv����;�-���F��%�P���{F��4̅_+Lǜ4���gu˼�ٶ.��+;��Vj��ٷ���doq!���EW&��9F���<�-b�R�A�����AaZ�Q�0S9�4K��
o���mVl� Q���4d�������>>|fFo�ѡ~#�J�M�ƓD�,�m�S��0��Z�Y@Čُv�tfT���ȭ�K̖��h���U���s7�,ơ�v�
,��ms7����\5c�)e�u�x:1�ز!���6uy��W�;A1u�Ώ<nqѩ
ȜAcl��n��	>����7��b8���͍ȖnT���w�\�f��w���`B�$%�>��RU��mM�#�T��) �X��ت�����3���w4|�P����ڱ��U�k�8�4n݀�^kܜ"�.T��6LX	޵�O�՗�$NwX�Ke�bc�Ɲ�O{7RJ��ue@n�����3f:b~�֡��}���x��)�5I�8{��$k��OI��1��鴝Y�X�lA��Қ�2�s*���=(�ܷ>�E���}`ȩ��q�ۯM�le��8�b�yRr����w�����FX7 �V�����*�p����#*U��Ϳ�_�� T�����\�f�?w�ܙ�L��L�f�m�	�a&ʂ��1���N����w2d}ɣv�}����@	kTI!,J���'%�X��X}��K#?]�tY�7G/qK�Q����Z5mvj�y��'���DΜ�kp�6֭�L�9".L�I���������� �i��TÄT1�Tik����ǥi�����|�R{[{'�*V��R2|�����mz,Q�5j�VBV��> ��Gy�T���z�C�1�`�Y�����p�k� �	�K�W��x�Q�x9���}�jm-� ��9I��UJGf^�7gI�7-wnyU@��2��|��\~#�}w���}DC�G��meq�F4դp�	�����h�
�4�dr�3\O7(��jA1,�����-8�1�;5r���Cx������[�"��M��#EaiӦ�i�w���9�o,~;��a�=�
T���T���ԃ��fn���F�ӍzblY�"��U�\�{���u`�8U��aK��:����Yc�ds];�0�n%��R�nut�[��ۆ��\��\Whl�����W� S�	Q�"nR��v6�C�s�%5��]V��ۉK{j�e���j-An����g�������*9�=��rطv�t�:�dp�;Ge���w<��zun%�j����ݳ�­���ۄ烮��mn,�Q��%��ͼp	�e���y�u��[�:x(�v�&�ӝԍa��OM�l0�'<�I�3�1s�-p�0l���u���q�Fֻ�Цl�ц���:���/��]v�\<�zܷY�v�3�
�i�k�Y�z�0z��`�޵1����?�K2m��1�5���0�k��z�y�qJ�d�Glb�,�>�i�WH���,��
��C�.�pՔ<ś��q��>����L,!r�j����,�=xfEY����\�OjS���A��lբ������K���a
�Z�r�T�%�1=�˥���+;:�ݠ���1�k�c��$P��I�x� ��&��
Րd�����ܮ�S"�E<�ZrOc�k���+x��_��QZ,Ҡ�2l4�!9�>�bː��{���8�$IF�6~��ԇ�Wۻ,K�Lz��g��,��^f���,��W��1��:$~��lLz���+�Nu;�d��i�z8^���������#gGr<��N�<�q�^�bN��%�sеwￔ�΄�͏��FU�N~��gR��>�Cq���o�r��kݺ�_EZ�F�~�y3N���r�	���{J��W��Խ�90δ��s,`��4��\�h��	-�y��m^ ���|�^G�:,�v21�t��`'F/s0�%�"H�n�חՋZ�|�I`�e��/�s&"���I6<��{��_ܪ���ʟ�
�VW�0��3j�p��l�����=$�BR�-..����J�^j�ؾ���\���|���,��D�z)�vB$K?��r綘Σ����{+�h�PA��6�Y)��dhi�/v�`��R�;6��ˡ����yLg2���l�;�9��٬�HU�Kc]�0dIJ���w��y��p�S�]݇�1u�@�t�%6����>f�4�V��e�tG�A�g�G�}ùa}�׶2t������6i[n���>��[�B�lY���Gw��7��N�<
ny�t������a��ֺ��u�����۵�vE3�n.+�k�h�h�����g�\�5HX�����f���h������:cFwq<���׷p�c�W�v���^̺�]��g�jCPD�9Cz�%{zj7�{�5�����\�y��V�����Y�L0ٮ��)e8�!\2R���ܗ�>�?n&d~��܇/��k�5�ɻ!#uz���O������!�?k�����A�Ѹ��W�[{%I���>&�������æ�����&�ZJ�˭�v�ڍ�u7���F�d�0���S�#��힛]�]w�kG������W�/p��4HD+_͡�4 SO�Rx���7��xC�B 6���؆%�Цl��AT�]PV�:�AB�,�U�y����Ǆ�B�2�_�6�Tv��_8_	6^iN�U��,C�ܑ��� TEH
ܞ �(�sg�b]�\h�����g8AݛT���g��^n�r���oٵf��j��[]��'6�0]Z�4�H~%匥�t��$KdQd!<�ɫ�<��mf����{F�źr�x6y���gFx�,p�������9�v?�ۅW�~cE��y��{�?[���0�M^ܵ���b���*m����.Vaƭ���
��*erf� 'A�RM��c-�.ɿ��>����ϴA���w�-X�iLF����&��ӥY�v��Ǫ
�˲���4���2ތ�M��>���W���T�
_4�rP��'flٷQ��fR.5�C���9!���o��.n-�á�vlx�U���$~@�8�}�Z���Ȗ'v�1��D���[E;�Y�w�.9�ڮ�s�M�(�v��i�6I�&F���F�~l�K[:�Ѭi��"�՟�����̵��!��4����m]`p�Q��t{�wF���a�@�a$]n��F�ʹ�ց�8������P������`B��Ֆ f�W]��Z�K��s���j�� � 5V>H�LUȴ�PK�Z��2�Z����>�c{&���@۪�'���5�����CY��:����y�-��+�`�[�Yu8;h}��q�QZG�Q���(z���������1ǡ�����YZ�k��3�e&®�&������Jn�fd�B�d�4W�+��_?=\�����ϩT���.��J��l�?L���5H�/�6�-8Qb����63�����o�;��]�X�_��+����[i������(�L�I�R�ZΒbor�n�6�۪m�{���P�d9�����ZC��;)qM�fԃ�H���S}gw�z�8O���FMՖ�될rӂ#ўٸf6~����~O�UB ��7�Lh���2� ]�)���U<a?HjƊ�?]��SoD�W��51��O�(��I.�Fxqv �9jH����Y��B��$����0SE��e�}D|G�|B�MfUe��-ʚDJ��h�VЦ)g�A\�Դ�T��}�ަ+)l���]����F�!!)�U�0��y���.����hz����}ln���N�yuv���Θ���ǬWoe>﷌ǀ�;G�8���ˉw|���#�u��Z�����RV��n��=lݨ�R����)�.�X��;��+��#7n��/)��+[v�]ѹ��\m��p�A4	�5I��]�ݦ�ݮ�Ѓ��¥�A��m�=�<q�T�6�4_����S���u�s����%�;I��S�z���u��#>�S�9z�K��d cֺ�6��Ʈ\5��hQ��]h�yv<��=����TV�����Hp�xKkJQ�8�*SmŘNn����K�:q�m�=v	�Ӄ$�*1���^�P��kٻ�x��G�N�9�������@����7��i`k|:
:EĈ]��R��V:�5� 3���F�P��rj5�dI٨�H�<��5�e���cx����e�c��S�_~���Й��5e��E��:���������0�e��5%QL���F�I��VĪk�}�ù��9I;Vo�W��[TU<��]Ql���9��3&�ޡ߸f%�5[�V^�~X������Z�A�r.�m���㲴v+˦#��ߩt9txB�AX��.Zb�IA���>�#兊����=N���_;������zӚ�EU�#��S������_��c���,,f0`��Q�}n�_q�0X�Uq(���A��Q�%���G;�/���5��7dܐz��sC��f�5�ۛ<s������1egv����]���\0Eh�ۥ��BBR&2KU%EeX�tRۨ�Q,����+p�f�2��k��uǏ�<�!�nu��/:�A-w[��> ١��`�Ƕ�&�>����xVi��&��O�1�S��]S���W��I�u�V1
r�۾��6��3{�}��(
��^֬X�л�b��GL��膶,&��5����v;rt�x�+F�;��p1���A_-�`h����0v��Gާ׎�3D����;�'�j�L@�(�H ��ޢ�A���kj��.�V.�9?����@�lX��>������b���8__���gY� �A���!B&hn$����֝̓q����e���9�W3��`�z�����5�s�>k�Ð3�Q�zɬ3~���Ʊ5_}
��H�Pv�eKl�}���3��W�_A��+���D��/=�fPcE�n���O
!�T�0<5L�s;6D�|.��j;X�[u�9���ݞ�?N�^�u1i�xi쀽n�̑�:��qk�k+`�)�.J�g�˗�뛌4�1�|�]5&�]�׽����K��n�S��1Ʊ�s|�u n6�Ƶ�껸����<iG{s�^�J������Zl���u���ל�[�mڡ혩,�p�hw��<��q�g�\�u�&���H1H}����M���'�3&1�u���7����@ܐ�4(Qs\z�(�D�oi��ӳJخ���9X>#>�R�I�?zRWWr�2<Y=vd\?.,��`Kyw{W6n��M�+�/."�%w\����ql��ֻ;U�'W�x�6n���]\�L쁰�:�-\��{a�s89hګ
v�!fv���s;o䦞U�D�o�Z�ㅰ6���	\b/,ڹ]�����/������e�S
]+�����ث3M耰��7l:7걭}Y�����@*��f��ڃ���כ3�]�@�U���B܅��elْ���v��;�#C����I\l
�t*E��+�l;b����a�����#����X�׻k�sr��ōr<�Ɖ��+yp��vo0�z��뢳�9c�x��eH�Z�
�5�N��g>��W���� �L$UYy�T����`X*��������I�]�KP�n�&���L��E�D��L@�<��gZt���ר�拦f��:l�ׯ��RTA�P�-��n�z��(]3��PQ*+{�R^S��:��[f�Z?�辯+�lg�!���\���iV���wUY��_����%zD�I��L���GC�֡f�{��[�����[��zM��t���z��������T�<��T��]��JL��{|\�C#K����!��ܺޅ(s����ñ���ř�	��mC��cĩ�ͩ��Eܥ��o*n}b�Uˁ�����F�V�f�-�a��4�ԧ�5�
T]_Y� ��=��!����c8���Co@��wndﺻ5�G7At|�칀��=rW�^�kZP<�;fj+�g;#/o�Q����7��W���B��볦Q
�3����z*j�n���!G���g��ƻ�N��?d��^��11�ȩ��/MlU�, �����8HXj���y�U����}x�=OE�n)�לEld�6P��:�Q��*x\Awb�(��w�&9j;YȰ�+`��]�0��(�:�F?Y���9�mma���e9i�����|����q:Z��K���a;�'��l�'��\/lj���'W�-�J�Z7*�� -��S�W�|{5����e���n�4G϶:�#�����YT��iY�S���sowK{���̟CE����c�\�q�9�m�ž�k5��xQ�F�I����}0֩���&Z�dP��]�@��i�#g�+�<ЦU��U��D�]�  |ЧM�Ie�G�(�/BcE\���V{E'���[s����~�A��ₚ!�f;5ڌ��F_%S	g�wt�JqZ����v�|��m�s;�l��F0>+�M�H|�"��ڥQ�H=�I�w�D�
�>!}Z#��*�U��~o��մ����(��k�B-��0k�Yۖ�}��4L`�4x,\0��1���x� �M�$C1�w	�Y�.7�i}ezj���H1J��ѩST��K2��pc�w�Vݒ��2��f�l�F����V���ʂ����Mq�mL����3[��w��}�k�{��s�}�KX������u�Λz�v�u]V{���>�0���)��j�Q��!4��Xg.B����.c-���.����'f�4A����Z)�i�ġ:ʅ.���vnj=������dƤ��LV���Vk�{"G��v��*Yd�X,�Ol��T����31Fj��A�4ߊԻ��o�C�PD��ܥ�-Q�y��5*{����2;H@]��ŕcK$R��\�U�����/�f���MB���f�%��q���Ī��f�
5:Պ���8g���W��mg�	�	4X�`��N�_��}�<�i�S�9�(DZ?=�\�O�X0���L�Gƕe�3<0���H	MS1��Ƕ�.�*M��l�_�����{Ĝ�Gّ8k^���'_$�7�}����7񂏀��R�Df�PQf���Z��~� o�nH.�mxT��ˁ�t�Y���;/�'c����
�g�pr�\v&Aв��or�\�%����e�Z���z�fU����i������$c(k��`�7T���0�:7&K���i�{��U�C=l@w:��;"vwMP������^��:svNH��n�m��o|�m�,�`�m�����Tm����<��9�r�	��oDg����Q�7�����닇��۷&�=l��zÞ��e��]vʧ/��z#n�/Or��BL�nR�m��t�������U���/@sv]��u8��e�/���/����n{IE�m�;�j[����SP��r`�����p�}*.sQ����t�<��6�܇e��
KH४��,���lG���ұE����b"w��P$,����b�.��	5����=r�˴�L���`�qo>:fR��n��+.�x�������q�.��|8+�f���J��fE�	N�Ra&��9E5/c���3{���-�R�u���BA���HAB�ˬy�U���&��\4�Z�W��x����HH�`Ӷ(SY��:�ؚ6N�j\���s=�̢d���|��xj�_*["�K���
��{3>���	�È'�=��)}�H�Kd���7k']b���D
�uK�0��[T��"�7�M��lnj���j�r�?Lβ����\T�ES���'.Z��k�R�g�O4uӅ�Y;O^U����k�y���aa�۱���y�y9cN���[�=�����D��]��d5N]����t�љ�T�2��MzȖ4��c��#��75?m��g�Yu��)�ƣ�R�*���Uz~C�'T۩W�~\|�g���v>�oۺ�_H��5�Ѥ��ʖ�w5�kX<^�����]S/��:p]�4�N`�H�Tf�ul5'Lt���.��G��N�tK�~_2�n4�Z��r����l�ǯ{E���N'7�X���g�۫�2��!�]7C��.�*��r���9u%��uu��zQ�No�;�޳�x��N����yh�b�{%�a"���
�}fX����Ϸj�؄q���n=��;��r��Ö�[Q�y����V�'2h��te_��aS��spFAmw��G7x�=u��K����R�҉�p��~�eQ�k�_Mz���m�����ũ;��A��m����(vo˦f�k�j#�79ٵ��e6�t�";d+p�ma���[J�����F�!�\P����~���D��8z��9�`��<��y�쮴\�'a����W!�%N9���2
l}�PUE��`#����yJ
=�B����yP�Ʊ�����l�`,�n1\+
�����5�=��#��֘��y��U�]�}�*��v�O�.�}e2.��`Eϩu4㝟Tv��UzC.9��䜜��,�~u��<�_f�$(U��&�$���K�Q�*���Q���4J�����Ku�*�6��<陇;/]��uS�D�F�A����E�[�٧j��X��{o�Vo͏Du�fn��lq!��e�C��n��>�ڵ[���+����Rn&�S`�z�-�wN�-}_]��`�T�����p��12���۬�F\���̷n��>f1GI���P��Y�)=0�7��-;Εr$6����&�v��Ϫ�5��{m�U�ɑVʘ�%�Gj
��.�V��V���C64���k}l����:�6�˲�H��LS9�)��yܬk9
r7�ܪ�X�yۑ̱��}��f'm���9�@[��g\����U��mfIڧ��1�?��~�~I@W��TJ�q?`^i�+w��}l��r�{��3���w+��͊��(���b�����Ks��ܤ��j�d��6�0W��(�I�o(=�Éa	hׂz�QG*�w(E`�%u�2��� �Q��ǽ[��JpQidj���J��(���={&mb����ъ����2�޹z\�x�88�m�b���t�5�I��~S��)�c�z�&�����@��d�_ &|(�=V������p��ζ��)٦C�5V�]xZ����>���q�)�<�2��f5طy�VO*]q�NZ���z{��������vx@=m=�-ܔ�8^+ͮ����t�r����N�m�-�e��U��>=cU�}�&"���$-R���V�;��B�����!X$�L���mɏ2�L��\c�fV4�a�T��=��jvʱ�Pp�t��ڍeֳ�oǹ�L�)����D� Tl&i�MҪ4qtnaK']�W7���W���H銱ۆ�����u#R�6�]k�j݋}�E�����7{Ǽz�BOC�#��"�]�
vu���9�5��S��qϸS�J�Ք7���;�4|����<�+�-6g�Ʃ�B��蹚���W���t�k
B��̙�-xALS6k��Ѐ�?!�Q�9dm]h��ݽB�w��M�Wĺ�wC�e���[�wV��{���N�!P0�[��2��ٹ<F��ѻ�,��2@>{z�#���Z�JЙ��6�Z���e��8jL�5߼~�r-w��e�&�y�[�F��r�_W�����Χ%�o^���ۓ4~I,�C2'C]@�,&ä�L�����_!C6h�*�!w�KQy�+p#�2��b�H|E]-��K��:�y��ذ��V*��Er&�M{W�f������~�*�n�lJ@�,6{8�ٵX�����۶�֘�#*τm�4f`Vt�za�Þ���y�$�U��VI�.�U�<mw��?2�b1�n�������u��y<n�h��a;j��Ѷ����u��m���:�t͌�v�Y��h�'Uug�G��q�-��Sa˂��8-�;7c�gZ_]����<M�g;��[>���M��u���Yz��EI#��r���x��)�Cn=h �ݛ5�n���u����u�N	����	F1W�ػt�r�V���!��<ia�^݃��ļu��!���{Q;��7fgf��NP�� &iC��b�[a��������b�)���䱘,}�"���3�>�R�xH�W����ڢ+��oʷ�����t��>@xWC�D:L�(��m�VB�F�og�-��`�+�?L����7�
�`̡�Ե��=���7�͏,�8X׹�HYT���pǜ��nV+UJ6��=嚮�[!z-&�N�Z����L��n_�������,f�7#d�N�Z�����h�U�k���6H������Ϊ�Ϧx{�Ru7���8,���6j���t��l@E ��U���S�8+��A�R���ٛ�I��!�4M����O��ޡ5l@&q�\ҫ��m��db�� �|��r\���V�Jت�f�{^27����K�8)ݔ$����{�%s�����(��� �/C:�����1�ǲX��Eiwjٝ�9�沫H�  P��>�%�O��z��E��t/�J��N[��9R�ic|�.'f��d33�n��T2ۈ�9���Q;Hsi�!��mK�Fۤ�������y�)!���Xp^��o����;��@(����,p9[i�śX�����I�[���0(EK��Q[c6���`w�mh��7����.�N�ڭR$h=��_�W��AP}6{��^m��czo����K%�뉙�����

b��q�	u}��޲ s�AL��j���R�;g0�C����3�Rp�g��9uPK���t�aʅ.sc��2t��Qi|�$�%])�	}�\�nH�6kEL��72�/�|.��?�bs�|��Ɓ����`ٵ\�a�>��YTo���u�1*��:-$��M�
�#�ȩ�ۘ-^�n�3���jn�PJ˓�OE�==�&N}�|�b٦)�#�]�؀�b�E��59���_,�e���U	ұ��c��g� \����\p]s'c��n8����lZR��⨲hV���1����?M(7F�S�X�ۦ����~V��� ������FX��D�^ �+h���%�ny\����L��`~�s0�ǋY�͊�^��2�$�=�[+n��v'+� +-��ӭ��I���.s7���cΚS82[�o[�&9UTM1�2�����[h}h�_G2����)��J�*�2�����E%�ʒ�]eS�ˤ�a�ձ��gw]��fw�,����2���Ԓ���Xק�}���/#�d�7�V�d��!p�7������RX�$��]��UL}���?U�M�2V6B��=G��>�nn��gy̮<ے�$�*gv�P�| }�5�_I��84bGO���l͉��̱k�z�][�k�@�2��ՔM!
9l�V�-�z��H�c��M���[z�s��۲Cs��v�5�K>z$���cQ���ɶ���c�YR�^��1n�j[^��XE"HR�6�͠��,+���G"o+l"W%�4��Ky�@�6Ԛ�s��&Qm���{a��)/�S=����w������&b��iϥ����?|���~��Gp���.E�	$���e%�z=Y�F�����U����c���������L�ľְ_yWS�+4�6�t��g�a�0���qJ�j�� �C ��'A&���?c���%,���F���Z�k&l��b����>@ֵ~��*����׼ѵb� |�ga���*�	-r�o�R{���<�U	�Hw`�և��F�C���ֶ	4��9Q�q�X�゠��E��oc+����l��:�U�D�o#�)��z�f͂W�Ë��:�f�d'��r�o
{��H���.����?I*���i���8���e���<ك.�q���	����Hwa���}�ξ�1Zc�u�HP��v��ý)���*a�����W�2�m��� #佭>ۖ%^5^�ͣ������qV1�H�z&����w;�T�q�v�iݰ.��j6�y�S��H릨��w'O]�R{���<�����u��T�œDX�V�k�t2��W_X�������cr�����B'���d�N�1�K��j�SD4z߽��w��¥�j3܂�R�*��ƪ���O������]>o��a1I����]��A}�S�C�Ib�i )[��{:Z����J�v�g�o�W���w+��0���}�j��AHd}��<羝+´g��((��qz�JG-P�J���A�k�>^mX��(��	�:^�z2
v�y�z����IL��&�^w�k%�҈c����܏A���O�Ѕ+����:ꋮEUD�7��}��{^䞚��~�5�#����MW���Xt5��F�VEK�a�CV�R��#߹<�H>��5}2F�g��o�����_���^-G@����nC�S�-y�L�۽����0��\[bơ6_q�&t�$�@�Wr�[j٥a�6k����5ӛ�f<���A�
�y&%kz���rȳX��L���^'S5M����ѵ����7{oT�n�!�2H���ܸj��h������ʦ�����1�,S��6��ٲv'�����r�d3���o���:���5y�.�{(q�Cr��"�Oyw�j�v�F���M��eeZ/�Ε�e�Ř:^�&���z_fm����ɷe����[�;�f���1�L�yg/���]�,rlVpn����������?}.�`�۸c��(6����|j�|�C�'Rn���,nW���,Y�iߐ�+ѫ` �I�*{l̺B��R�zp,T�j�+�w+	0(�ūU���n�:��N2�̩��^������+���ҕ�޶R�;:A�̤��ek���W�z9����졈p�ae�3@�� LS"&Z؂SuV����݃����o7�F�[Mf���f��:�qp�nO�(�k�+��L��/�d�5�R*�ՕI̺/:���woy�8:}v�6^��)�*���	�땷3������G&�qZv��ם5�G���@h*)�ђ�p�%��0�/!ͨV,�-Z���v��t�o�CB[|YiU�1S�qi��I�p�l�_F�Щ|ؕ��Kv6Ԫ�;1�Y�SUx&��`5�gʪR���oB����:k%_-,�t��]+٩�b�d�y~�w!�`�7<9�[��-�&�Mm+1�{u��y�\������m�s���Oq�ی�����z����&G�EՎU���[���<�۷vũ�Ϲ��xZ8��y��]������ov2���a���v�ur�����E�t�u:漥z:*x�!����5[��[�Sk[;���';&*[�m�uۍ���\\tdK���ӸL�[�On�waG�4t��1p���tD�1�
�:�ڑ�u�C��w�+Ig� j�9.�k�R7]F�3�`γ�m���m�6�^:�L\L;���4i!6z���W[/K�-��֜Fy{=c�����u��m�ϲ-n9z�ma�K��:�lWk���ȂvL\�G�7����m!ط>9���K�6I�C��6��rut��>�F7���n�Ku�ݭ�Զ��Í�nF���s��ͷ4�s��狗;�+�������Ǧ��Q��۹9S�v�]{k����FgLh�k���׳�&)s�K]�6����{hb��qoB��n�C����n�[��m�n�-��$�z�z��E�h�.���.v��<c.V�!���0b.{��}K�&�3�l�Н���dEg�s�u&ɰ�=�nx�V�5�m�)�sΐ\b�{�Ύ�9b�,x�����b�q���s��mfS��;N���ve��A�p9M&8=D�z��w��SSL�=DP-�o-�89�:|�m���v� ln(�cs��k���]E����i����m�3�upۋ;#7���k{jn=�ՠ�<p���뛅�v5O7c�m/H�Ɨ�x���p[�����x���뵱��nn����[�L.�����s�D	�Ój�i��)����6:5�5�w]f�Ԉ�/:y8q���yN��κz��nt�.��9���úMΘ.�^\���p��\Z�x��y� �Ϫ��j�;={x��Yle��q��sӁ�m�=Nv��;\Gd�)����Lv�=��'b玎�tV�X�����$L���a䞹�Wm�7mOJ Z,���S�"�u�S�D�+b��gsy3���S��f��j��������s�L�b��x�(6⎃[%l��9c���c�us�q�{s2�k����m��"���@R�;>�@u�n�КKs��n�lׂ��S1�h3Ͷ4�gdyt<���'e �6�|a���J F���wm��v�;<���me��*�.��e}[v0�	��\�H�ct�����OF���SvZ+H\��Z����}���ۙ�`��u��7�Θ��ժ�y�x|A�9S؟%(|v%�[�f���1ڃk�f��v�Q�f\����s%|�{�~T���Q��v��,IX9{�q4�
�S ��0�u[��{�AR�j�
�����aV�^F,����`�Y�gN�83����D �`�
L��m)�C,����/��`��|�k8����Σ��4U�M�.�언}�ɭUl�W(�[.��O0�&�mڗQs��ה��m�	�zܶ�y>��e�/|%xQ��T���������%��O����7S*�u���e�6]"�t�J�J82���&53��M�F���j�a�����Co&�����eF���y5�����W�b�0�v3�;6��I��l��T�T`���ظ�����ݦ�u�AwdL��s�']�.nzJ�)$L��}�����M!�O�xk��AA�#��s����c��ѩw��2ӥ�Y�H������n�;���K.�)�J��i�Xi�Py&ꐡ�n�;o�R\h��}a�����a��^&�"Z�WE��C�uo]ƨmH��LT��o���X��$13:{����B���,�j�c���W�c��Eh�Kf��X�c�=�}�0{y�cB��W"|XI+v�Yg f�����G� W��x|md�'�d)Uש��*���Fa����bݍ�EZ)�*��E(Z�aL�A�5Yۡ�͜�Y}Ƕ��j��B��<��H����&�79�7��ˬ�Xc�7uf�� �.�e&�?��Q��Pc�����굲���Y�Ɋ�*�w�6�/j!`�q]�]�}�<�4��r�L?(�l}{|��H���`^�J���+��Q6���[���p�ۣZۋ��H\��i͹;m���ɣi{s\�f2j�?_ߌ�����{���;�E����,B�k��+UƏ�C��>س�v5�Nf�q:�:��A�E!Qfv�_���3�}��L��ܺ�C郺��2+�l����j��S��*�x��L]���j��5��{r���T�k-��m�m�����W����ET'�Y/��'�P��H�{��V�����}��Ǐخv�J�`�͜I�9�V&e�ջP���]qyV��(*ש~>�Xf���).�Jт�nˏuG��c������݊�397�傖��	3+�ZT��3�K�ﴙ��o��ۜb8� »��]�^��\~�â����9��p[_1����n�d�mqЕ-�܎��F�^콕��HV�+�8���֎D�m�d�yҐ��,��w�5^[jܤfW��t�n�'�I�n��7�Y��hlcqp�y���i�Hp�5��a#qsʰ˝ۜ:��Ɩ[� t�U�nB�����n f�l�v�TQ>kt�b))���O�n�{֯�l�Y��S�n�F�;�j��� �۠)��rs���I��g��~<�-+v&a]V|�+���^�ܢ>KrN���V��i&ei��*����4kM*tS!�p��;x++����������OOo�k|29�!�/{���zq ��xZyy9ͣHQ4V>�V���U��(�F�'I6I�CM2��[�c��wurul���=m�̠}˙�l1X�f�}<{�W����R�Gpd���M�-b� �^�,^�� 21��|�3�Ogov�8�+�Vf���ժ������t`bv����6��P�;���&ׇ,kms7����hT��e.v.��]�Z���]ߥ�vJ��[�r_,���>S#�E�*a���ʊ������h]�b^z�
�[�x�ٰ[NO)F�3q�筻�pr��.�m������mA5%j�te
� ��ɽ�NLG�x�&<E���]�U��4���.�����{�xEW�������Bk�CQw�s��Tʤ� g>+fWÁDݭ�5I�d�ڵ�{�o�b�#|��"��9F��� 2��mN�î�X�����U�U;'�t���#��(�$���N|���w<�}7�����s��f:sӐ��Ȳe�U?b�s<gx���*y�����J�Y斮�\`#��6�&�;ᆯ�����x�8��t�T�j��V��g(//�.���=������R��Nv�N�qzD����W�sВ��AY(3Ҙ�kR4�ܚ.�[O�Cf��۴=Kk�&��h��A��W���Y	7���`-*6)W{�{�5h<��;y7 �gϙ
���:�m��[�s�.����E���؞��o/w{����*�0���_&���b�����o��՜���Cu,�U[��(�91Ҋgj:l�͑"��۱ҵ�:�M9�Qۮ�N�.�)�ݭ�n��϶��=����)ˎr���t�{v�L��Y�t�V�en�ۓ��Xڹ;T)UR&�v:�M9k��Ki�8�땧��Fp�UŞc����Jx��DG'&���u�NK��ո��GV�Z.���wF޸�t��g;����i�V��f�Q̄��yۮ.Ժ-����nu�����z�����}���J�UULD�ӂ(uU>��~r�+���o��0���LH>�o��7�#��T��ks*}�(������4c�&�*=��O@-+d
�%�F�Z�罕-a�fƝ�_�s�2�H����}��xpx3	8���zza�|VM��W�Vn^Zڱ 4HZ�D���l���E�U�WQB�AA�/%jo���X�Ej����U�,?L�ԁ�޾?g�[~>����X�h�'�;��Xt� t��An�
7m/j|I����}���w(�k��5k��ȴx�U����f��*fjF���y��R�ܻmV;X�UU����R�.H���U��)��T#<��8�l��_���3�_6i
:�N�8���(�4y;��J�{.��v=<��:��2Om�$�����؀�9d���tֱG��މ�8��y�]�R��䲸Ӟ���q�w�҃��4�R���\I�R��g�z̐߆���m�p��m<�͉b�=ř���.2�Z roZ̀��L>��Y��&b ���ڍ�gs�k����s�ΞփOx�6�k��]iM�������`�z	�*R;&nN�-,(��)6<�⿃lh��߭��`4��UX�Kͱ�m��<�R���bZ.�GP�����9f'4��i��� �)��,}���FA�Ňo�π��|nxO��t�6z�=X�y�s�]M�WaE�u�s��O^Dn�W���2��J�H1��6��K�x̸��_����X�����1'/g����ڸ��t�r�BK�mS��
ٻ�=u��(TTV����\��C��3�.}�U��_H����p��Y�r�-ۏu)�um�n�� 쌺6+$�8{N�r3^,�ܩ0]�['+q���Fu�����x�=��&u{�Ee�j�ٲzc����*U�>��Xi��:��E�{��(.��rU��k�	*w��E�@��re�]I�S�4�����
�-�q�P�i��OCm^̥Q���=Nl�h�g+ lդ>6X���&�-�[���c=�~�������
�RX6#d�3�]�����
�w�+Έ�q��Q��Й�<����X3dj9��WS��r��n��}3s����s^��Y;:[Z��x���k.0X7�hХn���.��J'�.8u6�t[��m6�+F&9�j��r�B�Ж�����vRE:��ŋiQ�8e�;Tؾxw�8}ԇh3��4�V5���{��6��`:И��9ɭ��Rxr�;d�w�����`��o����y�}�������b����Jq���ۧ��̘r���B!�D:!sv���Nm��N��\�}k9�m�jܛ�Ӎ��!��܁p#i�Azk�����Y��H�s�z�6�V�^��.��m�2�����lY}[�5��_w�^����c��}X�]�U���yf#Q^����:���n�������^�RH{��|��n��ˤ�v��E!��� %��Tgt����<e��*�4l��3R﹮Y�KN�{nJ�Vb+o�hV��ۭ���Dؗ��Q|�ܐҗ�Q;tUre��(&Lo�YW}7]��cv/��z���rm�S�|�O��>�^n�>����Tx8+m���7v�{lg�Ҋ堃�q��>zX���<2[yn#�=�[Y�`��`�X�ou�]n+5]��8)�5sr���Yem<��[��EQT@9�m��3;��WD�ɠx��Pڋ������<1�t;�	J�T�!�zU��r�B���2m����DU�\���F�_nvoW�t�g�>�n�l;Ó�8���T��k� �j�	[���9G�e�7���n��m�������b{ڪMB>��1u2���ou�K�+��SF��rIE�I���l��j��P�h���9z��1`5�%)P|ߊ����C�z�X}�7 ��A�C���� X�-�I��q'��{����ν��`���6|^�:Ͱj�̺ޞ/�[�.��őYh�)�t�H��ͫ���]~�7]�\��y9�����J�+��J�!���]�;xީ��v��KW x*����[']�nP��MHQ��\�ro=/
��w�V�0J�
|����povf׷#�bCPwL�3O7wm�q���)�U7E���2��y�e ��e��;��ܰsN���&����6�%=��hVT�һ{J�d
^vm9r�J%�ܶ���rr�{�}>�#�)�r"��]Q���qy841q��Y��(�_d��;�zyä�^�of۶j�����Iǳ�<�{w�c+��hL����o��5fێޘ�-XoWWk2-D����\s&�F�6����	�i�C�)���ʥlI��og.�y]Ѫ2�v�ԁc��<�'k�7'lu�V���I��݇G�>l�n�Iڳ���:;����ٰ�{)��z.���]��Lv�Y:lO7fK�>�cawAR�\��dj7(���5�d�s�n������w~YJ���a��)X�%��'�ͱ���=t�)���C~;`Z���[A!Œh�E��/O�U��nפ�����]V�97fh��P>q�tN��J�a	Y��P^�5�E\non�j�P)��#'XD�eBm��.}zie�'����7�Jqpwe����Ƹ�S<pX�m蹙M(����q���Lp��<@��T���3>��'<���x�n��
��~Y�:�7=�0�J"^��b��W7JUr���Q����Ye������L6�:�[
�&Xo�6_q���zj�n�^r�LͿ�@�C<͵JW�0�[-�R�q��E�V27薫񫵐a�;~{��i����㛰�i 6�Xy9���F�NԼ^��0�e�0˲c��]9;4��Ѫo�%���*�S�P|���\�V:��~4!�pN��l�jw��½�z;��Ss��G��5�j2�+(&��4t^U'���&,�������\�F���֥��bQ�׻��ϖ���y�v��`�C���ȼY�׈|�Y�����=��`�`S�}��h�z�����8i+��p�vs�s�n�ʹb�M/&�|�|�̵I��X�-a�Bd�͔���X�}oO�����x1yk���=Y���8��jp�$��2_�����l��^g�'-���S̫� ����x�f&��ɚ��u�&�{�%h�Ɠ	k͉F/�^z9_Cw�A]s��VM������yL�F�(��S� � $�0�I�W��
v&�ym��4��j�S�l�M��a C��݉ܠ���NSp�z�僝N�m������Uj�n*)Z-���D9�s��{kc46�ݫW]h`h�yf���)��b��.*n��w�n�)���*��Iv�\׾d�4���z����V)���
l	�ɵ�2��
�T�4�%��~X�	���
�mb(s��V�x������&���k��t�,��ɝ/�ϳ��=��mauc�幅Ĩ2�i�T�����s$42>�8L�n���W�'˵�N���v����xϦ'�kk��QfĞF�u�q�#�룽�E�ǻ�,n�N"�ZMtǊ\1���!#���;,�����n[��o'w�{�H��x�ܹ��,WX��;oBϛ�wC[�?�}�v)�[�E-kQ^z܂�L״�=w" �8��-ݷh`��3e�pBMْ�(�~ �gƼ�-�G٢�ԞMw)V�m��cЖ�W���6�hYՏO�&z��w'��N��U�u��o]u����_9/���"��e��1K�1�p\VU��x�c��
�.٨T�3e�b�,�M�@��c�?{�Jo]{�������"JBRX���@ӎ���ujG�
{���u����W�f��u1�^MiiZ�s����3J}jOبL
C*i�u��4�~�C�����!���gn��;��[�WSq��ve���+1�[4i�B�n>x�����̀��n���r
d�1�|�q����6�����k��+��n�.�y�Ӓ�M�� �*<�hT���wc��Ш����f�(_E�X����3��6-t��\�VH�c�vs�/礮��v�������;o*�[0�6�u�~��8I���t�����$:���w�;�B��v�8_V��J#cR_)�{�#3�T�2}ۊ�ԇY��WfM�ݻÅ�ʩͳt���e#Tg7���t���K��mJY���q���>�Kڔ�2�\��b�Cx��/�]�{O6c8v���Fn��l�_n|�!#4t�*u7�*~�c/l!XB�>�WH�WG2�4�I�ٕm*[���7�	/�t�m���z��\�H,i5�f�@�YVP��W�kt�7����!���_������$��b��i�ޝ��g[�s����82oF�\��u�YKYXE������Mǩ��ϱ������&��o�z}����w{��(֜,t�n7<��݌s�A�Wv9�>nvR<U��׹��ܷ�mc�Ce3��VHe�ǜ>���n�6;�SïqE�{�mz��<�M�y��Eh���Q�z�۩M"� a��$�d�i�k�t�Nw�8g��;:��Ԑ�ԻϱX/��Yn����4N���D����VX7y��y��,�1�G[�|xCQQ+���'���M�	�sb�Tj�y�쫣�� ��:�̨Wn<�)T��HE�[�|��4<�����r��W̒��@�,��ax�hD�8��]�N������^Y����e���F3b��{��:u��ұ;k=
�nQp-���$1]�@V$��¡��B�[��ۡ�ɞŨ�Ύ�M۠*!�+�q����#*V��y��>L>b���M��4 �o7����X���{"G5þ�vo���y��x���|7��At���_�:�e���2�8G���-���Ϣ�w���ԭ��_i�K��=��w3x�wD���%�G`gƨG�W!dR�-�_X�V���������M��:�ja/`�^>Gُ��n\w��D�B!���n�>iڵ4���k�{����q�$b�T" p#�>�ۦ�b�od��p~���m�↿e�բnRRTtS��9�����v���D`���<yz�PsuyF��2h5H�D �u؏�v��3��ɴ�Pޕ��B���i �a�ٷk�ܟ���ʳ�\��}X�)�B	�D*m7���2r����(x���ҵu�%���5���䩝yuf�6ɡBe�{\6�]z�]��m_�K�v��R�R
� NrmL��˷8d>���c�{���a>x;��B�����k{����$�3����U��~��+��e>�W��߭�:��٦֍���d�ND�hDl�3��\�6���QO ��&)�V�]W��_vf�)��X��o2Ɖ�6v}uϨ >t~1�P�[iS�󬻲�v�nzq�e�^�^�s�e��1�ܞ��pRtqV�I%�J�����y!����9��T��=����8`|1��=i�6���s��m�ln>#��5N��8�a2}�w�Qqh���;Kط.�kl����']�˷6��v+�y�fs�<�up��ފ?ӷ���@6�ּ��mq�%PlS�����m� �\D|�r�lxι\��̭��4f��W��VVfa�����b��А�9*&D^���Qܞ����oه�Q�,8���׫+�NZ,��rK$�I��N��p>�����8���\w�R�%=yd��-��^�U��5^�2�Hi�+7&��Z��$���m���^y�nI��l�4��������\0�q��Ir�X��~B�";���iӧ츝F�� #@&�(�E��Vn�/ ���n��V^ڧX|ڽ�����ғS�?g�ݔ]�ׁf�ۧ���\{��浛V/�p�� �h K�ӯ`�i�;"�}�U�8&�ڟ'\�Ao|����ES�W���������Qyd��\6�%�/�+����K`Hz�9�U`�R�lnю�ٹ�nR㛳&O���w�I�-����U�Ǝ��K������hw���4I�p��L��ޤ���V��ݹ�h��3/.b��:�y�}��FGP�#��[G-r��S}i[��{�fTEj>;Ej�<y��"܃;x�C�����)��}���W��bc�w�t�g.!>6���v	� �!Sg�a�.�v�.�wYG�Y)`L��c��i��*���Ft
�E\~^9�RK\��Y�i����,q��iI���	8q�[S W��|����)�a�_�<��kC[��c^{��R>*_��xf.��v�*�M:,�M&L����{�q�fwz�]
!��)����@�����ll£z�ЫM�M�\{H:hd�d���LpD�t�q%-���9��r:H��u�����%��/�C��;�y��7ђ4�$�8댤�ƥY7}��Z�ڧe��guI�"'�v�J�[rЁM��ÇBp�����eᰅ�Tj0[����N쳎g��h���3vn1%�b���u��cO׽��V`�YB�\ݕ��9�?g�2��a��n�M���0�Qt� ��d4±t�b�4�'����Yb�)޽ޤ��¥b��ʝ�`k���e��pM8g_���~R���I"i&CE�%���2u�WJ�{%���[��#���i��� ������W�ag]Na"sm*�6��԰�7
R��h�F�+��m��w7���ɚ�Q��R�.J����/�'xV�<��9'����;�i���*��Em$PpMd��rg>mrN.�ҕ�_mu��1�mݑ�>w]۹������^�Ip�~���=����r/�3Ԩ�
ԁ`����)Z��)�r#�v��/.x�6v��1K�җ�͂Ҕ���85d�Z��>�_{��Nm�[%@�+@;(uvr�5`u��Oc�Ry��թ�����,� �L���!]��ޕ�����0|d0,?�J5��B���w�gڸT��bʗ�|h�<;n^7s�����T�,:D�q�Ϡ�ͨNÏ(W{�T�V��>����Kg�{K��=5��$����&����V}A�VrmN��N�� �yo9��L�^�)�}W�b�o�悈:!�D%.��׃^̕���P����i-^��4���m3��i���< �g�?lםJ���	ՈH�_�{��L}��y�[�̶ϯ���}�X:��(�u�K"y;�I�qy��~kH{M�W�����9W��cɍ���B�l;��-d��ꨶL(/f�^�K���5��edI��}�%J�(��@tt���%D�����n�`�;��><�.ϰ�CkN��-�5e�\�tl�ve��P����-���;�U��R�˵���8v�`�}���2l=:������;�f�e;	���\���CG����Vgl�U+�r�2�[.�o���@�Ĵ�d�4�Y�<jxqᖦ����Xc-��n�'���d�$V4����Wǁ&?w7W���@A��권K��_;�^�މ����b��v����X��O�M�[������u"�E�KuhfL�rӜ|P��2�Y��i��٣�>�~�G����VRA�/��<��h��:,*($�X���c��n��qs�Օ���F��]$��On1�^G��8�lr;��yO6��SCN�9��t�tۤPI��p7-?W��f�Ė���f��)<�h\*������5�g�&��VXB�����,ggiN��@�x��#���w<��Kuu�������]���}��)_H�r})J޻(_ ���C����⮢�m�)v$ɓc���c���@o" [�d�^��R���J�x��B,N`��J޲	V��uk��k;\���%���61.�z�͋�whNz����� �=)͎M��Z�ω뜇E�1����Z�#�����ܧ��W*�]au����j�u��<��@�y�(U��6s�퍰x��q�����B�
x��ɺ)��^�z��	]m��N��רwmϒw7lt���(ǭЛTc����m\�gv���}���6*9ָ���]���X�N��۷���J��y�wnJ�7��k�����S��w�w��S�;��}~�T�����L9hK8v+�6�g��s�̦�&*���J�%�]2
��-�ٯ�!ñJ�Q:�^��j>�w��_����=E^n�]���z�f���c��f��H�����3<��B�UX�h�q�0�Mq���^�E/�cE��R�<�ѭ�Z���L���H�/����~f�O��R�b�2K@�mA
R*����6:��}�]�''q���\x�Vy����e=~޵��|��z�J����^m�w5cRJ�	Ae���=��zr~	5�_S���#��ڦ{��s14�W���3��m�_K6�{"x�݇ް��6�4Za���ζ�k���:��\��n^���\:���>u&��)��)$C
�L_~���m5��om��;&���uA{&q�t%ں=�aUY.�4d/�\M���e�Fֳ�K׈�	��0q&)6w�ز|�������6h��B�F(t0�ei�kq���u��%��WRPOe];yI���*e�b�˚�۹(#�Q*�].H���ڜ��us�����|3���;ޣ��&��o�L��x5�G�L�`gRӎ��{r�32�9geC`��{�1��$Ȧx��Hy�5s�������J�;s��f=��Gcn����+��mz|�R�Ҵ�y�XȻ6JchX�J;�����2M��U����X<��E��(�S6�B3��ȧj�f?PO��{�^ ���"e��[.��t�.'�ݧm]�Ժ1�};���v���Wj����{|�X���6�mV0T��v�M|բ��u��L�$Hnܬ�2���E����k����*TP�f����������3de�w	'�����;3�L�G�b��-�H���I��{ҶY����ڱG�P��c�(E ��o�z������1�Q��b�K���C��X��_iP���}�s��)����7̩�wp�RHy�����
PS.���I:㊕鼷~|�yZ�a�c��sY�+��,��o+Jy*�Yì#n�CG���чeιCzw<]��.�vL\�O���>�rmZ��{�;i�Ӵ��k���K���������%
t� ���Èz�f8�{e��Z5�Z-��r����9���Jhx����N�i�j�J����إ�A]��� �v�g�������Ub���DvQ�����y��d�4(��v\Z��ѩ"Q!P/��:�����!�3꽪W�ӗ�{��ˣ�ܐU�h9A�M!J�-�㛒z�q7�rt�-vێv!���ۮ:���.���e���-�¢z���Hq�y�8��pDc{Φc�f��w�zy�h���N�V���r����$7A�۫�����U�{���{}�]���~�b,�3@S�Ob��-�]��{����#r�Uozg���fk�%\����j^Wz��&�)�ڤJI��;�]��~�H#�7�
s�����i���کܵTYN��H�`��o��w�-���H��,A!���W�E'۞9���1���k��ۭ��X���]��9��[���>i���C| �u��ǅ*�8E��Ee� ��u혷�:�o&Q��.�z��=�t=�~�kۆl�-<�8wP�d�����q��{@e�������0�Φ��u�=�JZ� ��U�
�|��a&n�(�֟54E�Z�\�������ڮ3;�ix��1'	֛7u�g>����aX��~ݓ�3~��L�sl���v:��Y�Y�s��]�$nv��SQ����웳В��%�z3
�g]�ߗ��9��3iA\+���r��P�ᘶ���$���g{�����[��n��s�>�����3QZ]��7��GP�����jZ[%*6�4P��庎f`QW/<�p�y-��^.���>��\��u�ܹ��D)z
�H")#x6�6+$����6~LQ!�'�ͤZJ��c�̷MSog��1Db<����i0� �&%�jϦu@�o(���,^%A�kK2X��Vs��Ѯȅe��Q����ϣ�楼w�� �����q%РF�~��e/�`���aʌ�u�	١�a�#_�ˎ������z�N��]Y���߳�^����pk�)�j�&��"Gvp����ֶ-ۺV�'@ t�$�2�뼋6�@�є�V�-�����) ����gU�$"���J�U�̫�\��[Y�'�wS2U�[5Z钤zP ����ݵ�=Ȭ�m��y>�b�P��Ӳ��bqN��a͠��O�����U\����
��#b��6��F�ژ��[$��f ���c�i��Yw��)�`��{VjY�j�U�����[�o�`�G�4D��]A��d�0Vk++��]e<�N)f��ή<�`ˇYK��\vBr��]���#���ҏ�Xj6x����7��-�+��ƫ"�k���s��z�1�������q�/I����ϒ��;�k��%!���f��JP1��9�&��z�@�7���.��q.�[0{ip�gvl)3ц�m*e]�-�w��C�Z[h� ��R��n�x��k]U���P��ݼ�� ��g��xrRs|��7J��6����P�\r�|��o@�f�|�L;d��:��=�ee�9�t�E-���YӺX�V���B�!�h�(���dn`�5�nV5�Ynؒ�ˬ*�QZ���ٽ}ʎ�''ԃ|�mZ���ܭ�m{�>���z!r�v�Q��J+�0�7�`1yb�gu�X�����V!��y�Jڭ]�,�v嵵����.�0(�V^��S�i^����h+�\���:�R}��q�gʟWj���X]JD5C�{ӸW+��a�&�,Ɩ5·�-�꟥���������
ʲ���)C����Ut��s��h�W:�p��{s��f�����9x���v���ǍY�g X�s�qǗ��N��Rm�;��m���v�^�'��On[���ۣv��upA�4k'�\;n��F-�D^ɻv��+Gɱ�we�!�6�`��E��M��d۱�8���3���qU��{L����K���;�zx�K=��'�t3�����.�+t�����b8�z�k��x5m�۲�7Y3��O<;ۓ<]p��vf�#���E����r��غ��;F0O ײl�Mڦ�C�����X<��q2z�2�&��s���놮;����'��7���OP(^yh��uƮ��r�c�vl�Mu���=��g�]�vַk���Y�y���cԻ9�uQ9[����s���c�n���yM���y�ʤ��c�cώM�v��Þ��:����n�]��-�c���v�&D�H:�ˣ��h���.L�v���r�l��]��nN�x��,���c�Gm���eA�Z7S%�0�k����_�S��9�@&�C��k��;X�6���u�V-'T��7=T@��&v�N�� �[;[��RB旴&�c���M�.���n;�SV�v: 2�7��a���(��Vܻ׸C�x�x��]HM{�n.��&��'S�+����½t��N�!pm��|�� =�r'k�V���1t���g�����6$-��g��=��v���z�m��<ƞ�G]�xʙuOӱ/YV�M�
��m6��M�ss������1����\��s^hu�ٜ�9��u�WJ�k+�.�9��k.;����v���C�#�<r�849[o�!�M��UZq��9�!}qËn��Wn��-���v�9[hs�T�]I ��r��G.�z���j�A��rlzVu�s�[���η����`6�l�i���׮P�4x�na�<h���u�Õ�-�Ni맱��n�q��GS�0����7#�wcl�]��m�ik����]Ůs=�r����a���kk>f�������U�M��l�n��;sKQ��]K��"ûb�׊���{��9҆���v%��[��:_g,b]��F���^ڀ�GKs��i���v�N�Y����#��*:��:���T-�fx��׮7c��*��ϳm�ςkZ��,ON��v�����(�r]g�s���l��v;tW<�b�3{6��#�N쑎ܕWmgqt�GA�� ��w���fy�s����H��ݜ
�k��oL�!0߼��f�����]����7��A�R�A��AR-�We������^�*դg�h���v��)&�r��m�!"��^i�������݊h�}�/�+��6�ݎ�Ho���4��7noz{��8��~
���J���V�+r���睾��]]�^�c�+M�B�h�ܮ�
 �ʯfw�OL�����P�
��Wbt=�1f&~�-.��m�7�Q��X��V�E  �*Xr�����(�C�;��n�9�e����]X��b��3#��t��SU����n�s�����T��	WF�*��%Y3L:��0FSmp[
��t�c�*s���d^(�hƶ������z�o~����X��q{�>C��,��V����]҆Ïg�*�� �d�u�R�A�d�r����'���M�ɭ����׉�yQbbL��.Sۘ�b�Ku���Ub�5YSp%��m�e kCq��/���� �oa����V���B_T�৷#^�+��{��lf=~�d2��������2��mR�l�]��䱀BN���T`�\��}7;[w��e���'���LV����q_r�I�o�[��i�S嵕c�p%�4�(��l^m�'S�ۗ��<%���L�o�Y��l7��%FMf�������oX�;���#�Ā����͝NIJ��ˍe4��	���'�o�\�_����?�d�ޗ�i��M�����˙�;2���|�Z��=�ـZ>��s�wÈ���w��~��nz�
RZi���\t�DT�=��)�D�L)����d{dR ���&/J�	�_��*<��4�\���׼�,�{�~[NT�}��.>����͊���~v�#T�0�B�B'�TG����MwF�{�s�U�S<���n�������yT;��"��rok�g8ʂ�a�I*tC�H���q���7ػ`��Bt�;���_��Ww z��K�V��L�T��P]����c+�ѯ*�O46h�2j�PyּY�2o�$�o5��Hm뗄�"�a[�Y�\�O��e��	�G<��n��U4Y�(7���w��qI�f��'fc��ߗD�;31�t	$�>�¶��8)�V؊
��]���Ǚ"���'t����H��@�,�n0�^��,�r	�X�Zں:MD7������)�܌L�B�K�����Ջ��A��a��|^}�ETNYc��mYm�h�7Xp�Wc�I u�"i��z켗<�&�%��`&ƺ�\��=�3�a$��/�%�GY��pz{�J9�e{���n�h6�iۺ�-�uXK���i4�i�#�nL�x4�kP���%�'�}�}*x >G�޶�R�gzSn����7nr��E�1�L&PM1���g��fK��L��!\g5*��A1=���Pv*�W⽦�-;xԨ#� �D�vh���Է�ܫS'Z3����l�tb��׃.��p+7���/},� �	�eS3{H��դ����U����0�{7e�B���o]bW{]�X�� ʲӼ(lFUd�[H����roG��ۖ���+�0���
�<f��:���5�=��X;۬��Z;�8��.�.�]	$��ǲ�Ɇ��bх0���\���A$��k��f���Kl,5R��q��{���vܽa�]�k	��vU���ˣ�5��k ����3)��Jo�鼢X{��"x%y��6��c���~����@�m��ޛ�Re�k���^*���WT3(��N]o��+S�43��\�`�z뮷�׃
k��;[G�K�3;=�Ԩ%�*Jaa�Z߈,3AJ�&;3�A�9WYB�b�����g�B̧�Y�\����B=;|�*���.��F���Ku�OQ.�t%�-�8��MBo��b,[ �^,}폳J�^y}�c60N�t�@�\Mm��疮���p+Y7l{Z)7L�h�o����ho���cz{�՘�έ���{jZ��v`¬�(Te�w�t����O�ǧz�y�-��i���dt�[�j�a�r��^�j��{�cbm�YדT��^��U��^�fgh�l��/G�wƅ|�ѢRE��m�+�v��e��_5^��%�;2�]�y6�;����m��-�M���6ܺ�;'ct�^�nd=�vx�/g�����d}�g\�z�
j���-����Ξ7S�:֋-�u���m�I�/3��hNs��g#��j��3G����7[�� �λ7&6��Wov��O�I��	͔jz��z�G�;/1��!�s�6��#����+�`기��yk���p�
���ö�u]@h�7ᬐ^~~\_�[����boV�L�\nwrU�(�]�����ˎJ(׶4�(̆Z^þ���"wY�;p��$Sc [�n�^�g��YB�WO<�&~Y�g,�Y��_c����t|R�~�)of�nq(����}�L%��&�dMZ�8]:�b�g[�<�=�o3�3
�v;{���̈́,�a�����%�����o�yӪ/���X�Q�6����R]���E��:�x������N�4����c��<���v6�玆��]LGmL*e	ˋ;�(�>�g�v}}H�L��!��N��i�R�a�E�◎N������pO�u?�v�
,Y*�H鎕��!�Ghq��oi�x�wl)q�{�6����GGS�մ7}�߿���[��w�v���53�m�Mc�{��w�q.2��"��ן��:��*Q�w2��piQ�i0n���ˢ���]o�G�|G.6�ۆ�(�+�.�v�U�$�ԉSM[��<���օN���R���ˊ��6*�o�w���Y����z�]�z�����k��*�/%������G��m�*�d҂T��i2�SML��t1s�fy>�M�����������n��9��׊C�|�w��j�pߣ�'<����BRZ�/��}uO�;@�qy�^��Vn{r1�~ܚ�E��|���R}x�H��u��6�����A�� &��UEC���k��v�u[�Y�;Qr����%�2��z�z�����{�9�m7�}��̹��,Nd��b����v.��S�:KX���2.�]mf�&��6�z�ӡ��)�����A�� �5�ؿ�_�n�������7��z�����z���{��=2�Jeg�^�U�]���G	���O�>���DY�+�&��>��T�'�}0xj�|ڋݓ(J��Wt�y����7E4ʤ�2�I��TM�آ'x���L+���r�I�l���X�)�9����L���' Kد!SU��xz����7XeGX&��;Uc��h*V���Ge���mcƁ���~�	�ez�ZZ����TT N�x��M�9uz�+/�̽� 's��.�	uM���a=��^��s���`�:�d�Q���^���D!+
<^ow ׾�sv�@t��7�{�߇gJ{�Jp��ڬ���X�,��'	?��p�w���w��$4�@�F�lNB"��.��f^������Zx�u;�F��	��@�6���ג����/$�_���롺�K��(��=_M��E����g���β�����!�����<X76�z�<o{���V�q�$��{,{�"y�v9��ݵ��z�-����Ñ�=xf߁M7I���a���\|�xJr��bO��MAMV�X3*�x��?K:��:#K�� ��2�*ܩ�Z5�����s�r�m\ݽ9e��:�/S|��V�X>�L���e�V}z���؅��+�#�Q릗�(Y�T��E�>x#w���f�N����⬛�q��Q Ђ�����b���T����/1+4�h��%�T&vz�ӈ��2"%x|�OL>�w �Q��ln�fP�{�	.������7�ނ+r���2�6i�'R.�����᭳'3�h�����:�!q:S�������nNZ����b({}����f`�<���J��^��I��[�8��*��|�	�!��}O}ɲ�:.�n�l���^۞���b�?"{�+��Aڬ�L�P�U�� ��5l��z�z��ぉ<�c�'���IY	�]4�-��Y1�7C��}|��ӛCi�~b�Cw�<�m��Y�H�O�۰�yt�X���]�ϕ4�i7�e�}�pt�<��;u���d��L��u=Ǫ�/����Sz[(�p�;L�(�<�`�D��@�M�A4�'@��lr��:}�t>�ʉ5��+VNk�+7�7|m�����y��p�N�y����J�Y��'���a,����t�AR������������x3��Q��p\�m4�gi�D�nν=�H`k7����4DZ��'��C�x0.��,փ�٫���@���ܭu�'6f�r���J�ӎ�ۍv�0e�ۇ�si-�y�g���M[��h��{n�<
 UĽ)�r�3�q]���n�[p���8�a۩hCky�����';:��z�չzy����v�06CZ'U]�ݝ�Ж]x��N�/k�]��䮣5�+����Z�!����ޚ��a��V����<:�8ss���t'׭�����[V�{u��`�{���T���04[^��G/b~�$�u���B�	N�á�^]E�ϲ}�vJʉ��ɖ�A�$
=�-/IwΈ��{5j�r�V�~}�aܝ1y�_�ݒ��9�f�e�&��{��;�:2�.��K-����"{���k'��QՔ>��5ˑʿL�t�ڙA�o�����[��b�5�a�[Baư�.��Sr��%�z�&�,3`\�s�}q�;Y�^tھhμ�46�<�y9:�{i`t���RN���o)1n�+u�o�Y��a3ހ��W뗟B����!�3��lD}���?���<����,M4�m��U���5N���ó�{t��4b2�Y�>^+iRL�Z`�����:$Kṝ-ǡ��d�Y�C]���z�x�*����od�;&kצB� ��a�(R)�Vz5�z������3��p��5 �K��U�u���z�4�+{�~��wz��_ h��P[�w%�ܰ�V��8�}���V_
;��U��U�~}�s�{�4L�����V>ڼ�&�cOI�RNĩm�w����#=��ԋ�QH6ڥ@���&��0����h�^�Qn\�YʼtU����+���d�J�y��H9�\���(��)��@�e��t���_�9VI~������!\q��Wm�T��7��~�"	ߋb�E�oo��{�<��Z�Yߑ���u4M��\��k�o/ǳ��Ty��-��l?oVL�B�"I��T���w{ʀ&v�}6
VG��}=�ͫ�xy^���N	�l�ltjn{{4ۓ>�zl71�\�����r��*�����8`%A�=���G�J���C���}��=����GK���.�j\�}�V�/����JŠ�9�s�@�Ӣ(I�]X��.�]�����3{�\{��۱��0:�t���V�0\�v�rw��Ǣ�Cf�(���M�I�#�h�W�,�������R�]�P��W/j�$�����*w35S���8��{v�mX�h��v_3�\:�B��Xf|1[�A�=V�oh��EvWf�2���G�MU��"wQ�P�wOgc��]ksMi�9��M�����_�ۚab�����v��Cx�h�"I���dp��T�5��2��V���y��MӞM�M�;DН/A�y��GcO#N�٬ʼس+i��%\]��O|��v/+}chxG�wl�]�$Q�Y�Z��4��"Y~�f�4<��o�h���R��r$̉뷾t�� ����r^�#��J >�F~%�~d�w�玕9w�{��\I��W�D���C��E�)�0K�9^�a��}�'����4�u�+z��2p�b��>ՀT(��WR�B�[H���.��;i��rve��x�1��.�����*�;֩ĠS�x���Pþ�����]�s��+0g	b]�"�z"��>�Y8#���Q��ߛƚ�{���E`2hԎs1t�R�La�Ȗm���݆����� Ij���:n�ӳhR��iWD�r睙����UY���g	s}��f�ۛ����K���ǩ2��:�:	Y�E%�Q7M��+����+�H�����Q6���w{r�9�N�{����e����K#ܺ��V�0M�%�yb��v�ʨ�N�<,e)��8֠��������y�𤐙0�}����d͆u�]ϻ�F*b�����YK��G8q���F���M�6���fK�X�A��U�jM[���wKi�/iRL"V=�Ը����őr��Ąl�#Q�	S�Bm$�_���V��9�aY0�z9�l�>���8^�nY�F�e;.0Zubf�خY=��H�Hz�S�FR���M�٣ޛOٚ����gkW����{_u�x�ϷJ�7F;�of�ʘI�7&�җ��a�+]�<i�MR�X1�8��j��g������c<�ڵ�{���1�]���96��B�2��ӏ����L��*�}X�W���vs2����C��h?j���Ϊ0�;h�/=��>�R1�?���=�_Gb'�%�T9�sL��-��>>���#]��S�[vO��\ڦu��>����ڭ��y�h�o#��W���r��E:g{s�l�cF}��Xy�\e7�v�s����W�������8����G���z�O�����#�4RکK�.��̧mcƲ��󖟾��F#Y楢&2�̭�X�>����CUW���z{P�t������K���Ʊ�= ��Ƈ���a�Y�]"����ɭ|���i4�[b���n>�5׮������߫�>eV�wc����L5���X������P�c�����Z5��TԲ�%�`>���ֽ�q�2(�<ȸϠ�ب�*�G��~*�ER�W��ƻ\Y(�v��H��fuҥ�|0_XB�N/`%��`��)Ը�	��͝�U����f��uilM
���2�y�R�u^��#sX�$���	����:��	�a�|���-���8�m}�2�8�a��S>�켏��{]7w�x��.2�3̶��x�&ry��SE�a����v��Y��kn����{ ��}��������FWڢ+i�id
�MQ�Mh#8N��[W\�nՋ�[=lKñ�Q�����4TӪ�������!u���c��Y��eW����jY�w�����E3˟�v1q�;�mP�h��믢�|~滼�^{l܎kG~��[>k���������h��KE���d�T�����MU��Ź�ƈ���l�Kr3�x��Mʾ���~u�ө���:f�z*^�UW]��S%���M��[�k;sj2�-�޾ago���ͭ#1��%Ϲ�.=mv!�������$�q1C������)�__�L9�߹��%�3#�S���E�Yo�}�v��d����o�%�t�G_s{��YMK��,�׈�z-ճ������=�NT�j� ��&ҽ�u�?�C�F���)���l?F�ŜkZ%���v�f����v��J)��.!���g�,%�8�;�!��[sy��U��βw�%�h�fU0���MCݸ�>����Z�����ӑp�C�q.nF��{jl�,�n�0�����\�ǌ�=�#�̟c��ߡP�SD;�X����h��%ِ�M��ae5���e�����^��yWP��߈�����)�&U�!L�is}+dSڡ�|��d����\�FR�ӂ��XԮ��gI���+���ܐ���s'uݏ�Z,��F�s�[1=uY�I���aq��7�p�Ph1Y���ZS���{bܜ�]���ڹ�9w68��(W.��q�|�l��5���=�h2b�q�\�s�;HcY1�}<��oq�;au�]e���g^�7n�nSg1��Gm�^۳u�� �A�t{;���ì9��W�u����n^�x7��Ky�:�te�S�E��V��8����p�U��q���֋n {'@�v+�.��5(�c���r��Ŕؚ�v�i�+}���+g�#"�[1�[���g��o`�T�:e�l����}��M}�-�պ{>޻R��y�6jӽ����Oy��Ȇ��-��9��Z;g�����C��ޱ�UD�L�3.��X�h���*��ӰϪ�oW�')'��ƣ��̶qò�d�f���gZ�wԌx��e�[Gռ��=h����{`7�Gz�>v8��G��vkk�{��Ð��G�����s\��#���&��M|����nK	}=�Yhƈh��<d�ږz�XXq�L�����׳���<�5׬4���֊|��d?�9h������Ʃ�����!��o܊��e.]*���1K8�,��S�g8���k˕���UǙ>�aǬ���g�?0���������E����t�p嫟���9�+��h�E\o�y9�̭��|�F�*h���j&�\�����s$MU2��Qhƣ�C���r�c���9��z�j�3�(�]���VC���y�(�fD2*t�z3�{�v�z���T�L7�6��}�G!w�ꂪ����*��_���Q��F�@۳߽x�ZX��4�=�al�)�t�2��ݗS�kF_&nګ�=�=����"�Q�y��ձ�џ;�C>�r���^|x����f����i�!��}�Η�_}���l#�כkZ���1�J�Ymc�#2x�%�v���>+�R�P���>iu���=,�dU��D.��/~�}v%}���
�r��O[3�KM��V�� S��ڝ��؋�׳w>��ս*1ˊ�#�	9q@ �S"��fI�(Z�ߠ���>�EA��'Y���-kY-vૃƈ��}�Yיn��f@|���*��`,����!����H}H}\�x�#���D�M���ԛ؍�)ܟ\a[��]s��֩��B�S5�9�p�fl������l��}�u�w�A��dZ5��/"�5��̺�����q���6���M�������%�bi�G�u��;h�λ��.H�>��k��}#��Ѯ�KDg.�l��n��k���{h׏Θ�)��}�f���l!�D��s�^+���w����6�O�ݵxA��7�tꉉp訉��Qz�\T���c��2�̏V��h�'���5�5���vN�?^�y��,5��i��0�^��!Ϯ��}�D���8ռk�j=�g-�5�&Mt1�{�X?��G�U)�i�I��H�g��Nz@c�w\��s�͡�p���89�j��v�Rʊ��`N�|�.l�=������/!��ŅlkE4]T��?M���G{�O#{0��͂��s���ۜ{�f=m}i�0�[<�>�z,���.>d�X�=CuG�{��^�MH�Kdt9��Fr��"�G�w �"}U�s닦d�7�;�Z�Ó;��e5㗝�<��vU����Im�]����_9��A���Ӷ~��"ȟ�s�;����,l�w ��T��-��.��#����8�n� d���u�>���cǟzCZ �_�h�}�*�-��Z���ш���.��?����]��r3\x��bE��[�Ҩz��$�K����ծm��z�Yp�r��Ǹ�H�٨�����Q�>X�����j���Y�ՠ}F�j���ů��a��M���22Q�����E��������f�I��U*H�����ǥ^�y�{%��2�*ҏ~�\Z1��T�qs�.�|���}���)�*�.r�9���k�D�S8�t�1����g'�h����������溚�҆L~+b�T-�ޖ:g�'�cF5������}6|�})�fT�޺��7>���2|Y��|�p�Z%�D5��r�ѭ�B��rx�k��w�%�!u�'%֌���|��_Z���xr kZ��J]��f�p��^w<�0�]jݞ���ܑ�p�a��v;VͲӘ��#��Kf�f=>�<�p�<�L}��j�c���AMw`�7m[nl����e�מ���󶏮d��,>���+��#e��c%�4}���ßd�o�2C��.�����8I3�Ø�i�Q�/�C%�_��h�}ϝ��Wo�	��;����t柇��~��n��p#�F>d[>w��g�O�q���2>���s�����4g���<���=Ա��b�"��&w��Ո��#YOYMq��2�l��m��g���=X�R-���s�h{�-_��E��L_x[E��2~��ϕ�+�Z��Xf@u�Eg��z�%KD�E32�/����k����������ֆ�6�<��k�߽�o�O#컹�����ac>j�\�ٷ#ﴴz�!׹e2�W0�={�b�gc���kZ��B���n��?
�-�<�T=�5n�]ލF�l�*û�t��[l*@p�Gq�rl�������Y6���,0^X�w=��ŝ�J���_>�k�3!���в�M��t�a������Gb`����K!�d���}m�h�py�"���}�Q�G�9��W����Z+���jjh��/���_�r���)���p��Z�U�N���o���d�k�pm�lY�j�]g�n`�q�e�ٞ�8L���%Zl�ÁͻBqdtgA�-��~o?����Lk�;��c=�r�>+��Z:��4m�%���o�]�l�:�-X<t�4}�睇;��#o�֎��V墙�w�Ye�,j����1�����k{Q��}qȡ�ꪛQUQ�a�a��jܾ�,o��3�M,�qߞ]�{�>�+G��CO=��h���-ï�>�	�֊e5,(|�V�*�賬�Ɔ�����<KPr���>y�$��jr�.�K歄���f9���\jA֥��Q��"��A�����ܚ��~���f�����P�aq��,;�M�ϝ�kZ9P�k�AMy�V����ECJMQ��B��M��|������5��q�>壌�¦��1�M�g;��<E��E5L��g��e�٬��Z�~;���3_h��!������5�XH�=�-�8���"��t�j��i�V#�;PC�[���k��}���B%�}wH�AQo�׾������9�������SM�uy�g�K��-}��d��b���P}D}G�Z�������i�P{e�5�^fI��1=X=0�Gn������JT�����.D՚m��r&�Am�$'��s$�H]G�og��W�(�c��s��sۮ�uٹ�g�s�Kv���]z^N�PM'n���kjl��A���+m�OYgg;9F����|�h�6��^��'v�NuXnՖ�m�uFr�]N���nǎ^�:@��1���M��<*�ѹ7)�Z�ƹ]޴yy������pᮄ��r�<Cv���s����p���箓�Z
�z^�d�:n.�/5ڹ�z��s�lF�W\�g)m����R��V7s�Z�Pjƚ
OkoSqF�X����2Y��{|��Xu�׎�h�B%��}s�h��K�*උh�����;��F8k�逦�MW�|����C��"ab��cE��*`��D�'35UNϚָ��F\[
h���M��~߫�T��������K>�J羫,�7�Bl��,��[�P�ߦ¢1��m�L�[~���f�-v�c�y�}W>�5�Ե�>�����M�1�U54^0ֲ�m�2Z;�}��f�"4zaγ]�{�Y�Y�E5s�75D�pƼ�w0Ư�m��y�����S�q���f�ʘf�p���2�&ݯ�5L����34Z>�!� ��m�s�}�𥉉��{}6�͕��p�6	/�cE��O�g՟;D�"Z�KD���{�XK։z�9tϙr�Y�r/e����gz9R�Y�ᴌjY/^j��W?'m�	ҸKU(�K靈"��y�
a�{���kD4CD1���w�e}�-�>�[D4CÎ;��x��y�e>�$1����>��/8tg��}���ՖtV#J��*��jbZ��%ƶyxTr��IcUGdjSPD��T��ό��=�J�������8Ad��Lk5����T�i�K8�{2[�@S�=!�&�}��.�s�k�[E6��B�����~e������V��o���7ݜq�֍~�y�x���kG�g{[Xѵ��7c�Q��3��dޅ%��F �K�R�h��h���-�9]�ȉ�z�&�����7 �۱�����'{�2�Fp4�:�K+i���-�����SI(�]c�o��^1���53y;�63��?dC���Y�9k�;[6����~��������7����ذ��3�S�
a��e����gZϋ������i�����yV=&w�o����J�Z���D5,sS9;>�ю{
Z#�5��g����"��2��v��^����E�a߷��MGZ!�	aY�_}?N���ؖ�$:�X[��1L�2�X�q����(���?b
��f��2Xw�����Y�q�Z&(��ǰ�>ϝ�:��"����%�w���v�|@U�To=��6~���-�4g����#߉�>��JHe�E&�,�U�k�x���)�v(���aY�Э���ͣ�k6��,��q�o}��Zu�s�-����F�/Z9QL:�>��-l��#�]B.~��_vH�?n�ku�ۚ1�x�����{�v�+t݄�ܫ%�e�]q����릸�4Sߠ)����d���a[G�<�e:|�?w��y�<ԲZ2�c�nʎw�s谙���ݨG�*�)�����;kZ)�Լe�kY����i�5P�j�bh����[-��wd%�rͨ���v�3��'(����6��D��wY�k�g=��ƾe3��`9�o��q�?d�V��9�8Z1�:����շ{���9=E4��Uo�ətR�3Q�S5�kKE�Ͱ�����ţƥ���_2�͂�\�a�|�v�~���~���v���bo߯S���PԏZdw�i��q����b[�I3����$n�ڂ��6'SNi{���/G���YshK�����P}FҨ%7l'эU{�g.�g\��v�&
h��o�J��6�j"H��ь�̂�-�gWӏ���`�//����L*��wݕ�߻���)�6
h��k_���S���
cg�U�����wcWy�ֆk�;��"˨\hۄKZ�j������Rʚ�T�j�G���9$�j_j��ܙ�g����R��ʩ�������{��3����!�	t�d{3b�����Z�5��Hc\~ϧ�����W�k8�seղYmY�{=�ﲷ�ہ�;Fzk���.�n}a�1���{��Gd�ֻb!���ny0�q�\��=����"%�����}������Vճ���]�d���j�Ʈ��\�<����~�z�Q�|�ߌ�ǝ���1���T��;�ry�;׍q�j�Y-c"�??�肢$��SPH�h�kZ�t�L���>��?E�]9����}]���2�79'��lB�+t�cD5�KD�a_}�;�q��0�6VE�E��f3X�y�-9�5
[�G
�>��R:�A�iUDT�E���&��G~���c/�Tћ��d}�9�TY<�g%��祖{���[T��2�>gv8�j���SF���х����ֲZ7���艑éjbj\�ш�q�K��7���}�����h�s�w�	�9���{����(�m�&���;��Ǟ�R1�;�X7/��>�W����c��Tj�A{ƒ�Z�9�7EZsw۔d�.E{�1r�^ii���9�n�
C�?�ڃ�J�|��1U6���8��>_Q����7��ͅ:��[��=�cC��g��e�ԕ�X�>iq��W��mm�mS��-�jZ9P�g�j��<�+��۰��Wo��KU�䶋u���,F�]Erj��%����f�������:�]��Ϯ���U����rL�v�n�Ɉ���s��-Q]6vig��In
�6�F�!\�f?��j�L�T�#�~�	x��B+3)S-��zܨ�م��_\3�[\9�5�d�~����{Fp��}SMy��r�)�~{z�4�=P�k۲}��G91ɘD}U
����b1�1�	hϳ�-�缹�\Su��/<x�2�*�-=��cD9a,�|�� 3�wϞc�}�F;!�;kβ�g�|��ƻe{b����:�~gy�cϻ��"*�T�%5F#Z!��]3�����n�6����ޣi΍o���h����}m�f7�eTU�����Ew�;	�����瞐��"����c�5�d�
vֲ�7{�ϡ��%�q0�4���aw�&�[�|r6��Γq<귬:��p����̅�|�{���~4���N�3�9�7!y�����с��P�uu�{�����)��c�Dr��W�������"�2��s>�8�T���æ�"*�:ֵ�)�d�[a�~�-Ϫ2ڶ�g��w��T�2;�#�݋F����c��������=hsy�Pc���B$��,���g��)��nHhh=]�Y���s�NIq�{{H���	98�_f=[���t_R����Zl{f�֫�F��]�k�a:�>���`�\EIr��z�2�9�Gt1{�����3yZ�<��U�y�Ȏ�Gu%gO3W�I}㮡x�w׸�g�bm�q_mr���.��W�x^�-ؒ�)���d2��p|2�����7���{ɾ2�01� ���WR��&Sė� ���6�Y���+�A��km��ř_�y}���"�?g�OG�Ң�!9gj�WM���!\m��+E��������E�J���:�FS����XVaͩ�%}�9��Q*�<:W��0q)Iѽ�gh�n7Xo8����̻i���q׍�)�'��me�j�\�J�����\7�Ձ0]����Q$p:�����y��$��v6�̪z��]�n���g��R�8�������m��^eu�z�^�;K��8��"&��6�>΅v��n�j��a��Kw��C��V�L{�LZ,tC�VfN��ѭ�h�K�ݍ�Ti�2tP��+ea���Z������"���8��i�з��:%���ib���ݣ���m��-��s as�=1�+pe��.-8���0o�wX�Ȇ�Y͈Lpe
S�n����%^
�v	�Vz�Z{'X�j����کս��r��=���)��)��r�J]ק�Eo^�+�]O��n>f���4I<���` 2��I��{as�T��"n_-�sP��(u�����3xn�L���� SM:n�<��q�V)�fّj����P�e�k�MAt�쩻Q�t�l���^�ds8�����
�yu��Q�g�q�x9���fێK�4�ۮ6W����۴�]9�%vۋ���Z�� �[pV'�v���9�S�[���tq�<K��If.С�t��6��3<������M�lu�S�۱�p�n����ܹ<i{�޴ub�/k��sgv϶���q�Q��������n��"͓�<�pr#�<ZK;��`ۏ6\���N�z�5؞�ܖ��9��ڷ+����[l�p�';��p��6S�u�W��}�%��={��V���8�vʽ�m�㛛6���|c\�ŝe���lL��ru'Om���kSȋkkF�yzPH^�9��a[D>y7�ŧ7e�ll&ٗ�,A�/+z9�+Q�K�����cg��=H�p����&-�YГ��W�-S�rFÝ��»�f�S�q���]��cl`��nyo1�A��m�Vj�I�'<m��(�Sn��s�ԙ0{看s�-�h7<az�욷�z�X����l9�1��U�{&x
Ss��c��c��s����r����Ճ)�W����+��
�ù�U��IM��7d�g`��<vۏ<��g�J���nӝͼuU`��<W���(����35���v��7n�Q�{pms���r�ڎ�q��ϝ�DNF8��m�^�����i1��G��ض��5�Z��Fv�����Ā��9;mQvMp�wm��v��n���j� ��-��i8�Ws���t�p�}�+��+���$I絺����6�Ѷ��!�+��-u��u[��v<槭��趲q<X�y���Lg�����v�hkqn�]����m&�V����y�k��P�u��J�Om���+��޻����!(�1�ƃL�8�g�l��5R;sR���\����<�mx}	�-O�ǴV��Q���<�֝����r�s�uŸ�뛛ѹء�捄.�m�"�b���m�ۮu���{h^�V#�k+z��p��cswA�K�Ʈ�oZ+���q'�s�5���:n�\����z�s�t���*:3����)�L�(4�kW\k���;��=n؞.R�Ƙ�c[�ݶ�����t�cn:}�	At��=�v�7*�|^�/=ٗ�CΟL{:��ֳ��&�]��n���0��a��5,1`q��ޮ�]n�K�/)���n^ݳ���d�k���Ӳ�n��ͳV�xּ�f5�\s~��!uÍ�}6�h��.�XSG~��h��*��s�c�p�\)9�۵��y�m3�{���q�nǘS��a�\��Y|���B��!��)�;U�u�IE\e�.=}=P��ǯ:h�kt�c$��zb#�K�k)�V�Dd�\�ڙ闞z��KZ�h�Ǎgs��y���1�Bn�T������k�����;�ݬ��p��<�3�� �����O��~lLd��h�Ɠ��"�J�݁M��|��-�h�B%��ʟ���E�٦�>����r#��Ӎ\6���wK�q�9j���m}����Y�O�.�m}�)�~�����2�TT:sS5�q��a����rb7B>ۿ��c�S�u��E�
��y�Z5��pSE9a�{�Xz�xe���5��I{7��>k�x�##Z �D�����3&H��ڪ�n�E�ޗ��m��1��0���s�o�KD0�,���9���/D�KD�R��O-��=��b5���&Ƌ���c�XÏ�r��1ۨ>�o�C��7�>v��~$A��!
r��;huz�x�7lFת����7.��6���ʣ qZ6�e�/�W��g��X��0��}���ÍѾ�E2Z��޻^el)e5��Ƌh�����mS�2�O��!=�.kӌ�����Ѭ��ɹE��Ʉ\��|�$TM:�"���|�&4[�>ɯ�Gq���YkY���u~���~��X}����^ץ�Jl���U��ێwwO	Fk��f��{Z�__K�e���-j3)�v#{Ŭ&�)�����������W�� �w�������lJ)�����0����ͅ��a��amK�Ŵ{�޻#�C֏����foXu�Ծ3�Vg#�N�&�����Tш�SPSE�m@S����h�cR�sS��k��l�9��
j�}���'���8�n�3vkKF�C�	k+g�s܏t������q��Xտ�>?6�^��H�\��"� ��׮F�-��T�'k99����d��j�3n���d5���2��[����YA�֌w�����~�}�\֋�_�5�b�]B�SD���uQ q؊�e����Vڏ[d�z�?g��Ѭ��MW?5��G�O~��/;׈����mg ��s�C3��v|�*8�3���f���oӆ�g��~�E\�0��������D�H�\�z!.�Б���/d�m�{�yg�,����@����f��J����w�{��َ���O���a�5����f�8WyH�cW�Ϣ�䢟���v�����w�d�Y3\��E�Ӟ�w�6u�1�c���^���X˸E5^���5�}�pD�QD:��**h�q�虜�h�O�r�>�o�a��w��:}���>�L?�>R�?\��w	�}{��D4CD9aﻞvc<��Ol��u��m�yَ٭5�w�ܝ�/_��<�{4s��'T�M�C�a�ӴcZ�h����kS��F�<�S>�|{(����f�Z9��j/��������%��
�����,�p`�El��x��l��]^૽l��T\��kW^܇���P5{�`����#e$�&��i�Fh���w�3=b����:j_]�w{�vS_l"����kSp��|}󨋧5�j�UDM�h��?A���%!|�T��6b?��}R��?m���h���}Y�*#�֭�9~�E��gٚ�=�u�������_3�̧ܸ��h��{Nя�%��K1���CnVê��UU5����B����}�H6��~x�3#~��3�(�s��y�{�����S֡��e��S��_}�p�㈄L�d�k�������Cob8�M0��&<k��>c�r"^'OrO�n�=O%���C=>xLv;B�^�b�ݨ����q�l��/�C%�*he�v�]��SK;��%�α����Xc�^�V4[P���߰�e��"Z���T��I�����\^l�l��_y{����N����\F4o.=����ύ#�+�(���s���ݵ�T���W��P�C���ϡ���Ѭ���ɽ;�*kY^�S6�g;���"Z�KD�����������L"�]�����B�{��Ɉ�W�矚�E4x�{��GU5TTMM9*��M��2��1����?�ih�SR�1�r�����ߪ/��e��c\�or�~���K��������2~���k�D�w�B�-�s�ad�5��K	kzAlms�z>UK�)�����/Z��t�������{p�3A����ӥ��vU�W�+̶����h}�D��KD�E��"=�Xu�D�؆�@l6nܺ�]�"Q�;�˗l�Av���)b�L�r��������T��0v�T2�Yo�E�q�]��av���ȟ���	�X��M�!���[zQ|}���uU��<���m�an�rCL�a���kE�SZ�rQ,�/��_C�T�^��-��KZ_$���Gn����Ll��Bڧ�����.rSh�κ>kY�[|9Vw���S��nq�S�*!�����s��s��vv�	@�r����ޅv��puW���kk��2���o����{��q����{�6�e�4=�R;pC]�r�����m�>xW��߫ח���ﵢ2��-����Yֵ��v�Mq��Þ�ޒv\�L*M�5~�-�ް���Qs�����w�����M]g��̦;��3:��[�_6�^��{>��Ɖ|����h�}�4�.�G�7�k��j���)��5��$oND�)Ӣ�MMV|í_ 鐎sf'$�c
�9_o_ާh�u�a�E�y�O{�h�D2���]���~����D��Vn̈́�7��{P�]�O��գ=0cT�r�\����y�����v+B����.=*�J}����<g�˟��.+�޼>zγ�Aos=�F2i�ޛ>4KX�h���A{�
�u�2����^@?��O�W>�C^g5�vvaq��]q�V�?3K�}�l2I����虚��aƉi�&;�\"n��mk5����׶���sOv{�w���l!��&���1��w�a�Z%�-S�ʹM��6kZѧ�QMk%����>�����<�f5���=X@�tUϩ�>�^���h�>����ev]]tnf^��x�-�%;���/ޡF�Б:����ַ��p<�*<�d��j�<ɥœ<v�D���G�~��v{!�t9w3���]w'!�\[o)u�Z6�f�k)�u�ɪ�n<s�{�̙��	���#��G���סm	݊���kB]Fܮ[��'��<$���'C�y��qs�n�[eՂ��۫f'��=g���۴p`�/5���m�qS�1�ez�p����n3qt�8�s���\�Y��tb�6��-����v ��7/�ڰ��{\-Z��.�Ӣ���<�]�$�!�.#��4��Ƽ���~�Y߶Tzc5��9y��1�2�0�6��v,6Z{�>�+^f?}�V���"�G3�ɹzִv��S[�������W%e��w�y�1�[%��x�c�=y�"Ѭ�:�J��".��������8\��&�k���|�h��`�}��-q��������rq����l�_B֋�Q��~�{ݎyk��6��3��]�r�)�7,r��'ٮn���{kg���督Y͎2�-�5��}�4C������v����h��\�*�n5��M�C-����~���gr�܀ۋjYL���r&&*j
neԱ�S�kY����1�/s;�`�P���ε�A��v��w9(�cS������vQmu����y�6�s�}6:�/�9P�_��7�ka��߶l}�ǥ^�iu׬m���v�+c�YH�� ��q��v��d��G�꺫F4CEL"Y{�_#{<�[���_^O���q�3��e��[�-�}�qa�S������!���테������ε7��[��
%�
A�E"���i��>��;Cl���.vk�3���]��;nrm�<�F;����N�j���CG�/�ª+�}6�fK�\u��g:rW9�s�h�Ű��d�y�Q.\�)�߾�a�Y�g#~�����}-KF��t��V_}uh֥��r|�5,l�[^���i��Q�aԺ���ZӜ�-�2X}q�w�6�����*��<B��	ǗR��)�N2����D<�m&*ݮq]۹e�gn�����*lR�p'w1�޾�7|�zs�;�D�{
���g!��
`�>Ӯ�F_��2#Z!�	a������kG{Pn���jk��Q�ѵ�'����[Jؤp	�.�n��K�S��a��_w��h��a.YUc��U�Y-KL���b�y׽5�6g�{��k��֊r�;���h��>�>���L�������y#����&�)�Q34b���Y~ ֎�oϏ��n�㯡1ln�VSZ�L6S���M���-y$5M�-�{�/���_�S�*/��}�k���cGn��e\,k�nB)�d�ol�}ET��ET�MKqUXu�?>�0[D6�����G;���VB)��?]����_go&�վ�mz���h���٬�}>hǗ�>x�g��Ƌ��ʲ�4e��)�Z+��g���o�Ϯ�N�Ek28�@�DpM����f4�7�l`����]�:xN��F��3��$���a�5�D��nY��g��ߚo��a[E�"�z)��r�ֳ��z��HHj�ߜ�|�~����>`T�y�8�~a���ʋ��!q����k�󦊻|�3$��������n��)�_�L&�{^�8b8���ϫ���fLqq��,���{|�>jk��h��r����T`C�G*-0�w��c7!{��p{��W��i� ��S���|��t扚TTM>#vd�,�[T�fӋ���Z:��-�ʦ6������:g�|y��{_n׶�i�4�t����Y���u|yU�u�໺���K|�����u��X0��:^f���f
�9U�q�Ob�t�:�֊v��/��8a/�������kK,k6��fLѺ}�C�*��STɉ�qU��\�4}q�}�o':����:�h�����e�J��=ٶϹ7���Z>�"Z��P�~��
�ﰰ����F>�����yϽ�F���h��gk
�.4DT��%�½���uLĕ5Q#���k�|�P�v�X}q}�e5MS4�E39�=߫�����㿘W#��}�h��Ik�뀮�u�c���`-��9_{��kM�I�KR2Y�U��6q��r��c;Qx��ѱ�H�W�U�[U�l�������s���x��9�ݺ���ع��S����5�Ԗ�^>�ۅF����0�|�;h��p��S�}ʴUrQM0�s}�N�nw'
��f�GXK��\6�����e����a��a^���܆|L��S,�QC���q�;�-�ߘK��V}�b8ƃ������{w�P���˃{8��R/ d4���{��!���h��F��o����z���C���F8�Ua�a⋇��̎��ds5���5��|�:ly�3̎Eo��Z5�Ks���Ʋ{���/��j=�#=㾎T����4vo���k�:���_���z6y�U�5�Pu�j����;^�ɲ�J�sJ�����浞o�$Ɗ�ۿ�]��i�߸�}zֿ���m˨�-����󑫟�ݢ>�E5;.j߮���VQ�[-��>����ϼ}�S.�s�ڞl磙���)�1�h�m=���*Nѓ�jx��6�vT�5�z�s��'�Ѓ��F��^!l���=�~��b����Sү[j�)��1��T�5d��<��G&�o�_�я[g�4l����go��;ݺn�ΧW]�G'�y��p�㘓-�>��56�q�0�"ٯYy�ݛ"|J�Gr-_ᶮ���ߨ��VN�`E����0E���f�N���;���2��\���N;jL��4������������wu��]��ϝ�Y�B��>��[+У��ӵ��F�d!�U�ݴSߢZ����9N���xY>�}P��5�a�������-h}Wwm��u���{�Ԭl�9qت�>z�-��Il�rs�Yr�_�㓳��ٱξ>�y����՛ص�B)���5o����}�Ü�a�:xv��}�_�͸Z����V��뷽:j�5���~c����#�tE9uTj8�2Z%��k���Z5�Դw&�XK;*s��h�x�/3�9��P�|�7��r��,1�1�S�
5.�|��0��F�����ϙMX?��G���d4lO���xj��˩俾ȶ_evc7�Z5��(h��h��ޛE��E3��Mճ���&Ï�vQo�%�*�9Y���r/��k6w�f5��9�t�����)�Os�w,RXr�f�����c�c-�\����5�=�r�ϲ�[E�C6>ظ߫��꿧�ص�9�R�k�h����q��gv-�����-��K��ϯ�ݟ��]�� �Ț,:�4��`��;�Y�b��&l�δ��|��t������7�&@�{5���Β�\3���b�~�T0�{u��>f�{	��E�����#̵<@���:����r㚫y��V�k�KW�s@�rը=QWn�<C恠%��:t�n�^.��a�v7n�xݗЂ��/n�uv.��q���8�u���3��h_>��SW�����y�]���gk��N7?�c�/m��vh���6L �	r1�]t��[��^Nqn�����D��Š��vY��A�s��ݯn�sνrI۩�:Z��8�[�.À۫�L�8�3%C�TTEU|��L��w͐�Ͼ���kַ��)�����>�͢�}aM��_�rl9�G�9�"�i���L-�F�ٮ��B־eYr��
k~��|AT�Q5L���Ƽ�f���)�}�����f6�����Ó�y�K0��Y�=�E4]����Y�%����s��^{��b¶8�NXKZ� �ݟ��(�b�p�o����t��U2�#��t�}U.�e��x�g�]L��0�v����;8�0����H�S�A�m������:����߼u�����}:Xq�h������j�^���Z���}6iG�5^���E��8�C�U3Qh�p}��n��"{��_������O���Z8̚��D��
>��N��B�)���������a�Z%����w��՝��d5��nm��KP��Y�����D�M����kU�)�~���!�*c��yN��y�h�A��}����+�W����q�c���E�o��0�|p�l�,'_I��S���k�q��o��NJ־g���F5u4sӰu��嵷���;ƫu�����6�H㺞�$2&e�쳋����k��T�u�����G�ڸ��n�h�6y*YM�>����=�h��֩���)�?W�Sh�9(��A,:���{UXnT��{�{�oe�_�y�P�#;>��녭��kvԺk�9���[�P���^�Tg�˙5�������5�9��߱�|M�A�a�q֝7��Nܨ(�����|9���S�Qƛ��݂��f��T&��/�L��Mk�r�Uă-`����q�Y�
��ڳ�g!���CE>3�8��N��Ɖh�墽ﴰ���*l ��[�5}V>�4� ����4�A3DTI14��WM;h�K�S������/![E;a.\3��ӥ��8�=�5�ۃ&r�<�F���6-c��-��[���m�}�g�kG����$��2���h�����MDUU��A��-����}.9��K>o>��v�dk3��kF��)�܅���Xk�E4CD4r{��N�}Q�@S{�}�Ǿ����^���e�h�����2��}w���.h��I4TT�aOZ�SE�"XS��ϝ�Y�n4]�%��{��_�l�מ^�W�����)�*��O�-w_o�f2_0�[�m�0ѝ��|���ꃇ�1���U����?�������??���z�7a�eR���ܹ��ۺ�\��D���`��:��ls�B���n'[b�����q��ڶ[W�v�������<g�ͮ����K�S<ӿ�9V��F�r��ac��߶�,+�y����}�o��ao��[��zϽ�1�mkG�u�S��϶eÎU⦈�D�N#�[%�]4K%�����V���}ڞ�>����y�2��঻��UXq�B%�����c�+��W8Xu��>�ˏ���q�
��fϻ?z��"���<��'�")�Qbj�|��_}5�F�}��a�ξf��mk/"��2�)�5�=�}��_9ߦ��jϫE���{h�3n�X�3Y�����&P�;:'m�\�i#6�s:�yovf�S-M�\�Â�3�[#��[��y7-�p��\�k�ڶ: �|ի�]�� �x�������o$4\���d�w���B��Pf�f��^&�E��v�(�ȵ�l,e�����_Y��}�d��E�po[��\ú�b���Q<��;p'��5��WN�0wH�N�L�q�qֵ�������d�A�,���B�'_�y<����P��Eq�9������J@���6w'@��Z9�ufb+u*��q��[x�7��cY���r�f�6�E"���(�[Υ��e�Feql�U��p�����0��3Õ����xm�v�Hy�Zb��n���]�;%�8��'U۵3.����0�:>�#���V)0���c]@��^;y�*���5`+Cw��t��3:�%�q�'"��˽z� ۬[L���b���*$5k٠�&�FB%��^�)�� ?����=�j�}Ds��x���XtszC��m��)�.#E�v��M�d��[��ל�97�֭��J�SE�Z:!������[gJxrX�Ђk8�T�+�}�%K�=�Z3�W3.�Q���b�FN�k��TD���"ݹ�'=ϻ3��	s��fGڗo%��T���RD
=����PHyO6�m��l6�{.�yPTc/"�b��4y+1��ǲ��_2�E�'B�ؙyF���[�y�d3_v���&p�je(��|P만h���/]��9Q�a�{)�f6�������FK;QL�ר�u���| �I&Q.��g(�<56��N�vJ��v��~��ތG��r�fU�cq���oH8�5��
o�
�kjэ�����������,p�>����F{gf�Lq�a󜏦�Z^ɥ=���L��t+���]z�%�^���^y�5��ҩ�׳�iʿ�n.����ﺳ+�>cu��p����`��O�a#Ǭ)�@6k�F��4}<Ϣ�T-h�qY3���P�}eu����qv_P�UM�6�nbq��<�A������v.;��WJ�k�k�	�a���AM�T�j&��q�e4K�î��ۛ8ֳq¶�w%|�p�TZ1�90�zõ��l9&P��*L�)���!m����xY�hڊ�>�gy'=y;2��UQT楺��F�����D���c��q��/�}eǻ|v��n/��Y���0��73������jY�-|��ˋZ��q�?3]����������h������o��!�g��[�O�DK��uN�����5�k;ϻVq�_��:�9�N�{4nB��l�S��)1��v����=�~�mo�Ձ^U�kߣrZ����]�)�`ώ��B��aWa
*r68w�T�uZ��,�"����z���e���(�<m�V3K�ٱ�9��9�u�.)��A}����k� �fzh~�;��XA�f��'�B��U�\풛#4v=S`މ#2�⎿� 9ֶ�)|��r�yޢ+(��D�b��k{y�Uma��*��-[��E��_7�}C�;W�`;8�z�K�i�º�'��^�� �K��8��gWu�kۮ;�=U��0���%�����t��{[�iͧh키z�>�ޮw�=��Oa��Ґ����u`��V�y�j���N��5ػ�&�9WP�%�1����O%�_���}nW�E>�-��)�Qͯ\;�e�yx��S�3��k�3�/����
+I�I`:`�xr�̩���伸�ݜ8;�x�l{7��}�<�Ղ	�$	U{{���rx�v+�W"s�c�m���U��c��f�����ڵ!
c�v+����E���}�>Otm<+�t��p���E�+0����9x@��i6��v��)��|�{V'g�v}�6#�.R��WJ��35H�k�]-_k�c�-N��O�.㕍A��ܡi��[8�R���-zD2�Դ9
S���t��`ܮ	X�V1j\�^�oS�9���!}���ry��snMH���$��[}��7��-@X.s�r]��-���8�=G����۪�#��l�g8������^��t�l6��g۫fx��Y=Dv�#���=��p̅ϔ+��4'p;�����L�i�X=7;�V�o�c�y@��:�Oc��o�1�YQPӻ�N��LMd���k�n8�m����S#�o^;Z-�q��,mP+�k^gݹ�H�|����e`uX�XwlY��;q�;]��c�-�7gqs�ծ���S�lO.g�ӧE���~�N+�O�W���L�j�����0��o.O/m���q�ׂ���@mr���١B��I�Nޣ�xo*���R�N��1�)�n4|�Q�鵯�lv4�gw�e_���n�u���r��5�p"#(
hISIe+���{���+�����͈O\c��V��Oz:>Ӑ����`s�Ϛ�O�LY�2P �����Y��^�hW���[��sw��.�2� �lVnތ�@���It�w���#�Uޞ���
�t�I��M���d-#�X�l���J�אլ��vcE�vidk}�l	�I�`u�'��*4�#�ӻWV;r{[����K��]��s���X�H���L��e�,�V�巄_�[�6�R�xO��ּ��}ͱ�'��������ZѠ{�YȞ�ϖo�Z,�LJ�I�[|�v;����GI���Y�L�N^!r�bY;�˿�6(L�OO����V�j���3���W,�3~˻���[Zd��+f��QlK&��[�+�GL�R��-F1+�K]Cp�ja��yS~�-婳a�p[I�=�:x#�ASt�)����2x�1���龇{ �ӓcO����;��xx�K���������I�H�@�-��gN��Ӌ�㇯J�ͭZ�"����%��|�yv�x`h�C������%_�������)�������C�۱{������w�2����(�)g^��{�<97�����D�po�']5oN��֟��
]�j���ձ�ٮy;<���S�k�����6m⫢�I�IZ�7k�u�����>?���z�K�7���2���X�������������{z륋,bיKI�YŶ^�7������tjL�;����{�P-����ǿF|3P�y�7R���T�t�◛wk�q�@h<UmRM�¨O���� ��p������6n߂F���^�+�lJ�j�n�ݮ͇tF�$)���ˬ��K�<<OQ�.;s�ԝSv��X�	�+Zh�#����:�Kv�=���{���=Y��(�S�S�BI��?IJ��kg^}m>�禎�3���ۼ,bG=ݸ���#Qu���7��ݔ�ť��O�SU۶�m1��(�d��f��z���9c�1�cb���i��k�ǧA1Ou�ͬ[�-�<���i���;�}e����J]�\�O)l�'E��x<�i�n�;xNv��V��E�+7V���7N�xU�����W7�X����N���:�����h�0�黇��]f�k�F�&�N�l��M�Sg6M�o��y��soP�Y~��C�(~y�L�4L��h�\���u��*��i�A4�)��i����U�0�-����۴��ӡY3�,�Yt��y��5q��?*�c/;�}�~��rH�����3�s����=��Iݓ4e�B&绻�p�X���ʱ/��-	�/�3Z; ��N����m�M�g�P�S\L7u�D��g-�T[���������_��5)Z�1Os��Kwd������wa�4;�� �i�M6�eD�a���Z�~c�n��d�gz�ƚ�%��x�UpD�����,ݜ�����_���;�MO���5��<tv���{�=[���m���G=m�}#���n����`���7�Nu�� W�	�ĲI=������zQ�3�p���p斈;���?�YQ�m�}\r�Z����k�;lTf_��oT��LR&�{ދV��~jC�\C�����>��~Ă]����)��@QA��m	��A�n�ٞ���Y�����}5 [�*��]�I�R��_O$�̡��Ȥ�0!�I��}H�vy��o�\;f��0�D�zX����.�}��wB�Q±Fhb��.��H=sȶ�`�/0��F��[kޙ�$g=-L��%x�V��_�g�!3��>=o����Z �lc��Z4�M�.�pg��u;����\2�	�Z�5��+2��[p����B���%6�5MYҠ� �7O6G6���>��u7�9����H�M�������䀞͉�<뀰�@On�@gtmt%�F�S���m����:{�'Gkʹy0�[v6�:�
E�b��}����ݴ$������r,guv��淗#�Ftr:9�c$u�����us�Z��č�՞'���i����v��7,�7�;��l���֫�[vd�=u�i��v8u���m�;<`�K��Xn�A'#����-�=�;�����q�s�gg�(�˘�b�:#�p�k�Y�u������n��~�k����ۜw�=Dǽэ�.�;��;ނ����G�e��p�2��j��%MI&ǬQ�m��{}ʾ}�Z~P�s���Nwr�]nYL�髺�¯�{�პ�J�aۢ��l�)�_$۲m��5Ҏ��z��v ��6^L��&��vy�<�����<꛲*�9X��<�׿p��G�~��ۻ�G�9�����u�y:r��[�'�u{g�>�={�gVQEs��x�uy2�`�BtwT��u�a�C��?k形�D�|�_�*u�q��Mz����ד��W�o���X(�r��{s�s�OnzC���N燴�Q�C�.��*�su����u���3٧���?Ưzf\�3�q��-�Td�Q�J����=��f-�T����^+���ZݏB�$0�E too�oVG���	�׾���
<3�a���Vc�]�uu���8P�y87*+ى��[�����S��Mzg>wz���wƴU������O#-۬n� �m�<�y{)�;�}���;wZ��|�^�d��:J�D��I�@��K��;܅�;s٬�ww��B�K�DBo��^}�Y����y'(�ݔ��45�"�K�(P
�MT%�~�g�f�s�W�����tMYT���f�/��/��s#L��c!p��m��}�OUH��
���i�_ͦo�!��smz��һiB��"� =yG��;c���ǆ�7w%Cϗ�.-8�Ųd��˖���D|.�,��������i�ue�b��j�m���n����4�Ԋ�()%��0��l=�<��Ȧ�'��/�{<�z���k~�������h���'�9�W6Z#N�S��Ӣ�l;����l�yW�{7�C����!pB�ymO'�nMɽ�g�Aw�\c��9��P>t=�1���|������tT��Tl�rD�y�,��[ópF\�o��VWz�ݥN�(�=2Y|�M^՗�����z���;՝YFIRG{�vM�Q�1A��<U�������C[�ڮAя�x�֘�c�����9�ײm�u"��M"7�}Z�g�ﷳ\�����/���rY���O&�S>SGLC��Op��m%��y�^�Fn�V��|�4�[%���6���u� �+A���^C2�{4E,���[d�{�RD� �V���:/��)&��P���a�� ����x�Z��Ju���Vt�5s�{N�5ٛH��IPt(:lRH��w��^YR�pۼ5�gz�t�����w�	��{1g�؏��M����^~лʹW��@�&��q5G{:T�]s����|dtx{��ƻk��BF?G��B��.��BU���X���^=�ߊ��J�U����I� �b�7�Κ٫���W/J�����v-�}\�GĴ�����v��P~��n�w�U��A��5�������E{��~�}��ݧ紟*"Ԩ0��>�JKb�k/��� ��M���˿-��1y�?l��(
7E�I����ȝfJ:���Yy�l���U$sH�A�=���u����]5��8OE�4��gW+N���ɕ@��"�c%��\��])|Q	�N�1�U\�b?]�vC9�'��'V4_:��lL�[���{ҿ|�ѯrr^md�q�5뮰�k��\q�3Ofٷf���Z�
=u��uiɷ�<]N�M��h���Nzie�w�[V��yi��4��]-ص����sG�f4wҮ\���Z�5ꗈqh4Z�6�c+���
6�/�lyN���mį���o^�����tKӏz3�����מFa�d�3�c�ܩR�H��m�t�o+#m�p��y^`2Q��g�1��1x}��z���+�!9+V�'\�z���2
.�4u6���,
^޾<�0G�� mk�7�s�j�
b ��uT�ⷋ9z���$���'�R�)5@��Ŧ˹���N����NN��y�>K�hX��G�o$k����Rꪭ�T3fd���`	d��2�V/z,����)B��Ltb��n03���J{����d-G���Ќ��_j��s����ܳ���x�Tx,Kh�w얋=r���x�ݐ���8�}��N�)�Xv�i(V�ʋV�H���I�����
�e6�3O�]�kjv���B��%�TO`ɳzv���s�Λ���o����/��j��򖵚���y�%��L\|��ѱ�M^��v�-192��H����-���,n��:(���1M��Ȕ%���n�h��:Y%���NWs�}���etޫ�E&� <�#���b��e� �ѫF������Zd.���S#��H�g�q�}�2���`���K����%7�E�o2��v�U�2���wصRʌ�+q�n�[2�]`�k�h��jFr2j2���U�Ӑ��	�:ڸ�`��1F�Z�v�\�yS���t��uͶM�f����x�p\`��"J
if��N!h�j����1��c�o^���4���c��̻,�_���wr[���fgWF0��ͬa+�~u�%�M�[Y"mk��n��
S�]l!�|s����E�*�S���;{}��f<J�b�.Z��SˠK�������r����Vж�;õ'S�ԙt��ݡYqm����&�/�3<�1��� Eٰ�������И��n�3���2��Ռ���/:���h)�n��
�������^��g8��w��I(MFI#q�X���ua��=�\!m��	]��&�[����lq��t1���W��t��itq��2Hgk����l��ǁL����n��� k�c�v^�c�Ѻ����]	n1ڬ�֎��-��ۋ�9�(\F궁�ɋG��D��n}T�q��79'��063��{�F��E�]�xە=��݃ns=Y�9*����\���n\p<rɟQ��g��s��SG.4]$/=�����v��`ؔ����dQ�WI�����G]�Yә�s�GU�::�R�c�1����XN��VLΉwn�]<z�&�:x�̧��c�c��r@p���oJ��(�&.���c۩����q�⸔����9�t�8�\t���s�gJ��h�7c����n��K)m[u]��y���۝�r�Ů����;=m�oD��N�1�k��m�u1<���K�A�Nh�A��g���֖��y�Xe����Y����u<�k��pv�n�pm��:�^1b���m�����`��4>�Z��ӯ��s�7`}�{l&�RϢ��f�8=��<�/7n�ؾ\���P�m��^�7OM�8�2D�C+�t�*����Y9{nqٛoc���4�u����4��7l3�qŷa��4���6(v��:��Sk[�K�9��ۣ��k��'��r痷ۋ�=�s�x��TQ7\�v[8֔�c��Zn;`�c���mЃ���5�Z��vN��X�ŵƥ�y��Ό'GA����K9��Gck�+nw�Wv�Z,[�L��s�aU��)�)U��������rܓ�u�<pxۏ�Kv���%q��/Vg������sh�q��s�q���������U⹷[ms�<�n2�i;y�o8�x|l&Ö^�uu�_}7"�أf��5k�q�vݹ�6琗n�9�n�n8�:p�퍣��F�۔�ή�c�̠��۝�ó�h�c�^p'��^u�$��-�pr<��!��Y8�up�5m�\��6�9�b�:\YѺwe����#n��ҹ�\�G%֦�k;>��%;9v���X.�N��A��lힲf�cny;-�mǡ�N�'[<%l��j�L�۝���t�k�l��h��h�-�.��v���;q��n����;lꍈ'�Ӹ{�"\ѣZ�,ܩ�۬uz���m�m[�|]\���;�M�v�C�`y�o>M�%/;s�4^�
�u�Kv�� ���6��xv��]٭�]�����$n�l�����A��-9����=��\\�z�-���t^?�/?z�'=f-s��+nC�����/4\^�.����:0�:��P�y�\H?��*�A��{�i��\�i0�{���e��ѣi3���宇�L�=>l����ι��WB��+�����}a��H�Uq|��N��s�1�,���p�o�v-�&�u�K{�j>��ҩ�hk��׼�f�ʽ��M�㳥ֲ&���i��"{Gr�^\/,N]}��,�{����i�{vo]��o*�'��Uc;X��*m�7z��I��4�ma)��G{r��j��t<�v���2_�����Jw+�R�T�{٩�'Z}�ꋺ'�X��}�r��#��]umxE�M[X�@dB�����y�X������<0[�����v�Ln�:$����Q�v�i��+��%׫/9ؔ�9���d�>���J�ʞ}w�V{>ȷ�si�m�E�����)u,��O|sK8��f@,�ƶ���`��x;��w�1ڑ�#�1������֫t��-��z��N|����u(;#��@v1�7H��5���^�N�&���7�����.�#���(��P)Ϫ�r�BJ{z�x`�<0	���&1�@�1�rΣ��R�������)��5�ܩ+��uh �`�g�o��[E���?N���R'*#m��L�==Ϭ��Y�r���ιB�74?.�4J���g��U���z|�߄v�?+�>�X���5~!���a&�eZ�;�z�������R�JG�u�wC�\�ް�m��k��=CzQ���U�Q�dχ�FF���M:������wW�I#���������5�r�ZWA�����S,�E�ZN�I0s�h�X�/2�T��]�26O�����ʧ�E	u�w��Yr��+�υ�h�X۩�
 �rn�{�?DW�sO�ͮo�{Nlz�6z�&xW�!e�a��Y��8y��5*%o������ȤV�-%�x��L���o��-��'�yTH��ǞĽ��Sۜ�H6$�_=X��e[X6HVև�C3���JI-xm8hY�~
3�$��,xu�� b��+��n�19\[�G�e�e�锻����{ـ�Ka�@58��;��o����<oϽ���z�o��v[����v?<�_&�M`o�|��;�����$5�s�N�4�n�ox��Y��(�!�͙'��wc�[��t�/�M�$7D�Z�a�;��Һ��>�!��t���b\vc��~#�s4yy�(|I ��OVʧ��8�u]F	�F��Fճ�X�z�-'io[��/Y���ۮN�T.=p�hPt���-��=s��Ĩ�{��mֺi�ۚ�i�1G���'�73�$ �D�ަq#M&�����H'��^�x��}R��<��)��r.��֨��˭�Kǐ���y�a��=�K7�7ۓH×.�c��y�Q~��we{�u��(aso����_y�L���:p�=�q<uw:�5ך`^���[�+�(�[T�n�^r�ͫ��ی�"*	�����ŏV��xN��Of�ȍ������c��v[���Nk*���*���}c7(J�xiV��,��q	HZ���5�z!���'�kf<y���rdG{X���gW��G�+DV��9s�6�ťϾ_	�}N�e�%^1����=yʻ�dQb����9�6���֪<{R����G#b�ped����H�.E�t�kn�9y���;<luQGoZ��1mJ��0WͰZ-&FVkO�;�d���w�zհ9��:�z{�:]�7յy$�<RB^.W��t��{/�Ȥ�|�N�6����6bݾ�oS�#g���U������W��];��}>������t�h�U�X�碿Pi��'I���/.���2�8���P���P�/����Rrs�%t�{2�R��>
�"A�da"�'o��̳����^p��Ps�1�<���|<���X���tҮ����YJ�<��v��!����C�D�?6�Mw.��>}�,����Y���g5�������0Q"G[���Q���D�Ѣ�뽬��r�^�j�^v�֓z� */8ث�K0hw��3�	�+L+4��z�'�+��}x�K��ٔ�����yl��y�����?	NͫX.�ݗ�l�=z���N��ּQ���^ظ�q�zyLa�Iô�1�96(y��Hm��I��[�e��C�N+�*��r���<�M��.u��vlpV���6�����/n��<)Y�v�$`Skd�Ŕq�z٤�`v��Gly�tৃ,��q�-ػ`�e��Dt����{<5q�b�:����~�Ӂۉ�m�<�u���=����8 �ƺ5���O!�����/����"�YT�'�nߕ�'�ŷ���;�_ ��d﷦��>U|���z)�MMڶ�J�^���@��[n���9��g�yy���e�"3p��Gf�0_G��)�	i-�6�{8�$#�;�Nѹd)s"�#���1fO�R�r��\��]*�e{�:�p�;k�����yp�g�XP߁H	�~-���Y�:��05���ߪ7�Q�ٚ��4|2�`<�;��,�u��R�W,�;�~unJ3���t�'�>J�!�.胅05�|��̝XWS��W�z�z�::�ǒ�ym�v�e1�˞w۳�땢��Si�3�HJM2�!���U8��`�A�v��$�8�8[�W��jŒ�MS	7H���n�@$��8��,�V'���ZK׉��lKcjX�����"9~fy�\���k��X�6�@be�D��2��}Ȧ}����[��Ƃ2e�0p�km<qA���.���\�tz�k����ma��ov�B��ȍ�G�۵�X8SR��7��e':����1����\���ݛy��{����L�r�X{�7L��f-n��+����S�L�A6'�;�;�+o��f�C�3����*VP<��7�=������}�7R�*��,bA�oϭ�Pѯ(�8%}�gaH>�(��A�����#���9>u�1mm�s��g�
	m�a4�C�<���ۮw`�c�<|�S�}݆݅�b�����.�&�RI���toyS������6������jf��dik���M�������.���ң���ʙ)�h�]��)%l�vݛksp��=�N���Z��od�v�[�q����<3��jKd%�����z8<���{#��( ��{�}8g�M7B��V�[�}u�hB.��[GϘ�m�i5�7�g��i	�-�#W�~(:}��w��,�s��gұ�����BN>.��:1ڛ�f��w���{^uu���\V�����r�U�Q�)h�<> ���IK}[v��������R-5����v�Ք��Z����s�����VPdrIX�����P�t|�9��{)+֦�[����ASEcb��2۰(lmh��g��t�vL�vC��k����0�۾�B-���@�SW�*]5yf�y�˺�h`i�)����_=�Y���=�ї�������[�d!,���k��|��r1�߸|�8BzD�,��������ر�Nv}��ۜ�@��+lk��$w�Ҳ=i����i6l�ޙ���W��+��S-P�]�t���P�
LE�y��V���Ϫ�nrb�ٛñ�m��7c1�4�a S�t�u�iReZ�Co����/&I����|�FV�_=� ��[�g	�f�e�hּ�N�f�M�-���Xh�.���/�ýC}�hةJB��r�Dɺ��]x������z{�>�ژ�<�ۦ']R���Fc BM��9��<��%���&v��E�����;�����'X}���V��{ݱ�$�N}vf:��z�e�o����uy���E��緼���*n�1I�FT�V�B����je멘A.�6���3�-X���T����H�s��]��ņ�~��ӣ��k,[�3��
�.�X�%�� \����1WP���^Q.ޒ�R��|�� PE6�Z�T�W�����0�x�=�u��.2�~_~��;���?2ܩ���3v����g#*�D~�86�ڸ�N��C_��Bh��h6};�Tr��.�M���ܓ"�N�&��Pb-R�@@�D�{�JO���m&�;E��m��4��^�>'=������s��dw���|:��y���Mk�����]��:�h*tC,��l]��a)����ã6eYp��;.rݺKs���HKmC|�ڼ�m�]=p8��3���V+n0��t����n���p*���>�..b�����&y��oκ�R^�������%�K�]e���9OA��=Y�hQe|ӡE0
jX�ƃo{��l�w�(t[�j_T_?DE.�3���n�w�q��_����6M�i|7Fs��~��ӷa���[w�/bm��B�Rm��>:��N���s���zn�l?T��]Z�Rk��_���T)��c�]-�R��)G�eّ���+_s�6T?7�g��Ec�xj�*�!�{S�l6�^4Ew��H�1e�w8�W\�ϝ3�9om�95��!�-�	����m���jjJ��`3MۦG��틅{�qwHaQ�܈���:�I�l��h���K�wk�IǛ��c�v�4q���#����8��:u�\�l��r[�aݶGE�n��Aǻw\pOm�e��^� k���v��6rM��x:�������� �{X�o=on�۷b�r��;;�/�k�t�m=�#��nr�$m�����q\�r���L+�5�F�	��r+s�|}��y����uv�k�<0qc��r��ri��M����[����;���V��򹤮�����Q������ȧ�A��O��N��ó�L~L�ҍyK�S��}�f�dZ�K�)��4��z���Q�4:{gKn��@����[9�=λ��Hz&}()�M��5,��WڦLH�����}���6fY�;Eh�Bi��l�Mm�'�NX�3�slE�G���wl���z�*��۰v_�z�x|)��\��ۏv�~�B��fm%���8�(���~k5g�A]��S&m-ͺ�QӴ @��Υ+(^������ܦ��� ��E*L_������s�H�����n�*�"�	�q�wѭ�������-Q|��QVQ� >�%.)T�k��@A��\�?{�c1���
�e1D\��ꪥ�3�D|{�����;�n�m�c���7kt]E��������c�>��v.q[�".u]�^��S5%W�Qq��q�+#��������7�HS�_'<^I�_g��������Ox�[=Qy�5���AmsmY[��D-��KϢ.]�=z����|-��~�~9�C��RZ�	]���q��
&mbƨ>g��<��k�E���L`%��x��+2"�<k[��wv�p��4}I��g���\LM�!K'|�J����B��S}�6(��SؕA���	��OƘfޏ���U5�r�uPkT�ni�f��j{����J��s,|�}ڻ�^�2��?>��)2��T:�v�p�l�a����k8:b���-�m��p�jRQ�$��.4��H(_f�s�1CYwY�2����r���o��=ӫ��D��'rR��ݫ˅����l��8��w��<��_E���PѬ���mD��}S�U�l��ff"�IQSSa�K_�R5���-au~ش��f!��`K��T�#�Ad�ߦɬ�ȭ�z�{)�U�b�rQY������ׯ�Pי/�u��c祐�ur��{q�y
)$Ri���U��d�Ki{<�m�݋�Xx�1��w=t{��UX8�Ae��p%/����T��k�=eDy�����K�wkZ�,a]{��T�Ბ�Q�̱vGe2�]�v�|�t�t�>�t#���`��Ӷ,˭�[p�nܵ�B�V��P�8������X�y4�֕{�T�؞B9�WKKl{��O�q��:	�6s��m&�T�vl9��YU0���W7~�^���w ��)h�S>��Z\a����'��u�4��v�~�yuH�ӑ��ZƇ���8�n��Jo��XÍ"YƵ��T�]���)g}xь
F;�w{w�5D>z*.yeU���ܭ��k-���f�m���i�/7���1ϥ��"��F/����F����=H����żtt, ţeT)�Io�ݺ6n�
�r�� ٮ{]k��E�B�"�et�0�%V�^����7�JX*�I���*�y�#ڄ��J����D�kFf+ �웡.���^��	{��u}����A�����Ki��	ZXU�
T \��j�>F�d-�w&�o9 ���n��)�rj#���:.���bzI9:�g�PMgC^�n����&�^�m�	[�DfV���A����-��Պ��leu�]�!vw�;�wLό��`��k�⋕>;�j̥��j�1�jc7Z3ھez�h+)l
��&��\���Eb�	�b\g���zgX����^�e�r��s�S���JW`�J�H���n��C׽}������3�8b�d�z1Mf�g�6��Zɮ��ǃn,�r���Kk&��+33���r{+/Z�� \�l0:<�Sjx��a_��P-��ỏy�X�1^X�B0�]J��yZ�]�/�R���;EK����xoR��x�6����*�<�N�b�e�p����� ]�]J�m(5-A�N�y�*j&GY�n��t;�m������/����$`�_f�o<}�rҝ�0�&Y���E��)A�ڪ�i*�=I�3���|z�j��ū�)��$�ǣ>�0W;̱�[�*�V\�.�m�\�����2�O<ZU˧��uE�KlNW��96w�Î^{^q�����[���Ѭb��pOb���<��F�Xu��.���T�4�}/Ʒ���,�J�=�f��Z_4��ZW��}�r�E{}<��!�į=|�cICE5�b��T�-����X��)�bV��䥌X�O���i_\ѭ/0���{oܣ}���#Ȇ�;���x`��u��֊k�j�!�o��#�qH�㕅�И��K�-����,i�bC`d�O��U�́s��lJ�J��}�t�K��ȴ.�0%��L	aU��vy鴱�i�4���ce�(`\v���;i.�`�iG2@���kc��s��a�rI�*n&N�k�>ϳF�>�[�㱞gY-:�n��EY/W6�D�m�m,���@����^��v��$��!�4u���b�b5��k`�b]d�u���ʹ��Z�S{lJ�9{=�[����u��p`�>�%LY���i�ͫ�,6e4��!�
i����h��r�*�]BvZ4���V@���M�=��M��@k+<�^=��oĽP�1,vҦ��sq��0)�o��ր�WqĠ��o=X(��D5-#v�\b;���Ģ��sò�N�5�`������{��Ԣ�L�q1U**f�$�0���,Zĥ�+����T����q���T�t�1�� �
��:�bIcF����0T�KF�i{s:� � �-k@��u���ah)���M�KAlH���!��G|��:*�[��ꦧ�\�H�#+ku�ٝB8�a͜�ؑ���a-
X��y�`s<`KAM���
_�`�]Ֆ���q����9�AX]r)�Nm�_<�V�G���{^�Y�n�c!�[�v�	b1��:��Lڻ;�-��L���0��B���M�����x�_k�h;9(xЌbr�]�kHkZ[W˾��(�c-�и$kA���{
hQ�}�[��kM�Ĉ�(b�M#���G����J�RӮ�$����(h�H�2�%��Z8�V@.4��ܸ��ؗX��EW�f�T��u��%��CB#'�3��}��}��a��HvՇ�^ٵٓ����9����+r�dt\���rv��F���}
�����ww��׳=@�E�d����Z1y�,
b;>}}�4)pŬiŻ<��^���8�K�@�6"�r!��ޛB�w��̺��f�-4.���
h-���%��#{����@KZ����%M.z�b�H6�=Ӓ�U��2a���E��w.B�Y��\k�	0a���ia^�K{ü�Ci�؃Z��s<�Y%�rS`�1
�]Ǟ�����ZH� �CI�{�`��H8���q/g��w���m%�!�-/�5�����O��.2Ѣ��� ��֑��:`[[	�I�[�FG�괗Fj�KT�9)���!�y�`_b5�nN��JV��
h^�����xX
��W~�͋Z3!`��`6��J��Vv-xhZ�|v�ьE�й��m���:!�sU:�q�1��
}����<��J�9�yؑ�6 )� �����[�6a"o���I����"�	�H�"�� .�[6 �
6����ؓ��]u󷧼ξ�5��wf�_^�0C`�iH�S)�I���O��;#���=q�I���֒���הּbZ�sn�u�Z�l8ĺ�m����yî��~� �w� �~i�D4�7��Ew�6�:ì]i)e2w� 6+}f4�}��al�����b	`�ikAN�5��Iz�����_�wrW���VC�؊>��~�����a�t����VoL0��n�0��g>v�����DHF��هs�������ͽq��ku[�i�^��5�ɥ�e4Mv��<��/LpX79�1�Tʑk;�m�.�k��
9�WY�y�GChӷS��X_��Sݾ�ܦ��KGLk9�)ݻ���[,�v�	�y���7Zv<,��{�us�I�]����&u�%�68z�\���v���WZ��m��,���9|�=��h�v�������E��ș{%/c�
��y��)�\�;�E�=p��.R��qt��W.:j`K	iN���.�f����ف/��"���
b{��ϻ,k �0�SH��s��3��,f� )�0�ISS �k�6�����Oo9�g������M�)��9
؊hڿib���X'���M�v�c�Q���kqW�G�C�v�CK^�V�k��-kG�nz�6#Z=��{�n9���MdB5��o`��b�\�O^�:�k�[;R��w>���3Z��&�Z�m,`�g�øBZн=޳��wR1��B\i-��z[�햵l����+��q����RìZW���E�w�;J��ˬ%
��u�Ay	r�G}޼H�lD4w��g/��`�g�]iM�dؖ4�3�T��r��Q^�M��{���[Aځ)hD�֚�(�)�:���v�Mq��0|=������z%�%�Ҋ鉶��aֵ������5�r}�,؋r�r ̀R��^��M�j��(hP�V�p۸�����1�\s݋
�F0]�E���j�M
�^x#��Ad�*�f�
����[D�V@�b�G3�ኚF0�BTձC-��Z5����o��#���{��d�LR�7�IdCiᒉj���Zհ�����{��h����
YM
XW2R��=����_�L'�����g�k'=W��y�u����=�W\n�ۥ���{� 4b�v�X�mY��=��6q4u#�Xs����Ʉ�f5���؎>3���[ڃS-��d����5�L!�D2ؓu��=���;������}1>-���6@ư�{y�0����YlF0!�H���*j�sY��L<����*j�p>4kE1K7 �s��>��>�z ���1
9���j�|�$�����\�Ei�c�nf��܄��;�}��m[���3�;k�7f9<3��v��0W�A=���{��v���+h�BT9`e_�mC�c%���t�K,m�]�;��ص�8�+*z�/v���/+���y�we,�I�=��Z�v�`���zK�J�cCCֵ|�i6SA-'�睋%��qۆ�1K��F���G ����=�_"�N��2�ʾ�����d{�r�q��[R[���Msޛ9�Y6�@���K�Q�o���8�8�'e5���zO��k�{ϭ��r����׬�&�;}�A�21��GZ�"�)����؍h��D��:fc�SW���LB�H���h˄��g_�'�3�BX�7�,%��ٶ���V�)�x	m���J�Z�L��nzR֌���p5�̠��N`d���{\��k��uy�`kD5����\��z�ذ��4�xT����갋��/ҕ1G�Z\z\��ӹ��jV���G� PKd�#u����s n���u^˷:�*V]	+����Cb�L�w������+�)����[p��KG��w	]Bw�6��Q�[U�E� � Ư3�����x��I��b������H1�A}No�ۘ��-u�����֫J?����	f�S�%������Y�)a>��f��jK��ܹ�k_�\����;W)Qw�Q�̛Fu�PS=��i���3����X�5��h�<���KH����\s�a������of��^iKK毗�qz�Ӭ�,���Z]^��S��1\B:�3�U;�����A�5���5�`�Ny؉��0#����gnX�ư����+PS��hU�I�
_v%ƀƣ+�&y�W��c�ҵuޗHv��6d���[0�8!��j��q��HL3Q����z�Wv���?X�Hs"�[k�]��սI�,׉�wqV޵�]�������
�;M��4�]e3���~%�����w��1�A��B����`��zf�G�u(9�E�Ǐ����;�[�s�=�;~�.�b��}^�k�#�̭��r$���E8���@Q�ǭ}qPSb�z�ڦ�%�jɶ�mS��>�w�U��Xh똅{2�/�2*{�Z�D��2Z��iG;�y�Y�֭��|�7Ox��~d,����t�/n��n�d'v�p<��/
����ܚ
9պ6'�l�Ϋ.���\3��=zKH�l%�g������USMWa]��l���n�n�R�9}q�W��c'2}���{��mñe5��+�s�����8�j��y~�Ŏ����'����4��pzCvhi/���r���]k��pg�h�	�I��>*bྐU��oa�W_,�y��W���b�Ej���}�TX����=G�X�#�i
��2�1K$��7ER��**&�k�Z�:�t��U��d�o ڄ������1��8���*y;�:���3��g�����Q�z�?dJ�isqcH_}��^�9$�^�K&���O�`�v����+�vv�}�8PK��wO"�0KT�i�9�������M��jd!w}6u�D��U��<dC�n��=���7\����ЕZ��:t�JZ�ף
f�iz�Of������%2�L�h�-�a1���s!����e*1������ۆe�|6%���f��B,2�c�u4��[
s�U�û�#�n]6�k?U&yp~�wYB���vH�د�0��h�mzl�ak(��)|�{2�rT^X��P���Ɩk�>a��DSg}߬� <�!�kj��+�磳;�c�F'���l��FvL6�y^�yƷiո(�q�S�KR��>_�Sa�v`���J��(��Ƶ�9b���+���W��<�ɋ�[2^���l.�J�t�C���y:(���8��I�Z��b���-��W�8+��M��ͨ+�E�̘���%�ggZ�}�/�7�R�������y��'/۹��ކ9�����7S]������v�O��0�C�os]�>�v�%���cU�>{ܲ��n��ቂ���=�_�)��:���1��R�mUnѫH�#�(pʔ��!3L�Zu>z1Q����VٺM���nE�����C5��z��ȶS3�+0Wm��n�ӕz䆒��BR[�?XU�tp��GF���%�nQ,�R��$o�Z+n��M�>�E��~b�~]�;OEV;�wm^�i
p½Ɋﴖw��Xˎ98�d�"�'S_w=ղN.N7.{k̶G�/��=G����K2�yY�"6�/��W����4g��x�h�.��;K��aUa��ܭX3Jʺ����^�t
n�����mg���uxY>����t6xێrS�A���u�v��'V����*LZ�۲���m�N7v�mwVJ���s���˛�s����c�����칝9애��v��q�k��Z�ݩ��[�cf7[3\�8�g���Ȟs]�檹�ST�V�8xAN�� ��4�E�8�5��m���c(ksd�ۀ�Y�]ku������g�y���^"B��1k�[:d�>�mv8�m��]��<��W+�<�E����s��c�t��v��l::)��u�-G���������:�ٜ�(�m��¦3�n�����Ý����*'��58���D�0Lwo%�`��\��~�=��wN��yh![)X3E�8<,_���k�vv��ޞ5�uY�쫰3
��kR$ ?=��>B�@� �{�x�v�:��а����`��e�[�$�i��t����ߦ5��ɸ��=�>7����������eM4r�z�^��,�0�t�\�����E�B�@�B�k��2��SQQTY�m^�2�+���uX�	2��t���^�e
�g��R�\ҫ[��ob��]���'
hQ�n�۵j��vNT��Wg�4R_ �n�#�Z��X��R��¶��^�c��Y��4���*�S졓�X���M��D)��Ù�x�j�y>��+�2�}s��z���Xs�+�¼���Ж|s�s����ɗ��Nʜ�Q?�j4V�Ie���R�xZ�n�����C<Hl�4Rm������eУFE���f�f�L,�=7���|�y�x+��p���u��<UW��K�|	�H�A,�}�L|�[���;{jV`���jV�'�y�eqI��d�S+��7bY���M�ɩ�	jYN"�]����340sjg��Z㧐�����S�R��7[f�^�Mg2:��Eht�r�׻=��V�H~ٹHQ�!���
��w9]@K�X�	��[q���{��W��hX�ګ7T�d]�+�a%�����ػ����W���o�Q[���~�8�^���u9! l��I�-��+ �Óv�ώ��3���)������}|�ڟ_8���y���A��V�%���.j�+��ۭ���������ʋa����W��\!w>R�EX�)�EG��^rv=fT��H�{9��@>�Nȑ�b�ה����>��n{3ϝ�|�Z�"j9k�Z��x�<��q��/����8;����Rv�F&�{b���H}�ǗVFGF��<������%������;��.���D]���}+'V��/;��9xQb�!
Y�w|��abi��*�c�v{Pe.9W3J�沲�1Xˆh%��,v�n�����X!��=���^u��x��g81���N�`��<H`,����a��&r���YY����G���B�k��Q��Q��O=o,t�m�����9;�c&�u]�`1f��w����5-瑢��r�GhS�Y�T���Um����Uk�j�NېwM����+M�3��Y��^T��̚�'y��&E�jV�`�j�K�c�P��훮�E|]�8g�ςG!X�"Rj�������`T�������~Ua;��[{�T>�U�.V��9�?�/�Eϛ]ӕ]�������a���s�D�N[�ޣ{����$�M�����(����A��,��,��}U��.V�r�Pb�Pt��c��,�, �\vݮή���F�5�^փ�U/�N�hF�*'ܹ�}\���ڂ���Qa�>s6X�ŝ梸�^>�WY�(�~0���e��ZJ!-�୸�H\ ����8�Mܞn,�ah}�+�-_yP
�X0!��g�;��������Yu;ݪ�L�]�|����Lm��x��Ѯuo�=�Ȥ��C�����������ٕ�:�s^SYw8��\�R��Qgy�v�R���{~䘢��wu���G��Ԟ�(�l��+�PT��]��fI\{���Yu�Q	-cy�꘣S��={���S�^흀¥�>�2۽� �L���-��Wk���4�T��b���55�f:�I�����i��OA͎�RjVUҮz�IZ�T�����Q���Hw����l)j� �w���.*.���� U�2x�+�?lw�n�u'7�n?��R� i�������V�y��7}H�{��V�%AO�*����!���.nã�Iԛ6K�c��#�m�N�v.��vݚ*�GӭlS���p�n�V�F\��Y��1Q�8�"�.�Ip���o�[�� mF}=�1��Pye��o���'<���H������.�z��W�f+��W�C���!#����l|s�00�:���i*~�R� (����}�<]1 �]krM�?���}��K'3Nr���v�1:d�bƻuLgb��f�+�y�v�2�g�������[B�B)yý�mOK���c=��2���$ҪZ|��6��峳(%
�*O�;�Xܬ���䛔�!XU ���m�v�˦0R���I��Q:��
k�s+�l�Gb�"ȭ;�K>�����2�f`�$��� �$���I	/�HI@ I!%��I	/�$��� �$�����_�$����@�BK��_�$��� I!% �$�� @�BK�	$$�p@�BK�	$$�� I!%���_� I!%�@�BK����)��_��|�,�8(���1�0��l P4}t�N�E4���@mE���	
4P   �-�@��::  ��@�� P�m� :           �                    �  >�       l� /�}�m>���E�[��ex�wm���Ռ��,�� ��V�m���M,��t��{�{ٴ�+o3v�,p4�<y�Q�ef�eރ� t��r��,�f�L�s� �z�,�����m��=�])�o-\մ�m˻m���{� ���k7���حelq܊rٶqΝ���˻Fi�Q"��  @    {�i�i�;ǃL�����mm.\�.i��[m���e�Ӯl�r
)��vN�,�qk���lswh�l�� k�I6۝�Xm��{�s�� � �h7y���[`��t;+[j� ���lV������]2�m�8��٣Y�ݥ�ٶ�� �NU���:US�{''l��k�����������lȊH HP=�        ܽ�+G7(s[�:�˕�Tir�+e��oy�iY�� �+��nv�m�m�׼ǽ���k�˵b�nn����\ �m,i�=��7f�o,�P��T6oy��V��y�z�,S�q�Ͳ��u��4�gs �c���iX��w^��� ���6�w+�ZͶu��U�z^gU�lƳ��mhm��R��FW�        i��f�;�6���ݬ�ŭ�a�-�W����ن�� ݲ�Mk��lMmf�]��ٹܻJ�L�y�򵦬e� ޢ�[S�y�=��ݬ�
 
 �l]wi^*�w��T�RR� ���Y9�㛰�H����Ayd��w���/N�;�)dͲ�e��z ��T'Xl��ӳ�r�J^{�h3ɻ�7�rP��w3yΝeD�J h� xt    �   3�M[dU�Ή�׳[5�W�Ϊ���Rtǝ�J(4����iD��� s��{jF�]կ; hx���և��GM4oMُ;��٢٧�� 87��PִngN�� v�P� Gx�@ � :    o��2�bM�	� �t�=��9��,��"�j�&�۶�Ε*]k��^]ն�P����S��-�ҧ9���(���==7c͝�]KK˻K+k�S� )J�  ��"R� �� ���6�D� �A�~5 R�@ تT$h�@��$ʕ   y���^�m����zZ��so�~�]�{��{ݸ�}��~����w퓵����(C�km~aB�%�P��P��P�Q��ǏO�����}s��̬�qe#��~�7��L+�,X`(�3)��T�oU5`9�+>Pm Z�㭙�ڐ�7�Dd2�`�D�tFL&�M��1gE`YU{�� �+
MX\�۩��9��-���)����H�H[�K�����6�br��&l�vڽC�d�����zPǭ��j�%Q�\�!��u�.�PO^�V�T\�d��m�l�Ȓ&���o7V~fZ���&-0LjGSp^�_����mh��t�5�\�N:I���k"���*��m�L��(0H��n���/c�Q�����y�eő��['!����
ܤ]0�֬�V�.�;s&�w����)Ve �����j�i5h�hn�u��ܲ�*�I���n!����0�A|����(f�ZUj�̛2�Fn�$k/tu��T��G�m1�����V�`p��4b�򰛻m+��6�Yun�7�[�)��0(	+33]����v�������iWx�:Of�\�����)��k!���O�8R3Eɉ]�����ق��͇��c���"jk ��0f��4�r�MP��N�F�
.���f��`��x���si�݌
�	�c�YOpfA�T��F_�=D�!qJ�.��4���K�H%����DvJ�v��ܴbi\0�m���R�f8��Gt��=.Ӣ��@a�5���SIh`�36��,��Yn��3����h�-طx ���j�ߊ&,)ٺ8"��L�"VSUNl�������o�kF=�V���Mk�RhJ�&Q�w
ڳC�!x��2ˡm�e$	��3jR͍ol||��I��V���Ѯ?�2������4�������d� �Ͱ�w_u,�;nٹaų]�I&v�%���82�Ȣ{e���n�Z������[4G0ۑ��ko�rɊ��7��I�х%�1@$��!ܤ��3�JNdz�@��(B-�Y{
u^7�k7�T퓲����t��Z�eH��
$֧�Eھ{Ƴ�j[>
O6_��t��qj����8v��D^�Ƕ��1�w c��
�nM��j�M��m����,Z�z�ӈ�A&�ZI��C�E��X0,�jf�7Z��)]۬6^��  W���r:��򶋌f�{�O�Qd��P'L�"���7�"��IG�]����i�ҰZ{�B�d��Wt�(	f���B
7i[���VIRh�26�i�˚�i�0TU��F�4�k����{�ost�zwv��CP
�&��U�����ޝW>�i�'�ڔW�rdՈ�ԩnY�X�7ro�Rl�s`�n9!�9L5	UP�Nfi\�Y��i(��J0,���8[�&G49IB`��̵����;7[���7�����2yuk�x�ٸ�!��w��h�*���s.��ZZ�SC˺��X� 䖈d�w�f&Աu�A�N�sY^nl;��S8�-6�*�͠�T��ʌ`��Iʉ�00�×.`5I��(�@��Jn�b����Yc$�,3�H�&n�W�m^�z���cRG!
�3*���.i��D�r"�R�����w-d" �rT�~���8��l8~�F��)���� � ��%�f�c!!j�#�d��v�0E-en��n��6Ա�4я4F��;�"JzNf8%,��	H-ߗҜw��7��*���7��\t."��;(#�V��"���G������-�*A����Kqmf��O�q��4��Y�Gͧ���sB���K8 �c�W9�l��Ǩ�2��ԚZKf���2n�ȃi᧸�og٧�0;-�e�v���M�-��{e;%��9^'$d�T2�����-�V����n��{�E�d�(^�¨9�dH�U�1ԥ�[Qh�Dm��4��k�@QP�IV=�Q����sS~ɩy�Z��w
���*�$�m���*�{@Ȧ���5��(846�$6 NfɃ%h����e�;k',����Й���: {75�:l��g,Ud�MFB�FX�p|�i�'Ƣ�E�������]K��Z蔮�DIV	�OmU�ɒ�?�#J�;Z��4��)�*D�PSvv���l�lB�^��d�ջ�FmU�2��4��R�J�a�l3L}���\Zͥ�;��I�PL��E�ߌz���MI֧�6�-�E�Jӷt.f dY�.%n���2�t`�+4Ʃ��@���(��j`�M�aq��#zb!֙�J��on� Ԓ<˸C� ݬ�X�&�S{�Z�4,��
M8FtҼ�2�-��昱�!����k�l��b��Œ"��%����W�Qx,��i��6��͐���U��}�����	��X�IYj}7���P���FeO�7C0�m�U�w`n��F�ka:q3WBRd�R^� ��vd8#w@��3or:#�j�v��`�*˴bI��	��1�&�P��Ʀf��̨˴)�չj��J�M6^�L�)庄���F�R͟̩yAa�}1�T3b�a�f�*�įs`R�㽆�bn`�)RV����A%LeL��JQ��kwt6յ���^;^:-�l�>����� W<����0�7q,s�q�N�h��ۡ���.M���Se�2'��@�xĬ�`S���#�칅�/p�[��3Śq�7�2�+0ss6�@��ٺH�fn��&`q�C%�K�$նwF�U�C2d2��G��b���^BeY�TE;7�m�!�*,�Zi����Z,�[�v�o��l��x�v|�-?�@�m�b���rdB7�L��q93S(;�AޕI�·c�M`����	�|��f�nl*������˖�P8R%�b��q�75��m3��U��ۃ*�w+s,)j�w[6�+���ƭ�fĹ!`��FK�F�B�)D��R�6�[mfU�u�e��I�M�Wsp��nź�T?$�»82�:ܶ�ٛ��8�1e͙	��n��6�pӽU⛹��n����wKf͡��n�1f�T�F+
[o2}�WX&��bE�6m�`d��Q�s�FuD0�J���Ua��U	�	�R�8h�P��g5�N�ihwyc7QU�f����7 ۤ���t��cÃ
��Y
Ç�W�E�6��-�ˢk7S���`=��؞����f�h�,�b8���Zc�venQN�׷�P�nX����L��`[9�'�#z7&�zaoBG0b:	���哊�G��͝�v���(s^X7����FG��"�"�1�\�1	�d�(�;�5-�nZ8i˺ͺo-��G�Խ�ű�̙�݁�K`F��� b�r��9����h<�"��YٍQ��EB���F=˛�̆*(S0�F�d�$g&Td�`ef��Mc�0-�:D�f�&�ځYD��GV�5W6Z�K*�o7fE�
D�i�x�jט-eDE�>P�0b`�\L�!Z��Ù���P�!Cui���0V��Zn�]-n��L����m���0!J�n@7N�%��Iyf(cXib�$^m��J��!׹�qh��p;1JB/K�B[s�Fd��C5��ǸX3^�W��`�u�/&^�Rwp�f�����XOd��j5�e]�����Cm*Ѳ=Wg:��kǡ�j��jm�ke;[1nŕ����M%�*1�"F����ڔRW���ml�[�]��n���P���12���v2^�&�j������^4�EQ�P9�q^��9l.����=�+7��۩�P-]�Ljw���x�S��dr���[MĆ����q���d] T��D^VB���u5[�CRcL���q-�(P|2�n�Mݻ���[��aM@\����)ޅw�z��.eZU�i�{���������4t�8�8�ӗ�1Z�4^�Du(8 �e���G���լ%4Iɮ��#c*�2�������l�t�ɶ3cN�k��9�̗(������VӘѤ��j�M0^��X71х<��c�áQ#r�\��u�ر���#�kҮ�������{i���c�6�`�J�"�ۡh�.�/��hVs_I�&�{��ОF^��1����i�/��Hir<0� M�����@���9��Mr�q�y&L��X�bh=�� ʖbtn����BٛNo)���%Z���>��lM�3�VT��`z"�n�,Ptͭ� �%�&6&�X�4�ߝ��Y� �v��A�fA���,W-+*ҽ�*ɕ���Ũށ���K�n����z�M�͆d��� ֬�����KɌ��C�v�5la@"�U��N)�s*ʤ��J:�\7�cZH���U�d�#�ΊW���,�E����N�{y��ժ*���sp���f���yt�z���|X�א�P;�Lo]j��d˦�����Vc���z��G	R'6�4E����C-���n�{r;F3&�n	�b�*-��&Q&E�˷�V���^f���r�#�hfB���,�NY_h��r�itidj��G�W��҆�M��(��ypZ�`���B�f�2�͡�
��nS{R��6�G]I䳋Md��EL3U��%&.�7��>��#K뚕-ܥ�0�iJP�^U
���<����:�^[I���u��s1 Y����V��z��BDΜ�(��V��%o�Ͷ�Yyx�h�0�a3[	���ɡ�OV]�1��Ӽ���s1�
��V#�f�];�KHi�oU8�&
5�y���M��jd���)6�$��j���p�J�󘖹,];��s0�F2�3@�����h��*�

6;4)��d���G�ٚm��.�
Ȫ��;6�ܬj�+��	�����9�@��
�xVn�N,�M��k|��31���*lW�����BC����>�T�팒�o];��W���M�#���r�!CY.yd-ݛ�呺��P[hi{���)Q@��fi���f^'��	��F�P�Q����9
Ŭ[����X�ںv�#cl��1e��kh��dA�RY�.K7h�S�2�z��v�����������`��F��2+���Q2�$IN��U�`��r��k0�٬�V�Y��f��40�w�������-+%e5x��xe�WZ�����2��씖`w$cb�(��M��r]{��Ƕ�
5X���u���d�wk5^E���˶�շ�u�����1��tMc��8D�v�e�T�졛cn�n0E#0* Gb�(�63q舷�A�����sr�d��S�*�&CT�hfy��-cӗ���0*�eԭ5�&0У��2iT���hl�����iT��o0� E��TM8�<�L�kMְfiۗ��ˑ��G���@�/r�Q��YP-�ӵ5��v'[m�!էA����NL��3Uf�E�ʂ��-�����j���5&%b�JP�Yc����A��jY���c�)�MM-��+�Y���v�w�[���!�p���W�ht�����^��V�6�%�o3D��j�+%�B����ENāa�j��ړsq�Yƶz]�(�[���s*-�-e!�16e�n6=+Mo9@���k9�����V}t/[ ��^At�X�n��vG��6�E(��m�	�V���ksM��UmK!1���"/�0�d���ܗG-�ݒw
���bh`l!�.:tw1�}b�塋�tX��S(0���ok4�]�f�p�bA�&�Aķ+U�,Rr���pHnd��͇��ŵY.��˦1���6Af�ɢ��.�F�Y$R˽v�	S��y*CJ�76�Gj��"���O���f;��L���&;�uy�
�06\IY>pQ�hY����i�^��q�ۂi�G
���&�C�'"�	Y�E���DYd5gA&�r8M����ъ����֛x�h߷QT�.f*7�U���A�ncڕ��I�U.��	%n��cl��)�9�w��h�{{������%;)�XE���eݦ���4�\z����I�,�FX� �{��+f1(�pXIX¼Eʕq0�+Ō��"`4���4^���ea�������zE�Q�I4�e�vam^c�8�� �c%Z�+,��/JnMhC�
Yf��uu�^���V���L�@]�7��M�t(�̒�tm������/u�N%K0,���n���Ǌc�,ɪ�����/���ịn�j��ה��T�"�ؗb���E�U��b��ӻS.��J�I@��4��Ů��S%�XwM�$ &2&a�{ڝ`��	/�QN߅�m��]�#Z����
�F��F�Z�Cд֘v�����D�6�f-�r���1�A�^�M�f��*Y����#Miki��衮J2���IZ����������v3e��hVrJ���n̢�BˡrͲnh[1KI �� j��0]�k[92��8��wgU���pf�:z��D]7��9��
]��{��ѭCd<�*��j] o��r1&)Z����B�yq�с��a)$�5,�W�@d���!�ʰ�ܫ�h�(įCF��̂�ȵA��ts��a�V^�Z�s,^�Mї�Wp�od����H8/F�_��� *�.ˣ�#������v�V
�[����Ƶ�B^�Uv�ä�"��
�aJ�4�HZ��f�[[Um3�j�9f ���GY��>:�D�Õ��֨PR�*�U��$�����w�e�յ�婠�/�A�{@=�V���t�tѳ��s%�oLQ�H$�-��=f������k�rj�C��7T��;���#R
++(��ɀ��y9l�q��s^,�D���˹Yyʼ�Z�bX*BR�'�f�z)�d˫��jj=v��L�R,W5kMҊY�E2����e���a�-z��.�VPF����eYl��u�^�&Ho�n�1�s��幻�tekD���x팕y���wJ�xqM��YOEY��pe�Ef9��Kwڽ� F-� Gp�qfiJa�B�ʰ��7R96 "@�CQ�L�  <:��1Z�܂�(\��6N�Z�9�m�ەMn��9�0���cn7m"^��+���%�y�#-�pUv�·d�<{p�ָ�xc<�o-<�[��������1�;�ö��z#C�{q��>��W]rnH������GA����^�ٻ@�nnR�E����{�77<���x�ۡ�Vڀ�ɛq���m��{��8���gm��f�j�G+��]q�w==�������7m�'l��|s�h�ML�$�W5�2��:�L�&�q���m�T�]����'8�qk������;<n����pa 0c1�R���$��x�/գ�w�<M��BH�a���I�r���ژC����l	�\Y:�c�cQ�I�*��|��mֻw:�qƛ��Ĭ���\���X���܇x5M��^��+�6y��E�]���˸��\�:���Yc�U.��##c���;��B���g�n�6-I�����	��.v�ܹ�o\��j�*7i�oe��[F�u�}��2��.�d���{l��s�ݜ�s����h�^W���;n�����g]{g�m��ݼ���깩7��!:7���>ϑ�z,��`3�ڜ�Ghv�ڃ���x�еu�a�m����.����9�&N6ݭ���I��1�tL�,Y��d��c�۴��t�Q����<G*7�ĝmӻU��6�۞�z��:k)eGF�7k�	n"5��ې����qs�m#9m��t��7l�i�,�k���ؖ��.#��WFl��7��8�k=x��;wc��%�r�/l��.mC9��=Wm���+Óc]
���x8����a�Ѩ�C릫�����F֕�m���=�w^#K؊f�p=���;�s�b;'ŋ���x�Z��]�{��[=g[P�n���u�a�c���;�5�������[���M۝زF��ۤ�~F]�A�6�roi۴ڂ����n�m�խȝu�dLn�$=r�d���1�x��Ɨ���P�x�j��w#�Rܜv�[��;Z�Y�i'=L;V�Z�=�����;f;���6�^w�H%��
c�=�3��>���iܣ�i�'qÆ_h�Q��x���5��uns�.ڟv{<�ݭ�:ڲZ�c5ܨî�+k V����T&8ۋF$f���b�8��ˈ�C]����oH�v�������=�q{v�q�ノ����u�N��*v|��6��vcbxxwdě�MV�0��Wi+���uת�^ա�=�\H�����l���My��n����{g�tpn��X��q�3wl8�]V�mqkG[x�G���]f�_)��+��m��Z@q�n�r��Uˉ7gv�Ӎ����u����u�����j�緅�a�m��[��ׅZNoB쾞�;���<|v�\�k�.������/Z{��v㎷��]��zv���έӱ��B����q��9�5���\jֱ<�H��ϛp������>*/l����PI�1��+;�\� �M�hP���]�6.ݵ�\�ت瓞���.�7mƹ�vL�����sr!Ʈ�n�j��r��EC�60dܾM�c��b����=[�T<�knc{%{u�J�;�x���qL��]<r�˹{�:���>��n��D���6~������bS�ژ^Ҙ*�ӷ�k�F��T,�gk�^�q�b��Em�ܯ��S�v�wcg<g`<;��q�*��q�MA�;q���v��n	SFώ�q֏g2;�+���
i��d�`��ra�q�њ��,�Sc��8���ƒ�r�u��+7����s^�]l���p'ʝ`m��P�b����`�:]�k==/zmsγ��9�:x!��d��k�N���᭗Qv޷�����wk�1poV�9��(��G��]��t�-�n��=.�5�v��pb���VVgu{g�C`�WGa�� {V�L�l�玶L�x�8wd�7#d�C�[���8A�C�y�h-t�������=�wk<Z����Μ<�s�O��{vѸ4��ny=rV�2�r3�^�����6Si�P]���<��Ǌ�z�w�s�ä2�um��O������V�,q�����:�$e���m�t[�ppdܥ�X��۶�n۫�N1Y�a�+���tku�_a��}�c�l���Kv+ �@�F��cŉ��u�/U��m�n&L�Ѱ�g��}�	شݝ�����D�v�F�3�c�kn�n��]�p��xT-���8��ۊ�mWv��kpjs¦�j-�qٵjݼ�	��=�W�D�6�=�s���������LkM���	�ȯn�fm����5ƻ>Ůy����ܫ�h���>���� ������ɞt���N��c���g�.-O�vI��O�Jt]��v��^�k�y�>����;��sF�������Y����H����F܃���ۗ�G')ln��v8γۧ=A]�[�6j�]��.@�5X�M�ftj�H;d%�=���;sJ[a�^9ӸК�j.A�ڵ�ٻl>�ꛖ�=���x�$�e���k��q\;���D�J�IG����6R��xM��4��V�@E�w�3��m���g���\ JH5Y�6������e���s�ɹ�m��^�aq����`�Z�/v��u���5���g�wb1��WG��Z��o/rX0�6��k\g��v͎G[����[G;�r��u㙒(�(���l�7M���Y;S���U���Wqd�!�����m��m�c:8ܩ�VuBr���]D6���Μ��\;ۣ�k���R������5�c����;���\���0�Y�gܚ�4Q���B��X�����9��س'�m�����lQOg�����!9��ݜ]ģ"���t�\\p�ʽ* rv�I\���-�ye�viێ��n���x�Зf�,n8z�ݛs�Dx�*�Av��|�p�֣���{=A���}�umA����p}��A�_=gs�u��kI��ӳ������������z�\V��N�ŕ���s���麭��+�[%-��f���&�8�z6My�:�l���{m��-�l�vd���C1�����n:ێNqӍK/.�C�a�[>c���<��:�펜��`����� �-ӌ��n��>�\��v�@�w.�ƻRE�˕t�ٚ�7�5ٮ]��PX��P'򔬮�ke� �x<�]��<d���0�q��u�x��~����7���s=)�f�W����d9d��l���À�6�ۺrڶu���mh�
;���Y�[p��Q����;L��p����9OΫ��/� ��l����x��]=Wo�6�n��V�]ø���ۓs��KF�e��}x�]&��g�+gvn�sϵ��S����;i3 �q�a�n�y�90��"�;��^]��%<���<`F���a˥�6�d���y�5e����ɸ�=]��^�;�ᶹ�7kR��g`�����a�Z�n�p��}5�s�C��8v;-�^5�sylf=]a�W1\���CTbw[�4v�d{�|;/���;s�������K��y�P� ����w�_��:�����K��GמW��8"'���s�>�(����>x�Ѫ��f�H{��U�C���wM�n7=g��]#:�l��k����7���:�K�i�Ѷ�.��	'���9�G�Cq���:����Lm��9�E�b��#p������}[����l=���Js��k�y^ű���q��wn+�nN:���XGr��m<�>9�n'�9bfO=���ð�mi\��R��ۇ#Sz�˰=�8т1�$n%ǵ���ź�m��{nx�nM�u�\z��y�1�5͌�n��Vܝ�v�u:u����1��^�۫X�d<�8+a��i����n^���&+d���p
j��ِ��K�pv�=��S�x�u�N^�C[t����n��6�0Y��a6r�'������=n;uvyݺ7�h�p�c��7]�4��X�B�K�b�%ɶ�%!rJ���\�8�㔬d�6ln�����L\��٭���OZ,�|����F��6(��b������=��K��D�Z�Z�b��㛗���n�Ok<�֣U��;c����r��pOF,a�wK���a󻛫3��f#f�趭"��x��u(�C�\a[u�&��77��Ƈsm����=���f�[���(�۫��v���×N��kr���������[nN�2���V�J�a�����=�v�v�crݮzSu���Ѹ�d'�n��]�<�ѫ�9�<�l�J�9�M���mv�%ݻl-�v�c�8�V��	���V�ѶP��S�s�;g�����RZ5@�u�ڢ���i4^u�W>;u��m��P`�=;7'S��3�W8��2㕞cA���p����q��<�ׄ��8�ä��������%y6:��8��j\��v�Vܚ�cl���M;q�g�Eƺ0n9^��Wm�p�C����vy�U�6�Ƭ���=��u����
v�����䚎�nܛ���.�����y����zؘ��mv��xq�Sn+(E�ɶ��v���;̓��9�*�gtr�nq�/-����t6�$��/gn�T�n9�	��p\�[��Gg�Y�^�G��N�Vݜ�v��9֫:��޸� �6�>]� h�&����Bj)��6�����Asٳ���}N���m�0�,�O^���9�:���_n�Nw<;��؎�Q�ZzڻN<rWm���m��ۆ�ww��i�#��-�u˹�ғ���X��'di�v1�N�c�;dߍ���ͻ<:�&�i�<v�4�.^�ؖ�l�x���'N�4b�kI��v�v,���{r�m\ۯjb	n����^Ux���|��h�һWf�Lun�/= i�8Zȓ��)qgOcn6�p�Ԝ�\L��\J��=��[��X�q��wJ�h����0�y�j�N��N�S����;^x�ۜܯgGclr�%�>4�۶�=s�����&{a���v���<��jۜ0Gd�c��6Q��g�~�{���w��-ǮQQp��bQ��-̍�8�j]K2 5U2�� �/������Gk)�eү���N�7<$(�uF��zlVmo8;t��>ַ&yS3�F�H��;K��F�0bv�ɭ� 틝������9_�VMˣ<�dի�8㎣�==�,k;c���t������+b���.Ϡ�m<��œGn,�/�8�N�51p<ϰ>-髵�3�����8l�nM��ۮm\�:D	���l�ľ���q�\��;s"�twge��1+��6q=X���Cu����G=�[]d�].��k�d<�<��Ύ��q���9嘙l�gY��f�
���(���k:w[��-qj@���u��;%ǂ��G��{g�,��딋�;�mn�G;�ݸu�\�D�\cM��ͺ�m-Tq�r���������kZ��۱�9�.���l�[�n8cV�z�p�k�ŷm���ծq`��'[��,��!*�]��S�{&n�}sq�0d�GE�k"�W]`�-�'��u�:�NK+g��m�<a��ӷc�Rٲc�n�n[u]g�K��m�c�=.(�� �.�׎���i�̦CM�\�ʼ�֣\���y�s�n8��x9ή,�2Q�ĝ����.���ֲ�d��Vz�@���Ƕ�u�mk��7
v�%ca�ѱdݶ�"��\vu�-6��4�iu���]'d�8 ��:.�w��.7�L�m��^�oj�s<�/k��;��=x2m��S��^vu��sgsM�ɭ�m��<�t���g$9�<��^9����<f�b�;g�s���H��34����g�r�����ܙ���7��P��I�ה���Jt�6�����Vn�n��zvا�_펉��8 \6��>�<�V��m��bE�tV��]�n���s�y�CН���rݺ�Dݝ�&�qۢ�T��ŷHh��y7kI�G��l�<:����w�ح���,떻	q��9���h.g���uΡz&�s��>VSq��ezVNB�r=���}�R�~9E�I��Y�B�BH$�HJ@(��DDDD(A
�B�IBJ(P	*���E�,�H�)����:�~&t@�;n6ջvK�8�F0���"��m=��IK��g�#��$m��Z�۝�5y�����V2��s�v��#s�;[ֶK<P�yyK��}�65���`ֵ�>N���Wn�]�{Ƿ�v��k��sɇ�ZՑ��a�Fpv�gv����3�/6�����ψݵ�e{te�+}�ㄴ�cEOH]h������3*���l�c�nr;�"s���7nrw>D6��2ې<'γm[j�׶o��y�������\zm������YGR�ݛ'�i�77&��λ�A�̦)�3�����pZP�V��G,���e+ˡ=׈�ڼ�Y���I͂�Ե���s��
���{��ӬZu�����{ҏ��ݺ��88°�H LT\f��y��qU/�^_��=ph�@�B��A�$��䞨�T(An�~�Xԃ�"�y����k�$X2�9���82�r�[m�o�Xs��!��
X 6����]�+�;3���^������D�U ��YK1ο5�	멺S�d{Ju�Av�B�f����_�'��ܫgM!ur���TK��&Կ��s�����u<I��W&�n2�����N7[�8��ڐ7.�m��f�
ҵ[��,�e��O�s���d��gݚ2��f'���%f*"���Ct�y#�b��b&�X�l#�& ��3�	�k�9jnЉ�q�妐���,n�x�їٹK)�y�[ss���u�3r�,h�R��DF5d��xF��^A�1�:]OpZ�$5�L��b�'3aar&̝4��+B$@*�wE����C&.yC&�'�i�-,֦��[:���wn��}M^K��;�^��D��r\���3 �\���~�[��]nT�P�m�$�ӹ�l^��N��{U��ZB5�A1�TH�)R�̨��j&��^�9&֖w�si��V�<�ҶvR F�t���������{�H��T���B�2		d����&����ݥ�t`Ւ����"�}:VKE��f�IW����9:�X�x��;�e�=��˧���p<�l����N:���Wj�ǜ�k���/��⽹y&`�,X���B�{���M��_+��S�ɯ��0s�.ڪ�����$���ɯ8l��;�R�l�o"(ako8�n�y"DfԂ��>��q�#ӑ�`V�7T�$�dLMg�?�v����L�����nJ5�+l�v�C��:�w#w���cM��a�A)�����n���SO���\m∮!mˣ�����C��f�C)*����-��N�$��_۲�"��ݛ@A'N'#����aF!��V�H���N�ɫ��XdLK3V�7������1�=�*�8�a�X�˩�͜�A�a��w@�{�rr�~-$�V�?���'�̱��yb�U.���n]rE�U�XG^�Ckӆ5�g+f�f`U+�,���^�SL��o��v��hC��m1���D����F"����������������s�-�'��%�(�]j5s�H97��������Rq�U�ۃ/N�.�����e�:��a���ET-�Rҍ�8���xUzw�f�0ɬ����&r��]���rF%��ۗ�u-f�ɰJ��ޖ7�0���,B2��d�O9�=�-or���y՘i�7�b����.m�gВ��Ѭb5>ןW��C�
��T�@8J'T�nVs�+v7`�[y7n�ݘ�;8mw	�`�G&;v��k+v
{��<zw�T�:�A���+�2����N5�Xt^�>�kw�S���u�C��gZn�<5�7GqT�TH+桂
��K2D����//9mП�8Q�[Z���yԵ!�ʬ q\/S왪���3� �E�d�UM�^��-�%�������8�b�Oz�-���T)�h�5pu�'U���ݣ��d-i���odݧ��q���2��i����ܺ;Ů������]�A���^���o�XEɅ�U��e���8���|�і�d�e᫮�����Qځnh����g*��E5�ʼ�ӧ���^�ήU�	n���̻�GF1��mM�wۯ$�픪�KS
L7\��>'�e޸�����Ǡ�ɭۭ#8���.������z��i�sf�	�,[*���,���u�"�w{����f�Nx�R���:��'r)�>���Ģ�����͗����cG�e�3F�sw�2z]�A��J��JS[]��/H�N_�D��r8�� H��&�=��$�"��F��T+w{^;�o9')�d/}������:�6�Y��#�PK�N�3M��`'���U:H]��aO*a[�#3l]�U]g��ݸk��!)�f�����I�4��}��_�k�p-ok��sn�m:y�9�a�;m�]km�mn�^͖��q��4��.�ӃC<y��c�E�u��v�Þ8���q�睶5���d���[�ts�R7��F���%��nv:z����^�':L�Ր��A�Ǵ<��:-��8tBk������G;mq/��A��F,RC��q�M���+�����kv�H��mV�t��������\�/�\��/vv���n��!k��@���s�-qDm*qFL��\WG\����ۻ�����fD�����1����=�m�L�Gh�Uu��7鲐j�����M@n�)���}fF�-"E)�����Fd�ö�V0|Q]���4r aoH���Tˉ��qMȳ�޶>��V��梶{[��o���x�sX�b�YVq�!Fn�A���(��a��O
su�F�$�4Q��P��W��U]�Q�ZO*Y��~��m�ث��.�� �`܀�A�FR�w[
�I
$�k�*��V�����\�^�����W��Pg�u� ����W]�U�frG9��B���`əR$B�{�"�bhl�
��ɤEdVߠ�mZ&�n	�q��Q�N���7�R�җVɇY+cJ�W"�	��(�-̍����Ta�z�L�r��"�z��Q=&l�%�<��sIbZ�.�(��M�5z��A���^nU���'�Wa�{V�_�����*A�Cչ�7P���H<��-�w1R�\�e;$>�E�/��r���s�����U_�]OL�.�^���	�E�Ym��� �W�1+fԒ��Sys�n�n���đ'���YF+.*�"�UPRUe����E��w�KJ)B0㶺Ń#k��á9�T4�Pz'��7��9��,.�[A�B��3��FԵ��RQo7Bx��|哛�QֽƖk�7d�!pʗ�舟*<Vd�Q���%�v]v���?���fHʨ��Pl�Ҳ'9���L�����dme�VM)��fn�8`&�B0j�����RПJ�Ӄ���X;>�y;vz-��nm�C{Q���vvl��u�@\4�|[�ޏ]�k�m߽��ߋY�*�7�qa��.�*F;:��b�2�yjw��o�Ƅ�{�V�2.�q��쏔���P��jju�̔O4j��k5��ֱQ��Uz�C��N���[�U�,{}�i�h���Bs��|Nz5��)JUe(���y���b�T>�Ng{��D���#e�=�X�f�t�v�o=��&�:�LJӺ�x{�cŖ�VȖ���D���ن���1Οm�,t����%oa�j��fKB֨b<v=֤Κ�P��$�%&v�ݬ�*�v��FBYx�=7�<#{��Z�q��u&�oq"�� �V�n2�D9�;	�(�#�K��v�/I:\S�u�Y��v���j��ڤF7\�G����	���k��1ƽS"yT��%2�E<��"��]���b�6���r���4p�Z܆�{���kl=�{<��Ч[n:뫞�ܹ��4��<Sϯ�3����_qV�T�dB�����D��4Cz�-�5�^�˛A�;�y�+u�H䂒�����^��0m�Ɏ���:��[��1�xE�F����E�K�n����������X���$6�xq�E�F+P��kxa�J���k�N�Ӭ��l��vQ������9�ɰ�yۋ"�L옵�`�Sv+l%) 8����D^�Gw�7�I�>�d֩Q����T]z �
 1Q9��O�=Dj�,q�'ER�2$mh��A�174�8���uC�۹�f��@VՉ�Q�Y��1�;�@:ɫ)̽����]!��bp׍c�Y7� }吮�nk�*�.wsd^��F��R���ʠ]�c;)!�<�Pȭڹ�=F/W�=�R�3�C��.��[r���Uy����T�[Ā�����e��=�v:S��\6�\m��ym���E���)�Οj��}f��i-�$�H�@�W��˱��嬡m�ȲԼ�E���}rm�f�OCtN7K�$�- 2�w*N�Zh#��R�3�;5]z/%ɗ'f@�1ڊo��^�@�=3�A�[dE���H?B��O��j��u.� 8��&�.��l)cb�.���]�U�(�ڡ�V$�m!�nU�b%�2�����.�{7��s
�00����P�,	׵a�#��Em䫳����t��9�����>m�uXG ���Z�Q���Gn�T)��ABxE�{����9ش+ṕ������8�WoG���J���}�f���Mj�9�P����/$իY0A�ͽn�M��e�W��
T-lg/08���j��ѷ�v ��R��.��! *�j�ܯ	����I�������swV{!�5�n8�8���[��÷j.:\m[k�9� �m�X����Jj.��)Xѻpƶ��q�9����1]k�|������c��0��(��\Z:�	�D�QKQ��S*h��nh��X�ۉ�&r��Nk5�$e�=g��l^U:�m`u��������̸Q'r��W61�=���G��<%QŸ��ڻs�ǻ<�v�;v���s�B����o1�u�ܑ�{uڭ����gz�|�Yk#E(=��(�e�w�.�k�|͉�uVґj�>"=z��b�Jq/jf]�kfb��Re��E5�.�#�A0�je$���7nE�FHa�b�D^��q0��$I�/�r�a�������s����;�u��B�]#J��'�����q���f^�H�UT��s!#|苻��@����^6��|O7>D՜8S閎T�jV��MQ�i�Z��ņ�o����A�!ʬ%
���ǆ(��	����[>ћ�|Y��ǯ&d�����"J�c.��B-�05{�{sdi#�դM��F���|f�����a��-i�R���nD;/i��ջ��l�c �n��qO]b�q;� ���>����3�~�^��]E�]��t�s��aӹ{�\�L��6gXʧRumۇs9�c/j�6�l�+a�!bPe���U���ɫ��Qk�I��̑ló������1%�q,jDhc.��ۗX�#o�\�Ֆ[%I1�UZXlЈQ����q<��i��e�}p��5�n��驲��oJ6�*'l�هh��k I��r�:ݮ\�[�E��j(7�M�����x���L9u�ȣ���n!�F_pv��/.LZ&�l�d�D&3�fvf�\�8rY���̷ �@�
Q�z�p�y��s5lr��ңs�]�#-�x�2�ͷ�*$=��X��Y�4`���v��<&�^ٱyz���&Q	���9BimH���꭬o�&��d�:�z5m�;fnğm|f>����]�;�>=��vW^�L*v�һ�TM�iY����-$
8�-Dza�b�w)�Fs/:��"Mm�W��\{.��:DI�R Nv��f������q@���\���P}�U���m�r�<�u9+V��O/65h3ًw/�nŶ�GA�≸�i�X�r9{,�7���3tDݰO��{�҂��;wi�n�LDV�+;��x�|�u<ŏ�N���+���c�v�Ǎp�ƶ��]}b�62�+1P�"+1����\���}U=�ܘ��7��Ң��w�����[1�Ǥ\�P��MË�2���b�kZA�[L���Sټ&D�b0*�DB��-�Ӎ�T贴�č�N��&m�PY��j�H>��e�2��'8��2�Ti�;a���5m(8Sw��I�}�Xf�ht�ffW	M��ݪ���ˇ��9[bAq,f�'Q��c�Y�%ج8Ol��1�e��5cl����A}�r\O� ����p�>�.� �8�V)��.S�+7�\���%�X�e�l�qf�=�LR�w0'>�q�������1�[+�9����/�u�sk2,���@�5fV�L+<z?��-K���p�*!Ԇh��PwCG{�/.,=�xȻl,m�,;�d�ʇUEA�(��ce�V̭ɪs�}W���F��{Nx\����G�dШpB�|���{z�E�:�q�&ɖ��h7��^�ٜι�t�p:���FP�=\��6^��2���[��T��s#a\47dVl\^���jSO|`�"�ƾ����Nz�)ŗ�[sJ�0�q��1�&d�����Ӻ�Ι��I,�.Cu��)v����l������)�vg��:�gz�Uۺf�0J9�{@M�<�"�
�tEw�v�͇D4�]�����=���W�2�h�ʜ��z�����x{
�{Y���
(t0R��{&�U{{�	�8Q�Ѷ���0S�"3r|d���׸.�!qY��x�X35�i�xi�]�e���^uK�lp�y;��R�G�㸤�o��9���꼩x�4^�x�w"��I������7��눧cMӼ���X�jV�(�O0�B�t��V.c������؝�yA�h�5JE�0f ']�gefk�B�-��!���pd(����g=�f��]aL�o#L�2$���Pb�DH)����/*3�h��HCؖ�:sD�*Jw�	�s�˺ܨ�R�Bg�Yu�1��>�Eݨ;n��o1`i�ɁJ���g����Ux�7�J��yE-��G�w�u����6��t1td�&�I�^�XuIc����v{V��r0T�|�\�m�I�%��u��~�xX���:e<�z,]�ok��(��s�9N6�woS��՛#�f�niД�{35����t��(�{���Vl��.�\���.��8Ϟ�8R�|͝�.q<���M6���9fv{tSWu�`R��3��#Kn"l�lu�"
����y1��J��脮�z�#+���m�nml��Y�"rI;�F�(�룱5Xi�؊�SѸF��*}������_m$V�g��o�2��ֆFi�vH�V���ĞoC�.�X�*�^��p�o
����
i�Z�1�8AA�l�v��+���K`
�P��۵h��y7����z�M���<���( �l���YZ���[����ǌ,��i-F��S�]�AS�XE�[�J"l��%LvEPq�p�w�e�A�s[c����&��[�Е�坻On�t��L���7�N֊�Ε���j�t��F�!�����8p���L���45ܵ8e558X�D�c��n8��Y��r���\P�+��y��]M�~�m
�����&�υ�kdƁ��i�E��سv�}��G��D�yԫ2F��+x���ŃP<"وmB؊IBoRjK���=oI�V�x����kב���2�Վ���<�n=�U������ʓ��������t	&��1V��}���"L��W��>f��N�<t������N���^�2�K]#�Ќ�5ި�vIE �D$t���X|5��p|�0�>�����֠z�	(�����*Q'+�w��#YC.�h�o'o\�ih:5��iL)��pej������3dd��ں�(��W��&�
�!���̽ׄ[ᱍ�-ޓ�;T1@CdG@k��{�tή���Y��\��ra˯rY��(ζ
�)��ˡ�)�jn�;t����mHt�n9�K���s۝=z�v�uv5�]��N�`�E3�m��-�Q�Vtap���:�<{7]&��ۍ�:́��;�uE�7Ob�s��`u d�h�g8��oK��G6���<���ފuroZpel��K{6�[���na��^v��h5��	v�m����2;����o�q{Wd���)��ɷcj��k�dn%SE��������&����Q�m.aO&�m�f���w�<&�5=��a�^;�ҶO���Ι��4X�Q�GA�\�eyg�k �d6.��e!�|.���L��M�D" ��闗�S�z���̚���i͌U�/f�1ȡt:�DNT��kI�@���V^,���q���v'/��szzڶ3�p�=���c�+�&��$�0���%�f����H��3�ͺ�֑��'���d�ʩ�Qs�.��4�D_vlC#Ne�7����Uu=�Z�$`HG$�0N���n˳9RS�]s�g>[KI�]���������Ue��o]O�Uv�k�cT�1aZ��BY���1���u��X���\{�y*8��{�va��ݞՇ�fm�3ͨmj�}�+v�WYB�G��q�F��ݍ�	re���XM�(..����B�U�f�Ή�j���&x��0�,0�MI�̠��7<qSW�B��b����y��[��Ȼ�{!�����4���gVn�+�9�F;w����'��\�r�Ia��{nj���{Jn�&hVfN�X�wt�Qz���;�J�r�s)�>s�l{�b�Q�(=�!���i�@ܖ����yύA�qo]�xKu�����vi�rM���@<先}��0�Hp�"{w]d�Z�mk�/S�W���&��8�.�������e �sp�k 9������D��9c"F\_GhJ�\�3��ť�#l��RoO��!�K��`�\}�Α]��r}�&�"u]�1��m��0�D@�G�{��2\�9���z�a˙��v(Z��)���-b/�m�-�P�Y۠�gB�F��:�J�պ�R�����U����9��뻞i\C)o7-X����@{cѦ��\��QR�L�]mIF_?I�gu��A�5JX��fлQ%ʹ�,Y��#�ͳW�%-����*ж9h��+9ym?L��V�5Ӈ�j�aSx���-M���ki��Pl	R�)%��o{e��<	� �3 ю��mA��8������*��݉��l�C�H��y��{I&�xFr���PjD}���iv�J�Z.3c���.�v�5R�#�Cꫦ�!�����D�Q�ɫ9��Y�}� �yt`�xC��ya�!�u�6����Uj������1Q��9��mn9��2��"��QOɶ�/�%Aͪ�td�Cado-}�s�ɱ=�����-�Oq+�ۊ��C�s�O/v�#aT<L���*�e�:��J5B��QB��du�f��b�]�¼� ��=gkS�{x}qs�RN��$�vv^�'T��R���a���l5�x�aӯ�5<�>
��j\0�����������>�Ev�B;Ev� ��y�f%��#��0m]-����[7�;��E�N{k����c^J�G����3�E\�A�>�&a�#P{Zq���b�3��n���^͞���
��U{u�&rJ��� ���ﾜ��|��u���U�@�#fJ��Z�,nV��)��վ�d��L������Rz�*���.[9+'���i���2���ܼR�r��U��z�]�'M�*��ejb���.��|%U<XMu�o1:dQ�c�������M����-�t��Ρ8qc]�|V�S��֤����@Y�3�C�*As=�,�.|f_�Kv��tv����T@V�����8��Ug^���7��k8Ë�� H�նA8�yvݍ�c��EՆ?��o��6����Ɲnq�);qp����G*���?f�߳7��U�(����Lg��Ռo�!���@zʰ�_T�S3uw�T�\&�$U��L@Ne#�͸��?����뻮��c0�2��L��>�]s`� Q�ϳ2��Ɇk^t<�'M�<�\k�7�ܼumIo��eLm@	�b�ȸ?D&�=�ۧ����&�BjS�P��߶Z��>c�Ld䘫I�W�>ӹ��듮���_��%����{��Ow-��ވya����F�$�sjݘg�Ӽ�R��<n�%<!]��|s���7+�UߩJ�K���$���}Q4r�DDdIº�ܽ>�{�j���]8�<��7Q:$��o�"�[�H�.�����&_v��A��@�ó*T�:[+#�,7B�W	m�ǝ��V�IL]\lYV�������R�=`��S����B��t��`,B��Q@z���̹t&��i�-�6��c�6�ѳ�d2�R�ۃ���[�����cA�=��]��e�N.s�4P��[`햍On���v2'5��;���}�v9�YȦj�/by�ne���6�5��p�S�6&�}�,n���n+=��uE�;�M'���ۤ�����"�շ/90����5��dMx65��rq��҃:��ul:�ˢ��{$v����]\�s�Dn��gnە����&석�z۷�:գqBVR�['KN�ѕ�}!wtt�S�2!lm΂��q�3�̻��g���7�SZV��9�';��"��P`9�L�d��=�M���kUx� ]�u�iV'�
�fsr��#4q�+a+~&[��]N�I�-.�ަp4mD`BL�ݜ�����7�Vf��|�"Mte��I�4�8 !����������5�7�|��kܓڰ\�z*�N��vY��V�Ӵa�߬wm��FfZB"���ݛ�m�cͩ����2ۚ���g:�TDM����W��v�Rߑ���wLF�%������VL�ϻ�g����Y�oX=��g{��͜�{��O;0ְ�5#k��11�y�}��]���1Ë�c��Ԏ�f�wr)4�/ͪ�l@Z:�r E���<�%��-��J�:)�ӭ�����+d��CI��Ahң���<>=��N�l�%FZ��%�`�?kIf���a�SkU��Ir�j�o�~���F����[qk��}wŧT��Q��Z���9�^"�������Ui���eA�[̴�H�ݭ�y��ٻWJ�LE�i�/��t)�+�TY�O�]6,wBw�,��8l�^@-;�m��� �|��{�mč�I��@���m�YV5�AA��
�]���]�i���%��V�8�X%VV���QV�קU��zP����������M�
��^AJ/rV7{��j�"6�|�7)�N۞{�v�n.|���ݨ�Fلȉ}v�9��C�c�>����ӂ$-*�вҽ�ءƦ���3����d����1VSܫ.��ӐJ[���bz3͏=�y�J�R#u�ϫ�5��{���{� ���W�:�_�x��3a��<��\7�qəMJ��,/�ڱ�.L�4vv�@����P,`"FL1�'N�!K�6Z�Q89�y+�:Z�;���>nr��F�r&�Y���[�\]�n�4�P".f�$�I���M���=�u��O'\cq4w|&��^�	b/�m(����L�٣�$I��İ�͕�z^��吉в���;8�s8\�f\�C�25WZUB��t��[Q,f�tԇ8�A�a���H勃�Gp���(�Ơ˵P�j���E��R�-8�)B�x8��MQ��[��kd#" ��a�[;���+mu�|������� �Y��4e|+��&���φ��cq���sS8����z2��[��}��qOR>fH��&�vҙ^��3��W�1`p� RmsV��w�k�;cS尼 �۳��DJd�o|#~�΄7�*�X4Hv��g�a~�uiyt������[j���<�g�sθ-k� �u��zN;.ֶ��}p���ۊ;+]���=�"n�M�g.]���m����Y����ziZ�7_C�&N��������E�z�'t�6N�������J�Bk�02 ��{�S�R�Q�X�duJ͛������$���=쫭<њ��evn�}J�k�(�u�w�0[նm�´���"Y){�cV�wG_����]��S$;st��9�⋎�g��vq>�1��M��!e��%�/���^�$��
䢮�Qw|]��I��7�#�i�L|1]���V�P�Oa�/XxX7:��m%��,؏>��%���$
��T���$�'z)�n�8�����s.��P{�&�^��T[s.�KU����G���䣶�Z{/{�g�r�)%tN�Dz:Ƿ��l!<-����|1�0>��9Wݣ�3Ii@�zV�)U3A�	�`�����۽9��\k���,�@��-�NC���c�t�h�u�S�]#DC���zc;�#�N����^���v��{���h"��R֯��<��c��oRS�~�ɑ�I>�NS�DY��ݙ!�Z>B��=�dצ��=t��=p��b:pt�lr׍����ܙ��V��X�v@Pk;��.0R��ᬚ�x������!� ��gls����L�l�섾��uxm� P�˳p/n]f�\`~����M�Y<����b�=?=H�U�P-�H�g|V�x9U�+Ѝ�<+qV Bﭒ
)|����=b�*`��)�Sѥx�ފ�i�E��MA��i�)2�m��cZ�{�D5��Ͻ��k1]��C�jcj��$d����8�0��x���S�<���q��Z��7w��^��z�t gX7���֤W�1��ڷbww��s�	�;�L�\�v�L�N�(d�%��G+�v��6��CU{��VC[$�<�ѡ�D��,��g��B��	��#D�.����C`ݿ�t���$5p�����0�ӓD�b�N��j�f�	��
�#e�^��u��V��e�Q�H͌F6��E��:`T�����$�Bp����ވ0-���|�
p�AQ��]�d�f�H�s{�$�I70��e�Mٳ��"}��P�����$���ja�[��0�K�o^KTN�U�a�/�Igpփq0όm�[�aj{�m� d=Gm�����9cp<��J
ܑ����յ@���e���;�u��imȮ�Fh�����zĕbi�;��%��iNuB�oq�E؈N�>X�"C��L�1�3=����k&VӱG���N�-'7)���S33;����3��K����qޫ������ŵ5��L��R,+jK�³��r1�}ѳn�S��f3����
��T�^vE%�qXk#ܲT�R
]�_e��"�rY8�l������T���\u�ŭ��4�������&l�5��f�RKd�V�Ё���2õ4P�f�"�w�;�o�rY]X��6P��d]ēr��.G������u�Vv��f%׀�wZ[��_\�7��e��2p_�N�q�
���Vs���-lHı������壸���c-ݖ`�á�
���}P>�����<q�v��NW}�O2��v��Mڢ�R2�T!�V��H�.y2����>�����N�W�7��nNn�.D�c�WtF9������燎ݻn�ۖƲ�٢�Ƀ�[�@�m�l9����U����n�--5����g�N�/Z��2�v��ۗ���ʉ�ly��9lN_p�۶�Y=m)��1X����[;:�Eu�b-��z�R�[�%�6�b=y7,�&�V[��6��s�w<件n�ѐ�P�l0˹tZ]�,���R�3̝q�$�;l�����"����`�tv�<�6��Ԛ����qj�6{m�2>-�;]��3	�ۣ<CШ4n�^�lv܉lh�8ǘ\����o,����n���f�-��ۍQ��\�(G��n{��n5tGl�{a�x5�ss�����[�#��;&�n�ps@z����I��`͠�9��q�n!��;r=i��It�E�������&`R�\ClG��PH,��윛�ۭ�[t����ٻx�0�q�V�Sr�JVp}�ݻ_�q*����9t��3۲����ҞֺQK�;af��̺��j��Jv��峸�d��c��͹2���ںq;hD9�vλ�q��[�e\/4�RSd�U��v��ءnv�;]�0p<�S���ӝÐ�'��m�{!�§���T�=���!d�<2��`�I�N��":����n5�����h�)@sN.��mt�'l'�:v�Ñ�l�����&^[�ru�v�$V�WjDۜ����R�4�-��>�x��N�ك;o�q�}�b\��һa1�0��-�f	�Ѽظ��r\��*L��f���[����;s��g[�8�K<����c�nq �nݶ�6�0�l�=.7=�q t6��|s�\|�����A��۱�n�Ç�OI�����50Q�c�lOY1��[��Y�b��2;�͜���ln��c'��[t�]v�8�S�Q�t�i��9��0������� ��0�������n3\�f��e��<�����,(pQ�Y�0m�ۛ.�عȔ��vj2�l��L<�7m�i�����n�)���8��㨃������=Z�\\���q�u�jx��o��3����rdP�m{]��m#���gn{��1�cyA	���PR�J�S�b���yod���=
rnH�G������Q��n_s�R������^��S���g�=��{I9�ۺ�O%�3��v�:�u��Ì�/-�&�ۊ�ݹ��=�̺��ݻ�c�J���R����ޟ�MMK{}&vk��h��f�r.�n�w-˩��KR`�uA�\��GI��������e�&�q��2�\����W�\�e��g`��IX�/����	/���� �Y�d�5g�s���t!=+;'L��չ[!0�$�'�+�ܘ�t��]��1���۔�}]���2cw�G�����r.=�ɊUS���t���y�f{��s�ާH�,d�&Y�.����P�Tj��sn�Jx����T'}r�g��Ӗ=c�L`�r$��p��B���t��f{�D�,��7�����Y�|5<*�DOD�=�Z�����{÷�g
����a�ʊ�@Or���؅�b�>�ha�*iUPK�r�B���g@ym��v�f!�'k��9�W&|[:Q��Z^k�rV��`��l)�'}L���VФp��%�iHb�0��Ȫ��5�������7f��^5A��B�&�Tn;�3#k��ݎ���od�WsO������S�W*;r�����g>:���s�t���r�����!�b�J��ftfz{�q/:��W��V�V]ʏ�I}��MӀ]t��~��+���yuܦ9�e;ͦ��R�*8�)u�l��7+~Ŝ���41e���{p&h�j��"O8X�WAv�Ĳ�� (C��/B�X�>�h�D��E2�h]�c���;�W��^{.���^ir����q�1�^�2��$a/�\���7�wR�� �����:��$�p�Vf�����@��}�F[� �+5�-��!�N�V⳶�acڎ�QD[f����+��g����CP|b7]�\��wmѭ������;sv�el�oeسǵvԯ�D&��ED��ާ���|���*��B�/�d;Е�d�x�9d$[�y�1P��w�s"^/s������Y�T�|PpA
�(��ݤ������)ߒ��ɹO-�nV��{��^I^�X|r�w*�0V<�.���۵k����[\�H�f�<�ͪE"��[������{�j�J�ֶ��A��ǲ��-�5�o�Vpm�ͫ�uyn<��& (�8�Ӛ'7�v��v���l�'Yܛ�����*�ھgh����-�Nn��aR�����޼��I��vb�4r��<���1G�����r�9��g��&��	u��s�(��Gs�z�b���/�SxUs�kگ5+tNʸ%�7=��i�7�9�)]����f�3�;;b�T������HzJ����^�)*������cy���AQ�}��ξo.�N�9��k �HDEb*��3۷���ֱ�)���^�E[�˯=\`M��e�1���\�R�;K��c�־5w#V���&�FYΑ}��-�IYv�u��)���U�LEpQ ���JW���f���ҳr�.Nk_b�Ӕ"�mٝG&LM��V�R��)�	��d'M�3Q� 8�4n�X�ͽA��� �J]isg���ݽ{P��V�!0�W)�VX޺B#mp��Co��;g�UsM�/E[��vn�A",@���I�۲Z������|�N9�e���C�}����=&��^Y�������胐x�n'|L��c�e�b��0ɭ�3�1�<+Sɩ7�]{�Mw͌Q��2��mR��g/#l�="A�1O "��z]��t7�n�VF�TC�vP�6�gl�4&���`����]�=�53�
�鸣ˤ�����'y�}un;-�]�է��ŭ5�%
A�^B�S�1�)�V���xf�܉�9�9�:���"#v�O�X�a ��%t�{&�nq��lAh���c��Š�Bf���|�l?Dn�x7�,����1X��˂��z�[cw�R��:׻oiړ�m��$�fxP��:`z��&��9	��M�:10+v�b�4�'ED% ��
���:ݮ77�[m~=���ߍr����{BW�}�د�z�c�C��g�|�qc��I�|7nء�&=�^�5�>
; �X��Swk7o����%�vg��	ֶ(¤����:␼uy��X��;I�a��=�Z"C��ι������l���]�����@�s��z�����Y��OaG'OU�逌Ƨl>��]W@�P*�+��g6E#��ɂ����`����S	���ģ��\k78fC��qİG{Ng`ނ��oS��z�^\-��Mn-�w��rp�B�-�E`�`ۓ��들�t=�}[��G��l5�\��1�mnPi�0eۍ�[��#M��3�B\��t�wU�.����I�7�ͪ�Om�����T�&cJ[1ٰ�4dM��g�ם������:�w��:�V|$M�aKg#�d'��I����j6��x�6:Gsh\v�rZ�����x�m�E�����uvå������8�}��x׭��w2�kX��b[�N�N��_j2<�{Q�x��$V�"X��)){��û䦶���x�뵝E
:��.����Mg���m3�����l�{�ԙ1p@�N��e�
�o�$p-*����r+�k�]�1e���"'���U;�.μ-� ��ޔ�k�N2�wQ���c�����r�)jz���߸���)��,�I����g�P�;�A�~%_��1���D�XX�R���H�f����۲[4�V�*��
o�	��j�t	:]ڤ��Rgf^�I_FmVFu�H�i���R�x���jT�����3T�MoM�u���"h�
Oj�)eC <�ݹ>�'�g�UK���]Hb��{�M��U����s�1ޒ�w	Ԡ�w�{����<�(q�鷞˘���7�l\�SO:��P7��[>ų�8�dsA!�:����q����<÷��4��($�(���p��Gz�M@P`�z'�6P^fy3�첞��K��SP&yШYqb�y��$j������_.�^�Y�3���^(Z9[s�sC��1��
���T��`�*�ځ����\Ալ�-b�(�{�')�=m:wi��ew>���R-�z�k|+�*��7�9�|��X�8���o���%�� g�pJ����8�YWb͊K��j��ib��x�Y�#���c"��w�y5���]ֺ��Ðe����KR�J��.��.PP��C��H�뺗ܲ5i{f9�e�"^S>�)d��A��d�N��.y���K
��j���N��>ŝ�7��roS���x������T�GA�ܺ�R��&�gb��{<!&�MS�B\�ғ�Y���n�Wl�F���[����%þ��ǐ޶����j܏>��\$��Y7/�����Ð�w[=�#õqx�N���o<Y������VW?D���A�v�B�-�2���_s��G�+������of�;�s���u�U�m��E´�8�f'��#ٮZ���RY�~2�ڼ�^;^�b��z�\aY��ìn��ƂU�#m��<`��ګ�J��Zڵ ��]��͚����.��~�$����	��ZR�=�5K�#a��:{�m,�x��sK��ȹ 6�{vݴp���yub�n<S�u\�)�pbC3+Q�hU�kG�.�;p�Kٓ��5]�<���(��ց�&'�E�"����@����}��l���<�֪�
X�P�Qܥ�H�a��:�y^\-fv[
���uS��W��~����k5$�|��E�D-'����i��D��fe+7B:�R,\��s˰a]A6A���NȾ�B	�{ִwld���؃0!�tBS�}'�~��f��y�e���ɶmƨ�7=���5`v�d2{��dCq�=Z)6�n1�B��ޫ�)t��k����)�����y����`�a�N�O�)ijǖ��ɗٱ��[*@�!�y�yPvIcﮉ�1Ϸ�ڵ$�|��������&�~�M'e�yz7���w�kSe�.$߂�-n�f�����yC��mQ4�� 	w�ё�{���(z��3&y{t��M�C�R�[��\g�����}�;��]�_���5���Q�56�����&�����VcL�N����l�P�ֲ\.b� S+9L�;�e�.��]�|�u�2���� <�|��/��%K�뚗�W˺�	����w&�8�j����5�b	��4\V��Q���
;%\�}��B�Y�з���J�U�嬮0��_Cny8e�w9�����"g0��;�z㉖na���ӝ��z��w��q�oi�7�h)�ڽ��-��*{�X�TM3�מ&'l��"���v[���9����$:�s���+Vr�h���=�u������+^�-�����PX�[U���t�
[�"4�v\�fy(��k{��y��\�w8,4����q����k��f5�M���7C##�2)*�{��TW���kj��7]W�1NI���rs�)�;q
-C=K)u�9:�-�/7���\��	X�h]o������&��-�U�c��W�G�/'f��37)ߞM�!��yBL*����vqɒ�<P$�_҃���.�9
U�8����Z��9�p.w�[p�V1���d���xstvo�U:��)����;�yt��Z���ѩo�VN�}��5u	`��c���]Ұ}�!���C�rEMey��^���:��	��:�iʕ���#��C\�!�V��2�P�H�ާ�ײ�n)�蓓A�\�<��-u����e�<�o$�ֹ�̫5|�E��(
w�[��>�cQ�w++e��<�H��c.�O�R�K�q���2}	�۸��w�d�i�;O-O.�Y��uj���ι:�>�탛��ɪ�x��5���8�-�/e���]���(m�!]q��9�q�/�[K��)b�k���Й2�=����8�E����=f���:b�
a�=r�7^��S;��6��=�n9e�\�k
N+u��`y����ִ�ۡ�����#�ۢD$F����WA���vN�/]1;��}��||���1��W�Kl��%.����,��ٽ���yU(+�ŀ]t�gJ�4��"��O�wr���Z�Է=��C��Neu�B;="v�;�G7��.�(8-���l4M�=n���'xmoo�t�}���������]�"��L����bDp�f�y����E�r(��1[2�WQ�V���A��	!w�`xZ}�i�w�����K�T3r��z���k�.u��GL��!ݖm��%��2�=#D""9����j
MY������;�ji��$+} ��}:�z��eg�^Ѱ_��S���Ŧ�N���[�TH�ʷY�x�J�SP���hN�߯�ͽ �$�)f��0ٌM�[J��Q<)	 �k���W���hgyk�M
�+}ԫk����{_vݺ��ݱQ;l��o��p;��PΗ��C�Ǩ�:ܗ&�ť;W8q���R�J)��Ў��n�w5\)���q�Z��\�h���׎0�ļ��7G._*Y�y���v1U��J��x�h��::�%�l�̕�f-t=w9�9��8�*އ�-�F�*t��,(�2$>�3Jwq���c7I���2��諟f�Z]F豽KGnlsjb���8��:�g.�)Zo�d���ŜN��4��'���b~RJ#a�{����֎߾�Y��8�\�t��r��x���g������󉪩��tv*wf�
1m+�O9�fE�ĳ�3)r&�Ţ:����\�O�u�γ�B5$�hAi��2TT�uԆt�]iY-fi%b���3��6�!f�pSٳhonm��ۢn�E�e���'��v�UͻY���c�nU
�hRv���z>�Q�\%w7���HI�r!�SĜ�{��7:{�O ���r�ιx��+����n���Wz�S�I�t^}��q�k�A3*X�Y�{aP���q�\�;�s�sy:���r���㗞�ИTUQ!F� �ܺUm�y�]�koE���V^�\�5$�~~
V��"lk}�O����1�v�������O�NuT
��Nf��m�"Z>���33���v���1��xn䱎͟k(�x�nM�"��n�C~���֩�}~��^�]'>��B	T"���:flȘ;�U�����)�է1(2�#��mZ�Yc0]A�sնz��t��%}A�i�mW@��˝F�t,e����%���_j�Ǌ��]�&�V;�ۧw��{�%�=����QP�����V�-+Är�*�7B�p��(,�z+�0�u3��±�L��]�r�Y��x����=3���]t�@&�|�%p	0�*j�M��WS����kU��W;gJzP�Զ�PZE�̉b���MK|��5j�8Na��&��(�j���S%�� s0����6�����r'��U7+���U�j���چ���d��Ulw�iϵ�1�9{,�_]M3Ȕz�^fqH��ڽ_.�ET{�n��d��}���h�g��
۽9�V�=z�M�������b�t^���$�7;��1�ґt�{9��4��)u-q���dk ���W��a܆mDJ�����7h��ɀX�;��1��v��[	Y)�Q]1p�.S��廂^*�R��G}4dne�T|���"�j�CGon�uAj��`���UGn3۲d�e���rW=̉7���nv�)�ns1<��El�����D�k�Z����V��JT�Ӂ�L��*�*ș�ƴ�V�Qn�K�����!Ԗu֘�e��n���ԋ��N;�+5��[s�$�j]�i������9�5r*�l���#��w�]E��uȻ�q��/���Iӹ�__����l[P,M� k�T2]ұ�ܗ������ �=ۼzP��u��ǣދtr�"Ҏ��"�М>�
�gyiWnQ��>�d<QF-!�<��Պ��ì�sLP�+Q�OU�!�ΗOY3�'o�H�Ь����5n�Z��ٞ�|�+i�H�A鮰i��P#5�DP�4L':��Sݧ���m��v'�Af�:s��(���H4SM6�HՕ%��Fyq��L�G.�y<["�vA���P��پŮ�ޛ����1iدCxeږ�u�]Sߥh�ٔ�l	���"�32�]��v�9l�uu�>燋�]�v��Å%��x�v�M�u� �Z%�;�h�R_w3�5��S(8�R��x-��$�лqYP��a�ݯ	�HS�#L���'�n.�)k&j���[T�	�FR5������	wx��b���<�}����^4�����7Fwz:_�y��C�����oLKQ�8[�7��0�Ţ�6,D&���en�໹wmP���k6x����`qײg��%ʀVU��U{*��e����!�ȺmEVmĽ�5	���X)@%��0�}�������UJ)1���4!M�a��g�~�^���[@�È"�xa����n��hJ�U�o#i2���F�i�a��Xz�";r�m�$|�Xsv������6�dۡP�;-;�n0_)�h*���Ň�읬6��9]�G���H9A�w�5cX�{*�i7�{"�J��ᘟ��'�J;z3���S_<�'||���$h��Ԫz��>z�w���	B�h:����o`�����r;n1c1y�p�����χM0�1�Q	�����;�F��:�VM�:�qa��7+���x������D(eYh"H8����R����g�6:!��0�k2��Z..n:[ī*åBo�����
�}Q�|�#�WN�9�d�O�����oD��Y����Q{KN[ʚ����(�����[1��bd[!��|���y(�m�����ua����.4��8��n��U�\Z�^�����Q�:@tݛa�[�ʤ�C��Z���5��F6��L�}֤݄36�޴�o�#Y���~ػ��
o{7�<���v���^6�YU�`�B�]�yךfg%��r�5�P�_,�j��u�l��JD��.����򵊟E���g��>r��R�c�4z��SV��0'���v�K8&�|�S�a���u�����Jqb'b59+Tt���{ᵽd������VX!�7���Q���5A6�d��5�\4P]l���v&ϋ�[���:U�x6�a��q��맬]�g���D���F���1nm�����pt��������6�3��5��cZ�^�%�I�=�yޞک��r	{'q����s��C��0X�x��p�amHŷS�c�n7�v�{q�w.*�{O �xxenob��a������ٞ;c��m������+���X�T1�������(��k��LD��W�����o.��p��N�Th�����R{H�#�zf��IUq�æx��SB���ƺ^Rv�JK �P��{)"o��z�ֆ���8���9�0oJ�'r�n*�^��T|�x\{te����	I��[��j=U��5�����Qd�X8(�`<ѧA�
=�LL�̙�rvw�eb���du'���aS9xЅc�鶮�N�fM���}�[%���}�;j�=H��d>*m\d�E�S�@��=�4�����X���A7Ⱥ����Nv��6��ֺ]� ��0����G
5�JN�C��.��w��9Nqwp�OwFqU��&9�v�	]2g�Dv������v�F����<=��(>��U����>��!G,�:���cny��;��:��A�e�������c
t<X��0�m�y�۫F3�,E_4�b^�=Դ��ǹ�>�2����O935=��m��N�+���V\�5��>�
m;�G\��p��>s��M<�hkڣ�[��v��a=]�ӕ�=����M��M�.��դcz�n�+KF���hC*<�:�ԧ���z�˷:�7����}�Y��wb[�)0{ADq� ���8سpBZ���
[������{r�Mrs�z���9TE�R��9��l��j�nF3�Jc�D��kI��N���v�u�˪��a"�"c=7��U��ʜٗ��XpYM0b4�o23��As�T���u"u@�劎H���×�Xe��oV4�������톢�*�)��נ�+�pv[�7hUU�����k� ��{cѹ�n�}{ވǴ��I�F��>���t��P�B�w�<����z����j���H��M����[[>�HXy��6�U����K��̜BqR<��ܕ���60ێs˱	��-ޜ����ٽ7�f�bW�Ct��;~Ʊ�F�Ex�إ����9�s��2p�Obj��`A�[8^N&��e��u���4P���Om"��{p:	�����e�}{B�K��3�*�GlZsZ�<�3��tfܞ�Y,푩`Q��R�{�ｽUǑ�Sҕx�do9�i�6/:�q�2�]@�QD߬� -�Ym44�q�$3�atROv��b"ؗ�M\��齎��toJ<��uh)[�u,�un���(DFF�.��;���\� �]��Vu��c�Iv���w��1�$%�E���\]Ŭ��Vr2rH�ϙF����i+9F�^*��y�JWn.���t��f��� �~��+Ky;�ظ�K#�#���������x������'Sݓ݉j�< ����6�h���:����1EV��ڣ�:��y�Y>l�Z&���b���-.�b9���Kn׍�)��<��Ld�D�I6\��T	�O����>m�~�I�1��w,��O�YX�qrH�WG>�<�h�(��p�1UvS�A4��o'Web����/:�xF8t�=[-���ͯ
n���~U��_-t�	$Cj��o��ڦ�\�Iqi���3���},G��EVd8-�I��	{�oX���y��{�Ū�.�y��C9���� ۞�WD{T��5�ɽ˭[�=�!�I��_�)��PKoO����irpOuU[��v�U�0\��3%���D�N��g]zn��wi�Igq���Y�Z��	�tFB%�8Ә�ӄ�����1��lXw.j���ۼb���ba�ujV�!�2�����.�'��Kit�dڈ�\ўZ�]`�!�l;��`t��((Q>��h�!�����a9�����|�ad`n�L
���P�lc�+z�ըK�<�&���=����u�׮�����c@ �DD@lOn��؍ϫ/35�8�R�8�1�e��ں���r||E
]�s���X���w���r��N����>����u�n;�]:�^�2Ն�L;�S�Q���My�dB��@����o/v��v��{iza*ک;i
P��g(,�*��+���_�Z�<r��5�y�Uי�����2;wkpR���S�����#]�i�7V��P15^u�M
Ȯ�m|6��Q�T�2��x������6s���ڗyj�.��z�y��eaKB��G�*�0�S��J�Ip�ӽ�[���Ȳ�]�X�!حm�����nX�a6���U��6��-�5�ͽQjw�Uѩh�%,���g;e�w�zo;z�mї����x��L��e�0�,wx�]�Of�Uۻ�"a��NGIX��ڋW��ZU��l�M��2%��)�^����"�n������s؈�%e�ș��3�̥k8��B��w�Qt�l�do��t�	��d�V����S;�[Q�oKK�.8�rt��<G����7cr�ic'As'- �����;s�NR��[����Nx��ݗ�:ŭ�.<���$C�˲tvں��˸��Py�lc\kM�i��/'�ۍv-�l��X�h9��ní�8�ϡ��ʃ�	۲�=��Y�{�{;����︘���m�^�]�n��Pz�y2����=��֞�V
���OF���)෩6Dg���a9��c�m�n4rF��ɺ�pa���5�v�:���Ȭ��%�L�͞���=��,�~X�����&�����T,�T�ZA釆_c�A�<h�P؊Ն)�LWGaW��;d�Z7jh��b��]�=	;���۔��)a֗{yWN��<��3Nඵ���:9h܅���7����{=��lM��K!��,�\*�ۏq�͹yF�Պ�n��TyyS'N�w/�jr�\�M:�Wci��T���W���P�v&���ʟqH����in[���#}۴.k�з��8� ������۷]b���E��̝��S<���H��|��41yў���oc�������&w���6��D�^�=Sp�0����}����m���kc$bQ�e�n����V�1�5$���*��յ� ���c�����j'7����8���z�N8�r�V��@׽C%j�o����q,��E�5ޙ
9���v@u,^�;����k��zC���xs�/8�HJ�q2���8p
�d�	$�IfD�Ν{�"����j�O���2��i8;+&aGE��ȉSi�ӡ͋��E)�KP�ywF�^NW�'q��@�b/t"J�SY�-T�F�`̈́`iy�X�-�I]r���@��n�^�c��50�a�%gZ=�����E5�l��^Yg�m����%��#�X��|�{ҹom+����:|��]Ϧdʛǫ�
/kn;*td>��p��gt4S�@�a���Fa�:����u�I4��w^���&dtb�d>.���M���YCAg�.s_<n�{s:"�#58��6:�S��U�R�U$�5���)�{�oQ/�6���Z��lވ�R�2z�Z>;��|���	i�,��B��̼���{�݁zʌ���K����b�����q�(��������Xbɛ[1:�-�$k�ػ-`ᓒ���f�[��0�.�>�U��Gq�v���u��E3�'ӯ��=�׵)[�!{��*|��)}QU�y2��4 ��;�"��iCA�!�o�bQ}Ԯ�%�2�]?MJ>��$��n�Ҫ���,I�3�,�p���ڢ.��h�};���u�\�2�2(XZ��泵AI����i���D]��ˬ�j<a�o����:<'w�]ɱ�cձԶ��w��(�id�je��� �\�r#��& �F���,bn�UoN`FЖk�]3Fd��[�_����%`�f*��~���3R��k����@^c��FJ=�0�e�d��q���^&kP	M�Q���o]3���W���w)x��f�->`��R7'c��6 j�eٚ���.�}�Ep�����;��hJ{۬w�f�"�e�������ξɶ�2����36F�\w�,�i��ƍ�qzt�}�a�Y�]����p�yy�*s%b{�։R;E/r�v/q����l��E�T@� n���� ྫྷ���R:�7>����z�rAQ3���q\h,�6z`f�=l�y|g
��ˬ�!���VX��$�P�D�j�"e��Es�9F��i������*aI_#���q����j����-��T�C��u��O����z�pa\�y�w]Ѝ7l�e��ԑÙ��^[Ve���W:���v�!���zb���V������G*��������E VR�Uf��k�男�l�v����YV瘝H0�w*�2�A�C����c���Vo�F�^����7�.��.u�e��:��-Y@X*�͗��P����W-�]����Q�6�3N��Zc.�;��r6 _��UVn��{P;al�Dq�ÒW'\Q�� �-Ʒ{��mim����+w"㔰D��"V=��sd�J&��v�4q,�qry��jPd�_�.Z��}�����%9!��nT���S�3��ص���;oV�܈����u�;=7)%"��HP!`������fpz�Ӽ'E&z������]]�̥�gxri�p�{�4���D'���!�����yK<����Z�0��K���t� WN�p�D���l7��5b�D_��ɾ�YzVo�:��n���B����'���dzr��������CJ�J���M{N��Z�n��5�#�l�u>��T6! �1^��=�#�0T��Ә/�a�)�{�xl.y��F�oh(��T3nk��s���3��OB��|�ܗ	9�M@k��"{B珧0ge�o���/�v��jV<>C&����lzW��Q��ln�%=��S�ҏc�i+gn�p�L��;n�o"LH��㍾�,�z�%���W�E$��<����1�o�FBj�ቜȋ�s7UAF�Փ���)R��J��L�c�fQ���c���C�n`11Ep��uY���&!^l���"�`�e>�o�gT1�oq�q��(؊�3�q<.2a�C���U��>�ű��F��R.��CBj���cȹ�B��/&a2�ՇX�Qu���d�V�N�{/ZE��H9�2�4,Y��Ɋ�/\z@gF^��sv�,�Ln�4���c
����V�uqKڳ��ky3i�Z��2�F�L"�	�����Z�JE���>�b���f:tw:�I品�;xv�ξ,��EN3�ý�eL��L�)8�V��s�wM�סVVF�X����k�X����+u=��qwf;a-ۘ�T�xueRX�C��<�}{�]�$}��(�W�NY-8)�Vv�S�g0�3a��\KS���,;\�.�U�d\lh+�Cs�E
fw�Db��!/�M�SRdi��6K(Zg#�hҁ�h�N���3wd��2�Ā��.4�m�v*��n�tC6��Gl�a̝z����3�n�iv��D�1�fNǔ:��lκBc�eB;sVm������x� (wُYī,)��WE�e�1�1EJ��en�+��۸�����ᷩN$�^*��e��ϐ:st댽����1fh�t7�M�Ga���� Oli�W��m�V+r�e�[�lٌ�s~B����2� ����v�Փ������w|UW\�����Y��!����T-둽{6��^�*a���Nq�{�w��n�O����@��D�s@�ʪ���'\�ú�z�=pYzm����w/Gk��M��iV��`�Z/rgAi{!m�g{9x�d;WnӎU�X�r��w��70�à��ն3���n79ܸ�1���Ь� ڴ.E{9y���Ʊ��XL(J;�v7h�n���r�\֙���:�@���N�^9�:���#�[���.��G[Н;]�	�)�n��vf�ۮ�iJ�	�I̾���v����v��څ�5G���n�	벯��=8V�n�GK�'����k�[��V�L=mT'����c�׃��z(�(���
Ok����n�b��"GW6}uE�p�����u���"x{m�]n.�H��F�]c��)�=�[����@����a'�g�Wn��[�om�v*�#�Ҽt�5խ�0��Q�*\'cu�y��M���p� ���c�����1�v�����zt*L�s:+����Sm7e�5^۟/��܉���ce���v竔�vc[㊎@ؖm���n;q׳�����/0ꍊu�y�^�lO:�,d���W{q 3��w]��ڰ�`/.u�[Ǟn=v���C��He/;Y3��ہ��e���pc�(k^�4�j�ý<nH9�ۮ�R2�����n����M����i��6�yx�B�]��ˋjܚ��	�)q��t��4k;]��Z�ݎ���؋v�=lϭk��n�4�n׵\Zm�z3�Ѻ��8���ZP��GX�@2�\�Z�6ܚ����A���R�����1�k;h�[�圦Ƅ۫<r��V}��3v�Gn��qЧ+Z�;�y�;a��K�{{�-kuZ-�mv6��F8�)jB��=p��7GA�v�������٧7/N���\e�A4#u�5c�ՎN�g���-�ͺ��E\GJ��;s��p��nm�������G63�=ug�7���Rvݞ���6y|����v���Wdy@㱌<�@sr��OV�o�.��NV�j�"���<rq�e����5�s�pv��ネ���A�P�Ϯomwn7O��r�<��ƶ��\u�S��0��ۥ�n^:���;z��
���`Nm��;���)��8�ś�]dy��yΞ�m���v��lЋջ�Ypv���>����6%�nƎ��l�0��d�R�[�oc!�ݫ;sɵ���nl<�qòm��m�o:��W�5C�S��V����%=�f� '[`�������:�pf��\[�OE���ݢ���n�Wmi����@�섔����Γ[�|�K�q�~n����t(��Az��(�"���Y�E��l�Ĵ��o�1�*��e#V��@z�TQ���嗝��S�[=(LƝ`\��hW-W���z�w�c姞Nc�C�e��C֌�H�lB �li��;���6���ᅣ��1�
=�qlU�fVFmr��C��:C��Xn6�`y;<��U�'8�1��6T'B��q0Ŕ�'j�9\��{X;E���V=5YG��e#����+=ͽ�7u�J�c�,���ۇ$r�*B/y:܋j�o�ƀ������9
�����L��eX��lKj�ȃ9.O�q�UK&��X��)�`�p�;jj=�1��F��:#=e-�E�R�bCd96k��+v�Y�dj5�zҾpo���qۏ���d!r!�	�, Ξ�뺙�<u� ��#1�^�6�S��*>�]^��N��C�|��f�o'�T�yEԼ�[S5��6�om��(��F�8���=[��$�/�}1�<-�nZ{V���yu��8���sp�2�Y�(�{woy	j�ޕ�ʺ��\�86�62�Pյ�\h���mzZ���Uu
�7�>0���#FfZ�)r
��Y��t�=Q22�]�t2AY�ײ�B�P��B N|r+�^#u�����{�`��w5�7���̎�DKop�EC�A��߀�X������YiNz����b�]�r��R�R���Èf9��.�ܖ9�<����j\ǹ0�}�U��@/���[�����+��״(�*٫eʝC1{h7�ݟn�����gڑ<��4w;�^@H���}�cMLK�qy/R��Y}7�(-ӛP�Z%d�O]Eaݹ1�@�΢�Y��mmj���ے�5-�^�{8#�����a
'�^Z3�[�)��x��ƈ��P��w�����z�Z^,�iPF�񩵺Nq�묬);�1�Vp�B}��b�bT���Ày�?a�f�]����)H;#$�JIY��G���w��p�E���vo���\�7����J"�u���Ɉ"�樺鈉�8 ��d�k��$d��i���lM�U_�=�u���Oo*��6s�G�eXv耳Z�x�j95E�0E$��9B�s��M�b�����Ձ�����H�	���{2&<��OkTa�9�jT��8xL.�`�	�`�6vT��F��e��I0�ww ٚ�yz٘Jrޛxﰣ�'�f�%��JAk�s��2��r' � J���wl�[�^ڪl�!IF�i5��^���|�\c�z$�F�7ΗB �f��ڲ�4�goP�1&�tm�E[��ߵۮ��]y���ը,����]sk�f"A���vv�d�C٣r�J�vIT@��QѹI�o]ɉ�W;�kl܈�L��Pf�v����ʝ6:��6����^Z���؂�ԿM�◷R�f��W�Ў���ϊ,��n���(2�ޤĊ۫�J���m�*CS���ΐ	�.Խ{��.P��.�eu󊨸��Ǖ��4���J��1J� ��E����Ι���}smN^�T�2�~�\�,�Z7���k|����3ӊ{,Q��¦7М�r��?"�5�1�i�7�^��420�s��Қ��GP�Ƙ������N{���v#q��C{�-XRjC�@����Ĭ�Ie9� Ŷ��Ɋ�]*���JyX#p^QJ�e=R����f�VEC���YV;�cz��y���� 4�{�;U�+��r$]R�I���ݾ�W��!�X+(��=��o��������y�&`�$�1S�b��\��Ձ*a�c�w����ׅ�{�j����_]�_2d��
F'����M�0 w񜪗��S�Wb���ħ"un6;@��9D��޾���pŜg�����^(��w�t��%ˤ�KԹB�8)�p��GjzU��#�SZ�R��1T�/SP�0��"a8W"d��G�y���b���<؃Q�3��c�H"�]�4{��4�U�����&+̧C-�ld�s5��:���(��Z|)h=s��ў����u�K+��q�"WDv}�������Ss˛~^�n�\3N+���dF�T��Q�m�"P�/RtW"o(�l�d����2]���b�&c��MQ	��1\�K|VgC��ڔ-��k>�����gzb"j�MYX*��j�%�}�v�s8�M�u�3�@^��RHyw��:��7Լ�����=�P�'���{�y¶�R��x�����X�d�0�Cէ\ٝ:ɢ��c'�,��tpB�V�$��"=��#a�L�vF�����,۱����6����"��V�Y$R=�Ӟ����c�2�r�S�K(�x�t�^�kڋ��[7%�́���b������ݷ�9\n�m�����v9�;1@��N����ǎ�l�rX�dێ��C��j۷�wt�v����s�Ⓚ|�
�nsIlF�v7n�s��j��z�]��� kLr;�;k�[�&n�˜GL��k�qt�g�c���T��d͵5��Ѝ�5�x贜t;��nݮ[�Z+��և�Z�^��@x���p��0ۄ�!�)��&i�w+�c!c�������Д��_.�q*W�8 ��S�n��p����(�*PdF�pt�!3��m��EAp.z(P̵�uư��2����/�ck���4�71Y/w�Is��]o�OSc1�᫥��Vt�@����WX�c$u�:�i�BT��,�Ӟ�E���B: {
B��M;t����8���[.ISY�xڼ��>v)ׯ�*)�O�i��=��Ma�vkP��I��*[G
��>��:]�i�*��nsu�������ӏB#jGc�P:l��}e��o!T-@�oe�4��$ax�y��G!:�n�M�X���>�!ݦ����bK�Vn?>������g�<[���]Weέ���M���w��]d�I�Mƒ�8Z��lp��WUD��_���]����c�SK�p�\~�['�4Fdv�B/�h��jc`8�!Ǫ{[�w����ր��~���$
@���E��s���`DF��w3{���|,�|��;�a�ڻ��׻C/_�V]�-9��ע�x�x&��0$�i+�q
1P2�\�S�/��ڱ�є4>�G�,k2[
y\���X��b7eh3��@+�Dk}�Q���"�n
ze����+Z�2�������&�����q��ǘ�rȹ��Ħt�4/;ui��o-��7\�$d�j�Pp��oyܷ�
�iϻM[�hZ�܋�'1�=s�(F�@?c�^;D�m�����]�{�٩�����ߓR.��:�c`
��B�M���/��Z�g3`+O��q��t�
���=�C^��0b"'�ɺ�u�.��7�\y�z��j��vdh��JMK��-L�Qֹ�����fm���i�Y�ا\���v/#�%�(�a�	�u�e�!R�̮��Sۼ����;u1�0)��P%T�=�l,�S�0��^Cf[��w3}�Ύ�n��i�� '%n2�Z�Ӿ���|�k{�@����;�Q^��3�;Z���@	P�]U�`����K�#U����#�p�)h�xB����&��D�((P���@���ռ�nM��@�J��bmNs�ɧ浼z*��'2rb=�o25I��$�c .١U�Ý%�Y�lИ(�N"�ڛ��DNh�k ])s��p�<��	=��l�)���P2�B��E8ʔ���"��J�g�
�Mkz�������"�o�][�pS]2�]J�V�:�L>��Y�т{c)���r���v�������ŷ��y�!RV*bnmV���s���̐l�q]'݆`���%*��7W�g���%���@s����V�s!@\����T�UtAL��̭ʘ�GCj��'[vp�O��YR���̴�,�:A0b���JF[B�o��8/:��״d�V�0��j�#vQo������(�R�3���j��<��ay�{�9�z`K�1�9]�T-r�� R tH��ާX���0aE�G<w$C��l>��lx�7y�K�| ���W��R;|rj,@;�&��D��TsH
�@G���D�ϻR�d׬�5!2���C�-�<m9j������R�-~�]qd�$dl��}�����}Y]�-Dn�V�h�:��&�r�I���Tt�Ou	�3I�B�o<��,�YH�{3��r���Sj�_wci��ܳ&�އ�����7v3n��n�qKN���oq,w�W�d#�"�Y�X���(j�y.�]���ʇh�[�IX�N�mokt9�b�ff����j�҈Ƨ�����.B#���X,(�q)'U�F{r+D�r����]\�N>g��챶��I���+5�'5�;vF��Ǉv��^�c��
gvn�*3�E��#=Q��9ӽ��0�̆:UmG�3tS�>��}��՘��H�O���8��`�*'/*o���>�0
�(`ݒIA`��ƭ�¼Z�N:���(^
�����{�I���灔������o�ۣL���0B�tˀV{	���ZC�+@���t�Gq^#��a�U=��GC��e��>}#�;}�=���=m���M��LKJ<ٚ~	���vz����R��w5�躾܋�*")h��eM_&	ʣ|�!F��Q5���8-��3TЦ���:�&ha��Gz���D�1B�фʮE%����x���Y9�C��9�ݽ��7����QF�#�{�FU]Rד+K��V���f�2�b�ʰ�>��D�x�rdNFFsYQ��A�vq��N٦X;�B�ķ��L�C,�ą��J�,�q)�Iw�c��d��|+����Q�'��݂vN�\V܂�0u����i�Gr����g�q���\�{{����ۍܷd��4��7��k;���ۨC^�����ێ�v�:�ݗ��Q�X�|cuc�j;W'�'#�j�4��cz��*�����h+��s'8�M�V��
������Skk�*.֖�&5m��î,��]\k��t�ms���'�>M�zƋuS�Ѭ;�b���Oi�}I����&Z��P��z����9���;(��,z٪?���WrI)�b��vT����׼����}#���W^��i��?V�����������-ou�3��ދOeB��:D'(х5"a�ej�r�DVO�8�7X�d]���F��uÝ͑�	�-9�ox�sk]t���]��l�紟Sns�B�ȥL�zN�]%���]��c���=q�}���<����\g��� ��^��4����/w��oE�o���9�D����S̵7�Lgr\&.�.�r%A��YS�&d@o����id��#N8e��c�"�f��Q��.ae�yqp�&j � }9V�w�L����Z�Jϔa�y(�A���,�)�W�L՘�������A���0�T9A���a���i=�\��S.\�ʔ9����k��-��K���z��.�M�m���%�\:�pmB���Ϡgn�׻��=�W�h+#�l�"�>�Kf_UoD�e�6����X{�wt�;���E�˟$|���.B��]Lԫ��@����ze=��`(U����W�����l��7�����z���E����=�c�˭T8��n�N;ӵ�r�=���h2��6����~~���voF	���N��R�V2���g�;csg=�����C:�}U�F�7i ��l�j��%D�,�0(�jC����wYe5�����O"��Ы�����UU79Lዒ��W��Hr0a�gNF��mɗ�ض=�{�Ylw�KX;��ހ��6�����k��t'�O�k;���u���N8�%q�"y�0�@�`���	79R��W��+�t��5=us\�;�\��x�p1��}^�Ÿ��}�����1,����;,~���3|��4a�$�Vp�B���F���g/�%�����j8z0�d����g�9Y*dq��V&Ie+��{=�z��5�~>j���*���7�����e{���$W���7�v1�i��l�O��ڲc^[���T'A�P��_d̼X�.�%��Q�r
"�aY<.g��M&6�t_d!i�l���F��5�a��'�b7m+<3)����0҂POŤ��U\'��1F^�c���Bf6gz.�!p'{�]�"�P�w+�"D��\Jy��,���^�!��;QnY��܈$ލ7T*r
r�1�#*'	��9�gX�b��Z{7l�L麹�3�p���imfa�zv��Q�}ю(ͤ���V�h.���ަ�7��i#�v�<�Tb��P��WTt��+�F<�V޲�qk԰lˮ�+������vp����^`F�u�ٹ&F��d�0[��sI��̉O�ݜL����k�&�ϰ��fÜ��>���Q��]�)լ���w�¯:5���h_co@�ٻ�h�Ŕ3��bͺ�K�"yYC����4�F��1f,��KB��3g�NZ�a��U��Q�;��Ua�"��:ԉ��%`�y�vZ�n�	Z�2��Yw33%���۹��7QJ�w(��ͽ�R��8o�7����5�)�![ �C��5�9u;]�F���iKN�b�v����ݮ�6�=X�V�:2+���Uܣ��^�"kF��W�g	����ز�(,ٙM��u��S8�.r��{��Q�zv?�E*�:3k`ao.\&$�]9�|Fق��r}9fk���Sk�t�b,��[�3`��b����'8�l���<lމ���Q@e��\�x���l-��+��b�6'�2%�%���[=�{j���+���K���DB8H���u�r0�t[:��!k��eۃe
�bd��]C
3W*?-n�R���获V�i�KV
��փu�b�b��'��Umx�1��%���V7v���]�����'@oa�ʃ�!]I^��w�nw ��wNč7[�0MVj�F�0vFm=�=dU�`rd�ף1쩈N��Cw¸3j�	�7�<C��R�lf��(2����SM��ɇ��P����r�����tN;#�>���UIP��|�ٹ��={�8-X�.Iq�,UWm��^N2яo��ݱ�(���P&}ǔ+E��y7e�R%�Mc�n���=^�l��~�x4J~&��g��)R�,\Eom�p�Q'_M��bm�3�jm3yRS���(mJ�LȚcq���#���:'Y�x���kX�;��i�+���쵓g�	n��>1S6��a]�>Bbp�����q#s�z�aȂY���ӓ�F���MA�w�nuXns@�G9",u�"�������h��kM�lw�~�u��&x��/�4��uy�e;�f`��V�����9�^L�%Z��kkUl�Ye�r��UQ�$9cl�+���8{[u�x��ďMTD.�:�#ĔGK�f��d�DҜ��cDF���ɱMO(����N��q�`֓� Eֵ���x���8*�E5���t���6{O�ҷ�2�$瀱XŜa�m<J�cmp�rU�z8��D�*ՊV�re�,� ��s���&h�u����ӽ]�������@Vw�$=ړ�\\�?wX�9M.�y�M��	�B���o]��x<��������O`���!7z�R�#�옼Os��X�J�H��c֏����n����g�|}�jXnIR hYۅ���[��d�wWu����u�զ�Gŗ\���*!5$S�&Zsj���U�3
����� ��B�D!dmg���W������G��Y���;{Y=t�+�3��^����P#
�Yu/{�8{F>o�lK���XA�0z�maX�Z/yx�Pu�^rJjy�st��m�3'}}�i����3[�c�5�����W���{�E�
�10�j�]w�<�X�Ӧ��Y;=�~r�*�.��B����z5LO�yվe3�4򩝞�[�8������p[�{|F��D"b��E�)-a�B]�N��B�m��D$A+�0��&��r�N�M�n��f=P�3t�G�̶����C�1E������q�Ȣ����fhm��]S���VxE�T[.�/2�ITM�4�`�����
ٹ�eG��N��[;�M<7���*i֟'n��ɒa��U��B{�;:�ܽ}�S�%V8��-���Ya9�oX�
�rذ�7[;g��@�Pw&�Hn;l�eH��ٹ�[�$:��zkn��v�����nݸC�b�ul��v��v�pO�M��}xb�9�n�V0'Y�ێ�$O\Tq�@ �����n�+�Ӧζ�v��[���q
����]�]�\�G	�V�nV"^�n3=�� ,�m����pzب,���8�8ѲJ]Ms���6k�N.���t<3�����r��	��-NЫ+�=e�w�{[�T�`C���+z#�*��f=��-�V�#*4�^ǜ���Ą���w�7���)�wfง�'��U��A]�v���@2wik2(��<���4*��c�h�]X*+��q~�s�Oz]��� H2��-,9n�(`�gr05��>����Ư2��!T�ۭ����g��l�)���6Y:���U�)�&"}2;E��
X}7��4��L~���������:���W�r�|=���R]�I����ꂭ۳�������Nm��qo����I���M�1_Y�P5Q%@�	��&�ndwW $�ɔ��ga�im�+l7�D��]oF��딦w���Y"u�e�U��Nk^r�1�P��t��n�mù�h6�+I:h��[\���[]0س���.�G`x���t �T�n8#�zi��8�j�w*�j4��5��s�wJ���Q�$�*˼��$�oY3�U9:�Sͫ
�Y�8�2.�1|v�a�Q�������J����vJ����%+�X��)	;�r�9���$�!������i�����e8�V���5�j� d8�ձk�q������1eL�>��B����N�����d��˂#��@�VE>�(>���e�񆵯h֥�OEȺ{<�]�K�1��t[��h��yL�ɩbq�s=襤��`;J�mu��(��H�����7�k\m��ݽ;��.*$�ٽ�rS{��R1��x�e	�*�̡��0_#�W=��i��,Ъ�1�	��#!1�Bc*���*�ڻ�u]tS$Ն��,�������-f&�vN^��Ԃ]@ծ�;��\��I�f��rPN}����wޡ��Svp~P+v|��]�k��8���>OX��r�Ӿ}�ryl�i�u�%�6���<w}Q_��HUQ= ��,�6�2���f1X�]��Op���>��O^E���Ǟ��<XR)ݠ�v��������͎`#~q��E{��0�Grd��XԴ_�
³-Z�M�4��\�yee@�*��O�MD�;������Q�L6a�mf�Gm~C����>:��}^rQU��ELs5�@vs1J̞���)γ��S�V�%&�v)f�Z�x{�_=�zrn�}�e�=�k����,�\E��91i���L�vR)���f�w,.�ͽ��wK^Xr��3y��6)t^�u��d�p���������:���#���L����h\7��J�A�5�S�{B�l�}tU�$�z�c�s�{{wI ��7���\C�Vbb������Y�\�ѳ�J�t)��1��nZ�K���e�2�w��������*�u��\E��7�
&#����CڊI��FB�ݷ*stW#��ϟm�ܯm�p3ڍ$f�5gK�C(nPP�D��p�w�w>����9b}�r���j&���L�5��#��4�����������t�����<�I}\	k�H'%&��«�V�{�7��[��7^�Ы4�t�:-�����Al��T�.�x��z����ƭ�Ĥ5��u�[q"�D#�`8�U�&zs۽zžg=���5z �N,��9Ւ7je��۳KM���8fFê�w@������aw
/saAU�Všmљݽ�֭��*��s���Qb��v�4
(V���>ɸl,Ϊ��k��v�u���y�TYq�K���)b�j�<#�����!�ż.���9����quL'3��� an�?]��܌M���*&�*�\�kU�-�1A�$��c,������m"yUn+y��J�*.3�qg�W��B�7�˹�Ee� ��5���VL�SGݖ�P�U �55f��&��Km��.:%�o[tݝ�{u�v{sv�fyD�o ;n�5�S'�g�?��Rx1��pdMϠ�G)���|0���y�d��\/�����2y���x�e�Ue(��W��M&��-jnI��[�V
b_�]��G�^�BޔJ��[�O��3+��y����� ��(�:�_6Z	h�7(A(s��6����k�8n���"��%g�� ��o��X�o�/+�`�/��,a�w�E�Ǳ6�+uEM�"��6�]�$:�� ��R��4x�����.��V�K{��(m�YB�^5�m���E��/&�6�ω��_1���ׯ�P�H����Os�5G��M>\���z,��;ގS����YE='����>��C�6ƫ���(��V����q���.{��n����:J�m=X�����fg���ȍ��pt�ƅ�ƶ#s2�
�-Srj�բ�3��6s*��g8H�RS�!"c�g���[��׵����St[9�`�c���og���V�хƷk>��G��c��]
p�ɓr� ���<��v��Tnx�{t�c;i�cmOXM����7EY���a[\���헙S���֙��ϳ��8CK�<�!b�ZV[:�δ^�W���m�F�݌i��n�ܼ�v:��u�z��m'k��m��Ճn6׬og�}�B��S�6�������P�	����>v�����:`݈LB	%&������[��Y�y��u�~V�oB���O�㾭YG)�u��0���ђgnJ�͢9L�_Z��]���)*��(��<��S;WN�Ǉ������m���c����S�=��D/�-�S��~��IpA^�k5�s ���Ba��U2���4�PIm���]Oc6َ���'KQ4�p�b�ˢHE΋�N�g �:�nlD���K���v���
�7��0
�A!&�!�|N(G&�)�{j���첆F�:*�e�{�6�Ps�9��Gt"b"�!Pނ���i���"8�9Ζ�]��2Gi57mg5��yrE��־�aWmn�(��=�5E(��Yo�0�:�6ȝ����IAc��uڦ7�]�-�U;+Њa3F(ۮ�t�Ӷ�=L��5���pmc`��<���ܜ�)*�����^ߪ��b��ǯg�U�b�E��Ớ�%��t�Wt��?>z��v�dv`yse$�v#�j-�j�����SR@����'{S8��~Y(P5�I�q���ٲ߃~�L��3�&�f��k�5D[���N���i�zܭJ�����c$��=n�p�ƿJ�}�Zu0X���v="���1k,����:�R-̲�.E��T,N�J,��&*�o���ʈ��A&�BE7-%&	���`6���#��@* �I�g�^ۿ,:d�J����-<�Nk��Z^/�'At���
(B�vI�w2����s�r�re��+leF%h�\���Н�ΏQ�,Δ�n*mr�y�I!��|�5g�`�.�nLk���/_�Y�j��*Ԁ��k�q�t��^� r��Xh�o,5jC���0���X�����Ȏ�Zp�Ԫ!v��a�?fBo͒��TR�m�kA�s���<ƱD[F��Y�
��m�b��r�#�,!#n���\�3�1���wN�4J���G��5V3�Vv�A�0tվ"8ۆ�6�Y�rX�ŭ�z���J)]���"O?j\z���#�{C�ps�6���2"�;"�𱉴y��ݏc�/B⭖�Zs�T.��h��:iA�`�e�ۇ���;�0m�O': VP�x��V���t�=V��6L�(�2`щ���M̺k6s}��v����U�t*�ؐ\C�/�X��@.��"�E�E�Q�R��r���]*Lv��u.䊩�y�� ���Z0��v�缤��DKe�t��uiq48)��ǧ�f��:�>��k���Ҭ�.t����m��4^]�zE�HJ輑U���&�8lQt�b,��9R��v����z�vܹ;�|���E�-J��2nY�".�;a�crZ��C3)�a���C�{�n�����@��Z�9�rS�u$�A=��x�K�GE��uN�;�ɓf���眽q���LJ��Oi��=����.1�؋Ρ�7��EYJ���1X�L�!�ʹz��)�N��):�7����IJ������	66k�-NB=��h�*�;{��^c�xM�s۠�}�`���
���ߊ0C�x6� �љ]�ڜ�Q�Q8^^��s��hb*��+�Z�-�sA�B�����}��IDA���S{]��[Z��N��c@]���w�Ǌi�o�[�+�����P���!��9��k���*��yG,�R�ّ����=6yѷ�x�ޛV3joߌ����W�r1���|��)@��7y��`�-��y�o"�f���4�k�֎�ٽ3n���.�e���;���f��C4��I*%���D��9��M+e�o��;���c��t=\o<���m��ӇE���z�pNe0���B;<V)UDH���ip�7U�L[����v��v8ܽ�a�`���pg�8��\���	7_���o�^��דW��pVǼ{7���@��~��A�qb�3/n����3]WN[u�����	@"�2��]w�k�<�[�G���^cK�|�6�I/r$P���,ծb�dTwH7�N�-�a���"�͵;�q�zZ�Y`:&�$�n�)<*��%R�}^J�e	e���S@��H>�33��+�Y�هo��������k��+��$�B�0�� �m�+m'慴h����2�򕉸���s�	��[V�!VN��ٺ�_<�����l;�7�L��2�ɱQ�6�삵�T�KE���=�Ǵ��K����~�U���{�/+��>�
�l���&!�KR������0�r�8=���U��ؐ�Mb�j!�c������"��w�2���W>�e}�휞]b�_<4-z1u�6gUҰ�s�x�s��XR��J���dM<��1�i��x�1�Q����Rk�K:j�f���~�T�{;�ɼ\b���HB-�"�D��0r�٬�/L��1vU�gF�!ꃎ�3A`�:ڤ�䝹��Y�SC"��x,�ӄe��8�����"*!�_r��(l𽔼�Ek]�S��OEּ�t��oB"���,_bu{i��F�fƏ<�ۂ��js���"�WG5%�ٜ���]NB�B��}�����梶��8��c��#��k�v�]�ط���7��]Z9VxdŘoW-A|�֎����i;*��X��٢�|N���3��ҳE��%�6-mZU��H�g��cE�;̝ݽ��uv6w�W[�#{���c/ jWk�{�,���x��Zi�X�݆�Nz�R�Wz7pPy�t�v��T0�VA�	1]��v�J��}:\�k�D�� �Hn�.%l=t�e7���|M^�>�I�cj1jH��B���Z�.� ݀��=<�p���uΟkQ����5Ĭ��VȧwI$?v,��:t��xW_uL���l*���O�t(eɺ��7�7�8���շ�ʸE,��s�p�mf���r�}�f�,���v���7.wƀ��e����V�_iܴ�;��ۀ,X^���vn���ke�ޝ�6N�4\=�'3�&����O��ܲ�3;���B��fmd�h̵�jU̽-B���^�7��9oq�2����n�Д��j;�I�I�����6�����B�۱�I����'kۣh�w8{h<ݦ�����>���"��mN�=n}�,��ۥzř�Țy��a�	�^܀�����OUx����vZ`��=\��ݮ�۝�,����T6��Sqy��/X�`D�^��_]��ے��k��pns�reaS��n¨#ڌ\uo(���Ϸ;@ɳn�y�j��iB������8Js��v÷�(�;s�r�6�vDn6�,��:���/e����Ŧ�u��gn�ƺ��t���kp�n�lgog�z���<���;I��b�2Vc�v�7<=��s��nՎ�����q#�Wg9�[��0�����zqs�ƍ��;vD���s��{B��r޺����&AE�w���pn8�6Ӄ�г��{[!�-/�b.ۭ��¶��V�m�^vFĉo6���8G��웵q��`J^(�̛��[u`�����s�V�p\���l򞰌�&�up�n�*���c��v�q�9�=�+L��%�<�S��Ԟ�v'��ۯg�]tgOjWp��;7��P���1�al�8K���\�Ψ'�A��]	��	Ƚ��ۗjy�6��ؽ�^v�;��7�ýٟo-���x��-h���M^]�����Jv���fy��Arc��8�7�,�`;ܶ"Վpv�m�y��t��9���qb�zv�.�sd�z�oOem��V�O]gu��ls�Gg�K��9�(���
�� ]�&�=���К�囨��=���d��*���w6�밇h\���Na�pe0���p�.9އ�v8*���d۶�^�gĎ�շ�ru��qĎ�W�|�i �j��秛pR�:�ݝ�x��� ����lay���k��8ո����=��պWO��y�ޱ�e��-\�6�n��8�<E2�ؘz� =W[i7Z.,�^�m6�s�l��$�K�a�7;s�6��������n�����7�K�M�Fո'����7[��q;KsO/��Q�0��ю�N� g�w7e�4�������F�m��l�+l�@�]�.�n�\��WK�	_S����^R|ͭən�ݮ����$�౼����[c[O=�6�݇���l���ţgX4,��X��Om�L��n׆�J�[�[[5�VmG�����hx��p�ոzˮ:yW�og��4���W�������hl�u�]�.b�>*�ݸ)1wn{D�����<;�l�ث�bBu�>=ONn��q�nv��ˎ.��(�{uʏnN\8h���v�vf��b�7�a��65[�.L��]q��fk�Ps��3#��5[�NYx:�M��`�.���{4�$��lD4�d�vIj��j�$C���ȧV��-�Q���g��Zg2��=n�ΰ��M� ��������fZ����o��[ՠ���C�tI5�F����,���x���vË6��$.3	�y��;�ő���;����<��P'r�9=	ed���.n>E.�����y��4.�r:_t�r�$׏x�Ǉ�$����=��dH����n(F��ʍX�w�n�q���J
�:�A�!GQ�^[Z�X>~�r��'�!��@�����։��׽���������Y�Wjk"�KYb55�M ^2/�y�&��t�����kM�8�Ys�X��&�=�ƗA���Zj�~��{�_�'�;�ԥ�-�����m쏛�X�-��}���]��-~���m�\}�Z�|o_o�ԝM�_R7d��6꩖W67h�U�=�Q�Q�2�ZY�zn�z�q���-�u�޹5ƺs/[��k&�}yٝՕ�a��l���Rt���oTps���`��u�PC�����kx��=�P���Ow:�q
5�S��$U����>�e�<�٘���TF*�B@Z��y��8�%p�>�v�-ER��;Y���k9⧶��e��C��tGs�.�!�	�@����@��0�'	'D��=�ш��o����y��v^�N�C��&A�X.a�oH�ۉ �D�a�Go1�_Ec��ˆ�5�^���`8��C5�h�̈́�)�^I�/o"�{���DlM��b��}]r�!E�7f'9�+fr� ԮB���0�&xP��L4�$�*7m�j�s��ͻprF�S�5r����4��F��+���	B �mн��3���^��t��5�㗣u\m��3��ظ�)��;��0�¤�bG����^r�XV7
}!A�{�H��ﵪ6��p���	�
�X|�u������j�%�
\:���C�<��VB�&v�Ø�]��E��ѓ���
6H#�w5�D��w��a������g�:����1�^E(��ᤛ�w���.��۩���2en��X��ow8�����a������C��cx�}{c2� ��-�F�k4$�U�%�����M�� �d��V��D�%R�� ZF
l�O�6�ȈQ]��]YS���љ�c����0�W�C.f��Әe��!�ոj�d^��h��b�Υ��wuk|Q���6�h�,	޶�u{Is�
��V����0�|��.W�F���*M�"(�<�[t&=�(Q��gWrv)�\Z.���K��������n��Y��G�[l1$L�j�Z�Wa��i	�{Wi�ՄR�B��o�|���\S,|,�{�S]��&{��L��܊�F���.�S�#��$ p�J�ߋe��	���pcDS�=]|����6k���mC-r|��n91�c�DfgD����!�*<�M�	��s_��%%s&o��"��tp/�)�Ŝz�h���Nԍ�d�6���1*�8�I[Xk:aU��z5Lf�S��m@~|w�m)����r�k����G��lǋ9���r]h�[м�!�8�W��-�����ؕ��.�6޸������v_;4}Z4Qͣ�k@B��х����ޠx�}�Ћ��6V%���������q߈+�����ffr�OwX���ǵ:0A��7��p PG�Lș���(2�pKm�b�UY6*F�9\rmAFV�,�`zU���v1[��P�Y��n�Ԡ�'k�R7��fi��Ѓ=���9�Q�Ԡ�X���UNI�N]�����r9	#�<�\!t���k����Q�(0'5�m/��f���r��1���I�a�ɝ�^K�ڲ����f�3]y�y�;�`k^\���
�fpcP���NF�|���zw:��)�y\��qЭ��r?mnh��ŧ:��1.����w�;"�ә9�h꩎��S�l浚Ů�=ie�RI)0�~�l�k�'���i�β��Z��7�Ⴘ����s�����W���C�&�yi�+�+�	�ughD0KQ�Rg*��tr5҅QA�َ���U��0�7ʍ��=}\��;V�-.t��0�T;7L��}�t6Eu�)�V�rWkzP��+V1iZs�܊�3�l^�A&.��]v���[EN&��#|qM���Օ}���ݷ�{dy=|W+���^�����\�(W��t���Ϟ��Nkf���&5Զ��Z?®��L,�� ��c5:��%<[�n�Y��t���w&�5�2��[Yf�v�P�E������:����/2F7�ڧ�C�\V�W;t��cjM���N*[���+�@�⮝�/n�������xӞ5�<=��0�X���皷n8�쉻��oGgt��۝���Gn�|s��<R=�����S�h�V񺘫r�u۞�����惎�xxTސ���� �b��K��m�]���]�2tC.z"1.`���&�a������{&LN�6ۊ�s��S�.2؈
��
�J�v�g]o��&��jK�>ޭx3*#]+��k�q@C#�x?S
��g(�[��E<��ދ��;�P�D!�EAk��u�:/�۱k��Ke��C��uI���n�"�3K!d��m�9�"_6��[��I����gk^p
�r2V%��NqÞ�3Z�۝8܉��y��7�'^��i�F�O������Q������\�\u���nC�5v���:�}Zǻmf�c��c!+��ܚ�tr�aZ�����ؘ��M�Zͬ�3"���ś�+ڲ��kc���ʤڹ��=5�%B:�4�^�ꨚ��Q�<q��.A�ͷ�y�n�D��&��IN��\e��`"d黳�T�`���6� ��m�<�u�<z��x�v�
��[�>�Ս�̍������4��"#�(���Zwg:��*U�E3ʞ��BL$�w��S	<5ϻ;��2��oxln�J�~��Z�3���YAkrN�R��׵�;�YܵwPq�p����n/�]yPԚ�j`�z͆b�9؎<彙Z��6��90tD}�t�k�"Y��6Rw�' ҳ�`.�غs9���[k�ٱ�*�����NZ��u�2��Q2��.����b	����pfͮ�!�:�.��^j^��"�8`�ɪ�)ޠ�w;�#ݼ��M8sč���|���5*�?x�k�ڕ� ��Ú����k���aYA� [�K��}n���d�t���Z�,ɓ}�"7K�+�C��p"��F�����0��,�dmm�[]f!���YV���&۰E�.��l�N���ٹt��:��-	�T-�}KB��8>�Swo;p�ِ}�V1�RWf[��?s����ʻ/5�u��sh4�꧗�t��Q����仭��j��c��G\Id�m1�㛈f�]�dv���b��|�!���g.С�����+�E�z�\��v�*$�1��Vwa���a���e�Jl�vFfU�9)����~I��k�eVYz&QԱ�3qz&b�*޻B�!����@�Ъ0X���4_�^k�N=��e��;(i���}���>9F%{��^��=�Eࣽ�2�+@}���;�9���.��K^^S=�w���{[�ٔ/�t�)��^ћ�ܭ�c���{����,q.|I����z���V�fŊ�{Ȏu�3V�cK޼��yDI+�R 5�Ջ�wS{�5�e'uy��uᙻ�9�NrՌ�T��������rBP���N@�C��l����mx�jB+`XIAkj.�:�;��y�(ǾrM�,Cf{<2�}@漰{�Ȏ�Je���lG;93}��-uqZ��e��y��u�bM�=V �B�JL�َ�p�nݶEΎ8-���ָ��lx-��#�ӛ�>�<%�Id���ڵLy��q���gv٫޽(��{~V��G�A����]���h��뛍�ÅP����,�*�G6�@�_�JQ�D�R�ڋ �/������=�fM�A�������a¯��2ap���c�M�A?,�-���$EP�7jI6T4�0�f�W��L��X�Z���N^��l�Pn�JV�W� l�؆�����t�o^	�Q52����\h�Y��!�;�}F��owZz��7:�?[+���}�R�6G5]��]�*�\�b ��v�ax�lG�؜;;LN��YǭKJ���6�N��k�.!�j�f�w`����i!6���'��Y�G,c������ݻ[��5�{F�v�e��nn�+�XQ؆�	*$ҔOv�Q ��t��<z!լ=K����fjج̒*�R�N�����.r��=4Wk	q:�:�
��I��pf�`���M�X�\hvlY�ޜW86����+X�k����;�U�xUj{5�_[��5�\�s0�(����φI�e���s4N]���]e�~��T�Cg��MH�-"�7n���J�:���y��WY�q)]Ҿ��3kh��AB��1D���)��n�'��o:5ʾ�r>�s�5�
Z�t���7y̙S�.�9؋�K��H��(�
!m��L��EӜ���8|��<����ݑ�nuU�I#g0��	�8���^�F��y��6i��z�{��-X��=�gvK���vOiX�"��;��Ih`	D�&s�P�������E$��%�#M�9��LJ:>/�Jݡ�~l=�7Ԕ��f��9��(�z㆏ ���C5����8.�C�y�v�ߢ��q�֭�Ĳ���VY1���#r[�Q��t�%h9CB��ӺH�)w��^$����A�{1�*�>�/woM���wq�Wݿ[Fv̽Rs�4��	q�d�	�7*�s���u����
�PhnxyTh��:��7f�on��dی�ɘ�i驼A	z+'t[���gGku��*���;�7��qM���@f��w��؂~rA9�4tM��3u�0��;�k6��y�M�eޢy���ܼE���&�j��v_4�O�F�X�+�	����t=��A��F�&�uu؝j1��M:5�&�+����tkt��5��=��\ujv�Ux�ձNs��٦rb����2��ܴ���n�~���YŹ)'\���Y�N���|��}�y�
� ����V��r�Wr9ꯪi��%�pؽ�)ٙ8�C��3��j����M@�M}���T�D����5��+[��F���U(�بd;���3����:����#P����Ȝ���դ��)�"⧫�����J�k�ܲr>Y�X�I�R�td.G���ɋ�/�<83Z#�M���
l�o	�Up�;^y]:�����)�V�݁'WObמ��R��=�M�S/�1�\��ꃍ�����t=��U���7Qf��vm�?I6G)+(I�[=/}�B�DZ�n���U�����s����,GVlB�a�5I!L�P�9�L��GW�[a4�f��*�Z��+���x�m:�2�����\7LR��z��mVÀF1ì���3�<^^,X>�Um\���m�WhR�w2Y���֮w~��=�ʏ�������RDsNvj'�J�x_�s����9��a�S��E��Ƒ	�[w����+O��9J����vqQv���>o���1����ν2�[�o,���|z��U���^s��pnw���#݁d{s4���PV�/�]�a�a�+�HZ�Wy3��ﾥ�z�pbD�$*��c�;�z/��T�W/���(9���s�	�x�Ǧ{pe�T���너�	L$[f-���N�U��\yB�
��VYF<�X�/�H]�[	��sO�* wmr�tj�H��������Ή�J��p��Ȯ�ѕ(�+���{Z�۷�Ge�1L�S�j:!�9
���f��?$%�z�dTd!ـ�ix
�q![�1uB	�%A�V:�s�u< �'�d��t��kX�x���։Ke�v�U�	G����u�U��^ҙE�s��P��	��{Z�ڈq���/����瞘����kC=�p�T{���+=]��ZY,��4;���ռ$����W'�һ��Q��Ć.@8�{�y�	#i����<���6���x�ٵ8�Rn�p�i�N�6�����X�{ؼ�˗��Pgo�Ѐ=tu�U��1�.��P�ֳ�-l�SC"��~��'k�\�z���<��n�o`oM��P���Y�r�f��]&Q�w��Y2��N�г�R��ͣt� ������	\�� �Y��m��ץ:/s���)��/;������,M�Xn�UxUk�4�pQ4�7��H�n��r��Zi��\4��շ���8���zh.Jݮ�$���>�Sa�X����V� .�%��c�:��۸e�����f��$]<K,��2YRy͈���{��P�e��eN��݆���xj�������j�E��]�n_8��
��DB�5oT�g3���G@��Cs;���`-n��6�و�2q����7D���u�i��WppQ�ٶ��`f-8�=�\�]�����.r���F�t\΢/��$YlAR�k��;�u�٬�z�X�Y-o���3�y��r�����؈�D]�*"��Y�4���K�NX��.S�)�{��)v�e��F��̍��o;��]K���}{���yp�+5�w4�6mF7K����v�����l�:�)��wB1��r�5��os��vi��w>�;��G>6NN���̖Q������ާ.U��m�}b=2T6�\�����X�e��d9������Ԏ��]*�0VV�	�����MLm_�z�G:Lwi%��7�N|2]sy�jqƬw�e�}yʻ
f
5�-ߐ}\5����1}۸���rn����Ɏ���+��:��̴����浊â�\�nE�⛧C�#2NT=���:q���-�}���g�ۑ����i,Ͷ�FwM����`ߍ]�e�M'&TNی�{X5��G�$���z�:�8�t\��Z]�{�Z������l�
�)u�e�p�I�ܷ���,�����Q<���C*���Sד�����M9��7kY�Ns*Ȍ�A�[Z-W�A)e�
��LX�K��9VƬ9������� �]c*���:�B��6#�ֳ{?~�-��o�g�o��0�yxK���w���v�#ϥ��7�V��D��P�`��KJ�II�07�{KZn,�߹�j����v�6����r�v�*"by�Ҋ�&�m�\T�"�y���kNﱗ/���+�ȋe�Z����5�g�7���a�}n6���>&���"L�i��_cZ�W�HZb=���a	��`(�� );�����p�p_z��+0�Q-�(�=��S�j��.%�T��NB�����!LGٝӳ0�~�@���7�d�G�D�H�9p���Eb�duKV&y�A]�6m�p��z�}�&�E�6��KX�Jͽ6����v�JX萪�m�4M"�HZN�ő��ˋ�d��N�[��,1>���B�f�6��
<F�rF�E!����˨�T��\ˢ�Ғ��W�_D)�%�޼�!i��M�S�SW��~3|C`g�opO���>#�,���iUz�l(Y\�Y��2���9�����|B�D��"TnU�(��~F�Kb҈h	�F!������kۮ�ĭv}Jәέ��9��t����]i�muj�i5�|H� A�V�D�fHETfw�K�8xJ�R�DH�T����~5Rq� ��RG����d�&�4[���N��6�
<d�Ȓ ���ΝrN�`��8�T�����&O}�CR�)�%UKuJ��ֳXX�0��2@���'����Pz![���T�m���ڛ��8RG�|p��g�y�AF-40�n;2A"���#�/a��9k"��a�l��������k,v���\\m��_H��"I��"��y���t�/�[�h�2P^uY?*P4�Ǚh�+뿾�Q4B�A��Hp�}}�b~>�ɺ�T@}^�b>����=?qZ��mx_о��
��c�!]��o��M��!Ӛ���&z�TT�\��d�u��#�>i��u׆tǑ�kH�(���{5��}�� *:P�AeV� /w=��E�L�#>�$�s���q�?.GH���2��� A5us��ǘ�BH�(�wy˟�*[MU9���Ȏ
�BTf�"�Gy3�{3��5_��!��	y^}�L��mg�3(H�:#�O��X��y<�s����_R8�q�ע��M��[�]\�丑K~鿌}93?F����kv����s4,	+�<Ѫ�u�o��Ca�tm�+e�e�z�-m��V,��N�5/55ǜ���׭9��(J�(T_��at=��<��v�wi����5�k9�L;�ל{:{v콻�ul��\�y��6�^��r��u����#
�&�Ź�q/Y�y؎�z�n���m�w(�/k��	c��k��v�����g�7\vtf�^k�G/�#v�3φrv�l�ԝ�U���7\@��p�;]��:����[���Y�n� (�ul�<]�;_VRnƑ��]���[��B��vwZ���-.8r/'KmJ0QT-l������ގ�H(������K>y����p����)�	�J���d.q���	�J@�4���<�8yo�w���I	���ۤt�=�Z^F�h[�*!H�Ev��}I�r���MU<JM4X+!Qc�[���ߪ�`�����/��bV/y8WdH_V�x��ӻ �xI���� #V��j���|}^���X@���ۜ�u���`�5�?}�V�I!Ҝ��0uS�8)+�v�+2�W�S�̛b�L㍷
�BR'�)V}�����s�`/ZJ}RR�8ZB�W�w�q�	� �+��-��+��M���aG�2�����|8g�`@��,$Rh�SΉp@
H�I�{�uJ�5�W#N	r�Ϲ�v&#Z�$]#�劺,������j����O���ϙ�A%�n�v|�
8C>dQq�Eݏ�*>�{;V����q�N:�L�[V�4��y�\��QU�V�Q��\h��mX����
EV��x����p���5G��K2�m�m���c'��j�>���~}�#�n'���6D��r�8G�c>��E���=�w�j����G�ǝJL�=-�es���o�Ku�	��)�f���\�J�y-�ٝ&��41[NyN�d8��8�AԕNh	N�!�3G�Y�9-z�/�N	9v)���\�--pS��kH�a~�=Y� ,JN���Ր������/�">��rn��*) Ͼ)}O_wۅ���
�%��*,�����YE%����s�5��H�L@e�}�}DY�>#��9�t\r�������\�y��F�P̔�hRn�oz�B���V��_+E�n�k2U�u�����o"B�^8Y�e���u���]X�����y����� ��³�g�3������
�̔�_~�����H�ˈ͏��?�F�@��1�?c�F��ž���aEmR��ˍ"ܐ���)w����|�s�!p^��/�m��C��}�/�V2��~�J�����LS�[L_^o�k��l:ҳ�.�bTC���pɎBU������(�G��~��ЇŬQ�[G�>'���|�/7���s�8��C��-x\St-n���d�6 ����}��M�#�|E)�;鴤�) L ������_9�o�x}9�$nr$i��-ɳ�q�Bφ\؎~p�i��'T1�-RG���ڳD�Z�aM4�˓�}�|�gČ�NS"��T�ٮm����+��M����J��A ��z��}�@�Z��9� p�gJG��^L�CZ�bTGzՔ,s��w|>Y�)p�&�l	���b���q�;7qRY]5s.��lF'qz�[���
�F��v�<��}�m�����-.�vm*4����ʠ�����W���W1����MXSI�x_�_ �B��.DN�ٲ|,��z#���DY��o@���B�ܒ@7��֖f��ף�@T��@.���Wǘ��D�F�c_
7���!� �|�}g���5�d�Q�������
D��*(92��׽8�|����һk�>:i&�=�pŜtE�?���??�N�mJ��)��`&��S&�S%*�����x�!H��U�u��k1�h���	x|���d����׈܀�$�pt�¾����k�W�X�f�Ma���"�����-h�b;�u��3Y��nfw[!��f�Mh[��6�UHn�鬊Q{�bH$�R�>mD�jw�M�͡2$�VO�c��_5Z��8/��jH�1�H\�y�ɝ���Jh�������D��	5����c��4�9;}�,��du�M@r�mF�E�8}Q������>$�I(�x\��'�@=�Б���=�(�Ő$�O}��Ϻ���w��C��y�df�Ym�C#j�6��:�7?�V"�THZȳ�ID�ƍ�$Q���r�34)!^�K-��=����y���3����$T �0�m�]�j����ְ����Q~�{��|ؾ%ô��Y��R��t�wC��=7��05~�'N�dy'krF�CG����Gn��[ݐ�Z�2T]V���6T)�(y*���Ə��q�Y�Sv'®}�2��m}��K��}3�z(Q��Y�2��fdQ��>��)����Ef���0���.Z��;"EW��Z�4�D��9hF�>�{Fk�e���	�C%��I�Lt�%�>��w/*�WgԬiqWc(c�܏��UZ߈��״���#vK}μ6�x3�B�<(�EL=��#��e�t�(�(d,�����5��9�Z���-#��8�Z��k��`���3�dQ��; (�&�T�{����KZ��q����
6|n"M��Z���Qo��.#����k�|!Y��JȑӱW�u�zZ���b-Е
�$d.��}Az�?PP&JM�����]0O��w��Q�/�B>�2�kT���c�|}���z���+6����}Q�C�`J�s��KR��ir�Fv��g��筬W����g�+��o.��ln�l�]���\��G����:�uZ;�����(�MM��sG�tˬnY���/�_j��8I�R;��f�fض�M����Ϳ����j�,x�O�%�:�^'�_p�E�b"�n���n_�VO�d���$��Y�n����aMZ@�{70Gu��
6|7��}p�(�9�eZ�F /'�q(���UG�]8��\F����S�b�`&C���8[u�k�Ƕɞ|wm�c�p:���q�cG!����M�!XA�PY(���������4����;��w�1$�M8�\Dv��Uq�i
������K�v�����O�GdA	@g��Ad�;~1o��:.�)�2(L:��dP�s�_9���$���Tѫ���FB���&Q�������C�Z���S��/׽^<\0�J*܁��l� ��\��a�/���昲��*���|i�!�����$5�g�"ϴ�}f/G{v9�k�|r,iW��Sc��E#L ��7��آ�*�ʸ�%���覟�l�f��FT#E;��7�'ә�'������w����k���">�cK����%�̧d1+\��p��{ݬ�E&��ʪ#�e�_�PB=�o�Ԗp����2.�ϭW����X�I�ܣ�j�یn=�����
}d}1��s
���k�Ϋ��3�P��j��d1P�A4���X�����+9���I����	]������f&��Wđ�蹝���+��w��>���8[X8���d���GU�5_�!08�d�����A�q�G���e�Y�V;�L�r~�\��}?:��di��[��
M��-����E�I��@S�.ڢ=�sŇ֟���D��#�bg��"��|7�)W[��v�ZӪ�&�m��8�bBV���$Yر.:�V�VE���Ȫ��������5�|�W�o+�F�gjQ�����M o�������3�a�@�m��p�[�̀����9:�e����������c�ۍ�k�t��,��y���8��M���q�Z�cB�QES^��q�)$��+I�9�D�5N�ѽ\��,<6l�@x�h�	Z��GE��;���mWZ�^���-9���Kb�v^ڀ��������lc���-k]�ܺ���ݺۅPN�탙��&5�k��;���l<!ʷ7g=���srkC.�ப�:�j�I{k��4���f�l�J�U��кE�����,�bk���>�/���D�g�G\�"��UV�A��J���w.6�G��qZ��e��㧷�s��@�ߛJ�g36��Oy�-}.'ZXe8���ɕ�A���ʙm�6؊R�f�ap�6�D�y��UW�������F�cb%hq��>S��*<"jW۷�ң�)#��ȑ|�� Κ�/� f���}��h�".	D0p��}V�n�N�sϻ����/�ǅd)�h'�UN*�N�.\ӵ"!I	��e?�i>�|�@ZC��e3��.���ۛ�5�q4͖�ʖm����_hD�:DLv��H:��x�p��Q>� }qq{t��̖}�I�(�����.�n���_���Pn�i �+�$A�����A�9T����|\��8��}ٸ�]OSE�%u��Dd����Ր�Z_"�����[�Jn��N,i>@�d)�#�g�6�^yR����>��R
�(�w)�(����KH���V@�\u�M~����,��3� -�����#��l�>��i�
�w�(����z�zT����aQ�0�ad %��b��7����X}W �����Hm��6E��-�+ׅB�qf���NUZ��V3��4`ʘE�����N�+Gi0����uk�u�Mύj�WuWP�曅�k���t^T�Pāt�|����h���EC-��I�*�rk_{��ii�8L�I����g>��<�M�~�H�^	&�וw�GD�uE�IE���,�wܫ[��T >���R�=mX��W=�^  A
Qи���{X��Z|rl�0	���Ƽ� �Ø����W�	�[��:�A��Ph�c$�AgaEnh�f��!c`F�;P3B�ذ��ij��;PTTtu�\^�8�U��z/o;�3j��HG�O>�F����DDE�	>1���W*�{�O. j�����08�Ǳ������xk���c韻�u�����`��|c���SnhR5N�d�u�V��J�4�!?y����u��dq}���S��}�*�`�B��.\�>q��^�}V�_�_��A�|+$K}�ⵢ��ĳ�*��.c]ְ�x7oʕ�J%�M�Z�G_�n8T��,w�:h�jo&�C\l�$�N?W�M9���f,��P�a�L �����N'��E�M����Nb�������"υ	���F@�nx3�LϪd�0)I5U7Ũ�֓����Y�s��������	�T���|�1�7�/$ϸ�Ε$Y��� �=DmV���i³�%�՚I�N����Z��{ id�^�����U�K�ߊ�*L"i6���k6竺W6;WbN6@�T��������#-r��d�j��vP�U�5���X�@j"��g{<��R��82k�@*��$�*�����M� �q��$�57�)�9�����}=Eћ�|d��H�hJ���.�3�v�2�Ik��S�my�:)A�ZIk�V�g��(r�+��+Ə��ò���8���H]!4.{{Q�5��}�l!QA@�p�{}V�ん���bZF�:p�{٫���Tw�q��S�)����v�9���@�G3UxG�:�>	�^DQ�w}�|8��5(�!TI�G���������F��������`��aћ���bgr��M]�0uO{�&���[�)]���\��25��t�l�-*�r����j6�����FG�3~�3q�W/�h'���L]X=!z�xZ�1)H��Jםz/��`IEP�@��dg�(�)�;��ڿ���Ϗ���t�μ�"1|l��2|�8�C��N�FL}�ȉ8Q4��"H&�ܠ+��V�|�ܘ��X��sܣ���wU�:���a�Y��"H��8j���X;h8F*|�X��\�MI'�>P"Ϲ��#���te�}dUG��"��}�O�K��c:�n���e��T-�>�Қ~�]#�T%�EW>�+���Ws
���AM1U���i���=�ꮨ�܎��M
A]��Ӈ�����K�<3���5Ŏ�"1!N ~](�NO�,�����x��|x}1�.cTh�q�g.}W
����-�.Z�)*��I/��rY�ًE�+:#��;?(��~gqdY���h��h����f* $A��!��!��JjIeR��M<�x��4H��$؃�y9�UƁ�{۝'>��o���2f��<{���	.wj��O2Y�i����Y�q�QÈH��Y���ӢD���1�,f�ׇ>���eL�����&�~ߚ�$�=%�����I�8/]�-QO���G���!p_f)8a�fA2�!�����Y������p�z̬zO��o�x���"g��rs�	��@%�Q.=�k����&�܂	���d�C��kU~%P��� �{�J�
	U������Q�Vخ�"n<�m� 3��q��&ƌ� �R`���� 0^;lB�@*�+�����H�
g�rc��jY�!�cl��9�w�OO�p�ѥmѰ-�gv�%b��:�9w�	�#*3�P��ֹe&n��2��o��n@'O��[���{#���E�1i,dV�HZVT,K�|�<k�w�i�nH���vn��jA.m�-����@�Sȟ�=V� 7{ۅ�&$�~h���t4|+�@Q�?i�#O��4h��#��Ïp�D B[�RҟS_�ɶvv�X}$�,d����q�:�4k7�cq'\s���MT�\�G2B �J���S�<�k�an�#�+P�l�յ|_8��k�8�B�.<I�˩��H�L�F�|�62 &�*� '��t��#9��罵{�`�}zG��&}��-w�_ֆ�B҄���Չc��
���@4���S�۞z/�|`�3�N�iT����Ѭɽ<u�U}�G��~�~}DM�(�?��j�Kȉ:d�Hg��\�D��N�i�.La�4���x;q�߻6�8�|��ܷ��~�/3x�3�$y��=k�=s2�u*Z�Ej~�H��[ZAo�e�]�W��|.��3���zB�e���g��N�v\�x�p��^N�~��÷��O_��	>��"io9'��X}I?n�>��,��Ʋ>Ww�k%���F�(VG�?1�&��� �&���|(�1�!a����T�j���l�H{%�O��L��"$IKVEw��\-c[O��#���Y�I�%�r�	�$�C6�߰ n��b�i����w�iZ��]"~Ʌ6غ*!s}�J��S%K���j���8ܶ�B�� |.�� i��k#��A$,d�MH���Y��<��NG@���n7�Lfc�x���V��	���IߧO���0�H��W�ʋ ��=��>"MJ&�%���,���*s:�U�;����oVm�K��%� T�]2���p��*��Rͬ���ї(�յ�v����9��u�)�v>����U����j7t�#JnWS��wE�Wi}��.�R!F�*��k]�nŗW t�@��tӫSg	:NwUgJ7��o3y��'�^��(oW,딣=��n�z�-t��k��7�����>��N��8N��֞�ȗת�pl�j6���	%i� �Hb�w�V>ް�YD��w�v+q����G}+������WH�.��k�g�>��{MڊI��ۜ.�0�K�e禝e�|*o`fa��}�6�����;�Gvk�R���Jn���x�K;� *�d�],*�JW/�V��쬎P�J��$���ze�ur�x�Q�ŗH[��V�bc���w>w������%zn:٥ql�ˏ��,R<  ������l�&�b��6�G6!��ت��jg�d��)������V\U��VN\@9��V�n��sV"��������}}�%^�sFﻷL�1�5;se<�UR��-F��d�f]DFQ���Y.�ςJՙWγ]lї1��l�М��SN�E7:�v�4U�5Цi}�ZB[)ܻ�֜��K�{�7	�&`�w�fu��59e���k�K�(q��ÞK���g4୾�Ŝ��[$b��B���st�ͺ��E۾����}͈�dܤ��/�밸�c�$ͱ�f�ZyX��(����^��9��m��(۬iǷ6o��w;�k�@�'���"���T�Bu�hܛsn����3X���+��t�7@9�?�mp}۫�c4HS���g�s �<��b�u������8�u�v���q�6�c��7Lnq�'<��;i\���5��T�@ӡJIݫ.���l�v�ݬ�ƽ6_m��:��%�%A���n5�����ۧ��7D�v�ce:���mv�w ��G����ێ�ۚ���^�6��肘���}�n>�|��8oZ����i-��2���#.�ح��4�teq�z�	>�͵�Ϸ<�����+�kv�]on�N�9{v�{xn�P����'Ry�݀�==�݃�sq�l�=ۗ��&w	�ݑ��N9��ώ�����5�p�Y䚌�����=�q#qc���ΐ&ݽ�5�n���X]��ps�3���b{v�k���maÎ�¬l�j��eHO�N�:9��7`�s�e7s�(�Ó�92N�Ի#����Z���:0Y�.�S��r�7kq�n
�����;3���l�z�mg����:����uYS5�6P�+\���a�/[��p��'Z��l�6.�7:�ԏ;������06�M����[vη<���y<q�����q�6��e{xx��c�v��iݑ��G��=�'W<9�!�m=F8�jɒ�ɓrnuv�ukm���i�􁻫�(���z����<��[;��W\jݖ:���M��sڷ���[e�On��R͌�4wG���/C�f��2$��D��RY��h����d]�U�)�v��4.�n�x��NC�8T� vK�F�u�!�^v�j���/J@i�ܥ#���9����9s2���vK��r�7'��s�g��V;�vh㓧�k��|��30�.b�<��m���U��<�x� Sѷ�Wk[*T�S��ا�q^��[��m������'�ϮBy��^x^�ez�\v^��4t]��p�W9v�)ͱ�a�(�:�;���Ӟ��e��z��۶�=����Fn�R㳎.�u��q�n��N��'aںOg�q�o&� v퇴l�u�н�������Kg��Gnպڒ����6�l�8+n����r��`��n��Wg8���=�;�{C��un6G�p<#�`�vz��;)�d���&��F�P�ƪ�N�=��ư9�c�.6�w��n�=n�9����;rnm���Vqv�Q��w��<}��?��y=	��nv���뱳��u�:�����:����6S&�n_n]�u�u�ݓu���s�������ƍg��t�v��D(�+�d;��aF��:70<�=��>Ƿ�,4�}b��²Q��+"O��ɵ���$
!�ʜ*���i���{,JD6HG��꧷��`�_A��ţp���F� ����Na�dĉQ�x5��oO�t��;������.%z�qD�����[JC�.��3D�L���]W�ǐ>�� V�|�����U�A�ב�'�ETzH�H�wʀ�����,0�m_�T�Wy͛E58��Ư�{����{�)?8D��Qi6Z
�T����D�����D�
�>��v.FO��a`Ez��ҍ7{S#�m��@&z0��A�~Ϣ���}�x��ǎ�	��r$���>�(��
ih=�S�_]��]GD]�u�����^��r{#ck�Rښ���SU��p��Ցb�.w�O���'�r>:�#�)���Y�<G)��A�뀋�(��Yɸ^��[A�TE
��2,'�\��>U������w�OZ:B#vt����S�0�q��0�-��̮AU$�ML�gM�D��b�>_J�xI$s�ﾯM��q5��_�2'�1M��[&�}܍����F��pTFթL���0��}<�_6�HX)"E�
i�#_}��{��a|dUR�dQ�P��>�o�|_�" ,i�B�1(݈|�mJ;llc�m�<琺�y٣)p[��ʹpuKSr:��-�����ge�%J^{}�7��;n&�L��bT-�ʳ�^�x����T���j�U�4�Q���x�|��y��o�VYC���-��թ�&:��X��H�������T�1B"j�w�o�P���Q�U�ߔ�a+VVHLWD�ˊ��;�1!A� �3--[dNȼ�q�I�����o{��t,}YL�=�Ѧ���#u��N���p���ul̊�C���#� ��0������&uY'�P�}�R~�W ]�O�r��*����Q ����i�G� Gg�>��� I	,�'�y��Jl�1�����\c��߄n|�ƑMP�P�ӻW� �fvlXB�rP��0m?�{�p��ʅ�����W��ﯯA�f�aY�v�� MU<:}f"'�ϲ��]��;U�P�-	��n��x�!O~�Mr�n�EeVP���\k��K�@��EF|���Q����p�F=�I�D"/�_��M_��ׅɏq�ݕ�RY��a��s��Z������|���crk� K��r#c���������E�"U�5��*8J|��P��B�$R+"�}������q��?E1�.o�w}�G�NZ��"�����6Y��p� #E( Ү	,Y�0�8��t�	{/>�\��� �u�d�e�EP�Df1����wE�J;����r��-Dy��'���qkn��q�|y��s�R�V���Y�(^����Rc��"Ec��%=~ݯ;��옲d�Ɗ�,��Y�E�U�4���$�-�.h������o�:������<�|8Xn4��4t�J"�üV��$a����ybdm��1�����s4�0���G��Z���\�p(�W�n9�	Dk��_��"k�t}����P�2Nz�Qy�okÄ0�DbJʓG�/�VG�X�(����ȱ�I�	0��M�|��p�i��:�����w��z�	Ǆ\��q	�Pu-T9sU��5�B�I!�u�e��}�ϕ>�C�o�|>Q���|hU	�ܬl��>߁ߌe}��>���qa;ͭq"�h��i�<bLk��T���iٻ�ަ*�ȳ�{'5ŗ#4��B�����#�Wُ��m�� �{qT0������gz��lLy��8G��lƁ���A
�w�:��&���L�V��� �<�J-���9��WǾ�W���/�串�7,H �w�NBњC#E	:|���=���0i�0�>. ������goHV�⑱+��/���`��ީ�8|7G�D�7��0��Y����ܕc�J��
 5�*�� |ccK�É VZ����pҝU~�϶��z �d�����ɘߟ�>ݫJ�
HLZ>9&����լ�8*(�|�9��X/��s<g�쫾��y6ӕ55
�zrun'�M�����$I&��z��J�#{]�:a�Qh�7D(�/��Q�CU��{	p`����a�A� A�
Zd
ڟ�?^�Z���e��*2I�dz�������x�ۀ�!����K��X-G����� ���T"���_+�����ıL�Y.a�UT�j@�g�Bq�3�TAD]��3�S�ﻖ)�|�>ܕ$P�y=�<�/�OҾ"HU5,��eJS��M� (JM�"{4��}}�͆cLӇ��c�$�&GG3����,�÷��&z�&S%MT�.Bє& �9��$�0Ͼ��K�P���F�RE!�g�9�8RG��F��l�E�D)%���/=�f�"�D�!1*X��/����y�	'�0��
E��Ov�>p����`�!k妢|_����W��f��濾�����p�)g���,�yQ�羛��}년x�mȄ����^��@ftC ���Z�f�*��o
�O#�2���gq���Y͙m�ȁ
�)R��ԫA]����FEz2��F���&+�̧lwM�r�u0���u.�tzFPYl���m����b��$x�wf2��"A<�����4T�:B���_-q�V�酚"�∃�f)�p�P���
�d+������0�� ��tWd��,��	F) ��\痾W�� "O	M?���p��2�׷�*$"�"�G�P7b�D#����4}{P>@���q\lA�v�^R�v�k��R�ѩVM��K�oWi�ܫ?����9�E�(�rR����n��)`��1-�n�"�M����ڲ�8RH�I
�Ɉ��U�*;b~qqZ}�i-��A�G�y�}�S;�*s�	��/�MhҊ+K����|z,cO!�("$�$�D������+����'�YȀ>5R�EA{c/�#Q��8�*f�YhJ�����}7���B�. ـ,�|��"����:i]�,�c�Wݼ|M�l@dQ�
b��u&�jfU)�TR�f�D�B%�X+p����|.�������'�ٞ��χ}�q�T"�)�f��G��uY�D��>8��F�"�u�t����A��PF�ZH���$ZAl(Jϻ9�!��:�T��Ju4��"ﲰ�����_��?]�/����A����7:���bM{*� �v��'#��CR,��Q�a�'��?a�7�@�_=#�-Ő�L���H:�ȳ�^)�ۏ�2�pV.�Zx(r��*��5U�HL����kD7��=7�'i��
H�{���1^�}����߃#���te6�(�P��ޛR � ;����8>��p�����cq�a��&ĜG�	Ğ>x'c���WG}�䥊7�����[��F��\t�r+^;X�������ᕜ�f+p]*�ڱ���&��^��Q��<����IeL4i}�{�9sߞ��ɫB�y��K�xǱx�㝵�-�*u�whnkv��ۺ���H�Y'u��ca�>؁�h5nh@�۷s��ݮ�s�_O;�g89�H���ڎ:3a��ܸx�nj. �n�5a��Ҿu�r
p�{��Ǫuc�4s4s�-�l��ۤ;�}}.�mM���`m�kN7ܯ�v��68޻���]��%zY��ޡۜ�-n-ہ�;^�ٙg��C�/i7l�ۖ�%��qc�ϝ��ob��~/�<E
���q��/~�и�a����w�`&F]��6��o��DL{�|�Gt.�5�u�^�-�ޑ�GN6�m���}��&�j��P��� ��=h�%8*��Vߚ*]'$�I�8'�́`E���D�yg�:�	�$dt�vnGֹ������W~��׼Ԛ��$^�B�)����U���b^0�q�Ȣ�恧���a�?JD�J$�Tn�wL��U�ߧ'��&G(�Ĺ?g{i��	�E �!�y���"��8�e�F��C~>s�dfǙ�A�0h�B/���>���TWk�/zi���g˾p�Q{�>3�3��>DIހǠ�h�L�#�������s
�4�j�W�����Q@MU1�*j��������z�o��s߯���8kk�8�l��jH���g�oZF�fO�e�[mRt�N�o�w�? ��֬E��{�� �^�?w
�!D	�s�6@Yp�5��\�-i�o�,�`�m�+��xY�m�p=�0��LQ�5�~�"��|G�#�s�P��ђ0iu�N|4��G�yđJ=Fw9�u�7��5�b��\ԃxa&W~����B�G��Q,ۤ�p(Lu�k�?_s���O
��WDj�8ӠKSr42�E��=:�{i�Uיwa��K�@._@[\��uAdP�PT'~[k���g�~��zymQ5;m�u�d$��g��}��_�l��/�b�>T���@��}"���9�l�1xi�x;�ڏ@��:��8��p}�G��>!�&
MQ�J�z~n��]��),$���H��~�Mu��l�������۫^��M;�?��Ի5���8w���R?������D���#�u݃,�KI�[�A��@� ���Z��q�������4��L`ЁN��jرS�$���N��)@�}^y�M��<���ZhSU���{w�Y�R�}+y��y��KΧ� 8&�
��o%?�X��LӪ���'AM1
�o�����ޜXi��8��g���-,mk�*�]�����L1w�=���Q5�|�a�D��ﳘ�0�=-
�p0����ϩ� '�ݜ�O��h �/j�@~���0-�\���J�VP�i=��.�V}}�Oü��X�G*y:WK�h����h �r�R2��bʮ�n0F��]�Q@E?�SBh;���:pJJ;�@[�$����x�iz���5���$��&[�o�צ�"z�����T�v�Y7���h8ذVD�C���:�_��Y[G�����HY�6|A����=�ֹ ��ɮ��#�:H�7�b>Ϗ]�	�7�T39�N` 7�A���*�Lo�U�z�{�#��%� %�6~�XB=�;>��X��婒O��sƎ�yz	ƪC\�u��'6�n�շj�p���:"�92l��+_��kH<�[b��(�2	�{����jJ�LZ�IBu�������.H�P&X�!���D��Yk\�>��M�)�_���� c�B�ݿ}7�fې��	�� 
���Yov6�{��I��#%���C�c^~���	�m�@�-����rm,4�����k�'���$�6Qw~�31�=���1
O6�`����>f��q�0h�-�}i<��Cn��{���w�C���ț�r��?W���t#��B%���S[!5�8�5W�#��� �� ��5�����O�l���xr��J���Q�YV%"�s ��Na;�R�Y��!t���.�ٰ���Q�V��t`�����_sv���:�����mn`��;J��H8�=�2�ِ�R�n&�@ystm�g�Ԓ>��`�ٛV��]���`�cm��WMs����{�e߫����Y.@�H��(V�pT�?KsNfj
%�9��!^5��R���ۖm3�)b2�V@. �^S^��q��'�2#�=ii6�����q�z�&�(��M�΍�{&��Y��>rtm&Y���ڄG(T/�쏫�nywT@$�O9�5Z��(|jI�4-�D	�����~E��B�}
@��kqv�>cb<՜֗u�4�:~�j��߲b��U�IH��k]s��q�Vo���#�b]�xV)"�Ɨ�珕� ڻ��b���ʐ,L�2��Q���7�����1XЁ؀D�D�Md�~���u��湛^���0
M �#��֗�n�=�`���At�=eNj�ޝ�q�;b�t�ESS�y��
i��)�DI"�����x@��ܴ�@ vg)�`N���Y��E���%t�9h���$���W��g]��h[����#�sE��|Z�V綳��%q�d0>�=k��Ƃ;Xqrf_�L�n]'5S���"�k
+> +����e�x>�TA�A�f��?��|G�m3e�DT�b�E�
��0�1{氡��e��~�2�3�2(k���a#!�ՙ�j�֜^���ʽ��rĥ6�K@�>hX�rq_�V�%��7㉮�A�� ��B�Ь[����\�%n����.0lU�U����>�j8����B��?%^�:@˅؄���f�	���"Nk�l]�{��6 Y~��ZȮ� ���giq����i�6��v����ll���m��j�	X�y��%b�-g;�_H��5d�ng�dm8Sl��=��ͮ {�Hvظ+�lϲeP�~�5Z��>�!E�!�l��n�����nCҮ�3wb��Zh���V���iM�:л-��5 A��gM�HN�skͷc^
�{q74NG}�0�MK�u�@h��T�M	�&�1>{ͱ�UU Q[-pm�����=4���ȑ�8��Gיj�+ Y� �\x">��V}|�x�U�	�'�2A2I�3H���yY괾GM0��e�pTQ���_��զ0oE���Bdn�J�pѧ��;�F��\v�$����{4��6�� r ��]��c������N{�.�[\+)+��`�`�^֗Z�ziۄ�藭��vӿt���H��)h�������^�D
F$)pЉ}���	��*� �L�����pLA"M���/�}9I�1fFO��ó�fjP"�ύe�Rp�nj�KCD�%����H���f�F�E�>=ų~�c��c��8;�I�Bs��+�Z�I�|�PB�k6����uh��X�Ji����Ƭ���q�
~'���1G��
��y��rg��r�u4�QJ�K%��:��o�hk$�����~���eZX5�2��{�Z��_�%DD�Ҫ��pƑ �Fm�+��uV�w�x�裯d>�$�Gp�
��BK��-<�G�QI�jk?of��pT1.A��@�nE˞�r���|s�T���.fjj���� XE��1� �(��A����}ʨ��.p����CƧ>�Z��v�v�||�����wڤS`��%P����ir����)�Sg�cG��٦�	�� ����7� NL�|�:�vGd	���Q�'?YT#����:K��4:�jH��+iX�G�1f��֓.�x�Г(h��z�����E�����$Ih|�$L
>Uv��Y�7&~�"���	�Rt�҆���M��%?U�1X���!�ZQ�u~^���RRb��\�+j��*l%�(!��.���Ϩ]� 1�l�5ֱ��&>�	����Hq�tYYߚ��c1�ڽ�Z�^B����vCv�.�y�e6h�ٻ�́�ێ)ܙͣ��Y�k�����`J�6�M��ykrY#2Wn�s��������]׶�-׬&�N��s�p�H���;Ovy�kl�G���������ο���y���;l�[���<�d���G^l��ܴ���7Q�C�݆�>�������f���b�p�cD;��z�h�V��9�;��ծrlrubwc�sR�;�/���n��py���9M��L��ۨ��
�Rܩ&�ʪ^_�~I_�*HL�����/?7X�Z0ܕ�c�H�S,�3z8���ր��	ˎ
���޵�^������=�^�� �	9i�_L��b�wū]�!�I>C�d]���o?~�-�����5~~#�� ����N�&		Ǉ�_+���ϫ���ˀ��/}�b�p����?;�w��>m�kbB��	}�=��U�&���:i�7/f�%��}7�@������~�,q����5���ǚ[ڑI�F�!��i�k� ��ˡ�D0�x�er�����E��B��t���KV��N���_	O�~�y䏝��������s AYG+�[gI�NPbL%�3��Š��� �M�2v Cj��n��?Ѝ
8(F��-�Wm���v���N�m{�C#�r�-^�pf-2���G���A��l�,�Y�hX�3P��Y�id�ܾc�b���\)T��t�}ϰBє~n��4���R,�V@��̠ ��w���2���Ub�� 7�4����R������+��ڕ"�����b����i��jHDI�;����3*�Q�t"f=$�rZ�:)DӀ����� |a�K����ZR��{��^���\Ȁ7�����b�(��χ��_����oM��tvNV_��]x�D���� ��u��ƍ�d�pQ�g�+&��U-�uGd���"ɔ���Єdw�9s}�``�pĀ:g6�� �k.�yg9I��H$�ED�C�VIw���!�Ӌ���}�i���̮<�ܒa�b�g��rF1/�ųmi��jU>������L��SY�!��к� �	��{�s�F
�=?N��@��N:0�g�"u��u��qe���x��A��\�w9vR�x��>��n��Tr.?j���0��=�r�p�#'�G�$D�i s��B�ςT�{M)ALn���n0 #�	�"D�H���^B��w�>}�u���ŀIC@H�G�� S� r�j�� >|"}�H�R������^C��}J� Z+SN棶�YL[eO=V�6Nv�8�-G�h
,���ʺ�k�}�i�y��R.,��oi�ho��.�<p��η���.�E�5m���S�jL6�O���C�(0���[�M4�'�^ĔA�Gx,��u�o@@���XC�@�$6�
\0G+��� ��f�l��",L��"&��� q�y*JmQ��[MS5���S���>�i85w�x�c��4�Ʈ\ DzS ��l�3�#'��:�r�f���Ϝ|Icф��D6X�w�O��d��O��})L`�9���'k����h��[;�ŒF��T��	���ir��K�����>X�ޮ̑�hB �f{�� ����x%'s=پ}*P/�1�d�Є�$�%� �_C���v��VY\��Js#�Q�7n�Y;c��K㴋�h�蓜1tLka<C�E�Zm���M*$Ne�O��3�T�S`N������8zX���q` �A���pJ�4 *Y]�л�a�5�&��,M���u5�����2g�lG���ł�������Zb��Jm0D�*�����3D�\�L"x'C��f�<�n���U:��jjr0ѭ�R��͵"���G�8g�>~��\p��O��{� � �� {'Ԗ���]ُ��m��6Cκ�`�e�D�l漫#v��x�r��th1��U�N�m�JP�ڢ@��6�A��!m��O�W��T#�gP��`�C��5��s��%n�(���u͸��Y� �-��bX����0�����A�Aѯk� X�_yz֓����@�;5 ���lG����ϸ*�#�##�i�ŗ�^
�ūt?��P��2ֽwR���V�X�I,��y��柕n�X$����c�0�Ϗ�܈��ʭЌ����m�F06�MY�3�	�E�v\��q8��L�kw�ͨ�ޒu+��p�
�ށ�'2�i��;�'f�ϧs���&ڨ{n��דwvl�k^�말�ҖKW�N��%��hd�7E��v�SB!�n�xJR�dVY#���Ǫ�����/��}�Fw�"#iu���,(�v���f����V1j�;����,e,�1��1Q���i�o���ң������_A�*s�F7uz�K��I3ŦR��aٺ�X�t�u��9\�:c��x�ၳ�e�`]0�,����Y��MԠ��&�",���	��N�|j�l:�C����89nj�on!�qqiZ���ҫ�S|hV�h޻�q%$ �dei�����U�0�O5�[��op�*(V��uej�ޡ[�:�+/e��%����쳛��
���x����5���N��܏o6��Y#MD�Vv��:!V�x��i2E�vf�j�uסjeKSWK�������*�)�L�s���_˦w>�;x��K鱵��a�Ȝ�j�5��|LRh���*�V�V�w;q%bd�Gk�У���9n��!���V�i�r@����2e�t��P\-Ԣ��dèI������ lNdI�t��Kʰ�S
�{N�޺���Cٹ���T�CݹEt��>�|�خ���[N���;B2�sf�f�݋��������֘��{�@,Y�Q-2w�A�J`�����1�F�<f �L�?9�
�� ���*j���i�a���z��"	A�VJ^-6�낱�����0�mϦ�ʭ� 6@�^}�,��]U �w-�Ӳ�X A ��wٵx� ���& ��9�@�+i�{V���)4�t��ڪ�"B������,�����8���s{12Ӏ�%��@��_{24 �V|ٺSl������T� ��@$�2F�[�TR�=�R�q�kJp�%�  ���(y;�G���$VD�G���hc�����ޒh�X�0�#�����G�v�m�� -�#ͫl C�9�pM>4���Cj��N��c WŸ���6��1qҼ>7]]��\NN;v��ن]n7 ���uۧ��Jܸ;5��ѝ��k�����{�ffSd�n���5����X����0 ͍� )p�^�n����m\�*Ji���<�@pb R�@��m&ݷO|��K޿�f!/�{�>��_4֌�@�]lD�Ѓq}T-lB{�ʼ&�L�6�ڐ@���@��yG�U!J��Y2���@�2X�8g͟d��bch ]g��+��������k[���t� �Ҫ�M��h߾�Aݯvs#���v�P$"� �[B�?]Hw��x��N�-1 V�N}U��m�,��y{�@����}]�i=�W�;I��� /MMD�e�	���=����2���@�fj�h@��_(��!� A-����q�Sh Z�#@�  �*Z@�H���ｓk :��� ���3�g:�z��gϨR� F��A�~]Չ� ��EpaE��BKp:��}.�P��n��>����
�.S 
M�w�-�B����j_�Jpә�����6Zi�M8M���<�ɹ�>����=�9>�f�8g�4)� �%��D�ۙ�d�����"�H��b�j�p �-�;��Y� t6 � �׽2 �@�n.���?)�;w�哽��P����b�n�c7�����z��'NSޫ�gh�(@x��fL�Q�����u���wFE��Һ����TƂ}��^.��q�u_��m���	�o�ż��S2���R�&�u+���"�d=i*=q�4}�@���D� z#�1c���y�b�wR�*Q�F��q��\��� (���n�d�$�T$�T* ",��{V�	�g�q���2=�p[W+�T�~�2\v���x��2����kQ��A��4�M���sv�1`Lk���sv�4�H��D�E	)!6{J��U��n�M A	1D�}w�]�dXV�>BP=��s)O>�"�ȩ�Ӱ�m��n��,����Ք:Ċ}���bX'��I`
ͧ���ȭ
�IE�ks�_V��t�-��a�'�H�:Ț�� �� E�FǦ��� .���>� ���x֎�ppq�$��(��)��w1Z��A�֝��^m��Bdd�=rK��4M0sSp��BR(LRD�<����@E�xq�=����OU�b}�G�R��O���xq8r8pE��CP��:\,#D��\D��T�I}\�ͥU�*0����
(Q��ng��IjEX'e_i���L�tD�!WS��o&%�����ˮ2%�A��y��B��z�𤷢}Ff�DX�!�ZdZ"�w[�k�}���">!*!�}���Y��P����^�!n! .�$L\�hm�Ri�R�)mU+Q�p�R(R�f �>��U�-B�BbS�����)��v��gQ(��$Q"���ݕqf�T�}֬�_v���!h�]0����>�>�ű
�z�L��i�̺v*B��OgC٢�%�Zm0�3]��;��,Vq�-��1��s�hվP�BɲV��#�7�ʼ�ۿ�'�mgt콲�/W�ێ$���y���S��!�[��������PK��Wna%99�խ�y��9�]�1s��n��D;�w%�W5�I8Ϛ�y��݀��bm��R؍�kqcz���n=�X�m��M�LD���n��k�d��s�ir���;fD�=�[s\sv㮂h}m.��==�Y8�e��ٹ�����.�q����v���Bl�dg·;�c�n�ۘ�Z����:/�x��|g��m�:3�g�A�m��u���fj��	&E��?
!u��$O�+u�Bܮ�E�}�[N �"n�6��
��oO�H����..+>��s2��h��9
��Z��(���ϯ�`�_{�k�k�Dsr@!Q|U�'�Dއe�!BMSV���!M�R@���S�(��64��z�4� ��Q��%_qn�P�i#@�j�p�_Jb������مGy�;�Ė�)�����R�	 Y�L	�,Օwy� I�Eᐓ�:R� ꦚ�%�5U� �Ke�	�a}iT��e�ڸ�MD��� ϱ���C÷f����*�����o�B\��E/��M�X�H�
"��Jw�v�9�Q��>������o�_jN*'Q]tA! ��%���!�J��9����,�Q*<��b�p�	Yb�C�آJ��3{sp���(PĤ����+��f�^��d���r����Scz=W�$L�)G���b��Do���¥T�S3Rɪ�h	�j�J��Ԋ��˂�n�F
��q��I�.��r1��%nlx=�ɴ��RB�jE��aϺ���e>u���#@S٘�1\[��&'��q�}�0�4�5蒴E�"QݫLºv��.og2��˃�1��t�	�C��2�a���'�<k���[Tv�,���{L��GDmͪ��"�[o�@�˙H��빒.��f�,aES�JH�K�w��@J�
@z�2"�*��wmZ����w^�� "� ���}��w)dz��!��!*#�)W;�F!����D�N�p��'B�@$����/uZ�Q�{k��j^�n�#�O-3�DƋ˱7rf*�:M��Er�r�͍�z�A'����TOX���t�Y*��C b����n���Bb���ID3�2w�O��p0��\߁"+Ȳ���j���x���P��[*��i�*�K������Mښ�K��"$��ʾ��h���Q]sMBu3Fs���O_�8�K���j�рX��K�����q-G��\�q��#3���:��Q���P����Z/�Q2�]y�"!3>|)� y���L���UЀE�O�ٴ��a
JJj$���k�j4Cq�6�]��u\a�H%����j�=HBq����-��4��)�S"�I���"��T�Ԣ�j���#�Ȣ/�U"'�ܩ����2Ező�|.���{ �Q�)^�/z�|4��#́UZ��4���=�{�p�H����0 ���S����/�4�	��1G�>��e��u3k�n�}�j��n9���G/n}�㝞[�����=��p[��s������j�7RK��h^�fH���${C̍��d`DG{7������E�\*�
��f]tNnf�q�wZ8��R��L�z��(W�詵.�]��!V��/�$@�G!+�m-��؄�Vϗ}3Q#�G���|Wz|0�>$(ڷ#�뚟��<�"�� "A��H�=gȓ{̋>ӗ c��$ Ζ�-C����_7X)�D�&��FF����+�L�K�-��?��lj�4�w&��#�n��16)�}}���Z�����7%K��3k/0x�79�4��V�-��˧�	�_����F�ZӠ���r��׮ �ʵ�C�먯,�LU�X�|ϸȈ�9�&D��Ƙ%b��I|�t��H"m�jOd�V�=����t
}ku�>�A���\$���:<���]�)�+"��mJ�Q#�:���k���M� �"^^�h���D�gZ}���>	u���٩b�2%��� �]cm�̤�ZR����D��;�%������Gx�(��$���k߹<2��{}7"F'�U�D���_e�f�3G*>�
�K�&#;�V��� ��Ȑ���)Twf�K�J��nDT�S��-���"@�U1�\���҆�c�n�q�Mю.����	��뢻#UK�
E6���c�����2yt�@��D�k���7����P�˄�~�$�u;�3sJ�n�,�+F"�a�<��$�0�G�R���}3�&pd)�x��G�s�3�u3��LQiI<u�2h�!<�Ґ(��̡|�N�:��;jĔ�B��_;;��b�XE�ȅ��@W�����=���q� �NQ�Y�:�w�=؏M�|������B�����$����t:���/��^&�<@d[�"�[|��C�bH��Η�$@�~͜͹�W6D1=p�{����C�d��U)1C&g�9��@����7p,� mG��x:��NWi �,��O�����4��h5<Cc
ѓ�,v�rLy����ds����ơ�~j�]�)�*�� ��"�6|$Ζj^������XN�ΜQ��G_m�*�[wT�{�)��uՓ6��Y�w�n��z�L���dn�^`�OKL݁�"J7vޮCuV��[PG� a{��1��9��2�@�T@����X�p��ڢ~[(�W]��I�6*�O�s����+e��d�]�V�R$�x�g�_{Si`�$MKO���k��j>�|��G�5c�>����
3�39��.���u�ō�=�{r���mQ�n�n��mcaJ�
D"Ў��[iv���#��L�ƾ�݌�MS@'�b(�Z��H�{w���kX����I?8��U�@��bb�mw������<o���|j%�ժk1Lج��+��Љc-V1�I�j��"��X�ޚS'{�׌�b�03=[X��ʍQ/G����j�.y���U�&���R��Vk���&m) =}�>�Ь� ���n���I>iUo�j,�RB�K�]-<��=P�k�X��y�-��Q G;���(�]Ѿ�X[0)��|#ϝdH�� e�4gv��ͮC��1�-�kq8��b���)5�*0�A�z��V�F�g{M�,��Vď\A��S� � �ɞ��T$�4|�Y����s�����p�a.w��-�6츋�륤��7S(d"+Q���n!5�cM;޽�G l+(��Ӵ�WܪV�nڵm7���z�����=�=O0��فF�&v��v���\Ew��ҫ�)4�)�Ȓ>oyO�&߰�B>������.0`s�!X�*�U!�J4gJ�[���L�iM���,
�Fh�Y�f�22o�c0f4�`�H�$�:�5���\�P�o�QޢXI���63(_�����yә]���v��M���ϒ�yr9�8��|WA!��$�s�U��6�sO�C5�Y���q�v8]�Iݞ�/e�:���ͷhqa�<��h粯1�zv�ַ[1��V�ӗ�����]EnŻv8Ƙ����Ӵlɬsq�m�uzksJm�Ecq��O	k���D���Y�<>�v��2��[v�!�Yۥ�����y���q�u��[��fU\X·�nz�"ѶӵO.�n�ɬ��@8�3wB�Q߷�os��'�)���`��$��=��q� Q��b@��,�.�>�T]�a_..)��a�\�QdK��tȌ�m��G#=~SK�[Z��Q��k(ZWt(Q��o���ڍ��"+��ۚ�34w�-�!}U��9i��B��]П�z�E�,	�g̊�
}���� B�kr2N��{z: Gx�4���wY
�+R�b�[iG'1�����v��S1N�9�Q|�t"c-"H�k�tq�5]3r7��đ��S�Q�W0�2`��¨� Q��]y�Ա���|��L>+V��kd Aݹ*�5�;ʽdK�Țr�֝��`���j��}!QR &Ơ��'rd2p�>ۜ�P��2�ٸ�������y�#� l⩒��˪�Y���p[����֗����ϕ���[��&��5�S�#;7���X�R�4RGe�>��.�lr���iHw�+��vl�t�1��6g���
���3W<[t��<ݼ���\�x3ۮ,U8�tNYSb�IK�خ�B�U�5�Cib�Ԋ�E���k�^y�j ��y3G̲I����>�S��ܡ�B�s����4�N])��>&�y0Qל�&0(d�À�L��CO��G�@ɼ�y&�[�"Ji�1㗣�-�J�����;�,o0��h���;�-�z^�k���L���[�@J��2DtYqgRq�є�����ɒ��z��GȗM��hz�J�A�AP� w�������0�rQ�ʚĸ�b���8*ݤ����i�0���b�/�����cz�P�I�<���yB���sxdU��\\��m���W�=�~��X�� ��,�V�6n�:H�d��Վ�I��Ζn�"��`�a"H`�9��l�3���4�;��	-}37�yt�1s��҇li���k=���!���N&��Q��}.�y
��oE������m�ٺ]Z�#pF������<y���;�"�(b@����}O�VM�J@�LG�����_r5Cd9�ي�k�Ǘ�<��m�\�k��@$�n����Ռ\�g)��p��m[�P�
P���A���މl��|m�	'z���̆E�9b�X��g9�cDaǁ��sTh��^�2#ټf���&b&�j����V���qʠG(��	u��L���;\ējzkk�z��'����uկEz�Υ']b����w�L�TzG_^���OO�HʕQ�Ʋ�ݣ� � ��˄�zɣ7*�"N�o*���
a%�]G����I8b1nޅ$ݝ'
���P��Ol��à�� 9��jĥs]�-d++D�$,6+�or!V�2�s���-����j�H�x�����G>߅4�hC@�\��&��T���-$��ė��ko����ڊبv1f��QGy�ĉǏ�Q���\�����]�N�ۖ��_��|f�ՠ�q��~Uj4�V������ޏX7.lr�U�����׽Ԣ�fAY�S�I��E�##
u[Α���Jxh����{*����*'*���"u(�띣�ޓ�a�96ܗ:�"wY�kr^�kY�_����
&�'n�m^֢ݷ0%O�m�mZC�����pݒ��Ocj�2D��T�e��h��G1�~����B>>;;�w�c���a4س[��ͻ�^����y�_[0�b��29����]|d<�Ϡn�ȣ�J���Pb5J`�"׌Ґ��%)
֟O`��cF�r՘2�3{_u�2���>9s�o��k�I�Lp��D��!N������f��֔�TH(�rY
����0�Nw�oD�C~3��VK���`|��P�z��#�ύO;��"�7`�!ĮU!�C�}{&���8h�ln���e�s�d����E�-s�H�ћN��Ŏ���z1;'F+�Xɱ4`�;)�s�08]c�����ii����l���y�.��
�f��N�EW-��5����]����}�j��S�A�G�9�m(x�ڱȠ�+N R6	���N4���,v�����E�=]�Ym2�3<�t8��	�:��/\}���g�[�X�^�9T����]�_���=՜!��1_=:��cy� ���G.0#�z(gb|r,kh������Z�������gJV��r�
v��(�t��خ��K*�B��<�g�5�K�wkZ=��qm	I*+LNX)�q�gIw��f�����u�n��u����\Kv�^�
:�ϸeм������n��P�e��A�x�V�]�ƺ�q];�2�`��1+<�e�4�vv:9vY�H��h�Tڠ����PPn�Ѣ�Q�Y7�3�3"��[K9І�I� �F���"YT�l��[k3}_`��(C���?P�}B�>B�?����T�,��_�P��!�|�}��4!�!�!�!�!�!�!�!�(C�1AY&SY�?2��vـhP��3'� b:���t�

�M�Ђ{j.��3r�-�M�*��0r� 	R�W;��JQ
�SMX%]vȔ�5��B��Jv݊�ʃ���                     �  @           @        �U=4��ɧj�mE��:t��QOt:����s���I
\� ��P�t���z�{�:^�7��ۄ���I҆��	y5vi�d�x h($Qfh�M�M^0�^ϻ�h��'�  =  ��       �X {Ǿ��[nM< ��Gmݮ��S�:kN�sOm㻻c�Ӷ�v�]���N7�w���;z�5.�<Ov��ݛ��ޯ,����|���ۧnmCN�h�N�����        w��k;w�n�����{��ڶ���x��m�����g\O ��;�*x�گw]�Yy;�y7xޕ���s�|��_qv6k�� <��h��o7���q�\�<�=���n�
�]��<���]�wt�o&���V��� _y����������by�ֽkQ4i�݊h���-]���g�b�� {�ϰ2}��n�s�vww�;vocs�]E���jq��}�{��mKmwP�M:���9� �      ��sv�l�����uWko��YV�vx���X�ƹt�SY�ˀn�
��x�<V�oko��6ٮ�u�f�n��yit��Z�������2��^��k�����mV٢�\��(��v�����.������Qݼ =޻���ǜ���,���]��ջ;��⽛���o=�[�px 7���x�v5�춷�=�}w�;o8w���5�����[y����4�x  �    P �{m�M����m��=��'�����ޝ�n�7������ܞ by�m���ַ9ݾ��ﻷS��o �=&����� s�>�����=w%˧��{54u�UѠ���kږ��7P�w%�� ۷�4����ڻ[�w�w�c��v��R��%����< ��#E��s��,�v�7�1�����9���m��]�(�:�S�         ;ǭ��;˗y�嶶�9;���j]�է�<��ݹ�Y� ��U������wi]y���ڜ��t�G��מ�d��i�| ��}E��}�A}�m��=ݼ�˲�:6�ݱy��}�m�j�l/m%m��-�� <k�=���[k��#v���v�܍F�f�楺㧍�j����ux�7�qSo]��o ����]�ӧ^N�o���mkSl��Py�)A�Z������;>wv���T�� �~�R� 0�$�T ` )�bOEUA�4 ��j�@�*   ���*�� �MB���� ��O��?�~K����*�%�����=_g��,Q�+�G��5u���f9�g�I$I4�ВH�Y	!$���IO�I$I?�$�!$BI	$$?��������5"���j����Y��V�cUc��ICB����6&��h�ᗡZ���'Y�6 u�m݆��gnt��E��vӛ�T�&2�9b+h�Ռ[��oؐf,۹�)9��N�*�6۩(�Ř)��"Ŝ�j�L-e��ܥ�v���HMHot�;W�]ܒ"섅���nk��4sDh����+o2�Z/9^az*�I�a���ޱp̫�r���і[��5j��Kdm�Sm�H���b�[H��7w��\�o	�m�-,9d��֑8�;C63�O0�Bܤ�Y{�,*Ǵ�"�G�d�8-�W2�6�G�a���d�n,U����E�-� ��>7p
q�a��p7ZPu]-�F�Xj,g�N����p]f3�+A�mۼR�NX���8@�;b̸��v����Vok)-�cll�h�\V���jCg&`_k�#v�k2�\�A2o�*R�`�槈�]5ÕlF�rm6����F�8�ɔ�[�l�Ѻ��$����sp[V��X��Vh�4`��2�(nm,�L(����R�v>I�)$�ݳE$X������`��,�O$٪i-,X ����k%+UGu���Z	�P���W�d��whV�kL�<f����
d�Jt\7�h�%��X/(%� �i�nP2�[�BZ�c�0I�/;�eJ����ϙ3�Q��ܽ��킷u3 3QP
��ܕnaf�̣��"0�f���3k�gM]ģ�Z���i�ۿ��f)`�-�Y_'p��M}�ڇ5)��:-���5�[F�X�:��-+7���M;������ڎwU���d�3Ҭ�ۼ۰���m6��\&ׄ�X�8�����{%�J�=�W�>,�v]�Qcb�����尯��r�&�z��͝������Hb	/���b6��N���KU�<�X�э�L]�co-Pb�%iRJѷ��	�am���	5���F�:)SD��LÔC�b����I_۬�5��L�Gb��wf֦.n����$M�[@�E���a�»O���F�CX��^�aڀ�^%UO:%��j+V����(��HG10��z�]�ٱ}�e�T���\˶�Jj�����o.+Â/��؅t/Q��]�^
�e ��p�Dń7f,�U4�1)�R�ض�W�����M1�X�ֲ�6��&�����fY�^��wOC��"������m�b�I�`�j|酛6c�Oy�wV�v�R����6���KV���d:���!5�Uϒ-���2�5����@Ԭ,��Gr��Q�e���p��@;�b�Շ�ڂr�@�^�kB褮�#e$U���v]�^F]����Я����ƆXӸ)
3iLt�Wo�6IB�7���	����%�VԀ�2�h��ՠ�t'�emӍq��[V0;U�p^��-�ʆ�KK�b�Kf��+�L�Oez�5qa"�Y�ͨhN�Vr�L�V���Q��-�r�Mm*
�Ux̆
#����{�V:ͻ�Tf����U�����.�yM-��K�����&��SixԞ�=- fyf�A. �9Hc� #�O�u�A�%�ɳ�ڸ�.ȵ�`ݘ'�F,��h��m�eS���*����n�[R��	3Y�6j��W��g��]���U;�"T+Q�A-g6�H���*�;Im��f�VDs#�[��*m	�I�I���®��:��dK��'@�d˽F�w�Z�9p�ii������ۤ�aQ��Q*�H] �a�[��,��e����M+Ĵ^�aJ�[h�Rt(���sxu�s2�󉪙ˬ̫�n�ر�-���µ)dfQG<�P\4��Ukcoj��m�+$x�u���@;�Qi;oSDv�����-�n��B�k#�i�ܐ�P�dSf����r)�X��k%2R�đ���ln]խ��nH�.e��5�jab�!a�S	ͳ�k�7Im= ��۴��f:�4:h���kʺ-�f_t.��*��-�)�X%���z?4i(`��Hf����F�����*���ॻl�Ux����^�8M��h�Z�+��X;z��(�F)%�u�L��L�w*���s4 p<�'�*B�c2��5�3���5�޾x�P�������~����(�` E�!9,��u�;��x��Aa�L���F�F����YP�w&�;6
����IFN��ة��AR���:���H��5&����1|E�-IF�0d� q�v+�[R�i�e�@eb��s�8uD�;��-�b[4+b6!a�-�&����SF��0�W��S���t�w��ۻ�-���kf�"�Ŗ����:�,�u�)ޤ�/]���HvX�/�V�G2����.��� ����8�j��D�k�a+E�Jj57$��ѷtW�v�2W�8�I▆f�;�Hi�	�ȱ7\�[P��ڰ�ʳ驺Y70�aj�����d"�y@˨*i��,�Y�ԩcY�N"͡Y.Gz����[��qb�a�K'Ƌ�OqS4q�U�(���u(TZ%m�����غ��D7GĈ�{'UX`�L[{dY�L���Ũ�2(0*����ʟY�9gEa�	۷n�A]=2ժ�7v��ܔnj�(ۂ�WJ��YS(�:7X۔�r�̠tL�����L�:��ȫKU�HΩ���.]��v08��NUд�3l��X��ô��*Ri�)���<�A��8�V����]�ڴ�d�"b�*B�Ų4W4!�Yt�Rkr�/0h9n���H�ո�$���D��&-U������mb�]a�i����f�VG��+?cHL&vû��̚��A�^%��.��Ki�te�sq�ʽ����)L�4"f��Va-Ճ���v�1[j�0QY+oZ4�BhKٸ�6q���]��+.�vK
���Uh�0嵎H΋�YEobh氕5�@1�0Z2����ˬ�K{�M�7������!dTq�W����\t2`��z%S�c�U��gs-n] ��75;͔@`�T�!�7R�w���5�F+j�l�	�q��aV+W����2�Ѻ�e'K
�ۂe�0�����^�v�x#zJ2�-��hAtf�ٲ&Vh��W�eH�`B ��	���7kĻt�����ن���ݘM�A[��2�I��H::V��*=�$�eFn�c	�ys��VA��r��֔u�Fֶ���/%�ڣ�pk�$Bi���a��;׶�}�`Y���h���ӂ]Kʍ&n��ޢUl�"��ٛv҂�0`�w
��iMX�$\�c7h}ǮG����)e�֮x����5�3�q�����K��Pf��.��j�Y𚧎]���ؔ5�b��~8�`��{�e�C�	�s(c^�ywP�k��1��ae�y(�E�zuZB��D�V��L�Q�Rd�Q���4�!�����3!7�\�>[˱��r��fm'E�����9<�
�fլ^� 2��wtFV��ǂ4�X�����A-+ɦ�+Tf/�L~x��F�D+L&� �����4}���9k/v��&6�'�_n�?���b�tOX��5�r���k���>^sn�2Xo6�9�2i{�*��F��W���6S1��I�!	�@S�����S-L`�\��*�kbaz"m�ɉ[���ZZYWG5K�*��s{�$AE�����щ�r�D5[j{uU�}{���6��aV�	��ϱcC1�EQ���]oF4"]#tf�d�'�n��j@�t���C]�U��.�ے��/n�J���cn(啟,%�t���z-l��uyV2�R�w�SsL'P,L.^�Z�xQ�l�����ݦf)Z���)ܻ���wY�"FǬ㺊�ܘ��4H�U/E�IG\Ut����wSQF�@�|�T���1�j�`��:n�l�v�!I)f��BX��E7��,%��
�i81@�=�L�pcHc
͊�P�;�%W,$RY�vܺkVY�-��(�#�Z䃧׌����b�d*�4]&s-1yy���y�RP�ⵑ��$t���/r�e;/���60W�	v5߫a��^��2����E��z�
�V��44Xx�i���Շ�0��ע��T@^#��i�J��{hH����u�j�C&ސCүm�I�ͭךQ�R�ܖ��9F�NZN^Ȯ�+?RL(�A�N�=T1*I�!��n�l��[{�w7c�[��B�lC�Y*ʵ<�G�>�D�mZ�<M� ��
VR�HX���'�h��)�7.&f�����5Yt ��LdUp�̹�n�ЩKm�Z�giջV��G�U�ts� ������,ޖ6 �U��^Q�������vj;�|�:�voUBd��
'w4��`��fݬ����*P�v���u��ⵢ�NG�
��!�iV\���&T��J��')�k1~f ��o]�M«0�`�֚̌�q���q�׳>���j������+Y��]��3X1 ^�I
���!U��:�Y��9���kqSۙ�%��[i9���!Z�^l��cB6Ҕws%G��K�Nm�ݦVȪ�+u��D�NcWlVأDg�wvn+yX��.�Ѳ�X����aS.ɔ�P�r�j�ֽvBQ�{�-V�a]�2�=v
ǹ�F�h�Ĳ+S�R�JU��]����['jj2H�r��U���ܭ�k`Z���r����MB����tT�����"m��Y6a��[��F۽��+�EV�Rdʖ3v�h���n��P���5�RUp4�6�n928v�Gqc�-נ���[�)��Bc��ԣ���x��bl��0vV�\]F���e^X���f�e�U��ɷsY�u5��3�^һĸ�U�聵�;Z��s2aO[I�#u�yy��%�ތ��!V��\���h���q��)TE�o��B��V)Q@��Zp�|Λ�h����J8��{�a�k2!w�������mŵL� �$7����N�%v*
�:jڅ^Tq�e]�N%�6�����]"2�GlUX���n<̈���VE卡���(Q?5�8!V���t0c�pU�12ā-�a;�{Ui	֛2��%<�bg��(Zϕ�R��b����cL��Y��'km��u��^R� �D����Yz十k�ܭ�ۧ�,�ɘ.ì��MBc��&ܑ���YQ���BNV,�۽�N�)�mjq�U7���X�![l�u	�����w�&�IKɵ��@[Wif�	��^cw����F���� ��E�GoU-��V���4��
�3G{ �7F�]$CY�$l����zE�>Al�-�`>WmBfa.�B'��I2���E�u2فO�����n��I^b_&����2;d+;��qj�B��JD�R��M��kO�`�7k,��y�Qs$n�ʡD�Q�R�WtVB��y�r7[l�1��Yu�22V\�j`
�4��T	� �5��ʬ�9S��wv�E��3$pU�� g*Ej��[�)�ӎCyc�p�͂���Z^���&�n�+N9@3LXb��x�z%��e���f��mͳ�rPƖ4��"c.���q��/�c]���l���&ōו�aSњ5�*\AVf$%��2�$By��h�e!xv5kl�B��&��g6R�QC��wCt�k�s`�����&�b,�v�P��ަs�M�z��	ٸЭt�DS'K����R��:WP#�����˺
�L�$t-;[��
�-�Ӓ��]�5���1�^ca���n��I��;L��\Ȍ�j�����"i%�&�u��kp��閭��KD����֬H�v�;r"��4���y���
� YԽ�5f�Ν�TܹJ�z͛^�h�
��I�4T2��ق9,�A���E���ֲ8�x�� �df��l<�l5\L����SP�ҳ4l2�]=�K�
N�[�����M��OL�h,ŉ]���j�G�,�x�[`&Dl`�y��E���$V����"u�&e���6���:#�ص�\V�Q��u%�]7j���qL͏!�u�������ahџ\��S	��q'	Ɍ���zJU���d����k�S�]�{7V�aa�b�Q2��]#'k��o���A]⸬M��7 ��WukDٳp�BCy�z򠣬b^]��5�Z���:I��up��yb�$��1F��b���cKB�I������7�-�*�ɘ�c��Bo��n��v޳���u�Gv�a�A,9��hAP��C>��BlCC�t�R�A115)U�E�]f��V�s�*��86[��B�i�A[����]B�ɀ�OIJ#��2aV0p�U�����[4JN�,���T���f\ȴ���(T�yi�\Y�.ZjW���O��czңf�!1&iK�Je7-���nE�7;O1K��ӻR��A	/ƚmjW/p��/Ȍ� ��0�d���
�G�6�-��1Xp�#��&Z��N��L�SB"�/������,�p�+)Z�J.�Bc*�ԭ���;���{3d��MAW�f�i�\��݄Qb��e��&n�0S�0��t����WRa�f;q��ݨo$Q�f�	!FӫW�sB^#�ҵ�^,��*���yP�R�+wF�/�:�l�J�
���0�1m�i-b�GaM˳�w}i*X� #��4�L�}��0`f����L�&Md�x��r�izua���"@�o���I{�*�Y��YTի�fL8�iVh��`xʺ9���jɷ7UbµZ���+�Z�V�U~aL(��vƽ��5�@��l�>2�T����	�m�Ŏ�+<b#��P0�t�,t����r[��E
�$l�dj,v�v�m-�W+.]8����]��&y�Xv�%�y��v�6��m�m�bӠ����P3���ӎ'����竷;����r��f�A�m�r[n5�	��'�w\Σ�8۪�9>�K�!�lx����٧�7�y��E�������!�n�[��뮍�rs��y�G���[�=�/c���B��gqq�;�1�MB�<v�P��f�s�M������1�/��2U[��-ώ�7#����L��j�W;k�N݇�V4��n�v�έv���b���K���m<�W\v��c���������0�h�=�{T����=�NmV�]<�d냰#�].ۥ�En�\����7.�z��اkq��+xR��/ h΋r.�H3xz�7�Hv�'6��؈��6_-�r]�����ϝ���wn�-�u���r�Ψ9�^�Ȧ�ѹk)�'�������|��K����n�mX�#�OMΏf!ވ6���n�<V쵸޶�8���9ӹ��os��f뭹4y�>v�{ӝ�����K���������+�ܔg��ll���0!��������%]��3��|^M�5(p��!ݸ���Ε�ܹ�\k�X뛷N��f���^��3�^�ݤ2�v˯E�j㳺h��p���g\�]�^���w۠�h�狄��o><`21p5���N�Vݛ�@��kd�>{��*v�X�M�]�OnN�ei�-��� ���7kt=����]v"��<���y�u��mr)�-�����Z�;�\n��m���i�<�v̽kr����qc;���9;.���d��"-i���Ȇu��`�ƫ5lH箍�w8�Aݵ��*}�;�vqy���������tGRp%����I����6�{5uqWWN8Ry֬i�Ѳ=��m��n"[�Ca�i�v�+C�m�j�s�ܹW[mٶ�1V2k��.i��Ɇ���ɶ�r�$ۛ�^���<XL���sq*W3���k�<v��;��GH��۴�>��t������j��㙹��x�m��6Ȃ+mq^�\pi��ݳ'n1���k���Lf�<�e�1��nGi7q�y�	�<�:�Y�v;;h�u���l�N��ϋqho|���z��Z�n8�7gtB���p��n�ktg��kQ��t&:���[m��{q�S�p'V���=on�^�!�0��g`8��
m��ٻ]�6����x1B����na�{q�c�ݔ���Q�v�y���ݺa�L�hy6.Y��H�є�1<t��1��h�$K����w<De���vEzt<����fMv��6��I�u�Gd��,a�I��r�ss���:q�/8�׮4�]ۛ:t�v�k�-�Q�����Nnu���cƧN:�kWJq���m���y��b�tta��ch.^݀��-��kk��:tD(`�\���<��^�G\l��\�m; kk]�'[�%��0h��� ^_F%�7/�C�1��8�������pm�����c�����S,$��Y8����g�v�O?,�m�|�5���܅W6�T.{un ����qr3G��g���uOB�b�v;f5T���y��,;���=��8MT����;kF���r�aJ��9|��앍����O8{G,&������ެ^7e�%G=/<hl�)V��u��*.^ݐ:9�^+�����Q��mک<7nx뱊��e��<�{\��s{ttt[��%qo�u1v�k��Qڷ��'f:�N����ñv�P��)#���]r�l4��3i�E�q��\\@��Xݳ���n���vن�;��7A�«�uT�"q�"wn�n�rd6]�u���*!87\ۓ-�r�]�;#OJn��m��T�m�&vN�6�vM�;s���[�q��W\�ʱ���ݓ���S�>;f�j��1ӺP�Π��6��H��-�m�1c�/i�[��[�6���k���je��3v�펲�Y�������9�9��K�l�E��Y6�sz%Nۋ�\�,�>���nM�c��o\}Ϸq��y�˞ӻm�nw;������^��O�|}����͏\���_q�}�����c0d�N�묢Z����B�i��4��{6��/���A-{<mю}n9��VM�����rS�=c�9���S�����fzA2o��Y�BwlXz�^�Ƽ����ܯs{�u�=b��F1�rm�]���=�����s�{���.�����OA�*���8y�$�Ss�fN{R�k�H�$:�.�}��z��N�NX�:��_Az�g;��C����0���#�9m8��m����)�"�H��,n9cvy�۱��p�Y4��p(uN�3���Ϧ�Fc�/�{Y��<F�p^�ӹ��r;�ݓC��:׭*��+�v.��m;n�q;�9��nv�;qƒV]sx��:� ��ճ�=rn��h7^S#�z�x�Й�x�ӌs�9E�x�H�N}ų���Y!�40��,Y6��.��<��g���qA>��gn�\�#i۩�H觜 ��{k��xշ�
�6�ۙ���M���cM����ڰ�d�������{���1m�WWZ6����9�R�Ė�;#IrJ�]���<s�݂z��]���i�ѯ�D1o7�������ѧg���Y�kWmpv�ۗ����6�='6ty�:��sv,n|�vw;A��<����n�g��rc$����q]����z�c�+��Y|���"m��5�q�3l�K�qv
7�ݸ|����B/7luH���'a��^���okO���ϧn�&ȩI�{pH��ƺ�I� �M�-���K��n�Z2 \Nz�<֧�.ѫ�s�ط^n��sʙ���޶ J���{jq�^z�칛�u[ڋ��N&��c��N�V�������t<���%��3:�S�q�Z'Ec=k��uR^B�����U�c�M�`���·*��xqo(��f0�0�O!�א�a�I�����\�3�Gb���pn/t^��������$-ɧ�*���ήs�	���VÛ-�t�Lm�K�=�Q+���8�6@�wkAj7��x��v��%ʙ�.N��]�M���۶�i1��w�vo;ל�5vGT�6�n/Y�%�v�q���p��Ķ4�x\pݛ۬Y��W�T����v��c��q�;$lۍ��;�m�!U��'�n�p�h��Nz2�p`��.�H�½���^v;�:���qY����o�������]�v���;�Ő�nz;z���:�<� ��xǀ0k���ta��C�=GU�bY�g�.��7��-X�M҃Ҙx��Z���
���$d.�+�;�q�]���ׁb){u����� ��0���0>��ZZ��(\��Zj���lm��t�a���
�moe�g�Fxuפ�k�vӮ�^z�"dיv��҆�su�a��v�o-;�q[�6�2����ޞ7>�����l��-\����n*�+�u���۵�YGb������/s���ݖd�<}�~�v�mۨ��6��8��l��\c��G]���v��o<u�fzt�;s<�X�A.s�7E�����p�Xۺ7:��N�qq��rg�[��d�:�A�綦���v��v�ށ^[P�s�9nj�M��ݎ�k���^�)BkO��b�;WV��9Ŷ�D���dA��6�B\�<A��6n����7:{���g��2�!�k������ϰ�G=&a��*%�m�v�J��GլMn��[��]��C���6��]!��u`�Mɗg���gc�{��G�׻.�v��\�tK�q�1�j���� �vݹ���v���g�B\닗���:�[Qg�9xs�^vG<sCZzU��n/��jY��n�`�u�^������<��s���X1z4��/]frxg=g��m<��}[����U/l��J��t{�u{P{q��x�ӯa�g`�>Cyl7m�6y�\V�V���ڧ��P?�(8�Jm�f�{t(J�v�G�x��E6��3��+��n�9�J�O<n���a��DoOg��v::X����Cw9�gr�X�ٹ��=�t�{����h�
vm��Hc�p�훬�+���q�I�0�s�:bpr�����#��p�s��0��ż���5Z1�;���L��]���S�;W�i�#{vcs����n���ҝ�v�b�\8�U�k&ހ1VwEF�i���;km�.�c�N!�E�m��:8.Zt��8�On�!�v����E�Q��1�n{]>�o4v!^�m�kk]�8�݂v۬T���ݺ�&��k����8{��	�ힱV����������g�Y�Y�=8B�>4Sn<&�u���Z^-�g��=���e�-u�&�Yl;�>�5�b7�Jq�������:���=2cm�gv�یuh�h�soK�zƺt�c�>л�.G�l:�(��k����a���Zy����	�jA6�n���ݲ��E��P�88�Z�Gf9e��������h��K�TYպN$w<�@i3Z���9.oG=���q�n��wg���6��u�.���Ѩܙu���hx���t��~��zNO���x:��m<p��z9�)�|_o�矮8Lt�:�k�e7=�����cF3�r�u��{^xΊ�������V�𘷰+�A�ny��=Wj���\���<�=4]���*X���u�w�t[|�<}w'���t\{V��vk���o>V9�O�l��	�3��'[?W��8v���;�ݵ7�1�z� �ν�cg�Fˍ�끴���8�Jr�;r�so/�8�Y���1<V퓘Mx�7�Ͷ��m�bś
�1�ܠYQ�x�*}{r�݋���6ݜu�����b�垽�.�d;Y�4v{�[�ka�ۛ;v��%���A�uQ�+�c�G�_��� �	N�燶:����v��ѭ���5r�9�+l��-���n�џy�"=9�f�m�[׭�Ź4�q�a�N�]a8�v���u�����;)��=N]q�vL;�նQ�����9�a�}��\�n��\�:�یN�S�Pm.W�iV73���[�R @����6	I�I BH����z�~�rqld.f�E��s�#FvN���v��ݓێSv-[7]�nõ�h�)!�rv5�/���ݐ�a��f�mr�=��mF�K@,��x�iٝ٫�0m���8���lLd�qC��9�޴�ή9 ��p�E(\n'I�x�# �{�+��T�����U�iֻQ��l���X�jܷ\W
o^��=lA�kd�G\�8�y/ pK��V��`L�gu�0�og�@맱��b��<��.ں.�=���d[[֞�&����q����lV���8��\vw<�Î�sny;q�s�ٍ�] 9y�[y���bL�]7Z-ϔ��g��U���z���8�f�;3OnT���F�e�In���bν��C+ݴ\���<n��d������=��N��i�����LI�Kn9.��y��G��ۈs�yu�@[��m&=>��cn��{��nS6�v���8��{��s�����7&xy�lNyגs=��F��j��bN`�[���ze{��p���rcr���{sqW\�d�ϴ=��m�l���� EA������T=��ݞ-I�x��USn��g�:Bu����ۤ��t�/�Wm�糔8�W�gZ�W;�Ns�`C�����qw[��9�<)����"5�v�&�sb��>�E�l=<�ƹ&4;���^G����\���K=���<�A���]v�z8��ڷ=������=�m��x���2A�=�l�ח��T��F���6v�N�WlƼiCFL�8^b����C�s���bҗ%�51=����ۅ�:f,�]=>��؇��:���W����y]I����&��v.g��ݞ[[who	::{[��m�-[���'%=v��8}Z3��E-����.w&I�w���=ru�n=����b���enV�[����W=�� �l[���8g^9n��Q�Qv���v�a�ٮt�p�����Y�V���������>3\θx�pm��(�YHUe��@� �! �"�
��d ,��XH!� ۽;�*��([̕B7ye��s�`}��#��l�m��Ggg��\�q�5�8��;5��c	�� ����{���bwK퇇k��;d�8|\�s�mg&�7�q���vz����ہmŝ=�����,����7\۷�����s睳����;=����qr<]��.��bW�َ�b1������b�;k�[^z��N�ţ�U��ƝU�wq�W=�����=�;&ܧ����7��y�y�')��8|;jm���}��$��j��u��@Z������^T���I��`z��Zޞ�W3�3�o(1:��KJ߳z�ܫC��b���"Z� Q�4?���t�*�v��d�l֨<ß_9�a����<W^�Ob�O0�4?kH��'zA-�C�&ޡ�z�����A�ĖϪ��Hhb�dY�(��m��ۭ�aI�V{Z�65��Ʃ�2���+4�=F��yCJ޾��TͧW���>C��_��I���>�E!G�בkz��ė����*KJ�,-��.�=���I;˸bJa�ޯz�*]W�j���}G� i����˩�����E���ހ��]Y)���}W���̆��fT�������>��<-�W�u�V�χr���!@��>�2p�!�/��3��3���/���Ļ�щ-11��q]z�YA�:d�)�`��+��&i�:e��7T�h�
�%�R����͕z����[!�f���A}�4ҺV~���U�-
3/,��Y��5On�r��-Y0�U�̦��ng�ל�g����ǵ���=���llL�j�:�P�q�z�@�~�q���=�_�E����3IUF8�=p����ԃU1�uT4��YO�!�_}-f����<�Xbi����\����V7�J�i²���S%2{E�n>��Tj� *�V�(�b7C�ښ��*���[qdo�q4f�H�P��g����R�P/�,=�-٬����r�XEn	������IlY3- ��S39�p�+�Kf S>���/6Ͳ�M��wQM'}������I��_k�n����o*ypٓ�[5a�G�$��#��e��$,���9T{��MI�ݩ��UvKE�{u��l6�{�2�Y��{~u����7@�o�5<�N���L5����Tˣȿz���}p���{�9u���X��Va��a
���D}��+K�Ge{\i�
�u�#QOc�#du��[� ����o1�Ri���Xl�{t����e���X~S��_Zl~U�F�%��D��L3��⿚/ƪ���o+*�|�Y�����j����g��+P,�笘��^&wفS�ܢtN0��o���q�*�B���x�-/��L�fJ���}��V	 ����kdǯ}q���q��8xU�b�]�`�շt=��˺۩�[���Q:�v�ӣa���vޠ�����Zu��T<����G:e>Lyy���m1)�� C� �O��;1��m<S�xY��@i<���*�w�룺�4��{�Jd�O]F�)i�����c4Œ�@�;]�R� >b�n|�J'�����*�_[�uvu�j�A����f%������@����d9U�o}�����u��P���V�2}���h�MS�_tџw�]8ݘe��c��?&2w�|���|��&��T�LӶ�:Cj�{~�Ρ���0i�k���ez����Ip3u'���ԳV^�wŇh���=G�}q�6��u��<hkⷷl]7[���9LW�V��wUÅ����V��=�sf����.��?|��F�ˇ�
m�a�
n!�����`��b�-����{l�e���,��%$�{Y8��l�S���/��I#�m����/�4su�gNV�l�y��̶u�K�B�Kn�Y�篍V��n(����d��>��L�7��2��}$�S'����Qګ���_?^a�?B>"���̀!��^�6�C��gSm3~�qZ�s��8�'�ZKKgh�k�͗��lۆ�p���C��;n}m�qk��K�o;�n�ά�6�jZn|��F�dz�VzI����T
}�7���w�6�[����rȦ����&'�Al;TZB۫��X�VY{zVV��/\�YT��SI��O���e���_^]ߙ)8��H�G)ޞ5|��yYwy����u�q����b���;#�Hz_��}a�����_���ٶKe�C1˨z��O2�]f�A�=��2E��V���6�n�k�k5��w�W&�e3������z��8�Ww�=c����ɷ�Cnl��� M��4�8�!y|�.��_����s��ì�+�ӽ�Ѵ�%���'_;Kq��sn���W�ڨi��[��-cU��n^
�P�e�)�k��#�?t�������Q:�6�ʇ�}��7D�}tE-;�������@dq�6�2�6n����yݗiI�SږQ�hޏ+&�P�YO�ʖ�^:��e-���:����J��mg#�]+4��w�^߇�}<���D5��M��[��ٺ��X��JV^Q4�>��������ju�2�!�Q곇��:k��o/;��i���&�S��f�M_nJm�`���v�!�Ѥ(����_AD}��j�{E���Ё�� ��Z!Eģ�h�:�\m�nf�1��WXv��qڮ���0�
���ƲSw��(�����<���.��__��S�-�+���+��n� �}�bƊ�Bv�!u�;2I�2m
eP�;|�����5˳\�l�QM�V%����l�r�:>����Uh���1�$ɔ��m��_��{.ɉOɷ��|��>B�hl�j�X�/��������΋�g����#ܼ@���[�������H\��eaM[N�����24v�q&]��^���d4�5� �1X[+�����#"C�E��vv�V�M�H�0���ݥ!��I�����X�w]��e=x��/��[��RbZ�r�U�5���C�":@�~��P����s�6 �#�α�~­Q��5�>@$�6�Ǐ5Al�m[W�ރ���1,M8�W��Q{���Wl5u���,�Ĥ����O�>��)��t=1�U�1l̼w�i��b{T)�;��V<F0�H��U/���`�T��L�[w�<����jZY����B�[l��^z���1��h�K�5�\v�ɉ�J_��N�--�/6�ck�W���$��묁�;�v^�WG&�
0�/����8��]��C��>
iw�3�z=�/�=��owa�~4�a6I� ʺ-�������eD�[���0�������ɻ�5�uS��:{pqky���T�^��NSmM=AZ�v���v��D�xo=��:�y���	j�-��l�q��3{��k�rx��08k�t u����rj�rBu�Jp��v�P���{\k~|�q��Ʊ��m�}��]�-'�����=����>�z��n�g;qv�8�ό��E��/8�^\��uEr$��Y�p�Ԅ��a��T%�T�)�~��/�	��s�����t�!ј�է�}���~׹�|��R�@�j��[L�w���+�����!K�Pp���:^��k^��J톾�g�s�Xi5�+w�,��o�j�c��
LN0):�Z_��4��^���T��T�?}�/���]��)�h��'�8���yAi&���Ԇt�-V=��;�U���N��i��Tc��`�Ж6aW��l������j���6�-�W_`�����5�U$���a�{�N���g.������V���ʛN:��P��w;`d�*�����௰��}#����H�Y�ǠDx����V>I��i:�S���I���c7�o���6���̖���ӛ���S���d~�**3��+�õ� t��mV��[�Y�$�4c캼\\�eV8�&�3I�|���|��Lϳ����S2R{��u��{w�NQ�5��Pi8��[��V�oF�|�y(�)��e�����:g|�i�Hm��^�w�su��~ó��t�l��E0h��Nf�����1�j�ۓ�]��,q�Cun'���6�K²��
r�3~�@��:&����{�&�:ȧ{�Ѯ���c��T: �>���3����uu��2U��c�<�k���i=����/�gKdT��&Cp}<�W�G�C=h#�f௑����ΘU`GI����٪�c�~���A,<�v�%�B:;�+1;�o	�H�<��7Zu���5KDQ�n궠b���˪���f�]u6��4���}��N�o��m�M8�<�xM�g��5��/6ޞ&&36��u��N�±*��k1��<�U��5�6���p~�bM������S7���6|!��OF��c��Z,4��wL|�W�!�t�.�wu���8�&&�i��}���&��>a��V�ש[<]�Z��n�q�tW�|�"���{�_u��xW�T�ύmSOX�A��,�y�̨;��Mn�u)���Wz��v�(S1��)���S=A=sC �����1�s��b��hc�}%(S��m&bI$V ��'8ѿ����뼯���*i"��w@H���cY��Up?�E}`��s9�h9�Y�Z5]aĽPc�W�p�W}���I���RVz�&2�o�����{U5�`��I6�$��p�����X)���e]�n�����Y^S��6���'��TfY�i8�h
�{G��}�D1��cܢ9F�w5���8�д118�B����k7��]�o*�v��}��V6[�]�� ��.���]]R��c�Ja���b�zϙ����|�)�1�
�;h}��G΍�RNj�۩1�I��sz�hG=g�-�m���&�̭pݳ��L���;�cf��~�~@#�G��4��8*��g�W���:=��B�xW���C��ֻE�I�r��ӏ�Y��_u�v��Elo`������0�`�)��LQ�ٳzdr�*!Pѷ�^Z�W���U�\�&s�v����=�M�����Z�5��ke��=B�C7��kIֽ���}�'.�R��Vm���n�~mˢ�c5��K^�i=D2ف5�H/�#�&r�F��ֹz��W�����SU��i7Ty����LF�z4�%��
`�s��h�B��#ꂒ��^N��x��7&�ϯ�6b���-�K�:<�:��WZ)��.��2᷌�Ly���Z��H[L�w�L~{�ꝭ�7V�ɟQϪ��40]:q����8��&+������;r��u��L�Y�!��q�g���}
D�$-�f8͍����ʫs�\[e3�e�ې��<r�q<�.���˦�0܂�꣉IZ�������J����q�g���m�q��<Gda�+��0�	wO�1��7
�<��(1<���6�9_t�~(�g(-#�}�S4~��a��@��p��}G�����쐹n� �Z�v�yu�����wY��Y��3l1
��M����}�VΕP�1�u�r��W�_oٗT����4.!ر��ξC�*�c�����\�x7����JJa��b��Vz���M'晙S�[�n�:?p�*��l����[�*���T�ꆯ��!�RwU�V��~�|6V]��]��Lao����~�0��W���v��C����}��k�����<ji1�f4�bKz������Zuގ\�$N�8F�E<���
����kǙ�ʽ�<:)dp㉗gV�4ݑ�^�ږ�������.4wFaFKci��h��m��y�\3^e׈�n��>����͸���z���<�
�����}r�Zʪ-�� Z{+J��]������N�������ǖ;)���x�>~gY�����n��?f3r���@2�����AD �{L6�uP4�V����/�7μ�s�0,�qW/2�YvV\hL��g�Zٸ�v�᳻+��h�;p	�j'����%��US�D�5�6�j�d����6jO��O�a����]��޶��otxV0�a$���P��ǅ�|�����M��/I>f��Q�սgp����3��	1A�(�#%0Í8h?����J�y��_^�l�� sB9a�/[�d6�����QA�Vj�[�<JJ{��W}�d;U7u��S�]��~���jU�����*��wmyUCeᗙ�
x�;�%��L5��f��L�[I
I����f�A�Je�E�ܘoUA�ձw(�HU��&�f�U�8�u����T�6'=�&�q-�|3��+�5&�W۔�Wi��]��xK�0="�!���Xv����T=�1&������IL�b>ȶ;J}�>��:~��SУ����8�y����� �Fm�
�$ v?���f!��^�̯Te^�fVf�lj�H[�����߷�G��y�w��q�"Ťl�]�.�.j���׻~AK�I�<Lm!��h/;��KU�ԕ�ҡ�Y�6��}���9E�l��i-���^�5�y��D[���Yy��~(nBn�t����̙xÆJ�;%a�ʒU�쓱U� d[����^5B�!����
��x{�Л��S�'[l�y��n�ps�Uܼ���n9�������t��<��6�Eێ���E�	����4f��xR���b��̭���Q�����ڰ7��`�9��٠޺=�!�t�� 0�	[��7F�r���Eu��s'F���p�8Џ[�m�5����l�"`4k[t,Oj�9�*���mX�]b�kf<s����sۆE�Z�s�"�1�Xu�9��ƞ�Sv:+����u/��s�E]��������4�Ci��Y4����\�;Ws����Y�#�a���RQ����l�Y��W�<���oʬ16���΍���Q�Nv�j��Tp�������Y��ǎӨ���.�{f����
k�s]�v���[�:|�E�y���N&�ĞJ�4�n���{�AW�ď̉���X~5�G~��c�w���!�ٯ��Mj<ݝ�mť�5�]xM!�4����;��ɾky-�LKd�P3י���f���ѧ�檹�f�Jؔi�)׽g9^�eM�T�
ʖ�]���j�ə\DN�ꮖY�	}��ڨbh$�h%�}��I y��T��~T��|�z�����N]m�9�E6μ׮)O9R[�N�~<�\56���=x��[�s�yש�kܦ�i�M0���C멾��4�N��I�����X�,��՞��m4���׹�뵣9f_��J�{�A��DY)�k+�6v������Ι�g����i��e��)�o�{}C)�"����+^���iYL�Ժ��Y������l��u;��g�b�Fc�y��f���,8�ƽ�j�����q�l-%�ɞ�8�^+�\�:~��"��J����{�ɗ^AC�n��#��/�N;m��i-�m�}MaU�����Ưm��h�,��7��n����:��/���G݅q����ײ���m��P�iĖ'Z�{�oJ̲�!�4��.��(�,�;��r��nLc��|-B���_:�ŭR���y�7:�Kg�i-��[��wW�'$& �a��`�� K.���]O��?,���iR��1���Q0�c��KSWd�i�;�:���T��p�y���e��K��vG�-ϰ}\)��y~�M�$n�!L�q׽g�3��B���hן����89*������>#�_Q���B�������;��z`�O	�']3oP�o�����Cܠ��ɴ1�9��[�]�*�����Q�W�N��k]�H{�p��11�����0j��h�*��l�ZN�(i����l�m��2��z���g~�H��c���X~��w�ra��uJI���y��Ԗ�ڲ\.�F�ߵ܊u�I��|G�Hq�wP�묵�?[�_�3�vC�pv.�wZ�[:��X�q�/m�ܴ�w[&հ������/.c���O�Am&>���kT'~���9���_}��9��08��v���Y�^^I�Z�Z��q)��M�����k��5]a��V�z�a�d�n]V�]��e��^Q6�[Mi�<���V��{1�;���Jf0�簞qѺ�]3�oT{>��%?^��0�۩}���ۺ潽��j{
f��ߐ�g���[����&[y�膵E�y����^��7�bq��O��v���v��@�ԁ_A��i�F�Ǹ�ɐ���R��7GY��n[�y��	�W�2<O,�/k��v�f�闲v�7�\[F[.�V�rnT���Re�N�/`�8�e���^ϥ{1���*��uk��m���R{['Ȱ�76����������b[{r(�p#1�6�g��,���%���jI[�t���-�I[jʤ�^���(Ӥ��d�X�T���B�e�Xw^��*D�o���C	Mk.�nE��l�X$o.�7�r��M��m�BgZF�b��Jq���s6��A��v:W�����(;���Tsv����IX��E�L�]DU� �:�7d�\��Z���F�В(m��'�\º�*U�U��mkm�q�2����f�w|��g�	�[��Ԭ��Ec�A�n�'�G7�)G2t͢9I���L������ތT͉h���z�-^�u�
×X2eZx�36_��7=Kp���%6���Vm����H�8{�;�bI����iL���b��-��W��r���|��=i�
�=�3��uo��[�++D\n��cUu�XՅ�K�8����w��˽'6;P)�v+b��+y�_��[�&��T�����pG�j��*��kRL��46�gLw��!]&�F����3/g"�[Yۉf�r��9��>*�^�l����y��[е��~�wSF�Y��M�!A�|A�}n�,�`��7<mg^U��r��t��r���9�V2V�1Rpٮ�{������|unD��絯j�|��ߊ���?��AH"AH) ����Xi ���~�~�D��$��P��T4
AI��D�
�6��R
CuDaIU ��H"�)���
AHg�����) ��$��R
��!��
Af�) � ��RAI�]R
AH)�Eg��9���^Q��]�� ��) �9U0������AH"B�) �2�D�\����$�UR�R'�T���1���޼o`q) ���F���R
C*��RAH)��� � RAHeQ�M$��a�
ACL��H}˹=�=� ��
H)H)���RTAH) �v�i ������
AH)z偉H)�$���"AH) � �ղ���o;�\ʯW�$>� ���M2�
Cu�՚ ���R
C�D��R
r�bAH) �2����R|�I �q%$��R㯘��N4��Q9�mG��:zɉ � ��$�*�(�Ì) ��b�R�) �2�6��
Aa��[)����4AH(u%$�j�) ��$��Y�%;`e��D��Rm
�m2����m�l����3}7�?%$��R�R
AH)�!ʠ1)���[`P�R
A@������;D���R
C��ښ ���*�R� ���R��9�,��R
CUDʅ�%$���
AH)�_~���$8��h��(���Ii ��7tAH,-�$��X[
Nz�����Pm%01���Yl����=w��o�s���0R��9�nz�GV�:�vE����y���$�/��������6I�̻R
AH)�D��ƒ
Aƈ) ��UI��i4�I �D��XX�߼od��R']h��2RAH)UR
AH-�+ ���R
C*�,V]$?����b肐P���ʩ3����4�$�ƈ(��?T- �7TAH)iI��l�$���s�7�
AH){��el �D��Ry
C�=tAH,4
A��) �f����C�D��R
A����@RRJB�
b2c7tAH.��R�6�I ����)3���
A�AI) �S) �/�ϫ첆�L.��y�
AH) ��
A`SI!uD��R
B�6j�����II��D��H,-�$3��tAIHRAH)UYVo��w^�k7�\��|��R4AH) �>�� ���R� �U2[) �;�{��AH(m%% S%��p�
AH)�Q7�CuD}�bAH<jO�L6
AI�9t>�[�
AH;�e� ������ ��RE��� ���.�תZAHw�d����P��R�~�R
II ��
AH)�j��h��R
AH)mR
AH)�$���R
CU��H�����lk1]�R
AM S%3�D��˫H)� ���RU%��
AH)�m�R
Aa��\1!����{ ���R
A�D~d���R� ���d�]�o �W8Q�0���IIUX���AH)�w��
AH)��j�) ��mR�[.��=���*���j�) ��CvPW���H)!�w�w�
AH)H��AH)���ZCUD9^l��R�l�
AHr�
��bC�D�$�����&���������RTAgY) �6���
Aa���D�� ��$�MR
AH,�&sYc�_��3*��mk1�H) � RA�D����i!��
@Ĥ��R�&����o��}�o����aI �.����I���i��󎀴���R
C�Di��
AH:h��Xu�$�wD0���R�$���R
C��ݽ삐P�JH)�D��Ry
Hj���Xc
H)
��)1�6���Q�8��
Z$���tMԤ��R��րRUaL�u%����(��-) ��)!����P�V�5�{�j�3uz�U��2�v*px�a[���:J�7�	�B��R�>w�}F����S[tV����_5����><��Q�M$���o�;�JI���
AH]Q ���!���� ���d�l���Q@R
C*�RAH)!_h���7YyC��f�y��
AH)��v�aI�߮�
CuD%$���T��KH)�
H)
� ���L9ꅤ9~��삐R
AHz��βRAI�
Hj���R
AsuyD��R
CUA����oz�{���N�f�� �@�T�3.j�j���,M0מ�wZ�i��y��Ȱ�7�Ò��-���W��<��=���.��#n�Ek��$"�5���k���n����5�ה�9f�qw��1�+�y�؍��`������[�eEw*d:d(�l-d:n��H��5�x�[0��[��
Hn)�(m 9�K������~"�lt� ���9�C|ү|"��"������۱�ȑ��F��^T�T.y�~yg�P̲y3xmo�详�l����Yz/��̮3Da��ucd��Q��E�jES���"y��׶����7X�H�]����O���啦�W��G�V�����l<�Օd�IT�]�&xi�\�����d��t(��n���u�}f�3;{���Mw��>+-�9�
��UN�šn�CkN_��4HkU����u�J��w�#I�jmu���o)��;��j��Km=X0ګ�Zi渡�w��~�]��>�]�lE�rݲ;�jS�]IyU�jW���>v��g��6�rk���v�����z:)�^1��#츀���'�ϝ�Quhvzd۠��=�݅&���f\aL<�S�=6M���a���k��&��4cX(�n��GV�ذq����Gk��Ĝѷ.�gz�r�)�kc��K�A�7 �v�f���Wf���[���Ǝ�G\�Np�#j�`�t h&�Y���qi�#��G��ūщWo�D�������i/%[��E��R��Wb�#�J��ݾ��ؒ[�NW
p?5u���b.>������7�V&>,�H���5��nT9�=�jg`�wQ���u��,J���;$���[��^M�x=ڦk;lu�#�\S"�^�r�?mJ��&0�Ɇ��3�ܝ*O_�:�^m���~u������5Y�.�ۙ�����hİ��J��0�[Ҏ텵
��ɐ����6k�u��.ҙ;�~ц��&��+ɱ�co��𦢤�X��y�$���$�<��2�r6L
8'd��Q��E4¾XR�|���L�{�_#�dh�]A��+���f�̽��g�u�Vo�ѕ����iwn�1x��$�ى��q����$��rA�\��%Cn'�Rx��1Kߘ��LFY"A#(F�pc>�m���ط$���k�ݬ��ؐgD��ݒ�T�Y��S��f��m>��A���D��L�J(q�8�K^�2�w��t��|�͏X����;G	�8tx���W��b�{���{���mle����˥b�"f�Y,�S?W�;B嫦u2��^�S�-����RݛSC[��>���ٲ���IXN��j�o-Mu�`:�`�)�m��P�%����o�1iwR�3���к->��S52���Vi�.��� ����zK��O8c4��E 
�z/�;�6�Y�2a���T\��1�#|��5�/�� ��=c*	n<]�zh�֤ʜe�h#B�_&�)�e゠e���a@�����үIbP���%����zO癑�re�)^mj�tS�����7m�7Ȣ�J�h�$D�a �v�q���2��cQ�FK�0�:Gm�9_==�����hd^m��Ǜ�:�i�C�]��z'��onQ�b��İ���ܓ��v��u5۲<��9^�Y�(p�_�"S7Xa�E���с:��j���8k/�y:x[�a��In�=�Xn���f{*c�	�U�i��S4��N�zR�z��,FD
"NG�^Z\A�p�Jﲲ�5giXe356vZ�l��0�#R�@�j�V7�]�6��EV��_hq�;y��,��}�����֑mgG�V��*�z�J6_g\"�n���;z��3j
��v�o��i��9͗�vD#Nj-Ӈ�C�26S1�L6�a��b7���>������y~QD5[Y�u��������53v�v��k.�f��̸��|��XJ�d04�m�jk�E��Rʏ�8b\X���]#~'�g�Uʛ���n���F����S�5�μ}�ٶi�_=$��h�ݠ�c���~�p��٭��[��g���η(��#�����,%��6�8��6�'+��0��f�p?m�#}�`�l�R���10�Ïy���������ߖ�\ض����#ه�,>�P���2�䁍'�Q���=,P���F\��8ڇˁ���]e�%��q�:g)Ө��up]�b�U�U5�����3��A�(�����<&��Ѿ�ᙜ�������~�YL�������<�9��t�{�n��Z�n�0��T��fSzxل�����Ħ�Fݍު�\] /�v����as�mt�z�(ӵ�Uh�xx�_P"��{)T��6�s�/B. :Tͭ����̾ě����j֕+nᆉ��ד+q*�"�&���StU��{��2εx�Oi�1X�;-�p��$Ъź��ӞJP�vGWp�L�4wv��Y~�^�N�ykPy;��o�M�y1��Z�����aD��[�$��tlh+n�'a�ø㵚8[Nټ&M<{���`�6`*8��8k8��~�1r�K^�ټ�z{&}%<s�_˗��Y.����9�8Ǟ<u��M:P��M׶kx��j�F1���F����T������}��o���_׳s���DU�5{όP>'C4I��4p%Koi�s����W�^��o���ߠ�c��]��f�T�^y��OgCQ�Sݪ�l9#����<d?�Jhc��S�K�>�q.M�2Z���ʻ����U�\ӮP��WC`2�m<�[b���r0��L N��5�l�)2E�D��pUj����f�bՕ�h�|�e8�{t`U�)���H����*ȱ����e���[;B�w�cp�
i{a��)Z���V:��ٳe�q]o��n�T�Bd����<+��S������I�s��m��7:ଡ(ޟOJ�(��cDL'LY��v����]q��S�n$'��ع��;�ǋf}z�rh}2�.�����zM]mt�i �pt�8�6֧uJq4�	İ½1�q�88=��J�#��V9��nCܡV��6��k����N�,�h1�oc���\�gu����v�)Y�*]v���b�>�y�*�!�kn�஺Ս�Ҡ�mv1���ȼ6Ѱ�����9��fF��j��]�[n2ŮE�av碫�<�s��Mq�Bd�(����1E��s�L�������ϟ꺜�{�^�G/����cai�t�Ĕ���	�;}��Y�x���I;`O���"����14���D���*6��չHz�:|\�=�4r}v+0t8��u%���{,#��s���bf���5I4S���pXѯl�t�O1� �:+��!p������2ɱ�{`�n�R�B.�}~��[x��OM�����I+TiQ!U��3��_8fe��%\���:��k
ݼ���u�Y兄��-|(e�*��2eÌ������g7�3�󜱋0vKĢ�p �e�@w!�����ڗ�#�a��Cއw�)��2ԈA��t1|�2�#�'�Dc�Y�ض+~������L�����(ā�#��33��c[�u���A�ػ]���#�m�gV7#\/[-^���`�߭�&n�<��ng ��L��z��t{�˽�;��y-��=���r>}d���4X�@4��|�޷i����YZO)��t44.��L�,��űJ7��okZ�䙱�`���s2�ޕV{�r�9_k�.Ѱ��T;k+�v�U�yz{��j0vR���Ȯ�d��9�H��C�s�n�;ÒL���`�^i����DT����t��/���Q�}pnwiʝQv�����vp��<1�����чʪ�Acpk>����`� ��(%�>�&����3�fr{����ے����ɺy,-�gF�u�t̡x�B���f
y�%4!�=�������7����y��$HKi��I~A�eg�E7��vV�T�P7'�h'�+O���r/�{r�9���g�j-j-yY�(]JP���s�S��s�0z�X�94��������F��h۱	��\�˜��Ů���&���V�a�Bcq�>0�wގ�%�$B��ǡ�2^3�ʇ���^L-D��QÙ��\�]{��e�V���������FRt���ꊽE���B����j�u�![1���7�2~��c%��Y��Tz�rY�"!�Z�Lx�nf���{���~�-s��&�otm���9���<˿Ds�ҏaU�od��V`I�Ǟ��eGf�_l��w~gs^�����u������Ն��]az���KE�����F�-T�(4�V�I^�&������oLôl�>ʞ��L��=�({��ٝ�E�*�f�h�v*��#�q'f(xT�`�uy)�6ye�S�
-����$f7�����%���>�/,�'=�Rc�)� �Jך7Z�{��m���.�*e��Z�]��n��/@Õ��-���Y�� ��˜�B��@t
c8͗�w{�=�mH����U�wUo-B��u,���oY10�_f���9CIA�˗�ႝ �*|R��&�˕=}҃y�7] ������r��M>��&�V�+����[�z��=��]C�b��] ��a���p��%ɐeW�xfu藾y('mGl�]_�u���=��G׍q��������/�Ksn�"yX�M��G*�&e��8(�����8os�zӤըW���=�r��+ř�0�"Z���>��'OI U�E�s¯Fk
��ԡ]ו7��}h����@�X���N*ɵ={�����V���3�V�oY̼To*�ވ.֜���[ׇ��,Z�P��X�Tn���ĉ��NX�<�9�9�M�z�
���j�:��/�e�gs���;ς�>��5*v�����՟�F��q�ѽ_�h̬j��p��ZY���cT�6��h̹yԼ=c�A�qv|���֘�=3=�vv��NQk�[���%�s����g�����m؞r�_�ף��Twu������J����	2�pr	CL��R,ҭW=��zN����=��Oxl��J�%I%g�tTe���%ϰ}�}o��hn��wg���n��!K荠R�՛��>'r����a2V��qdY�79��{�ڤ�y�5�N�1�Z����yri�q��O���%԰��h�R�����nF��5�ܿ/D�	ء�I�N~G �&��w��M�=���v�4q�R]C!;�*�$rJÑ��B$J�R�YAL�~�Nȋ=�eA��l{u�p�����[��M���Ʈ����3�5��W��g+rOZu�ƻ+�'Q �|�N�����h��A��ދ��1�����s�)>�k7����(t39+��c4��5�swW�t�b�U�k�h!��J��lM�ط�Z�PS����͹���u�q���2]�E��jV6�5��E-ؾ��6"������Xب�^�(\\�������B����#+��ԩJٿ�o|:���o������Vj�ŚX�i��Cwvޜ.�E�4陮�'�Ly7�/	�u��a���#���>�K�.�=� фK��%�TX��S�m�u.��U�B�c���V�������C;��e-��Sw{H;٭���e�U����bU���6��׈� 8�:�;{8n)k޾�'�5��S9���X����1�`"��gZ��zm)�H!�k�OE6��*�s:��QG<���ܖ`de�Y�v˲k|rhEf��o�d��~R�|[7��M<�3TF��*������H���C�ܪ'��Ǡi݊ݕ�mՍoj]]��KY�m�1��v��<�۔�ߎSٛX�e��7����S��$��qQy_ekF[���3e4���jnG�Z����X�C&�69hl�oفR�i�i�Q��y�ѣ��Y2�u9�v��Zt�qֲ��Rds7/�"�;�����&�2rk�ed��u��	��3���Ez�������R���6b��/e���a׬V��,�%a����wʸ�8u#�|��6�x2�aB�ޫ�ד�wHv)�VA!�X�Wn<n0GM\vԾ
�V�fM"f]v'�Ƈs�. �[ڔ�k�w6�dM��<:5�紱3%��aVc��qoGnۚ_�YA�lK��vb#M���tR)��/;/X���u!�F=�nq�E��"�N^���X Nk���C��o��=��*��v�aN]��]��<��ӻF�p�rE����\�C<lz�n�u�H�n�������t8��q����{���<pەv�erѶ��qf�c��ݭ��{$�y6�׃���)om۫�&���2s�!�nzLݦ��ܼN�S���]�=v��9�v�;r�k�������9�c�y��x�m��ຏC��-éW��v.:/m3�Gn^yd�zS�����.�W��u�e+v<m����ʵ&6z��*���9�tdwb��j�׶:4�EMm���B�خ��t���ۧ���v�]q�C=��ɫ�fz�:-9�Z��nʝc���6�vsk��Z�y��an]'<�WX�mv0�Wj^+q�osd��a�=��<���z�WE�I�ݢ�vnv<�Ix6"�Pܒ:֭W�v�n�ne�y\s��]��/n�>H�mu��a�'B�r�vXuٌ�ї��nP���%�*{&�\\sN��7\s��ڶ�Tqkq�<��ݫO����g ��й��	F�t��̵S��� T��6�8�V;v�7u���t\tm�����!�r��]:�Gj؝�:v�u��x���Y!�cu>��esI�8���ma+t�g��^��ʠ��@"�w<K`˸��7�PZ:n�;Z7n{nGn3E���鹻�ݺ��1hm��vt��:^y6������q7&`m�#������.�u�x��
'IΜ�Fb;;���<n�c"��G]�n�;#� �Ӑ��y���Q��c�أ"S�g��A��k	�^|��{ ��w6��cG=N+�Yڽ�a�ѳ���ݖǄ���- cE{h��ú��}������㦈�u���䵸������B����q#Om9�� �:����Y��<`�\��U�b٢�um�b8�9�`�],�:�et�6�طV�zݘ�y�wf��ð��u�8pq�^����8v�Zt���Q�u�cm��)�<h�U�fQ�A�gs��9wG�뫃{�A��9�s�� ����Y�x��Z{m����^�b��]�y��6ʽ6�9���[�=��v��q\7�ۅ(�Uc�k=w���r�>��N�,q������[z�3;(lm'x��}ó�%��ۀ��:�{���/h7���I��ϳ���!����<��������ӫ/F��F�l�*=p��Жk<XL�?)q�^�sn����{+�3=��>`�3a��Nՠ?K%u[��3����'�:�����D���������J�s��k���~.�M����;o�$��f�; C[�g�g�v2��U��8��!zkͨɍtGQ�{���C� �;��P�T��Ѝh�݁�Y�&�Ne,��Æ��]��́����e1��4�s���FP^����v�b��#���A���n�A�d_fI'5|�Gss�އt��^m���������<kb�9�1��L]6����b'�1�o���7��<x��a�vX�s�ɮ^f[��VP�/"�ǎ�v�V]�w.�9ɼv�y��̄ZgS���4�H߲ˤ��
'^�=�麷�ؗ=�eo��l��ޒ�������o�ބJ�JF��}	� L�(pf��'��bW��ق��tE�]�s�ݗ�-�:
�)Y�S8iV�lT�%�I��+%�kF�4�m��[uo�a�;ඏ���[��Ir^/f,��G-�j�};#��o(�K{eq�a=�Y���f�hF�.�>5 ��I�w0��Q�Q��V\w|¨��Y�f>Vn��j�Xwx�o�ߓC>�`o����n�=�ss}��ݔ�J)hh��*t�M�jgeb��cz���u4�j윚.�{{�]��&jWW^
�|���р�ѝ�@u}�����_g��jޅʂ@��%#��"ה둻6�z�D���"��w�]:z��BM�g�y��{/�^څ���v���j�F���a3)?���Żq��a�ݯu�M���Z�-;sq�W�ŋ �!�'芈0%���nAٓj����<grx�e5w}=���%i�ϣ�^*=(o�?>�S�W�iS���g�os�4�h�B@���FwQOܸ���f��UJ�3�[�2�^5�)��w������V�֥�n,���4�Nŵ�i���G)Ӥ��I��l�q~.lʙr�m�F��FQ5���C�7��p�{�n\�����%�pX3�Q2�P��GDYU�=���cde���� �	a,�����ޙ#�MnpѶ�z4�hj<��[�ػ�ylu�i�XX�<A([8AMH�W�+	�I��>�o���W@ј�ό޳���x���I�1��j��V+��2T嗸݋iW�oD�� �%�a�����y�3At�Z۠�M�Eed��ؓ�2�9O�8q~o����;6!F#ޓn�4�/��|vMņ���]��;E� ��x�ѻp���ޗ�c������ӝd��%"�(4�S�Am���rRjl�v�KΎ��뽬g����8<kTu��=�>�ќ��������`%����v4����)ݾD᰸��)���qU%װ^�_[��ceF�f��~ȧh�5F��x}e
���!A��)θ�F��v�!}~�{������| h��Q��(�l�w^�3N�%h�[chEk>�+��H����O�pL��Y�I�6K���?%��4��j��������R��Tp�˽�L���/?o����q���gRB�@Dx��u]��J���ϏF(��o�)<j�e�6$��s�良VU��f�W֪q�Hnoq�Ա�^�=sa?[������ڻ�eX�9���,p{��<�w�iYw���+�6ȁ�qr?� �j�������T��B��mt�[Y�lc�Z!y06�g�"!����oz3��4wr	�j�����#�8�`�#*I
��
hBp�����um����ۜq��0/��H��W
9_������~�+wM�W7l���gV��s������"�s����w;u����O��y[�0A~�����9����уEա��ѡ��")wJt��CzwI��jߘ�w�N`��s�,��e%�ftԖ7oŦb� {��Y�g�g�,�6I����^�{�˨�u�X���+��MGy�o-���5��5s2��3���$�e!erP���c}+����x��;��>�VY���W��aJ�zۛ�֩3}��v�ad
}�T���L�l���1f���T�Vfk�}��_�c�硿�i�����<n��}��s���Ʈ��>��E�\��z�J�S��d|C�j�YY,����c����ס���ڲ�
@l��C��:�y<�"��Ƶ��ue�����7��r2�ţ�gfL��R}�*�=�V%���,�`��C�#�d�y�#��s�Z8^x����qлVV��0om	��B�;N����nu]�@p%tn:�n
�O��5b��X�vlIq�6ܛ؁8��v�G1��rF�kx�w�
�;����ۅ�^��L�1��׈KP�@\��Z�tJ�~_m�Qc5�X݅\��zp�΍�ZٲE��q�seD%ti�M��	C�7���0أ�mή��-��\�8�Tu/nLӱ�'�<�P�2r�X89^����[\�4Kk�_�[J��e�U�b��kF�q8T���՞�'7�~�l:�`��6k����^�z:�r���.��h���M��� �8a�Aei��^5����+{�Y뗜����ю�=���9
ʜ���F�~�DO3�s��pR�	�7OFŰo�X\$!��,��I��յ��ކ:��*�u��ʬ|i��8�陮�9�K�;�,��%�W�������P��9�gqѐ���43^C���D�ee�[;9��^C+����!%o~����߮$�� ���+�2�U�}��[;�v����ەގ1d$��)��[�,M��I�L6g=����B���<n��$q�bӞG|���D��;W�)��ϳ��/7��J�8�[���oW|��)��Ϋ\=���1P�X���oh�v�;/6��6z�rǍvUS��]F�n�U��`q�Ͳ�����gh�W�G;�V-=1�ܬ"*Ӌ�U'E��C�V���~2��g��˗�R�ܕJ�lW7�ω䎐h6ۧ��sl�;Mw
,_�%{G#��R��<����Jέ����W7���r׬PB���s������Z|�=[�bU����6����g��fGLV��;5
�c�!���Թ�;҂ˬ\]�{�����k�v�t*]R.;+�ǹl�ڴ�Ȍf��*]��;�n�Y溑��
f��9��!�+3E��s�W{{+�Eڞ7yo�������(�]��Ъ���1bg����ں��[
S�b׵�W���Hd���	�%މټ&t�r����<T���DCO�e���%��Vo��Q�x�
S����S��p�y��e�� x>+GCgd�RlH[�]JM�e�I���|fzy�r�>��uP��j�T͓z��Zq����^���϶~E����4��{ύ1�����x,���/zd�@�@�l�t锃n�ۭηnz->{�ٻZڌ-�����v����Ϸ||o���i�@����֦�V6��9��H��.Tټ��W}6��N8�n��Q�Ph���7�w^t'���z֏b�D�x6���v�ʠ Ej�J�(��m=�Wz����`�Ls�u#��#Y��,�� �Pp������1�L�!�L��@����������F*���$1�N5%߽�,)���2�_V�ŷ@;�7qը���4���:�y\铞=٘7|6�t�6c��St���������5-U�lP`R�۫�v�=��:����	�`��xn|��&��0?%x�3H����ÛI����wC���%�a$��r9��W{��[�����6�y�^j���8�q� "*���;�ܕ�\�� Xwxų[u|�3��[�VF�m�z7I�����9`�}�
̟n�3��i�R�KT\��ؽ����G�g��!����;6 0�{߼ Ʌ0�:oӉ���𱌌
��ی\,��֧�ms�<�Y�8�(;[6��G�Bl���E�ݽ���v6� $�9�ۮ�2Y1��{Ǘ�n*�'P�V#[�=��d�_p��p�ip��^�4�1����곞`�$0��A�,��%�c��ҝ��ӹ|��Z��qv������a扫�_�"�N����/.����$(r&nrŞgݴ�CP�or��Y�j���`hDTJ��|b~��F��y�<�r��Do�ΑJ>j�����v �W=v�_�����0��9`����o'��`�%3t�xSm�.���QR����ҶG�n{w�o��(]��3������K#N�g�4��酗J�K�<�N���j�u{�t�!��,�p�nb��U:���&�p=\�^���5o32�tW2r'3����rɵsB��Q�l�g'	/��z�G�;�$��	-gA���5f�%�cD����B�c��n�SP����ze��wg�c"�T���w;��� ��^����Trľ�mʍ/��ݜ��O��*��s�i@w1s��M�f��u��I���&WW�3����Y��P�	����� Y���ggsJ�� Ǝ�����+*��p��&�����$Ӻ��/�r�ם񺠮�2^��9a�.)��W�+x<M� �Zm�����m�d�6�1Y�}$��W�yu}(��X�[x<2�:v�9�pٽȗ����	��ئ�~՝��_x>��j�e�26��"��I�8	t8�#��P_B�xU�I`�h22���A'����������H��e�J���r�_��ڳg*��pR��<��ON�7oi#Ĵ�T�I�[��V�^(6�{����?O���Pa�� �����+�j��_�����^��;=Ky^L5�.�pz�����9|�k��VP��� ,4Jk0
:	Ƭ���f��ں��� ٽ�W��fM�ub4�Ͼq�2���*���va���,;}����̥��
�y^:�����ww�q���mn�܊/nф���ބG��߳b�jޥ�OD����9�����5�������ކ)N;$�x�3���m,6{{��c��y�$�&�W:����w7b�5��ֈ��ȬF*s�P;<ޞp��]N��=�Jvq\�V1�&lW;k��ݼl�x����r;w���;���^����Ӓ�n�X��ͨ�n�t/k��wO&;��9@��O�^�{W/,���
C���\k����hy3q�@]kn�2�ϳ�N�<�A�jѶ�Ü:����JZ�s�8�{A�^ ��l�	�ۃ����_6岯����WM�]��b��=�u��k�3�Em�K�"3������w�>�X�h�s��!���a?CdB6��l�pja��]�t*aH�o��OVܯL�H�_a�L�@M 
nV^y�	���	[�ݼ�{�f��*��R�;<����:�>��rMuuX>L���wkt�)�������@��VV�'(���`���ʠ�/���z3�h]�Q�E�6s�������B�`U��}h�W{�<�n�I����%�b}���;�T����R�(O�d&c�C`Y}>��yx~攭Ӎ��pYl���ܶYк�^)Ws�5\��.���NUŀ/�L|��⬆@���R���P�q��È������^�S+�W֡ bH�
�j��-�v��L��3��(�nkN�WF�eu��,c.6;A��>����5b�*�P��i������M�<�X��c�[;� ��џn6��	��Z�P��g��R��8��t�����2*� WM��#�>%^�~	ݔҴH���ImӋ�#�u�լ�-���wL}�~�EG'��2�"��?I���"�F�|ۊ��6~s�ݓ�u��`sVS#���Ⱥ������߽/Ju}�s
�z1er��������v�SwwĊ�*Ԕ��
f������cp�t��ЫWX==��
���0��/;oyo��
�"A���7ݜ^�l�Ά�owf��:�����r1��R�8�FPP����]F��Ɇ�"�u��5C쭽|倽c��_�V7�����_����>����y;{(_BI���!�� (D1kت/�G�ɛ��[�.b(�5Z�����d5��bw�`�6�:�&�bc������g������)	y�4V����[�QM$*)%���[�!���HW��>^�B�/3�.��׏�/��
�*���ɂ�bĩ�(x��D<\_q|���U�Q5����S�]�ONuo����- "4�*�.�3�ͬ����J��kb㺳{%�����n������0���i����8���h�Ɲ��ܯ-| ��-u�6>����^�s:�:�<f�T���=�,͐��%:��aR|�Qv�!����@�//��H�4��|kTť��;<����T)�YS=��*pV3Oٹ��j�Ĕ�)!�
��0���n��(�A|o��v���$@��n:F�K�v=��8~�ї�ž�4'��6�X�:yV�����Y���6lY�Ħ�9�h	�]MH��5.%y^x:�Z��k��h�1Yv��V�x˃�e�j݋N���i,V΋�^J`}ד[�孜���2/E�r�b�&e�S��+=�sGV�
���y���!�rV���V����Wp�W��g/Lօf�gM��u�K	t�b8��:�U�W�\]-
��9�{�J��?/]��r�؄�r����&�ݵ������&{3:��3F�뼮��_6�h�cd:�����F���n�u�s����w_��.�Dn�&��Y���)ˬKt��Q;5��	�/�:b�Ƀ�ʹv�ŷ�i!�~nxh���V��H�OQK��V��^`��+��\�"׫��g��������`�{�q3{��\�}��+��j��O2��5ٔ�B�f�Ea�\=N����5�<�޼��F���W�m�����U�Y�pe챮�<�{�M&�G_��<� �
�r7���!WeCB��/��P8�������쬎FHZeًN �����ۦC����7�>������,5�juΡ�.�Rޙ�K�
�����ޱ+	R���9�1����Tw(m����p4�Ma��"NIf����v_[CZ�M�y��o��HU���;�}����X��I���c}1����o���3f�c��l�|�'8B�s��F������v�`��Y��v�,�K�	3�X4�yM(���	4���TW�i���w~��q��wU5����PWy�ӕ�C����i���)�2E2 D�$q�No�_2��W�'��G7U�5t�^-��K�z�Q&�|�)���L��`7��_�������ː'g���{^_<Dؓ�]���aZQ$d�	�mz H��k�0�i �4^]f-�����1'[3�n(Rwn��D��k��1G�ʟ����`aȥKq͛�-}��X!�p>��3�ē|CM!m�%y����mϊ�݄�#�혻[���۱��Y	"�����I��^J��A�^�M�Ϯ�
��n?z�X��Q �����/�j�'�nા��!R�{}Z\�dB��&&���"�b������ꀨ4�a�>�px���)�z\!;�b>�x��R�~7�v�������L���ݔ�7�E����躖�(y��U�l��'6�V�!�bH&�&h43���k��3S�P���r�B���x'	E��}Y��`����:b�Csx�ٯ�����Ā��\k7�Ͼ�u���;���m���D�N���w
�0�I�h��w4L<�|�c��9ʌ�Ů?���B�\�IX�D`�aN��׏�e��#�X��CRx<�.*�]�:�T%�"zX�5z=!�U^�i0���	�BUq��Έ��1��.���SJX �:4u�������0}�
�gT��t�-��!(L�v0�b<�~N��}���d�)�W�Q��������ѧՕZ8��R+�3��]����*�����~H�WynĔ��jT
�B?�E@[3�>JGWo�������j��ڑ�cGa[����.�� I9�['�>P=}������La�ȅݻ��t�
VϨ�\��TJg�wg��[P�3)��jm\�%��>Ŕe��U�r���C#�ZG5��WѸ�De!�GD.e�ٛ=����/a]��o�� xJU��Dk�?RD�Duz�ge
�BB����u�4q�C*�Y-cD(X�A����vh��5e�s1�Y���yƛq�f�g�ZW�^V������D��KA��Ў{U%+7
Gz���Ť���Y�֝�K<�}
�r�j�p�b��"��㙼£���"����W��?���5��f:�0��������f��r�1��(���6��S�R�5��yhJ���7��]e�9�I��x�T=�7L����b��T�߰�-�� ��v�g�T=��	>�مдW�9�4�½Y�B��8�[[�33�z��;y��x�$EAx#gK���	[/6��^[��CyM���Ǯk�:�X�ʼϓ$C^�[���ɻ�ڑ��?AY&6���莻Z�sj��޷�C�g�k�M����g3\r��sƵ��O������쫸�וsv�gf�%ɻ8y�o�A�^��,3yu���Ƅ#>�7-�{�]r<]=)��B���J���iy�8X�tsF��r�=��M��nwq�8}����HN����:��ѮϘ�s�7����6ys��홀V��1Z���FG[���H�y�mxM�;�uO�y��M/63���a�VsA���oϜJ{�������z��Q���U��Nf+�C�LW�ַ��A;��	���56K�Z~����`!33μ1a�RE8�y��J-B�f9,g�?(�>�+�*���iҭYT�-՜b���
�ب*+��FB����DU�jº����oZ>[��_x����uLP�Ċ��U�)@�lY����|����`C�y�ʾ¾'���K}}�N�=��gr�nѝ�7U��{�Z�"A��zL��=ye̞���5�u��G��Ј��#�@+E��n]��U�dxgd��>��;DT�vhuKg.�4C�>�������8}���>���4��U��t�ǜ�h��g�,�ǉ+5Ȓ|PeG���>|�US�P�p�ᕞu� ���T�]�+ol���ɾ�QS_SX��7�׾��h�K~���ۨoE�j��4sU��o_��@��$"�D��`�h�U�ܸ�F�;.���]�{7v#���&�݉��"R���gٗ,�W�P�a���;��q�����D���s lN���v�#�!oV����x�� H��|G2Z���������6��[ ���U��^�}^G�����.����h��R�";��]ܸ҃)Coq\��k����g]$��A�3��p��w�(���X�f�W���>ꕛwӑ�i�Ok!ڣ�+H{�B%rȢ�ن���OWk'=z8Pg?w�0�4fGA�#�FD�? G�-Wwv��52&q�3ϻ��G~A�y�J������?x�9���]�L���^�̥ɛ������K���8�8�rs�v�p�{G
|>�����v#����k4O��[�p!Sb#�u��w5�`
L�U��%���5{f�Our5���n���(�\����+��̈��Ib?20�P�������m�~��I��`[���Z���������/�<�0����d��>�*��z1>�DM�g��K�|
����F��</Wd�^Ɲ�HF�+��ͷ`�ц<%�0k;{E�K��J4�I"�<�&�~b�yda�P=:���w���W�W��A�q0y������VG.p��z�^�����ř�^X���G�'�6~���`��K'�$� �(��*S�Y2a��e�Ψ�rwq.��l����t ���f�o�#�E@���ɐJp��si�ۜ�o>�Xs�j��E�h����]P���.&Ad�)�+"~�0!y�-`�p�"ʉe&�b=S����L� 6��2�����#���cJg�tK�#����ƴ�c���ŏC뒱kp�ne�!J�[��8�բ�)�ip�9���xÔ��4s�E �Q��;�Uv�׬�VZ�Z�C���R�="��ic'O��O�qس�O�X�>�Px�1��O�+t�`Ǻ�(�����&
397g�~m��o���X)#�dY+݃�K��{�����R�����ʏS�q��a��.'}`�O�@6���h0o� �m|���)e࿝f)2s���_0�x�0�3F���K������R�����1���j��#�ȝ/B|��dlK���'���q����e���f�����f�Up=�=��μ6��'m��w�� �i|!���[Z�a�iC�!x[�;]0/����߇��"_F����xWP�6�X�~�(x_�.�\�^����4[Wj�<�@�lϐM�c>A��WAX�yҖ!������O ,�N�[zj�j\p�����&(%�/X�YCD�����I�}���sb]bo�n�S0�.��
��TjK�n0�$�����>7vFR�Z���o��/Pb�\cW|0�S�
��W�y�Z
b�D!�2��?u��5}	 [��Af��т6�F9}���dR�f�K[~�3��T�-�WƐ֮{2�*��w]��x�
L�,`�~W�D"k����5�X�A®���B�͸-e�c	�؜;,�p�*�����N��[=���8�IK�Rh�V���k-��*�jr�<���Ľ��L"mс�Q7ƸlF	r7 0�š���k��.����m���D�8� \��7]�c�+���U\���Վ�p�IKp��ȪB;����=���O����A��R�3�����A?O�m�[K�W�����ez$:��.v��*v��lP�{��2��;����j��`���>5��C1�89���TR�2�Y�Z���F�_�,�C�J$�&�����Q�B�J�!�Wgb�a �\��P"Ѓ�e�p2T�{��������1_hM�0�͸(��v�+�Y�����|�f�B�8�E����1�ZU���N�:�]9}�U��J厩�o����߾k����IĢ8hX#�"�G6��ܲ�e�y��)��-�`�eo'�I���>ٙ�|����t/H&(DH��"�'��7�W��F��R{���	�
2Tp��
��j���{cOY�u��f:���%k�s��g���G��b1���5:?>�or�ҝ�4CW��Le�||p�j��,��MJ��Ty+��xЫ6v�EF�S3�=����<h�h-H�#ϬA���+�y}Dg�>��ě[�p�aQ�yJBW�����7b�OJ4�V�v���)��ة�̠�h����աWS�������Ǝwv,ͧ��tO;��o�b�7�ؠ��L#Ǵ�7�;8� �'9�/;���Ds�9-�j�^V\'Kls��@�5�V��6��v�[���7	lN}�۶��;F��7r�͵g�nۭ!���o����nG��,�q�5�p͕zźm8�u�x1�QQǎ���'^�Y�:1�q�/qwj�M�g�4�x�a�z�ۇ��R`S0�rB�H���O5�\�v���36yؽ�lc65��t�,t�gm��]��M΃i9�ٺ��<�64>����v�����Lɕx���'�bs����¦�R����߁!DwL
 C9�J���t�@�#?1�;i�lN��ǭC��4�[�Z��kQ!�<����T�ʮ<Ą��-���E!��O�~����.�F�}{-w���t�GK��c�V2�d
�׊�Q
v@C� ������,�
�Q��[�{	�p�H�r�mQ�[��ū~d&���#I)$��_4�(��[���S��f3�ϔdB(��|&k�)�^�[�2՜K����Gw� #l ��:�ܒ���\z_]�(��]�Xp����be�#����QyPքx�{���v{2+侯
��V�&�r�ʤ�"��O�л�,|��mfx�/6Z�TE��B�6?/ �p� �03�~����Z��o�}�
C��Ep�����M��Y�~�Ǖ�}�9_WM�g�}ժv���x h�gL%P�Bd�T��������ޚ�K�։�>��NB8.z7v��c�@��2���C��Zs�zH5�6���Z7����,�Nߐ�>o��yW�nV��)OA^�a�b򁀸  I��+B��1;g��;DUe�v�� +����k��Y!���vR�����qU��_B���a����]���`w�0��
O����fP�U7��%w�#�ъ��[��V�N�����$��d��+��$J�6�^I�g�(���� �>=��P~X$����iR�tC��1S��/�����}f�mv�S�*]j��,"vV�������%&n
�����uzkM5�	H���WД����K�;��J�F�f�CZ�R��]{�F�B�6�~-��R4$�W�u{t|~�:�M"��_=4��H�p��m�`n�1v1']sW��UdҸ��ov�>�|���Ȇ��v�;�uX��B��H۷`X�����^���K�,��R�{{R˽9�q.�|�:��1�rA��pU⤜B����V~�0�������՟�?O�~��<y�o�p�bH��yu�c.��;��Z6x��	��_n��E�4Ey��!Z }���nPq�������OO�u�9�.�.żp��ո��&��79.:��v�l�}v���H{N�2	r����C\٣��9����^(>��T�Sb�B�*&��kBӂy�]��hVw&���}/� �L���ء�@�01бG��6G���@:@zױΒ��NU��&��n����z���R�U�ox����ZV���`��'-��꽎yX�<Q�E��J��#˂:E|�8�(�n9%�hd)�J�Q��뾱XF6?1�\k�(=�J�,ԧ����S_�^Qg�0,0%����yX]��-�����s�vw�$�Eokp�$�[�&��w�j�s��7�,�J�e{{�u���'ܜ�0��0"��� ���A����K|`�(�@�"���dV~�#v`����qf�8�+E]��"�������j`C5��۟>^ m�˿9�~ ���n�;�#�au������X��]��(h�,�f��"9I8`a'���
H�XSu���V�� ��6^Q��Jn�!b��g� Uc���4�]u*���,H���8��(��#�!�w���ީg�6�p=(��G'#�s1��B����9�VOHQ��.6���׾�]�h5��\&�nO�A����݆[��5g�n��z"�Ո�ݾ>����@H�ءx���{�ev	����OހQA�Wv�KH�_-�,����� -���\OB3I�)�妯yL7
V�W l�����ڋ}T��ψbD�:eʫ��EX��gy�e���f���fL9��d�ߗ��J{|Oچ�� }є�@����e��Z�i X��ޮ��S$Q6�X~��t��0T3ٶ�u��?q��4�2�P~�̲��/uq�b�Cw��uUώ��������RK�r�@����yT���/<^���uk��ە��Ə�0!�]vX�a�F��A��]O����R��=����C9!�zV�|�B�%(z��w+_Dc5��{���D>��5��p[#�{d�;��fM����)h�.ßOp�Xz����s���{ʲ&5��f-��PE��и�v0�HW*�X���ӎu�'�7��+0�S9�x���^��xTA(�PWq���N�V���%��ބ*7��wL4� C L$����ӽ~�'ոIXH�)��i�ݮ�T�^�bס�h8Jq��8r�v��&QEe&Kk������8��� �jy%�X.��U��a�f1��ܬ=B��,��4kW�p����tgj�k{WM����2*�hZ���㨠�*����R���E$Riyv�|�8���+8����
<�7x6(�_(j*��e�N]R�v�"_ܟ�^"~Y�F��?�{|j���>���1� �R.����p�L����f��q]����o)V/�[�V�t���V��NމZ-zCNu�5�BZ{��PQu�7���lq���F���"c�t,�F����ɻ[�L�IM�I"Sc<�z�UNɾh	�DM&�Dh������?Y�(�.�����%�#����KHp��8{�_.;���N�gm�r�P@�p��ou��R(�FD�t�I�dC�>�{���u�����[P0�]��1��]�и��>���u�ފ��4>B���^:D^���*_g�!v��iX/bXd�QK��� ���۹�)�t)��f�H�q�E2Ϯ�{.�*M�����s���-�I�3�nR�{��Ϊ�抲�͙�շ�4�(m(�P�������U[��Q����C}kVhU�έ�r�
ޕ�w�Z奻J���j�9a���}X6�C�ׅN�����J�[%�$�vq�uZ7r���*ya��YZԚi��x�#6��@W������w� ǆ���.��=Q2w�i��0��F�Ӕ��O*���it,�~p�ۊB�C0��vn7�v�Bv��gT�SvW��9�����v��վߥ��H��z58������w��y\�����P�nZ9X�K}fcņ��qb��4�E[]���\mA�1Xo-�fx��J]�o��[�+J��w���]D�K Q�سv��D�Lhyi�����rMH����i���`�o	H8���µ̩q���]��.	[e����Z�r��A����v��{�dBڦ	m^����wVf����N�M�;Yc�2K{|���f�N\�ݼ:�۰K��4��`$-��+sr�6@�d��8�WP*汉l�5���Q��s��u��։�o_+I�K@GDZ������S*S);F���U�*�}�Qwa���v�uVv�ϧ?��Nѭ��6V��8k�F�����tYc>�D����[6�]vv�Oe�Z���`6Qa��#0�f���ׂ+�fjv3��h�U.?VZy�xR>G`7�V�ݤZ�^���l��I+߱3���觔���@7b��w��r���]������.�Dv�yw��(��Ā�#[�'v�e���;=�p�\Z���!���#�;��eL�ۮ�3�����Nqq����1����m��­]�ānLd��ո�{�]�哝��T�[N���X�|�v�G[�ŗ��+��wU˚b�5�-A�s���$�����5��FN��8�˘�,�{g�ݻ9�g���ۍq��d�b��mrט6���hsnݧ�CͰ��:��;��$����v2��z���g@���w/���b�v��%��+��­�Q�B��x.gD��=�:;�"7\lv�uɜ�L�yÃ^��x�ܳ�c=���Q��Z�ƴWe������+�Јӎ��cV�@9=�E�6=�7�M���-ϡS^L��tn�/_V�;��ًO8��Nm���nk����Fݭ�6��1��یB��;p�Ys��O�6��u�[�uc�A��!�;SD\<+�4I�۶@�[mێ�S��v�^��ѻzV1���t�/l�q­ێ;�i�\Z����Y�������r>x�I�6îln�%��\�OM��D���ۊ��:�etb��/=#[oZm��q��qмvz��9���r�˸]�y�������]��@�f���M�/ p�����:��CF'��eL�RG<�m!���ȷY��:�]!�Ñ�Ǣ���[�����V^Uf��5v�^Ć��]Ss\���s�s���s����i�^��{y��wla��^�>�k:�1���<����cO�k��t��ɤy2N7��On��Zg�����ݬ��aG�۟n��kgڭ����+�T|�Ϩ����[`�i��G�!l��p8����p�E�ͻ�������9�<�n�>�#qݸ�<Ẻ8��k���czŜ=�m�&O8�M���c�"ɁzW���WIr���vK�R���0��%1R���9��*������u�jzy�:�^	���s���s������m�Ɗ���n���j��ԏc�N��ke`�r �s�em��3���^�«n-�%�ۑ���E�n�Lݽm��c>�]!>�\]q�}���^Su�� �ڬ���f�,Ovn�{M��q��jx�ke�5�)�1��ր9�-����;v��d�y�����s�xX�c��9QZ�u��hU�3������b��a]����/2���um�Mv.��պqu��i@T���?�Ns�����f�cCϡ�eI6]�R�"�C�%������y�h&�n}K��%:�Af�;9R~s��e�%֛���~C���ޡɃ!$�e�83oeV�����5vw��$+�k����@����$o�e�+jGz��#��չ�Y7����D�:#E���ʃ�X�ӝn���"b�್�i�e��NC`if7DS鎦����ϯ(����?A\)N�'�:��~6~U�%�+0����,�o���U����F������U��}��M&�7��C2|IFO�A�V�4;;�6�\N���ʊ����b�I�5�ҩ�p�{B�o���m���R��(-:���CW����j��={� ����`yPx4�.��BI�R���.�O��s|���!����Y-zWY͒�:>����6n�Yt��B�{�,��On�m���:F]} imd6�#u6����_�o��u"�pҤ�s�c��)��Ē�� On���'&�6|��ѳ��u�;ۦ�a�f��q���¹���:��Hȃ��+uꝊ���n�T�HIHV���\ݡ��J�hQ3���;j�7�����׻"L���-���ز� ���W:�vhY�&'�G�v}�4w��ް��W1B(k}�zF�Ԋ�V.=w=�:���t����2��3�fu�uق�Rzu�. �~r>\`�8S��{�Y���Pǣo�gҥ����V��WoL�a��=Y��.��{�	/)�.�`�x�#'Ƀ!��k�?n(G4(�?U ��>6>�_3���_gg�F�!N���Y3�&�LUov����<��\��P���C���O���@|o��.|�5e+E 茡�1|މ�s(�xV����*��~�?w���܆�L鱹k��ˁ��_!R�c�`��k�"�ڎ��18Z?c5�`������Q�7}zݐ�dBF�J?;���<5N�Nԁ�e��ڻ�݊��HZK�v��|p���-�זN
�::��8�h��>�-K�k�{e�8�v�v����p��`��:�V`]��[h������@v�$��J�f����w��* ����c�_!�4��9��bHi�����.�G�Cx�'�f��D!4J#���ۀ����O҈g��Z��
}Q�a��we�.׶��9= T�׍�7��M��7L,/��h{9�#���X3��� Q�,(�dJ��?y�Hm�3f��Ob��$��f�P�o1�RTS��J��ʵy��7�5���״��E>��T��<��eYA��:�wy�}���S�I_|�q��sW�Y��[�����W1��Nٯz����g\�Qݿ�ʛǕ��p�ꂦޏ�n�eS�G�sd����(j��r����;P'��d1�Q,6S��5�^�����)=����ײ3�zk��g�p���G�>�����0;s'�O1��^���[�Ouj�"�0!־����|	06�T��b���A@h�0h�w�p}b��(z���wޣ4�l���ke%�`V�i��To�F)���WJD#i�b���N�ve{�5��~�v9�.��y0����Q�����N�;%�w��E䇂�l�M���vj���}��)� 1���ެc��>���X���`��[Zx���#�W'��w�B������}���=r��w �ҫ��k6�}����n���l����LT��
�sU:{��7u��qfZ��-߰i�^^v~��\	�|+ϲ8h�ޫ�ul���ׁp�a���J-#�CVF��B~�������8��3���'�߻|�tݕ|�q�+Eo6oV�׵溙����p�/�2�u�&Kb�\�Q�$.:.�2�C}�J�u��,nol\�����Vל�@a�E�&-?BA��
��EO:#��+��p�=?K�{�O��ΰ�֯�����%�z4]�ݔ�+��*��	v�k61�$�i�+�B���)J��k���su��˛R�⮻WL�>X#���0���9��F4`E�!rEXx��R��dA�u�Ԟ��--�U�� ���(]Ü=���+^ C)���N��}�!������h��x1N�=���J%	0�
�T�|���fݶ��dǮr�jq�s�Y����n�ݙ L�$࡚�x*��!Z�w�V-~��,�
����- '���+,�9����7�22����bP�]��qW����G
f@��6$pP�O=NQ� 	
R돔��5�����,ÀّK��@<����-�u��s5��-��3W��xE��{�d�ĴF�>��f)���^��b!�XMŻ��`B�*Y�.�`�1�C�¡�+o���6+�5ON���u��|�k�6��8�#�;�ˀ꽗� \^�Gj�7�pH$e����^��i$򲢱P]��a�u�/�a�T��ق�b	�٭��?�n����q�+�,r�����3GՍ٘�wb�5'`$�R,�	�HM��`�?y�3�� S�,����~��8����S�S�ߜ�����~��S�
�# U/eS��3�=�d��@��{��nͦT���^;�9�w��{'�Y�]���������-�W�u[�2����6�ڻï�%��eǦX�;7�,�t�E�o^�ٸ4f``����p�o��ʝi�ې^wֻ]�u�<��TF�:�Y[N��=ѳ�<��z��9��;Stvґ�ܜ�fX}�<s�-��]��k�5˳t��n.Y�TnM���w�yㇵ��'@y6�'9��$��[kj��_[n�<��[�Ev�n��b��p��Ƙ�S�*�*^�y�N�c:�Z��ny�E��{�܋�I+a���<�m�qW;�UV�*ހ�m�Yݹ��BN:%cf�Ϥ
�h��z�L8�RI1>2C\3�_W�8H*+��tfb�p�x�<
��ɿM�����)���u�Zݻ8zڻ��,T�Ӻ�O�F⚬�E�q�x�y�J;�D���_�Bid[�,���ڬ �&=��1�(���j\&^�gID��SL��c:��v�z�	���W�f�Z������a߅����4�R�M���$�#��	dU*#�����y�m���f�7~O�!�������r��+.^mցwټ��i���i],�~8l��ha����A����Z�c�_��O��9�� �ל�_ܻ��#xa�i�<��8FT_B���F�Q���]����d�Bt(�b�r*��"�Ezʚ�L�]��X��˭�.�*�`ߤŊ���C�%/��vi��E��G�����y��f�R����Z�%_m�3��ۀU%"�z���n�m�Wk�m����=�їۀ��-��������������;p�W�O I4Y����ƾ�h�R˴��Nt���7ȉSn���t�f��A�(�If���$�p�A0`��b#MXaV����5�:W��z�K�
�7�h����KZ�FX�	���{���b��������<9]��L�q�"b[沑.r*OLwy�a�<r=Wn�`Cdi�^�ԏ���k�g�tV��w����Tlsݒn�b�ξB�.��� R�Q)�3�;K�a��O/��}���A����o�8������U�FP� ?rܕ2��ع��W�.�v+QGңF�.S�ƛ��Q�����^�lF��c���a0��6l�;��1��*p}���~|��w����e���{��xi=�xwo39Xy���6'�U�0$;ׁ��<\����"���eRW������0d̦!8mSCa�-w�L���{r�[7Hg~��K�ieΕܳ�M-,�`���^ֻ��?e6���˸�oq`��ێ.�v��s��<�6*�nǥ�^(T)-�Ϋ��֤��>`�;��̛�f������_	3�_aaj�S�B=���w{�u�ӆC��v���A�/ã���"�N"�F8k9~�&��C|��>57޴{_Vb����s�Ujx��Hдj�M�+���w$ս����!�����f�������>)��%(����f�:~�������͹�/�G4��4�,�͎D7�5\�9ؔ��馴Ej�ˡ��V���t�mF���@��r�G�����w%u���>51덥��F=�cY��U�|����ѷm=C�GzdK�}��M�o/4r��&ȃ,O�m�ܗ]�i��"��u��{�/پ�7�q]��zޖ���6��8���� 7��@B��f7V�ʳ����� �.�#��qV���'P௝�cqAQ
�	v 0%3�Pav�Tр`�a#\�P��ǚ:�����B\��#�b���$"ʥ���h1E�tG'Lbx`�2e���Ge�\�N��f�Wc�۰�7m�8�w9�J��I����	=h�y���p����q%�vMv�l:}�媠PU#�%���'�ڼ���ܜ���\4ګ#�y:��=���-Iqdo]�V_}#������l�W��d�$$J���0�}.m�<zEAФ��i�o�:���M�:�e]L��MQ�����u����3E�U�磂��t�Bm�,YA|���d@Ē:��ɌңP����:_�h��H���՟o��F�c%�Q$��� ��׵x�5{�V%��~����Y��
�ڎ��@�|Bϛi�$�$vR)}��!EW�n�>�z+��s�?�2���}Y���C�=E�M`C�>���������<���g����f��A�(�2a�G�
��+�3�7�k"�uFR��7����K2��Xu��խ�fVCvuײ�ګ�_W��zCY��.q�E��P��e��]XV��6�J��pϳ�!��~���b�7RWoN��Ś~�k��<�/W��� �����v+�# 3b���mi��h�xݙ�����L��:|HF�#��M����;[�I��l]��p[v��n�D�@��3�Lh�:�в;���@�Ŧ�0�z��]g�E>[�:�R�!���lp�7���ͷ�ܩգ�V�f$CK�;�f@Y	8d��f=���J������G�Ҹ����!V*�QW����b�����?�.�s���r�<㜚��jv0;�M���; íSFJ�)�f��$F��v��������w0R+��C�_�Cu�F��禞�.���wj�|����q53,0�C%e�=���l� I��p+',�;��˿%��8�1�����9��wHWy{�FJ�t�_��U�3>gR�a}�Ч=�]���y�KjT�Sڂ��K���(�:��KM'"���+��4�I��=���Ȳ���^F�{��eb����2����_*��`��ٔ�]������K�<�-��N+�:bhOY/�U��'9��:�C�ڽxAx˫��HV���n�:����SُE�N�	�75��jƧ`;��*=S�L���#����ߪ�7W�w|u,��c�i��/boI��;h=`ݫ���:7e�rn�L`+�\<���������^��u�����{1�.�q=�U�i�n�,�i�ʪ)L����:k�D.��ˇ���n0�Ѷ�n���G�3�ʐ����q�%g"��ݓYB��nkm���u�v�)���{<q��F�M����.�t���d.�=q���m� �c���.�m��e�-F�p4wHgΞ|YuSv�g;�2��;N��1���pW���N�bگ����o���j�O/;��u�,U�z.��wJ-�϶GW0J�9�xQ�n��\����"�_�_o���6F��q��I ���0����{�@��
+�sz��s���,�5F�  G����$y�F����}�o��ϼP�e�o�n�W��!��Y��g2[|�L� ,�ӫ�=Ei�G6��V���S�h������El� G�8�����>b�״X�}�����rr�V���K�0Ha@ZqX����&ލ�(gJ^������0e/��-��n�z$��VR��ꆱjd1Z�at�z�yU@�܀8��F���#.BTE$�YZ4�A���,��C*�⎱Iҽ5��"�����K�.�u2�:qt�|xaB��od���'D��q�rR��v8+�Q��l����S9#��W�ؗ�������4�l�=?PI�5�����<������n�^��$0�h�;�U �'��L|�O���B�-�I��-:��+O��v^Sud2Ew�<�pN��R��UF�=��N&0nkӽ���nWt��G�(��*LT����Q�u��Ʀ2�i7F>�R��]6���R�DCyչ��˗k�m~�>�#n��#�4|a�ڧ�#�[��a��bAN�Oz7lgIε���Q�~�8,u��1�QX�2�O���'$�H)�^��l]�-����2I����Z*�f�-�������H�y�Y�-�>�γדc�����78R%jl5hbrKpb����Yu�yڀNf@D�E7e{�x�d2������ݻ�PW�Fֱ'��~ٻ�omU_E^
�<��|�H«6
���>�ǒr�N�����nb�Z=n�I8��r�@�> �[i��@��!����?��D{�n�����@w��[�	�P�4C_!���]�i�����-�9�v�r�s�N����D�{v����"(ɒ=��#Rf��,��+�<R�4t�&�|��[nv�0�R��}3y��x�P����tV#�VVb��t]:�t�!�ȰXL4��Gb\b�c�3�_�VP\��b�d�e�f��E����:Y��c+��{٬������C���'2:���k�;E��a�[����m�qe�^ �m�V�����B��¤G�Kf����e��v�.����n:���
7�u�$�+���p��/ׁ
v���ʟ RG4e��v�o���)��-�3�u�Q"��of ��_]%�-Z��S�츺NF$7����:M2�s��ъ��Z�ڤq-%���sx���Ν�ۘZ�jߥ�F8�i��G�N�6�fB�j/]U�����M�T#Z��v�+o�)��Щ�fjg�-�����b<E�v���Ѭd�g}����kX��-}-�U�b 
�Ӂ�a�ł���V�-����l�_O��
�jU��Ǽ�����i�˹3%h�j�١���{�"��Ŗ"�Z�	a_�^��~�/!,�L�A.����C�QZ�� l?��U���X"�nK>(��5�#��7�?n����h�����kھ�`8���OE	=��`vhЭ�)6�U�6��,!fA���CVS�5���g��]8��d�9�\C�n�q����b��J^%)�@���(��������ǹy�2�+g����e�'�<�����v�ngM�W��z�A���^h�N?*�z&Rmry�w:^P�e��ׁq�b?���9M]Kؐ��#i`�;�AХ
����b�0�e��+��S�ټ�r��b��&G�f���\i�'R��c�D���ᾗ�W��c>�+�Pީ���ûZ��Y�9\;��= �ꚛ6�<͸/���f��T�e]o��\����ӽ?'��R�ҍ�N+��R����{H1�8�s�`�:n_5}t���A)��:��k�t=�Mjֵ��`�CY��?Y ��1�J��ԬϰZJN�)�ϼ�[�Ц��mԼW21:�n��Vu������Z������F@���޻�;]-��aT�̞�Jמ���մ%`�����~���/-A��I$�6d&l�N������'�|��$wN �xL�tt��%�����i�v��W����y�˕�+=N�c2�����\kn�y#K�<6L=�㊜���u�mV��]�=NN��i1�(H�Q��dx��pu܎�xkW��o���V�d�_j�+�4!�z�_d�|ׂ��E�x��٬z��V�j���U�x�X���5�Ѝ6�t	�ՊÚ�cuq=��_��0!^v�U�����c>�y!�-<r�}[`��w��T����w��� lל�?0�����bX:^5�:M[D���\puq^�f{1���co�����]،��N�՝��`�)q=(4�Ogv�ū�T*
����ˠo�X�.�����e�K������.@�;�\��A�ao\��=��5k3p4����_>];W�sS2��o��,R�����wd%�Gnʓu%��4r��*��Id�f�<�{�	R2�s�'Q�GD�>�VqI�X�}w�4gS���R����nD-���A7�&XND�������+����79J�RG�E��֧2�t�������'!wxz�x��_}:�����{ ��d���̒�қ�
�;s��Z5���ȷ�s�`x�B��Z66���6�Ü���}��������_�?��߰�*�j��a��V����T�ٻ�;�x5�Ԯ�>�^��f���4�Vޝ�^��g��<�"sf`ff��/�0@�p�������yRY�����+pl���w��1���k��"�w#�),Zr�ʼ�X5���������z��RB�s���WYA�=�,��DH7M���[�7�}} ��G�w[|V7�]�v��ެ�b�_}��.*�v�A��b���][]�e����<�^(��5HS)�P&�)����?L��7�_�f�]�F��^�Eˮ�C���ov[�yE۬�dӮ�wM �ȯ�q>�,D�t�-�,+�'og����+(4�2&ήN��J2V��@&�
��,�t�EU1ݝ��f�v���4uV1`����de��oh�!$��ԯ
xj5�hM����=�ٽn�+� �o�d�CE�65l��aUu!n�;뭔}dz��eX"��˻�Z��H�bFG�`%ۭ[���;�s�5�<{b:�]�v9涷T�z�v�ƍu��m���T�m�t����9նzݦ�6�gp+!�����m��u����	���u���cAųvs����M�6wan�ݶ5�:�<���ۋ��7={un�%���k]1�DMfOl,��.x�F�mv�]�FWs�@�����k;��v�cA˩5Y��q��e���/&���/<�Ljw�w6p�6��6Gz�!��a�㇛������@nh�rЦЗ�(묨����ו��x�ˬ7`�Я5=�5����Z�
��eA0?��� ��n�^�aa]'��)@���	�ݵ΋ڥ.��'ܧ��\����z]��+
�\{���#5}�!���݂��Wu,nzC{t���)[�u�ݞ��h�Ejd�H�M���Ƽ���iIk���z�W�~�($5�P�uwof)~p����Π+&�K�`V)�K�.�d�w42��4�VBgz����T
$q������uv2��#��p�f�Y���i���_�_q�����E���X���U!���v�l���=�ּ�n��xO{�=�)aTۣ�i�Ci	P=
��4�<<j[�Xة��Y�e8/o���[�i�^=A�΂� mdK�׆�)�+zb���3~�O����5
J8_�(�	�n ������݌t�v wa��d���y�,�n�n�
��!66Ɓt�e�bI��x���KU��9���/s�����]�n�¸��IK=b�'�6��k^���oj���\����CA�4�y�B�NJ�������8_�u�'O+w�27�m�(I��]IAb�+�oc7��Px�Vë;$.�C�rL�e0&4�ޭ U��1XQnh����Hڮݘ	�m�����5��T�}�M��]�Z��[�x�Ys�]��p�*i��)�1ZrKAH��vr�s���|��`ݯ�'C�<3�a��y攭�*d��\�O�U�ZKA?kuo2�V��X+�0�qF%$:4�w�<��{Xb�g�'�`ۯ2k�uө�^��t�\U@3�Ûڪ�Я0h��4�;��oC�{���)t��⒫�6L)H����I�8����Ȏ{c�.�|�~�-	��w�!��%��=�~N�zwʴ�F�<x�:d|�pVV�æJ�X�6�`�6��8H1�'�tv�-؋����X������3��\ԏ;iܣE�2G;ږ���\KQ���6��k��fT�U7['��=���u��`�ݞ��D�/��S=極h���{s���S��:�=���x�yY�x�iܰ%9#S�j��ܽ|�Lі4cK��k{D�z���n��k���y�]`���v��] ��<����=�˥��z�eȗ���R8r��m��U�o��Rv��`��jӺ-x3Z{/ڇFn^B"�YG��N5~��m�f�V�LUL�b��%��i��rO�f=Acx�-6����<��\�w���r��֯���\��n��te�ɷ��tlf��T�]��IY	"��D$�)�ϱi���!�ף��e�^�ܻg}�����=xX�[Z�OeפU�5Xh��~��Z�����8�r���%�E;�g��gq�96�A�JJ�AJ�Ө.���{�V��Cc�W��e`��>�2�9�F�Q��o�������ux�<�cos�t��:
�Ik���t�/M%�f���{�G���v�O���Ϲ7W�����g���u�[�B��*Qo[�&L|�ѓ����eVY:��J_?4�xuD�~j��r{�C3jR�ݻ�0r�F��.�����os7Ya!�V�d������t��wٞo�'3�o+�?������'J8�kA�q��s4��w��S�T����O���2=�ۓ����˷/ΞvD�R�,y�R�u��gjF<�\�6�@�A�\�㩺~�'i3���RML=�e)��`}�ۧ�Tn��L�g��S�ʯ����ຳ��Տ�n�xE�;X��]ҮL���ܸ�*�R�+��۬�C��S|�]Z���F8��L���e�Ӣ5|�l����0��4��'i}�h���X�re�%� 6�
gP�pp��*��=�5_s�{9��y�u���Ϋ<n/�=�p�*&���ĮQ�*��Fj^O���e}��w�6x��[t���m��Z�n-���l�stq�N8λn����Ƹͣ��E�"!e	z��e�^�^g(�NV����A��lm�ÖgRy8����޷w~e!�J��bJ8���!�+�XEQ���i2���3mis���������n�Eyz<5ҧ�}4ct�_��c+j�՛��V\��.󩽢��M�I��q�ta �[}�cĴ
"�t��/���*]]��w��6Fx��%fg8�w�~POj�f�=���;׭$u�ӍI	6�V�Sr�O����6�`�,G�SY��Ƽ��*�9쭏��֖&�p�7|��M��&oi���j�2UExN��a�r4M�p^d��f�w,�'�fUAb��ԩ�k�2$��ʖ��X���h�ea�������F��E'�6�tzS}�ΗeL��V����ᒦ-ǉC0w(	�o<z
S{f[ e���v9J2G4g;��뚘����Q�/�l�0=v��5�r&�k�ֻ��5����\�n*�nܡռq�܎��nūZ��֩���v^����l�rj5X��p���{C�a{>-����v��\L�.� ���C2�wh����Q��y���p�v	���
8���tb��Q�:��m&6��8|9�MȪ�h��8��N�q�;n���:��;ldsz��� ��g��Ƽk;q\��r�2G���b#)�={E��<t[�z+G7�y�l�G�#��n��Z}�؝�����r���e�V�%��'PR�Q��ӳ�B�-���K3�%z'v��m	�%��_�$�}4QM�Am;�Q4>����=��7�iq���c�a��|�l��5��T�]���o��;�����"Zek[(�;���j=嫒�Х��)�S�A�XP ���o�ޠ�wuk���}�ےf���}�N?:��P����ޙ���𕊧yһ`�{�YW��u���m��d4�	���Ӿ{�~��ea�]��MO?f��%��{��Z$�yɃ�@��]Bf��j��ɃL�1�����nS�43�Ҏ aE�+�2���3.p�\�3��)8�^�P�z����Z�a4Fm���d����\Z�~��eޫ�-��z�yu���GH;.���q˜��N9\�<bH�ś�ogUI@V�1�q/]gW^;oa]O�����=`2F$�0�w6�n�mZ�l���V�s^ٽ�t�>��vѽ�X���j٦�u�n�����J�� ڷ=)CF.a����Ky�q��]��y��]�mvc}|$7>���=*�W	-cڇ���fR��c��rWÞ���q�?0���QWNIָ9�$S�oM-_4*�^����t��w������t��ߓ��IN)�	^9�7��(k��P)���d�"��� �ژ��a��ʊN<�+�o�[9�:Ǯz��-P�"}u�uO�估�T򪩏rM�1Iq�Gh�������דxl�������7|��0!��L���0#Y�� d|;Oun>ѩ�/�{Q�Q�w��aD�Q���^b�/=��Y�3��d�g/o����|[c7�B�Q���]�p`�r޼�M�m�g�|W~+����j���pZ�Lp�(G%�24W�&źNx5��3�aj�v��v�5�uD)��iH!�����,�� w��!]����DR%���)�ӷ�ƅ���ov��Yo	3+�k\���F��)�6-"UJ���3)���5<@�x��;˼���R/i*�U�{�ۏ���M�O��S�oT��n_T� �a�=��!A ����"nK&��{ܪ�{*R%��ٓ����-��x�b�9�-Q��ˑ^#1{ M��/W����V
#��ڒ��M��MX���K+)��D�5��O�pMs-�oy	��>#�z ��i����C:���@�B �2C�^�T+�m$%q�(c�LKto��f�����@t�m��Z}둫a�#.kM��7!գһ���P���of���Y!����]���x-^�氞.9�{{�g/'�f�=Z�����r�n��)|��ws����Y����=��W$�ن6ى�Ʌ� �|~f��G67�_Q�dK��\�����JGu�"�������E'^9�P�I���_VF�%�����}���ym�;�9�� *V�����et<�ΰ�o.�@�5٥]Џ��)���e�݌���a��80o�=�Q)�Z���	l�p���qΓxJ�ؘ��-䲙�����FS9��_�xk^#vG�k
!;%l���i"�M�fi���7�̰|=�;�۵]��E�3���:W���62���N5d�a���JFL�i%4������l���ي��.�K^�]�H����׌����i�|��������֫��'=Z/f���!�H��Ѝ$��ݛ�� �⣜�tNgffn�v�7�}�VZS���U���޾�jv�������7[��Z{�@�F	�>Ƹ��5��F��c�j�̓��&���^k@���{G8���u>�mi~�D��o��j�6�s�Z)����(غ�g�A7nWk]]���=�o���n��/h�M��A!`� $���G�jH���/VBk$y��w�V�l���Ll�~
�c�	���=�(4��Y�����WVh+���E�a��L�C�bd��"B܇x��I��j^},f3���}������kһ�4�[!%����c)�(.]�^�ȩtK���s�i���]�BL���F<rA�b�~�_]�1߼���{�c��R��݂�VZV+����:�|��bĲﳄ�0n���V8Z�f9hHJN�0[6/�yۭ�x����K�e���}�I]�٦�t��z�G7+%��Y���9��y[�Kn��o�I5��H�L;�E1zh�7'�r�=���gj�B�!�{=���۳�TqJ`�>��g��`�H��)��{�ꮠYZL�XjG��������/�綣f�vB�+%�K�a]��z��~QL�b���t����-���W~Cp{[6 ;x�d��X�|�C���m��X�a!n놓��������4r��M紬�]�e�9R�y��1���	S�ь��W�D�����X����`D�fme�� ��6͎��d}��5�̛��v�ѵ��0���<�ع\G��_g\WJ�Pf�`�q]�G��k��]$wfnwƲ�k��բ�j���ض��E�	��HɃ.`|��飣�b���S?�8��F�&�Z��l���:���8�ݮ�5�ځv�/H֓!�B�]���5������=j*�c��C4;n�H͌V�R���t�(gH�#�<�㹚ن,qn�;0�z��w��"��{�}�[}���er��B��Jݕv�E:�O��ذ騲J���ƭ{6��Fnx�$�*V���n��ᆏ���D7��0Az�q�gD�h+����G6�����u�-R��31mgQg@��{yC5[Ss$�t�>�Y�:ta�$�x��έ����u^�
�坼����ǲ������ЕV�z�z�f��뺜��b���9�@Z˼�:r����>�]���tv�Y,���W�2������b\�K�{��˒�����35��{�G7Kܖ|Z�����$�a��/I���T�֕m��W��VzK��:��0�+�f��eGf�ن�kr@X؏���D7��4#��e⡬��m��=�/��m��^���̌����I>i' �E%�/)���Bn
%�<l�٘��ݻwC勣a�pm���Q����rB4Qڸ���sɏh���nzK+�)���x�n��B��ͯ���+���8�F,o]�˲]Au�m��k,����np���<\�۴b3��koK���^��;OP�xf����s!t�ck�ol��a�����,[�/K���ն4vz6мG7X����4��)�c�H�+g�ٸݹ�@�v9�<��.Qv�w!��pv^��>82�g�4q�멻M����]��ջL�@=�-��k;��#���aӵ������s��}�R.=ۍ���x���9�.w=��0���O�Nۊ�k�ᎎ��SQ�V��68�n�G�v�m�c�^A��m�������Wb�ASm��<��1f9b�m��HG��h��U6*�(��QM
є�R�Ļ
�*�^7k���;v�7����IS�����[qjK�t�mh^���u���p]���]5���=,�x�X��b}�W	��=�vܽ��^����Q�6۱��G�\�m�ZxGp�ugҚ��ݵ�2��3��S��v�'�����q���mI���y�z��c�4�G�V�v7\�<hlr'��s���{�K�Kj�9眶��p�=�v�8A�!��ݗ1�\�l��/9ڴ��8-s�6�oc�rcq��)�n^���v�ޓ����
8݋v;��Br�ڇ��a�����q'ti9���B]�x���n���� Jqq�6���u�^K>����6���p�wur:۶dn����rjk�K�u��V�l;�9z�+�A�i�m����ܗ#ve���@�tW7n�u���m�7�ʯm�7Rᛎ6�9�뭃1�&䫹8ŗl��8�a����jݸx��9�w<�NOk����d�ڂ웮y;�·և�:ݞS�y��\]\��8�l�j��7<� z!V�e۷�"��-�;�wY�Ho*\=�����%x��:�n���yyJ�Y�[���tTGm�k�:��c�Z��q�E���ݺv����_"�� �UQB�⠹2��a
�\K��6:�=4=���[t[�(v�[ǍƸ����m��5i;�%��zp�;�7k��ok���6�퇖�V��祺�mq�+����k�V[vzwmדL�x7�����N9�]�xۭю�Q�U�n��nO>���n4��ut�qԘ��3�{z�eCG���n�9��l'�5uY�z �p�K�p�5P�_�����v���+}j�����S�������q��A�~����:W+M�̓^���1M�����i�?�W��9R�T蠄@�%��	�7�h�7�F�:;V"��]و0�su���ֳ(˗OԜ�v"��������K��=	��D�H8`��4fܟI��m�CܯE�&���lc�.�J��Vf+W=�MPp�շ�S
L����C'g�c�h��7�h��t�26����7ur�H��|��7d�A�`�$����ucؕ���+{2��QX7=����2��w�\�X±�����IsJ	��K���ͦ���&�sr*�<sQ��}��췔���j�����˕�t���+�js�un��e{��䃆5������d�A�YV<A6N���F�vw�Æ��m�6�H�t�y9�0�A��J-��C�=��W,�v�C�ly�{�a+��N�����p�����o�,s�wEʇs�ʘ[yބ��m�,SI�l=�K��˲i���v54^Z�^�Go/oDC,-��d&N�,��֢Ӧ���nu�]��O���ܨ�����{1��ř���gJlV�Av]���/c��������X��+��̎����{�Es�3��*y��c)&ME�wvΤ�q�}r)ۧ\�J�#��R�b�Vg�d���s�s�Zfl�U"]S��.O�.|�i�\d�p&�r]G�n�<����߆�Vg���nʻS���_.F�0b�v�P{��A#h{�т����ǭ-N���/�4��H�\���I4�tq,����}�4�!D��B/+<=��Ei�E<"���M���?Ǟ�X�-ӊ�i���|�{{���.B� ��9U�1���h�[���|ձQ�O"�(�����#�����ۜ\�38������	f1~���<�e�pb���C���w���f�=��p��6�ܞU�G�7r���7��m�`�`n$܏1�d������u���"_^^K�)�H�j�u�������{	����,ﶝј=��FU����n&�'"�c�ɯ���
���~�P�(�ok�^-'|�m{�4�Pi��dn<����X�|�!�TI�۱�t�\f嚜�v��o���,e@�z3uVme�oI��2N�w'<���,���*Z����ŕ�6���_eo�-�bۂ�~���:HC�JL��zk�w�ٸgC��[����G�ֻ�3�A���f�w�N��'�߁t����`�$�d���W���\��w,�$yɂ;7g�:6�_!D&��G��A�
���n�dK� �
]������&�,�$h��&DuIk�<�aι�۵�4
O..�=�mŬ��5�5
a \�����{;U���*��������O۲TW;h�v*G/{C����Uuc�[O�&2��ԏ4_�����ْ݃�V���K��Lw�)�F�\W9v�}��ʚt��d�����I`��:�����%�/�T.�R��6�U�.����S{wʥ���|�(9K�ݬ�Z�7�Ÿ5�I��{j��1�)�]�Z�Q�5c�^�с�.���D��AV��E�-\=����k5����9Qe��|j�OSc,SK�p�
<�Y���x��h�x��]��!l��]x捳|{N]����" �HoQF�v�y�W㛯4�x6��x�N��8�
���b݉C"-�dM*Z&x1L��N�gg5��qa:��4����{�޺�ç֋�զ��C���諉򔲶�*��m�������D�"f&YE"؀̆(�m�#m���;�H;��{uʠ���1�m�^����3A��t�	ߞ�vU���y{���<�꺗�����:�]q��o!!gU;��u�BT�po�����>�v�������/H	�-��J�������Z��+2����jS�B���Z&���m���r�8T����Fa��V�r�u:��n/3�f��x��s���.Lco�C�طU`�|�${�c-
�"�u��Ev� �ER�J���d�n,���N��MOi�_�7^��{x�"�)����Lv����!����&_/S��ٗ���U��`���
	>� �v<N��G|�o -W����6׶���꙾ڛD}�W�1� ���Щޝ/Ęl��.��yhR�T��m=����g.+R�U�f�	�3lVy۷�7����c�|�ZC�c�b��Tx*|��r�$�Y[��W���6�s��s�y��·�v�r�-��cz��ΦnkSێ����c�ymhn������ќ�����QǱ��,'m;�\��h��u��`�[v�{��v�8��M�pn�����fk��wZ�ۍ��nG�n�/CHi�F���0�}(���t��&�FA��\���w /[�Kg]�\uv�h�=z:�R h�'�����l''���\4�Pwmf��<i��<,���6��f�P�m���<]����?oZMm���vh��'�}�i���������3�yh��w�u����f�
m_K�-�-?o=���wW
h�+!�|(�
e�`6	��n�Kr��l��l��T��L�,�YG�d�Is��<3�/+b�����r%�+2�>�Eji��$���WYS�!{��qK�綅��7|r�=qUh˕�-q����8�F�����	���RáGP-0���)�E�k���w�-gw�3�ߟ�j��c�-$}�^)�xӓi��`�ݽ��,�j_O*B�֎U�4c���9��A��5�V��{���*����uն�,����Z)@C�Z����j��x�2�m)x=��5~��1Xgƅ���ZYz���`��6'��kə:Sw���qk���{�we�e���<"�K�X�����`��qaɨ��z!��;�vg%�>.Wshk͹�۴|z&�(Zܱ�lzUo��ψg�����k�����b��{�w$T�7������D���6`��u�������D�n$�l�����W��!۠V�[c�$]���w+��$ E(����]�^���,׷ؕ	Ӯ��ʣD���]y�d�m���q�v�*h��
�TJ�Ym�}mB����`��VM�&�OU�+w�CG/[���Z�Y��W���b����qOy���q#�9D�//z������9�r��,������������6��9��k�ވ ﺜ~l�U�|IJ�ޱvH4�	�i4�fe�?E��t��ի�Ƙ�-�t��[��2c���c<�}DJ~�KtSɻ��B����'�,:���G7��Zo��e��%ݙ�l�騶md3��܆�\�nݍ�[c��Rx3u֝��J�ʳ��#�����WDddvf2m�k����zo�Q����H��^�}�腋���V�B�a~�2�v�m����<����S�.�vx��V���#�Wsx�]zl�L�`B��]���/i��9ק�����6j�P�J�vb�ĒM���"���vڇ���LSp'Q��u�ͪr�VQ��I'���i�z�N�L��V����n���X7t%��S �r�F[��"���������]�ݢ�H��g�R.O����0����J�5�^���	�	�K�!HF���l�{�UЕ�	�7��l�Gv��_���I7j��D[�bW���jֆ �-�p�٪G*Il/� \8�T0nhcmf��{�11�CR-�:R�۹f<)w�U���1�t[o����
�KѹE�Ւ/�"�W���o�7k�m<q>S����n�w\���v�6�/&�W�&!�$M$�L0g�)"eI!�ޣ:�̋���.T[���0�O����Xl�|.ߊZ�ҽ�{�OW.ƪYˊ{\x���F*�*	a���C�Ç6�L�Mx�������^0�i�O5�[�T���������	yi[����w���a�ˌ��&9Y�Sa�/��ĩ��XӐA˺tCO����u�V<��#������U��q3�޳|�� A�(��,��r��3�ʑSx[2�U��c�iZ����cI�5X�ߍF�fΠM�Rw���x�>�P�^*O~3���%��kwB���uLm��Q�݅��ѭE�#Q�
T6Tx��=w��������Bi�Y-���3x���Y�����e>�?]�vQ�A��s���c�����>���w��:����ߣ��qĖm0{��k�ͷ-G�ze��� �p�����<���\$YB@��14l���x�2�뵝ohs�rt[k�{��֬�{zd�
lj>���}yY�@�3cs����'Q7���y�q�[�o�����d��-�2���]o܁46(��8L�F���	���P�I}���;bo�.RkT�}ew�b�cv*+��&q�KժPx!�J�6Rn��6ټ%�b�0vv�sA�GP���h	t��׆�K�
S�kC��p{��n��8q!Sld[D����!���'&s���	ۣ��N�-͂��0�Kn��7�N��q�x߷��Tj\��zB��h�w]����q�p�u�{H��.�T�LOe��fe�e�J۷����֐v�������6 ��[^}�u'[�p{3Ce�5�u�<jIJ��}�RM&+ze��΋����Ss,E���F;��D.u���X)e��{��(��M��I���r�k�R��eUڷ�?�N�ސ���k0E84S��5��:ۏY�l�m����V�v��5Q�V��1�.�P�/`����עo����y��������g�ڼ�nͽ��F;ut�=�Ev8�	�r��g�¢㮮�6n.y:�����������M��[l�[�:�m�`���Z��S�[��uŻs��=>p��n�v{���s�n��Z�͞�Y��	�hvx��g�3S�;x������;������=�r��c3m]��$*:q�yE��8�N=K;g������j�k�f�
5�ችܢ�=M깊��p)�K��Qi����G��by]��o~�Ь��ەo=\�n��=���W����Rw���F��P����]l�>���=�C��뭟
]�K䊿���5-���y}���[��C�����׾�8�Z2ܷ�xGQs��r�B��4F�D�F�"	2)%f4Ǽ�nm�>`�A�}�=)qcnrȌJ�݉�G��㊰W��5��s��M��q�}Nn�Ab��P�%H2�%]^c��^�y���7%�]�1��2��jss�V&[��u3��m��<n���D�A��T�%.po'Nق�=ck�Y�xq��\]�7�F������@�N0Z��ܑ��j�X
�]|���e#�[�N>��S�+*��>���`�w�i�|W:��)<�q�p����`�!JH�ͩ�x�^��k�J^�=����f��B�29��'wt��S\����w)������V��!Ь��Mi�� ˥f�o�W��^
��	�Ks����e��g���z�9�D�*{jʙ�ߴoLq�g�����j��BсB���i��N�cۺ���8M�<k}.E�L� D;��m����X5�/ʶ��̋�A[�V�%x��)��H2;�����}F��j*Ol�p�z�S	-�ҝc�SO���B�	^��=oyD��^*W`P�|�o�]���ߋ2D�'$���ӧ��)���I�%�;;��:iZ���r�uo�6�.���()��ݔ��R��γ�	"E��F$���G�u౹'j�Vl���ڸ��zy����Ml��rUvO
��DWU�!����_-��6o|�OKl{D,�+'����Ǎs�G�Qc���SF
�I,a�F�.�������/�U�lM�c��ݞ���'��C�1]�Σ��y���#��7�Q�᭗�}�������\/+E��W��U�H">��v���C�i��}�sepm��dDL��bf�Z�j3�h���~[[��:s-J�1v�QF��;��:��]�͙�Mtج� r!z��vQ*�*ɋjk�k�u�Y[�7�<��'�{�wV(��Pǖ�$��wswf|�|�ݿ�;��/3oJ����Pv��V��['j±e�R8���M��z�T۬q�Im���O��˖��X��ő\�AZ����u��n)�a˯]�	=�b`�����JP�2�:'J��M:�^aѐ�ӑvH����Z�7U�xTĹi%�S��;(��$Yj��w+�(^(q�m,�����i�b�oq;&,l�IT���t�R8����[���ۓ�%)��52`�V/`)f�0��k�t�7���l�̭���-^^�Yn��¹��[d�Ny���oip�37�=���h��}��>����Nl����8�ׇ3w.���kD=��=/�on�vKn�^ņ����2�ް�g,��'Ge3��"�8^A�RB�M���'\v�-��7X~��v�@�wU��n�W^��	�Fh-�F��nLF��ݛ���J�`�����̫���XV�Q6��YYƙ�K�����J;{;hmsW�-]!;!C��oe5�l��<6�+z7�)�L��&�}qoAXz�Y2�Ŗ�r1�k9��M�2�*`�K����=�V�]��n�z�[Ȓ�V\;���N�2������4���V�Lk��m_c1/�ozI��Dc�仡��- �W�2��/�]�&MD��Ca#��b0�Ḑ���AGÙF T��S�zO9pt�'�MCf��ݱ�99����xk�=��=�{q��Wff:�SbG�������vQ�Q(.<�L:�ʒ5VRSV]m���K��ە�(��!��GAczul��x�oOTd�2����ܦ|%�x���VlK�IJG3��.;p��Kz��� �g�r)�[�y�&w��]�t�mn7O-G������Vo����x\�Z���׷�9����u-O\�l��?VZL�/NF�[(X)(�i�$�F�t������K�x���Y�N`�9~+��A&�R?o�<ѩ*Z�׽��z��<�����A��"�R��zo<�;ױ�U�2�������oϲ����C�Ԫ�;�޼s����g!��w=�4�S-	M�q���Q�B�;�}�rm�[f��D�o����G�$/k���}�tN�()�{-��nU��7��ka��Uu����;w�p�o>b��g�㎶�x����jW�nh����PD߬��ؘ��|�e�Y�a9E���߫��5�Do��"�7�ْ�D���\n�g��⚯`Fc�b�r�g�GR�n���.��]�ru�x�,�.6�Ҋ�=1m�j�3
籓q拃���!qEƻh����|��_;՜�b.긯�n4���z;D�����Z�Iz��h˽���vo�&�`E�HFJ7x@3���m��w�t*��ʻ�;�k�YD�!wk->c��Ҋ�s8��e��7�<5vUM2Cn�Ҏ<��� ,�ҦRE5I&�b�zoL����9_����%����J�;mE�w��Ug���`��y�|���+�w��5Q0%"ѧ.K�z���&o}��%�m�w�r���a�56u�o>�h����}�{�+��!��{� ~��¾d�
)��;�Ru)bw��7�ǞBd0v�{���B�.�L��1tW���)s�'j2���ŷ|]D��P$m��*�j�졕��8Ҹ��d��H��t�jte�wj�-��1�E�-Ƕkw"M�Ku����}5��kbt`�$�go�Y�Y�︸㓋��?rZ���u��nCv����aw���6�×��
��{.���u�e���sy):�۶n7&��O�s��y4�ʯGm����ko�.ꍎ��ܝ@f�����A[.�h`u�':�9{v��[T�����a���Ƴ�zC�ex�k��YL�5`n��uٞ:�ݺ�d1ݢ�r4����t���۶y6�w7b��Z�>%;ED>}h���9�Z�"U�N��J>kv��+rۭz���Dvѷ��v�����ɾ�nM]�
ez�I=2w��$����VO~��Y�z����N�/˃���!1!M���wfݐ�<N��.����x!3�^
jg���rֵ+=��[����q%;��C�*����gAO���D�(Rl_}�Ѧ1o8�a��O8�������nh<��3��-�3'Z��G�uU��\�lQ�e�񁖠M�T
)wlJe�U��SC���}�m?"�r��F�ۮ�d�>�M�#��m�_?����*�LB�9S�Fu�g�d�~���|�;���1������@���v�n����E%O�t�1�;�b��y�¾!���xy2r�U��Ǫ"��DB���/���t�/���Zar���6N;��x��\+l:_�	��,5�3x������a��)1r���"ǥ;�B�m��]�ػ;�����C���*����6�� �e31�=Roft����w7���a�����)JK,���yNa�ǵ��'au�9�\�Q܊��Z��Pp����̅�ޒ�����bX]�y�E	�{���_��l�Ż���6����R>�E��^T�y�b�������e�,���e�$I�Q!6�g�srT�~�v�ٝ"�h��\����q\wG��ӦE�4,J�/-��M��wN����p�G��a��@��I'wo%�[��v�s�n�&$���}��{3,�<I9��6f�]��=]�����z����b�o���� �ch�aRH���]�r�CS��N���������k�+B�KP��Z�L7u����#�:g�{|��H�XH���X����l��s�)ãO�{<�g�{:�Lt��!6;8:�V��j���;�j�`�|��rN�$��]�!Zѭ����i�}��]��P��>�m���p:Ȝl�i��i���D��i��jI�ݝ��u��s�#�p�ɤ��kP��'�R�=h��)�2��e�����/3
���|16(�|A2I{��]�����#��Q�_�+�s��ͯ)7�<�"]��N�.:/��L��:�����%(nQ�V�.0Cp���9N�2�ܝdL����n�b� �[����[�X
�vm�(޲�֜�_��&M��G$��E_{RB��2D����ڷ�(m;��̛��=#��
{�/�q��x�
Y���~h)CԓhR�� :�ק�"�K|��HT�Ɛ��d��2�ٓ��y@��2�)��x'4OR�x�n�,�M�o��x�x�����Ry���؂���E��#l��ޱ7�qc�%��M�\��;bz��]sѠ�OM�|�{�u�i��Q�B��o���������{�����G���}-u�i�@�����O��Y���}��V��]�d�w+�퓓J�^�`�ل�W�^\�bfbm��FG�]��yV���׸�KĻ�$"g�|D� �b��[g=��v,�^��wll�ɒ[{=���������#:��_�?+ы9����q�n�ϱ���*��(`&t�D2�gH�{�v;�O-#�>�p��-��/>h���>��͋6�㍛���T<�����d4���~���K��F���f+�N�s=V�9f�q��˗lub���u�ӹQ�	v��rZ|ං�Ѭ�>YN�#�f�ll�J�Z�W|��
�I�*ŧ3���x�|���+�7�[�� nV,8������սsU^i~����.���yk��7���ek��S�K��%V����&e
b�eQwRQvU�<��{S���1[�h�� Mq�Hɣ'g��ɹ��(6�aSɀ�c����iѓ|��xӚ��vj���
j�Jxb#ƸG#IhB��-��h82��ǆSM�׫%�ͽ�ʩ�,����s���h�K9�ɐ�d�U���~(Ӿ�h�'�B�RD�PDJ��W<c��v�_LG�}m4��E�<p�R��H�#���޶T���HL�xR���1&�X���$�-Р[Vw���M�߼Oݯ�9{�3Z���"�y��y�Sx��g6��P�-���vlj:�y�7Ig�����<�Ӎ̈���}�9�L�Lǟ2�C��z���]3�����^��mO�D�{k����� ei��&A+D�ч>c;g'K�	�hӮ��we�"�.j����҃���+Y�$"cV��y+$u��ٻav8-r��G���6��Z�wb�mu�.Ď�u���n}���?'�p�y���v���̔��y{J�x��R��Ʃ��e�Ȩ�8��L&�%�1r6Q5A��q���u׍�Gu�n�F��tn��w^5u8�I��ݢӴq�yr<��#خY;1�r���.nwm8��;px�:ݨ^e�����ч�n��xp[wjܽ�+�$P�v����7'��%��D�F�=k[!�Lg��>�WXy� �I��	#�~��+xn�=���s�~��1���%yϥ�}+��vnq;�E����o�'~�3�H,0�*$��Ymw�9b���zW%����5̄�Ɔ�]FK�٥=�cj�Ezm��}��B��I|W��nG�n`8�\�7�ef!��f�s/��;~]�qg+ɣ7_z�Ǜ4_v���i91/4�ҧ��4�w���G�[ 
D�%�.H��o{��R]��z�z��*�b[��*R�!��|���F��C61%�*��X��=#�<�l�!&Zd��Y>X���6�d�v�w���i<5vCE�A�zr��2��k���;��n��OR��ֱ��*��55�\d����v���6qAT������u�p]ц�
�pP��Ah2KLw��'�x!��3�{[7S��\����u���?wm�����x�\f�\��G˽	�/�Є����TnE+�=L�y��і]�s���*�E޹�k��R�8���bV�{�.��Ek��4�UשK�S�Q���.'
r�K:YBlC3�v	t����\�]֨%|�ߓ��b��������D�����<8`�T�t��a�Y�'J򶷻�a�(��/��C�,:�=.�=��>��:(M�F�v6�ÎV�����mܸ� �*��i��/E����͹�,d��w�n�[��DSܖj�t��y��vny�]N����kfs,�%S���mؖ�;\|��v�c@	o���4�]��� �w�*j��(n�Mi�:�9��Z�<���|���rQ(��O��	�<�櫲�&yZ���Z�P��q�Y�`������@�������@7Nw[�x�c>��I��%�YC�m(�Ny�/��e�\�o�Ͷ���2c|�asXv`
8�E�nE�����:�=��!�ʈ'��HR3�z�|����S�y.�"�Y���;�ws%iU���f�B����N0��d n����;��>�.��>Еl� w���w����s�lYyu�qX�y�����M(�;n�w8'wK�0�ݦ�y���,������6c=o�:����aů3l�ϛ�F�3ݳ��΀��U��陥S���n�1���`l�!0Dm,��zA��H��8���k���$t�؝"�e��;���²{��6FKK�7��ی�-� ���hl���K_�\��k=;.�".�#ٺ�}nN��7���`u�r�B��	�z�����ef�jBZGg̻;5�t.�*����lv��ۓk� ����5;����8-a�q��]������ͳ�}k,]�*ox������\�opv��<����;6�Ǽ@N�9:ǻ�g=}|bJ�lϑ�9e�I��y�]��n�Y�Q����ǧ�e{Ģ�yzW��-W��l��U���8{t�a�܂�xX��#fHTMHo2(�F+��7�`��#�ܠS��~Z2^�YB��:�g�����n��ۇr�(d���p6F����SUeB]LH*�0�'Yq�0[d,C7��aƲ�wuВ�Y��~�h���^?D�����)�m�S*�tjs[�f�Tٌ�<�w=&�qMۯ
��N��e,O�N�t�rv�]KG�@�ݹO����9ld��k5����Y�%w�O����t�h�v�0��@�l%"V-��_Z����7ٜ�QK'v��U������0|�%1�����{c1(e睨ikr2�� HL�H"Qr:ZN�\Y<!n�X5WG3ǈ��y�W�;����3#,��E7�6%�ݙgf+Zm4�����_MĎ����4�^j�f�����u�X4;���[0�*�P�;��|�6�Ǭ��N�C������s8���C�o��
W��[[�.��{H����Yϊ28L���^g�%���(ڢw��K��w(N2��˘�ѓ~�ٌr�v�3;�I[���nR�%���H�A7i3Չ�m��CF�޽�R��Ϋ�R��\p��vGw�|	�����ܢ:�X�e�W��f�f��8
򎞎/D �fCI�0c؟<�;��Sg����Ot���	өf������&S�b�L\[�mϾٷn�b@с�l��TV=�r�n�-Ǖb���2��6�fvDn�JQ���w6��(�;˄`P�ʥh
�m%�T
!OR�o���M�w#�����'�VU��)@&a���V��6�=R
�b�ҝ�]+��]��7zo� ��R�b+�dki�{n�H�5�.$5�^D��L�W��^�z~���<7���$��b746��ڐ��^5�Y#w��l>��+��EU�����jG2�L�ǲEۍ�5�b�Q�K�V�Ǜ��@-��J����.���K�Z���T��Y08#�ә�o�L5��n��I�z����������Ι�?��^�6��Q�cKT�7r�*�	��nVH�).�]���ض%W.���*��0+����ć���� ��ӗ���d���lkI�;�:�>�\�D0!��d+���m(h���5#K��s}�gT�.�n�l��C_=+p�
�63�^wm7V6v�u�䫶v�Wۻs����[}x��E���
ؕ���K��P�p��n��Fg:k��=���y�>Ğ�m��0�{XU.5���J��m�JƜtSQүl�F�ܤVn�
��%��ۘ��y�r��ٵ��1�O��/�3j��!k�qj�,nk
�����f�ꂺλ�ĺ��C(�����s���Ò�דn���p�nos<�^ھ75+�|D�ɡ��\ӴN�^�M�Bk;{��D��'�^�k���z���<F�P�u<��BM�}�Iם�N�Y6�։ύ��61KQ�eK7���V�u�@pa-_���`���R^��7|�?[߿���ny�Kv�pW=�'I�pc���'�ݻ=���;�z��k?q�t�9ڷZ��^3嗍���jG/��'"��wVV�˙��h���8�q<B۶�k�gXu���kl��zo4오ƺkgX9�2�4g��r��n�p�`,�n���[�i���T{7nrW�x���]�7�qh�ugt�q=�I���x�ͅ.��-��<�>���ݻL�͌��sW`�\����m�9뱙����v���۸��=�v���v�m�9�=���[���Ӱ��R���1�{�����I(4[wggm>e�ǐ�m�c�3�9�����7#�r��`��f�z��Xv��Wg���=��9�;����
`�����'��ovi�9��8�V�w=��W#ru�;��v^�6���v9c�뎪w�}/�A���-���51ѝPAV��}U��.�������8�/��Ƨ���ج��$F�<k�������J۷mv8���B�=�����βr��z7	��c���s����^�;�<�κ�S֒�%=���fD����g��Z<��KE���Cd'�Vy
�X���by�t�H�ۜ㣎�u��k�=`8��&�s���96��u�����r�<Oa��t��0=�<n�p&C:\\��t��Zέ��\�gڰdPe��;d���í��Kq;d��v��tƗ�v��@�NL��ۮv�ڵ'[��V���;�n.�m���tK5�hֺ'��a�A;=��^��]�t�l^yݹ;\GKt�m�S���g�1�;��]Q*���.{XY��ue��MF����.-�]�;h<�}+�m�s�˸�AjpZ����omq�)';�b�+���l��C�8��XǏl��&�f�˸��Ѳ��*��(��/Q�v�8��B��b�0�MO9��sFz{;��]�Ma��7@lvǶ�r����z�yz��i�/B���N�cl��yY�è{���d����4-�3��Z펆�H��{�
��F	�c�{gK��5�z���^]��v��fv�9�ɽvrv����F���gZ�y�Ɠ	VA�p�] �WN��cq�FN��p����ֻLu�6�nP���rv�{<�{=h�x������q�EY�rd�`�yW�m�#�v�iy:-Ns�8��u�����x�vYr�M��8�&�8[����n.����#��a���t�i۫�j7`9���m��ź�����bH�m�/E�l펡��{��=P!kZ�-���?E��/�N��j-U'fR��!����|<���5(�����`�^RﬠߞG���1�*&�R~m��W�:ê��ge�b{j��69���[q%���P7��7G�![��ǧ��k;�3�a�����cHAI��*��C�'��}Y
J���}
��r�y�x3E��"乶m<���/����&κj��*�"HI�8l{�8�R��Mxs��/Z��6��kw]�7q��Q��.o�K����m����d2N9[˓g�C;zY�W��h2��������60:e����*b}[M�H��=��Y�e��}^ݚ��-jwqSHn�>�y���＊%�e�t\��th���h�E�۵Sv�m�Y��9��p�a�A(#P%!H�$��_C]�Q�y��'��[�A���-wX�5��+�sH��I�ۻϗ�1[���H�LO�s��Uy����핖�b����j�N]ɺW��5sw�Y_�����:�����>gu�V�J_n�X�K�;-��5:��Qd��������5
�^۸�0����k!�:tY}~�N.M��2/7Ǽ�Y�Iצe�Z�nV�Ʉ���.Ym9
Yަo�-[v[���{_C�h����|Kݒ0����d|�ǽ2����_=��P$�!��rW/U�HTݻ�B	Βi�����D�,+��?{�I"/_y��~�j͋�kg��B����!.-��H*�L���U�OD6�V|�zI�Gq?
7�"]��ӽNp�5=İ�έ8<�Sc�A+�,/�;^ڼ5�Ц��O��)�i�<�r�p�z�����y,����;�8�cZ�����o��pĊ���3��-��V\��'��m�y��Y�I���-����m�����EJ\dx{�Q�2������b�gU/U��Q�}��mL�e�MN�\~��Ec=E��enP6���P����vwG�l��c%RN���)�L��ST�� \d�Z����;.5P��h������T�e����\� ���r����"�,�.�E�c�r
�k�wOT@�',d���f�Y;���1A���-�ѯg�����Gxl�����5z�0����	��LRh�S%4;�Y[��^�����y���K�'+\�u��M�E�r�;�e���;�.I������Ԟ[���-$/K�1���e]%��J[���ƽ��XN�i7|��Ő&Оق�mw��A$\�ۻ��܊�oB�����������I�r��q���g��rg\���ݯN2��dܠ��l��h�Тlw�V_Kלv˔��m�[�sB��0���7z���H�A&���/�q�K	ꐌ)2���*��L[�{�t����-%�LFb=^G�]�$�l%��LŘ�Bȗ^�W��;h`�FKM��FHrر�S�ȡ[��~
��q���m�F����ͻ�^�e1��f�;���ON��6���B�Ǻ��)	1$�pm������p�~�}��9�m�¦�m�9��Y3n���&S4e�{�f��R�5��c]�|ץo���V���n�Tz��h[o���e�a��3� ��n��"�sg���%E��G��t���\˗@k���m������-��ىp�ǟtܼ�ol]i�_iHg��wtRCf�/Fe
C�Խ=���#K7���ZrX�yn�8f�kG�ܝOfQFEF��K$i[X��nk��B���ǧ�D�tn=e!ݞ�n�:A�KM�h/Jf�oo���	_E�����͝,mZGl�Ci5�-;KQ���c{3Kb�(�0�m��wT�9����i,�/�AA`gnf�Y��t֏��i?)��)��w�IQ}(w�������.4c%5#17^��A[�|��P���Z|}�r�w����}j�]��{��ř3{�V7k����C@�<���	3~5�����p#�f���͠��m�i�2R���N�v~�����]�%��淋rC����0T��xm�n�:!I��I5l��'t�Py�z�[]�9��$�؇���Y1j�yZ�ۨ��)Y��TB⻉W���e� 3յ#}�r��J���+Q��vԋ��.�륫Y(`멦#�:R��x]J��ܹC���m
���6���[�վV7��$�^cN�D4���t6�n�$.mUɈ0-����]�9��v���8w�V�>F���W۝�
��k�O��q�#,[,jy�Վ9-kwn��Ym�����s͉���˽�d9��ڝ�y�W���n6݌sā��滗�c$�܀�X�ɹ<q�K�2[%�`vn�vݹ'	`z3��Bj6�>�� ��m�<�[��}Gk1���n�,�X箬����<�ݳv�] ��dp���Ϋ��d��T*�!�D�&�p$�Ӄ�o)P�kk�~�763=�%���\br��A�}�8����h�_T�3�Y:�D��]��G'}���� S!��銱$�(�_	W]����[Y�=/�*�7��n��l~6��M9�\��%Z�IԱ;s�� Ri��)P@�`}��F���v��;l�5ގ���<I�돕{�?4��<	��+VJ�I�pv�eܱ��
�6ԅ��H��˛�L)G�.9�P�HUȭ�TX�}�ܠ��n����ԫ]��G�I,�x���$�$"(&K	��Y��ѳ�`)uAT��9��w�K�{:V	��������������,������󨻄ߑ�� �I�ȍ%"Da�vnx�f賺�`��;�ԩ�m�v�g)����k���(���ewg��t��k����� �u}�ެ�E��
�~�����YS�v�����J��L2��i4M�@�{���n`���k�5��� �X�:��ϞN7���[O+��̺��u��Θ���Ad�(k;j�,f��е�^��~��qf�1Mf��ۼ�`����f�ja���3��b&3\<	��po�z'}�ظ�:���}��&���c���Bܝ�=$�����t�DpK嬬��ޯ���%f�3$�_��{u��A쏅�����j"L�ƢaB#p�ͫ/pd�\�t���cmzQ�ܮ�8�l×���YМ;��^�O�5����8�蹝ueE�tCȄ\�B�(G$����$q��*V����]I���gyb/% 6�����eOe�>�7�v��W��� ~�cΜ}c��,���۴��]�O���v�<ٻӡ�p^��x�8�����d`�	Q��Aej}��ݝ)�aH-m,u����ˊ��y]hʴQ�(�r�d��R�����CB7����[�
�TG�э�����΍zX��M�qzonAp�<�Ϋ����v��=%%�(�^fTq6z���9x}~�,�%f!"9�
�����^�8�p)�Q�jx�-\����-,�u�h(�9�&Q�˻�n�P�i�]wz��źD�̻-�D`�m���bM4�
�j�~2M�Xˢ�ns����P���-J���oc�޾�<	��T�d�|n��=HZD�x����.=s�>4�50�ڎ2�銉ũ�h������+��۔]`��P���cqعy|�]�u\���z�%��;�I`��E�>ŕ�4���y/r���&,�kr��~�\u���;�$�*^¯]c>s�G]Pt�E������|�]=�v�i�\�t�v�<�A���Z�B�r$�#nN���{���MbҡN%gIj�I<}�9ej��:�Ƕ=뻗)��n��Ng�;g$��_+)Z5	��
�2�ef-J���^;'��:w��|'�p�Y��9ow��a�Sp�S�7�7��ީ�L�8ȧkpgy����%�Bԓ��l��&�����V�mR�tZ�L#�� ���V�����O�ĳY�^�ҋh�)�6��۴/&#Z�;��n���Wg��.Y��O!-wml3k
�:��ٺ�t7���ڼ4 �o1fV;�g1�&f��Q��L�L��J����t慗5�#.�b��]5������{D��[هN��6`�e�2W��ڕ��쭬�tX�$�E_����]��Ks��r{+�ʹ�j��/�u���V�5�9�W35��l�/I~�y\DQO�$��<��:�����;�G`�J&	Gvֺ^i=��8��rdR)�T���[��:Z���Q�m|"�2�_�i�/��n�(��u`��`[���엫���2��pm�$�4\"�w��#7�9^��~��(��x�bC�y�=��Z�1'+�&dps���Y}����:w3V����K`������n8���/&��+3�v�eyص���P�iw�)	n�^�:Wt���s�S��%=��uВ,9���7M#$Y��R���g��dC��J;7g����S���m{1�	k�ہ���\����'ǌ�"�� �}���'t��r&2E7�9��9���S1�g�T��x�����U�ؗ��TO�/U�8*�'�;z��t��o]z�����[���8�$����b���n�2�Ǭ�Y&��`;f��t�Pt���)��q��g�w|�M��)�j�bYe��X�r��'�ޫ&6���S���:suf���s<���T���Y��g�ͤ�wMq0�#mˇ������F~~V��H���]%�W:�:q�È�#�ۣv5Ҥ��k)y��s�v}n�FuGF�9�m�mTl����Ϟ�-ѝ���z)�x�Z��:ݮ���v
9�x��gy'\��gm)����Ns�y�����y�s�� 6�^��ֻG8l�h��>��Xi��)�� ��!�v�ܭ�+3v��ҧ�$�7�~��ԛ�0�n����һUȦ�|�E�[�<�UYB�ѱ|�㻧�K��籑�.�^���2BD�� ��|ȫ��=��+JWשּQ�]�Pwx�xù��ҧ(啻��?6���L�/�sn`�0�=�܁4R�(�h�p-WlR�Ӽg�^�O�U�ދ$�GEItw0o����?a�D�R v2W�+���ˑ�,CK�X��i�<���o�/|�
4�V��1����Pe.��hn�,<�L�}�YJ
�v�\���e�E+o2rβ<�q�8���`�&z�����<g=ڼ��X�9F�f5���ӆM������7�1即'o}�=��IR�����0լ��v��v�MG<���>:�-��Żd���J�hb�e�4U�v)E8��_{�ro�52����D�SUv;�uǢ��3C6���n.��ܞ%S�z�ٛƙ��WAa�*))&I��^��ǽ�δ�{�J��΀]�C��EO*�Viq�L�W���9]r�=�r���k��6�;.���E�Ȗ�}�S?1�y������uwT=�o�^�*"ů���o�Z>��Z�<sv�q'�������8�NiX�hM3�"�D�L��d�2����x3�����(��"+'��M�X�S�\���u�7����E7Gg��V����Fq�m��J�i�M��F�I�4E�;�=���ԋ�g/��Fb���1��jzCf����M�=�rRr�M�8ϳ���h��t�i�Kn��(�$�'oܨx".y��+[�iN�Zw��@{w�ͥc��n�8�h�
�v�ʼ���^�V7�IN�u���8��^���ٝ=&�bڮ$�'��8�uc��ݮǝ���4aa�2�S����ߟ����w�UϷ��N��vv �>X�0Ÿ���
�s�F���O���>𡱝����+�4_�P�$��dR���F�v�V|^��<JXc��k]`A*��]��3�N���S�1>�y*u�I�Ԋ�Tq�8Sڔ� M4*��������v8�I��+��I��-�RҲi���N3�.�:����6@�s�m�"�����=b1,��W���vw�Y��ii<�v�Պ�e�Q�͐%����R���ե�[���ۦ-�lj�6|p��׷nJ���+@W�E�^Z��Z��3Q:���@e\vxg9��l���/����
sv�s����;jܣ��W!�����U���Yhk;3�`ڠ���Q2�j�`8��j��وS��x�P6^J�d h�P;w�P�fZ�pT���w��7�P��
Q�v�e���IV? �h��5]�?M0��c�F���c�wP�gzgT��rL�Ҹ�v�{�#�D���G
�mcs7E����=O��4�e���z���R��Ɛr��� (5(��1e�(��,��x;Un(���Xȕ�fos�ʼ�m��T-�03��gD�k��W/���wϦ�Eo}�����CjȵG�*�f�NE4s��5&i�;=o*3������JFҧ1׍��씝j5����]�wN$-۵�������1�Z�5R9�3���[��Z�y�+L?Ji���f^�KEl��,X.��\+����ì����*�����$������c�a��oc�\�CM�����|v�t=��jLW_���k&������N��Q�۞[M���=�HI��#wJ՗��黺�t�Q�Y�&�t�E������®�z���ޕ�7�f3��L�v
ݧp�(ݣ9��nq8�SɦB��jT�m[�s\8fU��^�\�QNW掅I��:�܇����	e��"ӆ�s=u�����*f����K��v�M�Uy�C�L�VI��V�e�)x�C7H,>��p$�)��[�5�4`%�=g�3>;ל]�X&�U��GGZ̠����7F����ׂ��|��FMw>͂�^=O�p|laQ|���}^��'	e�E����Bfb�[dM^3b�nԼz�
���l%�#��־Y�#�����	,��}R�}�xӅ���Ƨ��|~�`�b�~������W���:��K��u�����e�[]m�sm�妵�Tܸٹ� �n�r���j�{���ku
Wf���Z3I!�/�_�Å�������:=B��r�3'�U����ߙ?��y�`ϭ�	O\�wH���ƙnI,��JI{�6W��˖E���b�#�=�}�1�/~�(�����-��ʘ�����`���ܷf��{�c��Nf�gzJ]��@e��@K��L�4ӆ�j<N�DN-{�\6F`P�L.a?(�"����`B-δ�ίen���Cy���<>���px�H�{2U�	�g������" �y���>�Pk�3~E��`�.�W�q=�Km��|�޵X�]\Nl�]�U���x�.�u����-96���[tPO/�a_�aU��i�����7S��+�����H[��*`3��wN�:�@M����W�s}�Q��7Zf{���تw���}]�7���^8Ǐn���j�uJ+���x)����{���U�h���^�㎕��z��o��M�ff`���2~�~�X�*����]Ӥ�ۯ��s�����KSk�3č�p�p�C�xh��k������GT�R��s�h�g�wF1�L�~S;����+�k���hlV�J�:[�M�*r'u��Uz���Z�ƀ�ݪ�ў����ɐ�)�nO}��_�"��b
]�+��U��W�k~��}T��ˡ�q�V�A���1��{�h��Q>�M�j�_ߪͥ*i�g7����o����~������W�ߴq-)_v���O�}��F�,�F��}����R�X�˛e�H��!���YѠ����c�^�Uq����{�~��]Ԥ'���+�\#U��ϳj}���x1���:�׬����8�b�^����}���l�WP���}�w��ǭ���·�y|��cW��S��� ��O��T���1�o�i��0(�1Ũq�z�׷T�w\�,bi]?��齠8���O�:�u��4!vu�G��n��W�:��>�iv�����6���/��z��e��Q��{T��tm�CArD�v` m~�ECgl'�AN�v���fU�Q��ڽ�������s2U�:1���*�1�y�������S;T���{�}�ٳ�:��1<�ꍢ�<����t��}Aʚ?V:{t(������f��>W��wX~���+�ߗ�ɿ�Eh��Q�����v���?U���+����~?^���mR�UQ�]c�faΡƓ9��v�M�ݺCv�����Ϙ��%�U*�~��2~Oݮ�G�5�}�7��|�������V����V觉S*�wQu����6q_Q^O&:}wsn�E�S�n�No���l~�E�a�� �0T�j{¿@ ��A�'Oۖ6Asg�>@��/�#%�
x+g���GI��N����ϳ%�j��9Vf�T�X�=9SS�
o�`^K^߰�Xy6�XG��n���z��k������<Pg	��e�Sg=]�u���wz7��=m�l<�W��b�b����s����ln����}�;���.�w�Y�Gi�*�:�`pg�Sn�`�=ς4�W���b�;t&��շ^��8���U�;V���ݨ;���MY�c�lvtG=$d��e�I9^���v��e�y�nk�0�l�����&�lcˮ�1���$]�Z�g�;X�v���Z�f���1(����i���N7��M%3;���4�\Jf?6�7���tq��F<������n�Q2�+iZ�1�ݳ��ҿ�n�|���_���:��*@
��DV4�ګ���W��ޚ>�������>?P8B+�0ia���;��s��$�UYy�6�z�^QU]mMr�iƉ�o~��χ��4;��i�E%��I��V*�s��ͫ�T1�U8�W�}�΃C���\Tr�Uu��+(�,T���~W�WႿy_���i���o��,�xz"u|��j��dJ.�����	֓����JM����i_��������%�O~��?n��Y��X���=������^�������oٳi��fy)Sn���kl?~�ϝq��)��~t���{j�V�8�~�,�1���Q��G��|���B����}�T8PQ��W9��+�Mg�ٴr�C��\�'[M����z@�\@4���D�l�!b��o�پ�����[����J��E�����_._�z�h��Яw��8~�? ��G�t�k�G������JF"�(\��v��g�v�o�+���*#�+�;��Sf۰��G�K��v}��AH+_B7���	��ڟqiQ�P��ѡ�(��ٵ��G~�l�{����gޏ�~a�|���Q���W���S���֍��RcJ�>�X��:��>��1��~�t�?���H:Uz��mYn47v5kvV8b5WM��r/3��zNǞ'����yM�����V�oN��}�?v�>�j���x�D�)��s�8�u�և%�J���o�Z�W����ƃo���iW�q�T�R��_��;�~2� m�7\��� �@R-Rp���CЯ���>�����Z��n1_>s����x9WM�f�uxn|�{V+�C`��Us��dʂ�������W
����$A�лU�sUn�p�di�Vq�O�zX>����
7��z�k׹XvR�����JR�ķBYWI귔s}p[�I�|G���-���W>U�O�ێ���}e��j�<}_�3��yj��2����?{Z�uv���S�X�t#_��*�)�E;���:v��c����(N(a�	z��l�"a�#'E�R�2�m�YT�������z��i����|� �_����?;Xa"�B�=<������ (��\~�����ƽE1֯\_�wu��ٔU���U�i}�3{%?bd]�daVY��k�0�N7N8la�P��,� Y��w��11@AV�M�|U��*��A�Y6�m�i�R���S�V�ܕ�>�_��f�#$|���X�37ٮ�}�/ª�� �:zV���J��ǻ�� ��s[U��ҫ,�]�=uU�z����8`�a����]�raI��ө��~{�ߵ~7v��yE3]�2i�FM��r����%�ײ�SZ��f�Eй��f�Ư���-]<�,M3��5R����V��eUB����˜������}W��_�kj~N\�UT����OA
Y�Un�ʫn\p��=8Gc\>V�N鵺=s�y�`Ս�f~DW�<�8��R;�v�iJ�+_�z�ƶ�U��U��R�{Vq���^�O&�U]��!<���������=�?^T�O��(+��iLt�M��Go=}4m�i\ޯ�ӷ�w�q���_�.U�Vՙyu�F�!�d���<*�31����Y�?�(�߆�3՚	_��+�ʈ�]�x��E+օ������9څ��b��e�����q���8�y��]�[�=�)���?�q�O�`�\=��;�%���U�R��x��Q�s�ѵ̦�
���+��ҽ��E0��!{��w߽������'��G�|���n��B�����ؾJ��4ѳH/�+���0^�P�ҲJrR�t�-+GL�!ZEvix�h&Vi�Z<��.Ue"�׼�{����ʦ�����S�Ǌ˩��D���9���؀4���������L�VQ�2�Q�L_߯����cwx�i�����j>r�4������ܸ%9��u{�?4ν���4�Y#�?Z���$�G�P��wL���5����� �7�,V��ݠ�TW��f�~�_X�D �;�NX�T7�ml˩���m8��oMٴ�n/3��^�T�^S��w���u����a�k��i��~u�|��Nٴ��SZ�i����/���g�U��]�4�y�Y~��eB���z�:��ۏ[�T���S�z��&���5�Q�OɎ"���Jf{nz�����v����R�A�S�s�d�X�s;��4�g��b��1�Y|�Ɨs�7������5�]�8t�z��SfT��tW�����X�
B�0$ ��[��s��ۧʚ~�<Ӷ~���3y�F�~y���>��S	���6����7�Ւ׈�����!�D,P�0�#��?}��P
iKfX���[�ga�ç�6@�7��J��1����r�~��Y���A���P��;jX� {��8�����E?n����w9�޿'�?}X�~k�����o<��������\��b{[O}�������s�a�^��Rd��q_~_[Z@@���=K�=vxw��~x�y.��3�n��A�W[�~�,_�B��/�S��׸#M>�]m=u�������~76�uL7������'Q}������u���7��3Y��Ϊ�r�G�j�[2̱�/1���YE	����&�楺B����~�éG+�Q����Y�)n��z��	�Y��O��5K��r�H�xRc�ji�|T����?@�t`�Fz�mM�ذI�o�ͼ0=�"�e��2�\����ej��D�@�k',�"���[��XW�I�W���������k4U`���U~h"Ȓ06�8���Q���E<���=����k���c�+�Յ��{�}Z(G|�x)\:�E'S�}�B��{��Ï>�N�g�B�PwP`���+����wG�S)�C�M:���/U;��Op�ZUw�������?���vVQL99�6B��hup�
�W��ӑg>�f�v���q�3�"V�l��~O?��16��\��S>��k���ܮ�)ga�0AX)<LS1R`����4UnMdA��¬�ŏ��7f�i_��x��߫�~�S����.���;�o�M��:��\+�/hi�g�)4Λ��^�;N�D������z;�=�t~�<OE_�|,��X��叽��,�����_��T���}�^!��+��ߙ��{��SU!U4��'�~�)��x��}[c^y����� Q�"G���m����V49xji���<�6�6�߷�
O�|<�~�jz��Jt��z����5���u�LLy�_<���6#�OȆT�#��:�4|~`�/:K3۫gޭ���uޚ;�O�M2����F����"��j"�A���#H� ��1�e��.��(�"�<~ض�w���<����k_R-��/�gս�{tm�M!���V�韻������[��c"ϐ�c��o��9��_��*�zp%��G[C�r�~�q����ܾ^]�Y�d�_Ȍ?f�}m��$
"�������t����t?�We�Zٚ��+r���8����W8b��O�������oW�!z�C3��o�5�|��|[�N��U�|:W�P���fto���ǁ��u�*�l�qe7���lM\6ܬ�f�@�K�0{�SɁe�&^�2j�g������X�ݕs�ڼ��lynn���z}�d!I|X����g�Ƿn$ʁ��b�5��7h��;��9wo۞Ȗ%�:�ɱo)�mu��#��[q�����z�� I��}�l�U3���x#���m���x��	>����>��m��b�T������!�z�����4�u�@j���Zx^�l�]��ݱ��=v���y�sn�!tt�	�=���vλO�v����SrgT���8�ɓC�Z���g/S��8�N���n�Ǘd��*)GO6i����ן��y���4��9�5��5�p��U��i<�O��w���GS��Ic�!�QYQa~���7�5���7W^��S�oWT����p}OS��W���h 
j�9Fj�矸���[1n�n�0�!��{U���O#�����k�y;Y��������Ӭ)�~���u��q�T)�Kahc���ע���ڔ�?2�کו�����*��U!���gJ�㿑����ʬ�?na�?8˟@�E��Ր7Wو[)1�1)*�+���l�o���6���w�R_��_�Z������93�~���Oz����O�7�:�h���v�M3F���_�p!�Xk@q�J��g�A#k��yt?#$M�����Ev@�{�ij���r���U�����������h����T��\C�>��٣�ݰ��6�9_!�����o5C�9�;�c��X��^�?W%�eފk����M���2�X��e��z6hV��MeV^V�N�J��|�?��Ti�@^������ZV+� Ek_�V�]Q�<����_m�c+�Ry�����4�X[��xAv��g�V����c���?��h#��w��=�i���!O,�:�V��,�F�.���X9��g�OB\���v7NwS�q�r-�::��sk����1�9z���g�Wݬ޿|k�l�T1�q�j�O��%�o�{�{f�����aih����<N/z��y�&��
�y볈�i����t��5ڔ�V�eO�lRމ��{3��g��1[r��:Υ�������������<����eH_�lV���rF@�J����;�uB����ѷ/;Y�ߍi34��߫���5�w�:R�tT�c�����mm��C�pb���
"��R�@~��g;4�����
����l-�q~�������UwI�RY�V}U���۩��K\�;O�O����AteEN8!q���#��m�3��k��������~���M0u����W�����p�c��������s�{��"~ki�y/�����H�4�1��H�+-/��h��i�-��Q��~�~�6,I	�F�	�w���Mj�l9���~�evf-��'��f>����G�r?�iG��]M��k��������o���Z�� B� 3�`c�Ó�wޣ����_u6�4Ŷ)i���?}���(�+1Q����ÁO���[���>_��Co��LU�)
�(UA�<������߻�s�P�<�a����¯��B+'�i�}f��7P�s�y�w�򧟐�eNU�杻�3־�,���3(���S@v�r]m�\�/k<w0g��n:�8W�YCh�.@bq$��x
���г�G��Ì5��{5�L^Q�4�ىo�w�}�5���c�y6�ܺ�>��Ѡ���w�Ǔ����;�����/[5��<m�x��v�(�4�����\�L-�Wt�fV���c=��e}⍦�l�욫ᕌm��y�'��"75��� �����75u5�a��>�~٨m�<��CL�c�/�����S��I������>w���j�
���u캪��i̻�ͅ?�]K�\x�nж��߳f�3ݢ�R�a�Uf��/{5��sZO��y��hC-�euuC�a9pg[K�����wU��E�^G�^ݨ:�RJ6���'��C�E�b�1�(-��mu��d�!����1Z>�<�Հc��=G��8��{<ý�?s6S���ha�V�i�:�64���ә�6�w���� ҿ���T��a"���>�r�v�4[�Yo��d15����tٶ|W��m:��l���9F���߯��{_���Dӄ@A����O��;��hC�wU�~�C/�_��o�i�����ݷ����,[��Ì⶛f:m��O����ơ�YwP�*�����N���EZ�Ҳ���3��WY�wTm�<g�S����l>�|�o|���6�]ϿV��z��|�ʴ-���Q�j�'���B��4��-�#�=�w��y��;z�P8��ݻl����!kM�R�HcJ���毻P6�K��tϜu��f�1�u3���N}��������V�dU���g��!�B�y_�W��\���sho
��g�*�A�97E C0� J_OS��Nĭ�jK�
�2ګ��۶<��'���j�K��M��SΥ��߿]�IvU�]�wG̴�����jZgݹ�������i6�&}�����Χ7S�������{��s�{���K���\�:�f?'���ު��啗wYyx�8��&0��u1�~�/�߷Z)8�k�\f���<��?Uvc��v��6E�V�/��_=��؅�y����f�����!�7��(��Uߎ��쥼ʬh9p����;v�v7�]W�fȄy=˾���Z��am�i�1�s�}z<���y��|�f'��8h3+�jz�,|C���ݺ��s�)t�J�������أ�m�A]��	�	��[���#���#�0�2���y�XZ�&L.=��q�&f�t��0~���9�#����X�fm�V�o�q?'�UHbRv�����KMr��\a�9p������os����<���[}��̝tj�\U{c5LU+x�Ӳ���d]��a����􁬳s����(�i��&E��2-�4./e�����W+���b甖R=A����ݱ�̮�Y۝����R�}��N2ߩÜ*��c�{Q��\1���@�����`l��#�]']�?^!~[�!��}��C���u��n�;�^셶b)��NP��3�~HR�Լvrx>�E׵�r�'�l9���{P��T߹�:�S]N�<�_
����1�X�tETz�}M�&����C�{��q��BV�{:�<�6BaLm��J��]՘㗅�^:1�O���cA�}�7�G��sڳ�0�|�~2���/�"�O�i�3��L��s�%�6@���@dVz��=&�T�XU��c)��o��mU�V	W0�RGCO�~�(��@0�u|�G,�Y�a4�V��/p�W5옛O7¡���9�����l���i1����z��A���5HUz�h�z�k�OA���)��ϝ��3}yg�����Z�8�0�w���cT~��Y��uvW�iکo��+(-�BU�M����gݽ�ʆ�R�b[{�`.�D�P/Y�w0�^���U�XRJ�c&��3U�$�!$�ܒH��IO�IJ�IO�$�$��H��I$I?ԒH���H��I$I?�I$I?�$�!$�I$I*I$I7	$�	'�$�$��H��I BI�I$�	'�$�$�ԒH�rI$I?�b��L��x�W.w�� � ���y�A߾��]�Ȋ���B���	IH�J�*R�$� �%EAI*�����D� ��$UAB���m�
R� )@O|T  4�E
��AJ�� HUUI%J�!JD��RR�EUQ	UUB��(�%JRBR@J���(0��    -�p>@�sqX.�nح���n��:ԕ��(�.�]+YK�mV�n�n��FK�v�&���.��k����6Λ��
%A/ ���j��E��ὀ     @   /\�   �G�ս�:�εe�9�׻�5z̖��{�ieu����vk��mo;v�ܕ��u\Kǀ;{�kfEz�g'z�q��;ey뮰η*���:w3[UY�s��j���U�uڒl��bǕ)J��     磩�ke�!�oOOy�s��n�󺶶*D��M��ۭ6���{֨\��*�����i�J��V��˭d���n[�@�E�����]��ps"AKl��R@(8  �Jԉv.�:-�]P� n��Z����tGc]jT�]�N�.�pɣ5��U[d�3��:::�vn�A�U�n��HD�8     7d�gUÎ\��h�&�]�'Mٝ��.�9�:��Ka�Qmݩ�T.m����l��
� a˶w`�c�T��I:����  y���ƁN���2�f��@kE��8\�A���{bfhc�ݵv��h����
6ó��l�Թd�;i"D����ITI�    = /1�l��pj�ّ:�l�뫰�.ƨR��(J��WgsJmErţv+m�e֐4�V��+�]\
t�p�
E%UN   �Sf�+��X�4���[t�p\-�6Ң��:tt:�2t�Y��-�Gu����us:�hN!��IG+E$�R*��   �th6������3�KX�7t�s���p��;�H-�[m+��+��P\�t(����8uҋ�eu
T�R�  4���,ڝKa���tn�m���j���4����ԁ� ��N�v�RB�4�κ:��{d+]�� >�E?LT�*�4d� C &�S������ M `� $�3Ji�j��Č��#L��<�ت�D� F�2hi�M2h5S� IT� 2     $�$	UL@h ��@���w��]�ݼ]�S���2��Z�Sv���>=�zI���6��q�����/�����	$����8VpEvļUEJ"
��4�*�@���}�)�Ad�$�TDU�c�Ev��P��a'���HLA`k%IP*
J�&�VM@*Md��J�Y+@�+!P�@��$�K@T
�DP� Ą
��� �T�
���b�� ������ 	XBV�$C	*"�H��I&$%@�J��eL@��T��YYX!�
�@�RJ��
�d��c	%ea���0�!�P�J�VT���a*V@�?���C!8���Ԓ�a,�@�2���!��Hk*5�LI��c*LIR�Xd)�:O�������p̾�.����ّ����\������7�?a�WM���3�2�/�÷���Rv�3���1��;�񞻔k���b.�T{'M�7�b���=GLS����f�����Nܧ�a�ٙk���,��tfT*�j:��;��861Ca?�Q��]f��P��3i,f�Ti��TG/cqm
���`+����8p�`�����Aܾ �?����Βt5�f���V��R]YF�|�{cu��8v;!���8���DKC:�~�q$������Vs��}�o��|�hz���n>i�<nq3/��U�)6��rV��K���G��R�Ь�����s6������i�:�9[4Y�Ws�+��{����dv16%���RC�`[���I`��}��v��du.���)�*�;�{PfK�Xգ��ۓ���_��Cv�E�9�����4�v�Qv���/����y�`2�����l:�T_��;��$�5��;9f��l��ŕ�[��!�v���\�2�\ޥ«iF}��K������1Du��i�y=B���BDtP�QU������e��vA�
�w�A4po���F-�R��`���#���Z�Nǲ`�W�W��n@�!C\YI	(�X��v,+�I���!�*�1�v��8�U�2;���TN`v�"B��\Z�� +�Y�@%KSj��Ak]kVT��47@c4���Bi���ŊM@=[���5��0�Wd��]�%���sdf�:����Y��̿����̿�U�Z0�Mkɗ����q�����]8�mK#O(V�UU��X��{*���r��X����)��stV�Ժ���N=wb����[J!wu�X���i��:ɶ�N�
ݺ9�+]��&=嚀1��������"�9p�@��M,�v��:o3)P#
W,[��'N[)��Mp"��rQ��%g7Q9��(��q`��ӕen^�@@� �ԖB�4~
�m<*�شi@�fG��f���ݍ���@�:#Ս7��HL�tX�M�a�C݂*°".����p�şb2�uS�vF!�}�̤(mֲ�����Pׇ,;)@�I�鸭�:���V�R�+eD�7v`�nĺ�3dE5r@���eF�q���;���M�͕+n�M(�ǵ
��i�PkێC�
��T�e�κݐ���F���W#Wa�(m*zfط�ۓF���qf�{�1��͒�b�8X�*�W����ݕ�SwEb$%�mE���K��d�:n��'���dGN^]��Z"�%�a��e�XFVV%����r���Yrj����fV�$A0^ѥ��{`Ԣbx��H'&���y��Z�j���ϟwe�P��Ȭ5Q����"�1�z�[k$H�1=2�oD���B`h���E�ܵ���G Q-�f�;����iQ��ģ0��B�۫���q�!Zs�n���9F�������\�1��+*�6bDh���]7eM�ǹ��4[�!`��6�X�M5��
�kZl�I^ٶ�[^�2.O��kjCr]\]j�:N�td����Q���)o"�e"�RK��}��J�,���6�ѥj��ې�td�!���4��x��H[UdU(0B��9Gd�1-�PE�$4�j���+Z7����bf�Ml�ek;	��V�d�ʇaڂ���'a�[���f�DMe�3jU�{F1Or�gN��C g>/�ӏ����m�mS|#ռ�8FE4�F�ӪCV]�q�aӻ����T��M¦b�v�iJv���uu���؛�Ʀ�wzjЪ,X ����&�J)�n�f��]�j��r�L=܊�9a0m�>��
���ՙ���m�J�3�T;2H2�ֽ��/Cߍ�:��҅l���wi"7]1Ͼ��hV�CXTv�jX��G�m�A'tu�ߐ�\#��(v�J�VcAś�.��O�~�.CdU��w��W�z,�!7v&��}(]���W���c�:��_`���V�������UNk9���H�C]�;`�Ռm񝛠����I���bh'\,;qh�0I���+*^��VI�.�N59��$���JK�ڼ"�:.e�b��)�l�z*
�t��B����R��`
�m���V���k�Lv����%3a[�>��m�7ǫ;$�aݐj�wM�Юe��ՙ��j�un�1�-5)`�)��[��q�����4�Mr�}�5"7.�N֊Hel�^bY�[��E��5�H�
5c�]�3s;/�.\�֣{2Z�mhRS������R�6PMf^*�S�R��'(��"��N�n�ځ{����#������*]��{"W�2�b��c�k�m��C�^[�r�R����;�����P�O(�8�[4w����HF�B��r���DXFa�滕3r�F�9�n�'�s�'�tH�BN����+��e��?]%-wvC-�6����A|v]Z���qo�5�WV�a�\+_�!bd��B��݊p�D�Z�B���ˍ�l�B�wP]0�HD�8���m �`�+#�S:�@��o�{��f6����U��1�̓t+�2�u������(֭hma�Tr�����;y&��{�h6j�F��;6�y�o��ddC\�jݘeL9.��ЌwG$kDXM��R2\�{�љ�M�{��&KU�6�&�hŖ��+	Kիí"�[��P�4�R�l*�p��"dh��*�\�Sj3D���IM��� Y�]��k��W8�L�&ӻ���GX�wBI*�r�7`ҏ�wu���*�����J�MN���'u�"�A�����B�:yg�U�i�׵Y���n�9{�S�pdBL4\��T��M��Pmh�9��:C�kr���,Ҧ0�U"�V\��d"VF��r��9�/dl�7iM[6a�]�Vc*�a:���C�����V�T�P�KW�Z�::ˋ�.j8ͪ��7�	Nm=�1^F0SZ�D�g`������os,ꤩ��	0�f��q�^�.���8�1��k5ʪ��Eȡ���	����[��w6���	�H�O���a�a�ݬNL�ѠP632����W�
��9qU鼖�f�́(����,�(�Ypu�\{��F�KuJ�UL8(�u��7P�OA��O6�D��r�4�^i̵�orj����,�,V��J�.�ŭ̠v�hCfs7v�(��;�|��c�E����9�Fa�|]��k�w�%�ަ���A;��<���4\��f�7�wJ���-iۧ2F���U�44��8K)fn1����M��.�U𠢷�V���r��c�`�0���͹�6ޡ���YVZ�
ݐk��1gV�!�n���ݸ'��㫺v�G��
�Q*Ѷ(�^��
���Hx�׻�2��fǌR�ƵʨE�qIy+�gD!���ٚ������w4����B��B�=��*JQGն���(��c����)z��y�V�]u�b��Ã�4G��S�b�f��&bU����-r7;�*�Wtn����L�jئ��	3�^�ce����*f,ɛY�2e̗w�;]mG��lҡW.P=ōz[V��U��ۥp�G^�ٓ.��0��I��o`�ON�k�s�%��0����hF�vv�˪��Z��Pi�0�@����tY�
�8�;1�O�jb�pp�j�%�r'��va�#=̕[��L���X�z�ο�}�9�D��p�JИ�ڔ��UƐ��� ݵ�'jVh2豭���n�n!k�\����ꆖ�s�XUcD�wx���0� �!�5 CP!��P �CY q��!P!�P!�:@��P!�*5@�@��C�}<��7��;X�f�Es���j@�T�mt��ƏkW�д�F�}V�!���wn���U�A��v6�k4���{�	˲^��>};Z�	��j�X�٘՛�wЮ�˺T���b�!٨��]����mftI:XN�ʡg_+���D�b��;��R��4��>�����D� �����W��I�SBc��cݓ�fي���K�����	���]]�V���1�dWIە����M�s!ͪv��S�U��ػV/5���2���{�\�nATh��I�{�t�[��u**���7vʕI��s5���ܣz�LFN�x��[/Zε6坎f�Y	�{����UOg��1�u�P�8�������a]G������s1[��6\w�ch�gH�'^�ޕ.]e0��x�k
8
���O�<`w ��]^�X6��GF*�~0fn�:Q����b��![�0��{�b�&�sqe~FS2��f���م�l�6ىA��u��^�D��*Х�C��쪥�+�cj�����r:oR�[�kvc�s*/��]�!9u[@�3$����0Y�M�
�M���`�v�`a���n8��B��utn��BQ��gvqˎ��t$���*;V��ZdU�k�}h�Q���P�j� -ހ�G�:hy2
�Ր�rn�*�Ќӹ�e�6mX��&�F2�J�P6s?���o^[5���GNʼ[�,R�Lel���H����#{�n�	H��Č*�C�1^e��{J��B���:�T��������Y��
Uv�S�QM���fl5�k��F1�n�հ�6�=Vi���kwJ@��������w3H�e��z~Ƶt`2��Kjm)ή�ؤ��a�{zn��

��$�Ţ�%�rĪGmV���Si����d���J8,���0�ѥ�ڽ�	9G巺�)=LGn�+�Y32�S�j��h��V#�7��m���ü�]IQh
�e�iI�n!����,�s��4����3w��i�0�mf"ݭ��!`�y{N���4�$��<�$hS��n'�@iy�Ef q��,����ʵZ���T&�����z��
��ͻ�K5ё(�n��&B�q�UmB�8Y7��p!GB�d��5a�ͥB��31�t�^��ڔ6��N�Ѧ2�������L���{e��M�ĻV�I��'��e��]츷�y��Sry/E�c����%ǹE7��Kv1�����2hjz�;�
;i|�w6g�Mӛ�;a:ɒ�kp\F2�X�F��P Ek��h)��ۻwi;��mE�P2�|@�XКj+��]��]��9c$-u�l46���f�[�*X7h�f�BS���-h�_�����#���s�y@Κ��&k9��ͼ���T����M�E^EJ�X'�F���X�:�:Yj6�@",�
H�x��[!�+ot�Ղ�R�ܺͱ#�2��������/f�L��8�=T!j�]O3.m<s��oY�y�2z����'�R�����m�>�q���ݻ�x��/3y{������I�1�Sp�9J��I*Y�^h�*c�W�d�1*�_��~X�w��"�0�Lͽ���2�ڷ=�}K�Vb��&�����b�cE*6K�3ZݽTxAzԪ��{Z��T�a�l�D�o\�6��jJ;��Wx]�������V����RR�me�ɔH� �kgi�&+f觟��M�i�5�w��W׻��f�L�V(^m:�O;ԃ����mEw�$H.��ԥ�I�.�B���LV��9�����'�\N���Ń32Y�SRc���ɴ&��F�8j�I8R&��gE2
�ȵ����L���2��2�,�t4�f�dU�%��@ԦA�a�re-�ɳ1�t�V�ܺ���V�M����wt��N��&òSȃ�.ؒm	0]U�RY&U�� �G��X��ƨ�"˰DܙGYOJ+q]:N^'g7pf��́7kFW�"���f�E�v���M��d�K����kO-����]bC��.L��	S�}h���
�_Q���$��p���R7�K]d*AJޮ��r�ftqfp���O�[�V�cA��8�v[�hܲ%&��}��O�s�U��Be���qwlG�e8_n⵲ڒu���T����:�^�jNA�j)��</.�ΙΧK�X�<Sm��(dŲ�Hhm�1��ǡ�Fۦ�¥8�r�z�L��ɂ� {���!�i�����C�l�&)��I�&�  t��=�%�s��UVݛ��|�n�.?}��h������Ky.�Ϭ����M�YW���f����e�9m�>���m���[t�gbܥuw��Y���#FswՏjٕہ�$�T)G&e%��n�*�t���$˰z�U���6EoN��Xթ�q�8��n�!��lꬨ�I;�9կ8�9�	ݹ[7�ZH���Z�n������+\��{�H���pl����2�l�)Q�,Pv;^��<7�-괻�K�u7�zFu1φ��Et��>V�,��꼝�V��43'-9t�+q�HѻV����͓����ޫYDE�$��;�ȷ��"��ݜ8��B�:rȊ�	�JG[��\���;jG�}h��Վt�J����%�ŗ����E��xv�7N�d���S˩�K�ЪvX@١xfsq�un���Kiwy��f4�{��	����P��G(�O3���^V�ZW���L�RR�T��[UU�i_�������E*Ԫ@*�US��0 W*�T������>8>|�vq+���@]�e1��
)Wh�>>S5*�ASwT7Q*�PW�A�u�jz�vt_����:�^��C�,RM)$�$R�6܊B������WeV��>��ҭ��Br����6�s�қm�2Ȣ����>|��UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU~����ʪ���������������������������������������������kT�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU_�U|������������������ϟ>|��������������������������������������������������������������������������������������������m��m��m��m��32�ݽ��WUUUU0RW]UEЙ���� *��⍪������W�����������Ʈvj�j������S�UUmUU*�j��V�g���+*��1+�U$�-���I$������U�Mo���털��1��fu^U��0v&tؠ�Ŋ��S7j1,���f������v/�6�^U��Pd����oGM�ԣ�wz�ڔ�왑i�%���M+��ڇud� &�V��D��g���TN��KCTy|,Ѥ\�a�}[�hJ�uy�r4���GL�{Y�����[j�+�g)���:���!���8R;VFg#��M�5�Z�.-]ī��0r���̜����zR{{Ыx��yc������zjrB[�c�G�e\����0�V���G4Q��n�lCC�!�ћW��j�4hHC��3l� C���̲.V���KM���R�\bb�2���ٴ��lv:�֨�:V�Π�s&9MR���	l����wi�vnJv󵹋��hf-�3�Ή��Pj�։�3TR�W����Za��G��e)�^b��ۇ�Y&�誃U ��N�~�����[O7)�)�k6u�X��ҷ���`��f��O�����lZ��/6��9�n8�_k�����oo�������dȰ�Zk��w����<��.r�\�A�*��33�n���b1k{���B�୤�S��C�������ּ;2��f��ӷ��(]���,�ޓU��LC��)�d�~{�m�]�;��8����͌_}nh; �9�"~��I�4pum�+�c�oVq�ݔ$�vB$RF��tŻo�ұΠ�&�2���d5 *X�͋��Uԝ�[�2%Ǖ�}h�shm���҂;`�R��$���OWN�[��k�}E0�c�a	+���A|y���݇�^f���Nc��S%�E���ՒվQ���U�p���N)I�o�ms��v�J�
���I�Ӹ��jgIX�ְ�K��2��P�}Ф�=���%d��glbLي���gr��XS�w"N���+K\^�V���B��x7�g��o�l=dW�:���slX��Ek�������3���̈5V�g�������,r��˲��ha�+�:}CL镅�����wT���ګ��Sl��ީ^W�L��h�ɖ$R��rܽ`�i7U�6�JN�'���H;�3��AZ�ֈ�[u�S��fb�Ij���A�7�SN�-��&sx�C>H�Փ}�S`Vk�M4�T6�fKMm"���QޥH�on_
�l��	"=#G5��� ���������� �9v<��W�r�4�t�C�	q5b����7Zۭ͜�AZ�ǃ�S����x��������X�j�fq' �uEmk�LjtҢ��9���ˇ>���z�ݱS�s#g@�fĺ�O�;Υ�sWR�;�K�Su����1Vh�D:�NJfbV�c��Z�����ӝ��d�[c�N�}����orVasb#fԱ�-��P�5�R%os�����g���NK�C}λw�Hg�v�J�6%oR�Qs�x�*�ˣ���}H��u��v�m�/Z��:,62=!�ѭn_=Zj���m�[��
Z�cfS3����h��C!�x�Y�i�frYvcM����&{1#e���^�+���4~廳�;0�l'�i��H�pM�U�̝fc�jpʃ��qPUR+�TYSq�r�b���crvᜑ�����t�p��M�je,�p#�Y�s�S�����[8K"�XF<Ǻ�:u�Yߠ2-�c�>��maǪ��!O�ÃU��K�nm-{�~ۺ�E�{����=&���E��9-<�,Tb���JN|h9����+�}f�m��1�[�N��foXa��NuY$���BpBbcɩ�u �+��⫵�"�\�-�Wu�5�RH�5>�2^�eJ���î�[*�UX�o�������C��Ћy��J]��2��QZH�P*2X�j���W���qQ���S��A$�s���0�4�gI}|�6���眆ʹ��+��j8�u5YOI4��ֺ������u]�!۸�θ�GF�-���`i��A�]��L7�D՘�漤)'����y���зƓXWYWn:%�`´N���EZ�8�kwe��S�KX*�:�Ru��% �N)��r.�i�f�y��$��0)]�X¤'_Bɂ<�' ��-n�h��u�:�-����̾ǀ%�8q/+�{8+��\%�+�S�!"Q�ν��kh�ţ;�n۝s��
�boR����U[�Џ�׈6�%�'E BuN�)`W��f�X���:�鱺�7+;%Z��i�uM�
�6T��:�or��'uW�/�Q�=���d��Vm�3��`�}�(�����lݬ}�j������Ǜq��[+�2�L/�px��oC���D3o6�v�.E��47�/y�X���gS������ _-��_.��l]�ĬV �U �kґ�'�{�:��<���f�����b̗cO��tA�
�ΙJ��x�Jg-h���*�&e��|Z�[���8aW�Œĝ7)�V�H�"�yQ��v!zoPQ�sCNі�7pl�y�6��qL|F�x+]���gUDkZ�%J���ɾ*��]�%���LwZO=@N��uj�����[�.��アs�6N�,�OZ�g�$���/�7�]{�/Y����3N��v��������p2�2X�T���
5��syM�ͩ�0>ʼ�7�f&9oj<�M�J��πn �o(���}l��CY�*���G��[�c�(R�&��X��Jk��G�3QW���Q�T`��0��z�'(+�r���n%a���+X{]')��]b6V������=�nD�]�*
� ���I�]#�Z�޻x�f�u37S�s�&(�M���L��Yg���FkT	���'���3O+ړ2��q­�����)�J�Q�U�*-����e2��ݼB8�y����#XK���� �^A�&FD�qʴ;�)��Y���܏L��Yk�d#z�����L=z2alE�Rba3�)���;�>�Vwf�[Ud)��c]2s$Ƙ$�r��������1�E�܅�mӥ�<��,�(0����"MB-�Ig�fQ�	j�Y��<�H&��ݶ*�d�Q49Zdr��9�� ��kxj���|�c?!S���w�S�DJ��r�
YM���5��霮�0�Ɠ�v��x靾���-��w� DXB/� ��x��f"/r>N�ֻ�Gq�ԅ�vL'U�%���9�#o�x��IUużŒU���܏�K�Egb�D��)X�LT�O�O�ZԨ�l���U��a@Ge�;j�\e�In+j�Tp��e��ķ�ٔ��ª������
�X���:n�M�!���C��W+2�����*�{y����Uz���1h*�8.�;l�[`S 4�0b�:�m0�C�9LwV��=!0e�� l���5�[J����R�&�Xi�x�m"�J��(�tp�BH����oH�*�*o�iN:X$H��U&�Yv<ۗ��l�ɲ،"D�Hő�h����(_I�k�Ɓ�Mu�Us�𵥜�X�s� ��q�s�+.��\˩����:�3t�IR�����v��ƞ�A[��=��/�����י��pй��A��ًZ�X'����v\���SpA\b��%@mi�-6wE��ZU�4P�	i�2��_�WM�nzQ�i$��XdU��=o��\����I�-Gu�NɵiU�VU�a)uN�؂��7�3)]��*��O
unskgA�d76�r���\L��)mfRb�l�@���CI�S�ҿ�R�5�P����]B���� �D_a��Re��+�Y�E�!�NJ0�����k�Ѕ&gM�5�eK��#y1�I{q��ұT��%Au(���%V��1��51�WZ(
K ��U�eA���^�����a@]#��y2k�.�8�6��V"��!�"��U]�x���	Ү��}o��-?*r7!��RmR�uך>��,[EUY��٭����P�ݡz�dJ��ws��޻]��`6v����<WmH��ܶ�P(�����8��eG:���z�^f���0�4)4��� ��6������kGt7|�	��kl�z�e�C�j$��pd<˭B�UHWgVJYF�hD2��ŷ]�Cm ~R�X��Fʗz�L�Ǫ'��m;f�e�`eQq��B�_]��Q��6%�wM����e���d��G�e+̊-u@�Q��Sw̭��trV:����Pt!%���)���:��xI�)�V�El�zC74ͫ��yb7#4�J�{�r��f�Œ]��'�����m6&mT����G	\Qw��^��Tr�fQd��	��F�+d9�I�,���|e_Gt����s�7@� xn�̙7;�^�397��d�snjP@�1+4\r��U��Qj<a'T%J�����@�6��x�&�L�A���00������^���Q�[�I@dL�Z��hmZ,e��N�A�`�V�$�kg2�����l%Aj�3�C��,�gv���vYi��1�69i2�U�]�h�{���|��C��������9AÍ�z�h��f�U�p��tT���lQ�f�
��WR~+��;4��9%�b��Uy���ͬ1��AItΝ�yڰ24J�.��Q|Bm�#�_gW���0S
tզ���Y�l۞"#��D�]��Ǫ� OE�\O�C6ew�5��k�h�Q�~�-�6x����:̓�H�w�s+�K0��4���>ċ6nc�]#Ŝ�GL�q����gh�ǻu�ث�c�ՖZ���Hea�ɟ�T"�rƢ�wT���V	�06�so�61��85T��+��c�.�ir4a��r�B�!�bAk��j��<Nb���J%"V�ȚSFZ��Ӆ[-3��s���o5���؛��7X��Y���H�˫�.`D<�ݒ�ԔFd��e��n�E`K쾜F��2q�&���_|�H���.
�޷i�n�A��iS�ģ�y�L���ۦ3l`���3I�� a�n�!Vd�T��#���2L�^�g+r�ϕ��n$P�ג��2TM �E�;�0u���r�k�R�6��$���Zl�8v�bj�r�5�:,X˗�&:�ęP����D�W����(=�7�q׀[��.��)�I}�.�<�ˮ���k�r��Ӫ���,o����R�Tђ;��9����T���n�vޚ!��P�+�ܣ%fn�rtЭ�6��ծ֥3m��<�{��[����\��(��'�]������X��듁\�Ԙ�p������˥m��հY;���t�U�0@��	���M=��K�o"�S�۸%\LA�K���E3�|�Ԩ��F>�V�7:�#��s����3�c*�c�c>m�q�z����c����� �p��p]��k�;wx���%[�L�+(�
�a+�3�.ӡ��u���.U�^�!������m��j�5c	�x��7�n��l��|��c{�O]D�
/�Rچ[b�:��'Ν�]&��ӎ��r��gn�V��#�ѳ����2P�_B��S��l�]���s����kmZf�e��q���� Gu%��驂�+;�j�t�"k�����)0�y#='��ne�UWQ�wB��ǲ��cZ�u�t�B����.�kI��]��R�����e�x`�\\޶k��P�P;䪴��Ku"4��H[�M�1FC/f]��M(�SHʢK�I8����ظ+�n赘Ĳթ۩�b�N`����e�Y��6(+P�\$�NE�RU���
�o�Y��U��F�N$C���չ!fuL���v ��f ]����1�9�%Hl#���ɻ�m�T��K=��,�t�.c8zUu쮭�����Zvܘ�:��P�s�CDՙ�w4AJ�P�(���+���ш�N�i�4P�M<��i`ۮa0j�o���Hr��]Jz�c��k����3V�A'LCU����Mȥ6E�ɄGU6T���|w�;�v~v��j�q�����۰9�W6|��p����(��d�����r�.:��q�T��n�{l-lva��6 m1s�ݴʹ�����,I!$�$ -M����` �t AP{���A[�w�?܄/D�H�
�����Ǟ�m���㖺�7[���u�sUJ���r�UUUUUUUUUUUUUUUUUUT�5UUUUT�UUUUUUUUUUUUUUUUUUUUUUU�x%Ŏ���u�g�9�Eؔ�s�w�qv�6�+�8��yA���]�������fC�N�[r��ly%X�q�m���tO\�S#���xɞ�/<GoZ9�Yz�9.�q�ν W�.�۬�wZ�\�ɛ�r�'�Jg=;ڻ{,�=�H�[\����\��h��cq]ٝ��]��gI�D�n����;����F�N��i�ܢ[�r�\�	����-h�gv����dͫ ���>%�q��n�mݲ����^m���j���ö^��Z融�m�l��
��R�p�"깶u9�
�u����^ӈ�b�v������f���4�b�\򑷞`��õىV��k\ܡpXv��wh�(�.�ꞻ{v{*���|l�d�<�tuۙb��u/��[�n{㠈n�n�7���M����e�iٶy�����	��8�<��֮`/W���{۶���C�EA��:�����u�;>�^d�gF:��<��-`��DP�� � ��"� �,� !��;3��s;���F�����Z����.�#�FW��gqԇ%�������Aln��-�G��c۫�jN{n��t�&�{7c[���I��9��Tj�p�������Z_e�L�sI�ݚ�������U��;";�n������p����rA�B��G3��_����A[�v�Z�d@��}a���(%Fڥ;�R.�6�v=��aQ:d��Ɯ�q�F���r������(�%=�9[��վ[��n�2*9��7zo8H�w��6���aT6���|��0H�/���Ԭ��{��̺�<�ucmX��*�y(V��,�ԕo^��^>�T��~�7#Wx�5.��z��z������~�եB�l�7�O�p6r-w��މ�齌M��vY�UaL�������sv�}�D�^񀛨4Ey���ȐT�1rnL�m��j�L��2iU��d�[-��kz�k7���9[s���k�-�h���{W�L�eMH�T�j�_�Nq�����������y8_f5� A�ˍ�]:3�����������7Z���<�m��S�O�1븝_mLc��~GE�h�z�b�/g�,���U�޿F�"�$�Uus2�F�q�-K�;����I�TL��G��dJ��n~O�����:��Ƃ��,���,���ѿ�����6�=ɬ3{E�#犞ߟ_f�5�T{C�!Ot���G��,k�����r�hx�vn�7D\���gc����9�n'x�v����)��������.�G1�v"�xwh"P5|�wz�g�x�)���շ/Ϗ��ـ��T3q��s�W3Zü��$
�Wѵ#j@R�XFGYxW/"�G_�9��������ս#��i�����Jrgen��4+o&[�M>�u暸bP$�r�{���G��S���{��.�юf��l@�I#��=Р޺�D�1�v�O�|t�b⯹g����^2����=ݽ	�y����h��M��D���xQ�E�-Έ�U�}+u��4�o���̉�L,`���O3*��A�Jܹ��j/�Vx!���!/�D�BNBa�2n6��v�ب˼��뤺F���}ð���0d
�?Y�7�.����v�.$=+=��^/�-{���+�ee�����	f%��qf۞�4����S���~^"���a�<7��G^ɿθܩ�uޫ2S�u��inx�V��#�����n3#	e~ʠ�m���{��zW�edQyH`�SW����Λ�ʨ!�}*�M;4^�R����Wc=t�I���Iv=i�Ѯ�Û�]�_atZ�nR[�n�"������'H��w<�:x�l<p�(r��<�^Ԇ]b������^�śF��/ѷ}~Z�8���.٬V|6z0�ʝ��/�B�c����+aJ��@�@�@�MS��gվ�>۬���ؽ��� @�4�R0��$�V��v^�s�>C��ِ[���O]ܿ!��"����H]E�����	�@����xz�So;�m���Ck�b<�u$����pԱ��v��4u�0��Aq{F��n��:�7��-�RU���$v��+��#Qy']��}�t<�.��T��rI�<���֦e�w�I�,�(�d��ަ<�F�4����0	V|��q�����oh�9����s"^�x�nm
�yMMU��o0��I�ΑU�y4��Au�#�FT�b"�������W��/s�;OSJxy���j\ڞ畑��Q���h�)~_��~fdݍl"��$�&���k����cr�<.>U��I���o������yl�|�~"f-�&*���1{��~��K�C=䭖#��h�W�\�x�[�ث^sH��3�3V������r�Q�|3Q��b:g��E�(���ː���q�r	*����4|e�h��w��?E�����9H7⧉}W���u�՗y\R�����e���ےH�
(T�G���>˻��D����0c>��[�f���#3/y�=��qCg��{~�����b�2��M��k2D��6��'�t��a8"=�6�pV�z�Z�v�z��O��:Nυ�;�����35��)F�i�w��z!^>"�d��Zaz�E��v"�%@�oۙ����p�	+����G}H�l�/�#rƁ�oH��g�3�*׳b0����s���j;�[	�0�
65˺��z�3^>�#��8�0��D���	6�m��6=�wܮ��2ݧJxq꼃�^�qk�<�{��)�Ɯ�/��qy[m���G
e���Av��'k&��F��T=�en��R��(�Kv�}�Y�Mp����ӛ��A-����mD�,d�,y�zJ�a:�b��-�AuڲxB�žI� ��7Eާ��g��^M��:n�-bZ�ѭ�S#n4����������������.d������@�:�^�\�Qvvө�Hή���=kb�b�ݼ�n�v,�=E�+�����+��.:��/E�l���q�9�`�ۮ�p�:#m��Gkb���q�i�*���M�g�WW���C�0�Ȇ�+�����Bv�ߔ�䨝GA���l�A�7r����%d�m׼�^�VP�'uaI[�7q��l�V��:��so9�D�݈TaS˽�V�yy���/�����<�����������E�!]4א�/:�/�7�ڻFm��uh�-.W"��{����z"�"��}&z�9�����Ai�!��Z�Z<�w7zM�l�}z1tے k\��lw���?�Wyw*���JҺ�#�S��v���������'�U��5�:zns���4GF�.Z�t�Yx��o�f�V!wŉ�n���tbᎵQeAs&	o�.�X��G+^�[��w1n��u��F�Ҕ���Kw���vzAll�5�s�$1]��Ъ�����;3o6Ze(M�3�}����{{sYң9F����݄��ZK^}NK$?��G����-��a�n������D7����P�S4LM���m�y?1�V� F���eA�����HB��s4K�7��Eb�nk��U<Yί��)4�n�e�"����RX�N�o^�cm֓�U;s�L�K���>v�6	rn�px��n�$��n:��ñ\7N�u�T�ὶ!�S��q��*�M0)	��S��e��8a�Y�؉�4��{y6	��b���2E��w���ڏY�-�|����+���[j2ё��3cۚK�=Nyx�z]
�ǯ}�a�C;=�P�E�K%�{Mz�ͻ��ax)k.
��E�܅���_�*�M�>�y,���-M��r�L��H�~!&��
[����CQJ�Bu�UJ�2����8�������mk��=P��lx4���t���*	3��R�ﮙ����́eP9�/��ӽS�ꨪ�8t�g<�l�'6h���ˮ�h~k��;^$�0�坏d��)��kE7E�g>�q�ϳ։$IC*P�g6�٘ݒ$:��F����7W�m����{��}ʍt�#��Xw��8!���G^PC1�y6�Y��ف���D�Y���;y�s˔v.tĻ�k�y����CV��F��Q�����J�t;���o�3�'�˪�3���nR!�GGV�-_���{�s[�,W��{�mv�N�T���\� ��-�s�	�7�MwH�P��V���S�&�FN��F����L#	9�F�e쎫6�"Wj����(b���ٚ�̅�wёI�=��J8`����$/�T�L:[M�J$�V��W<�nm�Q}����-ꕙ�蝉pѫ�{[��>X(*�6l<8{�����k�s}U�-�j��BD
�gg�CK���ò�9jl�ıf�=�����<%QUy��B��}��׵om;I'����i�[��ށ��^�𹞬5a*�F���I���Ӫ]�#�K�n*�`��Z0�2��IyQ�@��g`>]�EUM�����vy����ݐ��Z��z$�v���C+��T�m �-�����/���`T�\3����d�{Neu�j��>�3}m^|F[��[*�)��4�푆�M!��w:��ب`k���{g�Y:�b^vi�d�_j!}���|�{ޠo�RU��Y 2�fҀ� i������F�y�E`#��"@�~p�#)���u���ͬ=Y���Gsoc�И�t�ݎ��y�'7���Ze���u��/t��-$�9��U�e�����'R{fRF�O�ܫ;��woF���̾(��܆m��l>jz_rQ�{��{䫴����"�H�w��u����N���'����k���~6"F�6� ��aR��y�$ht�q��u8���.�<4q���E�$ ���q�N�F�F�k%o+��ϮxS��&:|�n=����HL����;U{��q��MC��i��MQ���L�r�n�f��"�5|�����
���D��Z(�[W��g�6/54�C�2��n�l�C�zs��T�4TK��������5%��0��{���ۈ&��%��Q�լJ�5P>˵�V��S�K����UE�LOɭ�{��G�bl*4�IH�X1D`MH�,���^���Zu� ����t|k��ƚ�6�}��fT��u��^��ϰ^a4�E��R�~�Jp)=�>m�9�B��z�h2�W0:5Z�˽�ۨ^9���a���O�~t��UZ�~��7�U$�C�jF��	�K����m��@��1U|+ym�ͮ������f �Vi�MZ�n���ӷ�tʬP�[���x���]S�� ��y�������*�UUUUUɻ;�ѣ�l���j^�G['o]n������]���8�]v�q*\n��O^Vޜn�n��{N͟g�=�>����\�����d�u�9��b�*K/*�ϕ`8�
�Ũ�;���F�;WW2���T� G���\�*.�-ғ��MD�w�"�(v*8=V�z�������o�p���kS�fK��K6������-�L�u_�g@�5(�p�T$&��Uj���{�ߜ܏�j�# �xD�v=����n�bE�-���:�F7m���Q�1�˸̺���!��+�x���6NF�3,J�����9���ݼ�2��z7����5 ��D���}o���7�����9Wc�����FN3�r��J�q�*���1Y�͝�v᪺�5��!���|��n#���Hԫԕm�%��ILCd�[M�+��<ney��b�k�0����uk�������M}�2wJ���%��/jL8g�;���D�T��)-�#8ĉ�kcd
#��v-���,��F	���-�v<�bWH�,ſ/>��������t}�<yb�ǲ���޿b��=�Fa	k^�&���ͫ��y;���½���d5�O����wWh�^�P�H3R���'q���#�B���.�Qu�s!��w2�h�B\���j�j������%'6�Jy��ŲQ88II:s�q�Msqm��:���͝�/Γ���	7�nB�q덄�kc�q��9+ۧt�L;�xp�
m�����)a�����1�����<�SB
�}�>���pJLSzӛ���&^�c]��HR	
��*Ubu�#��2C@�˭��ފ�y���=\��d=3�7����{�bz�\l��Z0A��P��*���	گ&q�Ň�2#a�$��d)�	�٬���\�<�1��s��ף���3sbd���w�g����U��w2��Rp��"5�WW�ե��nގR��z0���X��f���~������)8F\,s��)��8�� H���ж�2��w�Y��Ss��/�Z�N�j%����Bc)��:pW��q�{�iW�R	_��b$�Ed�������I��X7�y��N�62<����tF_��/���[덓�L
�����,ԛG��ha�9���]�=�
m	�m����Pt�c'	P@�K{_��c�ԉ�5�yu�R�����DD}Ͽ��� QQE ��D�{��k�w�z��Ԙ�Fm����eܘ�\���kp���Ѩ�u�w
���g��t�&IG[�Yl��W��N�����A�=:ݩ��In>�z�)c�q���꟪8�^�E6��\V'z�&Vv�d��TF��jc+� B+y���>�2�*�d-eǀk�U+�)�<��m��^�Y�����f�t��ˬQR��T�3���*Żӧ�Q5ؘGN�RVU=wS�ںr,�ר�9n�6:;�P����"+�]}�G�5�wkH(��qr|s3���7X&r[-�������d�
�p��>��@tטt�a��^�\��q��e�on�/�teG'���Ơ���p�\�Yu���\�Ll�־�왫6�P+_d=���=�i�]��[�+{7f`����/7e�1�ޱ�B5\9���<NVb��^ˡ�p��o*�⫺rr����p�v1�������oy�~��m��a}~�m�uȍ�fo4]�c�溦��ǭa_gL��V. h00��g�3�Qݖ<�&jk)J�d;{BsV^KH�[�7:���x���-�U�/4^�;gW',吭�\�T[�+��jK�6�,�78Ù�`��&��h_E�jY��M���W:�U-f������������f)��US�O����vU�W�T�@y2�]�
:�9
e�O�Wm���_��"�R�J�UU�g�U��UU!%QG�m�[����kv^�]ۈ�bW7&��Y����'v9���U��]�" x܇J�h��Ԝȕ��N2���kC�뢶���vL��t'c�b�%��{{^2bt��Y�\�͟78+���W��Z;u�gd$7[�&oa���b�]g/t�E��t{k���K\Vݍ�u�N��n�����m��[��r;�q�DbG�c�j���kv	��=�{�p�v�ɰt=�Ud�z��WS�a�79{r�>w=�ǇE�m��]>���^��l�-D�s�;c�w�p<l�nw%<���m��]�u��NwM���Ƶ�$�k;��hЃ>G�,�4�]�m۲�m�<c����K����r�qc=�ROiX�k�����箻M��<l���䈳-�G5aq��@`��$*����_���K6�|2*t�(��`7"� �����dɆ�S�ԉ�n���U�J��l�{x?.;Q�rz�n�ߟ�X뷉��$1���� !�T��J�|[�[1:�_�͉S<ڌ�o�mcn����O$}���K1�� SQ��!��Vc���k�w*:��0���㡱IV7�}%/��}�!4'?�:�u�ޤ�c�
�		%T���>;G(ES�ﾞ:+��C���8�N"�`���{Y�r�=ZvR<�[
�����D[С�y���;#%'�^�_
m��2)��{;>�̿n
��je|c��<�:�`i6�%�w���|�8��m�T��L�FKi_��)�N��w6���j�5B�,�[��_��>��j'�ڧ�&���r8�(�hw��o;��Zف�:q8����G���*�1��F`aȝm{6�&���ރ�.�b�ʂ4�#��n�Jʐx.��N�B޸�wsyj/����V�L������&a<�Pc�Ö��}�R>�p��)X�h�JQ%���tЯ��׍�jS1�!/��� ��`lhk�!�i�>~�τ�Re��y�b~f&�=��X��a��E���Wk�`�]�:G<�["�-=�9���Xa�-C���-R{ݼN�Xzh{�/�r�NKtxu7�ݭ��-�R�Mz���C�<'��b�2��:��Hs4$(5`;_\���1���&v"#���ǰ�XԶG�:`C�]d�y@�?��t�:�.@ C��=@�"�ha�AE	8�shZ����]ǁ~BB�aB2Co����~�8�
��ܒ8Ɂ��M� 7�p�\�Zu[u�!�Ը�̿� ��
���!�~J�Y����m�R
Ag��zJ��̕��_X�Y�?$����a��!R9p��)�H)-��+<d� ��� ���)i �
A@�*A`}��k'~Y��z��=`VAH)�>n1H) �
2fR
Aa�4���*AH,��P5�!�C�J�����f$C�� �1;C�}���/�)�@��ܤ��)R�<�wd���m�R
A@��1b�Y�2�dCz���y���ރ�VJ�R
AdjAA�N��)�0��
�) �]����+�<�A`t�N��$
�������37v�%d��P:F� �+R
� ���,��JʐY�� �1*��a��HyϺ�䂐R
Ad��y���|�ԝ$AHwi �>�& bT��) �j6ϐ+��u՘���+:��� �Ad�r�^��R�:I��!�a�
�̕���Y?!R
AH,��R'6�d��t��Y/��yh��AH)P��
AH)b�R
A@�VC-T�ä���R~\ �0����߿[ќ;'I!դ:��T��֤>�����|����u�I�AH)�R�AH(�`T��R�Ad�lĂ�S�����ѩ�{�AH) �,X��Y+��!�H)�R
AdX�
AH)l��Y>�,=�r�g�݁�R
Ad�V�Y�Y15�R
�Mꁌ��2T���d��
Ad�3)b���w)��f�!zۺAH,��Y3�1 �X"���d���7z��8p����*A`q*AH)�P�'2����8��B�M�p�Y �ѶAH) �,R���Y��H)!Z��)� �&{f$�?~��
N���~�s��@��!�fH,+
�R �>�0��Y �v� �
"ց�T#l��Y=eH(7��ra�pv���R �ZAH,�� �AH)��d=��|��E����?84�t�9�w�Ԃ�R �� �{��d����R ����? W�H(#l��_X �2V) �AI��AH,��`bAf�nk�(���1���
AH)d�jJ�Xw��3�
���Xo,1�R
IR �}�1 �t��}y� ����H)�����d̤��)������)��_3�:�ى��Z���}f$C��R���~.��=IY!ݤ��&2
AC�hv���i+
�R
�x��
AH)b�R'�ٌ��:@󮻶��Z9��}삐Y!���) �2��H,+
�S�H) �
Cm �Nq��3�g��7�\ԩ1�H(q%@�d~�
A@X���Y遯6�R
C�R
AH,���_������{�M@�f$��.����*AHm�
AH/l
�)���Xs��P:J�Y ���7�&$K�Y5 �,�s)�T�Y1�
Ad��R}� ����C�J�R%w��d��Y;��d~d���i'�~�c�w�Y<@�%H,��R
���
AH,풠,R
AH(ed6�
Ad�1 �>��r��-ߏG:�31>�xV��ѐM��Ss�(�2�y��j	o����j��2N�nN\qmu4z���1B�(��\QNI$�UUUUUUUs���۷<�[�Ms��裀���w2��C�qg��ͻBg�˷<z�����%]c+.|\�v��{\x�f���`+�G9��v-U������}`��]����j�ن]�6�@n����GN:��V�e��\ٷM����);@��R�I�+ � �Au'�\�{lR �% �{�Y5�[���������T����1 �q�D��X~aP��1��CRT��)s�����Xt��������Y/3"�Y� ��!Y��6�Ƥ�H(% ���H(�l��R
A@X�q%H,���dB����<d��������H"Ad��R���H) ���� �:����8���>eH,�Ь>aP*}��AIߪ�z~7�� �Lx�Rq�~`T��(x�b$��Y퀽e ����LH"AdN��t¤/��ۚ��m�!夨T��"AH,����
C�H)�R
� ������ɉ��e`��b���R
AHx�C�H,�y���߾<�7�5�R
A �k%w����
|�R
� �)�d�Y�1�d9���:eH,��Y9��h�Y �`T���Ԃ����,D��S�
�,�Z�&01��w���'�ʹ� ��J��
��� ���"C��9�
A@镬e �1�R�t�H,���P;Nw���u ���~|>37������+ ���,2����w���m��ι���c�6��7�7�(C�=K����ׅ��d���nιa��Ly��?E`���[ĿdA�p&B�ݔh�՟`xB� �L�t�"��X���1>�P���Q�+_��]͔�ѠY���!�A�������H�*6��:�ѩ� 0���%���ā��l��6�i�H�pZ�4H�	m�Qϴ~�k�3O��7i}�?@g�#�8uJ�81GYv"i�Q؄�����7��?�P�n�B��R��!�o-�k{��#��<@�L��A�+9�$ZD!�p�?D)�'���,5'~�GMm��2��3�Q;`�~Q�Vh� �r.�~Ҽ2yH�L�$}H��X���E�b#7�<��|?3���g�ŶV=ˏɉ�o�^�.�cG�X����O�>���n�3�{;�~.i�}�8��k<��.�R�̭c~�}U�dү^7��7RH���/l��v���C��G7F�6����f�|�C���[W��������Ξ^����sS�W��P� ��I`OQt����9QBE��?1�tc��
�!��r
��o�����$H�B�T�5n	S�ق�P��4s�Ga�I��4!㼰i�
/��G���M?�8z!�"�Cf�a`tc�����5R���W��]+(6�u�쀼ʮYΖ�@lH7��rWd�s��C���HWW3*m��`)����l�w0��d���	�&[g8(��o�g����,���䮪޵�ܤ]��Q�rn:���Fύ����l��4fg���*��]c����<pnp\k˯����}��w���~�s����������u�����l��f�;ނ��K�����Q�������[��CK?�d+́��>͂�v���,�9i�Fb2���8Q���g1�� H��z-֟�=�C��}�jj�������[�a��$�a�������v�7�y՘�쿶�Y{�b�~�v�uu�"��#
��Tv���m[� ����D@��c�m��iNw]�t�Z�M�<K����y�ZͮhQJۑ�K��-d58_���S}��O�s�I�t�o����l�#�<�?�*�~t���"�]H�q ���r��> ��)�	]���������z���Gټ25�߫�(G���#� �#��IE}�cR��pͭ��Y�Xt׏ɏ�3�S��A	>�&�ɞ�����TB��3áx���������B_���G ˻u�`�ˇes9��,�y��i�DEYB�؏�{J��P:|!�S�B��S��>�7��"�X�{
�~�?�^y_�6�i��dBa~7]�����i�t���=Ur>"�:O˗���*����˜�oWf��+�k�R�a庘�m8�l��{giP�g���^��}~��z�ԆeP����s�i��,���Ͼ�z>��󗇏�������k=[ek�>��.Ap���[���W�C0"f𿪈&,GL�ƨ�C����]u����w���K�8��4Gڿ��l?)D=j5v�MeN9���{L�YzeN'�'��*}qy�ˣ����u��c���.ѻ��p��b({eG;�Yh��~���"Ō�����^��\�V����Ϟ==�'����:|w�6�v�=�ʆ=����zy>������]ü	@���a�c)t��mWib�8K�����0�(���`*��Q���+�����"�,�;S6g�(������q��G����r1g��|�I��4��,��5�w��ͣ|<}�0۶�m�O�+�e��?ţ�U�%�Ì;���c��Ք�O����o��|�ѷ*�C2`���c�\���)�Q�g�?�������5 ٯ#�ĩǷ�W�+����y��o�bw�]��hԚ��,B�8�@�b<u��)���2�:���f��|�/vw痛�k5�_�fm�}\���9�0}������ ���e��o�Ws��B^W<�G�T_�Y��#c��!A�f���
 �&,>0�@F��!ڬ�_1/��ᥗ1���G���3T"Y�B!��4�߽�Z�y��{�|����B \�.ƻ":֣S�u��BR4�rb�G���/�a��懈dǌ�nx�憳���≈~s+�+��������������;�ߛ�" 8"�����=�ӫ�?�#�����؞��<�4��?���Q�q�����L��TIX�F�'��|:L]r���B�B(|D�*�G"�"#�ru�z�t��$�<�q
�k�nfN�wzo[�o����/����?wu�s}�?<q
�/ـ�����i�K򮡝�����(����y��}H���@��?J��&�1*�g� n&h����s�I��G�u(��M�d����0P�K?XXSį����`KkE�	�R�W��◗���̳���PS�3-+�;z���.*E�Xe��C�mS�����2:�$�۠����H`M�O��P"4�]v�e.(�}O��w��(�yay���lU����"j`wYdP��c�~`����D��L�7I�1����R�B@)S`�G�Q;LR�)v��n?k�%��r��0l�
�NזP\#�p��]^���ͫ�Aۋ��E�i�I"W��弱���r%v�+-��KІ�k�_^�.L۾O7bʆ�����?)z�Q�\�J㴊?$bG͵	�"�����c�t�pTd6XF��#@��t�y�m���t�����S�q�(�$�ԁ�K�#H��;��A�59]g,�d��l��tb'�E"�ק�y��3��c�T�1�Q�c!�E��f6�w"S`�� �vr��"ָ{����C��}�Nm^��&_���Zy��ju�r�-�Y�Z�-�qd�ˣR{���n�<��`���������y�:A�t�B��3����j�Di����=����1!��"����7<W�.��x�?p������܂�]�����X���FB�ƍ�b�Ơ���:,)1C�GȠ���6��*��>�q��8������x����H����)��i�{�qk:~�����XylƦ��4����s����}���٩�Y�՝��,?�3��N��/$��(�<AiRV�8y��}�<EȢ(l����.�ewv�C��^��~�ΙYZ����~J��b���b�P>�Q$F�0�U*8x|����5�����螪�@1�#�#�����}b� �ԋz� >"=���>4��F����T�G��ha���� #���P�釂�y�i`�_�����#(�D�����>t?{�ձCH�'<���ڷ���㿽��3�_ɩ�qK��>l��{em��������8~e|M�w�LMs�0�}��,��N�g�}v]nV�[r����t�1�Q�8��x�r�e�vnr�OɟK�w�wX�c���h4YID]����ȇ:�?��!�p�U��ԃ iD���
�!���n��k��D�,o��_/�+zc��)���ܸ�Ϯ��>�X��t�<AC�]g\�/���z�~3��s�	�>(���WuO�=�P��0X++�LO�w�p�YdI��N�F�S�0�jk70S̫�7N���;�e��ٮ�[}#��Մ9r4��8sR���~���j���������'��&S1���L�1�[�uns���(cv�]k2���ɤg۞�=	��p�Z�f�x���/���=�����z�[�kc���Ċ>l��=��qv�Z��n7j!��l��c/�z�\���.p^�C-���?8����������;��B���xP����Ea����9�_�LN��pX���"Dd�`QB;���b�����u}Po����>$���3DB��ȳ��s�[�w�������]�U��h����7�N�ܶ���Y�1��4~��~���[%�	8}�>��`����i�@����{��k;�m~�;��|�SĹΏ�1[�xG,������@H���y}�o���A����G�F��Z�iw01��u4����QL���,�n�y/W��=�w��
u���C��v;�.���wS���+�19�������U� �81� 3�1qF7òis�� �Ѥ��8��T�>"+�=FG� �)��L�������������v�v�;���s���㺙@��P��,��4"DH�a��W�ϯ���ѿ��ms����r���E1�>�Fb�\���#�Ɔ,�<��6�B(�,��dI��Ͼ�er��!�x�J��h>B�:3�?�����:p@`�n�����������3���ơݰ_6��VW���vy��۷&�Γ�T1�o����>�zMq?2���5����v�Ά�_��j�s.sx�������m����S�w���y|g��C�11�q���#D}��8@Fr���ND��V�(�"�:a�a��3�O�!q��-Q�q�5��v����͢�nn�::;���o�|z/����B���iV�)��������D�����3�հ��
����X��\����z�{�!�RU�]^��
���� %�� N0p�{��z7���'ĈA�H_1�d嚇�\\�ϳ<t�r�:`��6�:G(�XŴ�_���PT}�Fz�{��]ֻ��~]&�[��$}ʊp_Sv��E�2�u��ί�;�$�"'��	��q^䛕
�#F@�6�s����}�g�<sb*�Ɇ�[�9�M�?ˊ�<�0�c'���!ck���k�����/G�v��E�턹���h��Gi�����f�~Oܳ��+��~��_�/�~B�4`��5&���}
�c��$}��
?!h�k�a~��ozA���W0�i��T�����ںyw|�1�k8��V��>������0k5\�%c� �F���K���BCp��_BԾb,|G��Ɖ�Q���2���y�.gwf�b״��S�C��	P��c����{������c���>i#lY�p����o����Z�?����F���<�{է%Vʛb�����nn+tӽ�њ�_��~�� ���!6�E��P�/ ��z��z��8�=��pq?'�&�< {i�m~�C�@'�%����ڌ�����ۧ�aŲ��f`$�D���k��3���;��Z��-�!I6v����q����+���]��n!���n^�}xx�,�//r�J���O9���ϸ�_��0��c>���2�W,���}�7�oם'�.>&��eb�?5��W�����(ǂ̏����Y��j�ћ�ه�do� ���m�g���6�f�Nz:n�� �a4�_64���LX��"x`����<���>|}gܧ�ߝAC�N�?�#M��(��h�'ֿq�P���N�#�Q���hY����ߙ�J��|���o/�juqn{t���r9�F�����d	�6���]T�q�u��sq��Nm�u��\�&��Fq�mqwg �xL����r�>�1.�;t1��#g��������~�j�"
�a�����2�>�K����8��~�����*�:On�'��Ϻa���-�"5e�ݾ��	�ѩ?vǩ����_[��\2����s<>c� �Rb<#l��+ň�8p��]~�����m�G��Й� =�*�U���Ȣ�)ՕO`�,�I��g�b�͙3Z4z�CukF�y�d��IT�,Sm��F���A��EL�n�t*�����B����	M~�z��pk�51#���J�y�����[��6����Y����$@�(l�ģ�T��J����b,1�� ���׾���J�4S1 AQ�ā��q��c]@<F��ߓ��gL��ͫ�'�������'��:e׼�B,�#�TW�bvE���8�F2LCF;�;����~T����磼<q�>'ο��1�%g���@�S|�D�_P�>�>�QBG��S��/���Z��rΆ��3�ZeE��;w7��Y���w�Qw�.�~�?�Y^�^���ީ���~e��3�W��
�C�?0D������R+-{�UL3(��?���2m#�M�n@n�Uuy�b�I$H1M$��gǋ)t;k��҂�v��>~{ڿ:�g�`���u=��|�e���ٌ�|��핚��k���1]������C�1yD��l�!�����\���xN���1 |�wUEk��:�٧�'_�?���R����'#��gK��$$����m�L�5�5>��7d1z�[��ls���'�v���G�����EN�ML���S^&0Wn�~�O��t����;"�,�X��Ժ����<0�>��ň�gk��]�]Zo�G�b5��$�}C�{�`�`�A�(U��f/���pd_Rc��)ww��y`�f��'���`�mv���F�"��G� ��Y���p�����9��\��=���l����T���>^j8O�=�ȥq�Qcɉ�G��e[���&��k����G��,���v��m0��PA
E$Jp� �0�s� M��eD�E#�?�� 0�Ʒ���E�!�{�h|�!�X+���7:B�&���3��|��$E�P�3ݞyRH�6�&�it`��D�-і�V�82r�#��u@ӡj�L�/m��W{*<���(ޒ�c��Kl0i�N:�{��n)e��^����5Q�>0�3��6{��'��pF$,�0�:��	13UlY�	�y>_��V� �E�$}h���|�j7��9Y�Yh��|��(�>�$CD���hI~$�#��q��'�\ٵƏ�ؚ�}��6Q~��N��Q4>��P�t�������I*Ba��T.4I��y㗝�0�ō��M�ͼ񘕟�]^�����.3�����&�X��a��~C�}T&�E�>�"o9\7˳X.&.S�;�_߬��_��>4a�EX�#_}YiTy~��H�~#DALM�T>�o�H�CQ��GU��>8c��
^m/�	Ղ(̿����Q E�0ž+�gY=�e�������E"��]�1�ˌ�g��Dn���L"Q�5���lH:6CH3�$�Ssf?�?<��ђ�:���ӑ��DW�F8!�n�������`�'� ���I�}�9@�m�r��>CֳZ�k?%uƻ�3�#�������Yf�?�q��ETg�tM�T*Ȣ7c�	��'�d�v�'�<NǛy��,��rmz��i��MW&@�L��n�|�a?�����`:���D
:Y6���v[1HX�}"0X(�F� #�Tx#EGr�Ւ�v�ڪ�]x�\d�݋�ǿ��|����U��1}b4!Լ�Bc�=u������x�|�߹OYY��P@���O�
4w�0!p�؄#��(��
	���gd��"���	<�Mq�u��k���m8��}�5��u���t�[��ϙ^�g6��Qq;z�Ϟ������_p�r�f=e�ǈ�ݔ�#^�v�-���+�:H��?�l� &�+Q���0�#)Q�U������
2!��]2lO'g���d@Q�	��k�,�����Qdg �~��?}T��A�c���u�7�8���s��k��E��Xym�u�W&�U}5ݬ��FE,g3uW�����,��-��)g}¶i��}"LnK{f���Irqƥ���ޙ��C]����]�1/��� �!64��Y�/���,��	�:󞑝D�Â��o!�-Ƿ����2o�kVN'M��u�fu�xj��ofY����<������*�^S��2��`nj��sW�,/_[趋�#?:�Z�׬ntצ�X	1�������^hY����p]®��[����n
T�l���/�U�q�i�5's�x �TM�Pcgr37&]�êI/{Ge 4�}�(�]L��n����:����YO�f�d.u��\�Zg}۷�����S���3����X�R�WY��]�z� ��ou�O������9ڈWd�4��X������8(��9͋Fj3�����;)B�
���u���y�w�U蓷�V�ٔ���V�w�5ך�Z���v���[	��X��Sy������[յƴvZ�

$e]l�.*v��j����`�ɒӍ��Ov,/~Y̓
\ cr�����d�k�j�4�f����yV�oqɧ�y,���uWA�No8"�vC\yU0�*h��i�%*;p�Fo������ig'N]F��F-�)/�p< ����4:��dh��~3	���������U�:6쥵���
����UU�;�q5UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUqAQY��b-�K8뱎�{ ��6��1�n�>|����1�:8��Z�I��^��L`�eA�4m��;�ޢV7X�kud��%�IK�1�z���˺�p��{�,::2�7m�q=A�{'SXx8�0�����:��ݹ�T�&�O���N|���UN{o<u�<ӻ>���ݸ�R��Jx��p��n�[r���!����'uu�=u���w<������LZ��v)�v�u���7m'4�U��%z۫>�/9t�joF�ݏ7��뉺�����`�O�6����W%=�8�j��۱Y�V���oK�;�z���uჷV�jv��I�O����������]GU�=S��vz�8:݌1�,�m�ݹ�\]9�6�{�����vJ��6�/l��B�����[�	�v�Q:�p�v�5\cx��)�����8��%�h����3��pv��D�=�'^z�,ػ8{+�u��.�t�m��'=Y@�b	�;Qv�� ��۳UUUUUUUUUZ#��C�1�ݱ�l��=9�Iɘ�nNW��bƳ#pv�<>9S-��zޑ�`�v�X�F��N4*�n)�'�Gv9��r�t���n��s�<&��1D\�Ӳ�UYvl�)�=>Nڮ�'��]Y�%�������|%�qv`>ۂ��1$\�]������0�Q��b�D�,��B�Y�Ӣ�x��zq���N%gY_y�?��.��}��+�S�>!�_ ��B�ٌ��<0����L��ƁF��v~C�Lň�j$E�`��ƃL����F�6t�=����g��ڏ�ײ�e7�1a�,k��pn^��!z�F�/��������mQM��@��V��}��"�#�B�Kxʟ��R���J�\��Ż�C�4��{G"ϮVޫ" ���b�ܒƦ�O�>����<���;�Q�˽�S���s��*c+YR����3�����/�s���]�Ȫ�y��tä2��Tl�֚�->O\C�������T3�əN7oO��y��EF<ޕ� ���s��>�1<��I�D���H)2i~F�.�|-A뵕���1�cH�	M$�. ?�`'t�
1�p,27�姮rܧi����k�����ښ��̚�����|�����i�V� ����!��~#ULyɑ��H�|��9��6�ט"����q���;J!�qgie�̩Y�y@���N���m���tU�!Ö����R(E��L'|�#E�0�R[�ڎ	��k�h�����BDABI!�b'�@C�]	H�>�%�Y�� ��"��3�U֧�����1�?X���>"��XY�K����f�Ϳ������{t�;ŷc��a�`�i��m�r8p�>"��<����C7s����q�<~Ɜ� ������	�P����G��	��T�p|~l�����|E��H�}��m�W=��2J�u��k" �>��z�b�%�M[�')i��CO�B!�ш��z�MK�Q��h,�=�(3�rY���EZ�Q�ۏ�i���`���9�{߅ǈ�M��i����	��{<T�/v�ު�>3��ѧR�6��9E�ۼ妐�s�I=��O$���96\�>����݇�]Kt�zEy,۶�y۬�P�ޗ��a"�6�u!��|�<��h�z�\��q�|����vO�"v��$u����'���>�$|	O��88��K�ov����s�ܼ���+5�)��Ӊr���[g���^�eȇ#gM���	3;����GAC�DKT'�6�#М47��hB���W/�}P-,�0�B ��G��P��P�����|�ε ������a�1�E��>����p��&��)Q��EX�I��pza�(Ú���Zo�����]����q~m|X ��h"����=^� &�[��D�6~6p0�$
�#������N����c�ԗ�ߛ�����vu��;L���v�2���]O��o���g�x���9���*4���N��B(���B/�"Ϗp�Kd@��Rx}=~հ���q2��k�'�1����!�����
8bGoS�����<�u8˴^���\�����Y�7lͽ��n�մ�W\_n�c�<;��\%nݏA�>�`8h��X��&������B�?���#1i�B� ��@���4�*���Gp	��!��ǌ"��L���~��8�5�����M���Ѡ�e�u�.44��w`."��˘����q.ى��1y~uԊ���>�4�>jv�ۯ�1���'�S��&,n�Nc���#�B;}�&=��Kܟ�]��|�ϬX�!���V"~�k��3�����""��	�BG�%�Ewp�!p9!��N�+�nP���g��m���c�0'�N�O�1�C�G��(}�"1��>���c+3.%��5?2�C�O�U�*��DVD3��W	���wM�U��W�z�X��5����dFk�f���}����C�VD� ����PE�l�!�" ��ie}e�QD._�d@Y���dr�� ȼ�ϩ:_H�~�r,P�"�}��^h���eo	�#	�G�}��l�{&�غ��ּ#]:��B�eeH=i�e����&�T�?~8!i̥#�FǬF�v>�a6~@I���#��bB��}�����ʔ<(`�f@o��00.��$B {��JM>�pƥ����b��^0Cos���n}L��l�`�D�H��l|8*a���r_	����l&\@2> y��� �!�����<yJc�gV�Ƕ9f��?s��2����q<ef��d������{�{���F��ƣP�f�!�q@&�K��#$a�ГC1~��8�	���׾��+����o�]B�P�b�،B&��K�6G,�I�#>�'ňb��!�l����v���DN����9uz��-��u��մ��x\���E�i
�ن���(���K����ZN�6'R@�nFI!&��8�����rj-
����v�z�ʇi_�f&	��k8=e���~�^�&7�S������m*V_i��ǽ�15��l����`�I���z�L��Gz�,�T���$  ����?E�R�����w��b"��J�����΀�PI�O�ɚyH0'
	1(X��\+�O͂,� E`���ҍ��F�� �{^�*|���Yk�,�j��O�!v|�\:# D{�m}ͭ���a���x�jq�פ����ͥ�K7!،��
Oޡ{�%:/���SP�u{�]/�E�G�Yrf����L"��8p�#f����3U9���yGY�l��"�5�Ʉ>#��9�v���3��N{s�
�<��u�����?~#��b�!��B��˚C>�����V���O�,�ؙ;.�_/q�G#�x�L�%�a���H)JP�q�Yyo�� 08��:Q#�}?Q�	6��Ǟ���m��!���D�Y �&4�!����T;����ɍ[��ӊ�L���t����'���f���,�	D#H/�N�e��Eyq��FPL� R83{�Gw�k�Y�V����]�U����ث��;1�v��k�ŧ�h�?b���e�DXJ��/(��I��vǉ�4�Qن
�v��dݪ��c1Ƥ���9qIf3fe��F���M��]~�Pu�`���&��`B M�^�]�ñ����
(�R�>P#Ua�V^��H*"�P+>��{�~2I�}�dSi�%mUׯ��{��r����?B��Z��+kp���j:�.9�ɰԦ`�ly��s3��"W��1�2��A�sR�[U^��{	��<��u�iT���o>y�j��~D��A����\����k<S����Ў���g(�T�?I��ꛤ'�=b�R.mo�� �K�Er�Ѓ�/r������3wyGƇî��\0��P�;�@x��	`�x˾�U�G���E��w+�kE�~����R������_XAX��	�b��yz�7�L�wqr�[DL{��^��^R:��u��9������6Q���d�_x�wd��/3U����?|�}��ĺ2��	��p�p�T���y���U4��g6�XC�H�A�_@��1�'�LPH�oz��Ά|�ũ���EəGp���AP�%� 5�*��{�пt�>����F��}���]�*B��W�.�z��??P�2�D�Mм��j���L�ILD��{Lٞۃ������%�u�TB���Xj;�
>	b�s�vEM�3{s!�#"���''(�b�[�B�u�=�Q����8ݔ]~������������(�b��\Y�Z��_<�͵�����䄶��u</P���}}�p�SUUUUUUUUU��퇌�W��x�z�8y�=�;��9�}�\q����#g��k�1��r=��u�q���8A׵;\{m�5<e��`�m��&S���=��Q�ۗs�n�ָ	j���.�SI�f*�n�'E��8,a�iB7�݊ӨRSx�or�|梼��Jqu��\2��,�c���u��������.8����)�?�ą��/���>��Lk�[M{��1p]��*J<����i��kf����2mW�v<��P�OL��B}�b�B�]����g-U����}2/|�h��	���!�w�'�0��e��>"����}�`�^�VS�4�T�)8J+�����������r�ec�h�&�������ĝ�u�������儡�wb�+c���}^37dN��ts	�RtǁS�C��8��}�?��10�nz0��a罛�*���w.�!�6\��C.��`�����q{RU��Z��拓��wV��=�-��Wu%���qS�0�;��H��n��+{�'�ƻw�^R�y��d%ٖᄇ!2,���m:�\�A|�"��?��

y$.�_��m-ך�����V\�ǝ�������,٧t���ݱ����]�i��hUi�vZ���^���0�e��9�u�=٤���O��4m�����.����8�ݘߗL:��B���jQ7�1�bKi�Pl��2s��2R�n}�<q��o���T_vl�b�wݣ��S��p��bT�ڪ}q�Y � v��cީ~��-L��0p���9�8&U|�8|�p�ca_����S��b,���?r�n2���5�Py��V����nVR�eFP;��m̥����5rP����x#��}���g6��^ɹ�ʃy�\<t�;��M:���uњKc���=:m��]ih����ϒ�l��v�����?�����o��v�:�7<\#���)��nyU�/h�㳫��Ly�.�a����<��z����tUs��'�����M ���#�+�fG�T�c�8��lO���A�f�����8(��>��&Л׻�`�z6=g���I��ڤE���^��њ��y�M�q1.�f��z���c�q�b��t�E�
-{�}�z����t�b�3hq���.ʌٌ�s��uf���
����*n�E�T;u����Ur�I��3rn��(zO�wS�ភ��t�n����LD������6�qE#����c� �2�6���5�<X3�ꃕ.��ɚ��
 y�(̾�0:����.�c�f�6�
��S=R�|o���=�N�������q{���Ú��EWșJ[l1�c�A@��:�6�3"�n;�B�%k�9o�1(�l�"����>�9qX��3b6��3s�i�x��x��Bv����������x�o��yN��tמʪ�t����K#>�h,��1�1�P�T★�L���(�{���jY��ީO�)�\���'Y���=�߱�P�`xNl����ɯ���ֽpKS�\����(v�4����!z�f�y�6��{	�{�1�Y�Α���C�BP}0!s���F��/snST�u�_����e	��}7�i����[�#�<��"c,6�`�e��w]��(n�s&�X��a�yͮ��jW$ͭʻ�㏭�f��fd��W�M����ϼ��l��>�Ql�;�ޗnyW�۱�~�V\-�FЏ]-qČ��%\��K�G춨oQ��P��,/���)�X�,�d��k+Ѭ�U[d�$��
G�F��ߋ�'k����.DfzWa��Z�r�5�#WCdt-S����\N`7�1�Ab�\����AǏs��Xp�����G%)��06iԎ�.&DJ�'F��	Q�K�?���SUoVA��R�J��,�3Gn����qm�Ί�QJ`V����)���dI	 �U�O����/=�wѾ�A�F"i�*�v�֞�{t�t�֓)��͠���m���.���*���N���q�����zQ�ÀY9�v��3���6����t���[����E�΂\n�
}���&ױH��a�p J%���|�E_46dV��Vխ�"y�gOF��D�Ө�E{n9�R�4#���� 8�!������dl(\��M+�h�<�s����	�Q���x�s~�4�������Z�bd1�Y�7�n���اJ�C��*f=��a�R�ю��,��I��k�şw�����[%���t�\B �!�Nv�w���un=5�ˤ[86>q2�PQ��B�NJ��5˻M�"r. ���K��)�������B�9������E�a�@��J�Vm�7�J���:�}nMJxV�S0m����#w�yY��;tZ���}�y�7j�n_"_�'u^5]=�4�iի2��n׽����S�5�M����5����o��w�7WClZ�/�/L$��,e���"Ljn7�|
V��Y�>.s�]��}t���j�ð�%��y;4ꉱ|׻���B�`$�E��XgT�x�o�w�Cm�(.�fڂ����>�/�A�W<)�n�m��S;9:�]s��.$��М�p]>��s�K��#_�)\f-��2EJ�����sT�H����[4���6��߆��O6�4��~��d�%�A�X�G��#��{㶴�T2�qy�ஊ�!]����)U�<T����J\NM>I�������¨V��V��O�i��\���Z�)L���^T��kʴ8��PNA��`��Ѽ;����_<8�2�ys��E��m *�j�j���:�8�	F��<+h��^�Dv���Wm�3�׺Ƕ/��p-��dE:� �JUNj��	�̀SV�fd�hȹ���@�4�^Wq���}a�A�&B%$N(��Dd��NOzѓ7���齯:�O�ʯ�b��NY�K�����>�u"�aҴ����Go]ٌ��l�&���s�IM	�ĠdA~��U���r%Y�s��`��e�_X|���Q�C�&��rAW;��%}̏M�h��0��8�������tr6�a�� %.3�2�Z��<�L֓��Yj(_��S���C�W�nV}��������`bl�yk���}�w0LE�v�d�sn땊]���@r7Ep�<Gd�׼w_�����6���j���������5�kS����!�i�a��fm��k�����:.��p�8��@r<�8v�Cw�6|����p-��v�$�' �Θ�9�pe���ݷ� ��<x��s�3�W[Z�B�OHW\�]��OXsnw]�s�E�en��w�@"tIY���Fc��?�ꠧ@�����J���X~�+����V=�d�_KY����+�Ϗ�cEX��##iJ��;n�Z�<�V�����b��A���޻�����W�{��55�����A��;=���7[z�ę*9:��(z���]b�Ce�p�,(���9���w�����I�U��gg��.�bSٟ��?6�oli�s�]L�բ�6�LH��&Ǐk���Wݟ�����a|��Ѝ㕀�/��\�ZFYy���,V����;�V�x���mJ��3
����fx�p�EW&�@p�6����E���C��tsS�/��dS�6Zy�6�O޽7wq����$ˊwy0h�Lz�:��(�`�9aҞf��8�����H��T%s�7��b���%%�~o*�"[c%�Lz�-��F]�
��)l�>��R�o2��<F3>��hT���f�4+�i��:�n���]�g��z����!�o�v���A�r z	�~���c�6�y$��	��dyy�k���n�<s�=�&�h�U��8�u��fU;�x��"o���A�b�E ,?;#�ӟ	u�t5062��ӧ�S�0��:4UϰA:�+"hy)��QU.�ꇂ0A-*���.Q4.���*��Wy�/�*���SC�;���0Rlq���?P�GGv��J���G:T��J�٬=�����*�*�d@�zW�nU��Y�л��|��&�rlq�u�������z�i�|)���װY�E₹�f��G+b%�.'v�k�ۗ�M8�G&[����0yA������GnCtA����OY��d�jr��f�ζ�ׇ.!��j��}o���u��3d�������q%�����,:yp��@���%iUg	�J���E�#<�Ob���Q��4x����l>^��g��J�''z�߱;vzQ7 �|�kƧ7��p[���B���K;�Ά��7�wrAJ��m��}�_��f�A	8Q4�E2
/�	7 �;=��'��`������VOz�%�wB�Z<
4},��y��f���`��ą��X���W��lL�{�GOB�{{�)�^�����j��@�F�h�Ɇ�m����u��$�{�*D����j���R1��4�C����.���̈́��T����%l�k%��+�B��T�
���4����}�9g �UA}+���m����]I@[�ȇ�n�gw˓t����D������"Q���?#/���}��TY���J��J���P��H؆��q��'����-�zN�sY�^�JmbXI����h�Raf�����ؠ�t��B�H��{%R+���h�/8���݅;��āz̫y�}����H�c	��K�4A���� ��7�]���`�YFE H���4o�
�z6��H�J�7YՏ�Ȩ�
��e�.�Qr�E�3�м�uM%v�"r��]U)�AC6���Jc�D���SN��U���N�� �����������V��Omۭc��cn��uj{7�7�4r��!��U�<�dȦg3t��h����|/9[@]}�6i��@���vt�� ����8;�9�%��̗�6��]V�5,��v�����H��) ����4!�����B�ikU�xiM�uì�v�ܕ��E�E���{N�V$���N�Q���m�+�[�S1"�f=��jt�r�>�:�䂷��М*H�u*��{f�kQ�D:�f#�ٖ�S�
����} � VL���F�yyٓ[[9�Ƥ��h�զ��v�t���Xw���wOkE[�����X�(@�6J�7�2tnዲ-l�E���6�]���o����Q�ϋ�YH���+�,�fv��>��%�W�B�ɼ����&C�b˦^����5��[/qv_��i,��4�r���˹�A�Ҷ�4�F^�YEY������á�/N$ܻ{;���f�\֌�yqI"�*�8�U~Q��z�G^o41�w�i��P�bw)w�''�6�$�i�9*��jYy:FH(�*}��kշ�ŦU.��<ڢ���I�ȯ��7k�F��}i3`�w_UE|�t��K7Q��GC��r{V�\��תb���`�>��
�Hu�x�7d�1ԭdU�����j��4gm��UǮ�Y���B;4+���p㌿�o��ߛ��YLg�����RZ�jU�U��UR��h��q)���>،n^��c�ݫ9�����&
��ԞLj3�d�J(���=i��6��r�vN�X9��&����kdm�n��q��W<᪷�j�DNv��� 1������������bs.�>�����Xޥ��q��v�c]�������Zg��N��1�'c[7��7R/n�6��u���:�Uu;����	����Ƒ��zƌv˷��.�zGI�b�s>��y䤉�]��wm#�`�gq�&G=��w
Z����|��z�3ӻn��ۂ7	޶	���=�"���u�>�k�&¸��1�r˂ם��vLt�{=h��7 ��vc��TPy��Od�ͅ�tv뺅�I'ruݟu^Cu�G�nn��)���#�CCzn���Y�J|bO܋��Z�g��!'�����(�C�����Ki�	����b���s�����8`H"E4�&\�ى#��z�#[������;q%�EkY�Ѿ���o医*�h���}��,3���[��Ys[���2s��Q$������e$�n0"����;�&��8�r��z���Ao��J���<��L|� ��E2y&>�c�����sT�f}�3N���ƨ1�i����h��p�ݶ��{�k]��]��b'ݍ��M"I6�A8m���m��/��k����cx�J����:��T�h�=��\�J%m��j�E�n�#m�^8����F|;Z���]���0�V�T�R3p��k}�yf�01!MM�=Lzo�'�9((�ϰ@�B� ��"��/��`"��`������ߒ���YH�'C���S���-�oy��5wu��h�W���!�e�������iA"/�?V�X"F�J�\I��]��{����������b)��Y�%I؝�.�
� 1O�����)�د6T�f��GU7.\U�}q!#��$�L����Y���������m�73e�펟_bg`��e�~��n6��)	4%#�;w��]����U�9]����@�Q$�L�WL����$'PE����2N\f��;S���wO�y�f��g
q|��]����z�h�"�j}��?~�;:���ՙY��s&o���0$��9��xC�=�:��o�v=A�I��3 \����"i�L��۲�ϩ��#�{+�.뇌$E3�wR�0��-�Vm�i��n��V�K-�J_,'L6Vj��9n���k�6�I
�����R�\�6Cd�izuX�
8L�Fh�^��Q-Q�m�Ōi��=�[D|�߉�X�5{�<������{�1~���9b�|=j6Z�>/3�+�C3��O��s�^L80�c�B�ҿ? RDK�R�":/]=Y�nD�`\�XU�+g3D 8���x�VR��c�����N�=�6c)>"]�Jٱc�,X��z�`�I�a��ϴ��6#�J��!�%�2�����z�+��KF���0�����f��!D��%�A-����u��T���!�"n��Qb4���ӗ�{Z��,#/��(�>K;���JV�uӏk�m&�M2+#��L�-Ic���m�<�7�{<�[��]5[���wo���\˧%�����>$��V)��Q	�u򃺞�A^��ɖ8}͟Eۑ��I���@��+��2ڛ+}�o^ɗ{�M��6��iN�2�����c�4Zr+Ԉ�jR��>V�Ox��|�)0�|�L��Lc,�+�sy躘���s�ж-z2��:�l5�=<t-�NU*��r2�6'��1C�O�M�d�M�JI�Na�X��u��Z�J��e�޾�vݷko�Nē ��������.��>,�Aݚ����������QF��㇚qhsge5�N۞�]�Io[�g,!ʚN+�:v�糺�4�1�v�<yj�j3v��������;<��-�T]��D��:�-�����:3p��T�p��<ܗZ<��hϓ�]n��ͤ����dB�`2w�j	���U|��I]��h}��JU�۷��.����q.�{\x#u2�{��u���wdAI-*�^��\~+���"Mr�Ys����ؼ}�1��OHdK^�J2�0L�4XxS��g����t
AۯU1���O�y4� ���zb�ZkO��r��M�2d1�qvH�x�f�|�f�o��%�+�ϪEr�z%G���%/_^�
V�s"i&��ו�*>q��L՛�}�^�tw_�"e�x��S`C�7�^U�[��@��x�ʩ��z�[^��1}DI=�$�X簽φ_��|�?���=yD� ^B�ZP����K�O���*+f���RM�<����~�J�9��!��W�b�=��t�2$�0�t�(P�\M#.�9{m�n�L�T+*��`2��H-5�.����ʪ~������!� �%�O�A]#�jg��Ȭ26y�����!g��ɩ���}�n���!I3A�a���bݒ�-[Ͷ �� E%]��-�R��)غ��|�j��yT��&t�wi�G�f~M��;w�o����#g[x��E���m�ȹ:VΌ-�*.���D���Y�ht]{j���+�g���p<>p�7N1X۽��=��9N�ܰB�j��=����3�p���������9�{�^L\pb��{��<��j���Pظ�����+>���u۶}��݌��L�lb�]�Ndg��v9	؃����IXڳf6��_����_OS�[�$��0t�k����n����JE���o��hTi�:�0u0�g�П��;j`!��C��䖇�+ݲ���#�	��鐑P��E�[�̱�|�
	�U�d_�8`�Ic.�N���>-S�� �釔D�H<ۣ��BZ=�#O����S�a�?6��qDٜ��tB9��1D��[""�q	���JO���@�#�kA�	�/z�3	�{2��6���5?���̣�=#L{Qm�So�V��
�ɉ���I�,���z���_Ei�D[�jG���/B���U(c�
n�1"ی�"�ȰG�}T�D��g�>iJ�|�0+@�'˟�0z�1� �y�)�K�	/��:�V�s�gV�)��������ڡ�4C�t~9GE�C���c���cx0��|�2/
�_hތ���Z���$�}�O�q0�\��j�� 1�b�v_���aK}C꟬�D�J9�K�UG��H{�Ŀ�1F��~Y�k�ŋ��D���Ȳ;s�NdU��{��4}�����4Y-�$�����b�C<�○q2b-{d�*
Cմ�b�zW����3g��KK��HG�p��0j�$�H�[�
6�ڻ�ܱ��I�Æ���u���X�+z{\��B�M(!앳)��L#B�ɏ#�����H?S�4e���)+_(]x(^�s�ELY��$c!P-"�GH�"O�|��/�S����9D��,���5Q�Gq���=}/RU�4ʆ 10�u �����/yH�ߋ�~j��R�D����H]�5蝥e�3�t�n���VZ�	vǓ[2�-۬��~ǋP?]b��4��
����ϗ+�9�YN8�1��p"RQ�#��K�K�Xm'�H��&AA�}�;o&�8#cs��B��m�xD�E��+\\i���	qEBe
�uTP�Dr�X�ju�Qh<��@���|˪����O�Zv�,��չEA�ȓ,�$��/�6]x�$�����a^FqP%���q��F=����R&��o�^���pȓYN�']�^���2�3	}�����&o��UV&2���ܖ�@�7��ާ�/Ƽ��D�62�xo��z�*�4F��i<��4Ҧ�1s�b���E JϽs�#e��`�y��� $�E�#�@�eH�
�pZI{=�[�2] ������ o{�!(ѷJA�|l�
��d.����
Kݽ���b{��M�w>6�ۊp�i��1���=r�
:�vM�	lW[oqNIR-8�%�B�*��L�=�܁�=�8.���ܓM}L��O�ЦÆ�d��_R��"��T���<�@�p���\E��3�[L�n{o�IGV �~�(ƌ����y�@��\X�z(�����O��$�H�rI!�{�No]�+�=*�Z)��!�����ò����_�;"�e�����pLH�̡�����ca"e���Z(�jg����f��#˃G|�T̀���)�i3
J�'J#�C`�\^M����\W+~�{��CV����fWsH#/�p���<���f`�s�� ��ևtyw}�>W5��ي^M�2i
#�3�˳m3�P"C�K:jH�W�����Q����y�'�Yg �J��0Uy,��O����٥		sa��k�&��^B3�+|ÓH�J"_�E5�i �Äi��a��>���SfTP�&ʕ�En�����8>��2e�N�f�z�7[�xL���󠃥�E��_�X���{{�*D�0R���ؗ"!ox��c�~1�}���G�Y�5�V8Sϳ�x`C�=<�~��������o������Da�5t���GZ�v�߼C�ᆓ@޲s�5z��u�Ź�ɮԩm�X6U�:3��*;QU��d���̫�w;S��cy��QC�`kUUUUUUUUUu�<�v72�'b��&NΥ8��<]��Z�m�9O;6m��[UuP̙h��4݌��;��l��Tϩ;s�O�`�����:͸C�,��{n��3c&9�j½lKUe�Ӷ��sͧ��g�����ca�����F_~�c�R���{/�>q�3&�¡Y��~:?��K�X#�G�;r��G�5�"�O� �F`�v�i��Rk��(�J�;��)=i%7)=S8����Ż�d��X�>�[���kW�}X���*���CÜ~H��=�-gp����_i���4]���%,ϝ��КXD��&C�#1��=��9��6�k,�0I�_h!ߐs���{�]�|��uc�"gy��"mY#0�Dw���z&Z�O���b^�#�9������E.�V�͸���b8�H�wߛ;MP!#�a^�ۓ�%��'O��Ǆ
ҩ��H�u�N�C�^v�`�^O�xR��BS0��B*["`5��ɋ�0j�Y�ĝհq��W����o8�y����zsG�yђ�t�J��ü"/���k�X���)���o$�A��iN;,<�Ÿ��G':Dg�X����`C#W.�d��j)���t�ƮD,��J�cª�Z8fp* �?���m�B����߾_C#�����a�5X�#P���!�����J*U��l�7?Vd��2; M���`�ܒ�؅��v��o_<K�eõ�w���wi�$����P�AW��x�U�]Ks�5��<׺w݇WWn�Zmئ��t�y�3���5����I:�����śN]��o\�륳��\�X�7#0���!@ۀ��?�p4�W쟨DZF1�Q��H�_��%0*s}������ޯ��ו�>��"��I2.���-Իܯ���S�+a�:�j�ʭ?Y���1rm+���*'���n;�N����4��R�~�H��'��1(�ܧ�p����K\F4����?/�D@�Rp�(�����v�+�(D�@���İI�C�������v�jH�j�����jxW�<�El��n�[�ԃ��$?�d�:���I�W�&��1��dř:xD�����c_@}>��y��3�A���Ǖ��NyH���q��
�Kx�g�$��{<U2�U��y�8�·ـu��P�����i캪�	%�o�L,zv+��{.�8��Ԯ^�É{�-��aQ����Y��s�B��-��y_S����E��+��%t�ǁ��ݕCQ���Ȧ���3/�Þ=H�5@�1O���i���$�1h��ծ�=� �#�����Mw��H����p�pd��p�:`�������+�EG�*��mO�U��9��@��@h�tH��� �|M��0��WU����3��}��o�w�z�}�.y�ۍ��	��9G�D'F��<�~��a�p(�
%rS7z:�ʪ�=��Z}W��l�S�P>�)e�`𪾊�ۺ�ҿ�?7�ߛ~!��t�Q1�5$�������>�1�7:)>�w����q�@ �Q�qGq#�p(�R�Z�K���ɯ>�j�<�	\��nG�q�K߼�E/Ŏ}�??�|����ֈ�9�#ٷ�1YTN�t�w�H}U���¨Q9�;P=�M��?5�v"�o�<�wv�*i$�m���4W�Ǵ��h�S��ƦC��n����<�R%h����Q��zb�1���:&%qPy��3wd��<)V�����3�/)�Oe ���@!���rk�RbF�5���܅��5g�a�A�������A�B/���T�! -3�ë��{Ve1��X�;�b����h?���	T�A�9�9�F��o���sl�}7hۿ@��fN�1|s��OZf��GWWg�G���3������������P��=O0k�	pJ��A*��󑦡��<c�G�6�ތK�CC��ٺ������!��p_v�Uy��X��4��6�\[�y�|��Ȧ3�+�{]�6��阍�D7%��[g��id�
4�ǑI8���������	��3"c�k~uQp�tl�� �}�I�֍:���m��t 3��F_��G<����;�\Lw�:⌕��I\Ў�,����P!o����l�U<P��rHV�+s��g��5��ƽ8?ɸ�%	Q�K\Λ0�b|��٤^���m�1V��6x��TGG�>�8�[�P@n&�z�x��a#��Dm�U���Ic�3V�ު���{DL��m�x#e�|]�H7�`g����Tj C�N��Uj���(��9�`��8':�ٛ�In0tG�|=x����f�=~MuwaG��/�R`��亁�Q1I�~�Ҷ|���S̰�l�/�iK��+�J�C �P�D�(˩���>�$����`۪8ō�n(�
U���d�A�7O���\���q7a����E"���{f�)<3_`AX�,�5
�m��y'�Έ�����\p���.:YK#�u�����'�%��6_��I)�&7�Mڈ�X���[�T#��E�g���4|�ed_�&�_,���^TOۺ�<�g��y��ڡv
QM@7��|&
��Fr��F� �i�ͪĎnװ��l�{�P������|4�s���ܡb��x;����3�Pjl��E�E���Gί9��^�2l���y��uv�(�9F���ҭ�Ĉ�@Nc�!4{?\����؝��uDi�u�*�٤�a�fca��
]����z�<ڵ�X{3oL�)�-�B`2d����U���H�T6��.�w�Iv�ݩ����"�]��� W\��z��;��&�eq�ӇMν��r��c'D��{^�&����$��zÂYGxɍ;��[]�JB�[��밖3y���kY�9�c3f�p�:*ouѕδ�K]��3�]��)[:�������XW�J�ţ�t�g�(��i�U�1̼T��U�8��N˾��w6���<MoQ�k��T�VҮ�.��]}{f"��̱��å[���;�P�z�	�N�*�b�r��R��P�,gi�o����miR��uV�fN�,��t�;�L��h��E�78���:l.��d��"-�>�X@����JWq*���`�]O6P�±�Nk�.h������U�m��NʂwV�˶6Ԇ��z˺<�9�����v޻��C]ۏWI.�e���0�])ύv�͌w^�����=�)W�uu����p%ld3;�\,���ѝ�%�⫃).�G@��*�(iG( @�P,��$�!M�5UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU$rZ�`�\�Q$P���5ɶ�r���x����N���	�e,�\�[uܚ�ǂ�6�n�niլ�]]��;�EvŹ�ܥ�ݺ���vpt�/6����s�bCv��6�ۢ�l��;=[<�ϓc(F����N�J8�.��u�]�qg��l]����m�/F胎w�!,E���qV���hQE��<�1q��qɯaE���]�Oi�v77T�[b�qu.���u]YH]p�/*����njSe�����9\dGn�ɸ��ݱ��'��;p�`7n۴#RuX��g�g�'c/�1;�ۃ.�h���;�n�'<d�����,P� g6���N���w�u����&����5��0s].��r����yi����s��c��N(;.�=���n��vמ��["�)��N:A̭!/��<�3���&c�=��D�R�����ɞ'g�˛���q��;���Lmˇ�G=qp�I��=���F;.�����M��z�,��
������������;r�uظ뗦��q��8�bK�e9����:�N����cc���n��V��^�$`4�.��l=
��^;���cB���z�έ�4�Vڶz[֞:}���[c���F��n�1�u`[����=���;�7q��U��!��6e�(p7�_ .��ʏh�� \�c��L�B'ʹ��oOi�.!�c;]��L��NV��Q���,,�i�I��L@�oF
쫕�r�ý�
����@"'8��1-1[R|
�/���
Ef�%�G��-��'�jߎ�B��*�13T"����W,�#���Q5*1�#����w��}C7}3�f23���0)���#7�Hi�v����{��\vVXiJd��&�J�T��n�.E��?|��vBg��n�][�ގ����;��6Lx��p.�&u����
]�����j}9uv�.!�����o~�?�����6�tl�"���+q�oD�lQ
�wsY�a/)ۍ����u^-�G��^��w�C��������:$-���C���KI!�]�<0��dx�Εr�`��EXM�".R��a1y�K�S��3UI�Aq��NOOf����$c�M�Y�ñ][���i)��k^.8s�X�e��(�`}w^�||��F��{3�eϝ.��aG:�C�[!eS���|ba��o!���. u;{������0�]��/-R	nN��v�x#���-�R��y���[�uZ�A����7a�ѽ�t�u.o�I�/�kE���޻c#��O]�Zݺ|�ݗ�0�z�!�!�K���`9#��׋2AC�H���ۘu�Ŭ���r��.�(����R�ϳj��H@��Q$�~�Zx��4��Ĩ:�R#ƍ/t���񰕝�Ƿ�
�N9��]а��@UzD�kcQ�ܸ\�O�f���$㦡��ń[nn�)�ˋ=��g���k�	Fl'!2�5qFG����LV��b�������w� ��G��L.09T��ӎ
�5�5xl4�!	E>|gݥm�@��4i[*D(��]��Q@g���ܐ�7����Q�����Ǵ(�A��it�\��؂c;�j�����r�9aKx��*��'������_�LW.���f=��n+�0�NMůI>�^.���q�y]�^��<ty�#���]C���\�'P�0
��[<6�UFф/�{^d<���ѩ�AT��ZTK��V�d2Iɸ�t���1�,].%<Kz:��󿭟iS9I�( h�c��U4ޑ��x#�̏n�H�j��^̖Eu��C,���kr�&"0��t�a�C��)��c����u�������׬��R��;�3,Y����"��R`fލF��C��ei�Zzo�|�osm��;�k�z��-}Z��"�z��
p�9��V��֐�D��P*K\-��X�>�/�k�hB�0��Z�P�u���o�/�|�C!P��HF�M�`��0�i�K�!�)��3�D �{���x5�T!&��uTz��b��
ѿ��7C>�������݅��D�"��'ސH�!No�����<>Nt�
�
ՂJc�)Nw*� B�����G{���`���*�jO��Г�,�#��"���L@�/�xy�v&���^���5��j�;��⻢���SQ"'Ǭ�	�FSLl������5�w���y���[��9%���S%���P�Ɋ{>�n2$O��$�w4��/G�#�P�R%Z4ߘI�L���I�Y郧�GQ���z��mԵ�����u�x����{r9���Sl�O��^6n�*MӉֶ���Z�b�u�XγQ��.��l׽�c��q�Ҽc��Sd�����j)�Swcä��F��b��2�~J~n�^�%�l!,�">v��kf�۞ �\�D������:�p� l�n]��<e�*t$9��4Š�:�ny��ٗ`�u���2�}Zv��.v(��j�l�����BS��y�UgUVyW	����Twxuk�hZ���J��y�������r?��.i2I;�3�hGU�O޸�����T]�a��^x� =�2��K ��2���AA3�Zv�}�ē��Ok�����[n�gյ�ĥ�$�l	\v�#u��c�^�"c��-��-�R����f�n�Y���d������Vm7S�j��N�C��?f8�l�F5!�ʕ�uX}ǐ�oPd�$2N,39>t"w��~�Nv��5�3fh��}Ogm	ApDѺJGj��|��i��.)�D���ΦGqg�>���R��}R,��ͱ��*#��<1�:�	غ#������7�*�#
؋Ҿ�;}�J��u>����xAw-��(ާ ��q���]�:wٹͧ������a�  hI�L��-��<A����;B
����\5H�3#�#��w����̰����vc4�O��⬈ֲ�<3}:kpI��;��s�s~�b2���$��-�yeJ��\�F�y���V<�|g6����ӈ�*�Z���ӏ��Ĥiq�D��;i�@��P��q�G�#��^O!��m�P87>��=6v۾z����.����:]E�3x�fMΩr%m�����4%uK
���-��3��V�����������3y{-�������m2��P��0TLv�fV�qd���r�ںTKt��|��s��[���[l����<i{c9���wS�p��wcs�������띞v�G����n�λ�]�a�m]Z<�g�+T��%�g]��(F��n���lj��
�vMY��_I�Ʀ��}�t��������2�\�o�n�z;� ��f�~(�v ��毱z������~��\�/[�_���£>���vǡē�&�6z�D?���ގ����.���tҬw�z6��Ȓ]��&��I�}��*Ϧh�V]����0o���GbM53�:U=�+��2�8O�l�>�aE�;�p���4��BH'?g��:}m�}=���k�R�7H�j0X5��θQ턻�Pw���gн~��J[���8�4��+��>�SꑊjĽ���po\H|�Sm挂h������A��
�K�R _It(#�� ϸ$��ۥ��zX�{�)��G��Qt~'��>�� p����A�s[��G�yg�|}	J�HY$�1��hN�f�������ѳΤ��[��<<��-�s*z�w/m��PtyT�i�����k�0��\j�����/���N{�ל���H��ٙ�E�c��(��O�0��߆��b�����暽p9�֏��ǅ�Db坸2>������z�1W\��z�v1\i5n�3�q�\7�5r���ʲŖ9���ī����]�8[
0��d5�0p>9t{^��Q�/[�⩺��,�q�kq���i�R7b�sgնv��cR粬�',�ص-�p4̂8c%�#����byK��0z������}��iw�ڛL������~�/+pn��O[��N05�P�r���F	��i��:��4�'r<��y�>���B%�Qء�Q��z�ǫ���L�f(9lp�(�QM�#
C?\�vp�o�1X��c�#�����Q�Y�`�������q��G��C~��9��s�9H"cƳ��}4��p{�����U���S�qRM�V�3�?�
#��<��J���BN�u��fv���	Z&�i�g��ٳ��f{�!�������ǈQ[��J�sH���lć��^��K:����B��m�Kd�Xp�PC�9Ħ�����ըV�+�V_�,\k�w�C��gq��ӥ&��Q���==��~<�U绑�����N�O]�JT�J���PkG��*��(<�M6S������p�a�"6N��Ӻ��ʇv���k"ђع�����i>�f����>�f�e����7 "���.	l Ȧ0A������ �P*�&"$)K�A�w6}��>���{�u�n��&�V)D�(Q�2�XJo�3���h��zK���.��|�t��x���:��Qo3w|�M��]*��;@�����#w0o�ȱ
r�*�)�I��G�������:�["^��Kb��+�K��~o�ׇQs�ߧ�L%U�죖�����
fZ���wn�x�][ˁ�^�D��BG���E���,�Gjκ�0*
�[z!���h�W_��2�J�9�+"�L��EjǇr&G[�?��v4��
���w�.=9�ǐ��6(T_���>�����Ve�%`m�.C2����şR�L82SiG��L'��^PQ�-�.I�ꡚ��7f��v��c־���g@wj�;s����?@Dp����q�� ���]%�����[/��V��
*m�z��`gB�g�3;��AD�֐�����-�y�t�N2�]��'�8�z�M�BN�� �@����7���k�{��:���i��C�zpP�ٛ��{�0"��?!<z�cO�aAp�$��^�w!�Z=
�;�Y�V^5�onK�����ۉ�O/7��|,\{h�s\��w����0�>�+��7��7uN>��x<�Xn����Ap. ���K����Q���Mf�Q=4��0:x _A�t����Y6[���E���4�{�Q��ޔ��#\�`ח�y=�)$[�j,FK�����G��nP� �T{M�HN�Aa��ؗq��˯)�۱�q��Lşr��^�pބ�x�����v�(d��E�6�v�V�m܆i��Ƴsp�fAI!31%����}�Bi+���^�k����r6_�C�B����og�VRWJW��`'m��_R`�j��_��b!ߪ����B�V+w�P7��u)��=
�~n�
�O�Q<�R��A�Q�3U�T_R�H�0�Cݨ��|�r5b��i�;艸C���O鐠I����R�$Ct���`9l�T�dF�%���N�>����ȶV�x!�==�n�vCJ7&W�s�}��p�����[���}��n�������4S!D����0�S���ɥU�9 �T)�&b�s�}Q+�ہ@�}�NDc{��~O)������!xL1��i�	�h3?@Fc�-fD��n_q��k�n��U��@�C��q�J�1�i�:����x��B��Ov�)'Z�Ca6���iw�T��L�~m��5�~eTTz��N��}�R��Mf�۶���Ҧ����a3r��e����+�=�����UEC���������������j�L=v�pz���ݷ	�]��k;Z��v;���!&=qV��L��#����F�𹹀{�:1�.7[��l��s��m�6�$��u��n����8G7�����Gu7e�[�c�UpY��SۡN	9Զ�%O=*���:�ҙ���<�fA�4��-��[�A�,�(xk�U��7p���fo�u�7$S��u�-z d�� d���{�{6W�p9��F�lNn����ο�Kbtq;�����9������D��z}�����c�%d�v.w]_�ؕ�N0�M<��;��L��U@Q�K�?�<�A/_Θ�6�L�M
�E��ǺaD�b^��q!�+j3ʍ�p�2��	n4|��qv/7ya�_y[Y��i�����k/LO>�L�����,�h���������W��c�\ܢ=EL]y��l��n�����W]���F%��_��}1|ߧ�?q��M��@Wa�
g�{�l�n��A��
��:fXU��L2�ˉq���e�}�,���}�lWle�B%R3�j0�`5wH�,�7�V�J��%�i!�LIF������zV�=*-.�g�>=f�=�W�E,V�"z�=�5��(p��!R�&�}��I�}��\�#�	d8pR(*ɟ]L5K�WFT�]���5�C�en{���:�.N�r����쇺�We�e�`{�j&S��ѝC7y�����f`0G�+if�I0��L���}�ԱӣR݈0�V:v��:��Ǉh�\��j���X-�KO����6}O<� VȮ��`9�ٛru��Y��Z�qs��
^�NXPؒt��~b'y���^e��Ҭ�bSo�������U*��>�g|���6�P"�2Qힼ(�@Na���{���5���p�M��:
65P#4.�ܯ��~�Ջ������������ll\o*~uwZ�a$R?�Я��bb�&Z�N��I7!�,#�e�iV!=퇰����Ac��i�ELn�ާ�Q����w_?"�|�_��l���ߦн�E�Q�x3"�����sFEK�0��*���{@nҋ\�7��6%�j<����rc�{Pd=D5��E��u6�t�u�_������=�u�%A2��"J~kr��usJ-ۜ��vy�ۀ�n&^�<v���V��4}�|�L�g�,=�sZ����z�*��>���\�u>�d����5f6���t�;�k}��Z�F�l�2�C$/���wm��`<h��C��
�%}��eA�#�^����U�1�f�N����{�W8	:�71����ȼ���ŤDx��t�R("�2�2}u����<�?!�A���������~����f᥁s��e�^��"�v�T9�R�S����/pʅ�y+�Ç-��0uɇihc.�kT���P�D�_2�۝Ԉ�_)��c9�����Vֹ�wjĦ�F�Ҵ��n��c��'a[7�R��@4N���:����,����QP����K��.�d��B����1�]Jx�̦�T�o���b!¶�_�&�\�r��I�������v�*U��wһ�X��wWw�]gSX��p�+nkm��p�w�	�R��c���0u0�W1x:U�[Y�zDo�Rv��0�F�u�;���(����w:���q�P���T�*!�7�۸K���ʸ��w�~�ϻQ����̽�>aQG�Sچ�a 1W���\�]&w8,39��<�	�Y��Yӷ�^�q�ת�2�M�ۜ����إ}�ab�������+,3Wn��Y1YNF���+4`C7%��=���Y|�N��o���{�{{nA���Sr�Z�8�s$
v������ �^i"�v�ܜ,��ReM���p��W+\�u�&�i }�X�&b~n3��9����QM]<��Y"��LRZz��{�j�[�1�,3%&:Ȍ�7r���ɷ�B��:�l��+Tΐ���5@���\��<4��2/��G)���8�ϡ��jn�aƘV��R˝̽f�n����N�@�4����W�b�u�@�����u Z몥Z�V�U���
y&V�Sf.[Ul[��R|=�{u\,��3��U��Eݼ�wnM�lm�S�Ȓ�z2���v�a����	��N0��u��-�C�n9۞�У�;'^Zۛ�w�Fv�T��ۖ�n�*q�[v�P���u{\qf8��O2�]����m����g�9�oӱ&�d�=i	�=�]��R�c[=z�f�;r�wn��ur�s�G>��+q��Aa���A/l�Cf�����μ�1�+>�$�"0l�[��/���)��v�{��qƑٔ�7%y����_2��㸴�VwA�!���[��4Y��EQE+�c.*����L��ڦ��i��SGG]�\��	�Z��͸�ͷ9�.���۫+F�K���v�F��W�l��un.~|���-��mR�i�θ��m���_�t4xMeUO����������GX�(~ַTH~���FG�&
7� ~_~���G�ꃮ�U��A����fA.Ԋ7����\�+{�Θ%����^�is�q�2T��<E�~�[}�����yI��˼��uX�
G�BdfD�o�rѻUWU	��G���^�xڭ��s��(���vg�A3�I��|��w�O�~wQ׌���)J,K��k�Gfm!�=�,�!-(N-�v7V7H�B��r=�՘%�l4A5�-x1��aG����=Ų-�j��B@��8�;]��w�}!�Q2kՋQi�I���~��U��չ��J�h�j��g�����阮1�qz.�3���M��z���L�2�x�B�p˪b��Ю*�j�ʏ!�91�J�&��3�d�B�P�'�
�1��N��ޝ��/�/�k���S�ر�o/n���ߜϱ���>��N�]����/wG�
����б�#�V+���ŋ7��m��E�K��!��F���+�/e/��f뺠H���Tܵ���xcҮ���~����=wkf]�h�n)���J��N����]j�l}բPt��r�T�X�`�n�+bU�s.�����~�h�[��ʸ��h&lÎ_խkekeh�&����1�߮��Dl��O-X��G�*�l-��~8q�0訾��>�q�*7�]�<�I�F>]?D�3�6߾�<KT�{�ck~8>�ߪ��lc�)�K<t��^.�q�-H���m��;?1���	��O����k�z��GW��3�/LH����q����ƍ�YY����|1�Ny�t/s`?{�yLruf�|׏�\�D�F����U}TiįΤ���m���?b���>��Y>�ơ&)���@�}���}B��ۦ����Q�Ph�T璘�?��*x=L$��r��4jueH�o�^�I�H�����6��z۟,����Zd�Q��:VS_.�=��"��i$�x�z a���������5��;,z�3���-GJb�ۛ.n��}�?{���c�:��O�QP�f��H}��:��x�+��z�8� �sr2��.^^��^>��UW;�V���L۳��k�Jaq\mH�!JT���
��fS�b<R��b$�����ciˎ��#�#�e-|���y�t*5���\��
:�~�ΔDK�AԂ�0t�!w���e�f�ǝt}C��y��.(�H�㛐-�P5);V��(���(-ǈ�������q�v�������������#�/mN��Ÿ�Ȟy�nv6w30�����혌�]��\ n�1z��w]�ƽlnM��@;��l���M��Hh�޴<A۪���;���ǃ��l
\QU�e�1m�ۛ�;W.1k�3n���:�;"�\$�k~,��1;�M��Q��.&(2����*	�WV��s�SU��Z�ĳ���Ax�/v�눪Yg��6���7���Q��D�U��g��T�pょ�3�����u�݄�u�C����B��0uԛȧ�$k6�O�oLm�w�O$\=����#�VW�i�sW �*��4ww�����<��\xM���V�{�+����FY�Q��LV�e>x}0`�r�1�����ˠ�����s(o��
$�� *������gÑ����m�'l��Jg.����}~(�>_e\��
���'��A�EZ}AS�WB�}u��?7c��Z��_[�ݘi��,�Q�Ĉ~ޯ�e�,����g�8�}T��t3��VTN���\�lVx�>�3A��Fm�Cz���댘�\��O����?l�i�`ޯ��.w�ϟ�����|�e�Н `��f�h��vmp��[�>ӧze�������G�Oƨ.i������B�e{m�U���w�1;0��j�l/�:5���[OX�[|d`�(�e�L!^����7��(����7K^/K��vyvf�2����9f�N5��i0�S��e�ee���1�H:7jȡ�zR�Kx6�#$�@�n�9��5��h�v�{{%gn����O3�U�8�v�<޸�ܪ���n�R�o</4�[l�@lS�@�0H0��p� ���|���c��\]9ҕB�����{Tl��p�p�H��{tGu�lsk���B�� i��� �v!������gk�ٗ�~	}�:�𺪖����'�(�T�Q���
{0�⛑��w�wZ�zD���X�B>��eW{)�=$��8Rd�䙀�`�1=B�����+�����V�a��]
��B�v�܃)����sB�=y�y�����l�V� �5</n%��J���~�#Vs8���<�`vP[�#�`��}G�e�Kc�w
���4�.����3�E�xr�����Aue�U�+ʧy��S�t�Y�6��h�S0�qMׯw�O)���R��+��r&�hF��A|���Wyu�}W�����&�c+ގL��|�m�ݻv*��-`�@���%��gz����'�|��
gs�D������GOu-��Y������n�������ف�1u�=����g�T�簦S,��}�wCP�����%��FN���`J�s�C��u��f���Iæ����p��[l�����D�wY��rZ-��koidUx0��9�Რ"�݇��r��{��a��u������j}*�&a'���1���aFA6�����������z��\!¿�w����|�w�0N��
ʱ�
��a�Tr��1"t��ݢ�J�F�i�.+ǫsP;t-����bs����p3u�ʂQT4�[�q��g�^�JJ��a���V�A�_�_�{wIi��_y��ܹk��z6x��\�/�����!�������^U��γ(��m�ńl����8�r�^���>�;�b㰗Px�hC��F�MzL(��W�#��ocܪ���01���.cp�h�/>�4f�;S�#iA?4��>��x
��ͪ��sp"�h�8!��4B��������]?{��EZ�+c���N͌�Z�1w��2j��1�����Nd4���{��!�j7c�u572.3^X�s�.�4O�r�*��,#�3��'s:
�qB��<T]f\4S�Z	�$z�����kz��Q��������3ۋO]q�z�����ۂA�w:�v�]ji��Ψ|�}�U������G�c�֩����i<���v�
�%M
�˂N��z*ro�\����*��z��u&���;]�A�7����I�ߛ���Wg��I�f�(YQ��R��d����*Q���񧹒�8��[v�kԸz.�(���)� њ�����wp"f����g[1.a�X��ȋ��,oq�8��ҭ�$\?����P`�Q��f-��==�֙�
OB�m���X˟�����5`�U�s�V{0M�v(m��K�:�ħ6������ �%����Q�|�e�u��OGf�-I�!�g�0m�>]z�a[����8O]%߶I�����N:ωj}��U���MݡВv�D�Ԁ���̍�F�=��c��W��c�@�i��>�v8����Y�O1���D/Y�<�Ŕ(��",�,�\���s	�7�o}��:��s�@�[�]����=��.k�U��
�+� ��@$��D�et�{%���qca;_����<|v\��qN���*,�_6����,ъ�ii�Vz7�S~��}T�"KYz�.��RSǕ�2� ����׏��?� ��*'����Tg�Dh|������p�샶��e:}�ax��s�.Ouam-rD�{� �������f��&e�Y���]d���f����x��xoz���wY]J���t�[5�R5{����o�4�UUUUUUUUU�:l..���.���N3��Ҽ��U�CJ��������ՔCJ��8�ٞwPs�8�s\=�p<��k���q���uT��ݞպ���3�]�qjwWZrn9u�UvK�R�kp����x.R�@�Xά״Dy�����_>�x��^:Ѹ�����7j��z��&�Ǻ5�K?��z�{���V�(����Ed�-��",`�cg]�f��3a�
C�ۡ����**ͺ�"us���;����#��Dq�8m>��\.J�T`�®3�"�s��")��b���}����n�	����uǨ�����u�\=D��B��8�2W���e�}�p)��oQ�7pU
	����fyC8�a=��fl��䏀$��"���% Fx�~��ΕB+\(��u\�A�b�U���r��g�Ct���u�����fɖC��Bm��H���;ۂW�D��rVsC� ��4��U+.�8Ps��D��B�'O�;Skש�n��Q^5?+�a�(�U�FBN亅"w5��7��.;@�U▶�q����u�$�œ,b.2����	�dV*�[ېگT��wb)��2v��� �;槊�N.�R�C�=�+�3�@��U��ci����t8m�6�P�>�J�[��ZR�8 G��X��f�n}�zvyY���[��b�'�;�V��R�t�b�9��b�m��_��T.��Ӻ��5��W��El������Li�"����G�݆S��3۶�3�kg��P�ں��x�vue7
Whx�b��.L�[�5yr�\iy�� ܻ�	F�1X0��l�#Mw������?�P�t���y}��_�1SO�Քo���i�1335���V}�<�������E M|A�H��A���l��hM2����Y�{��;Ղf҂#�9�{�<7��+;����͕U������vՃ^��w�!�YPZ]������K�Z�/7o>�����۹N��s'F�!K�7�DP�cw�W���E}	�ͮ���9�Vt�<�Өs�T�t[	�z˄�8a��� �a��Z%�a,�k震R���L_TC´��}��O���p>��{��jf��]���D1�.~�2���}SE�^�J�H�dƈ@6�7j�H���Og�#�kl+�8ATV@�,<�r��J�2\vzV�����Թ�2�Ey�]��⟠1�Q�FQ�q�qΆ������U��S�PÉ'���J������{�s.����U=�*ڏe�/�ƺ������{�Kz���^��!�����v?zMhn��)���Ћ���(�s+�Z��OvL'�OꤧA��1��S�ݯE٧��"��֩9~��P��!�:�Y2ţ@��\����1]H�mi�8г'�W;��և<��K�����z�><���gs[M>Z%:*A�:��&Rk\
D4ײzv�w�0��U������H���`��HC9�nM�ޯEb�cd��~�����L>Hu����鐯��`�/c��5��{*�~ák8I�ʸD����|�o�	Q��zH��;�O�����5�����P#T�`��j$<C}�l�/h}���H{�J�u
��|�(`�ˤ�8	b�B�nڌ\�AW0/n}:y.e�&��`�p�tJ��q�|I�c|�ʠ�/=�v�>�xy��U��ħo*D֡sL�ui����;xWz�d3��)�����Z�<8/q�f:�.n�hq�����7��}xcOdh�*�Ջ���H��ӣm�yY�\6u.�t"��q�`I�	�k�aB�
��Ǫ.�S��O�gQ�³����U��MUGͫ�qP�ᒽ��%��]�ZԾ��TS��a�0��Gt?��w{w��Qn$�i�bp$��BL��ο[��/�ٹ�c(z;�k�v��;�B�H�8	q]��EE��w?@�kgS�3 ��}V:��s0�`W������u����*єýC���$�)�gNg���#7,<\y�_�����قr��q�0�7��O���"�[_�S��	A�&^��k�ws����u���7�ۼ5@�!h}���?���q�{}�i&s�^0A�L��t�a}�}Rv��'���\2��&���Q��G��P��迻5������M��aAJ,���FE���5��ۥ��a�f���
�#4�t���5�_�A��Ο>J���,�TN$T�.�i��2����OU{�d����M�xU��8,O�|j�U��5,��������$US���[���v����3�	�L?���}ϴ�sW>����1���	đ��j�;�Ep��q�*n2�;��fcn+��Ɇ31��l��Xk���h�yW�v�9R&c�
��@�(��[���ff�����B�'�.�R����������M~箽8a�����>��ұ3<;�ދb���o�h����+A����0��D8���q��2%س"oڙ��\c���[ŧ�1�u��:�P�����Z'���ݮ']�}7y�n5T�������/s|`���)�ͻ�B�N�������hn������nk�"������q)��-(�� r�`�lƫo��#X�x��j%%n:w]5d�&7�������#��.�3��!U�l���ZX���PUի+���3e���'WI7���8k8�C�]<��c�*�Ư�JE�p`Ǥ���ԥ*�B�s��RD4�=�,qm�U���!a��;x5��`P���^t��^���f�}�Ϋ��"�'j�e�̂���k�D�8�����3c������[���a��������R��3��UaTAu�q3��ښ8�?ȧ�|0<E�wP�i��Q����
h㳵h7w@ܽ�F@�aw.���k��R�6�^�7*wɔ�Km��$�:����FUl�N�7��d��Q��G'�t$�.&>6	��7U��O���m�����y��u���3t�;]M�Xq-ެ�J�t*�7:�䭍�)ֶ�J:W#�]K�镐�WW�K	�������s��:�79ҒK)i�ُgv#�,-���Fn�;�u��Y��6s�/����{Z&#(��.gI����'V����t� �[�z�mD�z�,}�)��An�\�L�W*�	��bq^�*{.J�kd�NV�)G)�«�
�u����[�6Z��5qgO��djG,��Ҷ�fB\��!=հs�9Z��������������������������������������������������w.Ǝ�����B<4�۞���/%Y�x:�;��;=\��4C3�gG� ����v��;u��yxc�M�Ϣ��F[/x4����;;fƞ4x�*���=����G0I����B�Ѱ�X��f�枭��8���\�N��×/l���	���<s�l����p	�@�q��k�;km�s�s�S�ɱu��u��=���u��]�����t�mDfʝ�����J8y��떺w8�+va|�<�ç\Z�۷\^I��[���\��۲jۮ�i�O�v&�ެۀ;Y�����:��kx]v��m7.Ʈ;A�8�O��od��g�L�s��E�z�p�U�&K�y��՜'\�`-�[����l��TTnv��f<s��n--��o�Ev�b���]��(�v)
��g[gN;����z�xQWvPN�mݭ�	�q��c��� <�8���t�9��v�B�6����w�C��ÐA�`��Uq�&ц�R��j�;��2�7an�s�6�][��=N���8]C�����Y;�٪���������m��]��[�=��.9�q�v�q����A�n�U��mB��3��n��s�3�.��M��F�4�cqə��;E�S�q���lz�j�n�VnW����W�9œ\i�;[������d��=د+�)qe�nt7'k�E�����`;_P���ΐ`Q�����_Ҡ�����bOH��N��v�yw��OM��2�J�7�&�o��Q#ޞ��ʛ��~ټ ��!��q5*���������P����S����+VϽ[3[�$"t_�u�h�;�꫌V���Bp����S�S�)�0����\
Ӭ=�����"�e��7��hLGaG��ɪ�q=[ɔ���-ҍ>�u�Aԉ
`5_O���s�O���!����u{��Ӌ����Αp����rn����T�'��4Tzq�T��fht-3��{�jV�Ys�E�31{�'M�O_���Y�ƙP�(�KkD�6x[����q"(E_n�{<��~���0����UQ��pб�n|�*��^�@���v)5��a�ǥ���o�#U�k�xm��n6�u�v�th ���8,��c��w����Fq���<��3�l�� �3y��]�_���
���F�-�8{��E;X�ߌ�Twq8�D�)P��vP���^����l�P9d��S��yZ˖��M��$��\K�R�s N��u<=���yr�K8���/6�c�t<��\��E�*�it�#��2	����t52z�m�lڛ\u��\ʞ�Ls��,a75<m[���O�\?�wξNt�'S�l��/i�!����B-Pa���olO9�jߥ�Ǌ�H���.$}�|�Q<`I�i���4e���Tp���#Ň�B�����)�ݛ�v��t|�D�����[}���3=cǸe	u�mA|N���ty�e\P���@��b7e=� �`�����(�H���(%�4�"H��
����]�M�g*cd����, b��O��}��^:ׂ��ͮ��tz7|�6�t\i��s�3�3N��\�8��|����܇��1V���ԝ��0����^-"'�GT˪�g��(co�^̃h�`�Hd0��yD3.��t�:]-YUX��I+�/��;;�:�m��N�����Pe�A�H���It%G�:�f5P��}V��ø>�#�?]+��wl�+v��m�u��Q����z�����A.	K�=?�
I8�NsI��Z��㎶}�+�����Z��D�V�����$�>Y�����1���^R�L6�,�p�sOi�J5ް�D�~��Xk��}x3���_����j���'u;z�����=�-m��i<�4�7[��ъyp$&2��h�#���L(��S�_9��b������tQ-�>����i	�&��:�L��.^�4�)�A]��wA
?Sx;�JpG_�)��Ԕ/@��������8e�ݻm6A��P�^Oq`�̐�J�c�3��g�87�	rA�>���8��Ҩ$%E$_�o��Q�ܫ�P
��}�ޣ���{G��������{��zU���0���?c"!:���u~��rZ�Ou&ԇ�lm$�����M�I�V�\�{hNl82�.4\B.��3����8t��Ip^&*\ms5lT�C�nބz��Qn�T��J�3]>�W5smw�<(y�����YaRp %�E�� �n����o�z���_�ۍ�Ճ%�������^s; S��\���u����:F|D��ى �D���N!Y�)	e6�_\�1,�@a/yL^�L_:�n|,G�҈:�/yϷ�Ί�>j��A�%xˎ���gCm��Z��K���ڇ�t�]��_���}���G�*�&�x�`��ɂ���ȴ�$CLW��j�L����e]��|q���1&;�w=�%ڸ�8]W�j�32�F�agcI<�.���LudLp�֍����:f��вNn���o��,g7wl�������5��u�6�Ao�d�V��B��ݎW�,���;7�����ܻPD��D��;'��h�&r�'y�]�BCÇ�r���=���ա�Ǩ�� ���#h��J���%,��lk�`%Wk����X�R ��i^B%�����n����!�ǭD��K�
�C�;ǁS4�˒��\:�Aڹq�koR'X�Z^�[�rhFF�e�q#�dO�B|�ٻT=�lr���B��U髿\�{��W�D��T5O�U�@`���R������d�D�I'n�Ї�;tT'�$L�$YZG]�9ٞ�h�j�n�@�qC�z=�Gy�òuRa��M��B�f���4�w� ���+&h�E|�@e�F���r�+o��@�, ��B@R1���e�i�^ln�Q���Tn�|Xʎv������h�My��l^�]�n�x���~�|���X����bB`�4�d~-��>��ut�F@ &���?4�B�O���S+gٞ��SÐH��V+>���i�9�ܾ�o ,�/�z%��\�U��f�*QF	��>I�qRӋ �_.T6+����5�@<.�i^w��LXys��-�����|�B[HMUUUUUUUUUV��l��e�-�G����Ѳ�	�ݱg{*'eJ=�zh���&]h좝��<i:xh7$)�$���-[n��d�\q�u�65�-�7S��HŭY�q͸��G���rd����氓�bT�3i�7ݓ�g���M\�Z����?p��;!|�D���Y��迏��J˥�����H]Cە�_��(���B�`l��$T�ͅw����jI1C<f�?���3�SR������6}�O�|y�4u"ϱ��ܬ�(�zK���Vy#	�/=�T�� _�Q|v���ٱ�f�DZ��4$F�(>vW�v|`GA�'������/
��MWc�)(I��mPωa��?cŤEbF����f	�Pa���ь���O�4ō�]fDFp�s�n&n�tNy�A��.�3��0����������V�ܓr�1wb�������-�0��<X�3W�ݵ��r��v��n���3_��:X�Ԯc���\��7��;��E�a��d���7�r��M�(�$�"��Ĺ ڵ8��ý��6KA1�����6�[��`!��Ϝ�(i2��Иܨ�T�X�P=��Lʾ逓�^�t��ŞY�zLz��-����d��{�97G��\09�]t��I#z����|�����QN����m�rI֋�p�)�ofϲ;"�r������x�jGQ�u�F�ʙ)��4��U"�B���tATO��=$
�H]jڮ;S�?���~zs�ݍ-;g�+���X�e��{��`6����*n+�.8v�;���G�m]f/%�� 
��DO��S������?��*W�_���Z>��B/y�-J�4q�Bn��6z�� =�]��l�n
��uΩ�� ���Eۨ����Xqb��u������q0u�5u>��o���=�$�)z-	E�+�9)�pC�,��U�-���UN�p/�p�B�(�2�aFDP����5.*���K��D�����d�&�Ͻ�1u���On��ΌLڄ2p�vl���a y����O��6 D�?��E�߿Z���0@y?�Ÿq�ԯt���#}O6� ~�f��Z����z����-i�T�ߐ򹉫�]�Y� j;^��n[p<��{��͢�s�L뭳D�M�d	�������>vU<�T:��O3fP;�;��P�z4������e ����9�	$"
�3Mh��d���	"��7�9<�<
\U�u!�(��2�b��T�FR��ǚ�-�`���C��U����7U�	7�?}�<<S�Q�K�eˀ��?i��\'��y>�Y�E��}���"��{g�֊}"S���Ȅ��y�����,삫pv5n�]1M`�]8:�=�w�h����3�T��˫��imɹ�~����ໃ%�g~pq�5ɝi[)Qh8Jק�u�wA�����(��#`l�� ��JF�����/���V�ڣ&��'�FΨN�u��7�\:0��+�߽ ���PD;�&�Ja
��[�ǝoyf��s�g|�A8�O-���?A��#�	Ed)Lb��^W3����#�l�HS�5�����=�@��$")��
e	
C'+�(����m��mu���v�D��9�x��^Xܜ��Vb|r;��o4f�l�&�z�:ɇ`/.{��˜���:!e_Sa7n��g\�n�ǪSpC��em�ENn���4v*>�e�b����ߕ����.���SK*�_�OK���yx���.���F{0FKn_�x8��ٯ�������ՙjLmة3�]#'��c*�{�95��v��}�G>c�W����c�W�m�M6��/{�E>���=���bY��<��v��uI�1l6�}�s�[|�s�'�/�5�<� ��B�;F&���>��g�����4UQ�\n���i��dAe̈���ψ��o�q=�\�M�̓���\�	� \v1WzS�W}�C˜��^������+���%_N��d�h( J�깯�ƃ�N�Vy���/�d,j�8�N�[tR�4D�.�������b�-��Q<�V���������T1�$��K�LͶ!��C�i�j�E�a�;'���櫪���+|t�"sgJo������z;m!8s�V�!�T��ٰ2V!�nf{�x$�O;�+pmG�K�2���Q��f%�x��c���X���N��q*-���jkMvS��& ����1�V}�8����]<�v����;)V"�(����%��"�Pq{��ϧGn�ϴp݋�E�'&���sd���������P�A��W5b����	��wv��@�X��|݋;����9�&��~?���~���k�f�L=fZH�fj�lOF(��!�����k�^Z7@]ț��9I��j�gP'+�*��(ա�ɮF~�H��T������{����8/OQA�|`D�>~ݸ�r>��ӏ]ч?"0�~��{=�NqC٨2إ(������ӱ!������B�\R�hQ�{�Ƃ�D���Qq�%�7r������BJ$%$�I$�I$������75ã����k`��cnP���q!���mu���n']�I����İg�x�p�=��ݵa�C�k�����x����M���r�m����-ͲE�a�\�Wq����c|M��v�̜�Wl��tt��G��@����~�OW�a^�1?���&�2�FW��wQ^��g��*�V��X��ᔈ,͡^�Q-1~���ߺ��z�=f���� S������p~����:���g���l�2k����8㍤=���u��	���;��1���$DR���w=���,��p�(�}�o������1S	D��Q_b��]>��q�%�14�w �6~��M��љ�D�+�=�Va��9�����Zyn�%f{;��b���l�P!�r@�I�
Y!��^<��e���6fp�v���E�XG���m�;<U�n/ni��Q�1��
�ڨzlH�2M�8����TϹ�D����}�Ww1�~^��R���V�������ז�M=��F,��=�*b���<ہ#�S�[���9�r��T�x�%8D ��m&"j޿a����6k�����W�+s��1�hKA�<gHܦ]�،^��5p�^W=�$��7G��b%5��IL�9�V]��ش�ƭ~�j�VjF� ���$.��|lt��G��{0��a�W���l�7�6�t�����5SLEk�A_;���L�gs��;&��V룖���|��m�X����־<�o�{S	���:x�Sf�$Nض�I���U�����lQE���EԱ�?��> WH����K�+�r��k�_GBN�9vrO��ж�_�<��B`�����c|�`S\xtڊ<u_mU�����sgl���#�z���b�z��2n�A�Z�D���-/\͹����
L��J���Z�[����߿��Tļ�*U]v6�A�����������E1�������!{C���ν+,�D���>A�~��}v(m��͎Q]��dk�Bx͎�%�1�blp�-�=�S]~FX
����%�ث�%��X�=�b`�4�P���u_����C3>��
��!�8-ٍ���z��^҉U�a����BB}��P���n�k����dD�;��U�t���'�¸3�wJDO;įM)�-��y�����.�r�|�i4�S �c�y�j�i����1׽B$S�A�4�l*~��=����/9�	O��4�	�0�ۏT���G����?��C`���"��n�uT+ɭI)��C}߄�,`U�k���:��@��3�R
Q,ӵ�����'�v�[��S�w�u��zsHn��c޹}��'�]<U��Q�μ�-�6��D��ιE�Ĳ'u���������k�cC"+��z5(.n�)��ɫt5Ue�"��\��bn��'�s�������5�z5K��U��gc����ws=�@
����a˚2vMd	�[x�$��n���-���D�׺s��rL܊U�
���9��N�9��#נM����m2��	n�Y�nf���)�7�hf�wq����t��Uq��Ǹ;�����]�gS���BY	�
�Mu�I1�/����YN28�
���t����fS�����)��:�>㗬7aU�h�U��4K���8Yլ޲h�mN@���\+D�W,i,f������gS��ȷi��,�+\�Y7��O������3����Iԛ[�����Xs�z����-�#�L(N�ܻS�;a՜0G7q��Ӕ����wt���4s�+�o{nX'�H���uA;����x�F^�!�[�焬%E�3��,8��!r�����u�5�S�˦(�@�3��NZj19l�wWw��Wu���<��͗�f��gZT�n�[�6��ig���Ҭ��m��`N�y��$��M��u~�|�n���7j[�ZqI��LV�r����ո�-�b� �W��#�G]UAJ@d)k%UN�CL��ԭWT誊�s*��\j���NS%s<I�3;�Y5�u�[<U�bB���uF��H<\�ݓ-��m��z۸3'-q�f��K��6�;6�l��'Z�����g�]�x�[nګ�vի�;/Q5�#:����\ývtj{dwOM������{�;W�0���z��.!n�	���g�����E�k�m��^պm^d�ʩ�u�������^��"fy_M�'���m��۠�qq�p#�n-aޏ�@7v
�#8V����f��{�v����K��ܼ�U�W�u<��.���!����ڟh�6�_9M�>n��}^.Ǟ���P�wr�Y��8���ьr����)[�-�f�q�σ�Z�Wdŭ�׀c���������?���E�>L�r3 Ei'7�oc���Tŕ�6�t������c��y A��g�zb��;Qۊ�NٝW����#��$՘[36�8hu�W�z\ѦWx�H��*�qpg����Ѽc>�o�f�-0U����ó���FSh�t�f���.|����u�*V>��+b�o+��e
�ɹ��|�r����_��[a���^f�$�IS�����+Q���9��	4C,��7�95��E���܍�91>�N+�G!�.7R�v�(*0R�Ÿ��}��=s�v��O��fH��;'d���D��*&J_�gģN~������	�t	�ǹvDݛe�N��@�R�1{�2ƨ��6��=��N����x��nW��/(�U�?=�<v.+-��f�ziY�YQw�V��2��c{��cl���%��룐��/��:��RC�+�������
H�M[E;�����2MFZ2H"��"[��PN	_M{���']�#��lu$�Nl�J�Mqx]��І�̨�[+�q�fɓ�����B�^6��&t�������<9�����:�"�[ESAD�!|�9�QM��'ӆ��G�䫷�#!�p�fj��+�j�3�}�~��^�`;��ͨjĔVd���꟮�`���K�+�ZF�1�Ue,Y��J��G L�m8&d�NNd0�'��e�nu��`����^�/Cq���Y݊ |�p�qک���m3?P;��� ������	S�AmQB��F�s�}apb�A����N��1$T�	�{ث~�9�7��\W�]�Y�=ۏEGN"�M�LZ�KZ�iԵUV�Q"6�:7��q)���|o��`_���eo��*��l�w�S�"���"Z�b�&�.X��&��4I���\Tv��k��˛eW�&9��Yb���s�y�����w�Y�j�q�ߊ��(� �)��A�B�i�K?�ק�G��D����:��aws\qЅt(l���k��}��J�p�U�$^D�g}>�QK���k����Ԕ�m�#��W��s�V��&����i>u��޿}�4\#�ɣ�3�S��QO�xx	�XvQ%NWUxL)��_ڶV^C��ss~}� �(^\[�N�O5��]R���{��Fd��g�^�݄j����������'�.y7ms�P��N3�2�7:�y����^c�=��*�۳�^܊���ʙY�^ݹ]�+�k�nŻe�ێ,5x�]��l�Mk�F�.nyx7���k���D��ʣv����v�g`����H&�8a�@ �?�9��,�E�9V�&�c�����������+鑣į���f�%���=cأeۨ�6M���z�Jsڄ)��)��F��@(�ю����^W��
���J�e8�|*���oܦ���Ro���<��.)�vQ�þ��{uRM17�@FLhoz��4Wݗ�3�լ��𞷟e\Yѻ4�p�&:�s�C�풭>��5y�'9�Yz��^��U�E��E�^�-���y�5a)�14�@&�K
��P�E`�꩎�L���Cd�-Z������߸�M>�w�"�v�����'μ�<�T�	P[��
00��k�.5��˜)!�	��L�ZZ���k�d|нef���L��mw:���-t�t��w�tH�S+Ƽ,e��I'��Q�Q)�K	�F�͑ݏ-�!¹3Wi�H���K�xL��t�E\I�s6`a��>��k7�G�z�߁�4��?NF�r�ݫ��9.�ݼ�1�"b��w��Y=I� _��w{n'ϖsY&K)@�Z��u.��C�əY}SX;��8d�Z�h��doK�9P:5sQ�V쭕�^f�5c�ۋ�p<)YOy��RƇ~/2�F#��-n���g�pu��&:�ێ�74�5�,�����������BW�w"���u�]��m������)��/B��k�M����
R��
��g�,�un��k,(X����W��}۰�~y�l����ԫ��:�{*B$��J�&��(`PVC�Qrk�96��H5�T��>/l������{2N+L��������ph�[��n���!��`��'�{�����۳���&�V�˂V�1��5�����r��qg������l���%[�����S�oכ���-�#�^�m�/�*B�S��=&i�G�s0����qi�+���A׭�Qlݵ�vL�;�~ȥ�:��h߰8+!C���h������;�6q9�pʙ^=N�2��Qn^�nIl�
.m���@����¥ڄ����E'Ύq�kз<�m]1��H6x��j��h��Ϋ?LSw�%9H{�}ºG�� R���*t�w]�⠉������b��d�Rc1&:�_�_oS�~��{� �x�!j��1W�O�G��L��z/��CM6���	�G�~c�����,�_3W����g���r�v��L��\�u3^v�ft+\M�U�-N�o�f�ˇD�-�lo����^N��Y��`���@w�}wa,褷\T�d#^wT3<W���~nG5�"˰DF�5P��U�¤ƍc���mz;1Z0����@�e$��(c���3�9��NN�E�\��v�;�jd'li:�o��^�A��?z�F��a����~j��Z=�U��&�ХVX����=�Eu{	k�z�#L�1"�&;q��7?q�Û��j�8�c�.����y7�����a��nNm�k]���PSA����I �e��bd���\��\���o�a�״�_�n�9C��Wz�0xP�������[s��t�������a+�Gq7�����

�/a5K�?+Ǯ��k�A������K���u����_z��}�v�ޣj�,��&ڊϔ��*ƿ}pe�ެ�F���p�H砞�$���x�ť�I+|�u4�<���ߡ���՝��F�=NK�`B��[�;�}��&�fzIF�,��hz�7���6
(��"�X�hm�H�E������w_�E5l�̘� �Y��='�\����ꆑ���L���7};�Sf���,AeQVs9)x�b�g	��e֡����X�i ���q~W�\��P��Sr�t�3���)�P	���`
�t���i��\o�j7�.7�(����ߣ;��P��d;�Ƌ{��˖�ڸ�j�[uY
�T�p�&�I�\�u�05�xkU�۩���(�r/n�A���N@:����i����q㸜�Ҥ��t!Pk{d��Ә�un��f���S-���SSL�	ղ���^ի퉯�d�۹1�ہ���6��'��F�����s�m+������>�Yz�������+MwCq=^��Ze�U�>�_&�+�w�T;�����������<oe��T�����v�3��[g�M�CʱS���$~���ޮ�)�Y���	� d�$	F?��q[�9�vl��
��z`a�����I��פ]�U�0	��%��j^���L�v�3���Cˤ�LD�*��g��9t��7=�yz^��)my��{��.q0���5��=q3&x�o����Z�n�*��(x��˞���Y=. Fד�1|�C|��!t:�u��;ÙQ�iwC.��3M^s�o��"-�]�/�P!x�u.��u)�'������r�UUUUUUUUTV�켵��[uDco5����k����.f��l����q�&��^�Y^v����q�94��ݵ�Nݹv�l7S.����9�<;�c���DAq�0<��b�y6��:�\n��k;���i�.;m 3��iM��~��	����yr�r���xK�b�h9Y����ߕ�Ib,?׉�~�	t*�K�W���ɠr P�L���w��"���U��2{lǣ����tf����d�(�P�خZ����kLx�đ����{:�9ȁ� �J�5�y���s�z��Ot�=UwT����	��ӊ}�F��ѧ�8���o�J�q�@I愧�'I[y�R��U�E8�ו�0}��	�����s��c�V�c��Q��΅���A8\���k��B�9��`���c{y�P~����t��cӣu/5�d6
&�jK�����t���1�N+Z�vݫ&��"8��(e�uf�WNLN�(\�.l5�^�J�̳�u���﯏�U��v�p���ݳ��]c����n��h�����;e@���tj��_wq��J:���0�dy�=_��~�f�f����,ĕ��%�XbG�v��Rj�s��¶$u/����C����lQ^����|�Ǵd��ON�YW+,_%�(�UțhC�7�Ne�԰^'���<�Ɩ���x��ˑ�u��ugW�f�6�<���<��|��a�۳k�E�㣇�J�qCSZ�ݎ�����n��!�iα:(�>�11?����ʢE�4�(s��c�)��.<��:�M�e�r��_�i��pᤓ��0L���q�;F)�\�g��s�5z�߷+�G��CJ��vp{:)�WW��^g+�Gx�b�MF�q=� �*~I��wJf�*\���!|���H��+ZxXr�qo�̌{Q�K�����1C׶v�D�iE��A����%6s��(�M��D^�Q�����$�N&�#$i��u���:P�.��=��EC�ᣲ�g��̵�쬚V@m‎�Y���>��c|�W��~�����<���3�/G�����S>��n0}����쁏����ϔwVAikް�V�̏v�q{i;�����sTB��S���'�jєӹ%K$����r�,V��9�����b�U�SQ�s�6�=��`(�v\;���eu�i�-'׾�^�YZ.�ݽٕ�w'#B����O�j�?r2Jsc�Gv�4B����8{�����������l��#����s���i����p�w�S�\s&���G��Eir3sT������a~B`.��${��w'f^�ils��(B�h�
� �Wx�۸�ت��2���<l���)�#so�߿���� n��+�5,$�w�,8\���eyJ�����e�_f�	=���b2��&�=?z��G��r�|�sߕMeV�����w�M�b�䥷�-�P��GI��K8�{o�m�ؽX껳�7| �Λp�P��	��!G�uv|�:q��;q��K6�G��\L��Q|�`޹����i_P34c��/k����|UO���8�:����y﷣|g<�F���ޥ��Aj��>�o��v������L��]綠(^ۨes�Fb�y�a9���\,���xyn��RUd�9��!��� �O�}o��bC������z睜������s����������]��
���Yn�����7�����̉$��'�"��69��� 0�L2 �&Cm�0�+{7������f����R1�S���Z��5ߴj�5�?^m��m�v��MwR�F7��ӗKn�w���z���"��S��Z�u*]i����q>���&`n�M���ؤ��z�P�iN�*<�pO���S�� %C��gRb/��L!���=�ʃ��������4������%�0i5X�>�co:�8����XAF~@�*H�pF�i}��=����2?o���Z�S���y������`�O��%��~ʜq�=f�Sd��A,��)d�	\&�����[6t_*`��j:U��S�Sv��q�
�����6W��GVE�ӱ~m���L5 ;+���=&��=X��8�@����?����Q%���e8�m��^�tjEU%1v�7`�}�ӲcY����0ɞ������Lu��g���L-e�7(�\J���6\�0�@˂)�$��2�G���*Q��%#՗��O.���Xuh�1�;�����	>��5W�t8$m_o�����Z�'E�dP�ẞ_\�-�2R��j�D��������(��O�b��o{�|7��ry�{a��#�m����/WGF!Y�Ÿ%ZWHI^�n)��tˀ�.����&wZܛ\㽸\�Wp^��v��jg ���7�����wu\��ɍ� ��R�z�����׬G8r���o��1���A��P�h�
mŶ�kH��nu=x��Mj+��A����׀S �W׀#,[�i$�ކ��Ӣ�[�̲;�F��zO��4�*��g�6s�uh�yi{��(٪�D�ǖ�f�V�D6�Y�wz�h�f�η�&�L�t�r����M��A=�ͪ
Z{��i�8u�3�Y��h�%�)�R��A�\�h*�u��eM"[ڛ�%�ŷ'h��n��9�3y�,�$fL���F¡z���c�Q��R����4�j��re�"8cm�cb�A��I������ì�t�.d�wҫ2�+^�ʬ�TA��Or�=��#:��ۜ�n�b��J��f�9h�>�qIѝW`C��\�|� �����1�sq>�J��S������1*���.p_]����KuVtAZɯ�ޗs���ޝ��sx��~�%�.pkt�<3;�W���ُL��MҸVo- �+r<�q�ͭ��)+�%j�;��>�Q^в�v�ө{;h��x�;@$u��e��0��ʒ>B�U���Dؠ;��e���mMkq���h.�z�d�u'�.�����g:�w����s�j�b�I2Hґ�#%�J$ r��N��1&�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUW�󭭺� O���'W<���u�q䢚�ۭj����<�Ů��+�vA��b�4k������J��¹j��j��=Y�=���v�ֶ0���d�Ū�^��ͯlu�lfMd�N�W�V���}֍ΌdCTq\�g���\�nSlv�փfƦݭ'=8���>f��\=����d�<7�.;�.�C��������p���Z.�pZ��׭��s���ݴ����r�a�V���Xn�0�<�\p�\���M&�b�QA��x�U�L�gf{<��[q�A�%�u�K�u's��=k\�s�^=��nݹd�j���5�!���p��U���x׃4�.8u��^�'�n���f^63���k����x5E糽n�Վ�y��<�=�Ka�����n��s]����u�Te#�13�2s]���5�=m1�.{6�ӷ/���.lt��h�qV��S�Lntaۭ5�B���"|���3z�s���vo�2\e=��T)m�����n7�[��2��7O���K�eU�h
������������>�����k�������u,.��<���㇓���A�֛�*����n��-��xËΝ��͢�7n%��c�6�Ӭ��IWYS�Wp�y�Ӡc��{�|�v�y{a��8.�c�v.- ��0���f��1� PW��m�Ǩ�mo��-~_73�/j�N�K{�w�����c�V[#6~0x�v�ؓ$�6Y(���{6a��j���yJ8I�1&;�)��r��=�Ξ�W~d
��0nR���f4[��=���sv�UU.{�fN2�"�?g�v�է�R晻�w)����XQ���'��R!�ս��J	p��Gk��Eצ�l��)�,7v��2G�d��Co����]s�Of�vg����EW���ʽ��|1�geB�0���%r�7=g�7ۮO���Â��]�I(�MFK���|4����ˊ�B�L�يDn����F���&7#tM�v�f�@�}����mK\�=����I��$D�j	b�c�������yR�#�M�?�jbQ�����ȁ��)�)\j���_!P	ܨ:��{�}?a����V�������}0Wvߤ������|=�u�g*�5�ǚ�s	���{�]��4����ާ[һ�3J���Z�9-�v��b��)��m����ֹ��Yu����'!j�IȘ*XA	�I0�Ap��n�̘.d�o=�.�.ڝ-�Nԟ���|����&�ڱӌ�{c��M�����P�	��'Ntv��?&��1��~���5����T��>���zzq{a��(fz�����+=�^�ف��E���80�G��cF����~Q���\`2�(��1Z[P�iោ6tR#�ꭸ�x���a"�F�KO/�"@7 ?���&{��H[ܛо6�c�b��mC''�������r����L����O]lyF�S|�Ti}D���Xz��n����I6p��7����"q{>H�� �x/Z��<9m�tS VIg�#��c���{���ޕf���h�L{لt$�g�x-��n׹Z���lv���$JDB,��B#-8c��5�Od�Ѹ�PI�5Ѕ��O�R������ul�`S�\�#QPtD��8<�ɀ2�+��%c�0I(�T�I�i����T�\߬����l1�F�A1�Y3k��Dak���t/��gq��y���];�m�޹��#2}���H��{�N�h �ׄ�y*��Ni�w�&3Oz���Ä[uլAj�YF��ZVg�9�l5X��J���|8�<U������,N�{X;GN9�f�j�]�|��s5i�}��;�FE#���ܵ�Z�J'y@�Z�ߠz2
��Į�l������
'�(��*Y5�u�����\v�ב�W��r�>Ō/��וA��8T��NtL�ʌ�L0��u��0���}�ŲG�V���l$����m*�5�?3�Q� F�;f_�A�RX8N_W7{�Z��G�l��6�v��ҁ���x���BJO�ixϝIQ��r/�Ftse�4�ɋ��	�В8�q&��K���u�1�n��P�EN4��tU���vzn1��+z*��r=��Q�>�U�>��`6�O�q}�:^�;����2w>6%��l\++�t͹[��N�l�-��􉡞�Og���V�UV�℃����e54�Uz�ы�}���IH��ڥg���^_�����Lo1��sY0�еܔ}���b�0�m�hlz���MȻA��-�R2��kF2:<�	 ��FK��:%��8��?������N��UxhyĈ���W��#��s){��\5�s�����UąRd.gm�ۅjM��U�wd�����.���z��+X(_u�W�i#�M��͈H�A�N�e��7a�,��!�Syq1�R4�I��4�(��s/��E]}�*2��Ez�M����)1^c��-����1[��W�>6�{�ϡ��x�G�,W�"��~���|��Χ��ٱ�+m�חg�5�S0�s])������q}MI�<���7��#��Ǫ���G�0������Oy���{ںpప�U�Ki��)����X����x��~ݽ�@x�gb�u���Z{���Wa�.����A�����q�v�{^�OZ'��G",'n�v��+�r�Ǟ;1=�5+��4"r�wW��ຸ٨,�ɜ���N��s��K,d����+m�l�z�K��*?u�������M�4�e�r�h����oAc��_&G$+�{^��X��N_N=�q�}>{�,���w##��-����'Ě��<Ƒh8`�t�U���D���Q){L�:��3��x�3��r�iۂ�nwt�����
c�n/uE�oD��6�Et� ����_E����e6V�y��('yݥ>���.�<�s��W>�j��:�LU�,���"���P�y�l�u:��D����rI$���������j^fѻT�@�uѹi�uf�ݭ������ �$�q-�������;U�+��㶕d�p��|��|�v:��I\��尅��c�onۚ�\���g���˷O�UL/kOM��]�a��x�q��(�S	@!|��D�8�5��/w��q4��'Q���V�*��H���X�?w��H��3MB�X�m,�=���SL�E�^�5����U�'�م���%>ѸLǲ��xh�4��33]]�ѕy� ��}W���I��w����+A�}Tl16�8��Ľ1����A�����34"���<�G�AC=Ó�b�](k+�������:CR��ߪ��[M�`�羍����;a|@1ȆQ 6aB-�ڀ(�s��F�2�u�����o��
��es3~�ѹwY!oU�����]���S9���8s�r[~PQ��2�l��S��r��0I�������w���
�p��'9��Vu�i\���N<g��Rb�z9Z�E������`�m�]5�5XU�l<2F����B)����1�(�X��s�0�~~Y��K�����ѓP"����"�/+��٨[S��|/��6qz<�ob��,r!e�L��}��S"Z��{���������������*��KA�k[݅u�s���	YG�ls+^�K�m�;1�VH�C����g�Ov�%��[��6h0)�1����:G^�Z�n���o�=��x�V���v�<�]B��!����=��N�i���͞x��	A��L�Tt~e����-~�_�Թ}�c��N�����[%��Z;Y���M���B�zvwгx���]y�RA	X7VD罴��U'^L�{\1C�M����(uh1^�-��-�6vp	�J`Lp�FG�}ˋ!O�m0�%@R"��#���V`�-i?�H�Q4�M�#M�#i=cw�΅c.X8K�>�m8xc�]�S5<xW�Kx�}V}5~��jc���t���,�S��bӎ��\��&�QB����	�*h��!g�!�^���qC�f�g���q��ћ��n�6[��ө$��i�RDT���N۞���NW],��>���t��ҫ�eOv�^�
�@�s���U�x��o���+^	^�;�o��[�~H[9P>w�
OA.��ݩN��<k��u��M^ 0a�4�g�$ƅǽ�X �g�n��9�s�P�؟K*��������p�C�������6�K`�߄�&�+�"��VI����ޙ�)�pT/�d�#��U���D����������No#��w�]�� -��@��Y\u���K����i�eNԇ�ӜO#D��H���}�R�.�/-N?����*7MR��Ehx��q �L2�c�6�9�vr��!/�7�$yY[wY���&�1Jkݳk�Gۙ;qf�P�߃uw� }�^�8�ߤ��G���y��|Wzql{��+f�t���V�$FfT�i納*�/v�<#�r��e��w��>��}�_�ʼ����Ѹuۍ���k�[).�ʛb����+������q���}���o2T�13)h=�֣�!v�E�:����cŔ8{�aE.5�^Τ�e�Q�q�9k��;�qUA>�*����8�W�#;�<;^�fg��;+����Q��o�b	��b�������P2a{�t�R�H����UQ���r7<T=�w� xuG<������]J0�_�5ó���yM��\�~����ÿJp�M��$NneC|������c��
EL"He&��A�∔���[�M��9�_V�t�M"�.����5\��U�yRd���i��Q��͛�c�:���frxJӫ�G�$���p]B��2�险Ь\b���4��K:f��U"�ES'��$�n7kV�I��P�d�1�4-���s��u���vruV��8��=�i�v�|��B�2 �㛅35^��(�MV�K��W'�V8`�le8,�H��Oɑ~�׷鲗0,��q��2�{F��xщ�t6Gcq��Y�ݿc��W{ͽI��
�cV8�g�{�� ���	��~nE(;Cxňܪ��%���,��w�x��;���B:�b^��ܛQ6vzV�,�-f��2�clP���48w��LQͤv�{~��0罕Tdg�:w4��^���;�fj�}>�����'��۴����n3$.�//@��{��@�����^��U��l$�CA�a�
M�?�Q7���B嵿! ի#�l��3�j���$���U�a\1�K��_S����^m^�޹'kAP�1�j1w�{�*G2L�W:ۍ���K�#�׳}�Tnh��58�E��2g{Oln�+~���w5;n����;��yG)ɌK�j�����Բ�0�� ����\����ά�$���ꫵ��H^��h�/�f��^ʈh }����򪪪���������@��7'm�_�s�\q\q��������=�Bw'>�n����N�x�
�ٕNw=m7[mͳ؅�m�ni�f��]�뭬�s�-���vn�x�hۂ�~����Tg ,)���@-�swb ���� ��e�YQ�~y'�O���^�(���d�qU�"]���I�hT	���U�D8��Y��#��Y_<(7�)����(��kq�vCW�ar�Dr��7>ʿVt�\:��.ª�����~q�u��V�vރ�oX;u3�q���:�Ȣ�*�A��F��4�B}I�w�[��Ǐ���;7n[7�42nU��s$�pw�������a�^(��5�z�nk�P�H��#�!�?���8��d�	l0� (2��?��cḼ~YQ��@im,Q���^�g�(���o�5�#����͊���{4Z$(2�]]|<�
*��nhp�&�֓>�(+M/��^��F������S1H��LE���{{F�_��*c��˟�;�byk��Ͽ��O]����rQ��
zu�۔3u�����S�̍��u���N�im�tG<ŕ�����;����m�l�|����0bP���s׽K��	&�'c3�\�i�^b
&���_x�+��\�l�!Q����k���L?/9VF����dVzr}�pږ�$]�9�5@YB@�;��W,^��U��H[A)�B#w`�m����w&�y�����Um���mt����x1w���c]������X�q[��w��'�h+�` �@6+#�'	��r�dB������
D[��F�<xV���Fn�S��n��_�/pw��wY�Xg^Um�@���2}f��ݪu���X�^�'r2J��)�eAT�zN�8}4��sڼ��"����-QSs5��9�[-�eU�8d����אstA��0$�j~I��	�a��pa'��l��Tz;S�l��0Ǣ��ky���)�(p�?;��gU�qݱ_�y1C��{�o�1Z]�"�(�)�m����T��x�N|y6�U_j�be}=w��ɚ�]�Q�F����MOz��(�m�CX؊5t������I$"#-�I��B����7;0�N��U���mva*Q�⯂�2�A��=}���, �:M�x��E���d�N���9Yތ��t^eۛ-��(��_f�~�\�;�8��H�1����gJ�EzOw})TfkW�x�y2���O3���K��j��C�|�}V�gU}{/��t����h�}/�w�F�0�9Y�}St��8#�.�h=�e�^���ݖGJ���u�xH��Fma���ZP�h�K��K~�-mnlT�.V�Z�j�o�t���e�Gh��g�,y܅t�!�_u7u����F�x�YyZ��C�}F�h��D��e�`q�
_:*�I�����]M\]C���M@p����*g>��ū�+OC�,�����=��D%ݒ,����G�jWϖ�V����s��+wF��ц��Ȧ�rF�3,n�% ��B�}H.�<�G���p���z9Ҭ�N��d枻�֛��et6���:������V���-�EKܪ�t��^�Y�2�#�U��gumWx���S�S��$��ޝ��zZ��͛$�W<z�RZ`c]]^QHk3'*��;b����99OuVt��eI1�I���8��Y�H�;j�	[|;9�}}g;�ɢr�ro�z��Y�U�]��;ܱ[es��K������da�I�0����/�y;�d`��J�\Zxa�賑��֎��t�<���2�L/o��lݼ"����K9�A�
[�e啒ce*��u+!} �9Ty���z��ں`G.�ΛaH��ùF�,:6�^i�	!�W[#��*pՎЙ�yLmvf�U��
�C��#���3��fZ-�Bg���ڬt��da#8eXY1�u�Ol�Z��p<O>/fʳo��R�m_4F����<Up�(��W���UJ�<Ӷ�Q�-��0d�gWi�Q���&�Nwd���F�^�%���5/�ՃWi�6�Rv�#v6䮮˛�ѷ��i�:�oj�f�1�q3��ȕ�tlӷ� Ks�[�;��x밶Q����Q���3�õȚ�6�C�]�;cBt��o"��e�� nnt<�tcQm��܏c1���`�^3=��mJy��Й�v�2x���h�;s�Ov�yN�bŜn�"��Ru��zWc���{�Lv�ŋiNz��l��ɹ�\c�r�;v9&�۷i�Z���uՐ�����k <���GES���x]v�jl��\�7v
�z91��QSE�3m<�K�ͷ���*��m޴9R�W�u��z�5��m�*��:ݛC�����j?7�;fk׃�$��إkc	�EX�li�$�}���cqP��O���
d2�оs+�y�lKr����L�X�a�K�af6�+;���T{~��WV\j iPՇ0�:����k���g=��R�z���׵%���h���SP
݋{ X�0߷=u?*�(���S�4����Uۖ!f�A�����0'z������z���J���tKC����`����g\k�ԢPV��"����6��g�IWm<aN^,�2�0�(�]s���R�[4s�ZhZA�8��r7�w���9�\'אh�A�dq��zH�y����ng�19�g���
�F��7��:'U&�k��g�yE]z�6����p|����y�3� 	�;����i\�qxb�&Ul�}����JZ%��F��U��5g=�y]�J!����.4A�EwL�X{G.٨)�劎�x��b�ώ�BI���h���l��^�_o����{�௵F1ID���L�$d�܈������]J�'��w�������e�]���KZc��4P���=c�X��	ŝ��9#�k8�lZ���GY�*��Y�ԯn!�J˹Mm�e��hf�v�s��u?24�us�ӗPm��(�wH��~(S0L";#8Ĉ��6_PF�^F�g�g˭ �mVi�&E�[wi~�r�J���Z��z�OI1���e��T ���:�zhS��@/l��'� m=�n4On�\W�h-�i"[���a�~�8�P�
%���Ϩx��uL��_T�~hFW&e�����}y����;"����ޭ�i�iFBe��44�e���G�3ͭ�x�ʳ�&\��(kx�9�n�X�+L�����3�l�Yɹ���Wtq�۱͢��J�A#� ��5��sb���wnB�8��7O�dg�0o{�BQa�r�y�ȟ,�w�j��dμ��E������>��\���o��V�kgZ�tZ2����]����X�O���VTa��9�S.֓������W�b��*G��Ӱ�da9�E�E>�W�>�_Ƥi��a�\:�
n���6��%µ��l��u���o |�R�>�t%� F��s*���D�༕g=G+8byguc��#~��`�`��Y��+�Vh�r��2�u`R�7x9���[��,��WpOw.B؏z�o]���{f����������p���X�p;lQ��@�nmen�c��Cv+v}TmI.��]��y�6+�g[��@�u�i�ی�n��]�kp`�KѺ��[�T�c��~;�4k�u�&;p�'Aչ4�KUM:�t�c�c!�\�7m��ތ�.z�(�]�D@�?~����19��A��)�D���F`u�aTP6e:ע-u1�Z	.�ع�T�鈚�p��h�e��ʱ�{s�LR����>*��Q�ߍ(T������<�Eur���*��Gf?���0l���X�ʸ8b��fύ�����e�p��ǔ_CB6G��1���*�s��9'g���%����l]�n��#�:�TTx���F�!&��.A��Z2�0����'P���?����|�����q��5�s����118Y�V�yMީA?A*�޺���
H�[���l̽��%���},m��u�����Ga&P�񡣅Ϩ�(��l�Q�f��\���$������q�gN;�9�w7���>��~��㜏:E���5U��g�����u�y|n�v@5��󽸼�T/�n�>��&$)��nH�]�Kvl�eҎ��ޢ��o�g��)W�W3�A�<5�p�4��}��a����Kd/��]~~!�a!_ ���y�9Jvu�h��1��?���=����w
f&:�JV�t�dmX��ۜ��ǘZ��QZ(>�]�t�q�o�3w��߭�����/gi���u]s�����y��K�g�[=�mv�^������Wg����cX��9��wc0񧋫l!.�7�wF� ���� j$[�������l�� p��C#5�k�p��Ʉ��W��a?u_H��i����,��'��Pl��:��^4!�tI�X=�Mn{0�V>d��W�}.��{���OPe��КM�Rl"�El%�cw��K��������t/գ��1gk�F���ޡ���1K�xr|'6߲�>
v�J E����l�=����W�ѩ��.!V��BNJ(6�
.4l���J6x��pk<�^D��8g#�W/�d�:M�zT�x|�s��Q}���X`���^���Ty~M�<�A'�D��NH�a)4W�˽*c�Z��sml�C�Ԙ�����������!�+Fd�b��h��,2�½=iў��Do�j69�H�זM���6�{��=y��P.� ������zR5�q�k� c��G`�W۵sxqX�z�Ӏ�����a��p����Aq9wإ���l��7ۇ��m��QEu���ٔ�j��M'�+��f����Z��82?̝����ӱ"���9>��m��:"�N;����Qsn��������^��&�@����)��;W�Q`=��z�[���$�JD��,H�\Q���Ch�$�ّH�R0�,&��Qe��ޓ�"v;z��ɑۓ�Zs2&e�wt�>it��
�>���ZU��Qſ4͘�ѱ��fWc��]+�q͆�F#W�z�X��{0����>�T3�B�y��`=�}G���s�פ�aJ�|���]�����S��f�,7��6�����@Y��q�#� i�͎����.{<��-r̃���_����NE���Y�c`:����3H8}��r��u�8Ƌ�.1o'[��i�S^�N_z�ŝA��������s�2}ީ˨�w"Z:��cƫ�ƻ�!`��M.���L�tųD�7��Qlw�sœI�HGބmԪd�� �˨�B���<n�a`x��{�_��£�r5��c�W�i5cW�=����.+6�#F�@�--��X��$E��`���*?bQt���_�B�O! ���)\0I-�l�Ko=���08�t�>�͖6�VT���1UX=RPk�4z�n]�wo�;�S3B��u��-D��-)gm��ҝG�i�^�3���6��Z�w������G7��un�*�t�/κ�o���i5�|��K�S�u#��3�Q���ݘ�2fl���|�N�F���*�!f4{�y������F}���֟+��>�$V�-ܐD�?�@�3��O>��g����·�L@�C�@���w�7��sR���~UDp���ˮ�]�y�]�^�^��Mb�7�>�U�坩����]���3q�3���qh�D�@*c��Kي4H��˝�����a�ۑ�0����u�.gha�X2�ź�JA�6��)^+�_����V9C~�2��A�,Tj�#M���zO������Ǵƿ[^�p�k���E�l:0��O��!RI}��0�US�]�aȜj	,L�&����(1{ݽ<�.�B�ےB��;O�����>6�3HU�����xn�П���Kp�w�2
*%fVy �m��L���K<�lu�T߶צ&6c�>K�9�U�_O�-�w��^�i$��~_i�Y�Ǒݧ&��^��%7���%Y��f���q)��)Sm՞�ӻ���Hku�f�X�=-u��'҅'8��#��;B�`�5UUUUUUUUV���	�N׻]��m�<��x���8i��u�mָ��u��|7x�l]Ռ���:�|>Ų�sq��uS���8��]C9�`�V�WJ�^CY�<��۶���'9�*�s���F�67:98I�M�m6��j���G���Ԋ 0���4�L�H8d�<�v�J������|��샰Au^b7f=2#�t�,D�?�4{�ƭ�8 �G�hyS���|�W�0q[��2�$L4��u]|�̟E_�v��;���-�g�8���I@�>}u�A�����	P�S(�p�Q����D,����x��9#��m��ڟ]Dp�}s~+w�pvC,�����r�J2�oͦ�F%�i|�;Vo���8�M�p�A���� ��1ީ�xF�p��3;�OR�(�Z�[�&i�S�'C�g��1Ա��0���mܓvY	 _�����R#����� �ռ�1B��}��\=}S�o0�_gu�^���q���A�'�{X�P69k���m	��J�I� X0��bp�8n0�9��v8��.kG�}N��r��Y<�7��r��OZ��;מ�OH�W\�0��VS���z� +�aP�ٯT��`�n8ݳ=���Sm�X[7ǑH��x<���.�i���	1,h,!�W���X�O��T�A��k���8�]rR���=�_l�}$A$F�BF��P��Ӟ����\J;sz�q&���Ѻ�l���B�@u�\mm\�;9[v��n�&�$�ext����\��
f9#dėP��㴧�\��+��\��y͉�J(�d�&�}tn���lv]�͇N%E=��������֋���Ϣ�9
7�z��Q�U��[mV��-v�9r���P��=x3���.q��f�u��
L.f�7ϫ_�'����q�p��m��o�b�~~�4`UY^���u������̫�'w#O[�	�-T�w��llt
4$�0�T\���a���<��gzd���Jm��5f�aMQ�>ѣ�������4㛆����3���ܿͷL��m��$�����PF��!�Τ��l�����Sh�i"�QY_�����'ު�n�H��`�i�yQ�˙�Q���˽��AI�)��D�wcӶ &�D2=�*����[��gS�9�ץ�'>�鎷M�Xٛ������Ia9��S�F$��X�'���f�(*a�{�+k�z�����`SK��эe�8�W-��4�����-��v-z�������c'�GH���J��^�R�f,ʕqvQu�wڭ�3���GNxʜۚ�D���xX�@o&4
)��9�wI"�0Xk��/#߼Yl�g�{�{�&�xS�`��tC�￼q^ڥ6���cl�Sp�����Os=��3Ң�R�C�OT�'֋��ӹ5.�(*p!��/1
�Ǫw�@���\8E�U�{΀^�G�n
�z;��$�SW<��B��s���4&lgD�ʀ<��YT���^�+�*m�\B��E�u��57nх�J-4�e� B�o׏�z�f̱�\dz$N��y�R;��K�ۨ��X+f��9/���GC]
���3F�v	�D��>@�����e��~��������A���R�r�41�op��]vLO���U�iF��^
�ڙϞL��	?��$~���tL��U,�Լ`L��d���r�]ѓ��r�s[]x7��e֗��'|���A$���&[惫4�^s�o�ֹ
���"��ז��J8b���8&�W[u�ʟI�&����妫em^��Z������FU�kﯪ�y�
�qb���(�nu�|��QwǤ����"���u�ͮ����Z���[�A͂�=���U,�'�ܪʪ�i��;E_�.ǽW��C¬}ۼ�L�*D�-��-�hY%���k��1]Or4��!+P q�8!B[�3N$����ug�&� �>)9�OZ�B&׺����.2r\�0�j"���L�qt��M���ۣhT[D�bqT�

B=�yl��wu|�Xߖ��Z��A3����>�<�SE���Bా?�|zv��*Ɖ#��o�cD(~���7��)�:A9*N�n�É��/ũ�1�{j`o����F3u}��o��/���7���՞��S��h�ϲ���e��2)N�7�dt�f��I!�NV I�#��[<W`�Ȓ�p�#A�E�V�+�Y�����t����������-�]ϛ�t���{z}��;�s���_�ŝR�߯Q�j	{^�\���w��Ѿ��/�n^�7$E�Z�=�p�+�UR_���9ɝ��W/,"ǃ�E��"deK��8I�kJ���L�\'�����AW�E�����V��?XE��hZ_|��x��
" ִBEdTBDET���
�EB(�2 ��T���"�<�L
�S+R��QUd Dp�:2=���t�����O�����?��!=z�ח��� ������W��B �
�Nc��:�4���jr��A_W�e��WRzt>�i���N'������"�#]�T@N-rn�|@Y]�!_��9lð�r9���{zPAZjV��s����$٫�N���xs����AV�#fS��\TA]� ����c� TQZMIyA[��J3
ׅJ��r|y���(p2
�M]��Au0N���5��4�9��7��Z_AY���3{PAZ�X�n�|��D��M:�-�
l?>�χ;�����``dq�hgт ���&�3�gq�Yӭ���g㡐��+É�aǝ�2�E���(���/��d�Me��)$
��f�A@��̟\��>, � @�2�4 4   
  A� @ T  �( 
P (   
�H�J���UJ%
�"*�
R�H$) �%QUUD	IH���HP�)AJT�R���$�R�(�!%xw�ʗ3RB<rU[����=I(u�4YmK��)�V�o[���n����u�I*ց��^��޷R�؅G{r���O^�{�EB������:I$   ��*��JU
A%T��P�ր  na��4P�{�QK͂�a�z������![�S��{���)[�uR���n���Nt���R
��*�f�0iQ]�w��4  *@��^a�tn=Ur{ە"���J$#&TI��c�P�U;�ԕR�O�Ҍ�{I݃�)#�
/mO{r��Q<��ޥ���"�@(c�TD*
*TE��SݸE*;��@�E��Ru(��n��"��  =�� � :�� K�����F@�w1�@ 22!T P
� 8�ª�� D+�  Hʀ�v � �� 8�(�Ω�� �F�  dr ��@b ��	]��u�� � �7�DR�
�HHI,{c�v9 
� {�s�I�$ ��� �@�m@P�`:�z$��  �Y� P���P�i��(A@� �t:{� :HݎJP&� {�C݀=�UE��� +� h=�� �a�@P�� ��/{�� J�  ��⒩dP��P�w` ^ �����{� p�K���!9  c� ����� p�y.� ��B��P�c� (����y$���� K{��s1��B�s g@݀ �  2G��8� �o@P��mJx]�  .@  ��*B��$DBT�sb���U���xڊ���EC�R-k��$syॻ�[o{�
 ��#�ނy�@{�E �� �X�K����� 4.�� {�� M�r`��	���<� ��$����@�`!�&�?L��dj�1 ��R��� =
)J�`���O��O꿩���qSmT��2J�P�$����i\�9�OH����af��?���K3f5����K3fLY�1bY���fbY��3��3�ř��31,�Y�ff,ŉfb� ����W�����"(2Ɂ��r�LN����N�)G����j�u�)|��Ѹ���]_Ҡvhc�4wd�d��iF2]�i[�n�.�Ѡ3���.ՍOi��ț��iu	fo��ep�w���yF�����\2k�4��al���$,�1P��I$��Zp 6P�q�� ��/]��j=�jX��,� t\9W���ݔ������UT~�ݵ�y"���9Y�� I���
��cg�>&�ȷ
a;��ŕ�FE
�J�wZ$�&X�q@,�Cn�z]^�m����A�soK2h�m�ƁR�ذ�
,��1@J�.ـ��v1�mZ˷zI�Z��Q�bΔ�Q!]��"��/nLҷ殝�����͠�*�f�/6����E+4iw���M+��\j���kWh;�F#�oF, 	��%Z��K-_� )V���j��5`��T���/Fl��^P�K���b
�b^�geg�H��Y��pJ5KR[*����'wsa�J3M[�x30LUBeR��p+%R͹���fЎ���5%j�A�Cd�׵vҿ�ХBV�TpSZ��2��v����[�"� WW�0�(-�ӛ�K͕t���m�Z�gX�T���_��[pe�ub%��,H��6Eca��3 P��{l����`[�=9�e�>Az�ƘF���$7��$�D�2fd�M[��ܡ0�hn���*�=�� �\2�T�b(Q;wX���2�'/����v�V��X�&ˣ�l�F��&0dcR��P5�Yv�ʃ(���9�P2�V!�������6������5E���.��W$�������0���6��M�G	F튶�jʗ�����"� �E*k�cҪ�L:�a5�̩Up�� ��l�F�֪�]Z�����ѷ*7�mlͼ`��[���*��vn�[Ub�P�vY�{m��������AwZ�óP�I]X�����wo|���jm�R��guڵ4�aׄ^��f���u�!�Uh�N�+�������!������О�橡UP�fQ\	��wt����S&���ѕ��і���K��J3Q.]H/3Z�͋]M`(�i�R "h
[n���Vx�.h"��2ޛ�-nä�L±ˍ1[&ȯ`7�n�"Ƚ����l�{�N��{p�蝚��ǫaݺ�+��W�駂�&5C��Q��sjJ�(J��t�F ǅ�n���M]������%�[�LZ�%�7�l3�P�����G�z���TҖ(�94��lY���9�f�nmM�.Z��t���6�0؞f��3�r��
��oN0�؁�[�3�mz��ʛ��ݭ֋t.��U�*�ɘee����ۺ�n]A#�+�,ֺ8�l
�Nh�A�5eR5�����nn��� 6�f7���9��%��V0��>��o��e4�H�l��z�z��7�)[R��L:�۠-�!T�2�K�$�ˇ)����3�wM.oS1|����϶kﮅU�v��T�}��I�V�=�s�"�k���9X�4��D��cx n#�q2]ĝ�/%�	I�ݚ�OcA���Ke+�V��ܺWAd�i-����\�I����&]A��Ƙ��a8ѷ���)����;������#la�^Y�t�Y4�,w�җ� Vj�-����pc���Rd�ۛ���;�Rz��ikS�MVU�� l�:e���P�wl��)�5|).�b$�ѐ�5�l0�����t�g3F�5� ߤ�Z�զ�VT)�c
͒V�p���֭ͣa+�fޣ�
=jp����~��c��;��PXʭ9m�e��B�U�[[x���n� �X�G��.8V���uѫ�C]ݚV^4sYK��֦�+3i�Rɴơk챚��@\��P�蘓�������j�VV�
�	/j �)LR��O` dbl�O5�̢��Hq�7h���v�RSw�f9�*���e����	���<��1��̕�!��@(��Nf�ʙ���8�U ��r�1�[t/V�T�g�,찙J!����t��o:؆��莌�`K�����5����]��v�g\���%^�A�ʗ��"�%�(�sv��e`Y�uU�r�7�Zh���n2�r��lx�r�N��/.��mL�!D�6�
d�D�E��X�,�Z�!+w5]'��kL���)������*�Fp3)���s-����\�W���v�U%�w.�/�gI�2K9�o.���Jպ.��Y���92:zufV�D?\!� �/)�M1s.P/�&�v�iJT+�g!V.�Ÿ�i��2M�sIWxՊ�i�{sU :J�1Q�V���G�@���Wi�u���x�ԫk~$X�b��q��=�1��q6;�vՌ/5�,

b�� ��7��p:5ŀ	D�u/2����U��vCwF��X2SS�.TT��*]Jr�����V�Yc�9�����4�n���2�I2���SQ��r�e�u�a��oF�к;{{h�x �ܵ���Mц(
�WALU&m�mI�����G:��tY��u
���UJ���(��.���U'4(>�dd�!�c3�.�jY�z!
4hD�)1n�V����
�nXaB�Ժ���t#X�<ݱ&I��E�kPQEk5��`:d�E^Y���	��ݻ��-�`�3V�b^M��Y^�7�e�M�Eߎ��,�3%-��m�en�W	��6K�m�����$�	RB #���[����Z�� Au����V��L���Y��3R�Xx��fZ8���Mʏw:�S������a��-l��6]�|�W%�B�ܚ�e��36��e��6ֹ�bm�z��Z֤6>R�K�;/5��	Q)n��� �
��܏4��NVT�xݫ����e����J�Y����]�Qf)a���L[%�&�"���_��c�=V�j�z���6�#�� l�"�Q�0��]��^��d�ɍ�65���ә����f�1މ����+f<;�)��T�n������X�d��BZY�w�<���4.^}�*{d:&ʳ��|��bw.d#~�V0�a��En���3V���ͬ�=eY��os�*b6K[W%[�d�m� *�h�hM�C�c隢11�{[��� :���j�EV�w
����h���X�+7t�5�IpM@i�)4���{gqTG6��$�P�����x����S����֊t�֝oD׎;yS2�ne
Ȇ�h�*gȅ�b�g",�b�ػn��r*�Z7�<��ɳ���.@��-�#r��dR�s5CwJ�2	q`�i.�5�l��������f<����4���d�4f���زm̽�3+V�WXB�j�u��]1�U����+(5l�ܩ��V�&�4!�
S�e��r�A�l��aeQ�P��,	1�wjb9���7jZ"�)*�E�L/.T��	iJ��f����5��t�wz@nIvĘ��@�U�kq�M}T��*�}�4�o�d�bH��v�/���5:�ĵн���~��js5ܥ*�JR�N�m�$hQi���i����5��s1��E+�e��.ΘJ0)��IyVv���wB���eb�b����h����Geʧ�+v�٦�ۻ"��y���Q��ڄ��M{#dZ�(r��Q�>�e�8�@ە��w{��^�9Pm`�H(+d	�F򉧘3r��kNaD�%��XۻJS$�Y���,Q����e�VFn[�N�6�jZf���
�w%;V��&���6�tE�ѧ'ښ*�P�=[��Y��zf��՛#'ڦj�K���'$����( �3-�"�[�I���Aaɫ`�-bof���� f��#����X����H��0��XV*�6V�N�j��摧1 t��p*n�U��-��%�6��S�Fé%e	��p���'oF�2�b��lZ�ǖmf����������#&k
�(�2��XOr\�-"��ӗd��(D��t�١v�:��l��X���$�����W�+���N�Ib�ۇ>��%��p֩�(�X(۩QY�-YRQ�n��vʻ_ Vk�t�����2`sn��Th�WD��S�������K�܅1K�d:J�������w��1�;�R8[ܡV\�W�b���j=E(JZt���SA���!��N���.�;h'�]�3�3%ˣF�U< �J��[��m�2n��u{v	LK�
�ĭL75�[@�u��2�9�0��5��v�dSt 4=�T��-,�Lq��h�[�fP��c׋
�.�l��PU(@��bk�~��n���1u�#����J��z�h[��ok%�I�֯^Mɑ�	��7u��PY4uˬ*�J�D��*mʎd�0�t֊�F	��/2��m�o5�jm=A�eř�Q��ő�
s(�6���eLA�p�ك0[��.�h�9ufV�3����M�Z�Ll|֝�m^P�4^R�m+��M ���kP�n�0�_����ˊ���6�[F�' ��b[�KR]X��^�����`unQx&���`����7�\���l��	P;��-�	�.�w�vo0 +[�We��de��6��꛹�y.���O]fڔ��6�I�EO��iQ���.�V���kkN�����ԣN�5al�������FVA�h�%lp7�XJPT������l�n;�d[4
HK��3~4�aP�I�vT�^T�*"[ �pf^V&���0e��)f�ó�,3��T�B�jCi,�&v-��k K[���w�EL�TL�̕�mG=p�&h�c�ܣ���vp� {7�u=46�0�ɚ����M��f������m_�1S�%�S+u��&[���:����A[7�	y�*h7��M�-:%ʘ
05�N�~�H1+,����+bWA���g�eg���P��8~��S"3skH�5���Q[�Vⱉ0f�x2nۗ4�B� �ݸ]KHm1#��hꎍ��e-�p���Ma�nC`^�P�?4�\[�-O����ȣ�������2Zn̈́�xU�ӛ��8-�ژ�b�aT�M�`���6�m�T���5Q�J�f�X�:4��5V�@|�Y)�����Lj�Τ0�Xe�tL�X�h��1ҵR�^|kQ	���
�'�benm�B^R_&v�+�e����[����s��3~"���jr�������m�ʁ��Iv˻�E+�]�m��Pق��^�)I���3EY��kV�� �qXT�): ��Y��mA�	���ۥ��V���"�.IN\��>L�.�H�%V�ƫ�X>�Z��d�i��n=w�r��6Z�1�P�el��-
۽[&P�*�����.�
�I��aH@��(����+�YOcݹ��M��-�
� ���h;{0|�虙�}�q���G����h�/���Φ�ݓs��J�sw��j6rc��vP�4�^��x�
�9zn�.r�f�y)��f$�u)��ֵ��5&���5"p��PC60��ub�k�%-]ɨS�����^l�~�#A��WV�"�#	�Zo#�u���{��j�� ���ߑR�,��@��7��.c�6��5�VV��*���5���gUI�����ᚔ�/jԠ����C�h&���Z3v�d�W��Z�v�E��-;�e����TT����5�ͨ,]n�=�Vk�lLY�Ӭ���!Ÿ�J�KӀj��|eџ�a���o۟!�ˤ�q�oveV�hTf]X��I��˹Q�U1�{tF<Uw�{���6�5%�Ad�N�Tw`�Ϟ�.�{*KhM���iiW���.@�[���u��Zsw7M(7c�n�� �oU����F�cXE��Cމ�N�=���.�]K��M��nj�>MܛK�%�.�T0)�EӸnb�l7�͚t]3��c70҆f�sla�+Qm�V�[�T�T�#ʃH�.�*�z&��\xJ��O���<!�K�-Q-!sS��:;���J�-h�P����BR�9[2��Qk�ɩô!��w5��50o7�~�a2�Yy%��V�r,�-� *T���8>�����X��Y�P&�mM��e�İ�-G(֢��3�YK/�$޵8�'^�1�6�5���Y5M�Kk��Wt�|���2�h^�k���q�(chj���J`�;݋�]�*���a�����S׳*��+-Y�];�%yYxm3L[�4�Xs?<�z,dJ�3w ��3V�p-�f��K�����0�V�dͭ9��M0֧� r�f`4+Xj���u(���L,��A�x�7V�x䩎�;��T�����F\ͻ�Hͤ� ��ї����O�����6�D�٫�x��0m��nj���#��j�Y6�Ϋ��9Rl��x�ܸ/MG�x�`���f�"��[���B�ن���A�d��m��SVj�ЍԳJ�
s	r�T�v���i�VW�v���Y�!��B����/q��+v�6K�sQb�k�E�6�p˽0iPڙO6fVTd�6�Β-�� �S˗F�Y{I�iSH1�r:kZ�����M�F��F[Ϥ�n�m����U*u�h̤�X+v�N^�5���Yj�T��UIiW�kak������f���Bf��e��Y��*����7mI`�H�ws&R�s��YtY,<KT����`Hc���Ū�d-���+F��A��ou�1Tܗ��bP̥�T`[fH.ܩ��7�5��2��v�v���j+$�[�0��n�:2��b��^(uլU/E�HVN��˭4lCeC�Y�(�B�`�j����UUUAN���MPUUU*�UUUUTCń�U*�UUK���eX\�vն�u������������kl�UTj���UUU�����ZU�V���C�5UUUUUUJ�]A*ԫT���UU\T�N���U�
����Aj���m��R�b�79�s�<h3�j��zx(7i�d#u7�\�����46�U�yN��m�:�ö��E�����v����<�*v���1Y��:�X��4=�]����x͉W���! Xz۱\6:�q���y;XL���5���\��7�d�W5��������aw
]��K:���M{<BT�=j\� X�
u��Sb�b�E�)�9�e��vK�����k��@a�e�\S�0��d�9g�䄻��[���]�;-f�Xxe�cn����R8n#�m�.yz��=�=yygH�l��8�&ݎ�1G$j1��ۑ�-1���j�m�&�:.Ûx����4�5�Ss�K�%xp�4��6:�����@�]�P8�9�^����M��yz:���]/5�^4`]�<�x�����^�p'q9�N��a�<�{=r'���vݣ�Ӻw:�ݶ7W-7(�޶�}�n^����9���|���Ɨ�\��'�@f�T�Q��7;m�c^n���Vٹwb����l�e88G���/���]���<:�vށۑ��yN{8Źz�>�Qv�yx����g��n$NN����;9Øe�x�G^�n��8�:�y����v�+Z]�%�،D�u������E\V7msƎ�oOFbmJ�F�U�����ǵU0ێ���k��z�9���p�x�]m�Ɏ��af��Q-��%���=�ve�۴q��S֯JK'.ݲ�<lC�7�xb�:��J\]sXt�sG��uu�q�eyݎ.v��[�u���#F�Ɏ�P�nܺ���#��<1s��t��s'n.u�^:�I������vK[���y��6�1�e�4�N2�%x�O8"�=�n�5�մ�����9��s[�%�<t�����jȜbw���<o\��7��qe75C��n.9��O]��0�zw-�����䣣�]u�ћqܯ/<���鍇P�deS7u�#�۞j󻤟D��.��H�u��y��\�K�Mt<]R�=�Rn4�=�.N�O6�Y�edY�k��O\�ֽc��9��Y(�nxۛ(�W��=Q��xx h5]$=��n[�2�ur���[��Eq�>g]�.�礽t�înx�����p�uF)ӱGl�K���2�dKs�����y���N�n�':�Du�u�2N؏]j���ަ�b���g�p�ݣ�s��'�X�Gi�Ł�X�i��ԍ:�ĸ9"ϻ;ц��U�	k��<d{X�6x^j5��k��������t���-·�����t�by���wnƮ�oM�nc&�]̀K�����%��bwC׹�8�l�k-m�c6�֩�� ��F�c��Z؟:��T�<Nq�A�Pn���۷Q��#�'��,�[n�'Y�G��z����΄�ɇ����v〭9��������0<��÷i�	��Dsj��i�uڧ���ܮ��ܮ�����F��<WV{=v_a+�;:+��^���D�=��D���i��cS�rq�t\	ksy�C=��8�̊��sUN�h^�m��B�ֱ�.m�Ӝ=u�ԝ�p�n�e�.���+�������I뤫�6�[�8����3��ݜ��mj�>�H�+n��"^z�r�K]'W�
�񵫞c��:zF�C�"�S��I7�ݲv��I�ڗ\��x�����s�g�
-��b�v�qzmPή�g�]�GU�V�W���m3�s���u���Qf3v!�(���Z�'Iե�����u%M��ũm K�w�`�M!�V��n9��N���ꀇ��q��&��k�5��[��#�]��f��v��r�9���;=2�u�\I����l����L�i�lr(�O��8�wT�&j���<vx�e�t�;�����ܺ���n�.�;=N��v���v�8��������Ŝ�W�V�{E�`��. �2���ηWW�+�F����.�v�c����vp�KONV��nƷWX;V�'�M�T2y�����U6#d����@�̽B�v�ct�\WO:��
�Y��2�k!�8;���n�i1�θ8���y�HJd캥;`�Q��2F�>�(��c�o�bҹ�=�VP�N�=�rg��c�z����wn�(݊q�'�uIԒ競Od�]U��n�ݨ�d�qp��G5n����Nպ�ΜW>�صa���b�y�1�]a3��4"���T[�G�t��=��sw�q�v#hu8��\h�-��ip81H���e�p��H\�\)�^�P�5��	���ī���e�J��ك>�нE�[��v��i{+݉02I�8ll.ʭKQP�^�'���g�jݎ�ܻc��;�CLZ�O	u��p)��<�6mpBv�q/E��7�ihN�\�q7*��qp�*���7+v�/\��M�⻆�v"&��J,v9���թ]o;uTfF �9�9���c����W���Y��ƹS�z�ޭ�r�Gp�ؓ�˱��%�QqD��[r�P��-�/���B�r�ק�)�x5�r�rOg�[�&�z�]����jkZR0��9�ЙW������B�N-�$&�'qnyP��)�ќsZ�c�<9��C��G�ڋv�J�y���d,;�t���<avrv�C��r�GY�nڐ��f��0h+�g.N]������Bp
t�ؓ��d'F���\cvN�qKGoCl�X�\tm�>���-ۖ��:���$�r&�F�ZY��kup�F<�໱A�@�9�]����-�Mn��p�v��^}UHWp�:.CL�������Zk/D�2���P����\z6��N쓀�h;d�`�z8{vc���dT}�AnE�r�6Ź�&����r�8���F��1ðksGN�sv9����^�8Ǧ�%�V��Q�WV9N6��[y�8�>�v�t���Q�b졵�.��3��unNy�4�+�nE�W��TX�b�w����uɻ3>0ݷ���ی�g���xJ8���8������]V����ӹ5ҵ�v(u`�;n.���C��⒜7(["��Ǳ��uѻݣ��x�Q�c����9��p[��ݧ0�{nʲ�� :���uѡz^���n-��=p��%�t����m��vۓ�u�������Zd��Zq�wk��9����;W��f��8��@:�G��r1��6{�1۬�<;^�g4�4g���y�2=.�)���%�7G@:�=����M����p{yp���"Dp��g�ۦ�rsČ�e��yơ�Bq�^Z��0�R�nW�����e�URƎ7S��W8�<�<�=��;����]\f�b�n���ɉ|��Og�9b�jz탵�9۪N׺�jm�\����rrH>j���F��\��c<���k��P�6^4�O��w<��c���blV��<��ә��\�e�ż�姀��n���mӗ��K]��ۺ�u�7P�lc��c��[g�qɂN֌����ؓ�[�(6X�蝮M�:�NN,s#3V�Cm�9]oU,��<v�nm՟.�t��u�ќP�����vz��]WWr"��K�v�6^Kv���E��ۛ�-A�Wy�`A��g���K㛉����s�Wpr��=��˜�&�ݣ��� ��I�	�t����j��'�w �,n�f�sv���Ղ�!��u7������f�ˡ�xz�v�4�z�5�q�M�Y�����햋�+k�s�3=���.^�yz��񫭹r�)��B�ut����Ny:��l�!�gZ8�ۻy�҅��&w�=������a�z8�kq�%ū���w�:7<��Y�A��#���Z9�ا�Nh����q3�81���*���y��q7U���ň�[g�������Vzi�s[V���/���'�N�;��*���:�r��eX��<܅oLck>x�NLP��n/2<�c��8zsu�pޭ�r��Sp���ӈ\��F�g@E7f�P�v�y�����jN�Kp6Sh����ݺ
y�тs�ǟn`�
�H񖱛ʨ.x9�k�Ov�[�-uT���
��n��[<�7C5��ݎ{��:��H�x�Ǡ�^n����T�������x^���d�f6���nM���]]����/n��n�g�g�`kb�;�@�ɭ:x%�i������;9^���r�pIWnzݳ 7�-�)t�q�F�c[[d�Wq���;sul; u<�ٗ�k�y����Ƕ����:L�ӹje�Q��m�ނ��6�@u�:,���=o8��ڻ:ݭ�;��v�>�4�9.�ڮ'ۍ��*��yٷ-�Wh�V��ុV��N�7N�=���a�s��.MP莼�[[���;cO�]f�d�%;h5�3k��n�\�eȰ�&���6N5g���n�(pE���I��)�v.��8u����	;����B�Kd�糩뭫x N݂�y^x�4;qԶG���Z��+�s��s�'u����vz�<��Zsm���g��Ns�Pb�/����]�Ս=s�S�J�:0��/e�Q�zî�ж�{lX3A�p��s]='T�rŕ��]^�6��#��d5HW��=�����Tyk9�ϔ�	��0h��s��T[:��c�#�M�L�N��@�Z9�˷!��؊2"�÷=i짉�V[���+��6���<�m�7M�)�7�̙vr�'��<�^��ց݈d��Vg��;t1���N��k�&0��ܽ�/3swn�N�q���wad.�1����̷">�*ϫ�{�;��h�إd���Gs[����jNvר7Uc�$4�t{q�t&���x����p]1a�*�]t�a4�.t�ן4�i����Y����K?�b��Y��31,�Y�&�ĳ3��,Y��ň1,ŋ1$	ff��Y���X	,�%� ŉ`ffbKKfbM.�?��?��/�?�n�Ȝ_X`���Z5��
�F��Pٶ��x������c|v=;�o����I˥Yi
��)�sދXy����>���` &��C��R�{�����3~v�6��d3",y�H��YV�i��n�6��ll��̀%��Wt�/��^VQ�h�B��e>���Xγ9-[���������f�U@�z�N������N�<��L
c�w��~�*w�EX˫ e�u����;�։�~!\�S�<�6S�~ 4��WT��Ȼ2��7h��p�1r=���={k�����mKW�aߴ�33�g�sM>6 o܀�s� ���㊑I^�ٙarb�R=�)�!8"�X���Dٌ�vk; �j���'��l�|-�t�@�t�X/Վ�pU�#l�Ǐ�A�ެe��	��x�?��dږO����30��ڡ8�+�oL���
G}�w�l�4n�w��ޜ"�_��~��[�[��P�^3,-�Õ�[�`�^�>�l�
�}y��z��{�:$4a��WkVȥᙺϮoi�p"�_�p���R��M��$^'���7��\�lx��tpm�Ը;y)��n�
E�ٹXK�ۖ2�ud.f97UG����nM�����ow��yx*��g}�
7s,�v�S����*I�މ�<�0$ohK��*Q��G4�W���㷬�.���ώl�1�y�l�m׃q�m+\n'=��|v�>�KUK������]��\y޶��Ƚm�rv8�3p`�r�(�yS���y�5Hk��v2�gm���t=M�y�9.u���{;��û4ۮB�ϝ�Oo
\������������=kְ{c��-��(��l�i+ML냎g~v�$v�B��'��*��`�p�%�R��D��x䕙����@�{I�������6�vY���� �z=���/
���d�c�G����̺���/d!.�|��>��|ZTq쩪I2�*VNװ�Z*�N�"��-欞^r�qe]��{��&�8����9'��2֫a`���p�C{>���VOn��v�I�c4�%xU4h 4�Z^17PK���1������M��mv�������0sR��1W���]�w��o�,��M�{N�PX�tBelM�I�w=.eK&�x�Y�V/0U���h��A�"Y.2��o[�=~D�u�dV0ݘ�ޟ0z��Y���o2l}rhKJ��#f��˕�~"(��W�J��g�P ��ˠ���<l췆�s
�
���[J���N��,�/;	+�<�C��@j!���ޫ�5w��{ Z9f|��]X�>����dy;��ž]���.}�Oǽk&�4p�����hVx���Ţ�ht, �h;��3jw��Z����3��9��j����up���t��{;T�+%Q24ē���ܷ�U�ˁ݃�R��׃:�Bfu��h7��Ǽ+l�*�0�Y�
d5��>�7��w'��K4 ��U�@���D]��DsZ�*�5��u:�Ed�d�����V�U��=�v��v�6���U�IU���K{ϻ��O���{�@���b��<vK,�~��^ݹ���w�)Ѭ}���}�6��]���#!��a0�Rӂ��y�h}���Jb`U�o"L!�9�\���ѹxƲ�|�������n$|"�ӈ���绻����:�R��%�m0�ThXM��^�[�#ӂ�������,tG�i,M��m7�5�*,A��a�+ȝ��2��dL'M[�����	�d�⤪����F6��:D7D
C�hY��չm9�x$[}C���r�ږd0�C�z:-u���������4IѰ���ɯ�����æpH"�T�*e�`���g<ge�ܓe��4ӌW��ܾ��d�^�0�l�Qo
�b�Pb��6H�E������J�g2����ʼ�?fi$�5���#n��w���s�3N���� �.2�H6�Mqt���0�ɫ-�b�Q���8���,��&��z���>����[�������%����Xq\�Y�`ˊ�(�:6��d��$�z��kN�Q�j�~�nV�J�Aފ�F���R��l��[��r�"硷����L��'�x]m�_�h��1q�
��L�cm粨������ĵ��v��H#���f^y�Q���ȲM�:+���x'�RQ�գ�i|�L�#�nUo������kx�DT�<�iT-�8���n&.��� ꋛ�D�*���ڡ�d�R���6(�ɜA�*)w�	��	��� ��#�
�l�8kj���xme���d�E�d���\��ԏ
r!D�q� �Z/i5;�>��|�^��'�tZ��?��B��Dv<r� ;ݜ!����Y� �8ȍ��38�hEfM,��,صT��h+yup��t��0}*�I됎(^>��{UT����i4�	ᄽ�.)%�A����~RP^Nu=8�Ga��>���6��-�A�1hӪ�[������ynV����-*n�`��Hy#��������!}�:�� O��L�304TIW�=>��<s��iv˧�����W��xE����v��xɟr�,]���Y��*EL�m�!���_a�K�w1��= ���߮yu<@��e��c�^�\<jz��)c�����+_��,QW�ͷJ�qd���gL�����lqh]�֔�Ӝ�6������`��u�tof;aXY��U:�bX�`ƳPE��f�ɪ�d��|�\W��I��K��X����Cey�S[M�T� ��5�*���Ű(J���存`�
��2�l�
�Uj��84@��uD���Ar�yS��W�� *Ē=wǔ*-�:����R���C��n�[a�fQ�&7
^��k=�-1&���c"k�a@�������JI����V�ߑ�^�����v�2 �;��֫�MZ�����L�
<�2<Y�!��H8&*&.բ�6��x��G�Eu���ف�N�����h\k	ѱ���^y�u����1�rf���_D�hu����~%�i��|h��P6��X��S��j4U?UB���2o��s��� A�Ã0�c�Ʀi�U8���mm��C�}��m�ReU�W��(n�&����X��#n{+8���0r�s�Ǜȼ2� ��>�+�wW`9F��"��J���vTI4KE����xf�ʠ*u���ͽӁK��,���p�A�	oOi;٘����K"qc%i#�
��e���NU&A���_M�"8r�k;IO��ں�M2m�����؟BW���J�Du6�ɛ����w�2�\�v�-%�<�FW����s^j*��3N�O���l�x���H~��c�]*���]�[��k�y7b�8�\���`5�N�	!q��Ғ���[hO	�͑�b'�J\�)r�d��:�O���Nf�?�m�V�5��S��Ev����W��]�tq��^/M��ƺ)��:n���h�u�v�&�y�Ӹ�%�q<kn��,r�S�5��/ims�����[���8�J�<@�[9�5�҆͜�h4	on����=��XR5G����ݟH�1�	V8B����9���6�3N3���լn0B;Y5I�UA�ޭbJ�E��s�����l�K}�+��<;tx�f�0D�P��B]?OkqH���-�͖�wYt0�p���r��Xq_�Wt뺹��ϵf��է i��(�Y#W��s�t��O���d�q�I
BJ*�:d�����-ӵrno�YP�nfB�&����gopT�����Xk91Ki�̉�24�BF��ffTĩT�y���{=��֎aS4;�*��h����nO��U����b1#�Dd����ǈfb�v�r�Y�K"(��(��Bv�,��Q�.	��%��=bȡ@�Ι.O,+d��ߣ��s$�j�8�J�����O�0�}6S��ľpk}g�,��ؖ	!�Xb����r�kw�x���� pT��<Q��I�q���L�X5�n�Y�B$"�2�R����8���̳�k-j+ң�����Ϧ�G�O�5w����=h�b�Vu�V��|^B�#A�j�څL[�d�EE7Lx��L�w�r��k��{}��c�2���vp�����K�r�)����<��I��ֳiƅ<&^LY�5+�jB���mt��@��?[9B��
']�u�(e������F����<,WaTNo�5����N�0�j�g��V3��6#�۶��x��gV��k\���:L�
�w�ӷ�C=�0���:�Ǵ�6��f n�{@�"�#�{ޮ��;��"���χܰ�;�����5�a�x�f�e��#P���{uF����:P�ߋ8��d��.`x�����}��v�T��b�����ew@��]�Q������Iඋ��y;�M�պM�f`�R��)QÖm����v<�ˊ@T�a�v���uq��|0]�ʎ�6u��h���Ȭ+vKPhоGo����n
\o�]��o+)�_J/A)��>���ȸ4᧭b�5[�������ɡ�!�:FJ#���ڍ����D�	6 ��V�8�Pb���%��sU�0sq^s4XQ��*X�NӲ�<�f$���MvmZ2�t��p�r�i�#��:+-N�/l���Ί`�Ze��I�n���M2��93���B^�;y�����"��F�@�%#J\v��uYly��g�aH:��m@V�[i�%�]�{b�"d��0��2u���0"�'�~U�֖�v{�C1Z�=�\��~[���O�y���q�+�����*�Y��� .i���.Wp��zym(`�7��=WVl�y�����ʞ�b�*>��~�mF������C����7p}J�$)�_��]���J��Vw��T��m	�O�9���F��zU�ichJ�p'1ef2fr�fg�X����}�@�v�8{�k����{�mE�j�{DK��Ct.�F�Q�<���]��r��(�X���c�hƂj۬>�Sb\QNX׮�sʐ�[b�#$b�~��d6�	�P15:lNR��:)�� ��@h(Og�33
�k�f��5����:�/E����3G�I-[�O/G�f튼����ٽ@`&�a���o<���E�:�M�s�>�[��u�[E�s�mH�jt�� 
����f��TA̡{K���/u�ԟ�5e�i�5���`�M�Y��N�x�ϲj(
l"����Un<P�� G�&�h�@�q���u�E�|��x���x�X��ዳ�\Ķ��rw7uM��mo�jhB-��Shn."ǒ�h�u��U~[��'q�%��{���Xs�lyd�L��|r�{���0�S4g+/(��QӷZ�AV��K$��C{��%c��:�� ��A�1s�^�t�5m��L6�ji%�Ly�n��p��$�f�\��..�o��ױ�w�Y�Z�cȵ6*f䕸��?=��Ja�E䦓̵�^Ł �B����"116�r�u�kr����C�BlcI�Q��P��.����/j��m� �����-;w��|�M�p�ʱV�0Ap~~�@D�mZ�u�`g�2��ս��ι\I_u�b"��f=yN�0C�H �'P�j�O��T�f��Q��q�qpNj	*E�@�����ylw��v{}y���Bm�����NͅbD�x�##L�칹L-!2��ӥ�+�qu{�J7־��ů.������ZL�r|๶�a��8.1%wULY!5�7n�Ǵ�}�#����B���]l�ے�+vuE�aJ�ȣ��*��Pf����޵:mGƸ;|S� S��p�d6wVN��xL,�"d�qx������, �E�l"�%�W;O�M�7㴁�`�Z�D�wu/L�(ۙ���2���vԁ+���v&S�q r��6(B�<l@��7OqG��M�-�
/�-�zs}
4屩W��� }���<*s3UfA>�s���^�p�	h\{[�Fk�X�p�7J��S	0)�dm�9�����d����QzL��)Q�B�2|}��,��c=ɖ/��U���Rͪ���8�z&pY�UR��M�������@n�*�u��ʴsRj�S}����-��g����I���q��wl�'��Ii�mA$Î^�g���մ������3u\�;�� w&;cX�WOUe��'���&Mu���PQ�(9�C����]3>iܧ�i�8=���B����=��ӊ�k�mcς^�y�E��{t�tݗ�I��k�r�H���Ne�[�U�����[�� H[��G��F������ ��/e��v��Q��t�ۖ�u2׍�xMw�֦6��'Ȳ�M1�TЖ�Svb��,H8��A^��*��3�C�K"p�����uci�����3��X&&i�"�7.�� s�1t丑Ed%�o���Qs���r�G��|�N�! �W�~KƷf����N'(p�% ���߻,wsJl�S���L���[f�i�U>t��Z�(�J�Tn�P�k:�v���������chQ�Ǎ[kd'�����y��eIԔ��6���Ì4�m�2dc���q&�@�5�nNH�}Weϯ�@���	��.ƊN�C�K�] 'l����틆�,�`�G���s�z��͒�w:�̣�� FӬgod�D7�µ��y~T �#P�!��	��_:uڼ�6���YR�#y��6t[�F�e��#��z��~��מ��~���8"�]I�io��|��j�Xy)�P�;��5�-�a@0�L�f.�ǳ� <@�e��ʹ���<#ǲ�ߕn���<]֮y[C�	���wKs��g��%d� 3h���7�cd"J%��R��X����3uw��|�Q�8���|����8�����U�ޛ��l�U� +�B^3����Q�oZ�18���Įe֟����ZJ����?[�\�޲�y��^���e���$(�N�2��_�PɝW[}��dV��������i.XRܮ��d(�u�wTv��c������jm[b����f_'�>�|��4��Nj8{o3�ten�����
o!մ�n���#J3�̥6�{���t�.ȇ�u�\�agw�Z.��g��:eX}&�����N-XX�� ��{O>Q��|ju;�+����޳�N��������!��ه��U�����]���3sVFb�L��i����P:�$'��[�[��!�Tm���K�UԾW��-���n�����ϵJ�u<w�觸��ۤ��i��eYt�v<{�C���yp����i��e2�j��ûx�g�a�=@*4WgE�����t���y��tx�va� �Kf0M�2�]�X����Я9\����z��cʶ���k|sK�z�U���7�^�w�P���Л���%t����U�rm	: �C>��-�i�656ʽ�V��݈����c��;���u}-�#��8��wI,�M����#�������U��8��� Sw���nX��˒6�xڭ���Ie�iŪlox����p���������k�n���/7���e-�{>��B;��n*�/)o���PוCb+��y����&������w�J`�t���eR���Y��3-%�+Eσ]Y�2^u]A�&+�K���1�BM"�d�m���5J��Um���S����P��P��y�dCam���������L�gnٷDܻT�ҾрT|�%�Z���s�򼽘!<�����]WF�-ѡ^{zz:�ܡw��ڵ�N�]cv,�3��C�]`��P�ȼn���ۡ�N�<���k�FD��gUu�A��[Di��g�<r��k�Fx�ZC��.����ܘ�Z�^�p���S�@��B���.���8˞S��eJT�4v:��i:�kG����i���m���;<+��g���e�nV�"�V6���"n��<K��tt�;z76s������S���&5[�s��%��zJ�L��s��*�\qc��X\u�+��0�qp�����`��v�p=JU۵YI�����t�z��ʜ]�5���ݙ�ϭ�m�����붐��R��n
���b�1����b���c*��9����ٞz���8$:�:������Ȟ�1��u\�
�r&�rt��u�Um!�8T��Ѯ��#�{�7hy�ڛ:ݻ2[���N������;�P�Kf���g9t�*3��aLG����HEvX����i29Sn{j\����Zo�.xL+���E�^y�ڎIx�q:s�:����<�H���Dc"��ǵۙS��g]V��u6�{�Q����>���8���ܥ�{'��E�[�;�գ=��2h���m�g����tXF���[Ztb�(��;s�5���tP;��;^$�b��Hp��pR!�N���N	��3��E��J�)pۗ�N����a���i8�bz��l�s�Go9��z��t�9-a�8���gC�m0�\�:Bw`���۰��*]O�:��w;.��pR��g
���vW���S6�nt����.�l�� c�<sr��.`{0�y]ŋĘ�a�퍈�:��N,�p-����y7Knvx�G�k�]��n��!�&v6J�Q��jm�:*��{O\k��b�Θ�����X?ܹ�h�d?	'��e�b_���X�m
����5���=��|q�������c3��A��1>?�{k�b�P]��Z�q�$���k�-�&b��������k�uh�����]$2�Ofy�&�8�5v��\�D�:�K$�c��W�L͙���ߴ���-�� SM%���1i����o�իu��4*$��ޱ�	Q3̂���J����Ck�G�}��\1hK�2u�JG��2b@��{�v��[>+���)����F�^�ϭ�=+N�Y������ ^L�-��LL�Jk���%�A1`+lţ�*.�!/�Qb�x���z֗�t��lš-~릾k>!���i���}DTW?���ʵ����h�����b^?vň��1x�ZTD��҆h�����G�c@d1C�/��T�W{�#D?���@�J.jif�E�K�ݡ����3� ����+E�ګ'�ލ�Qhܪ��kF1Z��s�в�+�4�.�F/w�{_3�/�3F``N�E��J���&b�EE`ק�k�J�bP���3q�-�B��1/�����%x��g��gN-z�K��P[�K�1t�c�ؾ!���;_��n慣��;[�n2Ш��y񊘘�%c�M�֔�j�����||%��1hšC!��.G�ْ5�%�1A}��k0~�;Ͻ����MƸ��	��d2}=V��L͘����K���[��,b�蒦.�����ǘ~���4&f��ե�h���>ڋ�X��\3BZ���pš)�k˾�uV�[S|ј���v�s����k�@�f.������-���?��z~��)�1Sb�L_��pHoҽ����hW�b�i�L��1l_��,\o3��_��ZLH�p�D�c0�>���=���s�B���$�E���{{���يy�%���n�٘�Ĵ$G��&/���b�߃�~<��t�kn?	*b�4�:Z�S+j�o��~3]�]8���Z���ġ�m�H��NL�ӄ�m ��4W��7f�f/d^(�v�	���Mlp�1ƇW7n��?G{��;��i.�$���9Z�]3⊉*.Ʊ�����ߵ��L̍�,U��-�-�$�\���kI��Ί���C�d����	x�!%�{t���J\Wdl����:)���{�!Pܘ3��ؒ��(
ˉ>ݻ�mA7���Pt�����f&S�w��Ԟű.���X����}).9SV�M��� � PK�~1S2��7�.]��Щ���s�8$�EE��_i��/F�13)����Z133����+ZJ��4 �����U%��߾-�.�s�\I�1 Į�d(-�NL]�洲	-��҆%��ŉ��fw�����ݟ6����i*g���}�Z.�ж/���c�'-N��*�w����#�>����1wMbw貉Sf1A?v�X��KBZ+͋�e2���������,|kͫ�T���>.��c�yyG�sS1a(DB�g%����}@šA%�ׅ��kX�h̷�;��k�}�/���Х���1AC!�h�k֨��8}�L��^�撂�Zس����Zg�����0�C�Z�����yD��\�w�Y�6QxK���g�ۢ��%[�L�>�P�,�+�
+��-L���g�gݳ>��F�,/��d���z1�� 6Ql	9��,��f�D��Ū�j�Y����T&K�&��6�0�S��V���qR�s[�+N��J�4�>�ҧ�wa\�P�� 5#�,Bi�@�GL�:��̦ �S4,H�%��P������[���#��uÎP��@�QSYй�;��P�m ���>�̧I"�%�1�gа1QT�Y�(9V+ų36r/z[/P���)�%6LO��M
d"j,:���i���kw}R��ܱGQdo�@B��8�`�𭜥z�������V��H�R^�@�zP�潻�����H:�mm��o��zi2)����+a�m �����F$>'p)Y]\�rp�J���D��V�l������,���9�Yi�v��kN��u���%�u]��Т%��;�7<�X��:�&,u��$C�6�Z[�d�	���7�j�JWI��L�[s�J����֘�����mIEP�rd�V��T���Dާ #�`:�pH�'(�ʵ>�G�t-�<�L����`�I;�},;$H�kBMC��3�# (��e)�}�d�fL���}����#&USP�$��;ʨ�wL��Cn�9F�7�z�"�t�Z ��okd�廈��{�HF�2������"��j�����,$[E�XG��^�{b���Oh��ei�����uh8u�*G��<�B��,��=��<�F�O6:>e��
����	s��p�f0�/_�Ju��}�x���X��^x�u�_��=Dn�"jS
?qs��f�ʿ����x��%�o���e3�I���8	پ~4����G� ��ʂ��×fh9��� �<o�A5B�묔�f87y�����H���^5�N��zL��r� d��Y9m�۲��
˾w���1=Fӻ~����<���h�!V�֊�&�)[su
*R��é�N{�� ��-�V�C:�퉫c�!�^۴|1�i~c�Xe��o1�ڬV�R����C^�ٍ\���ΛZ�d���5ť.wD,�X ���@���%fU�s�}6PS����NC�zh��D�+V�6�m��$ˇ��X۪ݭ1�y�"�na�I�k�D��7d�^Z��X��½[�N�X8^��Tk��:�6mS��nLh�k`�^�詶��s�)��x�Xzj�b�T�,*b8���O+Y1��zJI�o v�-��oX�c�y�d#j��m\4�]���n�V�ˎ2cT���.�{Z���Yգ.86ț\�3�u�F����NUҞ�|��a6�����	�bo��,-�͙�;	�a�p��~��. h���*����	�*2��T��J�V�a#إ��A@gQ�e�骍'�27چRԚ��@��8ԓ"��ס�4Zo6��wq�(րH��!(B��jP4��Ës[F$]�㾵1��w��o�W|ݳ3�!Uq��v��S���;][�� �Ӣ�(�*���+��q�`l�;{��+�-��1td�x\"���AP�#yز�gY���G��%/e�y��,����;#-���U$+�~TF]��ȵ.h�:�VژId�迃5� ��aR���f��Pø�h9w׭�[�k��bٴD�>j���3�Y$PU���[�ng�6ٻ�,���y��8k� 9�nj��ƫ��+���4��uIN\������s��}�K6�ӶI��֓,8L4�7
@���~���˷�u�AR����qfg�{�e�>S�]mu�Ӣ�&��ϘhS<�GC}^y8��\�0$V5��^ڪ���D�)��L�`��7e9�Co��: �@ς�#�*���Y~�n�L�~3�H~�ku�.r��"{|����]W���-;2	�\�I4��h[뽱�hҷ)�m�!�(n��k`8m�]�N��F���ݚ��h���ݿ?:�v�d�#!D
 �l|KP�3%�c�ˣu�#4R[�V� y���{5N�a���q���m��c��v���عG)]m���c��6W���Ĥj'v\|��԰��l�`�	܍��b^�<�C6r�I��p +5�%�k ���7���Q7���o�;;uZ�	
-W��IyJ��WO�IR[��a+q��s��j^n�ʱ�6'��:hB����%�n���凼nt oo�v绞���냩� �e�b}��1�����b�L���1��n}#%L�:Y�]�0��W��n+e[��4D�����N��y���^A�@C��A�n�)������f�fN��9!g���Y��M۴����MS�h!7��Hy'�CM�݆S���S ������.��
`[�6=��^H�.,N���!m(�5��h������Na���kO�B<��f�)���đ�Ꝥ�rp���
�Y�>y<0�j��___�6�أu뙦#���g���
c��Ǧ���(W��Nۮ����M=a`�m�PtL~y�{Sc��Y��]gyj׹ާu^j�y���!7h��v�������YY0�W{\6�#�g�a�+m�Q��9��yϫ:Y6�Yu3'q`;{Z"�e!8�^�r�伻ɚ�!��GȠ��97J36��ZyS��W��A�����̏d^��U�^���꣥������rF���������\��<�������i�zr� 1���_T=���l��������f7f�����S����d��%��e�r�S����q@
�����2�%��A¸���	L߳�6��D�g{�?v%�7�>�+p[g8ׅ<W�ѻ�Okdߋ��]�� ��O(�?Zͼ����-��f5ǵײ�sw�;o�ҫ�݁b>��l�5�֞,K�%�[�V��;o�a�|��k����Y�Dx!!nV_����f)*D"�����<��~c{��ͥ�WI�9K*�U|9�j��҅U��l��.
J����6!	�+�u��ZEB!�F�V0|�{���ߛ�}�cu�ѐp��Hqx�D����S�Lo��Q�� QncC�����O���Rfde���$�ZVgcj����~�v�cTʫW��^!Z��]#&���S=96�=����~4�{)
��׻ڽ܌iPLl�#��]߮�v$��9X�6��X�>���h�ݙCD�}�)�,�jPu��w\�f§0�C1�d��527��R��]J
�z���'���k������ɖ�z|����m#��d�������$�����S�ܳ�q���/�Ql��~�@�<�=c�4G�}�1P��,\�W�G(��pb�,0�z��U�i�إ�s�U�cb}�;KDemiy b
H6�Zw����P�м���'U�.$�d�~�fv�T�=�/���`1\åJ���ٜ���e�׬�PobX���'$��b^�^�o�A�}k����j�Nr�6�-�T&[�M���%vd��.�9��fV�+��\T"vѵJ�i�u{���c#\L+�\�Ӈ��Lj/�Q;���Z���h�bo����2�i�(t�~˺M�~��)q�Y�)EDPa3��;��,`xAqX�+6Y�v����(�T�p���='l���ײ`��ٔ�t��ˍmm����Z���k��Po73�3B^Ej�<%'*�8��{^� ^��??�^��ٰ�q�ɝ�rƜEk0��k��F���;�CV�A��.��N���+$(��̋� 2tʱ��Ԥt*)�N�Nr����OJW����7��ͺ���^v=(��]�4K[�r�YM�݀%f��^I����\>�I��U�1���d�8�;��g�t���U�x{
�#Ө��۞iZ��S���n�Z�^�N܁.�Əi�=oe������ݮ�}m�WF�2헲d�K%n�y=p<�u�/*��@�d�絎��z�ּ�#���60����^n����Χ��2�t	픍�۠Z�^�W��g���(�����K�Y�����~��<O�U���n^�«|�uN����-�o�����_�R��ǫ��8&q�uӲ��$�zۮ���^y+�\�LN�Қgh�| �תL`/9��ۍ^�9p�}'پP>GK�W͐�	��g�R�>d���ˮ}vk�f* /��Ω��G-��lܴ��z�j�@��Gv�q��^��MA���K1�գ�(7��nUzNn�ɜx�/Hr�6&_�$1��Z'bqO���.�����d��#C˲hح�Ю��_n{��w;�q�.��@�f�X�۹�<��C�=��v�\j��+�c�96)��6w\{4������m�zV{�����Q���7R�(�{�-�L��:��p���w�R|�ڀ=�ԓ�U��}c�]<�x�#.��֚bנǴhaÆAE�@Yf��mCB�Y��ƹ*t���=�І��I���5��9�Z��m�U�F��}������ǃ����)cpy��.$����i�!�d�1��S[�5�-c(j��&�A[&"��j�/م!���+jb����5��ލ!2�c[҇����.ܬ����i�13��O��U��D�n,�;w8WJ.��nmo05<'0��1u0v��3��Fa��b*��w]�瞚Gw��Ka0KFd���^��c�h��|�؊�Wy\2t���l�"����2�ՅOA�3���1�+��X2����ÒɳF��E{r�n�g�_�A�0t�t�Nyb��a�v��f�W~������-����`��Y�7aR����>��΢׵#~��*z�`�ܔ�\F�ѝ��{�3v��j���3r��|��A����ʕ#E��^�MՐ�̷t0ku��C��=�ߑ����8�S�}�Ӓ���k*���ώ���I{u?_�u:�=�߳��S��a�J�	��������j�U�Z1jg\Ֆ���@���T'�xf�?OL��)��|�'�{��3����O>�"/&���N-_��a�͝@Fx������QZ�î)���R�|w'��c��m߮$�yQ�P���֙��0fe��s6���ȕ��'l�Va(���*�=H�+�G�/���x����8�M2
t�0e�!E`Ev���x��9�޳ټq��V8�4��vsn˽���

�z{��.�yW<�e�o ֖�L�3޵��/��#��6@ȥ��G+w�{�y�y��cq�-�h�!��w�}�sl%x��5]��+0S{1�̩��m�(����3o��u�P\޴���	�H� �"���T��f�[X�N����kf�O{�%����aQFƴ�w�^�K�g)�b�az��=1^����;� ⅖�e���0vI8! [
�}�k�5O��Z�P��8#G�=�H�C{�DF�<;�f��J�1Uel���T����W��V��8���C��$8@ ��"u}^�i���]l���U)ys=O}��I�:����Ҕ���ڛ���:���fV�iU:�)3��6���4�O|�G��DAn[*���Ǭ��Z%�� ������f�{��p�>��ޥ�Kw�hC�쁟IG�c��E�̓ w/<�k����w3$�"sr�$�� N�b}��ǵ���f��.��M��m{�+�$���=��6�!����NN�v�ku��@���ᴫ�0L��)�{�vMƀ,�,j�a���2P����Q6��!@�[�rI2�s-˯�y���b��E���f���g~±T��W�{{��
w4G�7'q'/y^��f�����1YS6zyL/-W3��K���R+sc[�`��D�S97B=��W�U���x����ھ�y9w��Zy:�5�w����c����a�Ϋj�d�kUo0�/-u(�ș3l-g΢A툎������V�Z��n�)]���S2ٳ�,�]�@� �Wg����M#K�Փ�����w;�vy���na��<A�%�N��V���Q�󭽚X����[�G�\o��P*n�a�5t	Z1ggf��JŅ�^U��f%�<��kk���9-,y��r�X��*��/���ǑA���ݺݦ��}�\�8�<')��ڱZ�*~x=*:��ǵ�3���N[��ri,�}t���^�xo�{����`9蜙qH��=��[��{���|w7D�Gɜ4��/iU�b��4�`u3�Z �sm�l�M�Od�}(�-�[���<�A�7mcY����Z���Y��z{�����wl��c����CM^�y�W^���r��yʗs���.���K��[�je�o/:����δ�w��5��P�t�N��*���y��sĢ�.���Ed� K�{|����@��ւv�RnDT.������O>Z����ǷGT�C�aK�+Mr�V�����܆�φ��Y�%f�pd1괨�P�ݷlA�p�\��ʇ�h���+*���V$�hb���g,��2�J��B�YIE��A9���a���אh{sN�g��k�f��� ������̨�N��mZ��fX�ϝ$�n�ҙ��U�=�L4g%w؆ۃ����{f�vj7y���5�r�2���J敍+[�v��a�.����m4C����[sfｹ�l���z�y_����&e��eXZ��F<��-H��A����%.�j�WR������j�u��w��5}�dD���L\
�J��8>��ay=�5�Z0\�V�����U"�N����VD`h��s��-��uO��$��N3��w�q��=CG]��<R�[ґ���{$��
��'L�k�G�~~s�[����@6�H���o͏Y��B��aE� �p�Y��|Ѿ � v�_c��ov;X6�Yz��[8�"Y8b,*�;�	�e [����(C5}l�025��[YwP�����SLm�@�##q|��f�Ư=�Oov��%�|�üP5g�D�c��bA�?]�ֆ�>/g��P�;�2)�ۘ���x4������6��Y~s�q��P�T����IC��wu{n��vY8*Ql��6oVh��r�[D[�CL���;(6�ev߳U7�g��LmY��_@5}��mL�.ҍ�E����~Y��W����5�����V=��K)$��kz����>N}�j�����^�q�~��z��]�eq~��;o�����$ԋi�&��S�ڜ�;ώ��{�k����>�J�i#|�9&S�Z�0�\Nx\��lSn�� ��s��'u<r>=e5�킺��v��6�Q��e��lW!�^Od�{q����=M��.Gu��A� ���W/)ƺ�c�"}:ۡ�AO����ni�_]�֭��
7e�������y����3]Z���'n��<��n;o"�{#ڶ����4r�i2���j�sl��JGj"3��-L�b����7V����{y=�Qգ�lI��Hc(�{S�`�sg|L�n���攠4jq��V�����[|��/��d�6W<�u�὾�;]��J�I�e�'�i�R����*� �rٌ���p�^�Vc��:0��񫚦�wwx"����1�sV
A��(��՘HrH.Nx�7k�w���Z"�P�E��@�[M2�ow4�z���E!Z���:��Bٯ W�j^�K�*a�f�T��x>�|��}�n�����6�,8A+�D^pPlת2K�μ�����nzn�π>��U�T?p����au+tN��cw����z�Q+?�lf��U^�D�u�HAP�8]��zfg�Zv�lg8��&����h�LRǾ��R��8T����m� ���9�^�ߴ"��^�0�����p>T��4}&�+37Zi�iBHQ�mYy��v���w<9Ӿ�.ؿ�}k�v���lW���PmR��R���)�{�=�vE��N4��+�����W�-Rl [i$S�O̊��~r���w)��ڤ-{��8xR@]���u�pVg�<fz�Ýp�~v/����Uܪ��~��p�̣s��#ژ�%�e<�r�w�Xf�m'�����X�2��^h;|!����W_��N�0u��io�/@����D���aL�6�Ы�~�W��q,���A�BaUȇ��W�N^�^^z�E	I%>��c!  �E�Q���>%xy�g��['][�5������ta-d�)=Y�o�h���<d�i����j�'^�ﳯE��ׅuUNs6�ʧ��9��A�"�4�(�TX� ze��\ش����+�횜�ڮN���_��#K ���ȯ`�	���Yz�S��!�D�{�^�܌8�Q��$��]��C��)�K��a�gw�����s�~���~9�}�x��	�>��z��4:����3t����!5h��@E�n/xn�� ��-80��7��JU�f�`����N��9&y�����87^_�L�+�z񏲽�Φ�W�'�$V�M����J�W_���`"h���W=�>iw��z�u��=�7t^��4�볯�Y�Z�l��/"��d+&q�'�-�SPha[�B;q��m5	A�f5������/���W��V�
�z٪}��E��u'#��ent69�.�2X鷶����S�a���ܽ��x��������#G�@[^:��%ʉ�CW!C�sB����Z��a��vu�6�I�6�vFΪ}Y�c�$G�WٵҒ���%����l�H8�p��f��/�Mޛ�0N~��x]��apQ�噎u��СCEQ�M�z3f����^��Y�k�C�z�����;j��Th!��F�a�����q-(�� �b#oʆ�N֯a�1�}w���0�kU>^Os&`K�WY����;�5��?V���r�2��RJ��R<�.�q�u��ϥ���SI�B5b�mVڙ`x6\����4�ټ4\E���`U]�朥�t@캻��t���(����u�+O�>t�6���S󷲫�1���(��H�f���KJ|v�i��3�YC!}���{x{qͻwD
����=�to���Vb�9��j�o�o�+k�������S��b�uR�Gm'>����OMp�Tק�-��FN�<p/�J�9(p�5��ǖ�����j��4i���\���+��e�ϛ0Ō�f&|qhۘX��yj��ng���z�ZJ�,���]^'���<��M�yU���l����djL��6�.��/�'���k�c�S����7lA�^���в�Y�����}�-S�m�=��]1���s}x�"��Aآ)�\8JH����Ӯv�7(��Z�YY��G�����4`�����ԟxqua�v���eM���k5��ܔl�6������Ͷ�i۬
��\)��S2��ѭ^�ژ��_I�Ș�]d�P�d �\�Ϩ���UQ��	!8d&�h�l�Mj5��c�:��*2�3��-��
hd����-�I�F��>Z�0��N�����/�[�_Y��}�[��S��%RMn5[D�l����~ݟ{�x�'t{r��vc�~Kᵷ�6��:$S#�)E��}�L-?0�t�Zʜ������&��1ػ�f��B��f��RI0!?�BԘ�Y���O��P�ǤōZ�'0y�C���w)ߺ�E����F�E�'=��4���z��}BI���8�K;L�{��ȋ����{Xf����cU��:��T��<�QA�'Ի�=Z9��U�qm����P�	Nq�/R�|���%Q�*W����Z#��W	�Kn�C`�A��3��F����|��mZ{X(xֹtk��1�".�iHF��[	H��}��f=K�m���>��/+�sw��0Ň�u0�-�QՊW*>����.㭿`��T]�d?*�V��w*�W������`�n��<�CK��I���X�<�v�f����"b��0)��ח�#�d*�N���u��W'��5Z\s;$׷��]�& xk�]fc��	�{���.*�߬�^��R�̤�(4�e�Q�v%����qe��TdU;���f���
b�.JV�qЛ�����	�r��^�%�qJ�@�nΐ�n���]D��=�x��QztY��=��ݧS��[����X����\yƔ�]�ۧ���n�)�vy�}9�KO=�u���te�Ǭy�g��<JJu�����s^qu���`"�)?�%&�$��3�������WW����Y�=��s���Џ�6}7�^fi�/��p��92Lz�Vͩ� �#`��~	�UPZ�*1�v���`���3_�ixȳ{�~�CѹC)T޿!�$�\�"=�ru��¡�/`8F	a8HCB�	�[�9�n4C	E���-�fF������ax�۱%�݋�[/�4e��X68��/`m �D�v$9���'qlG����~��s�̙�8���mY��T�����ʕ��������ڠgڌ���o�}���x�1q�b�y�F�s�V)g_~�@j�������K��"i��Ƥh���.F:~�K��k�=�L����0�hAA�ω�W^���5AI�g��A.��K����2��
UOODd��g��'���ɏ��8��F={����������'�>�v�2H�[�a�q���N��𰚊�0�)���~s*�ֳ��8���h�
�1�G��cp+�����vRZ��x�ǫ�2�a���(��R��a��c��tm������b�U�O�{���ʿ*?D���o��aW��֋f�]=���B2n�z�ƕ���b�+���N��������9�t�u���q[�V����c�#*.��o)�G�uv�6[V:nq���F�1�2��Dz�h���&�Uz,xn��k�8ID��X�(ez�{�Ks�,G`抁����=v� ��J�J(��P;89��ug�W���!p�P`�K`�[`Q)��A��nSO�Ê�fTR�=���Sk}w"�Y��5�3t���+����iPuA)(�����f�\ߖ�|G��q��Ƴ�kh��)DS��Թ
a���gϩ����e�j��F�t���40�Wu��ק��-��6N-�_L�<����t���2�^���> ޿_���?��B,F���ʡx>��{�|�d�VƳ07اv�ն�e��}5 �a�Z�Q���|�O������<��;���n��xx�ae�tt+8��V@��ʂ�͝�>�n+΀�4tB�{j����H�(�h�K�Bi�{�`�4_{-n�]+!ل���UxX�o�k�ld-��w]�ub�rt��U�譊X[;�)�72��,د�ǲ��)�e{�_-��T
�j�=�S0���oq�S�L���vŵC�et�<Ϋ�tҧh�p6b�v{;uJ� �z�[=��l�v1�͝��DVڈ��S����I�^a��u�x�zk�R�*���}~�^�����b�*;z���%2�ۢW]v�r�vW��t<�ܩ��cW��*�נ���B�,��z��N��O��cڣ[jA�[`�͹��1��ќ�G����K�����N��u��wƽ�v輸"$�OZ{�KFy��P��T�v4�T�B���ԇA(q�]�����*��A��w]H��3���:���s��y�c����*=�1�.���Ӟ*Ę4|��׳��+�r��)A���k@1���4�*�tmﵲ[�h�2�=	ڐ�"�����WC�f@���|�`�$b�'���e����f��r}q^0��
a���V'���8_��^[��|�w��L�~
��$�}��l��g���vn�[�b��eH�6�������@�S�^�Y{���^���B����;�m��V�;=y_<�����x=Z�d�aa���cP��Q��H{ $�5�rl��9��vz�GB�����X ۚ��<w%F�L[��&p�����J#=��Z���$����,q��y�X��D��O;=<�r�K��ݕ^͓_�,�O���ܭa��F�oɣ8q6%�Q�b�1��*�,�$V
�u��)y;|d��*�����
�z��0�]��{�j�zv�q���.�ۉ��T^�:Pu�@y��!��%�������X=~����{q%����ʞ��gua!oQTqC2e;�9�չ�c���oo�`r��)��Nqʲ��hb:w3XW�������8+��x��p�L�7	L�b��ʢ��@ʰ�\?fn�B�7/^��d�"a��EL��
Ѯ�e4_^z��J�%|Z	7x�b@h�~�N~�Bv=71>�;�a^��v�2���]Mk�g�O9���be
L��'���zMuwFǵ.ɹ�ƢZ�I�Bl-b^�U�7��ծ�u�<��zk�M+�^OS��W_�IGl�:�/x��VY~|}~�`���Bz�.��g��~�kQ�rwo�8i�_&�f������b�O���2#c�'�嵶��#��T84�+l��z����7�M��uX5��%0 Ht��r�IZ��9��ۂ6��}�.6�mܹux�e�$P�H�
�Mi�5|jg\������Z~ݏd�̸�P�p�YPLLf�H�	���5���^���&�tVM_�B6�v�͍��d���)�O���;z= �^���khF�4P�l�9c�R��Z��_��ʠ����:�̨��r��/��T=���/�{���l��_G����+~[��`*�zQ�'ո6#��H���!{+��O���Q��nD��m1����HY�e�!�k�Qit��6���ew-���&�\��;#�7R9͂b�Q�:6���`�t�çn\��D��ع���֢�|�ք-Ԭ�(�x��A{6݁��;������ùc���[,����E�K��gm�e�\�ǋfM�vx��W:�ȩ���v��@nW��q��i�g������^����vz\�5ۍ:�R�ky�Ƽ�v<���Aʽ�:w�8�.T\�pw�뺮�u��+1a®x�۟'{r�u�-d{��w<i��� �A�YƲ�	��!�% ſHbsj���E��D�,�j���N��N4è~gt#f^���[3kGD�()������^ڗ�#�W]���%��·�Z?W�Y`f��t[�)j+}����Ci���kҗ.i��ޘG���.[x�{s��>�]�{�Ӷ��r���P���\H�Q� �t_Nc�kqj�7Z��d�\�F�ӏ)O\f3�������Ҏ��*9^w��=�/;Es6���]u�ɺ�����_l8��y�=�o�G���'0���S�^Y^��4�ܿ�O�g[{ ���ϗI�3^���ѵ����#�T�v<kڭƺBJ9Ok����\$0�Ab*C�J�nc���s��(�[1��5�;H&���}�{x��ƍF`^�����B���f��ޑt���DU5�k����T��шCa6Io�^,U{q�)Mͺ��¯�y�����$f-���\O���y*w*tA�9&<�*��b�p'=�X�W�9Y^�Z�af!���m����Nl�
״O�t�����\�8Gx�$W�gx/��L�t쮷�;gR9}T/ۏ˷��Bj�ׂ�F]��}'T7!6.9x���WP#�
J�lnήuضvJk5l��6�z�(\�î��Pd`�(P��Tm^��)^:���U"��w�)�w�3(WtYP쑊Ip֚�j�gq]����+Y����»uF:m�A��"���"ը�fJd\�MG�LDƍ���Zݙe�U�N��(>�%,��nY��Vm���i��g���ó`O1��<ܙ��%�X�v�v���7}:X��.�7�t�� MMMM��])�n�۽��7�빢�������Y�7��|^��f�'�G�Ѻ]B�eecL�Ž�Ьs��]Ou���u%Cl)e��h�83�C�� 7�>���Ay�p��b�9hb^�ݖ�^k�:���D�7 ����v��x�e�!��;�n�Y�\7�Q,hud�/N���,�4��v�8m�c�F�X�U�s��^̻�+s~�Lt�Z�*[��U��G
�ݛWf�M�js\��uۄ<��l2�D]n^�(��
p�EV��D�z�s�҂YJq�$��N�ٻh?�3���w�Jnə8�I��8ີ�3��}e�i�X2�ԑ�����
���o�z�3�:'{�}�8ov�Y����=8t�
��B� ��s7oV0�M�Z+��tVn����ni��Χ��v�sj�eN�4��SX���{`V�\ِ�u��(X��V�_3�ڸ�s��}�l�	4<��Z��~���{�X��6����L�@A�1xY��h����O�h��.�����SUU<���2��5UU����j�X`jv��b�m�5���	�5�G�����w=I<��=�'�;��v�ekW��/r�D]f�sbo\�V��㛵�Eps�3Kѵyc �t�Kb��)��U�<�a���3s6�n�X$Oqj�3R�S�E��n���n{Wat�7�q�����G;�g��XZ�i9yp�q+]��n�B{Z�d��jw0��6��d7Y::A�x{];Yۭwn���U[=1m�mȜ[q����Q�惫��v�f.����s��v9}�p��r<q_f�ú�9��]a��p�!p��R\WG����3Ǹ��O8ז�FC�O�Ec�p:.Z0��em[���V��Rg��];on-�8Nh�.��p�ҙۍ�5�[מ�\�gm��Ƣ�f{=p�ힶr�'\�ѷ�=�W�V�pnkn^����n�q!�rg�^$=�Db簼�ɜ�<냮:7C�U�u�z1��Ț�L{m�����%�ݵ����ՇF���<'=n#�;��\��t����6�I�h�]�byֻ=�=�M�N�=XCsuf��O[���b��.]�K����"]tN���l;��yWT�^�B��sլ�8�qݺ��c�I�i�gn\='��8^�p��1��ԛ���'q[������]-��q+��O0���tLÅ͸�]���0��=c�8��p��yOp��5d9���d�-�n5��ĹϙL���i��� "S���x(�ڷcu*�p��0]ָk�`۱x�Ӣ�mƳ5�7q�ls��}Q�Y�8v�aN�9�v�\�g��X%�f�k����l\�[�h9Ѻ`=G�t���G��j���{y'��r���dx[��Pv��ObG�������Jg�x�6����Y��=kuz�Lm��\j�݋�!;nz��֞3sG�8�fM=�Bv�nnsΎ��؞�^�%�������{��ݧ�\d�<C�����ѕ�=�gl�s�K1�Uqc���M/�1�csM�U�_P�;B�`�k	��4 �3X1�VE�ѵ����~zl��$xz�`��0�I%E�v��wM�A�]�ݧt�ѱV]�S�:�<��n<g#7+BڟLz�^�a�����(�O"����lH��D��y��;p�޹^�������߄�$��A��_�uN��Ȕ�y�÷����\f���+��g�|����:2�^�z�)QIhz��n��K���0�H�Ҁr̷�9�\Z��4z���𶃽�mY����߼��Ž�z�dZK.��v�z3,9V��&��g���<V��Ҝ�, �ټ�	�ޭ�$3\���� �+�~��[�;Ψ �߳=SH<�D9n���XH�U�Ҕ}�����ۿ0cؗ�0���}rw�(��PQ���}z�"��,w�:��O����tȊ��!O��G�=��v��2����L����\�hи�*�K�e��'9sy��ԉ%��e����D���xC^�B�mͿ8��h���Ƈ(66�V�7(��:��F*�B9xv����!Ba8����`\m�2�Dk�8���[B��4y�s�DV�h�Ë�I�%�^ɶ�fLu���Ne��V��iL�[�bt1��Ƚ�,��Aͤ�VUְ�[G�w.b�Y9Y���yS@���K�|�>���U��Q�b﶐��ZOK]+�����p��W���\L��R�k"��?zt�e參���D����SB�
y��/yy���M玅��M2�h'	����`�.o0b~�]Ԝ]�݉�x=5���=����9�}�s��i�U�us��N���&/Z��S���3�w��{C����&
(�h��� [�G��*o޸M8:gL�W��&��+�l��!���	 ��Do�u�P��_�}nT�X����>�R��I���� �@����r��[��ِV���&��=�u�S'%�ʥ�#\	B�%�U�!�9(d�k�O!��fx�VXEm�*��{^��F�+�6�{��D��7W�ql]<���~j�/W�vמ����<7!g����z�r��y��:�̑smΑ��
-���5q];�=�}>�S�簺��P�e�5��Z���q�n�Y�� ̏�师:	�
��'��
7�6�E(�Q{D��[5n�i�*��a�1+p+^�=*�gv��]!�x\���y��]�jh���=��#gg٠�T�4O�B*_�}y-���]��{-R/ؾ�Iȡiݮ��j�}�%>G�̕զ����Bp�J�We;c��i8F�i�tjoΝ[˝	�	{�*�)���nF8:��)W��y0�{�{Y��W%�߼�v!�MQ�qnc�6ڟ^h -b	��P��,z�
Ν^��X�����^����nl�;<���~�k���F>[���A9�o��'�ͣA��Ω6���Y	�h"�����ǻ��sZ*o�5U�<���`:�V�ǫ_�)�e�X�dVn���[^[t2}�l<�����>���1�@y������{���E K�A�� ���_�?6�}�m���O�O�[A�.:��woAP�ҩ,u=�Ŏuո��^p�DYLܴQ�gtյ�ׯeߺ��d�Ğ������v���S�O����O�(e��e9�
C[�@
��l�#�hIԸ�꺅�_hc=������i�+L���Mܙ3�uz�G5�;��+�����[ى���柇�TO���{�ƺ�����z2	��%8�1�nZ.a���׹{#�C��8�%#4p�t���k�;����0��ۙ^žةV�-�Z�gs�ҹ.��l��^ŘE֦<�W��ӣ�Ƅ�(���:y�3Z8UL�i<���6d���e��h�66��¯]��_�XƲ�z^5�����yV��:!�L�Jb�|tӽ�^0�Q�+�@�&�����l˱YuMz�9%N�R+B�d�4�=�m��r��m۴�X��ةDM\��z��u��DZ(s���x�YH7�N�#�b8���.�K�K0�K�{r�Vۍq@\2��!���9�,�!�[��GK�uЁ�σE��Gݎ�PZM=u��*S���ջ��	��V9����MK��	�9��@�m���.�.ʊr�\��E%۞�u<q�e�=s���[tn��gK�=N��Y��W\�ۭ�i�u����4ɐĘB^���wl_�i$Ä�	��cr�m���|��5ˎ]���Z�+�S;�}x���˳^7�է��|�7^4�v{���}��]Sޠ�M�YC�*=W�ޟkT	&�%��||v?�S}���7V{�"@LXs�DTg���sl��G\{�//�7���O�Fg�X���X��ҁ$�I,"-��ձ{��跽 ��F���f��Y�^B~��Crn��(yc� ��q(���S���ϝ��llV�m�D8}d�^�"}���^�j�C�Ѓ�TXH��g)\�<x�n0���<Wy<�� �o����Q#~u�{avV{d%J9ϧ��,����ה�ݎ�lCC^R�@|ҡ�wX7{�����!���s��o�����rUNuP�	�uN��~�7��P���y/kٞ�Wd[���"f.�Z����;��s2=�X�pl0��ϧ�I��̶�ܩ�nI⍩E��Mϻۼ[��k����6c��W�zf(3��9�����nT�r���߽my)��1bY�=f{���UnF�Ya�[�0��A/m��@�'�2v�O���+���U\��#T���=�p{�r��G�vQêp{;#�����I�Ks����z●'1b�oYˊ���]r���<��1ȍ��^R�B���segu�[j��4�y,���c2C���ӵOA��}��c=U)�G��hG>q�1
h�p��������i��OX�jߝ������)>����h@uP����{[Ctb�`���&W�+�Am�����uŀ�$�դ�γQ��`�sQ�����ҧj�t�QӲN�tѨ�
��Jj	�i�7w��5�<`�ʗri��
�B���Yq!u�iGa��e�±�+'z�|<�;&�w2��y�gK�`�+8K<38������9����"V����{�>�u.y�1n��M܋�]�UN����(��
خ�V[6�41ȥM�	~��L�St��ɫ�L�6K���{���
������4p�4'�1�U�����&��e\��wz��;Uw���늾��J��i�C�����h���e%0���$)GfT���[ml#)\�xz���|f:b�O�(���8���&v�����U�ߗj����u�������+�Q̲��i�ո�u�jE���p����.b�bC����R�;^��U����ʖ
����W̑��b���VqA'���>�\e�r,������B�����^��a����{�(�:��Q��Y��6�b�>��ً٤�Jͭ�k�����"録R�����c�MEQ^;E�2�A7Y��&�k��=��M�\�i�Z(�P�9��f��r*�cN 0nߧE
}/o��^�F���O�K]�b�آ��ϕ���{���3���N6Uյ�e�;���L��sxn��;&�^��9���'&�&6�X`sۑ8�%�����$a���_O����͚,X�� 9	�I�>�oXayК:��8���E�ʎ�K5���0Ni.�#�����	�M��p|�ulد$���F^ z��1��"~��S��U�l���=	�	"' �l�l���
�F:�E`�zk�����+Ʃ޷�.B�6�=3���N��CUm�.�3�3�k9d�4CIA��>�=���'�+9����k�O:-��;���NF��ݹ��dp�s��,���*�0�&�=���,=�D�`�8�U��GG�8��꩛��ܽjV��}Nz��%h��]T(�=U�,Wf:+#�r�Ȁ�(�D��<I���߽��[K���mz�';v������'�_�[`D%��:�w+�mz�\$ߦ=R�����N���d�$eR�;����4�v�ty�@h�� ��	�i^S��So}8:���8�-�����7$�D�mEM�i���Ʒ�{E���)-�(A��ţ�f���훛�LT��\�i���Ie���N.��� �QX�o�&j��k\Fz�"jT�V{�Eax�gn�w_(�C�h�"T ��ej��\V������ ��=�ņk�f�j�̟j�1M�i�"�]��V½y"���	n���{���p��[����<s����d�ae�϶�U澏�?Ҡ�Fߕ��sM��O1J�å/[v�]/ï|2��r&�қp�`��931~n�s��!�#(;U3#�8Rk8�U�N�}z���5��Z�u�ʋIG~�L�ڱ>WmO���]��U�k�l��C�?��o�`w7=�sO���Ws������8�jvk����("�E���y��S�4���Ji*Ow����e[�����{�K��^��)'*�ɥO�����}�nk�^k����T���Uz�����M��-�{*i����W�*��R[�j���e���@�~J�]�5� �BNz�����*5k֫�`
��~���Ë�.�c�ծ��ۙ����䡔���P��E�-;�G�����3�_������D�^��iXE�޻:�47n��j7Wf\::�P��`$�EA	��3 Ii�O��f��C�,�7�x��A\{��4yj2�+˝�2�ڵ�BL܎��O$΍���w�ӛ��@Nń�h4��ncܢ�ǒ���'L��`7i,�T�w��>���D�N	�$y�D�|�r�ܧzR~�"��Jg��\�a���1�w����}��]�l,��T4M���v$�����������5rS~��:�ӾT�K��j3M�,���7=��s�=p�ƨ��{\�[��V	�s*��V5�1T�=9#"��'���i��.*Y��[3�rs��E�v~� I]f�_��^�Wn������ǲ��e���ta�ݙF�2a�b�,�dl9w��Y뙘t��nV֚���{YFV���T� 5O��e�PQ�f��I��)�p|d�]�==����uc�ż�jm�K��g�έvD@�L�/1Z��p�筽����%�e�N�	���ɹ�N�cHMjq�J�ݎa��vXc�Dx�֋�us$�@�nM��j��z���[t�S��k'$x���x����N�n�k�#]nPN�'��s�hZ�����=WF�n�p��Zu�j��Ө i�k�@�靊�������	�,_j�����?[�/ܝ{-��:�����H��L�!�z�.�Gy�����Y+���z�n{�L�.�AI1f{ˌ�":UI=*�Ϻ�+�U���j��<���f�Nw�y�zf -�}&��7�]{;P<b
LU	���E2��s�;Vy�gHݾ�6��?�	,e" �m�`���	�K�-�i�I�)��M�O5�]*�Ѷp�q��nwk���ڡ�4�Hj�-{��j��/����=��S�.S)���=7� G����N��$��J�L�S�TMM�{�]�_���{�"=�(o��}e(ŗ�[Ff�xuV3�>�-��yo�ݳϞ�{H�|� {)?�׊l���g�U��������~����!0Jpn�+%dY"V��m�㣌^�k���ٞ5>>�	GY��z�|���Ԯ�x�/��S;
�������流xF�շPь���Ã�NC�ҠR�5��w�dM+����\f����*��FBUV�P��T�s�u2j7<\�#ML���9���u��O�;6k���
��y4��'PO*8�`Q��k�K���f<ڽ��L�ʋ����2�ǹ����i��bJ8�	R�M��QK72:��3!EF�p]U�p*Ԫ�j�6S��9�У:�ɩ2�A��h���]X�%p�pgm�֝M�u��)�R��_�wߜ��%��Y�G���w���=�N��{@%�Ch����Q�5�^���Ӝ!߻�����C��y-��y��Ikn���lPc��x:Nۖ�EơMӭ�N2�䃊.���T�X�~��Ν��UҧO� ��K��ݸzщ��:>���me�)ޞ�N0�.Ǫ��TL����fO�(�������q�(�u�*iA�{��ATOo����Ȓ=|�4��7�đ݄\�cя����w9Q%wnW���Ox��ժ�G���jL�L��{�$�ss۫��/m����x<U6&\��PpTS}T�Pf�:/�c �F�)7�N�̯D���]tZE�p������x8-�P��6쐎�[���b��{ߦ�����nwt�(r ��:K7�la9�2Z5�͟a
���"jc�
��>�3]>�7U�I�1Ԕ���7���f��D�,��FswG6�z*x���-��>���Z�;�4A��z����E@<A�I�ސg��dUF��4�������d�l�F����~�ꬩ���pI-`�D�Q��kQ1P����B�26m�A��/�7<�>|�QT�U}�j��M�۞wWl��V���u\IhWFM>�O������z��M#\���l
�}�|��6�Y���(\ɮ�(��:��;����FЄ��I�`I2naNW��+>r������{�=ź��X�E�GWhL���]s�ټ�������֣ۋ*g��#d�06�P߸��<��]�|�go�Γ��:�b�Ey��ɋ�_��+�niܤ���F�t��tב���W�:h9������vh��Os&@��d���[�s���a�¢h����/�d�&%�e�u��)]���q��f��:�F�=�*%�Tf��;"�'W�k���ߗ2�-�z�5�fdY�{ҽ=۷1v��Y������V��,�TLy>���6�`�79��6�����r&�)�y\��C�]LM^,F���He�u��c9��S�:����
t.6sD0n�C�U��S�$�(�b��z�wN���J��baX=�B]�FziyE1��+����Q�L8�f�A�1Y����Iu�	Ӿ}������g|z%�a��lZ���Rfoɠy��S�z��5��$�P��HS/���u�Z�Vn�Ң�z��k�*��ӖΎ����#����⯫�o�t�dZ�ݤ5r�����U�{�k��Ad.dO
襤������秸��	�au¯1���ގغ�<v���6�_�����f�S֏����\�r�s�*Ĭ)�\V%fB���{6j}}�p��F�"|�L]\KV�M��;��9q�H)�Rp��h���=l����O�b�*�����.��*��qT��ԕj�v�0&X9t�l���Yp���VԡQ������Z#��Ԧ])46�/�"*G:��e�F�Ae�w0;��
�\�}L5�p���K��4g=P���<B��]���n����2f����W��k�qY1)#T$�1@+��
��h!d������:��5)\ݜ�0�ip��ٺ�b�sc�����/��(%6l�b �I����u"(��_��y�,έ�{����X�V:�`�9��x�ڃ �4��mNSr�M�*R��8-�/�ʰ���n1u�`����Z5��V��gr�Z�j�`[�c�R�b�ǔ������1U�m�Ʋ���R�ԮuhAU��껠���3a���������x��u��Ab�l<*�[�sD̀RML/� ��q�����/���`9A���P�bMQ�C.�y
U1�z�f���{D�j�$�׽�.����n��2��վ��\����H���$���ԥP�CX�΃�&N�V�w-�����_v\��h���I�&�uӝ�:�{C��P��'6�,���{�
���/��B7��;b�U�):}��0��I�5oP�g�5֥���H۸33ke ���JM����	U���̷�Z�{�� ��;D�̠���gǻ��g�kE��W�ެ
�	ZY��q�iӠ(�S*�v���ȝ�'G����M��ڰ�8���k��R�w�*I՘.�N�sk�3׹(Z���%/ U5ee�j[��?��L��D���I��m,ԸhU3~�K�A���r[i�{y*�P�4��~��ߍi����Ǯl������l�)��4��M�?��z��<]V�c�Pڭ��ٽ��+���)����5���N4�g��&H�K6"WvMzO
�T�V,S��ƈ�f��-&I#�I�C� �P\$��))ȁ���g�e.�ţ%�ׯu����7�oz�����mFd{!�� �n�=g2�̟��MS�#(�+�VN����&IaCJ�
4N�RmU��dۤR�J��cGH�F5ȋ����Qp�2�48܉v�9���[�R�v�����:"+��撚�R��'��~�g�U�nˊޭ��sI��A�&y`�=w�r��L{9q*���n�q^59�r3:���p��*�<�ޛDIh����>k�Z>��w�{gh��eߝ"��H����E(�����v�^5W�ʔά��[��S��n'��˶l1YW�{6 ҵ2P`�p�> �Y)R�i{*�T�{OU��jMn#YX��nm�v���V ��l���/�/�±y˪5'[��U��ݽt��G����$Ƭҧ�=o.�v%rjML'�jX�t?h�Už�:X)g|K��IU|9LM{6�a��,t.5�4P��@0���r�x-��ژ"�oms���PΨ��ܝ�:������\KyVGM�N�g]�_j|.�~�q���i�	5۵����	w<�sg����TytU���eN�|�R�]�綥�^��:�n5r�;�X�s��g�\��g�ل��k��${c�i�b훡��3����>��Ky:3��;�h-�=ic%��S�k�{{Z懷]��K�:�Qlu���r�H�R�m�A:�sֺb���Ou�Θy�;A7n^��P;����"\/� o}3��n��=�I]�#���'�o
�U�#N9�NKQ3/����J�{��~	��(4PE�_I,`������?��<�9��UCL/z'�ʸ,s��oH�/b�g��l��vyB���8yc�����Nd��5��ʒb�/'��窹N�lĘ	P�=�v���L }��n�\(9��^^N���mq>$�Lu�*��Y�͋���Muګ�ZΪ��B%@ `�����g���з���Q�w����s,Ͻ��/9��~\��r���b��}'�Iv'�F�8���72��n�A��i�b�)i]�$��;��̟�c�iU���oa�ou�S�X���t���=7�N_�㗅Lun]� ���Q���}�\Ͻ���4چ�5Y��'1p�\w��H�=Lǲ1���q8�J�wt{�]7gp���{Y�z\8��A�K�mj=8r�q��S9��LϷ;�NP���99��|M��*'�ثxm���7
4od9C���>��/!Gf��?WL����{�ɼ�!k�<v4͟�!����`���װ�펶9���Ȁ��Z$Uj�{O��)T=�J���ۙ�T��r�w�[0o8��)�1pVjy�i��oa��d��Cـ���TM�-M:Pi��7h���sz
���;�]
�k
���1�̮�۝�m�qo>KN��,P���@�׆׬~x��owYHx%-�<�����ͅ�Cd�[E�ߖg'��כ[wIoH��nP4�W�>�g�(�UxX�
�s�S��4�#����%���v��Y�ԆF��j�2�wwq��yb��y<>�C��,��"`���Mnv;�gV�<��������@OU��^e����A �)'t�Nk���b�ݽ����0.��T�������b����/�=�CަC��I�m�p�M+}�v�R��W��\5AI�(+���v��]�Q�j�Y��]�*��7Y>��뭂�`�C�]|��zz�x�kM����4룳�a��Tׯ9mH��#ԩ��3,�͎`qI��M�$�P�G�v�s.�q�qM���\o�?I�.*n�Ϧ:5M����Ĭ�0�3z�D�O/�%�[��J�; �{1ʢ;W��M���Q��
I6�M;&��p����w��,�:�N��
�e�I�ڏx\���F4��]�Ł�9��5� �d{�1>�;��Iܚ�M�5����۴�GlT�#�ؗ#�N�x��b��9>��7x#����^X�w�6�q8��q��q�l��z��
ᢆ�������k������V�ٽcP�G��}3V���v��x��%B{�\����z1V��="�0
s��w
� $��s�EӻKFuq��^]��Z�U�Ⱥ�(���oy�/���:�Q�ƴ"�A����x�#XZ�\��(=�a�I�������]jWN��
�O���lT���nG�w]pm�������Ώaw���sd��oqbj�>�}�r=�D؆7�5��y����lgad
�|���}����٥����m?V�_ndb���˶|�N��I�+��]:�&Ҵ�deN�>v}���6�7՞*2t�u^I�P�15��&��j\�p���@a�$��7�P5[<*�Ge��|���Jr����ќ�[�������ۄwzs�>M_�h�wg��W#t�����ڻ�{����f���NvW^i�<`|��؟���쩯x��&A�^�����9�3P�{qv=����v�zh���R
a/�~��b�;��S<��M�*�\
G��s��~��/PY�5�`�CM����:�:s�8�q�=����vO�Lr����ʀ��ڜ#����k��֋<3mI�h�r4�s�M�6�EoM.��[wu�":�Ұم
0������Ǚ��I"�U=~͉�Nr��X���Rдv�LƮ�[����O@H��C,�j^Af3��J�m�*25�ک�1gb��v*ui[��LhK&��ZM��5�\�V����)^㎼bߚ�3�/{�T����P7�9�H��W(��q2 r>�a��}�S��*KS)�X.��	�x�?!�2�Lǔ��ܐ�V�����{6��ꭋ��ʵy��	&�y��NG�ޣûZg{�~�0��ὲw�{��|Z�l��.k4��,���:�/�r_��if���F��E�l�F��B�ќ��@����}�1:��waɿ]���/��W+#׫��NCg}�WS$ܗ�(����PN�o��_�q�2ZE�j��&đ�b���y�}�o�o%3�]���Q�5ٞSN�!�;���6����۶�פ��#~�=6D���Y�X�>:� �R]3��ЁE R@��}�UK��Mo��%̃��1������~�~����]��PQ�m��nm���[���kG�.9B�
��F"=��]���:����P+��]�>}6�0��(Vz������[��=�P�SY�y�����c��	��NF��F�ME��Rq�z=X����SO݄����f��:eߝy5;;(�t�Vx�j9;�[L���2~�@x����G=��\�h� �_eB=�W.z�v�J�Z���<�*%i;�Zzn������LX���<pv��僪�շ�
Jw5HՐ�X������{p
ϷN����%�G
�K������U`��������U�ۏ����ܱs���)�ʢ���*�r�S{��X��˴�.�`1i�C�����/qʶ�n����p�9y�jB�i�Fc�p�/���-���)�Z��m�U�����p{lG3ػi�\��uˑ���ϜU-�W4<����N�m�2vMۖ�8<`��\�<V���z�mټx������Ts�\-*������gn���70U�s����%݀�;� )�vW]������.=kU �Y�=L\u�9y����Q���u��I9�M��rX�O8S��k���܃�9��4�G��]H�V�����?��٦C��%��}s|c&�o�d+���y��BV���'��~��ޭTʗ����Av��)��������W��p�M����o�#�^$#2Q� Y���p���O=��UL���i����u[3}4�M�P�x�&ꦻ+=�%ߧFn��T��~i�7`���8T�TT�)Ym@膋a%�]yv�Yy)����݅娹E�����_�Є��$X��&��_
䦏+��C�\�6�2��l�ܽ�|.k)z�ǷA#���,ߚ���|�>�^�څy�����a����1&�VV!�cJ���_N���n���F�}����]u�g��
��	�Mr�w�O�	z�&�-SK��Y���p)�f{޻-,���q���g�lhp8��^��^�ը7OgM����(������j�h�gq��$R%Äaz���ʙ��g}�JKͭ���,���e�Wު�/R���)]Ro+�_t���2g7�Q9gM����7s�)�Cd�����%w�G �#���J�m��+�3ٱF��]e����R���\2}���<��2�C�����0�/u$I�PqJu��1tC��&�+�U�Ի:��*��̤>}�8�X����]r�{y��9�����(�Uj��F)��?��X�r��]��|O�l:�=i�{��J�/Q�P�����4�}��BI5����i�&=r�.]]���72�O*0e6��G�$!�j��鹔fэn춹��l�vg�ʼ�+��n��a��v�nOv���r]�f۞�K=&��XM�)ު��=g-�D���{�,A%l�^���΁���$���#C�^�!���z�e#�>H~[��c7��tQ�o��º�[�X;&��,�3��H,b�3�����gAQ����c:`�Y��Uд/o*�ƶϲp�w�յ�-ϩs:'H�5]~���.�ܐ��7���C6u�<+=��5,8F����Nw<��	�Ç
ckqf��G�U�-$	﷔��54��(�SU���ׅ]D���~4��}]���|�d)�[}��|=�4��I��0s7j��26Q3}�k2'Þ{�:�O�{q։R�$6{�n7 �y��[���d��%�7�b����V�}�x�h㨗�v�N_{�x�{	8aCh�H����NU��Z�tթ����Ӛ��)ɍ�t�1�.cwj��gV���ѱ�k-�:3���z�Nwn�L�2�����ꑜzm��tt����%-(�ҡz����3��M<��L;>�Be)Qˬ�r�{�Q�}�͏���؈�l�*w1S�K0)�������]go_j�7+��w����{����l�ףw�!���Ƣ��l����7�U�{S�5�U��N"��p��+���>5��;��yDϢ���iQ�Ig�7fd��o��Ѩ�4�/f�.ם� do|�*
m�J.͍�ާMg�C�S�YCt���^<�:4Q6�7�p���5�3R��7W��;0�w�bV�5�G��R2Nzn}S;�n�Eᖡ��Z����69=w68W��Z�)�e��g�}�~>:��g�:�������=��T�o������ޮfqR�`�� Vs�`�)^]�;�����h�Kd�b�����ySb�*r�/}��d�5�I4S�Y2�}���g�/����k��q�%O�z�uxi��1���RQ���_���FKGr�����3��XG�n��pZ��9'�	W~�0x{7�L�[�tԤ���	��i��̕�F=c�a�i�t/V�<pY��2۷<�(m��+�y�g��0����*���Gk�����0��A��$�N9�]���Sk��y��s�Ν�b��2��$�Y~�ō�K�6}sGF�L��Z/�q@���ċ�,&M1�C�RՑPm>4�S=+访yY�ƽ*X���r�Vu����M" ���)ϵ�~<�������w%�|J	��Q��J��pPv� �;e�l�U����t�b ����>�۬�Cs��l޾����EΗ�Џ�*���ԦǨ���}i4�Q��W�FHR&{QWyq�NL�U��/���3�L,}FF�W�B�P@�"��\o�P���wt�)^[Np��rD����T�#}*xv��x'R��=��Z:��4W??�x�`����Z���W~��x�������Uv����c^cwt�������>��n	 ���S��y#�{(ke���{7��~"���Oo�scROו�u�P�¼Hk���e�tWpI*"k̭n�_�>w9����G.��vК�Aq�7�Lz��uiY�nL��ͣ< l�i�Vvwۨ�=�Ϛ!�
�$%���w����u��P����_rY��&mp�{zܱ�hό�)Z�[��-�܍x�߬Ӭ����p��`�
���#p���U�K����y�����\{���J����fGmG<�!�s"����}M�ʒ�z��ˇ=���,� �`�*����nP��5������S	��1{�ũ���r�F�@���/{{0��5"���Ư�T��qu�t�S�<Ln�=u�>
c��-m�YթGB!GC%21�hn��ҫ�0~�t�rI���o�1����@3��拐�սr��os+C��[��q&g<t(���D����y%"1��ݍf�p�kMX�u�aY7���6�9#����wg�W����D6vk]��-�
,��j���,�ut���Ț�zÎx]��u���E�Y��T���Dp��nwq��Σ��<Y���v<�Yn��] T�l�c�bz��Q7f�۬\G4��Y���3rC�5���$.�nU8s>��v�L+A�{T�M�㗎�+�r;X5����k\�^F�py�U띷o�:Jv� �������9��}������)�__B����E�`	A%�O�H�e�Is���o2E.��M���+q�ԕ}[��4��@z�*�
�+�Ь(e���&����������]y`�\=���.��
�`��,`��waT�NtmJ�����뚉;�S\�a6�H-Ä�wnïe(%�{G	[Љ�Uڭl�r�-¶ܢA��NO�y]ux�6L��5.V���r�X�~�N���)��-t��V����JZ�&߭u�5�	�`��A�S���+Mxڨy~�t��~v;�zL�D�7Ƃ�B��Q�9�k >�G�~�N>��P��S��xp� )���t����n
E�����ޔ3w_Nuz���Ñ�3��r��1��fڃ�P�>�~��/�&�q�i�oD�u8�f�x��d��sW�ҭ饾�ǀ)�A7k�%�b�5Wn��:�;ԍ�M��e�9~��n{������$r��ᡉ,��ǩ�^l��Yo���{AB�9��^�\2�I�&�>��x�-oc'�,��63C�U���1��FH�SU^��k��v��i��4U���h@���m�<���V�̠5,���]����[&��:�a9J��z���q�V�͖w���+�3�4�c��\VSS�����7Cob5|�oh�6�F���W��s��cZ��]���v��eG(G d��1/�$<Λcd�v�u ��;���<vX��x٠����	S2A\h���c�V�78�������o�F}�1aV\�v��w�oeKg+0� B�0�sY��VPa�P���\l��[Q���LR���`�/I����tIp�Y�E��r���m�Տz9���R��˖��é���V�3�fKmm�[�Y'
�4]�L^{IwY�Y��W�7ZZ��Öf\��ק5��f�f�ܘ�:ݶ��0!�:���>m1Ef^��FfG�F�iJ���Bhq��Ȼ����(:ɉ֮5��j�ە��r����޷�����jh}�x�J֞�dW3]�}y��o��9T92*f�}�Gk0v��[$�;�%l��w T����PO{e��>x�h΍`�����G0�5QC	��jS�a!A�u�\弌ਛH�=uj��'.�8n���EӒ�k��QE�Ω�k��KlZ� w����Xf�W������V�K(���^F{��(n.��Q�t���Wb�G��M�;b� �R�j4m`����cf��p�ܮgT������˶,ڗs	���r\ǔc��Ag�R:���AM��ȅ�������4�;��:X�'z(s��l��;�n2������5Q�)6��Ym���*�*�K�f[yj��v�6�u\f�dMm�q���t��'�W�(�◕Þ�91m��k7�`��t=
�'����\[/�r����x�[�N����:8��K�.�\���Jϳ�밄�Ź�<8x����t��Z�u���>O32�8�1���xʻ���y��\����xv��Pu�lv/7�!\Xs�Y�ഽ���ݼ.�r�OI�8����9\u�.��p���^s��R�; \&抛ߖ�?}��=���n��wc�.���ɗ-���V9>>b�vs[W�.��a�<��{s��m&�^���iW����Ev��sԑG��s�^�:s�v���嶞��u�L�v��j^�-���Ż^�c�F.���,=�n5��<9��4�9��A�AژN\<�{qi��ϰs.�����[���C�����^������v���<�۟5Lp���	7{��gv��^v��[�u�ru�\���;h]�c��On8ѳ����&�q$]�y�@�l��*��;/63��֟N�T�n����{so��|w¶}C��+��7R��ye�5{�Dv�i�mk�օ�#�n��S�/��}���.ޡs��� ��5�gr�	�z���՝ǲui9��1aD4�cN|�{]K�Wi��	�M�Gn���vݺkk۞�W���mQtt�Oh�SJ�sKv�n�nD�D�s�L';���˗���\x��ZB�[���z�a3�mG-x�Z��]���l��z��Wa�z�{�k����bn*Ѯ9������b^�;�nΧ��']r7f->�ۡ��\g����ۚ�h��{v�u>��ˣ�{����D��7YP섃je�:�X�y9�3�pZg�g���],[�y�LKѽ��\-�8ݴ/^���x�^*Ǭ��l]v{E��؅���t ������u��On1�A�/^��Y����҃_neS��*�ۮڽu�2q��v�n�C��W��,�����L<��������ϊƻ����i�Rv��� ��A��']r:�Y:|�+�x�=L�}��ؘ�¼�mkz��m�ؚ�VF�d,J������|�H��޺^��|�I � ��N%���;wT����5+��lh(��3]]�.���8Ui�υ*-�h�ގR=�`r<&z\���iT�O��|PY�5���)H�o����o���eP�f�NϷ'���{�L��t�Q0+io�����Jx�b�8p[D��}恦#T��RS7�5� Uw��`�]�
�~�����!L�kXz:k��=|�d�b�O���
�A�]�de���'$߹=��z����N"A�b��Z���p��������>����TN�{�5��y������=Y]SX�|_����7UM�u�s���%�M1
\�E�6��Ǧ���PZګȞ�����z���6e���]��O���w���'�Rd��UvF_��,W;���$O��y]�kՒg��U^��@� ��a�"Me9��LN���+��2���s����	��?.���eA`
@��k�Wv����Ŏ����(C1�ˇ ��!6T,�ޮ�-h�&������ ��oj]u�{����[�
����q�8k�AT�\��
�*����Onߺ�{Wd.�E�r�a�" �D�fo�U�+X0�9r��%s	Fx���P�>��/}�����.:A�*���߯�;��H��Ԛg_T��F�Ih\�6*�w�����k���thN��ϳ�F��9Iu(Ӟ�����p	$�h ʹg�b��E���1zk�BUg鳚���~���v�{ ��2`X�g�`v�f)5�3"�ն�U�@�����dU��V�G����fM�PW��Įs5ֺ,�5��}�.�p��
}��Gw�r�t�h�5ҋ O�z}[o��984�>��׫[��)�������f0�wj|�Fl���a��	)~z<h6J�QDJ����(��mr��ۻ4lI��r�S�ՆTq"�����$�}i�sI��THxQ$ו�m��}�C74�����*�εA�}.�yܷ�<��><���f|�~_nn]0�C"其�b.I8C��{:jԷ)��ŲD6
(g��#=��=�sW'`����.�+�m�|j�[}Kت�2�-=\:=�ȯN�:�s�[N+ۧC�Kl ������1p�Y����^}'���>�f���˪Üp+��*��4��Q!
��۾���.C
���ݗTkٛS@�i�[@�0|�ȭ�����jru�[W�F�����`���v���+{F���w�3��˓C��컸5�=�u�h|)��Κ�n�ҕq6d�9u�;*檉�.sk��j�+;z�$baW��C������%�h� T;Y�Õ�|s�Q��i�����|uO�&{ٙ���3�a�l�x᭎�~��]o����v��YN�I%���ܑ=0���Ya��B��_��.���/(��#�'x��(Y�R���#�Q�ǁе|�e6�:`H��Ǫlo��S��Gz��x{�%�_Vi�y���"s֞�'4�z�ӂ\i��k�3�=�'O�qq�[��������df�=��'�/ Uuu�
��I�tDQ;�����-�7�!&Yl���P,�$;��G3��6�W��$��H�d�ʘe#L�o���M�ĕ��s�w�W$�(ǫ����j��4�:9��q"|Q��3�1��C��Y�3�쀂Bl�Zh ��Q>��j}�n,U`��
Әo7/��z��)�~��f�}�2߲V��47<��O����>����'��j#�0 lYʫ{�������^R�X$d^糒�բ��meakk��z*@��
ow��*���)��fH}�t	ۏ1�+���F�^���w�00��CM�G�)��zr�N�D�	Xb�X�3}ߐ�cg��~��������>�;�o ��,|,�,/C�,��U^����_�zq'�`��b*&p%��`�I��S��fp�������d��պ۞� �}�.nC�Ӎ�s�k����K���uNm���ʚݸs�`�;I�z���c�O���h�:3�t:8ť��Z�k8�p׎kԻziW33�ƨ�n�9��5�v�ys��]�]w�5�=��bG;���w��[�NDѭxV��E�He0k:d��[�KK���5V��ΰ=A��N��8:#��^�Oamq���Ǌ���3��ݵ6�of�τ����t{=��� 1BpB �藝!�#g�篢��N{HR����c�N��*��)ŋ9���YܞگY�9���P��I;|=�cx>��S���J�7�Q9���3F���JM���cR�p�N�O�:(G�hw]NB������5���k�x�͍��v76�'3�,t�5���E�q<u}�h��o;�I�au(�ᕔ�\}Π"��Z�^�k�2O��]yyy�$Ǘ�f�
)��`� }���Vk�͹2����p�z��C���p�,b*�h�n�u�8=�E.�a�G4�)�z�O��鬕�KI��������"Y�&	a��8)�4�yv^�:뗽�o;R��ꐏN߬k��Z0)�i�0"���v��wݻ�xTf��U��(��4�{>ߵ�d2�@�d`��饼wo3'ψ��o�y L�ş�q_�Nr2�$�'fk�B��>'bV�6�٪�h�^�:}�/�����
d�	��3e����<A���#�y�ݗ^�$P��Sit�l�E��ض�'`�}�wG�^����eM�ȝ���m#
h�[�CF�ߥch�2�~�mm������u���1<�ƞ�ufQ�1�}����c��a�Z3M�D+�'��&|=��{:�3���(�IP+Õ�1m,H%�mH�/K�����z��W��7 �_X^�aKE8`��jd���vvd�z2�sٶ7a�[A7�L��:}���t`�1u�ǽ5;�e�[ೊ����NPI�FU�vMM͞%���H���KXECj�F�ѹ�JN��x0�\�S�Gۓ4z3�3��<�QI|pM�C�'rL�UWҧ���-X�9���ٱ^�c��P��^�;[�~�wwy��	B�ඇ�Gb`�산U惱�:}�̟+I�Y���b�:�z0��G���
70M5=Q�]o�4bk��8�0��H��S֧"q��Ka�!�Ĳ@��@ǋwV�8���my	��D�u�ɑ�ax"��W�猣�o�(Y�8�Wی��͒$_#&�д9/�=�k}���2�
Q�t�G��UO�y\�Ku{�1:��/fzk�]/ee�������3Z��ߵ����7Z���c�k���&�nod��r%�<�ApcV��=�h��2#�a'
$NW$�ܙ�w&��os/g�O��\�EYU������|��|��YJ�շ���V�M2�Ol�񳚹cq�`�4�Lo���dZeX��k��X���-�^m�d��,Y�]��>�M�!tg���<&��%�v|��KL���"�{>2���roV��e'�yu���[�8u�1��|%�K���:?i["[��?w <E���3.���k���z�b.�h�'k����£��Q˜UgZ�)KoӨ^�EP����xX<֎�O��}.�oW���Zh2!�Sp}���Nm�ʫjf<|D� �{z3>L��]��t���lrNǽ9K�]�u�q+�Y�9�[���ٳYd�3~TZ�R��*��y�I�D�2��^���N�[�ݳ�|O�Dږs��W�H�.�f�{�$�����q��Eu7��)�^�����u����B���{�{pi�%�l�aO�TL
��ʗ��O�@�*��)�|O�Z6��Pf���{�h>�����]w�Fߓ�����=�!k�J�q}52��9�*��f�{y��L����Q�D�Y������DQdܿT�r��?}�]z"zm�:�Wrdx�r0��C�C�n8�̦
)8&d3	�c=G�ݡ7-gR����\_��E�K̆s�6����I��)e	4�s��=�����n:1����ʄ�|�����>��t,��C�Kԓ��9��y���źy,���{[&2�f�V*A��ugxVO)�������wU=cw�)"C��>5=y��&��n.͗Ӆ_�s��ƃ�	��Eܱ��.�(XC7��h׵dk9�J7F�a���l[y�![� �s�MŜ��0��x-UM��Rqsyfz��G8�8ϸIu
���W��P�����xΛ����ښ��1Q�p��k � |��-�~e2�.)j�q�Y�Uekt�1�x�;=��y�̨k^��ˆ_�Uɯְd�����g��G�(���M��I��]T�{��x�`eм6�G}�����t���2#�~�wd6����&��n�N���o�a��<�����������6"�zo$Z��l���{�n^��a���Qh��a�4Ϳ�?���إ�����g�u��_�/�քxYca2���["B����{3yS�/Vz��k��	�a�	�!P2{��\M*9�q(�Z:�O4o��8���_��l�\p�
��(���F�qy*����o<F�(2[J}�6���.����|�g[�|0�fgMW�^�l\�Nй�T/�����z�@�^c���y������R��,�e�a]ԝ>��'��և-��bp�}���8�E�}����#��;ƽq-�Q0�����z&�̪�ṷ��#ܦ��!
�q�ωɇ�.޿PΉ�Ne����'b[���%x휐\w-&{=q7c������+(�v.S�XM1�:�jA���Βp���Q�쎢ꦯ������勺�ei��;t�^t�G�v
���w�B>>��%��Uv�$O-s	�}q��n8wkex˹y�[m<��;2of�f�0q�:��;i�Ok�A@�@⣭��p�9�z�ݬ)�&l�y�J�=�l�pn�xϕ�c�����^7��� G��{mt�8=7f;.yl�Z�3�<�����[�^
��-YY��]\�F���aZ4�H���w]�8��2�G{c\؜+�:���@A�Є�Ԍ�+q��Y���j�j�?z�ԇܨX|��L�S�4N{P�h2He��(�Q�9� wѵ�����9�Cfܞ�����SǕa��Q�f������ӫ|j�h܎{TB�$2����1�[�͑�i����
��:^|����W�;��	Z���-w��k���岞A&g��R{���7��5u��j�+[���jpr����7l�]����v�mV�H�$�IA`�)�ǷuQʧ�:mt3��T}}w*�Չ�3'D�:�����&_t�Bf�.w�|�8���h�ð��$T�+�5���WT�p�� ex7�z���(��[��Nr��)�i1�"J�� {���B�<�$mqTg���!
�R{�U7ݠ��Cd�l"ݒG����������LW��mmz�6�N�5�) j]�}U\�i��8g���4��wu���r��&f�Q�Q�ͬ;v��i�e$m�8�ͥ����e�uR<`ܥ��S���ǚ��&A^�)�YG����*s1<Q^�c�6B��}��	��[I+�u9k��\�o�6�(�-�H&���'��X��.S���G���[ڙ�F���wQaxv�����ygTW��9}�0m��)���Uב�^��&#َ&�\�t���o�7��ù3��11���w���sl]^��2��=�}v�r*��g@2���*ܙ/E���ܬ�ʐ����!�ӆ����zn�_����{��=U>�U�1B�THǫ���.ú.׭�6 ��[�C��m]��p9��VM�9���{Ҵxeh���:�ͺ˞<=/N�i�t���o:����8��~�j}WH����@P�0�>l�I���Ո3�}'�tZ#��}1N�Mr�o�ؚ��s:��=�z��S=.3�:�j��u���G[�FA��r���.(�&e�	xS�p�.�s���7X'�_u�{'�R<�c�e�/����)���{� �7���zssW1�"��x�*��H����Q0�6ItY�UR�ߨa�5qk s-��ե��̕�pE�o��.K8����M�ͮc�	�q����)��^R\{e'��Qu�僔2���/n����<��B��Jn�d�=r���V�o�Q��G���"}���ڳfQMXuqU�r(B�9"�*��s�n}O<��W3��M��`��7|˂��i�o���e{\ug�b���NY�GJ�����QB)8X�2����TL!�݁ڛ����Q��B@��D�=���E­�3���7��� 4��"����ժ����(�k渁�=2�l�X���]�X}-��Z��kB�/ozTI3�o|۔o�����e%R�����H,v6���Ƨ'֭w�|w�Bz�{	��<z�d��nk=���48H�|�+���g9��k/de���杪��H7�jVw+��|"��L���{.}|d��GG$`��*i\��,#�w�yd�E�_f�I�����,?�?_z����ptQ��/�9Z���Iꪸ���U����v�PX�������N�I�.(��k\��0#izU�2�^c�^��57��؟.=y=_u�ٛm�g���Lc3R�HU�ݣ�a}ޣ����wWn�:��@?��H���8�^x;�G$z���n����<?3/�I�,+ӷWʀݩ/|w���W*���x�����
�Z�'CIRo`�yR��0��v�m��Lm��M�Kގ+	��e��.]zUX[����\�����S��^���YT�Zz�O\9���ǘ�L�&��M����cC���uˣ���Ǎ����zu���^+�^�U�GM`�;�n^mE+�u�B%��v��%b�]��j� 2=����;f�WRv�V��<�D ��xZSs�Ĭ�g(�������K�^5ϊmǶ�('q�<��Ae��p3	K/�Í��'��/�����$F��A��ǎ�ꍧ���엇5�n�;��GKXP�'�ν&�Ֆ~�R�%Ҙ�x�uvf kF��:vC����H���Mܛ��q�:ViO�tN��f��I�x�Y��'26$D���]�j���f��`]zMM���w��%�r���(���y����8�<*�j;I����	��zVs�{�q�e���o7)����4]hHe�F��܍E�q4����ղ��T뾃��m�Y�z�E��T���[�*j��cUݛ���,oN���v0�j4�1�B��o%`���z.κ5�_s�4p���z� �C1���](�S��ޛ��o�X�t�N�;n��h� [H��X�3�9oa�^𵶖���7�%ɲ�y��ŸL�s+9$ɫ�*�76�u�S ��R�9`s%��h|0�滋�^�*�u��[cu�a�p�ET�m�8�8?x�1$��U�bB�7*�%�e�#Mo�Z��k{�]cs�V�OS��a�f�mK��a�=������,�nƪ�'J�eZt�����J�;���sHym�IV�J�xU��V�zB���sS�P�Og�p�	�����
�l��ڟ�}=�d�f]o^�U����M?C�;nڲ��Z����۔�op�Q�L+��ء��i���o+�.�c1�8�)�w�JD�dB���B[��g�3�q�,��\�#j:�j����N��jV�0�Da�(�-�4o��Lf&V�7��n�C�Go�'7���7�Pw����I|�캏���=�C#�;�z'�ټ��|(r�<����l\*�bM���ul���ђ*�p>�4%ƅ��dE
ó��	��$��0 �	��,T�����9�����s���EE�,&f�ݝ����q�IiOf�4��%������k�m��k�צN����h�d�O)���7�Lm>�/B>V�'��,�0�K�����gW`;s\µ~����(y��C��
턤k~��[[������i�/ޞ����B)f8n@�2u-��s���po��\�{!m�{\OE4���֌=M�m=��'�5�7a�\�l���s����"(n�ݪ��帱ж���9[~;4,Ĭ*����S�m����b��7�'o��?U�Ev	I�[L���V���^�>C�(*}��Bv{D���h�<Wd�kں�:�#UU]���]�;� �K�<f�QԲ�<O]�{���
;"�� W8\2}�[�_^�-��������W��=<*��Qw�gx���g-ù*2��;6����A�tf��b�9�\����r �	>�3*aw�j]/P���E\�5A��U�kǮt�o2_��5�豔t��L��",�7HxVyz���V���O�*P��	�Yo�kTNګ���Vi]f�unC�/���L�UUY�Xrkm]��tU�p�%ܸ�*x�>�rJ���º�n<�Q�[E�Q�:r.�IҒZ�;�ۏA듂w\Z��h�G�{a��"V)MQf:��X���7��wAƳ��N��Hc�؎���w����s��eo8�Uq��qr6����V˭[�>un�����%{O���d����m�u�9�7;��
x�,A��f�穃fD�:�^1����>��&2�!Ԝ���1=� b��&@�a�5S3?^��9�*�kyO?:W�*�ω��� ����u�O���b��nNo��t�t�e����R�	處S��{r�W{)t!��y�HL6�`�C,�oԲ������0-E�仴�����Q���3	]-Ebm��z�;�˱v�n�wY��Cf
m(p
�)ÄQY �vlJ�g���\��EG�I+ͺ��d���z���'���>�����H턔�SƫS�R���Wۯ:�=�bìעvs���\ii><��燠v�>�g�.�����9g�%g���w�.^D���!�P��L��3T ^:n��*A��+����+�_�\ԍ�Q�V�=C�^U������ߔ�xw��5�Z�4O���2/�;=&�dܙ�^�3��
��,���g����9��Oh��W5��U�uB/��S�
rt�5v;�9�w�=�u��~��7Y��8�y�o6�{�O�b�d4�m����p5g6w�yL�>�>�ju����U�lN��n{�:Cq�*{�GA2={]y�6Z�97��b�
y2�z]�ތȠ�j�u�j�
�gPw��,��s�d�5�kw����)��ov��olT���&gzdS1�ޟS����&L0!`8&���+('�ؼ�B�5�\�^t'�M0c��0�a��woX�'��INv��hi��e��#Q�&Ҡ�Z����D��c�e�Q���Kݞ`�)%H����_ws�.g�q��q�l�`黼���A��ul	�AP���Ɗ�^�r������,l,n?Oy����f�����Â��c|9x��\;3�����(���MNu�lUG�bHl.du܎C���1�Lۘ��*���t�k����_�N�(�fmK�9�Փ��X��N��&֏J�b�eCWF{y������Ϋ�ѧ\%��?�qZnp���Yi͑\��̢kZ�=���)p���H��j�.nw�Y�*�v)i>�VTK	�p�}&��i���y՞�}��-@��(�v9���Ƨ��|���yR�}7��u��-��W�TUX�V}]�~���R���If�d�s�1���קۘ�{�MXM�'��\��Ή��C@
����A�M9�bN���՝��{$��3+s*��@�RZ-"H��;'���̼�%G`�����5��1��dzj0��n�P&Y�lV������{�fʓH��^�Ȭ��o�`�R�立Vv՝��F��s.�k륙�KF��6�`�����Md\E	��
�g��2X��u@*�;�ݞ�[�c��L(%��LZ�~b�G������}��Dw������T�*ߥ;6H�&O��)��]G� zpMrZ.���r��9^�Š��Re�*zu�)4=컥&��#2���1�C;kdi�]���+��q+���~U���k��U7�：���v�K��=��/����a=��n MBV� �������>:%���
�Yw�C�U���	~�k�x��χy�۬�����h�t/���R毷�J��2
0!^͍���97���]^:���UX�¯�y�AY^�����<�sȇ��5��Р5�MM���&�|l8Ww�n��IЯݢ'�a�
A6� �Go˰�Fs3����]-B}Ѣ��y~��6[q0c*�cM�>N.�Bɼf��&�\��\(m�$��a�Z;;w��%�'�㵢6�oªA�c@��]>�7m���Ў��-B2E���˝��͞*��lB.�yP�%ͪ���D5/��CX�@�Zg�x�b̩/���~D{m��hW_\����v�M3{��8\t�^\/��zs
oij�ˡU�~s��.��.k1ZEM[��R��V���ؖ�b�q���Yf�	n�U���v��}�g�F�J3Wa���#��/
>V����3tkN�݆�U�Uz�)V8�޵^���Q(z��~�:�C��w&�βc6�֠�9�2 l4o���O��&��D�_?�$�^��'#�_;>[5�6�n�k�8��im���(;x<25�	9�Y%L�pØ�K�ԧ2��1� ��S $_1wx�I��j�-NKA���gQ���U�(�����"s6���1��飕z#ja�ъܹ[�C�˺�bo=�3v�YXkݝ��|x�`�N�Hu�i]�Ġ���f�����;�G{�׼�*��`��n��v��@�5h�Gr�����GK�Y�v��ٍǲ�`�K�O_����*�om�+��{d�����~��Zg_&�ר����'��_s���yz땻>��J�(pF1��5�5��o��'��j��s��o4�\���������Q� J��-�>"�T�竑�֬Fӏ7�{m��$ͤ E� Ã>��Z��x�S��h�GJ��>���{�R��d��J�Μ�Wg�� ��&m��<Z�{p̚�V=+�I܎���6id�ӷ��N	$��C,ɢ#Õ	�s1W�m-2fHGmOb��Y,�]�rahGVT��WY�ιҞ�R
�2ƃ���V{T��q��r$����\u�ҳ�����|]5j�wG�$n:�X������x���A�|������5K���n���λS��\��JqŒ���ئ�=���k4��v�n�ۓI�P't��Tn7c`۞ط���θ��b̜s����u]���Yr��wgoG>��A�_)��Wr�mpu��5��m�֎ҫ']\�X�W�ɮv���:�$�;��pt�q���Y�F��0H.	l6�`%�ӽ�ɻ��үM�ޮqd��Y}�����n+��jݿ_��nr�|��1L���k� [V��W��j�����(ۃݫj��V��k�9䷤����^�sG/��Q���~������ٞfهwߖګ��(���m��qr:����d.��&�I�>W���4��84����9��&z(.7���E��s�rkG]33�)SN�<�]�ZT��q��t���3��a�=-�P�d��@^�˼��=���QРl��^7di��	jWzWx��˶g���g����k�(}��rͽ�a�&||��߅���sʷ%�V3[{�wϫ2lw�c�H�JPZP׼Gwm�Yw�_��Ɩv�rD�v;���z��1���/�Y��lr���V�@Y=��T��6��2����;ҩ�.,q(�` �n��ñ���sm��V�[��L�.7U^�;J�r��b��0��Xh�����>�$eC���p3��xo*��麡\ v���Kph�)r�����E�Uzt�&���U,��&;�qSb�9_�e.���G��zg���^��\��Ez�n?DZJ�xP����L�O4M��O�� �E���f˾��p����t2��p��]�j��buu}���k��e�&FE���_�0���-nW�~75����@|-�Ѽ&�[Auz
����.N�q�Ù�n�-�O��.�=\mF�!��L���^wwv�+d��[f'���B��Ә`�ĸ�f�6bs�C���;;�Udb�~S7�;��Д	Â�MȚ�F��^�=N�i�*�xRR��U�=�՘}�zGdl��A��\蕆&���ʸ=�6�:5 ,<�b��4+ i/�(��6�4����&��O��f���P�3ؙRu�oa����7�gG<�|����"xЮ>�ʲ�k��z���7��|v�n�ry���7s���$��L� ?�+�*�FWB���Qu�L
�:�{ Lw���7yc�H7�j�����K��Tv�7(#,���v��q��T����p'�d��B� Y���qWU[#��ťi7���~ԥ�I���ɺ08?RU�/�dy]��R^���	<(*g�Jy���$a�a�����)�Yx�_Z�kh�s�6�]k�z	��T�*�WB��u�y��S�`O6ƫ��j�
�$j�f4�bt��W���}�9}��"�9�T����Yλ�}�����m��ڃ%��ճ�Lvp�Ў3����S�X�t��l\���7�L.��*�k�g�`���Ѵ�4c�W�&�2�̋���=-܏nƕ	��$����{�.N��a������C����z�b�wh7z]h���*{r=�t�� 7n����?:��5��3������ÂI1��¸���N��ϦcӞCa���^�B�hhH9&|Mt�P�hr�X������垊����ݕU�v���y����e�pچ���ÅΌ	�wպ&Q�9JY�{��.����{2�2tz���QW5Uy��7I�����U����P2�k��;r��6��a��bk2&=�F��9�y6�y��@���4��r��o,cj��R�	.��ri<B���	.��Lf���'�	\�H��KYhCe�m�Hw�^�{�*�Y�SG�_��*��i��@��u�c��M�鮲���۔�z�v�¼��-N�S�����M>}�ߧ��*͋��.ӫ:}ƬO|��̷���F�˵J)de���4����ODƻ���[�9r<�5���zR�1s�z=�6�^"̒�gj�ƭ�����fďň]��v3?U�_�ˊ~3`��7�]x�J�S��u~[��K��\/�^
G;�6���zEz���KR�f�6%�A�m6G���&���t��+Λ3�e��Ж
����`3"�&'�5�F^X��9�;�Ѿޮ����>��(��S����GqfU+��z0sm�஽T#�}W����/ɷ:%z/�`t4�IC`5$�^;i	��RQ˨�w�n�§޹���i���p�3���U�{�R�\�/uL�ZW�V
���r���^����ڋl���&6(;ڀ3�nd��|ɗ��/�3�^���Qڼ�)���+ai!�q�j�3���}W��/��o��J����o#���f"�=+Q�U.q�C����x����y{�TŨ��l�Mm����] �냖�C�n�j=��k��=��l�T2�^ͣ���1�f�D�:
w�\S��R6�/���y�|g�F�W����
�!�՘׆�]:o=#��d"��*^��.�x��i�蓄z�㾛��/C�=��kg���=1K�����S�C#�T&����v{���r߭�Tb�aYGG�k���}Y|t�:�
$�2�M)ٙ�g�x�U`���k��}�C7ȃ��er��t�33�؞8����UI#��El��W?^5FV���#�d�~�7�^z;kn�_GwR 6QBپF}��5���g�j��
I���O\������g ��ׂ�n=ְMe�r�_��nWa�X�y���M��;כ�.�N	{e�򙎛�Ɗ���0����6|[m�ᤛw7O㮹��\�<���pu��^р޷C�<�>w�>��}l��pSZvn���NguԖݥ^��%O.�!��]�^CpnTN�{��.����Է�ŕ����H�׬p�;s���	3�(I�U��=]�q��s��r�sz��EN^�g�/Rk�gv�8�F�<s��c�X��]���cIJ�t�qW8D�(�
�*?O8��+�߿H�T�8�.����6=�.�uB_��4룏p�
E?�U>2}��>�6�V���u�&��Q2���w�\;#�5�+	���s9�О����*������lڣ�s�z9�L�l?OT=w�3�����e�p�H`�v�^NyfX�+'b�7�B����T,*����::������C��͙mT�k�Tk�vg����r��p���b�	{��Ϸv'��#�=~|��w�</ҸI��|wW1�y�*w{�P�%
	,6�*l�F�^/L��h�Hfe�n�>G�uכ�4��̃���pGa7��h�тΣư篫½q���5'b�.yRⷳa�\BpڡWK%��>�MQb��@p�g#Q��B������M��A��*������)W��=���v}r<k�.�D�[?U��h\�s��T�gs��(��� �>���;[�>�H����o�k|�H�ԁ���S�~�ݳPy�f'kz��c4�_v:��&�Z��9x���O'��&���{9v����}���׶��hn�wV��ӓ��S�2��¡ty�#ݷv���}~�[/�1�����ߍ�;��s��ַo9X��ü�K��.���E(d]�����7�Gc�"L�tR�R% "�O���U*~6�R�fr�j�Wk�SvK�]��,i�����6�lnֱ��.%'4,��j�FyP����1�wv���Z�}�,�˜�_|���:����6�&;޾�E�l�Ȅ��N�֧��sM���8��93�	�.���]w���R8q��2�v�1�VÝW]�ue�znD���k���q���3p;���n�c��*8��.���k�V8ɝ��30բ�n�&��z#��:�0Οk����^	���[JfSvo9[�p��{9N�ʫ�;T�����^��D�a��d��P�Y��S���n'��Ր����r�"��e�p���kv��͇��'�u��-�g��(��4wK���?�U7o1�vhf�"V��ǅ5�!U.�������h!���OeA��c�v#Q}�@�wW�7�c�IZ����v�>8^.(�����%7-��䵝�D�_Z|&&�nf�J��N�о��j�tn_e����f����>���U�W
�*�E%�{���(��5��D�hOx��0u����븯;Z��΂���h�6�+6(B�GP���z�m�(5��N��on�*�`�2��O��ylK3f�AN�v���dӿ}�MV��(bkQ��W0�aSwZ\��g*!D^T;�<�:�*����@HE˒s�U�/1e�L��i�v��RÖ�����ꪧkl�*���c���jwr#�'��uѸ��A0RJәH���tT��E�ݷh�;v�ۓ��==�ls��#u�QS㵻F6�"%��F$����Ʉ�յ۫Kv�{�مм����'��
oC헰=�g�'=�+v�' ��,���w.`�7��SWwG>���5����㪗�C��_N�K��.��m
���۠���s؛Ձ{.ת:9�v��F���6Cv�ug�����9��������M�n�>Z"O+dtZ�zs>�v��y��_�he9�W�m��p7pEF�c�Z�Vڮósi���1'�]���ݱ���f��n�K��dB����ܛ��z�GX�Nq�ۣ��x��kR�&6�54"´�*bj�&yؗ�q���*�Ͷ���,/���V�g��������Nm��N�>;=Lp���9�Y7<Y��)����,�j[��{ps��1G];n�Ĺ;����V7W��l�F� ��\��c;����D���;!v���8�ks�v^F�]�/-����by=v܈t�h��8�[OGNs�5��R��;[��\��n����5�s�:�à�����sKl���u����؉���׬�n�l弜N^��q֕�Z�s:R8��W���=�ڌ�HF��˓�u���W*����7C�sYA��(�b:�X����'tq�u��8���͕t�v^��-���8��4I�n�Wh%��vY;M�g�ۜ�q�4ɮݥ��m�fZMĤ�i:ǋOF��=��k�jg���7���յ����:�y_.�:�I��F�v�i��p�z�g���o�s�a槳���X�އ�q�x�7��+�Udw.�z�w%�n����Ky�Z�:����VɨA��v:}�v3���#%ݳ��j<��_|ܫ̧a7D�js�r��ay^Ve�ª�+�牭��%���:n�����&C
	��m~����O�����'�r�뻉ؾ�	�
 P�b�4Hת��u.βfL��%��\k9?~�>���5�[aeN�Dee�>|�#�/����n�Q�)�@ !4�A��n��Ǽ�j�
������u[����a�ٿ]���|,W��X���]f��o��R�GB0\d0�#n��H���.���F�/�uF*�"�Q=�2(~����(r�v�n<jn�M���p������vq�@ߎ�8h�ǏE=�Q���j���>&e�h�`ľW;�*`/HD8�E��쥧j��&���HQr Ơ�*���G��U��9�ܶ��&�!"�H�9s�rB/r�Q�c��u9�3�*��q����	��L�̈�U���S�d����k�z|�p�"O���^��;Εo{�}�Y`�N	l���Q��8�ǜ��o��κ�)x���������{��YY�+�(���9~��'��ʬ�ni�^mWf�5���^��N�Z
a�+���/<�)I���y����we��:�dzI��׶�D�Wr�����r���l�X��OV��kήq�wZX�vց$�jv��/ej�Ëi�޵Zn~�@N��������{�r���,���L�R�P�ݮb�Ɍ�{��fn��8m��k���@IR/�
��Ԇ�9o/����Ņ�ϖϤ���f�R�Dܭ�}�.^y�f���w��$��m��0�\'��eٿ*�:iod�\���P&;���'^
kٱ|��.�T��|F@�q]UG�Gp�V<U�wל�dg:b!A��D���3�j�4�5�6��E�^;ƕ��޹�r랙���F�}^����:1ltL�O��kUFrFg��A��˟b�;��	� ��$����#�[�����ma� �ˬ~8�A�{��uz�u�w�hm]?>�3Y�׽�S�*��]�PH�w��\y��M&\Y QE߄�/o����ys! ��/�n{}w;� w�93}��r��{JFa�ʿ���E�뎿a[	e�7B��������Sc< Fl�L�)��:��`�-u��nVτ 4v�^�Tt�?vQL�N�rεۂ���/h	�=8����5�w'�۲��S�'T����C����=�3e�~���>CV���m�=�ş�fgI����ת�U=уc�yKD�`��dnOT���~��^t J�'�x%=����n?�*.;��@ɃJ�q�ʧ�q}M�n9�v��,x_��#�|��G���IBp�Ͳ�;'<&���=���-�Y��A�Hҷo�R��+��P�i���M�hn�5#ٜ�C��a�E��t��^ݮD�A/���M�Z�7�qowe6��lG���bf�4����+ˆ���wNmî)�B�W�EP)�H�^�H[�Y�wn&V�t/-�>�.}دb�w>��to(	�m3�]����tW�<���}�]z�F{;���n���gU˯Ӏ�P��D{����B&��g;��X�`q旻���_��BD8!�k6[�왂A���hFc��7�a]f��x�����p�]��]���*��VR��@P��'��.�`̈́�����e߸��v��p�4E�_���M9R���z�0����C���q���O�o��@���ƬeBmLC��*Q�޻x�z=��By�v� ��ӆ�=�糲���,��Y����h Xe<�9�N{w�mr�����fs��Ib�����_	���kL8J"ZG�_��MO;</t����ev��zj�t��G#�ޙ乚|ϰ��:kԼ�[3}V������{_:ޕ[̅	Ap�,�\���UmH��t�D�_����Nw�Ng�ǒ�隊�XP�m�������휻7�c���T|����:}��O��V���/qn�@��a�uQ=�ڠ�`����w�����R�xq�h�09r�_N�n*D��7�Ϳ+�e�|[�W+��)����7Տ���[�����Ll�T������՗�9�i�!,Fbђ����ݨ>mh7�t��O�a�@w:�]q���S�����÷+�'t[bt�[���������7��B��*=��q�v��珉���6��oN睬=.˞e��9p2���h�����6�v��5s6빎K{q���ik]<�Hnͱ�WGAu�<��z�mk���zEaЍy�<=�����s��N[h�B�Sج�ҡ�e{Y�봊7lt�n�N6.z-��D�y�p;�v���7Ω�7��F��P��g5Xo=?���:���G�B.M6�}R��Y3=�	��W�^�Y$ep�њ�f���Z������S[
���+��=��̭ʝRt�^<�Φ��fs�;Pd�T6p��\�ѝ�e�fM+;�Z��L�Gmyd�Q?��~�7~s���/;ph:���(�v��t%ջ8����a� E `8-��^�6�$��Z#���$ߊ���l�@����%�J���*�7P����9"z��e{(���A���d4�>�����.��������{#�:}��,��fq�q��c˪��3kb�)�!�pm���v܎�L��1u�v����� �Ȉn�m-�cR��2�~�1�9�G��������Bv�*=�����х"���5t��ժ&��9���m��W��#�N	����Y����_�:gt��^r�;K�o����}��x_wv���U�=N���=����A�3뜞	Rs���QP8o�.�~j��w.I�!4�E�7ˑ��#��n=4f�����v�MC�{7�dx>����n���Aϧ�D�F������Z��}yE$���6���ͺ�g�:��	�w۫'f��{�aYsF"�C���%�#��h�0�')K J�:Sch�C��(�;�u���b�o��ʾE'��[x���W�v����K&��2�235��:�tsj�ѥ¬�ͲO��h����r>RaԆ���w�u�[��89���ov�N]ϳ�:.�������E�M����'��ʰ{D�EP}x����_M1�Z6<�`]}��l�W�S�{�5JMF
��Ay�>R<�=n�"�&h���Upn�x%7����R��o}$� sM&��H����:��Y�u|�k`��j3�
ºg�J�z=�DpP5��۰v�Ͻ�5�]}/Ɩ�̱�.qhۙ�M1�3�	�=��{�H�q���ٞ�e��;"Lm8©®�#����V��9���$���pS̃]��"r~9�S'Enw+m�]U�)#�K�+���� �8���^O۾���q^�;��>Oz}�i\^���b�����`�造|a�PP+��������,���>�j�Mk�r/�%��lә}����K0�5�r�w
��[FL)[�3w��ϯy˥���Ş<0��ٗK|;�pTZL#R7t,�q�+	��h�W.�C.«�q^��]�f�.���<^�3�` �������X@��ynO���C��T�;�M��i�I�vz�]@�΢�2}��&����bm*�׹a�:L��q@zx7N<�W��.���h�ԷE�x;�X��%�\Ԓm�5y-����k�}�,���T��祋��{U���uG4HȵyX��/,�����䠺w��awn�uE%�X�k�<���}�H�z&���]��f�#Ի�Y=��Y|<��o�
���<�"
a��5R��6j��/VL�n%MyIdFgiEϢ["�ܭ��4"�xe�Շ�s9�v�0���Y�Qmg�6]󴷩�Hǭz�j_��0��e��0h��V<3ՙya��l�A����8��s�ګz�rO�[�+�.g/f㸪KQ��SW҆G�)�Iķ����[��׻ <�a6Ҁ���g݆{sj9����w.s3d��d�N��ѓz;<�����ݶ��O�Ep������r�R2A<�WE4��Y��k��-0�Ό��3>ӞO!�A��d8R��s�����_�����jt���~t�����+�U^5&(H/o��a�9���9�hJ$3k��1�������޲u�E��J�M��,U-R�tJ�����n�Y�����F}�xM���iCp�p��ۤy
đ�5��LԮ��=��%q���eez4��p(�ދ�3�(��δ⊾�(�O9�s�yT�#��ƶ�ܬ�샮����p���QY�{pW�2���iV#/a�+h�z-�AD���?�����ZNZ}x���M�ۭ����V	K%�i�����n�T�<#u��;T`����ү�?O������J���j��Ro��g�uu�U�۾��?	���y��29^��"z�����ރ̆�[��mY�7�W�7�weH�(�np[Jq�v���[>#߭�=.o������'�#]a���9ӗ����8�I	罻���ڧc|���
�:D��7�X6N���W��C�g!�w��fh����d޸ʮ�m������=�mp��5��{�!�{v�'�B��H�X���6k۝��A|���03qxz������S/��8
�%��l�U�#<�^��U�`�V�𩊙]�I�qc�4�����2U���т h���,ͤ;ūV����&c�i��,�zf�Z����{�dH�f䮏dos��l7�j{���E���Y����VN��v��ݪ<`�'���.�7��5����J\�j�t}<��cTn���u]��l�S	/�V��<(7��.�I�K�o�#������^*�c�2��{y�g(��=ÜX��v��k�|9��%7�;���W���{��%ߒRL��&UD��GGC��9�?�X͐���6C�gyd{�����B�����yY��+	xü�fL�I�O��}4�.�ku�'̚�����+r����*�/p9R����j�T�g���������x3,p�����+��V5��[��vs^��[Z�k�Oó�����MOk����2����7�-��豰N���-��}�nV��ړ�/7�5��x���a<p/9�ŵ���q���:���ƭsm7O	�en�\GI<�5�����,� �����F�$�!���e��]pYMC���)أ�[�7l���v#�����n\���,Q��������
�Bux���>�Bq�\��o��o��N pRd8�]����R�<��s�W��s�]2�3�|����z�Y�>yZ���t�[e�Ҩ�HM��|s��zbg�h�ʧ(lκκܾ�"=Ó�6�)�iԇ5�;d���ҴU�ng�I�l?-��u[R�s����@5�I�d��T���������wS�Gs��a��7A0�p�Ew�J�d�*��+$�H��(7���
�3�3&}��q1��,����:�mqSy&�F,X�$��?�Ǹ�6�7H��[��CŭX��G�W*�6+���L�Ix�Z9[��-�h�@�Ϊ�`�sތ]�H�y��uW!�AnE��Z��zS�!�w�q�$�G7&��3ޙ�o�֑.�v��|�ϕ{�z���(5�s}�+z�8������l7�V�HkՖ'ѻI�m��"b@�9d��8�>7R�f�]]�`���o��U��{6m���9˩qA�W�~w��p��v�z�]Գ��+3X��4"�!����f�N�Qܪ��r=�+~۪T=��R�w��Dy��u�1���<d�O�]X�#���K�w%���wl��V��+D��	6qSsu3N��5�}�\��{�1��ML@�ۄ��u���Ij�Nsތ�7 �p�k�4kz�j��=Z�BO�k Y�D�y��7���#�!�d�-�@�����Ǜ�Mb5�����{�k�B���H� /�0��bJ��As�������C]����AY�j6��������k����8a��ux����z�9(^���%���tΫ/?j��=��Cc����}Y�2C"8M0Up�42g�"\����ө+�Y��h�ҀXH����L���bJ�Q��ޠ���J����+K�Rql��
[���NH0�>>ҙ���uz?-�nǷ�#@����9����>������'J�H�'^�a�����W�A|��9���7uV�|��7�O2EX�c=0.�ACq��:����.�]�k=oP^A�}���w��ΰ����"���{ԯ���[J�wc]�||�ޥPO�V���TV���(!�L6L �܎�0�b6NF��'�M�̏ny����'��TOٝ����j�VsZn�׵/���o�F$�3H}_+��[%�8���g�l�{��]�4�_7�aG�>5��u33�`3��:\�F�W�������ѹdZ�\r�v9������Z��x�l�\����>K�W���r!	ױ�ߦ�Me����w��C���>'��O+���ޥ#AW�^Bׅ���:W�!z�l\��WVV津X-Qh�����Ӛ�������+)֊i���ct��Q�]�aD�L��\��}w����wR= SA(p���f��0�� pe�\�,�x��jG�LWy{L��%s�~s���'`p���J��޾�&�ޕL�=�S����PL8(,���E+���竑��]��~[�{�e
�.���S��Tx�b��EE�$iҕ3����뼺�T�TZ�2L_�(���(�/���Mw� %k��D������̊��S��	6���?{+���q�2��{7J�LvD�u2n�vo+^�}�ǻ�t!Z� �z�ޟ7s�c�4MC��P���A�6N`�4�|�F2z�pb���Z	JY^~z�������l�U��
Yx ��̜5R����^��Kx�ƣ����tG�REy�#d�>����j�d��o�4])mlm7��\uEE鿖����BvP�TrK�,�$��H�
,6�N-՞�w��c.Hu$���to���>~��U��ɻ<dv!^N���+<��+�½<�֘��*6��=��y��ׄY��샟f�0z��f���c�6�"$�L�n���/w�~zGC���}����b��	/g�]'�}�L_(����M���)"�l��I;�#�����8ܼ�������>Z�C� ��dJ�Ы��-6��VmWKݦ,��0'iԷ������s
�b3E�O6o�WX
��a�/in�{-��@R+kJ����g[T���>�⯶��)�6/VK��V��'Ό��n�rg��	r�*��.|w��|�9Y7�ѹ�����0v��˛�}v¤�]��hȮ�N��i�G&)X�ȓ
�˅���wɻW�T̽����h ؠ�nܮ�i��Ʋ`_�W��wRnk���qj��!�l���`��a�N��F����<��tg_R����*S۬�፜��
�Re�љ5Ō8�9���˨�ؽ��.U�-kb��[�'hV�^�ʢ���b��n^;W�.��~�z]�;[{�n��Ρ�,�i
��Ӂ݇5�nU��[�������ZSo~�]8��B��y3k<%����`Iy��f�]��&wqˤo{(��)ɋ@²Cmܦ��m���hV`B��9E[�A̓������Q.zj�^�NIc�ݹY�{6�\�K����;0����ޫO�Q�[b^mE��Vm�Yjޏ��*Y�;��Z٤S��ٙ�����R���,vj�+�tX�Y5��M"��ӣ�TSwalh` A�r����H^�BR�߉p���R��Yr���g}'o>uCZ�\���|*�ڇ�80cf��g4?�-s׬u>�hl��-�4r1��j������%T�v���	۫��~ˢ�v�����L�uCsE�6���h���N���92%�5W���v��\W�f��4�fi�x�}�K�:<Of����yw�P�4�����2�<F-A�(&����Q:X��#��Egn�=��/ƚ�E�����E��y�Oձ��њ��^��u��F��Nr������i�؜�����h�-��!��63�|ga�x���x�q�=��r'<fX��� �o?p�'B@�xn�N��uXC5\xX~ݔMl�����'ș�"b��ڒ'6{%�����.M���}�Qg|�ښ��y��M��`����f�L�

$�E�#Z�a�����6�m�\�7�N��D�l$BN*X�>g���Z5�[ʣ+6�}�9���űG8���R�M=����(����i��]7o��+Ԫ�5-n�dW#���Q�95�*�{����2&{3�{E7�vL�qXÕ/'ϒV����Hy�o�ܯ7'�mX.r�:�޻o�ќ:[�!�e�Wú��6;��MOu��{]�U\�/���ˑ�]S>=s�hb�Өt�)1���R���~٬�G����<�I�=�dS���+�i�i�۶4H�y���o��)T�
7~��������9����.~�_�hi�h�=օ�	�I�K�;��E�P�2���{#�q�hޗO�F�ml�u�,���9Lt0��0�
.�o2�7ywF\)��s��W<{\z���B���gmĜ����jF]r��3�+~]���fM�\���l�b�B͵��q�n���s��-�q�wRI�ry�Vmډ��lv(�.�V٫��Ud|����#y�q�m��#�B�ˑ�9۳�v�0�W'M��' ��D����9�0	���p(D��s[��%�zf��{h��*����)ӝ��/5EH�����O����y����N�&���k�4��	�8@�G$�,�ɿw�GOj�]�V�_�	��=�:%���c�L��g��R����h�ܙ�=��Y�`ک�6�Wj��2����m�"�ܡl!�	8	����q3
��W*�Zjww���1cҦ#ћ��y��Vp��B���� �89�nu��2\��88&�HCh��i���H+}�/'w����SQ~��u,8�Bp�R��p�x�B�!m��Bznz����5W���Nh���B �O���lg���^�w�����c�rdd��zV��X��@��gV+�Sʼ��u������B ��ڍ��Uy��NAA	�P�B�n�V��P�]�w���V!;���=���@��wj�<ջ\�ȑ�n	���U�s�wŞ�#'���{���m{;�Б��n0���>�]�/#��VA���L��FH���_�>���As��+��B�ޜ�f����݉+���-=7�E]��8oܸT��98��('�>�|�$+�3�e�\s���3jla�uǈ�,��9�������ù�L�G�pz��iږ%�����{cϕ��3a��^�()WG�F�@�Y"�>���*V%,��u���t2 �L���5��̳�ƶx�Ԡzc�]K�='������e0I�0��VN���~��%����.T)uRo��~�I�C�ƺ���`���F�;[]�ӥ�ṁ��,�%CI
���{�aJ�)Qdej���t����T���iU��k����/B~�X�b��u�^�i�ᖉ)� T�F|]��]9>�r|%lzS=�l��g�Dd�<�ڑ�y�NT��8hTl�F|�j�+���v�D�N��^���v;�p`%���s$��4 ���N�	��]}���V!�8�i{δH�5I۟q+��n��7���.�>��b�xy�F�gt�	��;v{�w�8$ق��|�:�R���V9z}Dԫ�.��oWNH��S���{F��K'�����_A�o_���@w%,�y'���F}Ȏ�����M X
�Sq�0�bK�U<cwN�vyѶ�����E�Q��ͻ#�T��i��~Y�[ل\i2j��:b����?>^��<u������b^�%�?*��C�(NH�RD���i3f������ۮ������M���[�����n@��\��ݎ�ѻwf��Z���7�P�!���_����o�#g��{�Qkǫ���Ҁ�1�+
鬅%b�*�\1x�q��U��u;�X�������s�6�W@�G"�YF�g����m;ޏ�i4����EM�Ę�� q
��9��qp�۱-�XpS!���=�)���ܪ�Pry�WƽO�$>=f�k��y�V��a�rlɟ��{2{�'Ȝ���{=!���u���re�PS(n��l%��g3M�p6���J�3��J�r{�tGG�XދXDC5ő�����<`~�ӿH����)[d�nP������\eg�)}��L��JM�Wh|����[5�*b��3�~C���K�w��z^�o�S�L�i2{{K�/<��C��N�}�xhuY���=��K��P2P0SN�-\xw��ħ}���7}�ەq;��5��9��!xU�gzz5�s:5��S9�����UT;�^5��0x���$P����	����w��I6!4	l1`d��W���Kl��H���y�'b�@�� �wP@��n�y��em��գ�泠�z�.:P��A~~�G�?u�O�U�y���t�<�\9%v,�#���t�ٕvtmLM�	]���[�J+;N�����`�`���n[�������ŧ���V�a�7��7��,�Ȫ�u�ʙ���|�6�e%b���Câ�����f� �d�O�[I@P��!���^̏u��W�w�/�a�8��cb�\��?���7��/V7�T�SaeC)�f���J�S��{�D�/S˽݀��Q��R2i�y~�x�L*�4��>�ϥ��r��3�q������>���^;���ԷO��O-�w�����MRy�����c���Nyiǹ��Ϳ��TXg�a�T�nɦt���{�˾w�FM߂�I�u������g=�WX��{�R<z\��G��m���/}�`�$�H,��!���{|� �zɺ�ݽ�Z��<2'��>5$8��ޑ@ȗ���!yWj�*w��ʛDi��j�V?]"ys�Xs�zjg�d���'����ل�u�O�"���ƴ=ݏ�GU_�ڟ���������,���uv'������8�4�q`���� )�$�(M8�nn�i?�g���,e�dN�Yj�P�u��=#W�?K��#`mJ�[���*��0L �m5��c��=��yZ��py=�9��9U���5:0�%z�P�/5�?r�gl�{�v�d�sp��	�B�Wf9�G~�l Mm�b�mN^.�b����^��t;v�z��v��-�GVI���{��N�Q�~�<��p�D^	�K:Tϸ�[�햶�a)@d�"�-=g6_V�S����Ct���4篺�R%�E��P��V���^�Ą�̷�3#8���jxĒ���j�Y*�3�r�W�Gs"���d���co��N��wV~��|���w�S�3��z��j��|�{��v�<��1�&����\������sy�Nnf㞣���]R
�ۮ]��I6�j��u���g���n��5q9�{8x�ib�K;$��T綆�Z��8`x1�����0Ce�=���TR��u�^�ky����u�9��7G`��/E���W�N�ҍ�O\n^k$瞼�����1 ��$��Cd�����lz��o���
1]wt�g'�1��"�^�]�w}�� .0��Y�tg����j���>����3�nG�➾�zH�swv�*�@g�9�`�䨉������U�4yǺj��Γ��B�O/�__\*���e (p���BD��Y��^�8@i&��*�������sjX���F�D&�Gq)�G/�i��v�yWn� ��8H��0���@��s�`�zT�H�'�.�z��8z�}lE�C�]����C��t��v�I_��HT6���ʎ{�'�&�i&J�
�G��՚�2Ul�����L��K������8{cް�q��:v�r�z�,o�+�ǽ�s�tc2�S�B:Lo��5.�P9�3�ȣN*[&"���s�T��x���!�_�����*t�f��}S"{�}�S�AKé�>5�!�q,;&�UOT�1]�"�x�M�ڴ+�r|}���{:Oz���9ۂf+�����ڟ{�$lt p�6��r��l�t)k6�i��l���xA�������Ϭ�ѹVr8����똓b���
����X}�z�Ϣ�0r	]��!Y� ��"a0��9��ۋ�����Ӏ�5w�'�S��z�a�3��o+�Z<�2@5�~�{8z�<�QûG�P�V�T��ϕ>�"�\�]���1-����݇�j1/,}�����5�5��/��ԝ�S�PS�(\��no;o%isХ���{ieY���t��~�5��_�����Si��<	�kH�{�s�ݣ�]�y!V��C׆�XJ?��ًd2�Mٶ���vY�f�<�8���Ѯ�s���h|��7���Ҩ��R�"r)�>r��\l�����s�'*Y��j��[&���a<0���ҵ�ѥnfU7�gs!�Â�m�ψ�&v�n��c���/2"���ӡ��N�*���X5u���#�^{�}8�7k�j�K��Z�̣��nw��{�!I��#��]���w4lsj�h���6o_��9u�#�;�=�9�61�;k4�X���4��I���Έ�ׇU<J�(Wg�]D��2���?F��Y�nM@��g�e��!o����P��d�0�^�����-���"(l#O]fK���*�����w�ϗ�������}Y����;��]<�ڨ�,���9�o)���=�#2���<Bͫ��=@B�gո6"�^�n���[�$��z�7�N?L-.�a��Js�އsIlz�`�=r�s�����y��h��9g�v�V�K�`Q��t��Ai�t�+�U�sѫ�3�9H ��y�Ռ�.d�I�=EAe2L��.j��eI�k�Z�ծ�"��l���!��Z���'}}���h���*{ޥ��?� V+�Q'ݕbs+6��t����;���Ry�"DJ,du����d:k
á$d��V����#�:��]N �Wr�X^!ck��;V��W��U�r�h�[aǑXpܼ����b�D�nF���-�0��ĝ�l_�ySJ���o:eF��
��u�SR�<Ҽ�O�gP>q*��I���X:����O��+�@X�j���g@1���2�$�������������u�㆖�d��~^���c��e�SO�[=͔j�͗r��Êz{,�C��#Ff�|��:��t+��a��+HOL��l�Bz��7�ʄ"�	�k��׾h��3+7e��Zܖ�T��ג�g2fV2�g��K,��w]�3p��3��]b���lUE�s>'f
��^���vf��2���V"QS�>�ȭ�{8ƭ��v�3��V{���2g룲�-�(��9zx�]�Ԥ��_^J����"h}Ҽ�v�y��e�T�,w�rC�Q��,���;����$����yG�������[��<�z�v#�e"cQ��B_M�>�5M��*�R�/�D�(�B�-q;E��Vk_ߴ���~�X�o����e��W7V��d����.�^�f�|�c����V�fIY9�����#���%	'��4��i)?J>u�K�*�[�*����@����o��S��m��1#�5{N��Фh�4k���.����Ԋ�J�V�*}ݾ3kѣ�� �h	�m;P�ʫ3۷'�h�I�R�����]^z�oR�ݎ�Cq���٘&ͻ7�C.Rw�wq�%�o��{װB�P���c�f�����Q�E�,��᧨��|Z�O��שZ;Ն�+�r��S�
�'�i^]�O�w�K����	NQ��9��|�yy�N+AY*�� �$rtb�c�z�Q�hÊXI�F�(�a�6\z3h<�//b�a����+��P�T qJ�;t�����s�X�`���Y\I��;��T36E�5傫iV����|���+ޛ�W~�_s.q�,d�����va�΀���V�z]�'ps����ilmLq�ޟ+���wv����K[H��_�%���rdq

�!���xhs�۷�d^���GGLf��+�D|�.[���n|�V���7����&�<r�Ȓ;�x�@|-�Q=���wh����'2��3�:�c������o�>J~������e�62J���[+ٵ{��Nw��
	 �	�{�9���;Sյ��Z�Vi�kV�����=�#�-B>9�I�j�����U��B�321�x���b�� Թ��J>���<��R���* jpGF�H>�q#��U���j��/�7� �wۤ�`K����V��iT5v�׃��^Q��Z)1� ���̸\3�u�G���F$�xj&�&�r��7�����
��0�&�ޗ���tڀLH�j�m^TJ�:ƞ����=fu�o�~>��R�.Z��S�v�hv7�
���؏�X�6i��I#��K௭+�����ff�A�]MR�KM櫖`��r��0�+����ғƱ�^J�QF��$�8.;{L�ï(�=�64���)�O	�F/�E�����ej���q��%���h��M�Iu��N��	ww��wB�]퐞wC�G4�e��七-ʏ�o^{<n���F�N��4���q�g�@�]��'8����N��O���%�M��'��.z܀m���vy���&쾏��N�S���+O�~�_��K���~�㙝~|2}_��&/�V�f�{��b����=Cp4�M^��}�6��f�����{�tb:�Dr����{1z���#	���`i��]74z8(���-g�殹��C�;�vn�=gë����\�'�S;���</����P��yͲ�]�d>���ՙ2��t
�-�"+{T����Ą���2He�by|�s�b�6.T��Q�T!mR(�`�q�O�s���r'ңAɿK����#Q��jk�G�8S�m�\��6�< �Dw��#�����1�u�Nw��;y^��ݤ���������6��7 `���l7	}��̂t�jAgz��S��/�K�_pd��c��s��9S+�`i�<�k��&=���t��%��V����ͺ�s�A��i�B<��P�`Q��B����	UjH���XR�&t|�����,w�^0�l��bH?�V�ep��/|^k�#����G������c5s�D�����^�1�=��5�niJ8��CM%����!/q؜7��1�e��0��A��ɩ�G�̭��z'���'�It�`�[~�C}�5��Ur��Dh�\����~����C�����F'��@+�2L���& ��l�`{9]S�z6&�@F�f��x��C���F#�)�bQ�s�&,� #0�'��e��W(����}�6gL��H8-,W��{���z���K���-v��.��yya�d�Z��j�g<�֥��g�_VР����#mCv�!��]r9Pb�&(�I[P�] ����z]u����7u�O*�	�*.I�T6��Y�Vڃ�[�4�q�;�����6���D�ӥ���م>�S7)e�h�V^+2��Hŕu�Y��s��r�S �sm<=	��(��7ٳTT�6�P���;�;����Ś�3�,��K\o;�%C��f��zݔ�i�s���+����XM��Պn04���6m��0�Y�b~�W�e������Q�Ҋߺ�vP:��ce�f��>��2����M,0GV��^*϶��C�?���{�K��kԬ� ��D��ϵwU������`V92|0,K�fl�Y������M�lZ�/�a*��,X̴�r�)�	�;���̮�]�vYJd��7(������̮ͪY{�������wK �om�1&2nˣ�wL��8`Ǥ�\m�,�z����gK ��ҩF$��f�VN7rې�T���N �x�R���!ׄ��5����i]NƠ�쭮����o�:��0�sp�mm�����c�O��t�g6��O�fb!����kŲ��
���N!2����;E`ei�.ve��w�1�+A7m��cО��V�̀'*\E7ݮ�uL��t�ԙ���`����F�P��^��
+��kmڽJ����N�Wd[;��	ܲ���Z)�{]쫄p	�膧t'� D�PW��X�HǛi����h���j��t��W8��eB�.����:�<0�C�v��BwiZy'uyb֮��v�^��fw^�����X������Vz�l�W'e���3��m��q�b��\�X$܆ܦ���c6'mЮv�Z���*p-Ӭ�Y����Ͳ���4Fz5l�Y:�hye�v4Ϭ9�(.���Ϟժ��{6�W'����v�i�u���x��{mH��FkCcf �{9ީ85����s:�.��^�M��!��#fm�;K���o<v���A�n��v�9��'�{c29�.-u���	n���9ǝN��&�S�
�0m���x���͘��p�B�wPj=j��4��n�,�rc��ă���x3��Z]�1ۻp3h�sYt��1̝G�����`���o���R	@<�D䍒��D-Į�N�66�� �-Sv9����6X�2Z8ny;b�b�7=u'���.|K��E���^�f����3�ڗ�Һ���/V�q���y������4��7A6���o�紉�>�)������Q��֣��yўvV��,ݷ=��{��+����jݫ�.R��{i�8Nwhq�:��I���n@N�E�OL�`����p����œ������\�����j�T��q���ch��+�vv;V�F�GZ^^;�PC4�َÞ[���`�y�������qȝ��m�9��;�8㴪�<�^&�4��n����rq���:���mց�jxx�[e������b �#z�(���v�-m����Z9�^.ۧnuۻ=��|�\�.+�]�ؚ:�Ч[�W:��*7���u�b��A�8vI[:VnӹL,��Qn݉i�8%���j�t��@.�1n�C���{�ݤ���^X���y���琉��������I<��[�ҧW	Ӳ4V:����vV	�.����m綬L/C�X4Gs��6Ft��v�����.�/u��� ��Oq��C��Z=gv6dnX���]as���Z�p�Ι����Y1|~��b4}F�Dq<L{:��D�⑄�(i�7��9�|�k�7��Tž��zഌb�q���{�>�ߩ��E�CLa��P�$� z�1"�p���6��p�q��ӴW>s������}���U{���o�5��M"T���8-|�%_]�B�Q�~a��>���$DX����w�-/|�]��~�bv�	"&P���s�u��'{�B�D�	@�T��G��U|/�b]L�[�f��kb�ͬ�(X��#�#�UQ�J__TA��Vb�Ĉ��HC��D!Hǖ�E\u�U3��3�5N��C��K�g�����(B�%L��w]�5��x��߹߶�h�}s�ƛDrхrr	=s(�f>5��u��J����w�F.�L��">�/يB�ܘ�(�"�v���A*/Ѡמ�w��w��EE���B���V<P�c1wm)�����f��ǫ����u��@�E��}�t0�W��~�
�rs�r*
d��$r='�bޞpT��2�����'��Fbq�)癯��b����!e�~z�ِY��&�ށGd�D4}=t�����^��z�_��$��K��Ę����Eo9�Gｖ�+�A"h���c�!	a�׋߹�����/y3�,�����I��Ju{jw�eQ�h�g���I_~���4�N���	l�tք���p��]xQ
I�4�1�?~�L}��L�d�1O����m`+��b�P�9��ڠRsq�0G�G#����Lǂ\��B��}/�#�j8@�& ��3ޘ�D}���]�i��,�\ɈC���i��J��3����]���]�KE2��͙�"�������mXޙ6QM�K��A�rN�4�r�g�9nm�ֺݼ:`p�r:Y���4S�}�Z�Z��$���-44P��`��	(!�D߻g�$|��~�>`����딹��#�ۻJu�%�~!��Ι<�&{k�u�}�Ww�����NZ�Y�[��Q�y���hj���0��%�2q�������X�XzkkgsJ�:�1e��?��kc�_P���z�\�
?��\4�B:ŭ�ftP��ޫ4%��1.���k&��=��(��תG���zp]5���S:���iJ`A)�rw�7�~�w��?~3BLٟ��I)Ӫ��$���������E�o��y
bь��]�11�!���0��Og5�l(+l�\ ������|du��u����{������}��������n%�?Bd�����G�c��(��dG�o�H�B�lJ˯sY�q��C02	z<L�#�8��치�Q�1����m��ϴ1�2��MQxK�|_ߦ~����'�όRw�/Ȓ��!lh��~O=��Q%�y�c������<�gD��S;]���TE?���6>�~i�����Ι
`fC%g�e���k.�gJ��������"��vv��?=�#F��>�!`�,}���Fu�ٯ�DW{A�!H�ڇp�E��C<%��rywZ�9���{kC6A/��w���O���[K�y�Ę�m�w4,f>5�N��q�ǀ���]:bb�����pb�Oغ���>�"�1�7>'/���H�/!�%y���5�S��5�3�0�1pL�%��
�ew�y�o���Y���,B�q+ư��t�D�#SS��~�{���1k��b��t�i|QA/�������l�k�����YU�����`���-��睁�A�I	���)���en�C�{�~_�-ǉ���:gIEǞ�-���g�����!�1߮h^$�>�Ž���_k�����5���5��J�q��bg�����lg�"4.���Vb
���T**�8��L�C�6�b��K���u�;�_�<�At�3����(%����}�ߞ^�KB��%�~�(8��!����%�DĽػ���WO6$���֔F%�Z�)��ܟT����r������,!�ph���f!MW�*�ә a��2�m"���H�����G����GǦ��"s�(m�M�)l�p_�b���,R��QY��^	���>gs�R�Ԫro���v�:�dj`���a�.�����5�"�����g�b�y��3�iQ.�k����͉i?t�)����b����V�w=0x�<�C�L��139����ԭ�l}B������<>��O�����c23AAsD�(��e͈�>'��f`l�x���uߵ�N��3��t�ס.;3�PŮ�e���{z��Y�?V/�U�}Oy��-	7��U�c8/ڝ���Qd>��D�1:��^a�ӟt����S�	������c�>"4���"����� �߿%	�	�?�_���ߨ�s��p����>����i������K�38M�4fu�W~�祲~|�^���|Z�\X�$�׷]�_BD�4Y���c�\>Q������������l�߽��׵«Dv���,1�͗Fz4g"��A0��8�!��O8%g�鯾�oJEF<~�ɤK��F��8�c�$��.�j���fլ=x�y2w[��W&�uUq��n;[�l#�a׳=�����e�x_�b�g�>�2ѓ�~�ėϑc����h�j3���ُ�"�(�H""=u�{��=�^�Ψ�B�3�i�pBp���:g�N���\1񂷿t�󆍔��b�ip���>�*-�����16~���A"�d�a157�q{O�>Z~�*�vO�#��$}B�v��:�S�������U�t�fkrbW��u/��}��Ώ���'2QVPp�pZ1B"&9(����!g�ꇳU�=_ cjk�^ӿp��>Qb�����K�8UWwv�����r�!�_�"#
_Gݘ�~>���`�������!W��l?�aT�h�a�f*�HAQ�&/����&�߽��qѕUq�W�x��e�V����7ֺ(g��m1-&��i~�}����g����N0��B��L�w���F8˸Q��c�sA�y[Y�wI��hP�J(�Zg����c����R͹��Fv6�,Y���]��w�w��g"���m��%DR`=�Mv1�x�`�q��t�w'��ݛ��d�Pe�)�Îu�$����Zσo��|:�y����ۘ�[���냭�k<L�#������s���{�}p&�EҜش�=L��0Pr�{9-c�.:�ӌ7]���d�<u���l���8�0X8ؕ:7[;�4k<Un��ԁ�iey�=�c���=�Ƭu�-��m���y�
��w~��~�k���'��~���L!TE�`�F��za
O�&T���>]��F���y0�7	�-�q}B��'F�h��r���
�����B�Dh�	"DG>b��z�Dxr�r%����-�^t_~��iSu��]��jHz�u����+�d"*Js��ݏ��4p��_����?|�����s|'����XZYa~�����rE���B2��>S�1B40��L��6&=��?>��Fꮹ�a��]OIB�\���c�S���d�ث��u�JV�|_	tГ��;@E��(�b��^�a��8X���;{rE�"v���X�F"ʦ{�M$!��B(F#�p#��=v��,��+s~]^뫣�=�Zx���M�z!#�~Ȫ�xக�"�w����OѮӽQ���)��7꼟�yBe��P�1�5[��O�o�$P�Cб<?xBh��c��s��bb��]��t���_�+�=3��(���A�ȅ���O��ǞnM�n�7�]����]��7t5�ZJ';��U��F#�SU\%���b��=[&h�c�'轃��MC���5C�WX��0dP�L��>����vs0ހ�p͏���D��<���[&6r�4�/�!�q����x1"��yиB8@9Jlwb����\C5�����q^1=�g�P�Y�~�:����?�����'��Ţԩ�2HA���τ)j6��5�FD��\Je��I$�b� ������E�3��Q����˄�2O�:?}����@�?h"x��V&*sz�<$�~�~���5��/	��@	�(E)�f� پz(5�r-9[W��MS���][M��u^��^]��/��`��C�]v󢒡�8T�6�Ys7���+9���D���=Wy��?�5����kݕ�����RT��G�LH�����Bv;4��4HO�Z$z؂+��56�ۢeҎ&0P��C�'k]����&m�Q�E7�^����9k��Ѐ������g�Y�C�]�֔�G��A��ޞ���V�
�3��|L��=cJ���wk��y��Q^�eo;r;���D�b8��& ���{��Ӛݳ^��{�4�B��H�LQb��� ��
<�G��N׾��6�����XϽ��ď����q(�<��~1��d!s!Ht�B!���c����u�w������_�J���h���A����~�[j�U�\"6]���P��U!b��6�����������DQ�b��߰T~k�e����qJ�3�G�[:�EO�o/�(EbQ9��f���[��UXc�S�g���j�gH�(�rɃ�ЇOl�Q�n�?A���:�sihbu��f���.��3,��a"�%��=��>=]V��+���^��&�M{�����BͿL�����A��;�����#�(�B�Q��R�w�Ū���#�<a�Nf=h���\ϳ���@'����6_yxF�9��,��	��O�U��jkøx��x|[w<(H�[P㢫*�:��;�~�(��؉��+����H���DUa��A�U+��KDHn��ɣ9��͢XPaC�#�B�/�'O�jU�!5��~9Ȧ>��v[G=;����7]�}�>N}�#k�44��]�&{G��J�q�x~M��	E���������ݞ�)���yt�GG�@������Ј�==Z����P�c럡�r6��yk����&����&�����d�3��["���_�+tC��`�;8^؃I���<�v��0r�bb*�.� �+P�j>/��Y��S���1�/��+"v�Ku�w>1��ey�/g}1U%�����$D��#{��:�&K8􆙁��1�2�V8��L޷;�I�6~�-��>��T���Dx��J��wuR"c<;��%��.=1;ɿ���&��<R�E�I�M���ϣZ��n��(*&n��t����L#D���wO��������\�F�ǩ;��]�;�b���?p�j8�as��R̺���j�d�ih�97�A?�>U�G������}l˴l��&0.��H�K�.h�%�aK<�X��@��it�"�:��AL��m���w�zT�#��U��N���;A�Z�� ���߁~��1�X������ˏ{e�""�(��9̟�E��~��Dt��m�4�=o�(>�Y1�k���1��q��q:�E˾�f�oMeX�@����ózP|���_f�i�(Ye8j⤞�4��I��̩z�:�.��g%(�V8ߙ�Og&��pʇWb��ԧ���OZ+��ߏ�q��yy�nc��9�4l�y����/�0���μ�]�S�ۈ�!� �+���:]�։�� �"�Q������F$Cmv��+�����n{{9�ט��Fo#	2ʀ[E���ip�C	�~˜ٱ>"#��c���K���us1B,D\���Pg����n�}9��6�r6/�!OC1�D^���L��`���e#�g=~A����;���I \W�6�q1���4>A?fz��ۢ�3�����nC9fE!R��|_}��N�TX�a����n��j�x@V��3x������u�\�#�I�F˜0
Ϋ\�����8%v�m�j����?p��	uM���7�P���v�� �B&�zj�o[�&��#�f/�޸xa����Bբ4�Tr�ǉ�[O������wTK�:s��.p�}6`�`��w�{�o�� p8�E2 ��,��~�^l�����:��.Ȝ܃�5<i����O��?"t�\a�)>o<����G�M{�����r.�3k��{�x�ц�I���G��ɯqM�I�P�ϔNM>��ET<����
q�\��s컪k�!����<$X��K�/�$M'�y�W�{c��3�Gw��F:bdͽȯw7�	�}B�<r��������Јd�` ��"�#e^��6.��K
�c��B �G^.�����'��#�R�"��؛��s,�:�w/U��in�,Z�N���B5�������)��{("b��.`�]뛸��u�~�W1��S��pl{�g'�!(��(��=�#���u��r4�h|!�]�&0���d�6�z���h�]��?���H�M#>����NL�E�9�/O�����VO%�"C��w��\� R��A����ӽ��a��Ԅ#� B8M��\}Ԟ�;26��{��{qo��w���S}>	EbR=���f�p`�"4����}��b7�=�E����'5����U��J���n�I��J�:`U.�ࣾa���ł��u6~�fɂ��VPᛒ ���En��Ɋ�_M�h�aw����]�趾��,o�I�s��k�&@N��W`)[�][�&�z:gϮ������~��3	3r.f*�H���I�I�`I|�u�L���5�çm�]���Z�ѣ�^Q�h�N:C��-Gnp9�V��zv��t�k^'u���<���u͟Yu�$[���[��KD)c��8�y����k����=q=�R/e��oj������gRs�0reMlG5x�p�=���ZRr���\�)�=�ڎ
���f�j:�&�9m��q�����)B\��l������q���g��6PXhA���3M�7}^�E�_H�p�����/�wS��as�� Cp��т(!u���3QZ��R��D��,G%���P�;��Hh���7�4c��T��(a����>03���ί�h����g[��{�͌h��X#�j1m$>}7��$oFj$sd���.���!( ��2�<�D�dŸ7Z��^�F�11h1i�R��b�n-��E�1��K�i�;)��(mxF��v�����tb<{�䶵���p��Z?d$#�W،}=���=�����$d!}Yպ];�O����y���U�9w��s!.+= �����!��Nr�¤�b�{!MJ_�&����D�C�B�Y7{v�r�kB<�׻���͏��Ҡm�r�Y\;ޯ+��#@��<��םn�]Љ�фX�ߢ�(4 b�%:���UV ��N�k��A'��3�j�ЕA���Ha��Kk�}4c9y�H��;�{j�E�zʽ+s{�	^OL�ש��wK��/�A�m����+�F+ք���lؒxϔ�@W�D�_�}~˵O�R�%��Y����%��{�ׄ~�>�O_:�Js�fmb0j_�JQ"���:�at��щ7�;�fB��#��J_ZǺJw�x`B�Z���}Z|A���t$�����UkjR��(>�OpJ����r���+ٹ�4.���m 2�P}�)`��v�q��L���:���G���dY�J���U1�`�w8��79�z]f���� (�ۺf�8�Q��$:+R-�$P�#pqG����,�}�E>��<�����GZ�w�i��;׵w\N�u�|������Ej���"�"7R��:��%�{W<d�e�$4!�%���G���8w#D!�EFu	�UNv���(���iwueJ�x�q�Ƀ<V���������b��f���3
����3�eky���``���z�2�|xu��j4H�E��4��/;���T�?Ӕ�����R�|�����N�ˣD�"+���=����t>w�#y�X���
��q�]�	����끎������L�����{�9��o	��>Q�Li�9�+��џA)v���f�:�$��^<3A���v/Z���j��z{pw�mBI�K5`�#;C`z�g���{eUz8�A�:�S�W��齍�=��A�����ƒ�v��H�~�<j��&z��B�㊗��5�F��t�e���C��6G������]uPu�`�o/�d��}q�R�`���!������2�S����$9h0��)��%���}�ݹ��^E_��.���R��� �n�y���@a��-0]J>���;��[^5tg�VF�c�u0��L\�5ʜB,��C)��-:����L$X�ύS�64V����ըN�J�2u���{��~/�נ��J��:`CX�Tt�Q���O����a?&�GPq�zr*�7�o�.+��n�6uDT�5Hr�r�V�V��n��[�j���0,��<�ԅl�n����������$��}Y��/]^M~��ؑ���4��B��N��A�)䱣=�ɺ�liJTc�cǺj�:�8/	�CA�����>bg<�.�2fѕ�=%�Q��~��; ҩ��RO���G}�Q�y(I6�Du�	cI�����eϪr����k|����
����sO`�68P����9���}9&|����j7$�h`�����m*���j�zq���	-�Af�;�w��+/1N��exwJXK�W���G�fO�{YB��x�݉�Yk�G�V��,�O��y�����T��5�L/a���w���`@`��b����Q�>n�<l���h:�o'%���r�X�G���v�6oU�sƹ�Vk�/kg၌�o��ͫA+��i��ֽ"���9Vl�l�?b�����I�ׁ���c&�ݪnߕ�i�+�n�:��m���G���x[=���b�HjW\RY"�h�=�^4�j� ��2��ݯ9�L6��.�/^+�X|3�����p=vg���<���$�BhAl"�]לv�:�X�h��2�-���u�=������">�47��v|�XM̂��Z��f��8L�{�Yэ��tEA|d����33�ř�󙘖f,��|��K3f���K3f	%�3ft�ř�3?�fbY��3�Kf,���%�3f�31,�Y��i%�3f�fbY��3�ff%��3<�X�1fcI,Y��3y���f,�����fb���f,�����fb��환�f,�����fb���I,Y��3�%�3f��d�Mf��� �5~@Ad����v@������|�  >��   1��SM(���xwԩ��  	��� u@>�x;���BZ�Vآ �Ca��%vԨ�i@�D������r���A��UD�Q��9WA����P   ��IE���2��4h0�E?L!*�4 2  �  ���U
�觪      S̪*24�@    ��$�� 20M  R�1	��CI���z���dމ����z���In�j���@���*��EIj�i�����k}1�C0�Y�*l$�i����li�%-�������Ѧ;��,�4�K��i�����ӟ��ӗ��iԜd�����п���sB|�����Ȧ�pj,���h�%e�!��P�1�wH�5iX�9�Ә���`�-&�p��e:9�kR��t\�U�_Y4�1�7jl��͉�`�t6�n�f�f�B0d	]�v�^Ә5��x���Pa�f<���.ᖡ���I���ݓ�"�߄��mI����W�(�9�����+��1���&���Lw>k{kt��>�Pj�m$)��o�ݫii��T�L�2�3/�ͅ搥�-���ܔ���Su;����-�M�K�;YFK���Kp[�f
��p�����ff �,�Zh����V�@�NYD��h@&��˼`jÚi��F�^��i�ײ�jy���3@?��QȱQȜ�T��X��\<o&�,��+o��[4k)��7)�з[��՝L���K�y04�%vԍ��lV�V7'ת������X�� 3E-y�5�՗�a�d�nI�)���%�*���{6S3+"��m��ʎ�ͫʽR�Ry6��i�X��e5X2���,�˥�2�T5
�e�6�h���ϝ7�������U��R��<�Xr^�ؒ�T�2������I��m㭂�7)b�Qaϰ̼�c����\��䦷�i��I$����T��4�-Z�&6�aq�e����ϯ�~�o
�"1��'Qw3�   �R�cH����]s��2��c)5"��m7���-Fi���M
�0�K.qnb�st�,,�ct�n�ZF�v��n�k�jKVѮ�l�P�2�e�1մ�������m�SE��XK�i�\�6�.fB�٦�k���i��MYL5�%�a��h�l�M6��M�����WsX��m�DH\5�X�$��hg/3�*ְ��ج�B�m0J� �"������L�Y�s��6ke.��M)�-�%.�Ǖ$ҤM.LLB�%�q�5���L^`�&���4�#J�M���[��.���Y�Yu�S9r;��*l�ih��۰�8�m,�i ���VP��.����J��e��#�f���5ͬn�k���n&�T��%�5���7��
�Z�,�cF*mYyk1\\�N�sIEKt�jJp���۔]�i�2�%��b��Z�K�0�U�q����37t���EU�̀                              ����9�	δΜ}�U%֝]z�"�C��-�iٷ]�W�:��
`�$�eX��V���L�T��Ҋ'�J̅��>/�3��T��}~�b��8yr���0�C,�5��T��x����Mn�v��Q�n�_j�������m�Cf��䍘�w6��*���~�CoW��Hu��qv�N{n	��:���A�8Q��s���o���%�����SH����J�v i�+6��zI*H�,ae�}g�d+�	R���t�ҏ��[,���P��7%�(#D��N������39�Q�  E�xJ{�EZ����� �(��w6"ME�a]��6���j+���=/�E���z9l�赊�΅�O��Nٛ�˃w�P�x����D��8�"��G*�%g5��f��vg��}�ܶ1���c�)4�D��o[�.�=1�ƑIX�2B�I�iY[ �@C(Ye^�wyw��N����z<�9Eo��靪�>Q�R8�L=�"��1gy\�@�
>hi]��&aMP��Z؀(���P^�^���O��'J{�V���]��u��.M[j��
/&w׮�̱�o�Y����խ�i��x`�#�1�Ff�OEUd���X�	/K�%�;�/Ž��e��V]�&���t@��I �P!�1�Tke0U}_kׯ7�i`;�4̾��ǲ�4�3!��ԵuC���=�x<�:ko�+'��a~w�}��c�L��}u�m]�s��C!�e�k�'�pѝJg\�	����x-�SL����Ct^^��o���Y��i���I?m���w�c�6�u�J�-C�Zc!ǚm����%)��DѦf��W	��юbF6���Z�;I��%Ͷ&�孔�Y�`��m�i�
Kh@�Y��nb�KP     6����Ϟ�k�m8s|�P�w��)��-3���94��:���vlz/����*�)#�,�N�1�����UE$�Ar�C�[TG,\.�3}�s����5&�O�iK���z�H!Ė��	wYā���*�y&�CL�
p��5F�\r�`|H^��Hd��p�e�+z�0�2�X���&��r��
fU3#0���"�+\5ě`E�es�N��1�_����{�#�̝1\3\R���P�S&R���q��|�'3@X
L�$:��@��������W+�<-�I5z�AT�XY��[m����fl���<m�R}鸹n67�'[1p��[v�B���P��M��Q)��{��|�O�Hk�����L���a��xUhdR��t���&GO1��{co�� �Dulz�痱{y���9	|��ߓ7�F����`Q�؉�/h�1����^� ���y4�`S-;��:��kɄ�W�H.���cݸ��a��ZJv˺8��M�p�f�X��)�b�W�X�I�)>�������{]���_^������2����Xa��0�:���2߭Q0�(�3��Zy�Sv�i�}핊��N��P���S���n�Pi�s�n��*����Re>`R=�%��'Rs~�.���"��k �ӛ5z����ֳ�u�꾜3��r��q;��f_�q��MU]E�-�l�2���C*��@��icw>��!��q�C�ӼU�05�U�p�V���ۆa�a��>q�4�!B��N��9�L�^��e)�e&\�Ә�[��gU�[������m�RZȈ�ĸUVKe�ׅ������u��B�@]��_P�u2��Gn��Y�o��2�>�{Tm#�0ۄ˷��n�L6�-�7뾳H桇�a7u0�)�M��ǰp�=�0��)�1�x�N��r�f�I�	�T�<�_ًl��ǌ��I��6�x��i�nٖJ��m
�&R��Q\��D��ٔ�z�1�i��f���L����g��a���&k9y��fl��Ln���CtX�n�/b�,��1N��&���<�O���q���K��Q�5�{Sy%=��e���u�ޞ�i�H/��i�Z{ڐ�U�Ț�(�a��d�V�T�{gY�m������xG݊���� G��QU��ѻ�8�b�*b�w����M�nlm+��흅�E8͗]Z�;2�8�i�âp݉ۓY6���VN�D}<��DͶ���5�X||偃�X���e�7��sXI��2�<�é���I�l��ۺ�.�kT^�)�=�_����m'�Q�0�H�wXM&R[Ĵ4�$���)��)����W���~�0=��s��F]e95�-j�����c���Z
a<�M�{cD�;�&�|�0�e�n��׫Պ*�ۄ�e�.��}sL�)���j����-�y3���p
i�W��E8�Lr��Pϱqd�+4�[o(u�ڳI6�.�$�f��U��K�����b�q���5Yd�8�Vg��VO��m���V�>XU`)�)]'��n�0�U>K�RLb�8v��7��O&�3ʖ�\���}g�iY�$0�)��.�����x�k�\�4�x���I�C���{�3���0�������B����ղ@U��������&L2%.��9�^��FS��X�@e�`���kގ�Qc"��֒��Ofb�lg�SR7`��*c���l���vDY�"D_*ii^��.��f(.{]=M	�sK��ꊂ!B%�J��-�!�� �A��%��m�fmj���0o�f�߄�!j��E�����A�2���d�ޖ�.��=��Jr�y��a�9�p�خȻZ�#������]V~d��!�=vI�[��'\A{�F'�eLU�j��X�R�:�H���"&��F_<��1�������g�Va�`VOe�u�I����	Di4����2y�64���Fe��/q\a2��i�rӒQ9>����>�VI�K�%�}SP����bA樖���Bv��1f�gThCG$�E�LU��Xu19��0�O��@#`��0 ����	�BU5i����)5`m{*g�Yu1��	��T�h��!̱�1��y0�t�훳)E>7���4��P}��5�^�8�E���/}�9KɁ�=�Mȴ��j�)	��ogw5(Tu����$�݀ҵ�&�1N	)�b���=c`�sW}�%��I+T��+Í9n.���&R� ),�.f�B�e���[bؗ\�\���Bǌu@Uf��B���.!��]��S���	HRh2�3iQ�D���j,�TTؚX    m��m��¡|������=WV�6���4��ٛ�AK��i���kcl�Ⱥ��4=�3���E@�ɧ�{�n�c�9����v�&�(�cs:�mS^I��8!;Ԩ6��md7���E���z��vMr�i�qx��1(�t^>U�Y��-��[[Q��z�DJ�$���pB鷵����e�P.B�G��v�x=2ʑ9y(�W;ow�֞���к�3LV`f�j���a$�m����9���&�W�S~ w�:�蔨>�3ޛ������/+F;�23M�5XË����,9F���gD���VL�ift��/��S��{Ɣ��H>j�L���;F��`^�WI6���)���u��+Hy���; ��Fg�T3	���Vr�6�)g^�Ƚ���^���(��}�������V����+Y/���%��Ҷ=���i�C��eU���x"IC�Ge~k]�X�m�N*\���/^��.����"�6�BgA��0[��kj�ٍJ���(���q��L$F�R�L�.��9���+ڹ���x T��W˲�m�u�t�	b��Tم&�q�L�3ϋ�c.��r�[9�7��Y�����#���<�v�݃i�M��|��g�]we
��4�5��;�}��ӥ��G�}>��n9g9t�\���,�e���v�[P�[���*��}+��J�a�ڶS�ֻOX�ίU�
�TŻ��������'Z��U$����opubU]��F��{��?<~\|��Ƿ9�3_�w�"�x��f�-i�$��g7��;uq*ƹ���@�DY�Y���l_T
 u���S* )@I��2�G; l*��������מ��w����4ҫ��H0�z�ԓ��=3�3�	��:oe��i�}�Gr�K	��]���3yeGT�3���� ���ܓ/V�n�7Z�0�l�u3�mG��܍x4IT7n����x?�Cs�"��΀^'��E�m���A��Es�9Y���uF+N7a��Nf�nk�ȶA;��D�nMq��M-'~��y�g$`���Й3�+���+@�e<�<��󏽗ueU��0�\���<�vW�7���|����^�:�ܘ�\x��P�@��\"&��BD�m��M��`�+u<��,��4l_�fo�%�������+n9L��*���N<GB����3��`  Lt��]�`��jp�w!���BrUx�����g��Urj�9e����"5�!���֩�r��*ϖ$���m��6��"��
�
�zY4"�u�f����z��8�e�s\��H0��;tNl�"�S�\|Ep�|���*|}��5|L�
�Rf�z���O=�Fm�ջ|�O�?�����8vl���Ur�:w�uw?f�|.�-"m4��V��t�M�k0Λ��3νo]��Sb:�к��[,�0 "�h4�m���2c�M����=X�fʍ�	���c���O�v�L�mk�).p9qwƪ�?�Q�H1�JC��~Ŋبw����W�����!w��^�K7np-�[F��ֈ�"U�.��r;�Ɗ�{��yr������Ο]�a�k�����u���Z��.#���5�xJ�LD���eu#k�2[(Mu�M��JeRJ�ή�j���"���]��g���0�5%�f���!�K�6�J�UUUP   ��W�7�*�2ۉ���&D������ψ�ڧ#~��3��Z	N���� [�IT���]>r�
f��Aa�&)�d�[%V;O���j�7<�S�uL�/���B1�>˭Gl��z�Х��!}�!t�_t�[��,p��ٝ``g`��-+�]P����������Yق/�c��z�(���|h���CƏ#���2�iöR���wǘ���TPJ5�[E���W��%����T��3)y��D,�[�N��:�#���Lq|��ԑ�Nu��ɣ�-�)=��҇W�&��iG<Hq���� vTtx3�Q��u���{�d����EVr�{R{!@�B�X����S%�� R�2p0*����rЦ�D�Vq�p�Y����]������to�{c�a��m��?B���7��|��a�{�(�K�Z�޵�~�W����\+O��מ.ALK����,����<b��O�$w�R�rؙG��J/)hw�߷�.�]:���z�[�u��\E��ucq
e$�M �M���N�>��aW�Lk��'�a�k ��������V��ٖ��s�G�,vmq�}�.I�w��=3"\v��p-�j�z%���a'�|��ִ1���L	���)"���{5���b����3ۼ�%���oسN_�"gg��=	,7��:5�B˰y���Q'^I��N���Q*�f%o&���	ܟ^���6p�Qҡu]�&��wm����'blP�m���"l:ͥ�9D�a��d^�99{w�f�E�\�0ꛓJ�f������X>��k�[b$�|�����߲%6�%�^�8y��O=Eq�p,e�{mt¹(@�S�IXw���>��9��-�f˛.��Ynn�¡�)���# ���ˀ �F��d֝]2��ss\���{�9��ø� Ɖ�e�h�(G��E3|�V˗&�M�h��/���Ƶ��5���$�te&�Yٹ�"Db(=�B%��1�`��b�"�4��gj��i�����a7�i\�E�c���%��kk��V�J �	#e�6ϟ&#8�M\�Ǉc�$^�9y���%��m��ϝ���S�f��*��D��$UB��`�k�]�n�.z�桝��Q5C��1C(��,$>6
�����%$�^�#��vS�s6:��I�fT�]�:�fU[����I_]l�#��
Z��|�8b�4 F�#���O$Xs:l�l�K��<.6�ǭ�w/�W�y�c���X�YiV)燄��S�Qpr�H��_w�{
��J)`��kMaY��ú�2U��H�qqm��*G}w�1�����8�#CK��:SGl�Ǥ��J��}s��b˩�����|�o��(�\9�\o�תVֺ �!inu��'��O;��m�c�J�9������u�������m����+)6�I( Z)�m�BriÇ��^��('�z��Q4vk�s�D��޵�K	��1��k�p�o!����/+#����ك�r��X����ɩ��*�,�#9�5��R�[ U�Wm^Bހ�z��-�ޔ�2q��U��]��(��,��cI+���%�Z�Gdu[osn���.���6��΍(��u�5�+JA��,ܹ�΋r�5Y.�	o+� �k4f�L-�..�L8�B⹀����   ��}n�ʽ�(�G�V��~Q�w����k��U�$��YQ�`�ޮ�~�Gz��,�L�*5F��3U#��cת���l���z�=^km�u��^�5ڻ*y2[%.�ŭ"1�⪘��6汻SfclEj�{��X������V�>�]�!��,Vi�j�U�rc��
+I3��氷\��qŤ�&9ve�'&^��fNH��$v@!� 0Am&M
�H�t��i)$�qF�9# kb�'�ӲJ[��j�+`���bFm#8^�/����W���rK�We�/s��r)G �M�r:]�:ce�ں1=wl��h�WFzT��K���m7V��Ү*�B�ś��$�gk�XO��A��۽���@A=��o$�3�1}w5tKE��l�v*�D��R��!��.�V&I&�7�R��fʲz�3u������l8p�-��ox*�i��|��&�m����q��=x���vU6�f�,Nle�A-
D6�m�۸�[�1u:֋��;��L��WO��*!����l}w�^��w�!#n���!�˒�E^�t�։��q�l���8�3�d���sZ�ȢR�9��]	F���ċi��!.}Pu���fM�Ϝ�/y�Troʒl�n��г�%�騴�&������:�Qp���Pn۰�^O�#޳�J�����\�,�^b:N���̓J���f̠�E�K�u����6�8�
c���xm,g���էh��"�J�5��cGÃh����h_�m�z;��ڷ-C)�K/���D��m���(�c��>|mv(��{�}����Nb�M06�+`2�M������y�#]�]�]>�´3r �G���Q�w�@6���	�i�.�Ns���5B�Pvkn��&�Q�-d��K�,�g[����UA6V�ڙG����C�nv&Rh��08�-I��O���&;���).H���f;�۽��y8p�g6�ů;T@PR�{�ʒ��̮�Ύ��4����8��])��D�g��\"��P�i����!�ywL�j9X����>��ce-~��Gr�>�J$��yۍi���[`Z�Ȕ�Q$���D	�B����.9�e��s�U�Պj��(�3�0թ���GFWq��CH�Z���ntZ��7j��gڜ�(F7~�xN�N�����t�w�"v�c�Y���Q��V_���7�A�f!W٫�z�����dYs�ess�6�|l�걼��z��{Ik����6	|z��c��-!�i��|�p�k���������6�Ds=~�B�?_#����5����m����Ca9"������CF��s���l�D�5�.����J`��7��R�B�����*��WMYs�����Z�t�jN�Is9erb�i���>���LGǶ���w'|�w�{X���S4��w�-ig���tV���ʱ9�95���2���9��ۀ;C�*���a�x������`�Zw��V_4).&+EVm�2<L���#�kj7:hcj��]���n�ikmblpLһmyfm`W���4fl�ܫ�e+.�h#��X�ј�ڡ��a����b�D\X���      �=u��c+��u�����f�>�$umZ�:�m�����Y(���{��E@�*9Jp�c�I��{��ںn-R@=3�⛦�4M��i�Ռ$�Z�SA�2�@<��cZLt�đ����=-ݬ��ɼ�fr�^)���Z%{WMɚ�Z�����kӇbŢI������닓Ȯ�b5�uTdK$�*a1i��X	��p�
�7�C[B,%�A&-wx�L�1�Ψ޵�9�����c&_S�.h�HD����˷��7kp�m<�5��6�}us�ۇ����¨h�����{*O�u�.����*
��<�(2�y�� i��ĝ�~��L�k%�9^]K�}7���O ��8h�r/�!H2_Z��b��B����x=���Y�me(���\�v]����v����ls��:�a��G3�a�O[��
=�Y�ߙ՛� �V��6�(�PT$�� �D�i6�~R��f�`3��V�N���j�\͕zx�lpcd�l:3��#Z�T�j��0�*���R'��z��\!	h�|� �>�rr ���UԳP�7v.�I�_�4;r�����6	6�Ρ��Ft�g6Nh����ƃ��"g��bՐ�Q@u]*3
��`h榑�&D:���1_�,U"���ia$����#�_��bܶ-�N=j�Ѿֽ|5j$�>x�%`(:�]�T�f��J$&P��H�Vť~+�
Iu`i��}?��~��<ܘ��r/��뗧Qam�ߨ}87ɯ'N�}���p�SE��pI%���������_�=�I|��RK��Ԗצ�+��B��g2��^�"��/\����]_J}_�2X-��ѥS��v9qk���>O�-��kRߴ���-�ힳR�331��/����{s�c��i,L�Uk��Z���8��Y1�5�۵��m��9^�$��Ѿ=����}�zeлHpt��ŷ�_y1}����60�zL�%�3�y�f��@���3�<q-)�n����OC�'?Ի˽��s�ޟ��^It��?.��/������ķ/��s�d:�)z��I/��ߒ]�[�{=�i��h.��4�8+*�mI��$R�;c��iu��ς%-׆%��o��l��᭶|,х��|4��ޒK�����K��K���uOױ�_������x���*�n�4�Qv~o�/��9^�y�%��T��OP�_Wql�}~�O���<+��v[n[Ub̧��d4����'������T�{Z[s[��MD���㳏r���4�{:���O>8�����ޫE�VԸ����$�ňy5k�U����I.�wű�������Y������ew����N=F��]��BC��-h