BZh91AY&SY�w���_�`p��"� ����b6�}�$��U�(��*�+l�,�Q
�J�25EJ$��R�iD�P�$QR�h�J(��UHUR�QUR�Ho� =H$���H$P��*�BA)TJDH��(URUEU��))(��JH
�!{�e������h��Q<��-}�v������׾�G�nu���d���l��nJ�ϯ��V����(�u�y�=��f���|����y�pi���0u�돾B��޾���_%�ػYT�-���� ��	I-���}���}�{���U^���4���q��>ۏ��B�<��K�c����*�o7��q�h�o;���77y��y�}��r���t���;��}��e}���s���%P�Cd5����@}{ꔯ}����h�X����@h�ް������Wc�u�4���@����oCﶷn�5g�{�@����ց�k�뀹�ӭ��}�)�x<��Vs���(��*�UT�%�� � �)T
���r4>��n���M(�f{�݋�G��ԕ/�����C_e���`z�v4�7{�Q�}�_|�����t�ڜ�%K���r����l�}���٥�����A��d{P��T��d<��oER���>��I��Ǘ�CI�W=��}��m���;�o@��X��7�P�Οkϼ��U3��5�Ľ�m�*�é�}���z�.>�}� pP�dT<ШR(��*"JQW�Y7�}+���Cy��y�:-��w�mW���@������@<پm��lho�Ͼ}��K����>�폾à#��*x���a��ԟ����u�A��{� y�\׸E �@���֟ �8����GO���tPzDw����)��Ǿξ���}��P=�|UI�޲��+T�]{�}�/}�ǰj����Wn�^�:�=��*x�o�]ڐ�ޢT���T��>��"Q@�I<�=�S�_/z`�}t�g�;:^`K����mꇠ��}�������{�׭SD��4�7��t���A|�z�}�{��r���������G˶4y�xRJ�����ݽ���}�ܽ�/}�7��|m������a�T|��s��y��y���R^t}�����n�����������:W]��ry�4������>�@_}�f��ҒW��+XB
�A�𤄈 U���G��� � ݏ�g�(�t>�!<l /��GJQ��|�_�f5Q {����J�֪�۾1�ID��r��l�k��1U�ϪQ}�/�9�5"��;�wUS��;ͻ��WgL��| B)�D¥T� �h�# a EO���%R����   ��&B��TP    ت��*��0   �~ɒ�j�4   � 4�ҩ ��M	=SO(Ѡ�A�i���O��?������,���r���W�y�=�ʠ�&����4��)�I�ww>^�n���;���wN��>s�I�ww}󤓤����t�t�����N���?�$��wI:N�����$�����R�~�>O����w���k����_Y���u%�?&��ο`�L����C� �^�D}��G�@�˂�e��-������R��bowm_)�?F��k��G���l(:�c.���w��������Q�7_s��<����(��S]m�4�4����ʠ�[`Y��i������g�c'�t��td�d�w���:�t��fo=\�q�[���lüc.�h4�ehX
��Y�\�`"qƬ_ʖNC��zo���͎ǥ�AI��+\�e�t�7���2��YFT�4�#/�(6NUԺ������Nǧ��yOhPZ��D��4��{�ZU*Av�.�	�.oo2�y�IL����`��\e�!� R��Jwsea�u��|'p�*nš�=	�sIK��0k�K�2O�o,'b��xNV��x�U��yIe�2F��K�ȁůp�!��:t'i�P���T�T��V�)^�lm;��M��z�EQ�m����wNG�Q�K�嘔�l����U;ͥ-���v�c�p���a��jj�NV[@j��P��#J�*���3L�v�.�.����H� �1��T��ͱf%�͗с��W�s 4�E�/I��U]`�M��t�mѓM�j��f�	.�˭Nig+aZ����?��2�N#���7?�Gk8�H\����2U�M'GX�Ï�з��E؈XX�����n���{���ӆ��������ʳ.H�[h�+.��M-&�+A;������lӱ����M��pmR�E�
S)��Л���R��J�c��Z��+@��J8�c�N�Lqw.�c7j�	#����t���c�e=u����-�_�0v��*��ʪ��"�]P��)E��)��hRԤf	��ê=�J�f��iB2/-d�THn���F��)�a�R��En-�؝�D6�RmX���9�j�Ȯ������F�2RH9N��7h�e��t�_�̢5B��7(�L�sd
��t�a��jc�4'J���]�r-�l�E�z-at�M����������s��D���ԛ�������6����\F�����)���Ral�#�Q�nM jõt�����@=��bm�x��u�-5W�z8��t�0�SQ;bL�?�M�J�ƪ�O(ˏ.�ǔ�!��a�,�)m��n8��5i$2�۩*n
*�F�ݤ�F ���v�?�u������W&Q�كct�˽,XƎS5eHC-�swoc@7n�4ÙN�4!�3�uF]�o&��k��%�)��&�i*�uwA�����Д�D�a)֬urn��fٴ#P n'��h�	��WF��6�U�AĲ��M:M�mֆ<X �V�����ѬW��iV^���(��4a2��[5(�2jJٌf�k��l}+��~���pI�b� �!�%�V��2l�	ZM� eK0�:�
�;����E�ək2��5ҊP��w/�@�
0�O)(hMٶ���-4�m�jlh�u1���^J��f��4.�n��:��+i��9&��:��m[t�+�*Xn�^/I�����)tp�}n��F�9���=<���wA���ס���a��t+5��4�*Z�d4�v�JN1����T�.���!�ʼǺo6�l�r�`�U\�ia:�V���p��A�Qe�N2*X��멤��<�
��~��a'C�ﰏ��$|,VՆ����ƀ�\�'N�*�Y��S)��3�I�4�(Ʋ��H9wynh.V��VyĕY���+?k�����(l�����
l|�W>�k�IO*a;ʗ5;gea7�1�!W��E�VX5����E��Aj6��ůJ�6��(�4'`
�S�m,���]�f6.JM�R�1�L�݄���!(�
�̣@��]f�v,*���d��5��P՘N޹�6�MF��D(+u���̼�NA���o4�SbO􄃔Z�&�d�
������L��wZє5��O�nk0��Z�ICrJ{6�VX�t5��UfC@4��3L���p�XA��x۟�"�tb�ƃY�.;9(m"��B����Yt� �ܸmEW�ܥ2$κz�1�4�,��n�ڙD�E�M7 {��"�D��tT[��S)'[��ZCm��Cq�x�B���f����	��bb��l��a�⬩��b6݋w���3u��ҼH[����R�e:zФ�C�+�5s�i�u�9T��bG%F� !e�ٕ�݂%��� �ލT�q%�i�eY�z��m����n���f��IZ��+%MB�CkZsj=ɸ��n��R�5� �n^���r˲�����9��{7�vN�S�o-1�����`a���& ��]ka���V{m�?����0~v�W?�Ů�e��P���w���u��n;l�^ɂU@�f�����7�bٍ]�[r�f�"�'\�r�mZxqH�%��O\��n�)�5���@�f�QL�k׺���JY�{<n����|.�a�4���a�.<��^��Y�391p"&!���G���g�(w��G��~�(�?��:�!q��u�� @@��G]�+��������U���x�`��v []���9Y���P�
.�"]��-���d&=�-[P�� �lH��4���7U�,]G�2�p�X���/���+*��C^p쓪o@�f��:��������w5\$nh��T�w��x�'���wL=�uj�U��j�����d��|����Ye�/*�j護�j6�J\�f��Vijl]/vط���1�7I���z�Tr/�����t�6,��gf.ys��ҋ��n�۹�&ʂ�f�4�1Y��E�ݰ�lV�/�wAX4㌦�u�-��97i�w����M�n�3lN���m�I��w�W�/诱#J���P���pJ�2���U�$����M��![G	 d��q��j�WJ�
��7n��g
�$��L�y(��%ǃ$�m�Z4�V�Q��03A�ʏ^k�U0V��(Suw����W� ڎd���%*A卺��%ط�4��n&���:� �s^R���t�h3R�E*�٭��a�*M��h�/[T[{dE��JJ�X��5��A���̧w��JV��?dc�<�h����Uu�2o��}{K !��6��e5�'��u��!��v�;y��\�TF!�+j�Pd9�f��]X�kX#��Sp�,���K�w��:�]9GA�	��m���0ޢEg�ޑeh�ZN�PԞVm<j�x1쌢����á��������3Si3�惺��t@.W>�F��yY��
/X�6ic7.f��$��լ�ج����u��f-)�+U�ՊFf��ܧ+��:N��)��I��X���K-��U�$�9�
��L%�܍�]�A0$Qe[��Xf-�h;�ԯ����E;�D�:��yo����
�j����5�6���]��݊�^����u�v��+%X��̛��)3�"�2vɔlbl.��/��f��0ޏ),�NӶ*�O�+eOȋ
�����zR̘����=� �ɖqjm`w���6�;{�0�m"���˱���X�{����.�R����S#cc#��GK��ّ��ʌ ���[G6�e��8ؼZ�si��W��V9���m��.*�2�m���I;ױ��Ҫ����BY+yl�,�E�_�M5�
�t�N��NfQ��`1�@	�+v�[r�i��-��fs��tf%��w�>����V���>G�~g�D��!��'i*��UW�f
w:����W�����R�mf��u�(	cE
��*mm�����ч���VoQ	]�&\�+D
wMj�������`��"�)k��{�ZwX�x��w�L'Y���3-�Si"�)���R�D��vֿ�T7�F�ΛJ�v4���B��ƛEj�����ǚe�t.�9A,z�c&���]��`�� �,Q7���j�L�V����;p�/�?K�P���v��h��K��]��&C�B�hm��]��*�2��F�<;�$e^��C�9��(�$�<�Ca��M}t���t���,V?EEL���r]8��@z�R{�"(~�,�nj��[�g�Y=�$����E�Q��3eGET��7Y�{x�;d�J��`2Q�6#�	���H�����Q�6�]*"�;'d/�j�Y^�(�V�ɴXb�z�;��l"�k��h#��	�D�$t�o,�[� �(�������ǹ�9�x�Џ�W۾Ȱv�:�<��
I�ɄU޻l��3ˣv���`��%����&�t�����s��4���Se��>�{H�X�Vӧ�[aj�@����z'�O�Pf�SN��R��ɳ�V��ϪLv���4]4ܭ-��+t����E@9��=����6z�J��E�B2��2j��:2�īN��)����D*��Z�L�V\ٷk)Ғls.�2�7X��-�Q�Kj]��f������Q/��*J?��[��;���*ި��r�e�1[�8�yS2��WK4d(5U��ln
v��}k{���#,���]%^M÷�*�ofMHj�An�MQ�f[f�Q�tR���geZ��$p��<h��-Q��!j�T���/4!bG�6��ۋ"�O�7���X�t�.e�CX���Ւ����E�mf*����lܩ���|3��Q�CMX�Օ�Q��@�����Kuu0iض�K?י [ij�"�{�s{\R�RW
��'[�m]^��CV<ʷ-���n��OHb�^�J2�!I��n�qv�4�љX;��W�:h�G�#���/���c�|:~�t�*6��.�6����Rj��*�`�k�eo��,qui�1���=ҁ�mđ��ea���������	a9��:J۳&��5��n�F񌵈3]t��o�����s���鶻z.�g���2�dU��!�����񦳦��#�wX_7� �h�fc�$�X���h�[+�ߊv��0=����(���R��U:��M�(���&b��0����eƕs������r8�!�0f��ifud6N����r�"^>��sks*�9��y��Z,>r�<�N�p�ޮ�ݼvZE~7( r��E�a��蠺O��Z�#����OT<�.�X����=t�Vf걪�;�H �G�tp5����kj�����*�K���y���p�]�3;/MQ ���Ei(ea��qe��G�M'�gP��Pt��J�z��ͨ�U�2���<����ݨ�.�H��; ��ݚE�i�[!H�vtAQ���I�%�-Z�������o9���"ib��詠�aTX��@(EJ��5↠̹�{w���R��ΟQͷ@�%��ay��k#�]N�Q�U䐜y��[gqT$/,+���Mm,=k� 2�h����nL�W���(ԩ�ˌېU�YǃRK�	��-�����4�	[nо�sZ�%ԣE�u.��<uxJ�5j�0��Ӣ��-KCgpآY;�d2r��cf��3-�_�X�"<�����6�Е��O+]tQ���G�A�4�b��u��L��v�j%�@����L�eX ux��n��6@�*�HbX��0�sN3���Y�JǑ�@����.����B���d[Pk`>��ь�֮@,	���9����;%y��KI�Ƶ*��z�4�b ]9)���P��m�J-m��g�*�vG�ڡN���D���Ռ\մ��Y�0Ps��|�R�鹵�Ff87�n�pҽII@�0%��-����nnѳ���b�è�)9���2����
� ��,�w�W�5U�KP6'M���(�MZ��k�ی�v�:�!Z��|�]TB�
Tn^�� I�!�KW��՟��Dح��������tyL�u�`N�k[��h���)�CcGcH�ۏh"���;�Q�.�l���vr���v���	fid�Z!��9a�w0lXŽ�^K��V��C��G����?�Om����4M�� +�����e�rK�� T��G5�^��;]��#�-��x�
$D�9�M��1""��=�����4H����9;����kk�b.�q?�wv)/[О��X#v�f���C ����S "Xhw`��n��yyCCܿԝ�Kv'�������ऊ���[@�)4��OV�F���;�̫È&0��ŌHUٳwz����k9y��<��J��ܛnb�hLڷ=��]؋��hx��ۣp�u1g	[��Z�s�K�vE]m��4�`F�
%c�EBh��2�֟ĺ?���~��*�V�7��p�3@ ���hRneج���vN\�V�V��2ʁ��D桤��gn*tV~ͭ_�b����L���Ka��ވ�Wr�Y��0-4��2�9��,��W]m4)'�Z�{��n�r�*���m-f�8 `�5�z�j�LH�7�G^:�v7��1�H%vv�B����AY��@��,m�5e@�O�ORB;j1�m��r��A�ET��q:�l��L^eJ�{�1�iӵ34������1l�){o]X��Dy,2tʰ{��D��4�]���A��͗aPʴ\�,�0�f)����v`bV(�2v��s�4݇�k	�#VFO��ۨڑ�u%T���V5,9��
Jn��2�7h��ݺ �2��vά������u�����)p����ТHon��/4n�k������.�-�V/��"I^;FV�V�m��om�e�u
�<f��MY��p�ӻ�Yn5}��y�v��c���m�BՇ�_MB��ҧc��{ћU%ś��7r��{:�~�'�c0>�.��d$��XB�\D3U$�����z;z^�6�U7r�>�[�T/ �[����P
�/����F�w���h~�&#XPL�#$jIa�J��5U�V�&�|�3��(��TҭUTڪ��(������`������25U[UP UUU�UUO*UR�UUUUUUUUUUT�\��*�UWW*ґ-UUUUUTQU]UH@;UUH!WUTUU@UUUR�*ԫUU��j��j��Q��dj�������j���jU�UA
����U*Ԅ�I�UPUUUT�l�UUT�P]-UYYV���^j�'5mUU]UR�U�V�`s�˷mz9+/e
m�B�\iL��M��K���e��xų�n�3��#B�c�JnK-��:k �P���C�B��ij��a�W���7h�����WcQ�.9���q�8��F�\�<�nL�8���N8
[���]���q�8�=��9{�]vF�c�tNŨc2�6���2i�.2!h���n"Q�1��fu���y�.�XYl��Dn:�3�������5�.;Ls��m���*�K.��2��6_]���u��B�u������69�/[�tkzk Zk���k�ϔ�:�.�,��p\�D]�&[��6 K
�`mHِc��gQ�;�܉�Ixy=;[u�t���ڦ��>�:�E83u�8۪{mq��.�z�hK���x�>���|u��:��¸
@2��um"�ԣb\��A%��B�B]q`��a���XXp���[�CY)�W\���=�حs�(���`:�]��<�׎ڊeyi���h2���^D���\�=�utPttt�[���:�亀2�kbRKR�l���f�]�c���.�
�]��n�����t�1��:5�H�p���7t�L�Z��C	+��2�Nz	�q�c7"��^��8�)��<��s�
[���֌3Dz�<����gFeDl��ε� (FPJ�J�6�hM��M�em롵af�C$CV�.݉s
�P��[gqm6|�6��GI��m�U32�\��:��P��Md^B\	Cj:�i���2���)�wy��\�ۧ�!��жS�=pdm��nn�UӢ�r�l^�,��'�:ڸ�K��5.���1v1]8����q['m˥��4&�^̪Vl#�)fpe�iӅ���5��`����81٣�%�#�t�Z}l�f�5;��Q��]�F7[���"�RV^	����Y�����˄l,&��x���ks6�͠��]��ʆ�0z�:�����㫴i��5���L��3�l.8��jA�ս.ؠ���.xH#&^�.X�ڂ͓EDJ-�\��l����!͸2Yu�/���a�m�'f�=3CѮv����!NSNRuqIy󆐹ݤ7�8�3�&�n���ꥌ;7`[�"p�ԁ9'bN�\D]�׎S�s���Il;ݍ��l'.�=�q����b��&����n�;ta��և]{gYB���k�n�KRє�]<�Mpe��5q��Ys��J�,@ڞ*����h�M�$>:wod��׋]�D���gY�H$��]�M���[mV���1��n�rh����skJv/^� �&"�v�E�@��M�@�-�7j,,tiIb�p��
B#�K��Pb������@�ViHg$z�S1�2�=j3p�!�­l�P��n����FP.gi�9��JnݯGZk�s���i �W��q����f#Jl�cc�f������Ǳc��Ci���.�s��3b3u5r�n�n��Q�����k�W�V���q�{@�W��sѲ�en��إ�KF��^�=��=�U����Г��e8����Տ1�j޸��tm,'([�;��#m�<�+��ܓ�]s+�!�]��Xsk�m�!��Hм���F��.�y�����Ս���d,�`LqwG[I뜼���rUղFsn86�k'c�ʗXF�u�Gs��cF0�.��v)7�fL!�9f�0�r�n5�(����VZ�]f����ԣa�
����%���	n�	�	y-n- �^h���wAS�j���8]��Kh]ۍ����REՋrTj�Z�2�v��䲱�\��ܥ���Y�mu:�i,��	&��^]�\^��:��\��.32�R��4pd/l�l����ďDHH�3�������[��Aw�.�[�T��j@�jkl�	]�n�=��pޞ����"֤Qm����kb�]qk"-��&�2�B+��Բ7-lr�L�y��������$]ئ�W#({���n��k���8G���xB�X�T�a1)b�Z,i��ٺ��ڻm�������fԋ��<�7�٦�ps��6�qt��2zfn,/U�6��yC1����kV;2�L�\�e�(�J��v����\ѷ6B6]]l5%�v�Qf�Mԇm�չ��nT�=��F��֥�8ݪ�$w>�\r�,^����n�1U������6�hZ��any�u E��ZŖQ��]Dx�ɦ�V.�I��i�x%&��e,GZn�֧<TiL��Ȟ<��|�m]�.S����ڸ(SKi�P��l�R�VHYJ��1�j��ۉ�"
f�k�CU����&%�C1����������nۙ��UԺY��ӭ(�u�%$��kKYL/i�����o'���9q�t1)֪WW:3�'k��[��Q �(r�: �mv�Kl%���hJ6��봍�[.��X�B�h�K	�j�\��g6�1nQ��4 ٥�m3�����K�s��	�a���^�sL�/�NŖ8(����b�Ж�\[�M6�R�mg!$+�����r���u��vAe�Ʒ��lù2�6�TN��5������T�!;[��(v�:٢�*�*�7R�-t%u1TN���m֑���۵��Z�GM�uS7l+�(Bvۇu�uqϊ3-����ް��a�l�fL�lhW$�g2�ի�<\Ä���h��]�D�m�����f�l%B5�1�4�lWf�M(^ڨhCB�!1�9"��.5�i��F+�HP��{S�F��4�V#�3ї�٥��M��l1�h�&��:�1�#I��̖�&�k�iw$mls�`�\rG1���#�w�usۦ}j�7U��� �G�fY�u�R�w��c�\��lL��#�x��b���	����5`��cu��.4��5d��m��`�ٔ��F�.�Br��˸�kc��Ż���q�1������(z0���;A���e岄�����ے�ku���AP٫��=���'9X���)x��;�k��qs1ط&'I�]��N��d�)���)b����j�Mie��L��(Ɣ�%����[�a.�֌�XmBn5��J����y�)���٤<�!�j��1rAa�������6��@��Y�dm��C,�v	��;Vz�N��!�,���5(h��5�+�����&{Ln��b�4(A&��n5��0Зf�mK/.�'���vx�<�N����s�p�=]�C��nٻ5:(�pP)�%��:�f�cc������;i�.Y�/Ki�B=����n�i�����X܉�c�D���!����v��Q]I�㫒;�\Y��uq�k7��{Y�;n�����gGk��m8�"�(�b6�[]J\	lr��s�ff��f����p�%�-�����8��D�6����b�X�h�n�@����2R���l҄[�6��@0)���nH�L�Q��&�.uf��T�ņrh����sl���	e8KwK��H�AJlE-GP����G���;�q�ܦ֍��;��X�fޞ����Rl��[i��Ԕ&���8I�9�Mnc�ev��&-u��`ܻPLM�׀��k6�;R��a�^���e�M��̥�b�a�x��hk�N�u�����К;�)����������P��M�lf����ǘ��4�6���G�t��[�;E�s��'C��4��@�lk��-�j��1f�b.�����o8L��gG\C�N�7AE�ы�ktOlɛ���z��[m� �t��fHQT`ꃡ��ݛ�]B���[��cXM���wRЂk��
���#4֚�ie]�v�@�NM�ݣjn\�X1�wfKnvV\�n�ʋgq� ��X��Ǌ6`B�a�n�)A]SZ��UAj��i3&B:4*44<`��\�xq��V�J�ˬ��&���K�l#k�Yv�ˋ�KL,L�6����F�k9�e����01���s뫋�w �u�Y�+�p	7a.v���YWKt�����������m�C�qͽQ֗S���a.�G^*���<�R���Kn�:gb�Bۦ�ۖ�,��Z�ͦ�܅ݍ��5270v�r\q��^�6+���R�αHVR�	�X��FH��@�!v�C��z�7-�m=<��A'���v�ʁ�nxbۥ^9�8�f��������0�y%0��uٞ�O�t���[��q�v�c��W;�� ֤�I����Q�Sd���K���ɉeC&��R���A�΍[��H��6�i)[i,mu4��vG@ �D5!���na9���ַ4�+c�{0m�3��f��rH��!���j��;���R�r۶�ƺ��J�W!]>^Z�{ułvő�Ѷ�Ԣ�׹�W���X������6�C�l���b=1�`��Ҙy��<$��T�y1��\[2�
.y�׭�j�mڠ�^NH3t��!ۂ�G]q������w[S���;�e.��[u��ɮ�38��vٳ��NL<�f�2�bY�9�x��`3��^�lv�sأAa���Xެ��Z�4�i�#e,��F(L�*狻j��:��tv�kŧ�g����OH�B�ত�.,j�:��5Վ���O:�gf�h����nݑ��=Kal�4�bejˮ��HV�J����(C���L�t�s���[�i@�:�kI�XJ�X�c���� �V�]�n��m�.�[g�	��ּzո�
��:�=�jL��i]�ѣ����Y^��um���CB��$��wwz_vt�'I����{�t�����:N�N���g��I:N��.�_��~^^s�i'wI�'N����t���ӧI N����8;���;��t	;�t�'t�Ӥ���:t�g�����U��ȿ�ҿ��G���o�Ʌ)̲���e}��>m�R�O����&�� �T�W���By!(�R&�s��S9�A��}�ךg��.������^&8�u�x%�����R������t�3{a�u�� t`��1��Ɏ�ԉv)۔]}�g�:5k>�2��b9��y�������B��<��ԉ~�(6d�U�5��*�1hj�dHeNn�Va̅{R�)�u+q��JX'*v:�����
9�r6��De����S%���&����>�
�>ݘ�X%�+�~��.�V\�m�+����Vތ\��c��3��`�
�]4�+�e����w��[V���ٚ'l'ݍ�6��%?]����Q����+�w&�1��0z����F�^��u!���s�Zˮ��=Ű�};s�v�~qc���>�����E�[~�,׵5��$׎��ݙ�n<���_�+��E m���tVa����T-���1���Q\iv����s�[�SO�4F��]#W��.��I�����R�4��[lU�+�p��R�I�+q�����؏�,�#�]�w�R�)�^!r�Oq�-��tL��FQЛ7U(S����t ��+Yp�ܑ�ћf�v�Φ�;�-���=����4OR4����u��3m4��x7�dD���-��.�vv�m�,Ie��^0`�n�nB��l]�..s��nP�둓nۍF"��H�bfb�kV�P�FM.7��v�-�=e�$u
ݍ7Rb�ŉXT��R6$�sm������sP����'`����)��k

�(e��^1��%�����5�V:�{ �OO�������q�ªa�wW�}�3�a���!��cuRWw���B`��*���k�ל����J�(�{^�/l����]��JX�� і�`��m�%7V0��{5���Y��B� �b7/0,�W��'�U����zߥ�1�k��\�=\w}/�t�B"!@�#B�v�M�\�s�f�!Z/����U�[o`��G�B�L�Ý��d�S!���y�gyc���+B�X@�M�⢭�3,EȳuF^!7Y����OeAjm�e�Ջ�|�}�~z���;�yD��܊�U���e��h#f0Vk�
��w^�J���燻���p�G}�q~�bzM���+:��o2���Gq���7�@Ω�Y߯FL"B���E��e<�4-��KsMd���iu��c�rp_�����X�1wq��0�J��n�wf��1��<ͩ�C���P�72�&��FS��\$��[;l[��WJUX�����;z���<�*]�W�|�Y\�����Vy�$_
>��a$��\!mZ��:ca8�EJ�]���K��X���M��2Kc2CY��z/v��!�,�4�E�J(,��ɛ��x�ͯeFĭ��_�F�4TY�sj�	��8K*������Ef��xY��*)*Ro�����0\��ޙ�ٙZ=D�NL����X�a�{�fzt���w#GV~�Z���{o,��P4S��[p\u��^6dC��Y8�gf�s���z���d��̒�����g<֏�se�\\��	6��43щ3��r�V�P\%) n�Z�H#�S��1ݪ�킘�����0w�9,��sle����]��|��z}��_(������:�%X�M���Ӝ��O%9&-ܻ:їY��>��>���|�i��η��/S("!���eT�sL�j��C�e�ٙ����n�o��Y*�a=�����rm#����B�&�ҿɋ�IV{��lF���l�Y�Â"�̭؋%�]}ǻ��>�]`���*�~/��k��*|��ǒ��+&�5�um�L�p�KY; Jݑ'RWf��v=R���nrj��J����8�GLܔj5m����wfN��D�p႟�<�*3u�����c�5p��f��`
;�ۭ��Z�t�\4�^�W����fu�]l]�54Kh�к�ʿ��O�8�p�,5s]�J�q4MIo��mA�y~�7�:)���wbMR�`Ǖ�.����U�Q��P1�
�LB(l�Z�/����wj�|�ڲx��ܧ�o�>��w����7>�ϱ��:aن�7���U�V2���ʭ �+�PhA|�9C��=&���kV7��"޸��8c�����3�$��C��W�_3�Z��W9���u�]8^� �8�f$��P�≂�����Ǣ�{�A!)�L��8.�x�ۋ�\nl%z�a�di�]7�r{\]@X6l*�5�v���O?p���fLV��,v�x��,N��L��%ݽ��Qh�DsEι�Uc�f�a�U;W��g+
8�y����^��*%za�Qd�qxmXR��z�N�֬o�{9	��2��8������h6!7�΢[	槷.�B��T��xNJ�i���ˬӣEp����%E<�[f�.���5�����1QOo���ݡ�Y5�f����>�V]�yw�x��ې��3�V��^�
U��[;�߫��oIV	�5d��4��'�1vn	���x��j��F2�����xq��MQg=-�?���u/�qq���n|�2���j�8 ��ne�J�󭌵Ug�Q�a����"d�	^>Xw��:�ʲ���u���}C�ӎv�u3GN
~s:�`f�a$��M͐}o�_仹��>������7ٔ*�ε�Ѱ�Ml� %���ܲeڊ�%��LhU��$I4������]\���>�d27<��Zvӆ&u$���nXJ�'f�k
���	���fLg�7j�jq��f��pP����ݳ݆�l��
�<<����g��^��ɁMվ�/UA[��v�hi��D��#�<]hޱF(鱛��M�)WުjeXz��bN;�z^b��3�B���mu�f
c�JX��^��^�aA	G�|:+y�v~Ҕ���rok��ͧ�[(�]	Z��gz ���o(^�U�5�j�s�B;�7�fJ6����e���j���'l�n�4u��(��0"M�H���I$vsM��뉞4��7�0��8=F�����S�����V������+�)���sګ����=pزu��R�0�;�v�S��q��!;4����K�m���Y��� f��-L�ng�l�p�vn	��oYy����ã]���mt�%����m��a��/h�y��q�`9K��؈1V��ַk\A1�8�,&r���N��m���𞵞DCW�F{>?�wދ����o�f^f����bF�'��A�]z�Rt�0��I����
gl��[�x���K��8t�����Ս�pcS��ϫ�°g������\AS�!��F��@��*{+�
��W�}���:��+��ğs��;gr/Gf�C��<�g���㳓	m:�̀�Ԏ	�H
7��$kwys2{O�q�E״�����|k��ԇ���+N�A�6d"&� ��fAܙG$�y�^��r'�����a�R.b�{5p*;w�&>��%��ű	[���Qf,iq�P"�JXy-+�3�_�y-� ��h1�,q�c�?^�'�⟷i_i}��R�۴Y⯗�x&�������3;%��� ւ�CB�X�1\���t+q�b�0=�
	��ۙ��cN���Ur���TWY糜=7kP�;�����Kzt�^��4%0�Чi�UW�{Z��g*�g�z�׳��4�`��+���9A�{���u���@��Ѫ�Ǟ����X@�
�����*��F���|���;U�u����;0�c��S$IQ�YOL�܊�ƕb���c�cpR"�63R"|M;8]��_����{s	�.ɹe7
$T�&��]�V㡹�:w8�W�\&���E �lf��v۾6_�f�]�*M)Mcw|o��Og8S�&=���p�+v�;}��,20@E���ܖ�A�I���RR.3�*m�������mT/�'��g��K�l>�+:����=HG8�o��Ұn�%�a�(��vl�º^�y��k���'}�P���"��;��B�,l7ٖ�*z��1U�:-4X==�����N�iR	���e����ݻ��k&�OƽxaGm?˓H����Cv,>�[%����;O�v.od�{"ܬs$ø:��.H�
HP�TX89�W,:�n ��mЛ�GM+�޺;Ң���s����o��+�^�W�go�ER�jM�4Ey��kb�쀚A�S(2]��^��ףrǅ籣�ʶ�=�V�����GC^���WIQnf5-��-��N���䠢�t�A��0��	�܊��˚�jF�g����/3V�񌝕yu��������=1��{[mO�wm.�*$�
�Vܖn���h�l���.�l������<��-�=s��h4q����]F���֭��г\m�2�\�zs%�8��j�{u��r�?K��uAj�
����+�X�HW]�km�د�S�z�Q��I�V`�c�����߬> J��t3�=�-h�Ͱ�z^Sǻۧ�	B�<�s]���p����x���-�;Z��vP������*�5n�n�v�\4r��d��hoE*ub�v!Wڪ���r�n)nE�Y_8�6D���jd`��T6T4ZF_��N�G�g�Wb9�^x�\�lP��<�k��8�`�m���dK��4vԥ��gt���r�&�R�y��ɠ���o�ks���s
l�;���v�r�Emu��´�p�g�Ƴ�>{q�T��Rq6ӆ6a ���qG2ު�2��oa��0b�ݎ��k�4���+V����	e��J9
b\�c�(�y}���V�Υ�O��<e8,�����c�c�?n��Z�|o�oR��ҡ뽡�/��pu�xM�$�+�%4o�9#���4HT�?��{Ke�n{95�^L��Z`>Pa��f�2�,���Mwd�ѣ�o�w++(���4Ջ�6�4��������l�k�������ז〩�^���Ww�3˲�
����N�a�+�̳X���Q�
	�ʂK�:�f]���_�]
���\;������h_>�r����և��]�F������ ]�������g<N7`�ů�$]��-��X���}f�O��j/=�{�A�Yo=�n{��y86�~��hz�������s4������|�/�"ri��r�/�c3�PM�S������W�pWj��#n켏�����3d�p��]�rʕ�E*F�XVn��'I77�^��֧�D~w{(��o���W��c�\7}�'U�Φ�~�w9 QD-f߼�!�;�{{����(e�����3`d~�ҽF{spÞ��*ev!�#�fW}r�4Oz�eV-�}������+X�����cV�GU�����M-�ҫv�[�ې����J.+Wש��;��f�7���p��,5��=Pw8[�p3�C8\�m����ni�ޝ�$��ݯ��ذ��WNURս��vԮ���<��m�,M	hY*�
�.L��CXT�o�
���� f;���I�׵�M��oc�o����G��eGm�678U�p��X�Ѷ�pd��/�6�:N����t�:�m�ˁ%��Ï4%<F�]��X�%� ��I�F�%�2���+MZKk{h���&a�iT�CH�X���i����59��x{[��Q�8b����ȑ�@��ٔ���ZM�ѓ���9��Ś��){K�Mj�z�0�tf0�0q�ڈ��=l���E�
p�p�Of\և<� �-��%�r1ѯ�f+��5S\�ln0�BF�4��^D`]Ѻ�Zs٘/ܥ��+���3w� ���aeq��Ų�����\+�u�X��cet�WX:s\*�N\��}ĸd"I��ת�<�gKLv����ت�P�9�cZ�]q�ٿ�]���be��Ǆ�����i��a�n��M�E�V�wx.<���ǜr8�xh��Z�:�Ļ!�Z��<�L�Ԕ/+�P��Uа�L^��\��a����)e�t}��:��V熏�l����"�:���^��R���B��e�)�	@�ړ�6.7��I�Vd��9h��_�s{N:}�¾gn�m �ԝ�!Gq��5eK�`�ue��7�v�EEp�ٌ)D$��Ƒ�pL��۩�7����r���uO�yM�EyL�d�y����^�0����ܗ�3+���v�B?'T]�^FL f9�c�HfPF��c�׌]qf�9������y� �p���q����>v���dW����h��܃�y��ڤ�;ŹR�W����_;�Z`*ZՇJV*	��+�����5���VAL���T#f���CaU��{r��+��a����lQ��'�=�xX�0��s�;�*�!�W"�f�U��z�K��odG/T��C]���������Ҹ尬�M�\poK�zc��z\��
��� g*�2�4f-z݄��={�^�֔]���: ��tK�"{/;���wf�5�X&�6z��W����H'?�O+r���3�=�pS�jn�Aw�k��I1�hĲ)alK�'+��Ri[�ɑ>xQp��o��2�9]Z��bVE.�����ч�8�����O�R�B�p�S���]���G߷�L�z����h��d����] �t��k��u*]��/n�}���+�^��N���jγ����l����Q�an���2F���_�C������Q��Mr�Qo
�0��n���4�6��pS�4�5°�ѣ��N��ڹ{����PZ�_>ܼ��1��G_>+��B�98�%�, ��e���Z5�%zo�1��W�ۡbύ�9��T\���K�͸�����Cl��(c���5P&��p��g�
��	�Q1��s��&P���w�~�rma/^Z(-�"-n�KE�9���=�k�Ƹw[±Ѯ����|$K�.��ө������;b�ԩ��j@e�
�Z&�c����ha+m�2�i�$��)T
����V���kj�UU��
�*�Z� �A;*�S�(�Ӡ��p���A��b���a��XG��0���㋮Ր4���.m�R��"R���S��cX�BĽS˔;tmɨ&ָfy��)1�3����^�Zwt]8u�<�X��&�L"ѳ-�P5KD%fVX��.�6�B�grSϳ�d�:z���w�m"�ڮl��
��/֣���W]�M(l�����`�c����h����w����s]�w`4XֶZp n�]�ٍ�M
��M��[#f�m�X�@#��M�p���@8^�2�b2��dN�W!��C	�jU��s����(,n�]̀�cX1M�4�.;`�XWi�,qYԈ��\���^���!�F�d�M�.��l ��")ݴH �My���b{bݦ�rt�
E��&���R6ml�u�i]�c�l<�Y�oi'��2�Ő�57�n;]v���$'h������H�n;]��7)s��O9;t�.�*,-�j��n6��(�C�8��'`�\�+\�am�s�nhv��5�k��e�ʼKlr��u<G[��m���-n���[�/N,80s��#�e��4��7Zs���6pJЗuf.`���H����l�I���d1�'���7	���D�\rJ7f��h��ƅt��i���9��,#���)��㗎���b�ۘ5�z�]=�̥أ�v`��5���:�V6�݀�c����`B�]�@��6V�tۓ5�v����`�];e��f���/s(u�c�IK�v�n^��z�pj��#<�93�p�:##��\�cV.�78Mr����Ye�1R��F�1�$ԭ�m��Mt\3��l�΅nnnH�d�e���^�;Qî�LCJ.���(^s�Ǎ�n�vMc�d���N�J�Љ�#7s��j@�J�Y�-,3c(��@4V,JXj:�(��R驇UE�=�]�k��Jn�]��J|∶�N0��������}��n�w�"��>�"I�N�C�nl4�,�IY����r�]�6��g�~�����_���:��vm[��oT��㇮�j��X���f�[N$� ��p����j��}Jc6�bU^Lќ�Q�&�2H�f,�ᝮ���v	���]�,}l���˗�����[���h��[Q(e�M�����(C���<F��'^7�z�g<C��Y_���E��7�s! ��Δ��#7<{o�d$ij������{��ޙݲwa6Á��G�����|D;�O+(oE�
�e:����0�a^���oK��Q��q��[[{|wYr6�No=�*��{Û"S�kyFN�]`�2������{u��pYe�\�^ct��׮�yQ2Tq��T�\��u�I��{M���:LP����,IBL!z�Fq!���{"ņ�M0��ܽ)��s�4��P
K!Bi�^�=��Y	�pPFe�x�k�V_X��$�Y�MY�C���޷ �q#����}�����R/ٗ7�c+�lrf�s��>;�H��p@��V�~ �0�=�������VC1|X��3�>~���Ց�N�2M��[\�ՠ5��x�"K�3Z@.�H*�"H������wC����d܍����fy�^���3b���R��h�£��[���8lJn�����3-�w��5���{5jb�T�"���H7%kX[&s���*��M�E>�uӝ=�C7���|�;��
���)���;=^��7��t�?���3��~��U�M�;m�oD�{t�L\"�l�ѯi(�&[Ү�-zJtػ��$�$���K)Ks�e��ӧ=�,i���z���s��.-o�����U�Mm������y�of�hB��&�(��K��~2Ն����S��:�s  �4k�È���wUMF�F��f7*[ơ�>����벤�H-��D��ĻɎ�V;��۪��H<��f��z��(FAwʥ�7uq���JHHA���|�ͨ++�2v���X8Eў��/�W:��26��=^�Oe��!�~*�{0f�(lO��g��FQ��Q���ˡ;�&����wZ��f�s{A���F���)3�䄂`���$��`��K+u���ml�P$`g�>��$d���w�������
ά��Q>Ƈ]�8����)�G�W�������n�o�A	f�Q7vK�Z<["�\���>�ᛋ\��G����Ϭ�
�
��og>�a�N�W|��Q���g!\)���{<.���Bv�o�WH��R���%�a�G	��T^��4�L�$2�����Xq#	.Vf�N6u�E;�o�H?���(J��hi���3*ØNu�iv�BdzQ��M�yٍf4��md`*�5J��ļX;s0͏OW�mv�^�������Z��� sB����j%-~y����2#1h"I�����zߖ��ǡ�d�e�%V���)76aOq�C �FZQ���]^��*�j��h����S���e�^��'h�]���\��ƴ�l�E
�yבU=�&l	m-tO�~�=q�6��ō�](��9�/x��/�_c�̢Ͻ�A��G�A��Τ:��N������(������O����iS}r�����h��L��*�ĕ����v���Y{�+������Ӣ��F�t��K�n�k����ω r��β�:VC4;<�)�u48P��>��ڵ�}'��G�T�媡���C�]�b��Zʛ�oʄ��E�X�!W=yYƯ���l�l]��+�1>Ţ����՝~x���/'�c�|��Jm�}�a�̟[�µ)����:ωOuΟbyy9sDa2uA�m�ފ7nW84wwXaHpƠr�wq�֙t�Y�x�L��� ,p^ksw{�xu��ϡgKC*,���n`����0٦@R��w���=u�Z��[��s3J�p_�����}O�WH\������^�Y�Z�V�����-
κ����b^�J{�ǚ��N��$��B˥��ʙ�=��¶�m�OlΝҌ:R{xC������;�4�H
xE�Vr�)**��>�O��~孪�y��]�n&k�4�ݢ�;Ksk0@�#�^
�ձ��]E�;�n�����P`<s7<���j �a5��묾(��΍�q'ݰ�zy�٦���-s��`h��]iؼ=�[�� �S�����ܼ8���:������<֛����n\��׫L;z�΢�a{������=�i��u��ю��L8��|��B� h>�;�\b�I�s��
�0Y��},���vF��]%i~��+n;��E��7��f3�sJ�-�t�Lͅ�w���ey�P,���\�5�<|��v{d�(!k�8�y�I;�]���~s�AE�^���-mg�}�z��m&�!�T�9���n����}*)XN{҆Jd�kg(kބt$SE�申�/&���]�ڶ��C����nl�M�I�!&�U��݂��Ƚ@]���UϜ�JZ��3>2��WT=dx�.��[z�o���u39�э��
$*������ZB3����0�o�Y�9zk�y��e(F�=��Lg�K���{��m�'E��i�B�z�	ʢ'w-Ć�6�`������ Gp�aY&N�A�'�J�m���L֯m�6G��7�2�pe��ƪ&��1��;P�%�ۻ�D�-j�Hk]�d�ﶝw��]����b��,<ŹUx�od�(4�̀�1��4�n���y�:u�MG;�d��o�K�{H���}��Y���>��~��M��&��qNdQb��<u{����(0��0��¬\������+-��o�Y��N�W��'\��yŜ��������ϔ�J]�uz2oƍ*�ps	6�̽�澗xOF'r�� ���I�v��Y�����`k1N�� ��K�/�1T�LWr����gw
�32��Ř��T��X�K.��P��#�+\z�QUuj*��-4{���~���d��Ʋ�J�\�5s�m�؄@�];B4���7DrfB	Ɉ����4��f�O����wn��.��7�����@E��H����DȞg ��<���j�EWh�'L�̸4,���Z�cwc�E�����
<s�K����Q��|A�D���wo�q>飃,�r����W"'c���i�y]����K�v��M���F�z��%����{3�����|�[�Ń����\��<��(8p��O׮B�	樉�CO����	�pv-q��A�s��¶�ni�Y`��k��(�AKQ��k܆����y�����Gjb� �.����.=�Xy?;X}Rg�����z�2�6�c�e���a�`A�S�&*褑�����)�^o�U�"䩔��W0E�{�[���S>�mr?}���&�X���(�7�Q�ic0葧=�Ԏ����D�d�ro}|mP��̲&��qT���Ywo�V?I��dzA�T���en�����ǖَP{��uׁ0�\����O�N �`2!�y��=�P�E�t8s��͹s���k�,ƻ���ݻ�4��3����}����"e���^�y�@�Qm���FD7Xz��	�Y��[m~�ƶ,*d"�
=��m�V�W�ߵ��;5�31R�U��}\���;>JF��@�'��Y���U��ˀ��;��R��[����x�4eujր���0��%}��WG��Ƙ�/��뛯`�|�.\&�~��P��Fjd�[ ;*�!���l9���	�osrа� �͛��k>�,�'3�3Y�4�9Pg&5��r���E��倜���
H]�kŭr�\�.��-ɻ��n�zi��p�/ٰ�k��}2��{��^��aE�9g����jiO��R��ot��%�̷�a ���s�1ݜ�β���#���W����Op�Z�m��l6�<����@��᧌���ԯ>�1���&0,��Ϻ;2�x�aQ�JH�V�;'�/i�c�^���wI3a�~����8�����+}�m��R��g"�QƠn�
�[EDPƽ��e��=�T1�q�~^��h��ڌ+,���G`��2n�kQ�6us���rb�X&���z�C ��On�4 �������ڞC��/���2N�N!��|�V�)��x$�8�}|��]���9�o�iaUT��V�f��*��~��=\�[���u��V�\n&�]���Uhz��|��0��ero;saZ�D���4�|R��d��q%�l�CZ����GS"�V�;��+�uT�۸��v6�GB?��;d뷂~��`}%�ѝ���t7]��t�ࢌ�n3(�TS�T3��5�����U�TN߸�(#*�*8���*�ǹB�]��A�u?2ߵ�W��_"�Kr����˻z4֠��Q���H�8!�Ϧ��&���Kޞ����-��	�)�ә��W}>�i|H����=��%����l�N�v�>O�˃�g���e��d����p���ml/>ݮ7bvef�j��U���W	X8���_��о޻'�焀�<�(�:�\��7x�2?u�Q^������k�{��^dno�H�YL����z��&Ɨ��-E�����fmb7t�d�z��{��V�ҧg�`�d���^@[X�앗`�M|d����tn$���)k�e�Wx��ݏ��ByW���E��+�u ���
��i�wpH@E�%��:� y��mO�I"
�����2��ԡ�-1Өő��#΂�+�{b��\��u��ڝ�ǌa^f���������͔��!P��q+-�!(�_1]����EJ�/����W�L~�EuO+w� j�3���Z_�&������]]�:p{����ϼ�o��Y;�&�^��d�����������w6��tx$eF�UU�#T=�jH�ϋb�!i�qI�� ��r�9����@J�Fz�S����m�Qh�۾���)��[�x�yn�a�:ά�n�7N�����Sl�X��\Y��4ӳpy��Wag�|ur|J�kGU�IY�i�;���F��n}�x�I��9���`m�z���j����aIu�fi�k*�A�f�+��
m G���LCM,˳f݂����.�ղ�v�.�G	d1!����"��j�b�F����v)���c���'b�L`<�$��w(`8��3�Jy��B*3="�ݜ�Z����W�Q����mKv}�"��ť39�w��]� �hAP�R~d�u{�`���e!X����A�8����8�^I�zfo�C��p�6m��\����{$��u�1�Ƙ����D4���2��O���E�V��x�(�$x��
������Ͼ������#�6ٺCGUb"�Ѵ\p=�u�<��m����6�Ok��c|��9FBэ�JU�N�����~�W�"yC��^��+a?�+z���Z��Hn�auy8t&m�3���p�6�T�fٿvzXނ^���ܸ�1�2�!-�X�g2{(pow�>�0�a�J���H1�n�:|�0���P���� F�<�0YE�4*8=ϖ>�dd��"<!��J�3H��??��g�B'�,Ι�>�qb��y��K�+�� q9��j7�g�̥,���Wη/��z��S��qSat�
թa��8c��L������Y��}��O��<�l��`<}ҝ졑w�r5��ȣj4Q����ף��(��(&_T�3�{�p��%��i�Ur*��fK��܃�����:��wʈ��7�>��cC���-u�n0���`G�ygn���!X��(eܕ��%��x��:$�^U|\�SSՖ`Z-ŹS�RڃOI�n`䦪����
�2��l�0�u���@����W�����K����דl�>�"FB��#o��އf+�m�[y�����Ư�e;�)kb���,tBbU��۱1U�z�ȳ���=����5槰:3��A�R&2G�y�{ә�R�s\ۮ���'��I�l�L߈��{k�9��cF�oUw̨��xr��?]�y ���$�)�5$�>��ڹ�dr�<t o_��_{fj��څM"�/��s����v�vxh��t���T:~Gw��f��Pa��D��I��2�>;i�H�WJ��p��k٧f)�+$�U���W����q�#�$
���*�},�!����=ח���kUnzf���/�����s�n�"� ��jJ����2�e�c�y����(L�׼��}q��vU{d�o��~�@t�H��	��Q�7��)�g�i���B%����f>d#�F&	^'S�/�j[�����C1��[U�M��hm�����"��]�E�х�����̥�{�Օ���=��Uҕ:f'#(�սݦFڏ-l����>�3��ˑ`���&y+�t���ܳ>"c�/G=x�~�����5�ѐ�X�m�;�-	`&�:�a^���R	&�)��!g��;�H��;��h����z�������G�f�i��������'<������rTj'�q��`��\K�If>n�k��x�W����I&6�nZ��α��U���b��/��9�Wv}�n�z�,�a�'2l@b$A:̎�uW>}��V��a�c=��;*�yN������Ujn��s=쿰~��/n�{��6���>���n��`�J��;(���ʐ�u
��O��k�}�\�����B�H`J�t���7��K�NS~�'�J�L'��g�����{u�M8��9�Z�i��v!W�'�Q�@ (Aɔ�����ySyNj��C�,n�����������~n���ђ|y�GvS�U���f���g�X�}:#��x�U�I3��Zv7��,��o������Y�t�54㳀4�s���P�*�3[P�]Uu��sI�-@���ި�'{����:5����?x��U�wKlB��O�P�&2X�//��&,G�tLP ��0�.+�'oϔ(��MԢ�']n1�����2��-7�4D�G%am�&��Q���	���Q%x�N�۞�)�*���������n?t�Km҃���VFl��qa��~	���?m�:��W�B�_��5����
�:�+���$���s�"9ɣ�ۛO��3�D��U͹_j�j���ՙ<��9]�U���JI�5ڃ{�uΞS��%!���vi�^�U�l#��pa���p>l��. ��uU
~���f�{���JY�P�7�A�J��S�Z)����9
n�Τ���CJ�H� ��c*)���7�j���nf��|G24l�e�/T��l�um7����W6���dP�v�WMn��������t�*[/�v����!vJ��o{�u�S�4�Z��.��=���V�����f%��Vs�q�����Z���\ع{� c\���k$I�VQK/��Lθ��*����������$��\��\��I �x�+����^\��fdN��*�?L�;���7L�ł�j�H����B��w���4-	X5nS��Y�v�j���Ck�q��?k�����ɽ
E���m=CW+�_p�?���k֦����e�e����au��ٳ8c%�<��
�;�ÊĨ�Ғ�k*��²���<�cis=���t-���zh�`�^����Dfɷ��s7w/���5�.ܳ��+z��¢W�:�T��=6�l�:�ä��%�Ӽ0�2#z]o��*�y��׼nJ�α]��f	�\�Rmu&��>G��g9��Q�ޔ��*��mӗ�.�ti�8�?�8o`7ҧvUԛS���l��1My��VKDD���T<��Zm��y��̹]((�e��Ap�g+g_هbzeɟ���g�Bn�M�z�_R j��fc],5�sF���͜t-i�Ӧ�;޷A]�W�T36�����3
xj}R�)�cĄ���R�6uh��#�z�ƪ�2�H0	�o~�B��V*�`��Ҟ�@���V�U�A��.�P�R�{~��|�I��U�]��S��}�n%{����$�K���JE>�8�%�����������T���GM}.Q�O��zB���3�W�yNr������z�T�w���An%`N��4�<ViQV����wG%8@�RD='�u��Eؑ�E�L����O�۩�f��w7�
ǴN��GT�Z��fξT0�l�|���]����lx}��<ԚH��3-z\�(�]�$-�CWd�bVyu��כ��F��A��_���C7��N{���ǘ��$*�j��evnl��`�#H�݀�iu��������R���>��J�8�T4g<��B��k�@鰝��8ۛh�A)�=��q��n�E��N����t�|��eC��v���x%DX��fZ�[bV�����%���lϭ���}��f��d��Or��c6� �L�N;�:jO ��wFz��k'��Ke�H��b��
���������|8M_����n��z&5���PWu1S��	/��3���B�8f���+����y���\:��Q=�feXQ��u79ݩ"x��H8	!s��l(F�/MT�4�	,o�N=-�z����Q�#-���d�	gYX
�?_~���znS|�J]�M�	l�u��U�����G:�Ŷئ3� �� 2U̡��ݐѻJ�T�I#����'`Ŵ��yY�Ӯ���ٷSk� �7u%Eκ�e4]sFzEL�f�@%���U�l��^W��a"�OZej�[N����l��k�n�F��l'
��G\����@
��c������s:ȝ���,�'�r�.�f�\��Ħ�1���(��F�덈�a,�,��QE:���uve���`l��� &a�a>��1m/�O��~6�u:k�O�����1��rz(��uO��7�&a�pψ�����&���E�b�׈e]��u<��)��g"�{�j&sWU�n�����˯N�_W��q��𡪽��J߮7rH����z��׫p�~��R���at�$��3S�+j|��n��}����Sv.A�9���K�Mr9�K��@m�g�J�Ja�Ԋ8�)����g����4%��¯+��$WI���.�w<3����[�5[�>Ӵ,�e��ێ�Р�!HNs�
*��#�lS2���+����z�IT�^[�3�/Wz��'�?����gz�Eu��n��\3�Zel:T�ιs��ѵ�2���̈�
��g�A��s���ר�<���Y��&L� �y�%^z��8���#ޚ�lW +Ɣ��w��[O%藺��f͟�f����\̪����юL�@h0�M�*y�/_@�^[Q��PH<d�#�=w`���+=��,��c���앸_�g���a� ���%M���۝	%�B�`�SU�Cѽ��+n�7L�Q9U�_���q������߽�OI�^��+���Kf,�����A�^����{���<J�0و���!��D'eEַQ�MX�Xg? ��ו�ʑI{������
.Q�2�K%*�����7�� ���&b� �Z1:��=�g��,4�A�z���ey�;�Qg6�;��	�NӪҤ��A�4r^e*�`@�K�D�Q�È���h׵�6�-�6a3(��8, !���ml:4L!��]?.�xlҪz�X������Y�U��G {�/~ȡ������Ǻdd�6QH5�Z�NP*�(��L�=���v�]ڽ[hN�]����������{����\����^�/j:n�WPc�,�����Aǫ<C:��vnq��K��+�9r���8�.��/z��n����'��g�ݵ7��g��C���j�f���i���ɩ�����O���|]^�lVvh@q0a��IG�������������nL��wo�|.8��T6t�!P�����^����k�pL|a�gl*&g&E\��ׄ����t�C� �d|~ѻ�,����ZR�c�wW��n<�4�cF�鶆^x��h|L+�'w�i��AJ��d+�2���jM��"f�uO4�����T_�qw�|�d���9=�Vnt�ex���z����C�s�>{	�`_ �T�r����u��{i�8���M�q�����u�����oo;����:=��l]eϬ}TL�1�f_W�ާ�0�p"��w��3��y���DJ%�4,b'
�H�'��&k�N�Iz�u$����4���Y+��eu>�D��Q�<t�����ʆ\�P���ғA�M6�.��;�Q���4M�V�������ӣ���5O�x��3�Gdױ�G���՛����R&V���`w]�m�1�G��vJM�Mu�߸�(e S@���8�����'{�>�����z׶F�={��7���6� tI���T�"/3���>���3�{�ˏ��S�S}t;�O��<�O�� �n=�7�X����0�H�O�X��ї9��R��Ѓ���暴*����`�����kI-G�uGڞsܜ&�篳�3�<��TL�M��ڵ�4�z��L
�-�4`E�\��=^���`�i8�����,Y`z;u�3F���⾭õ4+�9N�m�$���s����s�>�W4����3�DV%	�>���27Y�W��｡/@\O@6yͺ���w YQ�^"8�f.��'r�Ӿ��:_�"X���R)8v��y6�e0�K]�ի���]T]��ۛ�]�G�ր"�Ua}�N?o{��xv�SÛ]��޴k�,��Bj�p�^N��E��^Vr���d��=�z�?�hz�uf�(]�T2�oʯܻ1�xS��n�;��^�����`�j�vm+�1�PmBuX��H��魮ꐨ�X����+u��zv����������z���[����J���9B ���=+��f֮Y���6�����c���4�[#�(F�;F���uӨ�g���iY�z�厹/ݕ)v=�����}=W	_r&T錬×G�o��7���ޕ&(����TU�d���ZF���*$���b���>���Z��[��X������D&�m��nPz�<v��ʪ~�0ˏ*<��f�F���sצj:�1��I~T]v���O2(j�Y�g�:�P�흾��^�`k��hLr�;OsP[�a�O�A���K�wW�_xvJ���9�w�r��7��C�f�i�.��e��6n۵q�9��w@)�~w9�GW�vy�ؾs������MW\����#Ղ/&-��kSy��AI�	|J���Y�����π�WS��7.,Y�͔d�B�@P�@l���(��.ذ���1R���=Uuהb�	�!���ϝT�d���Vr`��P���(�+���&��.%ѽ���'�'˼;(�a"9��`�w/�O�܊��9��Oe�r\��I�Pe�[�/v�Q��or�;f{\X��9[�o���C�/���d{G����5�'��7y�0���V���'�V3� o+[%ٚ�F{c�sd|!��@xl7����HɳYӥ�����5f��b�4�{-��vI�WIz-e�>�A�t���O��6z�_�[=�\�>��|�U_l��>	B%72{j?.Wi���"�՞6'��ٞ��b�R����s^w�-1t��w%�W.�`YBG���]E�6�S8r��X�G�`����Y�w�.*Nq�S�B�L�|5���v��	���� �J�i��s�X9�uY۟m�La�l#lC��\Ÿ`��Z(	�y��b+Xf˔	s��i�]zh�AW��hB3�X��c�m��L[uh���8�j2�.��������v�[���yp>;k<��Nҝg�ݣ����]��v��:��nqq��*��{rG��=+8���UM��㶽q�������i�����4 S�6߿�ʄ�G'`����#mX�O��+'��k�Md*&N�������U���A0.%8��O�^�����c����ӍM�6"eA����90ʇ��V<���%�qz3�ݲw�ηU>�4jhy�L=�^��OP��ģPy�7��F��%FV�bn7N��!�%�K'2Mn��e��#���F��9ӆ�?�15��˅�l!i�v�A�"	�f�P�M�> �PE� ��͡0n��\��xǮ�g����璍i��Kx�z��¼Ռ����E�V�krv��ؼQ���J�Qn:��t%�zD����ؙ��`�.�)�]5���Hg�!U������7�Jm���R��5w�n�}}6t�m;���z�.��!ڤG�UU�
�o��( PDЃ�3����>�ݹ/���/won���	k[�1��{R��K�&\���ϿN�!ͯ�-A$�f��̛��蝘^���'o4[y��%A^���Uﵿ$�H��2��WP|�?�O��(z,�z|�Ղ�mv��F3 ᷾\�r3y�������Y��
h�Ap�����}~Y�p��w�Sy7���WZlL�>��GAL��)�H��KJ����l��d8���ʌ��Z�σ�<f7�����	:vb�ŁKG۰{�1N�}mJJ�:�~��Gt�׍�[:u��!y}�7dd��bN�`��N�ʤk]wn^�wf�Bii�K�V�D:���w�>�g'0�k,*�/i��??!��Y�������zٞ���Oh�JT��T�H=�r�g��6���辊-z�����﷟���Ӎ>-fLX3Z;c�ta.v,�ke�A��%�Y-��l���U)�gv��N�"�֏/G^Rii���ȫ(K?_GٰT�_d_4��Jw��h'ӵy���#DD�!و�z�D�Ver� ���j:�_�밚������b%Hy���&��[Fb������s��=s��O^Р����̥�{���+"0U�{:�|z8�Ja �pa�h� �&e;�AH��Veu�X�\����;��:�̵Q)uWfz0l2O@0(����*� ��%2�$�����;�mI�u�w^��S
��/�7���a������;͒32��˩�#A���ta�ݕW9����o�j	zV}�*l�V������ǃ�s8��M��4�.�(�龨W�����"�A����$�R:���ׯ�LI���[��҈���J�ss�/�}�|N����-I>"{rO�k�|��=�q��UO����2gw|��򱌐 ��]B��g[f9SA���ϾO9~�	�
���g-z�љM���|��ݎY"H{�R �X*[���W���`9�v�X�G>z9��& �Q���맺Ҩ9�<r���W�ݾ�F�lB,�Vꟲ�z�����x��PG��nX�>�%N�o�|s���$ν|�X�]�(E[CFL�6
g)�]��]ڨ^J�yN�|�k���w���aGi���'T��g��~{I�T=���0�M:����J�R�s��n�����f�%���p�_>F�[���}�	�`��7���w���~���u�+�,�k����7�7��!M�D�՚�sӼSS�n�j�_ �ܰr����M�C7������ʠ�\��@������R<b���w�MǕ�k�zu�{�X��B!L��TﶽY�'����!�h�6����X�3���tσ�d���bZwm�u|ǐ���>�W��]��u�� A1���%{�[:�ϲ�k_v������ͧ�z��~!���i1�:�#�;�
*���4>�<s1Y�������#�|�p�js��V��^��m.�/_�����=�J����&����O=L����m���@
B�6D���8�)�~+��|���%ń����
�ņC�0�qB���I�B\����6���3R$�����8��˙�)�g�k=�N��!�������z���������J����N*n�ʟ��Ů7{�w�.�\4z�o?ni�5���s!_�b/�v&E��?Ng�;��l	@9st��J��b�M��	�R��=�3j�>��aN;��^��j�D
5�D�}릨ܬ�E�7D��u�~���\��A�@TGy��7X��/���n�[�*n�cA�[¸���$3s�5(��:�oOj��S�^����!�?�!��d����k�e+���xv""������zqS�+'�fS�$�Og�������zRg��{#���\�}FLUn���d��ZF���8�w��[����UA�I��[҅���F�y�7�y��ƪ��н���-�w����ϭr������ə��a�(S�{ٛ{)��^������ùy�л�^J����d��eV1�f3�:��:=g~�E�B�35Ѳ��j���߯�&��F�)�9����mVը�J�k��U,�3.��j|c�|�5�������i�C��PZe���ϦL��ޝ��=�|2�:�n9^i��`����3||�N-����d{�;�v-��`֦@�аsJ20��wk_��K�{����>��js�;�婚���Q� �؟����+f����-��I�>�1�[���ʙ~���h0`�C���\[>/�\]XœL�[u7�w�5�c�z���X;�2�6{Z(K�ذ�3ڦA�4�F<	>��z��m�c�25�<��7� ��Q�k���^�z�M���=�T�D���P��t���a��z�nprl�f�*�j���8��H^g�AGmX���[��"â�`=�;��t���z�;.�̄���Z�3!	��u�E��SU^�R�2��̳>G�ݻq�x��մ��ov�Rش�T���n��t�侕�rͱ��0Nt�����g�/��=X[�����4�\<������_��8Rn^sψ���7���ńF%}���˸�|tG����n(ݸ���[@�w���ٍk��Ɔ���Y5ϯK
���j[�����Y\�ؙ�砤�+�e�+U봀����b�:����Y�̔!I�M����R7R� �7��и��	z7L�� ��8����y!��ًD��z�܎x����·$a��iu�_��/��?e~��pP�$���3iC������� ��Yk�߹uu��_��D��ڙE�(��8"Vg�Y����s;����3�G�K=+�t?$ڗ)
�J�5b��.��w�y�	kC5dP��f�)��=�"r�C�ݶ�?5��93�v����|��S栖E���Yy�S�mA��IW��YH��Ew6U96��$��k{GB��ga)���}lE��ƨ$�����̔�!�E{�{@�Rx̹Q���mH���r=C��Uk6M����Ts�^�k��8GV�-=WuY�P�����Ja�QF]ɽ|��%;8g1oga�Ҿ��S����y��q��r����62��U1F���ދ�ƹ�P���+-X�(i����\��;{g��TOF�h�d���D��)�W(���Ε��ݚ��A̬��r��mT�I|��֫�-��O�Xt�-S�z���<�z��Oo�h����ݚo��0<�C��/���g��m�h���E�	}Y&���[�޾�|�u����>lB�Q�w>;$/a�܋$+�f� /�ո��ZJ0%�L�/������|_RU;�Ve�(�.W^��r!r@�36gP�V��H0(s��j�V�vb�V��*��;�T�.��������1C��'�ңw	��˩	Gз+�Df��!�𗵳��z�i��/�7\,U�s�]�ֿ0����@�i���[�47�M5�C�髣��֎�;J�$�����S�A��j3ܔQ�p�)�-��)���U����f�5�]\�y�'��|��+l�'k�YEI�0뼵(��@=��T��U���~�3�R�i��Y�m�gSY���&�+)���l���0��x� S��V���m[�-�Ws����zc����(�<Ίasr���MbM6�<8�>���(k?+�*��O/�&����4S�x�u�ǹ����=Ө������,���C��9�f���uOH�Ɋ�L�i��$��/����B��Lǻ�T[7Q�_��Z=.���,�X5U�2k��w���6�-&'\�s:�30j2���ED&C.���ё�>y�`�V%�FBz��`ªu���37;6�Rs�h�V.���*�r˲F�e��q��0�abq�g.�|)h0�6��n�h,Dq3n���鴁x���t���Z�;f<���h+�.���67���Х�ܳ�U����͝��\V
4�� �ѱ�y�����v��'TOQ9b�+C��;�O�ͨ6{�b�ܣg+��I:�����94����Gݰͨ�	����Dx](eX�jW$��ىoc�L�`N+�:�*u�fm	�;��nG��l�q=���;���*�����C����m+���z[o�V�+8Юi��=���\m+I��UUUWJKUm@J�J����&����*��-Q���HJ�FY�h͹ĳZ�He��	�$�Y��:�۩�@z޳P9�����7�m#t�XRP�J*�v��K�����\Ŷ�tl�i�c�5]x+�-0���x�l�`�[1��8K�8f��B+�^��ٳR�f�4p%fq����'�5�9�n�v���������c��Q���gp�Pl��u�k��b��ΓE�.�UԶ�R�r	��d��8^�bh/]d�8��5��a1 �5��r�R��lH�{=q�a終99�a[s�(M��q�4��c�F�:�����;G�Q���u�s�v#�D�ټ����gu��O0�Q�۩�Z�i�X:�tt�N6K��t��e1T��[IfZ�DS:�[Q-pv��Qg^1]��f�� Rê�NҐ(݆��Q�lWZ�Ȝ9�ݪ��C>��E8��ݰ�l�{E��pu��;�˫�8�-6�C�=�B�����*��v�pşg6l�6"��k^#vTl�hd�����m�f*	lѳq�V˂E�].��E�-�.l��܈��Mn�J�m�Kf�V9r�Oc�k�2��\(�۷a9�x�=T��sJnW�V�M�����wUp�Fd�|U��N�!l)㱵��p`�\��t4�f�5�[�R]��7�/,RAp��]BU�����X�M<=���ڱ{�W.�bkh5���%��Y��sv[�rH�u\��z�5m�:H1My���Ŵr5LJ��mX�Ҍћ���u��4��(+������$2��a�ljX��G�� �C&�h��$�'d�zl;�Gn�V�]fWiE�S,�݌�
�"�=��q��-t�ۡk���5Z����'&�pO��	vrwg��L1sٶ6�շYHLAճ����	޳���㓊J�Bz�=$K�7{k\�>�zh3�ұf�c�����ô�6����]ezQ��C�m�L��I��5��տ���_�W�����^O��w�{(X���B��l �ꕇٯ�0�276��>�ye�����e�q�+4M���!���@�8,�npe	:�S�ڰ�+]`�P�.�gU�{](ٻ��@�y���I���4���uw��dS�97����z������y*^_R*:8��:ݬ>���퀗6\IA�%��Ȼ��cKrK�{�+#�����_U�;��Z�O�`s���r��o{S�Xo'\Okמ���t�
��+޵|��|uzDD� (�� �>p��_�\���׌sϝ@���=m�#��ʚR�݆U�B^��eO���\��0�i^u�g<��U,'��މ��֠��w��=���e(����,3�����vuc�؇E�nF�lR��\q���fײ1�ɖ4A]�o�c�@��Z8{%lOz�n�e���IF��P�f}2����Jh�	���ދ��+"�<�|�aiד̭�;�Jb���ק�[=�}{
O����O���ߣ-!]X������h�9�~b�38t{���g��q�����c� �%��m�W��F9+0u.t���
��E5r����O�<��^A� Çp��\�E��/�
�3q",�5�v��Wmq��<�%��;ݻƨ��Y�j�ͫh���.��ۺ��K�1�S���������@{�Y�X�*Ig�Q�"FI�����'s�}��:uiT�y+6V���(<�w�&�D�hg:��]*xfW������OCp>c�η��"[��ˬ���n��*�|� m�R�{��h#��"B��T��}��ө��~�$�I��*�^Pd��g}~�z���Y'}�\�ʺ����T"�A@qޣ�\����N��ފͯf���ۜ���<+���v�;�%t�V�h>'�;�O�C��H�<W<P��*�;�`��Xg8)����uQ�_nyߢތCJ�1�[�Hgz*ٿ>�'����fꉫđ�V�tۗ��]��DD���B=^�Fx���[�ݨ�?ZHO�=�&߻�0������ñ?R�(��Wi�u�q<N�)�(�ـ��]�,-�b�h��s{6�6���p>$0��]�� ^�dw�WI3h���\DGR��+=���|s��w�9����q���C�Z��r�,dwAlCp�(m5���o7��|j�{7�C�ܡf`N�m��K�\~���M��&�m9�"3����;��R��u���]jҹ4t�т3Ն5��������̜"�x��ո[1��)�dÕ�zH yhIq�I���Qb�N���P��{��9И	AA����~���������P���뫯��nM{�����3:f�����
�rt>���� J��zڂ�܏R��C���$?�6����N���PUA"Zf��K{�,��d�Q%���W`y���]��rL �3j��Y���B^�����t�Q��Cg����][e����)`7.�*j}\��;:�X��oE�� >���q�9W�z:�������=���:Y�/�����GȾ��=�7�1/�U^ԯn�w{����HQ$\P��)�o,.��;��l{_x���s�Vk��&/Ф ��9�`�.�6+���o������w��m.E2GL�F���҆�'��^3}�H�F����)n}�l�c�<�Y���V{�w��p�zן�Z�hwu�:��1Wb��X�g�A{�`�ය���;1&ch�ֳ<��.w�ӊ���D�QP�'�Q9�:|<<+T�\�9��-�x���Xy��y|d6�P ��0�:��Q����%�^7k�[��1���*�y��=�߿u�Xd�9>�#��0$��M���U#��wJ����\�6��tĈ�����ϥ�/޻b�.��U����<  @�Y�O�Њ4���3iN��7��/u���5��r�r�5M|���%K�錬��{��Y������l�|}bj<M�������Uf����lC�6@�]?C�n%n���|�9KD*%m�L��M%�+}w������� n3ګ}r^��YL� zy���&���<<���!�]��k
�^wA2%+!	Z�����E2��!:�<�w ¼(�����_���>D�v+���`6z�oh_�t�mۍ�xw�����*٪�Is���4���Ū��u5
QPI�Ԋ���n��3=|�Y�=��*�M���,�[�����^�)���� ����4f
X  �D�i�:��N��g��[�ŮS����̷!t�Rj��f�
�Gn���ak�ۅ�7��]�5�p���[��������,<id�����i�����v��snv��d�{�!�`:�cv�0]qյ�룉j�x�X�-��F�2�61��D�>0a�9���S������{ж���g�7��/P@��LbJ�mweX{�Ĕ95	І�m�6���Y+�
���vov2|�r8 '�� ����5�&7�8I�J���:��bì��Y�G(�z��x�n+��uy;]�f�:Aj��,�����I2C��N%��� ��(�YY�g�� ���E/�<�l��
$�% ���2���!4m�^tmlAiU�=��!����_]����8���;3M�r΂�;U��{9rQ��uge� Q�d���U.��o���6�6h���!��/��Unt !��E%s�����|`o7{��4N�����¿a����#�]^��Ge���Au��=#�Fh�v���$ �W��l�DN$�o,��:kx���ո|D9^o�\�]�T�-Pe\��V���mX�T\z�&aW�κ;A�.�`��FKu�s`��]�V�q�	7� r���N�ho=���\��S��4K���՛�� �`y~�3����d�aVErvj:u]�X����M�/��Ԛ�I�r}�ϻm�e��Bp~6��%]ix�<��Ё�FQw����|Hc�=ǖ��yY�|�8hU�LkAn=����c;����;�ӽ*ź�Wx���9	��h-�6�cS�6:	\z�ŢI,�ʝP]m� �q�� �)R�fd��uG��=�Xb��2��\��M/J���_GҔ�[�~�_���4�s!I�S[*015��R��Hħ̣�V�W�%�Â�d��b�k�vDU��˺�\��ۃ]�0��%�]�(mA �a�xG��[Lp�/g�KKB�BB~�7��*\�|�M1~�u���w�������X·[:�ׯ�3�5�i��l ઎���*lzr7&�s2�Z�7K���r� %��VP�q�]�s�4=�1K[^�=�7�xґ/&(J�뇣)Sڷ�+��6,p��t�T��M��m4�u�Kog�hk�٭�X������}�p�
�2��v\��=�v�Ɛ��o��9W:펊�<�f�|*��Z����a_�.^㘥<f�&d
��U0N�	��Q8CQ6�fj����ʫ����KW�~�JE���c���*
^��o�,� I����:]�-���#�<�J< 
�~��wh�\�\ �r�,�=��:%5���� �{�U�=&�}�
�g{'�-�1q(��)���H�"H���ר��Nȯ���}~�Ӯ3���S��jo�*��À�P�6�$�����o�R���k���k�E���ѓ��6J\|���7}���������'������Ư]�z�q�'�Q�(�P�7�s�f��\|�h�0\����%;|�����2D�G3�· 	̠otTb�GU$���nR�傖�ذ�z�2���痥�W<787�a{��^=�F�5x&�׹�gU��r���w2��>L(�Rc���-�-�~0.��$߈3���N4 �9�q���>2-��ccޙ�#{�3��od�P�Z�9�1���'���L��K͹�}�=���m��֣a��	>$���E����L�$��Y�ԡ�Ww&�K��k��T�V=��Y�����!�`��wt/ܲ�)�_Q�nfd����<7\n�wU������f�U��Z���l@��4=��v�U]g���ayhH�œ�٫j���v[��٥�F��.{�]�h��s�e��<i��o���X�t�c	�޵���{C���Q��jpU�)ش���(��S鼕�,7Ѫv��c���S�T䜍����+��-{�X�nF���qݮw�)I'F}BP�E]+}��D��G"n�V,�aA�V��X��m��-f��Q+98{��gH0��X5VAF�\M�L&\�I�؄n��j�tj������Ic��q�<|w3g�*���wj�&!�c:S�]Q�����wc}��<bL�n<��=O�2�e���f�a�7=>���RI�E�pJн�;�m
�3{�3_��d6@�b��J��^��8�*��cs����ǘ��Cs}߫���}
��91�f)J��s�,��G{w�J[�<���P��jWb�օ�r���Y��:��M�G�dX3W��崺�Z������i�l_Vm-8�)tI�e�1��IԾ��9��> ���]:���h{�֡	gG��U&����Y}پ�|�(/�-n��8v��!#��m�V����Uۦ��^�h`xI������f�rdJa�r�_)�WnsD��i+�{}����>�'�覱�]�(4��fͪ0���s�{���k=��smJAQJ3{n���O �4�I�L!=�zf֎���rߞ�g����Ɂ��L�%2{�juo��;���e�zBWIN�Y�6;�c�e�1TZ]��^`�������F�!��0�	���Ŕ87��u�e�~�����`��ê�����;��j�յ�q�����\	t�Z7�K5��,�dL%)	������x1^Q ƞf�Lns�f��W�ĨAy�W.�W��Y04f��V�����檮W�#yC�����|b��3�o"�b�-V��|J�������d�λ���x`�L��p�+�c<�t^B\�l�r�Nx�ɮ7^�kac:.�a���&k�gڼ"�R'OU�me7kͼ�ܾ�L�&zT���,�ˮ�ϱ��;k�r������k1�{}ĵ	}%W��q�P�M��ߙݲ����Y�:��G�i4�mz�i���+��W:�s�W���>&1ٙ���τ�/Kڹ	��=�Wn�<'vZ�C?�^f��(~]�U�����a���"�6͌�D���@�J���RC�!�:f���k}\����Uj��k�4�vˣ�d�۰�m��cMn�̇pS7j�GG�󋌲.�s(���q�qF�ׅSul�*M�պQ���T�h�z�7[t��u:�5���r9=lb��Z��5fB�0�:Ҭ��c�@�	�P��P�=�!�뷵��\����C5����l���#f��B��X��"�L8+v;.�.���:��v�؀�"8��v���W^�?4F4;vQ]>��+�R	\���O�4�#�|�pCju���M59U>W/_��I�u�����Ţ�w���a�Xhw�?*�t�ϷrqE�^�w�|�o�Ҿ�Z��w-���Y��@a�a7��Ͱ�m��.s�et3����{�Ogܞ�x�%ô��k�k�)rvC�j�k��j���l��l�A$�~֖no��p71��$8(��;�ƒ���{�[FllWN���M{�Y{��g���3G^-��m�S�qy��
r�aڝ����s��qp���������>p�|�3��w��m�F^{���:=\�F�Ѧ� ���/Ⱥ��G�]�Ǔ�U���*��wo�;.뱮{7��)-�Uv���}�B�����~��lZq):��1��7�f�unO�9ύX5R�O������C��[�8�`/���/R7|$i�ƺV�{M�9�lM]?#�o<�f �W�G�X&�y-�[��n4�Q�L�X�`�=t�c�f�u�>{<u���pi�����h8iAAY���p��� ���fl�6:����X$'�W�^�us6Lē|�:��Rz�>����O�g�/��|l>�7��m���K���G�	;�B�{��܄f���'�ztlN��Jn�Z��`'�o)���E���#5�u;{�EXk�U	OE=5Ѱ�j��/n���$\B`1Q��;|z��WM���e[^{'!Z�g�A����zl�k�/HJ��d0�2�S4�'c2B��8Tl�����S]���%|����=�z�}99~X��ML7�����i�K$ɉ��xI�m{��Q�#��e^�Vs�;��;2�{�Y���J��6��HB��ذ��4ֿo��{}G�>�v+ۊ9�:Gs���ѯ'��s�����/�a��V�rs�-�~�@/�Z�ϴ�n�V���P��.M��tǷQ���S�Y�ce�}�`��vVʀ��:�����3���\Y�;v-]*�=_n�V��[2�3�n�?B#��1�o\��NO6#DL�Z����RN	�-�z�b�v��r�l�a���6���]"�ev���ьf������P��=D��|<m�<��y���O���yO�����Q�U۽�[N�YfM�f�=8��D�������<4�_!ޔ��s�HR�㬈yyL�0������^wC(y8��T:�^����^Cw�G{�*�{�r�����2|���[��wܺcqpbc�=�{�y�zYl����r]�ܰ���m��+rj{v�I b��0��MGC5��{�ޱ=>��A�z*��^J���͙��z��*<�eO@�_{w_}�%�jEJ7��U9��U[wy��Ksgl��i�Ӌ8���\�hVc���x�Y=�d�X���5�_\�C�V���~�wsGs}���D�b���)�������rZ����L�X��MՓ�z�ټ�G�_%��!���K<� Q����_��dp���X�8p�o��O��%w�2�`$�x���s-<zs}�v�'�<p)��g���/t9/Z��c�Q����	�:k�ˀ�	9%��������w�Bh�1Ռo��*s;����$�0����61w&T��oUp*냊5X��Q���g�2Ֆ� ��"s͙g3�M\j�[�N�55�B|����@�.}w}q{�9��i��S"dQў�=D�&�[�$�V����������0��Q��8�t\��]B�~��Ɛ�[�FDO�U���;3�͙�:�}���w}2�\W�̷��*ȹ����%8e��lS|��.DO��ܬ��}��T �5����g����W:ɮ��a	�''v:!:ognt\S[{B����ZjqX	�{�Umr�44�U��]����"��:���We����\���=��蔹-Dw�W�k��'Lp�J��Ɠs���Ռ=�O��( �(�c��q�?W��=�^������ݽ�bY �������6�9��R��٥�R _"�5�f��k��&�2Kl�Rp��\s_^[�r��Y[�uM���S�^Cl"J<�A�����dY�����Wtՠ�w\�4v�z��v�/#!��Ҋ���Ӥ��h��)[Z��͗VI�5��D��}�C��{�.�윝13-J.��k�S�"5��nD�(NgށL�#cd~p	,�-�9YҦ�q2�IK�]Md�υ'y�c����k�S{h���u�vj�����bhy��k��h��(�.R��\+�9۸�ʇt�,��M5}!��F�YY$7%�1�}����KV0ܳ�@���S���m!l��;���K�*-ox����p��Q��*GI��J��n���L�z�C���f��>�EEjY��k�X�4������
"�'Q�9۠���������.�]5D�쭝��=O��ef��X8F��0VvS.r����mu�oj״
��N1�T�zӳ-r�*�Gso)�]����d��w��t��޺T��u)�B���RwQ?���Ĳ]e��ݧ��K�K����8!]��Yzm���V�ح�yp
k�]�L�\�4zgb�wAa
�w�kQǷC�v�G=�����b���u��nc�Od��I�p�v�JжT��u�1�K:�*����l�=Z-+T$�bה���2��]��/fu�C���-��r+`�֌��Γ0L+�9ٻ])}����jZ+�u'0��Syەͱ�g5��U�v�3��ݓJ��U��#+��=5-B���n�"��3�x�I��'��e��>��i⁲+��x7|�R�y���b���+l�t�LT����h���B�S�꺹Y��r��m�AM�I���K:�+�ʪ@��<����r��k���x3�4sf�	��E#���jX�g �i���WvϰP�NJ���N]u����EBAn�/�K#p+[�_	s#XlנO9�ʶ���tBv��i���)���n�!�:_���w2��4����jT'�[3N]x��7��D��]��=��H����pR����4|����Α��~9u��T}�����B��ً�jm�&f�ıX�k�"��Iq!�+��D�(���~���Â�9�q�3�V�/i`��j�%9�G󯟷S�j�|8��f�Ǻz.�wt��킣�p�$2�W�s��){����Da�p�n���eю��T� �|��Vj�����0󎊐�����}�h�J;��nWS=��U��-���P��@�U�N��0�|~oe�P����	ʷ�c���]w�����Z���ӕ�bYd<��>���7^���{h��Ϻ�|�����T���A�㒞Y�n�~��+� ����x�Ju���E��	�s�t�����Gwz��-=�|g0�dz2�4��R��6hV4@�)X{tu���3An�}9�B��wV-��_U�Ӓj 7C��ut���i%��h��5<����۬=�rt[5=�f\d�O�y8N���X�tRC&� �@�Z^bЌB��Ґ��۪���v���z�6"L�0�	MWd(��
��L6;���4��^C
�b�:��Į�����qs�F69�Eh�8�l�ƳcGl�4�Ԙ	��&v)	���Ѹ�X�w�l��N�E���^�;(���
�^-{Ԗl�_�\�
�^w�����`O8 �{$_]�[�t&�P`����U��b��==�AP%}��*h���z�8�U���p�e��ȇ�[��y��B>Q�c�gՔ>�/�����5�qի5�&��j���Y���ن���FT��3��&�r��g�"gB�X����+͎�$0��@iº���P#7��!a�qU�$��;s�kF޼~�����-�>��4�ou�sE��h��Ѽ��,=�į!�gf�ѳ^H+s8�6-ҿm�Lӽ�F�)2�)���P*tӟ���|���_�a`w�m�fϊ��v�b@�<!���1~����)�|kr���(��1ۙu�=���21bپ��ز4G)���2~�ƨO�������v0�=<�ĸ�z�߇ga��/I���W��G�����-�e��p��4ݛ�-kԐM������ш�F'
N������j��͓y�2-�	�����GTu�''^�na���af@�uVhyol�\I0`:��e�!�k���1�Bp���6��D�휐��}��Mt{�2���n�b�y���}��hwŹ��긆{r�]�Ւr1˯b�J��{��o'��G�O%��=E{[�y�E����M���*�0l��
�j����a���������Æ�%*bفO@�(ǌ����xz�Փ$�[͟t�iA��)l4�0�juɐ�5]Ǝ^z��;n'E�|��۝�[�C��7l�#�8�#��mI�����a�3m��`RH��P�"����׺�:8�909�Vi���j���,'��:�����|�GU�@N�$���]����ci���y����<ov�����ޞ�~�!l���&�c#˩�n|:������=vϡ-�&���q�2T��a���z	CP�$2��W���᷵M�흶0�:�~ȑ��>�;�?����p�VD��h߹�~�qs�(xd֯��ݮ�N��w�Q�F4<����8����1q�!��A6���ݞPM���o��՝�G0��_t\�.g�;�o��T ��"�	�5Ш��B�^��q�}�/�_����j\�(��l��tA�����p�E����0�\'����V%�R�w���#�.g���@��Lߍ�{@_a�_�|�rO��
~�V���qЯ_���=�<�1�1��Y�!Z�{��ꕓ0��Ȝ�ж��&?���B+$�&E퓑�u�Ml֬���.�L̫�!���i��+��+܈i-iY�N7���Z������| FX��&3��mι�{�7�N�Y��D��a��yզ�.���M���|;
�)k�ӳ���f�xQ�M���o9�徹2�d�k��`��k��G/X8"�$#i��#R�����7��/O��4�:+ܽ��X���Ҕo͚W~�/�V���/kE5��o�H6�;ݲ����\�{�%׳9P��ق�.���M=3ӻ��b�/���Z����:��lf�ު�*�ma��R�*�Nך���5�/��ta�nz�ѝ�^L��v���*&��^�6Cv��������Hz"��%	5ėL�ўwW@�;4T���Yk���;�_���}��8JW�3�H�v꟱��(j"p�"e�}�������������|�ޞC�Dg�ƣ���tym�VW&�(Gk�s{�`p�I�ۙ��$���7uK�Ƀw�.&J�n�Y�����������,�-�o{�C�[;������Vj�|��gu��`������Ä[B�.����uI�u޻����g�O?so���|��������늳����Ʈq=�=5����i�h��p�XE���H���_3ӌ.�I�WaPf�j;W�v�Il�މ�Eh��W��s�T
����_��64��M0�,���z�%ؗ��Ռ�{TX�lמz�JV�1��~���X����E]�VU�H�����Z�Z���=���^�AZ�޻���'x�)l0$͈G�G�ȓb	�wUY��]�����t�4�����JxL	&J6�\	��L���D],���!IT\�o���+7�N�CH�wt���������3mw,2�@򕢹�e�?շd�ۅ��|�u��e��<U�|l#�n������E�`+���2y����N��*2{�T{vV���Ti�����Q��3���$痂��h��K���wuv��1}]�퉓q�0���E�`�Gf<�s�A(X�a�Rw����k����"Qs��v ��c�ַ0|X�ߩT���PȖ������6}�yVh�E��A�|v^�^׾����k��.�v�á�!A{��P%9�3]��Q�Cz:ޙc@YN9	p��nFHA-`��{y̓ޓĻJ����c�z$��#�����t��-^��<���B++0���;�;�<ZA�p��O*J���;)b�_��2kGfC_9����R�^��q��5�*�#���N̖g,~���ԟ���L	�����R�/^k����Ɂ�r����x�6��؀�iuYT��}�;�r�ݸ�B
aa6\��rM_���٥jy��e?��P�>(;���$�7��4��	�[.6_�S�4�rMf��eM �eze;�w�RZ�y��
�D:/��fvvC�����5�w�Ԯ%3~ʆ�>��kPS�vR�C�f�s�r7��:)�6u� ��v�E��k s(ރx�����p1+��z��+�4p��3j�R�H����s��q�`�i���^�5���	].���4H#�饵�X�=9�\ohK'���l����n����H�N�
�t�X)XT�miS\/M����q+3L^�1n��X��0
P��t�l�M���"q� �ǔ�6;u��l��:h�C���u�^�؅�[HKR�Q�����
��A��Z��Vm�{0a���a��/���I�9'ݏ�jx��<%Mu@�����҆�$�d�)5����|�S�r[y�tsk�\�/�?3�6�{���T�|�<�C�'����٫�Z4�_d2�8A�=2S�9Q$D��-ᛷ[��~�~����7��v���?��\}ߕ��j�^l?;�9��@�?R
,�yĂ���D�;E&}�"�&���W�//[��p�t�z\�G���~�� �x�0�&գ��>vT�6R��ݳ�S�ܕF]����}��v������1 �Ѕ����B��g�{��K��+����I��B������#�C-<�.fs��;d��d��\s)�t�N�K������+�d��Me�1�N�D��jy�a����z�w�e,6���Qs��j��tf�/x��v)W�}�z�3��4�ԭ�Ž�*�q�c;���4�6�#�Ϧ�M����d�.�ߋz��N%h���!��C�h^�+��z.q�9����䷑!�����צ|3�G:�Ē�r ��Vv���HÄJa�,UɃ:m{/{�ù{���O�&��=Y�0z�}��>��/	$P�Qg����b����6��l�L�%3�W�'ח�.�po��3������n��A�)����ɼV�S)>�͚�+�wnǙ���^��pe����{�(����|�����v�X��Jx���`���m8P�H���o�W2�T;z�s���3@���\s2�cE!�e���GkTu��N�`!9�F�(J�gj��n��σ�}�T�-ٞR<:}��:��Zkݝ�`�9���Q�Ӻ�a�
$�Z�ԟ?>��֙-�i�*��"��^�˞7���ξ�H���<U����tϦD�M1S�i`���Xw;En��,ì2�wnj��+�%8%0BLuPo��}�×oJ��2B�O��ە�M���>�N�u�&b�jȊ��c%�J/�[�<�VVs����_-�w��z�~�����1ȘЙm��w���CH��>�cD�*ۖ���^���O?t�iȑ�H֦x܏	;�+�+`�[9��Țx���վ�]=��V��m�L�z����V>�#)�o��t�����궖�+��J�B`gn��ř�O=���lO����R��Ϩ�����o�F��{$�q�s�v���^(�	�e�rѶ��>��[����a�P8Wg8/ce�m�`0�a�P�����l"���r��5v+J�h��:\���{}�i���L��b����b4[1��/r��#��aK�:_���w��0d�4��&�9{qJZ5�������l*�����V�Q�؛�7?!
�d�2�=����|��ⶺ�B��!����6kN�	�fd��{�7@>ʔ���S��UwB�a�?K��W�N0׎�\��!lh?o˶zUż�w|@~�m�o����΢:���>}��{�� �M�*|txk'�7u��`mƼO7O[_
6�Ωu��t󘇑�O��{�*B�Sn�Qp[��2w��<W<]�Mts����)�����v�u��i�����O����f��h�1c��W�G�'{ۯ��C�W|�=�/�����;�qY�{���{�X��go'���۲�"�v�M���}���|6̑Dak��(��8C��M�咕����:W�KøL�Z���eXT6;�Pq��G�Ot��/:η���r�g�M�$6(T���xyu��ϣ��|�b�O�ܝx��1�P�H�3/����i2}ʍ_4!���ln�P˅��lK`�5����Qq��nF��d-���9�U}M�<�=�*���L��[�}Ċ���w�Gh����w��W7�y�R����nD7�4jp i�0j̞�K�ZP�}R8{��8ڮ�ú��b���]�Bǯ�u	�Ǌ���r��a��ĽV_�+�4�|;b�(�,�E2�FB�*��wO��^+�`�I�g1$/2����tp�*� 2���n����h�/�Y&�i���(Ԕ���{�.N�$���{� ;�u���z�#�����J�p����z��}C�;��"���[��6�r����#���2�M����H����驦�j�w��y���@�z�6A�۱;v;��=碳�䒆7"c�|cEx�l���0U�j\L�U�3;�����f���;WD�X��v]��>�p�������1��z%�OQ�\�=`��H�2dF��vĚ?q�I/"�кw�V��s;�g����w�d��ʋ��WA�p	�X�I�����6ɞ}�����N�ٞ���yL�s�A���q����)����6z�]��\m����4�����V\��P��\�y"�ȵ�ɪ�r={>�ԠQ3�㟶d��6[ֺ��V�����2:�u=>����	6Ye��j��hG3h�<��̽>�u�k�8��.��Rl��]�����6i �_���[�u$ч�wT��=�ڂM8p�hC!�.8�~~̼b_Ih!t��|HLf�P`�{]>�ݻ�=Ұu�Bž�W����*��&�B=9�d�mO=ا��%��!�ٕ�FΥ>��2� �3X�%��z�ɏ���>}�I��ug?U�ٝv�C�f�L
��C���YK����Y�Rc�x�e�)]<��t��Z�Z�hl����U��9��.�z�uh��JҴQu�Gk4���;p�Q��dv��[��l�^��#b�3qk�t�*�Z�4n3��V��g�D��O5:�6�ٗ!�&�Q��b����hް��Ok<$���fȘ�Hg�v���jh�R"8�h �chXͭrXbld��.
��5���	a�#�8jҪ�k�'`T�鳢�D%e�5�hr��ַ@��3�Eչݡg�e�Ix[~���5yD���[}6k����2�sWT�^�b�{���l��;4�$6K@��h���Egl��K2;/�Q���t�zѻ�L�,+��`j���:^ׇ������~7��=3���J^^��؏o���n��xП%�ӻ���Ʀ�O�a�hN^_��Fо��t[�lq�YC&w����~����'�aW��s���[��s�n:S��kH"��� 0��>))�]����C�Т�'���Fx�v'��:�A*��Y�Ƌ��'\p;N��54;ݑ$��i
A��Fc��J�K�C���u�~2-��t����^$C=�ށ�)/dH�� ף�k�g)�_a�\����"�yl��}E��Fj��I��!���yT�Y�~�U�����%iC�##yz�y�d�uR�W���f���n��Z���{J����M*w=��s}U<vu[S��t��#�ۇ��zèG�{[�1¸f%Z��]�Q���X��ݵSg�w9�;�)�3��|=<{L]��]� ,*}ϕ6�B�!�OP��I	��!���}/��݋�ڣ=�(�C;�l�d��tN�#��quU��4��Ocю�6�f8�������~�l��+��+�����#���jRlVy)"�&�Y�����vE[ X���ꗯ-����q��ӹf���쭃a��� ��Sl7�p�SJ�t��ί�VX�%Tyָh}:�]Zv�YdXT1GW�{�o2����z;.����rѹ�h�GN�ǠW�-��k3��]��e������k�\�l�[D%�k�R ����xЭ��K���k+`�_h���Z���������,��SgX�&�:��.q� �n,��:?�r���#�+f+�G��\�'�ISd(&c������ՉQ޾կVb�S��k����M
St�V���mP�]��[��Q#��U�־-жn��?�uR
C�y���黼35r�v��X<��2����cT�ɫg�tu��V�o�
e����c�!��2�M�Bf����K�7��Bvڥ�f=�|l+F�3�X��-cz�LIe(޼��mfT�š��BGgn��뤎	^���t�u}9�2��@VU�3��iM���AҔ�D{��X�@ѥ?j��i<%��ԭtMe����x����{�W �2' m$Լᒞ1j�v�o�Ňw.�[/s�k.���HN�/�0���f�y�`9��%3�Jz�^wp���^r/L���s��Ἥ�mp��&
�\�7��w��%o16WqK+��7�8�ԅ˭��w��7,�eU�6�)�˝��4���7?��>v��ԁk���jZ�V��8)�&�RA�46�P*��)Ve���6b�VŃwZ
M>^OWn�˅'K��p��B����]+7/�̗���۩v3��'9��v��[��,�Ѩ1R�ٶ�ee��vn�"�:kYl�z�7n��-E�m��mr]���e�0s릩-Ù��w=)OSv�gEQ�ǵ���&t�0C-ZT����t�h��� ]��'�����jo���.��ؗ;B��R�r��6�m5�x�ڂ����՘�yɜ���QΖR�8�ԣ5&�6hJ�T�N�[Y�uZ�7A�@�s՚"��ZD%�4�i-f*�BP�f�+�٘�����Fs�ۢ�uÓ�E��Ɖ��6�9���p��UC�z�]����%d#v[z������+���)z�Jܔuǣ<�˴ݵ��]�t\w,���,�"�H{![�
U�л,Ňv�&��	�0.��uI�Ɓ	�l:�se�٩�ɐAm�ȑ���N̤���M(�q��jM4�s����m��j���heEv��c�\�Y<�a6�$>�D<����8���ֱ�R`��/a�:nu�;0e�3ru�ܖ�v�����Bsb�v�'���e�հ��턲�����`����1���,�N{,wV���NSs��C4�1�f�6�sa�) kK!.�Z�pv��玞W��*���H��j$��q-ՙ%���S@���#D�0\&�kSFե��SP��i�&�U�'-�0r������Yn�k��+�Vx���ˣ�����X�ec��:��ѱ�.L�* �U����mrމ,4
�����Ҏ����6k��n��ۧ;>��]i=�Wj⺫��:U������t�IY\�Yc�j�ɸ���U�&����3���]�����)�lO��Æ��㛑�]M4CGF�9ԤZ�<�z�.�)�3u�u�� �n֙�C�4�N@���_cahH��P�h�M+�-�1�)�����c^���n�f�sيlJJ�Vi�m�2MI�y�N�׫�x�>��Sʗ�Q��9K-��Mx@C���h{p��/�(�B�(䌬�.�q���]Řp�L��l,��0`�M7j�/]J$�	�4#3pF��;3k�餎^�UQ<68�����~'�yҟU�>�='����L3�.�����ѻ�1�А����u:O|A�w�S}��g�r�|�7�u��S3���lw[���	��+�3�t[��yQwS5�D��b����U�R��w��z4�t&-�%�#��UP/v�\��]ȸ��b ��0+(�&9	�å����}�u����Y#q�]��ߢ/����*ه�_t��®�f��.R��ne��l���a�	�0��P3��xna��v��x���70W<��߷i�۞Q��Vw���㞦srh��S�Q�D]5�_�=cIҐ�ZA��Oj�H�н\e驸4c���M�.�d�n�W�^��8�����_M�1�|*l�CG*8f����K�^.��/I��u[�&���2�@&D���\p>8���ggK��~G��]�����N��	��J��ش��ls����5��<�v;Qr?�}�ͯ&�
,6N���.�rc��^sr==��O��t���n`ë6plG�m���y�#�)�=��;�O��rءgU��?����=�}�G'��*��7��a�� �ݻ��ӓ�u�,��#A�%���J�g�o?\^q;�0hG,#A���;�G��p��hP��q�u�yz}�_8O	���u=>��+X�.��x�2���P�>�{r9�G��>�<� ��SsS��7�%��H��3�3hq���?�v�Y��x�i�$Cݾ����*4���x=3U��u��m#5�q�,�Z�d��ꍾ�e���\!�޶F��r�7x�	80Zh&؅Qt�gd�U�߽�F���7Z'�ۼ��I��vs��7V��z�la����Yu��vF�]3]oF�N����/	�o����m�s�ـ�G	�Q�e6$�5�t����R����4`��B�KG֕����xc �9y�Ɩ
��;�l�^����t��s�A�%Ő���U�7�K�I�P9�m�,���͑/����;����Լy]w"�:��B=E$�7�"��u�v*R��H0��=Z��n�Q��s��z1A i�y���:>�3��=�/�R>և�������35��]�Hx�s��NmV�f�{��	���r�W��\ZB��l�{�R�^5jBA��P�a_�Y\g7q��|�k�P���V"9yȣ�F�G��:����o��N����)�	]5a��^Sw�^�}2򆉆�
w�?Jѓj.�^wl�x@$�6t�
钳�c+1�}H��3p9�NBL�x�d:?
l���]���ڭ��o�u�I#T������yK=�Rc��˻��o�z�<�~�H��'�i��ʧ9�XPOt&I����,dnB���۾�4�9wn���<c�S>�^��m�᪈���/|6������E���(2��n�>pje#�}��ߪ70q�P)&��力�}��[^�r���}���v	����9��avWU�E_t��G�XbNNf��}Eկ�kӧ�N�/y1��uP�t����v)��A�@Ĕ*|�6�g�ɞ7.s��� �I����}}_;�_C�ݣkTeЅ��ێer\ъMH�s����)`��H�P�Ha@��%�������oYz��`���{�J܍wK���g��� �#����.x�+�����'�|�&��8���*%]�IF�hNe����[�u����c>Eq�3�f�ՂR�������M��tJ�S�'�|'B���MϬ]e��������9c�g1���0��E��r��㛛��W�~��:}Y7=��I�DJ��WI���Z� l�o{���ʱ�<o����������ۺ�G'��*��ޓ��Q#��
	i�A�u�<�r=���K��g6U�}������f�#�ɵ�L���_.{8wV7�Ed����R���Y��6��!^����~���W+BP����w����fQ'���D�
��$�,y��;!�eN�n�5�'��5��^�H�Im����q��u�Jmq��l2٣�-�u�!�&�6�Qj���K����8a�ae��J����{0V�-Dm�
9vU��96$3cD�,�!5�%Ѝ;Q4��R;7!4��[��Zʔ��ԫ�k �����ke�u6�lC��۵�̭��eҖ8)��H�Aa���o�!A�y%�����S$mg�����D�
�|&=HEw7����y?H�(�4)��5�'���s���;|C����=������M!��ÿ3<���P�^�$��߷����n,�&��8���z%w�p	������*��r"�o-�Ή����x�� Zݬ��q�]��:�!�٫�3�nD�Vz�[p�����6�b!(gp#���~�8xyr�7��/l���w���7$	g�����1�of)	�~�]�2f(��� �`4a�/0�~��ʒ6Q\eK������[�w�~fz����g�<_��-WV�4DaL{���>�Um���*�մD���{���L�a���^^J+D���5�~c9�2p�#�ؠ���ɶ��T\r��,ĺ}n���E�&��m_w�w���N�S#d�}�j��Bxw%�n�,�M4k�<�y�t��ݑ��I]K��Y&lk�����y.��0�O���{���R�険a��AY��q[=�g.��)�e�h�~!g��R��|ZOs�F	�/a�ʵ;�t}�g��'B�HF/�;q�>�x�����_TR]��r˙I�_��8k2�x�W��<5Cư���W6TXk��B�Z�=t��SpY
F��9<��y�K���ܭ��Lie���*l�H9��K̿,�ׯ_�I�m����ȣ�I2z!K�(גZ����03[C��:ke�nh�h;l�2�|�w/Gf�N�q�YL�S�*2�wnۣS��߼T�hg~^}�m��@�=<0�R��ux�|<�{�$��K�"�I�1!���w|���v���Zwf{��������:]���F�%�!�,������L[{~yS�#�ߨտ���G`�\���=ݧ�� �mϤdo���!�ŗ���8B����a3�[>خ��?!</�Y岂��<\���|~Y2��3^+��zr#0����m���h�&}R�4k�ޮ��.P�˘��[rZ�� w7uWH}2VZ���n��y@,�k�<0UR�ޫT��5��\2�yײ,\E�4�����e���L\_lh�^�ZN����W��Xj���+��;��`���}u�/s�Ui�e.�/5���Ax瞔�;����#7
D�rM<�Z��޹����U�c���}�z6�e�4��D�,2�wy����g��掗n����KL��Gm�:��`"��i��6�*�􃁷�1Ta�=�I���v�ּz>���'D���	%����@��b�Y�|��[R�Z�׶�ɇ�(�6jS�A�V$
^��d2��ݭ���AǮ��:�wO��L�9=(����(b�2\Y�+6�̵&��GV^�#��pE'�s�A�f�/����_���\����p�NÇ�>$굾=�B�����P��؃�0 $B��
���q�G+=�5�c�(�ːԐ���1U/���}�ҹ
������N�� �\{�g�ϖ0u�w�.�]�3���:^ͅϻ�ÓJ�-�(Ӯn��Sq2����ETs��f��p�|r2�ޚ�d��(?^��g-Z�+=�cy���Fd&�ZS)����
,T���Y[��г��m��A�e��}�]dv�r'�֞�DA3i��������i;�U��y�>lo�qR��wt��+�Y��Ǹ���{�Lڍ��;�sD֋KT���Ö����TQ_��V�|P��	�X�t��c�9���}���]ap!z�`B�PH�a,� �XMn�;A"66��w����8n6�����#�;��Lg����M�v��M�����N�I�SꓺfA�P��[�A�������0hZ���nB�lKlQk���r�7�kE����1�s���N%y�<�T�]\��������u.:�4�H:=��kK���yͥ.	�a����ϡ �]Y�;q��.���V����][S0�t�ܘ�J0s���Ps�P�4Z÷�/�Ú�#��uf�Y(hF�+.uڙ�pp�*n}��>G�ݼm�X+�p����;�p��Ϯ�s-�r�W[���Luk�439Zs��=��� ��a�B4�H��z���WOxZ�p읞�$O��E��c��X�
�3���,�lK��W��6�
4M@�|�L���@l��S �e.��a� ��
����[�`�{h�|�z��Ց�2�y���O������O����^�\��dx�g�Ό��E�^�X���m�L�h8,)�<���{�T��5MpC��Μ`ݜ#�Q�����U�vcV�Ut�Z���g��N�}"\����0
A�@��Z:�"�k��gz~�#�U,���9��Ic�s,�U�9ъ� �����'�U�3wr �M��.E�U	�HV�H��_�{��<���`��^�p<G5I����>|ȹ�5���2��w+�dvz��Q���Wu̧5�==��<� �-�~�M��v �^5s��hƴ�r���e��>h����:)�R��NU�=�]p�F��pة����gv�������b��So;�(��&Ba���좹!	��9�b�w�GF{�t���_��z�f�b?W{������
T�,I�-\ˣ��st��7Gc�vK@�-��6�����Y���:�3�\�ۦ_
�4�󌞴ːF�f)�)#
HxX�.�."C�\l0��8�5c-X\a�ft7f�k��IRl.�v���j�0Z��2�t�	t5i�Rh�`�zQ�n�Ĳ͌i�X��qQ��%�lVҒ�Z;�"�Dܰ�*�#kۥ�%9��u�.�ˬ"�0*���b6��u�q�an[GiFS�u�k-*V$%�]\�rbᵆ)-ƹ���8Ѹ�1����������_���u���$�r fO��>�v=g�'�beg���{���C(�C ����(�͍����4Z���T=���wq'W��>V�'�w��rf?q�)�t:�U@��Hi�١q�����4�a�/[��AW^�c��{O�c��#8n��ղ{��������t����,��rx���\��Ah�% �	n��Yxu�)X;�qZŋ�1��)��򵹎��~�3��ǜ�R�;汛*5��������� }\wԋo��^�Ũ���9�!3�웹�bs>��[��eA+�U&�ȿj�T�g��Pї*7����ٸ�[�yup;�qsj7w��b�5,^j�Vw�k��=���n��Wrf7�*]����T7"�j��*=�J�^W���$k̤_��!=�ϫl�q��lZ�WDR�ͬ�a�&r?���~&�wƲ}~�5�n>�8�g�����K�ݿY�w��5�F㑤�Q��b���0��un�������3ط�F>�n���c �Z�5�ѐf�<Ҫ��_��7��7��#+�a�$�o7ك�,����[%��= h�S7
�%q�e]ٔ�TP�n.��K��W޽��=�f(b�G�g��ۭIe�\8?�v(k�mee�>������Տ�n�<"x�T}1�=�o��(_7
�����Z�9(��L����&�h��}=�J������}M�z���m�T�/;�9�N.-���j���b�Z���|]���V��{Z���sLD�dp8W̠�M3�b�n����5�����%CI0���H�����o3i���x�Q����Ɣ�k�F v�roOd�Z!jsxL<��R�F�}�l�ݤF���:ȟA
l-qV/��䂾���ãk��>��͊��>��˿f:D[�=�W[Û�7�S��Gz.���>� �r���;�^�	 -!U�1i��*��{��u=��>���k2GH.ϔZ7���_�L_�����.��AԺ���}���K�T����DJu9�-Վ���06"�$���:H��\˜�GN�M)mFA�9UI,�^w��S�o^��q��M�zi}V��_�|36����u'����T�����a�8�a��|�-��mw+�93=D�Q��O�نŽ��W���Υ���=]z�v��F�٪����EZ5�/3g=$�7�75N�O��WTw����������,�t�Ҽ����'""���|�F��2E0Tj4�0���j�V;\�Ǳn*�8] ���B�$��D��8�n�;F�>�������F����&�8mzK������ۦ	5R���!��F6B�h��_
�7�Ð�}��V���ѴZi���ǟ~�͢��
v¾�v �f����VWg2n=�.HHp8�EP����
e,�xi��P��7�l��*P�u�Ӏ�3�^��-�T�3N���m��U��-w�Nn�����u����CO��Y~�7yQ��N��ϋT�kۛCֱ��Z%�{R��ԝab
�{��Z���!�_�����W�pu>����#�27|�7�j��_� 6.hM��V/���,�����+i���ٞ+�}cj}TC�n�.�_���Ʌ�R�k ���}U�竸�yr��_��t�i���� �jGv��c㥄�����q�_��=���X��8cc�fV�Ṭ�I�e���P;}R��Ι����]�6��jU�U:l]�e�o�z됅��H�'��|nx^F����*�:=�t�<�Τ.�j��-l���-nkm��m�wa'����*�֠[��nI5�{�|�U��s��������8-Q�6�Ӣ�ƹf�C��Γ�g��yyr�,��\*H)C����{'�6�X�7��V��0:Q�:c��&�i��ʚv;O��c�GM�ɫ�ͽ�NJ�rP�Ff��_#Dn�6p���&:�u^W<�F{�'�D2D��٫�cI=[7�w�ՐDц�9~�Y��]N��o�T�tq���ӈ��a��%Y:Ok��+�i7?)Ȯ�X�gi��O-����F0m�e��Vf�	��3('N��U��[�m=I�,·����{n�J1Rl�(��rv�/���5�(�外��:��s�ܶ�gaU|��]ܻsq��n��Ʒ��Ѻْ���Zt��S��H©f���� i�Npu�]��K�d^��b"q���oy,�l�=�3;���Y��k��,l��Lʽ\�<牚x�-=�b��e1ǵ����Ak%yJ��w�6<�M@��:�{S������+����R6)1�io �V�{2�M�鉾��@��ǵ�i=�味�GlgN$�n�ۭ�:܎PB,�m����j�o7��{�+�WX�%�Snm����$�N^�n�kT�U��f�;)�#)�;�6q=K/F���:9�m��g�v�V����{�wݕ"ȇ��w��\�Ws��K�u�j�e��D��;�^��%j@k�@�v�
[�ஊ�f�-�è�)�Dh7�!�x(EJΎ��ya��)q��:��V��@��q�+�+���}(�h�k{,��X6����Pg��jJq�J+��.�/.���Lw�+e��jB��2(˛Ҳ\���NR*�ou֪��rg�:%8�zV��Xޤ�&�K���Ƙ��k���PN�	~�Õ	wЬ�b��/�������]���'\5�Pp��tnݲ�:�Ԫ�b�.�Bt����{�#��fFgws�Ӑ<9Ar}�=�D�T�h[jr����kכ����@�7+�>y�4�I`��V�>7��t4�0_�8�sˬϯ�38c+i���\>���`��`��'$�#���x�N�Q=�U�<����I������7�� ��SDJ������T</7��Ɩt�{z�Ò B�F��w��L��i��^��,\O9جZ��pW ��W���z$ ��GuK~�{�o���Am���q���r��nz�^����&�b��(���jm4�+J[�^��F�t����'��q�/$t�[u����m>9��PL&`�OWb��?=���t��Fs�}>��2�T�a���y^޿7����[��M��n�^5��E�����j��ں�X��{-��,��5�{��<���)�ڊM_Q3��~��u}S|�hH���,�Ogj�Q0� @�1�2�|U���y�8|�[��{1��c>*�۟ʝr��[�_{y�W�=ֿW��l��}G�c-�h�A�G.k�O���y���	0I�W��ʍ*�VD��*��x�r��/<�>���{&iG�t6�2��B���c��V��4���Օf���*k1�уc��E�ʓ��iT�`0�J=o�b�y����C���@$E$�����iv���Q-�Gl��y��[�&��	���{�"���J�2�<�ۚ���s�*���	�.�&���8��XqL�[�;�'�͌��P�g����Nѧ]vmmġ���y���o�T�G@7W+�9��p��y"baj�>��R(������]��[pX�]���k�5��M�������#�-����~o�q_�/O��Ix�)q"��q��Jm(�D�M��$}<'/�%	-,�l�:�`i�����螪��K_*�m(�������d����k��_io�m�nz���uh���Q�FF*�y
��.�z[�������'�)1	�-Y�'�ל��=��L_F��*=�����~�o�B_LAR� ^�1�����[D"�
Mf\ٳ��ݯWaz�p�`�VC��йӖ�-6d�Vk�!@��x\e�L���x[ҫ=ʹQ�����~���e&�D�]z�ى��am򼭱Q]�$��ї[ڍB��j�e����xFr>�ܫ����;$r��1�(lv��[v��������4`rS��|Rʼ8m�S�bi���00X2*����tRU�|~�sy٘o�>17d�2�����9C��|0.�w��ӝJ�/��I0ˆK.�V]b��zOu��\�%`�:���z�c��j�2w�q��
W�Y~�s���=&w�}��Gٕn�!�V�x��Ꞝ2ﾢn�)$7�*M؏ioإ���u���q��N'��~,c6=\}&;��u�x�n�x���6�l����q����eG��绣7gb��0l��lU������u
3/��-#��.	������<�~W�ޛ��{��F4��A�܍���)w�����*�����E�l���WBj.��ǁ��;�ړ�x�q8H��Gi;W<\�n��p�Q}�׽�W���ʧGc�^��Ņ�HF���.���}�!�����P���k2�>B��#4������2W�MU�y���$�g����&/k��y$]�,����|���,����?Y��~��mϖ���G�A+�M�}�ǦsO�e�߆�S�b��k<dD�Pkw��b��8��h[�,�������{� ���|��y�QxuC�;p���F'q5.��G� w���.:�I%�ٵr��߮�}S�z���`�{�9\߼���z!�Q�&?>!3�{'�D�;��cx�3��E������^��G�x��&
-���� ̺�����3>��^���� �k���dSš�d�~�z�,u������U��Z���#����.O���A�>I��h�ᚺ B8l�i�<�ܪT��W^Z�n�\���֢�'lgzbj�s����!���4�%��h��/�R.3"ew[-9t�Y!��A���04�j'o3M`�B|�=�xפ64>�ɭ�d���xM�OYY�oI��V�D�W�f��k?I3uݳ�X�sj�4(�Z�6�jSv����J0 G+�|	���P�fھ���Utsv�dQ,H���[��ڥ�3����z&&��{��FτL;� ��Q�s�x���2��n�M���>���5Sۣ�g�j,fr�; 㝓W�����N
.4l��>���w�tg�]����7��ju����һ��"��V���Q|��s1�W�ǆZ����ק���9�Alz��`�de_x����`�fz״���D����������y78�ǭ`��ӱ�\΍ý��j�x�zm���d[E)�v8��;��		E�2�Az�2V?&���,7����~�������9#nIX<&����}�6;W�풠��`���d���اV��Ӄ��8�x����:)���@�B��'�Ͻ�3Okh�CDm/q�	�]��EP�vٹ�F9n9�a��Ą���4EQ�3m4�SB1	8%���ݝ����Z�3����TG/�;��!M��5/��.��W-L,��Tm�f}];�f��P �6��6��v}��9��lt�p~�����Rt_w��i�-�4�>�y��X㉁@�� ���H�?-�t��Űa�CA4����*��	���y��%�[�˭+�6-^�D2X,5�ͻ�a��*ڇ�3�e��v�g-V�}+��+aJaݣ[�_r��	r$o�36�.�.�<7��<.�m/oe��Q[i�������/P�AJ�eVm��$�ٶꮣ;��a1 2$���:|�����*�p}&���T�l��͞_9����<W���b^xO��K饄�=�L���b��U����3�4t��!��TȿF��b�u���k��eA�Q����=���Tiz�JqxMν�z<��\�p��Q� ܀wlg�/\��pĉ�c�{��_�1p��nPW��`2�p3�K3��n�݈��j������o��� � �@�M>9��z�����o[��g���B��D�$�s�n��!�vb���/Gej�?J�!��>�Sw�j��Q���������>S�s���/R��� ��㧒��q�4';�3�t�b��X�{�}9�I�en'����v8yN)��iu�	��A�|�Ӟ��vw�/���z���"�l�\a�s�� ����4��FzJ>�6�-��4�����x{f݃ݕ8���~��>6���!{;D�-�aׇy.�ٕA��N`S���� ����f<4�B�I�گU[����J��:�̌�}���*bk	��7ٖʴ�Isu���T8G �E�w�f��=��M.�F�ų�G��*�8���7\W����>�v��ԖŴ�r��[;�i��̎��pZb�0DE�%#lZ��,!��.�b�t����K�g0�F15���x�JH�^w�Ѹf	�U�`4�.i[�3Aїb�hq���ۡ�TI^�+��6�ƲjrK�m�06����ƻiS�\A�^����� T��^�r��]s0RJ۬Ҵ\�F0#[����cT��m2E.%6�p���N;��w?/��S"v���h��S�u^<�$�^:�ܺ��;�"�N&C�
+Aλ��W���#�}�5?P�~����z/?S�P����{��#��ɷ/�7t�{��֩�P3ܾ���/s�%��)�I8>��O�`��~qHe�b�Y�Tь��ǵvn��6�+Øp�	���2�,�ԁ|�N���85����<K���J@Sl4�Lv��C�аf���:�������d��d'�h���.��=۹�[D���!�$8H�����,�u����֤�zOd���7Xr6/�{>~�������V|g�f������9(��F2���{%V�O�3h�$ǖ���E�e��Q�� ��L������.nB����`Koޕ��;~��)�@�.$M_6F����]z��wiy�ޒ�I�P	�L���;b�յ-.��\��>�Ul7Ʀ�ץG�˘���k�P���G|_���oj�aV����CO�V$p�خ=R�]߼+sA�@l�jH�"��-���z�w��߅w���al���)���=��oO�yw�ҝθJɾ��7����k:��[5�C�s��zVܭ�Et�7T���.�����:i �Y��7�G����C�k�!S{f��I�C�}C�<�"�0/ވ�JA�n�^T)��;��/�����}�f���o�C ���<<��P����,`�6<�]� ͡n�&A��A�oQ2����,BV�M3�32�=vƛC�tЋ��f�<b�l:�_.α:��.���z)�n�\�l�%1������d������+���ᆆ�Oz�fΣ�_}��;�{o�X��K���mw��?,��	M�m�혭���l��Aq|�q%�uVmU���S��ŕf|~�w�{�O�=�'?a73��O8X�3������ry)���S��zX�g*��sр�8`(b�	�?>+��=�|��HѠ���/��>}լA����H��~�����*q��~:L�2�y�iđ��w{*�Ąq'r&���w��Ef����w�fgaR�s�J�)��:\�1�ު�F_c~7o�|�1R.�~�u[��Yp~c�	�{�Ӛ��yA� 2*�t��}�0�f�N_q�C����yM4��1c̭ҩ��FL���m���U9dT�i�)���w�S��po�G��6�O{'|)��Bv��������9��jV�X>�d���ꋖ���]P�kQ�@2ҫ��ݖo֌�0��1X�)�t���z�9I�eɛ��fѠw�.��)�9��ۇ�Oy�s&��"=��$�H�xx-���]���s>}��rv`�fd���};�W|$}�KA��bj��������fu�:��U)Ʀ��������W��8ܧ�MNz�$�KHL&�2�������m�(�L\�I˭��1���]�r!QC%xJ�ޤ�t:3�{S~,�^�s��m�����rH+�w:f�g�%ɰ���'�9@r-�%���aL�:ݭ~﫶7���-<����/�k��j���w�9G�L�"�"w�V�K��fZY����;����-�%_+ɛ[��}�<iwf}��{<�nfv ���lo+g%Y��5�uʋ���d�A*�K�w��B��t�:+�����<�`v-)��08`J�G��_�Ɔ��8�!�]c�>�p�G�ဂ��.��`[[Fdэ4e �l��p��඾'�%.ʭQ�ߥeO#�;8v5C)M�?��1hN��G����v�fn��U<qՒmA�=�\l	���r�Y:�?8i��S�,�S�F���8���w��ɟFp~���'��+𹙯����}�̃l>�?r�>��2l����Yo�'�'�	;���,:�%�h��C�b�Z�p&f��~��E�4��CԤ�}�.�b��չn�uRt�v�P܍��v�]�٢ X7Pʃ��)õͥ���5����
��	�j��b���E��1��kf�������D]��o��^����₀�h��d]I9��!������FN.���ש�hN-Pgl5�.=f�R�&c��R��Z�)�|0J�פT�A�0��O6�U�`9��%�!&�O�����A�W��	�=�SN�gZ�zg�zɱlq�����Q���>��������
�f�g}]�J�o��S>��o�WE�s)4>+�X&�Ұ|��;��!L�A��uճ]3��9�sC�Q���i��IHDG#Rm�ҭi�)���! �m"n&
Pb�	e(z�9s�3�#D���.�yW�z��i��} �,�M�,t�����3_���pe�����0�2���M�*]x}tm�w9|kI�=g�I��]_o[%�����(��s�M'�fF���kK��d���7�7ˀυ���#V���S��0�e��x,+�rC�Y�m����1؅i^99��-r4'���>~��E�/�ɋɏ�l�)�u��C}���/Z�5��7F�d�m<=��l6���Qךo�5֊�o���Jzz�`�]���\s� +���n��ߪ��a�Ɂ,q،`�
�n�g㲢9��qEq@���wP�t�RN&�-���ޮ�B��b�25�T�j�M\u��.�H�.����6[#.�u��8��b�M��h�=�J*�|_-���jT�4�[<��c�ŭ�&KqX�9�-4����[k��O���]�����6��N�P8�J3��0��K���j�^�f���K[<�`�p�lt�뤲`�)a,κě�Su,*4.c.kssKv�	p��n&�`L��`A)>�:$�t��ß�,p�"�d��:���<*�杴�$#�ML��riÄ� \8,�SƦ�/��qu�+��}�?���#�|�O�[���I��s���H�y�;�w^���w0�^�1�4�z�¯fӮ܍��Ԅ��)�:'Z��?s��k�-h�6o�{�v��y�y��Ď�E6�Q�"�ŕ����mk��0ܙ!�0��(�d�����e�ݥ{�~hr�\sl����^��f�U�u��{Ǟ���ezq�Fq5��;�sL���&�=��Q�25�{�F�w\}�o)�>o�s�J�f$"��8��	�5�(�#y��{�\^;c�=o���l�?_^I�ڡ����&�	��A��@-V���~���tv:�񇗔��!n�cӘk8̓&+#Y�n٢=�,�t�n��2�k�?gH>�U76���霾۪ߥ��#�	q �Sd�*2G�W�Fw2���|��K�z�����:����/#�3��kЗ0|Nr+�t��_���o��Oe��V��p�fe��w�v7�g#���4�ז�����j��N�}��K�s�n�-�V7�{��L
.���a��U	���Z��wƅk�g��[@�'t3B�=˩�e)�����HJƺ[S�I/�t4`�N����u�71.�&�i�ѡ��t�������+��Ir��7����𱹭�c�f��Q�q%P����*�q��	����y��2��\��R�A�iy�ՙcD�q�Η,�����g�R�wc�XȖen�(Um'�R�DNܜY�NkI����շ2�$X+���	j�F�~�Ȍ�N���byM��7v��P=g�ΛĻ�ޢ����oO>z�\=�e����/8�L��fk+�]�w�Q�C{�lR�f��W~���$sNB�H���� �Vm��]�ufW`��V���O+�ɕs B�(G�y� msVP�̵�Nw��2��mEڋ�����|Α�:5ql���t�ν��3^#�����]���<�g!�#4*�כv[�C�V���)�s�[}��A�fI��k�Uʇ�-
�Y2�R��A4������0��T����5j��u���;:�Yv�"Lݨӝ��
�Nq��LiV1N�9��h&��Hq:��U.���1��ekj��{���c #)�e�j�e�/`�3���Y��Y����i���L>p^pHnM����;ú���5
ʾ�.�ݐ����!H�����g3��k,w�xm�#V�ᬢUZ�kX��]N�5�%�R�zc0b<�4v���7F��{��q�E+��"� �܅3�M�]�ㆲm��//sJ�+��D��IMuU(m����U:)���l��*�Ԫ�UU! �EJ���iZ���U-���x ۈ��5�R��E��E�p�t����VwU�u��ugt�9�U�`�V67[�����8m���qֶ�V6�	��K�µX`��k��s�mٰ����Ovmu,;v�E�b�d��N"�N������=]�1<R��˥1v�d���7A���{nݓ���6N�"�S6:5`��bZYv
���(��7lRۂ�Ch:t&rm7ibJ(ꝥ�x����UѸ!6Ƹ5���Ё��Փ.�u*���5���&����F��9����U��L�ԫ�,��x�֗|f�p�3O�Cڲ��\p������;?������Ym���&е�)B\��t�N���s7\�j]e1�؜��8��	�=�c�o<e�8�⌸�>98d3���szv�R���6.����%��M	���k\��F[����2��]&��v��,��dR���Mv�Jl@uѱ��/iA���p��^��o��֎g&�6���!�oh3F�{U���gsT�)nh�q�!���kq���<p��n�\����d�n�[�Rŷnd�Ĳ�rhg��v����7� |n�]<��/	�T!$3�&���t�e�mh��t�v*��9��%���8ȡ�0�1����ph:-��[w"q��`��ݭښ��U��Od9|Bik�*�$u�E�,�`�3�A/��5�4������Ko3��=[2�p��8��a�si�����]�!���K\W��s��b��$�z��݅z:5�M1&	k[ۭa]ڡ(�[-�N�{�Jlz·�1jذ�V�v0n��^��ہ�PlU&7�A�X:Qz���&�̳Q]j��6��VT��]ZX�i�Mr���)�Z��9��7=�|q�n��(���1r�cr��`�;2��L���D���rv-;#3�� �H!3���͹�Jܰ-5��a�z�qP�Ȃ��B�5��l��]�/����ǹr��� �?3~��/������^���eŠ�[�3x�b|�e0,bL�1	-6�/)�[x�:<ZW2���-K��D�W� �����58a�x���:�� ���~��~�lXaTvU[I^�ίe�7�+�%C�$Q�45���]׫}�N���9b�0��;ݺ�����%����}��B�����ȣ4�E��Q���'�95ޣ�ZQ���h�`��A\m�	��/&V{�w�(��V���<(�ߜ���9I]j�����d���@�68�c��5��*�n�ڃ9�3	)��}�|�:&�GH|Ch�,��95�[�9b�>�HG���֟\��gϲ�.4����[�k�
�<�ȿlg��k�<'�<�E[��Af�3�|3W"�Ml�3OI�eV�Z�x�&UM�����PC%��x]�՗�ͮ���1!P�ot��w�]��.�[�]�s���.Qh�4��0i����.��Tb	aH�j��sZ�����70�J7 j�>���vJ�AJL a8��9�E�@mGc
]�Ν��VȄ�5�_�a����5a�c �YU�T��3~=Z��C�g|��γ���j�{[*xz���^Yt��Ѣ�*@�̮u 欝���̆RY�+�Y�ٲ�[��l��)*��04���љ+-����rW{«�4�H�e��''�/2�i��@}(a4��O��ʬ�1���ʌݘ��]��2�7���0uӿu6�Y[I���p��#�p�͓�0�A*�LS7ڝ��z��`L;�BDI�Z�u���zx��19��zk<�����]P�|�+NdD<�����.}hM�l� �h�`����J�7���}��c�4�nL=�zM�˝T��
���se[��f�{��Z^g%r���2P��+ i�}}P�0wCa ࢡ' :RDh���Uڪfem��г�\�nC�0m�W���y�[5z���|f��ΐ�f1�u[�������Ͻ-���d�ANt�f)%��o�Mf��(N��ǭoX�U���Y"\pCH��2)���,�Ǚ��%%���fP
���$�&�gw�� �?��O*�v��>{4v��>��|���?]�1��_��h˼����,��Mt�<U�W�,R^�5�+M�����^ʸ���'��KEZ<UVE^���\�i>�j��os\d�wgÐ`�6C]h�srul`g|����x��b����V�+ꕆ��ij�쬺tPL��Fe�ԏ"�BZ!��)C�t��d��S��*K9R5�gdeA�$mt��M�s�m*)`Q���o�ǵ�f��2,�fy���F��#���HC=����n����_(l6����,� �����4Q�x���,C��'���F���&$y�0���
��V��_�^*�*ϋ�{ʮ��`��	/��W�ʒ=X"��d�1|!=^��<�I:�%Av�`�u�7���@��}�3���,g$��K�7t���r�R��vU�җB�2�{g����n��`�nq�C�8
R�c�Zu�L�Z��&�^�H�d�5�5�
-���E��ˍlŎ�J��A5!U�M�u�����o������is����$�z&��c,�/���"S��k����I|$��h9��Uӓy闒Ox��SUw�{=%:|R���<:��#ze�I����Tc��^r�uM�U���*N�뛗�}1~�Irh �Yp'�=�s=;��<dog��g+��:��_����#�P��ݯlC2I�3]Ӏ��<�C��8rv�=�G,�̲=M:4׆'>:��_�[ʊ��~�V��w3����Ns�7&of�Sy�)��</n%�|��/Oz�+�d�FeiN/#VU������� т��5F0Y�	�Cnc<:5�u���͕9��^��R=5�����/�����V���qюK��4Q%$�� �q�7:z����92H<l�Ϭ���o"i������Y-��y���!��g�W�y�ݎĝ�Nup��kJˊ��A��	,�-�Du��c,��4��$��k��֣�9�j�/&z�خ.y�G�A���ӕb�I�<�o�ڻ\u�\�6�5�eٔ�7V�Mƴ)2��V���I�ě_%#y��Ã8�ng����`�S�����R�6=� z��I���SY
�&�=�vW���V�l�@@��)��Hܗ^,�Vm
O/������>ҖVO�ˤ�ݯ?��k^t���]^�P�k�wC�.�۩�&��w�)=���Z@6A!�I���a^b�=��8^�=ey��[�4��O��:���-c�r�R�a���AbW����ʏb6k�(��'���w��[t�Ë��(o]�o�H������̵m~O�Ͻ�vXh\of�䢺����C��V����F8ٵ�=�}�3s�m�.?g�o�� w�VU�͍����}�-���"���nw��69H�Qt�j�lna��a-
�3f���uO�UYp�+�{����d�9��Ä́=i�h��c���YW��(X�dŷ}쨆����қ��K�U�C�wdr$��m(l���T
���T���Pax�uܫ��zN�w�.��^9\��n
��͕�^l��u�j��WN�z+�TD�^�}lMGn�M����)�q<"�����l-����w(������[�v��;��vX
���B��\"�3�>�)�ѝ���{��Gmc���l�F�����H��Z�:y�闖����cGX8w����Y��͇���u�oA�SP�ɯxO��A7o����pm�S�WD�޴n{&7��	�KP�9 uM��`�˛��O��u����^�u�[�����&5>JZ@��D~j2���̾����K]@���>QBQ�d%���y���&W'd3��:�x�e�=p|'�c��>�=�h�?^��;^�������k��o�r0�o+��6��;��k9[�������*V�S��sѱ�ٛ����Q č��=��N�+�����{�r����3�a����>M�F�d�ɐ��;�ִ�{b�9�
ɀ����4��Y�i�Ůs�T�N�C:3N�Y��N�u���N<�}�Fn?oLmѿoo?v�@�a�%2��
��!v��]�=�N������a���h�����\�*u�8��O:�^^U'���7��1�ɸjo��ջWGӊj��[W��8l�D&	aR�S���ظ�l��u=3&��w�ac�?~̹���S���>^y�) ��zn���{5
^�yQ����h�<F����n���ab0̎��r��T�A:�W7z�D����ǳ�3Z�R	�2�Cn���o]��m%oA���m�(x9�E��%��ϤAҺ�np���D�YC�MFk�z���@~PB!Z.��]woq�w<�F�G6w��.S���}��J��lx(�S�udG��rE����C�9v-$l�L�}�������3;��F�������x�(x^j���lǻ׷�����{'�G�d.���w4g�wCn��`m�Gg.�b4
�{����U"=o3|8�A�u����|đ��2I���Õ�+9ʓ�~��*T��nᗋ����vL�7��_{�9~O'x<���=�G#���n���΂�5/r`\�a���6XfȼH����G�w,��ɢyǳ�mf�{[�3+�:���"8wdC��g�.G/}ѷ�/��V��9�|�lRǖf�:g���˾r�f�p�I7A����#��3Q�8T��&����玫�"Z�F����¢�Q�o�t+٭������tz'VϹ�@��NO�x^�Z՞����LHM��F��	�9u�4�PF��ڻQѧƺA�?)�)��m��t�֤0���<X�ȝ�f�f��d�gw�i��voQ_����]F��)�w�q��d�j�SƉ���	u��s;�_^�:���M��3e�a$� �&ۃM��Qx�]VO�)���Z���k��̆< ��Q�;�V@�����MjdR�Ͼ��ܨ��k'�
��|�xdޢL�_(h5H��/R�>��\#At�O�#�՗��&�]�h�\S�3����FzMNu�ř����# 2oo7�QXy�m]i�m?�#�����oR㵙ѷծ����m�W�U��e�d0p9�Yw휤��w|��?�.cD�}�w<�7vz��[*���O�:0�*I��-��OBĄS�b��d��5��Z]��y~]*��Z��޿|��c�_��������%{&6��n:Òh=�쫛��������4��ژ�{^�^�~#A��[C־�`���+a]��mn}ɻW&_!/!���!�rP����a����:x��B~�x���
�=�Y>
8��×|�e��q[s���&�%
? �����Q�ūu��w-�v��_F��/F8��bqx+��7e�)#�L�i3"��d�=g��[:qr��U�Uq��s#���g�1��\�w��3�s�|xt����qV�Do�}�'M.���M��W�)�0�	�V=�k7�u�v��P�3J_n�,���o3�'�r�5���e0Qi���}��0Ɖ��W�u-VL叴"Eƣ�o�}��2�0����������"�k�_���d�)}R8|:���3���A-��!�������'�j��Z:���︺��]����A+��S�d�މ|�q�J����U�.�.�K	�x ����]ׇ�ٵ��9&u��p�%]�9��/yRz�蔩RH�X.�ِ�sy����Փ�qq�v�ZNH���a���cT��Y�[�a.WM7#v)�e/��o���tj�8����S#���s����4������K`AڏX�m�eyݞB��0`�&�=��帵�����@����grm۶V�uLz�%�6 ӛ�:i����^�5�D�3�K�՝�蕛�����Kb C�ZPOj?�Q~Q�7���E�^�C1z	N{�{��(�G����3�8�i]+�J�U�x��7�}Su-vm��]04�� ��7�]��;'�ŚW���?uI+�-VZ��s|�i�˖�o��S�ǳf��Wy���D���!Y���|�>5��\q��u�t,U�\�o���]=2��e�����b\b�Q��N�M9琄%�;՞J�a�W�oύ����d���]����(p�=���'�N{�_����Z�gGŲ�u�{FZ
`Θ���+�T�����߼���og�w9u�7����y$/�0Fr���(��B.��v9坳����:+�#���p� (I�Iѻ]�d��Q�x��&�����&�|�Si�{���'�K���ەo��5i�*����7�^��]tl�F��G+��j�m�WXg��j:a4�_6�3�g) {uWz.��b�ֶ�0��{Tq',ׇ�B���V��:�ՃG��t�����Q�������<vqig�pJP�mB�.b}
ƾ�=����oVV8��9I(/Ïx�2?�&x�X/ō����b5�����y~g ��m3��<Qٙ�R]eb]R�������+�	2u�ř����l��X�����VM�)�%=�4�Tjf9�$��*7���&R����,��q��k5���2�Y&r {ڸX�kw|cW�Y�z�V�r�\���/8I��B*�D+�5qv�q�e����{u�Z������~�8��.�W���^Ɔ$.��u.9o_�([��˳���4��(�|<�b�7�%W��=��\ ��P;����9Rۺ�s�[q�i�8uO�dP��h_�YR������X�g�ɠ�*����'�lF��g�]O�O���G������.FP
���]]^CD��o��͸�������7�Z2P��@_wq�ې�\�g���ڢ�vD���m���bң�����Q�Fhѱ��P�:�x�%>]�$�U�>ǀ�PvR���*�6��q_���zP�0N�'�l��oz��T�K����|���i�0$��p��M+��z�=IØ4?�١O�:�N�X]ulE��aW!k�}}R3m+���)]��i��߫��-��l����2}\+�gk�i��)��1B�4���О+w��ҪZ;��)!E!��&��&�[�����	���{5Z���6������&���������p��/�Sc2{k�xk��t���/X�`���<���D�u�Z3j+;+m�]�滻=k��*�U�n� c����X��̵�C���Mk��1qB	U&��g����f�G��Q7�	���}�bf�v�~�����]W���X�u��ɜ3�%\�s.�����G�ji'���;��{f/����	�P��2*���.�5�̝,۩�a���{>"lۯ��ċ�7yM���|=��%8��\H���7�OE{�u#6=[w�HS�7�req޲<�(���VT(�B�BP��,���٢ܥ^_n4ϼHy�yۚW:;&�ȋ�r�����;V�@��!C��G,���y�<fME�f*_q�~�=�x��!�a'�$uTb�0׌�/�L�:� ������}4�p��<�����G�ݗ�.n�B�^�&7W�<jMv�����9�+�V+���!&����X��5�������|=�.��ز��u�8�0������;��+l�T1u��Y��QI����-���ԯe�3�)@��(ﳴ�>C�Y�s��Ӵ������/N���TIPc�x�&r=���vP\"�hԁz�2��~w2�<�(�8ݏ:�Z	�����^Yxf9�0R��3�k�+�V�wN��`*{����F{v�Vf������Ӿ���=(�|E����A�^�G)���ӿ{��Ak�y̺(ѩ�ɯ;���vV��{<�T[3��S�ɖ���ӭl����%�U�#�K#���U�����l�Tvy�^iާ��q�I�bQ؛��p�Ʈޔi[�NeR,h�"�yٯ�-㔺�ol?�]�q� Z��5��Aj�k7"�}����4#��)�c�pPT�4]eZݽ{�҂�3����>f�7Q�>b]Sh�\�_:8�<c.�f��&��o7\�Г�e��/�r�=�T��[�&�����)y�\fkozv��\�X%L�+X���Π:��uҭl� ؍���js�j�Lh��f\W"m5��4U�FoF��t��wr=�$�Z��l�.^o���荳���^����g�ٻ��iH��q��PTj�[6��]c�Ju��WݮSf[�խ�y�.㑫a[�2b�2��o��-B����e�� >G�-��r��Y��=��,�[ZJ[ױ�Պ�TMa��E�h��WG�$u����oS����!���]I��3m�놙33'�+w�&��2�^&m]�t�'ux	#}�k$ϥ�Ji����v�m��VۥO��^�.�2��d�],6/p��0i�4��k;�Z� ���V��Su�[}6�*�Ɋ�M�N�a���Xo���hƮX[�����]���_�5k��x1�ܢ5[��󜶄�*^X��T�}û��Q�"�i�÷:,�Cx��մ��y J�Qǽs"�=j`�m����}�DFc*��F�������=�Zt-��Ÿ�<^%�P`]I�{>h�y��hZ��C^����@$q�0Zd�������voKc�9.���-(�Oןq1.��!���daLgz��u`��vh�7��趢�|I�n�.�ց�t�XE��"���Ɂ�>����nl���Z7��"n�B�wA���=~;K��o�Vr8^O���r٤E��Ǚ��=28��Ɲ�YQ�Q�}���O�~����}��l%#-�IgF�j�n�]�갌���Z* ���� ZPa�`��`[���˩�GD8�Q���ӹ;��rnI>��_��J&��S<V�(|f٘�3��|_�n/�M��H��Ӿ���;����3Sz^��w��n���)��
���ߗez�j����Q�S^{yG���B�=Da�ɣ�_��Ѫ���$����s�yS�J� ����3��ҜCp�~�0�S�+�|�Z<��>Xuyr��q���Xw��w1y�kc�������n�֕��P��L�Ӽ%<��e��Y�Ƅ9v�ˮ�w�[�J���q�d���G�d%�LN;f����ra��w[���q��5��C/���cݥ�;pwr��qmW^l[3�	,4o\wIa� �/����q�6��r�3�����xedĹ�2JwN���I$�5h���g���\��M��t�kq%luRU0v�.!(@��B8i˥����|����[Bڈ�ٱ��)�pI�<X�a���d�&�"y�����Nn�#���Pb�9b�ZmG��[ļf��ؠ�=�8�9��&�J�n2��7OU������jB���`M6p]bֹ�U�&f�16���ZLt�"�X�hl�>�羶��}\w߿��hxd��}���^�o����%{j�C"h6�$�,���ߍuPn�$h�dh�7��vw��O���^�Ҹ4ld��^SiQ޵s��>y�N��s� *�=��c'��"0仪��./y�D4����)Ĭu�ŝʵ''��	P�e��EE��l���y��JÊh���t5r��^�'����@���ÄH-m�JW�ٵ��,2����L�#B�����ş)f�aR����B�}7Fdn�ϸ��'��J�@��B���H��o���uy��}��t��R<΋�j�6�}�,y2}Y����Tb�g-�p�Bu��݊����N��t������h��{+�g[PՏ՗�};{Vb�M4�2͊����S��VGl��TL��L��ԯ^�O����B�.2������ػ}�i������e{g��S�P^�v������[��2'yEZ���۱��h)�!�B6�H�f{�p�V�j��׶g�c�u۷vK�y������WҼrp�_t����70�n<Yo]�n]s�����C|)�H
�|�,cX!A�5}�������;��JW�(X�;9�{��t�	�}��0nk��-8m@i{y�򼹰c�O�^�"q]g�b��:F
%�mtv.���½xB��\��h&$�ñ&٘�$2Y������2o��YEvw�r���]ྰ�9��y����I��%6Z����Վ��}U��g,�?b�������T2�%t�L�n+�j}��M=7kɋ��p�}9+���JI�g����^fɰ������We)Y�7��=�5�|�?(Ў���3�/{#ruYe��K����ɥ7�0�cP	�h�@'l�]m���ZSO=�u������{vWg�ЧIE��N���W���-)q�n���k+�="WE���_ڎ��aLE�2c�<��Z�"'�v>���{�h<϶�6����Wθ0�T<&�&��*C�z�* (\��e>���B���L+o~��x��bǶ��&�&�/�B�&T]�<��\u��W��2|���u�&���>8u�a��Y��t�
Ү�L2JF6;/���s|#x替=�u������Ϡ�Tz2�8~�oT��O�}�JL���5�k�� E����n�jӷ;49R둈
�_@�*���L�lm��/Y�LtwƲ\ ���{�ve��&�.+�ѯVȄ.�����V��q�~}~���B�aU,w��$������#�^q��G�y']T@��C�36P���']�V��F�m����>���{�mw&��oG�<؋Ә�Dd�7+�����n�o��k=��[0
-�ZD>�-�@�[�������s�}�����j}�~������u<�fl5��:��]w����dFw��f�-�cЪ>8��Z�p󒾝E��]���k^���� o�!/��g�_/z�w2�2z��'/Ь���k�'��)�M%���uݻ��������s/}g��5��B:j�]i,vJ���04�ι��J�s�!�p�Ɉ/�^�ml:;����L����ǝc�d��>�Y��\aK���z��x�^N"Za�K��������w����,���B�]Չ���D�|	U�mo���{ۓ¢���ˆ̛��@E�l4����|+�Դ9�"�K+��G�xL��1l��Y�`�sqc�fIW��Y��]_ /�������S��WΙ����b��s�p�KМ����n�E����_��{}w�s�׺��\\]��)�x��G�K�Sޯ�p;��d��z��*� % o��N�n�b�}a�u^;�x���~=��c�+f,:��_o&0/L�X��F;�=Sy�UwGoP0�%2t����]9C}f�|�Xѻ�*Q�쥣��\l�.s]c��硦-����/�����Z3˕.��c�����QV������b�B�]��+�0�`~|�e"�b4�Q�%�q2̒�Kle.�+�fMNM���C5`b�OD�����=��:~�~uñ���6���t��6'������ff f��;y���5���X��l_��{/U٨�^տZ��>ֽS�zrO�48�q'�)���ܽ�2��X��zA����Tut���SH�A�ܑ�Td���~|m�A�K5�>�OyxAQ�;ܲʟ�ⳕͱ�	7�A^뺻��Nf�WkU�#� �A]�J��Zx~sfу�����y�G�4�ZU�g����Z�y�w�p�9-��pR��o[���S	}���;=ƳN,`�(p��e.�ԽG�v ���L�軼�u�ܹ�Sn�$T��9z��Ǝ����v��X13*ZbҌ�����ůƤ���`�lZX�ʚywυ��lp����ѕ7Sϰ �my�ԁ�Ƴ0�͆�ҧ3,�8V�Ҁn�v��D��sƘ!T��R����͈�^p�(�֋e�hdŷ^{pm�	Cۑ�B����N-�KN�V�g��v9y��ko$�f�X�1vrF!�� wߦ�T�l��ƽ"��zڑv���4h�
�og���J�-��lCH��D�/5϶������O���e�tF��t�������2*���]��Oqdl���u���1Y;�������l^ 6	�E�MW9ݗ붣Ѡ�A����Z�FuD��K�m�
�-(���kmC9l���F�q�:�1��W�ǫ;>*Wz��W������������qv��M����.�9�y�J1��$qFӉ0�z<~SȺ!��4��Wofd���p�e��O�"�\a���ˈ��;��D�^P�^�kw@��'���"{<��@�w�#@1jWUOu�_�JFD����ʩ����Y|u1U����s�WM�bzJ�k��Ƒf{����E<�B�ȟ�fg֖.��℩h���y갳0������h���v��Օ���Y7��~�V���L{�!��O��U�7�jȔ}�*���f*� "F�	�Ә�DCJ�q�n�c{4�_̏P�����v4z٧~������db�����W5'6hZ��Vǖ��.�; l,v^kZ��#���l�����zN��|r���7S�J�m��5r�4���d���T�8#S��������<�Ϊ.�`�m�fK��*;
�U~���Y�y�~^��'����")�e�-r�n�Y:;8�'��u>t�)0�l2�p� �L��͉.��o�'��2�g���{5k�ܝ��/�ɝW�^%�b�Go��]�#6D_�0T�)��2/���0���`Ͻ�$' ���"�^�������EC/�Y6�'���������_��՞,0�B@�
�ǟf'�U��I�wG�*%[��q����~@�;�7��ѐ���_6�<�-�&!���{i-㹵�en�;���H�{���//�Q!�̾�P�ß���s�kѦ3i������u������vQ~������e�Ç����kD�L�[o��է��
�W�}{��y�3�/�����s�2u�M�C�Z����;û[3�a����q�4m9]>�T8���z�g�
����VA�e��>7�\6�Pd��@�C����p]r7e�H��5p�A? �WM�H��2�Wb�;�&��6Q��Uq+�h����<�I�B{��%�����w�;�����|��5uM�rZ���j��$O�.ΠUx�p�[�����3�P��\��e�X�(��T��xV��:��ݱ՚�;��g.v�G9�����,���!�a��xe�Eȳ}��������q~#��s&+}"=�{6拟W
���У�'*Gg��}����.��)��e�H��ʟz��T�@�޸>�-L;˞�D�b�U�1b8N���^+{�Z�N�	����u:ˋ�5���Ì�m�H2	�
ܺ=:�̿-�'��=��+%f
�Z���2�)�����۪�[�#ܢ�}�ݪ[o�
�:��}3��ĈEl(�� �B$�e�ƟhwZ���^mw�v�q�a�0b����C凅<�v�1�\}h}�uF+�k���s=����}�=~���#J�E��64J�(l[���\yܾ����D�^��֫�ֶ~�����Ny୛��1�n�`�M�:V=Lɭ�ɠ%�1��!�?I
: �ޟ�#񍭰[�
��e{��o�R�m�Ld��nSV�'�x���/+N�[	E�
N>ba��=���ﱸs�V�?���g��'�xk�����Bv�T���!��g�0�f��q8ی{ ffӚ�i'@�h�A��{7\E� �z�{���{%���[%�R�I%8	ř�N㷵��s�L巵�lLΘe���;�!2a6�P��1qF[���=Z|��#�R��'#���c���Ƨ�{�,u�̯_
�Y"�5+>���G=�Oͨ?��g�#�Z��{ַ9���h�X��{+��힚s����
��\��؎��r�q�~͕�R�Ͼ_�~����.]�j��:c����"��� )�6@��`��T��(G�v�oz��Q��^��G2�#���R��Z����R�/5�G���,�S����m&yCY�3�5���p�	�3~�4�I$�2����\��>u�֥f�TAZ��q�x�e��n�2�7X�ۋ	kJ0��i��B��t�7yT�o�n�Џ�/=E���l��n���*��cGa�����f�*��w�tf��~_I#D���æ�>T��y<��|R�^U쭼�B�`�&�p��{�s����u\��Z�bF�m�և<�]�nײ�u��݀��\�B��T���O���ꯖ��n�E�>$�L��q��8�dN�3�`1OW-��p��F����/�E�tv{��T`�f��f��2��\�T��a�^\��y+v���`B(���Z���oY^�!���ڕ~P��5wD�wSl��F��͐������tlJ}tG�d�䥍����r���f�u��[���IRH��i��[����m�围����L�4Kv���#����p�i�ݲ�=��s��cI��ڴ�v�yx1��t��$n��Ќ�B�G�.YR���.�c�y�p֤b��0K���X&�Ty/m��/2��k
� �s{A��z��1�gKxM��YS6�
���s��R�hBʷ�gV�1fYL2�Yv���v�U�}�>w�ޔe\�&����(�������x�,|���D'�s�\�����"��$f%�%Z�N'�΋e��_^}YC�*s�x�0�0�~Mԣ6�g<f_��Y�ԯ��ϱ��W��`쌞�ΘR���έ���:�	</{��z�Z$R`��c��*.n�V̶����1K�
��<Z�$@����"X�]����8p�]��WDR�І�HI&Ci�]������j��t������x���)���^�O�xx��c�Ы����5���9�S{H���M�AG�����E�U�$�z������H��U_�Y����i��^��k�S�5��.��b�Dp�� ��=I��\>=3�a��Gy8`��d�3F/���G.]�F�"UU�`o�pC�T�d�B4p�g�h�	�`Ϧ�:�缢&X���p>ڿW�]�Y���5���s�g��36�'{�x52��F��G?�Dm��>wS���&=q���ޘ(����sϬ|DH�#�d�T�1ʆ���>�Vj�r�V�<�=>�����=>��� ���e �p[sh��7B9x��s_�uXB�
�Ng};��
��]f>�O��`��$hݿ�I\�3��fr4���>2�Y��;��|C�epb7kE��b:*KR�F�\9Zqq���t�0N��֦p�Nhyt��[��gii[Yo8�!]�S��a>W�V
�M��4E��	e����!{�:4K=,���T��9�e,�k�un^"�Jܰ�����[$n�+�dQ|x�M�}��܊�諐C�2�OM�J[�U���&mZ	�wf�BU�}�	�#g�iwF��XhR�{A$C|\{v����V�P��u�X�w2��U��[J�����[i���0ᖮ#��Pt9tɱ_te����!1��t�}��^L+�l�G.���dr�.w%�vںU�����ΉNM���_'�k=�~��������vS���uf�����5\*Nʾ��S 
f]���x���������;�D��?��#�նR	p���ZԌ��w`�n�|/�tVc�lgd%>z�gTf�n��O����
x�?��H�}Y���`w�3I�lP��y��mi���O�[�ʤ�e���0���^G���C�bG�Y1_D����l�+7bB���k��Y�+��n�b����D�79f l@��Y��j~|v�؎���^����W�4��_�pTյ�N�.0<����S�p�1��y'F�p�`U�ʥm.T f��,�ѕ�qEQnKΨ��L�w)<�W���楃�]�fq�v�5O��ky=��L��t��ڊqǍ�w��⬺̬*�rG���`��Tu�.d�P̬�(�\�umQ$�h�����]YD���T���S��B�5U�UJʁV�[]4�N�^��d5,��2[-��k��%/T6�KULЃ�F�B��0��An�2�V���ZG4�M�Y�8�W�����k�i�>���Y)�}Ce�%�c��W��-�Hv�z�k�Y����Jh�;�$��@�l�Q��\�vс���Z��W��bF����b8S�Ycmtd�[@�Y��ˬ����^�uJ��l31(E��W������ٝ4!3f�Z�����Ws��%�ҳюH#��;Y��-����pmx	y��f�zɜ-�%,�qnJ��0�P���+h�c]��X�7Y�t���&�� j�qGsv,�8ܮM�a���A�-�LGR�c��/!�Gc���͋-3�ȗWkd�%ʞ.ݺD���C�p���\�385��Ρ�=���-�1��v*�X5���m�k�)M�&l]��wH�xw	���+����s7c(�S�S\S�8䗶���.�lYy��.�aCPh���n������祥��]Mz�,����e2 q�ͺ;\����qɨ�QHl̐A%�x��Pj 8�rf�;g:ƛ�7f��h�������۳	�V4V9u�y:nH ����G�py�Z�;h3ic���,f,����m�m�:-;��#�:�M�;7�9zZ�w�7+[f6��M����!-q�����Ѯ��G6� i�n��u&�˵Hٮ�j�=;@������'@��Ev"^+
��˵�%*At"[��v�3v�4�Bm0��0�6a�Lf!A�@��+l�-bA$��m���"��h:����882�/�m'��ٍҬ6)�6. Q����d��pR:����X-\tzxn��ui3&�i����i�m�]�V�Gs�����!oX�m����.N�l�9p�sf�7d�=� ���uO3�����`�v��w���q�q�.Wz�M(���ڎk��L�	�s����*�w�T���B!`}�}��/��Ꮧ�;���M���u��&��e}5- � Jdx��v�y�?�}w[��V^+�K^����� ��t� �/!Ƿ<��q�.�\v�셫�GֻW%݊��7���7ǚv"H���#��$Oe����O�Q����(�,�=7���� >�<A z�������3���}�*��ZL�D�h�<������@�v򲀍i���� t��9�c����z�G�<���x����нڻn��>�A����o'�=����E�~c��+�!���QM��pY�]����XE�TNI\ C����F�9��8��CJ��Taf!��}�E�79g�Y���t���}�L� v�s��gｈ��#�:� Qd��v�g!�����T�_�����`�>�C�`���s�u�8���p�i(4<G��O���������|GÇg�V���{9x�4>'�p��t ;��gЌ?i�t�>�{;\ ����#���|,���#k��3��5|,��K�����>㗼��z�|V�D��"(A_/�@�	�{}��5τ?}Dw�����p��G﬏� 0�G����?P {���[���~d
 Y�? ��-�o e��7���?_{~��7z=H�����@2ӝ����m|��&�?C�۾|	s7W��͸�	���|�t���#���pM@Gᄑ���x��t�_NGF	'H��M��	�#�ͳ�r�䗤��A\�]��M����#r\m_.��?�}�\���A$����p�@Y��ᧄQ�r�s�x��H�/�����Ћ".T�ڮ|M�����E��Z i�
�!�5��u�������zh[/�7v|����:ݾx���ܤbش�(�	N�?��Ty\Bx	�����婎���t��;ω�}�C��Na*�p���l{>��K�|;W����'��<DtY��?G]c������T>���P��-_G�zz�R;�|�~�>���W�0�����A	k�w��YG�gBH�����x�#�Hx��7' ������P�r�Dz� C��.r�χ��*���Y�>*p��� C��kלּڀ�d�eR���Fqp��@���� s��>�>�������Rb$��c�>��6k��	*�W~^_y���GH��4;��]}�ﺰ�!&"I��'��������ˮ��Oi����C��h����]L!G�#rꁻ������ ^S'� Q��������t��������W�!�~������ó՜���W�0����P_}��¤6˼ʭG+�2>��t��� g	��4��|)���#�0��ڶO�0����W5}���~�}��sP?
#���_;tUHc���>�t7����L~�UY���_w��Ϧ�+���2"��x��G���с�Q2"HZ��#�6|~�+Vp��l����g����H�ȳ� a�>��żC9�Hj��#I	�&1���NZ��\�6=�- ؀Bi����dg��F/{}����}����:~~p���=w���|(2���~����<��hM]#޶Óg�WHd|�U$������=ܬ��rTp(��|㟾�����H� �D��JY?XWJ>�>�E�>���Dp��q�T�r���"#���?B>�3��n+vL��}uh���lҏ���\��\���	 e!�$��@�Os�|~\���	n(̑��������#�o�I��|�)ʱ�J۶O�nI�����wU�]�}u���X��n��R��[߭�8���~w���^���Ӝ}����|�b�'��Dh��$}�~��������r<D?B?i:F����8��ӗ|����}D�0<h������}�2��o,Yp��������W{�!�{��AaF�f)σ?�P�:@�wϾDG�~���~�.��wÈ�ywz��U��|���m���X� 2e�x��_Q?C�C�#�����p�� '��3z���p���_�K����p�e}��u�n��}�:@�_C����ө�G�9̟YC��~���.*^"��Y����(���������2Ĉ��?
{��&9�*�_��<�u,!k\F�Q��p��"S̺��z��$c�˰�|t�����I��������hMZ��M1rC.��5�f:h�B�G@�f\ۋ4���ڵ�evf�u%l.8�fK�"sۼ����@�!���a�j��?|+���@�r�?"���.9�\:�������K�e�G��o�c�{Y��pI�1�J�H�����#�Ha f�s�5X�~�`6���և� u򳂲?������@���L��u�>">8����hb4DT���]�W �{y��~�>��H�jw� WS���ʌDCQ
#�_����F�s*�Y]Y[? b�k��~�c᧤�W�6��D@Fs���������>d�3��d
����H@�>����t��r�] Ol����v"#`�,|:~"y'i����$�@T��q y��Y�E;�����p���_ ����}g�Y�hh�_N�Uc�ߩ���wS��%j�XLv���u�
�����'c�w�B�l��*�<�8nf?�1�/^
km<���#v�*�tSU<b9��Qظ#i����S;F�������\�ć[��3x��:(׷b��gn�]��m�rp��m�1�iaJb��9#%�8 �:���\.��]N +��\�����2
j@p\V����I��t���ۤ���g-p��`Km��1B<e6�q�k����bF��.�N�&�s�����z�.22�� B��"Q�T�H�t��1?�|��+w��$2c�>6c�z�PchV!����&�h�}>���2E�B �8�PG�;4��}d���� o�
��\!�����t�����L�E�����;Y����A}	rx��h�� PVoA|l�F��{�=<ë̚Rَ3�G�B"���"�n��r����i�\+��&D��?G|w��!�˚��!��C	il��=��q���N�t��1F�p� {��!�,���,����"�P���8C�}�8��v�X~�7�1�z_
@�l�	m�(�䛩qߪ�J�j�9sF P$Ѕ�.1�X�f��"��|:�$��/�a*�M�Ӆ�4b(}�ٷ�#*�=8�e�-r���-���(���N������$}��s��_0}���d�$���}��� e(��.]8�����2�����ɇU����B�k�9�z~d�I��D
x�I#ӊ��@�;�}��ph�s>dx�/��s������PCf]r���K����*�y�����z�H(���np���*��O!��В@{插�빽n�d� 3��/���=~�Ȥ?}1p֠�����A��D&8Lm���$|:��S[ˬ��>�5��'��g;���B�|4�z~W����������ӨQ�[��?yg˅Hw��/SO�U���LiZ����v�����y�S�����p"ԅl�8�?�h�wXb�Q���um��$��R�{���Z��G�1��_�Crx�`��qxRX�J�Ȣ>���4�{-���E<;|enr�ju��L�ۈ��!��E�l��h��g��p��c�'y��7�~y���f�����<Eb�a�w� I�W�<>��<#�>�g�x9�k1�"���1Dpν��7���e9ق2�������ڢOˌze/���Z�\ �(%�Z����[[p��҅<|~3`�<�d��F�����_F��7F|��H�*�m~�	`��@G�l"=�����y�D�A��'���, �g��n��Ë��SPx�K_L<R>���*���d��Z�ZP��y ]�w�������4},��$D������н�=�+
5����!L�#`�ys�:;�z��(�����#b ��9��]U�m|G��1#������"����V;x=fR��e���^����}��X���e�y�TD��cTǃ�U�"�/�{�!�YP�љ�xa��� Ǧns��� $f�o���<����������	��B0�C��s�}w<����FL\WY��d��!�þU�E�'x�ꙹ��PR!��$����� ������~�l�~����ϋ�!z�v�Z8] �ᚊ�q��ۣOR��+�=V;;Q��s��W��������I���?��pt��=�G�O�M����Z���b�j(�p��ս�G��ܦ�^�9������1sX��efh���.�w��иnK�_���Ke+M�'^v�]Ks��N�۱�iI���Yy�Kʗ	�T��z4m��h.K��$�4bp7 ��?pΠ���!����#��ڲ�}�wg}7y���SC�1�C���a�@� �ڛʚ?E�(Fa�$Fi�c�O��$p��k��S�L����4�(1 (�+�@g�/%���1��}��
��a�YH@�;6�Z�dc��"3�韠�s}1DO�~�����|`��WU�v_hY�7
���� �fe��V��9��Hs�,��`3���h��X�!H"��;�w�_7�ϣܭ�'7j���qp>�����|����h�����Ht����o��~Ե���nBT�����v�c~g��xk=YΧ��! @�(�� A0lhϮf���p��/��0}�i�Ȣ��,_�
�x˼δ60��ܜA�?ADu &�զs�/Vg=�7؜
(��>s�C�<��m�
�CX�Oo:3p�ή��@wC�cqn9�0�ִ���xv���qG�ۏff���@~m��o��۾]�G�_
?i�n>��=�D��#�ƅR�z�>�,����UXO�B�΄�W�*2�o&�O���k�����{�n/�}s����0����jZ��z��Q#)���R�[�U���z�w}Cc�^_d�t�>��/�9���1]��P���f
0����������ݼtQ��j�nC�$g5������c��;Y*5��'tEVf��78�K�U�z�\�;F��8�����ʾ�/����,��{~sw�$�=/0��|Q�KnxEGb��e����6���_v3���&���8{B��� sx׻�ϧ.��? `Rd���~f�]�N�^@x�Bώ<��;�<b����^Ǐ�b~b�޳�q�oj�y��!�}u^�P�w^^Y�̪c�^vEOUA\���7�������"%�����ML�S�̬��4w��u�yݿ���;7��ܝ��~��$8G����X���0E_�������m�&w�D��yyOu���5c�K4�O_��w�l!"�d� 1�.֟��K�ӛ|R�Om|�d{�e3�y��F���pd�5��W��g��;�+���^�y����uѸA����وc�W5�Tp�ɤ����<��s[�B'�p�^��mEj�mm�]׬eqw5�H���
	�D����X��v�9�WވY�g��t�!�!��` t��{<�}Ki��ل�n�p+�.��!�xz��T���s�~ ��OU�T�y�`0B#��I���s ����r��JzWF|^�Û���zQ��oyw�x�����گ��qnA�}1�v)D�>ʆ/J�����Đ>�R]~ɑ[xT%�ȂPd31�_�����${P�������v͊�q�Z�����L���y�s���݄�i�?�#;S�oU^�3�����oDX*���f��N;�EɎ眭mK����b꺣\ &J�n%s���T�w��[pƓ7n�<�5�#�hK�qX᦬������X�u*��mq�͡�З����C�fR�� �[9m�6ܖ�t��π�k]/ck;M�=�s�R�K�xwea,z�[�@%7����\u�X�]�`�C� �v��A�ޞ�v��\��ٹw6����HT�pZ�4!�i�E��M"p��Z\TWDGrm� s�i�[7�>�����^(���e=�ތ��	�H�Bxt� {=B���vq��"����48Vm�|�?p�f�fGѢT�!�M�������9�v��K�+�/v������ ��}������yy�*�]��7YUtXe/��ܠ�����,T={�U�ۯ6'���fN���0I��8�Δ��+lN��6��#�ɷ��J��͗��6�:����CV������}��~�����7\;�޻.��an�����ǘ.J�8T�&�$h���9�ɪ� P���<:+ͼ q����C�"��l6�f������n�չT��,xp��,G/OL���6��ƚ��%|һBȘ���<�G��0�gP�!",D��~N���९�v�'^竄?/6@�u��v�?v	t'�-�OM��]��:��-2
f4��J^<
���#5��<��i��q� z�zA?dd�յS��LW�8F� }b�_�8�֪9�2�5�d���A%�S�X��ڞ�n�p@�ѐ�%��U,<�<�	ϸ`�kT�����l�[4�f�X��r~�*����[�T��}O�l"��:/9�(^��ey�o"ह�<�W�����	�����\=�9�P�\�׊��QL������S.�f�T���ؽ�i��nqma�ؙ2���������!�3V����ų"�/M�1�.��tN�_Q0b�^d��BQ�ꗾ>>�J<c��Q�q�g�,u�Xn��70�Ԭ��7��@R��S�w7��;�x�O�{2+<c¤�޼k:fH:<͙�Q0z�	��q�tB&YѰ0�Q&P�#&%k��]|�ǝP���J����Ռ�4�H��5�վfl-Hs�����}��Uo��y��x�}"2q*�=�^{C>M��$_�Oe�_����ʘ�l����L��k����Lyw�Ǆ�����<Pso��q��O�_,��s!�n�+�DՋ������	�I6��E�OٺX��C�&T�#�*U��k��յ=��5[W�bw1����{��CN|5DǄ�V�岇����\��cs�|(QRB�6 ��]����i��y{2�E^s�������ю��0QVc��~�Á>��#�"��g�w:n+����Pt��S���spfz�3��1�T�a�Ḡ��?K���	�(��-\�Gi��c��?r�|F�xb�1�U�t�.����)��+-K��ڠ�I�"W�76Q�p����LK��b�������(J�N����D��/"o�}�V�~�% �+��h�*��*�P�v��#�T�n��}N����e�Y�o�}�"ۺ�c�=�z�ql��Y�]��ti����[�/7AY���n5J��D�P�d?�{2nVf�\R1c���z�N"�w�Q	�<}���R��3���T�H��b����zո���gz��݄�Z -�aQ��\�<��"ﳼ�w� �_J�������~�6??}nyT�s�%=�W����<%	�q�
J*��L� �ѨQM�bf`�h�!��{;��uL���y�wy}S��ޥtkv[)�s��|}48AM�{�����Jp�C�^����ٻ�aHe5h�|vfz �K��<�Nݎ�>���\�:����se�}�K���W��
��uS;�FE�oU�sO/ݑö转��+�!�*��mz'�w*��/���;�$L��iz
�	?�d�NN�ܻ�7<��9z�G�gkl��s>Xsj�ϛ������}���+�����:���b��p����@v��=���z��_�H�@�������(V��{ܳ�6�%���	UQ̫�2w�#%�n;&)���-��JH~@���n���>�|�I'I��N�I�ww���w�?��zt�wwx�y]�'wvwI'N�|�:wwI%;��:N����:I?�$�?çI't�c�wt�$�	�/����������t�/���������9����_����N����������$�'ww��t�t�������i?N�I��n����$�����_�����3	��'�OI,>�I�/�$��ӺI��d�;�N����:t�I�������I:N��~�=�����?�����t�t���_��~�?����'�����}ߔ�$�;�����~?oo������t�t���s��$�'ww�������I'I���3�z>$�'I�����%���#��6i���bi�I'I�������~���$�'ww������,����>�SY�I�ww|�7�~�� >���?*+��,~nP|+�ȯ���$�;��y��	>7��������:I:N����O/����]$��������������e5�9ӗ`(�� ?�s�m����%�� ����
C�lS������4 �[]�.3@� ��   ;��Lz =��     4i���p���@  d 5@ �P:+!٭����t }=     �      �  (  8             �  F:���    ����nm�=.���a��돣��u�}y�W���t��_A����5��(
W���ۑ�ǖ�=o��{�O����s֕�o�8����ֽ���ՎU����ݝ���v{4�����[`p,	����G��#M^�A��^�}A@�<������P���:
���� P�������k}׼uTho�v�Yu����u����͵�u����kܣӼ��]t�v�Z�n�ҽ= �Xnk��*^��a�ש ��֏]tj�����4�� (
��ӧ�ю�T��u�mѭ�.a�]*����%^���i��O!�ôǏ�=�ﶯ`h�c�k�ET����8w0�6z��{�����o]�ʼ<	�S���X(�: z�h   v�{�5OM5�����-�P�����h��S���=���������5�ݛ[F�0W���"W�.Ŧ4m^��ϣ�| }m������'���=���{�ݳ�\Lz tv��ֵr����S�s����M�=�z�{���o����Z���'�=og�ürn�m�K�OF��]���������f�\{aplw��*�^PzʶY�w<��7�v�d q�o���L�Ւ��. ̫l��a�������{C^�w��)�y�u�vz�znۻm��T<.�ٽ5{op�ۮ�GVޜU��*=ۛxr�3�{w=���=  Fyݺ�5q�{���B���v����^�V�g�K�j��s:��<���w��*�wz�y,ù���AK���onS�;����̌e���R��=�  z w�_w��Ei�9'ox�^9�i9���]��X4Vͻ��t���N�x�i;zq={��ݹ��ޕ�4�����^ְ��y�5 (̀  X4m���#p.R�{�:���t.ƃ�A9R��9ۡ���y��x:h�����s�2(��8@=Ӷq�ivz=����3�h�U  ���<�  �׎�>�j%�gx{�(�CN�ا��AÃh;���%������(]��`vʸcMj�4�pl�zzu��ݽ�w����f�s�o���=� 8b@O�*�4h� 4�ɣ��$��Dh�� 44	RM4�e6�F��OB� ��*I�R� i�` 0�? i5U(� 2h4 �$�"Uh�@ @}�/��]��~ߴE\�A��8���}�LD�)wS^L�\����B0:0 !Xp`�r�� �BK�p���	$!$�Q��B@	!@ ���BII(���������HII�+��@�BO_Y
�$�$��͸?�I��B@?ʑHT �준c$�$��	+J��� X*B�$��@�@5�*@���T�Y$��%`H�bBa!*�$�!�$@���$�� *B@X�c��! cH�$a!%B ��HT$��$�XBC���`�d����ĒcT`T+ k*bHbT!R�eddf0++�$�R���HJ��VV* B���1�V�J��V�*�T?�f$�bI	�I$� �I$R$�T �$���T��&!	5j MH@���@�Y	X@	�!$��&�IP�c *��IY ����ŀb�	O1�//�C����/�i����+/�Is$���P �����rIK
@G�����om\�yu�4/�{gJ����m�}*��j��)��$�I{�iE%���e,E���N��3��B��<	��D��rjg�u�Blÿ���*egu����q�)Q�?\2k��m֦P�#��(LU����J��Z�M` �l�6�x��D��ѰhV�Z�oi�b���dE	���\�kĪ�>쥓�k\�*�|�kH.Ow�u9���˟p��fv�SHV��h�FE��_�>&a��6"�(�N伩����2��>�J⬷��KE\�X,�ӌ�	�v��^�m����)�so	�n�,w{jU݋�
�r�jU3�����c�7n�]��$��R՘��jֱjռ�D�Y�p��9{pLҳ�����߱�7�M1TP�f*%4��JtUʬr�P*"e<��8T��`0����T��&��%�L�,��U��Ks/�"�jkr��ӡ3S�@�,D�f��w�yD�%�|�ܒ��ؗ[dlt�Y�#d�>VB�6U�Ya+�BaF�a�i	�>6j�>�
��|F}��"�o��:����fX��P�&]�ݫ���D���{Wq)�d�O5��x"��ubN����L�ⷴ$X�P�ڊ� R�ݝ�/`��eX��d�צ��c�d�U�P���Q9�Q�Q�'�b�SdS84f���VSa��2�lW�[�*�3>ә�v�^$C�vb^�XI/)b�Iye��f-��Ś5��@L�Д�/6h��d���72�U��f(�ۺ�4�E�3j�R���3/E�N�jޢ�k�]�U+�d�-(&01��0�d�(Pfa�q1X(#!&��?�Ց���iX�բ�^C�F���fGo5���d!�X�q!�m�z/0� i0rB�QS`��aNeRl,Tt��Q�b��%�3`�mM�,��7G�ŷ �*m�k~�D��ԟd:U�o��bT�P�v���4�l�/�&�S��
5� ����`e�����j!N�4���ʼn�cхt�G3e�t�df	+lEcE`�s�����~7QI�ۄhkHp}�!0͌���J�9	L<'1�㉖-�J�:f�1�P��9TY��p�]�����}�0��G��'������3,8e٘`\��]8�����R�N�A�rn�m��SH��yvr�ӕ�֡s2,�D����	���H/Y*�%�[��tl^�Zu�32*��
@ ��)n��i�f��	{�FL���7r�[��#r^�nF�Vɲ���ێ`7t��#ӫ;!gfݓ�n�e���D��-ǫa*��]���2��S5��be�B����3x�B޷��c���靶M:��~zvw��O;v�j[��H+H
%9�s�ǥ��.j���9[�����Z�%����]E��YL<Hm#.�*G3/"v7ib��hh��a�r�1X�kE�ր�/pf
�)ٳk[p�O ��+���[hn�1-:E����'�U�*��Խ� n��	�*�Yf�la���3횩�;�v"�fo=l���������а�e��r׀#��QY�ct]=߶�l�m���q^�cx����T�R��X����$�V��t�+,��t0T�ӻ+-ޛKr w�m
[�kF�E^])hK��K�e��uxb�ǉ�x�6�]f+�7(X
ml�z^С1ۃ)Lr�w0�R�Թ0��?0��Jr0���`)��u�UʱL��J^ڼ��r� :�(�Б�ߓ�U���y���l���vց��ws� ��j�S�2J��Qe�"��	������)�)�ʽɛ��輷Cst��%�b5�:�0S;u�!��Qq�QVէM`��F�n���[E�N������;�Q��xr���&����5{��8�2n�X�xqB��f�.��U�� ���������>�+��G1fء�ݣo�w�ܰ�3i��Զ:0^}nḇ��Y�2��Z��]��Ѵ����S�ζ��W�m�Ҿ�Uq!�Hq!�!�Hkz�kć����!Ԑ�ԇ�Hy������b�f�A�W�� ��+��tХ���c9��k|���*t�1j�N4�}�Og|�Q�d��_o��qa;2vgw NR��{�4����0*�6��y�6\@7.�KҪ���S���x(�Su�y�����Vj܍�L!�^�9z!�5U^��S�y�j�f`�s��ܺ�W���T�`ZoI��ER��36iw��@�i5�Q'H���<�/�|�:��s�鼾ud1��2Vm�X
cm�Rs9�^�;���@Q�n�%���Ѷ�7�Uݛ/~�Z"`A��*��˿G�f�f�xX�
�MM!uz�x����W����z����@e��˸��5ZF ��w���:��R�	�dvC����΢3��,�R��+1]L
̬�y`�G�k�k�)�,��6�W�𷈬pǗ�t��d<J�p��ܴB#��_a>���*P饍7N���~z��&b��²f�ҕ����Bȩ�#Kv�-n�^oI�R�	��Eg	;u�%t�wr��(��.ᖢbԵ�@ʘ�NQH����C�7,!���(�l��`q����V("N�`�����(���率�6�����\D�B�Z4U�e3���h���*=64�o E)��h�ş6)U��jAȱ��D�X�Z����,C����*�'fV��c"kw���N�l��_ʷT�4M7D�W�hh*o,�8�=��֯]�k�en�PS]h����@���[��h�rL�K,��T(��Ŷ�/PLYE�$imQ��3^]ԭ0��{��QEzoEf����M\�ǵ���6��h�iX�t���r��]�wf�Vą��j��G�ݺ��k��%9t�m�-S�. n��~��&LT�OFM!�'j���6�\l�����њE��0m��6m�U�͕hwV�BvC󴛊�\��:�̺n�-m�0�2�v�K�b�>72�dZ�^K�$�YW�t	�+M����W�J�*e^(�P�0���tv�T\;��
����w�(�ىnZ�՚��l6��ՁjM�s"�=wut�h�oB����P^a�]�Z�K�f����/V�Z�&����^n�f[30�QJ[5����F^г]3#ƯnI1���u����K3�%�Ō�H���7��o%Pe�X�e�WV��T��T���9{�rd�}��z<ꖷH*��c���Z����h����V�3곤`�L��	���ܚ�n1�r_��Q�O=��c���v��mȰ=r#�@�a~�(�0^U�f�VE�8�e���W�e�/5�r���&���V�
�"i��A�Wx�Ţ����f�@�����,M,hu��d~������v{�z��u���0=x���ƱG�8����Ԛ�2X�jC������f@RPE�2�I;�u���p}�C�>��ŘjZv��kLb7#*��5kX����i*�˱���eʚ�O�z��w�W�����l�P$8�XB�,�0��A�t���^�l*���0K����5f�Vp�y�$f�#Fn;bhH\W63���+V>ۺ�Џʅm;�m
Xҫ;k`�~��:�t�Z��9�
Jv��׮����Cs3�7kP"��`�ɳN��F�҄-�Yh��w`�����D��&�F�D��n�Ft
6b�-OB6��Rx쫥w3r�5����S\�7[�6�[,�[���*��Mڱqۺ�ũ�3�d����i���ذ�6�P�i��5�me�n�͍ԣrnܫ̖�G�ڭ�<dͣLd��p���"���\U������mL�X�������)�cӁ
��b���o^��c$WK��8��V_ژ�Y"�^�W����4hP�𫷶U`�QU��m\����aA��6�5�Q�Vlj#dsh��^-B�K��(��
X�7CL"�op�AT���Ҫ̋H�ʫR��*�A�P�>(�ZL*�F��r�Y_nds.k��d��`u�5Z݂���a-lū,�v(J��鹗bs0��(�v���ADZ�)X{GM��s\V���z,��㪵��ףq�ۄ"��QV�֎L���,���#T1J��Plj�bj��pdT(*j�\4�][��Z��;���I{�=d�b#�X*,X�-��J�2�X�edYb��$DA`ԅR��
�aP�-II �Q ��A�1t���r�T�)j�f���.$�ST�t��ut�{sq()�IĤ���*��A~
�n�v�75f<�!)��`�~>+���Lzu��Ւl�1-we[i��f-o6��m�j
	�ڵe��Q���(n��1-յ�Y���9���t�ZGm2.j�Z�@��YWU^rM�J��`A�Mʸ�ℕj�	�p!�����q�����[�wLCK)�NZ�6���4oi]I@+�w�T�Qys7�^yw��/��9�;�J*2z��5��H��UDAY&�9A�[���P�ӂ�6�l�`���|�2���g:����{Cd�g`��!Te�x2�[���6����w��f��C� ���5�X
a�Cz�<��g��F> �)�Y�]�4!�/r�C^G �C����)�G$}��zEmA��˚3���[Gm�hn���%f�Yxa�/�C�T�^z�Tf�i��q��-��ͅd:�t��,͗�^�86���[ô�j�
�B�ɮ=��`�[f��3�q�q��n���mMءAx��&��;��8,��]��/]m�Rڏ
� �� �M@�S�Em軛�Ja���.Q�{y7,�V������҆��Y7;i��J�q��G%�����.�*�zL.h�+Ev�+���4;U�@���ڹ��;�Jc�[Z�F�I����zkn��NO֠�f���hڳ��H�T�f�M
a��տ!!H06eC��h����v���"�K�9I��UE�M+pE�_�È�rpe�2pVo�V=��{Hm��x�U��m���
q�j)F�v��ʓ4f�*��W�ll��eJ�[���J�"�m@*$9�-�'Kg�8*�*�	Th�����\����%EH3-C�$�EH^����i`�V�K"�&,�i��T�!ųLQөbf�T�V~2ع��+��v={q\��~��mb��T��>�eՈ$6�7X̻�"+sjr��q�Wy���Va()�%�{�m�K�Ī;�U���ȼ��#v���ڽ��iml|�s aV���Nc�hŦ�w7M(��[�-ՃA�Y�k&=b��7[6="�XA;{BkӷY!7��2a�˩swI8�T9��Z����\�9wr�ee�U��)�y���J�o�KTӢeKW ��s&n1n�Ռ;j.�̭�cRj�Z��h!1��+(�m�fR�^c�*��v�`a�ʞ�G	�Z�n�Ţ`��:Iխ�^��Z�8T?k��0nEY.�a�$��+R�qk��-8v��,Cb��͛0#��y�C���h|˲n�2�K4����%�Y�[*B
�,��7�.������UM�4,�a�2�Ԓ�Ż��qȨ��l%&a;��eZ��Y֣����m�]�ә��$bpf�.i��	�vɭ����u�\�.��v�s$�hU�f����ۈV��~n��
�'`�&X���ǵ�����;����kڶ��`�Yz��Ү���Yلa�no&��k�%���O�6,B��	Xf��j�+V�p- Y�{�3�Pj��0�4�۬�ʥ���%٦ҙ����4ðQ䶠���7c�F&��N+wW��^5DV�u�J�훽!�_+��0�Q��{z.d�w.����%ߥ�wi���O��L>��[�WJ��`C�IG��㰊#(ُ&��Y6����Y��$Y��Y�R��[�/Mdz�v�CJ��43v�V�ƴx�7f�5yE� �o`{{Y��J`+5e�(�K4ܳ���EP�0�;�X�C��;F�����ݹ��7Ȫc��<®��B�f��*�h��vLE�.���Q�����0iP�P�͂��YP;; -ଓN�T�"�J�S�1�`*yq�]���1�*x�bu+aC�ֵ{1���I���zѹ�~��!7W��(f�:a+00�ȴ�E�1$P�����a�Q��G uLl��E��][!��2�8�sv�U�RwC��G#ٷd&{KKN�p��3^���"���2�Ԁ���R�ܥa0d�T���ź���.�b���vI[��o°4A���]��5TKf#"�D���B��6,+�TȘ���F�i]���*�yj,˲n�ͺ(���(˷��Xd-k�J��н	{���6�֋�6�*ܩ��v�3�/��yl��W:�boQy��B�2�0�d�щ�AA�Bb�;Ě 8�P�$�	�'w$����>�˾K���s���'����FQ�𪪫�UUUU�M1��������*�����ZJ�\*����b� �40�6P�j������������<�Y�nn��pq�x��e�gA����m�w���c�̾ίw������jj�%^��X0�X�.ڣ7e�2��-e��z�6��� "�Y����O��Jw�$�9bi���Fbm9�n��Pr�sZ���(��[�����;Y�s�uo{y�A��d���[5Q�g#V�R�L���8L� %�WՏc+T�
DR�l"��V�?Zu�3������ZZv�YÂ�Ζժs���c�e6��:fV3��U��ݝTW�j�f��Wq{V��Ĥ*�D	���ڰ'�b�&�I�סY����b_��
Yu$��sEҷ��)�i�ٔ�mg	Im��:��T*���f�f�&țۀ�y+�/��N�Z�ǯ/l�82�س�0���9��p�Ю���n��;R��֫���\��v[1��1v��Έ��v]�� �of2�B��aa�4��*���F��5�XX��/pd:��v8̭Sj����;TXz�{pnY���Y��"_
X�KA��!� ����9���U���Hu��][�y2�m���v<|)��������1H�l����yۗƭ\��)��51��;V�t���\uj��s2��c�V*P-cy���0s�1d��]�Bk�t�%87����J*̜�Z�+ur0��z�9sW��k=�y
�s:�r�Lv�&tT�Z�(s�Ƒ�f�'t�79���_��Ӿ@퇳�_�K��u��2魩h
5�ft�Բ�꽏6S��dC��E}�Q�D����Iu��m�v�ï�2,+�Ҳr�[�t^��
����: �O���)�헇s�ٮb�|���&D�J*�V�4jv*���aЂ4�Y��ĠN��2&�����SQR\����Di�-���[	��l�Ý�`BYX�K[�]�3	#,ֹ!����46V��H�x��v|4,��L��r^�
��ٴ!}�1V��k͕t�fTE�IӔ�y<�;}ojΜ��W�j�a�
�3Aĸ:�YܮЂ��9�5^�N��<�iy�p�˞R}ZM���sy����#�x#����B��G�;�Qe���g��z�и���3gu�|�Z/+�[+�<�⫹5+��FGד;fλg^f�iQ�W��m�Y ܖ�,R��Ü�j٬����4p\�Y�>cg�1A����v��K�7��v�@�`��X��X�&G����A�L�8 E�r�,�tL��$�wיK.�KǗ���f �r���W)'�Z�Q�*�tt�.v/Lc�_)f�A+:�����<i8]q��S�Vj�D��_ۨ���wq�d��u�+��N�䭽�Ts��}S��JhQ��.�J���nz�nG��D1KW8�λVccD��13��E�ۮ�쓪^�a��.�Z�a��
�n^\W\,Ϫ�u��ԋFR�Vp�7N�k3,�xb��ԬT�ݵ��CK�vE]�M^ob^ؘj���7�b��{�v�]��r�h=W��i���U�Y6�'�ԏ�(mb�:���mhP�y��*5�"2�һ��ohU���i5y-�f���b��7��.W.�t-�����k�9m��*˾��}6ዳ�.ͼά��:�y��O��RW	LM׬��)���@ɟ�kT0@apC��^␣Q������ˁ"�n��m���=(�(�V3�ӷL�B�	i�U���\�Y�]�A�����6Ŝ0D)v��CYS.z�i2I�(K�Z��p��e�q�{Yx�S�Z��z�\@m����m�`�ݾa�j������0l�ˌ@@��]��,���u�s�`KR*'d�+�w��+d����*bɕ�T���y�_��{IDQk���^���,��]7d6�Sr$e2��Dĩ%��Uzh�����sz�Y5�mk:hn4z�};�
I�M�'��ˬ�]C �;�5R��9|Ggn�քT;��A6�u����/�D{y@oB�O/xU�VŸ�p��7I�42(W��6Jp�l �#3l��::,Q��n����a��/S��M�u�{��Om�H���H5*9,�5tB�אn;��ǩ
�v(uȯ	Ǜ˴��;+��J��f|��X����H95�y�� �_u�3����
<�Ya-y���ӡ���OBź��W��2k�r�T��Q֐"ŹXs3�Z�N�D��4�͈q.���h*EZ�a�B&�Uok��>��z-��b��ǚ(*�m�:�����멃�7����)����	�_i�r�(ؽ#Y�U��2��F���D#a���թ�7ȴn��ի�9�e ^�D2��t��P�Xĩ�?�!w����i�u6ۘ2��ʾ�z�̧.�����R��*7���$8ot˛x(��U���$v�>'
��@U���7y����(�.䔵z��Ȉ[�
V3b�f���Ņ0 ��9ݪ�j"
Ȅ�O2,q��Dc�
��i�j�s3�"h�$SV�!���8
%e�k5	���0�����O�SE�!�Ói*+���`}�j��wEz[��T��ߜJ��V?�0�!G�)�R��劷�D�0EN� �	1j����[�ԗ��2�cl��P��H2P!Ji�9��L@AM�g	�?M��_>��<6��Y|<_���%��hxXy�ifN�~�����7����v��>�yz]����p�}�"�;���{����	�����|�'-Q���?P��&@�C�d�HЀ8˚�JKPʆ\@d��a"�-�o��tm��J�����	����tE���f�J��=��o�Է�*J0%$X%���ET%uS"q!
��P�ay����滯l�+��e���wd��%��Y�^�1a�a��:��ڛm���j�zf=�:��ä��Q�b�Ͼy�y�����-�Kn�t����ӧ�������Nۯf�x9�B�f�����k�ڽ��t��ޖ�� ��"��x�Y���Kg��t5��w��v��ؘ�X(U3�H�@0�Q
Z��'ZܸZ1���4:�>�ua�5�f�Mh��T�jn�ȅ`��}I�ݧۼ�V�p�����7ħd��Kkit�{f&��%ܬF�ˣ�a&����w�ˎ���W���ݡ	n�j_z9�]��m���@řh���qG�Ҳ�.
K}�7���(wX�Tfܿ.���[Ĳ��{�M���)����c;�m
d�vذ��I�f��Yf�ң,%ɮj�lƎ�b�dMg�Xk��v��l��{��{zA�@�����7V(�B4\!JLi]jl��/m��ZLc�%D�RͅV�|���\��^���@	h�����8g]�+�Gp�֍�4#yXA�b��~y7�_,��a���0JX0u��f}�/[qu�on�)[��%7�j�,� ��l�.�r&ˍ�F�Nm#un�|�,����^�n�i	�t��k�ځ{���s�U �E���)���ר�xatF��U;�f�Y*ڱm����f �,�Ѓo�5�崶���!
�#Ynh�qL�fxW���ջ-��ls�1#-:���@�L��V��V�グ�+�+�jP8mi�K%��vx��2kGCM ��V�u�hM�H��[7��f�jb�؀��V���͘�β��S*]����'y����&��٫�}��I��8YD��u�����hL<Һ�]��4b8ii2L��hk�B�g��o]Mˁ�ԕb��[F�d"B�u�̲��c��(���,�-�m�v��)Dʠ�1�FV6<���\��2�_��t��XM��Ёm��c\��!�(#�k�Y��^�xKFW��N�:6�o�]�&��ܷ��l۸���q�nC3&�_]M�t���K����pϏa�ێ�qXl��4*�k���ga�6�ƺ���:3M��������,xq��j���U]�1@�l�lM5Hb�^�F�v"�l�51�٬�i�\ۮtau�[��o/)�d�6��l�>�����u�ɒ���,R�Il���Rw]�����ƭ6 ����3h�٘��+f�S�a+l��������K.�n"Q�i�A�i�(����6`�hL�WF�C⛶uЩ���u��|�R�֑i.i��[yv��L2���YN��Z?F��u��ml�a24t��4�km�.f14���ݯgH���I�^�vO�f��c�3S6�i�n\�[����: �vw��)#2
�\��f�nĚ��Te؍�(V��R,nH��Z�x�SE���.����V��Y��	-��n�f��Ԛ�M.p�tZO{�Ҕ�6�S�il!��,Ch�mR���K���ܸLKtx%�v�\ɠ[55m�u��<��Yn� 283!Z��B����VU��n��@�w�^��*n�D�P����E��¯1I��`!�;Mt%�3V��u4����d��.�M���ԥ�4���M	V_�3���L�)am0�`��е��"���),б��*��qMh%��cZԘtu0�YZW::�[��04���n�:ܵ�Y�`��,�[If�i��d�M�cf��"\ˬ9B��%њ�y�&�4b��[
FL��vک����\YC`m����b��y�x�4�k)��\��,SRǎfv�J�#
L��mF��&�y�-K�`�b�Me1�(V��@#p�Wm���],(%G:�[�LD��	�]+LP�p���5kh�jk�.��fl4�%m��]��qx.�وb�-�K�5�	�lѬ�ue��6�������E�]m�MX�B�07qc ]Ͱ��ĳQ5s�Z��qtw(60��hU��Rks�lɩ�hie4�.�(5t��R\L�]L�X�m�����vc����]��3	�[tY6����lLݵ�P�����2Y6Œ�,5�X`+n5��u��m�ƍ��\Z��4�
V�	����s��hÕr娭"���Iv���6�Ka8���p�k���륉
&��flA������02�(�.K`��)5���^g�Y\�)f41,,l��r��Z�c[bm@�q,�v8!�^V���J�C,�5�إhk��GV[BK�3��"��(FYx���:���[
�Z̪�[f����Zŀт��xh�:7ji�M)pA�喷Y��J�Z+�Itʊ���������������������������������������������������������������������K#y┩�݃�`����&@U�yb9Yk<�n��nCu�����vn[�
��We�"�{����	���;����T7��^R�u����ZH��G]����lP� �b����bɩu��K�,�o+c|K��L��*hf`s��1j��)���,5x�VѬ��a$˳��OX��Mv���y}�A�ӝwVmt�r�+B��补�W�;�\�P�{�x
�X=�������ry��dW�S9���2R5�adXm�/��ËoxkYv-J�[�1�5�u�w�ԩo��KX� j�6��v\���n�	E�yˇTy�r�^>���+H�\]�TQn��j�kYZ���pk8��v�c.�����՝���J�{k�@D��|���J�N��|���}ӷj����X��enX�.Ι���ˌ��gO;�9Ňnc;[���V�lS��h[��-�.����� ����	@�9����ĳ�8�,�$����w����̽��ۺ����r�R^��޽7��T����mp�|p��/�E��In�]�u��3�͉��͹C�:�YoGU����X�{I[��;z��4��+��k�ub� ��4-A�ō,p&���3h�2���^
�\�ͽ��d�T�W�1������:�!Z��r�N�Mks��۫�]e��v�9��y��U`�0�S���*���n���
�o@���Y�n�&��Ň��G���8gi�飴=�8-�t�+feQN�u7���)XL�z���K��p`�oV�cHJ�V����~�h
J4`��au��gu��T�S���������.�#��wf��g$:��xmM��+Q	�/ul˓o�;E�&3�R�4?���tI�7�D2���pI��ݚ@ӻn�Q�-+7��Zr<쮅>�b`Ѫ����M��w�C�l��z��%����h-��>�Ϸ����! ���� ����&���@�:�!	!Ԅ$����Y!�	��!���HN$��=@�2H�k u$�H��@+%BI�!1 )T5���RJ�R�	�O�O�f2R��'�"��IP�xȾr��� �``�1�3X�}�'�`G� z��Y&�0g�Xyl��PS�|��}�1#톰���g<0]{�Y�;�Ę��UAT��$�����:�����'�ԇm���PXy�@P��>a�8�I'��+ ��g�:�'b VjT�`T�QI=HbO
���<I�zŀg���2C��*O�>O�n��c!<IXCc �5"�LI��&=�Y*u1:Xu�!<ef�M@���R\f z�:��~�Bx�Ǩx���k!X8���f2HO�BE�dԐ�R
����5�ש0��j$����2�OS��فE!�Lq�}���]�k���jI���%� ���
�Y!��q���q�a]LV0�k�@�J�T5���2N��ĕ��O�I��Ì�묶�c'\I�'P��"��$�s�RkԜI�i��O�{IX�>�<aS��`VJ��k��z�퓌&0���:��<C�y����=�IY9�L尝g<�JȳP���1��z��I��`0�$�J�5V)l'Y��p��'��
� _��a�ݠh$�$�k'����;������& bAz�=Hj������8�>a�����R1��2�ĂȺ�y߲Iԋ_�YLdI
�d
�3)T�'��;��8��9�L�:�ed8�QI��$�:�T��ć�$�P8�����@с���f2E |�	�$�I$��x�d�$Ԓx����QC�+<`�BN!.Y%@Xx�X)I�c=BN0+'��X���BT$�BE>d蓬�5��$�_Y|�XN� �&2c+'�9I:��O�O�jx��(�����Y	�Y!���@+YFI��	:���N��@~��*���	�:���RI�Ad�$�>@P��~��z�� >Bu��Hu�0%@/l��I1�z��d<���IR|�)Ԟ��OP�x��'P�H}� ��OP�7�|��,	Ę�$�'���j�@�8���2j����Xr��Ĭ��MBcz�u�!*(3ĕv��u
�� y����� Y���!:�C���l<E���+&�$8���夂�%`�J�5	Xo� ��
CPA`�߬��`�H[f��E��O��P5�bLCZ��B|�P
�q1�9a�9��Y:��C� ����A`(|�x񚄝�傒�m b�c���'9}a�7�&}HVzϐS�u|��ʀu�=Cd3��P;i%�!�Lg�Y<x��17��3v��2b�,}��e�8�βc>~gP�$�N��=HO���,����ϰ���|�,g�XJԅa�'���m�V���OU2���O9@�$P�CԊ@����g��ɮ�p��Xΰ1	��_��֓���]`T��I�^r���u�'��_:��|�w�G��Bz��a�!�9��(q��Bq����g('r�<��:�=O\�d5>OX|��y�VI�'+
�5��;l��n��6,QE�m�7�7�$�d8���f�PO���(q�Xs7g�x�IX�3�'6̭"�P�I�'�S�3����}��r�`�9f2x���;u*3�P紜Lg�zϙ�a��䓯ɼ���vMO9C�|�����&��^{d}�*0����� ��ݽg>��.ew�=z��f>�����g'��g�����P�:e���0f=Vc#��Ru���}@�����X�{�8��M}婌�Yĝ��w~��f 򞎞�]=ry���/��|�QjE���ǉo�9����ɯY�-�}�7hz��=g�
�x[�)T�s߲MƬ�C����{���j#�3R�`x��GċU�C�g��L�8�	�q��bu�ēRu;}��+�1�<d�,֡�P����Ԟ2OO,Y�?}�yOP/��Ƥ�m�k��>�J��*����=�����:�ϐ���~�g��{���s��S����R0P�U@�P�I��+�[Yݸ���ψ�jT���u���:��6�ϯSm8���B��x�>�@���ۦ��bOa�w���l
q�u�d1qZ����$	D9-.��:��:�'���A���yE�g�P�|v�r?3�<d���s�C�4C=�ߪ�ٶ�y�:�s<x�_�ݲ��1���紽ܗ�a�Ԙ�|E+|�12V���i�;��I��͟!�E>@���3p!�u�|����ݤyC�C�qR�N����!�K>��l<�2<�%�LO>�!�-�3G�<��p��^�CP��8�<a����ęhju8'G�Ԇ�;� e���0��M`x��Ng�$Y{�'�(�O�!Ƅ1!�*�`q�T�.Y��d�70�0�l>Bx�ߩ��	S��Y댨�q���}N�5���+�����8�05�j�Hqs�c=a�{i&$�>@�C���]�͠jC�$�Ro}�|�=�"2�@��Rg��;�/^܇k����\�>7|`F�xӐV�u�\S�ӌ�{���� ��37�����'��_���  >�G����̣2`}�� �?��}b������X�j'e\Lȇ�v,�m�@r�λ �T��)V��tf�MȆ`QsGfVV-���xu	E
��,�q:W݋ue��gt�DC���&�R�� P��Nb`�n��������Sw�����.t�{�wR�.�r�	���b@I��.j�kڜ�
�WT�g��q���X�:�q,��X��[��K�7�� �7)���c��2W���B���=z���x�8l��SpheƆ:�|dt0w%��]j*e�!ۮۖ����
j�s�,RIRϜܑ�/<�fS��L�x[m\5��7"�+;凨��g��N�s,Q��6�\��:
Z�n��n������ H� @��)  ���)�@�;Æ=�є2��=sk]!���jêK[�m��^�ޙ��y���s�?�$ā ��a1��,$���!S���B�T��"�<�	8����Aa!���R�5$�d�q��I"����CY Y$�f2|0�RjRc*I���ȰP�w�;��������ϡ�Qb���b�"���b�V���Q_�7�F	�X��*���0UT�X�
(�Q��2
�ͥ���뀱�֯��ȧ9�o~�(�OAE�<B�����6�b�j"�:���-r��u,Tm��UQF1j6��Ҩ�����9ث�Ug�b�� ��ᨱ�T8�p�b�,WYQAX���QbG*�2Tq�b��Xň��_ݸ�� �o���c�9���N!UQ�TF�*1,�Q`��2+Ju�p����7��>~Ͼs��+b�Ń�e�YG�DX���KU��F*��E#R��}��^y�*�,6�mDI�~�QE�UFҠ��8�EWm��j���**����˒�s�Ȭ�ұO);ݓ�����X���Pb+���*/y���DN��R�,K�1s{�1E{s}���w3J~O_Yv��l�<��5���:ݣ��m�QF*���/�be�xب����7�������hň �Q�hS��8���b��v�Du�
p���~�t��q8X����E)`���>!��Ԣ��S�<a�J���.DE�R���iQe�M��o��jD��Z�J� `�aP�9I�n E*x|��Хj��̽��5P{�1k/����-�Q���pY�Xcc;���" ;8�l�ls��ߍ�7;z-�����˦mcf�2�֢���5�s1Q7��k���V[F�1k̹h	����LK�c"�HA �7E\���M��[L�X�˽�-���U�-q�?yo��q��2�ݷ7<l�b0�)����e��DT�S{�9���(*���m�yC�f:����m���Z��ݦ�ǛVFҦ���нJ�[�oY�6�(p�
�p�@ɼ%�� ��(
��K�>�Ϸ.nf��C�Q"�W0���u����(�5;̛�Κ����'���w4Eu���G�ͅkw���{�e�f��A�ֺr�R����QOs1^}�Ͽs8�z��m��h�F�QS��&^ِ�eEZ����1��|7��_pإ�}��t�ˡ����^������L�@����
��/�!�?T���2��lE��0��U�������|�+<�����J,-ȟ�~a0}�� � �Y1_��aA^����m u <��3d�E%�*I�M���EmG�f�b7�c˺PO�a�J<�`nK�1O`o����w4��B ƨ����@�ۈaR�'��ܟSgOt��?���Ji�Z6���0��/[R�谠���ԢA������L �RQ�=��{ǉu�/9"]ڑ�v��w=��3e�-��HFCQ�RlZ��0,r��8%4�x�,5���~E�X�S~c�7��+��X��.�뻸FlԛxU�;���k�,��9{�[k�Ƀ����l�lM�u����ऻ�'�RS���#5��u/JD�t�/+˞j:�A����N�t�Pj�S����uɌ�Ic�*���~����x�>r�D{�.p��}��c�G�-�2�[T�v��V��M�����{ڹ Y�HI����Xn��a)7��E ����#
���̋G��&L@����$��cO��}��>k����,m�û�~���.��n�����/m��vLO��]��1<g�S-�w<�7��θ���܎P�.��cx�7+QQ������{��b���VT�>��u����+�P��Y��fC�)_R6v��^�bko2b��iDʛ��ᔤ:������&���"��"PU����.~������:7]Kl�K[�����͟3��Q�a|�e+e6���1¼��D6��ퟋ���_�\x�;wm+J��j/�x��>�۸�_6��V�1��s7gܸ'r������~���9���Ti��X j�$�g��m�C��z-���?���_�ۼ:�y��6���]M���
�e=���ܹ5g�Ԧ]Ǘ�'�M��Y���v�w>Ghr�+ ��R�`3�f���8��y鶅��K������8����4niA�b��b6$�ԡL4�C� �/+7f�����BG+/נ��/;A��� J��DioV�,���Ohj�yܭ�%�f��A����Ay���|ᭇ�g2�ḻ3�co�ѣ@�y?Y>�,��J�L�"�}�[�tɠ��G�D��/cƝ�tC@r��瘞vK*�I0ٮy���P�� z���*�?��ʛ9E�c����ߝ_���cg�w�a�Y4��X�~Gg�9�-
��L%8wL!�c+iR�s��ǿ{��<�����[|߼��U��z�G����l�������A�,M�A�n��~�#aO�Z��T�gC9z(}��J������0�ٌRӮ+�7��S��_��m�74����e�G�ɖ��3:R���XG�2�P���wV�Ņ��� ;p�w3k�;��-E{c�Yx�����K~X:��ݖ\��X�T]ݭ�M�1.Z�F�XÝq!S3�L�R��̭�kC�!6n�	K���MNNPf�*��D��,}iۑ� Hk��RH� �0�UF��%�Ub&0�y��(�(� �����`Q3P�K�bLoR� �>A&+ߟ/���OIצ��Ʉ5���v�Uvi��ٮ�J�'=��k|�NS���x���(� Ҋ�:�X`�o���v�J7��ct1�|4�.Ƈ�pO�dX�yy�:S�3�Q�=>F�6E;�g%�DFD	z��6H}�@�rC��uZ�a!@@�-(���%�?~>�.!#a�fA�5�&(�j��T^�L��j����"=�LN�1�	X��~ҟ�����^r�m�B���aԸڗ��-�{0�e�PmNKBQ0�1H�d��^���o�0�d���!�Pq8Y^W_{��HDx��2�	�����7'*�B:��J�(I�)�� ��1	
�u�:�#ޏ[��@"�u�$C�7��҈E諀| �Ɂ*�-K0~L����2`�$%(�co,rjÓ���{��#�� � �K6i�U��F�
�$�bP��뙺�`>�`?4gv}Ž����ov��_w�C���N#�D���٨Y2}+J:�ōԉ��j�z1��.�C�K³���"� �Q@��}�����*ne6�B����g�t���4���2&���e%� )���ֆ����F|��R���&f�P�Af.jj'⑅���2��MüH����ζ�嗇��r.�B:93�[+�=����1����Y�B�2�kp\Ϫ��0tԔvA���s7`I�	Nv�3�"�;;6�@$�{���o��D�]!X}t�X��n�ShQ,��Nذ�<��+m{Ĺ�8eK�Yk 3s*Y�#���[��0���m�î������6Ӏr�kqVN��ΐv塷��}Ն*,Z�@�]�O�(����Dȷ��i*b_���X��~�(����`�1.�� *v���iZC�֗C> ��w�`�]ѵ� ��^(CӋ��80���Ǫd�xa!�P�Iϴ�XI�G� ���ԥ�>�D m��U!!r��`R+��e�5�ǯ�ҭ�q�|`�Z��$�fk*f,!P>A��A`�B ��WSLF���J-��:XJ�%��:�,��e+�0�o3	�yѤ��â��\W�_��I6���&|
����q�xu���ߞ:��;��՘�	���zz����r��c^=��A��.��2wV����G$1(4C��mm���~��_7�|��,���w�$Y`���r����D�g��^��!�K-���� >(hBɹ������_��9 �\4�H�c�@J_f�M��Y�3_�Ӳ�S*�le��
���Ҋ*�4�I�+LL�,,�P�T=��j�X�q����r�+�Xn_�E�#�٦MlK�noM�YO̘!j�?�^L�	P��*p�!`�~(@(�,\Gd{��x�fn��" ��+�Y���bB� �%�R���o�⁂�ٝG�Z]yRg�7��U���G�l��1i&|�3�P�aF F'l�,V�-8ٕ�S�*�ỏ0@������	��I (���z�ټgS��̀ |F����0-�@�@E�����ɂ$�(PD�̱DS[�R���e�xf��=,)O�`=��xw�B~�����#�����;��Xs+�tB'&���c�	q�3u1)�[:�WC{ڴ[�V+ýG�{��s{�p(0�:ı)��p�)#���n<�U؂�ǮJ�u7���j(�8O��x2:�P��9E�~S-k$�lVʡ%G�Ҭ���С��PB�5Bq36\��O�Oc�	Ow)P��>�O�0����LY�.W���AKb!�17M�\
U��6���%59F�ſ�',n`8��0�Ƴ�����~�(�9�F�t91����g�v I4,�(a�3���_ A-?Y�@9l�(��W�Fa!(p��݄�E��}��g*���$C�1�|�@D�R��w��;��o;�p׊���o��H1��L��(S'�'t;��G�~�+ʡ�l
̆���"� �����+N�rj�FBIh(�*�ג�u�PJ��*�+�+�a�9*;���Ύ�Au�|�Ö�@l��İ�e��5f��o��6����`�a�`#�,Dhq x���v_�J�����˺�iV^�jttH_��p��C<�P����'B�@]6!
%⊑R.�#���ĉ#/v�P�C��'���B9�(,���:�ʻ]m{wt�����P��1
1v�s��^dM@Y��{١��l����3l��ɺ��ykj�٣:�=����h�Œ/g�i�)k!2%n޺�>��j/�PU��V�I��L�mT+�q ���|2f��l��M��W���C"L����[�N�+v��,�E�I�0\# �� !R"�(��}��h#�����2WY�����r��rK���E��Dk4����6�3���~�Î]�.���E�<W�j3���5� ��ff�����OY!Ԛ�<y�3��V��ݤ+%d'� �$���}ˍϽ�o�	�P�=}�B�I5�~d~��w!��Sy��z ���:�P!�c��~ܳ!���#%���Q(��:����}���k��Խ�����u���[���;Y��u��Io.��ݶթ[?:Ӵݖj@&�"�1�KD�?�ӷ]݉q��e�26؁qx;	�1e��YTx�hZ([i�AUhf�D�@T�z�ɏ8��$��i�K�2UA �Pݖ����jQ�	� 1��홢�^�LT�2T��(?ϩ���zoDd�fYN M!.�� ��0��
���ç)�,%4Y1Bwa�`�EP�$J�K�@SP+ͱ�Zpq��jb��ե��P�+ff��3(O��wr�����u���|��4�dp��=n��<��8�<��5��j��
�F�	"�V1Ļ�3�].�߫�����۫c����}��]r��!<+���F����u�4] z���O;�<���y�'�s�Q��ζ�A`�_϶��+�kk�N|��,�&�P�(��n��ԇ͐M��t�B!:�ob���2��9i%ׯ��`"LQ@�3��bUH��7>�8X��`�[W���b#��.�����yY��Q��A����F	-Y�=B�QfעX�L3pڒHYN��� ��mj�x<Y��P|Pq0^;5��{|)(�������^5��l,��ނChX�`o���
�P��%J�dB���pH��8r�2�?&Ķ
p�w���EZ�G�20^���%?���HO���Ӄ�B,9�B�c
)�7x(� ]��V��aeZ�Rg(19�4�ُ��G�m�51B�"H bT����f� �Y�Tә8����0ح�����~����租�	��>dĬ�$����?���z��Cԁ���!�M�m��&��!��a��7|7o?gr�y�x������@���}}�a��HO{@ c ;�_�����w��ݦ�d��U�N Hj}�E����)�>�x�jW������_Y��2=�y�����n��l\��qu�7��sJ�6��뫁�tWq����i�AbA4 �,Q~���@E��PQX6�7)�� ���q�|��Dx��T�a ��V#���Nm�rfL��4_����-j�K[�Qw6��9���~v�~��J�g��}�kMy1�<���.�(`�ٟ�*�`�J/'�XU٘e�EЩ&'I
�8��!
n�J5��~�_�s���j
��@�V�'"�kҜ1̼s��[NY�6,��P&[�B\ 8��c�˕�6�=7b���^VL|H����J.�+���~�"�'U38L�zVJ�7���c,�����^�f�̗z'f�I4���G����ka�M*�C��+�JF\{<��%���iJ���5*"�[w�j��l��bI6�k��0*��If|� @�������x�(��ec:7M�[j�j���U�Ȏe�}��l7ɻ_;�:�:t�k|�Ƽ*������ZNZDd�^fWG�	hs�2��6��jf��=l��3Su@�m�+�B��%��M&�~r<��T(Uө�~��\�ք�ŭ ���:�̦�Nz���^�T����`� �0E�[_�qV7 z���*�@�u�B��;�V)�Q���b�H��}!UTI�_ �f �6�kl͆�����۬�6�F��"�^�D8�����XRC����j�']\��	��FV��e�Y�\w����Ǿ]E��%u�S_|���83�^�xՆ�m$f��;���g�N��S��
���})�����(m��<�1�=K�@ �z,������w��t�d姈���EVĿ9�R{q��wl�*@X���}&����z�e�n{��u2ߋlz�G��3d9����[�쫨�8�����'Z���>3���#�Q�B2kS���r]�4'*��dP��D�O���jàb1G�U@�=w^�	�|�����J��̋*ޛ&L,j��i  S�b}�� �,�������G�n�m�ܞG·~�Y���F����w=�ėa�~����JY�[If�w�5in�}~� "3��BʚAzK�)�$-0��E-�{8�2$%��b�����(����@�	:�qeGb����)ĳ��;'CR�P� �e�,Z�:UL�XF��]lWԧs&x�A۬c����w,W���v�o�����S��e�l�2�f��k�;Q�9GD�����a�5�izV���{L�N��h����	 �8B$j̧4��[�����TL�d�m@K~����Q �{[S6
A�Ɂc~�}n�T)j�L0I�Y,C��v�\P����T�O��h��-V����'!�f��$��L����g��nɧ�TշBp�q[ÃI�`�/���踸��N �D٘��0�zL�*	n[��sH���� �/(o\�L
ЫƔ�8ly�>�]��fI'�_8Lis"jPrF�h̫m�<E��9HA6�y��(ɋPȊ���h���J�ۑ��.D����*ZIDK�r�B���ŨRp)�D&1���gO�Z&ADQdT2��J�Hc	8�z���7���|v�Ҥ�^).���4�O��&ϰܒv��6����ݾ����˯~�Qg�R(��R�O֢$E
!*�{W�@L�fg�e�"K>��>c�����Y�|gw*y�-���]��:��������,�6�'s3/f��xE:GGP��5�.�(���n.,l���Q�C�?mf�V<�p�2;d�Z3,D���IAP�<c��h���/�[ �VQ�~Y4���Aw*u�ȵv��z���6&��ޕ6��d0VϪow��&�(��IVj�m�2�:"���{׮�hn��ymY~�e"�ȉ��D�/����^>y�h.��R�x��f�����`��r{�@��o-)!]
g��ۃ1�K�+ �T�͹�zn��ОURB]m4?�R��9S7so+���������~�ѝ���4�P�!m]��1��i�f��}z+"�o�,��u�>��d�SP��U��x��a�7w�߿y1���V�\|&<����2@��[�*{�LCd[��䦪!&�t�3�q�����u��l�y@��+}Q���b� �"�B�%�~���V�6��(�E�*�K^���J#6��h�O�T�j((��
a�Ӡ�������*�[~J"��Mb:��ڙX\M���)�8�De��nW��\�|���J��/5$�	����ZPe.�(�f���; ���C�]�h�/{M�gM	�.z:蒖��t^����?k���P�QL��8nIɣ�7U9uH:*�/%�l��z�_��i�)�,��K�R��Y
�����$t��{�Y�Wu҇''���\w+�lբ��;Z�nwE��{��ܾ}'fi�e���>&h�����ՙۛW�}ʶ������S5�v*�������w�v�����}[)����(g�.���n�w`��o{�j��ҍ��-�(�КXpL�4���hG'�[Ɉ�y�jcX�J�i��:��<�nF8�v�+��b���{�;�Uδ𵙁{�^�=��(�Yw�)x�T��T�X��2ns�.qDNǑ�MU�0ǩ��d�ycM|��ݟx����4��7�� ���n9*�-�h���(�L�1%��� ���39X*�8DU��Hҁ'TĆdʍA(�#.ڶ�-���%�0<*���}�v�jƖ���w��{Y��'׷<bм�����e^q��;@�J�7F�T4ղ��H���_����q��I�@�i�7b��\�EOfd��t\ ��a���Sr��� ���K�YB�a�:"� ��}���,���V�lsbҍ0|�EQڵ�Ӣ=� U���9��=.��wP�^���ҧ7�*W��w	-nd(P>�$4AS��.�
�Ol���E��VM�41���
�{ל�N��Uj��P����e�ى�Sr=2`�eMJ~�8�_A��-#�%� 6�(39;���PM'�ciI̶Lg����`D�A]8����DJ��z�ʨ�4<�|آ�xd���"g� �nӉyU0	wס��B�;����/��&�)�����c^)���6dA- �/���JezL� ������޷:�����޻�#�x�t����w1Li1'�����v�!�
J�m� �şx�V�ܝ'}e1$��ae�{, .����;���&Z����Q����(AUD��$s�ίvB������a��x�KF%s.���W�:�W��VI�V�W:췬�Þ~�׮�p�YF�;�ƻI
./e�_��6�s�F�V�A�h���>�v�j�ڍڮ���:��
�^�v��c���v�*�.�V�Q#�\{�m��*�`	]����p��_]��w/���it��N��$�)��t�sc�N��K��`��3 1ـw�pv�&g>��tU����+[b��g������31�:	�b�3�_خŉ��|b�F�xU:J<A�z9u��[))D��t^��Վ%u�Ľ��ަ�y���Ftq˻�Y��;7nevSD�NYnn�W��V�;�F�PpQ�;�g��">P�o<��Y�\�Uձ5%�JM(�|��29�@Y�͘�n�b9. :E��U�x"�b�:�m�wN4W�*��uε{�{;'^9�sS���r��9
�|�]�
n���^撒�ێ<m.6�i�4U%�,�4�b�Q	�x�i�H��
ޕ�OU�����w����k�l��y:
��ja���3��:��,)�m�=%��Ї/.Z��K�$��ŋl��*�7OG6�vژ8�\��	�2�)M12��|2����m�۵���|#��=�d�� SU7.�GA�֧
2O�
e����)uw�ymj��5«����� /�݋�VU�D���]%mh���B]Ӗf�3n�����muG֖`����86���eM�k{��!��Q�ihW�/lRIp־v�]�d����%�z��"��Kdҹu:�?�!L'��oL���b����<��.:�aVP��djvL�ޡ����&��{&�t���������޾ܟ&U���e�{�:��y��PB8�ޮI�&�xw`*�8K�Ax\��E-z|h��'̘����S�� �.b��xۚڃp��=jDL*�)��hw��H!|m�E���w[���9�P
1t��"��c�k�T&.��#�}�of�����m;KfaS��ۻ/`J��:^ͬ��*��4Ι��iT��X6gB��5����ff+�����Q��6\̣77����]��n�{�fi��YI�H�]mf�tÎE5��\&J��e欩3�(�Hb]�%��ͦ���qF] �֥w=��-Ŗ��	�$����.cv����Y����(Hk�im2�f�X1��̺�,0�`��s�SWX�˚�R�JZ96孻B����m�� ��F`���@B�#6,SB��kט�^���-��sn�n����kh͒0�Q���0�m,)��חmi
�)LeM�ԫ��ĺ�l��8iF�h��؍q�u�4�]%�45���4�`5	A6hJ�)�f�l��&b�k�
�x�8*,�\ѳ\��:�٭�U�d}[of�oak�n��&�UUUUUUUU[m��t�L��꺜3��1��v:ԣ�.]�t�;q�m�WO�5�xgI;��AS۾�֗wS×*��ib�&FT�B�uV�ˈ��fٌ��3hb�uq�"�V�#�ු.d�ç˗;D��H����x$�>&����O��AE��K�E����&��C��`�q>N<N�y���q\��������zc<OR��~I����3��ʞ|��N{a_��f�o�Q:��?i��O�,��K�����A�D\���/��l�4D!�>i�1x�T�88Z�;M~�3��V/��	(U�@e/�_Rw�j[�?��.0�8�&,��l�9�a���-1?�*k?f�+d�S}�Ԟ$�c�7Ͽ܇�M�R|��RT����,~�N��� �-�U}�C�z����H�m��v	<�����r��u�d����~}g�z� ���Kh(}�n�����5��E7}�q5B��ND�MB��Qﻦ�߿zw����48��N��u�C��UP�B�g��u�Nǳ����m'����`[�8KC��J�+O�߻�Mg�5��Xc((x���Sǌ��{���u/.�S��X{��Y��������r�އ��z�����iơ�(vw �C���\[Æ�d�/��Or��1Z�߸	p�
v:]��[�"��B�*@b�;��X❵�\wL3��)�0�&'8�c��}�a���Z�s0�������1 ��~~�.�MO���*��`��)-�qPZ�4��-z�3�>��nv� Jq|a�)��󀻠A� d"	�A�*`�R6�du�H�ߩ�hpx��d-��������8�{O^����<a���<C�>N��������s�a�̤���׬�#U(|�|�Dn(P������=y�]��f^�������?=;v�)zEq�
Ki��Ǜ�&���#�,1)Ƌ�:�O�^����S���7�v���|�?S����OY��ML�&��]O3,�'S����9N���'�_z�z�����$���=��������7��e`���������;���b�^�&$��f���hTSZ�u=���9l��
��4��d�'�>A�!�s�5'����bAO���d��P���aXV"O��=�<olQ5��H A3=�����ϴ��'P�/��M��"�w���3\��f�Y��M�wpY�)��(������Ww���1>d���`k<I��~OD�m��ß�r3�̇䚒��R�s���P�?"g8+���2�	mOU���|�fT(��mnY����
�dϿ�GSg� #�@w2�=�'�q���?��q���k�?�����'3~���&���QCY>������{��i��+��ĝqS�J�!���֦��8��^[�:��T���	�8�ľ�A������fL������f��S��v̫����p��i��iKZh����`�Fv�;��&1�������E$(��x ��*.J��T��X��3�����b]���ns%{l���q���S��Ŝ@�w���l'�5;~�'P�ALa�8��Rk5��~����u��8�6 w��}��l�|e�ws�~`|����08&S����b9J�CӖJ������|�3�-`jOXo�y�����wdS�,�<�gK?0�Xk�>����E��7�j;=�dYE�$�{�����Y=��R����q>I��ۆ!��x�P�b��%f����T�bm�Fө�~�q�I��;�tx����>g>��Q�������a�4!�p �>����vL�f����?8�>f0�w~݂��nP<C2Πs|Ì�N}�>����|�j^o��1��ɛd��^;��3̦��PyMDa�w�8��SY_���N��èc�F�T�>dͱ?��}���4� A�";}�:ύU%j"�k@�>0��5�3i�aS�8��9{�y�gY��&=f#�+/)������^&������?_��������}�����/�Z��"�1�C�Lfm���:�{��7,��?�g�8��G�>� ��o���Aj5¡�Sf�ga iSB! �"���Z�$"/��8��?�?�8��>��O�<q��ˉ�(�}�����=}O��55�V�;������e����}������Lj��߳ć��SNr��(���E��o\[�d_����R�[ϰ�jC�e_O)���3���?��09�%IS��0Ě���>��z��Ol ���*��:H&���$tK�Ov�'���)��m%u?���<�9�~����:�3���N"ÈJ���/���/y�鿿����7e��w�t�^]N��-�iw{�k'53˨�"�3R�'�[���Y*Ki�
��v�(�d���: ����u�8�&#�XUgC���G�0�s�~J�,������|��0��g�8�+
�����Z/�&%װNb�d�68hqG!��qy��PQY������9�|	D��P��q8��fa���N��|CD��CZ'�e���O��M��S���(��<H���Tk:�j���)Ĭ�13�;��NqK��R������D`��>xX��ЯR���)nd��?{�����u1���:�d�c��aCS�Q���y8�sl5 �6s�g?��� ��<��9b�È��("O!���q�$��9�k"���'�U�r�򺧳��bL��hPg2b�#���{'+-塭V^Z���uZ+-c��7r��j-m��%0Rt����!=�CV����c�~�:���\�*,8(P���1�!J1Y8��|��\V^���ʝNg�y�d�y����dX�5�����'Sm%g��������Tąa~=����b$d}�9��̳�Y�$��j)KF1O�C��)+%N�<��\�����"�3�������dh���$�2@q>LOSRbx�%�~�����L(�V`�!���~�Xp�|��b�R���w���yho�7)���w0����L���Z��`�Nm1�r�D����Ԭ�d���qT��j޷���9ټ��pvo9u����gY�=q8���J�9������Ld�sg�X������8���:�I�O9�C���;�Io���&�v�O�k:��f�f�D]�Hp�8F�(,��N��K|��W]{T>?H��YI����^)��J�U5u6�3N��*���
z,���H�ڇ��x[���w��	XƝ��F�s/ʜ�M�E*�2�1�baP�UP�!�U ���*Uwy���v�>�C�ރ��TҚ�����	�������Z��#�Z��n0|`�|� i�8��˙�QMa������o�y�{16`�g��k��鈡kT]@=JEA'�Rr���#�Z�ڇ?h�I(�u�(���;��:a�[x�ŏT�٪�6�Ź,�n�3�S����ưDRiB�[2��g��m��Q&�[��>�|_�����Sa�\��}.��e|�~^˃��׬�/l�&'�ñw�뮯}n栎CE�^|9��&���S(I��#E�
�-~��̞���iT�UG��j�Q��^�jR��T�(�����-�����Re�"H������Wj���rrf<k�ǃ�\k�9��Bn6P��9���:�yRX��b՛(���B�n��S��`܉)(ɂ��FuV8���ʦ�+�O�T�^�����[�b��r�fSbGK��M9���(H��k�ɕd%��!��(6�S����6)KF�M��ʺy�V�b�+:,�X,6ڑ"^n+پ���>�=�y�yq͕i���;���4m��t�Hmx�0�ˊ�"p͗j[0�(q���_���e�M��bݲ�%�XL[vĮ4l�e.�it����͒ۍu̱ˠ�[m��2�r�:�~���}DP��E�
N���R�˙��M��?S�ϙa1�p̞�s����;Lz6�pط0n�����^��-߇<�f�}w�j�W�)e��2��X3�z{!����ĬN�S)�����I��.TZF�.:���T��:���	�)��~�N�2<Ldʼ��U�� bd�vّ'|TR�8#Ԥ�С�&[���m�֙w�
��������� ��u-�0��Ղ;R٠��ھp�w��
k�M]����N;��2+�s\����:m��[~@���4��]�� ��[��y���Uz��.3Ƃ��9"⢈=��k�4Q��ۧ49^��D�@'��Oz�?9�oSf��M�@�DP8>~kl�p�W�
�+��f�Ǆ�
6�;�����8��y�*��L�cNv���ʀPj�{T�
\+I#��Ϡ,sqphW=�&�*��S�eUΩ��4�K'�������!�6hU� �|�-�<4}b�h(�f*�)� �l1�\�=QV3��(��\�ŭ�M�CN݉	I	���w�swx��7N�<��^Ō�8�*�'����8���LlԤVL{ؕ�]��H~���uS�<��{��X��@���*��p�͕�Ф,Ɨ&�`ڬl���reZ���Zm�����k	C��UO����W3{5�Yֳ�iU����D��ByV�� ��J^Ѫ�s������E�����/��J�Pc$ԛ*̮�����t�2��<�o��C�+]:�Z��X""f@�I(1'�*�LL��騨��-}�u�CR)����h�]i2��_<u�IC3�Z���3�nZܻ���e���4�w�^mP�N����dw% 9lv8��'�J��y�^R���3��o5�C��sXCI�0m��s���vD�t�A"�$���h<��O˶��:`c�1Di��l	�M��0��~i�,1AQ@坱J���Nh���I̧.gˋUS&�M���Dۜ����'{���3�dF��dK[�!��&M+�O�[d�AS�0�9��K\צ�R 8�����,�Ȉ��u�y*�U���J�s�mk��S��1�Ӻ��7/yy|��y9l̡��d��C��Yoh�F�J7�"r������z���ekl��'|*Lͼ	ʏ3��`��Ϯ�����	�Е3O���H��(ʐ����Ñ�?h��ݢ���ja��9�i�����m�U��l[���O�~�N6�_l��2 �s�v���H��0��WL�B�)��vb�:-�
,J��� ��n�����8��pz'#ܺ�d�IRӢ�~�ؘ��C�#��Z�b!���$U�۵�D��j`��͢C�[��owy��@�K9�{����J�k�����dlQ8�Vy�3��-�l�Gj��ϡ$H�v�)�:�q��p7���ʚ�WNW	��	L!(e8�>�>U��s� �m���z���<��x"�p4ηc�~~H,�&|�ܶQEv�����UT��Q�$��"h��w'�=�����P�Y_� ����ue�5�άs�2�'�}�ξ�s���%uX�n�3"��B�-��)&z����6�0�%N9s+�	p�r�!U�S�W�ܧ:�P��x�c�J�B��9�0�VK�᣾�5D��s:^ndN��r<9۱�ӱ�N�V�v��������]���^!ݶ+9��܏�Z3��25%���؅�Pb��N�D#T��v�ӿ�R�g�ٟJ�7X$mg���.fZ��n��_�w�Q �A"��A�l7�<L �&�j�L�R�'qуc���t�L��ڊaPʅtj����\"�h�(�&0��{>������Aa�UB$��h��ӡ�~���Q@O"���1 �T ab�D���f��q}g���s�)>ja��	�7SF�˾���bULQ��3z���>gR:��l/>���c���L��O�|���:g����\4��}�m�kE��w(�#�E"��;u�*�Vv$���"�t��="&6�)�t�<`i�L�MM^y�/q7)h8� ��6�'f$�j&�&��S�ݟ6��~�3�Z����^�W�
�ˤ=�Dc���|�5�'�'�4��K0I�kbL������vZS�)cE�ipDy
Ğj:���z���&�s~��?��߉=}�p���S��8����y���Zf����9ڡ��|�@���+,�}5IE*)��2k� �����t��=�(���_!�h�	�!Ä����m��0T2�	�÷|��=3b�x�WIXR2������������:�_ `��,��.QT�iu���-�{;�"G�^9�͵+�z}E@���%x��W�^�L��ON�|p��4���,b�����`�A_�n+������Ȩ�v�����·�R��	ǒZ�}j��3���7���)݋��]�(�y�LI�qP/����Ks�S� ]4������lY3�r�nm\
��~�ӥ�R��d�j"�x Ȥ�^�0,�k6����쪂����h׺2fJ�-�9yQ5-��ST�1�s��ٕp���l�&���4v���~�-˟G���Q�֫3�? �A����uZe%>�T��ݾgm<Q�����̐*7�nˎ�^�̙�?n��O�/�ר�6��xF��|d�N{�@HU�!g��05��b;�&���X��@#���oU� �Sئ.�U�W���oo#`�ޫ�
�]�w@3�t���*��-9�'3 ����i9�vJu/#������S��@�rHSճ39툇��r��ثqU��ϸ��<�cv�Ȁ/$�.c��g۾�<��=��^� �M�$���.�V��%�Y�b����X�P�|=Xi7_�E���==o)����+8�ce�o�`ȴa����s�\���"�ѩ�1��fBA��nM�w�ՕH�&�Ԫ�UG{��T܌��W+��"	�e�!xՆ	n�Fd�1+~y����R���M�U�i�����J4�j��y,�1�J��)�ԯ�&"{V�B����宠����o�En���!�+j���t����f\(�.��*�<S�����ʱU�'*�U͐f.��e���=�h�
6��W�����ZaN1���"�N���Ya+W�\aW�&���5���v̹�UĤ����)x2�)��WH`�!͔�a3�1b���O���c3�%+�x�Ӊ��|[�,�Z���v%�^	��'�Ev�o�R���y�O�����Vy���G8;�м�9q,Ys5rK�g��Q�ʍ��=��ĉ��NKÆ6j���Yk��m}^�Q3ܝ�v���}w�˙j�Ղ"]�wSd�ق��ܲ�a���JRG�ƫU2�C3j�^b�����ׯqCD��!�Ŕ��v,݂���|�,���,;�{,�4;dl۷E
��@��6�S.dPq���BT� �e��ku�6�3<ݶV�u����4ƥl4̺��@uK��6�Pt�Yl��n�SR8-�]fk����᤽��t���s���C�7fɡ�r��_f�F�v2��>3`T����!�r��ē�]W����D�����0�xr��t��,8ۛn/�Ӝ�a����1�����k�Y��=|b���JX�U>+6ZS�pw�C�fBt "w�Q[�ު�i�9�]�u6#�=b�58��oǹ�k!�M��Vsoo= �>�2�p��e��,}2�{��l��}�>��\���F2߶Dٜ���3�v�@��Q�ʳ���.��X]i3�:�j����ͮ̚\dt�뷽I�%�2�J���6��k�W��ޡm�LaO�pH��u��l����4>(7޻�@�0�87}�\�!�a�����3��`� �^�~�)�M�����%H(~�����Mjf5��R��d�)z�}��iy��ɯ.�q�����&�P�I�������W����@�!Gx1�|�����6']�`�A2/5����	{/ҕU�ʼ���dZ4���T��}P$�P����9I%��wx�\{��o�T�!M�\�P$Ŵ�VN�(�0���&]+6�,F�O��N�LuSC|�'%a�+f��n��V�"���:�A�%t�ܵ��u�/13����Ј�v�S͹�~�sJ6%�ی�z��*z�k�~�e��W�����?���.'H>t��y��ti��jPj	Z&�!*:#Y^���H�&�D�=v�V&����)0ٿeby�5Gu�H=�-G�SC��@;��$�E�}�O.�T�7�y<s���e����NeL��%цK�1��{�v���5�Q �������c�V��l栢���!	����.f5�(u��ʞN�v�S����B���͎��ьp�e`#j<]8O	�.�����U4- �U��K��6b׼ԧX#���+n�Wt���Te��K�RV7:~� t'8�U�-ĴR�r�&
6��].Ldww2��O����SU5d�'�©��/֞"��Z�Fn�2�"{���$�  )��MVQ�ঋK��|'��O���Q]�]2>n�hR�pW������Lښ:�]��J^B{2�O�%Y5Nc%W*V��G/�+^�Y$�:������U~��L90�����f��_�>�j���T*�]0�I����w&4W'@����OTn.L�h��z��:�8JBBK���:� �
�03�4��ay���GH%�w<��2��Y�4��v��XI��c���*o�ϒ���9���E7D�'�/<��� �eY�юmC)�X�("hv亊\�����oƊ�9<P�).��k��u2�'V
���{�4�_T_0�8(�W�)�<�z��[&D#�T>����Q�pT�d�6WQ��6��V�ӹ*���s�q�)�T�X������ʧ�A\�u�}��M��-�P� �S4�fk�:�'l䴌TK݃��kU���^��4�{��김Tf9��ДӁ��>���\�)(��%P�ޔ�����]���ظ���H����y޺�Gr�1I%���>P���A�8N���8Bp��ۓ2J��IL�M9ԕ�y:"k�5�cˠV�=���r�Nb`|B�-�rʜe7fVh�3�����?�tl�m���������3����D��T��׵��M�r��U{��\�^V��U��ȶȤ�~IE-�N#���Up`�7��S۴q���6�xث�[Hq�Ճk�qiçPhA�k#ji�y�׮��Yx�Rھ��I:_.x��]`�`ǎX\pt[W��QGw6�k�~Ĝ�M��(xڲjC�����wnE.���ɹ5��Z��"n��N��T�^��D9p(��W{}�R�њ�^݋^���Q/�С�R����ل��ҩ�i����)�p<�2�J�#�h�������y^�nUY��1�Je�:R��S�U�"�O�V���O���������&��n�6�{)�˃5���3~-��k�d�fm�#b�?EgV8�ʱ�-��۹�����~tl�~��� ��9GU����(��sIX�9qHP��Z!
����bD�#���E=>ؐo
��VBi`�P3�LM'�1՞�����q4����(���T(���Z��<7�.
K�y\�����,�n�+����q�F� LGuګdCje3�8�7�m�#<��Bj�2����Zl�9]���"i��=��|�m�ϻZ�n.1C��~�ɞ�	Rl9髟�%�� !�a�L8pxU�jץ!\J���G�߾�׿I|׍4��[�jl)Z,γb�������u��^�1Or��W�ˋ9&gJ_�_ᐚ[Ò��sp�9~��6���OmuK�8ܻы�$B���1�5?W���!�@�u[��8X��)�>�SB8���@0;u�PS��QW�V9ywup%W��g�D���NS��*�c\ ׳Qrt�){JZ�J��U(�T9�X}��m�pG�7E�YpTH#Ք!�bhn{;[Y��.�^y6�9I�u8�)M��m�A��]k#+��
�z���S�8�@Z���"`ʏ��R�`���К�kp�h@`�}ok��	\����e�Nbb�.d.�������L����jΫ��j�� ���;�˽��У���˾�wE��w_'Cvu[U�%kXB�y��x)k�DDɛak8�ulDv�/���:���ս�t�H��(�R�[7׺0���L�uw�Y�И���$ߦ�R�[_�jsT�+@�֏��%�wtُiJ[L�uo)Ľ�s��l̩};��Z��T׉^YoGlηpl-�祵Q�=�+�['��"�=t��%ͽkR�ٙ�]y{ݗ�v��4ZF�`:��]j���:�U6*mU�+/(��t�iԥ�tC\��1�ʝ;G8�eKJwcgWS�k�˥�s�\��Q#lR��`r����{q���4h��r*�nv�ntX��.�Z��詙�M�E��ԩ�5�wRi<�������0�Q�>kӎU �<"�ص/Bn�2�DT"g����q�ڞ�+��ecC��ܱs�VAެ��:0g'���n��1�$���]s��{6������r��w]�]�p�XA�i2�Y��2�J���y^�{�[���!����56�:��K2���dӷ��ε��`���_,N�q������t�y�|�'���|�i$sv���=b���a�9Z��Cm�ݗ�cUܼ�5�j7y���5�r�2���J敍+[�v�m"��d*���z�P�!��:��zk������Z��K�YP��֓�d��N�Z.�b?f����`g��yo�L��i�S��*�����Ǻ�4)�~c�sqd���A�r�bI�j��P��T�,�Uۖ�.M�&ռqp&����[��j��F%b�qX�Ϧ�ά�:v�O	}38��0��os̓:_��j�˨A>���{�՜��V6�vri7�!k
"�#u>��k+d�0�g9`WdJ���C{3���B��=Yg뤂�'h��΢&��s���7��L�Ե���P�ɆӚ��|%���]�^^$��^Ef���!�Ucy��֡9A��'c�[���6���U�ߡ��y���'w�7�d��\d�Zf��ꙣC��x`���fדn� �zk�a9��u6UV��Ya^��+;q�e�M�*L�^��ڟ�������� ��W�K�8�&D-?2���%MM�u�L�7E/�f�ɮ�{W8�C�?XAAW�]w�5�FM5-���<��"̝qU�����>Ι5nyG�r�7B�T{w�Ov&��|���m��.�{Da�C�+*���᫙���J��A��0�IY�fYŅZ�{f�,C�Ei�LX+5=���.j�Q��b�nH���yML2��!Xry�0����vǦK��ӑ��*�xt������BH�$#̨��"�ǎ'z��\�v��f&� ��ۻp�'y��Ci.p�)�r�B���嶼��t_��<*��J.L�]6�Ii��L3Ѣ�gv��\&�+�j���8�S��\�*�����НX�]ln�黣h�T$杯ۚO�������������V���Ƽ�v}�I��z�)D$]��V)�3���H�޸����|�ξW�V[�A��:����}��a��k��6�{+�^���諒&� H!�i�LQ�dC�mۭ����~gvW��)�xOC~05��ʡ)�~K�M�H#Nk�ug嘼���,��@^LY�d�b%�eLQn�h�!�܂�Ŕ�S��f�N�QTk�w�	��Bt��z�TvSU+&ӿg{�,�u��r��gE��]�hL���'�ᑕС(���)y��U�Us̹VWyz3w@�kf�T _0�+l��372nyD��̴}�=Ҳ���+���ܢ~o��R�X)�����S�vr�Xå�#�2Z�D��N�5�t,�o@�e���pWԬ�r_M�|�O]�чo�{|��X�*0�I�{��ni��f�	��<�;&Ͷ�K	A�5��K�9�d6W��R� f�^t�q�on��/��cۯ;����͌��6nB�%T�v�i��.s�I
$�m�C}�jm�4����B���]��ϛi����D���)5y�S�����O��եWPU�T�6쁙��&ޱ��wz���hP����	,�t��ށ�xwݎ��R��W7�8pON\��ճ���m��?K����{z����	�Wҡ>��#}����n�c����!8[wf@)D��(u��o�1k��i�>�L��Gc��#�ӣ/nЮm!e�p��2�����>p���[��֫6��4`�L"K��
�^��)��_`Q�,wW�$�͊���:b���q�>Tg�Óp�I[* �wyf<үW��o�ԡ���!>�fT�Oa��FAB�c^�TX]uTA~�	О�j\���9w2�ӶQ�v҇	�T~)�ʂ����x�z��1�畱^ؾ�y!Λ�(��ڝ�	���j�M�p�\]�l��d��7\^�bW�}`�V]<��Z�/�N��j�"b]UЪ&�u��hD�̂�!�/eL�r��bL��l��l@���D�gHp��HFrw&¤�:�M\�WC
m�L��r����;�x��H��.M����U˾<������2�3��/s�p ��ܕF׌��DaC��7K�V�D��3�Q�w����0V@�ݸi5r�lQ�V��V��1a�U�r��AY�uՑ�����PWP܉���W>�*Ng�1WYa�L��%=*��/��C���������r�Vj����5�|grYғ�z�\��mZ�1�騹*����=�\tL��s��񿹦g�:I��e���Q��=��^u�P7h@A�č��u��C�*�/N
U{y{߻C�R@sɴ�o�-�LްwE�n�nW_k�=�C�k:r$Y�R�祋��������ˎ��_&����nIF�����R��n�z��FBy�����:`>�M@3�.M�������wbj��>�4�����-R��eba��2�����N8�<�
�L�9��ߛ=�`˨���|����h��PY+����c�r�(A���ߣ�C��hm�9��뚼��f�3a�=�`H�U�s*hD�-3B<��)�H��F�8�yh82JT%#P��q ��W����Ճ�l%@J^��v,�4�7RT(�5p����5:
܊N3�D>���c��l@)t��K�S�TF/O��T���pMm�VC*���ND�˿tNl�[�$!��6�T�\�/U D�(��j���&`/E�%���7�:�kOWt%5G�����;v��њd��2�M�L�=>�M^]�����+a(Cv)8�sB�W��Jj�(��z3)��K�%�*����E�N���2j���C\	 ��u8m�mt�TIS3���P驀�o�n��maNZ~�h�)�@�ۚ�Ty�0ټ��'"��ӊ䑢E5A]������%�<��`����5���M�vL(�/�{O1�ؒ��<x���1��9ٟz|o�T��@J1#R7�R��Y�4�C���O��G�s��w��yz4�p��q��%�jLzs�eUy�,2Z�KQ��H5ieR�����������aI��L�L���]˪��
6-�
,�p �S���l<�;�$'�E5�d�#��L�W`����y\ͥ�%Y}z`���6�l_HH۳��w_S�2�Q�Y����/Z+��hp�
Yݫo{{���B<����Ewo9K�<��AL�d�z<Z�c�������O��S�ή;���N��>�]��ע2b7�Mp�;��fۢ;�cM��L�+���w����A
�z�xzs�6�Ɍ5rɁԾt()}[R��-���+���3	Wq_X�xTKHsSh�x[�?��"�Q�S�w5�6\h�<VfU"�^���¬���#6[�]�\�����ʨ�G,�mp���WC�)S��c��©�	��uS�z�C�1Cź7���q������J�ޠ��K��6��pf>�}�Z�F����|5��^�v� �r�M�?Ifys*ʞ�����=A��[r3�by6t��2!�^���t@<#��_(.tˈ�M�a@�(��f��x2+NwƲ����T=W�k����V1�jX����>�2��L�m����Ac�^<��,#L���ot�3QUj+�bܵ-ک{��J��4oF��.<M��U��y�Z�*�_AD�;�=���E��j~*0D�	d�.l�͚ku�Ci�e�c�����{� �p���j�a<R-�ힺz`�=��r��Ϩ�ނ��'*S�vr��G�bs�|�44ʞˍ��p��q�nM �����)ֈ��74�z5���E�z&)(F}-�H@��0���7��\�SYV��&h�&��Ku;�\jh̊��uЌZ0À�+�z1dy��O3g��f�nf�J�y1(� F@0�Ek� �5xh2@����M���w��wd���;I%�ܹ�3r��#�m�豆�`C�u8|$ׇ�t�!� �!,�Α�ťh����|����k�6����ʌ*�E�N��*�w%8�}W3�%{���C=�Ts��Q ��.�j��c�2q�bX�ѓ��J_��ь�`�+&�vxb�a�YU��^!]lU�P6D-L�yj��͉��>�d�x��Q�P]��@���7�x135�X�O�'>�nI9�FW�o 'f)�sT���o3�o[��bފ8j�:Ȥ;GQ�������$�9�a&�Wm�E��R�R\M���p����F.�R-(~2=��T�	�ش���MZ�8���7~�!�n#���*jȺ�Ff��:$��AŃJ��!�9%Zp�\�^����=ھh����1ξ��Z-�K��M�q�U�����9ޝ#���.�C�^�JF�!"$ƿ5���^���i�e.j>"n3)����&C���%��Sȩ4V��8H8�)�ED	q�;/*�]MUD�^��d��oL X�u=1�}B��b���J����.˸c�>K��(�.�$*����@��(;�~s��ں�M��<]�[���)����>��,�C�ޣ���H�j���ON��c�Ď�v�J"��r�a�����S`J�!Ѻ/��z�cd��������7f�2���P�;��="�����3i+�+*h��n���{T�jԒ�bΞ���R��/�TI��p��M��$[�6�0�'��0���a���[e��7X�rQ��y"ܹ3�+�d�l>u��:e���n���]��Ϭi�ױ������;�ދ=|uu���m�\�i\0�3y�g�w[�m]-��[�l�X3`���C��]71Ev��&��.���u�`���kfX�l<ma��l:��������ڤ(`f.m4�m琉B����ܻM?نo�=�zf�&r9���1�1SV��h��Ӻ��ˆ���X�^<6$��8��H˞ÏO�=�� i���[F|c�yA���&��ߕ2��L�*�\��v�ü=9�S,[��u������^O�;���޺q��)Fq��$��D)\>��&3kc�S�A�L�t�(���$$���{�	���Ъ�-�����Bfۨ�^3Xd[c6_�aJ��r�k/|Y�S���'��L��ngf�W2�ˇ��iH�$B� d�|E��kI��}Z1U�\��HJKt6z�˖�]�~�����{�(VW{���jL�We8�Y�.�_Ќ���U��v*�߰�&�4�*8�֭��]��ΰ��^/�h�K�}w�ǺR�Lc޺�u�srt�X�S=�e�shp�����ቮ�d8�2$�}B��&��1$�[kՙ�v0&M�t̿\�rJ����k�Lv���Y}3�e̪Y�{+ŏ������� b=vW('(��v��r��u�Lg�|���>�Z㣱9���c:/��ښ7k=Xŏk|><cq�C0��55���.��0�6��T/b�_	�E!>h>3yB���gՁe�^F�x��l���_Eø� ɥ�!��&��s�BW����*V~
y��
�Ma<~ȼN�M�vi͘�;��Ġ�2�N*�WY"t���G��7N�����Ŋ:����;��3���Υ�� �g����ڱ�s��p��;�p���đ�6n�V�B�7��D�;:�[\I&K����2B��}��{�Dմ�%��Cs�a���H.���a!�c�h2{Ϸ�uR&e��;��F�e4�[_9+�n�Ҧb�n��ւD��<�'�F��=S_r�%�c��A-��X�ޡ%��/!⺏<.�1ckR�2��;�&�U�=�B��F�2��
 t�Ax���_�K�`e>��Nc�w0�vg���m?�w�����
ȣ��J��י'��y-A�\���cضh�X��+�0�@9�s�PnԋgJCt�X���BwF�睘c��������'@v�6��ȚG�+��J�e߯_�L'�0�TP� �ݳ".8�y7/B�{�4��1�_׹�
i�>��A	��.�O�����!�QCq\/M똢t[�v�n%pҋ����`H]��e�DQ&�z������y�w��
�@(�3��v,����Ua���r����E�	�_S����w�b	X��q��u�c�Wf��
�������B��a��I���:�U�<�A1P�����Ϛ����mT�L��Y�~���@̪�Gt����T�b�AEE�G��+�k��j'*�}<���ٰ���\�z�ʑV����܆��w��%,��\L[MP
���ʸ�n�A3�3D��r-P�P�z"Jyn�9cۻJ�ȮV(�*(��Oe�����}\�w�������x�T;�3T���FӐ.�K�(v�1�w�D�9�g+�o0�ؗp;t3&u�n{� (��*c�o�6�k��'s�ms�������s�]u�\��v,�l��1�
�.�q8�ˇ��X
&�1�by�L
�|��$�������$��~��~�A�3�
bV?r�?�yA�|�x�^91^��6"<�{����3P-d,V��ױ>�����Bn�P���^�^o�-B�+	s0��yb�Jd�Y�6�R�c� A��R/U�M�c��]G�G�9����>�6aJ8�n��H3x�I�+�͹�%�����Zw��B:ށ��k`�SqcmF�����H�rF	��TK���IX�],��9�mx?Z>��c�h�:�9���U�Bz���Q�����#����@+SI2k��4}$h�^�iN��2�����+T�.��\`J��� ؃��wE'|޷��g� �B;,���<JW<m�3��}�BL��zG�8b�����jq&u���΢�I����h�4BZa�Jb�0��	wo`�Q
c�[=3I9����ּϡj�SE��K�/����;=} ��-Gk9�ʨy�����K|M�t��(�lЌI7�++vk8wm(�&�F��'H����L+�Va�}X��7���ϗ�aD��amw��� ��^C'�$(�/����.�k�2h�z#�=.����CM��g�h�F0���:�K��Ρ�sl�n	W}c�UYS�ws�y��3Fq�k����N��-+U�86;+���|2;��O<N��P=�άNyי�w�޹Υ�k�OQ�[�R�u�'���=4����k��3)��b���sz+��=�+*bz)/c�3�%�|���WE>W<��1O�H�bC��M��+p������G�j�����CC��1���g�R}�]zq��dy:�E]g����a`Kų�@�V]L>�h���V���]I�y[��;}[@���:��@���xQ�d�� e���]����Se��Ȩ�*�0����IQt��T^B֪6P���v[�����[j�q�5(��2;�@�zx���X!R�qO}RhϺ3i�)'S���!���FZ$������r��ˀ�R����FE{o����w`2�O��E� �j��:��KU��~.zO��(i��Y�`3[M9;z<z��{��R֑���<j�+����j��盃d;pr��9��v�s��gB*dcp�r'�N3w����nY^��_8��	�3CDH��P��n�&	q'���q�0��.=x#�Ob��|�4�$R�Х[UV�9Gp��at��:�,b�ZdEE@~����R	��^aÜ X�g�fR����(>��(�Z�RI��}�ݩ��fW�BڙC���2}1(��7�Ѝ����'
�D��Q��gŨ��'�W�16�X���L�b-`�O��˓{9e��X�01L��'�5�.Nw_�&e ϯ&��Q]����h����5���Y�}�]"��D�`�ߦ)�����v幝��Q�ٗMww]aɹc�:�Y�%t	<��wr�޶�2v�-dʗ��1&kI��Y����1CV���6�5��l�;�[r�kV^hT1\F%��K� Ńv��SKE>)w7f鮦�n�f�9�mAՔ��X�y��j�����Wl-s1r��l�h,�I˿������(��c%z��#���mS}�$�޵Db��W\�5;��c�ǯ�)�ᜌ{l�.����5s�+7�O)"�t��e�E4��]�"g�mS�
�/5L���\\�/���P�=x��0���7��$����w�tG�g(�O\m+��<���k��E�'��h����Ϟ����0�f��b��/0OuWf��t��˯+��%�ܓ����k��׋��&T8)2ז��8扝>\$Kفޥw������P��@aB&����D,�Ӫ�0UMp/���Ŋ�I�������p�'�ܡ}�L��0����'f7#y�1���Er��/�z�p�,�]@�@�� ��m��N����E�m�9|�e*�xCKك ��*�����	>�s~��䯘�����{{I�_0a�y�D&:-鸐N��3]U�U�7'�q �K�K�͖�D����)��_�
��iv�4��w]I޶�ւ��R��/(Ơ����FG�.��+�|`��u�Iw��$���2�qW��!^�e��h=���T�+�B��N(�u4�t�MmO��K�T�d2b�5�u�n��L��gNC�1���(s]��)8��?�bg	�Ө��6n,YU ř��O���%g���"�A/����q3��znqB����l� It,��u�s�qmp)+;׍Q����Iv���ww9,��f�a[};�7W1�Fb�.:�E�z�,n��+C����Q-�ޢ6d�w�-��uW5&����t��Z�N
|*�J	��n��wZ�N�nBl(\r�կ���F�X�v�ݝ\�l�.�j�ӞmH�|P���]�Р���P�]��ڽSpR�u�@*��_Vn��2.�fe
�P�m@o���IA�5���F��]�j�:�X%ΐ�j��R�Y-6w*:��+����qP�_����+W���֜�Jk����Ʈ��z�~����2���vܶ�;��f���w�G|i�,WGٜrU���,��)݅��������u[�K�WWou��J���/;�����FN�L&ׂ�С2�Ȗ�zrVX�b��u��*�s&�{H��x��<��Et�K�y]�:�w0�Z��@p�F��ڗY[7���ٺ���۝�����k�;�BT9|��v:�f'�a��6�zĽ"��-����fR�Xժ��V��!��-�&щB�A���E��0&t-�0����=iJ�w��S��vu�e����Ժ�;��V�g�tN�r�p��Ы=V���uÞ:Z�
�ƛJ���O6�f����6�f��},;����8Gkr�o�,�7х:����e���ʝ�x1��l I(;<X��kU����s�g7����ni�gC�]*��s�Zs;���0$��-�+ǳ=Cq�:�>f�m2��X��6F�3�;7��a+"(��eǦ���}CUUR �a��� ]��jJY�R�)Z���Q���.�(m������^��5@V�X�U��ə�ʄs|Ft�op-tYܑ���5�z/�}/wr^��8��󻣶�����,�S镜�W(M9�D�
7���j��dI�A�sZ���hwb�y��w��YRX��T(qSy�&Q�Y�l�6d��n��y.G��s��a覺o_P���҂9J����F�zh{%�v��&ќ&��pѶ"�D�С�
�@6���Ж��������♛��|�=bJ�4��
9�?9��	ʢʨ%@N:���{���;�mΖ�RuZ�ʹ58t�n������g���]5�Gri��ڀ�r�FڈE��;�{Ӻ��ޑŏru��&�n�v]�L]�sYc��|ݷ2ۊYI�
b[X�4,j�i�Vf�ڜƹef
3˛tΦ���I������iܳ�kl���+e���-�c�Q��yw0�i�2�2�,�1H6ms6�1���V�4�p	��yu�m�W$B�-��̩��ڼںƥ��3�^d��� �x��c��sShj��P-����^��4s]�Yk2�U]4�u�b]��a��˪�يE9����ꌱv�Fe%[4&�s������ך��y��e�lb�[,��!��S;k�4eWZ�..f�Ʊћ#e���#Y���Θ%���Km�N܌��]Yx�nٶ&���e��[�c;d���,��38�Zךی�֔��C
]
2�Ș�s��1iv���kNm*�UUUUUUUUUUUU��O.�ߝ�������K|���۽J<�'ee {!�c"�ƬC��<��^EU�E89��03�u}}Z��}�m%��9��]vkt؉��C�QQ7�����z�6�w+1C<�ߞ�\���vúr�WRƮ	�c��JT��y�￤��>`=�Wctϲ���K��c�<5#�Q,S�[q���αt�ضk�3,���m�jW�� ���3 ���a����8d�/���΅\k0�N���479�+r$l?�����v��4!��t�����e�m�C�
���g'�?gs�I���E-�#3�����tGAn�Mg�yf]M�J{�-�E�<��B�=�&���Z�Uʮ9�8�%���SZ�a�"�H+MM8&u�9wI?V梥�пU��Ԝ>TG�Rc�n.=(�B�q�ow�2�O&5LI��u���ݺ F��Ǵ�s�ƙBff(5��%T�K����8�|%�>�K������q�}�Dy)yIПv!���b�z/�,I���x}3���Tr��Z8���TN�K,�	���σ�$l�/��aU;{��U�׼�HCVO(A�[���Ap�=.�K���є�/�\������}ÄJ����gxk�!Hk��<�;р3s����Hx�kG)�<�F'�ά0\-�p��s\߶�f��w�B�X���C���uFr��3(�:Q���3�F�os����:Th�2ȕ�m���7ݗ6�9w:�\��`t%�|��GQ��$J(7�. �54�`�)�����{ʏ����E�F��p��!yT�x����bU��'/_�+Kܩ�遊z�'������c�Jy"։�S���$�XyV�+�}�9��Bw�`B)�S�G���r�+W�U����Ė믍������ш�{�gX��dė1-�/K�X���E��Wm槏M�Í��.0���Fby�ܢ'yKL��04�a�#�XJ̏NZU��Q.�bwV�V�X�8dUh7�ZP:B�O��+23�DX�+NE����%�J� ��8'搙��nv2sL�:�O�G8�={]z|G��W�S�7Bvr��E<ȷ���*��)�U`��8de��$N��tcs1(s����Ċ�����4z0
��孯�_���+��Jl��(�W�ފJWf���fh�R��b���iu���dnɔ��98��9����ѫ^�b_�j�_>[;���V�NQ��h|_׻:V�P6�*�11v8��iԗd^Bu���4���i�qR�'T�Cȁj�6̈�����}ۤ�1����s��LQ�D�'˨����C�=��"���Q;�C�k]E�ܒ�QOL]Y�-��c�^�su �Y��^�_{��A8`/p���s��K�jg�r��5�;���a�sd���uI��[�E��?]�{>p�fʄ �jbW�ϼ�L��RVpڋq�ğsS�9n:���U�T�n���{t�P���a�^:�Y���'e]xd�X*7WcTG��?�q���{k�:;ǰ,T�<��p��^Ix�N31yꈋ�[�F�h�3ʻg)�d���$E�>޴(}�����L��'d�U�n7"ż���~������W�N-ձ�Y��V3k������Ȍޣ�����n�BXb^��*��+��*���ܑğo�Yۜ��nƮ���Gh��n쩻F�Hd�wCf��4jU��@��v  d(Gi��i��dy\����'#��~�����b3>�uY�|�n%͂����������FS�T���ޛ�<�`�}kUӹ����K�GQ��\�Dğ?M�́Ʒ̶mb�x���D���_+-���hoǦ�*�aC���Z��|��g	�d�j��B��X1�=詭>~����I7.��{����_��P�k�>�ZVK�#ih����w!ǲ��u�c���g�Y5�>J�ʛp��+�I���#4wyz��D�e��ږ}����37��i�y-� �Z>���_��&&Jf�Ǎזj�	���y��k[UffMPʾ}7^�D���"]3���",�#�a4ª=]
`N�h}餶����y�	$b�Z�L���P�j�|0�nTEU|uo��O6#����S��B�#=��Z:�C���ދ��J���>�hMLy�z���
�G���l6��qd��������"d�5+�QD�ɕ���(���/"��5��L/oH�؎Ӊ���ej��8t�ִaL෷�q����-5ʾ��4��t^zTlW�MǮ�,z�S),�T�M?_��1Q�Lr�tR�P1�K�
qK�}���m�yg�j��S��xT&�����I�~�8��8�X���,cY{�&͓l�'�1io2�!7�_d���5om��[���P��YfZ��%�.�(�˖(��ox��\:��L��R쨬��ۢ�C*7��#�eL��b*a�ՂA�)bu��۵&��nj�ԣ����M��KI�1.��v�Y� ��GbWA-co�:�i�V�tҶ.et�`k.Ū�X��w&�e5�e�uH��a"�m��6X.6��/ޚ5�?�!���ț��|��^�&��K�ө?�ҪTyz���4�r��������)&i����[(H���׳��Kʧ�S�!T�!K��S�2���P�D®���g�f)f��!��![����cl^U��>��ow�,��Ȟ�#՟T����[wy�)�U_��C#�Ut#r��	o�+j�>3n�����>�����r��L[,d���	'���*f���>�ؼفn^���w���vJ����$^����G�n]��2��gvI�E�y5�M��w1gכFn�kMcPb]�����u���b)���*ޫ��;�4e��'�O�%��\�(>��]�~'\L>�c�80��)z_���"��X#�'�b����{+ޛnG�Ì����9fw�I�
�Z�'���Z���H�W}�a�k�J��e�^f��������|���26���l�H�2+8��M}��".�L���I&�JR�0��.��U��x�wj��g��¯�}�$�V�f�y�z���3zKHa}������ɮ�p��g�)ƍ��ug�h6ᥰr<3����g:و~�4^�!�Mt��y��|�:Y2��w��Dq*���B�-4�8:�$ e�����o�}���nO����WO&R�z�h��R���[
��vk�!*��6�oB�N6*q�-�J��Ί����_q��C+;�F��ȥ��'o_w^�m��Pwpj�%�æ�����޶B�R��߸��M����0�N�AZ�����
t���Ë���t"1�7�}�Cq�w(ǥA���#XQ���C��}!��ja�	�̥`��N��gO��6���P~�wax�x�a�J�*����2�&�BwW(7������
=��S�dL���>�2C�_z�N}���Y���NxV�c!�P��9����ީ'����fu�m��B%����͏f�:�`tG�o=p,^�TI�4u;Q���O^�$*DE�zj�f#4�ҿ3���2�f]��-�toc�H��y����(�0/�~Rf�ea-�漢>�?,XV<J	>��R332TT��[:�>�m)64B�
�Q��p��V����i�_/R��p+I��S�r�e%��e��R�OU�=���Ԓ��Ws2���̥!���C�0���
ې(��h�q{o���j~�۝���""��V�qأk�ݵsk��|�D��Ԋ�bHr=�� �j��I[���F[w'Gu9����W�q3��b�Vj�G�m��Y���ߧ����Z��>~�����ڒYg��4�hU����f�3��!��U�3ۗ�~�}����w�+�lL��h����p`�!*�Èx$t;`��a�"�����y��g���K�7ݬ��� �ԝ�OFr H⪓gB�C����wz��o�U�U>��n��m�u����cbf�'mY!�>#���z�Er��[����ø_v��^�������@`�#�EQKfع����k���=Kvd���ʛM?EH�}��e���Dv ���
�*b*�7W��� �bu�ܖ�p�G@y\��[^�^�GT���W�����ANi���Нʩ6 o�'��6ؓ��$%=�5wr����-\ ̌�x:�_�@[��7�[�^ZÌ7{ǲ�zq���11�4WL�]q�3�>&h�<&�f��d30�w���[�貴�!5g,�>A+-��g�:t�=܏Ba�R�n;���������b�|��{E�S����Y�Ť����\uV�t�u&:Z�+���؊a@D�L�yZ�s���zn�$��{�S<��Q����B�}�Uz�i�Һ��,I��=u�z�g��t<�o���VN�GPV�Ҽ64��R����A�v�Ǘ���{Dln_�Փ{����ߍ�\�)C�����3٣�s�C�L�}7��7K<�~]�m����|�%ތ�:d�1@���
J4x����l�klP��7܊%�}3�u;�ь���čuK�S�,�6�9�0f
��F�b��ݺW���H�Lf�G��K�2͙�<���-�&�SY6�]���{jH9*�mI��~�{}��6^���ҳ�����Xohp����f�l �p����eQ�N�8`RY[�=T� �(G7���~���N���7~�G��(	��P_�[�[K��%��8��{e��/9�ݸ����x�n���ԉ�N��ə�Gg㊄`�	�x��{ݳ�ek5���;�7\���KӴ��N']�h]�ιi5��y�ѹ�c�^��T5AN��x���PdV�/��!�kc��c��WL�N�5�	�2C���1{�'�~ͭ[W�>	��?lۡ�0�Y<��{�HhB�]X��ڻ�	-!��I�
��z]���;��zT��Y<ws�̓�LІ��ו���%�_d��K���������Y�r�K�bt���S�n̮�\�ck��-���z�̯)��E�_��|�ް�d!��9��.�n磠��|
Jz���'eK��
vP����L&"�ut?^uV�PٷUf���^	��Z��u�1��:,Ϯ�
�%2 �M�e��)���!� ���Lwu�/���$���S�#�0��髫bk�Rǹ���f��U�7R]���^�!� ��G��n�����S�]����0\���ByN�� Ŀ�iJ�@�O��e�'�e�뚿sv(i��r�� �M{c��.]m-��F;���z��J�Ǥ�<���P�:�*ct�Q>F�t6��;<�~m���6�������\@��B�,�}�.��u������8`���l�;Zj$�!u�i�:��Wf��_y��s9��C-���BQ�[�f�8��s&�1��[��mj�ם�E�����8������!̧G�'֊�ѫ���Z����n�ٻ|�/�z,rW�H��dn�U� k&<8s��E�,hJ�x�F�4�����%�""�^���?.��y��;M�i`:�S[51�6�ڥv�j�k���Ū�4����M-�Jj5*V�h�ٴ4��M�[-ձ���y��++�n��jb�dʖf�,KF*�mʫ"��-��umc��@�
�mx��V-"��+��u?�2��t�-���lVZo�T����R��SB�� ��T�U�k�au���p���bCO� �:Q��V�r}�jf*��ʾ���A�����vT�נ��v	�(���y=��������aո$O$��r�s!h,�w�>�}��+^�n)� ���0�|�����7����w0�ؗ�P�Q�1�m��O�ª�ە��0����\R���3h���hؖ+^�)�vH-����Ƚ�8"���ۚ����ԇ��A�Dz��"m(cX��Y!m�y�)8S@��Kn�K�]�Q4W�6��7*��C݅Az}k6���Q�Y�Ѽ�-�ѽ��Q�)�z!U[�QyTh�\���6aN���N�[F��7K�Ӳ��bhM����kR�)�����i5r@���9�ziB�xy������r��-֨ C��}̗��`��Z�K'���z;�,���NQ��{9h�)�_�V6�S���J��p��H�kZH�[u�s�種����Oޤb�bb.{B�Lv��\ڏgm����mӌ[���_Ebx�.��^�[���q��S�[ȸڥ�Љ��|��7bR���(O�B��W8}���z�B[ i0v��W�GH�8�W]Zm��;�2��N���xA{�&�}]��s6�Y�H~�a��3��i
��&q�~�n|-/5��c�.[R/�[���n���tٸD9ꜚ{3F�y��Y΢G�!n�\�Ͻ2���g����^n�7h���8�Mȇ��F&fff��o�۱z�(�[�6ԃ+��(8a&��x��/�à�@ݫ�/�c7伷��Yqdf) �80�E���$�\N�p1�Pǌ�
�,�8}ފP�J�d�A��VM�ڣ�?�1�v���8)��-݊G�9(
5zO���2
�r�T��{����%]�����*�2n���۩t�K^�Dl�t
���	�X9��Mn�g�R譵8�bo�M��l�[��~1��|w1rĶ_I����ꮶwb�,�n�au��$�6��v"y�چ�Y�v��Fou7�Hv�0���c'H�����.e��k��Jmmq�c5��V���2˶9���&����v��+��dNQ��{�휨�=�t��H��#x�}q����>�ٺIuQfR�q�5�ણ�'�`���jYdU�������G�$��}Ez�f�%�Xɾw:)7�]~vCml��0�#VcGF�ʇ�S�f0�N�аF9^g�9l�#nd��[��e�/KP��쫨�!��աd�mk/�ƭn��(� Ձ�e �^MO*6��J���ϟ@��3�][Ʈ�m�㭃�a�5y�.s6�f�M�T����ʍ�̰7s�'ܩ�n3�����Нdn�4p���*jZB���:6HJs��
�C�Rצ:
A�E���cӴޗ�U�l�^9������[���~��i�r=k=���\h��7;��Z�x%��0�,�S1�fat��r}ۍ�:Հ�ۛ�ު��r�:�_�Pt�������W"�P�w0��!�h)���Z��L���Չ���Ni{���1���Kd_���N[���qMVW(�dpeL��Ф4;q������������O�c�ZA���fr�ͲXt����~�d"R�⡏CYL�7K���$��/�m� 0P�i��V����s*\�aX�ʞ�BF�Θ��A�򣻴�c���Y�:.9��fݓX���U��|u�au2һ}�[U�!%�� ��;*�i���p�.r�� �f��#ۇ=�P'�7]��.�}=������s ���_E=�į�^`&�LA>�=bҍGՀj�z�Ťh�uO�����ʑH�B�aX��.��b�A���:��4����/F?.�Cl�x�k|���f��pZ|��!d�j���m+�./hʱ7��1B���r�E�<urs)�!�>�@�S\�F�bՐ-���oٝV)}��F��	��n[�r�?��t⩅��y���+e��S��oy�.U��lP�Cv/L6����R���<�qw�.�x�l��Nl�DVm�P{�ũ*Պ�6`L�r�:ٷ�ܲ�ϖ��B�S�OWw*�G 3;�L�Rhm�_
6DT�u)��r���ˌ�`wՒZhnE14�쑂!�m\��+cD¦�D��Y�#�j��Z���Ҭ��la�F�j�s��;h�=��I2�ӜL�ptJu��%H�+0d��(�6��M�4U�9�3H��ѯ^fH�Pm�u��2����!�u��y�>x�&�w�!�ݮ"���勗Q��'�l�[�E�ӽG^�[����5t����r�㸶Յ��^⼒�b���N�'*	�[�^SFG-��`?�B6�CɆḐܹ�^��6n}�"w9ݵ�c�#c�'BМ��cZ��Df��I>�k	ys�	�����$`��{-�>��c�۴�5b�{(�������S�`���G3�oP���N�����#i�Rng]s���`2�n+����2�Um��s-ꖫA�|%�L��Q4�2�C�����wt�g�kE_M0��7��M�A���f/A5DX�[�B����(ln�pz; �����v��XBu�7��mpiY=Y����VN��u��w���y���J�A)y��+(�+Pg0aG4*Y£�q�u�h�����隻�����@�-��y�P�Cg��K���G3ul��u�Zq�p��L�Ob>�>b�4�كvn�tb�s�Ca�W���#�f�N�JV��q]{)J�SW`�E�8��a� ]��ݟY�e%ـ*ڂ��F���"ü�u�S������gnc�w��t�^�����n$�4,�qL$�r�l7wvK��;p���Zg�����F☂���d��b#'���L9�,9�%Á��jU�
9z�i��؍�	D�ז��v^*]��P��G��tgMb��N���
�U�J\�刜w�S�'&U@x��w��(��.��]�6%]#����D��;��\�������PO>t#9��9��q�n0G)]��rt'��2��@NҤ�o��u��1��l� ��->���y}�^��a��ҕ�O:��[/n	i �ä�H����ij�7�j�0zǯ���_y��!uz=��\^��m��á�����<�>TY���n=
�#��ц���s�|8՟f]Sy�7�'`i�@M�W����
�=]��FSʑP���`�Aόaj��"���-U�%��Ee,mᙻ�f1͞�u�5�,4�|}Л��|ė��H,�;��o�B��}������X�,�S(!a�h������1��G�e��]��_�g�֜���b٨�`<^�E����C��C����q��:3�C�ή��I�ސ�:�{�ܲ�=��� zG^��G[2;��6�!�
}�Z2���#2�j\	�|hPc�;�Q���X���i)��T�=�}`��
�P`zL���|`�Πdz='+g��!nY�1�"���D��e�+u{�#@��L`^����E�-1`Y���7t�	�[�Qt�6^�!?~^j�<*C��/pW��p�)S'rȸ�[V$5�n�9S(QYM��0���h�JfV��s��E��qBa�k���-u��w����I���n���Y��g�)_>^�n˻Wi�ԆȰ���)j��%H#�/2�s�V���h�ԄHA 2ˉy�`	�t���ثn[�FV��n��,���ʗ���I]c��k���Z6�ˆ����vl���é>���m�:�����*yұX�(:��g4�"�Tk �^9�����
���84,��4�]��O�~��rH��|`�@�|��V���Y�/U�~���'�J���$ݫ��]=�)�}ו�0;����{L)&�V�Ϊ�Y��Ç�v� ���������4RͿ|$�y�h`Ѱ#]x�:�ԄbÀW�!��E�#���ࢄ�r�.L�x�O�xw_�%�W@�u>���q�*��z�j��wɐ�
q�Ic�������D��&�.=.vtN��麻���vXӓ$����$%�o%I|�.u܈;ٖ ���|N�J��0N�6ק*o�הּ�kS�D���	Hy��pH���Si�[�iN�>����I��51��l��.z�6�,�kH����"�8a��ui���#x��ot���*���
B'C1�ɫ�):���b���X��ti�<��7�R���Fh��xS���싚Ňs��^�Z<ظ.k_u�wF��j;�T7�c��é_�H�}>�UWv�KN�O��F��G@aPc���JB�:�J���w��AɅ27	i
4'��v���by��F���h�%/h�&��j����W��+�i��hzBT�c����!�̍V��ߨ�:=�c� 篪�<nnD�[�Sǹ�6�|���/5��U�1ld�Mv�l�h�/��3�w�ѓ�`'�麭�!��[:n�]
��`t}�=�槗���yS}�Lj�fc	h�U{櫮(}���M��ߌ�P(����t�s���������X��#�L^�i��:�=�MG��9���%:ys�ދ�R�z�t���R��c�LF��,����T|�������SX�n�L�]�K�ѱ�;y���{-��,�vDF���>�]-�jQ�>󫺘!{�F����R_�j}�&gb@8�N�kA��b�w��'T������xH��{�E�� ������Gq�az��پ��ה�����{j{��g�Y�����V7��m�7M�WhL��*�PEj�s�]],�ys�����z{L�T�YDJ<�ٜ���XTBM±x�e!qF\Ed�'��u�-2�k���I��*`�a�{G��+�h�m<�D����RM;�zi�9�.ݳ�+���[��YW^#@ojpR�nӰ�ncBI֚�޵;v�^Z���Ե�;5hE�q�jnR��$H���39c�V�+/S�Iwӑ6X�b�i��Ą9DĬT~�جY&?M��+��eY��nT�t�R60(g��W,w�9��0���yYOr��)H��Գ�Z��+ԝ��ld�Ppi����lS~�ObJe�R��`;o-1[�n������e�J�qy=jN��6>����U���+3gxF�Q�gHy�fÌ��lYQ�hQ�#@�
2:yj�~���q�6ҋР��My/��D3���枓o��)ACy��愼����Z\�?��c�ׄ����71؎9���.�9��� e���ϋ��{�*�!�73�Jg��?� y�G�Es�,�2p=�\��s��j���4��o�ߓ�p���J�՘Uzy�������%>��q�[�`3�u<��
���c���/t#)R����[�Ϟ}��@R����J2��R0�$' ��f�|�Ǡ׷�T��|����u�	K�[�l�b��ү˟x	٣^m
��%. ���̀P� ���~UN3#��͈ѐ�}�W�[T��y}��Bj���:�u��$ߡ-1l_�@`��L�ي���[���W-��l@)��n�U}J+��u��@���+��I��"5��P�����1�������Q����~���!��k�7q�����pel֔k��ݤ^v��;�Y�9KV0����S_iWb������5L� ����cݓ9�S�;�ьmxԉ-oW�K���k���NhѰ�G��V��{7��@��;Y<��aj��tU���z+r�J�m���z���C���N���$�9���>�O.���*@�q-�r��xp�/%׊�5�V<�$l���~��Y���Qz��a�.ڜ��t�C�kΔdF�'^�m`�q@y�̤��F�qW �Y1�+sM�*
����3l0���[���ͼ�/ٳ���wο>x���e�ڋ]s�c����K@���'v��쫊�x�1�v��~7_��������n�+�\r���h��.���x�3��De��{vKJ�F�u�.=Oc��9+��)|q���W"D������]��~�6@�����a�w��q >�J{/C(VL9�=����e�r��C�����jc�O��n��,W�/T
��Cor�*���wPȞQ�A���d�+��]&I��{���"~�����uqu�*y{�:\|2�&^��^�۟d�|���Sr����Gr�Ht��-ں����L�ī��Tw���6��ޒnsެ�vl�Oj3g8e�ݢ�����f�I��m*4������9�"��M�4�nd3G���DFX���<YX#Y���}��m�kX��XۮX�QY�Mm��i]CFan�m�:�8���ie[�%��xl�Ba�͇R4���I���:�<�\ڋ�ffq�`��`����5�=ʠ{C��j.�_'�K�"�kˣ�W��3��C"[9��?]��9�U�����+�m�wF밑�?^���JRn��~���Non�yν�����e۳r�3\����~�.��������~�e�GM�t�NKZ�>C,K�qO�;̹yN��5p�e���L�#�&���=��^�H_�`�	�y��?J��pL��ޭ��%������sD�we�.-X;:�K�����u��`5����fa���ӯ65MUB͜�u
HԳԮ�:�@��'����$n�&���u���`����;[Tl���*4��0��ܙHQ{p*����8��&���TT��Z�Dh��x9^�3����V{$`c<�Rc3c��C�Nߺ�h��}��eLZ}13¶ԹF�5]m����O&��NQ��N}���F�[#(�_�j�H�6yE��Iݝ�@��{��E�y����q���[�p}��g�� ����gCΉ��iű�ਵ�\a���b�MO13�w~��j��D;f|��+����&��n5ٟ5ظop�aY��=·	wm����N���6�d�q<�d���è�ǘP�%K7ӎuNɋ���[���c��g�4>ˮ����=�z�ǧ@�\��~v5�/,��6
m���FL( AN=�ew���
�r��.@�Xة��X0D9s[ 3���ݙu������Eδt	�+���Mw�<j�ga�Պ++[��C`��{o`�� �k84��gx�Ȝ��%fk�ꉇ���:�]����7�-Y�a���bzO�z�E�q��	hE����5�BpU1���^�+��,o�BU���`�N�ےůӞ�es=�R���{�!7��c�:��b� ��UC� H*�cyz��^��l�q�4�a����Ǡʎx�f�;3>�%U݆������̭��E�1O��M�W������d��Çcrb�u^Y��QO���E�չ"�«��Y�J7���U|��^~J�5E$�����D=����Fs�a�M�M}u��
��RdD���5'Uߨa���u��"��J��܉<k#�D�u��HB�%@�Bl��-�AHm�P
㓷�ԺGs��_��/ ����Ԅ����Z7Vv�ʽ�𞴅aj�-�ۮ��v�2��Fd����83����p+���eJ���&��P�!�l<Y��:�h�\�&xWm��nu,a�9t:��xz1���(t�Q�X:#x?]�[^��{�Z�ҏQꈵ��̬\T�O.QG��(tr\ݼ�Q��f�/kp�@�����7�?^��l�[���I(����4G��]���������Rף �n���s�g�;���.�Xs�2�%�B�;lځ�z����W����ھ�u�&_���7 �^��ܸWۘ+ݵ�/P1/�f31�ju�1�[6���.*�8�1�������!��vn "o3C�������a��Gcѹ�fq�~��f��*�t�/˕��ǹв�=�.�<U��t��<�5_��++\"n�n},���X�{�����ARd@ތ��"�|�pVB�Q���8}wE��v������ɻ.��K����K�X�\rۦ����1����z��ԡ��t�Чz�H��m{׃�o
q�n�|�!Wа?"�fD�66
	b�,�y�s�S�N�@����pQ[��6myz&{��e���h3��f�e�_ E�[
⃷{��� z��^��r��z;���6O�|q�����Ҟ�]��J),B��'y��q+�uy�����`�6��zk1M��3Ies#�������}t5�v���gy�uu���ڗw3���1TJok�푌��F}=�
/����X0P�]��F���g*���g{iXY
��0(�h��}�p�.��M?[Ϫ�i�K���#��0ȧ����WGȼ�F	DO^ga��f�eT���Ƞ�Ʋ�펼W#'�A5~V�v6:�*槨x�mH�����r)�8tU�u��6�u�����Fsp�������Z��t�N���VBٸ�����\)�Y5�;c�l��<m�n�J$��%B��펿Eh�D{H/ )������w&̎X��K�^w�MfbyJ�Gc0%k��
�V�u�ְ�;1��b΀�.�������l�f힊���h͐�];i������%ᕪ�ۈɻJ�<e�B�R3O��~;�@���U�n]<�tC�R	�0��;���Y�ASko��~��n�2?�ܐ�zÙ�ke#�j�潣�`Чn�����{�1�*XjN
~�׻��KP����9ӕ���R��Nbc<j��~�g�$���%Yb׷��^��xΨ��N�2pq�b�#F��ȝ�Nj����������~��o��H��0T8	����Z{�'n��a;ä���uou���]`�+�@��:=LsP����ۮ�Һ���v�D��NA\oF��¢j�̜�qۜު�eٙ�x�n�!|��c�閠0�	�?
t��n�M
3Zշ�#v�6�w
Pf����W2�աeL��	n�V]sp��h�^YkBݶ��6�T�I^Cj�,�xj�:�Vh*�c*�c(�����uq�4�3^�]I����#Տc�;o"Ng����O����V�lPH�C�����o���=p�p��姡o���l�����!�^ٰ*��/�;�>�4�;wj��g��}}W	���q�$6i͗"a?�E�v��}c\E�J/#lT�@�]M;�mwz���c��M���5����cҷ�t�޶�u��3�x���{<b�E�}.<��[B�`[�D�B�{G&�V�.��RQ)6��g$��&�A]X'�>7�:�K,k9��<������3���VHr~�}��l��)vFŏh|��oOppfAK�>2�-[!�M���E�ֹ���9���a^�4ٿ�gg{�f}��Td�}���3&Fϑ��JE�5�+ހZp��b��ح��'ds��#��
��[~���*�b#|N�4i�;�P�jn��s}2gw�W��׻�p��dmP�������CR4>���߭f��x��l���y�C�Q��=Y����n%9S��r��D������)ķk��fP��È���=��LD<�{R�t���,�u�b����dL��q���\��Nh��t��b�Y��a%Q�8���'Z�Y/$����Ug�����M6Ga�痂���V���R˩Q�+��>�[�5�i9#�������(�멇`�l�g{���s9Q�Mf=���`�5;]��Z�u��+ =��h��t0��0�D�U8g:�5�tG;�b��4B�H*CQ%7'~Îu�Q5 N�.�� �j`I[�R����`��7(!�_]�18��lvEͫ��C1�W�,@aPf��T�D���v���}��0��7��X��Y�$1:L��� Rc�8�j�^m<�Ƅ� p�2�����q��6#wSO�? �w �!��J��z��ﰰ���%�@i��g' �t��@��+��p^V��9�k���;��i�E��{Vw�� ��k"�����`p#	tՂ,EYP
T$�r�ۅ�'�z�9s�������}�0:�; ���j�z��=�qX{�ǥ�V�ȮzL�wY_YV�1k%���[�^�gج�Zr
	��N�m�
#E��#��AHɳ�Y���Mh0l��#R���m)������'`@�ܽ��`���!�2U#�l3;�b�9�%#�CX�>���x����[$m'��h�M��r��r��T+�/+[=�ۤ���Q����g���(nj�\2�7l��j�@���qfb��bjVMf��D���.-b��=��8+���t:w����9vå�R�V����3�)LcX�ؾ>ڑ�_]��Ł��H[�����.&�ێ��<�b�:(s���tph��k4@zP��4Y��;Imv�r��.:�3�?��{I�Ym����m��m��n/�s}�n��Y~ V���T���T�5�	,���=�a�c9/_��+���ޫ�s���Wٔ�+��n��t���W��w�K�'[p�9{�-�v���F��`Y�P�WW/*p9>����2�ҚQ�ǆ�NK3��Vl�`Ҳf����cA蛏�о���a��eM���ش��e`�~%�d}xv֛z�u������c�O�L�����#�Ulн4�����7{dv�|�e�tP��QK.�J��J�2���J�S���0')6����3����4̽�Ͼ�/h��{���� ��`/�aU�I��8��brN��1>�{ua<�;�k����6k��i���Y���;z�]4�D@�[k��d�ECL�f��@�T����̏R���wGv����s\n1q�ۯ��9̳'F`c]�Ewm�fE�>��^��Ż�ֹ�e�ְ��n�Ā�Й�ƺ�idÇA��w�r��I�e/�&����P3�gqˬ/o{�K�} t�&��VV9f���q�ʶ覆�\��5�)i��AKY+Z�t�6Ȍ���3��l��`�SB�Y�5�T�y���u�)��Vے���8�����ť5a�fѡt�ٸm�kU�j��Ye�LFD�)m��:
YNn%�-%�+���i6����&.uі�2�cep��,Գ	2+�T�]434X�H-9�Bj�^&�l�ά�J��[���j:�1ō�!,vre����^R��jVY�H�5β�1��5�I�5t���hʅ]�u$��Sk1Bc*����������m���{��jM�b��"�*���Rvk�o,����<���ton�f5�XT4#v�v�J��v�e̡ck�R ��V�ޜ�����ͧ��9Yo*e�۱��� eW�l)����)#�@��B������з���������K'z3�;���)�aW}]E�kjxd7/�э���!��cho����nm��m�O���f��A�L�7&�q�2/6k;�#u!�XK��lD�L��Ǻ.�6|�ַW�Z�>�[����|��j�2E�;[����T�x'��U@��f����/�]2��,B޷�z�6Z��:�	�"��g�����r� ������y�C�����|:l
|��t<�=��onhנ���I��� �KkO�u	*���{c}��������j��Ч���n��n�7��Nbb
��ѩ���Eo�C�͚��^�]�5���Qخ�ɓ�����3��,�oC��:����UP���c��;?�-����r��u]�q@(�WWml�꿄V����SGUF'+\�i�j�9�[�	�<�r�:������Lsamxx�q���5��?}gr���
�Lx�v<�K��	�s���Rh
���7��dz&�@2)��`�iC����"��(�9`^���T�\$���Ӄ3fpzHy�T�flTzq���ft������U2Vb6�-:��]f`��5�B9Ξ92m�mP]���e@�GHvv�-�!h���z%:2����ni�X�V��v�]�INص\UJ�<.eHSs�ȣ�〽#A���qD��WJ�����=�M>��fWk�"6�M�kb뉗�Q�[���3&�z�Ȋi���4�{�v�G'���.��|�fë�E�C�b�x�:�%�1�r!7Ab��"g��r�=������U�*{z�������	.�ez��"�o+<���ݦ�d�K3�wD^u���&��}YQVØ�s�W}�	�������Ȗ�^���7#�V�с�}����;#���-����2n�|��K�#I0��~
�z)��ޮ����v�m.���FƠ�ДoQr�͍�g�!*��m�8��ͷݲ�N����ټ˻�p�]� ��	�h�����GWw佯��\�6�6�(��pΕ��b�d~�U������'gdr*39@(����/z�s�38^'L��=��j��A7��y>�+0���UHZ�ݡ6;:�8y��E��tA�cQ~EG��4}/�~��C���&�wkV����a�LZ֛ Y��
��8�jY̚&�읪�Y��������N9/NV+uKQ�u�9�ó��"X�N9N�z�����Fm����)�W��Ք:��	/<Z��e�`�Y��GtMf�P�}Cx\�2��Z�z�7����19�ځ�����nb��S]��Z$)hm�3�e	I��H��}B{3���C�ͽ��Q^�
؟U�k�1��1����˱��37Gm��V=ɭ�g�.	�pw��;��v�����,`�����-�+����'���%X�Bچ<W�ɟ;��BP��z^�3�e��}�QU*= qS�l�@�#V!��i�U/^�� �w:F���ޑ)_ ����z�\Z%k�]��][�!�Mա����V3�<�A18\7R�T���˺36����)����72�\^Yҟp3]ܬc�^��GJcզ|�e�ZM��Wo�V��=<c�0����2Յ�#o��L���Pz�	��X�a]R�UóFzw^�&`\-�O���^�)r�\ouXG�cv�J�K� =ɬ��`laG:9T�i*���~7����ke;��h~�N���`{������*�ӝ8���k�N���w\��ZMLJl�y�+���G�{"���L�5;��a�U�%��s0�ʛ]�W8'��+�fƽ��!8�N�T���I��=L�)'ǧ��xy>3N�o{��\�Zp�[����r��ίU�ab»K�^Tc��1���Գ�4�΁y��J)��[K�x� �*�e--�˲Q�g��+�m�Y.�-�^U�����*��{���#�N۵^=M�YxW�����YJ'&1^�X����A�h��8.��8͛�l�z1�H���L;�]c�<��L!�}���N7�:����6�w�$黹�~L���g���Ȥdi΃~�#ǚ$L��w?xb��YM����w����Z���֦�EI"�>ᆎ�C�9�0����m/1��Ag.��c�<�}Q��L���r�~��VlpX�wȣd�u�X*F�1]�Pƾ��"td�[G/�k&ը5�*&�S��p��j�/�v���^k�I���z���pZ�%�*NL*��&�P�����9l�jc��IQ�S��o��"�6_:��^����\׎��	i�9#�Ml>�y�����W ����"�oAsǩt>��Q4咽n�Zrҵ��K�\���7%�1�j��Z�D����5V�w�iW��&����ٛ;r�xӾ���Z��k�p�H�J���7�=�!K�w�K�$�aN�XB���^O�˼��f�h�[m`V�*]a�d��mT��yV�Z/6̑�������V����t���!e��������O�K�䳂�Q�ɒ�[ݸ�)a\,�sc�;��p}G;��j�翽8v끂iJ�tB5�}sʞ�V�#5�ᢏ�z*+��A#=�����E��Ԛ��[�B����O�fG���ۿN�l>֞�[��'�YU���o~�"�{�{ϳG�S#|3$3ޫ��������8�������x2zcT��]�״@��ͨ�F��/���OM7�+7�������֭^�^��I�M�'tJ8(�o�s���S>�O�M���_?������Ȯ3{���8|���īݺ��y6�M�{�_�1a����i���Dn���}IlauI{�:�44L�-Z��3��VM%:~�=��gl���O�l1s�6�����\�^���=b5��}�� /n]�C�e���(s��D�I�k!�ˇH�h����O2�}.���j�_��`}AU�e;�����P�T��\X5�3p������Q�M�ڕ��̚%��E��k���\�ڑ�7��_߿C�K7(`��]~H�_$'�*~4vV����E�vj4��˥�ǁ�3�y&�5��U��0�%K��&㨺P�@X[�+�}���&�EJ�)�ޘ��� ���]K���s{�}�����Y�w�O�$p��7���yS4s�R��4N�D�J�逛YL҇�y=��o;Ū�ξ��qYM�+�K�ѵ�S���6�qװ$�?��k(|QX��:I�2�qe|�{y�C&�^����˚y����=��D����X=���G�a����C#�Ό4V��'���Fb�&��|5�_ӈv�$�`q1�dh��ww�7�M=�#����pr�Qq�;|�j8Q�҇Vf��7�Ρ8�ξ���W۫�sr;��Ox@��hF<m�����D�_=��4e*t��B�c�(x�F	�"�;�w�"�ǻZ��1�,MNۙ�P�f:�Y[Q>����~�dc�i(p�j��*a�)�LO}�j�YQ��'����m:*;B�%�+(P-����w��k�v���7���L`�>�;0k=M�w+1s��q���T��q�o<j���ך�@>�X�co�g�q��+о�~gP��P��JMF��>�'k
��g���vs�a\5���b����0o��V�5�a��6r�W�+HD~Ŏu��>[�k��L�<͡�x�s�7"y�1��wP��A�/��f=��3(�9�����2k�P!%[83�<�iNR��˻6�s���9mg�Si_.ᚙ���(�5ƕ���g��".ݚ#.��7P���؇g��9m��~��ѱ�_U
û�x���7�ڸ+Y�tI��i�@՟���躯 �0dZ��p��~K��̲�h�(^�PJ�iS�������u�j� ���)�1�^η��J�i?5%lJ2���^�ӎ�l%���`h[�rn�إ�n9�g�/ގ�|BeJB���4GJNuG�^^Ë���p��M�.$:ߝ���ی�Ѐ8I��n�;�ceb�������\S�T�u�T� Y�RE�@P�8�VɳL�	���|���}����=M��dO�-���J�����xxh�^/�z�Y�^��
j�l���C�S7t���s|����:��ev���΃�ڊ�u밺�=��gЕ���'ץ1ξ�{�gd�lF�9�0�I��.�I��+��yYU�݈��p^�"��GH��'k�"���u��P��:�^��������������]*R*9�k�ݐ�`G��"I���������s>0*�(�4E�cmd5�nN��(�v.�2m7��J;�+y��V�e*�:�S�w|C,�����	�w>��C�QWW�`�;N����(*v˽3]	9�y�Y	U��J����r06���~L YKY�� O�����lݯ��匮.f6/Y�[3KD�m�Ɖ���i�(�"j̒��Li�i)�5�M0�jqt�JG"Ѽ�TyR� k�nffffNL[-pWv��VVͿ�f�Ѕ������������ f
~g�#BJ�(�C�Y�'�chA�M�ph���!7G;��.�r����"�&2Nh�/�Uy��r�P�j�2�)Bɞ驼!�'�;�n�	�+eP:����`ѣ�&��^����!z�!����PvPvt�[.:���Ҁ���������}w]�q�>�����虮wb������μ���ﴋ�ǩ���n�~u�Dq����U+��/��ڍ,W�=K��3S�9���~0f����ϩ���f��yt-��4�.��̣9�z�^�c�)w{�ƍݚR��|U���_1-�»S3��K�ՊUR[�k&�I�!�����ay�;��pCK x^�n�O<W�ڶ6ց�;P$�Sɓ����e�ϻ}s�V�0̲*�]���L����>2q/o�����.��ߎA�:���K�*�}�t�v���ʍM�drǔ��!e��w��P˻�[L���M��)l΃s�F՘�� ��n�
����:ś�_ۤp-�яonH�x-37��V�rd�owY�����VݱR��3�j�
s�؂�9$��ܺ�"���v���/��9����P�8y<Yݲ���W��`�Yq��'�ѳ3�|+�+�v�MbS�����a/;e��m�����κ+Ml]� 3I]t����U{�+��)�Vw;�����-A����I�kGK��4��Y�=3ۚ'�����'ڑ�mD�5���}�]�lZ���3�{)��aҍ��RI	�����%�/f�	�5��xe�}1�-x��"}������?k�\R�@8S��c3��o�;x\�w����`�-�x����++j%�⌄K�+1�QN�H̶������F�Hmҟ%��4+ǔ+���^-���v�������y�,[�]�y��'�h�D&����y�ݽR��U�Żؚ�ԆOr-�k�U�sK�����~�Hs��T�Y�ʞr�mZ�c�>[�稝Xپ��S:�tv�C6h"��'c/W�B4�n}R˷]�Ҍ��0r�.]3�u��>~Y�jPU�/�g���{7{<P]���g����>�Cv����6(e��C�o�mX��tˢvLtŀ�:ef�9\Wx�]Q�	��J�6�G�r�}���#��
#^�v2���Ƨ'֭aT')��M�Ta<ecT�1��qrTӔ��Q�W�0^����=kU�4f�Ϳx==+׶0��ȟ	!�/��H��]��������d��"�7����Ű5@�o���}1���ǥ��2�*H鵶���L��.Ý�u�ei+j�:���U@���쳽u*0����������U���Q/���%N�g1	�z%��157�[ח��^� '����c�FI͎$���38�[%���6w�nl^[�[�(���*�8ɿ��5�]�e�Zk
\{�l\�:դ�I�޻�	�|�ڬ5N���	��vx�F/iv��Y�a��Q���R l��~�? [�_���ґ	�4�!ʔ9��Je\�6}ӑQ�!h��yV�ZdP�V��5���uGU5$ÖR�3���\��#Ұ�b�G��
�R��N����v�ڶ����)������Q0/t���z�X7�WZ�oa�����?nVR��̋��a��P�J���3�Es�"c�8�bf�����PZ^�b�^q����f�3B�{�KhlX�c���6jֈ鎴��:���p�<�fJ�u�o"�S۷+5��o.ԝ��3�"�*Uǫ\��}V�rv,Yš�ô[�#FV���l����1=��t��(�s'r���+��z�y:�%��2�R��E�D����
?h���^]X�8~�#<1P!�:H��A�H xG�b2��[��Y���ϓܫ�l�����,<jW�~�]�	�����<��3}��u(^��@�xVq0����<>H�����֎����_�tU�n��b���9#�{�.w"%'М"�	A]孃���
�u��f��Ӻ�-,=Q�.q���6�8�hɶ�1�HUs7k0��
 d�L��9>��+ ֹ_My�5�F �6>n&R�mH�Y)\����&����=}N�Y�Xv4t�>�Qr���@�R.�t:űG"\;33+�
%@���vNUww��%g~�o�i�>�����ݐ'Ldf9H�vmZ{�4n<:��1M#�*�y%�Vr�M��
���]`v�*�v��jr�	HP�N8�Y�MM&����!3��y���~�~˝a!�$�!� �`��������$BF���������a��6[m�Z7�X̺���松�����jI�N:������Kw���>?8���� &���YZ�}���{�HI�����|p�qG�^y߶���=���J�zE��8��-��F�w;�k@N�j�nP[�[/7v�P=��L+��ء��i����KͮYv�����K*p����)��!t�˖�g���
�q�,��\�#j:�j����Э�v�^�|�5��-�0�=P���o��=�I�]R�龾�o!ͻ=�F\��╨o[��;|�]�<�&v�9�u5�
3
Z��c��}�0�6pW1��.�D�g7C��G7��:r����e6�ҴA��ɮ�x��Ƿ��%��w9)�v��R�.�Gh�˼˦{(j��ޓN�r��IsT���2�$�Ǌ�J���Ǫm����}
G�vk����c �zU��9�WI^<�����;�l�ÓA~Kmw��뗝�U��o��_�[m���O����Y��A<�8�G��3s������eh��V��d��є���,�N�:�-����ٴ�hcެ��=1��.�2��1ov��HG>0�fZ���z����Yk�u�Wu�,�;����Ǘ"�i*��I5�U���ؕ�my�x�T˺ �\��W�r���D�2��3i��X���7�S���t�W��^����0��#�<���KG���� �b�m����|�e�=����ad-��&n�Gk"}d�4�3��bý7h�D�ݠ��$�f�O���55c�_����6:׺��^t����$Ȩ�ث>5��0�X������E{
]�zۑ���{��<�8�;����g�͟7j.&�eD��Jh�V��͈yp�"���������:61d��1\�0�.Q��|��@?Į��öy).��:X�GT���U�����q�������J��\'����2�%��f��"��1�h.@'LZ��~�Q3��]eI�6u��1(�=�l���]#Ʉ|5#іB��>����2y�\8=1FSֲ���m�EY܈2$j�����g�m�)�!����xӊb0�os�\���/lA�]b������9V3���u]��lO׬f����!��:��^�KA� ��<���#XĊ�8���`�d\�.UN�<�ߪz�%|�d*Pel#g�b(<��3���R��Wm�D�5��1M��^�)+4��~������a�N��!
90L7}��_�+���5qV� Z�����[g��Ԕ�mu�rՠ�5kn�}zK�)��4ضfkU������,�;+sn-�h85��)R�F���0C,v�3]n2s:ke�٬,.&��������8nfoT��F�iPf(^*�9W �|[���Ut7�Gգٱ����i��|�HO����o��g'�;��|���f���T1��~���!CCtI�0O]<�����ުz�O?	]�q%,B�9qJ0��oz���#˷����m�ئ�[/��n%���˵k�Cμ�Xp t�z{���>O�o���F��y��eN�U�q#ZfPU/'�eM>ɹ�75��5��.�[��P/O}�-//����JT���&�6AXj�����[���Z��A�z(=��k{��3?l�,ro�A�6�z�*CG���jW�L�O����U���C՜WI��uIN�aN�.����Ƚ�I�rE5��U��P��G`���7����<'��b6�E&+�?��1����;/�,��L'�3/�b�:��eMo�����>�z��n�����[��=��hX�~�Y��&�٧C$����	/����sEVǈ�z3=y�I�1�>��Aۖ��}�r�NDU��ni�Vֽ���2떊7ù#o�|1h��]�C����
|�9�ݸ��v�7��$+�"�Y b�Y����P(���z}��a�>���G��¸)2{�z2=9����
���+p��@ɷr�1�&\|�d��"D"�h��� ǽ\� �����w �Ǥ�(��W�םGѹ!+�����S�ҳM�O�����yC Q�껤�������� ��N�턓�@��~��U��j��`�P�Gm��R�h��e>��2�H=3��j���\��ez��\�y���̘Xa�ԯӢg�H{������uVN���.�q���d��#�~Q6�t�����9W�#���|7=�w~l�G¼�`Y�*��31>1 z9�����튭�=�B8u-~���U��fefY��f��-�E��*���R���~��՛ ^B��C�ƽ�L�="��6#��C��aN�D�����R�Ԫ�;�%����(���gs%e�v�
�j��kT��D^�$̺#V����Ĺ�ʵ��|�߷ήPr&5�5��v�W�n3�|�Ux9�.�����)���;.�́�%���X���}p�Ű��/n΋�˺�Q.z
������.�quU9Z7�`+H�	��2re�[�����-TރY:�=Ƹ5����F����y��.��B�3֎���ڛh������B��=��ǰ΋�ӻ�N��r�P���c�e&kdXOz�Υ.�)�>�y����x�@��-�̾��_w�f�^���Ln�=u+�^=�x�Řĩ��٬�.2lr�]y>+��f}���g��׫=H�v�C��u͒���|/���ˋ��l�.˚[���������mERh��(�V1u��y~֢��;5�֖�ݴH�|A�Ż��ݥc)X����vg�D��3!�xLԈ�t�����evQ�P�m�1Lz�c:+}��m��b�2�*7:������Q�B:}cL=Ѣf�۔����ݍ�w�{��ہ�9j\l��ߜ_��
if�E�F翯,��<���m�]76�B����P��3$�g����x�UCNPir��k���"��-B�z��( o��deXdڧ�����M�ϧ*�*4��-���s%׫�(v.a�k��Ǌ+2��Q[�9��B�4(W��'{�w��L�!��CeT]����)�c�H�ּ��~����YuxƎ{���I��������V�,���{S+Uܣ�4�3$�YV'Cp�5�����l����ϸ�Sx��˻�5au(8y�kz����ʊV�+p����	�^|o��c��n<���l����vL2�g� �y�:=�Hڽ"�@�$c�=p����ȳw5<+b]l�dB�&�,�f��]g�z�����j���UW��� ���4Ζl{�0ȝ�Nϭ"Մ��U�1�~q�\;����݌/>�Jy1�|��I?�s��u��H���W�4���]Y�B�>}Ξ�#W���9Yd���j��8!u��S�貳?����\W��4!�x|�a�a5�ZV:%*��l_���>�_�{�b�=���~
.Fm5��W-A۱;&���<_�k-T-�;���J;�u��[&��h\��H!l^)59��.�#k�XPkc)�Qd�.ؼ�z	x��sX�}!5o^H�y�ƈR.D%�(D�|�`S�^$l�؅÷[��HuX�G���{3�Soc�sE�]9z�����E�.��~E�Y#��^���Ą�ߊ��c,"��8M	+�����ʣ����>�7����Y��%���7��o	�&\9�-���ӝ/�/�`jf&Xf�J�RPF�qX)!pdۗ�-�,�p�̦C�p���[��c��fܤ�z�Ӣ�U�����#���쉜��$�o:?��xt؅���v�	��t3�y��<��*CM��f�[-�
'*��yBi�ᎺwNХ�%���:Ҫ��H����Z���T�����.���v��inkJ��m�ە8�w3n�my��w�����t�}�Ǆo��r#Ӹӳ�I�{��-z�/	�0՜3�K���m��s���(�Q��q���ƭ(�k*7!N�ت��.���u�羴�G�KO��8i��>?�3��+�\�7""`��Z��[p!���uC4��\^��{| (�!ÀD�c�`��ۡ.V�y��|}���G=�鬜�q�|ite�38~���R�:�x�ĩ�޾���m`�[��Φ�G�nd�Ϫ�B���υ �+�R�oX���Iיf^	��k�d�-+	�v��K/�K�#�Z�Ɂ��0�2����=���5�V̙����Q��WU@zEuɓqœ[z�!C -���a��2{��@��I���Ք�	�Y�'ܠ�T�c՜1��4��T�}sls3��N9�_m����L�)șm}W�`�����11�<K¸�į�p��0��f��I�; ��rFz��A������G��{���so#8w�I���ٟ��|V~�UV�T|6Ez�n>����B�p,�^J��&o��c�"e�ek7vy�S�I�S��A�5u>����滰V���x��D�/ ��p}A�866RU�.�N�&��SI��l��*�<bqS9��^R��hox1�@�/�>DD��1Ǵ��>�a�����͟)�h��![�t���e�l/�L ��=��n�H�ܪ���j7���n�{}3��ݡ�Bw�&�<@u�&��I֖��.5B������{���ǖM_pu�F��ww��r�{"-L{m��e���i=<=� �Q"og"i*£t��8�"t��ӭ�C���z��yR�yq�l\@"�{�nZ�q��/�r�|1i��93�f5w,�]�{��*6�^m(&a�\g�>b�K���k��6L ��	�5x5F��k�V�{�T��%T�v�RK�z1M�z�������5p~��6+S�9
=O��Z%}����c�:��F��=������@_��n.��|��u���ϵ�8�x���<+� �� �<�h�6���<z|@�ǀ���39��e�i� 0�Km�L�mŶ�X|��O;��/�4��.3>�����n��[R�
��=��ꎎƕ���"'S_���O���vxۆ�ܞ�ON ]д�7�mj��ubbZ��[�]h���|%�0v�M���s�=�GO-Vqf�������m�틮��g:��o,;mC��J�1W�40ć�1hL�ݛ��[�PM*�V����~�у����OS�;��n��b#E�;P~$Ўv]���u<4����y�jJ^�`$�9X���ݡ0(L�����*H�2�?�������#u
$�q�,�X�1Ogikb�z1qW�Q��p�\ǡe�J����S�����6�I��{�صW�*%H��e��Ȣ���ܼ���mp(��H��1<��nq{x�:��ϥ����H��6��ӂ�.;)@�������+=xͧ����=~��kk�켚���+��i�܎Ī� O+�%�� �����L�O��+<q��T�[@W��¾v}��L(*
��a� H$���&�Gbp<eP}f�,{�x/G��1�P���w�TWq����������еed�B ��ˈ�>}��=X����MOLX���9�\s_�}�a��`��0
1���)�dR��|J30�}r�NW��������(/����u���%빰v��%{�f-;F֍lUv�Eg'`\��{�G�w:қ�׷�)�m!%mj!�\>� �H��5P"�qs��N��w\�9䥰}��|��Hc�NX�G� �x(U������>�!	�m��D,$��^��S��t���z�EY"q����!��oOގ�q{���ׯ��`|�tO����.��<f���jE@�A�>�N�l�����ir� �@H�d�^��꺍ט�FЛ�=�~�������Z�qG}��֞դi�sK�%��c�
O,���N~���c{� ��X�#��tyw`��騤*�Ӣ.��8�����$4���&���T�E�hͥ�d@��BQW���o�_3�yF�<KBT�u���׭�l�^v��ޘnU�A��u�Nr�kB�83�q󅷚��0��jB�����3^66���5��)�	@��
0�l&g���ِh���dA�$jU����m�1h�H&b	�;�呣)ك�u;���LKu\&W9�碷�=�t�5h�L7ż<��P��ұ"c.�x��W��j��loz����A�F����n��p_u��t�ȫ��&� Ն^!�����cVfMËE��uX�ތ��L �Z���;���޸h�,��.;o3�p�v77r�]Γ���-s��罾������\��W�����Ɛ�2����xM���6(��*٭���[1�k���RP�<���w1�f�����ݱtn�W�%3���mu�˭ۗh1Į�Koe6�m�D���iO�4rr1�s�������B����{;\؏:�<Ef��y3��8a����<��-��V�#<�4V��Wi5㋳�&ޱ�$�J��g���sv���
��KNt�=��wP=U��4���$����eBN����i�������!O�Y���x�����Gm����kL�Yus][�p-CũW��,����DOmV�wa�~^6�|�ܻ���N[�g-	��[+��g7�8�`�O#Z��9iJ�5�>�I�t�1��zV����oJ�N�f�f�-�-r���^��_<^���H2��+��_��|�k��-���]�B�D4,X`l5쎅G�:=�7�4���'�.�@B5�􂟡�s�w���}_y������{ŋ��a��0G��z{��z/��`@�6��q�F�4�b���N��1��_��[�gKx���&������:�d\{��z�]{l�A��gC�K;�k����Z�~��ۭ8��{`gm�*���3RQ�z����LlIƝ-"fj�0��XV�z6Њ�����\�J,��MiТ���-!�8���&f�0�U�$�Z��Vf'�"�8��v`�U{|u�L���J��!�.��6�[u&o41��XCw/��e���]%�㊲�(�q��U�:�|�p;���!
�]L	H��N'�2H�J������pٜ�]���y�)0_6�%f� �z�H���u�)�al��]#�[k4+��U�4j>��8ѝ�ƕ����!���V��6ice�[k�����Wi�y���3�ړ�������v�V�@΃Ӛ��N��G��ΰ��O���|�|�sk�l����d�@5e;K�ˀ=�F�DV��l
w0Tϝ�N�uG8�����@���1U�P"ݠm�"Ճ�-�����Z+�Ve>�{1�k���|U��zJ�Ӧm��VL�[l�ݱ^�k:��fF����h�O��U
y3��$��V�K�qQ�`��x�m�O�uE��RvF+%]��Y7LY[vju�r�nY�Em����L,���y"��YZ��* f7u�]�F�����GdY�n�
�k
����W�[���i�Jx�g���rz�[d[���j����ZК\o�a���:�r���j��Z����AU�����f%�kVMJ`�Ct�Lԃ��jcTR����=��pƋ��9V�b�;E���=O����*�ٸ2
Ov�;{��5h���ӿg|�����Bɂ��t�⹄��U�M�"�C::��ȫ���b�+��ګ�,��N��X�i=�<x����\]�_x~�g�2
���AC*�ld&����/���R�+!hfMDp����w��:�[jJyG�j$鼬��-M��5�ں�;�P�qlw�&ⱒ��V�(#+���iu-Y����[��ˉ���NT�^����%����'w ��gFu7�s��cx�s��=&��m_>:�۹ӳ��V�Yb�X;��
��6���M跪��E��C��໦ �o4+�N��ݘ���(t Q�I<חǱn��T�b�E1����gh�ٟ*��lSS��jN�cR���e
��f�84�H*j%����'h���2`<�"L�P�A��!��������c<���,��v�lۓ�
��kϛx�SnKk[�3ɠ���hfX�we���><�;ݛsCYiF���Y�ۃ�l�X&qLۥ�r6�J���������u.�`�r���P�v���4��1��I�	�5�CQ�C��b�\�\���Զ6kt�ԖX���^fٷ�g^���f�RkS�N���v-k�7r���ܧ2��ŵڄGCH�n���u���͑�M��-�T�q��ɉ�BJ#[4L�˥�Xd�J�gMUB�5�k�ں��^��ѽ�)�w,.�	��\�#��4&q�L���V�DGq�Ļ`��'�ܪ�a�I�mf�2��j.�;SMs]L���hY�\�lXlgj2���El�Z:5A[fK�3��Ǧ�ť���&���u.��Hs[6[X3b֦�s�h�Қ���t�.3f��V��f�u�n9�%F��I��1�N����m+�چsl3n2���ķ8!�UUUUUUUU��m��g��W�JT�����ѹkٝ��'kR�US�7\��<fU���������%]܆s�/.M���o<8���x.�:fj����wC��=h=s�ӪD���ff`&z��pVS��HM�*�,{)�ᒃi%�,��g�_?ᒑ�5U�7�9ܴ��F���I��X��7y!�K/jml_H[<}��g�C�O��k�4�.V����&׎E��>%n�B��3ͻP"d�EUCЯۇ{��~[��N%��!Z��.A�5T�m��f���3�ާ�}���w�� �Dԡ�v(G�ڍ�x4u+̸#���J�BeR��pm�g�k�;štp�
�j��3�������$�3SdU�c���[[%��#�;=�O`�=i���}���R�����_�\���Q���}�"fBZFW��e�eu����L3�ef��כ&�Y��4t��y(H�U���@�|k�mif�L���@�o�)ǩ�Z�쇞�:�^�Ȫx�GcI�?h���x��a-:��WQ9Yu��͐wv���1�.1��j ��0� �"w��%;�}�-��Q]&\�(h����F����O|�y�'�K�����!��2�\j?W���;y�� �V��{�������}��,d��F���r���e�œ+vc�Vňo*��x�tH[�jWR�HfRS5]���2;D��aus�sS����.�h�Oh���N��bm�[�0%��L�����S�2e����ב�܇�7��!�b]��U�z*R�}w֌ �+���Y�=ޜ�W]��ꊦnX���
�o�d׼Ģ.��'b��+���p$L
�\4!��˵�k�/dO(�ۗ���Sd|�u�1�_/l��I����f{N�u3���=�r�A��C��c���03̒T^�Ut�R����EoN� q����X�o�@�j}��:y�s��Y�+�~�yU4;�QR:���#�Õ+����3�i��:��15Z�?;��js�g�U�SNx�k-��13z-9��xc]1urÆ]pav��>�"��������ex�:�H%j<=,S���/�Ց�!�1�,e��ջzZ�l���Ce���p�hC%��9~�.�<V�Dy���u*���͇�.=��`~�뮴����j`��Z�����d뾧����<=�A�k�i���*���NR��> �H�3�'��Y��£�M~��_9��q�[oP���z#/��F������۫��5��[q�=j�+v��P.��l����i�0学^�����"��,�a��츷���v��#:]mg^V]ݽj�cS��F����6�Jvi�g��IU��h�5��b�2Jtꌭ�T5g�w3��1��嚍�@��VE_c�1ǌ��&�EnlP�;���B���~?�3���x���3r��:�'퇬O���E�Dz�ق��i��\]gޕk��e>���N
(q�����+wpD'�9�ݦ��h�1������05�G�޼��x�G���(�Wo�V�ʟN�0��u�K����h9?�q�;P?I=���j�YR����B��S���7��[(.�֤�m�$nr����Q����uz��'U�Gյ��^�)�~�ԩ{�P:S�~)�֧����㍄�O���I��2,]����D�"eS"�w��Wzs�k}r�t3z3=�GɇqճV��|0��L"Ő��3˺~r�w�|).��t����إ�̻vohj���k������u��ٟSB��b���2���ꪺgOt�������nzi��̸�y|:ݦw��/:��*e֡���N�������=����¹^Q�՞�{45���4�7�岶�-��!Ù\���z����B�IQ�*�j'Ra$�mB�l[O��u�ՃZ/~*�
�S�E�<�1n���Gq�� R�F��Y����1���Φ��dF�3�丬�Ɂ��d�R\B��m�1���ꕸDtf�p����,5iY��T�g$iL��6�t�W����+P��N�~.�o�y<�U�JK8��>����K����7���L�4JG4��m�]�Tgg$ǌ��J2j��.�;����܃�c�\���I�;��o]Wc�I�oE��3��R����d�U�߆���<���Z�7~_7k��Mض�V���L�Px�(9�M]v䁤jF�/^��Dg�������̣���������˧��Z�?c6�h�2+g��b��&oP��~����*^gy^Mpn+�-���j��*�G_(2�l��}��j������ ���܏A}��S�J��+K{�v���f(�M�p;�7`]���]�(F���[}�v�\L�32EN����SЏ\{ua�VΫ�h�]�,��qIU��4�J&���~{h��>:dx�Y	�:lG`�eί��M�MߏH�N4�nť�(`[R��:�)��\U F:�������"�r�.�Ĥ��ʡ-�T;X�s%�_TR���r�:�[�-ئ��>F���3���p����1�yK(��pU���r6^S�w�Bo�bȍ���孏6M�*�eJck-�;��alNyu�]��Ԏ��x<��Efk\x˪�5hx��Q�qRLs��s �Tm�#��z!�@Wk|�2_�������=��i[|6�����فilL\6Ai�0�WY���]�-Q={,��Pw�D�Zr(�o �߁u����_�%1�4�6����r/#3�^Z��͝���ȼ'�a糲�6ߒi�,�
4�)����p��ţ����^�J�TN�cX(�^H�̨�~�Y�=Et���r�	�Rk*��6"�c]�U�#'b곡�>����f��TMU;P���N�r)�>�-)�x�n���$ŀm��ׁJF������wF�ìCw���Թ�n��H��Uy#8�{<��(w�粗�>��ڠLS,�2gE��o0E(�^�o��{�|�%tR����u��Dv��m�%[�a����y�7��^Ҽ	k����||�v-�!e��7/,c[y�4��Rr	�ukPZ�_;��rɃpY���兇41��@�6������튭0�s��Jf�un�[��)t��Q�9�mlJܡ%^��/�D����@J&k*>�#�{/t�zF���y:��}p�:V��� yf�$��=7���S���fr0�����=< �tpkNM݆ۛ�\[��V�5�ϕ��@Fyu�f������Ez=7���T+n�FP8j9&eC�;g�r�p������[�E�d�4��cf��^gr{�P�(`]���i��í��qz0�LY�<h�5Q}�6�X"_[٨��R踝�/�Z{�m���։s�����rkv�u����RX���N��,L��:|���{] zs���О�܀$ҙO��=�ie��+��i����`@���,�S�.�GA\1:tޥ���썕1��gh�P�!��2�{˼�n�H��Z�㢆��D-��x�����c��\cJ1���?T��#Qa*R<�f
L�Do��KC�����i�
m�G��L�O�3	0I�'��M7�B+5���K�ʨ�˕������`�gD^Bډ�����m{�n;H��(νcn�_k���jmA{'�ވ\���f�5�nܺͽ�Ս�p�\�(�Wng��ea[ה����ù(M�ђQ�>�zУ��Q�tϱ�WJ�m����>Qn9�F�G!a�QX�D݇|���V�IQ�W��{�Rͬ�2ĳW���
�1<�O��ҭ�}�h�N�[:��H�S��/C�]����p�)���(��*��	�����dC�޿����0*���&aKB�h�~Թ~��UUS���ck1���?s��ީkG��}�rP��}�=���:KUR޹�(GR�@��CGL��]>����ɸd���7�,�����pǺnt�1;kk�}'l�Ǻ2�z�A�Z{�g.�i隞��k�f�Z����'��ق3�}�J�b5w�/%�K���mT5��+7�z�5	K�j(P���~bTc�B}��j+,��Α�VY�ƫ�Y��\�s!Yӵ���N'��G=;g�$����w���VL*Pڢ�隅W|)����O{-��}��ո���S��ڽ�����w�|4�B!<Sj����J�F_��>�</�5�މ�0��dC��^���?32����'�'���0ҏ("6���^�O1���MB�7wS��rTy���s���o�syr4z��}������{�ۢk�*�z��/S�!Ʃv��F��x{n�줍�����"�B�=���l�*]������0fERqqIr��s׼���1k�	�1��I��\�A�Fv������0�r�wR��Wu����^���u콖n�n�R��j�УlJd�u\��N��K��dm��6M��敛�����i�e���f8(ƌl���B�s�8η,�D*#r�܏ˮ���u�mjmm����8�#5�PMC��ʟ{|�k�n����P;u��M����;�X
�����NH���АD��ۣ�[T�b�c�����C��}Zڪ��>י^�Ȱ�o�L��UM̍�	��a��<��
��E7�ϫOT�R#o0��������wb��ߏ��k�&x��t~��<k�4�	�<.m�k�,��2�H.����ce�G5�K���u�P.���z׉���*jӚ�z�_����`G��΅��V�D���չ7�.�Q�:��1!�*�Eᨬ��Y�K���]$�TW�.Ts87�(.m��\q�qJ����J�^	��4�㽗�4'i��6"{ۗ��x�E� ʧ���|{|��1�V(I���IF�Uo�-�0ٛ�ꄰ�E��3�24e>�V�vX�ׇ$u�@����o�ZQ~ޓ7�j�k�MG�n��t;�����+���=ّp�����g��Xǎ�*����
^�P�j�4/#4�� M�oW�)��3!�μ���w%�r���[�A�G�1��3+m�N4���E]��Jx�ʜ[%�W!�	~��q�ƍoWoӇW]���L׹�X⯌
l�$��9gr��v�K������"?���nה�����s�!���l��.��9�w�E�9����v۱ x���� k�����j�?
x!,+�wO̃�n�}�������y��5������]�M��O��N�> qY�ƭ�~�e@8zJ�ߧv��ȡ!z*��+�̬w��<Yy|LxU��k���u�#'ʄD%bO`���j�*R�Wk\<���f�3���d�6p�>zW���/��@��ׇ	�[z��W�/��+�"�1��բ�}&.��枽KM��ռ3l�q��.V!������ٟ!�!ފvb�zױ������R��,ʆ2bD�Qک�.�J6�!7�!C!vr
ɕ��k����\\4s�譧��[6e�1PR�������n��MQ�N���.��}"I^����@3/"=�^N�z�,�E���y��>�P�����/��חk�{-���i�m$���*��¦�<�=w�5�h�)�|TU5=w��Ά�Ӹ�;�nm���u�[������:W��&�儅ɡ�G����]6�Fc��VB�m���NX������ ��	�(P�U(#y͢3� �����6��jH��v�}�6�����G!X��ً�
�Uf"�2Ь���2�u�a��̌��ޤ�Ux��_W�n�R�����X�\Fa��˿9��;�n��.0F�d��n��ư��G�J3�99\�̉��;��۪=z6R=̙������EKåT�������]׻Tl��\��
N�}	��?�M�rR`�nTc+�mv�zFuƕoB�!��{��D�}����H]1��[xpQ*)L+��A��Mh�5�ų��j�Ge��J�L�=����Q딽�k�١�Q��鉋�C��=Y��}i��}�;�A�(�].gr�X�"F)�&���(�EIH���+v�-�e߶>��U�1���J��^�����97$�;�/9�����1o�����{��'%��B�j���O� ���E��~����u��Ka1�պ��37��yw�^Qk��k�?g����ه�-#]J��Ș'��}��5���r��%�?y��l<�M3���<�'�'��@*�0%�	������K<c��U15wMWi�O��5�=ժ7������.>6!�n�l]4e�bi��3*��ϡ�,v��7;@��%�id�T�}�p[��cݣ�CP���:��Y��zdY�i��
�j��^�1d_!�;N���M>H��{�U��(l�y�}˨�
��a�/in�{-��@Rm^^-7Pr응���c��U��;�2��x3VK��V��-�"�QTXa�I�}]�^ܫ��˹�NЗP*UX(����)��0�+��.��j����,�@����`|'I�Ǒ���]o���3���s 5���y�w]
�|�j`Sy}|�>�˚VIv�K✵.��D�0��V�V�܉gf��kf��nݤ�"�53��](tfYn����2�e�^�َE�x���S.Y�F�ޜqc2�P�v�*�e���ύ�XCE��
G\���4s;te:c3����6���� �S�F�줵��C�7��G��/T��ɘgz,��]��G]%�b=]��\�5���ݲ��,�ۼ�e;�O9+��G@����$t�9!�e���V�z���<l^��Ek�N�)QM���� ����ٻf\[Vh�g)^�j�|K�/���(l՗)�yM�w�v΅�k�s�:>��v�˻�F6hj����C��c��M8��/�cth�1���5>�sw���e��O=9+;fv��=p�uu��p[;ՐܬYկ�.P�uCsE�6���h��6�9qܥ�D3$}�:t[g �;l�f�D��u��ԝu��Ƿ]��ջ�Z��7��6bI�<t�pїQ⭽�&�'���#:u�����ˤpY�\����(q|��AQ��U���S0N�_Q]�Vj��j�2%�::�2M�xe�xT|�O�p-w�a:���(š�tȤĴ��o[2����슺��]�V��vپ���򵷛�ȵb�ge�6�3�{#1�$;�׫�+su�^NPs�Ւ�˫��6@�va��qP��@izr��fu��I��j�`���>U$�v��}����u�hNl��.l���
��KDH�0�nc_/{&��p|����T���SlHu��G�
����46���\7���)H�^K�����u�kׇ�xQ�#;�u	�l5S�iE ��v�َ�����Џs� �`���6�K������?�_n��7S>g2��7��S��u�����p��ׅ������c��yjKt��s�;���+�}QܶP�!�ya�����<�^��Kʮ*a��6�Tt����P[�`!5~����4=ޞ�UN�L�9i�����?B8yk$ʑZ��9c;vryo%W[�F�W��o���=����F�ņ�[a��E�h��/��]�4n~#��~�S�|���w�??�w�yYF�s/)�Al.^�~��4!=�(��^�`������ٿ{/m[�;�2#wݹ����3��v�Ҽ���{=�x^P�OWk���[�Su~Kaü��K�]Q��M�������������M�U=q���Ob�(#S�a�a��"��آ)H�/T����'�wsR^�Zq��pvZ�r���Q��'f*y�h׺k&+�CH�|�oh]�������b;�Q��U��Y��ʄ�=p��_`=s;�)��2F�s�Y��wP��)leѭ���+"��2Q�i�(H%
]k��f�Y�N����T��:\�ͮ��mKH�B�{ާY��qt�D�
a*��yi��ir��#���8F��#rr�cj�mj�m(���Mh�NckjGis�\eU}����Ȣ�V1u�'tL����1�t��~�!�_�e�W�N���#G���q��/��g������'�7��O�랹m`#�#WFk�D�%��൲Ev޸�{ހ�+��3�-1�J���2v#z�޴���Xy�A���T��
�X�Й		"
a͡2�f"j��,��Ϟ��v��y<rO�5sc��S�3S�"ź2jL���n9���Qǆ���H"V๖<3���ا�EA�rZ\�,�.W��{�?y�e��k����������5{� L&�^V�z1_y\���u�8��+�{�������]�v\��J�[c#ئ�
��3|�MF�����4^���ю�QeJAR~0w��k����a�Z���q���v����L��ir���f���*��X��A�e"ȼ�ˌ�Q�:!�ب��	�ZΏO`U< ,1�s^��G�T�K�J�L�Y�G��8���/��d��@��]�D;Qk���K��E�=4�ub�}��@�*ʨ+k;T`��2����6���7%��S�`u��ui]i��u��^�=1��}�;V�e��D��vI]y��s��z(>*�ʸW���iNa>�G���ă����k�v����2��'Dq��WFhӕ�T�C���"O���4+��L��y�u�w��>��������Z������jZ�ivaV���Y~�����	�+�ɇ>�2�Z۝v��W��;��DOA���)Bo��yvG�D�Y�4�Gq�$H�qw���C��*^�R�QB�>��1���w����uaFv����L�9@�9r��ήf�*\��&(�(ڵQď^-�=QهE냢y���q�[�[���:����>A�)`'���<j�9$Э� nv4QR(��&��'�piGg�zx��P������8 g�1�Y���X�-�5J�Z��R���"�/՜���Z��VY��VỈ$��:�3j�p��8��}��8�2 XV����/
҆�U�j�ڟ���+�hŚ%��Qg��
�MI�"��۹ޣ�J�pAjflVE�=,��lJZ0�q��:v|��c��<���H�Ǔ��S�Oz����j4tj�w8�����p���3]m��R�6��m����b���ץ�R(j�����I���7q�T�]ۃ����Ǣ���ݪ�N�A~P��F���P�Y}��ݬ��� _p�@�{�`k>nC��J�^n��\�6��{{�E=���D� u;8����t������ewi�Cj�}�_V[S���[KZ5�얻���^z�f&��*qV�։�k#�F����e!�r�B`/�Ӎ|���}6�#��e%�ǔyMs�K�]`��ϫ�P;b�s���{�����Lƨ���Q�d\5m1h��=�q����y�3"��'t(�I��.{�?�c8�z�m)��hأ���%섎yHr^�W�p��FcÑ�U呪22�U�?gXw��h�H��l���X�VkΔ��vT��@���4���W%��zhQE�I�2w�"O�5����;1��|c�J)%���sg&���Wճ���Ί����s�G�$w*�ǈts�ޅa<�{��k��s�I��v>وq��mș.�XV�_�~��k����W�Ja���>�A]Q�AS�^�hu�af%>C�K��L��ʆ �8
-�B	�L��A Ni�+ml�%"�;Ü^ә}��J���k����c�tلP���-A�:R'"`��.��X���4+HT�\؜�O� 0A�sCx� ʏ\W�E5�ֶ.p�vġ�@xsgm�5�=:�AHi��5 �\z�h8�Q��G3w�[��B�K�4|9m��q�#l�,3�C�*`<�b�n*Vjm&t�A[0�y�	i�LɌK�����OZ�Pߕg^����%w`����bk#~�|v�wU��G&����� �V�q^�7#k*o
�?h����FI���{}&vm%���t�^�;A4����-�[7��S��P�|��"㙴���h�l��(#��
8r�ķ�Nu���n����"+�*�T3Q�1bt uT*�:Mgg������T����"I�6�G�ِc�a�
Dt{���1%�FO?`�_��E�v4� �7/�Q���y�jO����.�l�9A�i���J*�&�Ԭ���	熒|������J��P�h�e�6hnf<���L�
���ۂ�0*��F��Z�H�g�N<�J5�90W��v�O��B����z�f��8 (>ͮ��V��xBqX|�v�N�L�d�)��L�&�9Yn�+�z)H�J�~��Fg�z7�F���d��4��KH�Κ�g��7��K�Wvމ�]V��z��D��_3�Ё��-N5oz��GyL�fI�� 3j�T�lx�����w���]f��q���F/E=��9V]�1<�Q�Tc�Uu��r��.t����W��	�Y��pQ�TM����u� F�s���sI��c�b��FQ�=�N��a��*B[T����vM�|�1��[ԃ"oD�J��]�Z@�C�N��wOU�ZKvvT|͛y�m�ZB��]���q�DΣ�(�,!��Í�;(�K�. GR��&v���ï1s�\K��^U[+���3�/aӛ%����Km�.�$ۭ�v�P�cX��6[�Ch�L]-1w4a�b]�*��������jmA�%������%�{�(�JI�����p�"��貅j���,��)�":������kW�8�0���L�@�*�b7���oWuRčc��d�W��^�tF�s�LJz2N�"�{k�;Jk�h'�3~��R��vT�����B�8����2��b������Y#��~ZE�9ٮ��B��p�( �dN:�CY��[��o�������&��锔��s��Gv\)j��X!�.q�#�;��]��ڡ[C-n�}{��{d5�,z���� :	���P��*��ԥ��H��C*G���
z���PW�Hg8Ɵ��wam��Q�� ^D��ew�cm�nƛ�ޕF��h�橁ڮ+Vm�����F�t6 )��Ш�J��q��e�c�ON����4����`�p�l�g��ô�;SXvg͹�:x��+�0�냐��b�g��dcV&l7OuO��^�=�_$���S�)��C/o��;�Fs[Ǖ,�S���r�&<ź������S�zDt���YpbZ�i��x6�Z|�z�N�"�R�Mh3������>-W���w��@Η@෭;�$H��Qw��k����D������j�an����ءʝg�9�m�ih�P���-&qf���o8��4�U���n.�F�'G���^�����p�Ewv�#T�oVOܳӧ|}���W�e��=��m�3޳��Bȗ,R�%c�k�Fh���q-�`I3\.f"a��3��4˭��#-ͽ�?�����G*���	���o�g��T��m�K����A�
x���x��5=E��I9�i��ZN����}>)�4wum4bA��f�.���3��4�ϞH��u���.�^a��	�P@���mĭ���b�J�����-�~������(���g��6D�q�����:����Y��4�
�)�3@��n�]��N��*	F�:*��W2'z�]�[WT[>�a񓞶�*���,�����0�YGDuU7s+�i��e��0��UG�GM��S��G��3�#;��\�A�U�R��"�����S���Y0�����냧!�&�9��s�.d�/�����O��l�X�+�a^����TKM�����e%V���^���n��בQ�CȽZ�Ԧ��7�v�z��sY�<�AG��*}C�W�W�c��\1>�/�1g����YW	',0�i�دX5E��3��<��[P�ښ�q�S=��xp��WÜ����.
���m8��ڄua�H�E�\ؖ�8R��ek��,[噢����\�hZ���W�)�M����ǭ��,�e�������3�b��m��ݜS���[Fܹ�
��g$/�eL�=&tN�;�,Q�xVE.��t��D�CB]vXfD(���|������V����B�Nc�w9ߏ�ϥ��_��a�dז��Ua۽��~�ė������6]?�T�C�V]�l�bG��A+=����3Ɏ�.���
=����m�V�i
��F�ј:`$i@�����b�'�_�Ez=ëE�$#u<P&fA!+\��
I�0��wb
�/��Im/Mֺiy�Vsɪ���T��k�	�ΐ�6*��ޏ):�eS��g���9T�{� ��*�t<�̢ڽ��Q<�3�<ă���_^AW�lF���N����U.�Ma�D��@q��zt�׷c��Bi���X���;�p`DJV	�{d��{�G����T,<t�zc�U�w*r���lPH DYL%�I��.h�� e�IΞ0��Ʃ�3`��'�oJ���_��_�:&�B_�g����G6d�Q�jC��[��o��q�A9�������aq�01��]�@J��Gܼ�P8t2%����q�2��������Ծ1�sf��*�JW��nt�1G����}�c0=B����P�Γ�u]^��-�2�GbO��[�r2|T��o��]��"��Z������tA���Vd8��7�o�B�廙��idۮ{Fj���t�Cp�g&!���(��S�� N�k'�������9T��2��<��dc�BO�R8�C|�oW�B��(NVJ9�R቏?NE��l��8~w�K���>ғJ�A�
��np�>�e����m�	�}B��ٷ��ߓd��[K��ɞ4�w��ą�����������%��7�ќ�Ø)����n��>�YC�����'~bn�#�SWn���#lH�G��yj���X�G.�����MG�9�Ծ#<��9�l�EKsq ���2��4D�~�^������ ���1YN��9RPF<�lŹ�6)�]��n��>�sV@"�,�r<z�7�X�ZVKV[�P��Nf�@ڜg�؇5>$�ǜ�ɼgq�L:#�1�A#�쉺�S�h5����1,�3s��l��9o~6V�_��U'�ۧ}/c�}T9ȫ6�[���|r�V�_EJb����b�T?Rw
]E���t�O�D���-�f�hm#�fu�"A�A���s�"�Ș����7AX�#����S��q����]u"Ӟ�nzJ�����`A<��[/ª���|��"xx�:t�\�x�eI�o��\�o3;�y�5�Q��r�jʺއd¯v�=��X��S���RX�ݱF>Y��%��O�٧&s䫒�C�fT\��k
���3��\\t��U�#��3z�Ž��"�a�8p��[���y�<��ۍ*6�\(�2nQ���iI�-�(��\�BS\���,`�����N��c&����\�%e,c1T��
����i�%31b�6*��\i`U�UU�;1G%%>;��sw'�n����� �0�p�p&w�͌D�ͼjOe�W|���G�g�A��9>ܜq
�'��wC�橯VT�2�1��3�ϓn�s��C��YN�3��٘�]���`7�9�s|C��:J�W&o��q� _��U�]�w�m(y� ٜj4��#��μ������aG`�Ry[Xx��Ye�uJ�V�2�p"�/[S.Gx��2�$�s:!�*�K]=�A������u�nTk�˿<N�/{x_�b��4�D��'s�ˮV�ث!/t���,�U�Y�q7!D鳬����0}��G�ٙ؁�Π��s������˂O��ω9[B�pR�'�B��޽ɸ�tɡS�BGr�����tG{�E�N':r(�~\6�U�������7/�"S��KH`�!�*�^�혚D�燗Y9��j���m������W� ��m��#E�����yU��nk�ֺ�@�U,�V2j�ňa����ɦ�;�Rm9���l�>�-�vx��T����D��-�ې�<(N���Wf�Clo��M�a��#'���ɨ�Y�rU���
n�����bF�8�(~�Đ��:nj��IjV�w.���d�����Hv�.�w�����D�3�HX�IaF��Ÿ:�C���n萓�}Q���f&�no�W'YK�dި����:�~�]�v˶:�^X}Y;��j���05�mr����մ(;���c2��E�ݺ�c�W\�T���+V�5�H%f�(��]w�x�8��خcs+�@�GW6�>چ�(4L�+mAҭ�W8��A�d�K��fL���#V9�ܽ�|��f�ݚˢk���������H��!ݛ{�����eW�ܳ1�f/$q7���.�}���!�c�O������e1hս92Vk�XLW�	�y[̴�u�F��\�9kB�OY��q�o�H�kvv)��3i��,y:��=xnht�����J��ətO��9faP�>�0" k,g��ï`��$�����p*�,��ԴQ�e#ʢ��XC��4bіI.<��9�mRԦ��V^a��iHB��r��Ķ��f�T��n�C���l�n��X{��y�*ټ-�2���PP�Zj�&���Э�����_;x�>Y��ɐY�:p:9��f�Փ�1,�J���b�Wݛn��8�ͧpa���b�E`ei���ʴ�.���#|�h&����O
֫XM bT�E�?>�(wuM��t�ԙ��/	g�����P��^��h|*�1�f�m�ݣz�]wMx`��]�R��'@�wu,��BgV
�V��{']쫄p	�ذT��+]Tnv��\����wb�>�*Ͳ��9T~A�$�.�bGzOsZV�su��r�6%�x�ܧv���^�,��ю/r���N{�{7��x��s'ʙ�ǹq\.)�����Y|ְ��
�q�cqF��������BÁNPMn�"�H�]-�*3Z��h�W��ԇ0�+��P���ִa�uzss�3��ޟiÁjv�)�7i��������T�v����N��.�Z�BVK�ˮ�ER���3��bhR�f���3`���T<%C.eHp�J�e>%��,�jaP)�E�(G����(j��{���-!+�������W��.����+�1��<ә˾8.��~Q�M���.v��^S7N8pP4֖�.]rM��<�[�]e�l?.����(F�R��w+��%�v�[�^R��q���fF7x�u���]��W�k�1�,��Z|en�{������r�ʔ�T5X�֙�k-���R�U%�v:b���P���xK�Z��߄/w�f�3Lط�I���K1ku�]t
�m�.]c�ml6�F˰�)T��]��(*��ku �_��û*J:�.�Ɨ\r�k+�5-�fɫ�.#Em���ss��-�샶 ���Z�C��M5K��,��f�K+f�&x��H�$����cCg]~9ot�q��l���i���C]�"�kt���I�@&H&IL:$B��l	�a���R�CLJ6��m�ʰ�1��\�D�����B��\��(��R���+4 me��4`nA�&�'º�s�긥���.�f���b�[Bi��h&��UUUUUUUUUUUs/dۨ�.���)�(r��j��{+]����v���ѕ��d۵���j��T��C&�(��LY���I��b�[r��Gr�>�b�JCU�F�7j]��� � R��u9т/�Ud���u�#&�]�\�׮��O	�E�ܩ��Ld���2I_��6�{<w�$�D��x�Qq��㹟w'�@�S��Ѳ��pH��|���>p���(��K	p-*&��ՍP�������Ǫ|��� �%х|�S��x}-c]��s�~!�	�Bо�U0�T���뾬�lOX7��~ۧ��g�@�Q)����t*�V�����2�{=�2-�u(G���J�9�\�h��C����8�qs�uj�(�>:�+cD�u0�����G�4�ʠ��x�n��K��תCxe�=��W��$�;cԗ��<�7��k�5(����%�&{ʈW���H�]Uv(�_�f�t�M�.���uU"�ˑ)ӛ���qZ�S�;�Ȧ|�O&�t*��MWVMn$M�2�HRb=��\�
�����u���_njχ�10�ݘSU�J�]J0���2�W��f�BP�j�A��T_�,_C��g���w7=鈴�E�U�@*.��l\����VV��Uw�܃�'�{�3]�T4�=��;�cjB]=�LЭhf����vf�:x�Ő@wC/����;�-�o}���j��oE:ӻ��������6�2�k
��nI(NM�P��=�\��ިCj.>�y|���YHS�=k�ݥ�b�1���Lv��[J�z�Dr�Տ�JP�4Nn����m^t䗢���iV��y�+C�3]�������wgq����ܛ�IҦ�dX�oS����e̺{[���l8 �;O�~��S!�tx����VFҭP���Ҙ�As:�����Zu�SA�_��F����߄�Da��ó�mO��n���uz��'W/Bw{���!�6@2(`4)]GX϶P{��s/.杨|<�)A���%�kU'D��J9��6�Y�	�6f�Jz�_z��5��ӝiWa���1ZH��9
����$�9��A����P�@�5L���qO��oe�Z�����=��*y)�{�5�˾p���cQ�tTq��<^�>	4��u6�/G���
}'��I��2���ȃr��*Q�ԥ�
��Փ�g�{��̪}`����>��t	x�A���J;�N9����Q�*@Xjڝ6����0��t�ohǑ:n�A�Дȗ���vnf���{�{��m+��X֌�̰����h�у-��ѷBxA��Q����V@��m�L�~��*�\�& �^[���)ۓ���h+X�c�՛�w0��K#�'�)�&������|	x΍т6</�wx�U���WsS\���A�����[���f�K���<�Uu�:�bpB��D�r[1Ca(K6�콨�A�W���b�Ѐ��sEuJ^���B��)zE^��r2�wd�U�n��V^�d�7:����{t�������m�!�.�}]�J�`�JF�#�-���d��m����nu9z՛��HƸܾ3G_V��;���Y��D�����":\w��C:�Uh�!u��Mr�N<���Q�>!w��"�m��7�
s�������҇6�&t�;~
�Hf�_P##+9��{%d%��5�R�d�lyV��qN�Q�-J�<4�x(�Ɲ#M\X�׭�A���܇��u��y
/��B^�a���U�r/������܌�&���w�>�I1�,�L+T��Q��` r��[^Pwj�k�ґ�i�wk�����ˎ�b�U`OگۺX�h鋷G����
=�
J��V�!��G�8�&{}�~Y��<VE�e�11x"�RZ�*�V��c��>1YW4�2,f�sVs��zV�����SU�l�]�yh|5#�{#]��)������%.r�4����B����=��#��XH'm@����F���藹aI��]7^N�YNyr���f>�}*n�-��UX�w֋`|Zj�8U�[#/�D��z\�M+��Xd��!�F���_'� ͟E��ݡ^���;3[׵�����P�pM
�n�TR��5çܤFBw�+�_!��v����"�����;�(�{W����>,d�j�z�(�Q{�t�}�J��VU_OM��U�LËR�W�2�����n������<�\0�'�u�`�j��<[k7(V��řD͹�D��vX��Ǻ�N+�2���!��������_mۣ;�8�ބ��aފ9�}��ػqR#@�s�f�q�Ye�ff���n#�eI]hC[pY�kX�4�TL��-��.��);3b�klݱ(�ιk�h��$�L+��Q�%����6�9��͵Mh�|�|�02[m���k��e�ǽ��B*ã��e�g��Ƨ\��W��,�t;��ѡzх��{���n�O�uÍ�R�
���ӓ��2I�3���P��To���HF�p駨�6zr7	Nx(a�bJjvn��a0�����G�d�8��Rq���g)�C��C���D��S�P6S��ȧ��V���~{�o��kJ�[�3 ͡l�0T"a�i�!�g��0�H޲2�������ȸZX�6M�bV���-�q�� n�(w|�8�Yo�wG��)V��C�(Z��R��J[���"s����eҷ�E�Қ�6N�xTQN��t��G�~k s2 �jm��[���n���o)��'��u�T��%�ns4����2$��%oΧB��]�p�{����6�<�Ӈ	g����b��u=��|	�1Њms5|t���|�\��p;�1��;t��#u>-�RzJ�q�\g��~�'�� q�y�S�2�s`������'�E��z�6�{l<G+;�MP8�y]K��q�8T+r�P"�����I�lNA�{��r�os����P�v:�%-��OH
����q����(ɧ�'D�����c�j��XA��z�j��΂Fj<������|6�i['��c�9Q@Za�"�A�u:y��Qq�eX0�2[�(;p��&�bްqi�7���vo�U[m.�;��d�e�8hl��8&4��ꪗ�=�k�4�ь"8p�@���n��0�VK��zzoщ5���¼ZU�F])l�0�]�Ì�c8;ܮ'��뜉~ꚢ:D#b��st�q�>ѣ��F
��'�W�
5����,���{�:����!jކ��Q�uƞ�"�DC�{R�)�4r��/ߚ����mƨ��;f�i^i�s�4��D���Ad�C�P7��x7���P�&�(�r�#񇘄Ӿ� ���ϸ�0v�i>��b���h�X��,��]��J��)�8�k���1+�m�u�x���=`��;��Kܳ�Z$U�ԡ)Zg+�L{���I�4cYk��2�����J����ͤ���v �u��>T3�
���P7l�v/���{)�;#�B���gg��A�r�t6T�D���$:1>)u�["�`27gWi����y⧁_j�{٪
O��]��^��a���6�(jQ�>~ٗi��Ī;�⋇����lN"����:;���'��!�����3[�n,�\�Q�vvD e���i��\�ca��eಧ~x�<;�d���9Ze��W���괼�x���Ϛ e]%�Jk�H��1 C
=�#��"�� �k#�� lg^�s�K�ga�f�ڻC� t�}�/�Q�="x!��pܴ�ep�w5����gW))��s���n��Q
�y�.���4�e���Y+|�Uq���9��}�Cj�vf�V�߾¢o_�ye{sΑ�l� /��H�#�kY&�v�I%�������	3�m׆Nn���ʱi����2=�Sp��ӏ��ZrZ�d�$��}@��:+��)��j��&<x�nrCРl�SY���W�JЌ�U"�%�v�`��.V��r 쫌b�E�ܥ����/L���ڥ��rE3�yY�t���^-���}_WS�����[CE��C6/fuϪ��.�@��dԣE
��#}IUXV�)�c�C�����Hn���Ga���Ńk�������.�og��.S�K����n�P�tõ�;,m��S�Mh�w�T�s�r�����;��Qa�_6�?4�E0�0Z��.����GS��?��B�X�.R�䪗�'�.���9�����0p�d�7qLKQË/p{ԝ�h�j��,1Ẋxv$�0$�;�?Q�K��}��2�k3�N81�=���J�h�V���[�v�҂{��;�\�UY�#����r�P����vj�����M#��9;3��{]����"���pr#+��)p@�t.�ӽ0A\�����3F�Mb���Z��B�M����nbW��]B��-��p�m-����m:���+�����1Y�ę�HW���~|������컕$��{��%��VM�=� p/շ6:�Z;�Dy2��Z��/�F�6䜿zj��x6�DF�(����f�tR\,�6��Y]�-�R99۫�>�T�ϣ��+O�}�v띊�m-�Ln{3/�o,��v+�L���դmԺ4#"�5��)�C��X�2�rpe�Λ�ǒ>�DB.�����zNv���W��j���6�mD��ƽ���I���ntɏ5�5�*vZ]�l�D���J�`80��F %�C���������ڔP[��G�@Z�;W��1
��N�#��T��8��uJ�\�9��Q���=1���uo�H��Y�E�{N5�u*�I���X��8��4�]��rϪ؇�X�ő��v��
W�$����@�����S�=��lf����Jnn&|�����*�������	�E�v��1��/:��[g,߼����&��1tn]X�C;�1x�(���o{XL"z�N�,Ǳ2�����xvu�e�wp��훓�=�:�婓]�]��Y[n�@&#�(K̔���u.�����f�2T.��O���k�*9��V�b����[��+\�٩�SE�ܦ�ԅ	(��;k��;#_ݫȩ��ʕ�Sr�T�@�Y��!���f�Rh��F�5q�sb]��j2��Lg\�4�&E�i[P e��iX^kP9�gE�)a��6i���l��[��ڳ6�U	s��EU~n؎��ۘ�{i"V�]�&_�׆;�����2_��!"t]pS
�؏_.Nۉ���DǼ,���ʤ����p��\�B�84gΧ+.pTS>s��m��?T_����=Tu�^{��B�x��ɛ3��H�@�Sɡs����Z����ޫ�OK(�#���[d����)G3�N��^!5鞙H�lgXZMi�p�һ&�V���#�bv5l�c:�5��{Ha2�9�_����:��i�f�Ѩ�X��O����.�ѓ�j��*���&�/0O�����8����}t��`o�K��@�;���Ϳ#e�����W\'�E�g��xZ��]�E
���Q�p9�f*�½��>P`�S�4������$�cv�}�b�G=��TGE���hm�R\�GI���&�/sz} �d;�/7��q�������8q�04R��T����ͼ�{ub�Z7nb���[�ݤu4�2��؋�|?E�6Nuk�畸�9�ɰ��=��rD۞~�B#�V�fD��9��6='\[_k�#n�Lt�F���(f�F�L���bA�
��=���K{Vm�'f�¦�٢ڻy	Z�ox��j�d�����ԝ����WW�ۋ4���3ք�9^�X5�۹���7����Hi�f7�]D����9+��˭XW#&���A�x%��/��*�W���"��F擐zƣ@���c������3�h�g������k����W����v��Du����!����3����X
���m|0#	тu��(��0-�����BȬ�Σk%b�z�	֋�fn��Z�<�� vʏq'�CάAc��{]NE�^��Rx�r%�m�5J���F��^c;��9kv���tl���ޘ�e�"qe�Vv\ɚ��5O��%���nH� e�K�˟�X�=��`�s�x�ܕIٮ�KZ��q�q��(�l�vK��}�|���
z*oWm�q��,�ׇmH�,�Ƽ�*ڢ�"�Xɢ�Eʷj<6� Q�k�#:y|hUq�=~]%�W1�ˑ+j�%F,�����#�-Ȅ��ql��YF�R虬�+�h��ҟ!!yM�� ��f-���0���v����3����4��'DAH`��Y0EJe�À�H��.��]�u�/�U%K0\8s�44�:��4��Fy���>���,��N�6�Kh�f�D`�2��C2e�5��)3������~�kk�k1���i�G��_k�Juy���.o$����6���͂��:�r�\����]�ΰr����~��_6wE׷ۢJ�\wl�]���h�f��劖��}��s�X5��OZ���R�0�@����vנ��`��NH2����`C��=s����0n��N�ݣ|�7ϰ����N����~���X�z[�b�^&��ǎ�����-"eR�IW��ףI����J����3�1&�w�㣂Z�Άh\Yj|kҬ�#V���-�����*K�U1ڡJ@����}\/��C�'(Fm%}��b�	���0�*�'w�=�uǄشj�opLT���y�
���JlȽE���깘̐�U0w�}1���j��.�\izhss�
)x�z�^RS��-rZ&��C�A:�sеT��1��I��8�=7�˯
#��8�ĵ>�℉{$q����*���]�G��-�6�~��0ӵsu*�m�!�s�SgN�S#�P�.�f3��3K �����V�X=�U�n�D�q�Wgxr�Vw�Mug�wG��� ���ȶǱ؝��< =U=G=޺��^��9�WrUt�,�9G�u=�
��N��4 hl�j�=��{������"��Au,�vcJ����X��6��o4GG��W�[���[�U¶5ƴoZz�@�V�T����Z톖lN^TcV�־��D��	���ܼ��9U]^����9�j&�A�?��@�	$!$�fH@�g�g�ِ��!���f�BO�X@� NHD�I0��;	$�!��B@!; aI		�������C��v�$&�#�	!�� $�@@��n�m����	�0`����`/����w�����}�/����&�?wÇ�}�w����3f����������3 ��\`�٘30`�����Ho���!�C�+��o���~F���30`����?��/~C�����(P���a�#���������������_��sG�N�8ʈP%�<�r�%��1�x4цZ�[0�:��n�S�EC���j[O5��uSP�ײ���c�%MW��B����ٳ�vb'*T�ڭsoS��Oօ2^awyRÂ�̵z%Y��"�nm��m�=-kj-z�P�݌�{	�Nn@n�aT)����*,l��kВ��a6ah6���myߔ�V=3v��^u�V"��� pV�oku(�2�[&�R�%l�4@��Um`��c5�
��P�L2�!QJ�E��W(CH�x\�4lf������\.�P��q�L���v�[F�Ap^�t��̹4���e�^I5C�5M� |fZ"��LH�'t���G��R�5��s�52捲�Y�֥�����b8�^�Pˏ0V��#NZ���݈/^J���#J�w�k�*��詑
ji��V���PWi����x�z�'-]����
�v,+�@�xb�:�)Зi�VMm�Sjţ���u�Z5c�,JŬHT�苎f�^
f���=iPC�U1XlK�
sf��V5$u����j-v�	�{(ۄ�w{x�Sh���qE���RZ��oi6���阣!$��6��RӛWeQ�J��C5Ft�@�z*=�Y&V)&n[���i�˗��ku(i[I�ϋu���T坿�Ɗ����fGlV^^�W�<�6�����&tC3HL�B2�r��@���F][�5��EoB�St��e���TBr�D�ٸHŕ�;[��u�b�H�)�"�K[�j`J�aleM�6F2*�҄��%��;���s .e`&�`Ю��2�f���v^�732��"b�oysu�5
z�	�ԌY�p�,�Ő�e
����&R�1t�س&�����:��e��D��F���0�(8��Wz�fMcsdb�XF��;xt�j�@�%���H�E(�f4M�E.���۹}�|������!!"��B�@!@a$��HI$�����t@�Y #$��A�2I���H��0� h�����~C�Y�30`��� ����x�������N;��30f`�������T�g�~���s�վ���_ϯ�3�Gљ�3̾N�����������	$!$�VHII9��������$��X�>HI!	'3���aSLJ����I܋�����f���~��ə�3���X~_��	`|�l?�hq������Ɲ��3�����?��>����3�D~���������L��G�����C��/�x?���;m��3�c���ǃc�C?@�}�V����0f`�����+������ 30��ߟ�!�������e5��+:�u� ?�s2}p$���|����JLM4�]��z]�R꒪����.���W��k�UX��]�;f�q+�����H����*�ֳU5����m7Zze��M�����r�:Qӹ�8t�%u��k�v#ZS]��d3Y�u�m]f�"4��Wv�i���khҥ��
zͽP�N��l�EeJ3e��T��ԩ�n��      ݇v��� �w)�k�vd��`   z � �t@P<��Av��wa�(�i����Vͭ��V}��Ygϫ���$Dm��^�N$;�
��JxOq���P�����s�5M4�UJ�M�m��E"�T	]��ukRR���J{ڹU���4�ʊ�B���gZ�����Ν��j�m��(( ��`�w��� �����;�6���R�7ٷ7=ڥ�v���T�e#�R�ѥ���+d6�J�%����m�k���SDU��u[�زfc&�a��n�l0������n��ݺ�κ �fՉm����v����gL�Zs����q���i�U�5��㷯{�����w�����=զ��t1�.�m�)���{ޛ�mۺ��5�j^�N����y����F�u��vʼ�W���u�Z�eJ^����Z[�N튌�ݝz:n�ۻ���U^�Ǭ'{�]��l��z���et�Ol�eww6�����ף׻v�[t���i��Q]zS�M�Mj��kYs:WLoYp�:
��L��;̫Y�ժ���u�ƏN�[j��U�A������k#-m={��E�(������.f=0:�u�6��u��Vۼ��ίo@I�zӫi�C��s[K-�9����t��s�=�h�w<@S���/���V�[I�gF��N �zr�c=�maz�o<���ݵʝ�C��3ӕ�gm����:
����D��N���֪S��w`(mY���k�޻����+YV��҉_m�
4��ܵ�Zr�Մ��WN����������]�{��킱#{Y΍6b���5R��^�ι�QF�V����e��V��X]��ն��y��Ͱ�j]���N��e"��9m�jvݬ�ww4+���lnZi��{�t��5�ㅍZ�Y��{�{��]�Ov� uM��j�������ywY�j��k���iy��s��M��l3,/i�F���:]z��@.vpz�N�Q�{r�mF��j�U]�t*����R�� �����#sn��Oj�QvV�ӛ;�<���u�\bc-ۣ��ʈ�VW�N��X۫�:j�M]����s�ft������F��Ύ�ӮQF�%G���Z4���T�&��M�7z��M.����=㮼��ӷwA��Ӗ�i�:�񳶲���l>����ڧ�? 2T�A�� Oh�JJT � T�Sb5J�4=@ �JR�  5O*UO(��M$�J{Jf���'��W��|������l����N�����\!?ҵ9���f5��x}K�_�>�}����y������HN	!!!��	$	'�HI I?�!$�$dHHH?������
����e[��}eH�d�N\��5	���}���Fl�"f2�ĝ�#b��f�Ī9swe���q�9n����]�E�XI�Ⱥm'��i��u���J#dZ�l���"]"���;KR���y�[70)˳@�yR��!��*�@��b5*LŤ�#�X�Ct���Wl	����I�F%aX#������<}�bǰbů���6���8ip��SOoXH�����{�]FʄḖ��F�D.�U�$Z�ȓu3Me:ٛ�Ev���ido~ ��F�E���{L�T)d[4����'ie,9�������c�j"��6��J���/"tq\�2*�*���Q4�Ǖ�%B~i�I�nU�m�ς!z����[�n��`A�I�ϴ�Ġ��h&m(�Ҭ(ZY��@���騠z�R�yZ,�B�a����B �d�˭�C�R�Yx$�f!_W��*��ūX
ͅ�cؒ�w�j+U�-j��(:2w���K6OB�I�m��܋\R�s<'azF�]�������B��/��c���H�{�c��-�Vպ9CRBlu�^%���x�*B�����lke�����b�U�S�yV�Ԡ��&ĥ��V�Z:.l��X�ץ�:F�m(ֆ�y��EE1���LDU�t�'������q�on���\b��"a@�%$�/�A�+l�Nh�n-l5��w�����h��łKؾڽ��f@��>��>V
BhQ"�9�&.=��}�W-n#B[�[h:ܬݴ��
ݡ8��H��:<FO��f���?�ǧw��,.��QN�:�x�-�#��XCv����!pJ�q�V���.�l{���O�b-�{�P���{�s�������b(ň�*"VT����(����DDb"��
(���_��M�)�q^[��a��b�aY�V��" [Gqʰ�;�M�^(�:-�Ͳ)����R��yj����ڲ�4�@}Kj���ds�4��(�{�]��{��j�0
�[g&�^�u@QUI���̹����QK��$J��]�h'#�{T�t�l�Rn�`)����S-K�,�Aǔ	/�?�I{[�Z4�p�{�<Bd�o�bK��0�75F�4�7��U��_�.�Uh�k��������_:@]�ݤ�6el��
KW�:w�9�<�@ұ�(�R,"�� �
\�Sĩ�<�g��ך�c Mx�yZ)�c�%B��Vi����Q�EDQ`*EAB(�H��E$"���2P������5���M�5ofh��kzY5,^3,im'���Y�%���M���SO&��i,Ӓލv�ً!�֌�X8i
^�h�X����vf���'��C�fոK&�ͧZ��4�ڽ���X�ft�Җ(M��m]��[b=fQ X��H:Ȇjv%�͒

:�b+�^�6nkMJZN-�&���� ś����e�T�.���v�mݺW!m!0����OI�h��+�^ �h�m��`ВssJ��$l�h`8§�!�bGb��-�j 7u�J�*�n�3��FÙ{Q�*�"���V�,�R�%󬍦6�<H\�l���L�L�����Y���ۻت��;�;���@H�l´]�-l8��@����G�HP�Q4�=�v�ſF�L�u�3~6"m�z!(��.aD:�FҐ�7�FQ��{���pP�OVq]���^Fch�̶py�4F)�
�f��$ ����3TA7��5�'"D[J'�ʽtʖ���{i��Df<)�t�iR�yPĵb9q藹�@.����`,�x^f]�J���P/tŚ|���Cͽ:�c�`n!��f�=��Ȅ���?y"����7�	ؓKmi'zQ*�M#v�ܦ�](<H�f�yoN*��bbi�e	��F'ye�.�r	O�낞��I�EM���C{�1թp�"Y͚y��|�3����/M�t�UdQ�*���;f78k�� � 9�CػV�f�4N�2�%Br�Ԏ�R�����9��Tm�� r�T�C*弟Hs=x|�����s�53��܀��v�`�0C3sr�I8K�M	S&f���:�ư�]z)t�����N�(5������	�;��S-ԧ�A��T�]���؜�Va��w&��.S�y�ﯝ���b2���"��b�*ȫ"",(m8��Oh��U �R���Fj�?���^�1`�[����֐/Ix%�#un峔4�0ll��Ȗ���wLش\hؙ��M��ӽk�US6oY�.o���@�ɯ�7'n� <|޹�֎#��L�1�'��l2�<����"УCH��h���=�����&�����f����UH#U��6���4}E��͟A�@�5I�%2��b]�^��e�����CF��]��<Ϸ��dM�X̗˘1�i$D�6�ju������YL;�n�*b/�t�.d��rc�ɜl5��������@!k^B�r�MɄm�D�	Xx=-���'t��$��{G#6�`U��V�pmY��B�*}�Ñ��C��S2�Y������R�b:3L��K�Tׂ�$��`���sb�Q�ܮ�'��Սr�|��+!�4�D#�������Ie�iJ7j[��+��]���v]��IX��I�(�F�D��f�.��B��f���e����v���SV��y��U�9�Y��$�t`/��,좑Ɔ`���m
�	
V��+.���#&^fe��@ov�	m<�b1���5rT�X]=S��G6��g�Y���i(�0�'4�J94��[���$e8[Q�@,���AZ��K�Z��fm��'6��f&vn&����.Z�fU�N�SPv
#p�Ma��+�{�4lolm*=p3{�-��j���/.c�p��Q(o�M^�KS�V@�����B%hسP�yX�2cRh/*�FϬ7L���g�$��Õ�Q�DV]XX���f5$�y1jǎI4�Ob��[
d9�A�Wb
ISf��ee,��`x���A ��1�#$���	k>��J�o+@�V�[z]��%���Vl~SI���V̓i�bx�1x�P�!����Ch夯�5�8�	6q�5]�ٰi��d�.�jÛ��*h��yg�Gi#�FfZ�mZ�AR�Ewe�fVb��pU�1V��ʈf�Q��J�/$`��C��V�N�5������^��o+�3��	���,6ꈼS��7+!�l	��3�5�<�[�~W��$c�U�m9VU����Y�֥g�薀X17��x1ؖ�fZ��,ȭӬM�		=T�!H($۽���	�nD�.�H��n��
�y��+�*m̄�B:6��p|�4{�j�FA�41Id}���ub�R���+"U���B�mF�q�OP%��,I�0#!&l
��ׄ�!9�Q�O���{��������ʙ�w%mh;`����`!�U��!u�=Ǝm�NBڄe)&5��Ud�*@kW�nޫZ[O��͓Z�F�m#U�CV�4�,b�sqH&Bl�Z&("/F��/)�	A&�aޖ]�������VeCwy&���cN�alV���H��Lw�n����5'>&5���m�Z��7Y7�{�N�����UaNޑ"�L n�Q�!x(X�P[�˹I�3fe�O�f�G`�QrQ92VS��N������ڋV�Z� ^�fGB���[���F�,x�U��Im"��6Tv��;&՘!��n�Uq�Y�kma�,tn�f�mT�BL�G1M��) ڠ+jVlH�7,�i��\��n`�j���sZJc��f��k�Wr8��Ǉ<�p��}�VC�|�w�_5"�'$���t߅�¤oP&��6e4�����#s5�����u`T�ic� ���fGz�F�rtw)�%ޚ,�(CPob�yc�qk�0�C:��SyI�pΝ��.83�(�D���<C����E���[*ʕed��v���#癣w;Ữy��ަ�_o���+4��M)E��h���kR�-�[q;�ӭ)����P�-�E�P۬g(��Jස¢ˊ��XY�+��D��`�i	E���IqtS!k�(m�V�c�b���Ҫ��5I�(c �Uҿ��
�0��kks%L���0��5�Eݿ�m;���(����)�Z�<n�#�n�b]fZ����w�`
���H�W�q�I���j|��Oh�-��1G=�^{H�EX�0۫?=o ��v����e'����o|>�>�G�C7�C������\E�����
�X��[�m�{�����'���.Їo��WEh�'��,A`n	%4�vU�����u��$�A����K�fM��ʈҳ��Xb3Z��h�W%;zIt�ul��{ɷug8,����yqed 6�+ݍ�2�R�QK3�U��.�,��Hb�IQf6�sdf^��U�ٕ���!)4^m:����n7�o��;٣�/�"�'�����X;���{��!2��i�-f(ݤ�nPͤK�I�t��BnAW��n^���Y%7 �k^X����13��
�?jݛO2�
 �\�>E+���E���l�b�n<�RM|w%���a�D��M4@�K���J���mlR����Fl��cwx��H*��`i6n�F�kP�S��y	���GܺH�C�L�B�+b����2]D�&�
S����@y������]r�5Ji r

�<Ab���"(X$���eU���oq�Rz�#�`H�}�]_`���@Ru-ߗ:�9��BA<�v�m�{ɐXt:�[XԻ��n���˙xj��h������&���iP";���;�v�R�����2�/^�r�ۄ r�̵��e�wYOiE	t�"isPM�e���7,��M����L��R�<ZZ���g�9�z��G=�w�3��h�pe�9��\�T�.h�2�0���w�ۘ�[�f�݉��b�	��X�+�8>F懎kM.I�@(� �S��[1L�dƑ���).��0A��!h����� x[t�V��*I��zCǶ��V��a�e�� �ƅm�8l�LVV���m�Bܡm�����Ǹd˱�p$�8�bn�)������7�צ����aJɰ(X�)�C-�6�'`&t8�Z��
D���i�Joi���)8�P1|>zkb�bjr��*��un#k2:6�Fh�YQf9��]�ƯkP�B
fL)��4
td*2YZ�R�úUY^춪�;�+i�@�(�x�*���	/@W��EqJ���b�^PJ���d0�_�Ԡ�]�SKֈ�elZ�8V�C��0'M�`��ٻ�X������c��XVQ���4�l4%��8��s)ބn�@��0>�}�S���᭗5��Yp�FX��w熂���X)lP[VY2��M��W�*�f��j0@g���|����d�5f�sL;���F��4�Y�p%�i�&]�\c5�sOt�;G��G�`�6L^,v!�ua�g��F&��n�
�]��p8]ۼ�mT%�B�"D�1�q���ɡ�����+lA���
jj��jG�e��}��^ijԡ/T\���;_�x5/`�����M��-	 i��CB�fjzȬ��+RνL�v�RH�:����Ǧ��[p���5�pU��.�<�"%�!��0�.tV�ʚ�4�p��h�D=�ޯn������T��"ں�qG����9�ѢA#�&Vټ��x���%B��4)he�`�&붊L��f�<�[ ��[Bح��8�� -�t���f�G)����V���m�n0�m@���׳?N����Lr�鞅)��������.ö#�r��Wq��9�����JY�LO)�f�[h��x|�U�x-���3���h9W�,�`� �4�LW�}f�w�wMx6�v�ɍL%=`���d�� j�,4��S�,�R1���iS�7@�|
7OM�S�e ֠&[e�x�am=���]h� -�>���n�P�����`���9��!e{�D�½�f��"���e
�j�H�̂��ZV��ǀ��ݺ)C����Wr��j㊡���Ejؕ�	�G����?��}r�,����W�&�+�Tn�����0 ���d��Wwh�-��붌�P�9��O�Eh�(��{�/����-��c�~N���Hb`��t}}w�8�je�k�n��P���%�%����b��9O,�GZ�X�*� �Z8�����0$�Z�2oϮ���)��]w9��)v�*�׆�m��M�ĝ�j��D&ms{V�Q��t��rJ'�=�cu`��G��"�=�C	m'�9��y&�=}�>�1R�]׸$�v�B��n���^�}ӣ���qg��{Ei+p��U�q���Ew��{\lC�����C^��D-Z�\���ϱm���{�U����'@Y�'I�q�Y��=���
b�2��9���c{dqw�O��.��T}��lK�-ԙ��y)E��V�WvF8,vsNp5ף*`�9�Ӽm����|���}��k��V!Yg:kݸ�	9��q�	;N���zK���!@�Ŕ	6�5w;�xq�m�����e����L4�y֭�^������Zv�W�P���/]xz��9�����N����:m�Ԝ%+���%�]X}@�'Vr�k5�[�[�J�xwW�RWf�"�,��%�h��#^�n;�TA�����f�Zu`���R]� ~c�]շ��N�T���pX�)��k[V@릪���g'6��O��}Yy��e�`;o���d.�7i�v���E*s�0͌˰�Hw�k�s%�:򸑋�	Pd,��A����g�9O,,��F;=���C���]���.�
vP���-��:��Vr8���y������ �ϻ�]s�GSzb�E�.�>���jc����Ԏ�[���Zro7�>�Z��v��%�\���qv�zgb��o#�{�� >�h�kѡ�07�:ӡ]6V�h��^�r+����d�l<2�����v"����I�� ��S�e!���i[��u�Ҳ��.��)xc�BYtF]�.��]UK��O��de�яs~m+|WS7�n���kR<�U�w����;(����'��z5�֫�J]��@'u�#W�3]J�ꤍ:n�T��f*|do�O�a�}R��M+�%�pO'f>e)�g�w*Cx�Π��j����
F��V�q�w�,�y@�e���H�1�A�8Rqh�n�5�*�k(�ػ�{Ù��7�n���ҫ��iJŖ�Ϡ٫+��9�*�.�Ck�ch�5���\�W�U��a]��;&QZ2ݎ��}BDyC�h�y<q�[,�x!'
8�Z���N�{��	7w{Q1�k�6���=5���{�Z/ԋ��0�:��g+=�.p�ϸA�R�"��O,c�a�J,2���$g�6��ܓǱ�>�i�L�C��I���|��/v��;.?g{��y������y(��v-���K4Ľ�ӈ��
]�M�H�i�(�]p�&K�Kzހe�؛awˍ˭W/��h�P8���i �};����8"�V�%�����J�����ѫE-ǍÍXS}4r8���6�ZW�x3jv=�'.uJz���%,bh��yC�� u۷}��[W��i�7��*��.�)��Юꭗ�%v��HV@��hC6hh�E�Wǀ�)6�:D�F֫\�,H�v0�HٍWV�D��k�/I��QDl��0���f�Z�(���<�s����
��ysZÝ�vl1Z�V+��J��dt���g�S�;���(K噺/��$q�Ӻl���QN3�%/��(���nk��AӢ:�]�]M�+�3���n�ӲP�k��YE����wcH��:�l>u�44����w>#�Oj,]�A��;m�1��R���3��@vs�]�@L;�����M��Rd�i7��u�.��fT%�he
�z���ȩ�u�ʛ5���:�&>�b��6$�ѥ��b��Mr<��P�z�f�e�D��U�����K�燺s#;�F�܅�QQ�Κ��3N�*�}����o��,Eg�7����.f떛�����{�g	��nr2�s{M��B�=WB�:j�ʽ�����+�f��SRL�ɣ{E��&� ���\{ӛ��,�o;��'����s�9���?nOZe�N΅CXXg�3�������)��Ï�v����u˘9_sδx�RW�����mu[�vy���g5�����
mVt���
WY�˻"|�w���8�M����%X��;��׮�S	¶���͂����j�[�["*�Cp%�G��b)�ip#n����5ق�M,�S�Ѿ�,��4+17�w'�Q��Rw����Aţ�r��Y��iR�m�p���|^��,m���+gQ_ga:�\�lbY7b�&]�Md��W������-���On�̜e ���)b9�桬�D��o��L2e��VQ[6�9���-�[J<��S;��撳�J��\iY�"g_gH�th��%%yee��f�3]�|rT�@���g)Y�8��77��TW�vY���
�N��pk����9�)"yr�[�>�G��t9�=Z�/�>��#-7GN�7\�#�|f�uf�����!m�kv�ɛ ���"��pmS�3�j�+mԸ���w[�[fb�8�ߋi^r�k���\Z%�ͣ����������'N�t\n����լr=V9Sܜ�g�|*� a����\1u� �.k�K��Y1�w���K��OJt%d�lt��1>�K��ZE]䥈GT�7}�n.����6U���b֪�����K2�U�Cڗ�_1�nwaA<�P+ XCJ�}���63�3vBƷ�$��F-̗�:�%;ᠵ0V,��5�D���RT��b�n9G�/���g	��=2�_Z`[RN��c��_'\H�ٗq��׸����f�[�,v`9�Z|{�%Ivβ�R���P��#6��+[Z�:V ����NW�.�����[��:i�Hmk�ݎ�i	��z�����M;䜬����q-kw>
d���ަ�i+ki�ɡ)Q:W��e�Q�Μ�Q��q���I��3��v���j@N�َed޺��F�F�*B���
c�����;])دY�����#��/F���aF��u�d��n\�5ËI�C.�f�f�o����kU����w�V�]1bA����l*����r�J�
	��)k%��
�4���n�m���)i��ތ]�WB��1�	uݘ���JU�r�n�N6��Ǚa��EG��%m��2�k8�[������V�#�9�P�އ62�0�%lM{1hZ1S�:��.E��j�ܲ�F�򠚹%��X����������yT��H�� �Lh�4g\U|�_c9R�����^�'�ox<�����@W:㼨�9�	�T�����$+u����A�gN#��7�gg�{`9��\���T�3ϧ|jx���!��a���z<+���j�s9V�ǬdmQ*�o�n^?mYr&Ĭ/!a�.��'AE\+6F�f��-�� �[2����
<;�vӘgz)�R�,>�M;�[�2M��ON��r]Zr�>E�|^ȶ�
ȨI�=�>��(<
��I�Y�y���H�V�wf}�t��ɇ*�"�9�e����X��%����QSwF�4�QZ���Z6�s�{cxr���]`�7@�ݠ����
Â�,��3n�E��#��g.tp<z�Y5,�6��z����Fr���W&f�0)$&�� 3�*Y��/I6��{���;�_S���-$'��]>���<�����CtȬ������֟s�w���(��u��ke2�\�w����}S�,[A8�LL3+k ֗-��&G��&����wh�)�33`�}�L殣@�U�o�G���y���ʱ��-&J)�y1��-g������T�	TX4l:�v`ε�.��[�R���[�B�����NjV�PF�A��`�PoX�}��;L�'��ݻ�q3a�s/M�e3
�A\}�E>b���ZtԬή�h�Br��|u�tMb�2�$�D��ݛ|(O��}��tZ(w<�^��]��wd7�Z�g�'g�����p�7��dy��#���K5��$Ƃ��(����l�3;��N�j)�#�9��r��Ԑ��H�]�M#�2�7S�)\͊�ޮ!�y��%i��V���j��9�L�3���if�Rj�t��YZ����"ͭ�j�e�P�)�n�Q|ha�}�Y����>��p^�U9Vut*�X\��qL��J).�4D!}u����i�u��vts3�J�}X5]�+�aYuӵ�ωw��FY�:q�R/_
,�n(�h�÷|3jHo�Y��)��y�؋��n����Y�8�����̴]�d��J�s���h��Q�����}���S�nM����/dH����3�X��f5.n��33����6���2pSJ,m��.W7�T���P�j�Y�&w63
��Gz�c� ��)C����׹ء�ЈȖHT����*��>���$�׉��"O5-Fs��hVc�(�X�B��q�p�,un���=�j�aj3J���l��qRo)D�6��&=H���D9v/3zǦ��݋	\s�Z	�1��J{lqOh�܄ܥOSIވKQ[Z۔�����6��n>"�H�'9��3o5�&R.��KѸ�XM�c��Sw.ka�b��C�͹N�7Ɔ�l]�\�Ǣ��l��d/4�淊�6;�٪���+1B�.�..�Īqt���^B��w��1��3�Ԓ=m��o&ǹ'g3[�Q��l����Y߳奾�:��}7.��u���f�|o��WH�!�kNޒ�����2��eH:�#�b�ݷv�q5z ��W���6�c�<�p\z.�}�(&J=�[ٲ뙼��?�*Qvm��<�(��r'p�ҀS�$[g�o�)q�Hk�\�E^Y �N��N`%���V���QY�-s���QUћT�}r��j5���^d�u���6u�Y�J��:��u�Ԭl6ǴU��j/��풣���,��� �Ҟ6���M�+)��}���t@���z8�,r�3�nۆ�$��ʆv(os=����=����`�d���V��#�j���;�2����Y�0�_�#X.���^#�Fo����-�j\�YIv9GV9�M�F�4k�f�֎�Ef��+xpMlf��]2җz|�0�o�ٴW��T%2�[<�_e���yY����h� ��4����Ø�n=���)M����~�)R&��Ⱥ񥔑+�A��M�v	÷��O��X�sY�/��qX"���؆Zo��Jǽ���se�����볒�VifU�Hړ�^'�8��&se�S�)���kW����˕I�b9��u��ԅ�n��צ�K�tҨ��N܊l���=�x���0���F	ׅd��V�8pWIVYT�=I���)H9�������[��j�|����l�[���s��c:TV6�����w�ГD��еz����N+�n����ʋ�PS��J�veG������_\�V1V9�U��V��ħ&Qw���a��)�P��(f��m+��΍?-8Q�ژ�v�T,���!|�E%�r4���n�c9��mA}��p{M�]aC����T�[ٌ�b����7�m�;+s18��X� (�)�V��ClX�;G�z�4Ɍ��&E-4V빠�[�%���U�����e�Z�Mm��N�3��X��>���M���%�m�E΢h]�UպnI�m'W��>�fo.���Y�n�4-; �.�,Ts��`�Lc�.l��뮜]݀�q����X�K�6��S=٠�j�`�@W-~�"���.:"�ý�כ��.�o0'P;Mf�!OO���������0�?�o �Ǟ�����=�+r�h�30HQ;f�Z� ��7���f�M�˻������i=�[�d�p}�`����'=���(��Nv�
9ij�Dx`����C*������e��w{��V�F���+f`��ܦȏCtc��k�1�vuC"�|΋疨��7ajݾfD;� 9gg���\Mޔ%�Ǣe�/�Dߥ����%�CtC{I�}��4�xu��D[��ԝ37Q����^rӰsh;� k�4��U�.��I����h�ϳ@U^�	K�t�y��Y]���=\''�ζs̏������vCr��fu!�\��,J�xC��,�V�oN#c��5\���AR_
Rg[��Аn�H{�����vsf�gu��5���jPup୾�����[�&�b=���E�1VҨ5�tK"�tc!�����'�]a��%%W	�����Qʗj"(�e�Dzgm�+w�����snf�a��κ�u!靊]�!I�<\v-q�$�+ݯ%�g�p2��:GU/O[Z����72����T=�~�OP�w�	'8������6�]��M}+�����S�+�l�䬪����Y��x�Z�v�Ѕ]�nX�F�keJ�K�R�0WGgg_-
-I�����q�[�y���>X3��n��~��ױ<c�X�%;aā�a���L���	P���\�e�����tJX޽��n���kR��ogZ\vWV[%΂2�;�$m>���[�$[ڊRx��Z4j⿅��h�QE�k�`�k7\ʷ�cE�ݵ�<��`[���T=]��Uҵ>ŷ��4\�D��j`/-S�h�R�ݸf[xT��UPo��JZ���`��-N"��=�_&,S���:�3�S�/�#�1�n� �e���p��\�At�j�CoUn��v�1�"��kuw�!�CX-��IYK7�ʱ	�op���e�p+���2��eLn����̢9��@$����@> �P����=B��B@�5�N2'�w) [HH�`@� �I$� |��$�a	đd�8�B`	 �`Є��H0�HT!�Bd�c	���aY6�8�r�@�Bi����d�LP�BLH�	'�'���	� x��bC�x�� a!��bd���b4�Y!4�<@d0d��$�0�a6�iL� �@!R@�R���q���'Rq$6��Hu!=@<I'����'�i�2$<Bl��Bx��HIR��l$P1���BГI	<�L@&�`���(i	0�h]P
�q' m"�C�Ci4����M�I��$�6��N2Bc$��	�$*Yu�Đ�2@Y�AH�I/9����c&�6�=Ad�oT��:��1�ā�''Aa=�!<�P(�m��Ba&��vd4��@�u@j�1��Bq$�0��A`CĜd�� �
�z��d�&�u �a�@��TP�l$�!�� ub���	��VI:�vIX�.�x�iy�Mr�M�EOH@ǩ�&!ԇ�Ci�#�:�,���$� �+�IyBN2Ld��HHd'�8����l��H^X��E0��@��`m����ݐ���@�Rg��a�1�1"�&����a�a㴛Oh��x�q�6ɦd�I"�N3ԋ$�:��R[ ��:�Hi�:��8�u�I�!�I=a�����ISYHkv�3��I�
��&��6ʀ�(CyC�"���!���d1	�'RN2��LAI�4�$XcP;�!Y!ԝHs�IԚq��(IXx��4�B�@�4��d��;���8�Xq�9d� z�(J��-M3��0Rӌ��Hd�6�v�X��V�Ƥ̰�&�`oz�&�XOd�T8��>���q��)��S�P�)�z�I�a�!Y4�_/;tz���Ff�)�L퇩���kt�9�m�0��o)1&�\��=���x�a��یV��d�I]�Ԝq<�}O7�@�u�i�LJ����A��2�&8���7I��6��,4G�?��M"��$!�Z��6�c����讃�V�K��S-�Q0�<��G�y�1aԻ�&q(u'�uC^�\��yl�[�b��f3�Ǯ�G��7M����z�<,�;�Nu�g�;x�ĕM�}�t���R�7���־��(�}KO��G�������-��T:��ۉ�����0���Y�'#&���BI�'��Q��5 3�AT�A�B��r�Y��*�Z�6�z����Y���T B���:�������?\9{�TX�M��%'1��֮�hZz)}�e�7���av��Ֆ/>�%l���㴽��vf1�\wu%5(���D( v��S��
PGN�2���9dw��Qs�"����'�;+��*�:`�j���Nˬ��-�w&�9 �%�un뗂��Gzxv\ژT�\@�q
����P�(U��g��Vm�@Wu�"oYxb��$���ru�Uf�;.pj�8�J�hփqp�˧���֩|�HbW|Nf`$��[;FQ.X����:�E5X-5��G�y��T�t�L�P��':!��m�%r�1K1A[a! �%��W*A���d��B�X4�e@k�V"[xf��Q�����A�1�,��B?���vHAM[��|2�cT�LR\�V����Ӵu5L�bf&q�اc�/�$���-����N�-".=�E(U͹j��M�����ck7<+�����ʆ�շ��v����ل`A�,e�ٹ���!fx���7@E#�����8�5��Л��H2ֳ�(7Mٙv=\�r��(n죀���,��i�V�1i��o�����`�b�5�l�E��	���;W�DMD�#�|��EmP���ND%0rY�����꯾��R]o{i���
���s#��.R��!�%�WaV��}��z�is�5z���D��%Ag.�-q�vL�֡�kt��ȗ�g�3�v��b8�7ͣ�|;"-�L�̥�o��Q�o{���;j��.�~��uU��h�+��|�X.ܵ�B�Ջb�>�ym���%׃���e�>uK������9��ʰ����\�M˫��J1]��ɔ��i*�;p�Wݴ뻨�4�DGn�uE�f�����vE��䧒_1�PYa��c�0��]V�n�fՖ7B��i؁^f�z��C/jä*^���N�Y�QY�@�x�k!��%B�J����Z���'1�h|�MK��V��q��;�z�X���k�n�4�Y-���f�e�D�f�@�d���Ʊ���՜`���<ǭ�|1B�ڱR��r�]0Q}��XbwqY}B���p�t��1�R��Uc��7��h��vv��".��f��mb8����"�:�=�GA��i�sν�G|+�)2�r��*w�[���g����J�ƕ}��O웽�g��a'�	&�a�7HR�૛OX�!�mԏ`�4�����i-8Ò�ڏ�̔���A�������P���;����T�/��E��B�&�3%r)�:��̫�TZ����ly��\0��7�Q�%��
�y+}��2�ܒY��c���z/nw���	�o=����{���ϻ���N�VX�d�����0|t'/�b�Z�x��ݴI]���
�'Sge�I�Kfuu��;���Ą!�*I 欐��@�$�I �Bc�$�Hq P g<�I�$��&�Bc	
�B��d RA@�0��$��&�B����	�z�P2J��$��BbC�!*Bz����#Ǽ�r�a�)����=�w��;��{u����>H�QP[h�ЬQb�������Q5aEH�(�E��`��y��Fn�U$Rc
�#E�VA`�PPU�PF��CB�QQI��QH�b�0E��,X����/�EQX�7��E��Ōb�E��1Eb��"#"�־ڑa���u�LF1DE�+�dċ"��( �"�U����F"E>|Y��R����"��F ��[E,ƈ��EH�QϞ栰UTcUFcF-h��DPQTY>@�O����c�J���"�NR�*�!�X�P1WS��(��3=�H0�TP�&��g�DE#��X�#�QTVS�r����*�EX?4��GI*D�E�Z��2=�W8�f�Ź���(��Ŋ"��^�"#TTKoZ����E�PDVy���(�Gv�h���*0P\h��DY���X)DX
��@UAo.AQUEXz�����5���U,+�K�T>Ɠ,`������DVڑf{��U�EQb���TED�X�ƨ�U�*����4���gr����UAf�1UT��15娉|�`����)�QQ�"'֪�k���}�A=Kz��
���Vs!�]weƪ�U%jĶ�,VP�Jr�!+;)�	6^�ý��D��ED`�����i�|��EPE����l�4���F""��w��@�X�(e��*��|��M
""Ŋ��f1m3*��-Eb(�b�eDA+E�Ϸ�8��PDQ��Q)�2*�Q̤Ƚ�Z�Ԩ���E2���kQPY9Ib�
�j9�}�j���V�,*J�h�n�E����8�)VV"�"��7~��1�ЦҮ�����H �Gy�'R:]�
i��_=��|3^��}�1<��V ���풢/sܚb�A�+��*�V ��k�ƾ�Eb�ˏ�h���^4�bk*�E"���kIƬg�S�*�b��T=�V��(�-�Ȫ��r��>��i)T�Q���QD1*,�C��Qs2
E�������g�"9J,DSm��AR�LQPCMA~���TDF1��V��߸�_�T{��;2^T�$?(P4�@�O�QH���&(�M`WIA*>6A�^kj��`�0q�OmE���S栨+1ی���7��j�U-�UM32Qi�dŊ�R�Ҳc
���L�.��S��Jb�}���Mڨ�UUU3�׻'��ER>�U\���l�|L��U>e!8�ϳw�VP����w��'�f���I�QQE�X�mR6��Q5lX����Ǝ%�*��Q5}¬Dr�X��{�̲Ō-�S�C�Z���جS,��[��c=ʊ������)23�����3v4�m
(�ϼ�㵊'�ED���o�sUDF*��,�EQ2����nr3�����$��<=ٸ\�o�
,�}���w�{�=�X�yhn��UW�ӧEE����3�Q��h��Ȫ��*�heR��N�X��B����̘�f?:��"�e��w��
"�9���<�A��
�/�\7i�f/�6�ǶV���������)DD�b9j��,ӥ�QO�ϩ��K��lu�����+��������x$��"A�Q��_��|��<�GV��(,�Sֱ�wF�d*DVw�{���1�>��b��ɍ��B�J���=˚��F
���3�.���S�����i��UE�K�(��)]6y���
��H���A���j1(W�P�,ZDv6�>�ՙZ�Z6���$l-��}�*���1Ylup�}ٴQ?'����y�a̳�,q
�,K�pQ|�C�����^淺�+[��orW{�B&��UU�WM��a��r)��QG;��U��ek1��wn���b(�f�� �C����hw�e�a~#)X���]��|�-8/��IM���:��%X��{vWh�bД�a: ��ε����0�"f�d�t�$�o�H�� nN�� �2�v�w��uъw΁���#]a���M����ۨp�ݠ���x�{t��v�r"��dR�����1gmDı]�n�GטX�h<s��f��UG��_�u���[iD�Sݜ�h���� �Z�*����Tb&��=�Ֆ�91*J
>}�i�'��⪩Ʀ�R%�z��U��B�O�BZ7�wuY^�Y�N������ʯ��4]�Z�*��q\�
���M*���.�)Q�V��QEQ����SZ�ԛ��i�V^9�]��o���9L�Uu�u�R�#�2�Z9OnL<�Ԙ��+F:�ۭ2}��iLJ?&1|� ����7��=^�+�V��<�����WYq��뇞�������R�n�rj�c�)�wSX��C֋��袂��Cw3��6*��mye�1[g�8ߚ�k4��Jʈ��~�󋦊%��O^��緆ب��-�)�|��ٯ���/�D�]t���e ��=8Z�^�=ٽ��S����=����:�Y�q�u�o`�Y̪2��ѽ���Y,AQ��[�؆�k)ֱ�3�f:*j�
��%w|��(�ݾ\5�wh�D���7���}K����"���B/ [`�2� �F,��ۭu�]I�3}|�g�^UJ��'��f%c�����?a�+i�B����&�ը}�I���y�4*<e�a}��9�|��j����F�}q<M��!���(�ӛ��u���;�ɚ*V�(�E
}��k�<E����~qA�ΥXy�.�����ɛ�V��?�P4��ڄ�V�w�Ԩ���TLJ#h��F:�ʸז�{���7O�4�-���f�oݞ<b��~k�q�ʚn�*�5��.�q�X���].�]]eNҌ񨣿�f��:u���{;Rc+_�܁).��<��a
��1*g�oa�����cmR�Y~�@�T��6�IUX3�7u5�{���F
�J����Ӥ��"�R�����cZ�
���u|þ�i7k��N�.1j#�����kj.�ɀ ��{d�>~�!Y%풺���]_q��4TM��j���(�@�A�^皲lnf����I����\}�u�;K�/���є���}�4��ۋ��eyq�|��?=qD-/o��T�^�׻�1[e�S"�m�.v��k���	�O}�+����@�
c���c�*�w��כ�k0��t�f�u�ݕ۫q��nZ�źt�E��� ��h{������O5PUB~�o�Qϼ��n�QG�fE�˷݅ݩX���|�I�o���Q~h�lֶ�~
�r3�u��^4ǂ4լUo��MFw/uT��6�Llj�>�G]����&bUD�s�T�~jꢈֱOoΝ'�^) )�X���B�U �ԕ~�Z*�Ꮯs��-������g�c����|r匚U�U��+�[�8�`�ַ���%iv`fv/KN�7�J���;��(ҏK�k�8q��X�����o�����j$A9�֟U�x���dp�S��E�ٺndMX�z�m6y�;���{>��(�#'�fR��;���^H G$p������	 EM�z����]j��u�U�x�'�l�T�[o杨Ha-!B�+���R���$~̘���Gt�WI`�[��I��ɨy�~ &�v՛�L�	�%��ML�'��wk�Pp_&�x�R�J��Mf��5ڨ�����~�d�e���\D?(�i.a�Ծdw<u/���)���V�l�481����L��&C���$X]t]-�)[>ar܏6zk�B�;=F���"��)�����|�q�y��_���<��P|�_l؞Z%��L�{k�
.P�'�W7���@~@@� �$��s�~�:b�*!
@@��zET@&�9:I�c����Z妩���s��~|�kR��7�����T��lج�p$8�T�R���6�X�"�����	�>�b���ȌƋlm�{���c����kD�4�S>���#�z���R�ܺ91�h����̇F�"�Pv�! 
�-��x�3� 2�A�_/*h���ᦹF�p���c�d�<�x��t��=ھc��������2��i)�p�����_Avܡ�O��O���y� R�y#-�q�ݞ D�K���g��ɴ�\X����U,�6�D�ZMoW�s��6�t��+LV)~L�Pg��b�3-[]�Gϯ=ru*/>�`�O�{��U�W�_���,-��}M
J���ڲ�(�ۂ�]��C��8'��4F��{(B*� 
��<y�(�D4����Yv�Ǫ�Hq$Z[��+r�K��z�)�P�!�d��Z�P�7kT�DQ�S�+Ǜ����Y]�'.�����x �4Z����H�����}�M�FD�8Q���8D�|j�/�v'�,�Vb �F��z��3�ģl�/���F�+��y�3����v��;z�v�nX}C	Ї�C$;K�T�M��4U����!)��U�'W�ѵ;wU�y�7�&����>�}�ʤ<B�M��tE�<P#��Q��]�j�ٟS��{߷͊?9�b��)߰4_��~n=�ێ�͇�Пw[��>l�nXC�L��w&�xˣ�}���~��,�E�8�Ž�o9�H	<0�\̾���>���1��Jʘ��K���|���x��u�z.�e�r�<��¸�&b�uz�f8���Y�]���T!>�mu8��|�2~y.V>�o�b��F�ޑA�Ǣ�ə6������2� �?�$�����<U �+�~'�̈́Q~����C���[��/�GR���U/�9��{�D�@���	:���H�==�uݳO����{��K�{����H��VU��Y�k}�|[�YD�1��ѿy�v�֯ɷy\�9Ʋ�'F���W�����M�L�Z(���(��{;���%6�{�N��fl�U�ޠA!kuW8/��a���� �X>5��T���R�M�����$��Ύ��qF�bA�~a��?Zl!����)"!x܉*�g��&��X�-G��߯j����
"����u1G=�2&	#\.ω!��"���� 3޾�q[��*Y��a�K�[�h*&�1�O���~��5�AL|P(�N�N;�n1�r���E��̀E�Kڽ��Kq	
����l�3���Y�!���@�<S7�ĭ/yA��K��=Q�HX%x�����]����5�:�x�wd�қ(�%d�K�B�d��
�/��b��N�X!��0��p�W��Z��ڇ�F�̃y��p��v�^��~[��0J+�Z&�.�~�h{d�O���3����A��\� ��QQ���7�f�%�egv`�H��,�H�⏖]2�H�p��DP��>�ѯ%�8�u��$oW�4UzL�Bm�򕜫7��������
^��u|�U��k�&�Ȍu�(25����@�7ɷ-ծ7{ɧQE[TN�Zҝ��!7�m��(v��1�׸5��Y����8q<i���>�z��)L��"I �]>	�0�YF�'y/�c�_tL��u������J�@�T���A|G���OO��W����6/��+�C3��ɨ�6�an������auwJ�(�Y��C�S�j�ɥ�0���/��1h"(5a�����uvz��a���Ŗy_Q�!��H����c���'B�ԙ���NN����fv��4j��vr�eԢ���6�2�q,-y4�A]!�IIW�ə��q;.�S�~r���9�����A������N�x�r�.�M��ߗu±�W��ɵ6D�Ǻ1Xf��Ԯ�uy��=܀<!� <��Ba3�П(I �3}:�m��H!� ^4��\LWz&u�T>F�q��Da���%H�?(�$
�_ύs����Y<h�}D�����H0�D�+R�$<�r�ԃ?jX=o�EHl�
���H��(�OސD�P�l�Lq�$9��4CroZa-L��+Z����0��	���!���3Q�Y~�[�	 itq� TZ�J�����}�*E�MP���R���T4.�K�m � �=�\f�Ph憑!�������f������f�9CHjc�g���u�b�B7��`����W����@�^&���h��:�6�5A��@���o�E>_ݤ�/��]pA�y$�W[�]����Uߧ?SJ�sk2>Y�u��J+u�L?���M�� ��QCb鴑�W��
3$^�jz�(Oȯ��1�h2�˖6O��C�!�a�˾�WQ�p�]�uc����g�=�����Ə�'z�tρZ�O
R�4vΏ��
K��KAyq���P�(rA܀�PDQ��r�5�kHR���6�y����L����=z6�kA�K����	j�J��F��~�A�l���f�iY��[��?2��z Io�ߺ��F�l�^4ս����D3��%�}�X�#[<p��iz�
НK�Q�O�1Ϗy�GTg?�AR��o!�T�i�9͒I����a���.����]0�w�IAּl���t�,�-��_Ƒj���������E�i�B ��d�<�����L�JB�%�b�M�9��_��>:~�5�gx*_"H	x�:o��P�AK����<�<��I528ƾ$hfi�����Dx��2�:+���Ȁ��FNy���G$���)[����jw��o ��_%C6�t"�`�_O%cT����Z|׃(�:��_��f���RB2�{����|@�O}�>�'s�����!�f@�m}du '���h�|�<$��'�����+�>��l�冼��}������$�0��d��w��s|4@4�Ú��_��� ���
^��|6/�X��h��o��O�x��x�!�٬]���Tmԩ�Mֆ�L�%9-�d�ZԸ��k��u|�����m�����b�M�Z��=�|�ҏ��z��ܿEG�eе��@M5I�P�#;.{�ဘ�&�PO�x���i��>^dr�*�	��-���mSXv߭-�S�VPC�!Hl֎@��]�8/�k�k��� ���3�%@�!1��,~_HP�&����I�O� :�;��
hy⪐&�b�����N?�^~&ϸ�����.��;+n>]���;!j� ���F��wC��p	Mu����#Ar�S� B���wE�ֽ�
ʬ	}�(l $_A|�Ă������}��i�������7���o�!$۩�K���\�@�	��{��"��Ĳ)�M�-(1��>_U���J�f0�v���?逾h�~Ao?���]w_'Rx֯Vg�ʱO;(_�"���OȔp�f����	��bT)\z.�-���w:��|�==���;	��u�H�mal%����^�s4�1M�p�c��u��ʶ1�C��1�
"0R�;����B{(ʢl���^�F
�y���~Z��6Ft]w~Y$�������uT������~ e�d�%[�c�=�����/�^A�tV)9��r�!
b^�� B3����8����<W���ɠʍ5��@���bsd#�c�O�����"ݙ����z6f�����b�J�S%
�Q|��A�E�a��"�
>:����$�<$pS��e4�U��@���"61�U�
��/�B��'s�$�)f���
^'G7����	z�4����F�!"��?Y]�3h�
�uϩxcH}@t���ٟD#���"au������Ɍ��;��z.n��x��A��H̗Vg�AMvs���"��T�)�~,�§�_�c��l󌔛-у7�Q�Q��_P7�m@+(_+u����ܫ�.SӰ���"I3Z�w!���Hj���!�x`�HZ��w���}����.�p }����x���aM��s.�W�~| s�����y��s����T�>c�z���}����^���g{�c���>\A�:]^.m�ҡ���\���8(z�1`��M�{��]B�f�v�S��]v֡�������s������YE˼z�I9���Gو}�E�5�O��r"B��:%�d����D�P�� �^�:9|z��	H>�'/H��kȇ���wo���c� �C�L�f��i��ص�;�t�J��S/�`��\�'�_r����H�Z����<CLb�o(b��ؠ�A,��f��4EDQ�:�US��.���`�'�����Tc�O0�C<�0��<H[�BA ߼!�I�OZz�8tz��\B����{�H$m��LQj)�)𡀩(v�U�?u������X�{����ާpPj�*��M*��b^ȥ6�?��� ���0�q-1���X@�Ͳ�K螕�צ�5	y\�$]U�������¬0��1���>Xj��l��r�	��{�x�������;��N����!�I��� ׃t$���
 ��N=IW}eo���^0�7uu����G��G�X�b�s2�����=��SE�tp�Z�@�|�-��(m�tR>�m�����-Ƿ����y~��W�W4�������qa
�y^�����A@j*i�� ��橂��z�$y���^H)>�C�� 
�"}�¦w��qJv��x�ά��#db��4R	#ɂ�3��Q�Q�w`aH�>�;�Պ{iÀ�D��>��|f��B�>d�9(q��n5i��2T4��Qow��y�wy����~�h"��VQ���M��sz��?:�����_H���U����s%_�_޷�Փ65c&�(|)��B#{S�4�i�c��ŀ��Ne�ɇ;%OX���rp�?
�:�TI�Md�X���wK��Ek �@Uޟy��`�����U�r�$~At.�X�|C�f	I/C��e�cا6�}����ǻ[��ߥϾ�kާ�u�>7iT�����f�|>w��!�<t���׽��?l�X�˽u�V&5��홫+���7�i��ܦ���f���+`����4��}��.�C���)Qw��:}u�ѓO�k��Jy�p�k�2:�ͱ9���ϊ���`��^�5��! ���5U��M/�n�QN��g��;�tt!���9v
+&�% ׎��k�{PM[M\R��Y��[v�Ķ�Kޕ�̡�R��AE3c�6�=�%Ix�@Ί�|*9�Od�CC�*ƀ�{�t�Y��ȫ��TT�U���fi���W`�][s`�U��&��{�=(ȃ_��B.%���7���{�Az����b�( �ƖC>^�����U�65��D�xv�==��Zc�VfO^����_uG���_���T(T6��!H��l�'ɤ\��G��O̯�$�J��/�4!���ZV0`Ղ���bt�v�g¯��s��H�=�J4���f��G�S�2Y(_)*�ڬH��4~|ex�EA�B�+�>�V"�#2��m�-Y�^���ֺlk�t���Yꥷǻ&�l�r�	c��,�(�#^ad��+��D�n�笰JZ���W$F�8���*4ۑz�,V�SsA˪���O��'j!KxE��X�P�B�0�l�/�@����I���&(�5����8�Ș �5��RJ�Z�>�������M��΂(�MV�0E�^Tdo�ջ����$h����ʽb��� �N���p���>�\���= D�EV���\X��@�D��N/ʁ.�8/8�U�'-{G5�p���V]C�C�n) �����H29h��?4H��n݁NT �ؗ$4�V�^&��b�Q��J�A�E"Eq��\jg��g'<�w�q��v-2�`���,��L4�I��<�K�Y�J�m�0n�$�jVwt�5	�k�d/4;Yyc��(K�D�Pi�:(�b�oE5��С�:b.��潎�GM��ڼ{�íK��rhZ�q��C�Ikx�c�J��|�'c���F.��t����4M��Z��r.rXP��ў}���3�X}���ɝ��d�	�3�6'^U�����#�����d��CA���=��c#�ժ���L�@�1'��u�/��ILD�?z���nW�[� ~鲪�r&�!�ԁ"�@�+���ϻ��fc��[�k��ʿS�o�]^}�0W��M,,�����l�/��>C�&0t�* }��Z��0m�T���/�[�)ϊ������^A����jy[���®�twLv���Ӫd��9�%a,�,����Gl��V���4�$�>�!���
����
�s!�D����ۼ���6�<'O#y��|��(�צ|��)E��b�I����<����|B"¦�H<|Ƹ@�!�/<8-��5��K}]���eQ"IRP E��L`����L���axRB�����F�=�<7�!w��?�ф�t?Vny�&�0�cQ$p�y�����O�Xq��!��,����%F4U�d�)�Ǹ{�|Q`��P�,� t7��X;�)���p���2�>����iˎ�ǷM���@|BƉ.�?���!�dY�sH�!*�E��"���Қ08�g�;h�R'H��8(gBCWxw��.���[�*�`黭
��քE6�A@+)	8��R��t���G�p2�$,�'���R�'k��҄R��4ӧ��"h�_��
�׳m�W=K��"�H�4���LQ�E	�'ǹ��tǄ�"�:b��(^4����Q��$ζ(U�PU�B���MOI%E[[,�7]qm]����ّ��?r��cEF�{�N�O}��\�B�B�
D�ԦZ���S�"�A�(1�-��|���=y6�aN�sЃ�O�l�؆L�5j� 貣a� &n(ΊŒ���ە�JyBY��n�t�-S���
,�������b�@�\|+������R�m�}RuK�\f��[��`�[)ᷦ��@k��> v��s���+�X/v�p��?z������7μ#'�&o����$��j�K1��a!pﾍ����>��Y�H�J�
~H'��S3=f��*����8�:�0yh=t�g��i��^��I\׻��A�ޒ���{*�U�J�ԉM��i�&�k5�\+G�~Q�.Gў;��X׻�>0tU(�0m���2����XU�q5A��g�ި��\�jd|M)g�߯�(�ɨ�8֭�.;y�����=}3^�ʙ�q��ц{$�Ar�Y�J ��8� Gs�z[2�[�Q��u���G����	�!�F.a���5��L��H������V�Zk�_�:])��) (�i��&�Om:	�>��ZϢ�� �a�sH��ԃ�l��j�2��"����y:jf�k�"J<���;~� ��67E�睌{҃"+z^��㋾k���A+:J��D%E�|�jw�]��]����` �N��I�)+�Խ�4��]��#�rCeo�f�h�~Y���I�K�o;�w��ak��c���a����t (�s��@�
 ѢI�^��{_�%�gN�;����$��ި�>T_ȢΙزY$u �6.�^޻�i��@�V�F��mjp�|k���B���F����`yf-�@��WR�����K��2PO��#i�<h�@Q5�y� ����L<�:�#ܑ�ĤAQo+^���k����dt�% H<�A�}~�\����:-��SE�ysT�/��l�10�o�@7B�TY�h,��=qQ�$�7����/�� ���PqdRa�QyȦ{@���U|�ܮ$z�~��b$�a�e�twgn�����Y��<�*��L%�{=�?v{�:��q>��j۱k��2���X+�]: h�#@�u�f��0��v���b�����ʴ��pK]��I��ꆇ�O�7��En���B��x�K��1��f���	�/5�>8c�nQ�y��P���:���VG���׼{��{��WQ7k"��b����a���^�2ƽ��Q�o����*u]M�z��M�ajS��߮&��[j$c~~w<��k+/l��d�I��Oz����ͫ++03Xc�ee;�Q<�$��Ň[�\�5��%�$|ҭ��e^�vN����r3O%�s���~�4\<
M�2w� �U�
��"9K��;	�2��l+�Y�ՙ���V�̙`���h�a���m���K��3b�q�U�t�4�����P;՛�T�8G,�o�rA6칣��}��{G��u��X��v̸�(̓|35zoh8|���*p�J)PǰHV�����*]�+5�r���O��oxQ�MEq�.�#:���ji6OHӀ��gK���w��l�w<E�"]֏	�a�Ϯ棹1;N&���!32��r�cv��n#{m�)�+6S�Qs:�L�[m�+C�����B��k��|r��\�,=L�[����.�S<i�o���v��ьUw���KV<�T�C���7�;���]�[cF_Q�7"64LRE��!(:�h���"�<�t�?�����w�,�'�qӺW�l�t��WG'�����zR�Y��\	��;8�,u��c5��}պ;�\���b�ޫ"!e8{�^�ca�U-[����LVjc�b.�2�A�ǎK����8z]G�.a�G��w��״G�z��u�+���Ж�a��<���<���[V�g\�r��O��k)��S�!b-��9���x<B�� ��NZ�B��|��M��\�Fx^4�d�B�)N�a��ް7(�#;��zژ-��^b��vE���5o�U��<P�g_X��գ��,�*ZV��V%j�x=��!.�f9�`��*-���2�K���>{J�8�A�d��{yHq1�İP���~Z��]#F�S}΁�u�]\R3f�2��1⬦��X���y���[���K�Y�P"�};f��&�.R�ԝ.?u�C>��j��3ޅj�Er|g��q��5%�@�]W��������� �x>V���/f�X��WӬL��z�rw��-ns��9�|n�>j�K�3�wc����d�I@Ӭ�%��Ώ�V�^˅K<��s���b����ܬ�RHDN5�1P5##z��L|�oﾯ�ꪹ�:��c�T��/`�=�&%@����Pp��x�9]FwU�E!&�8֕����.ȃ�>�.�H۬R���;+z�1�9�u���ЂC(��8���"���15~Úef՚N��1~�^>��SV��&�I�u6�3gi���]k���J~�7E*k�+]�=�m�c:eX\���tg,5ˉ�Q�����9�1'{K�h8W��y�ݘ�N�b�>~C����+ѵ6;�ֻ��7��kz���f:C-��o�5����e��OP�߰4�N��Ӟ�Ꜹ^���a�-z��A�6wW�0g��%Av����t�"�Lf��M7��9;g�hsϾ�S�ٌ�����]��<�/&ޣ�����Xr&~i��n�M�=#�����s7��5�N|�2?z�S��I���hk~\5�Ƴ�ٸ����0�oiQC5E<��Vjn���٤��d�c����7��q���冝���j����弧���Ri�i9�+�4�c��c
��p�Q��z��ѡ�[y�7r�n�o���y���s�~Q��Qe��/�>M&�c7�j�Ci�N�j�t�9�i"��v�)���Z���C�f���A�ri�'�)��Q���p�PĶ���֩(�*�&���8������Ds����W���,��C=������8��/�f�v�����4�W�0Tc��&��'9B�tͼѣ����E��B������N/)�]Y��%j�O�k��|f�fvǹ϶s�d�X�i��y�)w�]�8���N��y�;��5�~�a�INoY矻6���0��*c�s�����^��J��ϟ����_5�_�������7����u��Qt§S7��9C���VS~���8;t��6����͟��cl��k���N���q�θ�M&����k��yv�8���������B)��o��@_��k���O����β�s�!��<�Q0���i�_Ͻ^��8R�ޫy��|g�7�37���_i]�B�M��1��1��5f5+5���p�N&e��hM!�̯���14��ݟ4N����Ǝ0��=�{������]�4�՗�s_��3���'�����P�uٖ+�c13}3|������߽
�]ݼ��:h7+�tj�T���c���2/���A�n?����l1��!��4��g�w�}�{�R�橯iSh�o_uw�bj�yE��Zg��8�y�ܤ��G)���ѷ�M&�۳�۰�֐�(���3<�Ɍ���KQ|[�e��B�$4�����������k��#����<	������t��O��3�g�c�m8�x����٤Ŀ���Rs�m�������8�s�i�=f�-֩t�&7t֩����4�����?2�ª:�9�syM����z��B.;���~�������gE�t��;$v��Y����̯��5��l�}�����3���x�e<a��m����g�c���1��d��k5�}͛f$����'{�����=�Pӏ�:�����4z���v�mި.����7dۭR�ۚ�_�����^��)7�,�*��4E8�'�v+X>�/�c����SF��˨��ZI�)�P�YƎ���K�2�Wr�\]u�rX�`r�t�z��㮽�����E�L�M�g�~bT�S,���B#��Ŏ-f�[\\Om�Os3�����DM��g�����n��u"s�{�oz�y�����&��8�=}�5�YY��j������P��c�a���~�N�B��2�x��=�6��=ι���|˻�IS�LB���_���o�^�pG�W7O�Uh]S��7L��i]���}�Y�L�ӧI�5��h�c��+x�B��A#P�>Dm8�L1�r�J%B�����xm��a�y��.s&�ꀥB�p�7�P�`������D��|tb��2���ſ�y���)�O���P�q������>�u���^�|��?3�U-��Ϛ~k�XV�"����ۓ��{IwF�~�u6�C����<�٠rÆ�bO�z�fn�L�<f��֦��x��������G���`���r�2�O�讗���>����
�A��׽�r�Q>�$���b�X*�=�Ӣ~�b���o|Cj��~�7CYG?h�)�R~�ٱ�J�~�vn�P�i4!����_����c����*�
��*'�|��mY�������u4��TQ���g��6�ٜ�7�jo��)Q?W��Uk��'��"[?ol���R��3��s�s@�Wղ�|�Ϸ����|�������!ng�g��
�4����q'>��=a�)���������3��S���i*)�>�ǽ�}��& J?c�6�����B�D"�`�Ep"��G�>ُ�g��	��D�����z{���}����ι��?'�YKoP�4��Z���εƠ��j�����W�)�L�=~��sV����M���z�
~Bꟓ7E�}ϻ�6�6e��s�p֨�n��EO�k�M:1(�,��q�Ih�J�h��_���y����Ws?d��~Q>|Mnʞ!Ka�a���I����/N�Y������h�H�q�q?%N%�~��N�f8�5t�s��6ʝC{�!�o�K��2��]�?3L��L�5�~�k�m
��CN��w�?a�iW��f14~���,����u>�7�+��#��}��yt�a���On���ǉ���Mn�zfM��V�\L���}5�;EY�����E���l�*ov�{f؟w!��hT�����t;�eN�2�Е�>��֐����K{�]�Ͱ��Vw�|�3�3�z��am%��=�=�a��h�6����3V���uS_���M�Y��'<�^'S��>�9�f�&�LD��*��k��A�n�6�O˽�D�{��F�	��<i��縯�EE�͙2B{ɐz�����:��בkPe�ew�o�;.�D�Qo`*ߺ�Klo����!��~}l�Aj�w�6t��~�S��A�WS���N}�ֺ�é��S��u���ۜ��u�Dq�o����VeVn��c��ú��M((�]���h�G�,���δ�4A���|}4�N
종���_Y��v:rݣ�r�P�pN=^��,V�b�x6|��w���6�/}�錂��[�:��a?�[H�񨨁��F/X�q���JH.�}�b�v��y���頊��.UЀ/(��j]�(z�.thiW;����-"�˴�R9�_HVz���#�4��T�g�v=���w���?l �O;��y�Ճ�_:`��-e+����c�!���(?%s#Q�+׶=)�'L*{���]ʍ��fj�kސHeR���$1U$Y0�Ί���nǰ�xwε����8 \sL�1����_ul���龺�u�@�w�?V`Y�Y,����c������΁m�����H"=�P�ڹ��M���(�G��|^D�ѻ�T	��X��?%��q���S��X��q�J=GJ%���3��5n�4�t{N\��Ǯ��>�D��R�8G^�*C�*%Xo�g��EwI����Xǳ�^�6���Š+d���Q��>m����t7�t@`�� �6��HO�'8ڥIf��&�]-eH�կ~����I����0��t���y�]^�˼��
2-���^{:,F!�B��'/NC���xuQ��ׅR�����0z
g8}�b��^s(�N��f���B�`�/
?�'�[� ���b�>�T�!`����e�Ɣ$OShH�_��۱a I8T�Q�8Wu�mOv	ϫ2����txя�,��R���}�h٠$Z�#^KL
TN�\P�4�o��'�����b��:U���V0'\�Ω7���ΡDf����>Aj��ۺ�{;�e�j��[�@r�nN����n�q֎����<>B>�a����ϲգݽ���2�|4]]��U�r$*[pv.�(�̜n9p:xȏ���"���{7t[��*2a�o��7/�Oo®oe]�X6@�(X�):1/k�]�?�w��*1 U��J�5ˎ���@����zy"\�}R���y�OC2\��~��f���q���b�lly��G�c{�*�4R4�Ֆ�!$Ho㧌�O),���VuW���A�v9�j᳓tC���u��-�{��̞޷G�4��Ǐ�m̔�%��B��ڼ�4Ԇ�yew�F�le��B4�/�f����I�C���q'�E�b>�7f�3
��1�a�)�?s}i?r�o�/O׾�u��%�q�DQ�%;o�����mme{ܦKř�}��ܥÑ"�8�|�k�h��&�4z�+ƕ4��r�-��(�����<1����wa͓rT�$U��Wl� ��+���a�"X^�sYxg^�/��V���B>���(�ǜC��:esD�	,��g;���$�?NA�7A�c�b��eV4���ù���L;{)���kX�DBM�֌Gu)�I��:A��d�+짼����k�ad�<+��F���񧻎?e{\��r�wB>���V���F�Q)������h/iF�o7ֺx<�|�1QJ��B��7co�_.>:��K4,cn�h�f��o8f�jA��ʄ=b��I��a���\���ͫ3ʱ[�n�G �u�0�/u�`4�R0������x�7��ݚ���ڼ�M7�BLE��
�2��*�8�k�,}���E����:>հb�
@��; yJ	�>�h���9�.e]��=Wr����:%�8����:%���gS��bP(ux>��3�q��s;b@�M��ZR���p㜱�	�Rc!��O�:���>�!W��e7������'��6���X�ʇ"6� +�ɜ��PwH8QN�%�]��y��ڏ�Μ�>8z� `�D�5�㣁�EW.
��x$�m�H�V��@�V�(E��y!c4	�=�m��oۜq����s@cQ�-i-}����=��k�Xvl4�/83c�Z ����
,gF'޾���='P5g�{s:�vi��/��v��ڕ�M�=$�A���.˭ϊO���v�QZ��2>�L�;'>ʗ8�z���2�Ѕi��P�Fh�O=��uiNy���hu��@,>h`�#�Z�j�gk���n�r$�m^;�x8�N5a"�#��5�R�h:��ub�ߖwq#'k�����3����ޏ.�1��W�̌�IW�/�b]�� �
fic��뮼��<��F�������:��۲���)�����!�,��V���ܐe�+���qg܋塖�4ѡ����<�C��r���'n�[>+�[�+Eܫ!f|H��.�w��.�;��x�ＮƶT;���n�8.*�ȊW]x�P}hZ��TD��������l�_�4�^���i�잻z>,�/�F)�g��nwz�4ܤ��{ɣ��Ӊa4��j����b�rL��؜M8�a�d0Ro7;��nu'��&�I!zF���d��0~!���z��",�7�tl#ڧb�슁�^�/׮s�w7p�; O�O�e��,�&�@P��ns(D�^��D�D^�J�_��@����g�=\4/oI�W,���0º�]�L`�b�e�Jw�r�ΐ��!���z����4Ġc���	�Z�rӻj;�����L�@>88xCR��Lp��	F�$w]���L�Q���C`�����u&��g��uwq廏�e7�j��M�s�6O]ؑ}�e:F�C=����X|<^}�2�L˘QOI!$��� �W ���%� -��sj.��U�v������x0gR�|�����O�J~�!�P�9�mm&	��s�#	#EM��a�n�"�#�s�TEzc�ֈ�}��6�HC��W�Nq�9^�̦LI"�s�4���T��_Z�6N5�r1��5��ҵ�M�EZ��z�W5ɳ��_�l��n��B�&��?��6����5�xS��{�~A%/b���@����M)��9K���i��t�|�`~�WBƴ�����I�%�l(�/����tAV^/������9���m����3�}��7�g�k��Mz'I�ׄ�^_r"ˍ]}!�,s�p��%@Jq�>n쑂i�����M��9&hY�`bC
^zߛ���׿�]H'��.vm�I����Y�����2�y�IV�>�KK&� ����YD*�>�u6�(��)�=�;��������n�k��޲�ܛʽ[Zg���B�b�����% ���M�.#��#:<^27��Fv���h��8r�a����3�A�����6�K�~����D�3Y�GL�&xL�I���+>�#"���x�/��fVQ9Ί��C�8��r�]P�H4�j��ʰH!�c��O�v�&��l���Z���hw[��y!��	��9���[y�[#�P�f�����+�'7�^}=u�o���O�~���WO��N�i��5���o���2b[;qfK��Sq��M�"��V����Y]����L�=`�=��k�a�^.v��5�u��95�i*����V��wޒ�].�)�(��b���v�f�wS�a���v�:@����jNZ�3�s��s��1�\>K�5؛��b�ae�6��?"[|�y���ۡ']��f�6N��b&�v$h�U�y�{FP�V�T���un���7� t�7�Ce~�y𭈙���^��p���`�K��CV	���<�R:��|˵Ҵ�;�_A�盯��"aj��Ni�Ii@h �S�>.�&ў�젃�I?�2*�a���/Y���P:�Ϭ��r6U�3vk~IO3����_��W~���*�k���r��y�~芼qm��]��H+yB�,N�C̱����������Cs.�*�?K���;�c-�H�ؐ)��-�5�/�8�n��"���D�V�g��|Vq�����oԍ@��O��zJa��5���R�6v@�8�X��'Rgx*��R�^�:�ǆ+�٧�5������<o�<.�a�D�3q���dc-X7��a[��EE>
�<�渡���7���&�t��k��b��	�$5�kee����gCpa�JNِOrz�68�{>=�^U�Ъ��M�H,
6�m]>��F��[�@����oLɽ����hb����S���O�l�"�����8/]px
:A�3qUG�<�D���-�*9e�k�`�R �ݚU�v�gY2v��Q��d�yS�����>n��6�=FN��Wn����hr��e ]��f������﫸Ɛ��Κc|bm!�4e�dzq���vG�0ֶ�[�9��+]��\����<_ lh�P�"��v�*P��#������{�k���ϲI���[=h3�1��u�s}]v V�,2؆�B���э�g�f��,�k��c�XB�5�߫Ӓ^{�����w��r|E�Cc��.}$*})He�΢QIzT��#�Av�*Ȫ]^��[]}����SFf\w�\��:=�`s�5!�Ν��룂��'>��
�JP�( �{O��izp���vExD ,:"�R�4f��\�Ʋ�${	m�*h/Vᓩ �%���]��p�����R�	)p�&��*���+C[��׷*��+�����z���V0��*�ڊ vsį ����"{�8������?{fϸ�V,���O�6�ߟ<�Ft������z�_O[�gm�G×��赴�i���"&?2��d�N�ץ�&�Ѝ�o�3�����:OB�y���ٍ#�-U�~q$;��)�)"73��� |m��h���ZyU� ���u��m���΁ţs.
��U��I4��gVd��Ya�Iz�����<�����5�)J1we��2	 ���7�ev�,ƐJʓ$��8�N�P=x�ʏ�vO#{��7
�1��}y�b��� =OG��ߺQO��|r�F�5d�\h�x��b����!���_�lL��﯃�}G�UȨ@ �l>�&��ސ�Thl����gy9}l��d+u�Ҫ��M\
u΢���ڛj�^}nv-��e[qX!bpb�b��&󶩅εNr�\�%C�\����^��9��⁫Ⱦ�wu��w5|�]i�]�Z�d�5r)uM<�n���w��n]r8^	��s��޷����Ik�K[pT�,]��k�t-]F8+�,V�܋��G�澢&|���� ����μ���E���]e$iU��������V�R��d��>���lWz.̽�����R��p�˲��^$���$F��Ӕ� 1�w�(�ҲTG��)�+�V�,�=�-��Ua�����G ����=0�taW�f?�LB��I'�猱ǟ/���P��|�5u�I	����x�nnpys��Mf�Bz���ս�\�׈�݅ߠ4���	WM8����z[�U�L���m�xO�����O���ז���������l���{0A4ߧ����
]i�u��ޯ�hR��U�y5�=��A�h�M� ���-P�bS�1���`�}�q�7E�?)�/�W�o���IۗHjo/��k�vT���R�#F1�M��^�����Z�u,�Z�KG�n����r^F�K�2��b���¬Fo�w�IW��A΅*���ws�_�P�����D,=Y�+��q�48�6V�^b���.�n7���N��#7�����P F�=���N%���cލ�<h�Yk2����@�-0Djh�"����#�O{o��0�Տ�=+^���Cro/�q������.�I�yn���,�p.H_�z�n�k��(�MNe�\z�$�ӌ�w���ne�x&��9&«Ṁ��0D�h�-��I\(���#�u�M�2�}H>%Ge[�������J�;�Dж�,*K9n-j�j��⫗1V�`j�)X����\ɬ/$IfP��h�����r���z7fM���bֺתGq����σ��ؿy�%�P�L2�RL*���:1�l!Mu5dP�u�պ�,�}�n7�!�;� $5v�{���#(��N�S�΍Đ��L��=�\7�r���}ӂ�E��h��>�\���fՔ�%�j��l*�t�f�t��:���bf��-'NlS>���g��G�ܡJWޯ;�yU�����CK¯�:�>�*|p���x��[��n�MS�z�'t.;�ۊ�҄Km�*'#���z*� ^$=�6�Y�H���~���;�R�^b��Yg;��x��z�:ܼ��b�V���gԱ�S�sn�?j#.��{��&QzF����t64_����ѻ�b�C���}��}�k�0TM��^�kj�x%�cu��)&%{7g.������B�yR:A^΢2?X�����SY��q��X��n��+�	����~�n�U��\�P��~/���@d^�t�E��������=����X�{kݶ
��W�}TlxQ��;�dy9W !�����%�s�qe�SG�=�᭻����)�r����UT�R�)�>:zvʮ�C��f�fVv��Nq���Y���:	T"䗅o�T�"��d�ڿ#�ub��AG�^�o�`�N�^Ї���p�fS��!U}םg�E`��J�
}��3��%���ʸg:WQ=��&��� oq-��[@��}]��WgǧQ]x`L��%�s|����Ǝɋb�y�\S�Pz����d+�D�c��r�����Q��b�-���sE�ڼ#n�^}X�},�����@\\̚��)�a^�ndt%�4��1"��
����_o=H��P�+�<�$�r��ؓ!e�*���a�8��g�.�y뤍�kr�����w�4�Ԡ�\�$���{�r|/uW�����$OOkh��|���Dw���j�nn!jv�-Z�ss���3%��k�����[~�DN%w;F;�%��Wn���ْ��F�[�L�M;3�Д-Wo-fkR�Hgf=t���U���Z���հ�AH>	+�Ƃ�󻉧���a��˳�"�^�5 HWbZ�E���:#܂^�}�Ds���������c��[�#��ϯ�pr��ƘX�n��BED[[Ȝ�wM"�%Pc����B�I3���u�@Jޡ�^�^X��PyB���\TF�9�M�G��m���8�-�+�7�0�!�2�c�p';�[����U�m�Iv�_Q��ۙ˪�!��:�&	OF��p�Z�1C7u3D�I�΂���5]G|�q�B}���uLnЧX�R<:x��s�ud���Mi�E��)+dT��f�X�V�y|�0��ɓo;A�-c���X�̕��:_]��n�&�o�Ǒs䀽evc�&��u�'���F���#���|������p���J��3ӝX���u�8�V���Y�o�e:ͣ�H���/b�ةor�Ϋ��e�i�S>��\d���%0v=Oe�]�����G6>�ane���L;�W^u�Zug�7����ƞ^k����v�k���%�G�ަdSy�у^ˇu��x2fg�����K;�능��s��h�L �ձ�,�ޔ��:n�E���p㏄zL����ٙ��1wz�8-|�C/B��*�!؝H�]�Ԅ[�!?j��P���Ø�:ܣ�,��N-�5�5�h��&�D5[��Qz�SL�}W��3���v������Y$y�></c��R|2��v�D9�\}dck,]w+.� ���b{���T�v�x���<]��{;H�}-e��·J��4})d��.�+����E$����u�x�� i�L���� ����w[��z�]+�x�Ṡ��KG:_7���q6�A38V.B#<m\�G+e�,�ޞVn=�j��n�^1co=���X+�=v)ڞ��差]u��J7p�i�k#��(�9��<��Z{�3���m������MC�i�&c�f`4�%Z��+Y&��眂��u�q���(�b��R(��YI��Ͷ;��̆ǝ�p�ˑ֓���ﾪ��i�0���}U1a���z&,>�������\�͞?]7LoA94;�8���:�4b(c���C��w�$�{��O���;�k��S?5&���yf!�0��'7��V��b}7�$�S\ƺ��r1m<Yc!�ʷcH�R�{]3Sm�cݕ�u�	d��OEy3V4������*��JI�q�:���s�j'��/�ƮfO���;/�W�]n1=�3*^�����ˀ�y�=��M�Xnzܼ�F#PMt/g�V�Si}���w�a�'�l�`�]Ͻ<0�"�U}���5��R�����힞���&>C�Xa.n��iO��=�LT���o�
�/���]v�[�v�i�s˱��n0v�U?TPXY��5xU��bm!}�S�OƇ��NA���7�?u������ /GE�jsĪ�|7��mwn�7�IP����z���n���G�J7:�YqeZJN�uC_�LK�k�Q��&�U��C���^��i�S��ѭ�#�3�B�}�慥���H���]O�\��s�nj���\��6ov�2��L=�y�k/Ӥ���e��o����V��(z)���y��K$�u@�7vHa���faC��{a�r�j��P�	�|\[�9��݁�五k��e/z��e�#��{�=֪���uʲL�v|(3D^���f��Ч�ud��ۼ�#�����on��mR�W2�s~�
�U��MS`}���b�}}����D�W���GQ��8y��:o�h���u�1�Э��oqh�L}����;2vΘ��^'���~�p�y�|�Uf����n�;����9�(�Q/�x��y�73�j�^$2X]�ԔXE�A��ΰ�����6����+Lr������qG��y��Xyq��3��8&���Gԉ�4;{M@|����ɺ�'s�-7���o�҈٫:��nR�u�SOP����x�+����IB��;|6��x�[jf/�w�ۺ#��G���1~5=]�uIт0=�'�Rc���w7X�l^)�!e7�8�{n�z�����7H�ڀ���B�u�s�����;��0�D�e�������u�<H����y��1���g{�c�v��˥x�_�$�y��=����=���{4ws��~����.p���u�-�d��ז}U����쓧č�0�u|�����g)K����:�C���=�8{Pn��FkҔ�nbr[��[;���Yu<�Z�s�vT��t>�#ً3�^Z=�	�J��{�&4փ뺞^}'6π������绶�l�qep����=�ǅ��ʽ�W2���ns������gS[����t+��
ڳ;`0Q�3�H�u���챗bn9�ؒ��͘M5�=I�C��n�@����O3�-����l�`�ȶއ)�Wd�a�*k[o������0*�r�����6R)dw�o\�1��j���m&A��W2Ju��e�������]�vU?k��7շ�'�m��\*��i�~�����,�c�ns)-���z�'3n��o�^��U��=�Tު�'X��@�s��U%W�/��2����k�g����.�7}6L�X���D���2c\�΁��i���M#}��d~ G�$���"n�Ognw��l�9:�%�e��K(4*��|��f҉��jY��i�3��z����kR*FI;�=�X��V��=R�y�H�o,���^#f��h�y�7�8��|15Dk�m�fT���-�%�hj}�'�ǣ���_��~/�KB8l��s���HE���=.�}W��w:������_)�^�ϣ[�[�r�}@��VdJ���~5��>�e�^�]��J7��}a�0�eS���A�����R���<ѷ^�_�-+�Y�[B��1s�-���j�*by�l�/�Bm�

�{euwCy��^	�tFFgu�S�yO�6y��l�� �)ڻ�zw0�\M׀��a���Ƶ�:�Y���g��B�#�����-ʘ�i�.̎��#�1aAv�`Ցc���j�o^�MU�뺅n�ڽz�d� H3:�F��L�,���g+���廋v�fn��i\�'��>X\,�wN���|�_v��v.mn�/�����!c<"4o0�˨��a}�M���9V�IP����}$y�G�'�-�l�ߙ)%t�����튥�F�Yox�����v^v.������ڽz@"6��Y��)Zʹ@��?���}�f���	����t���Z��&p�a�W��k)���u��M݋��%a��~��h�O}��{|�eD�k,���&7E�0f#[V7�~��&��`�)�������>��z��T��g�x��G�-�U��;Q׫����{{��$�He\����FO'����1K�˨<�t�^n}s;!o��C/�Ҳ�\��wt9��j���V��n�<_�rrp�[���f��y���N�~ȫ�5y����i@Q�P8����	I�HWn�o���ygsCg�y5,���E'�w��),��<tOU��ؼ�QF�o�և1R\�^�~������V�@�8ׯ{=('�9�]u��5=WU&0��Oq�e����y�A�|ײm�Z��T��S���=�:�m.�Bu��GU��I�F�RV��TIMnum��k̻����PcFu��U�6�;���3��7�n���1l��s(��*8�1�tcu�r������4���]�">�=��"sbv�g	}��۾HL�=�wжƃy�� 7>�����_��b��Q�S�_hk`�|�En���t���ߘfjL���2ק�L,����g���7���$Ѱ7ʷz�E���;�Y��ǵ�fl~�]�����$�x����u���h����nZ *���j�np�%��z�ߕ��΀��,h�Z��<j���S-yt ����<6be<򆒀&-P�n�%j�̺Z�`���D�=���y�c�Un��a@��f�p����]u�C�� ]X�e�Lzf��_�k�'��_����gJ�wް��}*�3�#��/i{;O�)? em��Yj_�-V9<�H~��B�M}^۫�����ٷ�Ū>���tUw^�����:�jv�F�ҩhl��x7���w� b�0{�Ϟ�%�z|���ӆ��C>�z��|7��^f�.��rL=���U�G?V��P�*�q&ݷP�����ꥤ�	ՓqY���5��_�!�X�gث�ƻT]#C��߆�57N�E{�B`>Q�R׏&2X�(M��#�ͬ-���"�]��K�'��{k���vt^w�ˇ�d˻dY��s+I�s��v��옷�YL�GgbX\4�.��ɥ��y�=���}z5ѝ8ҍ�JV���9�p��6�:���kC�,�[ӛ��(��g���Ŕs4�$�6RX�}l��<@��������M�"$jS�A�]gcx��՛���w�`:h�c:}�C�TН�S�p�:}�=ka��꺵�F���z�iR��\݄���e��ʃ��i�t����|{�W���:j�\y6�Q�
B��c��^�I��0>[�|���<3z$pu�rX�|�{$�.+�	an�C�(5}�	��-מS��t����l/H�=S2z�սs�s���x��VS��ܽ� �=��
c�d�=��l��<v.���F�
3������������j#Z�,�ض�U���*>�ʳ1_K���ӆ����:��N��;�H<=��o��;u�+�/ٓ5xׁ�K�8t{&��er+8�n�X�N_�]����ם�����,��G��=��f�hS\��t���A�D'�\�s!��B��%����(Q�c������o^����g?3�)�U�� ��R���DK����f��v�/��ۜ�.��L���x{r(�w�D�R�c�lN�[���m��=a<�T���������	U>O�m׏z��ߗo���+�W�=F�}�F��eOfQ �����oSa�/�/���Y�&�˺6�vw<\�-��EeF�8�&gڰ����D�L���=�]Av5&Xd��{:��|��F[Hs����@o�&��e�I%���fn�#.�K⺏v��%�{L�U|����g�;CQxl.o(�܅�����{���}�����6�h��y�����[��-m�{�9��K���)��}��8v�DIPg{q��y�u�QyQ�t�6v;������jw�����z�O����4�=;��{ sV��vv�yKޘ�=+��ܬ�v����<�~�����	�k�{a��
�3f�����6r�s�Sf��t�t`^u��{(y�(.8,^�z�g��z��;O:��z�7��]�R���(خ@3���U�ݹ�GZ^zg�Z����U�|�[�XW����vH"}z:�{ܫ$�5�&��nk��軬���9����H��I�>��k$�-��O�2�U�S�xW��L˄^.W4@ׁ������0���C��N������![+�uupWp�k��ʕ����'��y����(�*wC�=�l^`pT�/h��]����y�Ј0�$���Ĺ�����p{o[�$sB�Nc�]L��MG%������{N�8�x��wV�&=㤊�6��e�����jxt ��b��nq3�^��|Gwi��l��ov$Ȭh9.�OpL�����4p\���B
��1��xվ�H�+A)Y��!�f��X'��ĥ�םN�jſd�ܷ$�n�0�x�`7�ɺҨ^�v*

�΃�^-Pn^`Q���[��+��6l!�	G�_&������"�r�O�0Ns{x���f�:)�Sè�#ǝ޴_#'y˯kM]
�^Y�ZZW�61b��d[Z771N������w;�'��}�V��p�=�d�jy䫰�X���ެ�
���>��ǋ�7��>�]����ΰ,���^4�@8�0�<^�w������z��T�i��@A����'�>J��M����=J��
'Ǳ�~�ۺޜw���[pD�{�d�ȕ*B��νX�4��0�J����ϧ��-��^������=��ף�kp5�"�Um�a�I�y��Kwq��ce螯^wj>}��&Aܰ�����Қ��n�TU�����zd;�#�7�
+��L�xmz*�Z�x=�꾇��.��*�#.�.:�8��x�%1�3�찀����í�{�^����3'��u�ܴ�k�7���%��"Z̘kj3��@<+g!�X��!f+�C�y��U�ת�ٓ9O�
h(���v��%_�H�=�a�L�gV��R��,5� ����jt.���T�Yڍ��&�+i�l�j�h,�Qޗ�7uć=;ws\�̻D�,���lu��5R�ef3_��5<ɫ�er�<�n��1�:��ejڎ���ˎ����Y.�H�R ��%,4���+]ס~6W���� �.��|��fL�Ŝd�5a�Qp�ݯ�ٞfP���G�Ȳ����H=5�h,5�CJ�S�l���r��Vro{l����8	0��ꈸ��4A���)E~�W�����m�utO��dT���vp��r@zfi;;u����A�:A���HW>��s�����d�V������g���W8i�P{����̪�86k�r~�TOr�M� "�p:��ny��ד(�D*}wA9:�y#7�.�_�TW�)��۷g���{V�:5�Y�^?u���z�G�a~%�~P�nM���l���}�U���8%s����}R��^���<�T��= �@<����S��8롥��"/{1������ZW����iK܇��^ �<���5�p�0�Yg�����Ǩ�3}��=�}/͌7N�M
ՎvZ���g��'ڞ��n_�*+^T���$�V"F�zwQ�����tiߴP����A��y���GG�7z w:�P8���ɣ;q��Q������m�=��f@vV�g%�gn�r]l�����euEA��_D�l�7�gnS�LL��z]X�Ub�e��X˧R�V��3��:�c��1��_�B3����s���t^��{:HFf��~���=Ts�u7K��}3�Sk���Q�m��9�}_7p�Z�x{���O@hV٘f[�u��)�����f�Q��[y�ʕL�}ij�~Ŗ0����Ǖo1����܎���X���;���ug�������}�/#���i�'��y�[���[B�U[�j�P�Z�[��=9���ŋ��L��s,aǺ���r���!�-[���U��j����.{��oWKMV��wy���.@��{z�&����6�gj��Q>��ǭC~��>�+�4��q!��h���y���v��/����K��Ec�WL�K�ZB�Ї���SF���D/ee�AI;��߶���j�;�UH;Q)}�Y�U��M��z��?VzF#c��;s�#���
��eB�u�QV��(,[�k���|_��^|<:7��NI�al}�!�7S�.�h�h���P��}�!qW�=+�l|�e^}�v��X=I��7�loDĎC�,mn��g2���L Jt��X�)н���z�v�}���u�S>!�:�"s�OP�=M8���{�CIte]ޖ�vQ↣�YC :�j��U�B�IHV��̋p�D.]Y��Բ����n�dዅ���gj�Ѳ�!�4�}���-�>�~.�����ð� s�5���Dx�Z�8�ͣyb��0Q�VJN��ֻ6�Ю��)ݥ|6t�+��֨���K�>H(ě��i�9��Rf-2��_}���[�-�Szt}�o�OU�n����q�<�K��׿c'�<�2lE�i�����[Hݞ��z��es�_�����IjU�E<SXP��K�u;��������+؞>�8�����o`Q�L謡&Or=:�Sf�C����*d�z1��vS�Sd��Ʈ��s����+4&���9���/#k/
�P�ؖ��>����7����ZmH�ؘ$�����G:�c��w�Ր=6�+;A�xG,�U��ZKW>r����C�y;�
�̾��ht�N�C�����L���9c�r\�jT��QǼ�����0F�sg��Am6����p����w� M<w&��F�b���.[���:�Z�K��.;3\�k&��xv�IguJ��DHK�s��"�+��>
�<|e;�h�Agi"@���]EG1�f�6���g.���Q��o=��v:npX�\��F�Q����3+�5I<���L�^7�v� Pw�Z�JX̣pn�P,�:�+��ڋ/�rq�o����<����k'�8՞L�vC���J�3g�Ko^v�����6i�5m�˳\�m�wsX����|��s��������r�|��/p*E�4�G=�x7�i4�'�8@��|��t�*f�Qڥm��o�F�d]n���lZ�{]G^��A�u
�wA5C�� �)�[�Y>��=u�ѭE�&��kl�5lzu�w�J)0���V�Mo�)���D�ڱ����w��ϧ`�ɭ�s�X>Y�h��y ƴ'^W�<*�Wa�S�+�L ܃;w��;��-	X�i��l�p)�Dz N���k�ŝ��&�u���4!�� �U�ҭl=�9�\�y�)\���"W<��уH���NA����Pg�M`[����7P@s4^ԭ,&���+��u�u�S����tfnE�;�����������q�AQشwK�K����T�Qdp�V��x�s}�ݾ�Ƀ�ŌHa�.yɲ�q�zgIMِF21�>���
VwJq��>	�����#�xH<�f�9���vƕ�[�!fws��](l��K���ӳ�nv8��]��w?�&2��������L��C����,�
��m�̵��7bFCy���Ɨg݊�����f�p=V��b� f���)�m��t�|6��ɹ����V;��6�U	��&B��]�W ��Q��着��ޠ�ԱW�/�}>6�Ґ���\6��8Z��gʒ�*i#�*�lT�LSs�!%(���!�����sA�Ү���o_��z��]��ˉ�64�}����	�%<_Ʀ��v� _T����\�Ŭ����|��K��p�7QP�B���Kd��)�X����^N�v�#G��'��f���3x�8��y���fiڇ>r ���z��A���#��|���s�U���x[*ج�.�1f��F�s�Pp�:���{Ɨ^�� ø�` z���<Ժ-<�j�yb����%ƹ􅞖��P/o��o����RU�e*�L��w����.�N嫛�^I�V��x乊{�6��^xƟAW~Џp\������i1t=bD����yA�\M�ϥǷJ�.�dpl���`�O�l3�½���uʼ7������$�f��н�c�2Q	X�[u�A����2���;����3��5�
k��옼3<r�%�~��+��~O�!��7�;�B���5*.�i�>����;_mL�(p��
�Վt��F��|��[�!�#>UjW�
������=CW���g�	"[�J�#<+o0��zF��j��Stv�c#�1={���A�S��а�u�U���7V�9���fw\,���5�]�{�|�d ;�=�'l.CU��6��g��q2S��2c��VQ��:��W���6��9�d1�Jd�5��l,SWn2/��a���FKC��Q�L�^y�H�����_�%�ʀ��C�K/�8a�wg������~d_X�]/��b;6;�}��~�!t�*�UpH���6�۔���3|����f�D9q��$vݤE���ٳ\W�Y''��~��̕sQQuo_�8�zM���#�Fnϖ�oJ��~s����w�V�߼ekw�qVwp#З��R�nv�ޖX�5��V���I���#�Uw~�1ѓ:�L���޻�ǝ����}�9Uػ�k�n�vk��
���|�}w�b�:�!f!��ۯy�\1ew�;�t�u+ݥ��u�:2g���'xo,ұ�=yҹ_&�5����p�,��
�Amw���@��/��bs�u�e�~^�\�{�s����"�~�=9ؚ��[�,����u��]O�[�xWZ{.%dҳ^?
����/�X
X=��7�{6�2�s��:��a�����E֧x@<�2�
������D`��VwwZ�]\���дz0��9.��XmM�� ��uȷ��ܳӦ�g5�a0�<Z�\-3�82�޶j<y�gsyG C��O#�������2V1�����Cno[�3��D;�
ˑi�i������:�ι;s�Q��w)}�L�2���������u�RX=9��u���D���spތ�ŜF�N���m:�D+�� ;3��4כǸ�;�~��: Sy�1��&�K��S*�︤��\�xM{���퍵�q2>}���h���^<�vW�N6����/���
y�m=��}+��x\�=�Dcx_*���1��^��7Ț~��X3����`�G����^���J�޲Oz�*WZ̜b zW�g	Fخ���/���e�W�V5Y�kܼ�ï�~Q������k�e���,~�Bs�<�J�o�¸_eɕ A�s�~��ɚ}�������n��V$��c��3���~��esAZ�0�)0-\r�u �&V�h����up�.t�Ҁ��i	�1�ԉ�Yw����8^�W����}��6�R�|&ҽ�����A�+E�hǝ��½S�S��S����^iZ+��e>�����3&3��B�����<���Xv�94������ϋ�.Ў�MTU�îk<T��q�C���˽�}&��k"�|�ӌ�A��(����upkV�]���z����}���8����񈃋�za�x1L���3
�$����X�)���x���;\�<��S��ԓg";.�款�+13�)ޯ�:Ǡ�ՋǶ�y� �R��:���G�v#�=��G�rҺVְNѻ��EM#���<�$��������R�'�2)�b����;�Ěu,��Fj��@�h��V���w��l���~9��U�;�lG�tW�e�I2E>���s��VϺ��)޼?tC�̈�Q�E�r�=��9O���_=k/��zn#d�&�q�X
��+�Pp�篷�w��%�P�T��`�D�~Ķo��s���-�HzJ}��Ma|p�y��+��=��ڜ7;z�X��@�o������?!�r=[g������aC/�1�5ہT(0�d,JH*��u���w��2vQ�e�s�>����͛J��e/P�%Bd�X����A4h���ʽi��t{MW�v~���=d�����	����X������fx!Ne�TrO+��S2#@y�uM��:���A�Ӕos�z݇\�-t� �u��Y���ƻD��>ˠâ��e�k#3�:.\�nc3R�-���.����R���{�R1��C|�l��1�vekn�/�]�'��NZ�Y�^�W���P�}9���x�#��ޙo���[���sM�������V;��<��t���z���ǭ�^���쥗.�~-��yq}���u|�ޥC�����!=�uf� �=��̮���
��U�Yy�(��}��9�ע����Aċ�.1�;���{��>���=3ܦ��8,%'���������b����p#({��j�乱����˒J|Oh�5���X�?x�Tnis���7F�+�����^��)��)^Ϻ��<=�T�7+��񆌋lr�wr�b��(�Vq�y�[�PdW$<+���Vd�t΃c��f��G'�o�_�V��Z<�%)E�U�a�����A��jw)iZ�{B�d6�{�j�=\�Y��J���ϫ����}e�����]�+:�:Y������ʐa+G7��.���)^��:}�m�~���-$,d��YJ�w����=(.��I���`����`r�Tt�u����j�ռ�T�1��}��'7:'����~1:]�'��%]�3��٢⾚Sm�A��U�|���!�Xz�����,�^
�vݡeq:�co�u��z���+Qf��h�k(Is��L����r�}����tH�O�_:Q�Wg�[
ov�ame�y1T�GF0��X�o��a�R�i떡4��JK@�:Mp�;*���^�;�:){;Z�ZӾi��h{�w�js�]��EwΒ��;9oe��4
J@p��o����*afG�{��lx,���{T�E���?oy��o���`�4w��ut��.b\<��r#�7�4=��<�r\~����x�5��z������Ne�-�=*����P���o�/<����b��{7��,�t��Ofg>�_M�oN
��d���n�v�1�����|��PR(`�̝9�է����2���d�&��_F	9TH�|�Z߄���g�3u&N�^_�������|�m��hFC�3A�H[c���W�]�j��^3/���n�Nj@7ǘw����o��M�����"�wЍ�rE��[��@ֹrj͡2�w��I�>�>Z�EX����gv�{��c�b�t᧒7{i�V�ν+3�f��Y��v1���g�t�s�"2���WPD��v1b�����L��7�[KАF��d��G�r��ʲRZ^�/��{T��Y�\�u=�����r	%Y�棤\��i�԰�@zTo�g�y8q����p�v;àY͐D.X\��t��.T�}�&��I"�1}�˷�C�I��bh;Sh����;��� �Z�J�3�����Ғb�0�e����ݶK�l��������"�nVo��Z S�x�M��Vv���\}�&t�~�F�i;�����5�&%���f1�kHˁ�3��4YR��o��ײ���!�z����w�C��X��h�/I�2��6�Mt����d��j�S퉇���>���)���r/$���y���y�l�����W�'�;�+<�y�/a�����c,y ��}w�Ie(�9����m*o�'?y?c+��0��w�VQ"i��UѲ�uwZ���lp��}���v"�dpvT:��xr��̥�ת�6�������|��c����u_voZ�J�Q�����^���sr�R E�W5�kg/=�tνL�����a�׀��̮<k+�����Va��[��p땄h���}{ރ�C9R��m{��z��5&Z�Ò^��C�=�|x���m�8�U�����}r���ll�tA�;r$jJ�*�]ʄ��ͭ^OS�K-�Ecy�9���}�����g>�1_Dk{���)pj�x6wUv[�r���X�H��ظ>�:
��˗��k���9�)w����n��Y@�f=d��g������W�\�I�֔��1�����|������Tw-�����T���ב�rO`�MSB�4���1[���]����'F��a�9��<�[���O:���m<ך��w��������k����{ػ{�3�^U���NG�,:��]Y«t�s_�:���n��צ3D)��S�f��:���<��������|��<�۱{�o��l�]�܇ی�*���<�{ؾ'� x�4�2�~l,��]�>�_w22�fv쾮Ŋ�N��#�4�5��2[�svf�mg�U�l�����:��(�k���킆H�������8��~����L>���d�W��^�
H���R��5|�9��V�}��t*�8�z*�tө*j:A�*���;�Y���n[w��}nuu0I�#�R�]'��l�k��9�����*������	LH������6��6��xw�;�����Q`��]b�����ݦ�E0pL�R��ס��a��\88:���]��7[9�Ҟe	��2d��7[=��V�ZOp�%�)�6s3�|�_�ei(���9c�W!+����;v��� ����֧���b��{ʻhm� ����HG�G{>.C/8�s��]N���3*7�e��G���o�Ǣ�����ڳ,c;��n0�z�-���5���qq�o]���כݾ'`|5�s��M�b�q��$�*��t�ԺM�`R��!����~�2�#�u���:�^J��út���M�.��V5�e�=�x@�Éۜv0�)_O?xoN�U+����a[v	�ܝ�p٭$����u"�hz�mz����~�ۿDЈ��t�����o��}���#�o��U���ݹ���ʟ�L���F��>���{��P���(((?��mF���~��	j��\��xt.��N�)}���*�nY�����ywCˁ��/�.R$�dS�$�%�0�6s�x���������0g�ɕs8^.��K^OQ�;����N����.�I�~���䋺ٻ*�Noez)jXdzeNyjo%�,g�s�^V�ot�!��J���x�!����R�>���fE9�1#��'^v+�����	�"�Ԧ�^�}Eс�������r�4ڋB��c)\��R��$���_=�߁ٵ�c�_�toE|"������}Y����\�"Wd��!-.���]������#�Z@��@U �O�ø�N��B���\!p��jJb�u�d��Tr��\'�PS����԰ў��Q&���ў��F�`�r�a���ø6��ظ�S���?��yj~|�f���̔M#�&m�ד���#����_[uڤ��Z)d�4|�����Wr~K�ܕٟ�~�痳�.棫�$�Օ�\��.$e�[/=ZM�򍽵���� ��GŞ��V���u�����T�\v�+:�m�I�}AJD�vu����(N�x���������ek��K��W�'v��:�;+�9WG�?NE�*�D��.; .�z7ʴ߻:����oz�~/�AW{��U��i�)�q�!X.L��,��� ��c��u���f:�_"qg7ʣäU&T���>�M�E��7�*#?/�5�<�����6?o+��lCU�Bs��hZvف���/<%f{��e���L��B�D�?m�c��?���n�t8��<!��U9�z�i�o1~7_�q+��Oλ"���1�$�%=�-�צ����EX�_G�� �xF���V}�q�L\��e��<��;f�h���
o%D�u��������4=ۥ% [��Q?��Z��L��f�̏)���=r��v�Lc���3w麅ހ�檔s\^�������F��~�B�
��V~�V�g�-O��3�PU0bl��8���?���=�M%�}����W^��#�:�x�aab�-�G���C8������RϞ[y}	b2�Wj�l4���a�\	qC�m�=��rN��v�0!��Y"�9u�C�2i��3	��wM�kk�a$o!OU����n�=����7�@U�|����c}K��}����Eaw�2<�9Ҡ�o�M
�&�#�RH��^�;hd�ۉr5a���ꖙ��1�{Ǻ\�ɛ8d[�ԗ�jd7Y"<.�L9�M���⩦���۵E.����h�Wq���ѝ�Rm��&�K�ڢ� $��`e�o�L�����^:<�G�5݆9�r}��Y$v�d��g��-^���Y���%!�ކ�w��\:���R=^�p܆�r���l��0��Y�������/�>��n.�xji50+���od]L��.�q�]�W"�����u��Y��7�]��Y��ׇ�e̢=>�{�1�iP���/ON�;ԩ�k2Q�E�ct��&�����森��KA�ٿo��enL|{�h�s���78s��b<L�t/u�O����5i��@��9ͽC��O�h��r��M�Źp6V�M[�+����Vɼ2PѤf`��U���O��3;Yy���
��s+|�z-����ë��$����m�^��#ՆĽc^&��[ԴZ����r���v��y���U�{��厰9���Ƕ���F)&wu�[F�U����d�α�;Z�;4�J�q���T�S�j<�fl�5�D�cd�4�ӶvoWs/1A�ϟF�<߸h��_�>dZV��
#ޒ-���ur�j��7���%Ҿp>�ࣛ���P�i���4�/1�@�F��/q�J�(����Q���#{��fZo����H��{JLԐD9�N爵C�y,����o�3���5C]ef��z�n�`]�4̬�[.sK7s*a�nQR�h�!�Z��]G|T�^c��\��ﷵ�ۼ|Y̩ǛE<��!Xh��/)x���w��\t�SI��U�Jmfj��� h��z�];p1ͻ��ÃU��b�ctk�ż�#�^
b��*K(rh�h3��+S��8*N��&����KF��b/P8��:�g�:�V$��bm��kV���Wd�:�gٓ��ep���֓�G6f�6����[�G)���t�f�Z��I�<�.��P՝�w-�mk{�o�䤹<j'j�t.�T^�]{Ǡ�y>�a�Kw Y���n�6�X�ѭ�.v�^�}��X�(���rg����Ú�/�򣪎��"N�A���(�5V�ء����F)�|K��P�z��Q�]b��<��N�}Z�7�b�ܔEAͼ���Jl���r��|��έ�)��},��7� |/waʋ�zEH��,}� �y��;H?� �fl:�w�D��������>�GV�ާX&'��c;4�1ˮ&���'�u���mZF,����;�混|�`�Amâ��I�t(ytΩ~��9�J���#���K=�*p�}Zn��d���(��������^�Q��.���DX��$V;�dMg�ӡ[s�n_+�31�ZN���d��X��ri$f髯�WQ���X]&��A͏6�t�×8��G��Uw(��gYy��� o���0�z$#���EDBS#�v;6�*����I�4��ZK�,�9v��#v�8�O0W3o�͚�9�=�}�FuV��W;="k;��B�OG��R�0%8޸�$�n��cw���6�[͞���Y�ӱ4�y�ݳ/5na��O����V54���A��Om�Cď]�|�m�u0��n3��G�1�}��`���u}���{쩉'Y��f�ɥp�G?V���]U�'Y�~��Gi|�O~Op�ͯ_mz�V4Ϝ�n��W���?�2s`ﻦ�cx���M��d�ّX1�]#���x��K�x�G���ox\_a}>0/r����=>Q��u���0x�QX#�����l)l�R���<��({i�\m�;d��k���o9��@�dYX��=,��nːy�u�6��\Qq��r��z�y8�o���Y�����9��ѹ��hl!�+�,M�c�_XYV��b�M+��KK.-����v��{���8���Nھn�5}W��G���m*��;kF�W���I`��|A�==�<'�-S|x��+ⷦ� �S�7[����Wm�|���s����uI���b:�����x�F1��Y�����e�M7�V��"l�̸�+j<�,T�ͪ��윯Kϰ��VZj�B�S��쨲���؝b+�p������V�{�@9F��4"�����^�u��H����=����������h�1_�D�)|:y��N3���}�w�:ƶ����9]Q�&������O��i��3 �A�ȩ?g@�f&��e=9�CwGՃ1�j_-���]s1n.�Os64����z==ґG���r�\l���g��,�f+����[sʣ:��xN��M���NmS�f��ў�Ő��O.� �l���eE����Y���ث>�'0O��q�X�d��	��غDs���ӕ�֦�Q�N����dw��'���lI��k󕺣��!�u�zX*Ϣ�b*nA���4���s�z����ۂN_[끱k���w	9�Bwj����!y�q��;�;U���x�eҖ��o�迢�S%�L{6�56'�v>�כ�'|�s*�5J��Hx�u����+�i��+��ȋ�;��<1�#�D}.��>���_�����f~]�X)oar�������(�u�Rc�4�E����ō��;d�U���vC�5E��V��Se�������m�1x��_.��f�NE$����/3�d�QwU�u.YdV<0]��K!��`�tE�&v���a�����Ic��O����։�r��>�n�,�o�Wk���pM�ҹⵅ��UoB;�|�mgt1~�H��O���]��A� �W�{�%WNDB͜��ŝ�|{�o�G陲�:�tL���q��U���{�n��)T����V������j�0R̈*�8�? �ي�{3�R/|um*F�'�'<��1r�ʞ�~�N�V��{n�$�U����{+�%N��u{bwS�	P�XqDly7rk"��J�:����w=^J�Sә�ay�T�(��q;�;�Zu.U�fY�إd�G���;�]�~��4uK��ֵ�[�#���#K5Hw���ӝ�&9�b{���,��7-���fX�J���4T�y�q+��;��i�<hϼ���#��C4*^�O�1(�zshI��,����wzׂ�o0{�i��.G�΀Ђ�8�]���wT"�>�{�ў;�?��_%�y����V?��ܫ���]�у���虪"�7��("�o��]Ϻ%�N�wb��י��^����ht��~}�d�����f�Ƿl�w���J��c��!��#����_��tLV�+i�_�
�����ʒ�0Hǅ�3`���C�|�Da$cQ�?�����N����M��mB.�ɺ)85��+��y����2D��k�|�{��іu��8ܫ'ek�^�ږ��t�������fս�J�V!(.tE���{|�d��lya"8���c��:C��{W�*F{��]����]�^U�8\�Ъ,�X�@��
�#)R�r�A��%}m�~���}��{���&�Vp'j�<ʭG*:l�D�yꨃ�ٕǂ�Yϓ�Ƀ� +�s'����5y.���������E��+[��y;%�]����Cv���+g��K����t!8[|_�ߦ�ѐ~����T�7z�?I��V8�}�l��1��7����=E������MX��*���\k���ڷ;}\��cW�7}1��ݙ-i���+��N>��V���N�(�dj��w�o/��K��׍�r����r1j9VnI'~<w#�D��ƽ�3E�3W39q��2��hWd��f�`��t�gwD�i�����?��W�GS�p6"��>��)�2@�(0׷��VO������WV��Ҹ�����}"�#6��2z�.��l]; 5���,zK�=��*`w)j�N��Vi��o��=�7r��x&)
�����fK�r���9�B{+A�a>J�<��<;p�	��.��j�na$�z{�����6���yvzc������ג:��К+��2&/a`��5������i>����Z�3��zW�u�,�f��Mҷ�l~��n�����0���4{f9)�}f�f��N���&f
��xb����`��C����k� a�#�&����p��>��sOku��MQ:CbT.l�V��L���u&��͜*�7�*�������[���Y}g9��B��xp�΀=&L+�e0؊�N*Ur"	�[�\.7:������6�����/�wp��=�
�l��Bps����y�70U]���Ζ&{"��:$�P�+se\O���Rڳ6���IQ���yG���۟G|j#H}�`�Z]Q �)�����lҭɃ�$���n7wD*�T��"��nN,�\�"��цcKMLZ�{�N�+ԉ���b��<� p���%>�ˁ�������FU�ڛ�2�{ܑ>�غF[דU��)]�t�ܼpfu�G$Y4il�n]�4�H{����Ԧ���>�P�pG���	5��ו�&h��E\����9{��.�^T�B�|ph�Ih�tˬ�O�J��U�\��
��)�qڲ�c���LcF�Z�;��夐<�.��+:">~6.ULOB��:*46�V����y;���~�1x��QB��;�5���(<��9�A/�-�W\J��ru�����j9`�����d��r53 ��^S@d�b�}��f�����߻�[��u\��hd؀s��=seO�W���\��T��c�:.�֒����n^�5xj#��HJe)]��{&¹�]�Ξ��0��������cֳFnD~�$��*c�'�u��u��Ѹ�`��n-� ��pk�!yn���`��g�O
��%��2�L�-�zr�1���܅�ٮ�K��[��e�޵���߽����*�!}q�y�]s�ۖ��+��t��YJ$�.�yߊ"��]�vN�OT�ڢ+@1�]��g�$�{G���g��X�0��T��h������e?0j�şC�J���Jf7`��Og�:�~�6��G�>�<x����^���D�'�4?~Y�R9��;�}9�
��5M��`CX�h��VDlv��؉���<Vl]�GP3��gxW�A �#�v�Z�'3R�ř�gt�P��lN�or�a7�0R�t��Inm33J�<�?D�bϹ@�)�ỵ[�^�o��l輝���0b�Q{f;Rp��R/r���	NU�~�_����9R~�mn��������Q�������͋��qwQ�zfn���<����\�l����i�F-ݽUWP���k��{�uQ�����Up��Я��Iͨ�B�%Iy��1̖ �e�٦ϗ}�.�%7C��Ie��{\7\�!���eˏ�P4�M��t�(���4�޹9U/3�kj �b��p��^`����_���v!���}��q��0ߖ����uU�y.�)����:)^����G/�:9�Wk��Y�>$���r�P�H��;�Kc)* ���ۘ_����S��'N���MF�(XVh�w�[�\rm�ΜC1���f;=E��a��`c�Nt[N�]Ҷg8��/A���l���)�s:wI�������@:�9ӧ/�A��fX�q���sk��d�hA��Z�)�3Xu�*�t�Z�D�ʯ(�{����z�B��,9tY��t�߆N�	�=�~�o�3GrM�DQy� �o��|��&���j7���b6:$��X��U������g�7�ol]���}�39y{��B�ǜ�J�Ȗ�/�-�J�i��HΨcz(E�yT՘�������^:�H:ə�1�r���Ϋr�~x�r�Vk����]z
��ٿAϮ��o�S:�\_�P� q�K�p�2Y�2�����]��c��r[3�2�q#X1�&X��{W'�̼���9O*����/��|�]3�M�`v`�����M�m��#�z��Ru�Fg{�T��W�
���x���7x��&�h1<�����]K���Ի��i��s{� 0C���v��'.:�`e�9���q9}^�#x�b~��٢oa����k�c���v qxͩ2y���aLu��2w�ў�3Qw���B���f,OJ�	~��_^|�m�%w3�t�;�fU���8V�ud�a�{"V�*�%@Q]ꃘ�GŁJ5U�wC��k.~����S
�g�����=��f��������~��J��o:ߞx)# ����Q8��gsb�F�QC>b�՗]���.��wPs���9���e�A��R�V������u��r�n�x1-��2��f�vk{ok;S��<���6�u���^�vR��}7�N�+mW2ND��bX�h_�B<uUw�NWw�_�7�{ToP��ZȎ�C"k�ǎ���5��{�c1����EB�k����NJ��U��e_a¶��I�&�*�bRD��s�v��G���6��=6'���nEp5��H3��J�H�!�[`_��5�$�0;����o�_	����\�X����8]I�xN�:�\�N�]��4TU:�3c�lGI�QZ̜%o���ˉtt�s�GGE?m,������W���-���z��ƣA�ss�
�OK�؃3����_��<��D	xi�^�(���!m�yrR")�sG᧠�Q��%G�On���B�,R�26SS�7���y��ؽ�.�E�xW�WY������γ���:��u�؀GwL��}����Xh���J�{�$R�Q73��w;͗wZ��}y�+��ϻ�K�]�)��_ꞷYϊ:8�����X_�
jw�m���vi��{;X�DB^�t�^Z�D�˿yk�	�s}���4���4�ʹ=�hW^�����0W6�H�ƺS'}3&��Qb�.B��t��+�g:(�q�>�V�� ��m�x�W���ۮp�wq�Dv�������f:1#�p�`�ǽm��791ٷJ{^��cHفZ6�Q�c#�F۫Z�� �#�w4�����Su54�G.[�l_έ|�Y�	/:���1'�@	�W-f*!�C���3:�\(��W�ȫv2������S�Ssj�nb��� �6��ME�ڶ�{ s�1� �~%�.�J�����n�R�Z�I�d6Oc�y�.�A��;�h*��b�b��]���'{Ƭ����Ѳ߃�(�.�]:ݎ)�S[�<ۀnݮ�}��Ҡ��\�|��^I������c��|��x�Q����*P��(2�j�UyuV����ٽj�x�^�n����*<��5s���s��3Z0��Yqr�^߻OVI��l砨3^����7P/��R�m�xt���n�15\L�B���#=��1~^x�o�\�B�ٓ�9�^�6���*¯�WtD���j�	�ɯ�D������,��B��=.;O�l��m�f>��}�E*ר�膎W�r��3b��9g=`p��	���L�ï�kۚS�7٣"u�X='���~�<�&(��D�E���ެ�:�~��:�3pr����M��M���AYʄ���+CÄd�T�
�uu�b]H�w�e�rDz.+�Ԫ�X~\����7��iqfR`��Ig����0�������~�M�˥�����^�$p���W�U�j��V �H��I�m]��p:x�Q1����w�bLr�uv��I.�geoD�>I�m��"�,�|(��1h꺂:��z��֞�!ǂ�վ�\���f�Q�QP8�p��~��1����+Vtu.�^�ܹ�����A����d�u�������w��)I�Mp`Ni\Tպ��κ�,��J�@�z�ӄ%cݮ{8vW���֭�Zĭ����2�>K�Gu͓����D>Nv�s�ѕ�y�s��M3�rQ���y�󜺰���]���0�34��Y
0qs��֛[n
�ezf�hygJ/دj}�t��wD��u��)w'o�.�����t�5�����u��k��ҋ���:�w�,5!Y����ܜ�AmƓ��{���ꛚ�'��q��^���.^��P��"xT��eA��]�O����l��f� H�Hm�����I����߳��K��Jty��i�N>}D�j�1���j�B�.��X�p.��G���l~��+�]�
�Ad�x+x����������Qy*/n�efK�"�)���݋T%鉆������%��:��r�:���y��#K��f��K32��� �.�HvA���=L)�7-3���H2��2�ׇ�����O,�B��~1��J�ק`���K=�^N���Y����<�H��qjU7ß���F����ݥ@�L'��.�_��c?v�9j�+Y^^�O���+!t`��a��H9���1]^��@��:�T�t&f����`��c��]�o}������e?��<ߺ�NW#�_���%�&/���6�����"������r�W��&��}Uo�ڕ��}�S�qJj1�k5�d`��EC�p]�c#R�jp�Q��W�[d
-ۧYcV�
��"���e�J����O{�-�O��.b��UO-`��+��UX��>�%��g�&!�<(߱�ztV!�.� WN!�\��k���v��J�2�X��F�����i$�Ņ���4N�-�xQH;M����x��v��E��^�Z�gY�ﾢ>
� �x� ª��]nn��XXOP�B������|�|� ���2�^C�8Uv�)~��F�U'T5*۬`p��H�7\UeK[n04�꓊�������N^,[�:��Vr�!���<�f!�bK���1��X�ufdUHA��0���m���|k z�y���㠴#t4��DY<Jc�o�}��ǋV����֓��D�e}�������1��5�	�%��7��O�.u�����,��d 4U��-��ÚQ(���ۦs4wGm��.t�����+5\���N��x{���0�]ի���7)��Vc�Y���e�S7��|�K�d����^f��$�B�<���&كɉǈ�f��/80�%ڐ���]�r��խʏ��|KXr�|q�/��h��m�Xa-K����R�2��I�J!cKV��VI������v>�{�ȪG�` ����N�9�h��Avo5���E��U�Z���@Ŋ��v���=a�X���ϧG����h\e8���*��*sK�/B�K��[)�!%i :��R�+FA��5@R;����>5��'��I0�v<��QV3��w���Iud#�T�?J���=�m*�:��9�C��2�s$��K�@��fp�P�H�b��K@ ���@b��Y?ʦqК�,���y�9$۫�� �Q�i�Nf��d�'`�*b�tt`oUmԾ�T�f�0OwAH��gu ׸nѼ�{�l9�ǁ���!�Sg�ʌ�o��qvG�1Z���,�"�����>�t>{~	�je���<S�W�u��)����ZT�:^�O�ra����Qño�&w���d�b�pg�� l�x�8s)m��fȜ9%t�����Y�[t��mJ��1�Q����9�_Y�2\}-��\D�ur��Ѥ��Y��ݯQD��T�e6���԰t9��/�k��ӣ�M_d�ꈀ�َ��ٍ�u%�h�*���ɩK���[��ՠȐ�T�]NR�M:����^�\KI��[,����+�By�2����Z҅��ֶ<{v&�c]����v��0�j��p�6��P*sضj�wI[ܛ��U�F��i&��'$��ޤ�j��,v��0
�/'b⦺-��@�=�x"6����-�� ��?N�G��ܘ�|H+qE��ꪯ���ץ�̡�8fk]�A~9$�jwty��� �h��vC�0���',�/.^�ƾwm�
f�c�åK8@��zU�oQ�M끷Q2��{]��dz�13�l�n4u<��o6ӌtdǜe1��,��WH���K���V<ݬ���$�:�^�{':�N���=1��P�W:�&o�����tH���6�=<+z"LvM�����߅ VQg��AA�ނ��/4j^�k��� {��E�ֳ�'1�;����Z����_�b{w�Z�-Wf�@,�Xi�@�"+��C�EA�}��N�<����հ����#��?��#u؏q &�}7��r�o��l�&����������!r!{mخ�۾���U̓�`�*a���H����u�p/��u ^�j"����\�W�K޼��(�~�^�u�*��ov�����^�W�����^�sٟqo���R��O�6�Q����<s�^�����Gha���ҿd�q�+ݾ�Cy�/��v=�AC����\�� [�<��ͼ\�Q������mF��S]��25�8�UTU�7�bV�+u�[�����ͽ�y����.�k��m�J?]�+��K6�Ϩ��#�YnK�|)�mJ��G��H^���^�&��ב����q����α����VD��3�"�����;Pk���'���8H�ҁemu7ָ�G(4J�ڢp�O��Ek^�#[˸�\Vm9����o"!�2ӹ��g:�dUp8HD�P�ٷyZ�|/n����T�,��@ �y�⍼��[���N��]����ΩѼ�����@q��C.T�ɐ�>���Ì�z*s}������^�xM����Nn�ar�s���j�4��d��`���4*jD?t���A=����	������j(2k��Y&���\���\�ܧכ�wu��M�v�czb#�I�??W���5p��cGe�sno��@e��MH}rl�q�q!mx.�.q\�k�fj\�w~���=FΉ��=��z4x =.r��_{�ȺN��$)5�5v��q����3ާt$�nqu_Y}U�gd�VI%�Լ�Ǌo����/��>�g��' �۸�w���c�!��Jk���f''�M��R�Ul�{}(v��V�=>p1B��=H,e�2n���S,g�
c��;�쾳�������$��o
�J�Y��J�ֆ�e��tv���Cw)ҝI?��� �S�H�����>65��nz7�����@��Eg�듎�OF�3b��ׇ��[6�쿷"�K�z�A�^�>��pXݩ�/��Ƿ| Q��,f`�����Q�Ǻfq(���E��譏�L��GWA���z9W��L<u��O���c
��M��v&�Y�Ò<�C0)~�5n�� ��=E�y�h4� 93�7EO�wE-�^��t�է��Ĺ��""�pe�T&k�qv�{�31]}��-�B�XUhB)�a�G&Ȯ��ӤZh��|]«jQv����s3���[E�fp޻n>��X㢍������p.����U�bϷ'ڻ�]��FW;�����}�,���ݼ��n~U!q��2A��Q�=�`�R��+ٳ"'ޚJ�͙�L�}{�'��H6��u��c���Ts�з��f�I��[�:��E���JY:�Ѕ붸g_�x�Y��a�<�,����*�	��^��WH�[����D��� �x�{/^�,p^xG���zboO�zg�K­�o�Y�:��h�����*�d��/����T�}F�[����[��Oy�t��B��f
V�)TV�.ԝ��ћ	��[�	a�̞�yzn��y�:ĺ�VP蕛��:�ͱ^*	��)\h���cu[��@�w��ݲ��J烺Q��]q�.�{��V����Σ���1�L�$�����*�x�y��S0�u�)?{��G60��Gu�]5v5�{����ek;�秥���Q�1d>'p�������Y1�}D����:�v�G���}�}ە	n^N��tO��)G��Ȋ�&FD�&ܪ��(Y�)�w��
g�z�x��vf$�ddF�����kpq�B�@���Py���s��.��
���<&LU��ר���YU���l�mN=��t9��C�mt�L<8��9�3	�d^��:+t;K:��̝�zf�I�%"p&Z�çY�,��K$�zsޭ�X}�xgP�ˬ[ �*�(Hѧ��YY��^���oA}��]XȖ��N�e�ƞ��w���1.�;U�z���c�n��p�fK��l�s�t�H�9?\xR��T�w@���P���\D�E�]Rݪ��7���ݺ��Y
�� ��=�}�{+D�,�vjκ�v��}��ïb1{yw!>���b1䩬��7�̭�q�t|9�LDV��W3�u@��G���h���yߕ�ΈBH��x�����T���֍����{�s�ѕ�6'S��jN��ׄS��墴	��59�В�E5D��%�^�D������Uۙ��LDx�1��ɋ�+��1�]ޙ��%���5�z��>ORsǸW/PC�����{8�׆��atl\ǌUO���t,�w19T�t��9�~����;5qYy/���.Yv��͓��Y�r;�(�KGˬ���T�1ۢk���C.9
��o�����r���LK<<�\�e�^�^t��뮨�>�=�H(޸�+��45�G�FV^�8�ǉ1��tΉTq�պ�`��+oס��>�rx��7'��p��㓈��G�f���mLǫCV��M��)�M���M�^�b�æd���+�iߌy��p���_r�wA��o(����;4��A����K�j>f�H9g"'�}ڝ��%uA��Z�f���-�P��.�p�ϟt�8�.�w�����罄h���#|+���3hq���;�7�~v\:�;��V����V��J�e����XGRy^���~�r���L�Vyo���%N�^q��!�s�)j3�r�X}{VOk�o'g����}����Pv���ؤY�ou�<G������i*�c�9|�z�a��Ӵ�>%V �ƪ
u�)�2x*�]�9�uK^Nj:-�MIݺ��<8,�%��UR���g�'H��^�=���rПOh�g{�4+{���k�P1��U:*Ծ,_%*�uީ�[L.F���I�+&���Xd��g���W�z��t��=���"�{��gC�*!�=�ȝ�g� nG�����E���q����T}/~�u�z�<��tn{j���Duu��E>��5%aN{�~���a��f��#G�D�{F\�����NyW9����Ly7�[�GE�S���B�=��*�<�=5W��N�u)	u�Q�U��@f)�k�x�h����\��X��9������9��:�\k�{Ʋ��d�k�~��臏�4����7�c�U{.`�����%#��誮���"yAW���p��BN5W�v

����OD)R����$�߆mc�-�<0���m���������u��̞Z��;D�A��tL����jHThdZw%©8ki�ӓ�k��F�w��}G�u6�-wT�������;;6��kJn۵e�$O�Z�S�&�Yv;C������9q�}{]d�&gd��T����!�3��&�F��=�0e����<yn���V(껐_�H�0����v�mյ�0O1�5fޯ
����"�`Ƃ>��N���8+"����պ�9��O��)A�14cg��b�v��5����z���~���fC�ɜ�FPpȍ&����'M��Q�-�[G?~�����������7�ȇ�{�g~�n�9��oT�y��#w[�_�S����eɚ�D�}��]�>[�n�U�H��W�D��e0�آ|�^{4��Y�6��T�O�i����Φ�ڒb��[ޔ�EE	��o�%Xt=�8Ҟ�\��|�k1l��p��:��y6��ϳ�T\ȯۿ����Ot�_�f�t&r=���3�t@m�q\X�%�um�wZ�n�u�3��{�R��=e��S�ʎ�����*ja�����j�P�^\}�%׷��TJ��\�Ld�7|yW���.W��!n�wL��s�*QO��g[jOB]���]ԝ.�œ���'���ۯ�ۯ�w�,��5�ܭ�D3\�
���������Xζ���/�kAŤ^�YZdcR~����fT�k���慙�gKۭJl�� �a;j���Ԭ���2o�y&x��b���{��[�n|ڂMe�{opMO��s]`ΠO/��Ó=��N�~�
Hz"#�DǺ,@��X� �3k'D@��;���$��br�^g�Mb��֑�n���-�_���h�.����\����]��4�O���w�φ�-�H*�km$r�p��N�w_�����#(l�B�]��o
�&rb�"��W�&A��Sӗ[���%�uϳ/R�#W���t�Q�a�IćG[�)�nƫ"$��7�d_��p}˯>a�%nӉu����9\�<l���vϧ泹��zL+1�z]���n�!�*���M��a�]�&�t��O4�����ED<�\.Y61�6�Lz��ƞ�{Sw���7x3�v�g�W�k#��.�'j��5��l�;���v8�)]7ג�}�7x��l��i��vd�.v��v�<�lfMK�+uXi(|�����|"KQ}^𤃪�4�N�(?`����~��~�;(�f�Z��g���;O ��"��j���پs�����.�� ��x��T���W�����s�U�tS��d�Q��K��9k;���L��IZ�뻊���.e�r����^^QB�����Ԗ��U�tFg���צ�`P1ձ��`��S9�V�L��j��j+�6�mcǪ���8�C�^�rwт�%��t-3`_|bV�M.�2�E�Y�����K��YLt���R�]WSd�l�i�uzhL��pҷ����z=z�ᝑ�����}�G0J�hQ,��.j�G��d���=�O,m.�~"�]ձ��i�3�1ƪp�Y��ss>g6�P�˕{o��دv�����>�����`�uV�:X}�f3f�����/��	�!ٝ�ݮ�]h�]�o^�oMv��n���*=��#�+���4ۣ="U��5"��\���3x�egoW�گr�y��ߏYBf��r�Pq��W#l��<6�Þ�����*60���c=q�j{�33nG�w���\�G{�G��a6�LY1�}�D�?k]7���d��R-__�,ؼs�^�a��:�]��vUoU�J4�ѯY|V+�8����[�*7����f�(�w�����vI��<3���R۵�"4�b�G:�
c�4UՎ��Q�\?`tgEPYQ��1��>8�enE7R���C�@���A�T�#Ѣg��sivM]�ad��T ��H�LV�4��o��4�Vxi�mh�wT�Ѿ9�;O]��U��w��U�Gz�R˨&TM`ɬ�l�Oz3�fA#THԼ�Na�9���/FA����8#f��:�mz�9d.�V[��`�N��N�I^)�M-�{���0@
5�u֩N,ז{"�3�����oP��ٟKn����:�N�O1�;;�b�f�R}na���Ɉ��1n���5��@n{��{��D`Sq����	�6��?����t�� ���ӵk��<���W�ت|�6��Ӧ�1�;�u틵��}I�:��^�����uL>�G�`�M[}O�+�^�!Wрy�����{�#)C�*~�1�j�%
��xr��f0ck:���7�-w�k9�Y��JuJi��
sf���˒�0)� +밯�j�DnU�y�G�G&u�9���f{:0�����.{�jVL������&�LGU�==�ޚ��5Ð;�	>��_��ovn�e~r�~4�
:�ohb�1q��qG�Xz|4��o<I��gC��I�C͝�|�u#�	^'v
������#{2���[��qTr�u�v\�F�h��f����y;�V�����������f0ܗ3�����~�����G�ƞ�tVθ��t�x�\�����ʌ��n�Ɖ15{���H���펋�YB�R��ޙ�C��ٞ1-���F����z�D��/�ͺ�Ό@޼�:�WNlvUҹ��z�\G!_"��(�0z|4�t{%4�����yuЙ�:���AFa�%��\�Yo���X[����s�/�I�K�%��m���ޔ:�H�!��,��w/t��0C��J-�;.`���ǹt������ Gl�-����3vw����Ì��l]�oL10i�p�t�v���������<L�ј�|*-m*�+�^��,wj��\O&'�[�݁�`��Ԟ��ȿ{I
��t{V�,vi@ �<����f�A;{	GbѰT@����5H1$ۚ�f�i�&�9+���c<�C����]ǍT��;ڧ/T�u�K#f�;Td����D���FÆkl�5v��/[��P��lV��~H,�ѩ��h觾�I��$+�Uı�=Ώ8���>�B��*Z��s���=�97X����IWe����g�{]�(uw;s���/��uN���a�F�/����^R\��~˺z���8��M�]��F�`��_*����<�@��5a;:�b��+�dE���̝/+��e,��D�2�3#�}N�Q��9S�zLa����x�y��Zok,d�����x;�'M���'��a~�&0�����uӿ�V�&j��ƅ�y�r�礻��/�.yj�w�����O�)t���t7l��ܦ��-����]u���j��3^���*��s�`�>6^�j�R�S�"��n3f*�̲T��A#+a�j�U���Cۿ!��$6Ɉz��W,�!<��Ce�I��)�a����/qq�<@Zlꆀ�{�-�e_��.�m�H���.��bؚ��X�&(9�,�\dZ�Lُ/FC7T�pEy:/�.�bֺ<B���87�2P����-1:�{RT�g���y5glc�������U�#��ۢ�9K��Υ��$;��{�����LeW�T!o4�٪�d�l��C���P`5W�P¬m<�uԹ�uz�P㠺�����[���Gx����ʬidY[��˭����ܾ�௛�!�	 b�v��ϝv�����t����rd3Qy�6�ZPtu�����!�[ٔ��hu����m��k1�ߛS�M���l%Q']�UU� ���k�8�+1yik[�Y�_5�W���
�׫o�H|p��zR9C��#*���Q�vt��v w��\js�q�ȇ�x�	�W��#�Z�Y#ڣٹ�C���v�K:W_}�nﲰ�iŒ�)a�"8�u�OSފ�� ��4�P�b�B\�w�J\�B4&��N���.���Kx2R+�L���X�<�Hz�!�5�́oC�|ٝ+�ʙ�s��G���W��Vl��\�TU/\P%\:����t��� ���E������X��l;��9(�A.]��2yDWmI9_G*x����طV�%����\��Q���_��g=�ۍo�]�tO�
�U,�	�f���d�� �w��[�`�}�UT:��٧}�A=��i[��a���|��2��������/cԗ������i�JF�w�os���^Q�(�Ԟ�3a<8	ȔzwS�~c,�t�*;t��L3	We��GcWS�1lP8�+u���_�M�:�[�%X˳�do�(
Q�a�K�h���!����ٜ��vF*\+L�g�=95~��4t���x���r�3|� �z�<�w=�k�mdN���~܆���\�Q���2�땵���ͻ�09Ԩ��t����mq�A೗ۀ(�L���q�J������ψ�x����6=UO6�ќ��`ڏ:�7W�j�`��0)��2�-�9d�[�Ú÷y8��ϝr�I	۴����q�tY���Շ�/���67K೏G]Օc��щb-![pj`��:�ȕGP���e⭶a7�}lP�� F�`�j�nX�)YWnW�}P�(=�$����g&=����=QF��{��b��]�\��M��0�����<�V�4oZ�9��ָ����ªj���:��Ka�D3�doP��.n�ݦ�m�/p�
���6U��a����v��H�h=�9��ڱ�Ί����nl�J7��;��ڮ�V?�R��ӫ2���M���ݠ�E3�%����xk�P��n��y�����N�tq����&���Z�Y�d�;R�̜��*���͹�ZF�l�,���]n|CM�j���x�]B��sNd1i_u�;'^2C1N���0$2��1�փ�¢�fY쥃.1�1���W�}���T�������(B�5�=L (U�9&C���\��o�e��
��B��C�Mk�§K���Q5t�]�mH6�wL�l�M��o��}Q�R潐p̰��|�dmz����j��Z����4:�^�֫���w�
��?n�dE�I�7=�b�K�\��}$�":=}}Wwy��M���)&�"�~�GUgx�2�]G���鼊�_�c�<�Z�&�[&�7cj.�N'�Dk>��S5���U�ʎ�w:^V�s},�/5�r�W���'�2]���K,����Qb�ݞ�G�zx��CP��DǇ,򬾐'=�r����Q�NT�C�B�3��CSu��p��u��9ٱ�6�Q86��/d���6�/���1ڧpY���;�>X:�����^܄z�u=ؾ���)�8]H���Ɂ<�A<jrT��=O&}QB��.��%y��;q��p��Z�C�ش]!�֝���v'?cS���W6�W*$�����.�UkP¬�F<qAQqC�9t��`�6q^5�7�U�(	�w'�R����l�~36y�Y���+���w��3>!=2ډ����K���WΡmUzmuvM��2���V�na�M<�af����^[��o�'l���7�搼}��{Q�5��}\W�̗�޺�'����;�ۈ�&�f�owN��v�9��1�����r����T�W�v�
�l�F�Gk�LhE "�X�n�P�(�i�7[ny�$�4�*��^���S��C^Q���U�m����t)[�����j�A_q΋�c��Ngrf_����%��D9>�}~�J�Ɏ�n��g��W�
��ܟ*<ܨ:͋�:��wY�k�]b�K�>�M���U�0ܴ�Ǉݩr�w =�w&þ8y����}lŏ?#���L��}��Ƞ�M��b{�9��S���ټ#W��:ɿ��=M��s�u)�X�ǫv��`�=7��ư�6��yw�[,�U�<���!Z}C�	fcѢM�>���ϗ�{5\Izɥ�!�:mj�Y��z#�^[�B{!;�/�&���ۙ���g����pOpI�{nzc��4`��lgP��h�{��g]����i;��:��}u�Q�	��u�]_�=Ϲ���r�~d+��"B�oPJY���z�����4���k�wtB;(;�(�	��iњ����J�dǝ���t?Z��#����=�]�y������/?QTN��.�X|�v�)$z���Y�|T�� �ӕ���U�o{$�����ȓ�^��k+���`���L��7��qb^	�L�����jf:rp��*����U��2!Ĉ=N�ߪy�37l��Ww���Z:[���z:i6c5|ajFi��+7�%�Z/Onhmt��9�°<�d��dۍ���;m�^ZpaU���o�"�n�ι����w=Pu���4�ǩC��'T�.�ԻqX}f�����
@�
�1���|����<xo��(�n,bh���٣�AJe�������塲l�*A��9K��0�=����	[B�,%3�z�v�y��l���Hk=/yW_�m�t�J�ެ،�{�'%��^���fZnW'�H��GZ�s�Rٰ���07�{f�/�#TD������� �pMB�]���g�J�V�C�������Y
C�'L�bS�� 5�;�qd�����g-�5:�p@�١,垻����"�js��U�~�nd��OFӳ�=-{��7b{Mjn^��?��l��-usl������%���iÃ�4��~â�k�Y�����M����OQ�^4QO�2��3��m��:1���O/�n���P��-S�!R�d��xM>�{�W
�OM�WaB�`���o��&|��ǗAG|#�Dl��Cdpg�Ꙩ�I�v���9�}�{
��}���u��^2�;1`�\C��w��X
Z��ޔ�d���u���G������81y��v�JB{<�N�Qm�-к�W���sK�2b�^e��l��N����K}�a/~��d<��xo�4؄7�Cr64�X��!���a�̮C��e�i�2�� �9݁(�r+d�]¸o%�s���l[ϕՕY���˲*r��z�� �
��v��f��l�T�4���4䫬�^�_�q�\�Bи��2�(�wRީ߽�;;��k��EX�6� �����b�&�Û�K���!�~�Wz������"��R
Nuw;�P�4�+�"f�L�"�(�c�L#)�Mw.w�{Y^}�+O��&����)�.�bV"�zGk��1�UE�Rrd�?�.�8ߥ���7�_E3�G��9��_H�y����j:�}o��M��<�G[L�u�V����,]wW�ߙ[Z��ƀ�	���0(B�=[���,�zL1�� m���2x�����HE3�1 �N���~��#�Y�䴥5Y��ޚ��Z<{������e�D��r��ķ�1^%і:*踇�������w�Gvs�ۛ:�*��,(P�y�2ͷ���[n�_Aa�K���x�7�a�a�/�����];c�+e��P=�i�~��s#�k�����n|9����TF��9���=�~��3V�/r��e�߱m�d���b�+S��q/UЬ�n�ED�˪Ntn�P�S�40󭪛�P9�K�k���
���c;.m����	���N�M��s�����6���n��97�z(t�s������뾞�r�>;^�{+!e`�D��"���B�~M�[oe�/n���{]\8�=h9l>�94^5�Q�a�Dh&70�bb�+��1E�D0%�_���L�㫧�[���N-���熑���Y�g�^����Dd�%��7O��p��k]����.H���i��O��Q��J�+WEx�����b����FF�F�[��͛F��U)�Ά��[1.7��d��D�A⹡qU8'�f\�y߆�׮�e6]L�q�i��������^��ݳ3� �^����k{�0��9���'n�AE�}3��s's�p2�6פo�\��LW�f�sy�;,b�tE��R���?��*�_�.����y�7�8{���q���.��د#���+R	4L1�,�uo c�m�����{�;\i�r�.S������D��V)B����q|8j�꼝�eǜ���2Z���,gDF>�� �ވP��4�OD��:�0s;p-c�|��g�?���[CՃ�����mr�iD�픝�vm����;�r�����&�+�P�䔻���%��>�^f�\U{�G��J��W��s>c��? I����8�tq3�����:�yf�ZM�9�ޫ��7C�#�;1�ȸ��tM�5ވ�,vlf����c�k����l���w��zkX���:�T�z����"�V/:@�db	�}р}%�~��@��N+�����(y�����;��0��{e<8Pz����f��7��9�}sʭ�
5y����-Ih�3��ҫ�1vj1��kg��� �57� 5����T��T�*�-�;��/a��*^��;��,�=��Wf��ϖ'
�pe�̖t�!�粕�vO.��9��0�>*�zzz�0:�[$��3m��m�&#�c6�OnA=ww+�F�e��Dۡ�~Ք	�)t�n�v�I��Ὅ��:c��s�6��Ev�F砺^��3���T�4�`��\�^��2-/C�y_+��
������~^�q������"��%��.��3�d��T뙏>��Ϣ�橱y���TӘʔ���a���۔�����ל���X�~>�^�O~�}�����.3��1Dl�*W�K�w&~��zlO޵۪�(�ז{ވ�������fA�q
�z}"��;��lL9z:�Hq�w�"/�e­��dќ�;�]d^z�^�������(�C�:YY��!1N�V׈!��zom���j��C��qǕ��:��{\���_)d����A{.�;�$��}|���X�q=BK�*�j.���_�F�fz#����g�ڎф��/E��������l��{[9�*>(`�I@Dk�Wӗ��yua�/�n���W������"MwI?$.�� }zO�886f`��]D���4
zD�I�Z��͠���٦�
�(5�U�Z��e�ζ(*Z���ݵ��:� ��i�ø�	.���w�'�M��&_K(��T�jH��%�}�¾]˖��
/��۸�vJcЧw/5b�9���Ѫ�ϴ�K�_�����a��ݮ���~|��&
SO2������'%Gy%틽���B#�c�4{D�]|:wh��Gqnm���Eg��*��n&\���8������s\�;�c��%x����L�n���������߻�8�L�V&}>ꕞx(�����Ԗ#yw�g���8�z�����~�ӹg��������T���i�ccz�|4��GE}�н��n!�(���O��]J͕��[�4OL�Qͩ��o��YHɽu����X�8���{��D�)��PG�~���h�=%0K�IqjP�{*�fH��ԇ�| /���(�)�9Y��Z�R�p�N	�&r�	��0�ǂ6�2��"G��t/���Ldf����sP�Fj�9=|���N��{�}�w�Ř���v=J+�:�K�;O(<n��mگv����K���v��Twԛ��VEn�P��Z�-�MW���=g��	C�ו�b 4�����]&o��ɝ�9�YӅ��D�U��W_od�|Uulljk�<��P}MR����}�����T�e;�P���r{���5?f���7E��!�z�
���_4���΋�P��B�Dz���zC��Y6f�\�����O=\L\eLʹt]n9�@m2#���b��Pv��Bp9�n�J���#�����T�ʋ�p��ZL����n.T�ئ݆��wv�p�.���{��9�zƆ�)���85d��<���];�݁��s�+��K'Ώ�.Ǉ��^�X���f�w�M?+���&ǉ�]�"�[�1�k�.��+�1��/��_*�YQ�%����k���mD�P�)��k�F�`zV$f���=�e�D
y�r�b.?c��~���f�L�j���� �;Z��/�n�G��ik��e�I���;+/o��qj�*2!��sի�ޝ^��*q��;�x��2L,$ʺY�'g��жs=�b�m��#��^$�W�/��軔�OG����]xEuu8qL����:��:h#�X�̻��LU�V��x]nD�b����ʾ��"$<�ʆDj��3�a�d:��;¦�M7��Go����鍏�}(N#�,J��;���Ft���p�ƿṖ�������&�f�f������,�==�v=!�'G�/|[��۞�k=��̛�rI���}4GG�K��E���e��w�T&-���{��H��d�zd�y^,��x��Wh�p�쥗�݈�j3��ᄈ��~���T5}	��ǲi��=���]1,�~l��@��x4T�ۉ4]�X���K*u�h��6"�%��UM+Ex)������!�De�ڹ:>>�zP��
FiSu���_�>8ޤO5k)H*Ezk���1f�u�U�ywi �����+VMpMN��u���ݺ\�+Z�ƊW�}���0Li`��ӷ�j ��{���f�/�2׿~ƍ/��*<l�z�R2�@�������j���=d�q��V�hT�\�"��a���~��p����5���O����*���I������X�aa��5�/������<j#g&�m>�S�3ОW��k�F:M�C��7��2r����n`z�P�
�
�·<��K�v*%��6moo��2��^�����M�V|�=y��YKDs�N�Qsu[�\���y�U�U^#a~x�*�g3/ۭ�\����՝�5�<�KC��ۚ3'z�^8�n���~D�!�%&��Bfn�^;���QPژ��7�#�`֤��abo�p-�"�5:'^��u�ܕD�z����cΐY��ʳh��z���g���F{3w�%�iiK���`F�뗢+���<7]Uu�z�kF���
l�[���������/Mx�:�����w������H)���/��ڻ��aPef�T֒3b��L
UO-��A��cyy��O���6g���DHw~��}j�Q>y�����ML��� N��� �j~��!�u�q���{z�T��;b?��oT�����TN�:��y���p��ċ����:Zc��s�d����M�<W�d葇Fe��è�5=�qE8�Wû�*�����|5�m\Q3ƥq¸۷F�5WL�\	ʦ� {�<�zE���8�_�VCr�y��*!��c��1��y\i3f�mp�ĹH�q�4GQ�?G��b|�k/�=3���AuֺV��3/ӂ�|�r����v(�V��[%���jlh�}(-����!վ���`�_�e��5T��6۫�'.��Y{7#����a-M_��䷴٥���ڸ[���~?$��WY��<7�4~_����=f��*Tem6��tE�{@&�I�{C��^$��!�IN$R&v�u]��
ᆐ�v�;B�d���1�n4��]4/f���z��Ϸ�E7����x?��{Lwp�vD#Q�3.ΟY�Ϫ��Uu�����L ��tے��)܁��h�bB��s��v��Q�:�mt77y��o=��P���\����C߼��f��2�)�9��u7�(�w��1��]Ea�{b�x��@
��z����Lﷰn���]�_�6��b:��fviǣ�Ӭ������I؊���tY̷���[Ǽv�9}���]�ʱr\���\�J�}����Q1[�]����/L�Z�Ѕ�{�Oc0�LIz������3A��1��Q��N��4�x�	�)��(N˓m֮�&ٴ�(쟻���s�i��~d̂{%k�'Te�K��DQ\�S���[��k��N�<tl>gg�}��MI-��
OtWU�}�A,�E����$�l�*9fh�U��=�S�;���*;�HqՑK��1�9t�+K��wg+w���eǴ4Tg6��l^vV�=���_k#�P��k/��ӵ��9N+諭��z���d�Ӄ�A�y�N�Hf���NAݛZ�揄�9�!���.�gW��� �][�^�T�ګ��=-�_f��+�%&V����Ee��xsW$����SV��P>ߺ�|~��p̾�i�U_��r}��dE�.K��_W���%��W����z�g Q�S��7�Mq�
f������ܧ�ٹ���۫��	9+�#����y��^�\�v��,�K��&�5kU⏶��=X��ӻ���!npcd��m&��Jf��$��oU�O�K�x�SL�w����=fi��k��Qm����W�X�� ,�j3U�$xE�}�`�XY����`;]CǏ'�����k��c�Z:���K��t�X<N܉0��Ŧ�.�#DE[�+[������̋��q�<�,?>pU��1ܷõb\��6�!�n��4�����b�A���)K��)F�oc	�]ίS���.{dܷ��眩ky�(�n�L{�X�q�˹PM��7��̠�����KMẘ28�p�:;�A���bfo
�z7yկ��n��s�#Rv)�b����qu�7�	�ti�>#�0,����\�dgkVpڇK)���,c�WRz!3zQ��}Y/\��g��A&I�������s[�zt��|��t&|�;�5��s٦e�*�m(v�.�58�c����e5�k)'���r�Q�m������<�ّ���ʾ���z�wk<ˤ��O5����ʺ�{���yS��W��P�9��?>��"v���Q��2�����Vt���4�]|Q�u��Y�r\2f|J6�;ٙ7Z}�u��Ĵ�yL�sS���C8e��X��s%����X�@v�0���l�����s�o7��Z��a�d����r��t���w�wݵب�:�@k����0����p�j���uj�}��u�)ʋ��_�E��6���3�h7B#X;�͈V*]�6����ǑӶ �t��X2�蜆�D���ϒ�Wu2�`���΂ȸ�8-۾�u��ow����s�Y��i���Kl�sWmSӂ�G�,��6�h�t�e	̆W��ԋ}���j�i*��*G�Vs����:�S��R��[�P˜�i�������(>,�Cā܍,$���T�4L�8��Y�-0\���-q�Z;E���u�6XY����A/M-޲�ʴ:��3�,�7=aEc~�����X��]8�	�-r���ks)^u���V�l��.�����'��ϼ0�	����h.����8T�5�7#�������C��g�t��{b��7�żA�;�w��;��\n^b:$�2�`gs�Rv���c8����W���VJ���J�ݗ�����sl�GF����`��)��Oc2c��<�����7�rF�3��ovV�im� ���<��\|�!��V�x�M�F瘩
k�8L&�ߛ��9PN\DU[��h+}��N���j���6̫!���z4:�P�zW��e�5��Ӿ|���LY�S&��܌9�՛O717��刍���;�nقu�+���$�L�����V�n]�뷼�6{Te����%=9��G�_���#������q��s�s2(����wkV�+��M*7ѷ>���|b��Φۚqf�v������l9����N6���qCbĕz��۪��Yݷs��"��ɴufm:�ʡ	ٟ_M��Q�on�����8a�P���&��7b�rQ1샥�~�$�O��:�p�q��QJ�Cs�9��+Y�,�n/������?w0�:��+ۆGl�M��l�Z(b��N�lÓ���\3�my�C��������*��������i���J�U���z�(��)7_?~�rd���+1Σ�'�؋�aR�r�nnQ-f��^��q�7V��I�_N]�L#gǺ�Z��3Xo��V}�U��W՝]1�g��f�ߟsTJ�sbG���u�M8�K��9]���H��T�3�N1��حc�8��H��s�)�ƺ����\�a�^�Z����l�(��n2F�H��IN+kҜV��]\zܴ_���J��|��ꏖf\�yм,\����5��,t9�&���>'N��<;�1E^Y�	�w>ʋ��w'�j��ў�6l��U�����7�P��o@��|�p}*��y�}ކ�Y���w�rq���20���\Y^�wK����|ϴܢ��N2��(r\����u�јY4�n-J�����ɻ
�L��%�EO����@��Sw(�h�� �"D�{C/��s����6�0ꃻ]��ȝ�deX��})�.s�A���ɹ��ܚ$�{2ت��:n�+6t�
�W����V�R����.C˪���x��~��4�UώJ'�d ���P'o��\�v��k##d���#v��K.1��؇��8b��&���������
��m=��ޛ�������u�r��I�q�O����KJ��~��=Zn���oP�ݞ2ozW���s�X��v6Q�����s�G�/�G�?�Wp���ޔ�a$�ް��X�[�㰝���+Ru;��іU�~�ᮈ]�J��jv~��h�JvC%�/h�]Ѣ:��8<@����Ֆ^n� t��۲b��ѽ��OM�ha����J����S�w��rO�"�`زj����f���Y���`�6ՀQ�91��l�ߠ�{V%������\T#�����3��q����I�=��Y�{�Y.@뾛#b�Ԉ���1T�����{L�C�u%6pϳR������u���cf�^�p�8N)���9rl�;_�;�twY��[�OX�>��v�<��Z�M��X��a�Y�fNz"�EG<��L.�?	�N� J�N�<+4Lxc���ׂy��fM��f�w���
q;�́5{��,�E�l��a��Q# ~��a�4S�i��Qz���x͂�2"�e����Ѿ��~�\�[���m����ڴ~+Tm�Ψ�k�z�Ɵ	)�W�Եg�6q��XRᘴ9R�ӓET�:���h��J�(h��Nx�?QiMi���0���^�I�d���O���Cwuǫ��r�����V^c���-��O���D�혦n>&�c�Ǘ���+�2��g��]ڽ�s���u�{���,E�*���i^%S��[��08�4\8�"�1t����OL���Cn�w�n.U�hP�ɡm�ugcyh���N���'w38�U�"گF=���q8՜�ך!����ѱ��N���*�|R�u�S�]��W��
����b��1r*l�s6,��u�9ͬT��?�A�DN�6�Y.Vr�{���ڴ;��w���!!T�n��/V���S��2XI��j��z�����@�f�f��r�����t�����oM��rJ_2����Oi������҂��g>^·=ݓF_��U��O�gG[J��^5����l�C� �P�w%?Ua��|�������V��
�5�ƈ��5�9�sph�I�\]˛���bs�,�w�v��0.옶��9��,��xKڇ<�f��:�A�̋�^�V�E���;�ۮ�̣
�<�?�?�"/N�f�o��ҥ���􁜣Bk5�>%!�r]�>��'&x�������۞�p����:�Nh�QZ�������oNW�;����ʨ}�`ʒߺ��OMm~|���~��]��Y�[��W�Q������\���)�(���1P�+�b�I�-C`�K)�A����L�^tEtBҟ�%w�������V�c�*��˽��{Þ�Ւ�m��~�|zb}�o���O)��ߛ����$Ayf��#O���*{�s��sLi�jm��E2|��m�X�h\�k1��?cV���t��=��ݎ�I�֌�yF˥���EdH7΅T@��6���� ���#����;������nO�|w����Xv���':L�XdPm`�;R<_s׷�5tL���iD�;�[���9Oņ���H�}[� �±=*���7L�� ]۹��2�:�8�K�.^F�<O+-� w�)e̛���v��L�`:/�L7��K0͙߿#�?����:�k�H�2����=�7�G:�2<%H.�u{7f��+���̕�p��O	�����������B�7���;�#ɱTêeVlQ��5�.��̮�X��k���>v��20�f ��Q7�
�&� ��@��4M������k��k�=�63�,��OV�J����KP���9םnͽn�T���+�9,K*n���w?8$��fN�r�����f�z�G��_���7;��rluɄ�Y�735$�wB���f=��\�[�5=���(p�{1�z�m�>nJ�Ҷv��Vv��3o	�D��ȇ�U�Ԭw���s>��]<��5�A,�9^X���Y�w��7L��NL���J�0M�
��.���fbS��@Q�[MɄ.Ǔ��.ٻxi\Kt�����4n�ax�٣e�.+�N���X�=��"��:r�q@��f�O6T�q^kjz����<��	#jsz���x��mU�F��vH�b�u��O��7��Q�i��BR;��4n�*���cG�b{�&��,�I���ϵ�wN���\��+�:4��e�ز>D���\|��!6d�����!�ز���zmk��S��������ɔ]
�֪"����C����O����D����'�3���:�R��zu��V|�߹.�O' �#E�$览۷��d�v;�9��]L�^5���
����mr�2�-)�'���K�&g�Qb�D�忀��Y���\p���{�o<��2�����h^��穜�wk�^7�� 
{ >ɔ|�F�_#1���	kj��qh*ɔ'!	`�9%�p͛�k�r���Y��Q3L�=}t�W��v�t�������IcBg��WOմ27�Tf��8��z=���#�;�Lq�����5E��pA�R�ؠ�澡�d���5��7��+s���\�T˳Z+ݪH�Iw
�˜��Ei���1��8�����l�!�>�^9���W��FN(|#''ϯ��o���1Ke�f��*y��&Қޢ��rѬ�xP�U�7v�<���>W�!�
�~--�x8���̻昡��ɧ؟�"�G�/:�<�{�srN�$�+�I�W0��Ў���f��n�ST��J���Y�������3.߅�g�	e�<��l��KKjF���`X\n������X�:4������T�1N3�f�A��^
�7(^��<�w�)�l�,tt^U�p[��2��a;IWZ�����4s���rT{���g*�[I�}q�k��Q����$FF�8k�K����N������6OCxt���
L��Mikh���x7\L=��l��"c'�
�_���]�T��9��e*�����7�zVJ9]�9yB�&W���`:������ʼ��Y��ꓓ�f���?��N#��Ү�3�����ܡ^nk\�L����F�~������$.���j������L��>s�3'�vG���VOl�o-�g9u��<~�����ܻ�{ۙ}Oި�P���38!�qG�l�S8f:˪�<쨺��=|��jGuӥ�ιQ{�v��s���&�{PX�"d���2x�j��P��"y��L,��/���L��k����������Y�dݥwcs��Z$�G��0��,ɏi�j}$�B{{s��n@�`3��WR�M��V�G��n�~{��o�~[�Z'5��8�jΜ�v�"wZq��#��7�U��`ѵ��06�=�n]�;U��K��ժ�nvT�!��'ɼ`�m+�76��zk�+�{��h�x��(ˣ�sl�>�tUI�K��)�ZM�i���1t�s�&������R2�řr&�5�z�ot��9�~D��L鑯x�J{�:䗅�F���������,Y%b�
ߗ��>�.^��UT�K�rkN���r; +%����t,�x�% ��ݔ��+�e5;O�:�.9O/��e
�|g�����C2��6H뮕s-;���������#Y�՘��%f��դ��n��#pK3��˧ŷ|h`�34=���Q�-n��ެ���ѯ��O����>q���ǿC[�����1n�������ik��5Q��s&������MYF�?*�xo�l1��R��tmoh''0ȗWݘ��c�
�.�TC����dv�$/e%��7S�P��1P/B~T��Y����d�8݉�:}DS�	���G:ƌ&Gqr�*�3e-�="v4<�d��
*XW.��D�L�ާt0F��՜����R�Dj#�_���묯z����.�,gJ�ٖ�PL��JsЏz�M$�q�a�]��uZ���˺���W#�֧h��q�:�&4F̎��f�n%U �2������ҭx]-�y��CEWaX5v�gQ������O\�]�b�D��[��L�r୒�H+�:qB���T,�[�ݺ�$�2ߕx��ԕY1�4��ܹ���%/#oG'^Έ���$(06ʢ;X�[������GLa�ٌJ���ؘ�lě~Bf�$�d�s�sW@���kl�|�+ۂ+/��M󁏛Y��V��VW���V���:t-��n�д����ߐ�� =u�������2/��t�k�I��T��V-,6+)���+�ԃ-F)KN�/��SPvI3^��z��]�.��ً]*��Q�ܾ�[�:e�����ۨ�a��M�s���-"����5Gg'ڬ��a3�њm���%<.�,"Dk��תk/�h,Kc�i؄GuK���ف�xb��y
�%��^�Ǽ���M�f<��xo�=ޓ�^Bzj�4���5ԓ#EgШ�r��\�����*zU��uB���L�0��2,�W�Փ���Co�/�B-���%-�M�޹�d��:�ܜ�^���|"�n��ö���S7�{|j��g��zt�,�y�;�*�߿��nݷΝĽߗ���K=�{V���tN"�ٓ<�ț��C=8Fv18��boL�� ��N<v����J�fEK���{eF���ah2�}�����\	��A5i�(�>��0�C�<,�ܻ25�B�P�g�
�a����L���7�<w���u�j[�P3NkL�Av�lN�{���^��v8���7LWCs]���Dر����xǷ���S�Ӭ\�n�S���GB�^35O^Hr�x�Z>�F�\���9�o��#+cF�hS��뚾m`~����~��}mj:<�^�w/�Z�D��z1�V�N��X�1� �P��|�ZO+��b��A ���o�l6�~N_!��5�(Zק8-�n7T��v�����["T���j=LwbGD4�L켽�<�d�����������R�[�{���#L�B,�c���=FJ�t��w-�:&�r��*���&C;��|�TMR�z�iuw�P��ԑ��Ǯgt �򶯎�o�����=QX\/�!?u~���V�D��#�����yЦu?^Hd�͇��.�T ���CUN�4�jYm�I@��ݩ�4.��˂��$���w��}�ےk�"�{��R �2��+�P�%{��X�Ȃz=���c��3̝�kC���c�?j�ע�~�G��}�`�y����Q�kg;^�jB	`��>����&���6q
�=��B���?\���yȣc�zh�D7TA���G���3�=ٓ2�E���g���@�pɇ���|�f�b���vFW�.��!�mt�Tj�lݾ��`Wus]�c���9K�8Zxj@�M��.�[aߚ�R}�q�{������m���~3P1��������Ϝup7�q��� �џ�<7�K�ե��\tw��f�Z���^�/��k��J���@�BC1���'==�h��D�C���X]M��Q����T=��4iF5�������A�����ٵ��y�
z�;Ͱ�����.����WK�m�7B�B�2�Vb��r�A�`�)k���������V��=]��cH��{�����2S/�;�e\�΂�J�&�z�b:h�����x�Rت��&�=�:�-��f�4��{��q��x�ZJ�B�¥��m�݅�ǌ����nJJ`l�=]*f5���oa�W/;�, Zʓ�m�T��VX���8�9�g
��ʅ�1N�y���U8�󹽇n��AK�F^e�t��o%`ZO૕�w��-��"4��ßJ�o�l�w��5M5�]�֫�xpd{��H��7��x)c/�@��f��;O��MQ��s���3�M�ۦy��龻X�q&/jCGj��:ݽ�$���"��6�[BD�&�X��cx�¬�u���Ma��U㊞ފ��v�nC\���Zs�sO̲�QKd��pf��N��D��oX��+!t�G-�:�JȬ�.�!Q=\�|�=a�������K�F����9՝c"ޗ
�A��RWE[G��kn�NE�z��Y&ub�9^���t�V����M�V����m7����W8Ś��8�0�'1�Vl��f!�j�8o�����'\�!��ɻ�a�P�xa���r��5tNL[Y�Ic&К��Y�6]#����H<a���yQ+����FO.q�y۝��+b�ī���j���T�w!ѽ��d�פ{it�ݱ5k>k0&}�e��P�s��b��iצ+}�I�͹{8NIf΂{�e��v��6���x򴄀��xW� �'+m��Cu�ًT�%L���u:����ԣ/���]�n�n�h��z�Z�8�y���Sնbh�L��$=Х�����5V�g^8��V� I
�K�뒲�6\ujMS!V覬n���Է//�"�����CC��*-�o+��5�.ANwZ�lU���eP{Wu*m�ާ�ϯec����]�T���ggί-�U���kNa"��c:&��_&�]84$�;lY-#� 8V7َ;�S�D�p�I;@�]�=+��N�'Vp�3�'ҷ�bw��v^f+�f|�R]�`��7+i_Ph]��-|�n�Ą���*�������h�q�V�fu��ʶ�w��= �~f��|%i- 3�eڈ��=�e�w�l^�)Y��*]��<��1��*�E��n�k�mȌ�mj��{`;*f2�GY}t�������`�����=�X7�-�q�V�z.i��޴�{�6g1��hY���_Y�r��`��_�B�!�UtZqV�����`��F,.n1Z7n	�ț���3�!����V�و��=̓�M�*l�xo{�=�nU��y�V��j�m�e����w��0sW]b�\"�\�;*���n��76]EQ����V��9S� T�z��F���fi���,����3��'gF{��c����j`�z�ⵊ{�D�lnE�&c�j]���s�����Vn�`��'H�s���w�_m�(J���ݹDe�Ю�ܢpQR���?Ϫ���(R�sk,����L�$bڕd�)��Gl]��6���qS�{���Ȫ3�[��1`4N�73��NiΖ���ӥ�yk������J�"m�Z�!��nP��l���\qo�I��?����f����ۘx�����Y&� F\r�)E�(��t�_�i5N�r��JV
b�\��Y޷'$WgQ�7�g?uC�����C�(9=��};kVB%�˻��%��L��ĝ{.�r�Zi-	P�#=�E��q�o�V`S���*=Zy_n��dtJ�����:!�ȹ����N��r`M%��E
uk6�|��wPk�ۯi�l34U��ދ�n�ω���ƀ��J��P
Q,j��Ѫ�Kʫ��Q��rXtTxJ�@%LKoўs\[��c�$ټ}����G]��0|{1�˩�u՚g{ T���Ƀ/��̍�xs'�߻ձ�3��$�<ߣ�ǙFЉ�zyIZ܂iK�ʞ�䯎1z&������������8�~f��;ɲRn����^.q�\�o^�����1�R���8��F�5#k#�0Y.r�Y����4~����9�7~�9t�X�v$ŌW;Nf�t6�a��e3�za���VS�e�x���W�A���.#@Q>�P~pi�(Q7�S�.|���o��d@(�P��ݽ���TtY�6�=]�+w>�Z{�	��4�CѺ��2�5fj�� oX�Ǝ��Acc�uR��嗳x�[�������6���ef`�������M����O&-t�t^P���eױ��)y���[��Nz�����e�C$�|YsDc<�yonFw0��e�G�s������<�߸oD�ު NԹ��q�OB�Ւ2_�W�^�h���x�;.��w���z���E�����֪[�/��V[�a�1`���u�X�̯.�O�2�h��x$`�l��5��N�|�=\�7��{��,���ϥl�9��� QW9��j�9�C�r�&Q�ܲ6�:	��onϔ>{��p��œ{��^Z������2�n�z��~��dJ<�vx���b�T�߮���1�.��4b�1�⽚d-�{/iU���SP�"#G^w]ȭ��R�2�wnM���LY��WL�����2Q�
ტf��m�͗¯*7��J����ֺ�B�l�댭uB����<w��k��`�\{�Xj.6&��)Z�n�H�F�h.eQ�(�j�\�S�/����P�c�����8J������<}�mU��l�^g0�����Q0�5��+�2�\f�W;��
�w@n���x�Wf�$h{�r�9?]�k	�<���Ս�3	Ũ,��jw��bs�{cc��x��{��wI�O{�!�F�_w�m���«��6���p�4/�=�5�-(".Q$����CZ ��}��س��E
d���ڂ����Q��wG-/����>��|�0߲8N���� y�P�( ��*j�������7~܋㒑�]6dL��HT8{�]\����(tF�fnMzzK؟vRNn�����o������{l�|L��������)�+����z¿z⢢�oA�G�sѳ�h��6�;��=���*��V�ש�#�!��.��h�X}�\@ZsqΩݷ$�|�l��dK��Y �H-�z(�LX�`^��J!鮧7��6��&XXL�P�^��mK907W꾿����G^H��b�ծߍ8/��=����#����t�<�3l����}}h_@�ⰨU�B�2�������o��_�w�c�a�H"=��=O��%Fe�;��¹�^iH�:���ǝ�e��}G��]7���k�A��d�#��RM������xD�d�g5)��{�O�Fx���G{�!�A�ۣ�>Ӟ���4ؽ�w(�N;A��U�C���*�D���q��rD��$�#2��剳P|4TV�$ۿH�MQ���*���4Ӹ�ɇ2���UxlE*�_�"l�L�4��V�ӷy,s)Sj*g6�x<�K/4���k*��r
����(�	c��͆�6m�(N�C�բI61ԻU�����)m.Y��4/���Ms�]�t*W��в�!ID-�%����΢Y4wB�ſsw��Nf�&@[�7˴Y��U�R�+ݼ��Ͻ݅�d��c��H�d�g{7#�=�8���u%�]0aOp9�y6ps�5��׍��˄�׹���`x�ǖ8�����6T;!*�T���rPv^�<�b��������x_��q����_�-�!�R�h��tz������}в�Wa��ۇ+��d�fXV��t����� ��Xw8/%�~�Mn�r�%��*��a2�0&�zĩ1��H��lfпMwGTA�NW�)���:wA��;�2�ݘ 済r0;XFB��`��dd�Ҟ�\�yE}�NZf#�FG�w�F�u�"����8�^�D�T1ϴO����W�/m��Arlub���w�[�WonUޗ��Q)�+��	ՀV~?�Wۇ��Tn�pLw��/،��zxW�_o[���W��>�=rf�X��/iQ�~��j�A�ɔ�L��<��#m٬��1��u:�<3�>�cx_��<����U���3ɨ����,���/����p}�q%׊��S��Q����_�����-'\<��G��-��|Mj=�D�/��'w��M@Q��3���Z�.c̵�&�ײ��n���Xҳѷ�fX��1	��\�>V��=wi5{4$�K�e�*��̽����؎:�<K4���vq$M���{r�	�j)�Vx�F�P9�v�O3���2��L��q���޷L��*��:D�P��n�ư���/dz+'���Z��8���I�HIy8�3��\Ϭ����S�&��1��g�����iXme���s3z�\����;_q*@�y>�'��<5��z��ť��R��~����=q љ��Nm��3���(��;�EI��~WU��~U)���+�5:��@�{��w,d����9�.A�:�kn���R����2��>j%���>�n�g|΍�-��'Y{Q��NWt
���V��΢� �9;�J�<|a�*��Vr��ţ�5�6��]Ѩܛ=�Q�������W<�������g�ؽ�;��
0��􇤷���g�
�='��`lu`)`�K�s��z9$�wk��O���[�?E����v:��R��?wM
��񩙋��p>�1��x-�]љ���z�d�,�W��6{�c�1!K�������\�y�o�є�i����7e������î���	�X�ŝ;C�<�vō���Q����f�����=����K��4)>&��Z��j2:ߝ�f���=����tXI��^�Rqs�/c"�r	�l��3�8us�𫈍��֐.{ ����$Uƾ#��cY�cMXZ�C8fAJín<�-�X�ZN��2X�1zzicJ·��C\a/y��J�\[�������UyD��(���U;�|*�������9�n/w*=9WJN��돭��P�|���+2:��H�'�v�Np�����R�mm�.������K���Q��]���Uv�{����N��R�\*&A�jU�EGyE_kʜ� A�E�����Sq�E���ՃC��"jK�a����j_9gf�,�܅(%!�n^���v}��vr������\�u���.xW*���zYʙ��'N��$͈܈�.mΔ��ʃ�q�b��ބ�=��p�\}3a��A�C�K�ugzlb9�ֺ�;]Xf�������O^A�F����|�V+����g�RҢ{��5~[��-��?9����]C� ��{(D�1�ŭ�������Q�_e�*<�"�W�QfB$,��e���X�)�Gt���yji���>���5�'(V���P/$��l��»][�`ڂ��>�j�an�o���j�1�^m�*�gLa�0�+J�DP~{2 $��a��U���2y�]A1��3c3Ll���D�0G9���!!y3� Af�ɜU�����z���︖՗�j���Oe��MjrX۸�4� ֊�%a��=j�c$�yԁ�K�^����N�8xp�?]wZ�g����K�H"iԺ8u,���8�!���f������[9�stDoS�6�V��c��ܒ�r�3�fM��`���
���N���p�'�������̘��=6�����q=�u�_��MѺ=��������n�_�9��q��[X�{^#�L��Tb� x�95J{��M�̜�����<������6���t�o
�oa�>���{m%�:���ڋ�(��;�9�o�w"ך��S�5K�7'QU#F���_��Ʋt�������&��]�����⽕p��8�`g4�C�0��t��5�����f9�ͳ�틔W-s~���Iܼ��|WK�r��`u��*f�O������#3�#_�S��p��tRZ�+�~�,�e���+o}��W^�E�ᑺi�/}0˼l���s6�8(R>���r��lӏ5��ނ���>k��Nw�W��{���^�"��Uj�+*�`�L���uMܬ��!���������
�jgzue_��H�*'��������ֹ����ǅp��m`p��\h-��D�?f����j( ׫h��ˡ|���4$���JH��꼿,�s�8/GESy�17<4�7���9=�F�Q!�q����*d7Ymk?Y��hTέ�����֒�����@��~�;Y�(g����R�yKs{MMl+t�MU��p,i�ǧ2}��Zk8���`��Q��u9\�G��Ă��O����Ψ�,�W�y��:X�{��0o���q���W^}wve�Cw��ftr����DI[y���SxU�Z�N����`	ҹ�k�ͬu���N�Ի3�������&tF�fsl�������~�{��"�����8�����tE"zA=�bd�_J� )J^���;cnjt=//���=gg�0�`7�L���j����eX~�������0�c
��]�n��&����d��������Vi����W�M$4�"|�r��lO�=ao�v��z����N���k:�n�%�u!�����{v`f)܀sG���>����r�zq E���]���XUY͇�����B����@n���bsn�Ч��t�����9Zh��u}G}�Ν�����=�'f���7�[j���g���r �7 ���-bQ�)�&��*�W^^����^J��m��'��b�"�쳷:n-�c:��)��*���$:	l��p�xF�WJ>7�R���ｺ�Iw�S�t,�j�B��<�k�J�vD��V�o;.$�t<+D��Iz)�����.��������^Q�����gU�:���8N[��fjN���A�qxǐ�q�묻�{�{��+H`���u����}�16������f�ܭ��i�\1�Rs5T�y�W;r����T���y��m��O[����t]\��ns�z�8��W�&;��cw�y��k��w-��`Vy�Q�`�]�*&�퉭���|�(���ԭ����ٻ����W�i��6Js<'B�J�v{U�x�Qw^��uE�qp��n�Q����.h W��3���n�m���R��QQ·S�ƞ�e_�VU�]h'�d�Tp^/��py1�s{efád�16�E՚��
~��?^�Flk�V��{�(튓O#�'����&}�D�����%�ƪo�-�<�x?N�;�*�i!�nA���xL�;���
�q��X����Y�J�$*�"ÕY=�K=*�/�<zJ�^��M%.�!ڔ˄,ϡ/F��E��(��rD�e�ų�{*.,�F�{z�)ݲ�����,�Xu������d�l$mJ�J�4�n�fX�����U��O�s�U�m9�W�$��oږ狻��h��$ �$�SJ�3�9��I�yZ���b�����s#ƟM��mԳ���{fݻ>�U�� ���&qB�o2���X6���*�� >U�=���\2�zy�C�ʷ���(���kt[��fCt���.�]y�_7g4�-������p��1fV��� ��w���q�C�t_1�C��j�w�����[��T �� ,"/]_t����b;J^�D`Z���x#:������Ju����AK���.{��뻫z� k�r���VН�����t("!��K���Gӵ�����w��@x�nӛHj��I�9w��J|iǲkJ{2�$�yf���J�d6��ng��$u��s(�'��?�8dN�/
�e��橁��6����_�S5.�]գw�z�JD�^'��~T�O��^�����U+$]���,~~�J�x�~D����8��&Zq11#3"�d�9>e�=t'5dk��N���K�-�30�\�D@�z�)�ٮ��V���u�3c�����~K�{{V����إ���j�Mm�{o=n"��ݨ�����D�BSL��L�;՞�3K`<���)�*6_gZ������>��F�
����l�H%苮����B�g;н^Ov3|}�h�'>w��`���4���%w���W̽9IK���9�gh��ݱL�@�ś�i=peM���v�������g��yuG��A��.��?{\5�}:��lz%��rU�n]x�a��a����{ ��La�/K&:���Zwηj�)r��3���*f�u:�ʼMw��1wWc*4�b��oM:��K��6���v��-Z���ye�::�ᣵ�9e@}���p�����0����z���"�:f�Ӗyb��%��c������)#	v���9A�g�M�M8�	�TQ�a��n>�Da2�-��(up��l�+iJH�8���j��QFs
�\F�_�w���8���E�-p7�	�Ӥ�m��6#��mGw��B���ڢ�4�����kkf��Z�̼��޾t�hT����/w��5��bzüC%���������ut�nAC��Y];�>2;�خ�ji�qo��YƊ ��� C���Z��Y¦�\��o,����p9� i�Lb��s�p�4ε���;a�
��M��]��7r���.䐮�g�7|��'	����f+�e3;o�D�K(å)��er���Uep<{ֶ͇�Kqf��<�{�0R{���㽿9\ Q����k�#LEû����C������7�Vumpƃ�Ǳ.C��Dl�rg�w����ʙ�5�c⬾�J��k�`$�H��z;s,��^ݽAA��D[�f�Ǽ%	v$����AY��c�6�uw3�id7\GI�BPz���2QX:Y�{���Ry��x�a�!'p���-S��W��9�V�
�Cp}�m�sX��a�:�Մf��-n)́k;l�]��{|OM�9aN�n�Z��P`}2���;��ڬ�4k��y�jt�*�h�ش+)eVH�`�l��w)�c��+����A)��������N�ûQMe�O�B�Xo�2�Nk��TO/)���?E��V�#�#�%�7.lò��5f�4|N�>�S�}5��ނmbd��J�!��fBB�9B�p���e��kܝ,Z{�mӼH�*eõئ�F��_m��nk��p >Gf�����{����WWȡְ�/R��i�ս*M(c�Ճ������9�ե���J�l��o�mvs�Q�k��#QY�0���3�.���t�_�_r	��e#}���&�D�(��s�ۇ�S.É�sY]�R�jw��rn�eZx�HKfEr��$��m*:s-=��>�XT�6�!�0������#�,h�-���rg�E��O�3�۫8�.��eAt^z�y	0��X9��!��E��{�7n�g���b4i��ӈ�n �n���qTs7�:�2�ټÅ�"ʷ�T���o�;U)�L�q��d��(u�b*����i/�woN��.L�ۋX��,���J�`�j@;;yx��Q���P�z��tP�ࠍ�خڕ�u<3��d˜D}�v�R�
?=�kѣ�.�,��ڲa"�gn0�/^,����D��>Q$xB�wo[�{�)���bK{D���T�[o&�.�a��G�1�7-La���WC��[Vsq�3�3���{��#ވ[ں��8��-
v%"N-��Y:V�+�s�)R˧H`�}߾�ꪧ/�+�=��g��r^9b�,��2�TW�!�Kr5@V����BD��`���1]j�$�5j�嵲�q�=�s����v�KL���x���w���=	���%3�%s�9唆۞�!�k�}�==���Ee^u���9�a���	6#b;�>u��A�� �D�SԲ{vG�b��=���lO�)Mߎ�[
h1�A�]W�E���b9��*�2φFĕ�Ց�V����ن�3�ʂ�
"5foTF�;���C[F�9J��rڲK���6E<�H-#�$S������5��y�*F4�=��UW���'� �^���N�Qw��0�ڛ�0��{|�C��S�3{�^<U���y`��c��y���'-S�;WS���i��Ҳ�X�>9)��]װn���Piuc?�{�G-Ê�˥�)�׋�+�����g^�͹��Q�i�>w��>�ڬ�n��z�m��k�.���:i���g4dp�������I��=����@�ѽ���4 /�+���{ۖ�����1����T��懔~�Z����Nͅ�z+b���z����*�H{��t�:���SU5����qD��˃y���U��n��&R�L��H�{���#�y
*���6����m֌l������JyiR9�8�:�W9�`ݫ��:������}O9vu��;1i]e
9�8K\�f(����T)ǍU�X�
b{\��
b9o2i�}��n�6�p�Ǟ�L�}���HGZ�,�z�J�ɬ�+:�Vx�E@�<!�B��g��]�Z����b�m�'p��[��O��{�o�J�ඣ0=�-�y|��G��q��(������"3B��3��D:��#���d������V��v��^��p}�넽��tf9�^���zo%�p����d<����]ہ��G��o�?����'N�݋���Y`�T�K���Ӗy$���|�pDcUt��D��F��T��L�09��,�ʉ	��s�ߎ/`�x�>Y�D����KU�R�4<��Ov�~���v@ʿ_K���|p�^�X�֨�*s��{WM��.hwu�ə|���<�Q�`��+G�I� ���ޑH]a�����x���W�v��tN���S6��ku�����zؾ5���\���Ӯ-�����݀R�| �r�1��뫲S�!;�&*%du���aՏ+�N<��:2����y�l]
u�����[��;��e���M�lgusj��y%�����2we�k��y_r�/�}'�Hz˹?+�j�;u-���mj�>�շR�_+�7���8��v�kI|^a}����S7T�l�g@�#��C*"����G���9�Ta�ԑ�!��=z�#�\��'3����Nuw2<��ˀ�|Ļ�c� 칆4����%ۜ�~HY�{�B�/�+�ph�Ƚ�sܩ��h�yK��{����Yw�q8�n!���=����1CA:ϥo��ɽ���S�l��O��
П���a������oE�}㛯������i8��'Վ���>S�r�k�z�T���}OQ�F~��;�i���*LL�?�6o�����ա�z����{���כ��Y���n��=;].��A)
�nZ�Y���r6�$|��D�B���BW�c�\�?� OM@�J
��O2sr���Sӛ5�˞]��G���׋O�6� b^�j=�*E�
�k6��=X��=^�q�U&���lڍ�U{m�1�d��;��Y\�j!��F8딦x����+�9�x֋5�u���םAyP/5h���#�pϜ5Ke�â��p+vg��y�H�T9�zZʑ���(�|6ov<_���������k9�8��l�|:0X-�˥�h�g�V%x��ȇ��D~�^��5�,ve+"�w�D�'�=��V��ȕ ǣ�p���^��
��vX�b|��y<��յ�u�ܲ��G�@��5U%^���D�U�\���V`}����;��ܸm��&F��,���K
���8f���<�_)���v��Y��]}Hw%Z������`hԑw6r�)*̱�dV����kH����;U���H5!�w3k+��[��=�Qrq� �Խ��s�s�H�0��l�/K�~p���MM�k�����^7�o�s��n��{����H��ϊ�J�!Q֔�nԳ�mЪ�Fy{��QGgF�Ez�������!c�d�t�Sgګ �JY��cw���Jtq���]/W���N�����S"����Q ����w>όoD����������m�E>�����3��Tn�yj��^�Z2w8<���O�6��g��ye\�Q9S̈́u��Х���C�XA��hQA���94m�Y�����ʟ��ܵ�/.f�����G	�ܸ��o��� <�g{���Nm�ѫ_�D`�z(r�p�EˮW\K��9N�?E�8�|*�:Ӯ�S�H�2���:�S����Њ���J��0'qSaڪ�������=:�9uMuk�8c�T��ug��9{�gF�N=�f�3ae��q+���/�M�A�oTQP&8�̣��u�v�L�jjwڧUe�"��=e���a�*�mn�؊�����o��E��qm~)��W����OקݪClT�zإV��H��t+�;�AO�'^��N�,֭;����\�|\{���f՜�d�M�ga=u�u���{�m?J�ʴ"Qj����V{"g]���)�s�����syH�Z���Μ���=w�`�t2�g�&��:T͎��䋲��ׇ	��нA�U@��C?S��S������+��@����S�O?Ep����z�A�J.,Z�QsnjۿcB+��5�����Q���}	V�K�J����Y���#��h�k��_^���ˠ!�ţV8��	 Y��s��k�.�W#�HE˓�NÑ�ê2�Nis���g!^J?3C��lo��h�K_�7�¸*Ӡ�Kff5��cS<3�(��K-ɡ��j���,vs��S H�����G���<lF���f�n�-�k���F���t#�G�����?٢��p��2a��Y�HsF��ԍ�S��K�ݹeKΥD��G=�]Q�rz�)�%J^��Σ�N�ƻ�3H�~��R�Vf-=�#�
��V�]�Ijő�MU5�<%�_Wx*��</P�&y}�Z���\ӯi�W.Y��9�-:{;����ݷ�jƒ��:nE�ދ���#��Uq��E��>���̭ᐅ��v}@�ߓe��3���~�8�s�y�u���>��A�ؤǔ�~��<��G_0��jPd���kͧ���;j]�C%LAtz�4�=po�cznkǊ�q���`��w�rˮ��W+��;�K�3X�=;��]���d}��C}��`tyŋ�՛\sGa+u^�T��2Mc�=�F��]eǚ|D��i������mu���+q��+�:N�5	[�ٍ
��?FX�1����f�&=�0Qu�4)�X܌%�=qTM�2 N�o��jr�!�n��b�[��(�O�c��'픺�oaX0������)�g0��EA�
q�S�<zr2�G��d�_F��;to��������,��
T���o�S\�/>�"$��n+��@+�F����?�z+���n��6�F`|�{�y!dz�(I��#|�vye���퇻Y�(~qTSob�_�_���ɰb�����O^�o�,��l�Ȓ�Mtֻ��z(���k�a�x�yǱ�̻�w�ts8��F*���Z��z%C�h���f�OYw<��5��D7#=��#k�h^..2��md��c5���P�A�z�K��j�H��1N����)Xʈ�\p��=�sה!���^Z�'[ړ,^%:�&j�f���=*]	���nϦO���R�IL���G���݋��s��?{���f{�RQå��{Exp3$߻�e��1'ѝ�O�ŷl[7�m�Uԝ�ZlGM��T�vu;�(�ƃ�Y�j+OPE�e	K�{�3�H����J�4Rl�;L�A���u�����ut����ɖ �����sQ�}����;��O��߷���)c��'gic3��t�xc���S�Վ�x�k�W�&�^rt"�׽v��R	ėqCƥe����iJ���5ބ��c��b�o0ގcHW�2��P/�H��Ε9��U�nq��^�z�s�W=��JVnC�Xlg�3�t"`s����Y�<�	?�I^b�fߝZ�y������8h��~�����&30��3"vC0���LvUuhu.r�e��	·�^�����N �P[��Ѧi�6���&<Q���������/�r>�x©���Ɍ��n�3y�N��X�P+e\f�꽺���T鼾�?2�Z��������9��K��#�T�xgf��W�P��@5(v�N���z��ޚ�QsՈ��WLhaZxz�MC �ƚ`���"��g��q�υL�o��t�ԓ[�kF�p32����R�q1�����3��h�m�����^�[s��ue`B��c���Y���n�*W��Vy��V3^2u�N/�[A�2gU�6;ՠ*�x�'�+p���d��}QF�Y讘Q �g�ҵS�/�'M
��=@b�k����� n���1[�{)ٹ��j�$����V�f`��h=��8�:t�?GJ��e�Y�ɖ����s�����q6z�3Y�ڵeG�Ą�L�n��wV>�2������{��p|y5�"�������o�uf�6ﱷN�s%98-�e�giyx�(L>S��kcVQ��P���^/�Cfbb��p6��v�D����M�q��U�\uN��'��]١N�y^�������Eg5G��p��e�����t�=���N���WP �q울ޒg,�����6s֜sc6�X�m]Ϝ�����z�]�~)u o��f|;Ƣ5zP'<���ue�X͙��=������m�A����箲�MＥ�/�]Ý��HU@?,}�P�ʸ�,���44u�a�����J{F
@�4��7�F���c��Ǘ���흄c�}[���i�=�/3/T�$7r��&�m�"?D�L	�Uz�Bg!/7%O/�s ^������~y�@�^�SΣ.k;+�3[�����jS	���N���� o���rB�p+��%h�̦��L�Mo�ƻ��J�b����7Nkѫ`9�\�Vl�kff�+�U���e�2H�[��E�y�����W��z{���E%��׸�E�v��xull���ڌ>�{lAu�ߙ�JJ�/��#��y�Zsr��4/�zN��xz�~���䍹�z߹�W�q��C+����lA��r��y@��;���!�H���4x�A[Z.�U�Oת��V)�Wڷ����	[�����)�}��ݬ|Y��m��05�M���.mL����
�fa�{�y��2I�Lj���B�ōA�E�_kz7��BPE%V�e�Dʒ�H��[5w\j��j����=�nS�F=ZL`�ί��y�/x羲il������tH�IN�����W*7U�b�ӳ>ݓ�2{�|�R��a�>���[�
���2�:W������$LS-3����x���:���Mo�?1��˿b���6u�$.�|r�>�gR��H��s�����Mi	n�}��e��NQ�F��c6����s�gܦx�W[��|�Y�����poT{A���^$ߩ�y���)8��'ML=��L��w�и�3�b��Fu�-�uPyDd(UQ�)�֛�|�4t��ڀ��?m"8���Z�V�e�n�<|qS�Q��u�{�,>$�N�a��]���~�I�N�����w:��<�w��f,�S���D�%h�[�cV��R��V}�ؼ�D�b >�N���V'�P������VlQy׊h����enk�����=�:"_D�S�赗ǜ��&���5=p&���Ҏ���SLF���ҤΠ�t�׻Anv�8��x^��y����{��6���+G����<��A��^���zwV(ﾫ���s5�EU��� �,ŧ+�k����v.�ގBBt�n`��k|5{��ksrު9vx.�!�V��.
;��a�a{�#�^j�Wuc_k �6ҎD ��V��gf���R�n��0o3Q$���F޹�H���s]��C���J�_"3�b�'�9�o�U�qN"�{�Ta�a���N͸s|�2�V
Ʌf)d暡��e�&Y����r]�L}���htiգ�|G3���}_)[YOqT�����K�}��:�OZ�7"���@��P�T�J�E�vڝ���Ȁ���}�2�H�iV���]!���bݯs{�9E]{��g��cӼgl_��kv�cX<��k0!��ꎊ̄4�ȧ�Y؆�75a���;Z��1W��O�/n�L�H���}�O�V'=�bު�ۇ�6�VdU�C���W�dc���1_��i���z������v+�m{�OWq�LuO"��e�N�����w�q��F=�8�{aQ����S�Q�5W=[]!;2r�^�#�z7-)ɼ���`��ӑ���U`}Ss�/��=f=Iܟݛ�w�D)�{E	�]U'��)�8�
��`�J����w[5��G�ټ��/��}}�"�MX��(����f�8��I]��s�7�j�_w-�R҈�Ս�G��(2�������J��q��T��GyO']JyZ�s�+R����!����e�˼u��;p����/iGZ�ԛ=����뺋W ���}��p,���&P
_��E�����WU�ǜ_{�Ȑ�@����@�!$�$�rBIII	$	'��HO�HI I?�HI I<����b�O������Ҧ���o��%�@����j��pL��ӆ�?���
��)"��X�Y>e��R�Rj��ԭy�5���n|�E#K���;#�niP6!���>:�����$0}�Y�ԴK��t;��I��e�0�kkv�S̤�l���=%���(��؏f]ڏ`?^�B?w�����kY�Z���5�����=;'������{��As���Ǔ�0�UۈOM���*�kُU���C����#��eƬ���9	�s$��-��_.�?#����Jt-��S1�T�;��k��I�G�F�Q&k��J�L3Z�&�ܸ�)-�[{��[��^����׎`�/�fN��*��v�s
Ð���F�yJ�̹l�q�Ajrh��7�Kr�7�.f�Vr��X�Jo99r��{��88���'��*���D)��9;;��^ �QMJ2��l��,^�2�
���B^`˥��4��fACb��k��k$�2˥��5�A
ȅYT�p���t,����ude
Хc��hGq:�f���qc�)��"3�K(]\�Z�i�8��*±W�fYح� �C(Y�3Idk��t��x�3��V�9�W��)�L�qj�m��u	�413NK���Q�U��VV�y��A��K$>/,�^����w�t�`�+7*��R�6�V�܄nme���f�eP5V`@�(�L��ϲۂY�-^�Fݡ)��3v�$�`�ݒ��T��J�0���3Zɫ��I��{���QA�V�O[;[v�6.�d�.��f1�Pa���"6��c�wD��=YQ�姉̚���t���B9�O57Z!�Ѷ�'f��D��W��Ę��y�K3Ud�j�е�N�V�ϭUҼ?
d�ʦ�VA��
Y6� �-�&�81��i-�/2lF+na�1L6�^',;�M"�ٍ$sI�w�J�iec ݅}-s&*�X��|����ϵ�P�-�y�{�k��$$�HO���I����$	$`$�# !$I$�@!$a! ��� $FH �I?䐒@�bBII�		$	'�$$�$���@�HHI I?�!$�$�$�����HO�HI I?�!$�$��BII�!$�$���e5�r��pCd5� ?�r 	 r}�-�.�W #J"�EJ�*�C�,id�kZ��R!V��D�)��ڴb�b���V����NLĳ+X�4١T
@P�
)@@)�%U*)E�����Ҫ�D���@PQUT� �PAIR�J�EIRTR��    L2J)@� �w;�Q�w*�ݱ�������]�	�$ݻV�ݗ7C��u��Z��v�]����gU��g9z��4�����)<d�L�{s�� �`��lY�ݻ"����ٲ�ŭ�hۻ�����׍���ں��:ִN�pa˭lh�4v����J)P�*��$5��j.�{s�"�]�ڮ��٦����poء�mӆv(d��s���뵛z��x�K�]ݭ���b�1RR��t�i J��*U8�\A�9����Ӕwm�78i�W6a�p ;�����Ak��R��c-�k+3�m{kւ��ۭu{���S
�))(�����[<s��h�vm��t�S�{{;M������3Ѧ�vwtSs�ޝ���齷w$v��3t�`kJhR��H��@��\]]hj��Z�ᷬz�O1�w`���@�Dy�(ݑ�:� �B�A��kpٻ�f�= 9�@���-�����Ka�Ì���HbE&����J��{cs� �n��p.j0�p5��T���I�s.�wv�S�.k�48��Py��n�n�R����^�O^Ӻ�{��q�m�l�6�^�=v;�v�����v�8�PS����
�J�JUtB�x7�Q�s���R�f�Sa��Jo��-�s@����I;m�p�� a�J�J�"\SAp�9Af���T-r�!���9��P���*m�ۣ���w89J���M-����8��� ԥR � 6�%$�@ 4 &h"M�� z� T�U*  '� R�  � M$��##@����=)q]�5ı�5�'��zL��!!V������޳��H	$�����	$����I����K�Y $��t$�H$�������I}�Z�`�,���0x,�M���!޷H�)���{Y0�Fۦ�V�Q
ש,4�u��ʿ�1Z�-9Q��t�B�C.Q�Ӱv��ݭ�˼t1ٹb������X��T�@�+d:����NӬ(åޢ�ָMdn�F���b��f�;6��P{qE�x:i�H$ɧ��iZ���Iy�	a;���:�6�0*AHbCz��#�(��ƌAHq�&�b`x����@B��2��,����� ���d8�!ic$3�&�Q$�I��2H,f��x�]��+!ReI�$�x�� ��`�AM$6�:�+w��*B�Hu�ąHV��Y!Ԇ{Hz��Cԇ����񁴇R��z�ר]U�s�����m
Z��}iSL
2��)f��7�H�N���6Ú��^M	;VL{�hI�,��GELULy�T&�p���a�ku��(��+��GA�=�����אg���J�+j,	٣�T�mЄ���X�0el��0*y�)Vką�f�X �,!��Ia��CF��H�H-: �Z�yh���S�2��,�F���S5�*��+6ܩn����R�)�C�{�m�ܣ�RM�����Cw��U�1�1���:�H[å�޻�y�2���-��vj�
��!TfĤ�ش9K��6/`��CAI��X�Q]��wB")�*��&�JV$7o7���L��xP4�����I��U
ͬAS���1N⧣��A��H�1�Uͫ���� ��B����J���y�!�س�N�P�S(ૹu#�Í���'��Z�<)U��t/(����=`;���)F��4��s[4*1X���iA{ �/\f���W�R���M
v�C	F�@n�=�цThL�p0�f�6��y����1WA]�q5tV���7����N�6ih��V���Ӕ%]b� C[�V��ȣ�̬���dA#rS��UC6���䙦��C/i���i[��F��V����{S+��鉨�JVh!u�����0��hHF�V�V�ƽs"P̌@1&wq7�M�(�n����ֻp)PVl:E�y���6�ht���OD�-
.�ժ̐����A���X%n �Ɂ�^ӽ��F��3��s�6���@gD���"�V�i��F�����^�
+n��:�:R����Rn�L�L	���n~�cB��pV�`�%v�m]�Jf�2�H��ݛMV:(4���-صz���4�n���鸳c�65Û@���j��iѺ�&f�DD.�,�@m���ܻ��V�pa�m�(������ ���]�rf���k��-����m��N)^�nK���۸uC+�Zh8�[z��?� g6K��aĆ$��71f�E,���V�n�V*e뫢�����p�>�ދ��t22x��Yq箝6^9FΥ�cj�=�h2���n��*3��#v̋@՛�gpa�
`Ԃ-iESK
ӻ��P&�:n��aہ� !"�]b��.��iRR�o�R�s"�YF�KE
d��f^\
9����B5P1x�걢��]JtCڍ^��j9.����x��i[�NT�Ԕ)��m�3O(�{�V=�t]�*[���*�9�fB]�B������,�D6q�k)7wR��V����+DL�;�.�X�LҦ]J�w�<�ʧ�9U��i��iS��3vR
��^"��F�nS�q�����a���*r�N��;�:.��ͻ�Г~p{�`�ĔswO�؋�"M0��Y50FgL�#�Қ�g9��yw��l�-�!f6�׊^~E��
���6��ʘ�[*��(��^m���L�T��jV��J4Ru�b���jeкo2�97vP �I/5�����U�**H�ҠZ����T̎��)�5����I�F��AvZ��ye6	�W��B�F����T����O3e-���*���QV\�u�l�B)Qa���ה�Z;��@,Lb��k�VE�j!�n�H��E�y|�ݗ�k��z�4�<2+Zk̲�l��X��D~� ���ܚI�C�xoS�6t�<�ߊ�[��Qv���<����\�j"yJ"��E�C�L�w�X�@Z�?Z��:s41�cT%��� �V�8N%y��ym�wo���q�oi�F�ǚ�L
f�P��Zv�hY�mQ"L� V*�&��"���⥺X"�PmYX6��m�d`�s%�]Y�cW$:k�@C��@nG�i��H�{��j�ZU>^��oT�imdQ�5u��̦��p�����i&�k�F�Z�����l$�j�*Z�źJ��T4�[��,ا��(]P=�C�B�ۗnu�(U���n�x�no./��vww�7��R�L��(�89���h�h���1ՠ]Œ��t��֌m{7��܋����i�,�6MA��e�ګ���ݪ�*`[��hT�ɺV�+�v2^[��Yi�)��z��W�1�z�,�o�JGV�h�zh+���ٸ�m5)��j7h�A����^�Х�ɫ ��@䱴+fA6��\��P�*狂�a9�z020J��5ǡ����ݶr��Շi�ˉ;n�J��9�J���໠k�f�
��!�L��.�]LI���DnPeTf:ѧ,6Pd�P�0�N�&u�dDj���PiB�8�2�eVCoN`��Zt�Y��X�LU۩)�Sn����Ckb�_�[��;�U[ɓQ�B΋
�M'	JiV�!� �z*�Ц�%cCb�M{Wa�b�cÉ���ߔt՚SoɰV
Oc����`PGb��Oe�)�Ԗ�ˢ ^Z]����]�@������T9B��J�<���
Our�I
A	�MV��(�7Vwl�6�T�E�7P][���m�9x�fe$�Q���ZU��Ŋ�x�9�\L��?B���Zq��F�`�n/@h�R�a�C*�6*�<{�?G��ڂ���#�Orլ�u��6�:�~ܫ��wz�(�5)D��9�6��AF��n��(��@��ͻ�����CС�a:�~C6��B�/E&f7Kr�Vѫȳ1�.���j��ƳvA�[{�l6Ku������~	!��a��?��!B��ڶ����AaإdЍ7C3�"��ͻ�4hc��i�B�iU�X"0�H����)I�� Ua1��8/q\	
�J�b�;���PQ��1[X��F�[/S�`�EҦq�L5�!/v��Q���P��ۡ�#W�r#.&@�@�7$��4�r�����%�T���kJ�]M1
��8�9��{�-6��D�`��luf�,��m�,b8j�;OX�UEBލ�,%H��w���m�Y%Ѭah�T���C0��^�Oa��Vei;f5�lK��E��ЈAu��w{�w���)�R�i�j�V�Ul� 
�uy
W�2X��)��iӺ��+x��H���6���-M/}7%�72ӧ=:�:A޺nU�DS<�U�hKz�k���"(k[�������V�x����V���(��ihӴ[����*�ܡ�$�K�m�y?)v�V�)�&�ȥ��U�Ъ*� 㱂,U��n���5�g"�(X�EW���@��ȶ��n�ס���+:�`dX	�k��E���[ֵ�G6����j�#�~̊*Jq��Ce�v\�2����D
�JѬ�w�AAz����rhkHCk.�t�Z�@��Ym�&���FZ�� $��t�nఠ̘ƌۘ�Wy����[B��'s�"��b#n��b�"��b�n��@%�aܡ��j�iǊ��,��2e��Ni4��ʕ������մ�x�#6�4ʌޔ���ʆ�B)�h1&Zj��2�Y=�v���Ƈ{���:���r��EkY���/0�`R`�*�4��<R�4��L���p�������9Q\Ui�t�n�ƥ*ޛ�xpdE�Ziʔ�q6��������s��k}�x(��#�w~t�r�EZ���(��
���b��v���B�znU
�f)�{�3�8<�a�����K���r�2��o �N�P�VE��?��Q�_5�zʘR��2`�^Qؖ�b��V��P�A����4Q�-���赑��ͭ��V�W��A4�޶
�D&5�W�nwGb�VFu1R�6▍��Nխn�ŶD�]ݺ��&��@.���5!-��h�հ��E?�E�^�מkW���to7�k�<4�Z�1�iPWn�%Kn (�)Ձ$܍Q4j��sh���`��F���s%0*+��t(SHf��̥7
4*��)0�s��kn��T���kaWi���e��Pl�*��K�3�h�o�Z����=�f��x](�ڨ��T�ӄ��.�RoJ�k�9(�h�Y�j��#�&e
�0I3nf�1�*( �.�д�@U���5z�pVҔh��xsZʕ����A,��M3]���SEA��1��Я̢�kL����*h�Y���|�^]�5ti�$Y�(��K2�'M�M�X`";5�;ѯo��f��ovk�O7���'M^�ȣR��]�4��45�ٸ�"]2LTE1[X������v�v�5�
h���s}�E:�K�V�<ݩ��Mﻛ��P2��D�#%[(Vդ�J$%�gl�U%AT*�z�J�4̪փ����u�CpV߉�vV�"t]m�5v�˧"��(Խ�mІ��n�y��&Z�s^nً#��Z31Ʋ�t���uVn��wN(�Q���5������Qv�]���ʦ-K�*��	1*��B�(X��2��t�in��I�i�(�n����a��A�
T�]0L�K��]��[�@"�\�.�$ШA1Z��@_�vo�p5P�`*�N��O��2=���7-�:����0$�Ov�.�i'n�9p�	��֧153Aa�n�T��y��DUE�TQv�X(��Eݢ�4�Qb�εS;�
)�AE�(8�Qb�=eEcƂ��m]�k��kx?ER\�N�@G����z�6��#MI
����Ъ�Kw��lMFQ�Z�J9�<�v�V�
(�S�`j��40�Ҳ�P�CH`9�T^�@�ǌ�����7Ge��k��Ҵ���V`��8��3`�a35��S�����7��R�鸶��^_:�]�������DN%ט`��DL)���7��F��s5�@� �e,��e�7w����j�y�]�U��C�p�y��8 ���tb��v�T0|<��D@a����M֝�ۺC6�U:�e$�z�ս{6mL�7V'�G�G�q�t󗼻T]3̢�z�w,]�m�a�<͚�<ٮs6��5��kB)k���h�x�uy�7�SH�(��DN2��3K��71��p�ֵ{����w3����2x0���
C�NJЎ�Ksͫ$B엖�Uk����-�{g+���n��3�3���W;���3SV�T6[����yw�����Z���;�<�q�ؕ�M�j�V�_�ۀX�:Z*�\9��n��5/J��3Dr�t�y/o;��w7���`�	�Q�L�gf��9�WX]�/�Uw�[�Wx�8l=H]T�.�R�~a�cY1]!�c��˙��Mc���Di��㫬9��QRЃ��Q��"��n$*����!i��i(0����Wv��ƞj �EN;,fG�T��B�(�I�NaƋ�]�iC4��cQC�e/�YvwR�^�jP�M�����xZw<�|lc�wo��S{6��u�yin��̽CJ��b�)2�J��E5˩E�d#�꘢e��OR6�t��P�E�Un]�`T��&�$�k]�{z��3"Y��fk5��)�ie�or�``�e[`���lغ��<g������f�5.8���U&����T`�'�RC�����q�Y���a�'QV���E�Dkn�k�;�O/(�\ÇNqz�o��6t��n�e���o�;�!ER�Q����ڄ�D�[�J�'z5ſ�%AՉ� �P�k��Q������`��4S�4�U��ýG�ŀ�DA�I�-�+�UJـU��P��e1���I���#�BP%���U��f
��B�,����E�b���+�CMlh`�]2^١J���zk2[�vȠҩP�w�-ѬU5AEo2��S7Q� �{Z6eФ���E!U���L
-�w'B�f�����2�N��׈�tq[�ٗN#Y�j8�K���!��7���3u*�j7��)���L�;A0�V�+%�*�Yh�T��6�,z�ܩ�2a
�e���0�^�:�bV=U�yuOP��d���
T����rVӗm�2�D�P9���x��Y�B��2�%:�W�IA<�0!���L��[D�KjJV�����̡N����:]����%�]Xa� 	8����32^�<V��7�Dw��F�II#}$o������G�H�I�#}$o����7�F�H�I#�$o������7�H�I�#}$o����>�F�H�I�#}$�����7�F�II#}$o��F�O��I=϶>	�����8��u�s�s�PH�7���je��{$��D�̇g-�yֲx���F%#!2��a0���[���y�I'�,���E�-�gqa6����;1s�Q$�mr\�7��$���INCgvd�k�^�D�Kt��Sw���{x�Z��Id��$wzbY�u�'z��|t	�����Z��K��+����A[	$�+�}$��LK���m���.�%�
g6Ȅv�|�s��:K�$�����K�s�.���lL����T)X��&���o�R���<̕zbF���\�E�]��fV�HȦVqۂNp��Y&s&r�{�$�y1�����OI���GwYh��w���#m�vxn�Vf�sn�gi� R  �%Z��ٺ��"b�$�-޴�i����Wf��gPr�{X����L�$��$o������[��h�m>H����%����z�n�4��n���2Ӂf��HCt�gm�L��R$K4Y8�u���L�m$u|���lB́|7��#�NE��oz��-F Ԧ����6ۧ5؂��v*乧�������^>�]&但)7�p5���W3��#Q��K�I𛗍���˼�'ȤE�´���rU-�zQ�ȭaY\�KF$,[sz��d��7F��j����ˎ�6K�eB���[&��<��7�xi��5y�v��S�Oo�v��|{�摇���]��qkr��q���U��R���v7Y���obI,������;n�n�x��f%��^>ڶ7���ݏ��oe�9��xι��`J���r]t�t��I��ǁ0�g[ײ��=n���g�sUƞ	��Wi9�%���(
x�a�`��.9vzS��u�0�]3u�;0���p�;��k����N����w�e�9�a��Ѻ2!#rm�r�=��u\s��|,�lV�k9����k�;�Q�Ր�Lۻ[�+@�%�7Y�c�jo�YEGw 6uι�{|e��Whu�K^uJ�C�P�	�n4:��7MZ8 #������ҨN*y�ގՔ���/^\����#�:��4V�Od�5�B�	EVR��͘��ɶ�X8ڙ�n��;[ȵs�#z��[��w\��5��$\�=ͷ �r�nW^pə�ir�X@����T�D��s�R���"\��Ό�Ʋ�2��\m���7$��wn���N�8Zd���ݮ���FOv��Ŝ� �9.�1�a��,���Y��'H��ks8<;i�D��:�ۦ�ǯ �_N�}��H9##��]��Җ�Z�z�8P&�ݮF�'C�l**����ڵ��� J<y2w�"�E���	̛'_I�u��
�uCԓ��v����7s6��J�KNI;��E���������y�MR-�����̏�N�{�Co>�L���+;K��Qub�Z(�;�䜣��%˸��_���F#��|#h���H�]7$��t�F��Ϫk;��&�bĖ�%�I(�훻��w>���M��x��D�.d�L��wW�q�����'�;��5�ّ$�y��w�Ӽb=qy��ěl<^�#}\�.Gb�J�qW~�'�g��ƹuhო�ɻ 1�`y3��:~]�G�e�9�V�rĵ&:��TAb�fJvXʗ33���%�`G�"�oݷ����o�G��S%�ޫF2a�����$٫!�I�ѭATr��s��شd�%`���'<K�f��v�&�";���|��4�&T��7:�]�dv��΢�5��̒�!D"�wIuڙ�uv�,wp�oK�V�W�,W)K��֚��7�w��m�<�-E���5vdf���B�ٵmDؗQ�=�ٓ�(��4:`S���f<"�C���,�]�VWnǝ�JAnk�������QԘ�J�P0s|�Ҵ�!��5�I:
E��/66�gT��j��r޻�CP4����D6�2�g�r�>����(d���v���{�4*���ji3�6��+�0�_]��qk���(>n��1��r�����'\Pòl�E���^[�d�v���:�l+���=
o'Ԥ��D-�7����9'��1t����y�p����o��Ś�zJ=5�����Du���f��ڛ�#S��ޖۂ%�A��:��3��cX4�٫�y���D���BںX��C�����Ev�,Ǜi�ţ�W��d:39��F�)I����V+�g(:��hp��g���J|m`��Х��k�7�^�C-��H �8�\�`�&mn�A%&��+&ΐJ�'WM��N���(H����d���m����H��������eQќ	1��p_=Mk.�[�z�/@�����K:�]xǢw��:�՝[+�f�NE}�
ﶻ>#U�|�3�8����*��]m���y�rÍm>�{��De3�c�r�)�/8�m��x�)��M\W��-�Q�+����̺{]G�	�9;e�l�qÚ�Z�ɉ�u��h��c6.�Zj7,��B#��j�ŝ�\�v�839&�x��;*�6�ݸbJn���w���C|�wZ��4���(�쾤���ݓ{�`�oZ��u�P�s:I]Kj�X�*��"L�mu7�:^V�K��ʜ��:`��׫�:*I	y�B4��=�D�ãe���9o�1��d �2��E��L[��n�cX^v�#h���Q���,bT]��Lx��)�n���Y�u��j�:3�j��eb�N�;8N� $�,�-B�V�`��p���^$;����(V	��ܻ2��/%9���oP��7Ab�;�M��޶�e<Ɖ�v �r#�\+3�j��Y]�Xئr�ٽx���(��S|2���m0ӗ��5d��k�+\��x�%#�6�$���d�Rpv`�:��2���&��v�Խ�D`:#}܌�/�ݾE
v�E��\���n"���ƭ�b�e�������=v(,Q�C�MD�'��N�
>{Q��GJH64y���;܊t
�"�s��8't�,t+/0_-b�ќy��(z�۫k5
	SS����:6��wE��&y���L��eH��#]�6l��	
̝ɷ��v�u�#��ħo��Y���z8cБ��6�w|�I�r�.2�ݸ��5.��.Hƺu��x�����+�T^�'��u����Z(��X�k9P����Εd��
c��ko����ƍ�	��u<�gr��oR�tX�oevbq��.8bf[�R^u�U�^S���k�ŏ��z⨒�Wj��Xz��u�l��#��ib��s[�n�Co
H��q+�3N)ʍ�a��R�BV�\���3GN-K��,�{�K�3{�%c��C�35:���Zlުb��Or��\��e2�F�Z]7�yXt�{����;��k^��8^����C�s� �E�pT_V\��!,�헎Q����$mo<�yhIu1HJT�,���&S82�j�ۜ0#�j�֯�uN��z�̼��P�0,ބ�*�^������Rw��e��kH�u��v�lCI��\�\�Ժ���ۋ�m�L][�� �  �����r�B�Q]d��tx�ri��(��g�$ʾ���5!r0��N�=�
�F��Gf^�c�/�J)w�d��CC6�� ���L9��vz�w�|���:eJ(������x�Y�2�}S3)�Z{��F��}��MΧ�@}�wtq�S���-��M�|����2�+���e�+U�r�x�\��,����}�y5�`֥g4��P2�]˗7�vH�`KY2�w:�gqd�sm��Գ;'5�&N�̋`��\/(���j�T�d��X维OI�O�O&���g+|m��.in�Q���wnӍ\J���d��}�v�g�h�:���c��7�Ai*�Eq����Y��YV�p�/�
�{o+�SU��v_^���5.�+-���н'$��nqMZ���>Hx�b�Ɓ��A^��c8�	|Z15�7&\afc�Vb��VE՚wZ80��V3�����⫭�VPe
�O% $�ffV�St��]��������sr��8F�`^�Y�
�1I�4`��[A�[}������Zٍ����׹:����uW�2�Q���X�m��f;yb�V!.4ok���)J%�xi@'q�4��{���<bܫ|��M�c�2�Be���k��IݨTP�@����Qm�ڧ�*��j�^][yJ��s!�
��@�����Oh�S���F�ޮ��;:�F`��+,���I�[՞�E��"��v�bx)���|t���!<��h=��T���#\�8�fڊY<�ٹܹ�5g��6,m�E�f�+�*�y��:	��r:4��*�\�+C՛Q�����P;wO^P���a���{�R�)��gP�;E�NۤZ�/sD�E`�o���A<=]�17hk��P'HWv���ru����#bd�̤XJ������}���������Q;m�&m���6�{#�[z�wI}�^������Z3{�s��$�i�r�RhD���Z�ɔRO^C:��X�3*����漠��2��\k%�{�d�֫r��j%�(H��W��6�@V`[���Ewc»ٛJT�8Z{�P��ڼ@JM�h!¤��`���/PMV�(G�k��׈u2냸�\�
ɽ�)૭����fe�\�}Hv-J��ۜ�=�{W1�H젦Ժkt����ܣw�W�Wu���n�B����Wu�¢�p%��pa���SM�;ܦ���U�1W���o�����h.6:\v呖�<��ȭ����_���j��uDM���x���3�*6��i�T���,����/��y��{xeHm]�jOeMX;�5�֕����9��$�
���#�\V�N�ם+��%*��cݾ�Ť�;3���q�xL*�I�fU�=� ��'j� �n��ˠ���S6���kX�Ν}6'�q|��h�%��W�]\���u�]�ux������P��ڻ���{��f[װ`��f�δ�D.����Z]Ӫ�=�'Hj��(;�xp��I.��pc���{q3V%��z�*�%�+��9J��G)�
�A\t�u3������Iw|.u.�]�����ն_�3EhNH����*�0���%Jp恝����'I��Ѣ�:,�3�7���,��u�U�»�6�V5�z��(S��s���e�S[�yWr���\ܴP�%�=݃��r��!��ҫ�v�Dw'j�U����%��Y�G�e�yZI���L���W�	t�fk�%>���.^P�én.�:��On��Vf��_Pyp9�4����Y����P�7w=�oyPshfV-�����6�f���	�KC�b��we�h(ƫ�y{�]���b�j�ݞz���"�u���
kk,r�4�k����n���̛u.��z!%a���(������\�E�{��5��@;��.R��P7[Fu�b�q�:�U:���L�YXD��r�2k�Zki_�Sm�ѹo�����V�ٮSt�xD�UX��c1˥}�^�N#}W�����1Y{�ԁ`��Y�Cyv��39s�(F�������\p����v�S$ݢ�F����8rz6�^޻kK���YNlm椻���Љ<�c���!��Pҳ�w:Y�� �=O�U�)�.�g�9��n��:��֩h�@V��.M��%ѺKGH�0]S4�[�M��K,�6�>����:�Xj��lЛоwӒU�����TAu�ˆb])�WS./zx��EV������x*͵/vF��ވ�QK�p�cY�����P<4�sYNy��X��^a���Z��\��pL��2$L1+�����=�pVbCs���ͧ��>�E[�,��/5I�Z��k��n�_�x���%��g\�x0�	�������7��<&Ս;�5Q���7�p���FTwK~9��E-��\�2
ZgT޽ֿ4t�hg-�x������l��V%��s�ٕ}����ܾ�[�`d%oDjDi�f�ƻ���J �0���T�/���L����"��豨El"���N}ƹ�;׼��;V�J�n�TS
i�tn�d�P��1�a:�����3{5����Z5IP���v�э��=��`|��o�f�c
śщ)IcL�iQ�c�6��&� Vh׻�dH�3%d�3����q�����*� 
3����Q\)����o��)kN��̙��{�8��¹��3Ӝ�i�$u��h��Kr�*��]Xl9y�s�\­鯳��h��˰,*�Z؇Q��,��WA��4R���>*��w���=4�:؆�x���E1Om�lot�H���VC3E�ְq�����������o`嵜f�a�󛂕b��yy0ika.��T��%��e$��B�v���"�V�M�eڙs.v�-u�A'i��
��}�a�v¬�r�F�B����p�ZE��(g��Qn�j�λ�nGۃ�󭳆� ���7Ӝ훙ϡ�m�{r�δC�|9���U����ĵռ`}JcdP��)�C�A�1���yMV�C�*˶Յ���V;�ޒY���N_��]͗t4Y��6�.6=M�
��梭
��&���P+M�jV�J����4g[Fݺ��h�Ku�j�a_�s����Z��,�N\������׿�J�WY�qkX�XU5^�sp��>�o�#0�<�1#6.:Um�aaG����5���;�I��>]oE�8�m]�!I"[E��zė�HF�b�M��S����s�/n^kǥ��s*\g<Ɖn���A_�d�.7�k)\أKul���Ve��A���v�<�Ԇ��3rW#2c�ְ����ZS�[���Fp�x�Ƃa�TR�љ��T`��cաL�@��:���+�ƫ������(Z6�u�_h�+4��gU�}MQ�q"�]�':��֙}g��p����+
me�Mm��s{S���;�;�EO|��u����	$��	$�?�;��{��Mo܀C- �aB@IH�	�Y *BE� �m�	X ~��I/�������+B��5���	BZY��%��l��HP	+� LHr�	�I	1�$2I ���B@�a ��CL�.� bB@�Iq!m$ 6���HBC�$�Ћ ��$$�@��!'SH�@%$/mIO�$�5�B9@L���{��I��N1@����!*`@4���/�$XR@��l 6��`� uHM��	1�B�I+$H<�C�$�Bi*I+	
�'-�1!)�I�,	�BcV�	��*��0B`T	�Bh{|�B� ��
��[�B2J�yB�RB��i�\� �$3Ɓ�,�g���\�HL�`N$&�	�$%B���v�z�֩!�I��wVI����K�2A�0��%�A@��\���Y �!$1!��0��j��^jYd/��&����*l��!��1�3�"IĆ�&0R[@0�d�Om�@Y+"��q�&2B���LIi�Xt�H!ĕ���a�d6ZAa���!X@�G(I�I�H��W2O%`u��݁���8�MR��$|��I<l6�:�2�#i
�d�;�@:�ld�@�X�湐<a��H[���P�tl@1�L�[@�l��yhM\���l6�P���CyAI�M��i��%I��.e�L2���q�;� �d�	=�d=��*Hm&Ѕ��Hse�MRJ2!=f�\�i�=C9�GVT�sM��;����1f1g䚠("I�TP��x?KV�
�˴���6`����[�y0I�X\R����=��~dVۙ����r�N'�$ ��O��B� 	�{����{��w���{�y�	zogqj6��m�؇ƞC�&�ow:��Ô�C��j�6�����ٹ�ّQ��X�엻M�*x���Yb��D-|��&�v��+��;���ջBe���9�֘�Vf��6�Ǚjv1�}�yL&�2���`v�J�,\�[�B�ݍԵ!�����eѹ�.p�ΚL��s3[���T�+|��>�&tj���&���5R�-@�
�Y��u#E,�[���+�\�ͤ]Ζ��[�&i��T�{f�<*u�CS�ě�س���.�m�y]0]v7��ҙ��d�ԥ��]v���������YC:��Z��y�b��`�Q�fܡՋjvQg�^`��*�S_�X�ʔb&�u͍�̾�[��}[Ǩ*�|{����\��JʺsU��!�@Vs��2���c� 9��I儇ʻ��t��iU�*>hmI���;M;�vdV�Ҝ^�Z�ҫ���S��E�� �
M'�wm>#si�/W��o%���+v��ٱ�pLKqĸ�.�W꼖�^k��[:T��v$��Y��y����.��Eg�ͧ����B���
)�3��hҒ�+2�Y�K��Om���� ���9�gFw7_T%�6�����W�e�f��r�.�n;i�r�wm�F���ˈ�v��|D��j���on]��Rȸ�J�p�vvƻ�i��
�N�co!�!�����u��	����sw�9�?HHBOa������<��˗����*9}]b���]X�[�ܞ�cU��}�l�T�ZRh�5�<L5֔x��4����i�_<�4;���~�[��vl5ȳ2?�Wh��lTS,c}���*�X��k'l����3��W���[�m5>~�u�yxq��9g#a��O/G:�7o �
j%KHY�3O{�ܮ�P�&��x���Uz�Xj!��^{�_Q��B	��C�kE� %ww
��W��U0V��4��e����kz�%�v�ZZ�u	mT���n����)��C��;�*��pг�񇓫�o�}l��z�/6���bP����4��������A\�ޖyG��m���W꫷Ag�G-RufKI1Vv�p=j�E����43��5��k�Y@L��2�\nc��
H
,"�"bJ9��׷;���o���I���rM�{s�a5���7i�)7�
��|\���R<6w`�~ ��e��\X̷�)MP]s�fw>�C�(�i��bm���L��=k�U��Ix�}z;�p粯""�S\l�N�WO��9�́�'�ު��ʎ�4p���UU{��S{�lW�oRR��8�d̺ޙ����ra����r�����}C�o�9Og|�o�J$�5��rޱH�uܔ55A����*�V� Ї_�P��&�s��W�Z�WV}�"�VE�}6��u�-^VrQ=��ۗR��y�gII�i�޺D����L���[�͊a�9��m,��k��n#*�QԶZ<����S|T���*��hĪ�wd�ʨ��yb���;%��z�^�==�u|��0�]]^G;ס�m�G���̶��f�iY�d�2:a&�	�!��5�I
�H�-�/�ز��+�Za���g&��4�Y۳�EpU'�c���j��B���cU˦�InH�/&m�5��rN:� �2^%�M/��}6N_.���!{������J�u9Ƥ�v��k���b�vY��EtM.����@)}k��Մ�k�nK�Beu%|\y����
�{�~ |>ۗ�nw�s�E柊���'�cd^�C�_�s���sF��y���g�k��|�ߟBHh$������<C�	W3?kH���MIue'�����y�]%/���]����0r�F0>)�6{1"����4vז��g%^Qu �����fh�r����=U�+��y}}u"���O�F�U��R��E�.
�֗i�{��g%)��h�fuS+��� �s�|D@�j�Yy�o��G��;�{��<�9��o�h;�FVn5-�f0�|�n:;�l��:��8� q��<Qu����glv�=��F�}�Uz��^�T_P����ouv�>�o�=["��h���+�#gm@���f9�J�4��@�<�	'���|ឞgu�jާ9�޻�y�5-Z���tVV��N���@#c��%,�k�i�6�,A������3�e��UW���ί��t%ݷt��XUmV����s�����o+o�M��#i��>���Y���|\���H:���ѓg]��7܍�Ny���y��k��D�|w�=<ےD�d�Ϟ��4y�S6s��z�[�J[8詐�\��+���R�t���Ǯ���}�=���9�	
Hu�> :����>'F�*����.Q�-�߽�{�O����hM0`,����3a!�,}Xք���5"�}Y��
�F�J��W������K�K͢5z�qR��k���wZ�����[M-��7MT�,ۤ/��)�[���-�o����M���F
G�yV6M���VL"��&}��M��%񕙫�Z��mvP�9 sΎ� ���� �l�����u�^�g;�f;���Iijۋ��m�W���}U�M�{K��]��)ۆ�Ug����J}��塞�u�rJ�t�)/�(|roJ�ݾ�r5U��o���ޫ�.�m��z�D�I{Xz�Gz�e�j9tR�[���g
��[g�[��D!�i/�?HI�B��~f}��Yu�/ש|���W�K�c}O9�\�g��N�P��,�	�_I`�L5��f�{�z���{���ޝ1�p{c?�H����`䨪)���X���U*�TB�,JE��H��V���[m����'s?P}�[��S��b�t��cU��Yԏ1�r���7f-q�w�;��,]{J���]z[��V����rM��d�Q�ѫڲ��\H�1�U��u�,k�k'*��P^t��ހ�T��L~� t�f���M	�=�}��b���2������_�����e7Ώ-����l�y��j|[�#U���{��|�!��k���ka�oZ�����ȺO����3����vn�H��_>���c���ͨ�����}��U��<�ޥ�f;�f-ݞٕ�w
�'N��sWl�|,��f�۾t��}���ܬ3p$׾��s�&���+f�'0,�Z6��۵"�ʃ���+�/��"D���k�h�N��/w��=�x�_@���}<�5����|������w�;;��w�53k�߿>��y�}��>������4FK6 (���Z�݌ˬ����y]���1���S�I�p|������y�h��arp�&җ��a&.��]�;����[t�n�ݧT�7�i��'(X���?|�	��B��͗����)��k7���-Ì��EwVh~��Ϗ����n�=;O��{���!��'��6m�$S�J�%�Bz���=]�\(Z�]#gu�a<�D,#��_��k|G� ~���]�����{χ޺���m8��K ՁVKWlWZ/1��ΌR�H������ww*��^�� 
�w%Z�BOp��+�����^u����k<�oS�_�қ��nw���#M�ô�{kx-� ��]��6b)`o{�A��˯�lđ�)���wa�hP����P�Y�3���7.$d���
`��v�W�$6���.^H7r�y��~����s���!=.�r`ۇMbƚ�Ʉd�!R%��}�DS~��Y�Ir��z������Gl�}5bV��vJؔ�����W7��A��:����SE�.����y,թ
�O�wrL��q�ٮ�/"��@1ʹ�s/7��c�ު�7�w�{�ޯUP�����G���̎˵�lC:e�� �u�I�y��_%6�I���U�ꇻ� ([ }��'�WE�H���,�R}������]9c%j��f������o��z]j������w�����IC�lH�w�ܕT!����6ź	�T����{;C���e:�m
��������hj��	W��;>�{��7��sbx6�}P�.��p����4�#s"Q](�.��`�ե^�z���ʶ�c`���㉀ > a�{T�0�*�oGJvv�m�������oc�NDNU�;SU�{۰o�#�}���7<����ؐ?vᙓ-�!P��	QF�+i*��-�ڧp�y���U�7;s{��Z��hJ�qp\���]�yٴw��On�
!\wx,A�gG.�z8��rle
�/r,����\
�=�����9�������v.c:2�*���{:�s�����3�UP3��q�#�ڂ>��$�u��oB��̟�R̨Q��NJ��3��{��(��$�d �<���}�S�����!2�{2�Vq]�ݪs��m�YՌB��`7O���5;=��W���o~[�};��O<O����R⻯�f�[�2�0Ǝ���u��Q��"$�����y�zX��v4u�vL������X�ثi;��зu����r����\k�-S���F  ��v�0|9�l>ۙ9;��mT��Y�o(�����X�r�s}�?f~�B�K��DS.y�牧_��ӟmm�܁t���P�	�K]�����Uk��/�qĲ��T��Aq^�Y�x�b�6�����e��K��N盗���˜�p�ːt��N{�{��~I��w:?!!&y�w~�{0	���$�=�o)X���ݮ7�t���D��h\P�Շ{Y�{�{��|�p[�v�n��T�mt���J�tS��nW�t���/��B��[/q�NS,|/7+f���Xկ�Cӥ쬺�t�&�L�L}�:��3�u�rT3�z�p�A�2#�r��oh�2�>��UC�O��<��o臨>qï��Õ�fy��
y9M�c���Gz����HF�ܽ;�:eǏ��_y��^�׹�}	$���������{�꼯��wd�i:�1����q�뻎��l��9ԌH��r8"�}ذ�eM� >�=��;���q� `�8��JnQ�ULJ�9��5<I�(XVaT�����.
�(�Q*���zA��U��q�p>ɕz4P���n�`'�w�"r�ȵ���[|���Dzޙ�*_9sV��#�,�l`��o~�����7���y��n�9mԡ�û�m+���V����o�w!�ܩW�֩����r�T!�\�����=�:5���N_}�Jo
f;F���D�G���1G��Xb��L���Օ��8�#��V�l����m�Ey�|�|k۹X��*u����w�T.Ҟ8��m��r1��o}��uC'�݉����4���y�~��	^Xp
�%�,~�,���Qt�*1Tb��+��y�q�,�a�m�鵃s�t����0�#�cnkY���Z�t�{.�kՆ����Y���*#$�J�R��D�4�
��eT|n����2�EOJ�m8�H�fq�F�`b&����Di]8�n\T��L��6�}Ɖ1n:	�S
�2�ʫu��{��Z�(���9��'vj���7NP���.k�wte�\���`��)�E+�(6)F����Y�6�i��O7�L��}5��W3�7��@1	:�J�T��$H�� ��d�,��2�*B���#���7��͋��}���Z[�`o
ZV��0�Jw/�\��_<(tl��G4d�V��y���m�kw[ݖ��X5R���P��r�J*<��6��>6t���k2��[w��KUo�P?O���wI#m�����N���Г�K/z]���I'�%�))M��w���&v�=�$O.e��(m����D&��,n�y�im��/Xb�m�A�iz'dM�Êwn��p�A�K[�:3w4L��s�5���}�h7��`�x�m"�]R��z�N��<�5�-����4�7�F��k{5Vm��;��� �S������0�V��x�e6�=y3����4�.�^���r��3о��N�����D\(.���R����ݣ8�"cS;WG�^�؜���.�2'�׌��3��=݈�'�
_@�F��٧/\�yu�L%������­s��/]dՍ�ǐ�w�����]��'�Gq��a��x���+�<c �^�n�͕�$V���X��;f7|�W=�0��jÎ�Y��N����wz빌Y�ث���M"��ؠ�GN5���r�jں��[��h귶��i�8��4Uփ4�ۓ�U��JF_%���כ�^��#+���'.:���]�]���ptCV,ݤ̶QAC=]��.u	���V��;:���|�y���*���͊�p��� �bs��b������ �֠�ww<��N�����C.��+�]+�ڊ�*ã��bN��^t��t�f�n�th�7��w&�Lbm9��Ƥ��r^�.���h�V���z�7���x�ꜟ�u�-}�Vi-eE۷]���� {��Y��q�.Z�uuU��X�R�r�5C��0�/kq�����ơmt�ͭ����5��̼s
���C7�-�чDe��5�g\��z��.�J]�����d� >�t�[�O6�)���/8���������%�	ԟ�Eό�ߜ~AY���l��Q���?�z�Hw�W�Ʌ�=;����>����!ttL-8�@��׌��m�reL���ׄ}5���iv)�W�:�l��\�줰���>q�7W߰�ߎ�$`��@����@DE�$X���1�,QdY@@>�����Ow����lbƎ��-�T�.�q��
�k�<~϶�	|��"�m#V�J�Òw���T��Ё�����}_r����-]��-�����^Rw�X�r#rb���X�v�L�i���_|���O��
Ͼ��`�uU��4�-ms-�݃.>��{������_;���짯�u��A��ԕ�f�9�nw����)0���n�YB`˘��ϋ��'�b����{?'�$/��Te� LE�E�P�[��Pؗ�Q�)�voM�/e4z��9���0c�rm݄���ԗ�1��[��$Z�}�t�S!߾�a��5�2�xw�	 ����|��x��X���'n]N'�R���M�������u��C��&8]iN� �u���FLA����j4�7�`��v���!|��C�<��U관m���ֲ��xު1�϶�p��e���BE7�U��D=sd�����G�^Ǒ#� ���Y�p�I���[�e���1n�o�i׈��d2M�W������㵼������7q�1ڋF������	&2a�Jz~D8�Y�;]p���F��鍐���ʥ�p|:::<����t��Ğ⎊s����Z��l��%fF���> 
�8�d?H�\Ml,�Vv��#�L�S�#v�pZ��޵�#hy�߷n}�{�0�0���YY�OY>B��+!�T�@+�ǩ$�!�����f����q�q�>���a�ĕ�!4���4� <�S�N�PҰ��'YS(:��'���,�8���?����T:S���f�E�0e"���d�,�!e��l�z�}�31��g6F�6�0�����_�o��Ku�F�$)�|�@��xh���v�@�a�?:b\�wUڝǩ%F`9��C��?���{.�.���w>a8�� q��@P�d�'��=�<IP�O|��!��Y���H6C�p1*E��<�C�~�������߷u��$X>Ri�Bm�	�z���:��R_i>d�{ߴi6�qY%�?	?3�? �\ec��̰��ԟ&{�������7�o�+�c�$�w�����}��$;�$�'ټ���?%������=d�8�O����&��@�J�	�M�_����7f8fhJ��V��$^vL����5�Ӝ������^o*F�Nep�*M��ީ��|>�.P�D��dņ��O��OE�?��k󥪷H��5=/�QQ:wra�	�aN��f�R���\����=æ�j��|��׏��h>��B ��kU)�Q~�>�I��+W{�mI׶�;LZ��W[��W������KCY63ͧ��:��܊6%T]�UI	�pY�w5��}�￹�\��z�箿k�֔�%=��֕�1^�t�W�Uw�{�������"�oWS[+Rxr;Ɔ��3�z���P}�>E�B�����ٯLRf��Q�Z�D~IS�w��z�ψڗj��]M�6�c��	ZȺ�5���^��\~��cJ��uˠ��LӔX7f�Nh�Y��9mh;�o�����TK�O-偨�@�F�ߏ���y�i[���ew:y|��;���g}�l���x���y�/���'��s�`���lJ��4�0�	Ee[9�td^=Ѹ��s��1��������]i�p�C�Ǉ�����泯�q*���TW�� s����=	
8´o^�ps��@��wD5o��,�'FS�Pr����0�4(#�i|�Z���}���׬޼3�����#�\�Q�!Q�c7��̴�M+#yד-^+�U�s�1O�B��:�T.�٪	�C}8e���o��>����	�3�+�}���\-4*���;*�8lG�J�Ŝ%�LF����`x=��}������'���7yr����lO7�!7���.�4m��yT���{�WD5�ʪA��=��p0���g�g��3�}�k~���]����ߗ�<��g5��X��4�*����y�|�׳���o7�[}�}κ#*�_,�4�9�"������#9�Ž+bk`�;�[�9��v5����{M&Ԓ��_e�c���}�,���kK��^���s<��{�s�6�WU���S�s����/�/�m�.��ֺmO���3yu>�d�=����E�I��Hw��0ƻ��3>r�+1 _���'KF_hEF�{����[ߧD��>����G8����]��f����������h�H}���eN��|*y�>knV$�b�-jVFO����|%�ї��x�ń6�+xW��뼚'jj5����W�����ė|O�(��ջ5~J�Zz$MC�������Z�8��f&��3M�}�vV�ƴ�Zm���'"�@���A�{���r緳<�T|���������'�_��"���h�Y�L|*����N�����Kp�:�O���P~^�3�gs�2��^�fo���Z5�nE�]��j�owS�PX,��TX"@X,""����^f������;o|�|C3�oA>ݽ��O8���F>?h�G3.a��YtLiRU`AAQ`M2IH�1��HőA
���c1��)�2L�����E���B��V�J�BV��E`�ˇ��4H����v\��s�7Pl�Qu�uz�{՞�y�B���G��+̤U~����~�9x�^*������@}�PoT]����Bd�{�O}��=����~z����t7��2�=���qd����A�86�rY�;c�F1��]�&��`����\�m>7�_�~$ ���5���y��ԅUVu��y�;�:6x�7���x��L��_A�ݑ��#�V%�e��;gsϾ��{Ϲ�X]'O.n��k__��y�~!�C��J���N	���~���hA��y|w#�\ʑ6K��F���+Tm�9�K��Z6�������wj^�R|��5q���  +�^�G5Z�*j'�ozT�L���e]����-Q1`#�n|x�Hp�>�Qj'�4D�������px��1�mGQ�|> a����:�/�o�#hjg��6/���XE��>T�K욗}V��l��9D�����,��D�-�/�����}=������C�A#D%B�*6~��5�;F��t��\b��ZF'b�&����:.��꭮y۴=4�}K�_g��^+�IL0݌��m�od�\+k��v���n���_�V�U�B~vs��ܐ3���	j�cISs^�$jgy����}�n�W㦲���ߪ��	<�;���m	��n\� �doi��mi�Xt"�Rt��Tx*�5�V}�c��Ĳ����뾶����y7w�v�%�w�%��C)_�Y��(z
�1�ze3c��H �%��o��l�� ���ȧ�D���ZOq��g�8L�	4,�Y�Tf��Lny�C��|>����|E�6�T��t��x��ɨ`�"T��uJ�/��U<4	hۈ݊@��>��`nr���W9���o�3��z�����w���T>��ao�5V댷�ꬸ��Nݧ��cS�
������k���ܹ� ����$�|S;S9_]�`��u�����> t���.���~����Թ�F�,s��I����~�1b�^4(�hn������rw��󇉨�ᕷ�B���+�^E�������-eKLǻvO 5���oV��t��uԛ��üN��jNЯ���R�֣�:XU��phga�]�[�75��S��}�+ۧ^���O/�n�yϳZK ����TP;��鴰Y�oweW�;O��������w	ϲO�*���{��cC�g�ґ����_{���2z�;mr����������ֳ�o����f*�32m�_��g�~���A�����rS�¦ZNb�	���0gv(�������d���~^~ϻ�/�y�u����$�?H)~���G�W
<��&*��Q�7!�u]n�z�S+޴nb}�@ָ�./{�A��Ԉ5����|b3��[�V������k�!���g�GkZY=}��.�`T�ί�j}��ص����]��;)}�F
Xc5�~�D�F�7V|}��}�?8�[�2`��+�<h�
�J�Li�]�˗�c��� ��Oy����,�F������Գ�j7���޽ָ��mDU�H(�Bή���*��s^�}�8E
=��p�úߴ9�m���Q
:��мT�O=7���t���Z�dx0���G"W8�&i׻��`���/��..ɦ0�(pk�(vo��M��SЮ�N'J&H0|tm�`��黠G�$9Z��W�X'��E� �9�nی٤+n�;)-����|�i����z6"z66P��	_,����1�}�/ō)Z7�~���|`�����G���{��eW�B7���g�Lzc�c]�Q��;��R�^lO!�oÕ��\O�#@g�]}�G1�)�-{���a���N [����Q('"~t���[u�~ok��r�3�I�B{�g �!�'��~��3�׸�Æ���7��y�k��TD��?�9�m�#O��������Gt��� yҡ�&GS�g"�A���p�GE�Q]� ��R&�i�����7��	�K,
z��X�,(u����ȥ����_O|0����=�7�c�h��d������R�I��ɇ��Xc��P��~����w���x�O�0�>��Q��(,�u�p<�]P�Y4�!�>��B�6sZg��)}��P�1���g~)�]�7�2�%*b��d������Q\��e�bj�[�e���JSVPL!b�B��Yi�p�+��@Ę�b�Ȱ��1#kHB�,FS)VQ@�]� �c&d�dPa�����Q��
P�H,-l@CB��}��ߍ�]2A��\��Sz�%�v��ARCP�4#��������Fu5]���]&:w[4�wsLAV��`&n�m���z�b���|6Jܝ�٬��D���K�?S���������O}"�!8��v�b��0�(�BL�PG�wT"h�����"��*t�>����8���3��(g����L-�U]��1�?�)�]YEW+��A�7����&q.����J�z2t�wq`��7H��twZ��{�����6�ٖ��5��\���qMD{�����s��a����TU$=�Y>��B��Q5���^��S��
��iN�����q��3̸��f�����������p�������R|��@�On�z�E���MdHZS�{����N(�7@{�W�R�C�s-iqY��З�jq�? �B�< {x�> |"�y_�)������P�DsH�ŭ�J4���_���z�lVCf��}�_o�X�"ϑ�i��L6����V���K����o���7�UX���{��h �W#�5@^��k/Ү��ǁ��B>���S�����{5�[_}L��o�4pC�S�墴���)u�d��;�~w]J�\tJ�rq��=Ȉz8���ve7���B-Kz���V,m SdS]��I���cr��}�/�+j�$!�@l(�N�h�����<t�l0�Z�5�"��aN���h�d�ȝ�gwl��]�<T}fVB�Q�+�ؠ�c�j���C]q|�0�P���6�1��F\ͩ�ϕ��N��Ѱ��6{����rv�$+9J�u)�TI&;�X+���h����j�^��.d�SZv�U�AS�V�$q&$��,e:]Ԉ0���e˽�������Wo�l9�JŚJ�y�/De����7�N������͛G�Xs)K���w�������6z�wtks�锈�<�|����hT�LV�M��{)���3�j�nR!lWe�R�ytRB� #)�kgM����Ɏw����`�f`�)�RC��`�fS�R��)�(��u�y�|��gxkfs�x���<���y�<q��NF�[�0�v�!���r�ڪ�ëw��"��\��}��F{M��.^�\��3֜z�Q�b��I�(@ޟ5癜%�l�zx�t��������Fc{ӹ�f�����@��M �˷���ގ��-�[�5w8O-�U�@�!Q�-K�Z�C���{ +�ׇͳx��R�]�FºV�u��~��d�}o�$��$x����P�ۏ��u��'7�����;�+H�%-<�5��C��X�e�2tjZTlY�|������o-ɴ�������<�t��V��Q��^띣k��$�%e���u�e�\ֶ#������ժ��7��-���>�}�ܯ��'x�b8����o��v
p���h'�tڈ���=T��+cTTݼJ1K݀[�.�SV��SU��տ�$@���-�F���YR��Q�g;��6My��-�?lޮ�M/D�*��E2�sB�X �v���3���|ș�g�g���K�s����wc�ηd��Kri��M�Q��jII]�����^�ܖ|fq��Oe��v�4;2�n̹����qd��>{IÜ��;�Z�ׯr����Z��y����+eK���Y�?a��1|#�	a>�&��>�#2�r��@۷�wv���rח݂��j��`$�G{���ԁ�T��J����^R@X��!��yΏ�Q'?&�WF�e�?��}�p�`�i�rG�!��ҙy��#y���A��65b-	�|Nf�ͫ�S���]��Q�Z蠤Db��A�������y��x2�D�sziB�T�j�6^�-�^���ߨs�՚8�q��7yfJ�4�j=�Zъ�5w�q��)�㊸7�!���+�u+0�U�̀걯�M��"*GCX��̊U1����W�U�j|�e����᪾=��C�!M����+�q��2�wq���sw���0s��}a�y�I�K���^ip�����Y��=�J�vMAZk:��Up*���y�{�ٖ��$�_�1y����y#����QӡK�4��8h��*C����Y��I.'��^���ԫeV��褆,�4Dw�|#�i�`��0^��%��l*�a�)%7N�������[�z1DV!ć{oS>�{�ڙ������b�/��
�kםfD�z���z�$�*KD@;1�D�WK����n%�������P<zf�Ap�Q>U��5�e�B�
�s�p�$���>���+��w�f���XM�!z�|ȥ��=1�1�:���Bu�{�\*���n��ʊ����>�mF�,AJ�.l��Ĥ�C�1��C^!'Њj��\��X�l�`��q�u�Bvj}�Y_]�k��]��������0����b.I4jõ{�G��*'��¢1�.o���e6UP�y��V�P�y1��6\T�h{$G��ǬC�MV�495�DO��yN�Ȥ(�i#�M3�g��9�2�������wy�e��5[�{�z6Ҡ��9�(���n{�ѭM����Ac���U`�j��*TR�,1�J:-TQ��F[bQ�X�ĺ5�ȌU�1Iq�s��A������v�]����۶�u�'u�E��]l���5�tVM)���|6�ZX����AnW5]Zt�d�3	��(��6u'웡�[Z�/~���Ƚn� �B����y=}/0q0���J�#(�e͈��|�z��NY�n �WĲ�[��l��㨉��;�%O�h�}�#x��}^�����-Q�;�G�v�w1QC[|T��B�b��6������=q�����|�.}���F�o����߻3irD�^V�W��ZZ=d�G�7���=��{p�Y�c�`oF�*���ޯ��[�3����fZ@��_��u�e[c3o��e�ۙ�Fw����V;><[
��`�7H����īM��e�?H�Q��V�o9�,3{a�0�OJ����-A�QOw�QԄ
��-"+������)�X�X��)"K���S�*jq�;�P�.�gW�E�C�Ŷ�fz	!�|���W&v���O'�xכT&Ε�iL��|ᅢ*L���S"Z�Rgz�V�E�uU�ﾍ�,���g�"�/�)��g=v���V=����
/`J	T%B4�%z�!z	4W*Ue�oS�X�躼�ֿy�_=>�ku�
*&X��TEX�����Ծ��VU�|u⸒�|���*���|f�]Y[fF.=n�����d2:�z��r�VR�l�yBH��9�F^,�����Ҽ�{ީ��ޢc�쎉�
��
t�D
d�Dԅ�"=&n5�dpx�^�p�.D/ ��>�#���O}����-%^���)uoo~�G��v�C\��~���1y�H{��k�b�H��-.H3e<�-�ģ @�,�s\�Ҝ�ˉ4#�6	}�Mr٤񵊉�)�p$���$s�a>��� j^��uRwyG��m��G���V����V�1U���dp�&V0F����obm//��*#L�V'���O�Y��'�K��IG>})���n/2<�3_�#}�!/�a_�a�~{�gnD5�����&.���	oul��rѢ3��`ah�-$PGː��A��9Y�g�!��hCGEN|�kC7�g)\ߙ�w�	�������f�����%<�R\����0�"���=G]5ϫn.�L�#�긫{ɢPA<4�ϓ`z�/�i�m��g�kV�y�W>3{BI��3���9��;;���?BMg��e������G�9�}Ѳ�(�NR:�%<����$)�]��{��8�-�.�F9L�-��!(� �)���èVJ 2��X��:�C�z6M�,��i���O�*�n�5��:�9=L���]\%�4Nh���F��;G�ʻU�~4�י�u������^��~���.���-	�s�i�����3^�W���ć�#L�֛��?�m�M~��ӵ]�]�Gb�RMv��˻������Ϩ�a��ځ{����d8�lX}���ٵ,�Lz\�i������[kwXb�3��K:�����ύQp�n\�һ�����{�8����OZ-�ꁫ��>�Ԅ��| O�%�b�{��b��cwP\nB��kN&�榠F�9:�(�70}�}�Q�F�Ť����V�J���:X7�����CgwǺ�k�ߛi���O{��]	����%��o������;���Mg]�<� ��60�i��Kǲ>�aF��ρ��e���z�p��9�����9�v��Fک�G}��ަ)v�W��,z��{���L��b�}�vۙY3�R���(}�Z�Ũ������
�R�3�q����Z��!PA!F-Ea�dZ�
��Z-YQ-e-R1JD�e����*°(�T���A(�E!B��`\��������G{!�-a�Ͳ�\�E�dĻM�ܾ�Ki>/�5�8f]4n�*��UŘ�V���i���h<[-���p� V\̎(��M��3��I��I����q��@�Z�+DE)���[���	��m�7q"�7�t��mH�V����ڮ�d[���ňi�X>k�(l��f:iok� �5�7'�VE�*N��cz#��{�͈����/���u�o�y�O���jB�X+�/�|�D���J���VE�[�����6�cg�I��r8�K�4��^����`���d�S���(�%����|r��٨�/iq���u�r��T���Fw���_��zzЕ�z��\m!�0}��_F�Son/`]�N!��ӯ��Ll}�`�~F�إ���U�c� �1;�7J�x�� ��D�����I&��.���ɦ��~>��������;������~q��>�w*��M�Ud�l�8�`�x���8� ����▗12uʏ$7�g�޿���R��Q�b&.D�7���d&���LK�ɿo<t_f�N��fb�maQ��W95�<9;�׆#��4�"$��ۍ+w��
]�.%:V&����-(��W�K��׌+�j���|طb��e�E�na/�>�0/��.�S
���F%�������@�U/V��+}ĠL{�8\d�w��t����iO��wl��)����({Z�*<�\�y�ٟrf����d;��ҳ\${�'2 �C�������˯L��|~X�F)������KG
�=��rq(�z�Y�=r$��V�8�LF7��N`�ջw�E���rPJĲ�[Af������u���$�~�{�u�����}����:ȳy�&������z,u&hf��%w����^�53�C���r1flL.���GqY.7"	��� �
�ʲ�G�M ��&���&=�TvN?R��鲐�k����u4\+a�H[;c	4y/��~s/�����m��V}c�#F�����}��yp����C�Ar�Ŏ�WQb��� "LFV"��K�=�����p�_}ߞ���#�zE8Ԓ���JC�\���T �*�ۧ�XNX���2ĭ��N���wu��7-�֐\��]���e��ξ��]�/FuP�o�]Ӽ�����<��c��y.�vP�X}�8�� ��������O�
E��Y(�@�AQa8��Q�0���3��o^����.�t�X�_�Y�ڝH˓R�k�=�^�٫[���<3;��H�B|W�|������q7�c:��t�b��q�3���$1�_�K�QZ�+�uy�*^���l�0V�%�'�[ZD��"�mR<��x�Ǹ��|�%c��Pso�l�d���p�e���x�b�/i��Up��V��[����7/ތ�|��{�+�l�ꏦ����}� �R�ۿ5��?_;�3�h�G�㺘�<q�`�O�agl��*�*������,�ZiO-w�C�9���=���y���}ϯ^�z�k���?��A�z��w��i����-4�A���.��o#E�}\M3��u�:�)\82���b�x :����P!B�pI��~�����<��K���{L���%�K�@�<u��V��w��k�z�\}�Ƃ�B�q�x�A(�bG�3Ьu�/�e��˳W1�T���D�!
-�������L��Ҧ�E�_�\B�W��1	��Pr&{W��{O�^�]&6�����|�{�0����,��mْG�s��4ջV��@�t�j�=��D��(���l�/��D�b�wD����'%AN7*޴�����7�y���浘���sG���!�n�nk$lSXw:�8��c�,�jŌ7+���`������g }��E�d���������hlm�@lπ/D�CԴݯ3����U��q��z���S^ӽ��V�w.���ܡ�Z�|�|����@�L����Ӟ�Lylߢx�/6�|>	?�����aѪ嶾�]���g�⮮$*�N[�a�@�'��?D�k�^�ϰ_��u�����	!5�N`��D�G�I�!bz�:*��Ig�K�_m������p�v�3z�x;�Rd��ə�F��0U%<�Qf� �?V`�q\����h�>�]L���vһe�<����+���kv>5�{��da{'�7����sF�]ѿz����N�4 [ۺ�	YC��}��ǣǶ�6�*&9�����Z�'��[�鷞���kC/̎��U�z���
�5�k�ٿ��;��߷���k��@�@���~�u�����[p�8��G�H؄�/۝�G�>��t��G�K0��*�������&�r��FS!��W�YF:�����RB,������������=������w�2��&_n`k��u�J��*W�:��'oA��{����6s�}������W���ɿm��t1�vE��lC�TkV� ָ�QU��c����`�h��\ᄄ�,�s�^ܿ�o7��*{�C4k˫�h������ǿ}+5+IZ{.+&�0���^��Y�'�[�|i_�H��*����ͽ�;�y;��+�W��j
�V�χ�(�c-���I��0'=|/�b��� ȅh�70�E2�@�X�UZZ�,j�J�l��c%��FX���bJDF#X>A@
�f:F�k�Q�@�d��,��dܫ�y�j��f�Rs�uJ��J38m_WFUK�3�R��1��]Eb�ùs��]�C1��Hg�=y��ڤ��Y�Ix����|4��XʤXݪ�/��b�-��!t�f�R1��~$$��$����o'���Y鍌�}3�������^u\ݕ~͞󵥋��4��J�吴@X4����؜�J��UO@���ܮo��ݭ���|χm�{`����xt.kB-!�Q����wN�g�j�#lm�Ɵp��3tk����\�fK��(������^|>~Kg7��xjjN:=$�2v��/L8�^3d��f�f��+Uw�L�x��[=U�9=�צ5��v >|=���|j��'��w HP���x����WUD�w�l��z��|(���o}I��QSGG8�,6��&]�Ƕ�UAbM�{�Y �	 �I}P��H�ON�н�3�(dt�z��@u§��F����O/��!�䣮��`7=#Z;�q%�n�ݳ��w�L��*��� ��,O�v�׫�n���+;��PR^7��[��J�4�U�g�����fm�;.ufڧV�gh��:u���u�{K(6݊'�#��Q���<2����95��8%:���o8���{�y�]����+�;��il�#$bPSkF��j?^�c3LZ�%u�S7V�MASvl�r�;���ȪIvDu�T��;*Tׂ�򮳤ft�sb�0D!���,�\���˭��������ۛf#�:�Dt���D��5N*�i��X.��!a�K�bYa2��R�v�*�2����AM�W]ތMn�=�j�]f���,�?�*"��� 
�R�mcb��*�X�s�,9JY3(RH�i�k.�<yxk'Z��<�|�d��KsV��� �i�� ��M�'}�s�t��n�sY��3�X��ְSۆ�w�u��k�j�Ȳ�ӋԮ��ce,�6�Yi���=B��;��(���6J�[��p�6w��B�9yM�\�S������@��y2��bi��4,�Tmw����������&�C:�� ��#��^���-E���H�}$84Âw"�<����J�z��4������MΕ$|�jp5,+ݖ�^�m���'^��}9Y���Ed���X	�pũ�gٱ{u���c@fGC��F��������I�N�l���v��pT�nAi(,� ���c�*�]Ô��8�yݮo���WP��חϊODѦ��[M�b��&!��
��sVWg>���I�t�W����d�ŀ���YbXX��M�J��.���!�"����v+�i�<�c�I�y�8R�Z�%�1���)b�/AAֶ�׆=;�����Eyے��}��:d����j$�Ӄ�{�]��aª�\�#���K�rlb(��[款���
����InS���G*�F�3dxU��C2��a�6�&��3�=sOdQ�{�H���)�0?j�h;ZzWnto[l������
�6�%��� GSS���i����F��ׯi �mJ�J`wFu����&���)���hs �p&��r�a��� �j.�����AF��&�\���h�f�"��n����
���Y}��Me�C;/�S���m0�L@n^4w��K��'N����#N���A[],+zP� ïK�{\#���2��K��@�i�m���Pг������+�Y�c�s��;x�� �us�ĝ�������UU���Y��M:�}l��E�N:�o���W+w.^*��$�}�K��x����/-�s���G�:m7y4�7C�,Z����]|$�q�m\p�뚕�+{`x��#��"U��-9�l����^�L��:���ZV�έ1۲��DE��8F�����#$D�,3�@���߷�֮��/��6AYbT臫ٱ�N}hs��G� Zy'��>��d���΍[��:���}��w5�ˣ>�^Qy n��}�+p����x�W<Q�ѻs#�C��-z���7o�������D����xy)I��8G�ᘐ�j#�b����ә���8+}M/���E��Kg��#��k�<텑U����E�܇jw<g��]
H��)����{��L^F��^�Q�� fNw�)��q�,��0b����S�W1�'oR�8�8�dћ!٘f���p�>R`���]�e����i�7_߽UVj��������I[ޙ7�}�=!��r���<�_o_��{�`"F�����ƴSVFerz�yq��>{�[���+�<��j�^���Hkk�sfL����S��:�WB��e��Z;����G Y[�O=2���BH�W)�Q!�[SS�{��o|����1���5�}u�����,��ɻ�]FM�~��4����x�O"�:�'5f}Y�=uɍ�|^�4���Mn���"�+��߀��UJN8P���/�}<JV��Ѳ��O"� 1e&)�%2��q�`�m��E�|>�|�#O��=�����뫙ߛ���u$0$��tGw�o,>��Y���������˪�{n�z%~����$ýsTG�>��yG�B�|!|�mE�'j#�2{��D��N;�ܤ��ɲ�P�du�W_�=u(�C�̩ˉ|Dt�֎�Z�R�nc��y+��t�t-�3�����2>��~���d{Q�8�"�fB�m8@�db�����{�0D���V�vs)%gֱ�а#Sz9��EB,~�:6�����>�m���|>��Q	a�! -r�w�߿w������<����`X\��s����S�Mr6�w!��}�VT�Y؍@ئ�{h���N̚	���ȕ}@��:��Pe4�.y�p��4e�l�r4������2E�r�ǩ�� �qٹ�L���_�&�P�d�] ���� d���*���w�_%Ͼ7:cC����)w:	�B�쇩���EG�L�ծY�����w�>����Pv��^ �>$}~��P�tL(��INw�v�M�;�e�=�;��-���ą�R3��Q|��$c�mf�˅�}ίv�N���G��^B����xH>���_���ܩ�%���s��ftQ�蚮sp��>���$4úfK:�ax�C�`�I���sZ����w��#��{o���f���X�o��v��)g��?���V_������nˉ懼�"��z?s������@�P�����s&��F�'~�[�?qs/��(.��o���#8�E�1/Z�v�
~#~��C�|����0R,t��K��Z�Zs.A	� �"!��-3	1P�h�r��׹�c�>||��=�e���3\"�����D���q�Cx���tmѱ����_d�9��Vi
*�QJsr�E��LN]1��ǐ"ds�t�H#�ޟP�����ɟ\Ϛ[����D�Q~�a�����\����]s��b�����֙��<�װ����ۉc��u9�z�`��D�I�̥������U$"�E�uϩ�ɺ��H��ձ�jkݲ�������V���r0����7bpJ�~��K�X�.��"�`��^�M8=�8�Qִ�i}�<\j��(u�XF.f�Y�P�C��r��D� ��e��n�a��)�g�AcYc�j-�����J?�t���s���2�k^��B�\x}q;��m���Ǎ�����׷�s�6z�� �1��`A@�) ��/ߏ3�=��^}���-�%�Q����ⱻ�ƍ���%��Á��q�|V󇷲�<�B9d .���u�ˊ��M�M�Pa�����z�덧���;���.��#��w��3�ܺrjf�5�2Y#��)�I���1QfR�02��	��.Z��f�G�oey�T�6�ɯH�� t���ʵ�-G�&�Z��a��s����uг��u��E�ED{s1�M9,��q��)����{{�,�cd�Y���� _��<z::��Q���ΜEu-4�߾ ?|2�c:�F˕n=��z͑�V�\��\�T������0�5��__O|��M
�MR��z`��W��;يFl�'rQyok�����4#��\#�v:����������o{����ђ���9�Gw��F�AUF��<�G��$�q�>\�4�M�{lE1�>D�҇+1���*�rz�#���YL�:���4��K;�2�4�����1s�'�|V K��o��-
����oƢ}���`Ͳ�ݾ�NG��9g]S�Ob��N�U!��=o(�KN����b	��>m��	=�Č���{���2����y��y}]�?e
z+�R?�Y|^���1��=��	�P\s�wk�C��qW�,��ꐒ{�BR��w�a�^8�`(���H�a*EH
�"$��~w^������{��|��9X���o{��n5�Pq8oNάM�ޣ�Z��.���:��V�k�F�븕�zDK��L�L����_K�N%�������!���'gFG�U�R�_)ܕ7`V���CZY{�SR&�A��5Z��Ӑ�zj�G���W��a�AT�TO��������5ڙ	Sy�D����	Od�Wt���0:S��7UU��s=Lcg��y�]��y*;���>��z��q��	��!���9�y�cr�m�f�<xRd��(B���p��J�:*Dm<��y�2�����/.�K��$bI`E�g��񨘓�GE�@���%b$I>{.�j��1��w�i�~��|{Z���^ �c�S�]Z��\�%�����	�ۄ���6���0	��]�>�R}޹IY��S�ޜHx�����Dk����#s�9�$;��~�urz}��K}�/�2��,���.�"�t���U�By��.��Q�DhՍ�5�kx����4��g�%����3-~��=J���i����C�G�M��Ь��"�\3��%��T��N���ܮ��94��& ������
Z��g�71̟�t�Ml�VG3� 1w����~�Ů[�a߇�Ruʙ����?�:{X��D/^:���I>��H�����0k�R�S�F��`�>5������%[���"���^t��E��&�q�3E�,�g���Ҝ񤾢�����v�j������s��k8!+�ȟ��~�}U��h�F�uv����xj�;ο� �DV$�J�0��/33����O���A�����z!߾�S���e������T��2�h�0�3���a��J�R��,U����~�$Eh��"1z��,ۆ�"�.TVz�i| ��\3`�~��;����U���s��t��W�C�D�f����#�)�Z̖\�k��-��zܩ�\�(_d��Ͼ�΃���=Y+gG�Dp���D���`e��r�QV{�5�t��u]��W�5����գP��ú���)GY}ut&�E�[�C�!��.�i�2u?�ӈg,����vk�<0�Ãf\�ӟ�w��j��4�_rb\+��^�+O����	�O�p�;�N_Di��sꔞ"~{Aj&�A�6:k�=֡BɎR��H�J�!�w��6�������M��Ȫ+ ��@YO9}�����?�w9����k���f%��&I��l?(�����bҘQ�����Ξ�nf[S�J�^k�`�m!���|�2��kW��~��{$	1��z�^����r�{�'��nL��R:������9),�6ƾ�	��&�yyo�E���ƙ�8�5,v�Np5�7��B�N>��߳={��S�\�}�H{翿~�m�[g�1���NN�n�����|��u�^�T�)r���
r>%��:y�s��:p��xD !�z���}j�Yl����J�����<�1� �Wdz�72E;����w��&���^w�5�4>ʖ�)��)J+"e�r�b���b%�b���B�PA'��ony��ׅ���<�^�[�x��#��ئzc�n�Ŋo
v�(��Ϯ�dWJ�f�6�tC���^
g^,���Q�G����&���#�>���w���4̩��l�i� c��RkU_}r�'�����Ô*��+"�U�6�	_r�coF�j�:"c���9�$}������baNg�u�
pPg��U*�/�o�wI�e�R�ӝ��Lƹ�׃�X��"�{�O�L5�`��S^�@/+����Z��5�Yk�&�C�|�+��L�tT��vu��Oz������x�i����_n&{{{������߿]�!ns����;dǋ>�\v8Ҿ��N�PcUGP�-:&������g�q��u�=�.
��+�mg >�n�amnZ�{h^��9h��_EQ�ĝ�Q��F��bC��<j*�'}��7}Cc#;�!�,�l�lqKk@�q��ɉ�=��@���#b�i?b ��r*#k"���J־'��L�V:�_�;�2�"l�C�2�\��&!1 VE�,��w|��ksͻ�x{˫�ܺԺ$�[Z��gGM���N���s�^�n���ˠ�\�U:�g�5eN8%���Q���Ӷc8��⎧����9	GT6q�,܎��D��q󫶟��������7~�o�պ������~��|*9%��¦�8�]�ir��~/+�c�O�Y~u+�M��7�ong������=���}-�<�~'�n��>�s�I�"/�|��ѝ������İ���Eo�-����7���L��'���Dwv�&�_(<�y����ọ�8:	 =��?nי~���S�R=�8!+�{�����9S�Y�����gl�BN�í���j
ZiעrZ�GT�)�����d�㣯 ��a�������Kc�����Ϛ_��_s�jLj�\z��H�Vqj��)Y�f7��wϻ��H]�߾o������}�w���_q��~�΍<FR��N�~=񙏚_�����_v+�wXL�_P"59[ |�|>����	)�~���LW�7���(mm���݂q2;u���j��MBU�:+ w����6���� ��3Y���j �r��$r���4خ��ol�u�l�]�̾���M���o��i�*��������V(�{�u��8yyw��VIM�ś^�5�E9ٶ����V��C����Q�e.ٯ����EqY�e]	G�9��eu �hj�5��^���4�T&/f�p
�ߪ� W,�����G���55�ʧ���i���Vy�.i��뎬�s1{e���-�-�/;��c;��w��i����Wy��5N���#AG�b
0�1�kMw4�,��F�!J���@�5X 
���KC �Zy���k�2�o��[�7�C�m����A�l�wj��c� h8�]_�^�9=Ub�|��0�MR�Ւ{��ӦU}�H������ӛ���*6Ǜ�����n\k:��v�*i�_m�M��13[�{���ΐ�!0��m&�

&�����tr*���d�،;o�K�0R���;��"&��ōJ�Ѥ�`ȣi.��ti�Ј����l6y��5l�JV�0�nyO{<�na�.�Ӂ��`ͫ�p
�?��>���6�H�O,�#˹�L&W-�ޒ�ʛ����X�o>�k��#��{�ys��f���7�g@N��kaY�
�Ո�k5�hU!�F��x�R��6M�j�x��Uս7��G:b�^ֶ�&�K���{D���v��-Ĳ��r��GB��י��ۺ����CS�|�{`2n1ъ����/1v����|��S38p�f�k.�����nr��[��[�D>�-�GM�*��6f��f�cs�H�қ��r k��ų)��"o4�`�B��r|;�Xz�ǸΑsʚ�p��eem�c�!����cC�2�z���`8���ӹ�u�v�(��3��>W���qݻR�� ����)+�&�{���Ԥ��ì8�j�L;���kyʴ�i���9ܐ��j;�MPw�H��o.'ю�O_��{>e(eoY�umCQ^K�!VѾ��FG7ѵr'S�m��Нڨ����	Kh�8�v�4��U��q^2:��Q��*�
Dݍɦ������]Ѧ��H�G��n�_,�Uۗ[��m�]JĀo
�n��_9������{Fs�z +-�.�>�߻o����&WS�3�f�Z��c5��DL�n$���cʕn�,�l)�n�?	���]�ވL�Rx}����c�۵���>�V�ϩH'�L$vZo�Ư��?�U���=�i������;�u*����*˰h�S�RI�읗���`_7�f^N�� �h��֋�̧�T5j.�Fఛ-�u�&8zة�ğ٠��:�>��hwC���ޤ<p�E.�	�ژ�an�'
�f\&C�����;sI��=1��q�'���G����2���6u[�RlY��ʔ;���B�~n<,�wsߵ�k9��Qө�� �vZ�cr|�+k����Gj<kng�$��O��7N��/zǸ��ᮃKs�q���i�뢐;z�����4�� �Nsy�
��V��c�[�p�8d��w��B��^=�a��U�.מNœ�q�����a��էc"xU�^�����)P���߇ڕw���=��<�  #g5xg}�bc��c�0�;W>�L��TU�8�y#���R}6^�z�f�o�B��ZC�5�9s��/�����ŋ@X)"���&�p�q���73e5�����ׄ5�^j�DH��b��>8x)>H~��˟W3�s�Mk�Z6�J0ݲYJ���+��߻�5�~;�7]�����S�z��:�ٮ��Y�L��r1����BC��T��q�ś���I5��t�]^c�Y�[�n����O�MZ|\Q���ϟ�I|n�L��������r�I�M��Rs���諙�O�������.*n��'�
�at��c�9�K�}�7����A����e��ڄI�Yv��'Є�Š�JPo������]�}3�+W�&o�f�O8纯���|�O�} ���=�j�T���b%�4xw(�LqAn9lltu���k Ŀ ��<�������P��wpY��`��j��'Y�X��}��=�Q�ݡK�Oy�x븪X��֢ �L��s�5��� ��Or��R�����٣'�������F���1�}���Ρ�341��+�̑Ťb�5��s��tC�6�h��V~�ph���.[���9� ߾|>յ�����+d����>G��E���o!4�x�v1(j��Mh�k���b���Z�s,�X �H%@�Kl*s���_g����~w�����f`�C�h֊��t�ϒ��8�[OI铳8�r�N�lXr�BX�Ԣ��s[ږ��Ej�.f,{:$y`=��mGZf���'��c���^���!��@�g߳�9W��m��u����ݭ#�_��8�jS���k�ț����SnEמ��߲�H�0�����H��ٳ��e�@]/��<)�)Qw���]{��w���cu=X`�L6s�j����ȝ=��Z��:��$����j�[o�Zx�� �K�"�����ˡ�p�/%>F�M����_����F�>ź�x���wK-��4�g9����c��ӎ�Vd�^�>9ku���y��[������~�� P��������������oN��մxL��4�rkpO	;��裳{c9pc��N&���DM��A�ɵ�I�Õ�_z�g� y7���Y4��1q}~�?z�4��Kp�f���n��lȝ�DD��c�^˟W��';�/���cO/�'�}�9�>���y�>�YV)ĕ[iYI 0d��Ab)H2 �H �(�J��Y{�-;�w�����+��u��hf`
�I���C��R��R=o4�s�Zy�1DeZޔ򒝻�>�����l��J��vf�d[�ּ}��?b�����T|�!֊4�]C�E <��⦽}�5�ܵ9aÔ�`�u+S&�NE��� 5��z�Y�+�xES������:��Tu��3BP}݊��T�r���'�9���|)l'���̛�vr���9���lߕ���VB�Ǿ��ֺW� �L��4�]��w��&�Q��Z�R���g����9��g���9k_+����(�ڋ�.)t/|7�d�TG�:�`S�D2�#�S>�bփ�����"�H_?aX2F��81��O���s���>�A�f|#�El/}OKY �!��.�`��n�U��{�e�gþ���4�����t��5�����3�������OA��~�_:ߙ����[�Z:<5�
<!:��#yR����>�3㸢�֘�ś2r�5���xYP0�M)�u�b��!�+$
�Iae���2]�v�q�t��m c��&Wum+O;bf��^�pÒ�/������T�g�ؒ����iS�h/6X%�[�7j<oP;�:�L�=PΑ�A��ev/��'�"��U F������o</�w����2��)����m!Qsd�;�����YkLk�q�ꍫTr�ve��ዱ_UNI��ߤ��=�S�%�ɞ�>*i	�.F3��)�!1O}fF���2݂�ph�|P;��h�ffj:8%�q���� *����<A �Tdb{�<�=֟k7��S�5���C:q��v�,7j�3�_}Y����n\)���ҫCR�g]� |{�9�>pL|*��2|������Q;v���2�q�xQ[��T�L�3ص�N�N�B����cV�v� P�� �C��}?l�C��^����x��17�ěϗ�3�Ǝ��x�E��u�街8G3�S~�ϫ�uNR�}�^�4�C���IA��^/���c��o8Z�J�3pr��B����>T%cFf@�i�XA����7����n�H6��C4I+���Kj��1�Qȉ�я:�rV�E��]X�]��i^iK����B�>v���6�b4������9��&��2l�i����p���䵓�܆��Ǿ�}�pu�;g�+й1DϞ�+y+Ã�#"��Nn>�w*#���PE�N�1��$Y���9ˀ��Ǿ�6!��M6Bw���3�E��҇Nl�2��h���r���W�*�]R�˥��{*,�=��r�r2=����bE�/R���_��39ݾ�D:�xK��L���,'sU�|�?�J����v>�21��������ju��Q��9���`{� >�z���`.�f=[��	j�3<7�!An��u�s���.ʹ�Z�7��@�T
:B�>K����77	�K���U[��W���D�X1h'p+c�l�oHQp�'|���V�i]t`wKj�Ғ1��������B5q���q�g� ����ąF��R��
IY �E�ٙ�elr���^DY��������K<�V��AVqr]:vn$��7ݹn��Ke0������m�pk9��"gz�'���kB�{}�e�S(��^�'���P�;V�u���\�7.����K��P��Zv�<Wo>t{�$�2}�39���w�߶�q�'�r��ʙ�����M���|��o޷I}�H�}�_l�� 6���W�7��[;���@�l�%����0�Ϳxĉ�l�`�i�w�5�k����MV.��;<]A�[0��ْ����#�ME���9Fa�k�/���.��Z�{#��gT��#�оf�r�/���fK(���2hB���x顊�t]u᝚�9�r	y�>��g�P�or��f=���+�tT{�D4uY}q��ʑ��_tZ��_m7��͠�;M�̇��w�f�G��\(:�r����}��߬}��݉���.���DI��#BC�!R�C�-����Z�칯~d�9C1�(Zc%���{�>��k���vixb��ȍbY՛2Vz ��2��F����厈{Y��'N��6���7��r��.��s*��w��z�z��ꄪ�)5ѦVƛ���f�i� /��<$Vr�ŏ2bR�lU��'�K�M�GJ�C�q(���ssd-u!�Vc6qS*�oF�>7��]b���w��V\�z6J��ݱ�{�[�����<�.�qcT�w|�vk �w�kS�	�b�ȵ�n@�X�}�\��y���
�k�U� nO���BI7��"w��ߟ���_s7~3�r���}f������:f�c炴����p�[�6ʱ�D�1�;�H�����H^WP��lӥ�j����VĚ}%8�>>-��=�u}B�4���Y:��	�"jGϕ�U�jB��w�}�G�����;�
���C� &���X~[����sP�¡���^��=L:�y�N�w(~�5+��{��?EɅg�_3�o���O�K��k��fw�9�M=���tw��k��_1�~�B��R�"*0�
(0�F1�Ȱ�`2`+�!id�*H��X��1�(2# ����Fe��7�sO﹎��Wr�]��Q�%����z�ޔ�}`r��jt{6���C���;���C��悒T:��ݿ�d[���ݻW*�l�^��{:�����Xb�֏ajx�Ӱ��ؗ����]�&�V,��S�	?<}]���ryta��OQ���3`b1��uϢ�����TV ��!�F�����G�~c����l>�*w���盗ﯮpzgd~����m�Q29n�<!���ʷp{y@����,X�ĥE�Tw�V�M�WQ\rq�t� ��a���X�L���o�)GQɀ�Tn&�Z����xR؇%���,??3S	����U���^�����o>�$���7��j�]�U�}�y��=Ǝ���8�2�~a�������Ȅc���-~�q��7�	�$�Ƣ���z��t BL�����on����2�N+e�{ִ��>:��R OGȢ=����z��eWTg��s�1e5C�f�	�+t)���e��JQւ�^���.�^K���ڴ�`�D9�:C�ۜ���b�{y�F�;��][ڹ�%ic
�D�XB��z��.��yϻ�)�������פR�iz��D�D~�U>��PΤ�¾Ā�?sV4;Ju��|��\�c�k��W�|JX^�N��JI�Hs�c,6c#z�������i�׳W���e?' �":aJ�G�Qs)���vX�J���w��*(k�6�)lu�:<lR=C�d��~����i�*�%��ϳ���!�Qe��^����+�>��#|\�Hsc�ƌ�ǻ������'��(��ag��܉;�LNy~��ɯΟo�����	��}�9�� �+XUc��ۮ^@[,���Q��Le���"���5����T�_/kw��<�n���~��H�>��?V(1^�u#�13>q�ن"=/�<��S{	��/*��q���[���e-5�uˮg��Ϯ#HI8�3���k�O<��~n���r �8�R}4���a������D��2n����ɱ�5t�R28p��V��F��6ap���`o��s�#�V�c�רQ�j��H��^jH����3{�ѿwݼ��������g�+[��)�zŊ{WUwB��c6{�n��sv�r�"����y�M��\]31����t�Z;�GU��(�O`RuK����1H����Wf�Yd��ͮL��0�z�t��Q���o\����E�in֡ZjST��S�R�V�m�AX��ʆʾw�o��H���a����5̦�L��:�"�]��^L��&Цc�;њ�t�������v�y�7�i��q�{�4��Kk)a+* �=���7�D5�\Ju�K��C�w�3ovs:�w�"�=�@�@�ˠ��B���y��:���7�ng���[}{���x;*���
��],&jݹ�|�68I�'�xk��	D�ݷɫ��������ߙᇘZp6��X]�DKI����1[)7��Ε7���ְי�뉵_;�u*[��5�CJ(�U�Sw}�/zbK�0R���)�]`�Ձz\ްt��5�n�TᗜpB���kV�9���ލc[NLl����d�u7�JR�@��[���tvŻI�ut'm���e��H�}#�gcy���m���n�#'�P�"RV��@J��M���^���]�͒�36���V�U �E�k�ܜ��T�B������oFf�^l�/��|kyi��i��q��o�b[;+��Ǜ5�t�to�b�ɢm<;%�D�n��g�FZ���x�X7^:4��Vv������������V��k9��)J�8X�*��N\;�6�ŗ�S�Q����x��6���{XWY�W��W=�[`�<e�p��.�\}a�+���0^!�\�%��K���h}y:�H3)%��ˎ��m��8"�Nғy�Y�{p��f�-{8�d�'et<{{���.�26��+�ƃ(�u�5�څ	�}ݎ�I�/�:s�����8[���p;�3[�:�^���dj�u^�w�4�����R�Va>dW���W���]���qف�Yt��LaR��{�VJ�r��2p2�����*�C�L���l��Re7NY���}��{��so�^K��A����&b��E�Wf���4�1�JN���^<���V.mlܔ��W��K���t�t�ST�k��5R�mcη/v���^f>����5�w���QS+-G��\zx�;�`7S �r�Ư��юQZ�s\�q͕3�i���B�ιt��O`Y��nҫ���̹CkD�ے�ɀy
���v��q����D���{���S��>W�F�݉R��z�Y ��-��'>�ܽ-�{���vȺ�AZ�h�ͧ�^u���L�]:,��4��J�r�	t�6󟳥�O�e�cU^������]��Q��ի/����v�聻ާ,�WY����v���8�	�初1~�f�b�A��2ZvP��'�{��k��ao�Q�����B�;��'yt�����w�5q�]@]qX���[XK]+�`($n��yWK@�e���<�ad��Za�c*�#�}W�OO�z�fv'Q����5v=>��d3s�Ȓ5��vY�	R��l�#)�E���Z��	�P�U��U�[�|��y��i����@�[�oG�����m3��C�N�\��kU\��ᢗ���mЍ�c��,� ES��)J�>���'����w�����>��;�q
�iY-�X/�~/�/.xOt ��P}y��W�:�[�	=ї�+�w3y������|?o�s.�_�Ig��.��?k��2)fa���V�$? #�(�s�藶o�/U�r�Sd�d�oQ�
��zkgs�]���ewn5Ӓ���-�����uw\]4�Ĵe����C6X賈u�GR�f��t��?G�'���^����l�����;"�Se�
ޓ���W�x�r�FE���	����^��h�V��Ǉ�C�b���}������ֶr��`q�g�A1X�A�v;:iس�X�;��U�͎���-c������brl8�mUo���p�.��|�yt�Ĩ�	~���5"�W��ի�ވ5��VG��f�Sv����1�[��z��Τ拎�{�?FH�����ܟ�^�����zu�*ع�0�O��ڸ^�D�����r^n!C�e1hV��������p�|��K4=6�ܕnM���w21�ȸQ����h�\��A&'�97f=�z��-�G��C�撆F����{�3��o���� T��ۤ�0������?x���i�L�/*�O~�3\؅Q�?9��F�'y얾ڠ<6�ڈ�}̙pfB)��,ee��a_�e+�}Eq�&��ǥt��_q{e��:Sը�Z��gLg���R�C�����m-�,:1we��M͜3d��=ٽ�Ol�F�W���ѹ�Z�	G�욞�#E�x��/��w�-FUZY��R��c9��I�.���i�֘V�����PR$�t�/;���9����Ϯ��?D�46���e�k�>��#Ð�&/�K�X�=;qN|��'{`�C{b�`�G��Gr��k7~��8j�{s_���O�v�=�Z�K�ev'DDע�0ȋCC�]�rps5���}���K�C㩿wntظÈ�g��3�TZ�NW���2�������&}*<^Oy=̾�:ջ�b��V�J��}nBg���q��Ud��)��NfOa����!lŵ�>O]v���#ʡ��@s��E��4�=W��3���9��q*h�F�g{N�&�Nj#_S���0)�}��ї͞�����7r������!���l�+e�z���u��4cg3�wY�1�~f fP�K���W)�Vc,1���Z�ҹV�+Dr�bLLb4�X��R0�eh�+h���~D ��U7���,������oQ����GU��.�1U�y�8���v���p�\ȣ��Ik������^����\sp�4?L7ܠ�_?�\��@F-�蜟n:H6@C�͚x7aG2� H�H�0�X1	��k����`њ�:��Jx�&���\��o���n��������-����yK� ���|~�x���:�3��{ǖ+F\ WD�=�g}R/˼z�/#�P^Η�ڟyי>�bLV��PR��뙎�aҖ���� �dB�+ ��5�/~�\87��iS�R�q	a7Қ���-��]uF��o�z��i�*v��JBtY �*7��a����Z�n����U�|���I�{[�c��[�x�л����`�&��${��=���aN{��>�:={:�q�����?i�?	v�� M;B�:�\$��;����Tb�\�������(�s�Q����	(�bh�|l��Z��?X��\ʘ*$RB�Y�`�����y��>˫�5�MЗU�=S��V��������r�ǘ0�i�Z��Me��Gr�*^;�st��nVYM�a��=��!ȳ�
 ��@>���Z���|�DǥV�>�����M���̬�f+t]IY�T�1���l��3��fn�y@�Y��?ak/$d�Ǥn��!�@�R�T<���eQ�l��ė-��|��:�ً��8'qg-}��zc�'���vCǓ�gb��0>w��#�!W�����ҽ�2=4�e�:�3	��:h�v�:�/{��?'����t�p.v���޿��@�s�\��sf��^~��pa�������Ć"���x��h��	�Q��^�y^���1F!>� ,�ˬ��=Et�}���ꝏFx���{��S�"k��V�-E�Do��G��-���vo*�E�1mdHAn�0��6�8};�B�|!�iC=_|*���}�ww3*t���Y���9�E��|}�NJ^Μ�c"~}7#x]loWN�2y|�6"�T"h ?%��jݘ�V����U����(��X۬h�a����A�Pk��ab�U�֖b<�n��7:J��5��w�\�[;Y���[.��q�_�&J.2�rS�b�&��mh��������W���S= �^��_|�f����V|n��)��W�Ps�E�aW�n��M Z��e�#��~��VO���1�cN-�F��Ƃ|>o//ɸ����B��K��{�{��nΚ1�D4���㕳#SӑR|���m�ʍU��`5���+����W�<�E��~��Q�$�F�1��Cal/h�,f@�#,|e�֟�HU�.���#}F�-[k��/#־`����_С#�r�L�{8��0p1P2�n�g�Z�P�Z���Z\�86�*�s�r�Z���#��mYs#��1J�4xn�oB�L�������gp�z���x{�~#,]�N��k�:�C�\*�� zrh�zbϯ���<ǵ(ґ��+7���a��e���8~7��Wk���n�r�|7O�{瞚MD�2dTH�_ct\S#V*��! H�l��顆�k��u����v�fp���=h��][���s卫��c�j���I���,G1���"q��r-"�E�I������/�_T��ӂ���b�Ãy�@Սf���ɳ}v������}�>�8����ߨz!t1Gd�f������i�U�o��8/cH��L�n��H<��I�?[kt;���Ţ���W�\�kY�U�����1���#��  ;2!y�)��n�pP��U���!�X[F]C�O!H"4^��Y@��0�c���\ɗ�j���~�ﾁ�U��|1Vt�(97��NVMǴ�o#"` `�T�g�^E�m/�{pkXk��q���oc�{�{$ڔ8�٠�>K�P[���O�8��H�~�^f���4�w{��&:i��`���H�s�5��O9Щ���{�����`���c˜l㯿��\�=�����K~u�K�҈^rht�R�#����l�Y�:uU:oqɔı�c���ʄB!�o���j�?���!G�2�[RH�2\H4rVdf	q�P�B�,�
�dJ�/o5��u�ӱ�E�]��;8�dS��˷b��[')y��w=� ���`��}�G�s]mp7��*�:��on
)G�ٷ����62�~��g�z�_��>�]��?j�Xk���^yS8������+7 ��_����Gmn���	�.�5I�1�k?����j�n��Ľ7�g�A�K����4�\��a�B�s3�͆$3����a�]��d:����d	0��)��|6!�=�yL��w���f�,"a^tE�s肆�Ҭ�����Wfiter�S���9�{{]ĉ\���bR�2�mF�}�x ��A���d�b��3; �O�w@�KT��j	��&�6��(T�_�}L��g*�R��
��cxQr�1�Q0�5��<>���4}�׉�T�1]�����Ю.�Xw�Yu�~�L��.���[Q��,��5K�yDtC�޻���3��|����1�}�Z�:J��c$*m��6��J'�d@���CkZn	p�rTel����E��Q��J��K�k�k�<�s.���)�١1��O��H����C�<�)(;�}�_"����I;�Z#�E�sY��K�9���u�eS�񘂷�>��l�4w��m�H�Rf��������� ��"�_��o�1Y�2=>��}>9��/蓼s��ԧǬ� c}�Ϲ�5��?�:[#�����ع�+|�̘�����<�O�|�'O��v`�A��D�=u�X��w�p�p��=�=��Lؤ��8Qr���
���j�]* ��:�'rj��K�j��~���)�Y0�r:����y1�����D�٦"��t5�^\��\by�����4��@nc����Z�aC-:i�(;�̯ ��#�~����TY�fϏX�)Y��~$������_�uځ�z? ��3.�����	�]�u�cﾼ^��i����>�^|b�7����A1HKs�ɅS�).2�Q�������N��}�ރ���mgֺ:.ЉH�,CҸ���V�� O���,���;�߯�1M�w���ő ~_�x������:�n��:�7JY9�ν�<2�����r�P%����P$x���mfo\{����NL�]5�Mbnɗ}�B�+��G"��5n����XԄ^!Jea����R��Q}�L:~_�CmA�+gd��m���ky}�y��w����m���rf!\�"(9Y��7��be�(`UۗY�\��D�����,.Ux}����)v�0��/�Ǿ��q�誜���N�KϡʨZnv����P3V8��Mj�	
_G�	LJ�G�؉ԝ�-`'�7�uc�}�q3�3����~�4�U�7{&08�PEWomx��[�J�sTq�<��yT�J��N��~��5�t���B��~��=>��S�����T��X�c�D��A}�]J�Ӈ��K������1�Cȶ֭U8�úk:�6!�|�v��}r�0 �o�,�����ǻ�������=�=�&�Ť�p��+�5N��,�[��#�]�Cf���l�ntDW:�.V��'���l�̤��냮�a�ZX����y�"=���nv��� �� � � Ho.�|��S�ל{�3[�Ј����2�Gʴ,c�����=~���2{��O�l6WC�!�d��2�����Fr�Ŕ�E����w�p7�'-Kͱ��(�=�v�G19��-RK��r!�B��G--T/�JF�QW�g��է��
���s3Bq�/S�����ͽ�:���5����m9�a�%�r���L*Ƥ(�J[h�v��)�ҧ������gx]��13{�;��)���7�wn����&I(�����T�)��.���f��8oq9吩�sV���Z4%PU��xX]؝�:�v�N�����ښ�W-�������۩����m�<.��L��ֵl���3��w%�fe��߆�28���bs{�	����S[ͦ�&XX��\]�&��MoVlJl�6eh�M_S��*+Sm��!��37*�����=�p�D�E�y�nL�HTY�����i�5����0%4!���4�-�B��Z��9��Y���B,�xl��v��������^t���O=��nOeJ�0��Y��%E&�[�c.�\�uO|7�U�:�6�7�	:��uf���I'wI#m�;v������mrD�|�h�g�urDf	Nm��C��&�rg�����o\���͇nN��[�,c������l�Q�ɜƲ��h�T.��oM���4���d3v0'[K/���@�:��9r5���3k�,]nԔ�YW8J9�E��O�}{I�Vk�\�ɚ�|���g#Zx�פr���2f���{3�1q��֬Q���֭.���j.Y{Zy���ھA���-YywQ��	�����.5���u����z��"��.�3��t��·OXM!�;4��,Vw@�+Ҕ�uh��S3���u�ty}�#]��Zs�;i͝�� h�S�L�{vw�E�N���@3Os��hoEQ�C�z�-��e����=�E��j
@&U�6Υ��[v�7���D�[���c�K��"�_�Xsgf�u0Tl�W�$�n��R�l]���Zm�	y����K���'fG��+�w^�������	pg%��-U�ty9d���7�äF��9]�@m��*�\�Z�Nì��/\[�$ʎ��\���yS��-��vA�����k���_n��V�ٻ�����LO7(�1�b�{F��YW&���g;n`�[Qˬڎm�=̾,:)�)�ԚOp���D܊Z��J�(�޺燣��l��7�ojX��Nb�ʚ��5psx�~Y�ʜ[�2���1�:�:���q�A#ci�9���e��^�M���aq�W�1�w�sS�wN�t�<���vQ�\ߐ��ި����v ]*�/���gQhs�܏I0&��V�`=��1��/�W��<EJ��oF�هQ?��bGڬ�:-!��2b����L"�u�"�D�s/���V`q���]���'��@N�T��tK'�M2��L���w隧C�I���3>ֱ׵�^�c��p8�����%�0�m��&/��U�f<���g�4o,�h�{�w{���WY�~��B���.�O�o�����\�V`������P�`��J�������0H���{ڣ<ǽ�}Rq���N	�˹uq�����*��>��I]��`�\�K��W�B��j;��ً]��@o=S:�&w�d�	�@�_s�:��8sxR��x��dK8ȨM-�����W��¼*O��VW]�b��+	{�,]J�.c�V�V9��w��U7�q��X�w�	d��u���*U���^o�}L��y������W�aeD>�a�%E��!���=��s��<�69�{�י��)��u����;T2��+�S�8���SPc�4F��m��
YϚ�u�)��e�2G&�N"1e:瘧[�w;�s�T�PC$�ئ��.K�k)&^ĝ����㏷��`G��M7zȊ���K�v����v}>��1���:7pv��;���6�n�ނJ\g�%"��F�����+�,��z�˕{U���V�<:�^S��£vܓF4�ixޕ�}�Onjc��g1V�:�`D�˗^.c�ꧪ���f�sy<��u����;�}����6l�~��1xe��p�f�г�N�3t�Ss?Q��[[�̼�N̓Y�'O���V��	�;p!t	a��}�쌞ʉ#oVsG�`��A���ٞw��Z��C�*B�a�c��S����B7��*�5�w�}��׾
��ƻb|&��#�O%Ǩ\e�]x��qA���{�;�����P�NZSk�xj�Y��lG���ۭ�_\�a�`@d��Xd����Z�*,�"��c0�i�c���#-��ZQeV6�̐�@F*�XbC?{�m������\7�tČtVR6eb/
�n:����#���V�]]���i����,�$�y��7���_�+�;�W@�FN���:����Ff�HiQ��p�kkzܺm���ԛ���r���񢺺X�$!zr����ܽ߯��{{��/tz�F\��1Qiz/&�;�D����GeO�;%�E�ػ�©���W�L�C�龛=�ʑ��J/�O�8/��C���z�%/�;���J�#'iK��%�U�OvG�yg��z�[
���TB}���ҏ;�u�����;��z*=����{���<a�Fh&F������Ut�7�v�D<nCal*n/��E�Zz��!H2rlx� ��LTO��]є�g�t���O`)Qb<W�G�����Wx���Kr��C��p�3j�hnJ�����o/⟀}��k�Y\֯���H���C~c	���r�g�m���{f��=��W�wzS���oOi�� Zy˚���%H1,H��3_}�.��{[��Vk�EZ�6�N�W.ɵ�xF�ڍfe��y�tf${�'Q-�!B�����.ʱ[;t�vh1��"���l�T�Z<��^�
(�����M�å�J%LI +#3��*�Y�S��:�șTDE9'u,�\Y�Nwu;�L%i��z�l���lƵ�QV�«�×�.	�|~4=,lb�ϧ��p�so!��������O���֤TB��� 1��V��rz@��X�AooR�Yo-Ryj8�A����u�.�){��:�;��zQ1jx���cHC�8o�3.ПI�Yߓ,�!Ę/kb*���A�Xm��'��鎿� ݍ���\�"I�8uDK�;�l&gE�%���6{��}l^2<�xFj*���߰��z�zk# ؿ��2&o_co�i�yg����=����߳C�<1G_g�F�B�<�����4&��Gjb.�B����dx��hz�����r�?d��a$�'w�y�㯯������D���?N�/#⊄~A�缗�xv`#�\U{���1=�̭h�ަP�v��C�V�C[9��%+u��M��_�z�ڰ����z�8mS�y�yN���z��&'�3����*7�g���΍�������Q�e*^����Gr��C��G�D0{v�q{&,��K���,��>�Y:�<v�ի�����I�9q���gv������4�+-���H�V`4�ǆ8��K���<����4
6"����|NCM�)�F���&���ǌ3p�u/)2����sY�E-x�r_WXDO�����Z�T������>������ځ����;�K%�q ���-Ôq[�L�vv����k�ɞ��N�>�B"^��#)�����-S�Nlo���_ν�w~y}�n�r᩾�e8�A�cnD	]�ʃ�J��	�L�i|V�>n�d
����[���+��I��7��ɷ?\�}�~�M��03��^�fҵ���@��4*f!j��h�M�z��Ƞ��]�UN)۾w���uZ�Je�,-����jر
�Q
� ���e-�h���K)[�^��9�=�uP]2�X|3��[�(c�����]@7D�wz!�1hk� [b3���:S�v���c��m��뮔TKe��m���ؙk�U{�os�&������e։�tY̏O�
ߣO*������r��ED������l?D#�^�e�(�B�_�
�}�͉G\x���i}$ƌY�>��ݙ-�ag�=�4ʍ폽�y��%�]��_L���E���~�a���X���S�ߢ�Y��.�H�������tгU�U�XNXɉ�:
m1jӲ��d�7ȼ����ۜ�%櫞e�:Ul��ʚ?t	ت���z �ƅ份�r0��G��y���0�ј���7�_"�J��p�a��"�)�z��������{������h�1
@���J}���O���ε׆��������.��:ˎgK��ۦ�0�M]d�a��+
ի��Ε��"#�)c��y�z��W�,�p�����Z>�����ʞ�xD�n����z�8�O�q�
2GXaKd	I$E�
U�����N�Z�Z�k�̫�%��K��6�>ՍgP��T�8��c˘��nԣ�j���?R+魕|�^i�v�-��cG��C:�7���"�|��m�4`�v��c^�E��<\k��)}k����[���~��9��!��@�`����7����}z��g�.q&gVN�yY�ܷ�Ê��=	s�����"V�{�k��P����Z:�V����o}Yp�v6��j䰞G��Ԇty��R��L쇾r<bi�>�Ip��B{��$6�{���?$b�I����|��/������'����l㎗����3]!�U��v�J�¬����?]3x7秞�\��M���|מ����^��{��6�|O���v��k��Rr"��=�������{��O7�	`��-�̮��dD�H&,ƃP��Є��{,}�k��?�P��=���՛�7�)t$m!�L�)��E������gj�4*��E妝��n� �O�QW�TF�@ͱ"w/���'!�_SQ�(L�4�\�D!@�
�[V�,XH���3fd�`
1�Z�H�"a$�bL �&[������7q�o1���~����H܅:�]�fn@zvS��':7����7�b%zM�u٫�gp����)�6`��|�M�6NY*.6�S��D��߲����|��f���V8�����1����O�g�
�àx�����=�I]��u�E�8Su�sQR�F9���Z\��]jA�ϩt���Vh���V]�g���N�J��۫N�uM�2��إ�ܚ��G��ޟ����֫�JA_��ڧ�*�����7Ԓ�]~��C�[��� 鈺\|�=遹#��x�A��0E!��O������߻���{�������X�ʍ����X�=B���tH��vuis�:��׼� �`)>w�&� �51{2��}��c��]v�1��f��|�D�p�Qc������d_��ǐ�N%���4��˪�x�1w<�GK��sP��
ˁН?�x|6��\У�Q��ƾ������.���D5q.6f{��Cday���Q���({p4�9� ��̒A#�~�HRe���L����J�)����K���5>W��PE�h��#�Sm {�$iw��lnWYۣU��d�N�eugR7���}fV�7	��$k��.�ѪVY�f+7�����`|E��r�|�&�?Y�J7�d:�.L���&�F���%�H�F��ݜެW|BІqgTԳ��P�A;����'$;~�ዻ�ڠ_��/�DGy�_�!!��	�y����d�>����5����h���H�KO�&7�j�,�zJ��݋�}��}�7�ܱ5N.���R���m0m2��D���ΰ��*bYˀDF�ػྻm}**��y߬ci|>�#:���(�x���[����|~���E�!ih��ɏf�d���]D�\W��*#u1y�'y��~sw��i�;�{�%:����o� ���?�/|�����<:�^䜄�1�W��i�����< ϼ���!�C�9���=�ۡ����܅��	��3���"�V�|�g�ǒ�+4%I�N,�_zQ��Nn[� /J�aVh?����Y��#lq[��d�R��e=p�h��}��j�*3��n#KZ���(r��ԩX���$V�ۮRr�����%7���a~��f�p��vr���L�y<^r��H�g�>]BI&}�}�ا�.w���.��]�oo�fT����e�4mԠ+읷b$!	,�O��-�z�,��{��{��O���oߎ�d�A7>��������,��}�|*���g܉Ѡ�\�Or���@|{�xj��"���mWY��V�j;.����q���7���/����=����3���s�BG�άߪU��A�vK��!�D��ځ�lT0n5Yn���SO�D�ݛc��fZͳ���Ħ���L�hD�n���?��S�N>��7GY}���r���N�d���uO�9[3��yH����Dn��͌���U���@��X^P��i��ڢh�(�b�B�$�=�ݎkh���k�:��UD�&��,�G��$ ���+#����j����L��曦�/*�di��p��<�.=�Z��G�k���j5YN8z������5{��{J:���2��n��k+��Z��8�rt6�sN���Rr�@}�ě�A�fZ_�K�.oO�f�i
l�Hh�h]��&�#�8f4%Zb���[f��f��:�#at-s��K��&V�hV���4I�j�M\�g_jWK��S�bf��O� �u��^�D��`���.d���N�
�֢�������ƍ4�р�k�냽U����sunb������s�k+���֎�{�j|-��Ux$�1m˜�9�|�iEAl[E�����sFf��wu�ٗ�+����Vn�)ҨVnT4h�����c�+�׭ߚ���^{o��=h�f�L W���E" J�G���P��V���r��(c.qѭl�3Zq����wx��w9��1i�t��Z�`_�*\�mj�F���@i���!aiE�i�h�!�\Hk�g�dv�n�2�'2��d!�1٨�n%�oY�[R:hۍȊ�3Z�'m3M'�7�\JVT�s#���sr������2�SX{�S��u==$��m�ےn5�/q�ݻǋG^�����"��ϱTΏ�H�fݢ�c�\��7y���j����z$�/$��<#o�-�;��FNU`�)��ݼ�E�����+{��'�VB��g	}|S�5@�8�Z�t�.�MAHr�L�B��<dF�#�8t=r���nDۓwI2��`�te`�w.δ�Z�:8U7���!gu�U��Dmp�C���0,�jK�c�]ZPKV�fZ��mw�ڹ�+�i/::g�]�;��:��7u9����7����W=u�yk�,�Wo2����4K��#s��y@��%ӵ|i���A�Awh�n�T+}B^��o��@��e}�ث�f��V��j�ڷ׮�z��kβ��pj��BaCyXq:�̥�ݧR#�evca�l�;�gJW�
c+hI�lu�h9�Q��{�m�}��i4)&��9����Bλ4P���}�j�f����5*��Tw�X7�Q�J�������"�78fj��b]�����Z��W2ӳ(m�&��ΆeX�f<�J,��3��ʠ}��޼��L��˧�*v� M���`��ݜa�D�*j�)uE��X�g���\�i�>���aSÜ��;6��%Glf����ҷv9�ӕ�V]bWo��zK�9Am�NLƻu2�2!�f�Y�(Ch|i����"�[}�M�Z�1*S]t�=��[A��j�=���f�(J�/�UT�?���(d�6�O�����K���W�($V{�|���6\1���",�λSG_l����p�+�Bk㶤m��w]��]�C$����ԝ�����t��<�1��G�;W��!{n��t����mr
�������q�O�s믿L����}ퟏd�j�<|q�w�y�Y�$�ۅ�?wH[�2<s�1]�+��m��]�zVj�>@��> }����)��G3rxr�w���_F�ťI�w�,�7�W~A��Y��7����f��~[Yk$g|���q���.������!5��z�N���
��H�dy�u���$�wI�����[�Vh:m�_;y�4eA�=�f��4������~����=���~>'b�`|G�^cJ�=Aq9]�B$aߢ���o$��g|�k��#��ަ>'=M�|��W��+���^]��c�\R��B��;�={o1֬o^�F�R�^�T�>���1��} �_g��E��7�
���4�
�X���N>��UC�ꆼ���l�4:#F��i�U	L�����q,k7�8;-<Z7��K�[�5H�n�&&�9��Hw
�Wf~�UnjH�<	 �> �}� ��4��Bf���I�]K��nw8ٵ�x�p&d�@4�s�c�|XL�G����#�v��TwϪ/��Ii���XH�:v���W�>�=�*��ۆߋd���������A�TPC���#��S?,A��V��S"rW�~~���s����ɾ|��������w�d��ʉ>c"���2�3\��!W�3�e���N[Ɲ��\|u`T�,
r����hڟ����@! �{ݪi̡��QgF�����P��8ɺ���#���F�5���O����n���������Ͼ��т���Nt��j��Cަ�=�T����3f"�:x�>,sq4vᙠ��8��| �ULv`'��x�G��y1s�B#����puc�#\�VnS���\z�^�KiOp�q�Y�VHF2
�
�R��"�P(��U�#)@�FD�AV�dB�Y,R�H  �B����VIa!R����z�|M��q7w�Oi�	>�V�kސ��&�7����,cy�o/�]�&(2�g���ڭ+"R�r'-��Ԗ7��Q*MI��Em���ڷ;B:�*Rk���p����a�{�l�jf/�z�S�ۜ��b����x}�^#�f�[C�X�3�p�S��;Y覦��R�xc{��ĽRk�=���w�yny�洟n�=1<��&f�m�>�H���G� � $�{���T��O_VOQ�{\y�ؘ�+G�y��о�ů1��s��cظL��t.�^�e�Jҷ����jzY�lPX��{W3͜MvPY'8q�|���P�������H��"�*\��!RQ���.�R�Y���'T�Գ��u,5ׇ�}��;(jQ߃���L��f�s�����o��G�J�&Ad��l|ڂ�6�u��QX�� ���}F�"L.p�^�C����!"SK��������W��\ִ��%�wm��Z��ݗr�~�7��7��v����Y�p.F��$*t�ݻ�矝�Sj��H���v�_s����}�z���_a��1�q�dT8z���9ˆbU��r�]��jH�����l���7��|R�@�\xE�1�p��҄<>����z$�2w��NoӅ�_`��rdϣ�6&�\���ngp��|b�2c�H����-YR;Jӯ�AǛi"�?����{���;�@��e�R&7����F-N�|�^K���$__M�4�/_��>�~ޫh!ؒ�U��R�s�裺��������ujA����	�[.H?{����Y�{P�]g��J�5���oS�*\b�ޑk%2�� nW��x��'ދ1ީ���Ng�A�%�П�Uk^�� �L}�E��s�^�7�Ӥ��͠R��5_N��\{b��{��4Ԣ���ށw.p�0^{���PgECDa�Y3g}�Gΰ�[E�.�PW���BXw*���YҪ�~4Ҫ�����/��"��#G��9���
¥w-��u�[�~_h�,����ႉ��QBDD�aeB�C)w}��7����= O;�������eS���b�-v�y>R�u^8;v�	�]�t��>���v��%���q�;�}��P�;r�4W�\@W�q��ݔ/Q�������I~߮?�)��3�ozC����WW�ѽg\BS[٭E�������;��Yi����{��2z�NWL��y��,�կ�o�}�����ř�X�ť�H��cb�����RN�;��[�y[\N8gL̛,�R�w���1��Bm��+�&=��:�U�,���"�Wހ����gr���\8q��i�4���(�6�:kל3��� � "��{�~ֽ��Y��fh��x1���	�[�[�Va���M���1r��s�)���-�iF��nl�����;���Bqd/|;�0�d����� I��<��̽|��4�g�x:�8�a\��: ��q�<�*�>�w��4�ER�vؘfv��Aڬ����'���n��|�z�o�����q��G�~�=�9��2�!FE"����e��+��5�T�M�yBE|��x�=���ݴ)�t���.�0s�;���#��7$�s��7����۝���W�d��[�̉s��ސ	�ǳ�U�!�$���d����a�U����b�a��7�{
�'�Z�YӓP�Z� <&����9�j�t��,1�R�ÊmKTl��m�y���(�°z�%����<�~�!�4�/Δʩ�qN:r)-Db }�����Ƹ%f�,���������c�W�Gv���x�墼�$�}��3W����ȚϽ|9�P� z�����r�p3�5��	����l�\��5�WD癀A��b��}�b��*��*��	y����q�U*�,�7��P�q�C'�
�ۗ����{9�2ur'r���PwTҊ\9i���gL�9��'��	�pk��[>�E�:�9n��>L/�I!���L��d�xK;�bl���[uW�!�xl�i��v��c��y��I���aku�{}F��y��g3{��ߎ��mQ"­�H,e!Q������;(��	ܸ7�um+x{v�-�Δ3�u	���gb2S��9��n��c��)��!�x�uN�{��"/�KM<�w�3��q���ND��D��^�H���F���=�l�#"�"5��<g���/�d��J6B�ԃ6�?�����a� @�ֳ�?��}�~V��N}��ٙ �-���%B .��T�f��E�S��g�Rv�*�|���I�a��ǽ5T1{E��~ �'��v��!�|��]��bs�Զ��PA=���A���]�L�3N��NrCo����;NC�oS����3��w~f����Q�{�=̛��Gq�V� ��ng���b��hJ�R81�.V\˦�9��;�qb6��Y+r\�V(����I��.a�=��|�c�;�C��!<�6����6����5]��X�/l�9۫�u�Ǧc����<����㿴8s��?!$����_����o�U�UW�~R���ޛ�8f������xbT���hB��X�!�f�W*�,0X�YRUD�)j��%IVD�H� 0��P�i}��ŗ�gi�<�>�W& �f�*W���B����^W \X��9oh��T�u"Tb��{�������W;oWrQ��fm���^����Y���ݰ���x�-�/����E��Q_k��p����
�E��0d�%Rޝ>ۋ�����TYܦ�������VY��P�%��XY����n0d#��<��p�zi��7@�ьu�z�����v����Y#�P������u�U����;S����R�թg�o�hH���7ФH�z�K��燯��Q��n�LR������E�D|~���f��b�Y{F幄�0#�{܇|���4N*���srʛ��=���� ���7�D:��ڸ������mv�ȋx��7�q�6��K��}�[]�O��+��{�3�?~z����]�Ḓ�B�I+"!�y��;��o�<u���sY����;y #L�5[�P3�{�WEW����5Vwv�Շ��N�ٔF&l��f��|3+7������T�ۼ�9�.��;��e��9��R����F�;����1������ >��~�u� Wu_ʾw��ٟ�XF��q^�僛�{�ݑU�a�y333ӿ<@��QQ�&z�?D�l�3��1ճ���ȷ�K�Vߛ{[��W�����5c���:���Oݔ��nf#�;�f�[�:TU��XP�wj�zj���.��N� K9��\���;����v�#ذǋH?|~��܉����Wk���?}����v�M�Cp_Qc�+��������k]��sW��P���;�������Pq{������n��{����VK|�Vk��>2˓2)\�["����d�����x����p��4��\���v�))vn���ƕk��I:%�'�9����3yw#\��U��:�̖٧3��x<;��W)W>�A�p{�����]�!�ɡ�y���y�n+6a��χ���ݾG���]D�'��8��~���P��'��VǺV���g�aw�-�ٮ�FQ�@��ȭ�>�u�JYǍI�7������|go��`Q���1�M��T3�xӵ�d-�0���� �}�ѥ���ǐh�?r؉��ֱ�^�T�8�Y:n"�LE�v����r�j���Y���x�G�(t�C�|:A9�4g��ҽ��иڅn�����5z}�z٘[�>�ok{xX�Q� �߾���o�����aw(����ك��>괮J��������gmvs&f^.�i֮"�fY�~��G�t�}���϶:��g�VT���j�s��D^+R�;�V���Y���.�~mpw�]7w幷�x��h<U|̘v����Zw�.��%uF�\�e Sp���YXvG��e8�.�,��xi,1wqu]>�0Z�K�)
4�9Cb~*��Jާ���j��\]Vt�#6	 �@�s�( I�d�[l�1�8u�R�k˛��4�k �wr�|�0�.�6ٷq��_�`��q���� E�H�1��
kWY�ਊ�5\��&�4�Ī���N��z�=�9�|�k}�(��w����7�o�-߮.���r=ܬ���� �Y����u#�P[ ��4����ݦ���c1ķ�¯����e�d2I��y¨qua3�Ld�������7ǩTw��ލ�$��p�SĜ@����=�_|3�lb���9��w��Z�f�!�m����iEk(��+�?���8O���˯4����\�y��c���4����y��5Z��k�',Tؚ'sZ�y��6�3�� )��w����](���Lz�iv�h�݂W��5�Rɽ��!���sƱ�}#m��wt���ή�%�QV�Қ���P9��p�Y5&�:u�fp)bjn�gwT��^���T��@��mή���^��Ȧ���)c��9���ý��O'6ʮ�y����\�S��B[�mX�跚��k�BP��׽��-j���r4�ǜ����8t� Y"���\O��rv�I�5������oӏ����������7�"�A`Q��[#|x��v�y[��2�b��v-!V���{���S����m7dm����4ꆬ��p<�:7OFcz�.�.*�+��N���#�];���Pf��<Ƅ��ݶ�KY�c ��^n��r�n���bw��L�$/s��h1�F��I�}M<�W.O��84R��)6kH��d��v��;�8dЪZ�ľ�X�s8���SX��*b������IBt�y�\�L���m
f�E��wf�+]e�¯�"V�8�{�EH��g9�,�2T[DI�9�<\`��i�[y�zK2�)n*��YD��)�`R��YOr��gew)4,U�G&-�i�it��nQ�����c^��^^�������۵9\������5�E�u��	4a2]������VO���ڵSoY�
��;V^����dy��nY|Z�(ML҉�����]y �Jޜ�u�%��y��.��O���w7��]�9�VJ�a�u��y�b�E(n'�-�	�r+�s�|�+�j=�6�6��Eg���ێ��S#��"���R��T��}k�z.�t �W�U��S{�_��~��ԺuN8i�(����_-�c	r�8��Z�)C��-VX�^��牸�8���=}�n��}�u�^�#5$��W��F����|*r��r���|���A��̣�
��F?=l�����M. ����W�!{"��[F�n���N�����������R�R�jV��
Zb��W��x&��Yٛ7�~��_[ȭ=�P���T-f�yG�%c{�z��o�vRZb�ތ����?|�����v4��ó|�m�'� �Uy$3����y���
�mNj}^�58���֦�f|�T�~�b�9[u���y�����#F��T�B8�l�w�q���{�6��'.��廥)eD�Uuun�a��W0F��Qj+�����Z,--j��AD2�1Z�Z�XR�Y(�"���-�Z�AEE��U�@�?�ڙ�����޾�G�gY{�7�xS���n�>Ȑܙyt�up�a[*s+���#�>/:x��nu��FB�M<����J�h|2��:<�U�t�B�Ou�������꾒)kg~țղv̺�S�K�ez���`׾����'�M������|���W��2u�ѣ�3z�!]�d�Ve�L�]��@��!s~�tZ^�y��緂�,����3�J[S�̾�{�Gs<7F����&�Q^p̻�{�� մOe���j�UԌF��.&}8�����q�����ߗ�]m]!������A=���[�j��q�G�F���MC5�;18-�3�2�� SC�^���������>Q�=�zNLYYz�9Rۥz6>�������}��.�_��fF$PD����_)�|�����sKvsT�8�:D�S�{v���r�ޅ�}p��O�5)uW,�s�����v�Э��س�%�"V{�*"F�M]���n*G���(���.�C��}�.�x,�{	�X4wkNYG���i�a�[l�)}7���&k��};���j�:�ǾM��åa	��@���;��'�뚞ƪ�{��  P���͉�LǢG����+}�1�!Uӻ��FWz'>�;�q���.n��}C��A�b�*o��^O�3��(��~�Bz7T�j2+q�{�k;�������,k�����9�j�r֖x� �ÌOO�X������z�lT��[���k�����U�c�]�e��`[���Daw��������p���k��=�]��|�$���]-�bt��(()3L�y��|��~!xT�V�X�6�a��E^�&:�b�N��� ��N���%�.��qU��մΧG��YOTW�E�Ziq.�c�[�rr�X9�f�/�-M�KyO��ui�v��C�ۘ�Z�	��ꈡ�����.�N��U�G�v����2��v*�{0e�bj�S�Mt�{�����w���;o��rJ��+��Yv~�3�����m��~PRУ{�rj��Ĳ��sf7[Q���� �}sAo
���VvtL�HUE�����7�M�Y��uW8������i��3�|+�
��Cʰ}�_|18���sxc�y��OO�qɏr��F���[�&��X�`��  3���J�pYn�Z��'<�pw��#�4�.*"qY����^���3��_,J�S�'�\�&Ε0#G~�٧�=����߰�Ȼ)W���&c!iV(�j�e���k8{]�x�����j
/{1��ͳu7��t�NYS�_'��Uy��Fi������n)(	��@���޽&P3$���G�ј�=�G0��j�<���b��W���=���y��
�}�po��+o-�w�0} }��Z"r��V19��5�K�����4Eu�?y��/+�p)�˫�xf|S���aDw�
�=��|���*�S:xus,)jbx�����w�i��U�LW�3�+\lqG�u��_}�<�j�v2oT[��4���jҊ����J:���4W]�mNO�X����S�������+��>d���d��x��9=9�z��F��!W��Q��mh��lg�ҹ�D��O��πf��B��s�f�L��x�̔F��gv�Κ�͝��blL��|%	8'fI�xc�yt�[o�w��&[��f��#x;�sr�\[%Y�m�������c�r-9����Ck��\�j�<�UǗ���w\�m��CLʝ��\R�\�޺����ݤ�^���tnw���l���;�Rp�Q�ញ�z���q��Ɂ�^�;�{?V�ީ}U6�u��}KX=�\C��\�}����@s�NNm2�e�~�5t=9�Ջ���=�e�*R�;a;���ڕ_�&ϲhkP�Ѓ��}��6F3��m��x1#��/+� -����ք��+�ګ�|>X��W�O�͑A�e��W�N�Ҽ9�w��Oo؜��A���'Q�I�|X�L�eP�!�d���d�W����[mc����'��l�[�11��L��ȕ���>߅�_�OO�o��������;��o۹�\��~ֵ�.�ˬ�֝J�CX0�T
�
1�)cd
6�"F8R-".	s ��kb�U�Y*�R��+.\D�ܽ�{zw�^n��ٕ�;�[����q;��,R�BV��@����5��l�AN�:��}�oEb�i��������k�jO/�b�^��V{f�W��!_y�wp�H��='f	�>����T���	ǆ��96��/Þ�����/����wш�Jc4�<�[;�ډ�}�J�^e��}F�r��N�'��Cx":�]���\v�'����6L��26�<�@}�خ�g���W�?���s��vM{ҍ(nu��fo;3:x���]g9O��[���u0>Z�8�~�����z��U��8@�z�Ts��O{[`����,�]_S'�W���9�6In������_�GV�|\��ޤ�����b���E{�_��o�����;�|��1�VR�w.:J:+�J�X	�I����!���Ǚ��/t�ƯWzM�F�3�v&�X�f����/:�kjCk:pfT ��a 0�Թ�MS`Ǭi}yo������Yk�q)^������]P���@�/�N� �^���˷W��i.|s*��]doLΝEo"�{2u�Y��W6��/�M�y}�~_o�A߫xܻ�"�Y��T���������3�C�> '��c*kp�F�yj-����d�����SQ����_F���]��fé�[S��0֪�����=QE�T.&��0��������Ʌ�����[j��w��|�K�d����y(Q��|4��e�ig�<-��2���<c{mH��$�̓h�ٰhOqdS[ޏ��N�6���""�}V��l��Y^��p�W��sb����t"O�d(\ )Q� �*CE�ܣ�s��c������x�m���M3<�w��,���dtu˒8:���cb�뤜du���5��S75�\���6.��k3����ɾcb��d�����f&�cȪ�.`Ky��ln��6hU����+{:���(���բNT��b�Yz�����A�E_������^�t��ŵYՉ{)���av���\l=��S�Kx;=<�r�0)w�^��P�6q�����c�yq�}X8�cuFш�h�[��Eֳi�������-��W���<��u[�]u8�J|x8��F�Z��;�.gT���Ə��D�ّ��s�G�J��\�U�Jo%�)�6{�����Ώ>�ީ�,j��?�Z6�}��%}�r��w���H;1�œ����m���[�3����y��Xy����:G {MU�ִ㠺��$�ӌ��5@*ER��EXS4��}�3��6�ʵ���F_R����a�+���of��N�)6&F�\����,L��o���;��yn=��5��dv���Sk�yNf	�����<�~wˇ�UUKy���;Ɖ��n��|B�����~�)f�_�����Et�'���k�G���+��gOo�q-�O]��:����g�=Xѩ{�w:�12��k�~���<R��]�w�vV�v�{��g"���/	W��̙�;����^`�ޞ����칽Q^ڼ�J%���������O��7�dU���"|_��ba>`�tX��Օ����p�� ����~��Զxg9�'����1ڣ�vIӺo��.�Q���S�w�gP��G�o���J�#�m���6dg2T��u;>]�Z�↹$��fT��K+�I�\^���zp�g}7�jU�ޚ�M�w���d�?V�������51Z�WVէv,Ș?��[Smucα�0J���e�B���,`��*��!�5�D��zk��ˆV&�;V6��X*���/���chn�;�L��V����EMHн�+��U�y��kͿ]v3&��c1u]�iE�R��*(����G-߽N����p�@�N�,�<z� j�쯺3)to��o��;����Y.�c<d* ��4Sh��WR���f�s7�\A)J�Z-��c+Q�W2��7R�𦹽��9f��3�+��d�q� �to�P��H��*�9�1�r����1��7��<����S��UEnG#��op�m� B�R5e�����\9�Տ�����J=�)w�7����޶mRlve0D޵��}޹��Ć�U��jt,g殔�x�Аx�����{}C����z�|w��+�����|^w ֹ�I4�WmH�S��0]�o�o5�m�j�}�v�t���q�{�L�"A�2���{C��@�)	�h]�Iyem&�ȹh��:�I�j��b������bd�gp!r�V��e.e0�P)�L�|�����w�gL�2�\��,�=�/?&Q�N���m���y�ħng6_&.R٧�'��%ۗTgE�k�'���7��,��®�v�{�kr�� ��)���*�ާ�hg�;04����Q�Ho.z_[u���wG�;�s(�|�ݝ:
s��/iix�`O�pe��x�)�dnݧ��7��:kYw��u���G�mct�ݤ����h��Y3v&�`�ViE��{N_&��¥�yr��:S
�ى+����5�wn#\��O.�e�ӯnu��M�������C�4���a�d�b	[ >��Y���J���[8Sx�rtj׵������m\�pF�wW��p��G�Lx=����Q�ڦ	Ŷ쫫t��s��`�����v�0��!��7mŮ�uh4u�L�N�w���'u	��&�e��ͽ�L����+OwN{�]�XTŏ{��£n-*`{���w>���WI)0,L��� s�r�t���=U�{Y�J�$J
�f;�}n�o���<����E�)�j^ĕ:�Ri�wL�u��fAij�)�tO u��4e_TGʹIO�FΊ�h�2���7);TҥwvKP�o��V*�!���s��7��Ö/���&�#��)�;}QbN諗w��&�V��a��~��+���-T*v7Ŷ��N��ƅ��[�3j�~�vM�����q�$���Y���f)�c�q���v-𺘃�w؞����o���E������B��I8�����C~�,Fxö&em6�uևb�*^�Lۙv�h;A��h�# T%��ﰴ�tz��i�s.�m)�X��咶�Ut�> ����uwq�v�3A@����-2�������=5�i�v���,�h;��+�S�UKs�������q~��Ͽ5���[�����=?[-�|��24��]��׵n�/�)���3����=�A��|,�qOzL�	�ܨ��{o�g���y��ˡǎ� }��y����E��������f�	볩�u��m�'s�SP'WL�Q���C�3��gJ�' �>�U�"z*�Cu����r(�4�D�[q���%��:�z����Y���͛<W<�X��L�Ԃ�lmm7\wU�l���Vn3'�a5�-r����MC-�c��HB��Xń`K�hc#�@��H�`̶KTZ��B+`�R9� ��]����~ϱ���d+&!sv�l�j�G�.%fL�i��^�l����5hhM9�:n�r�a�ަiI泚�!�>6���ӹ\����<����w�/x�.�}{�m�m\��%h>�{�Y�z�(�b����1k��ams��/��+*L,����ƻ.���P�}畫�W��}��2w���{�����^g��y���o���	�f��v20Eh�;4f�׳U�{��^����b�ބ
�C����qڛ��쮵:mL.�����\��l�Q�pT��5��!s(�[D�jRt�����j�9���1������9x�؜�l��N�|'|>#|x��i��ا��:}Rk�����˓#���+���U��m�Ry�wL��ʮ�xR�zW�^Z����_:7�H,�2T	��{�9H��i���ʛ��N��ܶ������p���غ�Eּ��|����ܭ�]��30�����.]`�LV�Y7����U�sxu�o��k���|���][K���#����]���}E���|����[��:{��UqbI��|��"4/��߷Is�+Le��7��	��>F6���oRA��//����w�[��.eI��!���΋1Wc� g(�D��y���c���#ݝHw���|�Һc� ڛ֠�p����A���>��U��=Ӆ��O��_��h4~J��n����Pw|�V������7�:o�묺�]F�F�O��|8����]���"�e�ܶ�]g���yS\�.1c�\{s�ǽs�����}���)�}���C����gԊ�N�̣��}�����F.y�ǉ�IT>��a��UA~�~�]��\�t��TOxS��*������!�B�w���ot3^m,���@�2���#v�gu8FV���e�r$�G��.��I,��~q����������5�c�r�̗RO�-��	�ڧ�|4�{Ff�W����P��ٛ�]�G�~����d�U��g-�=��=q*��«�z�X׺�ڥ	���lɀ�U�v@�}k.-�v�<�)�s4s׋�VF��=�< <=�{�m]���;ّ!�d슜�i�g��9է��2��z�)V\����O��U=u���x�r���)��YT�7�������#xgy��'/�I3�>�fT�΀q�&'cS�m��ҳ�_�a����e}��G�U����<͏���hl�gV*c�?]{�����V�0D��#1s J�gV��'����n�\7ŤI�Բ�ڸ�];Tv�N�(�D����q/�d�N���9���쿝hĻ��x�D	�}8�Ͱ�Z�	w���WW�>CI�8����� ˜�3���5{�}���8D�5�X�\�MMp��Q�#��,b���rKXӂ4��|��|:q��܁����ƻu9�:�̑�!������h9��|����tSOj~K]Cr{��܆_vr����� ^Y̬���Q��;���X3,�ٓ���a�FnlC�q�6��U��<y�qR�^����� ��|��K�spx��<�j.axe�9����=[�!�n�I�Z��o���T�ή�%�=_?{�/2��}���y�f7�|լ8��}���ki�,�k��dz����ߎ�� ���,V��X��A`�	Ad�)E�{���9����nkUs"�n��s����P�)����b4{��)6�݇5Pf����ب��aJ��T��.��:�g�&��&���U�H��<����t�4�%����T�v𘽧O���Vz]�iIVo�;H׽Uy�r~b|n����|~廧(c9-��遗�W���Y������2���o�U^���/^9�*E����Z�Lth!=9=��j�uJ�K���W�9�6.�D��'����A��Qs�'�/ۤe�E���o*���فP�Ø�6�n�c���h�y?� {[����bg7qhI��_W�-���e}�p{�}�Ȯҷ�L��ԥv�����]R|[��5�./� ӱ܁;������;��A��iӮp-Ai�&m�PO�_s-�2�4H� �	RR �Da UbB��X�
_ws����K殞y�s\�f8+4s���x'q�E ��,��-+|�ú�)llC��y��-��壠��v��3��8�[S;����ª��,^=�j������@�P9}Jm���:�Y��De6��Nz�������?���c�Js_�*m��ܘ��z�i���>�_��=�T펚�9��7k�*�{�9���/3�6�{S�w�J�{�
2ɔ���rkX�S�/:�J�l�|��ܼ׮����@��K�gX��y;%�g8ܫ�f�_���U,����j{���B��3Q@�F��ra�O�d<Y�2�m��3�Ň)��ʟ��]b����Emn�u�{�ɴx�s*eK�P�������AG6�_���X�1�k&"����4L��!�v�I�������y��,(QYC��Ou�TK����dg06��]�"��)ȯ^�vS�ZeqI�dq��\M9Wب��ۦ�<�R�j�ڣ����2�I9C�f����P�ICP|:�N�z�Ѻ�u��i�a��}���U��=PX���|=�׮@ UW��){ʭr�� >N$�4sՄGz�i���u��W?�PoI`��QϱY82�C�H5�cz�UΫޯ}Ͼ�CH�}��|$��q}�I��+�$X͈-A�}�<4�ּ`�N|x�i�ϧ�&3@�1�7;�G��N,s��^�t�X�ٚ�U[��cT����v��@���.������<����I$�d=�{ݾ��V/�#{�y�<8'�τ��L�_3�Ir�۽I�F�u=���g�{n�R�������S������ϛ��8��]�:��J�Ms~��+��q�u�Mh��� X��HQѬ�3���T�������]*�Mj�����5�+����N��=��Z=�e��L��/*
�*]n���nnR'���]�ݘ�r����mS�{��9�k�{�e߯b��{�Є�w�>��1��у���K�:kEV�
NWLI��9��0���8=C��Y�9Ǫ:7n.���'��q���=(3�}Y�87��}������ }��dwumH�Բ�Lv��f�{I��;�+nel<[V�٠H��}�VG޵>��k��vS��{��wN_tn\���+8<\�f"gl)�^5�#Q-%)�d7���e�|7��'���2�ک	-�ߗݗ��4G�zn��v%^�}g�5(���}���2�`�;5�5�R�۔>�0��Z�xXs����w�7˟h,�/K/��U�d� �A`� �W<�z��wқ���9u���وr;w�8�v�3�;!t���2�a���Ǡ����jN:L�al6��4\r�IBڣo�1^�Gڧp��e+�����|MCw�#��>����~Fl�_T�e�t>�2�m��֓��#�wg��w��TUN/Hڋ�[�So/�ڽ��C�����7W�y�S�zc.�K�
�xɒ�k/t���j笑�Q��F���iU].���"��������H��ӧ0Я^�W�"�:�����L޹p���
�gA�u��^�Q��5�l�������\~  ��1e>���)��t9����v8 ;�G�JSn��A�,s1��L���X�:�٦�2��e�*���OR�����@:���9��r��V������A�?�R4�a��i��o�>\�N��ns5�ַ޷�'�$ ��� $��?� ?��HBO��HB��C$��!$����	T�$P	"������& 5���� $��?�$ ��o�� !$����?������@I'������������`2�U|� ή@�0v�v`�'�n�_�LK.����xѶ�קl꫚ڼ�z�[(h��X��ɶ�W��vg�8I~c.wc���t�!]{V��X�{�����ɗj�v���&=�=���<��M%<���4�h`70
0�I�c��nB���̈́�i�%�W�b��p�SMk�7�B�6��_��U�'lU��*6��4��7�kYͣ�,ظ�1<Q	v0$�� \�nUӸԀ�j�R�Ѱ@��{iģJ��k�bj@%1ݻ̧�[���c�E��jb�k򖭵��?�	H��@�I 2H �"BI	�l�I Y�I 	$ `�$��$������$ ���g���} BI?ꟼ?����АI�M�y $�� $����H	$��� $��_���}����$ ��=$ ��~��������O�$ ��}�����;�?���	 !$���p?��o>$ ��RԐI=k��d�MgjfL��~�A@���@ ܟ}������{V���h	��Jپ�-1,���
�QD%Kvr�� ����,�BZĂC@m,#V֚�ꀕN�%���PT�a٭��� �*E	PIJ��H��PDT��v�!��R��!A*`j�2*eH���5R�P�nƅ���qJ���YYjH�-�"�e6c[5LMT����`�M �i54!*��eS]sl+�Ͱm�kS5�f����������S�vҊ���f��U�Mt��2��-�BR����(�     k     N  ;�Z��ݻ��=]��v�;s��u�s[����o7�/k�{olۜ�6�{�����f���=�e���{����w���w��e�w����w�zzu������6ڌ���Vm4UR��JIR��ۮu�:kP����v���ۺz��owM���͛���S�]2�5�����n�t���{w�www3wsǜ{^�;�{7���so[j���=ײ��{z�����W��n�;76�U��Ҫ�[KUHu�t=��u�p�=<{�ۯ;ۯM���x�S�zr��ǽ]�z�j:m^�w��m���޹�*��JOm��o&�2˽��];�/cPޯV�J���۵����e-�1*T��w �Um���ɽ��f�k{����{���k�n�׬�#���:W^�oCޮ�����8�Z��]�Q��u�7:��[l��JX���]h�Q-���NV�{<w����k���'��t�^�i��vu�r�����p�֛a����=�]�vG�����ӧ���Wm����k�׻�zKh��D�I6{j.�-����V����V�a���t+]�cr�wnxy��*�<<y�ڐ�����;��:vw��ڼ{��^�ס΍׶׵��{�l���oL�������-��OW^�T:M�Vu�h�t÷Z���Qe�]��z3�e�T0��wv�{y]�Υ�t��q۝���k�������=�=��oz�׮�ۻ�x
�ֆ��TR���]��&ۗL���w.yu���uz��S�{Nna��]�-��gw��m��v��G�:w�s�-y�o\�5N��ֽ�{������w{��{��n��S���n���i��jٚJ]Ѷ�l)�s+�N���v��Gw����kK��^�v׳�hJ��{]�����]��V�ꚶMoa���"
�l��y{ݵ@a��{W���=�r�������zT�` "m ʕH � EO�0�R�F   �� ��T0 & T�T�aC#b*?�2ez�4  4�����I�#Md�I��2���;ZЊ�ln�Ɣ�G%�*(X# y*���ܶB��8��{��� ""�� D@���" ~� ��@"DB��� ""?� D@��d"DG ������_�H~�7M��W�C[��EBF�bbn�Y���c۳u����4A�Ri�pК�:s�o1�w@�cO�9���m�59�v&�� ��W�$m�Wt��%������)�R���m�����R:���9J�\�;���e�XELR�"���=a�B�2��G]�1÷Y��t �~<N�Z���#G����+����TnR)�Յ�̻�$�����v�ԼF����悼܈uݩ}|��N�F��Q(�G�w�tb�U���@��iFv�媢�1�B����P劒���j��٦4В rQ�тAH(��@P���b�csK��h��'��WK���b%���x��X��ttYIPAA]�Þ4z�ˬ��ĹH�\�]��ͧV�[-��G6�e��Ʋ��Q5ur�0H�,X�� 0Qq�w!l�bQH�y�M���/3�+���&�]�݉72p&����2�k���~q�i����͊Y3����*Vڵ�ܲ��f��Il�w*����7h��˵[sJ���Lܖˉe��r��-JPW�,ɇ/y7T�3��J�K���Z�K�;��0�uMoU�j���KE "]���m�C����=�b��+0�� ��oq�c�2nWE��f�n8��������}�U��Wi$k*`�|�8�����[*;߱V"����
�+�ʆ��2V����X���
���ݹ��QG;�󵜱j�i�O�L��D�[w�t�{���Su�DR���췹#F�i��5�}V�8�Z�,�5.����e0#�A�eb�nB���;��v�*m��]�je�����\�K:�[Q��Z&$���U3��WAMтte��[$��U
�`FPox�J��е�n� 1�.�t�;oD�,t4��˔1�^ٻ�Z�q j�$�PT�)5�bܡw%���mZb�H!#f�P�vua8Aw)�nn��q��]	Й�$�+ۭ��g- �����w-�WD�2�"m�Z�+A.��u�B\ PYA�v�2�2�+p��N�y��lmXy-2�5���z5�ͬ�-�:Hf���&��F�*�.d*��f�٧-�2q��r�=B�����*&E�*<7#�5{�A��Y��Ua�*�iT�ˇ����'S�EQe�ۄ��H^�Do��x/?]G:Ѻ�v� VlCoM:Էr�m�i��`B1R���l��O,k�y�������$5v70�2� 	�nh"F:�
�݇���k%Y��D�8�D޽�_���
d��:�J����Jp��t�a<s�N	Vܽ���^ҋ�]_r$���xAj<-	�܄��8#25-� V� m"�M'� �-��Pf@�WvK�������!��[�*�=�7l��UǊe�F'Ie�:y�vX���j%���9�wWJ���;�pR���$�B!��P%�:����������S�F�@"Y�A�uB�w�7RӐ,�b@��m�2Mɋ�k]����l�(*B]�`�+ �ձRR
�%(��"I�d�	����Vɧ:������yܻg(�!mms���(B^�
�,�9lCu���i�E<Q
��(�ˆ� ��N��%z�u`�)��x�Oڬ"ι��L;���*Ƶa����eѾ�����"�c
�v�R.4k��a]�N�@�f�2i(�f[wa��z^�Vv��;R����bU)���3[�J�����ܥ*eػ���:���
�t�U�^m�U�V@��N`�Ih��K��ų��֚�b, Dlm-OL�p̭;��m����J��.��X�1��j�ꡎn�b�_��C`�vց[�]$��vЊov_sW�;/��e�<� ��t&DZ��qf,�n�0���)��FÍQg��9�4ف����%RiT�ɤ��� ��)u�S��K&����I#L�Հ�h�b��0���U���(�6�^c^�-T��0�+Y�B�%p=��%7P�|te��/��`����[�.���*��%�ƣ
n02�Ej2:��Tj��G���:��2;�leᰮ�f^�`	1�F �	�0�` A0 ��@D� I�@b�H�� q�8��]N��ڮҞv9rl1�k���������� W�*6��ɼ�Ps�mt1_+`��}�$Z����0Btpx��� ƕ弙k't�ݣ�@:�Y/]%��{bJ�vee�90�.�I1܏��ն�+�v�����n�cAu������wK�y9�:=���g%���٨U�\���,�ĥk:�z�����n$�L�3 �5rs��*��k�q�b���e�Έl��ov8݋��(�H&�si<�*ӷ�)��*�[P���3'*���4��lI�;Rq8M�q��8��p��F�,[�P�Bm�U��i++3)�g
��r����aL�qv�Ƭ���s��Y{���a� �ᗅh���e�9(�GV�n�
�Be!VΪܧ��Jh1ٙ��oZ��J���F�D���r*1�Fްy!�,�`���v�Z�ۻ��*�Po�������]]���i̺4 �Ǡ*��nKj�'���76��J���MC�e�<���(ef��Z�6�H?��aʘ���D����"�IV,z^�"77+,ٛ�-���@�F1FcZl�nѧ�b�p�a2�%����C�e�U`&�1�4�5�
��Ac���w��=�鎵'9 �sA h3���N�]�MKQ��.
AP�D��H^���2)�R5�����D��X΀��V�~��5�N�±�(����n�̄d�+q�zPl8�^)c5�٤]�h�e���*X�)��,BtB8tkm�m��Yxp1�li�L��8%���HEwWx57Sw#z‵&XP��kn��㸝el�&`��q,m�V"亐��u.v
�Ɠ�$�`�B�(P��Eb7�[j˭��.�I�h����5-)��Ԯ��D�;z�*a`$v��j�Vl�#j�X�������1X'IW$��B�Z������N�9�d�D�<,@2� h[s-�{�[� `��m1��̰Mj�)�֥��CYb�5F�cùV^�5{����۬*P�E<�̎*n��@�Y�d`�n�s$����q2j۽��u ube��r�b��j�G���ݙ��y�D����mn�6�[([��PL���m�˦���G�.�E�&tRt��6ѹY(�tۆ~{�]�׭YT�ze���s#�[{W`U���4��;%�)a��9�b��y�4�Q�V�4,�)$5Ib��[t��[�i�	P�$�א�CFX�	��֖y�Ӵ!{� OB�6؛[SD�{��k!���y�cP��q<4Z�@�����P�܃C��S�f[��j�j�I�����T����h����f��%1���;�C�T��b�B��j=*r�����Ìf�ܻ��~�SQ�mk.���"�*�)W�]	l`�۹A*m��.���i�EA��[@�D�l�1�iT"ZJ�Tqb�P�dhW���;ɥj0�٬l-�؋.�k8z�ֹ1�c� if꘍"��Di�v��ǑӡL�֖[GnȢv[M���Xb���E�Z���An�ƚ���̬�|j��dfj��"#Q�
(F���n�fD�ܶ�.Ѝ������YZ]�!Go0�'
��Uf�J�X��U����Ǫ6���Cq�X��HŌm�Bb齅9X	Go&��	�)d�IrQ̔�C�Tg�m�M�X��)*�5���j��S)�$���\Y�b�wmI�c��[�d�T`VE�M�X`el�&�+
�,�����:�nZ�).�@PE
���4�h��lnV����L�јԣ���/
�D	�����5��5w�쉚(kr��W��_����n8�j����)ڕ�
����V.�ĞL��`��:�D�y��c92�`?��҄�tP��Č	Z�j�w6�`�A��6Hn$=˳&���j����Q�'�I�<뢨I{y��E�q��Z�����gj��1ޙ�sQ��V6�n6��cx���Z�0$t*�1ցK2�� ��5�!Y[�*z�ae�h��3H�x,;�"V���d��^uRv]A�-��2�F�v�j3z򔧋0JX,<ñ�j��a���Ɇث���������N)�4H.�1�Ŷ�1�z��gc�� J(�1ʃ5�bnfnkf��)k��q���u�6��8s2D����ѧ��+��	۫��;C�e�кR�қA�N�d9m�2fT1G.��r�c�CU	�H���;�Y)*�A�{�,�����K+N���4�r-J.-�Y����
�&�dM2��J��m�W*�d��uO1ע�n�Ab�"��J�{�;2^SY�up���7���y]]�]���b8��uvˍg�3�H]m���Џ��aUtgb�bZM)��IHr{$�D�MT�!⻍X0$��Pd`c�Z�d�c�:ۻ�v��YםF��{c(n��3ef+��s�g��*�����l�k�Uw�>�3�fZ���oo�5�d@��<:[����	��}nXw����]��|����<��������{ @�9�$ɋ#mE��#%F I'���%<*���T�yG���+y�e���Z/ݽ�4(�ĄR���k�V�*�f9�9���j�c���sh��>��
f��\w,��ڡՕ�u���p�YTh\�t�]��K�(�wQx�GNM�V�Yl�$�m �a����$�&t�D^i0K�M���o¶&oY����z�ɭDt�>�Bv�h^ԗl3sn��ܚ�]2`F�����
��|v:��u��f�t�d�(UI42�l')�{tE[�Z4qi"�������#S7w��ʠ/moፗ���� �륏[�:)�%". �nՉ��R���8Ƭ�4�ѳy�r7+R�!m��0@����R�n�]<���7du���H~�5TFe[܍��i%���r�I�&�j��2wa�bn�u��+�Q��ȟ��J��&^ґQ'Hl�ҎSnp�MYǪ�-V���y@��ݹd���Z)[��
pևP�I�{�z���m�a��w$M�J�7e�෌�0Q�Zɗ�)�,��c����\]�1��h� "]�ڐu٬i��%�֙����@�t���O/1쟡����EĀ9+*� ��hm���p��p���9:I���{�.�o.����w��ۥ�ki��S�ٔ�bL&�l=�#��d!*�CtK7�n�Xɔ���p(�m�z ��KL\��-�r��0mĖ���[[����Y����5��P�B��56��e3)�
����X*)C�b�C5~�)Qsrҥy�(AY�z�q~�*	M�/6��k^�����<�+4Gj�&1��DC��H����y����i]���9Mkj��X�v����x���4Ί�)mX��G+i�[X,�n��J'�f?����~�n��ǹ�E��}B�#D~Ʒ�tiP��q�]J�w�4�[�H�]e�����$��q�b �b3�ٙD�dtѦ��&��N�g�Z�p�-�X��*�e�[�������P1��v�k��y1�p5�x�rR�EH?�,�L@�;F����KsR�B��οΞ���֪ 1�4�ؖ�*�
��lZ�n�2P/a��y�k���re�[���r�B�1���f�5b���!5 ���L���3W��J�P4�Ur�T�Z rୢə���
2�m�z�ʚxv�j��Q�L*�LW���*��3*��0��Y�  �%e� K��@���~3Uk�X�)�� �# \�),e����੨�v���nc�SC����4�S�	[��rWE��c@��h��S8�.��
 �LQ�W�e4�Z8w3\Um���PU�m����xENQʻ�A��vm"_G���P��i
�yam,��L�H�z�Y��\�ܺx��ּm�ej�~��H$�SC+4[���V�Y����;cWdZ��[b�pܕ�;�sE�d� ����LaZ�����j�5���wn�(B����t8�4ɔ`E��UA�Sw�ZS�=�*`�A�eT�cw�k�u�2wS+�FwA�e�$�2�r��kZ6��4��3o.=���~Z���!�&;霝P�n���*DE�6�n/ly������+�ǘOdҪ㙕m�HD�#0KOeاLt�cډ ���nc���ek86�x,�����,b�ِ�;OY��oPI��$��#o
�n򐎲�݈m%�L�5�v����VEe(�m���P�%1��M���b�r����\��[�hx��(_���"J�OԮF�-頞�럱hs�%�Z��`��zE`�15)��-ռou�;����V����S��#I!���*#,H�Ɗ�����3wM��tjY��W��9ݒ�R��fU���z�ɶ���h&�j�.���lSn�a(/Ɠ9J�%�I�! �%�@̺x��,���F�З`b�,��t�4!�84;��Q�R���Z�Խ�RLIZ���V���d���Ղ��Q�Zh躀�i�.���N�$ b��p�fֻ��Z�OMժRɈS�.�)�i�DJm�l@���뫓��
�٠��ˢ�F`	�o03r�f���s6XXh�-f���ۧ@l�@���5v�6Z��X�jo҃a�sI���B����Ũ!���sy��LZx���!�2TӶ3�S�EYe#��]T��p��X6w�[�Q�[�{k�����ʺgY��p#(TY�"���w��d��!S�v4ep�":�g��u��/-���e�qI8JqIH$�S�:�UZݗ��v^!|p����ݏX.z�m�^<�:7$o����7�F�H�I�$}$�N��$���7�H�I�#}$o����7�F�H�I�$}$������I'I#�$o������7�H�I�#}$o����7�F��7�y�I#��wr\z�.L�bK�K�N���%K�����h��8Q��Κ�4�r�9���r��kt�S]�j�4�_(�H�U�Ӯ�Ww9W\���XD�wuI'Jl��ݥ̽�aH�Sr(������,ln��!l6ۃ�S�[��IsE.��N�:�����h0�v�v7cwg33&D����kt��@'��{F�5�I�+��"���
��[p����Ё�.�H���i.;�T����W�NჂ��u<��ڮ�z�����d^��Kv"��|��.�u�I̼P��*��gwLe��K9F^�����I�鹬�Ε/���y־J�K�ז薻w#޽S]s��|���0�	mƴި�P]ܻ1�����:K��c���i�zvq�n���`I�ٮ��B�R�vގO^����K��ԲѸŽ����)�*ŗ�z�Wj���������Պ�\z@���"a�Joto�i;q^�L�0�:v/I;��]ԇWn����Y{�wZ�~ݴ� <y��C��e�$�t�Y*�ކ6�5+O)[
��x�%;�|0m�g��{�9;wAot�t��}����`��_e1���\��i+иř�l���������ޫ��57vQZ��s[\���&����ѩ�k3u-���H�ǲ����\�0�N��sǲ�a֟6�0�3,�b�1;���<1�ɋ�l��%;�̉ޥ���	�wfG2@�7ŝY��!t���:�[36n��w&뜨��@����%��T������gi�6��`ʢ�ș��Y�]�ܜ�18r��d	�Fő����Lt��v��SA�����
�2:J���f����v郍oG·f��{�p]}}�ݫec_�����5bW5����$B��[W4;)�1�& �;L�����������o�%w}���>Wg�a+�yDaկ*u����׼!�qA|�E�s�G#i\�F��Чs�k ��zk�ѥ��b�n�p�핂�J�:��a`��In��TD}�y�N���c��JN���b`�<�R�F��J�����J���70'�.E�tFѻ��麩�C��Q���f
����ab �G^:����Xx،:��=�S�a�t�]�G1!5��q��zj.�{��ϱ�W�� ���K�mE�@���2��v��{E ����q�n��"��I��1S/��fj���-gWTL�#���v0l�'$Z��m�n!�u'�{r�l.��H��-��t�[xܑR����]:�{�1
}�_! 6�㴸P��3����ɩ��h�486�qZ��(�>��G�q�J9� �s�S{)K�l�O2Κ�*��$�O8p�#y��/z󙫝��-2�R.�+:���5d�Q��ŷ �۷��H�/��Ӧ��R���,�Q�M����f+�}��V5���1�5�땣�uL����:��P�.Ma��ay�P�f�L62������A]s9ݐ�!��6D�t:ق��t�zl���t��$��&�CY;R͙���s�3i:LMnc�̾����k���l5ʴwf�V�w4�W��b�ؤ��s�ӴTJ�k��f�tBOj.�E�);RW;�zMm�q��n뗦V���+B�X�=@��݇1`�C���]���^wq{%�M'�:j����\�B\���n�S¶���d�]Y��Ν�dU0d�Yw����Ŷ�����,�g.oB��9�Vb�ڳr���,��M��y���ٖ�u]���v�]�Oئ�ω:*�f��ݳ��D�BD	�oG,�O�6E�B�Q1^���<8t�;T8j<K0��˹8���o�O�-�Er'YOZ�{��D�5w5
��KOe�X8c��sDM���v�$�^޵���i I��ו\����{�R�Il�2պ�(c�Wd��O.�9�$��ft=�9�z�
Q��q�è���zN�����!p�bpnݥ��}�ܙ����Nu�Х�;�A����3�P���^�45��i�7]bA�"��=(HνW�5�n�S�oE�{y-U5vovbI�7���4Ѷ�<�]�̶��ԩM�+��l6�/g~�y/vs��Hٹ*^��z֍ט�������e�C!�Γ�8XX-[����W��"�f���1�be�ȅ�N�|{�k�k�r���-���q�~r|�Z2[����3(`'VU���*+�f��$!f�$J���og2q�c1�ӹΥ�&y�N g>h#������)۫�����$|�H <�1�hf����:�p�e������1`n
ZX�c�i�ܗW�$�V�;���h��
Y�:�u�Y9P�4�و��h��R����%e������LAr#헔���K���֟d�%Pv�g)u��{k��8у���c\��J=���n��`��U��Ĉʛc�<����t�J�_1Xq쬱���]B��\	y]4���fX�K5�H_Rӝڸ��wI��✅�)8��f�����q�p@/�79I0��c@��;�S�r�t@z�Q�W���c1V��󋕔���o2#�2�;E��ɩ�+�qE����"C�z��,8�&���6��QӀ�շ�X�鉖�Yzm�i�V�^�����X�ʜ�Ž����%��E����긂�ojS7xyDu>���Uȡ|�Gn*��{���/PK.�;]�`ރԗ^!-��F�ܞ ۽�M<J�J��r��]�����4�S�6mȶD�eZ\�e��ƶ��<�2X;G1�.d�M}������_���3ի[yo�)Zu�������� ؠ����8w\�صI���g��T�B��O7Ʊ���@b�;�%���#����C�� �
��9�>�r��J�@����wu��e�T1k*���3e�V�pf-AᆐW�:�A8^[�I\�醺r�I��կ1J�Z��]jK�{�*��J�����Ҽ���P,�Np�)�汜�9��9��u�q�r�C���ؗ�s�w�)�W�c�	�9]�&�s�!6����*�(\�s��4>B���ձا/X����u+j�&d�)��A�/nLo4���)%
k����5�Ɓ�O�t(]�۸����mp��m	�;k��0�w[��C�2���&p�C�]��(�����6���3��Y�:��ui"F�8*Ҕ�n&���N�X��{R�[�wvCܪ��/O��A�rp�ǠZx!��ܣ֙�|l�M���igw���{7��ϵf�Nw"���ӵG����a�	i����1N� l�Dt�)��%�7c���Γx~���c�cm�ٔ�B�o�uܩ�	M���8��v�ܷۢ��L�W	� ;;t�v�`މ��/Xj��X���y�WQ�*��ӿZj��X�\��+��.���1F���%6�1B���7�S:��lk��T��r�6�
v
����=�L�^m"�y��=	�Cen�Ѷ��
ч���R�cGeJy�Hخ��c�p`��s7��=��CWw���:���t��� ���5֢3\��{!�#��@z����H�Ƹ�-��� ����ηf�=�Yx�����bݙi�ٔv	F�����]J���?�eu�Vi�-�+@;3�G�Ĺ�M�F:]i]-��)رXE�kq�t�:0X���|z�)����Sې�$N<Eq��� /:��'
��]�ە���#���b�W�x�Ь{*v.Z⦲ۙ�oS;�GR\�����ݗ��)p��v�;��9�{_p�h���kd���	�Z�.�a��z����b�;k�<������gJ&u-�]ͬ�Y�V��Yz��*Qn9��{w�4fY3Ot�6�Q�hM�uz�kYG��GZ>x��%>��S�z�5�'Ij�&,v�D���p�d�A��md���!]�C�xS��˵%�5]F5��D,���hPꍪ�<�9�������`��V�Wꏘ���aLѝZ�M�GY��م_h�C��i�����>1kdX۫1�z;��tJx^탠��u�*PV�.�>޻��� S�=;��6��B�/�zt�a��K*�����xK�[��3���0Ha��=���Ջu�y�2����7�@@t\u�es���͋5%��Y�&{��TQ׏��-Bf��b�ss��	B�Ae�\�`��PNI`�i�W�u���F�+t��-�2!eI��m��GY�-��>�\�)�|A���H��{�R��K�O�)��աr$ �r���FL(�ѡ�:���l�j<)ʚ9-Mǯlr�� �KOt�C�����a����n�Ӣ-�
7ͳ���,�Vy�_ou� ���(�jLk�o�C�8 Dwqھ�f��v�|��R\��O�̱�O~���r����	<��B��Hx��P��'�z�n>�t�y�����8o��kD�W��.�E�n٫}4�s�S��[)�h���ke�#�xN��)g!W%#4r9�6���%���qC"�xv���iw���k�tA�R�쮇k���QL�՟��wSꔉ�F���js�Gpf��頞)����/X�j�wSw(�U��������4�7O�ʠ�M���A
�8u�MP�^d�[M.�6'v<s���ɛ����iӰ�:��LG	W#�d �Ӻ��	LVd�m(�im�W�yW\Y�Ů�!C�twQZ�����s4jS����]�Xh��-VN[�ֺX��-��y���t�Y~,^צ�ű/-��v�f�ٻV�#�t�M�uv_hG\���;y�������u�`�u�
ӱ�B����<G)b|�sشD�g
c����M�5�TF�XI'o0��d������8;:�� ⚴��ɵx��Uv�r�')^��8D)#�P:���X��7��/�i 1�Թ��'`ɚ7NJRs70��WV#ɫ2^g��Y��܍�[��p�98V0C�rh	��v�H�C9�r��m���֗8��������X�ύp|8�n'Ճ�8ä� ���J�s8���T�31���oL+`')֝4M����UvQ%Z@W�że�lvA�����pen���M��&�B�o	�������x����G��F�&�7�M�2�76ϯ+�'w^��A0���^⦦���onlj�'\�
�S��-5�e�SC	:1��`����P���/�Ve��͸�I�]����ܽ`�yz��n��7���].b����r�,�yA\����D�mqZln$��uv�h7��5� ����#��eAڃG��]��J�o��qQW
�gVRdP2�
�N�89��p^��N��
/�/�9�ȽJ��!ue'۝�⩻��J`��u:V������t����u�a=ǟ ����Z��$�To����ug\�a�,��2��;<S�α"t�\�����%��T#���ힾ�W�3
D�%j�V�.ɼ�h�m��=��8�A�JZrV�!sAN��]�PivwHEZ*�]���!�5����=�wFl޷m��,*fR��훪���L!s\Ե2�i�o-��5��*��ō��g�����i�
1[�l�4U���4㭈�z��ȶf�gH��%�}�=ԇ��P�a!�ѳ����8
���:G��<�r����5ht�S�S��j�Wt�![kt\�̘.n�kU%�ԋ�|�4���{���B`|�"J%��S+���r�1K*��N~X1ƞԮ,��VW
�&��Y#�]o-��f�t����!\�B�M�L����/C�Y����;��9�L�������m�A��soL�v�gcT"�J������ed��l׳�mj'��S�	gz���Ɗ�lp��k!ƙ[��2�	:�$-�����wS��J�������m������̍�Gm�6d�R�o7(����&��a�Z�v��P/hx�q: �@���j7*�5��2�	�1
��uN�ʆ��V/i���w1��[[S��!D�T`�0�!�:�m
R3�w[Jy�����-���ؐ�̫Ҟ��jI��.n��llam�\rtl�a���W�vz#(!쭸���4�YY��������;{ӝ��I����GV!�8��{C�g4L�X�sm-��PQX*��3Y"�	�����0�Ԯ�*�*Ċ7N/���Z���+��jeNm�ѵ�v�E�g�L��І��q��5�.�\��}�]9&�y`�]F�	�L�Z.�{VGen*���[��ִz�?a�I��ӯ[�B�
֑ʠ�_<(<�kb<�Y-�8��ʖ�S�(~��r��P�v�Y	�e]��:�Ӧ�ZZ���^����'P��F�D��{�km��M�X���[�,juVe^ WS�,ۡ�[j�v�Y�eH��Y��1;�khu��w^vky�Y9�MO)q:�BI�<��=�]� ��j��Gs+!���ۍ]��mE�>�;B�0p���r���w	��eoI�����m�,��m��9��m�oI����T�aܷ�p��Il��q�W���# aŹI\�˲��:+��G����M�}�CI���p�ɖge_�4�ŉ�c�S��醪��.�s웸�v	�grW�`�R����]��N����סj���v�Fay8�IȂw��Kt`� �5)�N�=�,	2�c>u��2�!�.��c�fV�:蚏�f�-�*D﯅����ql�f�<NQ#JQ���E3�Yz{�jբ��肫/H�S�n|4G���
�vFu�NV�̝��%"�l^�th�}÷��6��wI{{s���j�.�ې(J!�R-m���^��1d�� ���K�VH}z�̝�[�qh�܋�#آ�R�=���KP&�ǚڼ竨�!����r2�ƻA��w��W��lh�qC;�Ų�S넑np޵Q�3F�;�R#�n#V��MW��4�|���ϻ�7c�����n+��@""?DD@"",� #� ��?ш�1  %���w�ƕ���?�#m���!�����$��Dy9�Gu�2��ַ�2�H��6i��x���_Ksa}��Ԡ���l��;{r���O�9/T5��d��{OQ�}��,k�ONX��f]�I��ʴ��S��	�fFs����E2R|*���m�
Y8�`�8k�o5�n�c�v�%����#�2Â���,���å>���L�ۦ);C��`S�{���������o�2�$b��:�]N[�p2E�`�¯GuCd�"$��Փ����\m����K�0E=�#&{G[�䚜������#�b��s�f���˄�7��%] 0��;������Nc��y�X(��TH��Zy��7�6^r�Wba�#rI�~�)�8��wEʼ���:9�+��:�by����m.���[v��!��ri�T9�Ų)�tҝW7s-���1�+gY�g�W��UƖ�w>�9hĪn���Z�z�DB��rh�X7��V��_[���� �P��hOk'5�w<����5�E�Uj����Ib��ĝ�R�a�m����nm=V����Q��L��'(�*�y�?w-Z����/�������<v�)����
�Ւ�Sֳh�#���7��e���n,���o�`�&wR�d���V�{CX��4^[�*l�o�wf�Ad./^�T���哹(��,X��  �����?wЀ��˚(�RǼ�t��b_ZAJ��/6\
l;�vup�&p�*��7;���^�Ī��4�!������t�?��p`їk�<yo:�2�ɝu8e��Sev����.�v�%m{�����]��@:�;90)����X� aݖX�4�&�p=�냓W~�����nO#����~;�������8UkHk��6Ն4g����~~���e��LҡōZc#���$6ǧ�Y#���)������6�'&o��T�4%�6A�	R�#���Ȇ��M�C���� 6|�w�#H�����u�'Z�1��A]��&4&��acv�MW)�/<�C,��Pͱ��F���RWw���hWֳ|+T�\]�����͹�\/1V�<�Fl���Y�x8�q/��b i!�yƕQQT�ԎM�hxm�{�}-?�X"� �3oO�a�P�u�̯Gk��6�Iٹ}��F�����o��r������zv���Z�Gw�AO����*�}{oN�׭eO*�=`���C� ��@��� ��;�`2�b�՜"�J��H�&�YsV�.�/6Vё$HB � �I#�� �F���M	�g*�rIꃭ�1��#:��cYA�:*X�+9�N���V�N����|l��g_F:���V1�(~�|�r��ڤ��[�"O���N�c5�M�Q��K�Q�
g���a��@^���e�x�rB�LJ3<���%�����]�/��{=Q��
��NH�>�5�  G%�� b"��s�ک�w	�u�����*�)Я5 � �%�{�wv1��7����x���#��s:F�1�b�<����}����Y�R�J��sȽE�X�<�xo�7k�T��4�1қ+��e�w�x=/ǹS&�&R��H��"�ݰ�i�*g�e2�.�A��8;��]�s��s|�g���p�nT]����"�G~��vm��;rm
�g]=�c�������w!M�����y�˺v��;t���L���<9,��v��*����H�E��� %;�ݔL��ol܋�հP���ة
�ْ�0l���j�ۤ�t��[ws���W�O�lAu=kҨ��,I�k���'
�1� �,0H��F3��@Y�kjX��
�i'&	�R3�:Tx ��/��O-�j��="	��.T"L^"b�rt*�T�bP�s�T�kw��Qe7 ����ti����Ǹ�=4�OeA(on��vf<�]V��6�w��I��\ҖK����j�8�{��,鰨���y+���<�o��c7��$������f�;��I�]{LW�c-��4�p箦i	�i����Z�{��E���J&�s��)t{}[^�썴n�{�o�R/4DƷ\{�D(�v�8�1�z�f�ߴ�tuܛ[��V���X]�D����y��$=ݔ�Q����= ~vg�=3z���5g����U�o�[u$���cĺd����� b�2 y�� qb5{;�hz�P'���Z��3%j�4��
���P�����S��p�HÞ�������e7��˒��C\���,�4�~���򂖛�L1^�1�᳷�L��v��t3M���˃܁Д��_������Z�n��%�f_A!Y���o�Nz���0I
c�0��=@��$G�7^��gr�GP�"_+dgk���Ԑs���8#�y��F�G�~���� [��.[��Z(>@����t�Pm�0F�b�
�Tx$O�����d����y�|�M;ۼs�u�,Tvw!*�1Fqua]Vk��l"y�̺
�|��V�J�����YCLWu{>.U��� ( f��� �R�.��z*�hZ��U�>Я���������Q�'�<�1#J���A�7^WF��'|��n�T*Yq,��$�]y�٣w����A��{�Dv1ʫ/��w�hNt!sx�B�"�.V�ے�e]='�m]��>L�HM�84Z��^���f�h 2"u��]\�d���7��w�#���r�/g �>�7�~zM�B�"������o�Ҙ�(�'����+�X+��M~9UB�~��#k����{oҢ#չ��7xr�s]���A���~�y`�(\��Z�,5��2�2��n����4�z�3�rhd�	'h���� ĸ��.=+V;��*mv$s�|�g�ON�Shu�w�vJ��>=��:�1`�fxdc޺(��}����2�/�G�Y{�IZ�r�w��tϠA؁�����(�֙��=9�z��8��FF��r1�|���5�{�d{���=�3�մ����V�Aۏ�=�\�E��d�.�@"a6[��m��ܳS��ӛ�j_X�h�Yf�5�(�}:Ir��b��R��ݒ���r��d���������g�hxfò�6I�V����u�UN/_�-d���)�#(gV��eP � 5�GK筌�����k��=ih�CM��H�dn3�
 ��j����c�)�n�����s�X:P˚zn|���Ω�j$DGz�E:��#�W�C����2xW�>���[�6k:�:q�{��R��k�H����&}7CֻUJ`I,6 ��U�+t��a/*�7�Ya�DF��p���ݡ��p~=.��_y�ыTj@��٣:������]��W��ZJj{eNT�9~�%\�p���x�T��+�dc�~�}�U��[��z3mW��]��U3����Wt,i/@��.v���v(n�Ųh�qs|�m����#�����J���[u�=5���+BDd 0@�%����[�W�9�]%�D���3;��墛�I�
�U3��f����Z
=����B�Cx�
���=�v)�!´=��o��S�:�.F �oHdf�l�AH0`�� e(���|��aZ>��,��Z��s+��Hj������ 8A( ��0�!�P
 �bp��\��+�p���%���v�\��O/A���buA;�ٺ�,P��dR�]�n${WokJ��o��*$��Yz�x��=(��h������Ӷ�N2�5R�7�᫇E{Pj�˨s@�V����O�.���_��	ּEN�e�j"z��3�M�z�v�9b"1<e٠ 3v��u�#4��2��*��ׅ���������06�߸Wxl	���h�+S�]q��ih���R�"h���voyi�HwNn��V�ǥ^��.����k��S���P������Gu<h[;�Ҙ�8�)�G����:W���坯�+�lDj�%�>�v_^h�?���ƞ5�RS�-&������l�Š�%��*_-,p[�`,����ܩ�Y�=r��Pu��l�K�����f�"^𑴐Bs�����n�߰;d��c��Ay��DW��&���^VE%:T4�x^������\&�h��Ά �R\���^�vDD3�ޒ6{q`��uXY�w�&�{݅�<����Ei�2��G�|&.$�B�;�4k �I��4n��&^���n��v�����,u-�c�1p��	"�'���֌'�:��c4>� �X�8&�x7���7�>�������j�y 愴�׽���\�ΖIe�th�ֆ�H�c��g$�Iۣs��Usy���<MֿDpq���<R��k²��;^/ �M�*�������V�.2�Rf�1]}����;��nX޶6�F���cw'E!&�y���yP���u[����z  �a޳57l�{�%�i �3�m�u�k}wW(�J{ܺ��ۇO��s�*�7�P�T�����o���y*�ȸ`�MZ�'�I�'� �F\ph�Lm�{=�*�#I���J��$Ġ���Y�D"����.���0�ݕ�n�{�i�����I�b_!�q�Î���ќ�� Dq� V�@�zU/Eu*����k?H����J�uƅF����"<khVi�5���0��xj�X�/��Eu���o~&��;�U��c���bG@�I�zy!)
"�^>��qeM'{�v��!�2�_�� ɩ�և�7��/;q�C��9�$�f�N@*�^�y��N�er�f}���۰�]W��,�{�g��i2G�q�	Y&9��!�d!� ���*�t��S�#���26��خ7{�so��8�� 4)b@�:��f��:�N�E:���;�j�-X�]�ވR���o
G7��wς��^���;����)9�ێ�+�b�B�\���ʹ�D�V2��|�0|q�ީ����w�(yg&�F��T Y��t]`��3�"7V=Ӕ���mǌ3�^S]̾79K���?2�� �o�W�2����2X�=����g�������",��^1b��U���T�������*ͣr/[��,�.^ts��.u�#W�Rrc�)�ʹ�ݏ�R��b�&z���R���<rЬ�M�@� �#X���_�^��p�	�-G� ����w�!�<�_�4Wa��������Q~�Ժ#O-�ԡ5��Q��h>���!���o�����5+���E�¤�~�����z()�Y,�xR�4��0N��-���%�u
6���R�A�fw&q_�hu��!Lf(�ʛʾ:U1��� 7"](�&����FZ�!ޝ���<�V�]4�L4�����*d��˄�y,��S�r�h�`��ft��q�o��_#��`�U谔�p 3 ��n�z��cV��L�1ڪgf��17��dJ�1`VռI\���+sq�Q���9gu�ق7s�.0�.�^�v���\]��[8��b�7:+V�]������T����ſ�<��f�t�Vh�G^o0.��X���4�O����/n���8ۦt�Z���4�-Vg,��+y�}5�D[Y�,�I�\��'yMӊ�������/�{�̨v���zD�H��7��S(��?�$~�A������xe\�S�@�.��V\��� ""�GU����ּd�7�C������׫�5�Mڊ!��1��2��ѹkE!m��}X�w��HI�7f��䎋PNK���V�ܚ}2w~�����h3��@d�ǡv<�1r�&�#0�%�{���ã�O��aѢ��L�ϒԱ��~٘�V|�*�nyD?VUr۽��ښ�� �aS!��%Uzpⷐ�ꠑy�Ě ���<�[�2�d{N�<|���'՝Q���Q��{�XW��Յ�@�Hqn�D@�� w<O!�I�%�LU�Uy��-�(�3���̇C�ѡ���B0�������,3w,l/$Ž��(d����A9i��V�J�u�4��tzqN�1z 7*�����l^��‣�,���uvn�:Hw����6oZv+� �	�]���뻛�pa�a[��4����
8Inu=�Ȭ�zđ6��RB�ő<�ʎO�e��ڑ$z|SD���ӀGn)� 9͛��qsr��9hm���j���Fu*CJ�}(=]�� m*�4g�7�g;�ˎ�>m%�gT���"R興-��0>�o�xh��Z;��j����9ӂ��V&�]�o�s��4m�1�j��(���Zj��$���8��<�T���{� Z�4m!��gX��ns��Պ<x^r����9��K��7��`R���Tj@��(g����WQ���gk��>  �j�f�׻�o�J�)�W1@a-[���n^L��k8X2$�>����m��W�h���.!��A�v�Q��=�2�B�V��w�� @�E,#��%gs @DQ�=鈀�Ρ��ޔ��Z�)��y����k��Zw��H�G���zS��P�\'����ȱ��Y�9��#�Ok�C��$`����!Pis���M$,�`D1��+&��ܳ'�\���Z���u̙ǌ�\y.��q��H�Y�!�T`�v0MP ��ڵ�5wU"x '+�!\����6QV�'�6�L�孽��q�qEA�&r��ʑ�&������5H�F�{��H��)ˋ�P�U�YOo��jq�`]r�1�,�cL ��[�2�sCu���{ :L�A �e�e�ĀH���JSU��� ���(r(�C��$�.X(2!�.��r5^�(r�r�wAd"OL����N�sM��J�#VV�[�r��w�S)]`�7�y^����t76�P,m�9��㽭�0p�ͽu�5NWA]-V�WI�
�6_dR ��|�v��歬���`��rmt��(!W����I/������v���2�-Ls ��mRu/�b��cTC�3��.t#�AUĥf��5�x�НY`��d�2�&Vf�Q�� ��N��������^kt��=�%�hfi#1����f�w��bqK�'���MX
V���=Bc�Z�6���`���9�¨M�R��$
�0�M�-2*�����]T�I  1�*�@�I���3p��(eNv���Ѧ�M�l��(��A�l��7-{H	��#2��M����AM��l�14E	%��	Ќ�j�Y�q2^䎬��l��R9*=)�!e�,�:đ�1v�X:�Yn:��변�?ۘ�[0Ӣ�)��t�E]�Gl,�S�p�R$��*u���D\�jh��}EX��q�tH#���z?lB���V�-}�՛��i�zwwI&6�τwg:�q�줵�������Y���y���!C|�e�54k�
��Ыyl�z$Ԥ}�h/���h=@[���]f����z���)�!u�[J�e`2���8�eۀΑus��+�R����؄�F&�X�������* ��G(C:��9W�����p>ռ#{�6�}p��̊�i�:��ۏ���ն�*�d�2My����Ԥ�ٞ򾓪����J�V�uN���X6�;��LV�dU�-��이{`�.lQ7眨��e�ë�T6�2F �!-��-�L�\����@gSO�on]IY���j��z�F�2WwWX��UҜ�0�YĘ����mZL5d���b�l�#���E��]S�_$(0U�6�J��҃9���ν[�N�w�{���زK"��Ȯ���h4�O6�����U���	���8>�K�r��t^��H�4��GRK4��"��T�ǳ��gz�k�3�RP����+�^]�4����!�7��5��	+�,���o���eY�R��Hة�mX�g�TdU�B����ʝ:�U�b�T�C������|3P˃!���3&��zơ�V��젂�ͼ�(mnL��k���]�]�,�v΅��ԫ1�\ �. ���4�t�Z$��-`r��-������&�,eF���an�t�/NS���kIƮ3Y�s/K��۬��b-�I̝��s�����yPஷ�=g���\�|��������|�U�J3����֝����f�F������D��.\݉,��nq[w�9��SU����فD�#H)�@�!"�,�q�#�`2ՠ�H1e����@D�@b|� D���,��B ��3�Ƙ�yŃd �Z@/���7�����H+��0���0DD{D@�#�!&�`I@��rDp� Q��\�@Q�DIf�D}h``�r` ��Q��@�QG��0�Y�1`og�x�}[W�_>�|�5D�0�mDP0�(�I�ޘ���>0c�qh�1�(�`H?�b�� �!��`�1k�Ȏ1DC=���,ƃ�7�Da� "��@��ܰ#r�Y��r��C��G�@ @$G�3��3ɛ1�e��F �bM`#$a��5�T x���"4��&�|C"�ey��ȀH��!&K0��d�5�~���ovs�����r�@�2`h��B Y�ڈ8�Di�0�(�<5@)`q�1{y"(
"7��	0�g�!�d@$| I b $�`��@ � �$� � 	" ���Q�`i����"M F�,��Aw�^�\�P��� � I��c�& $<�] ,�&��Q�1�	d@&�N{��#��	qF�0�D]\����|�HdB1c-E��,�� a�5rk�iZV���Gϩ��A$�b(�0$�F0	H� " ~P$�4b�E���@�&8��+|�"� �>� �@�C �@����B#��@��������d`k�k�Z���7�k��@��fL�t�+P04�1fHG�q�oԈ�-@Q�@3 �>�̘���?�!��#��FH`"���0$��t��@dY�h� M�}�\���w'�o�$Q�F>KL	>r���D��Ř �� Z��f�" F!���"��4X� I�1j����j��i�c�ɘ�i�x�y�d LE�%�$I'+=���ʭNװ��<t�E���`�Ȃ@$
0���H�H*4�	 i�3��Y�b-� /&`��& F"Hv��*@
 ��(�@�D�M�PB<� 1��P���<���K�Q[�RU�*d�2i�c��Dd@�(!�<\��˟g�[����@��2���BҒk-":�����w�lJ�ˉ����wWITU8wA}�|���IwյԛsG&M��#9H^����P"�!���׷b4���R�/�f"L#�
0,��Y��ԀO��"���,���$��##EJ� �0�#�{;n�M=��04��DI@@�0�@v�cD,Q� �. d"(�%"};0#�x�D@���p�F,��׬�������	o�aDQ�&�L#�M`��� 0c�D�@fL@D@$q��$@&0я@���- q�!F!�����J"#�8��� �"9�}�6h�gbsB���f�d�1��0Ȋ # (y" -�#�
 I�!�n��!�,�H�BH�LQ חR@�H�> " 2#��p$��hC��/	�g{M6:�Ux2 (�!�H
0�dG� 'Ƙ�ס�YY����
 ]�t`@���x�I���6U$I�	� fߦ,�2 I@�d#��E�`(��9�y�~~�J M� �P�����Z�2F" !"��Q�DF�,����B�b0�fX��c�H �6D��f.���o�6�^z�x�� �\�Q�����#B0�#�2$��Վ"��2#�����C1�&T�<`qd00�@dB���b ���d� �8� ����р"}>�>ׯmta`Y��(�@$bC����" ��$2<A�F(8�ȁ��h� 0�& &ǔ ɤ#ڢLp��@F4�>ً1B1DA?0�x�1 ��ˈfL
 [6'+�]���@& $E�(���( :y� ��G�@�L@�f#" `n!<�QLe�D|`d�ޫ�`Q�Ŝ#�i� F�_�� 4������5���e����"1�6d���>j	�� a���� ��'L ���I��P(��@f1HY���,���F&~�P���0�|cLI��"=�> �B�
�>_!�C�2��u�̺��ٛzuD:ǳ�a�峆)Y�&d Ds�!��S@]^Pꚗ�ˬ��WM�`����9աZ��.lZ��չQ�*��5y�p#*�u�:�!5(n��	\�	�A��XA�x��8f!n��o;�=���5� q� �1@�F	���f!�4�]��B �!�I��
"	 ���<B:c� @�����DqE�	� #���Rj�Ӯ�����o����"��8�@��(۲��@����G��?diA�0>2 ��8�$x���Q&Ȇa�F�d����F8�"�`>nA x�H�HS[�{�zS���rw|��(��> Wyف�b#� #F�/��(�0LE?�D� ��� D� ��c�dh2D}*Α��a�oLJ#�#6E̖4�t���d���×� ���:���3�mޓ|�4�wzm�CuzJC𬵊���Ng��rߓ22�B��$`����ϛ��n�|�%�
&��;�k�xT�|/mjY�j��弹t����\1GJ�s1E�A1�j����'uw�S8��uo)�<GߗϦ�Dߜ�����~\Xm�-fe��
�[���Ͼ�f�9,>�W�ԥ��'�����(3�t��+:�mN��y��SЌǰ^�셃��$�UGu��w_w$i�r�D�X�$tw>q���t�)��2�4���^�p��EnU�%i^5����K�7.�kT�9d`�h��n��>X� ��E�X��?b��h1�C�Ƕ��qKa��T�s܆�{^�g�YT^����J*W�6ֶ�ǽӎ^r��L�;_���| ���i뗮�/HڐL�VD�h�1�cj~�Aj�#b��*A�xh�Ffl"j�꾛��h�%$��������,3���w�9�r�;˰�!r�وk����Д^�R�ڜ��k�G�B.�´�ĝ�T���J�GG'6o	Ԇm�⑴�]�Z��h��H0hw�"M 4ޤ�;�훹Д��bQ��JbrP#��F ��m��Ֆ�s�T��A�iB��լ��O01�>|���S�KV��K�1���%��"��ˇ7cF�6d���*��8�m�箛Ķ�F/#㶮	��ChV�ݎ����)�{@Ƥ]Gg4}u[����{ݖC^�M���'fw~�eh�R�C�R˝�M�¥�<���������:�����`�l��i�*ZT��VHѿj��C3J�	T�'OJ""'	����  t�ǖoVJ���Q�7��������)oٞFT�/1�֨2��8\ �ɡ+��#L͘��*�fgy��g�I�:��g[���ˠI�.�#=m�n\�?45/����NJ؀ k�A��W2�#~@����.�~���<A�I�ɻSm�P$eT?�Dɐ�t��T-6s�ʏVy����*�����{G'?S3��iDǊ5<��#�ȁV{���͏����>�����Q�?S�7�%F�a��Tᘺ䫻wk���yd׮�w� �>�E{w.����#<���@���	V|����-�HLt��ӿ�"� ��%|�W.�b������������0���ڷa����:<����ݸy�~�
���ȳ;ED9��O�U��q]ef����]+M��w���m�[Yl\Me�V�H��{�=�8#D��8E]9���\>�'7:��>8q�_I�툈��wYcԏ�|����e#V��	�w[s3�(4L=q���Պ�T�fR\d��.��c���iР<M�ɽ���r��
~TV�վ�u>��>�魯t��_  �$�~���8�W�f��:��#�Dq�,�yoju�ee�C�>\ ^����/Y��ʭ���/��V<3����1\��DD�L�B��۪��� ypu��^�� ���"�|$�1�M|��ݮ�#��{�"����5)�~.S���ԢyV5�hx�� ��vү]�3�n�Z�r9�;��M��we����W)�<��,ҏ{�~��tD v]Q���8xJg\�"�Vu�8{{�Dێ	�pT΃�X�j���sFd\C�N�S5�Ưи��x<=��xH[��唪���3k�. ��źgB��pM��� >�M!ؼ���piJ#*:�u@Y�WO�Wxӻ���վ�˓jx���(������Y���u��c�)2��cD��[>2;���&��|(u{� ��u�"3[�vL��R�& �A�H �I�H �$���A �0	�H1� �`�j�mp��d���O��
��UG�t���S�R���jy+F�! � > �&!��,��׹)�+X쳻t:N*s���yԟ*�9 �⁉�9�*Ֆ�fiR�b����~�n%G:s����ԑ���t_���?�.;���b�x�
��Re�憼����(-�o[�0jY�du50�.6�|�{�tb?���UR":�vg��MS3�y�u�/6DYi�1�7��n�f^���	��z�V�uk<A�[P"��(��� �q-�f��*�V:�\c�%�\뺧<(¶� ��X������B�����m.�G�*��)�'�c��N�UP����" �3�D�ey�nD@˱0�y����^��$lA�m�F`t�N̄�:{��}p��Eef��{���T��"g7���WR�b7:�Z]SV����u��$I@���_�3��@DC.����*����>�4[�X<'�������!X���\��/Ҿ�t��G�,:�B>'�����{(��Ȟ�c� �3�|��6�)���_���o�t."�n�r��H�Z
�L����D� ̵�$�Xe�t?u����6�^0���\�xȉ�o|FQbh��Q4Eky>8���D��7��f�k�Gp�Qm�ֵ�i�E�H�������1���&�7������ G�]�y�tʜ<D��y���s�T+�nM�J��fk�L{��Oh���P�\��@�~�\���<:�R��<�5ġ��sE�MA��M��y�˙�X��w�/�@�#��W-F��}���U<�[�Mc�Y�ZfwZ�r�9�D "	��@dC���U�kr�&6�ֻњt���G+p�,�ެ��Tr�tX�{��Go1�=AM�񩝶:��]:�-�&�N�{�[��/kp�Q�$F���q�w��@�
R�|�x�W���u4�%� 5���i�zT�{{<0��!��>�	Vݯh���I(
���X&��!�����ׇ�Ic%K��*�����5=��P��B�,�V�Z��������'c�̠{�:�QF	�0z�:�#5� RӜ��|��lOmm�7�ш�����S������G@b�� @aA���N)~�e5�ǻ嗻��}�S#��[�q�y9/��S�_�_T��y�F��sd�ZJ���6I39��P�AT�*�}0I�v~��a�-)�V_s�և��K�!�N�m��m�79Z��`{�˧��ū\1s����RlK��7'9]�t���x�Xl�&Ӌ�C��]�V�&o���M�;��>�m��|<֏�%���ON���'���9���PL�Q�Su�O�q�Ny[4�
>^)e�z���l���G��WD��zu�*�a~��q�*,כ�.�w(�"�Y>�(|>&)�S���6R���RW�ߵ^�r7ӓ�t��
D��~�!��YN�^��y���c�X����A��w<�r� ��W�=�.��6A��Ǣ�
��!.�s;@�9e��P �A�,gޗ+V2p��o
�5���;%�p.5��9i�}����q�Д\k����U;�V({{s��h�◻d@�㈒�����o�K[B"	���^g�D\�?y��_\�9�?$�ޮ��B���'�}�1��ҋ,�\.H@bnʉI�Q�t�a]*@��\�}i
�^ii��|0�ޭy�u��47	�G�gJ4" � @���j�7� �z|��g����f`��R�A�Ԍ��?%����Ϟ��B��:<��i!I�ˮ���� �����1���k�J�8l�<s>?K<�}Y�g�}�u7��x���j��Tzq�:��jE��/���C�1%D���t�����i6=�Ľܒ�ή�>���=�D�<��q5�hk�I!�́ɭvp��2���ZO�y�T!3�4T`��Ս{y%@{%�D���%���;Z"�z5Z��!9����`��$�&���3���_DG�M9�+�5ޯF��ί�
4��h�zK�R����gdOQK�_����w�#���� ���n~tCl���>�^����+u2i���R�;
]ҽpt���t��$ ,������e��ϫ��RO��0DD���Nޘ���;usdF���?��K|���I)������ i� �G��S-�O�	��%�\����! @[,'b�ڠ�~�XЬ��]}X��l�&�5q�J�2V�D�v�Vv�����XS
���Y���^��M��%���m�/'H��u˖)����+�����6!�DfucZ���}�.|�2O{�K ���J��>�S�rP�!UGP>F�4o?[�ݒ��g>��,�#w?b����S�'{R��D�vr��c�mx9�d&��\!��6GMt��X������H��j�J�+7W7��CR���J���W��aG���cb<.oU$g�z���0���
b h\�������?m�<��c7�S1��:]�R�o��"�ڼ0�dVo�c
m|'ڲ��$:�-;�q��MڟHH�x��jύJ����~i!dLR���t�4�mr��)��|}}U�#tf[ �䝍Lu��K��a@�@#c  ��)���Vf"�}2������Zɴ���S�V���PL�6x�{@.at�]ʡ.R��{�q'���@@LA�S�up�U��>Z	 J.��}�/��\���&�?{}����ځ��\�"ޝ:���Ǵ�ކJ";�HG��̵�ѨO�إ�et��n���wޡ ����A�#s���e�AKu�#bjw���vY����/��6G�6�M��%���"nj�ż���t/*�.�Fϼ��Q�}9D=���q?'��5g��n�z&Q��[_y����}���IF
"�)�"$/��U�zi PT��9�7v�Tq������v��%� ��@FԂD��(�A�@�m1�!��$83a��W�E�1<Su��)喚�Y���j��sv&��K��=r�gI�P�z���s��ZC�ݱ�u���.mp �0�M�������]�� Qb"��ު�0=ґƭ��5�����eg hm��w6bd�jWO���d'�w{�,2 .=hL�L��A@��T�O���T�u]
R$DC�H����N��D9g7*f��y�Ճ���!�nG��:]���vy���䇛#�/�A�����/�xK��;�m߅Ľ������׶G�""��*���B�,�Z��Y�_R�"�lUw�<�g�(�I�j�৕ڪ���r�gC��Am�v�� FJ�<��D@���&9hy^�m���(��ڨ���GR4e_k��h<��k�y�'�6G�s
SG�d0g��|�X5��$��S��䒽G�S$t��ػHo�9�3��J�@D����A9�f�
ZU��4���wE#u�C��]F��6�	O�31P)��A��^����l��N����S��0�������+
9��K�gm����)|q�:���ػ���SͿ!����{ai������u�g��
��S�:��B=M+-e��a�h¥����fx,��ޜ�����O���*�x����83�`%+�3�X���Z�<��)��O1�=���������I/>怟�S���xR���X1A1�dI	��ž~�λEK�7O���*�<�4�pI�uHб�3���l�D����9�C��[lTf�u�lw�g1�� ��+��j(��XBh��]N�pU$���A��	�n�85X���cMN��2��l^�-1��b��ӆ�E `x@�+�J�i�l��;Tx�'�;Q �|Ĕ�֙�2t�$�F$�!���	2E*2Y��c����"*P
I H*�l���u)$D"P^���B(i�/������g8do0G)w����:sK8gX1w<�㌍ֶs8���x1�,�Wg2ƌ��۩/_m�`k%�5���r������b�y�����/%=���5|���P>�Q�[�B#�0{&�m��+�X!�l��R5�kM�R��&��n�m�{�-<���ZT�����b��//�y)A�f����f���:T�$q p���GTԛ���u��h�Ǘ��g��d��R��윈�h����nId��R�xe�к=�2����;Qu�n��T8�U �#�l񈠇e���wUY�O�*Re:��mbV���DU�e
��M��̺�`+��] �b��픡\���G3��b��W�f�����X�2dK��f&0��d[��x7��0n���xT�p�<�������
��n+H�A�<m�����s��Rm�9�#��QR.�9��לp��G�Vry��g0]p��G{��X-���
բ�j_]���1Wݑ�Z��4X��A��r��X}{=7�U��=;�F��$��$<��vP�{kdg,��r<�
X�i�<�j���K�hb|���Y#w�FG��wt�,��qWfPȻ�S������1޳]���"�93���z���[�C9<�s��f.FQ�X[@��(3db���-���ދ�̢T�?zzŋ��ҕnufК����d�NuаF�ya�z���0����/h��Q����]I�#�7�+��J���ef�=�.��b���t�.�S�F��Dr���#�]]p�:C9���p)d�����Oi�6e�+cȎ	yqTM��m�o;���������EA��9�3kw����q�J��]rmm����ɐ�v]=8|�x�u��`r]d�+J/3a&��|f��q(W+x�!n�_6�on�l0OeH<ޣW��97y��]�B�+�Wa�B�P�}�t6�;^2�eY���I�e�Շ0�iU�2�����n�i*Vĭ�Wɒ%e�Zbq�.ΏCUs7w���nƿ|6da�T��:��8�&f�����(��
�t<�ml�j�(�݈"��V��]�,� �i2MPZ:�g���-�<=R�_�4w.���]�(�FR�ө�l��E��g(�	���wSĸ�<����Sl֌I���طI�zUA}oH��L�7`H%��&gn�ձv��d� �o1	57��$κ��YYyݗ��[\�TO����ɥm�V+b/R�Ȭޛ]So�tܾ7Ȱs��W[}fVK��<�R� �;(V�����ɾ�91M�H� N��j�
�����:�fu�c��صK����[Է �	�����^>�i2�&�O�Ǟs�b�$�+}�,��SM�����.F�����t���рJ�U���eB�7d�N����(Y�����_|3Q�s'a@���4��V�ٞ#�Wխ���ꢖ�D�#>O�U�+3m���p�f;��V��w����~[o�Ӗ���l����%Z͸>0���?x�8�!	���Z��$~�g���g �{ϒ����;1��U��z (��n#1�Pb�I���j�%}ౌ4~�gOe�ڙ>>���T���F\���lc^�����`�l�I�����1Y��.�&�J���BτSpk�-��߽�N�g>�����ڊy3Q(��l��*��Kcu�
8�MLզ�����Myr&�v4$Ev_s��3��CK���ҹ�ͫ	NA^7FG���O�)^�O���1�>�6jY;�����1���� �5W��3o:;�;���Z���z=n#x��^�������
R��)>L1��X�?l�_#�a��]�Q��:fs����^>+�W�K�{3�~n��� v��ܥ�iN��xoQb���Y� ̱��
�`�H0C�! A�I � � ��f�7�v�ŝ�Q[W��������ܬD�h��/A�&$�t�)B�&"	 �I-"A �E~l�A���S�e�Ԓ����Oakv-з���JN��`�������8o6暐��i�m_�G����g#ݗ�9*N:�԰MH/Qג��j9̬Ãչ��$E@��|=�|Q�ńZG����g4�G����})���7�iS|����1^��
p�U���[�h̯y�  �zn�Λ�$�x�Y�������Ee/o�s�D���߶�����¥r�ϙo䲼�D��YPepjIbR�@�:��R��<�dgسV��J�>�����sn>�O  �NG�T��]-L�Ks�(�A����u�kՋ�G	�����~i�����=V�e^�E��Q�k÷l��`x
܋���w�$9V�ڭ�T($�M*�������X�C� g�o�A�"����=�0�4�{��mS���c�Ϗ3�>Rc���O2��0��7&G����Ѕˋ2��z�cy2�_�՞k�`;��h�Ɠ�P!"o��w�bZZA �(� � �`���ut�Od�ym���+]��h'��׏��5�>�]c���5��^�܌X��NK9˛� ��&"f�r0�(	l������i����o���^�R�hc���AM���gz�'�R��=^<]R�gqn޶���F���oȳ}�t9�~j4	���b� Xд�����q�5���1ʌ��&>Ix�U�R@�?+�������o�5���㒋�q�lJ��j�?b��N�Eg���~{��"�;Zgrf�'�L/k��CP��Q�ї�.�.�u,I��G+hj��{X;�%Ů��xUۢv!8��N�<7��
<;w������h����2"װ9d�U$g��Ɔ���䲃�0R'�A����ah]�؏0�l,�Ц6�*�6��O�x�#���B�Ϛ���a8��橺�A	�M��x��}���T{���d���@�CYAW<���oR��MI`�[�J�����1C1R��kؽq��qx��F��e_`��^GD@"7��f�O���"��J�o���F	��ا'ib�	0������OOӚm�o��{}G�I��O�Zh���e^�m���)O������xq8NB��Id��F���f�t�h�C�ӡR�t�F�m��,N�};]rG-�4�7��.��	���}q�"��U�J�����g��9,}��e�D֜Kr�H8 �;1 �����=)����s��=�m�bf��P�4^��r��11�|����\�3/���UeI4Q������fZ���`w�$�6A6b4ē7��3���|�2k�!ޖ�����?3�~��һ�?��d��^/`���&�����T�gJhZ�r�A��(��}��B�����`��3���~��V"�<#�M��]�^d$��HĿ-�cJk����Ԑ7<z��V�#��(�BH6e��P@�ŋ��? }�����*��Ծ��h����<��L_(�3��$'8i�]a��5����Oo���[N�������q�9FN�x�.L&�\�(J|��ӹ��(��wr�)/VE��}��*�v������>��a%G��Lm���˃��f�y�.A���< �D�.)�(o{Ӑ$6�<�bṻ�-r����F�(%S���Ƕ�{f4j��6��!�|8�͏��޶�W�a��4�����R\�����GB��^y��m�����ZPt u��2/�'��'a;�1R�������Rw�dF��L��r��qUJ�S��ȹ
B���_�`�ܯ@֜i/Q��iE;x��v����~/m���y^E�%��Obڨ�>6�������p����t��� �����YJ���>�x�Ա�#��so�N���t�o�h��B��nq�̆�E�Wz��g4&kvL������׮zw5s�v����g�א�z�BѨՔ}Cp.tb�
�X��d5�2���T?L�:WN��Pb2�۝��o�x 0��>���"��V�|�SK���\�@�7t
��:&'&:L9�s�O�%��-1��c����(ރ�����Ú�:v �i��ޞm�v5&�5kW�|yP� �>��岦�o���<�8�	 H4�D�� 	�I�* F �F��Q�?T����o��gޒ�Rډ����k��A�H.( � �E��cZ�<��8`Q�S=k��W�WW	y��_+�w���t�&U�(��p`�btu�#Jc�y}H�ے��c��������^Y)Oi��N6��.���Z�<m��K"47mDb
�F}�����]�E-�/��L��.������K�6,q�ŗz#}5�}���>�q ��Ë�;�.#q&){P�%�Z'�c�)~�nj��v�!h�ӗ�_`�p_rS�l�&ȆM1�=�!X���2ˢh�%x�jY�cC��oy�* �"h�d{d�zŷ7��*]S�@��d9ů����3}��&�FB��g$c��^���\�tl[B�n2y���a���2��mD#{9����oz#�Mk`�î�F%�(皁��/\"�1�������u��yqi�����#�������Ѯ�}k�2�J�S�X��{��[��}�7C�;��v��(�K�ӻ+kҍM�e�M)(�g������K�´ym�P��v��k���i/Vb2ן�k�k�\����sE3�7���D�9�.D�YL�$�[9l ��q���穱y�f>ϴ��^E6qEfly�����o�����A_�.�q;�u�����İ�s�`��s=ǧaK'�|��1�;e��'�cO0N�}�I�=3^�51�p��e#K!$(� ԃ;wrEJ&�Y��7OoL]c�]�?�|��oD�,^�F'��t�@F����X�؃�`�#x�E���(���@8I��@A�� �;tbMc��v��F�ި!΄%H�Fb�}	s�ߐ�S�Ǒ�t�E��p`��1'��䱓}���5��>�+U_'����|2/V�͞5�h�i�����ٌ�',�u ����m ��n�(vrW�{�{В}W�Œ�F�7OW�N�/N;D(��̐����7�0c
�C��i �LY��A&���ߟ�����s�o����i�rOԬ`���2m���`p��ct�=7wmv�N�T��5��X;��f�zO���~�}��]'7+UCfv������k��o��vr�� $m�}��S"��4;�S6�X����_ T�D��O�E��ֲ֗�,�mEe�vh����>Z�HS=���r>kN:�#����E��'2��ȳ^n��'�aY`D�pG�� �m|�w���/1���l�� V.�>$�?g��S�l�y�u�g�U{���4:=U����:�q=����%�Q�%foOi�-P�&�[�K�����~7w��
y7�0��	<�u++/)�HS�0�}k>�n�(%d� �,m�l��+�@���/X�<��R�n�2kT��o;�S�ϙ��㭬�byq:W�ܵƔ�ǎd�駶�3��*�nO4�����9�:�{��ު��܋�F�\Ft�X�Z�U�S�!)�_/9�s(�~`W]��P��k3�m���}����H$L�I @�	�Z�OO�i˰�O��i��>��.�ד����>t����UUi�4����nX;�4�(4C���sp;\�,�q"�Q�Ĩ� ������px5au�b��l�ܫ�<s|s�����F��\�
�1��Іs7��7��0����ћ؁��w��]�b<�M5y1�6#}Ua0�:���ܣ,�y�  R�[���,���1��k�Y7�y��s]��|f�lڀ�+�(�KS#�~x�yJq}�����}����5�����]�Ou�����+����2��=�8W���_����f��8cB�c�/Y�/�C&&q��ɗ��B��s�� ��͑�wӑB�r���d�9��Vug�U�Gv)��uX"L
�}u���ƭo@�L�� ��OM��#h!�0���pt��ѧbY��y���U	&�H�̊�yIE�wW���׸l�,��s�u�Z�X�?+��gh�$Wk7Np�@�yw� @���2Vq����tsn�KE�.��)�e�l������� �	7ʀ�;c�fi�lC{�=�㽊���u��9��.ukf����Ū�_D^weK��˜�4�X�ƌ}|-Ww5t��`���׏-�s{wny�6���F�1�� �.��Ε�i,@�Q���0_� O<ېA��*Ӽ�Wn����rϪf�
� e��ov�[:�Sj��~�ZL����x�A�p�A��)�}��> x������f�	��9V�f�s<Wnؗ&uv*kJvP�M�Ǡ+��+=�y嗸�SϷ�Y�"����ӆ+�`�Hi����%�q i�m(�	*��_bR�X>�e'��;�
ɶ�HO�"m��N����A��B��XZ�I�s/������UL���e�~l��=�0� R�q���އvqib�������^���gOב Xcv�O^��9�1�l��{���?hR�^�?�o���I��������l��[}��oV}O�9��h	0¶��UO ��-%m��A�N��mg��@� �����l�ϟ�����8&��1Q�X���|�����;uޘ�;l�:Gar����M�P��I����,��{M-���}����Q>�TQ���ް�'�φa��gf�Uݣk�~���x��0�\Xq���Tʎ=����l�ɔ�D���B$�IK�E���������)n���=�l���� "T.��ާ��^'B����K�du\���z�]5�|�oefɢ&�X���H��6�c�R���N9cL�(�b�NNU�]�"؂{H����f]s��e1���\~[�\2���ODo37[�zh8��$>��È�o\3��5p�4"�¥lٙ��]�����/�Q/��;�X���5QP�'#��Pñ˼v���K7wB/;R_:��B����D
��\�?|�B�ow��'�2�*�w��gZ�b�}���	
���5���͞p��W���ώxk>�s�۳����*_�^�@����X�B8z�'��:��l �g��4+7�f>Һ�.z�Hy�w`��o�����G�4sf8��6WLuћI�i꘰��٣���+��b#�"}V�?z�G�Rڃ[�A����*�J9l�4`V��30�+���!�j�|����KO�-O�$v^�N��g�:���;+:�!���6�dj�[X��!-A��W�V�|>9����UD;;x��5?��2"_��j��ʃh;4G���y��/�rʞ�v�);��r���n]���Ø���b�&�*ANo��@Q�
m�S����. ,��f�)�e�J��H=nN5c9�r_�}s!��� �����X���C���kr/� �� 5�e�b�P�Vʼ�s�6_iE�1+n q&�0����a@��P�(�ݾ��"-���n�su�z^垩#S����}fb��l
�j��c*��;o�����@#�v�E-�N�F�-@�I�F<AdM��~��ٞ��#��[g�F������,S#ނ?\qW21� �7i��E���+�7�>��w�_w���sҽr����0I0H 	� �RZ��R���\�W�3?M�2���s�)5�]ED݌���v�m�}�z���}%�b�;85Ҫ�	ɓ�/�L��
�㋪b�O��֑�b��!ڙ}�ÿq�D2��U���v�K:�	ز��b� Yn�㐅3h�Χ�-�	�~�JՅ��_[��q�];˝T�9Q!�p�J�vx�=x딳�˞�8�� S�����؈?rV4�5��;z7���U}
���y��=<q�x/�%���U��v4����`4ġ��w�H�4��eZ�kI�Y��z����:<�G9挛"2z���� 0�D=-�y	|�5v�u�g�k2f�ҫ^����bb:DZf�����筱t�a���Ez�y�>b5��Ԧd۬�*X��B�7J@��"���T�mŬb	$�8jf=o�_��=2Qy]nx�� }�7�W,���DHc�*�����s��I��X�@�-�HP1���-��V���c]�;6����Π���^s�T�L��,K��F��ˌ��V �6�UwR�b]��H�-�`��eE'i��u��E�k:��Ù�1����{�l�7Md����Rf�XO��j��*�\��j�2]�S�,���HR����&�ʾ�D�[p����UCb���aM*N�;ȴ�GTIU���5z�H$i3�	��;U(�\��N�7^�֭*����ʖ��M�묹c�Z�h�3zvC���T��p榈p��Iu{��0���y�/�r�H��.��!�ƻ���s�;\CROd������J)�)��a�%�[֨���h[@ �+��ݎ�:g!fsc�$k�c�懓�qX��,�N�e��b�>�M9�{�����l�45�k�bH ��*�=��1�d�@AHX�B�x;�*;�vU&����Yک*��&/qB�E1Bd��w����;+b�j`8�4���J�+h]� Nhtu�@�Hp8�<�cwF�ePD��g����Kl�@*�A����*�b�6��kn3��S8Y�N˄8�_�ZV�e�0��W����oj�O�:�wa�1h��Z" �y$M�7��E��Ÿ5�kb�eҙw��X�ٮ�N%Šƙ��μ�!�Z"O��I��u��1��.�-�j�(3�tw,M��W)���:oEc��H��ihU�K\ܑ��M�pG�W<�IRCd������v){�*�LfS�k�=B���y����}g3=��9�hBV�:�#�Eq1̩ۘ�i�v[�{�]��Y�/:l=���ޕ�rG�aNd���ae���*f�� 7���3���+WW���YC@-����ݳ�/�Qp�:Q�s��׃5;N�0b��X�+���}�9�T�����uyrJV���޸�Ǻ�b��hs��\ڳ��;r�B��G��(/��twO�y�b��6�=��eA4��V��L���t�Y��خ�P��<�pÖ�ШF�bL��{$n�6�A����G�G2�wNO��Yy�S�=�zw[wH�"��%a0��̈��-�ua�y��HCy7[
�8(t��_lK��s��9S]$$�nd�%v��Z�1�VZ�������i��]�f�k4���!}{�K.�_�kY��h��~�'��G�J������V�2����Z9]0I�]�b��U9�Β.��c\�
۫����@aV��ȷ���n<⛗�1Y�Fҩv��u��K����X�����ԅ�7�AH�*�hv+�:��4m�%��XѤj]��.��6v�y��&9Zv�:A%�\z7j&�c&zy��x��p#�e��	�N��"� nj��ۦ���i0wzQ��]��M�Y&�=�7��Cc��NyW��ikx�h�6{��Z��O7�hSu�����ً�vc�Sa�&��h7�ܠT��B�mL+�[�]c�W|5M���YY%�ܷ#�����J+��n^{_�{s��Q��)e5���1�����=J0W,���7_	�#����Psy�m ���S�f#�=�>��B7'^��]���N�}���2�>F_\�g�2i��TPb2\D�`'�� 6�q��G`���M=8=�nN��k�s��z��{���)e��Q_C��qb6h�mW37�j�+2&u�R��n�h�a�QT�x�%���3�b"�����^b���]�����wd���k:��f���D�j�d�D��:����O�z3
kN���7qjц�7���s\&����lY5�\��>  �kGo^��d���ILz��Ǥo�yw�ع�a��8m�4�/N������w�Ӊ�}���X�����7���GH���;�WћGp�yub�Ji<�{��0���*w+Ƌ�l�2����d�a A����<��r�h�J@�7t�W Ʋ�V��{aO>R�l�ڲ�D~7�����S�pB�H��¡����{%��_U:O�h�;S�Q��������:����7�3���)��`��$B$��	"�0����S���f�Ly��n[bw;7'�@""�1�z���.lS4��ȹ�k�i����|w�(��Y_-[���vع��D���;U�͌���@҇R��ȉD�{��+^їÐ6�Noa����4�����f�_ST�0p�Y�ir|��>ܑ8z���@�f�}b���#��Z���/��dd��g���t��|��6���l�t����!�-])��O��]�[���v"�[ױ1��b���G!���oʙ>�Ouذ��u���ߴM�ˈa�M�,����Uܮ�ߙ�-�)r�o*tRO���OX��M�&̐������*��L̴������j,� �>n�|�n��{���d
�V8n����wަ��j؁� ��D��.C��	�\�3X�7+�,O�F�\@�CO���>��17TE|t��;3�3�y�˸�zs�+Zf:d�e�;��M�0�a��+��χY��~��6�@T��=���_O�:�}��:7���˗QՌI�*��V���`�ڵޢ`$� 1�c�E��\�B�t-V�`�@�l�v9q�9G��Q t�|�b�5Pw�J�ˈq��&���Թ��p]f;�0�G��\tc���ό��1��]���R�=�����_OM,�B#�y��N6$˓/ԟ5��G:�w4B� Hn�Z�?xM���RE(�܄UA�\g����kF� ��9b�8�����b�D � �0n��n�չAʽ�l�`ݼ����\5�owJ�/W+::�M���v����%5���D�t���(���w��h�d�ޖy��e m\w�r|��i{x��e!�i���>�=�9yR��5{V @Q�O����i9�Dah(�!t*�"<�r{�Q��T�
��J�xw�(=����=1����:���3Ѫb"z�bkc��5�9�k_��2-*Y�| 7���{޷$�"���9�w+�@gU2@�Tϸ*��ĥ��]'Q������z=&�B	�K���� �X;����/�삶�q[��zw��k��/s7��&$�QZR�V=85S�1���U�����ӼZ���(�P3h�K��l�F�\���Vs�YQ(��uR��u��й��>���NW4sڇ{��o7��%%����]��M���`���ɇy��m��n�~f���kg;
n��r�}�o̎���]EC�˨��O�����6��j"�g<��5�]�FÝ��wic�Lu����>�"� �	& A ��k�}��.ʹ���]�W9��2E�Y<���A�GUZۤ����{�\u�Y�ie���a>�'�?��+>���� �1 W( )���ܪ�ݧ
�ۼ"����O�����R.	��C$ѣC��O�5F�3�F���o	ŝ�/���\7��>�7�+[��������Ik�jpq���%��y>Λ�s��q���ϱ���|�N��;�|D�IZ�,F���{���=��=>��c�a��l�w�jD�Z���h�JuI�k%45v�;�Yud���(���2_�u����j�f���V;eZ���GD��!�`h����
%�wl��43�잍%����54�M횬)�l�<� �E w���]��>X���[�än���@�O��)���p�a��%�`����F`�ùz�|&��$�����]tD����m7U��zc�d���A�
�Q�m(Ҧ2�`M�3�6x̆@����P���\)���Y�F�"[d���U��|[����rBdc�ٸ��eH��gs�ݖ�*"F�uӀ�Ěc��d)����:%�����U��,A�����`�0H-�R��R�n;i*۬���n���ʒo�Y�26#ʹ�QqN����㘇wx�!E&��m���3β�ǈ`�IoB��e���g|f�iҞ��#v"*:�=�����씟H2ə�y&��P3=�߆YO��|l�D2h�0���i���R�_h��x�p�;ʾ涋��RF�|X�$���l��bE	�W��Ң�`٣o��`�fꍽŒ���W��:.��؀�5�:�5�`;��r���ҩYR�jV�{]0	�[�F`�f���d['��ےEc=W��Ƿ�l�;A���M�9�Ф��L|�  >�Oݻ[�j���c7Jd<�q8��`�ٶs�̀�C�4�Pg��g�Z�ߴ�L��.L��7��8��������O=�e��09Č�&��5a��
m��f����������{��V�f�{�㑎z!ǩl)�"�sT x�>ѐ���1k}�^�o0�6X%ꥑ5�
���mʍ!l/���� ���E���U-0!�`@����'0�3۴Ł�|Ћ�{�-²��׈�v�g�/n���C�$V%����z�oJ��Ƹ�s&l|�������në\�u���^\�i쫃$�!�� .'���Ժ���Z�2/W	�?5z��d_2�k�K���bąMƋ��[���	�I ��pb�y�}2�%��\p��>�|c����9m�f�y����bҷD�,<��&��O�s�et<�L���x�u)z�Fb�^aU�u۷��<���~������/����J�Y�y^}~���|�q(�` ��ʼ* � � �0 @@��o�j��>K����J�i����׮s�gX�ˠ  �0� "2��h�3����4_s�����S���Wa��������IxVSU�V��s|mXԹ�4��ky���>�zNv���-p:��.�:py�ϫ砌���O}ˣ>��x�nCb���W#���*��$�ɱLN�x�\KDt��r� ���Ea���d���|z/�U�?`��!�`� 'NcL�;�a�<�~�ܜ����Ga�m
/{�������� �#�o��/ۑ(�8Ш��'���� ��VVځڢ�E���0a�ӭ�5�e�q������|��EH��nY�^ҩwg�z��jqsnk��O��o.�J�~�dj�#<"#����>��U�5U�kba�X��.�D��os��]�|-��#t�F���gvgx�:��I��Q���oN�韼����j�s���γo�EYL���!%~pG/(:����qD�`p�y\���pdɺ�؉k�v�k�����Y���%�뗼�1.E�CD݌�gV���w�쌇9l�=+�w|�E�������d����4�_����n����y���J|s����R�M�b�bM�Է1�{�Cט���v^D��>2lA�4d�S��K���ޕ��p[��q���7P'��F��}�f2`|�B��s�"���c�]-*�Z���z�\gl���4�ݛ�ڔ#k:���S)�n�7F4��m9K���3��#�@�9�i�+�ҷ}�	�a�q��C)�`M�ʗ#�y�#��4�x�՛�(���v��}a��'�n�?K�Ր��;z� QR��7���q��_��A]3�����0��u^�ר�R%�P���u�+��qz S��@��V2�I��3c�6:p����>�~�G(���f/���Qޮ;� ��^YSU�sJ^&�����M��k��.�-�c�a�/�}�}Oh������y�X�'�_�d�_v���{o}�}l޷v��I�nq��#��:��MH��tJzl�9+�^5�xL\��緤�1���|j��WƑ���&#��ѕ�X���tR{t�dz>຿{� (̹��^er�m���m��0���/��Ƌ7��d�F��?q_���J˰���S{{�˨��l2�x�uή�$f5�e�wfy���P*o���Cڛ�#�v& �����4�]?00�^7��q��(���_;t��}�h:()��X�KH��_N��^^Wx�e<u��Þ��������mx��nM��M��AF��@d��Db<gD/�:�Es#KF��>i�gP� #	"jd��0-���V�r}��V�@N�[�ǆ�$��:,�ߴ
�:���[b��ۜ��tŢ[a���x�ʹ���ᓅ�tu³�9�㓃����O���J����ۻ��R�{G�{\���)��C���q�|�۴�dϛ��^�<��y�Yʷcb.�KзTu�T���YlfՍ̧�,o�u�h=��Z��۟�]o�le�F� e�����c��J�����׾ur��,�N��8'�9fA��!<�Kv�;��mcl��}r7�Z�b���ǰ��|b�@� _(�D�>�~��(�YO��^�Z��}�w�^*wK��U��	��v�\!^��Wӱ��:����lJ��΄�E�9L�Ƀ][���XG����wk+��7-#zo���ƨ
�n榷�B��'ķ��毣:��X�08r5Եaӆ�7SV}M%ߤ�t��C^�k��{�5��1<�Ӗ<��tv�K�<�����bw/vĐ�.-*}9��4ƕ�\�hF��D�dD�$��~m��H&"�ӆ��H����DL���X �q؞N[ŻMu޴�i<�2�p�aH$��$�L8 �@ �(��U:�����C�D	BZW�xL�(Hz���ݪ��m��PSoP!��v�q$ue��=��*>"��ͶKW̺E-:j�^g5�͙w��[��M�\~� f{������];�߻���I��0[Ȳ},R���"��UN���;s`=�O5+%Zg�Coq �7�y�m����r���E�b�������w-l��}����=���K�7{a
wit������[�W2��&z���[����cT�
��9��;�+�����>�dީ&k�Ve035��u8.��2i;���e�Wi�Ɇ�|��>��JoZU��[U/�!�o��6��K9|���6V�O�X`D?n�U��FĞ�\���-0ov��{���f�Ԍờ=jC&�^��W����Ʒ(��?l� ��!�"�+����޾��3{��(�W�2���U.�o!�pU�Nr�R�����[�z�U�*�gb,a<��{������zt�U���UU�����@���0�4�-�= f��`�k�{%y�oE[]������z���>� " �!5�R��F��>�~��t����U����"��PGb(�0D[@F�HT�׳X݋S�yư�n�DQ�+4��Uׁ���Cgm�*X<e@����ײ�u�n��s��ŁՄ]a��I�Ӕ�a}�?^e���c�A�{�)��d���6g�z~�i����?���t�s[�-��dl���ȊN���O?*�d�7�ׅf���Z�\\�5<k���l��G,)+�<�-��Z4X�ɼO��~���cf%�ڽ΢zl�L|��:�p>|y]�O��4��09��m���;�):�[�;[����=����ڳXW}��'@r���N*��};�|�߯�޼5��n����zKZ/��=3q��>]��ζB"g8��k~�EC�5ޭ^ �OzD��jg�č~�</hkw�s����۞}�g�jVf�����5����o۾��&�]�/n�0�D��[~^���柸B赲����e� ��8�M��u��xy���f_�����k�Rw��M7~M��=,�M뵇n�'M�3<L�P{�1�f���rZK�m�x{�s[�"gw\KQ�f�r�f�5�vP���7�2��)��趤�O�"��T]��A����U�]�Ƅ�A7�l ���3F���X��O+.�ʶ�T)����I)L+D	��[wܲ�7�ZL�L�R�+����nh�;�v�2J6��35���M����H$`�,,2�(�aM�͙��|Y$�l���E�5���L�q�}�x��ܫR�=�����Iw՗I�<�%��{g'V:��P�����m+tyP��8�m%Xݱ�4޶.�/�(�aC3;SWA�8E���n�C��̵����-]�L��\��q痥ʑ��h����Mv6�ȡ�xue.�w����C�p[Y2�OE!Ln�倻��Q�QF�Kt�P��G)�Lj4�f)�s0R<�S�i^m�B�MK@��c�q�/@����1k�,���2��f�{��5YrR�+��y�l�^L��tb�f��98� 1��ff4�}c�Lۑ%��	3 i� ^����$2��3�19M���:�R�fc	��Z����B�n:FOXx�-I�$`�aD�9�;�B��T�*˘}���o��u��#��I)�H�A�ZM�C:��=�V�,fv�]y�d��nR��S+>�R�@�鱒гln>.w#���qGk$�22C�WMu�Uu��|u�[Y�"p�{Jف�7UgD
���j�	�ԣ������|����m���ɯT�X�dT
�;��*W6�I�e��ʔ�t1�����g��v�Ԡ���CJ{}1�֍{#6f�ʁ[F�8PY7df�U88=�qHAH7��v�Ѹo#-���l��ٮ����:�m���{�c^,�rcz[�g�vͭD���QO���Ӭ��yԕ�]u���E����nh���Wv���ڤ![l�9�vR�4k�og듙�j
t��9�Q\ښ�o(�5N΄@�:2ե���_F�Q�cĩ9��b����;���u��V�M.y1~����}��(��Wt�N��e�.PԺ���t��r�W`9�Ê�[�]�Ο�l�o7!{��U���J�H7�;�����.˳}S���� i���Ξg#}�Y����ɽqkr�vr�,>��W@���k�xH6���m��u��Jq�y#�J*�:�޼T3����1�꽺�
ۜ�ۧkx�U�z̷"�dO�n_F�*�t��۫��r�%W	�m��r8�P�����T�m�d\6_v�(�k�j�.�)m� � R˲&n�kXmP��¶~�]���DH�Z�9��=��=�nX{�m�XqZ&�3���N������uvG�t�9��Wd޼������r$�k�ct��i�Ml
�t�UN��E̦H��P�Nk�����)���Z�j��	��7(���')p�"�������<椤��n����۩_~�E!B��3C���U�KLI�&�:�N�<vs��f`���B&�ߖ��U���J��I֤��"xu$㬿��U�1Y�fTCꪾ����MRY�+o[,*�WH����#W�*��p��X��dw�A����1���͉�{ �T�ښkU��*qsM�vL>]a�;'9�O^���d	"3e�Yej�eK�u30<_�����PY�_k-�ǭ��c ��l�C�b�VY�~$��j�.�Z�]KqB��S�;&���������zSC~�|����F�f;'_O]�=6��YTdX�p����:�����t2�^�����lWx�W�3l}�\��f�����b^
�b����'�@��{�J����I.�1�+��`�吊�ދ~y �\��nW��ӷw�����C������� �Z��?F�t�d��>;]-~����i��.盘E7Z���&CC�Dj�^���K������`G�9U��%�0Ӕ����i��ǐ�ṙ���WW��La�Li`:?�K�s��,1���H�[���e
�;��7KVݭ��9Y8��"6��5�6�J̓����]o�
W�:����ڼT�3�1Q���}�
�����4�x[�<�sڢh�d�ԯ|�a2���2ߔ�h<'1yv#s|���Yw��|ݠ����,r�O���e�s�M9��������6R7�aUR2%��张���fά�T��۫�#39�F�z�PS��гt^�a�wVxd8ݱO�\���&��������Z��2��&r�Y"�v�gz�&Nk�nT�w�1������(��ͽ��|���ɼ1�%��j7G���>�?|4E;�9&�\d�o�25Z��"|��L�ڽ��m�U�U�c�gA'{T�1[��vXS#��>sg;���,���-t�����h�����9��ifu����&���-�y�/*�ٲ�[u[��=��ʐ�` �`�̘��^�����¯���d�6]Jsb�Θ��1P��tS{���0$@�;�j�CRs�W��s-;���K��-�c��S�[p�C"	��	$Ɨ�y4vgI������� pF8���^��촰.����d�[��G.ζ�ݦ3��6�)֋ʸ��{�{�	���|��z'Cw}�u*�yc.�h퓘�.y�]��3y�Ћ꥽�Kѓ�7U���0�����u�7�@�>^��L}��22���y,ȗ�
������
�'�/���E��E�47�7��Z:GG�����<B{���@�q��ʔu2L�Ku̳�j��)��=~��:0_?4[z�TC��~���V�y�KS>��?;�o�sF\M�j���0��
M���L�j�,�����.�Ѽ �7�`��MvP��|��l����$ @0{��9�~��8������[i򘌞<�7��w�����ܞ���{�E�'�V+����
��a��2����4i����Ŗf��7�eb|RH��Rz}*�i���J�
�k@�lR1��%�k::7�n�*��� ���J)Z�"-G]F������mؗ$@d�#�d�	�0:]��K-]����.��e�ܲ+gHw1j���7Pp�l��7&�NGfc��gm����W�b�Wp�;��d.��J��vw�M���ص�7t�E�;�!�\_orS������]�Om
&�/F�X-'1��2���aE<��P��WXsz���ӳ��^N�n�d�3�_�J�Ү2Enn�W�r�@���Rn�}�����]��zJPx��b�_<�=�����_� G��D ���C�K�c���i��R�lg���'��%��_v�'lUp����M��#��5�
�����U��v���9��܃Į9���;#),k��h�1sv[w�n�Nf�d��RS���/���9?zn�t��U=��7�]6�A���2{6>>-�k>���L����w����)Z��:�#hK�E���ղwk6ac?Q3������Յ�@���[5ʅ�Ɋ���b�z#�6���]f����_v=>R�{9������>v�@������W�����*�*��$^��6e���d��p:�Q�$Ϻ4{�ˮ�>��4��A ��n0 EM>���E
�p%�#����x)%�7���P�F"� ZSIA����]��zQѕ����C�vI��:�na�}�ǲ?4nu�8O��'T5Ju����h^'ݯe��ʜ�7Yޜ�$�܈��u�7�c;��n3������q�@�w{�e�4(�G=����Evck�,�r���[!��/�w+%��q�HLS�ɛLvyi��g�תĩ��ج^�.<"��|^��b�>y&�=GWQ��U�2�tѷo���;�<�&��_��%�\Y��;ڱ�`+63&�����+�
 "���utn��,zX�Bu{8\���������n��u��EnwHǪ�ou.�L��k����d�=��@��W:<4A!�[�I�MЙ��ɕ�c�����8n{+��w�(������R�9�£�0�7 ��m��ޡs�\�ޠ��iڮ%ζ�n���{�٩G��F�͠�ZO�8���R��5֯6J�Ì�֟�Ǩ�D��b���R�V�e=�v������1P4Ɂk.|�qh�01k��x�($�N������ꀔ�l{��U���$h�`���"�dCcC@�h�3B��[t��������$ `�D�͈��{o��q�`/-��I#j,jN���Q\�R�EWEp���7gff7���{��J*��-� Ih�Уbz�Um7Jw��r&�4#f��!!����XY�l{��a�\�t�cD<
�T�n��S<?1�3[[t>W�T`Z&�t���a}UD?�����p>}�?WK��!��qT@�oX Y�H��3��>[�s��2Y	�'5�OF�"���+�K�g�DQл1V�ĳV<Jc_�es������˷����2��
�)Ï��!"�`�k*x.�ʘ��/���_��-=n�r5��
׹�T�����@P��6[���3&�GC�����G;���>����⻺(�T���h��y�jV'�y*N#����ۛ���U�y��뤹��N���=��c6�;7^�)�D����v뮊�]�����$K�إ��-I�w���1[��*��8�h�-�9�޶�����!^��Ay����$+���%훠�w[
E'2fl�n��fmWI�E4�H�p$A�?�ndV�K�Bt�[��а�6{N�˝ۦ������ժ����X�HL�[]I@�z���
D:��1�ņ�����^~�־]t�0��4��E��Y��.�h��mG(^cD�Z��>��SbӬ�}���|]Nc���ƫI��v[���4@2ɫcβ�z�r�\��̓u�wE�EN@�vN�뚵||}�U�J��]�(�����=$���5�_=����*1�_�%u��;�˄�w�*��/Ձ�m�|'�rxx������p��o�U�҆f�EH��5:I���l��;{;U�����k2y�VsЎ	O���5v����9Ḥ����9f��k������Q�ܙU4m�UI^�@6oNRq�q� A�v��l����NI�~���D�j����|�r�~�/�V��I�?^���s+�{x�6ms��vgVŕi��3��uLT�����������'�p���6������U����w��]���7E�9��^�(h�vƐ�1��yw֥e즆N���e4S��%p���=�Zs���w�tdPJ��fs���Ix]��9�G�އ��_ �#c+8u}��c83M��k�5Vg7՛�ñ�+-�S��'b4�3�����Φ�ȿI���[�}�� >��#�n"�sї=.s.��f�R;��sL����q�b��kw;>U^O=qnD➵.��`���4�T�E�����w�F�?q� &�7^o���X��T�j��i*_0݊��0�H�I��e��$�9��
�Ƚ8n��׎��s�A�h��ֽvz�u=d��~�R�3B����k�џ10"7���}���]l�Z�f��1$�Fݜ����\�Z��>�00�Y���fW���ݐ4��Y+�C/�"��Qr�̩�,Ly��6Q���fS6��+;Cs��g���4�YXɶ�w�#*���tկz���Y�f�O�G<�J�;؋�����o�'�����5x������ J�<�ĉ�U���!L`uZ�|����|��#M�Z�[�?�Q�
��>�o8{�?�R�3�0�� @�"0vm_e���ldw�"� &�RQ���o�s)��h�~�� �Z����)]����Gn�TL � ��������k6L̬ 9��"��k0\�~�]κ��4�@z��'-|�?���\��ogH;5�����P�9Ǡ��J�z`fظ#EN��ޘ}"�~Ң♯%���@D��2f����{��HU|��}s��?z�Q�D���,.qm������=Ҹ�[qϽC����Oq7�������S�g�(j��F�a D��MB(Lo�Cz#gn^diH�\�6�z�S�t��4�I�.f.��E�h��qdw�X�!�2���#Ӓk��f�&�����^ȍ"(�Fb�kenO�����n�Y�R��^�'t����}sH\V(9���,X�h�<U�J5M2Z��{&�/6�y�82�fdv֑1���*!��g+�Ů��7�{:0vʵ�u�}�lP��CC*��bEڪ�S1���o�w�
}z�(:�=L��Y���	�#0�w��0n}J�3QU����[�u^.KFit��P����Y��`t��p5]<�udG������܊ShbC���n3���)R!)�ģB�f�k���`�֦ ^���/�O����;����UN��y���w�V&4;�n�C[�k�s�k��/&^m����bvg̹/�9Uޠ�+������>+���Qű���׫��|ͽ<ᬄ��|���u&��ؐ�X�\��[e�<�(�+� ��o�����rS���
j��]�8���+��>��:���e;_3r�z\\-������,D�[;�,�~�b�K�yJ���r���*CԾOqk�����3�?j�x���lŬ�!^,��ڿ7q�~���س�����6� ;���z��Υ�S^h/�* I�+3E��9}��e�Dg(��j9��Ꞅƛ���O ^�������XXU&�vl��1�8<�i�)��l �vo�v֧��.�US?����yE��}�`��g�qʅ��y�]F�r�7F]=Y��  /Q@ n��<���d��^�v�f���U�)k��{�Z���|�`����Z)���[�ބI�]^�y��ŵ�$��!�4hF*�L��I�]l�l�ZoAf2�6F\�F:�\�����h]�t�3�q"j��Ŵ�U���1%Jk���M���!�|�AF�[9'a�ӂ򰼛�D����e�.�_rw�w��t1�M����	#s�N�z���0Cw��\�(��T��a,*H�����.K���`ޔ)mv#v�6��p�/������͡����J��{7�k���[�$5���iaq;�U�C�z^��)�7��V�էz�Y� ��I���yDqlg78�G¶�Yr5߂ַF�κ�śQ��+�*�p���#���[�v�rv��FR�Э�p��I��d�uwPKi56�,���r�77xD�f��b��:�IW�����xF�Q�� �nc=\�n���L��
q��܀ㄘnr����:ՁBt]��)W�)��*v��+6�}�T�q8�-A�1�m^R��B�bJ�ͬ]���3�=�'=�t�JQ���X�:
z�8"H\ݩ!����0'U�V�b�Y"�J�U���qQ�-��CL.�]�b ڣ�`6�֏<�jXUN�4h�*�@�#vw)����[N�%����-+u�Y��X�S�;�+�Z��F����$�I20�^v�a�8�GP�w׫Cݶ_p��i�:�0��s��� �����h����%��{���Wߞ��M����4�e��Qf黣��c8��o*�s���]��A����(Z�Ӥ���G�3��;�Vôgq�:R�䣱|M��V�0�IΦy�np`mwז����	��_e�����v��An���ɜ�lK��D)�����yQ���g.�Z)Ƽu�дu� �1`C��Ի�|Z�xi��]1��������vI��X����1���.]s�����i�2�cD
d��;����Z��x�\�:���Tmn�I:�����j��HVW[�у3/��2��	�p�4�tRc����k��&�^�	�K�wR�q*H��{�t�M0��Q�a��*Nwwڴ�t�lv�Y�VL����#�*�_�Zj�H��(���f޷�fB�h+:�a�Ѹ$!��S�������`��pѢ�Z�l�48.�:��������V���+j��%V��멖���Z�g.�O�
��Rr᮰���e;2�)��3b�2�d������yԈ�]�ܺ]���w�p@����/�XKcuµ��o3�1,B	� �����1)�	���	�m�p8�f������c��G@��6�(!���?>�ڦ�X*�
�5�/���ʶ���x;X�����;X�����H�j�@��gU.;�{��K�Y�[,���D��t�֖m٘�k9��rX(�ĕ�;lXv�d�IoX�\��ť�͠U.�֒�oo0@4n;���s�4n�-9�����~cy�ki�˭�����7c���u6`W�,ڣ��|M8�n���Uݡ�DP<kY�A�(MF���Fs�RK]���$��}�^4����P�v�����;?M���]X�3�n�o�I�	�y�΅I�3��{� EsS��:���"huJ�*�u�,ޕiZ/c����x���h�k5{($�1=^�ƺW��,���/t�7޹l�q��oLc������rыjcu�v�	�j�ŖL�o�k��n�)�7�ә~
"���/rWt��6&����p�m�Ǖ,ʏv�F��,�K���j:;&�XW�r������6��c�[�Z��&8
����ݛ�+�0@�lq��h�l�)�,��fr!O����P��ϧ �?��&\{�zו��_�n���D���S�vbb8���1x����yX/M*�����_��`�ᖗ}�����7��%���Mx��A���z7�w�R�@�>� z�g��@�@��x�;�៾=֢В��<���j/�9��9]�f��f�
	�(8�rg�:ඳ Vbz�R�C�w��(��%< {�'p��;;���7Ђ���ìJ�V�&@^�#E.�x;�\��w0Kj�����SAT�SC�F�7̞�f��P����3�F�>W{|]�u�;�ҞJ0BꨆT�5?�^�c1�E���8����&"�v�r�.�V�o�����7QYJ=�+8W�ט�ݎ�8�C1�^�ߺw�߹��wl?A�^|-�|�j�sn9@�����E��%{�[�X����ߖ�<X�������:�v3��xg'1�+���C���� _=[���ݘ�ˤ(����g�$�N�"�N�0F�wl�Vt��g�de�6����ݗ����'���ꀛ��l���(ހ4J�yw�B�w;���bQ�����1A���#�U���ć5Ci7�z�t��noc�������g�ҭ�PWD4(|���o^r�yݜ߬��"�7�@�>n�F�{�vkU�̷�B�k�,���{�C6������D��&P��(��m:�O^R-e:�Y�J���^��F��EF��R�>&!b��!$Iڠ�Œ�W�������a�J\�ton��Xv���g�����f�B�A�j�ϧ)�18Ir��=�+G&�inq��@bg��}	�6�^n��V�nz*V�+sY��jA��[���4tka���"K�BսbҢ�]hY���B�^�g�_m�4�]��D;���#�����z�_�}���8S'wB�����,:�{z�{�ػ�l��l�u���D�n�gݷWu����:�H�B���]w�ssx�����p��w�����H��H}�b�[�r�V#F���].���_� }�-y�vS�w�d�^U��b�oy����l:�܀P�s/�q��:�Tc)�;.+re>;��[ښ���HP��+@��D�\��r�%m�k�9܏���^����� `�@��Ա��E&�oa�;X�:َ�}�ϩC�F㧅�m�q���i���,���Y��QXA��b֋u��%�4]x�&p��`��>�=)�T҈�n��I�@�5A2f"	@�(�DIA�U�	<��rA�z*o,��Ys��q��Z������0T"QS(�A �ē("�$L +0ݧ��R������m��T+@�}�!�[Xx�5:;ד���:څ�/o�o��Ӷ�DrW\���k���t����w�^x�����)��3�>GK%�a`��j�������yQH���v�<�����[��[������;�cj^f��ޛ�+tJO��ո��x�9nz�׋1�r>�� q���z�F�UUxv�-��c�&u�N�p����.��S��7B26�`��qɠ;���<���Jf+p��Q�YP�/xw��x��U���u
ګ؝׆�Qfи�u4�{2����G�Φ�}�O��ٷﻥv,&��t�Re�q� q�yY
w��>X>Cv9��gq#�-��M2�]�^sLn�u��w-5��r;�*��ef�c�����T�
��  ,|�M������ܿN�=��g��O���<\ǆL�SĨS����e�w�>�7x�r����,w�7x��a5��hUl�`�&*C8g`��vf�@
������ɱl��nA���)��,V
8�]1�A0҈(�D�� ĤL�]n�T��h�)���gnM�Cf.w
��ȳ�;���1ec8;y��k
bpZ�)ޗn=Ŷ�ni��eJ��\U��Z'�4�B�]s<�~��?>�{��wU��[����H�m���|��̍��3:�v�L9�-9�B��.��G����n-B�Z/�@Ո�\�w7w��C�8l�S�K]�"��w���<ī�EM���]Wq��M\c�E��]��vw�H���8�֭�p�;1Wm�~�t��o,�%�wM��H�����^�7�l��!��b C�p >���
������o�f��Y��{ޭ��}��fR���%�B�=� R`�|~�9fMV�ٗؐ�2F����1ֲ�*j�	{{geT#�廯���}�e�m�E�9�؏"����ߪ�ح��'e��Pv9�4n�Z;�9��r��N#Da���o'h�V�xw������{�ګ���E��l�A�.�Aي�}c��2[owy��\33���9�<��gfd@����"_��V�ɐRYA�ș��@�e����6�c��,zƭF�f���5��ynpo����� �'=4�U�Cx���{�;�ol��
=�d#��-�!��ھ#&�P�f.Uec���w;�}��O�wJ(�����GAK_��բ�^-�v&�m��027קq��'�\�؜ꌍ8�Ֆ�*z%A�.�m��vv����(V��~m�{�4�՟c�
v>V_�l��wv���%�p��v��l��D�q���\�ή�����9>�Y�|�GC�+�s!{�Ǐ3�
X2�3�eT��FF��W���U<�@�ٙd���}��y�W��>G!�����f�������}��z�1槵KR��P�[��|i�J�����K=���c �%le�p6i]�֟���R�r��hB��ӫt��U7���S(/�q�by�]j@�m�v�����B�Z�fs�S�������ˍ�܌���W��<���<�-���sm��5�2Z����8*��Ǻ���WB����ߟ���_��|z�������=O��(ȂA � ��0` R�$D��4pnYD�ɳ��R|�s���"�4d���Fu"�DE$$��c�9&�ܱ�hN�W]���La��ƟRO{��f0�����3~�m&�����nb~�*b�m���Y����s9�={�O%�Ml�r�ixv�o���w4-��u��3�ܗ*w���#���0�}#��#��U�P
ٵ
n(O�ڱ�ݥ�ҚՎy�M߫csf��K���E�1t��I�,���&K~:Dp�F���u��;ux^d{����{�x�_sn�mT-�(��ݞ�S�&���/�5�61�j�n�~|چ-S��;���N���]"k=��/������(�@�z�^���wkL���uD)V3�"6�k�{�3|��.W1��6Xy��K{��R/��:��R�uk-z���.4�"���(�.m�7<��e�X�\O��"'r�1��#��b[�٤����W���w�:?Y�R�RAi��^�]��o��{` �X�>��۽���$�dGN^�_,�-���W=�V��W/�Gԗz�ts�3����������y����I	&�A��"#� 1^�gY��a�mf��.T�M�����LFQQLt�� � z���ͮ}�PKg雊�I
�ܝ�=۳v�+�7�g����y��\�o�IL2�v������>�����,3�}N�����;{�Yx�����
��/=�D����f�}�ܻ\N�+���|&!z��7rEP�zTr��Z}�+]V˙n�ʟ�R����	>��� ��s��SѭQb��M�����NVdf��z�)}*n�D<�
��B�nf���iR��*,�D�h<�e�"c�mm�e�	wn�N��{t�]�����f�7���Ҽ:D��觸���t��� ���x�m�!5��Ӌ��7�+�j�j�z��a�������i'����[=;��gz��Ivw'����u{y<�-�DK�2v�{���qi#:Y�Y�n��?5>�SF%�u��miY��&�	��~ū�S^F��>���{b�׹�ډj�D�|�F4�9�N�Nk�Ӛ�m�,�/����;GZ#9QQ����D±��7����q��E�P�T�bf`��z�O�kf�^5{�s�0�f�*N�K�7ͭR;��@�PF�  �(B0cC���i��Y�]�����5�<
����ܫ�<7�lJS�s3� ��|�y�[�9nw�#ҷ���Γ�j�-6��n�=3�����9�n�R���aX��óB�y�ٌ��@�ΠVp�>���jX�w[��YX����.���_I����<�`��m�F���.)59��E=<�q��/����j	�H˾�[Ks�a�f�5���ć84���W�>w��o�ie ������b�
L����f�ϼ��й�o�am�s�O��q��r��Β��ϋ���/39h�v۔3^c���u�%�S������>�r"!338���` ׫ٞ�9��Ut�s�#�1Q�i\�Et�saf��
��tR����Ħg���,�Y%����JIc�saƴ�Z����͸Ѧh�ܣkm�����4�Ƀ�O��T��s�9��l+�[�����X~��0�έ�����4!`�o�-����3#����4]�ϳ/~��"�1� ޜ�~�&fT�2q<�tN4;�宯U��ޡ�DQ���0R���ff�H٬��+��k��WG\������C;�Y\ԍ�I�k���6�f�$;WV���ŀ���lk���zX�͊�Y�<.�\N�j�5���k�^R�K����u܏r��8=7&}N�To{���}s��괎�wQϥw6��x{��7]U��&�fյ��%Pʿ�q�T�*�d����)��n�OR�X֋�W37��4l<nR/�jgX�.�$���jy��Ksqs��K�޵=��:G��o�[�׾��v�O���J��o�^J���Xsc�;��W��r��>�?a�'���	�W=6����L�� *��hGg]��Z��o��or]ۭ�/b&M �M��p};�Z����vT�'��٬M�M��Jb����̌��=Ό��N�
i��c5��_:��Ur�>��4DC0e�/*5��|l��}�3 �\~W�~��o{�r~��G��l��B�_}���92%Sz<ͧ7e���Lf@ʇ�H��w2��w�ӳD(^�[l3r1�7h��f8 �Nm�.�k(�C)E�b(N��~��к�L���C�5D��d(9N�wM�cw��i�����C+���A��۝r0Q���:��ݍ�*�*�bŶt2q�&(kC1#)����tG�w*��*�˽�Zk��D���#�sJ��ݝ���5I,��w�Z�"����t��%g�\�ʶ�c���Lُ��(�5�=�-�i���5=9I�I;G��b�h�Ϩ�[���巭��m��b��0�ak�;�v�Vh,��/�:{����:�N��4uM�P�Ի��c�:#n���NĢq�mGW�y$�sh��]�H�:����YӨ��'~���߁���ln��@����C`�t4��ތY��X��/q�������v�kl�ܓ�[��:*��s�F�j��S�X<5lD�ܒ`Za8U����{3���0'�CB�r����̙b˂�@P=�iP̑�W-�{X�c$"��Zn���2F�X�0����ek�n��i�GŘmOfL�"�8] 	!0�ŧ񔐤]��x6;g��H�p�H^J�����dw)9f^R(�7�
	U]��B落%D���&c&�B���gv���Gu=+*�	�o~�}ծ�v�+����$��$m��N{�R�A������#�Tǘ��=�����%t�����n��Q�fөg �8��07���(;��o<Ks1��p���=�+���G5��,X�71ά�f�ё��C'�]��Cb�@u�v]s}H�n�c[��J��<�xq��Q���(�V0;��3x�+X���WR{Ӑ���}fm�Jv��s7I�,mhͺ��*��}�fM�F��n�Jj��77X��R��c�;�j\$R���B�0�ylK�-���ܫM[P���ܷ�U݅8~��-�d{*r���8��(76��k�'H@�fT������B4�M��m1׃9��wIT����F��O-UkK�;�ݶ.�Y{���g^�\��x�]9�ћ�j�fzs;F��,h*%��:�j*
�=ٮ�i�9N��^�iN���L0?t`���+��: ���)}���voD������[�Ț�j�#�[�(+x"���kg:J�p��	��Fz/�����9h��r��rv��ۇ+�S��#7��ؔ��UN��;���K�������tn�!d��D�Dvx��53��c�"��Sq��"Fj:3I���RDB÷\�]��8��o�.�F���5����oK�;��$�����7�:�!J�� �U��'?1ƱZ�p9����ґ���:i|.���+q���up�XMIJ]j� 9.Y���'Fr6/�R�՛X9�l�y�%G���`ھ�����K�t��f�79��j�n�N��\34��ِ��9��W,g��;�o&g�~")U���Y)���Y_G�ͭ�3�nl��/%��L�v3���lCk(~/hSL�'������� d�<u�5�����OQv/_Zx�%�*����WlYbW6:!�,�{rs.c#y�ۓ}�ڍ�5��j�����$i�>��@���H�߫����urV_9F�u������~9�Y5N�
���#djt53�ќ㛽���n�n�MC-�N�Nl��\{�@��G2ətڮuZ9�^�f�C_Aӷ�v^�����?uc�+9^�wBr���t��c6˲-+n�,���4Hw�$�ɾ�c���[D�5OEE����|���N�K�F�3�#'��|ko���-۩�Wډ+���������c.u����^V�pg|=a���op���x(U
 BH�2	U�����u����U��dȻ�q]*��z�$�t� I�$ H�{���C4�]S5|FƔ�]�.�q�H�턾�z��z�̘�SJ5j]`k#���ʋj7�B'gf�I�zZ�%�5�������R�i�����aL�iK��9��|��hi
�4v�0H������w"���3�E�;�n=�{>ئt�r�|X���o�{���z��(v�̎bH�Z̠�@��߽��7�{Z��èٗ�ӷY�����uKr��=k�;=in"��2��ױsvnf�����S��p��R}�[`hZ�5��gl�G�Ǚ����������	��e�����>����iP� I]V�`�Ԩݿ�&���`̚|r9�` =r ��<��
��l�iwV5�+�h��ז]�6���n�+�c�j�����/�[T5m������/��Q�$�y��3y�ܛ#� ���w�=���z-������^ֻ�;A��Zz�r:ΧE�[�7�<�+4��r��k��4�i�"P@�/�� D�"D�9yNf���L�����rS{9:�d�=҆ցF	`�H�0� ƃ�ah`�qC0�6��	��.��;yn���p0� k%����n�,��k�K�"o.�ʨ;:�[���R�rm��:u�=����H#X��(���4'ޕ}�s��:�^Qաo]�A���������$��W�	���X����d��ϯ�D ?9����Q�րfj_۽Ք)�����C�k��ʩf`D�E�?��L_�~����f�.�Ƹ�m��X�R�����Q�wɚ ��=Ìv����ي�d�����!��Ͼ}���0G̛B��A��A���Ѱe��m��i���<" ;(�"FZ1˷��x�4+kc=qZ��uݦ/+ua��O5�竼CV%�͓9�o��5m�s����A��9Ee#�����@�5�=[7��<ç����/b��]o��n]��|��63��m�D�^�[����4�
<�=Cz_�c
�B�����W���c�緮!9��t�3g.]o�q�5�������5q��-��`������T�����؂�.�s7X��ۑZ��g���9���gF�0v	�ȳ�$v����:XY�]ӕ��nU�v�nh���*��ӛ��u6I��g���W܈�1�:E���ޭ��+��=��k�����4Up��`�'UΤ2����aP��\�������7�5�5^�����8��Gm2����E�f�M��Xn��s1Ytfyq��*�"z�������@u*�o>�oS���TT���vg��V�[xS�w��v�q�6>�d����]s��#�f�X���n�Yc�o)�9Cnֳ�k��7|{{E�> Do�F��M_Ӹwʴ/nG�s�1���hLe*ݹ�<�؛3���7�l}^��O��OC��O_U|@v��q�H����M�a��du��ھ�x�u�C�Fݪ����.���A�S+ys˹<V��(��8Ov���ص�a�Ck�9#�fs7���y�\�Jj�,T�#��ۯX�z�5�w��LҊ�Iڃ�r�Ż.o�<�s���L��'La�ճ�W��������g(_|�*%��l�Ń8��KB����ʹO��9�e] �*
9in��a����ٟ�� ~3a�Y�rP�;�ܵR�{��VE#.G�[M�G��}�F�ӕ���M�����_A�lPY�E��GK�9����v�!n-�Yw��}����%<�Z��zl�H�8X�ƮR8��=u�z%�K��#wS7�Httj��x����[�Ϣ�磳��g�uެ����s�Y9Oj���b���٫R�� ֭|��Eu�ڌ\ɟ(˳�k��ͭ�>�ׂ��U��u��=>� �D(T�7=��s�j x~ۼlr��	\�{���Y@n�Z�<����E㬼�3	m�>���5�uR4P֝��3gV�Ĩ泚��|gu3j;�'e,�v�|�B�>ߕN[8��F����f���@�fhw2Pv��g�3=yb�K�_W�956���mI�OA����{�͔��=������{�LV4J|��8��wk:�g��E��S|'�>Y�1�O4�K�2��[����7��*���l#u�Ws85�ѳ�*!;f�q��@?L	abA�0��&>H��4��t�u�j�2�o+��3�gR���sϒ�r�W6o`0E�1��N� �$�I	����P�#�

@X�k� -ul�u��x:��M��g�8Vn[T�.�z`����ZS#�
����)�[�IƳB�su{�PQzV�r��w���J'���}�����ݳ�#K�O`��uEj�
�[�]Lt0���Ӄd�gk�$�,j����-�k¿W��)�ڗO;dK�MR��^�V�V�I�<��竤Y��8B9\�Fs�D��g��Ք0D�d�𩃇�"S<�f�ʆ�08���7����~�TX�1Ȓ�ˎ����\�v����������˵�*�y^sϹ�I�J0fY�uJ��k�W	&����39��j��_�C���(�o��X��k�-�u,L��.��Ҕ��z��{	��=tl�>�����a�n�b|�gcRś����bΘXnhv)�l�N$cY~r�ϻ�c�z��y��
�rU���k�T���⠲"6�Os���s�����+���W�8�&������о��G�"�@�5��b���Ct�gf�);��y�yNݘ�0 ��ic$q��ȼ̌�]�K�URzp�K-ot��Y�k5��Nt�u�v�W�̻Jq�s
$����V�������N71ԓT����u&�;����9�wB���x��:'���lm�;��=X˩�K�j�q��.ƪʹR2Ӎ�9k���#� ���4:�c.u1�\�4��v�'���U}�L3��1�<�m}���Μ�E����1k_Vo}4��,��;�3���-�g�Ot�"�c�9����{ڶ�ݕ�6����X�w�7GB�d�9ٵ��B���Nm-������yvｰ31�aEu���B��[�"�Z�����y/�V��}�oi�[�����)o�3�Z�>X��j���I�Ҍ�M���:����|B�-}M6k��OR�Ӵ��d���9��{�O /G���<��ԕORa(�g'm6�|�ə�<�t�^v��S��{c��{��ٽ�j*��M�j�\�W�r�-Cp�#uC �(��1� �����+q�Z�S���1~�&�T%��	����"!&Zʿߊ!���`"G�m� $
�!��$C�L���mH4=�]6�Q����dco�.V�su�1��o��#D��o]v�L��lق�%*ʻ&Y���#�g����{^$��:��{��˲-�q�D�V���A�WN�7��2N��Bh���|'�kA�����v6c�R!-�Ȟ�jH�t?�,Y�&/j�t�ʺ�`���]r�~|Ӭ3�,tlC���\��Fo�GN<���r�O=��d
Y������|��1_V�������v�[{���k��O ��
�rmYY�7�������Uo��Ω���w+7�m��ߢ.e�2�e7���$^d�g����V6u��u�y�)Z�rfY�4C#G�� 
�K���mon�ѝ��gk��~�zz��|�)���;�X"�?b��3���O\�K��qF�TZS����U���E��/��{���#�ֹ��Xע�te
�B�t�y���起���߬�M�Z R� F��DRc&2  �t��t���8�*/�vgqbۼ�Ĵ�V�	 ��D
�t"�l�j�4B"!{��QAggGp��+.Ve�"�#�݂�O�]���\�Gam�#����l�dRsg��i�1�֫�a�|O���������m�T���󡅹�4�r+nDvq��=�gm�����\�ϽeU�,^�H���8c\U#�@�lξ��lh[G{��E۹l�A�������f�,ާ��]�\��P�����ܣ�ݺ-޺�e��}���j6���ټĴ�0ت�}����8&[��/N�x���@0]K&}��z�v���},�Ͼ���P����|�4̪�����(d����S�j1�{�����tޗ���	�2���Q�(�2�T��T�aunc8����W�����9�^�'e���" 3Ô!R�5�.��g�&栺0���7}�;������[��#�1��i���zމ&�{Q�ٙ�y���d����x�bc���k�g��M�їL�;�k>�-��=����u�+ ��+e�fiP��j雷'݂r[�I�c�� ̢�<j���t�	x��\�]���m�-���)�A�]/.�k��x+[������[�}�Q`�ѡ�Aܹ���ݚ�f�#;��|�X}�+P�a}&��E�5���/�2���:�JX�m������ 3S�g��<��ft��R��u��r�;��3����x�͌���]�ު�Z���6n�[��o�K|�1��=p 	� u^y�{ˈ�7��R� ��l:K84����r�f�<��6g���E\y�\p��	���bʻ���52j�1��S2���7z���z���f����t}��4�)z�$����Jω9�yr�oo]���ض��9���^�+������T"OmeF7�$֬UiN��yxf�9�B���*.
Z���B�OZ�������
��bMT<�}��b���t|�t���Y�/r�$�\M�L�a��vRמ-Sc.8�6�s34��g��⬨,�=>��wɮӿ5����xQS�'�md�"�/���4��[X���UO�1�r�uK�8���S����S&"��;4lX�TН��9��,-��	v�r���P���QTg$��W��"@Lͱ�����_Q���)@����8��mY����-c�	�pv
��$�:{�>��bDP2�I6UQ4�	@�`��@�n4!l\��%��ZA�FA㘙h�X�&	\��aZ�9��V��-����ńvc��gl��ζ/���	�g��=�;�:��SW{te���%�tvY�y���{���m�Fس�=����T���oaa���7��K�L����ݟ�Nr�	��ĺd�i^�S,���׷/�֒q�����G�7�`]�W��n����,��P¿5G����㮗WQ�Iq=�Vd䯶V��d���kwv$�����QQLs��բ+�(
�7����O�f�Z����v
�Ws�R�$D�s�Ҡj���x��d&���C�h@ZCca�~�l�&$+P#
}�q�<� QU))0�j�� �l���[�	��F��͚/M�*ٽ�����6l*;#'[4Mp���.�3N��	fp���Q����[�U($� ƤA�
�����9�%u���Ք)�.̗�e[S*H.�ƴκ��
�;Bӫ{W}���.tH~����H����:`��6�� f��"łt���s��L��ьG�U�Y7�>���rJx����	�Gw ���<��F�s��ߵ��	��g^�ji���/�^�W\H({�<w^��6-������vJ�z��䆥��{�w9�._k� r	����=����n��=�stT�-���Lţ��454�q���ʨ�D�.�����<tN�V-U���d�{V��FJܻR�jK���q29e�;������w-���2�w�B�l[��7�t���Z�z;@(�3���3��#�$�MZ�w��[��b��74i��\���*
�G�ܺB V�Z���{x41jd�
ԥ[��O��5��gG�� �������:^�I���Y��n��Z9J�9���n�r�B�R�PSoV�m=�k�J�=�X�>���R�!Y��Y��=�%c��b�ϕAo�J����p��� ����F�'Gr�Y�̎��X����7z7]z呐җQ�F�\UYb���e�
�,c����I��7���uh�2�yɞ��n�Q	;Acx����m�,��(���R�AQ�Ok���پW|)S�2�
��XӾ�i?� �;F��N��w����V�z�е��t]l@���atfƊ��yZCK�z :�I ��ѫ���v�Z�n��(=z1���\4��ޟ��j5zq�ھ��!'+$DZj��e5�[4�m��Ћsz,8��9s�fv�`Vx-'�Y��}:���9l�g�:� Й�-�� �kx��[|�8骕Ʋ
���~=�:��n=",�rJZ1Ǯ���4�Z��������~���նe=�E��=�7�®��ho���	��ɮ�:��zS?S�=�g�l�˯ܳ&u�6}_`�zu��\��~�]���	XX�kIj7��v78U���{Lp��=�{r)D �DG���W�q����v�<v��i���'��޾�1��3�x&�)`��<�"&y��fo�>1@��Y���9��Wu똉�OY�}�@ [�yS�˰�aGT�{��Ύ������5����V�l��sE�q�a���o*�cTN�S�5���++���t����&�C���a;ݥ��0��4-���K�G;v�u�QGa.4�^75�+ÔO�#<[�����=�Ow�D ��Ê�j]��#�o��2�����b�7��.��hD|@��*ex� d�Vod]5�.���Gj6pPZ�Õ�.�P��)j���+f�b�E�խf�bA"�0��cnwi�Ồ 0jbC��4�%�|��/� y�ZRgz��whČ�n
[�U�S�o�XY��յG>7L���7����y��$k�)!b�,�_�vZ~�(W��s�Y��W���l�����a�k��>��@�<M��B�\�V_��/5ݧ�GlJ�ӻͧF�_�։��b6*�Ϧކ��Jjĝ��Ly�M�ӊ�kY|��r�kJ;v��W3�Sï��xG$`�t��/e������Jj�Z�0�<9Z�ྫྷ����OG-Cķy��ϰvN�]��`6Dg\�Ә��`@�Ap�O�Q�����{��@���Rk�{jΩw��R���L�6�q9���'뢡�'(٫�8�oy�;l?�#:
+ьό���-F��]O5L�g��"uy����"�@�C�4���4�3��5�q�> �U�N��{ۜ��П+	r��ho�^f�
�s���8�.�n�CIS;��%�B!�@p	'҃�T'��ӷ�R�F���]���t/6k��G��KX	�bp&- �Pl�Vc�.m��J�5�^�����Wc1��!��sm_R�7�sB��6mZ�N��׸L���_ݍw;Mn�"��wߡ�}������f��sTwq[P�%�6���OӞ�G��E3D,ח��n�/r9�	��{Ë��eE	$�g$�C�붜l87^�9�n1�����5)4s$#{����ӻ�n����" P�W�8��dɈbN����q�N,����WSS��\u彃�j�.��*b���$m�F�g��w}���le�Z�b�H���� �G]��>�k�?O�0ʚ�f_��_Xӧ#e���x_���:
pb��6��v�AR&�MG@MTl�<�_٢����{��o�6F`���,�䡞�U�j��L�T��.��q�H61�DF.��o�����y��}�~��D�%����|L�̝��K�ӄ&{�}�߫��[�κ�o��Y����Ϩ�!v���ٶ�wCi��I���٦r=^W �R���ىduR�H]_��Z醫���8.2���¤ݮ}��$�+4�[�MųV2EAAn+�&;u�,�8'.�Kkt�wX�d:㜆-9b&vH�o�<�Z���h�]�/�T'�ͿU}�R��{_$}ө�`��Y�j2�"IL��E��{;��mc���a_3c���}Q�������c���=9�ԃ���B�{7T#&ޭp�f��;Q!�����Ok�ڎ�̓'or�=������Q��V�1X!(�3�޼){^�eV@`���Γu�r!9�;��c������ю�����5�q�}����G��\Z깲��kZ�.A���<�fb4o��a�(�k�+zJ!'���s9��ľ�J~��e�_5��(�ۃNA,���<�#-����M�8k-�%����>���f����$x'���r�V�8��<GM�T<�s�w��^Z���M����y��~�`۲���e.GG]���B�懺J}Q�?�_c�Å��ֈ����Ϗ\�A���x��@+� w���/�O��7`��B�OR�_���+YN�5�!CPp��ePΫ압}�n?���	�T�����Se[4�nL]٠m?�=��#��2���ܓ�j֓�^����b��}bf�=mO�L4r^꨺�۽ɓ-��{���J�W7�P��Ҁ�	gr��7��e� �Q�;��_�������� >L-� p>p ���g@ׯ�緢Cz>Fz7@|��y�I[ܒqּ-h��N�,ߩш��rR�����das��rWbٽ~=a�gl^wK�qY=!�b0�jh�j��ӊ��aX�9m�����ۚ���L	��9<����"/�t���P�{*���i�j����;�{��
�`.ǷY�/^�3I#��q>��߆W��n��J(z^���5����1xL�}�.\[��������K���!���Z>F8�>G	ɀ��٤b�����~�j6av�P���̀�uPW�~=�c�;�E�?tQU�V�e���l���I�Okߢ�@����c��X����SB$0�LIx�Ő7״p�u#�<.>+s�U�n]&�d$r�rݛ9�� ��PSf�*����ӕ�EX�K4i�p�Ү�ڎ%�qks�ʐ���%�g�}B.�N�/�����6¾\(�]:1���奾㜾�'����<��(,��3�B�����E��������Zw:�'��D;WVcM��Y�m�i���'h�^��"ޭ���z�X���j3�c��9��=�j� ��C"��q>��]����84� ���{٫�ﲭ\:b[H�[VEJdR&/Cv���WoN	�}��(���B)�j�j~��Z᭵4_Ik���A2=��^�5S^�#�d���r�t�]z�I^���>���/̭)�H7o�5���{[��鉍�x��f�۶>yy��/���孩�VY����ݫ��@�_w熳B˩����W0�K�����-�=|gG�7չQ���Ԫ]���g,�?0���{�F�J��S�c�S�5h���O��[�u��x��b��~5�����u�������x��;
c]��G����s�P� ���%����9�&F�Zi�X�K��y�U�F{��ѻ�i�Ɖ4#x1���¨�ss��s:�I4���?z���y?m�0۾ݧr�ʭ�v�u&:��L�q�_G�ƞ�{ݰ�nk��b�w�q;]ҀRsSu��|i�B�]�N��_돖v�H��l5���<� �T�0 �"	s[�޾=u<*�ێ�p��&mt�/sP
k..���m$�.;���;�_����l�vnx#g2����å���� I���}Vj�M�.��G8{tV�BY�ۚ�S�X�|�fZr�S��lYd����۾��������S}'[=���q�2'�ч�H~ܮ`���OoMC��sf��;oz�xľT���myU�;|��O`�΢��W\�����׳�9�m{���L���/9^v���;o�L.M�=N��"�N�q9/�1C_Vg��t��5E����9�B���ǋ�N����{z�g�U��H ˀ	l� "�0	II]��(�y��wRw�#���ן�m8;ya}�� �� ��H(� �`� 2 �b@�4�{�%Ov��Y<��������pv�Z�����:��.P9��w�&�����S7�-����HZ\��=k[w�ݚ�7�}�v]/�Sk�#�1�
�k����0x=����Ƭ���f6ݜЕ:�Y:X�K�?�y�>%kV��l������ˬ�<��/�M��q0��2���<",�����.�����|��ҏ}OS��~�g}W{��mW���>�F�zP
����N���v�����h���M*Q��<kM�p��8���N��u��nbe��#8��d���r��[�9q��ؘ�� ��k�	W�N��Wھد��YzG�-к�ź�4�>ghe��<�����mŮZWVc3y�������z˞��Q���O"d�FŴ���1�J�τef>q�Od��z�/��X�_�"/�*��k�������d��b�B�Q�%*ݵo�:�>�GI����v�}AY�..����#�:^Ϸ�	�z��:�{�,��7��_Jq�6CF�1 ]���pm⦌;�=�F��9G~S?_1�t>���@�UV����2��E,?�V�n�����U�������0�� �@��,�?�J�e^L�{�]��GI�'3����+��Çd��':Q�����k���ub��9Z\e��[���Ky{CQr�ܭQfi�Me��iU���+&z��#�<J��<����4�jн��7�"1hzN�UU�`��wV�={�Xl{�3�Ĭ8싎� }�]|t�+�W�v���eƈ��@f|���z���*FHU�X����c��jع�n�8\n�i���d��E��p��`*����m��Rx����&�c|"�1��P�op������\w�j�=��F���:�ەp:�����F�׀��U�Y_j��R<���܍'�[�u�-|�Y&n�.3���6�&���= ��s>K�
ax	����}�[Dg�9�G�Z�_��9S�.j�~��)�ݝ���9~�u�M`�U����{��^������ϡI>�.4��oL֥a�� �"�|�rA����]��yע#�=�r�� �mև|o$��Uo��'cs�v3��4���ៀ��_<�3x	�3���c�	�-�jc�\u�ZP�t�K�����Ϧ	c|P�jm�#��]�h��J[oo4�N�E_~�9w�}[����7н*�G�D;�l�0LuP<�HY�Z�	8��X:��MVN�wUw��Y�S)� �l�ѝ�����;�u�����Oh렡�fx
�|��[ӫ�.������݁��U��;��~l���o�]����}��5rC��ml�>���s�9+�.X1�*f����3�n�1��E�:��P:���w�xd}��}�t��������+�[/�IDwE�Qɇ8�RU�J�ec���A������((j�H��(�<)0Ƣ0������-��,�S�Fy���4 �Tϗ��v�|tJ�:���x���o���{i$�W���]/@�����8u�kF��$U�a�4r����g_eL��p�/5�� h�C�LOL{����}��˲O���ko�;�]A���r�ᚡ/}�����ȷ�%�_mJFh��͊w�u����Z&�*v����BY�����*,ׯ���usՇxO�*|5��5�
��������%�^]��=�xY�۔�}ĉP0��v����X�ca�ww.I��6��C3�';v5_���M��|G9�k.gQ��O�n�߾��zx�������lt4�J�ϙ�w�\���z�*�A"#MX@���2m��ܭ �R�R��V��`�`a�E[��!BtiL"�h�55O�a��	�H�Ɩ����;�Ui7e���uȖTՅS')�	ՄC9x	0\K=�c�cS1�5$��T3'Z'H٣���vFd�D�_!�EA��L4�Zє�	mS��1�*T�HQ�D�^e� �#6�\��BW[���zFu�pYH7�1���������Z%b�47��B8�ɛ;'q��Yo��k��J�"�b����FYX���^�� �L;�+kZ�'�QV�Ԧs�n�R=Շ���T��p�{��th��(ړA�˓�׮LN]r�zS��k�z�=w7m������c��י��Z@uE9�m�u@o���@�7d[�՞t�)󘪻zJ��31k�>#���C-b,��|��,*�/�j���u3b�[�#ͣ[���i�U�u!���8;)��`vt
)&c���}�m�αJ�Q�B�7Sr�$	,6�;Ś��޸^I+XT����"&jm������nL%H������y�c�� u�oV`��r�un��Tl*�&�`a�%=n4���	GV��|Z��h,���*��$��^d�Ss����P+FN�	Y[i<ӎ����s;�`��Y4F�� �J�Z�7B�$Ԕ��M
"��2�u�T�;?���2I�j��%�yBԏ�m��N����&{�7N�U�d�hLu����2�6�����/��;YEs�t!��6�m�Y�,&��G $l�V��}yzn�Y�[59{\�wdt�3����BIq����'�b���9q�����;\�S̗f��^2T�z��t�nP|��xv���-��
y�`�}�M�Y�Z�F��s�p�]}�V�lԇ2�y)5n��b����+K��s���kA��K��̀��Q����(���]���HW�`W���!�I̹H󺻡�Ӏ�V���om��˕�Ǧs�x�Z,@kш1z֌�a�ok�C�����\gY��6�v�#�o�	3��n���z�2޾��	����ή��P�'��9��2/��.�[ֻ^K�q����n	��b��|żDż$.��;���$RE�WC�1^�?�q;���Wz8K��)�b����N��F�Z��ʾض5�N���茨�.�g_.�C��.��5��9�y��v	D:�����c'w�Y��%�q��Hxu�~`���@^m�ن��<����X��n�m�}/f�_n�	�5�8��Y0�ŏ�8�o[3F�\���1W����7�E3��pi�62�s&:S:�ewSޫ��s:M�Zcv��972Ԭb�:���|���q�FEkcr�VRR.���tR;�/Q���9���!�]�쾤n��B+��]s�G�:&����r��C�E��`����s���'T=0�ݝ�bOz��B l����B�d�p�+w�?2L�U��ފ^�k������r�������y�q�^�J� �{hp�c��ѯJ���X�d����{�G_<=���y�|&�ʙu��2����=�����^��D���-{��0iKE�뮑]�+�/n�πOv�!�d�qi���U���~1ƑcC�q�l�a��;��e4Ŷw��r}3�ϭ���T���b[�uS6�MX�Q�6v%����q%�\5�����#��k�`��[,�)x�O(�k���:[t��C����� �CGX=�h����ܦ��ߦ`������6"�]�}�J�0 ���t&�nY��O�O)Y<��X�Xt��JEzK�.�p���>K�2��go�s�&��i�s�"��� |DY�9��!|���"���R6	4t=s��ڵ����b��
`� �><V�8xq꒑�3b��7>�v�s��lJ&�����C�ɽ�[�Gp;��'�bZ�T��[	��@��	�H�$�G�[�nR��e���Ō�s\jY�W���rrٷCz���b�J �"	!�r� ��!Lb� ��tCP  �wf�u��JcB�]I�ar�6�_�l6��-N̵��MÛ�Փ�*�%8�yՎW�q]i�ZT�Aس�¾�f
���%x�ә�87�vߟ��[d8�[�$_�M��m�Gh�
���g���(ɬ63
��ח��/���w�gpt����������W�T�b q�#��au)�7�r�A�����9�4�4wuy95�)����v�s��_��esy���~U�L.^�`���riQ�r�<
��n#�G-'�
Q���^gϷ�b4����y�GBZu���û��Z=�ܻ�����I���l� =کѐ��t�kwi��%����=����[<��#�))�����(^��B��{q�KH��~�~o%Ҹ�ɜ�/zeh�m^��y����W�xFŎcѤ���Y>�G�G�p#�~�T����JU��j���~f(rp�����b�c�VD��6L8�J�t\)�:��{ ��B6m�uuةL�Z���Zy�P�¡F�M��9,m]���K�u���UlW��A�Oy��QT�ݷ瀩����h튃.}��D�|��G�،z��9����R���@$jl�1#Գ%�.��.κ8�M�U	MV!�
��̓)�pI�E�D(2�B���z�
3#{|�Sl.�<y���V�+��:��\��A������nQʔe�&#��AWfw�h \�/���w{��KX��^ǝ� � ʮ��_@�w�k+�y�Sy��Li��@2�) L���G��������}q �M}���W&�e !\��؄�ݎ(�����y�#��Ff4�FJM�6ᗛ�ˆ^�7~Bc�j>>��l;�V+���S��T�c�J'�א�4§F���NU����!�^B�9�k����?j |`>~�τ����N��߉�#����&'�F�xb��?+~n�`�z�#�����h�PR�.M�n}��Z�t܏m�,�Z��j/Ӿ����I��4���P��Վ��m��@|��5)l�p!�D�%�TGL��S.;����Tŧˏ��\��E}�֙��˅�^0/�97~�w]�&�~��� ��9�2��H�H�ʏO�hk�@�+�U|z�����k�i�^��\|�'|��ƞEG�%�1Y��x��1Z+,�������Xs�C���,.:(��i�@����xT�Tc���r�z�g�?L}� D�@`Ao�v֚���"�]w+L�z��Ԟ�s,���@$QFq�@� ��6��V
�g�*��;��ŵ�Q6j�����ѻ$��\:����˓/���{���V�zm��ӔH�a:�X���sx!�`�[�y���?˞��2�Ӫ���'h�x�wc�^�^az�3a�ڋ�j�Ӳ�2����F�� �r�>����Xz%KoQ�$l�������S�ӝ�<#��!����ÆnU zb޷$֡��O\(�ٍ�z/�z�AU��w�&�]���\"t,d����N�R�BPV^V��`f8�q+'����>��_��!h�;ו��f���� �����G��3	`�����f�� 2�24�=M��@���qy
��G�mt��
e�ҟED%2��!V�#��X���;����y�}�zH�}pa�Ք�)�e��lѩy�p}sv�2��g�K8�Y3�/�/vt�1�8�ɚ���;'򛶅��V����}}V��4��;�g9���-$����5=��� ���ѥ�vkp8cY����.R��'��Bj^g�/��ct����s�7`�A��	&��s�޿�IF/��Vg�! ��ϗ��O:~Y��ғ}�+����n�f�әy;�b��@D@��IUU���O��j�p�"F� �;�,n�jƙ�v�Ǵ�.�
������֫��tα�����z��y2L�d�5�=阳��.V�f���5�w�w/��k{��X���x%N�Z��6�:��a��
�qs���n�2�D0YM�A�.��-��Sj��ǌA�<����79���3�f,�D`vz�ܨlߍ`�_G��#�1��� |��٢=���m�Ĥp{��ED�2��ܱ={F:C9w��L��,?��o��'d�Q"�Uxyʔq�mu��r�O!�ա-�n�g��qu'�ݧ�Z�L����ݶײy��v��Ɂǧ/�:]�)�ዷ2��(ۜ{������"߂��N�����vܞ��U�nvL��Y�\�I�ZyA�uҷ��Ȓw���m��W��}U��p�@���d���U���s��񻟍�+�J@�vm�
*!c���y�Iޡ���e�,�F�b��̢��o�[��j�@�S.�o�l�ᆋhmD��:�����cY�^7*�b��n�|�'�|�h���GO̞z[����t���ù��gȉ/b�9�5
[��NMp���c�t��-e�o*Y����3�&Z-�Y�)�C��f��0W�.qV(s,�V���{;��U�KD5�s�4aX�Ψ��������;V���s�芣��ѭ��A�+��a1��
s��H��L�,�Q`���'}PMr�	�Q�v�M1��Ѯ[�g���7l\�@r7o�f&:�=�8���!���L!���CAF$���#��`"���NÞ�!�(�TYΈ��5�����*�ɟS��� z����9�_��)���T���T��&�]"$=�Y�Ģ�>�UD�m�r�ͯ�i;��`���8"Vnn��n���!��I�n��؞v���%���hN�I��-B�i������|r,�� ݀MgG��㫭�䘾����c��5��7��E��P�|K�c	�j��v�F�.f�<�D�j2Q�7���і9��$c�Ѷ��ʔ��d��/u���~S��"9�e�dt��7��F\��Gt�X����>�ƧC�_L?n�{D+�|���U�)y���n�J��Q�h{�����]N멵��U��y<���_����+���'v/�EFn�s#H��gdfI=O��%e���7�k�D�,BI�I����$������,o%bZ�Җ�V��M�w�2UI��F"�(�A �"&�m���EA ���:���Bs�Y6�S�]��lj�Y/�WRZ,t��ijv.�缹�o	��;��������<8�An&q�=}�@����2T��;��VF%w�����~�P_�M�^#�Bw���t�K���^� k���l<��Qn�d�I�R��GRp��Υ����>ޞu|;ԵFN�A�s"����1��Gf�:Kv��XP ]��?^9�؀P�A]�����/D�ˋ�7.<��h�s��<�]��b9#iDF7I���,�A�͐�j�'�B��`�up�J��"�"��XV�^
y�=�x�_`H}�_��`}�R�w�oA=��}���v��y�&CW�꽑�W��*ߩ��J�� L�Gc�
�݊�]W5�E���gCR�zl��q�#a�2 Y�þ��\�I��
���=s�T�o�M5`�K*����@ߥ��[�a똨��*��W���}"8a�]�N�$�?l|��B3����P����P�QW�lQ��s�����>�7_�j���o�T�";��(��qw�kT�qݙA���+���^*�wd���L@DE�(�o�r�)��vW~���8�!&�eIA�j�UӑfHx�Y��)C�0S�d���P������U�Y��hb�Ekk�9� �=Ǣ�:���K�;���ѓ�� �Q��N����U� ]��n:Q��N�Η�w���eN���� ՊO����v3uTwҰ!^��}���m
^~�c�6�<��{ߥ/4�?Y\l~�]̷D	��g*}���s�{��v�K��K�t~a����9dö�j�����4a��fݠ �}�n��Lc\���W���(�n(�Qݜ.�q��K�~����w�GR�����]f���D��C�jS��;��_ݏ�#��j��k�v��h;�ڔm�����$3��z����ne �5&�ˑ9��Ct	l���,�'L�`�T�b�j��`�{���Y������|wF���Σ�ˀN�b7�n�ڤ�� �]���*�>j�~S�ԝ
n��ף�!$��ʋ韶#h�9�B>?w:�'��j�Ġ/o��������)~�	�/������)�T�f{�S���ZB3�vz�.�uٍ����s���ر�����R�H� ;^KҬ�'���⼯OR/qp�Gb������4X��W�/'��u�G�J�3P�b���wٚ�D�][Q�\�Í ��Yt@V?�H��\��L�pd��G���mwu�v�̽� ��-��x�ל$#:��f�k���e�n�Y{�s�r-�T�WU�(�4�'�t�BS�����%[��4��f�zT���e�zFT�> ʀC\4{�櫨�� 'O����P+c�^Py��^T@��6z���y��E��k�F���S��Nx��=[��Ɠ�z��E_�O�Wr�5��ɾ�v���5��uSL=?h���#�'>��t�s���"�O�7���	{�ʩ�Qh�S�{Ne�MG��Yo��ܢ&+�}9���O|�GA,�Y��ZP���j��h�ׁ]�E�HG�W]�΀�o�Z��:ʹ�彺�7���W/{�����&%O=0���\�̫��lՄ��_ ;`눞�{�L��Ґ��}�CF�sGT�2��ix�i��RtC�i���Ի�e�_�ξ�Y<�@��׎����i���hɹ��m<���Sy��9wiq�#l6��v'��U;��H� �dݮK)oç �k.x;|�3X�~�eߵ]<Tz͍�w��$7�+���k�ӣD�u���2��P�M÷j��j��	���@�3�Ƥ� 0����3J�`� ��9�h}=:�ׇ*�g��v�n�f�6s�!]ȼs��`q�0`�@@��K!C�jS�s,�d���Qw�x[)u1Z���A��#z.��\.��I��>�6�����(�����]R#jﻮ�W5��R���V����	�0{�sIQ��ʏA�㸹�d!���f�O�\��:���;tWz���;�{R^�(��r����v:D����;�%e�Ulō��Q�)M�с�Y�����z�.g��c��nn��v���d�E̲*���)�C���u'D9���[����va�i7���u���ZDSN.~�2 � >�9��?LnB�7A��`K�4مw��m��]���#X= �V_�Ǫw9σU�*8�^3>���"q
8�=�ۃ����؁"�u�o��nШUc�����Ք�L���>�����<���۳���^�$?1�Hq�Ԧ�(m�� ތ�s!��������/�<�umK^��y�"v����Q����\T���8׬��6?G��{k�^ER�z�@�[�|������=A|`m�2,������v�m�ъ��"��,���q=��<�܅���d��,�[�ו�^�����;�Ʒ��2����l5~��j�~������.��/ i�ӵ��V5��=ar�c*�P"Z�#�d�[�lT�Ϋ�ZkLI�#
�6UC �8�F�Q�`�z�H��!��!�"��c8��c6��{!���,6(f���ge�e�0+&@N��֫r4�pA�Z�d�j����!� �be�
ӊť���RQ�.:4(�Q�		!!MU�`^R�"�2L����7��~��7�Vo�1����-�k�� ĭ9۲��#*l	�y���뮷����a�;�}��KB�Z�R�޽�I��1W^!�2��Od2f��71u��@ʳ$�R��T'�$2��u!��z���Ȅ)t|�=y��sC�O���NsV��Z[����z��41#gLN���3��� ��d'g�[�s)���,/�VU#{G�3u�-�����Gu��鬕3�BW]]Ҁt�Yٯ��:{�u[@�����Zf�MRY5:YOY&�M�A�Y��,��
U�a��Z�P�����>�ʂ֕�S��h׎�U�a�LF�w!:CԌ��� ����2���%
	4���J6�2�����BSt!b��hwY5PL�%f���",I��A��*$���c�u�fcG6WN��W=ڿ�n�T/r&ȐY$�R�t���)JR�)9��)U�Z6b��`$�`v	s�4�Z�vS_��KD�y1j�O^uk�cu��F�5սnV���KN�<�7p#`e�{r����t�l�����5��I�>������XB��]H��j�Sx�L�N����4 �a5�-����4a<����i��#�$������!�̘�]q]�zm\�y��o�ˊ
��7��e܆�� e��I�� Yd���'�L���'ǡ�ݩ]�k{Z�����8=���ς�ǘ���1p�W\�[���v9S�j����W��rޜ����$��t�K>��J�M�7����T���S�v�^�(�|^��f=2��uBEEh��v����Z$�m��E�4�K5�W2�GS�wWr�R�0	;����b����@�pЪ����&h�7%��{)E��@,�u�k��$mov�6�ru)��EoW�WMolW>[{�d�R�x�)��������W�\���-43�_�M��2�AY1:�[��T����>�]�M��]/��Lȗ[�)#xu'�B�;��	sU�}��f���qI������v��uws]$뾊(�kO?x9wy(�Ԍt(���QS�4Zt8~f�F�о��g��6_�R\�s�w1�x�6���g���N��]��~������jK0�-.j��x�}Cm��T��˂^�9-\[{��C6�آ6m2�}����X�f������n�`�ԕ�bU���m�;"�lc�V�Weds�v��s4�s�|���hK�O/;��T:{u�"�wM�G��+c��t���Y!]��ZS����I[��CWu��O
p�m��K�33�t���b���ט�b�fwU���sK�aǧgr��8��$��/��mO��A�R��-ݙ�*�3k�����-�6z��	!*h��-e{�P" D
��T�����a�����k�$:�Cj���=�?	^k��I���'����W����N�涺2����̲y��j�w�F��;��z�`k#i��9Ug�K
����Z�O�J�v����p�ßbh�lsJ���Ur�6�[K���(\�d���T�>�R�[�y�;0�Ĉr�3��L%~b=��A��cȌ3�_r�5[��$�����Ft%��fa[�f�/ARU��\>��Y�/N@A�̼�xBq? G��Ч�B�FO<�l�|k�CD�~�ta���M�Fb����1�x>�/�_�p�3�V���}�H9��ҥ�Mx�j���C� <H�J5�Q�!�`�y������{W��2�Uۄ�N$�lj���l�����p9a[� �
\M�&��-t��2|��V]<�%ߠ���z�Z2BB��D���v�Fn�|G���0��a �p��(4 Pb1�ᩞ�kOy���if0�+C�x���x�x�mVs�A�DA'q8aCmD�b(	�-ԩǻ;;�/�ۄklDJ�cE���*Z�,W7:��Xō�=]���]tb�K;9C�y��n.b[�NYF�jt�,|cg�Hi�������X�Yܷ�Q=MP��=�����ǵ�M�#�j5�8����)��Z�m^�Z\R�K�{�,1��O�d�t�^V��,g
�jy�3P��I�Kс�,��p�N��O�Ԅ�@݊�b��k�f�D���E�� GkW��	���|,�O�3����� O})+Y;򛹶�wwE+Z�x-��F��Z�N��Ůz|�����u����Ce|�3C��)C�ͮ�ӑ>��h��(g�3y�gD�{��7=|o�����p�Aךݢ�B��;5�q_��3o�����:۫"�����8�Kr底�#[��v����ǒ�z�C[��`�p��T�����g�K/�i�[�Λ}rNSS�<�ƭh���ʲ\a�����*�?W�4�6�%R�}�\�{��'&����p��#�D	���m�>���E�[��Oʁ��M��Ɍ?O�+:�p����=;(�{�L0A=��xc{��&�:ܥ��c��ݖ�{rO����`x�"�"2��cS�C��}���@Y`�1���P/YDDH��d��k�%I#��'�*½��e��f_��7��|�^\�X���pZ��ji��ۄ���������p�|���q�cu���S�DRֺe�J�:�x�"sQ�Ӈ��E���Fy���$�-�3���[�j*	�~�M�-%9�E��5`��	��B��Tz/�Sz 9���l���nt!�(�-�	]&�&��:&9�\��Vr�\wCv׈]��'�%fæ�~s>���1��M����K�I=�=�hy��B�T9�;.����6=g$FEQ���hf �X`�K��p���g�zG~.]7&��*�C{�7Χ*�o�(]E�	�ڌ�����d"/x�+��S��S'�l�d�SRǳ(aE3��m/��1�E��Y��>���NrR�M�[��������>����5��1�������$1�+�="{�.��u�9�n_8�ub�vbusN��]F�dF�`t�ؐ����ߥ�<d�)]4^ĒrY���6�I�r�# 5Uoc�C :���ϔ��vsv����n�xTD��?j��T��g�� �ۯo��ջ�&�-3~�:���T��k�:ꛆlp/c�_^ge�2<p�G���8�7�l�:>>ֶ��Y��7��	A3��� �R���Jwi�cTt��\4Ky�3�҇x��5��s���Q�`���G,�|����3K�ȥxpѱ<�|��X��K��Ļ��s���D��Q�(po��ת�����(�P��3F������a�c��ؾ����ş|-e���0>��'�%�r��{4�3ϫ*_)*hwk)QA���l��~#g��y܇���>�U�E���k:���/=�9`f���5�jz��N�/7� �:���y�&�������8�܆�s9������G0�UbZ��������>��fp7F�a�C�Q'���ʚ�\��6'��S:%���^��1�__��:�v�%��d���7��b�Es��ԥ�;��Ra����Њ�C�ϩ��p�?\��1�Op�-|������0��7�DtܜE���� ��h˿�OL�0�3s3CU����yN��ڶ����;�J��L���$�1��i�/��UҜ��c:�����������W���-Y���ͧ��w@�"�F�	_CA�;_W,���&� �� �]�����Rz���&w}�$՞���3��Z���=V-��>~]��)��L�_c~8����a#Ph@�h������ܭ9<�+9�|�	h��^d5��^a�gk3�p	8DQ,!9Vf�fo{j��o^��>=	��v�4-4� 4��M�(����-L�z��{S�+�X��vI�/�xs\sZM±��M�d���.�ncb��/vfѸ�T,�w�x���O���������v�K�p�PܧA�h�������s��c��%��6eyU�y�=�`�����"�����$��-:������"��}C����:�GԀ߹�(�"'��N� �B�=�/�[��cOe٧*_��ݶX��¡�g��+�N�C��=Ee��@�x�pzLo�ŪNjRS������o,:]8�k�B���A�k�GH�6��L�0n��c�&�"���g]WV�H�\e�6}�y\ �|<&�ƕ4�3�f�,�����\c�������������n�ԫ��4�+^���D���0�uM'��o�O���;>m%�����c���7���)4,i��mj�݆o���u��٠���闆I��k��~a}5
�M��2=H��
�'�{VH��P���
�%	=IC�L���A�`�����uxԬ�1���'X��Btᢷ@n|uL�ʼ���<��|��;�����Hs`)P��x�I��)9��l�%7���;��4'W>�(�.��5ݰA �R�Zd
2�)&�gd�-��8�r�Ғm��g?Is����v��}n�����H�K�}�8Q�m)Na��sy�h��b�k[�+;t����ڏb}N������iX8ׄ�_q��E��֕��´	��WI���5���onR��n
��7�YaF9����%
��tIN��{p�hWB�튽���[�9���PL�k+j;�F��щn��n|�����_���|G�Ip�R�u&{�0��P�t�XT�hM^A0Y]K��dOO�O�?�� p6��Dq��H�>��u�]�ma3h��ڥ������T*��yu�1�fC��%PXp�2Ǿ�c)�Na:.k�)������G��Rz#v�Os0,Q͘��C�D����kX*=�TGCΝ��\cժ��	���A!��;s�q)����5�qG��5lf��:�r�	59l��tm	�vx���s�[:��WM�'~Y��_�g�=�������XVf83�2f+	bG���2=�l����Tb��$�y�գ���F�l��J.$A%[jQ�)~�Sh��E{�����>b�>�j�" N�O���X��W��@Һ�v�o36E�
�k���ʳ�7!M�"����Z������1z�j�� � ���d^#��sh���􆫳߷�`�6G�l��PkfLD�$�d���� �B �]2�n�USR��u}��VӺ��� O{�y0;�բvk^.�"�� 9��u�M?{"^i��f@��@\V�S�|�E�=����XQ�E��P)�2ڒ�Z��]^��2˦4	��Fm�3�=lYʡ{w���e���z3
G&S]�;;n��x�Z�&���\ޱ��1"&�i��^���S���g7��3:�ۘo�37NDM D�(�P҇�[j�4��RMSFM[k�n��5���1U"9b�cc���3y�i��E��6j�#fH"]|�	�Q��'.A���
����0��t\�ѡ���b$�����q�w��݄�q��aiD��Fi��Y`������4^A�e"�+��i�� ]�	����=w�9[xޏ_[B�����ZIG���*��/����[dS��B�4t| ��/��f�K݃;n��^����II#Q�D������6��!�jf:	�A�54�4�>ڿ�ek'�ד6{m���s-�`+��N�.�jcܽ.�؎�K��$����F��+�:ּ�Kk�����/O�L�wW1�z�n��+b�i�]}B�=pP�)��)K+���áU:p5`7ޡ�a���!����Og����̮�9���jd��=�m@���Ϡ�Z���l�^�Ub�Z%Gfc@!!��^j��AZc5��)��[8u�j���l�dԖ�x��#y�}�iGR�{�P�d��7{;�v�g���,ov�ruse��J�u��u�A��ٓt���Cm^�����7��Ҥ�[� ������K�[�1f%D�\N�9	k��8'6*�J�؋Y��\����1eU\E�Qk��L���Sv[�6�?��|� ��#�s��.�H#�����| ��@ ���[��Szkϸį%f�D��t��nS�-8���&�'6��� Б85��E[O��;Ҭ��`���#�)�p}Վ�}�Q� �?n���ڑ�B���|����B�}G�y���d'���Tϣ�do?Oi��\V�*Z�s�{e�[z�a��n���[�j�N>̾;���}�}-p�p*����X5RCfJ$o3�X�yʠt	����~��c�M�,�c#����A;Z �T��j��S�Ъh�J�����
<������4���< 
�gt{����c�m팽q��pX���Gi���V��13�ML��*U�S�2b(zD�әݯ�yW;Ѐ�<�↨z�͸{��<�F)�}�sh7C�S�IVqΩX����K�01y^���v7?಄��\x�d�7�g�5�g��k�۲�~��r�5��Xu!#�$��1�jr�,��nF�近Sk.�k�ٞU�6����k�_��P�7H¢"�'/R�O.F0��g��M%M�y�����^@��B�L�@�O�i�_���;25�W�c���_7B���0�/�����]޵՘��W��jD�Dh��*�DP���rfٜ��I_�_6j�=�W��΍���u���f�볦t�k�Eo�>	Ge�'n�ᚣ �z���^yS�v.ZCf���I�!����%V��4D��>ᴏ�,7y�bg���ǘ�_�����s��N~��x��\�P,���["�:-E"���h�	p�<�<ŷj�h��α3�E?0KG��A=����Y�Ds�0O��U|QY���B7��f.�>�id0�h�i��u�����5�)@�L!������e��J��X=����M���A�W�	�	B#O@wA�{}��;V��U���Y�Dȳ�\�*m�"I��vO�+"�=)n�T۲*gM�ex�)��[�x�V7��t`HS�X�!]��mfk�v�~�������HQ�w��v�r�K��ZUk뺵+�Y�ڽ_B{���Їs�5X%#�c�6ab�Ǚ�w��||I���j�2��u�zuq~;��� ��k���V��]�g���z:H���"lXJ�����>�v��sʑ3G�ғ�Y�?����	�H��4}.R�~�%��.�y��Y��w�G��{�4Q�&	���1k5�cK8h�,qJ����vD�f��nm�9ؕ�
q8:��ƕ���Vճ59��=��3�	a,v�Gmj3���'�>KP�Y렭�﨟GcɖB��󬏾��^P{����,��E��d����Ύ�~g���3�0�DU����);zk>��kp׋�-��J��G}���++�'$�D?}~�T6s�����>0{��&�sM���@=�?�E�}8dE|:��a�Efg'dqf�g)���ȁDD45B#�
�����}]�s5{>XRD]l��(��^6>M��z�Be�����]��${f(�"= -�H���(F�R=���s�^�=�q~�k�(zF�S���)T��^#������$D �e�k�-�2퍃���� G���Ǯ��x�3:^w:=�hzG��H�N\�c��	jgk����%W�ڕ�������$�񵕵=-r��5�G%n�ƕ��f#�K�����&���gUP_DH��b���:��ɛ�����#&�4�]w��ѩ��Y
�%d�ɷ�P{��4).>\���Y���/q�F@�
�jjݛLǚ�E	��LhF�y�y=����\S�4��7�N]�l��α�m\�o�m8�<a�����$����>������)�8qy����
j�=/�]�y��(��R���y�u
"�]�{C�k&��&�Fz���(y���ЀD���@"DG��F  �1""A?��?���� $ 	� (�"  0�� DD�@� �7�� " DD��� ��_�@"DG�׀������ "#�ë���������{�@ D@��  �D ?o�}��" �4�  ���R "#�#�?��߰�D���_� ��� ""?o�@"DF\@"DG�_�b��l�"D " DD~p�D���|�ο " DD��D��~�����Q#��� ������?}� D���$` " DD_�����e5�8F$�l�՘ �s2}p"A�|{*6ƲQ! �mD(T���Zd֥$i�IU�i����QJ�iUmf* T�B�T�eJUT�KZ-�U%P�� j"��%Ѷ*��BUP%$P�  U(�WZC�TJ5�����U��B��.�U��%E*��4��V�P,�*�@�kT�"�i�_M]b�RN�.�V�[j;�UJ6Ԫ�1QH*�U"�f�T�ʶ���I��XU����UJ�ݺ�+f�RJ� %MB�@   ��     ��d퍴�ݔ��%	T���UVf���%����TR�I�(��)T(�QV�Im��J�**�$5��	�T����m�AUYmm�R��(��T�T���v떍Dɩ�T�ՖT���5T��]�]4����f̠��u�E\�5=�Ec*(k)(%R*�J�Y"��e6�=2�+Y��f�ɔ��f�Qi�V��Z�̐Q�;�Ӏ�ݺ�]D` 2���@S���Z`6�P�P�p t.�ۡ� P���(�V�uC���݃@�u8  d�U��i&
��ȶ�
[h� ���$�m�)T�T
� �Gp�ձZ .�P v�MU�ڴ�����:0Ѡ �,6��]��4m���\5� ��l�
������ZU*s@5 +R��JΜ�f��0����@tLV 	f
aF��3UVP�j�,K�NZl�hP��-UB�%�� E	@�
� h(�]�m�h֊��pj�JѦ˳p� ����GJFVt�J���i&��W.4��6�;�0Pن�$� .�Gd�H�eEU�Q�D�V��uR�� i��Med뫔iv�]մ1CJ ��X v��ٮh[Jt�umvӋ�A�]-�;�05���l�S���IB��[�! �H��I�B��U��Ҕ�]j�r�+K��gnKe���wF6�5T:[v�n�ъ�cQqӃ�풊h��:�A=� �K=tP  �CCv�`      ���U!���E=�	)*��db"�����M*�� a?���A�d�xFHi� �L@IJi@�"�ؑ�d�7���Vi��9H
G>�\#�쏙���+�ϝ�G�`/���"#=#�� @�  ����"DG�@���" @� " ~���w�_�Ի�Z$�r艑R�ֶ�r�A�,y2]m�X���]�k2,c"�L,�tY�P8��-%���_�ɼT�����Ǜi��@��ܬA]uX۳��fFz���Q�p���i��ҋh�d^���-ˢv  l� ֒$%�u�ճe&1Ie�n�*�7N���1;�d�c�0B-�Y�!1��2	�h�,e�Z���6�r�~�jo2��Y��ʮ�� ��ٶ 1UW
�X��ga ����QY�7b��`$�^)%-(B�f���1p�k,�9+J�e���/�����P�4�QL�6H"-r�^*h�KԵN?�ލx��2����lډ�j�X�K)���IB:�x���z-XF�"��U`4�e�t��V`�T��q���
�*ƅ�r�����Jf	��K��4���kϮ�Ԟ�l�CW��/H���B��$+=T����F)�\؅a�h�#6���];���f�4#��oF/�yzR�%����\�v�M�Jf�#.��T��;ۉQ��N��T�=�r�Don��^�H��3J�m��n9u%K���n(T44��g��fҠ��hn�	��2f�G�2�u�7��]��7e����N��:�KáMބ!�U�w���n:V]1f⩧!��<���bM|�ͷf����)�oM �n���
�W������������j�����i�C�DZ�,�P�s��I�֔�6�io�F�,u[��Xz5&�P#�K6��l%f�b��pb��e��łO�V�=	Pt�k"�X���@��	r�Y���cӔ�e=�7pli��L`5��3D�is���HXB��s�g��{����h�؈S��MT	"�%�Y�B�kn٘\V��M��4�.�cI]F�5k��� �J�n�Uh�W�V̥rRř4ⷈ'[��Cr�I	R�A��О�B�!����*��n�b�1֌�*��(��t�7q��bM6Mj�/(9B��U���N�M�]L��e	��� a��$[�`�(��C}r#L0*J��i��tq=ߪWjV�Vs�)h�m�A�
�,n�V�i��&�E[��4
+p�d����ej�A$%L�"�^ea�siŐ,D�5�4�6�Bv�Hm�ٽ���"�~-zTD��M����9[��d�`��U	j�p#v�r+ݢ��d3��Պ�����-ڽjdCF������Q������b�ɳ)4Ҷ6�
�n�yiA��׊�ҝ�oq99|�,58���h�ȱR��wv��ʺz��B�ډŖACK�|r}lb��Re�Z�ӎ�a�Q�KE��
5�li+dct$�.�9˅t�ͳX]eYZUǷ o�(ۚ$�y��+g�	��#�UT��'PS*U�Tl�R��1�O�Q��e9�.,��C�e��ۤe�n�mZ�S�,�ǔ�0�7(�i�mD^B� �L�z ��˧��3X�6�olM��1�eaf�JB��[F#6lׇ5�4��͈�2�$�P�Vf�F#rލ��s�ͺ�q��P������RykԸ�ZY��C.��X�V�m56���1u�Im�Vk7j�tN���X�8�D@&�"N��@vK����HDe sY�v dF�"��s�mk�ɑ�ҵ�)d�IO:�;�����v���M�#���V]&6IDkgśA�B`3�Y4��r'W��5�-ѣ��W�[�	�ȭ�OQ���]�jʤ/*�Bi���f�
�q!��	�2)f%i��M�2�@�YpŔ��gm������u��:!*�;�w/�GΓz���ٵ7���l<_�F�+	�z�V����-E�QX	9�P��Ð�(0i��N���f�l�H�[X�gj�؛��/[̻��	w Z2]H�)���ơ��=��@��L�Gb�æ2�B�Dz���������E=Ÿ�\:Umŉ���V㽦�b�u	�F^���e���#&�:ku&RT��y���bN*	����R-�´m�B  �G�oem�]+Y�&,���a��ݙ/M
	���aM$�i˻���9,�c���i5tM��-���Lu�]��IHxl�u����E=JfVnd4�Y��9-�[�kvdR�ǓfZX,K����Bx��"2nͫb���)-�͚���V,j
��WB7�Y�:��20kv�(m�L��-��*­˦��#�]&����d]2tn��Yc]ej
+ՙR^��[�b6���Ӱ,�f�
�^���0bw��t�;���%f2�$����Q��t�l[պPϭPe�w���8K'5J6CW[	��.���ԗ��j��x���`Z�h���N�Y�y���*EMv^
R�g6���ML�8�������Y��V�wi��S�7�2�}�4��.��-9�����T �+�3/@�aX�2д��+u&�iXc�Ms�z*��9xAiq��\f�l��p飂u��F�ݡp�.�jӎ�b�1�án~��2���L	,5-�`@�"���M��Ү���Ȏk��F�
krn���Q-�rE�L�?n1c8�S#�[�I���r�Y���ʱ�*٤+2���o-����oe��q��2�l�
∫rM�6���"v򕖒LU���XS���
����v���e��@  r�X�Y��H{�k��VV,MnB�{(�/xVjb����K��PgwUT��|���S��k�Z�d:,�3Cf^�<w���@Ǝ3�t[�OVǔ1<���LP�
����6��Dz�bn��P��\vsn�j8�V��
0�k)l�GCcVrb�Щi#���-�Ǐo7�<"���X�]O2ջ�D���FK1�PbsZYY�I�Zӱl3K����Y�ȼ�U�1�HF���݁J-�p�Aܑ;fe�b�h�(+G��ˆÊȪA�|-�)�*����p�B���Re�Mբ+�� �5&S4�p��h[Ȭ�ܣl
c���t�=�@�.ٙ����ۈ����3�����4����0K�����H���Pm�y.ն��4	��WW��UI@ݭ�����)����n������n�W�R�nm��/@��Eh�f[�J�NT9+``���J+`�䎒w�R��7�����m�K1�J�rnXz���+t���ebu��5V4ˎl
BT���t�ܺ�gB$S�q�2l8�8Z���q��L��r�L�o~��p��7qRИv���j�5�m�K#-'�i;��X�.v������[��+Pr],��#t��ڍ�@
O.Ji������&ap4�\GbK	ّժDR�*�G�B؁���� �ܗ�R�i]͔�ǚ�n�FRun��-�A�ӮM�K��������ۼc�FثZ�����ƶ�G��AZy�
�(�����\�C5����ZG�!�X��a@́�ZX֚%�K"��� ������f=�yo/%�fe
 �InЂ]��j2+s,J�ݩBh
��T�fTR�b��I��3A,����t�Y8�eZSE7(h�� 32�Vݽ*hJ�*9C-�T6�-37j��r]i�ʂ�H0� �y�ڻݑ���O�Y4t꜀	GHb�fP�� +�;n�a	�:�s,��)�S��>��]]=���4�T���.��S��Ed��7u�2�p��mL
Y�DG�S/q�M^c�;�K��f��S��%��m�9r�
"��n�Ktj�vCus�����jي�lWPl ,QD��2m��H)�jd��q��l�ѹ�̨�(��ܳ 	�3Fj+�y���q!�FZ�q5,9�7�cXu��4.��N�����8�PB\S���LB���2��^d)( ��՚'�ŗ�#e�F�0�,ר*�n\���{6L:Z���Ú֣��4�a���8�9���W!�꥕*�mmǗ	´�cS�F�w���^
358]�3ACnU�+���I��Gv� 6��#aG�ha�o����v����
NfҦ�CkCtj+Dy���WF�] �{B�7���!J�CEe��.*�س,#���c%�f�KOA)Kb@Vn�,#a鄮��xk5�j��HѫR��/EE��+F�h��7t'$��������=�*�ժ�Lſ01���J���,q�+蠩B�/l�J\�Hne�M/�v���
�#�l[Gq$��1"���l�D��3E��9U:Ό����=�^���6��B �R���V3X��hcph�lۃ0h�
6]�[�KŹ�j�)4kN�c��k�Gp`u�o"Z�WN���v]mfh�S�����L9K!�Cm�D���-���[ugչ��<Wk2� ��8a��#��qRĜ�a���=�͸Χ��SP��R&��&�J�,f�����q�Y��%I#?��1^6�3l��ݰ�ys x���%��%�Yv����/4�@�%]$r�e�V�Ll�5f�OF*t�I0u��b�4Ç2�-���p��L��:صn�@�t-ӈɅ�̹��;�p*�6��{i��m<����{km�,�T��mL�ʙzĥ�%r�H4�E�N1N�m�;���H6��YX0M�W[	��$Qʛl�{p32^i����wCe�U1���ڷ��%��U�͌�?$̬Bif�S� *�#[f�R��������E-��"�\��N����P���.�wRB#u�h��dѺ"k"�v#�,����[�fM�W,H)f��L�y�#&��Icmd��`+i�J�Պ���Rʱ�����klFP�:��D�����Qچ	Z��KN]JѺ�#�GH?c؄ڕwAh�EԔoB�\4�C�D����l�F��j�����wIY���f��KL�0�[�݅(Yh��YƦm2Pe<6v��
�R�yt"�3Tf��n �BQ O4�a�Or��x���`*�1%�1ۋ]&�Fm�n�[�'�����C7$N](ϱ*�W���A��ƣ�qkm�9H[Œw�S�kW�����B��QYhJw�����nb��n�b������������f�p�4,��4���HC���n��Z� mZq�9L�2�ӭUo%Ip˷4GW�*��- 5�����i�eI�����F�n��,K�z�.���G	.��L��d���2�쒛N�%�(Gw���hU����@5�a���rä��3j��w&�ܻN��)0�a��R�(�m
j��0B�%:�bV�ͧZ�YIn�����5�(!XF-шUML��GD�dB<�xὥ�h��.��[�IBs1ܹ�Q,�w�ZY��/u봂��
pV`F�l_�<���D"���&[f�-�M�ҫ��E[q%wtZnS0G�G�PW�m�n�{X�:2JV9.z'/���RN�Q��� G4"�Qт��`�2�����+���r��ךnt"ƦG�&Eb��h���Ѵ4bx����R{c3���8믺]>��[�e(e�2�ڻ��`V�I���2�ŋ���j�g�����M����F먛[	T�wK�����L���
�j["��b���j�)��V�u	M�܏Nm��/�w7��ٛWO�N'��p���(J���{���%J�3X�C��lٗ4i���d�i��D=�f��ц�d�&1$cú�M͙E�2[ؾZ�'��F7��vQk6Ȱ.��0��n�]�@n�V�DK�+o{r5�7���#�H$JL�Է˽�)����T�`sq��K��iБkÂ��F�=E�� g6�"AM[2�-��������YF�ъ8�=6���ޖ�n]l*2n\cWl�4,��-����t�a9tl��fV���"jE����������
IG�Gf;���&0�Eh��Q���J�޼�[�, ��v0�kN[K*,!�賑�ɶ5���n��\y��kw�m�d�mg�C�1�.SZ�yM�ZZ�r����f�KxY�.��h�t�V�	��`X;�p�SV�C�x0)e%�!NIi��^K���`U����.�k4�F1�ͶŇ�:�^;57��e1b�j������ɂ�b��n����c8�:z�V4�gp��*Ѻ�����@Xl1d!�)���8`�fT)m�l�Z�'yW�T�L�x檔"䢡t�Ñ�&���L�v�n����n��1���O]`�M]�[x�������x �Ӡ����� $MK�j���gP�T7-�[��K�p �m
C�Vb�ө�񺺄�[���:�H�Ni�;B]�Q�X�H4:�2�T+m"��;{�o���
j���Ͷ�C�f��n,�vv��%�@%��i��M�_&�˵���z�E�X���R:*�Qzen�JYW�n�C^�L���h1�ìGr伍LL�km��f�>;#D���l��mT�zh25l,T@,���:iV5�ج��^EpSb�*I�2TY�*&��De��!�o33qm�Sm�	Ӻ�%O�����eTb�"�R
)-W��A��ӦZĥ6w0�aNn,���*5+t� ����!c[��lH�ܤљy����Y)�+\ȍ.�d�6�CcwV�6�nl/Z��m�ghФpl�q7E�NVh���o^Z&MTC�PS�#��$��彷�6�9��T.��"h��#�K���z�S�x�@4�$��^%ּ�"��X��4�Cz�rࡰR��С���z�[�a09���O*'Xc��g�� ��sZ)���$����[x��1��LT�n+�"����݄��ov��Z�/v�7m<�.�X��X��l*��`p�in~
n��O0V�r�G�`�h�(lP$\�����э�V�榜�jt��7�5����<vHL|�H�]�����dir����t'v��"��]�F�H�I��;���g���Ͷ䑾l�\�>�(�Ss1����]�K��F�H�I#�$�2Y�99'wN�S�uww9W��7%��%KK&To���&WwJ�����sM5O��J�ˠ��\��N��}���7u�}$o����>��ͽ�SV���F�}#iM�ǻ�b��l�|�x��o�K��w�srH�����I:7�Op�m�N��!i�Y_:����Zu�Fjm	/T��v�����>&�T�{�Xq��9^}�d*�_g��w���ê|8��͕����-,�NΚV��]2����Sw��
Jݖ�y:4lSZ4���s.oǪb,f[�n6�V�{|�`����,��4�va����c� p��g ����'fpS��#(���[��;!��:k[d��|q�nܿ�-�Jə>7t�����yd��.�$��c�3*wr�]l��M����K�������}]�SSOƓ��W�h�(����o*���ˢ�^���]]y��k����eX��;-�ѵ8�o��t�V]�jC��6z�m���廫剪J��𴓵��]��-Je]��gi'@VK"] |M\�R�OXd���b������@�gZ�G\��F4޶�N�ݡ�5��}�]J7: 0�S+vY�M��S��G|	2�
����H�Ո��-�+�*mn���(Mڌ��d��{u��ٝ��9��4�˽���҆亵��"l�-7�Z
�Z*�}`���C`�Ҁd;N�Ƌ���J�����p�b�	����F�[�wJ�Xr#�2�����0���̼��_r[˹k�m��];��ˮo�q���%(8q��m2�=+Uk��G^tZ�8k��얁`�V�`��@,uR��q�Ρ|E���]�����.�U,sx0�t�z��ZGtO&�4p�n��3��p,�2���YP휣��wV�;:�������dA�V�z�<6q�5uwWh��
�Ř-�K�8�e��4P�ɡV�W���Q��q*'�*��襡W=�ц�c޵e��%)2o��LT������V�#��|w:nˠ���n�ݴ���v3�:�m]�F�*�e�n�
�;��=Iq�m��DW3V<��<՛���d��ܮ�bV��»�4��yB����LlE���ol��t��q$Bt��4\�-��d͉�*�

w�"G_d������㕽\Hk���̩�����x�}igT$���L�rWp��ګ��,���R���Ө�շ�x��l�4`�/��ۣYpH{ND:��4i](wu�,,�Iz�e؍V����<�&36�-���ț,������f�|�u]"R=
 ���{�u�����3�{��rhT)�8��'K6�uz�K�)���v��ĔP�ֻ�����5y��I�M��Ղj�n�]�͇��@:�+��Ei([�puW\U�]Ψ:��X�B��S��3@j7°p�sU2k�'&�!�"^=��e`̭P\.QT���67B��
��5�6 6�Jt��2�y�bk��rnޒ�ruK�B���`Ք�����2��5�ԑ�o�=CmC���3h]��Ǘ-�;��6D��E������Z��㬬Z�;��S��k{��갽q^ǯCZ�k�X���&���l:���y�����oa[z�c����r´+�]m
�����o�v�ݵ����$�.���� ���5cYG��iz}$��F�a^�Iz<����l��Ė�\F@�Y]�S�;�:D�b��'�_Tu�V��K�,euc��o� �
;��Xpo�fv✪�Cn�Zn.r�)c�m~Ĭ�3m����6���,�Ru{���f�`\�b�U�dY6��L1dYWX�%�ab��Lk՚ro<OHyH(E�{u��9u�gg"���
�.�Щ��ɗZ]q��5�Q��"�@��#�U���lfE��q<Q�k��w4We�F��vp"��fj�O]����l��LS\W��4�ܣ/7��eHkX�§)q�xr7��]j���q��Hh������G�r�THje�j�ˏ�,]�ٰ^[���s���>q��g�ԗxD����o� ��ctWL�{�����aU.��Jz���mo=nu������.:�2]���h�"P�:��h��K��j�Hb ��^B���(�#/��ie �nKMN5�tj����Wk�l�K�x�a�t!��,�Tӱ)"�G�9���dd6*˕-�L�g~|	5'^t�6��=����V��h�/GA�;>��}��fVB�+��6��N�s�xmn��Q�s�e���WLG�b�{E�i[�Ǝ����F�ܒ�)��1o15�-w�7l�ܫ�J��Uv���K�l/M2�Y��off,��U���t� �H�2��)S�ov�=����.�4�NjVQݱ���/��#��m���oϊᝳ�ދ�jU�3|��΄���̠�6�a
y��#�{�
��M�}E7�ӻY�b���y6�U�r�b�Uү���s�]��N��;��w��yvj\/�����u���!�$
�r�ywH*;sN62ZWz=��3��\�&�C����j��6^w�Y����ڒ�Y����.u&&�:b7�Z×���H+�a�.�Œ��.H��ұ�u.Z��� �cVM�{���jun��6�au�f��i�Me�7�6͇�c�zR��
!�wc�g.t��8��;��
�}�i�����8%����g;v�[���\KQ��w\��Ojb��
���1rG
�B�S<��ڮ�X���v�p������݅2�˭'��yU���v:��S�Lt�r鷜Z�N���	�o��P�hb�,N!�y2�4j�k�K.��T���A��"(��N���P�,�t���ü'�;J�L:t*](�R�f�������}{��ʗ����u^<%<j�V(�z\Ǳ��%2��\�[���Q.�P_��I���gr��r�*�v�u��k�Vq`|�|��!N�;�5\�ׄ���%��xwV^!�Ցz�!�\�W��YK*�h�3���B������&�q5G3�L��]L�`��龜hOj�<��6�w�i��a:J��m!��%�bX1#e�Y2��ѥ|��y'{iM�c�F���`���u��]��y�R�È��X� �"x�%�C�5�L	wl�0ɴA�I����;�q^1��,���J���uK)�&[�mf>\���a�YX�������h�8���N�Z��F:��s
Aә�ok43�k�eaE���	��`��7s�Y:W]2���-���\MV���JvQ�|춧B�n1��Z�f
�E��v��D�*�0'A���FV�]��!5�{�����)���%o8��O(q�k-g0��]�˷����j�ZӨS���
X�!�Z&b�'GQ�wveZ,S[ȇ��szj=�L�J�s�{ ��d��� !��(b�R���v�4�U���ڶ�U��D�+;���*��]�ʍ<հ�;�p�p<�l=y�e�'`���_Nڻ��H�]Grݧu����F����,�g�`9�i��bJnf��+���x�k2��í�d��SA��ʕ��&]�=�Yj�-t�EP�ifaq�wn�@9p⋺W�],����t�n�4A�:�!W+w�o.�B*N���]�^�=̈́P5�Pm����D���S���u�c�8ز��Y�ۇ��+Y�s�"����sX��a8��8�1Ft��L�ĺ�R��y���Qt0�%[Σy���v�q��gEi6\]��Ԟ��u�3�-��2�R�]���lJ���x>Y��luv�2ʾٝ����3�[��S��JvӨ��&���o9k#E�9�67��fu��ǀ5��Fv.��n�����Nɜ��i��u � D��5J�ǅ��1+	��s1�4�=�xԴ�3 ��F��Π�+���]�LڤV�&s�:o���ݜ�Ћw�Ҿ�vW�,�ճ�8u�b�cw[w�"d�K�Y���SF�=�wM�İMvR�Hދ7�rs�9�T7���>�B'"����w6(9dV+wap5�^����c��q��z��0���)GLV�Ҹ� �&o�<�R�H\���_^��aU����s�g�a�<���[�����ا��x����:z���ڟ���ª=m�4�Q��Ve�
�;���l�{�=���ER��ue�ȭ��7`�q*П
i`$f�S%��X��q�n��;3$���������|�K�]���,�J�i�G=�X��(�8 ����.��
67���]�o.o�Iv�+B�$}�\C��0=���a-���As�7� ���h��8Tr�'v򂽮Cy	ϓ���X�5�WV��cٖ]��;�P1��Y��Y���ԺG-�x��=�s\�ל����;��[���)�F�n^J��a��x�����̍��%l ��۱��l-tx�-����M�X���՗
�����u���)���.37����̦��Kf��X��0�&����r��*O[:�+�����Y�l;X#+�1��c6┅f�~���v:���L7o!���bxB�sݥ�^�}��q׬T�����D��'��u�����IШ)+��]����t�J�PwSE��&���;�r�0�d:a639.u���ӧ�A�Ed�oy;�4��`pM#j�ɏ�ʹ+�`e*XG>��˳�ֺg,��J�30�*)B\��GB��s��ܖ�S��A�1�-�<T]�mm��Du3Bn8+$T��Ь�su���q�[h�7�t�#V7f��Ĳ�����b]/��/ᑒ] .��Y4�Q��h��t�]��m3f��f@���<h�mwk���I3t�RL��q��n�hF�IoM(��v�ثh][�V9k���*V ��һ�C��رN*J���WL#3Qċ��S��5u|�w�3����M�Fgr�hJ�ɪ�<9�Qל�9Vv�}��nX	|�&W�e����]��Ec��a���f�t��o|L��9m������2�Z�2t#�dvhT�{Q�!�Mk�	�6����Uҹ���ϥ6U�8�ĜTBYq��҈�-�g�ޡ���J�*��-fpٟ8�|m�:��nY]��ڧM�ʓR�-̔�nvTmGb�n�\��aL���S��t�U�s����v�&�]��ʚ7���*���S���Zb\!�)SEv��#�}l��'K�;��t�Х�����3��������Ĺ[{�Kz�H��l�Ι{��RZqc2�#��b�M����	,;�h�9$�Jg	X�I$r�"�Q2�803]F�^�@�I�tK),�b�<�+�̚�ti�z����(I}�3�2�����--E[�ɗ�#�6�\t��6��(.=e[ξ�9-�����G6��yy��Aέ�ε��nV�UЪ�n;j�b\��)?٬�� 0MQӅ^��b��u�V�xxJ��yX�ɫl��yF�5�Z�t�>d᷊��ƚދ�-DjW�h�:�:G&��0Y�f��\��F���'Wě4�SJ�&f�;���MmX�6xb����FO1���G(d�֧���a�R!%��7X���أ��r�V���Ic��VPWۻ������W�ƴ'����O����"�PN�&l��_Q����{7��
B�][%�n���w�Z"��)�HK�#5R���ՔXq��.:wf)jh�W�k.������<�A⾹�a�$^��4�JV�찆�W�Z�i��(K��y�}u+i��Gb��lJssw;�EY���4��K,&��L�M\�cA�{2����+"#&v��\�a�7f�q�YO�:ؕ	��t�[��`ٚM�Nk�����9�y���Kj5Z�[\��{2�MǖEҷ/���� �{���S!��Ok�%r��c�@��{�8�������m9�+Z��}~��^���o���4yC$y�Au���3{��gP ��pJb`Њ>)�d�Y���2�]�}�k1ڕ-��"�������� ރh_LI��n>wVL��X���o�l�ڸy	̵�^h�#�%[�Ț��\6L˜�s��N��L�ڹi4e���Do�m�A�A�'�w6k�`i���u�f�ձ�=���u���*�=�L�8:�=1���8�uU�m�C��t8r�l�9�53��ʥݵ� �+���z�f��7�i[�����n��NC�p�P���+zV]���z�᷋l�zU=v0=���*�T��w���[R=���/�-[ܢ��`P�J�r��`U��S�^w\�S�|��MK�����zZ�@�u$vZ�mj�5])�v�Z������#�vs�f��"H�wt���'���܇�/������䆡@�*���c�%s����Z>����$�G���mbp����D�����F5$�:�9g'��1oG�ƀmVӢ+�5GM�m:՛�b<ԥ�5f;�JQWd���}{ym*�(X�y�����kM�šx��m�� ��t2�b�x�Va��t�k(uueb)<Ŋ&�Y��c�jk�L�\\g�ܠ�b����8���Q0�8poQR����۹��Zz{�;P���'�Vv<ҽJ��ƊBe������a�W��sy�RX�u�H���u�jn�h#�\�U����c7����#���Ŀ�l��cz�V������/E��r��m\Ieot��(��	t���W����1mI	�MZ6Ke9�F�9Ǧ��h�p֤���6�ѵ�Q���	M_S�x�o��|��뗖�[ap�Л�K�:����;�{�<�m�2��w*�S3�Yw>�-�n�m�.�8a��h�4��V.e��;9���.,��M������G�.L�E�5�F�ݽΝV і:��'S�T�ͺ�-I=X�1���]e�5�Y�9��n�6��(�����̌��*`�3J�ܦ�g�mp��D�
�+vX��g'p6��N=+l�ּ�U�|bÖB��6S�����'Q�:�Hvp�dq�r�[N�d�;���s�8�� =" @��@�""G�D ~~o�ٙ��/3V~S�h�iQ�8�[�������so���8���S��=dZ|{Ms��h=u�w/�^�PB-lL���\�|r�sUnC�H*�,��"������%�Y)܎�s5qh����u|� J�J�;dn��c�t�O�U�Eo-�9������.����Wzֱ�XR��;V��%�J*�e����򰵔��m>�N��f�C����Z�j�(T[S �.�
��iü��v�P:���;D�m<(�N��|K�����R�%u�֥�&�-�۲�H�� k�M�L@9S��V�tY���:��3�p����!�!Đ�]�VY�R���������ft��Y��;��bc]8!�-�@��Xxζ:*��۬w}�8I�qY�V:�$<���A��+��ٱ`�D�ohl��2b.��K1~T�l8�wm�'t9hD�����k!�qh]��5]��xs�%��bKJ�*Ut͝j��թ�Ȉy���t-o^K
����,�Z��18!��pn����kT�t�ڔ�+s�P��h�HF+��f[�mv�ݵ�_W<t�@�����/��Z�u���&�*{3�6�DUcS��xiU�֒�2�ͽޛ)����M^�yӉMY8�D=�3�����'V[e�����i�DoC?Z���eF9��vј�ղ�e����e.�j�1��<����F;a�s��ҫW��:G�"���ʞ��l��\�M�+37K�3�g-c_�G�����tk,�2;�1�nwp��ge��;�[x�S+Xy�3��_|��ȺT�����M�V)�w�A���0�2�g]+�r�7w	�s�k-�<�Ӈ��P�<�\X����r>�S��7T���`ӷ�o�[�v����ul��6w`�=Z����^6�����Qt6}� �bP
��@{P� h<��f�]�Ǌ�|��:"P6F�3��(Kfx{���&��H��t/��<n��7�6�s��/�T�6�{=u�����w_*�j��n؃�z�;��{W�#�kWz�YN�8�7=]�M�Zvr�f|����U����8:��y�g�ﹳ��A��4u��o^��P�{؉����X�\�ɱ]����|Ϧ��1X�W p��u�}85���e�p	v�f��q��F���r����������h���v�d���b]�ns�5m��,nl
W����dz��|����-Z(��l�����\���
F�)�g�W~��uv���غ'��Yy��IH}Č�Y�K·2���O	��i�����פ��w����Q2 �62�M���9{u����y:�V�@���)ۜzGSu���[���G��^ZV�u����9�¢Y�v�6�VR�yA�y��¯�u�G����&Asq���d6OGV:12����r[ع��n����¸&�w�@~Ш	��W��ɘv�;���g3�ߧ��6�e�{�k9{SZx���=�gK7�����
U�_
{��G`f_�aڣ����==v�"�<�
���gt���0{���^}ڢ��8g�id�}��-r�@r�^���ٶ_�'��)-XVR���fW�W����h�TU�}��Q��V3�>3XL,j�v=[�=ݱ�9�x���P���A��>�h�7��c�i	�W�ĝ�y�d�k؜9d���RY�N��ƚ�'���YzB� )��l��ά�F%�f�Rw���2�� �o�W�=�5�C�lo��!��O���b��Y��xb��m���F;˫\�H#y�bO-�s��LoM\�H��"�|��;�Y���1b�ztyGlL~>���F�Q:��=��f�<�E��ł]��.-]%eS���ҵn��4��y�J������@{��h��->ʈ\����S�ʳ���|R�K�Q�-�=�VތGB4t~B�<��\�Cs"��:g��B�����E�ǈ� ����wn�;��1�<��@�w�Պ����7gI7P?����ZQR3zeƸ�/����g-V�gf�	�=L��[S���y]j�F$���#���+��{}I�>)���C���i0�����t��KgSB����rA|xw��񏶌��h��R�������Щ����Q�+��X$�y���"�罞����K��^�bS�2h�A>�=�~�[��0}��="�a��f��v����@�|llU��Q��8+��o��Bg;�����!���hҺ5a%ۆ�:����C���';tO>W6?y*��%�T�u�.sdoku7��+c^�[֕������SM�j7�#��+4��B�b+X�M�|�Y��C�jI��i�R�A�9<����ۻ�o��D�	)9¶,��|�w�ੋ���ׅ�u^���
��b��s������/+3���l��蛄|lb��ͧ����%^�YW��vq|��=pc��r��ᩬ��wO��$�
`���1 �;�U��\<!5�[��{O��l��}��^�1���l��CB�\+�b��l;��"u?
���b ;tV��z�ԛ�ɉ�Ro�:���۫}�����G:ö��m�&�x�(ŏ���紝h�r`����c6��{:�m���]EY�P���ݝd��x%|������H�}"�>&g�]5KA�B^��ĸ��׵���G�?�w��F=o϶5[�{YB��]\w�"٩+�Zk�X�gk	�sM�ă���,�����L<�-S�Ym�d��wl'[���a�V �ݼ�(`��wxw�q�zz�
Z<�gU������;3:>�}Z���\�9z+N��&��J�|S"��fc_�L�z��uF�`y����9i8i�f{�V�Ρ~��/���^��@=�{����-j������u;/O����~����3������Ѷ�F���#��]�OBS��]�"�IL��ﷻ��X�{���מRb�=��H�'�w�v��l���a�_��������.'VTQxLD��`����Ȕ����|�vu���L��Bf�s�?5�s�ךr���ر��Nk�C=�$���+ϥ�ʑ���M¡���j�~s<���J��3E5���g�۳w�(�{Ŝ�Y�{�g��N�h�?cG�zӷ��sŚ+q79y��[C�]��D�����\Xb���4Y%�4Nm��m�a�i�y%t��*�e�܌�p�e��z�]`�L5�y:���qU}W�n-����7�,���b�,��P�3Ph�΂�/-�F�i�A�|T(U��/�,���<GS���Uss����P�������r
��,nF����G�[���O��Z�{�>�l�O��v�zx�B��I�7���;_��xxη�3�u�
���ܱ�����w�s��yѾJ�1��0[��6�x9��Ҽ�׫�ݾ̱t����s��;�;Qi�����M��5��%JH�a�!e{��&<��l����k��}�A�����{v��x.�� 'i5[ޏ�_�^�+�����|�jN�m]����n
��K���"�:4;�+�W�q�x�.����������@�Pϝ��o�;W�onv������D\��p�[b�������Sv����=^"��T�E�����օf&7
TDy�J%�ꚳ{v
�"�({<�ư	z���b��-<b��9�lJ�(�gT��݋�ge�|�p����j|��v/̼8�[���/�8�ȍ���S��,�Z66S��/�f�����.� 8Z�Cye���KWR88p��n;�����K�J�0��%v^��/#��9G����p���^`�K/v�%��V�PM6�Wt0
�N;�9�v ���cv�`c%��Q����2�%o6^�O_<� ��d"�3l�I�ݤ`��_etb��}�����ԎJz�r� 4�q�+T|��50�a�Z��3�<�z�ޗ .E
�=�'^���s�<~C�װ�����Ȑ�Uޖ�}��Z���C�=��<k�Jŕ�K^���3��&xl�oW��Dn�ݔ��ԅr�{�^�&����+���J��_��T�o�ٳ�;��Ox;����/���ָwk�ȴ`|��Y��o\������.�1|i��u�TgU���KD[ơ�C�l�]p�����#ˉ��u^���.�⯍o���D(�)b���U��.��{V�/�R���Ő�����s��� ����.�Z��6.������g@Q��x�J�k�5ؚ`>.���Qd{�{N�a���Қ�WV��w���x�nF�h�/����禼����L��ʊ�M+>�:Wf���yREp������i�<0M�8��>�ƅE�u�pk?��n�9����jUK�^��A�o���e��qG}�x��������=��>�Yk�Z�(�KK����K ���s<n���KG2�u���Dz�sx�5mp<to�q�X/z�����v:���Z���.V�'R��k.S��x���kt$�0xN5٬�db�x���l�B�h�x5��ֽ�ڊv���M��рus�����vl{��T6��hq�;O��V�q�_��b�&N��{ˡO�]g�<��z�ʕ��� vݭ�4�?#�Kw�_�y��4S>�/W�偘E*�JU5���ftgF��Yf�P�jM7~"	�����ו��f�pP�>����O�����Ի��e!�u,MpA��h����A��O&7���q�>�3�Q�Z�;�Z{}���V/�gH}�3�ύ���D�hrU���[7g�6�.֍k�!Bg]�1t9�zõj+{.y�x�>-rIgY�T�75��f:�?������6����ZVd�U�� ���2�����|��=TG�������Dzɡam�l�u�)!�����Rh��*�R"�62�}q�6��{�3�q���rY�xj����̒�h�#��T��䢵Y�f���B������z��U��[[/7����.���*�1@��
�pMf�������VyQ���ON�O&o��;�foq]{;X����t�E��҅P�w��Z�:����xнWj͌WC`q�,#6��y��r����e���ŋ)�M�sB�j�����!�;���e�̢K{<�A5��1�Y�����[���)����z.0:0��#����uy��t�= a1;;U�;�P��]���|�zf?x���'��.�A�`P��[���rq�^I}��z�����%{g�p7��}g��!N*���hV#��_sL��VU��7��<��B`�,��f�f��ǘ�X��_/�#��=���ڧ�����n{'�|np}3{bs�+P�t��wQ��׎�ԯ3vk��z�^��\*���IAY�L�cS������.�K�\����:�WmX+Cށr;M���R<C:����Ք��t����y�H2��[��u���u-#���� w�po5Ͻ������<f�����9:
��}k*g[��7}=uh���Q�>(w�p�*�V��������j��p�t��m+�NG��c�3�^6�y�����7۞Dz,����[Z�7��9l�ԕotw>(���z0����=� ���~�r����9�[��*	u^"��pdwK:��i��Z�5�X��=~� 4��:�W��pn���H�8b�`7�U!�*6
��L���ĥ��P�;4Z�|.�(`J<+���R!��㧛��>7�T�uM̙t�wu���U��ֻM7�x���2�-���'zyE�&or1(��Q����N��}�,T�`�5���/���q��g3%[d�;�a<��z5˴NK��0�"X\���+^aTx���0V�*��r�D*߻=�I6|9篰G����3�b�c4e�!H+���;�΀�t6�{ڳ9OK� ت�X�oe�J�vm7:vM筫\�T�����x:�y�5p��6`�c��ֱ����7����]#���}}I�b\�߆q���v�֝~3���\"KwJw�/�T��:���'�WE鱈(�y��a{�F1k�����yf�^�Hv�Q�G�(R�upt�ŴJ{˦�k��Z�v>뉈��~鲰� 嫥6#�xR����/Y7Eݤʸ�9������g�abM]�1��y|�(5��*�Ʌ<���8��R��Dn:�%�۴��4R���X; �G]A�L���"�*��t*?:ˡ�C9�x��R��2�~�9��ٳ"�)�7�^ṱ�F�O��u\�J�hp>k��\�]wM`���ٵ����bѷʱ�T_�}�� �GRW<h��ko.��T�U�D�]#P�K-tw�U]1ݑ��ZnAYOS�ܾ6�9��sK�z���SS�/`����:�ws�k��ҷ��P[�AQ,Κx^��`>ֵ�j�é�uh�f�H�rԺ��K��A����h`9�gl�t���U�
��'C^mq}��caP��X��묜��]��5;����7ZĞ��Y/W���T���ؚ�{�)w1k�����~���������PoA0zx�Lo��Fw�q6��߷�yt]�x0RW�v?k`-��@^�G}>wk���r�q������/��-+���bi��{;�N1���Ӡ. �<Y2����͚8�G]9"�/d�r`�#��9y��@�tU1���{���]���h�*�&�I(~~�x=U����º�x��{�o��[�W��lh����d�e�N���t�Ue߼���wVIr���� ���/n��p��پyp*�w����ڏF�]qӾ��3s��������v�{KW��qxoy�����c��򼻏v�r.ã��lU�&k��~��{L<��f�5�?���$_���Ks9����ޤ*�hY��7���o��P��2�nkΥ�=�F��袏ԗ�R�#�A���sS�a��^A�.�vz�'���#m�&��v���I[�8���J���H�Q�s:���ږ-���V(�Yn��D�R>�p�hѮ�:�����1���mo#�J�[zﯔ��Yo������^kY�7�ћN_<��ӱ*��A��]��AsEȱ^͜5RWQW|t�<��].T��\�.���Kn�q��0Z��ں����n�Ѹ��GshtXi�)��U�#sy��γ�]B�,������#�$kN5��[�B�SP�}����@+�]�����qr .8y;�w�kpW5����l�v�b6�E�u�4:8ѥy�V����";�tj�b�fN�"���=�r2�(��2�I>����+f!@];��op[�-�Dl�;㥍Q:c���i��T�3�B&:h���2��*��H[;$�͑N�5�j�F-*ճ�1,�;v�`�CGr�5�ib�g[Ӗ�ѫo�gR��H�\"���ش�gjf���D�
�9|�:�;3���2E>2���0�h��N&������%����Y��t'����tq��-p��1L��1b[�hU�>�Z��K�tr^��o:���7Sҹ��\FZ��k#�op��Y{Y��o�GDyyD8��胅�&O�o�a�p$�F�����S��d���9��E��"2㼇�KB�w\�5:FE��ɭ�JC��ᥨ�W E��d#��s8�SZxT���]v�Yg,dqu�j�AR�D��"jMT4gN ��x1��vwwf[�c�`cGH�C�5�u]��3��v۵�e�z������^p���Үv�2���|һ'�%I$�Tmֽ��I��i�X��]ԑ�D4rn��iY�o��Xr�S����.;�Y�Vs�R7�-p�K����H�o,S�	�K�NG���]������G�p����NśS��ܯ�K+\��l�P�'X)+`�xӬI��k�uw�����_�.���{p,�;�1-r@��W�Ĕ���6�Ho5�hF��c"�D'�+�`*�1+h��C[��k��9X����EǼi�w9���i�W�\ �S4�kǑevS9��o�g!WF��l���d##���ue�ơ�Pg�NF7� ��g����CnJ�gt�;5����4�i;1VP��.1�yv�ʄ�|�F�v���u����x�΁m���4�p�l�5]��
��I�P�(� ��Sğ��y�Gԋ5�ek=�-�̰�[���}�v���ҧ|�bYa#f�t�D�%0�'�sB��n`T�;v<�O��[�{;�0Qޖ��_%w��u �F�r$
���]��]����j��ap�kc	�f=:�,�ӆo'N�d2���M]]w�k�c��P��iT�'�v;�&��W1������+��ASK��Hup�wN�Z�í
^Run�K��gH�!i�/8e�c����������QحP$w��1��L�[b��y`e�t��kAr�"��i�ȅ��l��w.��w��v���N�*.���w��7p�Qżv�	�6�e�ћ��a��K�9`;5�N�%!����ׯVd5]��f���կ�;�l����[�����q��e���7�"|����+֘����I� x�Pؙ�@"1Q�dQ�ف�.	�� I��ɚ,���aʮ�@�> �c�HF	Ⱥ$���a�� o�j{R��E������d�$���B(��{���(�d�'ԃ"��$�p0Ę �1�D�4�Di����hD���L)D#�,� x��w2<��h���?Q��_�n�_ԍ�1DB aF	�!��B m���(��R�N��ȏ�F<~0�/Z��2c�iJ�D	1�垡f��L����JDI��x��hm�_�*9�`$�)h���WsDF���<b�{������� ���c�h���~'�y� M��qa����$�0#����0����k����r�/��x0�cH��䈣�1&H�� � #��D|9�IL�lI�\b߮l�df�b��cǈ�];��">J	�"�����"�@�!A Y/S��qjk�����0>0���`|�2 �LQ�0�F	�U�J <C#��ҠQ ��:�8� �#1c`rPL@Di���I�Y�� �7VzDx�1� ;��߸��9���]���<Y�Hf4�hQ& dB/�ψ��1M�L3�E�W�Yf#�x��,�Q�E/&g�� azZ<@��&;�@��QDGb`E�0�;��}��-�-ݺ��20���֠i~��:E��Đ$LFE�(Ѣ:DYL	Z��'P@f>0�B(��0%&(��,��c�
!��l�3�2�h�2���/s������8����C"({&@�c��G}�r!R�	�-������$ɈD#�j 3di���(�@�H�<�G�3��#�∆Ѝ0��I�$����|~߬>�*s�������1����b��tb<B i/Ø�,�<P�#ڄ��j@�`qC��� >"� "0���j %	�E |`|@�D�#G�=]W�ed�{h�ۿʘ2�h�Bpum�]W��:p2V����3�4T�9<S�Yv��؛@�x17����`�U��w'WʆG:}g�u��)��{f�- �ۧ[D��.�+�N}�YGt�:	�sw5�1K'!�?l)>�P���qA.��f�*�8�{!7nnv�z��~�8�!�c���F�)(����#�B0� G�UmDY����Ig5�� !�������F� DW�� �08�hɋ#�!����� ��ƣ�@ϫ�s~�ٝc�8�QB:���!���-�1f
��@	!C08����a��4���� {���#��)�:�w�nV��f��dG�|��=⅐0�DG���0(�� Q�э����桘$	n4�(ǈ�nf4��d L'�"��`n����T
"Lq
s�Ȍ0������{镣or�w�vz4����F.�T��@��|��8���0<G�s��9+:cF�@�c�f "(��1&!����]2 F�#��Đ(� "�La�1�K,�ޮ`�N{�W�z��T�n��da��HDK@�0�T�@��(��n$ǈ�b%����DzІ~� ���C�4`Dz�i��4���� �0�Ϗ4DI ZP.�lN{ϖ�����Y�b<b6�ĥ ��`q �`a�,����1$D_��D|bd|@��D��2>1�Y~�q@���9�h��Dq、GB �r|E�T�a&3��+����ۚ����? 0��ㆌ_�S�J#H�b�@���$��,�H���0�2��!�0w�Lm�ɀg۟Z#|@D>(G���l��KFy �$d��0�7-\���:ζ}���m��1��08p�0uQb�f �& ��<c�JL�dC1(�[�0(�$�`%&��a�@D��0�D{�AJL�;�bL�@��^�f��м�DY�x��Y�$�(�� �$�0�3�q&>"�@ԙ1e��n�id}� %�bLa��f�G��4 i��Y  ��Y
���h��~��=��9���q��}�\��e�Vs��Z|�L��H����Z�Ԇ������Q�a{<�}FWyyHb=F#�ـ}���.����\�Ⱦ����@�]�oLfa8jnS�|��� GV���P��:�۬Ў��å�3�k	��'(�VӒ���\����9WL*F�X�:n2oF]�qN��z�d�.�jD����5=ݮi��?p�������4(*�Ԩ/o�� �CIS�z6��^*��������其�Y[��|vO�ӌ?{njS<�^>��c��XuUv�ίr:/-	k/�oVi��V�·�\����
�I�͌>����Y�i�)'��ஓ�n�8�ۻ��n�YC��G"���j*�e4��pHs�;��u̺�z���.��{��㰋�۳�4.n�o��]{+� ��h�>�l�z��ezY=]:,(K��zEeb���N�Z�SG�&r�b�Y�S>!�o9�CZ�1K�6Ňֶ�-�nǄ�Ǧy�V ����ݼ��z�Ջ�Sܢ�,�#��~�)�뾞"�@x��^	��Fr������s��s䩋�Yp��=d=Z*� ���hS��fW\RҾ����ǵ�-��7z�w���}�h���0c&.�\6Ub���tWK�n�r��G"�B٨��N��%�
ޙ�g�Z�W�f�������j��o�Wd;�׫kӽ�cǑ�<�3�]���6Lՙv{@Z��l��v����"D��k���n+ý�r�}2��G�w q�-A��J�յ�.%w�b���X�QvwŮ٥c:�=u��|wM�+9wf�����$U�Y��_P%��t���~�v���q��8�#�;.�6,�}Uo���~6�=~�znڭ���s�`Wg���/3M���-�0��Ŵw�� �xX�`5�<�?.b^��< (�$}�A�G-Wx���jר����c|����Dǿr�q^w�$�y�!6�3m���m/ 5[��+ֽ^"u_��_r�:%T*�^wa����t��Hq��۱������yk�*����`����l��x�&�޻=����qtD��xu�Ku<�ؾ|�=3�jz��������U�2�+���c�����@+ x�i�0�6=ôLX�����oޮBj泯bAG��0���ã���f.���)FR$ky���tvSċ>;���n��=L�h�G9}������c�Qx]s��^��Ҵ�OڊΞu�������k�Q�(x�z�WTZs{����[���yx�U`�q������{����];�3^��ұF�7iIZ<���.�YMmپ�k�;�pc�|^����������ٛ:�gx�&�W�ě�	��Z�>��*�$&���`[us�(lTCj����諸ͱdbv����̩ȭ��#��<�:�>`��*��B��n���ɑ�P�M%m��1+�1:v;����+ǵ�b��7�Y�jH��^�S���&:�d��iݭyU^*��a3W���
�\e�(�ޏ�K;�<�ڎy�V5e�=�Պ �����/<�}J���t_�B>����^�wsc��n��W�F=�9⯯����TC4�e�S2��㎳k7�~�G��t	0y�V�@��N�'�{{��@E4�:�G��s�~�Q�/S�B�]r����S����!�^�0��m�Y~bL��[w=�2�5�=��e�����6<�xc�5�`��$yI�YzVi��JL�9�t����=���-��櫻R�}�r��zXC=��B�T��S���L�#V�j$���<��Y�|8�`k�)�_R窷��HE�׏�o�ބ~n�o��m�DY%:2��|�-��O�x�B�q��g�x[�jw� b�.�9���kϜ�m��n�virq�;W���f�iۋ�����?"�q�Ǘ�J#��y�T��R�죉�U��༏�V��q�P�1���zP��9t���������{�x��aӖ���ۦ��"��������͡j�L�
��4a}eм˷��[�9>��c{�ӥŗH�d�4%����9lsF&��o�_S���h�1��-5xZ�YԶ9E���N�S��y��b���P�n���GѢn�����=�S>s��}��"����˛���3�@���l嗳ɘxBG�`z��q��z��^���_T!��Om[�AN����3^�N��o�-j~v�'o�ccy)6���Y�����c}�yK�zy��
��ʯ��ᵩ-��"<��z��5�Tq�ˀ�Ļ2��%���_� ƣ�t�m��~7g�{����m޴�����:���2�"�y96ܒ�n��������� �Yz����|u��
���h�'mw���P.�����S���_Wݪ�3�F�|+�$~;$�Ph]�}}����_y�:��u�~���������㑻��I���P��U��"u��j�_��*��=��01	�m����L��k�A��xߍ��F	a�l��?[��+�&᝵v� ��Pg^���(���5F ��p�L�Vki�����8W��v���#�[�K.�ϼ���`��gP}՚@Hp�K�\XV�z�q<���#Y���i�
��_�&B�|v�^�F/^�-���4�^�z������>��1�x���=m�����k�A�!Ν
Tn�s�X1N�r�����_d���ǈ1��k
�gZ��ۨ����-+�۶��wxn�oQ�I���]\�V���w�t��Y1�iu�:Χg:gM���Q%bq�yG�ѫ+�z�� �U�S���L�@���^���C��t+}Z��(OM�C��VzV��q7�ǳ�'�_�"J�[/���t�Զ�*|R����g40]X�hÁz�n�Y]�/���jj��7��E��L[�Gw䈄�՝^^[�=�ؽ����9����k_Ŏ�b�˖R�w�m������'�O��6o|G��V���Þ��絷��u�>�Vt�O�=z��,7ゥz�!'����&����<�gI����`���I�n�0�ַ%t�1=����m�E�xm]+�|�]{���;V5�<�=&��^�J���0M���g=ռ*��̻�z[�A�g��
��^8�/6�xsKu���}���4����OI�5�F�w��D�c���:�W�(m2�.<��U|��@�;0p�z��R��x��]�>�p���Tx�lHG�o̻�k%*sM�^q��^W(}��ǆ�k�b�~���.�N����{4s��y�)��û�f�v6������0n�m�+���s!0fO��v��4%g�w�����D>�d�I���+Z<�6{T��F�Z�7��.��S�WՓ3r�p��E�A4�I�D���-
Q���3�&�k҉�Vcx��\��y�n�*S�����#��N�J�3��{�-��j�lQ��b��m�9ܣ�ڝ��J���n:Z��o���ûS�Lz���������s�+��t���f8�����x�z�߆n��>L/>]����C;��M��]d��7WD�b���������G^o�w\���*��oKյ�j�@ro+��&�{P-��|0D��g�5L�C�/'����$o��e-�ʶ��s^�ܷsRd���x�Mx�y�:�
/PF�$'�����K2�.���j �ו���꣋��lu��f���I{�ꕃ�Æ�*����}<6�s�R.D/V�ϙζ.�{���*{��O��v.���<�<�	�]�V�W[nn�~T�]˜�L+f��hM�V��y�a~��t2���3U�r���z��m�lG��ל�58g���||3���T5��ɳp^�SOU��*�|N�q���*?'���y��崝�����;]VG�����d�'�)����m�q�˕0;|swv�:��w�l����w��Q����-�Ƽeo����*�ӳ��3�Y��H���x�]���+�������>~s�=���ޓ�g�H/�P|<���o��������2�P�t�x�O2��{��F�N�"�D.)�A����0�Q�'-�W�^Zή5 �lR���)DY@�9���<�J����x�KT�ń1��o��6���v�5�ٵ��J���(���DK��/�*�k:� ;�j�A�o%���ݵͭq�{o�/*l�&z��@�^�딴�C5j�]^���� ,��l����<�����C��5�f�$��u�_�sV�g�01��C/��s\����Uy�\T��0����^׃��<AE &����0�]��4�f������<Uݤ�ԏ+���������M�w}�|�/܆,u��H�̷��~P{����N�d-ׅ���f�;��E�Vx����ap���{�Ew��%�Hy׷�0l���oW�����3�/�-����_;�vh��X9�=}�<1߽7pI8x�tm�~Px�b��G������ɫ&�~"�?e�X�������8ZB��6����F��Jw�������"f��P(QCk^7�ZX�+��ޯ	P&
�g=��\lv0ث�ؼ[�oμ�z�<�zcL�x2<<F��y��,޳��L����H{���h������<�=:j{��:�/Vz��s܃�^]Ҥ)S�A�rz��;����&<}�V��Π�s���~���`^�^�F麼��3��AL�L=L�߸ٖ3tedʋ���+k
J�FL޼�:��e؏�s�eW^u�Zz��R���K ��w׫%.3d��#sY(���o*<����Zy��.:�Z.�����ǚ���(ݜ跹��&
y����=�q͞6	;��}{|[X3�g�z�Ћ~ո�ҷջ����B����q}��x��nϊ��OQ`Q�@�f�2{����y����?m�}�\�<��D���wOա��͜5Ti���t��+O�p2u���^nIa���zEq~����of���3��^�8ό~�W��X���w�z�WR�~j�N{G�����i�@]���Z
уޱ~����{Ȩ�>����zwm��$�n��=}���^O�S��\���Ƨ�=���������xZ�f���� jN�����.�c��sP�o����{�<��7ˈ���h�o���|���g�*|�N�����l:1</ί�oF8d({:(���ְ[�B��.������R�D���p��xڛW0%Y~�>��1���?y�kOWq������c��~�.IǱ�S��ҕ㝞A
�:'
G���̙��4�w���+�
�=���KH��'��t*�T�1e�G�;k�xYÔ�t'Cp��˺�a�6:ًq:�K�u��X�ӑ9P�7ǜ.ѕf��C�v�ckJiq����zqл��uĤ�,7�m����&�C�4���ރC����q9� 9K�aO��/)llA���Yl!�.�� FW!��B<;yq�u�{CM�)ms9ڰ�E��J�.�pj܌R��e��*qwVP�]�n���)3�p)I�ң�S��CW;͝ǳ�S�h��˙�!�l�R������f͍�hXOxH�#�m_U�S�S>舺�W�kd1o+�K9>I�s��S(�3�yGj�C�-���:�nN���E.��-E���z�B99�a+�ථ��ě@p�'�ʫD��z����(E��J�S�ڳ��C�@��9c4i�ٗ\�,��a����X��U��P}�V��(���v�8��Hv{p��j^V�1v"Pzk����5�tsɜ	1����
�V���=[�q�}��Ů��GY�6�[uc���&}ZBa�˺kԾ���33,����*9L�`��I�C2��(�0V�U�V�ƍ���U�/��2���")Ռ�����v�,��:i��q}�6%��A�L9B�N��걙i0[`L���`�q��2^��R��N�ZԖfXU�z`�
�:�+��eН�����f n�wn�C˜���cR��� ��O&���@�7q�G�;����-w�|m+���>lL����H�$INw9�wq����ۗ���(J���I�;2鄨�q���\k�\9Z�3H��)hy�Q��tY�T��!6���P���Z�8\iΨ��~�2�tv>��FLQí�\q36*�fխK]h"�K��%�QյBgj�u$:�a#o����`tx˻XܬU����E�͝H�]'>aafE�t�`��k�7[t�s���C|B���N׭�pN������	[r�]�6� �۴�1�ڛ�9\ >wg��gY�Md�K��s)ZN��J�(̝�5�3��1E;u[�7�	�q�t�G��{�gGVO�MQ��iT�Lӛ�����p�����iY��6v%�J��sy.�}t���]�G���.�#�҃���*^�S�2jV��]��l�͐Ω���R�����<f��4��u2U���u�yX�x��k�e-�a@I�/�T/e��(�����^�V%�>%D�bMdȲ��V�����w�E�{i�k�ǚ�j��Yk�;��n�{���UM����B������]�%��?֨e �;��y�&�u��[|'e��k:6�r�
��s��pP�ǈ� �͊�xnEW��	���K�*唶���K������ǥۺ!�kD��g�o2]�B��H�Q[��B��5�;$��X�6+y�Ԋ��g*{[��YW���Q�� =s��>�VXx���5NR��(���*Y4�񁹪������P�m��p�\����QR�ˋ����.u)ͺFc�[����Ԛ�M��=oWrކ.��OAOڽ|�zn��<�U�g�G�;�~f4�Օ��GhA�ߟ��}e�������=�8w�g���%Տ%v<�y]�6׎�U���o's�������L��5���S����8�+�̪�wi�u��έ���Ky�m�Y`K����w��L���xP���g��w�����r�xK�B���q�M.���w��_q�䧀vP�_x��t�o�ΫD�.�l̥��Ҁ��v3�c���UXіl�e�qyyu����,���۷��K=�.߯�Q#�s��0��L�qfܺK�ۺ�+̈W�#Zy�CG��3���o�ۼ}/���q��g��A;�xT[��w_��G�_�H�S������L��y�]�k
Ǹ�^�=����<:w��s�I�Ǐ�vI��|���]qڧsu�ʱQ�'
~O��7���\�/�|�}�Ѵ�v�֠��3�������㞻�چVuG�j��;u�#��7ݍYi��BYx�>"���O:��K{"ts���|�������s�X$��������uP _V�T�G_�H��u���LD���B���i�Q��7&�4X��h-��T8�/{��*��Y�(N��R>��e��~b{ļ���;���+�'��Ur�U���*��-T��<=/P�|4�D�=�����^���o��������h\�Ӷ�m[�}J����>�	���׏%��{�H��]%�ײe��θ+���kǾ�}�������\|1�7��y]��k֧x�ۨy�+&�D9�v����
����>�u'V��ъ��הK�;���J�U�T�����q�����+�㞛~��+��5�n�=�v�w�!~�q���n�fuz���c9�u����^<z��t���+���5�����ʂ�T4�ʐu�۔y�|���c]�C�D��>
1^�ѳ��U73n�
z�C�����ｘ�1m��QK>Oyt�*e���mKk�<��Y�]�?h���q���@W����F���*�������1*�\�$�L��#�<-X6:��J�~.�~*��YK��H�kO��,�kk�`��pA�z��k�~N*��L]�0��D���|����Yw+?~��Sn��)��,����^�	���Θ���c��gK�н�f�W��q\�f��ť���.�:-�dJΔ(�V�ѝh�6f˰Qu�|ݹoOj�Oh�ΥX���
Ȩ5�qu��,��nVݐڎfk����2�K2
J�Z�18�//��M��w>γ��6�Q�d�r�ځ�9����4%��W�g	i��T�W*统C��>��ˋl��r?'ٵ���أ�<�=���٬�����`�����	:%vV
�ct�%Z&�: <=r�����>�a��ǵ�z�����[�o�|=��a���<=������c��W'�����9�b��(Jg�ط��th=�hػ�z�蟽1|X�5�ھOӁ������|���d�{���k`ߥ�FX-�ۡk��m���3��t;���{r�yl��vһ���~�w�{|�t7�^�ۏӂ���#w��{gS� �|��v{��{6�t�~^ ��e'�0�A�=DO�}����M�p�+�r��Mfz��WoX���=�;޲�����"�F��K�{s:���OU�����m��^�Q��+q��ݞ�u����~�x��ϳ�;�i����أ�*x�`Q���3;�v=�o��#k=b[���l߅ԡ�ҧ���.�3�,��i]�	-�(M摰w%*�g!ӷ��v��mwՔ�$�[��+%3���22>�n��4��i��ۘ�dr�!-��c��������(�q�}/���Z�%%�$�H`��Ī�ua�Ν{b#��p�\cs��8oRfҭ���퉬������ju&�l�&��Ӌԫt�²��`!����{���
��`ϻۣ��2Aq���z��K��kت�U�h�B����^`�T�i������Uړ�޾�w�� �&�q�<|���������׈%Y%�`u���͏W����L{d���e�ך�����u��Uu�K�</ޏ�:�Wc�<6��Պ��r
(9�8s����� E`N�޲��xfզ �=��~K���S��JN�#�����v�2������W�(��M����q��[�R���Sq���]A�a�ԡz;���SK��ٷ�=S�Ox�c�:uz&�e
�����Su�y���{O7	�˻:;s���(犁{�N��{e�}*��>���8�L-+Îp<����K>�V.z�^S%wˇ�xu�C�ʥη7�q������a�ф����qW_Y��#�M���sm��:�<���G݉�z�s��8W�s��Oo��g؁#��t~�i�y����(��z0�J��;9��]�p��z\D�R�k]6J�k6�9�y�J0{��9�.�^I��km�*GS�^T�g�����J��U��{j�t��ƽ��j�S��Il˸��gL;g�һ�j���\���$L6Vp��n����N������;hw�ǖf�p���Ɋ�N/�_�`:���{���+b	�zgF��lu#�_��f{�������R���c��1>7�]�y']��d��ٝ��cWQJ���=���\�J��]�LU�[�O}�O�G����
N\޾.��8|4���N^���{�׼�����͟�mx���{.A�T��~(fۑ���v-������^`.�[�Z�
F��7sys5;'��Mz�g����e�V2���~-!�}�Ļ�]��#HŹ8c�{:^�x���6ssf����/
c^��۷��O��u5��_���s|]׽��(U!D�,OG��}�Ꙩ~�<������. uo��9/u��=y0zݗ�a+�o������ZT=taJW��F������y1	[�l��|��j���P����]��$��3y]OlJ��8!=ز#����>v|>ǽ_�~���E�LW�uJp=�%�������f�PU"Tq��Ř��^����}��Ћ�z4z�V��a�zT�LU}�=��y7��M¨z�S��m�UoJ�M�s��Ǭjw�%ü��a�x����hA�fzt�!�ٖY����v�f��7���l����Q2^�SZ��RL�W��D��*J����99�{CuS7�)���rzbGr���'j˦m��V{��������O��MZ�ے<l ���JN��K��rG]���\f��f�u����g�|�
�� ��q(��u���tX�/o{)?ڶ~�7�z��Kʲɜ�%�>�����=^]�����W:�$:v����y{�N�ߺyT�6Mr�����VO7��ڽP��XKܻ�7/���̺�#�oOZ�x��uFV��˚�Ů>��KYmA�k��������>9�ܨޯ�d����i�Vp�(�Yc�Jtza�ȳ�hW����v}��Í�4]p3�MT��|�]@*s7�S�q�\3�-�[W�+��`d^����X��e3��|�vt}�3����ax'R�ո�v9�Ԛ3��nc�R��k/�]w
+ʀt�Z,�ޞO޺h>��W+�n{Z._c]4��j-�ղ��'��w�X�������.�R�+ޖ���<5�[��f;	���zgBϻq�i=S;i�U������!l?��H�����V������"^G�_n(e�_w���W��v����R��c^��_��t�����,�;۳ͥ�)Jp̐���v!hz�ih���ZѢ�{�֎��ĩev�!��v@h��֮P�����i����{�-�9�`�	��)u��z;2�OMɣC[�8E���wo�NqlQ	j%�x[2wI�"���8�U��Q*�wӺ�ӫ|��u�+�Wg_Ng���clZ@m����y�~�p��ļ��%�?g%�`���|(�eϊ�"�^Y�'�w[�/u�޶!ܥ�;܅�ר_O	�$��v�<٣*�z�>�7kʺ�f5ֽ���ɮ��[3U��X�$��y��̙��{t(�@�<:��K�l��ނ���Fh���k�v/��Ze��AF��<�����a|}Ҭp>��;>����>�e��U��T]��T<���|�87�ea�~�Z�S�ʾ���jX� �"�b���][
��Sj��S�ά>��I����c:�5Ư1>y�4�̞�ϙ�� {]�jP5�W���s��bž~;t�x���������ܩ�wW�]��A�������ҷ��GW���.�Bh���τ�H������x����~{��}�a�Y����)�2@��岝���0w�H�'����_�Û�G�(T��.���W�#��sφ��o^���<�t��o\@��x�:���d�P��z����^H��g�V�n�⩃��2�%&rO�;�jX6��9B��=��.�ٲ�:om`/9we%+/yV�Gx3/f��.�J��;[�%Fp˼��Z�+�(KO{����5|��y��KK�3�tp�7 s�9��[��x]�:�B���P�����c��ً'm�}L=���~���?'ݍ=�N�>~�++}=�Z������e`���v���!�iz�T��{۰B�z�h���o=���I���}� `f�h7{]����]?jLgk����=~�y�?/kMk~;.��cS��%��x3�v�w"6#%z�z:EY����r�n��{������WzM��WJJ&+�z_�P�a����Uu�ίNS�~�� �wJ��k���`����4��{�Thvb��#��;��i��g=��=o݄K¯o�}=�ԗq�٫�ū3��q��nF�i5���_�Z���9��)�����W{�u����|)n�{�q�U�3��q�j�ӕ�u�n9�e^;�����S�Fʮ=~��k�g�`�.�Ϯ�>���
JlE���ɗ}F)�qL��u�AN�cI�>o���c�8��Ӣ�=�O7rۭ��kG�x��b�xa�^�4<|�{l��[|�f�\���]�]K+���jxv+pV�:�,��7�(�o�G��D���|B\}���m\��h�V�݊%�6������b�}uL�x��4�����/쒌Ŗ�e�����4�x��x3ߝ]�@[��;�<]v��<9�:%lc��j�r���9�֪ź�����(�ǜc3��ڞ-}�h��k��F:b�Κ�W��l٧�DB��^"��rp�VW]f� V��r��ײr��Y�H�xS�E���,�ɸ��*�g�i�:us�z�\1�HDa���ҩ���g�|m�;M�l�Ղ׹>��'7��Cx�鯯�P]����ߖ������+�x=�`Oz���4�r<i߳�����$5���oW��)����5�{a�^Z���V�\�p�쒶��ík���sr�}Xɧ�����P�2�z�OK���z��mX7\�2���=�->yɩfxx�|�!Vu��ޑ[=1'��TE�Bw������^���Fp���c�>u��l��ɒ����Uc�^Z�*������x�+=�n�<'��Uyl��wƍ��|�qk�og�,)�[��f���[K���yy(-��zf�+��O��b����}��m�?�RT����<ߚ]���
�U�TÕ�wy��׽�������{�&��L\�>�9�r�B�h�;f���X�g�v��׽�u�����v[~m�m�Ğ�++t�5uG-�tec��$C8աD�m:*�u&1b��]vR��sF�Ł5�5��P]/A%M[�Z��'%oU���P��T�Br�h�2,��B�@^�(9��k���H�7������o�/n!�y'-YZQ�����`{C5�=�Hh�<o�z�L���ux��_yw�I�:�ܺ�zǐ�<��|��g2k�ڨO��q�%��m���������':wG�����O=�v��}��"Cπ���ʍ���ݕdԉv>�������8u듾<�Lw�dZ�JT��<̠����k#�'J=o#����U� n�s}���~݆?ކ�1��Ŧ�7u,z��9���r��o�v��^��C;V�y����_�����1]x����.�
����=�ܷ�������Gk}�Y���zl������=�ٹH`��%�f�{7��i�=��7}�W�Ž�� �邹����L���Ƕ껍Or���ҼZ~�F�� �2�b/��A��܏��EW��b:&u�ܽ��>�j��z/���{��Ӝ�|K�O�A����bz{�3im���nċ�v|�-�a��~�_�QT���P�*�M�g���;��U��$�x\������c�z��hp��k��PgS\��R�Lu��ke桦} W�]k����C�#��A�4垼c��}w�G�K��ѮQm#�'Kc�mk%���P��8)p��f�V=GW-̀��@��H�����2y�gM��6��Y��
p�19��IShmu9}Av4�~W�o��y8G���UF���n'�j=�(���ld�͕��_v,i�;�wF�E�S�L0j��5���
�M���Ӧ��Oo���lnX"İ�[SD��5iw��f��7]�,<w@W��6k���76+�2�T�ڳ3�����&���S1��pC_=�qīmu�"Gke��F��;\�:�>ֺ��C6�(�fu����e�'Yir6*���l�n�t�T�VHn��qcs2�ɿ���>��ct��N�ٶ�G��A�ZأNb�|ݍm��n;9ٶ��#��\嵺nʐ,�c6�i��y�u�H�w>�Fo3c��n���o��&�&s]��a��ˡPL����Ǖ�,]�YQ-��-�0N⬗��,��5qa��K���^�K�����3L�qѰ2��ifM���,�t%�����_s����:��sʈ�5 Η��p�H�=5b4�����tz��4��}ϱֹ��}�*����٬� �[}�of��Z2�9L���w����\���oj�][��6:�p��);��"w,R����\��k�4�]i��X4�vf��Y]AnE`ͶEL����.����]q ��=�%@oP�:�*+[3�f"��p�=�t@��`��YZ�ȫ����2�s�m�u��rL6z�W.��<��,Ŵ�nZ7Cz���*���tSa�+����'j����oBvwq<qv�I];i��C_M�h��F�N�,k�;���(�Vу[�ҵ�n[��`N�t�w9�_����_v���E�cwUL��ۻN��"<�.o7Ɖ3J��}��,Z3;,�Ns���Dھ��m�O]�KM0(��B��ge_0s:��ӽ�:��]�9��7owN�)M�a��eY�m�DNAՋ�������#]"�1������&��{4�������QoS����m%'q��VdT�J���=W4��A��H�AL�ŋ��:�X=�b(4�.�WJ6��)��΢��R�_n!��9�A�^�v��v�s�V����3j�r��Qcl��'�i�[��h�2���������>7��$Cs�{��[�Z�t��L��Q�����[V-Y�+i�q�/	Am���)��3bO��x�C��74�,�j�=2��u��N8�a�b�k@If�ó���p��7W\U�'�G+��Tn!��[��m�S��<}��ː8q�.�i`��%�C���z<�eۼ=9ͭWHU������ι�M�E�+{
�LK]�Do��G��Ƅv.��ӽ��dlӰ��뭣
�*��Opa�m�H;�����V\Y�4N���(B;+�L*2���0�˺��C���U�7��GFv�yo5��ܭ�c�I�۝���/��v�lvE��,��-h��\Pϼ��������������OSP���nAN�,I]]r���L�|;�O�X�w��6��;�Ep������9�}�^������cBb9���	��j��)����q�K]���םz#���߽L�wyXےU7ȏ-U��������I8������Zڹ5^����'-����}i�gr�䨏C����<߭ߏfp�����+{F=`��C���UL�L`M� �ynO��Fw�_�_�}�G{������=��z��Q�+9J�o�����F�o���+�����>e
�uǻ+�g�����^az�8��x��ͩ����^�����q�Kǳ��T|��졁��?A�~�չ��\��5���Z�d��tu�>�;:|!�-\^���İ�ntO�g��>�c�Z���}vؠ0=�l�WY�r+�W��V�3��^���Hh�x�S�����r��`�������5\���f[w�D��<����2��get9�}B��HN������vn*~�H{/8�����q"I3�QY����'�*�*�w{}dp^�oQ;}�9I�O�3�>��m�Rf���e�z��u��w�c��	mj�D.Y.sphD5:AN=r���wN�޶Ì*���-��xm\�n����U�r���Iv��V\0s*-�J�g@�r�;�F����X�(qI}��9�Qe�d�杧��p.R�{�O���A�nv�H')l�U ��>yEoIӚ��o}�a��;���{���Ey���z圞�=��z��8�>}��՛���~7Z|軈�f6�Yg��h�~s�|�.:���W��1�B�ڲ��Da��i s�I�]]�����3�@�jҽ��=��X�O'���sn�<��G-��l��=�r�[��F/�yG�"�Ɛ��g���<����z�񃳖y_�����w�����8���-�s5��Q9��y��#���n7]}���\�ה�>>&s��۽,z�P����xv��s�tsi��"[��hr��ۣ$�!����֮���~���}7��坴�}X�Ӭ~o�%ݛ��J���<u�����-X�:�*�V���t�@3޴����������ϧ���}\�}�C/=���ȅk�>^7V�&6��[��T&�N�U���'�=�PP���`�o�c��N�{�%{.�#�p~0��>�C��n��מk}l�+EXa��#�:Vu><�.������9�+']Z���8D��W|(��gNw7���]2-Ц�\�-�,���t̻�|�	3c��%���B�M+0��B�A�6��^���t�u$ju9sz��CP(�Ї��̰N�֘J=��Q�F����=.�?N9��4�t(sk�����!�2~t���~[+�6]ax�r���ަ���Մ��M�����{y
�j潏�ܡc�1b�V��+�{7$���I��YʽS�\�X�@<�@��+��D���F�hW��w�T/|=�㾩�T�~�M����:o�GT�t[�Kxgiz��z��=�R5ڲ�����
;���}{R�9q]$C�oOE�4�<j�yݕy�{�R��
3k]{�T��gL7��(��,M�o�νH�N]}���=u�oy9���ǭV���V󏠉]Y�`�q�d����v���d�n%�'VI����	�ө0�n��N��Ŏ[���(�7G�S��r�>�
 "��V��ןT�b��W���~�?!�z����|��C�����csW�����%o��j���gWty��$���1�.�=G1������Z�8չ|:�l�=���d��]�x�^Q�u���{L��]�t_�׎�{]�n��/8w�n2�{U8���R�Z��u�!�Y�f�WS��3wR����KL�ӡ2�5�kU���9��;�f��T�+�����7��;�$���7tr���:�5[3:+�Wq�ee�e=�+I���B��0'��֜���8U���:9ϳ+H���]t>�Ц�t���A�����Ȉ$��Pq����}���8��^�x��C}�����Qk�U�@��]�w'��o�I�ܥ�s�ݙ��=F�����@'��<(���|U_z/J��uG�o4�ozOe�|���f�l�\�{�,�����}��墆��㌊ld��tO��	�]+N�1d3bO�ȟ@�n�(�����7P����B������zsWY��us^���#�G5�j�t�9�ϴԑ��soxe�~�J:�Z�ҭ���S�<�DLG��:��\���S��#ӣa�Ĭ�����}Z!��I�����'מA��+}�W�����Y�%�e�՞�[�V)�D��|Ovb�]����	�c�ظn��g��Gx�����z��;�Ԇ�M�9=D��yg��k���'�d�c��`鬁����}�Ɛ?fɽ�ԍ����-*���;}��"ؽ��g�c{�ǫ_���B�96���R���{wro�jk����D#�Ҟ�O����d*ޮ�jo��Z	SU�f�:�<B��x��B{;+��̪Y�10oH�t�6d�����ɣP��:��G��^S]6��bnU���$۾n�5���W�����q:Nմ�LRM���ϔ���I�Q��$��s� + J������V��������W���X{�^���Λ�C5F�ñ�wjWνC�[5vX�oOL]������tW�V_m���]u�Z,�U��"���� ׾6>�.P�p�m�O���}�G<=�wo������j�5������Ai��ヷc���v��qk�^��/=���aWVd83���$'�����M��"`��OX�V���N����qgٵ�=vC�[�v��l�ټ>��@�w����Ϩ
_3�]K��o>L��q���{�7���a�֖T��ݞ��v�r���T���9�	������O��F;<���� �Ω���+����~�z<��c�t�'m}+=��W�b�����<�����y�7�ބ�՞��S˭�5GO�V�2�.��Ҽ�醮����Z�~"����C4uǹ�ֺ�3�[>����+u��S��2�*E�L�X�x��(��L�#�i�:�����3�漴:����O�u��������T�CO�YL�q�巉{��7xz
�������jg/��xwbYc�J;��[z����4lP������RP�!�g��G����f����r�yψ?J�S�f<�c�+�J�]ek���>�S�J����@�Ĭ��Z2z�8�/��|�8�YO�ĖϮ�ZwƮ�{���]⹕�^Ӽ����[��,� ?rZ>��.����K�\�&�#�z�|��Cރ��7<?v@�~����ʮ�`#�O5��(h��p���ͤ[�����$��T�Ն��;Խ��:�>g�o� ���[^�x�Y��r���.��[Tn�Y��<��	����{[=K��3~����Ľ�#�z7h �3��a=VEdG�a�f/�u(Z�m�j��7��5�{y6���;آ��K[����|��o��}�_��63:��?��rZϟV���x��=�ە6�vc�ʀ�yzeJ�¹y����k���1gTG�'ڧ+���>/4ֈ�l�I�]�0v)Y��KfV__K�՜����~�s�m��������]���f�)��=������-��+�j7�ik�y]������܌�Y��A�xy���-z����o��M��u����FH�:G���lKx�B��"�ۛޖ��v��@��x���!R���u&����a��c[��,���P5..��t�r��f��ke�.F6F
��7��J����ݧ�^)c��a����q�W�'v��e1�j
�!�R�غ���e��aۺ��!��
�\�ۍ	����و#X4��:�8��>֭���_�n��xS�ݩr�E�_^\󎵳ޚ���B}ǹ�<{b����E/J$.E�s�$�C%C�yغ����H�6�}����ك��n�z�+�ɍz���˼Թ��$0p�]����YY�Ns�YK��dE��6�����W�J ����^���Hw�֕]�R�"�UC��9�[�m���j�;����������G�f�}�����r��E�3����oy^�������+p::�+����ͪ�q9���F��z߻�}��3u]�XW�i�.C�9��W�Ķ��Y��z�L>�^�2�Ն��]n�������j��㡉�v��u�Mտ��t�-��d-����!u�.@���Rqy==ꪘ�}�x�	��^���۞�F�58�Þ����Wsb�|ؽEk쯠��|ɣ�s���v�)�g�}��=��Ջ6��f������n������3_��g��t����*�w�D��6~�k��y�X~�P�hs���ј�#w�cd�c9i�'%�Z/v��p�����:�t�w3j�vp���I���з�j���y�̫�Ôbw�������w.�j�V��`RYv{4gQn�49��S�'^2�^p�ȞR���s�{f�k��A�	2s9��[<�٨�'}{���v"�»�x�W�oV辚�[�޵c	a� �s,L��?��(���­�m0����G����@�MN�P��#v�*-}��ى�v�D�M��XÖ$����uw.gn��n���rM�m�p����v)QɎ��C��/I�tv8���8 ��� �Y�β0�[�M�׆}C����1{ѷ�8�}��w^�͸7f�T��mw�e��ۺ����r�[��*���U�����'뱫禍dmJ*�3��_D���\�cX�,�����.�E���\Kd��I����y+Cݧ�m��/TF��ӝ�Т3�|�a�j{����n�ˡ��nơ���9��6��}]=V��s:���Hީ�����x�^����1'{U�p	�^\"���v��e^A�!���V�爫��K o�����a��n�&LF��h���+��!��h����r�k���}�m]{PƏ?y+�ӭ�4'$zٙ�"3�3��R��R�]��[��б��T&|U�����P���θޞ���X���L
Ob}M�~��`���,:�C�Q���/}���U���7�0�vsZ��ډ^aऺZ7��!�6^X�������t�yG26�W���M.�)����
��R��An�tQ�iӻ�G�l�ۥw]�D�G�@>�cG��BKO�����d�D%=�+���wa�,A���W�����kF �7�W]�y[��52e�-���#�[
��4I��#�a��W�5�cr�zϫ/|��<<1X����~���?R4��#�1�Sl��i�\�1�<dz!S�)T���w3��8I�&���>�w ��-m�l2�f�-�W�mS.�ګ�q�����I|rq�F(z'����Ȥ�A��9�KOL�92�f�ui��e�I�CNp��^S`S�]P�
w�;E+Ct��O��L�x�ׁ��q��-��v��'@��vH��@UC&#]�K�H���G��x\�!9k�N���@���wt=�W�]/���vF�%���)
{ � �_���7��N=wV�L�[F�x�n�k��?]�R>c7�2��3�7}9�����3Y<C"�S�(�����G|�I;�;���E�����8�n��uٖ>ps{�4T�DE���8{/mt[CC�C��y���W��
���Z�`�v�Fɯ���G�l�z�0�u�V�V�;��0���Tc×d����~"���D"��o]�=1�㘸G����p5��u6|#���ޞ��a���'�u%������oxi\�ڇ|���zs�}�97���٬�,�H�<���5�-_+�)�y�Gn���K47��usf��x4����}���'�ޒ�)i\SE����݆�nmɺ#��r�A������>��B_3��X&X��Y����+}�3b��"���`�[��xxT6L��-B>�X��,+��L9]����3�{.e��jz^���w��Y���b7�p,��.z��el�읆z�!�9w�<C��v�_�.G�OKk�j��>wQ�TZ��'zG�g���؊�.i	�S5����$ƽ����[�t����V,c7��Z����Jf�'��IG��	H��P!�����&s������,X��K�)�,�����Y0'�Iu�%�50,�W��j��\_GT�Iԍ�Y�f�̪��9�1�_��C�P���=��+�1��:�#Խ�(a��wl:1~�gcΩ���l����ꚜ�}i�`	���q�t���] �əX}2��_A���ۺ$N��}�>����]�>1]�ј�f'��v*i)9y���
�s;��D�:F�,K��}�nq�n�0<n:e���Gs�����[�S�3�������և;9S0Ϭ7��~�@x]�O�O�9�7��}�ޣ�W���iUyze;�~
�o8�oز���A��:hyϟ�"552d�-�Ȇ9�:�ŗ^�,��UnM}�2"�;h�f}*vB�G盒�a�)5���j��CU�S+i�%.شA�%赚��b�#�#�S�Y+���E�k7b�.�ۑ_S�r��!)Wx}�d<���
�m:�w5aʼ��C^e�YQ�n+	έ0�;�6�t�x3�H��1���+�w9+��΃A�{{�aOZ�)���W���7k���:ճ�J�J
���VSv��ı�q��&�S�mZ���c|�fK�e�ܤł«QP]X�j�́F(K�ڔ[9���ٗ�1q����#�%��Y����Փ����ZZ�9�i��i��{�cXv㹬�:5ܠ�ݼݒ��:�� b�[��Cɴ��s�3|ݻ�^���`�u��7����Q/�$\��Tu�����y���ࡣ��Ӻ�z�=ᵝc����6ڬ�gbR���O���+	����e�\%Ԧ���b���-��.�]9ҧ�؅L�Ϛݔs��]��h����="��ɽ��r�L�Ӆ�|[���u.��b�z�jI�8�΋.���e>���꺐���V [ĺY�P�7�������Р3�U�����zZ%�7�2o�-"檫]r�pm��h�i�b��{LTM<�2��Z;h��ŇZ�w9��
[�4��Lh+�pY�p;�4���f�T㘡�̅���pN�/�פ�����.-&����nN	q9Q����Z�[�aUʥ=�T��W�.����Q�����N��ч1`�掎k ��Iݗotl���܊ 7v�B�;��#�%n����L
��.��+���l�§e��kWx��ι��jF�B�`ޒ�)��8Ү㣨TS�u���ont���D��宫ݔ�b�&��La�n=���M�m3�]�����K"�X����D7E>�(��8�P��ڛrNۧ�znk�����Q��7�=)�S��ދ�ݳ��P���貵k8�wG���%��X,9�٨N��z����U�����˒���}]�u�PG�X���ip�B�9��s��H��Z�J��}����d��`�9�1��wO.��w��x��[K����fX!�7���� �*PI(�|�KV�f�ڎ��O-�8�4ԡ%�KsWn�,JTͫ����&u��#������[H�{RȔ�]�7C8�w���s�>L�%ʯ:�gr�q��bv�{iܹ�5#�Zu.���ΠKw۵�R��ǫB��i(M1�ó��`Ǡln����y������ز�7S��i���q�*�����ܺu��tD��}h��i]:���w�Q����F@���E҄36j��D���EQ�V�LY)j�"��a��8�� 7���jL��Ь�W�M�M�3�K:[���Uu�1B��z�����l�T��Sz(��ye=���+[�I�)��t�u*��d�K%�@R� \��Ɵ<ݸKB�1Gkw�=O�s�������Xn�u�T�n�f�Z���'a�5����|��hS�6�l�b���A-uu�u���^�}ZM��*U�NW�E>72���}{��{�һ�_/f�>�ç�P�\���=�w�L�'c�1&	0L�9�1���3)�l��ǈ�KV�t�v$(��S��;��;[��#(�z��o�F�H��f� z=���F��>�r�'���)��2a�ꓮ8�I�k����FK�,Wp�q޷-z||6��w28��٧��yyRvg9�u�_���X;S3�77-���_)z_e��kh��ܰ����0[���oe�g\��< b��UB�����[�sy.�v!������U̶�%fuy��H���sq�UF�у2x1�&�[0C�^�}�Fn��
�]A,��O�^kZș^��0��0\�i�(y����~wɁ�M�]�>o%v�9"u�~�� �����5�99t�ɞ�
!�z4|�]u�F+j�Nn�$p$�6s�;r�I�b��	�f�.�i�K�`�qݕ�����aJ�$z���vKd�s��PY���~����w�LR���=�}+�wP����ݸ�*go�;���#�3Vy��}�-w��l�^���[�v۩�sd��X���"����0���ڈ�q�e��Zk���+�)�굉�9G��ɷOR�nb9u����Yy��1�ښf@Wi�����C6G2l1��I[�v��\�c���c�U:,8��J�hDf��k�\r�8���v�Ww��J\zn,���鹴]���x��L�Q �:��@�t��{{[A��-1�vd]�5B��o!��\�	�u9^
j&Ђ���g�&}C6\�"}#T��s�n����Q��\��{�rjoTnmY����~�Si����]
cD���,ڒ0����� %yĹs[kk�>�'�Is���v��'�k���|���vxH�w�8E�2�g�Ys�i�ɡ;��G�W���4��8��h�d�#��l�y�x�TTJ�]���zp����>Yv�h��]��wcf�z8
�SP�3v���;�US�������2�t�9l<�t��4��f89b��#�R}E���kf�.n�W���%��:]�{Ӓ�$�h�y��{'�{���D�Ι��'4>숐"f���~�z�G��jU���y�%
���x)�����-9�wE��.�l�5-��9�K	ZrcX�'}{�X7(�������ȱ�B/oU�z7j	P-�D�M]��dI�\[fl6.ݶ��-D]��5��ca�ѯ2��ug��̶
������b�K*�s�6�����"�������\��(��ز�I}=a��Κ��=�d��㦍f��ɒS���&�7xX�'��b'���ƪ��#K�����\�F�J�5+:r/)��:�[S������K¸N9YQ��ܜ�=����P]֮:P�و�ԩ6�݂���bʖiRmu�űz�&�7%0��/`��޸bw}�D�f�v����K��kyݽ�s��?��nvș9�o�^���2��Ƽfe���O�]�'d����q<TT띻�8����x/h��.�[�:'�mtA�=��G�P��=�Μ𮻱h!k��ϸw[�<��DzPG2��ª�#���;�M�ʞU��<���tխ��tH�<ق�т��8˹��B��F:��m¿fnnk3��Rcf:�;�%C�.�a\Yg��v�XJn6m��fR�/ܳ�;���7�jjN܍Kͯ_�~����/#%*�s:�dfu�֊���mԐ۴��O���F���g��^P�ϱ��#�5-����U��ϖ��9�f�w�ZhfL�уH�h�]G�d�:3K�D�Kܲ�~�c�b>$��:h�J�ʽ�ĸ�#�\�şsu����-�ןN�g�[����+sj�����a�t_��R� j��s�9�����8��מn'Y���*o�Eza��/��T+���3�m����ʖd�@��/W�u�ܓ���\wy�%���ܳޯS,�E�fa;Ӝ��v��S���	�����/Ď%�n�:7��L�"�v���]�������G=����*��T+,ER�����g.hy�b#�^S�t�Ԁ�Z�؉�y�I]n��J�\��l�u��mٴ��p�ck�yI��ݔ1���i�B�{�b87��z�^�o^���A	�Wq`=�L�} ḝu�qV��sGNn�vHvK��e����)��jOY��'���(l�>���x�Ҡ3#�OI<��u;G� 5)�rk&*��fg?h۲�^�z�np��%�,��I=��E��%�o���]�pn�}����/�L9չp:�)�~�?UsS�ur�/���z�l���lEMy�]�tӤ���>��2�������[�Ѝqs+=����E���i���6���N��o�w�+���ơ�汘	ti���2b��7>��ʊ|�ض���ܢ��4�T�ș��{=]'�:v��\�u�qJ)J��2����Iסf�JFuo�\#�����ės��&^운���T�j�5��"�q#������K��hV��>��8(_�i
�54F(DhOƷ}]%�t@�;5�	�9��u�MRwꛂٮ��.k�gK��0G5OfP�}��v:���C��³�"�CT�z�2Xqbxb=����7��]��Fq]�E�Ś�y^����:<+�����z0�)�Չ�d�֊�r��޺���樲��tR��C<')�H<��Jf�	?C��G3�;9��<;G+�8`���rа����]�9�
_[�HgaQy�\�s��%gb��W[}�n$L|�`^��Ẹ3�H͇��'CH��x䘜��8/ �|�o�����2ʜS+�X�;�"��ν��7U9k�\���Q��s��'gEW7L'���jd�����*>��q���z�嵬_�eu��Q�<dY���^���s'w}-'�w���n�9w�Rn]��Ǌ�w[�[R��n"�g2�V�g��L��i-+{պ0��Gz�S���q���1�^�(�{yY���v�vsҺ'�6�i���<u{S#�G,V"=��Ei����i�������)^c����S]Y�Ʌ�V���;�{vt�3�TA�b+<��j�#����y�ސU"���n��K���;5�4�x��얹����{�X=�
 �����2{�;���z0+���Á�`�z{��
��*��^�̉�yj�Ք��G�D�j�W<�n���w*�XW�H�5��T��Mj0��^�v'71k��k����,��>�c3qw� ^�o|G��n��d�'�W�J��	�k)���}C�����Z��z��Tc�Z*Lu�,L�}��=�j���ήC�G�*ƒ���$�֜Wa�������m����,ǹ��G�LO}^4���g^���WWOpJG�.�Щ'ͿN֬
��rl:���lc����X�J��I4zU�'�w]J�.���x[����m�̕Q۝�_k�@�zdY�AI�J��vH�n�Z��7�[�����u��Ǝ_^�2�����.�T) �eb:�'�b�c�;t�C����N�ع���J*��.�펎�k��7��0��'Ly�N�L�Ҙ΋��V?3_Jql�^�9~�q��;w�ry��l���Y���_ΰ�U��YQ�1�-λ6���{��Tό�?��vㅄՠ��R׻��^GSU'j��ވ�# u�
q_{�v��{"�e�䃑;?�?;�"0�!���l%�>��u�:%�3R��6eFZ픓��Nnelcq�.�Ba���bs�� ��4�W _�xE���+�V���3W+*o�]��d���V�I���$�*�*l���D�fS`)�z�G����2����i2�ۢ}=�,e���'*�k+����3S���`U9�ᩮ\��`��v�8w&+��XJt�������n��|�ʣ��MS���N�v,���gb�]xT3�z��G�%�LL�W�X���V��4�E,�\�����5�Xy�)�Wo�	��gѨ�W�v������~�i�C���[X��&���8V��ۑ�����_յz8F�Dw�=��룳�v�ρ���f�~)�와nf�������r]aw�_`��3��Ȏ�:s0����~��U��3��nM]����^�*j>ӈ�lg7}��$�.zz���:�rYD0��-]���â����J���cb��]n�?7���Ŵ��dgs�7�v�j���751�m����6�e�F����#;5�e��Y���Ww�}k�)��L���{���܋�>����I������q��� �fW�q6ӓ�"��u8��9ߎװ/x�J�O<���oٹZo=ݱ4ن��b��
��1N�=�UmQ����A��X�/�(?|P�F^�}Ę�uO=^ڻ��w�~�=��P�mꘘ��hnȁ�\��������F.�j�^a��/�Wb��(c�j�k�vy\�b��*��s��G|�v��br�[�깨Ll�}{�����';$�7�
�o����2Ÿ�5ܲ���d�GC�3�һ��k���V����K��+�-�(�%O��`�ۘX�t�N��ZOFe�Da�G4 KTk kd*ܰ��t�/\�Q�ΦK����ŧ</�V��оU���]sW��{����8��ibZ�:"Y�w#|��O����{��]�K�ٜ��]����Y�-�{w/MFf���Y��l�dĭ%n��N�2�d!�ox��Û�Y�ò��v,g)q� �|�������n����3Ӏ�n�"��}�}�����:����:�ݮ�ЖD9؇p�d��9�&w��kD���=�ӕ5��t��+�F~��4��*r:B@��`�2�f7���0D��Z��Z�������2ϓ�c����T�:���Jѯa�,R�|�*/~C�ƭ�t�-����Nܘ`����@id��[ky��(�g+�n���f�5��Vr�yiμFT����~��Ni�l�,G����MR���7^s�t��_y���u��!h�k�� K���ں��k��B:�8��ڻ��3iP�x��I��4�g��Cj��#�8j����"ؾ7��(�=aĎ+<#�>�N���Mʎ�c�S�7��/�&V�K�������y��Ȏkt`�=�x׷���RB����7�v:���yּ�*���۾����}\�j���S��o7��ag���:���[�l�j�u�=L$��}�J̙�nc�Y ��G{��Le�G,������{�K�S���H���k�Y}�Oj.DR]ˢ��z�������*��Y��0U���Jʏ����W�54�Z�~ک�N�M>l�k}|��v���j(s���f���,Nd�*�UmH�_F�]=�;6�o����Nb�Ʈ��ʴ�o��D�1��c�T��eSxf����)���v���T�8���C=/��F�v��"Ĺɪ��Lݙ�t�I*������^e�?l��2`_\7{VU���z$�43!���: �֛���f�"k#���qᆝ��5���t��h���CY��B;='R�|N��a_f ��qƍ�<�D���u���:�*0��.��6��ws�l����Ъ
���i:½���af�A\��NrΎ��C�6w�c�V���?m�.�c͜�:$ڞ�:l��l��}�y��*1��S��`����o��:��-*��9	J'�{���o�u`�:q��'gxl��}Jo�@R篨����ƌ��>��/^P����F�GoG���'�~���O]z����t���g-�r5r�b'���{}����1sU:�B�X�2'�
���u�zS:@�/v0�<��nFϏ����`�D��2�>��F��޾Ow�[~���q6���%�fd<D���3P����v�ٺv`���&}��/���3{kww����Gs�S��%�Fn}�%�=73R�M�s������Lg���b�^U���z1e�p������q�K�Ƽ�a~$�>x>{�l̽�n�؝EAx��"�1#*���3�s�*��:�b�������B�z�'��q�$�s��ת-Ӭw�m��ډ��[gwvap���v�u����c��Sݺ�޵�or�����OPMi���WHT9/Y�
�w����f�ePsDE��_�GUA�d�����!o�!!_3{��!]%6=&U/ʽC�9�uGJmw5SǕ�L��p�C�u�"�m���g�ˇk���Y"b!�k(<�GU�F���iH��Guk�9�bE	�6�e�o�bD��t�	�e�\hǦI޲���y�s�ػ��1�:��M��̧0�g��%����N;=ِN��|�Oeޒ�b�x�*Ig.|��mL�W]�m�#d�n�dS1^u�S�<�xa��kq�S��uXf���3u�R� ��L����.�rl�qo=�jl�2��eF퍙�""|<z4��]N��i�/���v�=����ͥ����z���{=H:�4�m�۳�L.�Iy4�fQ�b{��-�s�9ɨ�N�����j=q9u ��}�x�����(o�ݲ�2#/��ܽ�z�4���;N3B�*q�Z�t�K�쥺S�t1����+*:��Ю�����̇�==�� ��ښ�&u�85[r����<&Yg�:���m�ܢ��8g��;̩�̋;[��^�L�[��;�6L8�ݟ�ExM��?���z:U���l��lF�004��Ŋ�ۇV�U��#s|�Ћ��ˬ=�~Y�ef�W�	y裡.?���ѹ��`:���߻��3z&����r��ξi��O��H-gM�;|] o����6�T"p�9AR+����^�{�.���S�|%à#gvu�,dvX؛�]"�y�N�ዿ��Gk���6Z(��,eL�&ƕڎ
罝+i:�J�c{trF�e=�h(��ʘ/&���,p����P�r��d��r��9�b>���y�'v��o�+Θr�m-o1��)�����P�팆uZ�Y[�x��2l�\ʙ2Q�V�_n��Wի��g�Q�)B�%���̏w��F�N�r����{�L�U�����rV�S
՝ik�r��{��Kf]-++GxP=�j��=�Uc.�^�}CC㪖��*�y��++�^l[3�ҕ8��zIW��!f�)Y�,j����Դ�FA��yܗQ÷Ջ]&���QR�e#��6��ӕ�V�
+����6'Zz�tvq��:���m�/\e*�J�sZ�<V�ʡupVv� v��]@,V� �cm��\���gr:mZ�a�E�@�e=H���"$�v�V~�(!0 u}Za�@�t�����2�m�r���݃\97��µ���!/mS��*u��e|�=��<d�J�b��3]B�J�&d����3�L6�7,�-�Ͷ��ܩ<�X�Ô�brIـN����]�o������i�"�9��S��
'K����2�=��[Rf�T]J��ɭ�5�&r��%����s���hً2�ti'G�bu�4] ��N����:-����NU�ٱ��l��#Ʃ�^�x��¯�^C��y�w�
>�)z]
\zE^ /_J�J��q��mvMݦ�7o8*av�v�Iֳ��쐅��d䊠�1H�	��3	Fsm%]\b�!�_�;��;xQn��p�*�����Ҷ���e�:����`DF�r,�V��w}7�B���qJun徚�1v��
Z���җ�m	C����Z���k�Tm͹)��yF.��rݯI]N�8��ĄN�P�n����z������w�ۮ�^����K��pj���;'�G��Z��w2�����h�8I��E�<�Z���ePw[aVp�:
�Y�y6G��8��y����1,} ���vά�ҹ��iYym��� H��_VL��p��^hJ�{K;�g�9����Z��t�Q&�c �����0�ouP�II92�.�;9pYwVest�QPOk6�Q��캸�F4��x��1��ʃ�^����o�z����cf�P��XT�0��nH3I�p���!>AY���I3�q_�+�.�k�!�0q�\;��OW!ۊ�-l�<��^�܊�ө+���D�@��Mb�#]ʅ������Z��N��{Y2�؟T��n	���T�M������XVj�wW�1Nd���1��+���=�G\��s(`V]<��y��S\@�Quַ���my+r�9�=)A���O5=9�ش:ů{���:U�X��+��WE��m����mV��u�c����m�j��v�"����4tpQV�j���ܼ��Jn�A�D�.�..�(�}je�����Sk�������j�ċ��<���]X�X�\����-_�b�����7I}��]I۳,�Z�N�rtV�S�kkGS�����Agv6��F�9�tR��ff!�g��=��$�wF�cc����>�q�r�m���DV�3�k�yճO�%sƼ�c5}�נN���xϯ�z{�������nD�[�)�u��D��w�c�M�}���Q٧=�*b����^M���nUGɭ%ψ���]1�.bu~���w�O��^��w]u�Z��w��P<��to�xZS�~�Y3�D��Ҝ�'��!���#'��*r�Xk���B�W�|�{v�|��yx��r��،唳u ��3x�"��F�^�D@�s��y�W[�}<y�����w��F$�l���h�}��b�w�\��ˮF����3��F	XL	��k�x��߷X����9��I��m�I̝�\lRȹ�T��yS�9��/�z����2�O���y$z�-���ͻ�K#bL��f.��=sW�X�x����ɞ�s,oDS5�+kO���yH��y��s]s����4�򗧤��#
�t+���>m^h��&�{��X�g�������~��ov�d��_�H��'~������[�=���˔���|���e͎����B�O@�Ha���y~ڼn(����"好�&��w	���S(�cAlޣ)�����x#���
)���v�uc�������A��$�%^e�-4��c*s�T�3�a]ƆuJ�+-��у���1ʐ��Yd���	ڊc����e�/_VR{����9M�n}���9����Z���tD@�sspmŬ�^�]�G�z繞���+�*�e��OS�TCs�dˇ�r��&�#,��u�s ]����r�.�W��0���{9�^�=;�B�+վ���iN��Cnb#|�'8!�9twI���^r����,v2��;c�+�={y���Ȏy|B=�lڄct���]D�r4N�˽�i�;rq�];1�b�%�)��R��
}���c���}r�N"�KI�Hϡ��P֎���=�r�j�wl�w�I ���e�[�͎�������[�{){< �T�/њz_��C����'WbQ�<��fʱ�̯w^���g�{,�e��q�������ES���}%�����=�
x����68{Ǩ ������b݈������w�0O�Q~c�gf��������7=�[�.y �cҮ#=@oL�N�̾���&���NX��y����#�=��m.���	l�F}7���b�M�UU������g�I����p=�m8<^�����|�cI`m���LY>w#�6�Q���&��Q*H�s��_Co*�b|,
X�:�a����6�t�Ė��0_��4lw�3��B+	ڽl��(�"���ƬnvrDT�r�[%obr� �U�u�.�!wwK�����l4�(SW��7�j.O`-��z����]���ٳS�X���y/V�Ѝޫ�j�hn�i7�gɻ��+kܥ�M�������CqvXZ3�>�
��O��
kz�.}v:�N痫� �wv:��K��kNx��3f�2��юx�8G�v�Ϋ�_��~�!^��-\N�gc���dW��ʜ�;>Y�]�f��;�UY=��Z�y9J��1$=/U%�&��tv��x3�P�b߬~~�����|7��K��~�ɰ�<飡��>��V顳��]y/LW�Vyh�U/*������;�c|ӵ|�;R�	���Q�y���\��W������U����=���ǫ�r���|��¯1��,���CN#~f"��g��s'4K���<c+&z@�O�]+��e�@E9�p�A;��K��=���!�-_<��g{���?	q�ݺW�e\u��'���Y�ȭ��>���V�Ь��W3ȴ��C�N�k�v����nZ�~�f��x]l�ݱ��GO�(�W>
N�m"�ī�l3�q��Ҡ��\Aw;W'��Wc\�C������ks���`i�Gh�g,m��ƹ���T�.h��h�pd'G�i�F"-aŧ�w{�gmZ�V�Y����ށX��0�� Zhud�9�Y�x�0s�mۊ������D��ݟ� vp`{�,�Ⱥ��j7<LՉ�ưOLP�f��h�ܖ.L���~�6�v�>����f"1���������:Uy-w���;b߂�*�#=/ w�E�=xj� ��;�5�L�(,}�dz����.!��mGG��CTG�l��=����|l֎yu����l��g"֮��{ZK�����G�e�.}�'5fy1��4w�zEX��'�l��쐧�}�a�S�Y��8a�Ѥ�O�=�`�w�[w�o��7ʺ��0��dUH�; 
�Yf(l-xfk�D8�Utʬ��Z�CZ���V����nr!�e��.�ˈ���f��WOuw1�l�S،���"��Ca�&�~L�2M����Ġ�z}����[���LlEi�;2���?I\�{1�����L�+��Y/����<�c��������=563�P1��ݪ���f7酼!:ǹ�Uut��o
�Fx���;\쌻�t�oe���ƶ>��ul~�(9�f
��f��>�13��רڮ�lo���Bơ7g"M.��<�
�������3�UN��q��X���6ǰ:7^8�9\wr��lpu6vӨ�R���F�T�v�m�@:����
;*�j X?V��+���M��*���B�oX�e�`��|�s�@1 ��ݶ1� ��N�Y�xY;������Um@�Nu1��'H��(.Ϻ���q����鋛��YW�u�,dEl{�b��A�;�a�M��h�KE�G?H�d�-����Ď�{�K
G��u|���T���c��)�i��U&�Զi7형Nk�(�ɹ�i�%��~�"{l\M*~�Xb�r�ߢW��' ����R�~��ȑ誯E�Ǉ*�[�5�J���b�'s��{��8wWwY�zc���"f0����9�pg��A��cJ}��\iq ֏T�3K���fN���x���zn���]��A\��䝞4�p�B�Q;�'����Vr���F��E	h�yߨ^���1{��E%O��h�^��N�=�'>ιu��K;�S�����w��t����+�U5$U4���V�Y+�}��d{��v���hy�����rhsA������{>�h5�|n1s���XY5NV���}�ܻ�{|���X��S���:�*"9��� t4���z��k����I"�*,SSy�s&wv�kL���༑r7A���D����
o��s/y
��|�uzڞ��
hI��W�S��f�v;>��;�j�}��)�5��!�6�m��o-�%`�4���r����j�K&�Ƥ�I]�AQ�=�%K=�����@�Cy�U�s!e��F�.���iIB��C�v�"��a�4�c2�I�:Ԛ�?������"sf)B��r�ѥ�`6�TMT�$�W��R�:�D�<QM]]L�{�U�ZQR\`1�9hjۖ�fέ�)[�����PN�J�*�+�Oi�V�+۾�3{�ё��������`�P ��=1����e����{�`(ΎR���\Ã��=�>
n�V;�S��_��_�<j|i���wTx���m�Q|��u����|C׏=���˽eW��R��[Sa��֊�����������EgM���Y)�*�/O��U��{��Oj2��8O@-��5�&�P�֕��1؟k�[y
"�e�֌G�W\�^@��gTUFO;��$
��ڇ+��ŞSjz���������.P�l:׳��3M��>>e�� o�޶��T�~�7r��Y��X���\�t��>�87E����Ww�L�`����.��9�e��-�셡���;t���R��7��5<�}'#0M���Ft���,wu@�ts��`)��B��{Tp�����%u���zN�;�td׏Jq��x��tgY��ܠ\**�����>���!��p n㚮��6�ͧ
��ƕG���Au�LR�Z�z� t��F��0G�lH��T�T�0�tA�6OkA��
�T����*���qޔX�t�Gm6�����Z�}tx��ó!��x�~;w��E��J���y��/w,y��Z;s���L��?]M�� �hX��-�]G%ʂ��>�{�U��V)p�5Ԝ~�ޫ���/��F�ݹ�ץI |����,_bh>��p�C�l�t���ǆ���X��\ACD�(�eKk/{.��o����{��C-y��}n������v11�0k�gX�'���FyDǊ�C:pb�޸�N8*�b�aX�͞��U�2��Q�pxG얽���x��Y�ɵ՚33 ?n��~�<_������W���M\!O�F���u�����o��Ej|�� �|#J�]-1�#��K�`���s���o��{�]�8����vp�r��1o�W���"���A���&��@)tZv���S�==��؟Z7�lN�A~���ƈ�t�{Eu�PNf��,�"ﻨ1��A;5�S��Gdi]'=�{�q=��o���fa���_������D�P1�H�x�0�w8��Le#���i{���t>;5��E?m�=$������X��t�
�*�u�D�Dr{㮌2��5~ݴ{����C��=�Ő1C�����h>N�+4U���OFLFP���=��˙�ȯ@���޺,�.l�-��gC�6Vh_ER��(t�{&�ó���lw��������2ܖ"A콰'�нnܘ�M����k�;~R�|�L��M�y�6
�FZ����o%�m��f�n��s�6�s	>�s�]�S9zv�`�2��*��;���,7���aˮ=cy?��~2�OV@1�����9v�����w}��  `W�k6���D��~#�1�eՅeR�S��}�ͤ&�o���������_{ca�^-�ʮg�T�M�~���T�"��x���Y��ꨈ���>�H�g��bϊꊰ.�vQ�]ݴ�j-��Ħ���x�r[3�}��3�n-L@1�j��^I]�k�o�k�皟�I\e���~ދn�{�����~�k\O��5Íq���,��>�u�
�*�Y�w7g�n\�e8��^)�þ�\�<�fc0OWM!nؒ�V�^==�7���Lc��ی�3]s�Y>�8�.Kxˋ*'�_'�v�o�h����z�N@��~1/^�<"T|+� o�x�Y��z�ޘޏZ��p�86ѾQ˝�!�˩c�니�u��E���D{W!c8�~,�O��iՍ[�H�i�A����P=��NS4�x�Z�o'���4/D�W3�S��sk߿(Y`.�CN�#D���ozc�ƶw�P�&x��A��MCb���m;�%�x�� 1(�S}�wTm��&�aȐ'��]K6L:�6e�E�k/ΦnT����p����������ܧo���d���+kV�'�����]�X�r��09� r�f��WW#�N��/�����wv��p���L���<�3��,�Vʷ��s�*&%���|QJ��~�w/6���±7�1�} ܩ��+L�2�ic3�Kۂ�����.y���XL$��}o9^ɝܺ
��EK�]9��K��]ٚw�з�l4Zo_N����؛�'xd�̍��q����B^�����Z��m�(�����=@`z��S�Mxqa��������"-:d��Wǳް�3�F��5xn,�f��Џwyt�����#�~����yn��K�*�[���s���#Z��i�/;�#�W��F��1��̕�B�W_��~��*N�GJy/�/�[�����=��\�ת�gzk�A.c��� OY�Q�}����ҽ��?]m�͓��s����0�Y��M�1��\G���#�ζ+� {~��<Tz'uwC�9v.#|��zs3'kF�U�M�܆�hjφr���WuT�Eؽge)7��](י���[��x�)�k����+w�ԛ�cٽ�N�=Ar=�Q��#3M�4��%K�ٍ�,�.�3�F �����}\=��^���I/%k2}�;�R�z�,N󭍯���Z+X~N��8��}_W�v�����.'<�p�cN�K���u�љ�|2d������� ^�;``쏿V��ǤJ�+�Z�*%��?,4��NѳsWxewe������)_/z*�޳�N�KI��>��2��/��D�����o7�Q7���c�� ��������b��S�=����t�Ғ�j��\���{wk#�\3�oݑȯ�E"�>5��b�$�2�;�՛Ղ	y�d��B�� 8!��#fX��,��8w�.����v+X{6�u^U��[ɳw�I�+��G�G��t�b^�_��'������q�;��l��w���d}�hGκq،�܊(�c�����8Z�����������'��.Dqe�Q�9���#��ER���`n=gu<��{`���1�#��Ԇ�b�3|����d�=�Zl���#.�����5H�=�cs8�~�׃���U��ۥ�{ã��G�fO- bZ)�1��{#�dCs����uV\{k��ۓ���)�^g��;�Mʺ�]v�TOl��Ǘ�T�G�~������T�Ȯ�ُ]Z�'�b�И�u�}kA�9a+�؛_kF�wrS�wP�*����e��U��U���r�W��ej4'W���Ж����qI��mE<Z<���Jf_.�1��s�˳1�ݍ5Wmv=�0���Ô�Qr[Λ�����ק]��@=o�>��P�H���:U��f������1���zy��L������͓�(�1&���hf,�9rs�G��N�U��e��l����y.͗ܙ�=�>�޳����'J�1{*{1Ea�{�>�|��@7��8��-��Ї�*���&f�I/{_.���{��W�GX#���K��W.ޅ���4N��GwxI��(�u  ��:�)���;I��k�!$��6k�^�ۦ�3�n�֏���(�}��y��cwr�=� ��Uu]u�6��+�/��z����ި6�|m�*3�K��˖�-���d����cEjZ_8K݆q��Cc"i�2�H��:a�y�����m=�ƶ�Bqz�����8�n�0AH��(���S7��E�V749����R���7��Oq���j:���}VQ���/��Qy+W	�t��������p����w�w}`[!uwn�n��D��&���6R��k������D­�ӛole�D�+{z(�b���mGn�������'�ϻ/p�V��F�w54��Z�M�O�	W}��,�PW5W�Er�m�3�A�s3hf���GPɫM�!v��r��sK'E�����I��zm������'��(<�ŵ�{q=�D���4j�]Esn���,Yu.��V%�I{��-gU�Ԙ¥fr�<۬��R��ȟ�'��;�>ڀ��]F����Pn��J��*lR 9wN�Ηc��r�W]���|�'x��E���R�έ��厂��zf�5�X�c�,���,�&�}C���[��L������v;%����Y0O�3��m,�p$�Ǐ�yz���7]�H��'2�f7..�'dYۼc��7B�7��b�q�r�Jr��������@wt�U]\]⾴]�N�o���M��u�.����s��^!l�/�ƒ&-2�.��s����� K�9�o�]/T�'z\�Tyܵ��N�}N�8t�"3����GP"���}\��6�ųz֎�ձӭW%&`|��꾘iŷ�<Y��tk��Kڣ�+Λ*���E���r��]f�7��,]E��c�[A`�bh�4�rd�v����[�b�_=���UZ�Oz�o������7����*[��=���Jn��Gp,��ȷ]���F�E�#��9���u:��J��#�riLZ��CL^���su�5����Y[�e��b�Q��fL��n�fT`��m+��R�����]�YI���j]���C|��]�n�K5�3%��cw#�Y�ļ%ʉ4�,��m]��i��/[},ɳU��
eep"��՝pp�j��.s�+B�����
Zw]�_?�*¸|îi@��6S��3�7u�ĭWa��� ��^�������"��p^��$����gn;�z���a��U�Ż���k@�2��"��\.��g!�±L�~|�p�2`�����R��m11���I��X�������^w��~yy<�ˠ���Y�N�S���ܪuq��ΰGou�N�x��	v	�9�泇v�#�v��<ʩ�u�W[��^>�sڻ�y!�s�-aw�B��1�k:����F����]���hø!�;A�6{���N47����ؙ1��������wz1�Dj���&;�g�tt�p�t�̦<�g�U��
��u�:4��̳�Xo|���`��e:��$L;Rv�ș��:��׺{��b��1�zUԑ���Qs��ݯg�Pי+�@��!l�am����w]�18Õ��{��ީ5Q����{ۯA9�j3.i���e��,��j��)\G���Ϟ�T�9sb�%b�7ڳp��t#^�kpn���|W��F�*/���ߝ(}���0���݉���~��~u��ɇ|xW38�h�^�]����y�yx�Yh�u���n���{ԣ�y���/d��e�ǡ0T��^��t��M�/�m����Xܲ�}"#��j܍KA#�o�0��f��D�|��H1�vs��s!�m��s��~i�������?Mx&�f�fG�v�qw�2�(�3Q�z�6Mw��I�gyx��Q�yE���X1J�`$BI�u��ڽ:i.��]8�ݕ>��,���i������D�oVݮ*;Ϸ��η�D���>�+�Kn������eu�W�!ޚ.D�挗�d�Y��\�
1�7�	���=�=�%�e�����I)u�bT�IL#��"�F�k��R��T%)��\��ڗ{���7N�ߒ��틕���h����YB�loL�r1كf�<UjH��l�K޺�"�͐ox�ϴ��*�{�F{2�5�f����z�ԫ]oOg��
}���l�8�0o���cz<.U�d�f��a��6r��rt?~�`6�������@J��N��N��S�kԱ���2��h�~u*�\ǹ�''�0�<iؿM�zΓ=��fxn��y��ּ���9Fe�����7�.�>�컈��h@��l�u�\����&���vm~s��1\�ҧx{1�&5�3����]�k �=�����򇭆�O�#�5tc������O�H헬��������4(}����n����}����ܱ���&��r��e�;L����ݒd��7[*�cuCQc��?!�{�2�˾��c�>�\�� ��	؝�����p�Kz6�T��w�Rw��X'�2��퀹4��bݨ��z ��R��M�2����.E���n�/_�}y�p������H���0j&%���0�^ 	�K�����5�B`�����8ul8����1`�=�^��87�})[�th����u�v��$H֞������ǲ��Dfm����s��Zr��G[��	��n�m�z1�U7�Rv�A�׆K�U�v[r1��h�t�n�}�7��(��cS�H�q�t4�W���<�CxҜ��3$���b��&#ϚŢ��|�΅����Y��c����?E��^9���]�5���b�k9ܶΨ��{k��p��X�N��r�F�|F��4:�#��Ð}�}ND�Ϗ	U�oݱ>�w�TA��z�\�}��b��^�T���j��W���lI]���9���ޟn@����wGE��x�+{t�9�;��^��Ȥ�z�zr����A��^��w��-�A�S:��y�ṽ3B��%+/F�d��z�w��u����D�ȍ�"w.�$%�2�uFo{v�^�D�B܉��t@��Ʉ��Ǡ��d	��'q���'�RlV��o*���M�j��Ȅ��K��&������v�0���}w����uF�{�AS��:梳#���/#��٪�]W*ڍڕS���tI���d*����]�"�[6B���M�����Чâ	�R~�w��q�^�L�&<��k2�@����mo��'w�]�АOӗ��%H�����wp|��~7�b�ȹ��L�������Tx�?�}��s��)M�գ=Q��8g�����ԫ
��I^�Q�5�½�y6����ו^�'}��X�'1w8V ���kM��;w0���wc�.A���U��lpY�K��N�%4vƷ-m�T�%�;t�ξ��/�x�k���Q����}�ѧiJ6��ZM��T����$��PWo+�x��Z����	�:fu��7"�_����aU������/f<P�B�{����*+=���ߎ�V��x�E�K�)S� �y����¡��ח�W�Io�t���&Ē�t_@�[���ޙ�T�l����1��;�=;��^�#��{��Wca+��3*��隍�*8r��� ,�I�<��:uS����ļ����:Mׯ���L �qv�g1����`𪞜A���u�dVg""C�R)�n��K����hP"�z���`���/v�:��Ox鋸��E��\������>�w�T�Ǿ��t���&MZ��pz��@�uv�u�-ne?��[���+W��F����8��;f�"[��K�f#)p���˴IQ[yX����+|�o���A�y�B|��"��w�������E:����rߣ��QR]�h���,�z���Ԧ�lU��U1W؛G�]ڃ�9��5��5^tO�L���-�.oH�r�\����5|K&
���Λ�*6|�V�М���ސGp�e+�ؤ^�g����^w�@O��](욓c��c2�r����$��j+D�X�B��33a����.ȾOV�*�V���*�5{ݟ �9�<wI�lI�W
,���l����9�"{�L����HM�u8�8�0do��Pik��`���hK���7Y��
z�;��뀅���5���زNn�5Q�Iu9w[��T�;y(ʰ���u}>�b0C�k�d�2偛`�-�Gv��<�{J��Ǝmf�z@�.z}z�G�m�]+���(�q5�2��y�On%p&�	��X����):��Mv��;쳑՗��g+ל�Hb�o�U�^�[�2i���T�]�t�mzM�]�}<��>٫V��ziN�~�k��^v�7f��꽈�aO���O�K�E�l/;�g;=cڧZ�C�Ba]�@>Ϭ�xT͚���'�;���q����t�8�<�"OW:�����$9��Ꝍ�m�>���>��U�����n�xV"�7�Mw��j��8^���L��Be���7�ɮ2|6���y�\�G�G~���k����ͣ��j���9�.�#�3f�y�2'���)q�R�Qg{֫��:gGU=�D��i��*^��l��(AWak#0��轢�Vk���]�>��OEw���<��1���Q�\�Yrs6�b\wN5�i��X|&�9�;pw�o����~i�TF+�ȇ����5�����s�U��I��9�z:kg!=�uG�cX�= ���F��LtD�!����@��Wz��^t�9{�2� "�+i�54�P�q�����qR���mW^e�}v�V��G��(x�9+ x�z)��#Yg{;�n��C����0Z��N�&Wp��@�6�if���	&�����z��9��..�v+0��;8j����;���=����Xz7���IL�����鈶�<��d�f|���72��r+Ԛ۳Zo�Q���	���՝Ug��P����+F������|=�R8fE]	�DAݪT��+�8N����$8�q��I���[)�,K�j/F�I�v�ίP#q�w?�<�����oE��s��qɗ��DA�rc�-P�NY��(3P+��ܸ���M�O�\O{|.rލ��x�u|���X�ˈ�3D�S��j6K�"M�xV��=�6��ǜ{�3��2��o=��T;�.;�fz6�ᓎ}�[����s�U9�{�Fhf��Q�ׁ\NԐ=��p]z�_\�D'Y�Cc�y���#�,����E��z7���L��_����S��7
�����|�la�W�y��V��*������C��uAe[J������s�e:N�3�'sK�l���;�J	�BIՆ3ו��7�׾�q�5U��b�8���'bo�#Ӓ�w�������:��һ�~����-�� ��5�.fb����7]���Yh�+�r����.�tl�\����U^+=¶��AX��C�{���Z2�u�T��YYhR]��3FH2�_EPW=�n0}��O}���īd$����ي�; �}{q=)��N�V�T��`\ٗ�(�C��\��.gs�q��J���ʾ���+�]�2.���K�Z]�,E���5i.��}Y�y����g)�狹��S�0D=�w���۾��3�=�O'2,��|��ߪ7I��C$�ʓ�����m�t�O^Hb{,�1~�>>�Vi8Y�%�zl�ɰ�n���[�۪9���ه�	�3\#��C�q�90'��ɫ�P��o�w����i�j�î��Ո�+W~R�qj�v=�b[��!�]2`Ll����ԉ^�V��;����8)������En(���OU_W	��Tӽ ߬���g�Q�G���<����+�у�W��/�ۄ4��A�S���.=԰Ec��R��"�1�ǣ���=�ι�v�`�{������\x��g�����91�Ҫ�>Մ�6��Q{9zhpys�������շ�1 ��G�1��SٜK���c�g���o�C�{���ԟ����s�\�]�_�DOJ޸��NKk���=��d	f��ϡ��[q�������s��	�9�˼J8�e����v(�}�M� ��<�����D�,ķۈ�6�Y��:H�K/��{��Gqǈ��۞x�,�7��	��ޝ���^�Xb�>d&Wq���ШWr�j�[9��@v�^�t#�q��K^
y܌���4J�Ⱥ�/.���e,7���]��O��ڳo5nU�R�d���;8��XA����GX���8�R�,���omB݋�㢝`tz�WM=�'R��_�u�ߊ�U�#֭d��˰�?{sG��?lsN�Wv�J��9ܭ�c\k�yP��H��2���r_CΔ��#T�Y��i�#�¹������a�[k����l�9r>����#�����w�{�74W^5ie�F�oٮ?��Y ?kBW�|��.�3�Զ7���.�)��{���=<�]^��f�b���9^ �~֜�C�O��q뺥T�v�vn�.���w��}N�@�T�Ig�����x7��1؁�T��׮��OA}r�<��y��,���kb�咲��z��B8ؾQv��q~5��Ò,�	��x��?�����z&�g1 ��Hc�;�k�l��tl�I֚��V�z��N~��y�T��	��#G�dMl-�[��`wT���4���	�u:,ϖt��JL��.��w-Ģ߬��O\�]
@�T&�)�z
�g����-z9O_N�Ȭ����R'��Z�x��窨�s��c+�1\��)�|5�A��!C�+�=�����+ dw����8%�{���[Y�s^�YN[��+������8��b"�����Q}X&".�y��w�;/a<�zp=��m&N�*-�Rx�4P�{�S�P`,`��U�3����M�KwN�O,�zQ�>ǵԯ����{��}�zb��)�(Y3�w��p���x�����Q��-ݳGn�.��w��.�w)�|Z�[�]pDd<�3���n��Mϴ���o��ۻ��TZ�b����F�q㦠ߎ̎/�&<��bo��)5=yt<�󍜫t�l;�}3�T^�Op��#'�_D:�E�>ghr.�ٱ���M���P������y�I��aB�B��ƹ"�O���>}�Dw.�/gD��{��#v폏��pS%uNUh�����G�4�'&d����V1�Q�b���XO2���l�ڤ�:�h�ݺ�*z���u��y�X�9,�jb�����=Ye��\�C!�Z�6���]d;�\ͅ7�m_Ï��$L������z���K?f��~d|�����i��{�ի��;��'z�1F��[U2e��zw�0��8-7=")Z]F���:���2�y�>����3/*P 5Yx�Qa��V
��eJ�;�u5�!?>���Ô?'SC�-��l����Wx�~?i���؊y���T�qF��s����c��Ek��SC�^�I4z/���;�Qkͥ!k��{S�}�ɿ��}t��?,�8ӝ&a��>3B�S�b��\K= �O�u"\����:T�<�3���15���Zs�a�7y>սw���-10���E�W!��i>ug���Gk.���c(���-l�Q��s��	]*�Qu����c�m=m:�zD�jq��\�C���������^`��ux�gF͹��d����Gq9ݺ��j�3������Z�c;�>VZ�%�U�o�����T.{g�c'�rؤ�K��&�`��6^X�C���=Q-?j�U�֍NR����5̾�iV��n^I#�K�4T�Q7�,!dw�<U��7�*b.ߌE��Q"�=4]<1�����z���{�Ր��1���q�~�C�H۟F�i�>��K�Qi#��Ї������с!��
�x�ܑv��N��)�q��;��;a?H�**��F$S2��2/���鈮���>�yV�TCէ<�DFsǌ����|�p�k�5�C��_4RQ��껒w�OX^�n��@f`�=[��Ed��O�3�^�\V��B8>�ѹ��f��Mfd��U](-�|�ס��.�:Κ��My�c����������e.��O���T�5o2*�f��Q���K����%���6y�y�K>�>�`8|��m����G{`@d�ep4m��=V��07?A��}�SZB�~���������4���^�BG(z�t|�&sٔ��7�m����S�,���|j�{r�v��xyF�a��}K�M
�{
��j��Db�yϒ������`���K�o_�pK�:x�J���Gl&�H�՘��DZ��lY�cH��q��.��;c�Q�U��d�׈�����݉\��XK76�p��Ш��F��l��V�ңMX����j����D:�>m-�@:m^���so������sG^C�9�n)-�7F��\9T"����^j�>2�e�YfJ�ܐ��K����Wq\P�ߥ�KM){�[0�V7ևwU�a���d�����Tho^C6��=���ĶQt�n�1�y��Ζ2^/���`r�˺Mi�vE�ۿA`�J2��9��*4��&!W��l#��۩b168m*�+��O��e�r��3U�]�����t����l�Jj����	����F���p��|�*j��ڛ��v�o
�Ƿ��8�q#f8z���;V]�oa�8zEmi����{�Jk����@4U;]�3���������E3t3-sHۺ4K�ˏ7j��tĞX�����E'�c�p��O'f�5AXX59:n,\oa|:��#Z3��{۪e	ܵۏ-�|
�Zmv�����ѭe�t����s��;a;ˑC!��f�ܱ'���
Z�J�t����/�Q<%SN�o�i������-D�d�Yt�[�y�fsa'cy
�\�
l+���h�r�=�Ba��银�tͰ���
��(��|��ju��;�"��'�iKA�N([|�lJ��<�\�-9��@t�Rʼ���^�nZ �Ҙ��[v�һ�.jh�'q�Id�tZ�s�7�ؽ.� 7N��0 	u�epo)*}���I\�!�t���L�y&�>T��2%�zY$���!�0�ŵr��X�}�ƻ�s�8C}w9�,�p�ɲ�Z�E�b
�u��t	��Kl�B��.�7kl�c���]�j.e���Vi9Ef�� ��g-��%D�Lt�s�fGJQE+ҵ�0um3z��+%u�ՋOƾ�;Q�,���*��;E3��8U��\�[s�أֹft�AsU��n�^Kǧn<��u�i3/���(;��DYͲ��ػ�37>cz^��v��X�wg9f�SxU�9�J	�c/� $o��� Y|�d`˂��A�8Uv�I��j����[N�cq*�P��U����،�[�Z��}[��b��p&w]Jr���:�rS����������Y�n>����L<6S�OPٌeY�/@|0��u���{���3�>�:b�u�[�D�̚���ɨ���1f�W���ҹS����Aظdtw�T�����;������:�Z:[�˸��پ6�`�l�B�M��'L���Iy�6e*
�Vrwi�j� szK�ld@�Ơ�/����l�6�� �yԟ6��D��K���	�(�,
\SC�Rg{*ч�l�R%vR�^�ދ
��f�d'"�Wg��ܧ�D�j�����}3z]FQ�I�w��ݺl/^)�7³bT�5zĀ;��+����P�}(Y�U�	�[|L/�(��uK�lc�F�������'Q�Ѓ[3G�G'7Gc4 N�P�juMиmb��6�0ܱ�Q'N����[q	�]v�ռ���n��ݷrlCй�Zt��R$��]S�ј9�˵NF����Tu�ؠ�Q���\�)9ok'q��_�}o!����,���n��U��v+��4���w�qrc����tS"f���7���TQ��]`�[>>ؚ�Ʈ�.�Vk�.&U�� ��;�Y~VZ��Kɮ����Sc���ۚ��@>�lU��Tj�gD8�a���� G8Q;	�T@�`��ğ�h�\"ދͮ�,�O.�O�$���fn}����"b��!ڍ����=�gú�*s�w$f��EW��O����������tN�r/��d^l+�uh���9t��J}�X㵷9��i��������1����cf�_�1��V/w�wJ�����\$�͹_t�n�ii��9;C�؀��LETg%,�uR|�I������zk->y��C���u
��+��$ud:i��\f^tg����g������O����gN���!��[nm8��mpT����Љ��{��Y�l�3b-�X�:,Y�.F��;D����?x�^{~k�_}�YZ�&�z��k� �x���߳+5e�O����7���\���o~��-5��:�Do-]l �~c����̹�<�""�'��&z֎C�R�J�=G;����M�D�#Asaӱ�s��x�Դp��Ю���^�2��p�9f�w��l\*���뾊Q
{%�R��ח��\n�g����m��{����lx��V�S�w"Q�l���g�����OvO�3�|��vD,];��5�5Smج'��E�~^��W|�K5��4�K�l��W�厱��}'{���}ڡ�ll����P�뱶t���OW��<�b-}~~qto=��M�%�F�ݫ;��4�WM<$�T�W�kf�c���^��as��f�.���>��P<Ϫ����d%�J�����BT����<��e�Υ'��t�GvUD\��Wx��Y���2���X�,Q�yǢn��;�[7����ݹ�D�#rD����G<�+4�^����66��/_X�������gO��w���+� �q���8�~Yox��lg�l�S�`�N���#��G/�z'���]�m��7=���#3��J���f�ոꭕ�̙��y�����m������D/d}���],�y�������@8������9�>w9>qR���;�5���r�U���8�h����O�]Մ2wO����S/Ϛ�s<#�kпq��c2=��.&�K�Q8�wW�n����6>�Y�l��d3'zS�x.���tj}Xȉ�ޙ�;<`�la�m��n18�]7�w;#]�`s��ݼ;n��Y�]Ʊ�!�EN�t;t�#<�K�'�{Z3f:i���f�J�Y˜��`�Zr����D*�A�W	����wAX�z ��r��]�����םҔ70Ҁfݗ���Y�R��e�(��[�CL0�$w+8�$u���:wNG�h�N�87�q���5��^�MOU�\�EK��R�b"�]'k��ۧ}���SYE�����D�-WD��C=�t�Ļ|�]S�v:�*�%o�+D��`�&^ǆx;h�K�k{�/�Og�G����һ&p�{;�(�%���������������LF`�ޘ02�T�ѻ�?�?��1�:�����Ֆ3	�t��GZ��bo����tV�I�� f�~>�/��ё�{���W,>�������,�g�bKX]ÔM����nG;&�7H��)#[��mo���(J�	sۺ���̺��W�������m�֘���x���Y�U!����X	��&��� R��Ž�)��Fר��e�F�c5��;ܱl^҅��.�^�3ٗ��wEc!9��{�>���1��.i������[{�뺸��~3�Ïv�t�',Nv�L�=y�&f�kV��1]>UO�^Ȃ&+�f���W�8)�ڥE|ᘖVץ��N[�����~)��n��sT��;��P$�#W��c2�=�Y�i�z�9�jۯ1�,UcJ!�ɞ��(։��*'c�7�rx�����C�%�8p�9J�l>�����ո2T�2��ԏ��C]��E��XxpLc� �2��$�-L�6�N��]Xu�T'_>����V�k�F�+��Cֆ7eY�M����~w���<S����#Ǘ;7�^u���xH�+pVv!�)Պ�(M��V����!j5�!{(�s9��H�����5�u�@�t�;���l�'f{O�.ř���e�ti[6`d\��f<jW,�:�۔����e�i:�G�N�MFz�wّ����J���)lﻸ���z����.���t�%T��Es��X:� �i�qbv�=2ϲ+=+USy�+L�S<f���<C�pu'���^�MT]�:3��%��C{�~�S���D} ���`�n��&�8���lb����؟������Y7%Fvj���9֪Y�~�S��hL����z��.�n���TÚ�,���iL#Q��|"$K��XFVd�Dp�{���U��h�+�>�{�{�뺭7׺����骠���2O��;�&;bfj,?(�"���тci$W+6��d��)�[U�{�k����Ci��np��'�0Wl�g*ƿ:�7쿄xp�:B���1V�g�a�@�E3RQ%F���݅<B��]��>���}���8CӍѯq��Uh�[b}Ô��7[u�C5m�#���q��:YOf�ZA�����p���׊��z���LLNe{�2�D�N��U���f�mS9�	5im
k�f`(��V�g�R��w8q�bѤd��֪}f��8��w�De���-�l�wv1�x]|��.2�mk�?4y;0�è��p3��Vc}��$�ȟ-:��YY�W[]�Tɹ#��A�_����p��U�>��13�n�h�_}�=W%�p��2�x'�/���QV�8��2�j�w�v�lo|�)���lߙ��o=ڨ��b+_�z�A��vq�����ǔ7�%x�:����x�3ȥ�^��Q����B��� q]8zg�;��B�;gB�}�\��{_�K���
s�w"s�Frn��������w��3'�{�{�fd�ߢ�}�c�h���.�z.Eè�4�1���5�4T��ܽ��ϓjcA7
���(�1�6&y	�Yx;�\Uh��{��&��t���ƥ,�ۚ���Fh��d�'(Eϧ��#2���3�.,
����l�p�Z���R���S�\6�>���^���ԆMB�Y�tԗ��&{1�� lu8-|�Uq��ذ�G��"��.
�n���=���1y�<Q�۾�A��CZr������o)�`�@�P}���6>آ�l
��k�fi�OS��.}�����9s��71�󏞍��4�;+>wVE�'�>�Ԇ��Z�Xٗ�W�w��g��.�I�1��~��C��qU�5�|�EK��9��_W����瞏b{��C�M����ݖ��k��jykhV�3A��v/�Cu��Թ��&�@e`��k�:̽ǯc���LggZ��C7;�������_g\8�U�ʫ�w5�B�=��ʏ�:2���8h���Ӕ^�bw9��;�)w4��6��h��gI�a����2������'�j�����´W��(:Nx�܅�}�X�/��i]�﹟�$z�iI�gV��f��ګ�'��b�Ɔ�c�	�f"�n���i��l�>�YB����"��ߜx���:n�K�F��M=:m�)mⳏ:+3���%�]F�˕�(��#6�VQ�I=�=�=�5{swc4(�7�yٷ�r�!�X�ŀ�v!o	<�3�Kڂ�p��Ke���i?\(
v~k ��^���щ��v^��mv�.]o՞{�-������ȓ�6vb;�E�Aȗ�:~��+ezH���_r{�5lv�}�*S\ţ����}�~Ό���e�!EsP,��ׄ�� �]�9���t��]�M���Vꁕ�c��e��T��)�J$��J����<��v1@N�K�����v��=K�}�J���,o�`��;��k�}X��&|��ѷ���|�7Id���k��r;|�����S�_��y繁�Χ����u�;�m�w��~�����wH],���.�\|&;�����M�}��f�̂l�	C�DB�f�UV��;=Ѱ��U��AYY="��C��B{C�o=ƀ�����R�߯}ћB����evkP�۬�%^�]��f���So�]�A�U��х�ve9���	��2b��b�w���]��o	��{l�y�$��u˄
�[V'I������IV)�`�T%���j��#�s1.3j��ws@�!�2C�P�='����y��������ہ;
e�5���=˸��Q�ʯ\� \rml�"w׸�������O�ӥ@�����<!_�h�oT�����G�t��j����A��o��fQh����M��VP��v?bJ9�\b��`ס=3�:�z'˜�ɻC�ܻ/Ez�����=>�[R{�}+��y���lG��g�!�mC��d�ˬ�y;�P�Ӫ�,k��){��[�b����9]z���z>��]��6J߼/�q�-�o��v��1��6�QI�>�KbWW�=��r���)��_U����ا1�p��/]G��9u���`o�S`P;z�rQ��k�4��9H��D�����~Ww}�ӂ��!�kFCȓMT��^|���zG�H�0	~���%�u�S����U%�b�yxn;���ڝj���|<���M��v%��G���gq�)�=�[��>,׷`�����䘸v�!G{vw���Z���;��~�Y�V���>�/t�4u\xR!z��qB�aϷޯ�+�r�h}u3Fcί{�c#g��Ԧx1�&st�%��7n{�-}U�{u&�n��;��_�S�~fP��Zg�U��#��>h�l�{n�)c��C���a�@+����yuf^<���}�Emkb�w0�QLI�pA�?N�	tWm�v__o>��¼`�AD��H3�c����|�̮�b�G�6�)�%dg]�Gx8��('�s7ok��E�4m{�$P=^�t���\gg���[�o�u\oe\�q�kҞu�����D�55o����~1i{�n�������"�t�8ؐ��R�/����U_o�{��WS\^v�=�cK�OPu�̈́��6
-�������Ԉ�6~׳(��%gy2���v}��[�ϕ`#��A5���l�� y���R��~s2�5��9�%A�.�B�S�O���������i��K	�ZdFs�����)�)� Y�\���jq�.[�)N#�>��Q����˥2�j����}���05Dw��A�=<ƈ�k����F�R�a�I�|:D���#���]��=�<��[�WV{��e{=b`]�|�q^�-��[K�
�%}w<s�Z�u���vz0��'ǲ'��U�uS�^]�:�N�Wq��3�fJ�m��K1z�j��h>�T$�A~\}�/�O��{��*�<Hr.�bz]g�ɉ��u��J\Α9�:�Nk�S��*���9H��s����'g@dx��.��3-�e��;ds��Z� .��G>�7Y�}�L�FZ�q�߬��Y���=��O\�_���9��ڹ\5Ո
'��n�*�S��X�d�[̵�}�����TUʝ��m\g8N �9WY���bj��	�;v5�v	�4�%;^�[̤IN���Л{���B��to��\�9�ͧ%��]��Q�[Zo:�u�_NZu;�Q^��~Uw�~mz�(fA�����b�U�W<���xd`����s��y&$��V��ߢG��{���uJͤ�6/)�F.��ch��4K�b�b���&q��:��vl��8��A��c�R��t�։Y����ܖ/E���v���n��~��^Oo_޺��%��R�8qV��빪�O+�gp�۹x�VL�E�'�kF�T���̅�=��Ō�f�]����Z��� �_|�G���D0�^C��w�x�R+7	e��H�mt�h��G#���)�h�����s�;�4:��V�_�
��(� �y���N�Bq������<"=XG3s�\��X��W�)'�EP��Wܩ���Ǽ�B|'����feR>܌�g���f�kz�kZ~�X`X�^��Y>�E�'����I_��@�qv|EW
�]<�/�o��:���=���k���'.�2�����NO^�X�b}�y��n_�ë���z6��k�UcϢ+"��jPt'k��}Ƚ��	������
�>��d��}Q.wGD�32Fe?j�o��"�>�=�h������z����ݣ�qxW����QZ{2��ɭ��{�z���L/l��"�%Ӫ�9@b\^T4Eק	}ީ�Ufy��j�h�p�2��0�:����������/ǩM����]	m��S,�ZC�ܫS;��K�}�nTSW@؎r���e ��FݽRWd��0�*֟!X�B�[�i5�=y���w�#v������kkK�P�����@�zYn>pv�k;������ӓ���I�b�#v��t	���#�i!?b>�u��3G׫'6�f��.2,G�FHݻɽ�j��x8�F́�)�U�&��x�|��u�ǆ���G��ь����&k7P�讻�M���z0�]1f������QQ킮C��e��l�I`;�ъ���s�5Q͐ru{2�NXԾ*��c�}�����M�c��.��	�7���r-�n�_p��۞�{H������Qos}۰��z���\R�2o-��n�.�r�_�Y��b�$������t�Ǎ<�!�?8ePR�:��{8.������+���E^�y��ú��aK>� 4/_�|�B*c/C�8�)�5���IQ=�t�-TONE�g�>�B��FNW��ʥ[��e�:�z]�c��_�E��)��|{�1H��)`��}~,/=�}��{C�^>	^=BߐS�[�Ͻ︀k)dѢ.�k�_R�lU�95"��ӷ���� SU�$�kz9��ĩ�3{�g�K�e�5��wkTn��4S��NF�}��6����_7�i���!���~��ƀo!H)�1�����Q軪���=ݭ�EC�p���Bg��%�P�ca��ƹ�躍璣WL�:���2��~���}��t5�V�Ji��v�tV��x{�^�W���[��i�y�Ua��4;�d��9���*c�mv�*ë�I[�tꝅ� �כ���:mI�l�|�kn1dTv�+����@rvI�6�����:&7��/Cm����9R�>�*�����ׯ��k�L��BL��h1R^��5>7��=�3T�"͙G�)Q{���م�.��;6�K/�����ÀsR��Z�t
��[�M�P���:]S��5��ݽ�W� �t�}\t��B�
L��J/�ӷ\d\aq�ZO_,z�WX�(�c���2�ˎ�V�}Ս�noAX�3ٞS���q�}J�Yc���s�thiI�+$�u�"���(v�#��6�+l��Bm�peA\�0+��@&д�bR6��!�,�.L�K7�5r�I���&��E����Ȳ�K�v#!<m�>X�Z]S��»2�J�q����[]DpGfeGW��{���w����ԅ�	&����>���.A��t�<��QA����H�5m��,�u��5�z�Kt�j
|�-Ǫd�����hJ����ZΈݽ��o5�����(�m�yFF��37��ӃJ���ͧ���e�v��N0��޸��;�(.�����B�k����9lk�{��f���C)Y���IE}BՌ��+���ui
,��r���	��^U�&)N��j��U�{���q��H�C�q�wL�Zo�."9�ξÁ�F��C++q,��o��;qpp�V$wk;�F$ͨbD� ��[��2p�������8S�e��걛�)F�N��m�LY���x &q�+{-(�[w�PKe1hb��/��-�_V*p�p;Ɇ+�����h���h��]��1g�8����n��+zP)f��ҕ�IAʴ!�7��TA�����r�ݍ�Ʒ�Jiv���OvN�NI�ࠐ��Ljۊ��:1��p���A�� ������;E�Z�G�ˤ똅��K���^;u��*���U�|5ɋ�X�kL�x�ý�_wGL4�g1��X׶2S{N�E�ȕ���k�=�Ei�ݱ���gS���<bİ��rV���4�z�G��(�:K��"�U\�y��rC��l�L��t8�=��FWhm�/3��޾Ͳ���޻��5�
Lz0*2�}=[�*�[�7]�"���\y�9�VM�+n�+k�\{�꽡9tL�&������!۸kxl��bw�xY�R�����j��������u�s#tk+���c��q��� �e�X�D�Z/Ua���8��K�<�YV�j�e	9�]{G-���a��rٙZ6�e����6��憋�x9��[ț���rn��ø��=�.ĉ��p�����C�ܷ�`�Gl���|J��rŕ���,�y��=o7~�;1�0v��CZﮆ"w&�NT�MG<��{���2�G�,���m����x�9Ҝ�o�#֨��w)ַ��b�K��
��J��F��!��������
�r6���[°�Ra���qn���ӆ�t�_�i.�@^=��?�~2S����W0%��ь�ٙ��]څ�=X-,�V�qu���݆}�ף]�u�XI0�h�4�d�UV����LZ�����I��V��
6�'=}�cy�}|��Q�\�'J���f��X�ܙ� � a�SV�(��|[��iL+���b���k}�ub��`�t�~�U�:U���n��?�뚆*!�z>gu�<�� ��ND�c�}�?qW��8�n�d�p���r88#׵mlY���/�'��-Q����Y��U�8�O�}�1UՁ*	���l��Ţ&��O������xLd�����?�g�<t�狕A�)O����{`{)]��z{Yb�U0�ř�C�p&�e{euL_��4m�z.������=~����������>�~`���֜����z����Wm�;�8�f������u$���k����x�eSc*�+|g��Ay��0�2�������5��rqƍ���5�oRS�vV&��F�^��똾�*_��.=��n����6�T./�%;���3'E1/�1r�ތ�c��87Z�T ץ��:����Kq5(���%��O��k$�ǝ
Ah�#6�}�n�pY\gn7���v�B�T���k��c����hF �9<+(���8����w����o�k��:�e�<)3�P��;x�v�UMZ&��S��y���K[ܕ��S��Z4gAY|��Z�'o�m4�Uo��<�=�Z�Z��94_�8����>���b�P�]���{T���P��W/�櫺�Cj&g�g��o.{��A��r�r���w��y&��<��1n��+�� ����r}�j"
#�;�c�#����;���=�Q��\G����o��9����u/�^��]u�����S�Y9��z�Y3�'���3�)t;�#��\�io�~n�wp��23�:�Ï�;�w���[�4�D��N�w.ǸT�GfD�xÞ�����f{y�&�t\���@��W�KP����<�jD*��G�~�懣dL`���Q7��m��؞��U����MN���wV�2�g������o�O��%X:1�KoS�J�q�*�F�3���Ƨ���2��������(H���9�1kK�3�v�4b���>�B�\�o4��mfL���CB��֪�y|��d��׾���1V2z6�TZ9�j��*.}.�\@x�w``U�<����܌�e���E/oq%�LD��x�[�O&yM��ΠO���7�.9�g����Z��ԫ��{y/UO|dK9<������>?T�ϖ9{v�֙ƞ�z9j�7m:�B�AgVh�Zz���
����$������cZ�gL���F���6j)K�4��^���Xy����ۈ���� T���^��u:�^&=7�v ��wZ���:��9�0�|t�&w���ɫ.���ē{e�e�z6l��o��d*�������uO�8�v:(M5��]�/}M���r�Kw}J�'(uX�)r��SzzBC2w�Ə?<G.��Y�LO����-s3�^�G�q���Sd���n ���3G�lP#��yw}���_n�ɳ7���6���'g�dVܓ,|zߎ�z��^a�[/ꖷ{7O����غS>��M�Z�C��xx�n~�ɵ~���ln�����fg$�=��l�;���Cd�J�nVR�����&L�̨U!8LM?"v�S�n���a��	�">��\��4V�u�rl	��6s��:��l�3ƀ�ǽ�S�
��Sv+��lO���ء<^u�3�� �������}X��;$�v9���D��H�%�Lj+W?2L��|����y���9+��=��1��j�T>��訏+��X��qww������~����PiJ�K�J'�����r受=|��-��
x�َ|ܡ��N���QN)��GW����/�_W����T�Y�?0���-Ǵ�x�_|4/Y^:������b��<���yjţe�$�Xίc��C�A��X�<٩�[kW�y��yJ�����;��]X�|�����6=i��dZƼ�T.��kj���<�h\�!����-=�������Q$�����V����f�����re��[9�A*��ݭ
H�ʽ��Gs�z�]�ڵssC��V��jo$���ޡV1�dP����P�:���I����"��h����j��Ѓ��]����4W�X�wkͿY�f�az�b+&�1i��M���;�߂�����-�'v[cwf�9����E���e��T��o*.�ص;�5�^S�=QU^����y����F����Dj9s:W^\b�o<�C{� g���ytl���>=�{��~cq{sK�3�^W,�,g�R���Զ��N]{{-�f�:߫��3^͚vy�����j�ϵ6�_[Y�ֳ�N��ڏʽ}�-�p��y��s�qT.FRnbAӛ�{τ;�Tو�Ӌݪ|�6o>��7�#�f�C��j�X��L�3{��8����>�ɭ���U ��z#ޮQ}oeW�rx���]��D}�tX+�C�-�{��~����/���|~�yٓ6��	@�ļUX��<��Cu�D}����+���>=�^C�����z�_��ok5�*���V��:p_���,D�=�8̝�Qe3�g��}4����v�^��⯽���;q�@��wG
q��Ѱ1X��]�΂?��P���b��gW�V��-�"]������/�y�=겝���z�ܯu��B ���}`�r_��E������Of}�	�[������M�}�#��~$��ڳ5�@F_�F�%�n�s�L��ŗ�n�Y��������+h��y��QS[�e0��]nv�2�*d����Wت	v�}���(��P��)��`4�-V�u����ƭq�)�%[�m�8o1����Y�O/����7�(���.8���i��Ipȇlz���]�Mg�j'3p�6�:�E��{�]^g"�|V�3�<v��g�G�>c�$|A�pNFАf���3�T;���]X��@ě|'s���&zW>�?U"���M��C��O�T�"�sgە���%c
��/��:�Q�ᷢ�s��Ska9��[�  }�Yv�Q��X��~�W#[�&c'��߸?n�N�ɾ�r..�l.�J2���YOv��u�^	��Ed�6�ڶ½�0�QH����oy9�͊�.���}=���xO��v��R��j��p�z��߻��ҳ� ��}ه��mP
Q���"��gf��+Sɝ�A�˴��~�ٙFG�]����ĩ둛k7:T��u^���=U;��gp}*VD>=5J���+�����v/��^�wU|�N��	�4���Tx�T[ɾÆ��vn;�;�/��WI��rf����|Z����4q��	�[w4�j|�b{�.�fy��/N{ؽ����U��gx'��M+��/�f��0ȅY���7`������ϊ����]&Iy��F����zx-��,ޒ-9��	��~�N���{�n:�����yk_m�a{3�P�A��Ź7}��bp�pN^�(X��u13]���Zd���el>v`u����x+�cT�C���ݏS��F����-�����&̋���̈��p^0�y�T"~��h�)
�N�Q�I��v /t=p�1�R���t��L���&\.ܦ��)֐�8U�H^o>�z�%cqL��5�\̤Z�s���m���i���4��_:JLu��=Q췭�o^)�\s�D*�ї^������<��Z�/�)!�'Ѻ8d9�O[>
��#l'W�w&a	�4[�=.�ϧ�۲��6��{_r�$G���a*���3��o�%2;���1��}�Ѿ���V+�P����F�¤�^2r��`�H��.Կ�����&��;f����L���ͣ�����DH�>�/�/Ka]����k+��kޞ_"�˗ NO��U�]�o}�<6H��~ў���g2��N��k����?k�+EM���yΨ���[>�t�����#��z���{K��$g�J�ϔ�����g�Dt��/_�{ꗤ�x�Ѻ�U����Y.m����k��s���7����J�g��ᗛK��ɓ�l������u ��]��h�coن��|.�T�5���\�"[1β7��؟�f%y�ґ]�$�?zgB�HD�d��4�.���V�k{����7�sBQ��`�^�Fm��=��R������}�U}C��3l�}�j#���p񩀽�be�z��^{FuP�Z�)�#GO>+վ�7��Z�����r*궧Q��4�՝˨(�E�X���é����N1y�zX
Yt>����[@�M�2/�pv�{��N�]<�d`�ե]ŵ�1VӷÓy�%J���#9����ۥ�� ��{�yR/:���
��ˮ�@�=*^Kr��P<Z�²B]��iŝ�gA�t[ZU��
�������[G�ΘJ�-�)^��9y;���:�*wt���Y�n�5���B[Ӯ��foZq��32���YZ=�D1�쏮�5\(��ّX�b�����=C��p>��7׀�Ϙ�^���6-[���B���>��� �����%�@�y�p_߾�Vrg�_k�5���=��ʙ��z�۬q��r�^�٭�����m8��z�ߝϡ�9��b<x�����ݷ6~~�$�^�CN�g�R���O�߼ �k"���յQ!�K����.��VԻeQ͏����p�V�Qٕ�ﵽ�����y��D���&é����������+�.F ���{���/�|��}��ڴOG��*�]�ap��N�K�Wd�U�R�(oY��3�{���m,����OjX<��b��]�_V嬼g*/S���[���ߒ��~X��Kdۮ�?�i�TU��?d�|zW|��w��9榙���
��1<��d��Qp7�=��hGn���>�e�ҽ�k+�s'�瓯�v����o����@���K�'7���q����e]b}$P[X�Cg�n:$����N���O>�uw�]��&߸f��FM4��1+��G��^ԍ���.�M�߃s��ȣ}�=��{����Tt��la����6�<[Rͺ�㓣4��l�aHٌ"������k�ܩyZ�^Va��70!���a�k*D�X����䋗}���Ŷ&�C�j����+��3/E�1f�|n�7,&�Bn������}`��F���.��pҬՅ��tt8r�T��.tckX���r�;\6�xz4QoV��^��cxx`���Rߍ�'� �&�;E+���n���-a�_��7�����}kXw�ǃߵN��3W�*��bs91�tT�O+Xź���>.����1�$�k#�.���di�q��]_����)�\-��=/k>9�o���t��o�{�ܒ9O�O=7O�<�ʽ���J�N� & ��w�Z�zogxǄ:����������N��[���9����l$kr�-m\t'�摌���*43��b!�Rx��`���5�uQ9l�z&�V)�5�M��/�w����oyR�����mzU��T���p��>�G<��ܓ�;熲�Gb��U��̑=�}e�]�򅤻�D�W>��M��?;��bA��v��[^ʯ{��_��s(��u�ƭ=A�5B��+;=�߮T�9_kƮ�����Xt����߭��|�W.S���k�~��A��Y����Ͽ����{�d�ӿ̈��{E8��ӽ�1�2wMF:��ԧ���L�]�������g'�%Ղ�o������]Zm���N:�����}{{+sQ��/�0'��_��������Ϥi�ݑ���˼����1�c�7�䍃n�����d�~��n�� Hs��!����5�lŴ�nԟ09��7�)e�D��kf��Հ��e|E��^Z��)��;�4!uՋE�26���$�:.�LmV�=�v+םO���m����]�������"���]�7��O5+gksBq��֏�i�w� nV���� NXy�s�y:�G��}u%2��2�,Ygu�(t��d�W%^�����ׄ%�@�t�]/r�h|j�C���\{44_����^c�KH�Iw�Ӫ�8�c���q2���i̹��>х�M	8��L�ۃ.��J鐫L����9z�B�c����1����b������X�sҮ7o{�p���r�/�ې�� #�@�t��ê�W��i~Z���#}0��--c�'ʧޯ� dGL�K�����;_}�Dug7^^��Ǥ��R�u��ف�zj}�s'o�z�m�o?XB���I��W�c���j��r�'����]�O
��n��N)���:^`z�&��HF�}L�ẓ����eP^��8�d�{��"Htkߎ^�w����3��}ױ�;�9pAmn��#x.��*Ԯ"�/M�����)bϭb{y��ULߏ���}��kG�>��3��_�n�}�9��S���Ϸ����ːr��O����@�I/�zn!�:L�`>8�D�])�Vf`{�)S0ƀ0���jI�����^)�p��S�6k�ܢYٮ�·<x��Ӳ_�4׾�0��@��h��le_�}◪� /���t�9��ف�ާqe���߁�Os�W_��r�(���f�_EY��DG�Ѥ�;�Sگ;���M��#dI�=t`���ⷓEל�
��N=,{�e�o�f��PVt��U�k�h��(s�g]oiн�b⼕�Y�)cȖ ��e��H�����E7�-󓲺��k{��Û��]�	V �	;u"�kd��Rg�b�J��^��-W/a�쫵���Ci$Kh�V=��.�f�3��V���1�y�ss��:�ԋy{e�i�VUn�"���!���H�b�]{�>��:����Z����Ы+��ιc*0D�p�1�T��M'22�D�U]f)e�����_ɂszܚ���Qן��c��0<��<�>�|������v�>�V�bnrڕ�(7�o��Y.��g��|"0�z��\�-��>pAM���栤�7�����3����"�/�]�1�	H?t��u<im���^�ځy��)Ŷ�eэ~s�v������䥔'�zvg����T�L:�䯭)1�;G5;���FN�U�x���d5�'N���ue岸��1��/l�2�o�� ���%K�5��r���Y����J[6C�ꫀlv�>�����e�{w&�:��нF�ju�ס���P��
�����gG.�R?$��?�.a}���1������CĹW�qU8��3;���dH��91�C��y���3��Q�k�u;������k��{d�nL�#y�b�e�Dj��Ya� E����3;}�yn߷>��[�[�3���w�����|���gm{�X�>F�t�*O L��T���^{�h5��""���N�Q �WS��X���(oz�}[A1Gβ��W��4��zs1��p��z����H�7������5����M���M��V�;��J�w87�m�A4	gi�F�6y"���5R������x�����\je�y;xY7@�m�H>���]�7�K6�%vY{e�$+��P;�%Et�宵u%�.,���[�;�w�����g9κ�7֞l�ڳ/�F����o��`Z�՘Q �ɇ�0�WƮV+��h`�R����ޱh:n˴�	�l,�����hXY�p��\Ò�҇N!:��"�]w���v�N�7̹�'�C�5+-����^�a釺����0v8�w^>X(˫��,����L]vh:�"��S9�t��gLgU��op9R�A�j	v�!jVy>�t9͠sn㫐�-���&.�3���D�m���ǈ�]����+-Ŕ�#����1+�̥�����Z�kI�u��uL���;E�n���Y1�c(ݾ��K[j�rs�M��w�np-���7]�l"�iS�ݴ�Ӻ�r��t���b�֯.�����ĸu���]FL�F:�e/;yo9wڲ�7Al9�_vo4L�ܴ�t��cB�N;z)ξn��R=��[n��1��-����+4�M�J�;�+��k�ޱ��Ŷ�~�gM�_RIwKE�|e
T�=%�]�����۾:�_N���n�R�A��R
��v����G��N�V�,�t:�<���W���f�>�kv�*�i���i��T��V�k�������ڻ2�	�J�i<˩����"�]�y��z\��v<rͩ�%�ۑ�=wG���J�%Ws$��ooN��Ĝ��N������z��,�C�1<��CVl��]6㤝�Z6"�4�n�u97u+{�	��R�����憭�J&m�1㐶��]��\�-AIcu����:.8;�At�P3Wd���l�ŘwB���M���4T �m��o3N��> GN�u�C$��K]yz)	\@�)s8TN�|�R�o�9V��mm^a�;ΐ��V&%�)钌���JS���u�Q[e��^���M�OǽK��Տp$�
��6z��P����r%S9Q'�,��q�W;�8fC�+�'J&�땟
X�t�70�
U��ا-�2�Ӎ)R%���rme&*W�3U[�\M��ħ*v���k7èE{�U�DΡ��l��%qC����]1���S����Rr�<���0��fY�͵���G�K��'�2��ػe��3/��ht�oz��A�;��7vT�|���ȷg�8�/j�#H��p���t�Ĝ��Woi���لK����5ܬ�cM"���8��q��]�H��t�z�f8s�#�ʭ1���e]�*om�$����z����w~+z�4R�����!f��.`k��3x��mQ�W۟
�aƸ�l��,;8�'G\UÅ=�g��{%�;I;3:TOE��2f2zT�.�����R����̴�l�f�݁�-ʥ��@c.����,DK�-�T#Nݧԏ45����9-TC:"���v�Wn������|��:��ɮ��Cy���V�:sjn�:9���eB�������mt����۝�7~��\΀g��ح wϧ���Md��3X0����IO,mlh�-ъ���G}��3�~���s��>�N���r1�ξE��:_]��}�Bc�]�
P��o��yl㈇���y��f85��wW;qXʫe�g��f�H��/aL��u��I8E:�c���V��JM��z��͉w��s7�w+�=V�a캨�y���B����p_M~����1¹��d�M�`gѲ�����v&ש�Ơ�J�~ߖ�W�ǳ�U��N�!`L=�����_v�h�~o��g��@y���ɠ%��M�#�~'�Gw�침�jE��q��`�'妪��!b�����Wp�ӭS��/_����e�<����.E91�W���	N��G�l�U1n�h�\=\m\�:k��N@^ ���ܱw���(g�\����R�G��w�?E�M�C��`7=Uko�����=�c�����+`⊠�%wH�rvj�LM|�wz�����I�e`qP�Q}�J�u���q��>mx�]���(l�~c�]3ן��V���<%6�j\�1�R��&ɬ��pJ��%_���_Z��#�c�ѭR��)*�m�oc��WD4�p���$x����;��6�N� �tIo�/�DjыFaF�/�Sd
ѿ���9N����ٲ�po��ō�7��^�@Km�}K2�7��٫C�n���Id���:^�ԩ[ۑ4vp��֥��kG�e:f���/��w�3c8&^]�+�-c{��S��N�.8 ��7-�r�Ku�M�hJFK��g;��h�~$�o����蹜�⯗V��͗�G	��v���Mb�RP�wF"e9�9M�al���f���e��}뉯�'��R��l���%M���R��Y���.�N�{\��>f9KgL�Ỿ��Wٓ�B��ks8���t�Dw�T�c"��m �{����2�fVӏ�ޙ�.e���`��6��;A?g�#��(6^���6�1*|�擥d7�]���]J����#���_7�"���d�v#�=Fk���eb=Fv��c���ә�smᩡ�>)RI�/�ҍ��姈���y�T��^~S����S��~~�5\4�q�7^t�����p��J�j�����Ǧ;�jg�W�٬�������6|*zg����������lS;�s��[��#��s�7nߴ>̫az�^�🆸�^�V^ȱC�"�-�jMx�b�9B?��
{̢c��ϭr�:�R1)���[�Y1�t������*@��}��������Փw*����*��u1�[��7����%T,��� �J�)FT�w����Uvg��N�جK��a��"�K�s����A��Uo�*�E}�:|���)��6}<���]�neP����7�5]W�Y����Y�^�U+V}&F�-Ds�o{Խ�z�`EP��N=�]o�*{6�	��u�j���~B[��`�P\`�|;�i�yZ���!$Uޘ]��dft�T��� �Y�����8+c3rj��#q��l72�u�St�U������	�'M����qP׼�^���9ox�2���a�/h���;����%�#Hr�ޥ5wi�q�,�t�z�/��잏y���q�\���^�c��b��^e+���Jy^��G��2�߅�[��^0#�=!��noa(��f/�,BQ�Ҟ�>KО�ю�ɿ9�~���k+@/��� �﫯G'���nA�ϭ� �:,y	��z��mt���O�+	��������O�b�I��1�S�+�l�Ӿ���ƨǷS�T�z;�m{�6(�3"|������Ds�.�v��$6>�6m�;��Q�ʇ�e��!�^Uh���(ʲ!{�8�ꛠ6�Fp?^Z����S���7M�&r��^+r2�׳�m^A�c��̯���EGp�{����`�$S���[�b��+'A���z���y.�%����z\���^ci'B�T�L	_j^P㈻��]uK�Ƥ���^�,��,]W��`D�8����{f��^zv�%�DoO]Uk���Ժ�?;��[�G�e&}춃&V��`'�r0��5>����*�8Qr�wb��*�������goz��}WxoZ3��;�p�A����iq��x��+�����Z��>����c��z=��{��3"�,v����3�u6��O1E�O�:�@�����x�`���W=����e�����X��g��@͹"A�z{�������w�H�=�/�{��r�~�S�;���t����g0�^+~^�6�p�z�P���:��o�+�_[D�����D(5ͼ�=�vmtL�l}Ke�s���u��&@�}���K�v��%v-{��e(u9��%T5�o.5�T6)B)n�ys�{ik�_]v�{��z�Bu�`��q�BS깻k����k_'���N�ַ���3�V�M�\xeb�}��5�;���E^cUE�dA�����I����f���yWE\c~�b�p'g��C��񖙯y�=0��.���{�"�Nu[�˛~̋R���i��H��';]4�~����,o������	}[�d^�7�����	rME�˯rp��]��:=�:&\B�@Rs2�XA+c0Z���3��zb>�}^=^���Ȯ�e��
�hb"d��_���߽Og��WFd�!A1�]��a�{W�R�d���AHΫ����^�~���v!�"~m��
�X�݈�!3����E9aǧ/��v��5�|#���k�>8r��n�z�߯=�g4�ά���{�L=Yf�pz�!�{yܚ�X/��q���wxg��\�ߴ�ڵ5��uT�.�9��P-��`�2L������ǖҡ_�Oa�ijr�<|(����	�B�:��ah��^`ev�#��˞~̟9����+T1���uW�'����Q�������L>����	_��q�������o�O�!��tvo�7N;�K���SՐ��=k[��=�� �������'2��E�Y9��ЊDuN�̣��v4�-7�l�qֻ=��du=v���'���_���"7�=��Q��$f��ËG^?[�S��)�Q������d���wed;���} 9��ȅ:�ɖG�4߽�T���P��%g�[ض���ŧr�G&��hJ���E�Gfiƈ�Y0
�h��:��ĝm>�+M���|$��&cYrQPU�����f�T�Q���u*'�	o�$��a+֩P��r��\ڎ�kܹ��ۖݿ��;b<�̑Y�&
�l�C��k�����ދٕd�n��q#>����\4;!_ -��ʶ�x���U�p�W4�NVW�V�Vv�Đ���e��{�f�~���tE�?��_Ն�~t���͑���5J��$z���|�y��G��%5�ᨪg
3�쑒	**�����=zK���U� W�}�jҠA��R�}�WP�\?[��'�W��]eO��#�O��i3���F�����*��Ϟ��Fr�";��#tM?\��M��U�Gaw��Q왛�="��}a�_v;��'ǚS����nMG�5�)f���!�}����WZ0�>��q��x��}��$�~rNƄ�����|��:+���F5_6UGʳ����E��NY�� ���k-G�cV`��n��v�yCF�)�*9ȓpS�/]��\���P|����DZ۵�ZǼ��]6�hł�\�
���ů����4�#�����U��,}PYy��d���T��L�л#�\�^�Μ��E��ؠ�����v'��TԿ)IC�b�u$|�+�4�W@�ǫ�q�T��.�J��_y<����xw%�^�v���>�=Q��#edq�33��I��[%f��/�߿>�n횅�?��`ȑ�ۚU*��)z��C����UI�{���U)lI�cI�3H(ԏX��O��*_C���]�(��ѵ���^/�:����}jڌ�>��M{�m����'�s�ہ�ٗ��� �ay��Tx�v�b�qb��(?�j���Q'������>��^�t��Nġ��Nth��^{8��uv�.Bf��/����/l��#��ʬ0�\7e�����#�����gpV�ca�$^u��;G��9�;q��^�7U�k�[Ą��\�u<�n��n�zN�]�����z��G�䘌Vn�Rȱ����wz�0����}�e���^�|:�����YB��>�f'�M�����3��fnfK���>�wJ�'C�l�����T=�ʨ�]:�:�åE��i+�;<���y_���C�V+�9��f�p��hhfb��gN^�y���y��@(��LǶ��i���fd�3Lέ�S�h�u<�B�c]~��uh� �1$��:��Г3�a��k�r�cﾒ9���$:�E��(Ww}��L���I��<�����G���}Zɏ_��D�^Csp�_{�M������?GL�����@%���Y�o��_�~�>�z�<��S�.(�o%A��g�:M*���tRrP�R�u�3�֭wx٥?d�}����5�����kb�+m!���9>ߢ�ܶ������#�#Ϊ�^('s�_#�X	��HLΪ� ��2"�{��64���a7y�V����EҶ�t���s#r���c��R��T�hd��Z�:%91w���Q��8�:�jw�IxG�5�į}�>�g��f�
�����>���گs9O����f�A+�ɿ
����Sz��A��ʜ!"�#�#���E�U���T�1�_����y�6΋��ٶ���?d��3�&�E���~hx,��P5Z���j���^���c�$���碣��nS��e�y���#����w)�Ǻ�V"��!��dz81~B��[47sWo�Y�t�p�j@��O����� �P1�βs ~Ǌ-�z���j�K��	eBR�GH��`P��W(�%��g�)��Z�H�0��p�/\��+Tqi�ϒ��[[�[�q`�4,��=ݔlZȓU�vw:���3UF�ݜ���A[W�a��:r��2���8��"�īS����`��p�6����Wr��W�.*3�������M��jaOza���߾��R�uQU��B�dӞh{n$���#�ְSC�P��֠�}~���'�n!�lc��lkr��0��/���Y�]������i1���o�"�o�Ҹ��!%�z�3��7e/�x��n"b�1���@R��/��s��8���-]�Ӵ7j����mEʥ�ܲ&��G*�G��G?��#u�Ǽ�G�a�U�ڱ%j�����ƌ��z��f��>��Vd�e��":F@Q�=A�\����ty�����zG�{uvhʂ���Y��	�&�G����΃\�cԀ��0�I�9Ż��t�C�i߮��N��0{�}r~�7~�Kr��In"=S�{�W����͒���dC�$#�Q�S����L���$�&
]�1:)i��`��Ԅ��5v_�M|q�DWGET�y���7\����k�}�9?kv�����Տ�zD��?xңH��5!}�	�:�5Lw�QG�V	Q=�+��P+j�dgΝ�U%��Lѽ, �\��ٓ���m�W��;��ՔF��g��Ő�.�뻜�\|�I����wp	f�*Gc�5��U��b�а���Q�=��'�&��Ɲ}Q�vs0�9� H�NL��'�ܭ9��I ��)���p3�h"��|.�)�k��~CXG��7 �����t�]��A����
�����{s7��e��U��w�<w�8�w\�Ck�O��2LI��0��2���>YL���H
�L\_�Y�Rɱ�b��>[��J�t�":������yF��πX� l�|��T�e/�����9{j��b|���k�*T�L��B>E�y1S�IH��U|�m�Ӄ��k�7V����ݦA��L����u#��t�7]���v�A$��X�z�&�a��Ec�@���]5j��*8Y����0չR�(�K�D����=�r�j��.x2�*�=�k�n��onR`QX_����'o4�g* .�+Z�� /��:�i��Ek�,�v�n��|=����� e|>� T�<z3 99kJ�1����=b��	1�Q��ٍ?"����Z�>e�}uvc.]�yg����z¡���������=�+�:���"�F������nr�?H?.#� 	F��,�#�0B�U�����C!�����Ta���eM�������
rݿ���|��RbJx��R}9R>�,�ܡF�� ZC��`t�ܣ��*(��] *�ŵ\[�S�F��<)�/�����8�P�%}��뷖M@�׾5!H���A��8���`�[�+"��Y1�	��{}t8�^��W�PM|c�2�|��`(��WϽs "(���B:|1f~����Z��D}H"&��~_S0�M���{�N�5������E&y��${�����{����˅}G׶b=.�a������zu��ޛ����c\+�7�8��{�U���59�F檒aT[��7E%��
�T
"vꬲ��Q<�j$��x����B"��� �y�h�EkpR"�'(ԣ���{�eO|,k����Ő�A�|ި�ɉ3C=�ϷC&d��<�0�km%�-LQtd���P'k�E�$k:�<i��n�#?,�a�J�l�MgW�Җ^}���1���ȮH�0/��"�<��Pt��K�"��/����08���@$�u�$m&qӳ%��p6�>�ꏋHMl��f���ϫ�"�F�J���0�j��f����W��?:�z��Wf��>x���2��m@;�0��D�M��
��_�Q��l��B�߳�FH��?)�f��>�:�^�^P��>���
>�� {$W�݄bv� x�F&�`���}����>_+�d
R���`E��z�EG��ܶ�����e�>L������U�T��k_~&x�
�Ԫ��i˄|�::]�.��F�RYN]K2�!�4+��f�95�Ѩ�b%���oo%��@e�$l�>Wd�qtu��SN6�+��EW_�i޼<�c��;(�uC����M�c3���o�}-j��dQ)�,A5�1F>*�D3��Z�؉��Ob��1Q�����4�����>�w��B(��]a�߾�t��(�us'�gR�q��/o����@��j�2A-���J$�l���136�>m�.�f�Q�"��\�~K�!�2`L�ƙ�?~Y������v|����T���rHu��]�U��*�"}��Ei�+P��9R0�#���=�kH��T$����G��G�ś���[�1s��԰f>2����G.�4Wn�3�XK�eex|�pkoʆJ�D�T������5��^@n`�%�/��fH� ��3�Y��懵�k鿩|@5b�#��`e�Uf!&�>��k�?�R5�eo����;��cH��gXÄ"41�
��@��=�dx�|E�~���0M�dW�*�䆑��O��68��<��6>��~~��1�D<bn0Q���
]vW�˂�Y���`��\�6Ta:ņ/����
�@'@V/V(��\G�Z���$ $#�ް�bi�@�͌��S��]�����}���Xa}u���+������i8D+p'�2��ه>�	�J�
�8�=�AU`}s�t:�<�=�r�|`���������Չ��I"	�}G�8A+"NV�q�G�r5�9}�]�2���鏨��D�3�1^"�,"(�Ѓ��!�S�&l�$� �=�#�m �)$��#�G�WPab`���&U<��T�4칟�W���ܿs����g{�P5��Ē�L��c�&�� ���g�#�zd}��I �ㄐFK1��#�آHDKI����19,C�n>X�.	�M��:׺t�	����Zk�r=�tD6t1ǱlUP��� (��$a�O�q^����y���?UC"�3'�LI�	�=1����0�a�!��ˈ�d
 ����%��&���{C���v���ߊ�}��,w�hH�@[�[f%{�yJQɹ'�Ӱ��������n��)�6:��A��ٽ���whP
���挾��C!��Ar仙.-i̖�ɛۍm��T9��2볖�]���7M�w��t���mm=�Π�;�������n��Q�ݽ��^��x��1?{���P�1��)4�sB�Z55 iF:�p�Edy������~�`|� �#� @�=�$Qt�l��G���H�%<�=#��'�NK�����|`{�z��I�4���=(Po���.>�Md"#=�ҭ��iT���=�7�6��bH ���L(�ٓcH�@e^2Q��U1U�����d1�FZ���Z�~�:�����T3'qL�� V�����R(�Fʁb}z��ȍ!$	�����2tz��|�� �Ϝ��	�C�P>�$B"�<�p$�1�Q� ��f�1��1�P�i����̩��\����c��J,�$;���4� {�$n!� "��b�t�+�B"�R@I��@*���g���Y����`=DJd�*�|�Q��@~P/���j�_���u�ß^_F����DG(����+b"�#7i��Z���0�RUޑ�a�`A�D|G5rHLH*\C iZ�B1PI�L����L� p�f9 A��!�$��F�J��x�X�W�����Zf�{��N�����D|@�@iR�@���1ﲦ ����P.��:B [B�<�.�G�DQ�QX��"}L�A ��S ���;�d� q�9���b=j3HG֠d� $�r5ʘ��ga��/>4+ݼ| a��C_1�` :��;�� �"�U�(�<��C1���>��i����@�$3@ӆ�F4�`2"1 <@`@�h��Q����C��J�D`Y��������,鞛���=u���& ��H�q�*>1���!D&���b5�f"�f ���<b!�F(J�b�F �!�D2"8�Fa��(�dGb���0���	!�b$�@C1�څГ������.���}ߊ�����`D�� A |@�1��}�@�D 9���:`4bj�D3��~"!���őf! ��=��Dx�@@�b ��p#��"�F��Dڀ�j x��D`@�����^�C#����ٺ������� �0	�* ���1$@�DDn( a��0�P��(�"P'rf�x��,��g�7�H���ܭ��s�� D���@����@�����"DB�� DDQ D���"��� D���"��� D���@�����"DG�@���D"!D@�"",D@�""?��"DG�@���" @��D"#��� DD~� @� � @�� ��b��L����:eO� � ���@  nO���F�u+�T   7�n[b� ��U H  �(R�(J�� �    u�     �]��:T�����6ҁTQl�
6�RkU lȩ�m���QESA�*�KUL�TP6� ���@�m�J[�ӢBA� ��kZ�'���ʼ��������S�x�]�6�.]r�AW=�J��Xq�Oyym���nP���˻e ��Ҕ天O3s͌U�Ѳ��˺��O{{�m� PP Z=����tv�

hy�򪪃��P����4+����4)���!�tP����У��{Gw\:�(zn��4(8�
8��ݬ1�ۺΊ<   ׁ�P�JW��i�����tQE�^&�)����Eb����&�'�q�錵7�T������m�{���kJ����V2Q�\�ck�{��M�a�Ԉ�w��ڦ�=�z��6ԮvWZ�  �m���@�ږ���(�K�UJ�q^��(�b��`wgzǧ�b�l����h�F��Ǣ��s��ż	(�x�(��`z.�[f�1�yeu�h�    ��HT*�*�l��	"-�AE�+֎'H���w@"�Z.{�E=1�������JQ��h �n��lVٷ.QN��[��K�68�)]ʞzT�{�ٶҚoz�׉��K�a  4 �G6�B�M�{���m��k�P��*s��3J(�^�=� �7Ez!ޱ҂�=犩U�k5��;�jm������4^gv(�5�GN�mh �^�GX�P��K`����6�j��bpɶI绢��:���{��M������z�b��Å�۽��h1l�ܻ�V���x=/X�=䊉���*��c�z��m�` �  �O{��S-m˗`ҵ7����)Ow��#ٶ۽�K���=���6���h�E�=%
w����o;���糽-�@�����דGJЀ   ok���%(�j�!P*�F�^:��ӝ��m��m���z�8��M1�[���V�Fnz4կ�����p������a��r�M��;�P��IR�������kmw;;+�    $�,N�cmy��m�ب�ҤN�c!/y���{������:{ea��5Ť�<�(��^R���w��������ڶ�n�(5�ܥWm� �� �TѠ  ?$��    U&�Sh��OB�'�T��%*� d  ��UH&�Jz@т=4�&�*�@ �ÿ'�-�������g�Mm�W�+"���W	�{fmv���YP�z�_�P��RP]��ʄ1_����P�8�vĨ�{�������]c������a�Ϯ��>������Q�w�<4�����3:�^�7���D�)���N�.-��<P�iYNk;]o-)���J�	��BmC�:9l�3���TJ��q�C�h��4�Z�vE�]����|0%���ēk���UWJ.�W\����F6��=�'�0�E���M.�r'-�B���5���|D�R�V=T�T}���7giTy��_�wX��Eh�?ա�a��	�[�j!�����%�'!�a�p�Ĵ�?	�U�N��@P����e�aWN���
�ʁ	��)	��w���r����[�3P��l��Cf�ݾ�ֳO
W�*k��}r[��
�R<+T����0k�����R��D\���Χٝ(ҘT�w�3��sѯp6�r�	�5��J��ѽ��b���-*u6�j�u����0����T��F���!�Ow���TÚ���l���=}wz�v�Ġ�J�01^�}�#�R7R��9\c�wJz����4�0+��λSW5��Y)���ufG�e����nWn@�W�Y�Ї0_^G��7��f�Eڻ4�һVJb=�ˆ��p]�"Hu2��7�N��zB�9�Z��K������'��Z/���y.�+ΧE�Ճ�[W�5��gur�L\���+�v�8��W���ـ�I�Y�ٱ�ݵ���.p�}W��Y�3�=9��	A�;U],�N)��w[�u�7wySVO\�)�.����ˋ	޷˝��l]|�����\7o���d�]�)H�	vQ�;�Mk���c6��9��z[T\Vn��V�G�CSP�YHQu�w�W�8%K��mq1��ҹu�m�r���Nņ�h�ܶ���ov��ch�Ë�ؿ`T��]��9T]'\�=l��شp%�-8�:&�ʸ�nRNS�T\4�qn���ܘ{%�rƅӬ��RAA��WWeW�3�������m%Ƒ��-�Ac[��Y/.&n�Q��f�Q&�7{KEf�I�!~9�Z�F�kFՇ�ֶ��]e$]�^���Yɷk&�D��'e㙲J8��Y�h��0rϘA}�=��>�y'��	��rD���I�pOӿ	㾝�I���I��'��rJw������'}"w�N�N>^��I�w�N�w�$�w�}'���;�%;��>N� pOӃ��>��x�O$Q\�>��"O��}ȉ"�)ݲ��#[\<9؆�fұ��i�#�6!���T|�Z��u���ik�7��h�T�N�����*�+Ž����Z���@ܻ�7(�T���J[ή�uu���[$XFa�}�1�昱�P�ދM�*�w�F�kK;�^ڑp�bx�p��)k&�ٮ�r3��6n\'�,�)�����R3B�飫C�S�:�Vܵ]}!�ͦ��9u(�D�ڴJ��ޱǭLο�lD�+���8�/�I͖���*s���y��9-kx�"�*u�����i)�!]l�5z�����	��f� ;5���a\�i$h�7�B&1����{8�;n��]hu�q)��[�[)w:<�''!+�����=�w�����]�f-��s��Rh4]��r-��5[�[�%�>/v��n��Et��ٺ�+z�R�"�D�6�e�̤��U�L���uz�5-��9���Vʚ4�%��
���Že��]���of���L�(X�;�8�{iP)I]��*�Ҁ�6��VL��
�y���k�b��;,���W5���+�kjm�Cg`ذq��pBgf^����&�S�Usnm�y�[b�t ,)F��墎��U�=;�E�OUe��
�T�vԩշ�h�m����T�]���5�:�ˋ4�E��b�h�6��c��Û��x>鯭֫꘡�'tQB�`7E0����Y��C�lљ�����5���U�A���P���r�@��b� ���0��1��u��N�7m�M�8:����k��D:ˊn=����A��3q���9���fI�GÒoOo����s
����R��̔�sF���15V^B�Z	�6�]E�Ք�7CX*��7y(�.~1(�x�D�euBB��3D(���3�@Cd���!R�P��so(T�ָ$Tu.�P��ՓMr�!J�Cr��ͻw�sẽ?I�Z5�ځe]�@ˍ�@FK���o9˩��f^�͹@[u�DP!�'s��2n�*{���;���pF���O2���:W�w� �f�M�`�q��٧h�T�^���Q�Sk�ך��Ñ��7?5b≯�F��Be�N�ᨬ�y�q��aG/f�v��n�˃D�7�kxaܼ��"���ցf�I6�f���ԩZV���ۥ�/It�V扸Ujz��Rۃm�����;�aķ+�}3k�����rpҷi�PxiI��Y�wߤ�QQo����y�M�\�!6��Ҏɔ�	kp���cv9z���[�֜�[t�Q��)o%u�Ѽ&�r;r�-�/U��fvi��DR���]yل�[h�,���.�ُܱ�D��wc:V�p�.���nfk�`��Q����t��"�~m^s&Me̎W9O�ӈky���v�-�T�6�8�R�Z9r�]���wF�-�w1�n�Y�ͼ�793�ޕ�n+u�S��a509��Z��q��G�9��#�5���̍Ĭi{�]�e���̽xN0�^�W��ñ���3o1<��+m�*ީto�B�f,�Om^�J,��rƫ�H�r�²e4Xt��X��X�w��1�n�
+bh��f�S^Z�A���[#2Ԭ�M���:��WmUn���0��4[4?��c��\k+%м�b��)�ٸ'�u���7dh���Ȟ��&JSlQ���3I{�os����^�����kv�V��j��E��m��ܙN�,�5B]�H���겙al�r�q��=����/H��׍�[�����`ܺIۃ5��4F���"e���,7oa�)`,*;�0�YH���Y	ۣ��!�t�����zA�u�a�R]����K�;h^l�q2Ma�~��_�Y�n��LЫ72��$X
�l��1tN�N\�/�;Æn�TL�WYÍ����
�fƦ�
���fc4�Ck+FT�o3Q5�U�̇6�R��������=A^�E��i�&��K�Řf��K�딚ޖ�n��x(�mAtS��tD�m���w��ݺ�q���+1�֊c6tf:�k-�nMѢ;-�7.Gk"��yr;SX�y{��5([{���k3�0������9Z��y&�o���k[����Ӎ�Z�4��Q5%����7�['ZU˻	4ee���-u% �^�]]J˥�{��s{�98�]�p�q`罂s&���}۷`��wZ�z�G�ԫ�41�2VD��p���iFY7h�]�R��|�BH��e8���[NEg!�C�Z�-���Y�l*Ӻ�otVm0�z�Db$�j�*Ɯ$�	�C-+�dGH�ՋYk2;� O������Qk��2�t?;�j���-zk<4��f�U
͛yg8���ɋ�Q�MRd��j�ci�X���!�[)���B�o4Y�[5��Z0$�Â�sVmZ۽r
�B�W��Y�Z��ͼ�h�J-��w%�̺kk ���WXTɘ�Z�u�L0���,�L&�kq^��Cj���v"�n<E�Sb��N�\Ӻtٌ�r�=�wn�t������6��=�H�8��T���)t�]�f�m~ܕ�b\�'t�d�<�U�BC!U˨�
'��@z/lg�O�Z����F�ɛv�T
�6�o�Y�o�c=�g!��+]�>��A�1�����O�D�DAu��#(��u��jΕX��z��.�n�+*�gH�I˱[M�+n^ܺ�R�ܹ5iy�keͼ�V�8��ɑ#Y�j�H5��75(lR2�����N*<�k��cq��a�z�K77HO0�K���,�y�Ӯ�r��]�d�3���n���d{��-;���Ж+7�-�ލ���0d�Q�P�9�7E��)e���4V����!�Z
�〬�"��c�n������)�z�.G13�qCn!2r�u���+*��.a6J�%�E-C�7����eOX֗&q_�6jǫAKX��{YsTi��72]�iizt����jf���ǵ.�	ikx<"��f�Z�{�r�7&f��Z�r�n����k�)�lݖk(�ɷ@������o��
�Am���x��nn����l���;a3�+��*TZi`��c��]���K��K�7�(f.�l9v^+���f�m�Ta�#�)C��&��\��(�G��y�����#cX��.���J���Y�v7s�rƊ���7�1���9NU�-�ۼڜ���8$�P����ޕ�u�4��Tͬ�r�b弸,^m��+hq���R�Nf���&�%nS-f8w-�Ũ�,ܫ��J݂�-R�r�r�v��	�$(\6jjxTT&l6+��������gh�'�i�s0T/I�ld�4[���&�rL?M�#cͷk��u=�k�sx�P���R,4yѻ:!˼��췗��(V����x���,�朠�Xp�qn�Cn�b��*��*��?av�+("rҨ� �W�l���Q�׼;��?@0�Xw7[�\,�]��ev꼻;3��23XBц
���*ˋ��#aei��G!,ke-禲�u@�)mc��ևY�X󷭐)rL�Fo��YV�:������<��ugQG��UH�B��+��\&��D��C6V��{���;�\iS�7���'P6-�����29{�f�qD3�(\��@�n]���ˈ.��ogiـ�ٺӭ��h����,���	Cm�Eh�7R`n���\T��qs�,���dV/lne���(�w �K6�C��d��?t("�}�W2�	Y���+�1�W*��Wc��g�B*^�ث;�[Kr�;/���Esk���� �w^��:X uea�wB�;I�v�J41�f3���԰�euȜ����¦�ܮ�d���X��W���<��$��`;�N٤9bܮ�ۂ��ƨvi��V���˷���u7ҭs˺޺ژ�u%�:�{X��=�1�vc��0���j�=�P7?.�(�����"yLĭ��:�WX�QPt3o6��89l�r��8JJ��$p��oI��;�ǘ�"z%�u~�.���̭!���ԫ�'��m�	'k����6�zf
�zPJ���Y1�߆�YQt�^YXۚ�`��(���F���㰭j�5������\:T�|5ޫ�-���W{�jb�
����հ�-Hsۣ���{��]��c(��l��A����0%wuu?F�K��6� [�7VT�u�ǣ{;]l�K:ed��l�Ǖ�N�	=��e������n#�(�hI�bO�;�q%�ؖ7Hv�$�7���W�:�0��A�V�U�}\j�)Qk��%�0Y'HB�sŴ�T��j<s��Ն"���v1��퉬���A�,����4^Ł��E�"��q��'s5;׶ꚿ(Wm<��:�<)����ǯ����V���(������;U��3)'��+�IX��٥i��C4��؉z�vWY�+�����l3��k��5M�t�Gr��ZC�4�%�ml������kb��ڙ����c�ߡ�9HEv[ѱFw���/��9U�m���eCCE;xd4T;���4X��B@to~����7���w���~{�'�� z���k� N^/S��!��mM���b��I��/�_fU)��j�z�����l�g,���r뮐gxo=�n��<?�
2cn�Q������Z"ҫr\eJtf����{��Z�+��+k^V6���k��i�Y�\h8�V��z�C�3:'F��ʠ��k:S�L�����o� EJ�Zp�ޞ�6u
�iq=�a���d}�3����*۶�qq�]]�%�]˞C��!g����\��Ն@�ra���^aY3ܲ6#C,pZ�`�J3�uM�9V��i�(!�S��1�����v�i=Uཧ.�S�Y���fVfؒ�]Y{�zvV܂�B;ۆV��ٸ�4@K����u���v��"�\�Q��ߓ����R�F�t��4F ��H[�%����I���&8�,�+yo~��"*�e���6�*�k,�1˒]e@��L32�K,(l�p�ҺX1d;RL��"j9'�3 �n�DB`ue=dն���#׈���!����v匵�7E���ub��c�[��v�**J�0V�X�l����1�i����_;fVvr5�8ˤ�$-��{y�kM��%<r���j��E��y+p�tP0�rۂ�����!ֻD�I]bB~ބb�2�n�os�]�P��ؖ�!���-!�0a�/S׵�H�9��o��̻�� /s�nx�R�Y�$�+v�3t�e�8�j��m'߶��Q�"�lle��.�=�X�4ج��YlK+fǬ���0r3���J�^�j���S��ڧZ���y0)�2��NV�c4\;��;�:n�m��럛k3��k"��Ef��m��D���=g��c��1S땽��{/�|����+!�=ɋ]hp�tqz%Ƈ~6Xݔ��+�m��۝.co^�z=;w��֤)f豈fޜo*�0��V^�N&����J٤d�0ۺӬ���r�c:cܜq�ul1���U�3%m�U�J����3'��Vmb�d^vyV�,i�����a��v��ږ��gh�Q;۩��!!ʘ�ł�Uu�Ъ���ވX��	U�8)��יq��C�	f3��<}8�vM����Yy�:cZ�"��ej9�B Vmf�W�2�ǥ�Db��>�[�������S����hCx�vF[R�v�<B�sƪ	ؘM�jL��oj_�,��q��Q���w��R��ͫJ�i��ע�Z�+,HY*�zն���Q�Y��ޑ�K�S�'3H�?h\&=�.����ͪ ��j�~�u�S��^;�)5]z���9��9S�n<ќ,k&Bj,�ZT!ժ���'�MU�P�S-N���]�X�ZT�Ƴ7&M��s��Z��6pj�u6cњEV�<��.�WZ0e�Q�`��%,�b�6�)��?1!832��iQ�J��gM^�b8]q�

���`3eGl��[Wl�e�]�� 6"3��%@@F��A
9��v�-�-�R�.���P��T �@
0$-�$����*Ԡ7+�T�@�9������n��|�}$�����7�F�II#}$o:H�I�$}$��I�#}$�����7�F�H�I#�$o������7�L�����7�F�H�I#�$o�����$}$�����#}>��II#u&e=X�V7@J�0�fd��vRm��9m��@����ekti�WJAp5.�PqW;]�]���f�\����=����C>b�_R�e U�ZtJ�T�ˬ+�U��) Ke�p`��{ ��Hܱ:�`��^��*�`��=�>|U]�*�U�,4�Uj
ق�v҂
��PlUղ<h"�`	��[OkU+Sm�q���O71!Wf5��7<v��o��ϙ9G��I��~��Df��%��VTM^e��t���x�5�4�mgv���������=��x��m1�v�!������.����ʸq(	��䴵�ݢa)�t��]�f�:m�O$,�X����1�ZE�48�k,iM���Lu�߯��{a�3��P,��gf��N���'l���n	9�Wn���Ü�z�ݎl9H�Q�{&맄P����yݦo���[!!�Ԡ!�֙j���On�7%1ĺ<շ*vn�O�������*1j,��}�������s�ж��ٞ(Of��g<� oWn�GM���vz�����������2��g�\�[[n�q�a>W�c���eX�.� �l��Q��L�PU�*�������h����D��Hv��|M�7�츋R��LT��mE�����"!/������>oz�
���d��_K�bU���{���I��ؽY��=�����3A���sC�Hz�[�O����Y�����Y
j�M�&�4�kW-��k�����d��&���z��k=�f�Q�4"gjQŶi�b�̢��K�y���V�h.��*od,R�&W�[2�z|<b?�����/���T{Tߡw��,��F���Vj�A�MD
N�HuYopwNc���Ѩ�ӑ�m�z���4�,���&��v+�6���y��pj�`<IG�M�[���6�q<Ds���3�;�=�8��W�M`�.e��n��~��c�ZF�>[����}6���n��bL0ѫ�Ef^nZ�@�S�yψ�P�k��a!M\��K�����B[Lc�<�zk�78�I+�[����!�`@���
�)K��rKi6��˞b9��f�,��6����k�;wkN�;d��d���G�B�)"���uB &��Gd�"��l4������9� ��֌@��s�FKk�;��B�~��e��-�j#�@���Jiz_J��\���n!{�~|����c��G�嗀`�=���˥�ٹ6�\�7A��Z��
i�&]�l|��a�� $���d������4�e�b�mHiaeb�)M�.�+���eK���p�h����v�knq��W��qût�r�0�0u�k7�z�I����r�3�J�^p��ƞ��qm�%�7<�Jd	v1-ՕKJg%.�6зF��w�}����bPٔ�f-������Ol�F�b-�8���|��v!����6�:�&`m� �le6�P�X��MK<cWq��l@��3&J�알�C-M����k������7J
B�љ���6(Х !e��K��u���]�Ͽ�<χ�E�6�D�)��/[А-�3M��n�1s�G�5�0o{6\Ö:�2������1 ������w�xK�l��x�z�L��3)2M.�X?�Sz� �TK���ϡ~y���Z��"ڿ�7n	�@��[Cr�y̱���ӎ�u	�vE6DW`k��oo�u@�l�ۀ��Pe]��5�i�ML][�����a�)mi����w�����TK�E�mʄ�`�l�RU����ۖ8.�7�|���â���v�X>�s�d6��Re����-ط��I-*�֐ۖ�A�j8vM���]�tvCd���g��N?r�矘���'N�G+Џ%���M���px:��ǖ�n��x���Y��P�utf"ۅ�����|��n~W��y��������q/}=��s{���k,�a�%�\�B�x5�2��ҫ��]���B�#a�����L�uX܄A�C�Ab�ST¥0�;0���������q�lrcd���.61v8����c\��m�dR).d4vT�պ@�/���Y�R��݁֍�%�Mz�h����h}2m�q��s������X�^<�Ӿ����xﮏ�;�B;��h~WlnDާ��޴9\���:��h&،�m���7OocXRQ$X>�����������L%��hB%Y�K5�K�gCb��Sh�i��F2��L摏�vP*Zc�&.�oJ�ޖ��=��+����4�'��c޹�eΰ��tP��=|zІ�.�$u������%Y
��<I��+��5f�w�>��W�v�ݥ���^
��.�lo��!Ԟ5a���|�s�nZ\k\rذ�rfS ��^�95�7\��Q��!�#�OJ̖M%������ɑ6�N9ǒ�Y���/;��r�Gv$븛���R�hYF�=�1�ev&���msf���,�����/F/�����\��c�'Q'IGu��cѲ7pk��7���X�u���d�q���|4M�e�L�O�y���(F�)Z���d�Cgܚ��@y�<L�P.��\�Tȯ:�M���%t��A&IZ��ۈY ��J�aX��!��	5��7T*�}/�k⣸�� �:���e�ʺXh��O����-��L6�.����|4�E��ؐ�/cRS4�5`�?F[a٬X�6�l ��mZ��ƻG:���*��7v�pʆ(U{M4�A�RS,V/�0��m�H,��E���V������kew4��G�Ty�.Ɔ��])3�����j$��M�����6�oh�S��r	;q���2L	��2�@J5n�Q0�|�#C�L�o��b"P��#28"]��m޲����|:B�_þnM<p�u�1�c���ލ	���}��F�ro��X�][�]��<�z�&� JkW��^���E��c�h!l��K�,��9`���2�q�>���������V������ՂCBO���S�_�-�O[=��f+{Vc-D�K���C]�;2�z��Q��7�FW�ְ.�їMM��L�%!5�Ąm��h@�n���ܿz���	�pu�7�Gwυ�c�
8�d^�]S+�y��7����|�+l��i�L�y}�)fֱr
Y1�u\r�a�y�qv�ӧ�_M���2�p)�rv��|����'u�/�������SO���<��@�l_�<���^�ߛ��%�����p�`붻�H�Z}�k��*�I� ��u�u���q���t��Y����%[��.�/_�ф�)�t��3M��r�J�Ŷ2M����A��� �u��n�x�Cݲ�k��:��#.#��7h��`�;aw�9_�y�40l�������_ga�ݩ���г~�O{A��0�1H�NZ��\�������t�o1x�M�i��禀F�T�Q�����o�|{�?&���.�!���˟�y��_|}p�0mjj�rhkRPȀ8�R"�P�K��޲�U��©O]�m�z��AlU�ۑVā��)�P��-<b�4�C��Fv~�S����Η�Ǌ�J�+��A46؛��g�}=@�3�F��k������7�|��TO&�����>tn�J;�zH��ǻ���>Y�q�,.Zf�HJ�<t�����NT��4����Mg�M�S$ZW����<��x�oºf�(hϛ>�}h%�xv{)fqJ�v��;G��vcu�TK,�����{�$����n3iJ�i��B��#m�b����4в+D.�;27�H�lK�i�@r�P�B�cJu��"FSS���I��ߏ|-�<r��ݸ�-�����>�`~��>��ɗ��Hۭ#7^3��齃F��?>������'���#��Υ+�&�0" �.<轻������l�4*���=�}�tv������f�+�6X_j���(�29HE(�����n���E�0s�mܛ��j5hE�A>ڰSZ��+&�f/C�wD�nnqr .�v���X�>�;8�3�]�L�;��az���@ˋ�ዢ]�������>:4��C� �&	}��^���e�qq��sչ��B9 ��]�T��2\�I�Y�����}���roF70�n-�٬�fB�61�ݩ�8��x����|�=��f�pQu���Ƹ��a3���uM��p��a>W�y��.J�չ[3*Bo��Ł��?��y�P��rWf�6�}Y����jݒ̸�e�T����6}�w�x�����Kk,��hF�qd�S���� ���|>0d?[�_��\�'q��S-�Z�gVd�pi�>l�7�H��lQ�s��w�>s��9�T�m�
`f,��������hV٘�fv��P!������a��Y�姢���L����]�XM4��[m ��4�!͹�e�Vf+vMɡ3�==Ly��q�z�e�Y�	P����������?Hπa ��6��t��i�{\���Ύ�P����v1j�6� A�Zi�6�n��,ѵ)����-bF��!�9�f�3������kH\��)q����@�h�a�9*���%�6� A;����nr���fl�[H2�;4�t,�mʹ�<OD��������o��:����%�G���� X.�I-f�R̝+ u��/�w�m�8��^<���l�9x�a��\Fz�Z�dcddɉ�r*T>!\N贱�b�2`�����e��n\���n�;�=|c��7}X��H����ĵm��Ƴ]a�L[�ҁ�T�9�a�%l1����L�[=MU(��53Uir7L�`��%qj�7lj�I���jX����{�����0 �0��W5��ln����ck�#q��kP�\�,�u�ͪ�l╎��|i}[,@��Ү�lt�ܸ��0�h�Pv6If�Y�u9Ҥ����d�k���Ii$��R5eb*�"f,�mBk��1��jP��2�n�s@1�c=���g[��5��Et���;����v�\�R��:jԆ6�8��̚��ٽ�n�����1 \Jh@2cY1��v�%5�L
Kn&F�r�\� �f�r�JL5W�g$u����3k�d�\�g.�4Mh�n�l��+T䠆�b���ɭ�WaӴ ef��v�W'v,.��	&�c{:�3R��コ&y�Kl46���Vg�n�F�ݰ�ut����H{K�w0ps�
N�=����)w9��b&��{2�淬��t��hJ*�52[����4t�*��6D�)�օ9�s,�Y\���:wt�����P�LZLҤ�'yWwN����u�$����}��c�uuѴQ�բ��J�^ 	����#���$��m���{�e��Ck7l^V\h���ЦԔ�[t�.�vH�(Z0��Zh#\���CqIe�'��g�-�bWkv�m���	�ڎL\���=�c��iF���9ؗ�ˇl863ub:dK���p\]�tvȬ0�ji�2���Y��Hq]�r�<�'G\�����=`<v �lnE�a.�\�
b�nf6�i�i��faE�E�a��4�k��b�L9�ٙ��R4��GV�u�q��,LD�r�`\a�뮶�����J�-�q���[�}���|��::��~���}��,�����@f�
�X3=u/cbSXa��
�Ocա�̮pLcIs�f�J[�12a���h1�]��]��ujݻs!a�AaG`8��6�b�M�.�ļ]���X��1m���dwk�i�cs�b1�4�JT��	���ˊ�׉��H�������f�î�i6��1���X#�J���S
俣<z��+p1`K�[�{>�6�u\�A�C�"K3�����*�M��5On����2�:��MrijlKF�1��o4��5���#;��eAT�`�<�۞'r\Y���7|���\s�}��U]���
�����s���p����9�'
[5�Z�i5��B�Wx7Q�z6��v�~.��<�Q#��,*pB���4ԝ��2:Xj���8�L���f�4]5��K�cYu���65����{)�tv�Kb�%�����)�τ�M�AM�y��/'�Kg�&̴,�U���G\u[og�#�����Ѱ].Ε&�
�7M6Վ�%K$eetE!J,l`�S��$��|oϗ���%y�|�fp&<�%�;����u���i��� \�.6����,����Ϡ��v���j�����\鈅�Ek>{o�fmG�"�`�q��N'4c��K�tH@��hpcJql�D�V���p��@���q��B�Js��i�!�3B�,dM�"�)ǵ�wg�8HlX��n�1֤����Μ��~��,`&1(���:N���9����.�l��$�,�66t��z@e��C,Ļj�) 2�B[�&e&X����te+N6��t"�P/(Fk����H��Y����uBW0�\�wB],f�-�=e�[˃r>��Ȧ)��c��&?�\o�v�����7��a��f��"�\�ZnŃ���qiv��,ۋ5�[c�L�,hڸtĺ!��:Nݽ��S�\�n��;���#�(����׆z���c;;�|��~};�������5��#Fo=:n�կ/����3�b̬�)�[���_���^�^����Fx�R ��@���}�V����1ia���W�y�^u�C�"B(9�:�O1[�;�y���WWae�{�Bz�Z�P� h�3+t	P/Qo��83h����.n�,j�z9� 6i�wIx��6��%���qU�h�����q0� g����ξ�O{z��ҝ��)�U��ƶ'��p�4�Y�謲�n�Շ;d�j�7Qɔ��Y��ƞj{�sҶ�������o�+�zb;�'N"��3	D�kc��e�w��x��e?e���$[����3�� �z�?����~kJij@��K10�Of�ł�'�����-`�Ŝ��uwZ�S�H��U�K@2Iݛwz��A�9�v/NhU3��C��B��wSۊ���Z{wc����k7��2n{���"���ͬ�N�XJ�ڳܪ��~�*��氟!p��D�m�d�Hĉ�x�5q�X�,�ʳ,KۼY[�HrՍOy0���DWX�B�� .e������xh�:�p�������==�v��d۩ג
'��z{z�QK`� @I(m��k�?d��h�`xY/Y��Ǖ1(��/��ӯ<MF���>�u�ZNz�~$��a2S��[���f�W��cZ�ӆ��9�����}���q@ڡ����~����|�������$� �~��{(���rܕ=<k������V�G���,�1Iy����R\U�,�-2�.����H+H7�bENIƲ�m1y~4ݧ�@6��5���DWB��mn1��U�R�]�u�%W�dv��������d�ֆ�afs�B���P�Ż����xh���q��z,��g[����,�yX�rF0�"���m�����Eﺽ�RCw�86aj�=�V�ٞ����6ϊ��ٸ̗���j���_ �K�o������{o�Y-q{�L?H
��K[�iړA��9����;�B۾��\]�b��}{)�e�:��\��]ށA&Qj��K37^��C�Q�͢5m���B�~g���J�rwŲ�c��QPz����k�8����צ�5��5��^��Q��E��~��2f:��Fb1�v.Ml;'��-6-��?CФ&Ĵ$��8P�W�=Ϝ�"�8����&���`�P&�`�4Qh���g�xl��ۗ)�+�gg����9vg�${���an�~�)�C�����oӼ�{�4����~/����g�G�I�WU�#T�!��PDƘ
�lX�l\&
	�tt�K���lv]5�k�E=��]�k]򟠜�|���g���U�f3w�dKm�Cʂ�]��^֧�qv��r�r���j>b�����(ml%_y��/oG��u؝�ڻ�t��`���>�,���nw���{�]:��B�Z@������j�y[O���%���e��i�L/ٴ+$�^�S�m�f��^��h�K�z��1x,�B�N	�Oi��u=��P>=[˟�����3Y���RH���{}�z��72셇���2{�Ab��[b����?��6�M�u���Rku��;tw���$\u��k]w�y��@�߯��[Q껽G
����}ܽ�J�E�Ν�5o���B(���w�{@�,�k���W��&�)��g��~'�g턷/��9��o|/��k���������G��CQ�i�E�t%�禁�E.I�Z�-����3��ul@pr���Rrβ��,����6oS��hl�0��j��3�6N��Ќ�
B�9�Ziն�-�0"w���f����L~r���n��6�k,�݈d�jM����#7;1�.�5eox�5�p�%�4��sCp�n��z�.a�Μ������c�+���K�g4��ΈF$�sV�I�v��{n����b��ޚ�A�]����Z�pɮ��H�<���h��ZQc�w�y�GK]�*"�!���0�D�9HQ�u�����RAv��w!�<N��}�%�)>$V�Q{	��qBO̎�Z��}��;�2�.M�EM�õF�m���54'��S�[��n�E�B��f�wYS�,��!#�b^�9׹Ն�9�kwjVU:��%퇤�J�-N�Q�М@�4oh�w�r�ftݼR����x=�>����2��y�Mٺ��c�<�sɻ����{�8��9vN�E�v�\Sr4Os֞DЦʤ�"C.�!�D���//'�<u�{��8��s,w,��m��!pr�#�����	����[���ݎ�b��ol�9��4���vsQ�.��+uq���?���k�d�Ѷ�tKj$�;s�40	p�J��hݳqiy�x^p��%��p�i�.�ߺ]����^.�����mu�ĳ-0IVk�h;?
�2��j{��y��}ݳ{���6�꼠�/;J�BҢu���s�����}P输�_�1�A�ͪ�g��@��uy�]ױ�Y��w�:^^��V�ޠ=u���6RCW��I좟��z�]�mw���J�<w�y��s�[�=���'��VY��t�8�:��h���f�16p�""3G	�n����&jvw���m�4���έ[�'_���7A:��z�}��~a�u��m�Aj9��.��yW��k$��l[+d]-ݰHɢj�n��Z	�4��b�8F���	�i�����z����gW<:r��4�hX��=K�x�����T��ǩ�<"�S�vz�Yu˸�;��qkj��}d�8��RO®�hmQmԥqjM�b	^6Ґa7��<�>5=>;^-t�ˊ̅�0.������Kz�z���x�Qű���N��s�{s�~���%�����^E��W+�~{�{~����K)$��9��l�U���s-fz������{����o�v�r�ȮWi��ͰwY�{Y�.U��z�5;�X�Φ-%�xK�����J�>ѯ7�Eg�H����ݮ��т� K^�g����ꪄ쵷(=�,�c0.D��n����nݻ9�kέm^�\o3j 9�a���{�E�d
�M�+a��f�/f�Ԍ���t8��0����E���Y`����M;��Ϧ=;DW����o3+v�k�e��тvS�D���O�d�\�,��`m��{�!�Kk��y��j��=�|ҹ}˹�}3/ ����~'y�{r����o2ד=��;��5'p�p��x��NPv��%e�Q4
�j3;A�`ؔ)�f����<���<�D���C� ��DD��׳Z��{y����^lo�S��^<��?`<��T�\�i�%�BfԔl�1Z��r"]���ʤ@^��L��}�&�sy��i��ǫ��C];��Y�^d����ޣ�u#껺��o���=�v���m=�
Y(��=�Iw�s����s~�_x������R�����~�Ѳe�I��X; xo ��.��Uac���ދ�w���6����(r���y�����������Ҡn~c�?	�Q���	�*�ͭ��>�h�u���+7  y���y��^��C��u^��|(��n$(w9��y[ya�[�^iV=&��NN��緫��ouk�מE�q����������G|�d��'4���mB�skL�f�`�|��xC^Սv�KGf��wH�����?��z�쐬Q�n��#��d#7g6��f��.�	#v��X�v,��H���b�c��O/,ܧ�k$���y6sv� s��=1�Y�^c�{F�]�.��-j��׏�Wm`������CO=�;��Y�s<�_>�o�_�^0��m�X��ŧ�����dWx,�J�����]���w��X�I�������Q���xu�W[��)~�SyN�r~�=�7��5tgRz�ך���`�YKu���;��z~�=��>qq�l,�
�u�0̂���&�������2�s|5���{�Z"����y�ٶ7�� $��e��;�ȕ%��Tk(��҃�KZ]��T�a�'AZr��Q�v]t��e�@4�gp�jP����#�S���m{.��{.� �۬���q*�}�w�q�G�|��r��Wz:��7yHg�|.k�g��ެow~��6�����ϰ���qsM�8��L�j���;CF4���1tJ�9�+cu���ÑO�7Qhʬ�{�.w�זm�M��|���ͣ6�5��<%����.��0�io����ʜ�9�<1E!!Q 4����m�s��E��ﴦ�-��v�ï�ɠ������M�}k�-W��;���Ԯ�k �f����N>uZ6ZJ*�U�Cn~�u�\�vdWy[����ɇU0��=��|�=�����{�f���s~�ZW�m��\���7N�m7��ۻ׻}L�B�ӓ3j�7�{��n�#�@ֺ��}블j�]����ڻZ�ydr_=c�A ��Af��Mz�[��s��<��ܻ\����b�K��O:����<�����yZ��ʖ�R��,��ȧD��V�G�-���t�4d�����(�^�7�z�fc�ܠ�3���躥1/v�>w[�����c�KWG��M�ǭ��+��CeU�W�����f8g��	N
�&�f����3�Bc@���8�G��#����̺.��z�p�:�e
�#�J�P��3���cf�)`�6��m	�$׉uԵ�ؗa �	q6*�d4	�fk��-%�Q9ؖk��zM�;����<8���x�U7�^Q�9�o��1ی��`7R�ف�k�Qnt�3���_x#^��s	-h��K�q�ۛ���gL�X$,�g��Ԍi��V�h���c��DB����h��w;Vc�pw6�m<�k�-��1n���)���C5E\�,6щ�:��&)˂���V4h���f{w�)���Ӭ$Kn���Sf��i�`P�}��O�f]xr��������t�ꇻ&����{�1Y;����Ja�pq��ע�S/:H-Y�Q	։���S�2te���;j���\ӫ��9����������`�j%b��K�'�γ�������iwF���+�������k��nml����~N�ms�!�����]W�&�M8��%P��ug�	��B�@#�{�N����{睪�Oy�
xNܸ�{�:�9[���h;�V�K�<-�b�=�w婸�TnOD��X��,OOd�+���p��h:�tV�e}Vx��Z�X7�5m�9.��殖�}y}3'�N��^�^#N*���zq�n���T5���b�E�t��zcXI�݈�:wM��o�*#�gk\�����RG�A�V�=�W�����m���ĶM�+�nf�d�,� K�����YM��z����z����E濂��WIr�E�M���/UB3�9�����9wK$��YP��Vړl�o�e�H`;����d�W�s��,���ܐ�S�\l���>�x6�7�n�'��lu��;�uBj�f�{��{�=��D�8}A3��}�1@ӊDl<C�m��d��.XQz�-��^�����E�	8@��N�E�6j��������{�;ص��0��gi�	7�޲މ�����Q^�]�c�Y�����;�&GP�t��F�M��Y�Ë\SDÜE�K���T����/�<�V�"�6��5H{��y�9��Ŭz�k�sf�|Be�c[r�-����m�94��Q�2M��?q�O̮�bl���=&�l ��?X�o=�.�z�ZZЙ����ʅ��_Ɇ��*�͕R�ە�5{���I���_��ײ�r��m���X���8�^����K�6)ܸ��3�*9â���md�;��<ݦu����U��\%�}kWn�{�b�;ٓjE����cF�檝���k�YӸ��h���T��i��ԣ��]0�1���w[3��7Ӷ�`lGZH�r7�u��Vv m�v.ls{8����QU��f��vL헳�5ڢ�0��D\�/۾j�[էY��u��+AE��R&Y�{)ի�Ƞ㑕�&(��)h�y���o>�&>u!��=`�Z�]뫴;��7��2��i�Q�3ֽ�9�q���^�]C���8V`�vs������[�Y��%������]�
#0�A�� �Z�[���SsM-��wN�_�8ko�*��Y�ٳč��W�ё �����;ǜ�+$�[�O�9ia�<!�Xx��9lWsx֮ SL�F�,'oe��Dh���/72�f����u�ɝ����]�,����&m �ć��E~2"+0��c]k=kB;,���^TW�lDa3seH�%�����w
�vUa3�ާ����H-�h��t��hǳ�:)oM]m@��Sk�t�ʖ�, W:�*�D#e�80�f�X�\J�kB{:��t}{Cf��*�։���l]B��:i�r�g�)��7z�ft��sQ��Kq�[z�kԕ+����z_P����Ś9;��o{���zcgL _��r��#OXMe׶S;e;�9�<���+���L�<`���S�W1.�����	˦��#�?7�?H�}&��i�~ݖ&�Z�f"�3{\{k�����k�񼼺�.��Jl��x\0F
 (�>Ϻ�G�y���k�o��z�����O��o�w�
Pr��A�N�H}&�q�V���)�toĵ��R��iY
���. ��%���HGѭ�>�o:�}d�FO��* ����#��ȹa$X�n�S+�7�2x����1z�%j�����ƴ�ROD�kVp �wd젺��7m����a���fz�Z=�0�4�|�[�HN�j�\KS�9"t���{�E�`H�o�p#��@}d2Q�G!�wb���_��?���:ێ	.���ز��?���ba��L``�'H[v��VDTĵX�J���8�fM0�-��o�fy�E���<�!���[0>������o����Ӏ8�.-]�$|O����I��I o_!Gӓ�;�MP�>�; �L=`�����ğ�O�]z?�����6"��.Pf.��Ql=�Ȁ0�эY* 
�8�:u힧�>Di�D#����@A��N|(�>��Ӕ���\��3D�ٷ����zV�1���1e���Es+�^Yr����g�ECWFCQH���DT4���K�<������M�ݣ������o������~���x��o(԰��4�?X�G�9��~�ʯQ��D&��>|4�ٮS��*4���Z��q�iu�|�e��Q�!I�	J��Q��4f�t��`����ٽz�	�>��v�L8$!��q����ȩ����\��+�@t%)@�@���B/��Ǽ��ݕ�W
��`�j���u��[EX�w�7]}KtO�\u4�wE`JYٝ[W���[��ΫV輩��*wʺ�L�����bH'v��L����GcM�A�\}�~`� syk���~o�����{��\h�<!�\{m�!��c�L,�xz�����+Z◅T?���{��qE�>��"T���2�>C9���d�Zzk��ۿ_o%;pgd��&���G9�COO����}�k��WhblD�3l�ElF�l�֗j�gI��(��ba��bT{���Qr	����L�{�qzH��}�>�w���^�p�N�P�{&G��"H���W��t�&h+^��#pG�6�{��6��Uv�'�'�������D����^hѬ�c�&J�Z�\8@)��LDLyȊ�I��4h�"Hb�!�ڷ�zϑ
>G�n[�[��$�K��$3Q��ԃ�hE�7 �\�M�l�| }̍�K�.���ީ����N�)ɼ�d�׌�)�<$�� ����<�נ"4���.F�DV7����;Ս���_�`��Y4��1����ƀ69X�o\0��>b��ro���` �"���������{�#����o�&�ڞ��U*~���|�ōė�d����0� �H�D�&��d�J�O�'��<�O��4�#�"O���S��7_W40�aTfǽ)�g���B�Z�ٯE~`4�����\i?��1� �9Z:���40|�-��}H��d�5
�Q�Ԁ�>9>t�"t���$�IN��ק7����N��<"O�DA��8�(���y��#�T^=Ǽ���|,�s{O��"�8�Q9���a������Κ2TE
�˜�[
d�S���1�%�Ç2�	��$�[��5��l���ƽ'j�f^�[����3�32��U�#�r�s�W��n�p�/�[i�+ˍ�Z�H��RǬ�<=�[=��n�b�F�[
.�\`5�Qqh�k�R!��{K�R�&D�]�������\�l6w8��` �im��ۅ��kM�I]���nN8�q��mΰ����r����q���[Ȕ��;#��q�N~B5`�,�N
�Bb�TH��N5�a,I���:9�?~����ک-��6��56�)�ԁ� f�Z���{|�l=��Fښ�क़W{&0�f�m�h�Z�L̕M�L�hZ���?	�t�������O���������O�>�"H�_�t�=���C��I�C�S��N�	w����LI6�p�4|� a`�F�@p�I�Zȗw��8�>��Qᇼ���A�j����~|��t�߶;�>�:|88�|zLI(�
��N�;�9�D��qp� a���I�|�z!�e� #��|;xL�cǽ� Ln���g���Ă}�G�9���y�n#ޣ� �� ��8�	>� �`0�0�)�%@��G�Yp�� l0�n-�D��(�S����>�=�"=헸f��%������\}i|҆������ օĴ�A"G�c�\��(V�{���:G�w=0˹D��S��Q<��7	�熞�*����?n�K�-�s�V��f�DY��V�e��8>�$���F}m#Rj�i-53w��U�E�O��k�{�l9E��/�ih�,�8����{5�!ɑ��#]���M��KI��>E�M��`��e�m�;��E�l��ӛ�v�>�Oݵ~����K5�Z_T���X�>�{�">�l(� A֐s��L4��i�. ���-�Q��-��ɠi�� �#���#�A�8����0�'�p��٭���@�ȕ.azωD*��\��o�y�Ԅ7ODET\�s$��@�x�#X:㵮<B`E�!J���iK�4� L��X��rI����������� �0b��n&��iI�"0��\"�����t@��,|�zHkO�9���a��TY�T�@Rc=�:@�\�!S9��@(�%��!��x�M����
!��h����ڟ<��7�!��-���pDm��Q���-4�D[�<S�w��v��]@��i�0j-c��W�&����69��:vΔ#
]B��U�w� � ą�S�鸬�ʢ G�|��ӝT�5�<��	b0�� S�'��Q��Q�+�x��D�p���%�4�|;�E�;Ϥ�hE$r�2������{���<l�*Z�T{O�,Rl�c�v�DE'km{)��DI������2"V
#O�����Y� V����	�v�^������ݘn8QK���7~���Ʒֻʡ]*egb����/p�&�$5B���"3�Q���}�;�*����t��Ͽ����Y��$�0!�0��ȳ���
����\�*;cz�My�D���;��1l=�{S��[j�i���o�[�N�R�j�Hz��	"K.@v^z�<�V0&O��ȷ	��a��P��*t��t=VH�oa'�DS>E�Z�,���2ofD�<�[+Ћx�"ϑE������������ٔG%�1�i�ņhy�YG��B �4vt25h���^F2�m��d�`J?��܋McX�o���$�K��@E�)������y߫)�x�ac��Hӧ�zT��/U��m�r[y;0�QW�t�8� #�M����C�R`�p��9�!"�11���݆�:�΁��t�ɉ1����{a���BH�"�h�$����!����x*j��aE�>��R������1��'�}6�@���#�x�v�Y}��F����#�p��;�MW,��������x������� j�A�,1���(�Y���);�ɼw������s�>v�twz�GA�'�GN�G��<���-�VѺѼG�;G{��� �i�3�oa���9��N��Ȯd*��z��Q^�=�h��>�am���q��Ϭ�q��`K.��#H�>I���[�$f�i~h�"Y��fhwP�����z�0Q�T�Y��]����,@�<��g�z {��DL�Nރ��D*�(����v�
"]���T8����L�^5nv��w����o}o�n�w��~c���t�m���-:����X�M9 �ؿi���8d�]��SY~M{Z&pi�S�<�ǋ�Xn��$�0y�ם�A������$��=Ԫy{�,�9�	�;��y>�ř�}p�v�Y�Uڞ;
��[�5O�UL\���2�h��p<����6�tQ#�Jr�Z��~o��w����{L�g�8�c���-Ố�K�M�g!�d8���)���Ï����by���
����^�;���i7�X4��sˌ���dy;7s�ݯ��(�a�Ys��?�	�}1��?NI)?�� K!����1� [�V���5��q�Kc�U�� q�l�S ��'�W�czT	�x2���E�4�-x� I�	}3�l3Z*��0?|�q��v��?i�~����h�Q�>��n[L<>���Q�>����y��n�ht,A`�#u��M�
�3��@��� ��n�W��i�\k\�_�b����>*tj��9!'O-����"�[Nܺ��\�L0����>i���Ŷf�G��x��C4�v�8z���6��� >�t��:�*�kՉ�XpМ�&�9�w���;��#[\m�D5�O(4'E#Gs�����E�s9��h��Y��4�X�>5����o���z�|ff5���t��/��>���� JdY"Π\�r�#���%���QCct����{�.�ϭu!� Y���;y�0��A/7Z���7��6�w�9�Y�b��G���$�D�����ׯ^}9�grYұ�l+�6���8�ŬZ$��Ջ�W�i��^%�X[�#WAn�L�k��'��D��׿��=�@����?�Q->�e�c���"��81r$�_�X��W���L	���A�P>ih凢��B2d�#�f$z����`�;�<㵊1I��/i�,�c��n�c�#݌�j<���]�פ�����E�g�t�6޹��,��S0�͸� �u0�*|KqDx^3�ώ�/-`M6x���ޅq��Y���( �E_f�G�� |�����:�����w|ޒ�\z�%�<}/g��Ll%d;�B�lT����`�d�/8>��Ὡ|�u�K{Θ �&�#�⧞Gn��$���<}g+"�'d�T�~C�Z}��~��I�|��UY��ZH�4����1�A'O��r�b��R�eL(�I>a�J�6��{� /�T�N� �C(��Ǒ�F�ƣ�
윏JoQ����A"O�S��ck��sdEmAS� ��ȱFO��"L�	±�xQ�8�@:C�A
و��9�>�m�oz��N�e�P��49��"O�5�T
>���u$��u6w����zFR�$�I����Tn㶙��iؠ�`\m4��p�Z������t]�v�<s�w���3oU����u3�����sk �*U�;�/ױXQ��gu�Y��F�7�����_B[z�P�ٛ#6�ףO\�W���7`�dK�gm%�%h�l���m�����b���
0����Zؒ�+[�m��bu��.)���@�Z����m��͈�Լ�f\PT�CC���[^�L���M*2�?O���d��N�ğ��χ�ZK�Y]EF�ke��m� hPq���i[��[�k��Zl��,�ft{?������+fѰ�Enr�ۙ�i�nԸ5`a�/��`/b�6z:8t��Y��x�w�)J�0����Ϣ��f�y�9��5g�U- ����(@�90���z�
"4����.$�; YF��o:��;JF��9�u�����8��ѓ�{��ޣ�"5�����޽v��q�4Oj+��i��)���Yr���6|�=�5��l#-YKw/l�7 J����|�6�G�CX9�"y��AL�gg���-�H��3�Ec{�:��>y�{dI�֨����}ޕ�����3w֔be�����ͮ�!�VƟz�,0�0�k�P#�ނ�G����f6��4`�Y'gfw��xaȁ�ո�;s���"�A>���-�#f���N2+�H�v�ߩ��������3�Z�������%����yO0Zp��d^#S9�#/���
]�m;��dA,E�~�xvj!$i��1�j.C	�2>��ΐ0��`�8Ͳ�Kϼ�����F�a��@�*Za�7�!-�`��n�[��?I?N��I������n0G�|��[fDD�f{�yi�k��+�^�
 I�T�}�p"�R,�4��b�s㍖�ط�u��oON5V8�~�m�o�{6����Պb� �磗���;��X��2�J:{[rM�[I�81���ܛM�{���������@ʶqe K�<�@�[����}��*�P�>�dA��	��TX�{�
��f�ǧwM}�`�v�o1�.I3�\�&�Y�����6E�!�x"��vHb�.�����}R�K�m�	�et%}�ND�xbH�0�?@Ǭ�~�,���mX�1Sn��v���m��w�X����+�-mg듯�z�w�xa��n����x��h�u9�>��d�X�>�m����|�S�0� 1�����,�,�|8�4�>��������Y�>���o
g-�[_A��fm`���"}��P�u�V(��,Ҋ����4_Qs�f��� Qӱn=���LO��������<��dd.Η�	nRGdF�h0G���|���޵t�-s/��׼��s�Zw��:+R�0H"�s�cz���&�`ʇ7�*�1��}��� �#ҘQ_n��y����T
>��q$3ʅ ��j�32$������R�G��V���DQ� ��1�~?ςw��{��iS�k��G�����q'�/��M�j�G��D�'��� GM�z/>���p�A������\ A��WR|�H��0�"9��T��Ž�y��I�![ٕ�R�f��������,=��=�9;y9�d�	�~�n�,��B��N�18*�
ynD����%_�ڏ���Q��h�"�\aEN#���|P>�a��"
a��O��9��en_���e�Ϝ���aǭ��[z�r���Z�o��œ��RI*+���;��k#��	 a٨zA5��cz�V4����G����Ժ^ f���v�&���$�0h�"z��|��(��&�Y��Ҡq��������/5}q'ѡ���d�#\�� �d����uzH��� �f���sÚ#���x�����$Ƀ\ʈ�����dGe{vV��C�~�9��fj�{�z����,-�Χ\���;nv�Y8g�:�lCP�w�is�:eZ���<ӓuQ�b\�c����� b|���L�x1�j��(��̑'�^�D�g�1b14�K�٩|�l%��)t���=<0D�4L'�v��l"H�wJ� � za� a����#�%��lxq�o%˜����t�E�z�!�����ns��m���Iv��xx����^�^�X�_���ow��t�UJ1�u@Q�����Da�W0��� Q��od�c��z��FF���E��κv˅�#��0}�	 mGc@�	��0C�Q��7��DS=]nHd���4� A��y�O��/☔��A6�&3��Ce�U�qf�met�GV��+"�`Q�.n��ݻJ9�f�vߒO��?H�L(�>��vm��
,W7�v1�|.���A�<��q��M�6�|�h�5J�f�\�A��}��Ac�-�W��#���*���a����Ar����cP�Zߞ��;����爛?O�T���A��M[;?.,/=x9b'l3���V�E��$9ȃ�	#e�i��Yv�%��dk�!ٽ'�k�tɢ4�+�&Z�5t����q�ß~]��D�M[J���[}��s�D�,Q�`���`�:��l$��x���`�7�-���6�o9�"�!�P�w,� ,��o��$�t�#!����+Ԁ�	W9o���"6�i���iq�_��wgf���67#���/=�͠�
�m-,��_�dL5�أ�|4��AY�!������H{)�.}f����NԼ	!y����|*&s�5�Hi�9\�t�b)�r��w����X`hWUv�M9Y�/�x���ٛ�k�7�F���T�c�����!�����.�η�d^ǃcE7Rß@"��ۻ�������C����N���wm��H�"S�W��j||%���[q�K,Ċ!���m�����s*��l�R5�����o�͟ǽ??����~8��<m��������������v>zp���ð�h�"�b��9��j��n���~���y�J'vq�\$	��6����51ۥ@ځ	z2��v��o�������⧟oiI?C�{���R��������~|}�INB��l��$�~�����	$�h�L�6��f|olÀo�Tx��:Le{Lcf\9���X�Q��R�=D�r�9����"�_ܝ�ai;-}{����9��y�?G �A(�rH$i�{�[:2��,�F����>L��Q�-��^z Đ��8����=�|y������;���?����E���kD�Q��Y����iW���]4���%�ćMN�<Fm3��w��@���߄��C���r%�|�����}�;�s�x�a��>w��N����{lpO���a1I����IaM�^��A�����m���]*�^�FB~f�8F-]�� cp?ؚMToVW���JCe]��Ȉ�	�H)(+7�w��;�F+[�?�qػ�͓6�K��{�]��D�8'�}��o�m�o^;w3^���\�*/K�[C�`	^̘��$����'����ny�X�ls��|�?e���r���K�a�iM;�u��iU��b�}7�f�fn7�,dͲ�l��Gs>���ax0q�U�ˉ���;�X��q۴���	۽Sz�V�q��W`��m�n���u��L˼����z��"�lg"��S��꽳��ՙ�8U0��ff�'Z�t���
��f0M�/DKp����㻤Gul_�[��������Z���Zʺ
��4ҶxPۙ���-�[�:H@�q��&���	;w Û���tV��tn��a�:N&;���=��~�;UB6�WNPKh��ڻ�sK�]h�Urm긵���tl��5oN�˶+X�7f$�s�;w�Y����|uڼ7��vS���5}ߗ>�����]��v�YG�Ӷ����$i�t�&B�I��Y�&~���BT8�b�aYJ����z.,��Jd��q�NDc��Wݣ�Yb�-�]�l�'ZK��)��x��f_O�8�YD�<�Ǜʄ��Uu֘j֗ȇY��ts�,K)��oS��z�ཱྀ��] �8dN�rœ�*��'B�a;��4����u����R�y�(/$���p�A�qt�*r��tu�J������N�yH���B���v"8f���x��
�xд2�Y�i1�/�2Y��X̍`��/��&���ꝷ�v6<����޻5����*+j�&1�G��-^��1w*��!�2~Ǝ8��K�V܃���ĕ�w��꺰E�V@4'���?��X�;N�M�����+U��n�����)�L̤.�8T��*���]��fH�0Qɴ!`6�DQ�̦1��Ke\�v�Z��P&Qms�d0��f�q����$���>����w^��<���k�`��Ŗ`��\�ϏΤ�U��0T�p\U2�n�ָ�j��ݮ9L�`S�.��k��/�����p�V��Oχ\��n�rom��s��0o�l���t��jpo�8Ƿό<�7h�
�m�7����;1��$����Υ��j50����u�eTt�v���ۂ(m�D���h�1��D4lҠ�.�-c.�2dmt����N.݂�V ��a�m0L]K��1��&�
�6ls���k��ڂ5F�3`��I���ґ�P�-(���u�0u89�URr��j��=:�:�ia�%�?�oz��g Mڹ�:���PhX҅h��]�J�cA12r�Iͭ�K�Z[EL�tV��]�k;lu��@Q�x�1��a�v%��	m@nTW$�\��e{a� ��P獹�;Tn�%� �YS)����R�/��.-�)4��0��֒�YN���=zz@�a1c�zLr^0[c6t�eN0ii%��&0?O�J�XY��\p
��Ju
&Pjd�VG������!��jS���w�7gf��?Zm<����Bib��<M�OK��n��X�5�Z��+K66*�I�Jpm���;��3㞎:�����8�T3veEz�Vd�"���@�F����G����c�MDܰ�����^�G	���56��6���t}Bj��`�-��i�犷cM��1��.��/�_{�k�!�|6�x����*_M�2�WV0��歎VU���f����.����^�|�V�$wiuܲݴQ(W8�,&�=��!F��ooOw�z̏�v�M��e��k�n{6�X��F��˹9�����4�.��:��n-c�G������:ks��4t��ff�S:"�&�&uijafߏ�}�;�Q�>@��+,!�j�ae��b�4�����Wb��q�����m��N���E��cg;Y��wl�u6| �xu�n�	]���5�$���O��	2H{a��%��Y
�ۭ��7�9�C�%�^�L���Qc�8�D��qe�}��l�'�v!�n�b1+���!��,؊��M&�x�+�wj��%]6Ķ�K�:z��%G��st��6.v�)-10����ٳ9����6��T�͠[\�6[�3���.93��HĘk
A2h@n&���k���=��k,���Y����F^�J�GJDKjk�)ae��V�6��sn�h9v͎�G7�P���yܲDis�2>ng�*F���,�:`��ق��Vz���&�m�»�{u��mT�_^+��wɩ�5O�ټ�6ئ
�:���\}�[���^��F��
����JO��*v���l/o��M�1�Vj��bS:1����U[�[{ع�8g�I�ii�3��g8j��2M{d��~�x�{mW�u��Q�)cr�ϏT��:�-�T�"w^em�2�#86����%����G�%E�`Sm����a]>4��m�Ov�f2�d�V���3�>��Y����',[����WuM<��խ��Ɲ�],��a;÷-1��-7L�23";zy�-��;{�����s������rÚ�<��QV����K�-��;��_I��s;����+xvzaމ�9�� �4ϓ�B�B��qrQ�]m����Ğ�M5��Ǯ�j�w]��)2�IL�"���ֵ�	`�`C.na�kV֛�ʕ�PEK��ʀ�;T����~�߼�6����M�n�n�eK��������շ���d��@B�Y՝	�6��z몠6���S�s[_}�����Z
��k�����}X��*�"�v;{Z-�d]pκ+���0�,���pq3v�r����&�uiY��F9��m;fܝ�D'/��Ac���WnV�ֻ5��ɪ��k��/-�&���j&�ٙ��Y�5r��
���fX]t�u��{N��G7y�r>{>��i�n���lk��,� ���ͷ��B`��rք7��\gVC�Ve���t@G=��Iݳ.W�.��9��9��JX�o6����E����\���������S����Y�n���N�A���N��d;�6:b:�@R�Z��Y�k��#(9y��T��.�e/Ɏ{Ļ��5��Jk惴�׎������p�+�R6�� ���睃.��V��	�;��y[;���;�n��v|,L%�;/�õ��2Ћ����|3�>�u�So<�#7��[���|�g�&��ŦBZA�`WC�m��\�&gq�[�y�۬�iI�v+q,p�Q�<d�L�@��ݤ���[�z��+܍R�c(ku�-��kvw*U8�f�<���<�̲h�yS�]�Le����z�':}ayE�2����t�i��/�j�%s�{s��I��z�se���u�$ ����q���.E�N��4��^��n�5���H��� �%lV,�$wk�ԫ.Eu�f��]@J�p/_�7ܩ���֜�#�w��n˨�p �~��+�!-ީ� ����A+Z�ٲ^��,2��;�X��k��i���ӯayC(�������$�v]u�eF�W#ՕέM���c8B�̚�"Z;N�b�]c��AկFq��4��b�Ql��ZH�)9d�d���CZq1��F�@-8e��u=.���PsD20Ί>1��{���rhR�$�ELT1����#5��: �@�w��CeB����4B�x����o�p�$Wc��	�L��6�k�Mb����:��V��&�T��B{�*��Be�֠w�������u�Tc�a�-�I��Be��r�j_��Cq��y�]�k�b���V�:�l�r�.���؞����%�a�nq[C508�ի�3��
3��xL�mr�ʸ�GM ��Mk򭧸����Wk�sa��4g�:f�.� e�]'3���e�§�����<_g^�{q���4.�V������"�r;CL�/	����~���V߹t���A���v)쌜� ��IB�V����ɣHyoY��G7B�2��6��՜��8D��ol��	�!�d��֞;g�"N&z:��(ְ�c��t�Z�#��0B�k�VkE�t�k�[�9�]���&5?����o���dj��i��gs��o���RAB9C��f���ցW�\�E�3w�|2����k�K>���}fb(��zEM?d���r+�w��6(�*�L�|�C��e8M^q���x����Ҟs��PF�.�� �]7�(�/8n�[��,��Y��~U�`>ͺ��<&g9��֩�oX��x��ʱ�K�o΋0��^7Fskt㰶�S��������+d�-�:p����ط|lL��^ō*��QDO����;��>��K��ٿ;�������\��o!m�۲ ц��a�a��r*i������i���-�I���
t��E�?�&�gT�+����J�ٷ�)k��:�۲z:Ҙ�O^��r��4����[Uj�TM�v�����p(�f���{#N�ǧ�&��[0�;�&����Ͷ}�=��"ۼ��VpO�W�#?O����KW/<��Ё}9�����b�ӓ���NX"����~?t��}'������O��SʹS����o�i�^���4����~�O��Q&�i5gO*݆Y�S���5��"��0NY��!Hĝ2ݹ�z8h������kSZॻ���rȆ�/�<n�ܩ:�Fj}�<�o\�7��㑌����H��YS�.l���G.�әǿS�����LǺ�c�.�vb�����k��"���k���OA��r�}���W�����}�\}c���y�y%d65��,��Q���a!0�/O/z���w�Ћq�v�c���Z2��+i�=��Y��3:^MEޛOyn�,��<��q�@�r�!�u�P�8te���A�)��[��y��ex�6�Q�.���x�[�1���|��� $vr&Ĉ�]+1� $n�5CD����*K�Yx� y V[���ޠy�%�LS&̳l��]��nԹk�M�nIHGWM�ˮ�v��������g�1���@�M��4��.e��.�K ݻk�n���胧��1���f�]I���=uI���m���˓�pqC.G��;B<���ك ��8)&,$��;�L\	�*NW)g�=���w���+���9/����u��לrP�����c��O��켫�����}8���o߯���/�}��p�/�!��>$czJM���R[�oL�]��\>��l�|DY�?�މ���H���c�7eq$�KiO-��SJ,�Hqj��k-���9���|ɧ��}Û�������m��wg��}[��a������flL�)��-�,Y���i�HW){y����w�����t�����\c[�YAn���)Kd;�*<�����/'�'�������Ď�ە0���5Z	Ӻ(3��;�D^dev\�!�q��|5R���Zd�O>�� �������a�G=���-t���W�y��ͩG?��k�E�`�1�ܦ0��[��dƤ�Q�am,cfMqԝZ�b�7k�~�d!Een��|�b����w�{�;S�t˦��41��]�U�&y�h��7uO�%������4�Wר�ݵKRَ�H~f󇂋L�1	�N:��ώt�Ϟ��{�oN�+N�~ߠ:�.~�f�Z�Y)����[�9Yۊ�c�V�>��(�Oe�,Z�o���	��8�>bU��6v���R���J4y���Wo����=��C�OVC>'��'6��db�'��-.^�����1��(�)h�-r�8����P�t��|!��ib�N�z�iw�cbA�Ռ�������	��J[_{���?J�ʚw����Ԛ�ry�%� �HL��زI(����rx�5۶�$�K\��|����A&��C鸒Z�_���w��d_f�du��ɻj�q��&�a�b	lr� �os��t�l^��|:5��"D&ȍ�24C�<5�"wc1�⶯��b����
+U�$�N���Y�nأ���[��ۈ�g����Bq9��H;hU�2�3IP֚���Nhv.n����s��g�� ����o"��x����V���dM��\vc�!�2�ɷ弤!�J�QyONk�L����((���Hݒ��h��`3��8���9�s����:.�jᵥVO'�#��?
��� � ��=n���\�\��P%�.h��B�u�����e?�S���.�5y�]OE�&��K��鮝�5����3�f��>�}�N�q���]�
o�=9�_h�6T염a�e"^�X�ggI���-�[O����?�.����q�6Gw%���}����_��Q�/f[�v�����}dl�K:޼���d��p�8d��.�bi�U	��lK�݈� ������u@����o��䞆�/o�ӣ�^J�f}�k�/^ �V�:��Ք�I��ڶ3��p�Kp@�����]�r�Q�-x/�6��s��iJA�&��=n��{~���gYe|���MA=��P>Ք�ｗ���֛w����J���;a96��h��V���8�M8�f��%�ͣd��mFZ� ��k�=�kfrZ;���F��9S;2�VO%n4;�90��s���k2ɨ���<�k��ѹ�����ګ:R!'gH�I�>�hA��c+�F��h�˒�|�pgm1+�dl��rO�Q���f/�C^b�������'����>x8[��}��8G�sS���rY]�s��>�kG3.�#��hE���c~��)���C�|�Ԧ����w<C*�Zj��q�C[ጺPA����C�e�1�P�m���	ܐ���;:Uv�������[��&q-��w>7	3�����:}$q�S�.���!����M
^]�LW31N�B\�h]]�[٘��.U�v�ê�������&�����$�HP}ɲ�jf��v,�W�����9�s�Gˎ}�7���=mxQd/;�iݒ��N�A�ңw��u�,�ʼ1s ���~���R�@-�H�����&-.�}��;�vۛ��o����L��[���>����7|-99L�":��q��������U.1�*��(���m:�i���b,�y�uԏV~>��|=j|� �f&�fI��Q��:C�:�����U�5,�$�i��J�}��[p��Y;z�얀YH@��@Ϳl)���cU6�*��Ʊ��q�Dj� lʥ�U�M��4)��*�S�HK8"�P��E��(�>Zz��Jp�H�qc1�V���c�rR�p�0�w��Zמ��O7޼z���˓��;���s��EK	��+�ȁ��^D�'�s���i���Q�"��ba�=��t\�!�}�s����X.�JX>�g�{��4��)~ّW�v�tMfm�c�xMr�Cod=)f��RTF�w�W�=���k��tt\�0��F��,�!�S!�3<�r���H�r�N����e؝Iƌ���Y[�U�Z�gf��@���<͍���tV+h�OЧ��	��tߨ���Q���������Ik�u�/�l��2Q�ed���.
�ot+��bn)$�tT֓��gm8�f�`�;�c�OV�|�0"ڷ���q:�|����i�}�|��۲jR�%qP�
�i�n˦m�2��+��n��<�W��˻��OzoMK�Lґ���c�,�x���w;�'i�@kg�6L�x��r�� ʛ4�P�(k�l����?��Lz�e�,�m�fi���r[6l6�
.s��� ��&:��X��tn�b��;{q��I��%��ѱn8v�n1`p�&O�3�mʡ;
���bdF�V1L�e�u1hR0mu��&��v��r"�y)�BPie�!�M�Sr#tɲ�U[j�����h̟U�v՛׿�ķy&��/X������8k8qV�{�y-��J��i��˖J+�U�b�n�����jG�Z�|Z��X�n`���� �r��_A:���~�����*oEjtݘ�������qn�3�T�y�^ O� �!�=��b�gkkwr`��]l�=�s���Ҵ`�
�T����{
M[�ݙql{iN���ta��,�z���β4N�5�M8���>[�ff�a{$�D���Cõ�w:��	8��9k��Ԕ�6�:������¨�7%���^�j��F��Ǚ�̦�"`E����|��mggUub���0���e�����(�) �C4�|�J�Hha0{i<�DlxR8ܞ$E8�z��@���*�#��Y��`ݝ�1n)�KE�9��h�j<`���Dfy�T��������B�d��.�jd�9�9�"to
������f���j�l�CH��Ǝ��Z�!>hί<�Bf,��T�"SY�rHR��3~n��
�D7�1~���Q\7���!C4s��j��OFt�f/V�Ɋ��RW/c
�{2d�|��1�O�y�*�2��O4&�r����2���V�[Z>R�Gy]W��<�+���`�3>Mp-g�lQ��(���ĵݡ3�=[L���@��C�W��I�Q�|w�aQ���R9�)���i�"S>3���Fh4m;U���p`��f?}�c\��v���Aҁ��g�D��^�g=�=o&��!��}��� �V�$Z^��ӻ[*������P8i�"��2-�_'Weձ�率;���Y(�,v�i5� >�f���o>�ޭ��x$�����Ch|S
�����]G�~̓��(^��E܂05�a�� �Ww�&_9�6m<�#F/�&������]���
iL!#���V\㑻`����& �K�����I�Sy�5�����Y|��� ��sn���e	�0q�U_�I�T]����L��>���!���ދ}��J��h�"86��ʎ9vË�cX��c:�J�1���w�h��oIo����}��R���qF+:�E���?�O옪�!=MqѰi��]� b�}�LZ<�����ɞ�ߟˍ�k���|�o�%x\C�(w��WG:�Rc
\%�Tr�%ύB�\��_ 
��z�:��r�e9ЌK\n�"�gbod��{��7i�׹V�f�=�������Ѯm:g���1��۳^7�2)�xԃ]:� �`��<2�oq1��&K�6l\�e���} M.�����^l<�ŕr��q�.o��m�u���'�-e* �ZTa�����3�͟��n�[ݻ��*�L��-�s{&�qI8��scUm��̃�oo�輸[S��
�iv�����b� ��i��!�/P����5�������.nr�ӚX>���e��F�^�^M{x-��ԳJ���SV�U#���M	EeFs���~�Hq��8�1mӉ:��HoEnM�3�J��,��%&oh�]����2���P�����a[�C�D�ݍ�ڂc�ʞw��v��f��{X��;��4̮��	���V��Uصh�v�����K����c9�g�}�	ʾ��@Y��{��kB��/%."0���ps�o:�>���Y��V��iXA���,��'�Z��
w&�Qfj��^������96N��t���9t�+vew-ڻ���˙f���D���(e�Į��;|:�rҩJ�����ǯ0gN�;���)K����o�UbS�2�Hv��.��R��jt��=�E��V��J+ �Y�e�#�B/�V�ϳ�����9��4U�i�2�*
�,�\�uq���Yt�
���uZ��N�E��P�w��֯b�E]�R��7w�Ks��{2�q��[v-���dPg���zs����宸��&�r�֬�݊�ś]Z�o]�_=7%_F��{��,�	�k+ƧF��$��$u{mwv)�r�������Q��oo��M΀���_��]�}{��	)u�2�Onbg��OCZ�A>{�R�Yl)6L~���=�>X�s�{P��$i�tl�F�;f�x�բ�NU���7������mC�&�߫&_ۺ(=��F%�bB�z��Rc,A�����@۔9������2mk=���v�ԓ����OZ�����E���?|�e��!��#�#H�g��;��f�C���s��y�Y�]=�Z�VXZHW�x���#WTn˸�h���9�И��)R���	�(�`yGל�j��7R�I�T-QΎ��1fЈ�jg��}"�n����R���'�N�W��OA���js�Ʋ���L����Q;e�4q{��խ�(���J&&oAel���Q�u�p,�;��3�ڢ��kBM�t�?vuK7G�kG�bf"�M�bCn�N�ׯ��"�MO
d<<)�l�Ώ�sP,fy(�݉���o�ۻ�Z�ԭ���xn�+����(=��{@#։ջ��7���7jk�{պV��M8(�F����՘��E��;������o�c+,#�N��N�{����r����Z���;F�E[I��h<�Sscp���	���E�ʀ����Q�*�*�i0�m�rY�"���Fk4Q�x��]�G,�i�U�T^�үW���P.d��s ��T��S}^����A��3UJL��M��5�$qN%gf��H[r��Ƨw���,�ŉfXO���ŝ��v��NtR���.+o7c��,��wӾ�9[���8ۭg��=���9"�b����=�Nvz9}���N���7b���~�=�u~/��=�Gq!��e�\�oίZ������賐��<�R׉��;쵮�7	�vz"bf`���%6�_�y����Y�fMe\�~-H���@nU٬�ϳ�jz��O//�4'���f� �5&
��J�1�W���=M�uy�j��"��[F�wq�C7��-�vP��E�&����=T�?����ݰs�e<���� �Ⱦ���i�����ɷPNUk҇��e죬$�ؼ��{��~�|%����vҹZ�����I%�����8�y�VsWݗΕ��c�95���r�,��&�-ו{���O�,浭Q/V[Q�S��6^��r.z�no�UpC��YCs���U�b��s`��2{H�W����w�h]��.���F����D�ꊤi�RA�d�{�֖l�'������F�x�g�j��i1�~�J����
��I�5��^v)S^:�9����z���Ih�'0[[a�L��A���:������7.�je�BS�������`�t��7\d*��q�Wcak���Ǩ2�\�+�
�KWE�H�2M����+�=��<|;��A�81���t �jEהu�W�y<�ӹ���޸,���8���֚�Bmp]K�����V��$�7mJp��com�u��3ٞ�ƻ��f��A�`���|�clu4 W���1��l�����׷n���u�i.n��,�z#�<W��W�d zz���Pi���~� ���f�9��)E�̘>��8��M��T;��o7]�Ѻ����o���'��uж%:��u��WZ���>����{%	枑yޯRE,# � ��T��fik=ެ~j�܅�N�)�K_��d��������"�[���b���)���%v���-Y�^N
��k������-a�*�-��s[o<MG��=��m� W��>�W^]��o�. N�M�Gs�|�@Ac��S4�HFO���5�~ԉ_��ӹʝ�+B��uj�ܲ�Hp�5�1�6I���SQ���,H�:�@7M5�RD����Q7�N�H:V0l���m���2�0֩�8#fz���C�m��Yy30��y�5��GS�G^w�*��8,ѻ�a�,N��ْ5��CxI)�&�h�<�ʘ<��I�pћ،	��0c%�U�ՏRz����,�*ic5[nL�qZh��4��.�;�n����$�Xh�UD��;b�jX��=ǗiA�ɞ��;�0dʂ�/6%	~�B"��-�>t���P�-XS�C�Οb��Sy�DO]A�쵈3�n�6��m�=�Q�)b�-�[y�ٙ��f���G�� fE;�:�1�nٕ�C�pm��P�(�.8�i�m���g��38�r����a������i]�+����4��Dվ��Ok��Aa �/��T��0C29t�U1b��b*�*N���xu��@_� 5/����y�/��x?ܽ���������_|��y�W��Z>���M"���$�kh��QEsx#�γ����m6���m����FV���X���*f�E&)=3A�l��c���3�1�_��J׮p=�ͣ�g��8��샘�{�zjSU��gn�,|�M!��`Q�fQ�^r�t.���%���Q3B�}����`8�3sFy���Cl��8b����.�O<1n�����>Z���^)���U���L�୕����2�[D	��[6GqbH���Ͼ3���t9:Y�ֺXVb.<ҕ�,M��ﳼ���[=��;hĥ*b���η3b�J��Lv�&�6��I���CzTsҀ2�����&��Ќ=��~�M�]��=<?T����ysA�������qE>�.�S?J֟�ڰqh-��`HyB&��q����ݭԥ�oO5��9�,�]mi�U��R�G�@Ù�Px��{6��]�}�Õ�m�����eί�^fOn�/G
�b�۹s�9�x�/w�j]MS2�L)Lu�'�T���v���� :j`E�[L�N׍y��pvW'KUbbBL�ȽӦ[ۺ\�삏3+Ҋ��طWQ�Z_n��%�Ί��L�C߉~�_{��0yQ�5`�F���e�d�M>��D���5ͯ�ˉ�X�Jq�=�;���k�ˍu��w	`�J��]�yHyYu�5��j��Wxy]!X,^���G���~��3޳T�����,/%�����~�G|���i,�
��Ǯ/��>�]�<��+1e�č��u&����y�i�u&�|���&����x*�q�J�q�z-��5�R���������t�N5Po��y�q��\��cp��+��4�B~tQ6�Ka Pi�)(w����7_�q�^�Gs��<�_�{KKΗֳ֫dG6f�S3�����h�zƄ���o�32G�:�GWTK�"o���r���5�`���rzk��|�o_`��y��].�_�oi���+��v>^�U����s&Ԥ�J;���<��X��߻����/�5̯�d�M�2�����gY�Ag�s�V���>��nL���,�Kd7[��;-;\i�3|�]�k#΢�aD���Bj<$���к�Ą�c!��,Y��ק�KB�2D�V��������MV�#���Ojl�7�7�4}��n��KJ��c�I�i�a��/�܎�/�_V̰髇�,�c�\c��}�w�wD\VcA�ע���.�33D���{Y�{�D���;GG;]��*\�]��
�V�,������g~�&�!���V���
6�� iq���Y������=}�j��M{�	�:��~�`+=_z.�#{�>��Rj�ċ��È�'�du�TvV+��ʲ�DVI��;�Ħ-��?�ϟ��q�I�v����|m�@�c,q��wfR��V*Z7Q�ґCq�WB��
anZ�L�z�ڣ��Q�� ����[Ӓ=g��荞��G�Z}ƅkz&��a����Ol��h}z�4h��t�F��_~|�lL�>.��|���X���ݱ��T.���hx+�>�:O&.`�۔���'
^
�%��%�,��i�nBB�r
��1��ܶ2C%Vش�E���:�+(��7`�r.0��6f�;U����k	�b)(���n��c�kF��mӈ�X�(�0��aL�[k�Ȣl?��Y�Qb��"�	�)(f��r�2o��/��U�%�Q�|9�i%�9���[>��d�o�j�*��[EQ�����_�ꟺ{�`�vwٟw�q5���i�?s|�e�� ���%6,�G)!Ȏ���ۙ�ŐǓ9׎u�9z�N��T��,�w����(Ԇȗj5L�n��x����4��L��M&�	8���B���]p�k �7��^k�pa�N��t�����h��s�����7E�|&�Ӓ��� ��A㮖�+�ɻ6՛t�2��?����:�WBق��clj3
&v�~['�0_-��\��@�H�K1\Mf� ���mJ<���0!�Sk��e�ѧ��7��#��A�2f]af��� �P�#d��h6�`Ú�.3�;X��Pv��K�lͨ;8���㆗hl��4�M:�+���=�Vͣ�`u͘9yJ�N�=�.��'=�qykGgc�
��<���7kI^����m���Ԝ�b�֬c43_У�5Y����-���HL��&�>h���o�� >�b�sHRi�r�����/t�5S�w�p}�ט�r6��L[T�1|� �5l�'M�����gAAû'[VweQm� joX�=�����M�.1�L�Z~3�"�F^�xKvS���2�C�z�W��9���o}��.�]�_x�\h�&{�^DZ�H�Ek��k+��L��s�m�-��Zk1�(|L ���Y2����З���[V7^\��yQs��.��,�=>������s)�9��\�;�-zЋ0���m����h��2�J�������5���*����~���>��I��1L�v���<�L5K�!����'\�NK	',�
ٛ�4p�l횊�n��W���YDlt�%ۮ9P��Z��i��n���w��2i��S���%�����(��OJ)`���Ó=^�k];��u\c��������A)b��c`�ͽ��)��ƻs�\��-[�����_������Te����ZS0�	nX���p�6�D!�˼2��P�:=���m6CARjk��Kz��4����T��q<2�樤r�!�9��}ɥ5���^3|��J�s�nIm�,�>Fa���a���3����顗;����eZ�z�Hy��,{s���E�g�s`�&n�7�ݪ5�s;�9h�����Ԯ}�xE��+(i��Q.*�Yf���/my�jk�ʸv�/cХ�����~��!w�����T�"�ua�f�![�X�ԭ�HݎR}�n���[n]�spn��K�fc�����T8������ћ�������U,;��H�F�2����c������쇳8��e����P�j:m0����& �a���=v�Q�v8�=ܟm��S�����(�!�31����@
�!k�.��_�\�������b`�dkY���I,z�R�z�"/X�]W�G��Uo:ڠf�WaK70�,�Y+p*�N�$�oE-�ǁn�<k��f��.t��gCVl���Mlt.�V6�Cd����t���n�{��A�"� ��"���锢�V�e�{'z�ޜ���/�znwLS垎=6�K=<��a����}�����2��y�`�˺.�&,�ϐo�7�3�$i�E�m���o4��ٺ��W=�����Ӎ��Q\�8E�o=�rʯOm���Όbn;�&eS�΃�d�b�I�MS�ȳ$9��זS��cp�k��
�z��g���H��Uݛ� cg�f,�b�٠�w,�.�]�HZ-w�wy�,FѦpjÙ��[y:�EҮK�ycWb�����ݴ��6C�K0W�;u������݆9�=��IN�łE]Ӭ�1�;4|+�t�t��f���oN�ґg�Ϡ��t@Y�$�ӻt+�}{��F5e����p�<������c�r2�x�ab�����Ͼ��\tnZ�?R� ����5_�#Օ*���=��9%���
�\S'�JOM��`����&���l�]0ׇ�ad3��Yuo�a��M��ckw>����T��̙����Y$]����p�O]s�-��RkQ�`�88'`��Gɖ�t"
7L��th����y*�O��ʚ�h{C�ｪ��׭��K&�@����
-�9�;؜����l1+:u@�n nNoS�X�<��mA�K8�Z>�.g��^���20ch��=��f���t��qs$9}�~W${��I� �ܾ2.1b��l2'T� Ʉ�5H-C^���lyNk1�˴�Ƿ�J�u����`o]=��}("0�y�]#�[9�Զ]d��e<
fq�3l��1�}�»���!�:j08�[�r$>���%3P���]�Y�B����|��Z׷���g$w�`��Ce,����D�^��޸�1ʅԉ���T�p�י���"��4Yi�j���1],d(Y�m�~Z-���Y�[{��V�2R�)<�{���-����8T�]tD핂�#`�&�N:VLj?���1���;��o�sK����Vv(��Q�S��0��ʇ��C����Bz/Hȧ�/�Q	��c�"��12�}�9V����5%ƴ�f*���&Y�D�u�46m���L'��ػ����1��sSM�%#$�A��Cut�]m�j�K�Z��ٶ�R8[�7��j#]l]�,��a;���Z������j��9}ܪY^d.}9 �ѳJY2�C3��K:�"&gD�i��p�9xE̋����~sL���\���Gȩ)��Ț�F��Le�6�0�B�ҋ�=}�	���X{���bQS}B��}>�2fM�jsOn�y�f�\Қc����0w��W����5���i+�*�{�+�ߙ +v�y*�3n��=�J�`�D��R<�4��l�0DD����ε�MLtǲZ�+#�-�i���?K���j�V��AR�}΍OE�3\������V��d���&�a$ }h�֭�M���'���v����+@�h1�ts��Y����{��Q+��;����g1T�I�mNE_d�殝zy]ʔ����@�=��i���{�9��_f��l'+�)�����T�f潍�/<����
G�A�tK���v�10"/1��|I�י ۠�QH�s���R�6�׺����Pv;O(�!:���:��x��7�ܥ��U��3z���f��&�:cb�ذw�u�]I��t�n��1�=r'�X� ���Yk&�U�:�>��e���wYnTK��t�0�i`�YD�5�W��u��6�l����z�ฯ��۟�s������M]��2v�D�J�ں麙�4xq{�w]��xnNx�U�y��۶��������L�_m<��S���A�b5Jd���}�ٓ%���r��u�rs�EU�!oaG46D�Dr��Y��پb|l�f;�o__�;L7/�͜+Oziy�]���'o�;AC{����LmW}��Y�\���C�`�3iݤ�R묜�ZN��uk�����3�6Q��b�K�U�ٰ���f�����6:+���r��0�Ǣo �7_n�;$C(���G��m%i���d���a��n��3d�V����&_�3l��=o�unr���_��a���aJ��:赥m�'M?�^�k��vܽ�J��bUs	���O˅�12��۷�n1�9`���	��"��m�:�pw%�4�p�33��CAY$�5�����a��C3o!o*���s�>����t��=yvc��j�¶��Ȳ�p���'J����A��l�� ����O?�T�)�"��Ǖ2t�����m鬫�h�h�,)�rS;(�nI�.`"Dc폤m��dQi�ѷ�y��]i�r��B7hz%�rA�`�����k��K��vN�慪]ti�.f������	�����=lD=/O[���xf�_p�q�\��m�a)1K5�ۈ�]6(����ss�����'v�غ�Ѓ%�[k�+v^�נ1�e�X�z�"����QͶǠ�u� v���Su?k�m`n�iHMP,��([����(k�c����j����JXEɜ3Yx�Z�	�iN������ߝf=*��ؗޔ1ޖ�h�Hv���6��A`.-��m�t����4�B��8"v{M�^U�M15�"�1+Mi��֨t�\{]�}"m��mǊ<�f��mWC�CFk �b�q�)��\<�b�z)z��~.žpU��B�0���ڰ��7����R��Vkޱ��yn��u�>��v�����8��y�, � �ŵ7%��(ڦ�3$uؠ��u��2n�t�$�u����f����.��7v�GZ�h!;��h"�6� �l39�Uڕ+K�k�hT�b7 �)�C��K������z%<�:�[��9b:�;M��������f�K�S�q��&��f���7��{]r+�����!�1��Ϗ|"�Rkm�(�i\���#B�X�dFmiՍ��]u�PI�X���d>_3	�c�c��2Y'-n�O%!�s-�����[tH;훖��v�f킈c�3��a� �/��y7/;�;��[]Seť�4�>��`s�R]��B�ЖX�2�6��%�6� �P�6R1J�)R�O��8��W3:Z]\6��nl
�-��5n�'�4�'�2P�S;{t��Ƀh�����c��7<ۦp�`���]�L�r�q,̺m�]}��=���۹�߫��}CY�z��61q�{��Cb�z�v�.��.����C>Ն8��M��(�	���,����Mp�6�t�Lc/\���j]�дv�iue!6�gj*��jy�c������8��2�p
���Q� �8��l!hYi�\F=�����6+��c��=��Ⱥyc!��:��]p�$�Q�F��N,��\���=v0n�����cS&+�J!��4n]B:�v�Fk�D�8nغ��%&`��F%�i���	11��i�-VX������{@��vأ/[,շ��w6�Y��&���d�,��� 4��m�B�Dٶlw��f�j��S �B]aK�
��]J +��nd��z�#������o���Wd*��Q
='y=� �
�;���8&�KJ�a����Ɗ���蘫n-��Br���WZ�����a�����'BU(k�=���j�i��U#1��k�P=cl<�Y�-�M)���=nd�x����14<��G)�
�zUq5Lܵ8[[�Q���-{���b�3����!Vcz�""\?wU������z>��՚�ה1�L�yŭ�܇�
���ƜF�b�:g���8���K@�h����E�r�j\Pn����ºWifi�Ι�"���)�~�1��sK�_�������G�|��ɕͮ�r�3��GЍ���o��5;㙍4VS�Н�Tr��-��3�r�Y��?Z��-v2~�y�{����	���6&�w��k���ΟF��R'
(���6�m![�e<�����.�1�cf?l�����J��ڮN�{9���)��\ܮr��:u�r�F�V=s!Pq���3�Ys�ˬ��e硹�ŵW����_g��2M�2�G�n���w��Y�Di��BOZx���g�Ǳy��v�
��צ�B��Y�%�Y� V)_�t`P�:}�7�('�'da(�41>DfF�WP�[8�>7�ӆ�1M&6�v9t�k*r��mt���V���hPn��8���t'v���څ���h}/pⰄ;��B���(�V_]m���'���<��o2��Q���$ʛnu딹��y�&��#e���-�e�\ku�1WL޿3$IpY��$������^�y}�v}C��U����n]o�Qus�<J0Y~��~m>��yP(�>nY9f�zIf��L&�}Z���شR(:��z�J���?��ў���n7�j�A�2��T�(򦊋�'�t5_5ax��Q�و��k�d�5b�B��ݲ,�����-3�i�-Νرg+ŒUx�z�f���"[�GsJ�>�n�}q���qɟK�;��M��{�AN\��/�!B�����N���kh�5�=�r;��%�9���6%�8�FSv�\W��̻�3F`Kt�e��pA��.�d1%��!w��g�y�2�U�{ݪ�I�[�I��T���+��8N�g?&���O?&����y��^�6��c�V�dGd�boj)�]�l��^d<���:�d�Ӻtf�[c�z)���?)��';�}���"���-����*��2��;Kh�Z���-�"YN�1�#�[�"�]4&Qcd�uGb�����S�w@��u�,�~Z&="��]oF���F¼{R:/�OU&v՗�ҕN�Q,�ϑ|{r�S�,�,���J44Z���Bu��]���@EW��%�s4A�:v>�|T/fl\�f��]=#�7"�X�a��i�b��P�:>%)뻫f��ɪ�Vq0��B�~(Y���wT��j�$wS��f�W$g���mjF�8�~�IT}��k�ۭr]��'u`;CѶ���VL�q0��K�&���-ه��E7"�ս|���ܠ��fJ�nv���g�E�C��.���$������TdɁ����#��E �2��ًf]'b��ϔ��" ���h�4�|��_}>��̧n-Y��!\�0��ކ��K�4��i����0�v���(閥�a�˵r+�9�r���������ߛ�����TѠ�e,B�ީU�U|�s���^����j�j���{�[�F$.��*m]��E�V�t�&)��0`�ͽ����i����^RR�5P�s2��"�[�SD�j���!�0����b����iD<C�j5|�dQ7�ܬ���}�cY���e�p�0VZJ]��~�UTN=�UK`eOK�ɧm�1SׄOk4	}��f�oD>�LD�C�Jaop��'�������c����:�\nY`�#W�a>&�u���"��n���:GA���<�L�w���p����.Jy��v'm=�{��=��%��.^Ω��ة:��R2��'N5gpǔﯞ��T��d���X��D%٘M���ٮ�`�cF-�Fʁ'��Z5��[�l8��:)&.�!Rh��<G/a}	F�ՙ̭�#�ȶ��L�c�Q�>�^z�.E���HC�v�J��yۣ�f�b���x������oC�]wy�k;\3͍0�L��脆�^�n�И�`L�l��J�Ge��R:)J�t��V�;��~zia'�ƈ�fOMP}eT��x�����8m��zi�ܻZ)@,Ȣ,IB6QQ3���m߫"�Bx2'�ٶ[���v�<O�����v���y�^U��~��D�zN�b�xY;�{� (ķ��'w�r66��"	<��u��jm��1����]�E�G[(���գt,��Y��鿧�U��y��h��%�ຆy�û}�<:�!MS}�C�vk8��JD�hZa���D�R��{"��##�[���8tK�)'�!���7jn����6�)�84�%t���r��I���T���2�]���@冷��?j]�����}�5�Y�~�rH����^����v�����'Wv}����g-\��imx^T&`�y��ݞeI�Ny�B/2�S�[	M���m�*'+�[�)3$C�#K���S
�#b��CR`�b�����;�Ab�F�ReT6���YEl�ɢ�*�Mn�i�k�[����cj�[}y���]֕W�gT����s�<4��n��2ù�b/v�;\\�"���C=t1-+%�v�ep�3�I�ߓm���`q��%V���hF]��m;Q�{Xa��%���e��>J��v��4z�-�:����
#��I���v;7i��e��Lsu�25�(T��˞>|��Ȕ�k7!;[qj�i��,A���K6�3F<]�)�v�5ܡ�;	�G�����LlkN�7$U�h2�E�r�n���8��nyx�����E�k���c�)>�&f`������vs'�ц�O����]/xu���3bک�/ӑS7�|괞v�\��巚	0}>�t����������{�y9	B�J�<(V���Cy.�תߣz���;��r�jc��ή[�7#.$i��l���|�I�i�Q^ ۴�D�%:��n��ݩ��b����� �9N�O��!Ϥ��`�f�N�,�"f�KK�1n$�v��m�y.�^��Y!)~ڭ�MI�D�q؟bf��%6+qy��k]��!��عw{�;�2�<�NE���xq&�J=(r*���Y��"�9���[I2Ҵ���bs�}{�����܆9���V�M����3����Ä�JI��!:n(��ɫוxz���h�;3��<$��t�B!�g�X�=r&�>��'�R~�-=rK	��Ͻ��ͬ��W�*�Qj�Yd���3e�
]M���Ɨ^�������Cݹ1��ǼO��EBe�5��I�$�l��kEWAu�Y���c�0��HNpPJ�7kg�A&�FL-�3����H2�vI��q�\�����cv,���t���'�S��"!�ӓ(32�Mq�3�ݯ��2��i�t|��
��R鸮�ۦ?f {k����qM��Kͮu���=�k�����۝+�D9���[���{�J��N�e�do=o�e<W)�\�^���c��{/�~�opi�[>n�������>�~�}�p������Ơ�n;Ot]4,�>��YĐ$��R3�Mz�H�|�O%��I�VoRW�ƠV�h�k^�mޡ,M��q	�v��Lv`^;�R�,+u��^��a* �\%P���l�f��Ϋ&7Z�'.Y��م�a�y�0�E�6�֙}3�]#����%��Z���V�~֎��7ɽn�ߏO��
�l�*|��U�M�v�{�uG\��2�
�Cm=��_ft�a������\��^'s��$<��F�&�����e�NkY���Y�1���s�u�_o���e��4� m]u+��!�Jk�nϒ�s.����#.����-����"Q>�5�oﹾx�Y8@,����zP�SDD�%�P�)�+ml�5֍�ц	6%r8��G��{�3�������3ђ�[Q(�֖�G<��
"�
z-Bkuw��O;)��C��z[��f3ae̍#��u��2���xxy���i�v#7�x۞FSK�|�o�Ve�B�!��4�ꒈx���/3���z9Eׂ	�36���㆖�-�:dz)4�zi��<��U�r�fT��ڷZ����R��M;��("MDs:��d�K�*�l	���쥦�^;k���Օ�I�橌��ƕvW�>4���Q�^w�k(J�r�t�%�¡��Q�L�mMf�f��0�@a%3P"=ʺ�'/Ա脰jh�Q�:C�!c\��=<�����Y��&b!�!�ٺ����,$�����Ѡ�ҙᜆ����d�(0X�5��>�9�?\�G���>��|�ی1��C��%GCF�HA�����F��^9��9�r��ܢ�ֆ�)S*���W@���Ge�[���1[��K��]��dL�Ȼ�N��L�2�EDt�g��>̲���MU8\ޘa�Ѫn��	���լU^C���洟2�]�.�|+��{KO|��Mw�.�� BB؏�P�ί���\�'^�]RHǦ�6�\��1C]����{b�N���#���2d&���Ɖ�Q|��>�r�U��9�f������}�䢢��V���I�4`��u~}�ܭ��}��49c�˖����|�l0�$�<h���!�[(�ٟl�����;3��n%�qH�|1�J 6��7/�Q�.�ɾ�n��{���^�q$Z�	�q�Gy�]�0�
;qЮ����É����E�zLl8-fV?^�ǅ#\�׽6��N�gV�fڰ,{pe�[xr:��;fq�ٶ�c/�]��WX{a^έ����S�����_>8i�.�o�������q�Gy%J�ݞ�>���	��P7(��=�oGD쨋\.';�$ɰ��Ϥ�,Z�5���T���6m�Gx��z�%�˚x����GD��(�lÐ���f�v٤rj������lm���j]Gm���J��YW��俥�t��P'��L�r#���C�{��>�]sM�N�
�Q��g�F���-��lVm宼��{[X/�S�N��aB�#!8��k�8�.���W6�%�[Oft�
��@Bכ��Q���E�V������7����U+�q�Q:��N(`2{��i����)��0i'̋��쓣��.&P���z�$���ۿ���EK�IH�g�K�}��5M�f�@�^�yL�wԺ�Y�EW�J��7�5�#����GYO{��j;j���j �W�a֬�F��2F�J�`���{MkaQ�P�ȶ���/XY�,,�XLnX�q���uUεu�!s�;�f��{�W�PPr	��a�n4�U�T���N���</c���a���s�?o�ci��3�&]�l�UN����"7��I��L̡;!M�V�]n�xm|�ޝg+���+�Gl+2�`TU��9E�d���w���V.=��Ex+��ޕw�]�4�{��eY*��:��ffo�p�����Ǉ�A���Ѝ�Ix:��O����:�3�f��E	w0�pm��3!r{��=g����� ���g��͞V�l��&Ic�Q�t�F^�GYt� �A$�Y���|�:{\y^G��<�f��b�.�4��ai\&a� ku� �Ci�q��~��-���n�	F�j%B�w4e�W+��4\�5Yy��;D�N�M`l�;�[���㬕���ۋ6�Ku��*�``-L�	�|zK��3/�Y�+�/�*�k��No7hoD��t��.��窧���^u�G&��g��U�ō`>���mn}\X5Tn�������[v�殺���d�=�1�>�s�ZM=6,��Hѯcr�禔vgEH���%�����<�p��?W�~x��ͬ��$�_{"`(*� �����v"eL��=\d
yR���>�2��ȗ�����Eu�;{�t�J�%+�������\��Ȁ�яJL�UM��	g��$A.Κ��7UZ����:�u��o/o�)�����ⳛ��u{�3��H��S}�-��nm��q��qr9���ǟx�"'�Y��(�-1��5m�O�ko*!�w��f�W����2�����wն�Ƶ��tPw:��Ʀ,��l�S�|şM�';�T��5�[�@��Հ���k��i�ݧ�����/�g��6�~/n��F�bl�Er��*��a\\M���X�I����S�,t��u�&�o0�T0wN�k0�3[CHđ1�=Uj�6�K8T;8	��G�t�ȇe=��Mc���rX����D��d���sk�>�9�����\_{���M����Z����>ڐ�QjFGG��:���oE�qA˶���x@��y.�Z��9��y����Լb=���⒰ ʷtZ��7$�<�|��μ�Q}8�l'˜�����%�`�f�!�We;KW5X]-��[���A��f���=U�+pe���G޹8>	?r�����]7������w�����L�#��|.����e��1	�I}�.��{mָ������Yh���
ZgZN�[�
�����]����v*$���������y�>�(���>2-]/�9��F���~�Ep�h1lP|П��~����Q�>9O�~�SC�u]�&N�	ȗ�uq��Q|��Cd�=�j��Xa�^�0�;�,�[���zhx׏k9���; 䮮%�хݠ��5�@�(�庡e��L�u!H+a������R!��&JBB��~�י�ѭq;�WEB���cқ�����JS�P�Qۂ%{�z�h�O����D3_"ȂSu��ڋ�Cm�"�-�p!�냑JVܔ1.ﶱ�g|gaë{Z��wŃO]��WzP9>�5�u�����WYDk{7WT���_dW������O�fwv�E#�w�������t����v&!BV��ԓ(y;]�&�M�M!�Ҳ'q�m��ݖ'GG��Q��`�aļN�����l�Y//n̔:��Ikr��͇0n�A�,�m�3:��z'#RoYl�)����YV#�^�sWWQ�%IC6,��J��*8w��?n��9�2YN��5���s�ݹ��h?vY�����A{�a<�h�#����5b��&;E>�S" b�47J����;yc��i����󻏮�n�:�!u�	�R,�c���	<����VL/;EN��l]����kO	-��FȢQQ�R�-oV+�i�h����-D�&����&���R����e�D%��\"MÌd�Řf\{V�˫.�L+�r�ֺ�S��iJYL����8Z7�S�
ВEf�xfԽC�~��P��f�:��|�gu���z�8�ޅZr��a7���)L2��R��b���jYg�r����
c��ԃ���Y�z�7l�����}�_wZ�W��*-;+�e ���� [�U�Ȁ�I�7��/ ����%�ڔ�!̨u�Ł���8�;M���N�C�hs�/o�퀎F(��|6�̔��F��htI'�9޽g$��u�eN��[���h�}J�bq���mwU��W��ҫpZ	h+�i�vJ���.��y�KVR6^LO7Z���L�$�rwiզ�Ʒ�[5*[k����R*���wn���>�z�k�%���sw���b�ond����^.��jeͬ��Ż�B��xuټ�sd[9��ːrn=�IGB���v+���w8���F��Iӭ�g&2�`���t�r U�S�P�d���)���~��dn�vȣ9ɠL���&=.���>�E]��� ��̜�Zovw��]�!�2rt�rH�.��+�o�+C�È!�'�	2؝4���a���[�[Т��7*YE�6v��-�;dtL�z.v-�i�?ś��'�t�Ī�/}�X���zvچ|���V�)�h�2�AQ���r��[n4�D�.}�l���m��D��@�l��%6��\�fٶ	�,ˍb&��➕��"�YEF�S!UU���w�K~��i7�z&+�Arc�&lJ�Ez������G_1\'V��v������H���g��ȫ7 �0��A&�����3�d��6(O#�
Ld�DS\�>WG?z.w.�wm��>�r��j�rZ`n�s���;� ��W��"{�G	������/�n�.�x܋HdKr^�	쓂ΚX<u<)/ gnvHjk*�$�v��֯7z���z��/-ǳA�,�d��������.0����n�=���j��k��mn�F9h0�5׮,~��;�����V_��.+�%A����q�����͈se�\&�i��hS��Tc���Jp�!C�!0�^*\���+2[W6��i�Դ�M+l�<7v`�`���O���$�X�����C��,�����nď�P�9Ú��׌�SD�"��3�2}�5����#9�`�fo��Vhx��6M�����5P�y;5I���/�[E6L���p�\xc��{����|ĝ�p�[��$���n��i�}[/�F�uण+  ��1j,l�^"�o0�������G��y��rj��Mf��&܅Uq��Ҳ�+�g�9�{d�lQ��:�\�m2�y���d��
7�Ia7�ޖ��;l	��q晘������yS�5|O�ނ�W�����N#�L����
�|��x����q�۱o�B������s��9�� �xk���������wZ<Y*{�R����0�����*�����U�Mg����W���nۆ�R#�MWG��Ɨ`I��z��Q�X���}��﷬7�P���������v�[},�_���Y�~Q�#��\oj�����kv��m�޶�������$仱�}m-�~C��}��Z�A�]\��k����N`��wȬO,����ctҧ���n�|�H=O�L�<�T���B�"�����[<�I�.��r�]��keM�N��Z����Riv5`mi=�W#��z¸��a���^�Y�+�w�w����1M�i]˼c���\�e��F@RZ�*���:�/=�Rb�9��9�a}t3��ݗk	J¡�B7L�b\���n"�ipE9`�4���;����4-#n���m�fWl�n��7:����P [5�B��X�Q�m�i�J4�8�b��'X^2���.f!0-��d��l�iG�۵<�m"ku%!MMF�H��mu���E��6b�rqj�&f�E0���
֎��d����t`�0ق���	��v��s\+�Ӻ!�2��EM;Yk����q�e�2��Vwuw4��<�F�ݥO���[Ķs��n�t��C��p����~jQ�q��G=�:�f�rm��_w��_&��얕�V��3�+^tNUY����Y�����OV��sY�KP�(ۑ����u���A��M�3�_�më����ɮ%�kB����Q����r�'!���fI���UUD��g�]ANk8�a�8�grN�`us���;�Ό����,Jͨ���!��T�L�GA.��9dYӡ���A��{�;]�S1�^�u�V��*��w���$���wȹs#Y�V���`�	}�>F��f�b�S��"T��d��a���}C(P��	;�N��o�Ar��\Cw]��8Ǩ
r���fs��+9|�j���� ?�O
 ��������M׻S����\Um���Q.a�t�H��m#uݢ#��@2M���'�.��m���=��5�9����jDۄ;	����[ F�N��:����ܾՐ�a�g��t3�3�q����� ��8b�T�4�٢�9��x�XΪ2u��2n�;�o�~�La������i]�T'�֕�ZZ�T��������36����w�9Ͼ�a�|譳�e}��:g�[��9{� 2�,�6WL�yEi���z-)C񇅎��M�W�T����U`N&6}�B���+���.^�-���7T4�1/���	�����3S�a��ٞe�����|�X0�������T[i�t�����[S�a�Nԇ���32�@���C�>0�` �����{MO�e൧S:�u� Ѣ+�oD���w7�WQ����}��TBG +e��re����qq����e�!�w�'�e��7r����	�A��b��ޕ!����oA��^��|�zãw1�0���y>�i_���� X��G�*خ��'�J�ت�+'�.�"�54Rغ��6�E0a������H�A�1�����6�*������uA��#��J\k�\s��9�=�ql,�:�jr$BQ"nB���6���;�4��h%��{�v�o��K�i�O38����Q���T3s"�����biڷ.b��l��d���к���&�m����1	��Xgp��WOˁ�����ְ��(�;��V�bݗa�e��zct�&�E�wgw��T�Xp���mٯ�;3Y�Q���r�!,TV��J=���s��ӈ_{���OvmG����t^{��d���ŋgWׇ��s�>��έe�N�|�f-��Ƕ���C�}�}׃e�-ۗBVe���뷯07��8m��v��̣���@{���ei�A��/ ݸUh٧YD靶g������s����.�ӧgd���9;4Q�./r�%��i�MU�Dl��`d��eGGZ��|�z"e���jx�m�\���X��a-�_�ClgZ�V��gݎڧ��.Ė:Ag)%>sy�u=J:$��ؼ��R�\j����ͩRzE4'�M����|���J멹{��]��i����bo-���������ߛ�����������WzA�t�c���c,�^���B��]n�)3��bi�X���0\���K҄#!�zz��Vl�8�G©����f�S�gZ̸�F�˚\t48E�˽���\8O�Kc*ٺq������z�w�Y�"Q^d�I���(�ߕێ����4���U1���������iڣ�{0w���7��n���p/�5�v�#>�b��ocf��k\k���pnVK 7��oFky��M�r�*�i�Q�$�������u����vjK������,i��RX�{ ��u���ms��*ɋ�����N�"]��tΕ0�\��s�����z:�Ϝj�E�:�T�"b�Kj�1Vm-�;q����F5n���z{�3�v;�Nd�DWS]���]�k�]��*YZ��ε���im$�x��� n��[���|��dMq����5T�����Mf>�q�t��b�xw�M��K�U0�<!f{�����Bm���bs*�3jb����n��c���x�2��ה���62u�6�-��N�<�ީV�M%�N{�'�s�c�h� Zk�k�k	��0	L�m��5�uƄ��g����/'/��DO}�UУ{��T2ƣ��u/|�r�%ߩ䈤��EDB�3��r[��1��l����o+�};2��j�z�2gv'A:F�tE�;�h��~��_tA� ��Q�h�VC�S���J��Vnu�WM�@�Z�Va.����޸��{��&�2鳠��,�LQ�L��f�����?��;�?lȵE���\U9t̟SV�^xw]e;�G��U�;Wث��� �5,�w ʪc.������ķ`��`��u
��d�QM�az��+�!��gY��tM�Kg���؋!ى��^k��ㆼƲ(�O�
x���y���!x�����չTD1�Fs�]1:p�vtbh��)0�
�j��WEO.n��T����L/���K�]֤*V�Er�`�Z^���6^Ť!�>P��a4�	Щ�l����V�Y���c�J��pչ�&����ggo1��z���'bC����WJ�����ܼgn�H�=��*�3���}r����񧓥���D��v�$���g95pv����g�#4ٰ��6hLJc���[����*��n԰��o�=|J�w9R:�4�t�RG;\E��M��}M[�nV��p���66�ދ�/����=����t<�/h�Ζ
ޡv�Zֱ���P9�ϪY^8��t��T�lk��zZ��^4Q�t,�#��h�@���"Oun�5�����Cj�X]C!2��a����^������;]��rt!W�i���\�u���ݫ�ryC�ˋh���x/ٗE0a�ϻ�7sOS����c�G]��Q�Ӽq�-���&�.�E����Y@o_*���e>�L׷�]��s�WHݼ{��s������7��=�7\��Բ��|.���Ϯcx�����s����y�4=r����]�����/z"2��]lo�&�����p��ͽ��>w	�QX�8;��92ݼ�L��lJ��
��&��]�p�5$�i�n��aT���8�;ߪ�jk{�ݮ�{�*v�o3�����웶��S���������?}��:��z�����DdU�������}��=�ww�]Nt�2��%�����V��&l�0�x�#�Q�t+HY�t3�e�V��uf�"�s�d�`�v,����8�0��� {��.�;i�ד�s�U�W;��78aA�l�\��C��"mFQ4
���@d`s��P�
�|~�b��x+c4+���mb��ٗ��r��n6�2��8f(2y��3����n�nn���r?���#B����::����N�������D��U��MN��Z���r�L��t�����9�n�������w?	v�K�+�˹G 8��e��u��'!e`�Ҹ��
k�2���ۯ��T�p�WL�U��\�V
�t}�:�%����J�ԭ�}H+7��6sV��2�l�c�*2t��Gu�I��I������W��q[7JCeb�E�qٯֻfNc�?p�7�$Ag���)X�u�H�QiTЫ�A�������5Tt��������귥�����:ha��un�q�rb���T��-d[�]8�x�M�g�F1�փ˹�d�(b:������)k� �����g��Y޻���X�8�FfeV;�<5��Ӟ��Ι���}�t���<p�%}���g���=8���ód�_���ֹ��HEE7���b�c (���&�ΏV搻b4�B4�#˿���$�@!1ᇗ}����'�^�~����fS�Ȧ����O8�o:�Es��x��9�k��&�M�ӛ�@��d��(��+q݈H��BvI��t&|�nb��FEr��6XgԵ�>�+�[~����vx`�$0�_LKSi{�D�������|ט�y�.w��]��:��J��$G�YE)��T��=8`�녛9/
��� ;��&��ӑ�N���e킌���۠q�Vf۽�-]��F��ӽr����i7�@Zr�ܢ���*�[}�L��7;��q�������z����(��{zV_đ;Yϝx��9����5ͽ(ܾg�סӕ��H�����i�E'�C[����n��,�	W(L�dMON<67kAQ��bGu�Vv:�{gm�s��-F���q����_/A�r�����LP��n��m�5Tt��ea����<���A��Y�3��sY�h�S�"� �����!�Tv=�Dт���1��_<�0�o��J�*���ө4�m��\JG�u�D�%9cr2i�b��G���������i�|�G_��SRz��/��ٹP��dr�8�'�#���]��c2�9oM�w\�³^�3��W��'����ݟ(VB�'+ ;�t�����E�udY�ڱ,6��1<.ל���B\��֢��c˅��z-E�LKL�8��;�Dk[��E��a�c��!E�vw}�J0�"�w�B�}��\����`�c��=|�S�^[��UxCZ�%�;4k]K&cZ�_U���VB7i r�$��<�ļ;D*憻�`�C8�^l+�}\�+5�ɭR��3�&0%W�-sr"rn�4�'+s�?Zi�wݼ�εKZk�<��v��S�5��4�ʻ���1�r�AV�U�O4��ƀ@��:ݨ5���t �fI��'�W���C6��ǟ.�3�+q�`��	I�r���zc��淮w���H�_���&���<�j��T�Y���꽅��/���D��؁����_�{��������o~�ٙ�Y$w=E�9����凞A�<o\p�8n���o\)�v�Μ�u�����=�m�{�q-�;�s��4Ojf�R�`�$	�����Wֵ��*����Te�{Oc*h57w�����h߹gӱv���B���4r��l�(i٬G�Pش-+�i�w�Q�Q15{�q�9	��o>Zz.�a�q�����G�(���y���!��ϻ+�ty[�0"ݓ0{��M����
v'���q�t� N����1\�$�⮷�!�2�m���8У:^���r����T�A������� C�#?B�:��ٯ=�w��Xs��7lL�H���<lпZ�O��RSxy�;��_���V��[�}���5�K{��'I;����GhQT�Ѡ?��O�:2�i�_׉۱:����^���4��S�VR�^�p~�n��;�iw�Q�
��)��r�9�tl����/��F���܎}�n���P��6���Z�-�5rf"���f�j��Y�;oY8l���gmB����t ]0t�7V��ei��m�J��;_X����s���i�$�񋴍<�^U���p�Fj�К�L��q
�
����U��:��2�[�9f���j�]弶�;5g#+��e�3�q�rӨesځ��6�P̙�h7 \�\��4\s�J�X�R�[��Xʳ�҂Kd5k5>��촄%���b�WM7��vD4��ܧZ�uȄ�]]�fh=�$��f��Ʈ�Gs�D�4� �H��Jl�v>2cE��W�oD�2�͎�9��Z2��6�IJ����?�abӮ�B�lSo���db��:����BV�E뼧(l��2n����oa�hܧ��T�m�v��֭V��];_E!u�u��tlgnt,�vS�mY��/���;���I�Pi��˨ܭq_q�sn�Y��:�X]ʹ��s��M�������C �U�Bv�X�m�Òe�I�����v�uK�F���!G��
o�]��-J��f��i2(ão���d쎍4,��*K�%˗�8H8����c+��pX�(b3/qK�2����>YW�Μ�;�e����ͧ�9P\rwb��r|dò�Gc��S�bH�V��[���y�D��h=�n�1�7;�8����.���O�.˧YBݓehȺ�R���;pk��&l&\��K�]ܳ*=��ɽ_cT6t�;&�A[2qS�G�a�WK{���{�@+ c����A�r�
7he��|f�#�F��H��=��]ͮ�:�1m��L�TYT�3]��d��R[vj[\8��3f�h]��4�s���!�n��>|1�ιK���hm.nM�t��븨14ue�l�^2�:U"����9�IvݶK��{z�P�/$��7�d�H�P��SF��N a��K��2�fu����w p��۞x;a��[۴�����w\k�=��rQ�3�؃��4���{D�ʳxz�~�B���jR[c;c�0ۤod`R̫"-�՗D�P����5�b7j7��Mr��9�l�K��C�fM�P�EJ]�vn���ZKs�va���0�]l�c���8��*g���qz��p�0mM3�e���2B;6@�Պ=XYHXv����Z2�\��޲�I{��$æԁB��m�W��B��Z; �ۃO9��mt-�]�6�t6l��D��CL��X�͙��\�����=k��n�ۊ�w駼�	�M�B��k2\q	l4WM���a�Vl	���֡�!�¦%��pMt�e�&�>���ƛ6/lj�V�B�|��<E��R-bF7Z6B�a�p��U��Ŕ2z��T�]�������R�ee�����mÌj�	�K��m�1u���� �߄��ԛp�arP?ۙ�f��f��@���t4\īW,�gY��-��n��H�������HFf��c\�,q�h�&��ۇ'=�ZWAnOd�'��m��q[iF(� K�q�L�l��������g�W�ƷlP��Cp���{5�x#��=��)�E}x���q�c$�1��X=}5��z��Ir�mha��mU4��%�՚��F�%���k���������Y�>���㜤$�nB�&�z�/j�i���1��x�$�F%U5��c�,�SRZhv�9άk��W��cQ�l�@t](��?!=l���8�wW.p��M��3\́��6�&�0#7^�¶bgg��h��@%t�0�k�l�Y[�N�Ol]pv� 8]�b���1qym=�� ��>����-�5֭�S���6���mțYi^����f�Q�v�jh�h��fc��]1��,�W�N�u��@�ee�܂ug��Ƹ���lp�0�V��,�
�R�Ze��G��Di�8+�sĐA�D�����tt�g�z.@?>O�v�4.Өq��G2��[�asip��j���Κ��TM֒���$8���ۇ6M&亮q�v�gp�u�pb�]��]�72�m�l5��LSM
S�US���K���:�_k�6��7S҃=���^@���н����}>��Of7^�AÝ�|`P�J&:�FFj��.���^own�E��ղc3��D�.�5sQ�.��U��GqQ���k�����ݐ��,D�*��{��L��?b[�㘾`4�6�}^��$���ߒ�4�Pmpp�c�u����ֶ[��͡+z5<�6nXMK��ޅ��T��Qk=�Xu���GT!���줐�Nn�[f:�4�Q�*8��t38@�I�3��g�P"�{���(���5�f��>�*N�{f��e�{Mt�1k��thE��8[�ؐ�=��[�n����I;�s�5�ȏ�р.qv�����P�mb��6:�|��[>�y�����-�Lṑ<��SӉ��a��?GD�L�T���L-fO�8�N�ng..�$\�]�6�k=,g�b��PX�R��zH[�n�O��e"!\W�N�>��Gz���s�t�-g<\�J{^:������˨�R��]Pg��g�0)����ғ���)4���a�a�}�I'D)l�T+@�9W�ӯ���{��w=Vϊ�����W楜��h7��5�jF�vv�c����N+d�=(�固�����9,�{�:>�����D���V4KЂc��ߎ�lez�δl�@e��)#���^��I���"��rV�04q����us#7���RwH�;�{��z1!��#�]�]���n���!}��qǧd�wW���f�7��޹�\��������)��&�k�f��֗w�������"IE
J9E��7���雋�p4����bm��qt����&Pw�a�x����ۖ-|>�-`�8؝u��J7j�	�	��ʹ�{ � �	�f�/$��y��� ��Z���떮��mG-Ʃ�R�BA�4���Yy�wѯ��if�����[z ae�"�1�W�]H�ȯ�q�_��蕖�i[)��AWnh��v��Y�,sh�l�b�4=�ͪ���Y���#�6D�ws�%;���u�uq�T��]�����;�·��d�II����q=�Q��̶�i�2+q��9%9(3��Œ�5r�˶��)�q��e62�i�"IƂ��)��P֓#0���sȭ�.+������xo�j�p�O��j��S\�[��E��������)� ��
-"���������m#�q��k����L[K�DF���Z�m������H(��8V�Y�L��3U��1�����`���n�t�T��Yq
�����ƾϨ��{ϻ��a�v�}��g-07��0N32E��dB��c�YG:��xL�>^��4�UD�rf��Ɍm���`Ba&�b�H�]O]���wP猜�눪I�Qu�Sr�_u�5��C�gI3�f.��w[���m������"!:��������Ŗ����1#���2��|��y��Y�t�\�;~�%�0Z��u
�!J(��DV6���,$a�o�q�d1rFR
8�(A�&8*�,*AO^�pi��㷠@���Z�:���&Q!����XU��Ҧl�b_M��'�K�����_�p�s�����>�
��%%�◚���ju����j�T�vQ�e��i[:	�BzW|�֎M���*[ۋ~��^�@���g�C�%_*���l7۩|^���o~�Ժ*��P�ıw��D+�odt�铪��{��H���B:�dF��Ƿc~�N�>�b@3k�ʲ����j8Twqn����^4���x^�FGla��]�0.靼�z��.�����\F'�;����j�f���^��1�qo�D��m[������Y+��PsVڢbdK��]�r���v���3[�2hu����[��Ut�t�Y��ί�mA|qb�T�e�˔��B�6,���o������|�yB-�~nT�	�7GN���d����!j��6�G���Lۣ��(�OH�]$����"#�ha�-Rd���;�f�/�j��xg�����'��w���O�8�8�8f�y������L\tv�:���WF�	*��1Kv8��.�z��[$]��t�.#��۽��\�}p��9k1ᘰ�����\�s_o$N�7���i�~�?��|�H(Joj"݈L�! �!�]�t�ˍgnlٷ}Ƴ0�{3@L��%jN!�q�����[))l�|ݷ���=�:3�a����"��֪�ĥc(~ �B�5�}�5J���錗]���a����!�C٦���F]��9�3p�ӻ�6ȳ��.s��O1B��6����ށ�7-0��;u��jw������8��}_&��Eލ����e�_L&e&�2=$������ ֪|k0��[�� ������{�C��6���Z�r��d+�R۱����NH��(�� 7��vϹ�ߛj":�s�ëc��.�fF���Б�㒛C������+;��,�YeU��pR��6�E*6����m��r׬&�QH%w.��yפ��՗���+{Z-��-Y�E����t��0\� Q��wX�z����Ï3N���v8��$�nI�Ki)��G�Ӳ�bjq�n^�6��w��w��H
٪h#,��q�i��:m@�K �F��L�kvĹ�k�@X@�����n��*t4׬n^<q]�=�.3��]&u5�\����γF x�_���v�z�՛T�J:�TƧ��sV.��9IsAf֒Y��\�.,�
��V��E#�{WiIGM�ٿ�z��V����u���`�+u<lit���Mkk4��=_cg�2��a}]5�Jg�s��սS��Tg�\6ws-g��g{��N����w�v���CTI\~��~�'�<�t{xJ�B�SSMg��!D9U�nB��?la�V?����v�^�=t�C�w���2}�����`�;�^�Qdf+p���V��Ǌ[3NK��w��/���K��䩅����c��/�*{�*��.nZ���[���)a������Ja^����p�v��e�������E"����A�t�Bێg�g)�<?s��s���	�.�}�>hv��5ߒ�g4.��|M^Q���+E�����{�
u��p�n�aĽ��;�vo����F9����v\�0���vU7T�mU�ރ2��j������\��c�g��kG\9���\��t�<���ZT�X*���n[œAY�<æc��O!v�:��u���ImbXO}�h���s�w�w��h�"Y1���cz0(�;��5�Bc'\^��v�Ι����,��<��3P�6e��Ӿ����2`S����ΕmYi؊�Q��ބ���6�lZ[5
Lp�`EG��TNW�ۨ���mۡJf�[P)q���\��Nƀ�P��4+�E�����T�w�E�szE�w߲�W���<L�i�`{}������Z�s��a���Y[��k�7r��٦�`���%���ډD���S�<�w��k��!d��\\NC��y��I�5�|6E�B6r5�k�3��l&��	Zc�NO�����:���ɭh�L_'`7hdˇ9g��4i����h[Uuwq�}���*c!ݻ�n&�!�EC(=��0��.�ͱ͡��O:�]�Wdj��w6��h���G[n;?�p��8п�}�w�v�����w��UR�u^���W7��x{��W�@����Ur�L��EuUM����ʃ��֥s�y�[�������FM.�Q�]Ż��ڠb6T�5����q�EE��hB��EmQ�48�y���L���fo/>�3Q��R=�S;+w�*ǖ��a6��䦝�A;��w�̑F�A3��߾nGa�o����������eGY[^wv�5�e�m��]�4§ʛk��̧�������Z>�� �[��vԦ���/�A�� �]���BUM����&�-ߟ&�L�#���d��7��MP��R[��T��>��̆�U��u6�+/2�TӼ�p��̦o�-��OL�ȵ�e�+e>�Zv�fe�� ��<Ȉϩ^_��Xu�~�����ƭBl-U9sDC��H��蜴�-�T)�s�y�Y��a�~��oz�g�۽NV��I}�ӡ�V�����gb#ן�X��(
��w�i,����q���ܜ�ᗝ�뉹d�vT렝,�V�oh��n����ޖ�����HU��3�jU[���P,���̞:^�f��D��z6��T5_7���[U;�V�\y���sojP
�MJ*q,�y�/gh<Q�VF77�;�<�p=�Pm����TpR���>+�w���I�_�8��{���ρ��'{<���~K�'5������o�f��KT:�n�Ң��Z���	��Oٍ[���0�/w�*:������>�o��4]�)wyW�d�U�]�6�3�<�}�ziޠp��ů0GM��)���w��}K�L�`^�i��o�]���o�fq��������ho�*M[�p������+`�r(�}�)l!�/L)n��� R@���fN��;Խ:g�G5��/%���WGR�E�;b�^�޵�=����_Ә�[�=���d,�H�ծ
z����R�;ǔ
�K�N��fQf�6�;�J�f�!u��=�;%5���nu���0���R��d :u���Bg�9Iwiؗ��S��6n�mF�;��G�뙼J�]��:���zP:Yҫ�}=sWsQrC���:b�=|�eq����;(�n֓�M@d$�oG9VOg~�q<����Q��K���)���àk�**F�S-���YsD1��P�}���4�����\��1S촳O%T��1�VSG[0*ۜ�:΋��d�5Lg!����F��d�@#{��=�5��<�c/m��xю��� }��k!S{�*���w�~����9FQv�w8.�ܺUX)�o/#ɛ�W4\<׉~�f�����Z�[�Ȍ�OP���N�;3�*F�y�N�,��7�n��^^��>�z�]��#(�%����v'�M}��_�AbZ{'S�}��6w����ї�a����ɋq�Q�����+8[��w"���-E��l��SyE���.��'�Co#>�T�i�%����ZT%�W��V�f�'R�Q�}ܪ��Nm�j�|���Ȭ��zs�������Gs�"Kk�{}��ֶv��K:.���͜v�@������DA��G��z��_t��8�������ǂ����}K@�4��T�wM��63��������R=ėP��N��D�Ql��M���)�������k��MZ��}����
iVwl8��H�������N���6����:3�ݗ����|3�y�m�6%��hր�&;YtжL�Vms%�ˠ���!��Qy���]u�6���c t�u���k��M ��+	�ͯb����2u�z;Qs��C�&���/7N��؉?����]�����SЫ��.��h:�U��<i��"͡e�R�!��Y�o���?�Ͼ��?ϯ�͗����}�5����=�y�����x�M�FA��Gl�6������[wr���9﻽z�V0��R����P��:���a+w5���G���]��VL���n��E��({|��p��*/g���t�;9��sz���p��`�	:�>O��!��
��W,��	�~�Lu��Xp��M}u������N[���� ;�(����<��`���gH�cn�
h�諔wt�O�q����]�i[Y�7�6����t�����{�)��^D��&X4╔��	Y��
^���ѽEƏOw��4����jN*�RuF��=�[�FU�RѲ��)g@��c��"7���h�Ĳ�u��	����q�h-�b�З��[�����Ff�[X���e�m�l"�R��
���+�1Н��b0߿��������Sܗ�ƻq���[��v��F;Q���U=��^/��k{71��D�8��۾�ܙqU��egC5a.')�;�r]
ML��O�K���}>	TW��ܬ��S�K~5�l4B�U,�w�͙��{��K��U��(5��N�V���K� �E��	�n�U��%�e�5ۥtK����*v�Wdڇ�]�ݎ��!��͊���t,�ngt&�0������;��{!�F� �	]�i��b�ZP�fJJn�)w3�ȩ�W��k��f ��Mt�Ʀ�3v`��|b$��Z�S�Ҭ�iZ<ՑeC��"�����F��n���������K](��� U��CmIT�v)�ۼ��\�(��D��WUV�pӜ;u>@���c�I�}��erV��l	Nms�91�r�o݃"M��;�HFXS�i�si���拐���w�,�n�r]���V�iq�`s+�0�g\�}6]�d�����J��<���#�MDh	�PmaJ�@2�G?G�#?JYE�|�̴�7�!h��J|8�'�ƕI���/7oa��m�����,���L
��^�P+�'���Ü��i�<��ڟɖ����=���r���)!^����`1��V��H;�����<;>�������^��Cjm0�;#VK�'���y̪g"���s��Yj�J�R������}������p竴&
�\?tȍ��o �Kq0�=�<��3�J��P�l.yw�v�Ӵ��j��I�w/����iųjd��v'	d���?+Ź���`���=3�.u*g4l��G��5�a�Qoa��dlMו��]Vro�b۫i����ۭ�瘻O�S��/��Ƶ[v��s)�lg-���G�/ ������n�Z.��}W��,u/ٝ�-������霐\�Ʈ����8�Q���M:cv]ڗeu\���4f��i���.ŋO����<U)|�[��8^���j%t�8rJn+��u��q���KT��N��\mX��0u�N�Z4�r�Lxŀ��z�<7�qt8m�
�D^�Q�d��~l�eևT�d�����T�Mj�����7[�L�F�3Vތ�j�j�"�ծAJmi��$�}{wb����e퀶m˫&��V��?���o<�:��1��(Nò��3���Ԯ��#�B�mYWڹ�.��y9�/7�(Ru�?m�;o0�}\�qw-�WϞ���T��]b̾EW,�m�İ��y�t.w���
U{wicڍ9*�{D�����^%�ӕ��i���α��-z�[l�{��Q�ɼ��c�v+�ۼU9�]��e���*��kgm�z�����������wnK�[�Xs�͇v�j6������r�[�7�_L���[��7�*Cx�ĦU����kA��c	��F򙓏"N�X7Y�j�}����tO7:ro��������V�I�g,K����{p.�&�m���=����ly��>�/ܣ�Nf���r��_�,�o*��J%܆D�L��v6���3n�:�:�8�Zܑ�1�1���P�AB�F�`_L�t'P,�Lz*npd�<4h�'%�k�ULV�S�f�pX9d
dK�d�Q��N�bjk;�g���1e��j��W�߳;s@�6N�JqA�UX�r-�fC��M&�#o\"r�7b�Z]��Q��,�fp�]�>g�*w]�V����9�W��vpk��\�Ic�?�y��Y-�e��>�{)ə�����E[	N�f��h.�)K ��,�V��S{�@�iMV��kr�$�I�1������}�ɰM��4�ڝ ��
W�R���s��Q�jb���^1���i���o^�DK>�3�wB"��� T\D��T�ۅ��n{�׸�
����M4��ZlwW="�T�ȍ�{���].����&Y�v�VW+����z*#%c�*��-ג��UYP�Z�0MB�N���8���U��oz�Nw:H���w>߮��ט��f��ʶ��^+�ӳ��کw�����@��q��J�'M�Q,�T[���)D{W�4��yɬW[�N*ɚE�#�R$K;�򯫞u�Z�8]e�-X��'k�wX܇lh-���l�,��V��9��s��o�����%Z��#b.t45?� ��Ȏ|���ّ=���oκ�J�{<�}K��_��1��:��}~�^��/�7(��q4�ƫv&�6��Z㵙 <��LR�[�����4��D儰m{���Y��_p�g�w�ۇ�}�L�;�꧲��aADu*�ܦmx���9߹'�����#�'-��H]��.����"�
�$�����k�}�h�G�(Q�>�����v����E��3[C�cff4����]�6�ت��������].�T�){S�g8,)�@�d��t/Z�<:#]4r���!���ɕ<Al<Aا�F+Ζ�SRv[�&�[���ʠ3B�vn���Dhyg׋L�IrۆMk��On����"+���s��_O\L�I�K�7m��+t���ή�uq,g�5�f�qQ��+ks��Okz���|i�|j�ݲ��G�o�Lɢ��Mw�&�e�������3�O�heA�eN�P���s��]���|jdH��+�31S��<���0��<*+i��{�-�1A"ֿd���c4S��s{3�ċ1V4V�m����8�80����Ms��\��c,��w%$-���8�pl*���1h��_g��ʤ1�]�ٝ��j��1��fo6ƹ4���=��p�G����.�6lp�����#��Q#.,77T�i`9��ٱy��7�>��V~��J�,��c���vYlL�f��*�-�@Գq���`�kq��˕s�����Q��^��q	
q�Q������My��m�ѕ��vk��*̘�n^� Ǳ�b��c֋l]��<�`&�n��A��I���;Bh,�理kM_4���UV�R���&M�4)��*tq��]�:����I�)�n]���[�7�?{=?X�Q��-�q��Og�<n�U'c�Pm~�t�4)z��/ �O�w��XL�r��Sx�z9�d��f��n�ץ��������X.u�2�A�:�x�6u�d58�ʸ��`m7��+�F�ÿeݐ�U5Qk�p�m9�j��w�x�-���2�l�{s�N���0�m�p��T��^?^{Y���O�T{�j�ň��f�z�k������$þ��� �c=?v�Y�����
�u�2�<9�ՅZ]�}/J8�%%U�P�!��v�����]����΄�2C�}"�62�u�wC���@隽�݃5]4�)��'�����a��*{�l(7W�LF�Bx-Ӊz`w����M�c�&��;o����lِ�&X8��� �mr�J��?�����:����)�W�[��6FT�s��b����0�������=��͚�����a^O:�6���nm�3pGd�^�Kի�-�9j;^+�l��M����r���s(�2y�7ѻ���y��[��Z��r�{u��/'Jyr^�U���M�7���c��\�S����]���Q�')��~_�;�gҐs���F�7�| ���� ���4{����u\
ʨ���pŝ;0rSMGI��o=fb˼�fŃ�j��͵|�Ĵ;�6k��܈���--��ܧ��׶���=�����YZ ��C�/Vy)[�i_��i��u�	䲻���w��c[7�����֪����c'
]z��F��p�Zsw��5�1g��.�h$�e����ݗ�ў�9���5r�|��βB.w��g���M�&�+���켦��:A���V��R�k��S�ɀ���iͫ+��J�����������X�ѴR�0l��sk���<0K�e���eX�OL�/y%zc^2����B�E��#�\�Wv'D)SQ�}�9SD[�Mu�;��B�:�T.�Ӆ�SD�w茱������_s����US}'��f���
ّ��(!���Е�UXK����Y��:�Q��u)��v"�,֗A�y9�6��Wz���5�p�m�����yu�߇����%}̿.s��3W0iy��5��{��ǵ�˞�m��{׷8�t�6���nS	����n]J��a����e|��a�+"�,�Ńn��cV~g��bN�x�_�>��ļ���27r�{`h�}�ƫ3���(���[qk������������7f�wvX�I������C+#1L��y��*O�tF��џ}���qVtZ#��gӣ����:�o#r��)�\7�)W]F$���r'��S�\���Y���z���c��X�Cf��B�c*�cR���(�&!ͻn��B���w��,	�Rf1�r[@-�,�h�t�-�P����rz�/0 �+-n�hډі^�}�j�/s��nc��O(Ș��i0�L�C��{�#f�����M鮢(��ӕ������S����7z,Bd�7��J�Q�k�d3L���`3]q]�&N�&s�6V�L}k�:d����ޥcO�������/YQ��y(�N<������33	�:[	��e�[\����dԨ����bb���u�x���oWW������##i݇;��up3���LuN=�XF�͠%˘uw�����b��v�ۢ+g��q8jͮ�ȉ�;8G�*f{�l2}��V���)�BK�Nf�d:�䌮K9&'v��d��X\��������ڨ��Y�	ZB�E��;�$��r�a]�rϫ�٤c����UW�ݘ��D��Ȼ�d��{<aC�K��<�,1��1�Or���{�8�b��[�cY��]�m�u5�4���fDla��u�;<���������u	�Y�v���+l(E*r��+%G�9A�=�<��gu<�S��Ý��T�tZ�=;�"���}��Lؼ��z��M���tޚ��!��빒|�V R�Q[��5Γ����i�|u%U�t������{C~�f}�'.��o��ԟ>���E�~�f�?H2�/
vv%�j��^
P����gt��)I�S�5�{:��9�v�����~�웡V�S'��i(�ݿӏ��O	>{Wr��V���76�`~��<�����ʚ�����独C�+�SR�l��2�^���2���ˮ�i�L!N[&Z�4Qf2٬��s3��k��Ɖ�c0��w�����,�Rz�*�f �M;��y�����I���3��/0�zl�T\���fK�m#�N:L|�+�F<�؝�|�g����N��#�5�o����N�븧ח�9��5�Ev ��g7�E�kuEN��T�����ԯ�~|�O�	Z���Vߒ����m��mu����kn��=n9���>s�;�v'<�2�v��ie���6��}�%��U�DK[{d�`�B.kH�ŀ�5'�B�܏A�'�pC'a�ÛJOv��C��2�qm��w��I|��[�Ri����zݧ�0p7I8M�0OB��5�{v�tk�<u�*5ݪu@O=�*F8�wqx:�u�ۇ)�(�c4�[�g'Q��4q�,s�� �)�&L˸r'\�aݢ<���:����?�v>Q�/�?�x��Njt��G��cr�a,���VefWQ�a-M�� -s)^��9u:^��^q���)��߻Ƞ�A�-g�[��є�]�jOk�م5vn�����Ә�����X��4�E[����m0]*��"1���m6�t����/j�
&���՜�����:�`��g������J�����f�C��Eu���0�%��!�#�9���M����g�jpT+)]�:ȗ��&"��FA��ܜ�����!�k��L���G��ߩ��T��Y�0b�='^nk/�>^�GЌ�w�r�ժĪ����+� ���5E���=���BO��Ό��Vx���=N�V�oK���|r���2y�ST�Q�!����ݱ��ϯf�Bڱb;:�B���ٌ*@ᦚ2��&�7'b4�Ɩz�f��g7�5�^��~��Wr�C�V����3�P�b#g����j�"ٔ��^��u�M��P��3j`�)͈��?;�	G/�KW���P���6�޽�Nk��T���4�Y�>ḿԃ>M�B��ckVb�[���#��P�^Cg\�'.}3qV_b6D&��ƨ���E&Ʃ�sU���ӵ�a�nC��s��׉��l��S[g�|�����L}��ժ6��U�w��dG�u��&�����0G^j�g��vy�ͭ�%;f��Fq˰2���&N��|�/��fX�wM{_��Ta(�*<�,��eB��L�N{#��Gj�we�f�r�~R+���V�P�]�#�uˉF�pf�eu�w��[���t
��{N|�}���A�F���Z�u����B�[�+:�����CBV�Ɣ�;�O_U�Qyݔ��
�щ��}\�u���nf����~���������?�ɢ�p;¥
��8G�v��=t�O]���3���\[MpR�	�W,�ϒt��c�DodS��MU9���5ތ�xѮX���j��:tc�Q82�x�w���H(h�ǭ��<�͖)"�u��#)�n96c|����ҽ����~�{��g��� $)��}?<��7S�O��v��r�A�os{�[_k�n���Ak�q�ƫ�uf֫k/���9N�v*�(5v;�l�DD�V!�Z�\�s��NÃ�wd��ׇS�P��z�[]J���J���Q�Fژ�I�Qu4-W�>�=iD��{xx��̚�[�Zg�SMq�{}/�W.��>�]o�G%��7�_�a���~er�t_u��WmъbLƼ����݄7Z&�����Z��\ �ڋcf���#���X�NY�ǌ0'B��prY�g@2L�i?=�x������\��gk��2}�ov��'�P�Ңje֌ĚoA��g��r%�wL�N�m�8�:��W���E�cr�X*Å�׊�!Z�MhV;s�«��A3��|,ݏN�MU�[%ݷ�R����d�)G6�G\�U��@�f؎��|��խ�VG�ߣZ��T�-g�O15U�gy+纸囔�mqy�{}������~��V�M���/�aO�w���9��m�\�]7��<=�����4�l�,Y��]æ%+wP��:�v2.Ŀ�A�g\��1�9�&��Z�i�|�+3&1�F�pɏD
�����->�V���5>�至^������5J��jeO����,[��O�.[��O��}+|Z��r����׵�.�t��~�*�_W�eɎ�abE�ݴ��{Q��fS��rL���b^�(G`'�2k��
99�J�����s�[]��-}x�B��e[�f.�l�_/��>�i*ڿ�J�c׷���Ș��-��5��ky��dB�'����1�<�"�E��f�ÞO�Q�K|˷�LQ�u��P]"���u�#".����v݁w1QL�6m7d���mb�^�M��^+�T(�kQ�'w(�d
I��ɽ�a��%Ut�nƘ�뀠���S�3��m/4�6�������E����d��/�����]�v�ght�n����M�ɦ�&hA�M�΁;m׵�¸�fV��ڞ�ɫ0��=� }n�T��l�������g>����>��Y�|��ڴQ�R��v���ĵ{;��&�ݹ�d���|������ʭB��;�k��Pfc"ZC\���hV��C�-9��+��y�魪����=O���Xm�|�p�Wȍ��;�m����Υ,�������j��usE��HcC]�7���%�Nໄ��$֦V (��]v��NM	����Fq&�����P�W	;ƽ�eA���'�]<t�1&�5J3¬�l��J�)4�~�b��Ӳe�@ۢ:g\��:��s�iۼδ^ne����v]=�˼�U�e̥yZ�de����|���ղ����w���ҭ9ɋjT�'����E�V7����]uZ;W��Q���U���-	]ֱ[�ml[|�/�ʶ���
�"�[�6�l/�<�n�u	���|��Y'.G�k	�ʚ�,�ύ]�b9ݚ��ԗ�3^	|*ٍ��[�w:�d���\k�l���ه&��|�ҕ��Ӥ��g��qǷ�&i��Y}��4�骊�ҩ��rO�5�QD���^���JY��33_U��']WW3T.1W��5�Bw6 �;�mn�$^G��_H�N�����@^�S7)�r!��L����6o\*��x'�3���
���Pʿ�bV1�X����X�Փycα��{�w:C] C7W6n*��s�V��}��T%1`�E�p����VL*�R�خ�� �qJ�7��˚B�l�jh�M]7;�8���Q=֠��:z�wji;{�oz`q�!v^�U���s;2¶��l�h��V�J�Ěf<��P��Q��P[I�ݒ�MZS����j�����~,���mi��̬�c�����iv�'U��ch�ʈ�����Y�|���D�p�����U��;K�;u�r\��P���S�����H6�:����N�mo�8��`�
ΙM��v�Cx��JoV�f�ȵf���w~u�����e���G�n��'��J�)5�P�K�UWeZT�����N��Gm�ڒE�t˫�����1�f����M U�<���lP)r���qE�XTڼ��WY�A2�qŘ�/f˚g,rVl�����0��0G�]���9 .lƽ�2�饨�E��k��0Ea�)�P�MW���V0� �ҁ�j'�d��V܎�L'c�[Q�6�Tڥa�޴K[fٮ�LJM�sChA,*�+�����|6�Ѓ�D�7�ki��m'RPq��!2\B=q��m�%4,6�l�:m] ��9�;31���ge�v�q�� �#]�N	�GK��͊:�S��g�X�;Q������(���jDm�k[4�0�8p6�^#D��WlB%�Y��zo�w&�z9LsO:�ޝ=\��b\�t ��������cP��f��ƺX	�[*&��e�9b�{ޡmۀ�)�f��zǯ!�dq)��cs��n��.Wˤ�h�,�0]�0q�]k�k3��tiW���SO���.Ya�]���|(ˤ�X�2�Tt�BV��.�wh����/\G9",��E�������!qkv���|;q��o���ǧ��L���N�8�KD��pW����2�̱?\�R�ZG	+�1� ���W(y�,�P��
����hI6�g��}
�&�c4K��t�����H1C�)zWY�����e
�!��c�s����;������Q{��<Pb�{8�����F�볡��p��L��b��ZxG����!�p�7>3л�e���z�fR�2�L%Fo�����aFkλMu��˥:S�2��%��n���.���F8��}3����p<x�wK�T`��ݘ�w`��u�;��y^���ۆ��a�CL%�Z�K4�(k 坊�� �3�>�󮲑(���R�,L�5a�],ԕ ������C,�OAһ�J	�ع"E�ص�����Y/7]O�F��:��_��J���ԭ�h�[q��J�K��[��h��6�x7Oi�݋��=ɥ�4�K-��2Z� ��Ѳ�]��]i-ͺ��L	UtB��z��[y�����L�0����Y���&E��~�/��˸z��ݳ' t�(R��j�ha����%,*5נ|X�%gtv���^*��A�<��J�Դ��	���e�������[�����&6q�9&]W, �J!E]n���fLW
Տvm��9�J������Mո�ܸ�HMs��Be�u�6�ދc��ߥ���X��U�x�Ob;W�d�vx�eV�=q�3�n� tc]]���
s�~���\ʘFQ���W/J�:4ؿ9wK,����qӴ��B�N�q���ܥ.�ר�f�6|���ª�m*�ڭY���}��u��{4������ɼz�=ѵV[��f�! Y��Z[��3*�,.�;:��7ג=_eO:k��Nk��|��䖻N�l�.�ݽbE'�L�Zxp���]��)ח{\��b��w���c!�r��M�0P1e]�p��;��M�3&��Ay ��H�b��y�Lo6���/��Jg1emBٵ2&�;M�uu��j".���36����଻�C;.�D;��.E�.K� �~�����r�ޞ*���;S��5��Dur�g���B�h�O���T�;�J�'m%��"{��L�I�8da?���;��#�i�Yu���	P	��[n����*P�j9��{��ۇ�����۹{������8�=�	�sGGs�c�ۼ������@/*s�Ow�;1��8b�$�֗�y���v���(~���m}/�̂���7�Q���ۍ���8�����.>)�c뼫\�;���}�ߑ}�ezfw3�+k���3�c���g� �&ۓ��c���c�#gl��Y��4���x��mv;�T��n������Y�sVع��~tr���������ݒ��˵*mY��9e61�]66+7���+z�lK�ҥ�ڼ��y��͏|S�5T�E�;�R+0$�����y�y��,ǣ��Z��Ϳ]�j\��8�Bf���|�ςl��7LF�NR���L��5?n�Uō�8�d�z�e�\��9~�D������e[�D4H�eBNs�4�Bn�=�%�O61��r����(����O'ǫ��n���Ŵ���H@�#�~u�f���vΓD�0]���[p����n{V*���w.�ʌЄ<-Z�g��]7)�vqTʚ��9�m&����ut�Wzg����`��oH�f�J��E��j�n] �`\�B��%�Yh��F��_)�^�_|<+ن.�s9�>�8~K�����aWR7�w�"^�V�a�y�6i�R�O�M�N�ΡU��p��b�y��������ΙY;��0+���-�6Y�U�L��Y����`J�x�Dt�̮�%�s%ZJ�yg��k{��6�$-�,�+9��'s��AP����2�=�"��ntF�lSkA�
,�	���ՙϷ����E�~7շ����Z�1��hw͉�ϙ#bGd��T���P�;��B�{�:�{�l�t\
�,��K ��ò���B�|ވ>I�wI�`s��:���+~�:	u�Dr�����b<ж촠V����Y6E2Ӵ%�)�%oVe���Цv�d�D�����}���[����էL.D㙑�ݎ��Túg7��v8�yއ7n:j����4$p��t��JN��S�}-���.N���L����gT��l;]�]�HSH��OI�}n�y��'@;/r�s�霓G��#���+�ku������x�
V���"hWݒ�l�W�ܺ�����/4ʇkl�K[�N�ۣw��;�_e><�}Ǆ<�[�I�Y��5�
}���x�[+�vn���՜v��𶞧|\�.������p+,���z���mr�\�q��}��ĨK`p����su(�Y[s͌����T���nb�E�LDKI��Ɨ��'�%
�ZҔb�鮳\ڰ� s���rN��f$;��ݴ��������v��6v�?�����~_*R������~�����lc���ٗ���@4zi��m�W"Ȉ���&��&���0|��o˅�������s]�}�*w��gQ�e[Y��(�*fZ:L��4F��7<��Vz6đ�4^�؄�`G�]�x��fL��c��̄����.{�������s���EQ~��z^�H;ɲk�sJ�]Jx�B��R��N��8-T=s흻�u���V���V�ܩ���G�>�Lc�����.���)�r���^;�K���T���
ɘ:�V��Q7a�F2Ե�Y�����d�sq\��6f���vdHu�^�㨨���{5zQ���t�3�����~��ؽ̋s�q.Mf�Ů-{dT��uU�큚:����g�R*U[c(~Ӿ��[Ϥ`�y����[���ҟEW�;^lRzku���d9*�xe���O�{SY�57�Si��U'ߨ P�8�nK���j���<��Jch���УE�M��9|�ڛze	��ݖ�}�����s7�&,onJ�
�J��2�\�%���1{͞��a����ԝv�L�]����q�n�N튼�]f] Z���fo�sN㻖'�K��-�[�5j �λ��m{9\*�n��3�M���;g<����#{s��������=q���.ыh�8���v�&�-�K]6f�e1���.�}=[K�hK-��SJ�^ݣ�b��Sm���HcPQ:]-.��3^{7.��;\m?�����A�m�R'����5�F��zݥ��Z��4p�=��	xֻkm-�`���́lb
9z�I���x� ��V�T)�����`�j? ]�'!N��.��`�Id�L�H������M�zi��J��Tv�!5g{*�Srԃ4F���]�1�v&��J�F�WG3j~Q5Rᙊł�@�U��73���bEe�q<�x�	��L�}Ʉ��IR.��G>�=MC��A����|<O�W��{��g���d��YA���j��]i�����l����;��X��X=�?=i�5	Kf]�l��i��RN"�u�������!�ˎ�N_�ug�<�nS�t�֗5b�S-`���X�}���Y�Q���?J��\"{7Pm�K��M�=6y��� ��nj�����V��9��w�g�#ϻ��K�ߥ]��H_��y����GΘ��&oA�Ϗ��æC0�+��Ah�9�,)6Y�S����7���ˉ���[�&]��.=�8��殞}9M��۷�8�B.:�덄�f�zcg�DK�s]�m�N��:�mu]��m�(T��um$�@7���3���4:6�,���7:�0�#�p]�s�S:t�]�
�ˍ�"�!Q
W(����zg��ء������Wg�׹4L�`�CVzp����3}8��y�6�zݢ��z�V;l�}�c�\�YoP����-�]���d^�y�#hf��:
��y靶ֻ�7�db�R�z�����}y�k�o���k���	6dB�I�����3��O��5�h劭�i4Ϟo��1[*�hq�ZhN3��B]S<\��J,����eK�1�?"�9wtĻ�I�j�b��qwX����� 2��]j�t9��=��od���츹����6L9��~����RD(�o�wgw�t�Z,�H�OҠ�x�>�y����[-��U�oD��9g6���p�Ir����!(�[��d-wz��b&l��)�����P�rc���U�<�`�Ȅ�͙cll;]��
�![��<�:rlz��r�+R�%+B$ ^_5�r��Z�Q��@{f0n|�K��� ��ya}��#Lq�1����ZF�
h�����oi]^��N�}�����t�l1˄����zi�,Y���h��C���w�2 ��Kqu��
U��X�>ˊi������su�[��,Nd�3���1�����zբȭ Q��������Y�{Fo��L`~����%f؏�������	�_* ���s)̷&*7&�ewn��Z��f]��]�ż�3��E1�LN������VR��횺���n����0�A�Q��ɩ��˟wѦ����iC�nY�'i����f��z��#��:��V�C����g:������.�6��-���^��d^c��g}=�܇��:�oD��ɽ��2����v}G��gH#M�����ڏ^[\��g�	�O��R��[.{���߸N�x���>ڐ����厮�X��~�z|���柳<�=����:�F�{�o�*ڷ�fo��r���
73�y�K�j�8�2]c��I0���]F�{+ F�V	��Y�3o�zeO/�8�����#b�̄��N��c�.�j���K���f��+t������%㳓��,p�wf������6�m�"Z�Z�Rv{�ܦp���)�MtUl�M��Ǧ��n�̒Nv�j�|:C�1i����|�y�xv\#��i�g��P�]��w!�����Z��]��r+�+]Q*eF/��̒�|w��䫳�s콞xvz�G���-c�dk����~v/}$�ᖡ�Q���S���ڦ�����=>�q���6��UO�
:_�Օ^���p���܄h�?�i�Ѷ�'`U��6��(�4����A�u�d���zBUf����5��t,�3P�g]r�
��͕Z�
Ɲ^����I	6�������6te_�i�a�!��;��xT3��w#|�L^dNK�Ñv2^z��S��g�<��3�oH����u���܏_5ڔ����>{�+��f,4ы�[.m�uT12l�]\�Ɛ��LQ���BGB�BY[�q�f�"���ZY��VgeR��2�U~��uz�y�ܵK�^a�C2�y-���1<���	ͪ�ڌj2��_2<��r��E��\��BSt���t;��5�&F�%�si�˦�\ռ������x�d�a��=�xكش��[N�g������U�ett@:�
,������j�l�Lfzgq=AdfP����6����v�Ig����C�O������NU�A�쭆�뵟���RE;�DB�&��#�:��WS��E�FQlv|:��S�ĝ*�i�
�}��Jx�㽞y꼍�WT���S;sìr���L읊d��ث��J]���5��k�zZ������v���"tMJK��LSZ�*�*����5႙�(���\GR��;���i�5}[-���3S���~�� .�c5;z�8M�e-\��b�=LWF��|b�����{��B�����~�
���t���ݦ5�n�B�y���
��N.�dc�JA�%���T��u�v ;I��u���w]$�,���n��ۀx�kp�A�4H4u�jL��Ŀ���=��v�-�3b�y8�ѯ6/~_/��\��3`��Yl	eQ��Ĭ`��S\`k���۪r��z��������Q�|!�s��� Uڊj)cW`hٖ`����L�9b��hU�p��!��mm�����V�q����Tt#p?�⛿`���^l
��4篓D�;U0[La��UE4��<�OMD�>a}�~��5��m�-,��ҋ7�e�/j�<��L�C3��U����K�9z��o�J�d��SG���?Oq����۩)�譼oG�+BHΖ�Bx��
�1����Q�o��)oCi}��e�y����� ��~�Hy��^��������$�»`Qo�?M��6��Si���s�ux��_o�C:��]v~z��m�kVt_��V}�&2�����ߚP���'w��(P��� ��4)���7�*f���(×{��ޫ�oٝ��/�HC�� �b���-0�L��N�ʴ�!�D��k�s�ʾ�6@����ITE?A]�ݳpF���{��b��s�sۧwe � E��)
��O��KW-x�]۴�Ո�*������^r	�v�c�O��p���>�u�VJQJ�,�i�]>����l�gݕ�q��q��?\	�����\M�ie/�43y�26�wv���W�q.��7�'Z�;F��m���:t�?��{��ǡ�}��g�E�.r�*e�냔Y�:�V���6�`�DEֻ��>���x�  � ����4n��y �]��c�v��΁�����\��������{���o���>���U	0N2�ִ�jY�i/�h[�f���e��bf
�n�y�e��QYɼNf�Խ�߷u#������_�������?^�?~��7���݋���������?�����}2����-�ĭ�ì��燤پ��u��@?{��˩Ϯe�:��776��9~dQN���ϱ��6  �8z���tĈcq�g����:j��T�0V�C	=���=��쭅�0'�i<r�`kzr�8�=:q��`�H|htౘ{�%��aT�ū�3*>���C*��[w"v����{���)Gk�v�К)u�r�
�vq3{��K���ɰ2�~�QWι^��d��3��1^�V	�옔�'N��d�L(eA�nBfo �B�\ً�7zx	�"{�9�Co�-e�Ӑ��({�8Ph)�_��U�4O��rJ�0Te��L�f�2��v���zM�p滗��ZMT�~"�.C1�:Bz�xo���
ȥ����Wm�G����ܭP�M ��RH��]jv�/[�f��� �xnu�Yw.�$؏;+���Wyb�8�#qԫ�v[�Э�\�Zݻt;8p�<�]�b�u����y��F�,��8���ퟘ�0^Vf���ޙ���Ƈ���tɛN�y��/�w *�T�����,@�V�
=n-�i^M��p����Y2���82�s�Icw�������j>��/��Y��1�Y��d̼5���ܵ���a�a��@�7z0�T��J�C��f۽�ܜ'.��H�r���Ӡ�<� �BR�@�\u��(��`�.�r0�4,���X��:�w!b�U�g	;ɬ��JQ{ۛO^H��6��`&��\�8	8��l�\Z��Lk�Qq]p��hv�pB��{��u�l��j�3�S�T+\�C��q[��'{ ���y��-�s��Ş�Nϩ.��Zf(+_�U�5oO��Y�viXy�k��w5��+��ո���L���ǝ���:�ɼҍ#��u+�_L4y	�e�%�l����m1�] /�m��Mf!u%�����*���t���ջZ�����jS�w��o.m:�U�w���iU��s��+�A5�xwc�
܇?�ފ�y�[[����_	�Bzt���I;�IW[���=2!$��E�f:�z0N�u�q�y}������d���"k�^���(|��[�)���ٝ���î;47[=��؞Ic���߰�؜Ӱ��魦3]�%�~�K���\�׿G.��=�e␯}2���r����I���zi;�3<�.�%�꽩x�`K�6MM�'�٫�У��~������z�J騗Ҵ���~o߯����_G��g�9�a흞h=\�����,��#\W��-#Dr2ku�cj�Pt�+�� {���ա��K�S\.R�vn��1WUsE����in��ަ�g�ݦ�A��B3J�N�Zj$��N�΋�:�9��k�T�X黪��=Z�+��=��g���t��#g��f�]��12���r��cz#�k/)ƻ������o�<���$#$���ص�c��CF�ry���{S&��Y��9CY��^�h���Y�r��B�=R/b��q}_�{�[�;��7���b$��{�[�_G'��a;��gE�:��-�;	\E�ٱ37��v��p�ZaKl�!0KH�9��ي�Ÿ�c�f�0����<vob[t���N�:;l�7K�m7��-�ݷ� gT�@|
�����s��~�����c#�(/��j����W����w3��3���~��W��w����<>�?d`�V��]�)��PS;�#��60M��%��.	`Z���4��lA�j�����gZ��HF��r�����dc�B����/�x}q��>k�np+�:X�r�v�S�e��p��b��2�ʋ3M���ʸ��h&g���䒣��,޾5��3i�?� =�9V��ޞ�_�{�:hz���#�۟2��+��Z�)��7`�{Vo����3_jW�aUD��[���g_����,���2���:s����z�4�I��׻¸9�7�i�u�����)>��]'�u��5�@,��,%r�i�Ji;��{���L/�W�0�ﱺ>zt=+
"��OL�ە��Ӭ�m�z���iќ]�׽H������g[M��S��Q�E�e�;*��̈́������Tp$/nL�Eh�M�:,E)Vё.:��đ�C��٢�eu%E������39=��;:ڈ�x�w�=[[W���w��%���p��C�IWm�^:���qݷ��Ϗ�_�S$��pypG���zmM�˳�ԗR�aj@�#k�U#�X�&B�Li��!�1o<����t�A���vLY�6[ű-rK�� �5.Ц��ǘ%��lq��
��7?����8��m�Mc@��!�zYt�icb��jC�ȧ.���`���W1���r�M�p�}!Ll	�9f�#�nJ�2��D���(�f6�bkE�����J;icΛ&�	�B쨹����m��.�ڻ<W\��۠�R��f����}�?��?�$�y�3��~����,���F(��=�p��� G��q�ٞ_S�x}AA����kj���M2�;k��f*����T����1[���dv���}�^P�6+�p&�����;�q���n`�w�)�|)�'gg	��� �L#1�>K�o�J����[�*�]���t��^���y:��@Ǻ��E��׵�!��?1ˁ3E�"�Һ��ʔ��M�!����٤!�/%ɓA�g��gv\�t��Z�<�ہ���1�w�o
W9�N[�e�p�P���5��}+��wmLA"t�^w�~�-�Yw�[c�{��&*J��7X+Yw�3Ң]�ӯ�1*J�\�"�᝷���66�U`݃]��+jV���I��r��$��8!%yʼ�����HP+�����?��D�S�4I�C.e�K�]Y۴�lDs��Ϥu�������)O�����ݚ�8r#�al��KSe�=-h��e�̣h�L�0���b������lX���G�����u�۵yJ���O7\���Gvz�+�⳩̴�f�0Ťexf6�߷���6�B,#/�-��I'�w�)�S��$�L��k^<&[cc"vT�]i�C���d�i��B]sTBc�$D�cn�܎��*��3x�@rj��R���4��hkn�;�~eo������l����k3F���AS��-�S��ѡ��i���7qS�/MLﻱ�T�΂���Nnn��л���zzr���&��W�ɵ1O�Ȗ�gh��oR�3h\4���y8;'a(��ܛ��)�,HO0���:2.zi[9ݎֆ�'fnr�WB�N���{���·s`��N�s��Ƭ��]#OLg	���w"����\]�nJJd�t�hUK����Ͱa�Yp�hD�N���[���*cfMѲ�D�5}��rT�n)���]s_3�w!���=��:G����3��%�o+<��W�T���4��o���bާ�y��03Z��-��[��9aa�4-֪��ͧ)�d�%��ڸo�~�~��qbw���69}�nL]�A��Zw8x;�����D<;{���c�jf�\��%�}��1����G=�� �G �����,���ձ5�o"���΂�(
o|j{�uN���՗3K^�~y��u��c=�~e���a��ex���ڦ���j&az�ݩ|�u�39Mf0��UOM�ĪD)=���;��E������,����,��[v�7�Y$��&�.���]7r��p������o�1�q|6:��\��.�[��N%�B�;���3;x;t����\���8���V*K���ڬ&�R�k��mp	��q��u�
�Ѷ�O�gY"�_bb��yP���=1��K�i�C���v�<�R�jP+j�e3Y�3������w>K�@R
 Ƀ:N�� �Ѭ�ΎO{�Ͷ'��5��)D��F�]z�&�Y�+,�{�n��<�E���n��~�,A���mmko[Z���Pu;.��sgk�xw£]��0�[��Zt�w��fڂ�hh���ް�q�����餡��j���&4��Z;-LT���^�OLz���m�L�
�\�l�P`��X���*|͑�[���}����֖��%�/݃��<(�ye��ћB�(�{����4�\yhŚr,������ц��a�M���qK�4�\`��C��]����{wj!I)���,Noy�G>�oeba��yu.e�ߴC5�_M&���u��nn���M�oG%�)����ϻ�Qe�$C!QT��P��"�D��e+�NYEI�
o�i	1�m�QV:��ЎJ:A��!�l�w�[vL�WE4pG*�x"(�m.�Pr�q͠�����镕�w��Ÿ]��}r{�ث�D��ء(�.E�r���Բv���c<��Ƽ��=��	-��`���r�7_�C�42E[�w�;$���1vd��sk0P����Fb�b<\�%���ͼ�?n��?c��h�}��V�><M>��s~��6h̯O&��6��"~�#Ru�h��K,�t(�A�8ꫡSyW�$2b�E�\�k��)嫔e�1~{�s��� �y�{���]#r�k(���8�{������;��o��1ѕ
6Ê�A�2�K���\�Ӽ���/��j�~�)����5�D�A�q�hJ���F9/B�����xd�(�P�c)\Y�-ot�Z3��H��s{��K��ᣰY\
#�6   ;������N���$[7M����ƒ8ŉD��=0��Y�}|B�@�0�S4�m�L����7;|p�;�&^�s�L*d���4�G[/�k�?}`>��)m-М��\��R�=>�k5Ёn����I���bP��L��e�s���2�e��-���Ť���vڍ�{�ڷ�s\g���Zu�R�D���3tA�-��3�]�5 j��Z�7������v��:Lqx����Z�����ln�d��E���\��a��<�Z��鲢#�[ͦ_!��K���^Dl��if�3�����J.]���."B�;YII�{���_{o������SE��z*�}+>�P�}��p�sK�u.��eF��Տ9M-U��wyJ��-���q�k}�d��؜/0o>�}�4Ż�Fۉ��kOw�zN{�Oسۻ��{���Ʒ}���~A(P�NY-�s��4��_���m�c���<�C;���ͤ�:{���Q����GP�|�2Z6��N�W{�w(Z��[�} ��8�wL��ky�r�jm�ոim�Ւ�p,]:�L�[���E{7������~ٿ�R���%̢�{>��V[�X�t&�%uB݊Ō��b�����1�bn��\qk�ǉo�����Lsm/�;�í@��������]k��]��9�}���:�l���E�F}���z^IL�H�,곻c��GE�K��#j���is{���9������"�n�Qb5,P�v������n��I��S�(���#��������oR*��{��	��!SNb]N*���݀ �<�C�׏ٴ�6���s(����Gξ���jw�����#c#*e$܏)ч���Y����[�ޛ&����즋k�P��,v�f��J$A����)|Ȅ�pf�v�99|o�\[�Y._\�(����;�:~|lm�||�Ko*�s>B��Vo�j���DS*j���Y��b��khֲ{s�/����ǰ%g0鉨�Zeuo,%���I[û���Ϲ~����Wۻ�5��$�������HV��n����p�qۋt�c3)��lM�Enֺ�K30H��t��NM*�;n6��̛'v����2B��Y��-͚6Ʃ3�o���B������8!�Ӈ�N賳3�W�yu��OsTZ'�SC��/�q�&��%��Ae߀�DY��,h��Ψ����Y�ky�K�Nғ»X���_i��<ɹwI�Ԅ�fW�}��4�m���9	���R|�9^�u��P�j�)�}�n�,�i72!]��8��Հ��%e(\�o'�Ժ�u3�(7�!/� ��l�@��w�ɼ͋��窱GQ�P9�x��n5Ȭ3-���&^�݉cn����WNs���fsK�rvw�u�D�fH�K%O��T��ݦ��R��F3/��u�x�:5��;O�YbF��y��9|xЪ������M��krA�)�vnV�A��V�79�h�j#r�k�C�m�B��ccNb����^���^�<Ng�q�b�t���wճYzJwR�fw眽j���ț��d״SX��3M���H��C?Y�x��%wލ�������]z8N�/�5#��x��L��n���ew��C*���e�*5E��\Es#՞���U���s�ek�~pyj�ٴ�^)���6C�A`�ق�{/ڥh�]:�ӧ�>�7�f��ND�勠e���Crz�����M����{�u�U��=�o�J#*ti�,�+N�<}.�ɋd��n���!�Z��`r�-U�D�9�-�\͔F^9$C�{\����[�,��B�C;��x���9)�z�J~�x�8�ӝky��,�μ��������-�n+h-����lc��Q�;��׫��������MZ9�/Ge���Ɩ�����jbǘ��sW����ؖhLu�>>��S�ϐ�(V���s֙��D�e�~�x�=���̶�۳Ѧ��{�A��b�˾'��6�;��x>��o�5N���������m��R���_�������Ș�u05��7o3o��=���`瘳 Y�p�5�l�U{W��fP^֨�ܖm{ޞ-eE�Y${����
~l~ +��z�Ly<8��ch
�d�{���3zڕc����Л�z�N���i�ˁp�j�fs�m�0�J?�a���e�Z_
�hHuxk��gl�:yk��5�l��OGYP�ĨA������O��������%c��[
�L[��Bv��yP���T ��T ��t�����5�x��{f�r���P
0��A+�N~��M޼%B����7�*k���P���A��(A��p�P�������^<<����*t�T �=>���>��.�n6~^5p���2�u��j��ߏ"�kM0T ۯ_��d�Mf"����;f�A@��̟\��g��PQْ�J�
�U"P�)5�m��"�Rle\�Q�R���E$�J�����
u����hA*�kgi����������
���@���TP�T��T�(U)@)QR�EPH�)I*�P�
T�PP��A*�钠	R��� R�m�)N}����i!�ws�v<�J�������7t�L���n���[o{zO6���t਽��S�֕�9�*\ꪉ}�։�׼{+Q��p�mJ�U��{r��K���>�m�ؗ�)*����[Oy�{U´w��6�[�36̯{}`/���U)����kz޼٪�g�:��$�'w�)����̔���")UT"	U�B�A��^����s�o}�Ҋ=N����K�FZ�� �L�����<w�IQ�@CwwTx� ��g���L�%�*�C��M�tH  ����R�΀�Z��Ώ7nEV6��Ң�T�R�k��h'��TFM�񂆁@Uy�|!
x}}J��;�9<�Ε@e�(���A��@��z��u���޽������EW�fXR�9�S�>�rA}`�9��qG�ݔ]�k \�TU4Զ�Z���$��P$*�wE)/N��z�َ�����b���f-�z�҉���z���{D��w�0�Lwj[� ���w��Gu݊��PUVxu��m�0��]ڊ�RIV�<n�&����4��J�׶�^{�ץ�c�[���w��o�q�cM�l����{�)#�}���[�̘�gJO3J�7y[-f�u��/�zm���U�R����)UQT����IT���S�����{��P{�����(�nx�T���з����ͥ����}�����oT��tP	�=B���94�6�V.��a�j*�a��u�ln���%z�w�B1�	b��4��y�( ���J�ok'z��c6j�z����P�u�]:���ye�{���^��n�1�U$ ��q�P����
���D=׶my�����BV��{ިi�V�]2�-}�|����z��W��E�;��q����=��Շ��zJB;�
.zzU�����f��еһb��H���^�����پ���{�%�Q3��UE>��Nۦ�o8��:=����{�T��ӧ�=�qKf�=�k��תU>���"��}}=��}��|���OG_y��w���p�ڷ׻��v�1�s��zR�T�!2�H�2 )�0�JT   5OdѤ�S(���H�   ?�Ri�J   z@��T�M0��~����~����y_���^�W��pn��8����P�>�|��G�| }�πY���������P�!~�	BIDD	BIDD�IBIDD�D$�DB�?w��?����2�Ҽ(�N0+�Aˡ�@�J�j�2vL��.�m90i���N�8-����{M�ueJd���	�[�X/Z�V��|�FX#�W��\�Ƚ�� �biy61Թ�\@+����PO蔪�N^���"�f\G��툩�a&�^��#@c�a��v@�[j�
�IkR9[�%��D��[� �ѐ@�1f6"R�bҮ�*U&5z�qT�^��sV���%��6iBV��[�������p�Ņ�bd��4�n�Z���ۡU"0�{�Z5�%#/�lԣ�Z�w��.���1�&�D
�&�� �E�X�* ��S���m�)�
�/k6�&�.<�C53#y�I��"V�:h�R��ǲ�+M��<ߕ���FKW��Ɉ�Lj�+d�v�-xe��w%��6���UZe.���J�@㻀n�V�%��-X����,ۍd�FR4f�j^�Kp��cV�U1��f��V	���{FU�Ղ�׶����E�i�4�P�FL���w�k��)���-�i�,��3��u��Gn�$.���1�[�iY.�4V[ D)^P�i%0�PVl�,+1�uX�R���ӎP
�6�dy�� ,��-d���B������[��х��9T&�kre\��R'w^�
��F7oI�{���Mn�S�A�9J��>jS�,Lڃ ����	F��`���^l�ֻ]��)�Ұ�TM=�Xɍ�srX $&�@0�,�x��c+�1mK�!�3J�<ub�֪e�2ݔ�y��*K��heB�ȡc77B����ّ-{�vAR��0��6��u$I��BA%���3b���W ��v���n��jb�.�`0���T��wc8�uTtV`��+��i`���b�&�ʚ�el��D�Z�.[�Gi0ret�s0�U ���F� [�h�:�;2�R`�7��FΉp:H���e�<Д���@*�
ɕ%;�ӌ��:�[ c��n-W��UM�"�,�G�D���UC�w-�7
&��bJH@��������0�w��kl�)�q�cwpTJ��,[�#Jr�JZ�.���n�uh�c0U��l�ٓB534�uM��5���P����^ǈe��o�4]6�[�G;B=�Pދi	s(!��<�����*CZ��:�⛙HkՁ�E�B��H�5Z�N@7..
(��R�@�6`4��i#[�*�]��.:*ѭ��b��D��lC�Z�*�e�;�4�Y�k��V�˅��˧6�+n˸VpA��%.�Z��z�d;�������F$��=*��TN�ix���P��F�n[���l����E�%�	���7'R��̫���S��lfʰ�H6m<�j�@Tґ:P���tn��"9��J��f�M�na(�$�Ls��jk&+4낮)�
T��jR�m<�^d0]������!�\�Ϛi��:cw {Xr͋ĴR��p�3V���t�Z�g��Z�T�aB�9a�7��t�/r���)S�4��0U�o.R���S��u��F�m�lS�X�Ef�ј1�6�ϓʇY�J�ޚ�i�ȫE�zr��y$v�Y��2�M+J2��L�t�656��f� r��L��m�����r֓[Ȏd�n�ʊEu1�*��8��{7B�䙸�Z�*��P�Ŕ]0��-Jۤ�+n㧦�]Ɲ^��%�Wh���0¤��U��(8�
4���kN�4��0�*���Į��R(�5��d��B[ؔ�rZ8�N��"j�Xfé��5p��jY1Р�G˸Z�T[�!���SsT�3�O瘢�4U�4��Z'wpdA�*S����R��;J��۽.��կi���@[�/����R��oh�-�Y��[V�қ�5��m�";��hnܱEкr���%��=8S���e,�M�D5EaV-l�Ml����N���z�=i��+�W$�F��vԕ�5-
�z4�j���-�6qn7�5�q �:钕��S�9�X��{X^�j�C��e;��iMԣO	�4Y�ecx`˃�'{	�O�*9�W�=�@�e�@�5H�5��A����Ű�i[X6��1B�"�;)���,�3�˃�j�H�H�I&S��M�91�8�Y�n��6�uy��;3t�aJ.�U��U��',LR��]*k������Rm0#��`L:���8ESю܆��6l�>�X��5�uʺˎ^�������˺H�d-��Ѩ
���76�# ��вZ�^0&)P���2�.n))l��Z��Un`;yR�"r��o5��X��eH��R,f�R��in�`�F��7���C0�(�H4���k�q�ܖ�H�O__�:��m��ۚ�U�ʈ}���>p��5j���ӥPٰm�EuX������3.�yU.$��k�.���S&��d�cǭ���HV�D�p��z2�p�ݸԴ�\TL+%W+Fr�:c%L?J9��
V⽩r�nVn+��$C�V1B5Ԭ�JfH�Uu��)ٵ�P�a���f�a�ҋ)�2�ʱu�v���������ń�xlf�*���2)��z��SvУVp'���[CX�����$��2\��kC��ˎPf�*m��Ƶ����� �;�uPݔaD�D�o�k)�sb��"ٮ�ɰK/�m�XiM�37v-2�`h��e�{6^;k���XB�`��X�jVh��60�[c.�aTBUF	?�w�Q��ڶv�i\E"C�.f�R	�� ����iSɮX��9���W�5�2!HVp�M�)n�s�n3�gD;㽟sܫ"�a��y��"�8vo>�ϵuW�U�s[���(+DWe�E$��gi{� 9C�#I_V�9:<�N�ҹG4×Buw���ޡ������4L_<��)�U'�$�ӈ�#�1+�dBrӧ��	i!]���RE]���Q륩�P�H�����RE�4�ap���fInK�&}�ܔ�EW�<�3�sem�f�B�f�%���j�Aj�=�H�TM�f��Qm`���;�Ze��1@�%����Ht���J�)9�Q�Z3@�2�f��64�5�g6P��9e���Ǐ!$����#YY�%���7)�7���-�x�i3q��5g3�pPs��C��o��S�/�Ƚ�"Xݳ[�ʕ�t�Ж�U��I):is�GER��Ni�T�f��8Wv��ϯ�� rh�Ѣl♟kFd tU��D�0�ři(1�c���)\�FU�nJ�Y�?���{P���5f�Ql��nbíS�p�ko(^:�.���d�!��xD K��w�dR�Q|%w��P�8ȣ�X�e:r�"�t7W��u�p�a:q�i  �`8jКʤ�MZ5���8��eB��B�H��R�u[&��7���hx*�ٟ�����4�q8umT�A�������.�� �f�lTF�,6�KU�G���Zf��򚎡�3FSڹ�^�L��@���0��H�29��ʹu-D�:�)	����5�F+EM{�T�k�Y�U#��䙌�b�V�Ɠ���d�W�J[n�2�T*Ś
2�!U��#�=	��o$Ƿ4)[\�6K%�ɒx�\fnUbc��]i��X��o@�j̖���+�Qv�y���.0�ˁ�-l��%j�CE]=�d����2���
�ȯEȎGӶJ�J� ��ԝ�26��*3N�8��AB���,�tl��蘚�[3c��N�xɥz.Y���
�X5����[3�_��4�Y�hV��]e�zc;L�Z���	�f�.�"�劆Z�,�d�謙z~������ج#�fͥ��E���X�ڙI������)d1c�X�j�k#&�ؤ� �#�V�vvlQ�L%���c4Ll���ٸ�䂮;��:jꮘ5�XƔ��KZ3H#�i�b�;0퇊ѡWm��A/.RP���)e��L;�cϥD6<p��7���4˩v��J��K�V�r�+#V\��N�d��),�u���vV�(T��MY��P����!�7B�J���ַiJ4n�L ����	�W�u�n`����HM���͗h����Y�+!�&eO���=����^�x�����;L7Ef��[r9?��J��cM��w�uc0�.�S�謉`��
������wu.%�e"$z�ѩ���$�[���4�hdl�q*�X��+/)��ә�v9��LɁ�
�T-�Uo#!��)D�b�wa&=D�dJo)ҦK�L9���kw�؆�!�/���M�6�����iyN��i�l�"�P�k\R=��҃*3d	R��I4kF�8������uHƩPzB�F��!7X/7�X�r�B�m,�<��j�h������&5�j[�b��-`����#���5ͫ�o)d�ɦd�u����w>��pY�f���,w���_m����ǂ1Y"Xs]����H� :��{�i�F3oq���.� YjP	�XQ���喝�Z�;uq^�,j�v��E9�AM��T�_���@�!oT�3e��:ٰh�yw�1(�H\���|eJ�6$���%>m�n��k�e�L����;�x#��{!R��5�E��P0��n��v�\�9V���
�������7YsV��hQ�X�(]�7z�ԡ"���y�,���\{��uFtW�RI���D
45n�t�������s+����L X���#a��E�5�7��ݑ���vFd��Z8������#E��1
�!nnCd@����ãV�++��k{m�kNGPKtr\���q�dH)e��X2*KJ�jn�v/�eYr��^-{�Z�nK���.G��7eZ3e�-�-UD�Mp@�SĮ��!Ŧ}��f�:NIb�^�7L�(�����E��&c0��)���fm��f��0��!@úq7x�L �CM��QڙJ��i�=��w�<.��JVpe��� ��X�B9��4J�53
y԰�+���U[��8m3���
v���ʪmI�keE�h� ie�b���9�M�{�Bt�=�$-y��T��1wE�L���[��t0�d8��fG���ƠR�-�t�-"�:�ׯEʫ�א�i��1dױ���t�j[*PڒB!��vr�B��ݷv)�v�1�7TEԸ�ٶ�I\�K]e� �Gnى�r�����F�YٚzZ��+�Ts�%�`J�2���Z�%ԫ2څ,16�O�a,�}j�,�˂U�~27�`#,�QRU��%���JfeXt�%1aN���.EEF�&1���Y2Z���xd0�`�ײ��f�>��t0µ1&Z�cem�{�l�7k�D:�%5�Qf�v���x"ff�ͤ2�U����j�2ƈef��bd^��
�4 ���n�K��;����>�ɫ�RQ �ӈ�յ Ј�;�y7̺L�`�{�)DIp{2GJ����3�Xp
�ZG.��/�щ��5G�t���㧉d�6Y�V��`;.ْ����qQܤ�Vc�`!�m^��FdA���4��O�R�JFd��O	��n1�5�/E՛L��sJ�W��H��D�eݫ�ˉ���M����c0����e�d�D��U�[Wn�Ve�F�pA-Ĳ<�d7V�˓Sz�q�񫘪͝�4
�`��N�G�e\ ��*��x�cZmu�V���(f��׃kok+$�C���i����^��6��B[4�u���A�f��RԜ1l�Tl-ޡ9�Z�U<Up�8�b*̷z[K#�<��]B���M<�1�+�+oT[���i �ͭ�{��t�Q���!�E�S������#���\8GO�(VB�:}�Kq�
��r��I�c�s�[�)��iV�KxV�p�]�K+�=�eXN_(w&
Xz����ֲcz�4��RY3}O��\��Guon�!X�.�I#��w��%�U|/Oʬg;����dd�n'y�a�N U�>02��d3;�Z�9��1rw�w�V��}b�ֲ5j��م���1U�3�M�J�k��I��wE]h��S�s�>뿨í��s%�o�V�c��#�v��.�-̔�vl�;/�V!�%@�aC���y��t�Xi�����YS�x�	m�M��ۯ�,U-��)-҅�u����v:$����2'�K �sl�#&�e�.dt�M�³Do)#���w�
��6�Ap��Ȫ<L۶4ZJT�Y��f��#gn[�jڡ�SF���AUB��͇]f�z�*U�!5�1�4�y�U-K�[��s��xI̺mˑjʊ�݋7+#6f�16�L�:��[Q*uvh�.ՙ���w�\h�
�����NX�QL;�,��b�hP��I6��X�h��i�6��`��DL"lt�7��Ԗ�1Qd�5b%�qY��	>K�R���1��^XE2�Y�l����5�fބ-�2f۹Ve ��v�L0k�l[�1�ź��]�7����7��۰�&�N� �(G��MB�x�@��)�G
If�2VՓ,�M��j���5棦9Zwg4�Ƕib'��Q�cr8��t��ϩaj�^��}0$��ncfCYL?nP�%f�.�ehA�b�l�3i�0�l�Vsap�^˻��w
�'�Mď��*d��^8|q+-���� �'d�;�PRo1�n�ڱ(��ArLV��Xς�.K�H�
3�!� �:	�z��j'�mee�9�|pn;���()	e-n�t��ea���
����c��z��!Q�� �p�i�ysp��f��Fe�Gwn {��f4�L��Ob�l+(����sT3p�ܢ�h�:��/�QI��+��T�r���2lcbηnݢV��U�i)2��;m�UB� @U��UT l;gl���3��)Օ�p�r�j ���]�ʚ��_�����#]��  50*�"��� ��������g[��j��-UuQSe UUUUU v�����l�d 6Wm�UUP*��fݰ.�Η6�A��,�C�*��i����t)�m&-᚜͕ј�lO>_<~X��{��|F�wj��d^��i��g�t60La�c�W�����ܯ9,���^8�.c��X:ml��5LDT���cf#����D�Yib���/VX�Ɩ�M��,�^�E �Ա���5���2�r+�s�����;a��m�-w �Lx��Sh����6�Z�k͕^���y=��`�g���ۜf����M����0[8�'������f8��<Xic0meQ��F�1�8\a��4�5�,��V-XK)kjT�6	���TB��	Gk���':�t�*��厗�5!�w�"f�y9�3�Q�u�E+��\)��Bk��4�sW>K�]��+��4箰���p�h�;RhPgq�5�q��e�j`�(h����H��8�祏����]ϚMJ���	�T�%ic�pr����܉kѝ6��_^ʧ�}��T?'6ǃͮ:�J�����b4|?s��w ��CZ^��6�G��s��{m�%&�p��(�ɑoSV�nw�)�>,J���g��֯lXkD���b��+%u�wX����%v:W"�%M���Q����fh͘^s46�vԮ����R�g�cb���w*�q���EK1ù#����fZAv���<�D�Ȧ�c��h^K�h,gZ�J�02�ד�3�f[�̻%4�mnҰ0�m3�85m�%`E���|�lUK�3�B\�\šL��6M#�e����&ׅ���p�-ږ�+u��b�I[>Ţ��C��7.Ns���x�qn:9��^ӵ�I��"&�呍�;8�N�iB�ʆ=��nLnэ�%NFJm��n��i(�]#>�-��E�M���]�EZ��j�f����,�..���a�v:3�T\[V�]�;|��yc�\�E�L�&�u�筷!�s&둰t�12��=;ҏAռ�]��8����er���a��rN'Q���-ӌ�[�7]֨���>���Z���v݇����Ӌ4Y�5��+���A鍌�����D�0�L��]���#t������;e�a���⥅�F�nҚ��7�{ŰԄy�PRf��kȮ�q�6T�L��a����h̵�-�/\�������+�Ѻ�x5��^�<��%�܋õ�J�e9�sճ�㷫;�1�1�]���Y����#Hv'&47j�7Wj�xt�Y�+\�f�	ۮ�+(�:�	��ؙ-#�1o���u����%w&]�kR�Q�����U@��<h��Jk>a;�t��خaC�'Z�Gg���7G��h�M�v�N@%�uF���`u�����É���C�3[]A�i0�M�l�^-w����u8:U|��\	�Y��ָ�t�<�ȏ-�K����w�J����N"�E�qu��e#��r
��ss��㹡���ם{PBG�8{�m�fKj�:�dկy�g��͆Vږ౎#���g��&ì�k����u0%������ֻ3"�:�p�5�MN�,�Mk����e���Rs7�&�^SA�7���/��G]��m�|و��;�z����T��=��l��v\ں�0[��HA������2�����/m�c�g���G�����*MÎ����u狹�u�v��,��tat����˟�Aq�H�����ixa��i�����*W\�N6gn�=���M�+�ʐv�J�Ʀ��ls�˄&4v�]BE©yKe��Z�8^��;5n�씺��ņ��k*-]�5H��c%�l��R��F��+۱
��ݯFS��݃���Cl�s!�f�\���݈ۮ6�����$_<m��0*G@e���!�S���,�mѮua!Vl��Z3ɍ�ɋ�	:&t0x��e+���<K�!tz�"as)c3��͢
�r���7_��ݏ����:��Ͷ297�Fu�)�2M��`��-�
G,_��kgD�i1�$�VNC4̼)����˕+3#:ݽ� mKp���ۄ��4٫,�:,)��IX����\�z�V���c���x�=�ʬ�g���S���.�&���B�vIHB(��wxWǅ�^[��x�<tteR���U�m+2�ްC�J�K�Y`ܢfn�;D�Pݝ9@��Z�{c��0ӣkq�nNN�u��쀴�Llc��u62&m^�7:bm2Knn�D�렵�rm���90Kn��N��	��^nwin�cc�f�N�A�A�%�5�����yv�19Wu�T9�6�@%q�����hй,��b�WvOna�cxz��!�ܞ�c���&�ħu���ސ6�b!���i\V���%N�6:���Z��MҺ�x�����,c�{H���lwmՄt:�6��h�)\ʙ�XM� 3M5tt�e�w�Ec����7k:N�MۡBY�۶�A�֠���oT�D�N�˺n:�qmǖ5,`#�Z�!Z��X́6c�\n�]/.��ټ�l�/,��YM�.t��6L�D�L�����a,��.�&�y��3�<�G$dlڗv�pqn]�ι�=�|ڢx�WX:��^�8�5sn�:]ʚ�m����Kx�=}�N��y=�vԛ
���1�Xb�P��A�՞��6�u�ZN�{r�qv�^���zB��cd�r��<��O<g' P.5������:�kO ]�	�9V�/�y�|�.��L8Ö��잭���d{]864��x\{�fgt5��q��j�Dq͗펱�Ƣc��5��X�p�ƴb��&{' l��f3��ٚ;5���N��R,#Dl�\�:���j,=�>3�{=��r�v�Kȑ>G�������= ��	;{r�t]�]n�s	�v�Z�njO6�Y�x�J�׺��јi�0m̽���5�r�Z��
�b^4�J��0*��ốzC�Zz{8n:ɱ��L�/d�6G�iwnݎ���g�H���j�9�-=(p����]-��es�;��q��ɘ.�%���<��xÆ	��%՟qo
;]�4�Pz�&�v���u��J�iD�MtQ	��	����h2�^`E��)Z��`���\J��SNU�m�y��L���ZE�[I�X.C-��Lb�v0�8n3�vHۇ<�;��s�t;ɼ=z��n	��Z1,v8{,DX٨��v"R��4 �Ik�Pvl�%�m#6��+5-�łku��"����%js�X�� X�Sq�2��H���gGCE*��7`���R���+��0f��Df.�r���s�ņػ05[u�)r��^�"0�ڡ���1\���Fi���a�D2����h| ��B�Rv箃��@�w�:�]Q������m�+^B%�jヷc���܇bt���ץ磮�9{]����n/Ip�z�sl��b9�Є�v%��%�J�H6�)x���MƉ�-�
c۾,|�uI"p��=����s:ܾ���U�;s����RX\F&��o(0��.{7�Ҽ��-�2�d�tİ��d�J�[.����r�E�m�/9'v؍���q�m��7\�u�8;(����A��sua-�+_6���u�d��qB �.�-�g��׭f��p;�7Fm�r/�֪4ʛ	4��#m�[c�qLpG�����6�9ݦމ�U��H��P���I�O�<n{
V��P����kv�����c�r����JL��i�RY�Abq�V�7@���ܖ��X*�:��-��b6VSJvKn��_'n4�[m� �v�	�1�x�Q�!˷<K�^���w!�s�\�Bۗ���ﶒ���3�ӧ;9ݣtL�t�J�J����y����xQ��ЙmR���Q\]��ۓ-�y�	ua��X����U�݌<n{N5�2<gMZ,4�����{8��ƶ+��3nC\of<N�y�Ġ�.WcsGuf�kf�#r�q6)W�2U�x%��z݀�<�Z��鸻0�l�v�R��s�Φr�D��K�*���+��=6�s�u��r�8Lt��Z�6�YK�0�sO3��l����rrr���+����S��e�Q��-�8�ۥ-!��8㎰w�n�u�g<�c8�c.��[��6�Ό��첣�CBl1�ulйã.��!�wRB�::C�ܴv݋�v�B�@'1N��:u�x��^�Mbs��c�؅Ab�U�M�Љ��S�(t�<���Ǯ7WY���������u�i�V_Y\�Fo�o	r�p���z�-���Ҥ^�(̗M�4e�q8ƅ㢧��M��.պ��\��f����R�mh�����+�z����w@���t��sԮ�sƸ�G�B�C���m�cu�G����Y��cO���m�lȻ����Sk�ç�s�[�I�v��[��[c�R�Gh�3э�8�4�|�+����83�mg0��֑���5�y�a���^���ħ/GeزV�<B��5U��
1+�j���'5��1��t!����#��p���!�..���^��x�:�cq1vM���k 
=�1��X����]*�(2���+��6�X�-��lJ��4�h��&1�$U�2�&Ĳ�V4��]r������e�Kri�m�iYG�S�ώ{1�x0��D�ٺ:4щ���v�9��dZf5�Rb�Smb�b#7�&6�ݓ�c[.ݱ��[��l̳S�Il۰v5�4�A�^(�3*r͛�<ӎ!��ѓ���p�;9mttv(�k�q�iu�Z�;pH�nI�q��5G��;��ƣ�㶐v��]`�+q��à�Vƶ:49n3�JYB2�Ͱ�\����q�|g[T��Y�a4T�)m��Ès�v�O=�sz5��/]i%lř��f%,��/�[�yt�3̷&�s�([���tL��ӺN��:��t�ӺI���P�D(��P�$�D@�C��J�O%ll��	\�d h�Xn��vE�H`Vһ8�u�)Dg'�����v^$�f.��܇Bgc:Y�ֺK�E��2�R�1��d*`�0��֗LMXh���= ����K��[R;Y�����iiA��k4Ŋ\�qhǍ�P�r����E��źx9�G���vܻs!�q�q�����;	�!�:�ϝ� 6�n.��{@�ϧ-�#��@�Z�Nx2���=�.c;�z���g�9��a;�umdm�:qO9����I:�^s�n�R5�Im�3�\������B�LǛ���YR[��n̄c�-mՉ	lՓh�9Y�-�V�	b퍫W�H�+s�\]�k�dz.��C��yG�<��v�=$�I룙�����.��븸VV�hqH�*����4�ܹ ��<]i�\�bއ�ݑ؁=Y��$v�T���댗g��pj[Ӹc��%���7Gk����<�b�=�#i}����ƼV�W$�^�s2�	r(�\3vC����X�\듋{`���qp5r�\�;n�Meb�,�y� ʘɍ%������ú���6�1e���S�p�&<>ݺɼ���i�	�^W50���h�f��@]���M��S3fƘ2�R案b,2ƶT���o��b�[�m��l�����rq��Jq6�9��V���o;�g��^��A������=1��C]�O��z5��ivB6��q��=u�l{pyO4X6.|�&s�4xP��Z����n�7evx;�����zc����gsp>�^�]3`]�a/mp`���#�f+&����P���kv@�-�"�7�K����/m�`�턶��y�l�2���r0=���1�1�x�
n�9��b�*�{�*.�5�7e���B��v�ME�۹:�����Yn����h�Ð�`���hcp��0X�{�9-f��[�Fk��8c7Gbcڼb޲����I½N��ݻ 9q���\D��	Hݎ��]kQ�)C*(��7L.%�"!B��Jz��ח�}4K@U�.2���7v��g`���K�ps�0ˍ�aa��IL�SF�D��x�.Ék-�Es�nt�;�|�$C�붃]�p؋u�����>��@u�m���;kGxɅ��u��=�]�@(�ڷu��jv[r�RXh��%�z�a���\q��K/]�gC��ݼ���E�>@�@��GNU��"��5���.��!;���w3\���!!��:��^k�ERIP5@�����T.���-:R�ݶ\�L�V�݌vL�$�x�2�O4�r*B�y���J��l��8~-��0�-V�wb�α�B�����}q+ݱBֻ�n�Q��үw�os!�H�\�_������H��F�F7&`ڳ�Ǽˬޔ��Ȗ{��JjYx���ț�G��7�ӹV��f�\��G�l�8e��h������/d�ޥ��k2_ޮ),�-��9�#��N��O�t$�o�z��/;��1���͸�'������2]�23���l����<���	ld����{k{�[Ooa��<@���E�ӗ�>���n�<B���j�L[έ�1x�7�D������9R-U{Yq4m�\���1v�n%.9��!(�!����{b�꽐j��r
�����{ޔ��y���Cٗ�&3�NAb������BjF��XW"��������/BV��h�Qi��z�L-rl�Rpf\�B�N��Q����՛ye	O�F3y]�\����ew���PB=�c��E�,H�T�v��ڗ4oݹ�j�B����}_�V��Wc�][6Cݜ��n�g�q����(��l�ae$>�a2�8T������Gi��T�Q�Ԅ��x�P�:_\���͖d��{pf��U8�X0����!i�TۙO:�L�t��[/7ף��o˨iY|0��'/Lj��<��XX�>�£G��W�n_�G�_m��.e���z��e��}w�����=�?>kF��H"��s�]�|/��
[,%{��=,����N��m���$ -��D/�6�����<=ke�]ɼcbT�]����]�ɶ�R(ܝ�����ޱp#�λ\}���p�y�Qv(N�9�Vo�����W���}y~����3��P�m��B2A*����{�fft=)%(C�8� �M��R�ұ%ލ���-z�Q��'��A�s��i�h�c	H=~�Z����4Y�K[�'���T#ԯ�.�i:����rS�M*;���3��� ��Ğ��@�`�[�+�tg-Xn^pbU�*����_mЋ�]ػ��yr���C�!k��P�1})nG(�{���vn��-m�|�v�e��:S�κU��J��J�aݥ�ޖf�4���F|�h���d�5��$� d'$�������k�}�%z�N��w�jn��%l�2�"��.��;�x.|\އ�qݖ�'�ϝ��ޮs)Jw�^*���i���i�T@a��U˸�ۍ�7N�4n�)�xތ��l���ݓQ4��z�M��m
����hI:
��&6����6"�譱�ۋ�������O:�>q1	l S���g����t��z��WQ�ֽ\��Gg\xv�'e��<J��};ܰQ�:���}�V��Aˢ\D����M$r9Vm��I����f��;���b��+�Ӄw���w�I2��C���ۉ�ݿo{�ߖ~m�R+s`G��P��׷I~<ve?]��S=��S��3�9�/��۪���)؝��ےz,�a3-�H��]!am�̭Պվ�e[kTP�}{��p��Aγ��1���Zw)��G�iY��W'�{�_�%`���"AFH���1�}�*�>��
��e>�"�&ov��s����v���.����~�ԊfM�M�0�7���d���i���4�(� ��v�k7:��ts�,��-l�����LV�.α!�N��%�����%+v-T}��~W-���j�I'�������Ď�k�0�����V�:��Ԣ"%�� �Yr&�n�(��={��R����W�e�d� �s��Y���[~�5!� ��|Rt=5�ܹ�oy�ǃ<��P�!.!	$ϥs8�>��.t�ܲf�a�AwMw}�]��{K�|�V��v�����1�~�v.�(m�X�H�����N�vr���E��(L>Y�)y�R��{�JX�\��VUb�ڽ�e��/-�k׭�)(���\ic�wVa���fu�auB�(ќx�e&�d^�j��w��gzT#ˇo���C��^.�Y�ٻce�u��S�Wf\�s/�Y�zk=�i�A#�1��a�U{1�-��:�A.�"��j�9sd��=	(�I'JFCݘ������t����T<]j�"�9(^͌�#0v�q���m�V��7!�xՆ�vt���9ϡ�Z�7h`���ۦ��cO�`.{o�
|�pܯA<�v�v����z�����]-��×�,�3�06�t\�tAv�����\=g�HL]v#��B��r�[��vܹ��Y^JCf3)��]u̸���w)��$s�x|V�ڔk7>X�N�\���v�Fl#�G��L3 �[�+3�kr�魔X���ș��ޜs�4�u;�c��Z��Z��2Mm�[ޔ��'!Q���hKW�;�u�$���^Z\���Je�z�"���[%���gR�ڟ��s����W0N��穉�)g���Ѹ��f�(y�cN���}�l�!f܎6������Dus��o׮gv�։4;�LtXd�l�\}�P������I�==���B|����) !ț*A����֜=���*�4s�Sl'e��~�2��"�]i����u/��>��6��&�*%�`H�1�$���O��yyל|�ٸ.���F�G
������R�W��L�&O�A�A�D/���W'k>��^�(+-F���#i���]������d�f��X<˒�ً�JDn3�a�@����9:ǚ$K��V��������N^�����e�қQ�z�}\+�[
��۴7P%*k�)�$A?�RAW�9�7��+�2�Y�,��+=Kn�NZ�W��S��mɔf����Bb�+u�ѷL�w>�9�*=��Ag*�$�Z	�J3���&���%A��ۨ�̕F�3�t�i��]:ٓ�oXyY�\0'�`�a�� {�$��]*V�U�c`���W�̕�}�ˁ���i^>�-�%�8ee�k#�](w��D%ռ�㔤Q�#��!�H-ˑ���(��Y��w���Ox*s�v�����$Il���R�f�����Ԃ�t��;�toå����a}�)��I&X횘��p����`ل�i���;��ww��ݬU�l���^m�Q�z�	6���랬���KBm���І���As���1 F7�KDck�Q��k�E�4�f�
r"��A
I����du�X����ϺĐU���L���/p�KK�d�Ͱ˔�o���؊*4��Ο�t�����v�K��vR���Ί�f
aW{)�x���<���;��N��N��?S�*#j7$�~�nN�}/'L� �=���S��!�z>}H��t�׺�y�v$)�'\[�k�=�V�,v�HZTF�u�����!��qww���"��h�j�훳�㧁�(�~;�[;���C��t�iW�+=xE!Q�SnOq��ܽ�
�j��>ۍ#��v�P�'�߻����KIv$�E��Y�糷�a%N�ۼ��n6�L�T@��Pf;�ؒ�^�َ鸞w���*�!�d�r��IF+��n��0b}�DO�n���Ȟɕ�������F�U|fv^���M��1l�5q6��YG �.��ȱ�[b��͏g/8�;a�0��b�c�;�n��5b�m�m�_o ��[�(.�:~���͡�׃��a���[��"ĎZ-�b�����^��f�3N��si�]*ƺG�f���s��͟@�Z�Fj�^ߍ�'/'����&T	��II%���.�Q�`��C9r��pۧ���oG��&���j���`w�~��zZgf�:�6J�6�aG��gOL�
�y�O��mxny��r���T�\^N
49�@��yC.���y�w�;��c��}G)ߋ����0�O1�{�Pjx+��o��x�f*��������݌D/�_4>6uk����7�Te������1)#�H<��;3�m���^�;k=oB�)���i��g�
�c&��e��w�c�ev+"�3�U��k�m�n��B%�r��Z]��k3z��\�
v���e�v�Mշ�Ԑ�[r;:Ui�~�)�_�g�	��լ�r�� �S9��Q�-����,���%�zq5�~��z���~߫�|ݽ�����/���=�����QDt��:%:H)�n�u*^=ԕ�k8���}=��~�z󫺅P�j[5^	��0��Zq!h� �|)�M��bW\ث�κWM�^�B�gӝ̆ft�	���T5�=K�p������oJ�a�Pn@�"�I��A�����69^�6��_��\�V��) ���G�ɠ��בǆM�z"�(#BFd��e	�Wg\� ���>�rc�g���78�G�JNz%���1�M^�.u\�O�V�7���=�(gO���o���S�W�l�fZ�����K_X�T�1��ɣ0j������HrwΘ����,�lk�j�m�m/(�m"�Q�dy�����.+��8�^w[�r�8���8 �h]���Ҹ��jg-��,��J�!������3��B�;����u��$6��^6���N�M���VU�Y�$W)�Qųf2����3�VÓGƂf��YR�����-���M��Oe��z�H���Q�e!x[Z;��Ng�u�t��5lQ���t/r-��-��e����(�%z�FB6��7.خL�sxuR&���H��DM��&��<�j����l������i�s��-��[��^�(�����,~p��
��Ax��bPE�Q!��w�^�T}������t֭��٨ia�.��w�T6O_lym�[��ӻ�ު��,���Aת���?6�@�r��8����L�ic�6wO,�����&_J8���j�&Z=���X��Nm�D�Hl4Ti��3�'�;�+~$�����wF�z���n���.���^(��/g�&�{�gm^�W��g���'FJ0a4aq�%����z�5K\8�q��yo����r?��O`ʬ��+MYў<���]�LV�6�p �Q�b�Q-��Wg��#[4��6�M��i�0v��zn�۬��8"�ґ�����F~��x�y1ת�41Bk�ܢ������!����wӥ,�i`9�������2�:K��;u�z`�&�)C$+0W��4[kk�`R_.������>o�5��M��t��r�.��o��"6-�:�]��7��/�6�hP���T���ݪ̊�<�����*�6��<żo�n�tm�<�����A\�F�|;',������)]Z��&8̒x��py�M2j����c�X��zk��մ�+���n��>������Ʈ��ȼ�y�ʷ^Z�E�pH���Q�x�G�(��J��U6,�tU J?W����L�[-�7��#1�[e�^���@�wܙ�x��:}�L�ͥ񀈢1�</M�����⋞z�o�9c�WW��g�ٓ�z��v�ź�9�r(�)��.��7����!�fmv\!"R0%3v1�8I�4:)-�vMYh1��Mg�1�;�����bD�������2�uM~%ذ�poRY�f"��
M�;��\��Aw�������\%e���Q-� �Rx
a���&���!����=��OA�7������d.��x�"�kk��g_�1\���i�^��u���ƚ0Cp��I3#���2#}����A���!Պƽ�]��G�Z�������� ś���Ct���e����j�y��u9�*��E]���keȈ=]5���L{QT����b�Fn�Wv7��m���-�5ί���|�9�R�8�T�[��ٜ(>?�w6Ŭ�|���N@��|v�PURZ�Iڮ�����,Pf�΢j��Z�>�j�v�7"<"�K����F�ZI�c�㵦7��"]� ��2�y���Po�,���%ie�t��L��� �����z�)���aC���ȷm҆�ӭ3#K	�l���=�EN[6�(��C�{]�(�Lv�wp2���7C�E^�{�WPޛ|�X�iKY������+�h/�ʙvI�H9u�v1i!�RY��R�6�Q��Ԓ)��@⠱oM���w+"�,֡�l7�bl7���rV��	&���ev���݅��č��O��/!5��lu��w:T�U/���b_h�D���Uة�m߷u�S;���n`�S.�:_��,]�j���Wrv�R�>ߓ�K��ڬ6�e�������wGw;�[A]���9�Gwt�CSu*k��eCC�3y���Φ�r����0(*��ǃa;�WY��ݭ�`�쵓�h��E:m�b�W!J�1��ϫC։�<Gz���>���f�P�	ifF�ո*�3;+h,�t%�����S|A����3#��\�_<�ҭ�\�V�z��#���(�:YI�/q��L��������x@l�9��*�����oS3�31��Y�!�U��<�l×vI=˯�G�ت���y�X8qQh��L�<��ג��h�涡�$�?Y��w;W9��u���M>�I'�{��1���aN��� �E̪�"�_4Q�$IQ�M�q.v�vo� w��{�Lk�G&א���R����0�����v�q�T拏I*���B�	I�x�b��n۵d��i6��ؑ�ʝ�{[Sm��,c�D�P6�PD[��KΠ^^Z�����S�%�ϸ�6���Tq�|��[N%��m�Wx���{4�Kَ�e��#��p*���B#Q�Y��%٩#3��W�U���xHB�j�`��3�j�, �t�_F��SझW�~Sj��4�?�l���=�Nͅu���*�G�R_�Y�����ڮ��NӨ�+h�^�ŎZd�m0��tmok�E�S��g}N�e�P���$C"9�U��(q�s#4��8��Y$����t��wq�GX�v7�^2�Hs�n�Dt���Ӧ��t�;zW��(��UZ�j�Ⱦݗ��}�fb�z�e��_�ukq�^0����w�o�y&�,+�|Y[+\ߪ�B�G5@�Q,��
�GN���O1T`�oES���9�.T�u��c�W��E��<��%2DI\���yK��-]cX�����<������ لvң]Hgk��@�hf��:�`;k31��N���ۭϬ�h�\'�"�V�'�n?BF�K�˂{Bz[��}���wY��#O�!�]���x^cF{�R劊4�XB�gP!�
-���j��^v�{��f�ҵ�ݍ+\�s�
Uc��kG�Q�fV��\�w�$�*��O^�%��r��c%��0G�QG�4��{�ѓ�R�]_���Ы�5c��j�t_=}Tq��VB�! q�=��!j7�6ܙ���]��o�m.=}v��2�hX�s:����H��K�e����ye�ԑpo��;Q����1"8�߼��L���)����Ͼ�ˮ�Ѿ)���ޗ�'Jۓۗ�u��r����'�ڹ���Wh��YI��8������'G��F��,*�+{�B�M��-euM�v�-q/Y%+��;���k����R#O-�%�uH�،b��e��h�B�m��o��a�ﻵ�v�,g�Jp6#n�9C��:������.4{\r۶�ܯ@Z���gK��KSCefl.Ѽћ�l�+{q˝�۩�k�ܴ!��R��s���&�	��[�DȚ���V.���d�um4��L��p��Y�wF��6�)�ݩ��)]��2��,��^f��ã�|<�c��ͥ�ʲ�l- ��X�k��$+�O-5�3,c���i�1�-��Y==4�ٚ'�=,��D�w �����E���n+��Е'א���P>���}�֎ٰ�"����֊�\Rԋme&�&��K�ly5ކ`�3���ݣ�$Eլfw��N<����F^��~����!
@��2IP1�ݫ��gm����\.GRU������^k�m�;UcLN���.�+һ-8+�h�$tI�N�5$H�%��xV��ԁ�N�Uv��݁��I5v(܊�4�\;��0nfꑟz-�\��KU���,������*A� ��\�{��̵��N���|B8''�Fѷs�����ط�,=�a��wU��������T	<I��(�8."�I9�sۦѐ�3�,�� ��3Z�a�1aM�F^V��c9Y����~��w%J�X���ɖYi��Q72�eQ�!�n�0f�����s����-��FlD��=|�߽�v�4}+G��ͿS�ٶ��([ֺQٲ.P4��B�M^��tU�y���%f�veZ̀��}C4�5�ʇ�'B���<���7����{M��;��:����ތ��ņ�gV����yٺ����4U�p��d��7$����m%�%�C�S1nj���Y�����z��ʭ��Z��vX����0��u�۪\ Ja��$��>WY�D/4�֪���*}*y�s�@�l��@���M]�;�C���y=L��t�w'Ev��*�Y=R�^���RQ���i�+�9����V<���G�,Ϡ�1F6n�eR-i�6�H������$~�M�Pr�lI��#u3��b\A��m�n��l[�pEg�����/�2E(4Á�%��Uh�͋ޫ}gM����ݷ�>qt�[��G�{X�NH��ջ��Gw�i���U�i#�B�&E�ȳ�#\�%����� �r�m�6�n���U~���$%�S�%&l\��{�Rv����H���徼�0/sq�Ӏ��qH<	��������::����X��a���g�Á�X��&�d�άp�kΨ�mh۲hD%`����Ncu� I��X�뚰�V�H��Kd%�r�r�ȱK�Wi�6��U4�뚏�����ޕ\�{/I�he|��0�-F����T�<�e*�����ڹ8���Jup�vʚ�>��C��K`�	���j��Gu���x�<�@}��
5����¾��3�?~~���ߎz� 5����ԩ��l���+d���Qvƍ��S���C{��!�ޯɯ-�F�`]��նey�f"�`]�.$	�.�����5SZ]�3J�2�L�W�R��|�v%^�"�SN ��I���f���z��>�<�e�T�+Bқ�<*��e��5	M�$�fv�������;ly��7�Ɩ�N��{����}��,n�� ��B��d�նi�t�X�v�PO�r ԃG{f��f��󥤫_"�)�gM��Y���G������ݬ�,r����^ry%^��)����]���J�0��N��]��R��^y3�m��h�y�9�s⠙[���\��7��m�:��D�~�A查�F���ڧ	�6�-T�v^T�#�!��?M�Uʟ("�g$�Υ�,�|h�zb�05�l�2�k=.��E�_U�0h���$�!q�~�.Y�.�݃�U���QE-����5vo(���6US+�� ��ɍ����C'�󠼙(�{2���`��e�ȉ��F,�������z�kRظF��u�й��v��1�$@��Q�� ��R�M}Z�N(�tN��&Ž�M{<ur:�M]�X��
����)W�j$#,��8inf|{��$�]A���ʵ8i�R<H����r#<}2�Z���y�X��]�&]�YF�,K�WP��D��I¼d�Mm���HK�>��}V�O��T�(ժ]@{s3W���Y��Vayү�j�<X�W'��
BDn�� �=���,	;~��K�$���1�G��KU]&�zpVrf�Dz�:�/��'?$�s��	�H�$�a�ⷻ+�����o�n��7�͙WM��[��w��>�D�����w���YY��{e{��a�*pҙ9�T���g:�R�m0��q\�ڌ�з�+�6+���:�`���Q��0U��x_�0��S�L���$�n�lqmnvۤ��Z��M�,ғ@��e4&�^9�r6�z��L�l��Ƶr�X�����@���p��u�0Zu��n:^s�b'�r�$�yњ:vꞀ �x�نH�R��k[z�Q��Gj�feэ5��g�on]F��7a˳�t��11mi�21�4��YJ!����@�����zt;v�]=�p�v�7��Y�2�F���b�,:ʧ��8��v���V�C�t<�����R�M��M��nE7�g�Y����\_�i�D��'��kw�kz����t�1�T�h�W�>��b�r;\��돽�w��})7�K.CM+x'[/��͊�^o�XR����5�_-�_�V�5���>�S����Oc8�����i�A�~���k�O��h��
$`F���]f��w�a�klLw��y��o�����c�z��Ja��jV���Oh�]n��e�ף���n��B;��ؘ��w�S3v�Sv��sa�3x�2��n���T���Q�A�(��`�PrAG1E��\�˳��IчYZ���o��z��w\{x6ͧ���^K3�P�V�V�� ��#��,Y�B!�5Dl�:�RR�&���M�R����\1e�I�i��¹����-�.��K)o���xm_N�"�ם|�U��7_{ `���b��J'��5�^zﲮ�Tm�]�3

�R7���+ZD]�1���Be���~��.8��w4��u��0ݜڄ��X������0���v`ȍ�����<�U���V-e�8������i����{�y^�Ȕ6hی�+��ǔ.>^��k'���+I2��H�JG��~�ѝ�,SP�5ބ^2^_�ɝ��G>��I��J7�4@귪9���m�G��dش�mU�4*+���n9��ϧ]f�J���
�.J����y���N�M
�6��͜s�nn��0��(�N$B
Ddr?�Y�E�abl�ޥ �.���:�m����m�..�$GƢ=�)��&��Q1�Ն��y�����>��2�7
cmh�R�,s*���g=�c��^��H̚��K[YPIf5ZIF9$�K�̩�v�:�-�Wc-J���wm�$�;�Q8ޤ�^�n�E��M6�i-��*�9�$
��{�����vq����H�/od�h/�Ԛ��k�z�}(OT2��&��7�X��GB�I�x�'ƍ�=�%�}�Ťެ��ݪ���e����XٗE��M���꒎�ڵ6�����7cA�A�YQ�(&�[V�=�Dsgg;pY<��'���*t!�8-��\��NC�謀�І�h��nI�,~�YC%Ycy#Hb��ܖ��ҷĄ�/y@y��C˼�:nIB���$D5:��y�v�6�ׯ����[�Fm1r��{3[r�"m�=���3�V3�����p��Tͳ^���(��Q�����/z���C�6Mye��H�������F��4��+�VXS�3d�j��+X��P�����&�g�{�����P�g�{�]��^�Z�k�y�n}��A'�:�g�����Z�9vZ��c/�P\c18�-���Z�ۆW�5�(����8����J�ٞ�t}u:�جa���3zǽ����C5��+����1�p0�@��qx�a�Q�I[�=v���Ce����H=$u]��jl�$(co�x�A�<3M֜ח�G�I$��jH�zcԆ�[��U��}��e���n��}���N#�n�/-�ίZ�Jy�Wݍ��C���w��:����ɲ�V(�VS�)DwL8�!%ode��^gf�����<�c������Vz�r��DK=���[q�U>LEO�ڈ2�-I!5�I{��}�e��B�������Imf�-Т߬���,�9`��vl�㙳�������ƚipk�X��f���@97=���]���s�\����5ˋ΋�l����f�DRA~�r&��r���U�ޤ�����@�v�Rrچ�v�;z�͘�mP-�Ь�;�<�(���B�P�m2NIhEm"V{v]����n�~��B�ǃyw��>��:!�|n�y���7$��Ps�?D;M�.D"0O��7%۳��;
�A'��^�hٲ�w��R:iGc��T6'
����s�F��"���!:�z��-4���K���\�E�~]ٛ�U73 �
Dcp_�ϙ�F�E+�ᚗ��h�Gw��Ӣ��ؤ\#��:�����<�~��p3�
�U-�I��c/[����� �p�����+vޤ�ޱTGs�W�3�6;HWm|E
ȡ�-+�y�i����Bq�ே��F���BbV]y��ң��%��W0�]S�L珷ϹW�-!I�$P���\-!2zZA$/��د�#HV�sZTpZ�r���G����)�n�կ.#L-��ZoF�J�R��I� Y-Ӽ��=(`eк6>��[��ͪ�Ԍܭl,�w,B�,��h�|ot�rзڻ��j�d��w�2�W$��b��~t�h����k�/����}_�iI�f�
y����H�̓�&�;���5nmq��� h���#9n��%0�7x�ꦵ��}�N$L8�LD����.�������WѮ'jY9��/pM��WFUĊ&�i��Փre���'��n8��o x{ zk�+�A��0N/���;7�bLh��T���,u!�=C�$���0�'�䘶�԰0i�Wevw=���M���'Ԇ�Q"�8���ݯj���r�ʾ��e�1�%�ʵ%�D�Ԕ`gs�cτ���㜢�ݶ���@y2�C+է���*N��
T�(bG�SR���g[�gf����M���]'c���$Yz/r�}�����c�H��ίsHѢ��Ѣ����AV�3R�}��V�06�|8�s+X+%H�DΧeހk]i'���'d4��o�b	��ׯx���&gSF��fU&k*�d}ם��K�fԱ2�Z�X��ڲ'RW��4ln���2woWN����y��:n��.��O"�yvEԄ��99�'\�w^������=6�H�ʽ}ub�E]Qs�X%��8���|�x��і����t
#bKs0m-U�ͼ� �u���t����e`�)ւ������}�9���ݹ�/L/�fP8P-�̎D� I+��jm�����(mg!U�@��VTȺÇ'I�jwk����ϳ�s�� p��\���d�{36)L�-eU P���(�xq�K^�W-�5�ƌvd���\�=�tؗī�8pyݖ���%oNyQ]tɽm����wq������)o�J�F]K�^�3k�W����[m��\�!�cûN�k�=F�LX��݇2.̓�a5i��Qk��t��5�U�4�KPȴ�V�ZZ��F�sKfW�Q�^M���c������x��jEq�x��y����`��`�a9����4訷�|�y���t�Қ��2�RɰB�Դ\my
���{cp׊�t���iI���[j��"6�m#I�Ke"e��k�:{c%t��_tu�ͤ�R�;+��,i6B$�nn�^��!�:��pJ��.l!��H�6+^ؕأk��^�/�/f6ne���R7:��\,��M��n�BZ'�u�aȀ�'�t�c�.:C4����y�D�E��K�(�[^�6^�N��N�N�nY.�N�.�0$���bMvt�@���!4uLE��aijSmA���%���n�WbiYbՎ(��o8჋��k�˥�'[�.㹶���Y�:����p��ṉ�^�ִnϴh|8����gCr������v�1�������KQ�\�6d��f�r�NJ�C��<������U��inýjv�",p�����v�)�k)Ų�@�8�*�θ���t�Q`�dV����@����ƽFv�}([g)��Iۣw\������tq���+ۯ6�=�aZ\�nM��ǎ��t����rq&ٜ��6T��8��7Ww�8��;D>5Y��Y�Sj�r��W��Ki`�J�G3D�-l"=7^��C��g��t�g��l�h
�1���;P����-�s/@g�y��u�2��r�C㥫6X��ok7-U�V��1�kbhY\`�q��]dN�5v�m�f&ZF�ljQ
�l����[M�d���/]���L�^ܩ�����z��pj}�3m�nst�]mv� S������� �n�Mvܪ<�m�չ0���\�]�ŋ2�N�
Fa��J���3�M����ܡ4e0$�9�Tt�7I�,y�K{Q�3[mes�a�[ڐlJ��9�m��۸�8�O8!��>�ncv6$�ێ�E��뫀z����Z�gsװ�zv6�91��nP^�힛<[m\�[�
�M)sU�GN��z�HTLJq��r��{˥c#�RB���Ƕj�LA��GD�c�B�h���x���=Ufʺ�^7Olӂ��-�`�].�rX��M��Pz���`Q�!��H#�#���>m��L:��uUzD�A̔����am�B]�����VF�
h�2~���x���`X6F)B
>��
�"m�k��`�,�)�W*���a
�LJI ���eֈ>��8l�ܾ��2v;��osݓ��-�{���U4���B�j���0`E�"O[R&e�j�2�ׅec�Ս&H���]l��D�I�G>�/O���8�|_	X�Y��V��B��i]���p�۾-w91�+�����R4CL#!���~��?�J/<������|=�y(l�k�Y�㢣��f����d.����a'.��4�=�W �\
j����o��y���&�|��&G��*"Ȩ��}���	'ɖ��Ʉ�\W���ण�Z�ƹ�7���ii�r_B�����g��,�տ���@3r|(�R	&@e�G	��� ޲مF���RX�E{���Z�-EF����<�Cƫ���;�C-ل:dm��sȜ����œ�ڔ�������ϲ�ڙSE�l��,���g�y{²��]5")���qZL�^��ł�p�R�Q�g�^	s��dw�X��a�BR����T�}֫lz{)���IP�-w��x�߽~�����B�N0N�+O�<�<���C���.� [润a�Kj� B%�S���WV1"P�l�/����V�O�]p뛸���j��_ikoR�N59�����!.�V)���e=I*Q�*�����d�X5��h���ۛ��G���A�޽i��r��1�����I⩢}z������Q�YM���N�[MT��±�:��U��@U7NvYb�>j����G%U1˔�˚[�H�h!I"�QE�su��*�����=����%����&Bt����|��0��	�-|3���q�tN�:P�皡f���|!zkڭxZ�cVG«p����*W��
eR3	T��|�� >��~�1)�ͤ+G�y��p���Y3��"E:���q[#���Y��YiȔ���Z^˞���X�{W~��H��d���}Ul�}(�8���п�O_������0�r��p\56�\"�R*���x�-4�$*{�ڢz���_�Y\T<��\/�}��"��_
G�O�괾4�$&p '����z/�;�G�d�m1��R�f}�I\�p*�J�T�
iMh�h7����*�0M��q�c�%c�Zܭt�ԓ�U!UY������^(��WM11���%G��u�	3��E
�uP�ϽU}��
�JKe��VpJ}>�(i&�-G��_;CNr����ld�O�Z���aQ�Q
������Ԣ�F
��,������IB�����f	p^��PfT��9�t�k_#:X�վ���-�t��L�녴�"����-�E|��KD��d]4g+���p� ���$!m����^��h�To���rv�MRī�5Y�`q�u�1+�T1Y������D���c�"�58=���9��4�U&s)x��)
8��n�~U��G{��gpfbݳ�"�U��녊���z��Y�Ծ;�|�,	�X�@��vPη�G5�/�|=�ت�eR�wi�i�u�jE�݀�������k�q�1i�j��k[��
�5?<��i
��L��Zp\#���"�n����/�:�z��@S�����Z"����?ՐSVG�ժ�D��JH�Q \"��~�bVpXE��i�t�I�DGտaޞ���#��d��Q��WH3@��y{;����T��6���'�'���@#�b�8�w}��j��"0虣�(��е���S�wޏ.W��{k��n5��h!Q�#9�^�W9:J��k�j�	�>��Z�j��1O�aw�wҴ�����}�ut��HH
��42W�vyv#\ME`�̩r؋t!˝+��YL���WS-7AHs(sK�H��X��1@�t��K�#�腃���[�Q�>�	��}x%��J^0�ƨ�(�<����-�=0(V-�(z��Q�.����/��v}�V�޸E&Ă��������p�h�S���!��U0�G�a|�A�l
=���|@�/C�C;"��KG�gqT��WU��{ٍ,щQBT}\�����qZViڣ�D�鯴xBϽ̫XpM��/r��U���z���LXP-��$]S�m�,��p�oH9\�֐�]�kx!��{]W��Hⶖ�+ ���Y��X�m�m�xq����p�:Q�թZoE�,���KE��h�>�{����
��v��	k�<�6f�t��.�M��B�N��U�'I�$Ϗ�D2�d����-��p](K���Q
����Q�\�v����d��,iW~繑c�p��F������y���C�'�t�H,U�C���4�גlJW_^�Wǒ�Ά�mpgxJ�|����F��2�kW��1�W��Ļ��<�ܩD�4c٢�~���i~�Bf���V��x��%�K3�)���X�f�Z\8G�[1x+��b��m�o^L<p�֗J|��|�9�s�k���^E�����n:�g��
m�Z��O6�\9Nے��bRG	�D/���p�����.7�H��x�o�Oy��~t�BFX(��ya�=u�c�y:�L�:Ab�ۇ�oRl3u�n�����o׻��C��=�f��Xt>���}ƽ�=Q�.�ܤ�`�����\�q���P����Ĩ���u_�G�ǥ�������
#Z�dkv2��7��Vڣ5�$Y�r�A�҂\#[!�[�����&H �IgȆc�wT���_�Vu��0�o.�G�-�ij����ȟO5\h�{(#�՜�%gƔ+���iv_y�[����EgN)k	s�ڹ��%�����<@�Do��?	�����#�t郪nfil/��9��������}�u\.���4�5]����?����m\,�-ض~��o����m�­��ZS�H�{ެ��ӡ,Y�ݢ����0��¥m|}�`x�xu�,T���IM4���ֺ+lK_
/�b�e�jLhGH�o߲T-��pX%`�IKċ���z�0�s��,�I��V�Xu���{ݲ䆛��֨X+(�߾`�j��2��q�8@.�J�,��*�$f�9<�T:�@�MVF�
ĸ`c�(@��r���E>lBvұ��)j>�v�'�|:>�O�x��E�E���b����4��j��ϫxҒϾ[6!$`ؔ���*�#D�>Jp��O�qR��u�}����}����-��Km�ߜI9ܡS<�w9X�2�h��0d&�]<��-r��;��f�wͷ�{6���}���.�c�<xyɮ�L�ny�Vݟi�oF�d\��yu��a�	n�+vR6j3$XS
ꑴu�T�#]���.c��sے���t�G3�g7L�+s�U�읈��h"(�Ε�`]h�Dp��)	h�MV2�M`�aă��(G*�[�&��]�ػj73ѕ�9�v���:�nRė��b��1��Y��T��}7�T:�����k�r۠Ֆm5�n�V��[uZi��J�0 �,���7�����V�(/�����B�(R]L�q�ڑj�~��l����3�P�<�#?w�p�E���5?rB	l"���`*��(u�bZ�d��|p�����L9�v�]���C.Eܚt�b�wʷϓ4*&i����j�bb5��VY���R�>��W���"u7�}�w��_+����׎H֊C_@���up��1æ־�T��*!�y�ڼ5�t��##	,ZE��v����ن,�Ͻ5��`,w�w9�T@��p�~"�U�i��S�W�[]���I�ҡ ��}V�}�RX!��vz �#|����+����}��ﶧ�u}.���A��Y|#u�,V�.[��I�/}�qZ�rW���b�!Ȭh�S���7��&���Sr��˩���M8F�՞��C�V�����KDȒ�8RB~���b_qȗ-�_�����V�GH\��L�B�is�år��9g9��H/��;V�F�ǅ�;P���Ҭ�������.fn����}����nnd�,�=�ڪ�Qil�"~jńgOr�@�䭶��s�?I�O&��h�}�aYH�M?��7Ӟ���g$Y�iq�f �e���9�p_e͖C!25����f:����?>,&�d��b{��v,Hn��3���|ƋIVc������n����T�R�*�����=�)ǩ����V��W����ҤXw�V�=��ӄW��E��\����f�/�����t���]�&�بپ��#*~/�{n�o�&�)���E�{�[0��@��*��D
�\���MT���d�,\#���� ,�ᴰ	!���Ͻڿ�������o���R�ª���-��z��C����#���z�oq�XC�{�+�E�ՃkA*�`A�D)�o�p�a�mS�d��.�Y߈do~�཭KqY�m\,#�r�i�e�hgz�=�V�[dP���*�p�{?|�Ϸ��V�Ud�W�_N�H�B��V����t��QR
jZ)UUV%g8�"�Qܙ�p�����`����w(lm�$��{��#����w�j�����>���đ�$	[�;Ŋ�9m����p\�gc߽V���$]�]p�b�e��������]MӒ�T��IT��}�b�.��Y�� 0���g�T�}룩x�;c���ai��j�wl0�i��¡T���\/o&:+ TP��8H��9^���=}#EGE�{�rL���l�H�ϹW.�R4ԚIf��`���(��iI68��:T�m�!M�e�n~�٫!i	��&o�"�:~�U����*~/J��w�/��4�e�-�ꔟ��U����xX{ZV%�c�.o=�X�v[k�b�J��?5D+���W�T�W�g�*A3%Q-�"-̼��#�(^d�h�ڱ�`��������f�ͨ�L�uɖ~��6>�S���F��%�
MB���V	i��:{-1;rY@X���{�VaV��,X}���^�,�$�?.����ʤ.�sUGA||.�*�.���ڢy��,O��Q'E��_uN	Q ��}mӍ����n���ݓ�=��7����h�;�ד���;��r���n�FǴ�o�Y�0����U�w��rz�����4��S7�"ġC�~ݧ��������[ǆ���;뫏��<H���鿽��{��zU�}r��.nd��:䢉N6�q9,���Rh�D)T0(��4]�����*DZ~��P�]��FW9�p�Zaƨ��ϗ�����Ի�W
E�K.,'M"�'�AJ�a��cѮi?�>V,r��B����V�z˺)�aY)%�=ꔆ5������_8쵆	X�& N{ܫ�~�VP��c��e�"�2D�խ��+�SJ8�H࿅���2%��9k�vwX3�����Y��ƽ������0����;`�d^6Mn:�~�U� m�ݔ��<*!m=#���V-��ݛ�`�lH!���=�ܪ����" �_�?Ɔ�t��#$�T��.�*!N���6�rS�fj�:�k��<�0�� ]:{t�	Yo=굢1趚���M8L[��?}���i�v=y��f�y�d'u)�@)�]��K��h�r�`Yb����]f��pϾh��L�s�e-!b�M\���z�� u�Br ��պUDuJ�g�n ���ft��kfcY�]5 b�f �)��L˥35]��	G�kV�'�H�Z��y�eZ�x4���S!Y%CFc�]}�Ql��.)N�!Ɲ��}n�����:,/b�N�-�
��S�+�H�IM_+�U�ڽ��:%��6Ib��~= R��ɥN�j�0\�Q��b��}�̞��r�$K:E}��n�Ȣ�iCZ}!:l�/�{�֐q��Y
���"k�}��#�0�G\�f4��Xt�!��y�P�_F��W�y?��S�`���u�[bX����g�K��B&J��_�"���X���}v�ӝ��R��fL�P��^�ݲ,b�x)�s����{!�/��y��}an�h)>K�)�wޭ\�e_J�HĬL�����=�����"�Y�N#H[�;RԐQ��H��X5���(�!��Ft}���}M9�?{�z�+��\�ǅ*I�I�)�7��f	{�M 4.6�i�D��T`���VťK�4��_�`,���}V2�b/��kh�r2�M�q�X��u#��+X��W�n����T��7��r�t�v488���n��>ٷ{z�ɞw���~�ߠ�%ƕ-|-���[M2{�眢Y1$�i�&}��+Hra�V�[���Ss>�;WϚ�|�XC$�Ϲjϲ�>"�/�G�{Á��p���	
q4�!I�5g�Y7��K�>%$�[�l�?oޫX.L�/�*��e-A_���#K��~i���fƖ�3�ѣ���0R+�Ƈ��&]U���
�rDl2ٳe/�OV~�>^V)��a=m{�u�k��t�	���Qx�W��V����B�%a�C0+�Y_�,����~-s??ɭ!P��(R/���V-�%��HtZګm�x��]:�T�UJ\�N��B�6�O͘&F0t�mP��q��~�,�E�~����ۆ��?�~:~I�x��śu�+�W��!�LF�:~G�ҫ�sՋ����H��i-���B绸\,�V�^F�}���%�$~����ϕ&�RST�%7T��0�v�sܕÆ�����Z����� Z�E4�}���bm^ҳ+��^ �����	i��ͨ�<��/�k�Ie���Yi|t��ƘH��xP���p�Ze4׫�IP��[RB����¤&��U%MUZ౽��iih��}����{'�����^ok�^F!e���Rܓ�P����\a#֙�Ց����F�a	���jļp\ �:�JC"�㧶�s'�=�K�����e�E�t����q9��2�D���JEMT�d-0��Wy~3�.�.��#�C���X̗k^B�e�ذT-�{��^�¹�qZ_Ӗ�׍[�
q¡��Kk���%gM�-��,KK#�5i��Wο��E6���� ��Y@�=<��S��������e���%��-�'e��Ģ(��:�R唞-��ƛ�AXU`��ڷ��#���M���l�j�Ӡ�i�h L�&�H��m�ὖ͗���ϖk�7f�̈��uq��5������� �=�4`��;�v�ɻo�aKн�!�M3�1-[i�bLM��4����iHQ����f�Z�{�<�iml0�a�kn%x8�n��7WF7cR\�IC!�30�F[�*��h.�v���,���+�l��{!��4^1����W2��*Zs��ֳ*��6F���E�FϱЦ��Ԧ�YHLZ�իvtf�Ii�5��%ݰ�ػG\*���,>�����g��k��`�[w���x%�p�B�af7
�O����o���F�J�|Fߪ�]� �d7z<�պG�����)k�wx^�WN,TG9�ـ.J���J�:bt��MM,����}0�ia��-��0�])���_!h�)���Osx��
��"��k�{+�|p��9ƪ�`nG���q��E$QbTE[��Q��q_��H��w�p���W����-��T) �tM�2b\�c!����օ�3�&���Y
�>�\s���S�{�ʹje�Q{�����-z�^�~ϸ��]8|%�����G������ޙX+<D�-���X����
�
�/p�R���ǻRM~�3n���V|�����M�k�uCj���~�CC��bZ~mJ�VĊ4�Y\H�~��\�T,7��O�a"G��V�S�|p�6��!�g��ߊ�=t�x�i^W7����pdr�mX.�8� �o�_��%S(a�������)z�$P�W�}�^+���](薿m`"!V�����裱��F�����=�:*�T׆�e��Nr�'��t`&):����5Z�k��p@�n�Jm��b�Af��/g���nt��W�p6�����Q]g��A$0[lN'��"�[��Pv*��X:�Gk��:z���TB�w�)����ن{�p�����G@�o�`d�ެ��8.ӊ󠖙���DQ���Y�\;� ����?$@�ؾ�X��R���;8�^���a	M;"B�e��HtS�T���0KH�J!e�˳�X����b]7�g��C��Mmܚ�d��=r���@\�Z�5X�h���|����C!6�>�'�����}��R�$�]��]�׸��	N�Ϸj�ژ�������d��8�W����.�|�DY�)b�H�g����G��dP�Ϛ�Z�xE9%��(u��u�AyB:��ϫU�mm,-�W��=�c��Օ�
��pL�7M[i�%4ԑDH��m��"Lb�s��!��zS�
hQ���|+N����F�o�ew��(7�B����!����,�(M����uk�p�M�Ƥ�;l0��b�¡ϔ��D�njj�-p�N��Rfc����7_/��~�Y�p�?)S㛫8Q�:`�~�s~��#����y�p���JJ�ư���0L���Uണ�����B��E�{�,煤m��+^"x�Q"$pT%h����3M�MRT�R����+,�s�iIe�	��}V�����^w!B���;��_y�έ+ܫ�K������+�5"N$]s�WAAiaƊ�`�(�$J�~�qj�8�n[��8�iI<��xw�[�p��6B�ȣ	��HP2� [�F��Z���\�2�L������,�eM��iT�sM�E�'��oYaK��[��՞$�~�U��7��y�9�(X��v�K��C��{¾�|$C��G�Q��s�T�{����]�^���|��vZe|4��b��O���}V�i��~k8�l�B�Y��?<"�A<���e/KPN(�29=�������߼٢M�c9J_�s��ǵ���)D2�;�=�X�:t�m�]~���مe�}s���"�}����tIT�]9 ��"Y{ܬ]�����_F���|��~����,�`�����I�TP悦B�id-�L�&�(RJ=�$��_���Y ���ƅ��f?�4M����wK�{���|W�}~����~���{H��	�^�N�d(e�˴�w��ѻ9Gm��(N����9��[F]�n�J�-8f��M��oԱ���#Н�r���K�����E��_�}�v�WfFsR2���hLN��`�8�N.�l�^�3�0������6�[3;f[��}�=x%�
�"���oX�X�"R�Vd�D��8š"������DU=V��Ѫ|o���ȓ�ٝ���k7�i��3s۷ُ�zB8BZ ��M�x����-�-;SM���ݣ��(h<�/L��95/G^>��w��!I5��EG�f��j$����3tܽ8�`�/�q�S��k"�W�tI��v1���s����;��>�w^����U�*�E���i,���b�{r��N.�M�O��+$�Tq9� t�k8[�s�^wp��ݍ�.b_JղwhPGv��!�ruU>:v7&�C�R�.�n�	�a{��u�.�沈�르K:�M���~�!��[j�BÁKɕn�u���2>��������~|2��V�䝸��k�*f�.<|7��ډ"�T�+����s����8�tٴudҷ�$弓%��l����At�bR�f�A^��7>xIblىм�s�fX�;�0���	��xkU�\�:���y���L_5X�I#��4��t1�w��UT�wq0�b���e�#�[��_���r�vظC̽}:�@�9OћIܸY�c �GNSٲ�_z)����4v������m_�}�+*�^2��ǉ��6�l\~TH��g��緵�F��P�TD�P�Ŗ%u��U�͘�c�E׹煦��_�|����� &�ᖴ���[M�
O3z�>�}�DR/����|D��%tከrE�k����yX�GF%#��o���-8,���+V�̴*��Q����p���Z�퐟��U�� �����)�Vt���
\є�Čp�Kg���Yl�A-�;��-#o��T�P�12�)1�U��%e߾���Oc徽Ց����0�����H��2�dr���S[��GMHE8hRB���U�Z�4X�e+ ���6�Q,�����{�����e�雵ҭ2竵�+-�lt�u0A�k���ec�۴�f�2��LsM�W���a-&�0Ji�!w������i��"�5�Dw!�7�U��S
P4��f�-m͈�,̤�y�V��ۆ���oˠ�G�S�3��N�������fpWW,$�H������'�'���!&�u4^	z`��+%gB�«w߷,XkP��j���]}���$���X��E%��ʹڽ����pVD�˩��?}�U��rz.�+Z��+���_��p��@]�=�v�4��O!w���z�%����N)�2���{��2�BC��K�����{��ZP�-��dQ+��-h��؜�� Ln�R^^
?��[>�x���:�K�Y�k�����ZY-��$0u- "�AϽw�	z�uZ�-_SK����j�&}��6�ʪ�JZR\#H��D��0�D�klvn�p�_����g��K�����ΐY^H��P��w��|��S>��J�¡H�-�H����� �<b*_��R�o�7�M������3�^���K��&���]�C7��\h�+/�o'�̸���&�t�����8��[��άh�X%HG��N�@���d��K���>CG�K�7 ���x1�X%��(H�I�c��"wX�L�"τ�I�n���j�-8O*U�_�b/n�#G�GC���S������xU�F�B˿�w�q8٣���a�ߩ.{�꿑��
U3SJ�B�SN��YX���7��@��� ��0�a��J廮����ٸ=н��.��R�2�Jn���4 �쫤m��b�1ȱ�2�"�I��ԙ�9��dQ�a�lӼ�q\-kl�[ͥ���`^�{�k�zo�k�0,�4�9~�D=��W'�}][�ns1�ÿ6��:Y.{���=�}~ƌl����h��+(�e�����E���Wi��:|��:2E�,�')L���_�j{ʹ��o|T�sl���lAM�em�E�M� ���V.mw�2�3BDtv��>�s��@�H�(�H��(%��e�����X}�1���~���'\��4���oG�&Ո��N��1�4����p�`kRG«|�6�C�o�9��i�@�45�]�
Q��j�|�U�
�B������s����X2/3ڭP�{,�K�])��/S��=�E}���gE��,d�iId_jB������q��B1qE#����#�A92nfy����G�*�߹[�0R-"�"J#���+)�婏����R �:�D)4�%�W��W��kF*"ǶJ�aX��/?�������#-�h���������"�J�j��'8�Ҫcd�*ic֑ƙ�j�E2 �[K��w���}���je�m{��H����&=�;�����w�J�~|�H
��ji�Sh�܉����NH/��Y�f�8�HQm�9B�{����ʣ�i3��BVC������n~��_�o)��~����,9i�}��2*���f�D����Q_S���u1�y�u���!m�ؖ�B��Yoϟ~��!�ha66vݨ���UqΓ����@��n}���\q՛Og��v�(�����rx&���q�1�'&M�s�$�kZ6�Q�3j�4��jQd�&��x��Fj�e��&:�(�h�S���k7T��!u���ŋ\�blu�̀�B,"ʛ!�`��xU{�k slmVqt�j'��K��G!�k�G.p�<���ٶ\�6���en��\�GG,R��^�n^acG���cs=v��8qێ���ōt��L�w�����`��B��|����$*�˵������H�H��Qtя���}���U0T@*"E(�i�������}��Vx��������b������x�� 2<�~L�C'��I%��&"�)��X`�*����(c8?3���
�0�~����z�>����`��͝Gϝ綖�H�,�D�Ih�,���.���WH`h��(K��6�7�s���>�����gm�p��>�'����qd�4�߾,��v�D�"��X�Ul.k\<*�D�,R�%�?��uZL��TY�\"�����z��ō//��u�D�<o׬�!U��}dj��P���kceY��#m��;"�LA9�z�,�|i�Q�m��+�3}��<@�_�ߌ��`24�i6�<pל��^ʒ����<�&<�ֽ��!|}�����^�D<E=�������V,,X�aYBɬ�6�
N
>�{j��}�![K��^e�g���Rߌ�z��7�m6=��Uݏ�Fa�֕�L��/_NzIr��S�&��A4�o`)!-�J�(�7��ߦGuh���7�둎�K{k���ȯgw+���«q�j�³����i}�޴�Ԋ��2�ĸw���,_־����ۑ.�)Jwӛv�w�����ȧ~R+�_��O���e錤�K�R�U����z�Od7M+���71Lnfi�UU�t�J�v��b�L��y�s*�f�$/��,��5��mo��������X*U�y��qZ]�]��>�V����36�!�)�� �߽.��?��.��l4��a��N�yH?*(�eEUT�jA�p1X�g�`%\|��X�#��G�w���o��~�K�(��v����Y~��QC+Un�g%,*�YZ܄��nE���LlW��3�]Gp-�M	����+���j�\kG��(��P𥉉`F9��~��39+��	$ٹM�N�b����Z�m6E2z�!�=�Q�C�mJ��~ma�{�N���g���,��R+#��]m�y�������Dw�V%�c L�t ��w�}�����z��@�������DV󞬅7�ZV��Wks�}�ܝ�~���5��ڕ��i�C�?]*!Q E{Ֆ	�q�#����$���s�_k�s�UH)*��\_�*<E�9$DqU5��=�fҾ���:w7�e��T���R�'�1DV}�Uƀ�p㮥*�S�Q'~ۨ��N '�H�SLY�o'�l�����K�ﺮ0Ŕ�p��J
i�����R(�:hc�����Nm�6Ԣ9Nz�R-¿s=W� ��G��b��b��ێ���AYz�;�wVzWÁ�SXL]���8~
+h�N<��_���ɶ��2ԑD)_}��_u�p����	p�K�+�ܞW�XM�}�d����m�)�]62a@YvJ��sv����c5vc�,�jb�+��cfTI�4"�&f���}�R��
��M7l#�~_/�*l֏'wH��B|q�{�V���"TG�%4xL�͘�3}��dӃ�e�ݒH���X%�+��d�;|��[Y�'	�p�2T�H�����iX��>t�x}C��U��}](X��!����k�p}}�sky����,�oe&Xψj��ebA����+}Bc��o�U��gz�&�FSH�D'�{-pCzB�}���6��.���
�$1�mg�	���)�L	���U�ΚxZ#��rF
Jy^�Vt\ 'O��:���m�(Es}��:��ȉl�*�����1?~�̆h��b)d��ё�"��K'.�j��ζ�ڛ��Ad+j�T���m]�݆�����-�gAv� hg�&���Ⴋ�b��ה��p��� �gݾ��˿��h_#�k V-8QeK�����<��f���6�z�������=WuY����ٸ���D�D��e�ұ�欟U�BZB�I�6%E����=�Y�7�z�h-�.���f��|���Z��W������j�����I��g�������)��9K��Ũ��3����	#I�&Z�=�j�`{�tAd*�sdb0SK}ϻM�5�+��UͻW�w�D��?�����`�>"�ϹV��"�e��+o) �������Y�t�.��1��&�\	t�_~}���^��D�K䑌��p�\4X�pW5]e\�� �j�ll#kt�ؑ�"�b����!��5K�
�C�|*G���^q�	�0m>8Λ�.4\>t��7�^�daC\t$G�W��'J������\�ޭӃ�w�_�������������)��#��9�Dv� mi�(�W��Z�*f�8�����ã�����U�$��Y��o��i񬿫9��V�%�<�f{�Dﷳh\H��'�V4�*��z��0����f���͢0d1��{>��@
$c+��<��p�r�� �"u�Yb���=<)��L�sUkы�(�[LG��$޿s���:\��
|�@E�*m[��� x����h����E�;�ň@t��߹���_�(��о4�B��mZ�t+�@����L&���9^�&���mԶ�����O�#���w%u�3��yj�5�d��g&.�8t7�I�jJ����ﺭ.��|@i�ꕂXa7r����ZE�8�N`J�!��߽��K���E�Wr*�����|z��U�������p'���	v�gX�]ڴ0OL���v����~�����Y��P��,#���6L�Ew�k�ZݗST�z���5�ő�}�DE���=�u^ 8�v*4�P�8`�yO�z]����o�}��82�TB�l)rb��z��1����n�{J���!�)��V�Lb�ܩ��Ϫ�����z�I>U_x$2B)��ջ$���E�6�HcX��1#���X�0��V�k(,��l��̱�?I��DK�Y"����N/��U�#O�����HR'�|���y���ե�|v�J���7�v���d|xRy�߯��-9+����F.��ߛ�mICB�ߵZ�a�5 *w4)������5M�$�eL�d|a�>�h����(�1t�_r���p!��|�x�ׄ�Rġ��
,��
��9~�+��3��B�P�<�g
`��;�@m��4�\��$�V���D"��]5�*�yuW�W�hv(Ɗ bD~"��-�p𣠵	�م����|�@b�VE���-8{�w��#�O���q��iM �s`��ۢ����/w�ˏq��P�8�P��J{�K��p�C!�B���r�\p�)��bbr�(Y����o�n(�`����#N�b�:'�Ƣ�w���|�w� �L/�V���~ҏ��+!{.b����Þ�b^�<)?>D�A���R����Z�w7Y�Gkg���Y�@R�ݤu~��/�Q�=��Z�|��,N���jȐ,����:�|�SP7UUK�oX9(�D��$�1g_6���g�����%�,ڸ�c��w�g-Z:�/��v����'|�VX�d�ϥV� Z)#�����G;3"�d
ɖ�	��Q_ǽ�kq�_��JT ��ʳD��������?Cw�f+���,��^Wie����
e������}j��k��Sb61���qՋġc�j�F��,��=_�*�T�C�m΂��v��t�W{vnL��S�v��"Վu���>�l �����,˗q��`�wkV݅�$�z,��ys��{�'u��:\���B��4��Ńx�=��,�7X�D�٤�l��]hk�w$?�<�Xf`�*��
%�0�Z]iSU�.���v��kv8�f��jB�iK��tʻr0+�΀�AF�*�� ��z{F{uN-���b�$+���0U��/,�b޶�Ƭ�.��1U�����y&���8d��+�
�g�NF	�^�YG2bEB�t!�ޜY�I�ND
�k�r�1�����is����/�<'���B��}�kٵJAK���V1�+��z�zv_��t�N��S���.�]0e� 
>D�B�u�߽|V��_�}���{d�|�ç��us��bV�h=�W�
����O*n�� �MU1�L߽V�h�&|�
�nI��dp������և�vXg��=��<F��:��#6�X���������$a(�ϼSZq~���5��ٟ��rcZ-m߻�q�l�qBL�h�.��T�0�e]� ���wb��=�';�6����1����9f��bE�~���x�+g��s�W�-\p����"�]�O�TZJH��"pS a��QB�B.����"��w�H�X~�Y?tޒ�~'�^�����e�ɋ��	��a��}X�?J�QF�V!
����eH���+V	#�yktaIY2��o��j���X�N/�3��5��%	�aO����2�IS5X�CD�N[�����z�o �T&C�	�o�;��Env
�2G~��$�?_欳�I��+\8p D����A-0FB��ג�q�Jot��#�;�r%zؕ	�;���b�ٿ��|9Oe��sYF�#4��S��P �\��bi3K����H�U���c�֥�3X��MWR��`�B���_>N����4('���(���x�G�J��o8�x\��+$^���lL)�wbgN+�5u0�����^��գ^�l���a<�z��8Y����`�)V�W�M���D���MR�#_���ŖH(b�8��Qv~�������*6��BZ/�o��*Tl���"�I�������GӇ/�����!x�n^cVҽ�c�a�*�S��wzwa��w�~k������J�~�5Sm~-�[TiQuJW���V%���
�S*I>K*�@-���έV��[.��r��}S_^z��H���;�у�8�d?�Oj�*UCMM,f�G��Xa_vhDG�*�}��Ѥ�1Yb��y�|��<qy�굇�}�On���#=r����]���o��#@�`#���xC���b�(��G5k�qEs��/�GN���X�/X������^��H*����dh��#��-o�H�9�����H���{�J�.�P�����\�[�d�X�?$� �_E��|h��w¬�2�����qC���#ZB�����<�;V�G�e����tU7)�īxu�M�6�Q�ԉ7'��ǈ�SZ�:IDX�竊��`�̠��R�(��P�D4q�y9���]��D=7��Y��<$�|Պȳ�]щľs�q�x���m�.��`��i^��_Ś.	�s+n5]J�d_��v����u?]Oec�zZ�����3V2�j�3Lܗ:�Y��5YY��u��͹�f{ &�:��<��� ��RQ����[�!���e�����KG��zZ�'��F��vʮ�X��U����򜅌��e{�U��۞9�*��i�vl�
��a�b�����W��f+����?a����Z|����h�"`T��X.�L�GN�O����>׵?�W�I�ǵ�����C�a��� ��^�u��|�j�l�LpVB�$�r��R��e��:s~�F��!�3��7�R��Gԫ��Z:N~�����@��E�4wt��K�U#�:USU�-8o�у���D���{���hq�F@]N��e���2�{��g��Z����$�Sg�
�V~�.��Ua���s�jȯ*o�|�A�yac�z2	��M�M�a@���W��w�T��AB��p��\�J�?/9N��mi3�|G�����W��|}�Ǆ��DO/��ch�m8n$��G%�,�C�?i�ih[��xv{�0�c>��w�:���@e�hM@�j���~���/�l��xS�Z��iY'H��ݫ�~�ӕB^=O�x��/w˒�n���`��z�YƗ��V��׬���鍏��Ҳ䉤)!3�p ���>��U��\���&f|��A��}���~^�v5�;WWY����Ɇ'm)$丑����֮�9Ӥ�YP�lEs�"�k���y�+$Y�4E�8\��q�#�n��I�]�?z7��c�Cv:��� �8�ܝ�"�\ۍ�\)ngx�4����q,]p�n��e�NisE�|&�r|Cǽ>� ָ/7���\a�*,VF4ن���������Z�vV[c5��	I�P���dw9kV']����}�>���������R����Vw�V��Ӗ�7���]߷�oW1���K�����3%�E	Q��[K���~����{�����Ø62��PKTI�jN{��lK�j�ipӤ�k�2a`/�$���+��� o�����0�{~�Z�]8[}���պyb͎
EI[�*�h���u5-��UH�4@�.�ڣH�x�V$�{��!i�@E�7k�%��C�d�߼/���̈S��3������ �<�?'�d��ۙ�jE�uo�HU���q�I"{甓/�0���F�|Щ T�J�]U��+�Bݑ#=�ky��7^���5�$�8{����Rǽ�U��~N*���d+��\>�i��q�&��^{ݫK+��֑��T��߻�y�<����)"�Gv-�§��Ø�6��'�.PC�Y�k>˙�I͇��'��N`"&R���`z�����y�Վ�)G�N5A-�&{��Z�B�4�����2d)2�D�-�/�����
)(A���s��V%Ӄ9�*���u�����Z	�|��Јϣ�](<~���E4��٪�h���x��X��Z�n���Yt|q�]S��YN6�P,>����{%��߁�� M]1j���rBh\eUS,ʛJB�i��0�e,�s	�t%͊��gj��Y�����j�D��iQb�;���Z. �1La	�VԋE� ���� ��ň#���Z s����Gi��F���z�1+���/�2���l(���H�PKwjֿ�iB���B]Ƭ�kH�O�=��Gj[�4椪���8'�Ď[���5�bF��_���
�_.�R�`%�j�Lʲ95UR)�X}�{U�8�Q{Ӧ�\"}��Z��|D�*�G�)U<%�u�V-mj$I����lѥ:��V�0�Ţ��{�~�G����Y뷽>^-����V�=i���}��8�rҒ�]��*0��/��������1�DP���~6�xwF��p�L:c�뫌Eo���Q|tb�`3����:��αvW�I�9}d_����}g�|�?���}>TJ-�ܸg��qx����b�\�_��.9�Ă8���)�>ʾ�֤�2�t��ՙ/=Y4�1����D||h�Va(�K�ǀ�>��,Y-c����.d�C*�:��j���|��*��V�Q�R��<ɉ�Yu*��{��7:�Jr���SUp�]z� ��zң������gE&	�i` �"o8ϣx�_c��x��&��n2�,�M�K�{֮:o<H,,�EB�}YJ�ڼ6[A��ß�\��˻Ő[�^���ջj��F@�s^Ƞ9b�	��
�oV���ԙb�K���_�N���s�8H+M\���חV��aZx`�mj㺑Γ�tK�Z.�A�S֌"��Y�)�N֤n��v�(�/��Vi����5��ů�:���fa� +��oq��V5�u�IN7FkR�u��	�m]L�9�]N�Va$��NR�\1�T�z(h��a0L�!N��-2!ٔ'w-�2>C��m�/Z�nnɸ�O�*�3S,���0v��jQ"1���u�x���O��ꖢ�P������F1\�;;MB�j"ڶ�=/�J��C
��z�svj��A.ӭ;���,���z����o�C��6���}=���RZH���sm�J�!�K�W�s�V`��c�K�r���.����mv^*n���y>3pl��n���F��y̻t�B����]�0���ؽs�}E]�W���vX�`�O2bܺ'7�A����t�ޭ�-����w�����b�m��'���P\
r�o���W���wd�{RA�� ��˼ɭ\\�Ց��)��E3~+%N�Υ�oj�Y�z+�\�! �y�h���S
���	ҙ��P\*�����i˻�r�keJt{��{0$p�{\U�+�F
��=�v�[�\2��8�V��17F�.��^�*?��>z��e�EBW��9��XN��W���jօ�Z���㝼����rxNÍ�Q�#�v��3*AL�m�.3��y6���s�yN��� ��.�73KX�V;K�f�v"K6!���=�xだ��;P���ta:��������g;M�q2�{t�\&�0s^b��R�Լ.����szͰ�j�pť2�=[5a�C7(�ˮ�lY�Z�\�'r���:��θ�4��9�8�4ltt+%i"�㧓�qt�/*E�y�78��K�V1��A�5�@�Fcc5�Y�kE��e�j�Dv�(ۮpq�h:�sIˁ�j��1�絣�^�Yp\�@t�YFi������c�啘��3���T�7���X�dJ��qPm�-��	�q�%�Ll(rbH��u����1��.C���/*ڞ�s�6�u0<z���]�h�ݐڵ��{pc�����nް7XS�B�vn�ݗ�P��7.�����!5ѕ�9-�4�s+ilu��u+��(�Ax�:��-��x���x���\�*�$Q��� �.-Ҷ5�4\ή��sl�c�|s`vf1����08봹���C�1)u:bS3��k,m�8� ���p�.���Ҹ&�2��(�L���{qg.{��X�t(�f�@�k��[5����<� ^s��m�3�lvw7+����(r�qigk=3�9�Ύ5�$��m�m��������N����r�;q������F��;>^��I���c�Ґ5]�u�qM)�Ԩ���>�۔:{v��;����+��<�7����Ӛ� �@� �Z���� m���-q������ti*�[rV�"�6�I��ډ@���V���#j����`V3Z6av�7R�#uD���GVj����-�٘-Z����;ie�[=B��%��D��m�H��BX�\�{<�9��^ή�g;�s��q���Rn�K� a��":���.������q��{r��]���p�O[��ޞ��[gd�L�s
�Zݺ��R�=���	꜎��:������N�F���hڮD]�Uqu�g̊V���m0=����e�ګ.ګicV!Z�b�l��7Vl��aȯ�������l��ܗG6��Ϸ!՟�����3sƇS�&ܫZ���&��֮�<�z+�ΣWl���1��@V�ܧ9tͲ2��"���jR���ے=6ޕu�],c2��ܦY�uءm�\�r�v���
�Z�����K�2ف�U�׀�[n ��KĀ�[ų�n������kW�ٹ֢����Tx)��-�������U
5�vɝ���E�Ϗ�-�:ڇ��~�v��=g�͵��=�����Y�y^��3d2�þ�������1@���:�Q�wX�G�!�P>�}���z��ν%���ذ�T����n�`�s!��앍�B=w��!�O)Fpy�^bğ4���@�9PCʕ7zUx�����������?,�Y�LR�	���
Yu��N3af���(�]����S[��P�I�6�B ��H3-�s�o˳}�e�q��iS�!�>�+�Mj;B�g���d�ۤ?b	K;ۿq}qs�*�5�6�IT�$�!�IH٩��iV��en��C��d���T�����3��luΝR���B�i_ot��ʨz���q��:+��4e�rZF���E�דj6^)m!u�����nhW�u53��S]�1F��@��:=�t:Wa��xp�T�����X����s{*�Wwe��8^�
�W=x�{v��`w)�I��3")��
 �8[rc	o_J�h>�B�fE�~�e�ՆsI�)U-���a�B�=����(�׷� �wGo�ԁ�H~�uխhɉ�IL�q�3��e,G�8�AX��my)^�f��N��;ט.�Uxގ��UTy�t���c���t�&��>��T�������Wt��}V�$���T�9�)��m!��u>��z��Hȸ��Qb�U4Gy�c�I�a���%��nD=�"�_�GsO���Z�Dn�^�B�<b:���Pn�nƎۻ���Rƶv,=��S���d��mT۹��O����\j`Q��i��BJP�$���ÚLvC��zg�p�q׋g:�������l�&�׋��|�REV����`g�{��Wƒ����R&��V��%u[�C6��^T�v+;;ͥ�pg�-(�s�A;�oln�l)�n���0�}nj�[��#R�z��Sd��C(zz�<[�����r�|�M^�g�	���h�)r��F �����җ��~�^�v������:	�_&Y7��!R3>��_Ki����<�du���{���5���`v����=\M�|>c[]W�^K0-�)Q���w�W-�.�d���t�6�;-FUU��<����{6��L���)��g�I��ǻv�.�V��>X���C9͈��I���}��~P�{��z\?xc�~�N�d5fvܵ�U ��PƓ�
M��h�qD2���~Yw/2掞��_]��>�O��RԹ��Sn����;�.�} �e�6�;��:Q:�(טq,��!��4���2AB�F��䘗�_t�U�r��1Z�5��-�-b]�.����4o�Ґw�y�,��hW�ַ����0��!��˅�dAteY��E�֢�v�X/+"af�ً�0��S��aF������c2,�V��+)0��l��L�P��I�t���,a��}Q5��w�p�{�&b	;4㻌��aKW!�E�)�,{g@�Ջ�\���/��&��ۡgR�'���vr�T:k��&pL�<0�]��x�MS;}�x����Y���Y-�fH��VVH���9Z���F�]0k��sF���ڙ��r��E/d�5K.�??\�0��d�fRF��g16�a^�ܰW���B����_�rG���F����%{ǋt@�}��������쮔����3�'����X&[�#���Yàj�G���ւk+�(o*v�]՚�B\]1%�M��Z��Զֳ}�^J�6J{�$���E���W������%�]
�q1B���c.��M�n!��?+ҽ��C�����|��f��#�"���*�o)�|w*��*�z@�ai8�f�(ms�I�n:�p��n���k�9{4�m�lΨ�� �-���8_>�Ɓ��fQ,ofC�m`IH�w��n�1P���{�>��J���z��nI���h���&l�����t�tJ�+!���1�B�)��#�����
�_r"���ԅY�c-^8o}ǔ��I����9�HQ�}�|r��U�G�t*G����șL���H=��S�����v�R�ҫb�~�m!O	��:o��cu��ު)�֒���;
s6�y��D���obo�}{����`p��� �0K"�wadJ��#$��c,t�y�s:};6�^Lxl�n�м�Jx�E�͏$��{��3�C����LV�}�������0x��������>�t�vEo��i�lA=��8�w �ձ��Q7o���P²1�ӣ�3�z.�s�{�l�}��g�s�:󇂀��ŏc��Q����׼���Մ���f��q���/%��<�R���w��\�����b���m�pFP�$�D�;�;qn�d1�s�q�ґus�>T:�Lum�`烍{���x���v����1צb%��4Mrb�!�e�q�!z�/�(m�T#�E����fP���������h����5���i���Й1�e�d��Ld������u��n�v�* U�5
āf���,�9�b[�]9S�{�r�h�r����\��k<[srGke�'n��B����\B۔{'":+P�R�ˆ�Ma��f��4Ѩ:bYq�fPF���ɋOOI�-V̾W�iU��9J��!'�{��k���q�˛!pN��]'�cs�2���޸�N6Ӭ"�fi�u�z��o4���	L�:�����I����g��8�'��>����֭��J�E�{���x�� ��O�$Ʊ��d���Yި[Ӽ�)~y��<5�}F���Q��������F�3��tin���6/��o��m��|�'���ׅY˺Q���C��xYB�8��wyT��ʞ��S�G�u������<1�CU�R�B�զ�u.:	fKR�κPP�%'2����IYrkr�o��F$Tևλ�Oo���V�;���B���U!��?{h{3/&��2y͂���~ڞēQ���W%?�#%ճ�a7a6,�"ۍ3��V�R�l%,u����ю�U�s���k%L8�u7�8�l�FҘ[y��>y �yj�/o��b	�7;����-�|&m3
���+�:#.�0���v^|7H�|�ˎ3��<�ה�Sܘ�J��$j��H��#k1݊sK�7]����&ʂ�-ז��˞�NK�ǲ0���M���@�˛��/=O���9�.�G�~%0���"�)7%g%��"am����,��l�邪�9}Dj�k��iJ��sȦ�Z�k��70��������F[0��|�g��Q���W�M���|'uJr��El��U��b[
���L���xQ�������ǵ�.F��e� ����p���'��B��j�;�(/tQ��M�Q�웵��*Y�)��!��J�&��^�<�iIh�������{��_8��lzuvm�e)bYf��C��'t��s�r�
-oaԚf]e0\���m7'<�m
����J��&U1y=ݺ!�<b\=�BEӺ�����ܯ��ub�o�aC5��V�W_W�dP2��I.��p}���̸*˕��������J.;}����e��u\��_-�w��c[k��}4tG��tB���&��DF_'$������|�/��Ց��0N�d/���A��+�{�vN������u��TT�a���0�w�����2���wn����B՜�J��뒉ב+�����������ȹ�s�@����~H(��$�nA���*��߸��ў��n+.L�U��׸B�k�3L�Fg�~ɱ�ٺ6yJ�R>���ㇶ�QL�66-�D(9;�}�8�v�>ϼ�%��]y��y�*�I��=B;]��^�p���q�ȇ�⻡Q�Rx����;v�M��:��>k|�]x�z;tt���`28�epK�	�f��\��k� � �p~��T4	}�`��7n�`1]�����%2�-��M�.p!Fn%~ݘ�zq: �i��o�z0P�����brO�RD�Ot��uB����'�fq����׹�؃+������C�r�h��rK�4���D�)��bU�;1#���(�ޞ���3���RF�1��}��Lrkw�C��W�
�L����lC�$�*N��$�l�̍�nK��=�VBTw�%ڶ����[�<�7�IyB,�>�����H��ݲ�^�����:(?Ss!;�B�������:��}�C|��Ӎ,uI��-W���s}y:Q�U�J�.��dA����݊���ر[]g�8B{��3��>&񋛔���I�u� ���`��r9=��H��s�^�y���/:�dU��^�)"��N4]���bU����q��ҙ>���]o
��S���Y�c
D��6��	����s�Ne�eHE���m�4�W,Z\���ޮ�TXh����V�7�u%��s�!^�b�j�~-�*Dz���T�b���z�0V6H��a���xWN�n��|�I^$�p&���-�	1εT���L����{�,��c����n�F��{��8���F�hM�x$��^
�U���`޾���U����B[���8����� ��B'+_L6Md���l�k��JkV'�Q��w�^ܼHY���I��.�UN:	5'���l�:�]v׫=|��qo����ԟ��c}վp�(�3��t���$�S��}�ќS1�j���Rwd�~u6�����{(]��cNbr5!Gd�2*�dk����A�E͡�̖p��(�5��z��_�))8Ó��,�m�*��G��ߒ]T�������y�$ƛէzP�݁Wk/o)�Z�v��@�o<u�TȺ�Y�5$t�޺ª���v��wi�ڈD�Ѯ\]m4ͭ]4]%�����(�n�������ɇ��v�B�2�|7iuX���d�shF-����,�WWM�m�:�q�C�j�u
��d�:�=��ν]3�;&��Wlk����q`j��YR�]�O`���5]\z<���RŅ���Y�F(7-�CAs�r.��.��p��z,�ѡ�e���hZ��kb���x �!��f),p�3�f��� J��\y��l���d6���GQW��g]�K��+իPȤ��j�&��b�{.�Q�iZ���;�肭3�`�#��
U��{`�ٛs@yR!/0���9=F��Ce3�f�:�DeЭ���.u��U�j�\�����=��-��~�G�0B���Y3�G�xy>�o�����'�y����iyT��%�?Osuu\�]�$���`u_`����L��ཱΖ/o���!���{jsٹ��Rt�kc�i�؈��RAV[��F��]G/;�;����%�/�[�~�����F��w�c�"<o��.�ge	R�tk�,Y̬fK��+�Ns@�rD�j% �y���58��q��z���OP��x罷��o�=�49��7���7�ë�8�N{�D�A)��1�q�mE�Bs�27u�%�����;Y�vV˴5m̰�]�۬xVhE�Xj*����ϰǟ�j�t�{�
�eg)�]�ʼi��x�\.h^�wi�����������.&D�)�܎�灃�8�v\�hv"P#��0�<�}ٕ�sYݛKJ���3�I��3me�z�L1�t�uD�}-f\:�j���T���m0V1�Ӈ.�hEx�0Y�J�Ny��ө�ȟ�3.�/�S'�w:�m⻪绊�e��s�g%�Yp/�f2؍�)f�Ae{���H��=n^��'˜ֲ\Z��η����}���-s@�.��G�9xA�:{�A�}ℍnA��H]�;��l�>Wb\!��^����y�6���XA���^̘y����b_D�z\*�`�m8�QFr��Z�ߦg[��z�|_D��|4�J��z�����J�I�2oxM��IUܟ{��+=q��Z�[$�7�'���� ���"�6�tj,��-��2Y-�և�n#nS&��ѽ'�D��H�z1�W`�o4Y��7P��ڐeq�	�y�Ƹ��*r򳖌b�W<m�d�mv�K�������$S!8���36�
�U��<�>�Cx}��yv|E��郚��+y�)"�6����G����x�0����>D�m6��H-�k!p�c���8okѣ
j�ó���S���Kk{���[�>�7A�$���*%�ʕ�g����?diP�ޗ�Z�Mؖ6
֪�f��1�mb�p��j����wݷz.�ScS=�
b�dÚrX�k
gF�jԵ,�m�N��]9ve�Rf�G�O��|�l��g4�cS#�Y�N���~��� �V��Q�4�s�h�sw�X;a��c�7n*V\;$k[�U�(����Y�g%}�-	k��]3.�JL#0sHnu+�eǶ����q�]l�x>�l�YBR�����6��-R��>g��h�0�Gw��x.�l3CZF&:�|֫�:j�N���k�ξ���{xy�����5,�͈9C6�xM�;�i�R�ʊư!Qs�m,�*��4f��u_���WAQh�LW
�2�;R�ݼ����4b�s���3E��>'�G�g�C��F�^�vnFu��Y`�,��C�eeg[z��b%���o��ss���L�bs�Z �[9�.���9�=�ȯa�[�xM�aN�)E���s���H �ѳc+FV=)����o�q�CN-թ�����6�B�50SzF�x��Ŝ(��5!�/Zw^fc�X�z�:��oz�$�Z1��t���[4N���8j�v��8�i��۝q���V:ѹ\{bƬ^KN���:Z0Kh�t�;�v\W�vc�'>J��Nl��ھۆH�C�����%����@�H�}V�p���/�-=�9���zy�=W&��A�?.�$,kOF؜s�5�6Աۧ/S]׸-&)m�}�+�Gd���7��T�\�Bn�*H��hw*Od�{����g�-����KN9�V�vl�FX��y�ç�&%`�w홃�dE��
�X�1y˂�d�<n�_[�9d�p�#�G$�5P��(��3eJ��;�ؠl��aJ�9��;��n����=<J�4���X�~�i8���?�m��6����E�M���:�f���]��3	�j3v�����,���L�me����@g��>��X�ǿ�?^�`��7>g`]���I�@���_ه5]/D�0�o��w���0U�Q*��n8�����"�^���|�9�U�s��R�x9��^���i̦�1��W��h�~�n�VS1���~�ξ���7��ѧ!�	�jG�_!`#��wt��#�QaumXԳ�sEu.�9Ӈ������+kn̩s����6vVr�6f��-�D�E$��=��^^wB��
�+{ةL����߲hagK�����v��.�QK��@�Ō�7�;r���ˬ����h�����~\�<ԄO�,)��ԯ}�}���Ժ8�g�-����Z7�.�:���玏W��x�n�݁&���#o	5�/Y�wq-�[��,�R�\8r�}�w��$*�V��}�c��X}jc��`;cň�o:����֮��!}A�2�R�)�J�f#1��d�KbB;��w,��h��ČJYt��{��] ����O�=��3\����[��6W�o������c��ms�U�����Ϸ�=ތ��gP����bQ���/���Ǉ$��!q�x�6�r��%���y[�7ëq��c3:��,y��rb�N*&ڴ����t�Y�^�����~o)�d�w�*��;�g�≵����9%��=������)C�Z�*	}}|h^���[��Ie���]��2�q���N�\�V�z�P/���27[���(�j���}%�ń7�>�oN��=��hT;��~H�[/�{hm��m>��Ym�]/��	rӑD�d% ��%8u)�N��y��ED��Ӑ_z���/�^����^p�2�m����9"p �ޔw/GU���o.E�EQ)�s({
~�}�w����˜�;*eV�Q����}�_I�Ѩm9EM�k�a�B�Ǚ�$CD�o��M���IV��%4�b_;Q�r�-u6�';vfh���{1��n��n�#�8^q�v��R��Z��ka��v��c.(q���dj�ѹ�.�n��������Ys��̱��˲��F� ^Yx�;��3w"��<q5m�[r9��f]��mU��0���@���@v������ry��`��nB�\,75���cG��"��k%qoְ�unl�Y��ˮF҃+AHV��h�WK�e�	�Z+��Q�S��]i5]/�%��Wt���X��[>����������s���=�v-/�+���I�J �29$��ч�8o/Z��t����Ȑ8�҂�����^,"��&�M-�.�D3zLV���Uxk?\����1�Z��HA�ݒr��"����V�W�_�9����8�exz����vBo5?R;,�'e@⦄wQ��}!�&����Ay��ֵ6�{Sc�Dh�S�y�O-ӏ�=�삙�@�ۘ#Q���;F_&/�z�%�@��"��Vd,B���2I���5�;9�°���z�זī3(j��D��t=�I:=|oΈ�~V�&��va��>�V[�0h�g�~�ˀGԭ��6�2"�x��]�f�)I=�8�]�<�&��� bK.Y���b-�kv�T w�_sP,���^�1�==��j�&[]����Ӿ/�w�҉ ۝l�K��7��~�b���[�0K(w�*T���^���g7�̸=75,e��C#k=�!��p�*Y�<����2p��Yk��7���*ͭR,�e�mA]�S�ιP갎��B�g��zs��NU>�e5���Z=i�n3U��q��JT|K%Vx�Vlu�"%� �:�{ɘǖ��
�~��OmU�/��{��z]�}�\��Q���)�_nwPƗ�r���L��6`JI
�&�٘B�F^^kKo�p���}[;vB�����T/�A���Phk�Nۛ���%DK������ټGb�wv�9����HȤ�ǘM���^�*&U�R��uFKn�����әk�����[w�.�D� �Y��ܪ&���*NP!1�4ꊚi�v�d�<d��4[p�o[P�Z�U\8f�6jw6P���%�1	}:�,Y�R5WJ�>���uZ�'A���bY����OQ���~󱗝���^Us�ẜ�T���o1؟'kj�:���w2"V���{κ�Mp�L�΋(�K�C$����~a���X+
�#È>3�(d�,����5XSGy\�X}��`T�ԥ���^,U��m���V�4OH��c��������m��EX�L���I/D�m��4�5m��ջۅKx�!v�����<A����R�y�΋�#]}.{9Ꙉ�;=n���R���t7���^R?ڣ8֎�d�©L4	��3�<��1u�{��2�����,|i�t�l��5��u�z�l�n/�p�!�!�yꯜ_2�;�B��[5�������I�L��O=(j����}��=���o�x�2�����Ju9�$ǝ�~�����0�p�����������gvI�)rJKE�2r��o� �����A��S��w���k�`�!Jѽ�K�1ߕ>��(j���D�)�n#O�RK��}���z�ncݹ'���a��r6���S����C-N��l�y�����z,��o{�����	9{ȓCB*0v4�%TN;ш��S��ZdkA��wb�G�D��>��-����>��y�*eW6��=rv0�-ȴU��|��"%��}G��v��O{�`��l֊vQ{�4�e�h��}����_{ʻ����}��Ff�)���g��خ�7��C|�6N5;�V���nf�Z+.�;Nm��<e�F��'�[hmu��Σ6�_B~��!�_itM���>ASMq)�Q$����}ݐg�s ݫ��w�{���o���+�y��꫞������bc#Dm�諺��m���{��"����q�edL7��8����]�l۝��z�TvkF�B��߹L%vR�V%�{�ہ�"��S���J\����q�r�O��0�>��~W¤�����O{(f�+M�P�\!�e��N=�U/&�=��3�!����.y����'��c%W�3|�iE�DP�6������s3�v�f�
�]�M(Z��m��dի2D��;�s�5ơ	�٨�HS�Pǋ�kj��o�qgk]���m?��uE6t����Wco��a%�>�Ĥ~E��أE���Z$I^I{��`���=�?o���sAOf�W��0U}<f��z���fk�S�z�n��I��䉸�'$�IW��eY��s�aFd����N:=�p��ә����.�G�bcq��R��+�qFS>RG���on���{�a^y�O�m���;��N�L8�%��r�v�V��̰��+d�hͣ���;u���5�
���BdL�l9��N�Y�ˣ:1vे�#lR��[��Mvc����,��Mi�a:��9і\DΆP����_d���X�w*�2�uӚܪm���s-.���v�i��fc[tD�ܻL؎�[���B]2Bi�g%�:N\nMģ�F�[0muk��XXQ��D˶�в�ZL�7k�4d�lEB�8���cv׭�y_���0���
��b�����P�.U��5Z���F8�4	�]l�7\F8Ѹ(���18v�qc6�B�f��S�?w�ޚ���I[]�c�E�?H�.�ka�r�;O��RTNm��v��+N	��"�ߦ����$�Ch��xĩk���Y'{sG��%�AQν�}�!�v).���J���ѕ�(?Z������m�i��%�!f��F�ѲMN���%�+��3H��\�I<�7��y�:����O�[�k������������D�q*�7>L��yd�P괥����7i�Ӣ�(��e�c<�1W]P�)���W�v�;�	�}{۬�D�^o��*�\	:���5f"&�b�n9�=ݶq V�C[[F=G��CN�����Rb��k'.��JzF�J�ėZoX���:j��k���,D����\u��sc��`@<�\����Bl���\��ٰ�=s�҃W7��۞~��
�����L*yи�s���-+��Zd���¸pB���R	8sq>{*��Z�d�Z� �	i�xM�ژq��F#CVk��I6W!·nsv[F�0��u�z���\�yN��5�J��I}�e͚.m�A])L����;�ie����̅_�uٯkj���q_n{ή�OG�]���q��9��������I2 )"���6n���������W?O{|m��s=]`�h^��f$GH���Ϫ��M��$�a�G��$�j���Y��G�Ԅ���-�*��c{UQ}�}�=�4h*�����Y~�8�&ɡ]2����}��V�X
.&X�ė�I��b[����<;���/T�v�y�����T�.�#�O�tީ�(D���o�k���]˭Z=h0r��)!1��e"�e�����`krU��muvݥ#o�m��0��rB�� �ܤ�b�̙���D#2���>8i=P-�|��(������}S�؝��\_��µ�����($�RJ��u	�u,��e�:��=�ԅ!>�}inY��b��.�Gy�u��=����"L�V��/r���B�|PƘ{$.B�Hӓ;t����*��2�_o.�wNX���=j>ӑ��v�j�v0Rƅ�������n�*�z�A�],�3�`�G;.�Y��L�k,��oI��ۤ�M�1��u���ha��:�[���˚�P��P�DA�I�����:�m�6��G�X�}�1-��D��g��"�]�>3Y�q�>�Ooѥ�+��2�_>�N�d�|mFcq2�I% �c|���'[��U>j�yu����BOa!Vx��7��]�\�Uα�;�YAu�V%���U#��޽}��]��0���Y�P� ����{`^ӵ�e�sdƜ"gY�n�\֜���m�<����6��w�TE\��v9n-�"���O*��� 0�4��g6M9��O�2�ʏ�+�>���]J�mE,�&����i������{�5��dJվ��O;@���0աdNly���͏<&�C���@��|�SJ�I
@�d$��ʐ, ���J�	�<Z���xf�E-��N�w�Y@?ϑ�����~+��՘�Y�JMF'�D�!� ��͡dwX>7��z�=��meDg{:'6M��l*���>���ν��'Z0*++����]&�#+6З-��d����M�CUi6ܫ�����YZ���Ú�,M�d�Ӭ��o:á{#�5��q.P}Bz9�&5*�$n���ǵ1��/�^���9��9��9�NX�6�їf��ktU��,Ƌ�g��72���N��)U�d����$�o<�H6Z�n�`���[�g8�`���r� �j��e�c��Q�:���c�q���J���7������]���ս7¯�4���v����
�a0x���~�V�&�ʌ=OCe�讲�gz	4�C���*{*���n�h������#[[4���r�S������hs��,	{k+��]wjw�p�Etȣ�D)����!zwOV1�\�H,��3}ڕƳ=GFҠ�ZW��ۛt����zĿ4�����X|Y�	-��̉C�n�U����_y�/q����jR9��(�ݏ�uٞ�;�׆0<�.j�yɿf9&�[�%�B	mzz�A-ht�&��6�uxdz T�����ziY`xB��(�^�=�t9�j�h�<�oM�t�_�Lн��_5��Qg�����O�����ꤢ)b�O%`$HS���\���9J�g�༬��^f�4�N���'��e��Ĺ�pD'���Eg����tV�c�6��N<R�ֺI��7�噙�k��+,�K��45����b�%2&o�?��k��琕�F$Z܅����o�<LX~�w[z�}�ci�moHm�6��yo8��s)��]�rQDl���/j�����T�/�y�/��&tvw3�r�Jp���e1I�j�O,g�)�J�,s�����TsW�q9q}C^�¹7DQ�u�i�x֤�*/n���Q;�|}^�`�I~�I�g�B��A��6E���E�m![G�ݻAc��Ev��77�T�V1��a���!�|�L���<y�ܳ��aޭ��j�NP'�u��̱JK���f����3:=���b��ɂ�c�߷f���^���I��F�	i��;Hr��v���F�����eT�\�/�[����_j��>���^m�1fh�]��N����'M��G,���7nЙӏVz[޼�!N�}��Z�u��n��ɗ��q��
��g*��۾�:�ۭ޲s�m]�m"�4iĕ�����w�Y��t�ɘ�i��w]���qHi�T���e��jE��=�a��6r_TGOr����ëjT��'ap��1��M��5��������Vڗ�V�:�Ƿ{�L8:�/����]!|��u]���UTt���T@@�e
�h��\��U,jF�f������)K��<!��^NM�p�V�.������r�xuM[u;<A����h����ۥ�n^�Vz��ݤ;i�n�ܽ���U�nt���m �Ue�
T��r���Y�.�B6�t�X=��26�n���c�Xe��L�4��������'�=��{s�hO7hqz�eyK�I\+�n���dƣckp'n<<q��Gbu�c��9:�5�o<<�I���fY��nLʹ6��x�G4���r�]�@�S���a����v:�1�rs�&ai�P
�u&9�$�F�MI�oh\�ѯH�.�ƪ�cB,,�V�=\ػOhp3�-Kh�i��M�z��K6��"� K��u[d��&�/7De��؆��0�t,c2��b�A�,Ҧ�*RU�f�aKj:kw2�2�l�bC{G�'ew-�{3�h�;�G&S��6K�y�x�v:�N�{q�GD��pn ����^�u�γ��@u��P�uKƓ$�Lwm�����U���uM�b�+�����ŷ!��V#�Q8+z�볛v]+`��F��[��I�^P�X�K�Y����-��/(��8�
SCh����=B�e��m����5>-G0v�\�;��Lf�6��E�lx�������t�L�����l�Բx�)�u�[���Ü��{B�zõx�G���ЩO��ڨ<g�vy�+܏X�`������ɞj�7Hp���ٶdf]���+0�Ʈ��z,�1r;�m\��v�O�+�r�W2��s�q��xG^zn�ݱh��Fr/Xs�@���;����7��=8;8y:�
R#ƭ2�l�#j�^6�v�3��x[YǙ���n:�W�uG2�ɦq��!-a��O���/���4��L�샫�A�R1�Q�Y�2eR��y0��]��7�F�덬�`3oN��{d��sʤ��ќW�8z��h��͵&��q�5��`땱#YӢ]mf*��V'5���mb䃹�"��!�q{v����8��۵�0gr!r�e�(޶�i J���wo[�H��W�duM[��C�t���Vj��8Ě�q�k�m���ÎI9w����wc\ޥ�ZْU̬К�Z�.f�ڰ��G]�J��K��,��� ���&�z�6^3��헑n�f��!k�t�.
�v��t�a6��E
�l<ð(�tB.� �i�]+��s�p���)C5Ȅ2� i2�?'$�Rȥ�*���{[�V�qS�튳��s[uv��[0���ƻ��i���]�a-��7N �4�WvD�_)$�h^u}�'�]o�krp��!�$=/~Y6���Z��er�P�'�_�u$`_t��e�m23�	S:�*�Ù�����g�&��x�T��2���w�)	�!^��]5$��׻�q@�2���Ϻ�j*����]��TB9R:8t��)�}�ގc}ܗ����	�w����f��`�k�}�-0U����Z�PR�ˎ��	��sh��؄(d2��{�Lɢ�C���ʂh���[�N0[>����g�7?j:��W�
yR�J^�C�5l%I�xkަFX�oQ¢���(<u��F*����,%��tc�\j��_X"x��f�rF�15�'{�L��j�r�r!s��>�G_����iӿyv� N��^�|�Q�A��6��G��Zy=)sY��P"LJHt؟s�]S}��+�a�����`�����ɟ`�ͼ��;\��h�ʻ�̮�l�uJp���4�l쥎�T���PzΔsU��6;����On|�X#_zSC^k�J�~��#ɟ�T�� Y ��B�1�qՍ&�i�5C{���߱�x��e{ǰɠ_T�ov�=�P���ް�]�y?t�4Hu"FV�W#I���eE!KR+���k�㪻�G��J�� �Z�e"�^�3��!{�����hYL�l碁���c�o2�&�E���I �W7@���䯍�كǈڌ�^���Wτ��Rew,��a7
�{����_Ԝ�u�G��>g)<���<�M�n�L�k��h��U�[�qmd��A�+�Wm�9��^�N261�[��9��f�z��)ΖE�L^��V�uA{��*����s�����}W�J̾S�b�~�wxM���Q"\�3��r�
�yD�^	{m ��4h��{*J�>�I���E�p׭��_~����9�/Θ�>�+�X���
�L��p��j�<��W�l&�8)"���%�{d���y�i���O�u�p���f�Wa{�k�Z��P�h:o;+V6Q�k������(%yCi8p�qs�2�'�ƇkC=�IN;�>���Z7��W���XQ&�S��)��Ni�0��E-��|�On��톖{R��0�W��cy�d��qO{ϗ��`�ם}����ۺ���{n�,������2閹u�d%��t����|c��W]�yf����e'd*]��C����`�Gy`Q��'e� �-K��sG�f؎E�N!�T5۴�)n,m+�M��B�I9��N8�v���[�P��^�4i�p��[�yߧ1��,�\���wjf���G���ŸdYɡN�Kl�0�J|��A�ɹ��,K��@�ѐx,��T�t���+��t)b!�yb�Sw�)Y��{>�w/wL�I���d����|�m�%�	�OP�WBh3}�$O��v�b�Cxf��&�;�wmxy)&[~a���o�����GʟsXy�ʄ��ܓ�Z�0;˘�\]���X�p��޺��׏]�u`�>z��#�˪��C�:1�0CpL��3pP�C,�5�ٔX)k�O�*��ғ���I�*��jYx���	���'p5��ჸnbvz<��z|����|��T����߯Py/*C;��M~�0[��U�An�:�����nM}!�^���6s�)9�Q��)=K��I70ģ!3$�+�S0T�`��)^6���:����gO&IrL��6�"����'��I���R���1|�)F^���;\b�M99��w��_mad�P���˷���{>x�H��y��͈l��3�U�Y�O]�;���w������W�Kv�'�z*���x�G�ظ�cʃ�ס���9��\-��m��M1�QI�0��Ju���h�3{;�?xf��.�Q����W_�[�"���ҝ�����dwR(���N@�'x�dK��OX�����n�^AV�׊�sǻ0\C5w��P4Z�Ҳ"��4eW�(�<�a�=T��<n���0��N;N1$�RH0���j��ة���߹���^����9ˤ�8r�<��{�/�^�w".�-���7�3�dC��K��e�\��;���@�˧��G#�Y)S�����&݆ק�*?:�X(C� �6^�[�_���6{�z�=��_��#��Bٖ�D� �L-uun�@���Wh��.G��u�ӰC`�^���.wQ�֍�k[��� ���oS��qS	��k����s�� CX���e%��c�M	z��z���<�9����>�}���HԳ��뭫,���H��F+"�k�8u�%ji`�E��^��+ӇX�R����'n�јQL̶R��13���X�x4��q�`d�b�>��˃���l���E��%&JͲĮ�ζ�~���`U�XAx�yeu���VК~�G����\������r&�m�ub0y�z%J���>D�\�E\�Y�r��rŌz�>���ݏY��ɂ��lA~{�x��F�i�tk�<ې6-�l�,]�]ޛ�Ñ9@�rG��,*,9U���=}&��E�u���U�cZ�Z���Q=j��㔥��/���c�,[�������z�~Td���q��۴o��LOmK��=ީ@��4��F{�{��̈�D3����*һ�c,<�6�ųI�R�$cp`�d�J���\ԕ�,�2�^o�׏���b��0��rv�oע���AШi6{�PbRXjZf���-|�Wi1S�����5�,�2� ��a�շl��U�)�g5yݖ�LEr�8��K
I���8���5��'ǭ���<���*���j��oc�����k���ѩ.,d8� �㏰��my�j��u�*�v�n��~X���;ZwmjD� ���N�e�9������kb��A]�\9<��G�͇�H�]\&˔��:k��i�u�B�yB��Au9ɐM5S��&�uGc_yf��i��z���S��P%��W��Ē�I�I�O�WK��}g'�������K�)B�K���Ӵ���DރMq��~�T��oL����Q��7�x��4�G�$p^��/[�4�Ԗ�K!g)gO�d͒����9އ��Y�ʬ^$5����-������r1LVxV?4�� ,'&2��g���_y�;��aB���gJ�y�l3�"/��Ͱs�Q+�61%�[y%e���Gg+��Ϟ��4�Q��r`�a����lE^kN|.½�<`��]E͒� �F6M��͸�ȍv�R���8�IO:��=� �o�x�w���5hZ�[�N@�lk�(W�S��PG$ᅆ[��/6z~����:���d��u�.֤f�'��ܶ*b~fwO	o�ꍇO���΁����4"!�!��Q��@���
3K�m�
�`�r}�)*N̺%�wJ�]+�r�pv�oA�����i�G���gf�oM&�C�
;��|:K�4�
WKWIn;�F�yY ��m����$�	��W0�%A/e��7^�~�+���Ge1�O��zk�`�_<��6���w��|��5!�xf�O�l6�ye:0�B�������T��qq��л�3r	�^���P�ӑ��P�$���fϟ�w:��l:˳��6kE��2C��6�Ώ���ĩ�k�T7Ѫ�s�~նs���Q	$!!�"I��mϚ��1���8{snkri�[43+fUt�-��m�"P�㇖���_����y�T�&������P-��"��h>���ە��[;6�wR���cѢ�b��H�\�Ee_�2��vȷ��lu���؏i"�죻�Ш���X֕���;�Ћ:_yp�����#B"gĖ��]<������i
qM�x8�OG=O8uH�Nܸ0o�0�2�U��E������@�3�#i9�J�e]f�*��h����n�9f��<�z�|���� �|s�t7}8�u�w*��-a�(5鍭����c@Ew2Y;�YkN`H��@q���m�j�3(���{G�y�X2������������e�Y1H�)�#��>hu�V�X��9�z�F�6m����{4w�e��8���U(�=Ѿ�n�b&0yy��<�<�YM&�>
"��X� �-h�#e:�܋Z�$�v��<��nvG����@�Q�=���g�>��*�H��-,��F�=�~��������^	�	�F�vY	F�$L�!��\.�{(��0RN|ٸ����t�m�QO����IP�rI�V�}�7����b��R�؋�7��yx���C[* 	��$�4�֓-w��������%,>���D<��~��<w��ͪ$���^<�������̦/���-�d�X����޳�r<az��c�
I�#������}�2��\�h�0����`�>�&M�dr�#$É(B�A���-��l����[�|S�v��e��\�l���J�憳��e���+�b���W�L�|�aN�=���Xv@�����d6,������l�}7�:�Z��D����ba����w)����:�Q*�w��_[R�7!�ׯ3�Y�]���I*Ů�ݳ�*�`� ��)���n�F+;�v�x�����5Se�)�q�F�]d����О�7c��9�g�t��d�.��;8�y\�۱�kXt��{K���ֹ^y�w@mmGM�9�I�U\b�CIc-��	��+�+��`ǣ
�.1�/1p\�Qs��-�ax]�n�M��4}�%��3���8�Ђ
՛l�[KîA"]�5JQ\��2�k6��Uɡ����F:���:)�	�j������U꫺�g��#�g��YR�\�S���#�934����kU���0�`V�W�VJMƣ��nJ�nqpw��H����xg��yۼ��{�B��;�6�~D�����"���ScM-����Fr� �R�!F�k���_`�QˏA��ҍw��b�K����{ޝ��e$�wAv�۔�|�n�Ɉb$)@��9`nb�onr�ﴏ;�*�A!���wAV8�官IuӔ���8�?J�� [��Ԥ�fX"�;�|�L�M	*I+�����]�/$�'���f�����"T��Fn	����b�6G7�R��T���֯UT	��]��C�[(�a�����#�mN��Kͥ�U��^e2��J+n˴٨5j�$��x��v`��NԐ�t�0�&WS<�5m�����[�'[�����V=I�.��^�A �-��%$G<�����t:ŧt�E/���7[~����4�Y������U�i�U�r�\��\�Ɣ�'�,�0�|غl�R�ԏ8|w/���
���2�n������Ol|{o��>�3�Y.�#�:��T�t����u�5E�S#v_u���',�$��ۮ6K�C�8���\�#&�i�x<H����t}�P�^u:�O::}��^��|��Ci�X��*�����?&�o���s�ꎲ��x��IѮ_�.�<��~��s�fC�m��Fn�CNͪ�C#�6�������� ���d�G��u��TQ��hP;�n���_x]�^N�'��]dp^b�(9{˂����8v��zݰ`;p����)I�h�`鋴��3b�#A��-����nm\��#�Y��g��r�Ei��t-r�i��]/_I,�2��ΰ�i�.0\%���}�Ń}�T��[ѵ��h�B_X+�	y�4h���F[/>s��G]��ݢa���;ƫ*s�vL�p���s{�0��=Y�#X��+X��U�@LD�`0��Rc'[��͕Ϫ��i¼:�0q'_^���{ch>Wb7J;nNWÌ�})����r�������7ٲ��dɇ��֬wSYc{&���a�|�G4�2��fڃ���l�pq��q�^]���8���ө�*j��Fp�s�HR�y��8+�-L���'��M�:�#�c��5>j̓�VF�k고:ػ�7nW��bk%�TI��{��՝(����h;�0���NV0�ҒsQ܉�]����鯴j�ǎ=M�藅թ�2�3�Zu���@�#��7}7������sM�]�¡ʭ �Ĵ�����᭦��Vx�1᷋h��K�j˙�g8�T�nv�l�X��*�eB��Rt�ĭ��VL˻�㧪Tѝb�oZ��k�Kna:0��I8��e>��uG{lmc�v���]��@}�����
̪Q��-J!-Ȫfu�&�Xq8+yVHm��wM묓;�/�Ǹb:m��s��^]
b�B�KB�L��vt����P�z��'}�{n��ڨ��p���_�@9\�r,P9tF�����.>�v��o�+�>�,m�d��ySh�њ����.���ռ4��=D��x�]��A_4`�ga�H�ja��u;���q���[ݲ�l?GoS��Vm�TJTBv;o��ۻ��	��_p2� 
�*�+ST\��q��ev=�}lY9��M[�5��ج�����0]Klu���1S�Z}Y�oe���!��=yެ�;"c�},|�	q��d^��j���u�6򜥒퉲�^���g�a�Fy����s��j�8gMy�s*�RwR&_Ÿ��{q?Q��:]o�S�-�=˽�&�j�=�
��y߳ز�J�h�Jە��n�y�3qu\�_�o�zl6���r~�jys��Ϟ$�_�X�Y`����3�|�^>wB���Vp�Q���=/#A�k_�ר�%Z/�pO�JDT�:��q�L5�涓6ه�F�Ey��Z&��eX�0[&BnA��볓�Kޒ�^�Х˕t�õ,�ޖ ۭ��Iz�]U;�2GOsl\��4�+�WrcF����Ū��e	���4y_a1�!�����F�����x�/�Yy������w�W_cv���S��b�悒��N2�P����c>���4��){K���-��<�i��{r���dwq4�H^zfe�N���*��ɬ�^U�"Z1�-��p��1���Ŝ�\x��X�y�r,�V�T��{�!�	�h-��~��{5	<hB��7�uԻu#�`�,�����O[(�E����"mF�rD��ys-��:��ת�����N*�^��k�߁�B-��k{̥��2AD���z�n���+�jP3��\њ�!p�,�ĚC�v�����U��]������챞��g�Ak��[M���f;]4e��������Zx��m���e��jX��9�p��9|���n�^*l�
���]�e\Dc�����탮z;�;��;Q�#谨 �P���P���
?�?&�x"<j��ng�o0u���
�����Bǒ9�(�J	;�1܆_C�^_��ں��0J����xHS�	�􄘢0���ȶ�m
��4��%�6�^��M�����ߏ�z7��땏��<�2�w]�epOo\-�P"I 46ߩЇt�B��Uu]�VM�op{�!�\��V<��;��c�R3���),m8��/ʳ��;<�������q���b{���4����#�!����֔V��sr�|-��w<���w#��o'�f����(��M�S�lV۾���w2=��j��ã-��;2�]�/F_l�e^.ډ3�L�0�Q�Rnܬl�=N2<i;N�Vʎ��	u����▊�z�MlK5l)���N��<��]��;;½cxlv�jLrpo.�7�������p,���:�x��#[�lgZ*(����=<�e�zG�;<�+���K�)�ޮQD�?>g_ccɚ�1�F���e-�涭m����yۗ�Fۛ�*�c�hz��qƳ30�z��S��G22�'X���/���ta���N�c.v�on��Vy���yJ\D͗��m2)[q��+�m��f�6�k��94e�1օ�����΄/�vFgj�A�똫����{�0����v�v��n�%�w��t���t�Hսꭜ`-��G#P���_t���=轵% G��r����
��tI}LV�K��7.����%�	7O3�/+�|�r��C��aBC⣁f]���꧞[����&��v1��x{�0sg�o{}��$�"�Sg��L�x��=iYL.-�L	��E9"V.��gW\�&�o(y��������6�Fti쯉��\�߹A�Քut��H/& 1��ݫ43�A�㄄Tp��*0c>(f{�S]h�������2ͬ����ng;�Z���m h���3Hgg�HjdX��Y�S����6�)ט��l�aL�ZՆ�0�ٔii�z���8��a��hj��˽���}��n99E���R'����5�RlTK��4�<��};9Es�i>BD����~,�;�Ul��Q��'��E��-;C(�Ś_��lD_r3�j,����Y�5�
u���.�"�m�B�K=z���-��q�N+ԟaҬ�7+�l\�v�3�7N�~��tM�:熲wp��g�=.�� �< o�*X���j�\�	%p�kN�~HZ�d��#�_W�u�a�	Y0��p��H:J��qw����,����X	|�)���$���S*�ﶍ�i�^��N��Gl���ð�܂��]T�r�Zu�`��pO�����4�r,�L@T,?qg�hHq��18j��$3{0n.�i��K��õNS���j�n�X�}PG�)ҽ���i�Z�P�w���?��J+�=�n�me�av[G��m�D���glsǑ(ћƷ9����hܝ�%���F�*Ax���k���s��7׹s��"+WQ��=�`��Kx?#�B�ջ囒�N���½���ci��8 P�Ɂ�p�݋%��.:��uGp
c���w�/�K���*_;�	�\W���k&lD���s5"��B�"%#
(N^�
�o���Ƶ��
@>��������npΘ.��������Jdv�og8#�u=@}DK�l�	�pɷF�#�D�|��4%�`ѕu�v_��.B[X]߲�h���B�8IԪ)%&č|\�R�)2����lhŅ���0u�]IX�*s;��s	�=o����A�f����$��*@L� �(����wJ*�y��˥�}���f�z����7z@�}\�"'_`�FǬQ����/KO����/af���e� ��]���,n#��-�ۇt����[��HL���d���k�PP:��IG��z���L�C�?<�o��Q8�^���7��/��e��m3�8y@P,��E�*���B��xq���(ܓT�{*R�!���{���+E���g1������K��$#jH��h��Z�k��F+T��]�}��.�������l�ȝ�lTG:��]���=���yS��1���[�VI��fx��V�v�i���C�����)����.�jQ`�V���7��R뾩�t\�%Eپ�A�gn�[�A�u��h<΍�CJ�w.�E;��<eR��F�ѽ�kse���x��c/E���ĥ�)Q��)$�g.m]\[��ڑ�6�t�o|sO��A̚,QEٿy�s#�������$I�ۖ����d������M4�Xān��V�^aq�����oNQ��xyq�ۤ�Њ�����MH:U�����~iW�Z����v�Q��tK����6��4���?H$E8D�.����<�J��+�>��ϑ-����7�����qP�J�Si�׾��/3:	�V�f�1o���ҳ���K'��MNkkՙ�w�����%@���rAz���:��t�!o�:*��i�Jn��{�=�|��:�շ@��b>Ӓs.�M���jt��%*��"�
֊ZѶ81ä���OZX<�����v�z6]l�gV}�c��k����	�vx����c-]�N!5Yg�3O��x�>U$ ��H'$RM�)�%��}^�*(��c��U��G۲�U�M��G�޻�6sZ����fh{=/H�h�6�
���H79���ݨ;�+����KI7w��W2�xU�ѻJ�8>ifN�kWo�-�jo30Z+a�c*��7��70�\�D���gr1Ŭu�&[p��;v��mG�A�n�c�-�M����j:��x�Cfw/����-Is`v�4��:T�l�nY�a}�9�=������6��vM�>rvȎ�:�3��.���U
��j��]l�5a�6۬��B�gX�j�vb����2�-�^z�{R1�7vq���
O<��n�2���f�H:��	���vƖ�;)�Z[��H�/n7.�Y_��|���-S�Du�"Ы����eO��W��Ѱ�V<�v"�r���s�'F���+q�o����h,��>�D�d��� �x3�UT��L�K�{��ܾ휞M����l�[��"�R�}�Ϩ�+������٦�Q�$���6���N��ׂ�'I��2,��7�<d�w����wmm�h���Ki,������i��Z�|V��?4��n�~en�۝m�_��
��;����A�T�>���_J����Tt��p��:��k�匡:�%�9�8�a�̅�#�R8�@��K�N;ꗦ��KE'}}^62\�[+�mN�-Zv������̪u����̨��np�l�d�����0k]sS�l�W�R&��a��n=����tY�8�$�RG�h�Vc�V�*���>� �m��Ž�𷲯Z�����d.�^J��a�8�$�^�K��e��0H/
A^�_o\��w֭mm	z�}r"����΅4�o�
���4�,����z�fG#Ŗ��&�Z\���;�GE�F�52*Qڔ������ʈ%{(_cԏ'��r���7�y�5�Lw�_�ѻX��t#��^X�D�$���wq>N��j�����9�^tr����[b��;s1�=yL�z9J�2�
�[ŷ�L/�~gO��>��^�ٛ.�1���Y���۪�ͮݛ�y"Sa�{��1��%���$��n�D���^r���{/w�^0��?�08F8�ٹ2��we1��K�֟��o�^�r�����⤅�#�Q�~ui��ǱV�Q����?	���JA�-[s�nK��d�K��9�.0�Y���3a��l�0���6щE����ϟs ��NDֹ8^<�Rg�����x�iճ5��+|��D����Z
�d)x���i�j$r*��i�QN����Q%��(�[�v�:�4߭]�������<�,�)f�m�>m���T|����pCq��I 7e�V9����Z��rT���j����Rg���ؖ
{�p���e��5��ں�Iޥ�ۋ4�(%,;նq���;qi�b��oI��sN�brBZ��P�j2okӽ�߮Kʖ�ol�K��+�e�^�<��CrBNiԔ8�r$Pw��weG��7���V����:,�֩��z���{�&/����]�/
{J+O|Q�%h��q�)�:F��*�w�%V�r���w|틈:i_eT���ž�w�ݢ�a���z�}.�y@a�*G�>��y,�GL�a5��b��N�M�N1���������n��A.�:����k����7���X3(�����[)�B"Wp��]:`�C��e��r�M ѹ=^Y�ׯ��O��_Cz̳e#��OI4��T3z9�Z�g���޳9]9m�l�����S2X���,���k�6���|2ab��0��s�?��=~���EØw�#M�w�e�Fl��^��v3Y�Q�3ܴy��Ko��ѧ�QP�$����
�����+sN���t���7$���(5ɭ̳�=ĕ���������`��ħ�1���tk���$f��{fk�f֘n�!��t����5�h��t�_[H���V:Ӛ�����l��^g��$��oZ���i$Uh,�� ��c��Yy+3煲�C��3�RG��S����I�j�lU��m�ޕ� xr��^��`�����"h���*��ܵϲ[�[)v���c�r#UF�Z�h��P7%��Y~{Y���(���/dn��y�^Ht�������c�=%��]�}����t%/U�t�$�v�2B�H��̾�-�Q��(���*����l���zk���~�>��fy+HKُ���}]��w�_�\o�?Z�n]����ޯ�r������e�Px,<�þ�4��,=o{�뼖`���{�qX¼�j#�Vz&v���W�r���9�٣�c��{Qws�\�^�E��m��m-�9v�֛���vK>��b����bǶ����>�_�*�&ߵG�ƾ��������e{$�	5ܱc�0�ӛ�_�^l�/f�/d�����M��U|�-w�[ͮ�mk��˛C<��X`Y�9mwu���<7��F%w*RJ}I;��{��xD<�H8�Za�z)�����iy�ku&�Q���o5Kܯ���X����
 �k4�:ht�wMâ��&l"����6�} ��զ�f%��i����yY��%����
��1�D��а#c��p��H���*(Ыv�u�.��V\��9�ї,M���ّS$�0���vQ�5�9xYokiۮ���]�|u�^�ky^K����E�8��
6�ZH�\��T����ŘU�Y�Sy�FM��hܕ�=N#�ÀϜu�U���MݵM�Jb����In.I��]�*�;�n�a�+/�JB:��T���[��{[���V9�R�����w�oi���d҃�!&wn�ܦ�&���'jh0�v���.�����nr�x�t9��,�N(�'`���ܠ���"�aP�}�0$^F$��Ms�[s.GW]�Z��2����,s�9��W�fT��RK@�8޵]�ܩ�J,ӳ�WSo_VYg#v ��h�2�8keٚ�D�2�:�X�z�C�/K2��0~1�R+y��XWLWGB;��ü=��m�P�&�[�r���`#90�6h�|�U�39|�}P�{�5��A<�����R7V5����+0Y2ݣ�\v2�	a�ʫ�6}{(��S������[�&�*�J�Z�(��fj3��u�aT�&�Q�Uv�v!V�d�Y�������;�r�O[�ޓ���Um\�9Q�Ŋ��jmj�S*�Ska�-U 'm,m�8�5M7��<��w\ƻs�G��/h�K�jw=�dwm�{��J鬚2Ť4.-��7
�p���ݞ�����#�U��-n�\�r���5H0j���n.��3�ڬcX-�!�Q{8J��1�LkZ!;�����H&�y:�ʓ�&D��c(�lVZ6�/Nۊ7Q���x��m��E��9(1�6�5�a�dݐ%����i�#��[]�,G =�4���<��Y�s�E�4�ȉ��v�Is;��g	���%��άTmt����1Ԕ�!X��'�4��<�̻�]�M��o�niƺN}n�d���,0�(��"č��0�P�;YR�n��wj92�ШE�Ǔ:d�m�N[V.E6g�2-��OlT�۬�C�����\����v���"�q��jC��f1���&��Ci���Al�u�[�B{Q��m��<|�Ҧw��ƚ;O\�nh��s��4Uҭ��7[(�MU��\,fٮ3�-�!�l�$TN��q���EG��n`�ڮ4ѱ���X�[fQ7k�Ba��1e���:V�{L�il�{ C։V���zm�ʓ�H6H��i�Z�%�.6�of�\�ch�Z�������eM<s���ez6�AW����v@��u�7a'n�y:����3��R|#�n�=q�֝Ǚ�=d���f�g{��Х�X�]1�o>'y��qA5ظ���M�5�6��kf���#-p�Gh�oh��Re��$ݥ�nTq��!�6��6Q�[��(�l5l�m�}�'+����{n�)�;^q���n����(���!b׭3O���.Ye��<e��y`iy�]0;u�t�hJU�ai�sq�Y��:_=��f^-�7[U'T�N�ܩs��;�5ө�Ԥ)(ư���,�a+�܉5W��{q�\����n��Z^&�p��Fe��pqm:�;AhN�%�`� ��2f ˥eq�[cV��ku �/i.����Z'sn�ù�����ہۀ:�3[P{rF���B��e�B��a�ɑ���].���A�\�p�j�;��K�9�ԖzwQc9CZ;g�e+�-�4��݂��`����I��m�R�'n��6�ƌ�6�DMEʹ��Zy�<w`��]>�Ґ���i�H�s��[���B,�|��-͢ٱs�1GV�-�נ1�3��*F�B�A�-��f(
)^R�2贼�u�!�e@Z�(B7C�܎�Se��Tg�o�K���:���$�J��ol��IWs����n"%����y�8wg�
4y^)�H�J$!3� Q��n�N��u��\���z��T�k$�����5�Q��:���t�ux��1�����,8f\�WaO�rE"��mCj9�m�F�g<�L�R�S�^'�V���|΍����	����cn�[W�e��(�����(I�� �O��.����Lo�G��8)Jۘ���o�E�)��k{=�ğ�xu�,�n�����?8��$n(�p(J	�i��ޒ<��>̵.I�l:�������n�׳{ٛҪX+��U�w�qm?�������o�{nRY�k(�M��
)7^6��S�]u��h��2h�k���t�a�ͭ5���&ҲX
>oo���5�������eqU.��ʢ�q"�M��m@��7H�SMÊu�ǵ��o�gW�a2���1�d
I4X��V��0�`�_��Y�-G}�j��Kx�/��7�Ir�TeJZ^F�^��X���ͮ�YDN�E]�`� f=un�0���?w���}�۲�A�t�kw��!*��Q0��Uݹ2�9����f�yy�^�,��,F�r(�28-y%��Au�)�����J%uN[��o�B��fߘ��:��ȱ��X������q�7tRB���D.JY�FaiH,%����%�����L�->���.�]>�K��+rA�]B���Vs��������z�te��O;�q �(�J���i�깗���3p\�1�5g�<ཾ)߼䁋��|�#{����^����.G\��
!#�f���W����FKR	W#,t \�U@!R�b[e!c���kl��0�K[�҃�4��6{ǟ?y��x���f6�yY�yל��YV{ׄzE|S͏0�ze�ztVFxBކS)��(�4l������3����^�U�;!0#��Δ���=��A}Q�)˩�����w��o�ތW`�Vp�@�Ǽ�V�vđ�"E ��j���-����4����;��>�
ځm��]���M���PSQ��P�8��P`݇�t�F8YW\E1��*=6�ae]���֘�i�x���i�mt{�>���D���f+��m:�7Br�,h�����eL�Gofӥ�=޵4��ne�]{=?��s��vq�7l<����g��)+����(�M3b��vW����ߟ��~�_�T]��"��V2֗ڙ�^��W���p6S��6�Ǎ-�X����ɻ��+�l�@P�S#RS)4Ԧ,8et���Ǎ�WP���Fn2Lѭ�etKm8=K���X�u�4Y�˹Jʼ���f~;N,�CY��G��Q*y�&K�Z�#EBX��Ir�S)���}0ʞ�+��~�Hc���>�����+��}�����}&�v��8���zڞ��9+��9���l8�M�N933+&�&w:{c����|Q�N)C�V���μ�W� ��E��n�~���~�뒞m��?O@ƃ\��\�w�r��eK.Hi�K�`�_�y�T�Ѯ�H�/-���W��KZ�#������<5.�YCo�U�'5�9��̄^Z�c+&N��e@�F^59	C;�f.���Wb:�wm����V�+��]3=�K�w�/�j7�`�'j2ҟ2���y����wƺb��v���=������৚)K�=�&�y����Q��7��t����g����Rz�L��3���i�en�-�d�"JCYID��n�If+.(U˖O䣆p�(�o"��NŢ�A)�����xd�F���yCrh�zf@}-��<�t��^�q�ڤ����D���]�!|d�Odd�P�:��`��]wzŷ@A~�4���f{�K������pņ��h��Hhg�H��A#MB�rL�-D��Ur��Ϩ�L�Ʊ�p:����
������F��;Z��:&��MX�����:1#�
Ü/6!AI	h��p\si�\j��)�z���٘����h��u��ϑ]ϕ���o��{�����W���oÖ��v��{;��D�A�$*H}~����i����ݕԮ���\�]��Ӆ��0c�݂��1��ܳ����B���9��.*݅��ّ�y�VN�'Ȱ����e�=�t����iM�Lk{�]��yk3w2�Y�;dF�|�sf�m�H�0}� �܀��6	���]�n�q�u��,'���a�b�G�pڳt'��.��;p9-����ų`�+�=Z�e�����\�f�����m��ʪ]1�!�e�a���m�����SS��.�	����dl�Zs|�b�qՃ���^.�gkY`��%Ý� ��_|c�T������+mB���Ky��]���m9<>��D������<�ƍ�W	v�v��9��Y�]�F����kv���L]�[0j��+�-AG��g�m����O�?�Ǉ"�x�`'y��K�n���W����>���4�"�: �oS�0������P;�ֲ�,·�Ƹ�\�wZ�KT�4���G�^�v�D�'����N�f1)�Q{@u�o�?^X�\H�P8��mcC���.��M#����o�t�1�Y�*����^��_UP4n��y��̱�s(d�F�O�M��$J�ں{��4��}��+��OK����TV���^���K�|OUY�/{VTsz���W���&`I���Le��=g�vW�W�,�}N��\�/ԙw�cܭB�v��u�z��=O�&u������o0��������P��m�ln]qn��4b鬸�9e&k�X�g"a/�{ߤWE���c����m����]�竳%e�X_kY�lt�{��r���$��z7�ZPT6� `����h���uGj]�0��]vQ�+L�W�k����m�Sn�sv����wʍ�7�jч9vf!�q\ۻbX�Ml�6h��ş`ՍlJg���Q�d���N^ټp1�	���~���H��3l�o6�o�D��	�)�M�h	ra�ϒ�g A@`P���E!�Z����U�'x�Yq�%��sV�yܷ�]	���J7l$�秐�ؠ=l�`�レ���ÈsL>J��R4L�Y�"C�[w�BԖ�t�N�HMy[ـ��f�t�B+������3���Ǟ\����{�u��5��!ؘQ\W��0K�)!.{޵j;�B@?Jx;p4񽲛�zǸ�m{mb�Ǧ_���I�^��_�ꠃPY���iw�y������^�����n.Z=̑-0J/�,�0���(6�)3�6�;N�9������9^���Fc�䃸����^����S�Z�����<��\dtu��b~��˽";���T��]���ξ\|CۉFR8W���a���j����Gz-LWU1�[�&�%ݨ�޷c�%+W�.��m-��M�XJ��P��j	U��t"DII����f�e���^��ٵ�i �g�}鲂���G�QOBNS�,y�<e��5}YtMdt�5K��"��s��ۨ[�!]zy)I���?wQO���j�Dfm���s�c�"�~������b� �����6t�ԤPþ���K�јTPO��8��B�άj�w>C��Q�W���+˻���=ްhvq��>^*��ye ��Uu1y��/�����'���r?w�~���� ����N�J��evrX��唀������O^��ڦ(�W����]�$wu�r�m�C
�f��h܎:�u��sl��gU�B:e�P��$�8�5�@�W���!�ҲҺYs^J��RV�gȁ�\���UM����9�����ĕ[uG������=��yB�x*rAq��YfŹksfOW�Eb�fʴ��[�(����~���Z=��9�;�#�=�T��P�*�Ow�j 4$�uW_�<��ڕ���o��ӡ��	:<�����4���.G��[�K��6�r�v����t�#Жf��ܚ�!l��њ����)�"B2�-	RAy�� ����zsSЇ�8��*���tQD���q�#�w�e�Mxu�=�z�2�g�5��S�6��-�k���ݼ���Q���}J�l�h���#\j5���:Z�e1C��Gzm6쩜뾡��@n�`�H���K)��w��B�4ف�ʒA����3����z(@��U��ۏ���.��w����P�\�2w�^� ��wD`+Gq�o����+(���D	�$���ͷi�fby�v�6G���e#3���]iYb.r�QqyZ��d=)}���X���>��梭[�X3-p��\~'ϸ�ݗx^:�I���k����ڹ��{�<���!�"?5 -ɾި*��#����/�˶�W=e5�[�[*��,B���eje���T����J��֮?�eC#$��pZ;����w��yv*�<��vOOa�w}�|����U��\!�q-���D��u�d6�2m��1�"�"���7ܱM��e$Wo��ђ�����ـ�^���5�=�M^��[�vo��;cco+
�yiy!/��d��@�q�/e��r���}���R�7)v���~��6�k{����3N���X4���p��D�i���o�Q��x>�3ZF�4���<����
��a�ܻ�32�3^L��gK�/ �k:�\�T�׏U��@��o���6@I�hGfTkR�bls�����ŋ����ml6.�����h�RL<����jC�'s����7u�j�s�nkF��˗F�Q�6*�,mW	�.���u#҅���m�b͕[yc52Y�[*��XU3(�6�#z��i���X
���Y�Ln�<�72����.�=	�s��N�S�]��pM�c#*�&��])\�aּ�7)���-��4J0�eR!c(�k�؏j5�(1��=��6:,%�z�IDRI?x�l��{�~�c"���&3�.�8�6�^�d�-�Y�a���[�#&_�~P��Wf54{%P�NF��9|�ߚc}j��/r��\��e�{�� v�GJ�'
�T��9�\�L_���4�>�Q+�bS��w�5���@� dp�������oj����2Ҩݽ*�>����W�@݋�V��MW���Q�g`�J�#�F~N(�d儐�.LO�R�2���8���L��k��k��[��.��k�l�
\y^0����3�	�]a�Z
��v��a�!���.(
d����e���"��'wEY۾��N=7P�݇���d?g�Ԙ�ղ�}x�D�s3 �寪�5z�\P=v(y}�68�-M�nk�X<5��CK@��R-(�	]�����J�h��ds����g���Y%������<c�J���Wr4.zQ��O�e�]��Y�~��w7�q��<�׹�fr�ePR*�MQ`�o�N�5�V�{��kX��>>��|֣X�|��	_R����*�&w�e��xl�q��V�r�c�T�����j�����5�ҤY���9�:���p`�v�6rv\�PС}[a����"��"��^�Q]��tw�}�RO��wBx�}Q[gLL�-�'Xp^:"��R~���$2��[u�3��Z������^|�t�g1�z=�(#��_��G��eQ��
��/q�[��
���2&�L>^�C���<����	��L��]�2�Z��g���Ugs=�ͤ���?`���~�1L\�[6x��9;*o�V���Ut�NQ������6�=Ug/�x�0�@����=U�x[����}	'�X���ų3=��L�{6��Q�����0��Gⶪ�В�f%�c6n�f�Y\6N�9��	x51#V�M�E��0-�khB�\A�4�e��g��|� ���Bͼ���'�u�{���C��� �+��+����,�7o'�C0�b-?&��s���ب�N�
�ȉ1Ěl!#�W�Y��n�?����}b�Cx�u�3�~��G�=�0p�E�+al�����8;;tW����1������wY����G�ŕA�؟D�9ĺء�����������k��C ��������=O#�0�a]�_u��l(O^�Yظ���͑�R�R���v3�V:��0��vUvq] �݊���V���p�s��B4����Z�(��³���5�sx�%�p<��u��m�ɹ���[B��L��i0]ې[v�#�#W���q��l<C�|�|
�ٽ6���������y�����,Z޾f�Sz"��a�SV^�x���5��*m�ڿ�>b�K2����XC`��Z��;�ޱ%���eY�r��3rVr�0�õ6�P>{�&��u��j�j\�Y0YS���)��s�o���*��țN�I{]�ۺ,\����\����o�d��op�|۸:^Y��d^��wvS���-1���h�"q���� ����{s��ci��l�\G�明gP�I�<�Sp`ʏ�P�[s벸v�0���sGe�͒��.��m�7�&�bӢ�݊9��U���H�%ޜ�zwv:�kf]З϶E�=J·r�=�O��wqѦ�ޛ��S�m�y5�83u�B]�ڡa�s���D���i�w8VS!d֯J�;�կi�;72����+�s���@Xa���������`F.κ�*�ݗ��i1.�WRU�2�>�v��CR|�k�";+M}��d�偎泊�����I�z�*~Efރ7+�F�����<��� �'|�B Quv�U��vS�ϝ��F��{C�&͝
)�6�����-�]XU����Ms�\cq�Q�n_�vM�)4�[���q��N���a�ݹ�G��`��uk�1�ܪ7��!}�*����I����p��,����wB�Ce��I��t�d~n���3�}�?l�m��W֯����SB<���Ex:������zM羷�_�e
h\��Ջ�B�sM0�2�Y,��������_J��;1[-\Y�tG���{J�6������*lx����3}
��C�+钀�(�(b/�����{M"�\�B�T��"����N_�L�i��K{>B���������㿘�Ş��9{q��z�Uzq�{u��f��[QqY7"ݹ�M۟�Th(�z��m�x���X��}+�q�?���{^q��c�Scg�Q1�7/�W�3}����A�٨ԅ��_�7"�q@C��5b\��\�s�)�*Jrꪶ8`B8�(K�WƬOg�_/_��<>�@:��/��i7��@3g�~���K_@�w���vX�0)��U��VZ�D�z�gz������?J�[�aD$������> QE���׼��´��R-�$X.U��7�����z���r�h�)e�#����p(��T�bJ~rtYS_��Ϛ�j\�,������3-�b�R|�R���J�eo_f̜?W!7}��޼�_Y�n/�4D��(�{H�������YC�C ����G|���z/Q=D�<�	d��l�a�;8,hwՓf� SH��ċ5]�G<������@]"�4�̰�9�8�^-��>�/6�\M��ő�T(�E#y7��Bov1���=N�g�t/~d�ޔ,��"�#�=tӾh����B�������|H�%�݂�XGE$sp�-"�>��,PR� �iDxv�٨ivt:��d�(H�%��F]��BkZ��0Ú5���+*ӕ�(�*�JBB$6�7��FEh/�=_f����b��g7X�}��hG��[��� ��Х��>߹g30����C���U֣�y���<�a7b���E���U��^�U�W�j>Ɛ%eJ��D�h*�%�T˚.8r��"o�Qd��>���`󳺉�?
xX�>�~��t ٌ��D?|!@{�R��Q�)�DRC�j�|������ɭ�<O�qx����oc1�B��Q�eU,m��X%8��E]������(�U� V?��Ϯ�"m� ��4�lff�uO����}ҍW��Gѯ��:-��������{E��~�@dQY잲o[��9�Q5�{�,��bA�|��~��-���Q!&,��U�  >8Yw)X��w-/��i.	&pQҏ�G1O��ku�%-\�p�"�9.�v�-�,��|�|-��� DB8Eϯ�����!�*f��"�#�j4M	P�HN���Z�� N�]	*!J���_]�3R���jb/�J���:��:�-C� ���I�>�w�}d8����A#��o>�WM-�X4��3���)�B1Yۺ�V�g*�(�ެ�rs0.�΃���uݗ�T���WN��ڎL�x�z�j���kk6,,�n8�v�hh�7lJkrW��/n��z���sy9{mmh/{(s�c� ��n��j�y�n^4t���0Wa]l'.�O�O<�;o4э��GYA�s��i��s��wn2�WVV��e�e"J07�qv�\j&x�g�ǖ�ں�TF�Rh1�5,n�R0�M�ݕb[cl�a+���0%R!�ccP��k��\a�ܖx׭�m���=y���el�2�m\���!B���.W+M��Qk���*֪Ir�iU5Nj���KښJ����x��&���|/����~ql7�֞|%U|aTx�.�������j�^=�����!���s���]��K�%$���jb͟�.X՘�m�$��Z���>�v>���"���n�{KI��Շ���}��.�=��*��P��ˍk�������,��V�
��Q'����8���@l�tR��ޛ;�}�5����W���**���x�VY\jH�U���,T�T%�b&�\��_ �}��`�QG��޺���8m�v�G�3Wó�}�BY���=oX�L�������"�BC�S�E%���%ϸC���a��:��*��>�V+[c�{_����)�Gݶ�Ys5bKI�	ZFgf4J�D/���qC�K���į���-y��2��t�f<��W�f9��i�� R=��:������L�GlQ�e��b��3$�����N�+sy�q:�a�Cӈ�)M�|������ғ����(]
����(�߷���R�>ם�������p]��ZA�c~f��Ё;���h�?u�7bi�vYA͗(Mr��ĭ�D(�h1%�Ý�@���G6��h�m���!�5�[�w�/�MKPЖ	}w��7	i�v.BbX*!P��*����h�Ɉ��	�%_~��:�^<k��8��>ԐR+��#�:X��s����Wq�p��PG]�{�M�{�i^IQ�;�����.\��d.�zP�G	v�tM3�{���pީ�N��h*x5��'	�;q�$���:�∪\�_w�.Ӧ��.�՚��>�k4�[����I�C����G��e%B\�N+@���H@�8|j'�*�����\"E�.�e��{�.�,$Q<�ֳ�Wo/>�4Eł�:��y*9�!�\�ʕ8ے�'B�ރ�E��y���1�愸Ӳ�:��.�H���E�}t���yӑDtK��]�NM���D�B�%��(S{�ܬU��."qĊ�v#����᫙�R��Y�ݟl׏�B��⏨y��^|0�G:1I�F���tB�Gg;�;���ʅb��䨪�ޖ�l���L�T�ej!G^��bA�k��f���m�i5������}k�9��\?}3p��$�ґ �*:s��׼�W��Z��ZDUrb��	�r��Պ��XaQ��D2��h�3`{^��5�,��B�T�V�9f3��y���N���3v����nt���<k�!�,�p�\a�	��k���ۉ�b�X4���F�*Zp֐��ݖ ���^}���m��Q$�$QDr�]��j��p�݋���[�A���jL����Ԭ��d+���;o-:Ԇ8��A���J��ӿh���F����LuU����a��`�V���b���z+y�p��$I���ެ[�"Z������3A��Dy}㖀X�����<�<G����
Ӻ���#�C�'ɽ{���ZJ�T�����owׯ�a��_eL���~�_2z�n���j�z,b"�l���?q�Mi��^[Xb�BH��d�(n����+Z��t;-U��=�E���������U�I��u�8v�'�>�g+��l���ڔ6/v��ȰK_7�^ʹ�OV{�����!����ф-%�(� <h�êzuhKN� �4~ru�fl�R_Y~�R ������4ȳC��F�<l��>�U�Dh�j_�^`Y�m��h۬C}�j�9��>MP���gZ�;��j���AHR��B*��>!h�ET�˷@��^��V��8!T�^u�{|Ӿ�A��g��d�>�8��� 2>�*#뺾��_����j�|k�K���b�De���P2l2+�6,ij�ܦ���M�Ѡgb
U7Te��i��a�c�j*���4���bL�ߦ�}�Z�6Z�TH�g�~5�l������pʔ]m��|��2=�� Q�X�/�?a�|h?�!@і/�HD�JH��:�q�	�����ʅ����ѐ����"R�U$>si�d3��+��<O���*�D�����=�~���A����V��W$.�gW�Nđ"������˯�
hT��#~I���K!�d~��}�N�~�C��f�������%|ǀ� JÙ�^��~񳣐=w��\��,@Co$gU�6���Ⱦ!�}{�>@��ʊ�Q��-�N�@DQ�r�S��W C������J�Vi>d]/�������� �T��r�
ń�!�D�.�Fk;�v�^��,���)��Wy;�#U}}�*��T��uv�]��u�3���3{TUn�E�&�[��h�|��j���~ܽi�y��S�Y���.��!5!TԺ����e� C���+ﰍ4a�F�j�G{iZ��-䠪�~A 2O��QA�k}���=+�G�l�v;F4Q�>)�d���1��ª�qEmT�w,�iH��\;j��r��j\��ؙ�9�^2�=n|�/ha�
�XF	v����}���+���^B��J�(�������h���ݺ��!�f+����}o��R��	�W�Z�ꐚQb�Uz]W�j�$���&�H�o� ��
�Q�4MUL�T�;�,�s$��\'��X���+������g�^��O�������� ���^+Va&��>0���Ǐw���������>��]�!|�Ё�<�p�dh��H�3��/�d�cJΑGj+y�bz�1�ϡ��Ȕ�oP��E�z�~��q�hX�	p���l��:�gi�	������u�c~ϼFb���4
A�͕�i8�rJl�x��6�fɻ�b����� e�
��8o;��`x(��6`Hp�c�Z,|�� ����*3�V��!��#V�.sK~�DU��v����~k�&��f"!���r��#�WR�H�+�T�&�S��3��Rz4�z ��)�����k�8�aQ	�����~����N@��SU��C�L	��s���ղ
?��fy�1i������2W=E�K���fo��U���1*t嵷�{o\\˻�nh��m�/�,��:5iâ�_[\�X�[,�и白b!�p�(�\[C�n0p�U	�+���\G�m�h�E�r�Kb�pA�.�ع�Q�,&x��8�'S볎����h�l��]lI�	M]1�i]�h5��	��͆籊4LF�v<�.$�rwa�G�|o/c�����ϵ�O�pQ0��g���ש�wd�j@b�VSfUl]�M���7��1���7%S���V޶v-�@��,�`�ڴ��2��n�Y��JU�ii���U0��1Kmŕr˗�Y�7�O�?�߬,��޶��X1��p�D��G�I�M����BV�4G�P�;}���ѱ٥j��WtH��c�d�VhO{�Va��qC�[x}z�����] r���~����@G�ӺU�T������.+K+qK��"ib�����0(W��dh��0'vY��W�����T~��v�� O�uZ|�sz�vң��'���WӋ�N*�
��2�lY�a��p���tz�Ɛ�����Tċ�{]�ԅ�Bd���ul�2�|*�������T�4GȆ���y,RN`�\�L�F>c	?|غ]F �i�S��ݡn�O?'��;��6T	?J����7H��c"�#�QϬ*�����@l7�;�ҾqL�����n��7|9W���Ј�� |���x�C���LX"���XiS���e�k1��~�)8p�f�W@�%uH!��O�ax��<]�Y|��{x>�5�n��^�DX1�v���R� ��@A[�2��>`��?�>��������f|j�I&YJK��{n}��C��9�zP@%{��j- �K�,NT���E5NS��~K����p�U�Z�\'�L�M�b����&R]�DJa��M�X�s�nU���m:7�5w	k_z��g���/�H*w�^|���/y`����_ߝ�pu2���?�:~l����������h险�H��}�9A[\p��Hn�R�_n�Е�
`�;\�3��	C��nf��ŢQ7���t�*�0��8��N9��3�-�@U�9����cI��C殪�T���8�gD��W9P�أ�ƫ�|W�Q?`�.���^�X��@�x��W�o�l=h�h4a?D�#��W�,V>O|���U��/.	;���d�W���0�;��x+���ME���w�����p�u�_�H3�z~� +����چ���Ĳ@i����CDF�#g�z6�.�{�Jg��*�ȷ�a��0$oR�H�$i�d�ib-ن��vLu o��J�(v�������PaNA��p�=L�6�����e
?,d"�%��_x����2����]��{�/�x #1�Ѝ��+Pꎹ/]��L�}�gB>K�?`��p*�~R��,}W�]��_3��c�B�����
�%,�Sq���~���Q=J�G;�� lh��ٔ�9�j��m�y��d���ٳ�M)�����~l,"�u/���6!������ʝ��}�]��>�YH�0�p��z=Ns';��]�X���D�bl�B�T։����dF�uՊ��������(��i2�y'�[��<��6�ݏƮ�ho:���L�{ow}�
@Ң�󡾅��2{�x^5T mj�I�o$: ��|G�a��{i�����";��X�Kr�?u�Y��9����.4᠎b�ax�,?
�`.�x* a�7%m�@^̂��9{����v؂���29�����+Uk�FiBg)��t/J U�l�H���&��v��;y.�B��������P�&c� p.���S,쒧��<�+����HsA�Q�\��9--"�}�+(��u�C1��d�v��dģ"1�XDY�{m�00�Z���2�t�/��u�3�p D	$��]��쫆���D�G� ��8��$"�%d{��j���ەcۨuc�M��/|����kBV����C�^(�U}7h}�����G��v!wljڒ��@�"{1��̥�Y[���6��E"s��+���x��}��#B:fҰ�z[��@��
�G�k�;�x�<��)w�&3]�a��&�.;Fx��zN�,�w=�Oh���Zð�H����M"�uU=Q��U::pJ�����.��x1��*��D�˴9.�,:	�V�U�+�z��������*�q��]�m��+1���C��즈c$��L�c�y��l��iH���\	�+W:���deJ�]�6Ia��u)3!?/7���8�.+ B$B����}� �b���J
U���&~'e�A�Ͷ�%��0��,�޿�_�3C�����[�a4#G�G5�M���_6r�Y��wn΢��T�C�v.���;��aB�5��PU/�x���!!�H�I`{�C��MI�}­ @�����SpsI�Uy��23J�k�w(�$�<U:.�B�_U���g�޾9&���X���D	�|�fN5]��ƉXP4���މ��أݹ*�4��\f�h��rZ��SŇ4�������#�gJ�s��!;�ꥪd�}��q��I�ȣ������@�.����SC�~��u��jq����g}n�^�|�� :��_{��d�HE"���m<vݳk͚R7긶r%	� V�X�3P��i����#�e���͸��U��Ѵ��R�MXX˅�U�m4���={�װ�)�h��k��|�`"O?�@��(`���T���wk�IW}�~���/��fC�u�l��d�ct�hU[�����q�ʉ�
����]�d��.���g{} 22��MrD#��s�s~�kEکA�j*����ϱ$Ք)%F�?s�.�R�;�s���u=BE�(د��BD��J9��~����R����i �뵀��=�|�	��_=���qrtfV���6</zB��(����Ȗw���vH"FQ�'�I[��!,N�X�\��,(��Bɾ���E�f�7��sⷮ�sc'c�T��ǲ��N汻P�Q(�D��N�������g�k+�q��fD"͢�3�|�1�sh\�jªr���P�$�DG�P�$�DG�P�����������j������%	%��JJ"#�(JJ"#���$�DG���$�DG�P�$�DG���$�DG�(I(���%	%�%	%�P�Q�P�Q���$�"?℡$�"?XIBIDD~В�����!%	%���������e5���|�`S�� ?�s2}p#A�;J���( �]��@���  ���:�WT�Z ()�R hR��b� hZ	�Nڂ�h�( ��@�"�E
�%)RI(DR JBUJ��)J���T�@UP�QH($��
J��D�@���UUa5����ҳ{s��m����I�r�K�wG��T�K{�ͯa�mKu�b�A�w�tp�޷{e]���T�����ga�V��eP (�*�v�'Y��:�p�S�t����
MQ���[-�mb�6�ê�\ZQ��@�޼�k�T�
��+�UB��
��8*U�HQARQTB%E]ʥ{{���A�;t���u�E�;�l��H7C[`���l�i� ���F�� �7*���Uhe�ˌ	�8� 
�R**�k���"� =�x�	�:NME*	w[�kS`ۮ�c��QnTJ,��U���� V��5�EN���73�h�  
 �ꀕU �"�(PD��
��G���4��ް���t�� x��<��˼(Qyւ�(D)�4f S�g@��(���
 @����A�P��g�g� :��a� Ҕ	U��y�.�y�8��CCA��TJ����9��
 ^` �� <AGl(rk�{t K�x)JxhPz �a^{ ����0t�X 
<���
 ��
�PH$)H�D�
��R��)�ԓ�wIR���-����PC �uT��P-��"�,[a�ZVCJ"���)JQ�(J�t�����Z[��RU
( E@�Q.��	�%Ps�WAs�]�[��D����z	������Cu��TWv:�N�=xC޹ճH�@){h Wz�$)QQUQ!%#r��jRU�:�Cv8�R����w�$��sT ����������WzϠ��l�<�����'m���OGwu�h�$�@+h:� �hy۠�aA@ 8�AN
�h]0���#@v�J�K����Q�ɢ�i��(���lkM�9�mۮ�����v�u.��j����{0���`��BeJ�� �EO�
JT��  ��LS�UL#��# 5<ʠ���   ���*z��  = BR��<S���_H/��Q}��`>��y�9�䚥��{���_33j{����Dd�r�E�!DF�+�r��""D(��
!(��!�!DG�DDB���DD(�QB������7��'�>+��[�Q�!�+�8��̵Q�h��,�:$�И�Y���ϥ������63X:��B �Q�{��g���$k��l�7\�%{�J=��C=%q{�Hmz���`�����3a9w�يnt�z��/W�\N7���P��I���q����q9ݗ�0�:,���4AXHb��1�f���$�����S�kx7����w7�UzU"��x�Ɋ�ǘ���Z���r.�p�	g/`׸k������z�&B��6�ί�A�y��~էn����N�9ex��Nܜ��"�p0s���n���雅VslR��?`��%��),��t����5YMs��n�w�+n(��0�::��\��p�z�-��1&�_N�ѕ2�,z��w;�d��g]Q=k X�vs�
c��'u��v:m��og�GOW�������WVBJ~�b��ڭ�R-��!zH:c��j8;�E��JS�*ӏ^���3:�ؙ8`VgW��8�	.�v�R�&}�n����b�ގ���l��D��Pqf���޹.��H\�H}�LUr���W:���6�e:�W�6�>�(�p�� �yQ�aR�**,�d=��YǤgu��֡O����Ǻʥ`�u��$Θ �C�M�ܮme���۝;W����?d�9�\�NY��`6�VO�$Oug*P�q�$w����:/.]}��^���N��~�'I�Ħ]f���8󨫤� �L�p��FT���l�m=�n�٩k����غ���5C���.�x·����YcV���&IH�:7t͛�Ak�;�l� �b}OT;��l�억��P*z���)O[#K��P�v0ݧD��o�&�x��E���y�KٙK(І�z'NU�*+�Cض"p�њlYF��=(d3[�xI�p���b�W9s��\��S<C����ơ휎�1�����&!�p�
�q}@�X�9��YxU�������kx����[���S�i�.N$��L�7Gl�&�(M���֢���ݣ��eaa�h<����]��� �.ưz���Z�J�O�I����La����@�s2�TxT��X�<�7�w5ʍ�@ї<\�dC&�V,՜U�����1rD�`��(Rd_x�Gn��6cǉ,�ukD��n��Tn��{Yb~�[z��9^{�aWa�	��=���P;t�i�S}b۸��0.TK}�Etm�ɻc0�zA2�v�Ԕ�5K/*T���1�O��	���"*��c����[X{V3VK�i#.��0��Į֏+�H'\�nT��6M����#���D�����Xt�:ٔ��zޔ`]�Hpe�Dx�]N�8��ItG�u\�6Pz��du��j���-|����eJ��#��cv�s����>�v�x�:�.۪"�
-%AOc�x^5%�������$2��=\®�	f��nP�q^�:�;�4L��R����чc�S�ݼ3S�7���!��x�uG7I��bV�J��\�D}ETLǩ�w�W�E�<�c�@�	�a�>��$�0�a�v#t����b^x/m�ʈL��Ƭ�UwV
r�>[���[�ʪڲ3)���`o'����T�"���{1�3�E��I$�P����nm�갆�D���q�q�f�e�[�\"�oTS��œ�gJ���Y�bwRu<Bod[h���*�s�/:�k"�R@�ὤmQ���	d������8$���p|�Փ�._�+�^��@ݦ`6n��q8�WHlj5�"����mݭ�)����L�y�6-��[�+��T���E����l����!�j&:3R����q�S�I�,����U$�]�Z��S�N�u�ҏ@�q6V�F�΄B;VB�m�,��5J������Z���C$�B��������$��kqqBn��#�����hb���z5��7O6�'�n\�,�]�Е�9xb��xĔ4%����7��Kq��k<:IF^�t,]�B�:������˰IuLA���&���вSz�,"T�.�D�7�<��KQR�_>�_�$^�wx��zj8i+��I�(�K*HgD�X��Ō�Q˔���V���\���s;\1��j�h��7��bw�~t�PR�B�bv��e��J1��2��q�v�wu*�@�q�����%壩���vx:e��Ԍ�ǥx�V�D:w&�{��Bt����F⩹[8�೘W�h��QV�dDB&f�%�݌����]w��x8�]�zcT��r�����$,!L桶/
���Ӛ2����ht�Tb�()I;^
��j�ViŮ���N�A�9k�o��5�<��Ǽ-�w�3Uy�7�I�����'T�G`��]�]����S�H5�`���w<��>�����s�%��.}p�[�^n��Ns8*�x�u�1�œ2�cg�+iqD��Z����;�c�4jK�=�0�=g����3W^���Q����'3X�! o5M9��ݘ��goQ�Q�5��C���u�]z���,]1�ػ��%��/m�]�{��q�s�3��ɿt4Ƞ7�K����]S�{;grɱn}�q�y�1�a�Rb��mY�#�klBh���(����,.����gc|����s����w�TV^�)�KÏ]��fnIi��O ˠ��t7�#�?$�Ie���:�v=o[HX�Uw+�hVp�)!Z�O��9E^lr砻7�Q0JY�bK ��;B�]\v���&~���0���7�Qr��*[5�Ӈ�qs�M�=�n0��/��5�1(rr�y(���K�-j���N&rM�B��Cc`�kZi$��� �3�v<%]Qɻ�T��B��7j�sN23���g1'J@c���7@��El$�s�4�)����ժ��B��S#�V�9.�pl=׮n�;�MĜ��7�9��z	�˖{�Q�UU��i�1=P�Ѕ�;#�v,�o]��m�ٯA�X������w��ג9C����^� / dfu��^�D�a 2�`�'J1JI����0CZ%��^L�Q� �h�N!�u�;���6�+F쿂��P�p�gUs���MR
��U��$8-�F��%���I��o�1�@����g���3}��l֐|-+\���� �W��<�[���C-9�wC�vSgB�5�4��p2f�=ٍV@��] B����s�O�Jh�{��iT*e�7����t�{}����]�\�(�+�v����䕼�WN2Ԥj�ʹ��]㴞8�9)�T(�� LP���Z���z��ڨ�rB�.�it�}Ɋ@��5�]B�s���vWJ�.i~�ӻ �������1������Ꝫ�12y5U�_�,V+Ё����)�û�ػ��>�\*�)j=�qQ�ZνK���u���Qhu�[/�^��w���rw��sy�%R��;��H���.��8A��M���h���_�vK��A-mس�TE����B�)?����B��at&�kؐ��6#�M�`����'$����qN@��	������/�O2�@�;)K�).��5�Uj�Ȟ�J�xw佴05�"�Q�����a�3z{�s��Sws����]����ιR�k5��'.�ŭխm��F�<�;�nMǂ�^�&�-=��q��n]s��nY�WLI<0��{�dW*�6%fRE*Ʈ�mN���v���GAk��.�d�z���{Ha3(�f����?q^�O�V���">�.˹hԀc�Ōn sSȀ��6\�(�#_h�QZF�5�#9� ��0�0�mv�Ӈb��vq��d�"%���:j�ڈ'�"�n{������#b�^�J�������h@XÕ��v�qe�5�\���XV-��=;*+(�n��>ͺ�E:�Z zn4��@���Ú=��2�����f􄗯'��7+.�f�W�Iį����/'E�e�'K��5W��������*��4��Wl��{���;��*帼�q�`�Ż��<��a�nv��Cݟ�y�|P}-z�ZXm�S�5������cSRM{�<�$�����;��;�{BQV>���~���R�������Iu����n�EMjG��L���f��V^L©qY�^9n����Z�qD�}�6E���{��\�Z�k5S(��A�H�1��̓l %�a�s���0�d��H/y�,�8��H�����A��j�11k!�j��]u�Ux�9�/v��Af�qv�j�Ӎ�F�k;�K�}YD3*�LB*�L�<iSDr�M|';8�˨l^w��ŵ� 1e���_�z��ӱ�9Z�)���4�W�%������b.���F̚nJ(��7�G��a%���f�=�EUy)H��]RYI����W}
A�tv��w'u����Y��"��$~8;���\׷ܴ3���r~������p���;��GƉX�N�wb�@,2a4��y^�m�E�ݖjl%W�q��Xl��o���"�S?��2���O��ۺ�[f����p4�[-k��e7ף뙹�1�K�N�4:�<���k+��p[sw�$㋍���|��CNl��Jf��y��c`������&̈́<+�m���}b�*^�uE�9Dahz��'�/�݈k�d�f�Ҳp�ԁ������y�)���A�FM��6���"��L��y��m�E!;�s#��m�6j�L�j�ob5��H���a-Р=�����p�U��/h�'��n.b�Y����n��>e=V��bu��	-��{�e��S�H獮s�Waۡ��w&Rj�4c�M� А�ᗡ3$�]��/g��/�-�J��G��d�`�[��-|mf9�&Lj�uHvЏc�_æm�k[�H�D;�����hQ����&ΦA���؋��Dp1��v���>�G�N3��j`��7r\�wT�����]�cy"g��x/�?�L<o�+�sܻ&��	�)Uy��$��x�y��>�m�\2�w��Ku�
���=��l����=���^N�䙠�2�	ۖ��Ww����jN۽��k�Z�f�-���0�0�i�Y�,ٛ�`
jf��nn[�z0�h٬T�:�_�����y�,}%���\�n鋊!��׳[���R���� L��J���1��0V�'�lݨ�w��II�8ʆU�M�1�_%mi���¡yu����b�5!S�nn�L��7�-R�i��
+9�My�����Q�d�r ��Ǖ���T]�M��G�n�w.�槐��)�f�V�8���ͩso��ә�L�E�R�͙pE&���!Gc��f���oI��S�1(��3���	��óv*u��K �%�6����t��S�"�v�EJ�]�R�`;�M�<�ĳ�dj�=�>�:Aȓ�N��H��a�a`ZMd99��t��Gӵ�����yj:��cԀ�K�Rϟg����w�D��m6=x�!���-}��ީ�/cNf��T�+�6<�u`�8�(��x~��!a˪�g's��O�#5f��9��h|���R8�f�GZ+Tu����/�obBʱ�)<W�X��TW@گ�ޡ&,$���i�pgm2�z-iD8���W�W
۰e�BK1�%W������4{k���'TzSvRO1�j(u��n�1üz[�t���P_�i��2�%��Bz�u�ù��z�����c�y������	���ô�q��8����@ծ��/7s[%ۑ��;��M����K}�<��T�k(����]��A�Tk���������� �b�=	p����*y��Ic�X��K��Ӷ弐�����6�Zk��A�?��o�#O���8p�f�ќs�q�&:6��z_�5Ll�\t�x�O;S��K�+�f�j�[�t�-���Yo�)����d��Y���E�	N 蕚��op�3���f�k�6o[��������y�^�˛��Q�rbqWgn<24l�Z8�x;Y�������wrԶ���nj:M�mB�{�^�(L]�OQ���)	'Y���LW��wݛy�n)�L�5:hq�V=����� ��Lz;:	ӻr��QюJC�[;nFN��Z��;`�|���������82θ��Q��K������:�;^ü?XU���˰S�,���g��Q��`8K�I"a��C�;G`��l׻�f�G�o�D%h<��x����fͺ@���6
��n]�t��qՀ�{v>x�X���*��q��@��M����ä�)�8�ͰU�3S�WS*��
��`k��[�m2'���M/�^ޓ�!ٳ���/a�O�g�8`��b��dz�BQ��0s�1�2�jŇ�cYR�N�F�v��+	��wvu�㚢k�tw�����xd��͇r��Б�;X�Q�7��E��Gا>zxƩ�ɍk;�خ�*�4�CC��!�`�縜���q�- ����yn󈈺�::�"gk����#�x�ʤ���`�{��'7�S��E��{�i�$�&�/���N �8^���z"����gS�3�D[�nlB���,{�U\s�T�J9�W��W����bz�֟�T��	,1�U��#���n7�t �V�8$<�H�a�q�r��)��X-��u,����������c<2�%E�[�ʂ�[�V���r�v�]Tv�#@C ▵�ݡvh* ��Ͱ%�8�A[l��.�*���vx�eaٍ��맺T��Ů���K�um�Qψ�Ʉ�yk�f�����vb�f�(5�[����3�cW�ȼ�S�ێ;D[�X{sڷ2ܝ�8��'�V��n�ᱮ^;p<ܝ�k�f��^��OO��W/g{/>pG6�{g�{����ܦ8 �a�c�Ŏzz�ˮ�H,�y&�ܛ.�4C)٭���p��n47��PvS�,C�8���<����1:������v�5J`�t�����/M5C�˛rD���6���R֮���Le�w�tQ�r�1t��A�����i.G.�`�q��LlB�9*.�6���R�)ʃ<nl�ŴF���imx�U��#Cq����D��Ȳ��́s+�v١k����й�X���*�����c���\����[�B��g�u�,�)�ZѺ������y�h{U��2JYLAᬽ�]/B(`bk1�R�SV"���6��P����zzM�������n���gq�.��t�ۤuۀ�YNqqi<��M�V�:��GfZ[���Ğ}[׭q��4���h�oM���N����8�Z4e�Ú�FX�����c��8�"6T��J�r#s��#��{oY��؝e��t�n�L:���j�u��{��7LEլ�����t��x�%�
�,��gJ���;v�squر�wnʉ�P���I�P��ji��]J���`ĚM�t��2�C�]��\t�Q]�{�'X�'���k����ƀ�n$�<$Y�g�-9��d��ۙ;	x�Y��D��:��-8Rn���8���ĲRiܣ�.(5���\s����o]�ԭ�k29��E�a0ʚ1ں���Iq/p���1Z��][�'v
���`zI��t�6^��)��:{�2�ML7���+m��5��f��ߏ����Oi^|v��x\��x痵ۋ��sl�ڻyy7\�q�cO=:Cr��Z�����x-n,0�\CS�<ᴮﬧ/Z�VK�4m���n;c��,8w1��]Fh�]��R�ʼ[S�"&�9��\=o_?a��tC:.�
;JM�ir�l���Ş��J��{��/�'nrN��&�r����[&L��s�;����P�]+H�4I,!q�i��h-�*�g��]�1V����(�:���i����ݜl�n���ㄲ�����%�&Pf���5��g.{o�.;�|=��]0�϶{:XLY�h�0��XZ5��ʌ�f�����Y�u�OQ�n>� n�s��s=�ے$�ˣ!J�N�eke��;R�e�ǰ8MV�
��5Χt�����uБmrq��:6j)Fi�����k�Ema�X������@��-�V]0��'�nVgI��Ƚ��E݋��q���ݹ��d�j�fmL��Y�$��J،���B���,�ce���2�cs���V��Nz�m
\)���I�v�%�[bfBV�4᩵ ��<��ok��K�wv�����f���.軒��{��WkI�vH��ֳ[n;�E�8�;��A�/d6��D��h���
�J�(�Fˁf��"���]�Mf�]���6�s�R�Ȧ�Ѫ7C��0�KZ�. -v�%1-<딢�f[2Te����Z_u����)Į��5ute��V��E�aN˞���#�%�'l���KXg�z�zLˠ�T�e�m�W(ͱs�ΧR�s,�IP��Y��-th������i�Y�.z��>ÌC�[�l�
�q�ˍ&÷�L�b{/<򝪁�#��立p�׍��V�1J���� 
j�6k���Kq�,(dGc�x�[\X-�Tv糑�F�I����Q��bc��`��A�ZMxv�x�K�l,Ck@����5	�ԙ	�]��Kvnc�
9R�a��f�m����HјoP��`9�]�볹^א�K`��c�A��[m��=�q� 7mq��J[j㉑�����R]`$Q�.IP���I�+xXR�8`�JC&�O���nS��<��u$:L"��6�c�;L˂�D���h��,�F�XݲBT��1XF����n-Ύ"�I:�����L��am]�ұ��X�!LFlX��n���ͦ4T�nc��TO=p	sĸ��y�y79��N���	���������jx�g�M����9c�%Vp�{X���ɘ���j��k.�m�4Z��sK��b+q�c��Nx�{]&;�E[��/Zkb�M�F��:w�Cz�j�mȳ�s�x�V�]��b�4e�3kh�l&&��0���l��<��u�t���m�D\��/-��><\3&�E׫P!��3"�F��n���D���v��caԹ�����A���8$��4ax�3\ո��0�Wy�Dz����he}-�]�QӪI�	�;�q�i�iv�ػy�r��W�^�
x�%��h�2�i�[ۭ���"ʧ�M�:u����wN�8��-���g1Z���7#����\s/�U���=�y˛�[�Tk{[7S�t�c�����䍝I�8xL����:�0H�\.��tv���]�����im�K��܇m��1΢�� $�V�{i�<l���~������7i�<v�A�J�Ƽy�2�SX��W�V놶�"_H��u���n���h�[��	L�]ɓH��[#n�J+ݲ�۷�����x�������pt�aή���*4]���J��Tk��>������baz��9����y�y=m�K�CY�m���3�Y��U�Ω	��q�û3��x�)�&g1.��N"9��ĳAl���yn�#�Pg��ȗl�҇n��2������gq�b�qn۲�K�i��n�n�V�5!
`]lf�mc�g��7���7�K1���{.��6ʬ���6{si<,6�Qe�eּvź�h(�Si1\�z�J�H�Q�&���2�XKsHCh�&y�N3��e�ҘM��T�a�j� \�ks�:[++1�b�`*\Ճ.VkŔ\h�w�=���q��;y\�]nt�8��n5���F���;���8���"�:2��{�v��bU�M�Z��<��;n�x8̙��zv�DaMv��k���m�5/�w��ҬѰH��f6VgK��fؖIk	�\b�iŸ�;/�5��>{:}%3�G
�7學m�ݸ�z�v��{�8����==�۟&;ra��tn�E�x5�1Ƹg�b<�=���5�bۗ�Ų�$��9u������V�l�HE�Z��b�o��Bh�\5؜\o��8ҡ9\i�rk�+/�F��T6�i�k� �3[z��xEYe3�(�Ӭ�]��9���g�.2�,��6θ��g����Gq�5�<�y�ģj- �ՃF03q�m�"�]9� Os�Z9�\Oh��Ũ���eF�6D���⒀ʓGk	i �YB��%�6FD�p�ݍۍ�:� :sL�gEZ:�.З�@V�
�㞬��nVjx��܋Ćͨ|���G/��rC`�oC۪Ƹ�d��8�ȶ���6� :x�{8����xS�������L�=��r=f�äf�ۙ��r.�Cr�hx��ܘt]n�f�㝹�8�"�Ϣ�a��sU�l���W(�m+��S��9��nu1\!��aˬюricm�Y�q�<]���.c9�n/���%NwAp]���v�O���X�l:�BI2av�`8�.6rs�q�l������n��g^u�s��䣶��3{6[+[�v��]a�M� �^��϶Cu�z�u:�aAl�Տ1Ͳ�8��=�ʰ��n�#R��:5�i�V\�B�$L�Wp�vp�T1�t�à�6�K��Hm�bҴ.DX\3�6jک���n������x�ŹL�Eǧp���֝���	vPɽ[�K'p�d{p�q��+��uX�h�م
�Q��-8ܰtxʽT�q�_\�׾`8��%�[wgq�E�p��"��꒮v���3%�����Ʈgb�#����G��EW�`;�ѹ::q��s�yn���<a��a�8R*1���M.���'�}�u��zyƼ�8t��=a=�z��mX��a�SF����Yn�p��֑,�����8�!��� f9���D�8��0cI��3hs.�8V��V9y��fG��˶u2��iGL�����$��ˡ&h�k�6�Xz���7��N�q�\��b��M�SU�0�J��#�c��LYZء)��0�tA�}� &a`Sv{,�pIc7'�^({qƻ<�<�:��C#�q�ۄ<C�J�"��,�>�㮜.����9�9]��6�n���L+�X����g��y������ӟp:Gv^�:9s�%��&G�`�#ru�,b�X:�kL�xУ�b�(�l�+�WC�ݸ���f���)G("r�XR�5EaP�7qr2�T���#��\Fm�`� }�S�xԾ�M���Ӏ���4h�2���Nd��HK�Ȱ����!����Ƈ6���À;qv�����:�^GrOrv6(�lv낮;���b�jPؑl�f���y�M�ƽ�]�7k��U���:��\�W���	��Z�p��a�޴vK�����YrwI�zЅ�<&3q@�%sk��j��A���Qr�.�h#q�{K�Lv���(v���p��=\v	�J�v9n1ev�&sy^nv�ۋ,nC�v8������N���z�잗��Q���5���3B]kz맅Xf��b�W<P�@��T����؎W:9��c��hu��k(n�0[n�8�yl���n����kv$x.��ظ�[\ֹc�i��Y�K�+$]4g��'t������Z�p�;�-Ɖ%,e��5V����P�4���Yv�s�m�{%�R-�r[n�,]��v#c#5�8�@q��to���蟘�f�,���ֽB�ı���#-��������t�:$����;g����a�٥�(	mۥ2��J���DBQ	DB�B�Q��Q	DG��DB��(��P�k?'��_�!�C̓�e�r+�DhJ�Ȱ+hkt%��^�XR6k1U�D�H��ԣ3��]v�癜�u��Ҽ��������c�8�<��9�l��: �{W����ڃ�lV��.&�)cRU�D�e�#��E-Zi��:I\
v����n�;*h��,����Ѝ�h���f��i�&VKʪ�/6�3pl{�n�=)�/l�=���ɬr�,�n�Z�v,:w`���.v3Er�p�\6#���8Aݴ!��>���1ttip�]��O`�A=���p���f��m�9,ml�z89r�մ��0�� ��|҈�L�ު���N�`G=����MG�V�Ӳ랢�u���m{r��z�e�S:6h��T')rT6���a��i���nN��*�qб%��e��:À�%9��KiL�� k�Z���F��b�%�A�wS��)O�y;���v�ԷHY�͔�c�h�0�g�t��'K��d���9�����{`�K�9�=�[\mh�;=���rȶ�&�<�/�8����B3�5��--��<��1[TtH��.uI�@�t3K�`G74�����%�,-Ik�2.�/hܜ>N���E�]9�����=RM�u;��q����������$c,ۚ7q敛[+Y�Z���]��r"[p;78v���Gj�ԅ�T�0 ���׎�,�nS���%�� ���5���fi�9��h��Ҡ6hhLKM.R��s�eOcN���)ͥ�tY,��p��d!D�4e�7�秃 ����=���6�B�,�6�ƙ�6U�u�xnC]��7�@���W�kL�c�������gp�̝S��$�,$�Pԅ��bkfu����VGen�Ÿ�QO�ݝ�s���)��n$M<@�8w�����^;v;O���s��4\�s�+�sr�۩"�0a�������%(��:.��*�CYW1Im��c7�`���[��$p�U�K,�H\E��99'9���(	 ����B�	B��(��@���$��JD$	$�$����$�%��JD$�D$�D@B��P
(�J���m��%��#Y���e�BYu��&�T!E5���Ғ�g(6���;b�n�+x�ӭh�C�!5�9)t�V��V��X�8q�����vy,�;�� G�1���7E��װ�����5bѲgEt'����V�VƩtr�6�Y�f˶2���q	�5,���Uv��mv3H�H0[�����yіg6�k������W%/M@�<=�u�'7G7'>��d�r���*=����#���s�w~Z�p���E}���e{�j��<��Q�0
z�m���Wi�ߧ��W��C�F�su����{�>I"�!�
���c�3٭Mm���{��;���k_Y/y�5yI�����&�+]���~Tآ�C�51���"���]��i���|���'��B�vs�`�	�߰����w���cx1N���Y�*9��V�}���~���k������vw�$�߾�1���@^���7��6O&sB��kK�����׉=�߀�f���Fm�w���I��o4�����疏p7=��7�\����|s��ͪ�u���A��`��W�w7T���"B�b�p�v��U��.�٥
�2�lC�7Y2qr�& �,z��D!��N�-���>ڧ����=Z_;�~pb���t��,s6�A4�Z��7�`+ŽRtM}���wT�s1paEq�gp��(�/zb{���0��^�(�"ɘSB��>���9���>��V��n�G�	�&zEKz<$��6Y���ۆ9�,����)���:I<�<Y�Ǌ�Q�]F:��/F��ciu�f\�R��� ���9�w�|��Ӓ���2-PMYj����}}���^�G?�ƨ���}��P�x��Z���qonN��woz���@�Xa�)���7��������Ts��ǈ�>+i����Z�TI���������o]�;��z;+������������)���mA�J��|��f����Q�׼����BkO��秇��Ը�VǤr�c;P8&!U���y+�Gm�^6M����C��]�h�h���ޯ��g����xP��l�]A���i׷�7]���'|XH嬆�nn�� �P��_J�[���޹~H�����%��a$��IrC�ե|j���~ڼ���Sx`^���˃8m+�C�~^��dA��ڲ��A�J�����X�3S��[Öѽ�oib`�q� 2(�K3��w��Ĝ��Գ�Қ��o0��ŉB�X�&��*u�VT���CC�QE�3�׈��R�l�w;S�^���Z���v3�z��a{y5{7e�����}�mj���3�Z[N�W�[�8u��N!"�K�Z�����뺗ݔ������m)�WǒZגwr����ë�p	s+D��sI ��:�{%��|����8�1E��q}~��Y���2h��N2�RH�s{���w:����}�b)@�d�8�ozBy����&m�I���ڽ(o��F����ջ��x����a��1v�͎E���oK"���nܾ3sͮ;��,m�U+e�U�.��W*|T��UB���ߨ+��L���l�^�@��Ǡ�@��[��'�����^u/,���/d�.H�5I����?�@��۰A�nA���O�޾K2��}��ezՀ*7y�Y��3�������9_Jݺ(��=�I���Z0%�&!��5�w2�����HW.�3Ѣ���8��4�����j:&�V�5�f�6�d) �8YRI|\��æ�����w^
�pj��T�[��Ժ��zW���)�zl=��5�\�z��w���퓄��V;��i�;��K����v3�����։����F��?*��V�2	=�ͧ���o�݄	$�#RHv��T�p�E�<{�%b
�d��pW����r'��f��J�Ť�A�������������c��cC�5ׯl9�K���������ҥ#��W+��En���c��Jk2L�`0D�J�B!�gǺ}�y�~v<�<L�z.���ŃO�7��{�0��,���i?[z{��|=<3�"��uK���b�B�p1gK,O57�]ҡ��5����`$"V�}���(ǧ}��-�U�SuLe��n�ܘ"��\̶��$��&��j=�Ç/�³X�t�ͻ}���L�:i�B?y�I݃⭙!����Y�s����Q��Թ�
J8��>�#j��O���Ӥi�:�7*T����>��!M�Uo���zN��K8&���	��PW�8F^��F��m�\��Qڽ���Y.ܯ����Y�:�u��n�C3}�u��{���գ<7%���;�8ϰ���о��������F��ݮJ��T[:&w�?{ۜ=�}� ���{e�w��o�`��zvδ_�K;ޒ�~�	96f�Ұ6�C�kɗv���Z�	�����p��J�2��fsun�༮ٖ��۽)���7�`÷�����ƚ%[�ֵf��Rb1e����+D�+J�hM�u�����9v���a�GC�pm��nI�X���pvh�"=����%�ςʫ��V�}�sԼ�6��R�.�Z�Д�c@lf�,C	
�5ʟ�q�����&�tE�W��W��h�',t�����ݸ��"���+)��4��W�?w,�o*ʣ[��w<�����`v���~S^n���]Vw��6f��l�"b6N�t��Q������ONM�r:�Z���j���~�ʒ�=զ�êp�P9�0"/v�I�D������@�M=Iz{`t3lӉ��af/��Ȝ|�9��>�����������[��}m�Q|ID2�ݽǹ�2��$p<�T�l�]�*�z�)�h�A'�ܭ�/w�B���{�ʠk��-���~�|�O5�u.��aE�0�6`a�w���9"�)���xi"�36�u����dqP��Ϊ�%�,����kiн����O����E_\�@ �w��A*ǜ<�rnJM��Y]g+�+�܎���sXN�P�KDFQČ�+��v��u�:cgS�o��9gӆ����gu�7������w
^�ڨe�bR���ƴ�(83-�w��������T�J��x���+/�+�Q�9j|U8unӹCۗ;/��i7B���9쏯�}��ǹ�4 پ>36�ċ���]-O7�l;ެ�$x��kzE?8<q������r�����uǥ����T��s�U�JF\��\��`&�3�l��W�ڗ��N
]>⧅��@�k>%����%�"�~����s�0��w��\�|w]�d>�xM��.�����M���t gnP=o��p��a;Ꜭ�L�E�b�iB`b#�8�ZBp�G���@Y����}�����c�o5mϳ���g���À�q��S��[/�Ұ2O}�ՔAn Z����\�k.ae�R��
��lb���ݛ�k�%h-&Ѫ��?#P;��������䓹�Yj��4��ݕ�݉�2o��������ʹg-YZ]i�y�e�(�v#:4�~'C��;����M��)v�����Ӌ��偞���>Էć.p�K�|3�`ąm���{Ֆ�7Ɯ �C�|��4ZQ��R�%�,�(���̻tGR���y�yw�w���菦d9T������	۰t^�RU�_��FO��M���CS[��[�O.��=!swe�@����E
Û-ԇj���G��&�k�t1ۛ�����ꞌ����h�$�Rq�7�:�~�b���{�����s�?aۯ4)j�Y�*���C5����D�N�(���3��Q3��BL�"K�d�"�T�
���`ﶮ_K�'/���+!=�ۣ\�/���Q�*6!��`U,!�~]�a�g�o��hc���;�=un�W��.���s�bU����F���Ҏ�RV:u����s��A��,Te��q�������������K^W�Oa}�I6�h�f;!����δ59w�^fr���P��'��>�9��I'�nz���W.�O�]y�KN`�3T���T��@���ڥp�nU*�rޚ �\��O�ᬇE����QΦ�~�_wF)�һŦ�X��ǜ۬�+WJ�`W��^�'�z?��2@���Y��x��Yxd�ƙ�(Jq9��Wx�k��W�S|$��o����N�~�U,`/|5�� g�x��f�����tFO���C*��ut~���o� ���x0R�1<��^��|[�u�uv��<��5+�$:l��{��>ݲ�Vׂ��ѳ�JV�E��D�PZ2�r&!n/!x#ڂ���̊�
��D�I�yg���5%@d~+���׼��	�˳k�?m�b����4��r�W��{�|wW4�fq�����B#2��A���K�l��GW�^�-m����MQ�Q�(jH���?V���|�S���߅L�4��p�o^�{���#3q�9��H�4�V��L�E&�_!8�	IV1Gv����y�r���7�Cٵ���E>�nq5�<2�1/>�U��b���x<֝�	� &�gɼ�ZǮ���z:{����Ʃ�h�tD����{�J�Z�z�|)�u��MU��iZ����&�2����h�|vN���7��.�uAsRK��^���{���2���q�ew��
>�1�.��b�{q��#DB��CF(��z�x�|����T�z�ٻEL��p]#�eU	��!�;ϸ.��p���?nX,�n��'���
;|���x�)��
~	�K_�y+#E�zӯ*�6�%{�}��h������ZfB��6���6�b�1�p�&�J�v���OG��MӰ�0�:���%�Y��YtR[�2������2&7��5����r�9����K��f$E�ɮ,n���j@mn��lgA��B�f�м�C��7��L�I��8�� Q�m���Ar�iTl0�SsKU����6�:6msV�����5�l"�%�'^l�)��jlJ:���1�]�7<���vy�k[pq�������3����vи	z����Ymx!m-�ҥ�Ef#�YӘ{��"ݭ�+�ː������iI-3�L���1//f��U��>޹����?eqBŝ�^�����8Re� a�f���s��{6;����_ �K�hI��&h��F�����|�?'�
H�����μjr�a�����pr�1#mE9ϰ��M�S!�����֟5��� �㣲�dɄ���խ��C�U�=v�Ow�}����n7!z�o����T�³�/��W���8��	8�?g���>d vy��y�����%��D$�F�x*�{�J_�1>�E�c�U�@��nD�?2��K��w��{��^���R~�fZb��s���=gk0�F�N>��E�{���-a3�4�H�"e���`�+���ɶz��ƙ�����;q����ŵ�e����y�=�u�b�~�޹/X֡����d�f���B��\���O����hJ�#k8T��ᬳ�*��܇Q{M""B��g��ٔ�V��#;�z�-�փ�D�{���ח�~�Wlÿ�M6`��n�o6�~�<<x��,w��yz̧pm�	6k��on$z�֟c�Lc^5�N�thiU��(��uY^�G*�Q3mX���{=^�tC�Q(�P�,�#�;,}w�5P�a�Q�F��n���������,g�`�^��r��F�d�f�k�[T
-
�:��&`a�w|��w��xq�n���P��uݍ_�(u�A�7��)jW����o5��Ȅ�z�8b��8J��_J�7��{Y���̥Sm�Vt�1b˭+�(�*�bl�(�-.�3i{��GG5܊y��V����A:<~��yq[:oD�~i�L�ř��W�)�M+G�0�X�ea���k(�l+�lpl��8��F�U'�ڛ�u}�c�ֺ����[���Ww�:�U�a�0�z�Dѯ3~5��g�ISb،�	���H%u�C+z�]:|#)u�yU�-E/U�u!�5�����P��=U{�SUv��<`i�ȴY�¨�Jr��RF�6��8�
J���^���A��=u�P���� �]���R�������r_
j/����1��_;��K�.x-'�����wQ^����dI|˧^L��b�6�-.X-�˂ь���Vx�$1�.�xoS�I]�S����-�������N7����#�c�%1N��v���{;�}��B���������������y��g��c�<r�n@�V�d��;g��6eX�~�o �~�uY��7���y�>����t�ɎʳD�;��Lq�iz��ke���!��b�'���Y6��V�z8��=��r����1a��{W{������:����ϔ3���]���n���۾ǂ�e�O��v1�6/��~�������L��g=|�wlQ�]Vj4w��y�:��8������Lc�3����{®&/xZ����K�`&���8 ��FR�Xt���D�w�w-��[��Ͱ�0^ӵ��{��5N~r�ؐܛ>�)��ӎPsܵB�7kC���u{m��ޓ�������ʏȟqV뢝�gh��]���g��}�U�kڽ�;t�!7�䙦�*X���=��3�����p|t��99����u����y����x�۰�t�;��`Wg��<�P껃�x�����o��u��5+�iN��N��Cv�Kn�T�9��׽���{������;s�{�����2cܛ:l��ܦ79��(N�ۧ��F����ɣ�|��(��׿e��ǜ0�qy��{�F�b��n��q�Ό9k�ӧ�����o����-z���I�p�9͇�!��(5y�_�*_��O������+�?�ޭ�-_�h�����8]N��W}O!�n0Y��tG�DE=ے�����suѩ"�a_�mڒ���'e�km��>��o��ِ4$(����#97�>\�EJ]@��B�t�(���4�)���k�e�ҒL�9>�����7��1�N�߾�K���-��p�rK]e�L�X��6}J�T�fc�n1�%�봥.f���XUYngѸ܌i@�~���W�0@F�L+�	�.adHjL�.��
����ö�iZl7�u��YB�D��}fT�H҂5"n:��ں��-�.Z�=��-���f�^�w�яY�~��l�Y{;���Z��tp�b���JI��m�c�s�Ja������	*3��]�(A�������|�P��oe{�!t�(����vY��[�g�'�~����f�-H�{�X3+K��ڶp��� w��.�)�}[��M��6q�W�.��[d=�D��`6�D�K	w�5���kdz�u�
;ί�>��w=�R�[��sc����R���A��uk��{�G~?.��N�aܥn�&��e˻��xzN@w�<���!��ұ�vS�qʯM-xc������*�X����]ũH�0Z�!��7B0Q���t�̵�*;l��Y��Fk.̠:�k�j2�:���	��ys�k|�̭6v��ȼVEW�Y��~=Lq���Q��(݊=O,RA�9˶/w�[�?g�#)��	�5�����U���t,l$*�~�TRΜ�/�����j���)G�t�<�QAgN*z��fӭv��zv�D{.��bv
N	E��5�#��=h���"���	���y-�^[���61E�=JkQ�B�FWS����`аE��K����(���'	o�vMÿ��!���7s֯K65��t+j���4*��j�
�<�����9=��Q��<a�J[Q'���83@��K��ܮ-���A�v"�s|&W��_���ζ��T���>�}�Q		Z]���ORpu��IG�fQu.�c�A=�і�	��w����(B�L��VN�~�/G���+��1=K�ޛ�;n�"�K[啘C��b3]����nCgW(گk={p���ugr �83�!��{e��u�x
�')�;x0��Ɲg���P�S�\m���*�h��Io/61�n�3݄�:��:6ܪ�ɧ]�{3f��t�=�8:�`��u�\�S�y��gv���7h>�F '��f:m��x�'d�V�؅7T��4�M�½��5I��U�e+�mət7�p�ң��|��nw3��=�\�pZz"�حƈi�!e$+��-������!>x�_GQ$�<Qw341��L�[�)�{x��:M�u<56��!1!b!$qA�Z�>|_Gh_f���im4yV�)����$�(�:����|�0�$xwZ����s��^��z�)qV��j�JH�j`J9:��׊~w:�d��rb�"_�u���x�L{�rY`�ksĽ?Y9�̂�����%$�j�-ϋq������4_�f���l�ۧ��X��Ez�������R��<^1I�s/��Qk�*ջo�Z��-H��ۊ�.��
=�y������Ss\�aE2������:����Xʻ�/�Di}�ԯ?�G�S��{7Bܳ�P�Y!B9�d�&5�=���R�;t�+��4���$��Y���U@0���w��&�7.��6�)y�믳�`JX���y@�p�S,ǵ����F�FI>�ֈ]w���)�؍Q/;��[;��/��W�,��V��s܃�X��E]e�37V����ғ������b�D3{�C|��rְ�r��,��>xғj�#��,����=��/���2���F���:ؘUH��֑}y�]Y�	nϠd�V���M�Bi�W�H�3��I�򪧫��{S�:�&yq���y��{�5�����j�m�0��f]���$R'h�.�ȅ�yƅʬn���*0���Nr��7X����'�H�
c{����0�
����$VW�8Pe6a"#��빟Vz�~��[N�������'ʲR�c��x8FE&���;iƼ��UkT͟�p�U]�S�<�Gݮ�*F�!��
��&�a�udu����v1%��ںW�𛡶�6����P2�țN3J�A$�����Hu]��e��;��a�IZ�({xm~�J3�7��cvo�'A�w�4�h@�L�BN?`�ř�����!k'�u�_G'l��j��������2w�!c�U>)K�zo	2Q'/ʃ�+�Y���Z�cQ�PN&�/*��R�������F����#]�f��G��m���膵�0��謘6m�>O�p��y��(�mƗ�w����o�y`K/$������	�<����DUB`���<����&�O�7�f
��L�)�Z���"1�&
JD�F��~5�}F�����!+}�p��A���4M�x��
#H��:�G����O6��g�.u�Ir���8�
�D�$����$j�)�l��G�F1���)QE?��Ed���[��*P��<������w�A^�뫭ʋ��9Oy2�H�VH,�mˀ1��8�'�$�k�������!�
WX��h�8���`N�����TD#��1<�)�7Oݳ���8~H��w�������fVנ9�Ks���>
Rf"\.I!��i�LՍ$��(a�٩<vT�R��'�R��\O��F��'����y[��;��i��#��/]�,>���Pɵ�<��m;4xZ�����47�5�J>o[��N��*x��cA�z���w��f����}�'���- �����>�.Żr�c�[߁���蠕��dlK,w{5��?{�S�G<L�NЁ-��bަ>P�K���&'_x��6o3Q>���n&����-M��x�4��+�{�S5Ft��ٸb�n�t��~=g䆈۠�	��u�x}�گ�9���^("/��z�N���f��J�ߨ�N��/��.�@�k���(^}
����佺��q��PhQ,6Jԋ��f2F�`!���ؖۛ͘�L�a�Ll4R�Q vG3�9����v	\����H�1pd���E�s��e�n���o�ҭL������䦴���p�h�����M�����~�P7��0PuV�����8�,��LNG�_Q�/�[���>=�y��2���}W*YV�c�V �����}!f���xw;��/$M!x-yw��4��a��"=��m��׊u�|�c]pSLߗ�yĈp���%q�:�E��羣r�ɴe7u��S�('I]�8f����]ޕ}��+b��]�#�R�C�]�!�R1QQ�D�߈ܧ�ư+��'�n{9���t�q�Q��UE��u������v7��#"��t���f�r������r-��Ûd-��^���%]����X��_��V������]:��i�;U��9�*ݽ�s����j���v׹٘ړj�6	��+;L���� �uy��f�9�<��lX���e�Kc�p�\7S���]΀��˙�[��!#��X2v+�Q�@��m��qIk��I��*im�ó��v ݉�������f�#%�v`�h�l���w�^v�
y��])��D�3��K�(����g#��9հ�9d)uL�Ѫ��-�K�9�5�0�lu�d&�q���~5W�Ǝ�����\8m���tA]� ��fM�LMK�RY�1�jȤPp��QW����������3R���Դ*�e2z�r�.��X�Me�k�Cb���n�I�P��m�Ɂ��d���ʲ��:4u[�v{�z�<��^rQw�r���y�	�o��k�R�Ү6����^>�yQ������&	#I$�RGg����w���27�����m����6^��y;������]�X|]N�u|P��*y>.S��M��f��|�������a�����ׅ������ԣ�:�"�*c���E#G6���<^�]O+U�)Q}2{��Mvëj,����x��પ�E|mG��ܧƴ�����+^k�6�)�_���ema��]��[�Ex��!�iV�.�)# "Ag'IxvwI]x��ta�uʹ�k��k�d�P���Hj)�iƲ�<� ���ߥy�|�r�-.RqS����ٸ�c�hWh A;��H��� @�����-��1|�R;|$r���+y�x�[��L�w���9
:�4����왫�|$���n�u��y��v�$�qob�ݧZ���m�y[�#[�ۇ�H6���2�-N
7�tQ�?�}X�{m�ȷ����y;Hl��+�~�w4�~�Ut��.���F#Q�L26C[�"���ˡIE�F�D����ݷsn�X<Ye�-��=1
��([o���}�&�BF\���6���ho����d�$�U9�9�Ȥ��F�^��U�P���(/eh>�n���������Tv5�D7R�~�<wT��ߟՍp��c���x��Z["Y�}���Rʸ{�pVg+�Z�FU�L��ԯn+̜+�eq	����l�lR'*��ƒ�6�%`��u����6s�Y\Jn���]gx0�R[��G\���χ�/e(+��.e�7G>�Ť3^�d�z�Y�׍ft��?B�y��Z�n7���ّ�!�$��
�k�����i��~�=~��i�[9=ޫe2��/��V��R�w���uK4^�鐫��.����,�U~�	��i�І2Lq���	���`���}G(=�J��[N�cc�v�EE��7�
�M8�z��N����4�?5'��:&xw�O��	|0��nP����NV+Gq�ٱa垃����k��\�����\2ض�<�/�`fFD��$R5�V�~��ԑ�ֈ����<i���5/�V��u����E�^�u�7�*
Ͼ��~��菓�,�2�������G���S����d��wbh(�r��J7Q�Wg����s�"�
�<x�]-wyH�m�V��A0�/1"Zi�	�y%m[w<�U��C���nAp����.m/.BTf&���4AS�N�ک�WZ�ìڕKm��U;p�NN�w�V� ��w���\c[��0q@G�{�N#[�6ґ��p����DJ��ָ��_jE����{�<�Ϛ�
�$�xr��tH^�)��d����n�CVE-�J[��H8�,#�I�{۪^1�,�z���}��t�s����o�{��R�5�[3i�^��(H�f�j8�a,w��[����8�ejs������}ӻ���-+�ٳ]Tε�~uV2ic��v�C��G��}�+��oy����<��z�$Oku�.z�lҒR&�:r�{��NyK��f�ei���ز&�U^��>���s����.�k�/eT�U\�R0TF`p��X�@f}O�^���vw1�;F1=�Z[����Fv�A'X�����Q%�u�����R���0��������`� ��$��W�n0�[�#"H�h�x���t��a�'��K��;��m\�/{������}'���N9�O�H��P��Oy�5'�Xz=�f����bc��B����pͽ8}�n�ֱ�q����kb�2��n`�}��z��W�����������E��GK����|�}n�;��%|���Q�|��hE/a�}B0$��<��mS���*Ȅ�|�/j�+���Ϗe���A);-�^�<�R��I=6��ׅ��i�窲g�R*�$�Qh�:>������j�`B����k�v2:�B�9":W[�]m5~4Y��*���oί^�o�S]� O�� �L�&�
��%�׼��ޏP�g�����x�_g�`��[�_-�0t�:��{��C����4y3��e?xf��#�}�O�*K���;�ْ���~6m�����E5n'�*��u�5�r��w<ET�Mv�4����wqN]�o�*3�&�LW���7{%Q&���Sb�`�G��^����z�??ZC@EX4�����ۡo�5��'�{k`�N������
��/j��Vm�����=�J�e{z�0>-��ޝ'�����\��"|��.i�K;�ɀ�ӱyS�/rNm�&�ϪM�2���Sն���QX��H��7�U��-�T�&�t1�۱��9MZ3`3��W�g���oXC����(y����^xU�7����5B4\���yl��,���},��!��q�#�f`�Fãj�ˤ
;kJ��L3f�ո��^�i~[y�O��^i<���f����v(��K�(k[�N��2���v�D)7�YX}�*?��EVm�t�t���9�g<�qg�k�E&Ǵo����IՃt�͝f��u�ޛꍼA5��	��k�1�O��ş�o�霡�� ��C���@��d��K�����Z�i�~��^�2����s��#YFq�:����Vї�ی�g�NUSS�*��#��&-+"T�ϑ�O%���Rh/)������p�3}��/��/���'�r9c��	搨�>�~���Y���G��ȼ���3���c����L��bz���م�޺��s�}~��xQ�;�e_=��V腛=�,�3V{
O���1,�<&���M�6R�D*��ûU6:��a���b��)�5�{_-��DY����J�Y�ro�k��|�%�c�������( ��%��&����I���GnH�� sdȋ��� !��x���tnk%JG�W�YiUK�&��àK	Y����- f��;�LgPpnNq��t6y�/1+3ӧ<#/IT�t��Y�v�)�p�޽o�D#�\��K����d�ۍgcq��G�#��jĭ�3"T�T��bX�t �s����ڹ�Ck��c/Z�q�C��.���n�<`腔�����:���=]��1�l�6<lf�v���g�kպ��?-���호��=�9�.��7Z�j��u"tu)�e�l⭱t+��)�R:��5�5A�� f7۠��V2d��\�8�l4	b ��E-#u���nn��b�.�Q�a8����c���?��v��1qز���s��n�gJ�C��l{�cgQ\un��]�E��.�fS5��ܒ�(��/��mYA�1�卝��ܞ�{��㬤�iH��#Ç6
묘�:뮺�t�&Rk�Z�G�IW Dc�bޑ��/��\���6���ɱ��ɅS:�\�\v��-�x,䵟b��ǎk/O*;j�]ͮ��������5�sL+�^X���xyk��i�D� �ݴF۞Ny���H��ہ�^H�F,�(���^n����U�X���.�T��i-��81pk���qpt�[u'n��rs[���>:�p����mie[[�e�{��%�
�i�s����v�N;�m�^y1v6�`�5$��Ʌ��fɥ��r�0ȴ�]����T���,����GCB�L.�K6l�sZi��&�2�X7��F��ӧn�8�	�sVV�;	�^��).�;�������IK6vcĕI��ˈw�����8 7���g�C�re�t��۲hn�����I���ضn�]���X�ÛB�څ��<�|ܒU��tl����h��l��2�B��z�&c��GT�wZ����)���8�̜+�<��g�p�q��wQ�;7��CQ���5ai7%y��3u���C �J�m�x1���%VbV����R�!F�lm"Z�Rd��3J��gn!OnB���un� ��[&ܛ���P�>l�|���˺sj���K|%�w�1U���vk�X�Y\]6͙\IC0�&E���\cGG��7n��3�'6�Wh@+���YGEV���%�6I�A�FH���ݞ�IVocs�lpG�6n�H���)��tkuǎ#�ۛ\��]s���X
�Sp��v���Ѩs��ù	�伃}���J�T!����cF����u�U&��?����Z4}�G��[��3^⾼��`t'�[��O����cK���Vӑ�P8�q�l����$��}���>�uL��������e�np4�} +ˠ3z;AG�f�,�U�������~�N��A�	 �!��`[�V�^�����l�2_]W7�z9v5K�,���[��o7f�)�Aw���Ld��.G��3FEE
H���o=={;�Rͺ�l3�:{��Vf�m��@..�d)���:.��uؽ.��8#��"��dU}\0�m��n�������C���Bm���g��`���p�r/�͚���ƙmx8���7���Ү�����9�f�GW&P�R�US%ETdn ��:[D[R�`�a'gA�t&��Yǎ��g�v�8�� #^=�??�=��3�����^��^_ >�3������ޤ}
'o�F:<�.��vvL�I���y��:�`�a�Q���c�\l��{�����nn*��*��^��U�uJ��{{ۆ��l�����x怜�����'[���ԮÞuY��K��eB����������7;�������|z�u��6K���Cfq��}���]M�,�~&��)��Z2��o�ĸ�����K����&�+ܫ��*D#��@�<fL�˰,�a/5Q�Y��
���9�^��4Ld�ܒ9=�����ᵪ)�w(ͷ�����t9�yA`�vu�^�3��/*�T�;��O���%��^~�M����W�5�baB�R:��*ȵLve�V�LS"�
Gnc�I���^��C/$g�Z�%yu���}�]�a����{����|�Ԙ��h�*B�%�2"P��$R&�\X��K��׭'5�ru�u1.��Z�2ɍ6ཻ�v~Œ1�Uu�.VC���� }�O�(0�0�w�z��iɌC�g���2���J+�Σ���5	��p�j�h���룱�Go���*��c�HK;�%
i�e���{b�M����eҙ�^��ڲS9�2�?y�|۽L����<���z���#�hű��	~3���{�e�4���$����thX���~g:k����ȳ�<��@l��!̡g'���{'E��듌������,K��Yr�=��i�J�}���$ZF&}5��ő�d���Sd��s��q�G%
�}}���+��3�eH�YuU�<S���5�����IϝѺ�� �M�ې��_x_�ZV�N2��ۏܻn�и�W
/P��Tt��JQ�Y�:m=�^^����8��aG#�p@����~�}�b�"��/�1�wۇ��}��&�	��pw�ô�[�Ķ�� ����e�v2q�g���C�Q;;�
M�bf9��f27&����O[:�*ꩯ��޿w�uƞ+��@�u�~�o�+�[�	�U��[$xn{w�h�%��qXb1%$؅�X�G �:q��~�~;��D�#�.�_iS�wk���P���;�^��d�������ٜ���OVuv���[��BFd���R��,���/�P����u�_o�Knws�{���t�3~���	�r3}����(h�y(�z}R���E#�@礀���8k^���S��eն�����e�������n�sd��<����e�|���������;�������އґs�N-ć5�[�#}��c��l6o��7���)kܶ*��n�Ȏ���y������������S٣�Oe�4�m1$A���x�솣>!���v�6��M#:;�U��d�jis���~[<���̙�4�g]Նn!n�#B����M��<�S6�(���I�ź<�Z'��R�d���-��j�t�S�ٛ�=u�������I�O{˹;�Q��ܜ�ӑS�PVa��7F,>���'昳�5�.&")��qZ��\��í�
uH��"f���=;R�4͂�4ZOzu#fٹ9��]��0��/���0٫��W;͓nǽ�Xh�*8�8r�j4�!����A��s|y�p�O��c?|]$��L�O�X��G��n���U��,tA��1"R,~�?M�8��OR����j{İ���E|��-��mv#Y�6|�EC�Lx�X!.��{~���g��=�~�ͲJ�ؗ�{��v�������ڛ���ʗ�������K�����D�����^򒦛7}�Dj�n<��=qp2���O��E��	�古��c���Ϻr����Zc*ڛ)ў���{��X�����E�7{�i�5Os�v=A��@��m�L�.ݩ�tE�F������n�i.7m�殐3WR`��g8�j-�x<SJb٦�X�u"�1t�`���Y��Ջh�W�k��ٛ�Y�"h��k�܃Krv���ϧ�w=t=�78�����˱��p�!���:�{�F��s΢۲�a�ؤ�T�3�=�Xݨ�9Ln��֎t��d�+��Bf�[�m�
�I��\�k�2r��͵�$zl���;p����m������u���(��4˳f
���mz9ׇ�Fn����(ܐSf��;�`���!��oI�nu�5�Ā����,�!�d^�|E���~q4Ԏ&L*Hp��d��k۽��g��#3w�ݷj�����n��J��Uvh�+�����}������Tj����IO��6��u����#6��ao~s�ӇB�����Ī~���`k�;�<Q�ձ�Ղk�&I�NNm��}���5�Xwg�^О{�=���vX]�v5m�g_M�O�{�o��0l3���rVQ� �%'�1]O4t��ض�Æ�J��s��}4l�G
=r�[�|H)�>()���.�Mtu�k1�� �)�k�y��^�y�j笽�D�s:DP<Y'��*̺�U��2��޼�mVN.��7`����l;��q�dύ��>����QhJ�٥�b��Lbi��Ԍu�Tp1���q	}�_t6���#�;�U�E�q��f��|���ː��`�x9�W��Qӣ��y��z��39]�geA��� w�w���9�L^Y�{���J��{W��n0n��O+#�׺�]y�~��>OΉ�	�ڴ��i�x>����ݠ�KI}�����nz`gb����ȱpȽ/�ӷ�sT��<|?59�<�t���ب��u����l%F�>�j��ӎ�	
���)'r$)(���V�<80YqHB��;W�3P|���y�\�d���(���<y��2U`�_��Hpu.7�����Mž������#čy��V���;��"i�����K=���,�Dk�k@�����4Ʃ�-�'�#`gy��&�Оx�����쥚��Ob�4JC:<ˈ��ٷꁵA!˺��?yG����v6��ў�z����������:�p�і�+s
S2�U���F;Bշ��%�t]l�E�週�ځ&�U��1&IT~�Ί��!+��4���j�a�w��i���!X.�wh�ϵƏ�S��38���G��<� �rD�fH�p㎩�K����'$�o�g$�0�\+�]�|�,��I��]�����9��>�>�M�9�L4�L�B17�F��*�U`�g�D�T}{�k�O7#m��ЙZ�h�C}�*�
�z����{��|a%�7N)��o���Јu[��ѓaߴ�=D]T�N{{޻��)=�^"b.�����tL:KsW��aFڒ�n"�SO�!���v�oH�����'nI3�}��������k|���(R�gV���[^y�fh��r�:t<�b�n|�M�!� �!8�{�)]uUS���l=7���]��U��vt2�)-�J����%;�e1�]���{��i���ق���u"{}v�^���2����$b�\8��iQ0��%X1��,�c�V�����%����<���Js�+]nz(G2�B����>�	�ze_���z]FwJO�~&��
�O����*����.�T�/��|��s̴�-���p'��������VWzN��]XUt���K���x�,��kI+rȥu����y��ƪS2�sr��{zZ�@ׯ���?��1�&l�Q�8��"Z���Ӷ��
>�W$�^�������P#t��s	"�P"�
�7����uj�r��֡�?3��������I��X������Y6i>�6��`����d/��(�L���������픋�� �=L�\�׳C$���N�j���B���7�{s���ڼR�e6M���x��?��0p �<�� W~[P:�w?E��*���$=�W�m���R�v�^b��{]��#7�'g:���t��dq>�������^���e��	�72�93[�IwW.� �s���ΰ`-��9.ȥ�w��ӓq*G��<��Yi���(�e����>�f,_���}��g�S�/����߲׶ꢛu�לk=����	���j!�B�N	JGY}q"�]��_�L�L愿3U{U�9{�Ԓf���6�y��JE/"�k�7U6n���[ׄ��#����O��.��k+"d[�^��uU·yׅ�ˡ���
���m���WJ_�?�;�KA�@�i8�E8ݜ,���Y��9���o;���<�q�2�{��F2 ��Z�_<�լ5׀��_Q��r/dN�y1 H����a8�-��A&���ɧ�<>���E^����-�u�,��!���;et��z�9�V��z'7ñ{<�;�|jƵ'e���xD��<�(�5����^��u���_���OmZZ�Aƻ�3%YY�v�U�6Q���m9h3!l�۬��:��9��
?T����Kb$�Lj�p(�t�e��X6h�QU�W���f��\���ԭ���Դĕll�G@��s2��Z��H8�Z�4��;;E�۝WK����ؖ3��Kf�]R��G�
j�����5Ț�m�7���#�����6��@�h����Eخ�J�����⢴xAVʇBtgm	�Nl':����0<q&bُln��b����"��MR�@!��i��Upݬ�$�y�}����wnﾷެ\���|wO}��݂� yϡ�<�-�|&@�c[M�]RW�q�x�An�U��"��F&�jG��s§��i;Y����-O��'�Dm�//�a�{m��u˫lM:G��P,��1>˥�A�W�o-�}�4j�j@�jD�R7�.�l��5Gܾ�L��kՋ1��!�ly!�n��#�Lγ|��U��v�r>c,l����}�r����)ז��O�9�yT����_��`����΅�w2d;y�"E�z{�f�y�u������Z���T�$�E�d�7ܤ�z�R���Ym����랽vo�Lgh�w⾓W�l{|�P����ū��X�_�H��vΤ�_���
�~�L��&�L�ӈw���,�n��G
�ɫ��R�\d{vV�T	ǅu�۴���YQnr�{�:�ӯ����ﴞ=�xG����������"&'�$���ҶLڰkVl]3c����K�A��Y�Q,\;���Kx�/�?}��^ܛ�kZ�߮ߘ�����<��t��G�9��o���N�]�к�8�{�v(��9b�$�P�k�|��gv)�1�w�w��R�<�B���W���}v{���E��	�>�)U^�ћ�Q�#n`Q*8���qz��(����wݒ�G<z�<���W��,��}ZP�t���ݔv��Ӌ�*_cL���x�����RH�p����y�>��o
º`���{���?xW���Mz1���nZH�I���l��!|M���oОs�{D���Ɏ�!$wGoť$1ȋRr��Ӌ�{o��~*ȣRᕏ|ݥ���q)b-c�w'b�o�R];�bkT��DU80o�FY��}w���X�-�&�Qx"x=O;�vx���Hݻ�l�֗�ĉF�ܙ�0�0`�����I�m�?O_�N��xxʗ��}�����׊�n�ʐ���Uה��S˸+��R��P�!��e|ۋ��$��J^j��Ϯ�e���>L�Piwt^{�c�B����䫙�3������������0^Ep�~��ޟ��f�h��JE"Q1�(��>M���S��oH5*����<��[��)c+y9���Ue]<]ڲ��F�?Q�v�}�Uy+R�LU_�6��6회��uG��Pw��^Qջ�?Y�~�'<�0����Cdv�ɒ�ۜ�(%��d�ېs�a��}���夢��R�Ź���_{��&��=��Iy����'��:��dI�bۮ�^���S鯡,�Z���������6��ޞ,GU���^˂u+��w���?�Rxt��3��ָ��Z�@�=˻7
(>�2g^>�@8�n���YҸ�qgyn��/<�^ǔ,����jzq���th��l��7�O�{���Sٺ��C�K�����{��u(|=K�D{�o�G�sh��dk��彾�1FYl��x�� �*��dI��Е��[6��1�r۹Y6z��f�i�Gxn�L�%G/	���bk��z��׭�"j#p3Iy뎴z�rѕ4x���h�˕��{R�u�3�;}�P҃.Y%-����d���0.=���)�%c��i��R[���� <=�k=������,l��
y?�ws|���5<��א� X^֚>I��̭�A����;���ioW���X�Z#��דW�z��Oğ{�n{u$df�(Ȧ{;i�|��=���^!���E��J�!�~c�vmb�� ���;/�����{xo���w�N������׾�>~����ԧ{�,�[?��}����4���ȍ.�F����6�A�X��o�CJ
�ݧq�P�漍��~߾�_{>p�i�T���}�&]��>���%�#��K6*�דּ90��&������ϰ��z��\!������k_�߭���w���
��47�Ӟc��� st�T��ys�s������9�	�n��H9��:��?����Ϯ��X>����n=p䝅-o�g��IH��^G)��=\[�'m�g�C]�PR*�YB0�	A(�4Bkcr�\�J��ߧ��d��Ϟo{�s�:�sݲ���S���"{����nw��!YȾ�8 �O�ٛ�Hb�y%5��_1r�Q�|ļ9\�_gl�����O3վT�j\3}�ם�C��:�+��l���.����w��-����jh��ƖU���k�K��'a8 AH�$��0�{����2_`��o}��~��k�����+���9A���Ԫ�����^�9o���ʢ\�DJ���;��u��v�z`�MO]*���w�{�9ܖEusR�$#HE'�z[�|C�\�e!!K%���|�g-w��{Ӷ�/��Hݞ���m��C�ۼK�<���=�ȕ��zg�o��;<a��u��Ѯ�>�w�Y2$}cЬL��Lm�{��r)uK�y�TI�"�����2�L}�_�c>n�4���W�d�T`�HoVy�0��d�=f��{�
^	�K>-g]�չ��/l��M�!�U�[gZ����fmД`,ua��V~B�D��/o?f��"�߹E��yx����u*�ѿx澾���4G�X�rt|�u~�*пU���	r��8$�P9#��+(�r�"�u]w=X}�gx-'�ܛ۾�1�zڢ$J};���g��\h;޹k0��d���j�8d�Mu�ݧ�}q�
d�"R�4����}��!�I��z�c~��]n��0N�36t���oU%ꦽ��*ߔ%U�{���%91��7�=ࣛ���B��k�+-M9	�~�t6��G�N����.{s�op�cO��w�<��2T���8�KPA݀�G��	�[��W��_a��H����i.��w�r��O9ƪ���Ǟyu Boc�EK[�z����I�罼��y���q�ƲIS�{��fׅj���)������i���y�H�fx9�y�j9���cܵi� �r��1������,K��M p���9#]���.�v����X�h�n��jܨ�T��a\�WYVP�.���MC��ӭBn��
F����*���P�ȅ[���#��d��ps�/\6,d��k �j�,^m��k���ׇ,[�ر���A��qB�<�㰽I��gNܯ\Nl��MuN�GWY��^N��Ǳ���j�'�W<[d��.kU�ό���}%�;Y.q���ƩK�ۚj�$)7�B;JU�]�C�^$5j���"�7��1�'~���Y�ƈ؝#�W�/��
)�Φ߽����F����5}�GW���ʐQ4�r��$�CQ�$,�2#������W��S��ծ��Ld�½<�p558~��WNw�FuJ����â�l^���5����ˈ2�i9�c����,��r��f|T���﹅��m>��wO*��� :ƨ��%v��!z
�"z��=���V��+s����$�%��`�$ǅ�Dü�n�UKۘf;Y:u�y"u��Y�����q�3sJWؚ{	��]�}�xH��`��y������U�(�-D�fB$�G�ҽf_)�|���̔���z�(����q�	e
�V�<��瞧[��ۮ�ޑ�f�����^}���D�$%���p����W���WKt�v�h���A�O������AȊ1D�]�b�R�#nj���uDf,�!?�y��ɟ$���_N���מ?������?<�Yg��[�\�(_x{
2ѐ��e�!��K�+e����?�_�����ԹhX������;w�X��G8�Y�\�FO$��m\Z�r��<�����pv�x�x{+��{-M�>��6,��f㤔1t�,Xo�vƙ<���	���Ÿ	r����/g�3���<'ȵ�ݜ����ԒB���˒8s��U'�:;��=y�^��W#���oTi^�{�>� �
���]|�z�.�t*W?P�Vܝ�hUr9�E
��T����?}�]y�qUg���G�TL���c���\I-��+�C��R��K7��/{g��]�墳K�H�Xޜ#aF��R86a�����%�]
td}���_����ǲ1�@'E�����ϗ������K+s9���1M�I�F2� &�h�e50��"i�'�۰p��!���,��ؙ��Wl0��.���|{=����g:��Q��%�sӺe�A�s�AΎ}~k7}.����_{&����Qy}����%1�i����Q�>��!P|��zvqφ���h>��~.����0}��.��+o��Z��~��c&���u���ǹb��A���QO`��!�\����Ӿ��t���s�FӇ�Ǆ�o�g+��i�̜c2�}�h����5�9��d�Y����Y:��^��řN�Z�L$^%��G5}�}9�
���6N��F����������	�cx������;�}�v+�}��x+��h����b~Qm=5�l��h�P[��yt���ls8qN�f�;r��rV�M�G�I.�z�a�\(w��0/t��P���2�o�
2[�+�B����l
�ͩ��2#��V�DZ��(=O5�3=�y[��N"�<C�֯�8=������w���:�	�
k*�gCMI�2Tv3q۝2$�sq�rj������5�N.��ep��8���z���������̫�ޤ�XA*%�'��ذSO�����/���Nx:��-F��+�4�m�V��D�����rIS�5�n�Ղ.����칔ܺ	h�~�+8) i�}�`"TJm�|O�-g�l��(+��~�)z0F�ܑ�*�t�&zoy�f�:�8��_;B���KA�zﶝ��Է���a���5(�����~Y2��]�A�D�1$D�#�߁�#wظ����>��fz����sWHO^�!K"�́�w6%��y�$��u�:�)�B�؊���(i�~���c'�ñ�g��t5����d�?_a�4ۜ>I�25����~��;d&)�`�_���:�V=�X�ɲ�\����1D#JG^��Un���zP�3s�K�{�����\�T�՝oM����Z�w��~��p�b�`�Y�}���n��$pkh��/M��Vf�]r0��`�Bb��E�����h�ī^Up���we]�v�L�%X&G��oi�OX����ڎ�*̇���"s:�ᱽ�@��_m_y��77�O�PV2C%��Q���>�v���������4MÎ��H�'�����[}*��۬P�V��^}`�<�NjX�b�Wтw�q �EG��O�~Ν����-=dǛUӝ~��U����]-'����G�帶n�M�_`�s}{�>˒9�A�N���r�y�q���^�k�o:�lS�WϬ!�h��i�[����*-�^��qX�֪^z/g�Vg���^����	N"�e����tY��Ti���ӆBH��+�}V�#�~���Ԧ�|�����?7�H&��c���n���^n�J�Ķ:�q�Z��7��?Q��<�~Nx?� ��ޞ>؊�Ɩ�}��y,�y#�ro��M����Z��y��ZJ��@��ID�r9#�;<,ل-�iB]h��h7,�& �l�Y6�s�=���i�OdA�]�Xh9ф]J�۠)�;����`�^ח9��*E���)6%�`�膺jT�fdZ2��:��+7SD�s��9�iU*�Ⲙ�0�i����DK����FE5��N�Ks�M]���q8���l#0�"����;o[g���;-�g��N�䎷9�<����]�&"q�i�����0+��"�f����u������u��X�p��y������N����[���!�p8���>�b6د��Y�}O�sj�,�`.�y/�o�\����G�7���<(n�&z�g6q�dƕ�!����u�^U�����/u�ܯS��H�ꅮ�+��y�QJ{�Q�&_�2̑���yN���}ҟ[e��1ӆ���zz:�{7�xϷ��S�2��?{�h"|Ϡx��T����d�#Q������6�6�����>s8���/��Hoq�^�^Č�g�	�u�X�+��e��>��o��
�Юđ2B��$I�'�]U�k����]>����4�⟯e`����ԻuPUnt��{E�A�I��Z�O�|��2}�ߗ�f����|�:�ѧtm��zډ�s�WnI�=�\)b*85��U�9���{�X_Oo �9��}�w��g�7^o/�;�x�Q�y�{�H�%-oP�h�?~ӿ|T�u��ό�4�U�8��P��#���鞠sM�^���ѓB9b�����,�#�1b��Е=Ҿm������	�fQ���v%�кt�q�ь-��I�۴{C�7x�ɰ�H��Y_Ff�q0׌�menu��Qzx��́9��*�����E}���}�|a��dH�nI�)D�״�iw�]���,���w?x�%��F�=�굺&�:��0?$�OBߺ��xͅ�ٞ���֎������ ͕'���ٗ��
W�����f�؝-�;��m�oK��z��w�#z�@����7�b��-h�Ħ�*c�#$[���I��N��$�ժF+����}ֆ��O/c�^�����I�����yx;�^ץf�]�;f|D��h��a�X��	f�XP �q6��ϋ����.gy:3�� Tn��.3�
?�����0�;��k��>ƚ��6o�p�ԼQ�u�������q>�ڕs�$}�Eu���q�?w�%�es��=~�Ņ>�x�
��Df׻��yu6�V���1ud
��+��(h�^���ϽT��}ߞl�p-׍�N�����G�+qV��N�$e#8��a�ǰ㝝뷼��{�R���Vy,�,��-vڷ�c���)�_��-�϶�) �{�V}��޺h��Iȵf;/��)���V`��-�lμ�m�n�)�ێ�͞R:N���z�Q�}=�w���Ǉ�Nϔ�9���"��s�|%�ż'�=��~9����o�.��+����rG�K7���1(��Ԓ:�q�/%v�_�*3|.u��5 ��?O�.{U^7�{^�z��2_\���m#�4-w�i���u���P"�%���8@�\p��U���<%[�eUl3��bV<C���&Z�"b�8���ak��qŐ��|��j��;^voNX��{�/<�ˍ�ex }#0��ǧT�h���dϠN�pT��;*���s�z�,��UǹCV�8*I�2�K���d�of��������}`-zG��-��,�ϳ�!ky�n�-Dd�q�{�"�&}n��Y}uU�J��Os�hOb]�T��h�u*�X]ۤ�Oy�O䚚�D4vu"�$�r:��!�y�hK5d�X���{�6�O��\�ȼس�]�ET����{>�e��`�U����n�����y�2�Jf�U��
.���י�&�oŧ��%���jǩb6��~��kOOϵh�{�e�M8+�_��_T	����y�e_�H�����O6���sy��r�r8�J#^��5WƱi��E_���Ro<۷�<M2]I+y�����6�53�X��*��C�Y>��~����_�͊Y�g�Σ5K�{N	��s������l���
�⮒��Yp�$�Hbέ�
�t�r���眵*�u�I�r��o�'��U��=�+;�{�φ�	«w~ ��+ ���p�>>�U�t٣�=?c�f��~���Y�p�=�����2W������Z�]z���D
˝�(�]c���^>1�|PC�{��p����)B@Df$we&�L���MHn���bӵ�{ϔ:ȫ��4�����в�([����)����ſ||i�<f8�D�`MdW$3�^�ؓ��$�ƺk�3�}o͌�ˋ~���{F.z�`3��~�G=~dޱ�>�����G]r#���� &I�±q2�ЯS��毰y�:��W5]�^5�X�w�{Iպ·��JR����7���\Wϝ��b�Y�d	��]"�%�u�}X��ߋ��}��9���뾻��zj���,�|׉T�h��]#�C���R�S=�^��{z/{��2[�e�,�`�{r��߶��(?i��$P�<��[��Ԝ�U��pUYZj�*�E����Տ{�qe��)G�[��_���=���n����oҋ�z�a>��a���e�1|���;��dy���\�<<�_{exygg���m>���W��l{(WS�[G7���3}l�-����k^vok6Q��������]�IG3���§�F�~�9�4�3n�f��<xW�k+���������Z�B1�Vʞ��(ί������D�)[瞾[����zO5��p
����|dܩ�Y��}�Lh��zf��9�7��D�����.��?c�}q`�����!`鍛��^!��9�x�ׁ����Y�vn�������ǰ�3��@o�QM5�����.7� ܻ;���U{��v�0�f�7��/ �^yAsw_�5�^qw{�9q��qT��b�w��Z�U�K���:fO����s�w��rsǿ_qM���u��+9���|�I�]�ǽ�R����R�O`WGEc�t����|��$#���s����q�M?��?a�>�����$�%c0�R�������q���l'���s��hp��Wtc^g���<{������n٣��7Ǟx���Y�����22�<���R������c�]�=���O`_,z�&9�ڳS�)�-z��`�Q�ߢ�`^�J��x��d��w8X��&s��z�;unN�8�I ��sS:�N��!�;�&���H��k8�K��;�7]j��քK��.���[)FU#a�n�nJ�L�٬��pZ��(ٗܜ�GZB��6�v3$�%[D��#���qރ�Zin-*�\�<B*񆺬v��������x��C͎��u���@�\OZ�{7(���<7q�
�ax��Rl;r�؈��i�j7=��l����燗��F�r��m�/����1�R��v��2��* �mnf�k���ε���ڃ2U�ư��y�CY����37LFee3�Z9��k����۠Tۆ�n�u��2�0�,α�Б��7W�B@c������B� Ke��Y�­�NU!F�tqې���G�mqasR��e3��l�xz�;([{��n�t��a�E��'�!`��^��<܋:mZ��5�9:������vx޳�ޠ4�^p׵j21ʯg���y>9筫�a���,9�n�]X�Z7�1-R��-i�I���:���ZpY����v�*�iL����ӛ��<��6�vtk223d���a��i�8�U9�HH�n8�^0M�6��k���X��aR�@��,Z���ї�W�����y&0v�r7�y�<Çs���ع��h�2���n0kvݝ5X�k{$�'*��Q�����mT�ת�������ϱ��B��t\�+4ڛ@�"ml���m����`��7ʌ��m�Z�}��	e��d�,���
Kw)��P��ڶ����cH�Gj�g4�fY�+t��"ǖ���vn����̍#���[hN���,ы�b��ц��qʊ�7l�����3뱊�`S��5aNL�9�q�k�P"%�B3J�������r�{)��b�;<��$�$��&���.#�;���Su�-�=�����=bd^�OX�Y3�8�ck%�r�m�����\��,2�QfݯXr��n�;�)�V4���n\<�ۯS�۝[�s-�͗�]�GX+�v��۝��
j���=����vN�z�5e�c�ժ�ѫO\�On+n#`���ǳ+{N��ݺ�<,�z4m���h]��+c;=�Z����6���f�b²���R�K�F�t3.�1s0M��7&�#ŠK$���tIr�J*��[�+�Z���fe5J��FT���3Y@�c�U��V����q�k��݀w/�<�t�x�܏�q���t��!����j[�3V��0 L�	7m�Ӣ�=e���E�Z��K22�K���
J�����~$��)9;�Z�
���T*8&��ٵdh�Br�e���1�{�};
j��Y��`�0��8.s��k {{�����Y�}�>���P%��Q&�ɾ�TC�>2�|�2(Za��Q����R���H�"�2���.u��V-"�R)������O�_�������w�+ދ!��_f;�훅��
��D���R�0A�i����-4 ^T�Ӑ�*"��+�}7�[@o&ma��>�^GN��1�ې��=����e���1\���/����>��p�p��y��iM1*)����3�}9�p������$��J��vȴ�y7���^,�9ܞ����E�P��j@:��y�,�����p�.�h���'W���d�~��:���ԙ*��/������	x����=�*)i�&�}�|�9 E��%'xүg����� +:&*��]}��
�ي�qƉ_����V�{cy>{���fl��g�;�O�n>���SL����s�_�it��qB[��3���}a�����s�����⿃{��1�k�bRYo��qb^�6���=}B�%t;,S�>s�y✙����0����8]��+�mtɧM,S�d��SU�W�os�ڽ����tr�c,�[���h9���
JJ�1I����ȧ�:������N�TxT*�6���Z��t_+!Q	�>wM�߫8�$ZB�=֮�+8t����xC��]����]�c��];����E��)�Oғ#v�Y� �o��S.�U:tL�L�UY���g��0��H���(��~�p�/�eO̮sj�~�a�/I��pJ�E뾥�=��sx�4_._��m�q�7G��4�{��P:�+{U�������y�s}�sf�j��3�7W�_)p�L���G���x@w��K��H�&V
ЂO�ʤ��{z�)���d�tq
��a}�}V��ڎ��3�_~����о��EK���]��;v�;C(g|o������K{?	b�U�����7�#�W��L����B�������k�f�q��_+��{�j_�EH����'���y[�pROZM���#�r�Y��,��Y�K�?g~]깕3.�L)S�����Ǆ��l�!^7���l�J��__��__�
I:O~�U�4��d��XG���^Wj+>��Y����w8�k�R�M*���tZ9j���9���?����K�P�����d�X�g���d)����E�m����'ϐ��8���E)*�d+�Rt�����@��;���qgN�&�/��b��w鿍���;�ٞ�RI�Y
�C����fI�'�*"T�D�1W�����i��w���1�-��T�uU{�r�׺�L�����Z��D�!j�O�15ف��e�:9n��R�V���T[U�mb8J��,!2%��&*���c�ZB�i�.�|+>'���7�B�<
����ps����}�O�kl��g/�Xp���0K�U��g���ӂ`-��N"�$�5d+���US)Ӫ�7T:�p樅Fu�Y�p�s�;��:.=�����ܭN�O0�M{�b����ss�¬N�ϓ��q�hSJ��{V�/�zD�ϯf�	r�m�����֞]�����}YE׾��!������:����Fh ��ԟ���T��l
<D��b���j�����1r�cde����~��kE�}y�Z�<Q��>Ѱ.�C���|�U�E\����6~�ai����ײ\�<�w��L����wHw��#�p�9�(@�E-��Y�T�O![ ۛN�^+
e��`%�L�<�f��	��������Z��\�:)R�U@@��M��2�������I����,�GN�j����}W>��IdX��1B�y��s��q�W0��Y�0J�E^���M�53+��"�u�VᛟrE�ɫU�h�����_8�!-$��֟v��`���f[U�wy����v�a@-B��=u�a�� �IBߌ�-�g���Ҕ鵐�|�~���e�Eg���7{IV�V�i���!Q������sφ���{X�F���,~ƕ��Q�^�}�]�=���]URMLu9�u�n�8��f�te�p�2����r&���n��a
��X����Yl�����֓�f�рa��{ϝ�NĊĬ�E
�S�۫!|�1��,��q��r���ߵޟ�A~o�֞I�g�7��!�,_{�昼G�xx^=��Y���l�7}�&�n$�Q�Rq��:��[,�FWe`�\+���p�^˿������;y��E'�ғ�S�z�a]�(Sn$RC.���iN'm�������ϓk/U���������_er}뙵�~������}��:�M&�n"�uU9�cm�
N�@��;�b���ڸ෎����UD���
hn���'�H�Q{<�ZG��M�\�Ĺs�D1IB[mt\�N��}�+VpB֤D"\b�ʱ-'������U(ML�T�-#y��H�~Ɵ��U�R�bc��>�Xaf���+�&EA?n{�{ϟzV�#^
Ed�*:�ib����ό��XT��ԁ~=����YؚP��^i���=n���p�^�1�����G�
�����n���{�ZAW��ۺ���{��hcu�w�:%7����4�]�T`8RB�[��샲�ĳ+�w7��K?]z���V`��?���m� ֝Oi�����|W�~ɚ�2��#�)�|���Z|t��ª}�����\���\�Z�X՞�Җ�%�Zm���=s�>8Si����7t�����^�ֻ�gh	Y(rpD���t�qe\��[-����8�w�����2Z<��˫�6������/�ݕ�p�N̈��$O~櫋ƴ|�1��0�W�fEu�������ؘɧ"�v� �v��T'���]*jϾ{�b��%V��熉�o�,#����F��������{����Ĉ��SK��GE&������i r_ں�ϫ#�}�[wS�ئ~|�t^!�UG²y���h��(�&Y�Y�ό�;�
D:��LK��b>�u\��^�u?��ל�2�1��f���l�~牥PG#E�rX�}^��N�"M8IBy�Ӫ���aGq�X�"嵴�}�s��G��ۅ�}�8.?J%�^��#£�\����6cᐬw2�*#���Vn��d..�M�vF�[�}��}������j����Z/L��V�K�t���ז�Q���r�xg����f0��iiB�L�����p]��VBt�M��Ϫ�Q!s�+H�+y�+�O׾^p�s�-p]8GP�RĬ�B�{���1̷.ij���=K�d��e�n��|Y7�������?�k�i��d���w��z����Ͻ���K�}�\<-��֐c5��ߧ�-,��*!2(��dĊk��ˎ
H�ܞ�7f�!
��D�����'��.�P��.���h���z��P�_�u��Ź����#�N99�u
�-y�ɞu?�=�ﴝ�g��8U��н����ζz��0$������º]5Ʃ��+�u�<��V���B=�K>4�]�US�1�mmܝ���;�w;�v^��N���]�/+��He�od����;M�d"�,�\Q
�.��Ǻa<s�C��6�.��q�wm����q��Ee8�	�^�uh�	��vn��#�#��cu�uD��m�u���a��u�9����հ�%�ѻ���Ɩf�mm�;vt��[oEb9�tgU��C�y�	���q�VJ9k��-�.�iO�N�<���,Y' ��dg���h�pTtL�52�b�H���j��3�²ĎT�w��FM�ƀ�~�z���*����#ㆭQ��),E�ܛ[�S���E����I�������n�Й�E��}���H��RC��	�e��],K����K韾禜{�4�� ��Yfz��~�p���|����tY ��]��m��!���/��m����_Z�>_J��/�H��x$�穹�v��p�gr}|�����������1,o~�}��Z.u�e�Oy�\`�����qb�A¢$�2>�c�ί�xE�E�^۲+'����)!��-{30�謅��V[$�)��o�N�(NA�F��)��cR���I�����<K�k�w��n��;�����}ܵ���SN>�cȲu�Zf����]!l�w�V,B[�������Y��ܴ�oݛB�e�����)#[RD��]���A�Ce�O����14�K3��}�\.��I�>,�B~�/}/�0�w��N��>+�VX�vU�$[���.�nn8�"G>��,W~����m�����_��Z{v�j�z�^��5��њ�ِ��Iq*��RY�VVۓX�p]Kv�!��h�̪�?���ڙV%$��%h���*�ZXkh�S�ۅ���Z-4W��<�|'�LYm\�N��O�{����d��勧�8�"�
N�M��7��1ol�R�Ƕ7�<gN��?n���1A��,��+��yU�LcJLc�>�E�����k�t^�>��]�n��&�UI�/$��#^Z���2~�O���Y�Vv�A�W�h�<����풍�u�=�wK���W9ǩ�=Y3��G�p��-(U��uڲ9��M8���.���s('���N%Z�pJ�e��Y�"b}�Yn��B��ܾ�D�����$B�	��3����2�3�E�rw[7�,ח��v��]��w����d�϶��N*ɍ���z%δ�Dgw:z~�U�S�ZB�rL�*<{��+��/K�߳�8Bw�ms�1�]�e�)�@J>�I߸j}�1�r�*T�f�%g�����0�S�ڐ	˥�����7߻�,�y}�y.��Z��Vԑ�5\h����-£D����K�1I�)	}�F�~~fr�4������O&D�F��to;�������KY�3P�w<�����N�a`�uJ�Ym�^s�f�bRpCa�M�}�J�,[�߶�;��}��/�f��KL,J�%&B�7�~�qP��k�Of$Y��2��y�0�.�Ϧ�N�+w)Q'�|�S-�~�?�?_�8��GK��1�n�������eR����f
�G��aef�5����m�Z±�(���%�)#�R�[_���f��7��-־����)�r�P��
�}ʵ�w��d*)$˯�ٴ��<3�_����"���Id��O\򘤎�7�Ԉ7\�p�N;��}���Rܧ.�S��L�;ZF���*�	X�Z?g>v�cz�z����Nl1Y�&0X*B�7�p��&��"�ϔă����8B����c�38�B���v�\9��oof�?wp;��ETՊ�2�-���A�1�Mw}_l��cyնIH�;�e�����it��*�#��˙������w
�ִ����^��}�/k��.x�� x���n��qj��m�ހr����Wo[�<�~�}�6J��pG�[�}&'
2o����x����)��x�c������Ҿ����\�یK쿸�Gfy��ҫ��6O������!�<A럾Ӥm�+"�W�~����}''徯�јEs�w�8%�I	�b�I�~��-֬�!��M�
Γ.պ#�_k�������.&��z>���+g�#���\����Ŷ�X�ܩ9�J�4S����r扡�
����-#<��\#��b�;���`�p�&Aa,Ɣ�"�~��?^=��KX1o_��3{�f��������6�'�����X,"ϊ�R�u���gjH�E�	a��LRAG{���N��~�����{P�v�Ja�7h�d"CKͭH���6ҪP�c�4ke�ݍ��eR�`h���*��s
m�Z4T����ѝ���E�"^�P��n&v��aW)4V�S�
��ϼ������9~�>�|B��EE��E��|���[�<BY�E߸����uSg6]L�F31��g�����K�K%�I������h��C���U���/�+$���NU��;��p��
HL��TH���ߞirBە�`���
d��Z�8���w'��^^�Ͻ�H���X������tۨ*FM:���q�>��KH��ȡ�ґ϶x�aYϮcGW-2(\�v��\��%��\��Y��΢k�S�!p����W�y�����(�!]��:!gr���ER���p�Vn5eR�塚7��k�	�u'��Mn{6rĬ�5>q��82>9�����ò�Ӌ�~0�ȱ}\����k�5$H������{=��$��TV��|#�f���=�M�r��ߡ���3��Uѫ���Û���Z�zd1��{�Wܮ��{S�I5_j�Ƒ\.����.�����>s&On�Y�1�1Q�z�yyz��,������0n�3T�u�-���8����yǐ�/�J�[���L*$s_t����<r*jY��=M_2zx��2�y�O��-U�WHZSiH��<%뿹6���h��k�Y���S0���{��?����ݴЁ,YMxC�\�5��7)v��[�v�t�US�u�V�щqjm0��r}��@H�s�a�=�3��&���t
:�R}W0��޾�w����
����2��r�E��?k����^��>�O+�%%�u�bU4�E���x�r���������/'�����j	�A�"y����I���g+e+"O^���Vr�^��^Ǳ�G�h"����g!5����%
��sڐ��>.��޲�)�m��q��NY�w��.�'��jK2^�5ό�x��+�t���S?}�J�I&JT2�J�w�޸TO�5�5��ZO_�ٿ�pS��{j��R�s��tN�TG�j�՚���d,1���fo�kE�>	�g�Yb	7/���ڢ7Z�"ϳk���>�G��~�XԒ�Tܪ��������iV޾{��_W��Z�\�t�\ ���*����}6�A\�E
|�e�"m�+���.M!?`���Ŵ&$~{�߿V���Ϝ,��\�����<���LZ���7 �LR:�Ո9���m+'�p��P��ݛ���D�O�R��}:cwݱO0���yم�p|��bU�e�dt�["������{!O>��� -7�{S�,"��m`w��>�ﾣU�?��	��`n�`�q���oW��tj�vAw����tx�̢���F;9��� ��y{.l�՛����c~UK��lG�z��t�;ih�c<c���4vԹ{1/e�a�j�>��j�����tu�ݡ��_Od�o"gp�򽞻�=��e��-�^0Edɳ�h�3hO.���r�r�g����c6x��0�����+7���Ӡض����u�ҽFu&�r/��;��åJ�R�@�nYv���T���1 ����.$\�a��ݡ�a�M�Ř̜��x5����an����]�]�xy�b-���mU>����I�j�3���)�oKR&`��cmċ{�
����;����E��y���ë����;��is����;9����߂�%${�;3��N}�M����']�k��sz���4�����P�f���;��;i�-�|%d/�w��O�ߗ�=��no���!ؗ��
�Og =�y݉i
�Bg�Ϫ����!x��$��� �bd����X���T�`�����]���+>[�{���  �D���{�~	�� �ot�1�������&M8�\�&m}��T�E�p�������ܾ��F�p�GD�����DR]4�s)���{����pI�̕�^8D-�߳����R�1�c���_�����8�t��ֱ��Z]3'�����$�H��0��#����D����E���8ԉQd'��:d{_o��X'�T��LS�|w�Vl�H�3��^��=�"��E��~����@�R�jB��]</&�U,���)f���|�;��p���G��A�������8_�=����S�
E��ҥd1[n�||+��w6���->�D*���rmwp�B_N<+!igw�_����Ki� ��*j��kcM��8s�S\�뱧]�nWI��ԫ�ޜ�Eڥ�\�ð�������'VF�u�iP�dU������tT���Ɖ���!`��P�uށ�W�]���Y�/{s�!������,s_l�R82O>�uQ����!{��Φ4�(�ip�'Tv���ￏR�hj\-�P]��p�ۙi�"�,L�g����	�-�ݷ~m���D��}8���z�^�q�8�����g�����]�v�c�t7��f���n�ɾ�]Zu�{<�Uon��i��0�5��߽8��w��4M�.��P�F}��ԋ�^qZU٧��
�	I�t8�jů�}6��N"E�k������WIXb�zC4���RG-c�\L��6�PQ3N�ń1I
�->5%�e���h�%��! �g\O���Ĥ��څg�����b�p�Ku�;з\tV�`��i�"�1�|����P��5V�U���]K�LU
jj��H��Kŗ�~w������4��gx\-><�෢[�Y@Y%Y�_|�j#�nW���L��B���>��b�-�X`�-/��է���p��x@�}�Z�>�u�E������O/%�_���E�A�i�%G-�b��N���. QdsQA�ޛB�uU�u��G���F!�De�*p��q��}�Z�Y�/��@�Q�|-n���
ψ�T�*�Z��ki����K��W��t��	ڋ�jϐ�f�M�,'�on�k۞�Lݵ�
�lq*��)�'����Wq�vR�+��Vi|�p�)���\�̉P���ϻY�t�DN���	}��V�s^����>gQ�>�1���	Q;v)"�9����������҆Y�n��n�#N ۀ����6G4(���,�Oo�_]Z�pOo���ߔ�y��$#jaH�;W��	����#��ǐ��������i|tJ��J��򦴂O��<Y���E�;������+Q��
L¢:n�\d:���(��USUX�#�b��%f�c�%G����i�vjb�VBb�l�������Y�^&����Ԕ}��v�ݵ�.W��ok��}-Uy�=��+P��Ӈ�ڮz{s��q�s�B_�ڼ�+���"�]I�ۇ���(�xp��s�5�ӹ�G���]���W����}�t�����5<kR�=U}�ԼјZ��v�g�zC��nӞo Z;ӻ��y��Q�:�Ͱ�3�nv)�gv_Q��s�,N�0�j���>_�u0�G
f�Ȟ-Ƌ�nкj���X)��i�=�k���<����{Y���^v^{������L]���B�m�Fe]�OzU������l�$��g�j�Y整x����z�u�U�O��rx�N�����ǥ����m�v��CU�ա�N�Td��Un5;½4�%)��}?\6��:S�7cy6���Iw>0���~������|�L��{7���ﶨ����[���5�f%w�v�����ނ���z��_b����<P�r���6�� �&�0Mȯ��Q����w��*g���+��yW�+U(EJ�o6;U?��Ahi%y]�JZ�xc�*Y1��eq�J!�ND��{�L�뫂,&{-��y����Ud��2�\�}} ��{x$ �TH٨�J�=ۡ�E5in��GhR�(��uc�F�Oe*А>f{7�4��r:���<�>,����x���jG$�.Z���{������x��Ã
o���ղ��7�#Zjk��������+
�W�U-���}�Ġ�.M�ov���f��n���Y�b/k�E+h����qn��Me����V�ZO�*O�g~��N�zB�>��V%�x+,X���p�����˅��١�K�����]����#��n�M+JN���R�i��=���>���z��޷��siV?q���Ң��!��_��H�n���őB�i���[��M�ӑj ���ݮ�q�[���u$���,�c��w�Ջ��{���]8��G�ߪ�a���H�!�4�/�!v� TI2(�rk����S��SB��՜;ߟ�������|)��G���#�V�Y��ﾩ��ٞ����h����-���ӄt�.�e��Uo�<�՘������H~e6T��(]+��Ÿ��ŕLnVN4v����Ӄny����&�ᶭ��yQ�r=�B�k�[�׫���ߪ�Zܒ,��ő�]{iY)"�~�@�aQ	��Z�3����"nup;�MS�ɯ�����6��i�j��d|-�����m�6�aYrQNu}����eA�E^�>�zi���y:�~���6Ydn�O۝Α���t��?eeg��O� E��k����<XGT�JTI�E6��8T��>-/�q�G%D�����F���p�^��잞~���c�x�"��oܾuw���ME9�����Rx��X7[K�$�Yw�j���iO�z%b=Ͼ�+�}���u�TE����~9w�zgܟp�HU9��fx�e���jľ0�ՙ�h�G�S*f*��ԴK�_�s�ڡ�T�h�E:�����K+��Jλ��D��T%���_8d�pӍ�[�"g�e��*.'3>�������I��1�V�ƀz�j�JX@Qo����[�}�����r��g�<�1�Z��j�c�o�F��ˏ{�c�yvll<k^�m1�J����G�ζZ��ۏ�~�Ξ�,/y�M�G��B]�
iǛT-#�?fy�J|��8�NCh���H&0����iw��.��o�.
Ĭ�����/�Z�r��}Ʌ&	I�軎�Ӕ�����x��d�U�T%�:#N��b�|k)��TP�pKT,#U����ޟu���봷G�xM�F��f�d���Y@K	��y��lU� Gd�j�M5r�"ԥfU)N�Uu}��''LŖb:I+HW_N�����p訅��Ж���Ns�9	��I/�¡I�&w�xs��!V��E�afs�z���ب]�'m)	~9��ϊ)��RKu.��� #>~1	2�$���I�������<���&���G��Z_*�r����r$��1IZR`�����/4�d�`�T|G�q��+S��i3��>Oa�Q�	i�ʲ�7�<�ŷhfj��O��=�l�o�ojH�i|�����\.q��v�Y	�㥕7}8�
{)�Bf]���k���.��	wsڭ4|-�e�]���QB��_���I(H�bSN1Y
���~A1�LnF�)�@=XYE@%�
���k��y;K���i��s뫄k��8*��t��sKbNsj���Ey�Zizؙ3�Ǐ�|�җ3�xTu���+Ϳ�y3����v]�k�f9Ɨ���M�׫>���{:c��֫�*�<��t���	�J>�R��L'�ߩ߈(�ia\�j(W�<��<����g8����{���8)��J�p��4�g�v�˛=#���l�"YK!M}}�MG�
OSM�iY8��*��wn{:)���R�;j�H�A�ý��ž�f�G��n���2�;������<9i�a���uJ�Pڣ����J�y�3|�fB'(��j.f�J�����Y�n$yI�z�'��8Mn�&(
�����y�;���f+����M�n��ln�֌ 0��f�֕�b[��G�mq���tCFh^5���l��+�f�e��O>OQь����U�ʠ�'tg��y8sx��n���E����	,vp�JKR�����VܢF2c])Y��k�6��c�+ak]2ʂ�ie��^mg=���m�kA���K4en%�B82�f�)���R�*ڲH�f�7n��ㅢ���{��x5�B�"��c��w�.%D}�X��c��e�;_}鸱ǻ�sVbϷ�5{�B�V� ,�6^�%����d.����d;M2��K���3(t�:e��Z�,TP�.R�*8��>-,3Z�z=���o�3����I���@r��M�qT��!�HRB���V�#H�P��%+����l|W��m�z�4؈Q\���S���	�X��35E��=�T,X�UN�K����p�\)8%��4)��}_f��Hbs
��ّ��M����	a�s�]w�>�����i�N"�ټ-\��f��5r�ؗ�y���ꊧ.9	N9/�#�YB0������t�� Z-��S/��W����-+(G~����ɿzdT+"|ՒF��W;��1L���t,��J߸��cn�ɵ�p�]�<�#�X)�wvI�cM�j�%)c�WH�5H�B�}~�܉hʧ	Ӟ4���k�����c�YiPq����«k��Vb/���ľZ�&�p���͛5	}�W��֤S��8RtJ��Չ�����g�q\)n8CQV$��/hzx�Ͷ����i�N&�tA�J�!4E�j������qH^�+!I
�==�Ӄ�&.]�s�*����S��=�ݛ�~;1�Y	t�Dş}s�ش�޿���ۭY�!x��z�xXYb���8Z�8.�GA���h��+7�|������T�I�ѩQ�>}�d+��k�5"�+���>����s�^T���Y���F#��RR��VoA[k���4�+i)����|I�g��>r���(E�ѪK��.S�O��_�|y��^�A�B�k=�b�~�+��#��t$kS=���NNWH�x|���/pK�o��i�8/�����u\���uϐ���ό��g_�{	�%�1�1��_���]�dtF\�������T���i���%$.�_,����;�ƾ�e��1W=�<Σ��q��9��,��/L#�pVf��a�Y8�;��U��~$�#���7��ϯ�߱ �M��g|�X������m�υ��:h��7���z%�ED!s�P�m21��\x]��\-/���o��a����xL���4�JZ�ޮ}Y\U���#�o�]�T��g��^(�"�ܿ���j\�U �e��-;�6��ĉ�K�}����z+\	�*�����}>}]R����>�Dh��}�Kĕ_��ƕc�m���4Hz�m��[��e��vaed�ۏ@��1w���������hgY�K��]j�-���&�cu�ۨU8�E�t�axM�e���Y٨sGhH�T���7%��ї?o�k��|�E҅bVX�����x�8T*/�),����oLK�\�d��l�ͦ�F���n7�_ů[���"�/�62g���2�&h��Iә��K������UְK�>�]�k�pW_gj�'�/WFP�f�TFww���W*8/!z�TX	nU�Z_�N�Y�%/k�+r%a}�jj���b_w+8�U�3��-�a$/zu�>�}��T�%M6K�9�q��Wƴ�K#D��}ߺ��t_u����W)�ƚ*��vo|\/�ݯ��9y��K�<cW�U���+Ͽɱ<J�V�,v��2�(�DA��&Un�Q���/�T^���V�5\JLyG��� C~w|O���:�s�>M���n8I�J�äabVƨ���n��Ri�s-ƢJ!w��*�ꀨsCtT��-!H�A&�93����W�Vgp��4�5��n�[�Ĳ��n�̿���:�=#Ｒ�B��5�K���������&(�E&⟴�����HW��ub�~׿>��X����/�k��R�EU9t��J��r�Qd+>"��|��_M����ċ�jȲ=-P����~����}��z�|*8G��2��5�,=�������Դ��U��!P����g����*��Y��U�����>�'�R���޶�Y6X���t5	a[U�����e�����fĻf��K,��Z&��о���f��i����Fp�9�U=��X�,ְ�ii����.f;L+��8�g{Jţ!��g��T-v���"���VT���B�t�-����E���N/�HE8L��T& �^���6er��������׻�߾��E��*���Â��=?�=�>�O`(K���R�W��.5�J�Gb��d'}��k�93�8)$�$_q���Z�&xV����Z~&��5�YN,�G�w��vw{4��{��=b���s��0TtT.�#L0��9�p�]4TCo��/�M�Ϧ�JV���
�odS�O�����'-�f��W$}[J��+o�X���O��ԭ^Z���,���~�]���_ϝi�0&���H�k��,;�ܝ^]1���v,�t�>�կ��Z�
L!}n$��5�>իK�����6��n���>���.�O�ؖ֗��K����%=���YJG�|���'ע��}P����L�g����N1���7L�n�/�<��!����W��'8�_{ռ9׵��B�ǯ��N8|.�����fcKO�/��UiEBfp�|�g߷<�����8)Dg�쵢��xPȰ�_rUSD+B��gĹ�WD�w���u���;�W߈�ϢdIh�jH��=��(�>�����ZRG�#����V�'�[����/���V�����eES$j	�^�n�W�Y�"3qak���vѣ���Kv�-ȥ�C&�k�¾�/{����"��fN��{�'�����7Ͻ�b����F��.������*w�t4���fyk�;H�~�v/�mC��-¾}�ZZi��Ջ�5b�<֊����I�Ea�hE�w,�^ug��œ;)H�_�ߋ�����L���Wc�Y"A�9i˂�6��-$�!P�"��e}���j�K��	������+RFk�$��|���Rre����B���53,��9m�a�`P�I���t��}�qC�m�,^E�>�V`�,9�������_����a﹪�˜����X	P�~ٲ��Ū�Ɛ�o��+#�k��>��.�eT�ە35S�@GF3¢��˻�������}:E�L��kH�5��}n�Ze�jD�>�B���VC	QB��gŮ4�&�4���=�-�����8���z�L�rR�۩VB穬���J�u5$�V%����<-�k�T�)�����~v�#J9̘S����	A�߿~7#��yF�����
Ԥ�2'�@�$R1>���VF��_M)(I��g�xp�pXCX�2�P@�'��P�8����U�z��5h��%h���Q���`,��^X0��{�����]1��s��Ϗ��v�"^*�6�¢�Y�m���� v
$m�3B����Ǌ�u��]���n/:��\bK�(��Ȑ�K;��m����b6+��+gEh���:]�`熦v�(.�^ʹg;��4�kQѮh���.�����9.%�K2����[d�K�f����t{WnD4s]�.TK�ng��V�e�.���c��V���4��IӰN.7%��3�&�:�=�"�:���ҘM��l�L��+�;�W��9{P�SO`�7T�.��A\N�۬rk�Ӫ�GD��%�ϭ��b�h�U��՘%�Qc,�DX��"���\h�����rV��4���'��H�_y���p�x��q��`�/sܩ�ZG ����>��a�#5b�[�'w��7��mΔa�rm+4�'N?O5�s܊#�i	�s���Ki���GP���%n����zYg��y߈����&h	=�\Y|����#J������Ng��<��쳫��_o<�2�*�2*w�.	�ݕ��b�Eӆ�}���ギ>�qƐ��n��3�x��~/ȏ�	ۍk-�`;��D`��i8�g�+K�\�
�WR�,�����f�9�)����ia�pF<�8�gX��SL���\��0�Z��������մ��)�����`�R��B*j�EB�z���j"�K��VB�~�K3���.�x�J��>)�uu�a,ϱXw\u���-N�ΉicVG������*]2e��L�ё"�_����$%����|,,J��
���1ڟ}6���8T/Z��婎������ҏ�en|����X�xB���+���>:�q"�q��V�����\rN��4�Ŵ
0��h&��Á�!�K,�[vG(�T�bRݷ��������+8A-�e�h����k��:"�ˊw ��f{��଺`�TBb�\?���K� V*CB�+nю��}�i5Ю�{6d���C��4_ry�k�\� b�¢3STB7�g�#��"&�wy�������z�Iy��/D���R}�깣2S��Y5���'��]+S�����f�Y�^���|5`k��<�^|�k��m��s�uĂ�Ej�1�;�~z�X��}�x�D{'�
������"u��oU�"~�<!Y�}�%�M%��yٴ/�y~�s}�g�f?/���yQ�YmX���sz��uH�&f����I�=sn�;�"��+~�/�Z/9s���~��a0u3�{x�pZ}=Un�K��\��ܧT��9i3 I�^�s�[g*(JD�U,���S�q����J�b�dh���<�p*S�2S&JS.��x�'��W�,Vgˋ�5�>�����>���?�_�t�a�V�\)&k�vn��f�Un'�2����ԯ�9O�bq�bUԷ�d�~���!}��p�0_#��{z�!�eQ0u�d�T��b�3�O/;�{��Y;����Q_l��/|8�Y���b9���y���w���8���Ր�m�ߵ���͞H����&ۋ�^ij���L�a���[��O>�\�?���K��asr9/`�[Zڸ�)��j\��.�](LK����b��*����s���5=VF���a
��7"Y�Ϸx�I��Y-�B��s��_���&;nFH�[m.R��ϋKﺻů&�Ti
��ak��o�Z& ��*0\����|���Jn�R���EM,J� ��8.+�i�H"�ٟb��[Ƴ꿳k�ߧ��}�e`�^~�w��\jH��g�&�Fg�}V��E����i\��0Kw>ⴤ�p�3�}���nw��[����ݑ������v��jU;��8G���N��U���VZ�4ZEJs�L+̔߽6�]8B�|hW������&��F��.�n�_��,�=���!��O�r	�G�#w���Ny~����6=��0٩J�d���Eq�b�>�s|b�8F�Ec���,K��[�8GT%�e5$��=ke������CjYTTb^8&h����[�}~ŇgWR�#��zn��"M�`���d}�ߝ�z���&�KK�ӿ{t�
��Si]m)v��zs�Q�^����	uN�X��i��N���Quek�\��'���g-z��4Toޔ���2���h8��'�ȯ���dN������履�U����+"��E�%%�J����������i�D��0����x{a�[�NF�k;��4������FX6e^��g�V����ɰ��ۻ97p1.���c�n��@���J����ϝ��MKl�Ϸ#��>j͖ھT��Z�2�z~�Č�q��jA�*�gu�&��׾�pﷻ���������~���I�eh�Fg;�xzj�=��١`�]�e5��/�_s�r.�*�'!(�S�4r�'����dX�����ic���/�?}u�Qܼ�U4��|E������k͙�DxRG���W��;K���妕��K����f�}��G���k�ɬ��s�Z|%�l��O��!�	UB�4�uF��I�M�I*�!+��K��uk�h��f�3
��lGo��ڔ/��b�y���3}����\��n�]���p�M�S�miW��8b�8^���s1w,�o�ڧJ�M)u3�"�r�?^7������Fu���h��Y���;�KE�S8,��p��7��^Ͼy	���qN��>޾O��l��<!{]�f�s��|e�ǿ��<��;Y�C�Hw����K�|����9��������������wbw��?M��[�"5f���,i���t?F�h��]Ǐ�~���������8�,�
��jȡ>��V�h%�3RD�S����ƙ�P���)�$�o���9MH�YW+����W��5�^���¿��*�`�}�J�.WW�fғ[O�ً0K �/}���yنtIז��ZSzD��Do7Vs��M�
��r����4�	�0��A�m��#O]E6��y����:B�ڵ�sZ1hՆm>��i�iG�B�Ҳ������Ɍ��ͨ�Ya�����ɴ�pbRD❥B�;Ɩz�Ϟ%sKT����8b�Y敔GŐ���;�ӳ"b�����j@TBﭟ`P��t�I�c�.^ϸ�i/qАt\=��5ʿ��,��.��cs���@S^��4��{�.0Z%E��Y��όKٮy�X�n�u�e��wU���D U̷���Ux��SJ��dX�������f�z���d)o]�����~�ݲ�f��3n�ҭ�kmt�]��7���g�}�c4\��g��?g���	s%��&��g��KM!�B�������L8B�Nx��fH谅X|��"�jjLFN���{�}�u/&��}���O��ZGG7W~�3��2�&1pZ���Z#�
����^�%��[nj�	z���s�:C��m%����;����f�'W�N�
L#��8TBdxE[�S����K��tL�;_
�#�j�³D�T/���o�\.
ȑ2$���f��Ⱦ��d��O��Dﳓp��~#�!Y��Ҡ��)�3��E���JV-���>�n���Zw�J��'O�r��U8]Q�Ŭ�w��I
��:b���ƣ�ډwS�6U��i�kM����9���m�+k�c	�����}N��sf<��-�ʕ���-�,��=�@��~���	2x�ǫ���.�Q����S���xX�#]�7�{���g�� �5,� 1w������L�|{ur��`���jB�s���Ń���Ǖ9Bֲ��QoQ����x�Q�{��.6�k[�,�/ �^�4�owc��9�܇: e��E�%랚�:B>��{P�Ի��h��m"���e��p��i��C��϶��~���X2�o�:jc)W�5�j@�h������װ�Z2�z�U)zr����׏�i�gcұ�	�+�Lz˨�ǲ�*
g��	2�:R7+��D�u7��J��g��w]J˷�{+��7;��ꓻ����3�]��1w��Z��7|�η�W�x��=�o����_��'o����v�vv���,��Vz�M�4J÷nD ��;n>���Zu���M�9���*��pj�퉄��{Ї��� O^�3��[s}�ˇürN�^��e��k\"�vi֣�˖j�IdJUh�{O��o혶����S�b�/��U媊T&�2�����b�^ڣX!�]�ؖ�u��5��\��yJ8U��=d�?Jɽ��M;�Z5�g��!�=����|�H��~���8]��l�f�p���3׹5�0قyaba��J/3���K�I�z�=�qx��ρM�L�~��X����0j�; X7���#sj����}�$C���gX��gCM��U]k�<-��-jb�RX�� �d�6�NPf%J8�A�/)6j]L��Jl��9������$��-��9��:퇳�xur��vĨp;m@g��F��rC�,�� �a�i�Tˤxh�0hmU��]�6`���eX|XݹǱ��̈́���9�aylZ�ۓ�$x�*W��8�OK��	��q��ƞ-��v����"ae�|��K��T%�7S؂��7�Ѱ������Yr�Ԝ�æ�6��lCsVBY���_��t�延���+��S�6MQlr�8�,f�'��9�'n��<�;\���<��]��ی�4�
��R6˵8���%Ӟn��GV�4�����z����\z5�<Sq!���D�]s�d(��烲�tvU��9�i)�z���	�|s=3����ͭ�urD1f,��m4�(V�A��2�e�c��ʮrf�t6��G+���'��#�T�vsp@
p���wS�lmP�
�:pY����Yǳ�h���)�n�r�p�d)݈�RJ��g�b�,�jQ�j�m&%����lq�/D��շ�@��^��qB�b�n!�,�x����P�,����j1o
�Ln���37O����͹�[�3��5ܲ�l4�i�mV!��t���u!Em��,��5ɇ����;��rv��I�����t]�{t��}���!v͇���hvR����^��/���\rtW;[�'W
7;x��x���-�"�f���{�py��+J�G%f��y���[���K� h��.��2%�I`���R���Ʌ7A(�MHK&�19��J������!H�ƗQ��\ih��r�tFgm3��뭖,�D��/;l컒A ���'��A�G �jy�x��vǱ�nk�j�F:x���vsl>����h���J;֔���X�##�Od�Z+cU�Ysj�BĚ��m9���`�f;��ans��ގ����<xxBܮ���ZP���,�t.�vL����.����E��>c�;��طFd�@vw�׮"놓�۶��M�d�˭J�x�j�ӻq��p�M*ɕ6^�/�3jE7�]��mǴb�xL��B�$��42��u�6�V�X�yv��Vs[����/m��\�1X�fP�D��ݲ���]��C��Ql�p�&�f�r�����xle{�-������>��4��-`C
r킗:�"pv�c����̔��N	3n�4��
�m����}�DXE�͔��,�׽6��.��Yш�"T.|��٪�H�8Wo�4kq³�Ǿ��^�V��~Tq��=��\'����
��������ݰ���Y�����}cdm?���2��)I�^�E��T.��Ƥ���y>�Z@'�>oT��;���\��H���߷�c�h�۩���f����g�+�[칩��9�p�%�C���=��R���S��17XA�yu7ҝK�.��7���4Yy��9��B���2#��q��ɍ�M�B)���/	M�!r6��e�¹Jj�py�^{"�k�GM�>����p���}�����Rn{�Hg��{���o�M��|:��@�p����e�5Wd�{�%��G��P���+�[|*#>�b���&G���U��t"� ��4I���)�����ѧ���{y6��lu����0͸�h����Sw/��ڱ���5xZ�2�[ll��N�Wܺ�X̩�؍n��[�Cz�KE���u�����N����ҷ��~�ޡ\�|l�,Gęn&�(D[�{+���W*�k�;J˨�L5XQ:Rޱ�o��=��<�꧸�I���|=���������x2{�����{r��پ�T����^"�`�N#��}ސ��~u�:��ď�Z{��[W�6_j=zv��A��
R<�.	�p�Mk�:��zv8�������i0��=>!�~�����}�|��d,���"`.��\���^�r�W��7%V:��>��.a�0yj��i�n,�T�W���~����*�M�T�5�$�1I*����Dw^���Viͪ9�2wu���;�O�CO�����"���+��s�U}�f�,���3����}S����G��,����C+ fe,�[,�@5
�]vI��ehƋ32RN�^������z�_UʪG�fQ�a�5����X��cB�{؅�Ѻ? ���4�;�H��糎����p_A�]q�q�9[G��j���>ݫ��^BG�vy����(����R}ޝd����z�������	8�Ń��f{.�4��h�w^Z'��'��Ofk�G2Y%��L~�XY���~kؘ��[[�V�E5�~]�ǫ~��2�Ņ�3Ajq�ٶ'��<H ]d�X��\��z�^y��a��;<ru�Ah��&N�㒓y����7�u4�n_���Ϣ�v��\B�h�~�o����p�}���޿{�[�����&�������������Qk֞Uq��N�jᲥ�˫�7]�GU��r~�S��0n�e�0��4�w�~�|�b��\Φ����.��r���� ����l �݅l��Ƭ��\j�hM\Jܦfenc3�(��|�~��]y]u�Z�ܹ���c�v]�+����nc~�I]v��%9ܫJu��F�q����؍�Ҥf�]ٺ/5�b>�f��C�L�ΰu���ݲsզ2K?~�1�M��w�������7�Q�~��O¸mp��[2E	pE{��5������4��y���M�RFiV�����,�0F>�4���x���Ǉ���B����0��%�q#��p�'�z{���|JX��s����s��byJG��&���E���c~���o��r��P�c���^tO���L��i{�#lK��95�cM��4{�F���;�}��.!�j���>}��l�8�i7],LW������$��ʼDy��0�:�e.;yWn��7�Vhu���>,�EM��R�Iμjk{yW�=���J�$�3&��ŭ�--��$4�`�a����H�����ػd�����p�9� ��ޟ������5"�ŊR�;�{�g��dv�\l��z�kad��G�r�M�3;�m���rOb���\/��P��}o�؍�u^��ޖe#��F���{z_Uܹi�u��}��|���P$$��Aq4�N����/zY�_yW�kʔ���b�n	�f9�ϑx���~�nԫL����^u޾�x~K{w3����� ��$S�m�T�%^>������7���A�4�m�?R>&_Y)=��c���5~�z�%CV�0U��W���`���6��4h$�8p��	A�`���]�|=�}Mo	��:γ�'�4ʒ���<X�A��_G� 8����ݐ
!.���}=��{��?+ޥ�뭕h���|�a��u��;͸,k/1�#�w޽����׾[s�����E��%�K]vM�2*g��Q͐툆�hE�Qa3��[�Z7L9�#p�U��y7Q���n�3��#S51
��Տ%�^H��x���l49w&Kj�\G�4�#b��&	�van��,m�CvHփ	g���.�қ��5�8�/;D;�vP�Qy���wm��b�g�n���.��>�hNۛ��kヷ\��;\:�����)YB�e��L:`Ʒ������{Ft�Q뭳�D0<;nP�=x���-m6��5�S	s����@�`����%�$O��|�f{&��^�R��c�2�c�~=<yg" W����:�G����Te��fT���w�5�&E�8�g�v�{]���5����E���+�:{%�x��i4;G�w۵���������;��/".d�I�,�h?✺���zz$�WAx�ʡ5F:�s��Vxe��'|O3W�	ﾎ������s(�5L��2E�GQ��L�q����"µ��s���%xז����l�|��D��{}��j����us6�<��%��u5����S��\1�#���ʩ݉�g]�=E�ɕ7���?,����{��z]'����I'�����ٯ��o���(�=9=�M�X7C�Z\�4�*ݦ��z���E��.�A�w�&ahK5�KRŘ6C��u��Ĭ_O��-�������k?Z��_l�s���]�w���"�DԖ���7��aR930�ۄd`���s�E���_��sd�9:ϔNkG���A*s ����'|m<9�h$7�f/���B��Q���0�\�����~X�t45�w�7�w<��>x�9Ѻ5E�֮�6k*��BmgaF��3��X�~4�D�J�&G�A����U����l��j����O�D=��μ���g����H�@���.s˗w���X���#0hF#@�m��`��c��ҩs�!����^6"X��)�9��1����ݬ�x���B8����@ِ6�q$�$��뷣�o<L����̽t����[3fR������������p��k�.ofC�߂��۲|+���eV��Ϻ�����vָlj:Ə��g�L1ԕ�%��]*ֶͮ��M%�XA��6��!H��W�x1A^�~���9���ܜ�{}��P�^&��&EW���������`�������q��2�u�u@CUT�����N���K��;�.�ڜ���?<�twf���?paZ��{WMDj^�)H̉����Ԏ�%�F<v����r�Cԓ���G<v,����;���
�B���>�͔�ܵ��=�<�|<cD$ލɣ6��!�̆!��UƲ�Ɓ�d�u�[���\n�+T���17���}��iC,��^�ba%�(*u��]A������5�[��E��OjZ�����R��Z�H�X�h��oc߃�_��?�S
\���jB�L�K%8��n��S���t���Z���Vd���L��La�y�w�N���LL#�OL���*�KM6�8�	(�-/��Ql�ư�]�1m�Lʒ1��(W��Wb�*E��ʒ(��T��,u��*�j�zo�۵ׯ��k�F���-�lԷ��y�����{�Y)�.��i�JbS�������ݩa^�f����A<�yҾ�ˑ_xev�e�eFm�QӋ�շ�;���$���SJA�������{]�؉c$�`�R�4g�gIr{�y��ᱣ˹el��Y ������;�Q�Z�Q�]��і!��F��,d{����c�|��N�b*�ԯ�ơ��|�rSr)D��cF�i��?��9 �j��۲C�=ٸ�-(�}鑂�P��R����N-`�c��tΕ^\�����V�	6���)��so�$��,X[ǘ��o����Oj�P����E��}�k�խ�w�mAf�Cҍ���T���<��M��gX�뫋�1<�؝���q��*Q���iF��5e[�u�P[��)��Z6DU���,��[�Ϥo�9�9 �H�~_��P�$㯘^��)��������N{�lϨ��*I�lD�����,���齖d��O�n��Q}��=�T�����zr=�E�r�;a��r�=3½�Ǉ�VS���8���A�b����2�/�r�w���/��7s�٧�E�'��zNB�E�*o�͚t��<��wS�M�܆�#��5�Ϊ�8v�b�zυ�}�����h,|)�}���{�Ԯ�RWŃ���h��S��!�u�Z���n2�q�SI�s�{R�{����i���;ɽ�~��ʊ��z���=���Y�o����u�c�5������fuR�v�Rz���(a3�^��y/d�gQ�_>��]�<Z<ϱ����"qӍ���lܙK�%=]�h�*��f�h{���ڙ��"ͶG��#ue�-1����j֑cչs��Sε����T����@�P��7!�4A�x�n#�֬6��riAmZ�m�(vi�٩s��^Qâ�ۚ4�4���G@�&�j�9�Aú}���!�u��]�Ƴ��s
p/�uV^{u��^���n�P&� �x�8퍵�5��l�]y��Uӹ2<�.а���pɳ(8%�[�R��@#&�˩b6�x���#дk�n3�x9f�D)l4k�^1+��M�[�|}��F��E[���}���:Ts�u��(z���d]i���bXS��=�3��Qe"�IDIݔ���?E��S{b	�����R�`�=�^�s�Ǆ������t}�6'I<=��G��=��W�ԃ�F�jI#r;�G&X%ys}�>Ï6�5�j�3�o;�DK�×8o̿N�H{kܰZ��(!D/o=uyIqoy�1���i�#�9���}v��$��:��I�_]�x腈����X~R�}{�U����~��r8�_���m2Q
���S��zٻ6U��r��)�翾kM8]�R��O�S*���Y8}��
Fw���e�S|����]Z�wC��T�F�x.�/8���gK\��<n�(p�[��ӹ�Ԑ�(��0irW��'�'N������_�z���ړk�-��ק�%�8���L.N�;�|w���r]�Q�$�'!i�k��O�f��o��}�j����zlpS��I�V�V���a7�71�6.;G	~��g{��z��Y�!�y�.^�I�B&έ�3��~y\�Kb��б|?tO`�-��0�6H�{����-`ӹN���L@c��RGc=n�����������#*���L{�oNs%(}dZVŵ����nM̞��u��4�����0�X�EM��}���9�~16�����c�z�:�z�rW�n��f�2%�N�!Ӫ��Q�z��#�>�PPcvG���n�z��e���z޶s�D�@�2�I�w:|�(�v�g�ܵ���h��j �����^��_ru�~�^w/��%��Ʈ#&Qۭp;t݃��n0/� &����J;/vq��N99h�n�jT�^��+o�t��ߔ
����B�i����g�n�w�}��fi�Z�M���2x̭�\��(�a6a-�aH2���g*���[Q��>��]��5��F�(�u�vN�������yYN���m�t���u��W�g�*$a�e�ɴ��ݮ�qU�k�K�O�5ޤ����L����)j-T�}���W���,��;���)��U�J��kj�����U�f�I�*ڷ�[>Ǐ^]���=��i���C�<���rm�˻��P!�c^^��n��^�pA��x�-����V���ǭ�Ѳ����r�Kúʧ����aW�02rTf�����f��K��w�ڵ[���9�����M�{O01��Ȑ|�Ů^Ӊ+{��H�Cnz�/Ϝ��3��X>�4t�9����7T%����I�o۸kp���{h�����vb>Wۮ���4��$��kݯX���_�l�J+9w�-E���x���@+��=�
�,�uIp�s~5��A�A4d*��<���rh�v��=w���!��=�d�+2_u?�������}�����+����P<J]啇�T؏���ikj��iAJ$e�3IIY�K�����͓c�+�`٨�^W���Le:�ўx/f�٫<�h��ɐ�b�8.Y�h�j��	��6t^�J����{��Q�m�۵Kixe���3T����G�ti�߫O��	�j�wޛ���%�~b?���սo}�W���[��L���b����i	4˦5y��y�I���M�
���NQ��{޶o�ss�[,wk��j��{du:%o J�Z���.��7}�1�]�}�͎W����X�E<����p���Ѝ����l��$��o5K7}퐻����}��⯆��cGa��f݇�Ҟ�}����^��:3-{ː;���\��}��x��Q�N�k�?��O}���᣽n����R68aB�;�ٔ(ZL��!�xg�{�2�H�}�����m��uns�l�����8���/�����&��2����٠pb"��D܇�M�	x���z둽9TX�NMR[�֝�fh�\}WSu�ڮK���U-��H���|���g`����ZJ�W�:-,�1�WWX��̍LC`sA���0kXĕ�飃l��J�w���\�\�?t�R}������~�,��B��6��[H�<�j����|��1!b'"wla��;���=ޙy���ݩK��%"sUQK���|dp�1o]uZ��|��x��t����q9�I$%p���d{�z��u���Y|>��}ׅ��[st꾅��o�}��`x�ߚZ��s�x�^"�I����AM�LQ����C߾Ť��G�}19=�&Ñ�������P�]���@������'VV�W��x�K�i�b'N����m�oV���"5$��s�0$1v����/����'p�muL���Of�d�<�{$�{EYex��G��ΰ��H�M8	RB����N��^n�������A+�V/��f!�%*��7��s����G�G��u���}7[���`5�n+�gn����)�V��d��Љ��m*]uæ4��U��2����"C��㉝0w����X^��E]�Fy�P'��+�����^q��z,:Z��Û�S��av#?H��8���6�[�}|{�y֎��o���պ���/�.?T��|פ���Ԗ���4<�M��X�������{�9 e�E�r�l��}~s�VfS��]ls��K�����؍��c3�L�AJ^��~�[<����C-2��GqIb7z��F�I��Y�ܽ��nJӷ]�=�q�-�ݔQ��)�Ku�T��(p��u:����a]J`���x�8�NFڑ������W!����w���"bd4UJ�x�G�h�B�UM������)ל�E�Q3qגeM��d��Ru��X,�߆V���T<8_�<~G��v����M���f�i��������_S.���w��c����./�?�T�hX�a�L�ך:��v���u"^iB��,[�Ǝ,��ۭDh&s�-Q��	I�[M�3�a��V�P-)kUn"@��<��<��H�8����N�y��lv��c�q7n<�9�8��0��؜�t&q����-0�}��X�l'[S��8+����氥R�-���f���b�.�;X72��c�hv��{�<a5g�g�ބ�<����Ƣt��uAїŀ{{K�N]!�@�5����q�{Hs-�ܽ�i�I&�d��6[�"��^����/�<7#���ꯄ�2#&�w}Y��t�_��\�U�����Ok`� $ �AC�+�MVK�vW�s���,�'m�o�}^�ϗV>|[D��syq���=Y����L�U�i]�����0�a8�7N<��[��o�D��>?>
ˋ���di=�q���[]�5k���uk;�-�b8����V֭ʝ{H'��zcL?O_�=�K^���d��.��W^���غ���7T���q�%�Z���lo9�[KD/��PhEH[�{1S�ȏN�.Ǆ�t���/`�}:뺽ö��f{�!~FSٻ�*�Gױ����R����'��v��i�����K��v�h]���ۭ�!l��;cg����u�l)n�k�m�A:[��<���S�����e墫6o��
���ݣ>1���6�)c��AaR�ĿoF�I1m4ˉBB��D�?*�z��3G�>����p}z�*�3�����>���1�zsWk�b����Y�B���_m��پ�w����O޿_��E�_(�:sf��Ͻ�R�~���z��|é^ucn��=r����>@�ı0I��v20�0K�� ����s���aF��U�u��O��}�ҍ���z����Ͽn����� 2�O}��ϭ����]{E���o�ǉnj�p5}��x}O޸O�U�TՉ���b��Ա'7a}���8̓�=J�d)#)�$�]�`�x8����=x���p�)Ƕ./��|�������P�k�8�mq˒X�9�.N��x#�N�-�q��se��+]08ܾB���g�l��u��<WG8��R.�i��_.>=Toj�:��H���m�J��8�y�P�;���wkR�I�_|�ϛ�a/C1��"�%8k����w��W�7U�������پ<�%��t =q���'�hf����!x�2gY�8���#R-�bz�mi_X��v48p�x򍣓h��B���(�=�%Uǟޘ+Z7�j��y �U��ك��������o���h��Ys���xu���qKy,�T%�G��"���U�p�M�����^4�,_�=�ӊF�P4�r��Aխ����}z�2g��ޯ��3����}�j����h�ή�i�/,0������4\�D��sjn��W�d��9�5${��$u{�i'6ҫj�M��W:S�n]��Ŕ�ӏ{�:�g��!ں��.>����GZ�R�R��t���J�&���͙H,�g��9�B�}�n��{R�T��d��8�RA�vcB[�n{��t�Z!C���L����鶏��I3v���m־ξĻ1���N��	JC�P�n�Of{=�㩎�A�VU�R	{�ț7�J��^piث�ˋ�F}��Į�����Q�����3��-��H�M����(�&wL��mCY]Ҟ�*�:�������`�`~ϟO�#"Z�y�KR_T�ԭ۾�Cn!L���4��`˿�鸆��4��F4�Ww8p�h���f&���~���gN⦊j��*�$�����ù�jAU�����+��k��dR�׆�gL�kw�^�|iF�N���c����\@�('�~�$�Կ|��j�Y�Ϡ�6T�Pƍ���+)̝^y�^C���������dUGN�g�8�b=~.��K�,έ����qC"Φ�ت��-M��$�p��z�n0�v��l]Q�F�����K�lѸ]��>����B��L��w:��wN��y4������}׶�X���Tl������eI#-4[e�6�\�B�݆�K��V����FI$�}g������������}~�T��ϖ|'Ȭxw��`�Ż��bUz��e$q�I�ܓ1�N"'.�]��\��wϏ=��w�ϭ��uzRL�]a� V����R7Ty_7���pĔ�d��z=V.�AV�}��,��Y���<�"g}RoI��k(_{�;�ެ���~�8�����gue��)���Hʉ�eI��st��_ê��K��<��ĵ��7�_�w�o_�e7��_9�љ�Ɠ���9qLNVU�C���i��fĪ�x�{�5�}V#T��O7�Ǟ���H�������Q�r�zѻ*g�g�����6���x�R*]�p��:t�=�F9��-�v#P�f��Y�� "afM�L�X�����a-k-h�w`mK�%bnU��c�$e���:O��ܨ��Z��Jq��6�r�V^8����*�L00FQ��L�	��K]���1�X������,w]{(󋝠���!����w t��z�0�"���[l����&�!1��5���;1M��`A�sa�ɦs�H⮚LF$*��I)��F

9	����O��ʻ���j���6����]}7��j�ۆ��$<��F�p�f׎Vx�u�r�S�q���8�0?���
��*uWD��_������pX�!z}� ����߷�yr>��4�r�(�`���}���F^�ta��[���NG��X�s��pN�v�����z��.i�j�W��l+|�=��e�د:!�kx�@�D
n,�������Du�V<���Hٯ��1i�O�>���]���}J���Cc�+��Wv	�����1j#ꒂ��/����d�!���ڧ�}-����(=�U�N�^�[�l� ��\|׫�P��
}c��c�}L��O_���gS��M4�:[uY��Ψ$�˹vy��mQs�-�m��JX�2�464dO����ٽ$�}J�gz�b^3�>[h<V(8T$�wz�<�OJ�x(�ʡY�r�e���M�]��b(PL�qe��t��Y�,�W�x��tcv)��U5~⊭�=Fw��������l�ϼ�۱6���܏ڶ?)Ȑ^�9�Owd�Ş�!�0�t�+����i�9˴�qaxߘ��S����s��Jύ��������.�@�$i�A��o�/�?"�(7鐐>��-ai�k������u��nq����&�K���.BQ�6��;�y{N}���g��K�%�|��|֛�ͷ��vqWlcd�Q[h��{k��8��[�'ͥ�FYHH�v����]R��oNCL��DyL�����z�\5b��>8�k�N� C�G����9<�O�����@8��d�n|b�8ӑz��8
����>���I���Į%T�4�b�Č9)#a��q@�M߼��&}F��dgu�������z ��*�_�aۧ���~ıT�%��|��2[���dDJs7�an���}�*6��}Ι�lmԪ�5|z���bu�T����J�S�]�0VV���i���d�%IB	�	Hk�{���R�g�睘}�\�S�N�5�{<�W�n�l��ڗ;Q���	t+��r7�/`|Gt���Go��xs�������n���]�Vh���w������y�����{���5����{[��R2��?}�@�]3�����}����c���5��KZ1����E�'g���#�
�����c��χw�%�G�Ϊ���a��F�N
�h݉�y��@���~��@0d\E�4�H�7�� ^^��S 0��0g�׎�K؟~B�;z��t�`Ƃ��0��*�aa��\�p޹�v�\�j�76�VY�=�YQ�݃�x>]rLs�9��so���۳�en�����3q{��P+���Y���[��|�R�&�x)���n�x� 		�/�G�[_Rv�S}�����S"�wDS�x���B��{�j�Scdwu�Ua��:���s�]����h���"�rG�w���\~�v�I��P=�Q~S��rЁ���g�nɔ�=��ؗ��qvl�W��^A���	�*$�JԀ��H{��yrd��ٗ�҅>œ5�'U�@j�[�S��A7F�G����w�����=p��G��꾜��}���=��uC��*��ƻ�#���W��[�޺}|z����v���!����P@��n�p��_nc9g�i1�u���A�#"H")H�m�$��_��1�뛞�d������z�\����㓽�nE9w��i�nݜW�� <w�y+���!a��t,tIa1t�c5s��ݢ���s�N��wm����S͸�f����E�忼|���\}�ڋdzߌG�~�^�_7�T��+�<��K�����#c��7�bk��K1�1���G~<���X�n�~���q�7�5z���'о�-�Jד�d�{N{EEx˝�ݎ/�PֶI�Ͻ�0{5&2�M\�'����}�?u�D�C��Omg_���<'7utw��ך7�	1@I��w����ӿ}�[�[RI�+�JF���a���9��������sg}y6�M���	G�gs�}fI�I������^�����=�F�}~i!a�̍��8.�\q]-�*�t����q�\2f5�읏��6�n���vcޖj����)�?~1|oi���H�?�~`���kKv�񁊳�^��<���.�հY�s���V{ӈѭy���rӧ-y�G^^�.������%�^�^�J�*a����M�;B2��

����u����?����<;u��%NgD'6>�)9��e`�o0���DU>wq������A����=�a��^!�|#��x�7=�z�O���h4`�ö���5��?Cs�������O{�Х%~�./c����%8'kFV��.�Nk����?	��s�+�4n��=6�ޛ��_}w�z����01���Q�����T%Ii��Ax�=5����@�S�ׄ5���c�&��$Wzx%a�y<��j�?e��F��.O{|�������nb���C��{s�HI�١�4��w5�3m��-����0��=\�L��%gC�Z�^R� MK��Lե+Φ��~�<�2��M�7�n�F�
��w=�St<����Z#����;���:_g��W�B:|�!z�����7��n���Z�ܴ���=������<d��g2��}��r��2�#�_�x�rKz������>����HtO#��}C���n<ǍUz�~R/zc���з��	礦g�8�eM���b�g%ۇ�^�lO{o����k��t�$i٠J�8�S����{�@L=wlz��5Z��&�=�ڼ���|o���������^ͮ��͊$�{�7~���b5!k�nc�^�'x������~�nT�W�������]��l��	S]�0h�y�k�lذmL����4��h�%�IkH�u��������a6l�
.�l5-%��N7EšD=����Yi�爜ݴ�\��������\j�{l�^�˧vX�ٝb�t)��9�]�2I�[c�c4������Ne 9�Y���Վ�����3��P2#���1�L��,P]�iAܱ�.]��H�W��`�k��m��6��$#���]��P����F',ŕS�����p�;�p���0�n�)7�����u4V��٭ �ᨓF��,,,��i�Wo8:4x�O	d.�>�ר�s�}����c���u�V�m�0���#�]��m���i펓� }��`-�s�;�N�Ի \<�h�iI3.I�u�lܬx61�X�m̢(t\gL�V緌����Yc+�b��u�8w7[���ZY[��v\v��㶝�`D1X����2�%X��6Cv���g�=l����h�\��y������3�p�FV�^�8m�1.X
�K� �Kv;�s�Cj��l�ah�m��.��LG����z�j�Z���\]X�Ŗm�`;��-�ԤM��l��%�{�N��d�]1��VWX╠�GH�bn�V�k�S8����i�P��x��x�5�q���*[��y��N�8���-�:�a��u���1�kIa`��")9�6��Jl,4�1X��WGuyf�bi�]Iz�{Clg����-T�d5¶�Y��⤳r8���k���E挖XaB0Y�9/��R�R���6�A6��6'm����\�QQ��Iec�B�6�dлp��3�:�e�/c5U/8!s���lqA��lY_u�
�����BL��Nvչn4L�:��s�`�n������m���i�'k=z�ۈ��ӹǍ'=.(�5ݰ&u���K6sc���m^Vڴ&������l3�|�c�+mlY��r��ę��s�r�c[�i�E�����۰�rZՀ�,�c-��m[m��$yt�q���u1	EZ�S�ݦr�,"�';���/G��=��N�94L�)۝��e6xޞ$�C�p����=.��0n���Xһ��f�����GLļ2�ڸ\�F�dв�)2 ����֦I�� t��ݻ���l��q�,mNX[0j�p�)�,V61���ι�)����Z�1�ں�Ηa���9���[L�z�=g��eЛcP�0�U��R�f��q�T
1�`\2�]�d��zb��_l~��Xs�[r�������1���v����FA��꼕�,J�n�]F$�P08��Q����=��L3~�	�{E������o�i���>�O��*So���������P�uZ�Ѣ���#`� ��o\�~�+w��x�~'�㺎 `�Z�Y*���:m�|>9����<�.�>��ظ�XD�FF���d��kzg'�}��KԀ���}q�>�|�����w.����kϕC�s=_��󌱿~t��ߊ�k.fZ��N����-��v�̹��H�=�*�u�j�����!g9�&�a��S�[^��φ��6̙��Hh&�B��#?H�q�5[�e�#��2ד+n����<WX���6ˬ��Ke��H"��H��{_ޚ<-�\���*��NM�OY����x>���c����+3��/r��e��9���(��>�mm��Q�F���Z���y�p�I{��8DǼ�n5o��q�Jh�;&��W���ە�N���+�ث1^�FG
'i�����,$z��l>߇z�0,}����r���?O�ف�Y>>�;:�-���.�(���&�	T�5��w:���)���n�&Y�!���h�xQR7��Ͼ.�^�����HMjv5�}'�(�L���#��W鲰T�jj]^�3R��د�]R>+uxT�d+�QY�z]^T�5��r.��kC�Kl��0�q^��ah�c��R#s�J��7Ҍ�^��S�ޞ�4���d��'y�^2�#ݺ�v�(M�݅.�R+�`�6�	�����Ãr�6[��	�����q��b�\��2��Hx�N��h�4����rM�H�t}�M�&Ͻm���6�=&<��9扲 ;U�l?��E���<,�-������:U����\�e�&O����T�dM�rü/>Dӫ���Ɨ�/�o~׋k�ko<��(�Ċ3p�$���c�1�t��9�%��ݤN��=x��9o%��Ş��K~�H�����+$>�<oj����xֺ��g��#��5�o*�𞉗�a͌���H��73d�^y�I1w�Wf��;��@�[�W���Ɓ=���v��0��^��{��u���ֳС��z*>v��Ε�ٝפe�����WK)�Q���������ӽ��^��M�!�}l��eV:h�u-wg�8�&@��,��[h�o;tOUU.༩����u��yKU!���F��@�]�W����AE-�G�!2I)�.1�!��]F��cх�Ø������<ܽ{\u��r�r�����i����.Z��ү�[�]?Kky3�o��׋��50�rP�)��p���c*l���6���$"�Gi �>���>P��Dҳ����Do�<��ǹ�U�k^wum���ؙ'z��[k#W�w��_"�.\�a����EN|�����HV��O�f��=��p;/~�k]Sq��(�B��V�t�Ɏ�H='S�A��V>2�:ka,�
1�A��;Xڶ�q�]���[�{��Þdb\��s�o=[��V��<��\6h�2�KU�[�v̇�{�G�`8׏,��/T����N���]�%��\����O�����[��wx�⢊�Ϸ�r܉.�!sh3�)ҽ��Xu�ޙ~�Y��zz؁�?w�U���g�ݢ ����%c�77o�!�b�	0Vlͩ��k�ݨ���([�Ib��2n��B5�J][Mg���@,[��w;k/bæ6���2�e�j�>�����\�rv�jϝNįwg���ʘ�<�S�f��Od�7E�v�>���x�2A����Z�SM�.D�iH�<�ﮮ�M�����;�Bfu�7�)v��k�(�μ�jTw	8&����D�����p��o�e[�ݬW���.$�P8��*��V��}�rc�&�S�jvC�Y��͞��:�Bv|�%.���^��O���gV�d|1`X�C�7��:�ߔ����E�c&*@�j�֮�����Q��G���ҍb:�5f{�N�kA��|aڭ��sG&䑤�m�6�c�SNJJ��qɑU7�/{7a�;w�)}��N��N��ox:������'~z}ضh,f�vvX�V�z��'8��)�~2�v/g���իs(aIn�pƫ�^�twD)��Þ��{���ww���M�{��^{����p��q4�у'
u��C�b.ӍGci��\��<9�2`�ŋq���6���I�\=<p��ڠa^Ӭgn��=.�n^���<�H��N�{cC��{�� !�x��r�Ӵ�m�:�x{)��1q��݆I&���Z��=�۬�vrC;5��N��m��"Z��X�xk���m�q46�V6��v��Gq���w]�=����(��S���r]��_mvy�NX-d�h�e�-Ք��ѳ3��N�j���*��x ��~~|�?�;�w�_�D�N�
�K�s�·'�dz{|�Uz����s�t�C�G�������F�8H:�r�gů���z:A�k�l������;;�>���GUy��ΰ�-��V��o�¡��w>R%)�T(�{~~xY3��$���im9o�ϋB���>Ȧ�Q�ɝ���<�$;jq��~7D�]	���:��"�@A:t�Mo�t_�2��F�#�����ܰL���:;���g_�T���mq��򎓡�f�4��k;���D�r���_y/XQ��&#-4[��n8nA�}�
����u�R�^��n�ً7�H�ÂNޓ��
�v�j��w��lW�zV�^�x(�AF��;%�x���z�4$���l�j34ׂX�Z(�v6�L;Uk��fK��瓭>���W�����ެ�tc꾞^�S�C[c��&^Au�ɛ�k�0��X�x��}�3=�E#tA� �Bc�8}r��h��wϪf���&k=�w�xs����C�>X��z�����3��/�~�4��记v�lQ�پ��y�%:?/VQ�ĥ:�)C��z�
��=�lȵ������Fy�����&kT4o�Xo�Wo��Ca
�oz���|ׄ�����FI+���^]�ם�W�~d"����o�^V�P�w�=��gt#�u ��bv��wP+-���t;���Ӧ����6'�'>qH�-yFL�病_6]��C�/3�ͬ�C�5:4B!wRvh{|ǈ��+W���.o���wM����N��S��B����ɉ��p'>�C��=N����?Ec���V�3�Dr{�jm�3�[�uݤ�^�T���Vu�#1?�"k�6��;��(H8T�p���v��.��u���3��v4LN[��$�6��S�乔�nxmwW4�<����)�;l�@���V�,���ξ��,�[���a�P�:�og���[�^��x���P��>��E�e���JXy���%\alū[�'}{����n���g���}ה5������aCc�K�^5�NF��+��\��5���0�,�Y����B^M���	������e�eM������"U�۵�t�$^�I��f
6��@\�3������1v�����m&{�m���#����ɾ�-�;a�ֳ��`=)KL�o�����M݇��+7_�LB�m��H^�U��?�ڳ���{,����+_uӄZ�����v�Ai)n��/{���D��K��Y�ug�����>y����õ]��Zݡo\"������ꛫ�S��X����b����C��!�HL�?#���z|�����׼�����^W�d�f�¡w ��Dr\��ݫ��źM��*�Ҏn��ww�;�k�eص�4m�e�8���Y�^k2bkn&��8�lp==&��N�fm<I#쓿�x~����&��U9��1?�ǻ/�,{��^��<�~?������r}:H}��y �����>���}�a��/�w��w��������.A�f�ωf�+谢=�9�0�GϞ����/8���W�
Z���'w���Ǌ�eٹX��=�� �d%4$eImK�~�A���ŗ��(�'UWGk��!�f���i�۪�V����a����=�$�dUM=іZ1�J	r/f����[����4n�:9a�օ(F�LUļt+e�V��w��P������'�p��o���^���s�Y6�|h�{~4�}L�f�n��U^&��柘��);9W��M�e~�>	��x{��-T�7`?����'�}�?��~����٘��Ԝ=�̆mHIR'$�:������4/��k�ȗ�P�͸EϸI����S{w��˩����$%��UW5@[A9'�<�в]i�7�o~��yzF��En�+�E{	��ð�wv�ڜm�4<���*b�	�Ơm�$.�
�t�����{�|�]�b�ª�vzT^�bk�Ņ�y�h�V��6��wr����]�V�������r(1ϤNCv� ȥ����dV�W:�\����Ԥ�i��۞��t�8BL�mu�5��ˬڭ��1/�xΝ��=��,.i���v|�?0��77��R���3.����l��}9e��y���'|����s��w(�y�v��|��̬��H��Q�Z���
�r��Z
�v��:���Vy�=��y�R@F�����VmVZ�B��)n��q��x��Tt\�#��r��Wu�<������Nm��|�X�nZ�g��c��7�e��ߟ^�wɲ����2{m�3�诳�/��a���_�k�Ϋ��$.�Y[39h�E��d�����ʘ�ž�u�I�2�ϐͻ==��F�26��¥�w�p~�%�d|�.�M|�:{r�x01��h�E���p��~A�N�S�����m��4bL�m	jҼae$�t�� �(U��ue���K��5��v�*��.ˋ���5ۛ�ρ���5=kΧ�����-�.Xab�KBRh�+�i��Mlj&)u����2)Zˣ16�G�������;�&��<���]eS�9y�8p[���172Ea��t�"��*���;v[��tqT�k	��[���`�:��ݚ�>M�x2��L9��r2�	��me�t;G^Ʌ<�h"m������\b)�����7iw�Q�����{�q���8���}PFVd�z��W �j��-�/�םA��e �I��|�M��A���!�)"@^F��o;'�G���C��Nf�V
?9���r��}6.�3�a�/��e q�C��y�8;�|����Tr���"��>�UƵsǫ����;jN���s��S��z4I���1s��גǞ�;�F��?eoG}B�6d`.f}Y/�L�df(���f������y��E�ϟ���Ӥ��6���@�'���~��NV��=��3s�<']�����Y���<�ZK�gO�O�mq5�y�wpf6;͂D<Y��E�aطaC�^�`�7�	��΅��}������ꐂyl�{�H���L���z%$r\�,Q�z���>���."�maV�5���s.��Q5�XMw;g��
�Z�Au�}D�(��w�xz8<�fdy�Ѩ��!JbE��Mud-(n�?
���-6u.�ȑ)#��󺊵��m��X<�Ǣ���R@\�6eH�����]�!��[��{�uzRE�g��%��^s0�yO!�e�x6
�ާ�pJ�p�!?��^ۏ|
�E��e�cj_u�{��^��X�`ag��v�����{���� ���?EPO��u�C��p��]\n��}KWF����~M������yHgj��N�5�S��^͟�4J����U�uӣ�طN�s��<Yk���q߶.�!D�5��22�r�^#i#�*�|tk��ڽ���P���ܦꁹuET�UFF��N����=�r�#��qZXD�H��L�	�k�.︹�p�ٖ-xm����~~yt �Ӳ�>,���0;}�/��my�ܻ�����~��7����F8g��y?u��2�h�B���+����1��h�e�4+;{�I��l�	�Lux����mع�����@�覥��m�����_3�}�J�If����	�u�:��.W.��I�Q�ѭu,!��1����3�0���lB"-�w�hy�;�����oDW�ɵ`�T(�`GNv}�֐�q��*'�2 ����9�\F�Y�}���qc��ϚT)!H�[��]�Vai`�
�ʤ8���Q$Z�0�4�M�#H���Un�^�K�[�p�����2߯({9�IYB�!NN�X(fB�l�UY�,��|��JD���|ɴ�ZZp+��S�U�K�He����z����tꂓuE�Ed*���OSR��V����ZQ0�b]��U���$.�%�g�]�wyn�^^�gs��U	���;mm嫣�v��Xh�spq��ƒ�u�Q�=��6+�C�g�g��{N=�SsҔs׀��W�F��3�uN����ywrˎ��_hJ%��6c{�����{k�K���ʗt�b��[Jb�9dxd8�&��Y�bj�HhX,�<KƵbdkB��h�z������N%^�hF�#%��j����'�Yz���( �[��z�1�nΓ�gm�e��*����4zV���v�H�X�x�.��=۪��U���,�{G��U5���T2�)�1k��#��0L򻣗P������>$���H�D�o�����y+c����������[���<xO#V5,j��������<����s���9���K����{P�θ6Y4�+�{^�m�r�Z=%:k���Ϧ6۩{A9�}ǐ�l���n+��H�y��W$��1d�����냈�����;}g/g���G�o�`U��s�����]x������,%�,m~\?y.U)hs�:�Gke{`ٕKѓ��0��h$�A��_�O�6w�4�q�̳��$��;c���SE%�7Hw��Ӻ�6�?l%�p��R��_��j���ԯ���^����R��~�ck'n>�~�y��u��vH�{�����4#H�P��ow�T��{�XLq�ׄ���Ky��m��v�R�k{rJ4�]K|K�i~���ޞz�g�l�7�ܶz��x�Ԯ�|�/}%��=��O�-B�>��z��^��,�"��=.�<�����:�k��"��=�蟬)����3k��L�0{�[����w��}�Cih��M��0c��%��*���a��YN����߹t�#>b&��U"�gZ� B��ޞ��^f�ݯyF���{�i]p��^K"(Ojc��rm+�
�hkJłW�u�h�7~-+뎊:X��D��<ӽ��~��%������"D��B���$�{֪f���ܮ�ԓ�:�����I;w%�]}����q��:�X��qB��a�u�=����p��a	����
u�^��U���50Oɉ�J�ƮB"H��V��a��/SS{0���sf���}��޷��b~�����a��DQp/U^y��;�����bFʑ����ƴ�"�h�����p��5�ő	X�`�D�K��x��G5��+Ƣȉp�S�z��%�$��ۋ !Xwh�D��z�KP�Ns��N�+����I8��Yt���։j�Sn"�Y�Z(�]�=T���$	r�&j�BZDq��
�B�4��Y�%O۪�i��Ԭ|�vK}I��o{JȊ#�p��wxZ�Â�҅�v�
W��(�n�9\pbQBJe���V�w��0�.uǟ������H�1	x�����{����,��@��s�$8�:%�ĨP�IX�Wf+3�Ő�4Z(�X��Ȋ"��y߶��F��PB_m���p��r�=;�\$,p�m(��P�s��V�!�+��2,�����O����,F�4�3�����Z�QdE��N����47
{��w�Ӣ�DB&�)"j���!,b�.��1����K��\��ら!+DQ"K�m���{���wJ��̍�O$d����ٸ}�vi��.i2��{ye>�g��譇.P梂�]�#-T}ꧤ�;
�P���[kh�w-�'"#U��\,٪��_J�Iˊ*!D����#�s���9��>�����J;ƔP��;���IJ�2�2�UM�%wg�Ӿ��k��.���,��BV.��EKII
�Q7���
��aB�#�I��ۯ;�DX�K�"(K)�@�*�wD�'�3���[K�Z��8�Tܞz�jy��:^�\M�)Y�����fp65�&�ԃp���M�3�;��ɂ�p�rmN����-�ME�O��X1%��"E�4�Jk��H!+"#HJ[��o|���w=>=؉F�{�,F����o�B�N��DI+ώNwe��iߦ�/.fBf�*uά,":E���a�h�B�s=�q8K��k�7��='R����( +�2�gfr#}�RBZ$�H�	I�Z$�w|Z��Rࣂ���$H�
+��w5�	h����u;�E$#\.M���r��P�EP��.�n�rtBXB��J�BR1+�B�=}�M�\�)5"�X�7�A�'��$���]�tQ�
�Y��k��zW�.��i,����2��#�d±B�Dosح.	-W�IP����K�'�ח��AM���M���>D.
&�y�V$���};�~��F�-DW'z\B�Gu��P�V(S�O��3�sj8(t��t��JIm&%'B�=�."H�	H�ܕ�%B�k%�u�<+C";7͛�^�X�I�HJH{�u۔T�D���S�T�#Ew)Q
H�$v�ޛ����:K�h�2�i�j9sf<����D���[#,�.����q�fʟ��)�)넼��ڈ�وZ%�JJ�BV��$B�^x��}���
�%7مdt�$X_����<��9I���'������~��ġs���HW Η��bg�E5�&Zw�����8~�9�z����^�7tE�Y��l|�#ve7��v�y�0f�'9^�Y��[��n�����hB�;B�A�ˮcw1��b��.NX�;@�ܧk"c@8��̼�A�Ŵ���be���X.]364FЗ;��<4&�Ep�JA�eڽ����t�p��%�[r�덫��J��\�ȏ�p�fWu��=�k��p��w���u�\n7NV�m�[k��^hۑ:���jl1֍��i���
T�8e���3C��
��m�K��ܐ h4�ی�RT�T�$�""cmB�DE��]�>.��.	�R�����O3�w�Z�$pY�%bQf�*�<�jD����*}ԨdB��+!�'�8(O��v��#&뗂��P������5(�CQ���^zIrwy��TX�"X)��v�h���2�{��{��A*���\�J��)�	�;~.!o=uDB�(�R�)p�}�ͪ3��B���0V(\�Es3����J8(���﯇v�.��q"TB�r~��\��ˉ���y=���U�FΚ(�=�^�EW8Z�#En� !0"9./���0���M�>4B[n��߸�7��b8(�7\%�5��j	��!r�\!P�I{ٸ��
�	M��,�s�s�}�6275���I!q�|N���B*�~�}�W�m��
&��u�L�ξg� x����@����d)�sU��x�!Q��H��	�L(�m�URmDH�I-{���+� �~pr��3��D+]�Km������������b�V.r�{�y结�ta�D�H[�{��4�b��D����حgbgO��;�k��\#�VR!3
H禼\(��R(]�d)�狅>q�.	+z]r��Ih�K}���;=��@^���u�;e��WXo��B�}sX�6L[�n8��j�eR�Jʦt[��K���aq�)�'��l,�y&�}���7���/�:V�q�p����&%b�^�jW�H�e�!Eq�{s����S��w�;%uP��G���0K9��]wf�KM!Yb���yn�.��j��DwryxB�y퓅��9����c��^X�ݝ޳�ohbٯ�C�w�M�	��R2������V�*�A��JW?!���<�m�|�y����9sw��W^��!���YW*0�,��ķݿ\(��"]"�kD��rm+"��!YWɅ�
	C���aH�ݵ�>��c����-�Y
�p������fTsos�Yruք�RBR1/u����j͗+�
V%�$�"�=����K�N0LK���5_����4���e%}�����=n(���*ӄ�Iv��-z�Q��D�D1%$׫���_��+2a��{��ɯ/�?B-��C������@5
��ZW�ۊB��)!+�o�����m-�I �tCo�C7+�Ҧ�@K�߽��B�W�gOlI�W�ie4�G�6Dv�pV+"�'R�S2�M�USTZ�r@%"�j��n�^�Ė�L�����I<���{��]Kk���pI�u�j��B���Z�-�bT*֬��"�w�iiB�yc�)�1%��6�\��V�Ƃ��m�ک�i��.�$fK*�2�X�]U�H	�aR�VY�03ˮ�hMU�j8E�ryg��N6{d�����3J!*!{��4QbW�f���R��t�imp��9�ኟ��qm.����"E�i^�B�C��;�Bg�G�2�;��x'"��$1$��x��J���v�����gKNM>�;���Co�%�#��.
��;�p]ޫY�L%B[֨QX���ee��G�-8��`B�D�.߹����$!���u��9�q"�o�I�$*)�fj�U	iF�'�sd+�>��ju��Div�P���ܬ�w	�%�*��oǵ9���+R��y�j!�{�euK�-�6Q~��:%M���:�
Y�j��9�.~�1�w�y�f�7=9�����n�9�����0A��R�g|\�j9�Y
Żsc#3���ܙI�����FE뫄������&�*B��H4R!a
��)^��W��ٝUN�\��Z.�۟g7����#n�1*!)$^��k��?��"�Gu�7���^$��W��e�s����O";^��d.y��NB���t�w��������r��K���-#M(��&L]�W��X$���4�G�N��9�R���ܿ:Y��K{� �",�����k�-*}ʈ�<G�5��6�t����[sh�dOfb|���4O����EQ���$a8�cmuղ����mW���8g�K��]�����h�d�Ts�[���\��'לגoۜ,������i�ESQ�xB�/	T�]��f���?=��y>����\o2_/9�
}���r��-Y"���b����	�y���κ����;f��I��ydd��EG�b�4���j�I��e���I[��Ȣ��J���j�We2,����4KH[n=�s�'T1�"�GPiu ��u�?x�����'����)��߻�#M"�dVh��L("luE��H	�N�mĜָr�{�f��q�p	I-+�U�sK�\D����񐨊���Zx���%s#���)m�)_}�U��&�b�8��Jťy[�oɮ��[�G��'������޷��ߩ�I�]����r���`�S�*��"q������r:pTG��Un%{��"�X�����K�a �����Ur�����m��v�zޞ[��9�p�$˾C��ڼP�)ݓ�W=�nz��S�ԓ.�A�n�����h�(����28C/�0��$+��$�ɡ9�C*��B��,Q[�(�x3=�c���Jh�t� MT�M�9]~����OH�d�<G;7���'F��b�TDs�w��M̐���beDI�}9���p��=���M*�C��K\�ݛ��Ȕ����ˍ���F��du�n&괺��7��|���B�[)���_[VF	H��ib��s��z��./�#�TF�*"(%����ٛ��~�s��I #���ط���Tt�"H�]��U$6�	��NCC�Mf������!��:��f�f<�;��] ��?
?iν6�hvY
��5�����N!I
���ۚ����>��s9�"�y�q��\���K	�PQ�z���f�cJ�\��kޝ���Iaf�j'���e?.���o�I%ʿb�G^�O]	QE�۪�:�Βu-�k�d�g�u�,��*l��/ƕx=�n���+��z0��=����\�,~R�� �_�d^����#�vB�N7��W
�>mZ7��Xi�}�N�Ȓ��1�y�˻�k��QƓ�W}��#��2FOd���{ߝ���vf,�/حF	&`��lVL�"�gT�ȹ��ܷ��fؠ3�OV�"����I��eGg�TE�چB�v��{�UN7��Z-ӏVI7����s�����?Nك��?��{��Q����`ZZ���r�a��y��o��L9C���?$�>A����z1n������&EOṿ���=���:y�)w1<�OJ����5{��s����f'��%������RM���I�v��v�mkñJ�$2�y���!V�WW��J�	s���|/I�����:7�݁Q��;Z��l��KX�����K�]��K��r�Hݨ�,�NYVұ.�F�a-n9�ح��ay�\�B����M��=�ǡ���;�	�����>\;VH���"��M��!��Wss���DDv���Qn�+j�B�t@�c
J�Fs�>��I��ZU�}6����	_>�?wex�1�*������Ng{��Gk|�->�mimH��h�_s�EN,����{J����U-�ҩ�sA��H](�2�QF'�>qb�a�,�ڕw:�E���Qh���7�ݘ����_]"��V{U���"R2=��Qj�|x�޼�򶗯��* ��/�^��]s�v9o|,��h�>�����X&l����F���Q�)]��^4Jo���O:�_�����s�����/��TM��.k�ґ`�{���1����w��eWKpL���N��˟B4F����8�]�x�-����j��*U�B]����}����T>����sT®s<ZU�J���Q����=�sua�3��	YJ���n��uy��gW&ef�o|��v���]�'<�ޛ�5�1RՑb�5y��{=�Ƈ̞ZY$>4|���f5^��W�&)���$F���Z�H�jȢW\P���_&f��E�h۪47Ba��u�*�M%]��mGX�t����ڃ�ɡ?�e�ԬpKP�j����7�E.��k��ɸ�F��=j��i8'6�ϵ�Zh��[9[W��B�z���,�79[}���V�4��U٪J�W���N������0B�m)�
p�Eպ?V��Q�@J��VkϢ�����}�|.s�����m��;/&��z�����o17�q�L �J�r��3=螦�ؑB�吮�a^,�'@5�S��~;���#��o�[���ʩ����'�P�'��B[�aB\�N7to�}���ݛE�-�F�3=�9k5@&]�������=�ԝ�{��udIo}����Ӏ�O�=�Z{���/�x���lM���3*�?~{ܾ-.6��$m0�g���Q"�MAs�lqqD��P�!�� H�UN-n��K�2�7_���ދD�����2ܥ���Z�^��M5^���ޥ7�~��vf����?D����c��kJȆ*"E��'}��D�Tꉗ3EMU���͚Ÿ��oű	h����o��w��Es��%OiWZ�J��b�R,�K�*���׷Tڙ�SN��\���<�P��+hG{s=�w�o�yϸ[:�q��
8�.���+��r[�,Jۭˊ�sp���Wmf�1����Xܔꗣ�R�J��I�����j�w+���°D^���Ғ(RM5D>�|K��/V�P<+f�@�YE�۫�w7?����p�=ߏ�Xa�c�91��7FS��}����Ku��u�����{N���۴�0�Dab�Ug���v��ցG��~g��z�����$#�n����,/1v���h/��jԂK����=f��ll�q��֟1p�5J)�zs)Ic"�~�ՙ����b�|_�`[�ɛ�w9h�l��]�dJ�l�Nq�o�����#ag��n�rl;ޫ$�w�dp��o���2������.��w;����y�ц[T�[u��S~����Ш�H�.�Ã�H�MHB.�<s^g�\�͞�;[;�b؊;�=�V��5JY&����}�?}EJ?�QӘ~n��YH(%�N
lvo��!���4�/w��Ӣ�� �\��0���Ks�=R{���ݮ�w}�����e��8��}Ր�OyǈVE+t�b�^�${�[U*�v_�}�r\aZ�!�.���|#�tUM)Gj��w��6%"L����B����'
�4�R
���ˮ�pr&�7n{�������zC��d��ώ]��h�Ȅ)2�O�����T@�ZD�Y�q^�:��jv*#wE1���w�MM������}b��yٞ������He&DL��%��gܭb�OGG����cr���Le�����N��/�axõ�'}4�q�ّÎ�OD��)����VIx� ��V��ٕI�Ų�C��{wE���֔��\�7%��fZ1T�s�}}ǰgi�8xp8H$�{/��{�m}�%�5����y�	��ƯgyN�i�v�/�����̫/�0���D��U���ck:}v�[y�+ȧ$�!�'pg��\-)���ϵ�釨�3wxV�7�J!�Fu��'Lk�?%l�*�sL�n�5�r��1lkTW���ںk�N �g��R�x�v|q���YE_}K�˂jw���~Qn����L��*oɗ�V��Ŀ����޽֝a8���=�o�k�Pj7�w֏��ŕ�!"��m��Zm�Ct�T���
�+�x2y�*����`��O���".WUgo3�U㾿U
�+%��bպi�����ޖ���h�	��<F;,���Ũ�K^tfv��u��#.)����D��Tg�ÿ������s{���x�!ސ�F��oTĪ�I<PN#�e�%˻6g��"\YT�in
2���Jf�d��0d��r��2!#g�+��:��f������J"���y}/}�U�����ۜ7>&�ƮZ��w,�#��Ȱ�X>�B�y��]0E!*8K�'!��`����ҏ?_%c9J0�m�V9��#^�7��8'�v�$�w�^��S{wB�x"T��l��,4'�L'"^X�R�����2�t��3T��ߛ�lK;����r��H4/syͮ>�b�7�շfH���T����z� 0%	����$�O�'��/�9Dg���O�0ֿ,E�T1]�U�Xu*E�7Y|�+w�US+��!DG����
"?����
"?�DD(�Q�"!DB���""D(���"!DB���
"D~��!DG�DDB���""D(����!DG�"D(��DD(�Q�"!DB��Q�!DG��TDB�����Q�#�Q
"D~��!DG�
"D��Q�#��!DG�����)���p� Mq��8(���1]��P5ZM(  ��h    :�4 t  �t��;�� t�� 
t  � �(R�U(""J

�� (�)J
�
$RJ�RJR*Q%H�E!P*��E
$�	DH��H��0�$�)*!H E���M�o<}n[.�}�����{y�������}��_n溫�y�׮�G��"�6}���iﷄ�m��m������G�ﳾ�S���{�e.���֘�֖1[2-���ku��ZJW����>��2��1�})@}���������n]�]y�w��}�;g�n�_c�n��vl��RD�^�]TO�a������:��W.�{�z��57׹����r����m	�6o�*E�I"TUϞA69��|��۳m��{��s{v���u��;o�v{c�Ϣ�/z�Z�����}ƨ���ۺ�����G�oB��]�>
��{t}�Gϳ��c���[0�1E������s���I����US���;���EQ���oӵ�E�s��J�g��Rp�������`W�>�-�z}�}���I�)�J��|�T
U��)PD^��Q�k��J�z4��(E[��(���IR�
w��������X�<��m��f��ꩶ*��� ��/g��c�m�/���u+fZ��6�kU|�UU^�y��A}�{ґ'����f�����6��^0�;5q=�<�Ȣx��8��k������lz����}ݕﳡ@^��jD�j<�*�J�$IJ� �  �;�  <� >���|� �>��X  ��U� >��n{�  >C����` =��X  �]�U(xE 2ϰ �g��J�P�UR��}`
(q��  s���@ t��� �� >���� }�ް� ��}��U| �b���y �������  w�1lШ�[l��R�$TU)BE	*R�  �ݟJQ���� ����}�@�[]�}= |���*<W����Ϧ�G���^�-�1���o�y�{۠S���%�}�Oyܯ��`�ϠJ��ʣ�}Š
 |Z6 (=� �^ P� }����|� ^X {�u� <��>}�ڊ$���J�M׶��{8��wm<�Er�N��y�s�����8)�"eJ� �@T���J��� ��2O*�)��  D�2�S	*   y�R�h0�0�%*��z��C�?���C?�C��R/������G���~�^�gns��Ί�"��� *��UN���� UT*�*�*�����` UB��� UP��ހ��UQ� �TU��}���ҟ�0n<R�v�Ӈ'J��.�-X�u�� ��k�N3�\��j҈�Ƹ��v���xg��Cy��xw[䱑�=�)��`=�W=8H|*=���`aO��M���(0����a{���l�*L���:A�(+A;+�?��ނ�����}܌�a���ކ���k�$��K�5]�z,�:p�ow�����=�$X�FI����M�ݝ�� 2��+@%�	ÜM���ⓧ\���C���Z&u��%����ّ5ݺPv��4���#���ŲvÇ�s� ��^v���FǪ��ӵ&K�c�U��r�?I={��w����+T�!{�Չq��,b�㡦s��:G{�160��]��luP��.�`5ð��o3�M�jgJ�nɪ�HE��O��V�3�Ķ�zUt��u�/�M�v�i?v׽���(+���	�s��l@+C���T_X*�����}������/z����X�=�^�'j58�X ��S�1�Gz�\�@! #A��o3w�4��K��w��g�Uj�)���sf&��F��/�v�^5�C�	�N�9��L�NLG��^�ǚ''0�Þ~����"�d�_*^]�1'J��"A���#�����9���^��
Ov�Y�s�H�c܋C�d���}8�����/�^�<���L��	㣚�c�{���
3wlsO���������u5�*X��%�L�i�;��]Kr���5��;@pm'/v��^����0�%�w��,e|���V�������p��Py�0�ĊF���w�0�R�a#Bѡ"˧x��v�qD�ti�$ɗ����F6��XԹp�t���Y�.3�y^;22�1�Ӭ�d����Wt����K��WT
��p�:�ڤ�b��F@Gg�j��4;z�ݛ��gK���h*����A�C���u50^��=y�1�N"�]���	��ekEkz���`�1w'MqW��Nɕ��2������<Z1oj�j��,˃{`[_s�N�ys���x]�-we8�I�R�Pޝ؆�xlB!����h����2���'���l���y	�O-�u�;���;"o%�1l#��bs�խ��Z/M�(�)8�����������j��-%N֮��Nl�����H�v�(<gV�]���:��Ü��l���㼹5�90@_�>Nq�sM��	r�HWR�/�#\n��=�:ձ AG�t�^����Ɩ��N����Ϋ�� w����$�c�0�}���t���3b\
T(�N�������lή��密���B�O9S[�Υ����s&@>��]�j�s�GhO{�����C��r�g����~�I��}on�]�7��Խ�m��=|���3R a�L&�i=�%�tM,r�l���t8q��7�!�)�6c��z�-,/t�B�\�xSp��7�������s�M�C��ô�/�Ev��s�V�i�'�9l���{�ܖ)6�m�������p�f�8ܿ�vr��#spp�;OB2��dܰ\܂$W �2�GFr=v��s��j�.D6������žq�A3��1�0�k^(V�$pS�͕��Գs^*{Sûp;�C0�R��{�����5�yn��Q�lڹ��yn�p�"����i�\ޅ7�xL�n2�OY�6)�B���0=>&�� ��K���1�Ԟ�%�}�n�T����7$������o�硫̨��e�[�q��v�zr�es`�&ΐ�����nAڠ]�tL���<`[F#��aCtͦiA�a�=>���û.p�7)cY{��������V�l݂�%�.9���|'n�S��Θk�&�a��	�Zz����ݼ��w6ㆡn���	!յC�8.)��zV�h ���L;��<�y����! ����6�j������M�(�0HJ)ǹ��.�74��$[��h�ލ����	gM9M�'\rq�So�7��޲����i=�ɩ�h�'��ش�p���YNt�,#"��0�/NO^/>�^��n]�p�	���Ф�t5��r��b���� U}3z��ǜ�����:l�#�p�|P/r���X�O;|XO�=�blWy1�k�6�o��ʳq���mzK�'9���F�KG=[�Zҵ��P�ɺŵ�ݦ]�� Q,s�'r�2��넥hX�l�%b���v�.HOɋ��q���Uz9�o����U��)��!�8���k�F�l;S�Wy��o;�0�t��hޅ�9M�`�7v�q�,�<x���KQ��اh��B�/o;�f�ĳ��9��;;�O9���ܡ��o	R�����gx�q7�qi�{�G��/���P�u��D��O��U�B��S�Tc��;�P?n�����P;_q����Nnӡ�{�8�V���R����_*B2�nr�F�\5"#�Po!lT�Rf�jZw��e���ū~2mʶ_l�<�0����m!������*A:���|���9{	|�7/F��'��Hs�T5�k��
Y�7\5�R���wnlK�[�p"��M�V���$9dHk@�'�с��,HUO�ˉ~���tC�����,v�%��+.���7�])�v+�9���������Ծ��[�gf��/'}�����Ӹgl�ۘn�5��wW��á�b8�����9N��&L���Ԟ�9��W�w�Ԍz����	ط�\�NU��f�BLV��;�\��i�Ww,����c9l;���uQŗ��4�U�n�?3L+�J޹0=ʂ.���72��7��t��n����q�#q��{`�k���_���b���if����Z�Ѱ�pl� qr�fi��� ¨��YE<y0��s��w{ SMb�15)T�tvN#6DR�H4-�ӧ�R!^¡���;��zқ	�bYx����ǋ���A��F��<8�L׳xt�+9ћܽ0jїCxN�čx}r��T�xL%� �B��up��;�Vk{zՇ6<=KŚ����`�U�2�nl	��\���� G�j�`�+��f�h�d��(�ʓ���s�wJGuh#:99��s��MQ�g7�*�hk��N� �sҨZF,��B�K����u�溙N[��LS��p��jFp����R��"�Z��es8Ѻ��q�&ad�J�k�������g{4ߎI�����ķ@'x̚W=Ntȹ9�j��gxB5u��z������n���&#IF��8�I�)Ɂ��SV�`qgk��'NS�f�$��i���h8���J�z�*9r�R��\'�o,�3L�K��NC{�C�ũ���8ҝ�%�����T��ꮲ���x���ݒ��:r�|jYۥ��5i�2l��89C�*']B輔��~�8�@������M��Gf�J^��G;ς��]O��8� ��Z�r����N&i[)�U�H�8Y�k��+���{g�]��?��W��,��b�>다�oc�%�f��S��y`�mޑ"o刈��v%��b4�Y�\e�O��򢡪$���m������{��1\X&Qjk&��&q�t��o�1��qps��f1n�w������s�a���裭�a���bƜ���-��t^<�ev�[���8�؁�m�Ʊ�,�k�Z�S�#c1Z\�S���<����.��V��wG��	nu��];����~�q�j$q��Ey��#(�x7U9��^Xz=�赱qLI�F�A�!���I]Frx�O�ڒ�<mOW`��۵�w�qY�g2��y� �aF��˒�l*�ߺ�\�ɛ;��:.�q�zXہ��r�yL"�w�콠	`�#[w;���yES%�ytn2�.p���c$�.�"�cRs.�27�`��a��h\�RLP�0�0 +��w@�x��l�]���5v��9�tl�]�'&<�+G�p�ϩ3��	�99v��뗑��r5���E��aF^|	��u����l���7��' q<��� ��c�w���n��wt��J��L�X1і���������cV<`�7�����Ҭ[�L��Fl�p�|8sNL��W�T�(��[�i��mBP��S�Oy�=n�q!M���Ҥ��e ��3Vp)���P��⳷��ޝp����=�R�\����/�3�[�`:�����7_r�2��w)��,�޽VV3���c�i��Z\Մr�D�t�F������ �Y�yM?0QnI�jѶ�@m����ʚ��@С�:{�v>cB�P!ba.�^�-��<��Y�+���sӱpm�$���i�E��%�3"^Q�5`��!��^&>����&x}'�ÆP���ۜ������2
.*�H�ٺJ��1���Æ�b瓳Cq?���=iY�j�Z�ܽ^ْv�aĐ��{�v<�*���1�5�W=����fl����|�G��>��k^�K�����v�ܼ�D��c+:�ӽqޟ���4n��6R��
 ����
un^�,��ׁjv/É���*�#�41�����q���p���R����  2�`���)�n�7��p;���8�Y"�KoL!aw�v�Bn�q����)���J\���6^yU�9;)TG�'*�F�h��tZ�0���[0�&֥�U�	I�꽳�[��@؛鋿* ��%ϦMsV�qD��If�,Z�� *��Ʉ�'�xz��_wN���	�&�H#����(tj��oVN�n�VZشP�3��6�!�B�ob�U�e��CA����	R�ghƓH4�Y�"�0F6�9�5m����ӹM+T�+E�X��/4�y���ofOΚ�Y���;k.�09��4�[ږI�w���	�t�1˜4�)�Z97 �.۫{k�]����H�G�v����rs[�D����e��=r�F��	ħ�L����ޛ�8Ü�n���;���=(��8L\K�����0U�NB��tbȷz�C-����-�	�䄩b/���X���^V�j2c� 38oQ�=o��1ǢnscA���д�Ǉg.�Y��wI���vP�o�+r��g��r��0��#R������Y��p �r�'�u9��f�U�Z�6�A 1!�nl<�7Q��y#gQ{�uI��]��(����7X�sT[g�Pz��|��O���n	oMk4�suf��v�^���X[ӱ�Yn��p�ݦ
~���^�r����h��sg�gE[˓�È�ݵ�R�z�x�D.:���7�n�
�	{�1n^d�t�	|��Y�J�o#t5�ٓn'K��>��$ap���"�O8,����n{u�=o��p���k6���d�"~���L/�3wK�o1A���6��O����a�i��8)c�tѕ�]ۼ�3JZ���۪�&��#W^$=��"����:N�L�y#�7�����#���m�f�����˙�A��X���;&N��Z�Z�c!9խ�:+N��a�0m��Ϳ�u�����tݣY����~IuWw��:����yV��7��q���oJvwߕ0�f��8�����-�r/*���.�݄�I��Cnx�w7N3�E��S� ��*8����"&y^�7�^hw@Y�;��X����V�������&��,'8�MY�s�k���U��n#�-R��:I�{M��t���`�&(2~�� #��>����M��śrĪ�n�����؊ˁ�D4m����#����e�QڵbB3�@X `^Y��s�bgLo��C�=����7x�.�f���ٝ���i՜чב&4ыl�~@�0�Qw���,�Xz��Чv�a�C��L��P���z�����G�[�^ɈI!m����10��������X��@�����"�,`�%"��Ǫ)	۵�\͵u��q8)��w<&M�˶d��<N�����6��Tf��N0z��1N��l��m
ί{Y7�l`]$8ރ��of�he��ܨ=p��*P!guRn�K5�i���j�:�,�_r:;,�����T�l� 56�ۉ%L�Ƃ��fU�F����uk��e�ƀ���;-������g9�@����q�ΐ�D��Ay�/Mjq{Wg����f��v��G	F�-+�ke��(^�lבE�ܓ�ӜF8�[+�XwEƨ��]�f�.������lZU��.r\:f�k�g.�7 �i��7.i,q��l7&�Z��_����vl9%].���tP��-�o�~�{�On�F@�l��5 ���f�
�\��=�L���o3 q���zz�����,Ɠ�kK/5��Ķ�'��l@�[|��d���@e����S��fx�z��.�
ۅ�޺�"1��-��l�M}ԽѤP�N͸/��Cw;�]�p��> B��"���sl��œM��:�7�o<n�K`��͙wnp�:`�T� ��pSI�!��OB��1sƫ�8��WQ�\9̀(�N��u�-��x:�n���Kx����Ht)�G@j���Z�z!XҴ&� t��u`G\K;�9n�v,����]���7�X�������t��6�c:��4gXyb7r���ъ���"V7��:��j�9t]��Qѽ-�,��5��'�}O#F����ʥP����B�B���*��m���ӫ�L�%[��m���;�m��V�gf��"�uJ�J����)�
�����F��quة݉�V�����T�C�vͼ�S���-X��۲L�C�
]�.x��ƋV�g$vT���<:��H4��r��ͷb�� [�����4�,bLm��j,V�r���}�E�M]k5������<a�Eq�[\��ܢO��KY��F���ϗ=�i�HQ��ů]�{�w\���3���Hc����,�0G�>��1q$V-�����+����k�lbNfIj�I���Z�P��i��\+%�I��N8�g�u[���g��L;&\ܶE�����s��0��u3�be�L�CB ��2��p�&���� ݭ3��<tE��c��v|�s�WZu�ȖLm���=;I��V̑����A��#��˗���Jg=x��]L��k�BZ��%�UZ�u/Wk�W��g�������݁Iy*��t�4��h�0:h��&TٻcB��c]�D��YI;>�la\�{e�V8�ͫ��n�[5<�󃥬3&�a��F�WP-q�qg��3�n�te���3ٛ��9mv�[����7OT��)V]e���*,����d�v���nӷ*S�w]�G�<ɑ*�<�E��)�K.[@u�k�K��7X*��ogn�8����l�sMu�N}�Ӗ@���a�{n�d|]8���$.ȶ:XU�5)�͛D�ճ1�̈r���۴�۴)x�ĵò��,&πv��(�ɗ��+|��J�vjK9��{a��\/=��H��m'b���-��廧�(��,:jfn����3]p6E���sxu�aJ.*0Ҍ3e f���n��CrNy��\:l�w�i��A�j�m"��`�K��b�[��^�Cv����ck���l9����:�=q7X��U7L�v�1�3j����v<o+�NH|���"hv⮎:�Y��<q�×1j�v����4��:�]1V�lm�#�e�.�Yk��u)��cۭ��f� �'Xt	��#�� �[D�`��;)�n�1��=�$p�t���]��w`M�@�b�D�8+��9����g�[f��g�U��kn�#�f��l��kp�e���K�.�����jLEmc�[�m��nA�����1��LOBϋ!ƚ���Kt�ʋ�8�ĵ+jv�gg�+[��ֽ�i�uwT	;\<>x+ť��p)�y8c׭�4kԅ��k�a^ ���14(���:�i�Chº�&���䫛5���;28����/�e���;��.P��ݞ��YY:��v6�#q�3�:�k�#�"�g[@��:z�X�mv=p�:p�nx��4���Ƈ3�	�C�>��ծ�XNE��bR���sV5�'�s�ܤ�Lc��^�'��Tl��<q�[j��w@i��Z�4�:�]�Z�q���S��M��O*ݣV덌)�穸 ��v;nFY���L�Z�Ԙ��m�s��i��؅��*�pY]�ЛFѶ��vș'K�v�xwTȏQ���#��Vt�Fk��#���k�FW�Iué5V�܃�c+F�;�+�tyɇ' A�k�<�ݮ���״uɪ�Lpe�Bn%9튰cv�sAm�م�Rh��ۣ�؆6�s�g#m\1����k�^�C���!bĐM�k���H��]S��,�>K�ϓ���Q-��p�v{<�Ս����ۓ/n��6Z����WG[˶�j�kn�f#�y�q���	���6���<�g��c�ƴ��g�b�<<�:��q�
��v�Np<h��P{��nL�^�㪟s�pV����l��-�B��3XfVjE�mm���gӓ�k�x��ޘ�F�pqhK4Inst���)Һ��hV&c�R�B�kn4=�a6�.�\��k��`�Z8v�H�e]z9�sŻ�I��c�Ƽ��kq�!�s��`g�p��Q�`�D\Ӯr��t�ە+\Mes���S-,5#,ɱѹ���<�%�� C����$�����kM8���x�s�ZN]��OgOb�P�f�oc�N��pQ�:^����?=ǋ�Om��k$�	�<[H�[u����P%��h�L�ǞU������p��nD#���J�q%�&mY�S��;F�ڦ΋�XabH�4��Ŕ�i�ֶl�����6	yD�G�Y��9b;Ny�L=�5�K�X�n1�
�c��n�^$�w/A*���r��?����=<)n���c6Ό��	I��N�u��.�������<>�t�7��m�h'n 6v���]E2�;�*T�"yT�-[Chۖ�s.�*e�u�;�燵�"�6{]v�gGmϻ8�mH��2���W]��W�:.��&�c��5Ŏ�%��䭺��5�wl�X�B�6P��-9��aX��Gq��%�f�sv�
niĆ\�E9�e�iN̸�ҽ��e�[\v�h�={z�ڄөMہ!�/\Ё�˦6�a��Iyfĕ����GO.%|�ト�\$��v����y!Ҏsc+�*-c�mi���(k�Y�y��_<�Z����<���8�(�j-G���حt/i_U���[ƈ�^z36�4�-e[n8쁉���٘�����ʵ��z�*�\���E�n���vV��姐��GQ*c�oE�����ׂMʾwB<dzۣ�ۋiCu���v4��Vm�ve��u�V�0��Sݭ�.LF�\o_/��g��r5;ȮڮLZ6�$���(f:h�^�"��e�)��-�Y3�Eۛr;[R8�ٔ�UN�$�6l�.&��s�<z��]Q֠C��{[m]����wCBa���J�)<�
Ǳ	 �͕���x���<�.��ƽw���y�v��.˻a�V$C:X�su�֥�lwh�K� ����V�}�9�A��簄�]a�"� b,���a�P�(R�[�5	cC;��d��f��J.��w���/t�]�Wm�/��]����y����;��-l���R�6�S��r�Z��,����z��ןV��3��m�)���U� x�ɲ��$;XBWF�����f�N.Ơ��S)�Vk�9�lr�l��a5�gKZ�k-s�Yr�bD��C;Jj�FYJ$R�hWvn��D�{�x��Mf���^����W�z�Vf��9�35v6�ڌW��âk{Z4�:܁7��N����=� �&���n^����MHY��Jg.6���M/gû;�兙8���Np�Q����`N,vꢠͳ8�0a�Z.#��f��h��<J�ܶˆR5�����/2�Ƶ��z	��
��	Q.3��.�&�wB5ܶ��K6�lct��v�E\���
�����=��!�ܞ׍��\���8/\���t�<�#e#��=��tv�E[�<qB6]��a��^�����l��c��Y#$�v�RZcX�m ͂�T�0��ɓ/<��"�[-����rf�k�g�p��m��v!C��y󗋱����&�̗���C8IRu	�+sr�����;�O��ݦs��l��q*���X��DW:j��o1ë��a(��P� \�6����Ʈ�&�:e�i�i3j�2cOs,<��*��9!�L`�M�۶UD�f��-����Hf�)t<NYv8hz:�kh�&�m�v�n�l��dUp�q
t������Ӷ3�H�I�\���r�=6#أ�΁gɚ���lo/*8u!nu�;�{V.�$SS6��6�J�+�l*��vzۯn&�Sn:��3*�%�S\J��Q��1�����{mGK�]''��rT�A9a(R�������i�sq�g	A�k�l�zⓔ��؊���ޭW��ֹ��۵԰k/m��	-5a���Bl��e`S���s5�Ų�5Yx�N�Ye�(2ŪjYbE{[my�gL�D5׳a�\f<i�2�e8�H��A�͂�eI�bl�q),Z��W�^L�N����v�����:�n" x��=�9:��^���"��n�¸��m��,�m����F���Ыzm�o�M�p(�wO'E���tq;em�y.�jB�n�N{+!a=:wԌ�[mi*=u��#�u����K�u��ysz�E�4Wu<wk�݆���v˺��f�ӱq��v���6Q�9����6�Sۄm�ⵄ֍�R�eM&jJ�4�*�a-�j٥a��6���u=�+�Oc^�v{]���6��,���Z!Sf��;nR
��lʻ��-0�S�1J�K�lc!v���l�6�V�r�[>sm�fj�eq[��3��)�г�t�s�����x��'Y5�h.|���̨kn���\��.w4=!��.�K���ms�9"�������&��q����m��Kݷ	���Cp�U�Q�A�e�F��9�쵍�x�Yv�Y��GWQ]�L:�Ð��wA���t��Ms��Z�K��Ttjˑl��RR��bJYL��Y�K������Ϋ���UT���y6W�p��9�	K���֭Lu�ns�t���6�Y�;ګ��
gY�ԛk��͵bE�`Ζ�;q��4۹�T����r:xh�C#��Ok���Tz�>�.wI�p⬼Kv�<�Ny��%	m5\��4ȴ�	E�!4+��#3�	��+�1��m����Ƙ���]>�'�nu+�����j�۝o=�v)zn���d�Ŕ�fŰ'����#�+�k�a�;s4�h@+\˥ԡ���
�T�����}�nN�7mm74)v�3��_��Y��4�s(�[��hmk
\	��8G�����I��mѱ(jf�����,Z2�V���b�J�`yi�=�;�/9{VK��|O����u�y{.�ܮ�����me�����Ȕ��\�|6�4[a<�Y��_-��*Gu��ru��A���[��E�.��2ׇSBX���JXha�]Iz�mas���0���ॖ�SYb�`ٙ�����s�=*.�t�����ug�g�^��؛v�v����&��+p[vk*7DH0��@B�
���b��T (UW�� ��TE
b��������kT�8�j����3Š'�^�75��/mث��`�'�`�v�Ш�s6΋�㳣rQ4[��)��H��c��q*+	���ň�;���
�ə���*���`���9g=7k9Z6���C)�����P�l�v���wV���5)6◮T �1�7b��Ocr�롱��X�jS�Ku��b6�vv�4�;u���wL�E�	�ⴥ�8nq�T�n���%��n��Y�n42�h.#55al��p�qv�{r���D̉�����`������2��i����Ї6cå<vf�n��"��=]��F彉y�SrH.s1�V�Dx厇A��;u]���2����׫V���uV�2��+.��Ta�4.�К��MnJFV���S�+�v[R��]w5n�ʝ\��g"�kZ�i�;t��#�h7���koi,l(L$%�=���y�IJ���$�M[��Þl;���^�y5.��2�&������݀�4qc[�t�!��Z�V�'��+�]�w���웛,��x��f	������˫'[��c���<�h,plg��1�,��Hh�c�l%��p�l�``������z�l�X�{0s]����ܦ�(l��N�tx �˷$�!���ʙ�f+�5b�hi��Ra�����u�!u�k�p����[�켱��XK���7>���i9��;;:;�	��3u8���@y�9V�0��k�=��@�s�֖�FьY��.�V�8�b\��eR[5�8���$�j��.�F�r�bZcbie���CDs�`�y�ƭ��t��Q��m�hV$�)-�˙�N1�p4Ԅqn�X[�(��D�d��ӡ|U��z�q��F�u&_d�Wh�zֺv����:�^/�����E=�8m���x�ݞ]�n����wp<�J��{rE��в��	4bM�i���:�js���-6Y��L��]*ڊ�1f\���nl�|�$��'��w@�t��t	:wH�:@��N�:wt�II��I8'I$���u�;�}�pY:3�l���ې�U��O�WWEn�Ʉ��Ջi3�s����s��I�z�̆
��K��\��B�L����������H��۶�]Op�V�N�=�OF����X�)k"�įM��S��e.�tЙ��R�'g�v	9.dN�ǉx+��6��V펍��<u�95o1\i�s.Z���iz��&��٪��w��[��`��%�d���P�)V��Q+k͂qcXYeHX��(�������<-���թ�0ޭ�MP�)ۋL�Hii�kl����.�t�U2�N�)2z�^��������g�ӑ����Imn�9xB���F��n3㑳�P:���:�H�F4"Q��l���NuE�0#Z�͊j��[�E���7\�M<��z�X=���6���\�$6&h���J� �Wb9W�[�/.� M�u�[�)9���V]I�Q������Ki��w�n���lPHI���@�%퍊����:<��Z��%��c�%�61f�%K=���,��A�\}�[�������� �e��wn��=N��ɴ�;v�R�-�"�X�˲akku�V�e�.�+������8;j�������8P�9w{ &�(:�����������M��xc���H�aH8s�8^&gq����s���v"���5���󟚽w,���<+��'���h�}�W/���&��ѧ�Fp������J�K�60-������/�Q���:<n���/��`g,���>����M4�I��2�73ч�;5'o7>��j���i��Ồ��7p���?w�����fF6A�<������3�xF	!qJ�I�����lwn�W��w�~:M�"���~j�#p�B�)tjȽ�V�M� �p��<�}2�J3H��"�M����jX�y�3���/u��t[�-�E����o��M���Y�(T��%f���G�O�f��a���� ��w��+m�a<m&�z��M-X��Q�B2����v=�=ݵCo+\{L�1�7tBƘ۴����=-����G1�=��#�a�;n�Hƴ8�q��GÆ�	
w�B�{u��;�d��#�i�u�`::C�:pALŲQc�Vwy���S�L�H�)�M -��,�p�h���%��CQ�_a��Å��1x����Ë���{�wR�]���[��Vj��ٷ�M*���1[�n�o �st[��͹��F>g��0>4Om7����t�G�'���QZ՚6ݡ�/�&~W-�}od�ܞ�@�����}L¿f�P�Ա]�:!��r2�"q^�V�:�g.����n��,k�(K)�bf��(Zoi\�<hTB����Mw�K��4�Cē�+w��#�N?����y5!�lm� ��n�����`�tU� ���㞇&�0^v7g��
�6�ӧ�渷]������+�x�4��,���>�l��fꁳ[wl�11a������7ww&M��w^�=b�R�r�25�d6�D >�y�H�D��L��h�f�{�;�u�p�"����9�{mK�d:��ı�3^�V$�Z�&r����&`��K|5��y���ޚ�C��oq:N!9���ޯL���H���${�x���w�T;;���٬n��p�;��b�ҿ-w�K�FF�}dK(�`r@l��@�$<�ޏh)�%�ja2�"U�׷�J>�&�"�%�m�0X+���d��/E,;�l��{`�:���|���fd�a���duv��S��5�W�zD=���wvY ������ՙsj�6�hW�bovӫ��H��($��e�m��9���o�\�{���y���I����틍��%�;;�qܬ���	m�3U�!��Ied����1����2��x�).^H�k+�ss+�vq	y\�sE��T.�؋��A��6죶�����Up�d6�����,+*������wuy��"N�Ƽ��[�?{��6=:Y<Ov�"�����7>$u҈MI D4r�q2ٯ\�u�.���x�G����S�[�Zy_)���.��9� ���݃������[�ٯ�2��B�8�svT��I�v��߹n�F�G�+�~�FkX:��Ff�U?[f[~�!�+�����8/$զ�dX�e8�6Nj�N�Vƭ�̸�x����� 5,�k�q�upG�O�mp�����\�G-[v.�X�po����ݯ�̏t곘��,^�rA�#��38��Y��m�����k�j� �k���-�WF��)kCuϤڼ|o����T�q�o�
	2>��~�`�����mn=N�6(Vf���*9���zM��>��k��Xy�1^�w���P��R��,=�Wj�o`�U����b�k姶Ɗ�lN�k
��8k\xG��\\<_��~1�-ֳ�Ύi�u��a�Ô���	z�� ���i�nغ���(�x�[��j��N�96�r��=������1�����jY.��[-VF�]�g�l�αY����U�Wn;4�H�w=�.��[��3�j�Ft�瓧���L�F�M �ު�F[�bY�l�GsnѨ@J#�;�.)���nPڞ�3rt��QN�ul�^}-�ӹ��nk���w�|��.�M�%�=��[��v3�5�SmzԳi�^ot���]��D[\"dow�j�C��ǄYX����z�fD�HNim!��x��1�̹�;<���������w}������2A�Ibܽ�<�'��Z�^<�� }�t�m�a�#R8	i��Pc��=�e��٦)#�5��1�Sc~˥��]�u^=�xK(GO���wެc�.@�cw��j/ɡ�ƣ&9�v��8vI��:�4��3��p�ĥzԩ��z�_e�2{�i�?���׃�I^_�������n��v���ͤvf�����*i5������� w3׼���O��9��h=3�զqi��'s��8�z��M�}�آ���U!��y��sgy��m��F���帝�06d'=�PP��hv�V;y���.�Nz�;fh�ո�Ú�5q�������F݅��;W��o��r���Oσ�$�W��l�sO�M6�:��3;�eg�I�9��~"B�1��]�x+,��[�4�����:��4�Jb��Cn�?]ڋ0a#CN�^�ߎo�
)yJ�м#X�����,
�KtvA�v�/	�y����+�ǌ$.�D5n����'��~�u
P��͚�;�����s�Ӧ�+�|��1�X���,5IҠ�bU�YTQ���Ȭ�ȶ_�i;�vM��A�̾�F-�	��ԍF�uN�s4�[�w��ލֹQ�A`���	a��Q��ț���v[�ao�����}�����A����,���
�'
��X��y_g��A	k�Ppa�;LF�m��rL)��D�Q�b�(d90yQ7/V�*�_ D{=���T�-%��}}'=|�~J����{�Q�b��
a�|[ 
=K4&5����u��͞ y��F���#�5/RR1#Q�rFj�wn��20���;�,;��Ì^�&d�
c,U~�)B<�螇s�z&a�[�U��E	����x%�[��{��켰Q~�lUA��ׂ@IX�2�^�y��p�]����Um�٣ݕ�z`���<c��=��Pj�t�T�E��NCY���l�Bf�w�p�8��_X��b
S�f�OfF�d�0������R���n�h�W�z�3�\�6Ayx*�Þ��we��3�^�٦�Zi�Xp��n����I��bY^)�|��>��%8�)ɣH��7̖Zz"R�z����9b>;^����|y��K���>�otH{}�kw+ʠI/�V���R
��Ȅ�[�^,>"^����ѤdP�VV�2����˹�"7�
�V�W��n�Ց\����֜z6��b]�:9�rΝ�G��!*6�%,�źl)��-j�l\ږ@���r8G�c�ۍ���*F�1��\��Pe���v� �����W�X�X��E!�=D��:���i#b̚�ɅQ�7��V�PhZ($ȡ
)DD� �s���A�&�i����46+&b�Ѽp����]���ogb#M��ax�g�v3��!f�z,��nI&Ad�I�Z�o�x����cE��}tj�v^q���N�%:�Ox%���RƩ.�p���h#_D�@��A$��I �����s�7d�}�άB(�N��T���4���hZ���ݭYkw�J��d��"L��$����xrk��z0v_}��\���p8;��a��w�hGEdf�#F��4K��������	~�_���-!2t�e�!����[���$JK^�>������4m{כ�
��&/�A8s��N�L�x�FK�S��\�N�0�(}����������,ŋ�ԪC�a���aZ2�Z%�Vz.m�d�p���9vש���Ӫ�Ϭ=���+��^�Ȭ�6�N��a&��7gqya��Z��5Z��f�D��]����.k�}�����B@	&;ßi�[�A�<��ǭr��*"�*O\�bg�wQ��(��>�F�C�w&�H�;r�`��^Y���Q��I"��X�]0�ޝ<���s�+��G��_;��88�D|;ۮ��9���i����1f]w�WL5ny��8��&�RExB!O<!�{���՞��da��5�N*�a����i���=�Äi���%�x\q�Bw��Ѭ<%�*w�Ю�!AIQ��)� ��!�*�n�������Pؗ���R�y�.���tQ:��F�5y*���_��Ħ̒���e��D�
B�XU���9o�h5�]f��W�2�!�`��y������!'zx�Y<|��4N>��E��,�xf�m8�a޳܋}��?x?��I}��EuM��s�]��nW��Un�E��+�s*1�R��w�����`�,7b�c�Nx9��j*\8{��]�T�j��!z��ixf����tNX��p�q�5��U�X;a3[�_;���f�� }/]՛�����/O�6�i�p�l�B�D&ۮz-�֊ζ8�#d+�ɥ�4�Fm�v�S���s0�N����*�M�=%���<���;QY�x�tW������nwiy�|j�����p$�m�$h� ���o#�O|�g-T"gB�ݎ��g3
�!!�'Y��m��a3T[��S�{ŏ���e���?zz)K/�ʅ�Y�W]��a��[�����k�y��G�L[��N�%A���s�龜>�F�|����˞į�����әz����2F#�0ۋG	!��xA���J��~z�O�y	z7����֌�����>��jX� �#t�[W�h8�H�ԍ�̒s(�]`���o��Q�����h(����4��>�s65I`�����z��st"�d��w�$��\����J!N0�I���i>}�WSn\@Nv\w�_��y�sK�FU!�`�i�L	�����=��\8�;��Ŝ�{\P�U�L�E�[�mfe&,udcd�u�����]��ٺպ�h��Cy%����ׂ�8���l��Fts7�u��h;�m�S�>x��L���f��d�q���ƅ�ێ�^ls����!q�ID�b`�U��1U�quc.Q57u�R�^�tl�LR1<o���Nuh�h9{۹|��0=f�r�g�٨�$�v���F�^>�mWٻ=�b�΅w@��jy$��9ۋs��]{����u��ʺ�GR�遦�ٞ$]ZR����`1ʒD�I)�05N�mt�9;��k��j�p���R=Bw|���0�d��~��Y�R����� �-cD#W��c���nJ)@�����Zx�iZ����6�������Ǳ	���o��g���Ȕ�$~Hs�������q�I��`����M/�s$[1aT;��U{.�!�W���n�;�
���k�+W��, �{ٛ�����z�����O�ku��~e��y��IlM+��l�&u��ɋ�����pJ�ˢ�m��ɘ�q]kq(k�'��)O�&�b�j!i�C�7=�R>D]�)Ьu���YF�݂Ɵj��A����׃A��}y��,�
�$�M����|�Ѻ}�I��7�tǍ�/�xK=�y�|��TT�{�,��b������#�1��>�3���>�Y9����1D$�d�l�M�&��S�*- �G;���)hd���gF=s���{Cr��c|ǔ��ɛ��s�����g	��M`�>�y��̀h��y�~��;�6h{�����Qb^%D׃t�7!�R��XwX�t�Nv���yW���&!ꁺ�F�{�6>�p�g�v��6;>3�h�_]�p��pz�v6�a�����=3A�`�H�	2�ə�T�Z�5h�,Ts$n���zy�;���\L�p���x�]���˳�i��<��DT׽�k��"�f�2Y�Vj4�^9�$0��^�����5��{���7ɥ≻�lΰ3[�9vT
�~�$�՗���6�w�p�xu�CwQo˷ϱ�D;F���=���H�se0�Wj�Ë�����p�x�d�ZR�E]�f����2������⩱u�E[��[���2h��yXb�O_aŅ���9��|�\�7����{�r-��)��h�en�5�`LxѦp[z�l'5���Z�o$�⺪�c�+�1�v���Z}�7�f��|q���8w�`R�s��=�$�wû��'t���N�b-	q�M�2�t\�@Z����}�S��}��]Z-އ}u	�����8nu���*q����<1�/���na��oi�����~^����1on����݅�9��Q�˕h߮�/��#d��Dl�w	�h~�!�j�p�=�����aޛs��ⲭV"�kj"��Pu�w?n�vFB��FNc�c���NU�d:��X�*b�wmf��e�(����n�6��2#�Lo\�"�����]>���z5ux{��F��s;��/�׶�⋴,j�~�w&�]�v(�) Ji!Qi�������Ճ���[��sw(^�(t�0٦GM�d$�l���U�R��[w���]��nƳ#;���mX�	�D1��Rm ���kB��!��1�G"'�VW}ߏySߦ�_%���f|�B-3�_1O��&�+a�%
�LW�����T�CA�BZ�s;�J�#4�Ж�v��[Sh�]�im�mҕ�-uP:-1���Q�E]�G���R;�����Ǘ�O5���9d�r��I�*���jǠ6H��(N&�4���7�����q��H�R�m�Ԛ#�O���y����"�;�zp�;�;4:�i���u89��g;���3 �_h)m��D��M��8B�(V�V�Ϫ��	�	��h�ih��ݪ�2d���zy-�
l���0}��C'4ȻS�$-���q	P���6^;f��{j��)�R��X͵�&�ͷ���Z$�ub\���͌ Y�T�'�Y��9p�MoU�MO��i�zZ!�c=on��̛�H�c���4m��%���k��d"#�/3�л�M|o��#�n<{��qi�����٦�T��vٹ;ş�$�(͗�O�n|���l'`�7��=cW3��űS�H�����q-mSǩ�I���	#7 �t���i���Ub���l��#��v���y!��Z��l���%��a��WiH[��};�Ĕ䧑�`U`� AC�m��^J���^31nݽ]��^z��=���n|�X�&�/��՛��,�Zt$p�d,��-����!��0[����޴���~z+�*�.U�k��v&�I�e{�T��3�ӣ\���� xm�A,ל�y4n���c��"B�i�y��U	���t�݌i�Ll�=/9O�f<%��H�v�O����0�43��Z� uc��N���q�t$�F�h�`�ҧ�gx]�x�w�,��Y��YJ!���@��C�U���|����h�P����O<wpV�Şk;R0���1�����F�@{T�R����fd�����w�io2�9p��]��T ��,�z�FgŃ�&���*����ܗ����޶����17�ta�*�lOY=�킹���;��.��U5���xk����w�pxkZ���@N�۰�]�����Q�Ή��j�����h��A��/k�B��nWm{ctN�����g��[��0^s�S��2�5�R���͂Q%�W�˽��bW�j�F.I�6mpsN�xw��<&x����ą.]B��[�/N5ϫ�ؽ������֮����y���n�7F��qty�pN����rE����ێysm��=�����ױ[Tn�q�JF݊��w;��wKr��K�^���Ϛ��
�vn�hq�!� �JHN��>�y�1{�z���J���zEc�\]�W���&$����\+��P�9�/2*d[\ft!�Y#̗-8�p���29�/2�u�b�8'Wv�|36��!����7>�H0�|c/���p&o�ґ���\繆�W����&�N%��6����j��a6��,LR{��z��#��x�f8zA��T+�|͚�i���1
����${����ة���c��Y(&�:�k+9�9���PR����3�c���V��`-l�hF����{q�a�`#��aL{Sٛ�|��y���<�~ʟ@t�0�ZƦG�>$�����n�E*�h��ؓ��p�غ�uOm�Ƥss��N�s�LI�e���1A�v+ �=5�G�d��:��[*�D��$�a����v�u��Wq��>����8�!t;�N�C�\Q�h23p���Κ�i�<�pet��
�S3�ـ�@�ᾇ|�xָ�f�.���4���
]}f9)�aL*a&��� R�m�r��	�[7YC*�e[�B�7[e�P�H�]���h���깍�8'ӧ�u��G!��d����^������=���-���
�:��pY�aB!}簞ß?+��ݖ��5�j��{)�����IF�[����!����'L�1��ANHFk�*��L0�w3�4�,�H�g�D������{ez��>�z:�J'��y��W�.�������盋��4�(�E�B�.��k��3yӚs��&w}zG�VWb`#f����V��a�R|��E��>�ѓV�)���U9�K5��e��~�A�D���"�t�c7�e����9�X7�>0D<k<��~�*�����q��?����/����&�
�)z+qH�^k;��@D�M|�ŧd��I�^c�g�j�6yeø����]+MvWj�1no}>����]�����N k�)�y�G��9@o&��X'^^鱮��X>�V�y���9�}J�d@<2���D���ӇP�`8f r�����e�M����S�y&c� ,L�|C���i:843��6�5\��0�V<�ۣޣ��x�:!��j|H�Q&X��#;�.7�FP�ɰʫ^m�����������䲽51��8\��/�D�2.7~ �����?c9�{���֛���H5���PG\Wc�0�.�9C��	�frd湚��wW{wP���,w�l�#1(.C�֩�QX�,��<	�R�/D�mu���l|}w�ˠ��@���!W���T|����H���rp�#s�kF]�$$J�6�mH��w:v��ft�`ɷ~�Ø�om"����ovxJ�7��An�PW��B���MR����ϔ�t�J��r%��I�ѩu-s�իPLYk�7pk�Y읞�zΕ�áe�����0�3��|�a��s���!�pECO3��{�)s�&�y.�)�^�tE����c�!�T6@)҂�M��JzM�gV�K�w[�x���e�1��(����{��J�n���4(F�x�Q;3�!����l	�H&��Q����x4���I��T�+8�e��u�Ί<�B�y�G���"���0o:��y�|�+ƙ���w�Cti3�P�q��m�/2���.���s;�O_$�rЄt��������B+^�;�����LXt�j�~Ǚ�!�n���)�%��O��^{<}i��"C�s<�,oe�� ��/0Z,�3��sGM�Z��o�#v��w�3��%����<q]�뱦��L8eY��/I	m"�,6ݼ��RR$��� 
J��w��� �~����uk��辙v��%�T8)�ӳS�О�=,����~#$�%��i\ئ��q�'���ϡn-���<۟m����Ҳ�w\�n��Nꕴm����~��>��p^�q���UӾ��X�"i�N���o��K|p`c�,�gy���]���Dvи�2$��\qX�L׌�)Lx��є,K�))P�ɾ1A���٥���x��~^Wk�v��
�_��o��3��D<��FJE�D�8�q<Z%�X�&�u��0G�
�z�'7-�~T�HG 2�uG��(��V��ߺ�	�Bu�2ev�M�$�$H��G]��9vі�����C����Fs�fA��>F�$-��f�n����D#����t�4����)/;(G-EMĴ���C�_pX�\4�{�S��n�xtn���Q|�v��PV#�����͕M.�9Qf����#*Έ,�`p�������I�=��VE�w���"m[�Ŧ����9l��N����2T}5���-�Ż�׻���
4YH&�L'����ҷ�*ճ��xmN׎���]�Y��n�w<�g,�v�m��o�J��D'\���$���3�"��!ZK�m����'oh�,�dN	v�W���Ip�8�MtF�f����H)-����Q�:���N�-Љ�3�Irx�[�t�i���zJn3x�0Q&r��&�&m҅��M��]��v��X�p89�R��lu���r�i颖l�6'��ݐL�cr�N3o�ӿ��)ߟj��>o�Z�4!{��^xe��,��I�����=Dp��vf`;*#���#2��LF�2G�4����u�ϭ�T�n�!�E���N�`���V ��$V���oc��ϊ�Y�ɽ�|5�)��`�|���:z-@�0��$ټVa�#�c7�����^D�VD����P^����c��MjZOd�X����V�g����.�
�\c�0�m D��in�I���n��▏MfU��^���hAD�G-|�y`�`B4���w�Id7R���]�
(���J�-cn�x�E�d{XY�N$H�q!�]�c��8��+*�b�������|�}4��%Y�`��j��w�O��C��)H˗Y�]�-��'���t5����bv:�a�suHqK.5���c'�z:�p��.=��<�5i���Y���'a���IR���2e�M��>0�Rn��$�X����#i�R ��E���.��<�x�ɋ���}Ĩ:F]W��}^(u�
$����4�q���޲�^|阁��6`���dJ��S-�^8�J�ް�T�-+|f
(��{���>��@m�eu����k7~ɞm��]A�
�/�����	�-: �)�_�n׻S	�~CF�PQ���"�������*��n;�z���T�]���ȡ��YHp��Oy��)�Y�j])�	��b�w� �5=w�������"�"7�q��F��_�ʜ}���*r*�>"�f.���$�`�RM�����˼���d�.-w0�3�O�Fχ��5����U��株��Wg��5^b']�ޝ˜����Q��)S��FY�e�IPvKLj骱-йݸֈ�co%�4�1.ڬ�nX��v|���H�e9���SM ���M�1��^�Ɋi�{�YQ���ƘH{mʰ�LTv߷CT*E�E4�i��n9|�����ɝ���6�9w1фOb��Z�
&��������sEhB���;د�U���}��`�4i���ӏ�� p��4L���4�
���>͸���{�?[�C�p�Ch���$�?8��S'3����n��N}!����F喭�LhK�\���aP.�l�6�������!���m�v�p.�9'q��`�;�|4J�)/i�dFS�U���_�t�g(a��j��J�����ЦßonzI;ܝ�`�� b�u�^WX�$������"`ybeq���NBI	� ���@/�������B%�r�ڰ<��۔����kP�� !ञ��z�=��7���u�2�_�Iz����A�Mi+[.���Y/V�����S�˭�]onh
�	�b5���&�=�]��C��YR�h�y�{�Q��ފa��9��.Z�CAhn�o^<��C�O����?�k����e��C�ޤD��G��w^��{�PTg���v�����4��L�)X��咀�(]�8l�G����{�Vn ��vf�K@ F��[���L�CިJ��K3�U��#f��ؒŇ6M�j��r2n�j�bXB?6u�h6 �� A����'��8��4��]���+x���{���ɴ`��m_C�w��:�8���qTZ��쫲�ŋ��ي�88
��h��k���qVW�斶�<���w�δ6Z�sv�5z�q&_M^�$=��vs~�@s�y�靏q[��ߝ�f۫�M�������(���鞰P��<)�cWS��r��� �D��M�f���/�+�>{����Kc���g6u�b�ےEc�Ƣb�fKyU6B��l�r*�Wsi�fn�ݡ�E�F��}~�0�3�}���LAa-~�靌É��Cwϳr��D{��,xC+�Aw�Ø�C�f~Ѓ?J��.��"~))7v�+�콞���$�C�xO�v��E�MhW�-q�l��1V�2=�ܮ��B}2z�C�L[nnj:��'I,�|�S�;o��Ԅ�EK��kc�.�Sp��>���}�/�<�����)�;-�>t��,��8r)i�ȩ�0&=��I��0���������@�f� �a����4T�[�b�J�D�K݉5���D����:e��
*Hq�8C�s���aBRj5V �켋<B��߇_������z0����D|�kr���cW��(+>�4�_��N���HR��P�B������[�z�a&�j��E7�b�rX^��Ӯ<��@�}�l��ON��������^^�r�-�z�tY�lz����ƽ/M,&<6��X�4 ?��2"e��!u7NA��G��6h=���<�zx�9�ƚ�Ϟ��ݾ�x.ݬ������0���Ǔ��|������A���zk.�=� 3����9Y�b�L,��lE��§:\��	�d��%�,����/u�wE�Ӄ>ccj���su?��k�x��S���A�=jźC�o�<{�;��vOcy��}��p
o�B�'N-��|;]�⬠<�Dɣ���o��yS�h�c��{�_�O��K���'�Z�]�T���ɓ4�/����:s��E�{tLs���~=v�n鹫�,���<v9<�3.�{��q����|���y+�'��g!�#�����K��u��Y&��p��79j��m*mo\3W��F�Yܼ����E�n�ݞ�r`�[$]⃜+�e�0��`���.�{����[�ѧ۬�&�}�����T12la긎��>@�nDpV������<Y��n���A��D�x��xf�@j��t�ny�Ѳ�V�f�z���I�/I(�?Sժ?���?��/�B~�I�K}��r�F?3ǻ�/�k�j��W{yJ������ 1��0��g�o��2������F0����I>}2xX�ᙡ��x,�hac�-ᖻpk�=�һ��#��F�����jq�4�c'��8qu�2o�`,�0�o��|�ی)ݙ��4��ڈ���<�C�9N��C��ܲ���s��p�s�6bz�d��ɳK�K�0��n�4欦��Zǭt쓭��D���i��NPۗ��rf�p�o8S����g���\�u���j5pk@��Ub\��-�q�i��r�Sk��s׻G����Z�9.�uӫ	[��f�'mM
��I6{s����۶�$�]��KY0���-�l˵���ݒ���=x�:��,�̜^R��n�Lu�8�`���m/]]�u��bx[���[�Xz:��ge��㩎wG��Z�N��]."][J�B�2�\�emӵ����+��k:v_nU�y�μ���mڇ���]��`�v�̽����z�m��)���3�S͹W�c����/�|��5�c�4� 8))	{dP�Pkzc&r77<q׌U���m$iӓ��vDiA��ƀB]��u�c�=���Y����q�0��9�V݌��ֽ�w+�n[7O��p�]��6�{�1��wni���Ͱ�m6��Uɲ�� �kF7C69���Q�/]<�Ờqlb���,�j���+R;Wnocrp�P�8hy֚�hin�u�t�B���a��|���^I�l�m�nm���7f7�4���qdMۋ'f����wn:��ĸ&L8{]yi�ɋ6��c�.���O	H�tK�HV��B�x����r��u���V˖*"3W;Z�q�׋���G�[O\Wч;]b.N��6I�J<\�֭0���6�y(�[
n���y�[!h)1�0��H��PF6����ʹ����	�� ���+oF�s���p�r�쫛d5mD6���5G1r��0V�p��qȍ=�#����t&�<��e71`�e��[[��ޛX��J��[kf�D���P�"a� ;D��4&�z�������zܠ�i�h�7��Tb�R���A�?���@��)Ҡ��t9ҫ��]Q����&�U6���Rdی�K�PLZ%e7%r�$�-�m�N�Ma�Cm��XYe�Rl�*k��g��#��j˃���c�'�����z�	#){�v���+l� 9���*����-��M[�x�28b�i�棕�]��%������WB�)�.�qr)mʏGF��Nz�᮱�����<����&�Ll�Q�v�!W'b����=��>eݺ�&��)���t\���QшS5�Rq���q)�Zqy�(j��3��!]J|��=o\�*�Y������RB��%?rc%���6�K�a�,�J��S(ЦAI7��}�J7rFq�r�OB 7,mbپ����C��mG��*pX���U��#=.��Z�����#���SmB�[3;g���,w	o�z	��YAp�t�ĈMf_��Ss�k[�V�nX�b��s���~�ꑦ$|�r����$D(���ffw��]p�7%�W�~��n��y�8b&A�M����M[�錙~�O�w�Y�"�O�t������A	���R��ĝuF��v���j�Q�/1����Օ�BR�7d�=Ym�iW�ֽ���*�N8)x2�z��5dHb,S%�.��5�RW�j�x��iuk�V�j:�]�����+��;a+�>�߮11��J�}k��Q�F���q��'�lѣ%c�T��?^f�_v�
R��\Q7=~�؁�؍Ge�^7� ��6>���Sλ�G���g.���f�W�f��.n��s�%��Q�]�L>(Y���V�����G�n��vw���X-
'oV�@�����c�FD���z�[�����N�[�q�0ވf�OK�)l<����(t6CÍ�������U�e�4�AjGW	豞�
Y����zy�6���-C���̍q!=rD��D�n�r-�׻�-ط}��7� �Vcd���G:��y(�r�!b2]�E�OE^��y��ҫWO�k�Z�р��rg����s�����[5�*cG���n�5=�������J��fx��,ыY�+z���+9F�*J�w�������a"��Mu���v�F;F5�$˯�mj�dC���=���A��n�0,QT�2�_�)@�4w�xʨ< c�6(��ǝ���4�9�;���Oei^9�W��b_�7P|�4!J��e��a�	�vx����wB���s�^�Z8��b��88_4>�dC'K絞����O��!p{�m+|�c=ӥ���Q�{}�i�Q��=[�7�_����������b�����jl�%]�Sa'n����d �~}��x�^�6�1m���ռG�����h��˒��^�;��y�m�M^�к)�`�4�q�>a���S��Ǉ��,Z�i�B�:)���|s�;kS�����ɧ_������9����$���O��ߓ;��5�3��+��E�0İ�fH�*"�EH�r�x5�o1����(Y<_�!\S�V�s���s���K4ӂ7���]g]*�]�p���^11���]5���ͳ�kq<2k�(9��g���R]A�3��+!4r�R��J�.u�D����#���m1�5�_pf"N�^�ɡ]�jB&��
���ф}���q���֒K��bDx���<,?7������k��>�IS��|�;a*߄}�
�g�ז�cV��W��k���<۟W2��Ϯh��$ˢ����k���*��9Ҹ���Kt�Ó�9��-�.e:�{.���
t��]x6�TA�9/�K�m�󠛤E���sެ��W��s��4r��B;�ظp����^���3Wdě��=�g��v�c���.e\k��|ez1����w��6�W]e��^�I���p�}�cί;��2!�u�0�����{�u����w*D������F Q�����U>��KiT��n_��B��F��kЯģ�����W"��W#@�m����GZ���0����bs�s��W{�Mywn А��y.�7b��h��7��Q��׆[�)�1ٜ'��~Qc^����8�^�b$un�X�F�LW�kBy�!���E�,� ����?5N4�WZ��i���&�^̤*�6�b&Λ
��|NZ���s;ՙ�*�c'�j?�M������Bt@$��W1�H��cZ���R�W�_�9Jć��Z1}�X�1��ۨ0����k^�o�32��<Z�6�D��Ӥ[!* ������sEh3W�*��㣦��G/ �@S��\M�p4x���D��l>C��6;�*a"��`�N������h�9R�k����N��f;+3�����^�hčz= F��)/��u��ȧv'�:. ēw2��u�@Ji��.�q����nvC���;�Έ �9��� 9)�|�+�{�=�U��X�0�$�wP�e���4X���YѺ�.��"�.�ܗ&=��^�ft�#\�u�J�m�fjl��aًї*��^�l�����s�E2Ä�X8�I^{u&!�;h�c��\�tu�T6�S:���L#7aW�>T)\�v�lL��lmҗ��m��g�x�:M�F�n��af���l�,�M �WtQ�N��"m� ��P���F!̂z��k#Շ=r��	X�A)��<��mZ�X<b����>U�����M�.mʋ������D�VQ�
�=2<�i�L�Gj{��T����Y;{�:m��/ejqw����ڙm�����XA��!�) �+�,I������5$�~Ռ�������u�{�����+p�Xihw�l޵yE��,�&��&f扱���)�`��l�g�S���bwR�mV���RX8���C��>T��/5%c��1������u��Xf��-&g��:��A�-�ׅM���Jl���%n�^�9�rҪC�_U��e7��5~��b�,�w�:���674שSmBDN(���|��󱏙kp��G˖�8e<���L���i�d��e�R�� ��M�e�[4���
�6=�!���h�����hӇ=`���.�)=Җx2=�]¯n"�1v�Rڟ���2��y7Ew��r�GX'ښ�xQ�]�!������J]����fV�*EM�}�̰��[6��VХE a��U�E��u�_W�xz��/BO�����R��Q�ux�݇t�c���m_��s��	�]`��'�e���xe��M'co���Ǆ?N��o>�p�����Z��}����"Ҡ�X�E����M���l/a��XA
���L4)4�O�Z`��H/"�c��L�Q;�m��s1	�4��L���g]�fK�_�τ�E�^�r�N�H$�`*t5���;2I�:֛ŏ��TY�M��jc�VAaiCo��}�?�1��oZ��>,S����a~��5{�)^���g�i�)����}r:��n�xgv��|�4�W���n�m^[�ܩ��.����P]�H�d�]�;1�󂇳�o��-�)�L*Hf�GY6f!��=�C���rF�X霹���i\����	�04ZRp���'��av�z����b��}�PY��i������HK�v�����D�6�Ǯ��4�*B�26��	�A�Q%6Ýa��C3���+֮*(h��X�
�T�aS�ל�������ހ�$`��0j~U~�#gI�dȑNH$�]x^���9=Vz�?]7b��S�Ԉ�"���ܭ��zV��QX�8��^�zw;J�د�����`n뼯D�{�E��:/m��p��F�s</9��M�/c�t��Ox�O>��ro˘[=�N�.�.&�m��"|�BAK�����;�z�9���+ Q_|�j�a��V��s	�P�ţ�p��[վ�؆Y����Z��4M�
�`H�4׫=� w��N��Y��x�y��6.��Ia-��_[����I��3��QS5���{}u����LR|�z/<55"���I�M�6:�'�n�]gr�.��E���e�#��l9����)"�D6̤����NWd��v��z��� 4�g���[���v'�mC��ŕ�y��8�W��)*���J�)�:ᘽ�=q[�Ȕa�T���j��=�e�)���W�#~�Ϭ�f;ۨ%N,	�zX��"5�/ff�.U�p��6K�OBj	�6����	m+Wi˻���>�<~�߷����Xny}O�JɯWw��^�\:Y����1)t?l�lN#$�H# �/:zmB���g�Y�����q�K(SEu��R�����h�P��[u��>ܜ�S�Y�<�^S�3t5z3�&��������������+�����C*1vR�"8��-P�y�U���{.��Z��Mߒ�1x$�,��4T��29 �e�|1���Ճk�|+3�#�J������
��my�o:�U��Lݮ���b���������[Ysu/R4G�e$�٦����ֶ���WJ'��%k��س�J[��H��a�̷~~��<��0ż���M?0��[9���_)���Vx����״���O�Z��ۇ{��-���"[�H4�E�Y�s�O
��Ǧ���PH��ٽO  �U���֮����Z{۲�=FZƅ졵�s,NWfxճ/��@� �0)
I�F�J>��w����޵��k��1��+Ac��CNŝ+ ���K-�ϭ�ޜ8��\�%2�IP�d5qs1��y��n��ߋ~wW
Q�ŭ�0�"R�l��.��ε�w�D����0�d_c�>9��´y�j2\`�3.�ϟ�Y`o�?�����y9��I.�%N�ȡ����1gZ+��oyK��>�����c��^�(ӯ˰3�йي�uyvK�e�&IM��p�|}�'a�ϱKk���I�5#K��h'�����L�np>�L���U�y��~0H߱��2�f�q�i�7��Z�[YF,��1�
�I��.BW`�tǅ��u�[Z�Մi���p��vɸ�te�5ʤB7��>v��<v�6�qu�A�+��n�^7;B�����7�����v^��uϪ���,5٪Lhk-�k33��^6��n���+�8����5"	ʑ�F�4h%�:�-��َk=��FV��74E&�%�V\:2其y|�y<�X��˹H͢��\mq��͋��E6.FS1�b'2�9�f��L�*�|ecF�?l_�`
�^��=�i�����i�wx`��1�Ƚc.���/<���`��4�e��a�s]0a�_�?�U���=�7�ze��@�% �_�>4�~Ÿ�x_L;�����}�:scu)}}����Z	I)!�!�@�v�YE����Ж�H�ND8T�����k��'|��SRmV����7%F���ו���mRM��6�h�����)�����L����=��zZ�q�Ҿ��Et{R����}+���E�M�^�/ñi ��&�(�	2�u�)������z��a(,���3Ma����\��y|��Y^.���U���0����&] �)��0�1M3um4a��&3kfͭ�׍<�ۮY'��[U��'r�٭;��r��K=$k\z��x=~�~q�	��}}mnSJ�^�+���39~�{x
4-O���_Yl�<���'{7�a�h%��nE��X-x��՛y[�L#�nA�
�V0|v�6HTˉ����[�3qh����*��+4�R�w��Äa��$��{-B&̧6����.�t�'<��'#�[� v����U�H)�� ��E�4�����wE
 �ۦ���y��f�Cޝ�6��;�/�����Q[���Inz��<V��%��$�m��M4�o�^��BL��e�j\��/��) ���;�����M�u�	9�������FoB]�z��>��c(� %�Sl��9W��T�ɋs8<<�̵OE�4e�=�66mn�#V�f�_�Qk}�Ͻ^���F�	�L�X|EϾ��5p���-�ZYe���0ʹ����»o=���';�9G��l��v��T���|o�0Q0-�/�}=K}O�s�Ǖ䚱��|��dW�%2�s����8�:�@�5�K���e����������D˘�5r�Z�R]�u�'s=��e5��jX���Fp�>=#6�K��1���d4�m���S��������6|G���.��uG9e=����*��ʚwd�;a���2輋G�!C}�z�y����%_[�=F<�p�i��1�% d^���q��o��OD���[��� kq�i���a�P
Y����x������u��\.��S��2�9ڍ]8�<�+9޼y���L�^��x��*öY��O΃���|<��(}�~�k��p2�6��e��L���3=%u�+��@̬��O����4��S}8���J�\lj�g���U���P�G3��o"=9���}C8�t����̽,v��g�>�'Q(�>�vf�5�`��R�,�4�V׷3�$�<6F�+[�������x�g��5�?����j���4������ग़&�+�����m?b�71=#nH�k<�X�j�(V#&�±{k���Ijwwo��/�z�y�J>�A�ط���9}��^���s�nXǪ��#���y˸�AV��wo�wzG}o��$�A��׌w ,��Z�m��U�#Ѭ�W�1���xO&x_ �w��fh���=���/U����ލѺ�q��;� Z�Bd��ϳ���ڭ��^���<�����}{���rq�'wapx��ǒ�%d�Ψ^]�1��`z���u�]�&��(�\n�{�h��w�kJ�>Ƙ��{�+�011.Y�"�P�"�ٖ=��?^W|��G'�f�M�ʴ��'jmH6��r4ǺA���rRmKoe�g��餩�N�"�P��n/m�2��}���2)����z�N�h�w�:�� X���;L�+úR��QT���<�'�4�t�S֒�7�kȭ�=�������~���e��=^��,u�[��a({�m�Ƴ�lq��_
�==�D��E4h�2�g�c;����9�j\l@��S	��]��:�R��O�)`��=�z�n7�h8'��y�r,���<>��ϳ�٪�r��c*�l/b����X,�Z�G����B9�	�-u�8��pܼ������[o��\-ٞ�v*
I�X�S� !}�Kgw-�}s����T�A�
�,w������M�_���-&n����Y�q@�{���
��΂�,��ZN5��:�o��m��cz��ړ�'��������|݁��اmN���T��i����۝DI��ɧ�oee)��P�Q=y�*N����yl*��Uˇ���9�^�緫�Qt�a �i�W=ӮU�U߭���q1n4ho�W��m_�>���V��������(��;us���;)ɴ"�z���,,g�Wo{j�ۭY�}�H�P"�t{�V�B�| �k�R��|!�|j����>3	bL��X�&Fc�X���*���y�qS� Īd��GP=L6��I��[�N���/���T��!r��.#մ�X:���c�E#��-����=�Ɲ��}W�WE�Q�Y�֔���Wem&64�4�a���VSF�Bj��v�"�nyˮ�^���������䡾����:[��g��\�OW���;�V�����4�ۿ���%��nY|��N�á#��r�LI#�%�O�L|�̠�k�&��g�`���L̦E�z-����x��S�_�������w�eq�{{�}sh@Z��$��%�=vm�N�l�}�^hSi�#�W�씀1I6��]�vשy:�9�Z�NaB����3���I��Q���{��ޙ���Ϣ�{��>����k ��{���T��������of{�e���.}��/؆�{��;#�
�q�E�$�(��N�mY�)���z��mm-ǤŞ�i�s��ė�K�˕k
J��h�<|�TV�]�r�����pc1�s���{��Uς�31a�İ�,>������Ƃ�)=�a��^�L��_X�>E��'��|���%��8��\6��R�������q+/Yq�^�jU�q�X�B]�2� �um9Ȏ��3�<�����Vۘ��}�ַd3��kX�$J�9��j���V�)���'��m�D��Oj�}�n��U�]m�E���ɋG�E웗���v�d7=`̮Z̚���:��:�'��||Wγ�;��"���ݙ���̆D%J�aR^a[���oE�Y&u'�W�Χ�L��F��]a�3NR`M���_d��x>VF������b���T�6�fg������M�k�[x1�]l�
=fh��⯪
M(&�@ړSe������yk�H��^"-�kX�������ݙs�8�����^���1>�E��K��� �ۮ�ѷL6�[9cM���N��g�B�������^�2�ve>��ڶ[fm��4� "�M��`�����F�����0��e��kG�H�4rU�jk�]�a���yz{೐�KC}��.[�J[�e#>�l�E�l_��Mx�����f��a֪�T��wS�(��Ѫ]jT�{{��5 Z8��G��2}�o�|�l��lYv��,Բ�h�G���.8N@ܮY��rY^B}���=:Ҋ��3-���fF,���9��n����F�39w�*�=�����y5޴hwRÒ��ŷ{.ffq*�s{8�i*hi��-�ͧ�g[i��u.}�X�'p3�J���vt}��X����*�_o�o/uY�rn{%�A=Ċ�R=�����B��/V�����^uޯi.t�э��yv仼�U3�l��a�9��3�x�W�Q�˵!�=����~q�Q��E&p" �&��c��b��V~�i��zj�@e��C�㝉X�vX��k;�y9�n�ֈKi�II4�6o��B;W���zQ���g:��8Q��%��y*������o�Z��5������[���ދ��戁1.&���8�]J���`�W�nKΫ�;x�AY�PWK�Q�<7��bC��u�%��G'��&��={~-��pE|̻.�m6�	iQ��Ʋ�4f�[n˔��J|��[2����X��� &������?�������ѕ
Oth���K�<+�J}d{�������׏J�;ٛ'=v���'K�ST�)�[�l����{�7�f�T�Z,+�����ط��L��?C�Y����t����Ep{�}��T��e�F�
|KSRI����H1\z��E{oX��Н)���K��mة��c�o++�����c�#m8��NY �C��_���z�n��k�|�W ov~��s���Q5:y`H��&/�,�E����hw,��\��X�3��D��(I��g�)�Z_G3�g�f���m�w>w���%�y;b^[�c2)��$oҥ�����=�d0__`�H��0($�i��e�<]��2�l/R��'�tx�gk2L{m�7�U���D��������ɢ2�Ji�UY�ҽ�w�uҊ�{ꉎζ䧡܉�āO�/;���*;5�cG9q9Ԫ%�=����D�y�/���{Ŗ�*��/� �h�t��f�IeL�`W�|�9��r���K�_��6��d��*�*�w�Vc�n>p��ч,�n����ٺ�8�0�3���W���vt�C�b�tz/v��V�o�r<�@�#-�bj@�5oZ��|�y��AV/��U��J¢�h��H�g˭�,���'>
��(���PsA���m��qca������P��ǒg:Ub��u췋�a67Ô���$�
�$)�NK�[k�Ù�P�t#����#϶L���7R��s��e7m��t�mou�v��3�"�{�n�k\:�n�a�V�_��t��/kȨ�;{�%�o�?�l!��*4SE$�U�����pz�v�/�Ί��2�FI$��_/��:]�mSn*���b���m����y>�4e�r�y{�{�L�����^�g&#9(���rjh�fcf�+5�En���iu�ٍ�9��t��I�B)�QA��K�)�t��;���v�x����{�j��C�fi����<6���>Ѹu�1`ٽG�^ǋt~�7Nв�*� E2��u�j�I�rX~��men�=.�c�y�[��
�x��t)��S�V��;70�W^�#y:��p䄐�)	E����=���}�,�((�M��C�����^�����.�ԧK��̹n���"p�L5���dl2�	�M��K���s��a�.�1��Q�ȡ���V����[���Rٻ���lܘa��w.qUzJ��O�H3��j),_ �^r}g4yW���_�8�o8�Uy��j�)#���A/!o��{������)�oɠsi}�>�OlQ<�õi��b5U�?{ީJ{^���"��H���^�i^���1�:V�G�/h5��3@R��~o��W�����gF8�%�Af�5=@Wv��u��n����,���.#���e`��w=��l��;fۻp�ѕ��m�&A���]=`�y�����9u����v~c�]N/WrWWnо�7	ڇ%.�X,�[`�;;1�ʹ�C�$�)�k�t�6�K�hi�0��,%����HX+.���V[V�\M��tn�.�s�SEv��8Y�u���6�x{;��^�MK�Q�������c%�n�����$7B7d��l%"������[��F�����������qi��J������w3�),I�y=v�X����X�⩁A�d�������Yi_�od||k>&��p�f���Ut��[m�Z��J_r���37\4���5l
H�T	������M��q1f'���:�zx}Ky�>�@:+��x�Å��`��o��Wc7@%��0}Pf��b�A�(��X�Y���K���a.k|TM�����o�Z�X2�gg�O���m1~��������eh�H�V�pWP8�%2Ke�������4�u9-�z����i|W%h)�S�FLҕ����Dw�i�evE���)���������x���2���i�%b�U�*�x�v%50�Z��v�cl]�-m���ٟ|�k	9��v܀���\�����>C�/�~�~�Lgd�yh^�f��7�X���f�z�o�^�$`�Vant���rI��	�Z:-������]ӽ���-AU���I�[z)�m�`�~u��?]�ǶS�;/����;��7<���Ss6V��immn��KŤ���B�(K��O.Q�ҟ��*�_��٣kf�TC9���jG�l�]��wGA��{��f�6Ӣ�A��`�n�MT� ծ�ҳ����?>Â�*補�k�u�.�ڙM��w<^�o�6Y�������R$Bf��pw�Lݽ�;v����kܬ������'m
>O.�nM{=nn��yѰ��I��ӭg+#��2�wemoi��'@�M�&��X�Iq�Ќ��S1��i紳���I%^��`uo��w�r�/�sT���l٤l�
��o��h���]���:�\�3���mstj��ųMc�j��u,h& &�u�Jm�.�l��������.����k�����x��i�ՙ۽�yv�ٞp��[�
Y�l�H��Rt�d2�MV,u�����dǞ��oF>��*������Wxb��o���+C�[ѝ���6�>�}aԂ��s�������%wcGa��o/�fE�f��Yt=� Gi|;r?f���Q��~��fWj}.��*���;���m��j1���k��k޶�f{��t�s�=������b��Mރ�T�E�{޻���Ud�S{��������>c����,�P�R�K���%�9��w�q�J�˺�n�ݧ��� �$߾])W/u~�.����������S����eI3L�N��l^�ǈZ���3��m����n�'��~�h�}q��F�+y|�*1 w>F��s��ߖNxՁՆ�1i8�02ZLJ�ݳ{5Ql��X;��f�'Z0��B[��!��	��U�׎BL�w;�U�Rww�U�g�T�R�Ǯ�:�l>���63��׳�����ݠx�JtCZ!$�j��>�H�%C�+���ʋ�]H�d� �us��8�X�����҄T��چ�Nޞ�/�zh5�����(��F^��$�5,Za�Fn��t��3�
�z�اl ��n�z�×���{������\�q����죙YG'��n���M�f����t`��S��lT�󢗧\��w|��P�	(�s��O�7��
y�!��G�R��ܸ��@��Ƕ�珮�,�7uk������z�M��Qv6Ti�Y6i[&��|��X}�l8��(8﮺�x"B}��>�sg��k�7n�s��M�rr�i"@8�6i�Tڕ���ڨ�[�$3ieW����΢z���m1RSH�O�����v��CM��^���b���y�{��\| ��-��]��&��(2�-c�+�6x�3.p�ѷ97����(���hdޘ���ֲ�;]G�Pve�9�Z<p��,�0r^K��o��J}m�{�𻸛[}cy�(��H4 E�"��W˅�=�5��0ׇe�gkk'���iָ%0w]�~m/'�#����EE��]�=�2=��1�j����T��g�/5�����o|�V�s1^/$Z��b��u*�
F���#3飲���t�d	j�Y�c�3lX�h��s�
��l����MN��0�y��|*����T�v��Η�d����gNIϳA�Stm��.C���,��j�,��xhS�3;�ߥq�����:�'r���pMhgc�6������':w��j�T���`\S~�α@}��=���ِ��'v�����'��(\9�2�b%a>�H˽����o���9e��f%������3����^>cS�q]��u4yX�ѹ���@W��G������;��&��=����Y����_'�v��!x�V[0�[����1L۬�a��[��j��d�>��1���"��ׯ6���\�������8�׈c9\���6���z��ҏ2W����F�#�O8/2@N�׺&�����jf������g�>�w&����a{_]�9�F�5�T٣���J��d��r���q0�����K^�Fϸz��.�m��r�"<�&���3�i�`4�Q��r;��9쬝�~�:�f�0��3��^�[��QS��㛝a7��~�{�LsGt^��@	^n��ʡ���(�D^�p9�]��f{5I���I��Vjrf@�Ks!���Gk��V,܊������d�1�|UE��ͽ����γb��,C9<5�4��5������ 	L��^ob�d���z�vw��n�����V�<B��.��P�j��x�� ���6��vc6���f��_��}�L��3�پX��	_,}F1������3ԕ�h^}ח�Γ�z����x�r�zxg����_�K�'��WJ��W*�-���2�>�#�%쩾��I���o���X ��L�A�g�i�F�Tr�wc�*�{�=0�Q�3ǫ�K�=������뒯fn1_�Õ�eֶ,ն�ۭn�iY�ݐ�y㭳K ���sܼ��9���3���tt����l*"^@��f���B)�����6��h(�똥���������5B�/ZM�n�1���+�]��qp>rZ��&*�"{M�eJa̷D����	H�uSvvRլ˚�e���Gn�޷;�,W#�#6��P�wV��ΪQ���	��4Q��y0���kd�s��0�b�ޫ�6f��OXf�.Ź�2tҐ�q7]��<�.�@b�F�[]F�%�Hu����c������D.�m�ż��$����M�ێ���[�d�X�/=gtg��۵���3.�nfGu�]����)<M��k�V�{Qm(oT���7-]-����)�n�\�U��n��s׎�s��vyw�P��^�z��H�<�GH;�4X8n:�6%1����+�SdLQ[�U�ix�E��4:
=�lq9�ܔ��^�p�oM��� ���n���@�t*�c�쭹��t�"�8k:���ö���ׇsՅ�!�:D��v����p��I��I"�y���gctu�5�q��O�n[ٔ�B�<r;�`ť��\���yru�#&�����.�<�	4�q^�Xa�,�&��ȫ�����W\���H�WS\�21��2�uN�n<���A�m���<=CsN;v��,3n��s�2:�Yi�1,$x&f&�����n1>��ˈL�d�d��sKC����e����\���-���cVP��{�q���WZ͖�ڸX�;��@3�̛k���ˡ�m�-�c&��.��m�4�i'�U��>8���;�n�AJ�i�l[��۫��#��zD�n8���Q�����{*<���K�'gLݻl�\E�Z�<�	A���%;�����m�q�l�B�Aٲ�q���crC���ݺ;B\$;ڶ�Y�ɷ�KP�۴�-�w1�(��=�^z�4��$���`�u�n㌎���<\�2��(秵�ʵ2�Fn�vů��Ha��\��f�SXu�-݈<Æ��]�هe����b۝�u� �T��i�im����wogx� ��Fk;��Ͷ�A��f�E���
�J�r=���y�Uq�!4�c8i�h�t4�5����-� At�҆�in�i�6+R`��XT�JD�X�q0�qs��@(!�occk[�᪌&��d�&���˛l�������7Eٻ:�f�
ۡ�	�W����2�TJ$6���r%�s��11�z���w/�ߒ;9�y	����I��wi/w�m(���P2����A��u��DS���v��2��Nӽ?6�5���Nj�ˍ�NRbF���]�>����.s�a�4�!yJA����y'��R�'��S���W�t�����՗��v��˲�ű*�_���V+�>ם�G$%�h�cm�K�k_o�	�~}��0�����7�a9x���+�e������n�f
�s[�{ޡtY�	h��%�e��ѝ�2ً'a��u�Rh�I.�Ն�(�AץJ;��ɞ���+޶�3��<�x���?:�4)a(�r�,@��ٶ�=�Iլ&��H�-��I֚+�1���َ�]^�W��|�/����y�m��@�<�~�~K�&�&����ם���M2�:���W�v����~T�����%���nH#�-C	Hw��Gs�l��S�/�}.�5�;W�}���/Z��.�+D�]����m��:��/E醽O�e�٣s75�6{�y?M�J �k�w��݋a^5=��
B�H����Z|v�����e*mtj��?(�Bt��xX���N�+:��"��7
�W����^X�+(hJ�|�{{̌̆R�pP�qht�F�B�I�c	@���|�6}�[�<�әiʧ]��<{@�8��bb�v4-���`�e�<����'�i�j�a$�L����O���et���N��7���C����E��6�����ir�o8�t��,�$�	��gE������DJ.]����h�3��l�ɶ��dʭ��X��nب�$M��۝-滚��\�曧���Ç���y�����q>�ʎ�i�V�r��|�����'�����Ѷ5@�o��$��)��/�)���!�����ϫ�'�w�7�4�PS8�jo��B�<�s���zQ	�ݧ��#N�DI���?"�w����,z���x����[�,:�h:��[��%�$���д��l�`��cz�
��xgg)\�1/����~;G��L9p2O�����,,�����b�&W��-��8+G	q	�m��{�*a@ȌԨ�N߼`ٸ��׮6!�R��9v�S>w'X�����s����]�|iq+���@\l`�}+��PI�	��DaG׾U/+���K�T_;��k�����s��J�ǪǏ$�Û�`[i�š���L8�8ځ�<�`�Z�Dze9�Ƒ�ɰ�����%�<[S�8�f�h=G5�;x�h��='7e�����������3��_�/�k���kKG����Y����!�zK\���Sd�@7MSm_�<��)Dy�u+�Y��Ir�@!ɸ<��ycK��o_��y��*ݹ�������#ݮ�XN="��%�  K)�������1Xɽ�u��/�/��=�2>�|�������~���s��_to���G@���(ӦXj{*�����^7���n��TAF�۹S�5Av�ޱ��ǒ�x�);���y���V��Xe�ZC|{�Q-���E�y)�_<�k�`��W9�G]��;|w;6�<���f�J����]׻>*����$�a��)����"����K��/�=����s��8�ΐ�"|7�{JĆ=�c�yØ��^�/W�0}~��~|�����q�r�b�˘�$��!�H���3��7ie^il`�v۔��N�"�i��=i���w����7����xW���7f}���h�7 }R?w ���JC_>a"�5M6�"�N�vSL6Vf��\���fÿQ=�ir�]bk���w��k�˓%��*�k6�|��^�����[r�Q�y*^+5@o�ud���.�DXˏ�7�+��l�A��Ѽ���떗y�]�G�F��H�&Lr]�ؼ`��2�g�ō�蜲�dr�ϡe��Wj*��QS�*R��Kٻ�e�<wЧNCr
n>b/���ެ�Ȣ�u����K]��s�A�{mԓ�-�6`�����o�����e�}_o��rv�>��G¦5\=���8�{b�)<n{�s�N����+N^�c�¾��ܘ|�������G�>�k�x�=�Vfv���x0�E�\i��n1����V-�'��ic��;n[�I�{B�n,��]�n:����2����h]��i6�!��AS���m�<�����q��0<6��Pr���+e{s�+��עK�ak��G�Xr�y]�b̥�N�2�nF�]��e��ë-��c 4˓�
\�ƶ7&M����#��[[�+�ө(�*�كE�˦�vo���y�Z�sE�z7%�[+Su�,����nn�+���0$�akl����k*ׯ���vN|�-f7�vs2��(�T��>�3�V��ԜN�RZ�[f�2��;����]��"����ϲs�S���M��k{�%8ǾŞd�a���x����佟#w�yY裦�z]f� ��*ʑ�a���U�C;=c5k 3�zS}wS~��2@�e�ˇGKQ�^r���ɛx��%!ȵ�-��Ui P�o��8ػ���]uf]׷*>4�Epc]ݯh����=����r���v:�8���؍�R��h��9����U��	5�˦�Cʤ9b.~�d���{�:�cj�/��V��9�s�)��<���Y�>M�M�W������w��n���=�騋sٗ�I��{tf�64����[k�[�����/\�3�t��?��]_g�ڱ�M=�9�6n���4�窙����[�#ia�>��*�M6Bm?mB��|J͙]�n���aT<oa�f�t��Y߮~��^@l/ǒO���x�K��U�C
]��ף�n�Zg���ǘ&I�{r*և�������T��d�7�ז?�ZhW�,��UnM~�ϯ���}ͺ�?U�\��Pa�)6{��N�8��i��#��õ9�|c���F���ϻ�߇O�{��ig��ڗ��s��n!!l�Ĩq��Cecӈ������OVz[ض�������`������D����让�R����R�"�.^� ���M a�{!]9$ߢ�����ϟ��d[�µڟ�Q|N���/���<��ϲ-��Q�U��-j��
6	0�Xi(���i���\��������E�sVcmr[�-3X��X!��CNK�Ewd滾�ѹ��S+�7�<9L�6��6�A���vxc�c�����~<��Џ�/�y���	�q^o#i�?XY�>?�l��L�=�����A[�P�N����Ku�Խ-�v5pu��ם��"��[]��2��1"�[��`�����su�ặ���و^Dk�5���<{<f���멣+�Y��_��s��h�&�x^3��0N\�Kd���I-iq{���k�Mz�C�G�̄�w[�\J�u&( �L�[u��V'g����O�w(�G��C�!� K���.�L��彗���'��g޷�ƺg��O:�a�$�����1���F�'n���΅ �Kk�o��yJ沞-�eM��D�"F��G���4���6�
�[�\���-ֱ���v4L��a-/m]����^�iD ����ZM�ܾ9��j�#y���z�m���@7������!{�ҥe;A�؟�{o������yun%���-$�I0cp_<�@���<ɄR���.2v�����co���W�1�»��Z��IΞ7��Ǳ���}����8E2SE�Q�"{���[���%`{m�?]��xOue�j]B�3�����q�[�]䏽��3�Yd"���aQ������A�mv�-60��Ǯ��rmz�{��o��!_{��<�yMJ|ĢA��湕�^�'��{l��� �%�	�ɜ~s/LF����r�{T���D%�/5f1�r��y�����*�-*��S`�.�<�~��F������zǹ�Z��(���GD:�.��y?n7���ܡ0S��*��m�[n�T@�b�SrA�yS�'��k���Zv�4��unp�������6p�1-��g�,Js��G3�w�����3���ܞ9w��ɝ�E��m�j,g;�gS���EpE��Ie2��,��&ϋ�}�Sq��~A�����j��r|W�u7ܮ�©Q��^���+ٛ�*�6����w����陈jŹ�q$RE��n%�B�+�^I/�y�ݴ��
v��#�=�Y<���D�-��k��mo�*FЂ9!�<�o/����
�c'�Ļ$W眾:=�.}��kAxF�7]v#�,��R!z+�{�.���㤈[들��,!6)Ӡi:����]K���2GFt73�5d�_��~���S쳟�������k�.��BE����z�W�$J�um�Z<O϶�m�����w�:ƭֵ���N������2ʢ�61fC
s�Y}����n�z�4ʶ��D}�};�r�Z�6H�s������5�C����`a�j������
⛩d�ed�I^I�<��nҦ�vHzq�����b���a9۝�ތ3����ۗ�V͸�H�v}��]�w<T]/��ͺ�-X��;1�OUx�£j��;�ɘҒ�&G��.����(�$�7�K���N�fO�W�����h�Ϥ6	�l����F����&6�ܭ���[��:�=�m�<�<���(�C��/����c���0��}u׋��{ :�WT��]�<n��+y[��V&�|���a8�nH�p��{���-�5�W�_�]���q���V;$��^�������ny��0&�{�/�ʋZ�%c���K���]L�� ���3f�$֯��ćtLm�S��̦3�G���b�?w{��i�]�&��R6���GnwآR�b)A���30vL?'�|`7T<�n�o�S��a���vW�ʴ�,��K��
b3GV=��\�Y�4�Vʋ�`R�â�d��j�$�٩x�6�ڤ�L�O����_��rC�
/^�����'zs�1��<0V´�����ٜU�Ƶ�Id$gi��$���8DŲ�۳���d�[���A�����qM��jI��D�w;�w�*(ع��Z�H0��.=��Ju���#��]��R[|���n�y�S��pF�
e��N�W�®'�s3O/}�?a�y�x����ߞ�)G8~�ӟV���E�Υ�����4ґ:ʵ �O�dQÚ\�w�\��h������j�f��W{dZ�՝�>�֮�}�ֻ4깪�M4�yx�b�C�����fSr9�g����ཌ}y
'�r�=�cE��h��a�d�j�����[̞m<]ϸT�p^��x兽�~�.�B�B�m�eJ$Wq-�$D6Z��%�i$�i���ܯn��]]�pK��}헂�����7��ֻ�������K�;}�]�����A��1x��"�q�<D���O���W�a�tvf�s&Mf��ˑ�G.<͙�ʜ�7�t��l�|fV�t}qm�s�����Jc���!�`h�H�k��I*ř���&���ݿ���� (�n6����QH�%ҎG�}�X����4mّ�u__a��%���2�S�J�����'�٤3��z�7i������<IPFZ)F	$��K'l�=�5��{���x�-����&Im�ڵweo�W�>�̬7���$s9[�`�[\ji���}�3V�F���V���G.�Yo����K��m>﷘��~�L��ƬK	Km��u�w���xN��R{OzՆ4�p9�m�5}��C<����觟��$l�x��ᝦX�~��]=�ߒ�գ:�����-�y��~��x���'5[]���\���d!�HG��y!����t�����G;�޾U&�d��o�����[Fcĺ�s�	>݅b�.c��8\��Ɂ�1u۹]rd��.)Ϯ��O|��8X{���d,K�/��1����8d,�c���ջ�8�2���!�,��'1�^��Y���Oh���
<M�WC��O���u�x?hqSp��T[�x?��U��l]o��g����g������3;��T�X
;9��C�Yr���Rz�L�N�dZ){�y���-@��h{��@��]�q/|Zo�`z�x)��w�lӆ'�1J�*�Ts~%Ѹ6�8��`�g�����Ь��L��go�����=s}�^�2b��E�=G�ͻu�5%S�vٙYz�v�נoс��%)�km�}企5nS�@�ܲ?X��~86���j鋽��=���N����l1��k��ѧ�j�xx�[�T�,y��e���� :�w�o��M���[<��b���մp�#? ��gc~Y�[��)���|1�[>�\�.�7�����Pܧ��g�-�8a�7�p������0���_��>���a��@�S�`�Jv���ԱEKwbD\*	}�݁Z�C��zNayI���:ٽJ�̯��P�s<I>ˑ�YzF��|�<��E�F8�̭���� �ŵ�v��wFy'��.�5���I��I:l�H��{�7��?��G=hW�������y@�$E-�˒��wk4���ʸ�BEG��s�5�Ƿ>�잇r�CR,��m��n��9*��r�=�d�ģ���Z�_���ķ���/�Vl;=�^�_�d����NF���j�����6�y0D�+���R踗B1h�\s��J7W똸�+��\�m��Jl��`���'%{~}	����ܹ�m[���GM��Ne�� 3�~tO�0K{��ª�e�T
d 2�"�!&ԓ�?%�T��X�9��{������Tȭ}��u�+k�I��wYC�ud��E�%�`���vW�T��/�
*�dS���I����w��RI�n9���|��ȡ��!���ͩQ��.蠇�����.�Ub�0 -� %H$%�or�/�~��$��nG�E��}&�l�1G-nr�*~�ڙs��Fg|	������ɗl�MS�֭#)��dq�j����SO�sA����¦��<}�h��Gew��Ju2�:`X;d�契/���L��f.��i��.�l]���u���ߔc�2G8#;t�ON���yR�*e_?���51�z��ǖ�	g��G���?~O�l�e�@	��uBh��c
���n4vN[����8��{uZ譮:��8%��i�#���#۴�7��o��K���.r	�����?�db����.�q/�^�����>�u-+�L��^�2E~��t�,���<q�V�mzI���H�*)Z_������p:Oqd�db��v�u�1�΢�s� �Y
�n�<��7:e	[ϲø�I�2bO���==���j��y�e�Q���-���H��tӠ�$L�q�}��_g�za˺\���K���c�����-a�^�*��v�~|���+>�c�Ax�C	����rwl�ffsXW�פt+��=ت�NvOQ5~tY�W]��2G˸���!�y�5��+����yM3w=����s���x]� #�����-��ӕoc�`;������b-y�07�.ķ��-+���^9eٕJ@� ù�p!�b@e�ؚ���6"�m*��h����;Dl���q�Su�)D`4�%yq&��j����L!Zggq!n�A�
u�;�#��T�;!y��B`1d��`*�L��Ȉcu��c8���r�F]Z��c�vz�F<�|=�b]m�6����U�;b�[�:N�u�õ�v[��q�vܡ�5�/8/]��snr����[�^I���Uk���qČ�!�n��Y�vc�����oc���+n[��̋�-E	T�e��b�Y�'�����K6X,gw_�����L�9��a�͏0���)��H���놹c��o��W��h��nH,f�bA���f�gz�O�g�[XW>��	�����u�Z��,�Y�����b]X��3±���F�C2��"��)	Z��2T�G�<9��o�}��q�hy����}�{d]ǽ��ϸZ��-y��f^����LQŭg��u۷�c4_��lc;ur��
��*V��ި��Q,̫� �w������Lm�Ƥ�d�ǜng���mC�H����_����?*�I��k��y��h�������ƍ�|~�=�R��W��>N�]���x��Az��w��K@���F�Fز�, �R�]e4�;4�.3�T��5ԃi�A6Q��!a��^^�c��䎺�� �_��/��:_\R,�h~4��ʞ[-v���-ߧ����%4~&�SM�DՕYW
 �R���j�0�����_O{Ƈ`�7���{�N�n�Og�C��e���֏l3f)}��|}ޗ��}�2\U90Á�{N��"̉���I��1yxO{����<1�x�OYސ6��Ȭ�*$�Z�~����GQ�I��}����eNݗ�i���m��Nr�]պ�[�J��f�h]~�מ���s��J�v��F�	��D:)&�������Gr߮���ŗ��ke�u���ޓ�x:Q�R���ɏ�HSG{}���`�������=D�#p�Si����aˀ�^P����fPu���o|<W���ܹl�5����D
�޾�񋻏$ֵw�-�p�іhXE$]K�Y������Ƴ���b�-�L��n~c��mR�J64"�r��z��y>��3��\�67yL�[�:�K��c{��<����u\�t�#oty�����(o-(�D� ��L�����Vݝ0W^3YF��p�v�r����3�M�^t�[t��(1�͹�`yo�헖j�.�@�"�F������ޯ- o��,�h"�mn�
'���{�E��뭼YsǇ���x��"~�Ҥ8�;$%�\�l�|�'��/��麣H��]�5���d��Nnz=L�W��R�U��.��0:T&�m��v�e+g�7�U��5(��q�AQ\���e�r.{S͇Zʁ"����ܷ��P���b�Q��^���r䕼T�z�
�mg�χ�tĚ��)6۩��)�d9<�^�7|�{�{ SR���n2���#Q�~j`�o�y)]���x��s��
8oߡ�\}�Jy��6�سP��,�s�;�{d���r��lP�h��Ecep�i�sz�z��-�7�=�����R���%u���׺�m�7��b�P���o�5�^��^�x�K�3٨p@�6[4K4��x<��'�{*{Ger���1��ٌH�;;U�?g��N{�#d��;�ە��ו,�*mj��ՏkA�i�鶝t��"����P���Rl�{�c�_���.�׳,^�|���U���=OU��)U
l���B����Z�<�,S�%�n�g%qYTP��O�꒛���g�k6��{}MO�e�����{��#F�����"��V`�<8ltM��l9ý����˽W��.��Ï�kMó�)��H���U���QML�ot���5��_�Z���6�!�t���f�#���I.SN!N�>=�?O;�;g�jy��c[�zՇ^�ύ�6E��K�����=qV��t,��S���L��o�׈�k���Zs�b� ��W�Ֆu��v�'�{����3|&jK�#��AI��b�as�,w���Il��f�8!�h�.��";�-�{"�l��H��]g}_58�+�ƛ�x�l"Zu~-�nL�>�|� ��$�*o��c-���L��;�]�.�%h�7�_	f�#G�2��B�o�pU�h�'���u/P �*0�\�pV>{���Y�$5�u�j�ˎ�܂eJY�����~���Le]o�!��K��ڿyi�m���$���b�K+{wبvL�{�s�]��n���%����ܻ��w���S-q��&vg�8Ubt6�|�R�i2���t���=�+���/��I]��L<���#X����Rn4pf�ұU�u�͹�B�������6G���HS�=�l��}sݝʗ��6[�'%jy����I���6u��K7.b�5릘�Y�X`Hۥ!�X��9cw�IKmM����ܹ�۩�Wc��� �n^\k��f.��ځW�N��g^q��X�Hx�^5�b�F7%rB�#�{j��c���q�5	��zh�h�f���:����k��k#˻g��v,-Wh-s2�\�d��\ƻB�hi�ѠT�q��XQc�i��O�y��4�!�V���iv���MmW�κ���0׬`�ru>���˰9��ܕ���i��Tۢ�Rn�:��U��p��.�\Ӗz��51�~�^�z�'��=���(=�u��q�.���Vm�D��D �>�@N�}f�m}~�0s�(
&r�[[L=�<��^[vׯ޼9���%%�p {��Z�R�	>��rE�s?��gמ�A�|
�<~�8�n�Vo"+ؽ�#��Jx�������lj.h�p��Pr\�r�rV�}Y�ǧ�����N��o&9Q�.v���'2�����|���L���
����^Ǟ��ݾK]^y`]��KH�g1ٮ��2�X��m �(;qB�z���[nHT�N��["ݮ��
_�4�v�GK�XS�7@Y��f��쩰�&q���~y;��1�U���X�gȓ�댶XI��u�F�F���!����&{�����j�\�cr���v�.�wNg4}���_iߢ�+PY�ſ��o���o����'ȋ��Wma�/�)��M����]���f=嵻䞲������u�ף�G�����o��GqI!��HTv���LC�Gw�����e�}��;C����w��|�E$<�_n_U�ю{g�ԓ��(�q��\�}0�x7��	����1.׏��}�'
�l~��gx�=�E�) ����J�2��f{����K*�m4���BXJ�LW�,�{�����(\�q��nM����G1E��ʻ\��em��R��=�'Z{u�[q�(ݭA�Sa7])�i��!�B�\4k�^$õkń�>������&�+կ��?]甀Ɂ_��a�~rH��
��Dښ�"�\6c�(�X�6c�{�nv�^v�7���{�N���)C��[)�:�<��j���sr��oG�t��a3��-�ȸOG�0xg~(���,�خ�Rgx�J>�����MD��A��]���yԮ�e���;v��kr`^�~��,AB�/}�����7[����g�u9j���o7N\L������|cۚ��"��Q'�B�(�I[��H�$5o�MAߪ�ǰfMPN�[�'vv�i��s�_��;[5y�Ϯ��#-���lu}�R�Ȧ
�A)��*�v�2�9���	"Ǝ�2Bt�W��v��N����.Y�{��y^����ޕ�ׯ`��w���o�\�^*۴E������z���۱3��VA��� YP3�/	-M�L��$�wO NM��x<�H�����ܸV��H�	�����p����	�����a��L�ݱ��	m��6�E��!���<���7OQ�|PTe�0�GV��hrw�ex�u�����]����b����	����<�Ƕc��c(oz:e�Y͠�����̬��\h��Nmc@��`tZ �HiBi��B���o^�5�'R���7��W|��^~�ɂ_]L4�nң�Hp��w ��z�����_A0�:���>��g�u~y�_+);����ۑg�FS�&����A&���΀���v	@�E7L��w��J�Xzs�m�p"���HEyQ~Y�-}�Z�S/����|{���mw�㏲�"ASGK
ԫ¬U2�&4�)��Sqz���9wUuŭF`k��[LەX�6��&�D�D����
lZK�G}��I�u�˰�9z��e�Oq~��w�.=�s���~EG��߼?G�f���SI��Jw�.����x�%�������!�|�,��:��O9D�J�;7�6G�OMn!^���&��A��%1�����w[�����eԲNks8]u_:�yZ�|���$*MCf��{�aEy�)�i�ˌ����(Vp��B���e6��6=�7!��Y�,~��ǀ�<s��<�뇽�=޵��u�%iSH�E��i:�<h���u{�2�֭va��c������Zh�PG�_�R�w4x���斚����ڞ�����Ne���72���f�P�	D��ʅ�l�`�?GT�;�0�#h{����t����t%��ˀ���}/��xX��vI��%��Y�f���Ԉ��:���{WnY��_���4��7��^��vj���j���V��xr�:&�!%)o��ㅲg���|�K�6������ZGOE�y�g���V������S�����~���z��P8���?D��f�Yl�ǯu���OƜq�v�e��.-8���0o�I��1*:��R���=�j�����C=+sA,XZ/.-~�@ˬL�N���=[ڜ�,?h�p����	�K�=q������oSs��_�i;g��Ӂ�.[qlZ�� /y��T�}���캽�^[��v�������3�tR連@�Hn<�9�ػ���D�5�\��}�̹�>�1���ǎ	�\80�^��g����v�~`駫�r���ԣ��o��^��o���;��	9�Z�u2m��5D.{=�;pg�7��پ��`��O�c��Ԍ�LR�I�u/f����~�Z^�o@��;�4sT��]�|��)L����o�����+}�P��ynA��q;h����2[��{R�����r��]����t򘺾�'���;��=΁"`���sЫ���N�sͻ�ٸ�=�^'�;�uW�ׂd쁧�_w�Kf�uO=�r{��\�.[�kl�٨Ɯ
��=~n����gbPjv\��������cDb�|Y+#�=v��ʎ��Jxf,��\��ܯoZ���L�T�˲���ۮ�j��o3���n8�t=b:����1E�D 8�Sd˘t��ۤ�Z5��Z)���{m���V����ەa�;�=��6������q�c�j�q��j�9�a &7.U���EYhz,����zC���h-�)ׇ���A٤&2��d���)TP��GsO<v췊Ӯ�4n;'(5·n��ٝ#��i�5Ne � �[c,u���ɛpt��\q�W����9��G��mH][�(�c#�s�L��l�\.��e�7k��fB����&A����h;7��z�[��3M��˰��J�/3��A��q78��Ҷ��2r��)�,�F)FF�0��i%w2�r�e�8#MҘɳ�`3�Rkm9
ח;D,\�P�u{m��LK\�s� ���]p�uöah��ڐJ�#eJ�Yd݀ںYYw1۸)�{�z+{K<彰���.�k�ю��7�!ss��){h&�ƣ�!4U�6if��nn�'��H+S���wT��k׷H$Z� w"���R>�8���6������ڗ9d�3"�[u`����<b�\��+���5P&WG4�[<&F��V۷iGlt����{ s�9+��j'Z��h�`�x���v�y����0.�4��fUt���K�ۘ3aQK���9��\��887��(���!�`��8��,��7��>k9�,�Q�r�����d��w7%��n�sϒ9��4��V�L�W8�X�/�ٱ@�&�$�!h1{Z9lvn�hf�W��ƞkPT�`7rzy��6�f὎zV��1�Q�-�B'��<Љ�0�]^����zrGN��&ή�Gn_v���qŐkë�u���n�Ҁ���V1�2d��f�x��%������&:��;=���s�d�8"��}TV���u��]��=d��U��[]>�5�����)K�kE�ڇG�).�M)�hNy�q׭��Eٞ^��]AqS)n+[�9�N����bc��WW�kQ�8�w6:<�,���w!gG� s��5��.n�a��Ѷ�;i��<��盧.����7g���{m�f��vn�rܮ�����ױ�0gb5 �x����s�qh53��N���=�z�2v���$s���t��v7�`�]0v�\�/>��g��5�<�؆{k�ÞS�D��T�k����\����rK���m�^&��qf#Y��춆�[c5�Ӵn�x���(՚�K�[�T�ҹ�Y��z��xB����m=�;	��JEq����y6>ܜ�2�wYV�Ԧ��ml�ڲ��:�������iIȄP�e�[���$�pgnr�׺���c�R�j��g|��K��X��P8{�`aㆴ�۟+d20��[�w���r�P�Pqh<K�
6cN(������h3dEC��h��!�hr!���G����'�!�}�Y�jD�i��T>���l����a�7|��4��fT,�"�p�/�HGQ�a*Hpj�5췏>�tק�gGDr�a�FdCZGqU�de�9��h i�І9�g��qo��p�#�Vh��1h�?f}��C��E\"�|�����j�m@�	QA��i�� �����V���cHæ�4!�i��`�/k��xn��p�j�E����b�Fzh#���f�hO��,|�i����!��qPϯ8����ז�0��m� g2�u���Aknl&%�3�2d�䌗n�-ͱ�#�Yf	�@��?���[�{3	�4ͤ42Ǿ�9CH�BO�k(��9�x.��C5z-��#M���`6����$��}j�Gz��5ሟ��WCH�Tb�hw���U`�6�L8�C;�La��3�+�V@�����#�y<E�v-�ٱ~�O��q������g���� ��Iw	^k��,�3�1���n��Š�g�^�A=g�n�풸���:�Y��[�U���v�;�t]�z�5�P��H��{�;㦃7�l�ϯJ���{�������CCXE�=������E$CMB��2+��At0�?hnc�Ξ;�_�ut�f�h���!�w���w���i��0��f��c�&h{y��f��[�#P��$���w���p&�,��Z��PM^��k���ʳ��sE�G��,�f�4�W߷�t;��B�#�^':@���7P�4�>t͐���߻Ϋ#��a� Y�UtE����̩l�!)�:5��� 3f���N	y�t4��:~�C��v��#�_˟>����f�h�n�R#��}�ЇH��+!ٷ�H����da��gۧç�����г]#"���\?A��݃56C=L����M�	h�����:ONԏ�Zۚ�u�ķd�v�.�鵹f��pf��OO�Jt�����Z?}�e|I�!�]�����8�>�h�����a@f5�W|l}ם^?��N�dx�(@��49��V:kM2	��s�v�X��ߊ�FT�F��kHf�4 z��g�����v���ϵڐ��]�dE�_w��YCMp���B��`_��U�頌���< }��69��hM�Fa�v����΁M�m�:OQi�N7�Κ��g�M�dt,��;���xUYuW3���E�ן+}�B�#o��|<s�׷!�|0<�^�G�(jx���I�w�{8�g{�t�ѡgs~onqz���˹){�E �`�Y+[��7��ǀw��3������W4��=�^=���U�|�ҏ�T7��Q�B�c�|�	l�-;k�O�^�i ?<>�}���{ށ�@e�(}��]#;����P�a�������:p׸���3r�>V	�"�H��¹ݵ��p�@��߅�4O��U�CC8����2�InD�9=��t�k�Y� ,���}Μ��7ʮ�4��g�S���w��}αd�l��4��d�٦���*�@�-���s�+��A�������?̲;��nz��,��\�Qڹ�L��v��z١D��2K�m㳧��ź�L���9n���9B�����ӿ��J�4j��+��VkH�A�f�O�]�J�և�6���^��`k��|��������F����0����ί����.$G<,y|:#j'bF�Qŀ3ҍ��P@B��o>YCH�p_���+O���h/M�t5�Gƙ��yW��i�	᠎��.�"�?�XF��=����i�#玚���0����r2S2�H����Dt���"'����<���a�9�%i��� 0�ώ}�}HiN0�T���3�w�/stt�����G�s���B�}����N+�#OH����G�B�&��0$`�$ۑ�#q]	�������8��ߺř&V
�U�ïj �i#��PdW3�Ck�؆�5����t��h�q#_Zf�������~��wVC�c8%�T����3����Ю�)���ӈ\^r��E�r�ҹ�kތ��ّ�s�����*y~7Cl��1�ېiM��>m�F����C��,�I!�,�da��-�����C��29��+����<��#^#�P�gX��+�|T�g�j��|k�߸/�}������5��kMwk��/��Mv�7i����V+Q[st]-^�X�Y��J�V˓��r�;˘n\�w׿�=�h2q�	������EC�á ��3�t=�:�qtٮ��_��a�=��������4:p�ψ��ϴ]4>h0ִ!����q�HL��ЈaEH2��.��j��C�WM�I'�w��|���>��y���9�^v��\��0�5|y��aIj�D5�!ޕg���MT
�$h/��`�V5P�+7��}�X�uژ�Cd�DK)kJ��(Ў)P�[�X�bO^�P�YA�Ϲ��<i��.�L!��/�C~$���vF}�� n^����� !�A�71١�ⱦ��['�9��40C=����X,�a�� ��\5���
/1��C���o��iG<�N{~𱧄t���Z�������J{��`t鮑a*��#۞�\�b����~߂�d��#�nh�ثx�@3D|l֑d��s��E6qR
83H4�!����G��|�5�CAw	�.��#Gyܝ���b�p��t,�GmT>8|g��ޮ,��	����AO����W;`a�}�Cu��2חk�o/�� ��w��+�������It�Z�һDǬo{^G6M�s��眘�|��8�d�v��`}���������@��5��v�]h��\�5�cVk-�b0��[r,������ϐ���v�a�^0��+�7=��Ѷ4�͛���,%ڹ�l�4���.i��V�f��Q�`��wR��s���i��(��@���]qrG%�x�ls
t�Fd��uc��^z����Xh�:�n��2Լ���c�ַ"��UKs��FV����r�$��'�������S8S��N�Z����s���G�-v�m���벽�P)�x�֏ �PF� ,��͂k	 "<j�n���bu��%�Jh#��
5~���`?gÜ�fpvkγ^"�f�߸���{�7��i5��B�O����(hg��p�Q�77C;BϢ��Ժl�>�.vo��:7x�/N9n�Y��#����A�>��Zh2��f9���u�~���������9�+���s���}�F���O���xϗ�m�B�c·�{	I)'���=�a�G�0��e�4�Br�s_�+��uІ�����uO%ne��\#ǄK�U�����Vl�#N� {����-;�C�k�n՚dY�g�8G͢c$�nC���!�׎�]�5��7{�} !������� |���hdU燐���%�U�M�n�6|C ��s��ѿ,�/a��wU��>$�@�5�P�|m��N���p]qabp���O|o�+���h3A��u�A}�_y�
J_�h���Vp��`�+v�Ձ����@�:h�=�;�8���53��Տ�0Н������_>�_��a�Ts��tƱ�,]�����g��n�wl��)�s���r�\�Mb�qv�h|�����M���hk\#�,�o>�߽:��uYĄ4�����]���E�x��0����0��Z��V:kL �OMY�"���}�eZ�,͗\{?��	���Uznoj�vG�h�ݯŌ�zF��g������*lR�p'w1�ޯ�׆̵x�k�= #p��R��o��:��,�^f#KEEu+�Hs0���F�MD�u��� n�гL�@�b ���Κ��P���k�6:k�t�/Z�9�@_x8k��ahk���Ee(�bN8�� ��Ȭ��<[����4�����>����Y�i�/N�HH�GM�u�k3��u������q#��>߱X�*|T8��kÞc�Ӊ�L�`-Hq�4�A�˶��|�8xb�t��=���@���doP'�}�7A�`q�4!�յf����� ��'�?�"��ri�*�<h/�;ǂҭ5�i�����C� �!Q� ������G6hCA���߸.�#���t�����|~�}ly0y_.w��p�F���4,����vy#A��%|��h/}}6BtлT�ņ�"J~�:�}ߊ��m����#t�IEɷ=�j��2\y��S��X�9�qnқ��k�۩"p�p�:k�h#|a����N��^=#���0իt=ht�g>㾴4��C?b�+��b ��~6��Ƽ\�np�<�������U��mI�`"��{=X����vϜ0�uQ�d����(p�o�xG��o��چ�-Y�*���@o]k�3L�e���}�;��	=5���b�C����47�>Y�c��'i�j_~�OXI��ъԇhp�F�C9�D26�u���p�F��ܭ!�k;�x��>0�O��� `�3>;����r{S��b�Q�}�"�nL�����+�r��,w.�[�a0��\m��{�D|���C�p�V\˹�ÜE���f�����a�d�bЏ�v-*����G�a��I\DȔ�M�"�5�F���<�9���@�F}�wH�!�z ,�������7CF��7��74:��;G�֍$��t���xx��Y�顽�t�Ԭ�4T�f�D?'����(�e���CM�9v��e����>�8Q����!�p�8e��.��S�W�wq�5�$D���Kj�>����ii�C����C�r�5���t>�V�dx��K���0m�{�f0����c� u.&{5R=P��h1V����̌!m�����X��~]�3A�Jή�����OXv�Fc�j��?9��p��B�h#�饗�+��5d3�<��_}���7։.�y��G�L�B�ۢ�5��A�X˲4��_L��.���)l8�A$Z:G�XB�}п{~��f��@Gh_��uʳ�#"&�Q�0��IC3]hq�P��^{���#������C$�Y:p�4'��}�q�K�_/�<h#����0Ѝ��i��]5�CC��� ��o���`p�	�@f(�#Z��XvD��b��:h3�'n_�}����C�^�Xb�C���x�٬7�>Ⰱ�t�߾�X�֚ŝ���S��,6�M8�����C�E�?�W{�� �2s��GD����L�?}�]����N��j֟�Ή|߼��s�&��w8~�9���/6n��p�p�	�Y�>^�ܽ�h�tC�_�ǻ��ss��^_��U)I�m.d��s۽�����o��R��@x���8�����w�W�*Ղ�!�wT~f����Ĝ��!�"�#�_Q�}��i�M20��B�<�����{���櫡�A�7�hY��K�X�̴>#��4����c���p�jp�f�,5}��\��cĞ7p3C��3�J�Viv2�����\kb�\c����\%�:�E��%�u�6�"]���O���q|@�0�:ٛj�@���#����5쿸��{�]���Z14!~L���E���n�������D����@��ZG/���\#���H�0�8G�I���L�`�Yq�R)��Hé4!��!"Ͼ�f�a�ǻ�]w�>2	��U�B��D#�;�P�ׁ	��i����pX���4����+�8��L�-O��g���� �Ŏ��P����6!�(���!�jn1f��D>"����e��BA��g~ߍ��|;I##�M[����ދ#M37�/���A4Ő<w����5�C�5Єa���}���B�D�-A�hp��b�s����ӓ۽y�K�:n��*F�Ҩ3A���`a��G�*�(��?qX����4"�&���5>�`�"=��+1�GƷ5г#�h[���x�MHCF#JHpY��f���"�_٢��Xj����m|�����w���+�"�5��>j���wte4�C�0��\4:���X-�#Hpr��a�3�ﺳ��P��*�oA�~٠�q��FL4����d	Q��Ŋ�戏}���t����������X���!X���Z�h�v[���P���f�����*���5ѕՙ����[13�n.j�m�[s燋봳:$����Lכ�����Wn&�.��n�͞�vx�xu��Cu����s�v5��a�$�m�;Jc��rG���1r��������cn���6-�&�[����`�Skn������Vj;v��VYx��1�1���r�Pu�쁺�ЉjD9���J��N�R�E�9�5ݷ3[�:���n�	ls.�y��N�]��f,�];Y������!{�!�{��x/!dx�4#M}���t-k��}hY����g������|ht�����_����5�ZE�ƈl�f�I��<>d�d �TR)P���:�b��7���a�-{+x>W�����~?A�����{�Ô//yt0�!���"}��>��B�5��dC[��Ň���v+շ��Cx��[�i��{���S���ZŸ����I��g�L|4O�>�;�$3�B�9��ZF����]�7Ct*ӻ������@�g�,E��mo�@�_{�ߍ�5Q4�Y�7D�����M��?	cH����ѺG`x��8@�e��o�_�Lt��?s��t4��rQ�A��5߷>7\?�_f�8l�j }��E�6t�Y�3�����uŤ�N���5|B4T�h#C/�~?.�q��j$� �Mi�9g�Vp���p�4��>9h_2=_u�v��>7C��(3P�����+|�hC�҆�@m���M}�獎g�C�4_nP�N�f��1�}�9"A�l6H-%nyƬ�v�\���\V����Bv�pӺ�wK�S�#�GI��=��WH�x@�����kHƃ0��h}�������C]!�e� �g�����/��Ƶ�F�w���|a����M~�����@����B�WH���s��)���`mô8G�0�<���,�_�+�H/����ȏ�d�b���o��ǫ+�)����N;s�mlC>�ޢ������BT��zf�$v�n��K]��_�N��t�qPdLU���t;|t!�$T!��?n�� �<4��,О�0�����?��������x٤G�s<K���6�$H���]��0��!�BN�~�Bht�C,��a�L����jp���!�5%�������NW������ZF0Q=*�a�s>X4֚	��;�A�_| B0�ƌr��; C/R��f}���$c嫿pXxGMC�Z����s�\f`�5��*�� 2,�8@��V�p��X�=����y�g:hK��`��6:�k��g(��B.�CM?chY��بg�f���g	U���B<;ל�����z�s�m��r!}����o�H���(�(�	��xk�9w8,a(Б5�>@Y��ߴ���x��޿���>�y~�܍i�8�,	v����0b�l�eur�u���썺���qk�1�(���x������,�K }�ϲݍ5�{Y8���aE�^^���8����Ϯ,���?�,	4I�X��ޟ�i�� YY^_]���t��=���HĈr"FH˒+���>�A�H���F����!ͻV=����߾��]#�[��">���~wC�Tt��yT+���:zh3A�$�;=�;�b�H���G���#�M#�:i�Z��}�J���Q�.G�HΡ����Zt��3x��VaF���3Bg���(Y�@s��s��&����۳�S��sI�JsS'��3.����0�:>�#���V)0��� �7�ڇ��Mb�h�c��O�5��^�+�F&\��[�6�T�n�m37���VK���ի8y�U�2c���5�ԁ?vi��6�[�4�� Y����o��˅Y0�Y�3<�Y�N�Ŕ�N��T�^o{���1��tgl���!���C��Uѝ����=�}�n]��Z�
�ږ���^lX7-�^W�m�L�(���}|��*r����J�s~�7��yCfl��߶Gٝ����n�%��W%���i(<+�Q���>��xk��zl����Ôe����f��}�,CAά����]�S���Nȩ}�!��ܗ)�C����bsi|8�`�mYD����D<����RY��ʚ�U������e�-խ���:�W�	F�.��E/Oa��g�-�����{]0,��h�вz�Ѿ��ۻX21�6�$�
nCy�o��_��/�L)�:���K�K�=����Ϟ�b���׆�Cj��?�||�Yؽ�̕���dS��[��LKt�:�?�ɒŽ���i����q;�&�	;z�!^��ށW; �զa�J[��ᨮeI���Ǜ1��o���_O�r��r_ZP��;
��=n�t� �͋��=�F��?R�qLg�!}�V���nb��xa�{����.wLk��if�}U��SY��I�w���8�c{v�O�k �:���<!�K�09&q�K��C3PG�s�M{�x��h4!��{51��&�=�J����>�>LD����P}��0#I9h��p]��ssy(Y5R���t;��B�
г� ]�8l���@����c�,�p>�Џy�b�>��#]�B���{99�$�'e8��4�f�4��;�:zG0��1�08p��go��w�(������c�	y��G�#�H�Cﳘ�kH~!���ޣ�����`�(П[ӇH�B����P����P�6�b�\�u�.Zk[I�A��ڰ='���y�7)�����{mB�2�XF��H<k��Y�4;�g��7P�֫�!F�U���]��c@w��b�����gӻ�!�;� ?Xd��sw�V4|�����F�����ѭy��d��j(��GMl_,�dx�3���cz�%�ﺉY36��Fm��C�T9�}����CBڠ�����+�:GO�,�?'��47����k�L���}�w���r����T;�G7�M���Z��>�����=:x�!I0=���F���`BH�ʹ�O���L�I#>��aWoޏ�k�><��U��a�w]#d>5���<�=4%��c�����n��З�1*����0�f��4����o� �&�7��t0�⬴�5P�f*���+���B1GMCC޼�X����6G�1o}x�>��ޢ���4��9"@��t�y!���SE@w���I��O������-)�;Ѷ����r`�V����F��	�${2˱e_ǿ�u����Z~$�bf��6�F��w~)4�,. ����鮚�D3L����o��u���A����j��_s;��wP�9��F�Ԭ�j}ߺ,"2-#����"��V@�������\4!����P�3p���]���$��f7d��KU�6LY��g���q\�W"E��-B*X�+mge�L����߇��>{��Ko�{�4��44�������ȫ��,�H�B,�=����}5h�'�⚿�3�7���x�ր�+5d|������*�ڮ���)�K0��RrA�4���,iǇH�G�w'��i;�|�8g�'),�����h���B�D���Z�@�g���|��	n�U��]t������g;hp�GH������Q�\)�8I6Y�C5g� 	�|r�|l:G����C��2#���j�"�+�A�b;��k���>j������ә��yd	�X�&�߾�>U��#��6Q{8h^}����2F
*Hn��@fz�Z��]�� ��lf����,��=����C5W�g{���� t�f�������NX�ϣ�U_9L +��o׍?_ 49'zmk:�����!dK���ϴ�4S$FԐ�5=�Y��d����8xm*��4-q��>ߐ�k��E�÷�O�jݭ j߸,�i��E��42}�n�5���l|k�U'�q��z'f����j��9��XA�N���*3���_8�-�{Q�+͂U��A{��d��w�.��-��Uүf(T�z���+2��2@, ��]u�跢l�U�By���YtW\���ob�pƻV��lruD��q[�/EJ�x��1�;�eD�o���-r6ځyl ��lٻ+�z��yM����sq�ȮLKg	s����W@�;K5��(�t�P�t�A������fQ�Ksf�[4 ���]�P���wn�$�r�]�^N��3T�]>���1:�u۝b� ��b�g����e#4t!�CXȴi�u�c��V���˰+���k�r�=���hZ��q}C�^��,�	b��2��t09�Vhs�����/�<�#�j�!�ϡ(t�}��9��œ�ps\f�GM@%�\Sz�Xh}�r��|b�	=ޞ������5��ޟ���t��.%��t4��b�gm�V��|@�p�~��B}�@�4���C��+㦐!���0֟���t���}�Os�>��x=5�2�d|{>�D�A&�=&�*7��H��A������h|�V�ӎƚ �0����I'�z:8hCC�n+���-q0!�Y����b�a��b�Y�`�����ť�"�3�2R�o��΄0���_~ى��3�g��}.��'��]����\!}ٓ� ��:F4Ȇ�.�������Ad�),�%{��w~�M�k��:@f�:k�﻿S��j2b�$ydi:Y���J�E�"�1������8�!�
�i}LQ[;�h�3���!{������CB�DѾg��k���w��`ՐECC��y�#���t,ױj��r��
��������S���F��L�*�׷01=+�]�S�Q�U���)���d2d�v�����b��d�(������j�Y�#��1�|���A�hpӊ����x��[�-?��9�:H=<�>�f�7�٠�uX������C���PD|q�����1Bd�(a�b�,�8F�}����iz�8�^�����f��]�$�&b�KtY����
X��s�k=��{�O`�!#�ڻ��v^�w�Xc�f���c���+����1jN8@V�����]iB�D$��Y����_�(a����{�`��>��@�^����Gw�8_�?$!�	�C�{ǣ�6qF�eD���kHf�<��`>���yC�?!�f�	�Y�#�
���+�D��f��.�|�OGM|GM�|i���c�3��@��iܿ�W�>%�k���������|��l�ak:�p��-�y_N{�Q�5Ú������/�VhCVC#	#�}���\4!�f!-PDY�M��`{˦�;m��3��v�w�v�~>�C�{��&�ޚg�k�CB/gխ���A@Y�š���"&@$	is�_	>_4W�1U�	6!�E˞����KvO:�C�!dY(�Xw��VڸB5	 }z�������t��r���!�\���Ϭ�>���%�̦�0#ND�j6�ܹ��b��`z�qp�\dB#Ls�.z��`�A�
D6�NP��7���>#�!�����K��\!�@�*��������l����AM��0����X�����4:�}{�}U���rP�*��h>��A&��H�l�-H�G�P����,Ր~���)����s��3A�2P� ����.ٺ4<��p��6p����р}���;�N���Hӧ�G��q�t�	����wW���Hk�;j��м�rE#�E!MÔ4�F�#2�}��� i����dz@���n�A0*��}�N��Q��l�|w-�^��y�cH��G��'��ͤ���~؝���zb��a��)!����~�m>��1�
<0�G�CY~�;���4!��+������U�C�T�B4;�����I
H����>�Ab�.�cvp28@�E{�Ct0��@���¹t4���<� ����8IY�&�����|��h p��g���tu��g�[������޿�P��{v��WhZC���~��H�n8Kb!��i�����#H����-�#����fϟ=�c����ٜ�;�z��XD(� 3�{��`}�}5�0��B>6hw����qPf�C5�f�݈{���-�/�����l�[l5�	��m.-3���z�c�[���vw@汁�k�ݖ�͇�P�(�"&8�C�-Pg�!�������@�!�A5�A�*͛�P��"�wP��:@��������Ɨ7���@x�!6Y���zU#B� �Hf�j������HZR5*H��F�����6E���Z�N?���'�9\>��7,�"�yz���*Դ�3NP�A��~ a��P���+G�W�'���H�Bd���5��ә��h k�N���'��)%���,��=j��y� ���M��J9��,���\"�>4xouPF����}�X�F�/��Ʒ~�v0�XH��?b�(a�*���>��k�Y�؄$�hd��$x6��2K-�#�k���гo����{�x@�{��U��!�@�"6!�8���tcei��?!d#]�ύ��Am�H��#���;)�ߖ����^�s����]���&r������P8M]���Łö�pdw�5���"�Z��{7f�@M��>���0w�]4=���u�Y�Ü@��DFH�Q�#�Gߘ�0�Q��`YF�?}#�|#�pІ�Ȱ�(�x�����_�n��	��Q"�7=�`tyP�Z�f��=�^PӤ	6l��@�rt}:�蘆���L䲼�[v�6���p�l�{�s��T��[Xdp���|�x�疍���C�V������L�@��!D���ߎ�iy��d	-гC���|F��׈�Y$CC�y���&��Fl4:�i׏b�<k;���]#���5G:
hvg�=���[�<7O�?�1)�T��y����>�]��:ތ�wn��+���o�Ő<B>,�8kT�+��]��J�j��DB�Nc�]5�!
@{4-�_���z�e��*�zd�Y�Bs��?3a8(�#�j��H�0�:lL��s~W�#I!D�,����������A#﷘}.}���6@9���M�4!�B�f�w���5��B�w�0�5{|>)+E�$9!�=��^Շ?ChF�|΁��|��j�����t���8,׆u��Lqk��d7>�^ќ}4,� �}����Ͼ��M�o��kH�vexA�7�Ɵ�_�zW��D�"���&�����*j�����kuP��j��ep��������V=�#����a���� ��� ���V�4�4��|�k���H�@@�!���5s�3��/�f��PC�K���PC���ռ,*=��V�N�A���q�_�Mۥ,�o�U�����`Y��O�ͬ�t�&���4T�A;��=�7Z��P���f�ƨ�����͟�7ϟ�]s9�B�;6�Ƹ�m=c7�9x��!E�WoqcrVƹ����r��H�&�\��ڸ��pe
Ŷo%��i+r�3����8�sn�^�3a#����t�+Ԃ{v3M��}�x-;�J��{f�gl�'����CY��T��:�)p���d`��F3E��D�D�1[nڴ�dy������J�D�8s)ZE��m�5uV�v�n��Le6[}�g��~P��}��;��r�Vh�.�#�}�����(Y�8�e�qC^�}�c���y���D�اi�y�� >�&}A7��+�WMkHf�D49�8�I%��D�$�k�3���20�#�f���ن�uz��w�WH���Y�-x�)�7C��5��Z�|��L�D�gDU�d"�C��򱘩f��S�}�<@��!�4}�ZT�Ԥ�L���'Mh#�@Bؽ��}0a��k�W��<hϯ�#k>}�s��cg|xQ �����Z�h#�Z-a��ܖ��nCr���О�O>]�Lăf�)��C�t��l�j��A��G��糮�a�!
 zib6�z{~wC��#Ol�6��� qp�������;��]q����?L��(p� ��� a���~?yI�ܩ
R5�VD"�����Xh.���#z��P�x  �𿽱r��~7C��=Zl��IӜ�`C�|A0Ε���k ?����4��$�4;y�0�s}G����=�^�r��e���[�{c۞�i���,���s���c`�f��c&�\�q��@F�C3�00���خ���G�n��ͷ��>�]	�YDe���t�|�8��zksq�菳)e�4:~�~!ua�����~X3�Y�C��"F���3�Q&�F(#.G�8l����� Bا��VǄ7������C�G���%x�ׄ�fk���{{�XE��I徭c%��������YP�9�ӝ��F1���7N���l&�[/��L����z�	�ܺ�P�$@f�Eط�q�~޼�< 6T?yx�~Zh}���a����c�ƶg~�׍{�C=Yh��\m�������T�, Y�L� C�_��4�5f���C���oҽ����s��!��m�ϲq�/}��f�GN�6����w��B��k�Vp�4_��V/A}Z��,�5���9$d��l4��>5����#�oy�'�WJ `����Fg�ǧM>:����/�n�z�5f�,Ѕ�Xۿ��@���hYdA#3W,�O��s�|k���e�_D>5-S�C��>�������hǝ=8"I���Ȳ=���|�G��"7U���ٝ�H���y���i^�UЃ��5����4������gz�i�Bf���,ϧ��i��ˏMA^g�}��i��m�Q@���� �P���k/��q�u�6� ��[ruy��IΝ�naD�E#*Q`��g�|O\��a�7~~_K��iCB����}v��<Ik�(l�͐<ws�V��I����
��p���d�29���*�`a�O�a�c;�_΋��]&)8r�4f��CϾ�=�o�<�ן��顖��5��^t��:h3]��4!�޾q_ƾ��;�5�j��f�����ԏC^�e���B:j�Ag����%8�e$Zr�f��hv*������+��!�hN;�HE����w_uWH��Nϼ Wv.�}���g\�!�bɊ�d�|���Ԟy���jg�~�K޾�YH����J�[0z�u���n/m
>��;��|;?�t���"�3��\�	���-{���WxY�f!�����HJTq DNH������=���FK�������@�5����#���g�)d|]��!���i��4\(��`�,qpЇ��,��t�K�h=ϾV;�V��[�f�б��i����j(��ew�����~ 2�|�,x֑�Q43ے����9k_!�<�'ܾ����~� i��4�}|�����~#��4���`�|���#ƙ�F�9ϛ���Ϸ����Σ+c��mǙ.�"Ogv���>:��^]f�����6���#�xx��Fk�.�����D,��}�h�G���he�����c�C�"O�f� 3���f�������@��,�������xzp��&@<p�~"����ɢ��]����?32�1�% ��{���5'������a�c��=;�1e�滤G�]|F���0��ύ����k�c�����pX���}x:�,���B�X!��I*<�1:tXM8������+48~ 2K��g�P�3%a���Uf��d?����#���w��>6sǝ���O5Y���P�h��b��=��h���f*ᡙ��hdT�9��C���`����i$pՏ��43��~/h t��]x��xf�"�͞�9k���:i���(���|���_q�/� q"t��r��]��p;����̆]�":pf[e�:��X(�O{��59���~�)>�(�G�:�N�{����{P7�1k�uUT�U��v��W��@�z�`�Zhh��>5��=�V���.r Q�rKIŀt󊴋4~@]�j�}�;��FQ�h3A���zI����t>����adrв6h/}}Հ|�a�G>��4���ߎD�6�D=��# t}�{�wۘ�\毆6w��rA�3��
/S\h�h�M�4n`�u&Q����^�3A{mF����P�d4C�,�3g��Z�k�YGMC��W���u��Vl�~
5g
65i���Vg���&_>4<z���S�?g��c�>bύ��5|B� ys�䗋p�"�r��<~�@��L�
���wɘ2�8�����vu��C2�<@�����0�qU��T���a�]�o�X<~:~8Gӆ��O1Y�ϸ�nD�p����%2Ǘݐw��w�aw���ZI�tJ%�[p�"0�#"$�<5����j��;�ҏ|�5R!b|CZ�k�g0��.�j���>�~~�d3�S�k��@{�oM����g݀a��^�}46��=!��H�j���*�>�;��)��$7Ct�B!߾#�}���@���w�t0�zj�	j���~V8k�
����>�;�U�N���6�d&������+;������6<k��3�%4��Y��&�l�
p��w\'ˆ��kH�A�<�ſq�5�x�q"0г_$&}�V��+��x�Y�7�� #f�Mj�~6�h"A,���?MÆ��J:5_!�h������Wӹq�����b�'>�D���P�xjOFw.�ױ{UǓd�1L���&q[���#�J�W����/��wG��l��+0kJYwK`��a��|zٟoxN��۸�n�R2�b&׃�5[tdmq����Æ��܅QM��t�??#��%M�%�n�������vݞU{dĕx�g=0�{��L�3v�Hf���k]e[w�hR��?6��5�C@����	�m�Zoo���7�Sj~}2���-�LY���ݜ��|�^�<�g$5w����t���l�wiq)�I�L���ϧ$�G�N+��en蟷�K�88)c��lء�yLK4��TޙJC��Q���=a��pȽ�O[��"�w��rb�j��7)-w|1�'d���������+��z���뺻#�&���Ӧ��Zc��1����4m�_��=M=�VVy���Ȏ~���ZЊ;;�o��1��E�������y���;��p���d=}��7��2z��|S��{�/q���;��92Oe��ܩ��/�ۃ{s)������42��p��q��k��j3}�������;��eZ
��#�n���&��(٧v\�$�L~����r��+�[v	luV����v^z��{|��33p�W�:��㑻���Տ�~9/�!@���Q�|Xc�yog�m�y
|��ø\݉Uҡ݆%A�Cv;�\�P`�*�e�h��-	�~16~!�H&S-��Հ���3�<��t�yf��n/0�S�r)im�-���<|I��CKM�b��-�X"�[�套a����WYk�!�E�)4&LG[e�B_�g*>�s�h�9�͋���w��nQzy^����M��-R͊�L��"FV�l^ס�y�g;aû\�\j�ľb.���CZwc�m:�TXT���҄	I�MЋ��oC�C��Ӻ|<%Q%���f�S7[H�X`Җ���x-N�I�ܑl=v*�a���s�.6����c�L���lX��渺�,uב��[6ܠ�$�ҡ��
��\�P� -�@]w[]U�F|n�7=h�<�d�T���X9�е�CMr
ˋ3��V��"���d�e\(;��]JQ�;3܌u�9\����ݶz�]-ְ����a[���Ű+�<��ٲ�[���$9��>�ōҗ!p�8V^"�Wn�>9�kd]��_e�u,b��)2KvV���!Nͮht>���X<�'-��K�1�m�͹� �HBo&8n��P��+����{cT��Էuv����1�hiinsHԮJ镖3m_�<r�����Lr�y���P�,5m�Ol���)	�IpY4��R�vS
,���r�/CW�؂ꕙ�M@�k����Q�筈����
���8ψ�e뱸s��	�2s�.#���+�':�\6���U�J�:�a.�,��M��[&�9|��ܶe��w
��;,\�74歶u\@��sG�[a�e���J��a�)�V�K��6�<�u<�||���.��z$�sK�yw ��ڎ�BU���M�:�qZ�sr�h���-�*d{q0rM�k�ے��t�l�M�,�m+�����[��6ͣ�WEm���k�N�mr�B���;j3YR�-"9�iMqa��].����b�U��a�nz��E��I�E�o.y-�=gq�!���h���=�7%��is��BmX���f��r����m���z����R��q���G�2��(���9:@���W+ �nj��y{�ap���YqK�]V6j̀�T���Z�:��(ʑ�m`��z�:7T=r��r�+y�]��e�p���!�E����I�&����kx��/U��FWu��8�@�(���7c/Lj�F�_|fn�Y����`�����H���w/��]���ܼ݃��"m��%6ڸZ�
��F[�)��Ĺom����^�4a��qg.D�f�mVkZ��mɢ�lL`T�dl��U�)Ε�^���_���5dY��"�w�ŃMp�D4���B��կ�� �DE�屆�M?��k�.([}�O��.#Ch#C�/�y�#��L�6k�4=>K9�G0GR;�8V���ϐh"!��~�ep���ًU�d������[Ç�߭�29��]20�H��47'�W_�M2!�u��O|��/yP���W��g�����5�����@x�<!��熯�~q2F#eGP�h7���Y���wCN��4���8Y�z�;��e��#I���勣��0Ї� >�H��ƅ�� x�/~�c�CǤx��촀�A���0&�D8MA��i�u4!����>�$[|N�����w�}>n��;��W����s|#���j��\)�Z�9Y4�3�$��V�@U4��7ٷ��X�����s�Af�c��f�;Ɯ)/4z_5�%<�I)���^%�&b�!z�/8$�>Z�I��HZ�n�4tw� 8r��a� +3���-����:,���*j�%39��V�4�V_�<ߚ޵׉TAzu�TS��D�+ǁܹ�t�P:�$�&����$wqN�� ���^^0{.�a��m�����p��ai����sF��=�3&i߱��gW@�hS��3W����~X��@y����=#6LѾ�e"3P���pT�Y��xe�IoMV�%^]�������y������=��)XSyj���䩮��m���lAISY���Nݱ�2��#�Ж�O�{F
��]����rLt����k��cl1q�t% ��'��
(� ٙ˾N^ρ:}�_]����5�[8�fW��4�w�U�V�+	ظ%7�GKs{~�g{.C��EҤG�)��b�+'� _�{���T ��n�\]�M�u�лjg?z�'��y�]יV�-��N�x��>()Ѭ�=I��-N9x�av�m�E��a��<<��ۃ�j	w�y�n�0��L1 m��D�����y:�i�v�p���Si��֙��)��T'V{�r�[*È�;��^_� h
	��@�e������ᕁ��^�p������t^s}��FS4�����3�u��;A�ִ��/ 3���fbJ�XtN�t�L���'wz�Gu��y�M��u��pcf������A���b~�Y�{��U���������Ԏ�3�s�S���ø[��(c���Ɖ�uz^���Z������f��L��������
���qd�]�y�T�߁��5�C� �f��+0l�?M\3I�#����i?�^�Mq_k����;q^�K��UE�B��9��� t�b:N��&"�}7��/�L)#�f�P2����W�Ğ^�=v�F�@�=�y1���h��W<��W6Qe�L��:�J8�����0��Y�۲, K�B���.鮦���@%A����[׺<M��ڸg��>i���e��)7�N�L��(���xܿj�wޞ��Y �+`L�E�H�ټH�ٓs��+1[~�
��u岅.��^��w�f*�-�6�o�����z4��Rv��&�F�DW�J��i5�ֲ�j����8ף�f�s2��mu߸!�}"���8�pz��XmS�P"��Z��0�Z]?+��z�L��:��p�~fk�	�����a��������0��mb���x^fLggo(��=^tW����43�<z�r�b9�0�>`���`:��[@N(�*�<2��6&�y�޳�L9�;P=�n�B��X*l�ϸ&*�Hpk����W��9���m~�k�4�=�8K��ӓvz���7�Yh�߷���B��(ؠcQ��K���(��@^��Dkb9�ˋ�"�h���y�M��\sP�&��Qu>=|_y���K#�p5d�e�T���ez���z�md֗9�{�`�4G��D2\�2�
H�Z�wh�7�u�;��>ס�/xg7b�̸��B��Q�����Ղy[:��	^�kp�RE�GU�����$HT�i�Yb�/w)w�m����|mt�M9�r����$��w;{��Xiӥ��y>�9�I���Mo������θE�+�����~�]�����v��bؒ�v�C]�ڽ��s��E��ߗL�u乿n�u ~V�%��Ml:��^���4���C�]_z��ꕢ��Y~;|�f�WP\�rӀ`�v�i��⽇�;�i8�\n�hw��/Z탅y]���R:�5��Si���ݚm�}�k�KzM�buD�z�X{��D��p�H�A5!�-2��[�m�Q�n�S��W3]nݬ��c���\�Q=��Z'#�\���yKfQ�U��e��mr5���'��p�Hq�`.$���.s��q�a����k�<�uvy�����]�ٗ�e��[�7��T���1��)��\
���<�C��HKZA��Ac7mx�W��(u=ne�z��8bQ��]+@���U����vH���E��&��n���݃8�D��&�9�\z��k(r��Q��l����?��ߔ�5g2��;<�d�{r��r��o=�uh�~���/H�_�y�hNʬ�Bm��m�TSn���`��Ǜ\��3G[�cǞ9)�E�2�o/^�����9�x1��V��{ƅ���"P0�	$�z��D����OM�ǎ�v(�㛙�
�k��]^^�޶3|��{����g��}��$7�F�L�RE��ޡ���.�5|����j߽l��?�1��?v�|�l�x�獬{��U���}��{�Yp>�r��tCH�%i�tQ��}�w_���2���W�m��˵�v�
�,��s�t�g�th��ʽX�k�OZ�S����>|���mKi�ZBd�7�bvup�Jd�\�4ODb���Pm���j����O4Ku��ԛޖ�ڤP��9ܦU�y�GR���+&�g�K9b��x��^�"nřJ'��o��2lS`��,��Ì1�o|1��/�㦯���]�Vo1�5��Is̎Ӈ�v��
.;�ܖ:�HB��s��x�wz�Lz����W��$��)�*a�|q>�	C��kwS�f������	2�� Ϻp�g����_+�F{��~~x@��*�5l"��G"���F�ۿ��:w�g+�TOMqs�7��׺V��W�(j�K�ܯO�����n���z=Fo�C�~�8}��X�@!.Qj8�A��ƙ�x�õ���u̏�_g��#H�R��\�g�uͰ�j��^�P���.��; ^ǋ����qЉ���v+)��(���*�29��:�o���54�u!6�앹k��34�I]:_ZR���y8�b��b�"�_ރ��N:N9�K�[�},���1c5e�rU��Er����m��ܷ�v%��j�?��$Ѿn{fp� U����8xF&���Wpʵ���	~�GE>���<�XE�<,��;�жX��i£`缮O����}�,�U�{0tj����rǀ��S�S������c˧	S��ή�^�mE�j��@	�Ū*�t_0 jX�����;��g�d�<rT��J_�r�����'����w	��RW�M��we1N����Ž�,e����C��;���CR�6a�cN���[0�y�����	�Q�7C�έ���j��X�
���4^���<�gB(2:'��:�T�cNI30 ��;{�1��shc~��nU�����C����Ǎ|�{M�h�`(��{�e�nz����c;��v:c�v�x��&�RE$����F�$=�����v��������6�ڭ��C9���:Zwj�S��g�z�`c���̇}�o5޼M��E3$bBYk��\�kOE�8�M�p\�Jn.G�������3�n�؇J��D4�&�ݾLS�#��<�K���T��Ȕ~���
��J?.̏-�{;������q*�޵(a�X�3e��|�
E�cD� EH�s���eë��y=�/��W��^�-�n϶���Ūo���@}o�ǽ���q%
Sx'H�|)P���o|�L 0�r�R-|Cb���]�ٞ���Oޗf��=^Ӥet�j^����w��~['8x��r}�F�ܷ>w	� |�	�R��w���~�w���mw��������|9Og�P:����Y�p��1�v��/i�4��>Z�ֻd�.�{F栌�07휀~ro�}�\�������
��!'���|"
�*�A4V�k$�?>�{�c�>����@�-+!�e�H�mJ��s�1��nD�%.>���,����V^_���EH8e�f÷���B����wp�[�{U�j�5�!\J(U.6)�{t�p��u׬:�JW��jݳ;�,.׃�vr� ��L��F)p��=��gsۢh>1H,4緜��E)U��̝�&z����\U�{�8������^�e�iX:��'�Qt�E �I�.$0�|F[��O&��C�2m�2�y��Ξ��ǰ�V�`<��^��d��^��7]�҅bm��lK��{{IV���>��HH��JI���A5vw|�q�;Jtvp�׾�y+ow�M�r�w�w�o�G��s��[�=Uj/������i�J���L$M]�l���s`�g����U�8]P��뙝����L�����"���;���>����~~�\93}�3�#�>B�N��*G���4���/����KX1&L�/�}����]v�7��C�
y.�9z�b�SZ�15�����}�囶�ꬶl�I��mI~����v� �@�g(�D�m�QG�nb���0����L�$�<}]��7_��Ӡ`IA�Z�-̠��1Q�d;��O\O^e����.�jxϝjf8�7n��u��{b9�tv���v�U�g����4m���q����<���-��/M�Qr��� u���H�2���h��"��GvR7�Y�E��C�a��]��5׷5� @�7�lq��fʍPضJ�	���{i]�ݞ�eJ}�[�.zz������ջ���4�%b�3��^o��cJb�9�1��۫�+�i'��]Y&ݵ����Z�����໩fN�S����������s��e��޻�q���}t��o7V��}\��-�X`K���6����x��~��m��Wh�>�r�Θ�����mn��<^�����t"�aL��{���%�ԏ�zɠum�*�x�y|�3��,��H�C82��4�����wʙR��w�~��Bb���4�6���v��7��QU�w,I���"�3��{
4�1B�����J�����ڽ����_�ҧ�JpADU��*Y����珦q�0V>ݻ�ۺX:����%���^�X�>7����!IR�ҤYT�m�&��	�nL,��򱛛��`o����V�!XݻR���Կ,��V��)�~ZS]'�9�͑Wq|���)}U ޴t��*y��-��r7GF�H��
�uǮ�K��m�{vwF������q�q�G!w���  N��;���w1�����Sx��ԱQgv[w���n��C���۽�DVk�\⪜�Y�o������`�9�+��}d�TN<���aPp�����s�~5&�����3��m�{��{V%*�ocI��ң�T�Oq6��}q�9����L��d�A�拭�8���:8e�þ�]@2�z;�{�'�t�58���*g�Uk;��qg<��Z���V�F�<��zua�Cdю�o{��!�Y<$Ո3�m�ʫ�_B�qD�������+�@�1�Qt������l�`a����da��s���T�P��p����	��q�e�Y��B Y9/]���g�Ê�����w��#�A�$a��Ȯ���m�fȨhn=�-��?g���|����h<U�ju	e�w�@��\�R<,����Y��T1��C�i�jEA�3�y���N����`C��lt�$j�� Om�]�"�����~ݗC֫�p՚f� #�g}ݏ��M���F��v�f�/�����u�M���%	\��Hn��3�yn�}���\��ӑ�����7=�i��T��U<���������EcB�^ܖ+��!�"� s%4G-�s�,~�~<�<���<F$�d�s���6l� CKP����*��ԑز8kH^�����ULW���X�c���`x�����"��Mhco��c��6���`]���]���F�H�j�p��︮�H��Ù�~k@� �R#H�@�ig�Ĥ-9B#��wPx��:�6ES��e�@j�� @�ވ��݊gغkVV��Bl�nƋ��7_�x�U�	~�F�[�A�}�z�Ce+��q���F��=	{��E���wn;�Jv���߻ڊ�u�ݛ�;��p�3�!�г�9�Y�b	�&��ɯx��W�X1$�
�|D��qoG�� ?K�ѷP�qo��{�g)�]�ɣ<;��H17Mz�x��:_���Ϟ���Z�s�S���w+F%5���b�
:�����E�ń�-�9�97�y��i'�D�Q���B���a2��S�wr��C������x�c/� ����]�>a�Tuć��ۼuN��c.ֳOm$O$��j���hY����ձW�|�����r�^�ۚ�Ӥ�=O'�T3�R��6^���-m�?~}��h��޸��X��z,,��m��#,����V
h3�Hty�-=�s�E�T)Zl�4K������m=��~��H��X��ӕ阤2܍�G����|ď�xz�{k,��Q��,fG��yn�F���</dyix:��z� V+x��]��Ԙ�[�Z�Փ�36�5�c-A�ϷB�dჷ)R��0����xO|�U���<��Ū�-�Y��{���"�Wp�qw�g�p���o���ӮW=1�1���S3u�!���1⤳���e��g�������)�$�Fr��a�� ����6k�Wr�m]c�.<[k�5-��S#8y�����iG���Կ,�Ayo�m�}O?<Q�ͼ�lJ�H���k�R����L����C��k'o7v��c�<ɷ[����� ����t��@G<et�:Etn_�� i�"�#�h�V��D���#n9/���\"� 7��|ގ_Oyi�P�B�ozl 0���CC�4���B���+�s�t�,���6j��7U��Y�Y��4֟B�K����0�	�w��pj��5���Ot���'�{A>3��h��nYB�� �* 2(���,��iȪD��;7|�CݡjsU���*h3CC}�2�-��X����CmP�a�D����u�w`��T0��j���"�\=�%�Nm�!R�㭝ƽ��XE��۞Z ��ڜ����S���a[axn�l]�ͫ��6k���� {� di�!��^�v��������N�IN�ܒQ;�$I�[����!���P�A3��t�"G�Z)�Udp��@j�|��4+���t-�+᪮�MUY�v��󪫶/լ�[�R��hVLР�"�5U�w�,WM
�<:a��qf82����4(Y�dU���}V F�TAMPDf���OӞ7U��P�MB(0�CT;����f�� U��Y��u�/� "��T��d�d���~|gݍJ��Z:Ab�p�:� di��C%��ƚ�4��C�Up�B�UT5Kf�g�ج
�A��tС������ ,�P��hEw��+�Ei��j6� ,ЮVhT"���)�1T8hW��@3A�A�0�3���*�@C($���"�f��T����O���C��Y 	�;�⺪� &��  �U�X_=�b��4 M� 5\"�5@3�*���,�U�
�B�4<u[�\#MUw;ZM�f�>r�Q�����>z�a�Jk"��y�®���)Gvvg>^���s-Lt���s�c2���vDp\�];x<<"�����MUt�@�N�};�����&�]�-t�vp
�B� x���hU�U���_�CMt�  �dT"��@���o�4���rX�4 �hU��j���5U^��Ь#40�'H0�=�5ZY�  M�_Ж���d(C@")��7���}=c������v��^G�Հ���8���y�\����E֋w�W,��ZL� j��E�+����(CR*�f�Y�1����b���B�u
��H�e�"�d��(sU
dV�B�hQ"�� �s��uXh�;�=���n���ph 3U�	 "8EC@{ۦ���R j�2 �?J YEP�k�<�r�i�ZB'��U/]U���Y�,ШY����t �R��y����������T�����@o  �P�2�!�"����`V���*� R,С��`�9~P P� ��{�݈.a����؇�g�ȓ�U�[��:|$�aޓ�'M�$N�
�E��v(p��\ @=B��5f���Uf{����B�f���3���ߞ�PDUx��*޼Ạ��"�yi���������_/��q
j�Q��N�����Ƶu�n�L���� 0�^45A��m�i�|����j��ߺ��"+M�Y$ =���B�����oM��h�*����
�H
�o��5CH� C@��T5I��x��=���f��9��ӤP� ��4��
4 ����t`�E�J�n|�����t�IB���H���8E�M*B��hR"����{w�({y΋�P�͑C�P��T)O{��&��8j�E�쎂 YEo׆�H�5����@a�!� �9�����V����0z3x*�MZ<��|n��&����ŭUz�^�w�+���.K'�xs�\�m=�*��Bщ������8f�|��k�K�����#-�4�9(��C����@%Øz톭�e�wPS�ݵ�<�:���U�QW�d�N.,0��:��ޱp�a���ݡ��z�k��V�M9�<�)<��A��7.��^�m�D�v�VO�u��n]�Z��I�����tؖ*9-�)nѓ3A�n'[�vjh�k��)e�2�ˣ���X���`9	�����J��Bɵs����h�I5?�x6��t�gv��J�$�hnM��؅����t�N��1����P����H��Y�4�@z��`Vj�j�ЦE��]�@���[������C�Ux��[,пy�j��7}�`!ZG�ńP���vC���0Ҍ���q�h�8hw����FT�U\���������{��C� 0��{9��W��!P�G��a�V�D��wT1�EG�ڮ�V��(l��hP�K|x��sEhB!���f�����thk����;ӂ|"II�%:s���*{���P�X�
�hhn��t��o�*�I4f�7����跔�U��\��^���Ь4��0�ƻ�`w~v9�:�EaÆ�mUEE/#�#�f.\���zw�c�'xt�����y��>}0�W9�u]�T  ��.�� ��ٺ�
�Ƞ�
���@R���cH�N*�hR ����SG/�XE/g����+ "4�UV@��h�[16b,�������dS5P� �>��wP�u
���]XQ[����^���z�8�ES47�� Y����q��C��U����G�аh5��׼j�H�fjEU��2(�X,=0�L��_�}}n�i�K�h���<;]�n�(� 7\y��1=��&����m�l/&��p�#�駏�T4,���uXE�3�V*��Ea֚��M }~�t������ �K��}��:�����H�w# <�管�̽v-*DU�Z����L�_Lƪ4�(t���d��oM�F�������a��7ޞB������ᐨ�����̓�R��1��F��W#{�q�0���Gɍ�-�"���,�Js�Ы4 h4��M�E@����5��٠9���M�c����9�C��YD���+�"��^׻�|�}ա��͎�������-5*HH�Ɓ g�j��:j���<� �^�,��a�#�V���<`2 �
����;\��=-���q���^�h�SG�"�^.�Bҫ�w=����H d��&��2��v$�i����@i�DR�w��߽��J�"��A!����U��� K
���=;�;��")�@�j��w�W@\ F��Q��y����,@=}(a����I1 {	)ܟ���6M�Hۆ���MT0�D49e
�9�f��P��l�a�Vnxs����������}�t����4���y`�}�`�u�(C��=����q٢C�MV��S4��T,֚�-�ºE�X�y"���a��2	p@T��K��;<��=CuGoAm��;r<ᎃg�1h��p�]�����@f����c�5B�@�B�#� }��b��l� @�>P�X���T����v��מ׎�3TȤEvs�w��ҍ<�T�@���G�r2�F�l@�Q�#�@�"�j�cJ�!x�_w�,T4�C�i�ɵ�+�;C�E������=���f�І� ���뺢p�DC/�R4x���� b���Dw�Vq	��/��ޱ�45P���k��y`(��qI&Ui���a�Z^#��܎���Y�q	�&���\�WU���1�.f�����+��E�g��Uo��07�
��כ�<g�'z�xK����nL��	�R�����k�l�R-���^�i{qf�uU���2q�����N0��$@g��T4�!�Ek��"������d�Y0�T��da�0�j��G�ݿ6�j�����p���5'��R�dd;
��-ᮮ15dCL�W����5��4�2!�.L�A<=�D.zq���!�&!P���v��C�hi�l#��!B�w]5\+��6j�;=1�#G�h'3Ud /s���s/�,t�$=@8� i<�s�WB�c O!f��&��U\�����x@dR�,�x���t�9z�	�l�njB���� �ݶ:��%�Y�����F.��xWMo R�evM1��,]q���(2 G1P�jw����4dd��K]43�s/����<=4,��")�P��٢h�wn��^�wUHU��T�a$P�{4ئF���Bo!߳�̑��n=�>Ré��)�8�)��)�W��f�l/}��Wa��d48s���� xE29wpV'�+����f�2=���y��Y�+�<CX���:x4�GMX"Os5���R�$�!�� qo{z@�##s��c���f��;��jݵ`B4�ơYw�������H�DR�{����6)$8@DEs�C@>��X�+#NW�zC#��tn-���G#j�p�x�W���z�[��^�����Y�{�99�`p�5D�2�o=�+�|��2�!Ԕ�2�ߍ��.���s 7�w����}d�b���
�$�b{48�U?�މc�dE-�;Nd�T��`�!ezX��EL&���OM�fe`虞^c��L�k�8ＬoS<,��G���CG����'"7�\D�@�Shq�<p�U�6hCz,;�bw'%.
���b����C4�s��cMiF��ň>�s�'Go�SQ��F��AFĞ��U�KI��#X�BL�I�q����ny��3�n��_d"��tg)�Q�5x����[2���O��"w�zէ�����H框����)���^�A�a��p��{t�a�:O</���x8@��E2 J�{{�]5���[�����)?�Lˇ#����|$���dT,}\�f������η~���Y����'Z�)>H	�;��������kᅄ �>λ�(�6��s�%shq�z��`�q#
nE"�����Y�A���Ω����Z�f�+�VH��p��������7��B9Ŋ=�+5�P��s���3�j�����I�,�LtTA��ɤ$�h!O'2u����xD"��uحH��h��+���ł��g�Vj�}jq�z*���g�;����=��4����ı@}@S�TSǩrd�Pe��))P�Q��%�H�f���`YK5��@g�i��4��{����A���4k���z_��H���tO���]���J˄!{��u4mk��Z�f��us(9�����GAA��ύ����^8����r&.��0n;ڻU�Q���7)V�liЛA�KAA��ktn�i��R���'h�%e���4X&C��U�r��B`4uyKY\�u6�tIfu�º�.V"�eຊۻA�)e��[`�R:������4����13�R�3�2Y��l0Xt\��.k�u��ǐ��F�ptmWm&��Y��<�:��;	�H%�ֺ6p��˞ڻL��͕ڸ�{C�]����4YYH-��e��
��������uڎ{.-ؕ�'b�b΋�W���dlɈH����v���n\۝�v��L�+�{�@�I�KK�}����^5�B�:��z,h�3����#{�}y�%��[6�����!��b�a�֪$Z]yY�rF>I~D�
Y� �/$v��q��Z����+�ٵ��J�=�F���|��Y���۱��r�"�K�wA��~���5b��?�'Z�h�b�����S���
C凪=��A���لV$�U�n��	�:��]
�)�̒�F��yX��N! ���le{��V�޺�<n�	\�����S��
�)iT�`"�����`jbG�C4�a�<��戓Թ7��$i�PRxʄC���{�L�K,���������Bf�� ���dY�O��7���@2;���)���L�de^8رb��c�gs^�a�������kэ�v��)�򦊪�q�L`l�o�U\�fI��w�C^4l�B��1[s9,�Uϙ�^@"�n���+��Te�$f+�t��6�%և�	�wl�u� ���!m���nt���Ǽ���V8	�bh�E�j����}]����Ub�\[�t�7ޞ�\}pxr"�����BG3y�;Ѐ�N�2/k�����DBGi�	r5�x�j A���9Z�fsZ'��\��vP4�����"��.~w�7�q>��d>�z�Z�	�G��mA�|#�&�T�ٲ��u�k�7�V~��8�U�4"��U��)"ާN�噽~�V���K�<�C�$����g�x{��-�Q��M�xGp*�Я���Vɯz���]�w�Y�~�>ʓ�D�Ȼ�Ε�n�+���L(~g2����m����p �����!,8���eɴ�*wx����o�/T��q���Ͼ��A�n�4�fA��]@���M�R^�r�^&��t>IZ@�B��|��጗.�����$+4�N�����ʲ�i��Y}�w��VK�)z��-5LTN��l���) �����9Iؾ��5 �d���l�8�_p>l�,�I
@&H@6�w4k��g6�&�Bh���U���-��̈�ԃ���������,��˂gw�:k1D*K�y*��F�h�(Y�sx�h�zǇX}0A<�B� ̀|-Ws�� ��9v�:=	m8���K�{°i�ub�Fi���d^�gWt��WPd�Z.���6��EF�+6��.:*��U��^��Ko�@YLq�޺{V�q�C9x:�Xj&�0@T-�V�k�2�������}^���S�����}��5��JxG7ފ�Y�����1Y�^4���4������n��]��0h
>�P��e=��Z}�Ir�C���/���nߙ\d�8���X���n\����>@�B��!$���P����d���.ݳ����X�B�4���3������ѽ�Y]�[ ^)�G��f�&��س1蝎���¥y��0Ɯ0�g1g��{���<�������12/�Ok�V��-��J�B$!D |����Z��)�_���|}�Ά�Fuy��$��|��3���XZ�g�ϭMѸ�X��{]�v�O;�	�uc�\�+Y���9�*�ym���y�צe�xO�W�G�ڊ~�s�J���Q�ca��ۻ�,_gen`F���s�qy��dPn�	�H��e�ؿ�_@st�z-���t�j�R(e�9{����n�o���=;������H�u�V�#O�c������_���^N���L6�M�x9pT�[:�wL�� ��ޕ�gR��sO�����GG]w�3�߼�!��v7IS9�2fq����:c�DaA�$-���6����[��m5�g+���JKlwfVW��|`�Τ�e-�msy�Ֆ����w
51�f:�I��ZpG��ܧ�'��<q�Y��ӧ;s�Yh��h"S�!lfP S1y\����w��,b��U5�4{ۆ�7�Nz�/��H�}�
�N�ﺶv��6 M��{�Be +b�J�R�'�l�53���~�!�{�%$�>����Y|���qd1сwR�YJ�2ũ}jJ^T����Y��CQ�w���=p��1��luϱJʸT��(���Qn�,����Xi���g�Q첩��W�X&�Eq���0P��7��<Z��=	�ս Xom��^�g�Ё�	�$�h(���ôű}�·�:�^�f��o����]<�w�.Y�hPk���y�+�G����^��f�"����!��`!Q�2�Wz�4%xّ���!^��X{3>�p8����f{��i!����b��#J	��A%�e�R iI7)���Mׇ�����݇�ݷ�&[ڗWsֵEn�R����<�ho���K�$HB�p���X��[���4�a�>|n�[�A�P�95S�V�$��)��m������UW�� ��U�T ��UW� UT*�  ��U�� UU
��( *��Up UB��� UB������UW�  ��U� UB��� 
��UW� UB�� 
��UJ� UU
��� *��U4 UB��z 
��U_� UP�����UW� UP��� ��U��(+$�k!nƯ���k0
 ��d��G�}>�+E @
��kF�Q��HP(V���@�T���WF��@Jk@(*�m�    �i��f�A!_        :                           � 7�      l = _<���ܢ�圴hF�	p ��[�zz��[/;��m�7.Wi�l����)Q8 ��nsGUm��v]��PT =���_t���[st��H� 륖,�䣥+9۵�����&˛����� �:���m���h����N���y�zU�%P$��)�      �  {ޱ[mg;��W���T�9�s*�vd�����yÈN�-�n�ڭ�l�s��jRtYE�� 7X�m7sb� ݘ"��T/YU�q�ulj�\�+�E�� w{j�[y����fk^v�mlĢ��<�bv�V���5k6��8 �]нfچ��Y�o3��h�p�ǲH-c��śl�!E ��         �=��t�&R%{s:��=������Zk��n׮�Ej �6޵�n��ض)�1U:Ү1ܬ�!��6�a�x z)׮�y��SY���s�m�������s��Jֱ[� �u�6����dي��2�٥��E���[kL8 4):�w.e�ѹn�U�ֵɻd�iV�5�i60R���P�n  z      �SK�<�\5�V�]vbDG;�JM��vh�p =΀���N橭gE� [���6�7;�N��� �m�i��TWZNv�i  V�)lý� �'�t�-� w*��N�+l���ZE&��n�m��l��v�[0� x���G�ސ{m�7����-��l�T6q�R�b((��         C�x(�t��`H/=�G���-�w�  �M����н�ǀ ��h {���Q@ y y/m�7b�:��A6(�t�=< e�@QA��:�e	4���5�e*� Q]�R� 4 ��@�] 4=h7 ��h(/Y�E���` ��`:7�f ��("������ <�����=z�LG���M�@��i�9v=w`�)�$�J� �@S��P�� MRP�T�5O� ��O�*�*   ���R�=M�4 ��MJ��4 2<zY�]�fz��;��p��5�9��c\9�˟>[\9�ݪ����W|�2Tu\�x��P����?���IB�ҡ�P��T!���v��鮺��߿[�0���V㺕�.��4[�^c�f:�cy�/{&,ڿKjG�*LD`��1�!��*�f jy�
ռ����%S�E�c4�f<Ym@f�Z,ł��3Z�uNm��b	�h�Dq$�]����L��16���VH�a�w.�|��-��=�7`�,�jn���M)N^�O�	�h����lȕp/"�R�b��퀲ȥsr����D�#S_�a�T�(����Lkْ���W��]<�jd*�GoY��^4��,�ɥ;êFl*s1�~	��䮣v��[c�(��2��&��yBl�oV���wa�~U�dڵ�0Ǝ-���)�h�7^��\����[�EE��n��{�,�0�Ż�jݽ�Tnٯ
�l]Z&��m����qb��Zb[��sR.d��*ѣ��qJCQmiof�����Mr�^��̽̒��c)@�8ˆ��tkR�^�i2u���n^��f��KW�n�-���2��dv�<1PL�gNRљZ�G��.�{5������&�n�l�3a�ن��V3)�n���3,3a�+jU�`:u�o6h���)R"��nF�Ț��m+a5I�O)��{�`(�ftʎ�D���84�VCYф�j�e�\ZBo� ,kq���L���e�J+�(�m�3���iy{m�hV+�-����4e�1:��f襹�m�ݪ�t�jԬd�I�"��3w@#S��0��ǖ1!*j�v/ՀLt��%��fL��Yy�.<to�]��l����28���JN$��yZ��=�rY͡��]ٚ�l���ѡX�	��75��0��Yn�fhGc�5k�2Y���K�6�t���X��n[xC4��Ndf��]\�e]��q֛Օv��Bmn
,4�#�nk��?���s�A��&�h��M$�l9�Q�����\����Cy��m4F����w�pk�n>���+�ۛZ�:Ŷ�f����=n��vn�۬�K�x�Xk	�J�ӣ+=.+�y~I�As�[�+au�6�E f����+,�%�&��y��h׽P���1b�ڤ��ͭԢ� 'ُØUͶ3�D��&��~i���,�0�`�Thf;x.�k�a�7,jE5�2|�u=���ld)�Ny�
ul4n�X���%i�r�r�A�U`���7HШ��,Ր�/+2j���S����q�ZJ?x���oA��a�2��Sm�&�� ��ɕ�t�[���95�M�.b�oP��v�W���zY��o
�+�]�M���!�;����Wx�.e�_���-���B6Ӷ��՛��9@�㺻 *ifXݬ�R�m)�,ܭ#Tb��,܇4�1��D�r�bj�Mc���I�7�ۋ�Z�Y�&-R��Ò�n�nՎ�G��DWu�R�Xd��tZ0й��e��M4Fԧ$;Re뫗v��,������Csp=JƄG��0��=w���{$��jc8iD����kU-������"y����e\�m�N���4����Ƞ{���2U����ͻ����敘A�yb\��.涱��f�J�����
�8�AZ&n�e��X��t���,��fsJ:k�Ȫ�f�%��f�rި'�N���}���6K^)�xf�7S0S�f�ĵh�x!6�\v���M����nL:�n�őZ�Alb�V&A�d���,\�&*�ʬ�:r�ʹy�;řu��VS��(q�Q�.�u~�%]л�aE�Ga�)i:W.��sJ �RY�A^��Y�B2��	5�� SuH���Jyjy���~E�CS3=�f]4���ӗ�5�x���oj�u�4h�6���Q�3�YڅT�JY��5��nY�laȶ�1��֋�5�\���i�1V'ӂA`b��%T5m�j�w��ûn��ȫ��:�2���$���w)]ڒ�6Z��s
 S�� ��j`tr8VVB}y-��"�X8S�����@�5pbx�
ȯ�2ݥI�MZ���f��5�*�937jmM�0U����=EZ��^�z����3p�p��yB�y6�{��b4�X���cGq7Wt]�mEW�d��ԫ���p,�MT~���*�Q�-
W]��4t�S-��
Nٔ3�i�ݫ�*q�c�v�S;H���� ���;�踲�"*V�l�ѺUgCW&�VPW��4ڸ�Ё�T @ɽ��V�#��Lx�af5��b���oD�m�nL�2�Fk(T�ܷ�Y���#E��]�5�۽��cm��^�ޫ����9
�v��;yV��EZ��cim�ʛ��a��d�u*-b�V�աg�Tq�
��x�[�pYtq�lQu,.��`�yW��v��L��X%�O1`7��9�#��ٙ���.��0N/{�8}L}�*�2L���t3k6�ӥ�n�͊��%\9��H����!��jMM�Ž:[^��[�R��;U�vI�dn�x~����j�=�b���f�n�Kŗ�=8�qT��>�MKM̷xVa�1���P˸��Պe��v嬹4�nAVCچc��a5��jX����.o+����~DF|�iN��ԫqZ���Yw�q̛��-۩Cj�� cqr���T:�6bVn�p͵i����O[,��(]Y�f1l�]]���YJ��U�c2��r�0R]eiӴ�c�6�3rf��O�����8a�ft�x*�n�QIF|⫤1�AXVչ#ͺ���{�Y�J�{Yf�q+��cu��Xᚫ(m8�c&Kb��V��%v�RG.��Yw{�����1�2�,�29P�柌���D�q؅�J5{���K6S"����%n�d-��l�ZrY�����cF��`W�]�2�O2q�hXМ�N����e�fP�qdn,����ɨ���$�:D���W �$���S(p��
\F"�V�M#9jy')���'9Uv�TH�T�5Vr�&"7]��jN&�3,�2֗3kNw\�]c�U�z��Vc ����1m<�S�n$�K�{6��/VL7��H���Qiqf���V�l}��[���LT�w�ެ?
[��G�^TϷ�3�s@�r+��XթfSIj�����S&j�#{���Y6�j*(�kZg-Լ��*��s|-�jh�)�^�JZ>������tP�n�੭����^s rF��K�.*9V$�	���1�?<��.�ט��sfi�B���'2ފ��])�g	u<j:���U�t��������nd&c��,7����f'����J�Y�����l\�ve�t�ؚ�<c2cm?;ē�)��k�v�.�����V /pWZ\�"&�t��3-
oh��d�qx�ױ��Z�X��F�$���(�	��:��Q:YbPR�~yㅠk��w�-�$���5'v"u�rK �Y4J
���!�W3��UzɈ6fnDe���b�u�^�Y��,���Sup@K�odU���%���7A!��r�v�!z����{S��Uh�#C,��{��(�x�&����W�%]?{!��e)��RP�l�d�d?%yA3WO-��<���f�,P�2y�=D�f���s\ջ�$��7e�մU��Uڀ؎����z��V��۝>ݺ�{�q»31�~��M�{���B��d���;�1�j��U�tb���q�Z�r��җ��[�*�vyWT �rx��
*
��6L[4�7�ˣv��R�MLT����Z��3c�>F��?H��)����c�h�4Z��3ѱ&hSw�0�
���L��g���(�he^����؅8-m�8M�5Re�E�ac�Q�O՗�1سb��QR��
�K,��Y���Wx��D!&��#��a�(g��Z��IF%խ	�̆��;��P��DciO�YoEb�w���AUʸ��T���Ĥͫ�l��6I���Oj��:���FԊ}*�������(kY�wP��ʏ0U��`��[��5Ѧ�n��<�����-n���.�=��R���]����Aj�;��`���p���q�T7Kmk�J�"jDcŭ�V����|mh7�R̒桦���pO	�5`��E�bT�M�Abt�ˬ�`�l��xU+WT㛐%"�Sz�-l5��n�cVwi�X�BPܡB��Y��ۭO�*T�V*���&7r2�<��h
9��ˡx#��G2�7%.� Ԕ.Xѓ~�Z�)�y�,�<ǯ�Xݘ��ђ�%*�Ћ��[f�`��ّәJ�uM��7���t&&�T��FJ��l��ϲV�y����
��&/������a�e�-,�w�
�rԭ7��8]L�SY��:��H�E��L��X����V}V���H�xA�.����N��oгuk6��@ X��T�� {q�ٻsh�GZ�a��IFϝĲ��̖m����!�1)��YZp�AzČe�>�*��i6T�Bf�r�����lC����o!�f&!�����2'�z��Ŝ�'�T֮l�L�1�٠�?
�U�`�t�'jV"�VXx�>�ʐv�E�K@�p�7%��yIlóe�ظ´�V���]6n��r�]�J\�,ˡ�L���	��"Mgى�AG�t�i���F��jVqk��J�if�Uȣ�k5f�����h�Ah&�w/-h��.����ajPf�q�g2L���o1�MQ�Y��Lߎ]��f*OK��,^�IжD.S!�ڑP�N^I�b�b�k��6h*7m��c�R�Դ���XڃN
��+v�&bǐ�rQ�fe������& q�+~v��y����mح����7m�SFz��m�@�8���w6���y�����$���1�CX�ta�S~~��ٖ)�4�S�5	�͢��@����67�&�ճr�Goaֽ�YD�)o�S�	�w�Gԓ�a�`U��Kpe�Y���[�&B٢�e �!��3;s�ۓ>@���]2S}�`:(�����D�Z�ˑ����A)YE!6��d��=�8�n�V��"
�
&�ё0r
�*5m=�z�a��x��p=*f[obM\������w|�2�$�O����JsT�k�8[^R��/T�q6H�u��Y�q�[6k��@�D%��#�h�m	=W����f>��W[��)%�I��X�nV�I�5�|�0P�`�A�1��Qm��n*�����{�s5vF����V�ڋ�Nb�"�P-|�[�ۤ�^��7��kp�#A/2��:�.-YES9�X0m'ZU��u�GS�3h)Z�]4��bԁ"R1]G���&������V��y����d2ɽ���j���6Ju�a@�m��3*J��n`�u�n�n:oJ۫-#%�cvP�P�JCe��0<6[����6B<a]��n��Ѻ-�����)�>�(�H-��F͒��oj�ݓ$�i����Y�f�4N^�������3d�����eƅѿ����b�-�6�%�O��@n٩i�E��.��,�� ���u��`�Z�H4Yw�G�dۺDf�����M[�����*��i�X��9�U�ݒ��#6�NJ�fcGV�u�G���CV��p�ϕT��u5���#�a,��
9F��&*�eԗ�vC��n�D(���n,�W��e�W��k%mۓ@Xsf�7T�V�Cv���X�i%۴����[AF�n���$�U�dA��P,�晻sq^ЃF�3"�*A�{7*okNغmݍ.�1�����-%Mm�y��Y{vqmmgr�4㩚D4 m�6%b��5XٷW�]9Fcl25�)]պV̷1!c*M�shp���\�0`���y6޻�
e
@Jf�)�{"�"h:��ַe�wf(�3*�m?�B7nE�e�.�PM^nnb�a8N �Ru���-ɲȸ���ٹN�x*� � �Y�XpZ�O�biӱ�$*�q��2��e�׏N^SU,�J��� !�{6j��ΝƩ�r���6mg��P2��r�iLN��r�Pٺp
i�����V�.�`��weL�pr���ES��3A흢u��7�+��\�{�J!�fe쫵���ۺٛ�KAH�M��fU�}1����v ��^����b�q��Y�;J5ʶ�#a80P�5x0v�R_�k7Vsj��l���L�L�{��l�xf��V�����kQ\[�.�16D(w��׋AW^p�&��Hc�%ad��潩S!R^ݻ����7����m�N��f�X!�w�l�<xd��1�[ǘp���Cw
�n*�Yp&1�H�����S �y���r��9�=.f�j�C�i����bnf��[��uJ�Q$�l"�ms55{�1���WyZ P�s-�he�[	�J`�K`I� �e�C9��I\��V҅���(PU^�y�p-�&�t�37f�b�qM�n��������]�����
��X�W��{2�2�6�E^�4*�G�F�z�\Unn٘(V���i
*�\��ӌɕ�ӌ��̛n�F�K���w/��E���][m�Oyu&������m�[X��X�ٷ�F��WE#��{��z��C FVd:&������`�j��nH��n�,X�,DwQtҲ��BY{DSt~��%�������,����,R��ZKKbN�gC���{��j=S�aG/43��P�i�1P*�����Oٍ�TX(�Qe�O���,���'6���
�{,�&L"�������ZSXҞ-�e�Ț<'U�P�39�[��l�Xq?����ڶ��h��6�Xxc�O+#N���
��r�.�[t�Z �O�0�$+�鵂�U�'���|8�+���U��EJ����v@̰^g��[����֖L���,�3ub���X�"B!���+�e�g0͵#�e��.��¶�ڀ}j��Y@�dY@3�Ң����fL�߳HU���'L&1�0LUn�V�U�cB�.];��b4��XuJ{2P��R�WDV�Bն����M�ͭOb����׵9gO]�w�:up�2n�����F��Z���(���7cv˕Z6�x��:���473r6���6kr�s���n��Wn�b�8�ܯI<ю�,]����F���2�Y�nMx'��%���uAs�5�6x��Q�n8��!�6�]t��]����<G�fu�}�rR\��Z:n��w;Ge;mvݸ˹��7>\e����;��۔y8s�{[�r��O]y��[l��b�]S=��ރ����:�d"N{�2���WE��/i�'p��g�q�q�B#Ɩ�۝5�F,�Gc�n�Vz���r>-���ٻp_v]�d��)x{M�n;�͎֣�9�"���k��vv]qΐ���n�ގ�[��f�	�ma���w��N�M�[p�p�Zq��ݶs�;wiI�۰�Υ�n�\q�nO޼��.���J��v4nl�߇q}���WZ]ێ���lr�>�2V�5�{l��k�8ymۅ������ы��5�����}�"tz�-�u�n1=�HC���ٗ!QU��'j�];���lr� ki�&G;4v�2ѹJ�;.N�gî8�?{�"�m���}zcp�X�lK�nl����ㇳ�n���a'��b7
�[.�n�ݞ1�3�:�M֎��Ϸ���P�Ic��Ө��M:�#&�6޼O���]��%��mt�a�8���xl���zv�L���l�s�7NR�������	�grnA㮯:�^��#�+�b9���+6�O��^���[��מ���m�x�އ>z�&.8{zxu�p/S5j�n����8�\�n��^��pcy����:I�d���j��t7��iS;'$��(�1�5�Xqu۶w���/v�;
�#9{$s����]F�EA��ӂNz�����혧�]Z��k���0k=���yNs�O+����nq��4��o���[�n{ά��D�')��t9si��wV��n'l��
���j2]\r��s�݄�`�������7N�]H;���%k�زt=�c��:�Ӹ�+�&*n�3=���B��W8Z�ۀպǋQ�oCn��]�C{1ۮv�4s�pk:5/E�n�j� unuƮ�JES`"�T��T���UM�=n�l��6n�e����f��]�����=��=���u&�{�g�6��=�q�75�sؼgEn���gi�n;dMg��Ƀ�g�:�>L$�-���\�8x��%�I�C���p�}�ێ3�ck�k��A�xN��'�Ť�\`�����rn4�ys�cf;!��1:l	W�i\UWO]��3�ٱ�`�v��:CvZ�ʓ��n��{nݞ ��3v�	��gv��� +p��[\���ո8����J���ǧv���v�ݧ\�m�b{M����.ۈmջXm��t�:yېN�mG4���h���;�,�	��p��kc�
3�ۣ=v�3oGTv����t�kd�'�Ǵ�r9C1��T�<pOD��x��]����L��x�'�^��k.��t6��q���Om��u˼6s�u6�-�������Yހ�tvj� /D��6���q�H���yܧ-�##1���ǡ{V5���hv��d��y�N.��Quv5;oG�~;c��?r�l�p𗞷FǇ��X�^ߍ�;��qۆ�%0g�.���E�(䇝��, ��l��n�W	�m��˭;��.+��;�D<:��d��r�LX'�8��%�gu���'���s���;�3@44T6�\ay���v�^�����۵�8"sk��n;M�a�g�on��T&��q�u=I�*��7���9�km�y6���YP.�8y�og.�P�VNM�v:���Y��$�N�q�pZ�0�E��5��:N|�&�w�C�u!RqYL�&nnԚP�o.����o<o:l\g�]m������!�-mulu���rX��i�v;Dg��7W'�;\N�ѻz�9�h���s8\vr��g�$�8v�Û#c%m�[���B�=��o)yدP�78���e��0�t��ֳ�[ngL��q��<��s� �pt�^׬��a,���q��u�SH6�C��y�go:�Եnv�qĮ��GR�۰x��z=z��7m��ݵ�<���mn;���Pq����Y��k�8{�7m����iX�n0s��m���d9��#`vv�,��H�ں]�E��,��0�cm�[�4�NT��1�ۉ^6��X^v�<�5nvWv�mp�*�v��)v�0?���{훦���Gr�`87[��g��O�ƀ�l[���8@��u]c�����v��7�9��l�T�ޫ�LD�(:3�<p�۷<�g8	�<�I�^�W5&��c�1��l�ݻ��t��m�OFq���[�;[5R	'hۢ��:;i֮�؈��l�홳��Y��[P��܆�a���X�]��#��nM�<����v��)��lcx]��Ǘ�5az1lRZ�zC��:�l�yw"��L����#�dbK]�k7E�\cq�W	\�m螠��vN��&��1�^7;��0!FۜsGc�N3����kn:��]>�38ݎ�"ۯ���w�]��e�ȹ�O-����oU֮��ɻ��񓭹���U��c��nN���mz�����`;������Fݻ\u��@��I˳�����{{{��u��q���O^1�����pv�\n<9�:�8��	݊��@�n�MZ��{s[t��\<�,���(c�{p
:Ƞ]�q�Ύ���c���ކ��Χ�ӵ��*�l7o]t9��=�:ݮ�)�F;sN�ɃQjsڱ���(y����]�qǊ��_�N�--a�+ e������nKϱ�qsg��rA�sbIX��gs��Flv���tm��
��z��oQ�O�3����/�g<'K�F��q��d���s�K]��.N�	�xOZxn'�w�'��q��'i���\�K��9����H��	�+5�����j��Ȉu������lO��wIs�9�bP-��v�y���&����r�=�
��[�s�y�Gуskvd���k�s�)�3�n��)�wgv�s����n��n.�j30<X�WH�3��wMɎ�xK//.�u��*F�s��T�m*7�y�G�=��t�����Y㭝�\9;j�!���tBd4�z��XkFtN�X�so�hx_|m����ܹ7�^�3�됭UѓG[qrmۯ���E��-x<�렚!�S�ڀ�dhf�%罇��Z��n����=�m�w$�<�����Tݰ�_�0�� ͎��6��wFp��u=)�nv���3���.�3������ū�F�����.�c�N���p�;���G����]�x^��/c�ٵ@J�-Rb�rv�J��5�WQ�8��ηf�OѨ��;ćʘr�Ons��q�ݗ�&�yZɗ�ȝq��]���F��kv5<��3�cZ�K!X��A�d�s����jH��
����v{�q5�=�!�+v6�H�u�I��E��\�듶��s�1�n:@�i����z��}�_pYϞ�Sex1��Ʌ:�D�=���B�ƨ!e�����m�y�w7�6KQ�[u�k=�z!ݕG�L�b���9�]L�\tok�ݶ��ɴh��ځ;qn�f�n��Ye͍�<�A<F����k�:'��N�ݻvg������̕�n�����]��k��=��{
v㭍��ݒ۝�+�=�K�k�{[�|������g2b6�rbM<�Ӽj��rm���s���cEq�5����m����r<z��mu�m/��N[��k[q����&��lF�\�{�Nv���b3��#�vۧ��>J4`���͈���۞���Gbު�'�S=��srlCџ6�:
�2Y��1�uarHA�5��G1ŋ�"m���=F�v��m+�b@Sq�L�#�bkPu�l�U�(�����l:Ŏv��y[��
v�x�9���c���3�#�6��B�F�\<a���u`�c��wg�<S������'r=��Cr�#n��:rE��m�eVq-a�h<�qn�ᵬ[[Żu�D1v�c#���AM����g����2:�{pq=�������+�878ln����ė=��p����v�v��r����r��٣&]<��N��M�8��7���g��[o�X���P�Et�L�=v�����[�Ƴ��z���Uu�>]퓴Jٷ@8z�x7W%��Mlu�ZMd�l<�{7g΂�;n��xv1�앨�bM�*�>"8��H]Au�<I˼X�9�%=ɹ��_?3}�w��`ۧq��c�����VN=q
��bWsF�=Y�k��g�l�p���x���Z۳����q�|���㎸c��rv��{�ut�i�9�ěn��nۛ{y�I"��n�]u��=��+��;�z�f�C�<��0]�:�>u��.��[���n6n3pڹ��Ի�7%99^�5���un�w�ʍ���+ʜ#�8��@W9����ڔŃ�_s����v��n��9��9Xyv���v7����m���XEM�����p1��|Y#�^����tb��!���;ny'�E�Z��炮��M��=��!�;�n���M���gnݶσ3�A�uRiǂ���Z�o9x��)vvy�J�g�N݋s��u����M�ݎ-��-�l���t�:R��������r�u<�>f�<!������߃�'cip<�=�_V�1�x	�0�(���y�xc=[;�nn���
��t3�q�1y���/!ᶶ�v�p;��2�S,�+k�Ns�� ��+��w�B�a���
�C��$����֕UMV�n���q1:�e���]C��v����r���]v7��Z�ϣ[��n��4���>4�TNR��[��GoV� ���Rvx���g] t��Pvyw����N�=S���v���;���ʹ��lr&�
���d6f�`L=O��t��k�q�$�0�uj�{v�.jo3�ی<1ŵ�8�Z:y���vM�[2����m���q�7��;t\�/4�eK���T���L?�J%
���⨇��CZ�s8�ݭ/�)���Rp� m��_cA�{K���9N���Ɂ�8�wF�V�-��/�����a�N^��H�r�݈;v륍��tqq���۠�>qs��q�Q
��6q
v�^9<����mG0g�����;	Dr2c��������X۰�����nw]�M�l�{iù��Q�Q�x�Iu$���[vz��@^:���붉1`����� K��6竄kr����ڻ=�B۠�cG�o>�[�g0gv�;mn�v:'yؕ�q�ޖ�ol%r��:�͙##��n�v;Tƕ���rf:�ԯXՔ�A�.��ⳞqgdD}�a��hy�w��hצ�m�����8��F�����g�:5���nx�ힹ���B@�m�����<�܂:�G]���A�I���Wf瘢K�4NŲ��h_A��5�ݱ�K�VP���*�ɞ�Q��3��v��S���Δ��kp�yy���Ž��*b�ˤ�U@��9�m�]ԧn�nö��r���W[r�� �T
D�m�ҕ2�g��[3չ���v燂�.趬nfڷ!�/VE��ݓ��\L��F���{;��>CFs���vk����{Q�Һ0�F�ɜVn)��8�7]m6���\E�r'�:��z�-��B�;s�tB>�l]���k��ڛ�؉�a\F\�j�sbMwn:����5���v��q�Dmp��6|=)��]k�Y��G[���z���.����;vv˻���q�)��g-���k���(�����ݑ����u�޺�J�ά�F��y�v�ݮ�#�6��';��-�-<=uf:�;7<���������V<�d�2����K���rI��Ja`�����m�sg��j��g;dc-ֽ��\z�`�,����ُ/P嚍�\И�^�*��m��#�ܱ/;�۲j�UtQs�����d�Ü�l�{p�ˀ�,��:�6�^����t'3lg*O0�<K��}���eHT̈��%�3 L�Fe�f
3b�P�(�I+���]��HH���b�w<�6;qy���s�@�vY�c���x�鉭�x��p�N��n�;<>��q��k�:�kpZ욹���n6��[��8�oNB㧋����ӎo=��"3�n�^������S�����n=r�^m�0p�k �Ŏ�rr1�G���@�k�=&�vzU���v�wbgzܶ�6{g	<���NA�s��p�:���wYҼ��78y�ۅ6˓���{(�0�Og�&���)��S2Ե ���%���i��p��sᙓ��A*��b��U�`�	H���Iʹ�*8:·w_9dh��4�I��9��Y]�)4L����E;m��4�.i5I�&X�\+"E"XP��3H�蝹ZL�'��we��z����V��P`���y6���-(�
��}U$}�g.k�!��%��4�<��xt��g�y�ݞqc�ʉ� �#��6x�6��Ks34�QtN�m�!d�R({��!/���Aa�\�LV�q.t�bS�kO�sT�D��Q�j�±D��4������X�!vjdJ�B���+�T�]S�D�M"n0Rg-�F�g+�s�r\ sϲ�`�Y##J!P�G������0��RB�D��gH�a)8�P&j��{�UWNe�P��ͪ�,�6�(�\�?	wZ����Knqnv���n(��P�R`�T%���tؘ�O�Y&�Uv~�)n�{{S�\���ϫ�1�3�&z���
������u7�&��S��k������Tdb�zo��7�g�'��d��'n�ɧ�F�#�+��\>��ã�m��h�C��މh����m�ǃ��l����O*d�x��{/�9HQn}�,�+�.�u�d��Kz���V��e�����G^�5ۉ� ��6FuZ�J�5��:bS.<y���ߣ��Ŭ��t��W��^�����4�t�C��t��& `��W�u=�Á'lːPF�t���)*�d��ו,�z38ލ�T:t�dN�Q_�mQk(�dUQT�tL�ݞW-�'uv�蝶��VUo;4Ѩc��T+D��WV;�I���GEN�=������l� p�*��j�����wo.�s��r�苼��tB��KM�]�ԀѮJ�]���2�J��ݔu�wCf��
ʦ�H��E��X�Vз�~���P��s;A�)���*9�bKjB�}��M��}A-���z�ٕ�,�|�H���9�ݽ��qWr�`FU���t�85��y9�8^���lch燬�3�v)�t�STR�KG"�U�r��^k��Z�Q�`��ޔ��P�o��Ż�mݦsҽ: 5sE�Q���ҿ�3B�-P�L�C�Ⱥ|��)�un����������q��m��"ײ
�i��?ek��Ets�Q�֐J���H|��0n���F�aI�;�{�ǹ us_�]��kڝxU�fls�<)�ԧ�5�p�;���ʏ��-ڶ�}ӎݓy�طՋI�����=����E����5%^�X�ʍD�ܮ]����ܠ�Ky�R������u"�H���6��[rm�� �^���xݱI���&�nJ���tF�te�	f
qە�L}2�,�+�>7�V���m"�l"V�?Z���ӡIjV`�v�RΔʏ[ܩ`��[�;���hF ��k1�B�:[͜��Wqq��P+m�49fA�۶r�$l�N�Ksq�ӹ����Ж�mn�VJ���	V�Ky�o,�-�[�¡����^	y
Z��_3���Eګ���
������j�w�]ZQ褝%�I']�����s��e�dc�T���1�R�^��Fn,�7z�GR�9ɬ@G(��s�>}�%���܊�ڪ�d���N�p��r����w[��T�m��ʴ҇ ǔ��4�v�\�����V+��(�����V�d��Uq�i!��;�����O������"�K�kO-x��eo{���t5�[�xٱ֮۫�Υ��1ڞ]6���mʲ���σT��Hԣ}{����wK�'���k%n�ٝ�eAj�S�p�	�@JL�ؚ��:��Ҧ�7Pxs镹�]���W�R<�o������y��<n��hiע�o��SQ��M�&7��zU�cq�c��Q��~�nn�,X���n�m�çN6u�f�J�vf�Wl�`�M�r:�p�Z��v�J�rwfCy~�9j�O�MM8��{yZ�n&�mv<���V9l�fsJ��qDpem�g��p��i
�e8�fjĖ6��B�Ul�}�ז��qܾ)����e�*��J���WwY�TY5��&p�0+����?x��yZ�5�6ﲐ�Ϳ>#��1%�'+��h�ķ��Z���f��&��Iw�7n�8������^���r{:�D[���/e���YS*��	60���f_���1�n�v��d�4�, �Jt�w��;�]��mϼ+�Td�aᛡEv�ˮt����N���M_��2���YܩL2+ܾ�Hk���[���)0�DY�])9X�='a��"ͳ�3ŷ��=�{:.�Y��2L[��37���!fތ�/.g��ot*�4��H<�g]��Żnw6����y�8s�v��W����5.yNy�ag[���s���c�	Pz91�9�PݷV��>�q8Y�ڭ8mvӼ�έ��۸�qɀ9S�V�p�{�m����w�E��3��`��c��ݺ�q'M�k�m�n�1ɮI7gk��������#���/��}&+����OWps�$ï7;�u��y��%8���y�����;n��
mkv`����&��t�έ�e:�f<�>�u˄fo�����{��1�_�Z���+���14'u�~	����G9Hج�f��9^�m���v%ػje��$�4D���c	����m�X�Wu}���v�t�d�.��z�N�|&����t�Q�C��F�Рl�
�N�	��}��ki����ڛ�5017
��Mh���
>��wk�&�B�֪���e"�[h�EX�j4���z�Rs98��c�Ps�fUEWsBWt����=�e|�+���oد'���'ee.���t�,��Y3��s�H!o$�����g���n]ʳ�1�z^�x��@�]ִeӘʾܭ�դI.%&�9��4���NG#�R�qO����\k�&�v�����s1�wi�+Q��ӻR�Tv��1F�-���֩�Ȃp�\��t˧[k�r�f�14����P��+Ɯrԭ�O��$��RIC�T`��c}ޢ�Ѧ�1iM��<��ۭ�ltvĖ#�>������m^?c�C�f�:�{I�H��n�8]q�c�ln]=��3z�x ��,�bh<�`�+%���p� �W�]ׄ����� ў�ƥ���W��i�[):�H�P����=�˳R��py�H�WWn7S6X"]��&�6{��ۯ�lX;����1]�k����C��>���g&b���;�]�\���� r��YwM���Umܢ�M�]ܯ�k\��R5ie:��%����fVgZW�X�p�!b�n���#���\�����˜�2�oO4�^dS]�ZK6�;�$�{�j`�)r
�5�K�s�S��ow{��l�>ϝ�B�����j%�[�՞;#�n݃ٗ�Lt7o]�l���=t�y��M�3H��M��[;����Aۭs�@$w�~�!5�fg�������j�TA%����Zݯ[n��	
�-�&�*)�$�uＮ��y�v9�qep��o��<�hus�b �ީ��������Ԣ~�EǞ�z�ۅM{Ͻ���4	�Ձ!c����-���oX�Z��;�':}�b��p�I��o�Y�a�Djzfn�ă�����6;���O�jT��O|��+x��'��[$�ޕ�g�s�_X�� �2�Gq��*]^��/�k��F�M����J�/��[��Mɨ�sA_��*@��V��s	:La�b����w�K8�n㩢�<86[�(n�����	}����۱�����A8\��F(�mV��W�t~L*t��o�{ʒK�e�n	&�<:���_�^��J�c�θk�{vN^���3�,��JՎ
�]�Ҙ��L>��q���h�ª�D�v��~!3�T˫]�v-�3���o����v��g)��\vK�ݮ�*p�T�5=���~����ڷ2��zؗ�y��z��;�����{�Ӧ�Ὂ�C]��W}��u(]Cα�����{�Z�������J��$E�;K�GE�{m��˕���]"P�X{Y�n벳�H��;���s;�t��|��ߪ#��T	UUzU�e?rn�E��xʧ�i�xlo��Y(Z��r���/�C��w�L ������n�h�W%��n��b��B��U��I+�ۻ�)���" 2N��C;ٕ�s�$}w�th�yG�E)?
{���\�7bl�wX�:uJ��|9cF��>�Iћ��#N�83y�L�N���`����*�G�|JDm��%�b�I�h�Փ���h�y/C�ĳɛ�e$R�mO��5����ؗ}��Y��htGMl1�
=p,�I���w` ��wK�U���b	 �=�t2�����n6y�uAM!�x}6㎝\=��4�]t���C��.f��q[]sr��Uq�[��J��T���k�5!��ͷK�R&�؈X�̡JҶ9���-��;��c��h�CŊ��ݪ�wK���X�W����M�:��L,=����)˻4��)�������jn�vIղz�qx�@��賺�/�4_�U6�t��q�޻
�$�w{��I�4A����Zo#M��*ĥ��:?an�!;�.� �j�Ҵ�����X�rk��=[o�M���;L�j���ۺHf���()���+�{��S+��Vo���71��|�$M)P@V�����ӌ�[��p��ew��Ҫ�#��=��}�$퓾W8]X���w[v�n{>���-���M���6�-e<a�����~Ҕ:�<,�Z�^�Tb�Sv߰��k�>�鎐��)6�_�w��� ��ȍ�nP�c�3{E�k9VO���.�Uvo:w��0Y�㖮�v5��Sw�v��6�&�SN�'5�V�0��u<Ǟ������sn+Zz��v�ی�7,��0(�����������qŔ�ɲ��Y�g5��=�����׮�u۟H9�&,q�Y�3����q\���jr����MC{n�����ۯ��x�:��"C	9˶��n�	��;rn4�&���铎#(q�u�byƶ���|����q��ҧE��o�Ep� a��L�7�<�c)��y�,��n���C��%�U�h Em��=X�yX� zmZ�v,e��_!^����H�d�L¾k��I��*'��z5�c(=y/�fo!ֺ�V����ӽp�+{��.��Յ�	����k��h/����am�^[�3׎����ѣ����ׂ��TeR:�e
.�����ٺ�µ���T#=��s���fw"� v5*+�4�j���z����)�M���&Y���xy\��,��'��>\��9�쩻���k�>�շ\.�K4�� 
-��-�o�5A.�K�+Ɨ�����g��+�+���뢚�&Ǚ�L�M}֖8�֤BƂGP�>�N�]�G��'3�۫���j����#�׮@�p��9�	�,�]�<�Tt�u�v��W�[�`�l��S61?p=Y�71�OF)e�15����z��[,R�H��+�#�Uk�����T�>�;|�y�PV#f��&́&;�G�m]��C^�e�x��G�^'����+4lM��E|�Pt}��{�_��.��9I����_�����%
ՓG:��^!Y��>O$��`CVAD6�L�M�}'��i,�\,zb�z�p��t6�ִ������4��:���cz}z�;��H�P1�Yu��P	ܑ��\��|R�Ԥ�f��-�)e�s�cgb]>صź��n�!�Q����qXJ�qY*�TV9s�8M�'W���[�B	�����a�lq���[��;޽&�L�����>n�t�Os�=���U��:���N�sn5�uɢ%�/k�	��]�q�u�jd�J��H�k�)k�g�9�~I���[�͡�5{�g���;<���kIv��s�U�t������w�"��܅��XT6[V{$�Q8�}ά�~��)ڣ�=�%S�`ண��2�,*���]���h�VJ�t�br�c�b�۬�}y,���=�X�xo�;Y�����v�J��`m��r{ ��ܼ�u64�1��s��&T3d#,+j��g:.s�s\�����ގr�u�r���j�4f�5�f�n���!�I⡵]�Ox�:�z���|WFu�\�9z����9�v ����lw\����y�����N��V����TX��3 � �͂�j�D�m����m�y��[�����Y�IM�}���+�F�e�|�lӲ�DV�fww���S���J��$К����z���Ɲ�|o7^і��^.�f��Nյw�A9ӻ���h�3:�*�r�ҩ�����>�n��Z�
r�u�l-�Q2��ט1����ם��śЃ��k�v�3�,\��Ӗ^��Ӓu�Ӗ��m��V���_<���Y»��%�+���wV�t�P�1q�Z�0����d_h��Z;#ǌ��u�4�37(!�4MOq+{u\񽞲�*�j#Hdʴ��3ݏS�*�6�C�&�U��Q��^�2��н*7w-E7X���$��`*�M,�wg��b�o.�>�W;\�OH��.�e���#(�ƥ^͡��ƾ�]�"�qe��j��s]�],��G6(oH:��/����/j�4�̖ep���\��Dݵ�dѱ^Q���u�.�s$aF,���,n>ݼu����x�ԍ�<�]��M��v����c=r�^�ܕw��9+�;�밟��Yâ�.3^𫷄, �p��v�g�AΚZ#7���m�;G�ٸ	��J��J!m[�N��9\p݉�����k\�����^(z��W�J(P�I�	(�#>���I/M[��rSYfU��
���7e\wj��u®Xm�N�w���Um�s�.��`�*I�R%"Q����5�U?�������_��h�7&9�p��'u�Rʹ
���R�']8��O4�����l�8��Y���G�t���I`$�I��"�u�5��]��ƽ�&�5*�(�̛��:�d^��y'���J,;5*�����3�π��n;^���n�{z��p�#�'\ct�V�ݺ�`v��.�7����<�8���[=�U�V�`���6����=2��)�u}'ڳ��lY�5,$DCX�U�N=b�hW�g�|T��X P��0Al=0���x��Rʶ��e�佱X�)��(!����m�i����,؇�]wܴ�m)sK��j�Q��)��9,��A Ӯ����wey��a���c���r��TJ�Zk�H��v�I�^4����ز��5���F�ZYR�Z�$t�`�^���ћ���{$�69�5�U���o'5�C�G�҆'R�Cu�nK��w5�nW'�O�M��Vw<X萕�ywS<���f�P�3Oe�8�TӒ�	<��V�9������=U�U��+x�)�kz��]� ��CY���\q	��������ܬl��fw��a����Ny����rZ�!�L�y�h�X���EP��2S;s��i�G!kjW(;h�q�|m:�ݽi�t1k8܋�S��Ǟ�]vyb��a� m��ʈ_^��ʼk�R6V�=t၅/���eܭ��h�������NC޻�t�Cnr"RM0��������QV�*�Q��z�fI��X�;�\�5S���@ת���-��C���q����|~f�c�r��q�n2RHZ�a]�c��U�{�L���Hq�w��5��/=ÙR�31J�f��,�%�y��,ӷ}�=B|
�T~!RD����S��>�Rй�9~�b����'�H%{κs+qoZ���1���u���nZGErz:U�ua]ѠH�Uۚ�zGZ_�۲��]Y��V�V���q����oy��ݹu2d/��n{�V2��`Xu�V�*��V�.N�xS�F�6�屭�f�IϘ�G"���2�'�鬝D֨��S����F�+E��gR�����{�l���E�7\v�X��#"� �n6�c���8��ǎ�F���2�X󀝻+�ۨ�\�n��l\���:���0�,hMbGa]ɫ\������`x�
��\��Z"WUAcw���?@tJ��8B^];��#�ƪ�9V��^�n8�=����ּ0����}�����3�G	=�t&뗖�����=�$��Η	�>%�>�\xy���2<@�/�=)G`[�	ؤ:W5��h���'���ܽ;�zݭ8�Ͷ��d��!SI�uѕ]ߊ���7Sմ�Բ�_�x8j��%ޙ�(�V{�(xJ�\��>=��%�������h�!\Q��S��s3���U�kU�t^9-ۇħ�e�l���ɓ2�_�����L���&�J����[�X�ڳ�dw`يK~r�P�v�Ы7F��/oRpZ�揟�$�H��/F7�f{�'%@�Vmo+Ũ��s35{1V�-
+��b&Lٽ7wO��;q����Y���4oe/q��o���J�x�����8z�}g��Z��0w�p5o�]J���H�4)ʂ
�*�<����צ�ѣ7�kK�c(�˶�*�!&�
���� Eμ��mL��{PL�KA�0X�#� ݾ��Kuf�-A��T:�s��z���Y���8Z?����d�E�fV�!bn*%��H�z<�`�[�����ӥ�t��gCh|fs����9����_�W}��">� Sm�}�v����e�KcY ��`�J5ۥ0s{9�X�^vsGm�O~�&���Oq˺[&y�A�2���,�� �A��ܧ��Y��h��4��+*�9V�{#�2'^���?�ଽ�~���@u���⡆��ʧ=�k6��Чu��(n�յ���%��O;ӹ���	�ǝ`&,��v\��f��6�/j�]������Jt��;�M�Pw*}�M�-"�VJ��ʭa������ެ�3jm�2�ۣ5���r�fV�S;��"�Oޣ~����pSP�b�϶��B�V�h9%Y�=5����w��9]�Mgө��
#��2� g��ڼZ�}+x�E�<��e�Q�Gn�=R(�%�lu� ��J��9L�+nA�+V�痊���k�ۆY��u%��*�[��Z2�����3���&�"w6�Qd�~����Q�=�[��6�꾺�������or+ٗ�����{�mC�R¹S��u�c���md{o�Z+�v8xԏw����Zh���=�S��W��$��Ǜ��x�/k<r�zҼT�g_�|�z,$�Q�M�]"�̶3Of��d��~��("�뫘�����^���ݍ�Q�݃���9�Z�e�'��v�fV��㰻MIZ��m����ڼ5љիkN\w����KN�'��`��7B7���g��RW���}��!uk���|����i
�WwKa� �C�潺��/��v_)$�<ԟ+��֫�>o��>�xN�����mu{�׏�6ϥe�b�e���J�����͹�׷�L����ͅ��
�Vu�����.Q>\6�3�ͫ��o�uCv|���\��u�.Go�Z�<�9�i��{\q�=\��n-��F�7hj��cj.�ӎj��N�V���O�o��=�5�*x}�q�w\�8G�RV^>��k�;;E-YG�rMx���#ޥ�x9yv��\�0�4�*��=BjԬ��[j��/�JB{E�G}�P��Z�ɦ��V��s<�)�QdW���ҝ�R�xV�����m�S�&�+�C%��pY,�sO��ӎ������E�T�M=6-�U��pJ���57�{O�yU�Q-��+v��ӹ�2���XU��q"���y�$e�L{�=����t�]z���[z��r!����t}Q]�&���Ɓ�%X�^�eY�;�았;�V�lZ�&-T���u�� i�EV-�op�Ʒ9�{G���1rh5u�W{�Y"�a+j��[����+�{���!�ٗ��7�s��X4�5�S�*M�ו�טEwZ{v�#�:�r��Y}]�#Lq�eN|�Q��Q��fm[�����dyy�^8��gl��lr^^��N�S)���o��{��'�W��Ewod���ѳ�1_w���_�����z�.�^Δ�Ի�c���`!��R*�Βm�,8���:��~�i%423�>t�UE��펶�OL�f�ޕ1x6����+�޹S�s�����lV�n��U4���@�>�JF��f[i��
���o:(
��K����m�y"�+���i�];�vc�溕(!��/ZKb��Z��������.��>�sg
���p�/7�l�6k�$3�$frX���=�pf����s(�j�+	$+�V�q��7�ݔyd�|jS^u�
Ρ�4�{}�2���#���'q(���W�ߊ���`�u֎����M
�-E[�|]���uA���X�#r.�T�^�e
��j��S՝���Ƿ��ݽފ�L�,�:)P�)LG_^gDRck�7\m�� ��(5�B$�S�]Ĝg6ң��˱����u{u���7k���ٙk���.^�����v�<�'��3��5�c55٣�z8���M�,��4;L۸�N�5��]�R����q����6�;q�Йn�f�f�@l�ػr1�{on�NTl�]�:z=D-á�g�Gg��m�K���Y���Q���]\�6��v�kz�l%�-,�#M���]���%�x�nq���*��"���WS	�@�]�<؈�1oE?a����tm���&�<�=^��oѤ��LU�=S�GA$Q**{S��[L��A:D�֞Ӳ���y��/��q�̤ܘo�����խ�g��{�M�6i�.swpZ��o��q�7+*��-��F�M�5/����𞰼,Bq���8nVm7���{�Men����J��1�.�I8]��#K�h���SE�{9>#4�F�Z�<rvl��3�r�*]9sS�4�����.'���yרM���O�Ĕ�6�̃/��>7Aߔ���h�AL�����Ûf���Ǘ���g��B�֮��Pz#��F<cyʇ��O����B9����1nW��z�O���;�DhnBJȭ��)�an�rA[�y`��;,��˷ls�S�O�LE����j�x��]�Vz�K�2E��2�B�<]V�����~a{�bU��;��P�k]�ZH��n� Q�[X_�$�u�W'��B�Au�ea��oە�̡Px��i���1�j,5.��J��5V��rձhY.,�I�W㣝ռ��g�^i-cwz�qw^մ����L�ף�'yt����Ȼ��TO'������vyV�I)è�d\�Y��Q?�RWL��z�w^>Y\�%ҹ������EJr�̢�z��=ԍ��O|�Aۃ�۳I����j��h�,�rU�L�5}'7I+ �k}���{�Nǟ]`�C^V�{�W�[V�|�fG�	Yc��)���y�w0��Y X	�E���y�#(ۜ�9e�[m��T�&wvuwAr)�;:�]_�9�QѾ���,��Y��+C�)�י;���버j�t/	�n�X-[���d���cv�����E4[��1���!25n�D�8QdW�;�R���k�}<רZF�Q�_6�5�b�\�N��E=��?LK@�M�[_�_2����t�pX�~��Shr�y+�^����A0��괇$�s7dako������Y��ǚ�K��B���L�IM�Im��y��m�v?{S�5�+���כ3io^K��
yB�lݴ,�N����y�e���v-eu�]�M�ﻃ�[��}�q��RA��Qm�9���g��5�ѧ�c�6X�|�[����Wb�ŭN6�y���:�Z⩨Yl�֚��,��=����Oq�Mw���H���z��b���{��V����FF�x�&���w��.�m�?���Gǂe-P�0Ss���>~9��{+����7S�-�W`y�R�ɾE>�yu�ž���b9����ט�f�
*g>Wʥ<�¬�2�,� *��ޛ�՗z�;��3�mcosvn|�ׇv츗eN�܊rti$@�4�c�W�3�Wjgoo����s������Њ��+s3K#&�i�w7�zJ��g�V��O�x�EQ����'��D��ݔ��[�5�t���Ϯ�A�{����^j{y��z�oE������ϫ���c����}����g
Tp����ښ�$�N�
�ܶ���2.�/�c�4]M�[�S��݉vŖ{�n��+�V�*V���'6�d�����fb����TQA�Uwv�w!d֬ �ex���Gx$�ۛ��ױC��;���u�n�Ξ�^��4����k�F�N�F]�b#� �QWݗ��Rm�6���jf�@��f�ͱ5U��ˮ�i�t$��U�%�H�A��Ɔ���U���S�xWo{�Y�1EQhRE��Y����<7y]nd�S���z�!��Y�&�t�U�*�X���,�B}�=�<��8�un��l��k���H)*q�ٞ6˙2�m=nqBq��&ƫ�����\Y�ͭ�i3b&iMKt��)�- �s�{�l���;�yݾŌd�9~�x3묧O�Q�Y��.�P��R0us�ҁL�4@�A4�n��͘W��Â���_�$ �������]��.�j���mʐׇ��/Sg��޸9��ݺ��WV�L�9��4 �|�m�{'�W2]Ύ���ڜix�?3�训�t�H��|����	�����١�*r�Ϫx��m�W�#��)�IN%�S�B�v�a�;
S.ߣs��na3k_�����3�*V-���pW�����Y�jIG��W��R�D�z̩<jz�
���t=N��fw�w9z�]"h�#�>~������^�^�;r����<��t�c��.5�xV���׷��u�Z�}r;�K��m:�#�U����w�X�wθwn��@�
�\��(?Q)���b�OC�@kkP�&��n\󞷆7�8�|>t�e�[vt�(i�섒{����ǻ3�l�'�z����q��bf��
.��ne���E	}���]�����s�$��I�q�R�uH��3$]xn�zE�Ie��Vw^�#/�e�1����9�&0���К��񡚎e�[dum���m����޼X�_>th�x�!1����Ѓ,���X]�/:��CZ�J_Lv���܈�,�hH����5.�N,
��c5���U��D���<��f�V۷�����*�㮽��ݠλ�[v����ѐۻ�/w�'^��v�f�D0-�CM�vQ���TO���n�_Y}]�ө���8�I��v��������^E1Uݭ*�|�44�b���w7�Co�"m-��n�&�t9�r#3��My��\�V;Y>����Z��4�n�n��mՍoj]]��t��l�vc�v�׊��甥�2��uK���V�F*Ұ�t�$�t!��}3U��/f���NqC�rnG�-JUz�,{P����-�.�@�B����d���ͨ����WԵl��lL�$u!�@~��lO~/2�{5�-HV�ܗ�̝y��f-�Xq���)of���<�.�*i��Y�B:�4�V�U2������%�p�ڶl�m�F���b^�шh���[%���ǛŢʂ�v�b�6�V�����L���N*�QI�`��fp��]W����{�	F�Ŗ::���F�7=���NS��Aj��ttހF|\b'=ĝ��n#����k�6�6���ǝ`�$�m�{:	��c�(��`��t<?�/�|��Ӈ^��z��p�q��x�;n�۹�C��+z�+�v8$^��dg[���Tv�Gl�����'oZ���eLs�hwn�{n��vܓ�g��c�v�x�:�����I�q�ݺG���,NK����nn<�q�8�:�������97��r+�:�p�˧��˶�ڸv����@c��۫��쉝m��y��:J���\8wK�;���"U�Y��)ŝ�Tʛ��6�s���z��.-����;��uv��{�=�=��^��c��˺�k�m�6�3�zU��{q�a�v�Z�s��xZ��8�v�=�q�K�ܸl�b�nӸ�&ΊޞޮcN�������h�:��c�f���b��0�b[Vy���I�el�lh5ŸP�6��9ţ�]��%ǣ:�.=v�ι�6�S�,Lc�n��G��;>�V�%�p��s�d<�OX�&`]�;��:�[�g��ڶ��^h�1�u۴��ō,��lƍ�hʤ&���;��vGql��=Hq[ѳ"��`˛s�v�ٞ��L�ɷY��CĶ�g�8�9�l�BF�u�{b��ݠ�x���6��V�[Z��/gɺQ���	�ZUc]=�-�i�ab3p����D ��W-���M�t(���Z0�(1���{t5�Ru�cqp�Lnp؞!�㵛��sc���v{�#����p��u՜m��k9@�z��қ�g[sV8��uç��h�]����c�l�E��U�tvv�g�֎�`'��(].7�8v����]V&xG*8��xܹ�'�ݸ��i+�cH� �uc#��H��nw��ui;qq�s N���>;�v����%.ʦ1�T9T@�� �n�Ҳp���Ս�p��n�������0��e!�����b<�q����[��0\Gl���n7F�����-�9��ڭ
�CRkQ˗A�\��j���I�n1��x/#�L<8�D$l%��Q�˹g�7&HM=�T+�f!�z3�r�l�W�/9�\n��vH�)��K�����g��)��ŀ6��"l۴���b�`�E��q]����q�lq��n^�9���7�b���rK���租�S���	|��v�u�ʽc��$Z5\���;s<��ӻ\�p��:�[<jV�y͕qx3���
v�ycn�rkZ]ӻ�F���Yg�����dH��!~CǞ�I��	ٛ&l������9D��]z��]���=.竜Rou�sU�j�����U�![-�h��>��H���>�r�+F\1�u_4��Ls���q���򩛛��3�v���;YR�q�I�q�&HH�
,����d2H�&Wg/W��M���qwy4ܔ��hс�(�;ݙ��!�+��f������=FGDw�X�
�I��q2Wm^Ύ9Ǜ4�^�d�x��[.�*ϝ����MW�	��~ʔ��{.����%�ee�j��X�Ê�Piߪ�FZ��X.��q���f����s���l&�v�ן��wnn��S�U��y�¢J�"�l.��I�S�����3�n�  Pء���3�׈Hہ��Y6@�<�B�O]��=+uD"�;i��]�猹�r�kmlZIVv����%��T
�.����Íd�^�,6~�^���r�c'��F�h'Ղd%Y�32So���{ݝ��o3y���A���o��	�*�+�z+D�{�u�+/\prJ,2j5�~�Vm��[uo<X�3h�B{0�ScO@aHбV=���SQ^�?	k�2aS6����s�2�RK�z�N�G*?��d��E:��n�a�֡�r�
S�[.�x�B^�NZ�5�򱕙���RU�7����D�_�n��ҹv����=���N�TYI��Ōu9gL���a�>A�V���Q�*�����j��=y��G>~�+�Q�QJ��Ok��~����g�f��a}C���'R�-�(&��gqh~u��;�VW�*�Ȩ�]Yӽ���+,�������}GNu��s��>���G]+zs꿨�mͩ��{;�U*��U"
�S%\ns�.��ĝ��堻.��m5�CX��^�推�.�i4S(�e'W�K�IPw[��+�G:Y��+R���껯(b>��z��5$��w0+�ϥN7��e޺��T.욗��{��;��;)-\\V�*9#�y�cM3�iQ�O��s��yև쎺�ܽ��ժ�v@EM��/��K��=�p2����T�d�KԾ	�� H���U�?�Z�J���mJ˧�+ ����]Z��۝����/Lݖ���W�������Ӧ�&9�<XR��q�#͑���t7h �K	���.�;�[�'����O�dJoej���:A�W����|��� ��lQ4���ݧ�E{�*ϩ��J3�u$�x��s��
���%�.�����A��~�8�fx��Kcj+����#C���J�w��z��K�+�hmև�լ�L�=WK�ŤJ��̘��g���M`�o{v��ISL̔��s/=�0Y�]8ECE���x�����:C/=m��clۧ������g�!M�W��i	����Vs�L���\7���׏�`3-�"z��{�H�c_t�f]E#�;&u�/t��;L��^��C֗i�����jbq�UҲ߹�i�}���d����:�aob�?:Ͻ6`��ܣ$�������y�,������o�����w�0p�� ϳ@�M"X�ٺs	�"ԛS�=�O*�^���/��m��5�L���Mݘ����o���C��7Cq-�=< �P�T�/X*�Z��t�:���ԸJ~���o�W�n,�z)B���	�u�ڳ�����6
�8w3�rk3���t7�o]F��7�aا��[	ɵ;6j_r	f|`̨�TwF����W�@Ozo_BCSGw��{�h[��+[A����DV�FB'eY�V�T@bw�����ž\�{霹C{��z����������M��0�1�y��ye���grQ����>���b�fx�;�S�nq�<o 8�˲���5�ӹ���|�$�m	��A�w�㿡
���4g�,�p�-[1G���=Y���']���O�r^󿽏NA��5��Q*���xz���"	V�%e��Uf��V+9��q�Ҭ��R�06��+!�?"���.J��$�{��7*mN2M���(=�ƍ�� ��ӧ��Z>l��W^v��kP�G,��_����:���n�_-fZ#�ܳ�o��T���GV.g�|�2�S�Y&ܤ��%�Еmm45�WRrjͿ.J��\��k�i�[��eٔ
�+6K�8p'�멎Z�����s�J��ʖz�:�Ŭa\H-��`N�
�Ejr�������A�������K}@�r��F�:Zk��w�J��w�(��w�k~	��o�J�����z��3
�Y�Dm8x��;�����P")�0�.w���kJ"��o�v���f�@��,A�n�-��\���YEk`+ cM��
9���st��/y�nL���s��rt6	ݰ�<g7	-��v�l��;93�[c�<�x���[bs��,�i��ϒ:�7��ƳۊqQq��7;dN+��۸�z�Ȼ	�23��Bu�=�l�g��9d���Tg�����ɗ}�5��\�o;�VXLc�y3��l%�[�����&�㱫��g��w=��90���`q�}s� Q]X۠�9s�-�9ö��i�]���S�>�s��4
X�*�S��I3�e{�Y���u�wO:�<:T�2���\�Lg��VFS5��)�⫄�� ��b�Y�$&�j��2��凤歲\^瘲��.�?�C�������O\�����T�<������F�>fn����G�����L��H�2�13�p��:�XRM����=�}*1V)$��NP��Y�MA}��歚z�mm��K�{)MB"�s�+wD�R�U2�/�%�U
7DZ!viM^�c]5����8R^��]�G�0we
�o�� �[y~��]�͛w*�ݔ��<:�u������X�Ƈ&�����u��_��*���뼻&�Y�ή�@�UH ��gc�h����0`{�ִ�*�X�R���]�{�̑�����c���1U��jt* |fC�i���Кt�b#j�m�Q��v㍞̼�8���m7'�j�ݺ��\PmؠE:��B�W{����#�����Q���|�� ���Y�9&��}k�fì���$��p�%p/�&{%�x�(��XESm� -������.oy?��]J�x⸬��e���m�v���]�C��Z�)�|:`cߦ��|Q��K��IkgA�6��b�$���hqo�$7�1���4��3Ƿ\�W�O�S=��4E;q�[�>~�h,�ծ�pW��7�o��5;k&A�?*@&�d_�t¿[����Y�2�7ד�w0﷮�'w.�zA�{.�u��5���=�(�S}�.����o�5ޓ����}&h��>m��K%(Qa��Q4kUM�)��d;�^�ax������+��^�Gs��Uh���t]�˽�D��Lg4��n���u�i�A�)a��p`*��3M�	��m:��g*�+u�7t�b^{��uU��|Xu�u�}[殠(Ţӆ�����f2�����y��Ύ��ln���fu��g��o�Cѿ��(S�YUVBV�����Ǟ��1q��M���<m�~�{|��km�\]��-���o��l�U�{����v[��}y�+��ج��>�Nt���aYc�P���mg:��/#u�tr|Lb��F�t���u�F�z������묌:�dӣ��lF����cmy4h+��W��K>�����ye_��w3���uӵu��i!�hȸ"�9R�K7�bwDѩ5þ��g�Q����m�:���켽� ��_�i�ESt���uv��'�D���+�)F�Z�{���b�2�E��%0Ų�:�P�������K��i�<~W��M��nd�����>ķ�����Q��q{i͍���P�o���:����%^�}���T�uX�ާ	W�ъW �a�l�9����VNfQU�^����f��+��M�33���d��*������vQ]���V�pXӈ�᫨�#~��3��A�GK�]>�w�D*E����ʳzrt��)�Z;S���M��C�u���s;�x�2���:�;���F�+�N'Y"�J��� 7U	l�s����F�C�=�K`B��f���]F1>�RJF�f�hW�z����|=Z8PtV=�讽���2�!V7�`x�l�H؝��bw]���q�);:��d�KY�m܁��!� ��jV�k"��^�$g����^R<�Ox��XF޹�mf#s��{��GNC��U)S�;	-��f�Mt4�aw��M���8����,[[x37�x�Ch+4��3 ����Y(AR�u�=|!�F�u]�#�aS@ i�S����B��F8S��>����]�:�l�T�O3�F?7OI���U��i�+��O�<�u<�wE��{--r�O�*ʩ5�
(h��& eY%7�#x%E�g��̣H��gV���&R��kbϓ�6ϧ��J��1*.�@���0���:F��i�V� �G��	`h�]Xc�y!����v��O���v�pt��]Y���W��=�*yo��kp
�o���Z¯rd3C�x&�9��y�v[��g���������n�W5�"5��N�k۶���n�[�}��c��V�-�)G�4��P&k����QLF�]�8z!��};'jq���U���ƙ(W
z׶��D}$�+;k���x��4�_:�Ɨ���jw�#�t؎t����������)�tДd,N��{�J��f����U2Տ�H�w���Z�$V��kڏ��V���G�Bn%x�?�8Vo�����$���g'�k�xf�F[ �^�����?{�m-����z�8��a�$V[��*ˣ�ݺ5��SͬF����U�h�����ӿ?M��h�����[�S�����'����M��`��Շn-�>?9Ү;>�-�ȇ֥���1,,=&���N�q�>�H�
�K�V�2K��r�u�KT�zKv�vS=�f��&�}t+¬[���w�=�n�_w^EYnCf��J����u�m�����-ˏtѭ�����܎zZͧ�L�%��������q]]�%�)�e�������۱/4�O���X�ทq�][��4/m�峴c����}��C��t�wgO<��v�oL���{n�pm(��s@�k;�`Ŏ��L{>���u�ڹ7�����6õ�Lk��׶\N9��;:�k]z|��q��@v����1����]��q������\v�	8���N<�M��1�v�n��eѵ՜��m�uQE��H&��s��n��^�N��o p�5�;�}vg���9;v��MnQ��WL����]v���ض����OS1�Y�n���(}ߟ�]�����E�{>���@�c�2�{�Ƚ���3�����^�LQ3�ww{k��>�_�b��:�㤰��U�i�o�G� ʩ�mi^cK߰|�fFg���B�)f���*�Uj��@q�u7�}o�l��pp�������v���,�a�*�i�~)�y`*��}8K�U�/����u�]���T�;�Y���u��2��%e<�ʎ������T54�W�9�5���R4�\��-��W��
��<ܨ�%D�����/���D���2�6ŝ2�_�����������T��$i�*���m�21�T�ic4��7��;�=$k��!a���,�	U�n�E��x�I��Pݨ���d�	<|^�h���t������<�x�W�P	R��t6��n.���G��:5�k�Qڌk��-�GҊ����Z��v��[���o��c��ɻ�vG�Y�4U_�^���ba/�W���:)��j��/�3M`���Жj��n�ղ}�*�y����e���L`���.wM��qvfչU
�����v�jb�9������9�G��K��d}ۼ�)�2�ِ̫�5
P}�pұ)7�{�^M}b�5o��g�p���w/���7�6X��L�p9|�l���xJ���r�L
�⾤[E"�%�E��z��61V=�S|�@�a�޿x�^��<����p6���f�Nv��x*4���Yɇ�w
;���]�5���Ϩ͡X�RѰ�Tf�J�k�|�eߗT��9o2�����*Q*�]�n�6�睳����Z7ܩ��1�o��=��ڟX��c��{㥚a:N���X�Y�#bߕo��
�@X�)��{�L�端�8�m<> ;��>�h.�ީ�uե��EARoz�ٕ�EU����X�7ɓ�P%u&�ޤ]:sù�����'�){c��F�cm�u�맞v78����[�gu��uc���ί48ƻ�SE^b� !5K.��N����N��)4�����^0���D(��AV=;�����W  $R��c�us�r#@j��R��9yI���\T��N�� �����zT�ڛά�����*[��|;��U����O�k�Nȉjj(��*���E;���I�?M��&T�O�GR����l��׶��{f���ߒ��̕{3���^:^gVk�X�
Brw(oe#zeͩ�y%��r��U7j�1�
A��ꅝ���6]�FS�W�\ط)���7J��nDk�5� �j��i�ùN��Ѣ��D y��N�)�����S�x"a�jx�%���A�}N��}6�P�����eY�s���^�׽s/Ir�ɕ�C̗�>5������+;�������3v���w�:�Z�5v�E�!�X�x7y�/|^l��V�F͂���!X=��L�exq�&������&�*6�3��t����m.jخ�c��׼R�r]X�84vU�NL!s�w�+�*��`^�0��ajt�f�� ��B:�+9��{�7W`�C2:��hW�9|���n��˸�!�]��!Q�W%�����N��-R�,:�V�]�erUnN
��o��w:�n��B�-�l7Yyӌ���Y\~�G�$��R����z<А��ƻ~~�{�M&�G^)�j6 (�["��c�U�B��N�|�Ej���4w+�W�2$�%c��_�#[:�/F��/t��.}��M��8b���r�V��'sE�}�m䡸���������q��{1/�B��:�T,���0!5��%�pa���ڳ�ח��]C�|����s����$�[�g���mr��"���e�ے�}))�Iy�p����2L+�xo{ �mͨ�k^�X�q7iц�2�-�w���|��;L��FW�A�U a���ֲ��Zq����~��5��<2����1牐R�@�s�Wi��m�L��n�0uE�Q�]�f�u�A�Kk�vo7kv.��Z+R_ ��{�%*�ȫ3�YW������}���ǁ�SJ���)�S¼���W��I�"�L��dL S���0ޚx}�'쮐#PV�Di �/�gI3�ٯ+ID�������[�٭1|VO_��CC.����yQ�����H��2omqq�|�N m4mڲ��t���;3��^�{o^�۵��E�����H2��E����%��/�错��)c �@Pt��]��=ژ�;���)���P}��]���j��D!���1ˋ,�}t��{����m[i!)��]*T����03���{����:�s[���Z��WM���Ͱcj�&N�����-�]��W�1ݨ�^k`�N�����s�?6�l��$ݫ.  ��Y�g���-��-X����6�>u�J��k}ҭ��we`��Uu�1�~�T�:��ݜr"a��t����f'�53�|9����c��G�6*�Ԡ���smL�l�/Z[�v���Xzz�"w�-�����,�����{c{LJ�4R�yװc;�P�oC�u�W��cL�$k��]l���2������`�`ToH ������Ǟ
~\|A���-h��(��i�a-Z�^��b_Ht��׷�M�
�Z�S�eO��zzg�����_S�u�̂f�zǙ��YtEɜͮi�re�4ؠ^��;#޿	�C����$�V�u�1��"nw']Xӄ�=�M��`ݜ�S��H���yf�Q#��K'���BB����I�y�{L�t���X����	T�X�=Y�����N� �m���;:�v3���>��Y&�5t�l*�g�_*��W�$��=��'on�l���Rd[У\�S1k��Q5X�F=ޔ�e�d@9w^�����$�6��P0�R����Ũ�	�[_�u���Y�رW��>��p�l;�]�(.��o�x����|��!V���������O�AT���,}�����^�U�F���y��ɵة�I^s���5~7�_�A��g�}����ʟD���_R
�C��+�H���O�:�z�r��"��[�m@�R%��e:�Z(�e��f��\Xr��iIb$v�sa��"��:���t<(Q�;U1FN�׌���:]���w���.��?'h��g�]v��������ύ�J!>�B�끼�f���^�BW�LX��u<�Ŵ���ە��v�U&E0n�8��4ՑZ����A���߷�6M������Y�W[�P\4�m҄V��h�v�8��f��3;nn���^ں���lr�z���m�m�Dެ��8��ݳ��K�v��H��2"�W[kG�RZ�3/e͹���O`���۰���P���kh�{���׷##��n�;ݺ���K��;u�mu��۾��!�m�]�GϦ�u�nri�b'`��E ����cW6x�Op�8���o/=�ֹzV�4�غ�s<U�}���x��X
�ۉ3�T����S5UO�D_ٻ&,o/�{�+9�o]���ls8���STWY{Ƴ"�$߽B���s{{�UbT�Av�2�8��f�5�{x�I���22I-�G���B�4'xI*O�I�=��}b�����v����Â
.#>R��*�j�B�<6
�tr+~�����i�D�*B�h���) 2�@R%���|�dq������=�6j��~��@̾��������:C\P}��/���S|h `o�/�]����K>$�
���O�x!��?}`�V}��<_-�w��0ݪ���}�+�19�n��X�0��V�:��� �(�^l�V��!�4W���~ֵ�a;X��Z�Z��VP�	Vg9���U�l=�mi�WC�Hs��݅��t�Q�/ھ���>�Ul2�\9�_}�J�I ��J-��}��E��k�N	:�+���c/�(�k�4v�]��v�By6<��Ȼ�h��
�i0����n�z�}%ƅ�+����Kb�OGY�[j���dr�{ީF���K�̩~�(QYگ b�	�%u�
��ڍJfd_H�3@6�y
�X(���]�����Vh�j$�,�x��j2�玠y)��m�w��ΗR��	�4:��;�u\��E��\i�qc]�<Y{p�EU'�~��̫ݤ����	��9B�NsoN���ٳՃ�2� �Z)ne�?贈Ti2S�?*���]��3�M&�w-�D��s'�ψ<t!������jF�6}���߾� ��\�/���^q�{kA��}�ob�n�BBM�ߢ;r*[) �]�5U�,�U�vב�^�KL�"�Y}L|c�X������-��a��9t��=�R�{s7�`ߨU4��~���G��L5BV�A�L@m�,�����i�)��c�����{�r龮;�|��	Ts�`Q����u��_G����Ҷ��oe]x�"�e2$���6� �%M�Qxy�Yױx���c��뱺�0����pk,<@��в�8RXଊ؊BW���.tR�`��PT�]�4k��m���\�2��0ھ�O�����M����y���h����?(H���}�y0p�pN�S1���z�n��ᒢʞ��>�rg�9��.�7��b�S��4y�\�+�pe3=��+E{��^�R+63�wt(]��[�[C[��}Sp����$�NZ�-��aP�Pг�߬w]\h�z.����^�ASM6k��d�h�ƅ����:z�oX�:Y�ү�ͧCJݵՍ�bZE��v�/����U�z�ۼ��M�����T�cs�>��ꕂ�Q���\��~�jxةx��B~�R�v�|�m4i�uy��^�LV7Ԗ�ZC���a�v�w�d|{J��c���	�ޫ�\M���)�ü�����f��T����u�]ו����|��}�a{E`�-RD��u�:�����ޟcX��V
>�f�Ǘ�����ހ2�O�}��a+$|�|׎��W��?X��{*��a�o��ZR=}�p�+M�h�UmG݆U/i팜"���pl^��[��7n�$�,gJBiˉn��O�4D�D�NN����.5�f�����9�I���v1/��埽ǟ8e����cT0�*�z,S���R��$��ޤkST�&�I
�y��,q.�*S�s��K��V�Sߘ��At���u���NV��]��[y�'��B��k�p�m���y�C��}���AP|�d�Rn�T,�ڿV>U�dn�;VԶ`OWW/]�E��&�X�bt��9��׵��A�碬4��q�9\�~Λ�LI�ҝU}T��)��D�L�	��A�{vW��cT��CL�g������߇:d�NT٫�W����]��]�o���s����ǅ@�*l�6K&��ꥄ�\Ƙ6����� �+otK�*o����W�n���-�oo�r(���^�\�W��Wp��Oz6�RJͺ�3�>c�s8Ag��vU�r�U�P�ˡ�~�|������y�ucfۨ(����k���K/�((m���0����w�v�
�,}h���������Z���;�:U~�,X�,4�I��s�����c��%#�6�6��,+�P�s�S&'b���F;)T-}�K�5�b�n��w�p��%�6�4���ҥT��{��J�s����J��Ѻż`�VU`��w{�����B��ɿy���l�C��o��Z��Sg�k�ή�>�1��J�{�o�S��0U��ť�q�5���h�y�m�ֽ��?
�7�*�� U�A�\��mW���Q���V2�ՋYȆb�z�!�;�T�䇍Vʚ�S�_���w����Bo#㗽�+@���+|lTO�|T��7K ���K��ɋ{[�����R2�߱,��ף�~��K���L�ޡ�������o��X�A�i��R
�R�K�,�[��rf<ZcY��Z�^���߹r�RD!�;Ղ=o,��;}�WY�$�>U`����>a<��`�� Y���P�V+:�;�`=���0`�PZ.ڬM`�h��� z
+�y��[�IF���P�5^X0���VQ����n�� X�o��x���w&��U1v����'V�{�r�y�ԯ��W�ۗ�q��Xݼ9��74󄷍���:unlb�9����÷:��-��[�Xx	�9t!�����ۧ�{����!��L1�<���,7��n��>�n��(v���R��z:�g5͹y׎̜�糀[z��;@8V眆�n�y�\��,q�<�(q�g���r�lqi���q��/4��ܶ�*R"�����"A�ȝ3�\=��ƺ�\eŏk\���n:�
��om;�y���%�m���kq��ks�@cEL���ԊmqUv�X�W9�SxB�UV�?��þ�چ�����x�i�����+Z����~����B�*t�(sU�j�ݙJ�
����&�|� ¦���{�M}�"E��U�V:]�o�_� T{ً�gc�d�(�%K޼P� �LT��;�R�S�|�T��zV��3v��)r��R`EB�G�~p�.[\n���U����q=��u�����i�i�ceE�Yvh
�P�؛�`�X�c����5�sC���S��{��ϸ�5�j�5:yE�؂��Z[u��I��\���˻еY=}YDSE�*���c<0g�%e��\�E[�+ECLt����23����ԧ�現��{��Q$�����VS��D����GӞ\��ڻ��v�ug�[?dA}�A�i�t�|����t�ǻ#<�v�˞�zn�_����rW@.�C#U�9�s�;3�%��i�=�W,M�aF�>��"뵖Z;����ð� ���pk�֎Lv�I��I�i��C��>�kT�n5��*y�}D�M����]����ף=���K�����EVmE�x��ߪ��YI�C�q��-E6�]����q�+W�J?r����[��L).-��w֭���`�}��I�Ru�;̤ Yo혆Tn�(��3h[xj�m��z*f�WP肺,q6���^��ts�=f�ά�ͼL�K�l|�}�Y�%鬥�פr�1G�:U~ob�=���s���tM�Q�r׺����ͼ�UoU?|t̀fo<:�E��j�}*; |������^樽�x�k6�*U�ee���*��J�U:��|t��߶��L�S!L�\�+���>��Ŭ33h +�dޫ�u�\*�v"��{�UN���{��W��r�
�J�8Ry7on�twR��=�t'�+�z;p.�K�I����*�Z�oy�O��pk轿nZϘ�>�i����KMf��w�+�XW�VmhШWx��:꽯0O��#,{^1�Y�o;�+�#��35F�������vzw�P�'(}'�m�1+��J�y;v{z^l]�n�ϗb%��dRtE'@SI�p�h����j��~�g�S[��_O3��8�}�Su�xwue+�8���ڱ: �H��:����.zVS�k�&��X����J�E2��RY%��Ɨ�晗_k�Xo�`�tw�cq�s�c �V�L=�K���V,��"i+�7��+��ֈ��?k�Z��T|�:|�%����nׅ��PnX�"vٟl�*�=mŮ�s���DS���5����׎����[��y�F����ڈz��� �܈jr�n�(.�t:���o<����zz�^�eլwK�6�����u�a��m���[����s*��L�Ҧ��|��k�S5��a{�͑a,e���^b?���v�y(��'��*5kʨ�|�aHT�����;
Ss^���eo�}L&Xu��y�r����ˮ�]V�7ڞ0��餒n�_�O�~������a���:|���S���;�B�/Ւ��U�e낄5H 1����yB�4ct��� c�
h)Җ��mI;כ�����g�[[j��'sW�#xN�<vj��b�O�j��~�v>��⫐�皘e�I����R���*���ԫ�Yо">�z���}�����ݑ|
�R�f��+\&�4�0�S7w�ӹ�*X�����.G�V�֨�Kٞ��d�D(����ܙy[����}���&r{���Th��V�n�f-i�O"w`Y5�^�+�����`��%[�n��V��[���+}j���:#��4�a�J��߅e�k}89t!U	�z&���ӟ�s��h��޸VP���>�[�y(	��|�STiQ5PV��7�r>���~�G�D�)��-6.��R���e%� 5����*���s�X��Z�-�t_V���j���3<2)�����N{���T���#o5 �e]#�60��Co;�k�֠3����5>����Vc٘j1�[ɕ�.�;ݜw/�w�rw5�Kn��V�͛z��{Ŕ+�{i��h�,fڭ��8�jo=�K��X���ms�N�F���j�d�<�%��а=�p��N�+�YW'd���;�Ə
$ح�z�����L��Jd�����,��5WX]�{������{�t�5(�P�ۛn���gǑڎs���l�v�z�39L�$m��'dhUD�R)l���)��q<Do�@�x�<�]�w����j����}���L��f�����>���t�yW�Xɜ�l�\W�:�X�*���A���^�v����W>��k����s9��h����=G���L]�Og�dQ\���ß
��������!�g��M<tT�_w��ap/�c1N���Ŝ�t�o�LxU[rGdhv����х۱b�"�os���ԋ�R��~���*��{cÈ�3�ٗ��C�p��J�՝�Y�U_ :����n6����g�t��L�BV��hg����ｙ����M���w���3f�AJ�u��$��^rJ���}V����	R������r����ka�b滽x���h��~[ M��h`�b}LQE�]�����Ϸ�i�1'Q��]0m�[�^�Z�,SMU"�r�2^=�ID�7��D!����>�ѻS�^2k���b�A���Wn��,��sV�q��Uv0o�p��*��%�4��sY%͖&R3q��n�����t��Z���%�ժ�;��7U��}v��6�r�k���&�������X�z���ǥf�ʭ��*�圪�0����vqq�}�n�ث.\�A[t��s�GVX�,�8{��DFgnl��f9q��N,���9��+.=��%my���ז�^T��o-��Bɵ�B��v�E�L��+��F�SU��'a�����Y}�%�Y�-���XlELe����%ۧ]ph��#'	ռ�iF��ne^˛��I+��m��]J�
�Á�\@��Kf��7�C���Ѵ�i��D�	޸���Y�ةgoe\ژ�0:�P�J[ۃ�=f^�=bEr���F����K{]��,4��NDF��ћ��]��F!c� Ȟ�]�ᕚ��&�5"�)�m�p����.]	�H�9O�fL����n�7&���X�5xY�&7v�>�da�U`��&�7���
L���*-̹3��D}ٻ�Y� ���/m�4�}�F� ��\ӕ�B�����y�d	�I`J�lc5�Щ���hlD���+c��8r��\����̷n�x�x�p�fM�p���jcp��0���h���VV���sP|;�U٬ڥ��������:�ͺǔۭ�J�a���\��h������;{.]<f�֭c��.��ɱ��p@��P+�>W���?-ҝN��iÖ�vFW���N�#H�B�Fa���Xŕ��ۀ� �-�NP�Z$�$����v����s�Ýn�G6�N��N�3Y�u��b�!�85���r�q�/�c3��6�6^4� ���v��paz��bvX6x��;h���1�im������M�=k���q�8��C��D�P�ٷ7��;X��������0�*t� �_���B�یz�9�k>j:�g!�n̻67�M�v;v��Uμ��+�nG!Ӟ�z�q˕���|�O[	��v����cO�%���ۉ�rm�0t��s���Żq��ؗ�tn�zn�}�X9��d�r�gm�V9��s�h�Ľ����u�\�+q������;�ywV5In#/��3��lZ� S �`�)u���{oX�<4����\�T���<E�$@(ۛ�����.�㝚����^�;r���><��6[yz��z�ntp�[��u�� 4��b�.�pw��Eՠ�^�oqvK����^N��7V�]�ֱ.���n{��S��\V$1N�nv6�wt�u��F���vN5��k�7���7�N��h��\:��pf�OY���О�x�ng�磭A�{��\��7e�v �
��Nyn���v8������9�s�pNGmO#���k��cuۜ����]� Cۮ2pK�r�nɺ-��m���u�sn�5��<8�:wk�=7'u�d�%C��f6���mm�kF����3�5�=�Og����5ع��$�V����A�];p����l�n�6�l�\ܖƧ�x��n�y���:S0g���]�7qr)���׷//Y�vC;!	��^8�7��\쬳c8<͇��WG;���fݱ�#���]d3��^y.�NS���X!פ�b�A"��]��'l�d����/o�c�Q�s���^Z�g�U��#]�x�,����۷t�q���:��v��1��`�㎝��X��n��p�nwc�;t�؎�#�/���ۗ�lۜ��F%�h���гeC��E���.��۶;tݎ�ݫF��l��;��d�%���ɖ]#���-����r�]�������Gv�ͧ�ƹ�wP��]v7gmGVR����·A��v�XwTnζ�us�8m=qƖ�&p�xKa�1�x�V��۝um�ɞCZ0����;t�ݠz���)l������ý.����79�,m����s\5%���޴u77n����;�n4�pף��tpp\���[�Gkr-{q^3; ;���1����4x�h�d6��ރ�8y����s`��s�%�ݮ`��*T�*�D")�ɚ<���ڿz���_���l9;%^�g�&c�j�Oh�U��	�K��d������X�@k�~��E[��b�"��~n�=�Y*�j�׋i�$[uz���2J�Gk�eh^n՟���`�1�48\P0mz7�����+<�-8%�=f�E��JV��5d�Z�|�邎&��-�JK3�>o&�W��W��*ל��p�=��AT^{қ�� ���㜄&Y��
�ws��K/m�t���vM[��e�>��e

�˦۠[lF*�
�k׏��u�$��9�U�h?)*�S�ʯ��Q�y�X��jv�Y]��*���>�C�9]�%���ͭ��2��KUpo��Hu6�Q4"�����_r�������>����G��1RK}Xr�8�m���qt��s���;����*#H�Rx���+��Ҭc��Y�g��S�c�&������0,�ݣ���tڍ�@�5Hv����s �c���M��v,8�Qw���b�0}L}7��߷�޺����7L0���<+�����iW{�*X�s�w�M,r�(�=��AV7�rNQeQ*R�
M��"P�Wa*U�R��&^|�8M��iY���מ"*�q�}��{Y�o99B�"��qm�"�-ͭ6��]�9�Z��Y�pEgt�5-�u�� k����;	�. ����ޤ>�*��z���>�Ea�o���U��n˝z�cՂ��Ymc��C�Β�NGU슍%��B��RWv3���W�:f_��o���ͧ����~�n����vV�k~w�hє_���p4']� TY^�\�*#���V ��^l��F"Tێ;jŴͱ.���e�{�z�{:��Y��3Ċ>�0T�4���sc:X���2��Χf& �*�7�ֻ�k�˝:�=��:��q!�ܧ�[�"��S) ����R�(���s=�y|fz���6м�=���4��#��.Nܹ^뒡�^�T�.����Ѣ*�-�[��U��ez{9��hFs�+��$�+$V8���m�1	�&���ksuu���a7^����q�V%��`�@,�%�5�x1s0ߔꕬ��E*�Wu*�w'V>��:�T�u�OG~p�y�`X�����t=��M�ĳѾ
��AMJ�KM\�6iLr&����ZY��?e�&_s;l�"�B�7��<C�}'�bE,���d�E��A�
��X��G���`�V;ѩ��a0)�uv��)��ǰ���<5��¶��U���c�d)*b����#+�I�i��,��㫨���6z��@�k@뭝�XhK6bՁH/��<�En�n���fFz�2�]��ΤQU���d��F���]"��4�eח���*5DU]WZ��acr�(@:N��n������Ǘ���m��u��S��	�m�&]g�|FV+�Z���n�):�
����ʂW���gT�_J϶����j�M:�%�-�j�KM�;�s�f�.m��-�E1����9�)_��e?g���Ⱦ�-�|%P�5�F�����.�asmGm�^�5�����N&��ݐ-ڼ�d)��5�v��tv�띙�A�t\�`��*���T�8�)S����w����-*�綔��˟;���U���4��s2�'ޕ�yY��1�c�* *;�g�;��yPp���Y��I*͒�X
$�O������\�0eS�uG��w{}�_}Z��x�ν�K�D-4��ҥ^��>sY���n�O���j�푙�o�E���>�U�i�*�8�'��k�nQ��X�E�8k��}��q�o�N��f��	�ʶ-W�⥧���(��n�V� fC��)p$2a�[�׃z�A߳�Y��� mp�GM/C*�;���<��	f��͊5
Ҫ+}�:���֘��7�&iڈK=raa������AwJ-�s�p:�I1�ˤ�ĳ���r�4��B��yco>�zX{�-oiҝ�7�oYǋ��(��{�nǱک3pS��S)�Y��+G�8D�P�Х����W�w��'ܓCW8�W�c�F���oY'zu3c�Y)�X���� �iߒ7��V�#
���羦):��i\��n�tȪ7GDQۦ�Y�h$�ݷq���ҝ�M���v�p;tV��+�ꔴ��Y*�"?yp��*#VB�n��Lpa�o�W\��M
�Z�Z��3��@��/�������F�VN���}�!�*��F*H��L a��/��!�G9�Ҿ���Q��yڸ�h��.�I������.�GV*�C���V�#�����f�CKA�ë�&Ǔ!�I;%&�qZ$ڽ,�3��9�����^�bBo���7\���\*�V��Nӄ��5�>�z�T�v�´Tf�0<��j{}�D)V���k�T�i�/P���>� d��uN�4��x�!�q>M~ ��-�C�ޫ�2�*i����1�,�{��Ղɿ�u��}^Z1r����-�؊�i0�n��?s�)
�N����]�?�v挱��o�睸_��\�*Y�52@���T{ީ2������ߘ(/��A޲�if��	߅j�u^M�̋�e*2m� K��4U]����i��d��ⴷ5#��H��֤A�}0�#R��{+jIKk��F�B�M��5�86촽�S���k��׀���я5ю7P��֝L��n�Ynr�1�쩔!�]���.N�v=K�ov�Ǒ�ۗH�a�`��Q�{[\m�f�c��M�l@ۘ���u��rQf}<u�nw7n�kv�q���U��g���hv���S�ll<���\�Kg[a��ړ[i��ۛ 1��u<���cc���#u��y؎ݦ�狎]�GVݻL��ƌp����Y�t�r����m�f�ߟ���*�����c��uK�`�6��X�"4��^��S/�jD�Ժ�Yn��Z��c��Dp�)�;���u��7ic���<$<(���׍-<k;�Ρ����<$P@KFw:����*#���ξں�~B��()觞��brxIы�;�>f�<%�醨6�d �WW�L:����J_oJ��*ΑQ�zU���?��V+���j�z�������$!��ik�`�s$�m�$3|.��A9��}�TZ�sm��|~
��A�:Ȫ����F��Δ�3�_^�����:)�qjf]�]u_+��>W;���\��r_QE]�$nQ)$J�6$g.J�*�}| Y���R�U��qo���9�>�.��b����������������|Ъ�� zCמ��/v����`[:Y��!D���E�u�Ϥ9��붮2�]~�v��7b��KL�5$Rm~�i��s��߼b����[���5�ەy�����f��f����X�R$xLS�V�;^��� Ə���F(̬���"	LK�oN��&�5����J��B�f4�菆4��H��gD𭤯1�"5��&���6	�O��5��Su�[��}�SѪy>}3&�Ǣ]��^ވ����k��T��r?^x��3���
��ڷP!Ϝ�)�/��]Ɵ�1���:��D5*n�I&o�R�O2ث�;�� r�l��^w�|y���5���ClL��>�ח�����g�y^�U�M1��3\�y�Ѫ��Dm�K^���}#��Jq�Z,
mR�$�oD�*ڱa�i����e�=�~C�+���nj��W�ks(^)�[8A-bh2Bv�E/O�i4�i5~M �gO���ս�{O��v9+����N��S��"� G�� J��]�y�<�+_�ا�9�쳏�l�m�h�{o��OT�˜i��8뤷�sz��k�ױ��	m���g��[��a��LANE8p��v���Rnoa,|O�^*�z��|W�����!q��y��'#�@�n�ʙ���:�j�'���t����E��������2ٞ3{��<,0pVL�Џ�6h��JC���v<�u�^�*Pd����F��Y�]b���sJ@%��/kE`�TV��(֑��?I2�Z4l��#�y��Z�u�u�Ru�gEwvb���%\�uÓ���{Ze{5�-h��Y^Xk�e�bUf���{2����'v�������&�8�¼���U�y�.��g�j۠�ht�uj�����˜�a5poz�H������[nG���\���2G�⹙@g��+龼<.��(i���h*W�K�*Uf*��J�`�Y)��Y��]�̫��5*�	&��Est�)�� U&�]�����^��y1)����]Њ��|ki��Y_X�Y"����ƽ�Q�XW����c7��65�*U5t{,d%�x�'�	_�N9J��v���ڒ�ͱ���uک����Mĝe6�p���P��՟�h�:O�7/�jY3��RG��'w�����޲��3�{�>;y��NjxN��{%L:����x�m&�z7�W��h���jɥ�ۭ7{칏���yH�:���m�3ܶ��w���s%����N}q�{5�GBU�5�5��_5�V�o���T�Y�.o��9�nm׹�+h.uK�P���w��2W�&���}b����o��s�D`�zK�~���Α:�g=�A��Z�����ގAoHJ�^{���s�n�)��y�]���U�#���� � (�->�}3�z���
��n�v׭��S�w�u�e{t����C`��h��>���a�*Q�n���Z���e�?^L�U:��W[Mv�.�l����T�d7�x3z��W��+�򿵣�.����G�7v�v���S>�g{���s�SݭG��z�{Xb�j�{���o�d*��&����w������1j�I׻/$�/���
��@E���X i݉9���lu�h]������J�X�Lm:"ڤ�U*��	W������[��}�Ƽ�a�R�/7�3=�ᑪE�{ˉ��H&�a��>"�Ո{�C�]o��:x�R4��� ��-����$u7�t1՟Jm�$b�ܣ b�ړ�X��ӕ�v���`���>��Ho�T��v�=�W��)Q�^�&�֎xӌ��v�9J*J�"J�ods�W㘋g6��f������{i�B��ofz�F(q�V���m��^M��]8�|S��]4�g���ѧ+tu�E+3���� Œu!?O�FF��K67�v��� :7w�g�r���VԊI멶͋&��	����pl��ؖPwX�*���7^����B� 4P7Y*�-=�ܳ�fʽ�{����C7]:��خy�4���t	�x\���1�]�*�7��ȫ���wX{UA���F��lk����쥰5�T��o�"�
��F��Xv�����ّ&5V�7��Ǻެ̴5���w��h�[ލ��@��_=���>�ݢ���f�sh�55QH������/1H̸�����m�n�]��n�M"؋5�C��u�{r�����.灭��}9��ے6�ݏ�+���a�ru��N�*f��`����6.8��=�ׇ$N�����:�ܛ�i�b��3�`ݺ��m�lA��1��%�cX��ݞ���!,�ư���z8�Tb�p�D�������:���i�ƹ'�V|�Ʌk�����cd�4����7k͗���yw8��^��U��S�礙�O���0m���������>�~����G�_g:cVU�oK��̾�&nFnӄ�xf`�sM�qCh���.ㄨ��������|�mmD��{���~���<�F�� �O�Y�Ky����*�=�Q�V2qJ�zP�Vk_M~������"���m>['�`��:�8F�q�w��7b�y{z�����g]
z�q7gS *;������`�y���U������O�L
����U)I�ٻ��y�`;��N�A+s:ĺ�^�q�m��PB_����E^�r���Ⱦ�+{��aak�]X�/a���q5�qiX�a-hV��o�2�2�w���j|4��L���/�l.����ӕ]��������CK��yU��y#mO���4W�|G���߅�H���F)c"i�����k�u��#�vM�'O@�v�����^�zi�`Z-1��5�4� &�N�r������y��SW-륤2�$��G�v>�-Os�S��d&��5�u�7`r��M|�]�i?[@"lq�V��8nl�7�m���2�`4��������V[��䥌yF�/-ҷf�� �j^��m>��>8٧�p��]h����>��idm�W�̾�Y���ʵvp�n�@Dy�ǌ�������z�=��{ܻ;I�B3���Q%�� ,�%��=2Vs�<�+՞��JLӲ�e�g���]c�\��*H�z��:��ڙ�m�uJWy:n��3�+��q�c�퇥�F�X���&^i�rk�g�xxw!��S�D�`���}J(�M�30|�D��k>�]�i�<�����z?�u������d��z��t�ks(���F��t��ޅ�eC^��C3Y�S�o�.m���i�&$�����Q�����76��d�Os{���!��ia4�(�u���M��cAEmns��I^:=�.�ԕ�l�c�z�]!�� J�������odnOf�<�a��b��1M`\)
"�����OT�#zn�/(VU�l�{�K�q�]��s��6+j��������d���u)^��T�OH9��Fa�|��ȀäCռo�L�]e��+�����	�iu>�^��V��S-�AXJ��eʱ��S=��T!�j�*�^�M�_6�'~}��G���,�ת��*%pLl���@r��]R��*��\;2����qZ�D�c2c#CwB��}7k�Z��xkm���n|�R�[����(��Okr��ٻ���,���B��1����f7��N���`ޱ��"��u��j�(��\kE��*���W
����bP�qx��6}R��=��:�6�1���3A�]������,�����v�7�"��k�m��b�w�GC���b	�jR���{œ�����Пs��ݹ��n����	r����1	�����J����
�/.nvU���f�e�:��e=��
��5X�70�9��]��tj����w=3��n�[�[�gi�铺�Ece�5����)�&��KEm�r��Gݸ@oywǺ�����T	)�fֽD��(!;A�>�6D+{�i*�5�*�k����&������ɼ�d�)�#i��Shr����W�3�n�x�0p���x�Bm�_���9S�6}t���NG�.���U�T� �8:���D�^[�&�hդL���e,�;��}fo]<פ,�G��<�[�!��%���v7I�u�n�[-�s���ʕ����QLMo#�{M�=���𮊅�m�2�wW��s;�{ϥ��um�!�W�g�Y�x����@�Q�Ԛ.��B�z>+LѶU.�]B'�SY%
�;��9t�
��3�T��{Q�S-Nۤĭ�j����|�q۸���+�?}7{�r�f2 ~EP3�ҷlK�
��~��T���t�tKT�u�nf�׶����ժ��ߌ�zk�k�>�ژD>�O`���ys��A��h�9V�ej�Az��P��0`��+�k�W;vID�nʕ���P&HE3u�Mx6�����t�>�B��U���fL�.u(�ҍB��}�VkƩXǜ�0xV�֦�/���z���;��Sc�ݜ]X��$�gu�3�r<;M�
���ѻ��ǵ��v�96
����I�7���뫛al]������V��IF�J�����ܙ"���3٣�z�_�
���5��x֓4��]/x��brA�ZͳL�^�`�?:�X֎��}S�zf]^����)�*tޢ��83<ӥr���>g�׏o�!�����׼����#|w=�o���iN�!���ٕʘ��?���qɦ�<~vky�<����wQ����r�w���z�?	����j�I*��~��%�X�IR�x��ȳ�k��̉���o=2�^�}ta��+(ֶ���}j�|8D��O�jXd��a�;]I���q=G��w���LV��z�����x�H6iA�<}� ц�����k7�36�+�c�������K�x�|�	볭w�*�m��y��˦���=�\��+���g��ǃ��<'�kD��]�NF��C���];��������r���ֿ����>�~��P�� اôu�8���Ez�]�b.�8�7vCς����x�Y9�Ѷ��M	������b�#��~{��on��Z��+��szO]�EBOyG���-ԡKn�\iB�Nv���l��Ɠu���~�Na�t�_��d(��KhR	U�����Ť������	'�n��.Kd�9�.Oa�}G��0�f�P��
��J��`� oBJ�/y�֋>z�;��#dMT�$�N�"�n�t�x�{��c���:��;
����ǯ_��}sG��+e԰j�k���㙡Y��<��b��� �gtQ.x*��s���/��	t�u���b{�ҝ"�D�$\����A��,��܆Y���U1J��z��'e����Ե�]\��hC:���N�b�KE!e+��;sͥ�d7�
���+�I{���HxpVk�9RXϔ�R�<�6�髡Pg"w}��[�>��lh� ��׏��wsu�$2	�A\���A�aj�S"�4����q�۶��tkq�9W����|�s��骹k�\��qso[v�U�EUq��(:|'j����7%�cj�K�(!ٞ���/U��<��Onʻds��ڷ[K�ŵ�C��� ���8�WrEv��<�ݫ�D�*�2��8� �m��4��s�����	�{=��ۮ��<A�B��zx5$Y^ݶ��`�tcG\΃���s�x���Ԯss�	������1�V.:�H<�j,�����n:�)6���΀cQ;m"�mk���N�u�f�ݳ3Y�-۝.�\g�Z�Pnds�i�6m��K{�߯����8Pl]���V��u�L{�s�����*l�Y��j�uh�Ϟ]]h�j��v�ȾC�QU�e=���Yn�qs�
(�
Yi��c�n�����*a�2�W_\�/�z�.��/�ߎLh2B<���N�j�8OZ��ʘ�F��x��~�"T��~6�f�nјlM�G��P�����Yi��O˚����;��G,VY�y7=�_V�z�4!o��>u�Ą;��}V}��9P9l�����գ�ʱ@.����S] X�-WCh�;m}�k�D�?���qߋ������8�Ȫ5��|}=�JG���\WY��ra0�u2
�T�hgs8iֻ.`��Oy~��t�BL��`K�#
���;���u)�~��*SȽO�[���z��^����R�v�u��z��64ԀHب��� ���k�2�*�+�['����`��^6q���L���IM�nz�S��8����} E�ʪ����1�&�����*�R��oq���փ齙u��:�K4ͱCe/�U=S�i!�ˑ��������)w���i{Y��1��^q���>o�M6�5R��#^���K�
u�F�{��hgpt�ѴC��k��M[6'��u�����h�v�aE�ެ���*w��w�HǢ��W-�J��!��嗼}V/��,߮��T�z�*q7괍�v=U��<���%lR?v��P�?{��ȷ;�N�dr�Vλ��k-��XX��K4�ul��{�	��)�Km��^�kͨ�M�r�|x8V�����V5M�{W�P�s�ʴ-(G�c[gm�v:�~�c�(����:�חԿb�W>lx�*�I��g}&?�'�x���?�L����/�k�Ӭ[�F�,�qR��Y�����yM[^w������A�rQ�U�m�r��<O�-r�#��+G^]��r��vGn;<s�:��ubK)�p�=u7=�2�l�\~��^5|�
b�	򬚬�Ezb�����Ӛ��۫fWDa�v��TD��F�xf��oƁ��ɷ2; �7]�� ���KS��=�]�/+~��ۜ�ue�P�H;�w�������v{�(&��1?H3ZzOX������N�!�[�,����*�W�HRH���Z> ȩ_�r��*.^���zhܫ��߷��6P�3v�q�Dצ�ik׎m�~��{�־j��ĸ�^b;����8�CO��Q��[\��m�]W�[A`:^wʎ2g+<}�E�1��ޏfz�*�F��C2@,%�Ϸ{�-	ի��+=s�NT��EP!x/q���#���J�����yC.U�1М����zB��=�<}�!�?mu�0�����(�g2)�3�r�Y���oJ
�ʭu��zs��䲂~Z'�/��y/�D��4�g���_bo��g2���)��\�PC��_]Rqۮ�݉�s�*�f9��ϛCgs�y�εmqDE0ͪT�0OeF�]�*>�ʕt�#�eJ*/���p�$�G�8OW)H�%�^VA�ھ��gQB���^i=}�1�tv��KV�H�m�D���䜯 �ʿvm!(�Fr�^dϱ!HW�J���9Lo� g�V��7*4O�zu���U�ʕ�	�v^PB<t"Wł&���գg�;��	�u`ҫD��{���.���f��@�W�Z��﹚מյ��ʱ��ᔲ7㎢�����<v��AX��A�ǫ9 |���lQ��l��6�mU�f{���ιB�&���<��<r�����޼\� 	�r����gU�5��]�I��w9_�o�uZ;B6r�#G+��]e�bM�V����dr�[�Vޞ�%�՗��[��{���d����5�}�ً���(Q�'b�j�,��!.0)�#����/ ����'|��Py���=��z
K��t>��_��dN�%��g��>WB��hڞ��.�k0nZ$��v��g��vi�0�m8�Ϛ��g�ߢ����������j�����c���V���]�<�;ޱ�^[Lt#UyF����{P&{�;�~6�eb�&��}��U��q�L��5 �v�f��EW���⢴h��sM��O�97��:M_�  Me7�kI��¨g�w�P\���׉���D%B�����ӛW�G<��s��n�b��B�{}K֨<�i��uu�f*��x�-���WOK]��v��;�w8[�Lkk\��J슧�m�L�7o^f-�4U���Ҽ9N���P�񝮲�Q��W�x��xP^>IS\{7��佗��+C؟�cjݜ�Ȝ(YIRڶ��X�;�x��6�t��w�
���N�}����0]1�;�ul�|������϶�)P��)�7Vo|�j�aT��>o�Y�B�l4lm�'�vqED��n��.�4������ղ��S7j���k7vm���q�ph��i���1�Hfq����lp�'��s=�d��ٯ/[c[��c;�u��v.���(�i4�kP#K��� {c	չ�m�d.�;;�ѓ�����e;<� �s� ܂�7d��l���,:�\&�o�U�]�$Psl�hwV;t��v�j;h�.1[<�ۭ�{u�ӛ{m�n�!a�d6媸�N�s���6n�۵u�=��; m%�ǹ��q��qX�㣞v�=Q��`��B9]�3�f��k>�`�[���;��N)wi�oAt둶��$��):�J�Ȥ�v�]�=��q������?w�"��*��:��M��ݛ|��P�W]s!��\3���Т�I����k������^p�G����SA����4�Mw�J �kj�$� ��x���O3�u�}�ә��ɺ�c��C�k�n�l��ѧI��i������逥���fU �Z��^��^�{c:�W8n�kK���8�^�燣�\�̩4�"n|�u�]�<+�6�	�d��m��g%�~A�����YT��f�v�r!��*P��3�Q���O>�pd�*Q�M֢��������
p��)|�\c�**eX���.�[筹��,5���L�Ѵt+���6,�M�w�Fo���ȩ$p�SY�}}ꁚ1�}��йdֆ�[�c�A�����F(���tf�;��P�\e��sϷ/A�t�ؐ�z�]ܡUd�|�vS����"�,��g�rJ��9F\����X�٬�/����%�.�����ޥR��eSzk~㊸�x����G��)SD�<<i(t=�}���鸶���+J�6��3��l +nw�������7G�Du
	LX�sy�å���)g�K58=u��ʹ��Sx�����Z��]/�x���r~�Eݹ�jG�·V{�{��{X�,�.���g�M9)e�FX����F'�G�z_&��]H���}�Jά�<��3f��u,O	t)L>��׵^s��U۷�W$��1�`"�"[NXZ(����l�r�yu�xE��jʹ��n�¥�HD"���z��b`����e{�ԞדC���f|�����؝3�n��BA0�Y��E�+=�Jz��Bz�fH]���.�w\��^R�m���Y����?[E�=��߂��S/8�y����]k͋J�('J8�� �a���lg�����[����۵�;}�[bm���HӲ�I_}r�Z\MZ��k����
4���6�y�o���BR���q<Q�@D���o����9��w�m��� L&�+�[�+_�B��������A��e�uʰۋ��Vy{7�N�����[U��ZZ�"���uM5t����+��&W��+�KdVƘ�-�'9u�.秭��ߜՂ3{��ŏ/*^�^s�kY���'B���ur�Tnzw���N�kɚ��9YL��u۾U�z�־�����K�u�i�dJ��lf̲Ը��j��z�;��J��Z�Γ�Jݺ߅$Z�`�}��ƨ�O�ۃT��.]q�fݨ��F�m�WZ�*�-�n����~r�MB���+8K���o�6�b�5+n�ld�g{а>�J�+�^׀�5Tr(,���-&�x�iwz��cJ�Q<������WPW�w��*�S��~��k��_KB�4�ZGyr[�d����e�@A��\z��/��U���^�����X�u��{n:j��m�R`&�6���-�W
AL�*c�\��۱¶yO�������Z��uβ��YZ�b[~�맰��y��cv#�z{�ʣp�L,�5���@5�&�z��w���$�*���t����u�Y	r�e�/ئܔ��(�����@+1�G°d�71�]�M��a��h�gx�H��vCp'��+�Y��0(�ҥ�_ ���Y�hr\sud$�9���Wx�g
��S�j�ty�ՈWdp��l����a��<����J�.��/���
�p���s��\�A{5w��'�YqL��0� ���ȃ���gt30@�b#�LY~wX����:�.������}�W$���Y5j����h��ojp��]������2�쭺t�֬��4t�M5I�*I�WW����:���79t���[j�*�K��I����Нq�i�S���ּÊv����̻������_�����H����+��=�-O<c�c�.�� � �N,�64:f$�L;��Q,�h�	7��,�⫮:�a��~��*C���\by��ulr�]�m�dW'�zZ+ͼ�g|�[�P�^�+�W#�LNR���sW���sY�Ҧw����7�x&������n�����:�c���)=�_���s�;�V�v|�޿e��}�g��hYZ��b��"�i�/���\���ۺ
��Ʊ�1D�G�_����a��։B�S��/�v��̱����k��!�t�-'M��n��
^�^��%\Kw�:z�Ϭ�g<Y��#X@�r��	��-^}��i
]���w������:#swz\��ҚھqxD��B��/��#�~�.q�I���6���<�p�Я{�nO[u��	��y�VY�<=�7��4WF����,�f�j�'o�zI�	hh�idgV�(VH7I�j,k�
�J��I�(�O,m�{��Mj�&wv�����w�r�>6�G���-Ry+��Qdv�Yef�;�,���)�^άV�T�/v��OI%"�����ߠ�&�	�J�W����L�|-]�Ż�nf��MԹW�	�}wCA}���4QܿL�1�|�m��d�7�A&V"�����	�]��\����k`�M�]���xQ3'wI$��ცt�;u���o7�e�I�k�)R"M�CN�;�����I8+ME�"�Mt9c�M��M�v{�v�+�R�s.�c���q��e���P�F��%�X�c䡅��klj}6�[ӌ;'n�[��Vn|jG(�����ߣɉ��¥g���>u�}[�ms�3/����UJ`ަ�N��p��Y�[��� �!��Z)]��[���5��['N��R��uwm����fVEƄ��Τ��Αwx��rOq��5j�0���ͩ��c&���k|�c�;o�(Z(�G�S���O5't��e��7,����!���'��Sx��,���7kCך�/Ξm�]?#Y�+=�%�{�� T�pw+�\�.1.0��������j�t�ё�V�6����p05�/yq���ֵ�9�Ngc�Ѷ��8�r��:%�k|�iP�:-s*?On���� c��>�/},�jV8�$���O�G�פ�S]��^�iu�\�VwQ[g;tؖ%.Y���);[qƬ:^�9a�2g���F���[�Ehe�2q�C����|�����]r۾o9!��{�	�u��c�8Y��\l��x�x���v�]�7��6L�M/Y�\��q�:�pq&Ӹ���U����6kN^���q�y�0k'/F�v�5�+������%���ɒ�m&�^��n�c"�AӠ�JD��H��av��1Θ�rx�V��Z'(�N.����uo+��z�f��ÈN�7��w�gv�8ݎu�x�[��x�{f�-�t� aw;aw&�g:v�C�#ל��+b�vu{n�E�1ѭ˽�H/y�V��;qӚ.Y�{^L>�Aɺ7NGdr�n�I�#ә ���mG��.��iK���띞"EK�Q4�����UR!�JE���
x� �PN�f��sN8�]�p��kY}��N<��:�z�Y�/�+�);�6�.n�\m�6�z�[����u��x��d]�۶y6�������m���O[�9:�+6�ך�Ȇqut l��W�Y�üK��/pӴ�G�����棶�]�qű��y�����7k��׫n���䳬��Zm�:LxA/O�m�[���׎�����nYx{�g��=w:��-��b9�)�-гWmm����=k��yuW��\�K�����Oq�N۬�n�i�:6ܑ�퇀wr��3��/>��Y�]��Pm�8��%P�s�0�C/o ��=�κ=]�#������:��6���>�V�swU������8Pw��m\��u�%ψ�W�w&�b8��[����O<t�.8�qőy��m�='���FG���:݄up����b�6�ǰ���8޵�o4��ֳ���k�Z�{ n�ܼ�ZD�S7�i�]��'��V��Op�WY�Rvh�n�r��í��]����]Q�`�n�f��9{��{�8{>ǃ�!�Yn�ۘ���c`�\���Og\�{^���n$絺*c�rdm��\u8<GK��(�y����+�u�Z-�����Kfo1�[��C6�݊K67)��8�m�2`�r�G��;l���q���aï=�$g��&����8қ5p-�6��u�۝��ݳK���s��"�x���.ػs�����+v-�=�a598:��hx6;����3[�az�=[��kZzmٻ$���Ac���MKs�vz�\݆�n
�'Gq��⹴e�ܦ�h���I����-��ɯ`&�Y� 2k;����q��뉧[�N(�k��Z��ׂ�s��f���qc&z;&���Aƹ��ޞ�tr�U�u�^�6��,���glw�}�������b�x�A��- Zl��l��G2-��N����I�B���:�Ǖ����f��j2k=/ܳ�{�^�����é:�. Q�4�w�ֺ���V�H(O!��A��X X�Iz}�����˺&��3������.�sV���1u4�B�^{o%5�wO��0��Ks&��鞨z���-kzkJ�n�c�U���������.��5�#�Wv���EP��JG��>���Ν�z2\�s�1�IݙB�.�AQ_U�=\ I�JE+��E��\dX�R�K��1�~>g���)ٵw��!eH0��m���ʗ��ck4;�o=��vbA���O����R)����s�[C���}��l�A�L��zS5��^ūa�V3Ӂ��Uզ�����y⤯U��GnI�5w��6�Ǽ:tJ��c���8�2Z\��yi�8�㒹���hy|Z�:�
�VӶ��]P�6L]ֳo�%{�Q�A����.D ����x+��h̵�>�v<��2��7c2ʅ���-��$��喭���5��h5�/	<�JQ{/^��r�����^�y0*��}��G>�H3
��z�r)g���N�M���U�,�ԝ|�gd͹�5ř�� �����iP�/�������l���ko��d��y]�g���.A�۫��"�����,{�N��J�Wm�ߘ�����QD<X˧���2Y�b�Y*����=̇__���N�U�ۗ����G	�%�����@�Lc�:���S)�DI�ټ��QL���S���"��n�OC�E���k;�=��Pn�e����k�)���,��z��K����=.��j{F�P�dTLt��͹��5v�K��ԩg���6���U/��lRy��ޏ�� �M|��U���.=�V��&�%��H�)�-4^�Ͷ�Es�e�QQ1�:���Y+1�����η�F�%�$��n�p���%�ޝ��.�=n
*���Au��_�����fv��뙳Řy�g���@��tD��x�1M�4D�W$�����u�]�L����}�/FB�.��j>��+�wf�'�d���l��/�V�ݝ酒��%!Y~����#u��i2�f�l�5��*�%��]�]ʕ��ޝ�C����X�z�(f�:�p�Ʒ�c�0���9�r�'�Vc�@VPH�l��Q���p��� S:/u��Y�&�^�f_Q�����ٞs)]N�d{�+Wu24�gV���4Y���A�_�؋)�}�ڸ%J>��ơ�s/|�t.ݾO�̿7�g��.�t7�y?v�o�����JN��LJZ6�4,��� �ܞ�w#�ܜ7sٮ�R����pУx��Ӭ$�^]��QX5����k�8�b}���|E�
�rl*(:0�9�q��ZK+�ع	�F�mѺ+]ntr	Շ�UaB�D"����'9oup���>l�{�s$~�1U*~�n���+��K�o�@l�yF=ܶ���zO)�T�,��+ 'e��~Z����q����i��c(�H� ��Y�d��{�\�Y���f�ZE�K�]�pKίxf_/7����z:�p��n����+)e���=%J=�Jg^{�Y��S�K�:ў�<x*��zo�m�9\�»)+;�RO5�\�+2�whV�%���+�����M:�{S�-�;���By�3s}�Sc}Y��\;�~��v���e���{���%��Oy���F���7�anٸI;3e�e�EV��ͬ�6N��f��k��L_b�Z1u*����O�-��Gqۿ��ꑚ'jޚX^�Ч��E��"���K=}�����b��'�e�,�k����t!�&��'NN��q��PŽ)��8)"@�	]o��:ˬ�����U�:���{Zq{�8�$d�:�(���Ȧ��³��۪zC���c/#\�s��ۧ���l�[I����U���]��z�Xm���:��R��O}�kf�b�����Bs=�阓B�GS_��)͐ۢ�ʱ@y(��������s�|�Ю~���}�>�#d@ۥ�7��V�5ŋ��������)��엋ǹ����e ���&à�u0Eѻ��r�k�2
���W�gw�Vb�E�iH˙����X�t�uƍ���L�}�ݣ8�F����e�HJ�)Zj�v�hS���U��73���sڱ��V�p\=�oe��}�=ZG�<��Q��ۗ�+-�x��w{���xc��$���n�Gj�P�M5��!�%Q�{�Vo�2v�2�f���V��K��z�K1 J� }b�2{�A�v�	�s�f��r�[�jc���O��T�c��Kܗ,�E��o��z�pH����5���E�����μ�X�|�޺��M-!ұ�b��T~>RP�E��6�����C���M��HR}�!��=s��WAs��꩝���l���!�GD�Y��<�6x��Ѷ�nK�3��j�ՍVk�.�b)ǐ��G��;�j��M�t�h-���xѓ$��X<n��@/Zr��c�@ꔸ�͸Dd���2dͼre�ٷn�sv�M��<j��zy�v�ۇ�=��:��g<m�c��>��9�b�n�H.y�[�5�ϓ�[�8LTWF�����]�6�Js�R:�qԚ�<�8��./?o�:��֚�U#MR�-Ӛo�s�PT�$3n��:�g�*U�~����^{��4Ly|��T�K��y�'�m�]���de�����w�'u�F���Z[+�,��-�T�A�ܡ�8]�I��t�m=�#0�:u��S�ł�{�V����B�NA֜�f��L����^�M�������Y�}��o��^!�	P�����V�M���Xk��?L���[���s��z;���:��|�$�i���G�S����'3��my�y�� ΢��ޔⴭ/ȹy��gW����o^� �KM�9�J�g]UR��`G\���vr$]�]�����K�)N(�WY!%wKǫ��$UkQ���[��*W����.��/N!�0k�.�7k�)�lZѱ[{j�2V��񺺲s;���+[01\��]u�e۱��IF��L�eX��:���}f-%��>�,���RX|���ƅJ�޷��]��y�k��DzEd��5�������*&��^�m�JH�MIKM��-�h^��>��7����3�^ƾ�*����a�`�6_��û❌
p�L���0ܛ�c`�luiVKc2�u:����+H����	����N�*h��5�c}~��W-|$|M��T}ք�2K�t{�۴��x�$�_x�z�{&���C�]�?�yX~�u��0M
�b�IG�`�ٽr�<\i��{N���Cr�J�T~���j�[ɲ�z�
�J�xFz�$��|�v��st�e��H�S&g6�A��{�Vd�K�;��m���~}B�s&e�~���G�vT��w���^��9�x��M�����i��$v+mX���Z�^�4{Wn\�6U���4�k�:��,:+�Y7�Ϙ�̨q�ub����^8�������Bأ������>�:N��XG���������:Ƕ�v��˷ct���b����!۸`-������0����Ҋ��z��;�f3䢈8]�s��;�N�,7�|���[����s�c4�!��W�:��EP&�ʵ��m���\���C�.�`P��d��j����H��d޾�a�԰��}�xT[2���V@���-h3��;$���L7���v�Kj�	Y�����!+�K�\���*N��~��st�+}ap}K;F���x�W�3�]���k�N�ΠViӸ;0�w]�so�m�@��'��]�w��ҴA��;�r�o^�����6�`��<�RtJIPmь��iji��ݪ��������@n�\�~��e$ޮ�x̻�R�������[�(m�o���	��4		0�MQA���N�M��U�� �#V8�!;9�o����є'%^����dswzb=9t��ޙV�nkH� ork��g�}D��M�i8K<uפ{^e������VL	��]O'9u�x�X P)�Y��-��H�}|{ˎg�T/�z��^�z�I�Z�.��{ϟ����L���D�����)��}��[^zU��H�h�U� ����5�JSk��vOw�Kʢ�b�yT9�K��z��qG^��e�xm�?Z��	�/��{k"H��I��y�'�T
��G�n	R���c��}Se�v�-L9QV���fe�y����p�I����/ܝ�w6p��1F��7w�d¥m�K�}:i�ܴ�[i�g�xz�TG_L	��=o*�}�z:{�~��b^�潾����T�. &켃3���8�5Z֘2��&�u�֞����n͋��@˩�M�4��ٹ��[%���#oN]3�}���8�RY���H�h��@�m������FU��N������w��z�kEY�/d�6������l���jX���1�"����v׳T�ڮTvZ�$�j�m��z�Q�!���K�	����-���\�:N�y��VJ"�%vOY���ʋ��IR����M*�j���_�~����k��+U��&U���}$���ߗ|0Qm���M:̼��趻���_����N��G������O���I�~&��@�F��=*O?�{z�;௥���VaM�e��*�M1��e���&s`�����ƞ>~E�D^:}X�P�&�{y׽퓘�y�����x����k:.%����
Jsqƣ�W�ۜV:A��h3���"��)%�:��˔������}/�j��!�/��$5��\���N�仝�Ȇ��x$��F�	��������W��Y]��bּ��f���y�g��ǧS��x9G�]m������݁�B�m��1:���5.���m���o���C�~.tH�Cr'�[�h;�>�<F6�K�t��k�NV�|�v�2��K.��$c��@?���؇c*Uƍ%�����n��j6N��v���];qˌ��ǋu�+��V¯Yk�&���a��\��.(�X���zn���P�8�;���q�iKې/{u�5��ri^U5��nZy��mW�Ŏ	�2�ݥ�*��r[��6xLvNz��]ga�he�8A�ܜp��i�;ft�u��Κ! ��غc�:NU����{;�Ŷ\��Hm������7,�W�]w>:x�8L۫�KŬB&fji{{�+�o��ϑ���+�]�S~7���W}�?��~���l�,0��Qm�}֥���kb-h#Tj��Z��roI��J����e=��w���k1�>�;|E+xw��U%����A��.:]���1^*Z���V��ƟsC���*^� ��r�n![h��7�Azv�#��&�++{���gWk/r����=�V�Ⱥv��x����צ�.�{i�2�])�	��lF�����{T����z=�GYE[k�n��'���`Z=*{3XJ�������v�`<���^�|/���]�[v���(,ڐO���g[j!�<����ӧ�{����O���wz���Dʕ���ށ �k?������l�O�,K��;�h�I��j2�n^�-պv��FV�Uv���UM<ǎ��_{���g֗�';�&x����O�{d���ow+}��Y��3������ٗ[9B�$��7K�n�~�E�ju�ٗ�����!��b<����t�)Ķ|�^�&�k��_��PZ��&�=�R9lcSڀF����n�t��@Vf�K��0��[��R�z$��㸸��Te����%on��P��I�B;X���:ܱ�N�a�hSm�r��z��[;���>���{ט�����ܭ�!�m�B'�{���T�Xs��e���;d�o���&�tuy�Q������;A����T�ߛr�W�4滊_E~�?M��,��:(�v�S/��;���F�o���V��"��W�WH��L&�($��e*}Z��g���U�ݽ�S�������vOT妍�(�?,��_gb���\7�N�;Ȋ�UE=z����'��O��b��b�k��øc`s����<&�s�s)������Z%����Y*��ח^O��I�!��-������a���=�����s�h�����e����k�m�w3�7�ק&V���o͖��n��m�죶�6X�Ot�c��p>wI��{�X�3��]z+���x���Jy�]0�oY���>���v:�c���s}Z�U�)#�	��$��L��ϝ���ti	��S��[��O\C�ꭂm�xI{�^Uw\ۇVL��.�H}�;�I�\���r�5��4�َ���hvAWh[j*��۴�1F��OQo������^��Ϭ|��0s�Ut���Lڽ�L�)4�N��c��v^+�q�T�mw!)���&e+�@����1ۡغ���cv��{�B*	Z�s��B���=��M���U��o�lL<�iU�i4��M�F�T2�>��:ur�,v�wKE�:�Jy��os��6�rn^��^��P�?X�3��z�;�,�՗���������wϣ��ʖ3����\jQ��Zrg�m��������b�:�*��c_(e`�˺��-�\$s�,���Sg2s�`�l�:����-�V����;������%�kT73aܳV��a��R�3��1Xr�l�������^����ĭW&����P��b����Y��n^�!�v6��[Fo.��#�gb��6�n��2iQ&ѣYRzO[7w/�f��D�ۣ�ɻ�����^)(}�?���X�9T�[�X�--��r>۫4��;�3L«,���3V�6�v�nv��aɕ�`Df���jvwS�%��wҏ=��a˰x@�Ĩң[<,����doԩl�M�<w2��T�^L|�bGћ�������9�Wʱ���i������D�ՏQ������E,�8�m<M<�k�9]�o4�Ǩn="'+8ָ�(��ńw:��2�.Ы8�&�my�]�WM��r��p\ڂ��)���f�w~�O������y��U�M�߫8�����}<z9��mv�ʔ'2ڧ�i�m�X�"u;l���]Y�����a�=�k�3{��\ʑ� �w�$���׺�;�@-�e�<�#�;ܐu��Վ�.@e4�A|��"ٞ۲��^�*;/;�"o.|���w����Q������'7<����=Oҕ��BإSQ���I�_�qF>4����/��Ѹҝp���ۂ�qv��@&UMTKT��;��)�ԪR���%���m���^ֽ���?~�Yͦ�k���=��¬��+�ߓ�K�:�T_���ƨ\*S�D QE���9I������zu yx��N�Ď�yxw���ѤԵ.p7�������׬ uz�e� y��͈m%pI��k�L�1r~Y;�<���}�����#�z�j��;{�n�&x��Jk.#�������������T�m�	T�l�5����n��{n��<�,��;�r���;��+fڅ�KP�1��ʱ�Vg�8cm�D��0l����yZZ_ga������(�2s�yuՕ�w]֫�|a��(�;���{����ӎ��mW�o&;�@A��Wb:�]�Wc�T���-�;�b���<}~��r�)���/�\���^��݄]��"3��`ɗF[~j4�!L�מ��i�Ǵ���n;'[���8���zMu\I��V/z�M]Z�v�w�߬~_����\%^�RG�u�Y0y��y;�k�a���j��i�hU��7io��#|�z�O/�0$�AQ��ڻ-��r��t����rT���ϡ�̛G�S�7q64��Y���8%�hyY+&����ha�R�R���r��0������A,E9�瘃��^۠�bw�9��n�~�+�Э#�ج����4�V����X��վ}��ɽrm︚"$�i
��JN`�̷���OS��ݳ�v�{���N���;	g>���L˓d�^�h?�����c���`5��]k��ص�x�>kk��4	��K�kJ�M =�ʫ�e�����;�+�&�dF��S�M���R�v}�����!���Yy���1K��̓|F�7�Vkm�	�6�CQk/Fl�9 �@��4'��Me���J#/[ݔ�b/L^͖����˥8�כ9���P��T _vG|�6vg<�ڵ��=�S��� ����$�ќ�'lnK��şf����<uԏEnxv������_8��0�c��!8D�'9��u�n��q�;`s�M��N7/wc��&��>Yad�cj�ް/Mͺ.�I���\��s��ۣ�n��dcqR�5�z^x��۷mű�O\ny�m��Xڄ(^*3�ѭ��a4�.7��F�9�-�v����{s�}R��+���N��y��u�ڪ������V���?{����]����̹��B�r�vov!a�����[�>ov�nE��;T*]��;}S��z�h:E�R�o����M�:>�Lk=�|xk^�?-�lu���~ǢS�h.�eyTH�ޕ�$��ޮA{x8]�(�ւ�IdJ���������XY�.�G;���K��Dc��s�B�'�xM~�|��x���S\�.j�ݯ۶�~u��3>�b�ƽ��N���ֳ��>鉏L<1��&�	�J<�b����l�?S{�E�+/1��ch"�v�+��N�"h�|F�m�~;VЧ�f��WDߝ�'��m˄��s�-�W}j��Ƴҭ�2�%u�{���ĕ�uZ�@��&���rt��9���٧:M���bM\G]M�hx7 ��R�	�4��V�oO���>��	���
����;8*����w�񼞋�n�N����:H��a�ԞՌ���X��<�F��.K�Uz�"n»�:�fi�w��Y{��[�������pBMnJѣv��-��K̗V���xx��>R�՞U��[�p��1�[�ہ�I�myyp"����9���O��L�s��P��%y���/+�T�M�Ѡe&-iT7����3xg��JUg��:ī鞗v�>�}b��;Cxio���]�<,[WJ֞�&��=Z�[)*	�	5�w�|�cy��۸'{��t����B�O@6�m��w��o+no(�PJR�~}@��eؽ-'�^�P������\j��O�S�k��x��}8X�M�h�a�a�=����zR�C��}���K��#��M�Qm�V���WH$�Z`�X-qݮ�0��:|�bz7'���U��p�[;�k��H2�!�~e ����x���&����E��^�\���^�.(���ED�]	�9�gW �)/e���˹s�qq@�ŋ˾*t�G	+;�k��H�g���^!z����t2+�rE�+���{�q->����ק}t禧����o[�u�j��	�YUԓn��b�p ���?m�o������ھ���ԣ��~;Ӏʄ���>�a��y�7Fv6ݬM������g|��@�}�C;������`���X�e@,V�RQ�+y�����ؖ��S*X��z{o�.�X�x��%J!H�"h���Mڴ���B�;��=�]�3@�_��y��meN֪՟q�Sk�|��rkn���d�����<ǲ��U��lZ�z�HBF:�IB� \k�y�{q~��M���/��9�~��3<�ܡ�cig��0#Uu�8Lթ��>����|�]��ʩ��}��r��1����7-:Rr�9ge����	�8�nu������8&��*R��.Oz�^_���-ɦ�(M����ĻM�Ň޶.=��i�	O��;�|.��nF�����8���Gl��I�k)�_
��R�ǆw��h��'oe��Q�a����б皑 W_��/�*4�{�o�>�bU�R�)(�%��G� 6pw���)r]ג׏�>�����fZ<��]I�qu�=;ϯ.�Z�a^�d�6�2е(/R�7�E PS�E4�&���U�r�Uy|�7�4�ÏqM�ޮ�B�w�ņ��[����e�{�ul�Ix�{��sv6���ݡ`1�2Et�-:y7��ur�Qn��Ƭ=[kNe���cA�������4���\�Ӛ���G9ѹ2-����"�*nT�!(�۾'��t���S|��x�'��RyNj�A"�^��v���>�Yp���ҽ|���/�����K�z��b`4��|���C�x����S�#eP`�U"Nͅ��ڃ�ƞnx�vSK��\-�5���Ѹ*�	7�{Ļ�^*]Y��e���Dov]�����2ǣ���y�y''F�P֯���J8��B�ۭp��f�3�d�lk����%��O�4ڥ71��zLC���P�z�e�b���
~�Vy�Y��u'M���*V&Q��L�e K�����n�?z��X݅�'o���k�&�ٹL��ŻYt.�D��q��f�������:S����m6�]�^�O<N�2I�u���lM�b��Ҏ(�x�����Oq����L��+ɾ&������< ̢�}Ǜ�ٿ6�]H�KV��Nf��lRkާfnp�So��R�3����Bl����Z�m�~�k0��WH���S���>�{pDG��߅A~���K{^��J{o֫�}���\��7.��RU��t�MQ$�W��.��u+yj9�Aγ\ɠ�C�ВގY��������Ly�N�c�*� 2���*�u�x��ӻp��q��My��{<���#k��޲��7ˇ}�l��'ui�짲��ۚk�)pOv�����.�5y{m��\�}�+��]��ԏ�U�V�k�:}��xzrk�vl���$h��>q������]�m�����Kar���i�1�Sq�<�a�j2�N�33�����c9���g�6�6狵�v6U�ҽ4�ݧ��4[�j�H/+���v�nr�4���neg�f�T"j�R:��EL��{�^��/�۔�᫕�~�{)\]�[B�y�k�O��
�V�s����ԝ߽��,���h�m�n,`ۮ�N�����3Ǝ��K��9�t�r�5Pb�Я0����*z���.�෎����G�
k=�8��7��x�ѐ��J�%��7�b���z�N��
4�Nln{�Sj�~\�[o�VwA��^���M��H����	w,޾w��-4ۢHlQ4YM�Z-�]����ܵ�ӝ�����~�=���ȶ���2�޾F���w�g���L����r�B=P��gz6m�mN��H�T(3�e{�=KǙ^����;}����:��	����c���/��.���{f��Qa]~���d��aӻ�:�W�=�#�EX��@����t��.�=��m�Σ�9ޤ�H^:z����ۦ�LT�j�n��5����RtM��n�ZΙe�d&�w/o���1�{����z���OK�>�G��~�hk���w�v'�A�K"�a$�I�ƙ^PR�<���N{��B^�O<��������ܚa�c"��z�5]l��,=}Nm����y�L��wY��ѩOO
Ղ��duΆ�ϳB����a��oh�լy��
v�}��^g��g�3t�/���v���ů���Z�d���;�\~��^y7P�m��	f�U��S\�	�[�w�%��Y��]�[�و��G{5�_��n���J㋆{\�;:��9�`��
����^�`���~DO��c�����k�ֽ��u8S��N���b(�%%�'� 1r���tܕl�&W����Y"գI]�%1PZ���Ჟ�N�v��L5�Z7[�V��dP��כ��r�@l�_;��P�ϛ���3_ٶ�ѹ���{ٓs�����:ܿE~mX��{b�M�lke4������Z�]<��P-��B�A�Knz�i��<��[��f��<�Vհ�s��]���a�W{8W}G���z�@Wp�u�)⊝�R��%-XUE:�r��m�[@o�kH�y������,q���N�s��4��7c����yv3>�����m���ep��{�����$��t����ٮ`�/���7i=�ݔ�U�s����N����F����g*��X���G�F��ւ}Ý�ZOM��豖m{+x����KF�Ι�q�G��]����X��$���<z�v�b�>��(�WS5�g�u�2�������v�D�٩Zi����KZ9%^[!�;=~����YK��z}��A���.�N`(�bw�8�k�b��-��2\ȸ$d�9<(@af���SI4'�yTA��w/t�	Zv�{9��|ja��Z�4ֻ���oķI�}�W7�>=[<�k�:c�T��ڮ�'a"�*�IP�[ho��!=�������۶�]vLXpm���� �_�
�Tji���}�&s��z���{w�&��+��^5W�q���k:ᚮRc���A�7u�bߵ���VB[Z��bk��EE�{���9ݏ/'aK{���Ṝ(����L��;�#��2��m�ޞ���N��Z�`������"��%���P��ajr��Z�׽�5���n����N]���s��>�o��>�J���EZ{�W�����3V���|���zc�+a� �G�?���M{ն�T�����|��*n��M:E^��~F�ėnE�.x�r�Y�h4�h�	�hg0 ���dĤ��::����r�^XJ��q��댳�V-�֗�����ڜ�'.w�1��R����Ã9��'��N-�<C��P���	(US����n\��۞�@ٛ�oH���8O���ɬz=ޑ�<�y�>�J���<�Ħe�7��/!c�d�*�W6�t[m��9n�{h�ꙓ�#`=�v�/f���lI��l�qm[�߾��t��ix�.�{K}L]���Ԧb5��J��5\xX�s��qz�T���"�j�nw���y��ŋ/�ai��-�t貛7�+X�lu���Q���U����hp�\�)�����n�M�l�1����=U?k�~�Z +���:v����sp|�e��T�A�O,��C!����l���}��pL��o�^rh6�-����53-�rx��{��{V:�R��V8ZA1��Yި��85���|��V1�R���?Z5	���&�������\#*�m\��lA�������o��L7cE�סP�e@*Ud݇ �{��%Ǉ�ʮ9�x]+oW��k���K��øw	�|$�&x%�q�U��'�}�%M����[X��Z�����ˬy&-���Ѩm���ب��ީ.�9G�A�Ck���	���X���U���6�u�o6�"?��e�+�x=YZ3�0���V8X�#9�ǻY�Co��� \qX�h��7E�.]$('���gr����ݓ���/8&VCz/6�Cht�}�e��wiʆl,���vS<�mmq�T�p\FP���ʺ���G�݆
���2X�&�::�f�!lj�Վw.�VT��kj���å�#�ѷ�.�Z����X�V5wnX� e��
m���C���U�0�	u� v�ξ��K�Gg.f	bB]���G8y����H���uu�"&��:*X����l=�O��24�f���l)��d���aMܳFc�]n�{ϙ����U�E�_�l�\�bw.�N+'��Ֆ��L#R-X���զh�V �íRr���к�8������t�z�V�>�f�%&e-�s�㵕�$��u%{�b��_7]{�q��������vx��S�,�4U�u����:u?�����#׵'�#ԉ����5,��&��Y��n���~�r�e�-��n�+�8覣�Y�Y�}H�n�Mc0���+�	RE�t�s{���iLڝ��ٛtvw`wMv��-\�J_Y�*oV��
)���(*���ݱ]�k�7S��5Նt�p;���,����4�B�'���.!����gY��v�+��i{}�������	�:$�{kʳV��z��\\��\��]�czv�R����=8m�eёq��t4���[��1�0n�7�E��R4�,�o�wб��cp�z�`��/Ocv�x�M�է�Wl�w��b|=m�3�(ݍm�=�k���#�j�봲̸�R��ևMgXb����1��va�g��;N�h�Y���;��Ю	p	X�ۖ���g�݂6�����m�$�\�q��v ������X툮�p��Y����ă�֐t���b�8s�J��
��B�zq�}o����nc$��g7l�U1����g��mˏ�x��9�g��c���r�.#<�m�����rniM\��{iMk�����������!���X�,���l#^�;ځ��N9�������������v��y�kj�ܼv9�����F��̱�䮴%�xu�F:�N�;ϒ�w^.$wF���ޅ�;�m�XnƩ�豾.���y�ka��y�oV҈�k.��ۀ-�Wƺ�A���]woj�7;�u����cv�'ZD�\l�p�����3�8����v��%���snl��r�aݸK��x�y�dy��k��Zݺ�n�Ru��3��a���	^������IS�nڞ�gmX�'z��y��ۨ�/n��۵�N��.���v朱r�8�.��k����n��2����W�Í��&��5�n��H޶�N������zx�.g��lǎ�竔�<��WN����qh�f�Zw��ۭ3Υ���h@�؜#���E[�dc�C��ʛs��Aw�>/m���q�T:�Wm�q��V��j�6w�u.�wH��˄��s�[����rqԼ`x�n8��;�i|�j̜�+�;���T�i�2�*ݹ��<F��<���Ÿ+6�l����c�;ۧ�Ɏw�E�96n���ôn8��rGk����Ǳ리`C=\�/E�y�=wEm�a�)��l<�
����0��z���W��-��j{A۳KW�YM�v�[rIY-�����l�.盵 �;��K����Ί\6�6�ftP���x4�V;:z�r�k�$����ֱi�1ڀ�X�vu4]Pi������ŝ�4�;�����1ǳi�fr/��\�ֱ;s�s��V4v\����ԉ�7��{In6[H����o� �gqf��]���.�.E��\;�Sr���lt۰'9v���3Zmy���ۭ���cpA�v�G`s�M���p�]���;X���[yLu�sp�X�lm��^=geC���z�[\��rA�<����c��kx��.�]m��.R�8�S�[p�����LX�y�<M=�3����뱳��n�e�a��6���_�}�VXs�8+aH�������{n��R���WZ}3�<.u1��m�C�?0S(�ϼ�.(V�Uu�gpr������Yˀ�,���6&��=�&�.FG�汅5z�����܌�v���0 8�T�T��2���>}{|{��$�%��Ц�N��!=k*�=щ�l��߼����ή���ױ�o7�
r�2ة�����F֛��|�]7j﮸��{;�ϩ���RtLd��߽�0K�p�\"H�Qd�I���p���)�K�l�W�<���.�����9��\im�VH���"�(��&/R&�jBi��T�Ƒ���,u<|ڌ4K�c��/�Kh��j��1L|�f���$���q�-�S�K9ۍ%�'E��8F9B�}�+_�
�	H���ȵ��v�S1�N�4�2+�o3����2"�楪�@��q��9{c�z�1�f��{��8v��`��V�Փ���׶WS��~������$�&�	<��z�W�i$�<:*��m��EW���μ�^��O5}Lp���8�a��_5���[�����!PА|tM��{=��D���t��t�q7f�4���܀���G�[���]</���u^��D�{���pO�S}�)�7?ݡ^�'�ohհob�F�J���6g�%�"�����ٺ]���ڻ'DG~WG�]-�kx�$��[�ٹ�AH�MgG���*�U~(�#�y	�9LJ��%!�T��*�k�s�%o��^K�:Y ^n�b����<� GZd{}z��{����]8��[��"�P⊪�KR������q�g�����KK��͟[�#���La
ł��1�}��ғ��T,0Y�n��:�w��s �W��e�����U���U�j���?���tf/���z*�����!>z�(��:R檙UO!N�4�T��p��o�q��߸�U��}��=�|�ښ�v׹ɉ�+�w/�f:)�L�G_���qZO���u�S�bX�ߑ����:%}�y�� �j�����<� �3/�\ʩuHuT���֑��ߞmW��f��x�"�5���_�y��)ɻS�?A���F	2���^��$q�F�­�}��t�Bۼ��}��F�m�V �W{t�?*��+�h>�oJJ�z��F��g��\�:��+'�0�Y�jZ�O;Bv�G&%��#$���Tj�oW�Mq���P���~�}�+���Y09��഑׾�y�ญ�"�5dN���K���j:ϸn~�n�_��Kjn��>b�b�p�@&.��������kq�-�l���r���\���M��TD����X��c]���.ǭ`�ٲ�}��S��	K�ep�TA���b��!j��g�X�!�q�Bß>�¾��Ĵ�
Nc�1+���j�ګzعms����֪n�v}�/&�'̯}�C�)0�*���T���Έ��i�{��\#�G{1d)|��%���9�
�x}�X���s�Q��֌;�r�:����òf���f�>�����AԬr5�m�i��X���sk,4�K>T5����y��(7B�;����o<�Zp�$��=�,#�v�P����S	�8�*�<Z�i�� ��p
#Ւ���b��~b��L�'2:�^��|�!� /�~�B�ǜ?
�f�8��֑��"O�"��� W�x��_qd.�(_SεmɆ_Җ:�:b]:%Ύŏ�5^�;�ɴ:�~��rW�z�Q�� c稨?�h��V4QI=��#f�'TRi��&h�Y���Y
��J��rz���Uy��	��*��U;�����g�v��P��Uh��9TV!u��|�x�*:E
��/[Rw�M/Z[��ů���ǅ��W��%�fl�e����y����BOs��)*�ʃ�l��<u��۫8��ۭC����
u�\]pZ����L�"��a_��-X��7�)X�.��{�\/��`���2V+k�ُ}~���N@�Y���m��8h�{zZU���{n�Hb��]��K��Z/�����{����i�';>4Kp���.���3*�T\-"���m�J��%�w��p�Z���?�E�;EB�8�x���(^��.D'-�Ir��~��Z ���H����i�>��Y��h�y�.��/�|+�*�XeOi`�,�l�o���7RPɚ���x�����	ZSf��g&�iU>C�����{7����	n5e]p�L�P�/����ǅ�7�v�{��_�{Ϥ+:%�i5)�� ��V/���V���,RQ�g�s���+�JU:EC�eUN�����B_R�1��I`�����\-#�
s�0�]婏�w�� ���Ǻ��ho�4�K���ZTޓƕ"H����K�~��ƣ��5�*0��5�.w�5�6h��S�n�G�՝���Gq#G�-��_(o �mӰdRo�`���Y�E�؎EA�����Xp�]�X�q>�ҢwՑ����e��R�_��������y��c�){'�[�»���j�.�U�����	��ò|����g�pٙ���o���7�Պ���!P	r\/}^�-r�D�v���|}��K�s��~��v��]s��4ډ��0��۳�@�s�w[��n�N��7c����ڸ�TԔ��JS�UGW�8��v+�W�)`�M�o�K��
�^��h���l���p�Bf¢Q������}��K�!aBR+��0W.z�/��r�n���)!w�h�G����rU:�����j�c�1X�,�{3�w�k�]�}d��!���<j�*v��f~��s�K>��0Ջ�U�J�q���Z�[�
���}ׂ���zgz�`�!�|}3�J��*y��>x���oS���Q��I��ǷHĺ:v��0���狅�
��|-�LxXB�k|�xk��{��	��d->��{�O�/��ܘ�m>�wD+��{9��v�E}k�O�1"�x������;_���'�N��:�|>�ưW4A�f���V@�Ob��2�Y�����Vgs�?B�t�8�7����k� �E��'>�ugb��4���Jo���RxIX����#����	�{��i��\)��^�*8t�S>R���3N�sSS.��h��!H�����{��5�_-4B�H�E[ʖ/w��FGs{��z�.��UE
ȳ⭤�7[�狅޷�����bO�n�3�j|�q�L<%dH����;��)�Wc+�4z{I���J9�n�d��{cUF�	�ȧ�7��0�7WY�ei����Τ÷y\�sj��F��B�1%[�Y�=����q�&`L<d��xJ9�����!��7cg�n4����i�[�n�=��Ӥ݌�6ꇶ���{GN�����6����1Ĵ��۾�ܼ� ��݌K6��cF���<��r�������`�j�4��%W7�; Ύ��C!ےe��+$�[�;\����n���,:��hm��፻[��n���[����)�l���d_>���x-�[w]����m�˹�m��GUU�չ��ܡ\�]u(E���Ȧ��ӡ��N�U/B�	��C��b_�������ҁb�}��
A�*t_z/�c*F��{ ��E�j��0	u�v�纳�Tw������+,��g��g>⿎���/kK��M?�B�����f���%����	��q�Y��R�X���ww���W�:����S�� }㻲��pJ���k�3�8RGyr������i]�꿅��,J�2�j$�p}�]�Mq�)#HI���zx��
�;)Q$-Yr���u-�5UT��32�Ǉ1��ZG)��g;�p��ℼv�c��)��~�x�`�}��$)b�]���>�:Ǉ������z�VF�QϚb�i:v%���iq��}p��eB�I9�I��|��Ӫ��d�T�<��L�b��muq���A֔��W=�Yh��X��N-�g�{�^v�F�=����ӇVh^_���P�m��[L[T��M�����S�y����S
N
�jm���v�H�t�J���Nj�xK�w6V��|8P�l�}.��V�0]��2��<+{T�����Og(^�z��V��������4��o��N���S-1z�YB���+L��;l\�%��m#|��4���G
냑��Ƭ�M�B�������{Zq>ۮh
�S����C6t-L�T�&pK���Q�L�h��n��w�EX�Y�+!I�8ׯ=��*#�wr�u���7՛ř���8�?X-���t�nf�Ɠ�}��N���K��D_2�a.�O�k2[T�b*+-y���\���v{ژր�����w����'�O~��`��Y^��f��ˁ��:kPS:��ߕh۵���6��TH9w��y:�g{�s����D4�{^���L�~�I"����~Jq^	����K7�"DUT��*:�@	��Ә�M�랉Y#�e)�����/�9�©��Q���@��i����h�ξx�)	����,�+}>���NU'4���h�Eˤ�7���2���n��Ϛ|i�Z���J�JTX�)��K�)U`&ץ� E���Av����^4�����K-�*,�~�_#�o�} nnt��5GK"M����g�
�T�,�r�<���*���V���2x��ޣ�2��W{���K7yW�D�$03딨�,�a?V��\�
@��t֬�>��W���i�e}Q���ب�8��-s�g'��EC֮X+�4���氌~�>)@�TE42���@�*�VE6�SJ�=m�}>�/�L��b���l�=�K�p��w�=�_����?5�z�PL��Rc�R�=�f+X���A=�6��䲛���;���z�:�Jq¡p�ڲ�����WwVa�N�-�����T���&���)�d�7���;P��Ԣۦr�u�G��Ҕ�u4v,XA樅&�ŉ}�����x���*J��@)����])}^�,�.^�1H $'/��믽7%ʮ�i�2��Y޶-���D{�Η�u_M����$�
��PL�A�G��d*I���U;s�΀bd�H����z�z�M<���7ɹ����4�D��BT#�'����Ɨ��V �3��C�g[���U�u���1!�Ĉ��A^����>���!�{��۹�����=�"F�p����=UQ4M��N�^�G[�8b�9��E�93��睯jp_%t��h�ݯ�E
�q�6�{�`��¢=۟��$��w���2���ֿ5��gtkQN9CWo���2�Mq�8�M^̌K�b =�3'>��H1D�s���Ěi"��j�xd�t�ˮ�ۋ妰W&����\����N��gu|1O��U����/?/
�5����X��tHO���2''�c��#%6�MhG:~?5�ö�?#6j�z��P�I���=:2�_��f��T��g9sq����q�ج@�Z����is��f�PHu�%�4���{��ٴ.;��ݜ^o�c��$E8�� �G�=�I�NZ�1N��PV��p�����*�*�?;O�YX>6|����{s�Zx�����t*L!gAd��V�|/NS$�c���V�Da�i_��괃�x_S�B�u��?����|8�\.�t��q�zl��w���zYeA~!A�6�$�g��3QM˶����;l����Wy<˝�r�!%�6iV��]*��4�j��~�����
ΔE�~}u��H"�E���>l �x!_���>c�z~�Ղ�p�
���g��:�x����s_���������U�E�Ф�j����k�|ː"�R���>O`�
U35UR��Z�0ZxVH�Q�����ƒV�}���{�><r�����{�+����|\U���*15�&Q;9v�g�X����p��3��
���~�V��4H��ۛ�g��н��-YbS�3;"?(���U�fi����;%|w4$E4G1��1E�R2c�G�ƺp�5gߡ�o��IU1�gޙ}���ӢVh�^n�K�|:�}�x�c4EO5z~"���S��P�> &�)ib�{0
q�H���i3J���Bt:��%�|*!I���l�Ok;�ĺ|x���ZLഊ;ږFVL,|!�۪��󴨌#�Z���3��b��ܛXGHb;S�+4�������Y�����n�P�/]�F�y�ww+kf��:��Ӯ`7��L��X(��Y}�����i�I�xf�[�rA������"D�Rr%Z8<�0�Z﷾jC�UT�T������_��(JD�q�<�j�8��M6.�m�!-N�ܸ���nv���5]�_�H}ȁ��P���w��Ջ�'���>�e�pTO��sܫ��i�H���6b�c��ү4p�<����[�U
��L��G#���Qs�=Eb��/k���ݘ�&���G�d�=jN�$���-�R��K��ǲ��6�}N(
�����k�(���f�����x@i/	�LJ�%�q�O��=�k�t�u��k���ks���«t��Uc<�ݤ���*�ף��C�4�NGUZ�Aò�˒�!B�I߽���7߉��ʭ��4[�}�ϗ�q�}�ϞB�i2N��KH]֗?t�x���1P�,V%~N�«��՚g&WFBآ���U�B���:jH��s��Uj��j��(uKx*裆�`���R��"������ň"$U_m*�BΦ�+���rr��c�2d��:�?U�{?I,�©$�/����V��P$b?��Uh`V���	��װ:P���т�'霖2+ۦ�yS(���4Ru4���HG�lL}����GM"�`h�����+�-ֽ�	K��I�'.5�}6��/=5��|�reh�:�T)���V%Â�
����>��Л��5ti(ђ���{������	Y35Z��5x�z�È݁h�,��-����z)�Xa�ұi�۳���}"I6�QD�6�P����ht�݊���ix��Dz�����/}��U�;J���4���R#�K,�����I��	|�*�L��_�U}��ͤ�H�[I��]kS�Ы�4K�68]���.��������X�}�i�:�.������_Px:__�6�Qg��4�*����+�47c�V�`twK��ʉ��Ok&�n���Sӎ�t𝍦�Ov�y��[<��w��d觋kp����ok�ysr��K��&�t�{R=�ay�u�f�^Թ�=�L�=�I��8݋��r����]j��{v̇QBc���z䍯;��9�m�����Z��4�/c]��>P��6K�n�����؛66�^�"\�Jt�۳�h���n�;������kh�z��΍hu��E>s��g��T��|�ߥaߘY-���Z� �g�v�'����#�6a�����A�����LV2�S+�J�_�e1_����b�ۢ�|�_���0|�y��v{Q���keVZ�TA�L8.Әo�E!,�TЭ�o����c���{�zv�L4_r���������{�6���>����s��G��m�*_�B�>!�l.��ᢺc���7ʫ�`��ΗHS�^�Gݮt��HVB��z�Zt�4�$�U�8ሗ	�R�����_r�����>p�G@�q��M�S�{�.�\,\&��^I[�z�_Amsۚ^�_r�`Ä�P���/{�ۡs��!����Zgn��r�u%6�MwYL}"�g�x}Sl�����,/yPp��9۽��+�p��&0��E��8\,�5�Y+"M;.@�jϫ���{;p�C�L蔪i���g9�Vh���5�����YR����\���-�e�i��T�T�R�'Rۚ��.�&��G��E��^��;�v��֐/��ȳ�/��|+Ea���_�~�#z�K��Q	�-/����0�|"�dI�(J��ם~��xa�)Ef�X��/�R���V��j�~��m�Ѳ���c��Ȝ%�6oFՕ;��T�b���76P��w��]g-��Z:i:����^�N\�%1A�K!m�xP�4����`�L{4�Fqg��q���+ت��/���˻J���y}	RƑ�������pZ1-�V���2P�/��H:N��K
BK���v�-8���Ս6��KW���}V�E�/�z5l��z�{x��� �d�%3����40'� �:�z]�`h���e��>y�����Ϡ�"���EL�	���[�����w���l��X��&�3��Ր��N��3)�ALm+���q�i ��*R�)�}n�Q�k�����~F�O����W�$�u�0T*�ӣ���SPj�h���.}*I��։�Ǟ�`O	�f� GZ��֋J���L�a'��<}쮫ZEq� "�m����\��ɪ�^���U�&����1�G(�"�w�VS4~�^n�dU
f�b���Lg���Z�c�D�2�5Sq�ѡ19k�w�5�W7�w����c������}��ئ.�BJ5V>����V
g�ũƤ|p��@I	��\R���X=3�2�VB�I�}�U$���s��1{��Z�ى\k��XÍ�e"�pL�v����T74��T)rUQ���d�dQ�tX������+o�3�<(CT���Xrku����^m?�r�VG�SML�|�G��Z��}Yו�v0�B�3bc�R�Q���:ڔtI���!h��͆6@����^�>�~�o����#v��Rx���N��ۘx�8�Dwd�������A���N�eIUG�~#���C'.w\�`3�o��ub�,�0�e4Й5\�M�>�z�i֗K"DHg��v)�g:b�_����׉ϧ�<P�Ā��I"�_s��z�!�z�/���Y͟	�\��{ddV�D�k�k[�d��ǅ�,	7��r�4\3�@��z��!l����v���o���k��>��N\>���/�*�=l@�Zwԯ�p.��t�]��V�.#�1s�{��B���{���H}ye��?���~�ҡ�KYN!�` ����l�.8<�����:��B�#���M%L��)�Z�LG��c���w�X}T�k�ߞ�4�R�@��Fxa�ɵ�
�3a�k��.c}�Ԥ���L;�v�0��O]�/r��^Z�L�f�Ͱ�L[�3]�%K�JS�w��T.�he	��D���h��Z�-�k�Ce˹L�7q���$�7�Y/6��ks��*�	߈Y�|X�ܭ�������^�oy��_^u��͝�*v�Z$z�r"�c�H2ɉh�/8%�70�o���̇t�n��7�˷�s�$��n�$��hCiS���9�÷���{�wU�޷eH:lo���vC0�їo��I��<��Z ��P�a�2@�|U<�kVG�^���v���f���m�D�U.�zD�OGe,�J���d��U�v*�v�U	�9�pL��u�0	���lN����:I4n.�p���W�+G�_7�0P�7�����V\�\����SvgAy*�vbo�l���ʾ�ٮ�e��J=��VR-*��Zh<No-�*�U��w[�9w��a��u��}���\j=��+�����v�Qe��Y�6��ġ�gk;�����ѷ��JV����&b/"���\CU�p���Ɗ�P��Y��U|�J�F�I���[3ge�}����i�sj
�Ƴ�ގ�iw�(v�`����E��Ŵ㿕�h��A��腉<����ȓD�ɔ�C�	M�p�\�ղ�X)�+���iv;vw[��[�!�+���X+	y� �-vb��[y����������n,�G��v��z��ٝXt俜��7qG�������u�,�:gX�VQ�!+U�Ǥ�W�Wi�mq��Y�-,ku���;S�q���}W��W.���%T����
�F .��i��S��s�4s�N�K���RS�:� �#EE!����|U8��/�Y������G<9�Ja��A.d /}�+x�t�Abp}��#`�cN�ڭ��`��	�7��"0e�||�
;ʯ��R����������L�%c�N��?x�6�����+�%$%��ib�7���,I�p�`ϱ�i�g��$u�$�w)���	X���\��_sI�~��^u��/��g��8��R��xT���J�+��k���$SbR$�K�*���i`k�GM�ˁS�����Y^���J��֩�M!��xm+uĹ3�;P�&��{Bo]���	k��mWm�T�ED̄ԃ�
��	��]_��&K�X�A#��4�go�<ﶳ�	�8�lB�W�A'����:�,=_LP�{�7I�xN=�������|�j���.�<D�*q޾.ʞ +糪���^ԫ�ʅ�;�Vӆ����0n�-�UUĴ�}��+���<}׽�e.~�q�6��������}�t_ �ʪU.(]�����_�p��� *#�j��)��ƅ��q^�ao�3�v� 4o}�����
B���U��ll+�}S�O�uϱ���r�[T)FN�}u@��53RڗSFF�>�(-�ɹI�BO�޽Yda�=IȬ|lA_uW-�,z�-��ｫ ��BAC'=Ω��ܟoݭ��V���d����ŀV�2&�
!5-�@�4t�Y�n�F����L,E�b���N�]1L��P�\D7ɇM�4�\j�^��S��{k��u�朰~Wk�k��+�b�'i� ƾ8W�s�� D�*(M���u�)�ՙ�͑�ׯ�`�E!�����!���Ǿ���=o򱗉R���~.�%EJ�<{o^�E�0�}��wJ����f�:&^z�Am�nK�&oۄ׫�&iO@�`��w�@�P�t��h�i��{�7 kL�i� }�O.���&�;h1�UԺ��H��#��d�@�;-"1�y����Zt_os.�	S�Y(�Ka�}������c=�ݓ;�!>���Fu�E����xxTL��+�Fs���z��5Eus���|��랴�S�s�Y�)�$�<ch(�LF��3��WG��k�G_�Ki�-��@�l����8E�v]�-�N6yuЎ1�����'�뗷*����L ;�Z�m�K�X�-����E�/�,���N�.��>��V���@������i�
�}�X�������W4���[�G���b�٦��o{9����L 3��ƙm����v�l�3�ξ�JW"�H+-{[i�>5�� �E:�D3��$]Vx� @�b��W�_u��B�^������~�=�k��5LJ�E!��c j����	� D�B��)+�L!T������^pUE�q���F@JNՏ�N�Y%J&���- �;Ɗl@�.zJ@���m:���x�q�nd���_C[0��M{�f9�r{�τlL�P�=�;>�V�W�st��r$����9[�,F�|IG����L��{��*�&>J���"(`��E6X�sB���P�HZ�U�o�~�9�o�]4>��ɯ�wSo��ߟ� @��%>sެ�`#DqŔ|ړ1�DP��9��{�"D�o��7T��p4	���,8��q�:\�}) 0|C��g߰�ܿf��+�f������* �ܒ�
F�2ܔ1?���z���K:Kf�����&�Nq�8P��M��}��͉� m5 -�(�s_g�zq���7�Vq^#�j`�SM��LAD˂���k�`.O%M�T��j�>��<qӠ���LSR~&�?O�+;�g�?�O+�#^�d�Kc]�.�)`͒��)v�_�:t��a��nԼsR	�%��vG:�­YlVm�y/���c��������T1۷!vz�k^����u3����{;C�N�tܚ����������g��4�g��ųWn_ϻv3���|i�|�,nלk���u�G0�c�.km�C���ǟQ8�.k����+�i���n�����ʴ��079�^(��:��x.����.�Fz��n,	b%y�ҙ�{+�m;K�+�g�)�������^0>36�3fL��wn�}v0=��!��q�\��L��Av�n6K�j�:��^mj�{\h�S��� ��/�d�h���O���X�#�1�Hcd��j�I"�W=śi��|4���gL��4���x�����}�f_&"�w6�n�"��җ2&Qa ��vk�5����b�y�:t
CEw��|f6,̥H��H6����}k�_�Z��g���i�nu��0%���V��4f}��A��2o[��|��s�B�pS�1�5��!s�H;����4Tv]�n>�4��׫7LӾk�|�9���y��>\��:��GC&�&�7����9����䥪�!�ѡH��m�S V&4}��q�Fv�b� ��@��S�S�՚���n�4-;d����«�H$����}U=���]�Am0��M�K��{�W����9���7�#�k�ۯ�3_��֑��j�)BF�WfT V� �MC����ַ���]6󨟻�س�|tS��@�[l{)���&g��t�	g;-���r.c� ��AY���H��"h�:��C��)ײ�Avevo-�����dj�H��"�N�h;YTaT�Ó>�RLU6:�S�V��L��'N�o�j����w*�7��<-�R(C���� 
�~�ӷm ��l����>�k ε��L9������r�._��y�/r���Z��Qc��bﳋ0=�T��3�
�(�A�A3���X{�L�~/��5'ߏќ��
!��S(�;�X�Q��]�m�X�k�|����/ki(�r�IT��S���8���pKM9�^�������Z-��Ӏt_?o��.�9XF ���8`e�{���{��Nn��kp�dpSw)y�:` ������q\0&�)�UI��`|'���S�%ρKl��uT�:͋��*k&�prK�`��V$����������j"q�m�G��RY��/�#�O%7�"oM�,U��V;�Ӹv�{�L��]Q.�����9Z���fR�5�^�ߜv��w.U���j���ne2���!�r��3Ŭmks�
cT"�]�M�v�]5>��W��`�}���&�?�����}��V�Ѡ <�$�U'-�����x`��Ӣ�@��lH�R�J=<���>��T0_�J��{m/��}�@�s�M3��#��iL��}���/���=�k��1)��@�!��[�3���c���}ɑ*Vح�bMǷv�(�L�)6S��!iF��(�U+�޵���?/ -�R���_|f�9Lb�Y	Ķe9~�1^X� �\�\ʳ⎊ĉvK�B�{��K�)�q�6Ϲ^N~|�g���!��;{��th�
�&+r~r�Jwد��UUʚ��E9�Rӄi%E%�V� T���O�U� փl���l.
�|����}��>��7s����Dj�!B�@#�@Yв��o��`�~vH @��"�����l@^Η�i	�����J1��������Qx
�W�-�@C��+�b�{c�Ms<�/��f�]��Y��۫���M��#��n0�n��u��iG �Y/�'h�o>��z�b֩yЋp����L$����q���v�H�ֺF�G��D�_��,K�_w׹E;U+��=�g��D�u��Q��k��ьh 7Rh�v�[�XB�y?!�F̵4Rr33U�':�֘��bd9��U8O�{U赳�'�+���9>���Ux~Y���Db��ng�`���K��0l]q'ޭ�k��o�>ii�+<i��)(T�]��wܪA���zr�;��!
�ּ��zk���ÊI�9h�!�ՙ�~jq�]�#BS|��l��=��eRl�h�%�����VJ�yw�8���0��[�9�0`����x�Y�u똰��V�*d�;p��"���E�6�k��Я2atl�����͝ Y��p�4\:Z�r+���S<�!/[R)�����ש�81 X�	���J�� A�m�🢓U#��R&�İ�xL�&� ����̻ezu���.	x���# 8��
l���)*nZ�c_mx�+�(�qd9�R���MNe ��ٸgƋ�ɮ��b��tE�����{��Ϲ����5�EBdnjV���_X�[�"�&H��ɪX�A�m�F
�����d_{�ǖEg��OM�Y��bw��x�=�fg@�<y�V>(� �}4��җg���!��!��=mPfR��BD��g��u��)%KH<IC//=54�6EԠuM69����{-±y��M��qM�n��vtu��^ݚ�۶��1L�K��yW1H�?UN�4��*�~��83�y�f���*�.O�����0�[֨RtVaH�zy�,��=s�7˧7�drHRp_|1����|$����ᎽS�t�@M<(�0�3�� �&G���jP�t�N�53E�0�u�>����ia��A�,�?�T�}�Gb��ި�a��x
>֕oo�,���
����;lF���zU��n�WO�����4qتDׅ7U��en�� ߞ�{�/�"�U|�m}?LtV+@/N���*���ӑ�SUF-Zdz�*<%(Vo���oz�-p�d�h@�l�_������C�h��;>�߽�Ԟ<
�:i����20�ʞ�и�zKlVE��=��\1_���dj%J���LI����5uS�]���eRj��3KcE��]�P"�X����k�'�!��3qep�(,�pц� )CU%�����{�aB�e8�[�.4}���b���Z�p�!*9�E}�i�-�?¥.�'�x�8.����«AUx�n��n��f�݉�S1�ʺbU�o�vP���]Fbc���+{u�>�稱y����<q�d����E��'N����g�"^ANT̒�˚��a|��Z��/k�Y�k���2\�8f	ph�3��gm��Ո�����{�ǟk��$G�d¢%��ǅ4�K���,Zp\!M?��	?�%�����aÀ )�r��&B�dro��V��{Y��3-T7TK�J!�
�qu�X@p�f��{:��s�oo
i��!���6�A-(�揼h�5���v.7�����F}Ͻ�Y�����$B�f�MAt,�й�����]h\�
�m&xXh(U>B��YPV'7�ߙ���v�w���8ܡYd)�BO���812/>څ�s����8_yw_!��6�&�D���p��4)��bg����B�㿖�e8h)���{l̼G�&ٓ��L,T^\�PcO��G���ֈ>����\(�i"�h�Y��x@%L��䷹<<+���T��,���x]~LV����Z\9��p�P����+#3�sUR���UJ���5�ͬ#�Y��C��:��z�I8 T&P�JQD/���p����=�$o��¨k��m�Bޮ��[� ^�wL�P���X��zH��e�b��zԀ���U��:G�\���dqq��9��q�>�.�T�M5[|OZ�-��r���}Rk�Ô+Ǉ� ���d-�^�U�	BD���jŽ���9����=��%%�V�ڮH~�s�0��iTg2;��F�V���������Y�>�!����xw�[�}��ƫeH�ۜ�m� {����;ZT�E*h�\#~r>���9G>kD�{�x��G[Z�T�OL�^���S�������O�Y���߾W��RX�i ��a��eX%�D��p{Z����J��<f"�d�0�{&$TP���2��k3�{��}��e׼/y��u��mn6鼗`���oiT�F��F7.��v���w��(�}y�Ng'l�ɽ>&��Ų��&\�Pu�f�j�d�G�7C�O�-�P�2J&���n{j.�ٹ\Wh�\�s��zYs�;�����<��;���>��=����ݾ���-�=L�6�v��;>��a��C�ɹ{{ෙs�9�\�-�,���%�A��U���*���Rk��[��q��V�xە�J=ۨ:Wm�-���9�t��n9&���I^�v���d�7k'�v쓍��	�cm!��AB��v�d��:�8ݝ����*��>�}�[-��.M��sUJe�UQ�+�|�"�N[�ӂ�Xᣧ~�>X������
�{:D�'O��3�W�Gÿ�$"Ż���L!�s��| ��w��+��X� n��N���Ӟ�uZ����r���k��T����G���ObE-K�[H�k��"��B	!��&�w�;��+�!X������W�HS-i�ޖ��h�D�¢$罪��/|�r�q�ae�������>B��{�*er��T�����=^�?����n-�>}��J��R�au�k	*>Wr�"�¯}�2q��M$,��XF)��>�^�Y����,��T�m�ޓҟ����8Q8x��s���U��P���-�f�m��>t�h�w0��s��,�$�����n��JY49����XĪ��������E�+_@}泮�r�ϕƋ��(�h����L^#���p��{��D'O��Y�|����BB,��Y���3����Sl}�P�ݩ�y)��B�p���Rt3�$1f角T�$$*R�%gg[V.�fWd o��ϧ�V���1d)��`6�����<���;��B�5�W�W��IpR+{U�	��\+vR����Z4�^�x�yq��W����fk��0x�>/�������=(pp��������sًbۊ�������v��i�.�t�m��3E]S*[5K�]#�I
O�'�F\<>�����ތ���TG	D���I�/�8�=w��o6~�*Z�| �۲	����W�߷�st�Q�J^����A��B� Z��}��lm&m'P[Hn�����{�K���Ԙ�FAIm�]3�|�ׇԜ��E���ܪ�s�X+EC��vvF�5��y�k��L�-.�ww��&L�W(����xj5��j�eթOtl���U(²Rx�=m{"EZ����C��?�S��>�B�i����'�c����mY
� 1_��i4^�!��1IID� �}�|0�p�,������勠p��S!W}��{���]Iʪ�6
�,�P��@w���ӂ���$/L�B����̩�_�_����p4W�;�5e=?W��{[��E��TBf�E�l��|\-�
$޵&궖
J=����ISU%2dTURϟ���Bb�O�yB�\�����n[��7�}�y_�|6�I�}�b�Z���=�޻X*�|���mY
��'��<^+�=p�Ϛ~k�D�]w����Z�N�{d,�}���K��� B�O�'33"��"���sJ��ɛ0���9T���s�W9^��\��PU�*��b�1O������wײ������<^�>»�� KO�{��V���]�Xo�W����~������,�����~��o$��_s����5�7^3�S�-��x�v�7����i�xs�0ܘ�mj3�ŝ�凎n보��`��Q D���.�s��8�Qv�;��Yy�����G���+(W��?���r�i��5�\+3k�_->�q���|���EG��G0��VCwڲ���{���J��jhuE����PX����k��h�^��Z�Uƾ�g�:�ל�$�Oo��=�J-_%P}�}Ő���(跫Ҵ���=S�Mخ�h(ׅA�
���Ѐ�
���2����GW�^����{�ZxGZ����U4�7-R�.id-4���F���)�*w����j�!s)��/�_��p�2֝�xj��¯�x�I�̰)h��[�;IA8��u�]-MrN=6Lѧ��{%��,f������*y�(-�϶��k�L̛�>�V9"���k
rB���RXC9/��y��Z�J�訄��������7��L7%0��K�Y�\D��=�w��WE�3�Ď����`�%�����LK
��a�o��I�B�ysÂ��z��U���B~�DTb�l�z�b�}����V�ܞ�.>�V	P������>������4�2�jn��ƼE��z��+����vx*!X�Ē���h�u�NC9�<\#��|��ta	��O�.{�X���)'딭�,^#2~�md̯)"�L�t�J�ޕ�o�O�z�?rN*PpD���z-�:�']p6U����_e��k���k�3�WVu���R�UMJO�)��*���x�a[럝{��#㢿Z�	�]ُ���|o���Y.��Q �	�ST,��~1#��Et����a
����n8.OM-5�sPd>X�s�e#�T(����Lbfq�
����R,��{ݯ�����K����W��$�p�F�[�+����AY�CU�C������KK�&tTGu�6������a=�}����5�G�Ϛ�*!��[�U*�4��9�����T%��%$w�<�}ǉh�G�N;��$^
m�o���q	p�'��yT��ຂ�Mmm+K�HWO�T+>+�^1��5bdi�"�%t�ǂ��Ĭ������M:�d��=��.K��1o�~����X�^�f{�|_L#��#��\2�f��__�_�5?0V%e�x��,�����9��	T�>����f�%�19U�˻ysi������۾7�U�u�Z�1�#a	����U�u��p����)n��o=��~r�9T�R��Q����Jt�R��TbXp�y���z�E
���;��p���n��{Z����V��#��2�GI�yw
�<�Vb0�����=!Q��*�]����qb������'±i��y��Mky��MK�t0�k��nÂn�&{v��(�<x^w<�,�&P���QL��j�Q*�Q�\#E�jE�Ĭ�IX�n���IB�}���=�VϽ�1�`�/k�C�
�z�,�^�i{2�̮�#�k�{�KH���dm��V�\cq�.��T-#�3@i@'��hs�J":��2��q����8�U�o�y�}ᢄ|�M|V�����A���B�Hd�K��I�UTG��Z��`p���TB���jH���ug޾��!�	pb��V�ڙ[&7J��RL�#���EAZ>c������[��W��\)!��¼q�
ͪ��r�������F�rҕפ*9�*,���0K��i|i)��qdX���5ΞV� ��UT������H��(r������_לYE�$I�B�r����'�R2]@�`�t�U�f����9U�u/�����p9�5��4��V�{V�M!b��*F�Qs���}�)uPԩ(����+��"�E��߻˅��$�,���`�J��ѹ��;I�,֓|&E	��)���)ʖ@Eq�'�g�t�G�e4����B���T!����T!��C�*�J�?	P���C��~ҡ�T!�tJ�4�l�B�P���C�*�J�<�B�%�J�J�?�(+$�k.N� "��0
 ��d��G|.t ��;� 4�%���	R� j��H(֍�vUh���K`5!�5A;dqiA �UED -�  �  P     �     AUJ (            y  �    [�KX��[�6m�n�JQ�a�l�X���L���=�jx� � S���]�tЛ<ON��vtoh�����W���$7�� y��^����Vt(������� �    @       wX           �x ��=Mm�0����[t�Xt�͝���s�{���̻�4(WJ/W� �@����M7�� 28�zx^�m����W���僩Q/ � �2��@      ���ƅG;�U���a�j�e�:�h�nw*��f�� ��E���*N��v�4�X\YWY�cr�KZ*� \���,��5*�;�;eE �Tٸ��kJr;��Kf� ����g��j���jդ+mqg@�KE���=Ҁ,]���;�6�s���Z���4�L68��Z-�`*�P�T.         vtl�s�$� �ˊS�lM�*h·.]�(*� =�zek[��m!m�����Z�7.�kf�kss�m�*� vW4YM���[(��S��KcD�-��rNٱ��.S�`�\ ݬ��[��v4-��ݳli-8������TSp 3����s�$��[7;��ŎnS�md�\�T�*�t�p        �v���[�T��Z�r�st:ҔW�v��eC�k\����4�1�v,�ݶ�l��nضұpt��Y�qP
���R P!�ܻ��a"��r[i#��C������5nn�m�V�1��)w(8kU� 8�&˙�l(���D[m���$��wm�ա�@E7
    
 (Q@7)�9۴j��s��CM�뭶��n��7 �uhӉ�	I���0U���m���`� ��˛�GY&�EP(T�tɹ��ִ�lܹ\V����(.�,[70�j�\�� P���N�-h� �v�Z�;e��D]��t5R���� �~�R��  �JT�� ���iCM�� 4 5OƤ
T�� "{J���� 	5&�J��` #��67u�>"� �T��(�F�w	Nc���)�[�83�O��VVa/I�H�c��:�?�	$	&�O��I I0� �@�p��� I I$ �2@  ����m�,eG�h0�ԕ�g��B�U�J�
09��ҽ��R�/a�7t3��p������eRm=��e�u�{6��m���A痭0rX^��+=�U�r��7@��e!ٖ�ZΛ�;�ZP�e�y[���ucx�T��yb�ۆ�0��3"7b��E#)�.��څ���{�P��1fI�nj�n��9-ǂ�qVI.\�>)R�Knf������w�l��������Cc)ǎM���H]�Vė%d�����X�$�*`��a�ǵ����D�Q��A��f�7�$��V�$�T��;���VK�l�E[ը`P�d�'�P3)Օ��W�8l�=�n.��$��?Xa��CF76�v�km ��;��ʵ��n3�d�!����m钭!�]Kz�m]ͽe��(\��o�W#و��6T��h��|I��]Fv�j�n�rF2� &eف.� /$��S!*��/O\J�aucؓ�<� 5��}�>�h��Yl�ϝQ����Ȗ3�j�9���X-��3^E�0�0�ѡ2´HXѼKla���Xڶ�ֳۂ�G;�f�4������mJV�6��]pW����q;���8�̆�{�`���j�P`ǻF���K*��kk1_li���]���[��C��Pq�T��UT/ufai≂A���a֘X�QU؊�yfR�8M�	6E���EcT}f�T ��M$E &",�yEB�(i�
N��|/��l""�(� tkx�'%Ы9{���i�c��87DoxW�]�Úۗ�o�&KטIע�7P�y1�7"��ѷ.e�h�]���f�ϥ����7ZS�[Y>���JK`�ӛ�f���6w
��x��e����B��Wmm�ƛtLZm�{��b��O-L�D(���[o@b���"b��Ʋ�J�
��V0)M��ܤ��m�6�GY�p��t@b1^"�Ν�M{t���3+jo�Uj��Q�n<b�fh3a���<���Vbn��)kA��V`a,��h��#p=*2������
͕v���Yl3�\+&K�Vwp^QIfG
H�52�3�,	���2�\,�^�|�faK,"hR�0R��(��Ē�*ʁ՚k@��CH���qnV��Qb쬭�Vl�\M� У�u���e�&�d�[��ʖ���%*�ͅ�xW��n����j��D3� �͛P:b��Y����kZ�]eɏn�ڶ����5��7�TY��1�V�љ��X��ժ�qt��Lͦ����M"�ᵧov���H�[��L *\Ȯҭ;�cݻ�e���<�"º� S�1�6�Y��U�O��v?�V��D<�DP޲�U��7��	�Ԩ�� V�5��ӆ�z-��7�c�@��=aߴ�.�F��#\�E'+�oS��u�l\9�Y+m:.#�br��*�Ne�$R�����xnd�Rud6L��O5,RG2��7��d*�RBiQ�n�aTr���[S$b˦�ϊ��O2R�o��
�H�%�*ry4S�ueGb*�#�W�&�lgr�v�:?jEn���%�ѩ���^M���
&n�P���r�k,y����F9UpK��x�N����[om���EZ��[�M`�K!\Se�M1�p^ۗplST˙�V�d���#Ou|ݍ�cqd\@�z�%�l�{F�R�����H;���HS��<I���p[��.�^���[X�ΰ��*�X�8��Ji^
�L�S~^E�k<�^ŕ,�ԜT`�"��(�oYȫ5=��m��2�PH[�U ��x��@���C3�O 
QzF�ӷB�L�̕Xُ0�������bZ�"��j-P<Vm��zЇ��X�J���?&j�K�B�:��:����_�Oa�T���*�2��W�|7G�Z��4�sP�:�QC��`d���T�H�^�T��򞺧�mH��5&�@��˽_��Q�ݽ��gX��ZŲڔh�U٘V��F��_TN����lQ�s��˅��[�K���e���ׂټ���5��~z�J�#Pˬsv�c"x��l�}Wr�9m27OLn�j�R�p�}XoF�LVlcNK��r���0k�{֛��V5䰕��L%5��\ghۺ+�;��̅��+Ɯ^��~6b��r{�6����jz^,�Ĭ1 jkL��t���n��͢�{VfT���KV�,�jT�̧��U�̑�D�Vt���j��KgƋ�X��J��E*����X,����<fŰ���WY�H����H�k̰&TlSY��b�Vh��7�^j�dP �ȅ�aW�2�֡��S��ե�V#��Ņ
���k��(�e�Q�/-��Q֭��r`;)=�v�ݡ�"��� <����}��񼍡�sQ��kӒ+��I'8eQ9��l�7��X94�U�)�)���{��ݸ���E4��bL�XbY675[6��5u�x͋.�W�2��I���z��,�<
�o�H�V8�d�3D�&�����Ŷ�
��i�i��{���$`�a�ZW6�D���6s2��-f��$.��Ki��3,��%`�H�˺GS4M]�sE�
�In�șN��j�!�����N�+ez�5s�:�|��	+r��K�YEު
�ҽ;�k�2/(-���"h�v�4����x�������ױ7�k�*�OTf��q�1o=�.��i�C�5(��Mp��Z����C�@[��|�
~�	ta$R�a�j�6�]ْ�Ҽ���N��m��V���)I@�yG+�A �T��q��	�4,e: ��9six�j�upФlMp@3o����P'D�ỚlK�fLU�7��8/)(m��~R�_��3�(\v�O�3�:T��n^Mt�6�l��31@F�XPw�Za=ɷ�5*�am�2S!�
!�lPm�@�������7"�o^`�-S��l[g���!��hT;s*f�i3����%P�W6(�,К1n`�gj�*���f	��#wHMT�7�OXr0���\y0��>2��k_�&�j��x6æn��R��hG7T��K�8ePk%��1����+5}�61�!t+dǨ��1�a&َ��m�{�N��^
�+&�U���7v������\�X��3(݊U�3d�u�C3ed���[�m�q���H��bgQO&����zu��30��㨢ͻ�Tgm٘�rE�����hz�4 U륄�
�~cۍ)kR���^
����Y���X��_�l|��	�MX���n�'��
a�;�p�-'c'P�m�?���z�[�øi#[�j*�9t����9�c0�/���Ĉ^s6�2���m,�M��)���	�a����9)��ٺ�7�gw&UӁ�������5�R�OVY@��Q�0 2fi[���|(Nr�kw���nU4�,��^(���3>P]:e����Y��x�E��BAU|���.�72�ʻ�L��-�D�h��@Z.��Xd����u�eMXp���.,��ɶVB�r�w̖r�E·夷�2��4p	�V��}�&�����+z�3Rf�A�?��.�����*"Tն*a�j��4�;��A����1[�@�֥nm�mV;r��E�Ln#WGEn��	�:7Y��.d�w����7�p�>�L�,$�o�ݩ�=˨�R�����f�E�C�%N�u�o>���WU�)��������en����5�G*٬�%}�^̦�/-�O�k��){tN����P�8�����BN�E��Ӹ*��]�5���)��:���/3x�μ�!�I&Q�.�/��$5��RL�K��2��HP{�>!t�Z73r��rN���]ֺz���1�F��u��ջ����jɪQp��KĪ��i��oQ�U(~���<i*�
�~_L5S�:}�#9��M(�|�I�&�3L�����2�t!]��*�ƣ����%_l=K��Ҕ���iveA�[tk~��/}�tS{�>�ȴ�/ZDk����1,_3���@�@��Ǌ����ܪ�z�ʺUk���>��.�h��ի����*��+��
ޱ�i�(�T�Մ�hRV�b7��;.�T�)���Y�F��W���[ʗV�L5!�LjsAb�呙c�./5���t [Ku\���3T��ۗ��-n),�"��TU��O�M:Ӵ��eK6dFa�i�cv���|Qf��r�9Ǧ�U�W{M�+.ӽ~�ҹ1���`�Q�����5c��q�7F~]Y��g9LN��I)k�k��@����)�"��-��q;f2�֞Sf�J��F�W��-m�9Wi4	��{��c'kJT��۬�b��7*]�8�4e���t�|����BlV�S ���gӧGT�np�ò��Pm
�yF��Jc=�z� ��P*�c(�z��Ԇ�� .��r�yY���i�R��b6V� c[	�N�2�-�	�M����^M�n�hM�+ڼP/�<��!K�t��r���՚��/VI�>��<tJ�+Raq��)]Y�/*�1���6��R���f�����1�Qyd�8� ZG��yR� ȱ5�Kt����f���+!Z�,�����b;S$�����K+�R8k�ӬJ��5���=j�M6�B�5�Ś5�X�s&.k�斩�!�����M�!�e�w�d��nc�el�LώB��n�B��&�,�H�j!tpL�l��
�����W��,��ݴ�K.���
̉�V
	D]K۸vS�Z@LW(���ehŦ��6�J8�S�fD�-�9h��+!�V��l�#F�X�(T�#S�
x�^Xm#���k��vP�viYv�ٽ%ꕰ���������]ǈϕ�_���H�IS���(���&��{����*Hl�+h���� �����2��E̺�(�M��l�d%cr����!	�r�h�2]Ԉ�sqjKN�����e�1���E��+Y�V�0x+�ƌ\xI]����9WA-f��J
�&�M�X��QQU.��@U�ѽ[��3�R��XׇP�r��b�o��Z�X<� H�R"�ɕ%X(�Z���Jm��F`͸.��V[`c�n\"�"�F�^���j�Z�y�"̡�X�ԭsMdwOk�s���kغ��>����U�䑉m5�t�LV2��˹{齛�Ä�u-�R�Tk-�k� VG��K��n�\��ŵ�)fb/���ʙF�Aj�3Bvv�r�b{vՖɇf��kUfA��")Ͳ�5n�:n�GA�P�'Y9t��O�eL0I,mj,�oM��l�(�Ê�� ���Z%ӵ>k#J軫[j��:�{��Z��W��gh����2��F�9쬸���}��b�K?o�C��{�����W.�ꉉ:609ڐ��M[߶�����-Z�\����g�:Y�N���)J�c�@���-����{ux�o����yb�VU��:oZ��Y
dXU�W�`��nЫ �V�ܘd�'th�}���mf��U�K0�]e�3��������m:��Q$�&��$Y���7&<��mk���]��C�N�ow.��5�=��[io@}&�ln���b$r�!+)�2�X��h�:P�+�g)eƔ�TvXrW�woUH�EѨ�],"Ťr���6e(�{Ef�%�����R8����f�`��[|X�8eǆ*T���-�s�r�k��xݰQ]se��ց�iW��yɮZhw$V�v=�p5����]�눛zmލ�����'n�G��F�F	Y����X��^��#�i���5��b?��"-��d1��nVXZ��h��Q"*��u�s�����֒�5�����dՂt2Ѥ�GZ�3kT�h��T�
+];��dϮ����IQs%,�&�ͻ�ۄ[�scy��k^��^��D�r޵�aQiZ���2��*0�n�v��cыmԛ��e%{�]�5�l�v[��;,�5.e�L���\ϳ�h����yC'��Tkr��u�"���_K��g�E�J��gl����K�)�����R�6�񬃤o���2MU�*���5�I�;d�(��𴱉���.�r�ɫk��S�3n�[u�e�()+�h�}f*���+u��wgg]z6���芷����ڙIEw)���^Y�pk�Q-H������$�A쇓H !"&��`S�"����[�j�+���6��
M���f��x��.�į�T-,Ö���_,yJ���n[D�X���^�F��m�-*�a`][AL� ���(���0��������+��<O<�fՠ�2U�pQ���eǭL�v�;ph�d�-:�L��h��ިZ��d�[6�;ǩf4� n*&�Yj��v�h��5t��F,ѥ��%��^D*�,b���ie�>f���+pܨ%
{L��^�d���dä�M�P�F���ۡ���D%&|( ���҅?!y<����:!|F"��rG-�[ãp��e;RvG�*
�^��{���ٲ�h�0utN�=�VȭF#
4٬5d`���Sյ��B��2n�j�mY��n�97i�f���>���3EΛ�u��k�ާC2m����2�Qk]-�Z��H�Ö��9OG^�Ǝ�ɖ_Gx��6��Z:����֍�8�xN�A��WQ���Ւ��6N������j[R��
���bbbn-Ɓ�wD�e�̈q*+V-����q�0o5��-/����I��eEF�SE�_΁*.����&;;y�V�״�}fh$]+:0�f�m_��`b� �w���h8o�7�n�9�U�8�V�u_ Z�aa.嫕V	P A�F�@�A���4GAcl�I�Z�C�Z��tYF 
�Z���UT�Z0U���^8�-��)��@PqJ�@@N��.�0jU���2�n�U^��#������V��)�C��
�p`�V�*�
����vUj����9a���������jNl�uZ�V5�R�c<��3�m���Շu���{�ݽ	�u��)֓�ۆ�'<sb��M-pu,h�r&g���8���U�c֗�l�ƈ�[9�8�x���[s�a\�4��3>�#r��"�P͹�j�nM��p�suqn�,��z���q��� ݕ���\�R.��v��;�+�k˖b�%R(�T�$��cy�aqH�����i�qBi�d��`�EK����zq�o�5�X=]U��	Ź��nƸе<�I��q^�tl��㐮�����;�n�hV���*��v1ǘ��쁧{tOA��v��p������)���YZ�"����n�lo�ڻ2xd�;$�͍�6��Ü�!�^۷5�۶�<R�۞�c��J�=gQl��h���1ֶ:��s�w]�1�9��F�{dW�ɄM��7|? �ʉOmy�Vp�W�َ���o ׹x�,�������
��bˋ'[���V�Wl=�����l������j�uq��L��'rg���r����l���~�m�f��\�x�n�/��ʼ����z;��b�b�H'F��1�={;RF6����lFN�眜R�r�N�j��˃pn�۬��36�g�A�s�1��C�Dz�A��Zi����an�k��\{&:-gz9�uq�X]�䎊n�q��r�'q�qmٮx��3���i�a�n�'H��8�cڬ��;��m�7;�U�۱�=nÌݬ�m��f��vMph�e���u1p�˂���6����pe�Q#��K�r�	�n4U�tN���<�r�E�+6y ���G��9{u�9�]�.�f9d��������A�;s���5�4r�gs�q�U�c/Z��\v�&��n�m��!:`�Q��E��*�կ9����GmN�v玷.��rE.�vj�˝��>����]=6��Y�܎�s�L�Uގ;=���ۤ�n98,����^�g�I�ۦ����M<��ƃ=�«m�2O�p\����wk��`�7:�lrBy�:)�Y��ɪl=����z�籷�%jpu��6��𗞶w;���݉���q����g����;���F��o7`G���g�
`9��ݒq���]���U��'�<��G����9�n�K���w��v##��G@���-�]���Ӵ��X+�u��a�0�Ѝ��sѳ����u���^ӗ�Hc���6��pv���M�ջn�[1�;���b�l���v����c�W�9�k%�u�ݶ1�]�3w&��|����H�=�����T���N��V��h�;iic�[����<VĽ�3�7g�]���;��pr`L��m�6�';�8^�[���㫀c7-�v���R�lUWl���`�!�|�[�]�9�< ύ�b�w/k�s��۶�[�n��=�g<�nKv�զ�6�m�v7[� Q�������rv�c�z��z���h��\m �L"����5��)�29͘�ɇ8��,<�ŝ�S�3�cZ<z紧;C��ɞ@이�ܴ�n9����v������8��,������`f�>z��tfs���<�=�n�^�Ջ�=��ݸ9��<81�x{v���Q��0�=�փmէ:p�������Fݞn��^����v��f8uFp�ۂe{�g��p�uk�g�<��.�-��s�kW'Οem�\g'T�����ˎ�ʷ].�w���Ι���jQ9-uB8H�L
*;K���ܝ�N햁xk���8�֊wm����Y�7��난�}gk>Ů�Q]�	n�}�<��L�lv\�=�ێ���\{����T݊�=j���t�5
�j�1Ɣ��ɛc����l��`�{l��ۓ�条�����j���qƠ�Ӷun��\{y�x�U����1��� ��x���'�!:-�u�Mm��>瞣v�7nՇ��[.�M���k�ض��{Gn�)��g����.&��ݖZ��(cv��%�k;+�q�3�ݴ��]��B��切k���0}�>�9\m�ԜQ�r���2�l��'����l��v.�[�ۡ�t�s� ��uٟ 0���G-������ݓc�v��p���u��/lsvD�W�00nv�p�>�n-���y�Ò{Gfz:y������&�]
�ש��y�=�\vum��B(x�M�z�U@��s����%)�=���H��.o3S�2Y�Og`���[�ܾ�BV�묆�v����vn���X�qt4W�<i��m`����O.�9�/u�׀ӹM�ۭ)k�vvG]�F�d{+�]��nt�Ŭȳ��Wv���5=rY�ݳ����|���J�aϫG<�6۳h�uz�7i���[Ō5
�nP��Zг���8��u��\D����[��}�r�\�8[ç;m�vqp�;s]L�6�����#aݖ3��q������,#�n[�c�y�����t��vт���&ݫUc�{�#Gn�nԇGO[spgk���g�N�ul�v�๷om�Hvѳ;�:G���z�r\[�7^N���i�ON6v����N��kc"&�u.�;�[uN:�{��}�Kg���Vy �#�'��8�.���;���<��ݜ3Oq�ㅎ�����ۑ��Ԓ�1����2v1�̎��WY�9 7��J�	���I�gs��Xʛ��a�J�2����+�}:ۮ_\��[��]�V�k�!A�u��t]��t��f}�[���Q�_�8:"DWx����л�0��ݮ�8��B���(۸�UD�7�;�n�`�}q�_;r�.��+ET�&6����u�f@��M1� :��u� o<���Ǯ����þ�:vF{E̼�
!
֠�
�bd��iW�gg��m8��ڻNM\s��mWOml�.:cɍ���ۏ9�	�/'q���{k�K�۶���y೸1�ۄ���w�x�B嵫��=��.����'4�kvx-��p��ܲn�6�'F���!x:�s�7[��#z�\�:�ǧ�+;;��ܥOd|�xW.���Ϛ�j߅�����0#����&+�i�C*�B���aP�kc�m�d��r�6��m���X׏JN���}l[V[��XώK9��N1E��K��)��ڻuw�[�����<�$�5�Sm���NH�Pv��mױ{;-h�˂�N<t�/B���m��нۛ)ʝ�gx��5��gٝ2p�c�)�����WR�sńN'�7\r��=��`��r�n�L]C�\��/.7V�Ҝ�gą���d��
�HӇ�\���W�X[.Kt�M�pU��Q�V�+G͢8�r��E1
Yz:� )¼S\gX���m���v�q�n��uzx��8�Gt[O��z-�:��\�ۙ�;b��^�9L��ٍ�XD�m��͒��л��� �!�SNv����!r�����ݧp�>�2e�.I׏lO�Ӵ���.<���Kg���7+���v�ڷD�<ې��Nf��<�O�S�Z獱�';�N{h�ۢ�ݹ��	x��x��O.�x5���m1iZ�l�0*z���+	k�d3�n�4���aG%^<�pp���v���3^�<�S��e��cV�v�|oSױ�� �<t6s�!�.3��{7\n��x�(�=r��l`lfvv�s�.�J�$��S��f��mvz �[��{hv6���j7��㮂�՞H�����{N��<���y.��;�2u��םgۃO;Q���g���V^i9���C�;�����X�Y��&Y�i�q"$��1i}��ݜGg&:O<���#^�,t�Aۈ3�]=�V�Ɏ���v�oײ��#���Ǎ����g����v��y���9�m.�
��j_n;[t�k��Ƹ�.�%�/S�prL87j]t�c�"us�l�s1�Ǯ�x�����wd�vul���:4�o;�]��v�L�	�Xɮ}H���[Ԥ���䍪
wYn1�����Ҫu�κz�����T��YwQFݷo9Ggv�f��)��n�X���=��v�����SIxp�+CɄ-<]C��s`��s������Gm�Q��.۵�>������[Y�D���u��[/kuUk[���M�&3m��x{v������nCWg��Od�qճu�:$7c��}˷l���t7\nn��p��-�݂h�zsQй�A99y��kq�vph0t����%t��Վs������W(���U]�;g�����L<�#v8��3�(�|F�}�ksnW�퇎���b�������X���p5v���b��vƤۘ���	�u�����椻`mɆzp��
��a6���������z��9���6r��Ŏ�z:'�5�hݘ �����g����f����hr%Wn�1<3�f���},�tmy���.r��ůX�0=���g���a7c<��3�3�-�rmã~+@� �c��}�/X�tu��øݸ�;Uv�m��vN5v�����q��n3k��tn�m]/�mv������g��ϝn{I�;������zԋ��z� t�¸�=�PC������������c�}�	�ݛ��n�Fe��n�/K��k�{nπ}�X1��v��f���j�m3{v��7+�q�՘���Ԃ����L��uu��]��d�z�]��#��G@��N3�mǶoa:%c<��a�ݻmd�G]͇Fmm���/n ��y��|��U��!�O�[$v�����[��^�9��ڷ67k*>+��:.����Dј�����"U�81����i�n�8����\�W'kB�9%��.�.���V:�����BBC�!����P	!O� �@�0��@[��)�o,�˻�̻�N9k�cu�N\']g5T�Ig��.a��ɕ������{	��;Օ�g���ہp^.�1�q�>�z�X�m��݌���˝٣���gu��i�+��g2��W)�]�JVe�rf,j��q��{m�ճrI�g�<tq'�a��Q��7b�����g�c��^�<1m烎Ѧ���1ӻv����g������,�C��N�ݮwK�%��v�\��)+�Cm�v���on�ڹ��'J��9{r�V9n�x�wVq�'Y:�E�����k`ڍ8���na�vòrl����<l`��ֻp데n�d����t�s�n��sF�R;l
V�{Zғ��H�ggwƢ��d咮On�1�M]�#;�9�ۗ�����wn�f6�8�]����z�f�lc�t:���-nڐMt�3����iջXG���<g�r&�m�ɋ�5���V�NL]��,��R�v�{f��Yq8n�q��amv�8�c�n��å0�W;z�׎x�h�ŝ;��f���-�0�-���<vW�-�����m�t"��.*�8N��nݗݲ;7m��t�i/([� ��ɹq�F���[�\��v�w�5����[���c��XG'l��zF�\u����j�O'�n��;�0Ŏۘ�9�SG�yb��6ѭ��v�cK���\J����ѐK��^�<�s�6����QI�ѹ���=s���Y�ݽ�m�5�rl���s��i�D>����&��D{��5��g:؎Z�1%��ڄ��z�벆�nc�#��Mk3��]�yc���ڛ�Ak�A]q�6����]��g�n;�q�7�@�dzi�^݌۲�V�n[�\�qTN��c�m���7cn���/'x�����e��N�'�Uu9��˳��cnr�v�y���7<��,���k-��<�6ۣ�82=F8�^�4��Q�{uK=���@Nt��;u�A얁7&��DU�J�,l�?ɀ	@���)( I E�) $BM:��]��ի.�wCɦ��H:3�&@�n�y�'����c��<e��\�fh�;GE�q���\�śy����͸��kf;��vp�A&\n�'m�ڡ�^�;W8���h���z��]�o-��:�Tyt�D��N��٭��^y̺Ǜt�ā��C���r�8��im�ڞ^Hʗ>]Ƿ3�������^^BJ��#e�%	V�T�6-"�.{�	�UL=�we^F�q�$N�e�8ڼ݈�y�*����J��}�=:�  7_����3��)�4�sbP��1���>>��f�'M�Y�b�k�~���u������G� �òd[����`>!ɷ\���g�R�w�o�lv�Ap�[`�!��aЦCe6o;�o^1���]�]vg<������N�~g���g0l�}{��-�7�^?�	��E��M1LޮpIy�7�~�K�J�����u*X�g����"��Mx��WP������מ�@�f���H%E��/�����=�i���v�y�V����#N�&2���$F�x�-�C�� ���k�*���֯Wl��s{�8����v�/w+M�ՖH�):�P��<����@Dk<�J9��!��g�d9�nV�'�Wd��5����91���Ι�pۉ��٤1�ک��9d���u���U`�)��S���V�Jψ�`���{�X;�Sۢk��i�f��Sy�3{�o�a�̧1r�/*���L��W�Y�#�s��"�`e��=�)\4:ٿ0=�n����[8��<C�Bhu+}�˫��+Zu{�}�Pa�`�6��Y:B򏈆��֓�;���u�)>������z%v�䘆���H|���8��4�j��n�<�l/��g�;�
H��c�v�z�ɩ
 +@L|�Q�D��°v��8@�x��koo�sm�޽f��{5L��La��&&!��a�Y�;�e�`�2�3�ܪ`�@��<HS�{Tf�\~z�ֵaIh�/��i�p�֪ab��
H��P@]��i�T/0����S�2�}�a�i�樛x��.i��u���y≉�@z�q�;a������ �[�gW���NZR�`��߼��*��E|kƈ� }����H��k/2����L���7�������3Ո�:�&��g���L�vNg.O�E����T���Ϯ������
����3L��8ӷL������x?9ޛ�W`�x�0��F�����\u��9.ۍ�c�=�Zw<�pv�;!��<��ĳW���9uOs{|s����u�>`=�1��[�s|�I�_&%3��1&j��Y�k������V(��¨�F��Ԭ���%���U�,:j�~���mJ��n�2�i���2c�Mw��n�����R%�dU��<+CV�/ջ���~���Í��!�<�11C׮j��u�)�������k����(V�|��v��Y������V9�'V�ﹷ~.�ۦ��f5y[��j�gP�QI����{d�}�I��j�mn��s�s=z�TJcӴ�*��u����/Ji�M���0��J�U��[����'f�ҦE�x^�H�Z�*��e&�h=��ʾ��_�oq�Yt�<�*Nw�>kt|��RV{ڽ>g�j��L5z~��X�Q�e]�l��,4��h�9���́�|��\��ܟ'��0�e��xo^̇o�LЇ>/O�K���v��`x�������:;ҥv�}��m����3�6�,�h�Jj��A�i�"@3�{;����� �Æ{��VxԲE��T|�|����~�k���*��ޡĔ�0a������P�6�į�/���05������Be��sg4�><[��Z��I"�r���Vg����)ü�:��6�ǧk`ݻu��9 ���
E��K��RC�9�r��gף�2�s㿨��M�����2��y�E���V{٠����έk}>�>|�$��&ߝ���KzÉ�n�"�OM;���Ϋa>t�2�ϓ�)�,6��Y侕��ՂӜ�;[�Yɏ��tL������>���5���(�Ϟ��c�=��'j���MV�bC�Y�a�d[iy��N�/zcA.χ�
�x0SX��?NBI&fU�Y8�_��4�������zO�q������Wٗ��0�4o1����뿽����%���ϛKv�7��:x��Gr�������s,p`���%�s��"�i�=w#�,�{W�:�}Zw��m]Ctsvm%������ S9�'��i��s�����j�a5V�*����F�<�˴��)�K(ŴoG��bǽ@�U�[P�ѯ�_u�2��a����S�r�^�w�k�M����Փ���}���T%�jÎ��c<��m.��uM�mf�fQ4�*U�����נ/yAªsT}�94�gy�o���]+��薇P�Ͻ��P,��@yyV�|�y���^�'Xu%�L��6�*�~������0W$����^��٤���K#��\�����qM�$NT2���s;I�
|��I�Zm�i��I_U'Y�^�����v���*��8�3�N��Z��;��~{o��&!L��γ/|�h־���>��(U�Ǌ�]�n�i0˼�8�y[N�;ʚ@"�W����0ȅ�ef�&+�����[~��F��ٻ�����ߨ�M3J߽�f��6���wjbe�޴�?_�Rm�>f�{�e���i���+|���~�La ϖ�B��x����Hg�z�+z�lJ`^��M0��N��z�6��,������ͺ߻W��6�t��u��CU���
C��w�;++�>ʗ��q��񫸛]�]� 5@���_S>�>�U�t�}%}����q�l
|���8�)<�{���,��!l�9찮{�40���d���t�ak]E�j������	�`�� X���X��G�I"[�R@��O����N�ߜC���ݜUN2m�w�w��/>N-<&U�W����ɟ]��ic�K��w�wu���U$����W�$�o}��6�M]$��Q�)y���9�M���T0�,�����׀<,WWG �j;ǃ��+�����M�nH�]Z�չ�s���3wyn,���5Ԛ��-'�ݶ�@�3g�%v�6��;�90���{<V�Wu�Ǯ'v��ݽn�ۧP+l���q�F�J]Ѭ�W���t��v�V���7L�u�k m�Cu���)u�vv�����q�.v㮓�)��v�Z:�裂��}�mv�y���ÈW�����]5��۶G-s�3���(�va.�H�=�x��G6����.h7:��xLW/D�O�ŀ;�v<EZ�]�t*��mz3]�nx9���]�}�Y�w�~~�O����<O�	�5Z��$4����b�s���y���߷q)	~��l��޽M.��x�f���y<��e�ʭ3�z�2񆾢a>���C�����)�!�F��,]38��Rn���%��>��x����}�N�3�e��3|��k�{4E"��uE���;�g=g��>q�ej�޽`W���X��o�@zW[e>k�)��_Қ�W���c��=y�N��7�뷾���8�N�����ь���3U�����b�6ȫ>�}}�@�S��u�����n�ϙ�m8�yS{�p���4{�woZ�i�)��_'�-�R������n�zk���Ɨ7!.��M�d�����������ji&�j�[o�o�6��kU�v�}��Y���A�5�V���Qe��ܣ��V�.�3�i4��e8�Ɍ6seՎ���.�`�^a4�'�c�֓hi�t�k��o�M�E�%';�W9��;m��R�w,��Ch���chY����3��u(����0�k��a��Y}����t�7��F��+������)�I�m3����o!ٸ�z^���L��3٩�|-�M�f^W;T(
iS亣in�F�������2�������'ڠ��q����Lzѫ;�5��M���Y}����5�9��|c4�}�����hiq����V�Aʄ� ?�7��>����!�k^�{���Zk��[�@�@�Cz�^���t���;�T�yB:;�+1;�g�P�����t��V��Vs�W�e��8͐���n�+��f�E&_�Èm���n%eCwS���;z6�8�W*�oU�kצq:���W����y���V[6����U�IUv!�`JL�m}��8��]JwU�)9�{	�۾גbV��J֛B�S���b�Ut54�>Mo�k*��:���W�Gg��{;��̬�-�A���Ff\�cC��FӿWx_G�문딤`ܤ_u���I�=���o�-����?^�3�G���,�u���?{�;�.q���7@VRϳ=���ԘͲr���bf��u�u���ﹼ�u�z�l]^�n���&��QV�,��CI/7�W��˖%�=��8z���5�k�0J4���!}��O��6�N��}V+�>"������c�|�(�S�y֬3T���g��f�Ki���M�Ja�{V��y^W��/����3����xM�wlEֈ�]�GS�91ڬj:�n�x��Q��f;ߝ���@�䘅_����Nv��AM'����̖׹f�|޵]�mg��������O޴U9��}�ʡ�T�W<3)X=���k�RZϵP�W���4Wz�V�wW��U�|�H�0�����s�z�*Z&]]mH�Ϫ�?!���8��v�Í=a���'
����]޵�L|�q�;ڧ�7�潛�ZN���D��%iW�\hk�ٺ�IU���`�^a4�M3IiY^~C�8�=�f��7UM��>L�%4����M3M��Xfn����i���n�{RӺ=�:ls2�Ub��q}+���Uk47�U� �T��7����jkw����kޘ�AH;�6�7(�&�b��*�
��{��'Z��ǌ�3�V޶��7���[L�Qf�g��qR����k0�X��t��Q���C�i�ȍ�S9�NwW�B��꯷Aǯ�L6�s^�8���w~�4q6é��>�1
|�}��%��8�'��W4�_Y�d���k6b�S�1��q���-4��Uu��B٢˫p[����'^��1�U$(��}L|r��}Z+�8y`�fz��υ�v*�9a���C���!���5����1�P[:�u�5�{%3\����_y���L��.I|�Ǿ��V�t壜7i,;�{nt\���8��գ���on�<nx���9��׽�{�{��N�O;��N:�S��V�����[�׬O�]m�4�w��=v��9u��v�����^�_s�γh]�)�RƳ��h��>ޯ���O2�gگw���N�,AJ�
����IuY=����\ִg��3���7~Ci-���u\ʜgS�a���WՎ�c�빠؅1_V>M���|a�W��d�W*��|��tKa��_�G�>jC���a 4��Ȫ&���Zv����m��:�Y�u���')0 �W�}~��|�rk�������o��y�B�M�uh,�k��ɵW�.4�=U,��ni7m���G��1�����-}��Y�U��"n{����k{���r�ݠ��sU1�~�l�P>Ͻ��<e���=�{w���7�*Ur�v�w<:)dp㉗gV�e���H|���v��ƈѹI�窥���r�YA�ر�U��g&�sMݘ�e=�eL;��lZ��[56����o$��Z�J��|�ȶM��������te2">��v��O���E~��Z?U`�����]oVɕ@�����gע�P�r�T^�۪���A�)�~k�iP�)����]La�!����e��;vl�N�v�]��c��:1�7l�uuZ�%	s-{�u����S{�{[KN3�`�|hG���Zy���ԛOĆ_���<��g�4c;�}H|�08+�V�UaM���a�1>E��OUj�yu�.�)�p����x�5U�����{.Q��|�ጽ�jn����V�>l����-�vk�I�f�s����oF8����;��ݣ"�O�w��ɗ�T�[��yS�Nޥ2SI\*?}�����LqIi�>ַ�L��6����8v�����u����R���ҾC�[�C7����1�e��A�Ϲ4֞?���Kbu[-�V@y��h�^}����T��pR�>�8?�W�O0�*�1&���������1�f�m֩�w�����ۨ{u�"k�Ym��6�cV���X�@����(_��!� �X c�:��>�]g8M�@2�Wu�W�r|��B���n��GP�u_��a�);�o�zus}�r����O���6�N���A���u��m�x���hqӭ��k���;�4�?��X��:��r��=�q���On;ၽ|>*��r�t�X��p���w�y*`Y4c�Ej�/�=��\hY�l��Sh�����-JM�I���ͻmx�v r<^ӣq�F��ٷ[�ln�L]z�;e5ocpG���Co�'a/-:�|�Z�:Y˓���X��蹹/n�^��᷹���{%���8U�mۇ��k���<��ԧ����˦9�vՆ��rf���l�!c��i�GK�9�8ꡗ�q�q�E�`��+i���ێ�͡��\�ӵ殩!��rE�Dlq/$��Rs�՜e3ճ�=]\��9���-�z�ɂff[�����-?s��!��ZՓ���:�Z�ɤ�=���P�
L�ώ �UC����+��]%�V����0P��*��g���
j��9G��Ѧ3�pq��j}y�L��2qv��B��@�{����kes��Ջ��w��,Mc^"�5�mW��q�`y)8�����r�n����_�Zi��ۛ��7xY�l��u%�if��n��P�u�������lq��5�k	�1�)���	��j��6�&>�Nt����>�>b�c�
�kWA�U0Ĭ���5}�΀�,ƛ^;�[�5�n�hAiRl�4��l����z]��7��o>tU�'2��i��7���4�r�M��s�V�<m&4����{��^�gn�8�N��&�}����{u;���C���}q/&Yt�7���I:�����ZO��`|۴ַ����=��_V�o��i��9�/S�-��Ql�^oWǉ�U<�.���=Z����J5�ֲ��S�gTV�׭H���؍��ֺ8ʁ;���3�	���7]����\v3��)`�F& ��/��u���1m�ү�ܸ�oןz�q�N��6�M&�^x����Nu�q6���m��*)��{4o;���ֺWu��a�1��L�:�|�Cl�*�u%!׽���[��ʲ��̹Y�z�%���-4�|��Y8�����f����GP̵��鳰J�r�&�n<T�Zq%�ֽ���ҳ.��y.�;e��ƺ�=+��.46��' ū�i!_c�T_�E1����y-��g�í��1��m�Y;u:�*q��3ݽ�$�f�=羕W����q�������pfEG--�R��}g�M&&)�X,�����ՠ��}��e%3���No���;�9���a��Pg9�u�y�.��N3YS�}�4�R_*�B����P�o�����M���P�U�������[���n�����w�q���Tޫ�{��d��:'ܢ[�Le�a����;m����EEj���k��9Y���6Ȧ��iw"˝��9P����N�/���u�ˤ`^�z�}��q��P���b{��u��s�5�f��Y�y<�MeJO!�޹����������;�ߓ����1j��P�>����V��}M�;}�Ʊ�{�s���\y��M�Ǡ�nu��6神ɝ�g��8�v����jF���,�JT1�>�}�j�a�q���� m��w��3EC��H{�WJw��կi|��UOS�)15����n�i����������n��b]SW�wyd��u�_'^$���z�)7���V�0xUY��+��u`��L3�
KO!���^�Z�Ĥ��0�׸��U��U�˻�����r?���>������T�TmT��4�����I�j��k8�������V]bJ���o�:8��E�!M�U���;�Q����S�1L��f;��oH3��1A��V�%�­c<��)��D5�v�%5ь4*p�����y�ȇ|�'��}�(gbo�&(I�.�g �W<:e�+�r�f�0d�[���3U��M���0��F >9֖�8$��{�a�^�JJ�VU �j��niF�%�F�@*`��h�L�y.�͙�0�ῶ�WW�{���M��vo±1Y69t�޽��B����2s{9ת�G6��y3�oD�}�*˧e�>@i'Y��$+@���Tk�d�����]F�*վ�[�0��z�&Kc����W��e�	<�&��j�Ԭ��G�(6ܙ&`lN�4ay�ھWI�;`ˮvtp�zV�m"%���W>h�tw%(�Κ(�);�鲘�Bw6�Gu4D�I�R�Ր�]�^ټ���s�f{�1��Y��J5+6MWCf�6f�#o��c�����9���^�=,���W�p	1=�l��qyF��6:#Bu������Sb����&d�Ǖ�&�9Qf�/TP�W�8�W�`U�-��.V*�WK�N�\&b����fc�d��
*[q���v�
�R�E\�}�ݕy� @ɳZ�S��0���Y�k�3o��ʙ�[i�ˋvWw#��BM��Y�d������؎ï6������Ҏg��^ee�ygf,YO��+����$ɓ�):ܕmڛ+CLnz��uk�+8{��1���C�蘣5Uڙ��3��� �k��s!@�J�E��|��!1T;���|������M��SL��g�����ݢm�?v�Q�M�� ��bs�W��³0����&�)$��$9TAH,V�
ATAH)�]H�o���p����H)�	�) � �~e0����;Z��{�I ��$c%$��ʣ�
H) ��� ���RTA~@�� �����4AH(i�e�=˹>�S�D��R
A
Aau�$�UR
AH)>B�:��
AH)��w7�
AH)���Ă0�
H) �7TC*�) � �����w��������*���R
AHe{��'���
AHr���R
AH"AH) �*���S�@ZAH"II �����v�i�.�������>JH(z薐Y4��Q)
H,� �9TAH) ��b�S��RTII ��
H_��F������RAHv����Ii � ���]}P7�AH) ��$�/]��O��
AHg3�{�RAH) � �RRAH]Q�
b=`P�R
A@������bJH) �=��th��PR)��Hr���_��R��s0��R
CUD��P?%$$��-���Rַ���)1
C�) � ��RZAH(f��� ���D��Sh�RT�S�$���o��뺽�z�?���w�6嫔�����/&��h�.ĝl����Z�;gn�۹f�	�^V6�be�e��
AH)���� �:�AH"AH) �.���S�~B�TA
AH,>RC߻ߝ삐R
~@��$~�Ii �5Tq�
AH/�T
AH(JHn�<���v�X[
H}z�&�)<�!����T�gn�)�[H)J�i���i!��
AH) �s��c�$���{�V�%$���{G��ܔo:�RM$>Iˢ
AH) ��0����I� ���R罣@bRAH)!��
At����RP�R
AH)� ��n�R
A��ZAH)!��pmR�fQCv�]f� ���D��R
AHUQ ���FM����T��� �>i ���-!�O��h��Ф��R� ���;��~7e��M]@��B��J
AH)�h�O�Ru��R
AH"A`5T��) �>��{������R%��D��R
ACݢk(����aI�愂�R
AHj�:$��$�����F�) �꧘RC��As��
A� �����;ꖐRUR�R
AH)��u��)�) � ���Pu�����Q ���D�Ì)1�>JHj���R
AHn�j��ř�\�fSYyF�)$��(Hv���X�^$�') ���ʩ5���R
AH~��) ����Hw��ս�Rb�R
A=�nLH)!��
AH)�o�=\aI��� �/��i ��{�h�~II�M$M��D��Rb�D��X_�5�����a����Q ��) � ���i �?s���d��R
A
AH):�$.������ �̔�D���Q�
@�RC*�H��
H)!�_?Q�?%$�ܰĂ�Y)�tAH) ���$;TC�y�$�� ���H)H,��
Ag̚�����G,V�����p��R
AH"AH. {��y����Z�1��`�R
A9�ޯ�_>�{>��R
AHn��������ik�Ѡ��1 ��U�Q ��B��@����
H/���� �N��
A�JH) �+=����R
AO S'�P�R
AH)� ��B�
�@� �������v�%��$���u4AH)+�o��p!��-%��R
A��
AH)� ����C�=��ϻFn��޾��w�ת����l�R���*$߮h$	O�cS2 �`�K^];ƙ�:sڈ,^x�?i.�#B����z���
��"$��׾����8��ז��RAd�) ����R
�MeR
Af2S�$���RU?2RAH)!�k��o���9Y� ���Y?3�D��j� ���Ĥ��RU%2�
q���P�JH)��P��{���W�R
AH) ���- ���H5D���H���ZAa�
H)U�Pq%=@�~�h~���:�&~���� |���@���z�ɶI�L��{���2Ja	i� �HpBZ�$�W� ;��wD-�!��dB�Hr��ѻ�G���eSF�7]�7	����zfy4Z�Wn�]�d�;��L�;c[���r��RII��� ��!��
Aa��Xi��.��S�$��䔐RՍ�H_�� ���������)��䴂�HbJH) �l]Xm�$m��
IL�� �����w�
ACI) �o�R�
A`~i �Ԝ� �aI ���P<��ʠ��ɉ ��
Hg5��d�����{�۳��\Ө� ���R
CUD��RTAH)�Qi ���Y����^�AI��-�) ���X���B��n�UD���Sl
H) ����.���I �;���l�k
\2��3R
AH)�R����R
AH)!uR,R
AH) �N2�|�o߫� ���Y4�a�
g;�r�JH)!ʢ
��8�M�m���R
AHj����) �9�o���Ԥ��R%�N�Z`RAH(i%$��q�3�%0-�ԟ�I ���X�H)!��{w�
AH)��Y ���R� ���^�) ���䤞CWAĔ�Xq�$����4Avþ�y��R
AHeQ �`RAC��:z�0��u ���R� �P��R
AH)!���),�F	eU����R
AH) �ީ-��$�UR0���Y2�) ��UR
Aa�v����^��)6�$�2[;tAg)? RAH)��-������Q��)�����P����D�ϙ>�9����RAH) ���I!�D��^��k��~��H,
i ���P����J`SI �>��Ӡ-)'P�*薏��D>� ���R
C�
AH)� �� o�ZAB�RAH)!z�^�AI���H���ܞe$��R
C�
AH)�l��ì)6�H���Q���X[
H~��|V�XᙙV�f^h��R
b$9TAH,� ���R:�L����/]�~�ܛֶs�N$��R��I ��_����) �O�I�d�L
H)UP>Jt����H)!uD�U���H)!�_�րQH,��L��j�) �4$���X{uH)UXf��P4��P���R
AH{[����
AH)UR
A`SI!uD��Rd�RAH(������+_Hn���RaI
�>ր������1%$�*�,�%$��{D���R�Y�u%��Rq��S�$��R
AH/�N{���*�0�����>�JH)!UD��X�ZAHj���R
C�D��R
%$2���Y>�Ka���e��9���d��H)!�3|�1 ���R
AH)��� ���R�r����k>������R�on�AI�h- ��RAH)��
�WD����\1 ���R
AHj�)%8��Je$����� ��%&�)��ۢ
AH)���r삐R
B��)>�h�E���R
Ag̝�{���)3��R
AH) �>��Q �i��
AH) �.���R
AHt3�>�c�ƒ��|0PZ^��3n��aS�e7���c-b�yl��U꛻�qM���Ƽ`���a���/Jڟ���A���7n�_F�m�:l��P�l�vcv6��1������J�mv����,nk`�;�h�9�q���{9���\q�\3<V�
w>*���	�mpݎ����]�-��I\��R��pR��ܼ��g�v��E�c�[Z�v�f�!�ݼ�r�V�6�Z��Z��q���m�y^�юN�A�#�Wa���*����ԁUm�;X�'`��D5�۞T�bkZ"�]C���p!����E�(m\�&e7u��~ ���@����,����AH"AH) ��u&�w���I ��ƙ>e0r�N������Ĥ��R&�BAbȿ!�!�����Q�� �����<�a��ʠ?%$>� �?~�d�) ��N��6h��Rq
H,��*�4����߯�P�7���6�ƅ���>������Uv��Y�n���t�1-��:z�t��[�U�ue�wN]�h�z�x���O��d:����Q�:f��HS�kZu�}�y�׏_�QOY1�޾�R{��bc��N�탕!�罳g����u��+�<BD5l��[$�j���$(��4؇��o{@|���5)��r�N��h�Mn����T�[��4�0�Q��*I��EV+��Z(��p�k?h���*S�A��=��SlĶq��e�L��S|��ocb��퀷��‎l5���@���M`r�V/�Ծx��,�ڨ|̼��r��ݚz��4ƫ쮞��q�aZ�����)�h
��ͳ�,i��X>6��*��1H.?}��j�Օ�\�@"�Q0e����G\�����u�m�������а<m5�ә;���}��1�Ƥ��!lZ��ޭ��Rq1K��)�v��&���s�\Xy%:G�}xN��8W[.o_����&�4���4n�X��ku�v�nq����f�G.{\�w;57��78�6�U�en�G�
Lg޽�4�P��_�i�>����:�9A\�Hm)w�r�ڢz��gN��o��O���1�_=��!c<��������Ϯ�V��
J.>4=U6��]cƵ}�b��_u����b�o7y�0�j��</�D��ޏ]:;!�՝��Vk̏a�3:��k�g�3��`�u���td�p���J�O�*�=ܾ�COjz�y�����Ҧ��v��H[*���r�R?}r9[@Ӽ��i>�����@)�βe����}s*��Jy6�m��+�-���i{��1��Ү����Y���w��"�����{��C�����|���z=Z�(��b��}O�y>��-�|���&>d���V��u&�N3�:�P�e>��P��ֆ���.�_�l�&��?v�]Ǜ�v�S�w<���]O'Xy�Ti���cT�z2]�>�q���Qi�����8��1��>�wN:�ް+�;��}D^��֚�o�,k�y�^}�q^*jڄݣ�83߹D��?}�d<�7��S������K35���^*S�60~�&}�S��x�,����<d.���T�j�{m�����/���P�����w[γY;����i�YY�+Ek�ĵ��Q�x�U��r���G$񇝮�\�bݺ<��Ֆ� ���on����C^c\D�~�oRu��LCJL���o��}��&eL��i��{zm���Ǚts|��I�uo��޲�Pě��qX��k��5�_2�)���ǐ�Ja��ύ��u�l�����\49�
I�T�����}��L�2���^ឩJ��,����s���'{�sΘm'��o��h���z=���� ��C�_q�|��U���`ەwY��q��J}t|�����뵠Ӷp�[n��4�1��ه��+*����_��u�RY@]�5�+[�/	�FV��+F����i�wn�N�cۘ��ѫq��'���BT<6��M�k*�ެst~ʐ�7��nq�Hc�OSh��{{����=a�)�=�ʧU�����lN�Ŷ�m(��Zjg/}�8x���>�޷�+ V���EU�*-ꡮk�3�Κ�8酸^V0���N�w�)�N�M!�w~��
�%!��ݽKC�7�\�꠾~���[r����2�'�c�J�c��SL8����h��PUxl���>�����s��������PZ�#�}@�=��W7s����P(c�z�R���4�am�e꩏�iXX=�x~��AE
�M�¸;^��n��ٮ���
O��/&�� �\=���1�@h���E����Z�l���}�8���U��k�#�>L����t�0��g��яv��M'�en �i�5a��Y�'�-�*	6u���ݮ��u_	�z�<�U6���SHi���ӕWn�-�3��#���n��
f��/�W��;{���3W|�S��ڝf�Z�MN��d�-���Z��a�}�s΍���1�����6��_�[���L>/��+[W�F�k������+�<��%�(�U��@�K�q�5�V�˾��s��q=�QO!�Q�i��nW��:��{�ԷM�;�w�9����m����׷�}A�?Lqj���e��Q}��&��5Z>�cUJ��X��S�v�a8͡�-�^��~�[mV����y�~e�fv�&�GY�kٞ��玻R��$�>���ճ�j���!H}dx|��\�����6�<�����ҫ����\�hn�r �̂f����]��^K��}��%�3b�R�����$�-9R�w��R>�YS������*m���m5e�uʶ���ͅ��WF8�%��O%��־�)o)�Uh�1UU�~�IK���´a�}Z,}y��?Sh�*����l��l1:�H{Z�գh�Kg��>J5�>[�Z��Ȏ斳��V��;�q�tg��ݡ�:�I����-�fN�X��v��^.���l�G{��8��!�W~�j���T��,<�(�k�ߴJ�O2y���ԧs���oW����z�wZ�7D�1XSy��VW�Ri]��}�z캾�Ĵ���r����]�pO�P�m9��!nһ�9��fZm'Xy�,�w������1-����s�)�gȣt���!^�wZ�6�u3�<��Y[����n�N��vmoMX��0��ڏO�}_�O�>�u�z�y�g+vq!��m��_}B�N�9]IN������t��Q�k9���'v���^v��y>�}���ٓ�Ӵ�/�Q�Z�����媾V��O����ws��=?��ؽ��o3�k�ic����Km��2��G�eS%#_1\Q���Va�{w���Xu;�_��SǾ����[����'��n�s�F�W����z�a��0cN�Q�E6����I�;���3MAz`�}�Z{�La�Pq9�;y�a�M�h�k0���L���+;��G��R[䖏����m)̻�ai)�j����{9�1��IK�t�������&tqe�9��H���ɚ+��2��<r�X=�&׎�p�uv�l���)��
h.��Y�kn����bN$�|��]��\W����;���1�������s&ܤF|&y��u��iH	cQ�6`C��W"�]���L�q�r��l�M�E]�Sy��g	��mC=��Ƒ\s!����<|&�ݳW2�=���;s�mݓp�S�ݎ-�x�g���{u�Hy�[k�#F�����ݦ��P��k�9�����e6J��)!�p��e8�"g]a�DF�nE��Ƹ����ܼK+���N�y�t������YG�`���LC�e�C?P~~M8����ѵLx�մ����]g>(�o|�׸s��c9B�C��!��_���줯�"����ɷL�|�5zd�߯��!�d�VQL�z��]�U�vX�^`�$���[ֽRm��߯G�H*k��/��6���ܯY�Мz�k|�r�3�(w>��O!�n���o���Jz!�<���~�ܩ�8�Y��p��q�]�~��؇��>��&�K-�CLr��{��Gڣ��I��i��{��a�<�UVdUL}Y�X�����C�<��̺��9d�R{_뗶���uÌ�!�G�z8\1���{���2�8�������Rn��EDHQ��/���>�@W���s���r�V��2��}[>I��M��oVk���(o���r�gY8���e3>�~tt�P�q�44���=yv�x5�z�F���0�����WA��N^�����U�Va�r�2�!��������M��
U�ǘ��C=�^��}PUr<����)�3�_�K4��_Rs�l�I��@�_Þ�h̢��r�]'.���a���.n�庇�M���$�lPQ�B��z�����j�ʶ�H��θ.ٹn�!��rH�2�kN>��k��*�M�?������PP�j[�ɉ���;|N�i:��&W�{u'��z�͚
w�����w݇�M��$߹{N?'�Y��f��@c��m%���˲�B���/D4���v,hx�2��{���M2MX�MJܤc�K�0���"�pV�84d�DV��^�Jݱ/��sv���'ˤ$��I#�U���ަ�Hr�������C�s�tŅ�w��������U�[|�7��
F���
�M�E��Lyړ��Z�sw_km�n�ϹF���)\k..J[ʼ�q8͉3*�N0�|�{[�:�ޣo;Jm�v�ӏX}�o	�uQ�}�]�<���٦b��R����6ϝ$�U'��ֹQ7�8�LB��4�;�瓔(�E��w�b�c�����٭l�w���i�.���[�6��8�TR��c��:�8�W^`[j8�z���C�����c��-V�������~gR^�_��Ӌ��/qf��#�T6X��GC�2(�����M5��D��go����8�x���ۚ���*�m�o1��!��>A���S���)�۰�g�c6�Nj�'5R��:�~�ڡ�ތ�N���ZI���L�y��ݝ��On��/�����v��H��ɥ���N��ǻ���!׌Ĵ����8ͳ7D�5ûÉ�|�����;TEǨ�I�L��}��}�����V���3�Ps��]ʊut��n�1���7yUkyN[�v��c9�z��ء�1���~��/�|�[~5���=�o��m6�m����4�8T�E�l<����}u�V�u8��f��Kg���y�j�g2i9�����P�}��g��}L`����v�!!Ynb�Y���,�Ȧө�����I��Y�+TSz*n��RR��~t�E�����i\ssm�*+����n����Dw�R�B�0��gDGG)X���׹�nHYYԒ�Qk6���گ��,��3����W����B�{��f��=a�c��}�r�]B���q<���؅I%��5�7���y37�W�>���̪��|��R'��ˇ��n�r�v�M������7��N%�ͥ�}J�01����U�����ׁP���m�5�F�~p�V�Kh�����Hm���˾g���z�xUV��˭��+qd�Ϭ�����S�۽�i��q��:���;dj�Kf��3��V�3��?QÜ�m������o���OePH*�D��v��=���s��v��T�ǋ=v���������>�s�Ld�8�c�ך턕��cCK=f�^g޽L`��ɤ���[����'��)�B��-�����+|��h�{�C�F�6��'}��o�����[��
L��*�y����[���^�hjژ��z���]��g>�gO0�s��CWS���W��%%�Ze��>l�.=�U�{����UU�~��vdv����5�輪�k��|½˚J6P.��>�֩��],���&�P�s��i�|�%=׷�A��þ�f���lǎ7�\8�|��{��ѭ���P��-�Z���h�r���0�+�s��8�=~w�
�ٕ˓��ލW��3� =%��ў���]\�ߟ�m��n�����v��9rJ�4G�A��������:��U�Đ�Z�h�a������[��<�閥���P�ҪsS���3��νz�fi��:=|�1�q�K��]�h*d��J�Z�o�K�\��Z3�U�����ĝ��0�wܺ:U7��q� D����4�}m�I��{{��}0���3_y� D��j�w�}�/Y+���>M�'�4����h��)-���_$��+�'Z��;�]'ɦw�?j}�e�"J����8�􉉃��2f�9��G��cgK������e^Ⱥ1�Ks�����UB��Ul�\�,תk�!&��E�������Ql}y��:�V{���i�3�r�a��y;�y��V}��m�^����ZN��Q�wte�����auT�*JO%���>��6V�-���&�&����M�$����@o�gW^h���g�)�>�+/�^�GU;�4��L������޽�̂�6�} P��|>�˷�6+��ou�����`�\<>��x��t���d�H�����F�^�X��6��ܝx��>a��5���*uz߹��7��1���&x�U���ZZ|��;y�!l�l�����?s�s��>����e>C/[w��|��j�^e�z�񕮢>���+�r����[�(��H�*"���s�+~�4K�[�����$�w�U�����B���ר�~�1������޹�|�f0�޵e?]i��#0Mѱk
*P��^��C���l�>��N���o���/;Zx�%�dJ��sEx/g���8J�>��LTUDT���NU5/i���T�}`.NS�^�m�>�a����/�Ny���O�;݁֡��[83=sv��O�ѦR�W ���o%��VdR�ނ��յ�syY�A�iY&.�V�Tf�w��9v.�.�t�"w���[k���:��d��owA,��ĮYۣ������3+,�3[���m�:gD�K]�s'{l A����t�]J����}z;���ËfX�5�+w�e˘���3F� F[~<�����)z��C�JU��kE&+�W�}�� +<Ew���0�ͭ�1R��eN�Q��N�P�Q�󮱎�����n[W��;����P�����WMɪ�tl�s��a�f�u�o!������g{:��r	�S�"O�k�.�tf�9]�R��k��7C�ob��t�l�x�T.��m�VB��
��;i�Y��^��+ɤ�1��k�K��ܑ��5��E�k@���ďoik�0*sm�C:�
�Ly,�՛���v��V���9M��36�Z�:=�h4T��f��9�M��wj;�)T��W�#ׄ��^�0�m"i��Nlm�6��m�
̀7��}Ho�hT���x�*m ߴ,�8��x����f���&�l�ю^,'��X�؍�;"�1�u<����dP�淮��_k�c#ϟUȺ�G@�S��X=���Lp[�^A�Md�ًtpe"2�.#::8v��6��)t��cr�w>��j*���n��Yn�T�i�|)]�o��a��7:�K؁�.��X�A�!$���%�j�$�l���)mv;m���0*�Uw�ۧ�+��x}�v6z�Fs��z�4�-����o:(㌟T��e�O�ۛ]�������]���ue�{
mdyy1鏳�����anu塃��9���ı��'���qG:��m�����]m�]�!���)�AtpuaGO�$_9�9���X�lyq�^G�X�7��sd��{=\���ZNͳX�Ӹ�Wɍ��@\
���ɷGeNM���c��:�^��W����O=ղ��V�Mj67Y�z˗A��.�gu;�[�Q���u�sE^_m�v1K�v�l��<!����5/�.����m����שy`.ۇ<�ܭ��j�(�GVݩ�Ǝ=����	ݮ�<x]��ybLݜ����vw6���YҠv��݋dV '"��4`/��DM�C�nl.�|L�H��<�]�\b�7bڛ���p��n���M�p���%�&��c��s�����]�N۞wc��6�l{�:�6�'fݻv3N#ՕwT1������G�gDٶ�)�˚̆� ܼ�̛b5�����n��ms���$��/H;��:yu�k�pm�]�Y9�E÷L��JۮxQpp���XnJ�2n�rm�,�\�����Wj�ydqEu�!�͓���nz�ڶ�!m؍�n��m��׍�<;=�-xt!ۊ����s���1�v Ӟ툸=b{f'�פ�5W;[v��[�1��vn�<�΃vzk��5��#�O�� �v��g��q�v�8z�̝n�J���s��vv�Ss�Ͳ��@��nN-�sp�ɵ�D���#��4s��nN��G>�,�g7>��sbHu�:}t��yB�e�v�rW�k#�nM��]g`��׷#�ݲ��k)���H9��m0vC���b���v�^�ή.����q�h���w,a�.L^�y��'H�d�{1dwAͭ��PY�	<�8�����-G.ɋ��
�n�H,t�m����GnNt{v��kkc�kFv�(�<q���S��g��:랰���20X�_\�67
7���fg�	�G#�0��n�^�E����w��z��t���Xݞe���TS���p��Xo.	�J3�649�<���Ԅ�j���>b�b�v7�X֫��s����Ʈ���Ge�Y�v(]�<'�m�4m]k�9���fS�hn�,�3-F)cm%i;�m����h�d�̮���=�9�ݦz����Ӓ�m�1��u�]=s�Ƃ �yk=��Wb��s��[�1���_�����_���m}��"�Z����A=UHV�>N�u�T�咽u��-4ͦ�w^��8���o�r��H���>�פ)۾oXiMU	��R;@"~xlQ�AT��"|�GBH�Bih�|�q�'�g�[�lUeB=�Uh�a�X���P�]a6<��ƙ��<�fj�8�{���[6�۲m-S]���KE>���IN�S-yA��[>��E��kyo�ϯf�ϒm:Ǐo�?s�:6�]��)A}�N�wP���n�ﳽ�N����`�vNe�Zw��������z��|���n��ꅡ�9�v����0Ӽ�3i+��{���,Ӷ�����zͤ���v��c`�[N���H��6��w�/��ﵣ��8�-����hz�f�Xϒ��ݠ=�~����ͳ�|�Xy8�&�Hm̭��[O0�-6�����k�>�(N��t����h��!�A]ʊr�x��9Uei����'Y�z�&�Zg�z��1w���d��~M�'��>"�5�a^x�Kսe�lU(m._~�/[�wy�޾�ށ[K���qq�H�ϥf�x`�h�h�J��DU��1��t�I����F՞.D����Ax佹���:�lEP���a�����[9Z�E�����,ǫ;׋Ԇ�;��g�Ҹ�74�v���\�ev�-��ɪs��G6�j�W��F�YB�O{�R~~����4��*�%�3�ЗY�X�,;�oX+�-ҙ�-�dE���V5.�4iv����n�93&ݭ����K
B��5�X)����w�K�^ɜ�߾U�{��3�h�Fߘ2J�c\���Yޣu����Yl�IB>!�h4����|.��*wh]�c�"i���ή�u�e��b��V�������7,�[�9og��w��+��2�F��3{��G=�N�[��5�Db��İ��.�`�f�f��`�8������{d��d����ޜ�r	�u�P��:��ҙ�U����A��;�kԭ��X���{5������yn�ĭ���J��Ǿu����;�?�דr���K���h�Y
���X�[�N��ܼ�9����De>��j)`^���޽���+��b�c�T)���.�����������ݾ4��Ys"�_�u�~4e�bU��.��N�I�x�#��w�J́mw����P#�/�f�s�K����5<�
ٞ
{Hq��y���*I���=��(����U����V�s\߿o����������>��L��y�I���>U�UĐ3�m��ehW��$EV\�\�-Go���>�tk�]Mp�w��� ����8%��c=�J��;�ۈk�񋊝�v ��Xt	m�w�L d��*�;2���k�(�e�^��ܟ{��v��6�>��[�YB����2���2����7ܛ��w��E셬`�a5���n��M.M�q�h_>2��o^c���9ػZ��pQOf�S�I��U��^U�|��$��wZr&�6��A��"?�M��<طC�y��b2v���v�O7*�����t�cb�csl,����L����<�M=.�⽈E�Su�Kh��g:~t� ��o�Є��|�qw^�w�o�5����AQ�J�� I���g+N>��t���J/^-ג�گ�@�<$ͅ�%�#鋬BV�w��őE�s,:��z79;��x��wlB(
�L���'�ZyZ�:��<��Xګ����Y��Ό����������& U1�����l����֙� ﺂ��
��R��󡼻�ns;M��e{)��{+@�GP8����ZN��W��ɣ6t�ӯ];D(G��V{��z��W��]�v*�8�%cGq��Lhi�I�F�J�Q3#�Cu��={u��O+��X\8��v.��Y*�onZ�����=o�5�ge����	Cw���ݍY�z�^�C*H���1/=Sf<�M��K��y��N����粮FӭΎ��j���8�cq�xlN�)wSۮ,7��8��cGt�uI�J*G��I��]�vJ��{�Eߊ�^9�ko4z	�5�w�/7o!���C�u
c11�`��gpn:��]׶�{�M h �K�q8���)�jS*��u�����{Re]$J��MC���V��
{�zci�W�k��;0�U��n�B�k)3���65	|��Gr�`����v�xZ�=8�<�w��}6ի�ʕs������P����<��E��� ��yՃk�b�Fb��u_׏Ȇ���2�Ќ�s�݅��c����~�}�����Nv�aN�$8�\��@���,ĸmG���Q������y�ƅ��0���Ѷ���}Y�N�o��{��f�{�Z��EA��$������*Ͱ#�Ǔ���6���g
Y�U̬������Vv�R�"��p3�(m�J�
}�z�o]�N{��E$R�	h��H8��m��ses�k�l�y�l�գ�U��A![�9�#��hr�nQ�S��.�nm��ץ�}m�ۻ7q��l��mf;N��6�y�c.&Nu�=��E������ٸ��-�lp����u��a;����i�ns�x��u��C�)�;oe�;9\��@t64���j�ݎP�\�]d��9i:ڸJ�7]�&s�۳�Û��A����R��!`ɶ���oW6ݎ8�rn���غ��5��tMֈ���w���U��s��qL̒%�%ܔ��S&l�%�(���s�߾���PqtP��{k�O/��6��J[��rV���:D��A�k�;g�!�zcai��ۈ���݊f��z}�=�������1̆eI؍��Z�6�㽨;I�5���@"�N���y�T]�/�n��L#�,�)TH��ʷ73Gmx��ۦ��ƾoR�]L������Q�t|4�tW�N�?���[�=�c_%�כ�#g���^r�Wy��)p�f\'Z�Ы޻����1�iK�'����/.p��x&<��rZW\� �Q�}�+}��(S�Z�T�*��Pd����|5�������Y�gt���{<�H1�}�=z��=�y�Y�}O�;��SG��=�����ݟ<
8�n�̎Y���wRs<�P�k���nE�p[X�L����?�F��x<}wn��CZ�Ӝ�0����^���^����1�:�u���N�u��#��e'�����ī�>�4�;SN�Feퟱ`�M��w(�6��]�gn�@�מ�ZpF�.��ǀ�r�t�{��]�\�[9|K�#v�.����v�S�����ɷg�E���/�躗-tg��V��igɹϸ�B&��#�;�X�d��9l��Ԏ{sf,����L��*%&��4�6)�$wn��t���=��=��p���v`j�_+��Z7T4o����v�����@-�f=�k�|w��l�B����ΡjP��()���̶.�xwK�e�gw������o��f�v�{Gr�ڎ���ޮ���إ��t��Uqt�)��ߧ�㻽���'V}.=k��U��[�v�|�~�A�R���N0A�v���v̌���痷��xT��ޡ����u�N��`�2IFnm�;<v����\�gρg�AF,E�l�흮7qE��,�b���z�8�7��<�ER��k�^#��y�.;SN��c3+�^8 �^/��VT��w�9 ���f
����:7�=ʅ~�O�A�)�PXl�:;<�g�^���s!)���3�\>ը1�Ja�.���*��4e��ٰ��~�t$ 2n����Mv��Y�w��X���k���q���~�E�[�zz⼞�kn�/*)xC��>��!��S����R^�AmV�5{�AYB���}�X�*�
�Z�<*W�6�`Iɵ��k���9���N.�z8kS��� �i�J���7�U����E�Q芈i�D�i�z�R��G_�겺��y������Y����N��u����,:�8�x?1IJ`'�b{=�Y�(a?/e0:�.D����L8��Y�;���9zq�j�r�ۺ��f��B���~�T���v_x��..@5���s�z�Ѯ���P�u��%�޲V^��;+)s��������D��c�.j��O�z͠��OV���Һ.����ޏ��(s�\\���K��
�fpndv�y��YC8�5�kew����-����� T�WX����{�S7�9����|�a{@��{���Ps��5.�l�nKn[��7���_�٨�%�0n�������j�o#rWB�4h��aTF��K�J���W�K��4^\�w��n�J�V�m�_�oiY�(���lV����J4<��aR1��kKm^I��js\�5{}�B����i��e�������b�������7�ޑ^�z�hu�3���+�� �^S��P{�m��9���T���k�w�Kas��G�3[����ԫuϸ4����o�3![���/�[:��nر�Y��m�CM\���l�߆]�wXK�&��y��L�-az;��J���vg	U�D��nyſ�QBV��#����u�4	ؖ���K�[�b-���f�y;=�q���H*�����W��� ����]��`ϳS|���xW#)9�;��.�|�©��v��ܞ���n�w!Tm��E���B�u,�9՚�}�H�E�B�+�^��E]߁n�-��d�����}^bX���A�欟h;Ĭ\����;	����^Qw��+�������u�ָ�{u�(��>�`Л�4���m��2����Y���#О����~J2�P��W���2ǳ��4��h�;����J��
ܿA��*�u �dn�*�I��g�*�W}��N�~�r��k=;�i���p�S�3�e�Fk��)��oJs<̨w������)|ic�����~���@�Ab�B�����е�~}1���+&�h���T��������.�ܐ��5P�v���4�J����d'�f�6�b��P@��f��5�u��Fw|�ݬ<4�ʚZ�y��Ʀ��X�}+��c�5�s9��2�"�+.�q���f�[��e�$u�±��-�Gn{v��yYܚ�:ܖ��S��Rjn�=����Y���i��yx	�lr%<�yZ5O>��k��P���M�ݹ�;�gbwNv��݃�q���ݣZ�qZ�n6�x��hٗ�N�3����ng�^s���5vq��/�q�ݎhENgv8�f\-��<;�v���n���Y:�<��0ŌRrഝ�����ڸ�;8�=��w[�:6{#��R8+asۍѸ��Q9�^��e��f�9XWm�����\�?,���Oך�y�����I�/�|�ޏ�6j8{�z��W�WS��86�Wv��x����b����6F��݂�L�F��o�7�"j�q���}�yS����+#G�w�B�C�I~Οz͑4�T7Ώ������*Ｒ�sÅڻ/�ߟ��7�Z��R �������¼�c��0[�����<����[��uE*}H��l��7�*yo����M5J���*�w�s�ݵ^F��������0��\{���u�Y��X�uO�{��T�usw�}Ǝ�j*D�G
���4�3(�cw��*N��v���Ɓ��D"�N�=�LSNB�ׯ�����g�}�����A�R��s����Y������W���b�}�}����'����'�r}����L�Q��m��K�I�[EYFlR�� D{RNs	�>ƼnV�1V��L�L�Mt�GIjaVβg��vyS�IT1����.�ӽY��:���Y����쑬���g�ѱ��T�=��z�)�v���
��(��WW`��^f�9k���hHk�����wQJ�nghu��+����坍@͐�֝����K+�S�0��7L��QYcO�����%Y�w��P��&�z���$MHw��ƵbT����r�"��z���gV�u�o�L���1V	�-֊�E�z`��ݭ��������N�{+����D��=��;��d��X�+�dسW��������VJ&Ôw9� ��TI���%ך�n9FSUoޔ��xv�`��fG���C�B�׼�y�t"f�,�c������pWG*z{���J�^��K��H�)֩�_�WIe4��>����0șW���)��[ꜯ�}Mk:#�k�K죬������th�S��h&�z�����s6���k�R��?�t�?�	ѱ�i���k��$Z�ݻvv����d��U���H@�/���uv(�IW[����W����Ytg���:��G>�/K��y��Q�.S�j���*��k4.5��ϑ�J�I�n�+��ï%��}���,�g��*��/h���ګҳGO�X�Wٺ�#!��U�o09��ܱ\�>ӣ�i��X�W�u&��|ܖc��݉�,\ܛ*l��n�gt��p���;h�'��#U\j�/|]O${V{����`-U�5��t����t�+|�e���5X	Z���ܱ%�,��vl�w�f��ݷ��My�z-���3(�ʞ�8B�t_Pr�-��t&u^���N��R�}̚8c���;gt�p���H\�w%���C���t��룷e�l�Z*Q*s�����~^�z�5��\�m
ώ�¶�s�8q���ޥ�v^�;3k�س�O���YޭE�A��6���� �W�t�k����l���	�[��x��e ;�:]L�fH��XΦi�Ul:�4%ա_Vc�M�n�� 2���4�5R$��]Y��p�.����:؃����GP"�[�ۯc��`�ג��<y`Φ�DC�ϊs���17E�Z�a;3b�]E]��f�7-�� �4�LO����mٗf�L�˾	��hZמ����f$��l�|��/��l�}v�lkB��&��2�UŉE:|�WC�%v֔�{�-��VYU<kT��|�Z!`���r�j-��Qٚb��G36���t�=���坲�wd^;Q\�L�0K�a���v��tƐ�Z8�`Q�u�R�E�[��	�y�Y�������xV)�Z��]��^��Ѓq;�Y�=�0&���eH������wr�i6u��c�wa!�f����4�|�������������w!�aU�c���;׻�푰���v�eH�}�*���A<��Ժ��k9�9�l�������[����J	��7I���s��b�����=�+�k����u�s�B)M����er_+~��w]�=5�4���`�u����%d:��,[�yq�����NZ]��w��-y����/���i\���`Ǎy
�Oˎ'�%J-n�Q���n_�(h�an�.;b�tw�)�뼏? ��]F���Vy�s\���ۭ���k���ѷj�'�|ӡ��������?K��*���]�ڜ�\�vދ�t�1���^v��Ƨ�J������J�o�ۺ*��*�K4C�fT�|En	��P�։Z��6;E�S��Z5��]߽�>�zo,�/Us�Ө�L���QYA�O���>0!b��ٕ/��p&ܺ�+��n¥�D���Z2����O86��L�\5���y7ښhk�昚�Ͱ7�cW{������*V�n��!���Ǉ��{�7˫ˋ���)g��h���sX�uP.���Uy�����_���Q�^3�+����^p*ŏy�k^m��
Ѫ��W8�J�c�H�LE����6�$����Uƻru.�K(�{L	�6]lʄ����]ѝ�u�Ы-���c}���<�ח�:Cc���������yx��
�~]���VH:�	E�Sn���xc��8;P�+5�)	Oû�.�	���&W�{�*�^
#�O�J��99R<���eZ�XH�����m���K*4�
�i&]�by��/RK99��;7nv�n�ge��I�[n/cX�M#�M2z���	�P�]wR��;RƏ�L_�)�"cA�{��#;�5ξ�J���w"���U:�K�ں��z�E��G[:���]��em�Y���:��/d1��9�9��)\/���!�{r��K���,M����.����}[��x�q�np˿'=�<�]jϠ�u�|'cZ��C=[�z�s���S!���H�����S�E��`�;���f�)���w��J��[?|�˙��A<r�ˬ�e�� my��n��褝+�������4f���o���v�.U{�����hٍ�>�@̀{|�Suܴ��]��Њq�a��!�;����m�Yg!*��4 ^}�����9�rP��\���4E5>fd�+
��=s�;P^���c�9:({��Q1��L�u��=���3����u=��P^����$V�{X/��^Μ�K�Y]oa�n��]fm��RL�u/�иe�]�=��,�A�ʊ��qv�p�=��E�f�E�v��ы5v����l��{[�ܢ��um�6goWL]�ఙ;conP��+ebroD/#\I�q�΄��+��]�<�H;c�#����N��Ni`�!��{G������b�>{�w��o\q���M&��Y��oi�,B���Ρ�{j��'�x@���۞�?�?|�r`���5�G�����:�ur�q�cL��4�^y�Qt�� �m��}]9�!�FJ�!*�����Y~\���
���f�?=�z����~cptNk�Y/�{��U����.�,�β�v�z��Wr�77zU��f�)�]_��m�֤�~��sf���sk�}���%��}�:,oQ޳2�l_�|��޵�ӛ�s���̶�ے��W5a����#����6�>����>���
�i�����M��m%k�睼�r�\>�[��8�]�Q[t��yx�7+���}���:l{�tD��]���/|oܻP���⒮Z�PU��s��D-�Nx4M�dr뽡8�d�V{��-�טe}���������ez�|��o+˻�y�y��3Ft������*�x�N�@�:�5����ђ�'/yTTv�Z�\xW�޴ҵ}���^fJ)��ܧ�.�Y��g��+6Q��a�^_�6�`��&���9�'��b��l.�p�ƚ����\9�/7l�<۩�vl������ظ�	z�Y��߯��E�i����ų��������g��Wi�}����-�S��U�9���){����\��L-�|����B��!T��y�N8�j��y�y�UV�Oze�mCM1�T��|�VT�ل,dPQ�4^��ʿWe�k�e,�}�tm���}��8��]g�	Xץ�|�Ϋ���<�L���f�b@Nv�o����:��y
w�Q���Ty�)gI탅v`�~E}��EP�&�A��xDAh��[�4z�h����瞥Iv�9����fr�{7:�CT���}���RWM��[w�S�V�QjmЗ_i�w�D��u�\�+~qߖ!*�C.0�%l[*��7)�UM�E�Cw2�_pw���s�-p�ѥp낰S���Sh�R^,��i�8y��p��b�WWA
�t��c@O�\�n�tyfC9�*p�ު�3>���L�z�%��>޾�O���MSi}b���0������(/������]Xz8�l�{5p�"�ix�</2r�hU��� �	-�姧m����<S��B݌���c����N�h]Pu���o��41K-�0���p�����o�zV��K�P���m[�w��A&�B����g����>5<��c�gW>��ۮH&���J�i�G�g����8��{=��S�%���{�U�[��[����J}B���i��-T5a�����k9���Yl�l�z�����+{ʣt�Y�f��2��9�~_FǊPi��F�,�����[[�@/+k3r��l=y/���7{�㗹64�5�.1-�A!nj�F��u���gmL��ԇ݌��#� wt������YA�q��A���!�U�|sW��W;��8xW���u�Q�p���[�A>X�e��e���n縚51�B����Cb�Y����=��>�U^z���&�~��dr�n� #QiK��غ���e[��tǙV�>�u��z�zm_v���&Q����;����x���];�]7Uk�#:����˹z�e�>�����SH/��iK�����Nl4�^^	�˭ʏ]�m{f#W�j��9H�P�-L�ދ��/n��׋>����(}�F�~`*�~��#�t)zJ�j����!EI֫+>�w�3�X�!�tΎ5[�n8��Z�~�Z_�o*	}�s�N4f�0`{�+�4���F�w�}FV+}��*z:�mѿU"Mg�>��*K>��w��y3�X�)�
��&��%��Z)��yt`�yS�B��¹�ܫ��{��'­Ԛ��2�����8����.UZ�S��͇�W5��5����7d+��[+����̚���~�ٝ]a��yܛ��7��k�?Cs�r�]+�f�S.��{�����ƞ	���G
4�ci�L�ܜ�I�ڜ"aK!ZVj���&�ˌ�Ղ5P�	�j��6�'ٮ\B�u����x�ײ��ۅQI욬���5Ӕ3��:��<�]�0�2�4�(*�OV���O��gM{+�
xo9��)U��x�)�����X*
^!Za��3�l��������,��{�4�AE"�k��ή�v�۬���g#���j��4njz��w;�F%�;d�k~���xSe�&̛�m��/���I���}ґ�<~��L���� �uX5~�Vl���Y6�J���о�53�t�eG��\��CꝤ�DKK�.:�e}�F���.�2���&��Γ��*�d�*�|��3��+�ݗu<k�{�hR��Wl~���uͫ�������l>�0��������Vӛ��k�%uԿ����%}��T��M���=����N=����V��G*��%
W[�;+ݻ���>B=҈ҫU"��L�Z�wAqJ�l袥�=���n�Ъ�������uww p]Z颩�-s<��}2���,���m{��o+y7������=��w�OT��uZ�*vr�"U�(��V�4��#��j�/���)F5�sV{�����R�o=�8wv���E1Q�Y��z�^{N�eh�W4s��ݭu+Jm!�*e-Ն��ݼ*�����ɒ�p�l�+��StR���
4/��S�_�zU<��^˺��b�=I��H�MZ�\uV�c9�-�@\�PCHB�7#b �h�D*��ƇmZq�pV�OOn*���;n�-=�\��������"��:�]��*Ъ��		����s#�7]��cj�Z��8H2n��5��->s<Y��zmN��
��v{���۔^�H�nМ�.��P��]�d^\���3�Kc���@�n�1��>�_h��l�v�C�f˶0:Cos�\�N�&�*�r���.���ظ&v`�i�0�Ő��jƤ���y�ON]�������)�c�nRP1�=�=�US�k���^ʎ]4�]u�xׅ��͉��k9�,�O}�[� �rTɮWۭ�DU��E,��ڍ���ʗvҞ�R�>@V��fjBlʛ��燥eo���d5��M[�s�%U��ʯ+�Rn����u�[�}ʭ"%"w�a��^ń�c�UA{�HzT�������r�lQR�l�9G7Ş��M'�W�U�y�+|�W���y��ׅo��B�X^�]H��	IN�X�(�c}�D�sE���4���z��Y�Z!*����THy|� �L�Q��{�.�,�.nFe�Q5���=�k2�Щ�=k�(����4HD��ΙM����E��ܕ@oԗM�ߍ�ĚDZ�ÙYޟj�u�Ay�H�3,�6w,�"��}ͽ�S��^;��ǁ�(W(m׀��b^ 5��rh�����ֹv�b7L�z��:�9=Ηq�!�N7K@R�*�,Ͻ�w���S{N`�Vګs7{jS�-�'%
���%>����{�n��5��nQǷ�,yN	�u���u�"��	bZ(QZ�s/�ڙX(��V��� QyP��O��a��ȗ��M�6�-7\�]x�����Ρ3&Ǹe�n���o,&��1רbڣr�YֻH���Fx���R�	��Uw/��ϩG綷������L��߻�=�R�~7�*�X e��X����Y�>.����`�X�E
j�w�Q��e�Id��e*��x1�-���֛s���%���t��ӆ��&?������j���Ά �u�q���V-�g���h~Y�aŁ
�V�قu�/�	�b�k�>~�w�P��s���������ι�߉�D=���
�ת[؅mO�Z`��g>W���j����B{���;5�~it�&���n�=��}Ρ���ѳU�R#G�Н�o��V���O')Q�e�FY�||=t+E�9a"	s�J1]�v�le�b����gOV�;RqZ�&�'�F�;p�l��S
�UAE`��՛z���,V�%p���J�e����&*z������@e���ڋ;�d-��{�ݣ�nՉ�����X<D�ɣ�e5*�O+����@/g5>�yQ�<#ٷ�<-[��TP�Ѝ�f�}����S����i�G�Ц{�*�qǞ�G����ױH���l����H�����f誘������>�,!.��+
�T�'r�5!1�B����u�'��xou�ݢI��u��+f�忱5-�.Uwf��F�����]��������gX&$�h˯U7��溾������o�+c'�&���u��4F�8XZ�ism�������ƀG�_�i��+T:eĲ�v�<�C���Mj���tI���C���oۚ���<pS�ɏ�U�ZJ��"ZE$�kn�q�H3m������Uߐ���r+:��f6F{��ά�c��W�xh#�a�͹\˳��~Q�E0�t���{�{����s����z����:�s��!ۗN쓉��o� �&��J��XA�ι��&^��zUͥU	S����4��U�.��X�yD���t���7��g�_��Q��Y���\m���x��n�v��
���Y�M�h��͊��8"�J�:�G7�2���u�u�	Pruz��%F��G��ӝ���Ҝ5b�x�?��M�yx���i�c^m!�I��F�4R��qH��+K9p��z�[=
���#����1��߷�=��}�=�可̦>h�Z���^��/��4�e��W�����sO&Q���:��c=M:��T��C��:�T���|p�w*6 �޺�}bC�/�Ujӊ�{ޔ&�#T��5^�+�/X(����e(z��+OgEkn��1��$��k�
J��l6������ű���ρ��3]5�T<K�}����j.']�����Z\��^�	�=��2�V]K��#}���}}+��3=,G�,]nRח���x����U��TS8v煕j�8����o����yeB��[b�sc.���\�z;p7vw7l�9�����[���ӳ\>�����w{%u���^^=u�>۱ϵ�H�o{�:ư.r�:Բ�~�@��g-N[�*s�L�w�}�-#�	�Qkm.<�4kR{�Пh���2�y�h>Ն�Ky �֬-���4�ϧM�w��N��d���_e��h�w��\�՞��V������9$���]q�hk���=�*VA�N��_��>iYk�mϽ�9���!˲,���A)'�u`��Yʒ5���`��X�,�A� .���w��_o��[�|�޵�]�z�c��VN|'����B�n���J����­�/�vP�tUA4_.8����X�K>a�|���V*sX�J�?�_>L�?��߿~8���L��f��/������k������b��T���K�P��9�ܫ8�G�t<��M��仅�6|X�,ה+w=2��n�,2������}�u�bF��co�U��u�+76 ��۲U�~vAۧ�s���EQ�:�J �̣6(s�m�h�B9�/��҇J����A�H
T��d!LY��ND5yն*EpzT��lwR򮄙xI��ㄻ7	��h�
T������4Ӗ��k[�����dx���S�DsV'�J�/��Oa+őO}V��fPG�^Y���j�^��i���0��ۊB��u6ͱӻF��p�p]��S@%q�"�"y>y[�3�A�w�kW�h�
���:lc�Do��M��>�:1j���7��@�3�3^�8�[�T�:*�{rr���-ȆY+
��oѿF����Щ�z�*�/jG)mڍNՠd����~��Y�Y�h|S�^��klY}�3�	��'V����P��E^��z/�����<6U��v�m�dEѮ�a�|�G=�/]����ӸV�W�%^��>���=�@��]�CZ)����BQ��T�T�&�X��
%Z���t�k, ݵ �^��j��w2����.�Ӭ�����x�W۔V6Pd�8�b�ՕH)1�� �:��aG�Z�*_�?�4�z+��e��x;�4��٫/<a^�*�F�1���B�!�P0�.��n�a���i��tjr�Ԉ����H<��+��/[�� @�f��T�.�W:8�E�PwLQ��43wK^���֙����ӗ+���x2�3��ٛ@U�I&�#L|�T� m(�����$�$&�k��М��&ɝG�<S�N�r��Þ2�.S�=u�\n���i	Б��۞���/n�p�k:��mϧ�$�-��Ɠ�38�Χ���b�t�\]���Od������"q���c���Wn��ma���u�۵�{3��<��85�A=�x� :x.+��щ�-�<�x��\���x�o)���뎷����N15��v��H&�㮦�����pV���
^�l�&��9l��;���փk�-!���먝��F�u�sq��3��v����Ƈ(m�'5p��l��K������u�Wm�6���mqrs��8�n�bzz�w�5�z��q�b{�y3���w��xQ�M;���=/�'Wmڹ�)����x!g^2hX÷7L�i�w@�l��;�U�w��vCf�;��p�s=��� 0�rg�σ�5�{��ͫ��:������z����tv���{����s�x��v��^0���D���Rvx�bŝq��ԁ\"�F�rAv�v�Uo%��۲+�`�n�ȯI|kG^	-V�vx-c��'l�=gN�5��ᷮ�vݗsQw`��E�ڕ��qqe�c��w��&t��g�W���5[����a����i-������ܡ�jL�
r\��-�!y����ܝ�]Hm��q��������ٷ`��<pu�wvk�I7��t�.&�㑃�k��=4ttF��t5�h�^P��nx����[��2�y��������8�qX7;]
mv��u�$,n��0t��d������t艠�nͱ���q�`��5g���$cs\�{7�2�%��m�/��7�n{a������n�y�\�������u���*�'��o\W��Z^��u�-�7m��f��b1�Ƶ�y��rq�f�%n��T8��.�(�-;cm��<�A�83�Ʈ�S���:���]\���>��"s��}�g4U9&���`�;���mLa�Z؟8�@��61��9�jEbfll�Ӭ�B�XcupT�x.^|��`}N������]���*<��&�{v���E7e^F\�m�l�qF�yx����T�C�il���3��'&�����7�onz�<����nkE��ۤ����.ەCQ�8ݣ�L�vP��ӻ-p����є&:$��GpW���M�;O�Y֋�nM�#]��Wj+YX�j+jb�+�X}쿓$�h���O�]�F��䮝yS��Z+�dg��
���W^�Y�_d1=��.���K��o{ҕ�{ovm��v��K~"�L%��=����]X�;��Y|ies�Ӻ��Ӕ��z���{��fS�v��^��_Euf�"��.�7B���O����}b~�֝����@��T)�M6.�z�A�V�5t��)x�>�U�-4��#��d���e"0wY���[7,����WA0_xT�b�<�ŝ|����L��iG-mǥ�{�K�sQ���b��̩���f��ޱFϲ���и���_��妕���t�i��f�&x!�dL��!��{��Gke$�M�J��)%��Y��m�m+��r��e�]�q+��)�8;�M�o,f����g��'�mg��ˢn��ŔM T�^^�S�J� 9jm[Aj .�\
bc!��`D�`qh�n��9ݼ&@�@r 4�;퐁W���VE�H%X�j�A�+O<�&����Ƿ)j�	^�%5��\����+=%9٪V�����X�YC9"G���E���}6�5y9��^jqƙ[0�U�wyn!�H�RY5Cua���om=�"� �+W̗Ld��Yû�
0e<�:\t��b���[�$(�����eR�����1��z�q��g�g3�V�K1Y3xV��̭�9^��FI��F����v�wLq�3z8�q�~�4��� ^%��=���5k��Q��+��AbX�*�wrϽS�U0�gov$y�s�VT�T/��xh�p���(��s�$G�y�}7���
�e�7��ג���+��Ui�4<��N�a�41or�W���L�q������Jf16y��gE�=Og�����ً��)�*f���j04�:TP��}���{���UpJ7Z��o��ofx��r�/���K��-�7\3ø��EvH�:N�Z�5� �ު�g��Ey|�r�B�Vz{U]�l�s��vk��.�{�����c�;ٳp��C���U'��8nrCY�z��G佽�������}�b�����Nw�1�2��۽^��4�����:�<{}��i>��B��y�٭AtPڡ\P�7�q�H�F��綵��������_;[�㲯O��=9����j(3T<�ܜܫ�>��+�����\���V՗j&Y#(�&��jx�۵�G�^	U��BYcn�����1��zj;~�FC ��W�o��c���S�Ig|�������]�KT��e'̊{n�W�XR/z�'v�++t)��ǈ���~�(���>�,͗+�wmB��]ʓD~9���	��1J���>��_����� T�K�ˬ2g��^�.鵛J���Ϧs�(�"����I��Ƴ*D�"��X�b�f��&U�����<�rdfإT�e	MMf�t�Lh���AW�Q�yϼ/�d�;�xO���fT��51c�wsѹ���-tu�L�������/�+u1J����A "10F���9�D�x�_68xn��j�G+����`�F��B>�(����>�~�~�,W�����F�*��yK��R�W��ހ�kD\I�Ψ}𼿞�7�A�u��l�Nk�Z����Q!B���(�H�^�9�9O�W-V��|�n���9������{��`]�u���O|��k|�;���4k�*�Tr�r 9c��ۛ�i�*Hɢ���N��fVz�ܺ'\y�R��:n�♕�:�6��[`j��l�OL��U
�Ǔ�_3�R�:���k��WX)��_sf>{��q9����?����i�[�{�]�[ֲ���>�TF6�5ݕ>BfGye�v6��O�%ݮ��������%�z'=���EؕbOnf>����[�n ���w��F�Iq��:9��ӖOEv�=XT�a��D�ńOW�f9��F�h�Vn��1���6��/�ҹT�����K(Y�O�ջW~�%^/=Iy����^j
v����L�c����k���XS�okF�m^���Ҩ�V�<d�B{q�F���3��c��ή�7n��A��*�ݍR���P6:[����XO����ۇ_�j��}��պ�ON�R��X�e.L��+���F�#��w�p��~��u���:�W�x�J:�1P��)G�|��<W���.G���n�}��:^���*�*sZ!�m��%�?b=�^c�m
����Z�z�>�;qj�oF����i�`�5�K�% XA����$>�S��>vlHi+�̸!��x�ޔ��i�s���a���������
zp���czB��ٔ�w�$~���r�	Wİ	F���G�&�̾4}��v��3'(I��up�qi8���+��m�D�ow�L}����(����ݎh��:��HS�Wv��R�Y�E��^��/��W*�}��2�٨5s�̆K��뱷p�R���:�L5V��/����h;��w�X��K�4@�Fs_:����s/|t��-oF�qWb�f�kl�{G(V@U�}o7�<�W�w6�U�}o��Άq׽���7�w"Ԝ�%�q�ode+
����֗u�������۲ (�euǐx����b��,��W=�yK���6$ǒ�t�<vV��L�z�u�hU��	�ݍͯk��g�=��v��=�E�3��7g���.<�]�ή)�%���M����m�����X��=�f��ۘ���z�e���oY^�9�m�۝m��θ3�
cq�[`�q<{3JE۝1�p���Ό�j�=<s1�Ӈm��u�^��ܻ���ܦ^:�TwTr�E�D��(� ��ŋ����ڗ�mP��+��*߸IS֟fy�f��M����*/?���^���x������k��Gh�v��򜛤�k�U����ֻ�Ë����l੧~�p�z+ �T�6j����R��:0QB���o����S�����L�u�		S����W�̙���9������je��]u�� ���:q?>ǔ��E��\�d�mL]�����T0�+ڍ�s'�p�Sh�q��;2�	H��_�2[SU
"蠁TRA%Wę�>sq�[m��{��7�;~V+k��Mt}6������>�➯;+
��>�>[IN�\;Ɛ���s-�fF�_%��J��(��$j���`��Ո�b���kn�\F�J�JZ~�6��הQy_'�+ҙ�9c���.�̷X�����{�X1���M���'�C$�+���%N��u���"����t&u�&z������������2}��ļgn��	A
D���)+�d���3���U�����7+4�_R��t��ug11Toʞ�"얨�F\�	ѬN�o��wN���Eߵ���2�:���g�ދ+f �Ό�6$;^�-jx|�k��&{Aٖu�c𬰹"�})M�{`q�H]������*)�y���ލ�J���1D1I��������'X�zgL��K�N-���a��O+�9��F�Rt�-�|0�K�\~^4G�����|Ʀ�oN^Y���]k���@�>�K���ǂ{@��t�Z�s��S&���w�ȴ���j��"���Z���ie*Ѩ{wO��=�Z����<,Q�S�s����E������I��I����7O׆|�}1�m֭��|G�Qg~�Z8,���o�k���+i�O��g�4�.�n�Ǽ����v|ŋ����5�^�t�J�����<	�-L��{���y��Sj-쎒^`�w��lgi��փ���/n�笄�Q(��_2J�9O&rg��z�m��CyۂCۂە,���w��r���rD�U*6�
�)^������0mm�4�ŚC�y�\�a����~��Qu��襩Jwg�.G��\�H&�z/۸�Ihg��nQ�ȱ@�*M6>i��(��������Σ�7Yf�BU�%"�}���������P��ϱ�����RyweM��}:���Q�:�x�g�{��j
���(�֫]=O-�1q�ղJ�k0�P��9�2b^J*��[bR�6kӍh��ӗC5\�����?d���W�>
V�E�S�s@
��k�q�aTpfW
�6M3�V`�C��ɪG�����d�唳���L��	Y9�O�gژ#��N� L �V��(����v��y_��w��-q�b�f�䏟���
O�&M�R��~l]��-&��Y�:��BJѕ���^�,�+Ů\�x�¿��|��#t��ȴW��jU�ޤ��:�V�<�N�:�/I���7�.�ow�]p������նJ��������X�n�C[��Sgu�qs����B>��X�).�^J-屵�ձi�u�$搃=��t<�^f;t�I>���������ʱ�=⹯T��ݍ����Q9L��jxR;r��k��i�9���϶��fV߷)���O�i59�Bu�[� �m
�th�^��^��i�����
w׶�z~yy�mP�����O�*]�`فx���ۃ�՝�xB��g���E�U{�ܜi�9T�2�z���_Ў�H'�=�L"�ge%�.�G������<�wj1�],@��ڋH7��Y�Y�fyx�
�H`����>��7}F��H��Z������ӽ��7i�.�.�j�ƾ�]����U�����T��������v�g����4T��(�6Z0�#겥�r��<�r���N*Mi�4�H�]�k�K�b��㖺�� �j�}t�/���L9�7��2���W.�EeZuX��PJF�[��g�kg�����}*Q�*��Z�f5���F����9;ՎQ&������,���7��\��ž�Tm`�YSq��AJ�[z�&G����]kl�F�;p�a�v��;;t�dnd��H����-�����q�g���.��WB������@yem�t{T�7J)W�����U�W�Q�WC�}��X���֗w#�_�~�T�QKX�J�1s�\�+����5�\�!�ەgږN���{*W_����U-�w� 4�o�M���R�j�z��D.�iw�i�'o�=��-�g�C�&$�;�cR�Ab���j���ey[Lva_Y0]ڝ'��{�ocԪd�5�+-2lu��Zx�y�Y��Eѿ�:Z�Ց��L#(P!SH�R��JJ���OnدoǱVy{)��T c4��yLĺH���W5~]�a�S(�Z�k!��7�rޫ�^�W�ux(�=4R��H4�W�gx|n]Q���y��{�Ճ|����1|}���>��+IB��U��ꕃ�
4{U^�X)�g0jkƎ��R�N�^��\�y{W�#/up�)
ѩ7�Z!,Qm>�&�y[;nɝcT5��W���H? �[��!�I�Ϳ;&��aU.�F_VT�0ot�$��� �b]���<��ػ�q�u8|�q�۴�h�gnN7kO8���z��s��xͭ�(�ŧ�9��v���>x�c�b�pm������>�v7Da����<<;=Hty�vӟs�Kƹ+t�C�t��ؐ�Ѭ�H���<�6������;a�;�V��T��K�����X����4��C�ɸw��S�hǅ:wa��WϬ���k �O'*�QWK�/<t�)�`Q�!��FI��s�o:Q�w�c�ʡ���=����K��Y%]w��*[�/�@�ϯ�/��.E�=Y֑^H��8ڒ=Y4�]��>�I����ذ���\�}�������ug����t���h�L�o�^��]����f��&�T{ج�;�`����`��1�s�g�o��]�N7A�\y<ռ�M�+�!X,|��u�jU�+�[�՟u{�u�=b�U���R���G_N:>�:^Wf��}���en��b�'t�k��YUr�_]��e���>(��Yu��g�^���wZ��r^�{�ڥ�C�M�]���kpfJW�E�y�XkwPʔ������n¶ �]}�;B��vnc��}�a;��'F>��=�y{Y��ש[X��X�n�l<�%���[M�a;;���(R#-��4�Lڽ�7��sQI{\q[Z��'ն��9�h8����q76&՗�wscXx?�TѢ[c�o�f��.#��ڧ��Jzh�*� }׷�}�aH�~h�u��ޥ�����Q�U�2�B�E�<���A }Fj�26��u�
�Zy�b>�2�*C�h�������nWt�1���*MT���C�h��jiW��q��l��k7����v.N��Gw�e=��8�܊i�M��_��y����R��6�@.��~��wB�n'�Yu]^��C�������Y�����}�R)(HJ]s�w�^F��2�^�L�f�M�vl#����j�9A{�J#2�>����b�����}�[��w�>˝^���@uD�N�J�+baY��
�1볕b���s�>"6����ᶞ���M�竷����4PgM>����^9������U
��	�����4��w�=��_�kմb��n�1�g�J���,w�ԏ̚b�B�}|�#��.yA{�t���+��b���j��`WO�YTPnJ슶ޡΈw[Ct �:ݺ��:Gn _b狦i5lA���(��9��_�6�����$Ɛ�»�����55�r(�ڝ�o��w��z�E#yB
c��US����;�兗������~�_���e��;^H��"��S����@报�}�w!�s���b����B��L�s\��85uOe�ȼǣ��{_8� ����?���{QS��,���wƱe���i����;��{��ԫ�^w�ˣ��W��Sk��S�
J&��e�v'Tѩ!*�2;+XD�\ٌMV�gge$:b���S��ȺNF%c��8(�4���0^�/�j�ԁ,=͒Ӄ��\�摓KX�Э��.�ї�nS#P�!6;{��4���Fr%2gf�VAt]db���D���K�\2�]�$¤wy�=��g��X����I�!�l�}�Nr9����֪�_�0[�l +kU���F]�"�V*кLk�8�4���ۥ	�V���9�\���r4��nd����ŏ��Wq��qS�E�qV6�e�p�Ġp��Q,��5Cj�;��[��6��B�m3��-�V��*�≋3^�Χ� ���v�nPoQ[R��ψ���0ZܼX�����j(��*eXn�R�a���R��y�j���VV�fL[���2@���z�1f׎b�:��uPC=R�mdaTX�;�Ւ�div6��SMCrʙֲ�7�]�����K/�����,�6�t�E��5�)��۳��mcr��4��7=7�g2�A �,4�J��2:��!IS'qEW �f����y�r�ڋ	�)�f��t(ѷ�^��e+���W�GL��.�qֺ�t�I���Z��Ťʄjn���[|Kݭ���ŗC�����e�Z�I&�/k({^S�0���ni�%[)�SU^V�z�2��[�g6�aT�7=�5𱩅&R�y`�H�4�\y*d]{R�K��%y�Č�L�{+b,G��G>�h.��f��9�X�\�P[53u˷u�0�J�����'�jЯWp�M�+n�`����Y];�^b��Lh�������i��y·�]��~�q��c�	VO�G��ܮ2�f(p��_Tf��>ɄCy�
^���/�$�`�7$�M-ǋ�=u~��r��� ����V}�)��7�y�,�� B���V�5�ook.�)
���;���z���~s�g��dS\,|���"���&�Z�%L��,Z�6�vywmv�:Ƅ��Cuug���xU�m˝܊�M�I�h S��rʓ�������z�Ҍ�=�[Q�!d�|iٺwv/��{L�S�ƶb��é�/)m���D�n�f�����!�F�i���:����+�K��T?9U�
��Y�ҥ���|Ǆ���S���&�5`��5����}�����'���U�ͽ,����Yʌx��4�d��)�8�C�ֱ��,��û(���j[�2�mz��Rŝ�F9)��w�ϛ}�r��%Uuw�w.5H�Bt�*ʿ7�%���c�D/�� +3\�>-y�:�[3���V�]g�1X*h4ׅ���R�]�!�@�w3v+��h�׺�q�AB[wl�7R^�~cok`��ww��k6yܰ�yfXd�������c2,����_�]+�E�T�{���5���l�h�M�)�[ &���A���;�O��0�#J��R�u��v�4d�������0|�<%ﯽjU�͆w�q��ayKs>��O��k
�,�u?����ψ�"���Zv8��Mǵ�m��N���{c��u�����t�<De�l�p�//?���z���i����n���In����q�_ѳ&F�m���o���*5�\�V�h̦�"�4�M+���k'��1q�k�� �z{��������e��u�bAU��n�Ѻ�ǲJ���(-�_n�a���Ey��tj
�1�6vye��.�uU�m��b�܎���@娔���u�]��r�T���K�~A�-�؜.���V�������8��hk:�Q�Us�תze�+�P97��(�2@�N��n��ޢ��<F�]Yg�؋��m�<r�L�������������n���rvU�j���~���G�R�Rh@4����yĘ'q���ۢ2�����uw+{�EfE�WB
g����(2�p�!j����o���V� [���y
�Ѐ�@�Q$��.mE�{-`b�(2��c�� �u�e��k�]�%WXa�yҋ.me[�.��ܘ�,F�r�zO��o�h<@MZ��,�)S�un�u=��ռ��{\Y��1�}�٤�����=�s��]b��"���9��r�u±��0��ְ��_m����:���L�Y6NW����&}�a��vM��'8^���q�Wi޺띁m�;�4n7c�5؊S������[@��+�Z�Yc�����9�jLope\ygM؜.����lf�������Z�c�먐2�a�Y���y�\�x�F#s�h����ݘQ-�G��`�R(�@���1�����=����+���<s�e�����Tj��;�����=(=N�H���_��
����ya&�c��^�����Yk�E(( ZWO�w�&�z�N�T���
�f�	�ͨo׻�n�SD�ܾ��;��a�X��t=���h��}Mh�z|�e����x%V J���ؕ{=�fJ�W�$6����?#ƯJ@yv8��=�ۺ��,׀�n_�hW�����g.�	��@E!;}����M�~4�-��4�;�~�v�V�w!~6�--:�ŵ(�P1����4�����"'�<e��r�{V�Z������۳��л�៾��Q��i�Sy���*		k���W�vZ���Iʽ���ޣ�O���|ٿ*��T}O)���� ��̚���:�:bF��	���G��~�
���%��譑�*Pgvۛ���E�ٺd�T�er���W��1���t&V�L����l��ÛW���i��Q�e�y:0��_nVڗ����(C�װrx��,gH��ʼ+����
�i�H�<�oąI*`4Ȕ���&���ȗ�΄]_�`����gĽ���6J�6��u%/.��t�慵�{ӡ�ct�	�nE ,gU��ܸ���μ-������:k�m��u�Y\��et�:�oйO�}�)YޜA���pno���uu܀?�a (�Ա��%d���<=��g����fiS*���)��Xj�U��^;�s�z���Em��Mɭ�/��C����Z4����j��s�ㄆi��i�Ω~��4y�ODf}�X]2�`��=�]{�ʾ2�!V'+��s�m��o0h''x�k��fPy��om8O���MW����~pD�u7<��co������۽�N��8�2�rަ7�xw�0R�(�J�e=��%�a�aw'��J|�5�m釞���r_!��+��s'��u�G�NwF#�M�y�;cn �n�t��/,pG�	�i���K���5M��kR��%D����^�Ҿn�r��y��ϯ-����$���XA�����<۲�7�f�Ƣo���z�+~��Ee�V}���]�K{��e�ݴ����viH�2ÞZi��z㮙�}���*�n��O�:�Ri���WBo�?o�g�v;�+Cr���럧7�s��w�%{�BdҶ�':,��G�[ ���2ӰG�:o����֖皖h�R<�*�k*�S�(�X���r���+�+�+�Fp�W[��egu���Ĭ'/8e��u�+ʐ�ee�)%<���.���ͻ���� �E*�HS��O Fj��m*�(�=�2W�*,���w��_m���·��F�mTU�G��ܞ>Ũ�@��ߺ�J����e�z\�{�٫���4��Ti*V���y}v���S��4�]��mb�.���ՂN��̶P���n���~�1�_ng'j����x�B�['A��J���۞�e�7u]��']��n��
��w}m�ɾ�{����M����kt.�>��z�R��5�ٍ�v�� ��P���O�E�v���
�OE�r��bpM����'y�C�sf��u1�d�Y��J��j���ϟct��{zT�+�-}A�}�~�=���s�]�~�U>^�,�<=��*B�����nv�+��kܜ�n��E(%���ަ��=0o���xeۊ��ƱFϣdv�Yj���LV�K�0������o��,����q����g�lz��#����P�[� ykt���g��iŢٟW�J����\��>�^7�=7���>��Uɐ!��ު�rX7�en��#���4�<K*P��u.�	iCJúСO5dQZRӖ�)��w�{;xw��z�f�1�N�������)$��[߷����½�N�W�7���^�[�r��[���}���Qnל��!���^�Έ�C�M}t�_�B T0j�h!x��}��{o�)��t�v���L�)���H�tUĢ*�%©0�B��~�!����{
?ƿ����K�ۢ*��b�~-�Rm�����m��.�wt��/Ֆxn<b�i��9c�a�b�Gs��}��qF������͏+�f��o�L�z]����=���/��c"���}�*�V"�����f���ow�#,��noz�X�%�7�g���߁$2��Q��U�Y��@U]�ss]g��y�#�q�N��b��/_z�{�A�9W��l�X��=eg�͙G�˷b���H�D &�Pm�*��~W<NW�ҁ$͛K����ٔ�&�p�����Rj=M7��+���_��:�����f��>�V��IQ�&Ong�]�ؼу> ��9��0�p��!/2�+�`�+77䊨9X߀��h�;c}|��7{*.�g�;�®�=�s8�}�n�n2�+����~t�jn=��S#����mb�
�Cv�$m=ŌB2?[
�7�H���RU��,wO2ș�'�e4�nf��W{:�%n2[%����S�wn{u��Ѷ�dy��g���v���SO͹�s�;�p�K��wQ�.�y�ڄ��nh���[��]/n]�J����7�p�f�b�V��Hk���Wn޻���f�G�.]���94Ly��J��*Xm̓���[<Ӟ���uuU�����D䱵��u�����:ح��s�m�k��z\\\N:쌡����9��M�nᓰ�p�:ۡ���B�v����z���*y�XO�I`����juu�n�<���u�u��/J��T�yR�e7��"�|����grgV<� ����Oo ���\zn5�x��L�GA����o��b�8�ywu[���Ÿik�y�5��@0X`l���~_)�B'-���zo������14;��Q�ͱ��׸�.)�im���'�����r�C�����ﶪ	�]O����*n��;��� *-U�ۜ G�'�Sk�vv��{z��*��1NF>I���>!'O��H���O��U�d�e����F�a�C垵(0����獪T��n�Z-�bM{��	8{6hׄ=�oٵ�ՠ�l�d�Tko�*<k�{��Y���f�l׫w��S^��9f�{����4o��xcU[:$g�{�z��裔��`��~�:e��:lY��v����f6nވ��D������,fF�6��i�`�v��-&��nq���@�o��Z�R+R��1q�g�&��`t�
 ���7�=�]���^�y���0�_=[D�򂴖�Th�����{0ؿ_S�c��ʳ�u_2c=ٍ]rpޥ��D�'�4�kG�g*��P�U�z��>F�:^���zWv�_Q�2�N��	���c���u�Ă�8*
�G�T���ZZ��/��Cʹ5���)���WmS�̨ʜS
��I]_u�/��h6���W�$�@C�����NE���� �X�k^( ���U�yTdG�旦`��VwX�򈞻�P�'D��4��z<Q��i4ZTL��������R�jʲ���ξ��{y]�2P��[�_Z��n���y>((,������3�l>�~t��z�˧N�RZw�4�0�jк�Z���dssw�;�,��t*�R��~z0��/x���7�
mx����o[��<)���{Z�]�:�G�J,D�dw�5���3O. ������A�8�f;p��eŞ7:S�5�ܺ8̂6�5	Q%�1�iE�ł�̢��cr�>$}y�u��n��ޙ��l.ӷ�~U�OQ캊��e%K=V�(��D]�%P@�f�M���.I\��~w�p�-�����mAN�`k��&��2��!�2�.�ފ�vfv/&��8���z��
�Uw�W%�.��u�R��,r��#mI\��;�t�I@��.���wR�no,mt������Dz�W��]��&��L;*A���;��E��ݠ����9�k�>�z�	���2�w�cs$��w��w�RǗ	�d9B�)b^	���M�����䐥n�6���4]�}�������2�Xkށ������|������m�����gfv�0���8c�I<����{MM����}�+�*$��`>��}�C�����L�{�4P�_G�LR�/��Z��ji�kg�G��o��yo%�Y�X"��������l�Z')ͅ�z�OU��^�zY���mn�f���Ƈ�F��X�m��t0��(��t�D��j����s{ͩyˬ̏�
30c��x�Wc��o_]C������/��Mb��a��l�t�7ȼ��0�>�~�Z�Z�R�A�K���6�b�[5^)]�G�:}�+���)�{u�o����٠J�VW�Fk-�Ҕ��������F��}W�?�X�y�Z��� W`�йE�1E�f����e̱�
;HDvc��R,��Ŝ�>�\�k��{�J�E���+w�j���b���дZ�_��{k���3GT�k�I��>_�G}��)�1��`�Fu��V�0���y���8�J�̝�|n�]�s�բ�k@�Y�$�J��L9�r����⣝�i4R�����N��}�	���_9��@��/K�$p���v��=�%���)�I6�G*�T�����p�z�������g�~�}�5�EA-��չ�v$@K�р>�J�5%��>��7� �qA&�EnW��+�X��D���QEd
���ks����r�oQ�|�v=����k�-a뮙+i�Ͻ��&����cGn�{Av���1el���ç�ef7O�wn��eh2�ό��wb�;J��]�Q�.���F�7��ĈIB�!��9���Ci%��p�wo�����~�Ւ0�[:k�b����C�+&eFB{�{ٯ������:[�}6�}�V�_Rd
):�{u���w�4���Q��JĢZ��V���%����^���}�+�ȷ�eJ��t8:b�rrY`�@�2�	�)6�2���,,LO��om��Ѣ�ǟY�\lu	�1�"�]X�����L�����,g�ɛ;�c�Z��4��,�^�V�n��$��/&h�Kh�I2�'����nv��Ln��I������Z�Z=(��q4�G��@ƯJ5a��D��nqs���a�z�xQ�(/j�Kc�7T����
c9V��T?v߭��t�z�C�d#�2��������lOP�`��f`U���,`���H�k�7qN+S�h�<E�����tR�w��jr���C\�y
�r�Z���Y�.@�Ηf-j����َ�%7tV�N���L�9}��{�/�̜�x�ū�M�Ҟ���\�#ݎ[���u�u�T%[5�^<�2R<ԸWIa�{�[�C�T)nmuW]����vh��a;)0e�3pFw��1ytt�}}ڦ�ŧ�Ʋin(𛞸���됋��1���8+=������fݚ�v�o�5�a���8iڍ�E��� ���]t
a:8:}����ǹ�F�l�0wd���l�Hl:��̚���7/-�Uh�*�|}�9��ܶ��N}s��/��N��^j��y�����4��wq#^��ĞA���o
��9qC�3 �r���؅L����3���"���\�`� Ǧ�G��9����dv.���|*Mزt�9j�Mx�%ޫ�v-<�R�kV��W����w>rLo�6�ZN�,�b`UqE}+i���ƕޱ)c���#/]JR�V����������4%X��:f�
�7GNW���̢Ǽ�c����B�� D Kl'�rJcp<{��1�������	��Σ�{���2�T:e�Z�Yѹ2pt���w9_.041X	j5��*��{by����9gע)ٻϬ[�u^��Ө(E�!>�Q��KW(Y���>��2n��.� >�J1��t��djG,��Ҷ�fB\��!=հ>o;pmkay#����ǲ�0S�s�yw=pv+��c�d�����3�8<mse�Q�i�cnS�F���v��+����uu�+F����󻋚�4gu��$w\3�g]�r�۬x���Gl����]����/5�"^zy�k�N��^�\�㶻ob��
s�Q���C�����n*�p��^�����gi��Ⱥ'�Z��N�\\��z�U�����G�ܬ<�mƸ�]q����{j�Q�yL ���<�Ʒ�{��y�F<�۷����tE���a���v3�' ����-��6x㹭��t{p=p�SúۄL�nώ���쇍�D9yu��:+>�\��F���cF����;���1��`��PfT�=���R�6.ģ;Xpr�v�ᚌ���E��H�=��ZݫY}!*�a봪:0�s��F�Ǹ%ϙx�!��63�Y=v�ۉ�W�cr��� ]�p�z�l�-@;md�:��R�'d��-z�y���l(��׬�l���hIC8��c)EkB-�Ď^��m����S��scA���y����x���۱���G`ǭ�M�͓:\��6z܅qeev�s�����]�m�87��[�c\Us��t��4]����n���눺��FC�@fĹ�����a�	�\�\����8�v��]ls�;��.����o��O=�]�-�9�βs��n,�Wl���Wcm�q3�h� �J��9�nlXq�+����,�#�|������ҍ��k�k�8�Q�K��&wm]�ۀ��JÇ���d��,iL;mk����N[F.���և�Mt�m�7*^��v��m��n�pc��R��q�C�ۮC
G�;�û{hS��5�8ۚ������ͻ���ۍv_M�����7������Iď-����xk`�ñ��o:���5�rܼ�j�7�۴��6t�ѓzC�/T��l���-m�z��gg��:u�sב�����^4q�';�n66'^���k&x^�l�콷G\�v���;a��58��crwݎg@�<</
�Q7��D4�� ��s��rq��
q���^�pr�N�6���R��9�^�*����n�F(�� �yü�O#��w�8 .y�խq�,�S�[h�c��].���\V����G���/E� P����ivh�c7v�R,�����[PJG�bdR� 
�i�F�9����t�*�g:�y%�Isy�]�t�^
ݞ�x�W&m������9�9�\.���!�;�Z�P��t��ӫ������hfg�s�63`�+�<@�˄xf=j���>�����hr۳�,x5Z���bx�Gg=�i'ů8(�O�.<1��7�֚���3����m�FD	�[�n�ޱYf��'��IU�ܩ�)Qk���J�tw�0M5Z�_W�/Ql �.��N�㆐�GǷ��R�ʼ0V��6>���Pf×�ݗT�{��p��L���d�t�;�)ޫ��V�-L׍k��1N?	�C��J#����[�������qIG�#�V��]�d{hms��enw���� �U�4�*4�3���xz��u��F"�U:{��+J���~����`�wg���h�����w'�Ӻ8e�Ws����9�]��-A-߻�HR>Tu�9����c���{ƕ�˾���U.���s��
��s6��5���������E�p�E�[wYg�T���|nτᩢ�Ю��n�&�u���zힱ�l&N�����e����7�*啻�����Ú�l��,V֩��/wĝ����^� {Wu�����7L�QxW�I��xWRɉP��q���ׁ����;C{ٞt���2IE�D��^����}�w��1���qyתzK������p��^*�)������v��]L�i�@r 6H[���9�W�W��MYO��I�t�'c�%b��M�g{�m�~��1<����z��F5w���&�w�T}D*g$���9�#�*��I�6S��i��dv�wƑwn#n�()�r��"���%��f嗅���G=��;�qK.��wѺX��c��d���U�z���)�n�(�j�f�](��q���ku��xϘ��K��O��z98���[;G2�BB�jP7�Y��4����}�i
�3�U4���N�c>���T�U�ض{G�0m����/rmAB������TV(� ��ܥ��,t�D����g'���m]��e��|����9M�x-�"tŷC+��/6v�vN�t1��R��!�Z ����Mޜ�Z��V�E���ށ}S��#�Y�v��/E`�R�N\fƽʸ�[)j���#�ҽR��M�6�/V�=.��D�������٭�H��9�q�����
ǯ�w2�熷���cd9���T�[�u/{�] kЈ=��b���(��ɢi�e:�������*�|���*m�=�x�l�!��'��(:�F�ovT��!��g��U��7���� 6�]v�	bH|6�/�M���&����w�Ԣ�I�'���ŗU��/Gӳ��1J!��u���ō��켥��J��	�)8��mb�o]��i���}$�PrO�j�4T�w��V�F�qe�|�,0u��`�s�ˡ)�uQ�M$�3�-�U����� ��0JU�z5i�h���q�瘓�ՠ��F�2�x���L���~��/I@��� P)��*�D?C�X�����jZ��U���V��/6��y>{ݬA��O�*|\�+q�\���F�,�������]ߛZEjV�#e��͗M�2����k���ɳlZ��w��kY����۠N3�x@nl�=�9p������DϬVLxQ`-�C�5���Ad�E&�y��?C��Jyc/�V_�~{W�G<\�J��}l���w�|�9W.����
<�Yמ�x��h�x��]��!l��]x�aٮ#�/^��w�u)�/�B��������;�Ƅ<�G/�d�^��C�V�"��z�
D��*T�LeAm5{>ʋ��d�2� !�[�<�V}���3����q�{E������Y�Hn�&*Ux�W�o�['n�X�y�������{��|6c]GB(̪n�[/k��s�ԛ=�z�u�۫�»��8Oe�)�t�����?;G%rMoy�߲r��w�����[}��8�d���V�RF�V���[������=U��@�yi���XhY��O���UCM÷���؃��Jܙ;��ɹ{�y�|D+w����^F����{={���3�����UA�ҫ�ׅ5E|C�7��w;����(�w�x�l�:�:�N��7��s�WL�`o�z�|��x�M�+ �[i����&��HV&촸��g�=����M��{9<���_Z����I��l�]������K���ro*^.`����.��[q5�\hs`P�.�O�����p�Is��x�&���o�G�8K�f_���3j�x�٦F$'���(�����ȉ
�5{h�uu�R[ȕ1�p6��VY�r,Rf��E��	�3oR�n������pJ�絥i��Y.vn��70*G�^����D��h�#����!'LQ�C�W\;�ɍȮ�r;�x6�8�څ�;ۓ��J�{w���*Bq��<�m���<zS$ny�tùn	�P:�s�hN��:5''b@3fz�u�۞G;����	p����٣`:n;1Ӈ�Ò^�����ɱcvu���^<s��e8��\*ds�d%1�g��s�F������/p�z���3h�#����ۏ�v�fǴ^f���zsd�sfz��w3�ѭ���u�趞Տ3H��i&�6?m[��Ɓy�����;��k%�}��<�i���ܷi��{��+���
�=��7^Sq��<nbl������%_�<�D$K�o8�o�����~ӯ�L�q�G��_~t!|i�y��<�7�%)��������;��j���3��&(I�i�˛�������Bf1A�N�e���TWP��4؃���]����T�KVx������b֖�����[[�);� ��R{2�ں�6��\�.Ƴ�
$G���o�oe����&p�y�&�
x����;����e3ՓV���V_��n�+~Z���pݾ���&�(�������9uv_5F��~y�\��T$��p�;]�i@yTΡ�w��s��괐l �`v�[n�;�^;lR�w�qlcE�����9N��^��KN�H�܅G�P=�*���\�ks�D��~�~�f1�}�1�%<46�~{��v��@��{�!6�9�f$m����򠤬��T(M���z1���_���lW(�GdV�a���D���:`��u�������D�n$�m'+l�O�g~��	�Ϋ�OA�g�^NE9^phmsɢ���ו��`�5������h*G��_a���a����yR�x^n�Wg�[r_n��"�HW#`��Q������	ҏ{�=rG�k��v���*��Y����t�u"LJ������=��Z��ne�?oeA�D�*9Gs}��Ղ��~Z2aB�V�-��;�h��*�c={����u��i����jn�������_����dբh%L��^�w�jw�k����c4߱̿.ӯ�+}��?[�Q��4\���}��/���O�u�E��g�������q�eT��QkR!��szN݄ݧ<vMέ�9vv��s�f^x�N���W�m�P�}��dW�ƭ_5"+<�'R�vqo,?$����"O`��+������̿�^� u�%��[�ֽ����D�)�{R��;r��g������ɹ�����Ł�AiB�=桲s��"�\����h�^�h���w������U�(*4 �H&��X\��R�N����ޒ�y�[��o��Űpz�8�k��E�&G&��`@��yZf:Ym���">i��h�>�)���w33�lKZ�=�N��%6��ثƺnP��S)b�x�ʳ���Yȷ�6���l+bm_� ܏|Y׻�h\��Q촜O���+m��թ~�J��
x3��i%������fa�ۯ_�
q�C �Ն��h�L�,��b�iB��ד�<�z�o�x�����u�_�H�1�����Ŭ�H�V�f?f
�a{<�t�!ܖ�>p/WS�5����ͣ�R1����gZF̼��|/���t��y\�ƭ͡ո��][��j�|�ٞx¼���Q_+yآ�]&�L�g�������/&[�}�6����{Ý���i���/Y
G6!A�<���xk��9��ϫ����;Q��E�Ռ�Gy�0���fgʥCC8��XX�K���sήҦ��z~��T�����~;���%������d�K�<7�vo`��4����t{�n�n��i��=�j)O�M�Ʃ � �6�P��6�hSlʑ5����}~1����8Z�OM�j�PwJ^{�:sj�u5��]��+�<���#�ؕ+��{�GwX��X
kl�ڊ�P�r�1�r�!�;@��:ȵv����<-=�O�-���gos���$�#�o;����Ĩ_���J��iQo�~@$[G��ҕKn>�~�dg,Z�?�uX}0}gJ)Ӯq�t�Y�z@��N�W�rz$=^�x=��#�e]
6 Dy����.�y����C8�n\Űv����[�:4.�u�LV�d���Y������<�i�<� ʍr|�;��<w����y��흑=�d��k����~��if�������rn�UD:�Ԕ��Y�*�6���yd� )r�}�7S	^v(�\���_d�HX#�?�>�;hל�{ӳ��^߻cH�i]
%PT!(_nN\���L㏜*7��eN�xԹy먺���.��C�+}uk}����� �����@�uu�;��''�W�\��8��A�C#{��qQ�w]��'�缝������vfn��;>|��+J�\u�[~qVP�z��M��Q����
^'�����~�^�>��-�H�1�X��v�<4��K�;
Tuv粉4����H	�3;��{�t]i�nn\A����0�����H��m^m �B���]��ĵ������y�U��5�.ӣ�����6���k6޻f.���mv��z's�Wf��d���w����6.�賝+�g��Ɍ�5��,�ȖmY� �e�p����$�(5d�G���pN�y�r���ӌ�m�̼�B��\N�W'F��W'a�q�#\s���@.4�Z�δ�ӻ���v�����zz'8��r�s�g�v..vX�R�x�z0j�u������&�͞s���]k�u�s��ur[�R3���]<���lmw�.��Pcd�&�����������Z�p��23���;��K6y%;i����#��\ʊQQ.���ݖ�͞�PtR^Eb@���Gr\�{^��>��3]n�K�~�8���F��-Mn%�uز��Ru����������s�G�'91j>�/Z(6���q�5�b!2�P��86����(�
���x��>���c������Z0�\�j�kŦs�{u��iem�����=�OE�z�nvWT�q��x(��씷o�n/7�׊�Z����_A�T�*���� �����s�v(��>�/���]׻u�J׃�j��0�nw����m�RΆ��4�=,3v�B��ڹ�v�B�*���՛�+k{rs�l���&�mdWy�V�I��a�]���ף��nv��wc�an'k-
3_�����1�2Ƕ�[{P�f/u���8{��Y�gm�z��HT���Ֆ�{����}��Ǿ����׹�H�ȫ��y�	�Ac��n�"J��C�F�R&(��{�O�8I�%�A6{�ne�J"���j��T��TWy�~���K]�oEֻI�6����-'fȺ��}65�P0J���|c�U���z�'��O{l�!�$�;�D/*b��좫��H"��bͤGt�xܽ��~#ɷ@����PU�����Q��%X���G���8f#
{�YW�[@@?o$��[z�>���:��gC��>ٌ�����f@��*����xJ()e�C���S�.�{��6����{���.����D6M2ټ��I�[�c}y�e����U�Ɩ��&��e�������Vq�ܵ�Y¼<��)Y��pW�g��ߝ�8����9y�[�^,�7h�*ٯs�&��Ewn�ɣ��;���q��0c�ߏ�oE�1`9v�ګ
:C<!=��=���9�Αq�a�=�pV��%��9;�g�v�h9ǽ�X�nqHT�ml���ն�Y5;Ѷ}�/Wu�Y�Ǧ���g��B\���#0�Gr�_;\M�u3�I=뱹�[�����ޮ�(�-b�T��U�TI 3���#��l��ㆴ��d���\w�W �}����w�w�����iE۵.m��:��^.�7���w[�>�;�E��;ktVX��e��f����v�}vŽR|0w���PǸ�I���^@ߑ�<���q4��
����r�|5u,mmГ�ҵnWR:�p�9i��ɕ6��[|=-S�r��:V.����5�R�8���\���Pj�S���NoP�mAb�@�h�R�V��N�+�o�!��^ÙNE�u"�o_׈eV�iSR�	,m06Nڻ����-Z�.��xE�;��9`����SNO	�m&�*���];�Y4� n't4��;�n���Je�eyyVAW/�,F��+}N	��e%\�V	�h;�{�,5�rj���&͝���^��c�r�#L�ۭ�χ]�:dXe]�9�m9t�@���G����̄�؞��/��w/�VHR��wM�7�r�L* ˬ�;zD����Ϋ��q7��3Q�n�۰���]b�,I��|���)A]95������ժ��zc�KΑ3�ڞ�I�Kݮ��e��I㇦��fv�����*�Q�2f���˸	%�����X���/}��`=�krV��ުݷ>���E8�uH�7p�x/z�g	��zS@[�\נ�������i��n�^wu��#�H���u�����6�_m�ĵs��!0I�Rk����x���A�;�鸜y}mѼ�S�mW#[��L��毻y�~��=��vxϒW��e��0�b�!�@a�Rgo���f:ģ�}�%��<����互��,���Fg��U���ގU��x���Y`�{s��J������jH׶I�|Ӂ5��K����{�Ӱ|�Wx��\�����ݏ-Z9}��{�n��{��Cuv��Þ�	�~��u]+�̐U����^��8f�,��pri�����l��s�-��&Q�ͩoxa����o��Z.Hb&V�#r��/}�5�g�-F�������N�U����m�O���|�M��?�oߠ�*r�y�ٹ���0��un�Y��Q�fx{HZi��o��ply�厈y�Ar:7�z��h��隕��#ο^k�z �,j!�rvjZB^^b�i�:b��W��G�*2�rs�\�s|�ǆ�R���5w�S��j��3�|�A4I��m�׊�n��z{��;�b���2Iy��nN]��o�eo[�bo�㽔N��;ze�hY�^t����A��h�
�a�Cx�{�&�E|.�yX<��٣=��Q>��I����3EYO
و��O�ک+�Z/MҜ�m5D*t�4i�ו�����8�zJ�ϛ>/V�������o�x'��
�g]�����:�����m H9�Q�v���4��\u�4&:��gk�]�<�y���S�u���l�����G@�t����6�DN��,W���`���4{���I��+;l�AP4�����U���{\��rt��P�͝^�:+�`� t�h���� 6��Gy8�wU����pS��o�v�c�� #3�=���M��p&�7)vCĺ�ފC;������P(W%E$��
gӵ���ˮ�]�����p[Nm�Ëܯ�\�I܃;������	@z�i��s��J��FU�\j{oM��(!���.��ܛ!���2��㘖Mr�ʉ2�p{�x�k۸Ǖ��4�a�g���D���y�Pd�_O��pXW߂p� ��f�V��_�2��.�s�q���hՒ{��O��'�;�V����y�U�!f\���zl���T��3X�VM��غ:�T"��U�Y��i�;�{���s���a]����qg_��(��ڻg>�=LK�hm�G>��ɰ��
�k���7�ڠ�5�M�|+�Y;瞻Waݴl�rF�^:�=�J�n����M�v�)Y@���3�u�e6���^�OmN�7\����ny�W��q��ے�9g�PԂ19x�e��=����8�nmǎ�x�������n�y3VI��f6�(�Y3��9�=dؙ���kqv�S;i�\vۭ�A�m\R�$��xݮ�j�s\�����a�8�ul���0\ф:�㰜��*�=�����:'m�$�qX�K�~?`f�.'?~"Z��r`5���,�Vu�_w��!O/�I���7.no41�:ķ�\����qw�V\+��9E��E�`�+����.S��V�����2�m�˝<��bm�����#i�^n�t��������_vxe�(�)S���	O�⠰�50��r�i䝚�w�g�fʘi�~���ګ����j����������~���b�?�]�r4Т��f���jfs��:(�n����n�wc��/ҕJ6���l�[�g�:G7�<���`_���Di`�� ���g��nJ�Sl���kb�P�:�v���ܪn� �^�/i��T�Dyڹ��2?�/�q��yy/G��������tª`�z�{H:�1�Si۫�;�c�ۛ�x�����m�6W��cm�Br�^�sY���7������$���#3N����ה�G��c�W@z��a���l��+���ݛ�t���Q'[����3���QTޞ��ٯS�v6x�tn�{�%`̩�S�^1ǃ���Z�Twr�l�6*�kEen�m��"�k��0o6�=��O��x֛�Y�f垞�ˢ����o���^Vn�D:�s��M{�;)�v�����5�L(�ɕ����*
)=iW�̘�վv.k����_���ן��G%���У�83��^��oV���w�2ƅ< T�g�];��]zM�S�D+cr�N�7��sU�~+(��S7���{D^~��w1�q�nV�����%3�R�رtw|]2�=���x=�IY��u��4$�h�m������q���4»�|jX�}�B����Lc��q�3�N�z�<�̅cc���^!<A,�2�����m���eiR�X9~�1��<bOE��a8���3n�<�g7\go`{m7&�.ծ΅�vw�m%��2�6O]�����Si����<1XA6ED��w�6�/O(w����c��^l�j뮦�2�`4��qs�����{润�qTV\s}��u>qȎ���&Fl�A�;f]�}�gh��Wf��>G�@H*�җW|<QV]��z̚����[�����[[��$���nGE�g)���>�	�*���X�\eÐ�휧)��3�f��J������C��7h)�{���Bbw^�s'�y�����G�Y^�c��(r�%I#V@)� 	�m��Q��][C<������?RJ��^dZR���cw����ݛP���憓Ò��r�/������Km�MEd����˭��gn���`ko+찥�T3��z���%���/:�ߕh�.fG�(:���a���j�$V�vlsv�	�d%�V$��Һ��[�v���ѽ�Y�4� �G�/�Q���=�~�J�.�J"Лwrݧ��j�����]�w�9HBs��u~!v�;���,tw_U�ծ�v�F9R�M;Kŵd�W \<4�.�	�Y��R�it�pC�rfv��
W���~$/�:�d�&fe��2��,`��tM6ﷺ�k��{p�!-���jw������=�e����T�O�w��?>�[�y��p�G-yo��0Sf�	Q���f�k��^�7�0�6���3���!�÷�#廠e��G���O���[�ߞ�Q,:Y�s�vOm�{��Qr���]Ɨ#2f;���Q�e,s6�Í�HS'����ܣ���C��d�@��ی��A0��PN� ���B�БWw�]���QHoڝ��{}���3��M�a�L�?7�����`�k����a��@ĕ_ZY\�D�}�]tv�[��n6��#<u�ydדG��͹z6��m���d��K%u�X+�>g|�G��ٲܥ���}�A���0䕷4Thp�?b>k\5��4��^��UAH�Fۅ.f�y���l+$o<��*v�� P�/˃W�i;[Gʹp��L�J�>^k\16O����Ma�;����=��On������^С�3�]�{�i6�p9��'��Ri��6s�ؑ��7�AY���3�I{�v�	�cmݼ�X�ˬ�b�b�*���"�l���?ߨvq�ܞR�I��=wi����9b�����\ys{|�Ǜ5�VX�b��`�o<��q��w9�c]Q�9�$�w���	ܭs��mc'+����k�T�K|C�=5��K�骏�4|A^l^m�0Q�遺X;���+Ӗq�o�'ƃ���9�t�l�o먋��9:\���ǘ���Ž��Ӧ����xHi�A?f2�dh;$���<5�v�-�vO����;U���v�Y�by�Kf��w:����۪���۳���mnyz�t�^nR�m�Im���R����z<m��N���W��ٕ��^�=�NĒ�Ʊub5:̮qm��Y)x�ܜ���Bq:+��7Syr�swW�:y��{�����<��pw]����k���0�ܹqmgp�7v;�p>�ast���&����X��x�T�פz@Q3ۃ�gg��a P5?WФ��h�5�_2˭g������YX}�7���W������B�4���A~��Z���T��*�{3u��T�L��3������낌��B��,�x�H&�A�e����&���f��;Yi�%bƀ�7��H�\@KSQ: f��H:s����t��(��o�%2��Ҝ\H^���5����5�oD�fOSK����RƻW*�ֺ�Ծ�H@�A������W�	�@E�=uv'@�=�;�����H�L�����:f�kz�,��d4�.�Oy�! X�6�ޟe��2��ř�ɷ����b�+)��1^f��R�::X��z	��sR�I�Bʼ�W]�[���H�䞬rk��v�S����kǌ���n�M�Wn:)��@ϷZ�fZ�_A�m�+7z�lI�rJ`�:Ͻ[k�/v�4߸k��j�wBשWyKn����<=�w]�A~q�0�e~�3���u���d=�y`���Sy��<�e��:G+��9e�I����\��7�����l頰Q��s���z�C*�
K�Ds6<*Y��,!^Lz	�:V
�*g޲��~��`h��s�{|�4m�]:��)4��n���}�د���BBfm����o$��9Y���ԝC�l^�N�����}�E{f�מAt@��x��M
$؊�Iezr���e�7��"נ�o�a�G=uY9��V�ޥ>4� ��qs<��N<�b�Ι$�Zn��O��]��R�!����V1\B��6z�dT�i��ޛ���_fY{���Y��T��Xy x&I4��}����x�c��up�N��%�m�Hr鬛n:��R��M���6FJf�\�\�i3��weP]�[\�g9}'�$W�E\�	�qf�I�]�%z�%��j;V�raT �CT�$�4Ale�KDm؛�����g�2ΚEr�k#��?'|ua�����,�Ƴ8�w<�#��{ՠ4�+�p�ܽ;�ƃh0Io�@��oh�
7A�v��N�9��L��/�t���$�'n=�Q�Ϭ�G���ڮŮ�j[��;����4�7�SH���".ﲵ��x9JUÝ7gT��Z��4�n	,tكPzw|G�әb��;�]�KM�ݯ�)ӭ�e�Xm1�G ��2���荻��v<�6�����d�j`Ͷ)�ݩ8y0o���3���D�mmUݵf�kcկiW���l���)v�s��i�=s����=,7��l�L�
�h�p(��|jϼ�;sw��v��)�-ٜ��ߤ;=����Ȭ�ҫF�Tt/�h0��nwO�˵�����G7V׃��nL�=�N2lÏ�#��9|��ᇽ���A]���=�ڱ�N����/j����ɛA����^��ܜN��0�;L�WS�FVX˰yI���!�\a�U����#C�wn|2E]�`���=�1�Vr�Ȅ�l=}�.���xff��7�wr�#�6U'M���2�d{xm*��~��[%�A7������]c����>^����&��~Ř��w�����*v>�H����v�8O-h�M�^��E�"��y���ѩhyo����B䙮SҳORlYG�}#��x��wy�����R�}��f�O����`��l6T��yao0uV�m�ו [6����9p�rxO����'P*��[W���`n�Y����3I�J|�� 	�d�K���z��yԻ���������~%i�C9�L]��3G6�M�/�m����ã���#��qԑ��v��p��bn��6����YF�eL�7e	�S��v��{>�C���&Q~��T��;ǡ�d�����_+�аfl�'�X��������AXӁ7;Μ8�����(��o2���wJCy2�����N�O(���ϓ%q^�}Ol��Šn<+��ʊ����Pt�TKl��\z�,����Ŵ���
�Ω��V�yJ��p�wUwn��<rt�Đ-zV ��u̌7�f��/�:c��A�Rl�uz�^���[��Ki�^��r���7�*��z�̺�����wݰ�g�*�ЮNs��_{�q��3��sjz��F9 ����R��ml=�1����n��6�B��St}�|P�P_�2��<�z�����j�쯪-Լ<�KW���r����p�&ܢ������"�g����Yͣ�u�� �L�Qaɫ"qbՅe�]җsO;D�òP���aIu;/(Ҝ6�(Wv��̜(���r�o��2V��Vƅ7Lc���VĬ;R�6%sUd�eVP�c�~��懬Ñ%l����lnԇĊ���/�a��y_�b*���5uCR9�f�=��.�j���.��(U+T�;��WhQJ�{e�Q.�c���g�V�2�Af��K|Za�'v6xZO���L��C�V��1����^�\�ntcw������9�<�!��)]�����d���Y�����놖B�߳,=�&0�ͳhm�ƻ� tec��,4�Y/�#��.+�9bC�]�k0��c\R�B�-�m�yr�-�rW����6^#��5���Z �#_W8������0�jM��7z��X�ms��� �;x%g��zW��zQ�E9s��/F�"���_�Ia���exؒ�I��B��5�s,,V�t-E��U�������S�e�L>Ad
�{۵�|SAV4��h����3��P�����Q�B���a��,���g�����bJ�͝�� �IC�{��@�fn���4M�X�4��K���k�55,m]����Sp���gv�/���T��U��z S�6B��V��N�n��a˚�C3�&��8ܽ�%��H9�Œ\�&�	;�ҷ���:�Q�/�jv�ANN2MKwkSnY�*�}d-��B��c����r��N��1&���x������h��۝�bus�v���[�i��A�-ֱ@`��\�g����j��iOa\Y��F�2<c�SC�1�{y�w�cW;���n9��=���g�.�);E��Q�m��-�OA�l�s��ي.wFs��|���v��&�M�n��k�"�n�t�̑��p�Ĥ3��x�j��<�1t���K��5�+O���/3s�9�`3ps�g��9y�㒷��l�nqh�"^w#j��������F�dm�q����s�ݞ����ݐ�;G�#�����;\�At���٢��-���uvמP	-��O6a�zw��=�6"`���ڮ��O�:�
܍���.��{�ڗpb���H'�]Wn�ujBԮ�
�]�x��݅���Nٳ�b��6�s1h}��uiKF۶�6+T����G^�q�=�ewg��cH=�95F��=���hf�n.�{p�n���n�����얳���T�M\Qnܾ6�fڷ70�v�ô�ct���8���˷Pnw=FnW��:܈��m]��l�V�{��ճ�v��t���}n�c�=@tk�.^�7\"�룎���:t�ƹ�Pp�۲��۵b�N��'�T�a�s�]u�&��t7Z�'����:Օ1���pWgs�)o'=��S�]��fNC��K�<��C�3�uۍ�謎�GU�5&�����I�#4E��{y����h��O6vz�벥�X��um�q����\��0�Cq��źOs�>�5ۓj�Nn.}=G����Gt���q�2���صgOW�YѤ�순�s�n��v$�q��{M1�]�ݙM��;�@���K��Y8ꋮ���>����2%ۍ^��A7U����u��9��Jov\v�܌>-r��v�&'�f���8�,��p6���rA�;�#v���gcN<\h:ų��(��S��^�p�L�d뵫��+���/]��Y��p1+�lc����16��Mf��p�Y�m1�v.n{d���L�嗧��ţ�C�Zy�sCn�\��0B�9H�� Ճu�<M�;jݸu,�����Sh緆O=����{�]��t]�U�]Ǘ/C�L�p��Y�����gs�Vϊ��#vD��)Q�T�����h�s�_��0;%��9�g'aۂe��\ka6��	��:����#����Es�f�n.݆1�;t�n�=�+�I�s�8^��<�ON�u��u��� ������i��;��)z�V�H�-:�+émj˘� ��mQg����g�YT��q� Q
TW[ ;����5|��>N:�d]���4ӳ��s�䥙y~y��D%H��p�ȶ�$�j���ͷɓvJ82�(���<����Ez�N��&�M�-K&�1�sm�O��q��|Vyz���$k켃}Zr�mRm�4M��egv6����Գ�f_����!���w�jhI��"y��(�:>۾�����HpGr���0�+K&�W E4I-
m3".��/�o.y�-�7.�;��� ��U�Z4�1��N�u�ŏY�a�c�vVc-H�@��f�Ps���
+{u#�v+�����}�`��E�Q��H����������bV��s�h�_�~y�2��K�㝈#���v��<�s�ƕ�-����)�Z������n��@T��� r��0�׳Z&�l|��o�9"\���cQ~{�n��]/�;]�����p�ީr��.��]ӑ�@�WQ�%����뼅R u_��F�-9����t:�'�q���67���rZ�<�Q��;w*��.{Y�u 7�Sb���aw���2G��})`{�H@)h���7�O�zMw��U���]�^T����꿇P-S �>%��>k8T�^�'w<�^�]�yVb��Z.��}Vc�<L��׵n�7���Z�����W�B| �,^�9x��R�l�;�q�ŭV����^;�>�g�u����A��c9Wp�;�1���S[h<�(�%"`��ǂ�����3(+�%�H:AP"ޑ���s���'G4G5��s���Lg�\��+�8
�A8RUA"��\�-�����|7{c��.h�w����{��{3^��/n>���:de�ec!�.)� �D�` �m�ᷩ��J���;}��T.#,�_�nt�B:׶s�[�C�M��'X�˽![ޣ	n0��1�wxkSrkS��=:IQGP1� ?W��̀LR�Ew������O3(��rxi��ayV����u1�D�r�:���6�r�Q�g>��o��.��;#��n��_,F0�����TN&'���75,���n֟Y��^�w����I�t�<�X��}��0��HS|�?���?-U��?5�ϩ�,����n�}���\�H�G{Tp<��w��hi�R�Z�c�ߵ΂��mS�.�0^VP����3zp/���os�w�+Dc�ɒS'�t݈��-�+���{��ѥmgR��*���%��^�.�]����T������e�jކ�쩭�i�$2m��u�#���{-m��x�u��h��W�6�@�ޏtR������n���~�ڝ[M����!7����;ޗW�s�� �zn���������
���|z����G&�y�pi�-zL���+ ��W����U�͎n#͒�g��Z� g1^Ly�V`�,�9Q�r�z�~�:�}}�t�黖6J�S[�Ek�,>Ii��m��	����qz�sϥ��A��ct�J���6��1]{�wSGn/���z���y���W�� �����]�gw[̃����L���[�׆��F5�\:����#m�Ŋb�/U�b=B���[�]bw!Ͳt��'EEt+]������1�Q_V�/b����;�s���d[ZZ�E�)eeqߜ(^���VΆǃഭq[%
���(�!��^�XF��^gw��T�yϣ���38��Yz^��g�Gt8�b
�,2Cc�������^�n���g����&�dSZ�ʵE%�u5la[�\����{'�x�;��9ݾ,���ճĞ��נ��.�f,�=�4so�w�̒y^�:8
�1��>�	 �
�Dh��>��k�d������(E�X*�@<��c5n��_��;�M�x/yo�OӨut�=*����.To���ܿ �D�3�{�m������M�e�1�d�������̵P�c�{Z��u�h�Y�7���tYK�ӓ2�ػ��b`��;�c�f�#��]���U���َ�د����u#}�.��uױk���u������*�r$���!��-���Y�X�L<Q�l�njI7�ǃ��Y�4
���C;���MƐ�V���La�^ e�JTۺ0)��P]��iL�
�p*^P��ʽ�ʀ�E�J�&w�//,ĩ�ȏ?��r�x�,�%Zz;�'ĝ����w�Z]VX����BK�CR���r�jչ��1��g�	���msv
�9Ŏ0���;)�Yў�v���r�6�^r�nN3���f9�l�Db%������7�h�Yݨ�7GI�a��5�����-D]v����pv�z9M�����|#��]�Y錉�nI�q)z����r�n:�۹8�U�i���v�y��y������mI���d������źM�]�qq�ۦ�$�������0S��n���FȆ����P��+m'?w����E�G��M�R��_��+�\��Z7�=��2WfV&�[�y?e�Wkm�v���Y�-._�ԧ���.o�|y�hI8{|#������������n1�ݜ�kݽp*�s�,������M�ޭ��rԾ>Tp�K����&���åh���gE�7M�A�3 _x[�2�v[�g���vs��˭��k��(k=��W����!����'x4%�`ёT;�S��U��Pޔ���)��(Ύ�GX�b�~��D����w�7`}J���i
~i(��c��H�"�wM�|Yӗ�+����[wy�P�U��ϯ��V&}�a�'��lc()$���^3�N�Z�5��ǉ����=���1��M��܍���3֣3�F�\��;��`7�v:n�����w����
T_u��^��Q��ӟo)k�
�{���3�]&��k��Cw��*S�N�z�t�@lJJ�޵���UN��L7��� ����b���F��hS��sr��n�)�p&�Y=�������\̫�]^aTϹyK(�L�z�Fo�z���׸Hs�����ӞJ��уn�V�\�����d�s]~�j�j���q�@�b�Jt��|��gd�5H��vE�-�vj�m�SϽ����5�;���R��e#́MR��Jf1l���^�,:��I2	������U�םݽ�R���j�Z~����onϓXk�	�\<{=���2#�ۻw;SC��s�Sww�]�q�-G�q�=�9�6De�)8�T�
�mɗ��?S\���B��u�A�o���G�#Ոy�	>���y�9:�]{~U^�8;>pQ�����E��쓞�pݸ�	��6ts��$�
��6��s�.^\���Hn��[p^R��ӔOzAnR�f���6��o��X���ϯ��`�U�7���!\p��x��.9�{�+�h�]s��h��>|m��J3_����o.`.��ߵ�V��ܓٻ��Od՜��jt�ɠ�*G�TE
G~G��Z� B���i�*��G+�}�<6ٲ���v��s3y�p�H�ʥOC�O�m�AF�/*4�������]��	��@IW����=3���G��}��oű�eะm�#�|��;"��{�Ju{(jߐ_:��%3/�v�Nn��̨X�7��m���{�^uw�b��j�,9��ex:8��m���XW�=t+���	Wk)��ꓕ
�d����M�u���v��wo���[�i^T5��	�A�~��߷�o� ��|��hr�ķ��1Se���6������;�߽����ۄ^F@;v��9��v���l[.��N�^{+��vU��e2�~������52�M�^V�g9�����j��ֺ���:�VV�HB�����"�͸���9�J'Ķ�� �oن��޻�w�y�S-ӿky��{���Z��x�h��;�fb�y�i���Y����~uq�.s�^照1y�署 v�[#v��ͦ�Z���Z��%��E����!����\�U�l��o��;��~}^*��U,N�/5��9�s��>-غ�;f�Y����}���&w�_'�5��#��Ӳ7c'�:O*�� ޷L#6߳B5�@d��gGJU����n�p
hM%<M<�`��e��|c���v9]�r�0� '����
Bʜ`�\d��%�����g�x��G{1_�Ln�1���M7G�Z �ה}��-H��V����S����vŊ��,�Er�߁��e����iv��{[�z����;t�˷vI�¹���?=���	��~�Kֵ��i��:{\ĽIq5���wO;����gWz�Q������zi��м=tŬ}�C}��`�)�P�|���7��]���z�����x$=�C�OzW�����K�#�1Q�V�++��yԾ�E^{�3���Y��U��j�䒰��p���θ��)~/#>��=kϟ�^���^2�s�{x�W/(��Sٹ�m��+K���h�=�#���H�H�����e�	�Uh�I��wce�EH�og��� ��=��}�N�$�(�t-��[���G֣��̙�|3��A��n�Y����Y^�s	bF+gE[^�7�{<S-�V�.>~�'S�:_���J{FT���'r����%>�-�{o�jM��
ά�yՕ�*s-a�V�al>�c�Y�t�fuBã�Zs�a���[��$�k��������n�����u΍��>Q�{�ˍ��y���C�:����m��]A˸�n�6�87+ۜ���n�����7hqp��׊y��ݝ<���jz�g�N�OA\�8��	�����u�è��ݫm�;�F�R's���Ø���0��D��7 �"�Qn�ػ1ƹW&n<�I�;7��;�l�㞓p���Y-+ųͮ�8��b��Fy�p��s�O6�"uغ���4��JI �T%{�3(��`����2�(��ܱp�/��H$�y��mt_M�H6��N�����j9�Y�C\���S��d$L(��K��m��Ҿ*�MnZ"�ZO���7(�=5�,�Z_��:��D#�2zC�z��x�.9�m��]�����E��h�2�'q�h^���k�����l�~��H�[��5����x淙F���Ku�;�d���M�^���WPeRK��K��u���k�їۂ�� -�w7��4W*��w�L�|;ˏ���j�QԩcP�}��z����m -m�J�z#&߳}�͹�}f�{L��S� �[�7�j��������H��lKx荒��i]n�I�WR�m:�ʭ�P��Ei�)�_Dތm����n���3۞�����֬�S[�0��i��M�CGZ�u�;�{j��S�߀�#�g�*���Y�Ju2)��(cTE�iPE:�-��=뼙O �w��8%n�Z��6��QS��V\df�����ɚ��@�8^Ռ��p���hSv��*��H{��l���9��	�󯃁�ʁs��6����w��a�%<z��g���;o���o��Q=���F��0��m��8f�3+��ܿ���O�����<����8=X��*�vY�Wu�~%��=�I�w�a���*$�lPE6/-���[}�#jN�Χ~�x���'U���9��b���&+��B�/<Qd���R�׽�w��<}�\�ו����X�-�'���:	��:��V�!a�B�	7���OkXȤl��ّ��H�s׮| ��6X�������9���
�;�L��jnn�{.���w�=�)ĒZN÷�gK{\�7i���\=h��nW��]]��24~�	��4�_sW�� �.��VN�E��t�w�^;O��Y:�>��W�s�_wy�譴�W���Y{P�߀M�۽A�B�}��O��Sw��ݫ�ѻ^9�:�O:�b�ݷ4a@p���2�y�VΝ=��4p�}�$W�]�i��﫩^雚&ei�����|mS6�N���&(μ^W��a�j��u߸�����w�/�V��c\��O��rnl�V��0u�$��=��)ixUt�� ��;��T�5nbɏ7��;�5st Q��]u�α4�Z��W6r$0�+��Y]���9��{��K�/��9#�� ���h��_�Q�D�+���
�u�n��|w�ke���I�x|p�Rj$���J�5Sh^�� �ɸ�W�0hz�}J�J��d�k�٫�ҧ�4��yZ+Lmf!7����_��
(�@�+_�0��#ۣZ��w��E�|����7z����{��,�*ig�If�4P�ѻ�t9)Q5��l��R�+9�7�'�6��r�K4,��P����ci%����g`���P���r�/bX%ɺ;��9+4C��2�n����޷D���ׇ�L�sF<��I�"Ǧ>�\;�oU��x��i}-��[�^Nj�C4����i�D]���,�kΨ�M��H�$�h�h�\�����Q<w(]B��*�!��z
ʶ!�^�I��뽨I}��2�F�d��(h����o�uf�kV7fs�|����6�M�X�T�9����S[U�m��T���-)�zT��Nc�[��)�W;
��io������d��%��ۚ(�tLu�|��[Y�j"�v ybo-�{2�Eک3��Y{l��>�3/���T3<qfG�8u'�#�����k�n�Й�t�:bç`�@Tw�%ڄ�%�Q�x��b:3��Ky�4Rǃ��C���{8s�{�pY��� ��V~�>X����7���q��v�7����Vr�^헣*�$-l���3��bz܏|��qʊn�~��U����{�^d��y�J��-�>��߅��/L_o�'eU��>�����mhX�9X�]�f�б��\��זxl�Z�
���DU{�6dU��o|&���}�N�S�����T�f7/��^���|���Ɩoz�c��e)Xꊌ�ϝ�(�x���֖#-�k�����ٹ��{m� G��`ESD����ƛL�^{Ϛ�6���2�f{�(ͫd�4��Z뺞_�ww�1�tIf7��ҥ��e (Q;ho��p��VX�����2Gޞ�R��5{�u�<v�@I��_�R+}�y�j��c3��[m环]�!/95�T��D�������s�U}���<��CF��>u������/M�{>��6d��#8%?X�x�*{K�k�nM���P+���X���Q��(�G�Z}l��ώo�Uw�+C�o^>��5'G���˒���׼-3~�����!.v�U�b�xz��e6j֋o»"7���v�/�R�+�<�w����9S��o�*�n�.�S����rb+���(�7`�u�[�D;�'�y�8�K���q�56"�݊�iu�ѿ�v����O���-.�UA�/%����ER)^�]��_OW�ԅ�f�t�y���i��!Wq}�F�s'g,�
66�D��]cy���G"/u����=Nu�.���n1�m�lW��uF��q�_N牝�k��&�Ъ�N�׳��^7c1h^�r>�U���k���U��٥�;Dm
��9�������0q�9[jk�m�>3:xH���d��,�ݖ�;=�X���
C}�f�')˒�,Q�]}�I���.�҅�;;=�X9#�$�	1@2��CU+?%t���9��X�㯐!3��7/L���a�S��C�����hwS�ƭw�Yh��gC>\;���;H_�i��_m���X�ZU���{&�l� �=����kHLxSتg�\����\`�ȗ}�����4��7��D���K>�b�@(�~���!�s �}�]��^���w�kJ�+�_>�*�uPD��u����y��c���V�%�h7��M��u��ߞ�h]�i�������F���D].N�W��.����U�y\.�j�.��/�ūܼ��������� ��\�V�ۭێ����c�M,�냐�K��
S�y���ݞ�r�ڲ���ֻ(�=��yY�5����OF�[�!�J^�	��lq9�46;vޫ�]�z��=���\h�a�.��O;����*�������τ���q�7�
��q6��`����N�5۝�ᶹ�g�ۛ��N�Q�i�uo\m�CӺ��T�%��s�c����L��l��[V�8��]�4`�mǃ����`���1�]��\Ĵ���El>a(?�^��[���5���q�K���WRw�-�^�#��t�G�=��}���J�rYAg�FWQ�|Zk�E[ˉ��u[�FnT���T��Lv��x�������C�)��W�&pxu�����#�>�|���Z��C/�	c�'��+��qo�{f-��ga![V��1���?���9�ڐ3�#מ���mF�U��.�Q�+���/��h��GϫV�Z��]�8��/
���W@�vuSkn�׏� ]�	.��&����(z¦���{x��E>|+v��U� ��z�yt�<���Myf��}Nn�^�s�O7W����)B�{[�:-]P�S��WW3�ý�����bý�26�|�.�ݾ��TU���ŐX�+z�xC�ܫ¸��7`�>�^���F<��K|U:�������}>$vx�禢�k���rt{c���2��;X�nqƎƭ<{Tv�!��u����`���a��K~���6�S;�%��N���X�l����ɹ��Ob����o���K��B�E4R,�M�~�vC��\�q�AIθ%{��Z�@p�liYK���}�42��cb2q�Gh'**����"�f$2�7�\�J^�up�c�L�2ЯjLr˓{fu����Ι����2n�{�GjD� :e�D����?�wU����C��UYD+`5b��������W W��Q���q9EX�{�t�r�>L�`۝�
����d]�u�l�.��1D�-6�	��ۀ|g�R]��QŎ����Ʒ��uy텊�Ωɑ��+�: ����=(VrΫ���X�a��t�)�z��ܛܶR�X*����rNg1��0�rCZ�	�f��}�v�u�"�r���lT�%���K���3g�.7����[�5'4�-���h��ݡ7�ݶ�H-���v���m���q���c����U�,J��_�z�.��_�;�n�{=�P����y�\k��x����Y�-��n�a@�e�RD��Kֶů���:B����Wu��p���F��+���V�⫖Ǣ�Tȩ�]w8��_k&�/�M���]{3owO�!T6��Ä��
&���k,S)Q���Y}����Ǯ�]�ݚ�޳'	ڽ��E+���n\�^��pQ�(� ���+�+a��<��^��{����j��^�򚂢�^la�9E��I�����o�Q��^�|�"�iF��rn��+�ӴK���ˬ����)�[��o��{�����yl^0��x�B9V��J��;���̗�Ʈ��\�� m�[WW'!��uE�{pJgCWf��!=�^۳���óM�IZ�r�Wzy���9��ѷ��Ӥ����z^־�*��,�v?���b�98�H������������n��x{^Zf[Q-��ݨ���<){}�����Žm��잲��]~����UX��nP��@�g�b��,S���8P`&Iem��{r�r7����3�mQ�^UD�f��W����^y|���9Q)��X�:�����ui0��v�߯e�Y�K�@ʹZ��!Qh����"kO��K����W�m|�7�쐻���#L5]��V��k�^���+�/�繋U��l�����k�JHQG���f�Q&Ac����rT�]��ԫ�B��.#[z�4�s��_\J�U <�`��тQ��h��>Ą��v3L�!H�E���r�J�r���4�nmZ��~c�-� ���.�`Ƣ}�ć�����N�#Z�Bg�4a%Lۼcv�]m쐏X��\�7f�z3Êwq�����;k�ģ|�ịW�[��2��{��?w�b*�Bd��ѕ�ΞMԲM��������s\vG�c����z�����6���P8����ox��wp�j�m�X���M4��<G��MY+���^���K��Н��=6f0��Yl��̑�i�(8���Wx�ы(�W"op����&������v�I�5�1N���w�KS��~E� ��x����~���4�F�C���ޛ�'[�����g�fzd~~Cf����7iH��G��3i���I�	0�$��z�!վ��S����;�^��!�?^7'Z�Ľ��Wz\e�'N�:��4?I�y~n��.�Z��]�v�Yib�[T�w;��M{M��á��r�#O���2tV�޴1�Mz��}��q��vS��L��z���yGZ
%����gt �]"k!��nS5u-��2ot���t�wIC�	�ww�A�1�Ġ[�J�]l��y��q��9aB&K]��ɿD#�{����G���fɟv��g�q�ru��tp�δ�`W���S�:Ƭ,����>8�\�5���y��#v�@f�ٺ�=u�슔u7)gn��}���k���_l=0q���zsn������v��hܾY�M��ǈyݶ�Υ7g�;�8���#�+���Ξ�ps�L�z���'�����ȧV�/Y���:q�n]Da+k��k�w�r۞ހӸ�S��+�������Rj�k7�~�B)�g�p`��gYyn��pg�yn:к�Y�y3�=�w؇�8���HR,��D"4l~��?~����f�Z�3B��Jⵛc�{q���j�}�}drV���Ľni��}R��-ew(�N��%a
�+-�z�oY�yq��-ױ�\�J�q�;~m#�|���M���A���H��+�K�8�	ne���YT�D$�d��_+���yQ(Zk�w��'�F3������}�G��a^���x<5�"����׆�����N�\sg��x�!H���[w�5��w|�3�U�_u]`��5R]��{��E�S�Gi���i�lE�^QN����l3]�\���{�]�qw/^ú��6�n8j�8v<�I6�;7nD<�y��$�ݺ8Z����g����oHxS��}�B��#�	���Ց��u�ar2`>�|�\���=�Zd
�E�A�ڽ�f.6<��<�pq�.�^�W۸n�P6k��":�E�Ф�N������a�Q帽�q�<����$}n�-:��\Rh���R� ա�ӭ)��]�ke��_\���[ƥ�y��>Ǡ1`�¢�h�|Տd���ָ��"�V�lo���;']�ߐ�]B�g��xw�Q���<m���TU=�կ<�`��k�$���3E�.n��*2�M�A%��f�2���wp;�&On+����^�Du�G��g��R�h�g���n�$ƪ:Ƒ���O��@F��5>
45R���3��˖"�w�pQ�n*�_�jt��~\��z_b�7u��L^1�W����v+y�uVY"n�2�Y[��3��-Q��Íp��p�؜Rp��n�Z�%��5M���������a��Ư��%��&	uepTF�Y\t�ǣ/r�z���L��O&�7�_�i�6�^�4n`�&O��z���uٺ����񮞝��:���3�h�=揝�S�i�'&�(� 4*�T&�,$ߏ��}�zr{���Kx���2�������挮��uޛ����m./��N����MOv.�60C˜��S��rj�/�!�Vi��j��v_`�I�ն��זѭ����E��.�%�(�W����I�%6� h4Ǫ��vd�^�����8w��>��@G�.h��u_��dZg���b �'���T�XZu��.�����U�꫊�|�6�@w3(TÍd�2�)N���^>����k� R�N�D��p��پ�DX6xm�Jr�^�]�[w}R�Vŏo����>خ��Wm.��U�-	�%n���^L�x+'\����Nؼ5O߿���o���{�t:���\}�Y�;���96���������x�"I�N=��h+��;D� �P��g:C]um]��*ç��HV��A�u�5/ϳUj�Ŭ�6��4wѕ�|(q�fu��|F��4P�Ao�H���l��e��%��T���,�������w�2��v)e�H��n{`|����a**� aڙ�&��C3�h�j�������[����mA�tn����R�g�ua�KV�/HD��]z��"���m�V�
d̲k,m���MY�u;{y]�X��uoc[���w�V�|��L��QQ��ҵ�B�^� r����H*�K`� �n`���asש[��P��d�8����z�'�u�a"���sw1���裎���|��WaeNp��,�;TR�kA6n{{2�К�����ۅ����3���s&i�4�+m�e����@����:��ޖ0��;�!Yj���M-��<�#+1�9�d�1a�I�%�����`��85m�m�؝��X���y}��Ĺ����Q��]��GYw��	Nf^"�&
0�e���"��i�y�[��b��%{m���<��V/nĵ��v��+�ޙ���r��4BAK���ogfr�l��{�\����A�9G���;,>�h��3Oo^�z+j\d)\��\��4���f�Ғ�j�KihR;`�Ӆo�k�M�*����U�oeE����;�,���T&�5k��5�� �@����� ���@$�$�$�$��	$	'� �@�����@$�$�� �@������$�$��IH�IH�I I7 $�$��II��$�$��II�@$�$��II��$�$��I I?��d�Mf8� �~�Ad����v@�������n�w� � 2�+�R�����]sấz{����Wx@k�U=k�U�y�n��D`t���he��U�T�:8�e-۔92-�uW'M��;0vuo�   ����04�00�����"T�z�H��40���1��=U�A �    ��T�Q�      z�%J��L�i�&&#a �DLM'�L��#i�z'����=}��Dl��{@DH�����P@\�X��e�2��i���TЀ؃��T(�Ā��O_�z>�,k�6=�� �{���^S��t�^/���@��	7���Q�G����T��٪��%A�$����ȑ�0�7�����9Z��yN��uu��w�x/
��7.��0U��l ^��r��|�W��2CW�%�o[s]��-h��G溙��*�Uǚ2 "r�H�����B�*L�K��h�r���� ���/u�pƨ�F
ĥ� v�T�.��s�z#m��hg�_b�*�gN�cIVJx���7,�s)	Wg5��i�d���z������xseu+9ۜ	t	��jt�B��Rߎ�0��i���k�D��� �+���D��f�I��G՗V���
*�Ed�'��ݡ*�f����s�Y��$=D�-���⋽=F�PHc$�$�����/�#&L�F�= �pr:����:�g><ήw���q��4P                                                  m4P               �                                                           �����wd����ݶ[$��ZHeI��
�"���n�r(�B9j�X�jĥ��	���Zv)ii`��cD��%���%���QF�R��Lu�84B5$�s@��*�:�R���KlN�+U�QXGQ���R�ґ�AQ�륵�ˉ
�8�A[��\�qH�M�#��f;[r���"��0�n��e����-$a��#������`�q�Z���Ed��QJK^i^R�v1�+�X������L�e�	�e��)S�[+��+�PqF����~s�k��؈��Bt�}`M�uk�.�{ 8��H( -+�Va.�D����ޕmw��           B� m�          v�ڹ,�i�90H�`Չ��8�A�F�0H�#�tv\X�]m$-
��vKlQ�cZoIcS��9��  [h 	n�۵vٴmV)�B���ʅ�����4������k�g�y�S��k0x�������nI6r�2�$U�o�w!�T�݋�I���<����H� �L�'�rB�r�k���ߣsxR�n|���I�����`r�U8�T#�*�U�}[� ���,� po�g=�gM(�\�R=��s�=�^�l��>y�    -'ͼT�ݙ�m��%(�����f���i�]΄�VKb��uJs�$� 3�tי����y1��}=
��iC=\q�>e��2I��<F3�p�� 3�]e��ws��Nʉ�ٍi#Ab�ã���ܓ�L�C�ʑO���IA)&�Ĝhӥ��JZ0�@�����R�]-�W�x�аh��ʭ�%B���;8�:���< �  ����X�T���$�#�\k��.�����Zē���d���-]�|+I��k/��i�>4��ٜ��Y`�6�%P-frRs6�3�\r���	P��x,i��M)��M��Kڕ��iW�Ĥ[��Lʉ"TKh`J�s&���>B��	�3>GE��kj�)���~��Y7��A��#z�Ú����Yb�f�e��]FR,�N��2���ff�Mv�"`�u�]�$gjso
ĤJI�u���+ӛ��N>�Z�f��fĹa1��Ko�e���Zr,\���BR%%���B��e��O\p������]n��    f]�Sb�#vZ�AV�,�3���1 �8B� � �� �@�J� �41<3�0 ҏA�*f �
�8s	��P��4-�Y����n�1ʦV$ڍm��P�1����ｩ{:�]��w~�)U��Q�K����JF��&������7��K2��Ӣ[�!*S.��]P��I<D��R���'��)X�u�>��D���۾JO�
�ElKMu�m�4��s|��N3P���	���&5�u�j�ϸ������a||��f��X���ߍI$"o�B,d��79�P�de	@�D�4��E�"�T1�#���@   %�R˥]T���S ���-�E��|	��.�R�@��d��t��%
D��jh��m��[��n,K��@��e̅e�3����Hs�F����W�}M8�%�k�xMF�|(O��@�7sU+bo�cO�vy��U�eדmF�'��nC�c�2�e%g����&m�tKo��ү��F�Ǣ�{��2Y!4�X��
F�-	�U��P� Ь{�3ӂn����ː�D	 Xv��`;Txm#Y�Z�j�Z��o-m�d�Ÿvixx\���2�<����'qX��Q	+��<���W��V��7�Lv犜��wj����)��S�� Y��I                        $��͗j���ڵr2�`ݛ���"Lq����\w��vTJV�i�	 �a#i�H�$��Uy�    �u�� Z�e�K
 ��ǅ9أ�a/E��8�%�sR�J��J7�J��bN|3�<0��bhJ��(�!7�m�,�62o���J�����(J��fPb!(Jy��q.��(�&��t����(w�%	JP�'M�dJ��8�i1	�JR�%	BP��8�����J^�JC6!(JC��J��M�hJh�bC�t�S�J��(H�o­W����d�V�c-a6��X(J�Pb �K�q)BQ�k�.{hJ����D%	Jo�	BR���I�\y�6��"w������p�y��t����)q8������nX�P�%	BP�%�Q�'�.XU���(�)J�瞚�=kFugFtl%	BP�.�2��7�	BP�%�9�K�J\N!)L��%	BP��BmÆ�%	JP�%)N丐�b��(q$�>YBR�%	BP�%	Hq��v��<G#֮6�sN{���X̜�$�r���Qxd�J�u.�S�HxZ�q����vfl�l�      �2��Z�I��r�� ��Ƹۍ%���L^��ĺZV@%�t⡕�p�&q�hq��-��� �))3�4��q�7�9��D�X��O��n	�l���{��~<!�:�� v�+x𛛛�d�ȡ�N5��*8X�]�7s�}[�<.���^�K-o�a{���"Vp� ;h+��z/ZӜ<�V�8,W�Pf7���S��\�ECyJC�����摍c���
:�^2���O>���Q$��m� `k���y���J�y��o
<.>y�yG=S��x       	-�}\��f�D�p�)���Q�'y�e��𵲨׭dT2}������F����<���@�6.4������3Th*�Y\��JE����J��7�o*�+� }̵�K����j��x%��[xZx�����H��Ͻ�2����4)�2r+���3�GM���w��<��}��oOZ���� ù� ecE�J�*J�RH� ���#�����6~�.k���˒����I ��b;���S3'�V:��3O��)�EK�I$�   %�wֽ]�M�%*������>t9�N �x�N�|eݯ
����R�B�ٚ�o�';�>�wѪ��睎^7���2��Ģe�2��������sF���׍��yq$� �/�����o�"�J7{|i� �{2$��vA�,�7�RTCL�����:�ta�{]�ݝo]羹����    ���ƥ��j����'@ɣpF�)�J��9D�1�<I6h�x|��{�=����f'"s���N��
�<՚���#}I"JA�wYbJ���G�_`���o&��2���W$�� ���P��kqj�	V;Տ����N��\I9xh���]��x�g}��e
�=��h�Y��U�;���O$��9�g4s���1���4���;8���]�}9�S��Ky                         )+f��e��*\��nݶI1����e�%خ�mP�NRJn��,� ;d���-�sd���W��:�    Y7kR�)b*Z� �+MS�ȯ���T�φ�422�N�p��wBO��H�H*�z�oM$9ۙBY�Dy�vqux�ĒNY&����!v;�,t����;��c��"'�\v�+lq$ *�>vV��,�cfsΥ�/��������$��M�?W}�\�b����m��2m�d�s��z��o     ����$ͳ4�m۶�U��e�}�½T��
�V7�3�ɵ{͜�.��Ĕ�Q�M��Wu��Q�6�6�U�^�2��t�[x4 8$��e�ŝc�;������cqffbU3��+jc�vw夤��&u�����oO_�ޓa���\*�$�%*	M�Wm�����2ϽG.$���f�J��=�����I��ν�   �][�6�Eɭۉ��
���S{�s1I��cP����]�C�|���w�^$�2շ,��;:��w6��Y=M]��'v*�x�$�!))
���kn:���&rWnQ����,@�8��'౑e_�ۚ(�Z�A^yp �
|�����g���s�%׆M�i"JI*,��|�3T\i�vn�c�{7{��]2g�kwԑ�9�sYq���+�Ыd�d��׾��;�|q�gsf�{�    &ډrk.�=%Ի`I$��m�"v0�e��v��d��]eϜ{�vi��E�}1Y�r^M����f��\�oj��7��I#�����N��I���u ��s0r�	hz�EAJ%EP�EH�[����E���ױh�]�s���^}x�$D����ƭl��t<���m����s���}����x���^@   ��6zdMM��d���b�ۑf�;�/�j�n��Xv�fO��W_R&���%(VȜ��]+�:���y���b�g�qy�{��#"����ewZ�零��J�@!���zI0%Լ�u;�ƍC}�0���n��1q� �������Gd���$`��N�{eBe`��-"l^�	�t&�g�JX.9�{�i�`o�٨�:�����Y �,��ޮ��	F���s�����o                         	��.�Y�ܛkw2Q�n֋Un���K-m��Y�,��wQ3J���5��1p���ɜ��    7m��u�ˑ�u�2�4F����U�t��fVe {�ڵ�Y�ԑ�����
1���mm;�!�mPf:�||qv�e�#D�Ԕ$��en���|��B��~�Gf	�Y��$�#!^jK{�*<gx��X���ob5I:�pݒ�<�dS��E�N3 �NM��29ZQѷ����]u��sp�7����@    ��Y��lM�*m,��J��I]�gl�b��hC��_ck �v���Brnf3��;�9J��뗇s��w�����Z�$T��MU��L�p+
�֭��2����x��l�o�����DJJ@99C�eݽ�JCN��b�ڋ�M�HH���@%E����a7wU�O>l;�=�~Oh�y�(���I$�   عg�G�ܹYQG
 �AB�Zm��Fכ���O���~�����^��d�XI���L�m�
�r����_0�.��ՙ���;ԑ�%D�b���S�ғ2�*4��|���h�E���<;�=�N�QT��p�Ι�*L��w�W� OX�ve��_�o���JI*	!��^�;4�I�YEr���a&w�ZH�
�+�'�u�oV�6�Nݓ�Y}9�1^s��g�f�}����    %ݺھ���!��ͷ�뛺5]�d�>�a(eAF׶(g�����䒔FJo�oa�:b\1�H*�a�������LM�VM�zF3n8C�����A�t9X��9�MQޭ˃v����f��.�V�੼���iӻ���#���$�"���c���Z6s�M3[�{��K/+I�@��b�ȒI$   -�[ajm�ѹeP
�	�o��$���s�ŻA*%��'��=�$fBS)ue����N�I�پQ��WS*���2�M�$�JR����=�9cLoWh��)5%��|n<�A�&������PJ�V-A	�ohc�t��]t����j/t$��^����2��|:!})�R���Pc�I'��*�e����g�Q��uE���S�ծ��Nzgy�I8��                        ,�Iwn�m��ݫ���&H���%*�mY �P�.$��bTN����Ys~q�    L7(�ʴ�����M:��V��O��sN�Num�\��{\�	BJNuۀ�@$����&��0��Vm���6:�F*TR��^wN�Z����zk>�Q���̼Տ��\��R �6N��\oif��
�᮸4�l,�ƥ?yq$f k )^I��S">��\;iu'��+{R���\I    7v�.�]FZ��K(��۰;��)�75rN��M�o��5b�뷄���"d�F�zWD�}b����\a��rיp;�8�P�~.w�I(JQ���bJ�UN��y�	��؄���"��&$�`�9~}�w������E�ӱFG�0��+ �Ě8h�9�����rdj���9��,�.қzRS���I$�I$� v��L�&J� RI(�Q�r���٘F(oKńpꨬ;(�F�湤��J%�@�)F>aK&�7$�f"m[����.��L��k��a�_b$ҹ}�P/*Y�^	��V�0�v�T6��`(n�H�`�Nl��WyP�1��ӜLX����I&�M�<3���k,c�9��_Ǫ�H ��V�'�4�,�6m��WvF��M�_Ń��og�N��gm�ow�    YY3Pd�*̾�E		 ao�^�ā����ѳ�=���
��I$ ,�L)��4�ּ�1�#ɍ[�"�9�yq$Q�^خ�=�݆��b��c�gH��I"�7��3H�SŰ�-��s��^��$w{a&��XN*R�,V5>ʛ�$�����-�̻<c$�   	&H��$n ��� [`6P��.-�k��U�	<��h|�p��t�F�cA��-��=�:�����H�����
)�'�$��f�@�6��I����e�w�;IH���$��G,�vr	����r�3^��-��hE�Z�D�I�y�1en����u�d�p�	$���m]sTPQUU -��
 ��{��ª y�?Pv@�M��9����`���n|��C�9����΍�օp����p��H�� ������q��>��	��`�1�g�oH0:����si3����h�����5�� �����s�h#��� �@�9
 /���#�������������=�A�"�J ��́��iI��0�v���\r����Q�?�t��:��$+x���A�j����oe���T �2��g" �|p"nWރm� z�f���k�y�j��:�6�ǡ�Ǳ����G���Y�@����k��T�����^��A�w�� ���>a����~`~�E���� �L����x	�?`M�?{��>�o7������ ^�h7�څ����= ����~����HH��@��;?q{ ĸ <_�0�n,�uT� �`Auu� ra���s�Ap)�� ﵶCB:�2��l3��<����x�����@� /��=J���u }?���?��x��� aT�;1��_�y(�G�9>�|� ܀y*���=" �;A���}�8�`�� �^a�[���,4�� a^�֩�^<6�*z��s�v�� � ���h�]Kc�z����)�� {��4�}��G���,  ��y���b��o_o! �@�A�c ��XC`u��'i�н�P��	Èm��ܑN$4V�  