BZh91AY&SY]g�_�f_�pp���2� ����b~ ���!��$�*]��A;4�/��JD��J ��R��J�)@J��P�B���@*�UR+u��hP�           @(     H   @               �  4   P ��=�흷�7}�;�f���w]}��r�w��]�:������݇� fI��g���ݮ��y���+�mxǑ(�l���Fx �o[�o]���(����cś�cФ�-6����Es� �ّEzx��:(�^;Sɢ��{b����[�;b��Oc� s{"(���Y�"�ũ���y/���(�̼�E({�AA*�E�    �   ̊(��z㢊<l�^{t>��=7֣�,�J${�  ��%
1�Vt�YfQN�tQ�e��s��+ף�27< �}H�͋Ϝ�D��^�%Q(T���K�4	W���QEz� �E�7,W��I^#Es��cF��
U}��/1�@Q�x x��(�j�d���h���ދ��^�gw[ɤQD�ހ%J�tȼ    t     x�QU%�s���R�{�|ϧg�:<M���X��]�Գw� ����]��ܼ_p}/��[|qv^`{ڻ�R��y�� }�l���.��7m�/,=C�D�*�&�S����s��ۥ[�cx ��J���7M6�t���:r�w<�ҵ�o< =ڭ��;��wnڞ{.��`<]�v������{���D�      ����K���v�+�����k��Ҟ�ݻy�
��� �t��m<^�ezz�(��Zg��X٫�� /ZR���ڐ��)v����Ku��{�/mwY�g�َ �����޼^�vힻ7N��t�r�we(cp ])�ݼ�k�F��${i[ϸ��G���{UIUPUO        �>����[^N�5�Ww�)�˶S�=��y�ֶ�z�� <Ҕ��W&��w��w�S�g��]�<OvҖ�;� q��(��JR唧�I"%T��m��u�l%����� s�ҵ�Ϲ�};��K�a�����>�vS>w/��{h�> �QJR�i����ϣ^}����2>���7�t�:  5<���i��F@��A����ъJ�@4  � ?��IUS@i�4�h'�T�4�T� ���@	�A5O&��OD�=!�G������ �U 	�   w������/ބid�=%m-�̚�3��6_$��7u�y$�\�(�JĄ�$�<Ą	$��@�$��i}DI'�)�@�$���`~�$ I$����I/Ȯ�W��^~��OW���y�l�7,A�P�3,Y�VZQ�0>Z�f�3��:޹f�d��b6���4��$q��$ѺKEW[�"��1B�Cf��R-��a�رtq��3���Q�5HD��>ƚ�D�P��e���*��s#�mWZ*�,�5]'�9)�\_+�*`�w�f���*VtWq��\��7���&�/��S=�(U$�n���v��ߎ���ƪ�.�nuܣ0u��ŵ�	XOh�2��v�b.�V��Ʒ����������U��	?UX��.�a��wQ����a�4;����D볒���r������k��<�g^ھk_[�h�F��s:SN�5g��y��~캼:�?�i̗*��(�ܧ��.�����$B�R��,����.�h%��G�����e�5�q��v�<vhm<o�-�.�Wn���v���~z�,�T�o^b����R�I�Z�(�b�4"��X�aV�3D�Y����K"�*�R�krS8͗@�Vfݒ��Y��%%z4�\�2M7���iː��?�<e�W�A�^� �E�m�4��'ނ��`��.��Z�X�qcr��蓉�4�66�����ZVGeMi�=y;Fa \�g�u�hr���z̲���n���[�w;��j ��D�726Gwb�ּ�x^�Z�B��`uƟWoU��z���,R�I��Ҷ����3WIfD�FjRT�%�nfoLJ��Q-�t���Q�9H��AՉ{WZ��Z�ͤ7P�4��fj��(�u1v�㥵��̼�.�~
�eI�5JLi��"�7�~�p�H����J�v�`{X��zrl�ּ/$�e;d��n���"�����Ą/;�?>x�(1���pՉ�V�:%���IE�cg�����]s0v�;V�[M�(9�����
�5J��x�
um]I#�����!�&��������O^nJ/b�����
�]�X����2]Zͷ�%7���R��]ީM������L7���Ӊ�,Mɢ��V�R�Q�}������m�뾇�S���w�!u�ܫx��6*{�L�V8p��%��,v���]�� �%Gn�����0T��)ڼ	e�XlS�L?8OZ��ft���N.���ٹ�2��8ÙEe��o��M�̖D�nl��l�x�-��,6��I�v3���7��{�3��2͐�eT�d3MJ�i���ݔ�k9��,[5�-bٔ[dM�2?Y��b���fY�j e��ܼy���+X���-MpUei-��lʅ��2�Y��H�S'���D�m�$ۨcO&�dQ�T���<�fq����Dvp��6R�
U&mZ�wGH�"�JZ���4	.��:��\�W#��9���Y�Stz�ͦ���E�u��j������tj-���W�t�V�J��q��V�s<�֎=�Ykx��Z<�"� ��t&�if�l���6�
�3l��s���W�Z��S�QAq՜�5^�����~r9�������������q�׷΅G(���F,YSD�37\�qRE�Vr���?h������[��k+�5�DME�u�]�B�fe~�?_mK�h�eA�s�EMU4�p���XH���)fDH�`���2m^涂��8~5
���GWL�OmU��D�:��-��7�]v�_Wje��*o�/3����*�Mǐi�/m�L��v[c�wg�ʘ���+c	�,
��Gl-�Ȫ�a3��Z���Z<�x�����Գ5ݫ���������/o�K14TY��NA���XV�P2AdC�hY�.Ŷ�D�M�q�O6�&t���P��hR$�N�)���`��L���t����Ή��q	>�*p��TB���@Κ�����Ś�s*�=�i3�!�i�X�Jץi�T#&K�����;g.x�9�ֺ:(;���� U֎��3v\; *�{yj��5m�i��Ebк��6�7��(��3�1SqOR�:])U��w3�a۲�]�Y�:M=Ƭ�T���9����ݦG��)Q�����9�>1�ܽ��D�b�+��� ��o�C#�"Y��ABV��^�$Ǹ�̺W��Rd���Z�]��]B2�ցq��L��&e�\��8-n�R
W��%p��'K�j.ѢQ8��Ϫ��t5���sR[�Nj�R���w�иS��^ei�1�٫���A�w�H�t����(s��I���gM��C�i4��s��q��hmf�;�t�]Y�U�쮣�^�ʘB����E�m?<Җ�.Ɋ�*v���	��:�d�z뺃��R�-C����I���2>��It��MB�u�U����i�x
�Z���Vu�3�Ʌ��W�w�#v���3U"_M
\wI��'��Z�������č6�,���╌�R'�콅���Y����\iS��Z� G�ylEd���pu��WC�p�%����o&�hR��pM��W�⵰��scY��^ey��7�Mݬx�9yab���H��sy��Om1}ثgZ��kI�Rt�Y�1;�j+,���.\���P�Ÿ��զ�w�So��:�E\�t���K���ĸ����K�8Du]G�T�xk�4y�ro�؍�k�ć�B�s�t�1Q�V�5�[J���i�o@u2��%=�&ST�d��$��cx+ n���P7UX8��m��%L3�c�7
 � d�ԂY��l��yA;ڏm�]u(��c]��F~ٗ@ʠf��R���Nh����s�sOg"���������\�l�p���^Yr*t��ͦ�0K�ڙ�SoV"��+^b��4�`6;��px;�JIoK��靶%oY�WFu�*�±�jen5()��t�L��m�2̵����ev�\�jk��Z�~�{AX� ���yxoV ���Rc��`m�(��MB$��N�������m;v��R\W��BF��
X�W�)Y����w�=�*��Z"Ѹ�rn�"��Wt@s;Ql����J�*�-��k��F��,���6��7����d�ޗ��^ԫ�J��ն�:��/��,�8��q U{Ws/,C)a�ض�+���V�K=����זX��pU�%��K�sf�f �`�3j�Fٽ��	���6�ˈp�c�wF�X����c 7�q�P�<�`ؙ�u��o�7	G\c%&�B
��V��WCx�Z�̑���%)U_�D�.����X/s񳜶w�4n��	�I5k����^fpᕤ���\�3u��~���hT�U&Tz7 ���j���Y�$���ǭ�ρ�.b�����Z�0ѫ�l��[
��k��M<�y/�X쌙(5b����+���,����	�L����5���b=�3�V~qeJ�\�q�ȏ� P�5�f4^���]����,��m����+*v���ʚv�7�/��RH��'k*����e�X�[��/�O�o�r�re�f��F��W��r�'dÍ�	�-�8��Mي�����Qf���U@#k:)ۻڔ���W^/s~�a�a��-��I��4;�D*8���t�	�\0� ���-��o�f��b��+��4��-]д�r"0n�x��;��W`��g�7�L�t��h%ǻ��v�g�8:��M�L��Y�8����v�:��k�fG�٬{	�p!�P(ݨ9�e�H�t:�%���({#;d뷮����D�s6��_����T��^aY6n�\˚ƙ=��	q/*ލ�q�:첢C�DWav$hp7�qj%N���֡�-Z{�����]�7UȪ�̨��
�7E��ܖ�b�v��Jq��XɬS�Ics	P�Sɰ �v^��� ���� �ŏ6��xX�ӔAU$�r�e�r&=nZYQ��S+4^(��[b�W[,�kh@�z^ v�{2��0Rl%&"�(K����B"����&I�Sv�K.��� �!�n��4���h��+V��Õʗ]ti�52��p�ə2,�y�+K̧�.�D��cU.1J��+�$�)s��@��]��塎P�&���3@씮��Y�-˰5�+Ѩ%$@�HlG���G���:k�Q��5i�Wj�Z�I`Ҵ�eӄT�H�m�rC��Ich�3�
������z��e�8VS�	U�ǳ}.��7�1��'j����X��Ir� ���yQ���0���	}w}Mau�{C��8�z�su��6Ri�N�+�V�	�<&�B�r�#�X9��:�"y��7SD��Lr++/���#Xwv�mL��[i�y�f
��7��Lmd�O.��G�N
�]^*�V�8����;�Z2�E���\���vg�U���:	��h�Q8�r�n���p�s+MF%8-3��t�4�I�e�U�ē(�Sh�*��/r����s��
Q�Xx�+�sB���4ʔ�7Z{a~�Ol�a�%�u2	F��Wu��G)�c� Z�H���^�65^���e�T`�M*͖�ԬQ��ڡ�E����H��s5
4	-]��L`��i ���F�ʓh/q7�"n�Kkj+�M�wW6�@*�n�䴳?,��U��V:yݲ��u�+�vv偪]ҋuU�����
���jѢ�"[CN��;O"��M��R��yj�8�td�i$o� E+�Ց��xL�[ I�g�QEr��t�K��\]�ɬԬd��uf�bdѥso�^9��V���f�%搕B�	Ձ����0ݔp�e���U"�i��+0Si��Ha���x���QV�3@�mn���U��"�GwM-�3]]dʻ8/�Uu.\%d��w��ښ5�v3+*��pG����l�Ml6��q;���J��r�8v�N�o[=�-�T�����ٷ{�M0IɩY��U�t�\�̸*V�*� ��,J��Ƿ-n�dr�
"a�wZ"�!a��2V�K����!����Ųr���<Ibv^��?s�{tx�o)�m?Ƙ���i[��rQ��=��m�pP@*ۭ��e�������ݳ���錰3)���ft��
f�,,Z����Z���~աuj�����WjJ�ZIo�Y)����3�P�(�2��t���`�%���}Y���;z���gP�T:�R�7��qK�.=���M�Wp�6����ݭ��?j�V�B��:-���`u��U�yi�x�(a�n�eS�g��U�ġ')�'s�1�9��A]�ѕ*ؕ[��̴t*|�M� 	Mz]t��?��&"0�H����=�`O�Wߘ�ݎ��T;v��0�S��F�ɽIɋkz :�P�R���%u����N�]�Ay����.�n~f-
e��U9W���G̲�`rЇ���W���k
���Pތ�1�W`���.;B�4�1
�cj�,�a�:)1x"ɺ�f��j䳦�\��R�3&z(��CwqaT��i�-J�$�.9��T��3�ݩ��9��ZU��A��D��H�C-V�b�@GN�ˡ�[#Vޚ�U`L�&G�n6Xn��4�Y�;���-�~h����[ŵ\J$VԵ%:[�ֲ���a F"7{e�w�[�XԸv��c5�Ԭ$�髐8�� �1�m�;��뵩�
�̬�����m�*ԧ�V�+�G���w�Yd��0�����[!���#N�+5�,�,:$�P��X����,R���!B�;V�~XV��v�d[Ov�4�Q�S0��d�6��R�];��  D�R�x�k�y�ۛZ��?���Xe�{��Qb�*n/��^��;wcv-��U�����+fm͚�11Gy�=�]g.j���kE$�!��w��0�R̙h\�)q�ԋVF�����h	mS�w[e\�8���Vf:Ք�5�����&�ŝxj{��$8�9&��,׊lT����"�i���L6������5}�Ԩ��h�U�R��a�[t�b��0��$�Vi؊��$I���&�on�xp���!�;#����m�됍��x�ؗ���'� �(wp�c�wj¥j���e�+���nۄ�.��l���oC	l�薨�̨�ymml�.��증�/+&�)�k&�U�Mؔ)i7[(R���j9#�2���㗉5b�͇wohr��v��w_Q$e���k��ʬ�����Q1<P�9b��6h%���um<�E�'AH�'�]�o/+B�e�5�a��U�1�k#5%eb�x��x�gl�,�����(
C#�h���+ӫgu�0�P�{npd��mSKy�u1���߃�(�43�d$�������3��ܮ�/:�$z��*owj����dU)|�x]Up�LK:eeV��S|�x�=��i�`��?b��Yʱl Wn����
�;�_�2�:�9&#�)]l%O����M�;�Y��>�~XPA�xVfuѧ�	���P`�Dm)@6M�����Β����uԩp��7mWwm"�9�9V���S%!Uwi�M�1%���J.���H���u�ykH���:���E�0�)��&�Yw��7,�h[�����@hۋ��6��H4��z��X�]��!Q|�/��D��Y7�I�tܢB�P�ӈ TI
�!x#�L0����9Yf%j؈�),4��yݚia��@��jK� � �>i�Z��G�B���:��\�*�R�p��������;WA����we�O��h��1kB�����۩�B�t�%bҨ��i�)���l��C�
�� �Ka�Q�b�&:�QN�A��q��.��FbL��`�KE���n�8��Z�h�Kbu�.2n��^=���~bmn�`�������P��W墪MN�p��������Ʃ�I��!8�<��5���U;�d����Oߤ����z�����ķ�Pvl��3l�v'.��q$-�9WN$�R̨2��3u�heffXj+9�1�x�+]1��n�#e�&�%���յ�[��Gqk�ZEV�~��
�mU��i@nd�ãk6�n�Wu���L����;��L=ݼޕ���ߟew���Mܻ�?�x���������$��I$��UT�[UUUJKW6����	����認J�UUUUN�����R�P�@U]T�UT���&�-���5���*�mWT�U[WUUPS�ST���e���ԫ,R�uTQU���j��(�-�R�UUV
ive�@����R�UR��`6�),�S�V�j�V�OJ�;rEI�ɳ�l@5����sV5<�\��A����q�}W*�URQ��W�Z(��
��W@֦{�U��M��ę�sUWUʰ�sʁU\�5U5�J��T�3ti6C�����WD�UA�6��ER�P��4�(��)�j��j�����V�VꭺU�Z��������h)j��
���U���&��U��V����T�R�+*��趪�Z�Z���4�UUUU�UUU@UHI�n۠{d�/c��l���۴����۞K��=���/3�Kgg��p��VNv3���������$�@:^��\�1	�ls�jV��듀ێ��g�:�j�����v^�.���w��f骞�i��m�]e��s�vL�O>��ò�.��qa���ۥ<���Sخ�����i+���i�{h�S���ʛq7��h���9dM��]��=��ۧ*kv��wZ�C����nj.�Sm�l�ۦv��P��۫��~W��7۶�n�s70n�m�1k�B�޹�붭WX{x�/-�ێ��hv��73a׺;�l�l�.�9�xz��Ύ=�5�V����F	3:y#�e�T���Gܖ�-ץ��z����<	�8����:�|u��}۴����̖#�o���Ȝa朚��n鱙�.�m�tx�V�:�Oog@�_DD�،L%�v_7�8�f�0�z�y�ێ�����ΨB���)����nÎ�pP�^�S����
{�N4m��=<�{Y�Ps9{6�
�Į�t��jp��\�]�ks��2S�mXٷS�N�Y���t�m�j�����[bz�Gc.Nݱ\������؎��	�ӄ���k]Z�4�tu�ўۭۦ��gN<qឱ�!���gcr�{<['[xE��x.Q��g=D��w��żY��E��-������źY7 F���WG3<���G�n �"��(<�k�$�盟Oe�t=��5�n�'LY�>y�ݹ����,c���*��n%��s\����V��H��s�NGAm����E�vl��`"����^�Օ8�;l�;_/���wkλ��l��6��HGmɝ/&�q�K˫��=�Q86ݺ�T��Ɏ��8�r9��>`k��c�-�v�2%��:.��v�4�8x���G��o#l��M��n�v�c�!�F��[���l�[�%������s���m���/@.ֺ1۫��)�ml��v�>�Cr�~�n�N�B��5rvQv��^����U�6��H<byn׈��+��1��H�mX�3ƙ<���ǎ��$'\6��&���j����.Ƈ��� f㫝�A��l=Qkv��P�:�$UZ�?X�1%T+�b]�9#u\��cj�ky�F�dU����9�ۥ�W�	VG�%��89��Oq�ݴ󸙌w9���O���.ۖ������¥�G(��S۶�v%2t�[c��A�ɛ�xrvV�x*�q]f6GV�W��A�P��
��pP#EP�2�$�+:���\�խ�&��q��u�9m�;	�m;���{E�֮NS��f�e�y��i��v����c�{O�nV��=mr;c7���ع�M;K��.���D\[���N�i�_lv��0W���ܾ2<5�K��s�����@Yg��ל����ۙ���M�y�s����m�؏ [�f�\�'��\s���]�v����!�km�u�Ϟ�}i��Ѯ�ΐ�O�帮�N2��<�r�q�5���kzY]э/��ˣswG�1Sn��@9��:�:3[���!�]���KOj�t���׭�n�h�7��#��,g]����'1�+x-���S��T�[��=����r�ʱ����>��+�okl*#&s<	��h�u:��Y=���X�)I��{YF��ywoJ��=]�zt�m�᷵V�j�Ƀ��[�2�wl�Z�l�vZ�;o;��ø;^�Gf�mb��㳭\WOFA6NړWn���msG.�F�Ÿ,Vƃٻ� v���3��MΟlk��8�m:��X���qe웭��q�9���S�S��;��o���s��1��װ�pnw���wa*���u�n�c���y���ح�.�}�����,�kzBt;V;a!��t��7nFP{��k��t�u�N��O=�8ܨ�ܽ\v6랯N�˪S�s�;��
vYx�k9�#��9�#�9�x�Ŵ��\�5�eݷ9V�;�ӕ$T1�� �-�"4�"�5�!@-M���%th���㱙N����v�v���zjmu<��Vͱ .�9;-�T'a���i�n2vm���vn{%��+;�:A����r��F}�h���v�E����wŵ6�r8S�/jrަNH�ۑ˫��ٹ��ݕǲ�۔��n�u�p�B�=�v�¼�2��
��m�nH��7�V��:�nNH�8}��ш�ۅ�<ܶN�]����#� Rw>�K��睚ocù��	���-��������M�6α�ʏk�A�۫��mqs n�97WWI��;n]�=�nTD�k�U�힭�q��c����|�x�����yt�:i���lc�:-nWp^�N��N�#t�Ƨ�;�����N0L5gggm���9N�Bt�s�y�,dq��NKn6�`ŋ@��ٻ]V�d�)2�-t���m��q�(�k�s��u�	���yݱ:۷����M��:����y�6�nڻh5]n:w ��R��F{�����y��<�U��62�n�ˆ:ݪ�u�4:RI�-��:����m{-�Ss�f�/v���uq�2�g��zKsWkj�Y⽇<ZQ�	�
�',�(�ڈD�W���i�2��N��{Q�;�)i㇠P�uv�غ3�^5��x<B[�t6�s��<�u��/o+�Şw�g� ӯRg�}}n�Cr�~���=v<� ���J�k�rU�R�{u��|����.�q��'5c=�Ŷv�Y�NwSc��m�om���l��������7>��ͣ31�h�<W���"���pd^��F����b͛��+�o	m���{����
�L�ݧ�5��d����ۊ�ͳЇ/f�pd��g�ݠ�$y�N˹��=�=��ѵ��kq;���6�_`Ajrvm���|�=�q�8�gp�'U��Ysw]���A9�Ɇwdv��-��В�ohv�p�e2���B���k6q�=zH���pbq4��&j�n:�n��m烷I����L�O]���z��s/$�gۑ�0mӱ���"��=�뱵����C۸�x��ש�pvܝ��X  ��h�]=f�O��b�j�<N]��3{-+�R�f3��>��p��e�����Au��1�K�4S�nۃs�J���t޴����Vh��<- ���,��ԅ��a��"&m�u�(F��6Ʒ;+�6Π�>o\n�T|���=Cq��"�ش/�����v��h�U��\�s���mö�mu��J�m��m��|��byܫ\ne6M�d�^�
��l,{pS�a�]���x�f��2��Mν��y�:㎺wh̺nG\�s��#��+;+����\��NT�a�{v]�֕��=������l�����]�6q`A�Cp�����qu�WZ؀�=o69oU<kW*n
z×3a.�t=u��F�v��o�v�3q<�c4+��X��{l[���v�d�b��q���[���5�-��t�$�Ǝٯ>��S\�Ϭ�Ïn�78�wf��+�b����`����c�q��o�'�ppv��g��Cvn�
�X&5ѷs��<�Z5��m��ғuHsܯ'/n^�������8㫶�N��[m�$�6�m�a�1���YN����֐�۲y��m��^���ZԘ�н�G��$nR���A<v�s�n�^B�H�L�i�y��Wo=8lb6�]��ې��t����;̚;�xֱ���7Ӯ���=�7&�tǭ������˵-�]�N6͇�m��+���:ڏ.��c��v�st��;�Zi㵣�t=1:3ۗ�K��z��5���6�ʇ;v9���K.�����;'ۃ.�#�cM�t��sĮ�l�96H���2�xG�����\q����o:�;F���ת�y@�ۮ��G�6��s��M7q��y�i�q]���[n�HGl��^t膜���	ۮ|#�m�Q�nlk�]�7�,��/v91��)��ob����c�8��h���܁������g��a�:�L���[���}BѸ��g�qϞg����a��*����u�O21��vMwn3�]�t��uv�s��M�Ʋ�ncj��V��v�v��u5��s^U1\��؟n`��۵sۖ�V��ݣ�.��u�n:���ub����=#����k�C�LSr�l�cF֬9��U��V��/\��9Ş���^��3c�{$-{��8ot]���n��,W���=�����1�<���O�N��j�5�SͶ�<^vh����s���s������ ��۝�ˍ��ٶC��yR9��cN�ī󓋡�l��m��4������6��q�;\��n�7s�\v��ͼ�z}�V:ⰨhLK��q���n�����B��0�3�s���7Uݮ��1\[-����n��]���f��U2m�s6�����υ紉i츼&k�9,7�qy7<���պd�F<�q]���0^��GW<��O!Ly�RW��p�x�Ѯ�p�����F�:���l������KrpXt[��8E����{��^�y�k�lyűۍ(����\�kv���ɰwG#.��;@�͎�ӳ�un�OHtr��4�l�����V�c87�&���7�s�ݞ�7N۷�O��k�Ϟ�s���u��}F{�9Y�k&�@��G�Ɯ�yub�:ˀ���xsz�W�/g^.�<$twSӝh�;'=����/p;7�;ٗ��M=�v�ڷi �@?�z}�.��r�]��3mmț�7h݇�^�E"��8��m{<5՗L즢�܎�BԹ$*�T�;�$�]�x��$�St���; I�! ��� $�]���?7��B��$�����U*���jjU@k=�"���
X�M���V�-U��@q-������l"C8y�L�$��e�qc�UUTmD���T,��j�4��8�����㛫fѮv.fI�1ێ�ѻ��3��]A���Z����,<��weq:7\v~����{���y��]{m�qU�5�5ٝ�џ[��W\rE�����ʙ��dwX#o<F�v뷐��v[�$�6.�nn�&�ѳ�Bzo;v�6���c=]&��6�unN�i�xS�������1�m��L��7\uT�cm�c�����vK�@�VL�GLr�f�l�=�뮣��ힸ�:�����Փ�)��5���z����n^�b��ǰ�Z�zҖ���N��6�x������➴�L���H7��Sqʎ*��Z�
2"�!��P��n�u�+gz�s�׌��\3S�wd���ism]\q��,�	�zG:�Mt�O�J�z���-�V����[ѹ���pV�[�D�v�����{g��d�L��=x��L�q؞����	���հv��9�1�������6)QMύׅ\=<=�3�/v@%�P���ӟn1�h��7g�-�ε��`��lI&�e�nQ����&���g�m���-�x�e.��\T���Fs1��k���won݇M����d�^�sݺ;�[3��XMHmlu�lm^�����Y�ֵ�J5�]�����rf^9�{x,n4�=��ո^������Ξ{79��l�/��㴽:7���.N�y�]g<ٳj�ק��;]nĻP㭞�����.1�L�mQ�}.*��u��f�Zy�+�z�mN�>:
��l�����G!l7a-��C�6*��LR��K+��AP��VA�n÷�0x�sXy���G����q�p@ݶ�;q�s��g��N�:����;���K�v7g��^V�ѷOF�x��;6C$]�΀�h��\�.�I�d_Y	���\hX�]6�l�n�:��Txᒋ�d�R9
r�� @!*H^E�߅Z6[�d���m�C�Ռ���t�����fI�t�ӛc=��[H���Lku֧��N�J3ܜe�v��z���[<��yRݛk\�{+C��pW���؋��8��q.%��Ȓn�0��=\�]���vw��r�l7[O�{�t���i8.��q��D�lq���N�Nz�����e�wj�8N���s�x.��������p(;xq�M����wS��s�=��YI�e;N��t]+��z��xe|�>s ��[�}7�"���qsHC��ĈH���Qc`�R���P5��\�u�ޢ�2ū�\�tʹ)ݔ�r�T�z�9�#6�TTZm�p��t�թ@��t=�;*&7r$<�]Eƻc�9��u����Y����i1���+Cq�+	)�0-,�+�\��b���EAu���~G�%����'��Bdo�/�6ѤS�1)6ki@�}K[k���Z��zWL��T��ܩwf�1j[u��y�V
K���*��S�zTF�P{a��
��ػ00�xh-hC\�-�ݛI��G�>�Yceg�P���MXƤ�:�"[L�B2n.'���n����yTuw��f5]�0eR��6U���f���ϐQR����aOtp]���{���fbCH�p�kc�iE�R�: ����V�v���B�'%��'.;%nc����=ut�*�փ�ei��gv�̏[�	F��3��&��x?�t!��~��MV�l��Y�e�WZ�C=K�*���
�D*�J��DR�~�nm����+D��ٚ�8I�	˥;?z���b)9�v-n�������8����E��5�ӻ���vL�N�vg�_w��UN_����<5ZV1U���kǒ��&4�'b*e|X�Ño�VC�D�7h���j���oN�2��r��D	 N�IJmmSB�ok��d�w�����C��Xh�h֍@Y$'���6,��f"���`����h�	k��gj�k�Op�n�����/G�x��ɝ�?A��b����Fص�J�~���0�|1�:Hm�	�H��3�9$�.�f��kz�"2���V��6���=`�X�ړsC��Y����p�h�Ei��νTL�@Yv�q�'Vr;/'._7a�1ɚUR�[e����uUd��y9�9�58l\���'Tj���v�&��.��,�}��x�4Te�j�44�1�>����!��d�8����lT�ƨ��u�^x�R��54�p-�T��1��c�lO��m��Q�c�<�aGL�����J�tw�i� �{{��?0G�����͞�=:g��t�����K
�@���Sl�F�];L�₫�Wk��q�~�H�;,�*\��b���-���ʎ�^�$w:�JJ����:v]f��(�e<oN���G��q�qd�pVZ
7	�2 Z�v�n�NW�B��d�t2�l�{%@!\��f�v�`��?l�zo
빜�ћ����T��߇��*�8�.���:�$�5����kwR�,D40��wN�-�в�Z�v����v��>��-U�Aw�ԫQ.��B����j�w��*�g�Ԓ%��Aم�_+��Z�>����V�V�M�ٛ#�y�R�m�kV�v������v�K�GgJ��ŤE�FV�Z����Gٛ����\'#��M�;DӰ�^�ve�:{Uz�Qn�\a6���@kG��Xvd�ez�.�uV�U�rVV��,�Rú�Z������:���Ct�e��e�>ژǝ[Y�u�N �c
G����G���~j%����,����/,�Q"����Z;+���'V6G,Q���eH'#��/P�2��6�4aH�6cu����y�}�%�k=|�I���vK+D��Ѳ�$6{��v�2q=�w/Z$s�����r��{�Kd�+ߊ�]ݭ�s%{�z�ޢf�
s2��#�3B�:oRy�-7��..��YԢQ�A�`_pp�+�I�r7�������*����c�Y���w�YSd�IZ��e6�}�?l�V���!�x_x?l^�����O��S���ٖg��DS�>��h���qP񙠝���|n	�X����Ë{v0���n/v�6	l�n�<�[�qHt�JL���������]���{��8�3�ÇI�k�v���bܴ�C1֧��j��YI�Μ�Aef�UJ�,v[us�'�-�[�J��F��Xi]SE���>Ǆ�T̥W_$F��׉VÌSW��R�%gj�޻��6[��]�@���*����Ҙ��9LUq<[��'�+��w�� Ey_Zm������~)�� �{�ˢ����5��b�Wvl�,�w`��$޿*�G�}�;ʅ!�A��b�vڄ`Nn��7keAf( �W�������������,uƝ	kzɼ6b�g{u��uӓ�s�)����T*�	�V{����g<�<�_�!���~Bd�-���9pM�3G��Z�zHͮ���u���m���vw��lh��*q�n���f���Ȇ���]#��0s ����8'��	NW\m�zl;ki�z��˞��|c�;r�����7Y��nax���Z�Q�V��u��M�{p4�I����n6�A�[�c�!���9J�+�*��5�x{Sr����Fu1+Ctu�:�ح�=c�m�d����8�n��p�������,v<�f짥{�z�V	S�M��k����c/E�ny�[�Ⱥ�i��pq�#�Si��p��ۃ{\7[����<�Ϸ]�����X@��쑟F.w<t�<DԦ*Ӟ�Gn{ϋ0l6Ny���?���U�=^3>©��L߇�eڿm��#ݟ�{�p�(Z��w���������ݐ�;+"5q��v�O��ˡ�����vI
�]�=���z�,���[�]e������;憘�\��N��tS���wTPJU��wf�H�%w�-��h�$w�ͺ�By�ZH�"�Կx�ܕ���=�
3m�@���r笛��5�>�u��X"Ф��s����{�Sw�轫�:���C�W�S^���3�,O�ױ-�O�z�8�ڶ��1A�`�� ��)�ɂ���[f5���r,��u�O%k���VcC�Xv����f�סyƈ�
j�;�O�2�(0��1�7�$x���ۿ�0J'���wh+�ێ��nK��ǩ8عs�z۶b�9�煵<N��F�Z�yN�6�Й��������+)h�;~W�l>ل�͛b/Ws���u��=ƺ���XQ�:J��zϼ�[��&��紩�^	g�*9\f;�_�^��A��B����L���}����Ԣ�*�fnW��
Q� U��O��X�x����1�{MY<)�rT
 6��pmԨ�4�׭�4��������2���ࢫR�H!E]�LS6������AB�gv�_��
Ȭ��[�3�j�Ï�fn��)�a�BQ�,�;�J�V�9P�e�gc����i��vZn���ӎi��[���pEg�yf�X�M���usu�=~�­�e�zIJ���M�6@J�ʻ8�l㰦�"�r�-j�}��D�J��oy��<צީ=3طjiah�[ӄ����b�I8:�Q�]��[+���x����&-��o,��\J�:P��J�D�dWj�ݍ�3�rȭ��Wװ"��{2e�T/��՞X��^��xɼ<��X�uܢ)�KS���Y�ј;;��\�-jP�uo��������ܤ+���/�Ѿ;���޶o�G���;��d�]�r���';{rͯ{3�0F�֨WgB��1L�j���1�̱"�O9r��Rnv��Nm��)��s��(rs�H���e�r�=�U��_�༫y3�^_"����L�n�\6ߢu��=�횽�\sQk\�3تl�WKk��Z＜�>��:n��vZ�8����h֊Z���~BnQ���HI���rn^#�*ˑ$!�:w)
�hj���8��i��73]��a�?q~�n'�Ziyz����O�s1nQqgq[ϻ��Ê�������<�|<��陝q�]��t܏V��6���u�vu��硢x�S��~�_�������v�����{�s՘'��w�^IJg��v�b�&4�D�Lc� ��6�
�+�J����OӠ~�5=�����j.V�~5Ǝ�6����/Ӛͩ��{���̅�E^�p�mգI���9u$� thH%v��}�[��;zit��:�M���a��%3���iΥ@`�3=����Oa�pݒM��!u����Q&V�K˝{�����.^%%t�;���<cw�P� _p��ź�iZ�BW�g�f�{�f@F�:���z�����)_YqXc#%�X	`l�֌�#m)�Iҩێ�OWP����ny��j���WUo�"E]�a$ Zu�Z�5O8�m�6��^����i�z�.�؞����zEr�X�2����"w��e�dB�>�6��h�Q��=�tl��Kw�9�[7ZpP�%�j�2�U�v�������>C��L�1zRߝ%fg~cX���O��;H(v˞h��:��+��(%��$��TlZ�+B��Wvxzp��ν;Eֻ�5��-%�o�[SM_�}m��U�yo�杷�o����:/��a]�
���
�)^���]㹴��q1��W0wn�#��&���\Cf���޴�r�B��A�Ј�_�t��B��?����~^��K�]�Eb'{��׿�:t����!��%�&��瓹�'L�sWKX��X��U��o\�cM7�W�w]\}BG�s'Y�=榅Z��K��ή�mg����W'���	����}?.���ɕ)e��:���t�Ȳ��R��_�nPٷ�t[G҈#����aX�����v�㝸�buݷ*��l����WM��jz;v�;����w�Nz��Џrn1ͬj��3�ϝ����v���̐��p���q�6"��l��L�&��ǋn��(��N�Հ3g�vBۙv�%T��v�Վ��9�w[#�G�]�7��1Zb6m���I�X�mャ	�ƻ;u�.�{ x���[�{s�6駵�Q��Q;c��K�\��z��lcŶ���I���4Xw6�և:���*n{��N�R�K�)r�� ��E'���i1����;���6��yE��罛�;w�,:��fz!��7#y=�HKV9eU����M}���X�Q�f��(�z���V��j�jc���L�<��0�_F��W�s�,vX�4��R��+�Zt��*²�f,%R%*o/2��õ�;��g��S���Z�Y�*b�K��Qz�G\b�V�L%RZ�����ha'$�[�0o;��ݬ������^zI)�y3å�oz��{��4<��r�V���̝�{��Q�̶��M��-Pr�׮�ٝb|�s;�pN����S׎�k����򏟳�OX���MunO5���uv/w��o�����c�8���xjP�[�e��ٻy��[�O74ʝ��Q�̳�^�F��ɿIgٚ7��,�c)�N��X��|UZXmݭ��/�ט���wRӆ)y�ݜt�ˎP��h��VM�,�v���-m��x��~��}������L���Y��i��h��������g]�a˸�@���-��d�%����EEX1h�*�\��7*�6f�����Lp�ܭ�������!
b����Y�����N��Dr��W�1����5�Ѽ&�5�i� E�N�߉���~2��Vy:�H���N�ܶNxc��I5�<�-M+�;��m�U�����$���c�[�I�қP,��@A�1��X�+B�}�۬O�^�cЍ+fA��f�gb�EO���+J�����X�e�(�\=��f� {�w�twӽ�y�[o�ǾG�a�]�_�u�ja���5�l�R'ץ����@�fh�7V�Ӻ����a�B�粬��^�:���h�=2)�(�U��"K;����s�fv�5f쀭��z}.�ќm���9Of�]��xب����T�@����H�M��J���X�5�Va�d�Et�����r�]��
�}�j��'�/32��G�
�x
X���p�@L��ZB�]����
AŹ�;��N��%�l��Z��W�ksJ�jv;Yp#0B�4���{ڄ�o{r��E�ʗ�U�cZ� [r)�j�p�[���6l����v����/c޵�Y�om0�w���qG��h�m��}h���s-�Y,�7v��6�)�y�j������& ��;c���vվb�� 8��Cᕹo*�m��Z@�n��N���QZ-#Yzy���<��K�xr�8��^��P��2��*�
�ĸ`թɩ��]X�o�lk��)b7-=���K���q4�욷����9����.��0�v�?ǎw�,��s�2n��wD��L������n�����Q�(�d�w/��h��������o\�`M�}�o�R�ei�ۋ��h��c**N&�"�RV�qT��:��gk*�q�?<���fF�c�|�	k�,qR�-U��Q�.�;?(b���un,�����2�٬��C�S);��%�IR���}ٗ�$��.��AL�YRlR�3��6�'�9�M�:��`j�΂G "�N��/,ot:s�:X�壶��Z#3���p�(-w�h��i
S�z�E�[�h�o����E.�b3w	�ӹPvD8#�l��RiYW�6w:k�ˣ*�k�g�uJ�iN̦��--p�J��J(lWZ�a{����J�Ё�S$�/��67]Y�
B+<��hȮD�w��;
%���xW���	cqn�u%�W:$�R��&?�ntp,�^�F�2�-���,q���9����56C+��32e���,�Ћf�zs�NFYB��(�r�d]��e��GTI��oVnU9��Oɩ"MX�p�{��Q��e"�i�v1�{�����V�"Y�Q33�gM|E�acC����
��^j���Z��-�-�iߚx� �_���<8!��//� h{�^�dW�q\N� �kj�AFR-�=JDJ��xh&�$�Gv��� �����?>M�9��}�Sw糞4�d�uQ�]>�n�6N��۶d���N8礊5��[�6�K:�؆�p�:d�t��fB��.҅1�i"Ko]��r���e*>fd��w"v{^��-&�H�H�(���N��9�O����2�]��Ah�D�Ȕ��$+�}fL��Lwy�Ƒ���,�R�(Ip�$�e9=��lB���P�b�e(�ތ�D"�-D>vv)�v\�Ѷ���&�E��P�u�VEm������1�*ylS�;�"����}%˙��x-zJl���N��@��,����O,D��هظB�ϻ6b����ޢ��n�{���v�X�[n)�͙>�c|l-��#Vy�՝{ʄж�B�O���¾|�F�ciI[PjNC�o(�,���!Vi�g�k�6!�]+�X4Ћ�K���A!�vwH)�C,���@�J���ۛa�
!5��I��$�@��}Qs��C����+F_{#|�m���Z��ep�Y�As�lĄ�u�(�,��. x6Vհl[Glx�J���S�Ñ����A������Z;� hF�e���Z����H�P������+}���]��U�)��'f0���O����Lr��Ϲ��@��Ȳ/k�t(�T ������_uDA�A��`�1����g�:��cl���!���ͩ�D��R�����N�UAX�Km�����rq�{N�Uw��+�TS
����*���xxe!�oj�o9w�|�>m�)�I�s��+]2 ��R�a�G.�\��2��a��Dr�|�j���y��boi踋VCn���&���g���c�#d#%��6})�;�i�C)fwӆ�ٴ,�J��4+��{�6l���[�O���^�=���u��K^���4���;#�4$᭚��W�78�O�Լ�}��q��t0�d�z�ማV����%Ћ=�x�6J�>l�n�ug�r`\� ,�����R'iY#�z����!���������Rs�`�W9��:��p����M*��I^���˵�2�#KM8@�E���A>���ä��}x�Da�s/�gPC�@�wp��a���� mQ;��e.���S|��V5R/ڲ�t��XMM�WC���.GA��G��-�ܓ��+b�0��*q����%�vd�'��pc�)�;[X��'�fێ�Nmd��\5��vC��'7Ȇ�t��:ѽ���ͱ�plqm�Mv^��H��۝�8q�;1�mnrGAy�n4�����<m�zp^�6^��97��y�rt����^�yrb��]�i�qv;rpZ>F2 �\r%�VvMۍ�g�G���n݇&��뭶|&�ms���Cl9�u[W\h8���]{ �?}���cnծ�m�a�r�"��4~��ߢ��$�W��<��wP��Y�ù�0���痒�*������a���l��Vƾ��:V���!���΁'y���]���}�4�W��,cRZF�,�#�0屠D_�h}���)[~�n������M�t��ב���z�-���S5�V���!�鹨cf�Ň��|F��1=t�h����e�#��)j,B-�98}���kB��齼�b�=8a&Y	�-��-�h�!�o����i��όF�����5Ñ'J2j�|CYYY��F�#�{HmTBw�B���v�U�Y����X.owZ[Ì|�qS�H��U��(�:���Z��]؞z��>�B�zϤ��O<�:gcN�p����Zr���Q��A�z�Q��ZR��۠��:g�e�2T�A,��]t��f	\&"�u �[�Syl3��~��Vx4F��W!]�*=��YC
!��$�\�4p�m"�Љq�h�y�� ʡ��/�g�����M��p�jm廸���A�r��v�hU��Ð���?&��غN��_I�<B�k�Nk����\03�أ���T�б�=�G�JLQ�Ȫ���8Q���d\��9��em��R����g��=�GUu1�-+��(`��>��.v�ڔzmtܾC����}=���rHrf�B1�*��
ԑ�u�)�����ve����3e���:<�:C[{�*1:�l>�
��>^j�I��J͐ei�|��hd9g�3Q�P\��3�"��}�/�(��p�L�0����m�6;-�7+�#0}��0�BmNv,1�Yr��z���u�t9�bl�B�%5L�!��@�uSH��o��Ed�]*=d_[I���]�zk~���ԎRȢ�ج��im[�Y?c=B:go���g�͑F��O�᠊:�����	|`�HG�i�gc�i�D!��S;�\����D6z���5���r����b�|�-���oҠ��ۚ}Ӽz>�ĈY<��ژ[9�A<;Y��e�E�F+���&v������.`Z S��d���CAC�wS���c�+���揧uֽa|%~���=\9�N4o!χ�6�gt���Ϙ�r�	�O.ܥh�֘���tY��;<�K�����Nvh����?gy���.�z�Q�B�y�Ǩ��Jץ݁���rƮ�)*A�Ԛ�z��ty�Q��$�C2��$Hv������PQ9S��$K����Z��tޚȰ����8]vq�#�bf�a���$7k-���7X��#M��A���dQ��#��T�{�����2	�8��#��d&�jeT��ev�ah෴�(}�b��z\�uF�Q�Q����^AM��w�mtw!CI�u�8�ƕչ�BSՐT嫢W���W��\�R�'��:��8QAm���x��P.-�/4#��;gr�E`��l�4���G61�|c�}��8r$ˡ����p�R�a^-���	��2�&�s���;;�8�+/o%�Q�AR��e(-��jB4P4�q�I�H�g5���v����Y��c��	�j�8��^���A�����]�f�ɁSfD��e�� �1�΍]kA�ps*�7�f�\��!�a��"O^NC�aM"l�c%���qa��d�2LN�r�T~]�w+bqE��#p�Io�ND�\��4r��Üv{A�W��6׎�0�e{J��;e�Z�F7-|]��dkj>6�P3�zl���1�ȧ� {zϳL��mb�%��z�F�cM;��K��&��Z`���N��SP1�� ~2�d�}ARU%��K^r.g9�MG��L1��Y�!��2ls�nǂ0��-2p��=��!���N�V���9X���m�k0�!�Fu:6\�%Pr:��b,��ɶ���ad��Uu4��8I2�Ba<�*}g�B���ڞg�,��HT�H���೏H}�q�C�F�� ١hY.E��z+#R�5Unٝ#B�6?�s=�=6x�/Y����}R�p.6�sYr�Z�?!e&�粓����A��6(��_8�;2��N��l��>A�6�wV��UЁ�z�̚�R��g<�d$V"����5խ�޷]m�)dЩ�(�|�x�I�oKG��eH 1����X�Yb��,�_d���C-"�}�����ZbAc�ٶ+e�.mH޴?#�Hx{փ�
���W�VAi	��Qda�5��cK��v{�$������&�*��Gl+��:�F���7���x�vzn��չ$��lh�u�v����(۲���6(`].��#d.�ʗ>�D��Ӎ�0A�맑!�EǟS>�(�˷#��H�}�D�A��ja�ث{mV��8� ��ֳ` Bׂ���l~V&����1.0��c���0`!�<�o<���35�@�"�:`�0\��ͩ�c��'���U�5�l���Ϫ�o(���1$e(/;�/N׍-�yϻ�-��Ymn��б��"Y���(KV�b�ic%D^0�0��r�&��W{u�L7B��퀂1u5d��$Ί���yϫ_��Y�a�G��й��mj:�;- ܯ*�í\�ϸq���+!�v���_0ؙ�D�7�f&�Ȭz,��7��ާ��Z��Jf��5�̞z�K,�"goT�M&��,����Y+�@UݕiYu
�[|��Eg�_/��+���6}�S�������({�ϲ;Si-"c% ^zy�q��A��q������N�#a!�["w{����GR�*U�͵���i0��o�<��W�V����.�]��j�IP�T�r��ͧ�t��wk� MM̄���K�j����d%Ha��t<�i[6�%�����teS��9|��ܽ��9��uO ����㰪������9�,y�yҙ{^�'B����'�xۧ���k�"v��_|��n܆����/�ס��Tw����F�wFq�>Qq���v/1�nu��������k����Ċ��˻�UQ/S"m��3a۷B�'&���Xɹ�̸�8�g���(����!Ŏ��w���K�tC�]�����j+��5k��l��1���Q��/Q�G�sMM�,R^��#g�Z<�Y��QE�AsD"Y�L�;Z䏽�,�3�� &�9���ϝ����~k���o܃�V���V��MK�J��'����6XU�����a�,�3�i�� �'��tt���h�^�`���B6Ͷ��=��S;��`{@u�ͺ������]!���]gMsq���n�c�eeo��̔Fh�
:⺢zMI(�0�����9�dA j���Ku��4�Nm)
m����fBD0���0��<lّ�|�6T��v����>b0��y���0�6U�SQ�G�,/A�2;��Y��r��_v4v�4� i�X;5���X�4�� p1��Ȱ�:vAS���
�%�1�7i=��s��'�d�]6`�t	�ݤ_�:��ӓ:�='��v��Ib��h�@J6H��q��d5�6#�� '9��l}϶os�oNE�T���V%6L������xI�q��[�e���=v̛��۞\��MS��O���'y(���h�Ҥ�Ai���?vA�S��ڙ�ĝ;a�m�q����؈~����&��;H��Q�Ư=�؏
墙���F�����d�rן�o��C�%�"Q�k3 \��KC6C�n+G��o_ǝ���j:���YQ�톰�)R7�.F�Mv�]yw��rM,�:��G�Zٕvsk������}��RޜQ=�ϱ��
R#D=�5���I{A�LkIrћ�A#)��4g.>�K�%��̀]�1�-�S��ڪgN�@�҉j���FyoN8DI��aע%��N򑘽F�x�=h���	C0���N�ųYd0��'g���98e|ᘴ,ǖ�5�/g����,dj�t���db�:~���t珃f3W���("���i��V�by�˂aT�ݔbI�2Q�]הɈG�a�4g@t�&#
���Ù+��
Ѳ�\�f�cV���4C������ŀ���k�;32�bIe�5m6�_�#^�ﰲSd2;����g�-;N�|S0'Ҫ��sP��0�!����ߓ��r4��WO�ׇ�����̗Jܳ��b������Y�9��l�\�LγH<��,Bĵ�E] �#!\`|<zg�hZ�1��cپ��l�B3�^��c<���eI�gz��Q��=�����^��l,uA��M-��ٞ5�{�����n�p�����m�+˦����At�Q=������R%���"c��$�����bGL�E�!�<�x�����$�/�:�Q�.ws�Y�4ώ�`�	4f��~��|k�������ϻ=���x̸�1��u�(�h���*c�j��,-�E2m���<���.E����5Rn�LNɫʛ�-�{�sdD��Q�m�L!n��+γe�
�ٌ�1m��9]b��.�]Ԗ�K�wq:��k�f�PX�r~��śďR�ۓj6���Ə��� ��8�s�%"�� ������y�Y
�l�.�A���D[DsEcՎ�������{/	Ҫ��H7+�fL���.0��a���٬�[" ��=1�G�P�d��ێm�8�2CR�=��/dI�^J�m��iq!gȣF�����Y�牁r౔w� ��Z���Fݕ�*�=iۤ^k���*r��޸�=�8�v��L�T���gg;Ấ�>�@�Y���'�>�BH�;�)k�G��1�ܤr�s��uӧ�ZE�zh�A �a����9�Z��kl��۔��8�,t��WD�
'��l���2��-Aޘ9�+I�o�,َ��چ�A:����A~J�8Q�}��:�mM���מ"�>�D�U{�l��ȺrZ���.Ƒ�����x�c>Z�*,osY�בsS#����23}i7ƫ�Q�`�TX�^-��zh&��x�,6�;�4z���Q,v���F��n��[�A�ꉍ�O=}\c�'u�.�g,�u \�D,#/ �c�
4I��*��'�X����y_]�v���K8���Q��3igI��"��4�B����ZGt�p�N%�5����h#�>jL��l�g"ȹ�_��������k�YL-@mOB�����\)�Q�\�N6��z�hF�0���0���/����G��N���3'�i�8�&���w�t�c�9s���uB��*���;d&4mι�>w�n��p���;�pk�}͝�iWU�_���T�����mQ˔;q�%��L���"	T�]�}�Q��=(Kw52&e����x:�9���۫�DYe$L��5�y���U�ҡ�fW�#�a#Ko�ڄ��~�Z�IZ!ȁ@Y/�(`�=BdD�������#z�-V�H��t:�������6�96'����� ���W�{���e�;$Cgu"M���5�p���k0�;�#L��"�Tu��7����V���"o�b.���H�}܀��!�� �d�f�ɛ�[0�yv'�2V��U3e�ҷP��3��uܧ�68���w�H"�A�� ������"I��2��L��dIF�.ٕf�'O bf�k���J���m#�I
ۤg�>ZA�T� �.��@��i�m�t��4� ��	��q��x��%^�9�I�������%���I��r�a(3�w�'Wn�G��!;z��	���Όt�X=U*!��_L������C�<M��nf��ei���L#^�7c,'�wJ�MZ������h�Q<��T-�D�o,)�ir�"͊�YW����ƨޜ����u,��_e޻�����K�)�j�����jk�r�R���݃(T�k�9jWb;7#��k��6��.���P�(�b4}R<�E�w.��٦�t��>]���7��/-,�;�JP�ƅx?t�s	B>�m��m�c����43<?؅%*G�͙\k�o`:S���Jv�r\��D\�s �%>�����/0�7��Ϻ��٫F�$U�1��  ��@Gn�7yd�B�Gz3f�=���e�3E���V���k�����yYD��*ك��쩕��	d��R\�'�K�a:�wYj��g4p��Xv�U*�/
�Tm8�+\O��a��5��h��y2�=�}K*J.Vc���P��;�.��)���+$�z��{*>�E�fj�M��������]�Aw���C4!���YKe٭�k�ЦC������6���=7ȧ)��kR��iD�%r�ʝ��D�e��Fܵ���݀{ƻ�@�VCn^$�x�)v��L�>3�G6�������'�F]#Y�d��ke7N�զ.��m˕:"2s��Y�nM�{���҉ڼ.t��]��s/F1�"�]�r#�R�IP1�]�nu6�zDknL7`k�y}���(�,�GB��d���d�wwwj��H�J����M���!D[5�F����c��t�[=�����vxu)����S�,�Z$L5IS��Y[l�U��j�/. �sfv]۵���!�c7�l��=�z�^�F�<�w<D݄��
l�n��Şv�x�����gq�ۛ�4طU'u�ӓqs�Jݢ��7Zثz�8��o8"��Ұ+�b�]��Q:M���\�9�X��m&���p8�wb5/���;���9��u���B��՜Jm��<i����X'Y�wX��0���e9�86�u�V�7� :tv��=4k<�l���Ӈ��qe��k���� �F�1�~��/��H��[�7�����ΑgNuxutc�'9�q��Ksv�]�=vz}�7���p���u��ݙC��7^d{�M=���ٮ���n���`�\���r���/n�li6���6�wT�\� ٬�r���Ij�y��{�k��u�e�/�7��͏n�����RѴ�����}`cg��9G��A�W�I�;\�x�p1�{���ZK��kwU�S�8�t;<�c�w`����vV�*��f1�G�������9�Aw�:|��a���N���6�����חq��qn�mn�rF�V�׌���:v;�DX�"���##V�w,�Ԯ{�l�������H�p���)m��u���[N�u�����n;�:��7Q��/b1�]'Jkj���rv�6�۴�<�����.����2���`.�wvk��u.o0����ζnO,8\�T�m���rO<Fby/Yx����ۛn!�=g`4:�6�]lOUGP'5�pt����:J�����%���(�"ݱ��yo1�ew��ev�}ӄd�(��9�D�3�^7l�I�;c���tW��u�MB\@]������cg��k]NŅ�xmֳ	ۊ5��c<n�lw�\��}����[ϝ���Ƭ-�bw]�-íbԻc�><�['/Oj������@�m�����	��x㴾���`���cs�l�6ԡ���+�u�i{m�&*ٻX�UUe��{Y��c��rp=�'�M�����[eG7=��f��ݝ��&��_�}��v�������Ӻ�]һ<l���H�r��ݪy�޵�<p�Wt�m{qq��[kdܲc6�X�P�NH�N
qĻ����W7�����=͌���nٗv�����;�&軶�O7��غ;k�/^��d���Xۦ�.�K;ѻj��88!�u��'p'�z�۰\�L�� t�mF�"E�\�l�
1�v��C7b�~;��9��B�c�S� YQr�~��Ԍ�>�m����$�u)��r[�L.�OlL��3<lU�hV�k�x|��kʱڝ�'U�W��ghK�RՒ&V�0��*��B��	����޸F�B8`�ݘ.���55�1!T�7����Q��"{`�sm�b�=���[�u9T#E����X��ܗ�h�}P�	����N^���dtɴs����0)�<sq�˕Z����X-�����l�����a�n.�
�?40VF�%������kK�l���O�@����v�+R�)�$� �l;=�(�Lb���N P 6�e��$�*�<�l��"��OH�iq��9~�,�)����We�&v�F�M5j&HQk��Y��n�K��o�;V3��2�����[�����wRځv`H0�\�6�,ov�xl�o��^��T���-��FےH�o����z�IѺѝp�t*v�	��!�ٹ����H'��9^׍��|�(��7�ok��HP�/��	=Q�ʮ��$<cIc>g�ց-�8�Um
�-��oȏf �;��H�!��#4�$DW%�R�+)'��)��v�&N5�Ŏ�c8��B��_���K��4����u��n�����/;�����C�r�!xq����v�7z�s��gʜ�N/�;۷F|�n��㹒"���� ��c^Cڢ�K ���t�(Ic����tlۉ�)1��a�>�(tY�<�#���v��d����3v��'
O�M"m9Ғp| �y��N,  ֔�p�v��A������	�ñIn�|>���h,C.[�m���Ku��qAJʣ��Km�Z��5�#����մ���A�{�>�\|.�4i���H/���9A=W�����:Q]����}Gc6��CB}&Kc���d�:�c�;f~��>@<'�}f�ĂEh��1%�z+��5�:<eu�����qpH"٘���x�CF�x9�7_�G� fب,n슫z˾��?��N#>��=M�pj��S) t�4cn�{(-�����Ȍ���T�Y���,������-��������aDv �R뷹��y����(���iFBwޔ��	��c�=�ه�o� ��a{­�T�e��&�sq�Ff9�MGo<
�U/NK�v�vj�D)&�P�<�I��@d��*P��.� �8\!t\�"�/������$���1��V�E*n[0�h��R��Rw�}dzȷS��O?�-�%��h�K\Xg�:E�}9u,iʐ�t�L�fK����(=0ڇ����}��l�;v�g���j�ꟑ�U�R�ͥ1ܭi��ž��\;�*#�t�.B8DF�ٹZ>�>P�l1�.���%�p���TO�%��b�(�'m��֚�::�N�[�8�:)�dmzK~�� ���&�I!7;�UwSHV��
��,m�#���u�{��z|`Hr�D�*�ʢ6IP���$x��]u��3#�q�R�D�l?��^$�&��ȷֲ��j�xF�2| ���.p�>�������2�W�P�
}1��M�����Њ������qK�����@��y�oK�B8���{0���b���`�͸җl�I/~�v��GND��<{٘YӪ0EvorO�����=cP��ؘ�2�ׅĽ�	��k�y�
pM���tᲆs"���Y���ⒹKA�Wm����
�	�����ö�߰��a����(���1}�� ���H4E!�=���xy�;�85�G\_v�u'�����qb!�Յ�uIe��0lg�nŁa��|𖆈MM4��}y��#�����)Q��Dg�獟53َh��Ml��!oME�`p��#K����Of+	˥u
*�����k�2n��::�f�R�X6�e����X����$���/2M'WHi1��怌���a�N���W��!��90�W3.���n�iW��b���Ϣ�;>PA�H���>+#�D���(��'��ՙ��itȩ�Z��r�A��.�ēӓjt� !����pD;�)��4��եD�m� 41myZ�O����iEHA���7�W{W�(����T�>�N��n�q v��Y�$z'��	r�Qp���g�Gr�xǸfgo�pΔL�@��Χ]m�瘄�r�Q�;+xesra;7�[v�vԍpd��R�%���o���I���`��y��qc 	�BNZ��`>%�6B%�ft�z;��w�i�E.GR)!k��gu��C���e3�z=\��$��ْL�Fuጄ:�V�c�::��F���L���g;�"�n e)1}v�(5Y�@�A������}�F��v]qR&�V�#N�E���C5�b�5׍#G�<gԣ=�gx�+V*>�B��lav�,������[��8F]cH��b=�c�z'z�A>�V��fc&����]VWU�F3�'yF��F7�m����bY�M�M����Q`ȼgsO���"uO(�NL��%V!>t;�4޳ʲ-�� 80�d1�(�T�[�ۜ�M*`M�׮�٬���Y�*d����g���� b^D�F�!�Z��"H6���,u H#�bZe*!����;F���0�6�q�f�xi=���-��L��&*a;����@H�%�Cq�/���#��m�C�6Gv�3��vM��0M6hb�]���Mʀ��Z��%�J�^���	s�e�˶8�O%�^��;\�I֡#����m��]�lEۍ�Wu��Apܜs�n+��q�/ܐ�o;���n۞��].^1�G��Oi�8�y�m�Lx¼�s�Mۉ��8w=�@q�ϫc+���M���x'��8nf76�@'�4'�)����o!(�ٳa����=�[��p�����y��;��Iv@�	��<;m�������]�F5ɽ��$��.���qfL���Υ�;�=�P�mY����:�c�F��}�JE�.P�f�	4S6��\�N
@��^�3Ւ�&l��p]��i���,,Nm4//D�4S#�y錴˭�rm��mM������D�NFCBX��b���q+jQ��f��=ۋ�zj�cq��'jS8���R'�2'�$Azg�L���]���xmy���u����7	��sS�n=��;>�]�r�}��d�rO>w4y�f��ն�
r��hj�f6d��t�,�vD������hj��\t��o��Y=[E���u�gv�4F!��2D�ڳ��t����=���I��Donb�v��d�cIm[�nzoY�B&\�L��R3v��Ai��4l�m��#��e��>16��v1�l��[o�~kF&7���>$2@��u���+8�v�6�E������hk�Y�6U!=��(�"O��[ęx��#QN��^�]v�n��W�^771��H�h^G^��3�NFA؞ �Gq��@�vX�>�$j&�ݮ$3GM0d�/sc0�g�� �[�6`��b�����Lg;��ͷD����d��M�}�qb�P�A��4�����'�b�Xɘ�vx�Fq����p���P��;1��$f6�[m�UY۶k~�ݛO+��4�i*[/��m��Gr绊�mU�)�2n.���\x���`�0��B�ډ�]竅|�Wº9�W��y7.eeD���Ԏ����H�]���c��G���D$���ţ�t
�:���k���-z�6��Q=�eo,���$>��!�z�ďK)���nE+�Ê��ŭ1z��H���U�0�]k�u1�\l
�A��sFj��z9j,*��-���R��/oµՆ�\Dp�Ě|�P$j]���̓��Ȫ�ԃtQH��ZՑX���L�5.��A=�9���M�d�P�F�[߶��r���,�ap�����1��I��^ҒNj�`j�wa��\75��GV���b���Z2��	%{�:T �A,�Zd�뀮3#&L_@�Av�q|�i�*B�ʘ�[ۜp8!�{-�IV$J�n�P��X�(��!K�� �$��b�t+Q]��酭����G&�#�/�z͟!���N"͠�&Y�ڽ���"�ד�8��`��� [sx��⎡��+r�-q�D42gA<���{l��k���޽˂,�Q�f�qXɚXd��,�=�O�:Bez��E��/6l�/�mA���9�x�}��F�3����6���bS;Тq$��!����q�Z�a��n��<����(�Q�gt1��������ƺ��t�[i������N4�_�Q��37 �kb�ݢ0嫍+�;0@�l����. ��D�����/��F�u�Y�J8GV�q�zٷ����/lӜR�*�@�V�2(�R��jpou��Y�Hv���Iԃa�w瀥z�6.J�|�/V��,g��xGd�8�>��#�2َ�wȕT�U�lr�}��o"Ʀ�9�馁&�r(��r������<x�15M΅(n�r�E�1�4�.E��e�gaGĈ�㦠3�S����ly��N��:��r�p���wQ�������@7�����.h���٥�6t� H�Y�u�<��3�������mvۉ�,E��TRc�;��q�#"ׂx�:X�T�$�D�1�a�ݾ`�tȮUO�u�KG*�����f���$mO�* {T��_i���J�\�h�O?���>��OK��
4I���,OuO)��Ԃ�^���w�AS��V5��Ke�p	KmY]"�t�HK�Pm��0�8EN3�a|��0��)��f�o) �W�	h[���k�y�r�J���b�3��4�%%"�\_�l{X�7��Vi:��[�Gq�8f���I�Ѕ$�A�5A�c�G�2B(�x"�L��8�T��t����w�n�.�g��2q]-enE���Ǝ�*Z��6�-ѩvf3q��ư�CBH�(��{�r�J��bdW?YhM�Jm�7��{���|٣¿���y?L:*�r�Il���6<
��2x���������4�	��!����@`}��Qg�Bsg�Ӕ�Dwh6B w�is8ؠ�(cX��γg_��pݖX�$lVr�C@6��
h�;v��G/:v�6�/K�r�<;��n@@�0���C^���9M��e;57g�V�Q�6v�W@p!�a<0�޶��Ќ�ɂa�Q��F:|��1���,�2B؞���E�k-���N[0��N("έaDm�Ge��lN��<'#	8�ŀ1�ƫ��MK6�.�AP�P�,{�)G�� �0Æ�����I���n���ӷ�.,ίq�|=x�F�A?�"�d�"H���*� �K�m��E�����in�xR�G����kC�Bf�I�=�\�8e�۫�]n3�j�>]�5��"e�G٬�������A3��Y9^�̊Υ^�ux`҄t&y��H�^b�,F2��2~��1��͖������k��-�N��6�D{[߷�;eNVT+U�W��==�
���ּ��ZQ�ȊI��T"�٪:��\Ic�9�i��)���5Sf!�,��{o�I�Gy�A�Rv^31M�ͼ�59j�&�;��>t5���R�.�w�讌�)z�ǑJu�}ǁ��튋��S#�bQ���?��b��=��%�t��j�1!�Uu.9��'2��AcMfC��j��ݲs� !2v�u���cvt�t��ψ��sY���w��7g��x�]F���{m���5����u��")i\��<��mV�ٸj��4����ƞ�0OmEv�=p���xW����]l�r�l-���9�OC�&4��	����
Nܛ�ٹs�}1>��V�'-:��m����;r��j/l�ю��r�i��<��Ӗ�vz����X�-C_�C��|��5�Pt������$�9��j�)C �����)ͷ��  �f9��"�ȍ3!z��4���H�A��N(\̈́#�RF8v��ljL7wETēt=>���������$�]�%a��0m�(�D���9�
d�����D�m�qW�N 	!�Hv'���W0�/��ا��5��>�1�
��j�v��V�C�AI
w4z�Z��s�3�<$%�,�~�*sk0�J:a�<)��m��?f��ƶ�� �0)q�F�댐���+�����������4�@���q 5+0l�Y$���&՗"�)P}Z�㳦Z$�D:��-Aմ;SR��$�!s��m#�7d�`^�lו�WSj��W�$(�QHI�B���Q�.���C�4!���͙�$c��RD�4�!�k�H�r�`��z�A����COudv�B�Ǽ��sSs��T��y�p�x����n�֔���v6ݲ;��k�qEiև�W�jbF���RUcq�e�W�^x0x�H��;M��,�.CUC�	2Q���mR@�"O���E��<:4IQ�\6 b�A�jW�����!ӑv�W�t'ҷU-U��l����ĻZȯ}����+Y�̲/�To�ϔ�,��%�a�=Ҭk�\T��v���w���6�y�xn�*���ՀD2���uR��=��T�򊸳�9m7�Х(:K+����S�N�s� 9#c�hE��;.���8��fr�l�M�r���^>��omd��ߴ�x��u>ɰ��=l�jF�޷��F�6I�ܙh����؀iI����q��.e�blZ^��4�n؛�0����&I �Jr(�OeWK@�Dq�Ur�I�&���~h
ՒL"Q5��hp�������/��A��;���<ڟD�����}QzHEc,V�d[(
�q �o8���vN,�	%x�; �6����=<���)!1	n�q	>%�"�0���ꁠ�:H	��\��;w����q:�"��cU`v���"ŷ'=^Nܞ����b�9n���:�7F6�'�[�a[ں�r���!��rȒA$�g���>Ð�G�`!��+dQ���2�E����_��o��Z�K�#�B���ZŐG��h|#�s��N�M�ݪ��m�^}���^0��n�|�����EM�2��z 9C`����hڛ�E��H���h�0�{�2M�H{IKYgQ�o�^#㨎:���	+�Б�E6��=��y��=� ��	�򟹤����A��֞,�;�v5?&���7��:�s�l�Yɖ�J*�%X�\�h���v�0��&�������hf�-����=��PTG�/����|��f��Zɠ���4�i*rU�a1��*O��"��x��o�`��Z*�N��ꄬ��>��m��y�%Y{�M��-��&��f����5ΘX�s�X���F�k|++��k��d$՜��\��R	3nF⫭Q���pƌ�okvn&�pb��W`�:DSgb���9P�]�N�;�jf�E���/��*�6�%,	V�#�����2�%��s����!	�r��V�p%�i�سo� �iw�\ƃ�郴���m ���Nn�/�n �nT@6����F`��:wlNL;�g�q'�i��Zn�s�_N��B�G�"[2]��J��4�빑*aic S��e�N`؀��N#5˥el��,]�oW��lnp!�ذ豵��F�sr���Րƍ�L�u�W�s��+ �$��4b����0��oy!X�s�("1�ث�OJC������k�M�q������ܷ\��2���Ͷx&��	�������Xn֏ݦ����u�և)ٹ�a�FX��0jv�"�A:��8ʗ�z�Ge��my	B�qQ��ݖ�g�����6�䒔v����6�k���4�P�y�:�6��EUʱu|%��9�p���S����>�Mc9%! ����<|�Zڍ�:��^����+�&yȦ^V'ol0"�ş<&�閑D�掠�� �u�)�7�0\��)LD�T(k!�V�e�jT���DE+�e�5�91i���%��|�4�UR2�م�w	�[I�}�s/?p�4v�b[R�O-���@W�z7u� 9�T-f�F�L�B$���9oCL���t�>��"����G{��4=&���w'�7l������-�O���m�v��[�ŗ9��qh�\�st��~��8@ҋ�t�[@�b�ñ�a���Ǭ�I+f��:��ݼ\X����Ӳ�:�C:B�����߹�-EDuA��V�T��bN�Dlo\�"NɑG�]�$���fD�#jޚduczH�Fj�n�h�@�XQ}s�-�Q,;$6��J����S�ނ�B,X��!���.�l�g��K�d�=I|�ɣݝj=��nf�Yxmspp�0�M<�����5���c~u���}�k�
8��-k�?T�r�Jܳ+����'��f=�!�E�4�'�2 ��$�M2Օ�1Q���&���>�q����d��|��QW�I�gϙJʵT%���z�&�`v��5'�ݧ:�j�8fnN��2MͲjѮ��E|dfm��ǲ��t.��x}��A0�Z�2�GN�섕�D6s���Q��۫q2|�����<�
�g��ݮ�E�K����-2C� D�^h���h�Єq�-����*Ӷ��W�_��۞]νH���iD�Hn����s�) D�V�J�g]�`��Rwi��[�\�2�/%b�s��N�.|�����1�M�Ij^DC&&������+�Ⱥ�2}d`�a��D^ո����[��q�
{�'7�l��� �˔�$p��=�M,���*)�{"�X^��Ƅ��[S�
<��fO�6HY�4���h�S��e����#�/�bWYT����p�,��=�j�Wv�)�0���(0�z�-]jr����gn	��>v!�jȇ]���1z������M+���.^Hl��뱝�Yi*��c�cB�f0�h��Ϟ�gI�X�vp&P�O�q�I �����54d���p�ܘ(�m"#q��Vs����Z𼉻��QrFGd�Q�RD��zoMC}���ƥc�MZK�}<�	9n�ć)ˀ0�LQ��}����rT{C�̷H7��ր�n�ޖ�8�� �#/tM�C;���`�p��N�<s*�^Ar�}�T����~�� ��.��59���M�xC�������z�/7.�<.`���Y)��:eͼFfg#�(ݞ��8i/��ŸE7;�C.ޱ�m��51�ix*;pEچ�sO�/*^]��]wU�m��w{�<q�����b�n �ǆ.�����]'<m�c�f.�����a�v���F��ָ�y��Gk�n��*�v��Vul�#oQ�u�Aۻ5���[�E�u��jܼH���]��5���mۖ��s�h݅�N���B�R�GYqK�^�g������H7Wjn�q�{duٲ7mâ:�r���l�<�É9"t�b���b�-)�.�!��<I�a1�&�ra��yG�B��<���M@�x��+��'%<�Y}�k�'*(pl,ax��q�X�C��%�+ i���0�s�zcB�r)�kk�|���Lh�I]ц����������iYZA>$?>�ś>�,��OT��K�q K&�7x�CE%�����='È�	鬈=�O0�/P�*�%�w_Lz|u���
�v��pp����h��%|kCY5�"N�y9J��u���[?�:vYH�%yK&���6������8��Ug?����b�යT
4I�Ԝ� ���P�R��wGv]1�R��s\�1�<2�Kݜ��}�]U�Tujٞ �,2������$��'|���9�*2���usH���A$�F����}`"��"b��5=n$��(�6}�{>�]|����c�S��u����u��q;����ancn�::�v� ��j�N�F��@qߤ�dP%��4.u�8}����G�;	:L6����N�OS�H,X���D���f�{qi��#�� ���v[M�DX9,�O�������
����*�J��y�úĦ��u\�
q��v%�t�$C̴��1*��io�o�'�`e��1v����0f���:�Kwn�T�ypԭ9��e��s	w|F���6Q�醏'+J���@\���B!�O�<� � �T�$��D3�w:�H���n�^�~a]�8_57��i{z	�!+�!T,��e��%��ިI��O�1����Ɓ5���Du����K�̶��Q�:>>�s�<`K��r������ �1	÷�G�y���_+���@����+�C�F7��ͱ&={��\�Ș�5��/��l�����MӲ';^ˑ�m9�v�ɑv���T�ٕ���=a�X׭F�}3��y�6��n��6����u��V
ʮX^��'�[G�=�O��8p2����=U<�ue;2Dm��ҕٲk8���f��]���<wZ�?m|�z�B�F�V�]3ٍ�E�+�N��s�:\��=��j��!��C���0p$:Qe�I�=R$��ĺ@������i�q{�Z�=���:���;9��EZ�N�A�{���ȭ�@vv��K(���\d�ܥ�h2��N��P|��s�"Ϝ��1T�M�[�h�a�ϽL�q��zR�71�����^X�ݖ�r"Wl��h\]>�3e��D45	���}�� �L@#5E�y�����x���z�ZUN]ɪ:{�k�V�d�@,�e�J6-�Ki:;�A��"͎Ӿ��x�S��ƺ�2M컂x�cAiCyFwkOn���4c=����Tp�\��$�ٌ�طG�#Ūo�.n��{�3�
Q��vc�X������qrM�	.oR!�5���=�s�S�F�rWi���8<e4��H��7	�$u`���w*U��	.����4o��k:�)�@$�F��$ʭ�Y=��4Lbul\XqԂ8@�Ne�y�U[icG�n3Z��a�!�\c��sd(���	c���P��X��@�TM�H�-Y�+�p��X��u���\����;�,�a��vw8�pR�,��(�늏a��9��č��h�z� @6Pԁ ݰ�k����N��Ԑ��-�� �x�5U�1ݼ7rޢ��{��y�*n2�,V�Q �J���2@R�����Zj͹��&��
P�'��>���"M�03U��Cj��0��jIx���R�P:Di�n塳YU~���@ٝ��!��I;���c�Y��Ǒ��вaƟ}1�G�6`� ��֧mpI2�޻[x������k�q
�.��t�r�!��F�rAfg>�Z>�f���A���'}������ؔ��ws^��z�BӢ�ڌ���w�$�.�����#m`Q�v�A���o[�=`���o� C����[�ia#����Q��y�X���;��4T�Y�C+%@qn�XV��7O_*CiY�vГN�;���]��Z@�%�aڣI���u�SW�*�D1�t����ǷUhI\��^��c��=��3m�ss;�0$] �րΔ-l�̍ǜh�����@#%��ox��aEϟzy�4�9�a�&c'�F^�jY2�3����A9~,��Z>-��8��m��lw���l Π�"��\���֌᰼�����3�L����/K#g[��4x�&u�Ĺ:��g��`dI
0{�5OJs�K��Rnaً�`����#��i��F��f
|�S��br��N�K,�٠4&�޽VE�׿����㾆6���q�9�����yY�TS���q�t�I��aF�9���m�i�8f��	,���$w�C3'FFXW%z�=���G�n���y��r�zLC-|���V�8���,�N�1D��0"m���đ�
�9ޜ�F21">x��Jk���E�;��'�"��9-`�w�4dݷvO��P��]ύ$zfy�J�.�CX�f�@`���y`:t�k��w'^��@�E�7B��dK8�n,,R��F�L\b#,F�(���[�(�izH���'_ۗc�����N>�Zkv�����P:B"oX"�)몀,��^�dghC]���HⅧ15Hг�����pN���h�f1[|��e��^�4��U���w���kt���uXԇ�X��t��n͸��V6h����\*=�a|�ݶ0��������vCѶlc�L�-��c:x�=����v�ן��v�4I�����h�[v�F�<����5�7F�8�������P�y11��60�խ枮֍����8�XW4�ϐl�q2�b��/O�)�۝v9�s�GFz!w�'m6;N���s5yz<P�4��x\�;/]��ݨ�Hۇ� &��Nm�P��,n6��a8�;K�]��>��H�H�"���"��X�߁֩�-E �6��E�.|�𜱍޷�������!�aB����+{h�7t�fE�w^����C��@;dJ�DaNc�A��|ݗ�}�� �2�m����د���5M�Z�������pSOEd7���E�t#_�Z4��G[a'ƫ�|���t��;�ٻ��v����k��T���U��m֏��!�#Y��p�f�p���c�	QO�0�Y��f�H����0��@&͐G]?��iŉc����2F���u�����e�+h\�ك�if��+:U��4�,A:l ћ��[0�l� ��|�:���DݾaP�:M9�5��g��0F:�0���@tDۂ���T��j-��!��I�,F���zq��Ҽ#-��u�Dsc��S6�^ˇԍ%���7�WVǠ�2S�0�P�t�sA2E���	G	z�!ݮɸs�����܀A�ԏ`[��x�sG5��|��i2���f���
��Û��C��-�U�]v�}�=֔ب������m�`wrvN��)ƨ�7����\z�(;���%��!�4���E�x'=c���s�4�R���v�%�N|�"���"�g�6�TӸ�p����j�~���f��3��|r]j
��_�*�F�ȯ�*�ec��w>���e��rU�����/�|+�]�6��Ƃ���Կ4�k8}�冘&Ӳ=v��>�M?Z]����������NG;۬���a3p��~��a�c�г�k�f7<�Reݏ7E��H���Ķg#w���ޮ�q#V7�.���F	8uL��M�L�Հ��2�zT<���-�IZE�(�Ao�t�Nq�C�NcO��aD�:�O,��2l�2Q#��q{N����1LUލK�ƀ��I��g�s�����2�mu�m$a��ю*�/i��-�Pr/������˪<�x5�܁���ݡܑE��-.�eKx5*0r�y��A Y���5�c�ފj9~�c�B"'T�'L���6��x���u�n���9�W\x�b���˶�58������~��;}��s�!d��;�iy�Ҥ�<KD�!O��T�ovq�S=ֆ�v'�Ԑ'ķ!$91�X�d�@^�`ᐫ�E_�!h��Ϥ�	toJSb"܀��,]<�'�j�V��S-.����w�j�ƏKT�� 3+�(�'���K��vv-y��i��8W����~_����֎Z;�c��vܶ]H�����k��X�K�V�Wm�"�>�0�D0���G�몁yތ��O^Y�Wת��ui����ٮ��af>6A#����0�DQ{�K�,��YA�t�L���NzE�T�(����~����o� �6�����KJ�fȇ�s��!����N����,Ɛ�9���w�co��=����v��Q`��i��3w� M!A�|�=W��z�J����6�p�Jx�D���+�ʭ�2A��V>XԘ���>��Ø,<����Mbb�B��y�M�钍�oIG�%[�!,@qB%����~���U���!�S�+�����B�[��*v�������Dz��@�X������ї��n���A�E՜dg����س�B����h>�8����I�D��Ĺ�\`Q�L�e������'�8�n��K!���$��\�"�YR���?���`p�UF*�ܨrׅ�p�Q���ks@���*�@'a�i���Y��琄f���ҾD�K��<���9ߞ� I`�'�}̜�>jڐ��ɮ��	�b��S?p��E��n���,D�7��9S�r$��L ��k{�
7܂ etʉ/�З��:/�1���%�\�'�y�I�d��H�s	ĿU��φ�����
g�gٯPI�#��#a��n0�K�����ٓ�D�a�Y.&P������G+,C����M���L|N^�m�x���yG�[�*����Ѳ���
-�Ѷ�:���̒{�$kqx��UzL�
�fkM{�]S��!(�J��.i�n}|����R&�@�A�y���g9���o(���䀪`�H���_}�'���5*!��v��鈴���{�=0�^_n����L��%*%N��N5���r<AlLg�:�\'u�.�݉׌ggGb�?���-�ڭ��x�M6}��s�ZF�|�ݡk��w۫
�mZ&[��>��C�u�\��#˧Xx��?�ft�=6-M��9�'hB�[��9�D�X!��^��r̵-�H&I� ���S2�x��6C��#�u�,
~��./ʹ�@�}�,���u��J�v'7��;�_f��$���=�)[e�j!��Յ��c=�D�n�V�_���΂,�Q=�ԦIO�d��܌~>�]��M43�k�hv���b:�z�`�&��,�BSQ��kޖ���,V�7d��M�������`�۱M#�X \�u���<��	m��(�7���b��H9D���jw���s�z*�aG_K��R��2L�j�u��ah���>je�4�}1�w�� L�R����|�95hX�ȭR&B�0I���gns�/s��qE�.����p��d2�G�0eqn�.U�л�K"*���.) �.36�K'6
Gv�]B��X��s�S���H8�\K��j�uњ�D�DQ̈́��-ܠg]�i��e��nm���;�!���c���'@�X���w�"Q�������cy�yu6�Z�eݧ���u�v�oV+R��(�ͫ-�498���8��C�|qGJVꫴ���R�0d�T���-�Ñ°���GI��,�۴����s;�nT��އ�wx_l_�y-�zm�t)V\�C $c�-w<˖(�ͫ}w`�I�����y������p+�g]&`;X���J�U�M���AQ�8���771��:�"c���mE��*Q��ZDf���O��ulX�Y����4$����r�j��O���:�nu�p�^����E	��ˎ���S���u�F����@��4�M˗�P:�v^6�;���/F�8VW2ᛪR�Wv���f��v�L�/`,�[2�iT9���[	�u܈�1CP��{`��d��m�qָ�ܔu��}z�w�R{��<.�L�պP=��U�o�W`�\��*�ۜa���7�OLi�d!n���DP|j�XS��[���Y��'$����,W:�29��Z�Sa{���fB�eso)�O;��4V�45�z�e^�dh�|�~U��T�%m�>�"�ٟ�fC)�(�%6z�I."(9��P���N�۹V�k��҇KA"�r�*Zi����I������P'�4����ɏl��az�6������K��,���Ҭ�����N�g,��FF4�*\�VXH��1�F�o(p�z���1��:�miM��L�h����������٩�,�W \4����m��f�y��=�h�ݓzM9��0�>y�x�˶�6�2��w[i��۷`�)p�[�9���ob#u�n�nwl�]��޸������g�wOaiyF�V6��o=s��î���oF��v'�lB'���ր�W�9H�*���`�^�rv�[a�Л{&���cY�j�$�����ћ�.t�e���.����3ۉ�=��)��&gӇ����Nv�H.]ϳ:�	sQ��;oi�=�\d��G�����n�ml@#ٱ�Ц���&c��*v;]U=�+t�<�ֻ`�{v4�q�+vy޻[s��<j�[p�we�l9݃�L���2��v�v:�s�2�K��0��P�7�9�}Q�w��)�f�H��%�+ŷ`��G>{n8��<�dW�Uu��.�ms�0���g*S�^7c�w`�tD��&mR���v�k��Ů��.ݼ=�A�]���f�O'Om��FԮ�AU��@
���6�z���u5;�ov���֨�,��K���z�i�n{2u�g��7CQ�=��n�Pv��v�.x�u-Qn����h�r��v]�j�:���ۢ�A�SkqZ+�.X�xW��]�}��3۞W:ٗ�8+����������٥�G{n/n�Y�W]�v�D���gvg����>dK�ҏ�^���x3����n�j��3����*��=k�����v���g���Z0���RDkq���mК���Ϋ,�c�%��s�{vy���ZX�֛*Wm���ӻL�\t�<*����1;u��M��OLۂ7h8���v�K��g�O�\C�]�kum�x��'nҼ�o[�nŶ�^�j�����;��4�y���:]:�����Nԝ�J��0u<�mv����lH���{)����3�x{`Ł��]n���<�� �[�k3�w�3����	����Fl�p�48�2��Վ]̶��d,n7��5�;0S�p�F��nZB6/��M��5����кW���ܲ�+a[�_nSfS<������e{�e��h���nي�sD�9D��㍛n[c����Am��A���8��GW�x1�kp��ֺ�m���J���]�o;q�]�⎶uI�r��Z:�����uf���[��q���M�!竳Z�Zfd]�����4s��5^8Nk��v��I;Y,�#��x���}ƣ�Kxv�"9T��0�Б.E�A��=7 `"
N�� ���sD����X�ϣ��]��f�DO(�0�j3W����Z��
��Z�u���p�Z�$#�!�y�i^�i�Dp(�.���\�j��1ħ�]�QG��$A_7��9M>�[�x��g�]�S�"�
ku��Z��x��-��%k���KH�q��yo9�����)����+�ۛ(d^M�EM0Ƹ�:�㎛#H�VF3�JI��Ts��9�u�ܱ��ij�Z�tN�%H��!>��c&(i&�/)�M��ｺ��%�B�<�u�'�M ���m�.��L�f���s��bb��/����ݒP�2��W��:`�sMhP׵�ze,Ὲ"�c�\�ke�CM�aT�"�B��b�ː_�zA�'�
6A�`,�����C�^�6��>��u�"�A1"^��Ѷ�,j�3����8���9u��&HͪU�wucj�%���c��a�Ou�[Bsf�F0rSQ튶�t[��fb�ޥv�/r��O'-�p@���ba���c:˂W.>�{�Y�Zf,�ƇI�a�5��e�Y�V�n}{�SLz|������@��poU[t��y]*�ݰ�(��hj�ݣ��`��\��g�sGY�laS�v������rŦ����{�N�^��(0��W���vԃ�md�xD�}ʣ�uKc�^0FOu@�	�M�Lgc`��%�wFПU�(�Q\�9-��؋�!��%���h�0�"@� ��fy�Q��
�q��j��z�mC1[�<��1�bb]��+��m2�E�(w�]�9pe��\����g7Fط���+;rQP�ky�Y�d�>xM��z=�
hY
��2oeR����>a��jZ�Y�+^O�������01���I�Ii����?+X-с��=w斸�k4�9bH-���v�ՠ�ƨ��'m���õ���� h"&��i��G���\��q[�YQ��\ƚ�i�Q����ttmT��
�;�mh}k�\�&]^'k�T�^������y��I�@��ϫY�Q}|ф�Y�(�vo����|��滈hW�%�W��YIƾ�q,Ջ��b��3($�N����\�\��5�
��e=��u2:-�Ŵ.��u},�;��W5���]y�q;���s�]�Z���X8�u�t�d�=�߳��zN0}�������!��;�}��U��V�f�Y1v��/h�45I��K�d��7�]�hsd�`=Cq�]��x�C��swV��y��m���zNt�-h��Tk�(��3�NIN�;��>�J�U�Os�q��t�{Q�x��[#4�c�y�ϭ��nA�3+���J�����˱<w�6J�ꕘ�g.�ۋA<>�f��Ss,;v�;��w3�}f���D����T�6����ָ�=��pY;3��z�78��WHt�1�y=�E��5��8.���̆ٳ۩�N���÷��f�'�a$V����!�#�Ws]1��{5��4�ח��}���:��O��v�Y����OQ�-}�sH���YFYk�͛����LU3��������^<贝7���
�˚�a��]󦩎I&mV\��mp.�=�/�P�!D��nlj�QW}�g��g&h��Z�����CD$�{7��Sݵ����s�k�u���D8vb���/ī�?q��e*����9���wVqnWp�3#,g��e�F��2;��fyb�����I�:o�_�6��mڎ��|�vqokf��՘�u�l辴zgJ$���;ñ�2�	�<���;�����}�c�|���tsl�	���b�����O��*.����9XzQS�-���o���Ɯ.��nZ�]�U`(US�.��5|ڳ�{�"33�^�]s< e{�n��3qã[<���+����-Ԉ��Z�\���K;â���u{��ח�x5���X��R�v�e/���5�͹m�u�Ne�1[��hI�;T
��-�=�cϦI�c���$Z�O&�뱘M�⃹�L1dR���Q�%��;�}c�<-ĲuO(�ͤ=�_ M���Q�jݶ����;,ϧ�c�
b�%�/�Mm��٭l�fė���̍��q��Rw�r���
ੋ$������a��I��~�h����Tu�T����;SȽ�i��ص���v��Ҙ��������f5d`$ffa�2��w�i��h
�~�뭟|��5������Qx'y����@���<-�rZ�����k(�f��G0�Ys�=fMO�6�˶#�`��"�5j�{�A}ݹ�9	C���%�=�u�4[������o�kq�G�Z*:ӛ����j�nv�e1���������qڽv�H�8�]���S�6-\v���@�ՙюK��µ���8%1��(��msq��-���g�FT98��nS`��8GSȯZ����p�x^D��ڰcԨ���q�B�Sێ�4n�u�ayz��t�%1��spsi�3�)�g��8t�*v�6�<q�3�F�l��5^6�n���piuøAr	�U��Q��r��Ѵv�v�K�Gc��#g���s5��~�ERM�}:��X>'�~�.q��h&�{��UI�$�s��+���w�;�c/���WDn��tUJ��sK�nUL2{޾�~�����r�LL^t[Vk�F�klN!�L-�]BJ���4k�(�v��;�k���--��[-3ˉ��T|�u��M���~��)��)�g�#@��w��L�<��k>�͕�K]���$* �	�Gcr2�o�+�{t��Uri�y��)���ſ3�:;G���5��.���<w�.�G*��-p�գ3�}s�S�Ν^�<�ecg*0�|TYMD�T���a�o�[K=�l�g5�):�}���Q�̞L2�lr:��vL#&�GM�o6�4�=\�t�=���wi��C4u�v��A(����k�?[P��]�:�o��tծ��Q���h���Ʈ8����x��M�v��K�"M3��.�n�*������;_˴�A"m��T�Ajӵ�mw3`F/L���,]2UM�yP`�TV�e,-k�n�:�v���������:N;L�ӓ>�w����K�oS��c����s>_L"��s$��ok�5����Ic�;��*܌�_2�m�ڹ��6���C�z�)��r��O3�`u��i�j�6��c��W)����7/�ty��'`�3;��C����Wi�b�"u��ޛ�n�y��w=pz���^�������w�iC��y��D��I���t��V�V��h��OhhX]����P/3���`�u�(Ǯ3�m�Ϸ��=��w���%J&�n�"��D�Y9�>����=}��ή]�n�����c��vǩ��啈�Uʷ�z��y���W]�yn�m���+_*�lj��G��caƯ1=�����{��j+��r�T�'b���G=b7�Yj{�����-�o9e�'��s��:��ϐ_<���Y~s�r�3\U��w�UD�~�Ƴ[)�d�P:�p�ڴ��s��_g|\V�Լ$j|�����7��8L�b-�jg�$X��k��j��@㿖��G	�u�v����쏛�z�P�f�I#ׄq����h΢��~+�ݸ��k똆!�W9�ngm�i7e���bB�r���xXٛ(Y�ju,v+i��̱YPӓ�f�������bs<���/H�sxd�Q�<���c��B�iO¶��zB*�erW��6cyY)�wՄ*!f*�]�YA�kxw��ʪ�˵7���ޱ�Bo$Սi���T+�t�z�G��H�qTƥ�H8��ws�Y�^��2��#ٶ�kG/\\6Z8�p]�.�$ή��c6y�Ys�r��k�8�k!Ȍv��S˫�H�9֣]9��h������)ڛ���!;;"�t����y{���}MWt�\�Jz��cm�����y����}g��n��h�[<��a�lq��k[DN�t����b�I�ߤf�tK����
%�s��)=�2X�c�Dl_y���k:�2(��_����O�d��x��j���9S�[%c��f+�O��̓�gd���ftË�B���绶��F�Ǝ:��Ʀ���Jv��p����-�)��C��]ø*��#7�ոi��*U\�|��&-�]�9R�{��Ґ�&{����0����\~>�
��>��z�v}���WLU�M3<q��앵ܭ�`|s�[�f:�����b�W\�0*P}��,q�(�Vг���7g�l���4��yuջ`R(�#U�%��{��Md�}��sX6��=*�h�"c�yj�����c�g�����|�9�Mj�ޛjRF����"+_']�z#0��"zXqǂ�E�Z���8�6��۷j��n�a�N�֗������)^,�	�c�yD7���k���Iֈ|g�;o���"ݱ�i����/���!�y�Zȝm�8�)=ou�,��q�Q,���%��]���hď�������tQ�go*��޼�P�iY�5`S���}
�i�4�<��F�a��p�����oz�b������w�&��L�O�;[�[Yd4��X#�[��_�:����D���l���=;Y�}n��d��v�\r��&�bX�h�S��dak���4�݉
��]KTľ��I]��"L����t���ӛM��2��?��T�m�gw<㭚�jz3>�/o'�������cб���mY��z��3�q�e��ׁg�v6R���y�&xŒ'�i�]j#nmI�61��v�M�i�k<�h���Qb[O��s��c���wCÚ"Le6��7\�"+qV�n�m�uΙKs�e7=Cu�ś�ls�mZ�ۢ�.Ξ�.�N�h���v��[�L������n6���뙍�M՞;4�Q�8#[���Ŵ�l�Ԫ�ڪ|��E-�8B��sƞ&�F�6���q-��1]�f�}Q�0����l]��E	/��=��w��OI��;�U�mYm�*;MewO��,�h�n�WNd��6���q�Q�����ڝ}��ʔ&��b��c!�N��u֏RJR���W���)���s��Ѡ�EF�̥xֶ��T�����W<YF4Z#�w�����0���X��wdgqz�/H����c�_+���b�o!�v�������N�B�Ѯy�S�~������Yƫ>��vƁ������ܮ�qߖj��+�w��I��!��4K�����B~�w��R��6{:n���ƹQz=��ZPfe
W�j�ck��7=;�+<g$lq�=�]��=�َ��p�E�c��E��y�s�mNb����Cj�z6���u���Ls��0������x!�H�ʕ���8*S�0���ȥ�V�cwr�dm�sg��N.���7h�P�9<5�S���hQ�&���iG^S]�(긎�O��hb��ڹK���-fR�2�!��.���oh�^�[���т�x�J�>h��]�$Y�TRD>f�����Q�X1�-*%�e��}����<Pd��[q����_�G
��o��J$�ԷD��m�j";z\\�ʜ�7<]홞CC��ӵ7-��I�z����\���kK�R��[Rmmw�ݵZ�$�[΢.��>BC�[�&��θ��չ�����kC��@ԕ�S�K-",�r[�sL�>���v��j6�o�DX��j��%���ݫ��ξ�[�D�������c8 �~襭��{gkp���v��y����\�
�%;k��{=x�P�ڭ
씮Z�=�g���;��s�#`ޖ��8b�uWz��Tu����v��S�\�-w[�xc�wL����9L��6�����gt�ؙR�m��C�Ti:�Lܮ��͆k��fK���.nk�o���u�4�#��j�Y�t-"m]�7�{��Mq�=t���(�<Z޷�ۜ���bM��mQ'` 絖#5u[�Mu�b�g�g�"�B�&\.���Er;+�T����7]���t��ˡ�����;"v�Ͱ�d�T����5]�&�,{��a��d�T���� w ���VbY���z���C.�Q�9v�̬�
S ��U�ܠ�UK�����雴�i�$��"���zTUܠûA�R��jY���˄�˔4�Aպ ��9����Jd,oU�F
�H^Ҿ\a�oZf��W��b�cĕd��)��ԛ[�c�Bs77��/�U+vv�����m[��m������ꭾAm��.@�k:���l爞;���X�{qb��.����vMVȓ�l"�Y�[w�i���v���6Ni�.�'Q�����d��b����&e����fKZv�iٺ�Q�r�R��uѮ��N֊�����$,	��Bb�@:�Қ�vm:%V�`��mNY{���$��
}B���8� ��{�ˉZ�jL�+����t���J�t�e<��6�K�: /\��niw]{!1�ݜiw�*���I}��9	�VӢ�n�,D�]�-��f��\0P�\�����W�Д���P����%�[�.���Kᝫ���Z�I���,��ֻ�2���a޼2�	R�4m�����y�c�|�������墂h�\����]���ҏ	��(ӻ����6]�����ܦT��"}Ox� Uްo��֩-�Xr�<៿���_w�.�����ٺ�f)P`��)�e�6�<4�5{���to�������9_���50�{������/^
�L�h�gj@�e�4v��\���xc&`�3ѡy�}3%�(������V�WS���kν����քr����E�޴8�N��gy@��[��i�ZYu&Κ�(�M�nv�2�ۆ;�7køa�;^��ulq� r�ckb����N��e���)5���Φ}%Dꮈ��FM���X%���+{/��.=M6.�݊�7���FE�^��*{�6�/����F�d� ��k�~��t���ً�O=F�&���ٙp�_��5�4���f���-�Ήo@<�hI���2��7`���ꣴ�	3�������m�K**����[v+ʦk��˨��VbV�T{�ef2����9������9�o��r%�]���5�w�gF[��[u�7U�-�|����ߓs\�*��:�e\��%��*d<r��)8�Mr���T<V��ucF�9۽[�T뵧(%ztr�!�!��הT��v��w��W�?<���l�|1/��l��h�Skz�B㳯�;ߧ��9��
�8%�����47q{g�\�+�����
$n�u�I6�<e�֊yD�:�.�z�������?j����m��]\GRץ�[�\c��:�G�/K��~�o�T�G���<&f����iv�.}�����hvMY���q3��Z�u�:wf���J�[WO^m�:�W�������<���*z9�rN��a�~׌�g��ִf��{�;Wb1��H��Ն�����v�Y���W���o:��}6c�jҬwȱ[u��:�Yh�"x�s��R�ˉ�������˚OoЏJ�V������,��%t�L���zg�K,ͮ+��r��.����r�ς����.���ke�\�́"S��H��fg|�k�[���}w<һ�$v��7'We;���Ʒ_;i�Z� l���~~��KF��r��Ы4vq�X��R] u΋�DA�)�s:���r�g U#�]�wS��v�Wm��W���<+��+7Qf����j�ѥJ�%�^­Uu�>���y�λ:���[��kQ/F��{I��s��ڲ�[�&V�olN�7k�����g��r:::��ץP�9��)vye����Wn������t ��q�nu����홉���<�q�nUF*�v����9�g�(�3��N�ݧ\�]����'�gv0�W)ێŦ����\�]\��mI���:{�t��]��d�.����=���ZeT�tFg�Ɔñ�X�H;��0-�.�v�����8HE�ϡ����VǊ%^�}�N7̞8��o\?z�_���wT�.��A2w+^sq�j��)d�o��7V���{ّ�yf�o=OB��	��c6��d���yn��Vf�����Z	�,ԭnB���֌���f+<���Z;K-�ed�A���{˦
�F��b�Ѳ�yaݫ&ś�
���ҟ�!�e�
5SS�|���U�vY/-��鵝boKUUY�9M&Fـ�v7rۣu<Ǟ�p?�|�����i��.}���~�W}�/]��/1Qὑ�¦9\r��[�8��Ƿ����۵�J�A/�b!�ܰU�{�C��������Z�=Of��U��]��noK-i�"TɼK�u�3�n��;�����l�W��nz`��ܱ���e��r(�������^�^2׶��1٪�?os^e�Ì2���.mi�i�Y�9T�G8Ƞ��q�f�gwg�;2N�P��gOO5�ݦ3ۍ����"�+^�];J��w.����*IX
��79n!q](՝�.�7*[ۛ{R������N���F�����<�ݦ;5�}�F��uGJ,�s}�c�wM���nE~��)%�W;��*s�f���3e�k�2ߞ��{��;�}��^����c�wZ�uL�b�l�E�7��+>D�Jһ��UX7c+ޙ���+�\��Ҙ�R��Y9F{���n�
�ꋕf؍糽7C22"U�KXk3�c�$��ڭ��%��[ke�/�3�Lp�V�J��h�������[�}�t�������b���ɓ8?@h}�3Koo������/�s��6��{b��:�ݭ=���y��m��uu��ѻ����q�҇9:�8���w-A�*�Aަ%�������w�5��ʯ��X�ֵX���Zv|� G�@J�@[M�y����T�Я�C���`&,��k�k]�]��O��$Ҙ����݆Wsh�v���cz$obj��Gdn��J�f�,au�v��V�cGd�4�2���Z荗���{�7OBΫ�X��cܑ�D���1=\���2͉�ǥ�4".���MU���,k/-���l�e��U3K;�)ϟkmq���T�?8g%�N�ڴ�U������}㕭r9*U:}���~�Qv֡t
�y�jލ]�8���z��t�pD��Q��q�%7t�WO�����8W����S��dc��t;���Yt}�D��\d�;њ�������?x�\�e�
5Z����q���v�4v�[N-A�Nxɧ�묉p�L3�r����G8��Q*i�4S��W:���fR����Kqw��v����ŏ�c�b�{l�T�grY�g��bī�y���U:����A�ړVk�[�*C�ɓ
�EC/��/�,1�S)���K��}]����3I%����Kf9���W;u�.b���ۮUo`��OLΝ���xlӓ7yt�����W	��hnA �8�`���C�eQYs�/��V���ST�?�1W&����nk�毽'����������G���P�

��]��V����>���&�Օ�r���T�&"�/W�0@7۔V�,��,;&
�&���_��A��ⴏPU�G���4TYm���=�8�s��'��4ˤ�=sd۶@�}�[��׳;���4|���|������jx��2+o�ԙ.|X�q���v1�͍����y�d������W���Bht���u���d���8����r���mV�<��\Di��^�ڻ���;e�{ii�2�Ս{��C�8k^]�$ځIzpW��Z5$��ӟ��2˵F�WON�vӦR皅���l�,X����,�����MɉE&b�j����V�?j�&&�M�~�r��S�+i��wMvd����etu	<Sf�����d�Tt%���w�X��m��e�I�]�������Sx�����G	ojo�޼+h��Z�O��AÉ�=�w&���H�ʬr�౽o8�w�_y��ȏE�u�g�\��kq�out�f�c�Ъ�3�3<��_�lD�I�F�+j��GZ��O�领R�����v�kk��q/�w�ed�^g�B�ޣ����3S}j+Hڵb�?�F�3�8� �l�WWm���Y*w2uO\㎺�����ނI��d�����O�\� �0���.��1��È�ʱ��.�8��5�f��j��о��;�9��.�W��wHM7=ki�B�=��fx���!�T�Sq�Ƴ��<�D�0�3��x*��^6���v�����ɺ��N<\�c��חc�V�X�͆�l�p[��um˺M�����\{��&���Ɲ$�d룲�pݷ@�s75#��v.��tZ�nq�a����UX�kW(��-eU�õŏ<��B��;�]���w4-{>��X�n�L�no_lE{�~�׹ւnnk^�.���=5ܧ/q�y⸹WXܣ�y{�2ێDx��eh*�٥M#j��,�c�_"`�<�/�o�yI�mf�H����(�7}Z^Kz���}��:�6�5�����$�:Qk��;����k�}��i�:�|kb��y��W�6��y�2�9=�lff���kV4��Gw�	�����p�5de�|�=z����k-�Gk�ˑ͖YLfțq�3jyU�nqϖ�r(%m�>�d���l�4T�<K�ƹ(8�,��Ov��Ob�Q8��\Z]u%N[K��D+����w]�F�.���m�"pt3r�P���o,}�H4�)m����ew*9"��vI�Iݙ�L�Ֆ���mW)��۷=W��~A��U�n��3�y�ۍ\�F�EZj�-��#���$�\I;U���Vk�,�5�r�^�oGv&���y��[��n�J7������o�`�~�9y��j6'-eUʭ���'|����A_�k摭b��I8u�VT�Ww6�-���
X�5<�}�]�=�n��Fұi]�>;=��.\�����I{A��#�琑�q�|n��k8����
�
�eKf|��5<���rp�o�'o�qW�Γ�,Kκ������/R�],{n�n���b�t�"�����Cy�h�;�*fY�.��p�Ob0k�r.|q�Wf۞�2�n��tW�/�PQ�+j4X��Io���d�m���n�ڥot�m�-�>װ�=ʎ�Sr5�0{��w��b�y�me��e�wb�b�nGS��W�]��Ŏ�����io������}˝�(���r퍳�6�D7K�uNa�J���^�z|�8���ש��2�T�e���[O���m�&�r�C�uUʢ�-e}D��s���5Nk9Y�+��q�ڀ�����m�l&�I�cؖհ⼻�7����@�8;]>�iZ��+�����/9uu.�7��ƒwQn��|�R�dY2g@�r�3��)��zwa���.��S�����U5˂��n^�;;'.��7(�&�Uu�C��f	×H�E�������e]��E�
,;q�?kr������
�n<�TG(i�f;��y��]�m�gv��,n����|r���$�����u��v��������ܘiܺ�m��+�]�Ze�iо�.H#o/��C�����S#P|�v�������XB^�y붰�-�Xw�o�����)
�6oL���z9O	h�@; AzggǾg���5�ă};�3�uuN�C��򚅪�;�a�L+�L�ֹj���g{�g�3 ��G;Qn��8�gDw�g9�������.�-��-�g�bN�6�.�9{TUX-��W�4�,��ա|_��E��g�P�����B���\�O1���qoh�.�yXz�;$�Wd�XS�����#��Yj�h��o��ҵ���;�o��%tX|�%Ξ�����m�����D�<g�΂I��$�ܙ��r_W�K��}E?5f��>����
�.0j����.����lT�������~л��'�_���X֩��p�����;��s��'T�6�\�ѯ-i�.k�h]>f)&H�N�8NY;��>���ןR��L� �wT^i�����Z�XZ�+h���m���Lͽ�>N�ʷm���#�C�6�C�y/�w9�M_��(/�8.��tZgr����lf�B^��!�of��^3ɥ���G]�$�����AlT~����\��2y}f����^�g}�����Iλ�J��c�B���f�p�wt�g	���z3��1�]�f4r�䮷��74Ax�A\����ג�����C�m�b��xS}��55u�fNK�8.�ٜ�gu8r��z9�r�<��|f+���_���5q�xL�Y@�޽�4T���T����w^n|�Ai��V�tm��V�J*��>����1�A�0���� �(9�b��mnМWWen�����'��խk9DP%*C�Vp�dÙ��~��L�-���b��LZ�
��:<�M-<���zw?=ٻ6��b9Y��4�k�A�@]p���*��&�vMNIbg봹fSY���6��$#y\)] ��^��i��j�_^Tx��G�n�R|���e��m쾡FFv�0t��ˌ|�c�3�3z���L.g4Mɫ������ÝT7t����۷4,�4�"`]c��ԼZ�7�aJڃ}3gf+�iY�7@@\�z�w;�c1�L��K6�S�v[� t���=�]�{�)��u�U(f5�^�+�K�։��D���K#�8j돜]�f��M�|�i�Ҕ���ʄ��Zq%Io2�²"3[�.�r4G�x���P��>�U���-�I�'6S�����qX���)��v:�n{���%ֺ�t����M!ǵ��m,�yaw�m-'���m8�}��m�`ãk�Q�dE��x��h����{��:��*+�H����X�Xɋ�xI��׋��<]�ۼf�"�;ՙ��^n�ʒ��(Wbl������wA�C"�e�g�_G��Hkm��ӣ��`�
�yW�0tV�����U9]cwC���E��ڇV�9�-Q�5V�sd�����x8�S��.t0p:�d
�K$��1PJSi�-�ͺ�W��ԝ�/�:������@ڥ�*��UILu�ؐm�� Uq�AU܍�4�-���q���n[���;Zmm�v��Ӆ�nKnj��d�t,@����R�J�'�*r��r�[m�9ݥv��c&�,h\s^��X�!��!���ms��мݗW^�nۓ)N�T[�:ڶe:'M�U���n1�Nz僴] o/m��<�z��.u���N9���{�_1/Et���3��5�]��{ ��'��N��Wj\s�ܒ�;԰��^�A���/l!�=ƍqή�VX#\�u��àd��a;AN�V͠����n��+��΂��krխ��V��cJ�ls�Up7���w^�q��x㔹�;v�r�ͼ�:*Kp�ɼۮ�)�"{�Z�`�64[Bm����9-�c��U9z۫�kr�Ǟ�`�u1�;8{g���$+�c&�xX�l�ƂNdu(����N;�mr�>K�r�-�/;�nt�^�}I���qv3�@a��^'�갥`jn��l�M���w��d�ً]����/@\F0W2�g[d�s��i��i��e�n���dv�@x���ۑ�۲�5�����M��/(�<���X˜�s�F[&(S=s�۶5��uu��:m>k��ݸ�n������ƽ���EhR���:r<ܭܝ�<m 1�)v�F�(��5#�mr��;��d�ǩ�;v޷b�5u�l�G]�y�bYSq�j��q��*XP^(ն#+ŃLv��+�.�F�����T�r�%����OP�b��̎�p+ҌP��ۭ=q3D
4�Jه��c�۬6CN�nLBv����=e��q��;qѺs�Ţ�kX��@k�� �6-�'s�C�r]��y2J�8�uk��\�3��r϶^���A���j��v�����ۯ<M=���#�K�r#�4@ڤ�8Z�@>��(vm�Ď��{b�3#�vQ�:1�1G�c�g�3���;�u۩�om��у8�gn� R1��v��C�-�'FF�v��g��u��c��t��[�����	n��%$^)Z��ml�1�#���}N��r=�R���#f�,d�%�-�7�<i��;�6�m��/m�Hx�^6Ӭ��G)Ԏې���g.Yv���V����I����!��[��@5q���ϛ���[<�����n�q���6흭�Z�B�A[�*�B�Et�WD�����V�ϯ:��l^��4��Wy�n1a<>���EBuֻc���Ѻ��r��Rb����v�m(W��%z��Ρ�
3�Ny��c�̉Ӹvwv�,=�ы{3r��͙���e��WR�vm=#f�w�t���jwΦ~=��F�&�[ˇ�ær��R�;9�pDg<VԂ�g�f�j���=��]�ԇf���u��e\U�Oa��.���1�:��d��l��x|;�L����C�J�f�w����n=3�����]X��F,�ث�0*��\K��3�/V2�6�����σ�`yK�+�=ܞ3�ͳ�ƨ�U*��zM�����|η�K�s��f��b�(�+c�r;Z��	�r�y[]\Bl�mG��y�B�����}jD�bsfx�立k�N镼�]u9�ڸ ̍=�߉[� �{ <���6I1i:.���𖡹�5�W�e�',n��|ܾ���]�}��(�)�X{�]�fl���a��,�oV쫘4ER�Mı�Mb���`36��>�zՐ���U�Wj�c�*�5K~�|]e%)�r���$Q�Q�S{)�z�٭ڀ�-���SEvgWb�H�_���}�La��m�]	��X{s�����aXQǡ�XNa���tc�W"�ԙQ�k�����׳e�b��o ]H\; ���s�];��<�Y)d�B��-�y��#����̛��˾������ә��+�_L�Sk:���~��wι�n�]��3�I]� 61�w���x����;M����sk�U���w���gԳ�5�{�`W���w3Y[,5���r��0,,���}>�}:��yܽ�����;��8񞊥$�*N,v����
2:���~�c�Ulz���Z㖒'��c�r]mm�\k�Q�{1s���q�C��E5"��ңJ�+D�J�z���ޞ���x��}�,�ӃM<���߆�M�<B��l��s�͓t�e
�S.�s�嘺�̋�L�כּέ�F�j{N�;���&uER���o<���W*�l�e��y��K}Y�.�}��]����z�t�-���i+B�Vf�cjo�kｐ�a�nm�yq�7��¼��K��-Fk���nD+��9�jֺ|r�I�nfP�Ġ�i���r�k�/s�iHٹ�ҷr�o���g��t�����A�~�^L蚻�k�� �q��%t���d9��xgv��wɛ���Wi��������TC�B�m��O�y�V��em��s�k�N��E�I-7�k|3����=�	S���쭻�9��8c{ �;�/{����c��G/��k=ES7_Z�;���h7%�P�(�$d�N��������m�٧��
�<���K��ڶ�Lܱ-�3��#�t%���j���Y���|�I�f�s��l��� �ã4:��Q���8D���E+���uڥ��߸���>����td�gc�Օ�6���ɮ�M⮮�`j�dnrx�C?s.�ݛz��u�Ubn�%��9��ċ3;��z�6�cH��ʹ��Z;�������=�7Qq�[NK��@��a˼�k���|Β-YG���^���:�9��ݰmخ6�q���}-%a�� ���i���be�w�Gq����?�؝u+�1m5�f�������iu��uj���đ)RO�Ʒn;ዾ����x��&�Aw�5��T�ݲ�{��3߾�5��}���O��,�Ee���=��3�G���D�'q�h߹1-�����F�$QU*l�v;�h�T�M�\m�p�Vi��7��'��f>�a�^���	9LK��fwn�r�4�v~Ñ���sT�jyUlc��O/5������������Z�Zx=�[�����w��d�vNȷ�g�B�9ޘ�Yb���'FtY����[�}�BC�����W<��]r���!dNT�,V)�5;��Y�0N�2wh�h{-��}&�h]��LU���7S���_6�]k�2���Ad��s&�^��I)�,��s���ú����q����4,���_���%��A�ZS�4�>�
�}���G�%�g���\�NYZac�Ϸ9�c罽���8/������;|vo�C��\瞋O�M5��S4m���W��(q���`�]3޼�����@�뇸�ۻP�\���F�ll�"��އm�z��`�K�v�ꊧ������x�����LR6�"��i�f��Y«Rd��i�wgp�\�ul<��m�����=;��;2q]���sї5���G]z�m��ݵ�XxX��md�\)�k�u��GV�؝�s��yeݔ�Վ�������n�nn�t�,�n�l���<�VVv��SV̙���7W�w
�����I׭�6n�ݲT��"�DlP�,�p�=�mY훒�s����|���2'��s�m��E�;`��nѸ �k�lHb�*1ur��B8{g;�ϓ Q!�0,C��_usOD�;�ʡ�b)T��;�t���gyQO��S�ٷs���Ӿ�����m])`�+F�#e�Ձ%:���張�w)�2w"�F���+��+~�����i�Of,h�W"D���}μ��˼ �tE�n�	��`����H�{S`b>_/�"����z�U��j-��B�N���m�Q��yF��vjYjhrK9^�~{���:���4~����Ls���k�m���w(�X�ꛄ��������SM&$�L?x��Eu�b����oj=�o9�g�D5TN�7�n�-�x��ο4,�Ȑ�oT����K��q�Q�4}�]v�\M�9�y���i����2+�[��z6x�0`��\����k��f���_����ھ��� ���G�ҭ��t܈�YL}۽����o������΂蓘p#fұi]���[���i��_�N�񑛵@��~;��n��Bt�g�%� �Ks���ʬ;�mf�DU�X����[���//6YD���%�7eS"�(��"�E'��u��XOHA�zw��q%ޡ.���7D��TNI�"ŝ�u�&�ib���_);�������j�L-VY�n�`��l憥�k��$�p��-e��;����V�)��o.�=���Y����ӳjmE����L:ߖ'����jz�s�w�9?(&�/cz"�T�=r���8.fN;��uq3�������ݼa���ds}y+w�aGq��K��P�\&_�u��k���s�Xym)Ńa9�,\&��mYOv�96�l�;9!�{>��u
\��{�k���0���j��3Q�kd^��,��ɜA�FV���vm:����Mw�`�����ll�l��*�p�b���)�ݯ�bqS�t��ظ���!�_���e-jN�w&��!�����]Y~��@�!�4=�NQ>H#jңv��J��X���_tø�Ѫ{��wv���j��@g$sS��E0��7��rV^S�23e7ʶ&=����GYJ2� �#����Ûg��@�2���EGlO�V����f���;�<��j��amF8���b��9`�AN��	ŋL�޾�%U�;�T������B[�{�Y����G���ɧg���>N-jʕ��"�tvg%��݂.�;&u�ۧn�d7n_-�ӗQXQ|��g�WV�f�V��ӣ�̦�-�n�V^��^�wL|�ӫɊx0�����?�ݻ7p2��ˣ���iϝ���fҘ�/���-��V[E+U�I_^�Xs��]h�np#�o:V��v%���ט���7�����~e����䨛͎԰�!�0!�(�Gv!��\�L�U���YO됣\.�X�h���׶��=�Y���v���q=����&�PE]�;l�f`<�����y�|e�·�����Uøc̵e���cks/7.��lA����^�`Gj�WT���<�6m��l޷b�z�Syݵ���2w��e��QW-ì�Z���?R�����j�ccTBg�ւ�ʷNZ(P�v���4b
v��czu�z;�o.��y��e��ήQ�|�Ա�.�1��O@X�B�"V��J�5_׹�����`�2���Pa���C���v�aS�Үm�˶O}��ũD��wt���W�Gkq���Z�p�˶��n����BCg�jWk��Q����r�[*��b������.�&u7�k��My�}�,c&�KOl�-�*�Iu)��ܝ��Ҳ�r+��Z1`��;�N�\("������	�.���ps�N�l�L*��6�wM��J3k*��)��X�GQi���c{����&���vwW[��#��)��C^t��,>7M{D��������d}Z�i�����R�����wWh7�w��u�����0A�q�]J%�����S�����6��udKgD*���#��rl��$���hw���}�	�Oi8��v�E�u��c���>oS���[S_kS��|2!��uwz�_a�5��/,cy2D�6�4X�E[�ǪS̳��"�g@�+���e��Q9z�s�dow[RL[Kic�H�R�%R�V�X��6��'[v��nt���{a���g<�h��L<ʽs��ln���l�=upv��;Th���a�V8��i�nʵ�>����Kv�\tn�ӷc"��q����v!��<�vz_v��w:���Ř.����u��������5�u�oX�{gx�������:3F�ܛA #����x��h�Xx{v������{�����e�9費sK!�|1����Z}T���_����d��j~~o8�����nl�m��b��P[��W���[��53��}ë���]H�Rx4qv!��r�����������W��*��t&�m�fu�`\�#z�����w�܂���!C����9�T8������L�k�y��=�t��a��bl-}�R���}��ϊusj�ެg��F�ބ0WU�F��'\V�17o9�S}���m�@(����cr�l��XZMھ|�u��v:�1��ٜ͖y�s4��������<��p����;E�:�^X�M�Т�h�ւ�ENOR���zj�����GfS�5�ԭ^+�8�iq\%�e�N23A#`XX����TA�</u��3��9:�]���.�.��/-�p�17��^���ɛ݌ �1��U���{�����ɞ7
�W{w�N���w�5֌!���N����Mn������f����Q���5ʧ%+���Dd��Ϳ��V��fяɺV�L�|���F�b��㨅^r��8�{)�+VNX����[�j��ǆ�����ح���H��T܅�m�K�7ngC�ES����K� մ-��l{��a����uͽL�l���Yƨə�b�?c�c�f���ud��}�����}J����l#e+.R��=��5������G���^�+��VJ��ӽќw�N��I��������%�1t*�����.��3�)˦��,n�<��]/Y��]���˷F+��ϰ�$�WJB��(��sg6����ږ	���*L�j�QY�㞍���ȯ0y�ו۳����Pmunz2��=mҡ�VЫ�@4텃r�����:�',��΍R}�͹Po&޶�s9	CP�G&z%WZ��Y9�N�Xb5����W,QX�m�qw��!����S<J��s{oi�9�b�[Nˮ��q��W*�÷cp��T&o(tR�흞u�X�ڥ���L��>O{�I����S*�Q<>�/�N�����қ�� �ǁqu�cl�6�T.0��	ߣ��HV�Z6��q�Ǌ�-=�S+�,��kW��Q��F��P�I�\Shme
�q���5�vGk��g쮝�͑�Б܁��ښ�c��X'V���@��J�6��:-o�|�*{��=�2�1(�8B�����N���,��ru�O�Ai��m��H��3��÷ts^��&�X�8Yc�2Hʴ5�<��YqZ�n��+nE�1��j�p�[m
흵�F�ֆ ��ql=]]��م��d���v�x7&aQX�u�aN��7*$E� *�.cj�-D���F�*Z�=��-h������_0e
v�޺/�(�S�9���7V�	��9�c,�T͙	�+Q�F.��:P��i�<⬸e
Ӽ�qh���Skr#2�u�eIH��@anJ�k7����:m��%�\�ew�k�˦X��lꮋ7,���x��k�ɧ�T4��9�+5NB;<��O.�^�sP�Y��VEQ�Q�6�#[V��Ճ�%����{�rg-��?���
�uZ����4�|�^V��b�3\<q�7���i���ǛZX7+i�����n�Hٝ���BA�7[hQZ� ��Z+NnQs6��&���_�̶d���+���rSǏ(iLU��^�4�GQ�5��Oi�v��q��9..y�.���F�� s2�}J��9�|�v��`Ǘ�wFb)*.��j����«z��/~�����>g>��ʖ�Q�J9ަ{w��Ի<o�"鶹���¦����Y�����M^��+��%g��݈�utb���xһ�J�C'b�:g)������T�Y���ۼ�&_�p�3���/�C��������tT`�;}���3d�p��c�:��:�ʋ�J��"�h/:6�@��>q;e����A85�V�;��m�{p�W�-
WV)_�T.�%k���|_��q�M��]�'�{����e�T���|��S�kkZ�ƶ�rf��sV;Jݐ������9ڟGS�8đ�x����c�MuQ=w���da� ���g�f�:�S�Sָ]���'���T��%z�"K��3s�����Ϧd�_V]�ϣ�O�z�ݧ厳��s�D)Q!2V�\��o�̜�������;����\������\�46`F�S�,�w����6�z7�&/V��"v2���NJ��Fݝ�/y���j��8��Ջ�zt�Y�(,ޛ��j�0�옘*,n����]���KC&pK2dAv|��ޞ���R�����5�^ �sN�8힇jv��;<W�E"��WO�/{/L8v��{�\l�ݳ�=]��xG���n�8�;4h�8�м��A�Yu��ݥ
{�����ۆ3���X�wW]SC�9V;o<]�?E��AV(���雚P�Z��a��7�V�T�}QI,�|���[k���mm�}#S��i��ñ�n��Ds.7�I��m��c�b��l�u(���:�;]U�-α=���;�o~�еI驕m�i��vjr70��)��������P��m�Á.�����o%(Xn��ѱ���,��!6�=�}w�˟�/�~�.XU�݆_����_o���ٯE�b'����J�Y����!�\�g[g��:�aL�w-��E��ޜ��p`�Y�<�|b�S�o�0��|r�B��ߨ�7vG�9�jb�mb�G��h�;n���Oo���kˊ������Q����lL�;�z����}���8�Lv1s��N�(�G-�[Nw��ֆ�sgqU��;z�lnƌS� ��3;ֳܔYɳl��I=��r��ω�X<!{q�ngqμ�w'n�V�Y%-�H���۝��{�Sg$o݋ut�uxOTq�l㵻�IۣgzM�c��:w7q��;\kf �g�������T�v�s�u���s7�[�����9���.�sR��r������,�7d%d��Y�G6����箲h�g�l7B=�w=dA�����shyX�~��ܠ?��L��QV�c�'<+h׷�x	^����,��۶�X�p�̣�Lh��+�I@�];�	3���<�}�2�]gS���C��\@�h�_R�i�Mew��[�IpJʻ;D��k�6��ڞ^�����^�{�Z	�&�P�����#c��Z�S�:����ܺ��b��4D����Ge�����xpB�BY�krb֫"r��T���X��]-z}����6��*ۍ��ޝ��~�|�٭��|ݸ��u�A"[Ws6T�5�7�6��1�UevJYm��:s��ծ�"o=R�T���}�<��oFb>��>%�s�N�Hu��J��`���s�b{ʒ�j��6��DG" E�ës:l�ޕ����/�nܦ�m؄.��ww|��awM>��3�=�흸�[p?C���o�}6$�y��]�?�j˺��Goy�9g�.��ϯ
��_�y7[e���V>9��lF��ܼ�<U{�x�V'fA@J��4�!�39>[8�#]w���oZV�V"�xV�=����oE�c�����5��+=,�7n;.����}���9�wL�Q�[d����v����_�5�wr����2�e��EAja��d;nT7��o����--��U��g��Y�
�*r�,�~|�&��n�Q�p��FTl?�,,�~���4\��t�*�̻U)�dͰk��t��OȚ4U��+��͍�	�N�#�WT�c1��e��J���C��<����Zk9�O�eLgK�s⫦4c4[�%=>�Α.��.3�k�G�:({k�,tu)+���6y�qՄ�YZ���QXՊ�J�䍫%�q^��Ӡ�M5�P����7�o3�ԸI�F���=m���Ͼ^kd.���{�i:�$��Q�$�J������!o�z���-ޣ�<�2�z�����ն�ϗxk7D�����}p���1W��X�)51�� �Ɓ�'�I�h���F�����f��#yb]���?'fb_1S��� ��MxaU}�f�U�juͱ��wB�<��K<`��ָ�4�"�K�>Z��^��p�̫TE����-��:nL
�|�l��KU-�ݬ4����ɉ�袭�n�n�$����6��o�{�n�xu=-���ڢ+�܋��or��K3G;gk���4�1�><i�)��AY�Hm���yg����}��2'�;�
긶FuGKL����[�n�Y{�Ѯk&T�	�+��dtD�nG�(yK�޻���u�Rc�Ք�Y�na�8�ἾZp��6H��@u�^{9��o];�MϞ����)g���'7v�^Q��q�/ϖ*зS͚��/|�s�\t]���X��Wgw��?���ϮQ��<Cay��a�;���Y�]k�f��J���^@�tj�g5�MƱL�$&)ܹI�S	�n�Y��yd=�Mq͍�p;$ض-��9t�2+����/0��qq2#��'vwE$�C9`�3䌅{�����.$�l�[R�����T�m�v��ݤ��.�2����)*���L���s�ǰ.v�"�\�c-��]�kF�7�	��٢�\Z�L��8'��ڭ�j ��u6��=0'�9A^�ó.g��!U#DR��G%���e��1���[t��4ݝ�F��9�*Ld3�Sv��N�5f��X�E�ֱj.Z^1������M�oY##�&)%BU߭�j6�t��:ru{`.���M���x�xw����!�t���˳����x'u���d戊�չ|�=�o�~��9�ت�ww��s�Ԩd8�7圱x8WGU�9m��8�U��{��n�Y���	�o*2�z�\�s
ʼZ�{s2'���N�WS�WX��ߴ�\Y�/2.�'D�e�W}p�����
i?(�70k����s�9}���B�'N�侩�h���ڛ*�'�!pR�	S��׬n�[������^Z�޳��oWU=1���[��=F�a��_j�f�M=ĥ���=;<�:)���ݝF���������:0dT�=&�/�zx�Nf��gP����G17d�jv�M��x�K+�,��έׇ��*_�r���U���"Z\��J�jI���N��=N�w!f�~MҼ�*���n!2n��f��Z�cc���0c��6͚A�-X]�]%�{LYz�q�ur9bKC�n�:��FZ�z۵���_�����ƸEXl\g��r�t�V�;R.�[��ۂ�q��������mV�n7>S7]�F]������vz+Z�5���cX�S�kGV��,�ѭg�֩r��Wyn�Sm��O��[r��;4gPaL�d-�����-�u��`����ع�Zݳqآ�#Hx(����[6	H�Xw$gF,2\��6��ێ�1,��YIf���f{���v'�����t�=ܦ�Fn�d�\b�`����W�ʮ;|�#e���Œ������',�����s�uBz���ZxN-�*��r}����F9�mGSbȆ�����r�|	t�60F��Y#�\�&r����N����l��%X�������m��7����S�7۩��X��T�K�;�~�L��B�>*�K1��'zZ�W��g���9�N�j�uvO.��B�;Ԛ���uN�RM:Ǿ��Ou���OzP�T�C���Ib��%��5q���o��e�d�Aͣ�����O����/m^6hV��1�{y���#��)���Yb�t
7�]p��]���걬أ.�w	w-����v�/�J'աGlXuA��9\DN�{﹛��g�d^���9�]A�}˧�\��ܠ12�V�C��ˈ��Vp�و�T7�G!A�r��m�pcR,y�9�j�V�����Ȯ��h���r�9Y���r�غ������᥼��o���2���la[x�lh{e�{Edy�<�VD,OX�]�1�kq�S˃7�坹��ٙ+jnR���K��t���b��8/	�Q?��$~/�1.�O���
מTT?s�h6��R�z�Y�ћ�q�g;Ҟ�-��H��m���k�e���z�����/�d�q?Y4�Rk���|�wM�s�j?�癵��2���6��u�?|T�M�p8n��3����ەh���k��$~z����߰a[�쟾�a�Nug�.7�������ڏ��kG��s˝Ƌ�0��Cl��%t\��⺳x�繸Vv�����kk��n�lRW6;B��+~�Q�k�T��'��zc���k�2�Rb��]�>����;Y�6jz�������o'�w�fg��6A�fqH�l�v��4=)}H�>֌x�XWU+���!������cg��j��qsЭ���njj�!�;�b���HZjjf��7�/��{�g,>�7���e?�9��N�^�u����U��ݲ�:u�{u�2�]�ї/P<��]M4M's�%B�s5�n�У�K�'�M}dY�C��T�y���8w�n���YÀ�v�u��z�T���8=KU��r%+�9]�͙�sa^olVӓ��T�Z���Er�W�*���9	�Va �f���nh�f���yB5� ڵK�w�"��Ce��q�n�NYQ�Tb���v��n)co�:|G���n�Ҩ����,ӝ,��/��p�cϋ�!�M����Z�vYD��w.�)d���t����V��o39��v�������u��-:��dZ�m8��of��ob��n�,grRvI3���ӁԵN�^,�8M�6.�%������_�Qߧ��������r2�$�k�fr�$p�O�2m����,�xv�NZ�noy�gM`�D����E1�~����Q�0�F������;e/S2.�'M���z^j��D��T�-��i��dY�o*�5��х��&�$��9ͬ���}Y)��S�gZ�.�+x^��.d���Tg�����T
�n˗o�[��}3�'�X��4�TY�Gbd�k��苿�.�`
����'�h�d�p�3�r�ͷ��W,�۲��Bj{�%���=ڶ��۷]񜗉�kk��mQk���яY��F5�\Wq�xdY2(��ˌ&6���om:5��j����m����b��۵�D���'U�~���,$���`Mx!��d�������I0�y�"�<��F���>��;Iաj���fwŎ�:�����}����������ڬ.�6��	�0{;q۳�i�yT.�j#��]�Oy+,�b*9Gm���rj�.�Yս�^��;O��M�p�x�{���.��W^��y���}�x��eY���ty�R��cp������D�U�$ܻ���O �������Xa��󦖡���J�}�b�u6N23�|�u1�_�~�<?�Wh"B��Pr�j�m��o��Ň�s5s�h<E��~
%B{�-��#�ӽ$�N/��vS����$l:�?A1#~ջ��T���VU��%��5o��BW%��9^*7j����X��(p�l�Dvfv�و�y\����b�VX�c����f��gf�����Wȫ$�v���ʫ��ۅ�" ���w�JjS���6:��'���oP&��D�:_�*�Le-G!�=�4�7[}�v����Y�ŭ����ή1e�;b*��Ŕ�"n�>
]̙Ղh�]�6������7;�2]]5��:���mZ�{��k$�&��v֋���c���ō�8�NX�wA�$OV��[������(��+r���t�NM�y�Lt��X��\��YQk�y�h0P?e!D�D)�A>�(��]F�o^j�=4dtxNB�=�S3���V�i��-T�!��[�uw>��,��ְY�ѣ�p�Mj�|�b��)�z�[2�C��=ON
)T_�nTT��¥b�2Ên٫β��VKCX��ٻZk0�JT�Z�q�oC���0_E��*��ji1H����*�=�/"C��Η�.|p��nݦ#�)A���1Ï��N��\D�n�f��]��
3��zJa#ox���a-����%j�s!����E
�̵i��a������u�cJ�O.��aA�l�@(
�ά���!�5�r�G%>x���3���e���Q��.;\�U��&��OaG���mV=p�O6ͼ��wǎ+I#vAEJ�J�5H�l���[c$ce����L�R�;s�j:��rn'ŧNhKV�I�����4��UV��������V��-�jM[I��a�,h�����Ǧ���ŏb,�h|�+�W[��d��r�h��'.�mDs����5����쳶���u�g�+�Ӂ�^.Ԇ-S��r���h��K�ǵ�a��,ax7
��v����6�[��w^wd;X-�x��:�#��r<O�����>�'[R�j�sm�y�p.��n��v�ۣ�Զ7�g�a��IV����5�.yqZ'�����u��U��z4�N�����.��k����-�n�+����n1�#I�D�n��b`ƶ���m;s����X��z�ں�70/�odrm�]�Ѹs�cj��Xnf�%�����]�ı��pgy�I�.�rv�h�Z�	�6y��ヶ�۔�m]	7c��og�Ս��y�,Ob,r�E��6;m�'��#rݶ�W�Ɠnn[,v[\�c�ZH�治�H�nuv��ki��=��;�(�f�[��u���!�{c<����w��ɸ��ZE1�Q�9�`��jQŁR8׌t��ӹ��Î��:�5���=R��a�V�:�q������Y��9Xz_Z!�4J*����n ���ݬ���<��NP.�BjL��,D�{}�}�@;�ؘ�{ZCΙ���N^L� �`y ��cqRjxw��\=���-�J;8��)�W�5r���k�}>��vU�7�Г%-�๵�����ŝ�ݎU:��Z�7�:N6DDy�K�&�g#�:|���	׷���)*GO9�nM�s��{e���4�筺N�!A�v��6�m�:�r�(6��gs����\v��)��7n`!l�7A��͎y���l�}Y��댪L���;�W\�۝�͸�}9<�����N8E���sݣn�V{N��S��q�2R�⋾9�ݭ\|�zyƸ�vY�1k��.ต"9E�&���y;tkf�8�A,v��ۗh�\��w��� ��5GA;�tsI�7�M����7nyN��Kq9�W�On��x֌�8ݹ�67l�.��[G��8�X�/�^N�yge.Kq�;͵�]s�W=[�J�}[��3���=�EȤ:��N�"�@��J�&(���ݚ���::�y�'c��B�g�ۚ.;c�hs۷q��b��:��Ń6���[��﫶]�:�!A�g��ݸ���<khl���:3m� wm��yu���Ն����Eg�]�):��E�Є.�%J.�U�����c��f��ώe�;�A��Սw���Z[g\o4]}�|�����߹�q�w��8F;~vR�h}G�X�~���.�jG����<����}Qr��=v��4��uS!}czC��G�5�]�fy�b%v�%QWe�j�O��E'��8�"��owv�J�����^�v�+��Ak��I$��s���殯ݼү��݄v�UdU�mצ��Ԅ�R��z7vw�?R�h]��؏�ݱxC����U_����gX�3q��\sϦ=��f[@��ݲ����B���b��[	S0�f�(�ey�S��E�������-4��e�}�S�؆���؈����8f.Ń�f`��;#���>�GgV�c!����$��;z��<.{>��3wt̋�N�x�}x�k��g�t�v�4�]�Oc�ۚ&����S=\�A�9��M�=N�<�x�c���H������������G>����_��X��P�p�a�Z�'���PӝƏ]QFͻ��6S�h�g��_c� .)��rQ��(��v�.��23�w`�M}T���F��o��t5���ݎ�A�m�^�r"��n�����m�Zf4�����&��ڥ�k�~_t���4�}�1Nd=|6�s�;T�wf���ɬ�s^4{۪M&�Y"��p������u!����Ǜ��,XB�0��w4�f\)�綕o]W[�H���SQ۪�K<�B�~H�]ګ�v�g�%>k����.��n�Q�n���m�Er��l���yC�ig۹i<�����_YZς}[ϞvmoX�m
�J:ӨD�θ���Mw�b��ֺ�GYAey��n���D������nw�z]���kޛ��%�Sܢ�ݕ�7csUV\�Sd�{�KZ�F=3��7��OMet�J���c�i�[Ҷ䀭�E��{��?w���]��ahZxM�J���{M��Xe5��s�47J�;�P|j�SΊl�:^��D]@��&�+%�w��2�n|"�~����u&̬���q�C�<����*�m4�_$l�.���/��9չ�+�qtN�ZX�m�YL��Z����zs�Q�A�<���b��{��۴�z&/l�Lk��f���Ny�	�����F��:��g05�k�{3�����gwηTw~�l"{!�i�.�N#Y�:�g��҂z���+�tqfom��JP7y��2���I��t4+�Do��<�ѕ;z�m�=���i�����,U<��{P���t��[=v��C@�l$1x�S'	�d�+<PZ��:�{]�u��g��� \�n����Ӌ����to�o����g�إw�vh<8[��H�G�Fk���bV���!��ݹ���.�BuF溇Ep����8d����~��^�ކ�4o$٫�S�������([�-X�+��n��w��N��vV�v^;f���ael���9B[Lnra�u�?{�\<�ѩ��^��B}����k1CKUޘ�U#t���J��KHu�����v)N�Wwoj����?�4��^aב�������w��z$ﾛ΃r���[/�}�:
��mҹ�m�h�5�1(�]֕Қ�a��o�R#��_hW�u$$=��q���n��� 
E�$�Z��و��W��w_G��W��uZ��Id��2��g2o��r���pƲ�C:W)g�h7��9��ʼǹ^ދ�`YsT%��cn���|V�a���y�j��u��=6�<m�X{.oi�#�`�:�J���-�Uc�7}�=g^�.�ԛDU���B��}]�2�0��{��ky��-����Q��kf�=���1�C|d7x�wt̋���1�nq�;D�}��9o�{��f� �Ҭ�k�S���G��w�9՚�Y֯�]�o���n�G~�Ye{\�"ٌw�͑n��R���$,zvZ�,��)�K��~�y�;F!ُ[U����Ul��r��c��lc��*��m8�]n�Kt���d���)Y �W>��p�'��Pq{&[9��>�뛷��z���}��2&��6�5�%�#V(�v�|��\(|��������G����ϛGaK������bf�IE����8�g3ɩ�����ײ����ԖZÆD�uF�f9WA�6�
�
���.KT�dd�j�QyH	���2RCzܛroq9W�8䨣$�Y�-Sn��vA9Uȑ�%C��K���&�utc8�Х<��νr�-���p��:�=��%�.k�٣�t��Z��cV8�ᬧ;f��\��h�md�=����m���Ό�tk���n�2m玒��]��9��q��Ӊf��t��e����\c�R�]�6ܽ��}�`2s�X�,!�	�7r�;�r�G=��n�8�����9��k�N��۶{uΦ�Ll�f�=``W��"zSr<q��ڤ�����֩�GX��|T2��֮k�k�9��]��m�-���Q��|�~��6�s�,Ū{�%u���u�y��E��Mh���nB�u:��cnr;]�&�#���4[y�v�ξ�Q�q�٘oe�^��Z��6'�F�H��ZV���ʘX*�"M>�n=	��M���^&�ng�>;��I�z�|�V#,'��o7���z��M�[1
R)[�0�ж�/���S�~I��C������Y�y<�����-}o�eζ-��/�}�=1Ԟ����q�b�7lqj�d�M�v��zv�����h�{Cq9vT�s�2�s�u��<�-DZ3�\g�GE��yb�����诞V�֣O��u׳�����w��E -�Q�7k�μj�V�(4kn� ��V)`�)#���-|��qqO�Ƶ��o릛,tى��6w������WP�Lv��Fm�[�t��7\�����j�(��YQ�-�����%3��;2�D���{��]�p7�]O6<H�� ���NL5���fT]|[�Ƒ���%��@�G1n��4*
]���,GY�Gk�ՙ����8�P�m�0�?�m��=a�T�<�\I�P���3n���7$��i%Q��r��Wy9���oML��{�.E����PC`'i���ˮ�Q��7����bl�MwP+;�%�I)��g!+�oշee�4} >q��Qr��%=�B��	����c{^��k���P�z̧�����rf�Tg��N��fpΙ�9���]���y��x+�1z���1��X^Z��4ϵ��o��c3Ak�v���n^r7�&��4խ��ٵ������JA޻4���c������$�t�d�D3r���Ҡ����
7�a��u�)������g=�CxY�n�{zǞ�,ѭjm�,��X�� �]~���|�Q1Yלf������V«۫n�c���GuS�c��8Dd�w^m)C9PUd6��������f����ee�E�<��{���OK�xj���{�l(��<��fj鴅��k%�\,��ޡw�LN����P�S��N��{��!��6�OZ�Hl�z�߾��۵T�t\=�65�i�˕%!�Aٓ��;;�ӻ�8����ߺMlL�S�O ���w�'+n�\�9�Se�z�hv|��귯4]���YNĦ,��F�]�ܻN�Hoo��u�^��Z߸���iy7�V�ulErw�b��xx�{s���}�.��B4Rb�;$�٢�kH�]FO�c6mY������z�Gel�2�ڱEKoz���w������E��cUWSs�ZQMfqw\�n��%[�yì�}����ǹliT��[s;���@�5����%�vO/��7�;m�".ۛ2ZU
�y�hQ�f�(b6�9�������/a_vu�ˢ�޾P�S�IY�JF�Ѳ��S���Mm�ڥ�]z���t�K=^@�x4�z�f��GY��Ő6&��yM�y,h>��p���-�������}�����&Z�hE���H��W��_�)��N��߾=W�8!rJ߼� �ϒo1]�,����*��5�&M�`�u��� ��攲4�}!�/�������F��e�<B�:2�����XÔ�:mc�N ��]�`���[x�o=Z���򱦇Z��+MB��:�޼w����Pi������o�gsgmۡ�b�����rS'�ӯI����\��l����q��������{/+D�t�j1��ӳ�k���E�Pe�ϖ���_��Ւb[�t&<D]�eJ�[�c��9m����7�U�ja{�k�qP��7-�vY��z��i}���y� "5�:�Y<%�wV���<��8��u�(ou4m�׬*ܾ���Ԉ���c�K�cF�rV튖̝&g5NEj��f�_,�vV��h��V�뽬z��Ξ���?VklvF�֨����7_���=��,�Ki*��G/.����q.zk��ɸ�|�Y-O���[��L�=u`[�aS�}�*z�YlV�f#�d�}���'	eQ�*�������V +�gӗ@�c��&u�"�~�HWD6
�ُh4�{n��c�zR�W/j-	#�'��zn<�K=<���%;���d�l���):O< `�
�W��DT�^����=W�/P�c=����<Nq�'�p�E|����+cn��Dݸj��&���
�����h^���l`�qѷ�;v筺/^:�}�]vd���I�v���u��v9]�r8��i�ļ��>k�დ��h�t9hx{b�y�9�"]�N3t�*�e �۵��v�k���QW)nv��n��� (�.s��un��k���I�n�)oOn"�{{l��-�ó��+��0s���n�X8$Բ�\�S\�[�Fp[���;����Ż{�q	Ƈ���-̳��V��]�Y�:N��|~�u|����dI�L�SF;'���tt��d���;]�6��"ʵ�k.`��q�׭���1�U�=��+��Z�*��k�(SMK6�v�<^E�2��a�F�s�?]���0B91��|�$f�fj��RLY�F����� =�8v�P(;��xn[�c�O���c�.�\yAm����r������?j�}�y�g��?x��W�?o�B�X�{>#2[lP���VK^�]�Z:7+m
��v��v48���E9����c+g� �����)�;\�CM�����?���E]����x����ldu�Z���c��-�z�G$g(hn�yT��4z&w�_��n'�ù�1;uF[�(4�t�.�&�Ab�p�F�p�����@�g�;g���q}ŭ�X�HuO�
���O�[���{�g3Y߮Ra���2����[��C>��tv3d6^��K+���J!���L˃,�9� ������ۤ�+t����5��e��t�mu1ht�=+6*QL�VF=�"��]�,��H�3ҵ�Q�y1���7KA�V�F�\�]���;PQ��|xXݓB�Y~#�Pr����i=�r`�l�w���{.߱Ousf�y�x�"��5����P��*��k�J�j�����ٜ�(m@h@f���J��oġ�V3������h��SM�0�ɿ�$��:�=kvR�$�����pȻ[��@[ڭEJ�Şm�>��r��ɜ��'7e2i��v�c���eZ��Oo��,|��:쑪IQ�:�T�r��.m歬�oY�.Ȫ��'T꺢�+u��Nn��ްӑ�]q	�1�I7��&�z&�c�=��r�]	Th�6v3�t�i�4����,s�X.�X�v���\	��ո���Vǅ+QJ�1��o�y|�5�m�|tV3�l|��ƹ�h����έ�5�4<�3<��dլ0�tff����z��YxOM�Z�A_��K%xZ�z�h薶r'D��g
avh]֪%GtB�8��Lg�ɻݪ���Ѵc��n,~`��|�HOw/���d�D���N��#�}�n.�-�i�(�o'�Εy�����s��j����M���e�|f����C�QY:P� h}��^�w���d�0�1��ԥ��v��-�o)����-�Y�h�0�z1X0�.wl��:�M��9ӡ2i���+p$D����z�0��Ό���|���o�����\��>f���|)�B��������MkF�]Uø�r��t����f��=}A��s	>w���^���C��%U����'mn�ſ�dL�n��V��"�5��3Sqt0-ˀ�N �M�*Ӳ�;|�̃����3O={�*Q\�[|��C�ZPX���ð˥4]��D��n���̻�j�1`�������d1
�R6"��Ȼ����ͩ$�N&\��m]��2u��Z�92���\d0A�X�V�޾�W�L�}; ��(�)ִM�q
�ğ^�*��p�HP�t��G��Ƈ � ��	@ຼȻ7Y�=tjՊ4+�JA����WL�M��I�ԯ+1k��!�X�TQZ�R���gF��FʄZ���hU���γ��؇���)u:5Hp�U*�7"!]�
A�uu�(tY��nӧ�ܬ�8	V�U��ns��X��Cv	��9�e^�M�]����鎶���q�V�����(������vۛ@vC[�L�qӼ�]Ga7��K�����%NJ8��Z���u���)�َ�̳�gwX��ϟ#V������RӪ���֞Un�I���H�p0�b>��z.g]�qY�}��iS���K�kCY���G7sg�ѻ��c��"��d�7+��M�kZA��@���w����E�t��]���|L�[�8��p�{f|v��1*����x��b������g�v�U�U���_��1�4���U'���S;�����z�Ẫ~����o4��w�-��JjL��O1��{jm}KD�`'V�Z���.���<a��$=n:z�$�9H!k�\r��m+s�:�â����9�3cyB[=��R2�#��O���9�ՍP�B�\�^�緸��Ne�V��ٷ��s9vNeMYs�ٞ�"�!�PΓ;;��d�(o4:�UՍف�ml�;�7>�5k�f��E����N�z�N|ӷ�B���u��9BCf����D�Y,Br�ۧ�ar,�ˎ�sk��<=�1ς�3��~�pu���W���t�X�xq�S(Z��0W��&V�p�f@��D=�z�kp���*�b���A��3��cE�����љ|���;���Hv�����`Fbv����CU�D*���oHm�Ms������ь0���ɦ������fEۦ���J2OP	eX�C:�Mdeh��ޜ�	�8��G��N?2W �%����kf1�MLL��h�PF��l�m�{�dӇ��x������ugv>
 �w;zO=I�uGj�m»�|��Э��`��Š=��^z����9-��nѣM��'n{-qa�fy��;�p[�q;�\��i�~5>֙רM��1��29��;Q�+3u��WT�'�Ј�z��E�#'��h��E�����v��:�$r�Y3�Ƨ�����<�)c��^�i���ya~�J.nw�_��b�wy�=Aǈ�xu9­շ"C�WS�j�B(�3�KU,��I;������O�Ҙ��K/]nL��C_\�	̖���v������ey0���2Ö�[Օ�׶)�6�I}�y�S�-�#��X�5�o�[y��cV�{��Ŭ�_3�c�cAaj]䇆������.�U��3����w`��}1wgb���A�#�2��wiX���u����e�o3�x�L^3�Ƽv;�����F�R�׾1 �>��q���������I^���>9جن�L��^ӽ��8w�5H�7ˁ��7U��כ
���J�!WMi"<���;V�<7Ej'Z��\���w�.ջn'cM�V����cʻne�u{]hx�6S���C[��l㜻�G[�V>_�rhB^X:�wQx����j���Z�0m�ݷm<��C��yN�n�-o$3]���<X8=@w3�	�سج;q6�]�@:w�D���S�7lttf�b������YR�2�'�]Իݐ�v\v|�n;���l\\��Z����a%�>��m�aιcnѱ�/	MFd��	�!�ockg̸��Ob�!��=N��qP�v��3���g�u'5�u��N��}���D}����g0+�:�ԯRr(�x(��v��&t�]�c�44�;S��*maS���>���J�*VZm�lCb�%�K��ϑ<�i�8Z/{5�vt��ލp:+^�V�p��i!�w�lcڋ��uCo������Al��Y+�{~�Ѱ�"�$^N �'��T����q�����_uݷQ{�\&���}��E����;6oĖ��r�m���*��
z��H����i%�5;��Cwt����Wk�׾oK?���G9TԎ�6�c.��m�H��D���s���N�Nl���*|�-��^�5럹��^wc�&�ԇ;*y�s�&�����|�J�>J��16�Ѵ�4�@F� cˍy~mI��&�v��P�8HXGR+�=�3�F�՞!q1�*��&Ճ���ų�Y��Kr��\]5�������uޱ+Y.�d�%���=�396�#�&Q��j�-)�u�D�H�ʭy����e�8B&\������-3�)>׮z׷=��f{�7y{���8��
`�n�z�:F��N���p�K/^����@��,�h>KFϏ�T�Ɇ��XQ"i�.���t)��*���i_~Oa�ʊ���?�
l'"�Mh�F,�n�zh�ݲty�5o^{&Kl�5,
�,��\�&�|������W"e/^��#š%|��5ݰM8�'n@��&�ɪ$\�s{OZ��rkZ��Z�h�9%�*�ן��og�2ͻ��hf��v���uF��s�(u�E7��o[��Yh. 5d�=�Э�bU.�-�ru�~uadE��j��1��w�a��i��I��I�McX ���uR�jw���;!�t����޷��Q�&���IYb��ٵ�p���}����bAf[H����ówn�b�n/n�Z��8����|!Gv.����T�Z���d+$��'�j�9�D	���~�3�;�0�!I�Y������}��S�v���#U�,��ҩ�����oU;y�E=a����VIfWMu�w1?��o�_4e_f�> ��A��'ܟ,q��
,�5�R��C���]Ĉ��aS�ͭ1���������p���grY���d��W���gb���H�ˌ�v=����$�n�4á�٘�z-�*�y,e��*ϝ�Զ&���hs"�����{w���9*�m	Mv
�e=�Yf^����걌�[Y��ʝ�#�wq��n㑸ް�}sJXZ@��fU�2��*��Z�Tv�ml��G�,4�ݑ/\���-֠c�aDC�1NwC���vF˰`�]s	E�Q�v�9F�(�),��~u.���؅_㶆IIa,n[\�򳖃�LN
.k��t ��\��d���y�=�4T���-����e�E.j�J*�an��Ǩ�q������|)�EJ������r���Q�v<�);s�}�Y9%��썝ìP�L8zV�mR¢*��Kykj�����ۙx�G�`\� �>���$��N-"��:�ʅ�4�L\C�KZ�un�P���U���Uw�w,�]]Iy[sr�Gw,���w{.ڲ�q��8���v�J5�o���i��y���g
;:x���X��K���	n�����d�B�
V�x�y��o���3���]�L"�o4	Ő�U��R��!�MƉ*��G<�q��W�����1�\���ך�9����j�Y%x�q��=�ch��z1��p���X���i#��6}wJ
�dF��ws�E�����)�>K��|�Y�|M㬇P�Z�>J��B��lP3h�n(`u x�H��(,�[��5l+U�(�S$��l\�R^�~�����\]�.��>'�Wh��;����NaMZ�Sǭ�8�F�uW��E��+�ꧫ_/c��v޷�r!��^5EV�87��p�����ŉ��_�a+n6��X\3���7�t�m۸[�SBm���J݁�.�ˠ'0ٳ�ť-�?�~��r}���z��=�>�1�d<уK�(Qg;�V��� �i�(�L�OlK�y�;�S�W\$�3';�.��Y��`6�(]7�.z
h��9��Q�l:C���y�A�^�4��Y�˔,�g��VE��m:k`�/]:e��f����Q�w.�e��#���[�^Yk�s�i�=��&��ϗT�l۝cZ9!�Mvd�s���
�\a`F�S��QG�W/=�9]�U�J2[l��l����`��6�z;^[��1k<�Ji4',�5�d<�`����gn7m��ّ��=�N�s�Hir�u��u:���;
;���7'Ȋ�j�쭯V!d��6ֱ"2��I咬g �d#;��+���V��*U��NUH��lW��6�U�..�4Q2�lV��ֽLF����U�Q�Ooj�W\^�hcr�� �.�������݆�]�h[��e��lp���q�%^�������m�r�GX9�����PNA�7��Y�ݞtaISp ۜn��=������tɴ�5�b^=e�8Ʒ=��G"���$� l���ۚ���M�ϧ�;�<$�&f�1c̼<su�c����.��;\#��	p3�����\����ͮ�΅@u����������q�>t��\�%뛲��}JuP5�\�Z�4�V�-lM��ڎ9��%m�k��X�Y���J�t���&���c��zϽ�2��7�O��ܞƪ��+&��zP7\�Y���K�������}�>��qq�+Bzϧ�uZ�,�X�	k��lt6"�3[�S��3Hץ��>r�YUP�[�WSM�wu�n:t������hL����ˁ�aڷ�3��v!�����8�%�+��s��z7���]�{����h�y��VuM��n�/$�9��JVa�[�7��y�.�͘&<g���4)*�9�V��ao�<CQl����~�Aζ˦�iW#qI�0�6�ھ֏w/m�T3����0���Z�Ɵ����Z}���Xa�IT�i��˳�_��8����)Ϙ�._��,-޳qr��ol��uT���\��IY���y��7�������}))
���d�Zz���ڈQ�.�n�6G͈+��B{��΃/c��sh�W8(�~����T�D?,��i�}rT�I�- 7c���h`��}��T��^�E�����T��ϽSKb�ٿ,��c���-��V�W$wiB��;5��Fg��9��V�;;�N��UYET)�a�}rTԺ������q�M�3������rV�%%b��1^mt��]ҧ�������5��En�>� ��e4����e�>��y�P�G%Q��j�q����K6.�]��fWH�\F�	����S0N3���d(^r=oLF��$i2�����J4���k�:l�5{�⧞ ����@rs���iҦ��1����G5=@& ���x�U��-����#am�q�[6�TzH��1�|kas��^� a�%���x�Լ	���wɯV7�=e�ѕ�^;yd��^��Lj;���J��J-o-����R�N��JG���B��<�҅L=(�r׸�K{;��H�CH�$���o��=x��g��Q9�2���sKs3j)�����A��7���CӤ�n�!�۵!��/�ie0ݵk�r�华�:�E��˾�a-�Sy�ݏa��G�\��ޣ�H	����H�\�C!��yN�s�q�[!��,�o��1�{���.uKmW|9U�r���T��:�P,� �]GU�[H�
�M5���$$v�?�gt�|����>��戞l a�����<��^�WP=9���,��3�	���r�d���;��}$ �����6+!�s�]n�=#���\{�r�{G���9*A�u"�2��݀C�"��oWsxn�4L��z�mX}�Ir��yz�?H��P:k!�4�2O�$�"ɷ�D���Q���$Q� ���m c�D/8k-\>��r�Tu;ll�,��oZg�)�\�R6{��l�>ih��(�|0��ީx��#�|W�>od��$��^B2��7�,���׽;��a@�,��]��Eܻ.p�˗.^Z�y��bu�_/Azy���i���"�[�;o=��%��'9�{��Q� (����������Y5�ݘ�����o��S��a�63�G�`{0��d�yc�t���ؓe�1�Ldk�;pj+�Mz�=w}� u/A�Z�ݳ�;�V6<,��ے�B�A�B�M�4z�*2�@��>E�>޹�G��>| h����"vF	�NbcIpP����`�0�c1l��{t�6���b&�ƪ֏�0�X�ȗU;�`4�mh�s����3�
�|�<�	-/B����Jwx�»lv'Q-y_.	A%Χ�y� :���
!a�Fqy�{��� m'm����>���
nܶ�^Z��El�-�����1Fi����w�3�����W%��r�K�4qƃo
r����4_3�v�����P ��ϼ��A�}�.���A��{:�Q�<F��d���^��݃m1˦��>&��5m�oV4	Hmgi�-�����Us�$�dUЊ2-���ifS�~�Uޡ�=S����4z����Ӌ���=>_lH�ن�Zt��zF�*���urVg���h+�.�+g]�t��,ь^� '��2��{�i��q��hXk�\b����2���Y�,���w�5��:a�Ig%�#,Z�y1Л�3��Ӡ*ժ@m��zy1]&��ݥ���n�۞3����qH�D$����%��ζM�80#E���x/lQ��m4_7�{�H�Km4�4��Օ+�k3��Y����F7'�}�'��� ����g6�|��o"4�1�1��w
��\��r�*J����,�#�-�LGz�� ���=/����t��q�@L�����P ��1�������uUd�>l�<��s��-@}銐�Z�T�qᣍ.���w�Ilu*����0�A|�#�@P��<�d"��%}��f�� ��6R�)�̵G���n�0=�	4�v��̼���F,(��v���-%�KB�_6��ͼ��( C���k!'��/9�ң�ax:^�=PQ��sp��rr06��F�6�ˈ�'99�J�r��'xy�T4J��U0�n2.CQ�vef�b�N�M��ْ6]�B��|Y�w���~3��~�@�$��� �$������
@$�}X�@�� �B�^\B@�X�@�#��$��0HJ�$!!/��2�� @�I}��o����;������kο��������:�}�����$�_���'��� �$����$�M�C]��}OC��?x�I%��y|~\A����]�~����ΐ	!�� BLBB؄�/Q�$���.Ͽ����I�+�<���Ǳ�I%��+�˵��x������<�P�I%g��|=;��i�K� �$�����i�J�}M��!I%�U���/�`�tV�D<��A�I�������O���K����Q��~Kg��B	$�=߰@�$��ǧ��}�����&����/~Y I$�C߼a�{c���>���$�_�U��@ I$��3�/��c��PVI��Ȳ vVV` �������;>杖�+Me�4{kmY�R(U*J%QUP��J�R��D�P�IUT����ء5��J	l�
T�"se�BW�      �                              ��      @ �R�zw<n��B���S�V۞���ړ^9�R�� �ZQ�q�؞�*Vwu*���׶��x wHR��K��U��Ƒk#{wY<Z�4�z�)' huJ�ԨW\v^���҇�];�u� {�U/^\�]��]rKT�mW�z�j\�!�[`I         ��^���]g��W�mR�ZW[Z��uJ�{� �ҽ��#QJ�9�)V�y�z�U{��D�` 6z�-RR�n;W��m�ЄIfԵ˩u�8��h� u]*�hJ�Yu�fH�i�\��T� {R�W-Gf�q7U�hr�:j���U"�P��Q�         ��Uq��.��v�N��ż�tSl��<G��Y�� s������U�c�59^�E/&���^-{V�E�� ������L�k9n&�t�d�[L�Seȼ��M���w.��8 �F
%�v��S��.��j(���#��5Q� z�m�,��uZ\nK�ɧl�YN������J+�ٽ"Rk-2Km         ��Wjm���4��^\���ܔ�w(��z�^#E.�'� �v�j�G�=�Hz�3���h���Q�w'�R�iKz� �k����ͻfZ���b���١�I<�(�����z&1Cz� �KZ�sr�F�I�5���q�x��ڙ�x�v�fحo< �����mͺ��ΚUg���^�����zw��UUm�(:���P��        Ἁ)�nY�y��Zl��vZ��F�Ŝ��mg���� �� ^�F�����ܻI��]�����݆�G��*VU� 7u�wG^#���v]r��EU���<�ת趭��`jz� ��Y�mūǷ*���z=z�aI�p u�w�4�@)�x z  �:<{ �� �z  ��� C��OC@U$z�  �{FR� 0 ��	=5M��"{J��   S��)T�=@��D�%I ?O�??&7��~�<#��2��X��lC�NNV)�X�˼J���kYe���rT�\�Tq*F� (P�������G�������qfC��pf�K4���w�ȖlZxv�8�[�,0ixniA�3l�ӏ	t�9�Ce�U���9RP�n��H�$�B�8721`�j��4�X��z�B��ϳc����X5��rӊ��Z%)�c�i��+1����v���,[hY�+)�G/!�IG5�Y�zj8c�r��)�[�z�ʍI�Ǐ��P{�Y��6�Ȳ<,��+b�;J�؀�y.!Uz�{C	��u��ݒj��D3C�Fb��Q�9�APm4�;�1ݍ�{��[q����B֪H����75`�So�%����X�X�Zu@ve�᧟h�{��D�V̳q�fSe�T��6J�{y�2�q�(Aq�.�7Q%�5��ś��ee�M�܇R��w��݄���K���ђK"]ᵓp@`�!��fb�$Z�]�U\����t{rP���ya��T��h�`��,Mc�]b�Pk6t\�PÂ��Y�C���mmLض��U��x*Ķ�	=*J;�@�8Yu���o(iǊ���>���%lP�r�Mr���V�W9AJ��UECKx }V+���9ɥ��05���u�+�h��@p�	Q���$`+颃�X,賵�@)���n�6����Ah)hL�����%dc/u�*MߋZ�A�����!�����zYPUN;���LV^�'OU} �-�<RN��[�4&�����{���M�+M�x��M�j4l՗��P�݀��!� w4�)H��VE�HKT�M8�;��Ppŷd��ݚ����zn�]�ŷ�g*GU�Z�"����F�$c�2��U,�ذ��j�%�i
�c0�)Yb��t��WVؑ�V3C�G����TҺ1�u�A�5[�R����n�N�!���41�Ͷ���^���-�!���N�Qq���Ηۙ��ꪗn���%�VN$����x�w$�s�WJ�mߛը3���6r��Xq�U�D'fb.��̃�2��E�;M`��+��X��f֗d��YLRv��eVn��*c6{�ˋȷTU�/��[�wv7k����j�Y������N�n�����F��W� ��^�UilH�p���t�鶻%���*����u��b�J�����+ H���s���ʗ2�&�N,�NV���E�40�4�֔�l��E:ځ�ݽX�����Z�ʭV�M@��Ɂ��jFm)W����H�k)+z- ���f#j�e�.!0(U�u�0�!�PPs�t-�y���Hcs�����o�u���o*�T�HTI)�u���Q����A�9�s�]��v�2�|����A��m�3|Rq���b�Bn�0iৡv!�UF��*�O����%T*/�%�ݓjѠ��j-�r�a�x���z]�U�>�x4���5��u�:!
����`ǽ;	���Wm#W� _I�2����21�;^^e�\Dc�ˊ�N,fC^"(Ǆ
��@9��Om�X�Jrb�zF5�j������\�/,����XxY�x��:�o��\���e�9 8���B4c�V�x*�_<���mH�:[���ͬy�f�Ώ]����4j}��۶V	�_�)X.��b^Ⱥ��n�����b����{FT��g%a�mᗱ�bn��7��S�;F$0�'֎����h��wPwB����'i K��T�ͭE��,Sb���t���[W�Hi=NKU����a����zA�ʂ���AJN� F>��v��5zc�sdϴԹ5L-�=$AH�N�(ʺF���o��T��5^|�}	��P(�+j�tKw��/]��nK�H9��z=����ة�%�0ict�P��r�n&��ђ���Y1�q���R����s�%a8�U �u;7��ie����%�y��]x�r7�] j=1[n�(2�ݛ���,\��u(�8�.�(jg�n�������3B�	7�@�ܳgwU�����fV�8b��*��v�3-Z��X�34j�ꗸ`�1�feY-��YXu�Dl�Ѱ�̂J�%�GN�U�a�%<�;<�挐ͳ���(J�]���+k�6�!	4�]���R���[;6\�/]�`�p&/]KҴݚy�M� M��*E��V�[-X�R̀�I�`ӢU�vn�[#YQ#5���w2i�
���SL�.6F]�XD��]�`P�eɃz]���s��mѡoq�3�Ĵ���ڕwpd,$��!�L�%�WZ�f�x��6��Z��ows*�!`�ouGJ����j���r�C_9j���9�����E�	��{Uw�^݅od�b!�����s��Hh�&M�r��o��@��R{w8�}�}�EBā�P��X;|��շ����kZ�����)-,��&���$�a-{��ͨ��0�Kn�Ra�*��^]��ؙ8�H��YE� �@ks�T7Z���QZ~�!~�, L�*T|+a��IVNCI��&=��c-�S-\WBAM����xj��Y�j�N	Lt�v�	E�Z,f�����T���h�NQZ�"n���X�׵iS/c�""CF,�v˱t��׃`Ģ�`���1�e+iUH@%���"���i���6d'&C�����B
�<��zk5],zj�䑘�ݱl�$5��T�2�D�y���Fbg撘����=�!/DջV(���f��*�0͔�=h�F���q�ݥf�f�őT��T�"�Y���/1���0Q68+l=��r8%���m�kDt��ȃ��P�y@e9�V	���N^[��m��:�YAVTg�Z�����M�$��!<�v�RY��Ú�C�����EWZ@�:�@жG����i��5Vi��A�⤵��i��c*�c�p��):�U:)�KIV������҄l����L�Qł��74��7I��Ir9X��cQr��!=+��p� ZX�ڹ�!�Ey��*��`��6ҰAl�+�rfD�W����[6�t'#�;��*4�Ը"h�+�B�ٻmVe�J���J�%7ubwz��b��i3�sw%��/dZ�L�D��)�GN��iVpϕ�伽�0E�-U1���+\�ν+7��!��ӯ�ñ��ReL���^��T����GS�SUɁ�{7n�ue�`�f\*�wR��:��";N�K��X�U2]�%`�i�=j4���O���fw�nl�Z,�-���/`znū�5*�l7p�vEĴ���8��B�^["�����d��.S����ŎL��yS"���70�)6R�p\t2���ʫq&^E�a�eL43.mU�u��NXWl�7�����������(�d�U���ݱw$�GXU�	:3 ��:]�M*��­Po4����T��n�p`WC..bU33ng҂���e���tϜ���T�$�i �z�ڣQ�Na֖�&�d�t2c��{(X��A�If�n]
�O�|⚮�}X�|s!q�]F9����|�_>=Z��\��[��.C����l_��5�.���/�]K�������!�cu�u��h�qjܾ	o
���F6��#ԏ,R17\6u�*`�o6p�ƻz ,{bh�#�S�4T�]���`���4p����H�4�2���k�*���f�)��7x���V"�5�n�N�ީC
W@�۰2t��Ʒ.Lȶ�2Ƽ)�����r&�Ǒ�u]XvȰ���;ՕT�&a��z
8n��i��]�$m�5ǹ�t�ـ�jX��=�@"�7�7d�/�nӨ��N��xPyvo0�+U-?j�/m��r���t�n,e��v� ]ubY��l.�$�&rʘ��y������^iu4��D��*5�0o&�[V}	
��0M�mҳr@�f�I�����.˺��zS@��D`m�p�E����P[ʟe�M�I;,����VDRȅ����#�-��5�H����rlX�9P}�ԕ��u7t���D�Y�kiS�6U�q�B��vM/Y�n[�y�\G ͧ��J&�m��؎ü$1,G��F�'KSM�7^ġ����U�?�d��2j�t�Er-5��*�0f�4�U.�6/V��:�1�F��i@ب1��ʫo�V�1��*}
Xv=%Y��r����T��c�0ޘ�����i��n���Ï�-��d'l!��ʎl���5�N�ۼ�c1d�X�\	������/Ra�[#�1���\��F��eێ�w��ec�h]īlugl� օ�Z�t�׮�%<m�n��/�U�j�vh���#-+��0V�z�ٯ�T7>A�"�b[(a��BښcTu��aM�*�Ԩ�[V�1��Y2�sۣ���D�m�̣F�t�wih�7I&b��K���L���XU���nk�he��(ӧLa��c�����n�-K�h޹^�R���]/��d�!�v2�]گ��y�\,��f\F�u]͕b��sm�H��OL�*]bu�Flt�m��62Q�++l;����*!'o%����KJ�{Ks]��dR�0hj#xv���q��Y�MP��Vf7���5Z�4n�ґ�T:V�tT�.enM%�pYԤXM94�4���,�Ȯ��W��gM1gu$���e���Eڷ��'�;f�]9D@U�t�M6�8]�z�v�4�X��b�˼��4@hZ���=8FmӘ��
ކQY�K2
̧r�3[�;�b�A����[��52%=�H�I�N�jI�w��r�W�-5����/Z��@R��FP���ʆ���v��f���r�ز�i������L}7
W��C!����n]���:E��K�kI��֕��S��t�V��6j=�f�9�֑{gu懹����&M�
�6v��Ř�0�5��@�N��(4e�ɘF#p�M�!�3oh�z��`�v1���K!zBH�:�R�s3V;6[)ۼ���	�Ňm�+Tct&P9bѹ�@ga�f��;[d��lmH^�ћONhP�)���])X5��%�972�n��ׯo!��U�(K�qy��A&r�[�b��Cs�ko>���sr,T!�b;Jۭڼd욱�DU-�O�0=@�fޝ5x+��M����z�g��O�u�l��J�,5��д֬��m]Х�n[q��J�����񸩇���$�ˬʱ��K*L:%���ks���;��t���8C��ƯD��i��W|��Y��Y��u�Yn���[P��i����;Gq�	#]Fb�KuY�Y3Ul�Ӓb��7�7a	qӰ��'buvYT�),[1aƱ[,��s6#Jd��}���U��h�bٙY����ҁu��J��=x^���C��d��Va:Jl�
���XH�ֱv,���=k&�lpB��*��׹�^Ǒa�"��٨�*H~�b��^�6(%ynb�um��Mgt���ar���U����m����ʘ���F�sd��v��ӂ�:b̊��2Z4��ݠ���5��6ZXr��ݴ��E>*[�l�=�#�8j<���ͶR�Ig�o��4��{|�U9N���\�����p��q�U�,cu��;�Z��4�b\�me8��U���{R��r�m̶*	�d$��]f�ǃ/R�h���
E}������Z�V`��5R-ʊZ-�*tNV]�M�oFi�"=�x\�N�Ÿ�i�"}w��E��I�F�9EG��tX��>������G*f�P��FQ��
��7cp�2�e�Yx�(�k-7���O����H�SZ-c�w+/2n;d��Q���-��q��R4��M����u��[��.Zuc2�OƢ���9����Uz�A"�^`���h<�[p6k�i�\���:��i/?�W}�<ƺ`�ѹ�l����"4�y��u�mR8��B��F�8^Y2)�C����*��J�C��B�`������x�'v��2Xs"�~"�a�Գ`̶�60[�y�n�W;y��P���&�x������Óu;Zּ��g �A�b�6�!)䣈���[�Bд6s7A�I��漩��Yh҆��oV�-q�q^Ԧ�۶�p����g*�|�-ѡQAp��h��MѴ�8���h�S%�djh�yJ��,���fn����۔3
�/,m���ɰ,&�bnD���j}"-���n81�zr��lG5RZ��6휃pذq"K��)��s>Zm���e}d�i��� �:��`f��h�4�j��P�7]���Aj;eV\�f��xR�zƐh�����<���z�wFƟ����4�ȩa���$�6(%W1��,����A�-"�&��o։�l�՚��z��,9���-*9j�a���۬{�(�-�9tX�M���ך7��. nc��ѹ��eV������lQ�V�0n����٘k�Òq�iК�Պ�(dx(�[�YWSM�84���՛
�˜��w��B���PP��PM8s�ϼ���?&s�[�I�U�/zgq���O;�Ā��W\�a���|o0��l"�����rÂ[�U�5�8�B�bF�!5W��^�Y�X��
�Zb�v�<�W�7j%��F���R[�2��и�+!`ܢ��n�ϯ0]l-9$)�����7��0E���H�.e�Tr� mE5rګ�x4Tː� ��hڼ��v̻IDpӶn+`;+U�L��n��R�U�;6�zv	������6�řN�Z,e	��en�%h.^2�\�A�Fh��/M�n����6�,��xk.����h�+`��� 
�f`\���Z�����v[�h�8���O��W�۽��n��Z�if��x�x2�jZya4֩6�6�����ZęD��,�zJ2K@;��7��6"�}���b3M��l�nlW���6�FU+���y-.����D�P��6OҴVa���J#��m%�ڃr��	�c`^�Wj�.ڷ�W�Deڡ˄>�Ue����_Vi5�S�t��q��RInIT�5uV�UuUUUUP ʷ���着����U@�ږ
�Z����U�y��ڸ��Ի6t��TV�T�p��sW.�UT����J�=������{<ʼJP�<��j55Ԅ����̠0��r��e�����/M��E� ��ڪ�E)NZ�v�%�_/0q�V�UU*ƶ�mu6�����^[��j�j��8:�V��j���j��̮�Ѽh����k\�ܳ�y���=pe7������b2��U�����MI��V�[l��;���U���М�l�JO7g�9wOv�j*u乮��ν�nO��ٸ�BV2s�O�ծ�oZ�J���,:ڞn���M��]�ZΣ�G��y��Cun��{;��cb�N�\(�G9���!pZ�ɲ��xzM���\֋��g�|�p��ݹ��=�!�X���3�1�b�zo�j*�A�ۓ�;vp\D���t���ڣղ$�X2mOZ��26��InWD�����ċ\�y��x
M̜gn���D{6ksϢB���δ��ս��G�Q��x69�0�h��1����@[_��}�(7ۨ�l�� �OWY����uǃ���m��caج]:�;���r��;;�N�ФH��]{����,�z�Pg�[��)z�6��r3��x�`\eN��-cs>:�'nۮ�Dtq<���&����v`�ر=Ogs�}�k&)	��vplk϶�9�%Ӯ��M�s
qs͎��UX�d�q\�wg�;�ηg���	n��\{t��pr��*&�$:���w� �1��������m&�s�PyyN&N6����>�w��fa�v�������O&��nDI�;�8�k�t�gn.wH�#V�q��V��]�뮽5<�8q�hڛ�c�����:�J�ѺG�i�q��ĝv��&x�9�1�������G!������j׈��*�]?��}�Q��T�[�#�ېjD�P"I��a�0����&r�^stM��x
���J��n�����O�n͠u�S>ܝ
���.��N1`���n]h�v�7ix7<�Z�;���9綺`��k;��p���'VE��8�C��yp�^8��y���ì�s�xp��}�צځvͥ|�,�-�y�X��q�lX�g�ع^�]Ձ(T�X�ݓ���z�c��M����]e��2wV��>O��;��[:�ZM]�/mV���M���v3G����87�	aP�;�-�ܕ&O[^N����?�Qb�����(��շ�mX\�������O=���=Y������m^sԯn�h{��lg�ݪ���Fۂ{<q���RR]�{mֻ@��v�v���sۍ�3q&��v��']���ƺ���p�,����'������0�{�;Sn�X��]@|��O}����Z�L�� �cs9�&�Xw'=v0\�[m�nU䶝�;&k���@�2Vm�9��-�
ع�l��k<m�wmn����i��x��ۓ�x��v�[���m�2Þ9���#�J�H�۶���U���gv8���.q�w�ze�����]�<� v����85��v}��&񢶇����������7sr��7�W�w�0�7$�u3҆=�X3����^M���7`#Q���r��p��=�a��]T���=�����:��r�͹�u��y��:zw]�C��RÎȝ
�Y�q�����]����][�x=���n�����gv��&�n����0Nx�gw�k����\�|t�Q�L.ټ�����ӎ2�6�jy��l>H�R�g�sq��	�m�6ŵ/����.�^���\���1�jn�Á��	�V�C��-Dd�7Cγ͋��U���n�4m�	R=d�\tq�]���K����m���;�����q��޻o��L9��s���c��vŊ�n
k5uM�<��V]�:���g]�r��0�cC�y٤���Q^��h�����N���6�/��|��N�l����:�n7�ޯ�`���.�oDRq�^g;��g�u�8���[�ۀ#i��U�mgC�<[��ڭRn�d�G9+5�:y�,=ĆV�`�n�:I�Ah�5g�]�s�ۓu\n�\����h���j��	�/q�m���WO;׎br�%�ݓ�ܛVѫfJ��I�뭽����E^q�r=�%�<b��d�f#���nN��9�q#�^mcIm�ܽ�m���.ζӴPWnt�a�H�6��N���v�or�:5�+�����=��oQ��)��ڰ�sW�v�o#	K���9�y�s
��G!<��tmv�w��1�ri��kn��b۷G�Ύ^��������6D^��ju��u��mm�����xZx��v�3����1i/v�s��c�NvvɆ��݋g�\m1ȼ�q˷N1�W�ݐN:�f��Qͽ��յ��&��"b�A���Q�C�,ĹǶ6�Np�[S���۸|��yu�ӈ���5%h����۶�rg��.O����_gs�Í�v7�s����7kqݻf�y�9�+�ѷX���t�:8�=��ŵe��S��m�T���kW-�ֳ����b�F�d�ron��v�n^�hn-�֮���S���H��k��	�s�2=�ܛYy�kǱƌ���a`���n[�7��KLp^�R["vkͺxܑ�]u͘kq�9tx�TW`�yƝ���ŎS:v�pv�t��{`���X��x!y7h[F�=m��[�݌��y�4	X8VR����&��97@/"��b�k<��۵�[��l��l�V�]�+Ʈ�;�(�l;M��T�7�{�lVu�u=\����=�Dg��W�=<t������x��0vv�1��az�Y�q�n��^��'�l�M��k[Ӂ���i5��SY	�w:n�������g=�X��e�P��mn���;Y9�5`�v6�Ϫ�ۻk���[�����ވ�M�#�܍ڳ��u���n�є��Y����{Fta���n:v�6�M��Ƈ�O�:<�G�R_��Q�\�0��b�r�u�����K�4מ�)��;Y���3��n��;]1���[AO�{j�71�ƣ���'����n��]F[Z�.��ƶ�4��ajdF��ݳrQ/q����؀�.M�43�lX3�n���v�=8�rzN���{n-��P�m�Ӈm3{xx<�U�ٽuD���K�\�vv��&�o����=j�n�݂�׸=������pw�
�7O`g��z��.8灆�~~����x�]D��Ծs�c;]���ا=8Q�8X&��66�s`�����`�\�ػLc��\��G���׮�}����e��`���n�+��ln��T�����t��$n%{n��O�b�cɺ}X���!��ԍ;�\���v�g�X�b�ͼ��s��x��B�"��yЉr:C�f�x\�i�#�9��O]`�%\o���h�`�n��]���6�ދn����\Gm�����[�z>q�5m��\t�S�w�{b�ݧݣ�t{�v륭��KmŢ|��V����=ipu�vq�<ۜW[j8����M�Q�;Q�-3��&�qm�8��5�Oln����y�x�.�-nɸ���bv�p�'c-�z�3lm�B��s�s�Is����uls�,�U�Z�3ˀ���{�'�ݝÏU۹c[���)*��]�=W��o�Έg{v	���l@s��ݮ�ֽ<�x۫wl.f3�r�\��Y�����������c-��ro7,��'vx_=�y���nq�s�g��풮ǋ�[�v�n��l�X���x��bw[[�n͚:�u1�2;d��՝�s�+�M�a=š9�m���ћ��"�j��5Xݲ`�<`�p�m���Ed�[p��b����t��Y�c�
������wW=���X�^ػm���u��`�	��xN;^Ks��8̞۹1�
3u�)�rӜ�l^Z0���wF�e���%�g���)�j��]�1.��J�L=�<��֞�nsC���`���=���L8]��j��ny���^�@Z�	��.����8Q�5�����=Om`��{lϾ����������s��B�x�Z�cpض%n'۠nl5�⋰�����į�v�����860�ñIۉ{��r�0OHvJ-��؟Z�O-��0X������3"^��]S�;O%�sv���4.��{]p�رɇ�'Ev���Co���$&�n��;hz��s����7]Qn}�����lm�Cы:��f��	4r� �xƄ��s�)[n��o=��ŋK�۳���\�c.f�Pr�D���c7�47g �`�'`�>{u݇�pt�s�L�'6�k�.Ƥp;�sVG�s��d�7i��繨�Z�WF����n{\��.��u�n���"���k�kv��e�&�n�GKiw2 t��6��}���5<)[�������b]H���{g�^�s�d�L ����N��Ӌ��0��.N����J`9j���x�n��dq��nu�$96B4�㧱i���k[�˨�`��;A���v���ֹ<E�z㋇a�o$1lAܗ<it�\ˮd�;y���۲�&�y���Ѥ�u�d��nn5�naQ��X,wn�+��Xݶɋl�8�,j���-���;X�p��vE1�E �'a��^�p���/��ŝ�F�K��&ص�F$��NB��u���[۷bڵ��s������s���]��Xs4Ml�����\m�ź����i}X��.��{N��I=�qӗ>zx6����W>�-ь��u���z��͠;�c�y��D��,<d�*�.էGn��ی��ێ:��9�^�sX�-���v�7 D=Gf�ӻK�s�Y�7:��y�G�p\;��j!ۍ�]�����b1��9m׷����]��NH��6���l�kU�EQ�{Jv\&��uv�y�=��-m�6�:;=|�{;��ۺz�vŋ���y��x�9�뵸�岝�T���5��U�O<n��D�y5�f��]�/&O]s�Q���z���i"b���H]H6S���8��7l������u���]��kq�х��C��b��{;o�q��^:�q9�GN��{��ww��=p�P=�)J�
D�H
��"�:��*���Dbn6�I)Ij��Yl��:3Ǔ@.�I��4���'m�B�Lb�mA�=�cm����w^��٢��kd}wds#�n�Xf6�F���{ٜśw]+��#�ansҶ�û&f8z;s�-�^ZN�Ђ��m��=F�쐖��s�h=��.��:'n�\b<��qAtO`�P�S�'ju��wl:z6O:��`�ü��,�8�ݣH�8���p��PC�u�T�v��:�Sk��Yu��[O<��M�]�
������S�t�voa�̼tt<ܘ�e��\;X�ڐ6|�l�E�7Wy{G*�E[�Ӄx�!���A8�a�8p�m�����8�F�i�c�N{y����n(��s�����q���Ny���ݹ^z��8ho@0Y�ۜ���[��2΍-��q��{v8�9ϲ��'Kͮ�@��v��Ё���N��g�.�V��&�6�{i��0Q+���n"�6X\��nf넚��ɗx��N�A�i��3�um�U�
p�چܺ��G/Gc���m�..�b.�\j�{<:�v�5=��7nwV|w^û\���E�u1����Spn��ضfw�<�����=������ ��c�m�f��Zm&��\<�I�j����γ->8����8��P�=���E�1|9���t����ʎ"�� ���+��4�/���]�C����i�\ڌ�s��c�(Ѧ7����8ۺ���0b��)X�������;;�<��ۢ��˧�vC
��(��o ��C��] ����^on��3e�\<�%��<K۞�y�x���0\�L�2�y����'F���0�qa|'G6P�3���Wn)���׌X͵���t�d�����f�v6�	Ǒ�<qpm�/g�β�M�]&���r�����cr��8w;�^�h�v���̴ډ��]n)�z嵰8��<Y�������m�s=C�q^ӽ��7s��v7Bu/Xd�Xb�.�A�.�.���u��N]n�.n!oi�1�ԍF��bd��� *��
e���엉��mז�l���eh�ݣ"c#ۋ�Q�!��4ظ�����;ʷ���b9Ֆ���њ�#��kh�쭮�7]v3�]j��-�yq���zMZ���m�]��@�1���:�8x��v�%nG���ò	�cg �����pmI�X�M��7=��z�/Lܸ�B��m�y�=�ǯv�t٪��/HP=����w���P��]�a6Õ�p�����d��S�&s��m��H�攋������ˬ���������`�)P9���_����!��?Q��O��$3�@�iƣ�"��j��;S��nw�zh�x�����Sh�5�}K&�k���n�i�]�s`�j��Ϣ���ן�Q���2��qoF�}�T�+��oA�l��R�ⷽ8.��QZ�u�6�w����qX��i)� ��7	1�"t�wW�5���}\��pr�L��x�N�6�|y���j})5��Eef��B�t��i(�x�
�DYR&��-��Q�[L�4[R59*�j���n4 $�TlT�}P�V�t�B��+e�a���M�vD����b��M�ɯ!n5��;<�����kہ:t�����b�����#د�Y�{��S_���g��nm{��:�k�
��dQ�ڼ�l����d�C��#4$q�Đ��Ez�r��6��d��2ż���P��`{�mힽ�))���G9�Δ�FT�����캜����Q�,Д�\��(��p���0�mfR�$L�R�jו�4�cM_��[�p0z҆)!)Hv��6����`��+�H*�y�o^h��~۩���!x���,������l�)����"r*�os~0��p��\�d򡦂��J��Y�S7t����{՚�Ki��N�1>�6�r#���[���s�]y�>��q|����%]��|�u��D�eF%���[bf�+da�g�����$3	����B��s��:n����ON�O[ a��� ��-�`�䋾�������}ǝ�ך��Gr��;�k5S���x3��		���e��f��L�o�&H��䓸�j�P͵mX�B#&�ѝ�Q�H�(�7�t��W��C��ܿ��f&��y�]o�Yq@�1O�h��N$1k�J���A��:�_�k�[KG��#�mdv��2�<|�-�1Wl�D�x�_CK^�(ԗEˡ�(���vÔ��+b��yXD�(q�=��w���;�Op�fJx���8e�g�T���JF��<[���3���u�պ�~���k��b���,��9f��zl����VVھ Q�w�l�����l��G�8�PB>[�S�q%�b"у�P�y�z$�H���U���#�[���@Ƚ�0t~<OB�D���#2&}�66��U�{�m5k��n8���v�P�?���|�DE#���0�	0I!����C9���(��b�<�	���V��<��Ƶ��\��M�n��<Nq��0d���(���B�n��"bE�n1.�[��|�/S��[�s>y�x�N�m����`~Q��53LZ���jFc�"�:�/z�"����n�x�Fp͕��n0f�R�3.H���ʦ�G�{�[Q����2GX=�zx�,�b��R��j�j���M���`yy	��X[�=P�g�D�{�+���7/]k�d�ٍ��͝�o%_V����X6J41�V�}���\7U���nN'�^n��>�"��x�F���C���>2I������W�jQ{P�,�Sv8���$`ø�䑳4Բ�Iz��ǖ��s�^\4��`����q�xCF5Uۖ��˓�[Ϙ�zݳ�z.�5�v	9*�؞R�
?�����z�wEx췣�����)�k.{M�H'f�vީ�y7�qmuj�+��Bc�����[�g�-ط�J�S=Bkov5�<��0���,�7��T3R�x���b���M�*@�A�>�V%ƨ�+�{҅�+u���6c��Θ\9r�2�{{z���,4��#�x��ۉ�����T0Lb����>��C�s0R�^A̒�.�g�W�^�K��W�ٿ�ڭ�s|���++��h�q�hr*F�[C��ӱ[������hf��-�'��1��m�2av�Z��ߥ�ڬ3��0�d�ii����.�Z�N�`xխy�4uAS��pQ�G�P�c8TCE#�Dc�fɌ����*�.I7I��w�"	�5L("!��j���]m]��T��۝r���mz:�r:;q�g�:�k��a#۶�\��9�n1���)�G��'g�;V:�;m:6W������ۮu�p�n<��A�sv�2G���{�Alh]0���ذܺ�����E�}�����l�]l�uZ3An}�<�.�WE����`���]�=����.C��+\l�:��\��V��/=;���ջ ͮN��:DV�A�&9;1۲�nɉ����\��k�n�����|~��7&����lN��M��+\B��FSݺ�h�ډ��ez�KM0��0brEyX�"��~w�g�E�Cbv�p�wnN�9}���_�`r��w���R�ޠC�=N�7�(��1rI�9O���V��_26��[8w�|��j���z��uUS�oń����N,�>��<���ν\��[�9g�y|�gTn����f5
�\��.j�I���ű	i0�n8/&d�iz�yl�bҰ!^ñ<~~�D�S{=hլ�����Qc�{��g#" &^��.����2c�[��2Pi�S�1��:�l��4ep��m$��C�p�l6/��,]VV�~�CK�u�}~�q���>ys2U/aS<���l�?c���D�@���ƶ���W�����]�2�aou?���F���+{�Ԣkg���8�W�U��j�%γk�����&�m��B���ƅη���2�da���j�7F��"e�-���X:ݗN���:qH�3�VhKK��
�]	2E���t"��ҕZ�W��FqY$=ًR��#9R�/h��!CbG
N,��I���7G�H�Oz<���._z���xׁ菈Dr�r��Y��e-����b&"��2�t�+�o��,�7�Ԟ�sl����{u������%�Y޶m���z��NYf�+���DQ� L���9!=e�wsۏ9K�Ӵ��kg�=vK��[x=��TE����M�Xn���3OEsnvz�a�ň��t�~|��q�!:�Q�<m�Ӱ/BQ1£�jE��ν�Y��@�|
�=�l�X���v{rd��t3f^?T�WR�e��b�Ϫz�
c�2#b'i���37sݾ��	�v|}�����N�" ��qv�����a#k�#O��cB���<��S!�)�{��h���6��L_�t�YdB¥�Ai���yy�Y�mߞJV�4WY�B� �|��D�����rY3�Vw7�+���6u�w�A�����`��w/��]lj�｠�_f1�ۏ)M�v�w�1^�φ֣�<��k;уחR�/uz�5L���
[�N���U��	�׃ q6a�b�v.�vN��:��4�ل�b9���I؀PDѣ0�E¤���v�ُ�<�fw�kL��Pw]�۪oڼC�l<�����l�qŖ^uvE�[�Լ��B��=[��Wy�Vĳ4������l��ьw=��DPN#)w������a4��qz�6s�H��׽�5�FK�CteMɦ����L�P��fܓ.a�|��I�/��+ۚ��}���^z����=�F�w��kϒ;34�|;-E��,j�x�o��*k��h�^<\t&v%+�K'D�)��},�*��R�kǵϸ�7⬉�}�������_��lRqH�`,�*=��-wR3fC�5��}ġ6����M����ĺ�Ww���b�S|\0��N����[n�e᫶1`��TŮ�uVwN:��e^W�v��Ku!E��*E�<��y~�[�����5�/�\^xT���%�^מ�o�OD�3$�BHw^�Ɲ�?k��5{W�� m��f����n��/ik��ݲ���p�d�b���%�F��#�v4������ϳ�j�<�ƫCtFݼ��<�:��u�͇�K]�^����D�J8�1�6���u2�A� %��E�ؽ��U�'�ޫ���Ϝ�n���/P��HC(���6V�U��o��q�!�-���8��j1>��)L|�Dn�U��$��x�V���J4�b���ԇDV�l�&�\��a�hS���U�)h�Q�]����/K����N9�~�t�>��BD��屍65@�*\P{>�����vn�ر�tZ�h�"f#�{]�</��h\�v�n��?m��tn��۔�S��@�z��u�3����{g����M�T�d�0���m�^��<��Ɓ��z�:�\�m����{����fS�����Z��6�<�*qC�e�޸��K]��;v9��^<ރ���%Ƥ��ŷ.=E�WX��N,/��� �muθ�W9�e�۷,��ެ��{�Ŏŵ�n�dd%#�F���Ġa�[�k�w���.yߤÉ�ȩs>X���z��xR��Cޖ;,�õ�����$�0��O�n�(����?z��j;��z�3��.c���/-/$�~�|1٧gm�,������}h�c�6�@��v��߽wK�̣}��5�A�q�WF���[��𘏫��z�Y#���e+�Cȸ�f1��#�lN�+�MJز�aog�V҂a��ѐ�^��6s�<4���T��P�l/x)e�r�g���8�W�����DA�k�=5ԯz��N��U��OF���-��n���ku����+n[�|%��-���wfEdD5qT2���d�s��.;D��MSځ+\v$ic\�]�ptz3��D�n*��5�޷l�GF�鞵Gud�F���oL��RZi��J�dma�6�+�P�	�" �R8��Y�����D�k��Tx����kE��E�n8r�gʹ�2�:������ē��d9̣��k;�WGy*Tڵ���>貰��Z\����^�����9�ٕ�w�x6���)�~�B�h�駹)"}��(��4[	�\qT{;|�Q������4V�t�v���O��kbv��M/�̷y�]��鄏	H��(�q���w��O^�m'�j�Y��<+�V�>����^ٛ��B�.���f����\i��#rN��5Sޞ��r�����;{�w�ӡf��X��S�\��þڃ_p�w� �n�\ss��f�����=��9���=ujŧ�1�]vxv�u6��z�M���~������+��+˼�Y�k�K��&�$��6���tǏ��$���SBG$�a�ʜo�������%�ʞCa�b�,?\�ߏybqS;��;��[C�;1$-�p(d5�3�v�z�ӕJ���W�Om�Wg_�R��=-�\���sA l-�n��];�Iʀ�����X��R 7ΤT�PD��}$�i-��w�e.ݼ�jm����ڐ��:�'������[�&<I�+1靳 �-���1-�d�/ �2)EW��=b�*�oR&���8��f�����i�λ�˲��&>�,�l�k��G9C�'wn�ck�����]Y/Q�;��V'IF�ߕ�)�]�Y�*�7����|I���񼇹�+��܎��\����h�@�h�W���$���u�j�ܠ�.�x�����/mrru�]��)zYdq�,�Dj��So���2�$c69XѶ:�o	Lup�h�>�o��y�AV>	�8kELf\I�8,�Ő$5=���;6��w���K���)�9�
9*��P�����R�J'l�IL�g�C�Ia��Y�T�k,�o�x�B�g�m��U�ln��w}��8A��������:�𡰻�Q��%:pq3���ow��d�'gIuhŒl��@����k�˜��K;k*P�2�y�8�7�8]S-�g��.���4���|�J����Ɵj�&���j�{ �mU�CN�{�-V��[89æN'X-7���4�ZQ�S�}��^�2���w]��}y@;���uS�=��e�>�n�,�cu�f�U�.�2�"��J���-��kV��G�w��k6�M�ɕ�ծ��9dY��Ny��G��Q���0@۾G�"���]�9�q�/L��V��\Ճ&���
�Q�d�Y%��/�똳*��:��Rl���"qj�Υ��{J�˗#�g��o�⽏el��[������M�L%���u��xm��A����r�����a�ܻ�Vu{�S�Җ���~�1����[�M̕�y�����*���	]����k<�a;S��+���^��㞺.؝ƹ��î�z�kE�⌹!n<�(�w�i�5�~��
�JX�{�`W,o�g�Fa猗�6w�y���P0�-�3��Fu��fwu KAn��^Vn˰�Ȳڷe�S@�y�o��B��'��g7��Z-���I2n����;X�?W��mîX!�_��2n\��!z�*�ʽ�r��0���>�@�"Q�#��#�zu{I��󹚳]L��/���ϙɾ�To2��2�5�N�B�>1CPEhq��"ӳ	6U�[	I�n��(���k�"����X:l9�]sc��������|6�UN�>�9ozκ+�O��&!NF܆�f�Bͦ���1J���=�uU٥*o�z��Fm����s�����X��F IP K-�M8jp�q���\�ME�n=�.��j\�.꩗sm6��n}2�#'����L�uꞖr����6�k%�3Ns-ۘ��ch��JX����$�I[�������{��1�^W�j��f���q\Y��{���͑X�#6mޏx�@���dp��>�w�vS�㞩4��z�Y�碔�^�-,�Lݳy����~�~ۙ���<�v�6�d�cq��웭㡳�~����'2v�Y�b�{%C{o1[́1k���(�Z�c$�Hl��)Hۓ6�KOY��nÚ��}{<S����#����y��r��y��!����<�fw�]���9�|e��ꭧ��֌pu]G�L9�g-�E�ޢ\�F�V�>��/,�wZ����se�Z�[i،�+[jMb@ർ9�[g���ug�!8��'\�v����K�𩪺�m��m��+��)�A�e׷6�&z�z��.g�1�y�b4w��L�G/�j�`�M��ӌp?��7�67��z�A�ƅ}���U��O9떶�qB<Z����Y<]���W>�m�݄��b\�]�6��$&�'G�2v.�Sv���-�T�v�G�;^5�F�=�lݱ�͕�5\&l��o��ݪi��^Zś��O�0G$�1����f�8��{t�YYQTF�M�N��ڕ��J~����ć_�����'1�XY��6�Y-`YCڄ\��1��.�=鲆a���w��r��ƀ��T�<%�\%�	fG�����ｓi�;��3YM�{��!�[2��c2vXҗ5R�������&8r��/�����{��;S�f3^h���5V���2�#-Y�u�vC�{��^,�\dH` ���2�m�<�v�k��O��}n������l��ڒ��Q��`��m�d��_���\I�c�DPh`A�ReH
{
l;s�ػhQ�P�e�q�c�M��l�I�q�F�h@�5!i"�=��?w��s{l��xΧ����{~��w�I!�,��ﾼ�f�p�1@��8�z-���m��ӾAѳq)��v��Qg��\�4�������(5|�N	�E�ʬ�ܵ��y��!�,������;�gE��Yz�����M������n��7(7�k���5�1mh��xJ͛��=�cK�������:���5[��Sɳ�ՙ�{gU�:ϐ�F_�c�ϔ�{r�����y��r�~z�Y��	��|}9��x��/I��ܽ5�ʛ�(��#M���#ǕL�'6��+1��"H,�l��h5����Ь#'�����}k}n{��5~������=�\X�}��� Z3�طU�Ե�M�z6�:��k��rbz��a�ww3wA�~��yk�\(��\�~ey����U�G�[�_��ɞ�~�E��>i����oM���sL�kN2�L��X'����[�vw�����{�Yy�^���:��M�rB�W��'�;��^�{�7�ݗ�v�������zj���K��w|�w��4w+��O3�Ŝ_nӇ�k�٫WjD4��K(��,f��p�%���:���Gx��!��E"I�$��z2J����˳�t�S��\�u�m\gv����j��Ց����ce�e5Nۆ�(L�p�u�=�Fw���/F�R�ꈡ:ɱlJZ���ǽ�g�ÙX�����Z�bd�|�*
�|�p���:��F�c�OV�1��p��J���\�'rL@�IE���w����ED�|����O�S��i����Uww��9Y��[&
2�
9d�ڥS����Y�>q<�l���;;r���VNԚ����N��r"(�V�H(�E7#NS����}�{lMtw�v��bv�� f��U�7؈��Į�M��*;��.�Cq��0�djHq��Qtߢ�NM?m�յ���.*{�F.K}��'�;Ņ�hk�J���Ҷ ��.�uΡ6�s�D��n����s�§Cn�˩U���Y�A6-�,�c�h�uWԮ�`М�+���X4��ձ�g";��pc�	&82�ng_��l�ք�����6��72�R�&&��]����my��/z�օ�Ȓ�8�a�I0EDY q�p��/W��5�]s�f�)�7���>%���	�G���9���W�	�'�y�L0�zپ``���*��ݹ�y��j�=|���XNI�b]�\}f=��=���~ڎ�_�O��0�8�r�q\����8�O�$�+�L���&�Q!�;ު�o23LQ�z�~�[��#P��+V1�������M�=�;e�Y���� L4`e�[�2���X�&���9�����	�R�t���c�2t��g��=��Tl7f8��i;Knw�noof��^�G��-��j�+P��X�5x{����܄���{��� ����v+ʖWFFK�M��@���RL�.���绂����nH�5 ��sU@޸�S�F\�za�μ�4!��q�-;�ʘn��\��q��u9x�������vי��xї��7�m�u����������y�a�{v뮻\ރvw�J<�ݎ%��1c=�j]�<�r�G��o^�I:ز\�=v��-�V�g����s�+���b��c�����u�c�v&��ތ��}����ֹ�!����֣(>��M�<��s��G.�jS��7clG�e���d�����Εwk��6�q���|�w���`��� �h�rڗ�^x�<�v�<�:�i�Z��ā�#N�o�o�O�矱n�P��[6g��`ѳ�;�ƑW�ʧUŖ ��.�Iy���alB�9,�Z8���@���gc^��V�=sɯg�����p0W?zc#��"��WGR5eHCL�sK����n�ǆ����JK�屿b�''<9ar�쵺�=�'g�)j+q�[r)$9o;QBQ��*�J/l��f��<�=�j��K!O���ɸ����}��ܸ>,���-��R�^�]������q���b���O����6	V6[v��yf������W�ub�q��'xZ|����.��z���f��s�5�;$��::����	�H�l& ���A�Q�sgweW��SqĽ����H�|63�>-&c��Ӯ��%�Woohne���G�V]�~�݆�z��x����E�3�ZY������T�y���2��@��<l9}V'+x6*>G&�B�2td�I�W���ڥ�����Ǽ�͔�$�!&]�ߖY��`�V�?7�RP��F1a��)A{�"�H=��]&p��w�R
X���c����	QRٻ�u^��cP�͈[����I��qɵ�o|p����-
�%�����+R�C�L^ڻ���7��aR;���fLʤoA��0##�C���˽{'�P��#��W&�,/�����^�Xb7�����Ū}ך���:��<HU0�Q�J
�`:z��\lDi�7I�v����l���Y�s�z@'!F�q�������N33�uq�cΘ�4��[4�nA[�q�.Ѽ������;����%���F7�j@6>�i�݋Ƴ&�];�l��Myn6��k���2>�z{�y� �Q�����nBZ%�$�&y�ׇ߯_A�ݶ���U���t<�NV�n�#�kCj��g��۵Y�B��v����ƸqĴ٣�i�&-�J��o;���[e
�/K��k}Ң����ׄ*E����0xb2Cy�˻;,z�ǽ�A�ڈ;���J܊͊�̅�O�{-��*ቫ��n���my��l�!a���&
�0�t�b�}Ɯ�Ϡ�d�n^'��zo�ޯm�[<ĵT¢��~���?��`X�����R�I��<M�Dݩ]����֌���7.����t����nK�֪u�w���u�x��oͣ�x�צfk`G�~��H�����O.�'�;�4�����Č�N����$=t��������ֱ3<i�;�Q�����r�T[P��~36ϥX��^��iؼ�Τ�ڎ�#nC�v�j3ѿgn�gPW�<�L]�-��+��%��L{�ol�ש��~�͒2҂D�.���xC��ȷ�3r�K��=d��!8�S�2�m�YR�1�:��Z�*f&n�I�f�c�t׃.�6Z`��N2���l��C�`hZ���}�U$�Dm-H�S���&nV-���o��|Jd�q8RmD��w�5��t�gȎ.�5�V���x�ů��q��oz%���Fjڛ����7����S���tЏ�vhQ��y۬4N�-�6�X�xy�5Ő��l���B|��@ؒH���.3=~�9ƺwW��e���Jzy��g�v��a�]��e��_�]�ۅ��	�*|�-���ɳ$�=�e�]S���sX*����'z���u=]���}��r�&-�d�U�����(�Qě���ա����k���R����+D4�R�mhu��[��u��F�67)�V*��Z�Axe�Y*��/|뻹��(�����kd�VsWN�\�Z���w��ϒJ�,��g�n��s���.$b��[�71�k�4���=!A�Tk����a�1�=�Z��b�x����H5ϩ,�I�����-Y�YTk�ʙ�����7��}]�[��Q9E��Fmǃ��mۡ}�Ŏ�WJƩΘ����8!R�u��%����7^y,��nlɛZ.`��ypp2�^ZՑ�s7C�vcṜb�t���w+1����Hie$.�=)�Y�7�����5�.�˜gl�cx�x�W�sc݂��S�A;��'��W�1t���+�3I֎ ���e�@Fp��A�]|z����UX6��ǳ,T�Dtj,��ݚ)ֻ7�!T1�q뼮�]f�/jNe:�A��ە��|�Є2kCY�&�[�0p��ʛ�.bP�	��R���5����02�&���ά\�Tz�4 N����feݒݕ�$�Tꆫx`���k|��
�c=�R��o�X^��ŀ[1�N��OY��E`R�e�ʑ�_fk�WR��x�ې��5���:���b�5W��8����M�e��إt�,7j)�����)0mf@v�<�7Gx��������2�-n�} ��
u�x�3(�
����mTiM�9��:�H_�y���f!c���X�ܻ��G.%�v���������g��#�c9����'a�y)	�`4��{L�K^m�(��b�\�ywzDa�l�kH:l9L��(�i�L-�����s�g��ՆKI���S*��(�]u:OW��M3n�4�4�(�Tnc;��J��u�55�\�[�|q<�����rg�m�M�c��+0�0�_-����������� ?M[*�MQ��Ft1�� �ݲ���)�]Q��r�'�!�Y�u,�a�S=���t+Ӈ<'U���GNz�����u۞|7mdr	ηt䊒6�$k�N{1*�A�j{=�X6^7mң������K�2��Ɂ��c���۪۱g���E��f�ӓ�=�h��ugp����%ʋd���鱎��2c��2`���x���<�Y�E��*3�{@�d���t�	�НW:�6s�ݧA��VFs˽���1v^C�7Nݴ��[�s��v�pF�>�m���.�����xw'4���#�Кrv��V�����k�0HX����v�I�Ov�2�A�ĚƸ��a�5u�cOU���n�n�"��<�\G����X+�lM�-��#ԝ��ps�7��q��
�e����7E��v�>M�j�9�t��w�l@�v��j A��N탷��u�y��m��6�r�݋mí^'%%�� -{����>{,�ǻu'[�nv�n^�p��;���^�^W����8ǰ����"֞�+�����;K�=���{[m;(c��#%�n�kg�;��c��{�o8r��"�S�e�1���ۍ�
�u�u���gyЧI��b7c���aY�k�vΐ�T�ό��r�+�tmѮ�m�O>wEkh�W=���W
v��Xmsz�s�ާ�q�ۭj����]nOOc��k/.R�s��:{j�3�z{�Q�c�`���&p��|0����7]�m���G^���r
�2M�˓�7iD�붮��6�|�۳�ӭa��k�L�<���ȼ���[��p��u��\�헏�:�'`�6��jW7]��ݳ#����<�ln۹�l���ڷon�石���q��Z��N�0o���7��8�Ql������=�gp
]�L2K�:�S��v6k��F��I�����Ke�w��̓�ڱҮ 4�M��͹�B�,�v���-ip��Ǟ�cQn�{g��ln��Z��uYz�VDt=��bv�ҥ;˃)n}=��r����t뫲!p�ۆ��լ=Tc���
���^	��tA��U٢;l��<B	��ͅӭ��knk��ÞЌ�I<� �>�tn�iCGX��x1�`u++k���l��v\�رi���z֌q�+-�{7���Cdn/mv�g�0��ժ{.�<3�Z��f=��f���i۶	��7-��-����`�8#�=�;s\D=]�b;VyL�����nx��y7r�%Y@�C3�ɛ#��7��>��>u�:|��.nqɺ�6���E�]�+����zyNn�28�;?�+���9ٸ{�v�X�����Q]��VV�p�ُ[�X(� ��q2��@X��T��fs���]����W�+խ�O��߸��{���&�dZR^=�~5��|���KP����.&}����噞y�� 5���&�&Pu�Z(�x)�c^������D��NBL�$�t�ݿ,���Ĉu^w3[Plҫ�m�L��U{{-���+(Z��[�W�9���z�$$��!r;�(�N6��Z�=D>��.`X4�J��j�u{B覥��5�9F:�W[�Z>�gj��.{�	s��t�ufT��:�S�u��t��ó�Wbv$(�X�N�»}�<PG��o�i���\��vV���l4gT����=|�&�{Y��1���5!R8ҟ8䬮��ʬ�^��So�u����'��2�z�cN�u�C����·��i*��8�����G�֛�·mM�meV�q����3��{�ȵ��:�+9��Z�\8�Er����:�"*É���qI�y����s�����l�v3G��K��~Ѱ�ᮡ�_G1��7!����kr���<�]I��]]Dޛ�lǝ�4�IC�-�2�jΠ���Ǖ3:���^
'.3rVm1�������+kr}.��V�h�K�}��^��LY��kV�:�S��w}��&�q���@�)��7W��p���n0�s���)��H�^��RA�P�6�H�r)PƤ��w�=���r�x��X��X��H�fYF+q�a��۫��f��������%H
I�v�C����4/
A]CD� Ar�gI��Gf�o+/5�m��t�}��ci��;R'9j�rG��w��_����c!��L@Ԓw��ʢ:��.��ozen^�\6J��0�(�"��s�0�l�uchb3��ao%s�o:���v\�z�srGɽ�]�;��*���"��0��v�zk)��9�L+�yu�������}��K�c��-�ԅL֪�Ǎ��Y�=��<q/f��Q"�����I��W��J�Imy�so�T^x��22�m�I�W��|fZ�"]��[��~�}��ZAJU:[��/wuu�ޢ4�~R��Q�K��wiT������K���A��ѷXǶ���ć-8�%Și�ۍ㝗�ٞ�qM��R'=�kկ�8�,���2/���=���L���Y��(���L�9yqw�Q۵7v�V�T�H$���jZ��A.�jְK���^�LyY����DB�r �(�p]�j��Il]��N#el>Z�S��G&7vo�=�C�T���^�d%.\�hjl0�Q���`{�h��y�ߛo�m�9�<�/B((��)��l����NEG;Tv;1W}��C��]u*���[�����q��x��z]��g)�Uu�`�j���'������M�%{Ҳ�ǩh��m8Ɉ"�K��Ģ�=����h��5�v�צټ���I�Ȱ�5�V�"�M�ǽJU��s���<�7F&7gyR�y�ly�r����)s��\�(��M�Ks\��rv��C0^:.a���L=��O��k��C&h���Do�%;�0�[��#d�d"0Sp��Z|{,On�u�yn	gd�כ
KU_/jp����,fo�����u���#IR:�p�IO�rp��wV磱�mm߽�hR���5i��h�;�Zy$V���{,^�P&��s7#�V]��k�w�Ɋ&�k�45�ɺ�Ķ�M�D!�ˬ��~]Y�q�~��֥滑�GqS���{h�g��mAㅗ*ϳtM'w���N$><״s ����<���4�1�BF,u@PJf��Q�q;�n�!		�ʦk���q��^H8��"�aX��C��=���N��u�Ź�r Z!�j�i&*����rGn5#u���l��em��N��917�=�\�;�Ϛ�5�����M�q�kn%9@��R�D�ca䱰�U1��\x�n^pq�Ju���5��q�W������Nm�v<=���{a�x�y�fȮ�����������*A�Ƹ���iӹy��{�.6�o}h��w'B�]&5� ]�O��盬6�]�Q.��Ft,zƞ�����g�,p9K���պ��y���]
��Ƣa��n6`����7�y����������&{�ݬ(Y��D�s"�^x=�e��f�4�R2B����ݿH��
���}Z]S�!�a�������t�0��w��C~~������<Xig
�P���H���sw�i	7�<p4���V��"�n�[`+�O��B��%�vȘpєZa'	q�3lz������Fhiʑ"������fN��yP�JݛF����/��.avn?,�����/r�HJpH�ņ�����n�J�[���">�3��p��kޓU�W��tn�ξ������&����6��@�̍Mת+��bݦ�����'���
n pF��5$�����~�e^]����͑���z�h��D/s�SARr�\̳��v�V	�j(����*6c�O7#o��`֕^���m?<�{�����V]��M�,��S�Z7��}�]�����1�t�|�2\�\�B#�k˹��T�8L(�M���}˛pq�gǶ��м��~����syʔM�|��~��3A�?HA�'4C�C��5X��6sW��C�]+]�Y��z�kލa�o��6j]�y]ݔڈ��j��:
�����SwY��w���(��Kމ3�Ϟ�Zwa9~��r�:]�r$�&Bڐ��p�Z��6vi�(|��@m�rޡ��{��T]��+��k��>�rXŘ�C��3kJ1�D�Z�rl>��	���3�^&:���mW�B�=z\�s���m^]V5���NC��l��iї͹1�q�>�.��f�j<Pݪ�{cx4I���K1��&����� �,��r�L��{{d�E�x�����%k<�w�U��!}޾���M�e%���-ǚ��^���!�޲.���I,38V�z|X80����;5>�X�c^�EpLm
z�w�sk��
t�%�1��-N2��&m��o�A�W#�wX�=��LR#�z��(����J֛F�Q�\�w{q��Ū�ˉ��Z%��{;��;Ւbū�91�56�,%���k�Nͩ2]T������p�#�Y�zr�jnz�_<�\O�+�p��K�;~��7il��������̰V·F�^p�xI��Q����n�A�қ��ng�m�c���.z��f�H���Ĉ�d��$9�7����-TlZ�'^�\�$��s^5����6��U��N7.�z�i/wU�y�:���#16L$�pv��l5ӽ+v���DB�l~�Q%q�G��o�3����y����OV<�gvSz���#1&fn���Q[�f�0W�=ZǱo��FB�x��9힩�a�����ؤ v�!Gb)#w��#>:��4�Vs�����=#{���~@d�0r`c>�;���ۋ߷A�cyXm�]YPB���4�I����>\����=Z��;b�=����&m�Y<�ӫ�����@[9�9�<��
�R��0M��Ǻ�kk�����
�z���\^��� �n
~^�t��Ԑ��-��r9���0�P��ZK��5ԕ��j9<8�^�l��9m�fNwgZ�+�#�Gx�pݛ�&\j8�H���3U��z�`.�;���S�#}=t�^N�=!��p>�M9	p�cEA�VL��������hJ�we�L�Cc��]�C&�����k/�:Fv��hb2�f8�m��a���W7Y��qh�<)�~������w�e�+w~�y�G!�W.�y�Ij3��,S���Ź�]����"��fە�{6�J��zj���Rn�a���7u��p��ϓjd�n�?Owb����Ty(��
���vy;~;R.�
�ڲe.�ǚ�%Gvr��؏b�5=���ŧ��egX���l���{��DY�W�uU��AE)*�).��F0��;B��[���%�pT/�����5�m�-����n�i�K���v7�m��V�1�N�˺�v�ݺu�n9]��:W���͍t����r�2k%�rY4�n��n�2a��yc��e���7F�Ӣ۝��l�Ʈz޻rzݻ7q���ƥ㤣��n,r�h�n�%9�A���kn����V��lV�b�^7�g8N�۳3�t�2d/F;+z��82y��t7I[���1�)�����mKn��cu��G�z�r��4<�mU�+�&~�u1�ٽ�{�H�nj~W��M�K�� Q �7�{�Jݯw��k�Zi�
�0�o��t�9m��0ݱKt��,������$���{�^6��ݖ3Wk���$~���>��f��H#rg�o[��Z6���:zfOe�c� Lnn\��O�֘n�Wy��{���Uz�_`S₉�[�4n
�͹5g#1�U��D��ѓ��	��e�hÅ�z�{9p�˵�q���)	,��/t��足�7��.���OٸG�z<���,.�wCr-�b�d �D���jѢ��m�f��v%�z盳�]��7n��n+n�+�g<�3��������H����$���w����7�١TzY&�]���ژA��k����o(Vz�y��$E"$�)4Of�fj �����A�����fI۱������f��]�L����P�N��8�}�l=c4�?0�̦N�N��Ɩ=X+�D��˖���t'i��{t��ڍ�O-���W2�7(�K �9�R��1�b`�!J5�I��M��5{Ahʓ�]��+lo�/�dF��,�n۞�=�`Y
�s�0���V���S�ĿT���o����0�B�o�T�YY}�(z��!$6���<�Z�z�(av�Q�$R�r/np�罜�ܛ��l25h�	��<uv.�KW���B�-�n춉~P���������.�C�{D�k�:�V��X⺲:���]����7#�u�uvaT����W�ϲ��^��JN{�ջ�Ʊ:�h����Xv��O��m!~�7x��U�K!��q$�f97$���:Ǽ�Ol'�uc�c�QZ��Y�'j2�"1��h6٘Raƥ��ǡB�]?2�-E��ɗ�0wl�D�*�k�-IF��zw��1x�#&0�a�iA�ņ���Z����*(0!��V��%\7��'�(�q8�CL����\9!��Yz��8p;S�ކ�����s�ꥱ����[e[��bY��8�oh��i�;7�2aV���i�g�3]�lR�Y_l����ۅ���Xd|Eѫ�&��*L�YQ��Z[�6J�S�-�Y�^)�n�+����j_G6��A]�C׋eKp:�u�F�um"�'�+G��{#���*ۀ� 5�oZ,[Cr)WRL{�]=�qFP�k�V,v�СB��j���{j�%!j��#�qU�Y��<y�:8R���qΧ�����U��W�"�Grh˦��b���+��b��>�+=�/�R�����[.�`0i8vO��l:8E����v�#�R����cSl�n�L��lGQ�'4>=�cD�OM���.uq�.:�/�����le���8�-�a1�3��#��E)[n��#kO%��1��v���{�]�4_8�Fl�p�HJg�7WA��,��.{�S;�#G)�\����ٺ+,�{�q��Fp��\�t�m�y��+;��`�8,.U����G>�2	t)��/��Fmn�]��,u䱖��f�}2W�+���YNuu.�Eq}�/e˫=h4x����F@L��č�i� �����U���\7�}w2�rgJӻc�Ss�L�f""S�t�/0C�tΐ2YԳ�5�5yX��-��_-���;c�M���f�u[���=����{f�v���+K�עC���a��i��Y�Л� �m�d,�#�c(ߨ��0�{�{t>���{V���2_!�P�9+p�w��?F%��e�nG��^�����fk��`�����Xv��ٗl:���������خ�g9�!��\E��$SYݺ�/�X���OCQ���K�Ss���d�v��n����B�%��-�0t����X� �?[�d����p-��Eh��\�{�c���(��"h�b28�D��6���'�_�n��:�Y��3���מ��I�,�����]z��ǴL}��IkD	4�1|Xq�s����rf�,ɏћ�{���u�8V]�cu=F��<�7�A>��!$$�#R+�f�b�ݶ3��EJ���lo�}���(5�|r��
ŋ��O�2�o9���@�1�񿎠��.���h���kE��B�{֛<h���]��w�0.�|��oe�K}�2���H~P>9B�7K2�Epy�����c�d��q#÷!��vuC�{(8C�nڻ��8r?ǃ���Vsٹ��؆C�:{+3����u�K���>�ܗf7]vJ�+77fj��|���j3��dǗ��x�,+�ӳń FFo�S3X�0�Bڑ��mGr<�3E��+�|;6�;��WDY��������w;�r*����Z2��È��pI$y��,R1���ꢰ�ܔ)�-�,a��TO�{�������f3|�.o��ȉ���&\,vi#,�﮶u�)ʻ�d�|s�<짍�=�D��B��>^&�Z�O��B���1�vOG��l�kՍx�R�<ky�x2\���Dvd����CuL�<UC�ь�	$:.\��Up�}\.��WO�DpԠ�|>G����&���FxE+���8��k/�]+*0��lzM��I\I�����V3��.ND��
�i��y��6�;z��i����c���Of���Wl�p`����(���=�7�v宷3�&���[1f�{q�۹0�c;:�n�r��uv��6n6��[�l��ÎwlR].�:�v�)n2��:�9.;o3�=�:�f$v�x�إ��ݲk�L���-�cM�n9뭞�;b����t�vWz�����,ibێ�vkZl������;*$^lT��\�[v:�뱳�B�eD�RO��-���y�~�jd=]��U
�q�Rce�ʷO��otR��1A��d��r$�*Z�[�X�����&f�;���QP�Eu��&5j���ݻ�bYy�ung�x�Q"ԑ#%n扱B�{���g���/�zI^��%�9���&�/ὣ3U��/2�,G	�qɂ^yR釔���\w}X;\�yiEz/<!:Z�U7Y�-3�5T���r�
f8�p)qǋLǼ���1gB�X�U�Z�g{;ڥ�u�}�^�i����;#`�bDB��nu����6m�Ⱦ�m������{�|����1HA�H4"�9��O�s��髳�w�4��K�[�Q�evl0:��1����*���}�&䊳��5�	p�S� ༝W���_����Wb�a_�*א�UM��])bD���Tࢹ5�[�w�1���6mdC���놃�c3T�yZP֙��D��]Cfޙ�K��Y�*y�l�JS���"n2	(�v���eߞ�LQ�o�&�]�审���|r��2���ǳ��R^C����""���_����{�㳆Z|���T��ZͿYJ�6)��7'%o=/^�x�bܘ^k'F�v��Ʉ���cQ4I��9&Fc^�ڔ�����c]��Vt;��{n��YO:���M�j�D7 ��'�]�q&�.��ո������c���u��W8�R8��O���>P&�YZgvY�f{n.�\溽�u�Q��ņVdi;"kw)�3X5h��y�0+d8IpH�.IuVp�?Y~��4���u�X�s|�7���o<s�x/5z�łx;�^�opb~(�!b6R�4�w�/%WuzfЬ����X7H�錶Ҧ%�+n��56Nu����E��)�-'����˟v��7�Ө�7��IB�g0r��ŵ���3���ܧ�βc��K�!����\5D0؄��pE3Gv�\�=uJ���'@��w�Ԫ�"MyP�L1yd�j�'yT�=�с7:^M\1�#iHBM�2�{yf�U�nN�*�P�d1#��.ݶ��K����{s��o�W^�OK�����P���XQ�ۮ����m�q�Z�k��p�8^��4��]:�v���3ìUo���~~����\On�~^�|�F�J��N�U,��-t�re^]��#��?F�ώn�j*�M'�Y4{�[�D��d�r(p���������i�ܨ�G�hm�^����i9�I����=�kK�3z�<vc��m��[���+���S�%��W�tˁ�Ò �rDl�}�c�o&^m���/'M}���ȧ ���f9mƟ�z����l�V��@��(�w�����@�G`;�7�gLa�r������O~���%��&��,�t�vKT��YK/�A%� ��0��t�m,��Qݸ�0�q�`�r�[�i����Y�+�������S<�P�h3�#" É�]�I�z{r�j�f����C<G8���;e�Z1��pF�e9�;UD׷Vo��}�.	5���٩���QYJ��q�����k�2���퍇E�(�d)��/iȻ�+�}u��&�C��尿2�yܙ&t�2��m�.j���8u�H5MF
.���~��^�گ�<�kI��]�\�|s�&�@�/x.��s�tM^�4[��b%H�^v�i^��p�bҸ�n�^7�hU�g�/���/�rSMn+�.~�Y������`��%2��|�o������]��g������,ي�۞�H�~�6�5�jH��="�V��Y!d��;�'�R=��h���!�._�2��nçeзg9m�v���<�+�[���MS��lv}��̊E$DH�"A"�1�v��x�����b���=��Ͷ����!�ڡ�������C��]*!�cp7m
r�����Q�� ��ǳ��8M�q�u��n8Y�n��hַnQU�˻v��b�y#u�ѥ�tv(sts���v�۷^]��Ѩ:�<w��m��lC������gd������=N���oZ[W=[�pu�"\WS�2�����pы��'y�ӳ��b���9���c�];�,e���/9=��n4�����j�q\U9��#��K@�b��f#6.+b�����{�6����z�e{j��G<!�(
��v�cj�xùO�f��^��[��qի�zzCs3��/Z��h���{�!VQ�u�
A8$H$ͻ�ۥs��r��S킲u��|�,lv�}k�ݗ�q�z�~*����J8ӑ�^��w��/p5�n���۩=e�Ejk�>��]�b߭��}���="RRj�`��p9$te�zw����`�m#կk�u�A���DgDG;^��bzzA�Gڭ�>�{��4�/�!�,�z'#��6��s�O
�i�86�3ͳ�q��\��L��MHc0�R��T��`��F�>�N�}�Vobe����rOV���Cَ^�7W�a�`�����Å$
����3��3��2�g�i]�ܦ=f��9����,��zsn���)[�ӫ҂n��v3v@�*�F|R�@�w�v�fNf�WU��'_���^��>�IX��Z]$U($�K��gл��1	�<��a�WyV�u���D֛w�����g#�r��R��=�X�f�I����&K�
�i��|�W���rt�K�&��Ž�қ�X�S4%��ֳ=�����8AC#�B����~w]��:��O,D�~�&���{���I{�J�z�B/R+%�ۃ~x���n��Zݮ^�;���a�z��=qM�Mv�<F�͍WKz�d��{��h��v{�
M~���v��Vy�D��ҷ��Sg�um]��9�u^�	�TO�q♞�f{�'��{���*��O�[B��h�Q;q��\��g{���x�����锐���1"�G�Zꓶ��T�%*Vk��7����aŝ��ww��u��Gj����rh]�W��`w�ג�R��g\1H�ڃ����іem���������GH���K�+p��Ju/��ˍ��[�'�pu�I�D� qDdPfh�6���G�1�-�i3�w��3!v�۵�	͔�q�f�A�7ӧI��`h�KqH��#{�=^��F�e �8�D.�A������9`m�f�M���0����<-�+�ZG��!���yp(c���\n�k)t���$�g�\k�{�{mٸ��	�!���r>������m����ZT��r{;�wa}#�ַ�b���<�H�H��	���=b�n��%8=�6���8!H���V1��y�{�Y�nP�b,-QL�<*�B(��jE����S�n���tr���J�h1�iI���cn�)m�$��c��'љ#@�%�,gw�y򄴁��I��\^�|s�����+T1m�9��o���
�C�j�jJ�݅�ô�)�Sy���Ǣ�^7Ǌ��m�CS'��Wݜzj���b��.gm���ǳ6���Ӳ��p� F1.(ӓ�.�|�X:�f`�C�YTS��.Y9&f�%�J��F�'1y���Fc���z{O�I�r��IĽe^}=����R:�ӵ�� �=8<Ӹ��i�ߜ��nn�3��k�O���]g>C�O���BF{w�R��9N_�>v���0A#e)M�L��y����/*�}3�N{�y�
��=M�ՆBoc��aĉ8d����i�U=��>�h����Ow�2	7qС����t���y���C�x�n���'�SٟZ����:���2�>��\����Z��M=o=��ܲ5	M�nrf��>���[�ϰ�.�7��]�ܾ0�W#4�{�	��1�b��X����m���zT��)slk:��V)����^
Y�/����[Yb����W&��ѫa�2'�,��%^B���q8i���u�Ek�2�<%d9m��f�ѳ4�������t�wl�T�ǳM���SVd��)��Ý�C��
��s�W%W�SE�ͦ[a���R�9{�ː�m���o[�;k�l.���K`��L;�k&񦌧{2��Do�fa��8Nْ�9��+xe��f:xM�e5J簾�<y�vm5>(=VMq�7I��*�rc�Gy�<՝ʢ�I�9̏�=|�e�������"�A������8N�z>��^.�85���ㅽyIWu"���C��:�y+`$E�bO��7F��u��$�pd,KD����W�㼃n���m4]��2�yV)i��zd:�#���yr����E�Xf�LZ��8Wh��w�{�HDýԘ}��gv7�QW�sW�a��Oe0�Na��9�,x�.�BG)�h��C��2+�%���<�8wl��1�wMC��|��śŭ����)1Һ��Ոɹ�+:�M9��X��u�.�3ru�6��7������y�ؙm$�q���ĐvF�!�@NTt7�0iS7�h���S��VkޛQ���V�ɸ��;�9<�� |�@���i[���یv9�s��gZ�܃�6�7����/�SN��}�����5S�;���e����'��&잺=��v��9|��->�;[��I�k!o\/��z#���$V���7�'X0̐!VZEw9�:�N+��z��)Y]`SIR�EJ��{Z^ �K�;dbHJ���7g�����8���h�=���nˋ��
m��;��� ��;�j�z[�����9�-�S8^x͝و;Y�殅8 N��i������8�;��F��k6�nۖ�<�ز��Z[�5�m�k�ҋ�t���ҝ\p�#�;U.�v�g�dݻb�w'k�n�<��� ϭ=����M��lY�Z�b1�y㋺�<�Hcgqڷj�݃U����gy�:�%��i�$H��]�lu�<xٶyay:���J�����.N��r*΢1m�Vϝt*d�8��&p=��=����)�u���B�y܆�:l����%���I���{W:��v&8�`��I�4��s���.z<Nwm{6���m'��,���w/d�z1���aY���n|�	��+>^�S��n���L�{�N6�v۲�"�3\wL��Xӕ��/�<u�v0[�j85�W��v��>y�$7&�mnP�m]�����j�Ϋ����ؓn�3�6����F�`:���v�r�;c�k��=KvU�y�c�q�ms���^m`ь\5�}Bov��랣X�w�t%����(W3���+���ۉ��Y㮶�cSue;q�� qݫ����뉭�85��sصe��\�{&��g��ٗ�=k�;��q�=���k�F+��q���n�k��غ��Ƚ�+�{,$�xӹ�\6áI�7Ou��h箻xS�B��UD�qχ��nz��#�M��C�GF�6c�2v�#��G����E)�B�Kk������1ï�.|��sSp�X�"�:�n�u���.��so<�·'���y1�e�-�.�.&�C�74n��O�����n;dg��\�<�睃`���X"���7Fɺ�]�o$anxe�e�v.��� u�ԣr��V�*m�ƶ�����v�٬k d�o(
񧵖�1/nݚ��2=DX�v�g�nR9��]ηkI�]�^��:s���v��;��[������;'S��!r�=�9��.���m���G����ư6X3GB�����u�tc=����c�g��ʜv7e��;sB��=��r����u/���i���Z��V{�@���\T�3��1k���u��.zq�Y!]�1Xui�O
�j�Y�9˹�3���|7��ts�9��	�ӺH���@0K��yvP����({/Y��`��(�ݲ\[d(��7=3n+��]�mӭ<�ʘuF��M��.9v�c��ݼm�'�V.|�t�n2�.�M6Ŷw��^Q�����#Q�W]~W����=��+��:>��y4��;��o�tl�8<ڞ	�C�@JQAqw����5s1�n��S���Y�wY�ȴ�Z�cK\��Ow��lK#֥7-��,q۰�jFS&2������nU�{TT	ký]OR�cЫ`�;�%��]m����e�<���'�B\���a�P ���0��]~Uy��XW�8��ם�}��*��fe�"�~�l�a6���/є"Ё�P���L��(�|뮤zm�p;'��^{+�v}�;5_#I �@�y\�;�ĝL�b]{\�uNw/d:ʛ���v���������+���^��n�Qmm�Y��釽�!%��o����%-���R}޲!YX�#�aso%{_]e:��f1O���H�	L��V跦�����>�Ǹ��_��(M`y�G���`j[(�\�v9�ml�r��)��2�G�ک3�f�K��|�8 壥M��%'�ԯw3�&{�.#;g��+^���w=�@=��\wU��	"�0)�3wM�=�6餃>��8��v�H>�[3��������Y���KBv��C���%"=޿5�Rڲo���c�z���LNlU�UWn(�l[�:��n���+����[MjD�Ƃԑ��ۂ�Y[�Z�rAwf��Ԓ��z��/��E-��ܗ�k�{u�4f��������P�{PH�0��0A2�Uv�ù��e�Hq]sͤ�ܦ�q�Tq�V�.��9
�dN�9�]��I��ݮ(�Y��O�M���ג�f�yZ�#I"��IA���)'��l��1%�Ɯ9��L#MB:���u���{�v��\8����Bp�����v�J��{H�H�'���zkarT�_5���F��W�r'2$A6��B6A�q$wwQ|P���H�����1l�g��a8L7s�Pkz�c��k��X����0�_ү`�UsK6�6ڬ;toI#��a��Vr����wܖTS��nq�ė���u'���Վ�AGKe0[},��"i�f���yr�D�Pƚ�:~da�6w9�&8k�d[��/ix�nW�,���J��||����I~�a�_��0��v�RyYrr�7qX��`�%�D�#�y�.�(���a�Z��*�}�;g�D-UgB>1W����+�C�0�#��u ��#��$'��^�:�ID�Tt_�t����(��8���DN"q�G\&�zy��.ޥэ�]di�`gZ�{qj;T�m�f	rx}�>�H��b�~���t�5�'�a�C���b�]31i��1��̄�E�#Y�n�Gq8r�f6u�?B4�6G{?�� $�2䊾�Ə��F�/��Qlڶ�sc�^����D:oi�S�D���'H����F#
(��Jβ�eV�E�+�0�Ȉ?~���Ԅ8��JG��8���C<�e�2d��Gݴ���o"���ON�٨>�1k/az�5K��z]i��F��7�s��p��m4��92������i���壈GVw�D#�l�!�7q��V8�$�t������I뾁�Cb��a�O�RŘt�*X-*D�K�v���,^�6s��\���]g:�)h(�EB�����n!����z�!n�=.���Ф+Ij�/��"f@�2%")8���f%�U0���i�4}cXI썷��Hs0,3MK���E�E7Y�i�(�[�"��u�p�A}`uOp�S{<����������γ��nJ����;��j�q�qv�^�Ż��p\�-%�"K��"8�N�!g
#1�E�j��^��(����y�3�/26����՜ӄV26�"0�j>���G	d�#��q�i�E��ҾÈ��γ�=O{��%*qg������A���0�S�P��Ir,�yF��N������k��|�ȝ����A�`��Pg��rF���*p�F���&�:ˈ�(�����#Y��k
0A�w���#��#��K�����J���d{�� �2���NIC�{���k;C7��ǻȎWH�>>�������v"���MǔG2l�.E�9k������s�6�Q�N�"���6�o�Ȁ�2DiH��h�;���?:{�F������]�E纔�+��g���)�d!gХ�[���:��e0���P
}ҟk�>>����<�2h����c���}�XB��.8�뤹��__o8`��!��Uqv� �ns�:c��u��H6⏻o8��A�KK%���Dr����K�v�$��A��.�=J���s:�Tڪ�.������xGu��qܘ�[3¶va�1ܧ:���68��;�� �s^9�ݣXݶ�t�z���ن�ێ6]�\�zsH�7Y��䨆���h�\����v]9���{݈૶�6�V{r����rH���B�&v��;NW�oe�J��g�n���\'nz�j#�g��ri��s�C;�#jMm�F�V���3�q��qV�c�Y�1��H�^~�<s?1�]ז��ϰ�}��#z��ނ,�3,1WS!�8��u�tC�"���t���v�M=��e��e�R9u�0փ��2�=U���k)ds7S�i�D&�K��ay��!�QD>��Bq�WN�v�5Wc/a$p`"�bwO>DQ�i��D����4���|bC��aӞ�ea�'�D�yN�:G.��\?�4<ʶk��oH�!�o%�_B�K#�O�0]6h"����|O��F�g�d]���(Q�,+�Gk����,�ۮ(��9.�9��8�0�w���p�����HV����������J.�5$v4��GMY�Ϟ�ih��,�~(g��4WBt�U4k&��ÂD�~"O�X`�O������oE��a�6����c��8�hF�jBP�� �z�sX���6͡���.!�㛮7k�5ͮ���)un�qma���G�X�_os��M�jo,br+����F�"0��S�����9�S��/�8�3�#u��ͬ^Æ����=�Ӊ��l&�PH��f���C��'��IO��f��
���a��W{�CA$Fr�F��'���<Ҥ+1L�jfc��`gtL�o�H���Y�ɏB߬Q�<���wt�,�J4}��u\s'6p�/�0�>~��[�q�{7��T�,�o�&��I9F���$RE���n��Yy��v4�(�5}d[����#��� qM����=,U�Gޟ�!�kT�J�ٞ�߼cq�����5!��0�jp1�+�=����3oz��:��}�I�aّL�bm�T��Q��ˉ:D�#H8=K��Vd��5��'{�o��2D\����&Yh���#��ҡ
8�D*�HL��p������l�l�(Q��6E[QD��sJ�E�{
4Q��X[{�s&sq�@�t�v�_����1�oF�.�C\��\u�r:��X玫i�nr��*�
?�M24���?L���,�څ����1�ǽ
�+=8C0�߾�>�S��}
����5�#���f.��[O�����"��]�$D@�F7r2�D5����>qB�>��mČ#oI	���aq�w\� ���f�8E���̦�iF$�VT����8~���9�!HЍI�;~di�B�W^�K�N#����cmt!��T�s6u�4<�4��bdi��3���p`sI�N�{o/���N�L�p{h�o��I���/:��.�8b��'v���
�Yv(L*�#���p9���C�B������G��|�Q�"����HH
q��(����\}�bl�m�>kݶB��p�7��7F]�s�G�D]=�[�mo6�q�G]K
f��6��ba�O0zoY�k"���al\%��1�L#:W�"�����!��a'�{[/ND��V���dK2F�I��N5�6_)��ܺ�f��p�2��!`Z����;�ļ#�Yq۞��K����`�#�ܽ��v����`��5"3pH*E��Y���3��{�;p�#Ma����c�|p�>SШ�޸`$�#�2la�`H���>���_"C�Z{����$��(!N)�8lt��.�L������4����;�7g��|��Y�L9_S �G�F�;]4�Y��3���U�x���+�&�p£��Oǆ��0�9�%����4՜����E֞�#�j��_�t�>��lI�O�	�=�|����WHᩓ��")!0Ƥ-I��.ۘ����g`2Ñ57̽D#����oT'����l.7�sdI������~��c]ͦQ:�7�l�6�Q���������oi��wo���%��&�)��1]d�Aܥ4adCCE�ba��$پeJ�>�aD9D�+G͟��"�&ك>�|�����{҅�!�O�^���A�m�����"#��sdw+↾������C�fE\Gg�,��2y��鶏F���D���\.� �u�t�V�#����#�=���sۮb�p����ظ�nu�MM9#���#��l�����I�$�&cz�oI�l>�ȧXA�{=��%�#�VYDb����4�j��(����C��p����F�`�WI���n	�*��iVK���y� �U���*�A��|���1�!�Fg��:jq!6��z�o�ΑKY��A�������ø!��M�i�nIb����I;�����oam��e����`��(e��Ŗ��Q���j���$�2,X�g$�4ɍ���a�ӌ'���n	Re�n��b�_��HWra���b'���k��Hy��;Mjz�zB�x��afUu����!�Cx��{(ݹ�r+��#�m�9�_=�Υ�A %#!QHpi�G"u2�^�:[�B%�y�۶*�i�a��.p�31u�^��E���wK���f#.l��7H��
�F�D��z1M5P\c���W^3(#��AR��*�&� `R��X"_S�j�w\vn:3j�BO��i�y�oa4�{DV�Z�����w6Qj��7�l���gz;:����n�v�oh�֔��M�sIbˑR���8��h��j�m*�[<k�X؄]��6�=Y.�G�]�v������]�����,�����G�;��`��0p�8W[��8w���wR꓉��by���s�v���n6;j�B�g���0�bx#N荎//:D�9�N8��l]6�� ���<&�nn5�8�v\�vv���o�g�]�ͮl�NI��ㆽ�Cc��c��'�|��磇h^�a$B�Y����(F�6cd'Ԩ�ͧ:����tˤ0������is�_�	��RqX�.�Ս���؆�i�64јɅH�S4�~�C�^�籽��-o(C ���`����Ͻ.����pA�Ʊ�3�Y�'���S�S`�F7�Dy^,ٯf���~84�	κ�̙�����������;m�ܫd3[�0����y]t���Ǥp׾=7�*P�#"�x�,�0E
w_1�/a�y��>�Ə��G��6��4}rã�����K��0,э˰��a�T��g���c�Y�1�\"��}��7Ȳ����c$"z����!dD��y�cg��vj���k�a��{�g㦬���|��}�](��<77a,E|�M�3���A���uf;tv��p�����.�ͳ'ٻ*�Wt�u�7=5��������62β���G�D�ǣs�}!�VG�_��e����®��]#Mg�nu`�[hu��)�~'W�\i8)�"ϸ����B��s��{`��=�'��yeOu���T��l��W���tf���)�^���|(c��۪6(Z�jT4����D�};�TUM4�]<�.��@��Q��R��M�Ʒ��?EDa؄����lc���_��]�q����D�{��O��_���c�ĤN�XF�8Gp��,�:p���Y}�j��:�	y]��>53�ש8�����"O��oUw[���F[1'}?#�d��(0B����Mn�λF���+�D�1E�#e���Cv���{�6+Al!��/��`�����edq�q�:�����l��b"�Ir,C�d�,��=[��
8ͦ��XQ���1�,5�A	oAjȏ{���-?5�3��O|�N��4�y�}����lZ���0QNIq;m��:�q��[��Iܓ�f��&�vcu�GQ����0�0A0�da�$?��Y|��?E|*�&C�z�Ǯ�^�a$a�.�=�T���~_"N&�}�j�כj��<Qx��p���¹���dMF�M7�#1Yt�"e{�K����}D���F�!'�!9svޒ�_4"�Ä4��v��6|�Jpc��,֞��~D.�ƦJ��
H��xI���ݘ�>�2�a��F�W��T����-�=�&$���ֶCű��wpb�8��.��Yt8a'{z��;˗ձ9	�9Sh]X�sܩ[W�I|]{���a۷)#Sv<|L˸SY
܎(��B.ܗ�&�Fo��_\���%�J�H�*�����|.��9�˟#���ƇC�ȉQR)���9!�I��39�Mŕh�rbCM^#��j5(��s:���=X5�]�6��f�g�e'(�T�}�Eu�6GO�a�nUˣ���jA�8T�n���L��s��P̸Z�e9��+��U����P���Ю#�62V�8��V������LfI�s�NL�B�v${��r�|�-$�����՜f�c����L��S+'<�
��dN��)�pa8��n�A\cu6QB�9�#���2�흯S�4'd �uV���Z�U����6T]��7/ o�g>C�b�Y	QZ}���.]�A��aHKM�O0H�$D1��v�/tb�}���l_=m4�{����Nk���.	zg̅�db��ʸc�˚��Dʜ��S��)GGd8)n�N�2�y����.#��͖�={_)M�3�o�d񾼪��7�G|�VkZ*����#5*$�Wݠ6pȋ-������+�;��V�{}I��a�A*���N�.��u�2-�%�[��\��X�f��ڝ�0^;�$��+/)�Y���c�����st��S{n�WuL{P�Y8uh�U���������v_\�X��h$�>���\�wy���v%�����v���2�����A��^�����!�V/�����4ۊ2SM����$��Y�0��]�?9�4Bx+ƽ��U��iF�qA�6�F�M��[>W]"��g`�n�(�}�kͯ}���KCHG��oĮ��J��)$p��6Q���2�9г"�QqxR�Q��a�oj�zH��-dV��!9��a�Yr��2�0�zY�G��{�D��Z�F�8�0�L�2!�Q����g֛�;֭=��[v-�Ovvɸ=n�a:!!# QH~5dt���y������0A�Fm�ة��>�a0�L�6Ibu�czm-�,�e��8C�H����H�p3#I�#�e|q��\Є/��u=(a�<4q�<��0x���!��aPDո�(E#�Z摇�q���d>�s$F��^x��{x���H��7�"2��"(�ᡄO�#ڽhQ��ʩ�9�����gi8k~N�z�j�v����>�q1���a
<Ea��;�����|�u�Ⱦ�d&R8Ć�Y�^�r���H}1�����t�ql ���{8�Dk�'&��̣"��1���\��c6k�d�k�����]Au`��%RwI=���1��S���)͊�Z���.��8ȫa]�V��[r��p�Z�t֌�vAǹKt��T��F�"/��������!�$	r<F��醰�Y'�L�?T+��PD��9
�Gg.��XF�d0x�ZW��h�"e��S���VNA�D��\�.���:N��.2D�!���Π��A�Ӱe�ۨ�<9��a�Y�uu�p�����	!
�]�Ն�Wǆ�*�fl,�2l�g[!ghf:t�0I�[Ά-��b10�]AP����h�!|^#���|#H<U�PX�>"�Z���.��I�4���Ӥa�῍/]��FV�:�[�<�EϺ.�{�\�������U,"N%���$�]Ѷ�rRC��$������
�ȝچ@`��S�E��qY�~c�0�s�<p�)�)����L}��Ҏq1��<��"����G�O���,U�N���~%u��B)$
D�H�!Ӓ,�Fj��g��x�=S�i}DA�d�d(�
4|��ے�"K#3(>��%�z���͝>�a���`���&	�!q�_q�XG((�jQ�,�aG1�;?���=�pQ�ʡW�����v��n7�a��=l��!���a},��~x#�9ԟ����N%�j�uY�,�}]�R��Z�Y9�R=�l�8-V����´��>�"��_Y�pgU�4��t��I���[÷�,ڧ�c�If�/]���\���K�v���ɛ�;۔��M����<���͓�;N:���v�Hnۓt�;��NoJm�Y竹p�8x�٠J�U#C�ˮʭ��Vu`p�u�%Ut8���;�<�3{Is	MʝqW�#�=�;�U'=7-��ö:�(�����zN��Om�4�Lq��ݹz�a��<�s�c�h�`�l�Ԇ�C�^��!��GR�1qu��NRQ�B܆)���XB5do��l|f���D�����,aƈ����3�'~�����Y!�&Cv?�+�Pt�l!�Q$W{�-���#�0���_�!�sdQ�v�88�۳1�{����7Lb�2�[	>�FJ�2*5�q��E�&y�we���bΖ9,I��6F/{��8k�}��0�a�c�Dڑ��� �U��;��+��5��Y�s屢��=�Y��h�<kmM�u�,�i{�)�����K1�(��;>�ȡc[TQ�T�et��a����YG�3�1��\����D[y��%y[<q��52{�aj�#�,�G��"E����
��K�7�U�W����:[<���'!jI,n�Ӥt��������Z��O_G�	ZVF�CO�3Kah�ػ�Cq��.F��O����d0�%�""��5�8=,"ʂG I����`T����Y���c.�c��6d���R�nC����ue��D��΅�"(�[NOt/`!���|�n���%MM�1�G��"gi�^#HBq֑���&��	N$Z�آ$Q�B"�wY8m��v��T�¤7�:J�o𱊱mi��o�V��6爫e4;����\�u�EXз�V��B�����J�o��őt oc1)�"Rζ���&���ا��P��A�鼞;]G����ul6�r��Yx����L��#��
�)$�����Da}O[Ѕ�D�6}$7u�e��p�@5S�18��Z`��4�E��D�G_>�\#M��Zzxk�c�Q,8\JHQ�EcF�-ag���ǈ33�r�{��r��k%����t0���ͳ�Y�W���0�a�&��M_�+�W��i�a��FH�>���nI��p���6Ja�S�,��H�oQ�V���	"0Nj��ir"H��o,��oC��Fuu2�,�xY�<�}tT=VsV�ߎ??���?�l��7�dd�ƻ]�g�f��Qt,Cۭ`��	q'�}��g��d�m�1Q��\���0����Oߥ֞���ْ��LoB��4l�]�抲�5lx>)����}QU�"�E8���V� R8#���A��5��-��t���EG�P��6��>��*�Hda��a����Pa� d�ճ�x���?r>�-w�F��u�&�M!.	��z��dI��ϰ���}�5�h�Rݯ˜���37kp=��"�[��y����EK���;��Si�ٗ��O3[x�ѵn��"�	X[�%ɥa}�p���}u���uޣ����$Y�$�'za��vʓ��l�����dq)}�ȑ0����EC՞�T�l٬i߈ԟ��s��X�q`��T����ۚ�H�h�PM�����#h�m�x���KЪ*��2ہHa���'�C[�ndp�(���dI2;�O���oa[�{��3��L���0x�T�����Ym!#H�4��ۡ��t��dB�צ 9�>K�����A�4��Yy���i�od8���{Sz�UƜ��k+��i�u��q�B���ҵp��F,�r?},i�#�U�l0�_�"H�d"���W5�S&4����6���\Y�Oa9F��ƳO�ϔ���M�R����eZz,!Æ����:��q�f�����A���1Mg��&�oB�GH�aJ�s���ҙ�|{���|Ѥa���w�	�2c��D�&�>�Ç�hQ��P�'����\�w`^2-đm(r�!��������7M��Q��x�>{�P�<l��\�V��n)#17g�Bϑi ��q 8m�6F���s�ϰ�'X��![z�6|ɇGQ�BM�
>�h({�c|F��'�t���y�̺�j*��n󞝽��f�ơ�ˆ�zk/�[C���<U�tp0Wa��Z�o3�ŕD������	�O���V�q
sp��Қ�ch�\l0�rm�3$m��XI�\"�W�=ᱦ�k�F2,�Cf���3Й5�9��>���l�-0Ƀd^�\$��!�p�:G��G�[@0�&W�(�J��9�mSv����;:��.�ɣ���r�E�5S×�=;p�i]��}���v�!Z�4�u��n�����"� �g_#�.`�v��E�oD�"t�C1�S.0�4Goc��C<!�G$U��0���(a�����[���ut�FB>ㇵfB�>��(�E�+�&��8C8G��?+� ���hi��*��ya��l�Pm4�2Ց���K�,��ĳG)C�MY��t�ٹ�
i��>�k35���C�b�G���K�a��9�%ĳ�@��!l�"�K:Q۟�:kE�a���ߞ�#H�a��f��0�܁G�#[�����^��>8G|>���e�鑤&�#:�����y�L�k�BC��jD�n"�'Mag�o�WZ{��>��뺻��>]����Q�_�z]t�5�@jw�s��"CP�"_���d>�0���X7�)t�maҞ��p�ҩK��Tj�Flm�+Eʓ�N�%��]�_Q�3j髾�6<�v�`�%���s*��fF�˴&[֒$���&z��O4����m����7Km��g�6��=�9۫���t6�{A�m��n48{.�$�C�e�����hE��>3¶r���n��H����<y�4x���c�[n%�u�70�{m�8:�l�K@l��g�5$��ok�Z�D��yl:0�-�����Omu�J(y�\�n�9�wVwmS�F*�u�
��t����S/G$v3��N���=<�vX�s�&��F��k)��l��s>fݒ�����$>�f�D5���c��0��h�Փ̽�"(���FB�4���rX��C�{����lU�{ ��Y�D $AA5"��e#OH�/.��eM^�@�R�!�y�5:���=�c�����d3�?�7�u�0�CH�O����<~c��Y�>7��߉�D�p��:|?w��?��C"����oZ�\`�0�%t��Ib4\�B-�fE��&VwB�0��o�6h�����	m�pI$�|�b$i�2���<s�[���4SO��Q��t���(+oI|�\]Os�'��!�̉�^��;��p�GY��_�F�NBʂnI<D?w[�\�ߕ$�:z��Fy�	��~!�4laڋJ��şi�F���p�[q&��Q�+�X�N0��5�a�-�xf|N�$�g�A	8�r�֮y
6l�3d�m�k�4��Mu�;�����DH�@�*IE�"��0�Dr�\�}\ݭfy>�D�d:1������^��	DU��Y�&t�8�`a�4�oj�äq�B��D�=��\�.4�bA
�J�k����o�-��+����{���;��X
d0E`�E�̗Æ��$�ۃ+K	
HZ13m]�ACf3a���T�Sk��M\qi%a��ežC�3��N�*p���0�"(]�l�z�I�,u�Aczb4�>D*��ML0es-����Yڏ�dOH\MO�q6�Q�C�?!�ȅ���+�rYaR`�;̂so�K[->H��MS[��).�^�$����jWt(��8xF��F_�3�&9`�lHn��4E�S�G�E���,-���C-���V�Gos�V�#�g�C���a�M����zO��ڲ��"��G�x��m�i����Yn*~�0�!$mN>��'ʘ"�/226m��S�#1�Dqd��\da�$�'��z�5ǈ�vbr��{��5
g��PZm���F�K<������=��"�8��b9,����j�C�;C�6��S��n�f(�1�����d(�s�"���0j�l�}�!��g�vg>V/ �a�nR�֟��.�~<5�t�1����@�MQ	�K����2i"ΐ�e��i���5wM�Wnl7�Y�`г
�8�E��'�^as��!�#H6��x�%�S��5>'��Fȝ�ѱƣ���)���p���	>�U��0��Hn���|��Di\�ܻ�lt�۩��I���Ǜi~�2�8l�jjEN59��ECaV!�R�0-�,]�4BKO-��Ji$�*�.�J[-$F��
b����fB(��t�"��oY}-^B�M��,(���������bW<Q_cϴɓ�!��S ��c����ܢ�XO�I�"!�@`��JϾWM,CH`ߐ���ቸɂBSf	���yaz,��w�<��#�ߟ�[v-�w���l�W���,t��D�������5����eY����p�}}?4O�p0���"���1�<G��:�p����M���]����
�\v'W�IS,DdP�"��4�G��G=�wL�&G�D�C��2}$Q�*7�l�ԟ
��4�Eu�	3u��2|>�,�l��>�߬�b6��Q�+��a'O&MV�_:ő0�v%PDBoYy�*�����sܲ���<p����S,����l2($��7�~��A�u��>)�	�ӊƑ���XF?��u�a���!�s;�\?Oa�Y�\DߍH��0�]ikHڵV�~�`hpՑ7�� TE4�iB8r�����4a`v�~��� �*�="����oA��F}��p�s�I��������C��j�g[�,�����X��a=t�r���v5B��!cd�0�Y��nc�Oz�Р�Q^l����xl�|4�Fu���]E�H�����֚�F��@�[F2\�Ht,�H�|���4F2}x�h����,"��ƴ�Q�P���Q}$gR�^� �0�[�ʤ���B�}Dt&���q�����H�q	$)�A��Z����lk���g>���wnF�z
ڕIzķ��QD�d�Vk�C�]Ϳ/��0C��tE�6�����0p�����t#=!��f�#O����L�,v7%x�j}#� �#�\����i�0����Ӟ������2
�k�B�����Vޒ��D�9��E:D�H~�Ns~V:k�o64c�!O�U��v�?(#0(ɒR�K�;��]�la�.O��8#Ma�}�j�a�[3<�S0{h�2t�J���ЁaFΚ!}{��:AJ����ٰ�!�(�i�Ԇ���Y��뾧tamBC�SxN��KtH�}��i�,�y�Q�0���oba1UЄ�"�D��*�v�lbd-��g:�[g�1x����(kЙ`�$	�!ψ�4�����f�ȳXe�$�����j��_"��AIsX�EM�L:�dS��Z�!�_i�l����_R�?*�N��	�Y8.�9Y�tWw�k�����WF願���&B{;��Iutĵ%�٘�2&XW��f��nț���8�g,M�|���Uԃ�Ks�=������vR�#�l�s�M@�ܢ��40`�ȲD��'��mf�L$-'�`���J�,K�x�f坏��8��PL{7�Ȋ���S���8^� �X�f�x���8��}��C��)f��¡�q;��]j>��v�]�f�!���q+�̗9��>���!Z-�T��W^"m��$嵂�n�s]l�:�G�Df��D�����5'��K�9�n1[IO�Tʉ��$��KK/�C�mm�w�%d�t}�����̱W6�X�����H��RKC�:�&�-۾����m�*#e����= ���)y w�ಱЅ76��AG!���`%���
MjgfI��~���Yw����I���5�ŀ����
Wpr �w/p�[�A��s��z�m��:U����N�n���v�Il��o�k�!��6�����-�0���s)G�wiS��w{��>|Nb}w�*ܗ����o�ؙ�Mβ��_(�Ҿ/��)Uh���U���g�E���>�w>K+`�c��[X^[��UK"/&�T"��^\^H��b�`i�j�}:�pq���;@��h�ܟTY�)��*�]7�6�^w��b�L����0�ޅ�e�'g����i�����n����]w4��Y��#:7��u�B�K	f�I5�۔�b͸�~����}���%@VPU���Fh�����vtc�g>bm��Vn���d�`=Sj��ol6꩝q`0�o�8��r�S�:��{s�q6p�U��m�2�h �-��U�����\�vz�=v�k;B�ۭ�l��q���$.�۱�yk�O[��z�]fz�m�\i牮C<��;u'^C��Z���p�=�^)8:��r�gu��#'��qÇ��n�[���;:��\���ˢM�N�`��e��8ۻ^d���]��˸�\8�`��g�pu��H�[!�c���Oc3��\�x������h�z.����oSn�&�5��C�������+�յ�\���M��睏en|Ks����ڨ���v*�G�շ[�u�C�y+ ���Ea�$(�չ�떵�����l�uS^yv�P3�`�v9��S�l��g�G�Փ�ln���v�-]�rer����wk={f
�d�6�#�v�՝��[[;�GBۉ;N�X;v�qub[����/=�������xvYg>u\L�c�>6y�8M7v��ϛ�:�
q���J���gZ�ntF��N��g>z�=��7Oa��Iպ7W1nz���pA�;]1۶:s�A�a�D\���R��F�	�A�����m�����+j�r��zť�7/WSۻnlY�d�+\�'@t�6*���Hv�7S�t�۲��=�k���ٙ�LL&-uk+Ai�jA=��:��y�v��󖞜�[k]V�_v�ދW>QM��C�'� �3B�J$x�ꇷY��&�;nX{3�j��pdv��z̽����ܚ�vz�\��wbw㵋m�//cuΙ]���3�u���`9�=vìsx�lnS�7l{\<9y�Bn��;8�gv�ε����kq��k�5��u���h[b�uv-���o`�	�g�5v2��8���b{�D�"��\k3���ۂ2��v��q��9��lAlS�ݱ�kf[�6�vi�g��L�����ku���#�%�[�����[��]7Y�;p6^���6�(q鍇E��LS]P�p��r���ڣ��(x^74#\���Ïg�en�j8�ut��Z�k���n�=U�yp�[���X��7^�l�3��]�S��i�x�U�=��mr�7n![����A1�9�	rZ�!�0On�=�p���mf��i�����;��W�� �N������1�{T=ͺ�ǫwZ���Tx܃��m��ay�O;m�q���D��U��7<vˮ\	ֲ��[۳�x3K)͵2qڻv2o'�����.&*��p�H��ae��:j��mC��K�|��_PÝ�WK���#��m��F�ϑ���q}Dv3q7���FY��FH`;����.��l�WO�Zг]RP�Q���Ʃ뎑��E�<����$ك'�r�]̆�P6FvliU]
��!����|���FUg1��ho4�R���U�:t�#>���r�E��P��K������gA�k��kRj�^��[}��>��6û�[�nA1!���O�\5��#��F��k��9�!VI��-_�J�y#I!4-�@�zbQ�|��f�:���ִ�"�γۓ�4�rQh��ƈ�g"H}5��Y{n4Q�(�L| �c���7nQ��ރɸ��0��l�5�_�>�]�4�jGn����ѩ[��JJ��) @�R6�)�y�d�Z������ZN�r]���ϳF�+B��uɳ�I�ç���"o�;(�xF���.�z�5>�$���@��l�@eN.[��Z��Du,�U�0���t��O�g�J�f2T��6;���2D���/b}i�!u6)}��fXP+��,�7�	���%f���g�ݗ�ם��:ӫ�qm�#�]��BSRpt����#�c��>����^:
�Y�,�r�RޘBM�E�AM�Q��9��2��.z��"����5�n�0�Iƣ�"�s������(�m�.r��N�"�NQad3!������Z�E��v|���a8G%]6�>��Ba"�h�aE#�:EDY~/{Ù2��8��Ǩ\E�6|�0DK�:J��_Ka����	8E���"}x�%���c�ޕ���?Yf�{��F4��@�[������#�
}��pi�0�c�=�T(}�(�4�����-Q�9Wp\y���L��?yr�9W���"<q&���p}JBs!m�X��M�R�&��W�ccr�Z��w��7]r���;p�i{�ͷ4k�a��)Hc��H���Ӷ�����x�4�0�L-�B-�%͟-a���q��pF3%�l��E�����cg�CH&���l��HqE"	�Q�2����f0��1]̅�$#���Eć�i�����B���N2r��ބ-y�C��������ä}ù]+Y~ǿ#_��}R��F��8`H��%�&���[>Dd�s�f�sY�ףe�u��K��m�~��r�F��{�sV&�"!����T��p1z����0������:��cч�_;B��*vR��>h�Xe;eL��w�W{�AZ��bt����o4��꦳�t5�W$�|��� 1���\#q����	Ō�C]y~�`��8B��|��W\�c����D��#@�r���k��c/H�ۗHDu7��j,F����)N�7��9�x��tu`^�fO����i�:�X9��C?[,;9� �GLdL]�!g��"y�o��.cu�p�l�laD@D��DE�
��!��;�c��6C[��2Y���m�j��N�u�F�3F2ˎ�]ug]��i3�=�ϵ��*�~��q��!_Y��KyРoQ'��� VNG`&]	5�lCx�����y#1���~>��J c"����0郅���މp��������
<G֒�3a>� ��wg�F�I��R�u�΅�5٣B��cx���1�܋w�A(BԚa�QG#������cC[B~A>X�dۈ4u;�.�3��tЮ4E�~@+o=�kת��ak��z^��U�%��S����	�%����#��f�OH�j_y(Mi/`D>�V65{M�6C�a'�=�ꍟS�6�R�)o:��x����9�n�������ȇ"��0�Q��0��CQ�~0)\�
y���2�5ۉ�G-:����t�0�d6��p�'4|��%�|�ӳ�Ѹ�$&C!r��#���0ҵ���#�\y�5�tYК>=��n]=B������y؞�\�i�"pEiC�O/�8h����c��؈n�D�ɮ���!�z�s� ���
���WnK]�L\���v-�ҧRXp\Tպ�B4Dc�[S���v�'��K�.5���8��<l�l��=5�d7<v�I��Kdݑ���mǝWs&5��qd:<#�{~i(��l��]i�p��8��\�Q|����I�l�Ʉ&�.sB�(a��C��M#�b��X>�a�Q�6�y�dZ1�!��H�U���Kg=���DA��D�xO�L��)�#��
�[}D#��e��v�6Tߪ�ße��s�L
S��d\�"��2'/���K���|9�|�d%0�i"�������P8����4Y�T�4�HXq��o��{��Iw�Q�-O`Bq�#�ab�f�6�P�T�9��V�4���D�f��g�K
#
)�!��G�� �{�{�~�fH�x-�%��Ψ�1�Y��8|��^I�(]��EZa�ޝ��C��i
ʲ,G�}Pwǃ�����2���n?���[M��4����|��>\�d�oNf�2Ye,=If%K�8��n�x
�rwT�*D�1#�)�Eˣr�0Mf��j�7lr\�k�� =���x^l��u�N�Cb�� �x�Rq�5T)��n1�Qئ"��bו��'m��!��-e�G�q��c��>;�lM�C�:-u��,�����y��#�u����Oc/5�f���97f�=���Bn�j��>��s�Tf��XЬ��r%���.�U��q���ۦ���ն��)�w[]��vJ��8v{<�v�͵�uc��s�5	-�]��*��ug]A���K&I>���8a�a?����`0DYd��o��a$H6D�����	��(�f!=�bGH�p��w�_�B�:ޡf�{�E�a1��R㱦����.{��+�[kt�W{ю�'+(���Qx`��}�p�D0��C 8E�mc#M[��t�T��%��8:Gۏs��InER+�Nؾ�!�c5+�d,�1�S۱`���D��0�fx���cD���d��k�+X�\��#SQ�|*�/af�Yc%�lQ#�3DJ�8K�Cc�`�7Q�g� ��5]�"�s)��z��ϳXY~`a�

)�%���~.1�o4���(�b��`�4��@B_d���7U��#�(������Ҡ���RT�L��x��GǒiBGL*��D��lT�rt8kް�L���s��R�!�Eǔc��$�
��ƌgf��E3P�}ǁ�$�q�Tn���~5�h�k:���=`�7�fd��=Kc=���U�7A�y�9͌Y��]`�F�$<,�����������N�,8r�[΅�#���+'z�6t��"��b,�`���z������,�֣'��&�̄H�4��������:/��n�і����)���p��j�Ӎ�ia�JR��O����A��eu�9M	^��_V���fFV��!�Y	�H������U������y:�	1�$�8E#aW�g�qFv��8۞�Ol0�m�ܿF�����h�g1i{��kdDK�B�rP�<l�:9Hb�l������0�2:��2��$��b�vL}P�u�VdQ� �0�,�?g��CO�Ld"r��ÊA�a6�1$��GZG/����?-#�:Ljk
y�M��ɷcU;�>|`�Z�9�1?\ �5�:Xa
��8�������6�sbt�!���#���D��%�ٞh�t(�d�=$��X$I���i#�����!�H����/��v4��/�����t$�}g�?�c�&�|>0#������H}g�E�;�si<bU�K�z.�
�Eζ�[��VRWn�Z��@��tP,���2mZp����ѓ�#�����h?�ŵd��DN0�&��111��RkiIc�},g�I����;��x^�2[�:a���-�$�8P�����4F!�/�WI��d��� 缫�d}=��Wm����VFȃQ���h��l5��O�&��`�,�+����`�I/�"������VW����20{oI��GV��j�@{��N<�e)h,��/.e,!�(u���`1�2勺����(����$�l�{\~�0�-�*��d������y5Z��"K�q�R���"���,2�����i�f����1�(�Zf2�G CpV0�1t��6X�C;Ӵ'�C��f8�""�s �c�H��W(@��Y`Ѳ2�����Mg�b���EM�w�߼l&�h'2��z���8F9�V4�"�^�X^���<�S��D"(9l!�j�A
�K
>D^j���l����.Q�JC��5��Od�����\�h�d��՚�q���+���VƸ���8��z=�7c���bY�5�����XY��=�BN7l�2�ϭ����Q�b}Do�ȧq��	�H�;���M[z���G�Y���	�HH��g��æ�uw`BI G=��=���k�I����^k��4�U�����o�}@C�I��u�a�Ȼ0��5�#�I��h��F(#rX��V~?|>��i}��$�멐�o1�'ٔ�]��N8���B�S��e�C�!8��\�&��|y�,����W��%p��j6�^4�2#Nl�=����D�-h[!da�:���瞅����E�����p;�@;7�tO
�S�e'+��t��އXGK��͖J��+iެ;r��	j��A�����u�}kd"5�i(��vՙ�������/����p��#Ǎ�(#�"Ϗڙ#=,j��E"K�w5��\��e� �a�P��!ag��gO�m�]*���;�	b�&}�Y�Mg�Xp�MY��g�Go�G1�� �٧/�.�'�ذ���F�ZƑ��ե�e�v���bu��P&uZd�dr��{�4���a�w���:o�g���8Nq^� ��%��>׮�B.���㌛��a$0�E��e@��6k����ͱ��V���!jA��$a$6j��4 ��r`����
6x��4=Ǥ�6"���SІ<~##H�⬓�K�Q5�9l�H�~�;L��̑p���ӂ՟Y��NG2I�{"��]L�$t���� ��[⎮#��
QA�s�H��(���B%����-GݤgfvȀ�2��6�X<E��i�X�~jW�Z֌4V�=�x�����8�~���ޢ0�5T�M�^�15�(�C�i���k���zk1�$>�IG��l�����{Np�"K��n��5#$0����9��Gyۥ�'�XR`��~�o�İl�9\q��洏o�͙]#��q���r�IxrU*?�*S���c��kW�޺�z>H�UG��ϵ�)\�V�ju���7+���URAIQH]�0(�P��88���Z�cl��c^�����O`^�����om��O9��;v)d��{�a�vǓ��uŻs�u>&U���
�3���w)s�	�m+˰�z�턡69�6�::z�fՆ�8X��7/]=3�#��������\��C�|��[�;\��ۯs�g��鐻9�e�+���J uF�7���q��Dl0㠥�ڴ�ɺ�I�����n��!`�I�.n[m�*�{p���,\�*>6���	:��B	�	�G������<k���`�F���)��<�
{Isg�pmms���+�H�Zg��$Y	�#Ю�8}���h�z�ˆq�E0ԅ���ᆺ�G�w9iXᝠ��*��E�"|��!Ld���&i��N>�ԅ��,�-��Ќ����'�^+!̽�8il\�F�R(�*�GC�d{�"ȧ~��"�X�QE>�e�![y�M���$~�l�B��Ʉ?f���x�,�!*����Y���8���Ç�_>%�� ���]t���}�����z:E�Sz�t���K�S������ث����g�6Xש��.�H ��`�#9>�#OK�H���z�B�&�E��8hal�7�G{�a���~-�"}�:�n�6�3Rm��a�����p�)u�O����FOO$*[Π��f��0��D⯞�E�16���*���=�`�x�wV��T6{!lm��G�8a���6�q�ϰ�8�)�#]?_Zt0��>7���]ν����I�:;(�����]۝����:a��=���{���|��3�Y�N��D��%�@����n�3�f���'�z穳�;�ނ�ތ�P�(�a.[:Ju���e8�`
j���Kh%:`,��H.;܆��n_Z��/SX8�Ap�5%i��7/9���T?�F?s�g�n���o�jl!�X�8���8𵦻�G������0��b���cP%"I �2G�Y�G�a
4F��(Ys�H�[M���ʲ*�׳D^�<F��Ad���L����#
0���e��桤-U�Waa���JXa�!n;u�ٳ�﹤#Z�p2�`$g�!{N�d|��Nj�Ab�E��� ��:x�8�"���M�9���U7[��^�x:E�f!��5��)�a�ˊ77�1�8�<�Y�u�v��a��]��:N��ָ���-YQ>��o鸌>k��B5�DY�t��«��p��$��y�g��%L�+��f�v�A��N��闎�i�]����x�C��N��M=�3���,���}���ߕ|e�>�f���]���B1D5�U�@��ޟ&:���#��a����*��4�!��9�~��_b��̎T�LM����fLo��a7½�%���HC��(зB��Dx��&S���am�,�4B�}�6F���-��.�{_u@~4��J"b� ��]�
x�������ζ���h(�d��t�{�+��UC�r�}��a(��*�b�+��D�y�$��[��{�7��a^rWN�v�"��[B���3����!s�6��Յl�'�kl���7�!�v)Il �a �y�P��O�<�r�u�ґގ�f6o}�%Kh��ZƑɝ�}��OV9;���֍��f�L�(�䝪*�U�-�3�M�d���R�,A�Xv쥷x1P}��͕�Н�Bj�zG�*Y��OY�Z�mk������ ��o�-a��͗%Jm�9�r��2\T�̭�a���S[��e��Ɠu2qa�=<�k:�������é�F��,*}5.�8�7]���.�rr���Kpمѝ��l�ł���W�V�*J��,/�u�xu٣�!V��4�#*�AP6&;�pt�4nU}����e��UJr��L�J0P�Ux1k{�jI��mХ���_>�㤲�*��P3l;��s���fVmonXq��efӗ�o]�H�5���Yϱm����\zD;u��ޭ#�,��s�[)V@r1�)S�pœo����;Dr���㳭S�*�\���\�}�k���H���\�:*a�to1��ɒ���m(n�\BKL� �`Z�fu�9�*b�u�ɢ�E�5�G*�m�׆�����1K;ei�5nռ�����α���o���"p-�+�h��d*�sz��u���z��}O�Ad(7�v*a0y+_N�76��ā
��U� �QWc�ز������t��yܹ�F�+���1u���Wo��2��7���sF����}��KQ#�V�~�ș|����:�Hq>�\o�[*e!h7��x��O�,��;��1[�E/Ņ��`�.�Cc
>�$��h��N,�F����{�f��Z-V����|G�����@�A���*�C�3�g�WtO�[Y�*8�kzA"���}V�5!Q����L������l!"��}��j��H�:F���#O�b'�v�:�����-��m6	�[��f;'��"܉�e�.��]m�ۮ8�ώ4O�b�$�������!�:_�n~��q���MJ6yY^�>�C��#i8M=Ő/	��W՞�a��l�?l/^0��i�X~�߭�����I#��B�Qh�F���gD�?�sS7�2g�js�Mf���q,�[a�oQ���l!��d#��yvYL����O���l��W�[�}�&��E�SR�N>�B"����,�4E��l�gt,#\H�6��l�ψ�Je�<�\�Nt�p��/L4�[&�Ri>a������T)F\��?�s�ײ��$̞
�,C�+�pp��I[9�,!n[��aw��bq=�ea��H���H�;�r����a��
�l~���+u��Ì����j�X�T�%��;m������t�!����i��*�)&{����^VŎ�}"�>RKQ��!V��>1�� ��Ԓr�N�5��Ig:)�@f4X���mޜ|��p"�x�H^�����OtܔM��`�4Cr�*�C���a}q"\S��0���DƄ�lڶ�� E�[�׎��;��.��X��n9g�rl�g�x�t*ލ��r���W�>�oǧ�dC�Y�DUd,���Y���
���T�AP�Hq���[Ζ5�{-8�% ��i��K1���(dq��6x���f�� �M����adT% �"�q����F���1�s���c.E������2jÌ8
�9�d��'l���mv��~��^~P���A�,FZ�4�C-ż���ap�"�H�����<7�V���4����K���c��Q�ҋx���kMf���кp�{Y��cL$�	QbG֚�G�{ �\6"I�4�,!�_�!&u�^��ϹEy[M�"Nx���΄
a��l�"�j1�M�d�]�
��:F��XG���5�Î �qȬa�o�izadu��#�\�����ѝ��&��L�ĵ��Q
Xn��BE��Vp���Du(�Ҷ�il�ɉ!�t�SC]�H<�A��ĩ�d�C�n�#��AET�pD���5H���W�	�l&:��t���_��T�����iUH%	I��)�J��{=�j�9�+tL4+��c�����^����,Q�f�X����ۓmMz��q�m��Ǵn�X�2]Cպ�\�훷96�攇m����k����NW:��#˓�͸<����g�>�XVk�vn�B�َ��n`���p
puc�`�]vg���
skoT�!ӎf3�o��o��C��3���qm[k�m�I�k;��NΎ�Y�����g��n��\����۬g�r��#���
��̧Y���$�H���?��H���1��p�C�4�"Q�q>|a$Q�$�"a���Y~��.��a�l���ZF���$�������E�\7$�ڼE#MǱ�:�ox̑�E�� ��a��޾a��D��d�h�>�7����l�`��o;�d,�����+�	��}��
�}Ap�$�jS�L�����Ylk��$�4F,'j;�rʲ"z�j� �c0j�����J�Rk'J,�/}��Ϣ"w�)�4�ՅEQ�f9�
F!�o};�Ŗ�a[����K0�ݯ1e���#�d�7����g2��u�6����{�@Z2���K�����:D9ĉ~�X��[*	>B8C����Ol1�+���X�H�N*��wU�=��S6~��n���%j�0#��	��<�Hq}ԏ��Օ�}���n�zh�X�v����wVv�F`r DE�|�٨ge�(�e(;EO��l�w�\���<u��;$ơ��#Db/"],#�|�OXG&ڤ�}��[zc��c�]Єsz����#x�QA����{!��{8E�^��t�i�"�"B߫G�\!&ʉ�NCc��^��p��g�`�ŏ=x=p:�?KkD4A�U���3ǹL���Mi�R���J�M���|r�I�L�\�G�uN���U�|yތa�o5���H߼������_i��H��jxyX�U�|t��-	{�u�3A����]���<t��]�'~l�\*2�)�!�LäkZC<#[��;���Z��a��דp=Ue�=c��@����54U����!"�G�����"��J�����h�"6d�8�����^#kh`�pqNLɱ����6�0�x���{:i*�^ma$5��aE�t�����dB*[ז�30���eQE���}>T�Ur_�SE��(R��D�EI��9לn�x�|f6��<��qUC]u����sG��>�{�W]<0����>��pC���g�>�ps��f�Z )��� �r���{U7N�ܡկ��7G�#:����e�;$��1�
@ܒz����F�2$��I��So��3��3Y̟adaB���Մ8�	�TD]�4�B�Y�~��ޑ�
��t�5a���Z
9p�\�H/�Mat�#{���+�\=���Z���O�Ł&�	4�;n�d/խ��kH�����k��Ê�ϾV4է9��ܬ~��܅�w�{��q� �7�sPG�QrM�DVu��^FA��FF��>�`�����||Х6�@'q���^��I/���\$��^��:�X5o��o��շǳw��2��쏆��v���2 ���S��wN��_��aGދ�CNFX�<�M�V^���>���Y�X��M"�BD[�C�x(Q"�Ήi<Q*�N����F�X�;�S8~�=�P�CN�M_d;���l#~B��(q�97I�SO3�ݛ·�/���$�ȟ�߃�SA�)RbGWz��>:��-����cL8l��!�y��!�q?��s�*�f�Ș�I��p�2!c����n�D��\�|D���|��?T�'ka/�m�	�8S��1V���[]'3cH�R&�C���4䖶;=p�YЕsh�?�������XQ�M�a�O'ی��,tW����}�c���A��X�"�H�l$�K�M��EI�h�Dk�B�|��
��\R8sH��6ju!�n�qBJ���o&�CHb8�k;��ӌ.�@��}�B��DY�L;�?2�a����mf�p����,�I�f���ifH�qy�C��Bw��WO;Ib�]�a=���'�9�Y�N8[@��-�O�G�]١����7�Ɏ��7�c��c"TVC���qAD��'$��͚�`���_+���>���ԃz޲3z��]��X�C�!#eru���R�w>2�zyf1RӵaH�`�.����4@�Io�s�ƚ|���l��zcHn�\�/2�ᣓqm�ǜ���2y�7Bg�r�<wVi\�n:��$�5�p \� ��!�!dQ�ڋ�#7��N6}�-�����DPQ¤�G�d��pl����@�����������il����,�s���{3Z�h�[6${��Z��l��9��5��y�2���;8;ﹴ��$�0c��}��h����x�k�g��M�Duc�6cH��8�a���bp�dF��#l�"��<���Ip�_v�� Ξ����[WMC����Ƒ�p������������Q�=��ٳO��2DS�:�i/��k��f|���yV���*�/�v4��q�t�Z���s�r�D.����2�a�nCl�'Wb����0���AQ�ɅO�4�s�v���ܔA�����y�{��c��;
��E+�{�zGH�U�|4ß4�14Q)�Ē:Eda}_�|0�DV�+F��{}ƁG���i��S���oIjk>��yW�͑&�� �ݨz�y!�VVz�BF�!���/ڳ�6�ó�rԆ��%�{'P�-�^����0�ae��w@i�a.�)��a{�[�!��<4���b}�\��֡�>��ӿ9���04>���n�vk�_<Zz|'��WW̩�F��6�Y�a|��=̺B�wv�(��y#\V�Y�Qd�[���B��}ر�݅�(�	�snZ ݷ;���^ʧP���*89��g����N!8�kl�Xye�VN����'��ظ,ݕ����˻hq��v����4m]�)�q����1���1��sp����H��=��ۛ���;Ξ�?���/}�=�8�b��
�F��{Yk�vz�ݚˋq�D*�c9j��d07`��.�qI���2����h���JTڞ�<=x^�����a�c]�\��yg��=��로zsm��1�:�o*�wceG��n�#$M�EBTj8��t�ӄ`߾�ڲ�xa��,�D>�&���2�GO�U.7�,��m<2h����9�+��|n5��4�'������0�L�I&W��zk�Ɛ���k��]�%(�w��h�u����ӧ\I�&��7U�3��@�#X5�z��4�������o+���>�_�	����ACH��!dY=�ݦ�:l�X�9�~8 �8Y�/����!��ī��WA�`951/\U.s�r�jA4l�Ȱ��1���JH�đ^�A��T�o��{v-��s�����C�!��}�j���:���?n^����cA�X�C���m��O>�c�y���1|����E��Ɣ�ACH�,հ�`���؟l5G�1���ڢ"ּ�q}o2r韊8Q��)�s�"ஐ�t�`�:|���}�PXCHg�[�s���az�
(a$��,"��k�#Og�ī�]��m;<�]6q��|���]���q�$$��n.��hٯ���S�/ǜ��P��Y�����ü��%�qB!R'�os��3�#�=7Oү�`��,#�8~�M��ē�G	@�d-Ǽ>=�]0��Α�ϕ�O*��^cV�,̤k��+��ȕ��	�gYWG�
DK��[V�����{[=\�<�)��_eM�x,嗙M��
Rr�߰�l�CO��݊�r�m8C�h� ��2�G���*�I+��&ϭ$.�õ�@�%764T*#$r#�����CV_�]&@`�ñ�FA���z�D-��-�6P!
"��� �������,,ْH��v ��_u,��E�ZW�T��	 �wd0�H�idX�\a��B�4��=a����KAs���%�8����	��c�ybB���'�������S����G�%�����t�8�K���I&x��l�8�"���󡦆ӂFcz����(��!毥4S�MB��|F���@�Uo��<xDs>Yߐ��*�ᆾ�;� �PFQ�M��X�ꋌp�9�lu��˳��FmUK��9���c���q٣�.H#�`���ݞ��F��k����";��<2�L}��f����e�sCg�g��=T>����_Wިp�,_d�Fu�h5-%��2D�-8�G��-�!�P4C/��T0����K�Јtu�E���>�p�\��A���j#bz�E0Æ:�Pb��F�4D.�v�AB�#�C
	D�d�/�$���c��O��zo`(�0W΅��pW��T!댧O<2[y����H��]
j��,?��[W�ɋ���9�3Ix�}eVo#�U���,s�u�V�$�AwU���y/����]:GKJwDǅ?��L*v�a��4"��� �h��bF�r�Om&��'�H�`��C5��΍iq���v�-���� kaDP:E�#
��E��Q��T�;�Y={Q6GN��S����L��$	ؓi!pǈCO����D��p��f�}x�J{�<_Cጰz�a�v=:�m'�jڑ1�<PB�M�0�N�S{����E�����Aډ���ۋA,���-��ݶ��RĜ��۵nD�[PZ��[��N�$��%BC@[a��?|G����y@�����p�l�7���Wнx�M3�l�R��7�bF�h������#���#4ns#L;�<�����C��zSq��q�Q�㡤<VQ�C{9_��A� �)am��]�tr�C�k��:x�3?~�CP\D=9�H9�p���5[1	e�B�-����"N���{䑑���&�I&WM���XoZ��)�+����=�2���cđ*�^�ļj� U�0���\���\ln��[�9��#�N鿗1&5�$�bH܈&�
��a��d^�s7�o3g,dJ��qE���(���*�!X޴���ިh&z{"d�dæ8��˝��̆s����ԂGn��}�Z�l4SW��\��gL\F�׋�@�_gusk+n�_n�x�wѩ)��b	��7�j�{�|�~��:GH�H���3~���p��H��a�E����CvZN�j.i�������TQF�Z��C��%���2�c)������U��L�k�۪,��.�g��UQ���[z�+�n�Ѫ���\k�D8�u����2u%�m]��*E�����-�]������39� OOtM���n���0C��V'�4�]��m����ƭ�2�Qy~D���$/߶�]#��ZC�����~l�Bh�Ā�X�C��)0�x`g�,0�L0�X3�l�c�`�g[/j����RPZmՆ>,.��လ�}���H􇁄��sݻ��׉ņ�|��%#�Cb8�xd(��g�c��9�Y˖�a���1���C�ϭ؁�]2�5��B�o�դ=�@�[�t��4�1�����6���!:��������EQ:�%�H��p���t)�� �pX�#���W�
(�;����]^{ܱ�u/�-��!�I�,����Ge�Af�����{�s���#�t�!���F��N6���
2G� �C�"���{�ݒp睤�1x�Q�e������&���U_��Ʊ��g�W]!��C�A�R��% p��ڥB^���W�]�u���E�{]����~�,��I�l�}�2Z�3��Yo����9�H�E�e,��.90_ʗ̆��C�kQ��(��Xo:�u�b�2�]`�S#GBwf�)�y�&��J���Flk5�[�<��vr��.�ʼ�t��\�����Whll�WQ2��9g�6��6�6��ΐ��sB֤^��W@KA뿶��yNv��!��86�L��H��7����T����&K&�8��p��z���7qo֛a�]\��9x+����;[�*
^.'W>wyN�;�������R�n
�Ňb�/��j�7�yx6�TAs��Dp��5OkuT�����!�����}��x�Q�OZ.t�㇚������nƺ��կO�h�E���K�d��i�yb��uڮVe�mK��3	�����V*�:�Y��>LVMZ�s���|TE&����e_��8 ��J�4���T�Sg����X�e
{�B���s7��1�b��k:`�z��x�f섭�ե�ٹ�^51ug���[ 7>V�]N�V2�x��4��h Ѥ]���Ե��H\��9�S�ӫ�3MK6�C_X�%�7�s��vMA*�&�7�+f[�áSշ#8Dd3��_r蝷�r��՘��ޙJ,/�[��v��e��oe�.F��\mN���L
b����m
޶Cx̛���p
�M4��}��Q�y��S�Z���J���	�8�j�3`AnʷI�[��n1$n`c���ڶ�7.*85�܆�7D�q���O����)��eуnwl��l�RJjn��u����{q<^�>��(9����qۥw<x�Sg��m�J^�ۣ����
�,�Q��s�gFI�n�CK��q�۩dۭ��_+;Ѱ����'S�>�>���;I��Lpkge�W�:�3��)��>�����6��xz-�Ӈ�&u��7��^��E�n*p�m��u�viWv�.Ws�.�΂P�x6�t��c=t�+�c�[�sO�g�GKB�p�k�vv7i�zzy�&0��t�FM�R��Ι��Z8#�7b�1�u淌pdx�e����%^q���Xi��͟=�V����e���c�'ѓu�'-/n������c]˲a��t�� �3��݂����|���g� x�`�7pf���Z�[��������v�
F# \<�۞���kd���p�gZ�s��c��7mm���<���Ѱ���{�q�5�$�wnŻJ���a��d�x=�P���ӎ�8��$��4tuɸ��� �]X5C�bx��4�xc�Au�[.'�Ԟ;v�.@ݣ;-��yEW;:��g8jx��!�qJ��rv��p�b��Wn�s]n�"<��q���ݟ(�&� )����sغ㴎����>YN1kv��6ʉ��ݲn�l���j�g��x�[�W^�{��q��ų��==�v�<�m1�)������V4qs���y��a��#�=��nw&x�.���4�Hn�ܒ��ͼv1����	[ZEԯHN�	�=rOW��l�`�m��v�]�)����m���1��Z�v!�`�T�d7\p�\=^�2m�ջM�����ם �Vݎ9�ϓc���S�x����]u�=���;{�t;��{V�7\�ە�}��Ӎܣ���umw����D�;*�4/C���	9`��p;�㮮m��\��ے�V7;����ׁ�S�c�S 9�p�b׉��Z������1c\np�C&���+��Z���|�ݏ'=�V���+Ƌ=��эU�������{6=��w�~�k�dy�p�z:�x��7\�j�8�:���d�<<P��c��d�2�u	���u��\.�2�m���e���E�6s׶d:���bk��v��8\�lxޝ���<vn���;�q���v�uO>�c�7-����ݳ�ܵ�Z���k�u��Ng������������c��w.�yK����'M�j�n����u��v�#M�@�fR�O�����8ɲO�C�`1O�+n��ӆQ��y��y�>#�!�|P�g��q�$B����ܤ=�<[h=����ҏ;�	'�AK�������X2@�PH�N+E��8�hQb훝mBN�-���t�>d-��1Cr�dn7��d1��"/�j$+l�c?6:!T1�*W�*��`����<x-<C��Q�đ$@��		"����+?y�b�_�o/�>�O(Y���p��z���*�L
,[�q�\�5�9dY�� ������f[�JqW�!�
s�E~�!q��%�a%�!�9�'P�Ǆqc�ѣB����"겫"���`5�"�\Y�� S�s!��p��?dC߆^*�w!�� �3���$sH���JX|~�~<D��>��.�I�A2܇k���oe6d�.ܺ,!d�2B���̖!��?����oVW+�I�%5�0� o�~՘puU�Cw�=3�0��,S{0�4}w��D�M��,�ZA"�m �p��QG"L\�77���8�nz�u"Rg�\��ע�2u{8��m"�,8���q���(��^�^6`D"�8���WT�娒���"�8�7�~XCㆆH��G����h��i#H�H�>]��� ���'\��ȇ�(�,N����Bq�pf�.7+�����d��p�ЙF�]���L](�uk|��,r���zGZ+��/�F��WϦu���CƁة��n7�F�nh�-�/�#_r�8X�c|��'�<�@�v"������PF�D�p�j�}���������r@�lHPaG���~W<�&Ȭ��񿻖��2�P�����`T5U��<�>�@8��e��G�l{g�P��B�#H_R����j֚O��u�p��y�~%�!iH�m�Ԓn��g#߽܉i<>�h�2���QC[&Y�pW�{vÉ:׾>#K~��t'/��7PY+���vΓ=��߸�������/+�CL��H�rIa�]C�KH�x�6D����c�ƃ%����K	\l�}���
[�^�F����5�	��ҁ!Z�/��W���bC�����j3�=pgmeD�pH�0ҍ�5lEs��N<�m��ݻv��ݎ�c�;O1F��H��a�}da�~⯢6Y^�}��$(���@���ƆY�Č���Q0�ur���zS<���|�$*�zA�o��DiZ��b�C�Y�(�Tp$d����(���/�����v�*�2$<	��<Ge�L���t+�_Y�.i�>�;5P�1H�YHL`��ֺ�
6B�݌x�	���;R�X'+�#��M)A$�>㐅GH���}:,ib��(�A�JW���ڰI�`��X��<!�])�.q�ȡ�""a%�lD�k�wպС9ڔ
�u:�7B���u�dB���]H3Jvs�s�na����B,�ý��|8c�*�D2A�ˮ�g�zx#��]�_�8"�F����r:E�Xl�X\�6ld?��L���'u��Df�I�Թ:md�Qc��6qC�ƌx;�n�${L3a�_�R���c>cMi�>8>}Ud("NE!��h��� "�h�E
�����37�
v�Uo��!����3Q;���Ug@��q��߆��V5 x�-B8��j������U���A�@�g��F.�r���n|���X�v+/��Yإ���}���Ϳ�L�#M6���<�m����aqa���D�x��e�`�Zx�rGZ�y����-�i^[i)��Ê-���r��%�NК��B�t`����j�Fe)$�x�c'�{͎ɯ\��s�W����:q5�.���q�<��Sn��e����+��G��ǨF�˖-���'H��=�U8B\�f�0s���`�%�����$)�	�Ax	� 9&�2C��[H���0E� Qa�"�f������6���<d��0����;CQ*���_���7��A�W �XB���o@W㐈�,�[��$[^/���|�x'���(����
����8����cdz�T�F��^�5��B ��e_�E��u�\d�~��xԜ�?)�	��9B������_ꈑ;��_e�<�W�:wMdTf%�h:�D�;�)V��֝&��;���u�_�M�gz���-y��8��MD	nB"C���V�=�m����`�±?��=+���l���^���W�U �2D�`3�.T�!�Q�F��u뭊����4��ч��s��3vV�Pɣm\��EFS!��$[�n�~`�<~6MW�9�x�D)mW����D���}�Ko+>�������M���lz�-����PE$rP�v�#�c1g�L+�ig�>��yJ�e(A�2r�U��:�>�� \�
[:�0`x���>��P`�=�J�ap�"3�<I��M|0z���ENZ�Џ�t���fm|X���y�!:ai��d�*�K}�������䄒���
��%}��}���~ѱF1�L��?L�E��� 1
"O���߽��b1��F{k�,|r]�K�M�}�ϓ�%�`�(�m�#�m֓��0
=^�B
n�k��U;g��{�*=�Y\��^(�RѡZ~@�W�,�^�{`�8����T���^kV�K�o�Mt�.�C�+���6
�ho�fS>�	5�{Zl5ڕd*v�կ��8vЮ̮��5vSĤ��M��	DR%6�bm�*r��	ۃ���y��[�ƚ�n�1{�(l�rF��N;��!�
�u�6�3��(\��ShM�: 2
�Ǘk�g�{g�{��\\�m֤�s���C�����v�c�b��;�%�Q�k�[Y8���=bˎ�V���hw=v�k�h6|j���}����v��<��h5Ԝ3���'[�@,�%�6��l�t�f��:c=6T��5�Z�I��H��7�䄮Kr�s��]sq����[X��WHMU�ϗ���B/��{�:܏�����VY�j�'P��k��Ϗ�Z��>~��ͽ��'��/e��,�caHP���>���5�V�z���Z�R1%c�e�Y
hu-����u��u��w��~Od�_˻�e^����9�-Ln����p���z�����C��B�l�Q�y�<��{�b���s+v����}�_V����gy���
p!n�]�nz	�u0�����}�G�c����W��;����q��3��z��T��Y/��3!z��/O��1���n�06܅c��޾���dUY�z��kd,ŝ#Df��b�H��c�r����@Kmc��2���������G�6�N`�~(B`fF�͛�{6���k�;[�6�1�.�f���um1����H��$M#�kn�#N^�x��Bz챋6���"�]�o������joؓf!��5��/=�	�!�'��[uÞ����6ŀ�Nx}[Ύ0����6�&n�q�`����=k�"�'����63�1��<����%���ǆ�V����l�m�l�^����}G*��<߶��v1�*�t�`�S�Piȁ�
�jn�g�&��QFЈϔ�2|2m�Zm#�-[�*{�fɺ4-��v0��dsf7&�mA���CH��׎�*�߭A�[	�`��(�1��I�7�������SP�����;>ۄUuy�~��mN�����T�r�7�w�9<�R{�w���k��Z�Ј�,�[��d=3��GMa��{iL �DC��dF�I�p15���u�U��Ǘ�6Q
{ִO���\x�v�byp�ڠ{�뇚cx�vL.���g,�&��r
UT�5�h�p��Cu�j���Wzl��j���c_!1�_!����}�C������}ƅ;���8`�B�� ��$/�*bHYh9"�.0��]Jz�� �Ry�#��+�,Z�ֲ�s�9�S����2���%����1���c�+�����߅�&.���H㱗d�.���Q�g���es̮�ۗ��O��3��t#�H{�!��Ž�ۋ&9��������-�����d��,��h�A=�
�:��`]39ܷ9���yli:7uU��ǵBoޕB�G����*ډ,3������j���_Vv����f��@�ѱ�"��ܸέt��s�����:-���e��@���;�`Q��;<���$�P�#��W���^k�:�M�6/�7+ޘi�C�]�*���L9oW��~�/���%�[��������r��g=:�� �q�s�v���<]���{)�W狏Cm����!:�R臈��
�%[�my�����!�n��5���5fHU���;k�d0��|�h�2�HU�~�AQ�$�2ŵ{����|���ڰ~�+��T���~	OOI���u�x�6���c��t� ڙ��x$��(�	�r�ɨ\��:禲a��_���;��z9�&��X�'+���E�;Y���;��
��2�(D���e0�9Y2Ux��6~�@��og�&�K�C�˃ivm�t������tjnT��y)g��+^�[٤r-��G���s	�2��,ޥ�L/����L�_hw��&^�������ͳ�A��@2�ם�ݶ�a�[���t��I8E�r-����r���A߭�Rp�FNL�.=����As���F嚻�)
�)�ޖ��X�ꂇ���o���yǟ>ߍ�.�؇�C9�nͶ��W3�e�g����C=T�w,�����nݹ���}v)���xVᯫVD^���~w�#����2 ����p��M�cE���n�p��^�8�ҫ#
_�W��aN��4ԋu�h��>|7��z@��"�35đ�+c$�R��AX���ۢ*]ڼ��N��'���?i,ax����2�(1��V��e���x��M9/��m����>�|(Ӣ�`ժ������W�;7��?F+��E�r8�DB�L����Ȣ�^���Z^�q�p;5�A�֯�U*�m?�d~k��7wz�D"���;ؒ���!|=��KPm)�F��tX����~`�ύ���G�� ���/�u�9Xc�4�}~�ln[P���jׁG�T����sT	L��"i;;x,���)��&�\��Yu7X��w�	�n�FTmn�NZ��ve��vQGk���`ee#G"^i:����ڇX&��M�"b4�04�a@����/�u�V�]:ì�^�G��qx�F�M�7[b��m����v3s�ݩ�\h؎M�xy��g���L����cp�lltT��u�r!j�N�ҳ�z�c��=�+���p��n8��O;m[�n�[�/�A�6�%���w;�89���a��;�vۉ��q\'���q�A��r�%I�\j�랎�h��}����fq��!v#�����pq��h��ntm
$=]����rg���s�Mn*�ݚ��o��������p%ǙD�2�� 0��`v�J���{��籠�{e�V!SA�q����>�b��&�8d!��dDď<7>�lv{7Z:a��S8�]�R�f�jqe
][tP�f���;l��"�
b�X�L���'i#���Ch!�{�EdU�����fٺ�B5\�A������q��k�s&`c�̪=ҝ-%o�g�zr����4	��:�F�m�ɂG#�xY$TR��wi�Q�֪?����^G���Y+H/��_`�4iH�Z�,~������J�W�,qF�(��f'$U�63G�>%���Q`j�I�cMk�ə��JaxBpɵl$)��ѱ�#(��&��(a_z^����q��M�_O&M����ܪU��v�{ggnq1==���
�e��.�t�!N��b����_L�2!7|wo0��w��Xac��:co�_�g,�"��n�=�OvN(aƵ^�j	����/pcd��![�}O|=���]���C�Q�`I3+2E�,[]3FԌ�����e6;+ /�>0r��X�b
ѻ�"u�]J���
}�h7Xe)Y�O�Ҧ&X}�1Ӷ�ӭe�ȳ�����S��Y�z�k�zY|Gw���|dlϡ��Tr7���*A�-��huYz=�~κ�Rzk������DnW�T7ɺ;�Ҿ�8+U��K����"�*D�M���E`iͦ��Xsr �nodj�z�^�*Z��<�/L�9.�G�6�Y�+)�6a	�V�,1�k�DOf�}Py�����X�||:Z)���#&̙�������ޙج�8�D�����ZUZ]��Wa�w�*��,o�.�k�/�����>8������C�h��ȏ&yWm �A��9K�QvR�ۚ����MV�I���Jm��(���sH�q�d�CHB�Ցm \y:>��" #r�Zo>��:E>b�%�T;<j<��m��ڶ���z|1�4�~@U��lFӀ�����Yv��eqZ_{Ի�"�JA� Xr�.�KS�^@#��qm���d�y����SL��"�
׮{�Qʶ�&ǭ�@�S�[-8�L�+S?]�咶�ֶ�������
#J�}o=[����^��2�N��ZH�JKʓ��~7H�e{΍'�c�^{&�ٖ;�;W[�G�7E�V7��vm�^�A|�wl�8���U�ZCwz6�U����8�n�ʱ����
F
�t\�WBN����9�;�ɡg!�W��k���w�m���T��[G�����%����ml�b��Oi�7�4#��D:�K#(<}�s�aO0����n���U���olҨ�wT�a}+�5���˕���XWH�����Q�K����V�5S�㛻��κ0�j��t휃�9�Y0w��o�U��Qb��m�o"��,�^��;\B�tZ�G%6���ө�쏺O�;f>yf�4H�8X�V�8�jf��xwhvdz��wq��]:�u>
�tHJ�oPa/��2��\,�}�*̢�ʙ�F$�W),η����R�FqծS�+2V5%&8@4_r
�+:��~Y��6!v�S�Ӹɢ���]�-ᨛ���}{�eJ�iݔx롕j��̫���r�L�~�K��yb��L�����Yr�J���\�2��ۥ4w89����Ê;�7��>�,p2�_rU���A3Ga�A�)[\GZ�KS.�ֻ�qV�Y��4M�5�y.���uÒ����k5���Y@k]e�7re[�/O�W���w(Р��>�JNc��v��if�:�̬�I�s]Q6�p��5z�d�9l�U+Tf뙅��*n��61ړ�G����j-�/��n�/.�/�^)��c��UFPˤ.]�F�����f5�~-�o������n�]78�k������$19f̑�qҳ^�����K!x^��z��(P�z-gٖ�㳑��M��X#����njy�)�8UxgI�cvƟE�s��+�Ш#.�!I&>�|�����#b�Z���V�E	�Ǧ�W���?�W��L,�2/�����! M���!tk�U�w]�d7�V�HB�I��@ȷ��Y���-�Q �kb�˙��˱���X.2b���2D���	W�X«��b��Hq�o���]�1ؓ��G�,o��1��iZDV��(8ͦ��V�{%��gg�Y(R�q:�!���-)rW��ʠn�}潸�<��η���g��r���ߕJ��M�{�p�`�+.���*8��W���%�_���׻<���M�
Ee�1#���y.�T�9]<El1�=�~V �4�c�޿�UyÛ�E��!r���_*�������Q1��͘���U���d���=.�}����@U�c����j�3Hׅ��C��9.үe�\|���;�F�ibC��%m��g��]V�nA�ze���>1���v_�6v.˽�.��輅H�$[�9�:�b���Դ5�vǦ]\��-!�Hx!��24l�RH�+
j.E��ѻ�� 0ϔ���m�큚*�Ӧ��N4���1T�/H�i��i?��N��ߟ���@���,����B�	�1�f
pB�!�mt�v<�nnۨ�3<	=SN�0Q�f��{���zkj�,47��|���p�*�y�XMq,��?e�(�޳�7~�D{�m���R���'���"�"I����c�Xu͕���ym��`���0�K|�͆4릏�o��f_���L,*M xz��V��G��'��������rS���I/�Zh�H�7^T_ʊ�M{�WE	T�|'1�u$�`-�P���!�����x�o ��59����t��(�rD�C��|�8E�� �:�c�����w`o�r��`�g�s4��ȴ҄�=kv�,�8���4�&��\�$
6�p��+O,�lk�`����s݂�$P���Wճ����}}����=u@J����d�2!�v=�Y�d��в����zj�_{Fq�
eC�E')�Ӷ�H�`��y����z����eл��ǈ�������L�%ՙ+�
��ݔ[N���gW������:m���&�4�]wb{���ʥq�W��E�cm<nP:��n��s�G$\ii�n��5qq�YM��s� ��\vݥ2�c�0�kך+�ݭ��=��3��X��uՓA�7g�ꗠ}ؕz�����x���yٽ��S�0)�vs!�ַZ.��h��t;��v�������펹��c@;����v�����Le.�k�׳ƹ��\���&g���pf�F���� ��y��;n���,8����Ε��},i��cq�`�vyء���m�=�xt��x"�͊"�V�Dq߹-J�:����T�/	�F"n	$9Zx��"=$?��U�S[q���cH�2�d0��Q]N�L�*�����m:�"08��;��i���	8���kK��`�ƣ,����ݪ�v��>��p�f����D8������lK'��rg��#�B[�5�?Y�����{�� ����&}�	ܩQӒ �iż�x���۹5w�߳3ՄP�*�k�0���KͿ�C��waUc��V@�C�nv*g�\a���#j�ɥsՇ8��G�@k�@t@�cQ��p��N)aH�/ˮ�cY*��휨�>�kV�8݈*'Ʊ��^�Z����F=���M}����xe�>Zr���6D�<!y^�u8+���Ͼ��q��y˼�/�ܖ9�"�nn���e7nzpGi�|<�P��]�W�[��������_�[��j��]�f����Y�:i�3��R�j�9�o�r��@w
 -�@e�b������C���p�
,9#RAc�J\~/
���k��T���v�?yǣ}�WB�s*l����"�/j<�sEηYY��%Tއ��bW�au��u�6&
��5mSv�c-��C��w���_v@�ƪ�~ٚx��p���tQ~��(�o��<V�&<�T
�<65��$P\�%X�
���K�~�u�Ű	�I�x����6�}�@�	�����[� ��Hp�V���qr� !.�߇�JĐDq��LH��?f](>�da�nUD���Ê!<<�bؐ��O��NG��z�a�k��G0�m-�Q��{��Fŋ_i|P��=IB�I-��ԇ �^ю��F&���.������0ø�1PI�G�5 +���U6i��d+�W��3���mZX
�����zx������ʍf%%�{\iݺ{�6�8^̀���v�ci��m�'���b�����#���H�c^��~s5|�NW^�����T����c:���0��AWXT�%{��p�����Z놹��)q�02���+N�#@����{�c��Y��5#�
o
4D }[3p��yr���Hqs������_H�"��[��v���#�0�`f�$��\��$i2�R8�F��@Y����f�o6�u*(}p��,"J��!b�vSca��7�����DK.�M�|���fP���N�HȷAg,�/��]�ʻ0ouo^�icb�^��_	u��'���Y�?x��U�V�T�ix�y�U�:ź�XjzP9��M�D�j䓀s�a��\����X��r�<�k��U���7K��� �˕f-�T=��3w��sᮈ*�]yG��Y;���&mWv��C��f�«9��m����Sr9��Vƺa
�����Aa2#��b��չȌPv|&�ֺ�یT��d��}~�0�x���0����Z�z�c�K�7Uy˰�J!��� ���޶���q�ݳ�qcl�sźk�eg�uv��/lkA��5m��k�Hx4��]`,�i���>W�j����������5'H�Z��9�w�o�'��l
���g�����IT-ֺ�J��Ӟ�	��mȡ-5,P|��,��~���6^�Ͳ$�>�y<�]u�Hc����Yu�p���:E*���F�-T��]���a���w��ƒ+|����qң�{��H�*P5 �����^,Ey�V���M]4�4�@H{��,f���ܽŦ��6 ;��T|��b�
� ����%�f{]�(CXƐ�xX�Ğ#�3"a1��e:�`��ki#,��b�4�}�Af��
��˞w�]l��N�5���Wae
>K
W>���MU���qLɋ-i �d��][h��Ǖ)q	�m��뺜|�&�i����{.�&�t%�Y��K���(f�y�r������j���bxU����(D�&"i���\�E�\!�5e
�>�b���5!�KH���h�wŏ�,
����J��>\�c(aQ�4�mH�z����j��04���۽e�M#b�!���37Cp�g���WE�=��� �;�xƒ�!,.�2b&F��#*��=�<x��`*� ,{��+y\t,���:{�$��4�50<��ꪭd36�����y�8B�G�)����᠄\!�l�;є�����m��`G��08��Ļ�*xz+�	 ?��{�s��*�X�`��M&8�_��j��.���A@6@�{4N &ϋ���fX�Gp
^�{H���Y���NDPaI���Tt5�#���`��j���Wr���5Hyb����� J���Ƕ؄�ڇ�V5�y�t2��H�H44��,4��^��M*��C
�,%��a�(��.��]��;w=�5!$�A9��h�����)h�݀I�U�]�G/����tt��{�xn�H�\#�4.�$�E���KF�J�hY$l�Xh*'��<A!�1�"�ܥq�@Y�TF���K�9�T��B� j:��,������]}_b���Yd����8!� "ŚZiI�^��+�M@�T6!����=���
���K/��bDզ���&L8K 6��/���(������1.���7�qXT�8�SnYh�^��q.*���$���v�q�F��RQ��<#`�gf^C�^;�Ύ``�̜�M�8��k �ۍ`:��3n^{\n�3��hˋ���v�E��t�t��⃍0��W�bmƼ�9jKb�vز^{pk�WnM�I���Wgc��Wl[ͶY�Uo	]�4u�������6�>�d�@;��fqّwg���wj'O>���vҬ�����Rʴ&a����]�ìf����۫�����l�V��וu�%�]�k�uǒ����qi�p�Ҙ���߮��G8�۬#� �+�cL�Y�7�PN�A�n�X�("@Y�����#"�T�+S,�K���g�pi�(0���5����,.RH3n�H r���tyl#��a3RG#�4��!4�@ ���c���Ú�0mU!�#ӓ��=4��0В�CH�	=~�cyH��� i� .�7��Eitv�)*�|�s+Ő0��7z�'jS*\8��WMpf��u\T0�U.�{���ҍ;5W͸Mp���R&��se��Ȗ��Wu��	~��V����������
�k���hw����*U�) �F� U���န�h0�rE`i�(l��N`D5��T"��}�t4����xjQ#�ẫ�h�!�����@� ����S)5V�4V�='��L�v]����j��7WTz@B��t���Lk�7���!GB(#rL���ToX�Uf��K��u�r�V�A�M3Cy�������zl
�t,���� �:@���嫠��U�V� j���Y�����A5+C�~`#�7/)>�˯V{�؎���TW_�6^��*���Y���Xy@�d�n2۪7l��3l��ivV��Ρ� �����W��nq�P$��C�.�CH��h�p�X:j���� L�6Cݫ��f�+��r��p1\"�Uq����=.��CƐ���+l *'�V֢!Pʌd0�p48(�!��h�h&k�N{�������,[�RF��O`�6.����mkn����TT�U
�rXÛ���j��\S��s���f�1꺣,���e�ʭW���4D�הizȫ��
@�9{��`����H" �H{Ϙn� �-"� �Ҩb��9�V8(֚�E���0��h"�4H��W<�	��*1
Et8F��Mm�LQ�_9�t4��*� RGUU��W�����U��y"N)�4'.���Ӻn��,j�P�P@��UK���b4.��R�$Zj��B$�������d�F	 �Y�KV{r�Ň�Up�-R�8�"Qhb��� �W��(����D4-�T!4��آ0��(֖'��p��3
��u��8h�:�tI�5H.��3#���,�#� XY8^�+
�G|/xl
���T/�A�;c��u�;*���3�Cf�PB�EuJ���E��D��C�hM44�*��r�X�f1]aj���D*�UФ�-��0������J]y�,�b턮�m�{bv�n6b�ʆ�^C�.�Sҝ�sc��9)B(�]�� ٠:ª�J��^g�s	�]��* 0��D��祀2�
@f�"�՗�!Yמ��`+��*�Y��E�j�^��t�vi��B t����Ht4�C���j8��G*@�-3$wCH�@�T9��0��4}~�`V�>q�m#���ݪ��@<4K���=��6 �lP�!��@� ��<��� ��VC ��T������pj�i M�u�s��<&���y\@p�a���+}��6�rK�� �Y�5�@�W�@0Iמ�+Mte*�Ah��j��A
��s��<�UY���n���~rf��2�%�=g
�l�ձM�c7���صSh�4��$���Ǐ�+(cE <��ؗh�z��ge*{f�|8��d��ܝwLQ����ƻ)�)�����M �
94E"( H�ix)�a'jEuCM(����;�$�T��ۉ>O���y�@48� a�d��U�� F{�����*� i<���Q�"��C�i��'��VsۺBM�\{{.�+` :���5C��$E[��y3��$P�Ĝ�8E_ Y lP�4���t�%�!�i��$y���YE�(���U烵e�<,�P� �M�a ;�LV+��3	�@p���F�D��yX�"�hV0��S�U�P<<F�������Nu�l���!R�K:Ѻ8"|����ޛ�j�CnO;���dڍ7C��i��{�{ݲ:$օ�׈��U�_.X���Xj���a��4��%���pV@�[ �MW@	�Y��N?mr���R�U�,Q\"��D P�󸮔HCM�QZh:#�WS�La�^<��n"�)8,���B�P�1�@a4	�,������57�����lzEi�H� �L ���`4Mi��4��U�UG���udW�,��@�MW 9��K��P�@��/@�:h:<j�����\`��Dۆ9V����Uf����@5H�}k4]
�/���)�R��}�L�| ��j���)[9�+��cS���,B0�������40���r�] 8@�c�4�MT4�W��JKD��E�S�, i��,�V��Y/w�4w��h��+�8k	UB*���ȠȪ�{<�U`#H��B��i�\��EWu���E�Uf�b��5c��gr���{9����a�\�^�f]bg�ʱC=ԭs�S�'f+f�Ml� ����Dl*m��.Bl�V��Y��[�J��� v��E׏H��ؠ8E�)���@c�[�|`����1���P h
��a!���E�WH�� �T�i�7��t�^�u]����+�
h�sqX�T4��U��d�oЄ 4�Vx���C���w���n:E����D\V8�-˜�f��hH��nJ��TeчnͰ�n6��(^n1�s���{�ߍ�V@��5UdP��y�t+H5B�^� "�H3�xn�t��T CC� 
�*w��uC���;c��a��r�"��5B�4�C����5@CU\4 C@W��?$p�%6�qX� PdP��P����>縬P�B�sۘ356�b���D��C�
�wO��P�*��U�(T"��g�, ��Uf�"�pС��*��f;�"�@WO�9�uWsy�PDP U�@a� :��A�@�H).U��Q�P�C�UBȪ�@N���8E
�UU�B�5X����,PH��Rǲ�j<0ܪ�E 4�j��y�+ �P��qP�R��K\���c��p��-0�n5U^��a	6�J"8r+���S"��3P�`�	��;�)�C���b��h
���B�
� Q5Cs��`5U��f��UU�Z@ {�[�`P�*� I�G�ۣ)n�æ#�	�\]Pj�wXh ~��0Q0�$�#��WUj�s��5@oy�+�T4<@� �y�;��1��_:��u	;aX�ZŻ�}r�A�3�
��%@�P9	P1�l%@��|�P8�%@��P?��T�*`�*���J��J���t�P6�P8	P4�����)��z�)���8(���1�|n�2m�Zh�ZS*�dRkT�F��%3-[[X�����5�fRV��v;2�E�Fؖ�+QAIm��fͦ���٬��   �  P                          @   $   (    ���V���^M_>go��m�_-��fL��6��=ݧ���z�v��������v�� =�q�>���g��׺�9��������Ͻ���|c���m����}�� ;{|-�٢�o'�n���;�7���s8���UUC� �|@    }��x�      ��� |�  �����V�ww���e������t/�w���+�7��|�}M�}���_ �/�b��j�����罵�{k�o�z�]����������i��g˒v��f<}�^�ȡ|         }_:�-��M��3�}�������ͷ�7{�u�.������k�u���{7m�� {�o��վm콯��_(�{|����Ϸ����|���sב�{� {�k�K����s�E��w<�0p�TMI�}�V�Q6���'�n���| �z>S-�ϼ��.ܦ�;�o]Y�v��|o_{�]-}�|y�K�ֳ�}�}������s�5{;ϻ��}'cϷԯ��6����7��w	UI�)  @     �aݺ�zw�V�v���	n��=���&�����S��� \����7��m5�7o=ݶ�s���ݕzw�R�S� ;�_pk]��m����9�R&�Z2%��w�=�i��۞�}���ܷ;�} :�_S��}W5��}�mc)n;](���={kl�� Jz����kݝ<myc�h���vw����^��B��
�       �=R�k�^�]�yu�o]J�z�/'Z�ݝx ����^{�{��������j���kLe����U��� �_m�c��n��o���������#{iyk�,�g�;�z����=���;��jV��+�8���՛]�U���@ ��ڴ�y��	J^��B\��-׍����[k3UA*�     �  ��G֕�3�w]u���E����q�z}��;��P�}�� _+֊(�c�0:(�ƽj{�}�������G��� �>� i������z(o�P>��>ڵ��
/��:*��<��{7w'� ��|�8��X }��:|��מ�Z4O���L�hx�
\ѡ��¼G�(x�B�&�8�������|��U/�P�T�@%*P)�IJ�� �5=1*Q�   ��U*R�  T� ��E ���A5%T���~g��?O�~qW�����Y�	an���� 8}�3�Q�E��Z>#Mj�ZQ����X�34��!�x�Ib���bI,�Y���I,Y���$�,���X�Kfa��K3f..�����'�OJ��k��M�Ni�����)��]��{��b/SE��v�[k6;�E����w{[��։w��v��kc+-�O^�Hn�.AI-.n���(���]IW�M��np}DQ��"�s����t����8�e����O�K���ū���p�n�ͭY|��R�瘱�1m$M� ��mH�<0Js�<�K3]�N����e��Y����p��V�%�gY��ª��1�"�ru�41Ҧx��p��fbڔ���4e5�#�*�ۻn2�F�u���y<��l>��+_��=�.�k��1��h��dvb��v�=����J��3���f�nrS�򷽝���q���C3�C�"���:�` �[{h>cF:����S��P�q͐��2��ְ��S���U5�U�bŉۘr�"��WQvm�Z܉��*7F-�-$�7l��D�,+�u�����#mG0���O@ʩ&\[����l�-d�6���+A��D��	֠U*^Y�G>РI� �sCL(���T�NDF�dI��Q^�%��p�.����y	z�p8�D�B2����v*^/r�Y��6��Џ0�sa�1���;��̥a�Yj��v����	t�f�ݻ�i]�p�.a�O<�f�$���n֝<{݊��CO[�u"�P�ҁ��-o^��^l��WN�G�HA����tO^��b����N[>��LCF��
lңZf�yJ���C B˘��4́K̺�nֵQR��!���un���W�qB�� �1�Dc���ꘂ
��dSr�׀*��@��@�e�AYJ�2�lJն8a��v���hK+����*��-�ec�>��7nK7�D���O�ur�!�*�ccء�=�j��}}Qa��)3�U
��7�+2@04�#���,�vmm�7�cX,$�me"�$�ҋ9b�"`6&m��k(��b��/�;�H�N�ۙ�鳎�/3�-���Tz#�2�*Hr�� $,N�4\E���&J�y��̆^�B�P��I�=1Ec�[�2�7iam,Jg�S���Nb6؅�X+ᮺ�f�!T���s[���u�`�=��3�-�j ��*�h���4��Z&G����B�K.G.`��Wy�ջ�TEI�U��wa�H�j�(��2��;�쩎�ݞG�l;1��)���/��ǆ-#��KZ9`�xtܳ����u q��E#�rSxz*ǹ���);�ī�-�v��$0��ۤ\��7�gKI���h��o�^�f=v���d,l�8㧔eӔ��R�˫)�6ܦi�X�J�ݗ�(t��!��Ո�h�p0�c��"e��`5���s��8�ڒnJ� �.+F2se��\�X@���
X�E=6	S0�H#����wV��"?��hMB�#ݨc�q��,1E�-Ҽ�*ڬ�K͂�J7�R�5*�����:)Lۓ7n孓\��H;W�Rgw�oU�nFF�X�[�A3\�,�GF�&���ҭ�4<yYWKpʌ�*�&|J+v/nzn˩l�vf�[1�A��"�m
{x�Ʊ��rdbi	�ekM�ȰcX�&圧�������sn�Y����Z�eYT-Ib��:t�S�q��ear����=5�r��ZU+�ޟX�`5{`�j�TV���D"��7Y!�{-��q����ਸ਼j6�Ëב���~�qҥJl��tn�I���iC*�&;�X���l7`���deVe��5߮)�ˁ�7�a-9�@Џf��ۗ�hG�A�Iә�͕`�H;mⳌ� 6N���`�7:��y�فJ\65b�jI����Iz�����wF�Z��7ʱ(�j���t�����w�i��"���Jƍ�Z����ڲ֛��-���b\`eA`f�,�i�t^'�m�2��%%��V�|���)w\V>��lnr��J�#�C��2#x�2lN�x=�pҴ%S�P^�_10��h�&�F	2S[��5}��Ӂ�!Ѯ��JE���V�b=�5���f2r�^�a�3.���0;0֪$���5�M�yc��I�mk�f��:+��QQa������U��@�Ȧ�ŜW#U�c!�Ƕv�1b��[Y0SZ[��4��MU��D��T%��Sf�r�;��&1��de�� x��ԨԦ�wv��l���͚���!1\T	���z�x��[/H�jLtt˱C`��qV�tBq�{��t����&��	�¦Ӱ�*��*�IBM�b���F쌖2���b*Δ�^ۍ��n��2���b��咐~�����������ȂfY+�4�w!<HUƭ`j�:/�a�^h�M�t���ԕ"2�-n�Xs!H�m�H93!Mˈ�Y��Atƻ�
wcE��AL����u�P}�`]�b�dѮF��a�PT���A����WMpa���[ek� B���՚�_Nə�pkf�ayN��l�ʊ�2mn�e��d�H�j����6G�X�PHQ*!4݇E"����-�Y�C&�-�4��w2�<�6:���Kk�p�4���8�� ��V�%K
�#Jl���]�*��w!����d�mR���U]G�S�4M[��w��P2I��ʡ�X!���s7+l݊^U�� ph%e�{�&^,a;ބ�jﳮi���{Z���=\�o�b|s�]tS�ic��m��2������Ү�Y��<���"�]rx5+ժ9Zوʵ��	�tJ���Ъ�ܢ�P�Ѻ�5������q���e݉�T`�B��"��0��fJ7�&�u��r!2K$]jq��x�H)XŌ;�x�A�ͅK�Z.��ɴ�V]V�҂���2�[�gE���@��K�CR�.������N��s^�i���ۙ����o�Y�F�6�^d�כP�j�]�&�l�&�j!e��U�YN�!'��n̘6����6�c-�؛�Pl���(�hK��彤��I�����̫����Q��9�c )e^ə�F�����lS����Knd̓se���S�Cj=@�ƶV�n���BUA4:$츋���E��4#�+_��v3��D�`}�!��/6�4��PJ��NE��=�,�1��L��SfX"VZ����0#2���yn$�'�h:N�h��]�Tq�}F��''s�/!w���J�)aWSy#��Q�"�S�+-P�ݙ�i�. �Dǅ�a��գ�����G��,��X�2hg�'3�d��MF�I��Ţ�:�s3&-$���ӵB<W�:F�`���F�,�s&�n�V�C�e$%嗌o!�JJ��,W rS
��Tli�wK�Ն�U��2��1*JD�uj�,�q�@�",]�6��r�v�9t�!�ڹJ���+zҗ"z��:�m��ca���FnVV-�d6-��h)I�[J�4�c�(�"�R�v�S������]ФX���Z��4����Wz���J��+Q�ʶiǶ�O��:UZv�v�+2u0޻����WM[��ȡ�mM���Y��5�*<�W��qw���X�0��֯g_hs��$K�lY��+6�B϶n)����9b�j��9�c<�ܦ-�m�5H4��.����]�#1	�*�!�4W����[틐�9C���w�R��Z�=r#Z�	��+t[������jա#�[5ynL�� �����)��5U#.�F��,�ܪ��e����ip�L<�9pg>E7E�������ᒼ:�dI�v��ܬ�dg��Ԙ���iOw\�eZ�M{��oڮY1T�]*�E��#6�UB���$��Ȯ��
���hz��2ǽ�>�j$y��r�q�����{�ܯx�w;}K!]t&G{�x�#� 2#t�a��m��6(�_l�U��c�V%sS���r%V�d��sE[�Xڙj�Q��y��TOQN�>"��]]�R��F�#��PԆ�t]��26�Z�z������t��S+,#j;���e�X���wʠ��-↑��Wu�t�;w+��9[BQTeGN�^��r��m�k��aa�S4��D��&�ƭ�y�
't޷Q�QL�@����w����)	���Mm0� OUm½����:�$�w���{V��Jj�$hb-��Q��B.��ٙ3�vƯ8+�d��(č_�imdG�ܷ4ZՁ�Tu^M�p��Q(��do��tq�j���� \�g���l��=�#�H�U�A�j�����'Dm=	$�w%����^l�<^�L�!�O ˻���:{����#�؉R�l��U��~�&�F��\�覬%���cuZl�ۖ�jKQ����ق�`�������=�v*f=���b�� bj�R����r 1� ��+s��锞���;����X����H���My�AX�ֹt���L�&[	Qu=�!;��|����|W#wv*���_2ku_Ф#Q7{�m��\D�@�^��6�sia�M	F�	ڵJM��.�1���j�BC�Sv+t�g	:r�(����˷/� �35㽜/S�|��V��C1�<���OVHmJ�2�O��k�]l�2v�Xz8'��!���s���F��kY@7�g4�7vd#m��o� �Va̙�����i��,�ʺ��r#*�Ht&��%�J���X�J�ٍ��VI0\�D��U�v��R>Q�ԯ4���6��&��:*eKz�.Y.�]k&J�����`i�g�jT ե�6�6kf;D���dJ92�"�Hym��{S|p^y=�3�P��ۨ)�ݠ�<�n�X����*���L�kDhL`m�p�3s6�jO,�D�y�EsAj$�MMcM��JۧT�1^�US2L�-������(��4�xU �A�ƨ7W�-2/l�Ժ��޶��-n��A��ۙ�pT��!h2h�n���j�^!�l�����(0�vu�ޥ���Qi��Aֺ��̄n3n����&�Si�8"��pfe��\���������C2�BU Z-MGuKh��1��a�m3�d��gX�2�����{��
y`掆��[�t���ͧ�WL���(8��m>9�v�`E���O��.⣻�y�t>��o_=�ǰј{��.q�Z�\`�U/e���m���R!zh�Bc����d��&�:�'M�3%�Zw�V0ݸh�C%E�
k\v�Dn�
��9��d�]n7��hyH��6��Z�U��:�{��(ϓC�⫭`򼔏%�RV*�n
p�l&�b ��D�oQ���3u�J-Y�٩$ZP�+�[0�Abu-;�z��f+u�d�IT�:�N�H�ܧ�#8q��p��-�d1e�6�ѹ*k��e��۴��R�n;������wE�w�3+^*�f+#�͹U# =w,�uI�S�(\"�f/X]Й���*�C�P*��Bƶ�����5���$�b#@i�Sun� �Z1��ٓBŚQf�JЪ|��7;����N�3',G��U���t��+1*���YY0<ݣ18����޲��4D�\�iY�mIc�$�Cvf�ZH71��l�4��bK�V�822��(̗C4����oim����[�p���/cT�[̚",�͑�D�4�[X8NY�h&�j�� �7�Е"ˑf���^'e6碌�%bx��p�\j�[�r��b�<cU�LEǵ��d��nXU��F��RPU����nY�����B�\���Ҥx�m:�ݦ+A�/qV�ߧ�iгoT9L^�k3CE�"l���N��i�.^�Ǻ��݉��sejJ�.ط�U�gkZ����j�nk6*���̷$K
{&J,Zʵ<�u
�e9m<�maT4�+�����1E�4�Y�e��ji�v�c*;3!�Ui��[�ȷ�`9F�M:�i�(f�pm-��h���)S�b�}��[���PKv���̭ǀ 5�t�W*KR6Q�a0`W�m��m������e<���aֱ�mCy�C&֗�0�M��*F/�ec��U1���5��c�]UK��ὔ5�j����⩬�p���37{��qp�v�.-T��b'�M�v�������M����`\S���S`r�ax�=t�t�#*����n[~� e��n�#�\��Q{.��j�몷�nf���b�$�MF3v�\\�,T{�)��B�Q���<	ϭ�����y)^�4n�h�U�ЦyP�b����xG��/SF�+T�e��l���vR/ޝ�n��̪��@i�(�whr<���Ơ��=t�B���j�'�(<�T5ւ�Eh�mI��{d�Cayk1�VCyWT�	%=Wjj�T�%'���Y��E$]�}kf �J���QE���_�AV�^�7���ަF�YC��#�a�WX�H����򖧹i,�y3�.'� �&�W��\.0��^G��v�b&��*�K�Wyb����
��u�� N'��@�^YC)hջC�������Vr���aRBA���m&K��e]<�]��U6�*��A�BHZ����rS"8�+)��b�Y� -�ʵ���B��4�j��Ḟ�*W+�9`v:��p�H�Jm��:�է-7�r��aku�PGrQ�I2h[Un[�́��Lh�`��U�ۖ�m��m���7Q�j�c����T��6�!b�ToZUGnzUX���*�6*������b
!a��{�Y����WM�Pm�OE`F����Z��Gmj�5
!M%a��:�*SV��G3��x�Ek�Wx�U�2�Yײ�h�i���.�*�e!e�X�Ӵ��,�cOc	�������a��b�M��3if����u���u`^��{� ǹ��	[��Q;���o3�	Ř��8���Ã1o��6���4��`Ma]�$�V��tU�UuUU]UUUU*Ղ�����=hWO=���T�pm��UUU*�r*�UUUU!5Ti`��U������h
U��+�-UmmR��UUU�UU@UUUl+lԫUUUUUUT�UUUV��*(�`�
��/`A�KS� �Ӻت����ճ�:��V�v�Rx)v�j�L�,�1U]`�`��n�Ԟࣂ����]73�C�M�A��7]T���v�U��ܵT�]At�EQEW!5VܫUmWTj�5U!5�*۵U��
�UA`�;kۮ���љg�2m��6,t���>�ն��u�LR1uۭ��m�p�˟񭗹y���+�r��Rc��}}�����-��� Y�1+�������j���W�M�M�Λ���3����9˭�η'��n0�f���ڴ�����Q��r��1�v9'Euj؎������X[��`�M�*��N4+�ԩ�YA��Y7<�c̌[y��4�=��n�ŗ����lp���:ױ�n�yM�<���]����\m���Y�ܠn4)m��g7ê=�n�p󷁍��<�gl���T��5��1��uw<�oBI<�[c3����۬/g� �`�9���M۲u���3�5�.���^���q�1ޢԽu�a�nkɇ���1���C��W���`�{��׏iQ*	ܝv9�][M�86��g���n8v��G���m���g�o\����B;�w%6.�V{vgw+��ob7���e��9�bF;wo+����}�/u��z+�c��o1��m����.��;=Zt	��F!@�Ҳ�	����k�룷���s��7�����Z[g��[��#s� 
H���XhP����a�uY㑎�j�t����5��g�\uו.'k�Yy9��q�X�'��������8����F�;��m�7kt��@�nŲ~2�۞~j�.�,�a�5��s����v���+��s�}�I�l���J_a�l��`�u���7%��^��KϱMync��:�ڋ���� �u7��qY�F[7;F�N��l���Wus�1Ods�z{1�6�0N��9�6\�v�!c�����0����یgle���y���r�0k����)���2ac��9݂Y��<�v���v�f^�s��m�t���O3��]"3�n-�<6�y��t
�뮝>�ww7WQ���u�X�t62c�u=�b-d㮴�: 3[-r:��C�A�̫�z����ON�'6:��]�I;De䋲q1��s.CB9/3�Ct�0{f.��^-z�pqX<;�ỷX���+�wN�.lkD�x�_O&7�>���7a�ec�IϮWX��>5�U�0+����N����݂�q��`[�F{]n����w3�k�i�Dv�*ݪ�a�࣊����R<$'Qd�4c��=c��P��}l������O�90�.8��kqzܘ]������&��":��l���u�5��Yzӹ.�l��͵]�l�lkq�m�e��]��u��2���p�t�o	���Ѓ'��y�l:�d�0@;m�x�(�$7��}��n��ZwAv27�Nwj����n9鸎8���vmsX��{cpF7S�Y҈ ���{5kTۛkvvM�M�]����D�q�G�.������,h:z��l��u�:����W.v�s]]ץ�S��p�<4�^wi�؎]9{i{lp�p�Ű�]cOOgGg\��c��S����w�k�v�؞�����i�{
#�2�^dާ�Iy�v� ���Q��-j��vs��H�ݮ�{d������Λ���)u���=�����n�S��Y繨8L�&�흂ѷ�7gתAz.��&v`}��H���h�����wd5n����%��p<r�O/]�΅�(�n�u��8 ;�����?_}��L����6Ƴ/7#�m��f�xy�k�l�><7�m:��C�;��d�ڎ��q��Xݺ�v�v�0����n��|s�����u\;q@v6�S���^#��3�Z�yS�.��v{T����t��<���C��5�� ���$�J�p���vC����ꢓ�'N7c�Ʀ[��gk\s۝v狜�Z]��[�2��͘�����ε�#<p؜j������6�{[��۞����Í�ܵ�(��D[-�u��Dۙ�c�����ڌk\���fš���`�����jA0��.�\Ҿ�u�����#�5��9[�rX��������;��ٺs��C�nj���2�g�o:��Ov�����#cz�Y����m�fmԏ>���ۣ����p.Է)'8[:����l��:-�9�ъ��>(������ur��+��x���pN
��}Fq��e��[69�ݫ�]��&�n1۞�*n�;1��M�{\8�Gi9B]�vҧOv8,�d�Ng���ʍ�B�\�3�8�מ��۞{<*��&(}=��i��3Ѹ�S��]r;�\j�;�Iq���:g��h/\u��	s��v`����"M{=MF�os��On$7nQ���Y7t�����d
�a�q˽��?�շkYwUՖ<��/[��v��{9^��˩�G8�^��ݜ��i�(�5�*u� �>�;�g�z���ۙ�#�ְ����no3�m���Ɲ�C/Cβ��OfD���g9�nu{v��1�Wc�2�wlI˸�O���T�}��sv�X�iWs��c �8�Np�8���ńrպN�T���,gv�%��<�v��m��h��=��:㜧`r�vd�n�@��6�Y���ÔN,�����OW�H<t��jt[�n[{rF�5�:m�q�1�3��Cm��mLnM� I��c'u�ѵ�T�4�1��hq���iy�,7#x�lRY+�5#m�����OhM�}/^�§o;���h�	�m;<���{���=�����_=c�j�e:�ݎe8tK8q�^�1��"�6�v��g��t�٫r=�R�f�L�.�ڸ��m���u����g�Pmz7������4�iÞֈ��.v_:�u㋶.y����$x��ֻ=c:�:.۷iN�جVL��v��t���i��ͺ�R�T��s��6w���烣�/C��\�'�qm�ᑁ������QζיA�v�n�xPۑ�]A6+���gp<��&�d�9�U��6��2^1�W����3�ck�qz;{��J`�m)��q�pw0B݁����
Dn9{Cv���=�緔]�=8˝�y��;6C�����[&͹hѭ�θ�9�M��ZÃ�)�u���[Z��+����v�ݓfw�yz�:b���Wl���Fx;tU�q��s�m��7B�<�XZ5b4�:N!���;���G�<�d炆Ϻlm5�+�Hw
�v���\d�=*v=�[h�m���ɮy�sh�#���<��HEۡ��r#糼k�㬸�x�y�:�-G ��k�7n���@q:��������-�;c�I�y��lf/ �����6�8�0���"t�}W�,�4�x�w0ܝ�c;q<߇�)�|�(�S�뮵u�=�����=�.����=&��]998�k�<��QXy֔���3�֮��л��mݣ�lc:���;�]�3<\���3	��۶E��������FsG9C�i{/8p�a�]s�7U�����a�r}vث��l'[�������kd��$�Yy�,��1��7N�v"���x�N����J��x�=SkS��[�����!�q�������dɏ!��{s׭�����oV�=�?\��|�I�6s�[�Sx�]�	�f��g���v�z;B���NSOc"��� �Ys�¦�r���huM���4���v��j��1v�w���k�.:�s	Êy;e���=��x9�ړOG���z׎t�!u�)�}��!���k�6ۧƹ0w/kb��״t���#v�vU�Z�pcr�V��՚.�V���:����ۙ���L�]ێ����=w<u�r��`���1�k�K�*u\��=e�n��x�s���X��zM���wl�_}�n���6����c^��&ޞ�L����80��TX��۴��1	㗮���#׶ �*��[]��_k}���T��v�X�ݎ���sK�np��Z'��Uۧ6����tn݆�7b�:��~�}}�B7�<c����Ŵ�Y�j`ְ;�km���ۍ���.��jM������ݎ�jy����6�f�k�6��&4su�;uN���k�^xe����/	��mngG�7�����895���{F����.���k����n��`�N��l�k�m�k���n�l띹q��X4m���z����![�y��e��I۵�sK����9���*i^�M��; �6����M�,����!Q�� �W���Q4㐒���;mܙN+]�-�cB���\���:���j�A�'r�zm�Q{�ʬ$�����87�-��ۭ�v���#��r�C��d5p���*�N�i 2ۨ�����=��m��J��vC|Qh�Z�>9m�	�Lm��e��Œ�,K&��g��7w#4����^L�Yݺ^��(���v:ڵ�@��w�s��bG>:)��g�o�����q����cb�#�.Ÿ�!M�9�^9ܢ[t�p�v�:���CS���mQtin�%�4$5ӹL]CT�ny����/�v'!{&�9�6\�m�+��nm�u��rwunI�.(���6�q&��n\۰�sӰ;X��˷�m�wY�"�lP�t�)	� �L��Fz�9�]yƱ�V�q�nس[m;%�v�c�7u�wp@'�/�w�v��\v�ڴu�Cl�$N�C�Z���('\i�2h�*���/"�e��^^{g��Y
mۅw9)�\N�[t��F���	�n]��[[=�^��vSs�f7W����-�u��i�wE�<�;��\;�As����Z�Ƣ��3]�%{�;<���UG'�i��jb��4�l��ŵҭ�r�b�m����h��<���@-5�Dݲ�1$�f,�_�,ĖbĴ%��3�f,Y��,I$�ff���fb������w���R�9�E�u6ʷ��K�3�*��-U9l�ޙ0J���Z=Z�uv�v�.��PnԮ��v��;�^�L��\�Z��x�\r�ܽʦl���v�#���H[��r��K���r�]�ӡ۵�^{/��.�E�H�幬��m���O;R��q��D��=��X�u�j��ͮ�C����\�����pz�CGm��`m�i�m�v��ב������E۝�v#�^�h<t]q�y]�)G���J�mg��,ۋ�nNx5������5ƭռ�۳ی�x���`�oD�T����ZB�s��{`���#<���,ͬ��h��7�	qە7i�=��P�]\��A�mŉ��h=srp&��W;m�s���V؃�.�q֜z�^+K�-�	:�N�����;`!Nzp�Xe6��C^;mu�pu8{]<n�*lC��\Xӭ���s�f�v��͞�)e�lnJ��\��۶��Xڣ@5	+��UQ M�%N�6ƭd��n����p��m�F���I���2\����RmX��c�;���Z���j�۶��n٥ض3sn��S�ϥ�OC��p]� ��ч��9�˸1WI80���[c@��덒!�m�6,b����}�b�8<��;8��ێ�=%�wV�A�+Ĝ�<d^�K�[���:7�2(��E[>v��(�]���*m۳K.�t���HrA��-�c��[����*g�p�RZ�k�lZ���@�i�7={d�dQ��/m�=�]`��7uk�C�:�݇B��'�郮�gm�� ��]������;9�z;��uշR���fܸ�=Di,��L\����1u9eONjfZ-�chj-���n^]�;u@�یv�;��w�t��nv�聦[��nv��]�����*x5�ɰkh���	�x(s�ã	�	�)��θ��mv�K��u�LCB�u�OӪWX�&�N��Qt.7`*��j�rhݶy�M�ni��wF������8��9�Bử��;��)5��Y�`�KZ�zLQ�A��n��ݎ��X���ث�Mٍ�C^㍞���t홛���zb�a�mp�X�I�aִ��co�睮�8w,�=By1��)Qa���![VPJ�E�^�����Fi7�u<B���h�of./�1<���{N�k�v��q�@sn�1���r�>ő�-��磉��<eN��\s. ^{��a�ps����>98^�+�;!�y�r���r��y���,���?�4�i���;��=��L�M.ďN�#8�`�dx�ohB-C:�+Vq@�"�0��`�$4jg
3BkP�E��u��NX�-�p���(	 �h.��64�C{Quu��4A�Lf���B���	׌��ߞ�F~ ���Ez��v��j"OM�i�*Ho�&��=J���_K�)#�WB�_~��[Km���5�u\�~%b-lWWP�P�)\\Mxky���a��so�J�Z�!��2����q�Y�.�!ٚ�'�~�nZ:0YŎb�6Ǘ�[�Z!���\0mt�Llk��oIh�\)��*gy	��}s�I�9ꘚ� ���}փ�`u���{�9�V�WlV��,��#M%E�+�`a�h�Qn	 ��Z;�;[w�^Vȑ��âP��}�x�i�]O�e�]kf_er��2̐�����1�f��=��u0��+9�(ӴQK�<��ɠS<�2e�v�<F��5v�Շ]tu���K� 6_����d N��[8=|��τ�pwMi���m��Ƙ�1}�qkA�lb��&iT�;�z�E���}ll[�5�+OObP���Fߝ� �c�ōHa�Dq�|��CL�_�������_�(�B�-��Z�7a�EA:�}�����ˡd4hn���$���r��W���:�N�<�YN�Z��q���q����*�$���y"NYB��@(��0�I�o��
8~�_z`�	p Z��3��^k�;DJW���.�׏�A�A.��^h�<Ge l�o\0��u��1��1d����!�]���u+,�F�m���B �I��݂U�p[�EE�6(�]���(Il��J�P ��Im�+�� �/2�����Mn���������y�2Q��E�	[@bC3mgn����Y}W(���+Q|�]��R[3�ƴ&w�ဧ��-m㕭>4C"�\�wn�T���� ��3��S�wU�6~$�{!D_����ُ��d3�D���GA ����o���"��%7d��G2��"�D;x�wX�չ��\vk�&� S�Mhi�@�m4a�9?Y��<�^���S�`����,��l=�"0�Ƭ$i��Z��������}�8DB#+s�{PM(��d,��t��Q}�5��8W
��Ux���	���"�y�R T��&�Za ����C�g�E���뾖�?#�;�ʂ��L���
#�,�#����*�|����p����m��ۗe�Il[/Y��\2�A	��Z�$jL�JR���l�$��[Z/S��t�K����3[��X��K��=0.�f�jMm��Nv�e���E_}��3��᳝&R�S~��$���q�D+��=���ú�x�|㲁��X�0�a��VۛB��M��_��'~��{c�U��r8�i𓼂��>umk�-�F҃�]�h�h��vWV��z���5�s��R�iR/�mԊ+mz\�*�0(���� ��5�
��sQ��ڞ=d���UF�
Mi���� �k��<E�q�>�}s���Z�%PY�
�*��RF��!��ճ��C���jk+��ov�=�OVa�R\��G�:
x%T�HWd�,r���#͍���}�u��A�!��L0�b�z�m(ѭ(	__Z�y�s�k�e@���~�q�3�k��'��~x�f2��7���	"�J��w��x�e����P�Y��DF�!9#� NN�C��p���$�e}W\�%���T4w��KT>��%�!{h�o(�'YS��5���*�[�IA-���kFqF��j��K�7�V�_@�(���HҏČ�u�%�B� h� �ԵJ�Q �h��"��R�ψ��Ĵ�@}u����\j0�E��Ɛ��UH㛥�=k�K=HY��呧_��E$	U]��bO�5��fzؒL�,�@ageZ�����Mdit�{6�d.�U��B�cu��;�iፕ[��r�����&sɵڢ՜4���B�Owu�D��35�������%E~G�X|�|`�!L����'N�p�@��Q�<_l�ufJ(�����jr�D�i.|��#��Es���ju��ՠa�s�u�G�ii�$������P����(�rB4��\u��n�;=�v�t9Ľq����n���W"�ӣ:��h�a����o�o�ҭ�(���}�	����a� ����UC�}d@ N 6�}������ҏğ��e�B�^�|h��4�*�q?���17*[?��3�~��À�6���q�]1c8��F�r��։��X 0F�B���-�u��G��4-}f�ְg^�U�\>bO�gF��Z�b,�Y��5�ر�پ�=��F$�_?o�X�*=�؇����"B�}f��(�L@B?r��O�~�#+�[�F�A��Oҏ�A[�u�F[s�|(ikc%��2N*�ߨ ��#H��*_1�f���O�8<x}���rܧ��Z24'����7��ؤ��TI��<h�%��� ���!�	|7���M�Z��}(��#�:��/�^��aGD�";����A�M3d<ix����SAUs$����/���B*��',3E�X�+u�2�.�W=Pf�\��c�xS�z�䞲U��M�
m��_#J �smz��-�]���m;��j��ӷGٮu��nv.���Ce2`�t!��e��3��7a�t�I�٥�gΜ�v�Gn��c��\'#Ƕ�ٗ��gz	�۵/����n^y���	�<n�\���Z����;3�[��u���a�;��I
p�Ŷ^:���8��܌<"۝lq��G&�����8v7}yn������K������j�K��ٻ��Н�}AO=�[��ltn�OQ�N��.5�N(!UH�_"àT��}���A���pՙ??�(f%�6�@bD��[凚�a��E0�D�z�1�2��ѝӅ���7�4���wn.�����sZ{���TqD�C"�+#���#����0Q¹7�u�"�<G���=�F"x���cS�Ñ6�����$9=ҸA�{%�.Mkn ��4�(<�UX�PvT�.6���}�T�doH�E����A�2͟W����H#N}*�-$�L�+�o6�8Q�)ʖh��V^p�¤�'�@�H�����z�;ȑ���}D�Q'!@>A>�(]�O��=�_
����B�$�G�(�H�B�ǖ��]vu�����r�h�H�Aw���o�l���l���lRۛ��8�f ����H�A���o�p�*�Ӌ-��gO��78���[�("�0�~H���1C����8��u!�3=:��>O�7!�%��2�xȫ����4t�y���=�u�!��V+tK�pJVy�4�͖����7~q��6u�Qb�����@�\��j�� ����������2h��d��i!���o�e20�3�M�&hʀR��C��S����� ����}��G7��]�z
/�T�ߎ56�+˴8�޼-�LB�[βVX�y�a~����j��SZ�U^ta'*C��*��.Pdʳ�^�"� "/H�H2
zy�ۋ���G��
�H^mݼ��X��`C�x���Lr��Dʌ$cqW���,�W\����|�BxQ�@I���t����}�8H<~��QF�6P2~�ޱ1Uv� �,ay"bք����q�ڄ�#�΃Z��ǾU_E^t�B�D����@��h�h6���P���>#N�,�u��H��_q��miX�Q#�I�D�GIm��r�]8sM�2��x�D�8&Rݬ�x�:jl0,�0`o�9�-���A�G~u���x�`��bV�p�q��$"�
�����p3�9�q�=�;]d��%�����^-��]�.gs�y����o���%u�>?\p�AK�g%`p�yC���d��$�@��#�hNεB����D��}uQb���sB
�?`���z�'��Ǣل�$,� �6�	!�4
_l]�aɛ�?@��"�~�CO��ޡ#'���������8hA���,����@a����a�(���Z�󃥠���Jr�u�C�Ԯ�2�ҫz�8j�J#oʊE���[,�c�[��E�jB*�D[�TRVlo���ž�ӕ:��lH��в��2���t�[h�(����æ��0�|g���Cd��~z�����ܪar���m�GB�g� 3D	�;���]I#
�ɢ���9�NGR��iB����I��d;B�-�@� V�r�G�H/ 4-l���K�i��$�h\�!Dޮ�vH�x�B:a]1�%�'{��+�hoFk�k�~������Mv�0��y�k����y�ؗ��B��Y��A8�F�4Z7`ܷOn�����V��i�I���t��m�~��ۅӮ&L���%VK;�����y�_x���$�@��k�G����B�2~R���ض��l_7��ut�y�,#z�g�fX�eq�d"r���[	�M|P�	��}gN�?#��M�T,b3�5��~����?kMЅO]��ƀ�P�Ct4w�����_ǥ�ڶ5iP�xV�f&�
BTjH�^ �8�h�<�d����|uv틿u
������S����tG1m���(!(���:�x�ژ��
�{�Wi
Y)�J��6���ܚ�IV�sq���='�r���C9��)(Y&��ݐ9��QTf]&���z������>��:��~~Ք�n��aۮٓ��N��,���ý;٥�n:E��m��T���j����� ��!��4]�P_f�v��<#�bZ$q�x�4FD3���O�{y,��
F�2B�A������@a�Ə���n_�dm�{(oc)/������$A3���B�"���J#Uc�0d˱�jo]v
Ųv3�,��F��Q��
A �>�Ds���f��K���<�m�[�9qAۛ����%���s@|=:g¦�w�=-��l�a�06AD?s��^ĺnvQ><�ޱ#P��W@n��:E��B�Bh3����oϤ�6RMȘp�&`�#�IG��&x���m����B��*
G��Y��Q~�h�6C8A�+c����U3~�R�P�6��^�lϳv����k���Tj"�mQd�($Ch���Aǰ0�4EE|�X���l+�f!�R��ڧ�
�D5��՜���Soj�~Q�]xՈ�1�g�m�x�tF{#w����h�������HKC՞���YD��u�C�|��l��\|N/�y@n���7UbO/����'A[�r�.�8�V*�r����[�f��_�.yb���0����5-NG=�Aď�H0�9�\�����u�hf����G<�����Z����~�> ����u9��������!"�ܡ0�XN�V,B���ܮ��j2S�%^��@��jڢu����|��ۃo�N�5��,�X�K��.�=�8�L�Q��R�����������9c=��s�T�"k�9�t��;;vY���ț`�;;D��=v�\>��ԣ��m���=��c��v|��<n|p6�y� 
�`2tu��C;Ol��'�����xƸ���9��pq���1��c�+�k7:��]���M��8�'��z|�`��,G)�>�p��[�qm1�Jnd63��ᇔ��[�v��cpt�և�$�	ŃNV�i�ВW���N���3_I���D'v����R��t/�� �#=���]�SڇOV6��},rC���4�� �$ͦ�-/?�ѱ��D�H �t�_r��N!g�K4��r���Bȳ�.�'�A���DB��z��Y���_��q_t���h��s�����6��4� S��bm��-��*��Ƹ�[��~�Z���h�!���ڴ�b�Q7wd��S�@`�ҬAg��T�����7dv�Ҭ���k�#��P�RT�d |�ӭ����s���Hx|�/���ԥ����?�ڒ�'a���WI��a��K���CֻP�gZ��l]3b��4mG�[0������ e�Evh�V-��!�Sh&����B
��U�A
�'q0��~=�;aIGǫ�Wj�ҁ'�j��K�����-�K��gCi�#�h�������X��tkk�Խ��0tnp�N�s�Y�cRv0�B�ۭZ�)| �}1xZ�}ׂ��"�BH�}F-/ԧ!��	#%��E��%��*aZ����~ԉEof�Na���-��m�Z��l�L(��4��q��{ ���;0�S���hE���O�g�S)j�l;	��鋞wc
�՗���u�ƙ��M��Y�b� ��%`��q��o]_Ewyni��D2&�Em��;�}���#g��ff�$�9"�X#��D�	ng�9�N�!(������.PM����>"HgȂj���$Q�B��H���F�DLl�~3������d�Q:���̴�#,!
%Sb��'q쯹+����_�h��Čڥ@�d�����~�R�ŧ8{9���vݩ�y��Ď�m�#�׸���OI��@���ܳHB͐�"�f��d,�wqk�>i����j��9�&�Q�	�Bm&$�ᝈ;�&�gl_T ��%PoS!�;��fj�޿Y��9B��%�֬Q��4Ҍ#�z�(�u8%챦�F�����Í�<6*�q����J�5�`�Q���Dn޻;���&���թyq	z����'(�\]
�t�_E�x"�h=��i�
���Hu�M��>8�Q�� ���S�ð�Q��dv�D��:�I IGQ�D����nN���%��8|`�CHPಟx�� i�[;.e�*����:���0�������p���ОH���s���x��_!BE�)2�.�gw�m�#��e�K}l��l�6/#�N��8b��o�Ͼ��,�*$xx,m��S=�΄�\W���s��4]�;�;W5E�������)ͦ�Rk��Q�kJ����hk�,�Y��%մ�]b���7ٕ��#��{�����CqZ�h�ua�YК��Qwu�-�IwD�5X��GVǷ�AY��-���gvQ�+�ď��j�=�+��"�-}!����w��q]��q�<�\�0�����4^�v�UPۆv�#�hJ1(���е� ��Å�gjv>�vE�!�ƻ[�A�C/��0�6
!)Y}ׯv�����-2�~S���Pcgo���Z�VQ,���H�Ռ����7Y]�Z�����|rX�u�̞{%s�,�(L��cՕv5u<H�\����T��J�\��v5�iՎ�u��ݩ�*}���3`.EcY���l
�P������fj`͜��1F�Qv;�MX�0�L���,����x�v���mu��׀�[�zւ0�YG+(;�'`5�e�9Ԗ�S&�L�c�7H�5Yᛱ_��W�����8;�|�����k�Jچ�U:�{�����P�i'��99���[�lQL�l��N���@�1r��;6���-�	s({����۴]-��`���rXF��_ ���*�FFF���zX��V�,���2�B�E/��otD1�2j	����}w7o%�~�e�/�4d&����貧_A=�=2�`�20jbv�^��r��%t�nO�tv��U�dHe�ET�q�T�̧|�ԟ�dxsk,A��f/�3���o4�ؗ���>1AdbŦ�(1b_��@�B�$ň1O���[ X���-��TX�b�I��bb����'\RQ��%�K,_����X�Q$X�H&�>��m���]P���>HQ !&%�C�Ͽ-bٚ3���1�b�&%�c|$6���bf/�Z �~޿iib�m���Ck�I3�♔��,B�#I13��ܚűb\1z5� ţ�KB�,B Ħ���?_s�.���c1�~�Isz��b鉋,B X�LLY�I�[X�6�/o����V蚳
ݦ���b�B��bf-����b��iAc ų ��y��m�ib�$�]2
�iQ*,[mb�'���TX�b�� xon{��T���>���e��Yq.skX�bP�Đ X�M$И�h@��X�bק�Y��Ě��f/�LX�>31j�%E�1h�Ŋ6��k,A����-bر.��3���L]3�(,@��X� �Ih�-�fC11b���k�����n;�<³�q��m��c��Jv�*f䍻.pY���k�nS���Q!sg
t�n�ww�LXĆ�g�PPI1b�k,A������_��N���It�b���<�b��bb�bGdJ4� X��.񥢋���X�b^3�Ab�F&bf�̆.�����ַ�jJi�Ō������-��1��ߧ����q/��/���/۱b�$I�@��z�-�������i%�� �񉊉&fq��k,A��&,@�X��I���.h~�Q�k��W�[ X��tH1��dB�.����itX�P��\11b�ߧ߇�� ���54��[I�#�b�KF(d3�n5�I�b��s�X�fp�b����3Fc4bL��LIi�-i?�X�b[�<�������pI��d X��&bb��%H,@�cY�I����vk���`bP�k,@��x�|�3SۿnU�p�%�b�B�c� X���w~*���PFF�S�,@�O�PX�b�����ɣ:f1b��@�-����[ X�f{o �-�����i8� Ĩ�\13�L��]���K,A�� X�|1&g�sޢ�,�n�3�-��K�4-	A($����{�Ip��g�x��X�b^1j4��ňB������ X�vw��J��b鉋gD�FDb_X�11eb��� X��{�_�	hXV�h���ٙ��X��L�� X�m/����w����,��ę���|f}����K�b�	3�(($��-�����	h���X�,Q��Fo��ܺ��b	&���Că1h�PI^5D�B�bء�Ęŋ����ib�y���S X�b����1|bb�	/���.k��jq��k�ׯM"y�M_��3�D�MӾ1}y��>�^t�ܝt[�.����;Y�qfl�7�
�h%f�B��^��B:�>�L!�i�?�{9W����,A������� Ġ�T]FAb�������-UJNJ�����3�*�(bf31��$.����,@�b_��~zűb��� X��LItLX�bL��Z13�b�k�'�?����fw��Գ�<,K�H�K3��IC3���-$�$	4$��f�K�iQ,�3"�fŚ3>޽���$�t��,[1,|y�|�1(����_�?��8�r�ǌ7�2t�]4%έ���+T��7'ݮ��VS��N*�9����P������y�� ų�KB@��I�����������L�޿��� \L���%�c X�LL�`$Ŋ��PX��=�s��[8,@Ĵ$u�bbL��%�V5� �-	ǁ����|���ZX�lJM~����߿=[䙋�/��3?G���(f��ą� ��^1b�2��q���2�X�b�o��-�&%�c5�LJ��bb�����Q�5�T
�)�q%�1b��PX�k,@�'�K��X�%�ք�F����~��-��1�fV�o�?~���k�������bb�5w���I��bf#�2����~�� X�)�}~1lX�mb�kd�2Kf(,@��撂�������.�1���b��b�ŭU� X�b\11b�g��|��ZmŶ�|d �5�yb��|��>1&,A��&,�b�k,A�����VA�2K+���bر�bщ��bb�Ko豋bቋ,_U��v��ؘ��f/�ň3�5� �ƗLTX�%�1b��8�C���[ ��.��*3�����]��^��mo����Qb�k,A��&,@��;��ŏ�'/�	3��A� �P��c��Ʋ�1b[߿uk��ۙ�X�b�I��� X���ę��&,A�3>�[�I?Zآv�J�n�౉�&b��ŋM�\o� ů�]���5�����b�k,@�13?w���[8f3�y�ϗ�$�&&d18� X�J	n��Ę�P��G�&fC�Ϋ��,bbHm+���ض,@�1&d3��&,bLJ�;В�������?=bر�� �$�Z1H�b�,]mbK��?w���w��L��*�s�ZIlLXę��&,A��5��11bO��PX�b�����]�c�����[���Ӣ��������F|b�J	�%�c �LĶ3?1rfI��wK-�&b���Ģ��,A��&c3�i���'9� ů���-��-	p����P�PIo栱Y"�1&bى�d3/��zX�g�҆.��|����A fcF3�&,@�1bm�A���o�[2��X���1&&��(,@�	1&,b��bb�>�����aL&�И�ȉ�߳+����w��ac�u'T��ue�ֻ/7�VұRr�g6�Y�:�</nH�ٖ���0�h%#.$�����Itb�ϸ��_��z�l�X���<�۷������Kc����.�ɺ��s�l��M��qұ.1�Y����ڴ��c�^!�kq>���ݯnD���oUt,�9�j-��	B�� �f����۳����{T���<s�Τ��nukn�&�;[�\gũ����9�s����<���C {�O����w��ݮ���'�����h��ѵ8�m�捞n�<m�2�P��۷1@Ր#� %"���Z�-���b��?�b����E�E1&,A��m%�� IV�b��y׬[ X�,@��1A(,b�ӑ-o[�TbLų X�_��Y�� Kq�΋B���LϾy��� X�& -��'���?
#�Ol��`�X��X�%���u��hHi�@ā-��LL�LLX����wi+�,���/��F�fDb�&,A��(Aa�D�kmb�1}g�ߺ�vH����\���[ X�,A���1Q|g%�/ͥϾ�(�*bf%���ϧ�-,@�m�^11ns��=m%�b��@����PX�b�~��q Y}�zkň1 ��� ţ�/��,B X�13�#߿u],@��&b��ň3�cF+�b�%��&.ֱ������]8,@�I���L������o�w߾Θ��X�b�k=}1*b�bb�_��>&1T�RۚX�b_���[ľ�.�}�t�	r4���cBLI�1fo��u��/��%�<��	���A*,bϿ4�SIhLX� �����#S���%����#4E���}�ͭ�l����o_����h�i�������\�W8,?��7�)HB�Dd��a�)G���M�:l��%+PC"~ݪ�TN$��$D�����VY���KB�6��Ga6ϼJ�B��?NX�f�������-R�D꒨�.h��(�]��ť�)��ha��|(t��s2�<���&`WP�h�F��-x��1eh��B��6�����a�LJ�"VM)l���L)��(���<[��x�-ێ����[k�ڵ�9�w'j�n'-�[(J� ����,e~_�����<Y� �
�H���Ȳ���O+�P�L��D	k�v�=�%����&q�Iբ(
�|�����M��aT�7ˠ8a�KEDb�Ҏ�K5i�s�W2}R��s�R�i�6�H�{u��p7:�x*R[�n";���[�Ӂ.���<b��6�*ǗWu��:٠���c]�)�Ꮞ,���r��mDJ�&t��#���#F��Ϫo(B���!؝��0!]h���"��ګ����D_M+�q��E��-��b�0��D}
/��wҚlƉLp����u���u��)��G��p��{\$S��D�������q �̗��zX$�L�H6���O�m2���T�)�(�c=����0S���\�P�GM��!�:���&8Ql���?��ѵ��@�rF���뀯I.f�s�!��q%�2k���u�cv�X�*�[l���`<'����`�!WۗoоX�!\n��c�O/��i�����@R�A�Ο���V� �JG�Q]��~^�'�7��~?7AÄ��;l����4$����^:Y�cG<kf����V��ldcr����~���y��k�3��b������%;	��ED�%{�]��C�:��|�yP�VM�h��A\�4-bl��a�.�H#Ԭ,N2��mt_S:���S{`�F�މ��(Y#�F�7�? D�zD�����!b
U�%�>]s�Q��"M���;};u��Q*�ArjZmJK,y�0��6�����V�hT\]yG�>��Η}�[7���x뇚$xAf���\{v��1�׹;:�2i5ǶRC�l��nk���9Ļ�d�a����J74M�֜�N�n��F$(!�<����
�Bg�{��#_�����^��%@��Gn*j�u��W����P:�w I8���&�S��C/�!gK �����E�>�D>�;�O藻��2�'�$���b��RA���	�"�i8��8R�v���b��I����d4��`Y�gK�ⴘ���B}R�g��$bL�*��]�"ah�3�>���@�ÐBUP>��g���cIYa4��kl��bF��y�{O!�*;�7S��Lu�.�r�h��TuR�9Ge~\]�{�s�L靗��:�D%�֘/�׸��)a%Z�Ȧ��tq�g*D�I�)@��t��5$0�?w+�xc]�FԲ!��X쪭#�<���4QT�}՘���=���o"rdi&wMl�$I��V�%�
�yJ��8�p5�XQs~ܹ�o��g-�b� k/�;�<��We�ml�ς�Q��/k������z@!�E����ͩ|���u����i�����i񄐩2u#���';3��d
���G�'�c��T6�?Y�M�Qã#��1�BP��=�Ď[�	�:������I�}�
5�ӭq|����=�� �`�"�olO��X3N&���*�<���Cّf�U�ݥu3��y�9��}*'t�+�������Y����2M콴0ڻ����8�"^��@')��\���[Z��#��8�/Nz�6��_L��G�/�]��}<���+�x�|�<�D��]@R�&�h�G��Z�מ��6@'-���w;S����둱�HX�Rȇv��;�ԉ�J����%�T���n�\!�N͸�y�h�N�9e��ƴ&[�{�iqޯB�+��I�T�����,��voL�yoz�����:B?o�h���`p�#����\�*p����I�i���Z:�����Vb�κ�Ƨ�
���ȘS��&�R���u���D 9�s���x|$�qR�{�H	^i�]��4:�I������������UQe�9^�)A ���ƨ_SD�_#%E���"��� �<Qއן4�����ô	(��$b@��S@����Zp�y�'-�}���NZƥ��I+���;A��vtԔ�w[����ǝ�Q��$�8p��)v�PA��$E�u�dB�e�dA����"S*���|�|�~�Lb P���g�fy�#-Qoo���ہ��G���X���>AV� «�>�*�:��	��c�8�D�xើy�cks� ���f�ץ����q)�L[Cp9�=Fv�����:^�XSF>{�fb�+�w�v�+ۊH�ߐwh�O��^�� �y��78���̲x]�:�(�,\b�[ISIp��L���r<n:��g:[���r5_d��DԼ��d��x�[7`�]m�5c�2�n����8�/�s<�N��H렺�r�/;�\�\ޜk�d�ۍ�vwa�5�2�;�J��l�ʮ��/�k��)�N�=��k������=�>9�]]�u�B=4���z��bk����q�v�wnx�CL��1s�m�s�k�Йn��mۚif��\U�vk��^��Ad���u�M�Nȣ�Kb��G�t�Ŝ�݈�뫇��,�����=~��u��и� V���#Iq�A�A��R h��WE���ZG�oZ �m�6�?���A��xH��d�%��D!2�0�$
�ܯ�5�<��J����j諽���1�>l!�w�&����߫�F6�؜1,��}��Jhd�}���@{s�A@�	4X-��N��,�P�k�xAGLZ���Ej����]� ����d���t�zR1��Nr�!���9Q͉ {{�^����Ĩ���ל�6*԰v۠8y :�}ͱ}�j����m�`���(S%(��O{��_�e|p� �
w�H[�aƙ'���i�jj�Ew�h٪����cPz`�n��n8�q�RQ"N�DZ���vϫE۲Э���4Ϗ1�C�85|6[�o�"�4��%(I3��/A�B�GMIբY����9d�݇����V�!��W�nb�;p0����n7-�=L:��nE����6�?x�%�ӻ��@Cܡ�,A �����7��Fs6�hx���N��;��Ѣ�"����FjY$��8�V��
��[l����v[7���"m~+����m:�nd��~��>����*Y=jA-��Q��+c�~�S�ｺ݇��PNƹX
ht���9��\����#+0vL���2~���6~�@�e�=[�"H�A����@��Vz3���i�<,ծM �pO����MգH�k���[�yt6�>~k�>ӗT��W}�|��jf�8�a����mUuC\�&AgE��ynu��9�;��mV2��F�۔�&�{4��ޱ��?:Tg�,��oh��FZ�/�ޱ6I���V�wu�E]!��\�<T��]U :�JxYG�o3���O�T�1;nh�6hZ������ۦ "�4!?V�[�CRp%�C����T��Mt�4�3��X��	��^i�:)/7��xa�������`��˧�3Qs�����e�
dIdR�:�S�����/[!	·o;'2�lX�t^�\ێ��-u�v���m8y�e����4`1����W8l��v-B�{����K���(e]��V�_����)�}^}A�NN�+r�(�F�� �,�U�L� �8D��r3D���O��J��8�����~���Sq��<�G=�@dΠ�/�H+A2F ���7�w�8.!j<#��H�����A��	�o�J=��^8e
׏��U
��d���h0E8{�#��fW��tEEZ���]v:�g-�AU�|A�86�s0q8�%�w�7eI6^輦����8��r��6ٲ�(N����yf���)�4n�s��(�����twW��O��чOʉ��l�$ gט!6@�CH�Vn���ѩ�D�R$d�]���D�W���LˣA����%C�3b�x����J��!���q��ZsH���R���Q-����{�"��:K��YcZ���gK^-�\[�B"#�Aq��TF���U�ݘ�h�tڌ#���xh�9�����M�ފg��$�|�$zwADiS_l�d���Y1"9k�F��,4�_�W���,j�Y-$c��!�}�Z���"V��Xo1\��Xvܱ���i�IK�hl>p4�au��7d���Y�R��l�X3'D�_wJ0�� $�1�)f����/K���|b�6�|���-��8�w��&���H!E8(` D�Ÿ���ͷ��zL�T+?F�*ane���Ƙ����Ҧ�:0B}���]\�?(�r��*/7����x�kN*F\m��Z%ӻz dB^h>ۻvN��(�%�7;+��$�H��h�U*j�_A�Wh��-��;��V���F?YD!�o���u�#����+��q�3�ѡn��8��:Q�����x�EП։�����4~�-!h"�`َ"�-a.�Ez�ýbĻ=3�Z褱��Wr���"\������w����z�̘�J�7�R]�m��W��0�b�l��诼�. �Ir#�[fi�D�*�n���X�B��5Fv��ޱV	���ĉ4�	��C�}s��ą�D�	��ھ20�j���� ������>l4�'�3e�|��WV�Ϝ\Tu
��Lbl&ݞӮR�Ղݮ$��C��P/���L=u�ຝ����c����<ބ��A��ާ0�1}lc����7�� :sE:?��1֧�>�+��Ãt��%��q�o7ů�63���({�x�[#����ע��(��4�L��h?VY������a�Ŋ-�ej�H�,�C�r��4�8@��ZD1!����,�}�!�h��H�C5).X'��DlYc��l3���%	;Oy�G
��Z�Fw^	�y|��~�`��#G�ˍW�
#���A,���S��ic����ʝ��X�;is㍱G}�w�4���<)��ŕ)H��$M��&ʯ�C�Y�%f�1,H4��\���`�͂A4C+����}��\Lk��Zcz*��9+�w"w+rZ����4����k4p�\������^x��x�6�'|��$���"�Q1:/�ٖ��d�@H�@�� �����7�����Vǵ�Z��8b�S< ��h�M�C����Zc��u���pCy4��W�ﴴ���Md�^P�5�kQ���r��6�4�N��VDo3Ꙣ:�֋Qt��������K����v�X�9ۄfε����,S3�"�\�}D��$ʜ9��P
�tS;&��}b�v�`�h.�Q�!E9g�f��9n����mEĈ{�*�M]�ӓ�K�?��b���;=d��úZӷ��1I�)��.�t���P�k����u��Ʒ���k1]�v/�Me��ܘ�UΨ��Ks}�a��,�"�J��˃t��V����٪�^��*ųlK,\��.:��<���l�ޑ
��5R���+TY�ON�n9+%��׍6tK�3�4�����������5gT�њҾ_u\KLi�J$�9�/Qގ�vl��y}orrA��J��V�Ӂ	Hv�m\��9�6se&m�F�p��K%���Vr:�(_�V2���x���s���E�[9NN]��<�N*ŉ_M��w�|�1 P�Ѯ�;�O�����9�FĜ�[� a�U�s���&~/xzI�
Q]]!���+Gm�V�;�4k��i�v�H�Uv�ʄ5�Da��uV�+�"z<u8"�T�:t憷���ȷ��8���)�����7�In��t�H�P#��'�ԩӺe�2�3i�ll#F� �ۀ*�E�S�#Q,W���i��T�c���N��+�i5�m���w�  �o��@]�j��lƨ���ӷ�\���m������t�2���:p�����hq�.L�O���#8x�r ��{P��ϼ�n�۠}K�<v�[�6��o�Z=������s[f�� ��3���l]�m"k��&�\�[mH�xZ�3�֎ń�y�y�H�[�f�u�Xr���dcOg:[�웦��!��÷l�mu�]���n�3jݶS]s��S+�����×�|.xи)���]�����`&��zl9�G%b��8�4�f.�)�u���7L�Lӄ�zݸ7Xy�&��c]j�0=g1Ks����ڼG���3 [�$��_}�}����F�خ=0���`��H���e�.y�N�l���#�p�[e��^��80�u��=��Q�{���T�g�/uA�7o5�n�Fa����6S�lw#��@c^:�9c�v���92m��^�l�@#��۝���ݸG=�4F����@�e�������ѽ]i�'�Mcj�ݷEw�0��z��lu�;g�zn�;�����ٲv0?|�o�&x�aY�&�똥m)�n�J��t��fN��>���{v�0�5'���v��@u�[�Q^Ǟ�[q�q�[��e{Z}Vt�;]�"��g���{�e��+g�XVڎ�l�[�n4�+7����i.�Qd�ی�yk>�\�%A�\a��*k�N�X�9��͵�g�9����x�;l×4Wi���Pqǣn�7tr���<�M�8ꦯm��&�b�n�6�)g/W�n�g0u�..�K�r�]sϴj:��}}��j�J7��cx�����c��vѻC�΅�8v��lg���'L�����{/=.[RZ��9����W�7csGm��B\W�ܖ���k�e�.�sU���O�fí�z;v�wlq�������@P�v���9&4s�9sηsuc:�N��O��
z΂�ڱ�����:p)N�:1͞��Vnػ\�ԙ�gv{Y�ml��m�ҏ[��k.B�n�qv�g%�d���qp�:��$��z���E�j{yx��i���\�l[����y1����u�ϋ���im\��^�/9Aԧ;i�n��%�xn�܍�ݎ�tWG\<&��QIs��y��:��]���3*�����1���mB�q��H��`��5�����+s��xڱ����<��{v뮃��լ8�v|quٷtr1H�ݒ�]��/4�:�]��N���i&q�o;�J�N�B��Lj �`^;b�0��,�Ǯ���[�����_�o���-Q0Z����E/ےث$b�A&�f>뜖 �a��Ri#ED��f� <�ڞ�� ��C�XY?KvD>�$�<�\��ʟ��N'#2FтG�8�%|J_v��˪�!�c&6�H ��,�o}|�]���l�Z����8Q�YGb�^�oS�f�1r#ֽξ�G��ѳR&�Ȣq��ag�#.j�g��ۂh0�(�2{�L�$��4�=SF�!�$�$H��7g�H���a�%:��GS\1��M_*�򞤷���q`�F�憨	�x�Ҋ�21Nh����0�(!g�}齣�E���H��6����v�������g�Y$aҥ��sX�3� PI
��(�AYT�8B �Uҗw�a=Z�B��S�8n����wC2W��0Q���	�{=39U�{d3ɔl��>�Ha�YaS���~��>.��[�Z	�
�`�C��98��la���c����<f�,k[���^�!r8#n:'G R�#CJ���c~˦��X����?c�ς':4D�`��Q�Q}qJ���t杘~�.:�V�z���� �����"�a�⍱!����:O��I��s�T�חf5VVV�;��½#Q���H*��e'ݹ�)R�Fq��Uţj��T��Ǯc�'i��_t5.1T&Z��7bdY
j��A�P���4F��1���4�>��.�S�n^��a�$_D�4J0$��q��(}�Kq�=��M�� "�@�'Z&����նK���Aϫ�
<2�y���}̐C+�h͡�	�.��L��~z��0蹦l`a�y�;[hlb��.���K��<�F�H�U�d���V��{#��QP$�u#
{��P��$�CA�X-�"庆�'D%C�I�[>^v��mlmU���_�>�h0Gh�<L��>H�e���8[����B��(+��erf�u�x�9)��@�� }y��D����O��D=��_I}���C��ie��X�m�q�4m7�9Ѻ/=���b�S���t��<���ⱳ����o���F �K��]�!���DG�z�[A���Q�д<3�n�K�`�2��t[*�!�?V�i���	�l�Nq��54p�`��Z����=�JV�]�9+�� :�:�Ѥ�9�^��@i�n);��%�A$A�@�	����A�!$��Vc�JR.�fQ�h�|��md[�*�m�y�x_P����#4��RJ�Du�5)r�:=�G�9�D
J�y�~�� W�
̽�/�R�h��/�(
B��+�O�uϠǫr��V������ٰu1�Cz^��������۩Y�e�*A"7�z���D���9��Ш���/˛�z�5PF�RG�RƊJ�_���Dk������	���'�@��^�I��P�oGkr`.�o�/����f#��8ޞ����g�����!(�U�v|���Er[-"[ ��m�����3cExÕ�`���[��Ҕ���$�ΈP$���6o�N�=SG`�6�l�ߥ�]�G��;�L~��o��̤��6�)�='���O>^���b-����==�m��vz�G=n��n&c1X���r|:��R"��_n�C���Z����{s��h�vU�0,���{�fQ�s�=훔P
 ��_Z�;���nؘ�1 �xw��GS�`9%y��%mࡃo��*-\���%�Ă�I@��:�AY���>�(�:WP�C�it��Re ��rq#�{�:�MRj��H��|����ev�Xʭr�-�.����W|��I;^I�V�_(��D1���wR)h�N�Gk��$(�(M�����{�U�_0q>=i05���5m:�nR9l[E �� ������H����E�D��@�R��1t�:�`��Z'�(�r�ZT����B_bV��|����z:AR���z�Nct���SSD��K������qw��&$S�T/]�ט'.�+Qe�@� �o@bYP@�cn�"�}���ٍ�+n'e��(�9�����4�Ǩ)�h#�Fyq���e�<�b��b��`3���WĎ��O �"�'�D�7p�$��`�� �I��
#E%�:*��b7���Ql50�>�ծ��,2u�{r=:�:�V�z^;����:��͐ɢ�n�����;|{�
��~7�8�C�&hzk��8bފ6�&T��9ȕ�E��[�B։����C9�YƗ�b�}d GW�����D�G�!�_�����2�4f�y)$�C�ŗ�׹�̹�̐-Ǧ�8���u��L_
!�(�A��<�Eь�mA[�l�9�clZ�r�T-��O��<X$�2�$�H�PIK�=d����h���;x����6�~'޶m�#'$0+gĶ�^�����i�LlvD�=�������ǩi�4�H(�P������F�P�ࡇ�6�:l�׾�a����P�x��&M����|hM�e��U�	4��2ƞָ�|k1��l�ɇ^'��J��v��HĎ����	'>�7rD�I�"�D�ccz&�����A��]p���ڂ�7� ����Ž�|���" j�	��W�.��/��G�����0�X�J'%h���ը�X��gUj�'w���Lr��Wa	��d���P+R��y�[.oQqH�Lޫ��׾X=�޸�R)& ӄ~��+�Dsb��IƷ�!�:��[��q�⸞�y�����/knUӳ]e������s۶�ݺrj}w$��.��lQ&*ּ^KnF�G��J��;[SGkn�n��{h��f<��C�^n�pmѦ�u��NRu���8!ێ;@UZ����W]	zbgm��m�u��n-&v&��k���i"hݍr���<:��=���e���W(.{m�z�֫�4]�)��rNw�uB�b�i���J!��������G�?'���P����N@���6�|��u�W����0���tu�S���F������RYd�x�S��@��`V9Ga�ZzT�K�9=�#��P�.�,Oz0l���ɯ��]�F@���`-\�4N^�Y�o�׼Ar% ��ۍ'��?�@�׻Y�<&��t��P��{�H|��,?���+w(���̋?	?\(zZ��J��i88U�X�X��������s��qS�B5~�A���?%��A�-U���W}�L#�ly���P@�l2�S2Ԯ��so�r.p��V�{A���͑�c�S^!�]�����xZXF�#\�#���i	����P�?��t�����W9.[mcU�[�y|m{E��t�u!�ڌ�P2g�������)��k'F\���umB����ڍާI�/�/�_h������!��fa�j�#��1���H!"%��`d�+EWr��=Ыg}�a�Q��`�r5�[�D����&�Bڴ"��j�ZXG"u��g�޸��Պ�lゕ�H0\y��	�U�������,)�]��n�Fr�_1I%sXs5�G�q�3Rf�Q��{7�'�VK�D�d����"~ȔY	%��Ybȗ��hr���Г2�G�<^6y����Is��/%�'m�.3$�X�/Fє6����P��^������bB���֡w��A���$�ˋ9}M}c�Wݛὒ�k��:��u\�B�����R+cX>�l��q�x��b�w.�]<�!Ȗ��U�*@Y�A��;�x�&���\�� ��7~-m�҉��Z�Ƨ���,n7��-��yyI,gv�3���<ɇ������ױ3����"̴&��C�����(�&�D}�/�z����!\�3��ϳ3�
��W׈���VxZ`�$I��))��Q��!�v��+�ۡcOً]׆N볘���������Zu�F:��+�W�wɌ�Q]�"��+}�T,����7"��D;��=� �&��Ӡ$_&Eۖ+�x�#�{�<����{�S}x;�n����9Y�fm=N���7�R� ��� 7��'Y�B9$2�kk~(wE�/˷l�3X�tc:ɞ��U:q�=K�'>�q�x}Z�c��9-�!�j�����2�ףڲY��k�[�޽q�V��Pu;ﱩ�Pj�W_7�S�����}��k��_,���v�p|	"��]�?2�ϓ@�Np�5������d��ù�ۗ+@��M�ψPbbw��?,nyoz����Xۀ�Q齼����Ɩ��li59q�7;����nm��n^X��7l��@-\���v�:��՗�~��f���)�����k
���z�+jȜ���Ї�{�34w_<�F�N�xݦ���E��D���(��$IިU�q���U�r�]T��=Kw��6�:�b'�_�I+���a���<�A�֥�4`I�)��w뽌6t��8o��**����K�u��>��kj^�B�]x7��	.� ��I�Q�;5���d,F��	H�����o��>��wҷ�����b�fJa�D�`�'z1�U��}i�,�����P[�kC��H�Ԑ�L�*���Ul�!�d�\�^ �v�^�� {�j��c�$�9�1�����!R`!��K���8�%8
:�g��O�tn���2�W�KW����=|�|�z_tPV�+���e���T����|#�W'���͍DZ[RY,����]�wj ���nY����ں�t����P���_�d9vb����k��p�L�T��@�?6�v�2��Orc�əU4Z�!����*��b�[�1ӈp��1�rx�y�0U��"��I+/{�,�75!Ԙ܅S��M�����ՁTX�>�w�C~b�^���a�t���4PN�x�O�i�4�#?0w>�n��(�]�ƍ�98azv�Rm��"�]J4y3���.����3���q�̳	Q.Id��j���g\��l�Te�rɞꨗhA�XnH��Q���+B��������Tv�����,�jih� �e	��i�p�"��f�Q!�}G�����
|=��:����_{����v�T	�g�v�.\�_:"k;�ae�����=�!��ΰ�+��=�i�#a�dWL|����wH]���k���{��-Ŋ\�Z
������=��ӡ(�u� �+��J��Ĝl\���u�qz�6�87=������]�M`_N:z�=vvx66}V���g#݁��ׄ���v���7du��lu=;��ѹ1�v�	�ƣ��{z�w��p�b��m��ع����@,�殏g�[�è7��h�s�Z���wGYK��>�m;Lָ��˸�����B\m�E�׮���/|l�v��CR8���.����cF8�r1�]ڱ�^7\�mՒݬQj8b����qB�*I?q�/b��W߬T�#e1.��
,�$E������Y�� ���C�%JF`�]%��7��|J8L$��5#���ˊ�ˣ��k~���z�!䫅��b�4�(]
�Cg}�i����:%���S��Z&I�$H#��n,Ɋ�?��r��TCk����c��Z�^�g�zeT�o��9��}W�%�����*!0�tæ�i������Ht�N�s�وE�q���ަG�uʞ/���t�d�vu�~x���gmOB6�,cU�5�f.��]}󌌔��[���l�{s�'�*F�?B���2E֧��(Ơ2)���ȡ���2�%r��H#��HS�r���S�1��`'\v����byl���`#YȤU��Y2�R��%\�E޵����3�>S��M	e�1�Bf����zE�۸L�[&�.�l��.��9�KטX�QN�i8�v0�r�V��o��6�F���<�59��rą�o&ehט�'$0�n��R*^WjЄJ��OMծnP��(�����aУ�/zץ��i�Ϥg���V~F1���ëݡ��qi)�;�a��G��g�\��z�&
�dM�_�84x�_i���W���̛>��0���2/�){BqӧP�zT_q�w��7�����v/E�P@h�~���6��`a̠o�#�5;�j�Ǯ��0�54X�@�6���q�cvT��f&%f�T�5�gY]�X�x*�tzNi���!Q�S���Y׍�.x�TQ��B���K|���9�o\*��6�#�FT��4���>���Z���6jK8c��A1#C�m��0�Ӓ(�ƛ���Ms�6v�*\�ލS�@n�Yz�H��U��ޘ��Z�N���$���Ⱥ�"N�ӗ�2����|�e7�Yqc��=�|��Fީ��āMG�9�LaQqد���V�0i?����]����ʲ��6�j�.M"�7�j��ڴ~�ֺ׃�f����v{9�%*+��,�ۤ�M�g���쮚0�,[���>���=��Lc��#��o^�=V���I�����NvI+��D�b��s�ml��W[��Δ%-�Nh�T�o�Ꭿ�3&��M���Ԡ|�6��&\<s-��P��̾+u�@���. ���k�{U��Ʈ�k!����6�nJ=��d�֣��7w&�軔;z鑪����:y�5��ф�58-�0��Ͳ�x�U�В�}��2�\Z�u6��w�x�p��7RL�]��{F�jP=��E�v9�G�^���T�[�髢2V��dVD�b�kG�_)t��\tj.���^v�M�nm�o���+_rރ:������m�eH�1;$�պ{QbCm��xv>�ᥗTi�Rd���S&����1�e�X�8�-9.��̋�s;���X����N%J.�;�n1��*ќ���2BUjKe%�]阙��a�RrI<]X(�t|�G�,'�Q��Q[��˶��[�hI�B�fJFI��7Vk-�٘�'R:b�ۼ�U�*�{�hFY|�N�.�3,̷S)�uow]�V�2���ŰD�sk^�v5�<�2u�iQ=kj��Έ��X����j�Ȟ�ra:9��1���kD��0��o$��st�l�cV=�;��9��'Ělo	[�����yܫ�\岹��f�`SC���u�/�s�_w\On����q��OgKܗ;0Z�9���t3rs)M�GiNьɽ/z��y��� ����.��z��s{J�Y4+k�UP�QZ��Hs��s��++���	��^ӛ��T_]��r��q����Q�!�>0��[T���Z_o������ڗ�{��َ�ւb��c��9s������f^e���˙.�G�{zJ�F�^��83�B�ц�%�#�B�;g�6� <�z��4�}���5���>kC�|������/3�S2�3`aw�|�j��UP�M�E��\3��Ѷ�{#��w`�
F틵�϶�>�Ngt�c�M:��.�J�-^�u�B]ѩ�
�.��,��N	�R��̣f�W3�uY�^�l���DT�T�^Ҹ압W=C�xHT�@b��n<�*�Ü��d�R4���F*�I���:�/2 Q�&lӳ�wKѺ���jU�U��`�ܤ���ZQ�	���CR�UJL����4'n?���9�ìVl�L��R�V����s-T����:�GT�BFR��*F�ƛ#�,G�n$܊�m�!���8�^���e��1�jΟ,��C�����o��&0�FC��� դ)H5r��i��Z���x���[�R����=V��>�#ls��֬�n�@�ue�nvV�ͻ����(S�t�澴x.8zWچV�� \� �H��"QXE�5ކǽyR�3ʷ-�YU���c�p�o}f�wL���oO\9{��-�`����Xz��,[�o���!��i�m�]�4Fo"�v�n���s�A�Gh9��v�:��ؤ�u�䳻���k��~xv��i8��a���GZ��*�;�G��W����pfV{������y[�<�BO��p7�~.,Ï�-��Y��;ޥx�ǪC]}����͚*)v�ޱ������"t�D�#���K�k�];BN�>G.YFImzK�^ne�'�}"ou�F��v�t�񯰜@N�]L�	������l�p�{z)���%={��_uu6J�P� ,��s6���]w�H�\}-�[&�.����ڧCE뵒��a�����}�Z���p�o�o,nou:y�cOm�Jd�0�*-�M�7hu���ang�*u��-�w�V�(�o�M�j���Ҩb�S��y�;��j�{ݾ5�P;i���u�X軕
��͵@ff�d�U+�7�  �b�V��k���:s��x0ot�5mEv��|�e
[s�tX�()'�/j>�
��f��0�7Q�ι�`��n�t���vr	�A���F�;�[n��\�<����a(�W��l󮛗Gn_\�F�5�/&���n�C�Q�Ym�b��0Sj,]d3���c���0�M�������q�)����\;�݁�/so&���넣l��q��1���i��F��o�8K�n�8�{v�/�
x�ҫ'�pj��q�=�e;v�rn�n����ҵ�!����N�]�#����F�]���o�/Æ�b䵪兖���r-o��߿���� ��/�F�t�t&a�}=��o�5���؇���!#HBl}.&DCMX"%OT�~��!?��&�֑��U� ���P�7*�Ɉ�����%)��fs��F&0��4��]Oc3Fb�*VoV�t2�6��u�<:UVX��a�A�&#�H\jHr����[s��0^�G������殘Ki�ѻ�-�ɾr8�"2!t\�ѕ�n!�Z�=��	(��ZnGCvf�jlh{��ֆ��oz�P ��F^^���P��曤P��3��3Z>�I/�R��P�/{J��m{$���s�
R@�B4���p�_C���@�ʮU�����v4w��0��l��=�����G�)#Gx�KVׄ�fy29�QB�\��G��ˇ4lx[��w��m=�7�������OC�1�8��loLh��I�x}�GOR��]v��7%�XE}Kjpk~�r�����VE2@�3��WkV~��������<�H����`�L�lì]��-7���7�|��pz�hcE��q7Ƅ�b�|�v��@P�Y��K�fз!���B�Ӝ�]hQ�+����l�X���S���xu���WLUK������ �����;��_g��ޔ�\�H��7���E�T�m�orF�����d�ŭ��s�A7�9���,�ރM���ִY���^�m�#�0��;�0\i�M$7���|��Z͘�_6`�n�ֿ:�jf��}�$9�=�=yt�}�9i�������iL6�E8��N�5n!ѥ0eq��C�^꺲n�_n��;ˏ���v��2`�4�ޜxu��1Tj�ڔ��q���VFݣ׶���7F��& k�[�ٝIێ|"�ػw]=��X+p猖#��4}������=��u,�&�I�U�3U���T�_ut��RN���we\�ǜ<hɲ��m�%�$�}�s�4s��k��D�A�6!-�
�ȫ,��TF��~n�cOӞ��<����˪#�=�u#@��HQ�g�B�n��F+�}u��$�6���D���Ѫ�ۇ��
���q�f�X��x���
k�J�y���v$��89F9H�����!�k7aK6�];�~��+(��]�'��goqQg��K��Ы�2z괞��ˀ��[ɸJ2�*(�-�����ń�-��Br�Jf�"JhP�������D�u��Dqo8S����3k�����ֶoƷ PV��1ʶ�}�N�h}k�����>��ّ�Z<\� ��L����O����w�X&�j�{�:+�U�&r��}̾'^^w� ��=�ȝ���m	�r��&yLś>��X1�yK��[��DD�!]0j����CAw �}t��x��.������Tf1�&�<u������L��r5پZ,y,ݹ�K��D�n�	�\��uc~�����Ѱ�9���Yw\8xSպ7]j�)���Uw_3�!���Ms�,�:Ȝ��#�'ϣ�"K�8�_������x�ۃ.�� ���^;Y����� J�xz��*8D�=�oE�|i��slm������6RM4پ"���?��9͎kx���f�%������@J����l�m!^�����L���W���$a���/eZ����e��/���#0�q��s���G����5@�>Xz=�n:��v��6o��·)�9�����P�ʴ$Ϟ��T�!��.����.�'�Huv�5�n���aHu^�3ըX=�Z�_n/��8:�����O�a�p�}Beq��$܁&cOi'uŴ�h��%�l�����ӟl]��V�.���n��76+s��.������>���g�u}ި�Y�<��/a�-��M��a��k�ϥ#:��%὘���1�XB�EE�[R�Z�^=jxoz����|��-����@aꗕ�!y�N������MOCʥ߽����@ݰ�؉�$�$E��JH(b����A]�iHD���_��*�y��x(e���H�R}u����M����y9`�Ow�̉��p)"�yq�C���c�4B���?M�0CA�t��r�*VUF�"(=:�W��3z�DVa����H��i�����.
���
D�ɖM��$�o}Z�v�-B���n@��͹���$LToԺ?�Os����c2(rm�ͅ#Cع9�R���d.Z�����?E��ܙ�'R���۪u��;�S"�i�Щnw��8;N�]H��+�W����u9��U	�ȧZ�ݹ�iƃ���8ɼJsDc���ϴڭ�l;��ۃ8�M:�/m����;k�cm���������O[��n�#%��7]�5�SW/M�GD-�u,�sK͗�k���n�-UA(K�$Ձ%�\��ڡ�� ����;*�M�G���{q�W�`��Su�z	M��p/a��S�/�ͯg�Lv���lsب�o�E���[�tr���>8{n��u���n�:��]r���n5�<��g��7]]l�;to�H��4~�B��������K)WN�	7\{���ޡ���X�DTS.*7��;�֡DW�fB�H�8b"���
2�-�v���f7o�˭O^c�L_����������s���U#�6�:�k��'Ƿ��<�o�c\�"�22�-���]+���@�z���G&̮>-�D+�è7k;�{w�k�U�w�1�R�̔=뱶��%��C
4�5����5�т>�����\4�ilÛ��)N����?U����דm=��'G�<;j��x�:��a�[�I�cr��vO��4�q&��[����=+kA�����ĵDa��l�;\<�r�������{sl�(D�e�Tm�X۪�Ѻ�x��ݸ�	;\{vz�N)�Tf1m\r2u����N���01K$Ӯ[ �i�P�a#��Ŋ�8n���ޯ �3��y��^I�Hϱ[�[)"���$m�Cv��?d��%<����]�����k!�-J���[[�ɻ�.���uA�;�j���kz�
�g��cX%8�]a3�n
�)�4�
3����"99�$�q�&M�]���Xo[��{}�9��HO|<l�q�̌7	n[V�K��˳!���/���Ϭi>�Lhgu�$�{X=��n;
A)�ʿF�>`�~�#A�jW{)b��)�TI'7
�H�����lT�)l�[��k��u�q�rL��+;=xK���N�{�{�u�D����NK\�h��V�����űu�f	D�=�-���S���Ɨ�iѯk^;0ʇC�o���LՕ)���~>��6N��D�1BA�(���@u�݉܍���h��dx�f+m���G�����`�E������ץO�6���x�s;���u�EN������l�[�da��G�7��
�$l6�M¦
&��K���$M��nA_,��:�A���k���ߋ��Q���4�U'�泤��a�.�ς�IZ��t�*Ij�g7.��>��8J��")����=:T�Xb���B�r喟�|nZ���U�Z��)œ�l��Y�yX��]nZ�W[�׍蘅җp��57#Z�IN75	�O-=�ݩ���M���Cc4Ξ�C���|���a&���*8kL�����Z<}B��v}u��<�s���e7]�d�bH�X�^fp2�����ک�t�ɃC�k�|XN�e6��4�H�B���Y��)[�V�ή�݋��3���H6#u|Nf�\E���엛��h>0Y'�f��v�~$oo�qS%c_�$��=��uu�`�HG��'Xr;�{U�de9n��pݘ��V�Y,m;)��eG/�������CH��M��v
B񊻷. nW{���l9�=珚����e��+�|,��Y�J��6�H-�_9Μ9��O�:����Љ��ٵ#4|{�P�L�̿�63�ߺ���WI���Xo�ZM��4�d�IY�F��w�ЎjS����3�=��n \�6z_z�z�����xU+c\�	��R0���1��Ȓa�[�+���y��_g�|T��`�C��t��k��^�r��w�]������"���U�Q�Z�ո2���KpZ7��:.������L%���ˀ�#}GC��s��v����N��:a�!|Uz���
Q�]5����~�Y�n�:�p�/��[u��T���!m�)�܌?(��z����[���F��/E�zxą�����Vu�8+y��=�;c���n��h�n�Lg��%�'�Ճ���Wc��V��a�6��;eT�iU�_L���;X�׼�-�˦ʾ�g�ʚ�����e`��s)2�2XE86Q�\vȨ���W�'���z"�Y˪z`W_Q��;��Ë���&��'{GJ�{�F�^��J�5ar>d�db$�w���뒺cl���Mc7v+��@y�x���&�Η���i���t�rO�9	�B�p�'&����ۂ�td��qg�}8�����\6�@�ٯ�N���b�>�tt3��>���[�&e��7ۓ:d~��}����?�Ih�	�[��P䢋�����N�4D�G=2�gW�r�\+r̝lq
c�s�Y[����b�U ���vF���V�+`$��^\ S�I���d�&nb3� ��3���1^���άE[K����[΃��}|6q�z,�EK}A���m��˧�Y��=���F��:Krܛ�}	�T�9 ����UR8�����Wen���i<V'+�X���u���ښ�Ru��U]��KY8G��Y��v�f�����68�[ի��3^iM����[j�������_b��P+N�0J�u��h.ޏ�u�uh�6C�����Kw	��]v]s��DE�p�lP��앓Ur�r���Rj����N��n{.�]���Ըӝm^�N�Nbjx �Ýl fe݃���P���A�7D��
�3�ڌ��g;�7�A�0rr�aLإ�D��͹p���zft�)����]�0���ű)�ڶ�m��y�OK����_�˺2�mR�I����wFQYܹc��ol�m;ۗ�Q֬X�cj��$�7u:��aSESF>�ծ�S�O[��2S�ck�g�@C�"r�p*���'N:;M��VM��wo�	M�¥ѐe�tls���w՝���z�ΠE�
)'�rW�]}���A.��Z�M0�נ����Y�n`2V)��	2vʻu�r�{OGl|��훬{z������[�3Ԟz����^Y[*�:Nu[}}�oFoq�i$�0yӖ4�<q�7�;s�ǇW#;�%���t)�T�8-=�a�G^k��nV�9Z��`�[Y�k������f�o���Zq��;�[q�2,-�l-Z8�.��� �%�&�"l��V��h0u�@J��-UP8v��������:�1բ�"�epl(��!����=����.,��N{)����K�u�3�lv7dWi�pB\�y�<W�}�7�����-v�Qv�
y�ٕ����qŮ�z�G>�Y�
{&�i�����ϫX,�!onN`��voF�=Y�4).��췒;�Q�ۓ�e9�RX8v�/R�=<l��(%�9�6.׊n����wn.���x�=�g=�\�+`X���V����PoqѸ�9���V#���)b���/��љ��
U�����ٺ�F��W���]��r9A4d Aj�p���rrm�u����G9���w'f�u���^Z�����Ia\�۷]]< �n����%�ݩ��8T1�ێ���#���{86�{h8�)�u��$�Uyq�غ����<���AƎ�ݝ�9��>:��n�Kq�{:Mu����F�3^��ۨ��oR�'nѹ��Aup�Yܔ;㷭�a��Om��d�t���v֘������t�:�͡�s>�t"J��y�m�p��I�I��v����;�9�N�-�x���:a�;g�+;�t����1��=�ƠZ5�'lr��:��#7�n!���V�6���*d1�e�z����F�������wo�m;+Ѹ��9��	++�\��y�y��X�64\��D5.�q�۷� ��	�}l�4��0��[��np v�έ�W.Nۭ���ټ=�mLrn�n\{f���{޷R����Mre��^�cV��=粻q�]�ܸؕ��xպ�.<�jovTC\���=:�K�Rzvmv�����rc]��;]q�g��M�������Cl��ujz��&��������x���x���ۍ�n$�!u듲�EUݵ�d<<n�j�3�3a7U�\n�7j�{i����oD���M��.}�F��td�[u��׶Mz������'�����8�f�!��;���.���s��M�0���F�7:vr�.�q�;����iF�&Gŗ��)�QEf콜�u�����D�*:u(�5��ǌĔ��vq�1W�s�-v�'�j�	���l�	�H�y�:��Lvm����(�n�.<k;ٶ5��8��s��
d�����1Ӎ�o�ݕ�۬Wgas��P^������wl;�����gR���m����"#���'<����ܩ�Hs󸶍A�R��
�tV�g��5d���l��)f��?�T��u��?���N+ͱʳ�b2P���h]�`���g]^�\X)}q{��	��6M�Θ�\x�^�gWe�\������^�]�p��C���7}�l�.�:����wQ��m���@�����.�!�	�FI6�6tZ�szt[��D�r�LV.��(+!��>$s���������<V���~K&�(=H�r�)�ho��J��2o���M���[���qk�Wj�#M���� �O+�n��~�o����0ƬG�<�j4S��؉�3�8w�ǬVv,���xb�5I�ul�]��<;��C��y�띂��&D���j�J��W�����s�Iu�a;�M닅+v�.�u\��ݹ��F�FӔ93v�Q3q�ٔЂk^�U�7���0��7�o ����)Y�j#!�{}�^�{k��=�r	�� �-��d����(F��|��{~>צ`�PJYdA�Γ&{ixj��ht
���/�
������뎸#ڄ���kH�yr�?�]�jX����͑yy�!�L��,]� l�{;ֵ��y���4�*߰�	�:�)�P��E7UƵ�"��whו;cK�s���yW*��*��L��3N��\!����e�����;�҉a�,��b%!��m��Z�Kͪ�W�<�rt��VW.u�/M�{S�]ZpΉ׌v���lܝ�e�?C�r2j��q3�NF�
���#8�(皕.'�Xx����Ww46�X��[�/�fNi��>����oMY���9;=l�-�I���kOc����i쇴�ek�fqh�M�s�N3�qQ4���,����u��FN��u��S���J��?i�=<'W�V����T�*�����0�6�M��T�10�Ȕ'z��X����71[�&y���NM�c����EQ��\������x��R&�i?�����o�x�=�4�%iq��(Nݷ[h"ǵ���a���m5���teֳÞ��`qi�D���凨]搉�iWbK�}��lݦ����J]Қ���n��t�Ɉ)+��E��� Ի�"�Y&Ƕ}U�;�[�Y_;���,H�4�����v���ժr>���5'1;�ޙʎ�lѵ1W�ozԧ���������n�j�Wb���Z$lG`��y��&���ŋ"�tS��LL-�2�m�J��g	R�^�Y�Нu���yAB˸T�s2�׈B.b>͝��"`oD�
ձ��Q/�Z��
��sv��\�qŴm�]�z��f|��Tm�?���_�0-���TU�~��8(��U��@ǝ���V����ó���	c�W���rw]N���-�v�<�%��0�#ˏ��]*�k��M�."���;���m�?m�I�q���K���:�(!F���A���A^�f�s2�P8J,�"��-}|hc���ǔ�zߥ�R1x�gejx��jwWI��;=U��R\(�^��B��ja�3���bi�����{u�"]-�����.�9J���Mw,X�K^��t���J��H�T�ӕ�&�
G9��ۮ�.�ܽ�`�RoQ��L�8�+��rJĭ>�cs-,Xv��)����B3g�\xa��@Y*@�D' ι�'p=]�<u���a��٣�T�����C�;�%�O���-L#�[��@y��m�>���[ǕR��mVE ���U�,����7#�ޤ�v�֎�7f�u��rmp��*'3+��00�|�o��C��Z�vD�Uu������w��`�I�*�R���#C��_\I�Iϣb!��&������km����u2�f�GpVt���.�a��2�I��NݿN~�G0��b��f#'�w'ak[��$�&�po��:"Ύ���fחE��	��>x�?gAiު��4�Wr���
��W2K��K�Sq�3t�nb=�x%$�9]���}�v/S�N�uث�O��E6qex�h��}��
��aζ+�a�AN�E �lD�9A���狞��1o�:�>֎s���ھ�����}>��K)ܺ���1w_؏���t��=��
�o9�S�2tf^�T���v��5u�m�[R��b��$�NzY��ʰ�E/=�r��l�՟od��H���I+U��m��M�@xݎ4o(k:6��w:㫝�]��-�#�[q^8*W��rڹ6`�o>�	��73��:�ڭ�����	�en��=c;V��;D��*���R�_%�嵶�3�\z��{� �bu�Lgm8k�n��n�u��ø��]W N^�,���7��u˻qRkzu�f�x��A��<�;uہ�����W���۵x��]�iݴ��B����	�X�n�2�&Jj�֖[)(K�K[N(ܳ�.��p=7}�n�<6����[�T��:�{ߕ��oQp�s;��Ã�j������$�,@��"���6�����|dq�E��#/Q;eɞ+t<�v~F4��3w&3n��e����1�9<����Ý�۰Zj$���YQ;���x��5�#��8��0|*�{�OJCc�Ȋ��p;�A�'|�3Ohf��5j���D0J�%�/�݇7�x���Ҡmչ�r��GX13F��;x7��;�^[�Y�G��}��ћ��C=�՘&9$B@S���ؾ`���V�+����yc�~��	�}�^|ژi���utg�����f�T���`����Ńua����ǧ��Ѽ���N��W���W��l�-����X]�\L�����ߟ��wL17x����.�i�_0����Df���5��GU���p��Y�����~u_J���pF㱨mE|��.��B�My$���ի�g�k�m��V�yN�������|z��Z&l�����0�j��'In�4`y���a��7�2�Uj��#L��Yb��!��\V�F�/8=�riEj�E���M�P[���A�|��k�١"��\:>���_���@�2�T����x�w* h��MA!P�arG�N���qGX��?��ݙS&����7�+⦍�t�|�\�c/��?}��+�B��&r�Ƙ�)wV�QJ��#	e��d̄D�Uo*7�땰$Ms5�5���'�`�s��0)W�F5T��<�ps��i$���V�M)	%"<��ٞ�vzGyC;��#�6�u��<�W��X^ ��UQ�6�]� ���-����)�\)�V���j�yE���e�s<�#������#D���MEI�,oNN��q]��S%����u���5VJ�9[-6�,�����a��A2�#9��c�!�BJ���rne:��ܤ^�$�k+C[&��Ϭ(½�K�%*7��tEdC�8��2�1-t"�(w\��;�0|�Ǚ�ɾ���z{v)�LFM���Z�X��������kAꝯ,�� �1�.�W*%��B�s�1s3����w�{��)�z;��gg�fT���:h=���t9�{޾�E�:"���,�#G	IǸ=kԼ�{)��m(C�+�/nɶʔ�9l�<'�"j|��화8}/G_A�B�'�Ӫ?A�u-Yy~�F��AŶ�mq��ms�u��q�4W[�\
�嬕n7[T�q���/Y�=�y��ı��)���y��R��M�I��ϑ��1�]W���_>R����S�}/� (R��I�C�����p�g��J/_���D2+u�&�幏�&��rƫ>��r���5M��>{~�
@��p�q��q!gN��^V��Cx�)�=�QL�#a�<�&���>�V+"]��Yy��%x�a�h���8��*�P��ι�H��1v<�X<k�wGo���]{�76�����:n��V=�8CI-��v�4��:_�R�D�]G(�r�Yn�Dq�fP;Ǵtυb��qX������#�"�i&�4��T��W��x���Q�[D7!���[��aşM���Y�g#/T��]{S�핒��μ����@�\ǽ6�9�E�������"����٫f�Q�yٶ_�M����qaI[�5JDTI]�����;��zt�ϝM���I�M�4N�{�*o�=�;b޼����3k#�]>@��J0�i6c�,^(@�q�j%Gثh�rm���A0D+��m�֜�O_N�X�Τ�AN�Ϩ��1�#�i�XH�E���G��g��uTe��Yc&.���*�7�y�P�S0����1�z����{4��7VF~G��-�18��aCM;�q���1��{�w�=�ee��{"�����z}N��[���ϱi��s"#�X�� ���1�r6�ތ�;�)j�ݶ�˚5���^j�z�y_{�w9�^G`��YJ+��wWJi���*q�O�9���X�:m,��ݢ���
�w%�Ab�[�,�4��l���챹�q�z�.�O=X�g��,�A���i"j���"����>mn�.�^6.N�uv�t�v�X�/b��Gu�g�8�z�;kr��{[-��r=�����z��}��˻�۶�v�[vW���s�2��n�cr�N�t4���Q����46ms�á��;n"M֠�{/M��qp�]��;\�z�뵳�k�l��[�%s��nuk�M����]�L\m�v^�c.}�76��]v9�q]�����n����m̃֍F7<�n�z�ԏ�.����β�gg��r3�D����?����c���1ܛ��5t[���~��l)�͐bf�R���f����;�]d�*������q.���z���Ŧ{2�郳A�������ޅ�j���u��w��q�l��O!Gd��&�)�Ei��{k
��'�yMu�)�=�4��y׍������ظ{n���(tՎ˾{�H!�x�n#!%F�F@ۋ6�Vr��k0x���'�z����=]t�ƪvD:o*N����R�a�Q��f�͗;̛|���Im ��2���v�j��$l�G��������n�e���p���̮�=�{��}܆:�����s݋��l�F���<�*+V����<�.���ô�ù���rN�8��S���h��=P)�yj(�>��6�b�ٰ망�ٚ�����z)Fi���o�=#F�X��P��RX)����7�+�ش39�O���.e׉n��m�3��´���RLi��8��cx�C�����d����u�R�8���[}�;����ژ�y�4|�ucv���{�܏�*�r�w��ڳ5�[=��7��V�V����}]�F�a����k9�ܶ\�W�&n�>j����k6��#��Kg0��=�;鵺=�X�ݘ�ܢ���sh��Q�%�Vߞ���۴����r&�7}q��=�t�c������B�d�ti�{�S�k�j���T~�u��f�"�m���|y�ұ�0�A�R�����3�"?�	����{L��p?K~�r��ԽOp�+����|c�O��w*h��%|nL���/=��c�G�pq���\ե㌌�fN�g�87.�R�m�_��������C�GNE��@�hglh�7����KoZ�Cf;��i(���	��[�iM]W:>�~隓�(Wl�^��N~ȗex��w���c.���*��:n���w���T}�ZE$�"\&�p�JW{z�/�>]m��V�o}U�����K/g��Ů�S��vFz=�;;oo{y.�WM�}4JF��۲ǜ6k�%y�}1[̤3Me���T�#8�oX �ee!�Ȉ��Mk�ثa�JNF=��i��7��eLLN;���'�|�����0��W�:�5{F�@�8ݽr!��p�%Wc�|��^Z�q.��Q<�r�RU��Gf�G�hd�"��d�3��g%]�ɬ�n��������i�����PKF�����u;5�Y�=�t�%},��Z�fT��n����$�������v*�_����\�T��;�{q6�86�j��hK!��-�� �vnu�3];V"����:�'L�
StV�|٘���� ǜ{Y��X̍j�@�x%���ݲ���i�L��
\��5�[�إK�]��֪������3Fe�UV�Kѱ�)�y��V���aݽ��C��9�����-��ر'��������M{��wI��J�n�ʹ{�U�
l��n�q��'�2Mಀ�$�x��΍Y���.�9���*i�&:U�\{(ͻ�uZ+K������߶�	��;���X.��Z~M�WÕ9כxL��T�P����=��O`��sinlRt�ǾS�;5U�R�沇ɣݐF��Ֆ*떨7����M��9��k��Z��#�A꒘�4XW�&���]�_9U�j��1uP3p�w�)P���n����]r�vT�?*�<Pi����Y*�m�������S���G�i`����!y{�t�]	�*J��q�/�����R��|�3w#��`먷E��4k�]��dwF$�&aI��ɘ��K��y׶t�{՘4�`����%�(��w����
_GX���ɫ6O�ڦ���j6i����V$⎝ۋ������vŜGn��3q�2L/1�s=Qb�W�BcrEW��h}3*^N/��B�{�kֶ��tB���{y1K��/�sd]�]��C{1��;�C6��|r���M�Hmşm�;T­���,�n�g.��25�v�̭�,����r[��fV�xt���M�ޓ�P�sSU�Av-�q�ƀ�Q��-[��fvI���z*�Y�o&�?%k��s�`��Yա�uܬa�CԱ>$����"���I�*��;����X�S���Z��x��zY��N~g�S�c������tUitȉ�X������ ���y��wҖJ�6i]L�,�{N�s�49�Y���x��������%E��X1,�E��O61	��ք���6W����6�{��Q��[��}U,�/f��t�~���|���(SݗG\���k�^�a�ui�n�	 ��l�����tk�]A���,c�P�t�a��ZGmU@�PVe]$������9υ�ʅٝw:�9�ƞ>�C����d"��9L�U
�~Y%�.}�UϏ�QI�!hIIɽ��g����0.�~�w%�D��Y��[�r�Gi��]<���Kz�ϫ�Éݻ]��~.��G�,E!(��i4��&�s�m�k��]��;_���y5�#Ջ�z+�Qv�wg�m�Xy�U�v˂h50&���m��eR�:�ķ{z;q���]��3���|s��ͻ�/�{ 6�=��{�3�n^u�"b��Q�$�14J&)"ͭ�7��|� U�6-��=�j����չ�u��"���6�;����F�+����ִ�QS��Z�H����Q�Βi�N�K������Gjr���r>D�)w���0���]Y����늪��IF��q��k��#�X$)U�,�l�A�l��K�t�1V+���R�-V��\suݶ�p�<V�1)��k��I<��m�lt��-�wQ.�x�>��������[��o7f��e;q��k��:�qx�yC%�uY�ܞk X���73k�87� ����V���70k�ۃ����eu����e�]��s�ۄ.�6�hU��Z]��vC��\��\-7&$�jˈ��V���&y��:����kr7~�\�y�����fz������=]�jm�Vb��?&g��}q���ǭ���v������ A�i�����#�]2I�S�"��	��9��;���&&gs�.gg�Zz���L��l(��*�u��+Uݳ��k�(j'�s�k��.+��)��Q�~D=��O�%����54�2uu��ѧD?�-����	�C�ϛ4w+E��ec�Ӯ��24���]`�3bs��Z����㣇?i�YW��'��iTF8���&������D4��3�J�-�N�o)+c�u60:���Rb�b�io[�ܝ��\�DuR�ESN�&[dw+���`��с��ӫ..�n<'^�uU��dh왍Ĝ���_}2�۪�{�6�����c6Zu��Ӛ����:m��=�u�1������EBҒ���k�{ԣ��[/}��n{lv��a2�~i�:,�7v��k�ې�����w�3n�`�.���|�O{��1d[���Ad�z�.̺�:ͮ��<�G�R�T��i�����䷳�ӻ=���"��v^�ڞYG�Qx�K�*"ZO��d�3.�G���=W;X���z2Z��!W	���}.��Q��_d� =}��3xֻ�&+dGI9G㙔�ʂt��I�wy[�nv�m_Y�u|�ʊ,;ǲ߆ͯK㣥M�z��[����/ײ��Y=K~�))�T�]�����j�S�:��W�_LG�:�q�ѿhz�^��}����s\{����4�=�GJ��F�*� i��Y��W��vǗv���V�9,�v'[��9N�޹+�K�43�T��e�L�3��ck��7�%�����OX�35����>��0c?@��6�g��S�=VqS�l����+�L���8�į�^Θ�2ƚ�S����Y�u.�v�#���pc&�QD�2@Rq����������lEK��\�9"�t=�&C.�=�A&N��E8�޳��YV��u�ġZ\wA���LYEl�;Gn3H=��.J��1�u�ָ����N��wO<<Ǚ�uX7c.��@������`�F��c�0Vq�|T��o��]k2��5L�nw��h%��Gr��T!�mw
㴶�3^g���`Q�/3��S�z+l-�n�Q=�߷�ij���0�o=��5V[Q��V��؎28�W���V��lB�pw/)#ۭWkv�)�:���7����<6����Nl�E�\�b�*?���%զz_J���i_�S�^M�BWr˙=�n:�$c�q�s���E�iY��^F��)H�p_�։�.�7�uI�V��s���=*���,��cdb�3�/4��p�Ԑ�����O�V{I�a7$��N
�5��\W��c�m���=����*{Oǻ�QD�㮯�<V�;�1oҪ�����1��B,��	Ho�V���'��'�r��v�l�)������ "��̭�t�UG7�9�E	q��{|^	���������9�5��t�磷݂��役�쳊�"�ݩ���K+�IҌe��7����*���J��3�FB��e�x)V�kx<=Ҟ�}��;@��y/"�:ʑ�y����sn�U�N��>N;�ZW�����R[1�7#,�+�G�a)jV��x��r�Y�����7e�m��}|�q:�-S�=�k:��4믘��j0����IMA+�L0�D��j����B�B����$QER%Mȫ���Q�o�
��e�%k9��Nl��j��TR�I�雘��zV�>��������H5�$��k�Su�%�#���6��6���L���,7��q�k�l�4W]q����aR�Ӭ�h�ħI��M54���1/�>��Km�H�MU�Q,ͭ=���w1k�/T���{�W����[">���.�
�%�Rleb�5��a�����x=Sht6}(�Uo��h�z�CqF�W��??�fp�7�>��v�|9���%Q��B�7��z�v2��xr��ʖ&�1�7/^"�'tY�%��҉U,�/FV,��^���?g�;;u[u��V��녱��;k�ݧw\4B�hd0B
� ����	-����x�sՉ�f���ţv.k7c��'mѫ��kW�ݼl�5�;��,(�r�/M��`y8;�,N\�+q�P���1�ν����s��GY,�X魇�Rlu���"��ʀ�h+	�c���c�/�ێ�m��RhN�R�4���������hb ��h�����χmY��4�]mm��2����FF; k�爸:��jH�	ġ2S�� ��:༧��x�G|��҅�IZ��u�;&��;<�bVT���E�]L{Bq��ae�a��[Զ��Wk��n��&�W�[�U���B;(��s�Z&6jƛO�����*��F��=���w����#"D�1����ۭ�uý!�,��^�C�w�-.�v	��Eڗ{*3�q%��vX�����Y���hv
j�l#$�&赹DMՊ�a���3;����c����^�TGv{d�� wW��Y6Z;C�|���?	�D�p��q��خiT+�o����)�Pqq�����ghP��]wF�۵Y����_6�n�����+s�O/���p�"*F�.'m��9�,��0�V�q����%*۫�EԸy-��8�1��F�Q�3յ�jw:��W��D���13^[<7܁����ݻm��#�^���#��q�6�B2�E�塙Lz�wM�7�࿕��E��1���Z�2�&!����1�٦������A�������᮷�k��,o�1�L��H ���[�G�u�`"�u+�iʷ�<�=���N���^�}��%��A�M���Vs�^S��i��R=�w�#`4��}2��ln��Ҋ���R�uD�	��wn|r�ʦ�4�b�I����EA�X������{2
�������&��^&�b����p�%K�bz���6����=)F�Q(��K]x�<�k���/�vl�9��v_�T�J^Ň�ʍ3N+\�������چ���N�����8�-�+ς�zx�ظn�uk��q�<�4���o��[���{E됼�g ���w���S�R��:�^M�{�´;�kl�~\{=[���Z���� ���M'
�<"W��CϽ�k�N��&��w����vA溁�Q�B���j��)TUF��Y<{CH�2A��Li	����U|z��{��K���^��\���!"��5��k�,�ѝ���B7;���]��,� }F���v���|��q*�KP일 �U/y{�=�����4�������m����;������ ��̻�̞{Ͻ��N��a&�9[2&�A�c���?]���U���ƴ��8�s������'�o�����I���>��!�4�yR�;͹�d��,���L*��PɫkT���)=Nz���nS�̢��¬u�t�I��LWѰ�	�	�P�ݞ$z}V��k���gSԯgj��f}��q�0H-ǫ�&��+B]����D��<;Uz^vƹ�mV؍��2#�/��ni�tS`����*m��ig'�,j��uU�cs{�t^ޫ�B��ٴ=���n<���W7㗷����IoK��q9�e����J9<�~�V+p��u:��j/��詳:N��:�;�r�:{s���gz�t�'I�L.&�Rɜ�ڶv/[�{z��]3ͅ����5sh�����a����;3��"+g>�
�2�$��5����i��:��}��M�d�;l�'����}-D9k��T�;ݣ�R�<���k�yWЉܾ�ҽ��qy��?�# .(�E�7�J��=)�ba�-�H�I!��)|{���{-<�=�x����r9�/+�8wS�b�Fl�\L"�)��n�gv�[���A�Ύ�vK�Δgdx�p�S<a&Mt[�.{S�Ķ;6�4?;����M��\g��l���"�{R�.oö������U=B���^~�V��y+"�ea��Li�����Qɵ�
�޾�w*1}�ˡ�w�`�-	�m��G�o�\!-��;���X;�b�)M}���_���	
���/��fPu*jM\����Wh���s<��vE~��[\���P��k۶���`.fHڑ�!���ֆs9Bp�j>�z��篦տy��E��h��/P��e��k��s:MvW���Yc3(���y����=�ܝ��b��g�U�o�ЅD</����ީ|rɉ�պ7��jd�A��ଲHé��=J�F3L��6�|w,�����8�	.��݈Q:��m�f�%Ӛ��B��ر�q�;�e�����kOۙ��+];+���:�t[|Q�&	�6]��[�!�X�)���b�z�@�mlۦ�fun`D��\�i�ڻW!�gqӂ���S���om�
����%'p�z�syPT��K�tz�M�Q�8]�QGv ��RsiE�_ss��T6)��U
*��,Z�
��G�[�Yݕ;Gڱ���YuЬ����N��iu���ۉ�3��i7L�����T톋�t��a��m�ix�0��Cd����S�i�6 fp�h��͂���Ay 
�f�y��~����Ȱ��T=[7�mhr,˖���0Xh1�4r�}ڹ���ھ�������uЛ�;ZC�5�9o{��p��P�* Vr���;;+���4��z�1qK�%��^�tB=��+on&�:���C����SS�&֛˾f�F��X����mF\�A�Ȩ��22�Y��C7-��wq���N������{��X��No"c7w���3����6�"����9�g�.��X��FeN�R�v�L�J�nt�@����5�7OFoΉ��&�L��s�YfF[0��\�x�U�\�r]O�Sجx��X����6�0�.K�f���*�r�C4h�{�uGH�D��g.��>N�9�;��C��l�Y,�e�ƜƘ��Ku�7��P�iY��c��4h�8�WrTR��+l�M��
gGRs����4qmg��]^ݸ�Uv�u�g��q�5��g�2>W��j�»n����[���m�n�F�) ���������2�٥�v���L�<C���M
(T�.r�m�8�N��R�Q�f��wV����kl�w�V�c�;�x���eu�������vzi盕�u�g6�8睱�7��-�x���s;�+x��]�����eո�]�ڣ��cy����u��m�7On����,I���5�d����qj9�����ɍ��ƺ���+�=v�<�ƮRMx�Ę����Z�1�tw'���)����2u��^(y�ΐ7<��x5C�C=��n6�mʩ���� ۣ��b�u8wb2'�,��ܗq�Jv;se.-N��u��d�F#X+���zܘwl�s�n!�U؎��7L��⎬�����r���bm��3Uڶ{=kz�����!��Xۗ�\/mc����o\!��F�j�����s��Dc�n���s��XDM�����q����淴��4[Ar�j�s^ ̆�Xv@�Լ`��s8!-v��u�̙�{On�wb���mnMn���Q]����p���u�#�h�h����%�i���:#�昜�p��L��������m��U���w`{^9L�b1D�����爻q�{;���x��T�A��秵����o5��=qq���r���
���Yec<��{5pg�TexKp=�m:�t���Z􋶺��m��M��&�5�6��ڠ�ۛy�<�B�j��t�w
�{\����z��r��;f���p��&�tx.���̜�s9D��X�����uֺ0��m�e�
=��͒|t_=�i�˸6t���v��@��Bb^w$b�:uɄ9��3X���)����Z\*����(�E����ZUn�pӭ���Vn��1�f�g8Nu۩7�5S�L�zN���kV6����{6ſ�����u��Y^M���]Xi�:��`go���Wt��;C�z݊��[n�h�F=��-�wq�0�݁^����m+����)�3��$�[�M����dBt�n����޺�{�u���1Q&4Ѻ����WRٖ�Q�Z�o��l��t�bm����.��5�M��/^"�O]�aە[��*�v�k�۴m��r�I���:��n����ȝ�
�|�i���`�ź�Ժ{\�ڊx�x�����e�<�m��c��~���?��]�B�qʉݎ�������6v�|F�U{fW-r�cC<�q���H�͡����8�-vU���9�Ú��[��p�{o��g�-�gWz�s�z��������q�?�_M'J'&���]�w���{;-Y�㩉!�T�=�=�䭴k�twn�̓U��P�^	H�p��R6�Yuz�!�zl�B�zg�b��/x��l[���<)4���w�®��\�׃�����Oɶ�R���q,wU���P�J�{�����n�v��-��e��E���]��.�ߝ�W�M6;�RI>q��@���.����qM�y�vu�Ok�\GS�:���܏��ofu�&�-]�|^�^U����[6�x��)(wB텳W'�Bondh��x��@�A!7(�1��؞�ն�'�ÛLh��i�כ�U����Ǆ�M���h�wF.�k8X;v���)�zD���[Z��6K���Q����tk��t�r�~��$nj��Ɨw_�Y�'2>T�w��}�/S��C1U7]g��AūqK{�+��&��p���t-)�!�\��{ P����Uh���GsAS�4���Y�,������uF����wnz��טz?f%��i��}2V�M�4����;��ּ}�d�S8�p����M#�aM.��ۧU��N�Y�kC9maJ<>���<�ۤ܅��q�7g7��5�g�lo�؁�������2HWy�[���[y���]`��=�:(w���N�dz6,�08�i8lP��������)��9]��z�Z�?Y�}�"ظ�6�K�E�tIƚH�D2E�hٮǛ���۵�Y��-}x2�ZQŷ�,^7�&�m���ܟ�^��eL��[�$0j�-��L��������mg���.��uF��9���_k��>"��E'��7�6)P�T$�h�+=���[C9��w"���Į,�GUu(%e_-z�lֆ3~�]���r^y�vI�P�,Ϛ�2e"ۏy7ד~n^�y�\1�3/ؼg9����kݹ�U��"Ʃ띓A=:��Ƴ�4`�7!�"�V?�Y��z���] ������Ԧ>�w��(&j@�_�L�k9o�ՉTS��Z	,����;5�VN�ƞջ1ت��gr�U�L{
��=���RaH�qG$�%�՞�Ի�WM��!���05r�]���Eeۅ��sS˯��m*ճZE����E��B�p����o{��e��u\��S���j3o�5�@���ͷ�=�;:�����y{�H.��%�!,�d$8�R�+�Y��YƝ��44)��]�m�`�[u�Ʋ���%�wS�o�\
�QǛ$��TH���R�v�V�?5a�����-y������מt�U��t�:.ԑ�l2Mn�fl�Y��ՖB��_�n*F%�ݺwXy���C�����V'���d��݈���ӎ��r-�H�Z��=�i�����88$26��IN,�imm���-gh�:�Ϫn_tC���a�tٖ�W�/������p��|�����!'ե�b�����8Mws)أq�����[����3��L��qE��nf�;�h�~ҥ4�ie�§R�`��y{;��D^8�����_�u�q��Ӷu�7�������k.���3��Z��<;8�M���m�뢶�Sx7�����mN�9��%Z
"��0�$H��yt\����Y0�O�<ӧM"+�o�����Qg���U��9Sz����RZ�XqƊp���^{�6�PΩ]׳]L��p��.`��<�n��4|#�Yp��}�Wv��R�UR�#~���jFDF���uve�b]]r"�-us׎xwn`�븱b����d�o�� ����vV+盗��X�.PƷq[�{���@2�k�n}a��|�'c�G3�N�5�*��+�}z��_Ro���G>$�;������o��~?5�x�Sah�u��d�eNy��U��`9٩y��p����f�g��v��ܶ���P��,���#aNWںq�u���63Σ��LC�p��^M�~��І]sm�j�E�ێ��۩x�V%�n���F:�K��nܨk ջ{9�v{=q�W����^7M��ۂG;�t!�;�nӷK�G\��u�;V&�}[N���d�.8y��_�qx�-�h�uՔ񨸸�V����m��f�Y�z���YG��TY(B�W�֩��l��PxG.�5�׵�p�17tTsF/;����6��b�q0K�f��{�f-鎢��@ =Xr����!U�秷λ�H��q�\�я%g�\�b��kH(�l������g[�Y�^7mN�Q兛/h�6�xy�S̡Ub��Z+RxA��z�����Q�؍řd�z�N;DeK�q�S�'�r�9��\9�p���&���X������P�t�	�bB$i"ۏ�$������᪟p��B9ճ������>��O{v�5N�cW�R�7��VW��a��&|R@�8�m�v]��&�G]&���A#��K.JZ)c$�#�T%_GV�@����9`�ݑêf��&;.��y�Zn��L{����4��(��ͳT�!F
iH{NR^8�~�w�:�x2��۱�vL�g^��^��j�QtA�0Y]
2�F�ww^����c�d�՘���K�y�ewY����ql&��W:��]�����a�ܜ�|�r35��k��C=l�i�� �.8�싙��[�:�v�v:ս��a�+�FO[۵n9&��i�mfs��� �6��aUP��Hm��$Zh\K�+�{��U}bd�^A�����fOo�����(l~s=r�C�g<��{�p!����E�)�s�P���~;��$������b��w^��F�$����Gt�}pe	~�����KK���'>H��_-�x�I�5�[\Ǳ��ݞ:́�6B�n5�=e��+�,��EȤp�~�<��ً5����ugT�����O\�F��wD�$���U���\�]��y�Ґ4�jC$s/�"����$��==�,>}����6;E��ˠQ�]Kj��b%֨�[c^�X�0��{=��߅&	i��3�rL�:]�WX�7�]z�q�ڠ�n{p�[-�\�_���$��2�T��,�}�VoAw�wm[R<4z�a�:OU��!�W��gZ�v��.���w��.�M�KT��>�A&X��&�$6غ��O�&�D���I_K�/q�����{�d7�N���˼d�U>ɮ
*�&d:�ך��F��HF�NTp���
>�yW�eZqn���OFnd��6>ᯨk�W08���h�=���'������p0(Z0�P�ťΗ��qRw���sy��;��R|˫g�e��FDĊ2 ���q�ޘ槞r������i�����q~;���u��J��iKfYQq�O��$x3@��.&��g�f���t�vcޗ�oU�wXՇ���%��i��ܫt�v��� L#OF�e�}�ެ�|�	A�m�N�T���s'y����N���%�.v��[��xk��{�wR�3e�C��ųI�o���a��]���Gez���ױ���y`�ly-_�ʹ����S<���M2�[�(r����;�8�h��Vc�o��/}c���\$�|�=������މ�0�Ɣ�:�\x3�0��*K��RKz�O�12сE8�5�����z+1Ka���P)�`�AZ��=s�}����o�_�.��m��|[�4{8ힶ�U5c���U�B�9��bOIM�ܚ��d�;����n�v������M�b&�I��#�0�ݣp<��r�U��z1Kj���{��V�+��w=��0z�~��%XxW�4#I�c?!��d����c%�lY�K��[��%�tIU;�З�Z{�n��*�P�����\E�= i�I�Z��M	��;�jMB�<�\њ���<��� Q���;���c2�%�*	��!�|b	��h�.XO���y?x̼��}�R<|�M87��^ދxp����f��w��g����$2�jBm�����~w�3�y����g_xޫ��W�d���T^���Y��{���� OإZ���
���bň\�Y�=��;�{��^��p�T|2��55뙇l���P����]s�J>κ^.l�޸R�l$n���+�pW��s�>���r���͸���nܱ�Ad�L6�mm6=��5�f��g� a]������ͷi�W��i�Z�w/���C[�
nq�����*�:U�����q��;s��<:Λ��V�Bǂ��㶜��]/X{�m�a�o5(�:=��G]s���>`dDY�-�{q����l�j��mW����ZͶA��W���?�f�6W}V�����fs讳��3�:5���չi$���BE�)z�����/?�w��˼V�fns6��i4J-*��q���M��t)���r)#Μ��,���8&�tK11��-Sףi^-��2�m��X�=0�������Q��V��W�1E�I$yW�h��z&�KVmdc��uʾ���o�}ӓ�2�v(���ʥ�uA�ŌmZ�>b4�ͼ5�rTV��X���z���9��Р�w=��՝r�K3U{BĽ�o�E	`��H����c�G[<��q`ج��D��Y/�9s�Hc��YV0����U�Y���]>o�[RA�̨RKJ��N����Ń6�.M�rD@n0�z@�L�i��r����7���y3���$��z/WW���qjC;��w�B���^'���Ήz�p��V_����!F8F��3��;'��f���{u��Өӿk�P>��foY���-5���m����Y2Fr�Y!u�{5IC�6u���V]�N#+��^�7���	�yLp�?t6��|.�b{:�T��9�	���N�K�0����޽,��ɒ��J9�>A{0��蔓S��|�C����n�M�������o�_��Al��3~��Ӭv�n��ɭzL�JB���B�ch �klb��ݶpo��5���˫z�m�L`�ÿq�<˳�;�7Fv^i�.@����jGR��F�洹ɾ�]�f{3����Mf�ڊ��{��tuHMn���DU�B,���s#;��|��|���FH0��.����:�Ju&�<�ک��e�cp-�g3Q���D��q��;�hv�9��ѯ���1��Z�maZtԏ��1�.��w���n���",cx�p���`1�BFI˼��g�ʘ��mE�|�O�R�N��}}�.+Ͱo�N�i��7w�w����%1�z4u[y[�19q��܆��3._e�1j!s˽]!�8���,�Lk�k��з)J�:mK����K�H��uv��E�ɾ.��a
a�̝kɵ�u��F����cP�t��IW;����Ρ���:�N��� �U��yE�z=��Ґ{B�+�p*�8E�uF��H
�]�7'
X�h}{�Fn�G�����6r�V�u���M.�b�3�t���8��jܵ�T�d�,vT˳�ҽ����xټ�����]1��xܾ�*���[�V�\0��x��os*���m���Е���$�l+��bݪ�7��(��%n8qB�-�Gmto���:LR�`D#z���nn��(o(��.�����"�֎꥛��R�e�f�mY<ܾv�Wa�y��|n����̺5��UBa]�m��g�֕�-�]�3�R.���r�s&�j�U�k���epέ��<�M�}˅7�.�j�;Xku������ޢ�"�!�{��		pf�ZM��\g(9K1s���qU�QcݘKW�^DE��I[�c���йi���Li�F	Z3����.���;25�i�z��n+�y]����<�tm(�p��Ėn=�tM�3��|�m:}s]��o���A�z鬕B4����֗�'F���'�r�0F��\�(�ݩ��:QT������D�0��I�J�&���`F�m�s�����l崎v,eT�s}�K]b�N.-������d�h�+H��<\�n��l�wX�#�no
y�a�ܣ|�g��dJ��+��N!/�{�n���a{����]H(wb�!rH�.�N
���s���.�c�8x����˕��.B�����c��ߡ������z��V�a\A��D��0���r�����Ժ��.s�Hb'ʢ�B����ݛ�:�.r��Ѫ������[�4�4�"�R4�(%��vz�b��ɻs-az�F��/Ӱ�V#BrsDe MjA��z�a�����o'��!'���'��v��e�B\X]6�v�L�r��x����N���@���}q�z��Nx�@���x䈊��vq��=��bӻ�X;�$�q�����	�����8�hĆ9���GDοO<x
��#�����m��+�Fvy�#���ζz�U^�4vSu]��4:Ne)"fG$Wh��c��Yyq�=�׶6z$f۸��d��5.��n��β�L5ٔM�c-<cՋ���u��R��J��nN��W�)�ENIf�˛)�I:�|-bk��Teeu��:��Ę�T�J������
���C�����,�W����عo5��e�+s�=3B�9�7�|�l�h�|�v���/Q�o�cL��#i��1��ڙ����A�����8�vah���Js�9�}[i/l��$4���0�K|�3&P���oX9W��f��Q2�*�/�XO��V���caVx�iZM1"8�q×,�>��^���i�y��Es�)�����_���EK����x͌F%]/���y�y��DT&Hܚ������9�hk>}���R��
�Hē8�S2OG�V:R\����
�uM&1p9�8�&���mrv���
�k�딗�C��~��R��,�WXY.��:T���j�1I���b�^esƦ(}��r�ťo�퍹s�Kg���J?b�-��w���]�|�Z��ivi�[�G~�/�%�S\�g3���莹��T��;��M�neTU��C[%�D�)D^�֣����y�ׯ��{�R��Q��a�H��d�/m��2�\�f&:l.v:8��]Ԛ��Z&�<��M�����r`{n���nu�ʜ�M8��TJ��	u�Y��3�.�ە�
�q&G��n�
I�hpWz��юнI���$v㋆:�,��j�v�],���v��p�б[��p�:��퇓�;���m�裓Q��c[���v��;�Ꞻ6g�=sQ��;S�1Վ,���}����=��U:U�'c��1ˢ��\spu�oXu�/S�w]WT4ۂ�����8|��>��I�Ȩ�9<noº`ѯЕ����;�x����s�=�2��ʱ�P)�e�Ip�#�ە�����Z�P�a�s�h��1�o�}��c/E*�zn����\�����fNC��i��-Rc%,�$����9�`����#2���PF)�2+9���������VKu�G�'3 �ndB��9V�w��\&�[��>;�{=tLd��/Y���������ƫ��}x^w4��͛q%p5I�J������z6�\t�����NAC�1�c�J�v���T���z�c��g�[�Պ(�)�����J�ֶM��A���t����Z��H�4��z:�;r��Q�Dq��O	��b�������ڷ]^���/����Ғ"�O��|�޼5x�P\ۀ��-CQ�yX���里�PC�
�nN��U՘
�Ë��oge�G/X8�Q�h'hnU��/
EM�9$�ؿ�l�\a6(� ̩�+�$�uP�A_k����7ϕ�.�2�z��ɵ��c�q����^~��*��FHb�����v��LnGlj��r��D��ds��݋g`�t�0�	�:p��A���"NI�����P��6��˹U�,�UܕؙܹO�������P����>[���-r
H�_'1�#�V�>�<�"T�M���V��痂��ۂ�uתtΘ������%���'��x@��~9!�-�뢜c��2s:h�v䱏=�\9��^9^�a�o77f7bY�o<��J�U}��6��ݞx&��\B�x��V�;ፂ�O��W��\��Ι�
��4D@�$��Y���q�t�J�����{�8�Q��ӛ��X�]�qU��cw*�/s�KRHT�:�돨�B�"p�w�Ne�,�Ⱥ�}��������k�ϭG�e�y�r��yMh���w.t]�u�oZ�����;ge0��Q}���4m'X��B�V��q���
G�*-��}[�ztn�=hy����ӆIai����o�K2�ٱ����#��ّc[%~��y��<9��h��z������BT��Ĝ���$�WbẼ3�}�G>��ڷ��sg���T��k���WK�7�C�ݬ�1D�	\n:pt�G]��g�M�pd�1qj�p�q1�lvy�緡��<k��Y��#o����{�^Wj���mָg{��n(izW�v��>k�=����ul�Dd���u���)�q�̒e�kzNY����:���[���v�d�^c��<�6)%+�/��2<�ު�2�����6�2�h�����;k;�<h�G���כ�������)���]��/<}�|�:Юqв#�C ���uy~���&�H*�3�o�U�� t��:���z�c[�~�5��ת�+�x1�����&�H��{p�p+�T��Z�;�U.p�Uu�{5��NBz�g,SaŜ�
�e_���+��fSxRw3��28���p{�'޳�v�ηS/�o-no��guu�G��/w��Y侎�q�'a)��F�v9�OLc�;�oBC���[;�u�0�;u��wJ��o8�ܼZ������r�\]UfN�3uv��vHk��.�I����:s����
׼j������=�eZv��{�����R�ұ�\�tED�L��qf��5�82�D�Z�RFmf:),z���x�Ž/�c9\�����tJ��/s:ܠ����8�D�"fn�|'��mۙ�W�x�z{�mM���;gl��4�����r��4^��D�RL�0�g���8�O���X`��a��1���W9��ou`�ڣ���V��|c4v��:�J>�")rD����|��c�0�.�Y��.�1u)������*~
���1<�3^pc����]�Vh��綕�j�b���{$�λ�
�=����I6����-gD4Dvվ��y�r�*�jaU}i����:��x�+�ؠ�L3iԢ/�[t�i���@��
���^��@#+)a����G"��=[ѻP�X�XМ�Nc����Ӱ���;��;c�vۃ�⛊}��[�	�:��8�{ �]�����8:���L)��(mtR�S7]��4��ts�6�v�kd��<�OO ���^]Ð(%���aM��wq��S�բ�A�����yӓf:3�:�tݷ'i�	.6f�k�z7a�ݛ���;f: �F����c]6��)4��A��ʼc�*?���Z��u1������,A��'�t�Ҷ�����m9������)�u[���n9[郓I�M�& ���7jh��N����:~��]�±���Y�s�������f�ӽJ�5(�{�^���f�O�!96,NU��2Y�ګ��Le�05�2;���֩c����2�gVV�����T������`x^��v=����ZŽ=�;��=�kEM�+ٴ^��*Z~���x�%���O�6��$�Q�=�#'A����ԊǯΖGW��Ǎ�ܻ�Ub�ӎ߭Ӕ{�����N�C�<ׯ�kK{����c,
(��M�*��]��	;���U�y�:�Fx�sH���CH���TZc���2��L7�`S��0��׷zN=�|�;��K.�ǲU�L�1�jJ�Ŷ�i�$0 c�pU�Lf�ᳫ�2!Ҳ�vj�5�1�:�q9%@?�6�4iu2�g��'��ghoKR��ۓ/���[:|��=���M��CTm�V���Z�h�bm��c��0:xh�բ����m�� �^�ⴕ�6��7�ȪPģy;޼=E��{��n�����9���<NL�w����w+o�`e�b�!H�R<�x|s���b���d�۴U���(AF:+74��q0erڍ�M�׏ۯ+R9Ӷ�ش��\R(b�Ȝ�۝��\s��*OA��X9W�C'j�ծ���.#x�[o�Uﮖ즟{r��È�g-��
� ���E�Z�n6c���\]^->�%�1��r��ug��7F`e���[}g+	�������C�+����`}ː)y�^��sN�g����V2���t%&A|�y6��%�`��`<%���g�Af�}:��%m�ǤG4wJF� �v3۲Wj�eN�PkQ�|�&�I�ˉ9��%\}mM��\n�\n�X�/k_n�V5�x��2�ZKY0U���5FHkwv^�@�@hڬ�r�U{õ�v�*q�f��n�	*��=7����k؆�统,�إ�T�������l��JA��7vIomoH���Ne�҆p�~��+s�gv9~��#)�u�D�֊9�����<����)�*�`Y��O}�w�ל��9v"t��%��֡=�=���M�p9�����l��ѭ;���ҏj�II�/�h5>���Hv.݉�� �
�q�lc;1 �L�8s��ve�un�l9!JC�w�*���G�a��{�E�6�Ʃ7�y�c�u/�J��H�������m�rٙ
l7�&6���]�E�]X��V^��m��v
y/$�G��gf��RH.�ʴ��!��s�Q����X�}k������QGh��d�V���8��mB�0�e_t^�����\�c��a��sc�{E$���W|�K��D���#�e{�]E�	���I��㾴�}�=C���<�^P�\�W�Y�w��@&���v3Q5W��4��Y��VS�0�C�v�(��69fU��I����7��}�_,lV���������E^K3ey�&��aQT��9�v�Qw�<�l;�#M#8:�(n�903�N���HU;f�3Q��R�{������6�adLk�D$��W6�0Ȟ�[����v����u�aH5'^0�V���u��������n�KX~�������we���Ty��<�e�=�3Ca���`�����7�M�;���4ggUe�����Λz�>��r�,����W݃,����s��d��^��I���X��3e�:��?�+Pݓ��Z�v�
D�O�)~X��^W�|����)���~�S'�"�� �A$������켙[����[U�g���Y��/�ώ�0��V�M0���������+Un�t�ɢ-!PC%#ʳ�@��F��o����|�g_J��Ϝ�;h��拏�iC\�hާ��>�m���<G4�R/�nk�uu�~}�Lk�����7g9��{�r�8�]�[q��n�6rWbBư����vȷL9S��R��U7�N�<������Aq���7�*!o��e�Ƭ�oh���Sf�f̖��IU)��#�C<�e�8y�F���u�[�ԯ��%lNvk��Y�4���IU���b{����v��`�U�9ö�k)J�2E<S�B��5=�B���y^�ج[7�J�:T;W~򄷞�۞Օk���^lBo8�ʣB��oy�Z�P��n꛴��[Ӯ��ʕ��n]u>~�<�ʐu�ͺUl��7�"�3kmL/�9"��7ն����t+d���BM���q�X촳��u4oxS]@���Go�9ݛwzi[w��9�<���=���2�L4�My�oi)��9|���X��qm�\y�ۏ��46��m�{[�o���7�_`�csnn��[p]�j���{���ܮC�o�Y�r�P�+��RÈ��6�w=;[}���1�^��0;v�ɘ����Sf�J����Fj��i�+�9r���P*.�ΝǬ�ʊV�咒1f�K4�A��7v�Tz�s�,�(���|��9�r��m�Q�� ��\8����l����p�Gf�k�҃���7AM�q7M��r�j<뱊�ˮ��ڛ8Иz��Gw��.���snC]��c�N찗[W�f����/y>�5��C�
�խ�g
��o+�%�Ҁ���%�ݱ���Vʖ�TD���*�US)��va�f���u���l��6��6�i�C�ٺ����c�e�}ڍ&����g�e3���ۺWf����n�3�v컎�.s��\K�-'�h;j�X��6���9�')v�����;1�\@�C�.`Lt륲;��ݺw<sz�ۂ�1��m�����C�½�,Hۧu�:3nu�<���պ��xCa[\oK�q�٤�7;�1���h(�i�;���'e��'2�rӮ'�9�t��uq0�rX�R�;=�]��n�0=�3�:��݋���r��\��x��k"�1���X��3�WKٵźu���{M����V��Y��nq�M�� �yN�ܬm�.����1n�=	\=��՞n�vŶӳj�N�;&���Z]���=��o*�a�a�6�.T��Q�̜��y��5���ݵ�[��q����e4jf7]�u�ka��q��Nt���0��/��������68��v�u�Y9�}�x�����=��7o:{G]v�(j�0s�?}�:6��.�等z緅R��9����;���@4a;W(ܼ͋=�.1ϳ�tK=���-]3��v��Ͷ��Ǚ�0�p�L�Z�̜ؕ��Odo[/�:�=�͸񝁧�QC��s�8�c�6}�bm�x�;b��y�T=m[)��8^��Y�ɵrZ�}���5����n�C�붎�	oH��O:�vOB����3�z�zh�9�JOsCokn^8��S���m��҇�k�cq������ƺ�i3����{n��ATWmѢ�M)R�2�
0E1��`��NK�B
��y�]���8��;L��s��g^t�˱n ��6:�\иw�MnV�8n�es��nvc�]u�-�\M��WFu�q�s��S{]����o5��L=�����;���N�B�p��ಅ�.p�<sc��Ó#��N��5v��m�K�:�8#���[��N��m��v�v�%Y�7�Y�i�Pu�4ۗ�q�b��@��d��k�e�����^p��I��V�ӗ��k�xWJ=���]vɎ��gzn���H��ܣϱ��];��5��i�T]rs��74[��r�@m�ґ�P�Ɲl�{,v���v�L���u���5������ޱ�絸�Y{�\���"V����oWX:����o��g7�ۜ옩�qov\;h�-���Ϭxx#	�My�*��w�x�A��7gљ�a"��[V;C�	���:�hAI�p{�k��f��計��(�H���s ��b�VO!��X�n��~�1�¤&Cn
�j�nZ��{��(g�nGṽ�~i�'����[�ѐǨ��_�||XS����ا�U!im�P&�L���v����t���HG}O��Ś�_r���#����͍# �z+��.�+�\䪯 �'�6Z�&�m�uc����^��^{�w�<v�W�{��פͷ%U����_>���w�m���cp�>qD༭�,���w?Vo����ֹf��OfzE۞��ޝ�}�E�u���y��]����@����E>�-�����fܠO�\r��r"���N�ݳ��A��$�B�P�0}�Fyv*T���/���pL]�~�O�o�b�&�jo�]���k�f�����D�PI"�	#*I[׻.�b�U�S�:զ�ژ��˸��Ԗl��}��e@��Uhb5Ӹ�IhTR_Pg�==Y):��W����p%��M�3�T|�U����r�L?-��|�{�z����b`������j�ˮ������8g(�$C������9��?uh�2��u`�|}���sS���ǃo6}>�^,��*p���7�	E��&ߘ~��W1y_�%S}�i/w��A5?Z���V]s	ԡ����st�̖�i \���S�r�Oo@��4r6�o�)n��U�zz��\G/7�s���ݞcc��O��k9��6ޕ��-%�1�de���N�>���+��×s�n!�X�:����.@JR*�]����_jC���T���W����=�߁t^/;x��Uk�^�}!��T���NG��Aڰ�<���yA��#�~��x,���uap��w�[�LV���r��^��44����B�ơb)`�1ʠxk\{p{�Fx�~���lŶI���0�y�˳(�>;��#\�w����3�&oN��6�`���w����f��x���ǣԇu�U���m���7��Ǹ��0�r�kz��\��XIUŦB����T�L�u�9�����!e���*g���)P�-ZnE�x�d�/������� q"|ڌ�Y���
�{��C^_B��ALG�ݜ��U�;Jw�����^����0�!�*釆��gmV)�}T�s���9bmj��p� Q�eq�;u(�x	���u�͖?}�������1��Z4G�:�o4V�E����]�(����gfnYw��iw�I�F���~N�Z��~1����}�3}��ͺ#���:�Sg�Q��s-���)TL�]gH��3���W�Y�B�1Yn����'Yx������9��su�V����ġ�{��4�����Օh�g{���OR�e����y�����ϝ������,�y�KQ�{��cG�^SY�(��"U����>W3F\[��nG(�z���4F���Y��1�'�7o��\��k�-���`-�i��Zp#�V��y���Em�4�u7�~V�`�r��?3�O�F���I���Ĉ��Ó��pqu�}�
6mH�$DW��w��x��lf�DN��g}�u�\~�8��KHa�N�k��㕅2��ڍ�F{pr�9��͡����\c=a��\-�X��՗%���ܖU�l�����6hWk��(HӄF���4d4vo�U��.��ZE�ޛ��#�}�EJ��'>�8�����0(@$r"<��-Z�Mi����)��r,�;U��b�RD��ע����蘙�	�C�?.��#�r>�SJ1|�{ލF��%�aL�gG{pMv�pF���[��}4�m!e�xo�~�߾�Pq�]#��D��>�OlAڏE?'~��1p�rh�z�f���&8�t�n�}G��o2 ����SF���4��+��Sda	Cda?��zc���_�I+v�-�^�E���o.��(�4x��,O�w-�ҍJf�Z{�"GCL�:~X������RFɈcHy�&��Ɂ�MMӝ$��诹��\��u��K$��N�*�i���F�۶$S@�q��)���#p�Y9n�o�w�2�"�f:�Ϣ#aII����"�}~\I�*��ӂ`�"e}��vB;q�Q��Dһ��q&���k:�@��3���sf�f%�;C�6���w_=��)8�xe���)��Rbۙۺ����}�]����RJcJR�Wʗ<֎��D\��29TdbQ;1�:����BjJ;�7'�,��wf�e�ǰu��y�#�y&�s����z��8��h���ŕ��r� ^7<c�����oh(����x��y�!�]pn-����������n�m��x-��mΝe���8��9�m���K�*��MTi��	^�<�	���^ff�N�9ٞ`۬��n�us�S�pu���;&�3vs�1�R��L����l:��Z�)�mU�Pqp=X�Bv����Q~4-6��o���t[u�(�]�24���_M��|��׸H<ӭt�����DX_w�iN����	D�g���.B�(�@ݯ���O��٨�d/'s�B�W	����D��6Qܻ�_C"A��$D&���CӂB���r����=�6�H�*�63����O�/����<��"�Lv��
E�d�>x��D~��
��	?W��g��)��1���=]��v��4��+��Mrz��<G�[QUz��2!jH_
���0Ӈ7��?�*[m�@�>�a�9"���}��1a�9J�20H�~g���'W�#�~�$�dAP�G{�b�7���aӷ�s��Ѥ�1~�_a����s���7lUҧIk���	�4�h����dB#7ŋ%oH�w������B��8`���l޽��0w�"(�>>�#�}li����b>��o�U�a����v(*��@g�4ָ�[i@37�68��v��m�u��U����݈$���8?	��?{[ز$����r; Y~�n�z=2&	9���:Y�(�^�R�����P-��������k�������_i�g�����1��n*���#J!�C}߷���K���h�|e�i��wb�`Ν��1�Uc���W�]\!A}�r��wΤvl�uKʹ�����
����%��;�� �0�|��ϬP�M�!b�V��K�$�|F��_G�lOf�P"��@��zDz'ۢH�ZL���%���&)4KQ��`��T�2wWV����%G���KS�3���-;\�j�U�T;���u�B�ׂh�#T�����97��:�k�;+�$�q|/Љ��߽����>>{�udi��~�y�>hn�X��?����+�)��]���,����M�h�Gv���蚼']���Ʃ�6��nKM��C��#66l�H��!�W/��ʮX*'޺�#�o1D{ȑx��^��*m�!���<��s�N�m}�����'!if����~���,O�ʅe�-������qլ�f�Y��]W-�s�.H�y��yfY��m8i�;椢��>�B�`�#܄=�֤.��&��_\z��zwL�,�:<
}�C(ㆡ�DN�j�~��/��[�k�p���n�f1I�[��c>9�\RU�V)LwU����Z��*7��Ά�Y�b��5R��� ��}���mKHq~��gJ;�teSo⽒!�D��0Fgq�i���D��.!X� PP�<hɣ'�����C"�'���R0�D�T�=z+�~w���"w��V�t�֨�'X�\�n��y:�q�}�Ə%�#�ݗk�J3jYκ������Gmb�#���iRX�O��a������Ǐ�(kA�)�(����`�`�4R-������gټpM#�3$ٺ�ɑ�B��:_��O�X�4(�{��R/W�P(���{�L��$MW|�������pɯ�r#�p��D䊆���t1�8}���P���t���i�ڬוRдp�:$Q���i�����~���
*e��R�����#?g����b��~W���Lq�&H�Mn���c���r��t��@L��j&B�A�e@;��#�K*"��8YW�/�8Q�d�w��M���a��hoz�M�Mv�����7�R&ߋ��:ß=B��d{�Z%�Gi쏐���{9d�m���D	Gǅ�-�ab��v(�u��GH��_��ӕFn]��^�����WOO�FX��p�:��=p�����}�wa�H�wkv���{��"s}]>���ȋj	m\Ϗ~�ٟ����=�o�#{��/)�Gc��%�kފ�?{VJ$M��^oz"�o���~�4_zD����hq�Q�藫
#;X�N�����~)@�i�HR98�ܨ�.�H{���В��#r��C��h#�}B8fm�O=��uU�
8�w�5�[b��+"J#] w}F�WR���N����wsE!Y�g��&:����T����j��f�VT��]�[/@as�*��݋QMmvF���U�.�奄Y�Jɐy�d{&��w�tjm��IV��>�0��Ң��X����Ϲ}P�ڱ���i�ӹqTG��^��3�@/=�AyBF���:s��3S���'1����D����._4I�Q�σFP��L��t�\�����{] �h��;.X�9��m��iRrƋlVB�I+��~BмR�n��r&�8|ԟ�P�[�yW���0���ǟ�ą}y�˦�����;�bC2I����z	̡�{[���	��?UbqQ�a%zύ���/��H�p�ՂE��f�y��H��<Bx���ÏFxL��h���'�޺�ٯI7�
�Ew����DG�{�!�[zI�����&�T"XI��MRj>ˡ�̨4G�^�6F�}����{��0�"�����2��l������P�Zp�D��?��6��?Ig��E!J�\�?�B�l�$�iӧ��3r���Tk"Lf_�P�T�	j�N��ӂE���E(�)�=�#�*���Iv�\t������'��k�i5cٽs��*꩸�F'*���K4��GW��E�"O���+�����N��?��)��tiԊ^�	p���ؚH������q^�у 
�sK���h_���Q�6/\�F?��'��%�oΖ:�QX���}��/�4����ۢ:k�]]������߽||�e
���cn ]'4;�q�dvl�[gt���Y�j�u�v�ؘX:q��V����D���ͲY����:�<��3�v���箹�;X�g��P�Q�m��ʤ���wa
��=��/S9{u�V�MmcPZ���LupAn]�8|�6���Z8�N��{q��7a�q���i��d�ڀx[��S�����\۪x(��C�v�^�c�a�Dt��ݎ���	�l�Q}��F��b&ӱ4.@�`vu�������r�{���m��Hlh��O��K��k�uE?;�m}�]/��'+�7��"D܈�<M��YB�d]����Eb_�l���Ϗअ�a�Ԇ���Q@�����7bh�1^�g��<3��GuD�2Y����"�}!y1�D����p�GUW��"����|��~��cU�����Q�Z+T,�_�4x�3����z�^��q&��*1������$		#�ѻ��'�g,�/�������j`�	�!�}X*�g�2)�v~Da�+�Ĳ��A�0b!]��t�h����qS��kH���#O����1V��ϵ����0p�e�W��	jȣ)!w��G���͢*ktx��	ܗ�4������Q��ۈm���ɇ?aS��۳}9Iˊ��U;X�"lM��*��8kņR��8�"�Z�����]_�Ue`�!IH�w���(�B��F�D� `�����z��W�j�ILA�lWb�s�[�3T����K0��ݸ����R��`�Z�'Kab����%�B��D��임ߍ#�!D�x7�.̬~FA�R�mG(,ѻ;�& �wYh�!J�ϯ��X~D{��H�?���А�"�2��F�"=N#e��=�Ej��>��Wz.��y,��M���A�q�k�l\,�$�o�������q�:9�X�i�QeuǱ�ϰo%���Q�u���-Ji3%�����1�#9Io��ӏ)����'�/1�z��'u\�>^��H9�D<d���_j���ʄ�[>m]�1��!�#��)��ҁ�� �Jf޺�9E�;綣��ֱ�~�C��������Z���)�J2Q�'�#��~f�!��E�RA_jTv��?fw�F��`���ڑ���"!�dQ��W�蟶/
#�g����^�j����&[쉽�s��	m�܂�ʜ����l4�d)R;"hV�����,�w�n
�M��AH��:�d�4D�4�}T�S��I4x.?T���`��l�Qd�_ �ӞR/F/�1�_$Bx*��c��/���	<���W�Z�Ԇ�Tm����J+0����Y�y�W�Mq`���⎍��V�ۃ��W��x9�]m�P!Q�'ߤH�$7�GU'v^y�o>B-
�9�0�	d�����MFz�}��"<A�>AǷ��rc#�5*m4)�ͷ����al�t���|.סA4	�{����Dwc�<!��sȐ�v�[��u)+��B�k�6_Xɝ"�����w@~�	��H@�+n6x#��N�<`����-X-��2@)8u�b����J&����9��"!�����z�
;Z��}�;��_'U]�.���vG�k��b���RO�6�#���0LОI�m��Wm�ۆ���1<�Utz�i����IglW�wv4(�EUa3�l�9�L�/3p��{���5����������3�C�6�7���z�a�CA-�EZ�Ra<s��Ҁ"�A��dJ��C9�?_4��M�*,�źZ]�V����s/>��k�E�lU�rZX������([.6HX4�r�5�ǉ��Y��_sr.��
�u�n��&��R��)�Λ|Fm&��Ȓ�j⫫���fv���X.�Y+1d+�ܮӞh�񝢲�p�#�7�j��A0ۼ�z��LQ�%j�e={Q_)�"�h�G6�p=yKJv�Q��u539�hb)x{:��jo^�^�DFq���]_����k9\��A�[�1<w�.5��մo�����ć��%"��S� �Y�jj��=Meݤ�Γw��tT��������o,��4�Z����4��q�k�6�*����l��
���ԛ6�&�������	`��2��eDʙ����
��&���;6�3jԌ4)m�њX�%L5Ӳ2j���3j�6�9��r;{=o.o7��YBe��Ȝ�7T��b�R}�"��+l13od�6�.��磳�u��+7�.��QW����Tt�9�s���x�-�+v�QĩڮE-�W��Od�
`�"}�:�W ��u<"��q��
���af�Z��*���Ç{�B�;����k]d���5�$��'���U��u�jl���T|�	�v���)Q�B��8������z<�y�H��~�A�z����zĊ���6�t�l*>Sr*�B�"Hr%j�H*�q^q�t�Y��W�TF�!rI-1_�H����ں�|.�v.8k�ؤi�VQ1|��
��<5/M禲����r��Cj=�D�������#dUϰM8Ff�}da�No����7[��{���-�P�����d�,M�7lu�3�k�$��[�ň������һ7�:�,�Bp=�|��I~������8E�P�dяT��8�"�R��Ҩǽz$O�,�d`qȋG=�2�E�_G������'�#���m�+G���`���?i�a���$E���C�L��B"�_��\/�V+�P�@���#���n�E�#H��DW���
8Cϫ{gE#�����;������?+-�Tq���a<E�����5�G�����Z�>��)~fv����'��Pʺ�#����ZdG���q�f������͕��g5���䴶+]��il�~�dI������rЍ�5�nD�:n��èL���~�Ρh����L�O���<�4�F��Q���f*�0�YJ�V��W�aUl('�F��I��Ů�Yf�jv��K��b�O�a�*UM���f��e���]fG��v��RԔI��>w4陉P��i�}�<t�0l~;z&�:I����ZC<����'�^�pw>ȑo�bGĔoPc�[��Z�(�E[�L�O�P��0�2A���܏yL�	C-1�Iw/!��oY�kA�����c��[Vڻ��]kWg$ujU�[v��9jn�������H�	���*Ԥ�}4�~�Y��b�F!�L�f�&o��G�bF]u�^��k!�#�u�����M�}�p�����@O��$�jDDD�j��u�
4D�W��+�»��gЕ;W�F�a3��h.gc�|d��fb�z�|�P:У�&�0I��xϏ$�moO�Y�Lo#N@b���:;�U�H�v�y��gM�	���ҁ:{���)���;��~����*�K�5�J�GB��ۊ��/� q-������f>�Th���X��Q��IO�1�x�C���J����!�ItE�_�}~��o��]�z�$ȝ����S����	��ѡQo)�/<�/º(�q��Wz��U�^_6~A"��o1�p'2Z��o�t蠴L6?s~�6�<t�`y���_��rݮʙ�R���YP��$^�$g��'��쩷5���A�0�;{o�#���(l�ہ4��yS$�$
�|F������نv�1Np��Ԏ]�zy�i��[6�h�����p.���K���v��m/d���na��l�k�e:4v�n�օ�t�3[&�p�i�<Y�P�W�.�uy��s��yHk�l�.%��ܩ���}���G;�[��i97/+B�Ӻ�l�m�O=r:���-q��	v�Rv��⭻{q��wT������Z�D�!AH�蕧b�>��cm=���Ȼ�z[eŧ;�s��<<n��ٱَՆ��h�.#m�P��k���Чٝ���L��rx�u��u�<H�Y�P��,��N\m����J��\�?�e����*Q~����6��ȍ�M��3�<�b�1�'PF�ެ;��{q֦Іm��D}۞�(��H��R��z&�& �ܫP]:Co��fM~���q������%�,3f�%u�rN�CZ)	5��l���C�x!�0bO�̢0�{�8��*�1���Q�ny�םM�ʉ*%�Y�Z�gI�֘8�yС����?ek^���)F6$f���3R�s4���!���E��L� ����	��"���j���}m����'M"��N�9:A��}� �Mn�e
��gU��DIi }��V�$[Xh�)���u�(i���	3���_`��d钩l䌋_fgsM���$.I1��x��}� մ(��I{h���$@0�NV�w������;�(E�e�9��پH�N�ٞr,�f����� �k�Xd�"�BG�z��5y��<AN���O�x�����X�;��.�Y4�	�Ŷ�Y;\�D�;�;VۗVLv�V�S��qG��b��Z�r7R��2YEr�!L��s��?*K+ㄑ%�ϼ�LF�fU9�/��ɸ��H�Ń��:E�G����̬?V{p�۲C�&�|[�CA�2&�y��r�]��3�9���c�Al��#�·D�vXg�##�b��٩���h+�Y��a�*\����M�����)L��,�h����|FB=(�=�20�p��Ec��&F��,����E_�]L�6D����A��^0l�륍z-8�e7E�y�Q�pTl�a7�B�qg
�`���6�}B~�BH��Gƌ�8'! �z��;���$������>ɯ:�/��#��RX�mӛ_����0�Q84���.l����h�҈[����yY����/�hbC���� K�W#��G� ��y���J�C�A�<K�sXq�Dl6D�Xd�)O��~v�[d��Wz.�P�P�?~Z��W�D�?������b�d�)�y�|Ef�Br���yȟ/��#�-B3)w����Ӳ�����2����uE��Vºc?���A�RլVfN��n�c���YW6ݺw�1���:s��G�͸^G�d���_Qg��u�h�L/�B�MR�O��v�$3ˈ���Tࡺ}���|2���8#:Oh�5��cH��*�!�~E0�E�#�㯴�:A��C/��#G+��g�ժ����G�h4}Ѣ~�k��<DZ���.���Yu�F�`��^��[�E�G����ӧ¤�i���@���Y,�lQ�Ͱ���h�[�^�t�K�@�H��0/�.�5m�Z��$�{�����V+L<Ѫ�F�rs��P�EW����R��u�n�:����]΄�ʚUhqwF3dO��a��:j�H�^"�8a����Gw�|ꦫO�XçަaH:UY�%&�"p�M�Q�����Ṍ�e"f�>�)��z�e$O�z$�=��7Ѽ$p6D<�zЋ�S�8��ǈV�
'�c�W��z}'��'|(QĈ9)��%F�����%>� �<�~B�!O���>�Ə�4�($��|�P���;�r�N�rȉ:�ўw�E�@���"X��Q�d!��F���֏�'���~�H�r�����w`8ۀ�\H#tm��G��ƅ;X�7-�;/7�*����8��K+(;S%�~�����[lEV)���S��P�� ��L�I�io�|'�ci
��P#���1L�#��I�8�#��~�<t�
�l��H z��Dd��"J[-����t��i�=�(ዞ�k�$��<+z�񝻿U�?v�b�~���R�)|�#��X�#HP��c�D�������Z��������^*�����	�E�Rf#q	0
+D��M5m�a��))�Q�?<
�1]u%��*�ehFQ.T=�:��
D��č�)�h��{��=+�:+��:kһ�l8p�'	��9���.̓��7F~�{���&��vI�&�ur��2����V��I�!.?DY=��8�B�>��xn���y�3enG�պ��uԇ��\�BAg��WNs�u���dsM��ʹ6�;S��u����s�
+|��>:�ď@��Z��� Q�i�D+D�;��G#E� )Ik��҅�@�.�~�Ҥ����(�_e@�6y]!����=��+��b��=���귔*CX�ވ�$Ǫ�W:E��$�Y�M����4�����a�B�	��@���ѹ�ٌun3v����c˺�ڑ�g%8Fd��$�����C�OH�����7��Ξ��/�9������~�*0���G̓�y�o��N;*"6��#ec�X*��G��L�'RQ�u�F~�cv���o>>>��?E�G��e�9.�~�z:�2���)!`�<�*�ӂ��8ђ0`�QҤ@O�� �4p�2�&����T��UF
;:Ew��u��R��L��b��}>�8��X��o�:4��L�2bk��.��g<�_l1P,�Kղ$n�@F�N��� ��x�D������#G(�	"�����mګ�#Hԡ�!�a����ۂ�,4p+�4���q���bK��a�zU�9��I��*��b��^k���&h��pz���:D�Ǟ�����5�5}��u��(�cH� 1P|�F������(��-¶�\^>GN�a�C�����י��u,����1��˶�ج�v�O�5M��4O'�HwM��f	�oe�lӀ�ed"b=�T����E�uc���!��L3�l����ԅU�z�@b˃6�t@|q�]��]��.��-��`{���*>�u��YfAN�Nj�����jhc�B���)Gr��^⫮��F���n����m�F��`:��y��Iǘ��'h:ӓw5۷-t�����nz�Ü��Ϋu�秌dY���ӕy�=ԋ���q��j�z�ndB�V�l6�)�����{r<�C�훞��x���h���{/@��u�4�ۥ軬i֎d/Uv�sK�ݫ�zԢ�c(�iap�6�67K[N1�t�cGZ���h-�.��=����P���˫�x�5p6r��K�EDMYQI�+n��?�?V�i����x$a�c�A�t� �O����BM�q"iH,��6dyw�U�R={�=�=y� H��L��[H"6w�#�%,f��_wyb�0b�B�7��B�覂���	�5�����K�o=�-'9����<����k�3YU�1~��#'^�F�hkD��K�/X�8B*3�/:z�'&4i���A���#�$j9R-&��[·��C�4߲,��}#"���b3��H���Y�*��)�"��ZY�kzOi��O�
ԒD��`�Hٲ_�EQGU9$�=���+�{ ���*pd�٭���-#�O
��}���E�ez|/��A�`���Fg�@�_�$e?�^�����0��R+q���]"�Q�h��ӡ���J���=}]�e�A�9�R��_��⍆�P�"�o����H�Af�>�G��8D�<ƿ����_��w�s"|	�?a�A�!�z��>s�$���UT1)|O��b��0Y$C]1�f���;�N��� ��&��p	�-Á��6��]���^v"��qٴp��Q҅N����#��dlv�$�}�~!i(��>��t0�)QD���Ab�B�鸑�>��͞"��e�;��P	̎�驞�!�AD�[)�zg�ɡ:~�uE�FD:HL��m,0�u[�Z���(���淇E����#�MG���`zey�M�ԳB���DFEk8��1��n)s��WC��j�c^�9�LX\x�Y��-���(�	��8Fo5z�~�:�v��UWxW�ϼ���d$�4���X�����ئ����#�sΫ��@I�T�z|W�H��TH�&u�q
Q
(�qG"��2H�^h�"N�Ɔ$jz�����i2{��+OA����n�D�_os$�uX���HFL�-F�Έ5�U��2��BsO��}
0�LI8�bĨC�4��/z�QR/��z���ę�rW?��
��Qͅ�A�KҠߦl�u�fPcs��� @�9��2����Ok�,�-"�=b��%��R%P�qU�ƪd�dY	w��^��	��ɔ�T��������@�_QF�g�����n2 ��8�yE��芟U��f��N$v9ᓃ�%xo�u���~B~�����t�ⴘ����oFݪ�i��nӮ��v�	1�u\u<��	m��?��m""��/��xj�ԣ$D��e ���3��
�/>D�=�y�yN��\tϚ��Z!#D#�,�V
����	3R�����qo�������8Nc-5i�]7�(���S>��k�^~G�^O��%��kXfN�lW/�r�@���9���р�plAz* ������훵B��*4[����A�>�k�w^H`��J �;�s�t��H!Z����l�{�qE0���ħ�d�^݁# &�&����*}�\/[��K�6�V�W8�ڞM��.��ʛ�9�{�ۙ�� i��W%o�u2bg��������޹�3���I6�ȴ5�$�6	�/ʹ�1��8K'`�R�!�N�6��!Z'
9*� _5W�^yܷa�xDU �� U�k̗xE�%"8��T~�x���N)��0
��x�6�N�DI��Tk���MzZ��{oT�|�70� bG�`�s�\����L(P�l4p*���G��fS,�u1��SGI������5^;�X;^��		���)��#�(h�G�U(��0�yYM���ʈ,�T6A�iz0y�^��D�$����K�t����m噺@:��xg%l�׌�n������sգ�k����m�D�+�r	���f��t�GE��¤��VW�
���$�a�$F@L��H�ehv��E`�����ۚ"�ʩ|�?�2Q�-��z�o�M���U���;*��9�2�����!��-"��{�G�d�*ϔ����H�[i��~��"�u�b��gH����K�)ϊ�&�jDI@��yM�N�,(�B�A�GAN=n��>��iy�;�( �t�8p�_$	JץR�2!���>�W���9q�U�"�\�B%����kfnZފ���<��H��'f���e�� ��4�｢��"+�GZG�82�Dŵ�.h�8�J�n�Ӆb�:��E�I�n�a{^�z�8��8�<��(Y��LP;��1�v�~=��$�G�Ɇ����?����>��&�`E!?}Fꭋ%GU@/��~".��<n��6�o�f.�<���v۳p�/���i�1t��]���W�d��l���M{�$
��)T�8�C&� �G�eh)}��!�)]�ZqpA���Y�wi�3��B_z���d�2%"9T���0����CA���_�
P@���R�&�ã\5�Ѓ08������i������6��s��|׼tE��)Z��=�uci�y��u`�.�Ĝ�mG	�#ywG�Y��U��-q�c�VYi�u���e|n�S�+�:��0A�Aݍ�z� �L��D�Ag�e �|B ��19�SF�����-ﵳ����A�H��$���B`�x��R�8����)��ȇ����n��mo��")N"������e|G$�ՇN�J@�v�*#�������u�至� @�H�~�Tx��Ј4��>��T(b@�V��es��)A�`��ɽ��mZ�-�$�o�o��	'�H��<��UD��
?>��Q&����~�����$F��E$os��T��Q�Ï�� ���|�#3�G�(!� I?n �:���ֱ H���M�`/	������ײ W~
$���G�ď$R˥"H��#�{��1#�~�4~��j�D�]/�E�&����J1�s�~z؁/� ����a��oI�s�T(z�:��%[D���^m/Vj ���߿t��O�(%��0#b�%^=�wO���7Kc��%��A��Ğ�1q�m�K��01m�_~��V���H��3��H3n�kh��'��~��U� �C>(ɪ�3��i|e�ُ���Zĸ:��I,Y���ĒKfg��$�X�3?�$�,�ǉ$�,���ĒKfg�,I%�33�8�Ib�������fff%����bX�$#31ff%��ĒKfg�,I%�33��$�ř���$�,�ǉ$�,�άI$�ff�ĒX�3?�bI,Y���,Kġ���3��X�Kfg��I%�33��$�ř��I$�ff��d�Me��80�O~�A@���@ ܟ}��s%m��b��Q.�v���q6��XTV�UMb-͉�T)H���� ���j�Qf&��U��� � 6�SL���>��    >��7�U՚�[M�m"Ece��([J�,�mmC%̒�־�X�kJ��=n��#Mm�eZ�U��	�����a�����˵������n�)������Pʝ�(ɥg�z�����9�������=ϮE��rg��K��{�:�}�Q�4ޛ���ۻ��ٛl��L�o*��US+p��B��]�B7��^�C`  W�   �\+;�ǝ7@��byZ4�w�q�FU�nz�p�7\���'[����{��˻%�r�
 '� :����s����U��m\<ܫ�ˮ��^�^�ʆ��{�}i��:�[����I5���v�D������Ɲ��o}�/}���j�{����fod�r��{�	m�y����愮�F)M��oQ"+�ǛR�7���t�����z��8��U��mR�=wP^T�תn���|�x����������S�i)�7���<�v^��k�}��c����;���m��c�;�����5i	i�wu���m��r��|Yz"���{^p���u���Py7�aԏf�k��}�F����t��T���oO]��ӫ����A/'�����g���ƚ�m��4]��GRv�f�a�Ӱ^Y#��Tm����|U�J���zF����8�D��N޻�﹡^�N�;��e��=ﷁ��O�0�{��y�ݼ���=f��T4|�4-�i� �@�G�f���+}�{ۯ�r}{��,n�>}��hb��1�����q��.�w�ˇݛ�,�;�
kΘ�N&��;`�kz7Zl�����O;�.��nyy�P=Ϟ�yG���z�+ُ\���
������!�O}���Z����n���i`�&��w���u�zԭ����_ �z���Z���'ϸ=z�{s��5��{��n��7�<��y4N�����m�;q}z�`�8�m�N�z�����wz�֛�{�}�����I�int�GF�`�lK�M��>�����w�w�=��9���=y�Y��:��^-��Ͼ���F����u�/�s�n����Z��{`z�� "���b�R � O�bJR�0��bh"c*R�5@   �?���  j���$Ѫ� 	� �P�%SMI��4 d��/��=�~�������f��S�m�XB���woZ�%o�$	!$����$��aB��$��2@�IQ�$	!$��� I	$��HI	$�Hz��{��?��e~�_���C� u��Ts���w�[��w&9[Y�-�b�!F���,̌���lm+*<�m�w`�X�x�V������&'n�ܺ�%ڲU?��o&
Q�TY�RRбU]��s���n�&�Q�A;���Nk�/D�[�r�P`fL�Cz�e-A3o^T�ى�#C��1-5n�(KSC�ڗzB��dYgeP9[a��
Aah$�x�%+~��mS�*��E�<����3:�s��o�$�۱�w�$;�Z+1�Q5r:�V�<��l��,�!�U���-L<�*5�ת��ƛ�+�J(�5����mM�|C���`6��iU֭�.,q�=�2dŽ��31Z�BmJuq��/@ ]��Qӄ뼶�X�eA,��(<xv���h��,�
��x�x��x�qC�ܨ.��t�ۈ*�Otj�HLvp�ϭ^�Ζ��)��"������5��7%�bE�(4o&���c���%����~FTEV�~'wk.��i�*lr�eři劲� fM@����c�4t��-�cf���jAǻx^�2
���5qnQ�\,9h�3���w]����!iizS3M<�>Mi`�b�ڎ�6pGn�U�ɢ�0G1�5�t�����3��X/#[��K��I�k��\�jm�!�XM��.C���6����e�^��lD�K.�!yf�8��I�<�0"r���V�ϞVVթC,8*��eh�T7Br�G�=�U���֨�=.dp�C&d(mV�)�����S ��p��˼Ѫ�Aְ��Ld�h�0�������4��c^�D�r��k����\�oO�Q;��A�ow	�Ʋ�0�2�� ђ�C^-:���@>TqS��lp=�W���ɖ��ΌZK�Tq�Yg,o�49e��+�/�b� �0]�+,�O1R!���đ���rJ�4�*���u�lu��4�j�8�ǨmU,݆�ڂ�C`ڙp��<B��F��.@F�":�*J J$�/3ÆƉ���M��"�n��ܽ�Fu����Hc$u8�K��N�@)]���F#1�yf ��+M!���F��xq;n�r��0��@r;
l��)
hkF�=/H�63.�6�f�C�孶�d]I&��ܒ�ʏX2����c,�p�2`�J+�<��Y�Ȓ��ú��c3mD�D�Ù2�ð-�k����z�"�H�w�i*�(�k(�2��F�+����g���=�w�ȈS/U4�K��̠4��7�n��řb�
��S�����-h2�t 7�N/w9�ꐚL��B�����WS�t�>k��i�'��(Id���l�T@30%�nɼ��e��� �[9'Z��`�h��L��V����+[�]�n.����u�]k,���.�&^�-b��4�7R:�Mn:4�N$�o_��H����f5^��;�x�N0��a�{�h�{��ۻ���p�<2����D+���W�|v���}����^�L*������	=��fnp݋._]tY��� $�]V��B��s���Q�F3��睪��Ht����|�u���;��v�E���5�&w]!Y���a����WM[Dv�Z��]|ٔ���L\���yd�{3\2�!i&�A�E����9z�����8�hi��w'����7x��$�*����3;I� �!�n��+d����i|!������D�����PuZ��=A�@�rW��e!uD��;M}�/�;Kmm+��/u!���V��y�V�W7p�!��Q�QU�k�o���\).����z��������4���\Aʺ�)�3��5����pQf�ʭ�*��2�f�T�I��pn���t��Ý�/;/o�Hhpl��3�p"q��;E�����Z>������\*x�uY{d��S�^|�A0�k>ϘB$���~��O��tv�!*�&������\���=�o*Wp�j2�����}�߸�p�Kʮ�86��v�����l4�<̡�&%mm_�Cc�V��?��ҫ:�e�T�
�(�]�dA���Ѣ�m>�`�����8;��Nq���dE� �7�e>w��Z��M��`P���smz8��u�7��V�C5�����8�
���J�FU�a3S��m��Q� +kT����k�Ż�.	���;��'��/k`��<�`r0�j,t�� ����(fUќ�U\[��s�|��,�j���_P�E��v$�3+n��o��LP<ǵ�"�I�i�<'��Y=V~o��P]��u9��o�%���d��96 �X����h�4��yB3��y�����dD�^S0��C�-ΐ0��O���oYw�N}/�����ǕɷR�!"�|�ںj����T���ݤ��Վ������=�d;��Bͻ�{\��߆�����#�c�2i�2���yR�)Q�n��J���q�I!T���w�Q�p�//#�s�-r<�1{[�@�kU�0���kl �4ްU�+԰�_+rn��1+R�J���Z]STm�t���Kln�U�଴��=��Q��l�t�V�;b�ǒ+2;��nel�^ǲ5U��9{n�nԛ�2�9j��p`4Qǒ�i�N,�Eb�F�9�ʰL�Bc��a�
�v�"�x��{N�f�ʳ�Rڎ�u5�m�ϐ����ޖ�w�ՇN��#M�����(�Y_cOj9n�*$Ȋf\��4׵��n�� f������4֪F��kD	R}�00i�/HO(n�Z�4 �M7��܂^�֦q%k�&�M�5��;Ud$v��u����epA��D�o�R�Iy��ݬu� )�ǎLI�[� ��m<�I�Ӣ�H�X��+�c��*�+{��t.� �j�G�<Oj�}T��.���ɻQ�y�^��e�q��ق�P[h�A�.�K{��5q�Gv[��"*Ɔ��ޅ&���Ǌ�[� ��=ݕm�!_=`���f�] #9�gm��Ow���sN�JP5�0U�sl�N�m�*��h�^��F �Y˻GHb�bl;m;z�����G[��W�vJ։;�*��i䥤�F��`�Ha�ĩ/v]@�o0c�@)�u!*\,���3�Lޅ1h��uw�m�2P��ITιHAcݗv�=�VU�&k��ѣR�XR���h�SLM]D�2�J�ӥ��;��7gl'�V7���kli�SU��PP�v:a�20��t2��b9��;+ �r�*�ð�!�%)(�Ś-�<�j��y�w�m[ZZz��˂Z�fH�S�J"��PYQ+h^�T���H
�M4�q;��9��M"�)䒴` kK
C-��<K��ɤ�L�X:�e�5љ/���?���B�u���2�k���Y� ��\y)f���Y��v�`U4�m�[N^)�zv�;���Q���I3]7&!SoXYCf��^�4��Q�#���V��1s)��Ɓ۷��q�Ƅ��"�L�Px�P��oJUhl�m�Y �p�S36��K����Un3�+l*$Q\�ֆ�㗚�6�1K�Ԑ����+@�K.b��2���:�U�ڴ��b�J��e%B9b�tFn�j�G	\F�r[W�1HӲ(q&��ٕ�(�Fj�)�Ř�.f��0�R(ĕຂ�*�C֥a@�/r��o*���XT$`��v����s:ګ-CT��7Xɀ�t���32iyi	P(XT7q��c�9���'�l��MmB�ݣ-���m�ŖF��HQ���o�ha��]��KSo^hEk��9��%</T�j�]*۳MU���)H�$�n1�r2wn��eZ=���f�Dv�<���KD�{�����N2g�*���7D}:��Uu��L�ݹ֕�{2��Z��P��6�Ky��)x��ӺK@X��T��+~ůq��.�X�F:��0���j�d�E���AX3r�aT�wf脛�6!Dk�qGe��k	`Պ��قP-���P6G���Nʥ�wT�0b��V�RQ�uw��l�6 �:��ֈ�S���`�RP�����rE"2���/`�,n��-,��c(��Yz�eԽ9[���*5���
ݫp7�a����Y�q�^�AݴP{֎�ı��$�S"�(�8�;�<Q��h[JI]���ε[�`��S�݉N�-���N��wE"��PMj�e�*.5�l��P,4�A`���)PD��M�J�%;7�/u���`���MDC+�
`�Fm)&��PDD^�(�� �*���AXUՆ�ڇ�ȴ��a�b�yJ��{��f����5ǜ��ҋ��b9E��tB��6���,d^3}�u�ti�]W��F�[z�x��m!C<�7� � B��R�pC��ڭ�.����"�/[܍��ů-�(��Y�����V��VE�6˃RHG*�Hf�7i��̲�h�Ek�c��� ���f��|���9Zcto�(n��MU"��(c�Q,�p�`� �P��DY��.���e�s�+TrVe�(����wz��P=RͭoV�x|)TQ�a����ѯ&�ݹD]�7RwE�7���k���T��1�dVo[k��&��7&-�����[5z��+V�vl��v� �E�ͬ�h����#�赪�]�f65;۠@ҭ��ӑA�iK؎�m=t���onS�Xb�k1C�K+j��(U��7w�F�����t�䗕X`.�1&:(�I)�O/L������ �Uwa��Q��S;�M�8�х�k��B��7"�_!L��RF�� g)H��6M-�/X�A���e�hD��Em�J���X�v�M���yO6�E���!�N$>$�H�|-0)����IH�R(/XR��
<�E��gog8��ܬ��Z��&�<�m�g~�F�e��{`\Y1ݧ�ڱ�
l@ʺs3-�A�{s�7YNʠ��KP7�#3e\�ջ�F��N<i��i��)�+L�Q�(�r�Up����Zaw���N���M��6���	���?r���hR.�`�`SH�J"��e"��
`Ci)�V��搦Lw}�i���;���ꑈi%<ͻfZ�7,�b�8B;,T_%�ʚ)ֽ��Pm���ڐ�(�Ee[�a�m�D���	(�i�"�Qm�];��S5l���՗o4�PE�4�����Ϟ;x�NY�={J��0[�6+-L���t�T�P+i�
�rRSd��h�v������5�Ӧ/<L0+���[�������BO�؎735��i�ʼZ^k
j9B�k-�5Ӄܥ���k�>T�;|;�|B�r�R&��L��VO�}y6Z��Z7�[�T�C�D�~��m��f���6t^�	x�F,;�4P�~D:1-���WSn�V�?�r�tv;JQ�P������`����P�?�A[�çD�bׅ1a��7��&�Q�B�i2h��v�S����`�

F֨.H=5�*�d�e�b���	��2�J�4�B�՗N
�k5lt�*�`,rd� �vVdz)���lSY2i��J�����o0Q�Bn�;�u�x���tV����*h�x���\12wf �.�F�N���b��"^�Y��PN/���9C�$P�M��e�8��ʛY��V�7.�е�/N�Ē�a�����&\bA�͏M�u������U���VB�wM�Rʫ9��6�F,d� ��N�j,�n��N��e�mSq'u��Lj4��)�K�4�SX�)j�՚��!�^��")�î�^��/5�C:b��E��:�<�C���!J�ܶ�����z)���TF� e����K��T����ڽ�����������"˓r�Ţ}+%<#�ݺy�"oH�b�L�HJU��1ƂW���͂�D"u��k�6����W�ڱ�p�M.�7F"����LJE�"A ���b��V��R�/Z�ȳC��Ej{�.���Э3-iṿ�6�z�]�e9+e��R����6�N.���:�9��� ���ѡ��pBE�A�c��:r�<T,�2�M�t�?"�K2��� 9Vn���@�� �&����=k_�5F�Лv!n�-��[�j�	;AM��P��]���aQ�(���ưJݲ��GmZ��$ m�zhl�����iQer��iU��A�(/)��5n�2>0�P��u(豄�ܶ�9h撓ڽ�4F�t�^[��=Z*���ɉ��4<�R4����cV㗸��"�ޤe��������/U�2�J�j|�����nbܯ��'KҰ�cV�Pr����,Ull����a��*&o5��饲R�Ic�iXs$T.�kE���B��eD�X'"ہ�^Y�T��K�F�M$e�h �8M�!E�9�v�XV�Y^�>*�p,�b�>R��M&%��m`��L��0�2䶲k1�xv�1�͸�{W@��
!r��q�hK�dn�f=���c"�4�i�
��&�Ң����h9բ0�J�]k�z�˂�[7,�5�[�w��2�*'���Ax�b�+,�F4��$so��h�;ᩴ���d�S9��;}�k5���+@#v��eD.�U��5[��I��-iZ��=�Ev�t7��h�Z�P��GD�2��AHm���M�y�	���ܗ�w.* �*���5$zs]�wQ�BYnVR���7�oH�k�ڿ�I���8�M�v�7c*����Wm�U\�J�ȍ,Uٱr��`�ۛ8vP2�@�Um�m����QU�kWm����U��1TU�M��v�@���6�U�UUUUv�UUU@UU�m�UUU�eWm�v�U�f�Wm�UUWm�U]�T�d�eU]�������(b�
���ʫ�W���
��h6�.�*���p쪮��͕Up���U�l�vV; ���*�m�J�n�*������dv�a�]��m���Ŗ����ʷX8��gL1vuWl��U����ݳu�-Wb�h� W��^eG%��j��]�ڊ��@�]�UU�m�(쀪�gm�JՃ�v�[u�l�u��Mn�vΎ���\Fj!���8�E�]U�ҫ/H�m��5�])!������i�ؔwY+v��4M�عj��.)m.]e+t�mM���Z����Un�.k���[�!���[.�%6�3[����B�m��C9�\t�GC7����3�Z�S7Z=]f��bk=jXh&身��YZ�ZFUz۠��Τ�VS��9;�R��w��6��J�wDe��;R6[4z�Y�֠j+i։lo3-2�7y2Բդ�l����f/Rݵ)\��Jj&L9�c�YZe�c��8�����K5��t����Z	�l6��̕���RҮ%�j[��k��ն^����3��HI���:�+1�ՎCkff�����È�`��YR�!f5��L�15�3��h�.t����}�5�&�
G�F������xhQ�f۝�_�LS!�������K-Su���33;RԹ=fq�-�k[T$� �� ݰ�V�2�����x�c�ͦj��cũ�M$�X�u�d��sD�R\Z��GB:"ON��Qf#0��R'�U��r�P�8ր�|CJ@Q.6g�W_$���V=���mS���0�$�"�^��ԗ�'�o##ߛQ%�@���^�t�q�H�7 �X�ۛ��������0�`���m��D�󣁆�9DX�q���Wȕ���
T%,)���	G�VŃ(d�q��p,Y7,�`̐l$X4b��u�]�(�`����f��T�d���v�r�S.�j�]�`����V��Ay�WjF���YW�w�a8�o�u���y�p6� Le���u��-�;�
Wf�
�wN��enc 1˧3%����4P�("�Օ��7�@	�8��X�c7e]��Ŗ�J�chk�j�V8����Uְ�ڕ��Y&B�\�|t���ȫ7C�(�H[(K�'y�$�M���
�5�{����c�2���](&=��G"Q8/�B_Ԝ�����\Q�oZe�����'�}bʻ�s��H���Y�e�KYE��� o�d��/5��31�Vu���=�!%�
9=�� �Y�K]��(U�a(��}ι�M���R����`�4e�2Wb��бJ���nY�mR$�[F��	@[�;�=�����:޼�G�Wl������ub�<�-�yk���Iˑ,s��RWN�A��,B��Ih`�h�� �C+o �6R��:���ua�@�n�m�ʺ��ǣW�:�e��4� $�ۖ�e�SOP���E唽�9�i�t>���o��钺�[*̙ް�p�+��[�v2ni���N�ǜ��!��W�*�����S{�m��Uaێ��zN�A��uV�âӴDy��wY��kn{z�*4�M���"��}�����jzRܟM�.ۥ�֔{�	|�n��^��ի���QP�\T΍����9n���@����D\B*����*�����t��P3�畐S� ݳݗ�%�N�;	wP��Q�U��ռF��n�m�S����9B&��o�tZ�J�76r��;�D
Q��j$zh���S������E������s{��kT�'R��:��Q��>}M7M�Ο��5ɦ�otE�S]M:��Rś�TM�Dq��O;�)n�f�<�a��\9�ƒX�+f�*M�m�l�1
�Ý��R�wv!Ґ��e�ڦ���w��s�2bN��3���OVb&uU�{2������|Z+5NڒV��Eq�P?�7���jf��h�[�K#��7�'��!��P�cp��q�rdڂX�ܜ�Aj�9�95���@�7�ç�v�[R�CQT.z\&l��t��j9EdV4���i��ӄN֩	}����fc�n�˨�t� �e�
���0os�5�
}�O#2���,e�C��'��̬ճ�aD�V.�*�qg��s�ŝԶa��(���+Mv�ܚ�J-�עb���K���7U�0�ufS��t��>�)K*1;U��I��[��܆Xy�F�R��P�ҡ�7��"�v�s�����o��$[~�cR�kȡ�]�)�2�6n��j����M7ZJl:]�I�}��1��JR����y!����.gR����*��a��܎��v�=��[K*&Z�hI:�j�{sZ���/8��d����i��a9��e��n�7��W@��C/rh�'s)C����UN=1����GL9�xc�A}�#���
� ��rJ�壐���p�f�0X|�v>x��W6Ƌ���N{5���[���}I�ÇWX������S\��M��c�5�0i�7���o@b|�����w��1���rq$\���\}��WJytGd6�����kk�ì�1���YKK�zb��M�P��j. {����,�)�3r��i���9p��-��(6�W�q�,`���hUT�)�;b����k����[�Å�`v_�+�Gn�qPu��s�]�İ�D !�;����#Jd6���H��ٻ\([���4����b��U`��N����C�)�m;@��a��jǔH�i\w�x�Ď��a��,.��d�u������k}��X�櫠 �&�b켤3��d6t`8M�;0��-�s.���W
�ƛ*�a֏��Я8�M��䚕&�m\2���B�@b�t	�n�,q8�7umG����Ь|���]ȑuIr��Q�R1��˞�3ؓ�J}uy2
!�t*�h>35���9L⸫�s2�����1����r�T�[V
��V�1��ϴ���uy���I�оy�Vc��X3����tjW��*ˋ;lp:,�Q;����Zn��lR:(�<�Fy4�2iWS�}�R������.�l-�"V�q�e�=�Mqpn�����hak0����+^���&kR;�t
���Հ�>�J�n�fw�\�do�.�=�x��!�<��k��p��:e�Nxz�����*U}h�;�i�q���9 ;k�B��˳�n�t@�Ր�7�D�,9Ք^�:�hݛ�cH3�3��I���D�hu]�G,].��n�m]<���Cj�Ss��=�i�t�U�Ƶ��	-V���R\a�.\���Qr��tf�7v��Q��K�u���.�!�6�<XR��A��(�7Fe��RC\!=�-��s2���Q�,Rz���g���v�ݙ�h*C�����X6)�X���Ld����#[�$y�7�t���%��gE-���OS����p_c֋���\3Ss��ɣN�s�wk�p��c�����V��Y�>�f�2�*�������XG0�mfٱ�
Xp'�f��F��=c]m��ۚ�al��ւ�괅��T�e�3m2��Ep;���/5��\iL�1DCκ�{n�js�LM����ꅽ�����b!<�Z��tC�� ���*#s⻺�ǌ,#D3���8!��,�T��d�w)+� � m���|�s�C�����3*B��hA���<b��D�WB�j�jKmS�,j�N �o'Tp�4��:���C)8�ڻ喟v�7���p���q2��pA��#)shw���q���Q��`d���:2�[���Uc��d��3	u�H�6{�q}d��Aa�s\=�]n���	BBʰ�����qv�:VKClT��08l&�ڰ��n/�H�G��]p��oKv//~����|8�3PyU��p��}�z�Pt�oa����_k� ��*�p�����C�)p,U-a�E�gp7G����&��!�w${�z޺��j�a5ʴ�Rv	�[<y��B�Ԭ�����Pa�Z���`JU7��tM�t�9��J�Ӫ����)cq����v[�<F�j�Q%��n��^�
B���S��x�(��r�M��%c�=�n:�'�]��Sz'SrⱝP�P�92q�Π�sR�M�p��Ց���} ��̤����*����`���r$����q\�:�`9x�0����R����m��R��%���E�5�*�Γ2��K�v��/f��ƨS�p�G ��T����2�Tz�h휃�wrn}���FPc�)��˛R�ۗ8�3�����D��E��a�c����Š���V��A��*K�=���Y�����ۄ��j�FR׃u�]���p�Z�L<�����-沛�w;]n�Dte��[A�h��|���(�/nfC�Y�\�D�����Ƞ�u�^�땜z����Ȣ���2�P�룱p ��X�� iD;ΐ��-Pѫ��YƘ[��ߚۖ"�w�9���&L��/5�)��H�,�����٩��@ $���t�Fb��V��FLJV��VJ18�m��(���y+k���;��x�����ІַI��n�GzU1ǘ�0fV�;�E4�E|dX�������P���f0sy�c{�vV�8���s4�p�לi�/2S�⫬�()�P����3�V�/#?v7ԡ-����z�ì]m�q���d��.���]��� U%솹[\w�GE}���W<縜bj��+h:�8�;\�GW����z����)��|ďfc�֝�,_���7s��חhpZ�-����~w|�ٺ�'�0�HO�E^��V2�w�nM�j�>}�ET/I��-<���j��@g�"�X���Y{�(�oQ�֛+@�!�7��)���Xޭ��
�,&�6 >+��R�p܂�yB��;��\�Oz���
k�þnG}�]YX9���_dPג���hlfՍ�I�z5�+�}ڱ5r���@����㽕��	�S��wD%b�Z5-�{k�(䇟P������nS�X>ci�KiM����3���k�/l�낹Iǉ޽Iދ'�`H����Y�rl��tR�B��ըpI��v�ŵ�� pe�:L�X�?���S&ur��m�4"��+j�.�p��N��%�Ruu�eB��Ț6���4���`�2�l�@���f� F�Q�q���c!W����m૚���b��.k��>�]�ԝ�[���T%��K�����-�7y�[W�5��e�Ru�9.l<.KU��Y�3�Z�VZ4����m�5���K���S�)]äQ3}yjfCǐ���熫����sxd��k��X;��<M�O�ҳ�3n�	۰�bН�M���;s�n@6f&e�{V�B;�{͠��*��qq)��t-�� ���X,mun�����*�@��;�;{����`q6�+���B�TQ9���Iɐ��lf�`%̡`�or�}�*vݮ,����/��+Eɒot���3+n��횓٫|`�V ��T�|��}��4�uI���(5[���� �ӆ�j���e�]Y��������
�'���UAGw��C������S�|j��ݪ[{�h���K)aa��r��+mZy[��7y��fC!��j䇫�D72T��Y�=jE4:��X.���q�?G�\�5�ҩ�@�6mm��X�Χ\�w@i��VN�r]qF��gU�7ȝ;+�ĵJ K��}X�H9��gd<��f�6.�t�i�Q��!��L�\��D�`�9md�#��o[i�ҁ"�\
ι�t|q�T:5��t�i�6�)5��Y�q�5b�+�q�K�ǜ��)���S2���k�淡��[��d-��B�\�K }`��ɋ�Z�Ol�D���=f��S�Ssm�˹����\�/vɕ�e�%q����䶷E�y�Ř�G�SSSby7Kb�U؝p�!�j [m6��t��8�f�F�cy�������,Vl���3��S\Sj�ց�[uA»Gf��[��NZx�'�8���J���z�-��j[��Љy��6ܩh��Q9K����m,I���;I��3a�d���T&$r�YF��E�]a��N�;���'�g�5�f����%sAw�n����4��)ҒvU�o�n�0�N��'��{M���LZ�dܗ���)����-��0oA���xwx̳��)�C�љc��]o>#�Y&��F���e�0���e���ni�<��l�am󙝼n��U��S7�#}a0��f��5�ա�H���Ͳ!0-����ea]�Ӣ�������Ʉ����Wۻ�L-MھJU��-��\�l5m@�g`궧	�㛥����5X>-������Ż˖m�wXT�0�A
�h_�u)2,:�d���.��A��>1��G������l.�k���
�:B��,���X%�2t�mf���@��	?�oD�MX�ObD7b�9�~��l!(UMUr�e�P�b���[��:�ͨb[U��SM'N�82�/' j��t��#�K����-�*��8(���jʡ,c�l��8Ðԇ2�t��ul�F���0�W]��{͕���I	$�!	!$�O�  BqBB$�$$��r! �^�7�v�L�s��:g3T�kn��*�m�ʸG*ڻ7�\k�B�.n`�`ꔆe�t-X�E�Z��,�n%v���Z�Դ�-UrZ�1A��fYN���#D�Ya�%ʑ l9�vj9�kc�M@CA�3�rʵ���2]�h���Ԫ�?���+���AIXxn���[uj�T�Kt�
}(k��*Te�0RE���A�:��r�J��{x����5W&���&E��%G��k�����I8A���Њ8��Z`�:�؜��eggL53l<@zm&)��R7\ I �^d$�i�B�#�P��:;m��4����!�2��Q�G��mb��O�E�a��{Ke�!]j������d��s���=[:!�=:.q���O	[4gpK{�8a��̍c;泣ŋ/0wF�6��t����B�\�����D��q�d�Wc>i
̳Uv%PRyQ��N�!�i.GU�͢o�D!D�G�����i�
G����
�f"���p(2u��'Q��P˴�X6��o��W,]���R���uV���a͋My�i��S�+e�@1U1�P�G.��fjuU�������0Tw*���*gΜ��ͳ�v�� ��lD���AWJػ��}��:T��J��<Xt�ib���M�L:�2�B���܉�{B�Q`Ѐ�e��ܸ��a��ܥ@�;�F�f����"a�҄TpV#
��k(�1�mGZ�#��*tE�)�{u-Y$�6�ƅR%4B���g[������U���Zb�;إ,����8 TuNF�o)-^;�B�"�&^�|��3d�n��8��d����e��/��%'^nWI��n��l`�z��o~�r��
p�yR�\1I��;i0�� 9T$`���/�����!��{�Xe�ffe�U���gU�]-[k
۵��C��$i�\����=���f�xmc_i�F��4�7ց�LA:�nv��p.Ê��-��Uil'�m��$+tK�)��q��"�x�a�����2�5'�Ä�D0��Ś�IB�U��q������{�����X���n�Y*����Vi�l���Eya�5H:�6P�TE^��[nz�ӈ��K�����l!SA?��=�C#��8�t���#�j��ARD;�HFݎ�����U��_��u�4�q�����5�s�D�_Y�y<�ͽ��A#G+��!1|��:��L�A�SU�����_�m�+;��a�(ٌH��Tc �f�k��駞N*TB�<I�)
˱�nf5�0%�26�#M�a�����A���SV_1�/���̌q=k�яp���|���+%�>��GS�����(x¢wgے���'��\0�<Cܷޅ}=�+��^<kPO*��@�����y}\��{q��4�2!ԏ�T6�bj�[yj�4�)<�E)P��tb�UN4bW�����g�3��G��	o۴n��]��E��b�N{=���~���z�7���#�G�F+����>���T�ݝݮUآM^n�HX��E�ee�/���]�����|�]b\-�ʀG� ����
�n2:��G>W�2�'n��.6��R��Ũʝ�le�K���f���� �������@Q(/��x����0�1�n��H��en��C�~i������/v_ՄP��۴��$�M����~�=��`C�b��`x҇4�<R��HU�N���ڈ	�-Q��?ojb^�"���<�s��'�g_�m1��p�^�;|^�;�F_/���3X�I��8%1��=�G�w&�3䄶AI�=Fj��=�%�+����őc۾Sj����N�H��-��/#��O���,�~��UGy0�k���g�������B�����я^�|��\��^y�D��Y2�m8��]��A-��[��L�I`7��Sr��h#پ��n�_<�t�7f!lmy�d�Q�O�xu��}� ��h�+<�'k�N0>�6@��W�W�3&�*!���>��N[��7I_�=RQ�}]j*,�[z�N��8���)���.��7�C4d��Yb
�+� ,�AÉ����й},��qx��_a���w���5S��3��5�Z����4��W��ON��B�=��v�Su���������]�:�}�js��:1}��d��5dh˔L��nv�#Z��}Q�t��|�·���́Ն���p��h�gw=����D�9B�A�w~qՎ�zZ|��ށ�pec!^B��6��Y�S9_�{8\:�A��UW�'֬u/v���pQñh9k�~�/B��c���ƴm��7��'vU5�y���Wܡ$�P&i�*������.{2�"��\91X��F�Q�ٝi�S&R;���*k��7���M
�>�C{�"`�,�Qb�[�m_��z�'��7�8r���D��b?i���=L&�_Ϸ�La��+�O^�S�zuj'K�b�3^ˮ�����Ѻ����X��U��Z���u雎-d�H��)�p!��;��#NR����(]Mܣ�����0X���;n�<�vq�Ux##*�+X"D$QQ�PcDF�}u��{\���x8��x_d�~�|E1I����[IP�Z���=
k�W&f寽ذNf�:��(8O|��e+(|�^]ƫ{���]�=}���v���!��+���]%�d|>�o��KI�Vy��E���q��2���hvb\Qt`̗���K'o�6�z���G����wzOp@Co�J�6-̧Z;Y5�eߜ[h۟g�I�/�kΊ���+.I�n}��
y�?i�X=�{�����E�*_����U,�M&�FaSՕ\��k���%FB������(�\PW��U��Y�ٵi���X�1�X�k+����8�5����Y}�z�z�PL� 7�%
� y�� h�e�1$C��'dl�S����KwL�F�'4g�Wh�e�WD]��:c���H�2t�J	����'��vZ����������9��C=�T���-AkB�,= �Q��pV�;
6�}G;j#6�!���~��T��Y[�O2�����2*,d��������ϝ��3y�I@H$Hk��7�_�F�}�1����P}�Ə?=M���;��u�G��?[7��wZ�����{0%e�#Qev�u}�v���ﱪ�o�t�n��*'c>���wƫB��{u�©���V��2uQ��e�{�[�4�n�3�9�]N��u�q���eU*M��5��M��KD5T��Td3FW1b e������Y�{��.�y$�IV}f�!iv��G���[�FU����`�m���Y�Ⱦ�Vrm��n��;ar����;=��'���V�����NB�M��e�йW΋-�P,�ID�Ơm�}�M��ֆe�G]҅:NȖH΁�)q����r ��k�K���Xa��"v�/k�OO�¶{i�����m�t�}o>���u��B��o��U%����6�0���EK�J�ڒ�Ni;;�=��xv��T[Q�d}we�.�0�a��P�B��������1zw���� d+�dƹc�/�mĽ\��Uϲ��ۆv��v�%H�/7��ԝq�|��sif��~�ۏ��﯍y6����S�߽w�t�P�WޭY��� Y��s)�gu��)u���P"X����}���ש޽��;Tc�S��;,u��ܕ+;�P0�%�u�D�"Ԁ�J"�!��GO�'ξ�����������.q�.���#T�m/#V�Zc*���B�f��R�~�}��G<��;�dC0:,߯RV	��f��K���:�ԛ/dh�n����[�sr���A`(�{0f��5�e�F���&+n�bfђټ,܋i9���Z�(��c��{�ȕ�Y�W0��F�/^-��^��6c�v��X���'����ݻ���x����sp�H��"(�p�r���w�
���T���\Q���j��nTl�e���Eh>���V+.�x%xB�Z2y����>�+w0]���`���������ל}�)kzp����	p�z��ޓvWg���t�n���p�p��o�C�A���tf?��%p���wQ��9T)z�ŕ��m���W�Q}��QE,b���d�)"H���$D[��í�a�H�"e7X/���ۤ�:��i��&� `���=�#��z����U:�'��ES�N/gOs����ȝ�gk3�B�&*���y�3!VOe��c��9�^�ޭ>������
�VO����h��<��J�����+���^��j�8��E��͙�LG<2Ȼ��3T��9>AĠ�>��+9�s����ָ4?��}�����l��]c39�Fb�=y�^ӣ�je=��s�Φ��)Q�:��4*ne�ɹ?�jJ��=��9o�2�^�_��_�_.}� �2{t�lV�Sט�����Q��V��g���2˴+�fesӴ�H������{��v�㲔��<�}>I�Nmw��y�쁸�$�	�c4������F� ���>h����l���P�Pk$WƔ�8��EH���z>kvx]%��X�<�ιȔD����9On�0PET���E"EH�PE��"��_�fg�����teυ���fϾk-v�|��k��a�1q}R���y�s�6|9]��`#T�����~�.Z�	���>ke��$�[���)��n~��b�o���"6�"���d�/�Rh����Vo��WB�G������@ש囓�'�*�c��2��A(�)^�뒁�����x��x�c~�ȗ��׫�g�F �T�)�Tb#���Ab1U����t������ֈ�d�ǻ]F��lD�<���Jo5�b"�K��%�����	@�=b�^��%�����Ίӳ�nxq3�0^Y�e���O16;����GvV׳7}�7�i�v���Y�S�I�x<�^uV��zE��J1AD�PڗVE�-�%�����.�s�J����a�}���5�A���5��X�KtDU����1�C�,�QSK>�A� N:2v4�j r}X/�ì�cE���>��ȃd1P��7�͹����,F1��j��v\�3 �l�~o[�,?�x��K#K�"���o�����=Q��=��{�n�{�݁=o��׉N����g��:i��α꯫�\���;���0l�̍�r���NR�\Q�Z�#I�wJ�fG7����X�/o���-V��qx(u�+Ҭ�S��+�s����| �d�Ĉ�����﷞�����>6}G�)�;3�OA����+�;�<��s�M� c$XI^���Yi�r�2��8�U�\�1�wT]�Zb�Ht�N<���q���2tٕ$�ƥ��qI&�mnUic7�LCSlX�e���BSTY��$J�t�X� ���k��a�ScTf����2f,�}�D�S�p U�#�eб�r|x���޴PNCq��완:�Q�x2�V�yr�ts��T�(On�Q��ϟA�uu�
��{:��HγJ1��E�Z��^B���
K�i�Iy��>C0������o����/���ѷ���(�dW~ΛK4��Cȃ�(7���qz4""���@����
,�g�_k����\I<���}�v�l���ǗW�(��"`A)�LR�&77��%^AOuÜ<���w��]��/u*�w�������t8�+�IJ+�%.�$�cw^�����N���C�Y�y��hY�[.g/�:]-����ܞ�c�{}Y�G�j��[lzI����a�"0��F#(р�|l�f�;0�1`(�QG�w�����}[Y;k9�\I!�@�fu����ǹ�i��)��v�aj<0��쎯�4�@w��ܒ:��д�O�G�G5��mT��=�}��G�n���m�Ǘ�:t�W��s���K�dP���Y��S�]�y��ɳ.P����iR�>�/�"��ə]���k�[������8�㷙s���v����a6ݗ]O�Cz��N�V��!���r	������C.�v��X�{��۫����^uQ��w=�61���&PDE X
��X*M�t�^}�_ښ]���>��9��OV  �*^��3�*uWӶ��>Z���.���{��Ǽ�-�H������3���k F���'�qj��:�v_/)��՞�}�|3�g�^��9d��cȸ���ZeeS�#��ꃍ�����2}4�u}����(Է������}#��Q���hڏS�g6Z��{��T���~�I
�s�y�[���߸^sU�w;���vf��0P�  H��������n�κ�������+5|O�`�|V/d�kk|�&���%��./n
�;�;^��j�c�	�	1�d��a��h	d&�C|���X锯9���8�_<�^[���ẻua���A~y�ҋ�U�/�.�䬓��-��e��tֲ�ә�9��#��0_�z�U�hṱm���	R̷.�y�q2������F��wi�m�86�》Z������er�|F�Jc
�=��#���izs!U%�7Y���)f���;��j�(Рp��7��nq�8�[e֜�m7��Z'���6�M����ɾͫ.��Щ]>G�d`��);��hi��c�e(���P<�4�	�R�QY㷆�ZCְ,����8���x�lj.��6�zI��2e�;��,���$�)�X)^���Ṃ��|�o4*F^.|y�����^t/�^�w��xV@��i����O���5����=���Kd���8���IT�XRX��FLJYꧯl�X�-��I��;�\����d�w�]6�>}�ᾪ�R��U�6%� �E_D6A����~$ilER�M�Q��;����7��m���T���G'S���% ���N]�9.:(��W���@홄Ӧ�_u0�.n�3X��f�] ,֣{�`�d�˂g��4ƊHi:&=��ŏ��2�K�zad|jd�m�l���т��,� >7�W"c��C@3��
�4|:�.�����Z�E"(N*��;Iu��z������oq�Y֖�:��J5}���|�2��w}1��J�u7�J���
��o,�:�o�훖�-��h�+��f�����ť
��ۺnD)���<��;,u�J8��M�+���i�5�zuq�C����Pd������\ͼ5mkwW� ������)�P��1r�j�䈴�*V���Q<4]Ohf���Z���ȳ����)��J�4s��V�V��!E��p53���V1p�B,��d	2���J�z���������ͬ�F�t[m)x�W�^b���V�.12�q��,�V��YWXC��S��N}f�4wR��q^�컆�(��z�-;� <�G/�s�ՙ�~���g�V�h�2�=�;�9�@89����|ij�(��0k�{���ORI��-�\{Nm蠞���$�6خj��_ '·���m���%$�OJ����
ví�wSN��z:Y����à//	M법����gM=i�	1�0��R��JwZ���\�Fu���ꝉ7�(��:�C~�����q�U�pN�q�AHLWԹ�+ލ�Q=��}���hc��욟,�@B�$�oԏ��(rT)�َ�1���#L_<
��hLժu���N���%[G�Z�A��"��
�)�R�T�)E��F)%�+���w?'7^��(��b� D}륩��	9��Ւ�D���W���ڊ�����u���/+���0��E6ǘ�F�Z�j��(��u�,�([�Ρ��}�3U𷞍�
U���7KEs�T�bZu���ʿ��Mc׶R���G$���=)驥�@0�=ʊEψ2�q�mN3�ק��{=#>��2f��W(�5Y�s�9�68�����V	4���>0:��Q^��m-&X����օ.M�}�я��I �����EI�Ӻ_��9s��)[�������9-��ČL<�tb�=�s�j0w��j�:��RB����٢���͙����$�(�Rh(s��/<��.�4�Yw��w�����D�]� ��sF
�^q��1� A��R��u�usW���S��z����'v�2�w���(�^-�n��w���v�o~^��`Q�q�ӎ�!zeC�q��kq�<���#ԩ5�M�G�><e�Q�r]d�z}��b�H��H[�u֩���m��R"�Ȣ,��k�U�}�XU]VMv�kq�#K�`-���)6���}5��� �H("@E���?���/��V�S��:e�΋}@h"e\�ᾗ&	��~�����$2%L��hZGӼ�h�:�:0�
Z��򷪏�zM�x\3��z�k�YK��G�Fj貪5}9퉉�����%9�}����#���RhF;^D�F.��ެ�v��U�:{K>� ���0���q��U�j�}�j�q{o���ۏ�ac�)� !�ʄQ7��}dO ��cri
�N�&]���9�E�]-0�ID�ǦI��Q������;�1�}��к��U��1�p���֒�hdX�ґ��Y��ߢ	6�K�/SP�_�&�J}�GB�7�r�[��o�V��W�SW�F�� 0_��n9���~���n_[�u��>sP$� X�V��y�uUM�IE�V�kv���;M�d����%
��4M����ĕ�}W�a�a���`�tFЬ��hͽ���v�1R2�̂![!��0V�H������Y2�5��^��.�0z�w]Od�s��s��k𝛃�D�e`/d�VU�J@�#H�{�,����}Nx�be�IEt�3��{1�H��4iZ������_7����_�sΑX(($b�1Q@H(�E�QA�#����_��4k��|���?{]5���h�w��Un�¥R�������UH-U ��i*J��Ϫ���8��D�]���396�S�zGz�*����Uv�T�%~k���R߭�E�r��ll�"l�hߪtF���>�ɗ��ܳ3�}$ong�)�ZO7?!"�����_�l�e]����}�O5W�4�����g�{�	�������R��	�?2��u
@�o�C��+�S	�|ɿ�r�O y&���0>?^��֍����_��;��߹W�0������IV�y��$>d�d4��'<�ϐ�8é�U@�B���N2B�V��̜M2J��&!��L-�/.`P����_s_�	�!��eCO��� 4��>���l�1$1���i��$��~����5�� C�8XO!-?0|T�\�a4Ͱ5� y';A�a'w���_����׀��Al��w��II	��$�M������~CwS͠S�Z�h3�036�,�6��1 �O0����JC䐮:�]��E[P�#�R��/.BR�V�0Rp52��BN!�P|��3(
N2C\�7t�oU ��C�^�P�KHu	��@����i$�!�;��9��|�!-�Y4���f�Q2}���5�ֵ�/�����x q�}P!�'�R�����y
��,��y �0���HHZ����j��E���Xi&$1�|�HKJa7�I���<�?i 0/�j���<�5��~�ٵ�n;�@)�(=ߞW�Z�n�;���炈�%<���tY�%Aۇ����z�<���_y���s�I��1J@8��s�-�%��yA>a�Hi�'��|�C�'�P<��д��
�0d��	��$�B[+T�}ܒ$�BÜ���]D�EEUUR#0�Ub'+������}<��Ho�y��u��@��!'weͤ�e$>d+\���z�c$�BBc�h�[$�C]�
���d��A6���_5̺����|�@|��H?�'�J��q��$��q�b|��@���HR�T&�!� ���� �����m�����r�H��W�Z����5��j���M'X2r�a'�!  }�u�-��a7��L4�m�i������HHm �HRP��+�	�3T�]d�8��i�|�i�}�������o��^�Ky�L0޿�� P7��:�O�����m	��RI&���(��W��@�L���n���4����Ϲ����L�d�`Ra��?!䁌@���0dך0��i�E R	Z�'�~�t Q&2~C�)���Xځ����HM�����ʗ�ZE\ N��x��Im�
�Ʈ��f�~�-����
t����XO�C+�O�	Ą��n�p4�y��*�qS���$�@�C�!=��䓈��kue*kZ���oe_���y������j�]��9f�*���kG󮝙c]�bf�F��&_�}W������r�+|/6�����ۈ>�Q�yg�.<s���׳�W���Ïv�̎K���[%'�����'b��*�VmV�q:V�m�d|���Y����a�H3�����̧���1�A��
A"
*$QQ ��E��o��㗽��2t�D�ѫЎ0Rg���t�վ�t��Ǝ�t}E��ٌ��w���;W����>�Z�Z		�?s%��3�]�,��',���:+�lК˘�6_�� �^�ֻ
�@I��̡%@&��RO=��nLpCv<���?�w���E�+Jo����~V9ȻQc~ 1��Wl�?���"��7���z\c��Gc���]�h�b��?ws��1����nj��]<�����'4`��� �ʬ]�Djqm \T�7R(�8�0��̩��;Փ�.���]�ֳW�����/U�Ԅ���# ���� y�u�vxs��۠ʯ������n�p�x@XE�\�H��}��ɑg'��f�2t���aJ3��}��Ĥ�eL3��ݩ�x&M����BO{Tǜ���^7�����+7}5�@�@����#ݡ ��z�BX�RxA��������*ġ�g��Xw]MK_vrzW�rS2����6��ї�����;�;�6�:魵�U@�e������ �A",E�������*f)���%ڻ귪�=�˴�	��#j&�^1���a�Q4�
`@P�b��ł
1BA((

H";�k��{Y�W����}���@��%e>�;[�˦/�"9�Sx�S�Q�+��H��o!6��N��ͻLUᩱ<��)B����H�Ͻ�>�܅7�r�ٵbb�mە�
���~&C\|^W���ۀ÷64L6=��%�k�"=��}V�Wy/Ê8h�6d��,QW��(�a�n$\3��@�l��/�X�d��a!����"T0��zM"�	��=.b�N�]�M�a��Ł�|m����D}��'\͟u�Z�{����/��g��h���&>��>�O��hW�f����׌`s�9f_�&��=��EJW{P��{�r��A�-�	���#�:k��ԢD��7 ����J��{�Ѭ�T��:c�iOx����;�=��G�t������ot�*�N��5��g��]��$�u���G�p!���k�B�t������ҫiPJ<��M��8�2�5dֽN��-Fر��Sy�X�ލ���+�]�+��) <Bs�_�QU�E�U""��B)���W���x��o5��~�_\y�7T��/������TxB'�X��շ^[_���Έ�4����WZ�W��uԒk:�>���Uv���-F�@W�:�X�א�Z-��`�'
��o`]X}���Sl�o;k���@[Wع.Ab���
a�eؐ��d2}���Ct�]9��G/�L����&4�P��9��G $�c%��vM����JBL����,�h��2�����BĹ��<���T���.'}`H���.��C�ea5~K�W��]���>����@Oe�9V:O�Y�N�ʬ�^�)���:����^\��a���><ihs�C�����c�|� ��<+E��F��gA]��Ԣ}�L��bo�0G;P0S��$��A�ffe�{���޽R����r������
e7]����#��&�ƝL݊�S::�p���=G=y���Unj�$�JEN���~6��X���Lp��I�#�� 1a��Kc󬞮�e�?��<�0)��� >����'T�Ri[��\��x57-�C��[���)t�Q�ք�<'�n!ҖlPV:�W��mzf&b���>�4OЈ�"AF ��U�o�y��k�V�خw[�;{�w����s[ޭ3��m�d��0Q�����ê9�G�X��v:��
S�y��z���Dߢ鷡��gya0O]{�{v=CD�y5NH���QV�r�ܹ���f+�� ^ծƔ����x����4�  �czEƫtQݬ�f�E�Hw9��8\��t��0Qh*�nɋ%9����\M଎F��ޚo�3�8=��!�g.&���z ��G�v|(m�N��M�~��U�a⒛Y� f�nZ�����>���+�]��K�7�|B���wQ�'��>�)2�����(붿~T&����%m�����U�V�������0�45T2
B�!(�j
��BP#��yo���s���"�/^=�N������4��΋ {��0��7�r�W�l���������6 �ޟI�9�UF�0uէ=�=�n<���z�F;~y�z��R�������r��}��G�dj�=i�7���I�|9f�xC>���������㖆��3��.mo�r�T�.I��{�*����P�9�.$�˭������X����.7���⾹qx[�7&��z/��g��qԁ5�A��������<����i�R����yܿ����*�`����V{��WY���t}֔�FƎ��p^��`ݡg����,�Bݹ2�.Wc�lqNȀ0�;R-���l~����kAB�bT�vg����
Z y4�M���1Sn	����Mh̾�@RE�E���B���)�Dٵ{��.wQ��Jt�=���I�G�$k}g�`�u���ԉ�I�	^\϶�I�2�t/��N�rQI�������ǜ�!uEϫ�({��l*�f�թ8F�rY"<G<�¯�(�.��C=;�=�U�����Zox/x*_}����#��K9��!?a�I��S�J���#@eOPs�!�ۼ�Y�d��{�f���wd_l�,J��1STo���`�{�#�Ƀ��3oG�|����� P�FG���:� ��16>b���~�"+��P�oo���T�8�����r��������g3�3M�;�G�t
�}L?y)C���SB+��վ;��Pg2D���,/�as6#s�E��^�q���7\�_/ڗ��h�C�6t���{�
b
*��,��,b�
8��C߯��|��ӵ��3"�(��B28�;*ǦTt�A��Sx�<�����9^�M�'�LV\L57=\����v������������}<�yCثC��ܑ� 9�M�>�#�bsk�*�o�'QaY�J�{g��0u���8�������!ӯ����w�Wn����@"�@��}����㑇7{�t^V-�V;6�6��˸�U�|�)�/qM���W��5�ū赴W���@4&e�1��ԪfȐ��,}NDeՌRB����Wt�J�.�d2�������@��`#�櫟��oW��Y�s;�繝p��;���3��A�92�B�m���4dp��fyS̐ze�;���xf;�xꢗv�̕Z�m��cك��?��3�L^��s��3a<l�H3 �W�L��}�͕���b���$N�Ì���o�QDޭ�2F�vne�����[B��p����`R���+���r`�g[�r� 3m�-��"�?�| G�A�A Py�v�^���^W��!�����1��o��O����5�R{�%�jv4�N�/	`�cG�o�"�v���w{���#3���S,�9�T{eiry�w���/���F/ӣc.�W�q�țQ���ďwv�M������@�+����Ol.���K�6�g	�?��.�74�ך=K�j�[����|#�Vj��{�֊ҹ(۵n������7s ��wbx��`(�֩Yf�(��w� 
xC�W�c�gf��w�ӴN.k;],��ݲ3Oj��{&5��^�q�h����-��1�GEB��F���iJ��=E�����Eq3���]h�h��0$G�Ӵ`C���{���N�M˿�������R�qA	A�W^�M)q�H�����jE��r�sN�vJT^0�9ݬs�f^�	�v��Q×ׇ3j���]ӧ
�y�.��By'��KzUMÝ�$/�����3Q�[\��5Wrѡ(U��w�V��b����T�]]�]��KW�_!8X�4�K�Ơ�5��d�P͠�(&����Zf�Ɏn��}��0��c�ָ�b�Vކ���_a�pl�j���x'�J�0c�x�u�5��B��Pt��h��CB64��E%�l}H�%��Du��H Y���D�Tv��rfs�x)Ԝږ��b��B�:��N�l�� ��J��I}�(4*�uO�:�T�U��˅-�C��:�]7KB���v�cWT^�?h��c�[.Q�n�e�q�p�a-2sT�����[Uz��	����B�{F��S/�T_!S�Z��4�/)Y��6e�g��fk�W�u��E��@�9��~�ٷ�*��cgD�(�"��+�ʪ��n@u��c]�e5�%������R�P�"�Z�e�t�{��9uє�[��Y�m��FД֌n0E��1�:2�piպi�Ej�Qz�����)i@�ee�KV֎��L9
[%�b�׬j�j:ݬ��_kX�[�Xճ*q�ƶ�,#�y��Qf�l�D�B��O��E�_n
�J;\Gh�@�q�5UW�e�M�T��'e*u`��[,n&���W�' ުyj��5��$�Nݒ%u��0%�+Q�1�L#qu�x� �H�G�*�l ��s3+RFۧ�IYo@2�F��.mq��;�R�j�sUlq3�ob2�S�R�F��$�U�\�{�*W]]ӻ=@X�ى#V)j��,�X������qq��7�����u�u��V�k.�%�2>`L,wmr�h���-h̆��nT��IeN��;XVL���&HL��%My�z�(�ڱ��p��+��H� ER��Ռ�ə�m�ՙ��IȻ��$�UB���I�F�������y�R����XN�:��u�K�]H��l�^��P{�W�W 8McL��ƭ*��TuV�ԅ��D_.oU�S%����/�Y*�;@��*�D�Vk��I���#j�7�6qM��I���2���x�0������<���F��M���8�1����l塃dY"[aj�����X�LS	ף^	�s��FK�%	1R�Za��h��յ��0�ֆ�dc:J�=��l�,X%�#|#t�dž\��o�Z͢��iL�����3�'i�(z��sH��T�����T��v\#ŀ_ q�9�ŖN�yrV=�K�TF�B�vT�\U�k��z7B�Æ
�e��7��L�f�66e\���o/1�S9\8$��X��M��"�!A}"8ZM��?s�������]$T.�L�{Z�� �;9�z�*��{��U1�56؁�UK���)���޸"&����V�˭UG���wX+CD����'�_�i�	��\`��UYV*��
��L��9�;pζ�
���1!�;����Wz�ngO����:��F�-��{��:�[�üjy�g�	X���dg:�����ꭁr�_NҘp"�b�%H���}��f�pE�k|�uV�>�z~���-�4�ۗY3�K�4!��݀��UB˔��.v⣊�=��t�*�D}��<��ۙe�ܒc��x�#i�$����ꉷZ*� #�O.�}T��w��m���ιVXu�����^<_Hțbg�k�ϭvr�@���U�pO$$���d��?w���r��>uY�s}~�E�}�k_o�qdP`��0A � fmPfY[u�EB��]ώ�iچ������F�X�#��t�v��N=��v�|6cUa�f?�U���1@�74�Pq�=����U�Rj!%�-�c4~����f�|�i���>z���鷽�τ�%�S4r0[s}k��<"t�����Z{չѝ�<O��ˈ��	F�l��:u��V�U2���z�� ��wc(gg�{IN��تZ������|
0A"��
���EX�1T��*�V
�#UB��EX���bE4
����TD��Q����  (�Y�3@o�c����.Q�:�Tͧ���h��N�_&JѶ�f�n��;ĭ��;��������^\�pՉq�"�N�*+�oO۾�!җ�י�'��#�7P2j��]7��dNM'"�r�]w��� ��6����ԯ0�Yw�.L�/�/uh$p� ۆ��������$u�~\H�O��K�����������H��w�(����5Q�o�Gk�;?�k�yXg@��%öBV��5�RP�S๕m!��DF5�����`���`���IF
�`*���}����k������χa9eζ���*B|bk�1�y�i�=��̪�w:��9���m���&��$mT��ЂT�:э&���燻>�yu~.�3��J��OH��O.��r�$��<�GU���}c�T��s�(��R�^� f�6	��q2[�u~:�@F^�-�9�o�i�E�5�:r&^/�N��K~F���^@�w���n{Y����n���Nx��s�|ݵ��0 �A"?}�D(�7㸔�F�s���?[i�v���9��q5��5�V{|\v2q�=Y~��OaK�:H�k���̭��9�ڼ.i���ҋ�b;�p�<��.�Kc��J��4���Z$%+�Ho6vN���H���(,�_�j���	w=W�;7�^��{��g�1J�rf�2����W�5�%����(����g���(�s�~RʐC����	�KO�M����Qqy�=Q|]u`�^''B���s}��@�#Ⱥ]9��Yi��_t{~�EQbF �H�$H�Tm��Ww�k/=�w���DD��D�eY-L󨜌���9]?��Q|�)��X�U0��꣧��V˦=��_,�ԝ7&;\�@��$�yѩ6������i���`9}��R&����gm`���3�{�M��^��}^��u2�g��U*�V.W�x>�~�EkF�D��1Fg+�]y� ���>��+|T��^��e���
<��p�����=� ��~ÅQu��̯�f�+��ܵV+��8�l�e¿^�$�dmK�@�}���P��N��Uѩ�Sf$�6߈���i��}�'H�rv�2���t�莚��`�Z��%�����e��ԕU�}�߽B�|w(���I�UNU���^%[�����õ�ry�릠n���rS'���"�؃{HM�����W�������z��ښ�O@��5O���������?c�*��}�CsM��FU��6u2q����t1y@�Ӽ� �=Ӿ��w�ݫ.D���On���Ƈ�_�Y���q�P�7�9�%uW�	���)�����Q;~T*�_{�����`C���f��l*��>`��}U~Kl����8��%
�*,X1�d>�>��l5����}){[�����w/�Ǻn-�5���G��3�>�8���Gtb``���U�}u"ta[4�����?;���D�O�UGc�;��گ}�Z2���>�A�1*�!L0�CL�8�HU&a��w&I���U�+�]f�b�χ��F�R���Su�A1��i�s� �4���3���,���=��~�z���P�1EF2 >   y}��dw��fhq��}�q����U���sG����������#�0�}����."�4l�g�䖙�]���Izn�������4bR�U�U�> |�QT�e����nI6��]��ꚰ�F��ڍHb��s��q�f�C� �����6\:��\2MF EN�E`�˫l4U�޴M,IV5�Ӿ�,Qd���zAZ����o���-r��@��[V~v`�����RH�H���xb��!s����4%��Ă��Hh���<� �?� >
D2�C��{�"Q���눈����Ψ7[>:��ٗ*���]8�;匎�#AZL/���*>��x�_TFmb��c�q��Bt8�(B��z�>�DTY���L껛���ڄ!�� �zbQ�ѱ�!A��*QA2s�z�-��k~��ʝ$��[m�T@c"��""�)U��2�{����9���GX�.^�j��y��zUhq|�;P�"��~ �NX�b �R������g*�?��ҿ%Z�5��B��A	���4̂#odHZд�"(l�i���>�TJF�8��eN� ���{N���&C�Ȩ��^_rpҡ�2W�Z���t�C|�b@�)���le��a�W
���ȠDl�:�����c[DՉ�@���Eᾩ���=D
mH��k�����w�N�J�����1��7�3d"H/ݰJ����񆎆����__��+���$�!��Ǘ@����~�@N�˟��_;����D�q�B+̸�2T�i>+���)�YXq�WF,4t5Ӣx����!Y�d@����/��B�6����|:�E)��&稺,�5ԉ��m)� P!	���B�4"���ŷW5�i��S�(�¡v\��u��t{{.��]o+�|&���M	�JF0cڤPX��X�b�F,&��"�n�o�^���,ͮ�uu��y�\�;�����5�r>&�&�=��;U!�t�L���F�/4���$VP �XC�������(0D�h�z�E���0��'�P��i��0F�p|��W���J�rb\E��e�0cǸ�j���يY�R�S�c#�^�qQa�R��ą��ğQjAX��,�PY #�=�_f|4�:��Y如�[	*�j�H�hq��}��ݡO4�c[�;^,����xp�7�8<���C��hh��!�(H��o�:(!�Ԙ`��B�Ak����[��B��Oӫڰ�"C��?Y�o��������L��������������Q~E�)k��W:/�� �������e��F�B��`^���Ȣ�x�B@�;��*Xm9!��,(��<E�W�#����(���ߪ��c�T�͎`�m���s�Q2����Xl���R���H�u�8,[��qf�	�BoS5��*�ё��(B<c�I�����(�#Z���uK�F�P���F���1aY��>�h�"A p-W/)��"���ER�U0&lA��=���G(5����Pv
XP�C�"1%	oJ�raDY��c�W��xTn艜�Ԧ�M�;L��"�:�;�ߴ��&q��$�R{��߉��A@�&A3-�T]l���.|l�X] 3*���ڶ:�S�[%�a����}���'yita�⮜3L�]r��4��O��(T1-�9w��Y'j�2�X���¹D͞JWt[x���ޫg��	�4��H~k��ZQ����ܱ(8�)Ή�m2ñR�Y9\�C�t����<�ZcA#�pG8"�A��Yv����g8Ͼ F���� "���O6����L~����_��?�v��"�2(��
����o��_V�t~�y�����P>J�3�ᑃ�!��N��͖�F�LF[; �(Þ���5���.1a���;43��a�}J��O�z(�a����)����Bu*f9�΂��{���d��ɮ��%'4=;�v��J
w��-���O�uԃ��5�O��0<_jb�Q��T]���H��'���5G�V���6SG	�˨�{��a#1 Ԙ���&9�$���o�%EE����,sɞǐ�ʇCȅ �#Z�(h�d]x���Ӆ���#u�DP6Q:�u��F���W_�)�b��ET@����a�@�j�؄YR��b�G���W/Q�B�y��<4Vc�1�[�-/�q���0���bMGZg�4��F�����@�e![��C����ZįzgB�6���N����AA���E��˹C��o�+�>��%�X�~1Y?6��b���� �u!��
�&(�(O$B���0�P���b>�r`���? z����+������O��Tm�4♞���o_{��V��I{Z�7�&&v+tNZw�\�B��:Xq��zɫ��*Nf�l��ńv5�l)mzf��Z�#~�Z-�����܌�(8�n�d� Q��	��e	`�- ��1�=l�'�N�{�b�e0b����R#��Qb����֞o\�H_��"1�x"7�|�P��{���o,��"��ufpa�1�\Q�iQ��-��8��Y��9�E�#33 �`�C=/�.(`#{�;8�ă`�W�Y��s1��L!龻����o��|�##�;�N}�Tx�����R@�B���b¿�� �
���.�>��p���Db�cZ�gA�1�3���RݵF
(C/���ȂD(�Mq�� ���f�3�J�H�gUH�а�_�}� qZ�l�,�O?�~��d���LDn�-bV�D:�0�o�Yb�E�I��� ��|DYbz�n��ܽ�sY��n�V�A?�7P���.�K<�GŐ�;e¿yĸ��&ڒ��2��W/�?�(�E=�G
?j@�߯��A��^��Vh�A%�>Do�x?i�����	E*Q(�"��~�w��<ET?� �"�~-k�8"l?K@��]Z)�Y�V@�� �� @��`�!l�K����pЅ�0�V_:.��
B�Gis���z���?{{�JwhG�ڄ ߧ�i�UH ��侇Z9&A�-�Q�F�aj�*�&u�H��>������Պ�TS�Y]�m:[ϲW΀��P*Ȫ
�
�
AH)"!��0Aa�^�e�e���V\�m��+���.].YZ��,i�B-�H�̌�"6�Pˏv����r�mÝk����,+�dz��qR�&�A��pJ�����X��B)=u���w8��A]4K�=�NK�'�����a$���Y1D�l�J�2�D_�5R:�����o4��}�m�_W�w�@�[��L���l�VQ�E+�k�z��4Zly-�jY�<�߮`I�S6�ʚ����Q��S���f�\�+���a���ῬR_Nm��)���>tɕ$�C�^�q��M���"A���TP�(�Z��z��q/ք5��|��2�h��5r~5���fT^�����gusF;���d5E}g�M/NҲ�?�Y��	t�M�
堰A�\C7
g�m馾ƺ�8Ǭj��Nyx��LL.�<��h�bb42��W���H�Ċ+��~p;å��w�Y��#9G��Q���E�`�Q~��knfگn�B��������t�͆��9)@�[0�YZh!�ޅ	j��65�9?/ Ϻ~�GρG4!T��!�Y?�1�s���5�)��R_��f�兞;�)rJ��	��利��k�y�e�ы��=&5�i��"$�#A~���O����1�������ߩ=<=�ｑU+����w���$JDԖ0���0�&%<�Er��d<}*,�`�f��j�V�Li�`������Q�S�ͼk�=�(�^�ս�kq>D�w��ep�r����cT`�XF2�B[��.'k���^�>k{O��2?~��!1��G6��`����!��$QdR�!�	B������*�#�G/z�.P��3%/��ov� �Cb4�2�2��r��������f�Y���"�^�����ώ��",l��hu<�qKs��d(�z� �nz�������vd��������{R��_1쩆��(NU�<�m
�.TWJZ�w�s�Ћ�|���}9.�`�Ϡ��������1Uᣣ�¼`�?<�M����#L�;�FF�`�6.,�j�j::��)0���P)]�����Y���,MN�EI:z$�3'h�#����N��d^�Y=(�y�8Y�LyBeثٴ'�.��*U��AS,ֺ�a��#�}�0>��7���w �J�z1y���x�d�`>P��&l��wOTD���P�%�b�XvO�2r���Ԧ��v�Ϸ��23�iu�QV�!�s�瓬%=ۍ�(+�Ǻ{����6����r�	��xp"����{\/9�H�OŃe<�
#<۲��+�>,�^P�B��3_�Ϫ��+6�[��>(��Ա���Xc���S?�  j��H�C��*6�Ձ�H�&�2�umz+9<��"s�nT.����F�:d�h ��S}�C�f��{/vz�+쭴�b�;]�!j��a��V+sz�_��w��S��@0���T�z�G630��a�:<ӭ|~��4�H����������z����B(�>�����C�T��/=.� �̐�i�b�}Wh��w^�e4+AaDib��ӡe>��q4c&�eHo���]h� �s\�ʒ�=�j��gE�X���1�ֱf9�����Hw ���Lv�&�j���n䂇`���U�#Q�Sk0���Sݺx�t{���F�u��-Ѷ�T�����<�1��ک�H�afR���|h �i&yk>�W)d
*D7�ؖ�Zr86����Bu�ߺ��C�6�Oq��>JH���n���У���f�x��;).ףp!Yo��6��ԥ��̷u����� �@�M�{l�U��s��5Y����Be��!��K/�\m޼��,�8
���.R�ML\�X�6� �}KG2#�ݚy���V%�+}�9[�d��vm�Il03��Y:�6�+o����T%U- \1-PX9�A����m�x]����'��ץj�r���Re�yye�%d��ۢ��E$0�6�ˡ5�����}�~�N8��-�#�Q����L�%�<tw���պ9���e�o���^��x�*���m�S�BX�M�Z5�o�@�� c�k�7�Ϭ�w�6{Xֳ0�
Ce��@�Im^��^�$	��Gm���"�|Ƌ���WٌbT�+'��Q�u��k���5�q��\��6�ِc�k0zSز�I���Kd�����JuA�]#.�(� ��ËXflj��J���ӫ��.�`�#"�2�5�����c�=G���M�n�t4w����۽'h�FM�&�Yǃ�gtY�S���"�ݫ�A�yahM���+&T	fi<�N:���.�n�,ʰ ܴ�����H�>:9�T�*޵*gy�ݝ+%�Æ�͌b�(;�Z�.�q_��#b=���D�rK��m@�����^�)�w�����rT)V&+]B�zP�7�[�x���*3O�J�����ٚA3��)����_;Z��6���i�͎��˱<���b�)+��i�V��3:��l5��ga�ݞf�uq%`�ֹ�كG@Q� �eS<e��p�wd��=�_$��vMUx6�%v�(�#����&�e./N�$F�ۉ��h�����N�<���[\"���u&sD�j��}@�]*+�����r���B�{dŁp��D��X�:r���шnV��;���f�;����QҎ�����c�]d�!�j<2����`"+��F����Ş<ʳ�hYܛRNT�����#협����:�`�؏��@Fdо(V�N�`а�cQ�G�(j�4@;�wq���G���QT`����u�6GF~p
>4�ӱ
:s�W���!��.�������h��~��=�6�ۉ����
 �L�	�<q�
����BD:To���%��h��a�)a���)(A�o��G��dT0���a������dQ-�1 �7ǎ:a�ҵB���%2���k��a�A���݂�0�\��;�-dR�-��I�YA���C;�y����ٖ�FAh#��~�L9��R�昤�D�<~9�\,ߌ.Ͻ[�AR_�u���}&&� �8.� ���GڜG����Y��9��3Jy�\@�R#}��Vv�a8!��<�tV?4u�X?];��^q>mD�iV#��#ϝ���	��w�{?r����IB��(Ĉ�+[���u��7R���(ު�����q��=�兀R+"HEFI ���*��n�}!5[G�7���N�B��>,����eDEJ[��s���p�x���J7LE�L��x��`�'�4:������g�®2�\ޅڀ!qC4��t�=D5��?�;�j�5���c�C�-�_}_t�׵���9�|X�ʖ�'�P�t��T����x�p�އX0�l%�|���Ŭ���y��P�w�H�Q�E�e�"X?msM3V_'�����!����r�����0$�q�/%K̇��1L�Y��V�c��j,H ��Q0������� Ne�z�,A�G�Xf��O�s����@��c�jwJ�lᙍz��YČ�L�&u��Qç�Q�~�0H'J6+p��X��,rK���{ tQ4S�3�5���w�L.�F�QB�P����Q�h�IHɳ|��r����u�+�V��<�۵��r�`��W@���/2��-��US�`C����D\MwuC�|�N:��B��ޞ|;��6����(p�b4�0�<�,����L�?z��9�v��X�+jV.;��8W��߶~�;�\�V����t㶇� 4�k�~Q�b����r�s7��4��4�YM�;{2 `�%P"�����cilR����t��9��O-qG��x"g�"�a�,��^�:��&�`{�-�ԡ	��b
+LUhO�F��[��G����
�?$�*O�z4�k�׸Uesh%��ˈ��1F+E I!, !��1��\�����Rw�H�6���OzGɖci�.z�Ԃ�D1|͕��3ư�1�H�2���7��F��P��(�!��}����L}�	�	cs�D��H�-���"�Ʈ�}����Z��۵��ҽK�cW�8~|#�S����F6\2?�`
�4v�7j��v���Qb��
�ĝZ%R!��mQSAwO�G�3#��� s�,;��sAԷ��l�7E�|T���]ՔjC;��,l|���׿�~���{�[���������T^I�
e]��gj���'#1F�.R����jY���d&����T8G����ɀ=�8�W�%@��<��ҏ����~�kVLz�6Y�W'�3���l{�-p]��h��	G�G;>?�� �L��<)O�C�S��$���]2�P� ������B�k�3��35����ы�1�~D� �V��G*�q���'�5�4��0�V6��%��rLij/�j�R`��;�v���t�𦮯�lP����S�x��th�0�ф����p$w�N�z��ܬ�Zh!ۏM�����0F�j�0���:�f9�Q\G� ��`6�M���� n�q��׊9�K�����$�?�<kS"��+��G
���a�*[�".��0A�`x䡘P�(p��2*���W�+1���p�?+>
0D;fD�u�p���fE�Q��3a(R����ۉJa�i�^V%��
w�ͪ,{�o{<�1D`�P�")���]������V?�U��`��+IQEAo�H�p&c�ԲbM�W[(�܃ �[�����=�o�=���|�_���i^~��h%% "9��Ub�d�t���v�|A�,>�H�Z�C��3�%�X[\],7�J��-�{{�Y���"ZQg�ES�-��z�\��{�`�F:-�� �Y��\/��&��C��^˟�LU�8Y��@��4�F���Z3��л=��4���]8�b��yuc�A ��fGwk�s�C�V�����ۡ�>Ol^XO�\��-�:�"q6���}u�Q�5�ak2�t�~0�Am�5��E�$��ם$#���*�?rlC"����,��ΔF]���0�7��{LC\��g�ɉ��16TqٿM	�pL���P(�Th �'�B��i"�� �(Bb�$����3��<R[��l0/�O�<�[<Y��nrHD�1���1|���;0��:���p�!���spL���	 ���sڝ{f<�U%�#
?�=	)iGuI���B�I/��å�-3v� ��i� �x_~ٓ�هKÁ-�&P�P���/��c�,SA%!���75�Qls&8	���0��T䷎u��ҬD����Ҭؔdp1�EɎ@��-~i��
d�}�s�]cM=���{��؈##"�U_����U[eh����g^wۻ��s�u0����=�k��~m�^������ ċUd˟����Q>NԺ�;=�o^��N5?�Z'!=޼~��g_7Q�|r�-k�ҋ.F����hUrf���+A��0�O2 ����@<�������� w�HV
l� Af��"�AP q���QBp����>���***c�ɹ��$�[���#@Ǒ�A���_�������$��c|��<� ��3��ӧ9���~0h�B����7*_��S�|�e.��Z��[(e}�}�@W�@���X=�T�'o>C�;�{ļ��gk�Y[S����8h=r��ؽ�ɡ�:��xf0}^	�he��#��'�H�Hy�9~taEꨶ.��t�D+w�:� ��<x>0�o۸r��1U��&W�$��5��w���W��svV���W}N5���xML(���V5)(	��"a9�B9b�@{�6Ӱ2��(Z`��M�
V��|:Mw��j��Q�8Q�J@�q�\ ���E�� vU)�0��ý�C�r#�x_�����l���Wf���g��%�(g�H!#�����>��F}�o-z]*�M9�9�G����Zv����H0 =��
v��:��=J�p�_)/����W��q�Ж͔�	&;<k���#A�P�V�>.�䉓�w�Ŋ!U��k^��g]�������>H�(�d@$ ~'�j/�vV+- �M�q3�!,����'?k�w/��?j�F��<�����zQ�1B������2ʁ �^f��@�=ʆe�a#7��/�2��f�D����5	� ��g-qQ���Z���t`8Uf���J�L����K��n��h���!q��O�D@͟��C������/��pB���jDH0( 9�m�{�t�mFx,���ֺ���~H��
R @�nuAvm`[�13e�&Ry��B��� ��-/f���0���5��C�k<|���R���S��}_}��E.0�W|)�]�+ed��L����6:T�8\q�oB���ڷF��h.P�]��z�g|�{�e� ǂ��&~�2�.��<�_6HV����N���q�GZ�L!�`�aaC)��#bh�X��=�!H��0G�I��P`Z(r�Ttm��H�(�@^T�G����~?m��ˊ\�ciX��r]`t	ݱ*�	�0#|��Du��W��a�K���A�M#���w�@mڶP�(}&DD@�8b, EO!zn�x~w��P�N)�p�f�l������������Q'V�S�Ш�!ÔR�Lk�;J��G��Y��kEI����ᇘXB?D�����7{Pȿj�gJ��g��B �j\�EPX��� �dE���
��+~����w]Db#bF�a �b�w����O�v׷BA� T�XP�⡞H� �8F�D[��P���B�l`���5/,q_�b���xS7��U�\�,F�P`p�F � �a���0$���gBo��T(/Nј��h!��=>��G�긳Á��D(����P����~�"5Tqa O���t|���@����M	�+T���g�UƇ �ʃe�G��� �;���R���#��� ���Q�x�������90���Cj��Q�0�_����(��BՒ؍(�
L����[i�oh�Mj�L'葌�Q ���tq��U�rN�����>�^Y���Y��Up�����Q��V*"�F"���X*��,X(�� �A"*����/����e����v&��]���`B�޴�c-��t��s1������+��뙦P��7��,,��wi��b��-�bt�6;�M���5UgB1����G��N���+�����I�ВUAT[���͑)im���r���#w�ma��/�����o|'� ܓ�B	�	y��(�������0���(�R5N��ݾ�� P"䡌�b����H�I� C0��&�Y�yJ�_�����O2�E���F�G^�+��|�K��1BϏq�'�V0D�����B��7�r��Z�#�)��;��g����K(��-�$&#I����a�Z�X"�Q_(w���>@g�ȇ�W�E2V� �(�`�
(��U�F,Q~��%��f5��N�`���g�ێ��!5WCL�`Qcֿ}��P�2�xN�"3�-aw0b}0�1kW�P}�E+L266D4V򪕢d���A�D�C`�A�<;�3�;,�H��S`<��~Ul���0���B����i��b��!�A�~j�6�ъ�8�~�� ��YV��������r���Y����04jT!���YdW�v�X�<Uy�qx�'�{���&e&]$!V�%z�$-����~c�I}{olM����pu,�_��*E��M"Q���2�<E�O�7��9 GJ6WsC�_O�v�'��Ÿ��flG�Yg�G���[�Y�2~�{>� N̞�g��,�M`}�-���Op�Ʌ~H��e~&݌΋�銸�ϊ�� &W�\ٝ�f����f�T����B�Lu-k���{e���
{��:�~2$���!����2�e����b����52�t�k��6�"����,D���,^����y�X���+/����)7�ĂK�q�@�}��5�Jg�}�P�~�OSOf���џ4���nrFG�b|�C�O(��=��p����g��=�\����y����W��ʞu�v�r3���uT_L�񵏌�ٯ�����|�ED��_Ui߱�t���b#V
�)8y���u����{����,7��we4������SY��j�S�
�0�d��V��a}d�B�L���)FR�.��k@X�8���T����{�mـ;?��n�#�n�|��Yph�����O<�ݧ:�u����챳�+Vf��x�e
-�*TX�;�����;s��A�MS���?B+���G=����2����ɳ;E�I��@J.&�����x��Q��+�)P�eEq�R�%J(�U�����
!�n���-tǢ�R���>)�w�f}���Q�tzf&K���m�(��Vs��ڥ2{$�f�pAþq�n��OީN�f��p�L��x64u���UP�k	�9��º�Dm-C�z]gv*+�npjMt9�3- �S3/Mu��=�{��q��Uի�v||��֩����p�I���&�1����0��>���/'�Z���$��W�����1�<_%Hw��**���q�4V�x�g�x�C��n�kn~�z9��hK�-�?�O؝��!���1m��1�+��x1��q�(`�+DI"�bE�E+}n����wy���Ϥ/���"
��x�[{�L�+�@Ep1"|zR���t���~������3Gy�8C�/e���L��2��4�� ���,��o)�Y�=�^d���#���'f�̅F���f����Q���[r>��\Y�U3 ;c<'�!:����pK�s��@�<k�����$���ڭ#;�t�41��w՞�|�y�|!����̶En���z�q��BsM�'����|�@���\D-T{:��u}Rb�&%��3ѫ��(����X.*�,Ty%�zm�ЍC�sV�f ��vGr�R���K(�R5��{��7��}<L�5k8�۪Z�v��U}Xgh85۽2����9Ǹ������V�����$�2��E>ǮEW���o��9�����b�0����-�ۜ����NnT��%}�����4u�Ӫ���4�[g�>�T��� �p��eX�Ց��P҉+�&�L1j�	��p9�/���H���T�i�a�m@�����`�(����`��k߯����oƨ��4�v��O̖�EDF#��X���~ >��+|�^��Wmu]b�R�f��a�w�&�iN����9^���q+��3�ѽp*CN��Ɵ?z&f����;��`�z߭%x�{��}���4�����D��Z���v;�G�!<�s�.V+m
g|i�֦��-�VdE��/`ߴ\�0{�����a6w�v�آW�v}��Зa��0k���֮���_O��C"��*�*FUR ��뚫����k���ie�)�m�=M(�j�_���|�_����@�"�`LmL��0E�]�2��F`�s�u
)�Y'[`�K��Ok�^8�4���Rň{L�tPtb����j�1�T1�Ҽ�1]!�������3'�Y��q��Jˌ^3*hKN:�La�g�-lw�yѼn�mV���Y܋�3�ޘi��ފ��
[���-���p(V�j�c�4��F���kk�.����t
nN���9F�Ά�u�S*����,���7'Q���1����]��ƫ��PQulQ@v��d���f���+��VR:�3��lhn����DJN3��lw���B��c��]�\�Q;�p]�1�WG�w�݊��"�`8��X�����t �_q�5�jP��n����di�[ӻFlře�<�.�Ա�K4�����n��gm�#\�ͪ"B76���"ŋD%PYm�;�[��V�PظvV<��/ZM��+H��N���75#��W�옷J��5�t�*p��W!��BTl1�%�Zĥ
Dh��P[�)1'�@P0.��v��C��!c � H��">���da�,t��]`4Q����s��j�����_0�6�h�-�������I�,�z�rɢ�V��3�QY	�w��zOEx�׽�@]�OMhe�6Mk$�u�~4x�E �N:��+/f��(R.��-�r�KuC>Y��4u�8u �"���G�OK�W�EW��!+�%�7��f췎�à�L�d2aY��:�4�$+�	Ԡ#u��,w}�	�:����1��l)���i&[qA ���PU�e�]���q�]�(��6m�v�m�7ctG���c�&wP�b�z`��p��f]3�5-�vج4z�"��b������h�1q6�A�-Yi�]��!c�4JGE�V�.�8t�E�'Kb���Z$Jkl[
ɺ�L������؂�}F��Dp�$�����.\R#).�f`���/a��ѭ;y��eÕ���p����v�<
�Kʸ6]����wvh��0��Puv��:��wu��:{sw�Pi�sy$�m�ۭl捹,�qrm�m�Ie�q��7�C����%�0�f�4/�_q���]���e�P��9.� (��4N��v�a��;��2dc�(�]�.�rR_�ӡ�@d���Ը��`���R��+�޲4���Y�^��@�PΕK`��e���z3|2-y�t�o��d�D��؋O���%40V�0���%wh����^+�O�>]\���1���(GPv�Xt�f����9��Q��7�-v�P�[���W�+�H�F1`�F�ͤ)Z`	si�7Sf;�	M����]� -+�pNʳ�<�Ȑ�]��������2ئ�cj�S�W��X��Yn�X�7,ԡ����<�E[����8��ժ���&N��� s}�H�BͤoL���(��]�Q�h1�A�a���F�w3XQ��U��C8��#'aYc3-�ͤ���]Le�fn�ԍ�trf1;-���%.L0{�dÜ�xPo�/�����tk��;��9�{��o&�C�_F ;=׉cW�/������F��c���$	ɫ!���6��Ԟ*��P��V�yN����#�R�t�,o'۫��;5�z���b[�w�4S6Ggdh��!��gv�w�L��ܪ����-5{���R.����v-��WR�R�n�]uŗ16.�B�k���4�������k�e97nu`¡;G�Z���N栮&��f:k=����w��3C��|���Z�	{l�r��(Nkuϵ]����c���¶Afv��KD��ڧk�͠9�;vw���{e����(���_��+�S	]�7�������B�)ԝy���Zum���+�T��D��'�'a3��7ݦ|�ߚ������<��������g0!�@dRA"H	AY��7�i��Y,V�A�AQTF��bo��ڧ�~�o�s����nZI�D��K�wʫU����D��ݢ�}~�j�uwlLt�!F�W��d�l��O��?M
���U��^&�Urqs�5�����!�}�}�h+���v�X� �)��(/�>�ٿY�X��Nfȁ��T�vHٳ3sH>&�V�$3��o�!F��b��Ϋ��N���]��w�5܂_nT��5�^�`�uo�'ȈDX�����S�j 讔%z/�����'���?gr�F�����'kB�Oi�Cχ.��o�{�|�}�ې�]y�*�$b��)W�q[�&'�9�^��j��D=\k��Z��{ں{�aw�o���G�Q_(̘�"�i����XWI�B�r�.)�g~Βa����'�&u��C�����T��8��˷]�GP]N���+f�MV�]�@y�t]س��JVi��[���c��1ZƂ�V�nc]CEn�awv�=����z�ɺ�+�75uj�^�y�9�szleׄ�޾��}��՗�����`1�EV,�1~����>��{3\�y��Յ�"AAR~N�~s#c���b��as�5�;ϔ�8��떪�pQ�>"Ӟ㜛ߢ~iR�߭���4�i�װ��3o,5ϕ.a�WW��8�B�ׯb���J�.�.�?ơ��R���q}V�r5L�w�l�Gm%��3�W�B�����X���]w!��M�b��3��sC�0Y�S�j�j=�(;b܉�%J]�}�#���o�"�M;�}����|_���oX{ᕵT��ی�H��m*Œ��-[��At���L�S����K��}���M	|� _K(���P#23�5��c���Ŷ���[b�\?��T<���kx�,�5V��܁�L-�ț�~.��/�*]^�n���}��ה�9�sv�z�H� dɱ�O�;�o��,A��c�F�yQP�:NY=?j��~��S��݈/���h����UO�ԟL�Y5�|�U_P��$9��j9}�ј�gF�w�T�$�i$�7h��X���O�Q�Z�g<�zo'loy�?m	�S^���y��� ��1���̕���w
���D{;�@�_0�#�`�Aa"�A H�~ ��s��]�s�4)mv��J�_l��M�E�gC��������>����ڟT���v��˙��UY�R�S���3�!\v`�d���>�s1d��7Ϟ���g�\��^z�����k��!'�**n���v�'�3	��'ds�t��A~��%	)�Dn�1'F�J�FC��l����z�Rfc��d��J��Zf������ʼ�'��,E�1�H>����9�C��������q�*Iۼ7�L��~�鞼�qC/�g�z����m5Xprⓘ+���pǶ���ksٓ��LLV#<��:�Qs�W;rS9gk���ч��mdC�� UÙ�MZ��eR�U-[qJ�f��|�ʞ:���X���ۨ��_ ��^�]{*H������>��ŉ6<�(Y�����&1�8\˷��L~��-�>.�yU�2
�Rs]��sN�D������<����q~ޛ�W����DH�"1E (� ��~���c��ݭ���v|�k�_J|��ݢ7FУ�{�.�����qtS��f	�7*s�LC:��QT�d�⣝����"��!�S0"Ga�t1#�O�վ�~"�K���y�*X{#�c��Ϙ�	�x&�B���n�m��,ٞ��̓*�&�1"PQ�Z�xnl�*rnBc����P��ؕ|>��؂�ԣ3�K�,�w<w�����s�ۈ���mzX;Y�w[o���6�JX��h�)D�B]ֻϠN{�w
��u�����d��gI�����fP>��*�]�}��M�C�I M��O�N_j�'�d���&��g��(]�Ox�S�j
���2��:L�L�ȑ�H�ͦ���P_~��cs�e��m:Oq}5��� !C:�>�TE���G��׆�z�X:F>9ro������f]�Nhj�8kYx]��\9�	�5C�ҪD!s'qG�K�.��w�Lx��νt�{B�,�ɞ�|-]�(���s�߹�`��E�#�Q������+_=?������������舏�e�ޜMb�IRw���Թ4�	�WP[����{g�m���r�:����b �p;����-A$ (b��6E$v.M@�([c�f����'g}���l��o@�fj�H�o8�C_��i'X ����u���
	y[�ZkI�xk����9�	��Ȇ�#7*�4�墹T��ծ��d�idJ�|�)
Lڣ_Eq2M�P���;�r��tWx+W%�R�h{��j*�J3棏z�V;eW��xȭ��R�c�z������~7��G޵�;%��â��w�(��ۢ.ĳKw��a�Pȣ!�<ꥁ���ῠ�R+�W��u��+������<wc/_f��=�����S�qD��!���2�*-�5c��`�|�����$HH2W�U�s}��}23"��|����;ٚJ&�0)�ه��v��P5h�;W��#�8'Rq(�M�O��ǚI^���`�W^sF7�gl�o+��Ay�Ư��""�ε�/��
b��;�oQ΄hȍ�^��e��s���T�e����+Ƹ�'>��*61�@F�؏C(^	��43{�",G$1�~�L���P��FQ�j����as2��Nz%�)�Lj����U��TT��$��Je2S*@�*U4��P�j��������wZ�����~��҈��b�F"0F$T�a��0�g�т��N���{�~�'�(�<�����6���R�I���UP{�Y��V�F3�&f][���w�D|�$�j�4z���ϡ�%�J�ޓ	܏�"d�]7k@�4�c�/��V�;�yޟO��w�{IQI��L@���BN��<�U;�~�8����)'�^������r�OFS�7ΰ����fna0�����fo�.��Ō��ŕn�FK�*}��壀��uq�n*;�'����yx��El�%����$P"�v���w�^��L)5�3BO^5=�4j_�ؔ:+ I�\���LHb����/w��EEY�����'��3�3�~٭D�
wӭ�z�hN��#
+?a�����}��St����5CB�]iL$���e�˜�a�Yi�>��)�Qs�9�����rc���Ǯ��-���.��Y��1��A�����Ī_��3V���O�6�'�VfL�RH�U��GtQ��Uܻ5���@6+8�.~��UQ�@b�(##��ٿj�N���;�޿r��~\|+�+�zt�<�˸#V�A/�&0�M���Q�h֝9�\#��xQ�g%�PL�~.�fy����+�f�K��Z7��;z��R*ӳ� ��X�+��<���׽�����]��ܖN9˺����jm��!y��Q;��� ���.+��4U����79GDLG�5�s�KX� M�&���C��`�^=���Y��FoleA"u�iT΋�\R�!�O�0�x)�5�M�!��Z�r�Z�Ӿ@l%]ԓ�{�Ⱦ���x8̱x9̕� O| �|7E�by��z����N��=�vd��Fc��WO�O���wZ_����z�x���g�F;շ���%Q HH)�覶h*�d�rU�����28ܚ�Sp�V�|���Vwp�Z~Ηj�}�}���կ�Q���?ҫ:`HY��QZ^q����(7���%ؖQ��*��y=k|旔4q��έÞTz«�)�yV<���e:��u��'���߼��TTU@A"�� �����_�˪�wៜ�Q�t�v�V;����0�1��B@<��2;8�6Wr���%W�Cq�w��I��+AH�I���9�,�VڔG�x|�c|'�{���v{�$ʇߓ��T�Cѽ-�ӎwj|�Bgu���A��5EG���t|{FJ��d*��Ӧ��"g�[^��p)(��7����`Ek~u��w7��{��gn���(ý�Α{�Y!����2�1���>#+���]������n�7&����4`�VT/�*�4��'k^9���+�8��j���_�׳P�&�Qꄽ����n���c&
T�nw��|��]���;]�`�F
���o�f]UV�	XQʴʤ�4PLȲꈺe++��-�0�s҇�)��T�yk�Yz�v�d���O�{c̟��9^�c�{�1�ĳMTQ�+�H��u�30��8�*�q�k|q>VOr�G����V�����5����+򭥀I��;�S�W�O�n��������feM��ނ��(����r.z��skF�c�\����֜�,C��?{�7�4̹[{�Uy�����(1B"ȃ��[3K��|��M&/-逕��y��~���n�1�b($H�P@?�Q�"�zz?���,CDV�LO)>����O�]�\7�q��{+��]��Q&<.8��G۫eI!:��w��g1��yr߇��x�!�����R��{�ʔt�
0��oԣ���������3���>�,���
O:P��w��)���
�bOq��Gm�1f��UnBM��K������m*��N��3ŵ�&;z���!n�w�ʱ1�a A�N-75�s��9o��̵����ϻ�zV9�ی���H-�:^�&�9�Y�ʪ*�Qt�j ��IH�Wb�N8�^3K9*R��w68d�"c?Ӝ�%�5�hE���~,t��O��>��a�2'!�`�������#�.�沄�R8}�ۨﾃ>�s��zs�Sy�Y��t�E~��ֲ2G�i����F=��Ey5n$/���C�g7X�U�6q}�0���,,�#�{v�𬁶f7��ۤ\ve̢f���O��Q,�$r�5���Q�F�	���1�U����{ǵd꾋���tXm�D6���ݼ��fƕ�T9�Vd�`����ؑ����������M�Q��]���K�o�nw�r�o٠��M/j������N�u�(�b,)UEdRYQ��~��	��02���I	������]��f�\���4:e�MQ���gh�o�K��}19�|խ�Ш���O�E_�7kg NLM;�1]S'�ݤ0@�������Y�N�Q��ZUg��=������>���L؉
3�8=ի�1|���&�n�mP��q�ז����<��}5�X�y__၏g�V8����
jE�~7-[;Vg�I�﫨������� ���˝qv�������lV��>)z�C]�L\d�81�Iռe����rEYZ��>2u�a�HҨNq�,!�k��4*� � D"��"W�nq	;��S��9����͋ɻM��wy(&kf�A�	]	�L<=�0�?����Lk�´\䫺�ѝ*maG"G���3]3NQ�x����"ͣ~���C��߀���n�=^�=�<���{I����I�X ]d���<Wol�����avwU`
�?f��ƣ���O�����x�ޅB=K��'�3}Lg�S.�@ GUȬEE�""�Q��^����g~��H_� �����׽}���CXڜ��x&+#�R���[���SY	���7�8�.���W/�Y
�,�NT�{[8����{�G�,�y���z�&`��|�R�T9Z:|zu:�м�9��S�g(ۂ:)i��P!��s��R�s�>��QL�v	�˺�$z�Ŭ�+�9�k/M̥�C��bP�E���z��E�Y��s%-"���	C��L��H�G�R���x��z�v'�iWm��L?��"'?�r:�����
� �Q/�d��a��ƍ�G����J�jF�Ͱr9P>����ܑ� ��32�[��dL��9ژ�tS9B��lq�	�	�����8�H\yݙ��c�r㽝	��-gN9`ٵא1|�`�3j:`Eѻ�D*�o>6�#k��%^*��v��1��dw��fd�mS��Yq�-�9��l9#�#���s2	�	b��I6d�@���u�Ѱ�A�Z�X{���N<�P6F��3`�B��Ռ�]�{���s�<����.7X;YGϙ�H�Zy���#GoW�ߒ�K�U�cD�L��Ae�^���o9��5�6�(X%�j��Tu-U�j'�lI5�L�ա��8:n����JD�������0t.��W|�T^�~T�����n�\y[W�s*Y���8��=0���r�}n|�i���@Ķ��7�ѻ��-)B�I��{]�&�n�Et\X���KT��M̶��k�=E��V���l��%_J"��(i(�%+��q�!�̩�?�bH��P�h��BꊩV,�����|9��y��U�ԓ�jZ��J��/
���m�}�oG�ܗ���]��b�ꢽ��<��t6���ʭN�tv�� �$���Е�l�8c��|�&�M��;�Uh��hR��Ɋr&�Q9g����Z�|*b�F��jyY�g�LX�S�|E1�0���¾�Nn&uȚ�~޻���E�^,���=�v�+SkBA���ѥ۔�1p1Q����U��
+VS��\�՜�K�P2p�q�В{��ݪ��;�;]1�y�!��/b䆇�S�����i��/쏺A��^��wv䖕ċ�p��S�[�F�>��\�^\{Ĳ�R��b��%Eӗ&Q�L>Q�!��2�����Yʀ#.]�V���s����8hW557ΆͼkB�v9�Ӷ�8k1�y�v��n܉�҉=����x�f�)�#1�|� �c��� �Q$*�
��vȔ�j@㯳��uwv
��7Ss*Sg7��P��UQ+�=�����{�*�)�q�{Ҳf���K��[d��亽�9ИF�M�zۭ���bb��w zk�;�fJb��w6`l��:)�{Wu��u����R�I�62��A0aY.����'u>\�r"+�֍�{��SKv�G[T�-�6i��h��c����o�H�l����^2҅A�ڶFԬu�q���u8#cNM��;r�j���[�f�z�bG�9C����~��iI9��<�fa:��R�=Ġ���s�|��rQ?S���U�OU�qvft)�	{�g�$;��pg���v�?�j6�_��|�;��I��,�ϲL�>����|�u�]t�ٺ���Pw���"��r���� tw`�;Ut2���s��	���K��tw��7-~� c�Ġh�3��m����!,�������\Y������:�č|�h��=^�u�!u<���w+�h������f*���#�+���P�\%��\��KL̯�0R�ʇ�n'G�����6r��3 #۶�^������)��HQ7���
�`���`��C?j�K���+��*m�q[���z�＞\��-�ӡ�K�AȇCo��ñc\����lk����c&M�s��T�e]��=H	S��~��m���N1������K�t�⣝"�oӮ��,�"�l�Nc�N�"!��k���4vOn��2'�2k������E��j
��y*�����������|�a�}�jSfd�A��hj!���� ��]Y3��e�����G�2ֶ��sߎf�7�H'��Ŀ�,c�k��}$k�Z'�g�.f-�j���KޚV�͉�2������j0�� ˮ�̏�������?L��8	&)>v`�L��MTb�٧fdv�i�||z3��fC��~ͯw��z��
{�U�}g����6j���̢�bj'۔�ׇ��6��)�G�.B�,	߯!4�"��b��.����|�X,�ADY����j���0����?s��{��#���Eɨ�ST�5�,��pd�����ʽ�=�t#�ފ���(^�A9#K�ף���}
��Z$ٝu���E����,�}�Ϣ"t����Ġq���Z�c�$v&^t�WM�0�v��C��yf�aXJ����=ٿ��d����r�Rхrr�_����U釖z�O�v��@`��noS��T9xM��|eٌ1��lT�H1����k�O�����R3�.����=c�jc&;?��U�p�7�u?oEץЯG�D>U��\~�8�|���?~���0%�����`�@Y	uҝ�����2���ɱD�WQX޴.̶�t�1�	Dr6��&a���V?�O�Ω��L�s���ܮ��gp$#��Eoª��#����ۡ[Z/��W,��g=�[���Stl���0�[ڬ��`�gFh*mSe8�1��%���Lo%K��+Ġ�B�#w���m�S��$��������v�̍���m�ފ6�v�ߢ �Ot�u�2h��5��.*MC���:<d\.w��1�c�6gew��Z��4r�S�6�1�*�U�1�JJ7N�^~��ATF��� }	Yܣ��袔�]z��%O����>����F��O��)"�W�*ҡɤdk{?6�i Y{Bpt��}8�l:K%g�X6�#�G��^3#�����#h��)���3�����+�-��!l����F�O�dq�;^��2'��F�:OGQ�@��7�<c���}�tJ�F�.�QcaϮT�/f��C��k٬
m�w������k������0��o���S�������z�>�S���S���^���O��(��I&@C��c�X͸֠�j�i2{���N.˺sE�Wg���1���P*
�Z4+�����F)}���^���\�]t�.a���Ӻ?n��؈@��T!I�����QQIN�����ql�1�y%�b�b�P��o3�����@�P��q�IHP%.���؟ 
�"b�������w+��5@o�w6l\�>?�G��yo�9qj��^�Y֠�q�צ�MT���cd¶<���u�|���Az��2�̀3�}u�m�px�1�ϋ�������׺c1Ȑ�����m���[ �Y_}3�}�^gxJ�0"�l�jnoy�B�"2(**��~��?o>��Y=��
�&��]E:P�/U����R,�w6�zC�}q���3�Ĭ���]U�sɩq{���g�KDɚ�ʂ�i�?^T(�B+����n_�>�:*l��:0'DݳE�DD��bk�w��ϖ��z�l��RAMx�&H�H�h	7�P�V�L8<�wƇiuT�\mԙ�1bs�O	g����h�����ק֝?���C���}G�E�F���m�����c�;����}M�8]��1A[b;VI$�SG��f�-;�'�ݎ��bet�żc<����&����TL{�bבA�U��1#�?�;c�~�j#~8x�����>���`^3G����{0���4Z�}mw�[����q��v<�E�{v���Y*@��,����y`�ʝ�Ѵ�l�s����˸$���'pmi�q���~
�k�É�#�vf��?7J�Q:���\���z�ߡB�c7�ݿMϳC��P�сi�{󄅄/:�(1����}�?^����.;��M$Q��U�
�`���گ7Ѯ���ܟ(�U��2D��1D3_�1�Q"۞�k���t������ �.=����~�ϻ��
���,����f��� a�4׊ʼ��?\c &�#�~AlE�Ab3�?W�nɬ(�O.�Gq�C��t��tWh~�����}�\��{��TTT�A-�"��خ�ޗw�s:L\�g}���/���F����f}�Po�Ta�ڀF?����]՟w59'�����Ȓ�5��~u]��޿0�dPTb��`?�3�%_�RH'_U����KE���O�jrӠ�5j�g��	b�Y���E�M��Q�HNg�r]دw�dßg�_���C�Nu	�)�2 ������\��sX�D+�vwu����;����]�`L�R���N8-�N���7qJ|-p���1�D_�{������^7�{�����M=絮�;����@d����*���:���#]}���ǱN�.>{��r��x�'Q��i� �٤���l�i�{�9.G߲š�\ڝ=�b3�%TPm��%�q>���n��fۺ;���{���2Ȃ�V2II��,�A��a�MO��4{�f��W9�#b �
1�APU���������%�L��U�>���o�bj������D�R�]��H}y�p򿻇;�ɶ3���z�O���#ą+��tHĦC�G�#���w����˅y�D#)A�v~j��Bw�Kǝ
D���|� }��*q���jU�-�>kh��?q^yeA ��� �	��{��F��d�LX����Q0WJ8�r)P.�H���]gH�O�s��ҡzN3)y����z�1�������}� �������ɯY��Ar�'szJ��u��w�*A�!6xg�Z�G���J�|�P[?J9�P͝T��ъ��ŭI��S;뛨�QU3�u��'�F	wx��Q=ȏk�>4����EEfu��fG��y��B6��-ݘy��L�U��l!@��gF�r����R��t�27����}Z��{��rf�wi�A���_��Y�9��M�$a$ۍ$d�Zt�@���1�%^��c!^���IL�nX��[ܱ�GK߸>+_˅���/�%8fR���I��l'	�m,J���(h�݂��.�?�@�Sa��6(�bJ�Yw�O+\h]	�����)�A�H�)�� C"��0�"�f7D�]�S�Qצ5��kڭk����ܿ�$񑀀ȃ��՜�������QU(�b(�R,���[̾f^迯��K�МH\\�S��}5�/����q���nc�"q�+r��NӞ����]���.�7�h��Y�U��z�ﾌ�`,��n�gv7^N�Ew�B�V�ލ���o����C,�����mr�-��>XL���W��xe�~Т�ù��{���fǗ�s?u�����F(��`��!���[��ܽ���y���ꤎm<X�f�z��G=��v��'�]��Sq6����u~��r�q�<|�E�C�4OU]�˭�2|)\���Gݓ������iKˣ�G�>s�廘r10� �f�b�LЫ�45�]"3`yq�C�ǹ���������W\�tV-�*
g����8�(�˶u�b���|G�n�	�3rƨ|����6��J��X�[�%ʨ���$ H�",UP c� ��o��=�d1p=��8` ���q���}Z�A#j��"���i�;�sW�>/��8{�NG�!��nO��.쇗#s�I���-��^Cң0n�K��&f�n�GT���t%t�G\[/�}ϕ���1�^�(%�G���ؑ�9��"M:�S=�٦��2�����=躛�%��y��%��=qͳf��㎈N�deq�g�jU�iaa<Jzꨭq�>� ��ʱ%9��
�b���C;TBT�<�U\^oTs����7��|��8w�xnv+Ӵ��4ع�x�~v�����9�|��n���D���A^�f��T�gc��Q����/�~����%��~L�97n^tV=Z�̄�2k�±���d,���g�DWz���障��uղbh�nƕ�kE"1P"�g�z���t��7����;��>�T������#����YEuw�ig��}v�\h�h�:��Rް�w���P5�^uid}UT����N���ݵo�� ��.h�]xX����iU*�;+���t!<M��彰x��G��H�h��K7.kt'�>�
	�4�����1��|s�RD�I���8ɷ"{ϻ0�v࣐+b�j�3w��=��z~����)A=Y�\�~~�G�k=5�s�6&b@��r�\V־>[��C(��ˊ��]�#=O��Mi�b����뚷6���{���xMY�̍@�]����8ۓd �5��|���"�u����u���ΘW�F�mP��aG��W�,7l�m�x98�fO�����n`T\N�����Y��;��t�����=9���QM]L��6���X�c};��FW9�M�U�����=G;�^�k�&�GWM��aw=N�����=f��3���{���o_��>�+��$��&�"�2�!^�>��s���7��-"��R2Ȍ��R*�^��A�x)���Ξ�hc�ag����墀�}�m��9s꙱�94�ǧ��X��y�HIāF��y�{^1��6�b��(q�v`�������ҕ�$Ɗ�ӹ;�إ��W���1���Yx"h�Z����)�\�(��n��+x���NP$ya�O~��ZnV{U_�z\yF_j�$$M���$Ȳ��()��-����fD�o�N�
T�o�ИB߂S���-4Af��Pw|�_{QM_�����hms�E�ީ�|�!~7�_�Ǖ·�]g���
��?W�������mR����=��B��fA)�0�[�c3;��s�l�W�%dT�9�<�Х�ꯧ�6�>���^���~�ئ=S������޹�ܫgY+�I�t\���~~�fIPľ��5WT��:q�z{"�sP���ق_V�O�
,ADQ��EIC�g��Z*����+��~ ��
����]U��|<2蹖o�tu�sitY�����b��n��.3Z�E�u���Ku�i�_�����e�n�V�v��Mn=��((��Nbvfm)���wo3&jZ�&g�hb�aB2�SJ�L���=��5�;��������|��jq�/s���{�G�.�I����<�.�A����[��r�NVJѳ��-	,uc����B�u�
sb��K!��L7ga4��8������A�L�]'$1%N��1���;��p��naX�G��f�u97|�9{�R�L^M��"`h�Uw3�q�B�#Ap�/V V���9��D�Mw���ْHx�o�R+N��7��*�ku��.��B�`Bl��.z�����Ϛ�ܗ�w�F�\R9�kN'�뾂*�(��q6����V�aE:=�^�:#�дӍ2��[W��7ÇYC�d���b諩�x������S7Dj���֝8Ѧ���J�It��ʦaXCI(;�uc�6E�m�������ݫ3(�S�u���QI;_G4�2m���탂sa�e���\�$|�!JF�
k�m�GLu1��m�L˖fǒ�;zm�x�H
<a����c菎NU8��&��ݴ��*ݹ�X���n��� ߾���L��5�ȋ��Ac��P�>TJx(,L��
��W�pIõ;�A-���nw�����]�SQl�-C����l��������*�L�U�--UUB�p6�K�[��P��[M�9�Z��S.UUҚY�iXl��W�È6�A.ٲR�k���,��L���R������ٶa��W&s�i�i!k(6�dL�D�%�-1���nc��; �a��JF�[uP�FHiK*�6�eG�7pQ�S<�G�B�I
F�U���r&����� ����9��ՙ�7������e�86՛� �@������1�yy��8�a��[�����]!y�� tҒ��F]�*����|�4n�Mg�o.�Tm��;+����՝٥ndZ�U�{�Η��<gG-����Ǫ���bX���l"����l�;�l�q� �K	Y�F���2��|��8+���@��6mҦ>1�{��$�����5�W=ssN�����s-%g*�B6��V-)*��v�hV&�ɢ�]����61j�f&r%��GA�ϲç&Q���sy�h�ui'v�]p��+��(��ۜf�t�+&u=��2��*Yغ�L���d�X`�J�:�w+�m��Z�������,�v/��VM)-J�����᫠�mK�Ko����H�o!�WB;a)��Ɍ�u�X�ݴ��r��9���hr�)�Դ聼���ᳺ���ti���(�]
��PF������Z���K��2��6�<�Ƌɽ�éF\@�����ݬ"����T2e&7��0u�KB�կ+�̼��ӭՕ6a�@)5N.;9C�8l�I|��m�a<�<� WP������ef[X��J��A��T�圸��st= �ms`Uѫ��<�eM(K��{+��b�A�8����Kܼ�!�������u�Tp�f�.Z����)�YTm�-Q�q.���z����noKraFn�����m�0'`1�:4��x�ӺY�M-���uͩ8��� N�&��E�n�F6���Ra�e������W��w5d��3ʭ�*<�k��YfB܍��X����F�����{�`p�n�[��~�|d\�q���*�u�̜^}s�o�8�>�8H�cG"�D+��{]�x�2��<�#8���:z����L��ZoCم����U�&:W��8���ETA�F0b�Üթl��컻�]�d�U�6�aD�'�g��euq޲2֐	���� E�}?���jn�=ӌE�G�uU���M�T�ᰩ���TZ��+;�����Mٮ�!�Pܛ����Z���n�!2��3�9�u
�uwQ@ ��)I��=z�kI���8�F*"" �2o��|�g*���z��Z����A� �}o��I�w�j3���#�L�#Kr�������J�U�� B�O{Mn�w�׃A��vH��V�׶�����ח��E�;/�j�~�z)|�%9�UWg�og>��*��LK�=H��g��5�_UP_}EZ������\� $Ր�Mξ��R���΂<�)�Pש�`�$X����9�is82s����r:����P:=���B�N�JnX"fz�.a�h�V�S}oΞ-�W��>kk/��辪�>P���,E3!%{X^��ok�i����{��X��f�����e�"�q"��P�`���s�|L>�}�~8��P���v߮�}�8^s�=!^��isd�Q����q5�2R�/��F�W����w2��N�*�J\q���	�Bw^�[^���u=ͩM�F�[�}�{{�n9!"TL�U��Č�r��d�n,@�`#��(�l	ھ�����O�̺b��`��X� PA"����&V6����v�ՕrM�<q��a�)��R���'#9��Z�F��>��0�>�h
��/��	7��vR�퉱7��a����`�J�~(�*?~�g�p{�.}4�b1��\Ԛ{F=>nV�W\7����1"��n�w=����l���I{P�C���{ �c�1y}p������pK�F��~�3�i�'����z�w6ʡ�n��P��|t@,�k)�]�^����~�"� H"�Tb��[���sw��yw��g��j)��Ԙ�u9s6�kD�Şx�S��0�߳��{�Q�Ki�ٿ/W��9�8�K���K'|�Em�#ﺶ�T�ud���n���6�o{�i�L������c5=�Q�:�Hɋ�o1g"kg�v����+d�5�}�u;���V��2�d+���*rT>}��b}S���&D|((�Y�AH�`�DX����������3��?~�޾�v�9���׆��͹Y�2�fKo͜�96L#&�]Wt�ԣ�Տw����W bf}eʁoݻj'Ew��ZA}}��1�}SR:2p��5�bo{�X6������2��޸���D��d}�_��]�ͮ;��s;����X�Y�}^8qp�`C�u1a�&���v�Vk>yٗH�n�!ܛ���1o�9՚��M#��!۷�6���¿U�Io����ks-;y�W5���ϵ��!�v
 �~2�������"�����m`W������P/�+:�|�����r6���*�"[B��,r��P�m}n|�yŝ�^w�q:�Jj��7�R�ʧUOl+�>
E�;�������R��d��ѺiX�w"����Q����Ӟ9T�oyIf�26�#T^��ccЧ*o��ڌM([og��OᄂG�*����$���|w
�������uڸ��#X��UTAH��E/��x�h�׷���#f��o��9�;m�3�~EU�^.�U;�K�9�;�KWd�~�'��
>���Ne��inLăz�\gjiApP�΁s_pk��x쿃��7�?�+��3�R���Qts�sу�O���C)��4>�����b4J�;��Ot�/��r�iQV1`��PdUQDX�1A���*��T�R���K��W��u�̮ 遀�;4"�aF��@n�k��nw�Ǡ�v��:�&p�f�C�:C{M�)+��\��m�)}�1�uK�m��sj0e�
s6���)/���[�cc��&n��Ѭ�A���4%�� ��7�
v	UI[����e��Zʭk���h��$���@� ��FC5�)�mO�#�ըW+�ܜ.��o���{��8�K��zw�19�*��lʹ��;7>�=og���0�ndGы��7۪�٪��CR�����tmKc�k��n�*�W��v�r&Ra=P�<qn�]_{ޅ{����4k=��w���۽?���i$�Y:%����Sz��F"�+��%e��>�g5����g�v���&B����<�W���w��L�"�M���K�Ɠ��p��6�g�X��|Hx����������5�{F�T�����u��0|*��V�
�hF0�x�j+f6cdR�)����f�l=�\�^������Mh���lUm2�����`�ɤ�fo�}¾����'���*eM�񎥮��-��$,<��t��~���R��e  �}����U�wt��sݮ�,ogq��Xmj!o�]c�y���C�=;��"�����M��	���?�R��Qt���cj{���A$~��ו��[-��N����@~�!

������3�l��L�g�O���U]�O�d�`��\w�D�W8Yn0{�Ŝ=i1$[/ol�J&[�ڗ��~勒
�EQI ��}����[֩�
�N�0b�"$@A]��W_k5�YW�j�9�ij���ŕ�\���-�������]�P��8!�Ss���r����7�v�̹��xs�����9��mgɥ�+%>���mD}w�O�g	-.�������3`����/5nF����@z���]e/?{��� ��o�����ےz~�����睅�}���#*���w��'����n]�۟3�n
6�>��{O~�ܜ���~�:�EG=z�H��*�V���_jqu]UW�(칭�|�x(�7���mɓ�mo�ε�J�@�����������ͷ�@b��N��l��L@I��H.�9�k��˱�A�ҷPݒj#�d����#�Uw�@�&��r�^e�1l�UϽ3�#���;���
<��lC<XNJ����ɗ�ӛ�~f3��6��O����Y2�z߿{����_��Y�k��r�AF  ��H�,A���x���t����!��w��"����#�GhTϫ�q��}n��ͨQ�*�F(b�4�8�у�{w^T��߫ 7��E���1����q�}Ϝ�ۍ7T
�j��C ��>�=4�չ�n$j5n�q�>�>�����u*�cy�'b�5Lf��;��)%Ti�1<&�*��~̿� �×Ns+ڥ+��c����P�t�y�j��Kk�:�xm�d2��%�X�g�J#:X+][u[a��������������RH��N�z�ʬ�V�N�s�󵚞�);�=�v�\{��ą�=�(�9��p����EY�u��j�S�ص�F~ެ�f�[����d·���D�ls��ˍ���˜�~��'&��|����s�ُW�n	4�6��4j<�b�c�I�:Tj�@ĉ�~{�8�x��������$��"",c"�����W�,F ��AD
��?Wu�o٬ѯo�����k�fy,�/�R�kj�c��cv��Ug�~�H�.����.�C�.�T�٬�W��.����M|9��-ЊF����{^�������v�'�b�F�ŋ�gC�x(S�1����6��/�'K�[kVر��<G�z��1V:�	2���W~���O
 ����@�ow
+I�\���7��s �]}戊Kr�V.T'�U��� � �W�����1S�}ΉVp�~��_�@DB
�]y(xEg�Hv�\Ϥ��ۖ W�����/��^��i.`Q�]�HU|�U|�VU�qU��딧Xl!��:̩v.�f���c�l�_�w�]�f5�r��a�*u�"t��$�W����,&�D)׹��!� t���=��&ӘCi	�"A��'\f�2a1s���O�CNm��y��۬�F�dꮜ��B�;ܓ)�R
�MN)�u�u8��5� \d�UugG_��Ŷ��I���]���W�L�\�:8��*�F��޺��T"��nb�#VX
�
���ל̗|
�HE�w��ݦ��⭧��*���t�Q�������Xw��NT�T��B�^z�{��3"��"�dI�`�䯝�R�+Ff��������Ѿ��3t�H�������B����+`����������Z��@<GG�����}�=�C�q'��I��o>��U��*���;����rRA`�|#���菳�%��N�f{���dO8ZZ;��P�y�|�srv�)"H�eHi�n���V��[R��Ҩ/{���t_	����)*�{7��?go��ޘ��L4C��,�S�ꮮ����wZɺ��̺�T������A-�*�ӵ`�9��U�������;�z�h	�E�
�dU��*�쓭���^6/8N�o��fKL�6�W;��J�����L/��xe���!��WOM�j��{gmy�6<v��n�B>>���d�X8�e�X,�ʍ����}0G]����
eW��b�R"��T���Q���U�g�7���`ƪ�^��] �So������o���5�̹������������dFkB� ����f�~���M�0�K_ .er+ˇ�ɐ6��0���}ށ4�e���q��'�U~���zߴBןN������X��ג0�A�Ȉz�f�4�!~�H�4m4��&����wU""$�F���A�,�ܥ���ԯe�7#� ��:k���{gkw2;�>\��A�����{�������	~�}���^����yP[�'�3�`q��2�~�0x�ި�[T�f�UB��Ľ�g��'�zLOF���J������*��|��d;���N�$��E;�ͧ�m�f+�yZ�W:�TZ�n��(^��BY(��*8mkL��u#�9�;w{�:3�fs�tV�D��'j���P�be�G��H�r�˃�`�m-Fd��jBh��b^�1̈́l�V"�JGzb����Ûu�bY�[��F�[�2�(�����t�;�'�q]�D�HT�-�XlP��}H:��lf�ŧ%�p&�l�b�k М-U����<)�E6i錬_V����ug6�z�:m�L��:���>G��Ycn-P�"-�,�:7�O���M(����,/q4��N���	{n��m.��8�8�EZ��,��Y�_5YL*J��K�N��)J�k�7yHV��k�n�pͣƟsm`�~݀lU���XpV&
���eӸ�+J�������Թc1����Ű"#l��y�{N��`K�@hh���ns���-ao��ƳyJ�#�~������4�a<L��}�}��Ww4Z�
.�qޭ��$�>��Bk��zz]����]�2�\5��iE��c��V7aj�5�r��5nQ&`;�yಞ-E���v��_�(J��S�:HHH�4ɇ9i���+^љ�����o	u8+z�c+ �]�?�*J\*sy�V�0b�{7�7�ûZ�:�t+f�R�YڝK;(䩪��Y���F.퓅]_ّ��+�4o{7}��	IGU�0��lvS��{��aJ�EK�m�(�}u����2{wM
��ro#ٸ�ՊVZ5�pp�ha����$�rd}R^-�<w%u6�U���w��c�f���;+�����pWT�k�zQ�2��-�ܜXv�v�.�EQ�Z�Xa��OD���C�[y�B[x��f���
,<E6򘜬��"�)%��S��2��W{d�X��f*O����Ep�o�s
�����]1k�n�{u�u�P�]��la5��O=	�8�n��
���E�%<f�{�2Akk��ym,�����!Qu�H�E	�!O�v���P�	2�w�L:���4h�KNj��a��]p2C���Z�F�s�3�;n��8\��-��P3����٧�v<��^�d�o;k���;qm몭���,\��g8r�.#�q�_`ᦳc����7�τ�'z����v�v'ε�@�5ϧR�uc�[ä��+󜩟5��s��`�wU{u�|�����	
��lW��~�Pł,A`����_k����V���W�-�U��G�M�u#���?�O���p��N�tCӡwH�����ϳ�9+���1q^�}��ޞS�c={�W7JsU��q�D�+鹄�"�����
���%yg�z���Fc�W����d�~aݷe�`�)�T���=ۯz)�+F�m�>�D��I�>o���ik�'<�~�3;�\��߄5�#]�%�5+&u�I�>U�ڛ3�G�f�e��z��z�v�,�����O�xf�x��_��0���l<�d췬�索a�q~U���8����b�`X�>��_���{��&��G���$����n���l��[�3���Z�s9Gu�_/Z35rK�1�QUX����`�A����S�+�s�W��̾U&ɖ�	P\�he�n�5�(��iz�5�-�=�����W�k_�/URR��Q� �� }�1���@|��W"��u{=e�Խ���q�w���<�'�&�]���G��0GՏ�Am8�B[��|]r�}h�*��;c�U��vӵ��:Z�;��{޹����x�-b�%\R�ރ}f'z~B��l�i�)�Ԛ+�˞*��^/����5G��\�����=�}��WT�}�Fy�a�ۼ^��)��^���b��=>�'�U�P��:*L���Qȫ�����J�& �H=��K�Y��U��� Ϊ��P��*y�D%X���:��EڼswR���'�,�|`%SYֲ����4g�<��W�{�ӊ�vH�T<љ����TX���#�o��:�l6��pW�/O�V�
��3+��pR�r�W<��p��Db��P�E�*���,R#�E�R�,��%�G�r���)�$nm��3�م���]z�F�4�Etir��;/����s)�Wv�8p�q0+,�r1�Q0��b2��j�P�pUa������`ǆ	%��MN�X����Q�ܑq70]�svt�	��t��DI��[&i0e�:u����,����<��lg^D�L��G��[���XxA������rA��uF�����e�ϕ�o~gn| �c�^����cbC���}�QT�L�ÇMYŮgn������I��UK�#�.�2/�B��v���|�����O� ��	RT(*#LC�߸����w������qL�>�q� *�/Z��k��4�����[��� �0���ɩ̭�u��U2�'1�{僚�KOX#�Y��}ꜹ�>=�W���lZC3�ʋ���r����ޑB\J1rK��E
���Ě�[fԙ�Y�������HWl]��s�y~�>�8̿�PUDH�AV@@��� D�AF(*�@AE{���>��ks�{�sst�u-?.�{���PaP�l0��^p�;Iʲ��Kp�@�e�T�O'Ҹ}��S(�l���3nu��2�8����AuDv[�.I}�baۢ�S��g8�4
�X�~و��s�c6����6Yn�-���VL�}��� �S�}]����l�U���X?9_��ķ[���m����b;�/=D@^��T�s��]�������G�s��� ,�VJ�］Y~���^��?d�Pj1-�w������wd�X2���/�HI��&�Uʚ�9��q�ͭ�[�k�[�	���ȿ��p牏"y3�r�)��S�D��\��m�#W�'}���t̖�=��}�p�v�s�׷+w۸ؘ�좯�x��y�gn(���Ƶ��z�+(�EF�����y�w�N������uߘ�}03|�'W3�*�)����yB�.���ꄏ^{�-�w��w|6��w�s��=75nb���d� @���㼜��9��
��{s5��;�=�� �ŷ�A����+��Չ-�@��ڊd�&XV��F�f��)�k�c~ s����ڐ���_������ݞ���1���m������
t�{�a�8�'E⹝������mF�߯�Ww++���Ow�@�w Џ��s;]C,YY�n<���9�bPF�	I���E�"�N%=�F�-�
9g�A*:�g�˻e�ӝǨʩޮ7�q�ըՈic��>9�?ޡ�%,D��	ъ��#KJr|�}v��W� �^��1������4g�WH�>�mt�	'e�u>D�rlM�Z�5�@���"����C�yӚ��YƑ+H��(�$�wy�kkU����X�����t`�=��'.(|Q�3�Ob$�mV�k�*���,L�D�����Ki{ G�ۃ��W�~ˮ��i��\�ї|��A`1Y{~z��f��0p��6CY��j��P+Nb� �h���Σ��ۨ�d}W8����w�G�wr (!o�	���WL!�J��N+�[^9;����IB6ɞ���=�4����W\��Rs~h�Q$iz��}>�����"��t�L�Ʈ�w���3B�!a 1���+���������_o^���j�jQ%_L���㲸g��G�2�(��9s ��)�^�[�{�<����6���Ѫ]�V��6M�:�f�?(G��m:�k.e��x�z6B%hn�x_6/,�j��s�u^z�^����D?Uk���ޚ=�<�ܸ9�x�p�xH�+"Ŋ1��b��QQ$F* �A\u��_V}��<�F��Sc�K#��VEOO@��đKԽBs�`,eǔ�v��\�#��9�ZV	�x��>g���@�!��}����[�0�OS�Յw�P�Y&�}�9*�/�o�[ūɪ�TUCH�e��:>�m9�V+�٪��:m���",S�mR���ʠ"�J��
��o������a}�Sw�wG|���T{jO��9d����/�$J4n�K-�5���w� �sz�#�Hc6���E��Ȅf�j��&�U���5+��@�A��UL�6�E�5b0h朹S�B<T�ym�]m��w�M�mN�Q[�n��޺c��(���|to����z:��G��X~ Q��w�/�^])�1�|W�5/o�^2�����"L��c�dY��`I�9
?2w`W�uV�-'k�R[��m?a��S���Cb��nm�_�����V}|Qꨘ�q��l�B���/��̞�[�>�U {a�Q�Gӹ0������ �
��IF��֣d��n��
W��
"G�D^[�I�d���:�D/7-t���/�A�h�_A�2��k�/kc�����Tb��%%c���m�����;�����p��#=/�N�t�l�y>��v��f���2�o�-l�7&���H@q<:�5r�/���d�^!oì|���.�#���ϸ6H�^�.Tslz���_`��Sv����'m좵K���f'Ւ���-;jR�`O�ge<�3��B��s�f��?7Z?�j�9�������y7+X���B�!c���� >�����m���~�1	�y:��=��F����,!��Pt�Q���R�w�/�t���y'��e��"��&��½������y��g:����N<����Ԝj�\;"u�ّ'����^��4��9�S��I��U�s�-�9[��ci�c�����$b
�M�����������z��/�1`*D`���)�z�f^]�X��0|�B��IUr1{a%\�M�>��3Z$���&�GAv���墼�3���϶{�M�|�su;2���}����XB�y�NG�%�r��"�ҟ]SO+����
ʠ��7ܻ���<,�}��t�HM�F�[�?hT6���9_g�f�7�_+{4�u�$���h��/�Ѹ��3_v�U�`�'e�6}|ga�6�����[S�w[�_z{�Y�v���u8���d~�֧��Ŝܪ�Q�n7�}>M�f�n���=�u���(���]~��e�c��v\���r���t)���֌��<V�\M�{A^����=@��{HK��N�
���&tj�izUGH&=V���$P�8�O�\1BKD=�����f�˃��ߕ�[LMT\�`D!k���s�yb0)�B�EE�P�,�X�UB( @ ��z��}r7V�����t�ME���D�'��V{�Z���\+��ն)����b|�� �����d����`A�u�����}�1�~�-��V1��_5ӂ���FE�N�>�3,W�l3�pZ�qy��g֭)�p�	����d�e�)���-x�L�}���)w�4z��h�v?f�!M��],�i�WC|/u�޴F/YĴTdDEEQU}T�0�(QT��C�y˹�<6O[�x0�Y
	y�L�����`�{��%�sbz=>��Y��Q�+��R�eFʷ�������x�Ø-غ��~��:���89�8,��1�Yخ��pԧ�X"Q��Qƽn#4]�*b؀��럊�{y݄�Y����� ��#��V>���W�s7=�q5����y��a�z�o����N�;�)-�b*�1��H2
�_ky]/���<�~��Ο�D=<��w���}yO>��*�k�_�n)�����xwV�|_���J�.oq~�����������g���3.�R<T#���DG��δu�:��R���c��&��}�I��7[)C�^r�>ڥ[�O����,�m�ٍ�����3Ɗ�Ssi��c�^1������ٽ�8���0X�Y�b'��[1��xKy�U�:�6F_�?��[��y�V��[�����4��q��H����P'�K���:�۳v��0�+�n�X;rC�@�t:����.���em^�s�n�q�O��N�%�J�*�M&��ֹ��w�jn��@��Wf<N� й�3�VBED:N�x�Η�:��� �R��P�:��f�E��#�j����؟�<#�x��gR}�H��C/gRŤ����h���P��B�!n����S�=�쩉�dg�睉��N*K�{M��I!Cy�)}��K��Nj9��6,�w-�� 3����$�YVʩx]��How�E��)y�"�f�'ۥ��P۔��|��#�����4o���n9�p������X]�
Zo�7M�ס�l�i�2�������t��r!��4�8"<�^�n�ޯ�2U�� m�Y ��"��3��:j��Ea|ڡ@���#H�3]h��~�g�������g��i�U60�̥N��
���Ԥ�MP$�!L 4��@�.�{sZ]Xo}�TV�ɟ>'ല��"��<V���)��jPw�)pL���z9m�B�WC5�B�Ub� H�n�5�UP��P�My�W�0��C+.��&�u��5��P�CYd,�
�Q�Xܑ�ّh��´ɜD�Q�cL��� JR�(*���˰概�eSf��ܭ��:�r5�*GmtW �D�	�P���(�0��\�êЪg��KtBi�ȗKqc�m�
�;�(2.zkFa�X�E�n�C��;6���s��X%�\�R7m54�O�2J1�Lq4��#��~"�rgG�]��ܐ!�*��4�;�s��v��4f�K6��0�����	�"��׆.:x޸u�N��,.��R�6,��5t�KD���Y���K��ufqg���̣B�ՇO�F,�)�h ����*�ӒU$�m�ܒ!�j�=�*�w9��ɐ��'1x&Q3��0K��fT��ړ�F0Ί3�Z,ӽ�-�A;�J���yZ��NV/��j�w*%�lz�-1|[�#�݌.E���v��$i����K�X��sݛ�}K���[�X����2r&FZ�ܫ���3w����Ȇ
m��"Vp�u��onY"KD�d8T�Fn4�V7�Y������'�/2F�v��˷�r�AW �H��u��>�09�th���M��)K����t��$�;ep�r��W���\2BW؆��iY�+ѕy>x�"'�kn��󏻪��ɖ�xF<k��}��W��cb������E�U,nL5w�Yy9�-X�n]�g�̛���B�U�>�Vv;Ύ�ڭ։��)Ъ�����uCx` ��w,Y�WRe����Dwt�Y��z
ј-l뮷a�A����2'��L�rѭ���0gf����i��ONY���RZ�����>#�ZL��9]��n��"p���-}��
�S�f�죻�k�T�c��:w�47�ާ���A��ɦ-�r��u���3$M��#f'�lV�P�������V�R���,��K�9%�� �;Kf��j�+j�vP(����-,b� �oLs��f�!>q4�X�	*�"�xоj�ὶ3:�Ӳb�Ψ�<O�yu�̾K��[��vz�,��գ6RȴXtvK�-�@�w)B�.�����;pLi6R�T$��l��E�5Sm�_;0� ���F�B!��������ls��k$��O���Ll8����w��}�p��:�NTMi]82^͍��yH�~5���yʽ�P�FrX��{���c7Cs�5��(Ӫ�t��M�}��h}� > {+���~���Φ�EA(��b��EH���H���k*h�N�6�&����*��N�/>z��rd�>`k�.��-+���m#�M�ه��7^��"�G�������*J@7�Q����D��b�h<�p0�� i�2���I�X��Ae��m�=�/�N�IpD�2	10�^ �p([I�0�p.��{�>'�7��ԟl�}�u_�jB�3�nIF{���y��{>��_b;L^��g���y[��A]x�� lΨ��5�Q��uLy[���xӭ������|�?| ~���.L��5ԑ3l)�M��R�[������+��<�H�ce��YB��u*[2f�x^v��?c��=I/�F�����B�({ޒ��e��l��W�8�/S�v��j`���W��=|LN�Ww��l�3�����a�{�Y$T��h�oW���b
�FD�C�����o�I*��|"5{x�w��=.2F��C��aQ��TU&,��^�Y���Z�v_�n�~x���{Q�4���X�S2ӥ��0{�r�����u�/ո������A(�o�!��I�)1nT�b�9�pf�)XM�4�0X��{?zsV�=�I�n~�{_��������(S�w�+�<�ȧ�}$.��cMۃ^�~��;�iu�_LׄwL�R�����2ΐ,�C'���Kn�DT�D�c�L\�����`�``I��e��݋�����W.��b�l��A?~)�s�qu��
r>H���q���#eo0U�y�n:�ԕ7������Ϸ�`�j��w�>�����Gw�sϛ���9�*.au�B��Y6�v&��>���*�]��}����5���R"�0AE ����;_��o�U��~��������H�Da#��u��c��	9��Z������$qw�9Q�O����_�͉8���d6� �_ � ��*���b�qv�
f�fSу��qˮ*1�?@+Gs�9{埊�͢CfΜ��M����=�v�Ey�eh�C��3��'����V��T�lh��
y�q�cUXӾ���8�⚺�\����4P�3?}��h�7����t��x�:�nF���
���3�
��ۊ�l��Ǎ�\�n��1b�'���N�b�cV�3.�Pۋ͎�W��XǦ�oW��r� ���螓/wj;�V_W��K�U@��R��1�����!1W2U7܂��09�N���c�f^�dC�s��.+V*��c�
��	��@�*�U^y���;}Lk���P���"��KtU�?
���݌��������������a��:Ҭ*��X�k~�VYV\��6��Z[�~s�/'��r���ať�R������Apŕ��d:;W.�v���u�h�;_U��v����Q��Y�)S�s��w_�,4}^��)����)�P�0���EhJ����r�#{=h��.��R,��7n$D�ݷ�wиN�r>�>KD27�Ѧy������F��S��vQ�e�ѭz�J���vg?N�gk5�Y�g�`G_���)����4m�!��V�]��x
�X�uJ��_�Z�\.k�C�����xa�	%{ڶ�أ���_�-lImg����� k;E��i&���L�њ9�q��� NL3Qe8FP��ݹbN�t漥[B�L�ҺpJ��k�(���U��D7��ZC���Q��r�q�%k�DQڷ ��6�h0��^��%�דV-,*e�HIR�q�e��7�)f=��-�����M[��P�r�k�����2��Q<�3�ު��q�Hi���"
���]�����O�d�[�"�k1��w��=�[����/L����s�]tlz��25�ouи�K=�l�-Oѭf]NGVtL�ɻx�W�Q0 �g�6k�}sܪ+��{���8���D�mf����{�y���C�z��0fDع㋗�����C|��=����DD |>��Z:�@]��*�l��=�l�"yr^�99���^?�q�)��:?*w��~�]i���pN���>ߖj@�b@SW��K�"����ZfaSi�"�}��Ep��q�1g���/��y>� �J�`�A�&&Tb���lg��h�]�5���#^Ā@?�nUS��#�@��e�Z�]b��y��*�# )U���)H�0�"�
E���+D�, UI'&�����}(^*�"�RW'E��0ɝ��*���47Y�dr�==� S���5�C�3������*��@��j�(�,�̾�@��ͻ����
��\줪����猿h�~���w9q�HY�{q�<�u��2�Z~^ɬ|���;XN����dR����P�ֶ �8���*��v��>�/��B�ǆ��x�����]H.�t�������O��՞h����eI�A��8>�B v��#ɝ.������ڛ
�G���~}���*�����ZsqLy��\"�$����4C�P�ϯ#r�1�_Q?>ɢ��r��r��eJ�s�+�����q��gk����[v(��|�61D�=fb���Mq���,�C#m��>B\���F�bp&e킂�����F��|a�Y �C�{�p��P���ܭ���k��ַ���DDb�X**"��*2Ȱ�bȢ�
 �DUU�QX�#U\�.iB�`72;���:�K�I�Ns�D�1Ѹw+/�CW���(�CT��\�B�vguw{OS:��䴐�R[K�'m�"���^ם 6OI�;Ba��gHSW�\z3E:wu��,��6ʏ_��zw��vz����<�_�6<�lgU�&q|�ύ��#i�����@�F��5�*A*�ƺ���1]OϿ�  �2/��_��;v�U��*z灵��7�0lQ��7'�a"�G@����y�홷cgKq*�,�k�zh�&K��Ƕ����h��2����돰�T����q��:����n��4t�]b��4t�ڤ_��v��I���p�U�����#|35���cH(�R1���X�Y�<�׵�8���B � G���T4�c���:�N)��t������dWE�9kRwL��u����זd�h�I�W�}N�����n!��҆첟7���+�<<{�i��+���7#V�"s��t��t�����(��4�]�d�52����n��Ս^u��!#ȗ�v��pk��յ�F{���{�wc�|9{y����14L��x[�-g�bJv�ݶ��װt�<�D^*ݺ.��X�9���}��]w^���",o�<{[s�z�г*e�C������]#��}�5�Y�9�^�э֪]�b���:d�&
�KW�C]3��'�c��)ф�G��V'홾Q��}�{����S�~�8a��i�=N<.6;|{=gqs��N����
Jcٕ���=��f�ͺ�Vg�[s}=������dVA,"�2kZu�'�u��j�>�m�`0,Q��~�k3��oWg��yٽz�H��t��uq՛@��`}Z/��=�t:6j{>��ů�}ejLَ7L�;lT�r�VcipF�T$�_@��\*R���-�*P\�b����vms�
��:T��0��=�^1&�@���l�u.��wG�v�p����֟�����[`��q�^`�#�˱M��f"���#h�0���i�p�����)�����x�ʛ��/z�د�Ҭ���j����9�ō\�9�ԝ��v�;���wQ�(ç#<Χ0c�S�5��.�8u�נx�jr�f>�����=�޻n)����ZZ��R���	ɡp�����3��<�➃�_�J��z�=à�)_���8��O�b��h��15��Ʊʠm�<՝��ʒ�;1kq�M��2׻o��!wq�s�#���:�ri
�sSP�Bh�<��~J=E,X�AAQ�)#$b�5�����;,a�yM�;�w�AӲ������[{*���;��R���G¤��"��o�	�O=q$s�Ӿ�I!o�$�\�?Ƈ���枱���3�4�z9�9u�E�)�w��;�Q�g}��{�j���AZt�Z>��0���S]5&gu�`���ooN��Β�6�U�hu<�L��y�S���<rT-�[,������U����
���5WtWV17� �s�[��]܉b.��ZB�De������ﺩ<�  �",��\��Yn�)�TȺ�[����
��؟��.k���or��tA�(�s���6u!�{!��H܉Bte��'�䮥��+��f�zϐa`�1��lt�ٕ�3?nH�(Y[�E~�i�mĉ
Q���L_E�i��2��-	E��={7������U�w�t����Z��EX�(#�kOy\��ܨ�()�E�����Xl�(���1�gm�n9�\��T��E\���ղ���E��v�o��_d�E��^\��7�?g�#)N��
 ��ʮw�&��ۡG�4����f7�b�	��A����yp�hڥ��k�T�[�74Ս��<-c,�����o8Tt�A9����� ���,b5�_S��o;1��x^�Ϣ��eW1�����qJ>`k�.=@i��0+yf�W0�
���I�ףUr�ۓ��&bo��V���(���񾘥G�W	եp�NZ8?<�JmEO�7�Y.�\ݥz���{*� u�N�l��sVs-^Z�#6�X"�:��8:�$Y	շ�.�F�]�UD�����=��&OX�A�Wqj��RS7T$�$���s)�h���Ʋ�a�I���? ��z����aPM�d�)�C�F��ꚥv�na9�<�yyp^@^�¶
�豗�nѠ��c�E]�A^hn��ټ!i$�B�a&���rU�N�����ٓU�>�M˛[�.�Q�5<�e$�U�ITQRBE��@�J�s;�2��멻���\��I�̺���>O3>!@}�}�qR/:����+&�4Ff�q<eEwQ8#YVk�o������c���p�[%�ܜ7( m&��:�Q�W���ܐ�o瑋;�?���+��O=>��³hfJ�B:y�* ���uWv��r6������7������B<v���uJ\�V���ě�%Ծºr<�,�V���e��澴����;���jq�x�u����u�9�9}Y�T�ɛH�I�F�sV��w@�k�2���I�G���I$�m^�k��Sʂ�.����༮.�w;D�E@P�����u�GOP� ���n��ؒӭ�v�3�Z����R��Tv��j�o����ĩd;;�a���k�/�ӭ}��x��,l�̊�sz���V�jܡ��ǆ�G��\xQo�ٲ�n".^�3��|:#�H�/r�l{2m�>V���]���[�UA��S<cI�\̋s���PQVE����1f��!�3/y$����tv�=1��+����Ö�eA[)5%��MR���6պ��&��	� ��H�wս}S-�p��-l�*�Ux�g)L�`Y���4tV��ᛚ��h��*�F��n����%�5N�f����HП.K���_G0,
.4�Yo5Ș)&6����N|8��]��yg�P�}�s�g� .�KoY�NV،�X1��t٥tk9v֎x���K����T�Y����OY]v:/��e�`�G��N��u+������=[E�=?���Іq,�I�} �bqG%��I��mb�O��?A��&��<�^%�y�:dU��Ot��Ҩ�9dU��Z�ћ��ۤ�=�=��.<m� �0eKV��k
n���R�T���{7�)���S�
��g
���VZ��oZ��ySY��+�,>����^4��1�9��B��Χa�����Y��@}_}]P�o=��9������3��"1��
 �P4���~e�&������e���7dPL=6�&UF�p��F*⇏'6�c��\�+�E�\3�)� ��Z"�/�
��Ux��'eۃ`��v�4��e{7'�o�J��&B8MS=���1�k7��k��齃�9��݆���p��[�M��ֳMV�~މ���XӐ`��Pf86y�݊�y�M�q�~�x�
��܄�UZ�f�dv��)c�'�|�x{L�:'����8z��w�~���;o��n�!�8|/�}�n�p�"�6�i�?�ߔ�^n����K��[��%�,Ρu�j.F�י&�Ld�K��v�:�<���ST��o��
��*vi9{4�����~�8[�aKԸ>q�m�>N���6�\�'Sf]-��|�_�|ޯ�3�y��rb�( ��H[�[=wvҪ*�H�I���Zύw�U��w��W9���+"q���Tl��*|O��(u���'e�T�6b�T��i�F���:4Ʃ�}tǮiGUYc���h���Z��`��=��HC�';g{&�R�!�z�v��\0��oϘ�++���s-��̼�6q �d!�8����`��k5�%��k�2�\�f��q�nZp�s\��3s6�5��J��ol�sH�:5��K�jR)wMD�a*Q]��G[� (R�FbA&��($F�f�rd����a�hj�z1{�v�L��o���t]]u�A*FuP�ܣ��[-����6�����w����խ����H����ϵOo�m�����=���oD
�/*a�dj�,f�]Aw[�����Cf�}�l������q���,�ٳ���}s�d�K�L�n�bb_��2t­G��j|v*Q�k�J^��S��TL[��P��Ϫ�7���x��W7�Yb�Y�A`�QR2]w���3w�~��sZ�>��2�������ޗk\X����V��pN��$������)/�z���Af�_l��qJ�	W�N�V�&ev_�n�ͮu�����V���瀃$I�ʊ����6l\�z��
M�Vz^R�Ӽ%//f��#��Sk�g�D�G*�7ۚ�_4��;�C�q�\%,��~��!�1��K����x�N�y��l��o�LEQD����QB1�cTU�QY"��б��"��E
B�E	�fw{�t���w)��Gz`�-�1��s�P�i�t��3�r���!���^���Ծ�K�^T�L�_���P��f��q?����Z��C�='i���Q뷅��<7øz��ɎWg��N�:'ZXm\���O���1�#r��d���ڱK���z:W�2��O�uxY�ʌ���˺�k>35��)�Ŀ~W��:Kp��{�G������$e��:�v�k��,AA��EX���FW���{�+�b&�me�q�`��t=Ý#W�1��@�;T�wu�PCl"FC4�-�P8�z����s����`�&��z�n�������6���>�����H��l��j�x#lm`�蔟��vV�oŽk>�k�Ri�6�./�z��I��^]b$��G�~?O�/eb4��������}Y���"�οBaB����e������G� 	�}�b�*��|�p��.�vV13-��O�c'Z`����1�໋=��/7���>�ߝ�S"�-����j���=���mW�T�b��rn���<֋L��v7��2:�v�᱃Z��{�#Q�CϽ˽V�A�/�w~#�v罿C[����n��_���F�N���ש�E`�PQdDUA2����������k2���QѴT�ےzG����9�nl��{�-')nl�\�-�8�����w�?(j!��٦�7����"xkt�~�[`����p������/��'�gx
âwƺT+����*=B�܂����u�:�}4�_R�>d�F�f�[�'jw ��\C���>�!ařY��dp����܇���x�����]�1����;���!����(k�I���z`x?�\����^ʐ�B
~���Sˮ-z�TPw}�Il[;B1��o��6�9�MYbk����ǉ�{+�t�[&P��&�@��5���UB�	�h�*3Y�g7r�I��y7�O�Ͻ�߼��N[�v�,HǪ&׊���ו�$�����$���zz?r��[��ה2�����;)Q�1��A�Q���n�DNuG��r�}�S�wډ5q��!���<ck�YP:�\�ɝ�PQ�\�;�wU�K�Cٙ���8���O���C�-���pit�����i�ʜ�����$��Xw�*�Nn~�k-��`��IԤ�c��_���T̠*���O��w�YCEC�y����˽����$���9W}V�h��S�z�ō(f��ml�c0u�TcΨetz��xL_1���׼&6}b�`}�#�����l��Ү#z�	����������� �*�����nv#�&sѝLК�Z��yx͍�u�|��_���w��v���ưv��B�,��in���.f�khƵ�u��rO(�*�ԱY};"��EE�B��~xw�ϰ7(\n9pݦ�:�4s����~����9n��z�����諾��8��*B�93�'���Inf��`A�T��3��`n�L8����a�F8*���Kw�Ɂ~5���p�(�D�F(�;��Mf�Z�Y��̡�E�`��Ȍ��(��try�ё�>�JS�7E4��-mOja��N�� ��]�|����y�Pqi�p��R(��U�*����${O�����=�]����Dٜ�6�8��0��7];�a}t�"����9��ït��hu�3�:K��'ڽV�^ѯ~��ʬ�Ua�}�U�u�)�}�K_�=�§�l�#7A�$��UHShP��(�E�K�^��Z$j>�o���_���"��uNr�'�;�${0�I��"`B�����+K W�#�mV~PyU{]�Cܲṉ�:�Z9�j��"�����%����U�T�g��z^�.`�O�_p��a�,��
:Yٝ3G�ف�Ɂ[���ʾY����$#g�j`+f6NML�
�,2l�T�Jw�*��Gs]�}����D�ATA"�,b�E�*��
���	�A"�ϛ+���s��ζ?f�V�8S(�Gq:�
G���<%��-p�]�	f�m�-{��VW���XqvMR�)�n���3��"�dgy�B��N�-�ujB��80�n�O.��yv��8Bܺ��߯5�E�I�h������	@M|XT0U
L������u�?T�>��~�Bєg�k�������H��J�uaҢ��u�D�Ȏݢ�R[*��5��PH_�M]|�������o�j��]�7|�js��]�7|��{�*�6=�x����æ����n,8W>�T~�b΅�B�S����Ï㻮n��[9� 6�)"����g_KS�,jf
b!��Z�=���nߑ��;	��v��u[P�[u���m5���L����'<������{U���?<z��EJ��\+��~ "���E�D}���j40��폢 TG�}�	�#o��_
�����V�����G�����F�Tw��vO�
�[��y
z4�~C�DS[�'���9�M\:��vh:�h�z
P��CFK�(��@͚	�
1Iw�_^����}�i��u�H��r)0]�bF�c�QVCs�h������V0>�(( ��7S���<��7�֪?O0���w�<P���􏖭+,L򏖒��:��tOUn�gH�ʃ(X����sʫ��G�m�E������}]٢���W��Ĝ��,�y�������w���콂����'GV��c�ٚ�S �n�ޑ����띞�UVA�����^�=�/�=1,!bx�8m��>ʤQifM�If�or�j�ja�;zN��N���z����}ؙ�a�W�&@ �I {��M�"��QQ� +TUl��3�S�v,�q[�v��q0ws7��H68m2'��]�N�+��72(��B˪�?oJ�^��Y�.�uq�W���~E��\E�e׆TZ��{
ۨ�p?���nᖤ[NO
�UV�����?O\���R�vf��xn�,m7���	2Iq��Gg���^<�d+�HQ}��é)��}��]���n�~�~Ք�
���z�0^C�K}��p�,ד�i[�u���a���1�Ẋܧ�?2��~3n�ݪХ�����߾f�{���")��<�#����-s���w���� I	$�ā$$����		�$�	?�T$����!�� �脒 ,�L���S�Y$ ����g?�^$	!$���b@�I���	!$�����'������N������������� I	$I T!$R$'�����HI'���r$��r~�����HBI5�_�$	!$�$	!$���IHI'?��! 	! I?�_������ц��O��@�I����-B@�I�P�$$�����/�����n�HI%�������ā$$���I I	$�����d�Mf�bl^�~�A@���@ ܟ}��'{���@ QE��:t@t� h5A]�.�:+�m\wFlٕT�Ptֹ�A�S�l

'v��u@R�hH�IR��+ْ�cT*����**���F�$��B��� $* �*P��"td�%T��B��$T�*�(Q ��Z��ۭJǮwm�޵�]����gR�{����*��[��;�*Ѻ�	����{������u��G&�uB����ov�ۚ��^��W�+V���kR�z�*�    �]�   @�� �@(�� �{�N��]���ֵ��yd=n�����Qw�Sq{���5z�6���ݺ�����ר+cs���ٶ�=j�
� �f�� �{b�����]��/q���e���;y�T�q�ޏn��b�Ě������������]�����ݽi�x�-�EkT��V(
��
�leT���{q���&/{�:wj^&�z��Ӎ�����g��{�;z��-�{����ݮ�zv�^��s�/y��Q赸����k�[4��)�*(��PR#q����G�;ݷ���'v�w��x�{�{oG�ס���^��^��/]�^�\^�^��鮺��o;=���o\&�d���z������%"��"���g]�2t�60�]]��{�ɫ;{��ۄ�t+LGG���w���ʬ^m�V�1��祽�Ub�{hz4��𪔼ӧ9N�t) �4v<��w�=�j�qێw`&�W��iSWs��޹���[޼zw��xΎ&�9븼�F�=��m��q�=S��U�����bR��*vw'��V���=׀�Da��u���mRE.3w�:9oy�����<te��]�L;=��.:{�^8Ӎmn�++�&fl�$($ ���=��#F�޽��l8��A���`6�0{�q�P,.��rQ�w�:=L[Հ�{���������Ps���ʊ��%E�`��q��<@���
K�x��������]�wW�Q��a�`27y����l���TS�|U?��J�   "yJIT� h 2F �ɡ��j�����2`��O
J�d   j �!56@��L�'�����'��7����%��u��/&)sQ�q�9�]���N櫝�� $����$I.@�I�! I�$I*!��	 �O�D	 �K@�$��@$��
��{�������[���?vݺ��1�	�����l�fi���ëw��^E�6�4�c�ѭ]�@a��C�N���L�Yy{�&oe�x�;�][�y�U���ז+(�����7���Vq�f�<�]����+��i���@Qx%g��iAuiK��c8T����B�	0���r�i���X�ӫ�)B}��=�Ӭ�yq�*ÓP&)����ъ0�xf؛��7|�\�)Fv�{6�*ܭwxiei�ۭ4[ʅ@�`r�+rְ�Rn
�%)غ��GP�Tj��n�{A�Y�ܶeYyt�L��=iLiԔV/O���{)���N�,��w�f�� eD�u3o4�&�	V�umm��AP#@^5�i�A��E�|��%����U�Zn4�4�)�!f��Z�	���K�1�F�6��waM�ѡz
dT���;�6VX�t�1%�(R�sr�^�8Pd
�
�XK�
�b��i��[�yܼy�Q��h�Yy�yz�-uj,fάGj��l�j]G[�5�{W�[��_���Փ�mۦ�������3[�e�l8�eй�N��qٺ/X+K���6��C���PEQ�����=�ݘ�jƗ�i7.��6�ve;՗7I��#5�
��0
̪{��E��)V��7pͻǔ���{(����E��������$������pI��}�kp��D(�WMMYF��T�Afբ@U-r�+4e�:�#�pvH��J���6{ۖ��&U�2M���+�n�dV�9������H����(I
�Z�U�zKe#^=�J�׹Z���BЬ;V�F��n�6�'�mmk��^����)��@����YLT����!�p��,�YԖ��r���r��e]I��9��n�������t�N��L("uR'l$��ٖ��SC4ӴV<�)ҳ7Xou�c-"��n���ò�<F[�[���Z��٦�d��Xd�u�e�n)�V�kv��Nʅ-9�
�$ڽ��hӸ�ۡw6�KM�y�
��$x�����e�33\���T*We�oL���L�o��K�U�yFf<��5f����T�u�4*��*���!s|��pQ"��fK-ۚ�-QŏM�L��Ud��r��'PB�^P�M�k5�cMZy5�6�"�r�COk���eXKw{�¨�YFEf�
�3v��`nz�Yx���{hi6W�^;j�����L#ks)�0�oKDmՠ)�E�$��"���Pnޘíݣ�5�QMZ�a-ȅ\ub��9f�[F@�Pp,
�k���#Y4��A�cQ�+Չ�$��qG�*�<�e�)�,�u��+ob�N�r�aFu���#�Q���u�$F�$�{{V^4mZ8�5y
�]e<���Z�Ljڒ��<d+�֖M����1d���MJ
mC�Kg-W�P~a��	�ӫ"bR/*e�3.D��V��{��A��m;�a7t���92�6���޺��n�.E�mg��Ą�
�����`!�8{f�n�6��ARf��7GP�����d�o �bֲ��7Oe��n$K7�5Z�FЉ�F�/n��h^jH]�cG}��ʛ�XwXr�6�d[�ܬq`Ur�Ng�]����ǥ)>���.�i�e���Q��{f�4��e����+[� �d���{���sB9w�ӽpT�rm�b%�*Ą-'7�o6����Эow٦��Y�o:w7!��M��5�fxSe9�n��fmo�Hf����4����u�6��4)�{tJ��ݬ��ͭ�Bl)�6pVL���f��2��@�y����n��tV�n�,xi[��L�l�����n�ܲ,��v/um�B�b̭�SDyv	y��c+�n���{I��\Ѹlє2�n	�H�L��zY��-��U��#tfFU�P5gΐ�\��`Zi�h�<�N�Tm�2�J�&M��V6��Is6�o5iZ:�x�������Zn�%Mǒ^U�{�[�x�yH6�\�[�ڌ�E��n�2U��B	�Sx�N��2��M����� ��b��ט���WB+[�֤��!WJ7�){*衅��1�KM̷�@ڼ���La��u�d9�6�V�PX�mؖ̒��h�RДA��v�g��+7/4�z�Rc��a�ZSl�f�7<�8C��z�p\�;�W�Y����v��[w35�6آr�YR�P�Fܶq�*Q�d�J��v��j
�hv#��7�q<�ٕ��X�D�5��6K̘�t�������Vrl@%d�H��ĳO"��j+�G�ԕ�x6�(G���a݅F�U��>4����U�+-�(&�i[)`uv��#�J�ǎMƬ��[6�ݬv�3gvEz売���j��,�0h��_kRk]Ү:j�=4i,�͢]ûI�3�;A{K�l��w��#*J$�9B��Хf5@٧"�5�lAx4�vТq�)�4JB��?m1E+6�]b6@Z�6��Y�Υjf���w����ݫ���n᭘�C�1 x�����Ve[ۨ�fbs+r�-��Y�b�duy�=���I�m5�/jL2��ɘ����	5��:��*���{��ۢ�nfl%�V(#�z����2�mݍg06K�(�C3L� 
��qnq�[demd�WWn��Ĝ�{�H�e[��L�N�h�F��
B�t�U�*頥�Q��Ò�x���Q,���໽�b��`nR(���r0����f�5W5e���JƥE1�[�41��3[iҊ&��	R�H`�+<�ւ�|���/3+oqB]*ԅ������f�`�Ȃ[	M���1ѭz�m�+�h�%B��FTA�r%K�FA��*���ae�Ձ	ٖN�#Y{�EJL([��&���jκ������8����6��-]WSF�k~�Gi�]�e0(�ɢ��Wx��5Ţ~#���m�Qd��᭔�Hȵ�V�Y�r��.x(�v������ar���E��5�5����%oZ:v��[	nm�5��#x�df�|׶�I붝��GN�a*�M�pXɨ� ,�Y-Ҭ��t�$���̢	����6��y����^���[�2�r�ɲ^�
���4���U+/0�k_���4�^ø������!��~�B��[f�9�񾱤�*o���mU������lɨLaSu{.Y�� �bw�*� ��u\��^��Vh֌[~������
�+J�M��\�gU�L��� ��K�7H�R�
��
�X
�	f٪�!T	�^z�"�Jc�7*�oi�j�����|F�x{Y��*�(�)��d����B������N�D �Y�ѓ2`��2�,�ä���2T�	�U��"�"� W�
��ص�Y���vZ� ���5��7J��z�(����LHMӌ�}�6q�N�[�(h��^,Uo{L�V��IО�1m�Go��9.��kV�\(��2�V�V�ͫ�aUK.��#�A��ti��ܧ��[��uz���o��Z����V8�f�"���7�f�kZ���	��F#7�8j-y@P2S`���2��&@� ^�cI�btFn��h:76�
�6&Ò� *�LM9T�J�.�xP<�/��f�lDPTH�W���V�x��ma֘�!�g	6�jfͷ�'%�1t��Ǚ��@!'LF	��K4���[�Nج�ugU��MT�U�-h��(���I$��v�������Rf�����4B�v�MH����@���%�h��w!H�����[XKW�hFt�,:�{GV* 余�a�
Vժ�3*�)�ۭ8���<�5˚�p��+�͎
�T R��1��FYys���d��� �V�$�"$��-��\�^<T��D�E9��i
����"��\/N1���T�X�p���wyuz�P��H�Ӊ�|�"���5!�U-Ihz��N��m��=هMe󽴬�#��8Vl��
̻1����p�+E��2c�3zux��7,Q��(Q��en����Ap݉[�+4AP�%D�<�.����T�.h9��p�`h�cMi��h�TKth��iˢ0��o�C�n�}i���mg
�d��[M�7~��F�K�S��ut6]�ݯ!�D��;��T`�5����
	�������y�KS%���{��#��*T�g[�F��Z��ĞZ�G��r~u��T�ݪ�� ���b�z֜`3�Y��������W7��n�9�����+n���݁wS\Š��t��[�T�Ե;�::�ZҞ4�����&�mR���b��(��*^�-o+�n^^�U�
eP��C=(,�VB���Hg)��h�vlEow��7w(j�tFVK��D��E@�y��B�R��/�n��|����&D/��*#Uu��l+�#p]o������oq�UW�CƅM9��7E,�2ݗ�t�gw;�˚�l-t�Sd8���R�0�T9OF�45Xq�i3Q���q͊�N_�[z��+j�T�����D��e�Luh���SEf��kj*ҬIf�ט�jj�5�sH%��u,��Mѕ��n	EY�VM,�v1�cG-��6��~��K*�U` w��R%�V��K���@X[��ݍ\�XTjl��w���]�//R�4�X��u㨶��#j���
.��t��V����1��r�n���2&՗�v�<`�(�*�
N�e�!"tʹ�ʬ��,�W�Yd����"�j$m�3pf�L�[QY*y2.�
7	+2��t�����u�G,z����^:�,�V��MF�
�ae^������un�Kx�u�=D�VhZĀ�T�W��T6�7�!)]P��L�P%�J.a�a�t
hM	K	˄���V��mMB��:3l֡[2�k|F	�"u�)��1C�^x�g_S˭�������`n�OM�	���x��]	L׮Ң�9��@���,a}X�%4M���>FEb�ђ�@C��E6���@G"nє�1��8(���W�ލ���ʼ`kMZ�û����s6�U���T��/I��*J$�Vk�X\9���X+By!�ƳO��Z�])ĩ�)��2���8������&�	 �#��kӻr�j������!J]��At1&ԙZ��0�2�bj�,\�R�&[��(1D6 �#"$F]P�1Z;v����u�b�%2n@�݈#���Ȣ��ST����9��f����Gu��8�ꪊ��1�""%�W*�G�F����3Y�.��B���r�г�a[�2����;�ZǾ�m�h�I����*�ڃ%����}w��An��J��{6�����+Nܥ�lef�˅b����F*�ɶ�Je�J�JA
f[j�50��X܇^Lmm͕�h�*����ʵ��ml܎�
�~&��Y�a��J��֭ˊ���z5��g���/2e%�m$NM�Wyh�冣�G,�
RQXI�7��L�[��J�ݬ,��Ơ�-�'��ݔ��ã b�5NY@�6�16��bn�sEQBr�Ȁ�5����E��{MŐ�W("Z�o^	a`v��D��Ef��:���7fۻ� ��n�$��U�[�v���w����-,+�(����`Ulҹ�RVy$�4�׃#��2�6��.� *	b��oҧa��0eʙn�Z�T�/rδ)Z�<̽�Sf��fƸ��Ӧ�Y��T6����ySNF̼Z\�be�]�*�
�`ɸ�$R�f��ݱ�sI��Ֆ	����!S*��4mQ�ݬ�tхeu��DG8r�m�Já�����׼�*�n�u�O���>bͫY%؍jF� 5k�oE�w����l���Z���6l�]�pl�Շ5[T�+��u����Ih��xP+\��7�i�X0�/C.��̳�oq�n���e������l"��,�U��T��;ow4�6u݋L2�ম�]�u�޷�p(� ���[5�T�n髼�6rnD�|�2��h�����i4�t�ֺkp�t�/%[Yj���Cx��G2;�X�]C+C�c�Rb�Oc�pM��Am+&���6�]�{��9*���LDi��U%�h�j�X��ќs���`�D���a+sS*]aw���m��o}Z(�Ͻ����V
�˭������E��Ee\Kb�w�#gU	��cn�]�1��4��w�;l�a�P[�B�k)�YUMn�-��l���X�������S톯����C�n�O�BDJ�x��ҷ��Ymk�]Սw�]�0��w[C�ԩz�x����j�z�������oP� ��U��[�O �c�ZZMo�l੬(��70@�ݵ�d�F\��ŋ8�MÖ[�q@�t*UBqa��3�I627Q�\&:p�˻�����ܒ	n�-\w/[�/C�^�2�0�G�6n��y��L=u�t4�A3yG	�����6ҎV/6��mj4VS�xPf(,x����ZkJl�uZt�c�\�"�]r�5���U��)!�%-cf��� �A���=������ܖ��m�)��5�)d���8v�z�0��WUo1�Vb���Ɖ��©�[�d:B�C6�fn�a�P�.e� e�=���k@��N^S��1V��j��3l��, Y���Z�K{)�����͌���J�cCUU���λ��d��Z�OI�,�_��͐�\Y%����A�̃�����z�.��R�j��Z�g�0�"�j-ب,2�b�\+k6��vaњUA��X�.�<r�8s&J��xr=�)��;OՂ�ҭK
�sua\6�\��wz�f��W&� ��s[�}�R�պ�-#*5��K��De�ث_r'1IdJ�v��y�ɽP�}�f8�_3wt�ֱ�]$�1c��Ÿ&�2�I[ӻ��ed�.�t</Z�c#*YkGyk�ɜ�r9|�1��ØV���R�m��c�}���*D .m�-�έXcs�=@&NV!eYZ�Y����9��d[�K��7�ݡŸ�zfX��m9���U�;3$6�\�|�TC�aֳ!X7$��ӟ��n��Ǹ6�q��+���nV�zz�_䓔솝��9���ն���,+78�:���7�n��۵ܚ��M�B<x�[!��sU�6G+}!����v�L�m�aJ� 9��[ջw֗hf�rI;�AmofN���]�e�G�#1�Wɫ7(�7xd�c�;����)��\�!t5ض;"�'�{�]D��C%,~tG
7nM^�����inl��m���ȷ2t�{��[��D�ݓ�inĹ�&�Iwt���b\ܒNIn�>o��B=WP���m����-�|�&��ũ,[㥙I���(yZW|M��
����ö�Z!�w�St�I��'e��h�J^�G5�R��*e�����Q\�l N����Xp���W�Y�oD�A���o�����դ�;fu_
f�gF�ZR�<�wan7�6�^1;״�IS.$s����������YR�;ۜ�ܜA2-��*��Z3��7Q^���V#(%��m�$)���A�xz��E��[a��o\u���\�>4�X�:攛���v��Lʧ|�8u�����n�^x[���oN��'_T�6龻i5-�㪜ի�V��d&$!T�u'�l���ַI��Ye�����m�Ԁ��o���M�m�Nܮ�!��PېmN ❹[��u��̢'fd�ku&���E�E���rƮ�l8�.�K�˹�s)8�-{gdx��2�tZ��I�7�t�-�@u�1��b��wD�������c�@�%���ɈU��f��U;���O�1������zv���\�;=Ȳ�H�9�-�Vҭ��^�x�Ĝ�e��W&�yl�;n�����]��y)��P�
ܛ6]	73�r� �˚��v;����J]�t��%��RK�ـ�`�Ŋ]�W���J��:c;h�׶FPæI��	C3�R\�{`4ˏ!*zB��w;�e���D�X�P��x*et�$��+*��ֈH)�vM�Q�5�J��Ǖ65gz��Ԙ��QKk��E�c��s�G�+����z���y+L�KBG�k��ZX�ݾ���l�+�5��[�LT'��C�h������J+��:e��z�2*��h��*�$4�[F�H%�s�rA�w���P�pX����	�l�q��t�>�۹�B���	���E�>"��6U�8M��)Ze�m.o��#}$�4���jְ�^��X��f���wX�׵�=�'���u�ͦ��Nգ�!|��(���i����f�HK�E�.���5�\���0��আ\R�v��BT�ٷvt������V�.�;ͥ�޹Cb����Ɠ�{+ebڱ0��ۂ��c��6������ٟn1���=��X�a��95�W6j�y{�3i��Ԁ���Y2��o86�cѠ\��[*�r�y7Bs$�]�"��L�ڻ�'�w��^��WCR���&�N�
R"�kE�
T9e���h}�� ��s�wI��[8U,E��o���&��RIn�i��A�u���Χ7N����\=m�Ȝs%ޥIQ@�bd=uW�3�OI��iwI#�1��M�\��.��ir[Z�Z�y�e���P�vi&P����KĘuʜzXt����f^p�3G���;AM���nd��j�Č�9l-^;ݫkFj�EG���=0v����ƖR�g��{u�*�Ȳ���ƪ�dGnw:;x�����=�i�[�&����9ck&��oiq�L���Ye����X|��>��xb���e�G��r�;�Lk���tȭ�`�
pqf�/�yש�TO΋�|M�Ϻ��h�-�-JW���	uy7U�??��3G�;����G��K�>�[��ۨ8��3���oW��G �7�H"Ħ�]�Z��m�޼�͂�U.f��D�żK�:u��Uls���e���Q�d*Gs$�G���dD�t�n����z\cfgM��&9}ݑ�`���L��u��Gt��
�&����,z�7��-�YJ����:o*���ADM�V�0A���>r�6�Y�� �l�ӏE*���l��gUޚЦW^��]2r0�N8&�ك]%�o��|���q\	u��iqr��6�w�ܾC��9�|�0#R�]�鲞1U�.�+6���pΫ��ԛ��0<V��(�֙�Z��67�E%�n�L��4��=��_J��Raa:Vhf��,:w�n�*�@�i�ލ���Uw&����0���Ө�2���-��/v�V�뜛�ou��#�$�$�])f�^��,�Іz:�jz90鶺d�X:�,e��rh��D��5;�I#}"\ր���6�o<�3�v>�G�siPj��2�c|Ɋc��Ż[�!���6��G	q70r�Ue�q�b����GH�5k�Q귷|�:5���)���;�J��]�Y^:i; �O��@EXTƈ�����]G�0��z{�18����vn�;�=-ʓ$�cb<��}#��y����ݹ�f���ˉ��{�{[��FrGn݇�A:��D��e�;��Q�ʅ��ji3�!{�Φ���p�We�wl	q�.� ��X��{l)u��&��0L�ӵ��n�6���j��e�Ls��
vλ��v��.7z/M8�9/M�nze�D�f�J�Som�9m5�)���n]�u,��a˭���j���l78�e^MY�{o���un���ٻC��{�,6��m�Q֢�!�n,�^f-�t햹$�V�J"���m<�S���h���,��k�'������<��gJ�J	I��Ʌ�fw=�ئ�[˒�Gne�tj����G[�i]�w�����B�����6��8�y���	��i��൵����Lc���v�^�(�E�e���[y[k����	�{�.�N̢w�B#I�����!rk�X�3������*
�s#C�;��LBb��y'N��,��ڣs��0EeGu��el�S�#�z��������'�Đq�M����K��qX��GAi�+h,�[�0c��+���7c9+1Nn`l�;���N�cM.�ڵnʱ]������Q�U�R��7�ZN�]��`[|�c��e��:�zF�c(�6�Q���<�d"ʷ�4]Z�/)�Xl��J���)�ѱL�{^ʄr�&ޗ-],�W�R���C��W!ur�%\'��0|+M�`Ƿj��}#�@��U�B�xt��q�Qqs[V����ʘ�H�D�R���t���n�^�7[�c��.)q�Pn���(e����Y�>F$=�/]r��/5�F:����:�F�Xo�:�*Rv9�f���Sq
��;MY�ѡ�Z���=6�|.Ć��3V;��4�hr��Q���a��Seuh�Z��V�ﯧ&�>�Zzyݶ��;�d��`�s�Ü��vp�0/�+�!˾f�,`b�K���Eu˰Ƒ'o@��F�˼��.J��ފe�CsVT��[umlC��!���@[����P�[絨��Ñ�WE\�23tB������K�Һ���Du�u:[o����@a>�;
�`�\�A��n��;5>�UE=ͣX�$c�-�p��A���_*�5Y��-H���3n��6:�Ю5��de@g^��2��!Ӛj��M�v�E�����*�P�Z�띠ѭg%��X��UŁ�5k�ijO\�D�	wW{��D�e\��6�tf�}�%\��]"��M�Eu�m�ٶ�w�ZG5�&�쭽�Ħ�����i��"���'U-{�k��S��d˲;r�i&��x��'z�(�"vggg��-�����n�˥�{V��9�i9Z�m�jf�4r�m������1r[B=4�c�wzA��۵�W0̊�/ko7-�m'�邶�N�EIf�ז��ʙJ[֞�i�l��p���n�P���xU��("X��%�ܽ�`�<��'s���#f�jp�V{���ė1eu(xZɷ:����e���B�b�¬��;7��d�]3�	[(*,����4�G h�^�{1�5��5��vB��B����E�L$-��ٷn�j}0]��
��jZ�;6����\Yv��,��+I���(�+��b���1:Y��h�`sm��}Sz�+ݭ#�{wzঞ�ZӶh�[��;V����t�t�j7�/�2�n��Z�wthS��˼�^U�ʓy�@�n[��3�s�:�0���[{�a�oc�ZYh�w5S�[6����sw_N[חT�G��NV[靫vR3l�2���l����C�lnIŖ�_jF�4y�1���fn����K��8�-��eʓ�+U�ѱ��Ss�|���ؾ{x����:��\یPڼ��͜�,�_N�J�yzr7#��)R�VH�rv#�K/:�7�<��麪>�'IN���EXWp�6�#����6=�dghi̻��}� ���4��h�3��T���׋d������"�G�����V���f
	�;Ȧۆ���:�DdwCn�6)3p�Z���o-V��]*�����]l�:��6�^@�0�K�/��UY\��t��m���-�"�;�h��d�'�'Y���{e�8��c��k�r�(F�D�j��Vb�7p�o�S���C����C�ţ2b��ݗr�ȭ�y=�;Odu�e�ɷ�V�F]_:z+\�;F��"ќ�;�X\����΅)�zc'����ыo��;cR�&GlqD�Lu8Lt�V�������V�[�۰ъȗ�q�˲�����A�F��޸f��5��'[�$!��5�J���"�5�:^ݱW&��yq�t��w*���kf,*'b���VSe(�S�eKx���%d.N�ݽ[���wu�,���k�@���u֌,QŚ2�XQ�)�[F����먡ʊ;\;vP�B��sF�OYd��.���ݫ�x��M��\Z�Ÿ�n��{0�<��r��^Vp�L�X�����bVBap�.�[([��yl��A[�w�i�����Xʷ[�;br'�H��:i���Kzjٚ��*:u�=���T�!���neZ�7o��pR�T���mi#')f�շUb��^�[�-��Ʋ[/l ��uEF�ŏyV�{H_�PKv:�^b��ZLٶ-t�j^r��$��՗�&I��̽�B�*��k|�l���J=M/����xX�\6�7PT�;�L�V��i��*(�*���oH�z����NQ��J�u�1��Fu�8c29Y�u���9�+�סN��k]�&[�i���[�����&�Nt ��(���s.�㻳�G��V���Xޥ���NWC����E�aVv��9w�ӝ8efDrJl��i��]y4����i��}V^�L�̸q�.�Yǁ���hmP�-ie$(]Y�¥	����ͷ�����dם�;�p�,��t�Ҙ�5���I9��jXӹK���8ܗt��,$�x��Z�N7Y��wdU��ȭ�.�
��-�`�E4�v�؀7֚�s&����M �'u(��i��Z&��v�0�4ok6�rX��Oo_��W�u)�]�V�Q�Iq��g��Z�̐n%�r��{��.�ӎ��8n!@��Va�<�6KШ,K�G۴�ِR�c�r���Į�Uθ� @��쀽�z��o�U��������!�Xu(��C��&��\��ȶ�ܳչX�D��34�K�c���,0rP��6���l���&jG��b�V�R\��2ڠe�����T�F�����	i3//$1Mǹ�%��fr�܂���vպ\+Uv$��=�vj��{�����8�rtg��Bu̥���Yu�k�gev����R�-�
����\�Ŏ�\-�Zḝ�j�ͺ���iQ��_s�7U�V��RZ)�n��]�G�%��=e��`�]]���]��ܫ>b5:��N��3y�j�WT��؅�yz(��F�O(�7��o�qB���8cf�#����]\(�#E�y�kz�ANΖ�>�H���}���!qS�*�	\���ӳ��n#�����y��/8\�]�9b��:�h���g1��yq��YW2�%ҭ�V-{e�wR�WF!h���u^�OD͖�X_����2�КE n�s�8����TP���G@��Y&U�8�P�Ro��56�i�͙z��_DX� �F4ಶ��eȔ�j��t�Sq[��ܻo4�\�n�m ��z���wt�%����S�o.�V�Ԃ�y�X�]�!�Hq���t��5\���w�MYSRC�j���덹��ڝٰ)'VJ6�V��d�/c����ַ�������,sxff3�xb��iԊ���IR�=�q���������E�wy�pd�dR�eI�FT��E�SB��Zu������e��zw��^��9�H$�Nn��D�f0�(90��I�����FӸj��5т�8Q9��kR.n�c= vs[ۋw��TӤ��֓���+��e&�I�F�"����s&�ۋ�;6N��7*՜�ҝJ��z�vi����5�@nǴ.�m=��|˹{��:<3"�:\����l��`)2��ȋ����� 3[�-�ܳ�b��Զ�����A��ە�n�e�0��S�����50���/k-�,�uJ��bK]��1��N���)��p�u��+�(�sB�+��et�bX�L���1�⹠�ߊwZ�;5��t�Řtʺ��)�g���̤��䠮�M*��Y��͌h���0��.��V�cW"D���Y�}� �ƜWWn:�K�N+�Bub�j��Co� �y�킂X����t�����j��ܞM�in��LTo�X�u`J6�- �$�*�� ��>��� I��B@$�I�&���	&�� � B�!) (I$�a	 )��$%$ @)	$����l X	I P	HB�$�RqD$�Bl�
KBH� � �(@�	hI%$!0 - 	<�X	4�$!�I� �B@�e
�� I���?O/��^q��4j��&�/�3���B^�':�:��Q�]��^�3t�S����'w$�vl�s;&��L�sF�xJ��L҃R+<��Γ���Eip�j����v5D�z�t�V���13|p���N,Ӻ���)inuΎ���4�g/��V�3QZ���wƤ�$֍�,OD"�ި��o�*�{�M��t]7�{2���U�C@h)�9�Iх���A�u���׿A��e*�e�(���c�E(��|K�U��nG�+�э� 9:ׅh�A�j�s�c\.��G��p���q=7��/�ټ��H�__$c����A�h����J��%�T��L�Δ̭�wpv�u�s�Izbl�*P�Cf��)W���#˭���8�쉇���D��1�6f�N�6�MQ��瘤��^T��%����y�1�ݭ�b�Nz{x�+��)�5W-޺l��N���읢��Rʴc&mr�[Z�Bfw��2X��r�ev�E��r�5v�j�ù�Rdн�&v��o�Á��\�� ��"럳��n�::K*"�.
�M��ΞΓ��ܭ�47��K�o���T��d�6ʱ��&���R�{�-Aձ퉯y�n룐of���ybߓ5v�1��>��ݼеtٝ��Сfq�mQ���.���0n��h\�҈�x@.���-��Y<-rJ`��٭Wvs��M���  $�$�ѮV;��r�}�ܚnA-Z���	�+uٮաSz]�����̹��Y����kl0��s��X\�|lm���W!z�W�.��\�o����B-n<x)���0���T�LD{���;�*�����R�OW�	Wh�WE� n�h�5J s��,�-���}\�Ʃ�ǂ�g�l%w�V�6�e�4�K�G���k���<ԩ�@^�<7��z��ѣ�=��\j�
�	h�W�2���:��D`];=a�q;��e	}}�U^ P��2$`��Js�`�+C�r;q��Z��@��a5{�U�Վf�j��{ư���CZ�d��r'eT�`7�*"dC&�b��7ʤ����rQ�$�gv�K�*�)�KR��`�N'�������9n[2l�r�B�p�[�Gu� ��n���{q�fc�RݻT��,���"�
u�n�c�/���0�ꮭ��9�PQ���H�Q"I22"(��0�	I�&t�G!1;���&OJ��]Uw���$� ,PX��o���s�sOD�	�i:�Y������J�oC�F�t��q��u�R�#'1RG1T]R^Hu-c�(�{m���
�{/if5{�,̍�Ǡ:�R��S��o���}w�.�� ݸWcM+B����Ǐj���\f%�MV�I#SF�i*�QJ�ǋ�)�m�[�v>���y���4Sb��q�EL:$Rf��{�r,�\���(��#w��b�y;r�]�:#�d#cpj#���^�@
"��7�W.�����g4�"�}�fZ��5h��F6 	�U��Z�"��ӝ��t'�,� �a5��@����m�s=��9�dy��ꋀ�WU�e�0x[<�γL1�
��r�nc8����7o�wL
�%RYb��� 2�\ⴊ%�44K]w_a�ʸ��m�3��-!��w���4�%�}e��R�^��dS��ȵ��u"�� �FBD#�¨{�wvL�ӥ�#�F�b�_.dB�Ct�լ�!VsNf�P��N��d ���h��n��9kX��cR���Y2��Ùf�Չ�&2�
��<���,���o�ֽy��M�v��/ɒ���Ado�[ܧd/+�(� �@L�¤���E3����z���l��׍��i
vl=�� X��cJ���2v��a�H��׍>�z��r����|ߴVqzH�9�%J4tD|�M��5��e�����*U޺��������8윝;t��Q�������O�l}9B�(փ����3v�'� nX�� �a��\����s.��׍ZJ��H����l��ש�\";}ȟq%�]�=�W��- ���j��vfZmf;���p �p�h
�g\s��{� a�r��`�E�\�X��j�s˺��st��+��E���E��AF �"�X�ID�sY�{�o�ݹ���$��A����0_s�>�j�*�Hs�&���=�t�J3\��5�5#�W����UU�b�G��h=��*so'$9�yȹ�x�gP"J�d�*h�XL�������R5ki��Y3�R\o\6��/r���G8�SM��>G�.��t��t�Aج0 ,k� 鎮5QET;z\�GN���\���r4�Лj�J!��@D:�#9V��Y��z]���븧B��,s��'�4(v�1��GB=^�*��2DDd��_�'�|�0f�c�DȪ��UZ�B�e�&��:�7 �v*q��<�z�JΜ��K�n�y#�;N��]�5%t1U�-=i�:g7o'Np���z�ߡ����9u���{+�ֱ�����Є��y�
��ȢRѮ��6�"r��ܶ6�.�=���]W�����hE"�� �DQ �Y_k�����]u����7x�P�� t�؂" �ye�Q=��W�^�	����\��òɩ��Uu��a����2��
�	���#��@:��S��`���+��J���ɏ��F�P�W��cf+��X�K`a����츽���_wPqF���t�#[�otey���)�M����Mr�����J��y�u��j���ku��u練����>�oUj& s0�� �6�W�
�\J�t��IĕŊՓ�	'\їL F	ư�iG����Ӷ������m?z�������qL��.�m�|�[���f�(�k:t׆�[�P��voYB�˵t�"P5R�Z�"���ʐ;���빛:V��g�l�]���ou����J�C�G�0�N0"9{h��8+r��[�t����a<K�Q���,���;O��5�vAk1ԋJ���;�nS��cujR��i)R�� jg� dU�\�h�2Fd1�`��X##$�0�H�ŀB��9��K�u�h)m�� �,�]*!Q�'+_&��@gSJU��YZ)v4ܺ�LE.���}%���f�DN���M]����0��	g[g�2FB�4�X�t9�wy����\J��U��e (H(UI�T�@W���^�v��#0}������'���΁,�֨u�{=2{n,�l�M�����\�n�n��l]�H�մ0SǉlQ]���7��z���}��],z�]h��m�ŀ�ǐ�([:#�4�8�<]�;%
�Jv8����ע��0X(Dd�V+&~���ַ�/��Y`k��[E�i��|�,�.{Cs�m��Y4q��ە��۞�RK8[����o��>�uk�z�V�(��;� ��d�� {����7�o�����46F��{f�Q�q�;J�!V����M:�����C�N�J�B2˥Yr/��jK��4�Bhhe�������X!(�
 	�X�@E� Y)##Pk\���f�����[�+�N`�#@ABd��&�I��X����*�*>HN���oe���*�X���'�Z�x\��ө� �Us±h���0S����.�6
:+��3.����^�严@TVL�$��~\���f��Ե�h�Wt�L��#��f_m|���V���K���Iܷy�$�d��S!R �E����{�｣nu����
΢�LP�tصݝ�������x�g�E1���C�5Ӟ5�,
]�X��wl�E.�m�e��W,c+�ʹOMd�3z�$5X�3��I!\{���P����kvMw=涫�Ѐ��GX�VwD0�����x��F��&}�������y��YԀ��s� �&k���2qu�y�wW-�ͽY����1�In�D��:��#�YEf%i��x@�o];m弝SS���`���k��.�/�����rף��d��<�1�C"#�Ab,dcAXA�#T`"
� Bm&�yE˔Q��{kn�
�sg,	�u�H�o�iw^�s�_=H��~�hg�^H��%�b0=�5�e���d�'WJ\��ڈj�5&
K�Wt)��HS���&Vc(�idδKo������U
�{�&"���/�.鑭�Γa����5	�wQ��$�Y;/�_9�R�v9K�.��HL���n�o�ҚvGl �r^��������SuL`�T�EX򂣌��b"�(�TP��*�Ue��-^�Z�ǵ�5vV��h��z��opDd��j� ����X�8�rp�p4�ɾ���-G�U|�v�D�ws\R��gGڞ^]p���p�ު�S���GH��'�����w����ǋ�
m[� �@St�:J�]�BqPWYJ*#R3�vcI��`�ݾ�L�1@q"=O[�1-k�,ӏ�N���Unh9���o\���@HQB��0� p�]�j͋�A�*��5����G�AR�ؤI�)�),���]u�!��aE,U�D�(@�PTX��B,X�DQTX�c#��W�y�Q`�"���Ȍc #d"�E"�2(&}�Ͻ%C�l��zE�冀xiM� �2��wLJ����$qu��8�K;1���V��{l����"\�G   ��m��d��a�}^�����{�mq=�!\M�[����[��Nޝ;.l�T�e5m��2�!].�b��HD��eǗb���G�X��8f���y�21��DTH`Z<< ����Yέ���X+lǇ��ޯzaT�=W�xM�no^���s��Wq�q͔H��r�[WlN�,��|qGI|�̢mf��ڢ���������뷵�%��w3D&^݂�v�p"���K���0�B�:8�S3-�./!���j��Ž!Flv��?�����S�c?�U�ߺ��]�=YbNC�R��ZC�q�ʛ�(�B�uQuϗ_v�e�q�}�k!�Tk��Գ,���Mq���ȫ ��� ��DI)�w��{�o��/��!HDǉ'{��}K��S�4�nVW��8�����������֢M`5�G:�>5T#��,HX޼�h��&
jK�yd���<$I �qČ_W���m�,�wQ�q,�h泿^��]�pi+v��>Y.��q/ىc�K[�;��]�EW'9ǝ�>�	={���Lw�+�v���OMX <=~��<R0������%��&o$ғ�AS-Dm-n%E���y���8^n�Ӯ��^�� ����u�����4\�ٌ�����59�&v;cF�=�_v�e-j��aN7+:�]Ī��r.c�����Pm��Ӗ���R��[t�U�F�[�l��C7��9tp�bhM�����?.W����D��F�JMk54�j�&[Z���*.��hB�����˔�V��[�ot7D ���{�����}X#0Qcd���Q�,�, �0"4(u��W)���[��:G`vg]�ȭ���)��9�����f�s6k��ծ0B���V99�e*����m,����p{@f�����,d�-��2|�+�jlUĔ�P���ݝn�ee�����񥋸�ME��������݉�+t��ծ��h�LBe�~�BӐ\٢t����YI�e��5��tŝ^q)�ŏe�a �({5w#�ەD=V'� �@�H()Rw�c���o���-�G���`#8��d�usbn�ko$�������`�U9. Bn骑W���P�J�耮ߗ����2u�Ze�M�61���ilt�V
�a
�*[��3@��!
S0��A�Yty�QvX�8݋�+ՑJrߵ�N�.�W$'�'7GN���$݊&F�N{ޑ��uz�i��]��A�θI�h<�)�<ǘ,Sa�F�Cb��c!��fY"(I���V"dB�� ��R�֣X�e�5N��JҨe�*28Ա�]N����}�p��4��#����;��)n��Æ��p�"�çD�b�'�I d���&*U�ή�uX��U1��ur[�;����}(p^��C��B_i��36��gd8�	s���#9U��"Ňw*��'L��+��IY��)BN�1��I���b.2u�LТ�0�b�Zu���V7�
�YJgtkm���x;u�����F��RڕB�uVQ�����!7E`�C2���T�t(Dd���]�y��I���x�j��0���/	aXh^�d�6_��S`�M:D�&	�|���Ee�(̥:����iuR�p��.k!����cR�-#1�s���k�o<�Փ8�	Hi��X����z�湕d�j4�ѹX���&�Z���+u� Ƙ�gIRER�}� 4`�[��4�2��3\͋�U	+ԅ���0 �G*^�GZ�N��j���#�� ��B�Gql���C:����-�+BMu���)We�R����]�6��*���yN�e�����Ϸ�4n���̻6}��Vz6kkD#%�c���9$��syߧjڹ5��I'r�rF�e�-21�'$�8,<�x�H�w�%<�\E�*����	1����	Sw�Kl�)ws�iP=�h	�2P�%L��b����Ǩ�(����w-��70�6&��w�nq���;�%�Y�!�3��}�2e� p�É��*G�̩u~���H.����,_;K�w�7T��]u+�t�����v�A������8bSR��WO/��nQ��{+M�s%}x�I\��O�3�xoB�{�����Y�)rͤ�	q����Ӭ��ֶ溋c��ƓҍX��B�*z`���r*�ې��<u��y��笵�;1��L�1��:wK�j	˶Y��ׂ7�
�!'ar��wh��բ���S�� :
����/c9gFp��j�4�(],�s, c��k}�h�x��m�d����$�n�����
��	@J햸k�@�	���	w1��a�z�^���h�[S-j�pT.�ü�U�-*W��ȅÓ��˨��iL����]˻Ueú즳3���L�3��Y�;	@���_ZC��f�WG@^v�K���.��'6�!7:�O.ÖB��	AU�T%�x����.���w��s:.��Ӛ!up񨖝�+����9�ۯ2�v�v-ӯf�}6��Ee�X��u��/i�+t/�7�W�z�G���Z�_%�f1�#��1��N�[��� �R�j5s%>a0���N�l�³�ͳ��7�����ڏ�|�[������'��M{�Dz�5HPs�M��a�IL��[�P��,�CL�Z�� K��{w'��C�1\�9d�>aM��0�W�Ϛ�il_0�ja�%3��.��_L^y޾.�� ,�j�Jm������հ�m1x�ӦC���Pӄ6�a�P[�JM�|�����H�Z���̤/�a�g�RJ���������}��fL���i-z���Kp�Hw�L��M6��@UTL�}���Θa�Z[�R�-3tIL�N�� �!�%,
d�$Y��5(��s��g�[�O�@���}�(�B"�`�Eb�,�
�0Ea����Wu�{��1�@PX)�4�0�i�Nv���yYBu�(u�'�D���Kg�V�]B��RgT["��B�)}��V�<�)-����2߷�=1�o��{L�KCL�{�
mz�4�L UT�ʖ�2�,W�9a�[3�:� m��:�������I���a=�����O}�%��8��ק|�|�x�iԔ�I�b�H�>�HV2RWyt�<��m���V����<��P-�h������X>h�Or�!�h[&ӹ�q2�:B��}��ֻ罾��i��u�����i��*��v�[}T|&�����l�ai���<�n\2O��:�X�)�~x��7u���ڢy�|k4ᅸ�}���}�oϡ�,���;��� ,ㄶ�x��R��/�2�X)�! e""�52̽d����Y)�hq�Ha�$�&�a4�%��U�JC��7�oU����1\���Kb������L��������a�œ��ݲ�RO9z�Ltb��Z4�کi���֐\|4���|��4�v�9�����CL�!}�ޭ0�����O%!�)��b�YP�e�d�<�b� u����z�Ц�]��a�qy�8�H ��Iƙ���Q-��P'�x χ��[�)e��B#^H�S�f��LɁ����
�jc^�O�铦�N�^�wp<�����Z��W}��I�:�����\0�@-��W��^��^�[�y��L7�@�=�i	�T0��Y<���i红a�����'̇Y��-�m:��wB��q�ͥ�	nZ|�e�+������c����r��C,ha�d8��T��+��i��d��S��qg Ì�6�Ad��"1X�	# �H*�g�oy���k���q��Ci� ��,EQdbŀA����e!�BF�u>{���%�I����L)��ahRM��<�ş0�(�|�>�Hi4���TX
u�Ms�t�^s�;�sת��q�4����y�b�'1ۓX�0�)ۻ5�����j���a��@��P�WuU"éH��<�&0���2̳,9u�/��Vy�����m����ԇ}S��4��l����O>a� 7G���~z��M!����Kr����wP<�O��7�RaUP�w�﫻�o���ZgX[�d�Sl�L�08�u%'�Ih>�S�s�a
B�i:�h��At�tr�CϙL�-�ɦ�i3u>e��<߽�ǻ�8�����Q�eM$�[o�$�f���8C�-��2{�l=�fRRN�Hq�'�q"�gVh�	��@,>� ��p� qd(p'.����8a��uI�m'en�o�--V�ɔ
@wV�Դ�WN�a��B�m��S,2�`a��p�)��{D��a�~�/���s�V����S&a��Q�M2,:����iL+)-C���Z[��A���@��^I�
r��ٖ�<��
kՖ�i�)��w�{��_��r��x�ӆ�}$��a�gqF-6Ì���L0�SHR.��C�U!l�C�7B�aI<�ou<�ҒS9tu'Y-��Cΐ��Xmi�B�@��/ν�]Qy�8U=�J�����=$8nc�&Ğ��윅o)b7÷ޞ�D������$�g!�a�M��r�HP�����m^��w/ Y��>���VX
q�M��*S]�~�6�>p���-���&sA�ӏ�h,�JJz� �KHy��P��ب����
�H�",X� 0
H) ��
@TPcDU�9��y�t�k4aI�(;�l�k�H�<�l�Q=T�Ӹ��m��Xd������(���B�1T�bJeX�,F*+�
iH�d�Q���N�I��S.�ؠ-�2��K��&� SI=��g���V��z�%�k����o��}2����!}��H�{����e�=�m0���=W	I�:�"Ȱ�j�P�8�e��]e$�:��{4L&�S
s�X.�(�6��wrw���LUn{?�U`���l��2း�C�F,P3��Ԝt�ڠ�Rz�	6�����@Ry�y^I�7�c�@
��M0�r�|�0�|�u7W��Տ�{��Bi�Sޮ�)��-�4��Jm�!׬�q��-C�R�I�No��a��S���CS)7���� y����,2:�Zϵ��{Ǥˤ��AI����1�2��y�a�u�3�S)�(
i�7u0�m�� �[n��[��X�l�0Ͱ�k�uxq�(�DA�=;S��U��@�Z�2�KI�$���a �E
Ō�����On��W�m/IPPX�_ڨi2�H�b��S2�*�d��e
�X����Lטa�T���7�{9�1��0�CM�j�I�S<��\�����-��-��
i
b����ʶCoXZkF���u�h6��L���agޣ�t�Qdz�#�����d}2���!�5tO&޺Ha3��*�ax�)���ҽR[)!���'�)0�&��^�R�Hm�'�i�g�S)NRiÄ{�׽���s�ϗ�0�L2�@�RL₳J�ƙ�;�i�Z\�l�-�3tZ
���M�a�L$�rȽp�XS�	-#ʔͣx$2�,d���.�����7����9���5��p���H�Ò՘�l�v���.�R�/�ew��u3mJ
��|e�He�g��7�bS/��BgU7��)7���P�Í��B���	8�e�|�c��az�`/3R[�a�L!�Pa��m�(���Q�B���@�U���KI�S:t"��*�����UbĂ��*����@H��:�7�}�ku�/�M0�<����r����M�����a��wUV�6�c����R��/���(�a�!�T-:�3آy2�O8CY��]����������nX
����ӧ٢�iZ��(a�6��O3)�-�!I),�4�a�)�'ot��)
O&�L� :���sj������Ā$A�Q+���F[�&���vE&Ғu����9aY��b�-�I���ۖi!�-��2w-Z4�x����1d�)۾�������s^��a%2�W(�aB�����y�=�S��`�JC��[�
a��On��݆R�l�f��5%��&P�a�цdz���+��Lz�Uhȉ�Np&}������:�J��`/]����`)+�[�e��*�`q�jI�$9��� Z=V�]�l��K`�آ�����R(u�m0�al�0C 2}�#6u����M� Qޢa�Ji�%���-��\0w�)��*���N戱f;D�Q6��[h-�^��0:��P��i&���{�ֽ��9�M2����;u=�Ȁ��%�v��{�G���J���~韽�W�������G��#D�gN��fY��U:���b�{F���u�u&��<Q��4���&#[���B�ojP�=�u����Q��s�x �cPUF1#U*+���U�� �QX�-�h�}�[ý��&t�->��N�
G-��ƚ�	����Yn��כ0=�y��N�b��7��b,�r4^�U%���׽�;�k����o�! $�s�n�u^��8��/"�*��`����w�Tw��1]�v7�T3�+(z�F0�	��2��@��Y�99�����ZԂ0�WQS�������Vr���+�w�2��_co2o;�9\���b[�J"�_܍�t(C�6Y}���I�̑3Ѥ��3�'b�
��b���u\�C�AGH�n#R*����]�A�Q"� ���"őES{��<��ꔳ�/$HT���U]���zj�ָ�ڠ<D��tܳ���}�#�y�#(l�=�L��aJ���nј�T�5^�/�J`�?}U��,j;b:��h�3�1i�I!��tE�b����bj>���]��C)-������g(�-�p̈ ,X�H��2��4���1!�m�JX�x"X�Y�?I$1E�֫�c��;�޵G(��H��T�2�"�V,b0TV")T�@PX��A`�$PH�\.3�v�Y�pƕ�Y��;�]�3's'Qh�E`�29P��2�^��{�4h��o'�HBD�S���6���Uv͜��$��!X�&#�����Ν	F�
P�
��簗�J�}�J��e��j�%��2{!�$�sf^B8�.�������j}˗���qf}q=�vjAK$�}�h��jC[�q溛;��b�x�x��7UAQ�;?0��w��#
yáSQ5[ٶ	E�׭��'�ި{ޯS��9�o��:�ؾ{�`AN����糠n7��Hc���6fi�8J�U"�۱DE�뉓yˉ�j��{:N�+&l��b��`6Y6�_~���o#�S<�",�i�v/nB�͋A��@V�j�a�p>��͠�(T��'`nGǦ�� {�%�"��HWd��b�k?������#���PF*�QX""2+RAE� ���������&�+�u\���S��PT�	��0V٩�G{��`�z�¦�f�>\'(����p`FGb��߷7n��&�g1�Z�p��u��nՃ��T�w��Gkv�=�E����R�/G�_rHC%�)��f+�����i��)�S��d��3T�)�T�s�W��Hz��eO$=P��ܩ(-J���#u�3���j�S:��3�c�N�ge��f̺��v���MQ�V�(+�1M�{ͯuG�!.� �[y^E�v_֑��`�@6���ޖ��fc��j�e�:.�AdYb���i��Ȑ¤�{��@v��.��:6d�;im��JKn�x{أ:"��h���o�q��ȩ%���X���Ί���B:v4��o�M�`�3S���"�tfg��:����qE�w"i�(TFEc �`"�Q*��@f����Q!���P�W�d#���e���ٺ��i�DBY�<B��SS$}�w3w�j�xxh�p{�ō�]��˅�*����N;Er�7_vHM! [
��Tt�ϯ��}�����G;hE�Y�S�l���-�'�����>��);��:
kZ!��9��ѡ��yJ�y�d
��;U�5��}����2�1�|�L&��5����oI��̀��P""C�<L T�y��f�\�Cۧ��iS}��6�0�i\���m��޳�D������)Qc�E��Ŋ��QR��"U�I���$
�a��)b�IDX�ټ�K�9���{ڮ��v+��l]H�jF- �Ї�p�X�Һe"�[��wq����˯Cq@���u�)"e�o �;�5���ĕ�5Nخ�7J��{����P���2GO7��\�hi:��6��A;5�&u7r����~h�;�0�C��^�f��.��+���.]7Nw�0%�|��ɪ�5.k�s�W��.���b +(Fd�E�,�\����.��n�j�-D��b �dE����Ľ�zM\��Ơ31@�u��j�l8r`eݴbԸ��j�su�M�`f�,����Ƅ��5�@	�<}/���e��&��o��X��`�w��1e��_�"�O;R�%�s��ɶ����**v��Lw���%⸰e��o��F�t����90�ڄ�{p2w�ٽ��ot����&G�^�(��6XYu �E`��]e��a�o9����n�[�)J^�f�T��Ϊ�PJv�/�Fk����)\��FۘeakY�=��_{ު�I�y>�{|���0[0L;�욍v�(���t}M�Fa�9f�Ė�'jQ/C��x�x��Q�u�e�C�T<�Y�-�k�fHq��}� 꿪�(��O���Ĝ?�#\�"黹HT*�K8][�	�.u����Oy{�o2�VRS� �/�t�
68�����بjճͼn�Z�4���BN�ٴQDb�DQB

Idz���O�_oݨ�j��F���m֩	�������5���gi���:���)��<���������̶(�P���i
8���;'\C �"����������x��r�-���YƱY��Wzp)N���H[w��}wZD�V1�kk��z�k�MՋ�Q8;c����� p�α��e�H`(B�A�PV���q�n#ֻvT@�ns5�׹rsܕ�`��V5��,AS�'>�>��G�D!7v[��g�a�[��XM�;O­<E��s����~D(��, cMU}��
g�������p���a�\�lZI|��\٘!��~�WZ��b�4�Gy�g�:؆�c����Ƅ�Eua!��`�2�/�g
���^�\
+y��w�qB�'N���B��x|�,k�Z<��Am����;Ы3V�!�c�bd������Hg���KY�o��ʰQFEET"�EA`� ��Ǯ�s��
:4e���z���) 0,�!��'����+���e��K��k�.��)��:��:��dۗLk�|+�BjK��|�����G��u�LxV"(s�0�xV�o�z�b� y�������������qG>j���c��ܢp��6��>(�u��D��@�T%(k�fJ?�EW���c�ǣ]u#��2�E��U !WB�,[�ͥq'7���`,��֬�L��NH�F:֍�*gO��<l�"xW+�u���h1�Y�I5���hnJY]H���L���Ԙn�yBJ�*�&�H�a��B@}V�t�����f]�=�)ݷ{�`�.Pk�h�;���4qz��c�\�u�r�ؼ��v�2U�
��L��]�:��gX�,:�^F�S{M�g�lSQ��
fB�Ėd�h:�Ai�u����;r��r��b��k.��z��&����h��n�amiԶ�=�qd+6�i̤r�΁s9}w=;i���׫�L�f�б�FL�]�a��:.ƍɜ���z�J��%!vJp�i*�q�d��泼��U�wx�6.�3a��K���e���i���l����(/n7yִH Q�ʖ��1�(h
%T�����h ��P>t�� xUA�22���E�O��MB �����b�3Q�,�U�5�d�+���"Ƞ��˗�E�3�]��
iP�0�"��U� ã]9�Q���n�ofm�Nb�RJ9��V���B�iQ�>$�PF�e���ul@�HՄ7���Qr7�0�ZUxW��|;]��J
L�bkE�y��$8_�SҲ��Xλ`���A�{I�Yh"���+U�����t�o�-Sd�Q�)�j���T�c�ǭoM���2�L�ܻs���]u�Bfژ�`�Ut�Z�znf9rhx�Z����oLW�j�i����PU�u�Y�a�p ��f�>�3(K�@�z���X�#�S�6�˾m��w]�jw4�}�o�F�Y������U<Y�k�̶��<`=�Q��7��B]r���`=�m�vޕ����������c~�f��d���d:��&��if�T�n��Y��Xг�H�Bv���+f�b=��F{�m�Xٱ�7�ܽ�*��,$���'ke��iq%�]�OU�9�(�����o�JX84I'yqɮ��,��,��J�*2U�Y0|�k+�*�����ēb�h��=&�f�Z��;�پʬ]w�u�#�D�:3c�oN�u3*M�b�y:�f
`�%X�e!ݕ�-њ�w!�ځ�g�/�Ŵ��]+i
Jޥ9�;�����wM0�N\�������J=}���nq�ٍ���C;mP76����)�}дe9�i,��Jv�˞���7��S��8�G��v��;����ǺIE��i.�8���!�vG�U�n%�#��4녋��*��1�LҾ�#��샢е]t�}f����Ӓ�7mnB�'������f����?l>'��Ѷ]��\-�]�"]?1�4��[鹲�ul'4�o4OA>���E���e��	�Bj�
/�k�']褍�J���Q�^�%G�/�ȫo����[��f멒-�u��s�r13��̷v��<ˍ@�u�\���X�Y��l_>v�j�۝5��h�S��dAI���W���U$7}1R�o6X�F��&�L��i�a��s�TFV�'t��qM���6�ƒ�j :j �hW���sj�{֛{r���]lP�&* q�{�ꖼx�jB5��B�܀�m�SgZz,he���eL�I�|��1	����MSm�U|��f��zA�iT�Ad(�|��UI+w��k�_b���5�^�UAdc$��)7[��[潜b뫌p E1��
�X�SI�9+��x��S��4fڹv��ʊ����q��C-	:E��ւ	�������F�1}'��N�j�h�n�:c�	Җ8���ąY8=,��aɆ�v��	;��u���ض%��;� ��c��ڧ�"�"�
(,�E`ꂑR���5Tb"�T`�(�DPUU������)UB��@U#1PDX�
���$TH�,U"�����������#QR!��#Ǳ�Y��w�=��7�lb�Y˻4�۲w��3���l���Wh)Fl�+��tx�:��]��'��Z�	3ս@١S<܎(�K��0{w�~�{����(ȯ��(��W���³Mr#8n٘�Κ�͚A��Ei#l�?�����i-����5״v\��].N���s(�,l���ˡ�*��^�x@�|��!!���}�6L�}lqҴh��0{�Յ���u �Df�i�5�V�u��'8���E�vۮ&�6",��Ehŗ�N��9�\� �R���(��TF*�0QA"��+X�"$Q���������ϢE����
0����ǘ�Z�APT�o�v�6&f��nce�%֢Ѿr5m����o��M�<-7do���^^_1��m����Ɔ�T*xx ��j��1���hrCNj8���I�ΑNځ�w��#Qe!Yo)K����}�26�M[K��Y�N��X�<�wb@ !�^�)(�Cc
�*g��z��z�o���Q���T�H�Ă�HS ��U��(fg���;��%8�
�h����V��I���m���z�X6��P�Mf7;�[s���뉬�[ksw���u�O�!F|X�w	#t�ۛ��� G���S�b��%��7�G��.�uq)9yC,�$�z��G��cz���y׮���S�=�u�1���Ш*л��v����ۘ�e�٩i�I���
&vb1�@�s���5p�a��>��`�
��@b�T(xU���]��ޝ�+��I���*��V"���h�EQ*]֚^W=Y�wn��r�0����m��%��X�&�T�6q�'���y������T��4bػ�e����\g>�gz��CT�����y��>Mv#�8mV��vHw2n��bj���#0嚜�u5%ƺ�&ȿ}�C�{	���Qo*��q! �ֽ!�`d��^�(ͷ�|N�@�5~ǽ��3�k��j���*���F�&7Ymd�೪U����I �IAI3�w���Uw�[��B���2{ ��g7�����m��wG�:ivu���ST�ԕ���]�R�M�h�<fW�2/���x��{S[���&,����Y�+"8�<�?��@VSo�e�����]��c'SsRF(@2��v�]��^�����W��?Y�j���l1�6�{S>����k��Ȁ�f�A4��B�a�9�,$}�v&!*Rdir� 7�c�*BCe,�< k�9�}-T�B�M����X�P�V,H�#|"�g|���#�h�|��J"œ������
�
���^�[�n%��t1ZM!+* �L�C�ˎ�Li�A�7��k���W����,��*�:Ver�s=g��\�� Y���	�z�f���
�b������`��F,H(����Ј��[�Ø���mK1���o���U@H0@FH�dF�I%W+��0q�8��t�,蕶W��&���9.c��]E/��O���h�����[v ��Uz��W�����_�^�>�y�v�wK�:ȋ�pX��T~��<㙶��݇`wz�H�zW0���8TڒR=Y���LNWksqI���ûj�8��1���w�����G�+�k�l|~�I..����d*U(�6��|QO|�=��t�� }_u��
�������v�d4Gl�t��H������o���fS��FDH�A��2 0PF1H���E$DQ�"���z�t���qx��N�G�#"-8T��ږ(��c=q���9zfsK����g�Yٷ@PGT'B'��hR�ʜ����w�,ye��ɵ=>���(?l$1- ��G㝅l������vǢ�޻<����[ ~c�9��B��J�73-#��x�]e5˨�=�˳+��wK�r����� *����U��c�ѻ>���p�r�����xvu����pI��x����J�Q����ё��v��2�Y�N�DA	rgD3V��#���B�AADF�JX*(���"
�L-	lH,�TUX�U
E���W�W5�U��7� ��Nu�/����m@(&򷨵ڕ�\�Y
ыFظJ�q�i�9��Kݷ�B�i����	�{K��)�F	�ą!
���k�$ٕ��0�g/���SV��V^�ke���;��v$m�ܵ@L5���:R�%���*���"��1H �U^*���'I��v�S��P֮U{��UUxh���϶� ,����$��LF�Y�E�f�
Q�;(Х���x>4�V�2H��'2�;�NY���g��X�\���qp��W��6|YCf��Vo#�nA�S����D����b�'��5���=���8���w�����~�ߛ�����>&KE���� ��z��"�M�(�+N��o�wX�B);����<���!農3�=���fHuf�f��'MO{�@�{�+��w]֣P�* 8v���&��1��m�r��J΃$��6�H��?�7�� �&�zx�C�9���^�Z���� �@����u�ԷB�\�\�.�A�b]
���N��R�^)VrJ�6b|�tb��z.̋�,�Ħ��Oo��듮���BG�;�ʆ��UwB���b_���|�T��=���Y����a�i)��H���/FT=j���:��}	'�Z���D@QwX�Y����eQb
�	2*őH�TVE�k:�z�b�3�ug$�`�P�P��m6���bujD��b����mv�[�yR��;�.rц-�@Xve�K
�$DuC���d�r�D�ޯW�`����HQ�5�t�7|�vO�n���T��`[�Poc���S  ��>�i��݊�b2���gr�7jd�9�;<�9�^9�WD˗�ok~��I+d��"�ȫU�����4m��뇅�F�N��c�$ε��=K�4x�Ҹ�9s��ϳ�Y�[4����}�ζ���w��~?G�)��Ҿf��� ������u��"U�}��zR�J΃���s5�u��5�c��o[�u���N�R@PP=U�b��v׳O���ю�������[��J,�y��y���l�:�j��[�Dk�IK�1�����1�
쏶jl�\aqS�N�Zi�w�Q 6m�����n�{e�^> R�E�����*��(��U��A��X�"�E�(�(�ֻ�V�w��w��_����tUfEs��_];�;[�Ph��hR{w��CݻI]$�1qN��u�<>��o�4�}�Fa�8��dڴ�e���O�.�6t�����:xdK�*��UV<0��%͞��g,{\�� e+�۾o��Y�u�_5d����C��zu�B�Y(�=�g2;��p�s M�X
0_JYv�\�\#�C� �Y"*��"�DDDD��H7�p`C�~l�Ga�f�sc>�֬��u�
]F3�w�л��%�!��%�Pl�"u≩��.:��i�*�Wp3�$+`4D�':$���N�ڼ�kM�Z�Λ����\K�8~7 �&f"D�f� ��b;�_w0��{4T �q��6 4�VCҹ���q���뛣/$:�DP����)*0`��DQ��H�F*u��HD@D��(AET�Jj�4i;��euZ�r�
���.w��m�-Ώ���� -��֙t����o�O��/�vfi�SP���'�f*�\��^�L�{��4�n�֛������r {q[����� ����>*U^�K�iV,VF��'�i1C91�I���1.�K"���,����}qk5K6;�|���Q�B��(W�W��щ���'�&�}M�ɑcӂ����ʵ����wGU2�x�_Q�ꊘ�&�c+BQp�l�|zM�}��x�Lfm�D
��FH,�dR3|޳ݽ�� �9hF#��kMv:*�#�dXC4�;���m�z�'����iW`9���/�ǜ#M�3�X���G�5�/�h�È�Z�� ���{��K�9-B�&X�����A�&g]�mm���N��#8iLK,�� ͻйg�\k��'tr�(�_v�EK5�s�\w��f��n���BL0U��dn����z�w���g!���b����(�UF���X
�����=^�*���p�o>�:���Ɉ�a���f�ܯ�	��ֱV-ʓo�f�L�2��I��V@�y+�r�����Y̗Ur��zh(M'e���H�r�6cl�Q/���i��t��3 b�f�67m�L�"�'��m�N�X��܍�<�Z5�O;	���ٳ� g/���3���	��7nK ��xP/��]Cu�B%��z3IrHJ�ithwK��	:Swgq�O=л� A�X_Uz�%�&�&t�����ux|�U���2�^p�y�9&v9������2��{�}e�m4֎��0l����N��K�H�{�(-
���t�+*%��^��Ϯ��OE����N>?�c]�~�H��	����.��-��k'IЪGi�I��K�/�3���7�b��.e�$77����֘<=@P�# �"1��"��`��C�f6��#܏�~�Ux�{���2n���|_%Lw�kd���9ǂ	�YKޗ����GBu��K��
V�fmG��N�|�>�P.�u�j�Y�|E��{@1ٖjc��3�N['�h]93_U]F�[���;�Sy�Z=A^s��c�
��Gƭ���Z��{�%�,��k)r�lP^���TԷܫn���:���Ω�7�0;�˾��#a��K��Gv�#)(/:s<C����@.�7G����n���v��(��mJu{�($_ΊqOn,*��0_p�4@���Ht5�2��*���2�GS�MQ���¡����y��u��E�t�nIq�Bʮ����XV��)r�L�ZQ>=�[�YO��/���qm;��Fu��*�E��	���H^�n�ե�;jK�A`�BW�'.ۊH*⩬��aH2�rL$�P"^�ҭ"�e8`h()2���z\��u}�#������
)B	"�(+]�D�x��(m
U8�b��s��^�U5����0QwwuwJU�Z�Y�*B�����QK����\F�FEX�e��}���r��7%�6.J���c�V��GR�]F ��0��c]&h��K@�cK+5wUL`T���L��XpY{6��\�Z4^0��Q��&�6��WX���Z�\��ͪ]�F���f��隠)�1���ʹ�e�*��!M��,�G�RL�L��.�P���m%�F��H���Bx�u�tWP�����e�G�*ʘv�6��吣��Fmv�]��fa[�W��fAi2��p���].��JɺF�b�q#S1Y�i5�л�yF=�
wR��Fop��-�p�jV閁��/��mE�V��x��]�"���+� u`�U����f�A���'t뫒r�z�y�(��4
���ݑ��q}G�^?��3�&SqR������M%�u��#xS��%��7�y��J�^��}���»4s.��� ���MlnL�1�]p���&���&����\�t,)��CO��kwJ�n��@��/o�wȌ��x3��7b�w���v�Ԛ�f���6��+���=��#���rI5�e�Jܛ}�^n�ܡE�5I��lx����`p��j��`��J�Y�o1�!A,�8esu���cr�-��0���.Z�F���t��xX���]N��P�m�Y����Ƨ`�[۷Ju �����o��C��"g�G��8(�-ٵ�i�-M������i���aW9�;�S�и�1΋��[Qb&����u�g;ޏ��9etX�}�@�q���9��;���~Ꝋ�P�xg8+\\ygZ�J�U��� �]8�kMI�\]\��mk�&�#��"܃i"�<bv��6��fD�y�,d�N#�Nאڈ�6MY�q�W�nP�6�	},�*P�H	��̸  e�x�	�`�w[�Y N�-F���}���ƫ)WXzg\Ə�?�bJ��o7[$u�ܓ�g�����H�N�t�F�9)	e�.L&�(�;0�v���⠢�t��A�zu����;�5��w� s��*���_<�:�!�KxI{d��/U�Ev���[�'I}Y˻x`Zf<l@bNW��^��U���G�B���z- ��(3��8\�q�Ϛ�D����-!�^k�7�xI�ǸL���T��:A���
#�(��	5��$�8�7�e��W�*D�j��ϻ�Kw7d�r��25�C)��"(��R�q�:�^���JwBց\ #QՋ=���T�l00ňe4+��$&�{܁w;�$��{ޫ�;��n�`!���Z/��f��$1�0(\��{����N���u�� ����~�c'�0h�w���\��T�� 1�0c%($AUu�7��]5���j��&n�}��6u6(,FEX�F2,$DX��X�0X�H�Xŀ�P�HK��ϱ:��c���>�:��i�'5�/��2�U>��wP Dt�s`E�w��0��薨�l3�=� B,���������n��w�޲����%��%�wvi��b�K�8�5"y�4f����e�2����2������:��3͸��Juts�)�z'�����*a�-�U^�����aۛ�J|��t��.Ɓn�Q3sU�r�>��C���3t��{'s�0�-TG�b��/����Uof���Rt�"v1��(�P����5�!47PE#��p���|~�P��ت��`��N��
�_-��d��Hh�Z�\�Sѿb�g�Y�Q1HxHT>�['�o��j�s6�0���?�A�3�D���������Â�&3B�r��u�S�M�T�Op����;[���X<*a�1�`�H��y�wt��^- U�ۦ0�mޭ֯����5w~�>M��I%EI5v�޽�:DR�D��`,�PE}�Y�3����X�(l<8��Vb��lX�`��#�LT5�Ye���}\޺�M`�W��|OvSW�HLVǲ�RtР�'� *��3"��ә�u���P��У�{)l�Y�Ĩ�l��.�j�L�3��]B�t��7]��u����K��9KU��t��c��Wޯz��oɤ�+�!�q�IAgU�3���5����~��@m��0�#ҹ �|����L�D����p=�{%^oLr�+fdMm�nQ#!��{���꯺��}�-|Gܴk$LIO啷Y7![@�R:s4k:J�>�%]R��;g�h���r=[��^C�mEm�*h�:`�JV~���:�����d8�}��e�C`ɪ"4�>�!am�B`^��]c#A��y%	3h��&�PR�LvK�hi#o�,P� 0����PUTDPb(,�Č�Y�DQc=�޹�W9���Ϣ�RD@FE`���W�&�����,����AS%�i6����| #�uV'�G�>��SdB�.�w���꫼��8�m�M�tۥ�g5)J�Σt�� s8��z��b�����t�<�\;�LL��{�W�����Q��.���
"����+6Ùb�d����Wr�\�d��o��;dJ��t:�=d��w>��[���s1)X^���A�n6�L�C�Q�L˱g:�x._���PؿFxn��`�mT;�m�8�-�f��ƈcMјl���Vy��А�V*��� 
� v*���9��
��a���Ɋ\K�PA��aŚ0ƾ��=�n|6v5>x��%E�Wwt��\q�]�
�̡��\��3���ް����͋D��rg��Y�����{y�"�--Μ77ro?[ٖ�޴۫\,�*�4�8�&>HhF�h<�X�� ��*���*)F ���k9������浺�ݚ���syML"*�<��<LI���0o�5���jZ��T+�:ս�؛:(q�6jT���Y��I��$����Leo��C����Q�A}�-���K^��D~���>�M�Ĳ.㹮���z7@�����Ԣ�����6B�j3�f�e{��=�y���ڛ7��3r��	BA��H�t�����iU���u�q탈ڋ�J�[2�lў��{ݔc����q�Dvr�9m� g��2�S<0�d�X%�r,hj�5m�����æ5�ֱ�۸B�(�+Ē]_(�����x�^�Ω�h�P�d�om�x��El��sI'��	�4��G�b�w�t05�y��ry
��8��~Nj���?ު����u������7���m`ٚ5�Vh3j]���\��>�#����D��'��5�s�Ί5I�=;�a��m��ʽ=W�lη�S��hcV�� ȰU"�6��a��E�H�`�Ab==��z����� ~f����s�R��M��c��i�R��]="��{/wT�r闌q۱�fR�yDtR2�@���6O��&eelֺ-{M@�C_xx�;�d���+K�P�j�w&��|O��I�O7gpA.���f�V��ف��HX�кk��֓{�D�q	�����9�c=z�W;-=]ҧb�}��̓��qҡ��wky4;�'R�=!�Q�Y�5
	��3I]��V*���V�[�\�$�R�zI�Zfe?��z{��
���Gs����i�Osl��1ۜ��r;R\٤ZX��z��NDv���S�h̲8X��qya٫c���[:�DU��Ԫ�r�u^#��N,���� &tᾇhg\���b���p�j�}Z-��#�v.-zGJx�)��d�-f6s~�B���[�R� b�ōtצD+:>
�u�.Z:jB��( (�(�,H�X�1��
1 �EAQ�oz��w>��w��L�Y1�I$DwZ?ʪ�)ֵ�l~(Q.7����!����|O�G3����nEӎ�Dt)K�< ba��`S찭�Z;�]ܼ��E۳���I��mg3,:
Y��^���@yq`.L��a�ߎl��n-ݲ�YݹD3���{B�	�sS�?�{ ʼ���ӆjXs�@�5�Vo]_�59Dخ�UUJ#	��Hֵb��+}�
ŋ*��� ����#A#���F"*"�X��Ɩ'*�"�����
"�� < =B�7A]��$��
��H!��yڮ�Ôӷ;k�rX�u	��r�����B��|���xgN�.Iv����n.�ܟ,ފ�g��w�Dv�U�����g&��V8M7-q;{}R��!r�}�&�d���+��t���a��*�H{�y����=��ޢV���@Hj�k���Ԡ�;�,�NO�ɠ͗&�NҪ�����ǉ�����	�%����ֻ]V(,"�F"�"�c
�
Vn�4ʹSmwD���H�Ih�%t�r����U^^3�v��=�9y���<+EK
�BX�q�|�}�9� f:�'�qS�w��0��p����j��Ƞ<��#�X���<��ԯoWe����#cX7n�LPz��`(d#y�c�¡��u��o[F��x^r&��@�1�%�`"h����}� eo��Y�qD��d�u���, 
 xot�\o��B͟�>�D3����@�$r��z��z��Yi�]Z�v��SWu�y!t�s��{{0㙽P3�+�����iҝʡ>�k �+p��7s��.A��1WE��N��أ6袜���fx�i��m���Ā���9�ɳ*��wX�k���4�A`���wV��u�|8�VGV�D�[ݫ|�;c76�-mޛz��ڝn^V�ͼo3@�Moe7��`��k��=UUU��D��,@�c�y��aX�X�DQF"-�\�7��Y�*��Q1L��{x����i]��F�qɓ�,�b�s��7�e,q]h��ٞ�o��;�y�:>'�����A߶!�Q�c_u_]�ġ�:J���L�[�3=8ً:Q�+�m�"���'l�dEq�Uk/���[ׅ��h�J�*�(���J
� )EQH}�5��|�����RN�A��s�&`�˽$�����e.�MP��u	�{��T������;��W�r$�v��]^�[�ó�&��~5��4ll���NL��^�.Uۙ�x�#��&�v2��,��q�]�j�O	�4�v�z�vp�gp�  �˪09�ǲ�p�-��n���N[���4qc ��}���J����M�=R���vo]ޯw���w���ra@EF*��E���dPX�AD$XTY����uu�=�ze߀&���P@`��{8��d,�BW,�a2-u �o��k���p�G�1��a9����	L{�I��·���/kݜ���;?~��D�u����D�Hb���-`Q������-�u���'49�G6�Uj��C��_"��r�t�
���e�v>�{��q��S���s����)j�:�gIۖ�g@�c�ȃ��:������ӻ��T{E͝;��j�H�$�:i�sR�{����s$�4Nd�*>�n���ԕ�����]�C���a
��&�oW^e2LȘ�w#f���۝�p�D��jTIf�ɼ�wJE�=�{�W���vs�e�`&�����y�O�>�ӝ��-��u2�D��r��˦)������{�]G�V���W�}��r�p��<�U���u�EdAX1DD,�������BF� EdD ��(cкq=wJs� �޽��-���p��G��TV^]�Σb%�1���=����טS3���%BBWS�gj�{��̍�l��t���Ed_%����Ed�yڱWo`�+O���I}�f_ �[�{ݲ�ò{]�ĵ����H���)!()����h�k��Nl��jї��c�ݚ��R%�4-nQ{�v?p����ƻ���㥩�s�#HA�}��v�p����yG��#�e�A~�zbN�*fZ��b��7�Sk	�ʱT(��@�3�" ޖ��E�r�-�S�Ax�hL�����St�I�y�dQ�}y��oo,�UȚ�F�[�خ��ݥsk��_=�c��v^Եt�ZT��U� t(4�� ��ow%#yk/q�P��1
a�Z�R(",��t�^:{@TR�\���ڭ���t��2�vՎ��m:f�f�]��M���Oq���|tN��*�]2[��ʏbg�j�<47TuX<������~t-oE�H�Km�n���]��r�D^JV�ڑ/Aza��2��z3v�7PaV���c=I�lY�n!�^�Gkk� �ݮ��Kr�Z�dH���I�D������C�UW%��x�q����1u��s���z������YR�����(�z�ӻ�q�*�.�B��V��*R;�lB������A*��U�A\�h������
��fڗ���w	l�9ާx`��LV7�6aĠ��]�J�t�j���`޺p��!�0���I�\��dz%-��Ҽ;��v��W@y]��ϲE��b@ya����	��n���ě	P�:��1��U]S��on��j��!w�Y�0���"S+�p�++[��,/_J�]O.�F�O���� ]��Uڡ�n�f����A���[�`�)P�>���?�����)�������tD���9�̛�E�����X]�[8⏴*��$�\1j�4�M
���Y;�Be����7qp8��ˎ]�eN&�������D'H�,x Wu՝�X7����j�lW�<�c�fl�r.{/���8L�'�HE�������AO�mC �b\kOky��Ήk�1��dvL�3ׅb&��K5��]k�U/xEd�[In�(Uݤ��ř���Q�J疣�8@�![��_Q��zf��F�����3:�-Bo4>%wY�s��"W.=�iS�mZ��`��w6:3Ю�j�O;�_QO�[�u��<BmL�/]�ݣ��&���w�k�S�>�1n�t]?�=d��km1r�<�ndٵ�s�����,�Y�q�z�Ź��^�ھE�z#U���eΉYz`ھ��%k
���#�Kg��{}�n��{&�.x�>	��Ps�Ү�u�#�0l�A[z��HXwmuF�:�;�"�#(.k�HQ��zF�o�m���-����ƙ�N@���;v

�G	�����yֈN�*�}���Z�c%S��P���.b�5�M�t�� A���.�]`64���P�{F2��+���z�������K�Ҧ��tkD�v�w
��'~}}�"��-�$c#!��*n���MBFR���eWo5gT�nڌ<�`�;]恄�ɥ�ϯ*&�k��{�>�|��L6u1l��w�{���R��]cU���q��]NՇ�0�)�nv�WŸ��8gvP��`�����y�5��E����:;(Tۗ����]M�s���{M󷥞̬���=zw�������X$F$$�����ȱ��	F"��(�$PF�Q@�A� �w /Gl��.�bLN��dGЙ�up�v+�:����#�V�r�:D��֗M��p�Ϻ��Ί>�;�3{� ��W&�e����ۨU3�r��a}�m!�C�tN�hv�5�RK������l�9ބ��}C���]t�*FHo�!��Zq�{Z�B��ur�u�杻����f��U�D����/���Ǿ���A�.g�:���uu(:�f����vc����[��9��v&ͳ1�Z:-���ϴr�;�O?�x{�(d�)hSD��Ó�_i�}���G�����)v7ye�Ģ�/+v��g+��Ӵ�WK�Qͧb,z���頂`s���7�绶xE����W�]����n���oP�+AH�b��)TD`(H���DFDX�^�Xλ���������A@A` �D#�{��F�):	oD�5��ۛ4/23��4p�ow���1M������w���5���}s��p}�{���
��卒*�p��[��K͵��P��x�s�}�Z&�Z�(aJ�5��˥�.���L�'��r�ogqK�{��z��L��~έ��+�U링�2�e�K�����S��1��9%�`4Ƅ��v^��Yщ�ɽ��l6uD%ε�=�k�����h�H|pl��dh���y!k�"'�qJ[ۂˎ��Jˁ���I!Ԁ�1�gw���󚬶^0uoK-����%���m��T�yB���M�/���p���钙��[�Jz̹f6.Gg+�r�:��S���&Mӭ��f�Z��޵��|H�� E��B��y+׽8� �H��DH�TF,$ T@`����y�p�y�c�\�sW[m�䣦OD2�)҄���]9�&�ٗ�&:*��r��2�����ԡ������~q��ړ;�Jm=�w���%�{�۲f��d`N���nY=����յ�:12�R|l�cFWSb�o$�d���7�����*�{�{� ��I����I�i�w��=^ޫW c������a��WIz�}��
2���hQ��&ӱXyxw���Ӷ��4�V/4��ɸ� �w��.K���gaΚd�a�Q�s�=��������y�j���흍��뷥��Wp4^Q�6�]\1w� ��A ���I��U �( ��P� �FH�UV@�"(�A"��(aI��վ��d2�f�.PQҵ�w�jM#C��+&f[�R���R�+��D�y��}lͤ�t��1����ӓ1r����W����3���뗴/��ۺz�y�13$Ĭ����ghԺf>����vA �^�ɽ�,��䗯\�[[�����s.���l��KQ|d_R���O6Lr�7Й+��4>䯟ZWã����,��Kɽ���s`����[Z��������w\n\�69�^�ٍ̝8��Z<6n�1�x���;�����%�s�c�_>7�L��;þ��گ����O�A���U/��\��=���*T�Du*�G˞�ɩJ�� ��t͝y3E�d��uJ�!��q�`\މ^�'�V�� W�=��
E�� �"�$V)B�xxUbm��Etӫ��1X�"}�W�ު��ߏˏ��/��@,�k+v�*��  A ��Һ˭xv��[V�>�WV-���T/�(ٗОw+ �ͽ��Oi���.+!;��A;72��y2�8�|��Q�b�|��s�4�|ƙꉹ{'<eu������?�N`�,��5��xy�s{f�jg3y���e�aǒ���+��Oe`y���yˇ}k5J�����o3����M�&T�k�9�{�Uo��z��P��D (2]�89��-������̃����hw`5)�5{�1�p.�=�m����5M��<�L�}����N|��IG��Us ����.�i7ǧ	]ь�&�7�{jL�������F7��Y�çǯ/r����K���}�Wн����hUI5)J�PDd�RHв���D�{��]��{��{���� ������#DTF*���,�1YQ����+1Pb�Q��k�֟p�J��
]��wgJ��K�y�Đ�XH�o-Ug{}���k�9���[]�tC�rܷ%�j�!����Z�����ێWk0�45��Ґ�zݚ��h�O�$�<s�x�k��fd�6	7�̵\�e۬?{�U��_t�����Y�ڽR�.V�X�78����(E����,:�]ƿ���iw�~�}����n������[Ĭ��kP��,��[�y{�;|��޼6����}��V�.��Eq�S��!�{�|zn]�F��Z��hr ��SuD��������[���w82�r&�������.��}ָi�*!o�&_M������\����x����zZ�c��uzY׀�H���cX�DAA�Q��
 �$�b(�,bA�{P��S�ϰV�����S`�s3�\��0�M;��ٸ�GʶÔ����n��p��1rW��S�P�P����,���Bᝐ;�+o9\Ćԥ-.r�9�7!��R�gd��z���"=��)E�8�eH���<r�Y����K:�ftj)�]��N��M��^���i�s}�b�'��nz��$۳�vM�`�Z��K�I�L��e��i�2�f�2��D��T+�U�߽�L������lI������OR�N�3M�}c�}bc�������Y�:�DI�RJ�����g^�w�zJ�sw�=�(���ĺoo'3feȸ��+��m���:�-r�Z�;S�}�3qV�Q��]Z�YG���	�%�"(��� �(�� ��P�Mc��{�y�t&N�`w|�3aT7�	��Mw�Y��6�G�0�T�V�I�#����|�Y.{��]�ۈX`��۽"؞�$�:����`�8)�W�e�u�fc���  =���*���<��Y�����K�U4YN��
m�Al77$z�kW����u#(f�n�O����ӹ5ڎ�S���ZK�!��m�j1Ӏ)����%�%���r�+��
ϧ�z_b���<@(���ء�����<����Z�0�������C��ś!i���ٌ-M�����MF�>٬k�l��X�>P��lo�y�`IK��|��W'v��k."��ѵtU\e��� �땍B�W�\��y8t�M�oT|t���-5��<]���@�a�i^���}���*w����g4Iv{�7&<��-K�X���c"(�D1$�
DA�����{�V]]�&`�Q@F��QUϜr����wg �Hv)"���9[�s���Tr�7}}��]��u(��ۼORGgY��!��z���V�)�v��<2�=����q�:���e����� ���sU�̼�+Z�7�����˭J
o/�l�K!�����u>�0���h�b�l�B.,�+^�]F�s�j��\�4�l$��r��ު���pn'y���Nv
�g0
�{����cg9�}�/��Vz���R�@����2�f�6�Ku�V��j;�]�Z}�ҙ
X\�M��cCge�$G��f��{�%oE��>0�wޯ{%w�&|~j��X[���x�ֱ``o�j~��֚}�K���jf�����bc�f�0C���g{b���<�k�sX�`����"*��@� ,"! �(��Q��J���ۡ,<��`�:�p�*R���S������3>���G����g{vܛ��}�f%�ڲ"�xx	ݫ��w�guk�N䬕�k��|�V1��;�\��;`e�e�^�|])���ޔ���Up�V&Q4�������ٙ�b����.��x!gKDPQ�[r_V-�LK�!%�.�ƍ�S�oV"�Mg�$�ۙ:�K�Gl�q�o�9�Ww�($H�(�DB,E���y���F^�����Η��Ky��T-��v�I[{� ⮌ߜ9x�OC����r��z�U�%��� �&nWs�]5�1�9*�I���C��;Qp�㫎wSԉ�Q�љޛ��&�]�c}����Z )"ő��,Q`�,Q�s¹�q�z`�9��E"0TH�2XLc�}�������ekpbp���]:i��O!YYӫ��}0ϴ��Pl��4�(��z�6�ĚJ�v�;[�R;���X�}UO�r���55�+���Y�L�	q�>3gP&�+WKu��o�����NT�8m�̙4����T�/a�.�2[�\�YN����]!�f盎��(^�޼��(�Yb�)vo�W�"r�N�J�^����K]^��_&/K��� �����C+٠vF�|%=5kUp �kጂ������y�|3Z���
����D<����Sr�L��(eJ�����op�� M�v��@M�5��R���=F�K�H���ݠ�詮�_VJ�H������nY��U��Ф�*D���[�t-� xe�f��3ޠ(��R����Ւ�9�y�-��t(�Tu$)
�������G���c,d��uGc��{�e	($��t T V;AN�х�r+�	j�<�fL�e0�-���	D�#Z����rS��w��l�t R�l���vk2�s����5>��p���7j�+��u0#�}7�9>ʫ���WY��w��{:����/9���g9�'|�ob;��)ɵ��цFf�R�Ce�4ЍD��� ��H����x�R�֎K	7�,T�S���ьP�iWV�e-�T��+ګ�}W��l�j�)���T[�����1I2�e�	;����x�V*���fC�4�D��&p��hZ�R
,�(��:uj�=�{���zV�̫���>ڟ#Ï@Q�g�c��Id���~7��bPB�D^�n�[��GQ�U2�� �;�ٹ��oq�-a���R��fq��[n��ސ���F��F����Ŏ뺛�� �Q��QRRR͇8x��Yٹ��;���2;�[5�v���g�ˬs���i����.�w�rY��}�:�JU��=�!����q�2�t����n�ܶ����*	���v�����0��t����$͜��
��_��/#�Sf����PNlܲU}d?n����Jb�2�<�xNIU��R�Q�on���(m�;��sh�j���ѝ�{��<��@�ՙ��$+�=������܈�9W&>�C�v/r��62�b��r�����o�;9�,-�����+�kԟK��:���L�b�w���$�ǉK�lMg�P�t���S�ދ�z��q ���sI:N�w|UZ�u�af�Y�r���n�b�>�5��H\뎯&j��墰U��L��9�mi�}���}�3[�}���e�8�����m��C`��h�|�,�8�NՄ�pr.�����3v��5�ʹm��:rgui8w�`{���wv���;�{of������:η�+�a7��u7gY����FU��e����"���Q_*��vһ�4�bo�.��FgK���w��:3��6/��4�.���s���N�皤Ur<Al[�d&�1�Ӄ0�+��T�)������X��N�$P�Khw��MMx���՘e̵�wU��9�-Սd=�M=��G�[�j��j�0��3���f�!�6��:&V���1]@������ke�c��|�m)�ģ�8�K}+�i�K�BJ��Q蝵��D�^Vn�gU�֚����ܙ����8�F�>ƜKp�+�b6"9]pƷ^��Ω��m7����nQu]uc��J�3.czHN��8m[l�r�ȩS�d���`oz���sea�3I�;Az��3G	�s��5�t���w}��6;���:L�vݜ�Mև�L}^�d��G�������-`ż�[(ΛJzz?��}���X��y�Sq�:5��b�0�m��j��.$ t�xx,�kw�]�b�DDb
�,Qb�PA"+dEbDT��k[���<ֵ���zp�9�B�˓/eN�F&�7~ߢ�sҶF�n>�K }�=4S�����־����Ŵ�s���������cʳ�<��/�,h�k�����I^ѾD��n������8�����m���NN�1���F�W��z�Op�غ�Q��F6���������dUz�z�*���K�֎*�n�Wo�쮛��v�V]���Vd��8N��{���$�,�h��㔍�m�8��C(��p<�x܃:N8鮢����ũ�|�[RË�}g�"�u�S�]l�멘�9��O�z�~����B>�ږ����_{$2w��f�	�M7�%{	[�A��cY۳�8#gi��pIn	��>4�sn�Tx1��FQ`�Ƞ�$��,�,#F("`��l{����zw;�~Ђ���Da�Aa՞�4�;~7|ϳ�<�k���Y��cnZ������s�3�Ash��~Μ��[�M̾�˙6\�rdb<iŖ!Gꪪ^ߧT��C�/�6�"�F�-�������ڶ���u�R#�ge��u�gN�3��H:q�j�{�����o,�220��P��z��T�M����Wt�qLܒ�3y��o�gs�%hgL���7«�^��������y�>��e꘦��&����r�ǃ"���^*�6�����[)-�غ��)�è������b��T��:Ҝ$Mёɢ-�׷�Xrg�:��������o������@�O>U`Of�����~r�>'�:7�y�<�w��K�Fuft8�j�}��;�W5��"�E�Őd � � F,��^@�*sd�d碧-��T����T+�B��[/㻽�����M�m�\�ZWw��߃����2f1r�ߙ���v�����U��+'TS���q�^#��|noہ����o�f�gM2�^�u�4��zWT�u��Iȥ���wvoLe�I- �:���@3H@�����{���3������}VjB F�`��ˤ��uR)��W�/*�Nrs�aE��<83�a^�
TY$��gz���d�jg;���髹/k����� ��λ����lsRV�cr����=��(ż:�Ԇ�uջ:i�a#s'f�s��H��s������T�p=�%�N��h���]���u됼��5�g�wR_Qaw��\��\��rN㓊�or\�U�!�@����c��T��h�d`,QX�T�2o��Ή᭤�/RdE.�}y����DtVkiM��O^�&��_@�d��={z��v[���it�����mB����f��7#��"�9(K|��J������=�B�VS&�o��}��v��s}s�Ucw��n�z�B"0F#�ΒG���k�V_>��7��^u��f�����r!��MpC�b�w`x%������9^�]Tkm޵��4=� {���U�� 0"� ���}��������nZ�n�lVN�kr��	��	�fO2��*D.�Ǯ���ﶬ,��qK}WY:����P����gQ�藼�vǳ��������y���.K�Ϝl�U.��� =�[}��4�p�2]i�,""���H(�
*"	wYۊ�q�n��C����H�TdI ,UQ@�X�"Ȉ�9֫�\����;�8���R����i\0�ܼsz��*c�'��G��l|��>��e�왮�f~�~�m�g����=���D�R8�5�uI��h�f{�ų���Rwo��o���f�
�M<N�x땺����$��$E$��Bo��9ϙ��'�G�u<�޷�;Oi50)[e����2�yp����ݍwב��7�4�j䊹i���;N.��/vZ���v.��^�t؏����)��|���8�6W7G!D�I RHL;Ξ���7��r���ܱ��Y�F�¦�۷E�4!�u2�n���r�nwv^-E��+��c��mj��2��n�[��S[Y:q]�k���7�q���>�o�\��V �A����"1`�*1�*�\�*�����2�sgw���﷭_�HȠ�R)��B���T=@yvo۲/���LRh�#w�Ծꓔ�����=Y�r_dޱ�Z�����)�E'>-��뭻J���6�-��ߩ�X�s��m-�=��k���܉_-�0���R�)��O���(����6��V'R@%$ײ�4�9�	��尕��v��ɮ�c~�W� :Z�����Y�`�IY��i��HWX�����&�{�����cio����#9�ӱɹ:�7z����������(e)!^�m��Y��]��&7�i�^�%h�Ѳ��4�d�1�*���^�z��m4n���i�vS����n���z.���$��𕣱��o3G\��;CڱiX��j����L��yF���t��S�����jf�*N������[��Bs�{����� ,��Ā��"d�q�}�u�͖,`��b�b
,�$�,A��:����s�3�>�TmmE�h -�*�y^TNg�{��t�z����O9����u�CS���e��x��V�K�q�I�v&/4��Wד�ݞ{�R����_}L�B~L�W�M���/��tr1���Ǘa���g-�����͈��k��}��QwR�2��Ε/t2-M}�4�{��$qk�����X��0l�"A�E!�0d!�o�I^�b��W�����ۭkS�����t]oMuGt;l^ciM��g������t�fU;��l��VA�{�FO#ޅ��:D�e���]C��o���X>�A-�.��q�v���}\v�'B��,� &NA��wi72�C�Q���Э�o����>��|q��	%�҈�HxS��k���,б{b1�
�@� ,Q`(�XF2
�E "� #"���X�y=���c��}޺�g��zi��ʜ�Z�k2R�:�:��>�A����.si�#�s��r�F͜�.��ؓ��՜3Ž��<\p�kMc����I�PV2L{=��tf�wU�b��+�|�@?q��AGj�OUVe˛{&ܪW��V7�_�q��#�q9?(�\y9T<�eCyz�����/;'w2�j���O8����*6��L��~KG��2>�L��ۥ�:8.����W��]s#�L]�݆������|�Ϝ|�g������:���sQ&�@�6��ecؿ��@�Kk����m���}���Y-�A�c�ԯO3����������z;��ʭ4+��ۣ�Sơ��Dt�ݡ�㖽H���r�+���*(�z���F��a��� |��`����5����p@��ў�u/cKjc^l���$��`�O��,E��>�7�ъ�＾��c�Uj�P��AQ��
�V3���o��k�^o��=���<c",�
d|O� ��c�{�KiW�uڌ��b��Z���H�'��y[5���q��;���w{�*i�$7үJ�N��ޔ8�n�[K�n��v�Y�ӳ.���vr��b��}z���>OL���l��&tk�*4�e֓�@�yB�.���1�����;���7e�\��宲ݕ����xex��~ T�]	��.��㌇�>3���I���:��j�����@���
cp��{��|*�ﻥ����]�ذ������q۵�#����Iv�Ǐ2|�_ʲ/��W���Ԩx
X(Ȓ
B2$�w�W9˧9�X�>بN�~$'Qw�L�I!�#������o���/�.��i6;>I������(�	�u�D"vRS���z�O;�bÅ�կ�紤D?��LƳ.Z�͹�_߮9��p�+����5e��Z5�y�!��L���o����{~ػ؜��wlz��2,f+3X�y��-H���" �$�a�o;�_3W���(�"2((�E0`�(g�IY�;uխ�ob~�Gf���{���[HNn��q{�ZÙ�{Ȁ=�Ȕ(��^�����������ݾ=c{9�Z��^�`���s�MmR<v�Q.��I�'�tS�[���;w¥W�q������p���'r�ѶD?0y�!�.�_m�yG���c�ٳ8���߿~�bzꠄ��D����4KcQ�So���V�I;��]b����.�L��g �%蛑T��K�����\Ɋ��������k��_o���L�a	�����{x@}��V�+h>Y�v8��06���Jы��֪�L����-D�EC��|�����J
��3ϼ�F�e��/�I�>?��H ��(��������k�{y;fV-�HVўӑ�]u�ҫte{3�Y�_��ҿ��������VR����%����L��i��S���{�^����ַ1X(�Ȋ"��V �`��^w��ƹ�<�9���2�ȉ&���4��w���m�>���fV��	������[���މb�8�3���}���:8���m}r�c���!�Ύ�Ҽ fw.6�z �Y��h�9Y�:P�*Ȃ��!���62�z�%KRz7;t��ˣ{�����`���sp��Q
2����5�����a
�z<�u�)���ǝ�(V�Aa
����Z�`@Gi��T�7�=�d=�SU��:��a��6|M��Kh ��:3�)�#`���B�4(4rfm*TŬ�]�+n�����C#:�g]
X��;�U�廹�͎���6��ʏ�t(���-���X�R�j�Ѯ.�M{EY<d�VРfM�������@b�k�*��}5��48Jz���r� ��)�P��'�^ݙs#��4'kxxۇ��3��N8�����[4�/�[���`� �6�f�d*��0Ղ����Mv������bVc���L&AY����YCwUH����h�t�%B����Ǖy����k4Yb�B&��oXq��U�1�UŊSB��E:�α���.�!%��)��D��.�F���EE��a3)Z��UJƮ��X�3��9�w#f7�Unzl*vQ>ɞ���
�F.]�9+Ui�)����ŷ�1���d$��Aw��F��V��kF$0����q��]y��]2�52$��N��H��z8�VZ�� 63~�5�`�t[Ҙ��]R�H;O��CÂp����ă�㸵4C@P��f�sv�8&�"Zɓ���w���&��B;�t�֓4���!/^��V-���e܋wn��]a���:�+�q]e�09�nvR���0z����&���l�KͭUv�rU�l��tw����-M����i�&嗂���6K�%�il�bbH�om�T9�N1���=8�K�2x����4)Ξ�J�����F_I�C��;����(�.�����޲��f��7��z{�]���B�N�6N�kE:䀸s`�h�N�ɫL����%R�8S���&^u�u"���-I��;��W�� 31.�񁻨T�f�6��>�;[��jq�Xn��]��3���%IW��r�7]��}����
R����g�˼�L��neؓ�nܳ=�X��������v��)�Fg�$�T�ȫ��Il�n͛w��gij�s�[��<�6�jw����|�^Dk��khpA��T��Zȏ��AKlX�C'dO�֫;u۱�m�T���۔�v�1����u�Kߓ�p���x~܇߅l�&�>5��}Q��i�u$T������Y�K6����y��J�)ޥ|��;W���)��8�>g�|��\�)gu���g�P���-ɧ���O�]	�����Z�x��<I[�֝�4�+]��6���Ĭ'�:�4�ğ$a7LdtE3Hl��s����#�Mv�KiG��O.��8D��nȩ�$ki`��S���Ww����8'�u�fv+��}��o��wxt�j�����s���6j��Yn����-�[rQg�u��b��^�䵴�#�iǶ����vYܖ�9K����{��k[����Ɩ1�ә�<��|��d��}QU(L$��J��6�Q[I���3�a�2 �|���^��=���~���e�����5�$L�����/�Ǳ����ʊ*Ȣ�PQb��DO�΋���Y���w��ߺ���1fJC��ִ;O&d�Fvv�y�磌��(��w�f��NY�<�ڋ��}���ȿ *{Bc��Eb܎,]�딟ov����lY��z��ë�[p+'�T��v��W�#Ao�$�pfo?7/S�tW��ѧ����k(���o):G���)���("�G���>0��U��*Y�bJD�ҽ3���H�A�d�A9�=М�4�����C��k�65��%0 �R
��i��0�}ش�v�e�Փ%4�327X��}W �]SIr���iֻ}k0�4N	��lU�~�����0}�]@�,�uD	�~v�ʿ���W�,�B���#=��Sv�����{@S���=�.P��G������Uor~���^�,�Եw�uk��ҟ�Q�A��ح��ʖͻOZ�f�9��Y���~��>n�}�瘮2W"L�g��mV锽%Gx4����[�{�9y�y�=�j["�` �A �1_x ��uͣ�_�OĞ�`u�mPיXL�0��fvv���&$�eZ��D�������DI��R�rW���cT���F�ݻ�zb�o�X�\�� >�]�%�|��؇����=��%�8����_R̗^KB��P�,ew�}-j�����Ȫ�k~��q�N�u��8xe�x����Z�$�{����+��&���7���Ec
�� ���E��߷������{���m��L0�mS���<n�i=�: 4�>���H����ۈ��Lk0h�����-�"�eڋV���FD�E��>]�6����<l�{��>���ۏ^�1��|n���{���P"��[��1����������b�%
��궹��M��O_fS��ut��Z� \�/6WC�z2����d{y��Z�w��}qi@N@?a"_O���(������w(#.��Ӭ�ŒJ���4��"��荦�
M�ϯ�Ā`��X��"��깞�ٯ����|+�i�y��o��>����3��,
�m�4�v`��H��h���:~qnO�oIO��{I��OeR��떘���M����_~���>7�n?���D�s��5b������ã�#ww��H�����ߢ�M?�|�N�Ai�k����a:��0��Ո����
 �0TdUY���X
��j�o�s>�s�c����� ,�@�Dl���/���Nnʖ�3�At�N��K���b�=]Qe���0C$u���������Q�������*`鸠̔/L��'�3������A��}���ϡC�t��`7z�� ���Ȕ��6��z��湅��W�	s��p���>��@URXv�T����vZ8���N���vodWZ\v�q�a�h�٦Eٍ�ˀe��)�'�5� �o�<��"��_�+n��^���\�o5)�ㇷZ]�-��i�F\J��=W� (0�$"Ȳ5���z�\}t�|r�v�v�����+�T%��/�G�B:ivD�_H�sP�F���ܡd��Ｉg��p��?�t�r�`l�m։љ*�jz�>�Qm�^�Ҕ�����1g��ԧē}��A=[R�otp�kgjǭ�ǽk��Z�rr��r|]�Ͻ,�e��#���kn>,j���Sj���S�6���)|.3�:�sw��qF	�u�r�0H�X�韺G�(���W�nO�c|�H��E����HȊ
�0E.|���>��p��jtͦJYl�'�:�w`<2R��Qc��ܗ&���Ü�mu,�+5��Oy]3c��f�t�|=��)��s'�s[�������/��!�+'�.��`��⌖p��8�!�G���:�5�\g���-X��>z+|˶k�瘺/k2���y�y�W�o"*(�Eb;iUG�EԦ+��PUAEA�(� �X�)�e� �5V�QJ�bȊ����<�򮭼��9ܵ�^�Ww��WzA{�L��,ݬ4��K�o{��S��aYN5�.��l�ڕ�0��}A�j��3�j�Vl^f�nlތ��_{�V���|@ ֢����ؾ����d�Jed�O�����rqɁ�B2<=�-z�<�@:Z/�d�h��lʪ����tʈu��t��(�::
��,��IS�ur>��C��_b��?u��9��{���ٺ�T9�2��	�2p��g?�f�e�%J��s2�N音t��T�T�]�a���Ĕ~�u���y��;���id�T� +@��{�TH���V,c���E��}�}]�{�>�Q3���R�=�^�PGĽ��#5E�F1ֶ3ӣ���*�֕*j�6�G4�.$��j:+i��l�̬;Xn{��G��$��g�x�6�N/���J��?����1�-+�IΈ�S�s��6S�_B.�|����j�Y.*��{r�����@y�4�EN��]���8M9�U�I+�~����߼�e��������#�X> �=�HS ,� >��1��o��i�o���͒X�.���ø�N�L�Pٛ�IOH#2��3��\��sF���n�}��e_l��حΗ.���tN�l7D3��֝�;�I�g�|�W��e��e�u����⒍�%����:B�o��C4�0�n'z�E|�/�C��T_o_��3�(�裵[E������l��U�겗����d��|������ݡ�v�)����-�����\e���<=@ (P��D��`��"�,�DdF
H*���ך�n���7w�b�Q$�>@@dD�	�o4V���}�u}��NZY:b�B95�n�w8r�#I��Rũ���h�oەCI��v��).O7d��j`J-��[�UJ�7�]O�߿y)�)�wi����!��Y6�����=W�|���O@�7M�}�򠧹\R#�����9��3Yg5��esT0C�+�G�����}��_�Hj �H�"��
����m���}��u��tNS�I�bv,�O%��Ф&�� o�[���=�}}���� ���s^��Ʒl�,�/zi���!z�EiaeS����}�)0�����uㅖ.�`��]�-��wXKhg5a�Ԃ'��}Ku�>���O�X��O]����?dU[w��!P�PI%\�n��������I+�Lw+����M+e��hܞ�+�L���,�!�
5m�[�����V׫=��&�%|���rڀ8�����7�0!��D����^�����1��X����� �TUEPR(�����z��V�����|���a3�|ޞ��s��!鲶�O��X��W��voE;�z�b�u<!8�����gv��NwL�x��<x��uF���_l�<�D>6���`���8m�����/e��K�}��3�u鮪��^r:������亚H��]G���ՕṠ����������x����g~�ϛ�'���h���Ō��f&�,�꾍�YWB<�q�[O����2���S��D�F�>:/�ίUU1^�^����b����Ysvc����^^���u{qU�5��w�:*:}��������5�b�V�_8e���-�(]�)\K����ѭ�=�E��,.u� V��R��|(��x��k:n������:�j�e��d���Zd�ݯD����}�X���h�>ճ�[<w��KCݪ�{ݹ���@�Jţ�������� �R"�)� (���, �F"("�*��H�����;�뛄OD})Ȝ�3��V/NݬF�ʮ�����A�}����ڹ�P9TC�D�"Y�af'�#;M���W�^Gn���}���M�O��x>U�������=1B��ߏ8��I	�k��uP�{d�/U=�ܾ���Ԇ��(�T@u�}V�m@�Pd�f�{�}�7��ga�@�Ҳ��	3�L.�� >�`,�RA��I������/��V<R��}�ۓ����j�_S�1F2�W��������uօ�:ڔ�m6���\{'�u�.��c��U�	m�{HF�OuP�w߽��~���+���������kD��s����e7��:�nk��e�.��9
 !63X�[����*�}��N�H�z.����O_�r��qvW>�Nڒ��]��lQ���V�z�G��Q���8�L^-�w:s�*�>kk�g��+��E�Xw�}���]������#I4A��.Ɇ"
)A��(�1AH��H**���}�9�o~��\�<su��]<�h��"������F�w�7������\�c^��_b|��#�,x{7���ʬ�lj�j:xb���y-�Kc�@�krJ��\��۴m޹�7�C���5�Y�"��S�&Χ���ޟ��cv�7���?K]l���z���y�36�/��l{*�ٹ�l鴅�<��M��ӶGl�]w&��]�������!��"�
7����{��s[��gcb����� j��G������c�0gB�R�g8�R����`I��JM�Skӷh�c�[�='m���]�����G�t�i}�Aw�P?B���;��T�1�6k�[O��s��2�#� ��}�90>X�.9�ө|6 ���|< �	�����z�&���kv��kqK��L����뉱 ',�}���Mk[�w]+��7�ՙ�v1U��R(R��_>n�y���Khe��m���>��"Y�I���5hx&��ZbeAF�����N����c��?V�U��̪����U�V>�����S���ԯ�:�����ؤUF*�0�)�B�H�
@D�`�\��g�zz�J��I�^Q���8�݅�[�@̪�����A��c=�;'lD�ּ��1k�����ء8N#87Kvd=������/v���|����:g+ϝ�<4m��9)��@�CV�����ԡ�	���1�UG���P絏���Q�a{y�v�S����%(�����x���}삄lv_����U���r��_J�Dڃ�\Ζ���_�xyd�_eޣtX��i��Σ�j�zE=*p��NMI�wtRC7���<	�8��Vӟ��8�wk��މ�dUǍ&��n(I�<�"��oj�1�˱��C����8)�Cƨ�F��EG�.����k���ZA� xQ�V��j�SCם�2Ul̩���J���[���Xls�d�)��ǐ�v3�7���%��n��)m��Lsq���������5��ۑ��ڀ�z�F�jK��@����E�Duc2��D5J�ًX�< �l6[�4]�c(�L���8�c��#��^p>�+���4
�L��9����)��U��$���@��@8uN�%AJAs�P[�*^l�̠��9�a^��b��C��~bl��c�i��^���t�uJ����qӎ�f�@k�H�L��9����7����o���%Qu�z+E�[:�X������FPy8�+>����$	�h�OYK�8�Q�E���X�`��Go�Hq�MʕT*��&�l����{�K
��D���ӓ�j:d�D�(��n˳	IZJ&UCCT�?*	�a�ˀ���(�a���l�hVf�x�wh��"j�%wt(UDʙ�����Nd���u^+�g�~�EW��,��KsQ��DI5����tk��CLcQC++��������F�����B�`o1��w/]���y�6҂G��ZJ�¦c�T�6�i7~�����3u[(��sM�}��M<
��!�n�� Z���Y�mQ����㎏us���mx���f>G�ɝV��f�}G85�������4Հ.����%Q����k�{���������UŐmެVdgAg�r����[d����,�ŕy�[`^e���[�ڻKa|(o��y��n���+^8ow��WޚyBA��S.��!DRkgP��Ǹ:�Rb$1!nw^���``:���,�u��y��M�FM�tm|~�G�35sRc��v%_U���l�l�RU��v���38��+x�|����-X���Tk��v���}}��̥�w\�t�����T Ɗ�(�]��Gg�][����X�Wc.0%iH�4�94�c.\"2b�|�G<[�)gv���"�&cjV��-�V	B_��r���\���6�[�e�YQ�+�.�[=�B5�)q�W�WsKv��í��*U���R�w�n�K*V��!೏2&<:7�Ue^���u\K����7��Qw�@Y�KNl��˖�
�);���U�!ݾu��J���4˓Sty$4TT��j+gF�:�dv�iȶ�d�CĮ�Ԫ�,�%���n�tNm��{B��f.�x���,a�9�N�+��Rok[�K������r��VmqV����pG��>c� �49�\᱑H(���#|Ќn������q9\励o��2��Ȋ�wUd��>���gC����at�����9'�=]�z������[�"�~����j�V^��+���*�Fʋ\.<���3�{&L�9u��n�u҆f����^���P�o.|�D���k�v�QT,,V�J�� '��� {8�'�#1d���w��"�*�"��X�ET���q��e}Z��\Ir�+�|,K���;kԒ�Rh�eT=��	��{E]w2E��nւ.�$�F{|}&y�Z!�V��2b�\��5�ߎq��|�d��Ҿ�MG�ш���bJ�`N�i�ɛS�N���zUN�hf:�����]T.ڋ?W��\͘��o����Q��ܚ��e�U(���3�;���
# DP�T,�����/S��M������ᇠ�u���D50���RU���If_*(�{w�c}�7-�E���{��v��p������}���}���q�佮Ȩ��?>3'����B0#�*�7��U����X��=[�pi�l���%-���N�1L�W" LG��[L y�~�c���$b ��$PQ�AF*+2,��Gп�,�$\��[}᳖�;f��0R��[iΗ�c�݊��幙n*f���
�Nov薶s*F�M��������nO
j������|@A�ȤQdA�,�AA�>�ZK�~��䟮��]P2P�J�n�]�jp|��a��N�^y�T�2d����`h��]��rv	���-��!�m�l���H�U������/��+���X��M�ѷ*�!oOP�^�嵺RjwUV�Xݗ	�p��SN�������=i�˱�v;LG}��%z�l������P�ݕ����O�$Qd Ͼ�~�q�ec�'�%���{U �oM�Y��\�ٺ��:�En�[�̚��>��W'�e<���r�3)���^�0��?��F��q�>����ʉm�8�#��7���l}[u#컹mL�e�;�c�;��J��=�9#�if����Q�O��/����N�wq}��� ��ʗv�o#��T��lJ�KŰ�/��? b����������M�)���R
DdDF1b�QY1#() �H0D�� �H�DXwX�.��vٙ���֮K0=�p�ͫ�h�N����a�M^y�s���E�{�p�s��f�eyik��GyP�S�[������^���M��ƪx8�R�rK)`����h�X�0I.��%d{�y�Q����k��Z����aө�sc��]Z�����Kӱz���fWQ�ϰ��t����,e�5�`#��a.$9j��h�OY�'��*�/hx}i���8um%���x_R`s��wr����;i_#�.�@Ǻ�D|�D�TjUE�2�S#EI
H�(��c:���7)��p�w��c�=^����Om\��-���y[�p��WY�d4!a�R���NN}�|�`lW��Br|�^��WQ�Ҿ���{m@_ٹ�$�г;g����{�� ZV5Ջ'����#�u�Ԥ���e�]�7���{��Lq�Ҕ\w�kC	�����uAibQ��,�~N�{�C8���$D�EDF
��*1 ER(� ��2 �P�$�E�"�T�ă�Y�{��}�|�o׷[�O*h�W�ܖ	��e�ţ�g�8�����D��3R�Q����eN3Fv;�ܙݰ,P��iݖ:��6,D6�u2�R]]���Y\��#�8�^>Ѿ����{Yo���s��8�*��>}w�蕬}̳��Cηp"ٙ[u���~F�`ـ�7Ԡ>|����S������'��Xͫ)7X����?f�ҩ���Ni�j�d]C}J����?�bK�� }�,7�2��䓓�ի�rk00��8W+��?xP> @'������	�Kcz�tA��{��|��<}��Ԧ�)nb`n2U`^�(Z`0ʀrME�}n�Q9=5OZmW��>$���V����V�oƸ[�i+���Ҿ���~��U���挺�!�d�O1l��U�mZ��^mĮ��qC�>^�P:���[Ők�Y�J�I=�V@'�$+"�T����,"��E`*��=�g�+=߫��-�l��ݵ�zBeY$/�ո�p�#���	�a֖�l`��AX���*�\$��9t���Gb}7�Ժk��{n�}�����| >�36�:���x�G�-���k�z�)Q�2tKx��J�{�i�t����\�ˍy��Î"�K-.�O��R�#L�F8�� w7F�������9=>&}�v�ܝ���{Iŉ��t MH�7�@6H�h����!���rOn>���gwn�R���7X|}֗6'n6��S�O)��� ,��s����_}�N��UR�ږR���	�j �0�����̻���9�U<�?����~]�f����v�Tu@	|`eg��&��Iu ��zl;=�w߿]}k��~3^���O�_��c͌����_q��y�&�dYFgj"9��F��c�1��N����)�o>DN��V�M�nN�\$�C����>'� ���=U�ߵO����Q���DTF(�`�	��A���"N�-�3��L{ݺ߹w���pwgBo�u%wLfrU#�~L�7:���ˌ½d�1�FS�C�Q��U\������󃵚������L�H<������}�/t}f~�l��"�L�ٵw��mE`�W�������F����[��ˤ�q�#%$�)^n�A>י�;e��{S,�����P��~�}�Kz��rp���E÷A��K�R�X�b�8��,��zˑ�E����ׇ� ��8�|dY�kk�fʷS�����}��j�x��(0d$�Q��s��^W�7�ܪ����J��A��el[䯬oK[=4P�i�Ӂn�V"KP�(Qx_��3É��p��f��6��}i�_�>���@>u��-�{�f�J"p����Qn�&���7����v�p��^�O%U;L�rM,:���nK��c[��O�����m�)�����6�Vp�Ø�8���8��뷙,D�F*�*1XE���QF("�E�H�
1 ��F"
ם{Ϫ&]��4�{��
Ȑ��cC?+��+�(�*v]�i:pˑ���+7sa�M���7�z$�'�3p;`G�9�5j/
�weG*C�ޜ�2� �q�6�B�+븲�|�n���rGo9�1��-`����	^���&�c;絰}���G*Uܪ�7qnv>X��7Yv�d�QI��q8��3V`т$`H7צ�F�<9��Jguf�8��is��,��T��,�!��7j�ՙ����B�&whQd��J��y1��h����O�B�o$�19?�~��C���v���ʬ�>�L�k߳�qUj�:;���1�H�iqb�,&_Z��:�W������Υj̴Jdf��LA�Q�Cm(����|�</��oג6S{��N���!�G���qX��gPO�ǃ�)[ʁ2�v��iS�;����3��:�wN�1�jW�3ei&��&�rW��X��)b$QF
��QX# P�w�y�5�i���7�4��Ra������b5�әW��� %�t���n�Osv�x�Y��\�t=ԙ��U`�K��]�6��om��u|�:S�0$w*
�r�`�7�3��?~��R䔨� ����w3W��W��vD�֌�%�9�)7Q�����F��h_|X��<pק�U�b�W��}��,�&q525�k��:������U�ukip��P�潬���\�"D��"���pʜ�ض��2�]�[ӤO~u�L��4�Ȉ�r,��o�Et����/���&�{�+�޽�����$�� $��{���^��W`���g�e��M���e�j�����D��(�u��J�OF����Hp�KC6�]iDJ6;J����N9���5R�{�p]����'�>�O�}��������0m3�#͖��r8�V@�KO��$9��:��k�\�Z2�����f#S:��N!��:�ۿg�_oݭW�j�*�*��aDIHT�A$��`� Jв+=�tW�Í/����X�F0�$`��E���@${��?wu�L]�ָFm%k��F���:>�3� ���~�a	�ز�L̒�zcK4�J��Y��l�2$��u4U��X�;)nK%O�?����&w���������U+��6�$�('�T9�q�x��ts9x��ZJ�b&����T�1��خ�ZЅ�6���]���3��/������6Y¶LhK����9�tn���}qf��w����S�ʗy7���av�ӏ3��ޮ�pM�+�����^��w��]�_�.�y �*D���fnCX���b/U��[G�Sas���@7"��Ψ��`�y���!݊��G*�+��$;���J��H;�����?,��ֽ$
��������X0'{7����S�ҴڀB���c�{��ȝ��u��[^��ks,�1DzZ�D��.������a�x�s4f��w�H"#UIQV �V,`*�"���PbF2X)"��QPA�(��0c����F ����+�=�w�O���������3B�uK���~�˕�e�޳A���z��Q���'�Q��	�U+ݤ�<9�P�Ηvk=��7r�D��v��nb6cG��~?�+SO���� u��t��]pd�ə�Y�32�^Qu��O�<K�>�SĶt�_��
q������Q&,�"�.W L�������K�@���b���"��"�.*�X��5)�*�"#H H$"�2)�T����P��~��5�Y��B�����3�liLm(�<��t���`ob�̡�b���s"uҕ�/������Ӹ	;�e+&Y�V���MߩH��D��u�����6\���@���g&��3V�Xɔ1X��{�R�������|�_MtA�6{�͝Ԗ9���m���jn��q��f�$�����򪃪-��(�h8�I�
񚴭���*A����b,EQ�+QA�F ��H$H��b�A�Df9�wOq;�����)��x�[$� ��� P$̒=�:�����?f�u�X�{��<�Y�[����Y�/w~\�ˈ��:��b��l��їB�W���=?}���/��u��s�j�צ8�$<+����Zb�_�׮�}�(m��s:�Jնx�<g\��QL>�r�	�S�m�/�;do�q�����d�+ӌt�,��4�weS[�g�g�wU��ٻ���s������� ��#�P~���ksu�k�Gj��:���1d޾!$p�� n����Q}4ScL�`�iN�n�� h�&۬�j{�YWZ-�"��� e���1Q�xL�
Q�O�.c�X���Zk#;P�B�ҩx��G�Yۺ�^��j��(����с������5��*���}K��]yG�槵p���l�d�$6�P/V�6bnu���V7&d8�]
 a�|V����ZU��ר��7�(V*t���@��V��6,�s��w"��ޡkM��E�լ���2��j��J���(zM���78�[Dʞ7��@:p���Z��v=@K�0NU�q��Jcս�t�D1e��s㴵I���P�m��2�%�Q�\�=@p�<���F��H����R�7y�7.�s�(��R��g��&}�u7{+V︽�]���;��gŖ��w�s6�`�#T�AJ�T�R!
V�F��7��\-�!Y��j�U�A2kȤ�t-��m�"�UI Bf�ST�W[t]ڪm'M�t��1��Ⳝ�PÉ���@d�@D��U��t-k�ʭ0jJkXlU
5�xrN�i�Y�C��i����b���Z)p��x�^L�%��qU�bϩФF�{D����Aus 9؟�t�eSu�)
��V[�H�wU��Y�oYM��4�0�$�(�
An�]�oMd1����hG�3ى!�[����FL�7l�&�Y�Uh���)�V��(��طu3�fZsP�XWaҥżv�ܜ�_
=�j���z�[�Y�E:1�}#�.��p��d{pC��q;<0^�it9a���G�������
�cE6�T�6; �7j�Ny�
F.�e�H��x8*}�����Y/��	���Ɏ!u�W-G�l�ب�yswC��pm�eKe�k��9��%󚸬���(��d��r�/t-s)��f����	����P�s	����k�jVH�3{°�f�%�䣇Gպ�ma{�Ũ<9!=I��K�o�g��낔�Ft�Y|-��U�.x���$�Od7�V4�&�[[B_(*�f��u;ښ��.Y�5�VVAIHȜ;u�����SֻOlZ�W�(Ǔ����(+IV�ʗ�0Փ�2�A�5� POvpWQ��+����r��tE�_��|K�gk�GoiU���M��	]�tĞZ�S6�#=�n{�e�U�6��y��-�w���^U��s�h�z�p\��_��U�to����*��[qM�x5�)ͱ.Y�V�f�e��޹ժ�	.�����S�^�w5���t�}qS�k���.��N�И���ڹ*f�����í�+�P����9�6�J��s'[D�\�aempҫC�ᴏ^��1v�CH�z�	{k�
u��X����������.}m�Z��lJ���b3#CK��j".h0�
-�ˬ�`綣f�	cQ�SQ�s�W���0c�|����co�߱�M���Jo9F�<�zz��&����G/[BmJ�2��f�G.i:8'y�be�ҩ��LǗݭ�nJ��� FER}��A��;�g��,��ԗ�7ܻ���(��ً'��wcIk�u��{׾������Z�ow*U��۴Ӝ���A�>;�r��2�X�r�ΖT�^�y�v/%+�Q7�z����,��[�\{�U]uT��v�k�՚� n"2*
�U�Ogf̞��k;h�F
@c""Tb� ��P������=���3R�j=��@ަ�	�T×��&xM'8c���q��:��J�)�S?RH}=�Δ�dND��%K�?^�6�A쿇������}�����j�T$rW̑�4�d���$LP�r�O>��x��yFV�+�/dH�KN.[m1d����&�ۧ�3�pƻ�\�b�u*j�x�'�ze���(��>�z�|� ]�xz��q�g�p�̗f����8n�,R7^5U�v�W��y�K`G��G��>7��a���L�ݴ֫�}�[�sG��9Ko:�X��Ɂ��#췷g�,t��ce>�;���]��(VV�mV���o��j;��k9|<����G2��y��)�� �_bG�OOg���Gm��}Ұ�7�.wU#|x�qd9��K�m:#��m��7L���/���՜`�3��K2։��g��AIV1VAEAf3�w��w�8����:{�:�"$*��, $`�g�Wv�VW��<ϱ�vW��PR�Y�p�E񡚓���;�͖�o7Y��y_��u$/��.������vv�ݖ0f{v����z�5����i
���JV�\9XxBA���m������%=�:�_Z��tƒ�C���)��)��,����y�s���ry)[�%�--ۯA�̍es���X��@>���5��g������������jd��A/*3T��-�!����/n^>z�^��u��q�fg��(��L죶��U	��v��/�;"��a��2�\�კ��������N����W]8�b�8�̴Ԋͪ�Լd d�������	� S���5�xu�����S�����Ks�����\�s?}S&�\�,bG�U�f�Pw�g&>�R���]��Qg������!Q]�n��wu�^c�ÝH�, ���Y�$ *�bȑ9�f���w;�];}}گ]��q� A)
A�{9�}��]�^�+z��Ȗ��?$v��qlz�;�ioB�uC�`u�w�f}.Ȱ1(/��$��뼷T�~2d�yJ�B�X�|�b��߶�zi��H�nk��>�D��x��`�XivxgX:jM�&�̥��I:@����w~]�":�؅3-gK+y�2�0��\�v��ܼ��{��$��A>�����}X�,�Oݖ�$Ϫ���M�t��͉=��1�x���T<Χ��ܥ@8��o�i�����N����yj�gkf[=�B��j�TR.�����=�#���T�L���*= ��մ&���R-왂�u���lU�|�b���uқv��G/)ktuWuS����^�{!�S̰���~���ͮ.��0"��ob�2���{�̫��[X||��^��wc2�c+�Ú�QV�&���:�q1�s���"^���� =�Y�ﾾ"�*$Y#��� �( ��5�ϻ��J���0�:�!̨��C:Ҟ7qA�|N�}n�˫�鋔���@�.��,��Ih��C�h��U[&�����H�+���ߧ�<���1Z3~��N���$g��zD�(֭wZ�fd�mD}�����#4�WLLŕJ��y-��6=:��H�/g@�5����?�|���y��u=-K��?�ws�VR�/E(j`�u �LQ�C��fq�ȫ�Z�f^��&Z}j紳xm�H���������Q}�ﯰ��|5\�o���D8QӅ�ߗ!�[Ja�F��zS�W�E�㵃}\=U�W��뺘�%ӽ��揈��#��ڼ��U4n.E,���X���T�5a��T��N��q�iu46步��f*e�k�2u�}��u��,R�����XC_�r���se�R)"$�#1F1���j��׊���;�{�Ʊ@Bsv���}����F��Z�|֭��-�v9�9T#��O���;�7szߺK4��S=���ԧZ�8�{��9�`\�suJ#}^�]����M���KҞ;�-5������}%W�iFa/�Ri{*�f'&�����pӖ�p��᧖ܭ�S��geBe�zO�eOss7]�Q��uCq"�9c9{��0�jj�� ��F0`d�,�9^�>][PM�<T
��;�o��Y�'B�Z�!�]P�ң��gn�^Kvגu/h�^�R�Rz��M���q��g�Y�}}{X���f��{"�/#nun������S?
���_=��Ϡ���lW\�zfb"��T�}�|��o����!����w����?����R��9����4�(B"�dUX
(�"�PU�ň�bE�DF0EQ��+DV�����"�d�EY
�(�D�0Tc�B�K�&�����9[�T:w���B�
�9\���/��R婚u��>k��\x�9�-%��2=�;����|�w�/�7�[/.����S˺{�L�`�5��}��x�Q/çuX�Ճ{����98�Ww�Gkt��U�"�K����P)n�2��wl�d��V']�d�i:��:kgb"��\J���>��,���*���]?gy�lAv���s ��v�c�!�0�GaL ���v��46�\Vsb�k�)։5ff�S���b�f��3	r��&��ު�;=���Ϣ9��TN&�u�'�"u)�JU`�Ov5�y�ފ��{�J#9�Qm��1\tK��+Н֙zi3:�i�͒������-�}�Ǿ���|i���/��{�t���v�:on���4�ʓ#Z��N�m�#��K����8�M�p��O\�gnK�WMHv�Z�,z��ppڝ�/���� 3�G�m����"(�c���cDQ@X�`���2� �QTEc"�F+*�(���Q��D�?gu}ʪb^�aƝq�ex*�ָ�����sw�	�b�ݭ�`�S[4�e,Y)�ض�T�q�&�r�wXM��e���)�=�Io���qІ��[���m!����g�f�щs��t7I�^��M(G����|�v���w=�huJ����ܕfe���8+�E嵶SK�I:&�s�3 &M]E�B)m�5ooO+���f����.��ۖ��@[�9�?�v��y��K�6�&��\\v]Ŷ�Wr����>��H�0��>(kk��Ko:�q�{��f4E���JO��u���4��� #%BO4 ܬ��9K�R�0�C�<��v����=iM'����U&��O��?�L1�H4ʀ^�5;^;Ҽ�
�i'�	Y/��v��G8ۗx(G�`�sPeTM@��&^bh�:�=x*���(��b� X���DDQ����3����^�b��k}�=�Vm�E"	 "� ��������F>6��'mi�z��Sk!Ф׵�z�z�����hΟ<Yx��f�/��,{i����ѕ'm�|���k�l��-�ֽ�|�� �ڋ(;�+�*�.��.J�c^�O�&��9t��'�J���j�\C�<߮�澇�Zvy��wt�Ls�:^\(.�©%�K������{hԱ�s�j_׮F�=3`�N�R���>��aa=wX۬����Y��~us��Wp����c�rס�D��@7*Z�Ԓd�U`��4g~�n��.��rg_��h�h���YrT��~q$��Gmq>��>�]���U�zv�Z*b���}`t<�V�t�:��� q�nPۑL���%�L�|u��P���^���j���n҉�gZW�dv�Ϥq�gW�S��q.���iyݫ'�fV�%-���>��]�5�<�=���|��nַ�=u�V� dX��R��Qc,g�k�v���ի���E��^`tT��DH��DA ?{��={��s�����K�ף�t)����~̽mfKl?{��S�;n�|3��$i/��]qPj�k����3	Dc�s����R�������|���W�$��wȪ�D��N��J�R[�͋�I�.�9 ��mG�C�������,ʁA�N]�7�}5���.�/b�HF�З��/�XuPpgC&И�y^��-��^�*W�2�,�!�� 6*~J��S���T���b٨������!{
􉚦�������OvJ���߯z�<�c�3,��Ƴ���Fl�#)��&Ui�&#��Ix6��U����'�u�,;�+`;9n���[����<�&"��t��nL��MM�8y���Hh�.>5:�u�lԇ��D�W@}M����u���x�J���h���b龁�nd�c}���}�8�;���TR*A�A��H�X���B"���������=}���1����:b�f�y��ݵ��4���R��k�K�AC'�;�W�ܤ��#C5F�և
Ӕi�Q����+�^�W�J�/�C�mlVGK-K�\��F������d����A�t���^�J��J������#6	�oXf�m�wN�\�ݲ�R�pR�s=f�<�����r`F;��k\%�U�1ngv]��v�<5���(m��d;�>=;*�]��/*�&M)-8�>�����W��;w��=���˽w�"���P�{�½᱀x���kDĦ��D��m�#\�B}�^T�Nx-�jB>j���S��/���)&��J^׈ٺ��G���s/�U���{�
ڷg�0�'���G�g�x����gn�cx���0��s���Iu�rT��֠P�J#y[���by��g!��'V�~�b��� �B1����������(*"�1�UA
	f}��ü犾{�Z�/�� d��	O}����wֶ�~�(��n�8�i�"�^�3]Iݎ��� �yht5�z�G|<��܈�8L��ب¹Cj������sC�$Lڽ���\vG�ͭ�����e2O�$�����c���M><m���t�	t�"�Av��p����f�n�ڊռ�W9�ә9Y/��5��U�UD�+�Td*Z�f�B�bf��F��'���J�-z���L��$Q�n�=SuV7[i�7
��)�Iݣ������'y0=V�]b �@�p���TT%hy���YF��v�c��o���&-����Ƹe>֦J\�^���:�3k��y�k�X�+8:7YYH�WV���i+:����`nO�RH�1Պ"�f��DTC�`a�B�+����ta��|���c4��ײ]YJ¥�6��j�pK�Mk�,���nkue�n]i�u����T���op8�9�M�V]�W2:��e��k9��AD�Jh |�!����M]�;�'j��%��bR$$�(^-0�ͨ�@�7*�U6��Д",i�����k	��TQbz����W}���E�cKz�����m��P�qZ��VW$)�5K�Q x��v���t�D��z��}��0`������(�K\f����v1��W�����ܚ37�^B�e��]���������Q���x��d�{UM�qT��ņ��C�T|��B��X(����z�}(�䉺��}rpc,d��rK�[����]0^�*-��U��2oR]�M�3���Q�%��;xmL����)����1bA���@n���.���<M<����ظ����xA�� �wB�Q8Ȣ�!Fs�|�sQͳܩ\
�2��V��<����'t���n���{�'������j:��#�MY��#��Y�s�l�;O#x��^�:�&��+��8�P��Xj��mM�Ɂ݇x�}���[Q0��\���ta��U��fk�e/=�2W>q�.T;������M�$t]31'.Op�3G����˾=�V+gx�]�eD*�@�	�U�Ĵ���VP�v�ib�l�!ɵe62��/�G��[L�H�KN�f�m*��A˰�����t��LavQ�37�<�\��	�n��ݝ+NR���T0c��5\�I�qй��i�(բ�wp[zi��c3�m����Φ�\iU��jw[+��C��39�]�]ǹ�\�s90�q.�^���c$�Ur�j��ĩ�r�ġ���jV�[B*�4�����Z�j���:���v�*_QrQ� �CXj�a�.�$��e�ձp)�vn��pn���1�E��t8��Go��52�&T�K�*�g]<�R+�ĭ�J�\-��)�:*fh�$��ج��+�8������7�JX��:�P��{��y��ٜ�L� �v�e\u(:JM����jқ���<kU=חZh���m�[�7{m8�uj�ǻ��y�un���ײ�����/��*��ǵ	�o�C���"��A�e힦w-�N
w?b����n�.I��qv�tc�Dmh�{v&�}9��tMոH��&���l/3�����~�Q[����6_F��^EX+�P�:��6��HZi��x�w�߽�p�F����,�ׁI;����<g�%�� �P�\Go�W�7Z2�v��
�؝S�Z��D��h�Ρ��#*�廒�3�i�gc�{��$�^]J��Ͻ]�#�`ľߌ�
br�C�T0�U��O�TS-Č�:$!n�J-Ԟ�-'ݗ��bBߏI�V��3��_T�S�l�NI���N�O��=��݄�J�Y�����j���P�T@QT*��"����oZ�w�޽~7ʠeӖE�iL�xFy/C�I!Ҍ��T����jpEL���챗vd�whikP���f�AkW��͂ܽ��'��k��Ұ�mnҼ�J��Z��^��8�������ʗï"�u�o�g�)|�P� �f)�W���{|Z�B"d�6T��s�!��ڟ)Ӻ0Ьz=�����v2bٍ�x'�rήW�]>��3����[C�i�{�x�Ժ[uRI�z�@�?~���x�� z>O��>��/~;l�U*���w\���eD�$F?� lnA������K���9zw�亂jx<G��n(�B4�e 9�x��H*��<�j�H^^,$v-㊒1��<Kje��CA�zzZ.S�:W��}A��+#��<:�%�%b�\����_jޜ��ݒL�D��R��[��Q�ERDa�U ��׽�9��^��J��i�P,2�4�����n�� �\3%[�*z�A�����J��\Λ~��G�dw^�Դ4�C6�����=����#�V��`��[�WF^�\iJ���g�{VZ�.������Y޻���J�g��O�[��.U���{5��1��@, E���:n��+���KVQ!;��#���9��2{�t��M�d�&�����E�UK=L��-ѹZ��O������r�^��Z�w���r��%GY�Ũ~�� ���������1�������V��+��-Jp��xh��wMm�Y2Ϟ�	����n,��K:�\�Y�R��;a�ꇡ���)k8�"nfYo)C�yDu|����i^�$q{���bJ8�t*���Iy�7(ך�{�zR�뾈%�D�CI��Ԏ���!$#&5��<?�����()E��bA����I�Ӿl��1�������7V�ߞ{�N�|U_{�DcĄ�J̛x��$�짆e�U�2����u�����R�`tUML�wvWh̒g%F&k�{Ή;�"Q�2�faZo�~z<HM��	����6�^��q��
�����������1-ՄZZi�'����(ؗr�sca���8��׽�s�F<;H��Λt�u&k��ut3p	(�1`�*
�(�DUP@U�"(�"�-PR"

��F�T�R�E��
*�+�[F#"#TT`�(�Eb*ł�H
"�b�X������U�(���{�6��Md���
�ЎQ�r�wi�N�xn����e��l�t�lQ���ȃ��8��-+�Yү6u	����c���we���c�'��w�L ru4�32q�>����g�'�+ ���ܞ��i�8�b�/	���<�Q�ׅ�U���C��֒����&��>n���/F�n4�S�E�u��up�J"���^V�3�3M�C؃.0�w��n������.����Q�UUΞ��sGWK|��­�0��խ�z���E��D�Z�]��:R�X2
,AE@Q��$E�c�����y�5���즷+ud���ݕ�s����[C׀�:�uz��G=f�^�K�_�/j����a|��G�j�s�W��:応/�vc�nЎ�!�|�;�"�D��Uq���j=j��o]�';�u^DBuU(��8���F�>H���M�\`����`��W=�pМ���R�[Ԛ@H(��� �"0�o$�y�^�M�4Hϗ��MD4�r��� ��s�{}��u�����U��6�w�Y��YD���O%�w���ՙ��R�뤧� ]-��a���t/������ۮm)ں���Ce�����	|p��5iz���F��@��\�'s���h	G2�.	"��Lf�^˝F�C�e��A�#sGl�.�?@-��mK@q�o�����V�k�Q��Z�F�^��]��R��
�$rU>i̞,j�]ZX�۹1w�fĈ1����dY � �7���̈#E�`�� � �7Z��\�*�d�;)%�A�3ڈl�A��Ǆf6R���蜳��w-%�u�3˕�.�׉�)�x3�j�kۮ��m���;gah�rG�u%��=1[$[!�K�8gc���f7����VɎˋ(�C��εrCub���G���:ngJ7�ϐO�&�N�5kk>�g��R�K��4t"�x��閯:�S�"��lf��zEf�2Z\����w9�F�u��S���q��J�\g���u�ʉ��h���.��'Cwu�ǌ;�:غ��X�xw��n�`gP�g��e×m�n����L��Ƕ�.[b�G+1t!j`�o�](�F8�9�}���}�$�6���}�h!]UR��T;�V�j�=B�.�����D�����@'�C�x��ŋ�6�(ݨ�mu�a�m��I��TE!@"���17�v��S꾢�]��/���qg��L�U��^�J�>��J��4���RUIo�:��"�V��~�	'���8�Km�����w��n]�Xk��=����p���H���F��i)��H���4�Ȩ��Z���b#_�@4��C�b���B�姻_Vm7V�A5q������U�_�bك�: =������Ը*�z�&�͓rw��9w_e����~\N�%��vvZ�p��٪�Svy��&�|\=r�;0�L'2O���,	��F%��P{��]z�����j}�;��V��<�9�q��u�`��v,��.j��}�^�i�/��}��e�Scֳ2�ٯ�=�ZO@�8U}��}���V�؁����Rm=��N.>�����+��_V�����0��\ulKg�41�������(��֞[G����k�=�f�/-�ar酊��Y�����G�| �O�VI��8ֵ���j�{�\���HȈ��H�"#RF0`��~Sۛ/*we�zn�^��]�6�9��B�p�V�UT�,�Fq���;��7����ax5,̻L�cIj�s��m���r��	�~�[X&���X��:��f�]�2����,����N�Փa���IhF垰8@z�Έ�n�@Dvr[��}�����xPlr�C�G�� �1���;�㭝лM��rh�;��d�vcO�mRޗT*�AR��X�GdԶ��3��⻉/�1���ا6Gj��NĖ,7utob�v�j"v(7��s��j�|�ovҒN�$X�����/R;�|�*��%v��hU��V34�e�+�	B�AIg�JR�ӮĨ歡��EZ�wJ�Uw���s��������B6{�^a^�A�^�U�3d�F���4�"50���sv�hQ�2�.�O��$�lT�M���i.�s�wG�����bDb(��1AV)�D�a �AT`�Fk�������x�u��]�r�f��d�^ɪ,FԪX�
b��@L6������ԇ��qv��}��w����F��Q%�������NӟW'dud�A������,��s�ʅ��.	��D�Q���%;� rL��+��D6���b����z��'�����t��q��츤L���^ï,	�乹�������T�����emK:-xd勛����Sp�˭�!�3�Xy!��H����>qun�(����<�=�Y
���nE<E�Oq�A<�W�h��eˁ�8�[�j�e�yF|M�\.�
�
qy7+�~���9N�z� d�O;���胁cY�g�j5Q���}:��-޼*���qiY�-�ykxV��R�����k}j-o* :/��\��{a[�6��A�+�C�2�Ȉ�M-&�4H�̀�gk.2:���A "�F
������$�-wW��άל���*:\E�a����bх�~��~����#���v�7��o86n7����Բ��h�h%��L�ˠ#&�,�8���Ol����Z�4����D-^R�����e�lT�������5�{*"��T�V��FA��F��S�[Hi`y��$��l�)�:�eJǊC����J��ؑs�)rU6�<>>�#�LwX�{��y�m�z��Ρ�%��>��mn�:v�9QvX���;������C��풜k���^ʏ��;]N���ҵ��U�����ԛ75�HOD��\*y�ql8�r������{b\��
#��`�e�2?Z�?(Z��ڑ�ė!�BMy���-�q�z�_pZE�g�xb��.r��`"|
x������+���:Fl[�E�flF��iJ]mS��\�z��L��O�V�8�d[JQUq���|�k�zu�[�Y�z�DV)d�,�Y���� Q�+Τ{qsr��-�+]f���:_f>$8@����N�uC;��d��:��f/-n�b�j;�J�|dxpx� �{;x;�Y��M�P�����$�B��vʿAf�y��{+�,p��Ѝ�����͕�����FJm��Q��jC��&T����SM��	�::�D+Ȭ3�R4!�W��R����2�8Z:�O!�AG8䭧���媢3���V�s{3^j�=Q$��I0�t-�.�T�+���B{�C<&��G�����m�LG�N��Oҽ�Ѫ�S�vb;��9���mL&sIYb�����a�>죜��e�걎���� I�P	 �O��� $���Ԑ�'��L�6 �(BH� 	 ��@�'�$ ���{ �	$��� I��@�	$���������$������/���������
���S�k�l�f����U���H���� @	$@�@�d�H@	@�I	#�I2	'��o���$��'��	�0I @��2	 ?�~t���� �	$όB�I' $����$I7��\� I�W�ݙ��7y0b I���I'�>����@$���$��ׅ����`�?�� IyO����nz I��L@$�_��3�e5�2@��;�� ?�s2}p$?��l�v�mb���;���w8��f��6ؙÚ�m��h� ;��e���32���uv�]��I�[��VwwB-��9���%e�6�JbU��!���k�����&Vcl��5el�[m�hTlX��SeZd3F��B��M%�Y�bԅ�֪&���f�cQ�        u�l����.�
5���:O[gwNn�Y��M*��h�    h   � @���  �@B�B��8��hw�z�G�Q���4i��Uo7��������y�����s���m{A�r���cխ��ob�̡��z�:�;v�mw]�)�����wI�M��P�Mf&�KMZ���s�{�q����5�U^÷��u���ʑ��:�7e�׵�<�����{�/k&�n�����\z�:=٪��ӻ���X�NZw�����9�
�=��e�/R���z�t��\�����l(kY�ic,ԫmks�f�W�����o9ݰ�#���k�j�:�.�XW]�݁��^/=������]vrٷ]�����N�)��a�^����+�<���N���kn�6����Wm���*�����R�l�i�V����d�v�{Ͷ�����=���ku�vh�Jƴ���]�V퍳6͗{޼���ץe�+C��]5Jw�׷�{��ݝ�[m��u�g������==�mu��ܻ��b�-�e�e��6[L�ֈ�խ��[7F��vs	Z��J����Zk�=���nʯt=�����L����M̻m��:V�.��۽�\n��f��^�4���G��Qޗ�n�[[�mS> �6�.�r[�Vf�l�M����:嵺s^y��3tn�;�o.z�۷K���{�%�J�w��[a����om��G�ͮ��O�=j��y�s�[�[Cۍ�ų�[����c���F�cG��En��ӺX��{�q�J�q�۸���]��5\]�z��Ⱥ�T]������a�!����뤀���n+ɪ�i�w=:w���w;���)��N�M�u�l���e��u�v��3-���Z�m���3WH���wS���n��kZ�u�7w:�gq���*&��u�UT{��W�^�ֺ	��9��2Ύp��ۂ�on]ƛ�9���ޛ��4�6�EU{X��ڤZ��Z�,�ku�G���v�\�ZF�����Ɨ����gI�������{��]�l���mz�p���3{��*����U�Sާ.ۯ9�z�ӻ;w�l[fkPi�e�Y6թi^3��tu�{z��^�w�����V�U��g^��v��o=�nU���<��k:r��On�۫��̖����ݽ{����rWO=3��we���[j�.�ٶM���	�3MZ����2��&ōm�Zp�{&���Pd21���1$�Jz�24 jm4��#@24 ����JT��d ��h�z��i� Ѡ�HR�B=C�<��'����/��~2?�{.��\\\��9!EU)�u��ĺ���D��$��^����v�.~�Є�	'$� HHXBB��a	O�H@� BC��,� ���$Y��*�DTTbȌO����H*Ȱ`,��H.���w��R,�YX��_�yja�W,�u���� *�s��jlL��!��@�%HQ�V�9uq]�ܘ�2���=���$DQUV"���QU�@FM��:�����l��r���l7�&�چ�޼�{���e��k�C.ꍻ���y[^�C4:Y�h�eU�6�8B�$�
�m±5	��=�PW��n(BJ^�K��f�����7���c���A`(�bŋ���k�z��fP+ ��b�ETb�s3�~����]�i��E�:��z��6��d:�,6�d�ECv���׀u�%�{��꣍������aZ̧je�(��̺�+vٝ:y��l����s�9�Hm�y�;����K!���m9�V�gJZm�2R�/U�Icn<�V�,��ph�FVe��F�{R�ZN��h1b��0�����!��X�eE<�G�(�l�NYESm}l�E�,��QTb�PU׷����k��dǮ~�EB��M�$P[D�1�s{Y[e�4��:�WYd	�ׇ�A���]-
aU���47�(��|}�f9�I$�"1T��c:8_*[A���;X�o�T��-�1%�e�
+Fke,�U~��V`��N�u�IQj�u��+%b6�j����{���7���P��t���V:�8��S��Y�uzҰº;����W�U!wPizZZƲe5��w0�6�P��EJw��4�qm�b���DH������}u�ޞs��2Bha)�(��y�]�f��Gi
�*��?UT`1��&��m��2P���!�z�wvX�[��&i�4 �UW�UEJ�X���44�.�UY������w�W��(
��,yۋv��6k �'��²h֔�f�0k��Ζ�ᱫ������o[�0�ә�߽��m�U`,X�V�EDX�((
��UU���u����w�YI52�/
q��n�Ke�(���¬�K3Q��Q�yoY�Q,ñ�z,A�mʗ�N
br�7O#%���hm�����r�ӕ���Z����w�s=��]溻���HC��,�Aa ��Pb�AV
ER)`(1TT����DĊAb���0UI`��X,PQb(�� �����UDD��QH�#1Tb�b`�QPYE��ATQX�#�XU]Ը��kU흙"�ȹ��vX7��5Ԥ��M��/R'^��PT�&������"N�����r֛��a������!E�^c��T�@�y����)���j�)�/%��]�t�8�T��#�r���N��[�^L�6�~�c�SJ{l�(0:�\Ux%�@B�*�Ò��d�k-ݶ�V�BF�a�t�ظ�f]`�f,ʚ���PIr�2�R�j��yGpb.�MN����d#�æ�̈�Q:u���6�m�<����%�E7m��X.�*mCq]Em���w0�rD5;����dn�Ī i�ak��Z�u��7IqB�Zq~j軕�#����{�bӴ+M�:4+sE�c*b�:h=�<6cǩ�h=��L[^UV�i�|�ʆm�����)�5��K���#u��
�1�oh$��7koX�)�ǔ��L�am-:CqZ-��n�wv�a�B�
�4���v�8e'Z�n+��6jv�+D�8!b���&tS,j��3y1��d�E"����B�ה	�dY�bEB���b���u��Ӑ��;�!R�VF�TI,:��$ʽ-��ӈ~:ʷn����]�ۑ-��@������x݄7�&��xh�,��\Q+W{e���qn��V�/l���U@a�$2�����v%��_�
��V�bi�l9.��K�hHq �E�䢈��)�E"�M6(u��6):��V,�E�q��ڑx���W-�R��T�j�ۣj�\N���4�n�B &Y��$e����2N�[v��P憓�l ����%�M��T*��'^�^��h�r�n����d�Y��晌ݷ�sV����S%h�4���@���[N=4�^��\Tn� 5m�ԋ�h�&��S"�rKd��Cd�lCQf�����6��-�AT��J�RT�;�v��A��*I4� ����f��p��[a�� e,I� ��2��Q;��p�ÓYC�a�ܻ(ay�L�.T������Y'L����x����qa�ɣ��\2k
fM�{U��-�Cs8͜�[/u�mۑl�A�Ǫ#��[�5��a�-�[�{�j4ot��Q��
�ٹ�1�O!ݼ55��ضD��&�ʭP��w\Z.���i�̱YL�xB�ʰ���j���U`ax�2�/҃��H��Ip]���ʻDV��z1�dk;�:L�B��}���]{�Ma�y& 0�Z�]^���?+-A"�fшL��
�5���.�63s�p��x���|o�}����\ٜBu��m'����Op��g����o��[b��f���yZ�#j��7ͽ9�����mT*I���ԱU�Aam"���
aQv���C�P���ɻ*�-�UQ���Ij��@�Ie��W�
̧�a	�i�pY[$W�Y��h�6�X娃���^�v��+���Q��F&�8�1�VCb��Ӎ���K6�i����I�B���M$�PKrd�y���9���}��Wk��YA�Z3X��@*������|���������E{��q*1�X����,�ci�b-IY�UCڸ�Ym2���$4������X��U�ZUb$<��HT�`i&�ԇ���C��1!��N�Hm��Hu��
��d��]��u�[����'��8$4��<)�,DF*���#<�Tb��ԔM�E��Z����<B�R����(���(�:��Hy�N��y�c��f[Ԃ�T�J�8��d`������x������vK�*�N��H�����5Tm�:շ�!���A�v�M�n�{��y�7׮�gV(�@T���U* �4μ���ZӍ�jZ�Nm���Y���5gU�XÈ����T,����ó(hq�VHbu��V��zj;*���R�5���,K��ޣ-A���R�y18��t�Ć3���k\4e��,a�@�ʖ��b�v�g�x��ڸ%Wbe�U�Y2���P�#j4eɺ�T�����R��Sv�H"ñi����j�B4`�B��ڰ=�C]h(q*�Q,X�[S�3�P_{^�g��i�뎷�x�rj7�������/���Ʈ�j��7OF�󪗙�C#U�-�%�m][�ԝ�*m��r;��
���
�c��,9jdaX�S	6^Ku�����;�zs`����E���Ʒ�v�S8�!�Rj�B^��[�z\ǚֽ�w�^���e�l턚@ҁ_�]4<eH�g���Pj��wiirħ���"�n6�<T���<�{�qV�2�ef��] ��-Pء�e=oK��>�v��h��(�zq�4սo^]Ksu���Pꪍ <0�PH)TJ�[.JY�p�-��*��-c���j��h�G<(7t8�e�HU��mP �ȼ�e�n2�ԭ�:�<����$y�����Kt<�.�+%��H�]���vc�ak(]:1�Z��J�0ɥ.��g�ڴF����Á����L�njX���-GU��^a5�9��[f]��0�v$�����d�:�h5L�ő�d͆�
�;��l��4�����bJ� �5��0a���a�2��k\XY�^�+*���W00`H�A!��+%�r��б�4e�"J�u` ,�ޣݰ�؄G��7̽�܄бUU�	Q@X1R
*1b�E"񒨊���DTT��""��G7�o6縻�臭��`�,U^e��ǁF��(c���Kg��0#��A����Q�P��T�u�n��:J�,#���ض�*&�t�6ZۏwY�fi���Fn(�l +AE@�9o�]��SѷT��)�X�mL/P&d�h��i��n�j��u%.����r��6ŭ���&wj��Y�ƮmY�2M2�B��M�����[��-A�FZ���z%��q����Tr��T��!��=��*�J����v�q+L` �tJ����N��^�6��T(�L�Jmb�^K�"�c`p܎S.U��%;��c����P��ƪ5MѿMA6�1XƳ��%��Tʙ*ջ-���-�E�EyN� �Wz��Le,�X�;l0�؀U�m�T��8�x'xww�bn�R$��٘2d����d�<(�"z�U2�FV���Nzs�;^�*�Y�ֽ��l�4�:!��2��z�8�:�� 8����T�-��0��M��仂�AZӥ֖w���I`@b16�2�mf��4���Af��D�o)
�Ч�f9��p�~�\�ݪw����=k��$�h��3A�U�m�Z$�հ�JZ� �F����n�MS��U
�T�c�������(�=6fU��d��I��h^!Bf���
j�Ҏ84m�I������6� �Lu�X6M�SN	��g�ۘ�6��kp�*{>��a�&��^��oZ�a�0���q93�:��-���n-�H&l�%f�F�9���{{��W�V�C�Z.�ee57GB�4�$͖�e��d�������bnU�N�jl��pm�~U{Z����T�U�����ծ[N9&]cn��-���D�xIIͫ
��2��v��T�Ĳ���R�oZz�0\x�
:�F�4.�u�����F�D���)̤̄�sj~NSǭ�fdh��4\ņ2Qb̋b^�4gUf�T�]z��Z9
�R����-Vj"����ݩtG��
EP�}��8o���f�s��vۍ��[���iPnU�+f�=kie�����)`�j14��l��X�����"�z+U&`�)K5�s����;��eQ��F�M;�D� !(�WI�D��a?��u��`�e=	ǆj�8[*��x򛳒�5^v��b�5NXE�����A��YJA��Q̪�o����:}b�/4 S��N��li)V�*���fX�.X��EPc0U2"gJx\��GzF/2��ZV��5Qw1����K]�nнw���˷MS.�I�SHZ���F:8���������̠ӧ3�V��,����ڻa�3['q��l�Z��zQܫ�H��*�%�V�
7 ���p�A�`�7-c�U���Z��NlK7BX��B�6��y���܁���-Qe�$���@�fҬݬ���n1�It�5�b�Qo0���*���{��}NҺ�je�ѧ�އ����B�1���Qb�PX���������ﻭ��y�P̇XHu����aR��$�+	&�ZC�y:��uVʼJ�q6��EP�œM�f��*�㱯p;�@+6ަܦ��v4)��\�XVo��*���� #��Ś9݉k�(�=�q�b�o��}/B_sM���7�.����\Lǘ�$#��@�x��N�������"ڽ�a]�{6�b$4�p;J\�`����:Z�q�+�iXh_t������xv�s�#6��c�6(u�Z�X�{�Gz�8_Q�zW^�Ve`3��ǆ��"7���e��e:�*m�|��ӬD�
�P�X�XڰO�����x%;�8$r�R.g:#�;������G"�"��5�EۆPZ��<x��q�kM�}c�v���#��Z��c9v�#+�9�:H�3&�=w]D�ws��7m7���K5��yN�f)�){j��pQ����M�q���1���/)6I6f�a�ƽ�:k9IS��^,�������q�E�h�Fs�wٔNuXf@�]�2�t�3��8!x�����؃�V��Ş����uk�
�Q��.���v� ���q}�Ww��A�".K��e�X���"λ}X�N��f32�Y+j-���+̽�ݒ��ؖjn&p[�zp���9}���jZ���ǍȘ���eðᬖ�\v�;�8��{��Ht�S�5UB��!�f���0%�a�4�7�W\6�)R��z��[�r�5��j����ů�r�o_n>řʳy�x���`�ݒs�`���Yj��YY'N���H���ʵA������#5���uL8�ZP��������N�M���u�;,>���c�0pT�w[����/�����z��P�o�ރ�U��9"��:Y�9j֡%��<3M����اXC�:¦��ه�� ��ri�RN.�W���:��A��iy�����4��,����y����s�(�=�]���#����G�<[5��̇��u7e��Yb5a�w�g���L�ɼpݾ����*�,Ё�I�'\̼=�N
jȬ��-�G���h�1�gi������fs+�mh�X�K���j�tˍ��d���uu�
�x��v���h�g�����j>œ�1*�B�G�ъ>���8)ٗ�m�"�;�b�/�#�a���K�;WZ�S �sN6a�XţN�A7���_�I��.d�uҰO�G]rY��MN���q�)@�W�z��!�Rf�;\j�F���ò�'�h�$�x3��א̚We-�t�lymN|{�`��2��s�j{ �8]�G�0��/��q��{�P�X<�;$_����U�l���V�*N=�%pͭ�"j	F���5��R� [D�2P=u�pZƮU�2'�
�xf��G�mH�� �e�pV�G. �iޣ%��3"�p���}B��˲�e��M4cI��ہP��r��l��y���Saªv*e�ڠ�?��0�爂B��������
�ga����W�Zb��(H�r���g��]�nP�e�IZ֕��l���,�[ҶP��]��qv^�Y���� �N�tgE@Z�&���V�2�vYJ[����K�]�<6�d�+����ƥ7���V�0�s�jƲ8^�{.��I�)o��g2;��nY�����f@.��;5^G�A����i���i�.�r��YJF�7�8�y���nvۖ)�i�X�<ѐ< #�4f�ZdUV�:iHR��Ʈh1$	�al���B}"�X����C���S�YNR����}�Ě�1f,�/i�Av;t��r���]^���ivs�&ǎ��rۥUޥ�w[�ؙ��K1���Z�:���:	����)k�vOK���Q�S1�Jp�K��V��Y؛BA������}uY\���OӌV�J`�Q�@�+������S2fs4�fؔd�;[}d=H�C�Z�\�4d�rm�C��O�P��=��G/�h���XMe���v�e��PZ�D����a�w('��W������c�м��hi���vk��j����ZlQ#H������ݙ�xۻ�*(��KVn�,gb�\wI�����׶1�sb����=�/�����	�,����1�Uj��u�DP���B�ٔ��&�
J�Y�ԏ���h�U��<]X�/{#aI2nˈ�,U�v֦>BZ�c)��� ��������T'iT���`k{'3X7`</(,x9����N�т��TU��3Ƶ���V�5ߊ커T���cmqg@�{�1;�\%��m��.B��=��/Ln��mĭLV��Y��ЂDq��yҮ��ś�ϑ��{��F���B����-b�2a�w�H�7�F�B�u��X[� y�2��H� �i��{r;I�P���E�z�
�����]�ǝ�'*�_h�.���f6���.�j�@�8�W@u�V�v4L��T��jE�6e�u��}��[��[\��u��i�(��=�i����*����'�a���u�!�vV.���:���
�	d�Z0�8�qƴ��O9��*AR�e!@sA�i�����x-�\�ll���ν#w�V=�ϩ�U5m��Zǹ�S����a��|�	c�� i��;�e,�\Iwhu>�On�,cq��Q ���\5#�n����07q45��U��֞|VY�VMȱ���m7}/p5]\�e���R����a%t�;�ι�]2�+`��po�w>Lb�}W)]9Z����0�.��W{*���3�	$�Ժcӷ5]Rgd�t�H8~�
4��ŜI);�]
��md�B�Ľ���F<�8��N�V�;�e8Ԯ/�c�a)·S�G=����+s����W��\��P0C4:��&�3���j:��e`�������P�K�!����zo�F�@�S�75Q���}�cǫ�"����@���6y������?3rt����Aڐ�E�s���0f��B�A�q�SD'-�ʲ�c8�2��zy]�j�ml�!���r���Ȯ�K7gGowi�[%+���w��X�Rq����JB�B����YI ��#,�{
�LrM�*>�D��~:P]�޹n��A����Wۇμ{���ɧVC�p9˚k_�Ѣ�%��f[P�-%mj�Kr�2��.���Yۊ���
�+(�)8�q���kw��:��AV�^>lُ�_A��INQ���̶�T�U����0i��J��r
B���X
c���7�OÉ���T�47�ڕ��v-g�mUt��F�6��EeTPwl/�~��	�Zi�.]\����܊f���}aX���nY�r[?��m�M��x���
S}4]���+F�rT�*,g �D�R�W] �`��mh^�eα�z�خ�E�x9���*�'Uf#�	�j� �L���Z�o�{VRĒ��=�~���͊�gn'|����F�����F�Z����;9pZ^Gov��F��nma�o4(�)Y�9�r�lk��q�WF��[x�&��쓖=n�Uq��U���sj�:�z����2�=s���/r�n(�]�z��m%�s.�	�Gc����0H�8,7������k�Y�zs�4�V�R���Z:SG#gdH�ۓ*��5&�bk'h¥�-����{�M��F���F����e��l�c��5�k5;'7���;؛,�����z:]�9ù֚4�+�_�r	R��#o-��V����B]�x�l3O3|C�b���I��3��CqT#f�\��nLe�)����E�y�&�!ғ�C�t{v���X�9S�ܷ}�\a=���yh]HM	��j���ƥv7��=���
wO�N�S���&"�׎���5%���ǎ��NW�;�_>ܭ������X�U s+p6��:�޵ϖQv{]���i<�	}P3m�)���Üz�P�^H��q���67��x1ei�	T�B �}�SY�қ���J�SI79c�;3�����ͥ4��35"�2�,}dݩJ䎜��*�9�JA�ke����R�oh��)�=���!ȇE +�
X�M.Oɷw��m8T��lဩ�G�v��DVmյn�Zt<.y-ii���Ŕz��|��z�B��äL��I�%��L�Se��j]ͮ���Ѝ�U ��������\	ђ�Ψ���:����E�=X�ʾ�+��4��θV=�1��Ӝ&2�� 1�t�;G89eu�֘�Ⳍ��L��}JÃV�NeJ63��݅��Wu�-E	���ЎG�q�E��D��¾UV��1�õ�@�٦���+p�OI�!��5:�bu9\YwY��w���rը�ax�+�er��w�2�(�]�@`��ڑ�"�#�\����r,�f�����ۥ�%����it;Z;h�&C���f����)�5-��TtsQ\���"�vb��󻰒�Ӓ�>��&���3<j����E߲Jy۵���?ovG�b욨��լ�κ���$&R��|��9�}�m���L\k�R�+�d�Ҧ��=�'3qh�ouq�Y�ԧ��jn�PFwGb��$��W�4��hB��C�|����P��TB�_T�4�w#�;�k]�/�F%nGf����{���a�Χmי�n���6W���<wCjf��P�j�T��˦��Ŷ#�hr�i������Y##C��S��@�U��shWd��޹�v@Z�#�y��"5�]��r�7U6:�/5��dl���n���Wi�S�鴨o2��#���V�A�&�*�c�����:���T���k�Z���^`��kw�+F�˦ۈ.S���{Q���݄��A�E�1��`P5�1�vS��)��
b�[1�7�_*N%8Hs�C0Z[X�S*��Z*qv�C�w;��W;������lؔ3˄Ɔ��3�e擼:�p���%����#
*N���NZ֛�Q���yp�[�ZGu���6�U3��+O�tSݷ�1��%a<{�
�I�С3-��_��{�9����t"�8�jg�����{ۥ?)1�Y�h�w`���h���X}��iǐa�1b��]���v+��E'Jۨ��ӽ�鎅��%4CO�Ԡ��d�a�o� ���t;�ꙣ-*�gvBc��5E��@��k�nݹ�gv{�����ӯ\e�|���A��X7&����h���qв��{�����v���6�2N�� ]�5�wו%�x���(�n�6��v.���2�V�9�7��Xv��q
���+�"�+�sζp�W��K��JZ�ɺ�7f_>�ݦ�M��k����X�困��[ ��fj���%)���D�"��*��t�V���($�g"k6�(�5I7;�A�MZ�Rj�S�Y��Nl���ۃ0Ы�COU�O���Vp}cZ6[R�R�j�i^L�o]���l9)�'$�`ES�x��{Lf%�\����0K8Si]�� 7-�1Qm���'e �Irw�sYw�g2�9��S.fY�9��C��:�x�U�7jo���b�u6n�g��)f+�M�c91�v�.��y�ƨ9zGa^+tɚ ��Hh�Z�ͺ�"}ưܴ{�1C�w+f
e�(;��md�d����!{�Ώ�0k3)�����<}II3��<}ɋ�[���璯
yk������/C����f���p�ne�`��Έ͸�J�I�+�b뾚:9t;*h�'ʈ�f��t�K-l5��5UN���}�^�:ߓ9�6t�[��Y����{�%
�:I��q�}C��cǆ�ryu(lF=�Y�|)��J�˘(`�HЪ�:܋0�o�yի�,��Gz�4*�|$��9�S���KA{\���nd������3��M�����)���! ����`��|�jb�S2��Lg3��9SwU�؁���2X�H�P��{�����N�鐥��G���9��L-a2]��T����Υ+��ξҙ�j�&�H��b�y�-w���ß4�,� W�Ki� T�Y�c�pf��${����e+����euS�3E�QB^��BZ?���'����r���cƃ�Ǜ��W$���7Y��Ѩ��Mg~��`#Z��pᇬnKλ��
a^Н�A�ILzm�sl
�(B�g�i{�n&������wvU��,��e2�	-p;1֊KP��+{ya8j��"�o-Pң�X��OB�k�p^;TW�����ͽ�&\T%�]B���˳}?f������9������u�KV>]Ϸ��Y�Y�NdwU9�]��S�?���wl�6�u+��i�,�b&r.����� �T��E��{+'Iw�]����q"�%XAu�Y�<g��<�t(�l��ĺ���m�q>�N��t�(,.e:]��7wu�&+�<f��0��U��(҄����R�Om�������q��O	�d��J�w@Q���2�����m�u�J\���N�7Z����r���r��"����!Zi�Ek����;�))xFn��r�9}Ǯ$;هW=�,�~�G�UZ��{�p���2�]��+:]wM����lЛ3�)s��v���\:b�&���3�ɖ��}J�8|zqS�_u߻�Ӕ��v�Mҫ���珖,�@	U���� &�M�MwXh���ƺr��W)�ۥe����WX�B� a��N��F�T��N��[V]��b/R����n^P��p�=�=�q
�&k��:h�|����R��5r�%;ݖ�!r�^�����B5u]��WDs>����H�\�k�nv0���ʝ�$0^B�f:[Ӌʘ���&�c��]���ok
��I�����&�,�Y��VO��]ni�vI��a�D�l������t��s���r�x�DDj��)A{�\�^D3i�%j�D�gu*�;,�vu�緷����<� @$$?�B��i	$8�H��	XB�!$�$�'�vB(H�@���@��C@�` Q! c$&0�P	��$'r��� �Hi���i o�HHJII/ZC̐�-$��B@/�!Y$>d��C���D��Y	����CI'ڰ���$�c������	�!�K$�T |��@�I��@9�Bi �?Y
2"Ȳ�(JG��C�	�"�i�`u �s�� >�^R���AdXN$�urH�����wd�E�A$:�y�Cܰ8�^X{)a�	���'Hi#� Tr�c"�G����;�I�`���hb���ɘX,��Z�0�!:�yL�0� V=�6�ꆑ`"E�a�RE�CI��'�Br���4¤�7@�>hM�̡�fM�
��kb��t�M�j�vɉ
�� �Q�d��&Ђ�D��eE��T�Ww�ͥ*,rȢ�4�]�gR
N��R��|�'ڻb"��,�"�d�I*:�*,�����1�I����ư4�۳L��5���eB)Cljɦu�YT��o2^��P��6�M�(E�aR<�LoU%v!P��
�R2fYj�u�&Щ:ϓ��R�@<�n�o�f���e�*���� b|�5�<�èq#�il�ÓT>Mj��m�jM1՛ޗ	.Y�5H[eb�jDv�0Aa��I�����<ɦs�$�w��*#>�=�:�٨�8�H(,�'���1Evq!�U�O��s�,���h�����&٭��Nl��3)X{�Y�S��!��.XVs���CL�
mx�fh�p`�j-�� t�2�ᔚ�/ib(ʹ�ɶm�����+ ����L.��/xg�i<��ʇKe����vM�}��)R���^ٴ41(T<� �Z
w�l��0�켳���f:���Q��*V~�ѯh����`q����@���ui��bE��3Ԩ��_��� ,�����9���u�W�9��ݤKH';M<ek�d��2�;�3yw��A��dc���ML�4j,4�X��T���|�j�IG01����3L��Y1�b�3�I��n(��P�q8�wnj����~N}κZ�e�X�\�u/=f,�]w&��]���F��|��3L��n�Co�۔~{�ӭi/4wv/�{%�oGP��Y���T���ۦs��A�Q�`wE��h<j��a�^s3,ۙLs�{���[��4:y��|�sG[�:ݽÜ�B�ov�mУ���ATM�9����O�J�\��iﹾ�Y�
�o�Tf��d��ɽF���t�z�*����SGy���r�滚TQO����
��*�
�����P��S�uzk}7٥N���=e5�h��%��z�Ӥԣ��`n���u��SǞM{��S��eˎ��/R��0���ZGH7y�Q;��Gܳ7o�5J�'u�tu*�r6*�u����+E����Y
�i�Ɛň�a֡�G�tS��3x}�zJ�"��
���uzR,����/mm���S�Y��oE�~un*m�����^�hM�4;O��hy��5G��p�#a����q���MX*��$m�5#���
 gccqXc�ELT�0U-Y�$����[�QLe5M>�ܥw�X�+4`�i��V�5��`,�U;���mr
1e��e�p�i��X�"qd��]��%�q�g5E.9���`�
��r�b���kV�ѡ���h���	rT�P�`�T�X#o2�d�cVD�2�Q���\oyDD� ~�� SV	4�Q����\o�k�f�j��F�ձ��Z�)-��*��ഺ%_���F]�n�(n�fܞ�=u�aE��+S�oY��y@�yK�Nd
�Q��|�����S�qt@V�W&)���kg��4���a�ۧ|hY�8h ٭_�}��`d�Ȩj�T �)sFL���£-n*,бj�o��pkX������P��gmH�PJ)�4��:�^�h���l�W�J�m�)�!�4�fX54�T�\)n��2�y�^ڽW)P4՚B�$� J<F��>MvB�0�ڃW��Cͪ��R+u5�m�+(�}ǃ��7��:�1akxkF��<lm��5A�i��D�]�yQ�_��,�r�u�h~�l�2��_�����Rl�����8��ꅤ����66X�G��Wb��X�+�) �
v��G!������ҥd*�6*���{ESƘ,��\c_}J��㩢?h���"5QF����ֿX�-E��ӊ����U��
�gD`!�?c�s�������G�e+Ν2%�p�N�.�E�߸1W	�_�R\駦�P�+���WW�PĀz�8J��:�U�%]�ub��8��\�-%R�F�"�+4ۢ&Qn7x`G�*6��`�3�T�*P�Qeۢ]3��W!�]mY��!
೐湛x�٪,�� \(����L"2tdU��N��*U�I�eV�f���0*�!�
����a��f��t�Vy��4�����v p+��u��̧�/^(�KB��6Q�/_�GW�u=����D��kT�Q�ت��0��M��������r��I0�ƥ�`VNC��%^i\#�V~hJ��bA9&޺�4�O%@�P�F$`�0��t3�T��2�!m�����W�K0�(�
�l�������b��,&s[�gt�*�

9�ƣ���uV�
b�5���u+ڌ*�&���Ь�}T�
�d*4*`wM�pTlTjJz,��$M���BD a�I
�d]�����a7�C 1�)���Y:Z:���i�x��۬7��
qL.~� ���GFb��,X�/iPj��xF��0�
���2���������q�? � ��c�or���gI�]�Y���.��)�̀j�fS�m��hP�WQ��u��ubبͻ�,AQ^�I�؎��^��W�@Fҕ:]���̂6l�n]�+�����fa4}~���wh�d��T�h�e�f��N�;�&|��eQ5-��WZ�eVD3��S��wϕ�=6n���(��e�Q�9���E��[ �n�,�i�;��jA�Q�R�9�t��f�� E lB*	�hJj��5�tD�顸�1^��fU"XGl��TԿU��쐬���up�\��i�3�;4�uӾe蕦/њZ�@�
Ȏ��B�N(���ӥc,�\�w��$�E�Yf��B��a���)Ҕ����aͷ�Mm�SJJ��T#U��y�ȧj����Y[��ͽ/ȇ�b��f�x��v�"�&�nV�Qך��؞�w#���`%;��M��&
�͇�����	'�����َc�W��pr�����N��8�37l�@�Z�=N:ĩ�F󁹐��m��Z�g�KYؔ����!�֛{)s}��;6���}��tŎCQ�WU�
X7}rv�I)
�}oh�ת��lgP���l��3��4N�F�N�o3B|?�ɹKrMDN7ݓ��s1��;)�{��yT��bf^��� ��UGć2��Ջ1 fm:��X1��|�R7(���Q!��~h�λ�8Q��C.c}�*�	p��݁�T���u�=���f�?	����Y��bkN�o��.��&1ͩg%.
�n����(���w���\�s��ϧL��]ɺ���G6��$����x����zm��M�X�[�/w���!y:��%�Z�%v����Q���s1�>�G,Q*�P^�����7�M�W��-�wL\WN����ca�w�xtt;zY��]�(��[B��7��J��|�v�24i]�·�)�ˑb��ҫ v�0�^q��c.I��7f��Ǥj�S�j�3��^Ց]@P������ؤsRZ�yP�J�����(ۙW�&�4�*��C�U�˓�|-)�^�,\�����
%^Ѷ��v-��ڽ�l$b�ɧf;��NҒܬӔ��V$��'fr�y����+X*���w.��^�Q�T�>ItM���w�3pz�+qlB�����������5�ߜ��К�sF�St�ͼ:����}Lv����B]�v��`yr�Z���`f�-U��{�7Y��Ӻ�Lȳ��}�a���3�>�3���H�!!�����0柴j@�@�4� �Hy��� c!$>Bm�,$�@�iy!	�����)�Bk�։6�8�Cl� 9�g�b�Mw̷z�6_�� T ���,�*�X��DE�DUX���UH�*��Ă�%TR*�Q��m�-�b�AEQUTb
�@D�QQcX#"��\EUTX��"�*�����DA
/�*���+�Ŋ���bO����8 ��E`�1X��U
,��Vy�eTX<K ��uq�U��X���Db�*�H�U�UV6�V
QY=��&��*��*0U�(��E�@U����
�
o�Ȋ,X�X
�����Z���PU����1QAV"\֦�T��(���"E��X�U?ZȬY"��FER"�=LVE7J�UgRX#"ş�UD,�
��Q�QH��F��db$�Ub2*�ŋb���<J�

�����X��3[�"��?,Hx*TiTQUH*�(����Ȋ��,U(���P]%D������,QAdX��dX���?�""��-WY�#TE��(�g�R�$b�
*DSϾ`�A�*��
����F,�b��Ub��PQ�U�*���X�j(��1X�E"*����TV*1`�(���
���@R(���Q�Z�X����1~�X��UQX�� �(1����bO�*��L*#��mbgn	r��EUV(�*�EDb��7�Nꂢ �#cRɤ*�j� (¨@P��
m�����]����s����_��s���
,TH�Ȳ",PUxغJ����AH�U����X��b� �~i���`�@PU�"����eb��UY�kKҊ"�T?Z�X��X*�Y:�!�sZX��EQ�+b���bȨ�{�kPTG�U�
*Q�PDݢ�W̬R}�kJ�"�Yb��b�t�X���d�(,UQ��*��b�S;lTX+��**�*"��R�DV*�(#}��V��X�
,uh�O�[h�As\:�5�{U����?~Ϗ��s��ڌX�S����E��weE:ְ�((��T�(��G{��c�<�"$�*�Q`�Ub�y����EeTX
&]e*ɛ�k�,�"������R�X�gmH���*,EA387X�1��AW�EUF
�kSB��~�(1EdDQa�ـ�(1UZ.�؋(1�jz�U>J� �^�U^Y��`w2g`���gèYQ���Q@]�<���X;�;B��iV*��
���+ƈ*,C�H)�b�����c���lF*n�~j#�Tb��iT|�n�cL���E�;�0A��*'iA�wSJ��(�UPED�Q��C猊�j�M��,QUO��xU��UUa��}��g�p�?o��w�k�=��UweX�-�V(���[|63�Y�X�����h�UElTV?���`&�ADT_��1�,k���8}�z��QE4��9����(�PM�����;��ň~�Q�������Qժ*��#� �W�y%z�þ=4������Q�ҥ5j�QE}��ٿ5wJ���T=�cAQ�K��EE1F)�����.�*�"�x�K(��
���q]�f�{s����GZ���h6+�1"3{3�QEE���bԦ�\X��3Y����7��ގNK�3߿�@P����0�����)mPC����F��4�EV"*p���TNk&{�z1S��)X��L}��J�"�I����]&"����y*��PY�LJ*�����c�QDb���HQFk��ۮ;5w}��1[���p����(P��\�`��u�2#�QE~J�UW�*�[U�~օ2�*�O~Ɋ�D�f��m3a�Pa��y�c��(�S�o��lU1��a�AG�b��`�������k&/�P?]�6f�gW'���#�����y�;fz�[w�Fє-p�]��n�$�ӡ��lA���b�Զ���G�+���?0_]�i�H�Y���{��c4ol�\X�5Ng���;�gL +8g<ڵ�U��`��ݽ$��)���˔����{ZZ��T�X�ܸ�QER!抪��UQݩ���lЭaE�aX;���UQJ�S�ԟ���?5=l�Y�EQ?4u~��ڪ�l����F3
U�e���1���#��~�[�|cy�����ۺ&���E��6��'}��*
#iC�*#Z����(����z3e����Q(��s���1�����
���0��,E9���QEcy�0N5}�kB���?S�1.s��.��/?~���s��{n�!֢����=�LU9i�جf��a~La�ꕂ��l�V�Z�1����ł"�늎�T?'|�u,X*#��R���P�fUU�{�1����5{��? q�cY�r�?�wBz�� ���|�G��?���
@
�U�j��i4�[�Y>vu*�:ߐ����A@G\l��H,{eS_���J�E<����L��Ϳo�����6_�Q5�osb�F,
u�
��$P�
K�F���:��Hm�o�>? ((�D��}�7=f�^~����wCRi&��9js���ڪ�W�+ǻ��0�g��w��ܨ�S汞��'P�T�����7�Fi���U_52�ם�����U��\}��}�7������V
��WID����zџ}L����=��p�(�=w��k�}:�m"/䔵���*�m>/=�?!�Ub��w��y��>f"'��V�_�n�x��;+���b�d!�5��,A�J���Mu���)��?~�B�v�;UI�S3[Ԇ�}�&!�6#�S�Qm��������T�b~�3�ZӉmE��Pt�)�G�`�v=S��s*���b ґ]�ϭ��+�AD���v���Ek�㸣�+��m�~J���u�s�LB�
������C�]5���o���Ӗ��֚�����>?  �?@� 上�;*�J�����]�d���~�XcB�21FҶ�U3����8&�g�X.�C����߽�q�V�g�X#��R~���f"����Ck����ڪX*�_�����4�� 硿R۬{ϧ廸17h����͋:݉CMb#��������Ԕ�Q���L�D~CI����^�kF��!B�I���/̯SlY�߰0�����C�
�Y���=���F����(�=Z�`����߽����b�ĪbѺ��W�n�_d�.�&�d��媗+����t7062q�urC�y��@�Q��X�M�3���۹�s�2[V�	P�o���Gm��PC��G8�:��Jގ<���A�K��@F_�ɴOXUAkT�3f���6�S��z*?S�Y��srm���������C�{�g�Y��1�~?d���DX��J���>�<���ڮZ*0S���k!�i�U��Kh�ߩ��o?oڛa�Դ��0�٣֚������Y>���+bq����|�o։ƨ�Y���f���0�N��M0gV�]��\W���{���`DPk��*4Ϯ5�1����}��hY�?oW��(T��j���a�Z�婿}�f'��K��^����"ۡ�zm��.���|�s��J���ؾ�b�5�u�+2��d*V}�}����֡Կ�f3Ԡ���7��ޞ���[Dg����nZ��.1�㷨q��Թ��=�8�����Tx}�>d�󙭪("���i���>��֟2��o^<���DLk#7����Ļ�U����W)M5ya~iD�~n��}C@  ��c�s�궈���%c�/��wh�{�~���M���+��֐���N?= 4~Q�^�[ �A�5��_+�ss��������Y3=�0���XQ���]gw������]���.~����X���n~�/�T�=��}W�X�NOܸ����~�0c�,>���uau�&���si�k4�K?7���v�/�ϙUtn
��WE>�ur��p��R�%`�_��������������ݫ�ލ �j�f+�y�{GSA�ʬկ5��|��ǩ��S�nXS]�7?!���Li?]m�;|xgR�� 
�C/�ƫ����j�4�\繭�ٴ�k�~���\f9.�*�'{j�q��*���EUUG:g��Ȫ��G��5��/���b�G�N��w4�gp���+�i��S֪�9��'{_kQG�{�<�d+�?e4s�&�T�~�c�*~J}���W�vVP�4Э��b��ͩ������t���a_��x��!�����`�'�f��t����:��������R�ˮ^�Fl ><L]B+��m4�H�3{V���zѶ�*'1��"ׅguC\	p�����O+�8�Y/{���B@Sغ�l�����V���H�?w�lL�aQc#Z,�gsz�?8��?~�;a]RǗ�k��8�G�������R��r�Nŧʂ$z�^-B�P��A��k�׃A��7�r��#5��i��Q]��#�f&�~���i?yTD���{K;�f��q���S4q0Y �S L}��ú�Dc�]��z�w��G����!X�%������S��i(���CUY���?}|�Z(�Z�3z/&����4$X�����Z&YkEXu�߿w�}�v�8wW���F�Z�P���t�Ю�0��ޡ�f�"��hvX���Vl�~�b��k[׹���;N}��{MR�͗�ͳb�Ǻ޴q*q5��"x�7�3]����.g�[�X_����~�׿a�o��0��
��~��iA��}����%.𘜿+��ވiys>������=�	���ަ��������u�d�>|/�����Fg�ɽ�����Ͽp�����"�ڡ����w�o��~�ti.��uc�b	���u��u�៙��z����Ț���aLW.t�yl��Ǧ��q�<��]o�5�?b�}��k����3Hq&���n"���?!��v�uT��3T��F�q��R��l�͊����`�X���}T%����IYbwyPt~�~�w�����S�i\���Li��O_�H_�^f�NZe9���Za��)8��װ�>NN~ͳݰ�?4��"k���?L�C����*�sJ&�����o�M��+��)�P����:�g�_k����俽fy��4��k5�^��Q��[^��@��tP�g�|���T|�w����ow�Ҋe���qb��m����xݗ��B#Z>�d����>��"v���,&��RI�r���?s?��)�(� �)�Vfs"~�y�mn�ٽγ��
�Ք��+1��(I�5���[D�7sŽ��,u>�TMR�m�'y��P/qk���W@��gr�v�q̓1f�S"��D�w7�r�=�
�jJ�OCO��4[����9a��6xd5����um���ͦ�z�`D��b���"=v��������:N'��{�ܿ����tq���<h�~³VoOv�.��me�9���^��9*�p�e�X���(�
5	^�U�yAv�$c/�W�T(Z�:�#B�"�����	��Sp�c���I��Q������~N��S?~�NV�^i��ҼA�������͛��UN������~ez��
q��C1���d�����Z^�1�R%�cn�n�ӿDU���c�(�L)D�ǒ���"��@h�p�,~ 
�����*4G��[����]�T�)����T�9؆�3���<?�P��I��~��hA�̞�^��ܡ�i��C����k��~�^��=����d����7ʏ@y�J��p�쮾6�Z\^f�wO��=51��g��}�"&3Ē�_='	%J�9g���`|o\�?4��*5U��\{-�3���1�.>���
>��1}g�2�;���=z38�ˣ-X���h?]	���f~����s�6�G���o�f#Ci�����.p�Y��0���L8n�S�����^�4pU�'"'�8#���|�����*}��Ԭ���H�fuKW�VV�x�u�m]Ң]#N^P�D��lW���u����~����QS���aǂ�9�(2B7�e	D8z�+�ឪ@:Η�qe���(A�����l����h���~�ju�W]�� �s��$}
G����I}aU�5����8�U��zq�B���~�P�w�r��Bg%�V�=Z#&
��KmG���>��|>��@�!	�B|�H�$�Y	6�$�QI c$!� `!	�'~a�@��'e�]�� ,���R@7iM�`u
!� q��@��5��y	* y�M��[��%d�� Ĝ@6��I�N2 i�����M?�2I4��B�,6��������0�H|��H;��+��|�|��#��e>�
��/g��5�n��%��Mn���fB�«Z�8$��GL<������:n�(������#d#r��t�*3kݿozvw��Vhsy��t{�ڪ�jQ��<o��tI���@-"�[��#�k����]�韍�FE
�+��U���A�eQ�MPϯ˗��2����Ơ�"��@�����[#r���iyV�ڜ��i\3�#�4�E������xۓM�?a�޻?t�.�b��Ҳl�C$,�@����xJ�U|�W(�y*�o�g}0vghw��>*3P�p�T�0��un����*.��4'�}Jk|��斛�`}��H$�x�Oa^M��3UW�2�����Ґ" ���!;+���'J��~��5��Ł�6b����v���iG��#O�hׄ4�fݺ;�}�����~ԅ�M�t}�{����/�r�i������z�9g���1�o^�,Y���6�7 /�_��<+�* M�@%n��W�F��E��*�K�D��i�z���g���)G�I���6�n�!��$l
4���c��]F��q7|݁䀻Ǵ�*����k�x��]o�����~�������;~��q�fj*V�����t)A0.U[^f
&�g�Wb]����5����U�˯��W�ܫ���/�BV��>"�&�N��u�D,w3�F�'®:@s���*8��wMO!(s�~���<ppWv1�����x���ѡd;�Ŧ+��C�0�M��>��!���_�iĦ�Y^R+L�D�8}9�E�َ�z�w_f�|��BHW׾���^z�0�������q�_!�4��u��P���y�~y�}�`?4@�N"��x@7�ހ�^�;ݛ��X/RO��=��0��{�2�x5JD[��8����g�n����ޮ1�,�0����+���uLA��x�K2�^S�ϋ��
��R�n���(��m�����o��"䫺pO�zȵO�^!mX��_3�զ�k�Tt���X�)O6�Hx r}{��~���r�3���+�y�*1�]IR�~K��*�j:��]ח�w�pS5�i�K���+�V��k����XH�H~���z�ַ��m�(:h.��}�,y�������H3^��ݍ�| Q� S�E��!���;����[�o�(+b�~��5d`8���j���������+ĩ���?��j�����~�M6�y�T��[S�����A�QJ��Ќ)iJu���S�W�����b�Eщ�.��$�W����X��ߣ�|V�&#�~��zQ���+���%yER��T�I�����D�U{G�^����^H`J����K�L�T��Xr�g��'ۆ:��\b����
�oU������@��O��X�U��J��+F!z;WN���7F�y�4�}y  ��X�B#�бS��w��Ӡ]Fo�\j�O:��k���S1�x:��\�=bQ
�����4~������ĈM�euz��pn_��a�������KS���(@����Q��)�NJlJ�=��0�Y#��أ���¥a�@C$2tV�S4�vLq�^5B��������w��{�� ���Ģ� c K[�����~��z�ɮ�ͣ-î�`gγ��0b�j3���O{ܮ�?{o���T����׹�n8�J�ik�4o6Bzy�;ۂ��<S"��xB�'
6k|e�o����H��[j�A@Q�	����r�vd��T�N5��d�5�II��FQd��n��U*.�����展b�R��=��{�*�m��p�R���ᰠ�� +��X)�D��*�T�ڷ�j�Q�;=�J���<��ʬg^.��Ny� �����CC�z+��,��!��
xB�|� �2���,&�p	
f��*S��kY^�ۣ�Vt�"�a��M�_�f�VƂ4+����˹�{P@�_"��rٶ������)�Sv�-� U�/�ÎVh�{�#_����?M5��==���iA��_|n�;�)���XhO(C�\=6�`��+��PU��m�K�:#��t����W��)uj4QY�_Y�h�z闞F��y�
>u�Y�����2� ˝V�m�\��P���[���)h"� ?
�����(= D4}�Պvc|���n��Ƨ�7[c�9;����7�~~.����Cg���G\0ȬE�N��ܪhM���4���­����)qu����C�t�K�xO�S�=�yaڃ��.�ޛ��_��j�+��W������!�S�ߝ��<:k��r$	�oH�����w��n0{n��S�������P�������5y嫂���v�����EY��:��ۥ��4lL�6o��]gO�,@�3C�ZءU�B><�L��t���ֽ �yי�.���.� u��k����^�sm@��)�J�!��B��/.�oV�"�����\���](vV@[#ӛ���Z,H������giw���G;^�!9����!���z�EڕG�m���.��C������]�I'�o5�˩N:2J���Q��}*��mp����;����UK�����Z���)���֝

���V�`��g�S�y��jk����&��>�$��+c�YQ���`czoy�:�P�MQ4x����9U�󊘣C�>��>����׽��Y����߸��Txwύzz�������]q�c�?�hq�>�`ogC�	0z�
��j��m�����u�Jet�F4*��TU��r)[	���'c,��@|F]L�c=��/2;H�^��o83	HJ�rg�U׏fx
g�2���٩,��F�V6_�����YY��7�5Lz� l:&��4��p�%�c�$иp��yes�bUw�f�pw|a�F�t�&��B�0�Ee��|��n'2�y�9̱Hb��"V��h#��+U��OB��-f�tm�*و%!�o�1Mk�l@v��䉘��|G�i�������7�U�̲}TUC+�k��Q9>İ��ڰ}�(�纫a��  �]�q�o���4dt_��H|�^�����'��+�yW7�ֈU��������d&��:.��?}�<��O�CJ�!*��.�T��
45���8�v7a�z��![Ʒ?T��(>tH'8�,!��'3�Q�W���k��/ .i]���Y]���'Q��P��5�]�7
X�-\~(w��oH�ˎ�p�yѼ|r���6��t���#��Ojp<Nj�J�22���uԻu��v�:a^����A�1`㻴���i���y:WDn�p�6s�!�S(�P�w��;u���5�X`�Ή9q{�ؐ. $F ��e�Д7�P�G�t��<=��/��o6�J!��^��|h�?�zd$�,լ~�	���K]ѻ��_:^����G+�W��0���;�������#ҁ�De�v":���CX',�Z�
�f���q�>6�mR�9����q��f�B/iΜ3�mL̊�P��[�7��n!����cн1v0����� ��)UC5L������.�h�K~�};�3G5l�20*3."W�}���m1R�<?짱(1@پ*�fo��2�)�(�l&�̇�ϺG��̠� �wxd�Q�_��1N�b�]c(+�z��Z~���4�'��R<���.PXp���Y���%�Svu��/�Y�5��F��^Ej�cՌ	�#��Yrς��4o�?e��M�ˌ����L��c�K Do�y�l�We�V��/d��Ԕ�Q��Д���T������D=α�������@�x�{^֘�F^&?v�J������/L��G�.G�������{�s����(
|���k�F��Y���}M�^�=Kj�� �����x�{��%�d6�uv���(k���E9EZE��N��L.�::V]��X��E҄�����ɍ�l�����tME��k�aܬ�кy�������up������]�K��=��z�K�J��غ�W�+e[P�m����;9p��ܑէ����.u*u�Ot�\ANE��fdU���ǛB�6����z��@���6���G���I��?K���b�j�wt�e��>�klW}�@��Qm-��aT���xw���E������yԚ�}�em_Rk�%X���fg0b3�v��ԫ�5(�/��P��t�R&�G�ñ袣����%�ڳ�,�n�Êʜ0. ���3��(��{ :���A���tV�R�lK�)s���7+R|�Ρ���5w��R�� ���b�n��}o���{���T�U���{OPޚ0��wf��d���4]�"��"�hޠ��ǩu�����\x�:�;��<�#T�0'�e�w��l�����ԥz����/�6u.���KV��L)˭+�`_�����YMY̡`q�o�̝�6NGhU�|�q�ó&��S��~�3��p}�/�v��u�6mL��X]���X.�-&����PK��м킭�!����z�	����]|�o'gPSmu����M���Zv[CE��:���0��h��ok��W:X�9�W&Iۮ�=}v���um�6*��������]ëy�rLX�=�X+i�2q�"}5p�<�ܭ���[w�� m�,�] �
���1T�K��\z�����:kĻee���\� �[X�`����ƺP���!��nK�q0��)=�ͻ�t�ܡ2Q���[�9�9OɳA�th��u��w��x�;]�̘����5z#��*����ۮ��X����Ft�.�x�ۗ��E�CA�a�>�V.���Ө&T�س| sW�u����z[�.���&*�9�Q�m��̺�ܹ�����$�2�ќ�����W��fqOVkP�]6���c�k�����]��]�|,˼�X��%GH�kT7�r�ƚŚ5ѷ�RJ%���ŷ\��Є%M�ي7�M'S�m����&�qdK:u����1w���6��Zrbڽs���t�|yۓ[�/�v������k�HP,�k+��s�4��v�.c�U0'�� ���j	�/]`�
Z���ƺn�Fl�D�n}�{�  !��e�|�7Y��ٺ��tE��W�ل፳���RO�sL]��q2wL\����F7W +vX�]�3��wVl��H�w5Rݞ7�3"�L�}*���'�*���g��܌�����>4�H˙�������Wt���X(�i|D��i���c�\Ai(���M{���Ԝ�̸�-�����7�?�*�Y�MU �rc�	9?����@%�H�E{�'�yΠ�>;���E�qbͭ�|���Y^R7^O~A�^�Z����kCl�X�u<����^��Jo�+�ۑ
E����E��}e�2�-�xA�{�p>�*A^ڢ��C׋:��Gbݼ��1�ϯ�Pϐ��s��ͽ.�d�A.�����D���(� �ؘ�{4���:W�q����#9B
�P�u[wI�(���y�:ԂWk���J9��v����1ǜd�K)�w�I8��}&Wwd���WE���}������mg��D�B��G(	Y�wv�LW�V5b"*��u]U��X��y�eÅ�ឳq���/#d|Y'Z�xwM������[H��jN=�f�^L�Q�d���N$�H���|ǶTeu��Iq>���9�|�X�D#wc����K��5)Oz}$e�)���� H�:�A��%��:uBFE��PTMg���G��x�����DNoU�Z�7��*�G��G�w+�0<�9�H@Ą�̆toQ����*��Vw���С��$�)����mEѫ�ʉ�O�9}:����k��u�#K)������7���5���_E�泎��s����k�"x=������Ȉ�\;�hT}u���D��_<�qܮ:f�LLW����܂*ە������$F���R�#�[��VF�f�Ua�w�u���;S,[�4���<w��ɺ��N�.�F[-���a���!t@wf�n4��8Rލ�띓7 ��/X�`_i*ޭ���F���q���Qsѷ��}u��g���ê�3>��=�w����ʑa���A�ֆТ��,�ϙ�(�|�;AM:��a�L�8RQl��@ۃ�;�N򞜵,�!-�ޔU�C���Хɢ���+�����-_�W4=����';����0�	j9��x�z��B���}���/��:@����^C���D�s1�'\{��} )��+`|�Ě�_}]M����&�>
���O�O�2�۳�cQ{/4;�h6��˨����N���cXq�>�c�y3<!"�;55P��@��8׽�TB���u��'��wG'�3��O�Ѿ��PTH��">�#�(r�qv��~�}��R�5+(��c���a���$�����Y�zء6.^?I�aM���g�8Y�����?o�LH�<r���нu8��[���W�%`�KT4��G2�_�I]�f���]���a?@��+���̈́��\�����J��>t���XD]��$=�ə!��\mk)*��!eBqp��<��*�^��&R�y��N��E�+���F>���BQ�j�M�M�B�!���D��
�1�N�qI丢�$ߝ���0Y$q��o뾠mQ��A������Ma�)8�A�(Q�waYu���Z��x0���c�*���^gcLWs�y���o���W�n���%;�L�^��Ao�rb�s'�Ջ�Y���I�u�ws��V{�uZd?g^�=������ũY��˹���eD�{]/M��N(��&h8��[��a�V&���r��ná�K{��%��:���F�͹m\��Ե���+ER<��ޅ��/%m�TUw��\kl|w~Y���
u��j�?CH~'��7�(F���" �gLIC0�p�Y|�w��[0�����n�a�Π�nx��F;�E@t2�D��??\#�Ą5B�_��!�
���^�J��"W�W�����?�~!��Թ��dS��H��� �ZŰ�/�[���E��B�(n�=*�m!�A�����d�
8��.ɼ󬴨�G�&r�r��s��*�x�0+�Є�㝺q���^��q ��.ꙹ�}��K"������Zw�/�B)��tQ#D����S�G3*���*�F4h)|����ŎԸ�+��4﮹���"�'���l˱�{�u�ڹ�6
۳7ֲ�Eњ*�@^l�<�D~�����,ʘ��ۇ��0h-��n��n������c}j6�:�����}�J���AS��m���2)+����0�,)��zg�4\;�!�ݢ�a��N��c���CwT�8L�c�o��e�o�B���`��%�Q�|*=���ҭ�NǴWH/��B��s
UA���L��UvH�M�cz��&_@�~��nU@���*u,f�5%��z�����MOx�(�����x�[j^9>��ۓ$��} ځ��S8�*.������LM_�5�����О%���κ�僀<~3}n�M�4"�9�.�K�{@���_�7��}\.�_����z~��a���b�ጵ61V��x:�_6��M���Rf?�Vմ��js�R�;*z�Ss�ݷn��ە�l�|T[;3�O�uD�/Vc�CB�/�lCֆn���,��]���Yƶ���,��3�P�� ��r�'e����"ѹ�l�o�=��������=�b�lS��⸸�>[�t�#�&c��V[���3T��p�U���mC�E��q�g&�n1+�`���8����h#�%�f�n��X�VQ�]����믾�t0=~�����?}.\]�]��=@��I��KɎ�.�A���}O��\��W�9�s���T�̽���zꃐM�8�l�[*a�y�q��녞�3UnVj潓Bk�'�f��Kz:rI�]=¾W������cKY<�94�A672n����A6q]fB�M�R��׷2���"��9!~N�Rei�x���s<7�<�ke�~�;���$�H��r[�lo�&9X��ae�G׼D��G&*^�Xf���<�K�=�)����p{��ȩN���?ֿo�z�7���]��d��J�7����>�" �y�@��f�azF�OB^D�7���.9�
�V9��U
:*j3˦�w�I9r�����P��j:�>�I���}>��u�R��˜34B$m�=\�0�$7�њ{++�b�;jpP�i��ZG#p���+������J<MZ�,�(]-�
����D{���c�"��B�[V�[
&��۱�aӽS��Q�+�����+[M@=x@����y������{�Aۉ�XWW�v�I*��.��5yG0*R��6GՀ�E�q��#i��WLò04j+Wp�\f�I���	�2�C���Z�q�Q�ܷ��y�j��k0=�������I�(<�/f%J����������]e_V�a��V땊8G�/�$���U�m�fh[
:];�n�����P̣ޭ��0^3�Y]j�XB��l����ݸ��{�κ�X�p�^BU�����轳}���"����	E����TB�L�G���~���\ǀ>��S���]
�Z�b�f ���N�f�u�_.����*�g��v��}�>�Pc\A��3R��E#�/!���3�v����e��YO3L!<i����_%�H�O�>製}5N�R#3�dߚ�P��!n��::�q��b�q۩�@����aϑڲR��o�_��z��hh�ez��n��쒳�?��	����M��L?�"�����?AC���T��ɺ�땪���ȡ?f��߮ϼК���f�aֱ�XG�,tcy���fg`���m}jZ������^TI����`���4Y<+)�Ms=ޕ�T�e5�Xyne^/(>sł ����o��dr�-DFgb�����18��]t7��cǼ(gm#>P�[J��t�s�s>�m�&�N�?'����q��Y{�'N�d{���'Kܹ�jws{�BT�����3��R��`�����j
����q����������e򋫪j�U3�tCV�`w+Of���[i��/�:ψ(~�����`��;����i�~B����^�d߷gf�{L޼8�=��+�)DW�|ꑡi{��d�(���!^�)���'$�:�$~	B���XDɒ�=ڬMY�o���8ۉ��Vw6C���~���C�ݜTʮ�:[�����lQ-'����x��+���WN�ӹ�������oks�P�$��qú�6x��U�W\*Gz;��]r�Z�unUV��c�.�<鯅�c��q�+���$n��ʡ\硽3�|^�U;c�X���]���ǶEF#�����%\[��kc`U��z���� Щ�]� ���ϝ�Ҹ������ɭ$7����k�z�t�z*�ꞙV@�<n�?,ʚ#�b�6��%0�~�fT�������=�n����xE�Z(-t4�����<YM5�V��8��Z�E��U1K��yJ^�]�sE�J�N���-�X�u���s槡����c`.�#�^P��U�2W0�N�vO��=W�Ϣ&Dmy�K�\�*\�̊�{r���dA��bb5/�u� �ɪ)/����ܶ��2�j�;n��P��tTv�/:HY;f�,$��,F��^�l{h�{��5�&�y����;�����P��r�_��W�ό~֞~�(/Y�1��WA�귗{���#��ݠ�����w{bA[l��w�t�
��dm^iR=�xgb"�.܊*�Q1`��S���LO�*0�q�]sF��:��MM���b����^�{�S_<��jʁl;�	��/����5�1��<&;�R�*����\���.0�Z��Ǘ}���OA������S��~���;�"��'uv��YU �O�W�~՞K����yƎa���+��<Jq��<T�Ay���?1�e��Ǟ2��y���`�
U|�,{7t�%I��9��hB+�K&L;�����f��Ȏ�	c�ǘ'�k9տn�=��î���H.\�uF{J�+�ΐ��6�h����x�_�w�8��\��{�Gu'�own�l�ᡦp����0sz/!ɡ~�迓���F�����I�炟��C����li�딫���ysz8V�ޝ�{�\U�p-v՚��NpU���P���a_Xx6Aw�j"=+�5�lI*whTE�ֽ��F�!�tgGN�J@wB�tV��1Z�k�s�EM����C�Xu��˧v�7�G{hݪ{�['%Z�T����;?y��f�H���V�����$r��)[�8��y
���W#gٕ9�L漒��M�٘o���۶۸Qd��tӭ����/`�#�w�W�Gu��3*ߨ,3�vi�v:��|��Ee��p�6D�]dC�N���>.C��wd;�.$.Q��3 ����O,.3�&��������;X�߸P�e����_g�)]�QLVaJ�F�����uZ�(Aͺ�>H8���f4v�r=��}ƽ�qo��z�'+R��YC�u[��4�맾r�E�Q�Ag"����I# �x)ܨ�f�6S��\U}zm���\���I��~�ɲ��5�����*C���_�_J.�����vN��"o*~���=�Cb� L �]u�|މ��4d�ag9�
��ʜ�͇0:^z�'O��ghsC�.�Oq����ӑ�[\�i�����s������v���~wh��<v�
pK����}�H�� �;��g*�ux�xV���F헫�81�t�S:R��k���gs��n1��H��x��ƜZ a���V��v]C]܅��Z�\��t{R���f�h̔�G��_f���:1�!��u������S�J&y��*I�zv�=�ь�qs�ը� pypHS�w���@2�������~`{����ʩ�V�J}	ǠHc����2�9��Kq�q�<6D�~tlf��e�m�X��}uA�����qK��� ��+݆\I�WKK��r�`�\��R<í�]��L�X�L�b��i�LY��K�p3~���&�ƅ/W3KP���Y'SٜPs霣YG6&�����'i�ﴷ�y����j�p�1z��ct�_��P���)4-y�'*��V�#��q	��̹��jnL�^���K[\��X�LY����P����}]�s�=���^���t�����'؆�)*��}c�� (	���r�֊��˫]�A�K�r�J8��_�P�otƾ�z��<��⢭�r_V��+�8�/L�yT�O�J��_M�Ĩ\�0��Ԍ��Ȋ��J��$#;�A�\�q��U�f�c�n�gQS�Dw��lNRD�g���׋���F_��������o�B����1��$A��j��=��K>�v�b�����9
F=�Wޟ�������ؐH�<��Gz}@� �]'��Q�&B��-n�,���,���m���KH�T��Y��{Ϊd2�M�[�jU�^cB(�p,����s0|A�����9�M�|�&�h��#I��W{Qn�ٷ,�E�T��gu��3��Fm[A�+�R�j�V��c�ń�ip�(�V��)�T��y?pbc����:�Knft�J�+]�	����w��X����`������t&�o%�n�*�Ⱥ����;�Fl��AnĎ�}'�^��y"��->j��N�+ؿ_Ɲ
��B�z�G{<�CU΋�,�oܓ���T��r�X��mC"ph���f ���k��j�Y��o�D�Q�n�^��y����҂����G��ه�_e����`���0Q���_���~�}��U߬�׽OM6%D�u W@��N����;�nd�	Y�.�P_H;�z� ��`��+�Լ�30}���O�e}ec����������
�Wwp�[7��Zyk��X���<���rؗ�hm(d�HL�^�V���A��o#��@54�W�f�	��C�0�#�8��B�V�w�
.5N���V�.DNu�9Tt�T/��*롲3�Ռ���7nOy�F���_.��v�S�m�	��S�F�иI}�Mܹ�u��L���ēj�FX��۱�DL{�n��~���-N�;��fMǼ:�1v&�{�yæ5E/�J?��/Mo��H�oK���k0�A*�7F��}`���~�h�������	��C���kA�#�oa�{dѭ�y�@� �`�ٮ�ʜ�5+o-�ρ�=E���X8"��]7[bO�SM�r5mp����Vgr��r��&�ړ��W>�:!<k �O�%*R��&������(�Ƈc�����پ4��.�u���}��޹g���p4��De_2K�������r���w'���,D4j[-�r�A�]�5��wc��K����案܍WZ���]��uΔҍ�� ���v�I����lݶ'Y��`�����9���>�;�¡���X�kت�T�t��ȳ��$�e�>[.�d��h�e뱚h�Ҹ�R%Y��E7��*���f]�K���-!��BS�]��N������h=��tJ��^�=@��Đ;
�˫�\��tk�1���V���?#!O�#쨉~[����4��2��'6�XBB]~N6���c�g�aihF�\F��YO�ϑ��a�G�̏�y1�=�����,j:����T� ���Y:B^��
Y���L�NJ�Q�<��)�E��`0<FY.M�H%���Pb^��'�\ŭ�V�5��z�!���\QΑ�a=���zA?N!�"uz{��q�7(-2���~�=�@�f<����-����q�shN�v"oT	�&�{6l����7�WE�����d׺��0S��V�����e3Z���j�Ώ��f��=3�K*���'ט����[����.��ְ�X"�.���C��U���LO���ϻE�����J���EJ	�V�q�K���1��H32�g&�l\Y�^��[��;�͎�Bc!E�N��������o�)��k7�I������Ag}L���y�� �hCaƓy躨�Եؓ�s^"�1�"ی��3����*"����3�;ԝ��$:�
�3�6ia����I�쵊�2J��aY��K�@�0e�N�s$��t�QV�;��=w��!۳Np�]F.̓���\9�8�c`oc�D=���T;4N�I	�(�-��k=���?��6ڋ[K	M]jL�k&=��a�IXS�ܹ�$��9w��om!#��y���L�ۅ�-�wD]Oٽd���+z�Z�1�o,�;�f6�rc{�]1���̧ï(���҄��3��HVP�C#����qT{l��Y��ɜ2kP)h�LWZMX�2M��cW��FB8��ZK��Ҝ�;�x�#�����ꚻ��*7�1�6{�\p\�f��F�X�wGV��jP#�)
Fh�ꋥr�;1>˫���9��q6T��S��M^@�y�i�\�볤;�0]ǧ�ܵh�a⮧-�x'��L+��lu4S��7�8e!ݚ9թ�u�VU�,/�h�M���!�ko�<st���ɑ]	�$˷�ʑ�y�՞��H��k�J�Y�x��]D��v���������N;�7����y�O+�D�q��ƻ�JI�C;I�	u*�%�t�<�˥��
f����S�k��J�d�x�v�:��b����+۶䷏c�2k���n��A&���*L'��ć0�tդ�c�fPj�A�uR������Y�ЗH����\R�`��1��p�i�{HW�
ݲ�}HkC��԰���z�թ�fA��D�0�;�����V��ޤS�W;�i�=� 
�6�c����9v��^v�o�VsC6�թ�p˸�v����64�c6�.�w+�`�6[g��׾�ׁl~9��:e1�Y˗N��s�0Ñ���ȧ-!)�PŸb2�qcҭ��C���Xm��γ��9�o�n]�ك�|�.����H��V�J�]�f�h��	����SM_I�K�f^o�a�j���\�hehiZt���Z�V���{�:;\�#8�g�N��)�u�(ε�N�id�c9���z�NCc�=�u=�+**��ק���j ���z���]]��F�r�|�ٕ��]�@�{���)[zr��!��o��jU�i�Nf.�׏\m�N�^P�I�9�՛��	r�I7��NM~!̭t2.�A�!�	w��?G(���y�x�j��72וٙ;j�LAl:�˰�Sά�_l�K'f����m7]X*t�mr�4���`���nGt��������s��o���F�����C���m?�J|X-��'Prf�/2ԑ����fvE���v��k�c��w���g�>O������Y�1�>��4=�u���V��Uf��-�=� 9��[t�'��J��Cj]�{�r�.uLՏe(�պo2��-N+F��Y��)��+��Ю-���";��\���r��h⇭�ʷ�7��x������;���<=������k��19�I��U*�$m�O{�m-�a(�h=4�#Н���r�F��8l۴5L�F.��/��x7,���~r&�yf��w�j�ѝV(�\V��r,�ȼ$tQ(]:�q�Vei=�W�xG�S;��oLu������REW�=#��j6䉚�p�0m+�^��+ߏ�y��n*��ә!]:�s%��S�2AϹ('Ҧ#%�_�� �`!���ʧy���S�O�/7�K=��V�T�Q�C����F
�9����m{�N2f}�;�F���D��=Z��N��B����=�Rs�f�Ò�R|�eZ��f�yY�V5}�a�Z�Ձ%��%(
�՟�ȩ��B�K� �� avt�?G��b�u�>��������3=	2���� ����9b�UcW�r���wk#�lI�Zצ��G矂l�*r!�"��v��l0�һԄ.���Y�	�����j(t�Z��9���rf�<k}9���ŭލ�?XZ�Ȩy��f���G^5;�sܕe��������Od��bM �����l�Q�d��Yʣ���3 ]=�nK�Y�7w�mРGy�B�G}��:��w�\+0�쾪��ؒ�xE-����ۊNcݑ�+�n̾�����ZB���7���{�yD�r�o�P�{�fj ;�����-t|�l'-��Q��_B,�Ȇ�ʂ�S�W�5w���u�T2?��l%a.^d�\��^v�;����a�܀y�o�uj�0�G�:�[q�͡ZPz��R�+	�n�<�Tؚq����v�2�����RV=�2�ЈĶ%�fL�o9ȝ���]�Ж'@����1�R}>~F&�3�!�1����Udu{��0j�eejޤ��4g�������5��+�|�U�gٕdu�YM�a������޵k�������{"V^����l��ʌ%��Tu�.c�f��=1-O?�ބ$�)�ڛe��-��e��r�qY�ʄ ��k���=�]�,���G/K��	�ϗC|/��g��G�z��\����+���ق��$��Cs�e:_?CQd��ԉ*n\��Lq�>�ћr�M|[���$�i37w�/�����L�ڃ-��܉��.^���N�|�O�5���o�����V|�v�w�Uf=�+��&���,ڇ�y�v��R�}� }��!�}�sٹ-�U��j��VCB���E���i|`�&F�W�ƪ�\����C*�=n���rV#Q�t@?=*a�`���[�����?E[͛{���f���y��$f-5������YS5�ѱ��7Wu%�;20�܈�c����g�������0���y�Ž�..��Ust+��� ��uQT��9���&����&6�����[���L�:��vD<^�̃˼�k�n^���@}��-Iw��,��m:�o>�V<id<Us�XJ�W딴_�3�C�0�vo��V��\׵C�t�td�|�Wm�W��R`wD��.�V�U�}.��h"�\��{�iG8���)�S�A���\'rlTWz{.��p�?M�6��&kr�K0��C�b��]�w���jv��TT��/[��t�ut�W�}6�#�sND�O=�| �wf��m�����LI��B��ػ�R��l�'�ٲ!�]�R��iEHu&�S���j�mc�fr��bse��o0ߊ
ȭ��T�@�F�[��wk�qa���J,"���N��l�V�J����W׆�b�sx���H������j:��.��3�	4�����H���4P�s-=���9Ddy����f2��9�}6��,ma�����2m1<��[�/H���2�2	Ub��C�����1���i+���V����aC&M�93��5'n�l�}<ڭ�=��̙�}t���S�Wzy~b3j�db�:�#^w�yN��e�}C�Ԏ�V�%�P�n7��88>��}�'xQ����.Ao��v7��?�m\���t!�ӊ��b�
˲�a?����Cp�rfo��;�Q��o}z#e���ݷ
6ϥ�l�|1O��-&{��mEWL�v/#w[�ȷ���8�����7����h�SB��u
���fn(1#6c��tbO���O��
}U5Rb^Mr7,DL�l�Oڗ�	�{lFg!h�����mҎ���n��{5#'����f�U?��De���v�&�V~��aX��Qky>�����*�SʮEiG��e�[�o#2�8����%u1�Б1��s�:����u)�,<//%^;	F&So,�<�[�xc�]nL���z���^��<��
�4.��]�S�c)	�����~+�����r�|���/�ۏdӹ�"�/�K�a)���=�վu~z��� v'Qe���W����3��,��U�Z'x�D��^�#9���}1�Дc�+�٘���*�׺�Y���=��p2��fU�������q�gƔ�~�����&E8�{2A�/�M����̭y��0�UC"bڽ=[��U� ��_<+M���kŕ*ߙ0�����0�7�[֦!��3���e;�eѥ�](�*�y����xȿo��>|����+)Ĉ3U6NWA����]({Q�{8y�i���g�gc���ys�83�	�x��n4,�M^�]�5�C����}�Z��������W��%�I���/��ogNVGoU��l8�������3i프5T�}��93#Ik�2{iޕ��_n�=�1ee��G5U�3R���w_;�������W�A�N���͋ΊI��햠�gU��ciZ4��k��ϝ=	�� }�A����׮�ek�S"�^��grq��!�@�s���j"jݟ?�g� r���ؘ�VE�_a�s(A�_^[��s���b��1Q8�R�j&Ƨ�S�T��Cbl�(��c��dX�Y��䛛̮ҌS/J뫴:xsq{���~�\vUĊ���\Oq���xm���{դfʙ�������a�Ӕnݷz��q�\�y�ݜ2N�l)�ɇ����NY-Fm;]9jt���������6��ɜv3���ӎ4q��)��H�<e6�ڇ�*[��{{��J{nz':}t1��c<�
ʉ�<�C���=G{k��覲ų�BVJ�I>����ԗ/��k���aS�k��?�����M�p �T��[>b������)�����G��fX��,�˅���h���E����p�t(@�$����һM�/�LWfV���	,^��������Zk͗��;8���~�~�ʚ3�n�
 ��Wڲ`W�bxp��(*���Vs��H��z��æ���*�Ӂȩ.��??I�:W�8J]��YaA��l�ܟwY�c&���dN��S�b�*.�Ly¾�zD�=�P��^���J�
����0��!+���7n����uvz���?&
���W����A��p�"E������������a/}N=��N�^D��7����o�����S�U�Jb�J���AR�˽v21�r�@��~{��3(H�����/0`�W{��k��D�Wٶ�Ÿ�����{V��;�^Zvy����t�,iF���q�$~��h.���\�����Ge��'u�n.�B�_����pL�ޱC{ޢc�{�#�5G���>�����v/�3�Ud�ڢ�����U���J����E���C���p�0cU��Y�s��_mc����AY�� Y�[І�g\|y��W\1W:��A��T�<�GS۴Y�7,sB��?i�}V��;�bN޽�ʷÍ�v�:ﶄ�:��lb4f�Ǻ�n]k�AҊ�6�:�>y���U��_࿨b�zi��y=���p�����|;���J�GjXQ�,;{�����4���2�Yy�[��|c��}^�8{[��^c�@��c���{2���\�ߥ�"�?B�&��v��$OݣZ���f4��uO{|��Ԉ�(�g;�-�>ҫ嘟�(Ԕ��m}r8��"���݅1�1���E�Ѯ��ct�/	��e�fP�3G���]uZ81����wq3,\cֺ����)Q{��r7�s�c�r�����&hŤ/m`˺�r�9�.y���;c����;�:=<%i
�`WnC���t���b/f�P�U�]� �t�w5j|Jy^:9�R��'��!�nX�/iWò���՚WW��V��̟����=Z�j/� �7����pg����j���>�����r��g��+\ﾣ�Hv�'۩�9:�����{�8�����>���]z�d>�JԌk/i�n��ǖײ�5O�W���wכhG���
t�]&�S���݊u�@��и���p��M�gڽ��G钴��loFg`W��x�a���2Ķ�]�'S̑i1��Ny��R���@��z{s<~�*6��U���K��_i[�D���Uu7�]Bs K�x�U"��;�bv�]yZ��<X���:~�#J*<����f��TQ�, X��N\՘��Z�oy#�=�w�3�C9Űբ�D'M�g����-�1<��$��t���2��t�����W#]Z�Q+�مz��(`��F*�Y����,gd���mz������ߨ����|����r�{����}\B�L�0�%<jLF��N��̚�q�$B<�ď:�=���rc��3[�4����X6�]p[��GtOmj��5UK��j}����H��#,ŸX�ӑ�cF��=�a��O\h����0"�J�F�x���"��.�����b��9�K{_i���M�'�瑩�9��VW�S۷�7$��S�d{���r���^@+#oqx�v�3��m��	F�3]�
���L���#��@��yVҬ������%�Mi�>z�Y��q�/�6���yj���@�m�e0�'KG�{��_}�𡅫�s�ĥ{��y�	^w�Ў�NٍY.%n��F�r��ȶ�s�N��p���X�iJ������#�H�}��]��/�v�l�zT��ъN�B����}��H��8�4�1[�B�^e�CC����uvq;̓/4�s�w+B�]�G�y�t�0��V�_��!�2����`I1��{t=N���q/U�rn4Uw1F37!>���wM�v��#6��D��YT���uH��~Oh�����"Ň���GՂK���� 9��C�ۘ��ދ�
>x�ef?ppfХx(�#m;l7��0^��xnE�@�]A�c{ѧ]f�_\������ r�n�mr���V�a��y�a���>5:���%J�k�_\-�'�2n�2�%�'�M]cnG˺����6��!��싔k"~��L��z|�A��7�W�����L9�f�n.����C��#k��MA�����Ϫ#��am���V	5[��IB�:~��xI��f�KP�>a@g�:|��g~+�nG8]0R�C{[�P4q<#�� ~��zk�k9�����)�hG�ttE�[7�}�q�83Z�wJ�r<	T��&l���������:���f����N}���:��t��
}��stk82c������=���~��l&{�ʃ*��!��h=ʻ��{9�9�E�	�)��~)>�7W�x�+���g��0�B�B�H�xn'��ꊃ���7�� E�f{�����n�n"�����K�c��.�i���fk�ds�9jE��u��y�ѵ�U>@\��\���عS_�m7�^?c�C������9/��O������@��ӱ/P�-�ʛ5�pֲ�_��M_��6o�[�%�}Q�+�Þ��+�b+�}��TP���քN=~��ʗ�.i��'��� ��E��Y�yН�Į��p��4#'7���6�P���26T�s��LR02nk���OMU�T�_�g#�^��#�z�s"�,t]�]4��A�\|o�U��\����L�)��mu/a�f��y��ǽ�ʕgy�n2[c�e_k"�t�*=IM��r�Q��e�	Oe�x�^X]\�1\m�S�:�Ś�D���0⯳E&���Y俬8|$�~��^i��|�d��Q0;[�k�OW,t�WNeWQ��z7z��Y��]/���6=⾫��мs�{
.��^x���s�WW��k"��f��lr���~�h��.�~ˉ����H��W\u�gQ��js��+T��a��0�9���Dh.z���&b-�������=Q�26�j~����J3� �c0O�����(EN�خ�ǕO����iJ���N���3�n���%�9w;�p#�WHŖ���{R���o�ͰǞ]h<����Ż:�C�h�3�����Q���g����4�Rwe����Eq�'ƣ|���K�|fB�-�O9���"����nWQ�bZkj�_&��\�a)���̣uO�O��r����\��U�3k�Z؃Oc/���]֜�I�pyBj0	�Q)�~���_k�<6q�M<r;O��ʍ�GfqQ��m�U=�B�&T�x��;'�f�}[� �\d~*�GvБ�R{��GAT��f��̜��21�L�r)i��Ϊ�_<׃;d�4�����s.m������i�}�t�Gx;�sCF�4P��moOڋ�t�?U�9���,�;,��rW�Ķ]�sL���m���u/S=3of�v(O]�x1]���Yg�L�t��fT�U��*���x٬53�r�(Ex?�x�jxs��sB����b����ھs2�U��egh�{A]�c�&�u���Hŕ�G�Ʒ��f��C�'���ƪ;TU��?�B�t��1�W��J||����Q�-�&��*�!�f��8�z_�����H��'W�Hz��C�"�����W>-�>�a�B嬘:���������o���>�W��J��j�s��v��w]��A�6,L���	����ԮP�	�V�m�eTv���������*u'����Fc�oǕW3�s<XQƾ��{+%E{�;���sλ�������0^c�h���t�^�xU��ӳ���tg��"����O�����y�j��R�4`tm���:U��9��-s�s�FEb��3��O�C�33�J�A�6����-�'�ԭ�t�։�3�W��f�=�v��u���)`�������u���|i+�̵�}���g������_!�C��֮����s�����Y�z<��A�xodo�w�R~�w���~���e�¦��F�4@ؾ�zɔ�Fol�]x;��x�@W��H�����0��>�fh��̑ٱ#<���9���*e 2�˶|`_D��ǜ>�v>o��ϗ'^��까�T����N�t�K�;�D�I�cƽ`�P��\��� lXsľ�;�?bo�f�+*#V�
��D7��.�Dۣ��%c���,U��	���ݺJ��)sBT���8=�0�U���<�Vo�5}ȣ��*�뮩�S��i�(ؑJ�x`����T�1ű���\���5.������5f8��!���J��ou��¦%��Ճ�-1�t��$*��0�		*N��j�:�Pe�X�*�t��]}��`��N� F�3:�oz�I�\����On=k�E���e;x+���9~�����d�|'`�t� �d������P���(�4�~���i�C��ͨG&��aP@x�ʗN�ؗ�Յ�9\X��j�L�SIm[�Z�R3x��(j[��~Om��'�!ٷ$�nҬ� oG8�*��� ���ձ@�T]Vgp�'w��} �e0��8%
վ��+�gbݕ,Q����%�C=����]�uN�7�Q��,^�
Q�>� JgzA�?M���b荱6K���L��X��[��h����w�p:�e��-�3�Cb�j�_ID���ȶ��1\��6z�ʜ4GG��L��S3�#��-��EvN&F�.�'O1�d��^3�wl�v̢;�[k������]ͻI��Y�ǗY����w*���5Xյ揯���Iܻ|�ٻ��Q�y���<l]�A3���,����I�]F�/���tWi��j��Ctv�]2��G�T0�n����6�7B]�EY��i�	���
r��Taa�P);�z]�[�t�z�d2%�m�����(�w�-���@S����_�I`���I���S�R�1SE��N!�l�yC����Գ�gAWan� �͔z�LyHz��Ok}���C`�.���?��A	LX1t|7lɜ����=�����VcV��Ǭ2���R2���Ea�����n���|�%:��ٷHӫ U�#{����dB�L
բ��7$WY���8�h�J[�û7;;d4H�f��,J�NK���cD�"J�2��B�zm7GS/@jݭ�����O�=S�:/xnU��&($�uR�a�M�eH� �%V�	��!t�1�+�.����=�>����3�bOA���[ �+kZ4a����:�LN���QBL{�}%#ώb�YxF���.�!z�B���_�|��F��
���(o�Bq~�[G�N�Gd�x�C���(�'XK��ʘ����f��
�!��R�(@�졂u2�� ��̬|��8n\�,�[Ahw�*S�f�I�Z��_�%*�u�A��WF�p�+&Uz��ڔ�j�\�[/����&�_R�v\�81os��ЛF.jh�s�� �����kE݌1�ׯ]h��
���Xk:2괍|N�jW=��[		2_ieW!K�_���fc�S{[�K^p{Zԩi
�*e������om��/�����6����/P�ל�˝a�偃t���a�^��Tn�L6h��Akp>$!����ȶұ̖���!����+�G��Y�a o����Ȼ�
�zp4qV��r�YK���aTc����r���TדA��E�ry)�y�Ƌ�;�.X�!C?�o���4�تkF��k�[��T^���L�:z�Ro���=��k��1�?�/}��|J�{aPg�}�s��N�`xt߭�Fj���݀��n����� �ֺJ�����Y��wK�}�$�h���1�	����He�\���⇻�hm��=E���$�YD��f��cqp�`{g��@}�,@������{C������nTς3ʀ���,���M�$�I����N�ª�_�NVc���g2:{pړ����4�O,!������]7�ڬ?͸�t�>���\n{n��˼�߄P+�جhk��>-��ްT5�J��V#���^wf������N�{"��}Y%�Ry�m����X��ߖe"mݫ�gJ R����*���4�[�dۡH�|<`D�`Gg���#�t-�h��8�
�%Z�y~>O������+8��&d���=����x'v�����:����^ډm��Ԥ��N/����{۳v}��b�x\����m���6�z���I���l����>�ϫsgR�M�WB��'�oN����ٗ[E�����zv��/���	zZVv�t�Ğ��u�"p�W�5��3r�3X�]����;��JP�\f��
��wtq+7��a˃܏-(;��Ro>�gW��T���p⃎~�ǁ��r����h-{qR��a;��gYǌ�,�i���:;�q��d�(�z�_�L�p������h=�����y�e�f�M�;�xhgE�ʅ��y-
N��_?p4��I3��$fl�au8��:$S��^�VW�����`�*� �..�߹]���ƹE~��:�^�B���F�F��w]CBw�z�F��R����ޫ�-��L��y�1��]����rW�{h�!�m�ro�GT)�����18{N��'��7%$=e��;���Ğ�=ae��J���R,��iWhջ�\'0�,��,N<.�y�T�jR���(�S[�Ǉ����~�~�Ӗ�lɏ�ƽ�?-��^pC%}��,Ӳ�W�o�J�Pz��J�w��ڐ�q�Vn��4�Im�8���*�Y��ӏ���(LS��F�o��8���޳�};$z~�!U����սX/�pV��c9%�]"aʶ����wt��I�����B�n�W��-�~ӱ�g�j�yG|�z��S�f� ��o��Cv*Pp�R��[�3j�	�@����7�p���Vk<�b�����t�6�B�����3�5�m�ӛ`���}^�p�>��#9V$(��</>բ�kR�p����wU��=�_k�.������+��7��rL�!������������p��Ó��:�(�[W��8�m�fL�v�Cod�p�yND�:�Z��g���6�4���4��%Ó��\���Pd-�	6�;�v��y׸+R9��B��q$_we+��u�S�R[���GG��3���L��fW��'w�[]�1cu2��:��j�pL�;��zvv����g�.7�ٷ�2���鶌�P�T=����y@����d�[x�8GV�cT���+.m�CW�y��1�c��V�T��m�?<�G��f����;��� �S0�^�,��t<m_�A{[!@Q^�!D.�&��5�B���+9��WU�T����N�=J��!��w%Q#DPg�+�^�ei�3|D��bp�3��X���$��]�p�����K�xv�Om�$���v��o�}ھ��r^���Y��}�j�v7����ٕ�UG�p���q^[����_8�c��[��(���jͲy�W�g`ܑ[FE��/��ͭ��	�����W�JE����]׈�~ ����ɼ/�n����&�)�fkZ]5�]M]�����a|�E��\(��)���}i�M�N-Ǐz����(�L텬�4�y���)LS�����/h�cR>Iԥ;�^����*��y�g��f�`��s^^�p��
q}��f��u��y���8��J��:��2HU��@N�(Ndיrf�ӼM�<���`k������7�9Uj�:"]��X؝��<�e�F��f��, ��<�n�R�1�wZ���s�^�[�I\3�Ӆ�"�s�?dԯy��7B����9d�smv�N�$��2����,��zA�f�{GGPS^�v/��s�U�>�INxq���y�o1�p^��X{�
S��槍��������{?^yT�߽r3�~��޳�$v*���O�����X�F�w���d�l�"�����d�찟ADo]H�8L	]��ރ���cd�]�9��(�&{�K�mdUd���y��f�u޹����2��{�Y�-�E��u�gz�͸q>�T2�cO��Z��Cʫ����m;9s	�c�ܹ��1@?�7���w�3`���ʀ���*��F�+N�g@=�f��"�h��`��{w�k����r��]�n췸�j�z錋������}J둗Q-�L]Ն�ܰ#���G�6���e��]L�e�+���
������5���Wֽ��p��j��q�#]�܂pF#{��ꚭ]C��N�D���E�ӥ��=2$��n��U�F\*r�ܫݧ��[U]�=��F\����3>�3�CW�'�PI��͈����n߂�(ߵ��<�f����#���,/v�g�2s��u�[��[���)��8P"��N�����ύ��PkԔw����e����u���x�E����&��H.�{����P#�-������LT�y4�]�`|k~dAs���/��?u��ҹՐL�8 tB�M)�<�j�JԔUf�&Y�l�����<��k��84�N�/�B�uf��l�`�j'���|�u�y&��K��C�kvFin>�r��$��'EI�Nvkࡱo�jf����|�������RO!K�散��>�xޖ����|Ǩ?�ǵ����o�>�V�^f�3\Lu����f���

�\,b�E�}`zg�D]��
}�������m➏���]Z���)�7x�>l��j�5��+��{>U�B��,���L�btv��!���B_��3��[ ꌋwS�<E(>���Z8�5�+��j�ȕ��S�c}�uQW�V��
�����W�s��-��}��%�i�D�V}�'�Ȗ�3��j2>>�j{N��V��T O�:t��L��$��	�5˯e�j��^���Yځ������ b���H�z�n��*�����kvJۦ�k���4;��\�`/�}^O`Kj��띶: ��D<��������V
��-FO�r5�Ҝh�� ��#}N(ξ�@��vj����-0,<�{,<�/��ߩS���`f���_;�ߒN�x�^;�5;�_u�G3NMv���=�;J8��`��V�����=��B�P�+��ɨj?*�k�o�AC�﹡f��>&=�=(�?fM��1�cB�y;S�W8o��Yn
�c�vƒ����:5��(RҲ����"�����5i��a������X�p��mqRϝ�O3�Cw��:�^{s,��vv�#7�%�{0��0���f�{q�ӡ��j��'-�m�F�4�G���S�i2��W^{|؁�����I*`�l����K�%+��K�XEG�77)�*�͵ݓ��N�$K�m_`�I���g.�e�4�L�1��iY#=Y]{Jn��F��w�N�=�=���"r�-ɾ��о�����n���}�S���ύ��HK��pict�5�9KQr���&���0pqz�=#J�@��{k�>���E� ۙbUwX��&_'ȋ�!E�4U{�<w�H�%D�qhJ��5%`_��@ǝ�~Y�H�[�ڢ�^H^��7Gn��2�E���`���Iw�ϓ�0Bc�e�t�G_Ϭ�S����ׂ:�9�"ȹ2Bq&w`HRі�o�5�O��T�wf���J�w�o��o��N;�F��~F��*��>r6(�1R�:yc4�9,-�f�צ�436���fC�u�����Ë1g�7\��4��:���Ϙ�?	U�5�=k���]9p��mX|k0��'�o�5z�KC���;A!�u��B0`��yN���/J�ݺ��Ro!N�a���mk�5=xs.��&�OOz�%%�����H����y~W����ݮC�ߏ�^ݙ��F�53fQ��r�f	�����d�Bν+Ǝ)����#�d�T������aj�[���c��c���P����;:	5��F����m�VAÙ�P��]��d.m�芤���k��\�!�������C;kMv��W�(t/VG�
m'u�X����c�AT(]�
����(x��yS�r	�(��w8����t��w�໒�R~U��Lg��a��!��o�A��G��3/=�pAa*?��:"rf,��ne@��ޛ���u��"%��qv�}�ț�{���x4���N�8��T0V>�D��U�������W~@}������;H�~Eai�V��řQ��<��ys�g2��"�̸~ژ�����U3�0��b_^f��΄�˳\�]���9�k�n�y�9.:�3(��kc;���x��Yk�=}��p�w��<)JqD!�f����v3:��@���DE��j�K�W����Z�����6��c��1��cŊ��˯P1���2!�U8��kn�;�hE�U�(��,�9��iUh�sW<�\5O�����WmB��(��j�":�.&�W�V6X��(w�V]��ϸ�+)o2��S�ܔgϛ�	��S�_1�iҳ
���s�%�J�c�H/zNt�G��-��^�l,�݋�_M�s��hk9P ��9rt�Ӕ�����[�w��3�_A^,���'�=�2��<8�A;|&T�6Ü}ƨ
/��Ęz����Jx%��yf�X��9�VT�[��~�-�.����������+�U7[�����s�fx��1�(>Ge�0�
>v�]Z"������s�.��Ű\���F�T�Ce�x��}~V��o�����`,T�
=�e'�^�ѥp�gw>a�����e7�5�8���.�n��y���3�;�eV)��Փ�q%�A����/Qm�e	���	aAr`:D+&���w8ug\V�c��gh���#ȹ�J烤r�h�ip1�����elvx��9����7�(e]Kx�{�M�4��Uf�c�%�y�t�9_�&o���MX�`�WQY�N��%A]��9F1�r9_(���;�Er���ǖ27���=�O���)�hW��2'�w�W�/]:�_	�hv3�,@���멎��P���]�32�x�υ�ƣo�J��q�[����R�p6I�,g2��V틑UF�ʿ�q֑��:�[�'~�l��s��yО`�n�EdQ�FU��ܴ�ջ��A��U_:�h>W�Zn��Gd>��(_��Y�Dcyr��վj��Ԙ�cj1�r�1=3�8Ρ(yS�.�fθ}0��80K�����co��V�dY��﮽�+v#ü4��bkzP�;U@�|e={B3�"S�{�cG>�y~�S�O��%q��^�j���čQsZgK�Rlnz�N��������@MO��K,`�O� +ð���*�k��q��x��#q9�Ej�p���Ϲ���:(�������(�W!�%l��e����-��TT�k���y\��Y�pÂj�:qw@U�a�;��ӊjZ��;.�����r��x�8��sRSl]���=�� �"��U�:����]�i�YG��{G�zD�}�<���x�ʕ��c�z[�1ĕ�-Cԍ����nV�Bl�����澏����Ò���װ�}T�[ʣ�ў���n>b�(z�w!������If���@�޸���;�+=�K�V��o���׌<�}����n�SW�9X��>r��e}^�2�~���{*f�O�*lU�%��
��N�N��<����y�>jx�7�����Ҫ�����-	D5���+<{�v���kz3�i��ݕ���_���^��_�t��S��L�Y�6{��D��F���ړG��Uj�|*�틵�F�ڏ��:�v�'�g5����z�:8V9�1�LGH�^Ƀ��s�L�a|=���7�}��`]�͑o�0g�����ŏwS����>S`��"�����[���}���ce4n��0�`[�Ͻ*�Blg��SR��5֝	ܡ��R.*�b6����F�[��7���_�������)\sA�D}�ǟ�@�*nn���v��ę�uW]Z���Y�D�#ѽ�$��<Þ��^���lL@��c¼v}e�d��猪`��« �Q�#�����5�J��d�W-�_����]��
�N7!JQ��=��j&�//U
�K�m6�:U���ÛF����:��wdǬ�2���3_Lw��[��Rb�@���%;��l=�gTт�׼&kAmw��{ɾ���1�`��گ��C>�s�c�5�]6/�W�6
���:~w�d���;j���O�ب��Uo��:�_LTֲK���T_~���'�6�^�s�=^�-muB����@�P�<��=���P�5>'8E囶�ƻ���p�����߁x{���o�;�ɪ`ܮ�*zb։=|�X���.��s�[��Y�[^��M
��1?��CՐ&��|+�cUM|�z�E�E��q�"�>�P*�̋7���ɋ��D;#C1�G����$�p�lK8���1��^���ed̃�]�&-x�k�>ߺBcvc��n1B s��f����spo�n�j���N㘉��h�J�6nq[���!+'�%����r{���b��y�T�Q�&vcΝ�O�G5�Q��wrdF��g��]�� ���k�3��w�vK���z��4n���muF<�GAD��y~Bt�=�hm\Z��M���*�3��T`M�w\�1s��rxa��Li�V���&�*=T

j$mSzT�L�{�(�*g��}���K�}�/_|��Y�K�{4"�8����)���C�ۥ�T��*�G.5�6�^z�Z�I�t�����a־n�I�ӵz0�}N��9���&J�=��+蕋��˿�Ӣ��F���ĥ��=*�)���>LCL���_J�)1�&�gLQ��?,������hC˸w��E�;Vf��-ӳn����%�)t��ʫ���X�����f<���ۆr���q�v�hwK!��ŗN�*^�9�٨�Vu��j�w�8�D�U�iJu��v�GZF�Ȣ�!r�#Z�PQ�{�8L�*��Q�l�7�����:��8)�[�rU�8���v�mL����̮����Ăݘ����(��u���6��[hr��,�]c~Mc'������[y��ხ��x�k��g0A�<�?9V;��2��6Kw��/֌��{��Z���d�p�sK�v�i�qT�os��rD �h�X&fMY� 1��U�+C��[i�Ԉ]�Jh>(�Z����r��ڬb�6y5�٪Y�z1�>&��i>'rn��v�,�#��P'm�O�q�8^�Vn�>Ѳv�u�L:�}|[��Ū�s�Į�������.9zvi'�@�����Ӯ]��S;hn�J����f�K�dk�J�#�l�i�v��oy�E^|�&�/�!c�t�c�]\5^�v�r�5z�t_i�O[��S(p�R�v��7��鎶��+�<��ɵBԣm�U$�}���~Zk3]r��
c�vVǇO�/�DQ(�k��7�]�q����wu%iP��0T�kh,��brͫ0��̛wJ��H��Q����1[Z��P]��4g=4Ŷ
j:���=\h\��wz��:�kC󻶕���3R�wc¦���&���I����8����KE.@�����h77��f�����(7\�$g�c"P-A�A�`���CB�K�Л֞�Ng��a�a{�!��ç�Ҟ�)nԶ��1�e�ZEQGJ��D�v�+��(��o%9`���-.~v�}�F*2U��6߰���a�*�TQ�$Wf�K-A(�B+ ����D�{?LW˶�l�^��D_Os\��d�BO�P�[|��S��w`���{�v�,|�x�F��rIC��Íڨ1V�Lu���`̡7ei�9�7;��y�������� c"c�2�>��|�mA�|���X�X&��Yt4L[�E���R�w6�T���!n���o4��w��Z��1�j'(78\�X�Y˹�4�:m)R� ���I�(��\��� �\�81���W4�@;kq��kY-U��0���]�q����ۭ�&'�aP4qͳY�E���wiݽ}�j��*�1�{�ժηW~s���6�c�
	����B���Y{���������0�ím���LO�����Q��m��v&�"eOP>;/�.�3m��M��NwY\��j��v[z,m��]4���K���H�RX��G	�nUm;��Ɋ���O�"�?�4\��%݋��K��L���ƨ3��aB��v[�0]�<�����#���#5�f�D%fu<�B�!�z�K���ZF��M��bw�һT�@���67�6�'�/��|> bݍ����lE,����C�K�S��ƛ�;
U�����`��^Mt��W�Ly�ˠ�Dh�m���^,3y9Xʁ斉x��8�o�-[�^�ř����N5�t���z��13�'�1;WS�#N�Ãj�	x�E��v�f���XVV?��k~�C<>��:Q����@K̍�+F�H0����o
��<|�W|�U����'e���ɻIx���vM��2�U��6qW��_%b�3�s���M���o�j�󘒧k�ۏv� ��p򺨬S�D���lq'���+"\Q��f��ѺN��3�LB�5q\iUw��cw��"q��/M{:&�z������=5JBl8s�>p��q�ݓ�[ޑ��	��u�-[�d�.��#���`w�ϼ���ž�ql'����f��F�;:��2�J��x0������0{1zŞ��H�2 �ݧ���Fw��<�/�	���6��>�!_R�.�5�{s�o2 �vz��Udy#e%�Z�Z;���X�m��W�k����e�dq$nB�5$3��N#��>�;�*cޭ��K����u5� �y�a�ݦ�np����]�:0��=
�S�^v"�I��&jȜ����-�ߟ��z��=�c��8>�N��5��kI�BV=��u��Nf({���ZSFP��$�d�*��U��Vc�㭸
����N�W)VY�E_Y�}o�*���"1�d7s��x���}9j���5�sV��������2�9���,���8�s����u���[�"|*�^G��\����S��%%�;mD��q�sk�]ۘ6�����Ўe~������۔��4�|w��|#�/�b:��*�1�����r_y�{�'^�/��mxm���{���@[���<� �G�����r\�47�3<�&�Q�W4����3ى/�Bʹ($;�]�=7��3:Hg�.fi'��M}z��w9������l1-�jm�ִ�G���]{&�2CW.�z�=��@[M<ǣ��@?��p��Y���l>�Ee+w:.aOVa���G?�����=p(Li35G�#�W�jx�aY��%�=��e�`�{��Uk��ڃ'��_ElԷC�#�oW7�c�ZrA~ى�!�}r=9r��gm�}�'�Х����;����b�2*�uI3n0ΓY���:�v�V!����ע����{�:p���H��=�jD�3]=�0\;�hdw���U�����o	$�7�Oc�+LL^=&*�[���.�k��T+";�'5qL��2����tif-W��>s����1f���ϧ���	�j�!��is"�ћ��O��'v�3x!s���E�iZ�,VJ}�JN�V^XC���1�m:����Rى��y��9�7��n��HS�_���#�W��i�wpr�� ���r�n1����$���Ip�z6.M��Q'9$�Z�ʗخ.�L��j���㹔/�\y���j��kJU��]� �"Q�b��~������hx�f�ą�C����<W��R
[�L�Fꤠ�]�7�$<s�U@�����Ej�x8+�����'-�̤R�>X=���H?�`���7��������l�$f	�R��ogy<X��O1V%:��Xo�*u�F��)�-�K��3���7��Kc>��籃�j��Ӿ�.��A-^�ݴ�B�f�(�{���i���*��e|����݋75���a1�m�<Mё&4ڶH���٢�?`��\z&�s��������d�*y�~���Yֺ���}����G��g���/.L�[�����"���!1�K�g�d��?,�~��]Q{�*�뉯�|��upG�ݵ�A�c��?�l�q��BW՗x�#���ȕ�}��}NEGT�W��=�J����)�]I���DĬZv����%��,��3�)I	�#�g[0�gMu�ֳ�����&.�M�'F�b�kf�DE%���˙����(Qv�ű���:}͖o�쥞��*4����_�]ޚ�A�������c"�f`�ܫV!�� o������.��ͺ|�ٷ�Ǒ�Aн�bm�1�p��h��ѡ�C���.����}
�6��잉�i��*+�= ݪT���5�&H&p����.�����A�C�-c��:C�7&w�L�Zv�����*���O{�
���51�Cٗn=g"����3��8F��ѐ��"w5Þ)�9[�i��3kG����F�.<�v�����b<%I��}��c0��{�Q��^y����ڎ���N�C⼼r�Ф��n���L�:�E��<���n��4��gI�\��;i��"EjL򀱰G�:��Z�j��s�w���L�^z��#5���ֵ:6�YH��^��.�u�z�╣�̽Y��Bx �S�=t>r|De�Z�P�;~*wϧ/�}6"�	�P�h�>kM�x��;����_*B�S;:�e�Y~�/�#\��O�Z��,�s��f�'`�3��LT��Ō8#}^��b~�`�h����������R�t<g��K�|ʈ�&���B��Lt$:�\��ڿ�����{�T�A�g����Aѓ�Ǥ�j�iK>۸b�b��d�6��17s�F��R�U�v���PB#TExz�$�	��!����X�T&|��5�p������}P<c���5>ޜ��u�ٕ�spWƍ+�G�ke�Xfu�t<����WM��YF+X���|w�J�c|ӳ��e�F��"3�s[�"���#[kh�W[�&�U��+�q��[׸Ds���l�AIY#�:eѹ��Ǚ�&�I��Ww��X��t���"�����y����U�iAw�΄�}��p��v��K�iJ�V�A��A-��6u+�0s�R/�fB���5M�z���ܳD�	U�K��ԕG��}�}e+�:d�C�Y(�h;�:H�x_Fo����Sd��m�P��G�W��h^_�v{M�`��f��O(ߋ̥O��b������������#քm4�[�s��z���M��r]����x���3�#ܡev���g��W�"�&��p;�[�lN�v��#x0p�^��vkj]��~��/�������a1J�:�>�v�P�uȬ�Z�"�R�͚�|(O{�Sn�Fy�^��7�9^�=��	���/n���6���tW9��ξ2;5�#q�[,�l�l�}7GӐ��Ģ�]�5��]3C���6�ޕ&��1y�8��ܿE	.��*>������b�F�:YX�򖏙jd�ּ�L��-�b�#B;4���B��̳���cD1��z�u�cw�|꼸(��l�=ۙSҵh����&}��U'�Rb�y��K������Sq�:�Ω� �j���C������Ͳ"9B7V�ծ��w�am}�"Lzb���J�%�#�;;�B���Y̔��R'�V�ᖢ���i����n܌`Œ�}O9���Y7��ʸh�T/���Y� HS[�J�:s����.$qofoR�:�(V���^��ٜ�����{jWO���p��*��s�r}s�ܷ�/��ݬ�9{ԯ���=8y��d<������uM�LU =�2)�܌����%�7�qf�7k4x��;�ԥվ��Nl:�n�wӗ�tՏ^v\��]��5SX򷂙�ea�C�N�
��wz�����$���h,�?eBȱԔd	�=#�4d�X�zG)�7&4mCQ��:٫we���({��IXk<V���3�ޱ��� ݺ8^_��3�"�>���>�Ժ����k�ܳ�>���<e_H����v�M�)0կgw��5�8H��у2���"���j#غ}Eh^�n/=9g^ ������&؊���m�*FV}"�b9��v�}3p�����T��ɳ��s���W��Z�4���d���9��̧�9�WF�w;1�W�tN�P��f���7�}���LT����Q��VOz��頱��{�;+����@�\F!Խ��.#.hJ^'�r�����7Ѥ��5H`�3�=%f�u@ʴ<s����jp�H땽o{�K=Zk��A��i��<Y~;w���#2b+��0%�4�b�V��=j�H�g�<�'\�>e��ة_��c�reŃٍ[��^�����IsU�Ru�n�)�2�`vo���]��������}��<P��5���`�e��q��F֗�;�ko�ꛇ
��-�lk['m2B�}�#���f.hew�y��#F��Y5��7�cR�d\�!�ǜǖX��9�x��;g`G�iO��ч�>mG�����7�}�F�o�ڵz���L=Y����\��E-�ڙ��e�֙��Z!zxq��7[P���|�|��f�Q������4vj��K�Z:W'ˬ�[�Uc�َ�S�t��y�Ca=@��r��	v��m�ҫrc����G�¶�03��ؼh��m}^�l1^и��#��F�����鯌<�O�黩;�{cN�g�KM��H�1Tm�.�,ط��L���oQ�Y�B�}C6)�w8^X0��-��yQ�%�C��]�+g�z��`Eǔyf�#�t���
�y����C#�-�7J�L��������R&���nغ	]��sE´c����;�S���o�핳��y^���kBWP�{K��[��uoH����T'՚#�5��֪͊���5�j|:ODm�R�Vw�P���&&��ߥ6��[3��ơ�}��yȫ��~x�k�U�M���ƆGEX��ՙ�"��k�T�piM]k�!l/NA��Ғy��hN9p��Bj7�cķvP��;}�jOr�Z�GT�K������	\�Ǿ�7����1��H��_��&m�e�U�{�=]c�;���>h�v�7�l�Y�I�[��9mF��^��0\��q�Q�k�Z��j���y{��NSSEG�����)n��ٍf�C����m�7֟,�Ҵu� ˲�:n�mpZ�ۭLj� �|�S
w���NDm�;u� 7c2�_��}X�;� ��Ȧj��F1�;bEf��9�S>,��������xW��Y+�d�Du�lb�]�S�!۸	n��/7&�1��~'Ͼ�p����Y��TZ�^������\�Ԡ��[j�~��p"Y��شs����.��F��Vծ]Ez�(�qK��|�fe�P�戳�e�^cTi���y����s�B��{+���r�F�����usN�OUd�ψ�u��D_ ��H�NdT<t.�^�ſ'�5DɁ$���[�M�:��b�[�X+��]��PY�â�	�AY�Y31༊���pۮ+B�}�����V�+�{��q:���?��\�e}�q����3C����Q����"���.;"���B�^w��+;aOÖ軺�*���fyc�0��
0j��
���+�
`��W���#ã�.׃ܿ;E˴/海��.��(�yւ�>�]���uR��2���b�4�'&ol���;�k�;dX%���u�GLEd��k��F��6��:�����*'ܡ�2���4�����\8�Db7\1f��+��i��+/#⩥��j��{ǟV ��D�\�u���2�ܧi�Vqj\���Ėy���ɲ^Yl,���;CC�<�u�5���Ի��E���=LnL<�zL������p�bg���9.C���0�t�[�,�F.�%q��&���ᡷS�9(Gߨv�3���9�ħ 9Y6�3�;ݗUMĿ�󜛔�*�g۞�YG�� |-[E�χ�{3׳��-�E#2������F`Xm�<�{��s���iV\g��)�:����yB��N9T#;�=�(x��լӾ�xA"���} ������у�wss{Rej��9�cK�Q�j�K�.;bc�f�m�Լ�#/��J�Ҕ�b:O�m�1�s�%�e���rn��}�{]ǅD��(�������˸"}�Wi-j�@�u��,
��I���UМ�����}>_Xml	�Q�3�ݠף�!�m��[�.K7Dޭ�꟎��t��u��Z:j�u��}I-�ae���T	�(��y��t�:3]5jm�/4V��S}��sw�vWק�42qjW�y�&�"W͋���+����&1���}b��5~&��|��|an.���ٜ��CvqЙS�&w�Y���LQ��hL9��)q�w哵
�d����b�]<E �o�)�"�-�E*��w����R�D��!��>�m�����'�Ҝ�5m7l�Y���)?M������J�坤8'߻��&�WB&�Q��ڒ�>�Pz3;���E`�[��؊���ݳ"Y��ɵ���y���-����ɷ�	��q��Jv�f8�-Ҭ�N��~ͥ|23���u5�~�X�
��7��ׂq�"������O#b_�q�����"b��x������] /XBR��]�ž�_0���<&�FRS�v:�yqc�pT��^�h�$�9S��e
\n����=�p����k:SS+T>4�P��y0�����ǽ�s�*���U�N���B�
e&�7SQ~�������G�,���	]�ɍ���-��S�g�vs����>�?����3l߽ܫ%�x5b�-�)�{�m�3��W�3לcoO�Ij����k��u�3��YY7˵� }��e���dV������oL G��sO��tXe_.V@_LjC]�d�9��Y�������F��l�&�Տq�����%�Pp���a3Yc��{��1�/���e���k�y�UW\�.]_�����ɤ{�i#���Wl�u�/h���n�����M�Y|�c��-2.�����\�M���Y"��IΑUH�w�$O�[�^}�\+� �{��|w�^�3��'�q��������	��0�
��ӟsX��﬎�;L6"%۫���.�yIbu �^"���a�e)Z#�+�U��aߪ�M�8�aN8l���������{MYPWR�$���҂��#j���3�
[�J�wJ�nn�p��װ+��j�B0T'@�����R���۔)�W���-v��qu6X��k�����;���x�j9t)����?73GD�5t���J��V��`B��t�hC5���#�����iy�K� |���'�
��6a5vs]�<]�i4�]�5�x`�v�3h+c8�GK���tT�Q��������۝�b�&���ϯ�H��@���'��u���`�ߝ*|��R���g�]��s�I!Ԅ�;M�u���In����-�	&�t']v��C=x���Hi�@���VO� �r��y����Z��^$�z���$��{Y�T�Z��0�ҽ�{�Hy+�[�I�~d��y��������t6��Y���s-Me�봮��u	 {���>��6��@�JU�GP0�2�1G�]��w��1�s�����Up�n+ԭ
���AUb�T>���ץl�ˡ֢��ﱻ��et�5�ϣku��o1�(E�US ��� Ҁ��حv^��{;�Q�6�h���eZ�h���uP�W)��涟 ��q��j!A�NY���^�f� u!�3��O�Hu�%��v۹������\EXLb�P��Έ�0��I!�&�}���w�`A׮g~p���=u�1_x�o�XkZ�a���i }�0��/n���g��~�T�Ƥ��.c�6�����ʟn��1��fk�;�ׯ5/Ym�h����S�q��fOe��mN�n$6�38�Y�/��{����٣����4��^�)y �z�'ʛg��!Xu�ٟ7
�웡�v��2���7� +� ���z����ًw�'ES�y�om�ᢩ n���Dأ.����~�ֆ3�~VxT�9����6���V������S�َ����{��c$'>���.��S�|�!�Pt*dô2�����]L�ut:�!`=^�vX� b7Cat��q7�gyx�S�z�n�玟���]k�I!D�.v��u��_�`CH��=���j�m��k�f���]�Wt�PP���1��9�ͬY'h�w�s�<0��xR�qm�ݜ�PI���H
�D�ǽlB.�B�[��s50*�y9.X�D1��5nݙ��R��z�}�46f�x�)�¶���w�M�7���pa�V�,M�I��Cb$�����O1�c�d�/����`��̝\P6��צ��-�KZ�YV����c�P�i�pn��8���up��a��Ս�
������8aF�*7�!�zM�dۮ6����Aݞ=����@��E��Ep(��gl�"]�B���p���]�]\"�eR�*]������	d�鿚����M]�ܸ����X�=�;�U��I%v�q�:�Ru��q/H)��j��_+�V�q���իD��ϭ���j�b��X.�i�s|[��Qf�K<���ڍ���x&sj����V�NrT��u
l�c8r��/.�R܎I�N,�4����̝gUm��ï���R]q���B� ,٠ �]}C7���bM��}%R������j�/��,��t����B�,���)��W~��Zb�;NI�+kc��_GAT�x�vp��/$=�,Wc՚9��=ѴՕl����S��T��{F���b��=6�mh˩�l�C�a�Gv��]�)���4�n���׵�:��.�cD:3�ӈX��b�\�96d��׿| ���&n�{w'2yp~ב��n��3	��H�i���wY98���s�a��&9_e��uN�l�z�F3���fT���w	�Ǜ\�v�L�h57bEˡ��~�G7Eԃ�x���Sٶ=��b��4l�������vp����3��	*�1�3j��}N�O �������2����)�K����_�C�Tq��MMu%ێ�+˰D�S�_��)Z����o��Wx��9���ɯ.����\��	t��3_W��D���[��S���Lw�.�+͝�H+�]=����M��o)�,o5j�ׇ�#�/~������8�_����"ݓ*�3�E��yY&����X��EOs���Ƅ6�H/r��P����d�y�)_G��//����v������
6T��a�뤦b�b��i�>6�?@�"��<m`y_zn�&���M֤���8��`��6����=���>.���)�&�Qg}.|��0�����O̅6D�ek�R:1��0�	��8�^����+�ŅW�9>�)���g�a��L!��EY�u:bШ��5;�h�sZY�O��<#��	^�b!��K#����y��>=��ŵ�ZhVr��l��LR�Z�F�闣�α�/�|��@$+ہ7(��U/3��S�pmkW���:֪0N4�	v��L���8��{�0TLf&`��[�Fi����Y� Y�+x'XGf�wF#Z+�	�j=�JX��ܧr����^�%(��wf
��E�S�PW�V�}�6�8iޜ�5��6�Z9��?10�C�R�W�<ԓ7Up6��xk��ro��z���e����}�eg-ta0��!��)�[m�"�#�j��/,!�C���>�f���qU���L��^$�k�n�s�2���m͙����r�g��^�=�ٺ�d�\%"�^q�s]Ӯ���G���h�B��ɍ����o�|�S���ޝ��׼'��@#&r��={����kxL���p)F�L;C��BؓV!���6D�K��TY^~Yx����P'w�l�0l@��qWY�X�3��Z��B�wڵ?��sW;.�������S����$H��*Q��g��q�Bk�ϝ_ְ*�=ߟ�6��*� ��Dg���g������!�e�/��(Z�QB�k���T�$>���fW���Q���sq�Lܭ��J޿�{!+^�[���e^��8�f_�DJ���>?/��Wܦ�� __�_���:WC�_;s �L2-:+3�p�^;�{"��!?%F'hu�z��iŭ[[�C`����sslͼ?t�}F�F̹Q8'�7�>z4Z��YE�E�z~�̣�P2g�i��Xɹ�J����\!�n�W�Z���Qw[�{J"EK��e�֖��q���5:P�aW}�ko[|6�;;�X��w�QXV�ٓf>ʇ�u��.����6ŧI<����[���MC����jucv�ƾ� j�J\���`o1θ7'[�}�<L����
�jX��r]�y��tp�'�N���w�����ҙ���8 =�\���1�s"owy؅�oqz��5�����a�D������5q~�����$m�tlf��Ƽ��H�X:�FV���n]�	�`����+%�
�}O�	h�Tơ�Ë����T4m�S4��l�G����nb��{����BS#3��4�U����o���}͙�_��k��p�d�]^��׫��H���k-	��o5ڴ=�M�{`+�(�w6'�f�d����]��s}�"=�x�)ޛ���Y�)����"����\��C����J�`z�c��|�����t0��Wv>�_��8�9t��ۖ�b=��r1V��������Y���q�c�Z�r�g��!�˿��f�t������΄���I�^��;�_����{�'$Z���qӨ�c����'<� ��ɓ�t)ގ��*�8R�5���.FD�#Kd�;@�Moe�]L�F����?k�Fhޫu�GG������|�P���ÞҺ|1�jïyz�Ji�/6%�s�rvשּ�D��8 �{U�2�U��׈>���� ��ަ�_8AuG�q�yQ����ڄ5��U��FDk2�s�)��0���m��R�I��.ې�dغ7t��rq���J�+'ooV��r>�F�xu�����g)�4�u���gb��;�6���`��K4Zs��ֻ}���K��Du��P��f��ע���3�]���N�Ȕ���9R������7��랊&'q��e���O5t�����1ƪF�-�4�r2��-.�W%���u�,n,��={"Gz��]Mr��^�-���/�*v��������yG�z�直uEY�2!g�����c:�Yr:N���Af��WAjn��=���RR���z��h��7N&W������j����L�;���1(@��'��8��2c���������u�KQ��z�=
���ϫ��l��A�p�����O��R�>��<��f��^�H�NR��
�4ػ�$�oFY�-z5����WV]w�7��T0_ו2��[�}7�ݓN--�K=��s��|���S�^�0�#��xv�Ғ6
B���Oֱ��8 EOP>J;��µ~��E�L�<Ы£�e�{(4+;$�x+����-�kA{Y3���E�f�#n�t7�{��Fʎw���'��r8�C��ǲ�l]L���`< �h�7~U�f2�s��D��a�j�|Ŧ���9�w����֭�fY�{�U��,,��|���]t��-^P�jL�ˋ��W��ک4m��huW�j�Y�θȲ��J������d���ثLh1�m��җ&���U�� �k0b�xǔ�뭒7Y]�>���t="���q!����Ɂ�㬒p~$I���ʽ+�w�o��Ӿ�П������ݗܠ�'x��0ߠa4"���T�H�u@�=˄NYPȈ��2��y�P�G�廕���c*l�
֏J^��]��!/T�1{��B���-ذׁ��M�����s��|vj�ػL� \�p�=�\;95�p]!�{��)N���3�RB۞�^T��}��F&<�������� U��'��ߝ>�8�ӑ�i�<���I�w>�_��4�����5y���K�_��ڬW��P[��Qv��^<�����-�,N�n�3˦nЋ9�2Ǌ��㙇`��
�`���Ƌ����_w��Q�X|((Z�t��ewy����4/�QW	��2�s���':�,��fh�3�R6z�U�lh;Є��dԯK��<<^!@�U;��7颯�F���~�8]v/\�^�b`�(��
��W�v�&8���ܫg��`<&w�'�q:R�?��z���%s懁����<xO+��
�V`P�~g�t���vt�
{ɑ]�.!ޡ^�oξ�]����~oE�g�J�ԉzq�Qt���y\�Bn9>�5s��B�3"�a�X\�i��k�(Q=ah�@��SY�N4DԺٝ��o�M��u:�m��Z�igK�e��֮�J䕽�3zݐTν�ĥw��X�]7x�v۴�gwJ%!�C�'(9;�����d��w��Kڍ�>����RB쏛#���ߚ����}ף�q�g�_��y����dՆiY�cEj�1�E�1�>�l���o��M"-��AwQ,TY��)ܹ���!1���&n/���'S�����~/5b���Eiu��(j�=g��:~W��ld�>�݊T�z�y�l�=�J���?,%�u�#<���8��D{~*�w���_/�6�;�-v %K'l9�oN�A��y��{P�: �:@�;OI*�]�q����C�3VuU!��?}q���Ȭ��gi��:ܡ��W��n��u}g�\D�<�Vh#�������N̨o�"��Ù�'YB��+'U<\���H�T61�,�KMHR_�<�^���̛Z��s�\�����q��F+'%���M-��($��X��W]L�$�Ʋ]�~����~�]����^:�ڴ$m���>U����2LK�ب�܅�n5��)
�U:���zg0����}>�&s_8`\]�e�s�C,v�b�WF=4 "�C=���;�w����'f����@�@�K�S~ɨ�ҍG���م���Lӣ����I1oS̭�bM�j�t�B���H&͜&'Yf�*Ǔ�-�	�ɵ�ȣCrh��vf.N�J&�]��R9j4��LM�Ɂ��u�ל�jv�鎺�!')]��N���f9N�φ >�j��<���� 1�@bǠ]��q�5�I����+�S؈�;�W������_�3��N��VJ$y�t�gX&���(f��럣�u7��7�	9Z��BZ���ˣ��[�r/6[U({g��������.�燵5�`�+����	�{��l�'j��ׄ4g��C�^�QT�\�R���=Ax�g���]�_�=�*u�3'���>үč����rY���l��}��5JDR����{�.dG�1���c��*ʩ3�J�A���<� Eɨ��{�����_5��3BKΏ��:m����=�p�����aIz��y�9�u��g�(�gcq ���X��$����9_��s_�+7}�����S!)�u9���lԤ!Ȕi�D���1gc*P��zbrǼ^n&%��,U�;�9R����������vx3�`Uy2nw4��B)�[�F�6(o�̴}u��]T�<�"���� �b憽�8t�ﮠ�I;��5��x�>���ț�x��0���Z�uM
���63#I#mnT�b4,��9�B�`t�s+��Ϋ�f�厃���9z��t�7�� j�<��\���LBl�{��.u�dr���\�+���a��m�����*���?4��C�
����y����yKiNFʍ3��eӜ�Gw�q�0����0�ġ���U����l���3ꦗ-���.ͨ5���x&p�U��0ʱ��-��U�c5�𼛩U���b����`��������1C"���_�7k����ߑ̒o�*su�(������6�	��po&/�TWO��im�:]�.r��^���QWy���vm�<^߰�u�����鹗�׆�wUuK'�}�[�~;�Sk�P���}�-S;�vg����Kmw���U��h�)tu�W��*oކ�[�l��W1�x���#|��mnQmp7p�u�_u�T:j�����f�,��].�:�<�K�U�6�w|p�9:����n ز�1Տ}rO
�
ٶ���߸:�����S��vz����c�	��q9��N�Ξ�<j��^��RS���������
��i��{;�V��5G͝�7�؉ƹ��ԅM�J\~���!#v^���Լ:p�?R�	��q}�#��Lˋc�W�ە�k�������(w�l��Ů����Y��4ڵ����0��5�kh�F�oW)��l�F`D���F�j%81�;N^�r!�e��sL�mvG(;|�u���`���+������<׬Qu}O����H�D�\�	�{N�fI�g!�
Ǻ6J�2P��a���j$�g>�:�`T�Φx��y?6�v�Y�:.M���y�Ⱥ����R�9��b8x�7�F�<�R
��&S&^�?��Rw�����b؁I:�Yt�_'N��(�5fkVY�/�=~�I�9�R;|���D1}�)QTEw=(O�����e�5�~z"��7�~����E/�ҭO�*�������4�51p�ݡ�kfdG����*�
��}�m{BBЈ�{Q�Ƶ3,��4&ܭ�j���g�ՍT/S�2�Ȯ���y�|�z�{��]����S�#.�վf= �.���]s�.,Ir_�#�	=�]���b��(ަ���`�Qً�h�3KSѡq5��y�Ķ��h_�D�Ԇ�گ"� ��X�S�������
5�51.yH�����W�����m^��Vt>c��Z�ղ�:�^����GE7�ǧ-TY��pB���W�U���6����=��t�ƶ�ovon�s6������뷵�%T;9��%�[�!�9���x�1
�f`��#f�NF��^\yA���:�m�qz!���59}3O8vW��m�`Sn�n�9�^j*��FnI�����Z�XaX3MHj�=�Ѕ�/k</����b|e̵e�®���D�!r(솸���eG�Vm���Y�)j�\�י�P��J�o*���Ӥ�d7���`�w]�3*� ��	˔�6	Ҷu����iN�e���21��)��1���Q|�����Q�Իkՙïr�O'B����)X�u��~�%��pZ����9��E��-gm1���Mg�e�� s�2u���*���g���
�C�������O,���O%�O�b���	��hWӾ�A�c> ��v)aU�`˵]n�޺��=���b�}���{���N��;#K���qYn��}q��S;�s����"z�5�g�B�&�lOH=札�j|�:^{q�7f�ʷdE�f�u+{U�Γ��_�.�B;gY�%u>�Cyy,�z����mV������`��pBd���.�Z�B�}��)`>�T n���hu�%z���G��z!�I\�MH�2+�_���=#I�=]&�ʻ��8��:�jx@��o������yn��ƻ�q ��M�����Ox�E$��^�͘:�C��Vg��&w}B���l
,�f�z��k�e6��g�կԳ�
Iq�IZ�>gn�1�*��F�NM�ݙ1E�h8�Tq�m@Ycr 8�$3]�þ=1�Cn��Df+���Y/%�ݹ�{�еگ��U�>i��>���7H�s�Q9������M엍����'YXk~�/\���bU�5��Y���`1gnly˴&���0��Hw5Q�H�q�(;��I5t�|8$:̩
$�;5��W�Z��Cy1,���zX^���\Y��^*OE>W5`��:e���d�訣ENJ�oM�#\*�c���+���@&D�-����dm!�����t���WE�ͨ;��h��X���WC%BF�v2x�V���G�	�v�)˛NʹɌ��u�};O��c����f�친M��u��}��p�6�w��ƻ�Bcv��N8v�RG�!����&�� Yy��E�ˍ;�֤;�׉�����7�dV�i��m1ae-�UpX�����M��{{רJ<B]k2چ��HC���Ѵ�&Et�������ɘ6�{��7����p!n��#�����Pݷt��l�<��~�ze��� (��F�	��;,sN��V(l�F��=�%�^�� U���ʜoZe�E�����Y��z����j����h���<yܖV4�rS�y��]Q^,���&-��wMQ��k�@uw.9|�w,���7�;�I�N�<W� {)!+��H�B���{}��!Y$�L���y���9�C\�un����� 5M�a���'n-lQ02���#��۷ջ�!{��)���zͳ��\W(��DӃYa������{�3r`�L��:4�'t��gs#���ɿz��l��s��@�U/i_&zl����=�� ���;�}�����3)F�۱�*�E
�v+�,�k?~�ؓ%�I�!�r�ڝ@q+}A��?Vq"��=J�.+�^Nӂ���jL��M1�w#����b�Lm#[r��!�	y��s�"�[r�����2�=3-ٵ��0��G�5U�]C�F����㩅�5�Jy4\V��K�-����Mwg��5�2��>��Fڭ�o�����M�9y|h�� �o6���{�����ӓ���r�f=�:t�c���-�]�~��1֚U�*���^�~T�0�)E(�_=+V���ݴ�Z��|��ա��
���{�GA�p�}/G)F�.��O�T�0vd��W]��M�3X���L�+��Xv�9u��Z��S���V����_j��YW!�xֲ;�.�D�ϡ�l�A����*�n��_�ݙ����9׀�q�{\R홙ׯ�Ùc/`�Ή�"�nM���D���y��w�y�Yn��=���\Y�t��-�4Ν+1���v�d���(d�i���^n�2�dH^�o�3Nl�Wòv�h�|��Ik��w9�s�b"�D,(.g
��r��O*�<k�j�q��yP���C݀��ɇ�T��f)���q@���]���ow�����Tes�vn�
�`����v6���#����L�ڄ�1�a0-i#[wZ�߹��- ��]��� 8�9��r��盹8�xr>�P�5�.�>3�r �8�/��f�As��z���$�4��*m���y-�ͤ�rgP�Qᙙ�ݡ���Q���i�}y����+$G��ٙ������Mҩ*;��1�#�������{´?��a|8����;d�S$����nj#�j�<���w٦_f<�g M��gB̥�!O`SN�9Y�;��ܮØ��B\j�Ml��Ry�5�rO۶}��G�ʘ���ϧ`���qv��Js����+|�ݐOf�j�:�W����X	��=1l]�"o�ф��:A��q����/Uwư�N�"�vk�0��bC�J�������U@�8z�@g��p�s�O_��c6=��>1��}�N�X�8���i=�}ᱵabzz}	@���<}�J�J�{#�(�{Ϫ�T��e'*�0�1�Ê�P�o���ޛUg��ϣ*��x<�����++v!Ɩ<;'�]-�o�¸��T{���;M�d5�Lz�f^�Ϫ����<�<K��;1���6j=pX.�����3ԝ��*<���q����k͛⯕v<q.�s>^����.,�Ӽ�Y����/�x?W|j=�*�Qw���jq!�bg�ބ�2Ǧ�4i�(z(�ك��!9UV��!ғ����*�'xḢ��b����0��Z�`�liEҬך�wdf�D(O��M��/�)��gd9j������eC=�L�\�0��5��$�qV�7#rc��R��:�ҕ'R���u?F����m��N7As�A��"��R�W4v+Rl��9]P���P�'Aݗez����۽�n�Ԡ%�K�R_y�^����v���b������/aY��YԚ�w���;�SI��'N��y�ƣ��<���ו�D�s�%�=�b��2q�3�H�V-�]�{4�X��x�;:���z��i+�O�7��xa5�0�/l�޷̈�q�z���4�_$[��|a�a�������ԙ���y,-���2�n�����kh慉��/qS��s͞v��赛Cv�<�AQ���������4���As�j��^rvk�4�,js��#r�`�L��4a�G^ֹ�K��#�=U�;w:}4��s�V6]�~���H�$:�	�wQ��!�⚞��`�{ϡ�U�(��U������Y)��N_�ˢNx��~���K�ث�t�C�ɘ����:m^�c�i���0��Nd�����pt���_�͞��c�ds�⦊�+5t����n���/�Ꞿ��^F�����r�FU�RG�k*1��{���	~Dα�'QwnȺ��P>�{V�����z.Y/�}�#v�lD�Zȿm�/N�Bl�E/�5���%uB��æoZ'˦^(��ݤ��ͳ�d����G�y��ܦ�Uy�y�J9DfSeY��;r��ku+P�*�5�kbjXc�܅A1efّ�G)Wc�r���P�{�u#��ʘ��^V�\f�ir���ec�gH;,�zn^솟&;~�~G���泧F
��Gn1���5�'e���$�/�8�#�������5ag���Aڕʆ���*��9I��d�{��qW>���f�{��fr}+�����+�w0�D�ᜄ�����Q2^���|�CPJ�м9E�a�'���꫎�xк\صe�g�=Zi��ǎ��j� =P�?��QwF�/{Y#fn��sw��9A��>�+;6�6,����]p�9	�G��vt��>g�Z�E�<��VV�����<��%�p������"9���bU,�!jhNLm/^�̒���u�o���ϭ���Q�V؇P��/�jurw^�SN�f���@�ܗ��v�+|��=�O;.+r^-���������Im�~e�eR�)�u�r��:ع�S�=:9�|M��xA�E3�Ad�� �勥��Cїu�y��P��ȁ�&qGA*�G�.���n�d5���=��a:ng�D�^m,3��(p���и�\�Ys�R���O��?5�/G�-)W��?>|��Wv�����U�lLB10|j[�6|��^��fV�u�����O+o5�kgt���BJ=uNL��\��u�j_� �=y�e3YS���r}!��v3F)n����P��!n��-��(F+rM4�Cy���p=����p
<�6�r��&+�\t��\ �?V6���gﮦ��s��z9W\�\t0�3{<�Jg;�Щ~�2�
�О���ˁ����^]���OTl�v��ѳ�#v�{t�^0���"p*$�g)��x3�k����%�GQ��;���Ƌṧ�Θ�9O3�!o-�����L��]�ZP��|+9q����3�:Y(�"�̎���4-�S�ؤ�(�齧BB�%�a����/7�>B��������W�A�k�/�����?_N��Rf���ލ+j����r��b��s&�Z�۔�W���m�Q�e�s�<uv8^�zUB�Atj�J�{"�=�UK_Qn�Lw�w��g����P��s�ME؝ֻ�\3;=3�$_Ns��9��#Ѯ⁷i��%���c��K�\�����l�?[����A���EOj�~	`��t}��#Q�V�`���=��*��o��P��&mE�~�.R����1��1�+8I��vUhjG+F&��}G�s��[G��
hU8�)�S�d��B�B<�+�j����Q�O��ߏ<|����|OՏ�O�6��mL�@	M�+.��n��J�ȬIؾƛ�Cz2OK6ࣗ��ҚN��\Bm��L�k��ʃQ�.q�(c�ۚuw�q�U3�N�����d��R{?ۜ����[BV�ImhUʖt�]��b����q�O�ؓ_RN����}�����ē�k�+7��5>ח?wCS!8�p.��K�>��&�1낉ƙ� �tz:{)��<�U;�5f#����SP�NXa��h�^ݔ]zs����j+�ci�Yo�׿K���Y5C���$T>v+�յ���+"s���o�tj�V��裗�rl�9qՙO�T��g-N����5B&�3��s}_)�Z4ȇ>�n�Ӗz>F#c!i�蚣p��E�l�;y���W�B�<���h��~#�ٽ�����{�ܡ�����1l?Zߴ|���U�?J�4����3�{�)G�t�����gWl1'v�8��~��z6%z���Gu֊��c�UEn�z��^�/2cZ؁!���E+�dGQ1��V��w��:�^���}�^KhC�
��VMέ��a�5��x1�(r=�V=�8��󮐫�:a�ͩ�TN�8�,�]�w&��w���O*��g���P�4���Ӓ0��|�U�S�7��M/M��k�8�P$J]��5��ڬv�t������֟;$a����$n[���ւ�RƄ��8(������s��՞�)�a��htX�qt���=w]3qh]�9��ALTغ�U��������	��W+�t�V�ġG2"�'t���k��	Vb�-1|$ɡh��0�b�F�o�Ѣ���/Fn��z#{}c_-�]�_�յ7�7{ D$��&�w�JV��_
w=6��o@������Y�y����[��ލ�#�3�Z����I/^T���fnQL�l{/�ʾش'C1�Ы�󳜽^D2s��B�g��䅝��������}Ȇv�v|�N��Z
6��~M������@2iO��M��秪:���+}�7�k��%j�ţ<*c���됢(\��P�잏}u���ʋ:#2c��z�h��1��`��*�{Q�]���Dz5�a"5��7�Z�~��k���_��v�FSk���jz|��F����`{)��������s����<�#A�xO�����e�Y���9�	�������4W�	��a�Cܽ�����c��[�U�S�#���TZ3�5��ve��v�!�Nϳ�ˬ����H��J��h��Ŧ0��]%����G<�1G>��G�H6Jp�u��O1�j熔c���(t��[oc��s��9��L#�LY�=��G��X��gKKc���tD�e^��ԅL�HK#"�J��e�Kٞ�ӝ��[���3]W�+�]�;
2�ˁ�{&�B�`9�c�/��{M�>�Џ=ڶ���Y��pn)��yS��Ǎ�o�~��S��3v�=�"�G�2�L]�N��	���?�c�'�ΈL�
o.�B������gl�V���o:�r�c	R�Se�(�Q�7*�p���0p��c�'|ˣ?b{㳞�^Ǌ�D�ߍ�8��HS��{��NĻ�2�-�W0#c�q�����;At�_W�cp��k�n,�!�7]�wN5%1>�^O'��W�\p�$��#��>��Є���dV�)W0�~���V�U��0k%>��ȉ�_�gc�8��2p�-*=����]��~cs�G�k����Q<�Z�1aA��N�ǫ�s�{���X�|� ��� /�?~[4(��<~-T��>�<�=���~ϝ���o�^"��T��x�D����|�R��/�_>�,�C���h+2�C���ԏ�ە�R����n`_f	Q�x��@�q�#�M^w�T�W��72 IZrl-���5)��ݭ��^��ϳ�.0vx��,�۷;^�u�rbDe8 $}|�dB�O��;u��r:;=7b,:Z���{��orչ�.?'����#5�x�Ǹ�g����t�@ណ��̭��_�1GD
�s;�&ދ�(V쨧}�Vf�\BAԎ�F=(��T/�u�R̞Kk�L�F�{7�1َ��-N���q6_%���`IǱ1�c�lD!�gv��{��掱�m�p$������5�΁"S�}|Ԙ)�Ӎȗ��S�MV��Oa�H�/�
��l�Nw�Mt��;Pd�w�3j����y�z���a/�7�p:�;���.�'Eë^���8˜lk�:4`���{���O����x��=��S��e��7��8�@�3���[�:Tzؑ��j�L?*�ѥ׫�֪Z�ﯱs�5�����Ʊ-���b�GQ\�by8�衖 d��֫�,s[��D��:u{���:e�;��m�rd��>�<����e���wg��W��}j�nH���#5J�K�ä�F���)0wn~*\��1|2���&j8���H��턫��w�>�S�׵ͣ��r�|���'�hZ�6nk7�Tb��� �.��C�(s���mL3�X����Jקp�Z*c��{�1�9z�6--MYr{jn*�/ZM"����9��n^˙���y=�c}�����ʆ�7��hH������9M�5ӂݑ�=+��_�W�pM�tEO�WbԲT����Da��0�E;�N19y�g�kgk�zQu]t�#�Z<�Wl�@�K�ULB3���up�i��:��̯ٝZ̶(,b�Lצ���N��wRE
���t}q���|��#[%n/~c�(�;u9'�m�0�"mxL�ı�Շ�G���U
�hyn�:��6���'X�)��ݲ=�,�����}	d.oS8�^pr��'ut��va�\�� o> u�mL����}"��ӆ�»�j]X���L�j\�;�ְA��T���������y�ho �ك��/�.���#S��t2w�JXhLS_dW�Ʈ���0���U<9�'�!!B��z�m٪��TDxt츳s�|�2+R;'��ɯ>`��a�[jIJ�O&�
���26�؃sΚ��(I��^�	�]+�J��
/�6h�p\�|t��麍�~�"�i�EjZ{�۳jDY*��E7ת{>{�}�99n9�� ��X����#����}FPʰ\���0�ޘ=_q��-�Yx�Pu�	���H���O�E�����k�ҵ}i5���.���ʸ'Ҧ�Ս��v7"�32u���vO_i��h�rig	���P�j���*=�?B�P��$t���󍄺=#��֙	aᘢ2�ma���
�W�?w9��O�Z�N�d�#���y��C�E�0��|�&��z�Z�7�P%���^�Ϣ���wj���՗s�P �F=�.��^��9��(���P��O������o/;|��(v��&D�������⤵\�xd�����T���-z~RR�b�����#M�<o�t��3��ҨB� �3�v����8ǝIu���3��f9tD*��]u,d�D�8>YE�3(��Wo7����Ϋ\1�fg`����8����+�)U$s��|gRu�Q
��I�0sw�k��Zq������b���AK�G>o�	��R�B�Y��X8�+�uǴ�u�)�5���a�K.g��'��J�34��h���ژ`8CR��v�˾B[�S5�v#oʽ8������T됟���<�0�c?UQ�����8�W׾Nt�J����{�^�#(�v־m�?U�V'��閨�۹�Kq���_zײ\��c���������~�ח��m�O�hꨫ6{�fj����Lhh~@�(�{Y483���Y��V�o��[G�Ϳ3��)�?烥2Gܢ�غvEŻ*�x��S��4�o5��l�~<M_s��/) ��4WuQ�m�^6�lԨ{l��^k�f*����$�Q�U;�:����z����͗@�{��'�;^Hg�oG�� �Q��~��*�s|��-D��@��VFh�DN����ɴ��y_M�=�
ԫ�X�K�O$��O���\5�Ξ�q=��F�����]^����<�+-E�������C��[��R� ��T|v��N(̓7�S�!�tj�����6�-?�d+T�}���'����f=��`��*�֌�K�^H�O�s�U}Y
��p�.I�]z8^�-v�x�m�qÒ��D�M�j����A+��H�$���5:����|If����)��GK�LmY����3rì��m��lk�VA�����Y$��Ҧ:S�-X��#;}w�k�b��LPf�oc�;�A9؀����
�s�����wҴ��p
A��k^=}�}[�#]���4>�uu�1�<�;흹�6�S�����h
10)w
�!���x(�2+o;^�-M�Ţ��F�UY/#�V2�����3Dlp�z$��a�ċ�}�W���
���{���]u�m�4d�\��t�_H�:��G�+����T��(�,��ޏC��@�#w`�6� S�R�mi��t^�k^6�/�g8E�jG�y<�0dF�sN��ܶ������
=�	���/C�ޜ���v�5/`��십*���*�G������#Z	y����X���	ɂ�=�Z3*J�,��mn	]�P��7ɱcɭQץo�N^�z�pr�S6�y9��@�.͉�Z���z�焵r����l�EU�͉�Vv���FM��v���3����6���%-˥m"��޶M������QuP�,�t�'�,�9i�:����i��vb�[&s_V�⼚�XzV,s�&����C��Њ��5�:m�V�7��h˽j�ܖ�s������+W]��� �������zˣ)�p�s$�g.�E���-�(��9f������ݑ���	�N\!��<���7y�{H����-99�w_fi\���&F�}���l��ҋ��|���%�r[Eo3ȹe��%5�cN��{��-
˖�y�9�c�r���4E��t�z�cpՒ�W][c���`�X�Ϫwu�3G;�ӧ�axE�۶�H�v��CW;ziyF��F������1׫w�Ҍ����N�N�\��:ePxt]�8��5�zhif�Mm�,�d�<�;:]���F�m4�s��o��dhLх�J�Vn�>Ku�r�72o�h���ۭܝ�ݻiq��|��tV�9B]�]�;�]��Ύ)�%[�������ѐ���x^�{-��5:I��W* ,�Sf슋ĩlo*EYC�%F���(SÈ�.CFWr����{�#C`Km���Y��w
�*wn�#��V��;
�I'lE��_a�7 E��ݧ�SmBB�m(1R���m�,rl�l3��b#dֻ'q��s����"�7{�P���Fo�Z,f�k.K8GtSk�.�L��J�]�s���:�V/aB D�����\���YF���x�GȐV�U���7�����w^���0��դ�{Cj�2��x^�5��ڌјo�y���膊���v��掀�F�ܣY�+���0�!�:[2Ď.n�|�\�+�}M�"Vu��0#�:�Z�¶E ��ڍg=�V[t(wp������������m;�ei�!B�t�.)k3������G�u7:��ދ<4�UG��c������� ��f�JP�v���R)gU0�U�~��n��}�a_�=k��" �6/o3С�ݤ��WZ�iW:ხ�;Î��p���K�Uؾ,��M�=�EsO��P�l�.�߆MD���3,O_<b���CK�\<�n�̧;�gV�7w����T���qg�A�en���:��w����$̍�Q��kB� �ûd��9"L����XsGu�}aí:�=��R����j��v񈾢�󩘄6=o�fp��|�����c��|w�惔�7��X�:�X�������ɭ�{=Xn'�T���/)����m\l�{pG���[����ʭ��u�{o�QV�ܾPglq4��l1��w���G�lr]�����t�[�:G߂�c�_w�+Er����)������ê��E�GI�Lױ��ĮX��Y-������W�V�\�,�׻)O����U����+��{Q���K�fo���­EVU�H��c%�C~۠*y�;ԜؚF�hN��kU�Ԫ�(�4�V-{ST�?G���W��!�4���3������;�I����`X���6�����d� EA�ɷ }��|�k��
�j��q�hg�Ԗ��]ʲ�	��ڳ����B���1V�1jq�.�wB5��[\1���ϛ���ygWn;C�Z�A@��I���Sm@�0��q1q܄��>j(���M;����h�9���Us�a�(��rt 6&�.uvO�x.��ۣ��z��<�v��91����=�p��Oh��u+'b*A�����z>zg�v��;I��j4\?zGC�u�D����N�MP/un����k�;��.��[�����Pl��Z'.S23����>;�����O@&��ٰ�}�����w�S숬�NL��Q��f{c��a���y)�*�n�|�j�z�ǖTf末Sc�����\
�C��L�F��X�Y�6����Ң��m���a���hYΨ�}�#8�Fr<<+���c�O3<2�8�Q'խ�Q[� [0+�9|�AK���+&G\�Cz(ʘ꣢�٫1����N�c���Mm)>�oؾ�5�퀽w��&��=~����y_��#a?���)�xGOnJ������'.%�X� �6(ķ�:�������E���ߚC�{�X�6o%ܪ��g�Z1}e�j��L:랄�d]ZQ��h!�'�͍O���AЮ+k��K����Kj���{;%
x�7Iޙ�����(AD�=�தs�;�+[�����;ٲkj��W+�9���ok2j�du4JYiVb���f�[06\S���9Cvv�85RUȎܨ��gl��ǸD�y4��~�	������m4�סy+mƫ5,�2�V9y}�x�:}ݿ��Z���=E�킌j��g_n�txj������:V#%z+M|�N�����jZ��R��8fVZ9�ٯ/��pC�pz��ΤO�\Ml�����H�	z9�B�rA}���[44�W#qf��Fo!��w�q��
�^�b��0�C��]cj���=��w�v)�そ�cլ��)ѫ�6�a�b�)X��}0^�x������%�T�`����w��	��^�ѱQ�]�Q�^���݊{�"�����[��#��;3I����:����o/"m"}�����y�qO�ƙ�o�(��x��pТU���ܢ.jxz5���p��>T�gxxް���ˉ�~cO<׽v.�C��|Yk��iB���[Fg`ϻN(>��������Q��.榇B����Y6�r�QbFu��ږ2��@^bd��+�3g��bZ,�W��x�uu�n�z�Y�w��.rA��Y�����K��7���~i����ȵ�)�{z=U�я�ھ"Fb��ΊN��ޗ�\��#����h�C��"�ϮI����>�(�Yu1J�ffR��op$����r±�V�4J��Z���Y��"�o!g��K�Q�)k2(����+�o��Αs����aۏCz�V��Mt���tV��`��X�]�R�ç������'Yp�^�~�<�f��=DM.Sֻ��e: 쵱#b�RL:[�h�}�N�Y�5S&=��.A�܆^�p��I�բ��SO6�P���etDS�P�H��qM%y�W�fTJlނ/G]޻Rݿz�o�/�.������A�4n��:��fE������Ց0 ^u���w�T�g1.�Q�PgOղ�`�Ǣ�WX��S���{M�e�uO�2&�l�;��b�V�𺉀�}�oC�"z�w�dzo��Z/��gX�����y���N_�=��}��F�Pq·q�=����s��R*�ieF�4��=�O���[�hYvP��vՊ�_���S���Vl�,m�����_u����]޸�Mݟ=�YU��fd"��"��(�+�Z-��r���=��-��B�c����� .��&ޓj��mrwp+���g�h4rU�}��dyhصݪ�1(TvP0�V{��2"� 譽1&@ۗ��,�X��W�Վ�6�V���|	�����<iĄC��ǰGU�~M?�_�u��Ќ����i����A�e����s��J���C��N�ln(�tH7j�$wSw:��{#f���ӫ�{�����[��zu:!�/��CX�71��f2�S��)�qV����K�O�:F��|&VJG/fZ��ʅ���� =Ф�@�����+kW�͸4ȸ�Q�o��Z���$B�1�(<�T[�}�{kn�E��S~�QZ�2�9^mN�����%���=���Nw��4�9�&e��P�譹����t�^ͻ����4�m�G�]�s'�y��]��S�=W/��?7@}�(H��/*��Y,���=��l�Wyy�n����h:n��r���٨�kX;��B�;e{��K�#���3,�����/�S�踝��G&�DT�|�&�%o�̪��[7������{I�x�xp�p�^�fOc�=3v*�H���� i����> ҬÁJ�c��������K���<*�{%
�U�`��NC	��L��~3��<���Ϭ@>7�����i��^+��o��~����Z����*r�g�M��j��V��*��"�5.=�Xo�F�����3}Gg�KB�`ǞK�G<�Yg�(\K8G�Z��/��*�Y�v!�޽�O%(�Q�5�;NG���cHMz5F�)p�m�6d���ݗ}�f�c	%�ƮcO��s���Z��-)��v�,�ǝ��6���Ar�=���:�1��=��'K"o�������˖�/�>uѬ��|��9��(�v��l�,j���c�t��oz� �s��q��~&��B�/&��ό�M^���9ke�HR������u����4�]���Q���6��L�O������ے�_�����ykii~}��V���N�zj��s��3U[��O��/��.��#A�r��j�4}���]��Gs�%%���V����㻘����q�N������e���ۄ�M��鿊��$�w��d�dv��=�'� ��x�=2,v��a[�UTv��0٨a��u ���>7k;��_^�o~m0��1b#��6���&�CU�ZB�鵩����MGd?������KH�\�][��HN���ݾ�6&��\�%��_�Ix��v��ě窺뛨5��_�y=�,h��6��áD�y/#�A�{�Y)���e���o�.,�M/��;��j�W���b�3;��>�b���Y�EM��C�����Ap/��Y��4��� �����'�s�;�5��psٸG�l�P���R�Z�!P��1-�*�m�����YK��B���x�@�M��f���1uB_��̥�H���^� �C0�WT���U8׻�8_j�OuCǡ;���v� n�0h�/j�>;̯_Z��Y�Vpx\Ε�p��+^y�F>
!Ȭ�Uh|;��A�����`[W�!��	�4���"�[6�w��Ur�gt�x��ޅ{��Ȗ���J�{R��?M}���ApU��\�[�!�d�f��+}⥊��m�=,��I�6��������:{��z5(�!zg3;����$�IþڈG|�lx����`����́��D)gՋ=>ݢ"��*F� �Azuo���$-���7��p�����v*=��IZ����T�Ȟu0ڵ�v�x��e��Tߤ������HWk�[��x���#����z)y����S�hY���Jb�$]Ww=�wҾ�EE�q�{^'��z�5k�ywX2�f3<�u�o��[��ܗ�
=yX\ZZ l�L�0�����}��Ӻ�|���J^�����;3��Y��q�
�W?E��F"�G��NvN�WI�ᧄ>��]�'�h8�I���L��{�5�O>�;GMɼ4�c�/ۭ},y3O7��1t�[��gb�d��]���k�!r�nc�_e�ە;抅꿦��������<����#
~�o��,+g:�o�oO*��w�)v�eȡm
��D�~�Q��nŇ�,V6F��[@��n��T�Y9׃4Vf���V��N.�� ^08��x�m�m-�t�%�mr��v�e�ĝ˒L��p��Ӱn�T�]�ga�~ѷ\)w:&�Va��Տ�k%i��+!��</4#�{u[c.����X�s�38I����ᾒ�{��^�j��3�\�)7/�:ShIm�U �-Ӭχ�{��*��6r��p�i��_L���P�1����4��� �W;ױ6H<�ё��L��1�E4.]��<9J��Ԡ���d�����&7XU���C9����7-x��U�5����%�+���;A��<�����+�N��o��WK��g�¤Fv�T_
��<��yh�cD�9���n�:݊$��.�@N7K���Ts˜�B�Gr��N���쁑*�C��r� �nY�dY�L�!����f���W.�sі�'/e��'���~�h�
��t���N�l+��i�ƴW�>T:7�,��̤�F%t��]�N���)��8/��?�Z��bݗ>��B˹��b�]�u���v:�j�E´��᫽�9��c�3N��t��9�&&p�k���'xLN�e^�{�~�� ��zs+�T�W��͛��̥���g�bY�T��Y�Yܥ�3 �꜋��W5��4���`Ҏo��O=�G���]0�]�h=7����3t=��un�q&˺��Dw'`h�i	����Jʅ���~�=�e��0��L�*���bf�O[��,�;V�jPܒ����,��!��ݎ�s�:�;������S���9��M��8�qi4#	��/���h1n���n��-�P٨t�3�����hۆ=^H]�̎�n�ƌ���ڢ����A�#݈W=�'�Elp��H͋J9�9���5B�����9W���D��hǮ��f��÷��~6|z���<��`e9��Kp���o�,�?S���ɞ�f6zI��P̘{[;�dB���B�G7T�6��#_��bƘɌ����lM}�"�ϑ�%\a�P�U�D�z�μ�/��QW�5���n��O�������.����^WR�F�T�c�����h�#ѷ	��^����?��5�	J��	۷���ϊ���V:�|ȏ&���"��#u�,yS�3f�B#u�]ʈ���H"�zn�z�(@�_�8`�<'ư!^����H�mnߔ�x���/)�]y<��g������aV����ب���SqN�u�J��h}��j�#+�s��Y��9u��0:w�ve>�+q?F;��z�w��S�����ΞN���S��w]R.7�˄f�6��2�y�eI>^ۃ�7J%E,9�I�6RĬ9��O��D�D�p��+3���K�,��0U�""�>�bݭ£�P�)y��������q�`�2gI��n�!�Y��`6OY����V&�Vl�κ%Y�i��I�q�@���w\��nH�3{fn��o�f��U�#�
%������LS1{}O��*Tt�ؽy�{,F��/H}c�y�q�ۉ��-2u���ges�ա�ƛf0yd��l��O&/]!��o�Uz��}�+}P�����s.��صQ�-�$p�t�'�q<���wnUd��g�Û1��_�T׭`�/
�J�W�n��6=���LJ;��Ü2~_t��5�����&m��5*��n�Vww�A?@�v�+��aƯQ^���sa`�������fr�Y��<�D�/{a�jv�IlZ�_P���ӗ��\����Gsq��8�^�ڐ�f��=���#�L-�����W�ƽ����F��3�jsUݱ�Ի��Q�-`�|�EG�n�hC�+0Z��5�m��y��=�ϕ�<~��k��v&���{+�(X��2�d��R��;Y��������� �?z��sK��z:���`2*25��JO�Ue�r�s�f�>6�5u��,�r�����{��zY[y�R���x���%����g��y}u>7CD��Ӭ��.m�<�s?
�\�y��)~O2�x$�����vh����j7Z5���SX��wR��J��'p�ib��a�0�S��텱φ&l��`�F���d���<���T!�mT5o��X"SFf�1��i�;��4�-��\�6��9��F`u=���s�m��t�h;�F���y��o���5)]+v��ˡ�θ&1�+�g-�F���b6�V�i��3�p+d��ns
5�\����׹J� ��T�2�܌e����p�M�a{�VB�vH��b�.⮾{e_2��֋�3�^'�g�A6�h~"��]��_�����LV���{�����U�MP��.��-���G=�Q���)��ژ�v����Hx��$F�qn5�
F����M$�ғ�0p�O�2�gB��n��k��G �ѕ�9��J��/7^�u��Y'bB�ˢ���+3���E�=�e�:���s7��pF��:9�G���z�����Nɉ�5f&6.���
t��w��#����Z�]���oE�_>���������g��6��/kLp�ˬ��������n�;V�\��E���#����_r������Aw"X��u�K��Աe�� �Ã�tT�;�-k볪r�Ś:`��e��κ�5��u�3����S�eq�c�5���Gܘ�;��V0���@�!Z�b�M7����'[.S���U��E*k*�R��d���Va�E�ūq�J�u��ΧL������-����5-0��r��L��+=3wFh�IRԨ�^<y�-h!�=C-����U�'aWl��f�:
:���;�m��W|��Ek�J�(.���a�0I��b�{$ӵ��'ۖ�r���Օ������RшS�F�$�7F�:˨��k���<����SHLHZ0���;�p��4�U�3xB�]Ȇz�+f��A�[�1gt��V�Hf_v�[50�c�=�d��LZlFެ�3XYM<z�8j��y�o��Ȅt�Fl=,]�KٗCn��C��w�9U��ɫ��gWv��GPQ	�\��f�������9o=�x�ƪ;S*7)s��;��.��od�6����}GY�2���M�wL��'.��ˁ4@���y�D�PɁ����ʗ��U=֕ �Ԭ�fc}�:+a���k��y���M��mb������U�{�T��[b�0@���!�\)m����H��.�d�ٯnfshVf��p-�dT+gn��/{0�B4M|1��r�G��}�\�Zu+��Z�
��]�řx��R�p�**fVh��������u�ih�]��0/�	U�X����2v�-B�S�n�z<yR�oY&m�8nea����9xؼ'�,Ys�9�v�E��IHE8�K�}}ǎ�Ks��u��:�uH��6��,N�T/hu���WO������7G@����oU���1[yKh��K�E�r�F�׷�����/��y_���iA��h�r�n��F�kKn�1���aEd�gq���;3���A���V�)]�P��ʚ�ո8R�Ҳ��9H���9t]B�� ��-u�����>�m�)��W�{�}c�<��E�`	�<��}{c�{d�G�����f��~�ALN^�Ó.`KT���Ꭶ��(5�,���n��3g�=JKY�SK;g�z�n&/��S>�Z�Dﻯ�)��Lؗ���OJ��߳�0BqY��2��b�3�E���A�S]a�5z��rK�d陛���<�A��DƲ�џO"�2ں�z';���We���[��.zI��^��ݿu#ǜ�;47'4s]2�*EovOfy��W(E�nUE��v�3�T0���e{�c�7�!��]��L�<���Q��6*�n{*����|�m=����	}���x�c<h�:�g��1&�|�����=z�+^�kȫS)�ǰW>M|桔_�~֯�o�Y�
�Ѓ��}>�Ƥ��mv=��w"�SD�M�o9���/�;Cﲦ�{Q��YvpT�<���^�Yy�l���_�qN�ׄ���G�w3�U�1��euW�)z�ܲqT����ᶓܹ�C�t�x�S�n=1���²&�*A\�jf����]f��B�D��þޙg�p�9��������X�l�틟4�7���}ujM
o��D���{�26����k33d15���g��ag�wX���:��� 5犽@�ݳ7>F��Z�����P���B&��i�[�RB�/�y���s�����ߏ�k�=�?,3�[��y4�(�ojLz^�ً�̽��0�B�y�R����f���Fg!nQ�m>+���;g�=+�U�}�"�K�ާ f�8�Ϭ،�V�6�g��� O?[�#�\<B�֘��������+*2�(M..Ī�R���U�O��vgV��8׉r�����u&v.0��H��簈�:��&�6r�8�7���޷�~���3�����ͳ9���R�n��U!Tm%+@�	�^��}dr��%�����_����X*VOYY��U�P���;�]����z(�N
S��G��4�V��s*�B�Omɼ�'*��~�cAcqfR6f-�ض�A��ϡ�9v���Zs\ܝCR�MΤ�^��q�5���v�J��J���W��B�w���'�]1*�J��L�L�9��Ҁ4CgV6�k���)[��qs��q����p�M��d�)�{����+���U�߬�\������w�{�$l�/�4&����0Xɘ���Wt�5�л���{Mm�W�����K0G$�\�t�2Χ	����!�����H9���=�S1�Z�r�UϷ��<���v��o�߭xRAI{#'�<ߣ٦n�1ȟm�^��q��SU��`���J�����'�r���:9琧β3*/råv�A�5Dgr�If�T�=�x����S�4�3���^�&�F�٦��÷Klݮ��cV�
E�4�܅�%C�l�L)��ݲ��߶��#&���b�.������]6�u����F:s��d!�\j�s�u��w:Ƌ7ȇI3�c�=��)��С�-��}'�y�KйrS�DEp�.����G�7�࿸wh�J#���w�^��̫�Y<�\@�ϯ5��"�=<�틀i�j�{݄^p���Ӷ�j:X缹s��Vt�:�TU�^m��;G�yc��&c�^+���_X�W�Ku��	�����+s�3ygTlP,��`��z�[Z�Y�Łŉn���&+@���3:v�U�.GT��lg\��F�W\RKн}��"�_�Ma�K��<�Toz��I;�e)Oe��W�m�a�:��$����������Df����;���t��ʵ9���X�<���^����*Uհ��բ7���E����:9�{�G攀�uf��Y�_5��^꿽��7s싵{�&x��
Q���	&�.�ݏ`iW��Ə��U��W9x�l��=N���P�L]�i[�+�1WpƲ����7���{����ܸ�.������� �B�*�h]X�#/.%�E^<�3\���Ո�~̼�H_ۇ����M­��;���O��eB+����[�׌i�Z�����׻��4Ǩ��\ȥAq���z��rޮ9��KT���s�:�.'=�!S*��{���4�g����ޥ{��ןN�O�@z��?�O��2xۏ�-jE��;�;#t-N�rk~����6�}#�e��0'�[�,�Ny�3��/;��N�k��wB{l�Ev`�ec(W\G`OԳeC�G2ب����T�W�UQ�6T�a,�9�ո����$��+b���*�'�u[ͥ�QL�F_o���1J�tIY#��-�F�u&�:�-�� :].~�~����ڐ6����p�pg���"��V�WDAu�f��Oݽ�V K�W/�~�qjOfס��wsb3ޏ���R57~�u����B���C鸭7�s��\a� ���E��鳱>�)�)�C���`��A���� �7�?tf��H[\Fyf����>��o��� `� �n9<��ȅ��lK��^��O�
q[��R	�ŷի�U��~>�;Mn?	8_�)*o޹ފ����Tk�]Q2-���ս5>��[�]}.�o�&��	���n��>��*j���Y�B���gTL¢c�o�٢}@�Z9����*n�g�� ��Kж��Y���������z$��ˊ��m1�;j��6~j(�ݤ�p�Q��)�aˮ���z��;����c[�.�l[z�z��mt��s�JX��3��r��{0��\~V�u{�:��	�y�F���\�%��-�k�w1���${BU��'��b�8�Bz3�;�!Sw�w!a��2ي�M@��շu��a�n�m�2m�=�,�j�Y\�p��˰���!U��T� sxZZ��&���"�=ϳ�J���ܬ.����^C�u�y�;hZ�z�@F��{_�y����Ϸ*����f_O,>�3���{�T��V�7��u}���.������,*Rv���{��ﳖ�>�he�e(�Lw��6�4(<�<�n��)��i%��̬���o�'���o<��i��fi���Ѣx�E��ȶ�_�$�B��=��#�}=a���+��x>�[J�ð�/��FFOL\��v鸠��#�$4����x�B�#S��5�z#�9�����C+Y؋�;חյr�G�M:�F��yhW����;^�C6����{�"�C�v,�U'�"�n>���ڞ�0t�;G�dn���V�O�xP͗���/+�Ǹ�]� �L�vNϛ�ׂ�u=�cc�[O"D��+���˰p��^+j���S�#�2���7��ߺ��^"�}���gg~ڍ �3�؝�܋�r����,���<X����5��ܟp�a�5H:��m[��XvU���=|�,��N�]ub���,γ)�\�~Ղ�^9�ՙ9ޝ��\��ck������mp��y����X�/]ut��\�mtUN7�xXjf������3�̹��.�zx+��h������-�5����9|maƒޚ�3�j1�÷W�9��/{�iv��cs���:5M��W^;J���8��7�}90��:�as�x5@�',��dl��]-מ�}��(��=���y�:*��䙰�F�#�%���g�Gt�[��Yr��x���#6�8����s?ꇙ�+�M;��Y׭t:�M-X"}gE�@��R�f/�-xg�t�e���Y��%<�5;A;� P����=0�.]=Yǁ�4�]�9���ҏ���|Mq�%�<�_ݹ^�y�*��5K��$��e�ʲ{�U�K��9,�����H�l����u��#f���/d�+Cό�U����ۚI�����_O�蓅ܨ�:���m�fr�M�ї��f%u��Z����kU\�W�lY|��.�M�g[���RW)Z�{1�Ǣ=>ʙ��nV: �Qoge	Eӛ��V8eL��k�dm=�!��H�ͪ���C�E�^j���A7ܧc��WW �v�r��oSoo�5�|���[�:�c�Si��cJ�@�**b����ێ�I٥�{QR	�b�/7ӧ&�˘���+��j9^�i?FH��Q�;�}~�o�T�Ð�z���m��{3��N�׷�U��#�lb��B��*Ԁ�1.�\����Ϸ͗�w��[�|�
�XL��JR����e��C&���:$���5-��74�ۧ�_vt�m�V��q��
���;�5S¦s��,�0:�2_�iK����ָ]��
����N�@�띉�2.YYj�f��������|����O���^w_d��t����������s���d
�A�[�3��1���M�����L�9�g{�]�$~�侘h����k��;¬��4��:����3k��{ѯ8]����e����7g;]6=��i#��=e��(t/�ܐ�D[#}�V�p����T{gTHFB�i�:����J�w�*y4�rr�cP��9C�B/���|a��/v;J�؂�d�{��^�KI�0&�ݺ�xܶ����Y7�����G%�Z�LKC�HAwT�@ŞOo����.{]��;>�˱hy%��NF&�޸t�2VB�Y���8�Ca�����B���p�j����:s����et�2�c�9b;@�1ޓ[�!T`�fn�(�g\��*��{�F�,��:����{��g_�<FZ1LF��7׆CD�{��|z���%�όW�7�P�����~��N���WHR�Y��<DI��Z��I��ћ��t��3}RW}�j���nO��*<������[v��z�wG�{��q%[�7~����|���[�ٍخ��:�s�s�J�����v�ѹ	7�Q	o��߭�:~2~���<�}[��8�{ޒh��'$(%>;�sc<��u=�]BW��uzb����z�~�o�g�~� ��(V�Bj�J����o}����On�畷]FGn�ђO��(����:�������)�������7c��9��'�S�I�.S6GF>v������;�>����޲dq�~��tvyo��Ώ>�j�MԳ?/Sn6�.@�����r�3�m�1,f��Ž���GdP�C����quޞZ�IR�[m^kcR��к���**���=�:�Ɯ]���b�j�&�܊p����A�s���ԝG�����OފF����K̳���G��U�j-4F�:Iı'R�i�k-ͼpjإd�7x|���]�p�c;ˊ�46kjx<�n�S3��V{v�Q=W��)������G]�qa^�}�@}��+x�؇���I\����#uhi�e�p�PN��E�]o�L�*#r4%�ܹW�~��fac��2w�J�p�S���sK����]�=s-z��{�W�Ny���y ��ޜ��2pϰ�ߕ"�����ך0��q��w�oc2�o8�~�ן1��:������:���E���7��(�������9uJ6�m�������~���u�ݯM_���5՝㥟/Iu�v*��gq;HSўU��5�O�Lwǯ��~��n�9��;��:���媊�y�ӡ����%$p��E�������{�xʫTyU���ǃ�-�Y�}u"=�X�;�$-8&+�y���Ĝ�F'�r�U��tƓ#�7e���j�/�]_;�Ov���V�ڶ��+����e��v�݊wo�De�wP��+;/b�b[N���l0��9%���7��k��r2��J��]('s.� �����G^�N����|���>��*�c�\S5����7���o,z��gf��p�<�����|-t�AWU$d�ƪIz�pFVQ�'`R6d9����yO3��LWq�Ct�r����ʬ[{kB�|f+����� �.��*��p�a���̳zy�'D�sݍ/�$����n�g-���^��v���
�{��c[�ŕ��eiY7m����Gm���}�h��K)h�:k�G�o�������(�2�����:N�5o�Ts���aJ̷ӵ��x̥x�5���+yv�ހ���g8{h�W<v���IjK�|�$Svf����Qy5�ڲ 㫴��U��tR�K�W�Q�Pc51�LМ�П8{n��)�ûq��"���N�6����7-@La`.�����b� �����$LGOXd�v�VSW@�M<�5����)v�5��)��XpU;��s���\F�yt��Z�V��oQ���{j�����-DngtP�^��Y3����ݢ��.�����+ߵ�`�҂��/-�cG}y��>���ݴ��6��9\�z��X��F�ѓ��,�;����vę�V^	�b��sV������;�xPDo0A,�$aV�}�n�T��aX|zɐV��+�HKb
��Ӑy�ާv(���P���eX�������+9E8*gN,|��`��ԕ�Gc.�"��2�ڽ6��=";D��.Z���6���v�]�d��-�jy�]�obgW��boT��,�����1%����q��Ȅ�
��-$.bٽl7�Ǳus�5(�xj�=�T��s��1sUC�>�+��YD��(Dd�Ǫ�Y���(��(f�S� @���գ4WrV��[��{��J���ˇ!9��8�yG��[���fIǱ;�KA)O7�@pV���z'N�����hfs����S�����F
Np�k4O��jӲ��W��h���FWBo0������Q�P=� %�2����������ಕ���oH�b�t;����p]'e�d��x(.CS��.;Z\���r<.t��Q���w��ŬѬ�1T��1,�凜���ɔgo�#坙8��Uv�c}[��� qƝ|��u#um T�gq��r�x��Y;����iu6h��6�]JCT&�c���,�s���Q$i�a����{'a�auЅ�{��!��rr�rqt�{2��/'gJzZ��hwY{�e>9���A�I9��[ŉqꫠ�C��H{1EB�YR�ڪ�v�3�;�9{vX��k�mg*���#@�F�#�XyeY���tN\����u�0�e�d��LM��B���� ��s~�Ue`�kzh�3�	���jL�Q} fµ�Ϙ�����ƻ*n3O{y]�U&�T�],T{ʖ]U��������r�X�~����u���,�U���Zz3g�����bG�U*;�I��yw��'A�����>>�f�]��ѵr"�t��"}��.���������R�8�퀂�CϾ3Ӽ�W�.ԣ���x�?7�m$;�"�Rk׷���*�:��2���*5���EoWޖ/���]C���{�[�8���1���s�-�N\��EM�v�Vn���7�H�gs�]�E�O���[��˿����Q<�꛵6�5��2(�(�[�\�0�e~9E�>�i�2Sn�m�]����F��̇�U{��{Z�k�]������D��a�fyU�"��8��{����r����^\�r�ۑ����M�«)��vwޛ���&�G�b�'�w<ٮ���ʡ�Ǣ;���רS��j dh���N	5�AR���o��&����;�Zԏ�Ԙx�׳)����� �p�^G��-W L�Xs{��T�yE��y�������H\p٢zwg�I#��e����Ց ]���w�C#�8*R�|i�`}E�.��Kke+�˻UҹwY]����F.}�uՑӝ��r6��D�y�&�-�d�:���"��za��D�~��vf�l� �Å��V?��wl���Un|��k�2E�v���Y�_����J;s5���c�NΪΟ\��~B�����a])�I�\ܟ{ju��}"9\�Gh��=+�,�ל�x�'�As �{���l&yu�'U����ܜ}���Oa�01d(At}B�������;�z���|�U�k�|�݊r��ǚ^]�ٝ�g�,��dl����r��^謯��e�7t�����Mw���~{�5��0��6Q��n�g���>�G�!�1��
-z_x�X��.���p��񅒁�e�zc^8����=�i|d��G�@��F�����'c�cԷ�t��U�6��~�B^�����Њ�����KQ�U��c~Nb�G
K���c�p:���w��=��gJΜv����ܿw6������v@�v�.��f)��,���ogH䊮�nK�pL��N�f{'�Һ��uʡt$h�9RL��%G�k�Tj^�6��"�jm^ӚV��	:��M7PK�ڎ-�%����px{;Aw�:_���@��\���(�P�=�go0;�I{�W�̕�W�ͼ�FOu!V(u�f\�|D���p��U���(����zl�U�����촢�^
�«���u�u���co��wf�o����柨�p�$���i�����U��·�ug2˩�A�Eµ���
{rR�{�y��\f��1���'��7��6����s�ߺ&Pz�Ǉ�4}u���p٪`e�3���M���\�㦯(u1R�${z�Qcc9�7��6��Ln[Z-t'�12�V�/=]�{�EI�[
]�BS��z����Ɏ9=ɝݑ���{���;FED�f��P��`�����=j��,�G9�{��G'��VL`�bfkb�o�����;U�·�]Ǻ¯?<�_׵oM�+އ��Kw�K^��Y^s2k�)e�zO��mZ�\�����7������!�;U��A�t�{�>Z�'�§���n��v�e�3��C��.Xg��;���T�t�p�[�Aܾ�-&6�Q�z��^��
�=2�-u�T�g2�K�Mo��5�0P/mv�o�7ï<<�i-4�0o;���m��tCj+�l��@.�������e�����+��"�χ��adw�H���'�r�L�5��wە���$�:p*���zl���n����m�|�ᚩ6P`zn��_�O����	�������V�|H�1A��
}��=A�M���ywxD�å�ڸ�J��2��`Y@\��Y�V�z�| ���z����z�R{�瓾����@B�t�y0��V~ʺ�v�{�N���[At�y�=4M��~�O�+�r��DL�k�1�sn�������4�c�p�N~���א?o�M�~8k �] ʚ��:'[!�-)�y^�c�f�����w�GB�B� �9p��w뉽�2��v�u1��w�W7�/��=LBy�Fv�[{�9���=�ٖ�F�I�}AD����ݽ7� �N���A��Cq��<�}���,T���𮭷W������x��SV����g��|��W�;v.M�S�4�Ǟy��k^�/��±G�WF�,���r��'����wX�r�.|�S瞺P
 �ۉ��(�Go��Y�-V*I����3���6J�%�F�Y�o��7���`�IA:҆��B���չ��_RW�.��5�\�v�w�yA=�X<F�j�Eְ����%��%깻_�^��j�F���W!k��V�N4Ǧ-�N��n;§J��8kg1�yu`�y��}�������f�_��F�(�fu&��^�����8M��΀�/���uA����b�$zub��e*��o�=%�P�5YԹ��6�:��{=�F��+�}'{�бknp{(��ϖ�X�p��q^�s�/g�do�of��wD�����9,}}���i��3���
[&#{��~Ĳ��u�5��}sFT��6'e�QN�g]�z�S���iy<��PU0�w�r����'N�(U��q���}M3�K�d�|G��tȯu�߸\���V}�!"�[�:�~��w�)'ʾ�߭�=|<+3nU��懫�z��[H�+[�֗��٧4s@yv���]�R�O�ڽӎґѩ��n׻�b��XĲ*�w ��ľ�ƴjA��ق �SXb=��+��8���tzr�9wk$���-�\�j����v"i�.��ѵ�+��,9g��;�����m;�eL���c��e�8˓�V�d���R(�c+F&E�I��3v�T2d����3�x�����O����:�u�Y�S5�Ue{# �#,6��P#9���gN���^�����g��x=}�c#nh,"�U���]ݳW�����{����ޮ�p�\�R�7��ח���Q�=p��Cs w��{:��kUh}=���M�it��Wҩ��v��1|v�yV�b�����n����g���S�
vuT�8��M��^��%�j�^:pEj��Fsw��[3���(n�'t�T�FU��e��8�܅�%���~�:fT��v+�WV�,��7v\<����cJ�g�"u׹�x�/�NS#�Y���N�`W,&��:"���G��AVg���Z�c�a�`L䗏<����x�f��=��'�SC�7*�ם�{S˔�w��u����3�������]��|=~�`��j&0d3ю&D3�r���%U�q��2�+m���X��r�^�F�B[F��7�j�{�Q�"����:���Z4U�ِ`�Ջ��J8w���pTݚ�Z=	ʹ�d`L��葫]}[�+H�z^+�F���k��^rM�eln��PUu�ɴ�k#s�1Иة��v���5��i��'��aσ����1T}��k'��)髗+�c�(F�sǶ�EL8�V��=�-��X{��ŲBY2���GF�{_�fp�Ei�z
�p�5_%�t�Fz�k��W�k�fu���R���cg�0-(�)��R���o��2�i��b�RϦV�[)�7lJ62������ A��A�C����f��aC���5~=��e�=��c\�##�?�
v�˻�5(c�Z���Ե<Wh�,��,F�@.}�B��TN���HEr�G�2�ˍ�Ys��Lu1{���:�MMl�gyB��.p,��4de�]ꙡ	��%�gv��,\NU�s8nt�����/c5z6)���:n��7~�UV�8�p���1ב��=S��Xy��O�����kO���}N����O+���괧��@Cѕ�:gq��Ӟ����o<i�˛x�~��Csu�s�뜺q���m^��x��v�򂧫v�?��v\��yvG��T�Į�4K��h�F���͏:]98w�5�k�V�%jl6���rf����_g=�z�Ipi�xN�m�5��YGl�u�Â%_L����U��v�r�q�B��B� ]tu�"8a�vܳܲ3�ӝA�s'������s�9�y���2T��x2�q7��u��o�'˶���:�A?�e�T�
����g�7��g6�/�G��:�w�NJ��]3�!lM�.��p`��B��|L�MyN�p���kۻ��'c�Z�f���Js K�2EF�'�C�jW���dLt`�t�Y�����,q;Y�����E�ɲ�,eG����l�N�C��o��?{���}~�:�Ԭ����~1�=x�Ȇ,w�q�3���eڷ�:;�³���F��۠�[���9sԎ�]6�}u#��[k(�&�!�Ϟ�u�w_�b��u�/�'�����^$���-�hs�X�.���f�x�4\W1a�Ȭ˱�vj�+���f�W�dK#��>-v�;���>�<{��tf{&>j�G��@�y;=<"���g:.�tm;�ȧtk:��+$]/Gݺ��<ȱ���T)ްڦ�Z�j�����dͩ��]o�X|8�:��WT��h!ZjsX��M݋���d{-���k�E�f���� �vdǺ���rVė�GRر8�8�`�r�eRk��W~���<������Iy�+�GȒȓ�4>7#����1{��,ܥp��ht�3�O	�Q����T�j�G�������yv����Q[�i�ԕ3�F�Y�U>v"�{.;��9y�X��cib��5�;;,s����7,�Ne���֛Q����N)fo�㵍�[uɠ|%ڜ�p�Q�����=�E��u$X�%�j�偛�����_�V�D5���h:����}Xjbh�Őpuـ�(}�{����{�Ox���so���kmJ`�r��٦���\M]��MFm��x^�i�3�!1k`��[ɘ�P�b�J��߆\7���@�Ig�u;+��q?���k�DZ�}k�X6����b��^�I�B��U�/���νJ�.�{^����o�o��Q�=�]\�^�h>{2uu�>�ߪ�v\���ty��C�ꭦԲ�ه~���dE�k<���������Ys]�����4#���oN;_uYdVVS1�#�yj��)��aV�V����Z�;�K�A{7����C˅��Ƥ����Jtzj��������p:m�C��V�,�u]�îe�N�P�X6LSc��B��[~�#�~��./�},դ����6'c�f�M��_,�;J��\^�B�r+'�~�������sU��d:���T�noL8��f�m?�G�*��/��%���;�Ln��$'�ni@5~5��;*`�"��v��CF`��#���^|�����$%S"Ss=v��O#2'�RR'\�w1���*s�L�;��a1�<���s��Yu�n�_�KuƔ+���sP�\Ow$/��F1z��s3�z�F���r�K�o�W\�I�{*�coVe���OQ��t�����c���i�b���Wz7�\i�뗼�/|7z%�B����O����}V_<י�`CG�2�ћ��&���$F7�ܩ�N����^�S��Q�0�٢B����������$�r��`U�]<����D8�ȱ�[����W���r����~Mn��~�C������k�����ʌ�W��j��@�����<�ƻ������(�!�u<���:T���]��C�ޗ8�1;*s�s���
�*$JK�3P9lf�/ۗT���R�u��Y7	�ή��2�X�[�۔�[{+�;���"�y�\ƭ��C��po2����]&���oa��V�װ=�3J���Z�P-9�R��Y���Wֈ��׫��V�A�C��)�CH
�=���u0�{1�	뾡�7��Y�U��eT�GPwu�u���ż��ddS�q!��D�H�.��x����|}��ߧ�$ I?�H@���$ I?�H@�XBB��I	O�H@����$�O������_��ݙ�M� ��ݴ�2(07j�v�Y��y$����N�+��E�#"�]�1�%h5�0���q�k\GQ?���d�W�N�Saen^�C8�	3(v�K��O\-�&B�*��V)�)	۹�5B%y*Ip1z��[l��75�W�$vEj��P5�S9TbH[$�J�T2޶��a�#.�©S�N��V\���*B
�l����U�붘��5�z�0֪��ʔ2���2Ը=�uW%Z����oNR�i�qe��D-X0�bi�e�����8*� �P@��3]ʳ!:RkJ�)�vF��4����(]n�L�n��y���TP���&ܻ�Tr�A�c����$V�[��GsZ��m�Zm]Z��*/n�`�e7V@̔�[wE0[y��70P�E^1P*Ѳ�Y�l�ْ���P�W�)f�dy�L��,;�.��*BBn�[0�ظȢ�Uܼ}�nj}ӫ��[u��\p�l&e�vDz��h�������Id�v�7w�݊�d��n���)GA1摍��`l�-�Ŋ��CbL�rdn��M15Ѳ��T���`��6PT��j���Z*��h���p���M!��ɠdpݎ���Ն��l�B�i6-^J��0I�Y�uj�m/H�z���lP2��V2%+P�m,e<�k3V�wa�d�ة�����jnn6!o$˦�] �m�c��v�j�հ�Ӷ�{�V�%���v�Ǡ�KW�kn<�U��a@��-�&Q�v��Z��QCb���K�L�N�j<��[�3�ą�(�4��k2!u��͵c#m���֎� Ȣ�Ne���u�{r'�z�nI�]ZWQe��"� "�ĩ�0��i&�����I{�9Xv�YERt3d�M]Ƀ�b�@�Pk�(��AJ�M�r����VLR�ǌ�Vu�d
�w�T����P8����L����Xv�����kًFm�(��:���~��:�m��U
���#���!��V�L���M�������0��bтZ{pFt���F����1���غ�E7��ȑי��ے
Tq��9���b(b��J���B�tC���j�]�Sʢ���]���*Wff�B��V�U�S1���A���fP�����{:��.�O<�&	F���n ܀(k�0�wCDh��:v�
�Y���cRI.�]]�E�hWz4V؅����IL�����Hո2mtCA�v�Q[J�ܸ�&S�ЅJA�r��b��ҍ꺺�woV��Ҝy��2��3"٫DûE����D��s"1��r�#�q�-
-ڱx(�Tlم���h��Xѻ��*�V��q������tէ��\&�d�7�h	�X�d�efVn(��fj�%�mc�;QJ�Ǎ+A��X�H��fk�-h���e�+IE�A���p�*9C7e˅o�lj�Y*V�l֐?U�N-�M���n��(����"kA��nkH�a#-�ŀ^���ɘZb��I�U��ki�,ꡊ�-��$
TmԢ˼z���r�V��:� 4�1�/�4�QG3��o��шH�U�X�L�q��Y�{Kl��m
�nE�awZR���e�.Q�#+T���ޔ�~Sd�J��Bn!���P^���E�p�5������<����p�q���T� 7tۥ� f&pV�����te���n,�@��4��P��ׂ��P՝��7	�.��7�^�bh���(Ў=Ci]�.U!�fK0�Q쳯ta�r��fMwS@�Wf��2�ц<(�qe�	��R�L-S�?AX��q�n%f�?���s��M���ˬ��]�t8^J�h�ڡ�JP�ۘ,�.Q�pfW���
�hå�r��[[�J�FG�Y�ĥl��8�2YY�0Λ����*�����$8�nh�/�bV�;���9�tu��6+P��VlgYx��$
�R@���G��YWPZ��L/45�R���Lh7��T�hRk�眺{�U0�6�g�1���RIb�Xq�MKip�A���{�!���*��%��X�f@�t��tq�w�[�̧������E���^UVaC!UA�P�v.��B[50���R+̣��o+ ����͊�ƈC8�dxr�A�����P��֛Xf]�i�ܲ��%/���U�b��hQ�Ĉ�,Cc�jV�����v�����pU���la�F!��7V�Ad��Y��*��IQ�dm���VP��SՃ�SCx.�
ժ��d�7���]7�hĳ�wmKt�)���e�3Q�f^d+?{��7I:�T�-��f[����V�9`���]��FV֖�I��dŃu9r�օ ���E����+ZBYoF�h
���"��c�&���Q��1]K���@���H=usF�4�X4�n�����$���@��	 �	 B`B@H@!$ `D	$ `A�$�I$�$$ @$�$!  HO��$ I?�!!I�a	O�H@�XBB���!!I�!	O��$ I?�!!I�a	O��$ I?�!!I�BB���(+$�k1k9j�����
 ��  ���B�|*q4����]��Hu�,v�r	�@�3��       o�^�� �\��rwwf������Ve�5�i�j�+5[6���6�      ��Y,��-�  um�+8  q�;��2e�j�mf�ڵ[k� h�{�@�ڍ��k6��2��Kf���W5�*͵a�fp��Auv�j�       �!���x4��9k�;�˝�ن�f���zv��+eϷz�*�9��M������]��k�-�W��t��W�{�˷�G���z�nq{�i�m�7W���oe�=iO���^�]7���{�wn{G��eV�����t�B�����  >�xW��
�����Р��`�ݗ�i���8��m{c� =+��p��:�MuֺR�V
9i�e�1��������7.�U��x �tuw^�.�� m�� �t�s5�ؐ(s�=m��os�+��*ӫ�\��X�wty=��ѣ�����OqZW�cx{��sve�ůh�X]���Kն�m�R�L��&�:z�D�B��xu�H)T;Ձ�{oE�]���X���:=۞����@���5M������fTUɎ�(= �b�[j���݂h��x���60�By�y.�9i�z V�����={��(���V��w[��T;{xg�ڀz3����X����@J't����j�5�eU�c�JwwE �.�]��J�Oa�`�`g�ǕIZ��mQ;]��:��ä����koa��E�p���]�p3�kl�Y^����u�^�t�{�e�����I^^������W�.ou�m�ޙl=3��K{��^<�3���[eU�MFh���m��*�;��֨Qz�κ�('u�鞬7�mb���OZ/mW��z�yN����6�nWC;�S�]��6�W��`6�[5����1���q �QYk@{�z �U�xk�z F%�@w(��C��o=΀n�w�T�=�ۀX�z�ֵ���M�v�-�7Jm2�����{�%����r��{^�.�uJMV: ��=�OME,��ɀ�{�zwk݀����o���z���fU%e-�i�&��)$�,m[+cA�x E?LT��� *�Ē�H � 5=1))3H�@ ���=TBR�C ` E?�*  &�J�Q�M�4����?��~�����j���D,�o��UN�< ^�<��̷�S7�O_���$�s�6p��HI�B@��Є$	$��B@�K���$��4HI�$$	$���$	$�"��BT�O������ū������-�Qi �/ʰZV | ^_7@�d%`q��$PyT�ŽjS���p�w��:A> {��<=� E��)�¶��st��i�!@Y���܏���~u�4�WKp*2�V��`F��!��W�I"u�Lӑmb�BV�������eV����*�&e{0K��ͲX ��N����r*eɪ��³۱ZG ;�WkOE �$���c�E��cN�;)�jB�+͚3#a��S�M�T�G�;�À�A׼�>m$�YX=��wy�Rg��O9���3f�t�5I����R�0�6DKS^o^k��7�LJ�,����<I��&E5�����Ll́An+u����6�h����xG���=�|FƵ~+��	`Y����vv��kVV@��,ߔ	�TN�6x�����"�;���i�*�G��������R���y�% �L��n��f`.»��YOےW����^�J(��2�W�o�b:cp���Z�Wdũ,X���g������tT�b�~���MH��#�h����'č��l��x����J^}������
 g�`#_�-F���ō�ޤ��j�v�Z��E��.�)B��|��j��YȈ����wFZ
�[�b���6�zI(� #�	���]�J7�1���66��吶�Z��L;)/G�C�%�h-�i�mT^�*=�9���2GXc��T�Ǐ�o}w��,��2�����>��	��]�,4��,�*1$�o��U�^�|���g55冐Sl�d$6�Z�7�]y�y���Z�hm���w/ޣ�d
u��9H��f�ysA/f!إ,����eBi�H�C�X��#�_9Q޵V�쬗p�bo�	��|V�aٺneK�6[�����cMl��br�Q����}�bbc���)ݧ"yG�T�ܖ-��͚���7�A`)t���u���i��Xn	 � {7u��Ѡ��h�oW�_)��;�`,��Ym�IXVT6��xǹ�L��^�c!��P��ŕp����C�K��X@��7J����	{1 wU��Q��if������帩*̛/+��V���<MB4�Q a)�� ���eKWx���X�^�8U�i"��Ȟ�dŅ"�ƈ�l�k�nb�u����UhiI���C 5�欚��j�I+�0��nԔ2�>�R�!���(≕��H(�#���꠬m��m�7)(u^�Wtue�1ұ-m뭫��4z H��0�O�!D"!����5K�}o���2���!�+g3.���t�������H,<e@Q`m�̵_MDn�n�h;n�4�՛�z��5�aJ�����>êX�.˗���[���J҅��B<	���� H��zt
�I3%��'�r,�8����-�
Ī�c�����+� �����y�{�ǽ�S��N�&��q���bAI�����w.����E���v�dN: ����S���2��j�
&�x�^�VA@G�b#;b�XH�^jfX(�R���	UǶ�`��(i�F��zπ�A`cY)mz��DKJ�Zج-�B���V5��k�(�B�(�-*"[Um��+,e�H���B�m���eTm(��J�Dm+[h�֬aX���zþ|+��eG���Al�3�VRÍ��(U���F|���:DY3a*� 9�faJL��5�yaF7tQ�D@��q��dZ�v�E�餰:�RJ�]k[)��ۙ��-:�F�ݠNZIZ��r��m �
#P�F����Z؃1�\�
�T+�L�{{p�+H�V̪�#	>|>���dR�[WM �,�/�SeSE2Jrn#���00V]U3 W�Q�Ɩ<�t����cǪkU)�3���Bh1V8�[�W�6V�0�.2���P��T�S���ɘh������5�wZ�Pfn�����<h<��&q�'q���bJ�Ǝ�,]��^���㮴�hd�EUQUQQ`�A�����I6ɤ�&&�Į��"�!�Y8�Hm6� tT�AA`�"
ň���@1��*Q��ڊ	l�%�mX��DMR��cdjcmTFT�+ �,^0��K"���B�������T��U2��c�TL�Y*�$�R���X�2��I�*bQq���Q�J
��ʈ�4X6���Kkģr�Jʊ[ED2�A���r؊cDc1��DU2��R�̴.4��&2��R�uKM4ESV�2��.[
��D[h,+DYZ��j��Z�-��2ب�PD���m��h,1,aP-��m���Q
��Z�LJ��QGQD�*M0�D�	b�"�Tb�HA@FJ�*�*��YYl*"�Z"���RB,���h�"�RDE���0PF�0FH,�����h�hV�PU�mT
���+Q�F��ce��ID*)X-E��b����R�"�*KJ%b��RF#-�T�%dH���"�Uh#(�EQdP�H"E�6�Ymb�ijY*��%E�"�0��%�PQdX�"��� �a �2
�4(�m�R
�dQUE*+R��H�ֲ���TU@�J�+%��-��B���",�e�Tkl������QZ	h��Q��bȲ$)jERQm��%cF(��b�����DT��DU�UQ,0ZءU
�V*,��#TV",����J�$QaU	Y
@Ad"�!Q@
��!�(@��XY	mP(�RJ%����DRڬYV�*DF)"�5D�)dJ��B�IP*�� Q�Q-��F�-Z�J�P�)ihQR�h��m�������+ *ʕ�� �I,�� �Z����[-�H(��6�A
����{�����#ɧ�+N0�+,�yu���=G��'��s��'?�����24�/�e�F�r�;�t�B=ܘw	V]�iA�k]�i�e;�[UE]��anh�"dz��TI��b	+U�j�؂KUK��[��[���:��$ӓr/<�i�#]R��c+#��:�j�CQ͚[�%�����E�]Bh�
m(ؼ&[ǎ]ӛ/D�Ƶ�KZ1�TnT����Nw���k�`x�ی��l+
2V����kQ���P.�s�R,���AMg�$ ��2G,��Ҡ����M��U]4DRҊ!mb�4������UE��U�P�(���6�eTnfz��5�]��`(,��0�P��qw@�X,��!X���u{�i�y��|�s��z�3]5�{�d����R��V�T񈕀ә�oI�R���:�����`i�11��-,T��5T.Xdd�R��h�Kj�[L��y��L�q���Y.9��u�z����b�h��2���mP���f���0�hB����qgꌙ��h�.���q����p�7�@�dF<��T�ȶ�l��kU�T�G?"�i�{��.C�m���L�pnX���i��K+t�Թ�B�Hc]����`OR���6lbv��ӕiVe���ݺ���(�yH��z��'�Rر�
ֈ�:�UL�R�d�R[UDJ�JÚ�M�*�>�}�=�����ͽhV�A��C ���b�]�}w��K3/Je}�#5��l��Լ�n�mi7�#�TqCS6�Q�۶����@Io%eՍ�t� �J�������E5Ct�K�@f4�a��9�	��b7��55�[MІ��"�V��Ytj�M�P[}�-�G�B��I�Pgh�v�[t��-k��N����7�Q*�v���Uޜ6�oDom�N���V�Mj1��l��YK�V?�,��o�倲
M������>����ӈJ�^ؽ1�Nn��b��#s̰ȻKҚ۔Uf-":˶2~H��Ve4��YGEa�FX֐����#E���  �^�!�WqV�6	�.1P�`�@�P�U,�B���[��&�ūn9,��/f]V�{����P��֨.#��*�v�Y�4kF�ZB 8��hcgtO7�;��OVV�#Z,����ڬKlX�d°� �#+O<��5�9��o������y�PuaXT1
��w���S�XW8�cw��56����d�	�����A�pTԑ��<ٲ��p�-�᝼��a�o�ɡ:�R<aY����P;lw3O6l�\���1��5��d�`[�y����[�Ú���*7�k�++�3Y{" ���ǋ[]��}�l
�Yl�.���:����^ܕ�mQ�i,�
n�ǉ��K�B�8*���GlV���`�ikբ��F�m�9�����n����ز1v�� a28�u��X3i�z\s%�����
-,bL���܉���(�kV�m�Ex@|n��z������K�>V������×�Պ�-��\��O���K_
1U�<�{���7��"Z׵j�&zY�P��U���
M8��ΡZuA �v3O1���f�b��Fa�i]���
�}l��y�~����$p:IM�۹1�>0)2��eJ�.�y��]��ΏtU=�o6���g�[��&X��V�,i���lJ�1�7r�=����i�e�yf��':�H����*�\Ìԉ�vk(`���v�t%�jɴ*g;�8`�z�/��Ҫ3g�wٙ�qS�[ҬP�`)��`�����v �\Y�ox�RޠΖ`�ÆQB'j�T�����ra�Q���Ź��f�8�S�Q7�K�90�|��S�	�_v�p���*6���ŋ\\��"�aէ�q^XM����(䕋�i�X��	�ۅ�ӖL��ng���q��f�����/�<�����R.��%8ր�o4�)���i�J���a����qG%�rL`�\�@�+�}���\�;����ٻ9����4�U�wkux�����FK���	e��ח[��ǞbF�����&v�k�L�n�1� rM{�m�4���u�Fq�`�Cv�)�ٚ�6c]���2���_M�|�s��&�.{mY�^�80>�i�b�r�f�c��+�fl
��`����&��U��H9��{z�aݕ����ҬUe�-���N����Q7����\��[�wm�^��N��)�g��3KzC�R�Ub���kZ7�/���V�تQA��5.��/��2�V�)����� ֆ<�朒Yݢ1�|���:�
�s����65�s���/v���)#[��L'csn�0贠׊����z����y��UZ�_/�t�o�ǘp�4K��c��/.���w�%i�Fot���]��j�;��g�d9b���	�2n�spb:�͖/��t�=�E�<ܟ���#��s����w:�>�Z���J��K��8Sm�[Aκ��B����Xjw]�&a�QNh483Q��z�QSѽ����lвz�.������|b��}b'�.w��vJ���|�ެۖ�G�]ŃY���=:t]y��u:]��U��tBd>�sIWYR��8�[����*�z^=�bT.�4P�����)���.��ƙG���lh�[�x���tea㏧Y��P�9՛��K��4LM*�u��X>�A\X@&+Dvq-��d�������$�
<�ڎV�j��ڒ�fq7Q���c%�jd'���]`�������:�Yҏ8�n�#�H2L�0�Z�Um��e�t�\��-�$	�����p��bL�#�z�{�L�G�it���D[�8w_-�L��2v�(�:'��aJ~�.s���Fj8�9�ʽ@��u�W@O4�/��zwS��#War�lj��k6���٣����ᵷ��;�:����[e�]��t�C9��U���!��ъ�-�#x����n5����{�\+i�Ra͠h[�H�Æ�ө.�Q�6;{x$�3S�o�.���r�s������Mk���x�y��
�.��l�[����ļ�𙀠+�Ӧ����ֺu�4H�j���`圬������N����b�	#K��\��U���Q�\�ܲju��;U3mc����	��X�����G6Σ�kֹ]i�/y�JG`��-�xtKNb�2.;k�ppGfT���c�k̺���q늺_#��왝1��4����7�J�6��\G������edpwd����.G���S
�$����3T�%ԃ���<x���ӫm{���=�I��`]B�=r��Y���>ͻW5���/J*��-f��B�c�H𱗿��Z�;׏�z�uԮ��Ѝ#��X1����]@&e�-��3��\0ԵH)�É�1�}��s �sM�Ӈ ���Sx��N�i�\#)˽\;��wXR/k�M�5o�M�2�T�1Ϧ��m����r��*�Y���I���R��a\�V���[�tyʹ�S�9�5.ڝ;�n�xc�C��Z�i���Ck,3�$�[}uq�ٍ>���2\Û����[v*."��L�ЁYHg\P)�t���*��#�P	���L�M�:�,��:�9��w#�� ���a��w�:���_Mz�-�(%�>�����ѻ\���n�[�%)��6漥ܲMy�L��Q��PW�;�˗�L�W|Y�Z��qb��z�����o\�uE�i�_kf�`�Z�up����Ш�����Z��Gl{�q
p��ǭ�,F���gm�KIwpي�#�r�ѿ۳X<urdV����⾮��6�v�=�tZv�_ju�DS��V�N�}��Iw��=׼y�i�c�e�V��t=g���Fxb��򽱋�r"��7�^N^�}��m��wzI �-�lT�%[Z�l���h[Vж�� ť��  ն��$��� M����M�%m��]I7e�-�h�-J[j�@7e�mH�m         �BH� dZՑ@-�C-.��]  `��� �,�@BȠ��   �%Z �m�m��.�m�  	 4PdR�V�Amٲِ�ّ@��B  �m[i���n��$�jd�� h�$�e���5��I�Y���ue�Y�QZv6̫m�)l�Y2&͵v��*� l$��#6ʉ#E��ZZɶ͓[m�m�b��jm�%�f� ��B֊-�@At.DZж�5��5[�D�-��lY�d��Wj�#7m�"V�M�jVY���mm���$�ۓu�d���ܲ��g*-H��n퉥���  B �@�  � �@      �k$�m0B�Y���7�KRH�Z�]Im��d�w[�d)�m0 -��hd��  V�ڄ��� ��4P0 `��  V�B �@��m���@��
�@( 0ZE  +@! h�a�-�-�k��m��,��@�m�RY7`ۀ
ձe@n� 0[m�]ݔ�&Iim��%��-0[hŭ�����0m� E�� 0Z [w�P0 `[mh�nl��n������s���ϧbV.!��K���|Z�� �㯌��h����\�+YƸZy�>8{yf�P1� ꝛͧ����aRN���/��i�7�EtG,������Ú���3&.�ǒ[�=wQ4�]�nG����v�4�_=�Xn����k�y	S�ZE�[�����/r�H�kT���Vq�R�]˱7���n�;�頣{���%t�C���4޸-L�!�JBQ��e])i��b��ɗ��Zj��"��k5����t=�;�Bt�zy+u�mI��
��n�l<D��C�`�y-%ۺx93�#'K�-a�nt�x&f��m+�pgf�r�H7�.�_ex���3�s��e��v�g�w�
�&)��sA�4sʭ�;�hSu��f0vN��,�6p\�hQ5���\����%*�)i|0P��Қ˞���b����˔����&o�S�D�W -.�7��Һ�Y�^��i_R�)��/����,�i�5�4�s!/���ٛ�H+��)ٝ����HNӬ[�0��ѷ3��u��G� �"̌��`gu�)��+!Rf	�+e��;7]�4�+{x�vl���a��6�@�[ݻͥ�*0x��Z4��H+��.��qb�F2�1�����[��yԣx��˶�vHu^&(o"O,���6��@��y���������K�ic&e��k���Ne��`�y�2QLr�x_p^��Z9]z�s(.��}�:��Q��B��t��ٲyݿo��%J��[�f��]ݲ�HK�#-�7eL�dݻ"�`    ��  ����F�t���e][f0T��]]eʛ�n����,�ی����Vյm�!wir�ۻvXnո�IL���6բIlZlF�[R̅m�ɲim�n�$�[i$3j�e��n��mb�P  ��Ԓ�ݶŠ��[idQ�Y%�ݶ�ڑ@7Q��Pے��MIn[4�Z�v�B�!��-m�ՕRՃdU�mvȷR�$I( � m�m����n���[�m�%�2-l����m�Ud������]��6��r\�id.ͩZ�$�$�۹d��e�� ��VK��VȓaWk���l���>��~�ގEN�ƚLbU{��\)X=:U�xkbv,���7��u����wh#�1�פ���\��/��B��{��)&v�2����\k�][��6���!rm^��g�CS,[ܟ*�q�5;+�_Xzs�j�����2`�Eo��a��}���k*$�����W�~s��$=p@z <��y�t(	gwx&{h	���§7ad��
�N��!��.�rz��P����a��X̕:]�|�q�!GG��l������Ύ�����u���mt�R��3vj�	Mma��V0w]�r-{�����n��qx��Ի��f�m,㑳7#�����`u[�$mlY<���ϡԃ+1Ԡ��u���ҵ�r�p�Sl[n�[��   $��RA4�-$����B�[��2en��6��e�%]k&��e�K�d��[E��4�nˋl]��S`    m��  �d�b-      ��                                 ��   � �  ��  Š �В��l��V�6�E��Y��f� �I  	"�@   ��-� ��͖���[&�腤%�� �@ �ն[v mˋjK�o�\>�X�1��o]���*�o@7��+r�0���hB��K,1���ܵ�IԽ4"<5�I/@<:��jw�+3��\ү�Gw���H5��s���{�i_D��;E��.��9�J�-�|�fZ����y��j��,��ת��j��رu�N���M�2�wqǒ�n��P�R���mL�R���,�Ɍ%:���P�hvTvɻ���:�u���1�x���˶��Ѝr�-t�L�J���\{9�_}�}�}v<�g��~�;������.��Mմ�t9�Wu�ŋ��"xwdv�7[�%�7�k�=N��a棭�V#����Q�@!�j/hŹt�Rc���9_,.���h�k���E�ńh�^n��5�r�P���m��){��s8	����zf<P�d?r��K$����W� �w.�v�v��0�(��<�{��0.�s]Z�X$�l]-AnS�;2�;a�u���t[Y���}��ۻ���c2�|�h�z,pw72��U��hY,#Ń��n\��v{ԥ�7��4v*�Bj���m�rP���¥�;���1YPaz�s^q��bt<}|T���;6��ػ��E�'��������v�zi-ڝ�99et��z��]�OM��3�&pF�����:��OEot�o�,�^�YE�wN]v����X��n��(K��1��f�)ۄK�E��VCE�M\ܣ�囗'Y�^$���u��x��ji]�g��S�����[�<�Ź3c=��V"mp�Oi���^ˬfv��0���Q�:[�0K�{�"9�N�z����Gc��lv*.vә����S�$���>���l`tz�
�)H��,�{w"R�՚�v�q1�N�5+��6��ܦ#��a[W�2��
��ڨ���Y�|��ԏ4c�o���*�,l��9c�\��ӛQF^unT:Wt�P�S&����9��E+7]���t�1q�#�m��"�]_�e�����{c[ݗy��A�oD�e���b��V��ӧ�7��l�g���/*�j8yiiFN�;%uD%w�ү�ɴw?9��ǐ=���W��Z�j�n����5LQ��}x9`�r:,��������3h��׎��,�U/�O`X'VH�Ut[��4i�V��X�u�h�s�O�jD�R�dЋK�$�\��oC���٪����Kx�6��AV��\.f,�L�	��W�H�TG>���>o&ʕ����(����o.A,��],�j�yP�Yt޵e`A�O��� ���w�9Z�P�M�I���[;�r#Ǫ�aS����0q�
l�sj.cr*��4��e�j靀 ld�tʓNM�&���e�����S��n��[#[A�6����O�k�M�9�{)�v�("�Y|��n�s�h6�e��o2�ÏK��܉`1uP�m��˝S�q�Ug:kT���A+�u^t3��2��^k?��(�T���HnIBz�	?���% O�AHI~��m$"��0!D$I.�$0H@� :��P�?���I!����հ!P$@
��IR������@�4�]4Hu!6��)8 y�H�m$�BC�y��aw�&�,�ܤ+'���
${Bx�4��d9�'X{�a!R(
L7�� c�6�,��]kZ��m����G�+'�F@��1;{���B�˙���2e�ߔ�;��7�bN彤����_)�<I����/]�̰��o�+�́D��.'�������m�L��GN�e�'�gn�V�({ѰrÛ�S;�Xs{�N�tv�[D9������8�5B��R�g���i���{qܚM�6s��4�=D�GD�Dt��)YZ��a�f�.��O
��w��Sl���Kne�K
��q�m�Q#{�E�_f?+�t���U�b�-�0+,���J�<w���z�y̘����Y���8��.R�nY�zk��uw�o��j���׽��Y:���R6�Ч���v��'���y��:�U�ʹ�a�3YC-�S��>yU��ȽF��'N~�x�1�My+3ݙg�w�}&}&���H���_N����@_b(�_*#�0����Qx�1V� }@
 �\7�5ج|@7���.\iP�W�%m�m�7@��]R���GJd�z}��T�זYv3�u��w�-�U`�-E���:S	21��W�n��ѓ�K�ފr����Đ���P|jv��'�7b��^�c9�	��d��Q���M�(��K����WPD�r�D��%���씝{����]~o-���#�V&�C�.[�4�GM���3A�������2��!p�ن��$�-]ul�.��Kr�t��YF�����hN?����]�e9.!�3���"���E�C��<t �Yy]M�_LZ�l��?���BUm��Y*vh��o�v�eX�.��"4��['d�j�@�B�r�՝��n��g� Ǌ�[�-�:���	ru�⃇zų����K`�7+95��(V"!���[���>�B�F�'iuL��W=�Jc`��n�	�Jv�X(����-4j�@䙻��W)w-����U{�J�h��G�[Z��X#l�R�!W�Ħl��"�u\[�oM�LR�3o�*/1�J���D�0�.�!54�u���'Z�֡w'������̷"�I�^�m�G;K�"�:�i: Ebڠ�״�Yr�,,g�+����-Q���	�˕�cHl���b�hi������#�T�Q�h-����A)��fe�]k��ʛ��|�4��6�!�T73�ӆ3ۤ�
Mkdi������Y ������}7`�}�B���:6)�(^4G3��k<{U�r+��͹��k��1\Y��֙rX�)*�]�S;�R���h�����\e�l�K�xJB�C{�X�(�f]��W��#GIeӆ��Hݻ����w[P�v'9�,�B��G�x��9�\
��5f&a��i�8���VV�Cs%p��j�T-2�E��A�y[n��)'��$��ZK�e�4�tP�%��lP������m۽d@�;Pe������ 1M���t,[B�P#��3M��2	7X�ڕ%U!l[�o��L:��c)���j�:!Q���V&�^�3�,�j���(�����n,�T���t�i$Rv�(���C�v�?ՖhmF�����m�GZ���A� ��f���9 �	Ի���4hL��ԡ6$�ڬٸ@�pX�K!�l ���'^ˠ[�GDYaw��l��{ɗ{���ٮ��'f�&��B@�<b�޹���)ShaP8`�h�*�Y��w�G��pYN������`�e+�(\��lKr��EŌ��p+���"Ƚ�ĽyFD��;xm��/���M�h�j�
���PDC���:2�e�[ˑ�B�6C�J�e��vfV��Y$��m��En����"����1�-we]�- �t�AQܚ�h��wf�T/]��XՎ��FT�b����-e������J� �v����rQ�x(cf<���JE����iw#mh�Iɒ���aR�^?9���&��3hB,����hrb�V�x1�U��]�ImL2J�Z�R���+l���d|�8�QV��I���(�,2�o�>�SQ�EpC�IbY��^��\t����<��r�铍�6=����ֳ�˞�wf�-���:�)y����Qv<�/(c�б�c4ֹ$i�J������R��S�
i��,��v�{j�P�R[ZI�5m]f���8�*3X���v�A��(R�K"3TQT�������1�%VP� 0��]�#Y�`�]�Vk+B[�C�0��J@%�(�6�f��|�Rdj�[J�.AOMMw�>Zv�W`�k�͖̅3L �ka�ؘ��ְ�嗵ˍP�c7.H�Հ���ILvp4�6VT��b����Y0٧�tV"��p�qf�M�KTag�Z���`6cx��6ffXam��V�bP��#/S$E���wyf���-{Ef��Ŵ�]z�B�����)?N��^bٔ��Kb�wPu�n[^�"~��fjgw-z�T�Iꤝ�y�X�a���*��;�m���]��R�������fmܖ�f�!Qe����֤��/E�K)i���)Yb1�d븬ZV(�'����;���U႙� �%��6���.F�l�A��]��c�mT��n��̑�Ԡ�P�T]Цh����H�D<T�k���ɑKvY7 �v�~�SR�F"�@��{Y�aywH@h��l�!�.��"� TEI
�b�-KI�*�tQ���/Loņ�lT�5��ۼ�É��J F�-�3N�K.�-,���ud:��ӓi�B�m���Z.Ҵ�꽛 &��������w����v��ߩ���@��wdM���\h
ٳ���e�c\��{���f�2���sn�I��5���{i��w(��(�pd��Y��[����f%A�jDH�َ�.���FlZ���Y��C�7GAƇVb�914�Ǻ��l;b$��dW<\� Yz��]w� F>8�q�~'�z��.=�m��;El���ģ�%"�}�"������W��].pǵ��H�lnA�d����uc�;�&S���T�r��P��"����%ʹ�2�wh  [ham�h  �-�� �Y1X�j*FFI�u4���̒	6l����#dȖ[�j�Ԛ���m�	m� IFܒ�$�P4P0 `�� �+�Э���m� ��J�w��m�;�3�<%��{*X��(7��K���>X�C)ܣ҈Z�v�,�F��;qwhw|��m[�;��L=�^YYj����<�rvݱ�ڶ�h ��-��Hf����d[�I1wB�XMJmq-��vC-H-�j�ڶ�ɛ�ɒ�n�66Y7�߮�N�ם��~���}���x_��M���A�{�X��r�:���>���w�ϲI�o.[D�f�.�.I��V��e� ��       ��[V� M��E�� �11l�nK�;�f.�c^�4Vz	�;�E������Rꢳ�wu�׃�ma��C>:��+['i9ibpժ핎f_]s�S���0nU�0EH*���\���Ǯ����W����)��͕3��2��=}5�W;V�:��r�����g��.���ܶ�6�3�w���6���w�{;�L�]	���1%7rj����7H@+$m�Z[��i������g�N�@�P.�*�5�Ӷ�b(	h "�l��Ǟ�~���w<��㽻��U|M�s4H�D�H� U��Z=�on��	 @ 4�����BM�$�x�$�@�H���1$�Hx��H`d��$���*H�H@�$��
C�I�$��Hm���CI$P�C� �&3i	�P�K儘��&����_�}�OX�QAV"�+�X.�� �EAQ�U��YTbZ)�TPݬPEUX(�1D�������R,]4E�(ZEP`��(�F*1r�*
�EH��Ŋ* �Qr�b���<�7J*"EE�*(�1����DA�*�+U`��Qc<�0Ab�����"�**-����EwB��n�EQ"���"*� �v������Q9��J���� �R�&�,E�,X�"GT�H��
��*�� ��X���b�i
�X(+�2ѓ-X��4@RcQV
E^�_y�5΢(�$PPDb�X�*V�1AQEQb�>@���EQbn�Qz�EU�V,U�(�D�EQ��X����%Ug��cX1����%��fY`�Q@QH�5bk��(#
r�Tݪ�TAUH��5�Ӟ���s�����pR"���U4���Ub[TX1TV�P���X�V��X�r�TQUTDD���DըŊ��u�LT`�UE��ZuJ�"��X֫x�1f�`�Ҧ��,4��dG��z��dQPDS)c~J̶1��DE�#�X�ݱ��ӹ1T��(("E��H��\�����TAV-B��QX���+�X �l� �)�X��ccO��1��C�
�%��ƪ-�DU��9�������{���g��_i(�����DRW�DEDYԪ�j" ��
�������E�VEDժ�P]ZșK﹊*3T������V�Q�G=��Q�Ucy�CN��>�EV*�M���7J0Q+Pg͊�h�9�Y�G1�ϭd�]�qr��EL̽5�IR ��?Q$f��1'߈��n���9~L��+
��RbTAiQ���U]��7B�6�qX�D��~i������1T�Vi��_=֕M�Ͷ(�({e��"+��#��b��#�UV�y��
ϝ8{gi�}�c�Q+X�B�F)���E�D�TU|e����GIE�cc"��_2��U��_�s�wU|8�49C��0�QQ����oF�0�q�g��Wm��FDƂ2�5��**��f"��q3�J�Խy��2��
��a2ʱ-=֌6*�Y_2��;���"����-q��Fe��-1���y6�}�aWTӈCꎧ�L{3<z3����h @ =��ɫ^�f���R�}�(���b�҆�CN����O��_�f���"�[���\��v�=�QrùQ���_(Y�*.��2,m>C�k����m~��/u�%�B�D���=-fܡ���v��ڿ=���u���3.L�ƌk̢�ts{5����O.�k��9���4�ȳ(u�*"����1�"*��}~ͦ=�+�__p*�(Ƶ[oY�C�)������Y�Ӟ��w����?x�eݵ��_o9#���e�ن��������컒2�5��b��u�����4w�}��
�W.��0m�5�g�ٕQ��/S��k��N:LbV��,���`���9�sg�Yw����0����P�D葴V��wo�wy�t��M']��1�VŨߓ�ҫ���9��S�E`֢/��{����{J�S����-���kx�����n��pzθ�-�����T�׹�H���, �L��(�Y��1��J4wڪ��E�e��Vsy[1�;�m��#��NAV��;�Z��V�U��;�㶯6�#��â�l���v����f�j�����	��uR�f���!}q?YL3G�1s�7��!�F?Ze��"��s �dD��J�9ߴ!�>I��^Y1���T�Vx�VLv�r�]kD֚�aa�S9�����'Ħ5���N�3�!�v{}x�ާ��� �P4z*�_Dw@�������n�}wY��(�o��\k�_��9|��Luj��S�pѫ1{�Y~w�D\x�KT���=h�AaPO�%ϳܠ)Б��c���`4��U����JD��@�+^��T^;u�w7n�ɤ׍�i���5V�N��~�#������,�X���C�e�~�5�6i���>}�i�t)�̲�7쁘�4� ��{e��JI���,��D}#ƨ[�U���񊄯'$:�(Jԧ9�i��CiS�i��/ֺ�g��oV*�"���g�<Lx��
�nyt�;smP��B�\!�?;@Ż�1�g��j�Ys�/�}��|�1�I/�.��氙��Jm+!�M�;����q�4�9�[���4�����$�l�YLg&�\C�]����䕨x�i�V�+�q��&}h.�����r���ώeW��5s���5����c�8��4�^��L�Y�s<C��0X9w�Y���w9�xuݰ���3'[�az�j�q�l�>�>�Z������~����i�"�f]�nDw��Lܜ�_?}�y��n����q̤Fx���wE�Ĺ.�\v��&�f2VUٞ{�z�)5��Ӈ-��ɽ}��[yq<C_Z����=�3ۋiY
�?3�Q{�^C@�?�s��}�w� ϫ�Iϫ�'!u�DK�x��,%r������欬3�G�[��t�|㈡�}��]0�m8fg<t��C��X\����O�p�%��%�k�q�~��b� ��tϹLG�`z�8óö�Y԰r�J#�}�'Qju{#Do/@dx�}՞�e�W�w�]q�>��P�W�i{0����k*����Qj"���Nsp�E}�H
��(���<����<s����֩�S��&����ֿ37v�)���^�}��aR��,�(��[�!���IS������	䗃)i1M�콆��37B�0�'�&V��3t��o��I�������%V�<s:���b鉼�5��ڡ� �w�˕�<���Dۼ�1>�ԟT��-Ю��T�#]"(��W?2T/�Y��E�m�<n%T�7C6w�K����X<̂�m=��I ]W�C�q8t�ƶ�����J�mX�)X2��|F�1H�yc~4G��Z}&��B�)��	*k(|���u����隦d�t�b_�n��3�Eh��GE2���7ݞ���ɖ�g�!��ܫ��|3�S���|m1)���p�ґ U�B�ɼhI�^g�|]��qP���^e��
��/.�[��%�{r��*�6�d2+���"vQ��;\D
��i�I�0q3�Ud|�f��7v���`E 4Հ�|Ҧ(�Y�sݶ(r{ݞs�l�n�6ےw�2�7�I�ݾl�;��>ɿsSL�m�`�g���WN>\�}��m<N	�Mv�~���SI�������U3��ĵdc�A�6�Wy`�;I�wAH������Q����L����� �-c��"�(�TP�(��O5*�:���/k�a��߻f4�ea��q!��IAp41=g-�ï\�j=��}~	�1�I>�EUb�q�cGĳ��]��>�R�A��\Q� [q�yH���uH�I��	4�S�~�|>�a��~5�>t�M֯
��GY����QҊ4F<��	�ώW���|�"*�Fx��3,�Y>q���u��~�>�>[�ǉ$���g��Զ����^�pۤ*��2��0�[i����c-�7T2ӟWfa��:��as�^-}���{x}c�4i�!
L�|�{a롺�)���>q�'��LMk:0��#�l�#Ď!�U��[�J�d���
�	����'J�!�qͶzE�{�1���M�ʭؖ5�+y�L�E�̈�`J lBCڻdݮz\�}�1��
��|�"7:t�D����kY��%#ܺX��jh�׉���퇇o9�]�v�raU}�"/���w��{��0Y���_�L���>�&e������>���@A����P'∖�.60��{�һ����)�9'vmWwA�9�i:���e��#�ru���tf5�=G�XX����}	�:����	{xf�Քa�[t�	vb���{��;f�s}�~�nl��ۿ�7x�Z�C[�no�=5E2ՅO�\rY���0���J�� 3-�/1� �����p�S��Zr��'����<cq��~���n��(	�6Yr�,^J�Q��@Q�nA{-��zo��7s���x�ZU�����$�X�������b��+U77�I���F����v����$~�+�I=7�ϰhq����%���sΫ-&J��{�x��P|Eڟ���|�t����˖�YD�����{�z[�W	���z��P����}���AU��B�>��/W�DD ��i�Y�Xr�Y4�A�`���9eo�g�j�@U3�$�G�4쬊�#�5�`�W9����B�y�!޷Gg����G8�C>���յ�;%Y�J��Ǝ��]2@�v�ɍ�9�h���_]�5��(�7�a�y%��`�Ǫ�Z����)S3��>��`�L�s$�sw�O�k~�˟�6�>�zH4���oU����A�!��(k�Έ0����B�V��ny�:�Ю\�t8j��5gp^� KA:��������fv����?e���kw{0���U���͉b����-& #4[Y�V�V赻�m�Z$�Iϝ���w��'�����7e��Y���Z��T}1yɑ%  6�$����t��m�Ԙ�cC�2��O���+���#&ő�&It����w����&["~��.��}ݎ�笹ٓ���pY���c����J��h�nگ�;j��1��N��?F��bJ
DE"��n1Z��,mO���ӻ�(��.��(U�a��p�\j�o�%��n�Ɛ@|�%o/]5o�GD�k�0��Kj$�+�c5�d`(�z�����t��am���x�O�l�}��߯�|X�"�fP�(膸t4��6\��D*8��>`��!E�}�,��>�Eq��zF/f[*"j�#����BUb�y��X����a�S��ѵ�0 �A�^��4@ Rߣe��sv�vI����o���3���|b,|��=�*j�P��(8͙-�y�ڙ�n�?nM�ω�5�=�|~Xl�C^D�`�S�g�kO�W��-���@�^xɮ��Ee��XW7�f�1�@�X��)T�?���Z)K[�i��%6s9p����n��p�MC��eqHQ��>� 5�,�O�B�~�`}hFx+���X� ,��k�W�-8��F�E$8�i6����l���y��y�����n�+�c���P�<iU����s�ZMYb��^�W!
Z@�z�Pٵ���<�x"ЯV���o����HW�W�� f�P�VU��2������~!3=g�n�d�#�QB�T>>׺�ww+��㼐8N�Q�����z���wV�� �!�		@&�{� J�� |���$@��a O����C�$0 � lV	��n��	'R@�J����d � =d��$�^�		Ϩ6����A 9�I��'�$�����S_>[n��.�۝����(j�w�l��0�c}ɸV�'�8Iqr�qa������n�a��wp�S>N=�О]9>�1����#iךv��T�o%򴬞v�	�((`�ۭҙЌ`;���Z�v��K�Y���3B�����|Ǵ>f�Ӄ���N�D3��6V�|&�vj�^���ϊ����A����&��_���𥌿�Dq{�hϨTl�F�88��d���/ku��BZ_H|�V��%ݢ�6�5RK���?u��gs��=��6�.�7'�b��6U��>*���d���q2����>lf+dF�*f-F���>I1�j�?@Qt���=/�ji�ZF�6�b>�X~"�i�� �8c~�vg�<�ҬFHg��D�)�(5�(0=C��b�'ڜ5K�LǑcD�O�T@�>Us�;����	T(������rK9����{{�>���>M�e������&t�:n�'����N���Z/Ƣ�K�����G� �>��b ݬ[/>���X +Qt����?��q��2lDj��_'��;��י�P�$qdۢ�:*>f��9W`�湓F*Iw_zp2��>{ƪ�X���� �
z�K�M�$�>dW�J�th�H�\�]j�H��)��y��7G�6��&������M��/P���v^eEZ�>�����`-C<�1�,�!��<�dV�M�E�=�n n˼�ڽ�͉�ᣰgb�Dܱ��5��W����2�d^����Iu�Hk�B�\ �{�@�sIn� �,�7�n�N}θ�i��Ș���i5��k�^vj�"ڽ��3Cmi����M]t$X�����[�����=J�N�僻�� X�������ĴF
(�PP�7���ѥ�4��)٠)+��<m�;R����b�R��O�ŧT��C�|/��|�Z~.ɞ[�>�o��z�wb�h�tTf��J���,;�P�y(���Y�񦽹
+qފ�l��jVx�*�5C��B,��q�2�����i�
H޶��hF��罨��Z��s)�bA��Q�`�doe|�
��L<P�q��"�֐���gg�3_�����Ͽw�D��V���2��ٕ��}���{����'~��w�q5�Cƍyw���IQ��$��M/!u���45)?f��v���ײ�����9���K�?z9�@�40�$��7c�Wu��lw�
������z׃D�RV�V����j���Y( 5�Պ���`4���?��f��^GF���x$8R~��M������S�u�����>�����^ץ\U"����z�����'�I���߯��g��2R�������}�ӟT>�͗p&uW�X��-�.�h�l�{�u���z��ϫ$�<��y����q��3��`Z�k��k 7�P�+��Ϡ��d"�z�8�������*O�M2(���Y>����m�<w����x��<���a�����fM���W�Z�[L��c�o+��>x�pF�:޵ծ#7:�yԲ�omA�I� nT����/�ݮ�5�"&ޙ�)���c�]�:�M�ZwS�	�5p����5P��Z"��|V<����dmY�m���\��_O] %��Nx�����n7A��J�.>��]Y���0ݻ뺁�	0�goj���֛CI%���.�_���C�nH���x�˻�ؒy�wn�>펫��^;$�4 }����V��2�I�����@�0��񲻦�~���߷����8�O�����ɳ�����p�
�Ӹ����(q }R�;���ok8ӷǸw��3�'e=^� ci�Qlp��ڑ'�xQ��m�H�#َ2k���<Yo�4���T�`ꥷt5k{�oȠV� ]�:��A��@m�Յ�,�C^�:�h�b��:�[S���iѹ�(Vz 1�����L�s�w�P�L��1�cO�ط�x�E�T�ˠz�b����^Jп�j~�pnQ�0�h,r�Ƽ�^%�Gԝ8a��"̑��Ӊ�+/��Ѣ�����A�(F��W�W�cob���,�wӳM�Kƽ;���j�yT�њ�0z�ٺ��\@��)���;gt��E�%�{���e���cq������-�7�)��v.��p�Y�i����m�F$0�I�ƙ9�"����	������l����i�{v��n�܎&�3b�{uum�]���i[m��)$څƶ�d��qE� 17d4W���'�޵��w�{7vl��IK2��������yy����  �uj~�n����/�s�o��׾��<��6V�H�997v��	�o��s����Z0=v�1��}�C���R:�Fy߰��o�;\L'��2`5��'\�� f�0Ⱥ��t`�%���G���) ���eUp�I1:���F�8����oܟ�2�U�h��}t���v�v�_ �U0|�J E��&��lg_��p���@u�3�h�������U���� �m�n�xFױ��<�h�-��6�l��%��Fi�S���{�1@�uh^/ƻz�I�+.�7�U�$;^>����)���bN��}�\�(X���m�:m-|M���j,r��,ou
B���B�wܦ��1ܵ\I�借c� W^I�<+����q��I(���M�ҵ?���XQsS�RB,��^�aמFjϐ(n�,�=��ѥ����.��T�ʰ&F���Y<���R$0Ef�v#َ6r]�O7���<����#�#e`�� X�����ג�`��P�F���Y�d*����Ev�_���㯽�Os��-5D+N��+��i���Q��kLn�lg���*���%� ^B�{XFϑ�Gt�ò��w��g��8��Xzfr��	)6��&r�+*I��ˌE}vN�[�N��5uݦ)���gE�����]��Y�S{Ǹռ[n��5���8g*���J��+�Xb)p�RN�~�c�'˙�}<���7_~��2yn�+�{��ܫ�TU��Ѳ8$_����"���m߸{�쿌?l=��@�T}����3t,�ҕ�\xU#�nM��*u�f�vo+���m?w]�(��!�v�
0�m�H�{���/E0YH�V\�Jp��<�!^>�:z��o����m����H��l�> V$�4����C�w+�T"mߏ��^���u�/g����ϴ��*Pth0hw*Z���-<����pB��d�.wޕ�`��`t���{��x93�;�q�^�|F���bB�o�����yr�i�����?rXO�-�&au=N�͟�����;��M���IV��ۜ���#5�b^�T�P�rz���5Ʀ��1�|���t�6�@
PV�&�6�v����h��wI���kï�V	����|����(�CqQ1�W�+"�Z��K��l�t�^5c ����Z"t���*<䯜�}2g�ϵ뛏;���7�>�~��n��>��>��/�D�EE�UCq���<����h1���\��y�d�-dߝ���Yϟfv�h��3� ���N;R�����`{߹U)5��V>=�0Ц�m	��2���������o��n��ҧ]EK�Ӎ�<�m^j*+��Z����!9����_���[S#Ö��"Y��r���^�� �R��J�p��rD!9�d3KW7����@��/�<gդQ��GHn`�����_,<g���g�|���Z}�*�_�Խ�ظ]%L�>���!��~�K�H�v��7��cp���s d�4����r�r��{k6""#舃���R��8��˱��wɌ���g��䕨NZ�C�.��	� ���f��L�������6(����$
�G�E�㎅�H����%Oi1��H��l��T^�!���*O��ORs�$�A�n�Ō��=YW��^{T���LPU�
봆?n��`q��u=�.o1u}�9�>y�D�p]��;h&{|ϹWy��I�}Ө�i���#α��w��	�`���V���MG�՜͏NI��;�B#��k}`A�:\��ٜ�q���]tS�6m�8�t���"k�\�.����{\�HA
��3�r�a<m�ˋ�v[o��7���%%�g-|�#�&��<l�r���]���+(�R&�;юO��d�p4Q�wq|�q��u�nM��ν�����+����*ˬ���A*7��Y�ao^e�j:M¤��u���>���_sc��kGM�b����Qf߬t�Y�����[NX�0vYts��$,KW�ffk �s�#��8�!� 0�v�n:r��;٘ҵ������&��w��QE�z��!�h���:���`Bü�,p]����y����-ڬ����@R�Q�W+%��TNl.Y�cK�ূU��N<��)G[� �K�p�	k���O`M/s gq����4c���d���ǻ���x�`vo�?� ���m��vv(*���:V�!���ҁ��+����Yfs]�ws�)ڢ��vh�9.��w���{�{�|�B���{@2!�Mc�hkŇ�I��u%G嵀i;�LM����z����s�}�i�������a�W��f���[��bLC���ӦSY�ĝLAU���y����#�=�����>����ȧ�2�*��������Ĝq�-9�y�@_��z�&����4���sz�^n�����Ý��B���W�LaQs�rT� �#.q���#�#닼�q��[g��������N��4�&��c*T��p�x����Hs�O���N�f*4L��5��k���l�x�����y�H(��!Y�Nk�6�V\�[&&\��w����~M��2��LT�|�x�ҏ	A��U�c�Iɞ��������RTOR�P�V���۬�+���q#��4c��Xbu%a��ϵ6�'���i�>��Z�m����.��=La�����q���V���ɏI����OreFuD�;sWЕ� �(;.KP���F������Z���#�s���L+�c�?&���a�����i�x��4��Z��"��Xb.3�(nYS��b��v�5�1=wˌ4��>9���̰�e��ܧ�P����yʃ�|��G�l��?��:�0��4m�yn;I�&w�&�CyJ���l�{J.٦��yt0��S"�)�D���ϻ˞��<OSG�OsdƽpE8��������<��S?P�����Qb����g�&$�v���i�1��i�����T��Kh��h�S��\�4M�]�L�c3���Z������9�{��|��uCuK�J9a*c8�OY�������]3I?&�a���:�XVW��ٞ������J�����o���	� 0G�d�Ch���f�Z�Z��5jC�k �W�񘂛j,����}�0�Ϭ��'�L� �q���iD+��[�:�M�XpM4g{�cP�>�C1���WM��u��������5�6�Y{a�L+*|��\���/�h�^����!y�ѭ�k܅f��[�S�L�i��9M�OPϨg�oӚ��{�9~OY�N�0���a�&����Ww[�^������|F���b4G�C�nfi���P��ydXmC���=g��q�*z㖁�_�i/5��N!Oi�/_���٤Y6��
�yw�r�:�^�I�]kf2fX����+��b>��ƻ�F.B�p�fT��SO;�N�q֜�<g���Lh���;F��`u�CE�<�7�d\���b�����ή^�-�b������Ξ{��@�'ۺt��J�}��1/�a�Ld����m�r�vfw��δk��봞�3z��w
���bo2/���*E��y5�~e�M�"�V}<�5���Y�7��u*	����G�+�A;g�g��B�r~� ,ؑH��`�b'�_h|��P�*�ۼ��j6��<CL>d�I��&�wTȞ��H|�QB�Lx�E�m*Ls�W�=��u�����'�s}����nFVn�I�IH�ShZP�����H�x� V]�x��9��� i���8�x�N�&��+��j����H��V��X}�����<�Ci���q�hB�H)�1��C>���s�q����yU��Gٿ�?���Y��x�`���b�I��4�sz�M}d��ٴ�>����:ͳ'��g;��!�Ma���;~��~u�E'U+Xy��󼶀���~���hn���l���o��Hj�����v+�~��xyM2z�:ͳ�,��!���y���ji�~��n�T*VKZ������.;�ﷰ;��m'���;_,4�1�ܳ:�1���|�H�)Y���f$�P�__�s�^f�xj���\g}���4�2fwN��i3������80��8�S�M�2�"���
�x}����`u5�>LG�N�`b��WԸ�x�֬
'�[Cg-Y�Ĝq��y�̽�j߼�����o�e�Sl�����u��&�;d��+O��Б�q�i�'�6�\θM~���Һa��D�}�n�J�$���.�x�4�|��k��ߺ������X��k�3%}D DAԑ]; lVV�3�~��T�O5N�"�_.�Ϭ6�I��g�*c�e1�=M81a������1����r���1��x�}Ci���z�]Zֲ����'C�`T�}桂c�!���߻�܊��!f����ؑ�p��"ҋ^����J�Ԭ�%�{�f�x"ԹkC+jJ�CI�!��{�<���?$��t<5����=��X~CSL�ްyAT*O+���r�\OY5�~�`T��ڼ��[�ǽ�hC�!��Y��?&�<@�3,���tq�'Y�l�M��Hr��Vy.��b/�~a��}�	���
�y���cX��ۇ^f�>z0؁Z�=��I��Y��
z�9���
w����yc3r��Bru�<zskz�j2�T���q��ʆ4�fm-Z=�
�)���mr��f�B㟛CP��x�w�v�++j�f 'Mƍ��%��PRd�Tmcc���Dv�c$�]����9�ɾ}�^��en�T�t��m�+�o=�=���˻��  �l�$\��x+��Η���+V#����0��\���畼������?��3&���=�<}��֦���M��w���ިiח�Ltɉ��Ͱ1��sWI�Syx�"��<�\Z���a�)ɿ�Ѵ�M&?5<a�u��F"��8�>����*�|.�/��_w,�$�
�Gư��V+��~�q/�M�w����Q��&%B�ٟf�ԟj��z��YY��y���}幫{�}a�4�S��][:����Ci�Y�6�����k�~�a��
�_�~�~�o^��k�<��_��g�2"bO�
x���LX~ʸ�I�+���� �߆���k11�����'OۻT%a�ǩ��i�(W�Я���'~�?5���o�Y�N�������)^#�&&{��L]���xܻI��4�*+�3Hx�qP�r�v��L���3�h6�V���{d�bu�e�[O|�\g�1�CY3��G�>������j����޻9�Oi>���V
�����(i�3)�M V��>���)�vq����Ѥ�q�����v_߽�$�6�eq���o�c��c���}^ۯoOuqP�<�y͜G���0�o<<�����y��>'7N�SIP��Vv�ĝL|C�f��3�1�>��ݼa��YQC��C��Y5�q�+11
���3�!�K��14ϛ���P�C;�0+�q'ۺJ���>?A1D!I�>S9Z�th��4}�{l�"OR��?f��~�H�5�߭�qY���Ľ�4]SdPR��^a:�HT:����*iL{�,1'���Lt�yd#�O��D![�q� l]z�O���}a����Ĝq1 ��m?y��پPFm5�Zc{��0�ɷho����$���w�H��S�Ԛ�f �S�̡��X���9˷䙪T�'xx��\I�~�����or[.N�&�j{y��*��9x{�X]֍zi���nP�Oɤ��I�����=j�X��s�>]R�j6�����%M����L}��T���t��8��
�B>�ǲ�DzG^j��;9=�v�����I��"$������F"8ʇ�2���
队��5@��紛ݬ6%k>J��������]g��XTs���y�d�(f���z�>z��Cn��ͧ��Ԏ���K���g�3��!�	��<qPoէpU^�Z����ȧt=��Dy�w��2%�G�Շs/%�ʺ�Ub����n�5 ��SEAƠ���K�j�Cgv�z��#;e��A��¾TP��֑I�5�C�w���p�ҺJ�wFi�q4�CI���:vϘc��fښa��o��i�,��i�6�LK�6�Ձ�v����Mrʕ�*7�t~�W��S��j��������޾f�<`b>��|�5و�#��|uu}��u=s�(�2��1|�=a댋��y��u}Kn��:w�w�d�
�E7�ZM.�c+*���14���1XT���#�y�n��H AB*��+��6�z�M�L��Tח�Mv�kXM'���t�gi��}�i�Sl�:�Ӹ�����<�q>f�R�ݕ��R�1ؼֲ~K����B�����}���vx����h{�:�[�?2u�q>���=����������M�Y����{�&�e~��6�Yү�L�(z���皕:�}̚t��7���t�é��'^�N�m�9��:I�ۈ�{��+S�Vm,14α���#O�O<���{��a�0|���4Ǵ��*(~2���5M��g��Nn�
��g�s��~zO��%Շ�sT0L}�"�9�h�����]=���5���Lzf�h�<f�1'?41�%a�i��W��&��VAyI^��y�~w�WԐ8�h�I�PКq �����;9J�YX�9�}a�Dqua���&'����a�{�3�a�x�G{ɡRT9�wT�����,1�����(u�Y�� � B@G���Ux��ʋ϶{g+ke�nE}2��'N����w�fg�߮�0/������Ɏ?�Cl��l4��~�3h`��Y|�tN�M�P�}�#�+9������XmLa�e<d���y���hW?5�d'�5�"�9�.�;���W�̊}"(y�G�G��D2b��"���}�_���[��*iR��/�K?��|��1ߞ�ϕ��\�.�Ȅp��V���B^�_Yv�{�T��P�kۥ�s�쏴�(��P�lWo?گ3׏�y�3d�������۱��z����(�Ȧ��ǟ���C�h�h��m�A`K�8�/�g���?-�F�����-����B�͜'�S��k�,UM��++��(]�0��eN7�֥��.h*��k�6�q��^�*�ۅ�n�'����2��I��9���]j��:�:vf8���[pd�����\�uȈw�莼ݹy�i3�E ��U8�&�5�tW�j�'ݾ��	
ipS�Ŧ*W��R!��.*�����7�D���9��w����TV4�n}eޮU&d�:S���Z>
��eI~���J�e�����,�7O݉�}P9�D�e���4��/�A��I	 �/�6p����H��+��9�����0���yY��������Ί�:�Z+=!�$���u�Cb���&H�SR�1ؖ%]4=3킘��m��Y���Q���K�i$���y���yv͝ �R�T_��˼RTR$T �G#����oA��o	�*�t	�q�{4U���G�����l��y*Cl�����J�W5Z�����&�@�!�ᬺ:��2��_C���JUOl������=�.�\�>>�.�H��C�U`0���N�+�PF&�B+��$�!�$<E��C7���p�d�i�<�m�́b
�Yس]�T��(����k�'������jУ�،̷�H��y���n{&s�-d�)+|,CtCr�j��Z�K�2W4�%ʀ*ڥ1h��jV�
�U�%���#=��Z<3��Vax���ɪp/e�m"���1]~�3^ݼ�^���$8�4iw��L����:�#(~%U��\M����]�Eaʗ����EG?Yn��.�N����sv��>�^��c��"���c{0��{�ͷ2���T���qBS���@:�'��-�{{���o֗��$k�.zF��\�ۯ2#�>[�,��Ec�o=�d��Z�`:�CS?�h�Y���>�u��2�_����uW;����x>{����s����~L����I4g�rZ�z8��қ�Ngz�ԍz�{�j��_y��� D$,�
I��U�9�(H��i�=ҧ�X�o�4(|+���5A��72�V�j��gE�#J�[H��%��hO{�~�v�_�}�8k�EU('�8�K��ġ`�%�kq�U��� �
8�0zR�؏9�'�Kՙ�e{�yb��#���c��Ҥ�S/��{��^�g钗�ӳ�>Rbl��	�QoQ�Ι\����Ҳ;�wxN��ӹ�����T��\�ma%û7��r�0��
���RXs���B'x�D��KY�k����������h���٫�[ْ��<��(��]�M���&ҝM������qG;-T��.� �P���pR���
Y�L =P율�3� �ǯ�Ύ�)�֨a��"ƾ�OE�&�fR�lgC�U^���B׹�azLbI)�L�P��z�f�Y7�o$���o�L��P�a8��:��7��Rt��vo=^��?4��=t��P����2�:&�;?�ɋ�Q/֣�w�L�ct��_��uB�nk��Uy�_�
�*�y��Ik�:�H��f�nXʨ�^����.��V�\$.M��l�6n1;N�t�mu��K�6�؝�lu]Dݧ��T�~��B�I!��*�Ԋ�dIn�T��ܶ���2HŶ��皹����g'�w�l�ԍ�k5�g|��מrOs�nZ  m�����~��_'}��ٻϟ}��y�E�����-��G���F�ǿ��|�;�I��ɞ��w�9��{���˟��L�L��5�`�Vo���xXS4���2Q�[]�7�}�-�$�w7%��^7��K$�\��K��6h��6�@ʅ*
?���h��al��6������#]�ׯp��q��H� ʱԠ��%��A�t� f���Rm%w�e7Y�h�%����ؽ�z��o��D�Y=��zSf�^����P���s�" �H�Uٗ�Ri�;ss�6��i�tE������ʪB�*׹5f�l��G���8�����yiu��얞CX�Y�փ(���Y/�A�����i���ma��z�g��ɔlk4"|X#��;�K;�:��Iy�ˉ�_�ި�L�^�w��7Пu{�.��z�CA�h�(�09��5X9/��ƈRU��EmE��.e!��>+Ǧ=�3�'S�U7W[.��&��N6�[�������{�3Ƭ��f-�Z�Y=&���V2�m��V �`bK���<;��?�6�"�.�s����sxM�||��v\I2��&��:	�P�bժ�.\�ؔ闖P�V���<��aʅ�^�C|[uUd�~|���^	pP��Wfͪ���Q�5F���gQ���
���	�t�]��ǩĽ	C����s9g�}������릻-ٟw���h:�Na�<1����*�p=,)m���Gr�)(;�|����%�c0��/�ΜՀ񀃣��˒q�x��gV�b�����s��#M�[Řf�� ^�$�n��~:�xU1�lN\�p�3r�؄mF�RP��_��nlA�&�Z�"Q�X^�r��_C��dԼ�TH�
/ĞO�iR�s��Oұ��OX$]g����"�R��\ӎY1�1��A�uC����e��	�J���É9Du'���oE��w��%�]=>�E}�{j����m]�X!�^������{�S��md��I�� ���Ac�E̡j���|̮��9����.Nuӗ���[���b��v�ؽ�լ�t*BKS��=ـ����F;��0$�n���Bc��cCl�!����d?#=V�G����otb��=~���]��a�Cڡ/��j9;��J�P�����v���j���ab9�MFkp;#B~�L�<W�̂s�l�,�����]P�^�gv7>�0	��
E>�LeZk�LL�o�����l���gҰN��+��
:~��$�gK�h�#���~ڹ�����E@j4)E��7k��v ���n=�~�-�$�O4�T�Qk2椾�s���u<��\�p�T�+�_t���b�fc{q�B���S�MQ�F7?dS�(\LJN�����&������ѷ�0�Q��C��� �!dFT;7K*Y��6�#�a����%d�+ŏ��_>��r�{y>N�K�(D�f�Dr=:v>�j�Vcŷ�`����e]ڕ�ps/���qȺ�ƟV�os/���� ��L�|ڨ�kW�|�%�+�̡�X�1��.;�6���{s�:a���(��͑fo+�Q����+F��aq'��᾵�wx%���bBF����Y��Ҹ�ez�_`tX�鹮b����$a�(x�7�M'�(z�q�Bob[�^�g��E�N��A7ϙ��&N�t>ؒ�RW�!�:m�dۡ\��c� BD`_(?Yr/)ow���g��fI�2N^��8��X�1����@�q;3�0�u�#�]�i�<K�,Ln�=��VI�غ�Ip��{���Ǘ��y��[��ww�g�Ofy�n��Y���~�č�u�36>Hz��⤃:�>���ߩ̙��)��g�3��k7ɑz^5�f|�İ��,��@V�n|$>n�ڥ�e|Ǫh�}7�T��E/�woW�%����3`��&��M�YO[��p���	�C� �ҸOi�s�o|*^>�w�+�x�w���v�"������B���WZ�Ո�I(G�X�%g���.�6������tvd7֑C@6��q��|'K��R����q�J�'|�K��'�
+�����~қK3��E�N���ԩ�K�V��]�ܖ\ukQ�v[�.f%5�t^3_G[�ե�ߴݳfY��RK3w����I:��ޥ�Uq����ۤ[�s��u~̈́�k@���b�Hk�}i�@Н/&�mt�V^b���c��#I��g�U̼ �o����jl���KY��.^�Ī� �+�Lg&4�g�ۖD�ʙc����͖��B7v�Jp��^Q��=iP��:�[�.�U ���-�V&I��׹���T�0} ���u	�w?eظ��S�W4�գcJW7�~��fE��ғQ旷Pr �ۿ9���۷Ĳ�lw�k&�V����� PXOA�S��	�KV��ߚ���W(��^�Q���3U5)F�e�:!#T�C=^NOX���5=�o�=Y�>�|nS�{���!r�2m1ƫ�ڮa�%��85��"KH˵.���,ڣO]������?����8��K�iN���{r��H���n�������CuK��7P��"�	K(��@D�
y:f�Ս��%D�RmWAT%�߽[amZ>�4]�c^e�YP�ʄmu�#
*�.ɸ��|�OX�W�����\�s&	� a���ɠ&{^uP�s´��u�.�W"=)u-�P�����R=X�z���t-C��;��(0��0���=iY�n�F�nB��f乂��(ӾqP�zbXu�stn��0.��m���8VG+�Y�����&��]B��H��u��r؍�<.�L\�e�/���<�W-�c$p$dR44����NX6J�Llj@IZ���H�F2���c�g�>�x����W
��v0h�:����=v��g��^���j�5Ֆ,���B~r�N��8"SO��ٴ�mA�^��W�x)�Bn�+	�̯j(>}�_2�7��u�d@�I-J��K�;t>�ڶ���A�l�Ut�� ��(�1^m1b�	�X��ӫ�\ށՄ�x.�����)�Ef�=�۾�zڙ2��U�b�{�@[���GG�t�_ V��z�e�4Z`텛<�nk�"bӝ���c)7�Qk�kFqĪ���'l�;l�22���0�걃���Ʒ�rU���B��k��S�;�ƍް��l��؂�*)���_`�ڥ��m�F�WZ��T�>/I�s�*�;��\呧��ذGȭ���O�����τ��5Ѯ�Z��N�#3�=\\~�ax�7��-[◗ܮ���+�3���iW殲P~:�
�N�n��(����"����޵l��4iI�M���9vĘ��'��n����>���R>63�p�w�^�5��\綻����>�|��O���}���=\�����H�S�}6�������y%���� ~�������G��[ܥ�Ϯ�������}BI�U<w�ܲp�����&ܚ|��0��l>���{�#Ӻ�t;ei��;�C�Sm��d�Z���FK2�D!^R����4�qn��5��Ƚ+z�!��R�mf�#���A�Y�u�Y��\K/�XUf1��f�c��Y��Q[	��ͽ�0��ٙ��]�.t��|�7ZK�B�Q%	A֤��)Ewm�3'J+i��}Pcn_��[�a35J���C��Wj�3)Mӛ�.�wp��nD�QE�i3�����nM�4�Z�d� ����X֒RM'm -��ْY$���n�j@ m�b�E m�.�m�,��cl��vam�d�$Ʌ�-�\�jI�6�7m�j�ɴ�n���k    �썍#im� � ����[n +@! h�[�-n��M.�,�o���m &���׿��=��rjrr����7ɓ�]��&۫O|��8>i:���U�8�Λt�u�(���P%��o����9�w�K��L��Q mˑ��l�jE��Kn����P4�jZũ%lŶ�%Xֲ�`�R�$��j#XͲ	5.�vn���y�{�������/w�{��Ҫuo*� �l���ߞ>�����y��w��h$m�6F�.�sf�b� $��        m ��,�v�[h�	"��ݶն�k]�N��w�A\Ǻn�����Y��<�%-����eӫTa��漘x�5�fj:�eh�{L���]�O�����4���"굹���O�<�s��7��GJ�]�۵��SR�ȭ����,�;;�)m�WrK6�ϰؙ��w*xn=�s��7�v�<<�=�goJ�W(�߷�s^{�Y�}~��s�;9��][E
�pKSf�YUf��?�����m��s~��~��s��f{M��Z�vK%���?K_^s�����ض� �$�a�\�St6k�������=���չWk&D�#��7f�ٽpI��ӌ\���DW�UmG���y*V�	����Dt��0��2W�v�c����'l�oX��=%x��x9&�ӌ��q�d�ƒ0���mL�����t8C���9�L�}�D��Q�,7ere�-��1���s�޶�+��Lm������KߺJ���bf�^�`���f���`���;� 77�1��;l�uDl����}��:��?���y��I�׻?W�F�,���ǙNr`:�<̃��p�vQ�:�Dk�"J�V� $����3Ȥ�! zu�J�.+a-OS�~߭1��*�MnL_��x1\�2B@�������4L���WO�$
ө��d�~�;��\t(��"
�sǄ%`b��WQp3���u�Ri�� 5*3ia7 ��{�7ת��I���5d'�܌��0�`E��(�-]>�x���m3k[B85���.sf��vU�ٴA���L��~�#G�`�����nl��L<��Qp���SRo�}vͳ$+c5r�~w��/��t�~$���Y�]�������`�C��S��O�/(���l��b(��+\���~����|����P���;��Ƴ8�@l��R���_ՠ�&`ay��z.�ΐ�SX��+�ҭ��M���X��=F$^e��u�,!��e�������>}�'��)�/V	WVæŋ�lؓ���]�qk�_{:�I)�9�4�m���Wm�&0�xK�[����.`��n���]u��}��ʧT]w���!^5�뗐��`	�b1Gʹ��#GV-F�_U�f;�9Ԣ��Z{�zV����E�w�L�
D�8>��
Q"
�P��
����Y���)��Ɇ�Քꉋ�f1>���^튑�А�y?
�"��L�`B
��C�f��E�T*2cJֵ��vR��S@��Yb��
�i8~�K.zZ��O�� Zc|p#L����
L��xG�� j�8�0�U,zh�����3=8����-ip�U��θ®n0�4T�~�Hk�E��o�p�~�O:5�(�=盽��l�S6����m�~��Bन�Jɣݳ=�JG��b7V���^����]���!�)��K�y;��YA�}�o�+��8�3�{G�1�s��3+.�i>A!�sY������O�e��dWQLm(���w�5��^{G���֮[�/��dWL&"�B��p�3��97,M*;�M���͇-r�=6KF�Z&��՛ob�vcN�i�d#�'ٵ1��.�1�'��d�&�~_,��r�~AZ}%#kTN�j�O��>�.�F<Z78��FŗOy�B; Om~�i;�b�;	j���]�0���ٻ�,���c��U�-�S�ӄ�`\̛9	�M�뎡�NN�԰Nd�uA����q^�ճ��bN&̌���,�;�L�TOuC�B��Ch��I�F"a�r!]�ݗ�{����G�^j��rts����l��F�Egޒc�-�+�p<�Us���� ���hդ���P��ݫFbazjhV{Tp�4U"w����_YY�����	\�|�^*�wy_\�X�W��6�_�w�5���l�q��;J���$��8�*glT��mK*W���䳩C�د�@��R����ߪ��'��	(���Jm�#���l��S'�,w
�hr�D��<�$�^Q�.���?$ a�9k�������'�BJ���Q}~Kik�ʛ�Θ���^�I
2h�n���S(�D/9Ϻ����"���x�mzz�g���5��
���ͫ��pŃiJҰ:��9���>�3U�������CG۶���u�N�b����0��^�� V1;�>R����{n�h�Ű�z���V����r�B��Q��*�����gb��?u�S������Tȵ92�e��P��6K'��g����F�^j�Ó�Pm��Rz���4�������xffFJFG��1�"/[n�^���o?�7�7��������yݛ3�[���_�|C��@n�G�@�����?if�Ḱ�K7+D�ESr�֍�ܗ='
a�^�����*���}l�s(�cov�n�@�Zj�w���h��Z�n�tjzx��E�c���)[M���=$����/�����-���u |/��&��B�^�W����2��e�(&��� )\d�9՝/��w62+YM�n���M�;%A��7WI��M�`�,�1�������}����*c@�H���M�}�d
Ҋ$��Q��"xQ��I��Z�5��br�y�0G3�I�.R��=���U$�y'5�+{"|<�����^��PH�
*�Jm��7�!��0��FK �r�%�|��0�~k��]z/�ή�Bi@MW�@���0e����
'f��dx��=�V�V�����j�s��A�|Ӫ��Q��J�ŦK^]�	�~�$*M3 rtl!�mı�WK�^��*�Bt��v˯t쟴��Hʇ��Y��TϺ����Wy��]������#t���o�-�JNu����;�I�o>M��g�7��=����?�{�$U{'z)�§B�:�� $�Q�nl'&�p�E�!Ԩ��kڮ#�>vW������?�+�na��Ջ�,�`X���ZOW�zX�@���e V�^�b��[Mqk�]��3$�7��N�<���)����L�������<�zI���������[��?��q��#�|o�L;�����N3�5�,d��0A>t��t�z�ﻩڼ��S{���Re�6C�G;qpV�ݏ̒ډ]��έUi;��K��<�������|��v*h��Ccn�W���he��*��� :I"׻+^H5���T��$���Ɍvܹ��ۜ�y�   $��������I���}����O��o����&�_y����շ|��f���~0'7K'���%N��21oL�+�\�C�I�yM����?�0���u��y�j��=>����t2���|�<M��&&Mǅ��EA���gQҡ��΍XK^ Gyk���ݿu��O]
�c�s4�6l769ME��o�z�7-�|a�uu�^��(����P7'&��;=��W=EYz;�񆬑�]�ٽ�,�▮_�\-O=�j8��"�=2Z��@{����N˒�}x�krW�Á�n�Z���AXz���P���5@�dC�䧖<�W�,t�G�
��}�k,�
#~OQO��8�� �0y)���R�`�w�gZ��P\&������ơ`��"��R_���
�D{�\�0��9�����=��Ms��y�ޱ�D�z~�u-��d���yG���O(��ޔ�]�B4Nr����X�.��i�K!���霫�Y��al�}��{��&���l�3u��"�9������P�Ee��{K��Iy�&�6%�\��X�n�q��8 �ʰ`��^��@�1Sk	�<@��c�1{�G{}KA0��0��TZ�����߇a�h��+Ϸ�8(�÷�#z�\�mRF���E���Q%K���7�9���8w9.ȼ�SW¯Q�)�(b�[lu{zeL꟢��kg\�D����1�����ł,?�z�Իɘ.J������(8�C��z�C<��ff}��#Y!�|*L%�*��3ŋ�*����~�-�C�^� ϣ��������%�@���~��yly�Gq;l5֏�Y��\��a-�*F��'�ǜ�P���F�	�V��|�>>��/�n�v�4�D_϶w3�R�,�S�,�����mAy`�1$��� �  F�i��J������7orfr����Vb�&�xg�
�Dϋʋ�F��]���IB����y»��{��j�a_z�B^|x_��W%��o����~4���+���x	J4�ڿn�[wy����7��o��3������{|�y�����?�,>�ǄA?
��=�ɤ�E*J�TӞU$�����Uzn�!�&3�YCN'��H}/�ΐ�O/}�mՏ<�ʄ��M7p	�^[BE�Kl�{�5�����l�\��]4�0p�(7��a}DⅢɍ^�� z<�vfZ
ߒ��(%f=Y�g�̱}����/u�zH�v��}��Ѝ&8ʄ�>Q��쉅�|2��2`��!p~ڣ�O��{�'5�����s&�HI�^��3?�n�k�邊�7;~O�@��n�u�n�[�2�˂�A:4�S6T��;K��Ǌ�zd߅�#QZ�W2�U1��zjw]w��	ݒ���aꎮ��ť�����.�N�;�;9GݼT.ʘ����f���_X�
�-M�/o�d�`%�:W�w-�4�_���ͽ�����݌����v�_7�{��j%�3,wx�QҸ�M�Ɍ@��Wq��:n��/�{���qx�iw�30
��+�7��h��P�FKjj2��B�|N�o˦l����M�{&�=�$	��b𪇑ړ\�����S����mW����bC�,�=�_f�֙�x�G�C»��3��L3]6o}�{��)��I� Gz5�h��(��A�M�T����ަu*=^ԡ�.�:DiEF09�+��Ϲ��<�ߺ��&mJV�G��H����.�4DI$u���p&��dE�6�Kf�tѱ��Q�R�ӎk��*�����4l�[� ��Q��%ԍ�/\TI��8�O�K��S��d5f���:�&V<��@��S�ҽ��Q���uJ��	�U�cs_my�o
�����=)y,�)߶���cY��XC�\uDuuٜef�h�Ӳ��A�������+(h".���П��[�#�F~�M�>
��-f��nb�Dzp6���3ެ����*�@� ��\:'��k։�R��P����z�dY>p�P�
J�qC���l\�Ru�:�3����y�Ð�DV4�.8�Q���`���^N�kj��k�x'����7|��I�t`��K������\~AnN-˴���w����ny}���RW�!�D�t)ِw�f�F� %hGS79C�N��5R�vЙ�X(�D[]���A�r��;}�7��<�w�[���w������]������]FCX;�.p��n�H��Ak��5�l�9f�o�)�g��=��.F�ݚ��l#[e�k<��Ur�Z������C�^�-ϵ�w�~�p��Ϯ�>̕�?8���k]��Jm�\�_�rr��3b���m�<�Md��R��x�p>�7�SHv��b8\V-����)$�2Ʃ�ʬ {��ۺ���;�+�wW^W�f��GZ�`1�]��H���G���.�HU���eyZ�Y���j�A��x�N��c�P�(֊�q�|����0y�����|�BwM��dx�K�����L+7=���1�ᩴ{�K�e�	�ʫ��f�ݟ�-���w��b���lt�n.'���v��5�?\�R@o�[��:�R����v�����^�D�����{N}��ʏTз���x��-&AF'����6�����mL��L��;�j�G�P���%/��ga���t�@�>�F�P%�!��1C�#� ��|M�^R�c�b� ���XQ1�H"�y<�Ϥ�k}���u]ظ4�����!ɖGNC�i���Y</�M��R��J��ld]G�H�9�Qa�n�h��<Fu�@^b�K�K�d�D��Z����ِٳE�  I-����c:���s�d5�M7rT�HɊƟ�/���y���s  u$�o��M:���t�{ l�3�Y&�-JA$9;l'	HcrF�:^�s�#Tq���2�1����+�|��5�~�N��5�
x�'�uf	'Qw�6�J�W����G3v�ˢao��0
��0�>M�=31&(ۻ��7�9�q*�[q~���x�7ڤ�#ɩ9u�̭G�E ���T}Wm�h��^�C�p�F����P�(�����n�ԣ���(���ȍ����־Μ9%u��񰀴f�8RF���!���m�$�.~�x k<L�ɽ���`�{��Y���ω��X�=ڡ�~�i3��릇�]��o�#�{f�6+(�%����.�ͱ\'`�:	L��j�A�j�g�����z���YR7�$e��\ T/��^z�Hd۔h��LV%7�<k)b����%�9�yMY�f�}���sJ[�f�L夎��(��Ԩ�<uq\�^2Oe8P6�|�{���.��p�cmNW�۰���iB�]x	m���<D�އ8��Fآ:�Eo��Q�g�v���>���w��w��-6m(0n�P�7s.��K�.��ܝ/�_=��ڻ�y�3.���H@��Y�O�]��Zd(ۼ�0�؞�:�;�}¸��#6����I�Y�9iFQ�s7��Kk�,P@�	��g�#DV�&5��K��r l�z]/c-]��;ʵ�|�x]>�Xe�im�R�,���I����LZ?
�I��{G%K�~�#K˻� @�(��U��V�P�0v/��cJ�"^�Ҽn��BC�$��S��]�=�D��ᦷ�'��s��yV�k�@"F���\���Z�d�Y'�AA�����Z�}����yG��@�6[;Z}O���R�e a�1xNԇ��J�`�|�z�V:9�N�f�|��1�;�x��oR�����.��J�k~�9S�ep���~�|uT���efl���H@e�����	��I$��P�\h�n:�G�)r��27�^�vA���moI֕];��vF'䗂�����N��2Ϧg
��T�"��=�[2�͛
�/'�^ؐ�s;V�۱ܥ�sP�&�ۨ����r�>�Z�sp�㝦	;���]�ww}$�N
�j�!㐽�у4��EZ��L�cg$�ʃo��z-�S����O�ӃYG��z��6���1�y���s���]���ovL�-����nm�^M�=�E�XG�ꅂ7�)^ICfaj$1�^�ꐫ��ܽ�)M�U����2���b�ɷ6IcwpP�b7�#Q��7�x�	��U�w}�,�f��n[S���w���v������V�3y�.l���f��+/�Sn���b���6k��{-^�.��H�,.�����"��.?m��캱���Ϟ�er������b�VǙJ�cy~+u#�8-�e�U�>�:�'۩��7c��`���9�H��7C���'@u�q25f˽�s�8�h��E��O��2�obY��CkS��q5c8�t�4����jf*Y�q�{Z"���;h�d_�>���[�(۶� ������{��:�,c1N�q��������7������qM��3f����{�2m�}��x.2��7(��:���Py$~�3�ʝ����f��Ϲ���W_ �;FJϭ�����D��(}� X;��T#	���xw���8 |��t4���q��\Y��_��Ikve��3���M?&w����{������w��s�'zn��O�M����a�߬>�\.���4�k�5c���=F�;�7S�E���o���M��o����'��o_���m�k�凂s�+5t��Oj����8�h�� w����)�ֈ�~}=�vzej�<�C ����p���ਜV�b�"zmU�:PW:弛�<��ۤ����f�k�_S<�es�`8Z�<�\o��]�g����xʼ�R�5�ѩ����)�a'�F���]�FrJ�i�٣r����t�\�������2j�3�ǏW(	u��F��u��i�6��JT�Q�*v�K��*�4F����g_l�; �y��:に�5_�'	��}~Q�u�Ȍ+R���[#@�=f��E^p}m������s,as7�-�Y" %�.��R�ս]�D��izHWWF� ���ޔ��P�/��YwYڊ����� 8�L-��i"B1su��1<K�:�ը;�����kx�5K�B���+:
{h��|z�]��V�@��ڴ���AA��Y-ٴ1�n�+o����ס,P�fI�\wºֵt��;s�*���kk���
n�:�:[E�4IA�&Z�&�a_J�̽���BQF�.қi$?e;:�-�Ue�%ebw���� sd�/�Q�j
�}�m}�:��*��U��0v��ę���Zn5���;'*��N�}d�.�{�B'��.T�ʕkj�Qv���}d��a<>V�cXX�Wv|�r�1�	��uxv/jIb�ý3'�Usnc�]�Z]�R*�!��t��I�N�׽E+�YԦ$0��g�KlnGz{0��ԇ%mB��+��h�I*�D�,�t���L�����A�K&��Q�F�v�i5�z=|��w=s�v���`,�>�dVKsxv�Y�S'���$��JQS��ZN��*�h�>�ܮ�o��W���FP
�*�,����䟟k�Ϳl��}���&@ƬS��x>e\2��+��)�/^���i@�D�����zc�{�'���>��Ȓ[ OfO�h7S}t��4�$�n��M8���v'p�ͥ�A�R:/�i�5��R;8���{	("�$yJ̚�5캪���C~G�
���iN��V��K0��z����_xWw��
�irglo/{�4ږ���o�<�<��ه)W�'���x�+h�4�Y�'���
���=�A69���T�*Θ�D����C�튋��#���J���M�=����4f����Y�lzz�p�~j2�~�e��d�+eu:�`����������J�#yάy�59 zh��p�����~<�2!�ijm��ȭ�	��C�Uq���z��d�3^�y�^���:*�oos���I��
��X�j3/�z��o�z���#��c4�^�XK;}۳c�S쁵%�%�
L���wL!h��@/ZU|�{&���e�T{rۢ�����Qf�����k��#=�88�1Ϥ�8��d�è��<��|���g��$���;��6s/hO����}��^&�x?Cإg���M�Q<j��R�q&Q6�~��&�r�5M	��Z�*ܮ~�tz�x��R~K���8)�*�VJY����{��(\�ics�cm"��>m&N`�'�V�򓗞�v�)S*5��W�ڕF��jGގj^4J��y�s�2�3v���t)�:�	��.G-y����N��|���'���J��7��eB9��^��8�p�������ʗ�^T�=>��3�d|7�W�KǼ՜^g~1B������XǸ]��
��z��ã�g���2�w��gF��@��x�!-Pn�sл�?t%dPRγ9c��;���(Eo�-�]]/I��� �R�2[ �ytD���Z��e����?��)O(�\�q{�=���������t�����.�˯B`������.�`�'����(Qw�d �2�S�R��^G��.>F_,I���K+U�5�ߥ8lc��:k�q���c{��`�.���06�Oqr�p	�4�h�*��ier)'Ho\�
ї�N,çy]��wX��/S,0խ�E��UjA%���̛�54Mȏ���~��r�k�9䓻�*l���um[d��g���3��<��d��m��m�	.�<�7n�ou<9N���Hn˨�mY&�mլ��yl� ѹio�#��dk,B �"?z��o2dv��/�$��vߓ�C=��=�X��K\����ܷg宜l��ʪ����$�2ʡ&K��mz�֯�wE<�3p����@�#&����y�8�;n}^��w�rry(c�k<����X*�+=m�y�w�6By>��w<��MN�uz��N^����㻉A�2z$�+�[�5r��0�Y� ����C�W�
���#����)1sjw��Y2����s�#�N	 �~�u�w�6�"%�6�4h���o�=�n���4l^��2�+9�K���z�b��3&��&�VIf�:��?�_�jh/��wNx����D��za\�v�����,/�?"J7�]Z�+DX�J���6O�x]u�{�n*\�Ng���g��)%���7���H,�[iм����`��	�Hk�gR�͓��z��IA*@�	(b)"K^��%!�{Q�����^od�F5�1Fb�w9�(X`�HnA���>j+_^V[��ƣ+�-1�Dgg�1�C�?' ���lQ�Q�f5Z"$�4 {<GJ��CC,G�i�*`��
���|���5c�S�R�����}���٪�(�UB2�1�;�"�s%:txP�k�<��H��oG�;�1��������*�J�]�W1wo;�P�W���yOǢ�\�+S�LV�x�0Y�
�-�S�
i�ֳ<�Ӌ��s�e�]M��=�Y�����	I�\�R6Q:7����$�HP5�8� ��f�k�۶���{J�	g'�'	tވ�5�G��h?Iz��>�K@y��U��
��UJ��=��7��[{���VM�P�8���&�+�!�-�G�kG8]z줠>��������?3�E
�A1���%�"�wFj�I%:H�=D�mX���ӹ���	ͷR�ӱe�{�3�r�5{JH����&t��Φ�:aQ���?oי��^V�ٚ���{�ۻZ�����L	��2��3F/�i�}j�&%.}I<%�n3��!��1��'x��oI'��<K��jv��Zp`B�͙��sv�t]I�F&I7�~��g�&"�e㰏V5�}�z� �&��J}��Q���[���^߅����k)E��^ű&�.Wy�Ϋ|A��"�M���&,ܗ�/�]�=Pp�4��k��I�G9��R!YB<ҋ�{j�!;U��&f��C��A�gAp��eȟU����.pL4��kKݪ����S�݇�����4ƽ��;M���z<b:|�w[��Y��������e�7������B3�[��NS����G��.�wi�=�蓠�K�~=�ͼ����C��`��u�;��lp8aK�o^���*��D޲A�Y)�ӯb���Z��[>5��6�t;�#D��X<�R��^gT��uO�%�~��˿]�A%A��t��rA�˛���{��4>L	'�J=DQ���Fݧ}��|4�������槀�N�_h�4�<�=�$�KT��P(R�Aų<T#{�cƇ��v��(�bƬƴ�Um��7]({��n�Z�_��rL�d�i1�m�_�!^��_H�Mg����T��u'���1�6T�G2��h���im��)r��ٓwlt�/m;IJX�Q�L*W�XP� ��ud��:� ���V�U-#^M��o=�<��4��_��0���	�w�6\��r{��҄��H�HF��_Ƀ�բ
��9�Y\����'���ZG�-)6ucڏ)����6Kh�e�/"e3��r�o��Ȕz���^�T�w���vg��P[f; ��=z�QFaƦ8!�>�Q�B��A���T�	���Y�/g��,�:%[�~��]�V�^��G3��d�,��H"#��YM�=��k�ԻSۻY�X�GXץ�I�<��d3w�ֹ�ܮ�O�������t�Rv
c�Z��=T����cU�PL7ʚ�j�.O��rBm郸��1���.�	����n�^��1��Bg7���y�E�PD
8��D�}������QU���o���yB��8#�����v�F���e��/�ẇ\`�F�?26~��`�{�˹,͖f���̶�������7ov��×�"6�F7�ػ6�8*T 'c8wM=|�,Q�T��(��zi���Ó�V�����h��04F�p���B0Q�XP�f�Q~7M��htPY�3y��\o����3j�V�b�zp�N�%+�&�ł7U�s�&�UW~U���n���Z9�rf�$���~�ِ��Ej��\hq����o����k�s7�7>�����)��(��7 �s�v&)}��Z��E5�4�1�7�>�ۓ�x�};CرDʖ6׷���X�Ɏ��&|��Gܐ�1��X&,�:y�#���x�~ś~�p�����k�B���b��2�`�|{:�f�\�(f�η
��{K�����śZ��t֑ºʡ�}0b �}u<xHj}��t��G�M��߻�b���rk}��I����{���5%b��ҁ�xi�_.��*�2ijW��Ɠ��)�I����f\���\�:�y�S��ے^�`=w��>��_s���gi�nEY%��mM6֢�]��M�I$�h#��D�+5߻�<��m;���KY&1en�C$���]�5|���/� 	#tn���|߻�����;���;��}����7���sZ�`'�l�/.&���ů�q��W ��ȿa�t��Q�~�mX�kD��ܳ��Ӟ��sC�)?Om(|?� ��o#����Y�O�,��=11�lٍ� ���<�)]�0�$�"(o}����O9a6*�{�w��l��/9������d����p�C��^����(v���׶�}Td2��.���xp]�f}^�U��Έ��:����/�I~q�����o��Ht��E쫘iUuñ
��m/cj}�Py,�lF=���o���9���œ����E���̥=ҷg�j���_d�G���¾!»V<-�\ 9-�B��/��f�*C�2�R�����1��\�ZXb�>}�̩�G(�f��f�J̽�fυ@q��8D�x{��a�-ׄR6�`��F�wÄf�Qv��x����d ��(E�>�M�������b�6�T�.z���^�hF�?9I��Ԣ���|�h3	`b�o�e�`L8r�H��l�����>W�Z��w�l���cU�c�?s��Ս�c�M�^�a�y�w:ŉt���Iw
�)�:��w��s�h��۫�J0��E��Q�{��v��r^�KH��^���h(}&6xH�����
��X�=�1��n���v:[��MȂ�������z��گ�J0Y�d�E��;��q�i���*�T�5n��|�_ug��ꗑU�����o����v��G�+��v���wY>je��s�m����ZW|*M�)k^�����jt�ٮ����E�j3ܚ{�F,����[�<���t^^�M����g�v\���w�o�xqV{�vr|s}^ez��֯�k���P�rg���u�th��@I_Y(�RM7���J����
/�Ǥ�)����	L�
�Եz�y,�9TO����}W����S7-�N���`��4Px���E|
=�[��}}�X�>ٿ:��鈧9@/A�=У�޳��c���=��ᇌ�6���� ���%�>]z�Ve{$Wg8���h<�UD��=��w G�u~V��i�{W����)�b�0���v�v.��M�HKYVW�Q��s��-!׏�j>���b�Z�ܨn��t�����K�r�xw��;]N�u�yq�>��3���o��a{øTY��N�>���1xD��s�C�,���Z_X��]����P~�t���BKӴ�z�d�6�]��k�w�I���jH^���ɾ��N��R�8Ѧy�a2LT��_#�{w�����vy��=�ەb�j7��x�������;I6�ji���'Awf]E�d�P׾����7��z�1
q*�f�U�L�:��ם�8|��;ޝ0ξ�缋�׸w�lJg�u+&^}Cғ�K��x��LG�5��[�Uކ����Srǅ�k��k��}�I�C���t���v�}�و��6Y�1[.�kף�a�GU\_�\{s�;���<���γ:��}�5''��E��|���s*�ey��e^i��4����g�9���e�V��N].�"ǳp�M��uS�[/�>�J$*t�3�.<��m�(���_S{ê^fOL�����D�9��wV��(��,�����'$�%�t��`�K�Z��z�(�*�Y�	݊c��۠��4#�ven�y��K����2�.�h�gm�#:��a��W����s|��g�����6�߯�j3?GQ�pc�o�K��]���}֠�60t�¶xJ>bv�#�8�I�ԑ�?}�x�ɗķ�@�c�=�'C�ۥ��Ч�"�����d���;�ŗ�Yzn�q�h>���V��%�nOON+�\+ffmLWu�@�>�k�wg?��~:�c~B!���bR�i�r+ �{/g�����oٓ�n�����Iav�Y��dw�غ�<w�����v���6/���gi�2=r:wc=��tn����a��!�r����	��6�cT����J�H�zr&���]����v�R�蛋��^�~�OA��yM�U�3�#ֆ4d�))����1�z�y�ֽ���ڮ޻����=���K�o0�4΃��fخ�0�[J7�d�p��b~�ه�@s�=P.��h#���$7��S�	!,�	�b,�D#V�v�LŮ8�ݩZ,+:9G��h�,n�r�ƺJ��T�؃Պ�-T����jj���Ʒ�F�jǦHpv��&����I�Ů�ۑ�l�2�ޓ�{����m�;.�*�G(�L:ˇ�3D䭥�J�k2W3%�S�ڂ��lɪ���6�b�[׹����ӥ>ړd�0�"��T������۬��{&��ѣ9a�~G��Xa�wp�/v����j���(56�u����X�� �u^rэ�;y�HH$�Z���e.I��ce�9�\�k)�l m�ݓ�'V$�Lgo���v2����\��-�h��c�֖��E���:���ƕ�ϻ�Y�r��{��:���f\�������J�'����`3	�v�c��;��9O��}
���4$(u��6��|\ЭW������2hh��]ӥ�`�1���m浉�ă��=:����n(�猰�{�-��t<ج7����'�,���7���H�s��L))���[x3y�;
1�R�j���(C�dK 7EG��;{��r�o&�r8ȮeJܬ�l��̓v���W̨�a��h������x4�;Y����Y���(V�N!�.�e�:�h;^i���е�z��J�{G�_��6dA�3J?m�Iu��u.<��Y𞷳U��$��D3�J�7�m���W'��1rܝ�ן����	v��3� !���� 
��d�6R7������wF�����ud9���v���\&�s�[�-�$��Y��9��V��f_:4�W;����D���A�h f�؈�D��� �V.� �ڶ���m (-�d&�*[��"�7-���d���e�b�-��\�&˶�-�Qc�\�T� ܭY��X�m�Kv�  +@! h�` �h�d��me�d�]Y0$�u��=y�y=w��7����;�Nd�@�M������F�������]��\,��֕٤Y���a�z���睽}ϯ�s�}�sgK�cl�c6I*$�Ʈ�K�n�m�-� (Q��	�Ki����n�������u�n�E�ST�i�{�R������F��{s�����N�;ۓ�S0�+����+�����'<Ȧ,f�����D m�           �bQ&�m$�m�m�Vƛg�Ϸ�m�,��P�3"m�.v{�LB�l�i"���h�5ԏe\Tݒ����
DVel@P����
�E����n,(+��<�á�8���;ï���\��'7x�
̘!���d���.��w�4���6:i����e9��[�����+��O�[�/�q�\?c߾�'~߹痎�l�%MRH���˦]��%F�� �3SMo'�������%n�7d?�ȑm�[��~����>�vf�s�@ -�����_Gw�Ns��;*�o.�	Ј	$cT�A� RiFcD�&����E��3eZ=Y����о���zSͨ���J\��/ۻ;6��y�`�g���uq��ћd���)/�)^�)gx}+�6����{7S��q��&�~�����;_{/?x��;G�Y��q�?a�͚{�jd�]��|�3�c���Uc7���5�끦�2�%�{w"}���>�{�l�N����m��O~�Gg�������3y}QQ�JAO�F���`��5,��f&���E��.������v%��Ʋ�'U�UY��15������o�Q���謝&�G<�����V�r�m��Ӟ8&���<�uj�MOvf{�݁N7W^(p�����gVP%��~@$�(�Bm'������!z9\(��o\���.?8i?�a��}�_�ٝ�۽h�����3 p��}�D���OB'���h}팳�h�i�<�2c(T�/h8���{)<�a(��x�f����(�͉iu���E�cx;���H��'M��aƵ3��ק8wvA|�ԫ������uoM*��cu����s��=:w�:�j�ϩ_�y~!x����#BW�����GF	�{�}X"����\c�nxQ��D��٬G����{��GL���_����пNG�R81Vwޞ����W�3|��Dl��|��������jR�(��ʗNܺ�';�7~ɴ�=��*��f*Vzdy�'�]��=Qj�3[��o��ɲ���L�d�z��8|j�uӾ�/j�6���:jw���'^~=߱ߛ�f�d�Fq�ݶH��nS�J,P�Ξ��e_��4v[¾~�}=�{��/�����{�Ĉ�2���~\�7dV�p��c����v�3;��z2�������V��]
�-z�p���M��K�dS�ޓ۾�z�uN�dݩ�[>)��0�xRD'�ڵ����#"��ĢT��4�2��.ذ8C�8z��d���֝u������l��SXRO;\�N�T\��b�]�������fv��:��u��gn���x�\jp����Gxik�i�/�5us�K�yFxXΛ���kώO��vH	���Ve0�vC̫1��p�ߠvf*6mY�����4�_�l-~�yZ.B��O^'�qҩou(��g��R_�E\z���P�����&�:�
��9:(9����멀�*����pfdȫN}@��v���k/��w�����(�+s�b/{"ZD�� &�)!��ȱ��n]������r����3�>>��/�E\��$�Ӳf�;_����"��·>�#�x�|����G�|"[��Áվ�j��'<s�76��~����OeD�ȥ-?z����EƖ�|o,}uf9M=�؜�x��_�Vh � zd�W�ޚ��{$����R��JW��	͓���r�{l:�QC"Um[�%o��lT�21�" �R7�}Mzw)�{(��s�ե5n������w��_'�����f�ý�����݁�K{�V�&��Ql�o0 �Z}P#vR�66챻�g�j��b���1�{��g*y��<m�f>я�h|��S��/��ZU���oZ��cq��uG��Xw�~\k�j�B�*~	����c���܄4�-���}��tN%7�����x|f��pG�'�M�cLʲ�y�B��E��ֵ��wuK����Ͻ�;�쳃��ޟk���3,+���=�*&W{$7/�9a�D��e�.�nQ#0����*/h�G?{򵹂�eE #�$���*G3hRC'�KۏO��Ξ��{r(�z
�\�s�H�_0r+�隡�|�v߶��v2�آd��Z1�k��j����gkt��݂N�6�K^ۙ�tN���������~���fF/�o�gޠ�n��:�',�������^W���FO�ǁ����j����rck���T���_�÷�ZW��huH����~�4��.�cS�ß'k�&�h�G��#�\�`����Nn��W��������߬�{Ѯ��P�r��]��j��W7F�:��Mz�<W�z21	F���7n�Q5T{:>�
��Y��\�v�F4��xm޷��-77f�<��/�ߥ���W����-��ݙ�ݒ[�dn�jh(���t�n�w9�}���}���'����ݥ�$�Em��͞>��^��� �"}�Y�;�����w/�6ju���PI�%ـ�V&RD	�m����N������%�|k�]������y�\y��ϭ���Mz�ӟv�8�}3���s��~��d *��{ه&����P��7/������3b�׏�zw�twv��.�tn�=��,�6�JB�ݹ����_I�;B���f!w}��_�"{�[�~��Jذ�^� �Uϛ��p����*UtH����Tt�"T���;�]3*r�IT�5���_�6��>v�4:���������mZ��y��cfsB��[��Y��(�v܋�
Ηr+\n䅁n�*]�5�I���G
`������n��$ϻ��=y��b���[2�;n�W���=��2nv�6�n�6]��K�g�R��5֦��" N��*�u��X_Z����	EA�Jf���:	��~U���O}�~��K��+��ќI���T�/`�­����5ò�Ow�w<B��VSM�S2������v���G]��XP{��s��qͤ�3�BtV�������x5�(5č��2|E���+��(��<��j#��ќ��[��]����gT.�$e�M�E�*H����7�uʻ�a=t|7��?hT��6���ᳵ0:=g�4�][��{;�M��mP���������n�u�����{��ͩJ�u�ﰧ@g�Q�8�ƓN�9^쮉�>��r��3Z6��ϦӅ�#�U�g��6:�xk�Oc���p�f|�/�������~C��� !4����5�o�=:D.�}����ѠE���S���G��|\���yV&K��mZ�$�"����� ]�+&��]�χ)�4́:�yS�����P����NfD��7�޻�[F�s&{$>��cc�.ޘ�}[>��=��L��w���������J�}ӱy`�����7$L���ݫ���Z�Y��-��'�6%��F�	�����T���o�z�,�S���t�Vp�:F������������r���{�/��_Fm�$��X1Ro���eاx(6�|�ܱv6�sYݗ��U/���Ѯ\�i�9��q$�+ =W��/��mmv���ԹW�w=�}��TZ�H�u��J���H�����f�Iŀ�5U(gb�sTC�}�j��w��tk�)Wu��W�y��������@�_E�a��g��f�w1�u]}�5�ό��\��7�G��.�g�l<�z�{$F_�mC�{��ۻ���I��kf6�!$KZ�`8��	��U[*��dmTy�Zt��Ev���P�/����+��{z�}1�*�ޭy�
�z'j�<���e{p%|�{?��w����f��}��S԰z����W�6Rž�','�TQ��e^�F`��a<Y��M׵�~m{dϙ]h_@��{*�X�5���>�q��Wձ�;s����u�w�0�t� A��b7�zjtqSuU��O(e��;!N�%�Fe>��������\�-�o��gQN�9id3��;�l��\��GF��mZ.��R�#T�)����*���޻��-�N������vYl�z�C�G� �	]���7��\/��S��mn�'��'g$zN�-9x���]�]0s@�r���Wy��G��^2x��#/#��	q��)v�+�����oo��k�5;�׋���H�̐�Pʓ�ӝ�(���6N#�_�?�_<�;u���w's��e�����z7-�}����a�ǷLn���at��e���hQCoz�6������{l}qRrw����<�gI�>t9�xG�`z�5�'*T�:j��9ڶ�`�����f�7�F+����.j`-�]tF��ڇ�1��LM�M@�v�'�m?�%�ݾ��0���NU����f��&���Щ���P�zbq(R�^�:����އ;��l;��V���I�G�^�PWo�ڔ�--?o�کJ��^��<��>Lo	��N�eO^��[	��l��xq׹�YJ��r�'&��~�w�������}�wh_d<�?,�ʭ��('='��@ݠ�x{Q��/r��<�^�Kڱ���ux;�kyL~ѥ]Zb�쾘�m�&�5�doB�r���^q;Y<��H$�m��m�����Yj�b�� � �bkw<��߹}��[���s�dd�Ԛ�Il��ef���ϳ����7�%  F�[k��z����X4^�.H�V�Er�&2U�Ъ�&+m�WKt��`���ѝ��en�+��XsB��F�p#��������;da�>��0�޲z`�q5��!����Zs�^���߫�_�n�$Ul�[-��7�o@����o��ϗ;9�oA���ds7��_܈u�{kƇ�5�ҷݜ�й�y���S�TVeR�?�U��3�%f	��m�J�����[��U�ك��Q��.��{��n_��b�F]ӽ���ӝ7��7ё�}!ǻќf�ʙ��k�/�V��'��
�����g�3f�S�Bv.�;9�&2��l�XM�l�dm9O���:gGJ�2&��Ӌ�=z�S�{x��wn�M�s˖U��b�_vY�*Y��~�����gwӮ`���(�;~���!ٸ.vӊ&&Lu�$�������2�����u�<��jmcp�{��\�Y�`׭�{��b��<��ʕ��V�9	�;�5��_;�^u�h����++�Ֆd��Օ��Y�������:�bZ�9�'ն���٢� Toq��n�R�� �J_�o��{��r_�����Flջ����i��V>϶�:�f��i�p��9K}�.���K��GC�/L��'Z|��f�rU�8Uw5���-����ޗ:.t�W�T�m�����wkLN�NE蹤k��~Cz���t�����x��jp�9�p�m�7�l�7} �oe����v�W֪���V�~^���88+�ê}��]o�����c��_�N��ui8�7�L�l��y*Q%��e&�����b7��|/��Q��Q�ʴt�_���Z��^͊��{����]�ؘ��k>�\ӻ�쭯�:��6���3��'v�S=ٷW>���Iϸ�{>����̙�-�y��k�\�'y~Sq����L�W��p����<֡�8!kmT�_L+ݣ�/o8꧛c��ۿk�+9ɶ{�̕���5(�Et��M�z]�Hf��n������m��z�U�t��^).��Z�-��sS�m=���K��PW V�F�bL6[��[tѩD� 8R
��{q��\��pʼq��rRܫ�m�e5I�b�:S1���/f�M���h�� �=�!c=]�6�H"w/$�S5f�fd�����:��;�9$X�}xpf�c��M��.�����={sjڳ�!��'��OS��������t�v��u~MDSN��ٱZ��s��r�;/k|բ��]�m�pnl[Z{E޼�L�Vǻ� �E� �M�s�'=5�y�7s/��<�ݬ�����[w� "(J�5s7���y�g�VI&{�!�2Y���G��Ǉ�ݦ<6&w�a�BG{n {����i��q��a�m���z>�H=3��vw=�3��%@Xx��,�޳�=�[oH�f�� �^�����d1�l$-޹�:��:�!.�֤ǹi	�5{Ns�Vޝ޹�q���zn�m����@��OY�=ˌ	��@���;N�G�� <���@��O~����
��	7��^�@'�����<þq/6I'_@��I�)�ɜ�|���~� G8/��d�&<`L z����Z�*U�^�����bR�,��L���z=���;5�{���I
�m�	�	h]�I�[༃m�Ѵl�%�-�{�������tS0l�qy�;�q�U��!�^��3�S���0z�m�^ wM�I�B)l�x�t�R�	�[	�u�i���w!��z�	;�s���]�6��^ѭ#D2��+Q_^)j���ۺ�5(Mo5���#l��5�q<jemq8 ^�n�����CI}v"� T'�w9���@�|qc�%7�b�˺�B��Y6BCK]�>ҶI���U�miwҺ�sW}��s�n�/����l�l.���J��v����Kul��F$�ڷ�]'|w.\�#ϯ�|�Q�΂S7y5�˭B�8rԵ��i�<����9Yg���uֲou�W;kx� @�,DVc�ǍȖ�o��>7�es��f�Y�x |���MF�_Vy'�����P99�U���L*�Bq>��a�̦��jZM�b���JV��Y6��łh�ǐ�x3��4`�(C6��q�]3E:��:��t!�-��wx����w�>�e���D)�6:'���v�ٜ���I)��<�A/�|���{����N�*&���t2Cwۂ$yAt��1���;q�rr��OE'��8�5o��־��0��C��ݫn����Q��
qޛ�Գ�ʴ�]�E�,a8��u�v���`���K�_	*��m�ս�k9>��/ђz�d�:o�Xv���	��������g�C��������L�{%{(�irUW�6��k���O���^���5	D��ƗfॸG�X�l�;���%g�^�N.��������m��Lڑz��x{��M�I���}w�2-)���.����o�me�7L��8ْg7�oׂ
[T�d�U�F��\��Ϸ��g��e-�}���z�������ǩyD՜��Y9���w�(AX�N+I~�Ìe�a���1�|���jؙ�߂���N���ܺ(���F�g��	w.��D�]}�y1��}�����s�}�134�}���#�y��~i��y����d���z'P��]=}�q�b��@����������ޟ>���C��_4�2�:���v�9Àޅ���3�8��{�\����2Qp��n��O�����֨ѣ��0J�m��	g��ԫ��fG;�h٨:�V-}ݧ�n�'���Vf.��{��]rNx�r���$V!UJׁf~u�����@X���W�U콳]�m�zŃg'7v�9�?fIj:�Oy�3�wj��t^[6��\m�<�͉'�$�D��ۿ��}���>w|����o["���5GW�'���-׆�#�����[���^Ӹg�2��1<��4Jf\�Օ\�M�oo]��,�C�_��p�;���0�*�����r���9�������kg��<��VT.(�{�
���c����W*����Q���f���tUج���M�[+b�e� k{LC\�-����'����
v������zKX��������<(j�z����ٹ��s=�ewl�=�&��/G�H\%�;�u���y�v�0�u��o݆oϗN�C��V��]��eK�S�b�;��{v��$#h?p������7^��YUx]ˍ+�S5��C�Z�t�=,ѷX7s�9��6�S۰��:,���20Ck��0��F&���Al��n�Z��#8.��KR4�Sj�ّ�6�T �d�m�~�y�߾�'��}�bȓi7r*Y�mi����z��m� l��.�d�9���OnG{�cGfs�K�M�[�r㚼ϫ��#3��vP���t�����s����mq���i��շ꛼vj�E�J*/��z�n��0��ߜ���F�����7���X)>���"^rc/�*zln���6��G��wj�h=���^�1j��+����{v�3�~�:�}�H�z�J�Ppdm*ި�=���=��{�SuW9��=�t722;���n�:)ƪ�KF6������A=�r�n[���	���l����{�g�nO)��h�?%UӞ~�BS�#=����Zנ>��:�YQY���%���s}TL�ű�����~��G�܊HQ�����3�,��8<���m�����KB�i��!	6�'W��>�o�����-l�f<��S	g���}Z㑩���S��i����{��(�kzAPo;�����Ծ�Ez�j����}c=�lu�'@����6|m��%n�����U�v1�'3�R骳L���1�g[������)��V�:��l4N�C��u=�\4Ffs%������Q���9RhV�V�;T�Uik:zJ�#�
��Ǚ�b�t���=2b\��G�8�yK�/~L��*�<�_��s����yx�=S��<�?G�y��6V�3؞ �o����]%>�R��U{ФwE���Kg=䔤�32���"�����-�(B> �.��ʤ�^�˞L)ou�Ά�*3$��L�����ݿV��9]�<�=a��+2�-b}�wMGA���sV�*Z,w�g�}��vΥ~�TB�v x惊�>�w�[��Y��.��r=*Und�����=0�p��{7F�=�K�R`0TKޖ. ���y���rP��.�D����c�XxVu�p���Fg�s&�*�W���iFߪ���u4�Tt�U×����8���-�ηn�]灜�c�<������<­v����?_���cҩ�cK��S���u����	'�{óݎp8z#��E�T��E����yzw���#bc'C����$�-69����n��jv\�����\�.:���i� +a&�k�BܼңY�x+��\rT�6�� e�]�ŏ�^��.���0�]��w���㞰{��~�^z��o�e~��}���Y�4��*�''�^H<��ny���O6��g�z5�[���8�>k���>��.�7Ս91��"�P�ɽ>�ڹc.%�K���u����dya
b������W�����V�oJ����Fn�V������m-��Շ�<�+��H�e���v�b������k�����>��m����{Y�׫���������xGc��s�Ԓ=��C�9��~�|,6**un�=1��Ui9[X���j,�eI^��WLX��KF�<L���a������|#�actQvzǣ���O�^���}5��l@�6�q|3~�Mg�yEv�ݙWb�+s܇�Ͼ�jE�k�F�-��9���g�Ԕi˦MTH��u �zw*�F�v�X��T�:
���g�����EB.iƫu�.9o��i�d��Ӫ�~9����l�9������Lt���/�,�-O�DM��w7�6n�]��Jȇw>|� �%�0u�ux��E����/��y�F�h�w�4{��Ą�>���;&`y$;!�c��I����}�.�z�9]n����}�}W>�����Y3���jU=7��;��/��3�M��L�6D�&O����^￻����������?�Ƒ�y�S��SV!��}��V���M���)�ʷ>_$�����PQ��߉]��{c�F��q���/��Q#���_c}��;�0�f�N�V��8nxwmym�nEd|1� 5;[���1�t񜩿�37_�
�X����۠�=*g��k�F�ދ����7��9��qؘ͍���_�eI��&(��(���_;u���s���{�Ca��vC��~*=��`d���S5��fx����g׾���J���;���º��H�{�Nz7�V�Y������L��++�=>v�mt��Y蜇�9N?%�V�R��9�ћ�0g�яje`��(UO!sy��Ɇ�.g��)d@F�pOl�� �Y�X��s�d)�dt!޸�v��n�Grs��1����P�����X���KR�DP#-B�sMZ������ l�X��[�r?~��l���U6ʹnjn�r�����~�mq<��<�� D��n�C�-�\���z�	��ݫ�O.�w|ݶ����o�"����nW謉ӥY�m]���gx^V�C�v*�	�͏S�=}��#�b�MlIiWz0��a�{����##]���l�}Y�����:�r��s_<�eW�2�.:��>�Wp߯8�2���=�rA�c����#��w�w�]�PO����$}W}������C�=�u\��S\NuF���־�;<���f�uE@�E����.W��؎j�\��2|I����k�o��ڧ�ڹ�g`�X�w�ßW�[��y����G�R�QϺq��C�C�ؕ�/N��ӽ���24�gnvn�bU5�?x�z�X2�ƽCu���qs��$Ӆ9��V�I��IpP�d]X������.���}?}�N�6z?G����]�te�b=q�
=���w�͙�z�ҩ��5z'���{��A�l�
|3�b��z9���(OҼ:����%)d�ź��VǮ�1ed�˧��Zn+�0�XW\x�"�������2^�Ū��p!tGU�5�[U��B��w��w:%����z��g+�]��c����NNQ\��R'д�AY�1�ࣶ:ga���j�����,���.��w'��y�z����7z�M��f:��ogX[�!u\K�)��/W�ӷ�9�s���e}���xG�Ӆ�>=���J�����^T�#nk�:c&-�u�!Χ�L��{�%r/�	!�)6g<<���|ڷp�X}c]��w_�����M�Y�e���WLN����ڹo����N���k��w���yػ��f�Rث�q��%�v�BM5��[�Y^�}�����3uWW.�=�9��g;����ת�y���o��N���T8lt{rw��:��+n����X��6�3��[�o�ݭ3B��Sz�r�J�l^���X�������;��+��·<`ʺ��R�K�n��8�D��u�^�ӳ����dM��'���]ɾ��{7f�f�ҩ�}�hg5I��$�ѭ�U�k�.J[�����Jт2���{4��˲ul�u��n�Y��-�QRM�tF�G����x}�}7�0v,v&�o{��k����=|�#�0[[{VqD�<=�ڟz���+�,H����7¨ϠCJT�b��l�����'���Ʞ
c��.��p��������aTOMeO+�e��ξ���.Q�]��e����w��Y���P /[pPI3�8&���M��Ҳ�6�\c���)��zm��f�0t���'$k����t�ڿ�4pZ�,u��o��t,�@�i	9��Q>8��z5�{�.�s�t�u;ѓ�OT�)��u��L6��z�<���T������>����P*�Ӹf&4@��&[�ح�k�ck��/j���K&���1_���(ٳI�}Υ~@e���}0�ȯ}�YǄȾ��/Qj��aY}E�B�]v�͵���x��a�/�a^��'�_��h9�^jٙ=g�;׶e�Ӊ*���Ee&
IU��D�T����Y	�q�;
.ov�	�vZR�.o���ʚ/��-^Wn�an������K���;v�Aj��q���<}au<����t�@��!ٶ�9ﻌ���\Ι��=����/zR��,hj'.��˺ف�de��G��y����&H��M���k��;�T:����>G�b́�]A>ܛ��oz>��{ӹ��+2�d��S��������o�yD'vot���N�b�ˆ��y�^�DE{!�0�È�{�������a���6$J-�����=�Y+wT���u
���r���ulHdcď\��`)?03h�p�Z�]�WЪ�6V\��.�ŭ�{\��7t&�at�~F�慨�_�6�W��{�8$��ٝ+��&%����=��O���i�{�^�U�&�!:���f���鸷�3�;��Q��=�/G����*�c}��>������^a�^mS��B<��˭����WNZ6�x��X�Ѓ�h�T]��F��]�b�n�m����c��ԳZ��{v8G{��>49�Cu�wJ�2:�4�`�Q\C/�G��>�Ef湻ʱ�vh���B�Hq�W	,�	�Vę҆��0����&.��NPݾ���k��d��/���K������Fp��w�nG��Y�:��m�5CcIPp��V=&��w�^c1�ι������yvޗG+�y��)�vh�R!|�F,\fh�ev��]W��e���&�Y�qS�xLr��=�;s�w�ө�s}�c��'�f������V3�GIN�hܔ: ��D��չ�
�o�S���b�c�)�kfK.P�>rڤ;���`Jҋ(�p!����u:����z mu���1�0�Ƕ$h�f�t:L�ߨ�o([��*������ ��9�,���v��s%X��:� ٕ٩�b���(�^2�֊��{��h:漮2��.�:�ɊQE�[�Uށ5��KC��w��D�׼ %�(�͹c9up�Ø]�t]�U��kw5\=�q���ɢm�j#+�p�u��51�9�bv�gtK*�i�;M <lb�G�iqĖ�iU�h�c�f��j�9}}��.;�F��7e�c9<z�M�6�d�틧,�pc�]KΗ�l��Q���j1���\yL�v��۷�X��A�o��9�=Ī�i�7���ҫUཛQ'��9�Y�`�[�k�6mjFE���f�2b�gq�G%�S�Ԍ [�:˭�Z���:�s'�-%V�dM
��y0<1��p�Ǝ�e;��#����-�"�N�n��k��� �=v��h����˰c��gs���=N^˹��o�2g7������j�5�-�-��mݠdPZEP �-�Km�m����\�6�74`�e�J�j�*���m�)�X�ݖųem�l[��Km��  �m�ۗ%سrm0�-im�@( 0ZE��&��.[E��-�Ah�4P0�l9���B��9��Z�QXt0���.�̛�Ւ��.uz�̤ 2ڶ�r��6H��9�P��k�ܣ��bc���}N����w��9KiPd$�$M��٫3r3f��]�A���m�n�Ͷ@ �"�Zػ$e�l�$n��ٹ2�O��ڷkdJ�����y��U-=`�������H�x+y��[�����;Y,�,&�I$�	 m���v�V�$�@         m[l��%�$P .�@�j�=��<��WR��VN��ȁ$���:����!�2�����^�z�|�`��G�b�Ρ��3eA��F՝��Ρ�yMRh���?m��dw�������n��|�i$@*�J3�']�mH�s����Pg�����ණ{�����O�Ӆ�9B��õ��y#��#�ܽݶ�s�}�[2O��K"�jڻ2�-�df�cwE`���Ykw߹߾�}��������/���6�l��fIV�fL����rw�j�   ����ϾK�3�߼z�����y���o��Z�܃�u?��A����}�Ù�w����huC?�@�㴚C9�/�ň\�X�����267/��?{N슭�XHZW�kS쳗�@[:�_���{�4��}�g8�r����vj|ꧫ�P��um��dP���E9l��e,�B]��>�������{��n��F���B���;�P�s����tlI�yD�٥u�(�/Z6���r��pE��~��v��]�Q�wM������?�N�TͭPW�׉J�D�����-�	=���]kbTC�3��k�Ҧ�n��7��%y�.����~;:��7i�V3�x��O�4�{=�g; ��������$��s�^U�˲�Dm�����w���9��ۛ�2�B�9��ex,v��y^S7ܲx���Cu��eo>^�t��}�B��u�ټ��c2�cN�	?d���8H����)�"v�w�d�e��������s�-J���/�iނ�.j��I���[�<�y̢�K�ت�\V{F��{tŷWa&�ٙ���������������q��S�I���_�J���ٟ0���
5�_��͋;n?�}�?�Fyr7P���FON�i��U��;�=[��k��z�b�*��H3���;֚��Ië7�[4t�J�S��+k�Fp畨��=ơ�������>g�v��nx���٨��-����Y�����
��۰+/^���n^�{�^��|0��2�~�<�w���x�u_d�����#6�#6�m����sy/p�W��D/����t[8�{���Խ������*��O�e�n�C����5���!�W�+��'R��q�N����=��r)��
+�ߕ����!�P�i���w6� _�'Iw�z��gk�l[ӳ��}��9��y�`�T'���W�<������lm���m�ǰu�6;;�V���`Xz9�'=�H��wu���[|$PNp���ȗ �]���*�A����@سȻ�#��쬆����J��YpT��X9*����ofD���'z���8�TDpt��LO�WK�Wg��v�k�\/"�P4�{{���{�u�jAv�zs�gy�8��S1V=ک������WM���1�^T�����y[���!r�=�q�tgo���z��soG7����An;���:)Q;y������r]����￷���[xq��S��F�>�!P�p����~�]w�ԣS�o���>�]0����n�;+n�=��C�{�Ũ#k���Rv7�fa����ϼ/��,~}�����
>zﲺ��SF�|҉�}[b4]}�]й�X,/������'��iiK[��ݿ)W��J���Й�q쨯Gq��0ޠ��sxN�,[�mn�c'�}�{�O��ڜ�5�8��r����_h�2��}^F�-��*,�!a"�+��ۀK�a!˳+b1Ұk%S�.�(��:�<-�:k+rƍ�����:в>���޻"�I���;{��M<�-�-�8��e^��:`ǫ��
2����ޔ��A�����9Ǭ�J������X��:�������݃�K����߼��H����y��Z���F�ܑT��q����im��J���t�xv3]y�w�p�����)+)jS޼��X��k�'�x9�y?�����i鹡^��^��>�Oٓ��;��&8�%��̉Tƭ��м&��MQ��[0�y��=�սay�g�l����پ�al��Jeu�ߞ,�#��s�h-S�m�s��p�����s�k2}�s�o�
�k]'۞�t �&�ng�J��^>��ώct�w�3A���h?+ȩ�ն����-	�Hb��vח�9Wp����L%����s��h����{uZ�b��B{��˲�t�Y�tr��o<���x���������k�.��V+G�ȩ� r\ؗ�;����Ҵ���}.�{��T��Ɵp�2�i��ic10��NޱqX7�/��j#i$��BȦ�B��	���3t�@�1�J�Q}�֥�+Qȍ.�h'H�ZI�	C�ry���d�w�m� m�mj�[����gbΨ��ӹC,�.�j%�:Z.7���0bb��"솻����Cʫ�v��_�*�fN3w��5ۚ�o��G�,�q��8�������84M_�?y��8{l��$w�7�O����}�/{r� �ڴ������+�1�Wb��u��ؙ���G��{��l$�Y�7�½�l`�qW�d/=���u�� s�Z�vX&�š�=�|&�ao����uM���ܻ��m�-�ys��\9�a]
,��LYqz�����Z��,��O|�mO:>��w�A�ZQ��߷����{���PN�u3���ٵ��oʵv��~=I	9��TMQUZ���u��쫌��W�\k�w0vg�;��io�?w���$���0���u3s�w�'~s�Χ�>����߯����'��]o�X�<fL�zʭ=�����>;�+iQ��n[6�Uָ,�iT�n��j�����id�i\}o�M�]iv��u'N�-dYKJS�՜�M�RT��	]�,Q��
A���w�B#ǚ69�{qS�NVGF�Du������V��8w�+�\z��@om��9nb�@�ދ����}��~^ƾ9���� �e
"7�w�3ݦ�����ՑY��"�k��׈8\�8r���,_O��9a�/]�0^��� �}��4�ʊ��w:�n�{�e�d竳w���������r�6?u�į\���.��cw�{�1u�HĲDU�����z�X9���о�x�`c��
i����z���^�ꀺN��8��ʡ����w�5�)m����矮�a�d���A7���v����_����SΣڧ�)̧�ݠ�{)�B��$�M�{�{%?C��}�﫷%\���x��8I�=���rĿc^{	�c�^s5ny�r��	��P����l,�{���K7ۂ��tU�s��$�߆���LzQ��N�/aiY7����i����h@����Y�ٸ��uvN�W�"��"S�NڰWJ�pQO*풒:�w@j�3���.�S���L�+�YY���ݔk)T�y�Ue�SIV2�/�셿�2[/��~���P�!�:U�c:�����Zhs5/<��Ѓ#&/Y!�ȧ=�r��L����߳���xig�<�v��ɮu'P�k�6k����Vi������u�]��}�,��WkgT��֕z{tl�j:�����u�1.�<������(���Juj�������sǠ5�2������7�����W�k|�R���g�~�S�2�h��p�.u��>[S��e���-����(}Bj�fe�jt��,��!���>��Xy���r���Oo2�y�:D�y{��l;<��[Ι�\j�'v�'���ڶ�������ѵ���z��e�({2����+s}ر����S�b{^�H*�	������N��kÌZjT�b
�cf�=��w*\�{�-�k"�*Ս]и���+lB�3һ"kX�EZ�^瓂
�Z�ǜ�"�����<��(z�	\�P�Dm%l�N��[��>8�����ȳI#掻�����P�>���d����q�����3�%�����8=C�?j�U-X
����hݷm���2���[����z���{��KL���:A������v�:+�����$s�	u*��;����A],����x�R���=:�:/R�M!�����k+8bbG���ޥ������	�B���i)ɾ�q���w�fV�\%}ζ�G~}7�&��珹fl����"}3\�o�<����J���`�˽7�jg�:ئ���`�{zFs�� ��Y��G9f"����~��Ҏt9�|_��g�+�E<̮p���T���+��}AY�����*�¨��~�Xk۹S)���AB�(o||�s�Y�{�P�`�X�q�1{�O����*-{�J'8L k��T1��1Y�����5�J\K�°���v8\9T��IC�%�B��^RnX��a6�Na����b�0�%4Kl4�m[kL�Yv7qEo� �dd�.y�'u��/;���=ݕ2.�d��,ԡ<g���y웳��  �vշoܶoŷ�.�yM��ГX��޽�4�)��#��k.��9cS���y����|�J���g��7͌��鸕wӀ�Q�b����GE�2���J�E��1��q���9ӑRL>�-�1�/P�ov�w�Ӂo
�>�Y�*���\��<ٮച{ϵ�i�|�%�'K��L��7�Z!̫�,���ǠJ�����l}�1���C��II}����M�Cɋ��Ή��j�|�g�T_P�;��b��f]Z��c/2�:�E!�~�j���i��׾�������f|�u߷,�2���Yh����0{����Qn9�	8��{܎1�ry8����k^����ϱ����-�����v�x��5��{���-9�ۃF[M�v˲&�;����rnΌUR>�N�U�u-q��%-����z��M�잿mE(:gO׏٭����
�(�n�� (��
���>��G��Ǳ��SK�5p����1������s��,�|dUѝ��e���K���95�j��/A� :���٧��Owi�U|跆r�t������`{��m�O�^.�c�}s+���#�s�̃@g�����3�3�U��a�7��V�V~D�K�P����6�v�1���<��}���{#7:�=c8+���ܻ�1ܩ>�g(b�_e��]C�=��	�_#钕Z���#�ءƀ��y����3Q��rw'�&�Sa�{��H�2�ڷxz^��y����#Ș�����qC�	��uïke����P�?;d*��7��3=ɣ�n�*��7��������Ug�c)�Mm��H�J ��*�Bª����C(��S��m|�q��?��-��od��u�\^K�?9��ef�Y�w���k����ן��хv����n��/�>�_to�9�P����?i�'Myղ�W�۾��WOUxu��J��+���v�̚�Y��?E�{}r���|���Hf�ϮoLu:�j���T�Z#���ΰ1,)(q6���J�{���TGnm�r�y1��_�5�z�qQ��9���(r�����#��ǣ�2z�yVz����~�m�fAv��e����W2��� �-�H	N�.�֛�/�*�/m��a`�A�k�;0��Q�B�	\��¥�,������+����R���&��{���^ʁ�[C��:XyR�]rf��Y�Z��Z�N�h�����z�b��%ߺ��y#��3��|��������u�i6A�st�pҙYM5�ZE<�dz�4�lVԭR7��M����(z��}ô��U����Œ1��KP&��RQ��V��xv�O��{�<G��23�b�7�Dm3�Ip]p�IMd�ث�gIP�u%�&[2��wȬ��5;�aW��+rm937�-��=ӂ*�slN*=�H��s�֫�v"�l����ߤ	�=d��y�ߞ�-��1�J�*60fF���V�F�
�k������kUh厅,�����Y��k3wM��k����!���F+��V�G���R7/� ��cR��0a�)�*��zo8@�t�4J1'qW<�$��eK��4}Ǫs�R�4���f��.�J��:x�,�)6����n�9�<3��ֲw{{���X�������u���X���Jon��](	���A����a��:0j�>-py
�U�'.Ao
'��RWZ�`�[����mh.Ù��Y��%�2�o�N�f�
Jc�X��]mk��
�(fk8���ai�W9˂�[˛��D���jn-��_G�{6��*������W�\Y���֪;8��\o��9�G�p�6}Q��u�p>��^�V2$OL�x����_Tn=`�-b�W�Ֆ!n�v���K}s;6��d)T��Tcq���K�t��o���E$��٫:qg�a[p�����h���X�(ST�p.��oK��4�K���!��
\��ˣ0���7��d�AQ�@&���8P&d{�U�-�<wv��Q��:�}��Ӳ�u�.����^bu�R�N뗧��d}������w�u��oQD틫 �pnō����{��|k�W%���s)��r�|�>�U�B%�<��w����om�eAZ��N��ɼ���Y�f�ҧ�uݺz��ȟV��$}��=&�=��}l8��5깅���C��mk\�&����;<�2���{���ly����}�]���ʑ�s�ز=��ω�X7b*v^d/�SwR����Dȋ\B�}�<��1����|�Vq�fr5.e"|���$"h�F �S,��\��p�ٷ�46���R��~�N���n���dwZW�W���9^�\����(`��}Ѿ}s�e	/+o�nRҾcd'~3���'��K.vr��,46o���͐�g���bw�ɇ3�n<*s)똿^ѧې�/�(΃K{�~ mzS��8�4�a���gF.���^	Yg����LOvy���UFv�:�:���8}wDE�i^�J�d��U���;�b43�g��u�b���C��r��W흷�;���$�+�Y�7Rʱ�#_<}S��,]�)��X�78ը�-�#�ů��*��c;��x��v�#�y�묬��n��:�I��7�oԫ�7F2b{پ]�c\r�v�R\x��b�>�uLOt/��_.΁�0��z7w��yq����Ў�6�{��.q��}�{�����}��x��uSR-_��M��<�lI��������vƏz�F�P��7;7���j;="�>�NU���u�J���m�������V�8��޵�f�d��=�Spcw��>���r�|V�3�:�:ޭ��v��96���q�@85{��R'���}�d%!ղ�ϸ�GO�^?s�E��sqA]���;��;+�T%�J ��ک�;�X�����|����3����gq�����B��ϻ��[L�/���֓�1-;���j�w���_�	ۜ1�Ӌk:p�*�;��Ӽ��GK���<��Fy�ʜт�����ʺ����ǎP���W�uwz���o܎9�WD�ϧ<j���r�S'0�b��h�]��U�}9� �}E�}Ë�oc��b��d�3�6��4q����n��6jU&��-�V��u�547R@�k��I#f�N��)�Ƀt��"E�RIU2�R^�>��y��3c@ f� �?�P��X�b���H�d�H��ߜ�N˻�$�v��y��=]�=t��=Z{�d��(��B$v��iS��v�p{3A�˰��b�Qkw|C��/�~���λ���'~X�J��	��8�E���B����M�w�Yr��f����4����73ͱ�nN���aQ��|�6AY^�}*�*�x�X^�=��{���ؽ���Z�.B�+n����?s��A��;̝Ǔ��Gw�J���U&,�"t.YX�c�s{�����m��i���^��bʗEg�
�F�gf���P�77=yt{�l�($�f�:7���W���uǥ��=WrQ�j�_\��I{���_W�=ݓm��E$�4�2�ݖ��s�&���~��Bo��k=0ph�Ј}��z��6=��o����N]K��<r��I�Juo���ۑ߆�(�c�9���ϫ���(_8�q�;�� vg���)ߎ��f�L�2λ�
��e�v6[�z`\�B�M䆩��&9w:�7���=��tUٕw�uɛ٠���.��T��vw0�f�3/Gv�|O}��z�w���kF2��=����s���r^WN��b`o�r�1����9��A�ñZ�{"����!�ޯ��q��]^�Ɋ�����cn4*�}L��UɫC���QWI�� �gs���P;�5��ʋ�"��V��y����G7��1
�7o�D:!�H7����].��{4v�pQ�]�Z�TtfS�B^�7�k�ɜ6:������ʞ�_�/mˍt��ۻ$K�{��9�v����K&^l��0{��!yL���VC�CE{����bx��T��Sާ*^���=�)����7Ō�C�%%�H�����o���i�~W����5���W�ד;;Z���/c�����Λ�I�u+c�8���ݙՍz�q�Y�#�.��������fU�u��^϶��w�x��Ϲ]ff8:�嚜B&��0aZ����+
���\����:y�� 2j�����\A�ü�RQ�o1ok�Ct�])�V�\s-�6�<ɾj�'2,���t�8���N���ѡ�Ȃ����=i�~K۷K;C�􍙜4^�W�i���Y4
�v,
Ty��߂�vg����y����h("]��n{����'�f��O�H4!SD�e�F��݊�Z�X��ҽ�Pg?;����l6U�@F�}NZq��jR0�����g�g�Ş�E�=>5��h��)�٩k��~�=�g`d�Z��=�\���{c�N3�/޳Z3�rm�����)��`�}�&3��� K��V��^វ�QTt���<�3%Ơ]4��^���ͫ�n����ou��#,�/���P����	Q���/�I���n����{��t5�W|�rT�1�kD�T�b:��r��k.����Ž/�g.�Φ�sdҚ�/p�ҏwn���͢��q�b#���K�f ^�k�uV�ky��^��W�׷o�yN���Q>��ӭ�-byv�-~���	��=~�g�ďl,���|��^LHLAd�A7�H�MT����}�o�L���z�Svetz�?�~�9G�Ʌ_dɝ��o4"����yz��[�i{ʵi��H�Y݇�f���{��%�uv{�w�Pj������l��\+�ϥ�zL��c��ͦ2��������ŕ��N�j���W���U�Q����������Z��ʖ�~�ü7�0Fܩ{�L�VO#x۽��Õ��=q�y�9L��s������gzB�n��{/%C���R���l�����ct5��O8;�u�d�~�ct��W}@k�SE�����H����Ǽ(�c�yJ*��r�%���q\eRZ��Ǳl�*��X�-G�fv
�m U�0n�>��z�8(.�ӗE��j�MlWW	0��F��F$+�{�q [h�\2�u"(a���d[-=��d���ϸ�7�_#y>B�L]h��K6�>�����j˪  ����I/h��LI��N+����lo�������6I$�k�����m&-�:�����meΕ�y<��9.�O[���G� �zW3����"S�����!ϊ��8WD�`ݟ�<^�d�Y��c�#{�铬`��	3�B�y�1J�y;3��k�M^u̸����.m��e�kǾ�/�5J*�ex��T
���׈�_����ߜ/�ն��:1��o�7!��o���s�p��c�]N�ϣ��wy04Z��7�O���z��ep�������h���]���g�L�){¤c�Noq�=���<�3v
ޖ��S����p��)F�X�8�g�ϰV�������E���v{d�n�m�qo9��~����_�߯���T��{�rI��GF��+5غ��g���x��F�n���h�L����Ư{j>�:���*\q.��=���Ӟ�L,Y�;���N��ڻ�<%c��5��\��7�գ���H�Nl�����-��\z���f<�G^��|Vu%�s%n�p���x�K� bڹ���N�����n+c{#
=��zf� 秴.�;�����z���i���\�[�{O��weM��C�^�ߺ��C��?"�b��]2������U�1���"��I��h�IK� ��Ή� �h�p�E2��ou��7�{-��[��{e]GW�g��_�@�{f�~$vez{������6i��(�wVM�4׻
�d�{Y.��!�3}�>I�ӝǺƟ&+��DClOd�f�U2�:9�4^B()|���7�ލ#�a�[��2��Y����W�{�+��޼�:�t�f_b�����xy��e+�p�G�%��1\��k�D�խ��p���&t�	�ȓ����B����h�+�A��]���.;.d����u���	�M��
[{�TP�^!Guى�ߺ�Eڽn�}�2�ls]r��׳`Z'97�;�$����f����Q�5�����70�TPmQ
c�L�����K��+�8$�D�9;5�1�c�d>䇩\��e�&[*�xf�ў����.�~I��o�g���\ìA�۾J�ʜQ����x�^��Ⱥ��k���T��i������W�۪9����Ꞌw?5��<���0��g�s�(��!��`Y $p`�IH�K����Nh*yӯ~ڃnγ�h7jT�c����O�5��ݹX_&�7u�e�J�+�W����;��|�F�"ʨ��D�B�ܭ���iӚ�nj�h���R��w���5�2F�K��!e�o}eW!��&�{��E����f��SÖ�׫.����g�u>��gp)�鍵�6ь^e�Y��ϭ$���P������Y�_��lS良����g�Y/{r��rQ	[χK�cuL��cX��Y�w�u$��hE^<�mX��p�#:V�޲��?Y���/���ޡ��$����9m޾��� �:x<�a�
�s��_������Q���}��w�Yi������!ܨZY�Ѥ������{�=����ٶ̳%�.)e���,m��%$B`�U�/܂��TKa�8�uM:3���P��MnpdJ&%on�!ۍ�Ҭ#�z�,����Q��7bN9�kG����=�U���ӧ����v{ٮkʅ����ҙ���"�]�lo���J�ᒰp��h��U�۳��u��:�7&uȌ��b���6�m?T��}.W]���
�wj[�3Ϯ��g�E�Ʒ��ұ�OzDR�����p>���������:��=];��ܞ��1y~�!��jS1o�<3�jĹ��fz�0��j� ��(M]�����2ٽ�2��
��ߵ�U9���upEݎ�i���g���o3���{q�r�D"J�R�Y3�걒���Vp��*�΄�NL�*�Ù(��W^]۾'��tx�\J�r�����F�.G@E�O+ܣ*�+�&Mͼ�Q8u�uؕ��ܣ�1�6zTM1r#X�QW]X�ɫ#�:��f�$v�u�X�K��h=g:k�Q3z�Cv[���iN�=�c�����2��'�,h�:�XxXX�����}���=����F�+f�'!����x�VWDcq�;�&d��A{Sl5�P������;��n���u�N"��p%o\}7����:`�,i�v�'��7�?����3b�i	z��c�����pu�٘�=��8�iu����i��U�#@uq`��t#Ɉ<�Q݋�,Zkvʛ�咪Q��\*q���U�1�;�S�h��sW'x���y�C��J����&ӳ�s4�'��<r��g`�:���n�&����Qc3�c��d�����/��ԇ(���>�%��2K�&�'0k��z�l����1���f��3v������fUǷuU���7Ye[~�w�2@��S�1���]J\L��͝�V�p�����{'f�і_ܦ~;ɺ"��ǡ�e����;Qv�[�g�[U�F�%�˔��"u�Fޡ�:#�r���2i͕�c'mI٤W	��?���}�Ӭ}�i����-��c���]�
˵����Ǳ��z5 t��ir�ZV�AD?gc{�Lr�[d�d>O={�=����O=������dP� KR��m�մI-�t  $�� �� 	%���ثv��a&�BiW.U�2F�m�[hVji���vl��I
���Y2h���Kj�Ɍ�576�  dKe�$���0ZE�L V�B��bQ��ܶЭ �-�W%�}�s���c�6Ļ/w�L��O���,�'�\�̏	{��@������v/M\M�r��w��p5���6>�Y��rI��&�o��w�$�6�b�ۺ��6ݫ��m��7_���-+w@�m��D�d��ۋ����w%�M&[G���s�<��0�m��p�.m�P�`ޓ��ŵ���V@��P�k}}�T����vm��،�u��[���   ��        EIj�Ԋ ���ܒZ ���o�����w<���m�I�8��SZg�u�[�ӌr
�����Z����;-��6z��t3&h��H0aT���I?ʺ��r%�a~�p?��^l/�Y6�*��ed�f���i�n�윯�]�,6�۲������e�HKc�݌(hFIBݵwc��燽��\������v��]�Zմ{r�̀Wf���ޅ��R%5 � �.���ɛ����d�am�y��7�����^����v�.�6K$���Ho���s�[<��  [l��ܜ�M����f��s���}��g�~ �M�\����M�N^K�;n���w?G{�^��O��\�qh�6�� n*�9�r�{�κ�u�S!�6Ԍ�ц*�oV�''�B��������G�^��ߺ�x`��b�&7��t�u�G$��r6���?����[4�0��X�ܻ�&�ǽ��Mtĥ��4o���܁��Ԙ�1H0����a
����׸��δ|V�#sq��!XTj�c~�]=���H|r��I�m����^�?�c��e�GLqƆ�Dj���w���W캒*{�oˆ�����̯.4'�7J�R,�^ׂ�FHޤ�+��z$ERA`ə���ݹ�޴s��x�����S}��ư��h��"�]yG^_M�R��!��g&E����=��|��N3����{L߿eγ).ОDun��,�~�=z9:�-�>G��=����:<�P��C;�2E����Q������2��@Q�cg�tOW�p��͵&u`B
	�z�\ �#d������9Y�b�������0;ek�-ݑ��w:,M�ӹ��g�.p�x���:��>���S��U�S�tN?YC��z�Yуi�K٘�����Z"��u\����Dŋ����]��V�� W,Dy�����{���9u��f�<ǗA�۽���ϥw�tϺ��A�Ǚ�=>����������k��L����p�ג�V�(��4�(xN�g{�q2����w�Վ�2 -HT�sW�3��Jȸ��������r�?�.�;��83�z<}��n]f����4�ߞNѠ)�(�g��q���{���]P��T�]��(� 0
�&� ���Mvy0.�$�4�k���L�o��cG����xY�'�Hg?R����yV���7�Q��ދY��+4E�X9��ީq�|�r$mg������=�)莍���W�N��"���ZM -y{�2���75Tqk|�u��e>1�6}��9�>�G#^�x�E�gD����&��������
�~�ٕ�Ǘ�ғ�nxaKdN��23wLӉ�����+4x�j�i�M #����RJ����+*d���$�!|�/[��u�Y�aV��ۺJ�޳%��s�n��3T䲖�}'}^ܽdI�c������֑V��}Z`�y�wlux��lSԷ�|4g|�rh}[֗�^�=+@*�h��(�s���WV뚧�b�l~��Ѻ�ʉ�oTz<*ο)�b�~�E�G=뾠����X�̻���R<���n��.���{�w�{͑�����n4�<�΁�wǢ�^HǊ*�`A<�rq1����Y��Y���^<
�������=��V��!�k�&�l�H�k��|�� D����*	��>��5���Ĺ��<�=Q��6E�����$/RT��n/����F��5��>ܯ:�^
���3��y���x|h?\Y�>�L�z�L6��u�k�=p�G�wM�<GoO�ǅ˧5�k�'|����WU}=*@�k��Vk����F��anʟJ����J:cv�$h��kR����BץȳIL����� w���~�yЦcGm^ü���^�l�z�9�m���U��,u'gG���^)&Jf�m��x���s�+\��Ǉ;�rL���k��YI�4�eoM�|�'�S���=�>���*k� �?_����у?s�Āi_��ʢk�at�(��q1����^sݷ��q�����P����ޮ��G����4�2 Ϗ������~����9w�v�����4�9�b�|lҡF��C�[��v��p(i��6���+����Q�7n��1��_d3�MS���~؛<�: d�� ��7G�J�@s��cB�>�OFO���F��2���q����b)�*Ԡt�����y�2�9w�*�h޲�\Ou��z�M�Z_��$s>��'i�W.F�۴g֠�5<\i��=s@�z�뱎���&���1ZHc�g��ܐ�3����!�L��g��?��	y-Z���b<���f�'|N���xh�>�Ol��^Q��.�[�K�5�\r�^�����"���W�P	#yM���Dxgu�����'��������v|G���O����ޥ�UC^Ll�Q#����n���*���{~�7/%HZ�E+ږ�����YhZ��V>�*��~�����y1��暡����l��\�����1�7�,�}�n^��l�n�m�e�%�RI�2�� e]�`���n�kyߺ����Ln��vo�nB�K���&�7���e�|��,ٖ�@ kIb̾U ����V����Q�X�����}7r�ݶ߬�/.���n쟟���9��@�����A_y���*�{��L��j�iܗ�.,�vQtbw��G�[6�&��G;��k*bǌ蕡�M��.nz.����s=��~9$xݚ��#I��3�M��Z���ݖʩ�;�X��=�/�9�3uM��д�QW僥WLW�[�Y�Fa�1�}���wJ�������}��0�Y_K[]�:L_�Ԩ`�j2/j*�.G#����䈭9��N}q����QOS�U�"�h�����(�ࣵu�D��7c�)��H�cw�}�i1�o�ud,*���r5�	�s�xgyvƾߵ�I�|c�ܥ]����>��V&qd� Q��P�B�S�N���Q�^�p�����OB�SA�I!Z*%u	�m�99wl#e���M�:�{�L�
��LZ�3Qjk���DmjYs��,|(m[��N5�B�~�,��G@���#r+���r���J6�D��M�eaĮ�=Z���ᮼ*�Ne�T�o6M<Y���z�[��&@�us��H��]� M��R�#w{-�7����E�JsD��(��pwot�)NM�@��2��3!�ͨ�&l���o�s��9�|x��UĈ��{z&�(��~쯰q�6�c���xu;�v_�F������Ue�/��MD���1h;��6��Wޛ�-�u����e���V��q��������^�u��룑z�)�9��p�q���,CjvԽm�r�����ami]������Gw��6�.}��pv�������
G07���W��ou__5W� s�x������~����띿mR}Sk�3���@{��c�k���rc�O�k� z�UO��?dX��.���ۻ.Րع�Z�ų�{�q�IL�爁��;'ë��7���Lg���'�1fIiz�=���?Uv��jx�w&^٘��Q���B18(w�H׺�l��n�OI�dV^Ϗ��`R>o�c�G2�k�=���Ns��W�Q>T5�쾁[�;�c'��5ElVxF�j3�m���ǊfGQ�s
��K������%u�^�m�=��d����s��z�L!=�<�Zؚ���#���[����L'Y�I'Q�ٺJ`���Gu��և������O�5�Y\${o�R�xrT��fp�2,쫜e�'��7����C�*~ƣF!Nr��;,\��2w�3����9�<��ԃ������wz3�<W_ht���N���)�q~�ܨ����c�.חC&T	w��`�ǟ[�����u��7 ��� /Q�������jo(�m�v�����z�`�S�B��{Ѭ���-Ɏ�Os�H�"�$�I#6���_������s��f�~���M�^�}�(�^�bU�9~�
1�M��wx_
��z7�t-�k�}�b;e`�.���Q=�4H�y#�+��>d���9�1w�T��~{E�;��q'��/��0�O���J�1÷k'���r�s.��:7��_� pD�J+������p?ݬ���x��v�qk�e)j偭�ˍ��� �QvbSz"}�,9d�U	���>n���;���d�Y��{ʓ��82�uc�b�93�@���6�:1���7
����u�A(R�Zw���p�f�aW��/]k���5��[ى��qC�ms�4f��*ґ��|el|�����\P�C��;F�[��c/�ٓ��(7m)nj���-g(�R�V�O�<���I��*+ϫ�.<y4EqZ��ߥsj�xu�h���X�9���p������~g����3���o�d���ϟ����3i�m����?ۆFF�On��Dy�9�Ǖ^su��0��<ezzV 
{�=�\R
[�=���5��׫}�1�w�f.���:Ю=܇�啛�Mg
�2�Y��A|�NB�≃��I�0����
��唔v�L�����W:��g����e%Pc�K�}�&h!çWxώ��Kl��7}~ɗNc;}G�O��x��:���V�ʥ�=��Pǳ<�|Z�R�� K�z�Nyd��\�c�.���x�9͇�f&w6[J�����l�/3f+A�#�T^\�{[#c�� Z������0*/'.�h��*a��W�\�o��N�y*b٠�Tvb�g��6T�>�@}�r����O�Yq���9�p��fn$3��޻l�=GK���2/Fn�t��.;�m�c�� w���������厇ݶ���@���V�Ӝ�a��0-� 1d�We���f�R
�6�D,��v1��:�̑we�Y��f�s��^��3n��[h $��gy�y�����ɿvI�}�������)t��DC*QA�f�� ��-#k&P���@ޏ*��ǔfkL�ѕ*�
�{(t�Y:�b�d����F�zՃ޽�u���,�|4e��t�}���0v�(lE�����\�o�kp^Y�F����kJZ��}ʀ�+W6
�e ;w�}>+�'��4��>�)��Rģ� L9��gb`n�F3%En=������/��&E�7
j׉�yMDɍ�����N��Pa�s�y����O2�FPw�~6O�$��/	��{�:X�}��M�0FmIaҡ�2�7ׁ��髫W�$�1m�*\�зw�Ԛ#�O�Y��Ԇ�,�	FEB{�@b�7�T�{����xg�����E��Q�ʌ��="��������lW���m�[-͒ۯ�99�[�����#j<��v����c�/j�����u���Z���;o��b��s7t'ŪT6pCS,q;�$j帶h�������Ҫ�s5��g�ގυO�fx��q]zN�u`#+:B��Q�~η[������n�b�Wp���2�=f��+yR°�<9��M��9DI�Eчk��9;v�9�/Ve�2�,��5\^9*�7;�~�L|ex�B�^@k,z�IdS1�F��39��U�w��Z<��v3������#���5v���fL�-�T����==�\_>���>�c;�X��r5�'���Kw��őس���s�E�`_@��pC�:!R���)�`>�{�)f9{�R!��_��]Ӕ]jC��y���i
힣E/�Y��{��i����w]�5�tg*܍��X�ލ@���Hю��M�yɏX1��p*�1�Ck�v����ҍ�+)S�y!�l(��S���@�7w~�C���y�w��y��d�i���o/W�#,�8,; B���j�� ēY��m��� #�z����y�9����ֽPi�D����!к}�D.ػ�ɿwT�����pz#t��.�w=}�3�� ��#mѦ'ъ�[&�?$�bQ9t��=��yFQ˷!���6���S������<NV+t`N<�$	����?b��)8����rh>-bo�E���b�:X�O	ݺ�px7��ぼ�k�7�:�]�V����d���]<��_앋v�r�u�Ս2sd���WF���$��0-u��G�D�V��u�`��l�2��'nuc�
ð��:)�p�9ܴ�Rv��w6D�CS��j�Dsl��k1�|��9g%������6���� �Z$���蜽��F���:�S��Aw+;	��ȥ�r�i���ٛ���Vs��"��W:+��+P�OXo���^FKe2�n޺G*�^�P���dK��t���'U�;]���H*��yp�@���V�Ə��]K�����諱�j�����,G}��Q��iA�� NX��K�3��ډ��-�;'U�a6�����Vy7Ehf�t�_;�,pT��Fл#�*\�p��A�ݶF~<�b]��9{
fVhŠ�g?L.�\��t*i��J�ӯ�*����{R�۾�'�ojB�LY؆��p����*���\����JW܂�ݮ!1l���w�P���r�,Ǩ���jie��"*M��bܵ*�&���Tf�a�5�@�qh^h�%�ǭ�,}rأw�p�CR4ŚL��܂�%+C�"e���j��!Ձ,��W����c`�o�fF��ry�js�΁`oLe� b�?VرaY8�p8kB��f���s+���pI+`�J���O���)/X���\I�:>%sh�u�;�JlLi����/��,�՘��]�&P#"�N�oU�حEP���wgY<v���]u�t�W�y�%����T���Ei�]&�fa��V���B����؆��ۊÇI�i#�.PVåcd��TEY�蚫Ν)G��N��J�md�.�i&ō��TM�@RB��UiV�UnDl�%Z���hk4�%u:ra	up;p/5{�R���)f�H�Wo&��Ua`�h͜7y]U�[���nh���Sۢ�ѽ�7�"f&0j=R�:�k�����1�;	/Gb�(�p�F�����:�3W�9�9��l�dK�M��6�uO��{��7"�����o��ؘ�������]�܄�wb��J�˹��,��@�>��ݽ��{ޡD�3��G�W\>ޙ!:j�[�'���![�>����]��z�s1l�7�l�'i�^�㸕2$���F�OtTh��Ν����i��*=������V���n�|5�R�#�D��tzmT�Cj(�r�����vǷ8��p�ޅ�9���L�gx�Z�ϔOXT&Li�7>����7�RE2CH��UP)"މ�2��@o�'W�y�F;���i,G���pU8B�cɈ|�G�Ϻ� �f�F�>��h�*O�|�uBZ(��)R|-0X���/��Ϳs%(�n6zT�}�jr*�x��C	q��̕����Mp��/�f�du��F?b%[@g/���HNb�/�w���}^y9 �����UOI��oq�>��op�k�$ә�96{u�|Rqgg�e���	��k<�|��.�Zԋ����0|O��Q��Nk��2�^��Fg|~�;z�f���~�rP�c����aa�s�*u-�'&&���<�[�uX��X�(~�i��B3��Uhy�%ۤ�䓢��^-���Y��&*��$�b�f�~��5��}ԻH6�FQ���vZ���Z6d�> lK]ȓcG�c�������7��
�2N��E��%_��2�T{+9,�/�ݍ\߷��rn���_{3����<�'/��p;.ΓEK���r8�}{-U��8}ł6���/#Lg%�(�}r�m��-�S�h�]j慂�՛�:�ޫ���2����0��S�K���Э��_w��a�]w�=]Gu�K@�t�p����6�y��)����GI���h�'��U�Ӿ�獊���)j����< @y$r'2v��9�u ����W�TƠ5�U�62���эh�鞫]yN�����F��B���g|��͘�"#靧�8��\oL���g���SW�fh��'VT���R�x��*v�^�*tG����m�^��~-n:DZ�'F����[\1H�Q̊����f�]�%oSc{�V��v�sm� �%�)��Uܒ���8���wK}��^��&p�Pν���������7�C�iu.j���e���f\m�U?��bn�őF=�{����>��n��ِ��5�M�I��{���l�ʒP �I%��rW�k�Ǵ뾆���YHJ���jA��M<��7,�m��g��f)Ac^�H>�=š�x`�p�0]g�d��~w%�=�D��'~�-c����TC�|=ǛL��}�hF��������sG��֊ӷc�}���#���>>�['�u�S�8�k_W����BϬ��|���׽�ǝ��c���<1&M�<O_����ߏA�v'�;�� Eƺ�[Q�{��3�Og�|&��K�(C�>V8N�,8;�\��;�@��묍T�wm�񭯅*���ُ��v��
[g�B6��_�0B��=[}�j�@�&��1�W9p���gս�?�yՕ�	9d�""d�!Sm@�o�����ţ_i�.6u�T�������^�MN�fW���N��|��{P)�D�ި�$b�3K}�s�g�s9�3fĻn�[6������;���ʕ㪄&Z�U+ �=�L���U38{�w-)�A����z|ks�3.*N�c�,�~ִeu	�V����X�u�<`y�ya�����g>X���VJ�T��N�G�k]Xzo�v�(q"�����̡��l#���[#�W�����C=�nj�*�X��o�c��F�&^��%�jB,�etg���ԌG]���(������E�C|��=�ǷTOj�Kwul���pm@ْ/y��[�S���|k@���i�LN��}����o3�z�_e,3�Ȃ��1�G�b�@��Py�g�!���)�R�6`�(��t6s�
�6/�}^��0��:u�j���oU��qy��T%>���&YCP;0���e�,����$N;�5��_�n*����������n�YǑ�R#��"���s��j*�e�I�Ʋ�3�|��x�w�l�f& lQ�:N��܎�K�'�V݇�����ڡrn��Sr+��;�ջ`�dV���~�J�ģQ3������ ���4L\޸�/����;^�������?M��$܃��ؐ��+R�Үo<za�f����>iC�.1]�z��JLc�K��[I�CD<�3\��k�x�=�}��3�����z��lx<�'�/�=M��>\�9��ۿ�p������cR�j��~��g1�z�
������h0W�{��'R0XX�,�+���5fe��u���͓E�Tr�W�X��n	BP�6U� �h�^r�Iö��f�ñtzT�K�1�=�N��}�Ů]��",�Us��'+�,�|sǮ:b���� >਩���{������ݯ8�����j�}W���l\��!1�@w�<�q�N�޼T%(
�DXc0k)r��+H�*�WUG�8O�@Lת���A~�v)�s~�ۂ+�!��x6w\��x���?+�S�튬Ӌ>3`<V�8��Si&�l�CO�9�9��IϾc9���'�����﹞�a�C���B #Q��>����m���=�B�c�v=ۥ�X ^��p��ې���:}j,�uaҮ޺�4S��o�o��Nݱ��/jU��c^����P�6&Vv��
 Y��59m����vՇ���W~�e�D��lM��]x�:S�*/[LFF'W�ܛ\�,�-W�F���iz:nյ����G"��p���~yhq���]*Pc���@� b�qX=�q������M���V�� �����D`���c��+����}Ǔ��uM:�d��˛;j=���;��)Z7;a�]���]���υ#N3���'.o":l�4��w��ü�օ���/��M'�4u�\��Y9��N�a2��e�	W��l�����7r�Q���jh�ň8F���ǁ�K:H����7����ޑԈ��\��eȢ�xЌ�T�#һ��=���Ω5�M����g�+K�&$�Dnڷ?�u�8�b��d]��ޘ�7��iw�W�}��;oV�۳5;�u�z�g��ͻ\gw}r!&į7�)��r"�����p
ӛ[�3NgN�u|O��힇k��HTiE�c�%m�2��nQ;�AwOO�_i�w�!#:,�� tϪc�������|w{�o�(n�;�}�#�����b���g4��4�����sH��i�� x����
��g��;�{LO�եmI����*ɑ2t=���}n8D���<�^[~,�Q�� J6�`9���we�nyi�B�ʘa�WpԤ	՟"C6�W�g8�θ��{lp�Fe��3�=1ޥ�m������{Z�
�鹊N�F�-�料1�x�r���v��L6�F_�ݭ컔�ņ� �7���&`f ����HR�v$�W���W{&a�|g_vo����1�ϟOe��m�[I �!,��V]dݚPe[V� c�5-��M��o���{�;m�"j�l��-٤.}��3�s�MI.��� -�E��{�2w��wP)V�Z;��n	� �I<�p�v?8A�����0�@��D\�� ��08��r��;�;g���h}Vm�Q���[3
�X:+o/q��f�W`���<O6���L�����u;�s�S+��+L�F�а`?P�\X�L�sC������?��Y�����Q=�~Y�Y�cC�QYѩjXc�n@=�o�������ڦ�1�[├��i�T�i�S�FP7�j��
��O��1YY�١�H>�y��]줢�.ZΎ�{p�b�����H��i�����vf��ΩRD��Y�l���7���#��*c�W�����V�.�� ���́�ڑ/Y�a���l��=�*wfv������I����P��{��jY�Eϯ��m������s1oV�=�p	\Kp���ɔLT�!)#�ܴ��D�EvX9�|[,Y����i�&x>�䮹�1��Qv�Q���<C�EnegF�U	�
 ଵ���I���q�(s���`�u���\��5��	�m<T�(gv�-����)�-���^�C1�D�`v8NYd��ٝ���͒N�M��̦��%�*I�=�k���'��0	�md��.��׼�cݓ��Gz|���}	���c��n&% 3���^�%�[�|��)i����j��̾�	����R8J�G��m�S���5�Ҕî� ��o՝P�>�^��n���.C2�v�Ǻ�oTb�z�<Un���(M����S۟}��q�S>��7�b��Yc�]��=פ�l����n���u��'�Y��c[9/V龟sſR�!#XXEA��+�2����և��H�=\T���d�=���2/@�����ߗ�)|�d�>�\����xc3[��}IP�����JO��u�m���>�ww�1<{���_�'��t9f�O<=
��ieHPp�+��C<=�y�^d��ݘ뢷qߵ!���D��ܙ�*����P��o��r�`��k$��%Ɍ�N]O�{�ҡ#�ϴ鴮(�O4I>�h�2��v�9�U_o�H�nl���](���R�����&�����d����^.b��U�W�����-���2�4�9,��:�?F�����.c�M����U��e)����чռ�|��ҟui�Ge���Ex��5c�&���ZA�W�k�����#���GU�	�(Y�^����A�
;3@������힚�w�s#�w�7�f�dǰ�����$M������ą�P�����ď6��]���ح3IF��U���lj}R��{�����
�E�����4,���ٰs��D���Az��(�;��Z��{�Ƒ9����EU
�?�/kl��Ͷx�q� /?}|��'���W�����������{��=��q}a;c��~xaN�l��=�}{'�y�~��P�y`�ٞ�*���c��y��S�Y�"�MGb]���}���duǏ�=��ћ!B���S�͟ 
�6�~�.r5m����sj@�J1��Á�٭������J6���#f�P�����X����R)�:�,�?�}��tZ?��ml�kz((��Z�i��]���kyV�U��G�v�˵��*+^����u��^���};٬1�C���Y0�śGQ�Ɇ�$5�0��(ͪw0x��3m�s��l���(ĸ�Ci�n�%G+Yu�-{;����l��"������?�p9Gt]˷#+�Ys���[�-ujz�vE/o�<�7���j�|<,�v���$���O�#�Ti�f���^��b��xv�{;�U�q��^�Z��iբv����<��o��?�+5�n���s��W4�=r~��G���������5^�����"<`�ڿD��L{��]��W�dP�G�ӁQ�������~Ϋ��yEr�S��ӨO����q�>��ҀB�	~����+�8k^ɮ�����:*f��#p�=�V���z�)&��Z����S0fOdeH��+ZG����f36��X�DYc��>&>pV��m~y;k<��	*V��uH�j��"3۳�uY��lO�cZ�㽧��.�v��z��gS]�_]x��,Iv�P���S/�v~�w��f����ď���M�D�ByJ��3�*�Mη�T:8
A:���{�y�Y�2�\���Ԝ��w�����\ٓ>�|��u>��{�;��>ˋ.��tק�-D���䌣Q�Ҥ#k8�C��d"�.�[9ro8K��u����^�������I�����ot�tp`ѼZZ�&���
*}Y��\�N���n��ŶN����ĤS�i�zME��?�m0��ݡ��R=��}���g<MԔ���Y�Ң���A�����Zv�k\+���o�����,�k�W������̓_��y�?o'���Q�M�o��w�d{�c��@��"�]��'d�+SeØ�-Ef�#i�;|t"T//��Q�u2
i'�KwL�5����{������$��$	I?��Ԅ$$��_�HI �@h`@!?ń ��	$����I ��@���IB�� 	������$�����$	$���@�O��}����H�{��b�������~�������/� Wuk�?��/d���BΚdW�*ݵ�0巧Y��ƃAͭ��V��j�aq0��SַQt���偵�V!w��4��&�n��S�NGz�\Y+C,Gv-�`��Rn�܋Q�R��t!��7ƞ�/6�{�T�י�V�{EJR�6�Ʉkпi��4�헷��+In6,�kICw) �%�E�b�9wWkU!R^��dݢf�#	8�zЙ�w%�9�1�t�ȂP܁I�[	*]�E՛�̑��`��1��n	�qSP�R�5�/l�j�d�wGc[�h�b��q-b]�Z��m��i��m���Ml���I�i(�L-4B���n�Um�����7Z�Mb�dl��s%��]#z�D��iܧF�6Jp����!0-Ւ�cy�Ϟ��c���^؎\�6S�sT��/J{�$�jM�4���3+�։������ۡ+(#ra��s4f�֦��ii�1k4$t�P:��'6�H���F��WmR��@��Ci�������Q)YVw+B���DH�r2R2�b��
ig@͂D4�ܭ[,��H�;j�*�f�r�̗w~ES���K�z�N��1�L�mj�TUl��$ܩ6���͖ �)O^�T���E*@�#�2�����k.�	kSV��Q]"&n%e��pb��$�OHӍ��nĵ7��a#T�'4j��f��Y.j��k�*��t��y�v`�4^M���[6箜��G�EȆ+RI�F,�U��͏,�%�4Z�Ь� %X�ܻ�d�ʸ
�O	j�\zVL�Y���.Pf�!o��׷��X�uQǰ-x��k�ke��y!l		�MZ"���$�k��ϵ^m��@�&�â���U��u���WPL��id���Di�dسJ�S��d-��!�P2Q,n-y��hR�oU��J��5��FXkԪ�v(5���h�$�]:Z,�����6��r�tr�G�j� ǽsdW!�+��+z�h�a[w�XA�K_΂�n�N@mi:�+f5�y��!:�0*�������B�eV
ݻX-���m�EF����Mf���%dɶ�4���R1V�t������� k{gNLr�J�h�R�C>شɷ�K`4c�kt�a��.��í(-'�,�b/J6��6n����d&�hZF�3�jL۠i�F#^Jf,��cn�0��f�@ǥP1k�j�YG.�����A���d�U��K(�n�l.`9�@)�N1OE,�snں�I5�v)�ݽ�rVf�Z�ۨ��0EkVcm\��9x1��\�Ah^�ĢN��!T�̩���"W���Dja��@�y0�wX)ڕ��"5� �Oe��
�No�2O��**"9�-�ɀċlځ��3pn�;ec@�ԑx��.��h\ϙ�pD���R�K˹�at-�����W9�Q��q=⺞�����9�˩Q�(m�Yt�.��;M�Va������:O&l-Ve�r��Tr�c��ƫP�)�q��o۳j"-&!ǻ�*�3
��f�X�&��qլ���M�t��M&��H�����3/�k�Xf�1�Ap6��
8(4�M4 ;购���Ҧb������ťMp��[4CwxJ�M���;��Z����m��)h�P�j�;�4l	m�we�E�pV�[���Ӫ�i��5���M���V"WwYt�؎%B�(/jβ���Ɗ�b�A�E8��l�40���wk]�#�ԨeZR�Kd�D�
ژ�h2�1���'&��7F"��Pi�aڔ��D���+�w�E=�)�eEc�OEW�q�#n�p�͢ɷz�JԜ�iJx��"{z0���gawlf��(���#k"ƅ�/(��fM��׳FC���&K��<ɢ�l���0E[$\�Fr�^5�k,dAӬMUC����VRi��4PY$�ٕ��O"��r�`��-���6�Rb���Z]t�R2`6V�pPt�]!�;�����0�ۿ�U;�I�L6Ec�SFR� ���Zė��Rf�kf�ܥxԵ��uMO��73[�)��ǅ�&Y�5PFڍ�RtuA�oN�	��Lz�hCR�!R�F�	v��gյ%"ӹ�bVo��p'���ޫ۬BŒ��R�Lfb�5�D�"�Mպ��#R��S8tV0��+��gF�QL?	z`�8��8������I,�9�\ݦ͒�^9,�K,�_��%����O�+rPb�[�u��f��p���R����6E8W觲
��ș�Ɠ�xYr���\����e��.0�՚ i�J*wdjH;�����3L�Cj�1�KV�n�+�bT�B-�f�����=��X�$����6��V����Ȟ�̖��0�`&�\�e�蘳.�%@�F^i"SmbU6dw���֑F�Š�U�/Lk`����ь�v���QSH����쑠��&���jFkMm��BDo�E�<�h��l�0cqg�1� ���A[l�ތ�y���o7�f�����i$$���	 �2BHH�@� H��IH H�I$�$��I	 BH���� $ `HH�$������� I'�v�����H��?x���� HI�M���$�� HI�_Ւ�$��ưHI�������sf�I@�O�� HI�'����$� I'�I@�O���xg���sG���� HI�O������@�$���@�$�������e5�l*|�j�� ?�s�m����%�           -\�x                 .;�H$(	@              (		
�$                  <@      hh	��Jۍ����S�j���ʦ��� w[p��F�n]S���[�E���6YK��d�p )��nn��jܵ]��Q0 @ >�� ���  >���6݇A�ݾ��K����rݽyG�����=5�y��v�^��;�Qj�í�w��)O��|  �      }�t�7��R���:S�i]��� `���^��^^�J8��-m�7u[f\ :��\��5����7Ϡ }H��u
�ںSg w��wf*��z�4��p^{����za�N'6닮i�w�yݶ����{��<   =    �c���������^f�s�׋���W�oo;���,sE��V��v�wy�ʽ��;�"p {����ܭ��=�mm9�^^ۓf���z� ���=�]�wm�ֽ��Uy�{ok�����n��(
�e/w��g���f���l��/oKg���:;��  ��    �5����ݽ�݇�����y���;�-x= ��U�s����n�w�^�e�x��mt�����ݶ��=�^�ӻ���^���^������s��k�^ �y�-<m�^�-������n�w�nU������w��:Z����ͯ/e��zw�n�  
D    PyQ���ҽ*�^�om���@s:拀gV�m�V������nv.ʜ{���O w����gv�P��W�{�ͮڲ�;]�K84u�lW;;�pm����mnwu �w-�� �S���j�h9�����j#��)k�  S�hL�R�1 ��L 	��*�L�*�� h    U?��f�T� 2     *{mUJ��	� M  T�4�jT�FM4`� �i��14i!�i���=#O��(�<��������~�_�G���yߘ^��l������@! �k�`�a�$�$�%��@?$
����w!�� �k��@;{d*I! �~_��I�P��Y�$	�Bc	'I
�BHT�M!Y$�$��bJ�M0�a$�V�Xc+$��I�	q 1�c12�CMI �d�J� T�i� C�
B�����!�`V�H�B�Ą�i�B��J�!�
�1
�P1*+ �!�*B�`V�VT%aX��@�Y%HV(B���R�I�&2HHbJ�I�	X�cI �Y`I��$!���	$�*I�V@�d�%IY�TI��$���d�1�$$���$�I
�,�
ɉ �
�����$%j@��$��a	+RJ�%�BVVcA`T�(LJ�BT$�a1��a
�&�������IH@4�2I&2I bĄ��` �!�������	*V@%J��!,���g�xmI��@��+;IFE��U5Hk
��OځRj����H)���~Ԇ�TYSYT2��B�V�V�U��!P����jW����L�6�T�I�N�+�wJ�-��`��̵�����k`)
�aRX�P*V�Y*WL1;CH�B�6��Aq`f���t�j�D6��;@�!�V)Y*T��ˆH�J�������f%ER�l��*)Re����@�Vc���\�ĕ�*�z֨�t�l1���3(U{aPĕ� ���XTZ�Y*TmJʺ�*
\��T����T�b�¡�
8�RVi�r�aZ2m�&$��A
�S�2!;a*�4�0�++(°�4����kE6��ш��
ZPY�Q�2��+.X���M3!�]�eIP�;IE��*ID�%��c�0��b!XV����\|r
�m�+ۆSv�v`hLHq ��$[]�V':HU�V�4��W|���6��ֲ�f��%gn:H��ߙ�8E�m���6邋E��D`�
�5c�V
F<Hib�E�Fh��2T�]v�9
�Յ�RQ5h(T�)�c0f�PQ�(��#w�y��q!Q�c6���4���Dći�����y�@�N%i���,�W�rY\HVE2�(ZfT�aFr؈,Rxԋ��1X�4�2�����-`�Z��8�:Hv�_5̼4��;f����e(�3����-��9���U���q��\h�b(���C�;Eěe�f'i:eH) ��N�PO)�b�i!�b
j�:݆(ԇ�P"��Ғ�U��4�p�`3�f�Hq���P6�^wL'L8����RbB���r�f8��leb�Hq�T	H�P��`�l@Gt*����(���x�d��T�6�2�S-�H�i!����P"1(%B��)"��E+"��l�Q,H��@Pc$SL!�,3UhŐ镂�� ��ŌU`,q Q	����p�H�H�V(v�Q�� �0��c	PQb�b�,�+UT2ʪEP`V�$�FV��VB�A	P -���b &R��E�$��E�aXt����E�����1
�Y�UX�N���@M��$���� ,"��T (((A`���`,�d���T�H,�A`((H� |���X����ڛ�"tf
=��O�h��i�r�gԞ�S��uZs}5啙y�H�WJ��R��ѡ/ֳ.��]���ﱕ�ߒ>���8���^�{�HB�ܿ G]�>W]�>}�yٕ���w�op���P����rx.���UC�&��k�*ږ��~��&���܂��/�v�U����(pV{���?�t|��y��9�k�
[j�[~Ԗ���Foι�.a��7<j�Hi��wB�U!�AE�V�<UJ�i�S,*ʊ�Y�v�ą�6��Z�$6��6���Ì*���Hv������Ѝj-�R��{�6�� �6�8���N�$�9�)�^q��f��vk��
Wq!��C�$4�R!��@��m�i1�a�!���HT����p��J�)*�d�zsT�!��ln��v�0yeQ ��%jm��Ҳ�ˤ*(8���W�`�wJ��8f�B$;f��P�*
<�KCb&�#��9�*��[m�J��2���
�C�l\��Ŋq)��L�\�S�2��.$�X1a��I�t��v�a�P8ʓl�(5%eDM��C�(��T�B�E�m��x��WiTCI�I+6�R^����w�gS�2�����X,��tкκ�q˛��O\�6�
C���M#�b(Xl�[U�q����F,P�ZPF���6TL���Vb��29�U�QyLąE���@oY�c)�ut�
�f@EA4�:α�.q;w��z;���$:E0C�h,��E{j�{���[PݲC��Y*��v�T*J�0��HbbG)SN��FۧLÛ�Օ:Iq�
������w���J�R`b(���oGU��s���:��{z�0ί[ֶ��C��l!���C��!��$:`f�L�}f�nq��I�@R!�AH):dćH)���Ă��@�zIޱ�:HT�;@�C���Hq���C�$1!�C�
��ig2�5�w���%@�B�;�#�HqN"�R�.9xʪ���bN0��f�v��$6��!Ăͤ�Ci�8�Ă��!��Hv�M7iq!ąHt��R
C��!����
��!�C��M$��j��C�����*CI�H) ���
C���8̉Z��V�Rt�x��!���$�<N�:d���C�Ci$*LGt�����ښ�RT��ʕL�Cj]˝�ul�eAt��!��Rt��X��Ea�PY��)�G���Xe��3�ˌFi��������6��4s�M�I�1e,���(���@�40��#YU�bC�*�ć@R$6�XCĆ����E�VN0P�<aQ8�6��,�T�TP��x���t�Ă�] V���CL1�yjJ�f$Re��VJ�XCl1O6�y���1!����d��Y�c-j�)�q�%M0��!�6��ҁ��$:Hx��C�Hq �:a8���Hv���T�V�k��g5�@�!�C��C���C��I�H)�4��4��C�Hc� c	6$bN�:HbB�6��B�L�Ӵ
�ąHm�N����V�Q5q!R��i!� �C��i
��C�!�!ćI$8���
����^f�]���
AN�*CI
�P+R
AH) ��*AN T��R
���!�CI��
CI�1 �d$1 �H!�
�T�Hoxu�]�v¤��R
T
�R
AeI�2�R
AH)� �*B��ԭ�V!�:@�5�M�V���S$jҒ�8��� ���R
G+D��i��fi�Tf$�����X�)��\��f�hc�RQ8��i!�m���J�,m�4�M��T�[�$�T��XVV)Y�Qa�V6Ɉ)1 �D*J�j,^�$4��q�)m)kƪ��8��IP�*m�8��8#6ٕ�Q^�5<͆�]b&al��bQjB�;Hx�x���8�S�
�P�(fˊVe� x�u-5pQr��T:�L�q�,U�eV@�eJʼ�v��[B���*�jj�s)��,PSL�I�j��D�e�ƱL��#���VZ�0T�T��p�ր�p�����@+���[�z�sY:]O:��!Rc����ACn��m!�ĪE!�+օ���x�bZ,I%��[Un�b����*(zʌt�0̫��SV���`��TzB͎�GI�Y�5Iuy�u��:��b�ڣ(�Z�b)J270�i�hqqq+cA)�GQ�[h�K7���B�S����0�I$:Hq ��q���!��C��i�:O'jcb�_(��R�jZ��y�kSix�1r�(�����:���*+-��ZUEm(3]�1�Z�,�1S2�q��)��J��S)�`��Xx��i�M��I�zaX��oĚzt�*b¹+�1z�k �Fn8 �1�L`����ek*҅�92���c*�h� ���U��B�;Ht��!ći$4�@�)�.��.����� e3!U��dY�V8,E����`!`�I��L@�i�;Hi!��!��ov�8Βv��Lh��$8��KǛԸ�j2��WVQŖP����W+w�7�M����TFv�)ݠoV�f��FE���+R/+Rc4���0��v��I�v��Y�C����Hi ����H�:Ht��j���FҌ����Q�DkKjv�L�!��X�(�1%W��TU�P�*�*]�bӾ��=� ��-j1]&e
# ���3
L�"��ң�i�6�zJ�f����I���3�ݺb��b�h�N��ˌ鐬�d�J��@s�}�`���h��q89��U��/�[�{���ؗ=������z�}c�=�}��Jå��;%k��v�ބ�۴�{�pÕg߷sUy���W<��?��+�~�s���J���e�[@-��-�,�z�J�ol0�̮�U��Gw����www*��旺�<���ow�9�mu�dx��ޮ�[d�����L��ˢ���6U �ר�UVPU
�m�����]�����Wt�
����9!+_�e��\����j���6���i�["�AF��v�$�?�r�)]eCj!Ec,��E#��ը�J�,n5+���X�dPj�8@dn������ូ�v�˦�o[�x<�������˴�թ۷���n�D #j�?I[u$���4�N�F��v�(�I?q4�
;"��&��+U0�J�t�������E]�H�u��82��2��q�HUUC�-ۮݷ6�{;g��*[�t*����+�������KA�J�V�#�����o�6�[v!��������W��U���(�Yl�$R_�����2*Ki�Ԉ���+!�6Ӑ���5=ou�֛ٽ�zX�`������U���B��
����
�V;b��� ��7"�~q�ݴm�8�Zc���͐K �n%��*d���qHX��r�aA���E�H
	�KGJ[jo��5*Q��D���q(���!�ح�[%3t�ηK��E�{��=w6޷=�y���wO:˷r%��N��;[��!�Q!Z%���Zu֝DE��
 V�8�cg�@V�Ug�\"
�-j�N��=�뻆W����׻��}�����ETl��;�p��4T��R8��? B�UH��D�K(7,VK�JۥiƂ�(����;o�t{oL��ow[��պ������UT Ul*����    �UP U@ mSqU @AT ��ř�ݽ[h @�*mm7Z�+[`  ��TR�@�@+*�  P +m���m� P�P*� ��*�*TT�� ���
�UU U*R͵
��ݲ�EP@    Y@ UVڗ1T���  �U]ZU�Cl� @UF�PS� �  dm�*��� �V�ۚ��Tm�UT�*sT�lP`sp��@����֯Sl       m�m��;t*���  �T�iUqq�� 
����q  K��*��U *�`UX�Mm�ت   ��~Uw el��z��@ VV���m
�TUU6@ 6-�^����/P����ݶśژu��     Up@    ���l�@  ����\�ݪ�c6�-��U�Pp�U [j� C��V��@   �      *�UV� �{��� ��� 
�  .` �d    U*��U�lG�  �AV��T@6¨��̦̊�R涶*�@�   �
�� U  ¥�ʀ
�   Skj�ujR� �   Uf�wYܷ����Rr̬{      m�         6�J� �l  *��    �
l  *�  �sTU�*��~���J� U      � 7īl���� ŕT       *�      ��     �  U    V�   T �@ P   UUP R�
��~ @�@�  @  @UT     �P*�  �  dݛ��r          P���u�{��[�~馾����Oum�m��� [=�]��m��fʷ6et����  m���nj��-� [6�P  ���T-����QY�U-�ep�ª��
��  � ���˻w{km[[yl�D�=������/�̶�Vݷ�7���w7�nݏ��� 6�Ϋr�r���;���%@on��K����ww��\�l��6Ǫ�� UA�J��U@  VɛgqY@  �,��T+(Wu�P��6���l�j���@ <�V����n��:�w~߻�ʷ꩛Z[�m��P�6ж� 75zU
�J��u�+���޽�2
���`�p��?Wꊧ��{H���YAT  �S�*��_���B�U�� -�PU e   T   U+m��  LP ��ml�'p*�n��[;�n�Z�T��l��
�]� �U
����rj��ܭ�
� �*�{��eo���gt���n�Uq��d����M�*jG�5"�K[��|�w�k^�������)��A��e����f�ޣ��V��ܶm]�]���k��;����j��c����q��7E)���ϱ�7w����wݒR�m�Wjk��� 6�r��[�;�/�N� �M�-mةX��H٠#�zL�'���w۽\��{�rGp�;�<�v�u��ٽ�ԪW�m�í��p ����v���*n��l�e�xVA��ڬm�F�+XUY#��4*8D���Jݍ8���~�wswn�Nq��2��5�U����[d����{;�R�s���i����2Gv7.����m����n,�,�$dd���("9�a\������*c.�Խ��mq��pk�f^�ݘ}��m�=ɷ=���ݹ�%{y�[\�1������z�P
����&[$ ܎R�F�CM��
V�+�	���$�\�8��u�b��7<��^5�����ݶƏ��T �0�6?̕;!.R�=���S�[��sUM֝�R��%OwV���Uݻ�1�����DƝ��K	�ݲ[�v�;��GN���{�U�
�[����[�gF��A*r��~rRX�P#D,�uJ1�ʥRI"�Q�ywUw/k���=W�)T�u.���v��mP  6���~`�,lVK�v�co��{e�뭶� +( l�U\�*�P@7�Y~�? Q�@p�
���� �m�-��m���j�N�S`  <m��P `  ��   ̀ �T����~    ]�� �� 
�M��f����7��m�U� 
�wU ���Pn�������J��P�  U�u�  )����6�  @   gn�� �           AT 
� T  �       � o)lTT   *� ��T���U p�R����S�      T ���o�N+k\�V��[fb���sڣq@�P 6(@�EP
�m�`�ŲĪ �  ͊ps6PP�gXP   Jl *�l��YI���[&��s-�l�P+%* c [���tϷcg�ՠ               �          P            m��  
�                   *�    @;�@����Y��U    
�  �     �            �P             x        
� �                    ��ܪT� ��    P p  
��?  +(�lָ� VR���W��*��   � 
�����Ի��{��  ��B�m�
�b��-� �7�          U    TU�
��  �]Ք��
�   P,� VuKd@ 6�    P  �   U���m�*�    �=�  ?��                  
���z�                        ��   ��         p *�  �~ U�
�gu                        *�             *�             P         ��U          @ 	�          U�           �    6��   w`          �ӕj�  \�� P��v���� [h*
�*���T�U*��M�Y@� *T �m��  @*��n�s�WuR�        �U �m�v��ij�m���� *�*��j�@=ڨ@U�mUW�yݜ{v�  �<T����d�i��Cl  
��w�k��q�               �*�         ��v[ym��l뫲�@
� �l�����Y�;� � 3�����Zd 
�         {�klolU�U       T�       .`U ��@�*�  s�`*�atU��簵��շ]k5����� ����n���o�������������r�XBB?�?����?�����|��v��Y�kZ+( �*���Q����P T� U �e@
�� ��*UTT�����z�v@ m��mU�As
�m�PV����ⷷ=�PN ���d m��@  f�J�Sb�� -9�T
��pT����  7
� U \(  ���@    @ *�w �-�T  ��@ ��Y�so����P� ��me*��7{wm�]�{gnC��������@�gT��M���Y�wU��k�x��wv�^� �m*� �^�eݶ-�]wot=�M]����{wz׻e9�cv�w:6ד��E��ٺ[��1��V�d�:�F,���.�ot�m��,y۾�l����tul�]�y���z;��=6w�N��q���wt��k:��m���l��U#j�ݯ/M��gC�û6��W�M�6��u�����ow�*��*�8U=U��]��ʭ��-A�)N�{l<WuClU U�T  @  e �U[@3Jn'b@��Af��� *��.8[k�  *�   P    ��Sj�UT@ �    <    m� UB�T��
��p�6m�  T+%@�T�� U �� UU   w@    �P *�YM�    T 
� T @ Um� �� �VP  `�Q�@T�ح�
��{m  N`.`+���uҕ+�   @ ��R��(��P  {n6�  l�� ]�we�O�H$Y	
$�I��G/�U*Tr��[��lM�,p��ʫm�k��l��n�*�� �@k���:�xiס|Ʋ@�d�i�������Z{��ښ�6�޾�K��^����]o;��ݻ�8�sgT�(j�m;���6��UT ��^�`T�Sa� ,�`
�E�[hV�ͻ��*�ٲn!T=������ڑ�$4�&����$  $�A @8�9$/X��s������g�-0�H�whv;�{ ����il�:2	���X�Z��P(���`�޶/z-�;�t�W��n&]t5��SU��H`їj�u�2��H1���y&RA��m� ��ՍⅅxXн�����T?�V9��ٯ(JΘo;O3��8�z7[q�`ZJ��u��w�����c��e���;���,u�4��Nj�5|o�^��ݫ�<���k���:;h��*��{k�x��~���|���x���2��n-����h�|�xKh�^im��� �;�v�����y�ͻn��� [*U��q;�;�]��خ�O���,@a�ʰwPv�<m�]tp(����LT	��q�{��=���?���cf�������Xp�^oX���yv�
��'
�4�ڼ�Z��/V��s��=��G�wV��7Qڈ�5�\��e��`�%}���*�>�Z@�ʝP=>޸�)/3���	Zv�I%$#��k�y��Vs�l���3���{6�ΦF����Eal��y�Z@�ᢽ�g�*\r 64�ƫ�xx�����JEgK2lt����d-�x��X
�O�V �8Oye3�3�!����B����N�KH�Ҙ���c�h��pn����%R�x ��OGB<1\0or�0��y!��W���,��@��;�hש�uֽ��J�of�v�SmT
�&���nW�����w]�Cؿa�w�	HY1g����G��a���2�a��s��ye^�NLq8;>� <�m6�$6ۮ�@Tɖ�A~1]x�ݪ�+��C�y (9vW�zS���0J��Sx� �Ѣ�-����lS�o�Q��ˌ��o�z�� �#�t��dݮ��	h����W�@{��t�NKO�Efσ����~S}'蠥Am�r�ZŤkYDQ_�)�t�՘k,�a��px�x���?��q�Z�s8;Լ��
���Q���hX*�֚�۬�귏�|��к�N�^)r��n/���+���{:a9s'=��[@-��2�eݍoml��������uUof��f@�mu�أ��A�m�*�C���^�>��\�M�G)C���2蘃Ժ/�v9��u�18{��]~��Y�"J8�P���Yͯ:O8�9�@X�Jq�:MG�L�1�κ�[�P������7���>��r�٩; Q0����8F��pE�|28�JK������e�4�j�(^�q�q}���a���o��|o?~׻{����h���T0�<p�[LZ韰�h���х�2#�w�p�Ͷ�D^�|���{��أ�{n��㐤��FZ��O�Jf�0��\k�R����?�ЋB��r��1��Qw�5���GkW��w|�zP$��7)m��#qV�݊7s��v��QP[* ��������7@PJ�~�Yz�KCzk��q���`�00����m*���Y���X�Kcą��]E0@l��f��SzW.� d8b�u�q�q�3Խ��!�^�����c�Z?�^��LRh�m��l&�!����2d�b@P��B�'�u�Y��5�o�)T~��z�3{�T|jf�AR�A,�H&�ALAY��I`�M24{vT�o��H�ƿf��ֺ��gYV�#O����;naƸ�zi�|�]
7@%եa`�ώ���'��úTz�|l�	�)奣X��Ƽ����1�����7��Xw]	�����hU m���m����B�m�����ueP *�﫽56�=m�E�UK%����P���~��ܕ���lv� 
��^�����ߓד�e�Ю����2m� w-��eOTw��J� *�(ح� �ز�� �UQl���m��ʮ��ـI���B�1��5i���n��Skh\m9��R��9dƋS��}?S�4k�g�$�./�|}i�Z�JE���Ê]{$i�u�'V"�LS!��`��ٖ7���g�й��)]���WO���k�~���<x�xRH��"�h�
n��X�M�N�8Wi�q~���nx��T7����?�;�)�$��p��$o��t4�.�M��d3n�rO>��s� �RiW�|Xbyɶ�%�����>hnJ�_�����k$g&~0�{���a�T�m2S-W���j�w���Vr$��g�?$o	�H8�����ó{/�hAj�5���7��uW[�m��ܖ��G-{����;M���k7v�p�R��Ŗwm��WuR�P�)�5����0ˏ�?L�q[�N�Cx�i��TF�o8�,�����<��$���۴-a+5^�q�{rɇ(~�,��Զ{/�gw:I�;-M��Ѐ	�]�(�Wabr�j���U�H:��fE��fE�<z1	��I��-/ݨ�P�+0.�pwg�L��T�D���n�b>�W���xD��A�S��وc2�h�JE�>��>6h�P�S:���� ���MS�a�&�ms�X��ڋ������J:r��	��u;�T���,����pX�R�vZ4�@�Mc�ީ��ˈ�~P���05�x�|Fؕ��"�Ly�\�O5̋|��l�m
�D��#�hol�]��e��p絥��*l[  �{�\��V�]�R�£�2!�9�Y��1��ٞ˅uP����g]�:���X0Q�F�M�+C+;�8S *h6�m�N�W��V�f�״��}�28�L�T�=�[û���ď&Gu��u/�3@�Ki �X��+%8C��9D�ݎ!��M�n��K�l���42�G�U�P�5��E���s�+&���m�i5x)�[�Ϩ�h�n=}���w��`l�����#�QRB�TZ|o.g:y�!ۇ�>����̔u�l�j-'�쇷����T��g������o<| �e��&���<(�ŉ6�h"��{b��W�j����U�ѻuܨ��N[,�Qu$���;��Ai{%~k�����B,�G\NSC�!����B0��w����!j��$���D�M�tS�!�F�A֯���֍Ý҂p� ���Ө��-p&_h�cma}d�DNY(!M,H�@Q�u����=�}�	�B:!�a��T���ކ�a���Ԗ@RU@	Km�2.f���}��K	�<��z�m�0zf{"u����z�8��{�m�%J�������t\xםZ��y��%�X�ZX���*��U�<0WWf�c�x)���[ح�5!�bO5�����K�޵�h��wrZ��H�d����w&�w�5�y�]��emR�*�USm�l[�m��OMOU��k�;��+/R��LB��<��3�0�j;E���ZsY��SD��e6[7°W���t�B۔�B�������^k�^���ss�z^,#��Pr���UKT&��>,��g�x�zĮb�`ȌYtc�x��Q���ܴ 9�NF�����-���^u�҃�� �)b9ܞ���^�<�yM�J_����<��Bn�-l҉b���o�{o��]�Yz �+���ydV�d�8��C}��0CCˏ�՗�c=��qA�6x�V�Y=.��-ō��%&�X۸ :����zkv�U�n�������
�  e�׻A�fǳ���@[ν6Ҡ8�y\ٻn�̾�.�ڮ�ͧz���v���m�Kc��U 
�csT��Qܪ�l��UT �� �U �� 6� w3-�J�;��_����P�Pm���ɽ����M��電�����ۺ�����*�5�j.v�W4������������dLC>,�iF<FR���"�ʑ�>I԰=5q�a&��K%"Jo�\>w">�;3"g,��rg]8F4�dM�~�m�O�~��͔d6�DN�u�?{KCIa���9]+7�	Ъ#F��������}]��U�mw��Ѱ�KB����5�iY7J��T��
�:��t^�~c�V��B,�,;�_N疟�?�������E7�������-��]����.s�H��fgK7\�3B�LC�q=��O���~�h+����Q���h��������ꜫ�����[h 6*�Ͳ�m��[��Uz��qx����o��#<���Va������vUD�[U��{�k||+��l9iU 	G)W<s9٫��������d��Y�w�x���t�	U6?��vQݽ�ü��޷����)�EM���?,pգxSɱ\��PՅ�iF2,:j��!���ک�� lq�}zk;?Qv�k�V��ֽH�[ƫڽ�<�ӛ�64Z2�=��	�9�X��	�6�`�%�[-5|+,��p
4m]�����`q�z�+���#յ�������!�e\M(H�\�N p�ZI�O�箇d���+��ɣ���9�����pCg|����s�l��~�(E!@ � z���7Z���ծ���V�;�Pf5VY�v�ڣv��,$�}�:�N��c]隸�di��3qS0���Z��ȸ���|�l�؅(6��i���U�Ow&Y|eJ�����D0�����_�<C�]X���f�L�j~қm��Wr��j�j�V//ܽ�w�Êᮾ�y���W����U�� v�`� ����!В! *����I�H@�I	6�&�o�@��$�N�:�S�^s�S˭s�w�������Wҡ�m&$%I&�R8{�wf��oL<Hi���9���=��Ri1�
�����$=@:H�a0�x�i�N�R���{�lOk1�{R��H�"GU���J���=�f�=���{�O}��IR;Hiz`@턝�
�i6�$��=@�C� O������q	4���6���!$� H]s E�������	�	'����@ P�M=0�,$��$�H�]�y�z�s�f�Ȼ����aP+�����8R��*x iз�n��t]���W���vL���m��Ӓ�(R2G-�X�Z[���{k6�=5�G]ݾmλ�y�j����z����]��|mַN+�ӭڲ�e���{t~��PA���b�����\5�#G�S�&�Bi�D���z5'���o�'�λ7	�I��&�:aS�Y��f���{�J���'�ǌ+�T1��\���N[�sYsFkY��S�AM��Sy��ε�ӣmd-����}���L��C̲
bT��u�V���-�<��X"���ޛ�d=�LB��<aS��纘��H,�ߚ�.ï}�Rm6ȥH���m�������Ϊ��t�L��˗.�q�-��+�����)��v��ur8��c!��8��z���\�d�:�z��!��H)��X(ed;�s�܂��*
mV�ٌ�V�0*s�zj�惶x��@��,���v�
>���2����tW�P*��������s��k{r*uUe 7v��퓶ݽ�n�{���x�L�Cv��34�����8��k$��Y���
���1�.��Z܂��+,=f2�AO�{���sΰ1=aP��lr�}l��07����l�u��kheT'Yd����*t��}}�WZti��Y��5�����,��0+ �v���A����ܚB��95CH)m�����ՠm�;�4��*�Y�:HT�Y7j����7
���L
3�C��7��aמy��;�̬>@�;I>d�|�U}��qֳZֲ�5��i�� ��&�|�z����'��I��ԓ��ߺs	�|��}l���T���
t�טy�_s:�W��O��P:eC.���l:�ߵS��g�OXVOP=�"����В�GKm�������6����9y��Eњ�ԜN y��t�=Vl�ie�= c
�����9�߶���nz����.����tʂ���>� ��$}!�Ғ�`�>�̺�����1��Ӯzny�=aY6��[ �l
��s�����m�ֲ��.k�P=cl��C�>`9N�z�}�}���$8�Đ�yy�̝�y��o˷=I:@��j�d�7�d���xh�y��膐��N�N�T�O���z����q*�
�V�Vm\����n�;� �R���wm�ۭM�o
�%�^Hq�� ��<aX��{����^H��YRx�a�9�M>�~���~eOXVS��@��4��j���_}��2[ ���11:aS����yï����/��m��A@�y��fk#�k�e�Xf:��܂�$���l�-!�T�o����]�4c1���=@���aRt�Y�M�����B�I��56�{l���ʓS����bd��_k�>��oZ�t�Z�$���y�w�6�][�֍�x�>��I=C���N�����L��OXM�l;OY5�Z��p��z�]<����k����C�14 c�1���9{��W�}�߯��+'2�:��x�H*nOz��9m���B�~Q�K��?�U'V�,����痻�h������߾�p�0�,��`Vt�����������d��$�
��*C�d�*s�t��_XT2�5o�a�Vy�'n�}\���5�M2�t�}��~�km~�k�vI --5�m~_K+%N�@�ޝ��o��i�^C^�V>O�Hyl6�����@m<@��eq��R
z��q�aP���4��H�~�,� +s�S��yO�|�A{aP=eC���ޯN��~��������T ��
���K�4ۺ��{u�S��{ll����   � V׳��<����fzۻU�lwg�����ekk<��y_os���=۶�����m�]����F�d   �.aT�lwS��;�@�*��l�P T p � � �PU
�B���_�-��mm�<S݄��UU�@q�=ٕ��˹�w�w]eݩl�@+l�ػj���3x�ֳ�{^���Ad��:�����_���N�Z�& m�'��S]�1�7��7��J���R
|�P^�T�'_g>��0����t����&�)YY;eC�}��a�_\&�*�
��*C�@�i��?o�ˬ�unff�����8�`��m����:d�����zn�W���
�}@���>��s�� ��*�
��*
O���� ���1���A�����Fd������G�A �	���%�yQb�<u7�c,ŀ2������c)	��A�4Ãj��?Q$��N�L
q�k:�u��֭�fjᙙ�����ȱG�=冐^#���K��j����P�=C=�kd��0X,�2�9i5��|l!�_XT2�ߔ�R
w�={ε�,�2�2��
���!O/=���#\��;7���$;d�9T�hFk3d����aP>N�Hwl�2����jO^0X,�eZM!S�&*v{��²z��aXu������&}��5�ć��SlXT��T���vw�I���`�z�œ�d�*k|��Y���u��� �̻ܛuޖ�����WwA8*�m�i�lmXIT$,����Km&��*���1!��'N�u\���T���S�e�
�����M�0�H)�(�`�q�!�sν��t����0���;�|�S��y���h1��d핞2o)��OY:q�����a�.f���i���bC��S��`��|k7��H{l��?}x/�V"�=4�VU�[I:����ۛ��NݯF���m�eִ�8�@�ƽ���q
�Cԗ~��l���@���T�- ��y�M���l�- �;��4���4��'���hwH;���ҭ&��(�����v�J;,����!�uH)�T`�eI��1��;��|�aߴ�� T�&��bC�d�*{���
��m��aP�)<�Ɋ����|n�T�-�S�h�`�gܾ�[8�~��V<��:�fH(�)$�J������(0aUf=��󗅿Ha��bڵ7.��F5��Ў�Y���i��=&��X�-��KF1^~���̋��ɝs�h�uWu7�8G�A9i�-����v3�����l0v'J-�I$�<Jx�VTk�1�Os=�i�ͷ;���� �
�[n��$nЈ��[$�?i7"ƴ���97����ïL����_��0��;~�t����~�w>�o�����h FĊK��d�מϜkQ��)�*G���0	���P�psyc\�?d.ܯ�Gu� ~�Q��Am^�Zx���b��y<+�ӡ��5l���������;j�y��sap����Lǅ�*��$!��)d�Z\x�ɾ�u�T�*Y���O����׳{z#�Oׅ�.O���CV������3�"�̐bR���?KQN��0h��/N(<�/�`�n���>�T� �.��=p����$������=f�N����쭪w  ��[�F�.��E�.�(+�7��	��b���:���(7
�S%���K(��	$T̡(�J�3�
̀ŸQ�R�	�+'� �"ǖ����51�r���hU�����3P�y����i l��~g����%@|Y���#Nחv8�!R��!"I��G<�٤}�q�y��l�ȆE��yg�-hb�
R����f�p��ai��d���j&���D�~K,ݘ��g���qo���L����#m;Ns��<u�Ֆ6!ƚ%�c�<C��qD}�a���3���,���a)�e�h�("H�����d`��JWs���� 6��!�ѱ��[r�")�?�5'p1B#8��T�f�2Y���U�k���G@�O�5ϒG@���'�^tk®(�Q�V>o�}�sg���6e��E��Ϋ�Y�0�h�s�(fs
��t�߷4{��J38 )���IIF`6lCf7u7a�"8u�	�Q��y�̣�}�Ɵ��}�y�c�o9˝�my��3}	k	T�FZoՋ��� �
�P6��7a�Hb��^8v2%�<Fޡ*�J��~��q3�$��o�i���o:W!]e-��¨��a�F�c�4�\F�+��J\~�!��}������v9��R,`vP��V��F���������������
�6���Ɪ�<�m��e�l��wUQl�   �V���{{}�����Y{m떴�U*�̥�G��l���N����s�w+L2�n��m�{��ޜW��U Ub��TR�h��� �T�Q���R� �� � �*UTU@�z��P�m�����*��3��G�~����y�9i{�۝�-�� `�U��^m���(�VX�ب�{o9<ձi?�?���pR��|bB�����>B|������}�s����
�%� ��vk�zY�:{�qUeS.�1��Ql����`]`?/.3���;,N6�]���T�-������>>�PH���'`F�O�xNԸ��UCC�{�1:�ԁ�(pB�b�;��q���3S IH)$�k/�3�w\]�Tn������c��)���Ӕa)�;��rӹ����g�r��# RH
!�����01�^r�B��=�{)��FZ���]��"[�Ӄ���o>�!�Z铓0�EU������{�ջy��˾�꫺�m����ګ��VN�,�ZRQ�
��N�E������?����dC�{X?|��f��>t�C���Wj�^����S�@��������B��oz���5��I�mj��'7��׮�)��ݗ�2F���]�ݙ���6��ݷy׆��L0�%�N�k��yu}�W�:�H��ܺ�{�����W�t��B���X�&� ǗD��1�tG�M���j�c==���9g�������ۘ�������(Ye-�z_'�Ϛ�O�\ ����F����V"z/�C*j���}s͸1���ND��q�S���g&�Ϲ��7�B��Ѹ�<�0�=v�m�V@��v9�D�s�G9�����[���]�xT��։��.��b��n՞�����k˺0�@lm� #u���kT�$(P`�oorh'-F���͏�
���x�l����F��v��ޗ&��������.P BR!AJB��l=sო� i4c�5FK�ٱ����GUŶb��blӃ�Pn_�w�V�,}�����$Y)�����:,H�f&��� �;�Sfx-ݗ�Z6_��o�E,Ţ�������x��#V,��-Т�������.����*��U�j�W��h�Y��Q�x@�bm5	�(�i-l»��5����6��Uc��ܵ����^Y�.?e�ñЋc���pGq�OF����8��:��� vKi]�Z�ۼ����z��]�۵ܲ�� .`�U����s�]Up���PZ��ܟ����ksZYgZ���*��k=!+�t���=��z���m����C�E6�e�]N�U�WI���F҇B^�sv;������o�o�w���n�$R2�i���h^�'f�6bxNY��N���py���_m�*��_1~س��*�4�]�K��% ����_�'��o[�&Tkڋ���ib cY�����+=,q��C
���D؞�y�޹���a��xG�H �J$D�1vX�	�5��υC�2/:�8-�\"�kS��M�}D���1Gs�܍��%�@)����|Ye���6{�黹�u�l� �[��mn���ce��%*e\��P^���/�����/�k�4�؍�����>�%\� !���;��3Hf����&���"R�ن)G;5l�������e�<7�~c�hۉ��@4t��̆�9DX�ɋc�q)�% 	2��T��4e��(��8F͉��Qp#�c���/Q}�Z���m���oN6YT$�ؐm��=C�Q
�q��<n�q�r�*�8E/LA��lw� ���}�֫c�bq���p����d�B�b�,w�:bC���-�����n�����P��7��twzg���@�$Y$!�V�䐨(M���'�`
I�N��l4�H3�И��Bm���4r�F���u�{�[o@?Q�C�~�������y�x�z�2@;d�M3��<BH��Xu���Xv����dw��$��N!<���'=�׿r�y����v�5 CI�y���B���t3�tɌ�+,	XN04�9�d6�R@4��2_)8��6�H,��v�g�4��!ى�6��Hm t�'o{�T]+/������!��m��m$�`��B���P)�6��بm��6�  6��`��P��M�H���z�*l��=l��T  
��T*�n��!� � �*��@ +(  U�.�  -�*��j�[j 
�
�� 7���  mP�
� *U 6��  � �T �   �      �� �Z������ʠ��n%R�KdV��xs�������v�-[kwd N�N ���U'y�-��Z�ok[W�*v�j� 6�    �U=z�d���zv;�n��ݽ�n�y�ٞ�ZQf7e��&2�-כS��tw�ֵ�1�-
춁I"�6�l��_nwgz�wr�����l ��khn�Cn��]lP쒍�*t;	Id�6յ���ֲ�;�S�7��wvٲ\�}*�e6ϻd/���~�mT�U=T�T����m��P �[����2  UU �@     [[P�U?�� �֦�ڢ�N�T�Qn� m��*T�k�  T    �     *s�~    <         *�U@@)�� -�T �*�  U�T*� d� B�T      5�    @� 
� �     @ ~�      l �  w  �� WR8�U��3j�TS  =��+l���UvH  
�?��ۦ�U�mF뵀 �f�@  *�Uʷ�t������������ 
̔��Wv��ŲMڨm���w�����U
�  *�®�P;���/j���?v��51BدUu��V��<7�Mm���-�Wy�v��n��(���l��M�YU@�mu�T�ue�m��m��UU 	�� U ��� 6� w [%I֕q��� z���SlȪn�����]��ܷM�{���+���8� ����ob�z�w���6!���u�R�dS0M�^�ك��΄���yd=���"ߨQc��~����*k�05g�ACt%� L{.���G=Q�s��#������Ծ}�Ȁ	�$�B��-�j?��f���_^5�<�z��>�b9���th3Li�������a�D�1��m�
$I)%4�?�Y\�E6+��5*�����ǯ?]�^l����K����<���]���ď�>�&fB�ED�(Cf�u��.��0);s69���g��ቅnc��0h��C8�ݣ��L���-������l�G$������ݮ��P m��V�;vۻd�f�[��"R��"����n)1������|�91�7 F�,���T�ʍ�}V߷�S��ue?2ѐ	k�B�}?0��N-����=���Y��>�f�H
C��ePT��(�Cr�В�ܔu�-
XH�rWc������9�@��	�5�T�u�6�v��:\����9�są���m��G�i��3�q�@�y?	��*��~R�ٿƁQl�ň1��=��^KSZ���d��� %-_>ؾ͕�̟)R�D�P%��ct�>�BB��J����G���,�D&�s머��<׉6W�e$PdS!��:�8S�c�@q�t�8�M�������a���ʛǲx聧���6r�V� "�P�n��0iٻ޻�V�m�w@ Sm�U8յ��Kkl��Ƅ;��L���/��W(p;�f'���e&��ϝ|<%�k�v���W9Ga��UE��=��5���ڎF�أ!���f.��W��H�7����Cf���}	#r�e ��%J"������� s��`q�9�:������۬`Y�R.�r'N�{)S�[1�d�TKW�$B1���I<rQ�Wm7�ѿw����&�E	J�z{va�	��zf�oC_Z�X0m:*nn�ٙ�LDνҠ���f�4$luQR�IB��y��Ӄ��Y�3�1�ӷ6��"8{&[����+�j��7��a��l-jI陘��^��{�m���Otyv޽�n�dU�-�<�Sh��E�������� �c���ц�xAt�L�:1���Nrf0d!N+�z��"�j�v�I)A)�$�@��0D0�5��ؼ���Hq��,sƃg<PZ�_H�r��_.f��C;�_Y�}�H=
A�c�T�0��C��tF�Fq��&cm�S�)��u7���͹�ϥ{�A��RX[d[H���}���o�qv�D�2�1�0��ܣ���7�P٦�Z
�H��_f��&��e�gYͥ��S��@��ѰR�$b-=�3��>�>Ǆ����{�N18y�h��Եèǯ =n��rM����؀-��Aڝ�_.����]ʾ� 6�T�P�wv۫���څ��v�������[������{^OM��[�g_m�+X�	%��T�FT����[K�����{n9ׇf6\sg/��\���2=7
����Β���R�SR��_U�y�{�OmI�T�Ⱦwi�e��:���~��y"�fPd��h�Ibc���W�l�M.�Re���RT�ܼ��h�3��%z��#��\bY�g��"$%)%%(�	�k�6�.~")�SK����w<��V�	Ovk~���Φ�,[�/��O�)��RS4�n���m;�˚�U���Uڴ�p*U �	Z؜4wy�7-���Wwm{e <�m�ޣ����ޖ�������s�ݽڭ���ג�v������mR�*��=��k�4�l���[%e<6¨ *�p  p �PU���W������/@.l���V�Os ܶe��m�=׵�����^�w.����v�[Y	,�_�l����>�f}5�G_��`*�S^�\�^���ϓB+n{�S�����c�fd�ԓD�\����푺��o�T���e�ަ��oL������@"�J!d�	D�n��N׃�޲龩�f��x��9��w��OkP����2�5O{w��W�	){��I6�gq���-�WD�:�ً;¿���s������$�҄���Y�k/��x��]i<0��ǣ�!$�S��q�i��J�'T0�g�o��Y�7
����N�ۻ�����Ϊǰ��E�P]�g����[���G�p0����N�Q�鋷�ȱ��]���L]��l8S1���C�=4�9��?���Zd�k[�~���gѵ6X����M�ɯW�Ȕ�e$H@��]bUjB�\��q@�5G#��	E"���Q�y�/���j|Kq3��ņ#Q��M�z�;���JF��o�k�ت����>�_��<��~�l��B7�/��S�w��
�㫭~���x_���[$�#�6n�6�M�q���u�p�Q5w������8��&�_;�e�P��`��[�禼���Ln§=	2��
�P�I����xm�|��Yf��\����C,2~r�b%�"Go_Kｖ��j:�ϵ�v0��PCm�;��K�q��ӹUml �-�Tn]j�I]#( 	�S[?�:��o��W�Y�>�؃�W�H3�Bjb%p��7����f�86�ݮ�@�͔#����F��+��sEG=��ɱ�]����b�m�|b�Ѣ��<I��#��*
^���{��y�<(o�k�ſ�w�kԢ�<ƈ�7�B5�1͚��Ь˓�YKm�S��5T�����˺//.�ve���i����'�j<��l��n��?I��Jfbz_[���x�ؘ�~8}{܏sS����{כ�:�������r�-��ۻ��ލi�:�y�m�m���M�ֺٵ��w:��ؽp���f����,���O�nT)ã���D�v�c��w��>1R~� -IcV�V���0��2#x}"�1����~���v�P�)G
4X�蝍�����{��2�I$�(�E��3��,w{*]R0d5(>0#
{���^9�4)�j���?k�N�����`�hm����^�Z�	���q�_hH��Na	��j�i�G���B��8��v!_g���r}�]��O�u�O�7��؝��������|#�s��8UhOI���L��N��k1�r�-�ܒ�l�9��D����c	-��ܒ����g���v��n�]�dⲕB;��f�m\������VT�!��@��!����4G�����%�=���G`�B6�E�h-����{����n�?�&�"��>?Y���F�d�2
�`�F��/&3�=��t�2�@�v��~����0sB+t��RS�V��\k���<
��Ň{4��<,A؝���e��UKV��X���2AK���S����b�oE��`�~��dS4��{�D�����1F�)"�$�39c��Sh����P�u��q#DSv��F<0-��72!�]�g���|�>��/6�m�ZM��n� ����Cl��M��Gvĭ���������U�����[6ޞ
�Na�d U�ei���v�ݵ��� ���ѽoCU���}gw� @6�pUQT[;�m����M����   �@ m��*�P��������UU� IA��FV���mZp�NF��ն�: l�+{{��[Vډ[�P�j��c�j98�����O�����R ٍ� �Gi��(��l�!ue����}��L�$b�8R����^lp�FF��=��[��窘C�B<��8X��������	B�Q�J�JG�G�G�>:]p�`i�6rQ���B
N��4G����<,}�{��|�"��������o���B��9��=$�Q�c�װ9F���G�aˊ#豿M&�Y�^�m���~��i�
B�l�[5��߾0~`m�A(��l~�_|UxF1l���u��0���m�ø�u�����f�:��v���+��*��lZ�u�g�t�.������º�БZ)���7��#��o8�P#+Fjg�y�ŕ�������a�K@@���P�3o���"����MA�EZ�-*f�v�%�I-�ȡ@(UTp���nYBH���T
�Ѯ:p(��º�ܣ��4~��d���GQ�~���ܟ�WI!ATW�m8�9�|�l![]`��֔�+ηゼ �}�n�߇���&��IM�~j�oN'Eda1��﾿��B���|J��Ρִ�f�]������ܶ��?�I�%<�ႀ��r�}1B�3$���d�6}�����;�s�!�8V�OzI32M�$
��lj�fm�e���wyY�B� ������8 ��j5���~=V|������rsO��R����&��h��j'צ�ٯ?���E�:t�ᡏ��EM�4 �&�?�2a�J�6����O��4�Y1��l4KI��l���a�AWj�e��]�C!_{��!#$���2���N��>H���3˄�۶q�CHi��$��HF ?G��.zg�Gs,!�˭�z~k77��Ǚ��8�H�6�{�:��I:`�d�l dY`m�P
��!�z�	�I!Y$�$�z�v�B��HM!"�Bcc$��v=l"�{f�:tst m$�N� ��IBx$�*i�!�Y x����I 2H@�$!�BH��!;d$8�q����I q$�@ Y$�B��@�	 �C����$Hx�(N��Đ�:`�$9c�ް�4�I��=@<a�4���&�iS��!Y\C�I�I�턇i 2H��m�v��J�1 � b@��$��Y׾��)�����Kn�isޕ�{��5hJ 
����?[#r�c���$p�f�Ǟ��r�^w�۽ʂ�����)#b��h��٥��^ww�M�����{G��ӵ��7+<�V�M���"�Ѫ���F+�ݤj)[�����U$q��Z�ڈ�QQ�����H%*m*�����h�B���~,q����{�ӝ�f�j?�|���ڵɍi���#aъ��iT��_^eGӼ�D��U����T�d��?6�*8`�I�1\m�c�̎+����a���Y�l����e�;j�p~��{��p
C!��Qp�=����>�5�;�k�E�oS�>,:+)z
���+�8i�Os��n�P m�JUwM�$$JA�-)���xϯԱh�,� ���<���i5�4#v����1�Ƽ��$��%(Z'���Q����)ň��wG1X�H��k�_v��
0���d"�R�R��1F�;��(Fa�^fP"���G]?H��w�ϥ�A	��a*��HYjx��n�9�*����w�%v�p���c�ٱ�B&hs��.�+��}����z2�羑�0ן�>��3J��e�,��T�������$CCUm�ˁ����f6\#����*5�"<̳pU3)�������7=���*��|�[�{
� T�u��+���aKm!B���ֶ��~��zG#��Y��Z�3c�\L��#E��Εs��s��z��@-v����1g�:V������>Ѭ�����ڐ�|�Q�D�:i��JEI!��������	g�]�H�-d�����e��rb��@��Mf��?���r�4�M&�%F�����o���@D��"�Do�X��>3�B��Z8H`�`t�c��ܭ�*��1����e������h�������W��4hW0xQ��o��[̽�rl~��]w����O+#�m��L�T�el٦�i���ب�`���Om��mP   �wm{hù�{��@����S��� ]En�vo��m)��]j���=��5�uW]��͎UP�US`��pT��w*��*���N U@ � 
�m� ��UU* ��6m]ն�V�˹l��T9�9.�oSr���Y�����j'�&�Yd/{�B�����������F0f��lD��H}3!���Ə_P��h������ m��h�	��Z?.S��!�+2�����w�YgO���s������?�X��x���$�D,��1]q|4X�x������ �p�Ǣ.ojz ͘���N�KZ(�,����t���2H��D������~�Mځӹ�3�y�����'����a�&[	��M���`=���ڜ%;������'�)_]��7���6�e�Z��.�f��u�m{����ݬ��@�-�Tm�j�2:���m�r�z~����y���o�=�V�s�V��qky����h!�SI��G��k��1~_�+�����p}�����Q���jR��5B�B�l��ꎷ��Q5ibJ�I����l_���cŹ�w�^7��0�
��92I%B%/�S��כ��]n���U����p�8�pڕ,��{H��(�e���P3�g��9�ޕVҞ���XQ)�YZ#˫���yc�}Z�;����澼����[F����|�{�����iG�Ĭ�2{�9�7w ߗ�{-����kdn���w⽻K�v���wk{{
�*�K.�b�F\�+)����?����k��V�V����<6\a4��ˉ�:�}B�nT��@�SD��%&���#MN�����utWV�u+{T51��v�9���p�$�)l�!O���{X�}h���O�O lw؏a��5�ߟy�����f�_w��{�ԭSD�۠�o�|8���i�@о�t�鎻�'Nf:Muz��OY��Ss.+��oj���gY,P��� :.���./��O'�oLS*�W+nWVa�_l�}{��_���*��@�ۛ��v�'w9]��^�;�Y�
��z��m\�[mz�F�F�W<�:z7���R�Hq��rx����e�*�  ���fT)�Φ�9���N����i�˻q�ިϮͯ��͊�� 68�}���X��s8dAEΓ���C7���7�X�|���7=��xxWS4&HGPl���J�X�ug�c�A�=΢@�Ǝr�kG
!�w&c�3nP�����jhC�B=�J�ʞ�y�~t@�WD�`B�I$�)b,m�C��9�%�����0�!Xb��8P�q��I����~�w���t�!�M�ꕵ۪n�;ۥ6��r�| lJ�����)P�u��A����O�E_o�4i{����5��V!c��m���:<�W�ux̑;��9$�$ `���L���#����9k�� 
J5��1�k�6k :#��4w7ބ&�{S���H��"v�@��[��?�ȸ�O}t�!�,�;>benu�E�~��1|bO��o��xC)MȀ1%3%%,�M���Va�G��uܙn�m>Bp�cş��3�|[�'$��9��y0lg�v3o[��(��M�&4�D�IH��WE�niW���f\$�� K5�/~5lӳ�W����DLxk1�{�S�&�E��)��
$�5W�u��Sc76�R��նۋ�Ӂ�݀,�� �u�Ǻ�'�l�^o���y�� [��6��v�[^��^�nZH�F�%�QA����'�{�͕��`  �U�e����ʠm�UC�
�e U;�  ;� �*��,����7���[{U�����Uu[E��S���T��O/����{l+��e�T����viH��5�`Yh�&.����#:�Mo���S4��4�P�6���91c��.�=ײ/ޖ#��{�O $�����)�"���SQYu]h1��i�PǬ����j8+:"�tlee�rj
�~X�Ͱ�M��M�24}�N\1+���+��UR�sS��57&5��{p���G��*B��H�R�s̏W��2�E��v{��v���]������|�s���rg*�^{@a�I�)L̙FT[}l�O�MhC��u݊k�#AG��Awf��9a��s{
������>��?�øU��]6��y���wn��2��sB�U 7w��J�� ��+G�<��ni����37Q�ci�B[sTc�"����}�X�4/^I�L�K$)	Qn���sq}�}�Jo�/ho�sm��~��
X�pj�['
�֙�^�|�绽���ݟ$�:E����x<��@��ԯ:#�ţU�r)�{�UT�mפx��
ffG�R��d��o=mM��OO9�c4
nf�b��/����ņ���D@,�����k������~nZ�^n�F��a�Mh�/Y��w���e�3nh����H���$�!�v��տ}��x���4��R__����o�UhS�9�S'+]oP��tٝ���w6����k������W��:���o��!#��q������~���nzc.w\������?�"�%dK*�������ق���q��r��j��{F)M{7d��9��|�"�@�m��D���:6/)FC��a�RF�z��F\�i�f,o����N�K0�n�А�a@��o��%/U8����=z���^t�����QE�IЃ��w��� ���e�R��_�P:'zښ�Ʃ��K�@��n���}��Eng�w��	��iRm���m�m��{3�yݫ���l T��m����[:�`YJ��_H����j3�����H}�K�H����oc��#�x��y�;٣Q��7���7����\{5�;�puk� �����f��Ρ�X@�����l��4�ߚ�J�t)�ZL�SW�?�hO�����]]�ܰ���1������{�����Cq��\�n�Z
0���ޝͣ�� �*Tx�ձK��X������c���?��j�P��7�'��Ӭx��ћ���JZ�)t���c�l�l�~�j�zԡ����{���`(����2�q��+�l��#p �mo�{�����n��ru��jۋ ��ʠ�m�imR�$�I2��Nt�y���һ�⯞!�aS��\��f,厸>�x�j����p{S'�J�$��$�N��mVi���5���G�m�9ˌf,p���*�C� e�)�n������I�H��
M�
b��]��\�\6]`�̏5�]_�t�7���}��8p�^�j��R[]�,��/��ÚZ�p�d����MpC�91��h���5;�b��G�=������{��U���F�����WLq�>,�V�r��:у�t�#�����1l��bZs]��F�����o�Ӯ]M4��f��D�˨tU��Z(<�A,��I��]u�t�#��$��+��W��YG{��ý�,{�����&�o���KGy ��������������` �0�́n�@  p�*��.cm� �[� � M�T*N�U��l U����l�ٵ�d��̎��*f�$ݸ�  ���l���  r]��*��6@U T�� �PP�[�{w;l� �@[ j�P 
�S2         P�@  @Un@ �װ���Y�^��묦��ةV��ٵ�޻r����*q�^�y�m�.aU��d�
���=U�OcB�*UW���N�iC��VP �   T�ڠU-�˙[��ݔ.��u����sj���&��V�s1ٻۥz͵��ʪ�]n�fU7{^��;�h��ٷ�n��u��^�N����ъ��\`�rA��Ԍ�[�U��f����i�軲m���y�]WW���;��m��i������Y��h�WV��*�܁���mk�6ø���*  �^������ m�  U *�Vڠ���� �M��@ �[%V�P�
�1y��R����w�  
�        �
��P    �    �   *P *��[hT��eU   r�@�� UP+( `   �    `U  ��@    P         ` � � s  [+d�m�m�  �r� ���Ͷ�Tζ�[�
�E��     ��ր+��6��� &�EP   
����P�Q� [b��U�kmk�̽w탫mm���t�U  
�S�u�uP�ƶ��,ڪ�2��\�w]U�v��w�X6�ys�ڲ�����R7U� a�(O�v���6�
웹6[`�S��;��UR�A��*�m�@�AT�P 
�T�
�v����� ]�l���u�tw^<�n�^�ݫ�m�	T;�,�Q�s���e�!��?0��K�i�Dx|ɗ���F��:8TO����!��X݂�I@L��6��f�,�d�	��X ���w�"��Ez@en�K~�,��X4\��Q��$�m��<�����>?e1��%���1��9ɳ�
�ϗ�9��M�O��-=�{`����Mދد_��7Z�	4����Q���t=��Qs�'�,CG��s-Uf?D�>�C� A�J�̨�R�c��C����=*�*��F?��t�������>3��W8:ɸ�܉i�[MPV����]xb�}���Um�q� *fm�idD�M���������ޟ����N6,G����@���Y}ٔ����e�ϔh��އ[$�?i ��B�~�#'��3+A�{�{^��:��4 m[%�DA��m���c�B7j�,�R"�K���3�iCc=��^縴�D�8>��e��:��j�u�/���Z����k���FX��B>����vF���8Ihحt�^{k�|zQÃP(/$y�.j�#����f���c�%��c���A�d#Ho�۞� �v��d�%z�[ko�|sK��]�)\%R�,����N'�� L{����P�s�o�BJ� ��e�E!��Tv}����mvVA�
�q]��ݽ��2��#X1[�o(��\�m-F�^4V�5�o�[�wrb8P�͊�B~�	&�$V:SH3'2#�>��}����e;��q�'�Վ �ج��:��Q�
Ѣ{�ԍ��M��y�J�ٓ���l���.��¡�
��]FlhMҪd#���ؗ[����!+ J�h##�_�3���#�Q�p�8�g�41�@�Z0p�1N�KDD������Mh��/ �l�P�n�D�a��)�4A�׬H���ߗ����WHX�:}�{��� 6g�+o��m�6�:�z��:�}��]B�R��*�@nwWz�]�{�ؖ\��ǿ����a�-x~�/+�_�+9[Ǎ~D�"�ep����X��Q3�zL��dKD�D)�� 3������K���4+�kG���>�kwc߯�ZU\.��#�)��[m�����>�C��}���y��-pb 4W[0;�C���Up`%�i
� ��˥���u����Z�8<{a��K-~�| ����u��%O�|�n�̻��/���h��62�@���v��ej6��+����u:[Z1��ua|t�\kݾ�<��Yf�˹#n����lh������C����w����w
�Scd�[[(N9����2��OЁ�mS^:ܨ��Q�1B�9��k0��+��q��E�#�����(���R�4�׻����ٰ>.�U38t�7
�,�㩷���*�#�HE$2T�.�w^�1�����0��IJ:0�5T���Up�$e����V����[P���^o�k�Fv�\�xϊu��>U�2��28�F�\� ��L������ǰ�Z&�������E����sK�������/���7�G�o~�x�������|�vc�m��m��I2n V�ڳ1�6m�U9�d;�Q��sl�]ʠ  ��6ǻ������.�vT�AWj�&�\��UEs��}{;���Ȯ���6�D* �����kd�x�;�l�  Kd   �  � �WuJ�������lՕw���\��A��}Tc��73{���U�v]��{V��sKt� ��WIi+l�K@js��<�ՇK�`<����\��>�t���D�����!���PĦ͑�m���������1�J��/�b���Z�m�[m�&Up��4xu�⠈��2�Z�|#~��!4���Cj���n�p�#�D��qBH�n!W�5}o\��n���v�`�yd�B��T�����]�N����*�L�	���$D����j����j��{+�{n�Ww��Zu�u���.��N������m��#crٵ�9��ۼ��M�QPU���j�{.X��u�����1���C�tIo�'bN{����Ma�H � H"St���wzU�ۜ9�t���|jK���e���&��*9*?:%���L	J"L��Gw�P�[V����_g��=n�-i��%�$��^U�/\�/��-�$X�t�[_O���r�����
��v[W~���G��S(^7����M��������|o�Ϧ�낾�C���DN*&RI)�$I��lh�A���p�Q�,~���S??���C0�s��N{k��:p�k����c��6�� �kC���������Ͷ�
�pU*f+���@��u����d��3�:1uP�ރ0�<�gO�S�i�#V��(��P���톏ŕ�=ߤ��i�hFZkҬ����b����+�h�9�ȮZ�1��u�D�4U ��	RBR�2���GQm1)�GE�ܗp�T0��#�Ն�����������o}*�=��nC����*��IjN��X��`:u�2��r����ӳ\�K��i���X�3�}@|xV��{j�������U$
�
Yj��c�c]��ӚbG��̠ݚ�p ���
c@�U}2V{{�d�b�j���q�Xck���?���s{m�n;����*���й�T6���2֝uR�!�s�>�����r��^1��bB�i�:,Pn�T��1a�^�(����U�5�#�<�2���I�f�U��*b�|�;��'�T�������]�mվ�2F�7�� �$m�wR|�`��f"��#սJ�#Qe�G[5�,����|ov8F�=�WRON�Y�R4����Jk�c�;�>��� �������#����ň�8/�nW2Z|!L�w<�`�/;��r��	 �0jRJ$-m�܎/}7���y6��R�s<�.��MGԞ3��$bd�x m�n-�ޭ;v���ۺ���� �(I�����h �P������ו�E'�{SJzQΑ��a�zc�XVA���?H��ʿ;��x��m�>���H�n\�]�wg%����3�DA$L�EHHJ�����8}՞��S���]���ܢe�0�'�g�j�
�u�I,���F�|��9�n���VI�#�������>�?����m���wH�
`�i����K���6���C�v�g��=�:+��c��ɮ�o!^��D��v�J�H�WԐ(`�w.쪣b��.c��W6��7���W��
��   Un��\޺�;�U�z�:n�T���S��k��n�ۯ2���77zݷ7��^�����;��j�ovv��J�UUQ�NU����m��P6ʪ�l�6�(
�@;� ]� �PT����f�̀UwwVQ�uR���������R��N�<ͮwE��z �sv��&���Ϊ�"$f;��oY�o�Y�C��kѺ#u�v��䥸���`t'�$�R$�H��ڃ��ҁ[��w:�CM:K�gݑ�ɑ~Z�O�oo�7���]�ܒ�J:�K!-4��E^_fY�0��=�1�*V&Lʯ��f�EY��}5������'E���J�`^1�Ɲ I����'����l�h�0��h��47aA�Ր=��K��t�*�Q���a��l�M7�-*���Z���ᬳ\�G�8+x����H�^m�{�R#D�W�J��+�J���n����������۽x���ڧqTV������&��;f��ߟ�\�l"8�2��8E ���DP��lZ�3��!��2*��$�P���iI�а֏]�\e	g�m�׫C�t)b��(_������ЖZFK:+HR���ם~�cA�)�dHu>?CDZ��6��kϋ9ٸ��+t�5���\��|t��;�`�4�S�j�Tf����C������]xR�xnk�!��.�B��y��}���&"�/F���o~���>�ِu��	�\���m�߼f �M�i$JiI�u��W�=4��i������lH��+����ۯuA������l�Rp ��y�wm]����m�Ԁ�Z@����6w���*���6���BZvi��"8:�8�������.�[P��mD�ޑ�����^�I��+m�H��6*�F���1"dx���44�|�S�r專�>7�Tm����g Sə� ����Y��^<���>үF�+x�tS+��C]���z�V�C�`�XG����<� ��Ɵ�v�s}{�/Ove2l����W�3���~6��U`;̳��[�C�}�u{s�	�V�X/����"�������%m~~���;QY@6�ݷs����[�n 
��q��G�^�
��������PC����deE"�R�I)+�D:�Dj(~V'�%TrT��+O��֓uI@mV��]�M(���QOԮ�	c�ݽ|z�ְ�ϯ=��_v�<��J8�i�A	�E$�$r�0_BB*��鐤�!|�i�-�y\"|c�~W0�wzfN��;�3$%$ B$�K��t�r^�`u�II�M��RV`CP:tt���3�ޜ���\X~�K�zD*]�I��	��M龧��n�f��`�ݝ����K�rn!{��Ꝕ!���&�I��� 9m�WiN��ǹ�=z�tm��Sf�["�����*����K+�ًJ�5�b��^�»�{��(�K��������㤒/ )*bRI$${��{ُ�K��.](�7k�=�o�F�ijy�r{�=���I�0�I��-9�Z��G��.���ݸ�n���������^�$Lf�ZL���9�ms�s�VT��}���vO�q�o]sN&�u��S�R��Wus�x_�{ca���(^ yAm&�m��}5�O�����
�=�}��t���<{�{�����J����v�����˝��nۜ��Um���� *�VKmp��T�(Z5!n}��fz
p�Zgg�q��{�iw�7�)��~����-&�A?�O[�����}��ֹ��*%*-sc��{�"+�L$e���m�M��=W������v�l�ڣ�'U���z�{׾�2E��d��h��2o���s��ue2�w������S�öd6�m��yyP�u�ճuVW��L"�m��o�/���p���]�7��(j���<�ᅍ����}�����Q��>���$�I$�I$�P�Jf��[������-�x���.ke�Wr��U@U ��Sm���/s�UEu�Zb�Ӊ��vc���ۖ�򮭻���s�%D��c���-R�Z�|����M���6��N�AܶClT�U
fD\�T �  ڨ�*V梪�ln�8�R�@�AUY�Ί� m��v�wW��}��v�R 6*�{6͏c��[��D��M���%�����_N���#�w�1�&Ÿ��� bDf�xO�J�-��4_1�koƱL��wW��r@�q��d1����-��"�Ǩ��}����ܨۘ�����2�P�@�xD��b6��Tn�x!�LƋn|�i.}�Q��*��p�a�m�O���O���� ޥ�d�ᖭy�֘ko�h��!�����i��x��Lb�ଉ����D>ǵ�w�ѿOF�.?��\N�@q�[M�a���8f�c����cY�5[<q��Hi��b|Z��X�����$J�oj��v���=��l�w*���� *mKB�B7D�$��۞�tXG^�L�)����H��y�&���lÿs9��ϻ՛�xrJ�%l�`S�_�I���Y˄5��&jy�@��f6����=^���;�mzUcT
 ��P/�����O��w=>���+��̮��8���LI32��D���ЖĚ��3~v��6����;\D�򦟷�]4O-鿫�#lD�[m���K�5�.��0��C�oMv�9~-�:�|)i�>"�v[ɚ3S2�^n|Q�F��듭���hY	i�5��������L�ce�G��, �^�ɚ�!g�+����^�<$+<&�3�3Jfe�2G�� ���:J�QDB7��um�n�5�P
��v��A�J�B�8]�W�}��g�0(�wX�N%��hT{aa
�q�=�_K�9�ɍ�p��4�2�
i�m]p�=�l>��.s���c�4ؗ��G�Q/�¢�!�!��F���ۺ�Ⱦ��gx�4�ک4����1���y55#� �_#K�LM����Lf�q5����ފ������d���0�޼�0.�i��H:L����H�~�����O����_�g@�7��AQ�lx`�M�T1�G~�G�G����k5�g����K0m�̚�|LN_Sve��{ָ9��E'Z5>����Խ��ד�g����m�i�Bmݭ�۷����^���wE{��� ��T��Q�"��Hp�f��>���<�U�0��-�/��0��c�o� ��y�{��΍6Z���HP�ޞ5�A���b~�
el[Wr�8�P��͑�GY�N%�g���U��Y3����v�% �IR���s�~�1��Meꁋ�Qb��k>1����斶��1�r�Lwn�مg��'�0��a��)
�W��T)R.�����`�u�jmՈx�B���/���0��|m�����Ueu���w�o)�A���='����U�:�V������3\!��{�<�а]�|6s�낭cG}����'����=�� e ��*l��u{$��{�wm��+$�f����U�V���^���&��%�aw�o��C-B.�v��C����se�>��2�TrdH(	D�)��88#�;(�5> R���ċ������O]OyЀ�S��E�%A+e�a�gV�x�z��;Oݝ��(�6����>j�f`�P;G`� �s_g9���6���x�=�5��E6{��jO������������M`�4�M4]4Zw�������S��r�F�U�B�wWMF���C�R�f�Y��Jc�	|Nc�g����uvl�hJIm��ݤ�	��w�ս�uP�P����m�J�� 
�*���c���۸���L�[�
�EB�JX4�id���M�&J��.��g-}��"�̵��(UU  'UUm�e��6�� J� ml� e�*� � �J��T<
�]m���c` q�M���=K7��+�:����]d��m!�0���1��T��Ck6�dJRIPDʞ���b�6��c�e���⡈C°�[���f���1��y�q�#<}��|x):JP%!eJ��Έb+2�Q�6χ���D�,��W�^�b�4D�vĝm��ɿ�zH��#��ʤ-�����
���p1�b�9:��ڠ�S�X�p�� �wWM_�z\�a�X���UT�K-����{'�M{��}��u�+&c����:0�X�M�p�Z�G0�;��,F`1[��s�쳡�0����R�P�K4�b����3F���4�Ň��4�p�x���ܳ��{�{Ƥ5���q-�d�m(x����+iݞt����{��{Y��U {�����R����~���׬��f���C̙ܖ�SUh�(��51�k�M[֤A�'�]�#����!$���YS�gE�1�Q�7�z�%o�6�$����jhV&:�rC�E�Q5?G%�"Q��V��g��tfn�lńq���H�&V,�ށ����]ȵ��vX����FKKcӾ1�
�R1[��m��#r�a��|�u�<,[�&ol)3^��$9�F�k��7��IY����>E��1JgÅ��&�;,F�.;5.���**��wwWi��BSu"�A�Ii�Q�jઃ��q]v�3���o�Ґ�y�u����Zp:Ώ�v��xL������o@�ҁc�@P-C8���M�6�wv�[��wn�U � �m��7���ǜffI3%(b�Me�s�6��6�qlՉo���Oy�w���W���o$@e���j*��|wkzY������� �js�J�c�t�bMI��On�u�ɱ[��w�~@`�)7tfR�G�qe� X�>�۹���b�2��5��<1�Ӄ��O<�g!�V�Y�v;h�Z����ws7���O!ZB���ڒUׅ1O>�e��1�Ɍ�)�F3��K��qS�3kϮ�8�uB���旲m�*��On����kݫ�S���5�^��bs�Ʋ���ג��RH��v�s�:�e��j�g�<��ӽ����ڲ��l�@-�ګq:t���w �t������n�7w$���u+�"���ڑY��L���߲$w���_�`�>�)L�B)L��,S�ښl�}�td�n�xC0�Aɾ�s�|�hd�wM�ޑQ�}�|�HC��I*�-an�����a�� �9�p1�pe0���f/��7�������A�sމ�v��d�\G��QH�TJ5E�v'D�+��>vT�z01�r�鋢�y�Q�=;۝W㹾^qۘ��X�.7&���(��R�	����:��:�Ϲu�ϊbD1�yO[h���<�*��쳳��g7�Q>GQ�̺�(�2��x m��p��u���-ݻ���p�E6
�:[K)mm8�T��u�׬~�Ŗu�s.�<p�p����+�?X�x]��ُaʎq��푂$F��̰��%4Km�ťw9W����TX��ҫ�1L龉�ƾ/�_�+�^��g,'
�|���xj��J����¨|lk:+����n��J�9Ni�G�̱��5��Y੍Ί�{��Z�jo�y0X%��J�)�pf+!S8d�"aUi���*�r�k:-é�LE�b����29���$2�F�}�/�>{�^�[����	�J@��U�$C���X�,1��X�78Xc�6���F5j�on�{�p3�����s���FD�lX>�T��~�W#<s�Bͬ��<�=~����]F�9��^ն�Z�y~�w��-��u�6���U��x�3켍B�f��Md������������b%Z-&�m��m�
�X�6��UN� VR�  �U ��*UUJ�JT�i[fŲm���d�-�[wU[Z�UK�R�UUR�����h� U wT�� [   
� J�
�[m��ܰCl�TTB�`+\�  �¨  �� ���       U@T  �   �  {^�s���۽�˹�j� *��%@]�ݻ��o(u�h��mg���M-��l *�Aub�c1��sk����w-�{�(�UT
�Cl+-����ַ���� S��u��w^&�݋��]nk�ە��Ԭ��a����ڝ����^�Ӯ�Ovy����v9��}��u]ݝ׍3.S�ua6��;{n�U�Öޕ��e�͊�赺�Ͱ���vw���1i��;�ҷ�R��J��	h�أp�(A���K̀;I�mTx+u���u�.� A]�Wce@�i@
�  �  �  UR�
�e��� m��e�dmR���*lz��[mB�*�ٶu��  �    T     m��    `  � �   [eUB� UU]� M���U    U@-�l  *�wU ��   �    �U   U@   �T      T  U  �  w  x  �Tl�%e�P� 6�R�  v��8[�M�ش��     ��jW	[��  e� U U*����w�ߟ������P 6��6)�qU]�B�9�V��l�����e-�T� �>��kk��w��UUv�ն6���;UV�ۨݔ�ʷ�9��v�3�����U�ve��볩��UR���[UB����m�� 6ʪ����d l�  � wAR�^�l޽��V��������U�V�r�TջmR�.mۯvݼ�� 0Tٶ��[e]h��"on���Ƴy�WK�6�xe�^,g�\�kߟM�cE���ܛ�S����m!A�]�E�A��PxVzfszf���,G�اep����y�S0C*��+w��Oyt��'_���:���Qic��Ea��p�"Ǻ�D��txOn�]��`ωs�jw�q,V�Bى>��M��m;������� �%)>������Ć��Q�lp�C���8`�i���7H���V�ߴ.���Y(�/>k{�|z���ƫ���b��3LR=��c��V��k��~�^���]kOݏYބ�rJI [i�>��v�u%�W�w7Weݩl�]ͪ�n�n��0m�	(�z`�n��\.�n9�bD1<�-�%�Ut����6u��5<�s�{�+N�P���;а�Q�.|���$����G��\���oWm�kY7ק�}&[U
6J8��,ɓ���Գ3���3��9�]192b�g���tЍW]hT�Cw	:i$6ۦ�f���8`�驦�<,\Ǜ������a�Y��Ǐ}�=>;;���O����<,�-
�m�5��\]���X�o�i��tm���hK�<���)���:k��d��˹�w0#�	J
T��0�ʛu��rٕйZ��޻<j\�S�t1�W:���Z��F�{�w'l�+Ҩ6�۵*�����۸�pT�*�n��Wl7nn������Ѯ��=���w�ӄY����<"_���щ�/��|hGa�jȉ�P%A�2�V�Ⴛ�j�s�*K=4�����)D�&8�8H�v9ǻ1���a��z&JD�$��18:i�'G���4T�k���͏1�&�ϢVL]yz�tr���S��.�,g5Jn�h�!��A+�.�l���xUU�|ztt�:Yϔerʱl��4�a�3u��}��^�5��'��Im$�d)k/=Xx��d��4�E�N����5���|�0��a.�"��!�B�Y����m$n� ��HW �!�m���v���� .T�m>m�p+�4�̔a���8��9/�Vg��KD6���ۃ}�ey_y+�|�0�-��E �3�o������/�nK�{-C��~�3&�b��D�k�A@B�u���m��f�󶙎6S�=N*����)��2�}�l�@��H4HM�s/�H�Tx���)I�紾��;ހܲ�����\\�o�;���h��~��/�7~��gOyZ_�" &[���뎙jl�U���~_M��s���f�ˑ3����~�����f��Pl�fۏRn�쭪w  ����ou�{��˝�FܙF:�ԩ����ۖ�f�[��Ƕ'�]�Fj�o6��vk�T$&QEY@&Q���$j�8Q�*X�1�/�ۊ�����9Z("nL��O��y ����
TH��m��`6�F֍I�6B�_y?�b����XgH�����b>�M}�>�����k-|5�(6i���n�^�k�>-�l6]��#7�
�0L���CP���ٚ-���3>��)���3���$�6C ���n�X�':�3u!��4�ZPXf����S\G�@nU�{j�i�ޞݻ�@�{M�����m���*U����g[mST�U�T��3lws� T  *��3;�=���[\G��*��\����kw�g;:(J�R��i�"Z�*���ɶ_nt6�5,l��j�R�su]�m�ܪ�R�8 m�
��_������ ���U *���v( l� )bUq�,��ݷ��l�::�uy���ɷ{h�*
�6�d	�8��� ��e�}j���Ah�>>Rc7�kE���Q��>!�[�&�����+I*8��A&���8`�5vW\�| �*��2�臱o-���f������y~v+���|�@�M��I�!z&y	kNH]e?̎,���d�f���eS�\ �5�X�+;����p�T�xZ@�Km�:M�&��i�h:�m��s`�0ia�&n��?,hW���,��ި]��)q�su��i��m�eJS_/��4t�,Lq��1)Իc�BZ�s?p�)B�[�Ԅ`�}&����W�-���[ �ӷ[.�w[vk���w@m� 'R���Ͷ񛛼q8-�Vp���-�	�Lŀ��mW�F���FVx��������6��U\��PI-�*z���5ט���z̘�� ~��ǭ����(�-0UB_�i���j�H"�vZ�l�R �% �q�����'.4Eng}8.�������z�=�7%'��L����� ���\7Ƥs��hq����X��
�T���g�BZ�{��r��}r�r�t)�X��g��{���V��~��w�#�ڃ�i~?nѵ<+��;Kuho��� �� Vm$�!���q�X�U���G�|��zk��#���Ά�ƈCFY�~gu������Q?,�+_|
��P�j���7N^�c���]�mvV�;�P
�kk��]^ڐ�����^qͪi���W�W��ح�bWL ��Dc�˵�q�K��Ώ�5�Y6�Aє(��]���a��z`��0��\|������b�p��F����H��W��_2u9��[-����i7�־*�������v����ث\S���r���C�Qe��dV�!�F��<�6�i0���oP���[�޼�RG�Á�z��|~W��� d�t�,�b�9��w�U�����+���U�T5i��������؇���j�ׂg�a����C�+��ܲ/�����U� ��Ok��m7f[�{Ew{��\Ų ���c�m��w���|�hx^m�:����uR�G	g���x~σ�e~Dx�����"���&2|$�*e$�"%S��Xa{&�1%�߮X�f5�^�g�W�>���]�������ͺ㟴5J`@�Jgxׯ����x.r3{{ۃ���l`�_�;o�}��#��4ϷĊʊ�B���������ۜ�nD_�C\�W!0m(�@�gt�2�P�7ċ��D��ɱ[��v�;����B���	JR	"H�2���,��Y�ˆ!2�٦$��}rc�k���'�c%՗}��CO��fj �K ��m8������i����4B'�ʶ�� m��Vڹ���VR*7$��m�-G�����E����U�����効:�b,1�[N��e�E�r��]��{�4�����Zh�T 	l��l�ǽ�Yش���y;�Q<|/��mTxX�;Tv i��ĺ#33��ύ�+�}ϯ=h2&Zb��o�H��/��Y�fD1�t��J�!A�	��Q=~�kg9���N5xx#}�J�Z: R�Y��kח{�����C�!��f�����k)Tp��:k��j�
s��JU�<4z>��_�I@�n�5^=r-fgYgvX�]Lt0oƙ~%��S�^T����}u>`�M�|vg�C��ƨ�z?�?��[R�� WM�s��wTm��Ⲷ���I�{���fP P �V�����������;��%k�����")Spe!%�pM4�J��!�N�ג�v�ٙ����m �s��Q�u��v�R�@����el������ �T��{@6��6��Sln 
�
mcm�������v����󺪷eݩ� �Sm�Vt�wk�f��V˫8~�ګ�_;p��p')��='¯��&�/yx�*Պ	u��'6'ԫ	� &�32]Y���nL+�)���%��{�u��Ʃ��U3T��Q �Kf}��۱w/e�s�e�ra˧�Ѓ�5�B��5Ѝ���|���Ӟ��u�����pъZ旾>=�ä��үX���:��`5����� x���OT��}����s���w����q���F��ĲJD�M���*���\��&�wQ�k9V8���*�p���~��>�;	f;հ����( V��Pm�I-抦���k{{
��d� mkj�P��k��)��#��Fn�T���j�Ү��K�$�9h�D{s�Ϣ����(�$�-&����?��u1�dl��y��Ǿ�T*uZѢ�K`QG�"(�~ �����&��4�tˢ�n�Q���薣��f�N]v@�Vx�!�{0�N{�X�;Tz/k+�$���%��
�j������X�8Eʘ����]K��̌�]�8��ϧ����k��,|�5��I&���b�25n�Ѱ@�,Kg��F�M.<r=��؇��>�L��bf̽WC�$&�v�4<ϑ�J�6�h��t���HteH�
��9��@�vL�c@�.h�}�1�*�^E�G�;5���߉1Y,���[m�7U�����^�v��� .`�U���m�����BL��HRmzCYg��9*<YPU���ؗJ'��F���ӓ+�v����AZ�u� 'A�JL��j�q���\�b�-�5���2�a�,9�9�Y�l����߫��i���gz,��m���]u��΋Ƀ��ѡ��\��_���}^U-3�/7��ѵw�^X��7�jg���tIԫڰ�j�-��J����}���w
��y�{�ef˙��X&�:�����q�RW�捏���o�+�۷u��v��6)�� KBN*�E)�lUX�pv��K/蘛D�Y�)D�J*�q�֛�hv�J�R�Eet���6⬌��mUC�`��j�Mm��]Ub�k�TۡZ4�ڭ�Y�
Q������Z,�Z+)'dlV��+U��bq��:|��U񹥏b�Z�{��C������a��:�JIb�[�,YÚ��P��M��"�h�E�n�U"�
�A1<��8O���i���4D��o���A��JIH�7a���:۵Qȁ�W�n~v�,�K��TB���Ŝ9}%��oz�zrp�{��4%���%)YlrgŶ��k�޻�븵�.�;� *Vur֡�ww&⒤�«!af�\�>?5�L��l��Hb��3*V�!�;���L��>}||��Sw�@�K緍s�i�8�Q�PtƎ����6aO��p��P�a��L��I�jJ#��$A��&�m�)�p!��/�F8xϺ�G�0!�k�1��q�*�m���ָ���<v�@
p��5_�y��X7���	�;g��Fz�'��{P�eq�;˹���A�I�$��������
��]K'����mP��5�p1�.Xc�dU�f<�Q��4W�w���Ry���}�Q�������y�?���r垀��n��t�Z��ۺ+�,��P%���˹��AK�8E��u�ƍ�ӊ+�10GS�U�1<zX�a��O���"1��s���d��m��\��5�r��U�"%��y�C�f�.|
І����g���{P�N��M&J���ǟ/
�ݗS�eN>`��nh�>Q ئ�/��]BY�{���~{��C�pv���T��X�����LߕzD�d��"�'��p�8GR���W�O!�{=�.�y�T���xփ@�E�Re�Ror����>�r���0���%�����x͝�M}1��"�$�I��ogE����F�9l�d �T=T��m�j��UT  �i*�vi��U�q�V0 ��]�˽��S=�ǵ�����|�uW�t�n�k97yIw6u3o�P  �۲�*e���6�� eUP .�P� � w   o��~~ ;��wS���-������:�f��+��
�]v۲�۲ٵ����@e
�J��I$$����dH|��:���m;����C+#G��̗
��7�x�/��>��_1����|�����P���	��5V&!~�-L�4�J��m\��J��`���5nt��}Z����td蒤̐�I	2�n�,1���~�Bψ�_Ij�Ob_�TN���\�*����Z>�µg���B�m�e4nP�zl���d�٤|�.P9�C~J���hr�폺�sa��z2�ބ8 ��;�I (RI)�ÆȄx�?��e���A:�x8�0�ި�u}F4:��l�Ξ���o�����l�V��Gl��7�]��w��Unܻ�� 
m�[�֥g\�*�t�_ȋ�uoZ��8�?�O)Tp�����դ�5�&�����iCO�y2�dR֣$�-ZX�O��k^̙�����w{���7����7�(܈*Fn���l�����[�c����Gr��#4��ȼ����C�z�4YưW�n����M����m$��X�KJ����Zt]�-yּ�_�7��qfd���>6k�]nw��$W����l��D4H&�xѓ}��Ct���a}�XoGѢ�Ɏ�6x��Rf�cŦk1I-/oM%������┱�m��B�c[~�Tܹ���6\���"���c���h=��=�^�/�Q ��W��m��7w^u�u	n�wEwR� "�)��2*� �#��wSo��^Ac�0��=)���I{ O�o>��4���ӒLm��6O�jI$�h��m�j�[5�9k���P��C��G�L�fx��㎽�d8ly��
a2PM�����.�6p�/Bn!w������ARf�#N�4����8:��H�M �M�Y��WB�h��{�f¿��N�U�<p�Ȕ�x��Y]g��Q�lQ�к�E�l����y �)4�6�\�3�Z���|��Z<!�`��WI-�[
�I",=�� ��pn�z��׻+n����ܐ�
�J]�rJ�"%�am&�5�3	��vz�2ݞ�knP�F�������rz���E��i�ШT6�����bᗳ����c�Y�W�,:Kf0g>��g��}�ծw��)I �MdVp��2-XXxᆻ��������ß�\.��]S*��t�&��R�B��x����|]],���x���,4�J��EpB!3��-b,p��/�!K�v��l��4oW�דCl��������CYƥ0x1\;�v�|u7PV?S�]|n%*��S��~����@�v�`[D�F�)���|:�����u�+mw/�~?M��YթT�,۞pRO҂S~f�K1�4������|;��mT~3/�:7
�*W!�X�f:��7������g8 ȶB�[$Vk�k�º��u	b��A'4�V3әp1\*�����i�NM����y$���ȶ2A�B�/5_^�������ؼ�=A��F���EX��Nb��F�8ֲ��9(c��Ƿ��n9��
�	U��[��ʺt�������e|+���};��F��C6�ObIGC!��L2��>��p|o�X*�j�~�u��D�ӱ�H�^FE�u��X��@=�ֽ����g��m��I�J�;����-nsU��J�zU<��2�;���U  *�z��ۘ����[[[�*�[�ָ�ۮg[�k�:��z�:�qZ��7S!Z��1D�q����{sj6Ъ
����il���]����qͰ@� *TU���6��`���a��*����6wm��@�5T�},���z�A�Osk6�<�[��U����U )�I$vISAd�H�s�m���f|�YF�t���j��@�c��u
cח&��{�W{ھou�D+v�kE6>�̳��qz�`��D�l�#�K����"�S��>�sMr����2SI��M_O1�̹u0ס���/�p*႑���8n�r��=�U�׈򷶞�C�n�m�SX(G�F@�1�G�u���`G��$A�Ⱦ�����z��_<w<�����MN4[BP�AYMy���q�����*/y3����+ַ�^���6��;�t�U�A�Z�i$E�V���4�y�wsN�[�w  ��J�H"
��Z4I-�^u�тĐ��f
�ŗϞ)#�ozY�b��=A��x �l��l�Y�ᣆY�N�����O��� �	H��Ѫ�Q��q�8)c��0�0(�]V���m���u�l@ю�񺂘�<t����75`#����Ki�h����������ՏaL×bK,D����!)qo�lY&��50����Hm��d�E\�#��Ե��E�ݰ(r��W�h�Y�WVy3ƋHm����4�.�"�:CW��&m�vF�)%��B���O�H�>�shw���UM�!��r?����c�L��M�����Ƿ|���H�-�;��Em����u>\�wwM��m� �Wsj��r�V�e���e\�*����
��b������j�֎=^���c��`�u��Lxv�$��'�M�Ы��ZG�����)�f>�-1�20宒'L]�!��s�'C��Ɛq�@��Gd�2�5ֶ�l���������tTp]w~�^ʜ��^�.�M�X�.h��a���0�D}$� �(�p�5�_� �	A���>���� {M��l-�Z!іi�w'���{�֫�G���)Al��U�:p����8�d���O�C>R��3�����;�վB<1�䭓k��n{v�l޲n���{-��Ő`��U��G%��~����w׷��,�V���i���b��(���q�\F5�f���xּ�Zz���R�$m���V)��'��O���D���1M5���lÃ�|���'���A�}���X+d�Z1K^�=��6�Z�V�"�-[�]Ɔ',B�*rkY��C��V6�`�ح80#�D�t�m�(�j�L��9������q����X��A{�8�g�p��~�P���O�D:�MP��9��>�����(�@ֿ��^�Di2PF����>fL�{�Oǣ���r��_U���Y�?����_�����n�*���sf�gt,�@�V�R�Sm֊[�l���3ʺ޾�}C���9���=�tW�?��o�k�=Ϲ�,�u���.���Yl(��c���ٜ�����x�{ٹO��������9�엓�]~AX�`G���`�Zl�����=�f����b���jiY�5Z� �3�!FΖD��z"y�"l�P���I	]C��6�g/�BzHW"8>�d�b��b�(ݡ���]��N�%sQM�ݕ2��m$D��B�j>Nd��o�iK�}k�/�u�G�E~�+�߀����ne�n�0��N�W[�������9^�o�����7�g���y� �SK{E�M�<��]��{����Q��G��6�3_e�n-���U����8�	�r�m��m�СTB��*GT
��� �A���ڨ
�P ꪠAT��� j���nX >-�UY�R�Ϊ�-�Te*�� /8sw@;�*����b�� *T*� ;�ø [ �Y�TN@+(<TZ�]][{��  *��T*��  6�  T  6�T    B� �@�� ��2^����6�@P�@U[M���v�g�������]z�v[�*��l�����mݎ�;�T��/�ln�4���U l �E��*��s��T�� ����wk�ۓ{�}ݴ����� ����BK�������~~�軷p�\��һ���׽��k��;���K[VZTD���6��`#o��#�5T�K-l,���r�1�W�hҴD E����B���q�/Pym���� ;�T*��[�U<�wl�h�7�yJ�� �T �   T��ml���@  ,k�U � VJ��YJ�`*�]%��6���     �  �    ~x~�:�    p   T    
�q � Q� 
�:�U
�   UNZ� U
��VQT�    w    �
� U U@  �� �         l �  �P  �Tkv���ꪪ   jܨ *��� ���ȏZ�z�*     ��R����  wn6��   -�צ��lU_�P�U� U]ޮ�&���^���`��n��� *�TU뺕7��n��p�n�ٴ�۬�/=�ݣ� $*+i�46�PlQ�;�;���7u�V��wu�ff]�P �mQYm���;��l�T� 
��  *��P�l
��UT�ͶFٳ��9l�  1J���T<�w}]z����ӕ�=���»�T�Y[j�j�nrU��j���Eؤ�%���I�e_@U�Z�_om�cG�l�>"�e�[m�-�4��.5��eXv���Q�@��zǺ˳��yY�d�n�����+{W2X�:D��`��\p��Σ�^ �b��S�ñq�\�g�v��蘻��c�1�p{�*CJ�!5pS��yr�I���+�H����0� �g�ŧ��}��ۛ�^w��]zs���Ñ��t���:�S�<Y��g���V*�5����ԫH�4�o��Iԋ�.���%]^�kd�S�����vӷ�ݵ�U���.l��dr��V�ۀmQqc����׵�5�h��Bx�f(p��9���X��7�Ϳ]*{��F�["v�n֘�c+D*T��z0V�p���ub���������~ݬ�
Z�%rK`Њ�D�Z�XT��Q�Ԋ�R��-N�j�LwP$j��í���\��j�8��ʳsMp�$���)5�0I���,���V0��p��YS��/��������&���@RZ��*��.����>"pc,9�^G�|k���#O�wCM="ȉu��m#����S�mY
Ke�C�W�~��p�7�X���f�u�lq�\�1�ݿ���+��ǖ$��m��m��{v������b��GwU.܀�-��W7�l��̂�.�m��t�V3��D�5sM`�D�v⣙��x�N'عB+�:��n\�v/5w�>I!�ncMu����7�9���o���vwg�
s����S���k+ �ت�4������wP��xR�Z�uތf�{�_gd6��W��Q��w>���k���8rRe�l"@���M~���ٵεe�
�Ǒ�:B�~���W8ׇ�8LWP~��W�oby��ȋ��򒲬+
ҳe=9�i�Iy�E��k�e���F��A��>��s랛OqW�����TL4Jm����)w9��<��om���v��p��`�۫[�2�X���e|�E�G�\cW��������5�sx�q�����?.5�</̑D��m��n���4ws:�0��B�|���X|l��d��/�%�Z�ލ�0`���,0�tE��6�_D1��}Э}^�(��6�uum���љ� m�%�����ʼ�a�M2�5�D��zfｘ��o�w�R�h�_s}�o�׾�E�H4[d��A�N�)��*Om����t���"�̞�ٜ�h��-��m��$7�{<ݮ���z���Y�й�� ���a��y�n��+O�l�!�´�#u����|_�o�g���:�}7�Z�>A�<�9�B;@�n���~��9��ĳ}bD8��'���n�	��of_s]������_�ZX$�$Rm�72�˕�씔��2���◶A�r�o@	�8�T�(\��z�?nr'�?4���r�Y��ܷ}���qZ�*4����&��S�II4C�����CR�2E��*囲������a��P��k<��[�7�:]����)FUWR�ڬob�T�l;��uJ���p �  ��X���ͻ�qb����  �T��75��ڽ�]k��׻q�e�X�Wm仧[Nn��TU�qR�c�h�l� �*������  *�w   m� �+����*R��R�r����;��{����p
���N��x�ױT�v���V�R�w��v�R�B�kR�o=�-�e���Ӝ�u-j�˺5�y^Y󾈿dN��XeSH�Q�[�#�,�a��Ad�߶xA.Mrb�ӊ{�H�$��M�hQ-v܏9T~2dlq�S{��y��3q������/��k�G�����U�X֞���`*L����ũ|0p�f��9WV�w
	0�X�?�F��u�lX���m�+"���K̃������CS�<�j��I��"��*fo�h���w[�H����@��m�P�QV6�Dg��"�[K��R��Uc2Ww�LUV�1��.rq�	q��j3~���i�N�bh��P���$�������k�k9���M��m�h��r�:^HkX7�Ja���u��O=TWZ��x|�'��W�q%��du�Z��F��_��7�^�o���A�1Ӕ���3C$��=�ͮN[�k�ދ��V�R�JZm|͆<��Q��1��v�9^��hv�����p9LW�sC��MfL(��A6�h*W�r�;�z�M��u<ɩ��p�k���*"�f��_�J����W-��OM��!$.��%b�;h9Jkk9~��9ơӚ9{`����P�B�ճ���bxrp�1V��^Y�J�ݍm�*�^î��y��޵m�Őx  %��I���XW$���o�a�C+$�ĉ���a���C��������AV����讧�_���I�$��-E:��b~F���,9�Br��_�E��/A2��D0�]r��Ԇ��py��wRRJ�A�4z"|r��A�l��	�y%D_~]y@�X�QDh����c�g��l>��I9��	g�C��i��D;k)�;������bjͷŞy��CZ<7OzZ.�0��aNe�{�P�����,�D4=k�m�ܐ���f@�h]��A�ͷW��ryT�,���\���\�{��-I����M�m��ۻ:X��{w���۶�v�mb����1��[�R7(«m�%��u幢.y{�}���\�����qx�{<�������}؟�k��d��%2ܧ�����\�˞�{��z5��W��sa�:��j#w~֞\�L˚0]���ڑV���8Y�{���{*-J �d��(2�%4�
�J��M�ݯ�3E7D��ޮP�p�!�ю�)���<_>�|l��u4��~if��30�rt��͎�>D�J���5aU��a��7ܮ<��G���=Cm�4!�G3)�,�O��JW'm���;��?����������hka�^{�Ӿ�s{{3���Wu+(
��m�W��{J��2�p��]�3+�ٍb�v#]_����#!���zt�gQb�Ʀޢh[�趗���3A�r���3��c�s�Q]Dpph�JWL��֋�b�݃6s�*�G.(��!��M����4eʹ��fy\p�P�hW��h�8�̧�b�Ƈ淜��d)%��A��n���*�&��С�<$�����U�{��#�`ؑ����jY�Y�:��:�j�(�I��*L�2��p#4�e����q�ܲuu�!f�n�SY�š|8f��8j�ӟ���RJ�W����5U*P�*�M�f�c[����5Sof���n쪶�n�wP�UT 
��`1�zyR��;�DT�n�U����<ޛ+=ڜ�kt��󫻦:�ݹ�v�[��<mA�UK� `�S��;��UT � [%e*�p ��m��+���~�q\o^ۚ뵐 J�]�T�AU��^�}��ݺ�V�s^��VAsU ����_E\�w=+�#M?�S�j%��b!��!�8��Y������\�o��	�ss�o�om���
0r��ǏI�<*\���K������k��;pX���Z��_C�*fwv1ã�uTt	��/5^=rk�k$�ƹ���qqi�+��GUp�D,߬J��禎ߚ���a��J:�ZXА�x{Ez���
����+�xs�9ND1�t���'���_���-}��k5����Ă�$�I��1�"��18E�0���J�B�����e��_�Nƻ$�4`�^��|�����{Nn��owMv�ok���$ m����7[U�J%l�<U��!���t'�qx�Xs�ÞF}����k��u]��iU��>.���`�RD*�u!��N�U�;�y=�׻}���)c<�%���-���_us��KG�#�O��$�`&{r���عt�\�qInyܣ֟wrʛ���,sH�Q.�m�����sr��ۧ�e�%�A��Nc�ӎbs�y �:��ΡYE�E��e&�R��U�BM����KW�}��䮎_�\�k6)X;���{u �-�i:m*�Rc�\��&P�keH�zm˙�1�l֎���ܓ�uٺ]1x?�����B������V��ֵ:��;����wU�˹�ٷ�m��f��d�y/�|C#1Y��������ȃ�c��ڄPKV��K���ysjt�͆80�!���@��K��\ތїOG�e����,���Y��9�g����ŭYG-�(Xǥt�r�:UV�!҄�NR�&=F1UnK�Q�W��gt�w8f�;8f5��,r�|��Ֆ�/f#�%g�n{�X�iViC�f��Q�����o:E�&�~+Z��V{����\��*��*w��=��s)߮��6�h�i4Y!���Ζ�-�ꂩT�q-�	�H4�q�m����V�m��8JA��%���'�޾�y����o:��X{��a�d?2�D�U��qQ�� �oV�v�^�|�{M�<�tH�������$t��SPChn�mҚ���Q.kR�0����b�"�������qjqɞ��NC�-Wb8Y �Cm������d�ވT�a��P���]ALb&�8�/Nr���c��ݕV$����<E5����I��+)m�J�׹�nz*�e��C�{/�3pP)��s�Ʋ��M����Vq���t���M���i�{mO3^{�C�����d1�UER�Wmd%ne�е]c�Q�X�r/zpE*�W�
�P�r��j��c�53w�V>nnE��I�:�U��H�)���\��V�f�����$#�-C;)�|0V+es��Ә�9׵,{s����ay�q�fa*�zm��/������ףZ����'l�o�x��:q�Mk`HI�'e��XT����g����@�x�M�������7V�[D+93�Cn�þ���M�h����a:ҹ�{�qG@�icr��rz��?�d�g�3�C�-���4c<BԞ����f+l:FN.�*����׷�{u�W��v�wE{� j�d�l����8V�i-�)�=�.�����\�$f��l~!w7�+�sz;�S[�~�������<$ lp�ȇ�q������*8@��\<Oq||�\w$��X���D�l��@�;]��rq�1{;��7��;Nw��������+�|=��s΢˜��o�8�N���UaBФ�ן8kf��:��4W�V����5{�a�b��~Ⴛ\�]{����#���cl���8ng#����Z�Mc�iSR̖��{
��w,I�b����|#�o����!��'^�>b��\�_~��~������,��*Yקv�6��
R��UC]G�@�wqR�U   *���ԫt��\�wm�o\�^�G�mKC���(5Xꕹ�kZ��v�n엞�\�ww[���U@�R�:յ����l�@*�* �l�  �� �� � �*��m��mvڕm�� �{*�i���XV��U��f�^�Ϸ=��mo`�� )��lڵ�s\	
AR�.�~ǽ�޶ύ.d�̊�j7P!�h���V5�X?xvX2+�ЕN����k����B�cu�&�轕f��γL�(��.�M��>���*I1+{���w�(�h�RFz�RYl���_l���х�O��$�O��o����^׽w�2l^�.�8l�tZm��u�t�f��T=�����s�[��V��g���|�{�`�\.��O��i��	��5vx�y�`Q�TS�]G"�_�!}upe��>ma�<�ݱ׼j��S�:��`mݻ��ٺu��nw=�]�w�w�Vۗ2�� ��R��::�p�B�FZ�,��Ƈ}�w8�cO����5oܩa����ԝ�������n� �i4�	B�i��d�íi'�u�[���v׼��=o3�:d����i����l�7%l~���}�n���9���byz�ևI&賈0N;3R�F�I4
f��X5�FC�~ܵ�B�zR�U1�dV�j]�,�B�A-W{����΃~�I~���M�l&��n���n�F�'��B��J��8,�!о�׃����8*�0�&3{�#�c����w�ݎ 6&�u�4��Z��~,���G����Ұ�}n�f�X�S��67���d��~l��]� m��p�qN��k9w
܊ 6�*U��c H 6�Q�$�uJ���⏼����#Ǯ�8C��ǲQ��,)ũ�v�4��4�iR�$�A	��Hp[�b�Ȋ��Y�YYb �dp�>��W�5�&�:mu��&�H�c��@��k�oK���;шE�f ��j�	S#���i5�P�~�Q��\Y���Zo�ڸן^�92q�\�IS���M9�ܢBtT��+ޮ��B*x���_�=�W�aq��]���$�8��H�sRv�"�Km��R�h���L�8F��R�c���8D����9�
b�:z�8`��B�դ��f۬��wvi��ut�w��;�M����JU BB���d
&���n��ƆK�i�1�̇��r�/\����3M]o��1���U�����E6�����Ϸ��ll�#_�b�r���ސ���]��;3l�uW�_�D��%QO"��|�6�wN�ZpzM�83�{�u�oo&9���`���=�r����B�TVw��˘e�gm��������1���/T�?��^߷����t�I��H:CU�KQ4��Qt*\p��Rׇ���M������I2�$�D��m�Iּr潯f��v�w̫��ݒ� �f��[�-�n��QiF��}[/��3!J2������4�;�o�/�ڛ����i��i-���<��{�5��9�P=�3�Mw�sY�qs;٨Q�Q�ڮά���ᆠ,���:���;C��c���ߐv'�{vp�Nb��wR�Q�;d��R�]c������,#n����Sf���+���@�
qjXgICo�uN�<E���T	�Bm%L��B��Ɩ�]HPz`����Y|O��
����Xp1P`�o��\��.��p���;w5��	�=�ܗ]����;��VU�U�6�gqM�A�uhw���guU    U�[��G��wn�U�T��Y�n�Y�w�޲��;��l6;�k�n��Kn�WMz����T  m��)6�����`�UU`�U AT�  l ��*T �m?�_��+����V۸^����W�$���ۇs��kwnѪ�v�-�@��T��Z�;���lRm&��)�<�ə_]1³Mt�H�PJt�J"6�eDԛj��Ʈ��Y$�RUu��$n�wDhy���T�j����v��j���jw��P�O*	6(W��)��WO�4;�C�8E���ZmH�GQ�u�l�PƯ�Z��D#8�\C6Hdv[u��O�9� ~�uUO��1|�3W������0��n4xZ��_N�ׅX�n����Y)2ՠZ���=���]��~�\�T��i��<�^r����Od�#>������@���[m��څ��]��[�|�Ү�@U6�P���ݱN�Gmt��i4[�*
t�s�Z���k���.І�n�j�p�qb����c�j.j?]9��K]�Q��y�<Ց����׷����+���yA�M$Ym�EdPq��L��$���%��
��xU�l�*
b���L#܅��ga7�C�a�#�I�d�m؆��,=u���`��d�P!��u�˲�
�X7�<��*�¼N��$8r���T���Z~����E>�
�t� �g�o.i��k�kj��\24g��)��ߕNȓ��#'�j0u�z@PN�I��A����ʐ��T����j�]�����ۓӧ!�����3IQ-�m��K����]�㫾��7{ҭysC� T��[X�PѪ��{�玽�_CwX֑��/����!��6q�3��C�/=��9\���S)��B�@t��˧D0�X���u8aGP�ÍC"��11��X�.�<D�~ 4Km��d�/rC�tX�u�(d������8���#��s�Z%o�G��?D=���MO�z�x��C��0x��t�Vs0ݠH-
���\2��e8���\��+�W5ݛ�)vMg!$!)�R���7�l�I��S���e�s�Sِ�!MA-o�q���ug��-t�A�ZM�m��9�ۺ��O]�N^޷m�-�@U��P n[wU�2��Д�n�Y�m���Y��U��|81r7P!!�f)�M1V4R�Y�d���_2�'P��bp�Q�C��Dە.������	=]�)W�\P0��(o�7��C��fe���F�lXM�wP!!��/؟)�׽P�=�9f����`����=M{<'q4�+d�B����Jn��5��[c<�*�](ר�H�>!w@�\�Ƹ�g$�j���"	�.���?����I�hb�x_{R�iEҦ�h6�7�<3JŃ���%k�.(�S����N�U��9�mQiQm����Z�xkw�u�gue��K(U*l,��	--eaTv�ѐ�k~�||G��F!R�ԇ��p_@���w*vxr7�Y�_M������LJHu�i��a��F4:C�����.�1�
�<��%SpЃ�̞��r\�{1��@�K%2��<C-��O܇�7;���f��Z����#�弭�H@#��m��Δ�0�_��2�=����5R��G�~�Xܾ0�#ǨT���!��[邏d�����P[t����S�R�<B\�R(�Í���:�^��<˖x�����߸��B��� ��'��`�O���$�� Y $0�ß�  P�L�$ � TI$�$$�����4@��d�$��Be������!BR�Bu��<?��~]�����{��s�u�S���Џ�~3��_����xB�~������@ ��2?������������������B����?����������������~�CHE	"H�A��I#$���B#	!!?����K����O��@� $����������6O�~��=�HB�3Y�����>��ߜ�7�~!���_�����! �������=��� �B�|��؄! �S�,?1��@6	��0�vT��������\Zw�l�����O���~ ����.F�X~�?�؟�~���d�B@?�������?��x~���߳�ا����u�����������I�Z�:<?��GA ��S�S�v������������@���$ !?o�?���p�p� ��~�����������)��d�R�0��0(���1 |x�@%R*��A!U��d�� D�$�J
���JR$QT

ITBEH)"B!R�T�I@I*�T�������H!E* UJ��@DTU%�*
� P�$��
�� ��A*��J�J��JEHI@��"�(B oU}���{�h/�ϥ	�O���z��U����W�����޾�K�Ej{���D�|��҇{�w����{Vԓ��Ψ��D���{cL��n�
e9�ʪ�>�t��;�ֶky�UE
SYO>�$�QQII !/}wo�7֧c}�9�ƾ쩽�9+ﳭd�ﻀ����(���^Z�ڭ���W��1W{�}�����F+��f��}﯉��������O3Bo�y=vS-6��q�%(�yΟm�RE�D��J6o6P�ڽϏ�S�J�^�,�������t{ ���S�SF���n����j�i�3��{���T�л����I�;�Ƶ�\��ډ�e�y����a�tooJ��S��eER���J�-��
<�R"� 	�_>n�^��i�k^v�Y�T
��4��l�}��ﳭ2��Ȕ��5/{�K��f��Eը;���>D����N��2�J�9z8/>JS�}��y�)�Av���R������Kl[+ٕ/]w�s��"Z��;��w5��z�#�Gz������V��T�yU��JN��gR��}�U_}[C�ϜU��o|*�}���"��}������Ʃ)��_}�"�*��S��M��m[��J_}駛���2�5P�Zһ��$�� (J�R�-��z������.�N�ْ�۩�N]v�f>>����ﵭw�����Z��}�u�Jd}�3�uUm"��m�X��ua���ϯ��5;h[}���<)4ʾ�w����eI�ۣ����ET�Ѣ�P�ﳾ��7ǟP��=���2ѱg��H��f|�x��]J|��y��Z��iGS��|�f�O�CӮ�R��O'�6�%=�R��$�ǧ�x��R}K������G�I	R���>�*�@PR�R�����2�/{�ƶ�Z������CO#��>(��O{����R=�s�}e]�y�޺� ���g�]����i��|H<�o���Z��r*�����x�e��m9�Um��UJiy��۴W���ԪW�׷����uW����f�_;�c�Vۮ��=��Ӿ�{"E�P+t�����s���:Q�Q;���}6Ͷ����z:����d�}�
�{�{��֫m�>��� �}"�J�ET����a{[MZ�c��i��}���O-{z�#��R�|���^��J/z��z^v�.������+q=�������:U]���"��^q� E?LT� S�F$�)   5O��5R� �D�*�4d��F#CO�	�UD  =�M2)#@h'����~%~#+�������S�����^�/�������������$�wwY��'I$���N�$��wO�:I$����:I$����t�I;��'I$�������?�����~���1��6ڞ#�۞��4S���g��8���<�?e�V�s���6$0�Q�I�a���v�n��V���L�5�6-)$�0�R�%۰���v����L�����~>���/��JWGʺJ������Ƣ��;Ic"���tI�B�tl�0mfc��
���t��5h���=º�#������jEvݼ�6,�AA����"΅j�D�o=8����΂�.81������qge����+t�朘�rz�aʍ>���In�x<���G�cp��p������X�
�d�ɐ��;��/$.��8��;�7�S0)� �����(��S85���;����9��%���ݾ�ahgH�Z�-eؙ9�O�h���a)RB���ʉ�0��S�Mu�M�0�nˉbq�6Y��`=s .�Z�����	y�
F򘗍�D��`�V�ŎР챷Zt���c���V��{�7(1v�KAk��F9޹2�,��,.��r�����F�=�!��pШtz�j����邃�t����{)��;��iܑ��71�'?Qq���G�䇖�І����T6%Ч��;�;!�b	&���!;ި�5��@F�8	�lz7B[��N�d�J�n�Q~�͌���J�2�Z6���^A�M2�2��=ޟy-b��a�/\�}�0Z�^7BƔm	�6S���Թ����YtB�z�t�`�h��l����Ab�UX�n�K�7�7Gs��M]�v��G��g��e@^�Q��iV��Va�\�l]*�e!��LWMv���螻�Z
qF�VձlF�Rm����9��w��F	�iS���M�x�woNM�gd��c����II�[� ��x�ԧ�Rrh4�ܠe0�L(	W�`QD�&�h�M��b����5����m%vrf���tĔ�a�a�b�I���3�����7�QB�bK"_�U�Ӕ2ɧ���I�	nq+W˳�4)������3�Z�w{f���f���Q�m�{�{NQ��5��u�;�E;�;N�+��K"��3WIͼ��.fr��]�KW������H$��f2��0�6��k��<�TDX1&1f)'Wb�{��0�C8*ɘ�^��ɔ�ӎ1�7o\K>D����^���G�x,�+L�����;��� j{��COX4�ݢ��f��q�q��(ߺrye��V�S9�6���%݊JC�V�,����/���=&z�R��V�OA);��%�fHnڤiFm�PbW�u���zX4Ǜ'nK��p�2J.�r�>.V0�R�خCd'%]�0734��%oT9|8L�t�MW��WA��D��JM�n�'��/Aש����3/"�$lǴH.���x������6/x�_v��;Yb����Q�w�]� ��%a���+�[iZ����� 7WӖ�w�|r5/����cM"9�����q
7�щu8���<������q�%f#��@�[6���n�P�nL��,��Ϙ)�d��cSqj)��ub��3l��n�N�0A��'*]ad٠��;Flūi����Vj�!�:{�*����^�r���!ۇ.��n��_\#f��ˈ=7�M�������Y0�Y��!&��ä�����pe8���@�)6�qf���Ň���RP�����8<@�I�i[q���ֲ淤:�=�\M�~��ư��C	u���CN���Wu�L܅U�Y�_^�]����(N-��+&��J��xc��V�o'$ׯ$��6��q��Z�M��h��V�[Ah,s�i�Μ�y��T*��r�L�L��]fnv��Z+U��,׈k�U&);#f]�~@�Q4Y�8��+�L���=��h.QT֛�[�e���
�q��8����Yl�X4�LXj�ܓ&�����,����t�ma{rJ�Y�h�ʍc�.�G�E�6��Ga:��2�s�d�}���v6�C�N���r}�^��R˭�hS������`�oRFTw@Q��b4�x�X�
��&ڷ�!��轛���D�&�n��^̝��a���6�^&z:�
��8�!�N���^�]\.��fȉ�2���O�f�KO�<Rplk��{�b�����s7S^n�7}I��)���"�y~�V�6T�rz��yS��A�Z7��<ѓ�/z�cX��);^��3l����Z�24Ld��Yu���-\?�����6�Lz�@�S�Li��K6I���G���J�88������e V�=�4ڻ3we�d�q��7fo[6i5^9N��pJu�)���)3m�ݧ	�*����5l0*�e8�	1l0n,עݙB��n^f��*���3�Sl��i��x��-�1�n�^�^5��[�{[��Hiw0�b�6��ɨhbG��R��u�;be�.J�x.6������U�N0�Y#�{Yp�1��l��%cuu��5���8�B��/�398�Nx`�8�O9��}�52��5�M��Sܬ��������0�(ش<!ޖ拿`�6�j�AB%�[{���)�F`$�"��,X�u�� 6�5on�gk�ǻ��y����CnZ�=�7c��7��1����c�藎�8�}�f�؎�=�jMJ��2b;b�/-DY3�̰�6�FG��ٹ�{7j���]��b4>�~�4c��`��NN|���pb�w*�O��	�x�ʻc��v�l�-����u;��*��I
��t�:��)g�#��^������ڴ��t���P���8U�0%_r��%����jɹlb��ѧ����tхˇ�3��;��q��lC5̘�cg3,ݬ��T�C.i�'���6߰6�����^\�ۺV�Ce�E���_�-.
�y�hTi����\L�j�
{ٽ�l����41��m���q���:WÈ!ny��a8v&�J�X�8�\����Go.����YV �CRv[��{t,uKG%�	�Ƹ�5?.�N��\�5���`��B^��=�ޓ�#i�{q�'2�BT@m&����j��48��=d����㳚-��k��N�r^��[a�s��-��b1]�z9R����FYvdYQ�A���<'*eܒl9�n�5���*7���Ǌ[���7����)����(���Tڎp�^h�p[V��G���s�No{�Q�2L�74��BR��$5%\���\��.�@���e��A�|)튢E[+��'kc���k N����-�9 N��0�P�jr�Ǧ��o����
~<V���E�{�WG��)����QЯN��k�Y9�z���=3��^9�#�'������4f�:ܣ?mZ6^*�2<(e�����p�GJG�ru�P�X0!������)���g#��n���J�I�7���s�ak���I�7�!]�^E�L`�����QŷY!���ich�����.Z�%v�ޗw��"=�_ۘ�Y���ݻ'TU�x��uC�%W�1�&�����Y�i�̧Q5�)Kg�.�ȍ;�r�.#���У9���8^Z��%z����[ǣy̖�٘����ӆ>�3b��(���4=�ӱ�X�n�%Q�3v�l��wQȣw~+grE�e�Grbhǵd󚶎PNR���V^�3M�#ժ���M�Ɏz<�SN���w��v왇#�Ϡ� C�H�ڨ�~�����J�POc��N;�D����we�Z:m+lK��Mh�ׅ,CG3X���b4+�D�ދ:��n9t��6�I��۟>0���:���a�CX�n��� ����FP���8�Sb��l�����M�޺&�M	(�z;\ѹN��;�OT�f��WWnq���A���Xz�E�-ָ��^���ḙP�Y�Y�_NŊrx�v�s���qN�H�ݔ�g8�3#p�W�9��A�RLk9�;tZ.�cXάԠ6=�Cc�|.ƌ��"v���s��>/�HP[E���w[�^�.���Y��8���בN.��]�+O1��{6���^�;V@ޝ���*r)�M�{�v=ݺ�r�8����d\�G^aDnZ��ܠ�d�3{�!��#���)ـ%˹�B�=3(��ً6�q��K���UL�7�
�2#��5�x���kF5���S��5��:�d��A��\#.yG�'��۽r�xf�9��;�x V4peCg15��{��K�"������u{�Ss�'����[�������,�Ѯ�8�l�:�C��l.� wŀ���}�G��!��{��P7��O`9Dz���M�<Ls٦��jxu���4���[�ɖ����s<e���y��!��rۭ�r�5+S�K��js(��p%M&SM�̭�o*�tN+49�wl��y�n*�9V^�4��h�N:P3j�u�9D�R�2�a��Z#��!+,.�ʺY�]&������t���R$?wM�3�!�M���Qʲ��)ƹ��l��7�9s�^Ԣ�R��9>s�c�<�jW��CI6$!Q	�z���E���?����ø�vf��K�֜�#nڲ�fƜ���<��g�٢��tX�x����3������uv+��Ny>Y��(ē*p�!EʎP�Z���k�d����]n�P�zh.fā0f|n����t%� �(]��"�P����=�(���-l���p=g�l��{�A˒��x6#"~kn�~5�L���x������˚��[�i�d�c���0�,��z�㴡����Iߩ��j/Ya73��@�#HK�4���99�x�������֎q�OT!�"��5us�cͼ�j�����.��Mг�L��Fӓ%�d'M�!����7���uR�XJ�K�[���Ɉ3��Xy:Y�9'1\���1rܿ=X��Mm._eR�r��D�FT�y���͉�2\X4� JM%I�V��o
��Qu eo4tX����	����tx{�E��i�΢7�ɖ�:��Ѳ\d��R�۠�����\S	���:�*�!���x����t�1�ݝ�z�V�}dk��`�2cƕ��.�[k��G3����f�Qf3(E<�����]�XP;�吅4EoV�%����i���	�ٛ��}��^3w$&�<�!6B)��4M��B�j��ғA$A�n��T�^��(R�h�F(@B��(���s��e0t媼Sh�`mh*�:6��L ޻�@c5mm+���v����E��k����v}�����i��̅��/̐i��Fo#p��Ýэ���Ε\��?����_=���P+�5��GtlӶQ[Gt��^7�.�)
�w�;�8F\qΝ�p��o=BI���H�S��oF��oB�mUʟ���%T�gC-� /n0��죵�.�%�JwT�̡������ӕ���d�D���m� ��d7 �*��̈́]ߡ�q�W��6`��(IW.a��qb��Xo&N�jx�-rlx�|l�y�d�R�GF^��WkV&k��g�U���1oW_��k
؎���SŨ)�ML��.�m����2�m7�%;��+��Mu<�P��Ua��Fm��	�AFE8��o��JWK����k�
E���&7������㓗p��!�Na�F��T�����HF�3w79�?;�T�u,Z��w���>O�CfCH�s�p<j����)LV`�����&xcZ|=��������,���=�=��F&q�m�G6y�Vsק��y?31�0�ݬ�b������@1H��6\��i����5��݊��żsX+A'/j����Or]7OP����J��އ9�����@7V�%.�L��m[Mk�r�A2i.k���u�4�z�Teͪ��p���.d�-��=_#�p_��/(�l�i\�X��Y»H�~;;�8���T����d���vo�q�Ē��rs��ѝ��A�����мwȞ��m�X��i�K�LJ>�B�m�N�����1�dxA<����	�U�*�V޶�����Qx֣��a]��<-+ѶAGs����Mȩ㝤E�᫃��ۇ��W�b�9^��b`�k���+'<�p9/SG#w���\2����u=`LQvF
���47�*��+A�m�\ݼ��,��",��"wm��a岲�G��D3f���4+y��=��tu�N����wG^���`�`�hU��&�Vo?;��[
ֈ����1���K8�����H�w�F+ұ�|��a;��V�S.8���y�hH�3�Jě�lT,��.2��n��l�dA�{N`��ާ�U�.F����6��jZ��Vn;�3`�u+���.�%�5N�s��fQ��˱kC�3�ya2�R���r[=9�f�&�eӗwi�U��ʹ2��l(cw��(�O1,�����M��e	��81��l�K�f�����s4N�n�N[��i�!x�Z+s`�hu�CPgo�b�ne�x2W�JPs�b�ћ9gAɽ��S���I�xkD93�yR��Iv�qfj� �m۰N{�^8&� �YuY7�����\�I���@�ɚE�fV�F��9��)�V��0(�lM���=4�c3�RӼ��A�7��wQ'ob�(��.y"���ݓU�rd���о4q�-{d �"���"s��ݣ���~�<iw��[���X�C�'1N݆;Atܷ�0���B�m�06��i`����d��{��5�AJEtsqd��W��$����g^]\̛彍ZHzvo�"�>�@�<��n�G�1��L,ȡX��a��"�%4 6�'aq�P ]�pS�E�*��WH�[r���M ��f֢ۛ�|�&� @��&vWa��
R�}�.cR[,��s��+UW)#T[*���UR�X�I@��V,� ٣p�q�(r�s �s��������9����t��;G))��(�����0k�I�4��G]B�e�&*��q�.�WT�G|�[T9�m�xÍ�tHM6��b��b���N����Ծ<�y�-�!b��e�(�`4�]�VWm����P��WhÙ�4vuyWLq�E;b���N�4f��i�둓΃��kã���.�Di�ם��k=��Vgru�2r�@m��9�v�Vl)��v�v=���^� �B�E��J��H��:�m	�j��,pV���� AƖ�1��a^��v4j��:b�Ā�Mk�;�]�Vx��cke�.��VX%-���U���!h��h�R�:Qz,���@Ť�h�Ѳ����h�v��*��
��T�u�=���m�Ѕ��cPc�1Dw2�e,ƕá�v	e�R�ͯ	V5�K�a΍�����}x��x�����s�iK1.}ാǪpn1�l�1�m%�1C���^ �7��,�<�`lfDK+�x�*�F�00��<�犻MB�v�]��򯶹|�=�c�e�&���pO^`��8;�Y��'m�'�.l�;���a�����l�1ƺNՎ�Snd�!V�1ǣ7�]M�T����`т�����ŕN��s�^<jX��v�]�m�,��n�%�&�R+IaK��c&�����ug�Cxc�ƞ&�J���1���Zf�`�f���)��[a��\'g�.}�9�+I'��Ek4�����:P囋�ъ�GWa�[SMH�-���m�-�F�-͇�:�s,��w�k��yM�����ت-���r�נ[�!�6V�7sQ�J	tkh�����B�]�-2^yG)Pz�+�����^�M�@�\WB��筧��#�v�+\�K+1��ۖ"bmt�fH�
v�6�2�1W���)�PƷc�1���c���j1/:z��ưm�ϪQ�!Փ�xq>}����[���=ry�mb;9Ez�Y(wl��մ`�q������W�m���p�^��&� ����3n�k ���If��y��n�����Kh�X��c^G�\�G.�v�@�i͚0��X�kK�����ّ	��j�)�!m��#s�պFw+Wn��d��J����kFl�c�X��114�ƂYCu�9�,�8Jxǋz덳��Vq�7\6��7�1�f�/n�+��`�@�Yq]���� �2��&к�yE�s��v#��["�[��]����1p�Лf(��=�����O'c����=Y�#�[1-��-2�-pK��*��+�\f��0�9`y���*�c�Ǜ=�s�싰x�i4�gyW	y���V�
������ю��z,k�p[t��8��'=Jd���C�	C��9���y�Ǚ9݌=��s�+��é�ט������ڨ�:�H�1i5�%�hGgjДB���ؼU%��=���C��m��0R��b�a�Z\������ݶ�d�
3&�00ۦl��&ЫB�X*J���Xu�n<LZs�C���NŝU�����2��/,��w]�����\@�c���J6�_T�Fvv�����Q���]���G1Ă.�ًj��%�	\�/A�M� n�;v[��c.W�wE�'id!�%Mwf�o�)��v�̏
q�r��ѹѣ���9�%��{l���oɻE�p��Ӈb�\�%��ý��F�|�o`�x�eok�q���1'�v(��	C;����D%�ne�;6�X� �@��QP�p����sB:^_c\l���#q��\�E�s��a,&	v��.���U�����k#TD�bø�q������N��lݰ&r��.2��)wC���n[���v��{� wu�b�ܜ��p����XC�ɷ��u��=%�N�*v7eҮ�v'�EюKZ�3g���Iv ��3�(s���B�9.v|�X��"<���'Bu�6Tll�8G��jl��a�Y/<�] d�t�{���]�S�	��G(��5$-�n;hݺ�^�@�y�C��#�n+��m:�ѻ!a�Uk�l���+&�fՔsh�����2�zǄ�kd�x�%�p2�m�;���6-ێ��9�g����i�3�����*��r�շn���9�y�s��l���Ŭ�xE�;B�'�ź����i��:�(v������l7�fp8�GD�YM,5a�7K���9��r\�Z��nN=�U�^��g�^6�(�#�,Ƹ�vHеkC�����T�]��ǲ�Ḓ�T3E	��2q,��p� �]�x��5
Vav�:B�1���WM�.��&�JN�n�[�s�g�l�;>{i�����8M�x�&xpݦ��6F�&�� ����GQ��Ep h��vG��jp�"=�w\z���nS��.6s˩n	:p:��n2�6N�v��0���1l�:�������;u����7�a�sk��mi�8�p�v�6#e�ft�=u8<������"��	[Whef��̘X*X��%�2/(\%��FWg�K���kA	c6+�	n�yW��kr1<t9���v�Y���7EsV�хY�*bR�����l.���d�IpX�b-�/R�K��M�b��Q�V����+���|tt�7�)I��<vt���Y1����n�b�,�a��Y�w�.�mY�Y����ɍk���vn{	��q �i���ʦ�����xu�xmm�	��C��6n�N���),�s�	��I��:�0e)�<d;Ύxp��h�8�7�r�s.�X�!ݵ,�.�2�.ئZM���:65 �cg��ɰ�g��C��5Ѱ����p��+n���,R�d(	B8�M�]-����ˊ%���¸�i��ԡ�u��볂��V&�k��&�x�F�e[
P�NA��
���0�m��8�6m�(��P�9�4���vʀ�Qò]�t�cq��죞��M8A�6痶9]����0cn�3&��f���=8'!�{U�(���2�lN�b2�5��L(�̻B��n��&�f���Ae�k�LL�kl�����ݮf�j��l�H鬳T��2�rb7�S;�$u�Q����^����kL�)P�YM��Q��d�����v�g�ባ71�=�׈��.����7[��O!��v� N/V�x7
�c	CWY���e,�n2(Z���/=�1�{t��L-�Z�X�&X�p�Y��u�q��C(�����<�c�����r(l��rXzq618�
���s����bUWP���.k�v&��j�Zh��<v���&��p�GAj���b̝�"m˟N<=�.���k($�X���2������U��v#v�m�H��f&����*�CR��nx��[�e,����I��\���]���/ғAX�m`������╭�5`͞�v Ch6&(Kqe�8\%z��I�:�N�q����l�w	�&z��r��6S n�^�^����k,D҆��w=�N�קN�2�뇓���,�%5!aAtJ4*8��m�M��V�n6�V�`Cc����g�D.���v0���x"��6��+X��=�BIƴ��g���r����pql/;�e"��8ք�	��iR;�6C����ͩ兏n��ʆ� 2�x�=i�s'9�w`Z5��W��˽��1��M�q��O���4�qg�.ݮ8�������yݎ���mF�#�)t�s.�Y^yf�e]�-I`�X��X�yƫ�����=�֏e�ˑ�MJ$�����f���.@u#aej�.&��k�㋊���f�`^ێ9�셹�U�U��(k�i��x�6�]����#��
�:ݜq� d,�P��3#��at�x{��q�6��]�o@R��nx'`!��|��`�Arl��F�'):��4��nחq� �׀�)�5�W<����䁭�
���8^g�]��q��H!�u�������Nx{(���1E�3-��d5�f�=	J��V�+����4������g/�E5i'+����z�"u���ι� ;љ�:�q.7vk�ƒ����]g�ܕl��V��a���VY��JRWK`e��k,��K��2��ٹ����䞣����{�F5X^���ל��\��
��fe�)ct��f}d�7gq͔�����e������tug��p�d�F�9K�/[a'=g��8a٭ɗ���7=s�a{m��K�p,�&��:r>����	q�b��Iϳ �.G2��n�e������W`�XSR��ӻ\z��$0m�z1�+�p�k�kn�]�C���6<���[J/+�(��:.��Ƨ
�kbl�[ 	ɻ���#��6rC�g��et�]Q���X&T���㬮4.fjG�h�	\-�䚶-�u����v;&�z�����;��x�2Yu�!sg/\k�=�>EN-ς*Ճd�]Jck3�!K`\�:�-�h��J��+&ۊF���GuԱMn�]	�<� �˹]����mBu�B�W��l�WF6�&�ْ<9|]����-{O&<9y�ú�8k�\�q��!�ĻK�q�F� ��2�GR�hn̙�ta٧�v�%�8��s�ݺ�&r��I��qaY]H�,��/(En�GNM������AŔ���������g�9�{bp�Μ܆�gȕ����!�y�]���aU�
)����Ŕ�Xb�Mʰ�	m����HeKАv�Y���KZK6�Ƥ��*ضM��HB�`)]4�&�s�.��d�r�	���H6��d�����6ŗk1i�Y�iB�
]O��t�N��?��N���'Oû���pN�$��߄��wN��t�I;��<�;�N�2I;�t���I��w�����;�N��	�;�t��N�t�'w@��wH'IӤ	�'wt��N��$��I��wN�DO������S���(��'���n[��Nv�tN[�Ud�%����u����k�D�y�V�`�kl�O�S����-SOwh������/�"	�q���O+p��B��Ɍs5b������f7q���؋򱆦�{u�u<y��?wz��!�\
*
�>1�D�e�@�[�[;n��h�uFh*&�]D� ��bt��.�\����ڱZ`�d��7�Et|����9�u�Y�$�&ֲ��f��2�h;���L ��Q�H���T362�5�'k"��NVx彿X�4�!
0G� ��'�<k�+Z��0yUS.���,%:�cm\E�+~��5�����Q(;;wx�
�}���?s�`�>�4�"+Wl�0�r��3�,�[4kA�)Bm������1���~�y��ٻT��??+$D���HX�5��ܯ�t0�{.4z�֧KH��h�v�ZT* ����J�X�yF���eH�k������8�i�6*���p�O�6�Dxb��8Pڃ��SN��q�^��Z7X�˩U�$�����6��
7hN�b�h ��2�.f��'�j��F٥���m�!�J�d
̗h�x���f���~�8V�\���QC���ۦ/Ә��m��i0��؍y�y��ڶ�R|�["r��T1H�`��-C������[/� Y����1��xNM��OOWX��J���mfҒ�� �M�6�E�=�5�[��\��N������7�k&�Є�	l�n���]I�%�x�,��c����u�g"�����Øc֓�vی�[.y0���wT��n��wb�1�Ա'7g�]a�H�8�v59�&�
ʐд�e��4�lE!k.�:�?9,�/���u����ƌ����e�l(4�bS���;yCo���}��! E����5�@Cc�t��喀�N�P����E��ٴؘ�f���d�{����d��f�l����m׌)z�>����;B��%#��4�����%��g���F��t/1O��߯	|�ނYeZKl7`�#^9v���^�]�����1�ᒛI2�d��ik����њLc���S��	5�37}��B�W�;b/LU��>�eb���6�h�EE;��	�N\nK�Wsú��{��99t����8_n?{.s'r398��w�p8-�j��v�z�`����W.}�(Ƽ1:L�&\4H�aZI���,�Щ��_^�~������쟙܀�?#�\צ�f��+f���U+eӺ�v�eV־��7��<7Ew�GkلaGJL�H���]ȢUףէ,�WJ��j-��xkvZرҞ8/v�z�к5����z��6��s0�s4�ccV�Il8p�p��V��v��)��S�8� �z�犰��~go/k���F�f�6�U��^��F��-�'��T���[ᘬ��k[;w%��u��l��c3�[�nں�ӳ1��(��f�0�%}����}a;���2A�;r��5��76z��N�a�ߙ��P����6�f\��q14�ld�Wj��$� � y@)I �Wm�d��h,��H�<�h򂜔n�V5�O������H�U?�ޣ 8����� ~tq�
��C)�X,l��Q��Qspl�pI��W�E�8�h�n���n,s'%���[�� �W����ɉ�(�, ���zgUI��z�h�$@�������=^.f{�6���j%py����5f�*ŦZH�f�����,ڑA�e�L��<oa�P�h�b��Ŏ�\1{��"2ɴn�wz��<�:���ˑ�`F^�J<�f*7w� �$��+���Oqx6�׻7��zίo��͓�g��g���L��������:.7����U�ʗg/�=~IC��;�u-�y>�6�	p�h+X��;��:&v}t��w��
�^�����a�O/g ��QJ��_�Mu+��_�����[r��c0j��B��[�Nㆈ	=�7U�9�X�|�m�ՠ�q������YC�m�p,͎0*j���m�&����g��ra�h��! aI&
M_�����P��+ql��_��!R�띳��i�<�k	�%��e����Ke)n����c�=�w����b���Km"�,0X��oT�޸��XXذw�vW��x#j��w�	�h2�P��雺c�R0��a��i��n��f{([�����ݩw�{j�Ly�DK\Pq���7�,��#+�wN�}Z"K)��. */�z��h��vj�1O�5z�����d;������g�4��{)N�}<�r2a��*z͍���UH6�ȣ�B��~�XZ��K&�6-�G}�}���֪q�y\.���+}3=���I��S�)�������x��34z��m#�[1��b��������� :��)0D
5L\\�8�ʷ�Je�����u���.&���9.�����s0�3U���h�j�?m�S�W�N>�ut@��9�r�9w�`�`����j�Z�쑕��ى�
2c3j����@n�"��!$�^�����R�ġ�]��k�`%�B���m��1c��H2�[��5	&��C���Y�Z<�C�\&�w��V/�{Lj�W�\0�a��5�s4S0�f�ض 4��^��b��iQ�fnY�
�>���v�^7���=�׈�]w:�E�ڭD���y[��{�IBp�-0c� ����[�Ff/��r𥫹N�p�+'i�p���л�$;N�73���<��T�d�W�^���\��d�חf�m�Ҏ��kWM���SO��l��p�|�7{��I��c��K�c�����ԏhg.Ŵ)hk�Y�}=9:���ŵ���(	�ل�H��X/a��'Ea{�go,�>�Q��#�n����[�)�/k���[�y�+�\�N�l�1�s��3�s)]>����!���E��{)��1>�f����4{��M��|�lM>�l��w(�W�u��~�~��L�6�مgznDc)�l��i��a������v��虣n.3}�^MznL	�@x����F7��-���	ѹ8;�W�M۲�q�����L�:1-#vsgl�Qtu����G�i�{�ɭ�0����wf�mfO�'�1�S��lKL���!$IB����+*��׭v{�r��(��}{~�c3b�G4ǽc��>���� ^J�#E��/z�/p>��i���_�)�����w�Rឆ��D�v�~�}����{�j�W'oc�o�_Y���J�ۀ��8�.�ț[�,�^s��/Jd��$��S�ݚ6v�����I��=��S'���`��f�EY6e�#.Z�VC�}{4o���B�����\���,���΋��{�*6+n�e��/�g����᳐2LT��@E�M��.��۳F]��Ti�́�h l���v�ַVR��5��D��1�U�V���ݶ�[n�gK��E��^y"�od[c n̙���[J+�q�����h�U4̹1���1юv��ohi�Bj�hCк;��kt��z��!����z�vI�P�֧۶]I���z��\�fK9
�'N�[����~?o}����x���ˍt�����ʒ�<�o�����)�A6���׍ T�u���n�{�-I6t�t����oo^������Ʋ�
��f�����]佫��4V�����)���^5���' ��'�݁
"�=��rM	��Z�}޾|ѷ�iI2�L][�`�`�g[����r�e듓-�pˆ0aA)� �5�no��9Q�<�׶��u�����)�ٻ������ҘY+v�\�gs�X��I���36����D����A;� �5�͜Yq����#8	2�å�Է(K����`{f��a�E�����\�l���p��"�E�h�%T#VV]D�����rIy�+Y�y�Q#@-�l�z9�]�f�2�s�/��J�T�6I�u�����26���-h�L�BЍu��4����P]`����2|5���J��/k��,,j��	/=a��� �f��,B)�ءu�Q��4ˀل[)p3��"�B�Lgr�f}�6\��G���I3�o�Ok_�5���:.�D��L��/�B�y������O-���yp×��,�c0,��������۞���F?r�Z5���?,A����n��A��6�}���2��-%s�V��o����n%�[��k���̊��H� 0`��i�:0������L�k��[f����j
��I��_���ʽ�;E+��5v{�?y�*[�o�^�qO�lg�q�t&q��r�{����@1��
��V��������Ѿ�c|�W�<�<��$4O��P��z�(�|���cެ{;*f���)���ͩ�y{ײ�����~$����Zg ��K�́��^]��j�I����xZ��ש�����{�n����g�����c��fB_�dڽ�Jz��s#C.4�p��^h��*��j�w)/:r�Yq5[����3��y��`��=�1�ޓiV�Lu)~�j8�w^9��I�F I��q���F\3�n�X���F�a����l^����O�G�7�]�T��V?m=�����-y��3\��I v�pzq�(+p����p�D��A@�E�E����&��{bLR��j&zI�pM/�a%�l���������G'��� T����xL
����]��=���=x��gL�Km��o=��ŢLj��`���/H�lTy�Z2���+#�8�6ֱ���K����
�����}1����w���VUcf�B��ku�o�^]a� ����k�8e`I�e �dfz�Y9�m��y^�����x���8�4���,�~O�v(�J���ڍ�bok<�nF8����326�S7� t\CO뀥hݵqn�#�V��D��s���9�֙Qa�v��\��������J������{v����En,^���w+�I'	m �m���D`Nn�e�q���U3'�Tnx��]�F����+�6V���\צ��i�.�<w���%�@E���������<�mmlƉ�{'[�`�~wB)K�聂�ޏey�!<}�gV���;����,��z���퓹�4���"��	f'j��wޞ�ٵ{��Pu��� k:yނ"|	6������q�r�7�vZ�s�:?�m�S;���箦b�X�ʣ�SWu?�r����4q��8��Myɣ���b%7�I8p�Z��ص��n�Ww�/~��$�V���|g����RZ��`xR���M��ݫ��W�n�l��i����`�	������V��y������?m�.���e�:"��Y.�j�zu����Z �Y����C�VOS3�����J�ϨFxѬU�.��1Y��z8Vƌ[��Ý��۱�>¢�Cem��o[�G�ò����;pT�}����Ф��哥�o�tp�
ln̈́��^\Z�Mα�7����]n�i��r|�wy�w����΃Y�7��޲b�&��������pj㽇V\8E&\5%+�oVgVhJ+=�U�����ZR�ܒ��F؊��}/e[W{��\�Mڳ����a��H����`���iB�NƈsE]�[�1��SOF��?�$����X�[��s���-�W�໐�����˟'F��тX��H�[���~ߙ�^wU9�Wm�;��3[�V{�v��A�ф�^냝�Q3n��������1�[�w7MA�)�2WԼ�tƭ�<��ģ�nDIy3F��]!�ó��G�6*$3�i��uyhi)�\A` �4�6�h����X��R�;i��;N�^ό�Oa�9Q��W�T���d,ѻ�3T��}�R�g^a�ߪ)�cG7�mG GM�A�Bi�ج�*܇�Q���o�>M���g��J�/q]`�4��������i�%cw�.ݽY:7N��NȿK8N^��v{��Yx¬�����r4u��.L�4���F��W�!��kk�4�^Vm�q�2�7=�u�FSC�H:mŭ��0��WCm��K�n��[Oc�n4e�k�mE�B,���oϜ�O,��$4�':ж7�i6]�5�Z���ݥ�2�闋�f@��3f�K�iƁ����4v�ts����A��0f��웫%����<��Tiz��h�4R;rv5��n-%�#qԎ9	L������8�0��k���eܿl5^�[�@%��1�@����i>�J���y�K�~WW:�W�U�j��Ւwwt@�j�d:w��h'�C;q��4�Ƽ��y��4�#٤�����{w�ɻ�k��0{��P+^�tU/FA �$L%���SO��s����V�}��)k.Kd8���܈+��|���_e�`���C	U�%�n*N�;���נ�&���
�����oxP�z�>�`Y̱�a��ڝW�<#s��=}Ȣo!�W��F������[�^�:i�I�F0���=*��?�q��>�"�I�tڽ�;�-C,�!�z��:25�sY/�d2�-�*��w��Jd�[�w��9�R��+�6�ϧMηچEa�#$D���S6/5�aˇ�����Y^�Z�SOL��e�|�n��i�D��?OE�޿W?�q����k�ܔ�G-쫕c@�5�݈S��f���dÓF�����(�{n��b@�B��ߦ���>���8�{s"���%���D�]V����Pj���3v�-��3Ѳ����z{�=7QF{W��Qj��}o����ԅ>���.!�:�-vQAR�t��x?0p7��\�o�7C�8~�T��܆���X�p٥s��S+�zBa���j@�ֺ��6f�y{t��.O�9I#H}̜�G��Ƅ�W�Ԕ�
9�9+�`��=�i�|ݫ�W�����}�}�zn����ge,�أ#�,���2WXf��5w��%�h��O-Bk���A�:Z��ȠȨ�ε9���ݶsS���?m{�=���Ė�����
���7;���9Y���䍛�gL`!B���+^��b����g���qDEv�;��&oyn�_+@%*��K-r�)ȹ�a̜�����5�c��wUЃ�����]=1j҈{\�ܣ�+�A(�u�l4�v^�-�]%���+y|���n���`<u6;��m��U�Y�c����k\��1�Ep^��2{v3�X�2G�|�����d�3@�qt&YtL�ynGL�t/�^�ʺ��Z��3�x�{բ�:I�#\�x)�3����®���I���}�q��d
��V,�G'��_��4k�q|����~�>B�ʜ��)lay�IyR`Y��l������H��b�Oo��M��Ӱ_7���3pbp�T�X���t�`^�ͽ��D�}��ci��.��2.����D̻�lͻ�$�Bq��wrI�潲�x&��C��#=Ӈ���vz�Ny�ѓ3_7�J��m��0�+ q�ή��]��RLʮ���LlMnc���܉��M�V�u�KfݖK<��9�(a��%�-S[R^�َ<v���>�P�B�cF�liH[h�,�*�k�l"�fƆ�Y�<1cI�X���,���dh�Ng��^g�Ö�ӹ�"����ap]�!�W��U�k6.MZf܄�v"�n�\G9�tR��C�;���&��)է:HXq�� ��B]�m�`����ϋk�{n��*pX蒸��\�'�8K;�}sT����r1{pd����ٽ����+�Vޒ�e��aܜO6 ۝;��x�f��9�<
�3@��('\���c����[�=Gc����^�l��qw8��L���[)Nj��76��j��K�{X9yQ��d����h퇂�6h&֑���J�y�[�u�v���jM�M5i^��E�������i����I��,I�9��Օ�E�CK+�k��ӎ
k�z;1�3;)s^F���Nn1�3fư`A�K��B�+t� �ڤ3z�tB�*Glf�,7h�K��[���ׁ����s�7b̠�fW�v;VfSXU��[eƶ�����ilu�������hS�=Sc9^��`Oi����vx�Ԃ��L�ӈ�b[mZ��d����'v�<6Fm͗����h�1��<��:�mz1�;��f���+)��m�iA�(K�k�3#(�#�2ֆ�V���ݳ7�����J%�<<� �#��95=����Ora�I&��m�(x�!8�c�R@|����fwklܘKQu�����
��<�6x�b;F׷� <p=���hI��wj.�]���'gxE{`m����[��ݼ��±��;sd8�ֻ{��Hr/@�w/1�+7.�+bn�u�bX4��ĻR�F�m�4�-u���73d��k��]T��,vÈ�@����ͅe���v��D�z�n�P ���D/t )s�U��5�6 -����~@#�*Z�fd�yk�V��-ۙP7>�@��P�	1j�w* ;W�|����5�FX�+���`i h��ͬ2N��V�]��=�KP��ɫ
�{P�eH�y�,�V=�b�K0LN��S����;��/�uC��::_y�xM�O���@6���k
�9�.}�M���$r�ѹ�`gP|�Ite���������x<Ss�l�xk�L�&w����&X��� �����AӁc�\`����PG�6Q�7��P��!���w9w׻k�շd;`��O���׺Vh���䕪|)l����/P1�z��fSP 8�U�%'��*�fu�,>�dU0ވ���3�b��z��9����g��=^�J��O�.���P�����n���1e��Ż�,�Vn�JH���-W:0�N�~׫U�U�����$�,cS6�]H���������;�z��9Gu=��}�t��J6Ɵk۫��< d-�@�\UΞ��{�̚NS�����xl�-i"o��m���{��e��18��cn44�fƚ�1��G�='o3E�b�y��6�g�+d }�4��a-a����9(����U�缦�nјohm��nw:n���8�﹇�f�ӗJ
���޹7E]q����q�9r���Jho3�@xeVI��O��n�Q:�
u�ނ��.��g#�������ɗ+�/�T;�P��G{��ot��H'3��� �+W�,��M+;�z1��O�x'�;�����/�]8/��D�6��;7�[��w=��ٮ��,B�*�,N�F>�ۣ[� ݂bd*ð�#^m^���X}���n�:WM�� �į�[����#�����8p���{׷�}�D��	��W$�Y#�!�M�l�[�R������Fĩ�T��ӗ��އ��L]=�,x=[�ulg�!������K�[̽��ς�E<�wỠCA��hD��=e+���p����~��1�@���mE���6�SJ�����fQ����Ok�������R��n{72}1���,���3r33nGj�E�
�W=@M�J�4���,{f�U�Y�H��s]���z���q�`q��̦k�ӛ��H��U��fm��2:���l�@�F)�y�Cz�uE����O�g0�5sK$��s}�v��#�Q�Kp,�]I��M�T"Rl(X��ӵ^=���՝�2r���
*j둌�����*��ā�ױ}.ٛ"�c�MxƚO1��J*�לi�'�S���*}�~�n�5gu�FZY�3ƪ���ոo&Tr��̬�H]t��Gs^�މ���ȷsV�D�l]���q�'hΐ�o�sէ�ZM�e���q�3臨�� sgu��'�_m�o)l���ߊ��{���v��߷��Iw��X�@Ʃd�U��r��R��­ �H����;��8#Р& /���Y����Y�
+s1Lj22�Qs���t�������ónh�1��&�up{��!������39x��#�X�m�k'}�j��l�EL8lR�n���>������$�"�ɖ�'���ȝim���t9�e�\�1�㧒�؀��,�n�r@�
��(u�o��婄8��F��ٚ��b}�H]MT֚x��ɚ�� �{Ėʪ���^ʖ�x �p�6���x�C9�3��W>� ��<֓��Z�#���9\q
%�bw_�}�yr�)S�Y#��@�����eIq�ιKE�]�M�(���l"�I�i���M�ڝU;W7���@�ߥ��?y��T\gL�b�Mx���]�ԁ�^��`t��L�WGT��.��}�;F���"1
U�>�� ~p�p��##�&�;��gP9ۯ�grl�2ɱ�߾5�Ztj|�k�\;R���_~�jv��y;�������
��x:��X���q���ѧ]�a�v��|�t���Ñ+�)��r��O<��v�;��ۀ���1HGd0��6�CXj��Q����y3��є�	�4�ꓴ^�����P�l��sH��i��K����ۥ���.p��y����D1`{�v	�����bs�rf����(G��NC��d�N�E
�h���q�2fk�L9�k��f�y	[f1���a��l�c�H�\k���3X�m?O/��@}��� ���/��(J���w*+���va���n�/wO��H��I��S��0�<j��:���RK�H*iƴ#���qՉ�Nȫ��3;�3&��Z�CZ����m�n#/�ͻ˗O����=WU37#�t`�G+0���;�^�MH�Ӛ���)0оY>\b�h��L�A�$&Ae��c/EcuLO54�)�Q��u��7sɭI>5v��ow���e�y��hB��"�@~'����[s걔�zO ���GEv��Yjj�s�t���&ZN	��W�3o��/K�:�dT%���۔�_{4��9���XZ9����O�t��@^�!k}y΄�?
&z�B]k��o��=S.k#�l�}��̤���6��!{�ec�wQ$����3�jtdP,g{�i%mΓ�X�/�״������O��h��Nmn��R���;J���e��� x x��&����dw�#O��X����n�ٶR��O\ϺXyw&w�u���<c*���)�mu{I���^YRr��s�@�H�"�d�u\Ӷ#G�s%��N�C=����F�W끌���Tĺ.����1cU]=����������O�V.����t��}@��K&�7ܯ�-R����Ƚ�c6����(��w2���|\�gc�+H�uv��/e��*V�ޮ岄�Ű�y߂G����g���g{Hu[��{zj�7(���ͰpI¶2.G��^�3m��E�D�q��WB�O�?����n���'����&G�P�K1[cE��+ʟ��L'�J
���/;�*{��Q���O�}�s�t�ܰb�d?Bɬ�,�Y&��%�c�`�s��wF�x�Id��"��Y���>O�M���Y�E�x�����j?�-B�2�V���Y�#���nuI�޹D�	�:��d��*s��3n�ح~���ւ�u�;�j�'�ʝ���]����r�����^*简���o��`oy�aj��e��)�X�|:��_n]��΋�d����l\�2�g�����A�����8rG���@�X��)���)���"x��Y���{�~ǜ,�<)`Ԟ��|f�m��B�{�$��vk�ˬ�۞��<�<wر�k<�]�L+�8 �)5�
\<��f�^�)Wh��"�����X�⟐#s$iu�����{�ྐ�u�#s�3@a�fMC"��^��F�3�����5�0!+���mo^T(���9�Bi4�)��=Ɵc#�	���t9=�`�%�y�kT�}�=�>��#�Zj�v�e��
���44���4�6��~0J"L(:g�z��7��L�
I}쎶
7����4"7��%Y���p[K*��$ht�$L��7�\Xt��T�^6��݉����{��՟!�%���n����5��Q��s'��҅俋�ӵ[;��U���jm�(��؃(���I���1n�]"�����̓\������rg_E���I���
}�C�[7K�{c���֍��-N`� �6j��	t�=Y2��G �2\6YI�M�rg~e[{�`���2�{��%p�T+����$J�^�ol%z�1��Mfrk������PޝGc���|f���<}&7��b�D�YO���hϊ��L6QB�	���Zz'�xR3���o�x=����R���J＾މ�+�G'�by�3;+�x�<�]��Ȼ��뚷�}�S�'�,�1eO��������j.eM�)�*GZ��0p�7u������b�-����]cp��vq�c%3=֑�R�j�	vP���n�_1����!u<����7�G�M�p��j(�\M�̼���pmN�����u�U�(�JBh�0�<��9.,^���^�<���=�׈��@m��*�ϗ����ryJ��gG��xNV+D#�~�Y{|e�!�ʶg�׽���,�`o_vtЮ��!��L�.]�^�(6��Q�����Ϣ{g+��(�Ksrz�pE����j�[��搷��&8�ݵ���o�)������c�3�s�)��p��^��k��́����p�$q<�W��������oEuLu]0�����&�d�]��WWX�;��v+D��S�飛X����+�ܸ:��|�=p^Å�{�S��qEq{Q}��h�+�}ݢ��>�;s��V��sB�Y��7�X*%�;�ț���?q�4d�ik3�6�e��=��"ӄ���MG�{����9Z+{<��,�+���\��$��:�n�B7�ӡ���3:|�sa1��h�-�	��Ѻk���|��I[b4v��	�J���\�edw���o,��+:�����S��=�/1����M��ޜ��|����$@f&��]���H_U�"i��}���5���G,|��[z�ml�ƽ�P��&I0�g�	._�{���a߾^K�b�Z-1�H?���T�`$O��%)�"�C��CAM3��n[��c�{s��sm,a1��[=}w�K�n���_(l��S�Xj68�s����]��<��l�΁�1?;wYv����@���.m��q=I�=[�K���؇�OY����}��淕�4o���cI����n}�>���.���ľ@JS�F`^������}[�w�E�-�y5��>;�.{��]VLg�mf�7�����K�ty�&N�X_XP�Mz�7���9;=xeF�q��Y�~ށ��W�$V^_D��χ���X�آ��P28�_��%�E[C��h�������%]�b��<g�.~��f�8�7զ�~�<���G���T8S��;�lǛ�U�jĴW#H4q���,�ٍ�'4��SvE�3� bD����jC0Xl��Ĵ����M-IA9��	5��Kx�Y��PX��E��{�Q��.R�0�6#RQ�F�+l�SYt��XGn�8������ϫsY��W���fH�N�`v�͎ݬ�6�Z0H�MC$pi^��:����lzm�.�rQ/R��s�+�7���tm<;�z��'m�v\�G�(�8��1��!���h(MEa���$��W6��ߌ�8�Xv����uo�w9S<�m~�̵�1O ZP�\�~굺���ߣ6��k^���I���b�	9K��W�^�|��T��5��#r��,����g�z)c��f��J�s�2`��=��ˊ;�З4��i���$���嘖�)u��t�|����5}�3G��z���P1�(���؀T?�Y�S�6�zۣ7����  �fEA$�pS/ݻ��ȩ��5�W�R��9��0G�	�X2�{=l;JY�qUQà�V�u+�j7��ͦ�p -Y��'���uoi���7D�u�U���ޞ��a�KFn��=��\@��x�5'"�gs������R��%�~3��U=������8I�`9��2/����"4�g=��}�G\|s7g���m��}�c���G��0�n6�·i��#���;<���qG��CB�&��F�{Ѣk@'땻��'��hZ p\$["��~�9@ʛ����j�-���-����w�\UvF^-X�(���Z�j��5���<��6�Z�׹�,��y�wZ�W�{��R���)|ҹ��}6{�aʎ������f%���N����k=]��df�V3,��>�Y�O���bj��;ĺmW�`�5���~�][Ȟ�;v�w
�I�^�6�W��}��B6cq�7C����:���|�t���Ϻ/x�f�NAk�U�ѹF�e__b��o�~`�k�d<${`���3(�\�K�Ы�����	7Ij��x� �p�?7X�p�&�6B�kj���W�/n�D�4�Ѽ���R\`V�k����N�8����s;���͜�ʓ���O�	ʾq�v��^����b��_p����p��Se�e�=�{�[Î/�ۍI`��}(�綖t+�rã����+�oyOhA�`�W8�P����雜"KZ����y��)�^-x�;��TӞ��}U5�0���+,a�I�!w�c���5�~�(yo.�-N�`p.�%�y��]��e�'��Wj�@��{*�q�k=��&s3�EO��\�Xjl��6�]�Yzv;��,��"�fz�3Ann(�S�ї�Yn)uw[����P6����m�E_��,?K�پ�|�e�W��5�/���Q�-�w��s�$`p��-�3�gh^��uZ6k�������~6��1��Lz1����.����v"�b#w��I��t����r�=�"=Z��u���N��n�y���׺�GKnD�
詼�O$w6�L�g�)�J��B·�I �6��nC�hnܧ�˰��M��m�.�"��=��=f���j՛��䣪^j$'�7�lV]Mr��U�F�VI��~ַ,g9���=s�X��̲�J���e�ۨw_p�r��Zp�O6s��s��W���Mޏ�n�����:���m,#�;��}�n����W�����>/U�������@ѯ�SN�U�8���i$�nf���&m0:��4k{zp�ž�)k2� ��Mv1k�nO��X9��<��t"iT��Ir�|�%��E�νu6���!t4l��
+${`�g0xGK=t%����oƔѝ�؟�܉,���LU�QT}�:��۶���jο@y�;�� ����LT`�"͜�=ĳn);�j�f�\d��M�T
�i�
��R���X�]���	ܦ���A�>�C�$�*H�Q�}pr{�~�;{���'�O�4]_dI���s��{�*�j�;O~�R1̈́dC|�:7�H
���m#9~mu�ι�gqoV3�+�>Q.{/�j@$�����\T�#�ngY���
٥�;6��Tͯ����x��Wu�\�ti��II�K�M[ñLjy��;��I��|Ǉ�O�1m�s�Xa�H��\�
�Vy˗a�����f�G>�G���nwT��9�V8����cu��ޖyt�>��ފʔ�2�R��R��n}8��̿(�V��[�}{}s�*�SԜ��ـ���8��L&�.VE��l�z��k��4���G�z� �Q�p�Vn��R���r���;ۿ��5>�
P
ߎ�9B
޿A���y X�)�a��7�v�������j�B��G*�[�6,�[~��ÁZr�O�D��g2��&gt�ێW��lQ��h�<��y��j�]uqp�q���Â���q<)gx-���{��׬+�lȮ8�7�4��kA�0c8�n�,[w$<�B�\�1o֡�@]�aܛ����{�o����uOf�n���|�P�Q��l[w9�R�������"�To;\o��;;d��%��5aq��b�����0�ڙ��:�?墝�hV��/�}ٵ���4�_I��GMK��v(��J'QR�����'�z̋���d�yW	�]�Xpu�:
��`��X�!h�Vf����A�p�-�Pvu�:�*��a�Je����H������λ_ܡ���V���ȍa`a�y���G7�wn�X��5�DT:u�WEA�w��M9Y[d㩻3�)�']�OO�, ���f��F櫛�1��U_Vw܏k��U���{e���4��y�.3,��0tS@�N,�G��� �gW-��[ܜ�3�ĢJ�)`�5cqBgO{���	��w��[~�������8��n��[��L*��,z8`(@�_<�D�zF-w_u�m����*v�8AΎ��7tJ��uEw�V�ށ�Ӗ�D��Hq͒�z�豮�1�������p)��.�\ŗ��p�OUaڃv��wi�N�g�+�$.�^��cȩ�mf��>~kp�ª�I��ogv/_��|a�o��
]!�)���ܖ��.�z�y���ڐ�r/�	�у�]Bb"����NM�d��<4��r)�SEê��	9�,�w_�oT�]��Ϡ�T�A�'��}Ӟ�A��g.`@D�Idy�s�^���Kr�|��똤���;��P)(�og+�q�d��4�-��=i���2C��d�^lP��������c��n)ezM�^��	���a�zy����N-�(���!�h�59���a�p�lG�-�]!w�ǳ3��A�7[j�5�.y6�֭(�ٲ��)!B�?y!�Tt�)��w@�k~��[���׏�Ÿ%ɭn�Ol��������j68$�6��� �%u$r�Efe��_n�=*%�K0/3�d�>��P��S��Ry����j�=ӳ�\�+��''V��ܗe���X(}�^��1yY
K�� <Z�9Y�廁����P)�h�W՞�Ys�>����ئ����Ɍ#T!{�s�dE\{F��&PM�Leó�фē	Vͻ��M����^g�ڊ�i8���*�E{��ֺ�P��Kv�Oc���ۺ�2Ľ�H������xՈ����')���ZT�����B�>d]Fn������Lm+o�ƭtY���^���/�ޥ�l�F]̌��q4n7���
������]��=���.�N��{�LGQ���]�W㎤3���T�o H\�	Ap�B�_PRsM��`�Y�v���!����r���g3��'22qoJ�[��yt���ޱS^2�X�$�;���j��d/�8b[��c��Bf��v[���v���o�vc\�f�rvڄV���le�~����.�6.�8&qP�̣�a���	\YYCVQ��4��z[Xh�m���ev �C�����Gc���#�9���'<�z�����.�&wil]	cd!b����0R���*�n��6�.�w�L����^fo%v�-͝�@:z��u�����+{V���ġF�s�3�R���LRu��-��W=��x����U<k��u�QK׀ڸ���j
PZ,�����j����xE)��P��*�y�����f��3=�=�nb�"A���[������IA_"<�4r��C�@N<�h>G�ͫ8+ҥ�$�!���4���p���c���^/oE*��g��Y��C��'Y�ee�.{�)��S���՞� ���ځ�J	��bk"�����Ĉ-�� ����� ���e[�������y���5�H�Qy��#o�ˆz�9�ح��X���x5v2�v�E����l���$�=�gv���g.O�G�u��ꋾ߸L"��r��ޘ�p0���@z��~�OX��2q�1Z2c_got/W{c �y�H�up	������c �59M\r]�����36}�$��7,vȫ���^f>�*���>�7DR��t2u������V��3�ȏL쨬��#=#�\ -�H,w�H�����%��Q�پ����.��@�qY`L�몙h5=ؕU��kr_��3C�ݢ:��~!i�t�_��{��jgn�`fJ������̷���j�M(D(�1	�f����E(#Rkd`����x:��)C�3���n�x���{w�v��yWi�5�<�%���ܫu�6����|tR�ev���Z���;2��A&�0���F/���]��#����)e#����9tBC�I}�s�Wh��4��d%����_?k޾˙V�$gz>��6R�լ�K+�&��Rs��s�9��j�^<��M�/coޞ>�^�ݻ���P��°��{ܭc׽��<+�(}^�<�k��t������_��B���\ɐ�h,�V��,����UL��0p�#L�{������@�à��d��1�-�8��ۮ����Ivd�dyNЙڮ톷\;���?;������������'u݆�o�0�J׃�oF���̜��:��0�[�� lf�M�&��r}��u�H��LXf�3R�������+[�H�cJ�+��ki�NF��S�H�P#i�[��VJ�38=���y+�VC�ݴ>�sϞh�V�c��m��;�whg��ފl�'��A��[V�T�/'c�����s�&���1�T�8�d�~0w'=�VD:>�k�'�}�g��3�޹���[-�<痳3�7����oDI�ɸ��K�w0��a|ӂ�
�{]��I�\�}��1x�#I�Ι%���2�8a[�t:�]O'+xB&���GFh���f�N�ӄ�FeAs��ʇ�Q�vH�De�L͛��n����f
 �(w2yD�p�p}=G��Y��gz]Q�]� ���kԾ��j��]�8y�(�p)ؼr���r�W�Th���Η�oz�����~�,��qXw�w�{g��Sγ��`F)8A��'��j�L�vMZ��ܜ�Ic�E�386�}kh������S;V�p�X]l�됍	�gqGe�3���[hi��zw�7g���qS���'�L�6n�|�>��?)��Z��[��5"����a�L�(R��R�<U���N�J����>�@E[+7r��8-�c��}},lͫ��q�}���7J�"��zky��ݾ����(�؄6���s�ũN`]Kb�b9w8v�&���a�y3���޽��u՛�y���+2�ʶsV�U�:�j����g�	�*�N�ǜf�JV�{����8�O3�u騺����%Р�@_+U4@��Rdb��2�M{ˢ:��y!�t�n���i-�N�Y��f��ݻ�:&�w ���4md���˅O�X��\�f��0�eWn	��8����"�.�C��ou{�xg>��H|V��~R�	���+�`��a��=���o~7���Zs��n��g����'͡d�dt&-��ZD�5�+�
����=7�+�	l@h�a���ź�fׅ]́�{��=���7�e�+^G<���Q�
}�$P���|�|pw��p�@��{ӨRz�h�#�����mR���˪M�1�ЌI�s�Q��pEk0�L��q\���ު�2��p5���>���R�[����j4����&]`M	��If������1V�rs��DճY�1	�7n����{�OR�-(���䡟LM��<96Mg�q���>�w�����j��q�O�_	����[-�6�_\��,B��C�'�v&�7ٛ>�1��'1i#W���27�`��=CԶs�P���݊����"!U,2��	�.W,F�Hb;�{s^�U#Џ�L�e��g�+1�S��0:N�Bm��ٍ	u*�W��j��/��`�1���`K{�RS4b��BF�k?����8�R���8�,�sV���F�N�"�!X&oj��.�=y���,�a����&p���ͳ篃���0(Y�����ｫ�|�'1��1g�W���nO?�4��]B�v��Y���|�k�}��"�l7�/.$�kɈ�cy��{��P�+�yy�f����o��⛎���Mx��Ǝ=S�]�s�k�<�F���R�P�r��it*��c<���L����3��t?�B.��
������[y�#�h�
�`���H�#�L�����J��sYz=W��]B�o{�n^P ��q!�M��m�9���M�ye�㤲�>���k��r�������Ml��nm0 \��r�ƈ����)��}'I���'|��'��5��ct�H�MH�8��G1Zg&����f�+[��Yh4؂�?L�������b��g;�_������M���"�-�	�	�47ݞ�"(g��.=�	3�7�9�K�w�?c�TwF�i0�J���7�!����K���U=��Cr�ɛ[�8�9�ySl0dݴ�f�&׀��nO{>��,�j�\k<�s��՟M��xɴq��N]�MB'���$KB	�TZQ��r�^%�K��vpg#\�{	.�Q2e��~x��=^���O�
���'��8@�~V� )���I���ٺքM�g�`/;U��7Ĭ=F���q0�Rl8j+������ݙ�9g=�M�PH�F�z��2y�b��W6u�@���[�����ْ�E7=Csv���k�dѳ��a��ɿ���3��hDv�����XW��"�cY� Ђ�A4ɂ`�Ym�#��=7�uc|�o�r�gS��V˻n{u��㮴&��Ѡ�Ӹ��	;�rE��^9�n��MѵU����]�i�pA���Y���v�g�:��=(�gت0�2����sţ�M��� :���j���g2�*����g�� �Q�,e�m�{e�M��:���;�{l�e�(Q��*�z䓈�]~G�	R�wq��zA\v �6�{U��+�&��ɵ�6j���U�<v�Tv���PE���j ��w�X���x�h��z�I��Y���'5�njTg�<�-�N�dҒ#�z[*O^�[�~���%��)?t�i���`�<������	�at"�^㘜�ќs
Bm��C�#��M����/6��YZ�W-�?d�G)�iz�P` ��6�/��m�t1k�J���v��v��ʅ�HNʎ����XE�R���Ms�VE�l��?���K�:`S_w��f`��f��$zT!o�������κ���`�7��'�9	S�ʛq#��׷2��#AIHn��NL��-�
w���!��5���ޒн���V�s��^۪�U`*e�\�6z�]ŪT����f\W��$��Y0��XԒ�K�>w&ei˜�/W֫��`��x�k7i����c�������N� �{���Q5}�$�ó(
�<s- ���ӛO��8LL��Af��i�\�M�נ��4�j/fD�^�ϔ�����Vj�����Ut�>O����w��&�k���X�-,��o�j�{��߸���uR�Ǔ�#	���$$$�ڴG���w��WK�'w��vK�Y�2{]цO�[���b9a4�ʇ�Um�MF�$Є:�otY���ͷ� ��DH}�ƂʹF-8A��͗�SI!��*�yt�y�(�x�=K���[��+^"�L��QK`��U���x���ʩx;�ݸ����J;�ߦ�c���̺���="�AP�v>����W��|���A����ʠƝ���T	Ncsbit�B.hw�����J]w;�k�lC[�=��YM��ڴ�qk)3m����O�����Ll���D�G	��]��}Q ޸c��	zݜ�ι�=x��uFb��]�󜩕�v���L{~3���$�hM�)�=���$,�'��<���
pDQ:�=���3M-��캑��0g2���V{��6�(����pd�w��A��JčM	��WR����"���C��=5q�o���J��rk�f��Y���}LI�P�Wu|MFO���W̳F���@�2.��!�N��/�5�UQ��z�;W��2j���8��I�٬����Kx����EO��ѻ͔� &YP��2OA����-����ݷ�$����*���`�B{Ӱ7Q	�!ݚ��~�S�1v���L/�{�V���u�H�,��WWL�WfU�+�0≁Ћ_�^W=���Gg��1�9%$��n�+�!��J� J���庖�bZ/4\V3����]]:�ǄNf<��o#�!j�y~� F`D�lbC�q+��w��3g�r$&�a2l�x��&!��ϣ<u�!�-�R[ӥj��Ɵ����OP��W�:T�W��k�l�ܹ�2��C����H3�������~�3�{�j}A��ڐ���bqA�c�dߩ�j@�K�8�W�f�O���?���8��ק|�`T�ഛ.͎��[ �ᬧ��O������{��|m��W�g�ۙfj�����{�{tP�a�Pɂ��B(t#2a2��G�6=�Z�Ψ}�q* R���{��R�#��>��i�=#�`�;���:k���1i���6�-�J��������ۏ!QϷ�B���I}5�D/�{k}��9��y�з�[�
8+�'������U�Ϥ��f��{�����2ۛ�61�e�#���9����}"��F�1�"I�6˼��xG4�	����v��aٮ���J��y��A��xኔ����o,C4�Eh[]�B׶gú?��RO����$��i��kh}��I�*���t"�oUMf�i�Tqm�M����>��\�6,Ǆ�ul����mn���vx������R#	���z�Xj��E�ZͰy�֪��/ �_L��[c��#6f��*;R�w� ��hB,�*�<���u��]�Kѱ��r-�����A&,�n�B���ݛ�g�Őyc���	W�(�{��^^�Z����)��lNu�ۑ���"@PAK��S}����v�f�r���� 	�DT�L���G�a��
�9L��P�&Fm��{{����w�$�%C��j�I3z_�܎Mz!�L�����W-I>��O�P����[�9әF�<�v��ܪ��u\a�#�\���2&�&�JX�l�����ͫ]��tsњ0Si�SD��Hu[=P��uG��v�,��R�7�5���C�}d+zbJ���!�3�l�e�S�b�/E��č���x�aM��+�t�A�kkZM�����+�I͉��ByB$��t��#Q>x�h�!	K���{��a��'u�����=��D�Y]D�ܑe_!�n;&O%G�����v�,C�i"��,&u4k��P���pW�K��wo.��	���������/�ffs�W�q��\�X}������02_�����zueD��Y�j����n��`[�6D�s�ٵd����	FP�� �_A�����g�
5ٗ���D*���ě@u��V����9rV�l��俻�6/+g�ߗ*t����/|�ۻ{nb��7
U8�߷P��1ܽW��r�u�^��"%��`1�z.�P�>���S���=nr���p��;��q�t�OSϼ��)8,����+;�r�m�c�vn7Vl(�w�����r� �߫3�/�+����N��TV�����O�_l�흵؝�Z�\]gr�)�<{�k9�|�4���Py葃*�Ν���;�2�n��=�x+��.}�:���.�/�.�7�3��A?���׳Z��cD���>���Q�%bI������B7R���)Tb����^y.b9;�~]F}�Wo?�<��0�*�.��Ǽ�r�]��������\ݾ��=z̸�mB<LX���J����0�(���L��D�1������,��o�ã�<��j厓�2^��p�w�45�M�����]:ڬ��>�rǇԁ�A�7;����{!�N��x�o�C��Tw���7��~�J���e�2[=����^�	��G���L��6�U��.�C�,Ϯ�������\�S]q<�G�s�9#��ܱ��d���7E�@�Y�U��q��5��Bc\9��K��|�
:S\���d�����s{�ƈs�-�X�h�v#5�,��&���;�u��v�ʀ��=�Í@�����5�$�1�k���2��n\�6^^.��B�k�b�˨�G;j�E���wg��n7WW�%%�]Km7�����Љ�{��������
DA��E)�{7�W��
��K�K�u\��t�F0@��4r��}靗�o~�<��>~��)�?I!��I�F�[�î���}�Ygmg��;��5r�FMF����{��{p ﶲ��H��N/#��٫���z�^���<L4�h��7 W'�&�Xf�2ꝧ'T��1�����9̉�E8`N��s�����"��.����C"��Pc{y�QȖ���,�Ks��n&�i�,�"ƅ�WNs��n���b0�WVu�*�i�3s��${��E���&A��}�����86@Q��D��3q<���M�+��|��ۂ�E!\d���;��B��|EywuR�a��hZ� d!��uقc	��Y�"F�t�F�{ßQf$�D�����Xr�*���ڝͰ�{�V�����3n�K99��c%D�gmJ5N"WVڣ�l8jmi��/g}�N��V7_.H<M/�[������)6�-ʤ��C���i՝�[V!����t�s���P	�c:��g���o��^�g2^���:�\ J�qn��uxN�[��S!k������h���A\�`$�m�.��w�ך%{ͩ��u����f;����Ͻ���0(�Ϯ���'�Hr�񻛅O=~�>$�Kp����=��kǔ�V���wQ��@����V��a�^>Jl^-nF���|gs5��YS��Ջ0lk�y\�͝�|�v�.��hn��w����r<ɑ��D����Y��^�c�o�	�y��Z-ju��<���<�ͷ��z蟧���3��ι��&h;}��pt1�+󃏩�g�g�=��sj��H�:���W�1�)OLw�rWVr��xnK��;�Wcʶ{B���/
k��{w�`��>+9�Y�Q�ne���z6;-���gw����u�-{j�f;�|������:�77ӷ�(�G�'����W�i�꧊t��z^�>7��#1v^a���`fpj�����Vڧ����)��+i
�*���j�K���~U��s���߅k��p�	l�|[�ۮ�D�0�1�d�߰Fȁ3���K�0L�t��2�C�)��6%pfX�˥�<D]�������g)��/�P�g��h�РD�3�Ll,���D�"��韰Gx�Ad���޾s%ƙ�6���L�]�G�y.��)���1��5�v��.�s�o{9��:��[����+��B����S���b�V�P�T����F��=��n�s
���6�H����<b1w<�\�4�U�M�.�;�x�V�$G���Ve�ŏU�j�ݡ"4徠�Wzۖ��E�;�k�Vx���ٴY���mG�5λ=Fe���V��A�m�#�֐(�L �I��7`]g8s6���4̡)�+�51s4P��u�7K�;gS{"9M vqj;p7.t��{t�எ�Φ��4���9n��\q˞�.����o�oaOHh�6N���E�+�:'˸���s�ӻ'�x�z�z۝O.�A7r�%�¶d�����{-�>:k�!�'W[p�YS�n����;0����� ��m�V-)Jc�����:����=t�ܻ�� �n"�j<b�`��e���9 �mA(E�q��"I�(O'd�7e�n�	X[H7YK������"rm��&��n�;lx̒!�j1�;3v�T�K���F=6ز���KC"�ԑNl�i)�(#8kt��r*ۗv�]
v�v��б�B��B�[�Ym��$V��H!��m�6U����l<H�q=�l���Q�n�E�Zt���6��G>W����;��狑�ӡ���=.����=�l� ��/j�m.�&C��.�#���0t��kfv����k��p/�9���H��:�n���λtr���c����2.��!�n�M����8��Η�;���5��;9�f.�'7Y�S���&"5mm�7�M�����	����G�N(�3Y�Q�sz�	�r�IX������eݢS��l`�g���vbqF%��(��3+tPn֬�u`ChS`nn.�����
)��7(�خ�\�ne���N�y��l=��`6JM��-ўg�|�c��$���S�I����Z3YT#n��u�n��nd�������<v�<q�4���V�i����e�]!e�Y2�@ƍ ���s�Z�l��07%��u��v.Xk��^e�[L1�6��	+�p�Ὄ]�gZL��a�4�F���<Ų��i`���Ʃ�7:����fs1\�jM�C
�Z���
�c۝��r��Q��$����a�u3�1�[�G�����Y 8ͫb��(�ښ� ��a� Z�0���P�n���w�� ���f��5b����f�O�;Qj��i0�\�D��ZCx�9�h��c5(`�õ���i���,3 �����-�!�uW1V�J*rt��8��-Ν��"$߭�omu��L�[�K�:�;�N�Ajֲ�*3�s�t��)�u�|�R�+�s��Ӿ�����`n�_�hA����֪_z�7)�$Lt�ƨr�:�p��ȕ;O߈�u��u�,�>�[�ٳ78�wP"=�!(�/L��glĊ�3�	(G@�&8��t�5q���(�rՓ�{��t�To�!�+�M��޺�������PZ�Wv{-��L��)��n9L��_]�~6-�x
Q��?�}�ͩɸ�[8kò]y�fo3Iѹ�ȩm�Il$��`΄B�Uj�Ճ��_�������^_E�xN�z�&|����3��/P{>����k�#���sL<�{�;p�O���~�x�C{8�(sa�p�M`�yN{@��߄�c�\�uA���%E���g^]���w�cT^�j*
����+ۜ�SKr'3;j�F<=��38\_���|r?v�@=5]�E#�-��霫�ʑU��и�+�\4�-\z�|���U�槥�	�m&�F/^gp1b:~�;M0�'�s�6aF�\�R $�m���qX��nL�fW�%j9�?$�MN߾�4u�=�c?-/�^>D�6ɜ��M��#��"ٚ���X�o�rwVog�u2����#cύ��˯;�����b9��S	���\�_�Ϗ���9Z紎>��۸<7��M����*)r�{�|�G������hCp�0�
�i�#�ϳ.f���D�N8��W��kjY��1��>��.��N>��jĔ��H9X�7�qP���d[����cn۪���#�͔
h�g.(|p�A�2"�[���N���s�0�u����#����=o�g[s�FG�C���G�#-�yd�4�*O4������܌�6���O��qD�*Gw���f�9 X��-�\����1�z����{ �޼����#�#�=�&��}11:��≎Q�z(�˻�a����}��/
�m����Fv����g�qU�jcDR�غ5^����H4�
@�����r��'�}���ݾ����7��P��O��9�(��
�Nv�a�.�U�3�`^�z�!r��Zz#X=��|�I+�ٝF � ��sy�9�)Lt�0�ve�߫�g���]0]3�j�ݜ5Ϋ޹�W��z�
�0�f� �Re�pDI�� �4�p�X�b]-�IY� �aM�h���Ź�N�	�b����{�F����r}���ʣ����"�\�ݒ��g����e����LA7���ºx�K2}��Vfw��y �
: p�&�/`���x��g���C�#��Q'��Q���v�qc�,Z�
�Fz4��_�����Ct��7V�x���=����tw�:�~zg7������~�B�P��p�"�:���39JV�=Uc��
�ϣ��P�[�w[�-�c9�AS���G�w�h�H�c\�5|�N��p�]o���qs��yZ��xF��Ǔ��b�s[�������A�5jQ{���&ŏ���a��<co��:�*��c+@Zd3�5h�9憩�u�\�l������(-��,&��9�lЂ��v\��j�4ߔQ�BtזiO
������۷�G6���`Z��Lw�:��!�F�6H��oy���θ����u+Ī����~��й��,�����"gv�����!9^E����u�
!�E�9��/Ov]�E�����n�ؕ���sQ*�I�'��K�u\���#�[���w�Z�~��!����a��f(���t'�"|D���Z8u}{��d�r�G��=-�;�w�;�;�V�VL�7����~|�#��C]ʠ6:.8�\[�t�3�`?߇���������g7Em�>�t��ds�C<�����U�NH�{���<��;M�K�����wP����4J-�4~��@N�����^��| ���Q�����F<ü���2�կ���&�Y3�s����?Q0�����`4e3�}.�ϪX�V�
*<p�>��Qb���7�L$���]˴f�~ �X�&��.}C��0P"1b�*����;���B�(��w��Y&�����C�Pn��\!iڎ�d�>��#��������Pn�G!��̍tĀ���uS���)�
h&V,�rt ��ɓ^��&���KY����2��P�3��c���s�Ǐ��Sgf�V�/9S�[�q�!�)^ִ׼+O(8�T��R�ݒ���E%��,rݜ�WN�>'�mT��`��؍�*�u�Nx�l��.���>N����ʷ8����f�@ui�h�;������(�v�x�0]l�<���;<ת�W���ḇ�%����	Gs����i+ǃ'mە �vs�s�;GJ7��N���갬�H���֓Ksv��2���;0aGPO�;vNZ㳷غB���p�k��J���J!�cd7��o����DD�?�]Q�b"g^���������տ��e�c��ir��!jLF&7�yn���7��M��d f�Z�w	� ���6,|���Z���ӹ٪�q��}u]x��x�֟��kE��t|O�y�𩣜�'�#�c�d�e��Ǥ�lj�b�E�3����d΄I�&���RAL1|G���T�[�u��\�&􏾌�lD��D��9߁��8� �v9%�z�	�Z��Dct��d	�$�?��`��3��O��鈒^�$�x�&}wBi���(ĳ�Ĝ�r���a�٥�m%�&�"�Q�(����H���|9}��[a+�ٳF�P�0L$�{'�f�5�ˏ�Q})S���Ս�&/e�+w���Wַ��Vf���YSZ�&k<�03HB��3��fJ��Op��E��&�~n�,[Gy�ݭ���~�7�����.=7��u�[?FA(Z��C���Z{n��kMXB��a�$'�y��}�iZ
�s��2DH^E%.�y�7b�03�z%C���^
�/�O�[d��g�#�q#�9-߲����w�~��b�(�{1D&1x��v�����ɑ`��3!�Z�c�1��Z!���8�%�_?U[��;�C!�@)���l�s�[�{��ٍ*�먜��b����������������v���X�Q����lQ�ʪG���P��wC;6��c�gk=��*9ٵ�)~��!�֝�|�ά��8�����F;�M��ܳT{�|x���_d �b`�hpt���E��u����(b#	e#кT^�� F�����$�C����tUG�:�'Tr���E��.r���ܷq���?_����?�]γ� �n��.��/c`f��ڇs�V��"�%Sd�-(gke^moX����f"�mɣ���m��������X�B�ݐ/�$�3�D���Z��k�mt��gtB�a�.w�Q�]r���F>��=w?Q�Gة�~�O��om��B����&I���LK�bs���BN3"׮��.�r"�zz�X�����d����|�&��7���r�z<yt6�%�\&�ϱ���^��&]��*��M�Ń'�����l�MK�K�mG�A�G���4d^�D�G�!dҮ��Y�2�9�j���C�GEϞf�f�x��Ș�F�7�i�>��y��cj�ؚ�n����M�K̥�Ud~�t�]�SB�.�x��/�7}CM^��z�Ԉ��`ne�SK3L��7Ͻ%4��94�&��^�Dl\3~��{�0�Ц�[b���^@��!'�w��W��r"�<�.��H�{3�~k�+��.�<Y}7�a�ƃ���l����bg'�kRz���/k�2�'cU(�K�o3���ӎ�`������m���T������M�~�0wu�6��/�C3ו4BġB����;�0/������`�&S0���[dz�F<��:�T5�	B�V;baP�64�����U��֤d'ifm��Y�F5��DY]]��E�u��L{O;��	9�b܉�����z��~?��ܽ��K�:{���/��+*b̯�m]����	QN=9�F���#�_�X_�^�����v�� eL���*�D.g���E��P[ ��-x	~�6O��q2���2ۤ3PBR�������ǷFe$H��6��5�O0��vV�՛��'$��B$hh�)V�&�A�tE�!�f�B#peu��#ݰ:a��n�J/~H��js=�u�=�#�� �{�?`�����o5~1����|���ng��9�밣�2�D�B�9�'�$Y�޼!=�-�jL�.B��"ѩ��_�B�����y��#Ő ��`���OB��-ٍ��]0��yxL^�zDS)n{�l>!��G�vb��!�77y����M�ꉆ�B�G�mw�����b�v|\%ʙY9�4oi������	�A�ᯰт�E娀I�®⯻/΢�A��0����4��=w6�"1�_����p��٢�j(�}34�a�c�}��n��N��X�L;>k`dՏ#ل&
)D9���kv懻;�t�� Ph73���[�ܕ�!θ���n�������yAK�%z���9� �|"ܦbv�J!n��0�]y��.�k
j�2�׳�ep C�@���C�1ib/�!I0r7:���1|���_we��b��d�����$�n�ɖ���o¬�8�&��yp�">�E���P��Іԭ,�7*dǀ�r�B&�!3*�$Bx���[�.,��>I����Di��Rn�#�����0Q��!��W��	�����qAs�D"ɨ�������"ď���nv;�^����G�&�~W0Ѭ�Y�k��#p��)��C��9�O�Zv̇y�RNVvh����.<j܂�>7���
��<��*~fwj��&<����{����Ь�	d�����6���9�ib�F��Â>T�ȍ��*�����7�]c�3>�3q�I`�����޻؝�3�0X �dG����%D �Qf>�?S�ɩ���Dp"��̝��b=u�|�>b#���L�2�>�h�+g����u!�(�< ��Ik�]����`C��zy1��;�P��#36� >��o�_����P�}��cI��~d�b�e�g���������b8�lC9�Mߔ�����Oơ�`R~�;�g�G�Z2KF0#��Ѵ�>9B����t⤽u�dǲ�2P��<�.��f��A?�0����HD\bT��D<'2�y�]��?B&(<,${7;tQ����sRd��	6΁4��k�h�2x�Bͤ[sh�CK���@%An(���2��?��"4l����h>�����?�AHdi��	T�2�&-}��T2r&#��Uq���q몡u�ot��8E$}�ف�*d�7��119y"�|  �BD%�Ewe�T��{�=K��DI�9��z'R����n�-��?p���v~t�uZ��?@�z~w�dCk��5�����j�#��l�ߔt��O��	�Q�����A��R(`r���h" v��dK�nr�ɣ��"0)S97��B"�FH�i�|��1[����V�.c:9N6�^�P�D��C�_{r�1��I] 0C��0���ЎiG>owv��4�7�KQ�[����&������]!���Mc�sYd ��V�]�����`�*~���N��Y���82���������	X���#+� �S!�.��hP�����+pu�h�p8�z�,���bܗ��R��9]�Q�f Y��s(�ن�;b�\,��[��"�4"���	�1�������V�Bu�E�:��=�ݡ�h�l,a��f*�j�D�8���Z9wit΋��{q�p�Vڳ��9ђ-�¤錺�aͺ�BK0P���l��O[������������2�;E� ��l�#@>b��8Q�q��*�����$�:ĸ�r�}���&bك��^(cDt���3�?Cq�#۹�M�G���Ht (�H��������՛��HyĜP�u~���s�ǈ��Z�HW9d��2��"�R���I�u;q��Uѣ��l��"{���{ު����F@�I���pģ�;�
}}����(pK��¸B�h����_6c)� ��Q���z�H����0 O-��~�w�s/�s[<�zya�f�t��!anK���#n� &@� 	m0wb$���� J�Z�VZ�00�����/�w60>1��d0*[��ʃ�mEl��P�AH";*,w�_1>O����8�|R-��f0�?�q��Ro��\�a��K2Tq�;13��R()�cɩp(�J���"�^fE{/�WϑQ�8]�a�L0��/TM�x|DP���A���{�6�w��#�aт�FR Q�W&,@'������^�z'5�3Y}�޹���1p���ݹ�,]V�C%п2z������b�8bAJ��Q������g��І��3y3����!�/.�m��wC-(H�Cb�"�r4"B��[�Ue������Zb��w�XVb2���G�4���������R���o�yƶ'Дb�����,b����1��|>�/��F�m��!��y�@,ÈMɣ`�fd/r�9�f	�H�D���& ����c�쏗��HJ��~�@wna����͡@�����y_e�w(��P����
��`�R���	�{P۴�5np�+����ҷZ��,��G%��}-�}Sʎ�����4�9(n�ɛ*dz7,��~��ZG��Vn:�C���6aqbۮ����g�Oـ�EC����!m�C�e�N>>I�o���� ��b��B[�un�6�s�۫�l�rYkrI d�Ǎ�1�{vŰ�A�,n��ۼ��'^1��� AV�OP��"�_sl	e*뽗�Sq��OѢ[���*�3*xצ���  Fr�h�L�Zw�<g�����{hDfg���O6�Tb�	�K��Z��
�N���}刈��`��yw2���*M�9��/9����pH�"kޫn��aM��������:#�M�a�a7�(��6X��g��z��!{3���\1X���a?L��z�c9�A��ˊh��>�)��C�̟d������L,?h�nQ����T-���P*.x̋�`a~j.W�=K����	]�t�X1��ٮ��Lx3�-ɿ�>�^��n,D���T~�1~�q~�dL� A�c�9��8q�_�=�����vۡ�F!ܾ��0���wE{g�"�p�~c�c��9���Gtos��@��hő����T�H0���� �Owc�s��AD FX����\�PCr��;j" �ߜ�!l���
��Z����Ai�쯶<T�{��_<���,A����'4T�U}�U꛻�:�N
L3��&-�c��"G�+���꫶j�(V�(�.:;�G6k��6`<=�z�����d��s��h��N�6���yc[�`{'�1
"75�]�<�����g�+: YQ�~b��x����b��|�V�c���cN[iUe�gW�|�д�NScQ����ޝV�*�ٷJaP��&k/�p���xz��N��	Z7K���ym��If�:�g�W�����
�똚M?��a�8�K��
��uGd�B�J ���PEe�"�_5DC8 ě�U�R�߅���-n|��Uw�yx��7����=�͜��Oaߟ1�Q�yڈ;����!�>��fc�-.BP���![�3G��Ȉ ��P��A���6�L��{�W��H׶c��fOMӿdVȽ^��$�%шw��.���J��*��I��%�s{��$Vs3">����f��Y�M�sA�ݦ��
��(�o�;�
���%$�i2�˺<�25�tl�8-������������ɪ��"����2�s\�	��(B`Djb �!ҕk&|"l�{'��/�M�R���0�z�;x����B!C�����]~黹RP��(+[��hX�W(���<�=�En!�&�*hA�2TU^���8Z4[B^�T	���8�˽��Y�m!5�5\O���7ز����@�A��)E���d��#,��轻b�i*(# wӰ�=nyQA$� &H_���Oi��9�me̳��諵��DBp!�4�@py�P�;�N����qł\\p~�?k��1���SE}	�=��{3�v�fTA�>��aǽ�,�s����"�Vn����M~����,0� 	E6�4~��+]�Ra�T�jP��nvFo�}2���Dĵ"��y�8|%9�w���H#D_�'Ԃ!z
���,}������O��؋��R�w`��hBpZn�f"�X�9����u� �˟����MvٺM���q|�8��FF,��ޤ��H�Ӗ#�7ɦ�mܽ�U�V<�[�s�t��V:�F���x���t�F��1u�Cv�p��_uy9S�+��^��[�P.��Q�ٵ2dQ2�G�w4)d���Pl���16�<�>Gz���}�x��uj��}��'d�Sz�im:	���]�y^��#B䢥<��������O��ɂ����t��ܖC��K��ŋ'%��8k9��2����PsO�v {s��	ǥ�ˊc���w.��$��3]6��,�1���\�w6��ͭ��^�V�z�Y0\�/�`� 3'mq���"K�Ckn�:�ʛ;�*ن7�_�va�h[���fە�Q�EM��B���-���y��������c��읗ʻs;f
.½N�����҅`�7Hiڕ�e�`	eE�����prr�M�x�R�X�5/��S,��õǗ�Y��I��s�+��<Y�h��s�&�oĂ賒��7����J�Ӆ�<��	o[���9�v��݇s��D�.���0]Qړ�IJ���T����g=��9#�{F�>ϗ��>�0�12)��@"�owg�xf�ǥ�fa��ğ�2m�O��ۺǻ!�:��8̾���m`�	�^+U�{��	ֲ8�7I�R=��=XJ��W��ӆ,<��҅�n㐩s�Yw��K���4֪w��o0A�1��p)E.��B�o����$�m ��14m������{*�\�����0���a��{n���w��~�-Ծ�8a���̧Oq%"�4VQ�|��[ԟ�G�����p��h�?<��uo+�@/���4h`�g�����q{2׮����A���I»9���5��e�0���uq�?@�
���oV�eB��&W�Kp�_z)[���Dv�)���mpX�GB,��M��6�Ü�����@����K��/���ـ���M�)D!�E\�W\B��G��&��ME�=½�p��E���9���N;�����r�y�khdxze3�����=���"؂�2ڂZ�A�P���j5v8��Wwe|-ۄ#�l"��gj3��oC~K?GO��s�9q��v�$�� �̧h�R�]u{;<���
�����",����.b�!��>~+�O�Cv�/(����b#����+�TM��R�krV Pa���Y�QVezDi�Ó�e'
�bS+��+@7�(�ͤ/r��}`77oY�|{�޾�#{{2����:�[��X�߁��N�v���-�sN�N�5�{�����Yt<O�Mݶr�o�ڒ7~��
I�I��LA�D��a%S���ĻK���2�}�8ʙ�R���=�[�E��F?'
d���%a�_G��'<W�L#��+FWf��2<�w��-�z+����V�<���W6!����C���%�HYh�`☶ 
�̯��T#Q�P7/��]a�_��UBX4U��΂�^Hې�U�,}N��б�V�K%�]���.��J�T�v��lq����.,��}�ұ�uE�:6ln?[�i+	��_h8͛nIx��;]ΰ=��-�P�*�S�ϋ#ں�k���8yXT��	N�L�و��2�WO����Q��'G;C��s��%۷>�v�,��=@saB����Rlk���תR�>��c8��=s��lո�	��L��S�)��<�L.�>���B�F���t��k}[tb�< �^��;p�X ݍ��Y% ��j[Y	3k7{%�%�ʚ�#���Gג��>>�a�W�yH�)Z�ΫU[L�O.05�h��$dcW���&���tzP�SH::�Dk��h�18��T��vU� ���P�kS������bO��7ƍ��<x���\���G{�0�?JF2,��Ⱥ5�j��22���L� x	�;���!93Ys�{'3R�F�7��$b�,�LtP�mBq���9�:/]nQ��v�@��y���]�`eCd�<3���U�|Q���Жe��f�����vT�;�{�~�y�8�+�u�1B���cs�����RjI�w_7i; �_wP�~YK�dJO~���;��e
�̕��R��e�|g+he������~�͚�ң)/�%Tc��ݾ큼���i��8��^\�n��ÎT� ȥ5	��Py�DJ}��5�d�۾�΂#G�ڄp댞��y5�O������~3�پ��ڛ��
�?iz��!����=0��ڝhT���Im���:sVJ=�g?O�N���g�դ��#��&Ƚ`��3.Ľh�ų�
.wp=��]����L���0����#�Gߢ}��LUi�@�5�D1k�}�f,ϣ��@@L/��D��hG��VA)U�����r)BH&�/�����~�/����2�ö�D�B����䀱�:{�d��P̣K���4^*l��=y�b���o��h�o� ��m�/�9�nj��7vG�95�	� �T���f����L�C�-�l�9-=��� �Y5��L)���M��͸a�4��ߏB&�X�M�\HV��`p��xXɇmmm;gI�����2�,�5�ӊ�E�դ��):��Pi� "�ɂ;ww��zt a	�H�cA����:#�G�³N�*�q�-�s	z	T��b����g=�^��K=�O(Nh��m�dw�w�ĩ��!NFem���-���^�?*ÙW]�P��\����Ω��(�k�+��5�Ζ���vvvO
��LC�P��x�ͯ!�8���EPV�8Z,���˓O�cT�-�#14�M,�R i4o평b� ]���0����J�S���8EY��ijB{�m�y���Y�;i6�q: 4�yF�{4se� Å���4�zfMm�2ﻷr}�.��&3�f�V~�Y�ci#���p1{0�(_���5N}�W�T��C	$��c��Ƕ_�J��R���]�U�9�&�
ý�#���W����y�-�^��u���QqUo�c3���{=�20gڈ�P�Nd���{%��tjA�p�H=������<1��؛0�}��3����FL\�ˢ"뼉����p�%d��؝�ժ;Y:�厌�$��(�Ƥ�4ZQA�I-��%�E��ힳ�3�)Ӎ���q'B�&�"/�i��=.a��d����^Չ�B!��z�ta_��]���>�V�$�uo�3;��\H�A��4�N;���~���RkJ%�����hJ�Q�^���y�gDϲ>==2���D㳏���q+2�Ǟ��6�:s[`�o�W"���^9��TL�M�ȩ�ɒ$?x����w��F�lx�{l�;N��f�<��3R�q�y0p���t�Q�&(D�(���^�{g7n1W�*l��Ä�Mr��Fmv���ݫ�}3M{Օ�d�keqBD1�/���kǭ�\�4��iǫ�������H�sە�iGevڍ�c�G��l�bW(}��S�v'�h�m#7w'��\��+���F�Q����8�s�f-�nGv�7>�$�7�k�K�a��
�H�eN�흜�3Y� G܏��}\w�t�F�q��A��I���n�C�c�;�q"{�7�@��U�dш�f��(����mV&���Y28H���j����k�F&�q�)��+{j��[hYJ��3繽�cv��k�wۿ	A,��>��E��<�]f�Dׂ�r�6�m���n'w�(�f V�
��$���{qIW^,m�0�!��pFhy�d8�w�~7�Z�p���U�pC�r��b��`���o1��̉f�mL���V�_x�rH�vE�3�y#1Q���Vhdnq��h��)�;A��pk+ܤ'5��1�P���)V�u�#6��,)�o���-M���9b��z������J�1�����X޳�u�S�uQr�k*�E����W|��H���"A7���{2�߾�<o�D�j�/MRa�%(&�G���X�\V�T��d��B���v@�c�|�i�5�nf�>+.�M����=�m�{���\T���vP�}��YIH��n�����͙��d'�;g=�9��H��yJ{o�M���w9���e���>;�C�L
��I)��V}�69	����h��:��=��R�\�������RQ���ި͌�oZ[�X�k=�f�c�@��f�{ ��ꑢG���+7=NV)�(h#�zM���K7ჴ"	*L��� �ݰ���*p��Gm���O�t�J2��#�1�Y�n�q�-ȪJ(@&HYz�Q�v�NC/ﾫɼޘ����ʰf
����۹��<;��F���0T"�A74$A�fe����r 
�a����:�p(�X��8��[[1�[�E��>Y����mK5�6��)
�:|oTp��~�̚�=k�?)B`�P}��T��aF,p���򷶕�tA�o$5[�테GU��
�e�L��;�4��B0�H�a�!�S������~��p�s��.��K��K�޽J�s�f�p�AڞjR�0�lh����Z��鹎�@�����6�Y�/S����bt�Mm]1�ܺe�H@hE��d�τ�R�W�����d�{�\��**��9(_҆d�^��n�����3DĎ��>"��f�pH�����ϧ+ø/����Jg(Pob�/A����Š�P�iJ�\f5�˘5�x"d�[vmj�!���iYAtڽ� �d������5���ا.�{bK�p%�k��cFw�AGl?k���ů�@`�Ǽ�w�x�hy�1�{i+73fʱ^"��J�@8HB��ZiV6��rck!iY�.7mrf������nDb@�<�ڎm���d1n�F���ƫn���n�T�o/\d��ق�{8�<�����F�pb��a.6�ײ��Kݩ1)�8�����jfm1�ea�A�����9ٹ]��x�x�ݚ_#����:ݺ{����c&��܆{f�z�A�{pu� ,"a(A��jB9��b��1Yn{0��Xp��`#O��$z�q�-�N'�������q�������[G��Re�t`3p Ǌ꬟��9�$Ng��UÕ��&M��������nB�S�/(�+��,�߯{���V��|s�Пw�тpüo�ݵ0Ɉ�b�١CLgiT�	�a�aU�g1�����o����p��27��e��j��EJ` !���&��s��I�t�n�A*;#4��r.�/+�۞Ϳ>~����8�܁�F=F1�"+�{����0�aSb��_Q���]�"U���<�3�2N�b���_a[6}Á!��E�>�Mt%�����E<����iH��Rr<恝�͎��U���'��>�)����l�"����PoP�P�����z+�*"t¢n[cqK�ӽ�w�Orf�D2!�O���8Vb^7��-�T����np�V �N��g�D!��ݹn���h����W6}��઻�:R�(Q�!h�2�%�W_�o��S��G���e��ڭU��9��C ����t�FoO�ѣ���9[�<����� u2�swަ1mr��3�q��7����@d+�6��sz����)��*��F/� ��)a#����ͭ����R���oH>y��NV	�w�W��f���}�L�J6���Fh����5�2\:�R��8P0/��U��g$#/���Q��Fk���۩�+%��~�	(#���g.�ٔ½`�I���9�xB��}�D�%���Fc���mgY�\C��'�k�ݡ���qj)�ݾ�y�Ǉ|�i��b�P^�� �*���"� � !G�����i���Y�Wz\O��Uk�	f�Z@��t�yͱ���W.'��0Y̶~Y��j�����$�J�#�k�.�����l�`	��33��ۉFKGA6�މ�e�S{�lpu��!�n�j�ʆ����s:���!AR�s��rf1��������[q_���j�s�zI�Qn������}���+�����߿�S�~��Mh�P��O��؃V���q��EƜ��BL�ɽ��ˑ}��j�s�������\f���gQ�*ѡn�vl��'�?(7��_e�h���1zN��g`�}y��[&����B�e�w����%�wuu.��w
i��¬�D�Y�������)�Ot�#Q�Ys2<r�0�ōW��S�2u�ݑ�&^�VZY���Y�p�'��鎙)]���O)����܃b!���5� ���u�(tOE���gn�9;ꇋf|�jKQ�.J�i���r�IW����k%��ݰ��B��$��eצ;�9�=�;VZ�&��w=�z�sg�t������Bp�-SQ����J����TNx@72�=�J�ek�cJa@�
&ׁ�Σ�3,�X1� ��ӷ��� l�U�����}�J#����2��B���M]�l�+T̪75�p$�Y��T[�\8�}����*+zX-
]�RՑ~hu�=R�c���3"M��&Gט�Ao|c�7�/=}�<K����=޹��w���3w蚉��h��*
���vp�Ia�s:*r���;e ���>EJ}�ՙ��q�G��[��0M����je����v�G��&)*x����v��#�����蜸3�_fm���;x�
$�Y�U�<ҙ�IZo.nխ����/�
%j�pFt���מ���}.�,�H3J2y�M�+�����0���
��:V�%=ܺ�ٙ��Q�:����1к-�(h5�w/@g��\ߏ�Yȳ���9q�������
��K���:v�ss���12-�p��O�ْ��q .M_&pd�!�>����+R���U�s��T��N!�q��D
�w�R��y����b�^��m-<�_�j�<��H"8r��b�����NE�±^���f��=ӳ	��:��l�=�P)�\��
]k���7�}Cm�p�(#��Ab#�i���Q�o �oj=�p�z����H�dY��y��m�0�:0s��x�
�s=�����pr0�H��jV==��$n,�3t�����y~w�N��(ܯt���8��捂%{&8���ɣ�Gq�S�����l�m�]�T<h�e�{*�A��q��GXU�&i`�'WL���J����]�\����N�w�U���%��u����Yg3���Ba��i{Y
3s�*}���%7
?{x�':ӛه��Ne�oo��݃�,Nl,,L�C�1�����.[�u�U��v���R(,ᘌ[�v�u3;��}�c�n�V	Y.h����T=SN��@�(c���})]��ߥ^x��|�����S������g�(Zbumfܓ��n����'�A.!���ը�L�̫��v�\�[����z�}������ʆ�8�g7��>��w�$��A�lE>���Mvz�領��f1��!�՞�W�<<�	N(4�	��$�mo�`Ma�'!���*=׹���^�Z���՚�L_ۯ����-G�O&���L�K��2<�N��nm����:Ma�9N[�쌽�k��<$2�n٤6҃iT�m
��؎���J�+��<l���ߝ��lg	ۋ�{ ^Mx8۱�,�#���m��$�j�Ӈ��,����Ld�0�j���N�y���c:��Ip�g�Ž<j���~���Uˎ&2:g=�b��6uN���݀�	��.A�7l��'���f�9�T�x)70y�C�%�g.��(��Q�ƽ��EF\��̘�k�g��-����ya�	��F�m^�<�ɤ\0A�_�׷��}�� =I�et
��Z�g���יM-����ԇ(��*$�h��fm:ۈҤ��)
�o[�c��^�i$n�ފ��wy�m>�a*V�{ z���1$uMfS�����|�)��PSb,1��4�2�:�bə�O�����"�K9uc˽~v0�}O��޿�E�hs��� QN�yv-���y/Lܦ�x��(G�UA5(�`QǴ.�(��C���mP�4G:w:��Xx� ���X`f��@,vⱻM)�Sh�t���ٽnȡ΋����^q�V�q�˩-�F����fe�n%��
%&�q���NAnݹ����p����<����(�Z�k
�l�d��[�!��o6��<xZ�G;#��&�؛Q��ٕ�&��������<��R]8�Ä�v1mѥ����ے5Y��VXA�kA�Z����z=�y����uj��I@��]]�h���m�p�1�)+�i?U�׫\h=!��FQ�SE}dLF�T��J��M�H���Hj�LG���6�W��pW �<�sZssf����Q�Awq�n�R:��A����.�z���rF�{��M�A*/��⊬x�U�3����7,rRDZ.3�#���r~�=F�#�Okp�㗪�]�:�1�.ձ^.��&�R�*��@��鷗yQ h��(��h��O��s��)`1���Dɯ߸������~�i�7 ��́��4��o�X��8����n%�A���D�8ci̯Z�:o��h���
���=u�R�B���\N]Z�k^��ҙ������+���o}�\�}�Vᣠ
������.Q�)+�ًG�������Rݑ�AGQ��vo�3Ҹ_��R�A+"c��G����J: �,��gz�qnS�;5%���qO,��I^mҫ��SM�CpH8>j��m�~��Y�R�Y4IH��0��n�N�B�Ǟ��vb�����	��mɤ�h��o�A���V�ƻ��E[�3�ϵ��/n����ܑp�
��b��/	j(OA96���D:.g)畈�X{
z��	�2ļo�b�\ƻ�"�5Af����?7U_� ����S��.I��u�	 e#�^9��Yk��ȇw{]+6F��h��c��F{�,�s���{X�nK��߯nk�v��Z˰��v�9�t��jV��]}'�����P��Fy�p̷�O�-A����溳i�p�>xn�r\�\�*�/n��o�x4FF�6�s�6���-�\2e���˜�;v���o���kqk3`�]�}ޘ�{l�y>�uʞ�i���I�H�%S���:Lwk[ꢞ�!'
�ò�=|Wȡ�t�֝*-��
x�M4������3[����f�ݾ�ϩ�װp6��Ý!d*d���1��䇐��Fq}�Ҍ;��axe�k�u��N*w,��]Idƒ/_eW���͗:�N��_ˤ��}m�6����[��ݡ'�O�������J���fR�L��~�f�հA�'ݝ�6���hs�Bn���O6M)��U�jGv�gOҜK��21}B��&rG�o�k�NO%���j�۳�b��ooJ�7}+C�4n�%�%G觷6e�����=�I�7=9�閮~[�������}p�b�z�޶ا��솎Z�������.FT�5 L�t��ۺ9��ag�,R{�u������'v���\��t0� 1�c�ӳ~�~����B{f���\��̅�Ժ�����r����l:X<����|	���rm�vN���n�~�����8��g[a:�H�ה}�ǫ�J�ż�ksq��� �f��j,�ґj��"�m�(��d�^љ�0Gi8�U�����=��cm%U�vf을�v�8:�F�&۷m�ôr�}Ӄ�<��&�<���к ;F��wx��,��X����&ee��i!��}pr$�<�I���{P�e�r�`7�Ri�S p��8�e� ֆ��l6����)��nwc����!���E��I
ȐnJ�!�Y�ɣ5i��K�7]�4٧WLP�f�nʺ9&C����ָʠ��ua�w'l=W����ʕ�k�+լ.� C�/;gp��=�̊�5kefF�+�!4���c#t�[e�j+�������΃9��k̽Y���s�`�h3&F\�[,t�zх�����	k�è��ңe"B��%� L�&Hq󕆒��� ��R�F6a�[,����7�/P�����6�v������0s���O��u����]�.,7���Mr�=s���\�����CN��/	v0q���/�x�v�z83 ��G8m;��U��d�ܸظ���۳Hr�*����֭�����W�#��x$�A����u� �[=�7J�;���\�f���l�C&&���f[�M���E����&�ysܛ��u�nQ��y���ݰ>^�;��f�3�s�[���c��N�`N��v�CBS2���J�V�&�HYf��]�j�i7��)��!� Lu��ce��5ef:�n����pz�v�ں�:%敓�3l��p/�&���5��G:$��.vЦJ�h��iE�H`kr6�[k��a|��	�!���O=���b���x1ڐ�W�R�p��&�����E�TNe'g=�b�\��i��s�y��s������pN�b4�,D��n����ۉj�]��uSm�ax݌��ƛ��'!�=<��=*S�r�FS��
BUt�#��Ζ&�9l��YL�X�, f��Sc�9��Yv���ݡm��|��7����\'ps����l�a� m�m�5�nFĻ<�J$����{���~���w��E�vO���ܮ�aS����i6��0���{S�7P�tm�JT/�l}D�}��Y�ܤ��# 4!0�DՁmH���8�4͞t�6�)��X�C��w�i}C�7�?a��GO���bb<��zC���T�ۡ�����O훉c<D�N;��8�}�x�^lp��o:�Ѱ69pa��f$��&%�W��v��ēj����T=�Z��"�˚��\�XD����l��F�����n]sr|v�Q��Ô�-����T��37�d�ed������QQm���F���6���wnk%/+l��v��weA������x�F��H1˔�Mg��ho"]�FhqV�vee_b����pq3!���{΅��w��T�gY�;��X6�*Y;��F'�]�J�ٞ5�$�y�Q&r�k��V�
�Uǆo�:Vo��sQ����o�4�����G�r���NR�3L�%3̘��wVS���8M��CA�D����U��w�k̩�j��]G�]�R#��7�ͼ�g%(�[.l���]��ң)U�������|�j�=~��|ؙ��k2%���G�.�ȝ�d����Bc���x?�����Yo[�_�$k����Z���M�q��!� �I.KŹm<w<�+鶭�4�=�7�-���s���&6oI�}��%֑rϮWAp�BfOy��*�Ǌ�ޕ<q|���r��e�'^* �=C0a�[m_T9���b������vf�꽴����	�ܖ��rr�y}�E܎�Ѧ�����@�ސ*i܁#�f)*w.�s۬���<YC��0 �a�1��pF(C�2���B#��<u"(k15���~�R� ���Bv��76�k�|�d�Q�_�d���,���D`���a�z�kky�v]�zt��OSD@L�d������/p���%
v���o}$��P��
�{�ݚڗJ �*.<�B2kw�>�<�B��Ɔ��Lݽ|��Gd��am3�9�̅U�'�t!��6�!�Nb�Ҹ|�k-L��j�5���l�ͫ/���.L9��C���?W��6��}vɇ؝�w5X^�X-s? �T�/�ڵ�}�!FԽ�gs��CG;�	�	���U�.=B��wL��u�y�^��eLXaSYR��8RVUmבC>'��������qB���:�Y�`�����N�J�q!/$2�ܘV#�}uQ#"���0XeKP�Q�pW�F%J<b]�^�+�PÜ�G����N3C&�� n�>:PX��n���vÖb��Ͷ,�����Q`*:��grٿ8�8�^4��Z�ۙ�/�������Z�+;f����.췤ҭ�d�Pv�v�ni��:RX"13��(Bs���t��	��ˮ���`�%@�a��I5�{-ϯ�����c���Ȅ�֞[V�殦1��N�8�-`2R���I������]63�1���HM�{�/|d��� ��wr�.�2G�:��3b	�_R��\�������ڤog�Im����/d#�����zTj�s����dσ�� F�n2�kί!�!��eʸS-�n�w��TB6ya*P����n�1����� :�E�փ�K��	��v:4��D�	��A��7<Nfz��ɸ��_I-]�o{'�8ǎ`��u���3+��kD��A�>��/o�S1 *+��Z�*��V#�X.je/M̈��� EOQ͈�?%� �3�	&�>��ʝC����;oDJ=��	�x�ϻ�+���o���ȓc,,����#���k�n��߆7�?<�bs/���V{3m$�WQ�tD<Bw�=�y�~���!���e�M�V�C��MvB��՟��za���ד2hz�뒹���A���*f�+m	uaaa���@k�ƶ]h�(Q������0��y�ou
�p0�6_l�3�ӣ����a�Tw쯫�+@Rt��{�K����N!x�d�ݽT�U�]�x����ڀ�S��Z��,.X�72v8�uw�"h�w:Kr0n|���.�ȃ9&�/ ��d�%%O���<�_�ewO�;�F q��^��f�6D�Z,!�\�����UuoAAt"��l)`dQ[��5n�ΩK!F���l"����S�zG��M{���,�<�!^�y���ge�v��ſ�j��d{Q�s�����Q���}�G#piE!�%��V�w�E`.�����r>��@����=��f��L���vO	�'N�}
}�#.��m��	{,����z{�\�e3���r���G�Kw����VL�o{r�X�sW��s���>G!n�`���cv:Ġi����ƚ���4%T��r����cH/F�1�T�3F3=e�6R�&%/sӦ6��6�\���m�ɰ[p�Xb$�� ڰ �r]�7ff��<m�4��y
�ذ�.��1!FC�5..4\P#bܢ��)f;o ����<U�N�l!���ز����4I�Y	Yf�m�`�ݻ=�v3�0�3��-0w�ub���E�|�����-�������ZMr�n	"B��-sw���l2�6�gwq�qG�NOq��F$+�6*�ޡu��­�c�2er�~�� A��̰����*�bi���r[b�5?�KwꚒ;;G��98g�g��D �$]�EU�܉\�N	I'ӈf��⫺�;'7��{
�1������eB�Y!)$�� ��3n�aa�*[�jJ�G{ �w[\�9��ݗ�?<�����T�״��ݭ2�ge��T���]K��R`���Q�"�chA1S��e�f�ulѨ���p�8i�U��vղ#	���P�2*�+�O����Q�gg���B9^;�D���y���Z���]��
���䆓��	���J���$"0�t��}�껭"��t/C 0�00�	�p=�dW��h}Rj0sl�va5⃫��[�%�_���y��p�����a}���5��&���w5Y�J����[.���xE@2���Ӻ���K���I����գ�c.��J>N��eb�zg�7�sZ���G7�'W��bϹ�A�@��r���y|&Ğ�ت##�Z0H���W*�6q��8P]%Z6��g�}C�����NV=�n�����*L �!�߬�AK�ig�]2X�5d���&�� (��Ya,NYceAm�)�3�i�Z��qN_>��^�mc�b�<��w������
\
�M��Uf�_7{��P��V���e]uc�����)�mc{H�ْx��om?�f���p��B�&p�n�=��
���]dʵ�z��۰#�������" ���G\3,�"	��	��`�,K�����7��kj�P���l�[��π�w5��ed/CY��S�.�ч�b$N�n?O���~D�����l�J��caq�CL�	G��A<���Z��xe���[�E!i��~��D�oL�����~C������.��,3��hx����7zft�{\�Y�幓uK�쥞Ǳ�C`�+���]���7��=��#�޹�~����MyY3y� ��;d}��yc�Q��O��Ng�)Ϳ�{�΁�(}���zVM�Pq��M
��s����tɉ�ɮ�W��iNĴ��F�Be�e��Do���P0S,�+��l���.���I�����Z!�d��TZ��]y���"Y�2�Q^a�ơnVhD��N*̈{��l\��ڍ��i|���8��[�f,u&f��������h���=R	�!�'H�	�ҳc��u�ՙ~Λ���<w>��5m�9��_Un��v�l�3�n\��>����浩��3p���z��3/Ύ�#,���v����"9sD�� \+���a�;Pq�����	c^L���p��A�q����ΎW�G����[ɳ�VM�9�(⺸�s�.�$�6����J�F���.��"���w�J歚ل�y�l��.�T�:Q���e�3ƀ?k��a[����^n�Ce#��U鱓�_^�43�v-e՝������yցw-T�w�
�b�G
`������9῿l��ݾܑ�� 6�M4Ӆu�l�6(�c;IR�y���o�P��ǊQS��G�z{�0�2ڸ-�9�_J�G��'�<;��צ�V�7�mu4^�:U�le�t3s���zڀ�`(M'�ȸ&��&+�ϧ��y��q�&'�Um^*�]<o%��Ǖ�H��,]������6Qݑ3d��v����i������Q�x�����$����9X	�
fmy�r����ѽó�;
;�������_��':�:�j�R}�{�>�ca���+^Þ}Y?z� ���`���{ۦFnv�Qp�4Q'��M8��f{uWb�����-�K���)F�S`�ݗz�@ Y�0��h/)g^���˻&i(����E�=��,Yg���P��I+��m��u���U# dB{��j4�~�/5oq&c7��f@���=��HJx�|A]pS#�͎�k@��ܚ����Օ�  �ltgb�-�뼗~���`,w�fJ�(��ݓ��N���v��!��3
ԩY|���dUgV��΃F�s��'B(�c{�l��[GM��mJ�r�8H�V�=~�*ʯ13�1t�6� z��z(?@��UoOb��y,{)w%�NU��u��vL ���hO����uq�;~i@i&����(��u^(�us�Ƒ������R}7Lnx�ĝyـy�$�0�g��xf��Qt��B��qdS\V{o+�jL�pP�+�iH�*c��p�T�3�W��ۛ��,H��'��-۠�\-IY����Ƒ�c�s����~�N�ӟtsrS���$�,�e���*�<*�	�\�n펕��v���j��^��YyPum�y�˹�L����[�]��Y�r�U��g_�/k$ ��w}��G��v�^\���p�E�� ��1Qh��߫�0���Y���������uI�?>���]z��a�R�y�嘝���t����~����fω/����ͅ5��D���;�Lϳ&�ƞ���I������]��T>��KC+���^��F���ƹy����g�7a6h� ��&	gs�x�ޭ�Ap	��nz����,NVׂ�#.r�g\onףּ�|2}雦�5܎Y��|�C�Y:��M ˊ���sUY�`���#j:i���Y3��7��uY4G��%�o���*�z���
W���yK|��cͧ>�mf���q���*�*�j#5��>�9u9��.Z�D�M_���%
�˹�.�u���Z�K�z���j��{���xeM���[�pG6v&�o'^f] ����,�K���DX�[�ۚ�`ҹ��M�]Ĝ������gkvae�cncUD"#
��[�DG����Wr7��!U@�ym��M���ք��T��,�Tn���ݍ!�)o�3(�7���+�;�E�{>�LI�F[��Q�0��$�YF1����Kc�[�.6I�X���a�Z���Q��i�oF�:��j�f��:��8��3�u�%��N�m�c	=!��dǍ�N��m�.�u��A`�׃W'/]v۶a�{�exU���1���v��ڔNQ���NL�j4u,��i�r0��8@�Z��ˬ�l�T��ul�7�^�6����W�Ku�w8��a3�q=kxo�
k͞��v�>=��W�0�#8o_�����GQ�D�)�3fu�wu ���.&�=����j[����'�������-�(�j����P}��"��#�~Xa��������jf���	�,�<�r��㨘�޵�'{ G/������U���켧����ƺ��}��3%��:A�j0�A�D�ˌ�=
n���G��6�d��<;fY��>��foR�G����Pj�a=�	:|'��w��{�<�I�ͽضn�P�۞s��O�Ogi���
l����Q<�R���}�Ūe�:�4ML�zS��y�3$�)E^��:��s*�v��c<���.哋`����*�Q�������С�6�ff�&�]�2,.�a@���_B�Y�r���y�//�s�׈O7�C�w~βD���FǛY��v]��Z�}�0���;�}H)��{��R�[�T(�z=<R�����^�a{�u�_�Y�{{O\�μ'���uN�3����==�f�p���4hy���UFQ�Z.mr�y�s޹˛�oȨI �d��F;)�������[�� ��$i�)����
��H�ӛI�v	���������7���냌 ���S����)`�EIB��=Y��omN���6��ADq� ��a��߅�jfꩪZߞC�����H�����0Jh�n�:J��ymV�[C$B� ����	lJa��Z��I(:"=��h�t,�s��\�p��1;���N�uW8k��}����8#/�O}�k̿����B^�n<E�_:�"s*o�j� gn�pr2�א���o{mm���AAp�i�|��f�S�'+=����%��{�r�RҠ+�Ǧ��k$��zkA�o��P6Nf7��Ny*�l@����X}���i"+��FYu�As�08d��c��J���t��T�o�d�u�v�;�b[�+q���u�.g�[�d[�n%�X���^�-^��0�Vcp;x�p���ːVO7��67��)��%�{�H��!j��"ski�Y���:�K�b�X��J�@��X옞{��f��ތ�=5��wZ�oM�:��.�k}�GA0 ��8C���z�n9�M�s t�g�E%�3�K7=��->��5��Pz��Id��8��d��q�NY��U��#��J�ͫ�ۋ�:n�5�"&��ܪ�K��-0P%��_]�;�)�����F^'x��X?��V�O�?pXP!��e����&�s����'��1�Wٱ���(PKA@D���sm�M_|Mu*��ڑ�<������H�C6� �M��.�! ���U���z61���N�Mb�ׯ��=x��Q6,�-���5�>B�ei{<�;��#� B̕
�p�/0��]���~�櫕��x8?8��T%t�R9�fs1��F枤�4Wt�fd��T�L�$��q�}�:�ӭS%���-or��3V�<��w�܇F�1B�3�vz��{�ˋf��$]��j�uv\:�w4�\�W�Q�5����O���umL���viH�C-=澝�i��[���k��X�\��y�*s%g��O!U��.��� k���2BP#9\��X���+ט���1���*��s���Oٝ;��9�;�6%Tϩg��� .�R*��K�4�{�N�c9�Ӌ>��2Nn���aB����1�]	�݌������S�vuy�e�0��lX���K�d�k���}yc��4��8p�sÊg�nn��4Y]ƥ*��*{���̴���+�zT�M�f��6Sro���H�����5���1r�#�I\B7P���c�e�^���us�M�,�tJZ_guw��J�M��0fnSZ�Y�)��t�ο#���R|��9%1֬bXWnP�X�3�i:���A)��2��<ڼs8��˗�<邜ʤK��u����c�3��'#�/M�y�i��_�V�~x[��߂�P��+2Ը�jb�޼�q���,���P��z���k�{7����L�5>��ͦ_X[���	37�������(�w�Ӻ��h�a�IYT��zw�1�z�գ����`�l�h�?����k�P���e�Gk��+N�w3ra�"ʽqv��w�(,���3:�~����]Vm�;R�j�%4ӊR��B��ޤ{�X�t�O`̙�{��k�l=�݇:�^Mx�]��*��tҵ�����Q
�R��M2hn��+Aw%�U��;9�D�w\�VV����0ݣ��9g���5ՓgLW|�"�/�/o{����܇��;Z�9��c{��5�'e���I�ͣ�����1]�_d#Ə^ֱ�5UH3x�L��)�$���[W�ǳ=&"�0kB�ҕ�sHE�g;@2k���L}����p@~���x��/Λ"rf��h��Ԡ���"Ӵ�<�,0K��=BS|�{��5��y��3m2q�.#)Fw�^A�w;���A?i�nؘ^x��
�)��RѲ�9,��s) 3�P.F[��'b��Jb��{�ޏ�N�"��)���u71�����8ϗH�e�Rs�G�fվ�\�;5ʀ)
����1D@dч����YG�Gf���o���uA2�so���V�����IL�P�ͮQmtƵ��ۻ�4Y	~rC�;�R0,�{VGo���q� ������I�۾·�塜�-��#sP�ճ��)�K�*�X;��G��v*M���m�q�d��݃��@CxpXLs׼�&��&���V^
	K��;��-�y`S��ߋ�>+�/m,K'�;1�f�0�Km��ʮ�u���C�2iO*�6{��z5>ԍyt�*��˶��3P/� �A�D�Mj����2���g�hZ���ٮ����zv'y���{����N��4u�g
;�+����!R�	&E巸ۤ�*8#	�i����èMq��>�f�x�S���(8*�m�T����/l'�����c�Ӽ*�Onc	��� �>�9ƷnK!N 裉w,��K����J
P�F��K����]:���i��|0�@���� �f�yG/�\m<��З�ud4.�e@̡e�a/�tfwu�v��J��QYG�M�JB�(w��e=���'Ĳ�׈���!�*mtK��$U�ql�&�E��$���_��(�nOm��5�-�M�g>�4pC/�$ǆ֪����X~���1�݁&s�i3(�)7}��c�����t5n�e�OfːM��e�q�
=~TүgA���i}�E��b=������A:����>|/���q�f���Z���uWw?Z�d�<��\f3�Z�
�{���_�L0�`!�$��Ot���``2䰩	����ٖ�E3�R�,���A�aa�j!�jO�ve�il}��|8��US����|\�������g�r;.��mnx��b���8kKb�J��E��8�b�"\/h�m9�ay����u��Ա��YJ�hR#uW%k��8�˱v�ui�h3h2ۮ3H�|�xy�v����InІ^s�ά�Ƈ2���g��o'i�XF�t��kG8����
uU���8����[��`��y�=�m���v硳���ƍ���3���5��eڋ�:^�<쁲E�M��C)��- �:G�j�W~���<�^�{צ��3�5�ݘ���oY�]�B#�|fj���_g�P�h��-qT0�ǱC��N{$���=�_@�޼���ob��)ZN���7[)j8q�\}Q�,Vx�2�\�k �%��Y��^�rFn��A�!�Yܽ���K��ۊ;'�%:���b�8ڹ�d(	�2ꢐ�����
�Я:w[o�k7gA0e�N%�AjӚ�y�4�=�i`N�u��zD��+�	T����s
(�}���"Z��v��Vem��lr�Tq4ل� �3�bI���\������+]'/T���}��0�D����k6���l�y�z�J�q�����9����=�z����ݠ�Pi�S0�:���՞��f�����}<�f�ѻ����7�w6���I�oTzw8n{�oV?c]��&�獊nL��"j�[�/n��ł�WMV�կ|�:5���q�I���z�ٙsS��m�G�Sf���uez�����ba?My�{�7{���O>��uW*bz�ޕ�nd��5���tt$�" %|�H
Ya��}Nt	������̝�-���/6�Ibj8�/a��^�:����X-��'ӵ�%H�]m��^���s���qǡ�\2-�)o�������hܻ���z�V��\�����F�5�v�,�a�S֙�ߠ�Y�k7���sj��1�]���Uʲ� G�Be��Ms���`5>�L�މ�}��!wp��,��4`�� ��v�rF$���I��]v�k��c�k���,"�Q�0���r>����Q��ǺT
��M�T2懪�Ș̈́����;/���Q��k�>;ǈH"�)8A*�zȮ����Vv{�ӫ3���زnf*w��v�!��~�̍@Z��Ӑ/��"+��[��]�}�<+}�Nm��2ˡޚܕ����<�����&g��|󙗻�x�
��G��S����1Kd�(�ϊڅk�fL/.	�x(����kۄ=��l�9=��s�S���GÄ�p 	��c����\޹ͥV�8�V���s��}�]���vz�X_?�z�g{^X���3�܉:1t���@V#Qc�v��;=Yt�v�DhE�C!����VPԼ�`�p�p�l��޳d�-%�V��w۽����-�79��syS�g-;��N=��j{f'�����h�[Z�D
�̫�8n�jo��k2/�Pr��P���3}�soc+�A��;��!�W������@�d�	�4q�p�]3�\�)��ꍟS{8j랪g����y/}�[#�V@�v�*S����B��a�_Ot�אձ�7��yt^��Q�N���j/��.�����*�(*���ݲ�o1�yo��#v{ְ��s�7�#l)ϫ��]},���sc�+���
���[����d���L��B�77Tw��F]�o��M����1=q�;Q�c3j�ٞ2�"�<g=7T9y9��rj�ɥ�*� �>�&��� #�u��j-�ri�x��~	ρ�W����N��8+��ԍs�G����Wb��P�K|yqɝr����q���л����>V����]������SP�p�N��XV�l>WU~���g~G�4�Jb��_��oǶ�;K��P������]�,^u�5���Pe�ݰ�	��:j8���w�����l8$\6��W\g�㙏v�^!m�뫾���5' Z}�o}vkL����Gz��	]6N��@c<�y	�'��bVr�h�y�S�y4=��%rIBH�>����v�w�j�1��S�Jw,�#@�2Rd�Z`�55�[���a�b�]f�;[��z�_G��ھ��'wt��iUV�[}/�O���:�jԦ�1Uԡ��Ζ�^\��o2 �'a�e�0�Q��>>HR��[t�޳&��(��z��
]�g�0�Z)l�l�D%�R���~o7:�h�ٓ�N�Soz�{n���J;�K-�B*�/d�o% ���P�$W
fL�zꏙ�2�%"���9�*k�mW�o���!g�^���ϥA��wM>�ϖ�^u������=�N�J����5~�Rπ�-+Uy���Un��u�"t��2���m���µ㡊�S��S93y�K���E�CD�B��f�EX��c�Q㑇��:���=Fy��Ӓ=XWlX��NÿU�?/W�s/|��?�����x>u֨)����k��^r����i7	�U144܊�m7s�;�7��	���`�<�jDX�c�.��v��S=�i�vx�ŝ]�3�ÛX'�a.g�O�C�����r�hz7+���p�)���O�eMz�n�\�xN�5\3��srcz�����+~�ݳ��g(�-���Xܜt\��y���9�u`�	@�foթ�*���I�7��aL��\]w�]�W�\{��D��F���nkwT���.
;4Z4͘�)V��cA��(��؂,���dME{IB���;�f�>����aYޥ3[�4��]�^�P�n�:Z;t�%Fm����R�y�a�D0L�B��Wb��]3ݓC�Cc��g"��'�񖂔wv��9k�:���N��������Dy� ��=�i����l�¾�3�x��Z��7�<�7	�Z,��"Tr�)��NܾBV�����M�y'==X&��=���Y5�r�<O)�zɹ���.w�.���������&��~��2�v�y�]��!��c�
�qBǰ���~���n��+q�^Hψ���x[k�h�T�64�vN�ݳn]�g6��`��p��m�4��.ٹ�%��}���u�[�){[�%���|KZ�8n3t�v�� :b�T$ˑ�.��X�x�[۞�z�3���,#hU��]4eR�̰�vk�bܘ���u�y���ۗ5��p3����=|�K��:s7[.N���0�2������P���h��5�<3'8I��s�8{���N]M+ߔr��A.D�t��dd�0<��$��$�̒�e�z�F�h#��V��8x����9B����.���¼="+v���%FU��^ݚ<z0���#��WO\{w�6~a4k�)w�J�2^`�j�|%; r��p_��9����rh�)�g�j9�$tG�9Ǜm��-�xÄ��f�K��ө܁�7#��]��Rr��5�ș�)u:/ݹ�~�c��x#�؋�eߨm�ք���(Sٙ��O	�uuxA������b�R,`�0�����7x��CQ���[4������s����s���%,��4!d��d�G�������6��#ׁ�Uٞ�q����emM0z�=��GR����9� ��}y::}}�ՐZ͛���r��Y՛\�N!�kۀ�j6x��sq�L.uq�v�`�iδ@�X/�x�
6��X{9B�ѷ��$)�K��li�J�����\��l�e$��ܓ=K7� ������s��\4�"����n���ї�{ᬂ��O���s7�֩�]��T����,�{X�K�Xd?F�FF�E��}��T�>��f�TVi���oV#�M��	G,e>Vc�Ö���*����gκgq<#���ޖ�'���	VZ���7�74Q��h|��6U��!���HԾ���3w{���
�v|�?���ZD�X��V��G;�;!n�����pR.G�8nvOc��G��O�:�T�\&A>j��ә�s|LU���PV�9YO��ۙYs{mϊ��dhi|	hCͲqe�5lG��R��}���� ;r-��p�6}����Uf�{��(OY��{��)�jB�3��eA[`�B�i�G���l0�P����5�<&.��OX�{S�1�׹v�h�a9o��z4W[�ˆ�Tس�]��F�5����6�,Yw��۞�v:d@4�z����ټ��:����^İe��W���b���yfe��J6iz�l��Vi�vrfG���|�&����!	�
A���9���,��w��9�=y�֯g�}{�ب��M�����J������CN�G�U�خ������ܝ&��tT�,�4��S�.v!f�P��J`�Ef�OQ�Wv��se#�qE����Set�4�  �@$[syW�L.�%�^ȹm���{�ma��=�W���~~mwe�Y�َA�������$��+�v�lH�ϖd5}}�<��u���qnJ�S��k�Y
��|�6m	U1>9嚭�R)�\z!����KA�G�r{i6�o{i���~�[��f.�	�фFW�I�N�v�����y?.��$xR��3xbzi�x_چ��se�n�3^w5�=Î����g7�*@ޒ�.���g.���7`��Se�[;�T�zx_���N�+�HK7�������r���Y%ue�={�薱]��/�T�"`�3�0�4w�I%i+�L`�y���L�@��/�	��<y@np�!3VȨީ}�y�Y[���%�4L��vv_��{���W5��<[�w�W�E��~3��.F���V�>�:H��W�Q5/��M#�%�d��S4�y���==&]m��ρ���F�l��S-e�y�p�����da�&�n��~D�;3<�{��l���Í��p�$@lM��<�*$>}���{�����[~�7lx-�&��S.�]�v)��f�Κ�6���"��i	*&SKۍ{_p
o�]#�])r����ƽ�?VeZ��Ok�#�%F����5.���S5�S+/��qP`� *�v����$	�Ӣ{3��P5U��~	d,w�;G\/ҩoyH�r�λ����Mh��y�ޜ��c�`��S��L��0������*�����VCe��H�+�_�z�8b<��vP��(��`���@]XΕ��װ�Pf|`����{q�f���&z_�XHN�_��V�D�'���M�/�-��P�(���6q��5dF潩�Ξ�h�\ϳ/�E/[�"Kw��=|cN��)�@�:M�|o��{+�l��;f��o�eۀ4���+B*�j�;U�-�c�|5�k(��{ܨl;T��|��%K��2��a%�8M`��m-ى��5C�]ڭ�]]Ac��go*f�Μ�n�u��jwN �xbw槅ׂT'��l97g��d�S��9F�\����=�S��	:5pr9I�n~8�����{j[��/�	��y
&C�J�`%�(�Mw�������*ŠF�����E^�y�m�xѸ֞##�\ӯ!���o�u�*m��1¹�D2���R��*���Ga��@��������.{_����{�2V��Ou]9�n�ɦ�V�7�lv����D;�sǱ�7���5�F��NȒ�ns�����H0fJ\�V+ڝezY��1g�~ծ��-\����iώ`49k��S(��ª�P�^ en,�����=�TX]��ׂd��WL����,&C)����n7�%�y�pHXB��M��H/e�eX��u��D�nT+�U�Z�sZ񷛼4V��@�A1�1d��O��q���x[��6/n;�ͼ�Ϩ=�u��c�xy��z�����>���˶pLf�7�@���{l� FA��Ş��d)h(	�0�(�wT%��WL�T!��9)ٔۋ�ki�~�H�5	tA����L�{nx��sd��m�tnw1x�k��Z��%�Z�ͣ�6�vԄٱhCK�i�/��㞝k�������秷<9ëx�*��Ѯ½�L�Փ�\n�bR���V����[Hv�M�-F�l�����2{���?�,^ð1��]���(�pk7=ݙevq�+@j$�J v�7��#�7Q�5��<�4���o�#y��k�p*͞Z�Ý[���|��Yl^ch�>��qUX郷Ҥ�*V������}��@%� ���'��*N�Y�r�/�I���l��S}Ly�h�D���L����5m6�[Q=g=r;�F3�r�H���2����i�&�K�:��c�u�@��*
`��k���+d(��{����ڧ��nBڵ����,��������r�1y���;�0r<hL��ra�;�ǪF�g��^�:��ړC�t|�W��쾷r�~u��Mg�b�h@��&O�]����l僮tFW��緯��~�#�e���(z��&˶��KP��t�@(�ze�a���<��hV�����n)�-�Y��\����B]	���p���b�w|�'}�;K)rЀ�+�ёي&�{g�D�A��s��ߛ����@
}I?<x��ȳ��M�Uz8���_$�D����H��.���tZ���68�&V�I47��)��TO�K#%U�N��H��y� _�u��\�>��n�#�G^B�p�%̲����9�`�0��ͦ�YӂC�j�z��-X�J�<��`v�C;]=oX!թP�cs��`�OK��\ŧ�ܾ���ߖ����m?	��\�N�]bDr�̯�����u=]��yǷ���b"��u�o4'�恓ܴ-ˮ�;z��������g�/}�%��v����1��q��ׅ�nA�ڴolfw&x�{�:V/ЁE����n��ʦ��ѽ^�x���k��;�>�j�OV��8FD�B�r�����O�8#ً�O��'Pc��Z�ẺA�oh�X��q/E�.;�7]+"�q����:�*#�[�N�޵�ms�o2�ች���{����1����ǁ�(h�#���\�C8w�w��׼(Upk.I�0F;e�ɤ��۷�7�a5s�c�ْ�o����gۼ���{��52��������w��
u`{QƮt��<�&˩��0,�K��S���ර�3��B+|F�t8��nOk��Wʰ���O79�����L���u�MΝ����]���y�sx�=����`ٱ�ѫ�� �7∙�n_��Ե�{I����j�hf������]�+À��Ӎ�ԝJ���u�y�h�@ǡ�=Dz/���w����[�f�p��9��_Hp�<�s�	Ѥ־���{��ff��=lV���x�lqY����'J�e��cn�h�{��$�-7��y�0�`Ǖx��vۄ�	�K'f�&M[N��E-�s�Q�St�ܸ��<�m�u��y�N�nd��ll��lc�\��u�����ⴋ���:^���Ri�n}s���<��c~�2��,̈́�آV�0'6 ��Z>?7���yU^fͥ��m,&1�̡����:Na}`%���i֭�ySDX������v����_g���D�6���v�*��]t�����ۺuj�\�I��h�3��V��16\`�!�\mRv,������vg(m�,�a��ݥ(B�W��l���K��M��S��z7]t����\Y�a��,ج���:V��T��86��]�d�ZC[�К]�jZ���K�uŉ	t&ZG8�4n�4m&14U��гk怀R 3���1����g<�<��ǩ���W��:QO�W��zOn#���,��M�)yp2�jQ�cR���(�zF���x�Q����V�G��;�M&{&e!�lŭN���v�X�Wl�h!9�̆��ٷ���8�Zڎ[t�G���y���i�ͫL�·�����*t0ҶT�Jv�W]*�!��}\<���@v
F��!�2h�����蓧)�^T9ݹ:^k�!��x�]n��$�θ6�R��	¦rcN�8�z ]�f��&���j�cI�ݛ�.txX$G����܀!��m��!͓!��n�k�[6+zXI����`6�[�"�v7��Ѯ���ng�q�}�/8�87�G8^�\��\Ѽq�ŗ��m&��+����=���sj��˛kk/�G���/3�����Z.�n-�:�]1,@Bna��--��L��:�xv­\�G�|=Iѵ�
�9㓳���dk�pF�g����mQ,f[��/�����0�<s���,=�k�G��ЋjcF�[Ma
�[VbK�Ie���� �yxxm�e^]�[���u��s>�Nc������=�c�0%��P�	�؀`U_����hT!̬IV4/d�y���t������3n���;�U2GB'3Ӈˆ�)�ߙ���40��0G�0a� ��9zq�q��z�Y�Q�r�R�F�ʹ�U'�����ϭ��h���l�3ɛ심��B�羅����&����+�]{5�w����W	l��̶�BW�y�(Z��X��Sq�UĦ2s�&w��E�r�,{Ċls7�5J�Rձ�9�����+ t�H�� �M���˓�3�H��@ c�+:&��څ[��A"j���m&msA�V(�g"K��:TWuݼ\s����:|\�d��j���������tj���`P�E����`hw7j�k��On��1�_���!_aL��vvϛT�gՂ��ܬJ��Ѽ�殷j��s5q���س*�Lx�A)�M�D�Ħ1M�����Z9�7�r�O.oZ�)Լ��V_��
���x����&����=̻�N�f�ʚ.O��X�讛�O]��:H��H� ��զ�����]�uճ����������I`��`� 7��C�5��y�u��h� [2R�-�6$��遾�Υ]�2N7E.X=�;:M[3�]$�
�����]/35���Q�b&`�|�t����X`��9{-��mw07sz�S��]]�N���W���z�J�_�G��y�횸Ɠ�ʟv�\��V&7tzȯf��n7O .m@P�<!�E�������~�����U�<>�wc��o`���W�5�^�xh�؃1�ڻ�^�l��<����n{�0�l�I�®��������5Ψy��f�VϺ�7�C䤛��R��7��g.ʧ V%��۹ٯ���cD�ǃ�6����öC����,�憁��C�Mm�;�vk�.ޒ�Y �J��w]eΚ�1�����{%�q�7\�4���'�~����W�֒��>�;N̬!��Q��S:,�~Z�&%����cɝt�[�D{������;���)it��j��]�	�p=Y����a]խ���
r��.koԙ���YuZP�Vz�����{�t)`�L$!�q�H�k��)�������G���PU���+VQ8A�F��������n�����)�q�9����#-�cځ��~�����g�GɥJ��zi35��'s��|A4|�9~�;`r���N��p�(E�`Ap�yM�̊Y�\�C+��Ӕ��Z*g�� :�0/�����kcsS|qgq��yh�E7��+�Ȼw��+��r��� g0D���e�ճBA(??z\���ˆ:fW�V�+f�-���*�Hge�k�uD֜6M�ٜ8y�E䏋��#�N�������Ee��ؤ6m�w���n4�W�B9��S'=��C=Lf��vz*��+-=3�G:ԗ;] Π�5B�21N��ٹwض���@��*���AJ;y��}�-ކL���7-�{��"�Psun��uo�9䖧Ǭfk�+��۟I�r�JFČ=Y^����Et'�.h8���B�����͡��r�ӓ���]�7��H^�*��nc�v��%m���X`�h�P��//1��~��{'���0�{I�L)妶w�BKJp�4`�M��7&��e:�t���7�O����Y�b�;�-E�[��W��ͦ��!�Ma,q�Dtc1c�!��>������d�d�`L-��_�I�CZJ0|�$��N�@dvL�n���J��f^<t��"�-��*�Y��8(���}�jv�Lk�s<<R�^|���0n;���W��������x��/t�sU(���<:י�u�G7x�)���I�c]��]{�ʙ���1�q-I���Ңݸ�U�X�����\U�������\�Ǎ�ʞX1�s��~띍����ed�[}�~���a�G(.�6D�צC�<�9'=P���*y`�dwEu_q^�Jm�Mz������n`��7�u��h����["gK��҂��ل���8P9�T�7������ƕ�A�W/�D�i�w���2�5!eڜ��ݠ�%�u��L
C��	eM�Cg�˰�QJ۶ڦ�ry݊��A� ��K��Z����9���اI��%�����%���*F�H+-�1�n��Sg���s�:9�J�v���q�����σ�����}�&⣩M���p��LncXmb4�H^��p�Ë@\�c&u@�Ii��F�5,��Ox����R���dϏ
fiu�f���AUK�bsۻ�2dј��M{!l�̸��ʭ����y�Y�/@��.h�`��"�4Mϸs�C��� j�3'��9��U������,�K�\�η]�a6 ��
��+�c��;
�E��Y��*��ʙ�_{K=��B�P��mAlu3�[i�;1��'M�\��!,����A���wz�J�w�=�3�N��Փ]�
�-m�WܧG^*UMA�ͨ���yV���èB��m6JaX$Eչug��z�$;{���N���a����m+������G k8����V��3W�|Da.�3`�[[�Wp1И)�%0lI���;V���a�/��L��`�𜎜nc�4��Y}~�o�T�@b#��Ջ�r����9��/����i�y��ɴ@P���p�f�ל������,	��u\M!�(P���b=�������J�no���@=�[S�c��@jQ}9S[�~%l@pKb0�b�-mը^0R�5��t�o����#`=U�w�Q��t���Vf�S�u��k�qC6�E*�G=��,F1~�=��^���/+����v�j����lT��GH��-egnPO�h@����+18�>�N��Gq8Ge�{�Jb�6:�CA%�rH��̪�t�dpW���g0w˘�́�IT2��Yf���[�����Pa3��s�������p�H��J~{����)8�d�lv�)��.ɞ�I��˚o����]��wS<�&t
���QCO�AҎ���B�n�c5����\�WAZ��Ǡ����}����	�����u�1�縆R7oR���b)�ۗo���Ng�B�'��/�� :_ı�G�䳹ɋ�k��u�����j�~��2�S��M��.'���2snnA�y��W'1Kw^�Gi�d������{Ɛ��ʣ>�7��L�-�����,��zL�yY��5j���J��m�{Ǯf�E�.��j�T��p�q��9�����T�96��Rב��-���Ȟd�+��4Wg�D�l������-	����}~ơc%!-�z_��8%V��T�����*�3񜻸:�F�%��V�9�]���y5��f�\�5�B��or�i�g@�eivy�׀h�[���г2�y�q˻]��d݋,�Zb�+6����^��fm(l�vZ>��uz%֞�(��+�t��n�j��˛=w^�$��B��|��~c��A�1]KoP�]��'o�=��M�b,����NS��]�q�<8��D����ɠ��N�5qݙF��%� ��0�d������l���p���ѕ`'�+�h��P�:���N��L��a���J~��;v����+yy���#<U�:ڑ��F�H�D )3�ʀ��ޚ����%�D���HP�:��ى�s�uv�OJh�:��f�Ш �x����{�=�)���IVB�j�M�r^����p!�m0�"�=��&ǽv�U�s-����=Q�M ��*�z�{s��.�Ml�;ت��y�qOU�A��8='(ɭ�����v��L��A�
Cݔ�U�z'�� '���e>�ч0�V�`�gW��Wq���SQi�L���Ĩ�5�ؕ!Vl�9��}�^������˽J������������D��f�;��)�?k҂�z����t,U���|��]������%�{�v0�����z.����  H(0�;��~�L��W�M.���3�&��Y�s�{ۛ dھ�>�,��NQ�o��<]nf��8	��R8�h3�G(^��xy�Jd�h�k_boz�iD����?7��g*�̙����@���^�r�\Z<�����z)�Jj��[3mPѪr������jJ��w�,�BS1	4-��v���-���p��"w~�}:2�կ�
�y4n���'Z�3��$���π����Ȑ1�Ʀo�py���xoV�1~�eG�>�~jR}Oڒ�XF��
γ���ۦ�/4�aG~a8VF�-VRV����/|y���Hr{�{}�+�w�Y>V7Pp�a�'tk��l�na��s��0��M+�*�xH���H�Rd��2���yi�1�=;�'�Q���{9���ݐ�u�u�t�Zk��C��A��2~��H�Aܪy^x��Tb���9U��.�5�@��ǣ��kt���)<��?F����N{��R�����e�t���S���a�>��0��m��Y��.U��P���!��Pċ1U�F?
u]~}T0We�z�\�#��t������F�M	��
�ȩ��vɅ����Ū��>�9��A�f<Gd�Qʬ��HۆE�9}���l�=�0n1�^���G�O���۽	$�beŢzyu�����}�H$�r��їɿR�R���vu�3F6��OR���Z���T7�3��t�M�_S�xٔ^�9/su����2Q%��F�-�<������]�v��#w�U�����T��ۍq	�4y=h[�b�\�Ώ��!�XUJ��m>���أ�{�X��q�(C�^�rV�	���L�Mi�f�M)R����,����K�3\
\�)����<,uD���y�zy��!����(�q�vN`�^u�-{nф8���Ɖk�rK�h�K���v���̲.t�V����>y���A�Y�Gpg��ay�[��a��sJ5Yy2l�y���zqq��۶��PnC��%�������˷-�U�n����;��욷�蚟��^fH����[F�y;���T2����:8���羸́ͥ
�<H��o���fѼ���Ɏ8M]���zM�뱄�~D��l��7��JT҃�e�co*T���ѳ�CI�A�ސ�+�%���=͂�j�л��`��w3w+e^O���>�<k�u\�D�>0�@-��t<oK�\����㗂-�{v�T�љ�b��[��߻g`�B���2�s3[��=�sw�������y��5���
�9,��X�\}��	2�Od�9��_��y�v��ER�V(|� �^�P{���ΜF�6�mL��\� ȫ\�V�m_rː���ȲI��X���
AlZeAp�:����&���^5/=�O�H��N�Y���{f��XOA���Q�Ġ�+=-� ��n;=�}��ލE�m6�R�h:��'Dy��%H�]���$��Mɧ8 '�wS'�)�#�J����k�fr��W�}u�(p�3L�7$��21�t{��]n�qA�����I�ȣR�9l\�]�YH�mJ�W�7'��[G�S���Y���V{�5�=c���l��ػ$���4W��p��y³w<o���7S��`�<y*Ȑ㚂ۗ�;4�&c`�yn׺*U��x�т�T�%�S�B�|k��nt�ڬ���f��meI�7���D&�4��{�zGD�K^Ä�]_�
ۀq�f�����\s�8魳�k�A�;P^\v�i���j�pa������K��4չ<c�~�;ז��0�j�L����d�SÃ�`c�پ�Vo�u��G�LBh�!%c��`_J�n+M,�#*���kgҤ�e9B��p)���^�*��pv%�OD�	̲��ުyz�s��]6�0�LM!w�º�d�ɪHX+}��n]��p�܋�L�B������~ɋ�^ҷnj�QT��g���ݸ�u1z�i�@�ӽ]�S�R"����	%%��Y�MdR>���_.����ݾ�'/���ys��X�и����w^���_o ���wOi�s�@h�Zdݳ;���=��yX��a*�P��4넦U��^�O3�h�mn��<M�-7=��x�E�NɄÉȓ��]0�j�F5s�T�D����C��AX
�cJ�yS.��Q����:�����P��4�(eB��5*F˩��	)dΉ-�t�f0���g=��<�[em�Qy9�<p0��/c��R%��>{o||v]Vf�vd���f7�^��=�7n��Uړ�n���m�.]�f~�\��oT�y�:c�+�)���h�׃��%�����d����?c��cSa)'�%KV����̓VЪ:3�4�s�e��d\u�e9�ȑ#�j����2��ւ��V�wQ�N���35���Em,{~�;�HkIi��@�C�k�1=�9�/'���ĘX�fY�OE�:�g&��8L�:�Bzݧ~��f&�T9�w{Jܧ��+�&��&��M�]\���~ $�%¹�rI$�;�pQ�´�M0	���{�=Wol�)��8 2�H.^ͬ�3iz(�@����7�{��ռ7�ǎ��=� tR"��� `��o�y�n^����ZxUa���@�O�ɖ/Ћ>և�X���W�?.�v:�\mGL��Q�����5���p3yx�uٟ{�:��P�%�3恴��w���	��G��O�f��.��$��B��֧,q\���iCRyv�{[vɊ��O�N��3���)�z]�7�a�4!��
��Q�.�`[쩺Y��cY�o'Aܡ��lh�fK��3j�j
����	���x�{3����t�� �mѺ�O�nP�#�r�!�i{��>���)A��N�R�_��np��N�=�0laji����O°�Ѹ�Z�"�nG��RU4=�����-�����j�(�q'{k�U̕L���g۝�	���N�Us͡�9u�J�F���S�m�i��[B����ҽD�6{�v#�2�7�9���'��g	{��ټ�[�q���~���h�k;�dm��Z��*��ӑc!b6��f�f(�q%�'�uW+�s+_adQ���Q�q�|"v�vd�x�x=6eb�����P�}�Ƙt����y�`~Y�S�/���<�ی���.x�V�J�]�xǞGċ8���e{gtl>����oS໱,^��w�)�g,V����L�s��`g+Y��l���S�L��o�@��G�z�"�1˟�iD����̹���n�%P�/)t��1�o�����k�ۭEu����Z��=��[.1p���L�MP���d̼h�H����Wsi����罏9��M���x������_rޖ�r�����7���Ҡ��s��`s�A��)	{Ӫ���)��N �
�hgl��9��V�gJ`��:v����̊K�����%���Gt�uPςO/%��W$�����M�\�m�z�[-_���;M8F�l;S�~'Q���vS�Vn�����"��k˞~RM�2�'�?�ͻ�T��t�ԛOx�y��%u�׵���n�Vgs��ZNQ�{\�6��[q����Ƴ�u��8ks�����;y���y��Jfl뱄m�[��٩����]|�Y*�������A�hгmW=����d@Ն�P�����&y�k�	#Õ�*���_Lk�>�7l�G{�A�l�w|��8�6IH� ��b�^�;O��A��dƉ�"{5g�h�W�+����Wpz����v0�T�OQ��n�yjφC e���G�l6S�!Ade��1��<�����b��N��>��4=��
&�.��Ȫ���ݝR /���4#5潺O�I&���O7��a�,��q2�X}�٩�-�����|�}�����������D�>���s�7F�N��Šc"��Z^�s˯0�P`ÂXD�����z&��5�,�½�T��{4���[����Q���V��1G�5�Qy9�f��h��!,aeP���5�	ɶ,
5��/�t�""@���o1㋢�nO��U]��\��g�]�:2���ə�]�F/ �cc@A�M2�&� :s�ü:���sv'`\�)��]\/ziHW��'3/H�E�J��ގ��1BA��3����._~`����T9�;g>�w���wXm�چS@%GA,\����ղ�\'�@�sˤ���Vn�����"�O�JI��{ӒK��;�,N؜���5\߫-��$��+�\�L��C0��X�q�e�oV<�~��1��J�M�*c�c_���l�.�b3�Ʊ�rR#SH����ے�	w6�k�uf /k�˸N�R+7&����׉Z��^��v3XZGj�l�%�6�!Iai61�yx#5�(^A�qV��m�,R7���-�b]���[&̀��qۃ��7Q���{)�9k��"��TE��b�f��͠F�ι	zc�ae�ܽ8��0  �B!{�w�O�~�c��b�q��T�S%s���fZ�R���^�m�6�PZBǍJ�[��5�
6c᳾�u�)��Ӳ�z���uh4���K���ъ��	^~̣ꜵ�=��i�h�U�C�����ޠhƀ�dtքt���9��P�>�|����{s�	�Yq��R�F�����AΘՌ^i�4�_p� �pT4!�Ը�wY�>��&�ߌ�9�j��w�
�NO�}�����;��JØs����Y�ĲRsE�(]����rq{�y^&Ub��W[,�`@����a��5Puy�j0�ڬ�����UVg�i׀��D�=��3On��6�Je�,����Nd�5��fĩ`eM�wU���s�����<�(���*Z�]���xz���n��x ��MR�8'Dni�Ց�P��*���1s�m�E������cL��ڬ�{n;��<�Eo/����1��Y��4�H~���;�p�y��ؽʺc(�Q/D\��:kp���	';�t�`ǔv��%P�e5�Ӽ��XN�v_��
�&gd�M����<���*_�eo��{>���p� �6���?WD��=ݕ��b����NN�Dk)����l��G5X����=�L�I��`��M��q`#2�х��Gu�k��ܸY��:}���7��"���;��Y8�'�X��m佥��p��
���鈪H�E%�p!n����RE�Gm�.V�M�R,��c�N��C�߽ދ/�pm<Ǩ��+���#��*#�P>�(4�f�G�����1k��d�#"ǱhE�I�4��,0���+9���6y����;�U��|���ދ�{����G��3�v�H�7����W��}l���Kda��޾O�[Y��oyLO7�Ŋ��g9�0e�X��:r�%X�	���U�ѵ4k�X��b����r��y+O���Y�{���
yWL�����2ƅЃ�ED��������X6<�%��Mڬ�1��F���1�	���� �wu��fR��9 68Oa`h�����{xk#��#l���q�3T��U�Ng��ȼx*�&V��r^U�!�^7���5z�����\���ˌ��M/LL��<�qm*��L����()Мnǩ����B@�	ąj�-�*Z����.���lW����%�A2�o�-�tl�E%MUV�c�����[)�0ǥ�����_{}�P)sɪ��D>\x���������	�m�DOo����n���@K#��[P ��O�>drp/.�Z�/Z#Y�3�4<��?yFD��x����0��M��%د==��������m�qL'Zә9RI��Q�nN������D�h)��=[
��yl�X�Ӑ-ںRn�3�V�aЂ/��B�t��a��a��i��'D���f�1�&*�z܊�oMi���ߐ�%��;��f��͡V3g�o/����7��Tu�}�7��A3�gM�.3ԥ�lN��l1��ˠ�3 �לp/K��o,xmY�Y^8}�j�i-X��o�#=���̔e6�z���<�C�%_����y����.\�H�M�^W|�����,ڜs�&M��7�gu��DǞ����Pz�_D����_�'m�F�/�m�f����*�IM�=�����`���<(��ư2���a�����o2�6*�
�3k.��ь&X�M]��������~��W*�&��X��f=�0'	v�Hfc]<�G��ײqJY��nz�n�݇	��4a'�O�E�����
���c�wdn�8��NF�y�x���r:��S�S�<����G��~9�:Ӛܽ�3�GB	�`"��;����nO,����^9�sn���܋�Y�t��O�E�zu���᩹��w(�;�$S��ٷ��Skmn���0g��/�1hA1��=7<lp��\�`��z]�`Ws�˖`�oE�w�='�51"����O��eb���SQ�7@e�	lC[��Tp^NzLr^ �G����i�o7}Y���`���֕h{Mx�5�iv0�W�&����-�c�w)m�0�J0Sb�'}w66�5�go+v�I��#<�4�;3<�؟kt�ɠf�Z���~^4l˰��U����K�xHY�,����}�#u�6O�X<ܳ�Ϫ�͑O�B5���b����LT�Ù�"���,&���fŞ:����ہ�=����+��ٯ�7��X.���[�BwT;�YOXwoL��+o��^w�.���گd�h@ƴ[ ��a>��ɾ��ܳ�n�?<�����l9ga��o���.��zR�U��=áU�;����p�QY���fI�۝2�s758!�_� ��.��c�h+�%���U�.�u�uߍ�[.�1�.�wrފ[�g1A��Z��T�p/aѓ���g��x���#�\}��.���N��l�a��mA.�Z������έӵ�%�Y{��֌�
����I;��4�3fn^��M�6*���gzK"nu4�<�&��Q�N����W�J�2�^̠,d�&�w���	+����6\n����? Yd�+N1�z��Ʋ��4 ���t��G`��/��&M3��Ƥ�ok�8X4������Ih����&u�����r�qveT�@�6�nk���� �Ṗ�;��u��_��n�\l��=6法���y�O$��Gnw�p�Y�uk7&���ȐVlL����5�i����m:�g\`v;����I�p[�	���vf��2y�:�aϴ^Cw��v//�����^-Ծ%��L0Ϙ�q��w�+*�C�4��v�N��P�,����r�U���/���4'�>�v�7,z7=7k�V5A��l틳5�	Z��$X�&��P�:��˝5ى��z�y�~?����VoG�&,-�%Y�e�]\�-���4�B#�����6.uw;}����f](=��P�q���#��c�M�2j����@*����o+ I��/F�k����܍Kb��R�ZF��g#�KO�)i��co�{b�W�����a���{�w�gj��^Ɂ�#����wR*�;Xdn�/O���	���M:��sO�omݻ^k�b���غ`�b�aak�J�8z�����-�~���� �͡k�V��^��x��`//ԕּ�-xD�� �?��<+ixQ���",����{C�/����P��j������L'gt,t�V��~+f$l{�P�<�^�kӫ(xY��	����*�IO'�[���fcd��^��^���8�$�R�沩��[�Ih��4��������1jc�vn�\9�܈9���e]?�)=�Ko�����>v�\,���tQ�g�!�;����#3)6�6 �[�.Uኯj�b����gv'7w`��Am�R�hB��]zP��0/F��Y>|���z���V+tͣz�G$E����̳�a� G'�4�,� B2L(_��+Nf��]"��~g���FpEJƎ%[ݵ7���YeV��{���z�^ǷX6�e%	���}��!xdŪ
(�-g����욘7���[��q{.��Y��a�00
�����2��� 8]�ʣ,df���C�hf)�w^@����=��\65��|�T���ʪG4�pkJ��9`畃�F���v�̹Z��sݜ�B Z�	h~�>����(���g��N<��^gl��v�l`5[TL�t�� #�Uk۸�;�m5�&v�L׍�u�w�_p�Ǯ�Ø=&�U������I�TD�������c��I�����l3��{��N�y!X:���g�����:�c	����_^wy4d���h��gA���/����h�[$��*�=��T���^^T�'���㼨ӓ&� �Qm�S�IQ�YO2�ٽ`u�9^�c��u�k��\�-�O_>{���K�^բ�z����X��c��M�\ԃBHl���Ԣ���2ۄ/� _� <b�b����E��
kDkEbt@i����!���]	M�Zw��Ws=���(�]�Y�p�+��L=���ln��Yi%�z�'�`��*89u�C/��s^����t�	��ʈ����3����r�`ʐ��r��p]�K@�^�B�E쇫}]��D�X����f�Q�w���sӉ6�d�@�<V]��U�=<� y�uo�]Z���is��o�0���^(�i������ӈ[CCxz��٧��,%�G��x�W��u�\K����ٝba��<28{:��>���K�.��gK��pa��[��5�C@�d*�.nkws�J��,�����ܣ�����<��}k��vq�g�{+�8�z�j➉����iW�k�%v-6�����鮻Y� �c��� ,C.2
��4ƃ��=L!�y۝�eA4wW�����	���@�6��m�W^���������-�%��p\<q{ &J�=��2��b�営|����r�.jpcܯS�0Lώ�46( s2�x��@�P�\�̝��ja^�w]�ֽ��]�M����gD�9�Q+m�½�ܳ�~��M��>cv�ֽZ��9�p�5��O]z\6[�2ԁ'S�^̔��鯢#I�J��隢[�r]N�[�O;�����\��[Wd<�& I����nlxY��]:;�����-yA���~cG��)�o�!�l�Y��+PCK���z�{�ݏ*Y�'_&]�N����;������$��� (���c��>�{wz���&p���;�"3ƻ=Ԗ��$ͬ�5���^^���;��zr7�^�ج��M���z���,�[�o�gx�X���t�
� ��D񽵘����~
�@P^$@{4�W�X�r�� E�]^�%� �#dԷs��!�y{�#	4�85xC��6�#���e�[LS�����OA�M�1�<;[U��Ks�2�0�<N6���ϛ�H���@2Tk'o۹SGۉؔ�-�C��7�7݉݁٫��G�_P�wA�[1��U��46�z�6��VA�&��d"4X�:N_�r�,��BbK�/�U״�]��^E�n��ł��nE�s>�z@�X��z|n��F�d8%�k٥ԗs�f�im�����2�9���"�])��K�$���ul�7K�bН�u�o�]?l� 	8���;�E��� /ͤo O`PVB�Hqq�=߅�Y�=�Fj��I)3�<�=x����ob��Ў�^�vQ�R1�BJ�����x	�<ʊ�W���b�cdݲB8阛p�:|=���
]�\�d
�[0C�_dy��A���q�]�p�c.�����;k!�H1�DɃ��v�q�N1��Z�� ������	��ϭX��S�\np���`��{@Nv�rŚMv���zz�[�ږC�P8�$`�+�ϣ�A�s��ݣ�@Md-t�
�Mzƙ�],ұ��FENTv��p���۱̬U=��w>�$�@|x	�y�=���<x
r��m��j�kU��;�{�]	/��������hs���5��K�;8�j�,�q�?jZZ[����+P�M����p�*�+݁c�!��냛-���Vک�~ǥ��- "u��;�M�t�M�ŷ�U%�o��xw���T�\���A&w\V����(�n8m������I����BN�/nm[g�J"�$rbe�a���cͳ��܃>�;�&|p�76��CA�^��xckxg�u
�ai&L�
�[�P"�{��疉L��57Y�b��A��~��4,����l=�)��;���N[��2/�wU)��"�TmYG�$]��M;y���o���.��7�\����-
o4��5P��ѓ�#4����ӻ9��yܬt�=���6��U�}� f�NL�(Q����f9�jݚv6�����1�jR�m�Z)��������u�u^�DP۵S��M�+�̹�T��`�)�"
a��A��Y��)�[��K"Sf�3"ױ d��;;u����a�i���q?
�������h�oTB�ԩ�W�ԕ|�7��� ��Nݭס����(����TW-3��-B^����~��^���H̾9z{��rcq��0�a���r��FA����g����Xް?wm�T��٭lYJ�a�{�������\���1R���ܣ�[�Af{k�B�T���g�9�Ļ�7<��̸)X1���$�;��s:[ˑFs=p��x[���u�|��s�$L�^��}���cʈ�g��<{�/���^�F/�6������r�^>}�vǯ�Z�.��}�O{Qt���Ӈ�����μt��W�]����wJ�p���H݈@�9�feuv�99^��a.ʥ^���>�Fe��լ~�����X(������w���E\,�s�h��j�y���εʎ��$��G:�8�S6{�x�r�}��V�r�p��;R,r�)���T�[9d���Yۭ�iH(������U��������S�4>ѵ�M��>r��6u�'wԉ��V�s��w�̣��ޅz	s�r�_SF7���D:�t6����e����[{:��hQY �hF��	to:�ǫa�|�'���o1lU��\^N���*��D�Gy���s­Ae�2p(��[G�y����ғsFv��<ݹׅ7��'�ɛ�1�I;7`E�훼�[y�������ލ����&��b
�G����x�#h��@�Uىj��[���%n�cR[T.�q�
C�6��z$$�ň.��H�f����x,�<h�*�E6#	��#pBP��GvưE�W5�(��������av��<۰�I�\]vLt����kbXA,h#�Z��R�����[��/��I�أ�'c&	 ]r]�x���H�:D�ap�SC8�c�Kz�fR�H�r�逪�lд�65�]�I�L4(@�ϟo5ֳt�[�q��1`�Na��%I��R�zcFcLd��CGf؆�j����h��h�W*�Y���)���A�lO��brˮ�g\V��Z��̍�,�!L��\i].�A��^��9���k/�F�]�ns�v�<�9u�ظ�iY�lx�m�f�*�`�F�l-�1Čvns��;����cգ̩X�m��PN�=/1����5����3�\��]��C�qu�
��<�v
�d.w�+/�TWV�FC�e����ڍ�#c-ڮ�T)h��[��ۛ9������H½��pu��Ev�C9��M�x�ۙ:y�l;����i�B�����ah�k\�+��f+�]k������f�&�'EF��b��գ6�N<�-圽a��yt�;&��{���2e8�;�s�!5ۛ���Ԭ]���&,����l��v�p˜�q���Ӽ�hWðR6-Д�$q������n��A���dL�whK��lA��u�*APM�䖁��e���mdoC��;:�8:�����K�#+Ad�U�x
9c���e!]�2l���$6/6�6.�r����gqs��r[���q����Վ�3����C�|L��/lK�qι�㎧m;�籗 vg)��r���K�.Mq�#�����m�ܼ������ym��0����']���ݮ� :y8-q�h'�����I͖W6-��	f���fS��ݩ���F��ێp�\[�r+��ȍ�vzY��M�6;Ggc=lMW�Ś�.�{lۓ�+��N#�<g�آص���Y#s�Nb�,�NYn��^�r����(���rj�;OͿ^���v�Vƍ�p	.A\Q�)20��U.W�2F�h1*��[ژM��'#pĕ���:rG�r��:�S`�^����8���1� �Az�;��5� �^��>���������&���fݡ�ݷ��h�m�f��UĀ��BD�X-�j��,[
f�'�sLI�R(6�;���i�ʦ:u�[D��3�x �Iʔ�ݜ��m���	^z.�uT�N�i� �@k�U�
��L���p�Fv̞����g��� ��[RskQZ�<�����Z	�=0�����j6\��Cb}���kf��FVӶd�R�(`�>~���Z�c-<�ė8$硰�MϳrhD:L��ߖ���S�x
#76��y�zKn H4�,������E9������\��ҭ�9���J]F�;�C5P��"umTw��ڇ�������F�7�Z]6� N�Ӧ��0��Å0ж�u$ת��9�����3���ҷ��� ��!4�m��v:��A���V�g��c���r�ј̳�!H��iR�Ѕ�;F�*}��ǁq0j�k�o5֠d�>Gj$��{iv]��
Z|�Fk�E��@<����o%���XC��������$�·�9��+Y/<�I{5�7F�	�Y,kM���`�d��LgOM7��nx;�x+�Ԍ�|�.�P#�Y#@�Vŭ����^��ļ[$�/d��Y��M�0	-���*-�^�d]�+�_^#ُq���׋kr�zb9;c�!��4��Z��S�P�J`��tp\��M:���m����΀ecv(❺�y�0���(1w��N�E!��ҿl��%״;V�
��g�ģ00#H���WlGT������(-4�,��� �8GO{{_W��Z�,ox��%�u�{w-^WXw��y��.���:��}R�T��G�ûi��c��B��^Vu"�!�l���G���&�"L�bՌ�
'u�m
4���,��n�0e�f�p�Ң�f�R�v���+���Z���K�����W��T�埼c�eA��n��W����^����.�.�W5o�|����SHh�1F��&lûB�x�꼩,�hk�4��[4�J�&�5d÷�*{wsur�/of�o6����ɽ2E�}���jgd�~��,�i2R$�b�q�P�m��Q����%�Y�䁡�bM��U�[VDxms��֮l������&�	˝�#�G�򞧈�:�"�kp����Sk�a��l�d 6����?2��<�W�! [�����5J���

�cf(=3�Pɥ^u8�љ���`�o�|�d�4ĥ�D��*� 93�ٟS��[ F^������v��@$y~��z3��[�둞IX֍X��Z���{�Hm� �������cg|��J��)��y���}[�U��Ŵ�W��VGfbʹ3��w�¨�Z��I�eA�J�gn��sq�� v �ۆ�i�j�)jn��MjU�9�Tm�n䌡姞�>����t��\�K�Y��4�5�A�*Z�5�n�a�0�bA� �MV��ͻ�"��<8qO��潘�=՝H�iʭ:���/D���S�ngS9��k	�6���t˔8{�v���b�V��͒�3�uݫې
�W���X��Ce�A��mmI&���;�q�Ua��8��8	&��YǮ%g�rJd��s��x5��ۻ��CI����H1�[E�/�e��yY����a��q���1>;�6t��S~�˃Ks5
�-�a"\:��^��g0�2AGO��f���6����W�d)���ޑ~����^G1�Ρ�8�kΡ��\v�C�8�L�B����zf�}\��7v���2��Ĺ����eh��.�i�5�\�tƘ���\9�8��LNx��>��|�%��d۱�<z9���pq����:��K�=H�i��5km���l+,��h��,�-&IBtRS�b�Ku̤�2�V����S��Op�ƚ������-�G�.GM�iO�+/����Wvn|�����r��+�
�w9��ny���������0ub�T�1�ٻ��=ߞ�T�잿���ے�E,c�(Rl��W@P�5�p�#P�'>�2�t����F�!R}��d�{r��gL�g��Od�������8�.yMc}��l�<�{	=��L�vqޝ͙8���2T��5[�tU�x/:3���k�%�� ��A�f�m�6�N�b�\c\� X�����������zgh��X���6G�̟2����1�!�A�B<��[�["�;Bc��v�"��0���q����^Y�u�Z�i���g����.�WY5s��EfF` 	�L�@��B�Ҹ��N���)b�Ӵ����x�n�ms���d�xٙ
[8<���{�Suuў^	4����x����Ԕٖ�q��v�6��B9.d�o��*s�h˜5�M�y˛����G�.�Y�c
<�p|l��I���z���>z�ub7G	�*%������Vf����a�T7%:%��E__��?�Kc�V�H�#,k<9#�8�\���:�-i��}���gXݹ�rԾ���Α����F�t�n�غ�%��*��L����4i���	)�^�Oc�Fat���m�����`�������8��B	pQh/���2ו�Ǩ��.{s��
�(+��۠�孔�bo�BP��uBjd-]��*.f���k�	}�Z�	�os�ʴ@x��X�0`@�`�S3���s����d�����>���\�ǻ�K��wk���Xx�1\�B���͙8�4GyM�����7[���r�{Q��y��4ح���t9��o1����Q�Qq��U�$��V�2�,�+Y���9s�k����A����P�)Ee�y�)X�u]��q�'��ed���� �xȣ1��B��;t�j,��A�8��8������^�$�d�x�cKe�<v�˽�{��}i~ˮv��2��R0m�=$nx홎��G.y0"��k1qZ�T_�~���{��²Nlg P�w֘����3��[��'�ak�7���e�Խ�z�������:�u�$ ��������)�M��L�P8l�e���3�,��6�(�rr�S����J����I�� a4H�O{kqYC�	��-��L�E���K5�Y�ͫΡ.�)���)��9 �Z�Sv�*WXf�ef\��=��ي�;vO�;���c�����U�����޿v��5����*<�70�n����8�W]�9v*�����ǒLA(�qЫubY�h��;\�NZ⻣�uГzE��;Y}6=�c�@���Pu?�� �j�'W�V��O֭m�����f	to-aqJ�`�޲���q�Úpl˟��MBK�B^�r����ρ*�l�XD�?(�US�-GD��jk�ڻ�
��Q�h+ ��k6�6[�m�V{��[Ԃ������a��X��{��^��A��?X��]�^DCN�K�Qz����������	�i�Na�&'�]��N�yѥx��3�s8gU��73;��Eoŷ��m��5�Q;�����ě<FfQ������d���s�8ٹͨ�}�N�p��QR�Ă���$�r�[[�9]�1�[�T�Į�4��T����E!@��jͽ���cD��G��ޣ�̜py�^n�۩�����-�v�d���be$_��/�UA�O/o'�]�e+u�2�j��n�7�g��3�{�7�1B�j�������͢��,*d�~��ȴG=ۢ+�a�p�����՞�0bΤ�fr��:��ۚq�����=X��r�w�9c�c ���4�U�T�)y/8����gׯ�l@�6[a����VXݨL:Zg�� ���h<I��ŉ�"����\�}����vD����>�3� F��^ë��I;��{Ǽ�mac0���1ݗ=�f��+�7#^-��M8Q�;�,L������[���a��\�b��PmAd�ʟy�N���r�	I���)��Vp��{�����ٌL�]H�����+��F���Kr)Ǳ����)4�e nR��W4���8>�ti����`w
���j3�b��=&��� ��kp)V�;7����"@�㭪P��;i��+��=~sZY겊5�jG�#���/���٣(K5"�R]4���M�Q���x����z�+��ûO۝��jgZfFRa�X�oZ.�M�l�L�cZ#����L)9��\`u�f���TƘpk�e�`=u�Rk-�Ϲ1ޏol��'<��G�A��<Vm���;e�RYd�ʐ�%�@��ư��ң��P�sxף�g�T�b����A�C�7g��9��&�b=K��{����>�7}8�Xl�e�#++�|�R��NA�k��3���-���m~T[��k�}u�k�#Q���y�˔E�7�-��W`��^'������G}�}�$��qs��<���N&%�0qa/��9���ٶ�w:3Z��ue·l�PQŪ�2����^�����Vclv�wy;��f�闠��;���u����/8�H&��sk������͆�}7�G�f�/�����e	�����3Q&�[:Y�5�8��E��h��"�a=%�*�;�.����A��k4��y��{��vl1��ؚ���8�b6�������:xw��l�q1��7�ז!.������^=%��𛕊T�%��H>��[z�Z�v3�t��v"�ʳ�A	9��t��seq�Y#ٙpK�b�G3�����鯳�v�o�(�M���ohN�U�{h������]�x���I�-�=T+�KE͂�61��wn�a��f�N���kP�d�Θ	yɚ�(��-�9[}%�9�g�� �"�Iò��7S*A��{>���.�X+\i�*��<ja�	�Ķ��tK6u���6�m*����!rflWŧEa� Y�2q��3'S�ky��]��r�/��e��w��K�.JF_>�cP0�	L�~/Ǔ1v-�����K�fu��*�]nVȲd�d����.��+�%�u :���r�s̋+��|��m�f��U>�g��f��%o2�V���;Sܮ���>�Z���q���L7��8�6c��칃)�V���;D�Ύ�oV��,iui�Ï��h���y�����7qc���#>�X
m6Z��,�V�쵽Ky@�KVs�� ���\���m�b�gp9���C��j%�F~��0����!�׊�zx1���a�0rYv�0x��ttE��|s�}7Y����f���%�BVpe��k,y���-���2Bo�=k1�P�a�0�L���$�	fR�>ذ|��_�
���	��6�vg����lL'�3�EyN�{x�繽�D���9p-���>�������Y[N����oiт8;Ã,X��l�4�ʾ�D���Q�"�mkT���˩4��3���k�o�T���m���w'Q�����xZd�����jz��N'I̛6�����Z��(p�qgu��=��3{:�)�[�wl�M⼤���Ы�]U�F�1�X�0l~g�:57�@o�i��V+w��]h��D�ClvՈ2�̼��d�W=ъ�Ye�A�o���^x����	�5Hg�*��\򐳝�%`K\=Td��p��)嫗���~!��e~��*D�ʼ������=����ڼ�����۸�9 ������iV���5�\o\�4�M@�x^#���/��$PC�	{���5���Q��_��se}1�#c{��<�^�"��q�ه���6={�Z�)6�����~����|B��\U��a����	� ��@�M�m��y��h}z�~N�I'ww�N�I'ww��I$���i�I$���I$�����I$�����I$�����$�ww~����I'ww�N���N�N���Ӥ�;�;��I���'I$����N�I'ww�:I$��׺I$��ǹ�$�N���:I$����t�I;����$�ww���$�N���:I$��׺I$���}�I$�����e5���<#����?���}����*��JW�"BEm�H���)R"@E�A"W�5AU*B^�     =
   @  �@    .�]��N����=�5h��{g�vU������j�aF�޻��c��M��g@�:7c^�� P�   �@   (d   � �� �  ;   ç^B�w@��X�
;�p#wp�U�(�
v�$�"%-s����;x���z�f��r��޷����N�t�{w�����zz(�:ih�Ż���K��j7Ν�Э���  i���pް�G��; �w;��x���u��m�)ס��w��z��Of�K�Kf*"�1o�te�W�Z��v�{t+ԥ=����Ԡ�4��Ѫ���O  �7i)֒�X
�I0!l*��^ڒ�L�^��<���	*�v5P��L�p7wn5�(D�������R���^�T��
�d�Ō@*�   ::Wg\�ݨɆ�1�)M2�I'LO^�*���*��+�U�T(m�X�Ĩ���U]Sl�f�T�e��jt{���n���r�aT,   ;�GX�tjWl���C@w�s3��)��!BU\w4 k��]i�k��    S��)I!&��@  � S���)C �    )AM	��ML��5G�6�mD��=��L���       E?h�*�z� �  � OB�%*P�&����i�~�������#D(T�
�����a���4�D&�[l�9g,�J�/�5�TiEA�S�,����?W�e����|�&d�2�ȥi��!TeVbR��.���V�v�i�8�q��]�֘�ߦ��ű��h�^z����=z:�M{7ק����4���4k���7a*چ�Sa�j���֐��L�Y�-�:x�U�@�����;��x/�u��eWiʎ�po�gL���&�� ����<��::}Y�z��q��;SJ@5����S�|V�˥�,�e��.��s�t�B�m��Jr>���!����N��pCf�۴*��2�@*!���>�����ll�U�����C�b�2�У����r<���ao�]c����`�e��A��MB.9Yt��L���WY�.��L��;W�
���2S�)�a͙4MUP�N�2�^�5.^S*�?�~7$DFvޗ[����X&Y��z^�(�N2�������ՙ�5��[Ŗ0���u��cr��Atv����8��|�J�e�Ē�i���Xd�鍿��حE�j��$����Z
�	����Jo��/��#�̹��	r�e�s�f�$
�ղ�yn�Y7�hj!��e^m�6C5�{o;,^�#/6!��hd������lAI��[-j��]]���W6��,h���s�+�4�mKB*=��Z+)��f��K�ݔ��r�zr�ȬV(ͦh��&�e��ر��ה��÷{�x�+,��OS4���QۡV�dR�e���4�ya-��p�6��a�e;�AcL�Q�4�i�ML����3"��udx�Nz�\���!���*�='U-�5B�|v�LT%+ͽ�5oqj9k�g,f�Å]�R��7�M���HbY�9\LT}4�*㫅��G&i^�&efn��4I��ޣ��<��Y�+��x������Y�k-�%7�R�%�,�L��i��ۖʻW0�%'7"��k�YI���ƴ���x���I�����E)bӻ2$���Y�/^hg��я\J�0�ߏ�]CO-�8E�K5�LX�"��G'�k�u��W�Eu6���gn�&�+(F�Ҷ�!���aR�Q1� R�VT�p*�qU�r�e0m��9r�޳{PͣYv4 �8����j��3d�)���6�㛗�9��[��X7H9�`�r��q��Y[Kj��L�V���(c�Gz�I��2j�1�`Ǩ��^c��]��ij`5k��|�v�U����x��o].�̖6˴�(�Ⰺcs7\-������8��Ki��YƬVf  ���sY�W�P�::5(�Ӛ�jh��q����l��*��x�^éjv���Qɳٺss*	����!r�l�1^	�╏1��ɴ����y�[%k�ǋ�d�(�d�n�'.ܵb�����o�m,��	AA�4�����8h�TkT�Bh��V��������3v�'�R}��C �N���;��<���/��t�{$ :T�����%K̟u�3(k�7�2��Fx���ٮB�2�*�0�g/�:[fkCvIu�Ụ���y�v㥒�z��z�
x�s"�v�ڥq�U�&���ͭ$��F⺇���j�=ui�T�4wvfW1���6�Id�n��[�m���FkA�u�t�;Q
���P�����F;36�`_nǃm^��Vm%�j��*;���x^��mk>�H����`����ƭ@Dv���ǚK.a[	dc�~��r5r��S��ؗ9����*N+QЈۼ9���ZpѺ0�1ņV��[��4��1���x�,�dV�9��MJ�Ű�{ܱ[�����n��H�F�b-P;�\��TP�H]�˩.�n����QH�fջ
2-�kn�"����u��Uu��P��6�%3Bź�V�DV��͎�Lw!-c�S�7�p�S���ۼ�s�re٤&fd�J_@�ë�ݞ�K��M^V={d�	_�I��V,��ވ,]f�/r[R�j��Z6x |��~�_v���=k&������E���Mq�I6�n����+n�Y��>� �����K������i9�M�Z����%�4]eCSƹp�ǽP�G�G��y�)����*9�+��Ǧ,����O�e�ϪA����p�gV|�p����T��wK���[9��|1��꼠v�.��@·P/��}+7���ɀK�c@�2*;>�Y�QQE�y�٨Qu�I�qI�>�P#��F��T�X�0c�[���ˡ�Z��6f]`�@fҷ1�.�ʫgsPI�X&�aWz7aӍT�����Ȁ� ���yB޵x�qЩ6L�/�fe�+e���Mowt7ti��*��}����AGUǈ�W�B��9,�j=��R:���Q���]�s�v�K%�`Q轙X��ٚ��A!�5��E�ԑ4rH�b�5�AYK0մ2G�x��<���d��[A�n��#���vp9Pb{9�78���\U��ł�]��HUh�����1^X��0n�2���`�3�7b У�h�����miӤT;p,S � Kx�U��(nRD�+p\�Ź�A�}d2�kao3m)�Q�-�۠�d�
ۄč�2M?Y�n�g,۽����0�d+�!�bUO�'�a��0�hK�[X�9�p�N�1�@�i���G�&�x��h�m���f�f�-�Ф.>�כ�,cyf��A�Yv"�Uw����~҂�4
!^v�ҵ��t� .���z1�D��<����wr�AmV�ؒ�^4�9�͡��u��VӾͮ���M��̪�Ҽ����|,��ဏ����%�3�1enȗD?L�%Q�N�yrt�^kreG���v慀��3z�I�S4��ڢ�Z\kz~&%�wZ�3������3�W���ECUp��EE*`��VD�\�V�O����~����ϻ��M������UNE�-�R6l����u�kP�\��^�^}�G��9�\b�� r��GEں���X�,r�n�=v��+���`Y6�g�gvNw�f妟٘U���,5JE���y�hr��y�B�G�[6�
���x�؄х�FL�X����\#�x��ۗ!gv�_��tB���=�,m�zn�}Zz��f1S��O\��n匘e!{{���V38ݤg42�c�:Noտm̝�p �۰]1X�!>1}��A�f��q39G.�4��B�42j�}��X�u�Ҹ��Kʨ9aǺ���h�eE�r����c6�#n��rfF�f躖*b���D�V3p��\!i��J�w[���DG2�LYm'(B�Fլ�z��m�p�o㤅{ob����L��vb��~ߣ ����6EX����a/��Ek�L�
N>�<6��\�:�gol7Cd�/@V�K�{����s�š'����X�R��L1�ǯ(eIR�uM�p��t�E�����h��}�U�Aȓ�fK�~Q"� )!;��u��3>r]+��|�1��>�]�"�� 7sgSoB�N!�����JȻ�7Dm֡�
��`���:e�5��/��}��"n�Iٖ	����F�,]E���֪��:����U:�v?�Sx�Nž����2�Xt0v0N�{6���2X��/c@XgĹ�M�M�p�q���ӧU:�6(������Eβ�G�Fb��ѽ�{:+t/�Ѐ������J����}�5�鷓7�䫗Pq�r�̺�R'UZ��b�ɗo`$�!ѻ���5��Ӂ@�5&\iL�r��,�O)�@��e/��^`�L�l-�j�:ch5�6JuC�o�������5j۷#�#�-z�1�σw[�����QI��@�R@Lj""1��n
�PJ��(Mj�W�R�{t�/KUU*�U��anT���<lV��%��UR�0[UUUUUT��HQ�۵��$`�6O;�RZ��%\;��6�����+���T���P ����X(
������j�j����V��U��vvj�OjeL�*ҭu+���kSUJ���ٵUu@հ�(� ���!�:4�W �mcT��9�J1 v�v���quRqs��,�F�@�\�u��`:�A't�&��F��l@U��n���ziG*+G]���x�M�9ΰ;d��	�r�l���.��VM��8��b���!�{�,7<9��n�jw�����u��s�7�����YΚ��{F��m�C>�-ŪAȣ�������n�Tb��̛����q�X�{�q=8֍n#<�)��ƺ��7V�q���ܓ�̔��z`��*ub��v����嬔i�v�¹ss�0ŸnE�3ڡ�{p�툵{�&۪����ю7�w#������T���=�nXȅ����0;k��e�Һ�������x{A�6&���nvD��=u��t��ۄݳ�3��d�Wp-8�m{!&{t��v��5V������[y�s�z�-��,�����8��d4��g�<v%�xuw�Ͷ<vRI^\�n�q=V�8ݚ��=�8[Fw=���)�LvD���c(Hڱ1�a:�#��`��B�X��cGl&��|D�m赭�9�y��:ssmعN�u�_mĩz{#<{n�^6;p�=[d�X�8���P"�1#%���ڎK�]�۩�H�7���1��x6-Mևy:J��էwh�:ə�s�n�лL���s���;���W�ݧ��.qX2D
hZ7mьsmM�{te�n۶{g�a�q��=�L��;��.�׬���mP�;�ō���c� �Ku�:�R\�x�!�U���a�`��\=]��L�����I^�F��A�<�� nQ6	5{�F��m7����p=�ë� �^N۰I�s�^7�.�nw4�Iڗ���C�=�]�۵B;"���;wm�8 6����)f�������{!�s�����n�9���[�i9�q�B��x� ��۶Wv�W+�s��GϕM9��-ӣ�������G�����dܕ+�s%ng͟$��!�d]��Hh=3ф��`�{>���/N\�x��n��
���lH%;�hx���_:���t،�t��Q�`�Xz�҉2;l�s��t�n�eCn�Q*���^ON�s�:��*\�H�*`8�6;nxa�<<���������������(v�6ۮz�
�dq5D�TH�D,@�=���ǻG`�z�@��u3���k�ی��5[�8^gE�grM�]kv�#^�h۰<yy�׌�sС���Q��Z�ݵ���GF���hx�n���m�t�ͺ�yG�X 7��N�َ�lb�ט��w=oa�s�"�z.����!-ݳ�� �;��^�m�ka�1����v��[�y;�==c;/)�p#�9܈z��ê��2�;�@�]���� ���p67<�9�Ń�-c��<On۶z�ݻ�w`�拝O;nzC&^�a-�[e��ceݷ<r�n�Zָ�y.0X���@��6�uBȏ��+��ܝ�Kw��ǃ����Gd�������oi�v�&v��n�ɳcW7Ok���gع��V��^��k5�9wv��5՗�x��ݸ��.W<|^N�'n��S�w\��O=q�N;Al'�!��GU�u�/�5�ܧ��k�Q����K�ctn �����@�\V���{M����{q��yc0
rx��d:����o��̝c-ֻٴ� /C׶���<n�i7��V��=�7V� <0�y{r�l;-�[v��9;Fq����D-g������q���hw"Ww���N5�s�N�@5�^5-�0#���kD.#q�6�n�l�u7:3;rc�����#cvn|�T�(^���bw79��h�/%�Z����ڮA�G#Ԏ�e���k�kv��gslh*��!�SP��hC� 
��lӶ��51՜�����p󺛋����:��e�N����q�s���DErq�S��c�8�|�/��۷`r�a;(���Ws��h���]*e.�|>��5����7%�-��uֈ
ۮj�8��+�ې�v�n<��K��7n����sXײ�uv���mGlu�-v���`�24v����u�@n���s��k�4S����(�֎8Ŵ�r��9Γ�
�u��u��ݵ	Ǟ\GYͷo=ig�ү8��;�nr�٬�rp�^M�vm��������f�d�J��cs�cN��G9KvOEn����&��f�-�n8��k[[�4E9�x�M���s���ʹ�"��iq�;:���n�+��l���;^v.ځ�Ɲ��5�{Bv4�F�C�8�8�7�v��c��t��ٖ[\����cg�;���iz)��En�u�.�n�6�;v�Wgr��ۼV���G���w^�-���F��Q�/WW�����l��{Q�a�t�:��@��R����N�[t�Ľv�tm�O��6�[s�4���uz]�q�[[���G�����W���<�h8�Sͻ=]R�X����n��;S�\��/frs�uǵ�Y�x�Hݫin������N�ݑ�5v�7;[���(��/�5v�m�<��pv�TVG-��o{��t��9��fbI~X����..}<y:�orW<u�]u�)�(�(�fbf}�SX΍#�J�\�UG�J,�2���+1*�)L�#0��	C1K2�&f`Q3%R8�3�[:�O~lR0�[j�I|��/��!aDY�w`$]�t���$4!�W�:;ޛ'��2T��Qn\�^A?҉�g�\1��e��n��g�;ơΜ\(����U�&�1���!�h���׺
��(�x���idiJCVq�Zy����Ny�0[��LG�v��_M�6�ߖ�pG��H�T��<�vU]��
��a�+�߂vk�H
��{�ϰ���9R6AP��):Q�)�	�8�������0/��E��H�M��n[gi�?G�O���㍭��{-�)D\���bDHW���|���y�ڗ��,�$��-�r�ɒ� �MNȝ+�'T��Cp"���R;Y˃n�o;�&�i�Ux*�ku�Z������<��Gc����	�|�]�@;�y@�>���	��Z��s�kQ��Q� �=w�1���z��;�}�?������\_��6�yW�e���=��#(e���K:���h:�\���Ԭ�kllA���kq�4����)��˺a���W�\q	û�g�3����ϕ�k�m�z����[<�v��s���<o>�fۨuPy˻5��];6��" *<Q�[���$<�E��Z+�xq|$���	�����m&-���j}"��q�Rn�������wy�|[K-�bt&"��`	^�J�rr��?VZ�g �_�@�.��ˡz�x^g���G� ҉E[z9�x������V�Dd�J�v��F
�YPZ2��*�����x�ݍ��� �yꆆ|���i��TAQLS��ܓ�<���8�~Pφ`�r�V���	HNd�t�WV)$���4�����Ļ�vxJlt��c����ĺG�'Dч%�Ҫ�~�dAy��I�����2�U����2��\/R��KY`�E��V���E�Zx��>�� 8�֩�׻v:C�Uٲ��h�� �~�N�1�îN��.��о�=|��ٖ�ٕsj�4IT��+r�V6i�EO۵�|���wǆ�YB}��gF���L	쒕��L�D�&��5eb��s����H���Ұ��d\We��Y6k+(b5���hx���B)\��A�HK�>��i�8$� �	ʄun�II�����|���LEGB��6���q��_H�/W^B����*���E[R�(�Q��Өw���#��;O�>��|�N��,�<h���m��C�jQC�yF0[��	���7�ސ��#H��*A��,4�*�m�Ql�L�.�1�-���3���M%Q��sfn�~��hf\�R�aH��'F�ͭ��s^u�e����ErGHoi�t{�OӒ�#I:�$ETQ����V'��q��]^
/`�jF��k���
�ɑ=�����9�8���.y���J�{�31D����ə��B�g�<�I��í�g��'U�'�|CH���Ѿ�H�x�6d'Q��TI�� ���u�W9���z�؎\Wi�-�Ŗb!����?=p_܉�V��nc����]G�Yj	���t�Cնg���������*�*��ܣ���k������=��r����vB�$�nWz������' ��L��Bw����iQ��Y��1�C�A���vHk��]�D���aM��[~�۹�{�o%&R�@z��|p�ы7��/�iA�5k��7�'�?��pdDOݒG�;��W-��\zc'�]�����Y�-��@h>�+�p�KiaRUH��
}$��-�z���b���[���	��^��<�lϹ��MI$��&u�B���޿�"O�!��˄t�]��>0x5^$�.?P_-��Нa[���=We�_�=��;��!C<�y��*�	&H�n.��[�WHD1}�_T�7��,�k�!6�=`�Yں(#����f��8�K��&Iz�U�̰��L�l]��S=��Q���F'���$ܓ1�&z�C��M�s��N��"
���y%=�䑶��r�S�����}8{f�� m�v2��
t� $����w��&lc=�VhzF�����7~�s8{�9�1�0A��}Z��!����p��䒩!�ʜ{��Bk�{�A�~������BHw
�g�+2�-��a��MQg�Cl�8C�٣ǩ+T|��{����e�ky#��1R����&�c;0� Nc�le)�j�+�{�?�����-�	\�w!
d�CA�X��h;�<��ɔ�et&�=�2o����U���c��;�;���	$�-J�A�u\��z���Lp���Y�ʫc���>ɫ@�g�NZ�׭��m$�U���ڎ�\�3�J��Q+YMU��J5����l�4�b� ���]	�Bέ`�}!�Й}-BI<U�{��[flba��~���=��h������������B��6�a9VI]��FStPn�#������5\l:v���,�g���nB�,[>̦��;n7X`]��c���u���<(�w]���=�Y��xp�����zVZs&އ��K��h�Xڎ[��W�«=��.���>�W��`���Mb���QWl^�fǧN�B~�+WW=��0�C�m�A��5FRJὼ^<�WA�ְ\=6�@��ZE�Gsη��ߍHjZI%��+��4�w��P٩d�����˳�C��v_[�bwI���N�a��Dz���ZPg2�@L!v��X�Z��tЗ�.���줥S��4n�а�V
��_M@�PE�1�&a��2�4˹��l�n�K���SQ��ggq�Rt��e	��&!�4|Bg�ުF���
<�)v���6�C1���n��$��]Q#Q��Z(C@$�ߘ�{��7�S�NS�1p�{�*Rc${�Or��2�c,,�p��%����x� ���ց@���0�a��cع�ܳ/��,׃���B��+q�
���~�SM��y�f�t��-��^�d��4����n��($��8�O�j�"EŇ'fw��	����X1��$�"�+Q����~�J6�]���q����,�k��zk����˺򖧐>-�h1�z�ҥ��^Hc��y�V�牣���Đ�G�����B�!#��/�X��x�f3����������GH#��_�Xͩ�H!q���Dyܗ��C#N��/�F��ֆ�sj�i��-4���;��5h��~���U�v�"��3����.��ML���44��B���0�Q��7�Gڲ����9_+>#�i�ޏ��OX0D~�A��j�I�fa���>�C�1i���FeN�my�=>��u0x���yQ4��:�,ԜZ_y�M/T:t�p��3V;<(����.���\��a�G@�v�=,w�>��(�m,�-G�{M�#T�ګԍ3/[@��w�Y�xۛ���@���Yi�T��r|K/�7�f��G�x��]:��Pv�W4���X��#v�����&3��ύ�:���:��xW��2dg��=I�w��5���/�w�(��z��D�$�Y�r�u�BH�>0�Rة
����~L��o�Ö�W��L9�,ͣb
�����p�z9�Én$�,��cdK��L�cM���Ā�!���'��ƴ�F5"nLu�F!�2�'<k�*������'f��{ʞ�|P�$n���a�Z(�|ח�AS��>"t����0��w%!f�9��1hxF)�G��Xڦ�[�W|[�A�v9��,����o��WN�<��R�=��K5ڋ�����l�3j�C����Pj�Y,�	�D{%L�z��5j����b=Or�	��A]��F���#�Y��,T�	x��q���O�		v��cJ�z��o�#��H[��,�͗����ڎ!��דv�έ�F$J:l����Y�ܠ&��Q�?@!��,�zma�$b+u�ʷ�_\���R�2���xFaa����q����4�p���Q��0�e�TQJU,$�>��9��]9Yp��-�k�]���n�z����k`��A"G+��r��V�ND����^T��QJ�禷��K��| 뜭�{�/ES��T��S�TV��W� �:�椂���Q����P���?y_�̮ě0�"������fӵ�^�P!4�jq~��7R
�:U��R�%�mi�cݹ����o�`�;�g]!�q{em��7��+�����^���Sh��<��K�l�@g}ZUUA9�6-���ܻv=ؙ���q!q����E�c�we-���3�;u���]��;]�q�X9�R��v�K���Wo=�:�n�:vǰn��ph��J��?z�}_*܂[�ب�_����Cp�dL���M�=	��h�ax��o��
��E�i��g°P8����^��{�����wm�6tI��{t��܂>�Ns���S��1�t������$�#r�X�yiFYj2ǒ�8i����So��:���-}Cc�]�R����k�e��F{�p�$��5ɕ� I��Å���t
$Z_3��<}e}do&��bB��f��y_B�1��_+�|2i'}����v�H��uku]�a�M���t� �iK�4N����Ô1&v���)fOx�ّ���)�a�BƧ�B:|}n�)^�V
� 7��?T�ܑrF��.6wH�2�z���T���I��%�F�Ј{���fy1݉�v�hff/��1��;��}��>5����,���ET{�`$��YB&��wttn�e����%�^Y=�M슗�ˮ�*�vGnӼ�����I�\{+YԌ
L�Ȯ���j1=9�S��oVP�����}9L�4�h�3�Z�e`�����c� �ˈ�=&K�*�;N=����m!7�\�^9��,��(�qv(�Jy�U��ʋ��t��ho\�z�ͼ"g
��?��c��-[���q@��`��,��W�z��%I�L���Ʀ,��e70�Kv=�z��*�q���N)O��j^��v�.φ�t��wD�{9N��-Ņ��@x��!V�/6�(��V�v)\�9�bԫE�����@�|&��4T�Y��+��H�kB��5Tޏ���e��I6X�(��q�$
4�H	�!u�sl���: 2A���Ύ���nܽU$:-�G�.��)�o<��ܦ�.'����tɴ�,��=��N��щ�;sr]=m����m!rs�dw^�]l��k1��2�fQ�u�J�Y뛓\��s��ѷ[�sur���K����y���p\n�WC�}Q����}�8��^w'=]��v�#�'�<����5n��9&��k�[�c���	ю.���$ǀ_V�4��U&�⪽�*��8�{u��8��ϲ�2���Bn5҅�囝���ɵ-��d�Bxv�k��ȧnz=�;Y��<<����$��q��gv��،�w]cn�N�]"�`���{:�OKrqnAk��t���̸��&:ؽy�݃�[V�����9�q�bx��rn�jH� ��^ñ�>:n��qp�.���l�W,⓻b�(�v�6ڜͼ��3�)G0��b�E�z��{v��k]G,���nf�펹�i�������w���m�DlL!p�`.�=�s�q*�Yb�l�'�R����f%�8 K��Z3?��P���L�`,bV5�7���{�LK��V�8�,]mb�gE^13�S�8&-�6+Z�	(&f{}����jQB�'��[xB8n��.M����䘘����FĶd3�P^L�/�L�.	�o��y���	p^�itXŞb����������[P�X�xvL�Z����sSoi _�"͋B����i%�b�$�؏�:*f��E�j,zy�b��ň1.�b�_�QA$ę���38'��׈�tX����V�B<dB�Q���6��ږ���b�[@�.
m���&36-
L�Z11/k貉^k���;+��&$��f&f���rd��v��f���b�ƒ����^Q)�M�J����Apf%���#OD��c1�^��Ί-�&(d�LL����K��V�=ߚ*����Ab��ŝFC��yE�'�G��n��6bٟ
���V� Ğ�)�-G���������(�&,P�������y��?n�k6S�$ň1^�PZlYE�yȿ?m�1Cr�<�7�(/��b[7C1�{"@���b_o�fk��B��^��i�����=�w5��<cpI��5t[��x_G���%\130��X�ϣ̂Вb��bbZ3FA(e�b���u��D�/Pb_��uo[Y��|$Ķ|$Q�bfc1��Ι��(�$�ilL^��6SGD�����8�Z�͙���LJ��7�b���*�Y�A�$�?��b鉙���jm=��n�%m����⁹��x ����b����=�{�էL_�Ƨ�hIAbm�bLP��Z�f�$	3bV<�g���,@��J�=LKb�lЖ����f-�����}�]9��4|�&��G���J*ݻ�&�v7R�gQN��kA��Í���>�@ozw�.Q�f��Ũ��	/��2���|�)�LP^pPJ�1�u�	-F����.�1&,@�fr��k�Y�S1<�NW��kU��Xļ,@�,��%��]Z3�KF/�LX����1��Z��q1ˬI.���:b���Y�}�X�6d1&z<eAbm��c�bJ�(&gߞd��3B�J33Ц���8 ��$�T�űQd4/ ���ٛ34C˿��I|b�$	j4����d-G�z8eоW�!!�� ī`�b���bf&-k��-	~v<Θ�P��H K�ڋ~ilK�����?U�io��衚3�|�/F�����gM�5�X�.���k�g>�4b��2��u��hY���P^�"H~��'�[t���kA~M���2��$X�)樖�� X�lI3�ň2�}���ٙ�]8.
�$�ȭk%�	"��:�%����^(�g�o}��s;Z�$��K�j�E�dqF��pJ��FAAb_���%��ŔI�s��G%Uͮ	lTY�_V��1Abٙ�k6s�ųBPX�b���t��zru���k�|�ũ�]�����VV�����~�4b�(pTf$����B��gL}�ţ3f|%��{�bΝ6$��C�LT[L�LJ����D��{38��3)�X�kf?_�]���x��y3_5\��|��gLZ13�$6�]KV&csn�c�S!�q�,@���Z11}��C�X�y�P��	*&$ϋ�������,�И�TJ��*/��L���?}2�bb�X� K��,^35���TK�����*�flT�/����)�B�4��լ@��}�P����~͟� J� e�ò:*J'�n��.��T!t���9��4��1&2ICLL��詜5�$ň1/��LA�I�E��b��^LbѴD�f\v5�1/NJpę��{��6,���9����Z�pŪ��bT��~��t�{y��g6҇MЙ�?P�o݋5�Ŋ�,�/������8�p��Ĩ��8����n��E�PLX�l���h��l�`/	��X��&,<�b��U%�b�2����&bg`%'��Z_w�.�\r�K�ر6���|��i{��<,A��b�K��L���13�%#LPYP����υ��bfk܋:omb�*e1p������Z038-y�� ��Z{OHzZ��fc3�K����KBb�PY��13BٙkT�O�C3�}��%��bτ��͉A.
�Ab�kb�kM����¦``b�K� ��{�߯��0�$A�`M��O����fns,��~�b{�%�)ǟ ZC�LP��#�g+IQ1b�b�Ή س��-��鉐LЖ�P�F(d0+^1C����ͯߧ�/sҙ�[�_��E�Pľ�~1A2�ZZ����ϛ@�,�z300lb���������m�����TP�(a�K�L��7�K�����p��AxH�lI1-�/�X�M5��&�[1300(�1&g�&,�߽���8�*��S�:Ί�\)�	^r,*�Z��š%�b�1.	�E� �E���h]��A�1$�Z3B�y��LZ��yD�����8b��(f�I��1��3�%{��]��G��z�ь��b@�bfS�ߢ�	}�t�R���В���(fx���vd3]y�IlLX�b�3;��E���L�W������o�~q��.nB�}Ǒލkp'�N��E�v*�uа{H4�� ��v�k��v˼��nܜ�����b��b����+w�H�>�h��|q�ݓ-���ݷ�l�p��e6x��L�(v{K��,z���|����o�u��J|-�P�Z���>y�1�$�֏"�lZ1��(,@��7_i�1&*1'>�;��%4����X�6%�@3>�������-�si�13<(,��=����_��	y�P1 ��(����1�tI3M
?�01h�����fS�$ň:bL��E�VQbq����.F��}�f�W����C�yD�1b�,O�pI�)�#[3=���[��ؾ���}�C!��ė�X�2Q��wȒ�� ��yE�1hC����`A�((��j����Q����F�uw)�.�	{�D	m�24*bP�<KC3��X�*f��f���	B��	tY�ى1-�my�X�3��Z��LZ[��{��1Aw_�*`'���ߜ��md�X��O�(���(%�زƱ3G�]!���ъ���y����Ţ�,@��LJ�b���������̢L̻�l@�F�F� Yw�%�5�bI��h𘩟��d3��.	Bf��Y�4����ɹXm`��01���	*&e �b�ƶh]?}���絞<b���&`,Zmb��o��o3bf1p��I�34(*$��Zk ����[3�r�dC��,@��n,���/[�{_�z�/��,�P�(f��~��9���-��q���=�;�[[��B�!˰Mh�gI��H��"�1�����C���i�r7"�*>Is�XJ������h�f]Z�
h�$8���������9�Y����(mtL^�f^%\��3z���2
��wH�X9�������65ܰ��{P_g�۪L$�whqrٷ�ԛ��6fnbc����v$��n&�{��KBd�� a떮l�A�QOh��L/���/{�Xu�1��_9$���fq7H-�G��bi��?v�<-�-&O6O0���א���s:7��n-rIh\M[cߘ�RI�>��j�9��]�	9����844�Ɓ���M��WuT��蛍v5��j����ęB�{� ��q��J��ƛ�@$���J�m`5�ُ֨ޡ��9�P�U<�y����<JVD$ڤB8f�C��M��C!=�Y!#m�1�8�F�2�ʼ���`qR�nx	.ϻ����v��И��ol�.���w����,(�_��A��Bz)�.�#��c���W�,�n�g��nj�Q�(d���6r���)�V#�[�^
�����=C�վNF��B��2�5>#�&W�8֛�KB�ԟ[�x��]/�]k���qwy�N���M�OZ��0�T8p���o�ڋ�TmAF�:�Z(��wu�S�s �~4x��E�yP����h�6(r��55�pd͍{c�r����$כ�����!I�������g�ٸ�uv5�W�#F��Ike]S%��¹]2�Ǡ��rgݙ�Ū��RS@�K=���.m�t{�CV�G�Bgs���l��u
Đc�e��.u	.]�\��P]���`킨���-x�}��9�"�d�IM]K�&�*C5m˛s3�q	ë�5�Y��%����T��������wJ�}��j��n��7Tc�ݥ�
L�<�E�WW��p�Y��g+�Yif�FP�;��w�t��	.\�ZE07#��j#�(����R �@��{�ˤ<f�Eh�cz��]tK��M�@O�[l��#�F�O�a�N��;ӲP�*tee�����x��sR���m]��
m"�=�����OZޠ��B��䱞�t]i������! ��nM��4�0�݂٦�=���]��;h�;v3:Aʼ��(5�"��}�������O�Y�@J|:��u惮E���c<��p�y�*�㚏��YV�Il�ڪzZ˓�}"�?4��+�?#wrq�A8ry>�XF$/ݝ�T�����S�U8x�Iy��$"��pE"+���un.�&	ȅ�꽪�ڶ�-��Z��xp����R����r�Ƈ�:�����3�a�Q�t][�>;���Ɵ��GȜ��^��n3�V��b��:q��i3H�:�_鸳"}!�D�q�[���r]q�� ֝M�#�&�:�̈́�,��fb�,.���p�}���4�'79E�`�ͭ�O=C�9���t�㍴s�q��g�j�!s�>{2���8v9��)���m{ο+������0ެ�5��x�6x\p�>DWN�����"�Y�`��'�
"�*Y�!�H���`��,�%eo�0L{y�
U��4�v|@���tQ2�J�|�#m�ӔnEy�,j"��o2�n����ɴUBC\����6�T�"�-}`���~V�'/�}�1��]��1�G�F�����a&X �j��v��+զ����t�KW�꺕�����G�s���-`PK����+�Ė�;HQ�L.VJ\E�}����9�7��q�S�3�����RUaQ%¯hZB�{��+�Y@�� p���~ Ai�囩xy`(��,��!Ң���^����7̢���^M���(�:�7k{Y�i|o
��a n��-P���w�+{7�N�|�Yr��s��*�nU��������u�����+�h��,��] ? +3��"��F�@x��&*)�y�b���S��˛@<)�v]���5��;��6DP��r�Q3�ǹY�̚�T6�m&볭��r����!2Nxǭjg��}ǵW��J�Rp���VZ�F̮a�5ٲ˲�㋸�M��1W�����q�y\#�$�!��b�����n�s" ׻�H,$G�'��08�w]P:���x�zwN�|L�Lytk�a�.��5�Z�!9���ȃ���*��IhЌw]K����4$T@|��O���z�BHQ���(������B�d�O{4����w |�^��(ğ�����2hz����5�����V�6��+z�;��r��<n�WB	�]Z�{olg��G�H�)FZ�&	*U��r֗�DB�Z�~G\�-KG�<�>�E�]m�˱X��D0,�ۘ$��y���]���<$�`9I�a�m5k�G�_�
/�� E'J�����J�g��9�, �p�=�V1��4"[Q�Ed�y���$���R�5j��%Iu�e�Ӳ3t�k�_$2���Bɼe[�y�R|A����uRh�Ad��g����]��ran� 0[�����p��/��+�EY��<��b������3�ݫC���Q��-�l�Vd){��j��W�S��F+<Ɵ���t/��2�vqH�&�e�Z���
DZ�;%�B�h5�̿V-s��[�o���k����̧0�L��lm�#��f�>B���i|p��OĄT���o*�JX�nI9��0��h>G���"�� �J[�?�����l:؏���W���I��5�A���c}ۚ��Y�m끠mA���8~;�]�T�j{u�q`�Y��﹠e���e�C�C���P]���+��WE�3KY۩ˉ�u]'�Q�R�A0[�o*�ݖ�;S��nf٦�t�g��r�ʴ+#��3&^��m��ڵ��Ϻ r���:�]��y��y��gSe˪
����T~��s�u��M7$�;���}%��	o���K^�[#���y �D�F�*�G�u��=Ы�N�$$))/e�S��X�a�ᇨ�T�?�)c��wx�t�Ckqw;�����{�ðegW��7G,x�;5�0̒���s��r�k�ؖ<����2'�\}�V����J���';���E�_��ߜ(�A�S����?�>0�޾�Zx&��2���r�����c�6x��"A$Z�C"�yh�g�B�Em�?�]]]�C�q���%)�j*+�{+ 1���;�7�����!���#�p�i���u^�tu��eIڨ��d�I�����².�*�}a(��-	UX~�"��E�K{R�k�#4��Z�#�K�2)1Y�A�z}�݇���료r��#,!VT��ջ���Vc<c�rH���P#}�F�.�DMvP��@	$��~���o��ԣ$6�P'�� ���M�I����oE�o$zG���(A�IEu�^�A����sg��h�zA3h�p�4H"�ٴ�Rk�O4����HWe5šXm5e���P2<�J��V����iv]L9��4$r�H�2�'
������">*D��Eƨ��<���ܼsJ�U���m��,�lo�D�>�+��Z3��
��)Sa�@m�L
n��ݵ��2��v�t��Qq\;z2�h1��9��+�,������;�F��:\Hv��v��r�7g\繁�B&�ܝu��q��z�mU�>y�]��+���� ʿY_���"{�Ӿ�n��]�DE�jm�&]��H�sA:A���#�X�r�#����������)|��h�ha���+]�����	F�@�CMH=�;v��w�؇tn�ʛ7���{wzZ8�1�E�QGLp��� �u5[��"K��=(}����)��viU]Dk�	?y%�MKu�ͪ�gr�ɣ9����և3�i�i���ɛޮ��
=M��ܲ8�m�$'=2ϯc���(�Z3��^�l_ڔ����6��1n���0����+Մ��6@�#>����jF�Bim�=`�|�+�Ӆs��h�($�%iLCsB:ς���k[P��F"�\^[��z�N�k1T����tJ 5�L ԇ�8�u>z��H� �/�����-uTf�I��V~�~@���*�Bn�zS��z��+|li��<D�V�^�<.���.��NRё�:u�GC�=������#?)o�R�������0Qt�A81�֞�S��;�:*��J�L$�\S�yïSh�z8ѿ>�?_�������"�Bo݆*+��TI��@srLAH�}k���+��G���\�OH�y�m��o��N���E������*����5��h�8��ƈ&��n-�U�]Q5VHо���W�·No%t@�C���U�isvj��k�b���+klx[K�ګ���'�yG�S.�P`#[�+^�;�Z����c�y��wfZ�f�yZѻHrD����GqX���V�ت��3��e�;��-�@��{G���}@�:0�k͠�I��p���d�� ����&��H��"yԪ�y
~A��$�J�XƏ�ZI�{�$ű	LV���)���]�,�>�l@���4����`�勞���H�hJښP��V6-!�V�s؊�^�+r��22��M��ncǩ�t/�uk�N�*��on�՞�w�l�7KbZg�ٶ��N����2�L4��	�v���z���*U`i�X�����$r@׻�Qх��A�D����x�ƽ}y���B\ۮyܠ�D�Aj1c�;gC��
��3��M�>��k �O�H�ɻ޾�u�1
|GBrd���|��0fa��-i`�X��=���X�Ҭ\��s���~���e���4�.�a�Կ_q/�0ً	$7^C��L�J(�n�g�c5�K�����{��c�:j �	��|2<�b��BjD�V[�k�Ur���
�j"j7�Ҩ���P�^�q�=�(��S'��g��dP��Ѳv�yz�n���'5�uQi
h���SP?�Ɓ�o����4"��b��˷�|�.�$��ыD.1D�l�[Pz7��y�CP^u $	#���y���^CO�+M��#����cH��I�C	CD����R5�U������U[~X��-_펹Bд#�X����
W�ə����?|Dx��4Q��S7���";]���~������n �����oDP�ւ�dƴ�+�|i���C!i	�p�1OLT-���a�ɪKV�m���� �x��,�	�
�{�{��'_+W�\� ���Jb��]�@:)|E�pXY�o1Ya�&�)�����C���X>{�c<F��}�����_�Mt�}KΦb7m�[��cBϵ9z��r͛�cy{P�~�zj/}�|i�#!Z�]`^<�֬$	ay�X兔ʪi��U;��Јܭ��j�=mR�#����p=��`.1���~�$��v����n��B���w |�`/'�dVدWD)�S��:gy�����H1"O�`����H:}���W�1�,�J���꣇R�W��/44{�ԓ1If�#��p�v#��������޿;�G�����U�>݆�Փ[��@�E�1�&��P��jfu��R?��$��H�ԑ
��g\�8�A]֍Π�J"��U𭛁>!s��t��-��cse:.@7Q��C����=�m<s�ؼf��u�c�m�
��;��7S<m�;<=n��9ק<��O	��tC����ލ+ؤo���zʾ� �]���uԫ*�C�o�C�V�H��ϝ17%���dVr#!9F��I��$�])��]�f'uh�vμ�vg*#H�n��˛2��8�6�v�Dc1�)=����8bMvm{�Sv^q=��n�n�c<4n���Qn۳�h{�-����Ut�
)%37�>�(JΊ��h48\HT�=�,:��8h���b`AM�ϯ)a
�H�BzA<lc]����2�b�)I�6���b_k�a���M��$ ��d&�<�C5m�Zk.�đܟg��]�ߝ1u� �/��'b�WС�h�G�w-/�?o�oW��YHت4��
�����8A1Q���R������Y7lf�5&����p"J=�bU�w�	7�"
��=�!"��P�/:�bȺ�B���=L+%Y���R�r�蹔t�v��~�q��Pi~m�������^9p��]c�G@���r8j���7"A�!�$ �X�pd��O}d�
4��}��<wse�{b	��^�L�:��/�3C� �y3w�tm� �K����~ �?M�.=q�Z��>4E��'ptQ�ia*��j��8˺$� ���-�-��U��e���U���A�byD�80׌|/K�++�X�bW��Wթ:^�=ͧ�GXGBBVU�
��a}�m�U�@��n��l,2����z�A���r�w��ڴ:Al��?�4BVę4H�>�#���b@{�@A�n끳�DB��Z>�B�I�W.h�nw[� �tOh(>I,E@��`u�
n��]"!*ܷ
��qH>���\")1،n��0m8�E��{;ח��� �4�n��#�q8�ƪ�d
�+�pӾ=����-ir�j��d�K�>����^�4�^��}>N��nAI�U�����$�L#��Y��#}n=�;S�uS���T�!Zl�,>�! �g4�ۧ��������l�T����OL�'�{.M2>�M�i��ɑZ���R&���}5o-�f�"��ʰ��,E['םbl��I*L.��M�����n�|���
[�*:���1DY�bR����#hU�N�υJ�9#~lq$"E���B\l0�Aewe��qB�r���[%��l��>�C&�\��e�*���A���8q����s9=ky )�PGJ�GХ �r24�jв��2 B8��w����������lgܩfx�^mU�Ko5��|M۔<4'��!g�*|��h��U�/�x�쮞���|��� �i�^�t��	$�<�C�aPJ ���.=^^�'��7�������ھ�*�$��P��P���wm�Ns×ɮ,ː�.ܟR��� ;���l,b�s(%s�"�����nr�XLG|�(|B�RJ7�f-����U���ȍ�t��_(6�|T�I�bg׌QT���c�<҃�hf�r�u�W���ICw*��A5��P��i�����	�A6��0�w�w0�b8�Mi��oS� ��g*�5��S"��|\Z��f�qW�~�����ib��|V���ܺx=FR��5K)�!�����U,g�n@�6A���Hs�lZG�d�A��
�	z��_;���p��� P��[
�j �$��w����"�F*�rg�/e!p���"A����H&��ݷ`�
�è�G#����@�h%��X��t��-L�&��%$�,��I�J����lǮ�".��z]��wT'mʫخ�l�[W��ѕ�ʹ������^:�"jYd��-x\=9�\u�nq;���qۗ9���h@�$�z���^����αuڗ�x�v�X��OI�`#m�Ն�yڎb{'�.8����-�����uv6���^<�P�KѶ�����ꢟI�379}�1�Va���ؓoaY��~�z;�A�����y�,G{���!��{)�Y!�����k*��<��R[t"l%��򱫛\�a#��o�;��k�����W���2I�7J�lz�6��{��~}��Py�
<R]��j�oyr1�P��φ�s��=��ٰ�t8D�|��d��"�kǥ��!#i�9fUu��f��5Я�O(��D�2�D������2�>�`��{6�X���pny4��U��"E�>j ޟ{�9 Z�Th�:)ޱr�D�gs:�N��&(��}�a�o:���	�d"���~�_�0�t��7ʈ�Qi7�Kp�A!vl!�r�-3�]�5'd
:C��ժ�AܙIiF�P��2�AI0��:u�V;�*���]uU�9g���	���[F��S["�W�1N���}��`;wU��W9wkghoLKG�{@w9eo)�\јv�VzW7ۺ�=ٌl��vt�ZD1�L��U����%���"\ܪͱ�rmeV�g	6 ��ūV��\��u��F�Uމ|�V]�ߛ|��.�YF
;5����۬8�D'�oT�SW(&f���D��u{FK:5WX�|�z֧��}k2J���5���C�NP��T�����}qS�f�[��X�^W9�ds$��:�2���*�i����6��rKae<q�u��Ш��;�pd��1H:����M�#.��w���a��N��ͱ+o
F�f��T-�b]c�NC����,��E�!�M.{GM��-Uڨ5R����F�i�ML����Q��4�UU*� [$S���CHn�W#Y��&�g�8j�[[�&{U;���ܾ��فn�q�C�^qr�#�ت�o0f��ת�Q��p]u�p�u�<��`�3e6g^!����Ň�w&2M�1X݂�e,�0���nN��ls�*��n��q�@�V�����<�#�Ѕṫ��m�n-����j^�q���#����f�z@�sk01=ۢ�KZ�a�u�	�.��k��=b^�Q�^��8�$�u@;y4�qW5'SnG�oIc�n
u���e�n���6ۇ��5���1���w��pz=��c�[e�z�<;���8ּ��{77�ݰ�;lN�ܱ�@L[lX��*��_�cZ������������ƧZs�Ѯc+��מ��:��۷�ni���88�
��Éֳa`7I�A�vs���9m��t��47k�^=u�9�*\a��I�m:o1�F�����k���St]c2�0m���hI6�т;v��Nw�<u�Wog�,��Uh��̳�����M&�m��y�TL�4j�BrQ�P!Z�0�.~<x2��ٛ*���>�}eQ�Ovsqq�=<;I�sļw��\<��#�uޟ��$-�D�pyi�C"���;����#��|3;wV��I,}5|�^��̭��^�� ��,Va��w��+W�6�)�A����aV:��\ed9fY��_eS�{4eQ<p����m��u�K֊�뎍^\r� :��g��}��+a-�|��8j>��z8΄��X3ތ��������Сf�.������$bgvo/ϛj'�;�����yh��[kADM��Ibl �?q��Hi9�����2�Ұ�D��[�w}��M���>������oI�;�Eo�r�r�󰌔-ps͓��r��vy���W�W=�GE��S�3,|�9�4t�K�"/��Y��-��^)!��"hw4�҅�[��KsE�!Z!y��ʺ3�o�����1$2�0�����"6��0Y�Hi��=���E_RO[��YJ�%���Lu���e�r�mQ�,�P��9w;�mp�Mz݂#��.��@ �&��P�
�0/S8P�:�Rm����`��^Ϣ����3u�>�(��P�MXL��'rgh^*�+�~�68I'�B�m�&�MX�*�+)���Z�$�p�\�^���\����ӭ3�76FW�`���`-��i5��E]�R����	�F������r���U;=� 6�堵�\��P1HK	c�U��ZN$�|��Cיdo�'����� �e��l�v����	�S�=�L� �$;�Q�`x1��@��x��Vg8���"��W���6�2��W�q�]��ٹI���N�>n�ˋ����㙠�9c�Ǚ�7L,aWO>�z��Fv]_-N#����&�]�k��a��t��(�T��i���}�����J
�k�Rj���yH�u$�������hW>���o�k�+9Q��8So���H��]i��mʀ�gpI�2�U�;hit��(?-*���gP��5���GW&��6z�mz��D��xe��J�7��!���Y#5��c��aM�˭�q�sk����"�5'��i���I��"{O����O�cՖ,��Rz�tM9�8zI �,g�Ҷ�P{;�fۘ�+#^���">���|\L0_^U��Т��<O{��d�<mۏ��@�-RQf�2��Xѡ�P�6���HinS��G��хj��yŜ	�co��oS�v�a3�?�j��|a ��iC[FMn�uc�W쯦}�+WCt8��wبd>�]A�w���������V�"g\t�Z��d�!��N��S���kPZ��f���������W/���M�E#0�k-b���ջt�m��L�g	ٵ�u���qI�t฀�C�FԮ�j��Eb�~�o�OEB~tG#��A�����H�+1���x��	h�*T}7�����Z�O�f:�#Ud��:"��J��(�<<��M�����`5`2� �D>^���I�J9*�0;��A�V ��7����Mv�Ϫ����xiJ��6�Qr��,Ia��%[r�,1�3؃�	�(~�)5�lz��R|V��J�+��2����c���V� o��8Ʒ3jj�Q[�O��PV'�BA��zr�>���4V��P�>��۸<4�����!��@�m���o�}y(�y�D��V3o�7�O�buUUg�<�I�p�I"j����(H��	g1ͯu:7��̑F���W���x0���.�4�ː۵��>�V�N@��7��kǉŤQ$��ͨ�?�%��Fe��@�P��ès��[s{i��ڷ�p��������G<����t!�b�2� !Kx�����L|&(N*���.���s�n�0JE�C�{���F#|9�M�L~y4�( s:��/��)7�oB.ׇ^���8����+���ٞXAlm�d+�����Zڇγ�뼵����ބUQ(�zt���!(������i�r.F/5\�G�<u�?w�
:��c�/z�5����֢?&� �*��U�0���B��u#&p.(��^����	�mx��h�BB���qE���/��u���) 5K<?z���}Up�Gg���p�)�!�\�MS���O+�`�ǳ��;�5}t��DEsΎZ�B����l�'JW�H�ۊ�t����v�Gv:���ż�q�������p���ao$e��7b� ��r8q� ��G�R����wH��}t�z���D�g��~��G���a�Q�C\����j��a���d�-j3�NT&�o܁��B�a��$`��vw���q�]���.��5��&ƫ�=3 2��8�%��ƍ)۳KL�%�G}�ԑ����z�;b]m�!b�y=1�AI
M^�լ!D�'ž��;�#H%C�凨|�s��Mq�2
[��(��b@[�w���q;UPB�:l.�B4�I>�܁�e���5�_�A��W�
&�){��ԼEr�N�?o��!��bo�|b}3b5-�eDv�҆��B�ή�B��Ō�U�Mׯ�����IB���ү�'Js��ӕ��)6$�z<<��4���
�fdo�E�����?/w3B�M
�(�w>�rB��r\�P�	HVSRԙ�Nlz��D��"�f����Ҕh�ZSuĕN��q�����5��~C�e7�YO�9>���THEg�%~ђ2iF1>�D?(v/E_B�w.؅'S���l��A����u��Ƣ�V�:*���؉$w�>�ޞp'N��(ў��[p�Du����1Q�����҉��{���V���Yג���Mǽ��#`_�
�����=��{ �)�r}�jU˄�t+M4�CQ<��J�s�wk6��������F;x�~Ru�ћ?" J�8;��$%«ӹGm(Ac���{��y��MƼ�������K�(�m���ԍ���[a�c5�4�<�d]싛yZY=��a$�fGlN(���ޡt��(B��W[V2}ވ�az����DM>�9[��jl|�����hJ�@���e]'v�l�N���h�ֿ��5�+P˴����1_LlH�0w��ο�XB�@�D;
�CY�Bͯ�?zo��e��t����~�:�=�$��w6*ՙv��i�H�~�I�٘Q��8��B�h���nU���l`�c8�vBn����<�Ł|6�p���]��=j��۞�y���ۦ�ٛ�Ǉ�.��[]rY&ӻu��3�;R'X���\��+�D��]%u:�-*����d&��d]f"��J�}ͳR),ҽIM����}���?D7���i�d{j4�����	�MB�Z��b�UsS�ԗ��+}�'��'���b��w�۷���,�����Kh[e ⨢t-���k�I���n��zЯ^���P&�S�}�|$�ӽ��gl% *���R��k�5w^���MQ�N�/�%i|�.d����{�2<H���N�ey� ��j�b��Zݼ>�˿L��ϴCÉ���,x5r�6[7���_]賂����p�g{�EJ;泞ck���c���L(��{�{��iӍw~�(s��̹ޗ�z��ڶ��n�`�2��f����e�t��u��C�2�9�<���Ax�������$�@�ꚢ��oU�Rtr���a2D�A�\m��U�L�������.�hw�2���<
�r�G�ixR��bcd׽a�{ޣ�k7t��u�/��E1��@��Kד��s�;�jQ�~����(Y��3�<5uQ\��b����M0=3�P'�X)���BV��������K�(k�7�Q�W[�Ϧ�����5V�$ٟQq�g����to�'������trI��v{�����//`|j\��z����'�v_&W9םv��3b�5��VF���E�%����0^#\~~o�n��Ƞچ��t�Wv�bf����Oo�:p ���r�����#u��)�a��{������4�"as��z�tҮ-x�\�����)�r>�ٕ�����!�޾S�Q�:�OeV<�>��w[�B�:�S炸������_�k����$B	����k�W��^�K;��
���Ӭ�����$���UrA� �����(��縫Y�$<���[Z)D��7Xr�@�y'����vh��^����{�C��̱�j�Ra>y}xW!��R��JR�p4v��ɝ�] ܁%)��n���`ƜG�>0E4_�z�B{ަ���|��_���c��![���|�#R���n`�����_�e8�5K���,4HSk��8���YGo�\
��3�e�Ӕ��g�e)=�Pv������玺�=R�m�N�z�IXe*����`~�/i�9��J�U�܈h8��샯$�x)�M_p�[eł��W2�ޕ�1���[1w��ͺ����Xl�:�l<� aG#��v�k:�2���ث�W�_
nt�����Bqo��^C�s�n��&�e�S���:!��#
ǫ�I>*��Z�첲�x�}�U�d,{�6Щ}v���69ج�S���Wo"���tSF�%�@���_Y���.���ml��d�W'�h��[=��䡵v�U���YX@:���T\n�N���nɡ���L��$��q��W�f�"�NWNF���>�%w'iV�;2�B�w�s�JI�ρ����>ߘ��K�wk�~p*���b	�:x>�����_�oĹ���f`�
�F{�>>T�d.��*���K�x�W7IR�gjH��"��+��ب>1:�B�!9�٭��&�l��V�ș;�X\�+)�Hv��D"�=��QYT}�C�_5�����#���؉kP�6ɇ�ؐ4J���x�i���ǩx�hW/�E��~�6�����Ϻ��5�]w�\�����AP����^����G��i�������gb�ϛ�1���wVо�Y;�>��G�
���q脿�耥ȟ��������׼�*�̇��k�<�л������ӹ�4�A�w5a6d�����4�����	\��;H]�s�3��9��r!Ŭ6�.]�i*޵A�i67<��ώ��r����e���_Τ;�ѳ�m�T��WcZ�uq�YQ�����y��5I�25&4XH�6TNsc��@O��<���3�����"�<Q��:���4�F��7cT��D5�Y�����R���~��&���z�r:�i�xNד�vG{�� F����E���Uۚ��2in��6�~���}}�:�`=^��p4��;hv��Rϥq��$25j����5����fo{�E��yn��ܜ�Yt1X�w {�p'���۱kn�ud��h�F��;X�CEE����[Ë���_��p9�&ꮖ!,��E�L���� =����m�����P�<�{��y�D��n�������O9�����G���@Z{.Vױ��������^_7O3]b.�Wvw@��]|���BJ�n�i~���즃���R�C�#{��o��=wܼ~8q��ʥMF*���Q��9�ƙ0 ����%�˽���k�����۴�>�e��L�꪿{�՗i�ӷ�}W�&C��p��j��u�gP���>�wBQ��q�Y}�@�N��&�cօ=�aD7m��@�uj�h���s��7�r��f��˱��R#$^Ъc�:��tl&643~����gv�Hdpw����ܷy���1�����������p�z-e{z��~�{��rG ��R����Hz/w��X�"�c�JD�%r�q��B��1���������n�oZ��u��8+��
.�T�-ћ��I��V(9���3������C��`�y���U?��(��O��IHoFa��фl�ʬ�y�Z�����C�W�]pY�Zr�OPOi\��l]ȶQ��{��nK�u�����Q�F�$O���A�3�ߩ
sճ����x ~��z���=9��u ��ʡ]�>"{qp��Y�u�2n�|sqK���
#�{Ά�^g�����n�]G$�n�i�"dLb�Z��;�bv�T�i>�Ǘu�5��Q��I��j���t�e�߳D���x�I�y+V&\}��*¬ߺR�~ˤ
<P��<\����ͽ\p/�];�LZ ���G%�hV/�eC��͕�
��?m�?6���oS�z�n������Z�Wɿ�3Q����h�t���U���3�=~�����OU�	���xy�������Mr����\��õ������I���o{���޼�l��hY5���e�}�íl��=�гAa^k���o�{�K�^��-�d��:���͛�,�ۄ��h)�{}�"7܏�GO�fXt�$E} eh%^w*��̸+�����v	�Tn,;�Z��j��{މ������=���w}�����
��$���?o\��n����ֶ}�|�x���P�uZ��+���X�K�0�&x���DqH���:�Vc~v�s���/)3���|�(�z	5J��\�@�Ua��`��<n@��98�>�zg���7^y�׍�Ȧ�2ӷ:�ظkq�ۑ�m��n@A�^v��yW��DU�x��jN-vks̓�t��1H�n����Qb��}�uAG��!�{��2B<<�d�H�LZ|s,a�Dܒ����j��̾��AXȼ�A��-'�l�{<�C�eN�t"  �����t��l�u�Z!+�=�Y�}��7q+`��䌨rg3è&��y�?����!m��uf�����e��V��Ф��Y�CA�D�[ڱ꾷�6?z�k��~��
��6���+�#,d�.���2�(�y����u垝��&l�X�g���E��'vGolɌ+ˀ�*�+�U��D'<Lg7w䧷���3x[��M��,� Z��J��sX��_�a����-�g�GV�Ț}��kX�Sk�r��x �~���%TA�ڨ�w|��襣@�[P��%B�14B*bH$���g���z{{�k'-��d�W�y�Z޿Ɗ��K��=ki��؅p��B���xE%mv��L��.�!'��YY9��v96�X�4}VE�� /+_�K�z����/��m\�����jߒ�'U�Q�Ű�I���1�pN�4�u�D���,_nj����to�
\42b�J��k�=������'H{�	{�in^K�(�ו=�Ut~��8�]�s\�uݷ�
�i`�A{@��*�� �*�q6�ґ�S��Dk׼��/����s���i�&k�V/�z�����V���I��c������4_^ǂ�}kT�q�۽̔=���C�]��X ����;�n_M�������V8Nͽ��=~��1W:�Y)��]��^�kV�i,����t�����{�\�<��a�8&/��\��=~޳�{��+�ݞ�S���.Ӯ��[�yln��Li!UǻٓAy�IiW-���f�p�����}��P�"����%n�KG�D����V)��W��ת)��˧���#����y�ם�݂y�����n���[A�ѕ,Kő��Ӗ�cpx�;P��K�*�.���P��L\��?w�=q�Q�T�㮮��Fm^�l$=�T����*��n�]��mc���t%'0�>�QŘi����s��ϊs�r/D��O�z.��	�K2�zkˡr�߽8k�Vz�xUҌs����}����arކ����{�r�!t�ٗ%o
�^5뿣��cV���4�w�A�+�~�-nv_<�ʜl��-CJ?��
-+h���aH�Kp������y�Ix;r3�p�݀�W�aW,��}���rኖ(rJ�T�Vѿe�9���U�}�^��nz�S�-�Zׂ�ϲ����^�wKGn��|O��p{p{}���0$8A���<g��0:��	�zeˉ�[���o�C�%���<� [������p���f�5�E;ڴhG��m4ۖѩ@vZg�x_<�i4]=�zM;�p����qJ��A�Gmؘ�����wT��#��]�m.�e��B)�%v���lOV���!�]Q9mB�������#�����û=�����x���b�=�xK�Q��(���z ���A�8�OW0e������8�Uدv=wz�JM_�MA�L�h $qH��p!�&�	L�ݾ+�w�Ʊ��t��~��ڿi^#d��V�(��=���̺�]�8��m\�A[���E�~�)��n_�G����2ǯiJ��vf=�*.�9�׹WY��5�^��::=��\@���/-��q]�{���2z�25�:��,���|��{qOwRRի���\����=�{�
�,)�s�6��r�+���{�R�?�;:��ę,))���k��mY�����������{�:{��4�䚽وG��]�l�ۗ�����.���&f�j�7y��(�D;7� �,�[�������^�X����vP2�A-���ewt�L�o���+�(�<s���TI�}-Q��K�U�D�0D<A��q���Sf�m���v*�y]ʹS�����-r�����ce��H�v:`�X���B���v�n��j�z�yq����:
�WmҾ*K�u*W6�Cl*��)��ev���iꆥ.�r�5{��mُ��/�����nǗ���3l��4�V��C��`�⼠�և�fM�Ed�Hv�;��fJ�r�:;*�v�2s,��Cs�ݢT���6�q�Z����/�A�.YM�W��6Z��UmR�J���Uwi�i#\lL9P�c:d4n�<08��uŸ�r��]wFs�w`���moDl"=9�U���]���pi
�:܏�{'���9;��\rk��.w`�í��\��׊:CGEr%Ԡ��ۧ�>g���ݕ�3� q;Z�+�cr��su=6��7�=������f9��G�ng,��ծέ`�sǛJQ�=f���R^;��c�l`��\���^x�7k����yym���b���;���ǽh��7d�.��۱۞������E�ܶz�/ny�����\�x�fݱE��V�N;�n��7^ٶ3¼���
���S,m1A�ۭ���3�ݶٌn�Mtl��Q�K�<��^7�.���ۃ/<���ᆜ�ۅm\n9yol��l���Vsk�@�:���a���k�[��V[��kďY��G��vRHɣ��TF��jq�v�`%rm�p�����cW4��c�8{3���qd�u���r=^d����7m���h[�J��?�����������0��s����;.��2�A��@Bl��?A
�
V��JI]��$���~}3u��^e�\�b�J�a�������&�:˙~��=��;���Ċ]�{��(��otWG c"�j��N�C��s=�ޯ�)�P�=\��Sd��{�,�}��O�pq�{%߳�ۆ�!�<�z��c*/]�ӧ���Zv���X{b�L�:��7`��죪D�V��Qj��ʽ�o4�cD�����F��������^�$"����~/�uv{S<��'m�]����!_.ݕz��w��Qn	��ܽ�4p��#W���0M9:�r�ߺ�H31<���]y���'Rጇ$𶏒��ݞ�<*�z�1{�Fr�Au��_;�ݨ�!�%S��	�'�mz���Z�\/��w[���\��ӏ:w�8�]���~-	�x�c�
�����[[���ԣlc�'�v�4/��:zn�r� �)�^�x��6h�3p�[n�g�p���nx�c[�����$��,�ɳ��\��k['BL�5�ȷ�8i�^
�B��������/T`wW�kVv�{��������(>'�7A���;5��b��]x{�
߽7��3�@�q�u�w�o}�w��V
U���}k)�p�-����ݳ�Ss����^��^n����\0��s4N�ݽ�^o$G�#n��<�������S{&Y6Vg��'�k�0Q�!�����}=�/���$�hX.Q���Wu�ޫ���:d}�8��yU��W3�w��ꔕ�d�$��9-��L>��}��o�k����7/��D�$�g�d8�����!{��i�x��������O�H�7��{6Ovн;o�ooc������7���D��2�L]*��/z�_��:WC�e>7*�&��f���Ԧ�7{K�V��E͎�Ų�㷓���v�OnvҤiڌӚ�u2j�[�}[�32��]�#�ܒ�К6��>d��.F�E�B�9�n����{t�.ӈ���{��nZOW<�K`՞-s��t����y�;6x5����nFk��9��!�6��LKrg�U���7��pKٸ��׀�$��x�nфS�GC����ڳ���Y���$e��ֵ�]'xq��ݦV�_�@�{o���L#|�09^����2C�����A���j
G�
�$a[tk��7<�x0�u<v�r�����k�z���<��x��gǵ��,��Ǵz&�J��^SJ��M�T�+�+�g;w��{��E���j[CC�\w7FE�F��'a��^ܛ�=�Ż�lr�t��p��.����b##�o�Vx��bɸ�Z���o=c@��e<�:v]�%����[树C�Z�����;��ʾy����p����ϰ�.L�&Y;�+`�l���򜎾a�<vOd�����ɨ�~<�RyVU}�ռ����qA	l�(O�EB���.A6��C�C�����e��~k}.����!@Ԭg1��|߂�4voF�ͬ�[+�Y�}"{2����ҎIitjƋ
�oI�l��wK��5�N�����]9�6��u���ϡ��5.c_e�t�M7�fi^�{�ۑ����7w]���{<�������L[t�Ŝ<���:)J
�c3�+��|�a����uɮņw7R�=Cci�T�8�:t
��#t�(�$�A*�s���i��%g;K���ذ��C'1\jN�>�k6��,���#i�Hk|7u�޷ͧ��YP��k*�w���z]b��{�8Lۏ���r����Nu7Jc�y���:�ߕv�����]aґw5�T���.��N��� M��ޡ+=�v(��ϟV�~�\���Y���/l�ՂOZ��-!	��Pۣ�ȏ\{�um�Y�G1O�7���v�o�������j0��oy����������RY��rv�����$Ξo[��z�������s6�t�S�JK4P���quwѠ��5��ۏ~ꉹ�~�p��I�<�.�ו�	l����m�ލtX�n�c�Ƀu�E`4�E6���P �λ�A��WܠrZ�߼�רVՊ�)籫�)<�g�V��,?mghF"�s�qR3²߹��[�"��ǻ��s�v.5��6�^j ��fivaL��gs۬���y�=�.֛E�e���pSi�{;�'�M���\9^��?m�畷���n�nP��iث��q�8�?!rc��3|}~�m3%r�я�4��}~y���/�A@���<w;�pf^զfռ/V��>�Kj%s���`�s�_����P�/�8�,�圞��e~&���-��>K��̼��;��ŴZ��愚z��v���(k���r�W�.W�8Oj�{�xM�ψ�WoN�o(sg��B¾Ҝh�#�3ݝO����V���L��!``F	�g�7	Xݦ����n]����v�����N�qKI�GO[���ֹ�!)��=�Rv+����+Om�Y�
(<�sapZ��te�wH�i�ln�ۡH�S�����n��S��HG�]��WT��#gܛ4f�ݣL]����u<�gy�y��qz�#��)A{�B8A���[4TO3xA��r���+��oKE�I �0���U�$��U�h���z*x�w�R��mQ���{�+�ܹ��l5�b��mb���V��`�w�#�\M7����zz�V��x@漞��T�#�9��p\���-������a̙�y齟3��Z6���!�M����s��ϩ ���(�<��Ď�K�d)���k�:NB�B3�`^����zڂL�NΗQ����4Zt��Mw�ûv����ݛ��;���p�ewh<¦z�T���]�F-���Șb|�ْ�)��&n��}L ��1�,C�E�IB���ޓj�;�K���:>���*�a�$L��u�%uvUt�3���{|��,0ޝD����)S�%�A�#�Rx7�r��w��������_U��a̫K64ڎo�,���C�5uKŢÙk�9��t+4��u�A��Vz��׽�Hרx�Ј/����p&U��ڞ*��;���/���h��W�6��'�K�KFY#a[&�f���aI!���&≑
�=�(�m��zln�����\��]��=���F����H�¨Wm��J�\�u�k�%�[oMWe�ܕ���� �����z�x-&G�P�K}�(s�{�dN����w��[�&;^�!9㙣Xe�7돎={w��bW����AZk�WY7���$�2��y1�ɾ�a�j�mYkf���u���h[ފHY^���tKՠ̹�~�3
�j]>�_�c���ϫ�;M�e��x� �f�Ճ��+`���[��@�JolɣK�B�u[=�~�i>6���A ��zV�^��v��M��u�dl��|/~��zӬ�IC�M]Cp�ͻ߅PU1F2��-� �Q/`Pg��E���p������Ѫǚ��8_V��~������%+�*f2$�)s��a1Gp�FTa�P�YOi��v��*��.�
Ξ�� �m3])!��8NԒ�_-�i�4."���e6���f������(������ݹ��^�89q;��r��]��Uc鯕c��X��Z��
�5�V��jwx�
�]�S��aɴ�5�m�-X6��]�-��.L#oGs,�j�P��:w�u�ru�n8;���T(��tCsf�`�ᦶ��J��tv7ev�Tvm����S1e�퉣g�T�;j��]^�nAM�Y]J��j�R󬌝�M�\�;�QR���1#��}�ԁ�]#$ov�0`Z�~������{���o�[��w�����J|O���M��~F�����]F�^��z�k��3<�
����Q{��%]\2�@g�p=�Ǘ �fɮn�u*�y!�[+���C`<���b���8��:�74A�:w����C�(*�n�U�m�	����o�����i�����܂* �q$H1Z7��+3qz���p���X&r�=���ߢ}0eD�Eg�#3tK�@���$��_J��)��~�b�I_��]��,t�o��5#N�x��E��{y������%xb@�Q.B/n�����	�/iK�ҨƲ���*��ry�}:�=�<;�;.�c�e�Qͧ!@ʁh���*S\U�=nSɔ�<��8�X׶�vm�ۭ<�3؏c�t��2^�t ۷Gk�3:CV8��n������\c�^|�y2�q���[[auN����rE�_�~��?*����">�t�A˅��ͺ��ӷY/�m>�t��`�̚Oae��ݚ/���n��C�U9͓V�l%ڀ�g^:-n��,.:��B��.��K�z�I�Q`9������{Z�yIh��]m��5��7Co�7�|)��.�{��v��(��� �b��;�Y��;�ubī��ɀ�|l���0���Y_x�\z������3c@��_Wf�=�ɣ����ƋvD�a5�{�E`���J��݈7¥��n���2������N�d�ݿ]
�����Y��L���m>I33w�n�C���"����arWB#�xY\<�����m�߮GV�lxp���9'[�и@c�=���y�t!����|k�;W�a�/��Vu�H;���]�H܄W�j�3{�X4/,�#"��u�,�//[V#z�^��\Ц`��T��vꪎ�M�ǉ6��	���-Y��#�(�[�D�9V��~�z����D�ѥ;���x@k�֌�؛S-���U�6)��>��W�/��4 0�tbe��D9���p#�4s�w��
��P~��/)���P�+T6��1�x�ByL�7Ud������v�J�:�x��W��y�\ ��<u�.�ѫL����А���t��߾�@_��:,���^+��ϼ���W��'\���\����VuX[#b=N����T����O!���G���<��G����ԅH���W���]��kw�\t�ax3bٗ�w�W5��\x�hZ�Ԍql7��Ԯ�S�t�d�P��d��?j��pц덕���~��� ��-n����7��v�ʊ^
@�
J A�����Gv9Z���]��8�Lg��\�9#�Y+F�݅��1��s{z�Y,>�l֩���S�R�Ͽ�|I�8}����7f~��ڕN�9�̈t�_�a����q�S�C�s����
��*vsVV��B/T=����c7Z�p�w�4�^��^v�L�
��5��a8G�L����%�w�>W��^��T|��`�^2_Gw����Ҡ�\f�-Rp�v.�xe�m�З��{V3��"��A�6L�ݷ�Sͮ�o��L���m��t*�M�]�1o+�]M�tV�5y)z���+�.�Sd��	�ݞ�^4،���<�?�V��9~�w�2C�u�th��J�{�0���d2)g�ժ�PU@��F*ۮ��ߙC��*vRK �ԵBQZ��y��z�9��9���õ]�;�'���yڨ6NM���͂:nF<���b0v�Z2��{N��qu�b��2�z7��A��x�h��e6#��4��n���>��|}���!�V%�ʱ��zLaH��"�%9�S���[2�7R]���2��)LY��4�ݤx�t�w���y�ms����c��rG3��RF�(1��`w~��*�cr.��O_�_f7V#��I6�E���Y�ޮ�)^�S���t�ܷ)WKM�Ճ�UZ�#�*���a��I���F��Xq�r����Y(Ԃ����+����7�5R{�:��̥��Mf�=�����
/vu��l��M���u(�sjk���y�C�t�́��rg�X8��u�+*8*w�u�#q��:w�h�x���(�|2��C#�g�d�z.��;�E��wwA8�Y��ƭ(�$R�C�R�0���ݺ���ѾS�ź��*nrJ���$���e�Ȭ�4ˌ;n�N�5���-h�$4���͗o���vu�W�%�ܧY9�A�x��ՠ�����<eyWg�ڲ����k�Q�HJYy���i���H�4�,(v{<55��l~�_�Zc˲�:x���;}�&���$�#�h��-�V�F�B��c>�(�q���(��zz��=������Ϯ:���l�[����V�K_M�����,�J��z�Iȵ+���j!�	���q���A{���I����W(�H�;CUx^��N�$�@{V2f{��*�fM�oə-m�wS��v
�a���n�[~Ϗ��k�<�^�F���:�2�����n
��T�+N�"rP^���X��V*f�b�oXҴa�F}<�k��׫n��d͋kdʶ��l�e��Y��ow1�E�J�ɴD�3^��XrJ�6P��A
U	M���H�������!�{�*��]�����Fm`rjZ�]���{�MVěə/��u�J�*q�
�6n�6hL�ko�g[A�����"Ap}�������o,aW�]��$�qv��m���x�e�#�ON�0�KA��y4��
k��Dku��F��,�v����}�������^���{��ힽw�RoNe�G�F�J�}���{��&W��d�i�p�]�ճ�\�B	�	g�Y�^��veObQ]���c�s�����"��`��\k��B��}�;�}����=wӜo���!��NƘ�k�j٬��Ax*4}Z��4��=���'�0񄂀ɫ	��T��KyV̎b��󜺼K6�.�}wh�UJ{F�9:a�ETB^
�1=�u�`�BҬ�Ґ�������0��p���9�I�s��y7��ɱWL�<�b8�)�IkrQ�;F�v�Uj��\�m\*<1Z�}l��km�;���Ny���K�
�ĳ��G�������>~��$��=�&Z��WJ4"��lxyL��vL<��ٯ���!��3`^B�����.��`Z�%ֵu3�|�Z����??XM���mtA�7]Vi�)�����N��k�8֊/�]�2G���r��@]�\ԥT���׹YU\J��^�N5?c�O��i�_r����JժX���Kl��֍�xP;��*��w�cL�L���ڦM�9%uwyVĎ8K���z�����n���J��\Y���yV^�$�h˪W/=�f�S���K�E����c�冴��%�t��-N�x��ӹ��u��۷k�����/,V
�7||�K�r���[j�I�MV���ѻF��F�Fj���v�g�5�P���uT�z��I�l�w�N�ޞ�8�2��h�R��eeWV����J5D<���+������}O����z�������J���B�*ZQ#u3v�w�g'�H��o�:n�{��VM���oS}����ݢ;�Zw�V��4��B���IG���	v�[@e俞v�a���(���p9���ʚ�J�}Rq��*�<�:*�"Tܧ���~�6���sF�7b��P��+{H'o*-�ʆլ�����[�rs�nk����B�4N�t!޻{�Ӆ�f��xqR�j��W:>�E�v+ε�^{�p�(<�S����� ��9G@{d�sM��э��;:N �K�U�U����3`��mؑ�:.ګ������hݷC�o�j�k�[k��X��f�n�ݓ��G���L�Ź��;��X�������J��&��)ֹ4�n�.m��k;���7Wk�r�6�w`쵝���"�'r�1ʈ�aX�n�w ���a(;t�}����ѻC�!�8ˇCM�uɧ)�����p��>^���`�;���FCx��q���붻ͨ6��c�yx�����������|��=�n���/F�y6��l]7m��nW��.���sͮX^m^oP��z׷�"�m�J��޶�^Cl�R��d�#�.7o���mb^Ʀ�GNd��A;A��g��9�F�\@�p��8{���vy��\��x���m����F�Pg!��wRb�lt<�kd����y�z�}wcp��κ�\�m�7�k����k�|�� ���ݞ݌bv�Z-��ݞ�gr�Bu�i�X��㋓C�ǍY-� ]�����{[�Ǧ��.����[��uϷ�]���Q���������������jҼ"�Ħ�n��w�����./�I��t0
h�D��$�H�%7;gpڹ}b�7�+yų��y
�A�r�	��KU�۩�'���0��{>v���b��QH�T�2�Z7-����Nv�f�f|����'���V��(��ը5�g*��8{o�=�k�;/�([��N9$��<�:���A�s<�J���߆Y�U��>�L�0#[ѝ��|�Ft�j\oG��tp����]"�������nmۂ-sƕ7T7Z�Ì�*��LE}��j|0s,����2��Y�k'5.�uf��x�s�Ӽ�$D���uV�z���A+�'>w���a����CA���ɸ�<
�(;#vG��WW��.�ٽ7y�[�K�i�"B��V�ɺ��>`ꋎ�a��ָ�n��U+; ��Òb�fwI��eg��ڙ�{�� �X�A�p�+"�������"��D�����]׫��6���M�V�����T�%!�9�g���Ri���2Hz�v�vʝ�S���J+>N�Ț����c�����^뗨ܽ���w��;�=B��'���.�eb���s�C1�	���X�s7����U�f���Mg�ʙ����p1}�ѳ�S
�g�OXU�kN�����x#/e��a�L�E�cG-ר���`���>��T�Y�j�j?D�

>�q�M>�l:]Vl]���p�	_}���g�	X��X�4T�XH�-e�v�&U,'yʙ'�:OoGii��30�R��Q��vWj�zڝ�&��Q沊��w)ȯu'�&�'�D"�Raz*ߥ��������b��*�ީ�:���|�$uw�;}6oq�\�;���%rл��Z��u��yÌu�9��
8U��R�w�w;���.�nV��@����!T�m�{0��םkv���pc��]�L;���Thn`1�9�q�%δ�ku��Q���N�sz��H䋺��KË۱�l����z�/�5���Eŵ�";(j�v�d����������9ÛK�m�X�$J+��9f�n!je��[@�U��UA'����Ϟ�"� kv�,f�J
�KKQs�p����cmi��#����j���M�Y��i��݀j��\Z͈�@�4��5�-�gT9��ۂ����#_~�s+�Wi�ht!��+ӷ������C�^����|b�A��,H�pH1�U�k�uM��Գ��;p�*��4�:V�Oz��ԍ���3-1lGZW4�Q���H%n��p�۽���\},���j�i����rGJ��d�u����>�0!���S�v��f�������H뵊��(��PĐ&a�&�p�W�:���=ݛ���+Fn$(N{պz#q�V����+�=X�g -h�&>;�o����U�YTu�-���M֤+��ec��R�G\�n�S��A�j��BN4���AmN�IL6o�k��9���at�ǵ")XF�Xr9a�����Y��k��g���@|�M.&�]�o���4�b���p�20S�2�`�r72�h�q��2�������{]�~�+�S�˕�V0�u���e+&�ڽ���lL�v����<t#ʂݝևu�����!���z�鴬,I��2�d*����6+�٢�v�&7@b�V6�hd|�"��uD���h�:���w���:���"�(ݡ�*�1�R�]G������nu��Y�?g\�ڱ��rn��i���4�mZ��o�208��BՁ����=x��{:r�&�g��9*ح������=�c��Çt=wIj�R�꩖j��V�%�̙�+9Μ;Fm� ���]�*Sup��=-��������m-|0�>hCB�[b�k��*�W_DB�}ո�����9G!2�t_]�P�WB��̗@�Ǯ��k#�M�U��i��q�FĽ��n m6z�^���ܧ��4w'�n�%,Yf���sn�{�D���<��%�n�ξ�Z�%
��m�ځF��2����ۼ����jQ��9hۍ���tm:�]-ՔTY�YA�罫\�W��� ��s/՞At�N�]�SE�]G����[JnƔН��T{�u�ǝ�}��<��M`�KǐӴ+���лU�
��ίQ��s	��{��T�;չz�]�Δ'ie�j4�"ApC�r���E68�㵠v.Ŏ �j�5w���˩�K��Չm`�r���ڮfwj���n��v��'mb�c����͋]ؠvv,��r�U$1�4"H5,AT�ua��O;�^�7���G��qki�Fh�MpZ��ه�����%�F%5��z-p�UZ�bT[�X�)#�����&1�1��F�Z�q���m�y��;�V�@��-��A@�4�S��ιo:�������mGR(h�;�]<��Qyࣉ�wwF������β��n�3�㫼��+���iK��OC*Ue퇽�gA��ߓ��5�����'}'T!�̑d���:-5H��������H0Af7u�=A�p�Ϥ�p�Y4��]�=Vt�\"��Um�%�i�@�l2����r�6��beV�R��s�{��=jɚ�����sy���s�8q���{5���ee8G���S㙙6͝�*��K�ߧXg�)�aK݇��2ݱ�� �޲����ug�9����B(�:1�l�{7kuI�U%{Քqc.�+��",tζw5IWC�/6�Z16*|�����rZd�ШM�yLolR� �Sn'�l tr�&.�3��&���߭�6���vv���ݷ]X�Wi���I�rM��ƭ�ݗ��%,�PQ���:��F���e�����Ty��`����]�H�{��ew:�.�PZ��ʵX%��щ��#/⍞�*�
Auw{q�Z14���Z�w4'�h������x΄�uN��p��N��oV�AI#�ꡫ�wF�*ы\\��c`�A�g͵,)$I��p.�84�n�F��[oe��R��M�u
��Za72����Nvz\ʼ��a�X2��ɻN�g3�3��UǏm��e�_nQ]�w��i1���Q�Z����e��7���e�H�ч���6Xљ�L�Ue�Ʒ[�j̋�A��\��ª��m��Z��ثD�_!�n���]�[��j�1�*�+^�99��iu�7�����6�}�ʸb9*�	�3������E�tH�F��8�)�5�6��"=8e����쭻X�Mص����K��k�i{��m�����*٭�X�j��nV\/���BF�otg�2gS�_aˤU%C�E�,�[x�[�Ҳ�)��b�>�ԏiY��2���%�ח"t�<�ӳS=yi<�7�c'�i������,�Z���HM������$��k�����õY��gqN�hZ\+���!8{���:�z�a�e��}Dk��
�/q���g��LT��c����ػ�^��FK,���U�o�VC��6e��&咽�TOTFu]�$~����7Ъ�[vN�~&d�4n��ya�T�ŋ���4ŵ	�����ʭ'p��>��;���];����(6Ƿ��O��1Tr�^X��8[s��/hn�A������;�3�KŔ#��V��G].!8+k	���- ����oHD��<cOuo=em]h��#�GV}��V�2��d�3'u�z����͊n\S_�/���;Q
3�a�KD����h�m*C�r�ݽ��K�Ϲ�"�ɀ����)�n�1�ujM�ks����[��f�rc;��l�Z�p��nO�T�ƌ�j���/��k����������]mt�k��}�E�pD�2�W��K��]�Y��l,�3�d�6U��tͼ�2�iF��s�-v�c/)�ێ2�YE���GnгI�X��ݗGeB�HوW4ƵӹЎ���!W�-�^�E�X o`�j��a<6�kb��9�bv*���ِ*
�uu�ޔ�S��:���U��z�V���M�&��M�u
�W��-��3p�ی�/s)�%b�S��]`���nի�p��X��M�\��Q�^^qK}��6m��1��7;��ݫ�W0�X��N�6
�]ymhSҪ�nQ���Z����j�q6�Q�C����RH$�F���>��L���\�MPNnU�{��	��貐�t�(E�ArL����MK1K���s�Y��$�-�pR��k���n���n�q�e��:�`�r�t�L�����Y���.��Zb�m��ƵIq�3���Ɍ.�t��wwڸ��v��u�6�Y� JG�Q�R�!�җ}���A^kK�PeUm�*�Y2����aD�7�s3bE�م���a�ش	TDW:�b;"ĦgЊ�L{z[�b��%�ۨ�7,�������ۙ�<��ʝ��	�QTuȷ��g���;NKn�;���=�%�������(B��N���"p���y�8)F���BXc1��W��u�F�Wu�y�o��kr��lxoo�J<9����5�S��S�����2���]���2�H�E�/Apq���ϯ����]��U�z��B�lк������Y��dh'�}}uǩ�ِ�)`�3wr��uV�d�M����ݟe�C�G���}�����\�����f���;�;� ���hk�Z�y�w� ����(�W��DI
(���uu���3sTy{�[��,܃@��F���D�e�o�q�Թ�9��x�k9[{(�ÇpTڣ.��G��3��X�]��p����7�u�w����]�S��)K�W�.E�Q[#���>r��l�
��U�v�ި�g�-Ą�v���ov��M�{��h*���%Eϊ�[b�.c����%ot�RIX��M̂�q `�X$դa��f*:H��v�8�A�K��`{K��b�U������e�
Nv8���/���9�sݲ� ����|���gc漝]Bc�b��E��]mǑ1�w/d�n���Y��f�vq��\��n��p,X]m��t$m�z��G���!8�9x̡���Dj�hv�uw�o���&�e($tcÕĽ�\,aը�*R��;5��VƲ������Jk���=�\`z$n7j��|�أq��l�
�c�$�P���4!0�8�
��uģ&L*Mb�:�:�D�ѴM�0A���A��7y�X#�aЭ��h$�e��Ռ��iA{�k��Tު��)�Xyݢp�ƚ��)�vx�RF�5X�.]8�Ώ����Н�sv�'.��� �T���wY!���كR�9ج�+��C_��<��j�5s��w�W��#{#*�1�w����rSKy�o*�o������Cᒐ9NI��R�O�,��0@�os4����m�lGV��`�l��+CM(��1mǌ��j;�q>��/ =��1O�pwc8��@��]����7Z��$	>-�ͤ��h��I���"�pe��u��lwN�.��-��@.��FSڜ�2�Z�	��:����l�o6���`�v���N#q?qk�~f��*�xB6F���m&!�7	�=�O�\Z6+��)��歍:2Q0���x�>P���]��]��4�8^�c�t�ԥ��a��m3�L�v�_D{'�P�R��XUM�דp)�e�.�1<�"���3��`7�$��|M]lP&H[�窫�yI^�ˋms�8Q�py�-w�����I�-�0G�Q�܍��lB���L���{�v��&�'3���'i�/{K���$L�V��_��?_��d�<1W:�Ϟ.�����A��7Z3vb�4w.xz�X�Yz�mg6��2�����gt�%"�u�Wm�d)?��$���gZ���:�v��H��H0��2�E��{#}�n<r�i��n[�I%�eX��X��b�o�gU�L�+�7�u�]�4ю���٘�0k�WVh�����{�;/��}o�!-;�4�ȕ����9n��p��/s[�]�z�3mE�8��Fڲ��a%�S�8䏼��\6�j[�#{�X�����n0l�S:��˒�(�r|ȏ(�ՉV2%^Xtb��d�,O��:�����Ņݴh��,\��C4����C��;;n������V��L�nT4���vUvW,z&�d�cc���ۚ]��}]4V�J�+v�֗=���w=\�9�wJ-A�Lv˷�̽���W����cu<�n;zbܣ��kimw)�����t�h�F���DLV �B�4���6�5u�1��:��G�Z�a(10�!@�'gz�,�V K44���IV����xɊ�*J���uؖ�Gut�6���N7����
���諣�V/]ݼ�N�����*�{r��fhz����\ӡ�ھ�H�A.�kr��H-ҒuE&J˪��Yj*NMÑoq�ɳ�6V�W���ɛ�~U�pd�T���+)�����c{n��<̉a2W*aA���p����=����b¾���z��AZX^s3��,�����H���bb�ͯ��5)��mqϏ��=+��
.u(L;Q�[����Ezs3]	�X6Q�b�e�Z�7fֻ4*J0"::�,��2�`���+	�^�̕���|VfH��<�UN_Y8�N�v�u���*��U�w0Ҩ2���l(�Qt��ggs��f�Y���)n���]bP�6���������*�f�&)H<�;x�Y��Ê*��!�NJ#���եt�Ⱥ�Q�V��;��˺ngB��|]��E����ޏO\���b�.</
�1B5aOq����[���L{���V�5���f?��U�b�]5�
��bBH�泗�v |�u�J���efho���F�D=W4웡�.���7�^��WJ��H�k���8�z���v�ڒ�GCJ��W]N��
v�"eZ�
b�E�M'mݻY��n�pe�*9�/��J��q�K���70�u��}�pU=�C��u�b�P#:�ܼ�;���{8"9�����X�ٳ�N;'g���m�t�t����nx8�]t�6n��v������g���f�<�-��J�O7k\j^;{&_d�o6�u���N;�{v7���`�;������Ί3��-������۝��{l�.��7<��X3��ͱ�G���Ln�h�&-[V���kvK�����v��ۭn�!,u��Anz��6nҍ�G���s�5k"w��Ts�Մ������֖��v�щ����G�&yE� i�۲�j�v�{R�^2Y��m:6����]�;���azO>�1��x�u)����F���n�#=�3�gs��3�X!���qv㸴��뚸�V������n�Y�ya서T�6�F��ڭ]t�v�#�+��1�&��ƬB�w^ݍ��Eˣ��ܮ�zy��ˮ9��(�J��E��8�v�t��xo� (�`P�߿��?w�ζ��4,�aQ˺�T]�:�7˩���R&~(�Q��F�ڴ%0j'l7��Ё�6��HF^�}V����r!J�Z���+���B���-w�2���쩻K�a�h�e��,pO���i�JÐ���,�ށ�cĥ+�}V8�%�Mǹ�����6���ibF�eID7�30�(傩bn�GB�Y��p�}vE�m�b��W$R�gf]��p�Z���&����77<�5�<޵4������jǔ�J��7��U��K���s3w;iɚg��L�ͤB�z��}6���@k澡S*��]=K7fXɅP�jV���J�6H�L�"lΗSo���S톍��^<�:I;=Я	��;�×P*ۮ}ip��CdJ�����[��Pl9�K��K.4���C5���N�μ��v���j��9�2��3y�
MWT��x�ߎD�!�G�
ˊ�/�E�"���n6�ؑ ��Z�� ����Z�\��B�0j�d*���d�\%]�}�$��9�х���4�نÕt6�X�0^��rۮ��E�є�b�1W3]�9��'i�C��V��s�e�Ժw[���'��m�3z�;³sVJ�`���ck{LGr�サ�����nU����������d�Wk[L���.�Z&�jA��8��v��\$O���\��ߓ�Vm��c���tGv۞ךฆ�0(����Htj�kf+7m�n������n���+�E*`%ٻ(-gY}�D�������z����M��N�I��֗f끂۾\��+w�^<��@����A���
�A���7���}�>47�/(>t�33B�����z�ڇ���h�;M3�݌*5�����r��v_�����v6;1�غ�"���5����{vۣ�mi��N2m�lk��F��gmߍ���h�������#�R]��pm@�F����]�󭅻mn���+Ycb�Ƨ������������k�9b�h�4������ՋL��\%ȽH8墅G���>f1-��s�q{u�;�MQ%%{!�hdYܬ�lݪ'��t;��	�l����ҫ������[�V������i��t,�#��:r�B��Th��朒� yD1�Xm�%HzP��B��Kʈ�޿�k[>���-�<�ɞzO&�X\�+��y�$�����{��2�KO��u6���^S�a�%e��!Rd�h�W�yaDW%�%�ӈ�W;D��!Iaev�5GE7Y�osp$�əy�DKL�E��vp��;)l�&m��{�Jv=}�����U�`����xd�X[J�O�}t���zZƟ���]�^D��	[�f���\(��%�q4���[`�*2f6��N�k�o�]l5R'yC�3�˥��¦�_{�N�Ȃ��@+5��_���.��K�j挘��0�4�B9��%E�غ�W����1��EH��R��]�:L�9i��c�|`y�;�|>���3�RG/�V���<���U�U��G
�QE�Aq5��D���]�����Ӗl�R���Ο�{���X�׶���J>�:G�%k��c#���:=��i�v�-�4||g%yw��,���^�X&��y��`�z1��e��[$(�f�8x�����<\@��w]j{�t<���5X-�x=�/� ��s���&����X��F/׼��{dn	M7Erx�xJ.� �L7���9b���X�&��w�dt=��z�q`�/���^<l��g��V$6���4f��~~uD���k��	z��av��l�V# ������l_'�����	�FMb�x�=����ٜ��D�Y\hgh�7�qT:��0�g*�T=�{Q�yT/|�Iza���C"��s:��yp-�"��/��L{:�9�U������F�ё^��f4�خ�B9mA"w<��Y�b��r��nu�Mp���.�(�*Y��&Y��r_���cm"o���~&�=�����P�!j�&K¶���(>q�E{�}�ʊ	���ެ�Y��_I�R���]^q��n�;[Φǘ����2���t�#���h��V{�5����d�� �~��e���̖F�bNtmi����@A���uE��lw�1�TOV[�T�Q_b���s�u否h��~@����Q�:l����|�&eߚc��W��k�������C�j%�Ȉ �Q Ng���I��m��mz��B"v�k>д��Րz��{�s�R(���$���W�w��\@�O3Õ���XX�Pu�OD(��jX��Y��8�a(�55ٷ@��0�X/RB�b��{| {iaصk���q��%2�Z���S�T�^�?]]x~�T?i�yj�
������;�M4��ˡ)Pw׬����A+%߻8�Vlκ��.��wf��'sф��DR�m[gn�Oq��Ń�{okl�Sq��cw[��s�ȕ9&�yv�k\��q-2��:�خq�,r�#cg�<�����d���]y�`���J)��y�E��QgG@:�,��_	�=��1�kG�U�aEZ�wK>�`�Yt=�!���aGy�١�P���vW��Q�){Z�Ύ���E�%����X�e��4Lh�����Þ�㖴��h	S&�f�.�׵x��7�?�K��?���i���}�� ��`��:zX��S�8t��v=�8O���qY�OuԾ��T�V�Y��[�Ǯ���U;��̡�@~���s7ލ�Ry櫼�F��u�͊i�f���"��.À�v�|����͙3���Yq��ʴX�W0�O'�����N+�y�/)J�Ǽ�f_	�\a?!f_���7�P�K���uK�k-���bx$���W��}a	�^�wcC"�-�_r���ۭL��W��%ݮn���S�m��gh��v�m	���49/��mG�u#'����%���q��ߝМc2��`�XQ[��z�:�N-�
Ж���Ε��Nr�|ېPk�w2��H���R�=��z�Q���;�_&����\Һ�݌�(NPV�L/P�nwxP����P�/�v�~�{�V²<Msz/|����pI�����ś�N���3SA�J�8t�l{YZ/z�&*�#K{|���9�:T��M�6�7n$XlF���n9�b��(�����?w���?=����9i�ق���5{���yC�a�o/���uyѣ�~c��[�m���v��yNgk�=�B����=��>c��i��������<Z�U���*�ȏ�I��C|�h�È�`��Y�<V/_�Ғ#��/5���.�xt��+p&y�r���L���\/�J�1sEX1ftx��R��רT�(��N�,�����J��rP�9�Q��ҳ����z�"���ϊ�Nw�pH�y�-��
��ΰR��}P�/�7*�<s���{�xy?.kn!��=�8�@G�`�*"F��T��2*ǋj�j&4��U�����V���p T1�(��a�+�פLUW��Ϲq�G�ߺV ?f4�z6Ikf���%0�YzڕkS���&�` � 1,Ői��*B��$���V�Otyk"W�ߴoF� U�����P�h��dA>Xž62�ZKM3�I��i�D
l���-$�6��y�JPtd���ۇ-�~����rk��>�o�<��##l��K��|k���5o��08+��m��	J�\|���=W�=��X�JR��W�L�ߞ�˻����Zc:c��z\���=1w{J��>y��11M7�B;W��\TԶ/'����k��o�����:v��c|��̳���Up��^�缉ZSUJ�	+\��k�xeJ�FײLX�莽u��������<QJ�R�����ò�t�j��(鎧�:uW��6�G������[L�ל�)AߎgM|v������3��֔�7S��w�3�����Ǧ���q�ފPsv�|{c2>^��=ǌo_�<\%�QPz#���_u�S�M�#�i�D������GSP�K�EEA�u�cQ�K��:xT#^��ۆ��)��km��4��w=�'͹)A��������"���#��u��?~'�z	���|�i����^ڞ����'����{H�~���v�ϟ������'8�.��7.��X��c�v��=A������OW���IǶh�PvK��o�N}&i�zz�#�>�>������M�qN̫J�a^Ư����}��J�wQ���������4����d���b�q�7�b�H�
[Զ 