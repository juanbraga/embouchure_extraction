BZh91AY&SY�c8n�߀pp���2� ����aw��      �@��    )JP(��                                            �          =@   � �   t� � E�  � �@1)F6P�FEV  �6�,cT,l�&,
� �,���*\�f�]�
�          �jZ�!��q��f�l�gZ�� S6�X�#�X�P�  � 1 ���8�@� �S���1 ��� ��X�ti�;�Ur�*�          j�AX�@́E�2�� 7q��.����sk��Uc�` ��'.��J���T�m(� �f������ŀV]WZ�  L�!25ֵ�iN�;u��          u:�q�����+��lWWJ�  �tr;��#@1h�Y�`\ ۅ.1��:�hP���F� uR�\����q�ā� ;��Nl�A��:i�лì0          �q�5fQ�v�mN!�L �ULmJ,�J�҃ �X )��LM*,��U]8 �siq��Yj�ۈ�Z� wZ��n�q���v�9j�O  ��d&�UA� �� T�	'��UP4F�A��        O�j�T��Rh�  h�*%M�$�2OS@�z���MH�f�UM�@�d�@i�8�tΩ�9Ni�;g|�Ç8k�n���)8�4B!	��H! �! ��� BA\�A	�ҏBA���DH>L��]'|w�2�Ĩ-2Zķ,
QDR�b�A�S ���E�))�Q�����0AXSC"$Y)�1T���Ab�1dT�
AH-2�)U��P%F��(A�$AU ���Q(� #�� 1���� H"#b�
�E�)!I""ƁT
`�2�S�RA`�(�EX� �"DJ��R
AhX5UURE�,b�@F1"�)�E ���Ab���VT���QbĠ ���Y �QH) �R4���
PTQ���dQ%1hXĉ"P)
H(1���
�Y��R
,X�$R
AH*����R�R
AH) � ���H���T ,H��H(,A�2H
�F*��`#DAE��
�"�$�$ đ����UDdP D,�X�HH�11�(B�`���`�*�b�E#E"�R
,�QE ��*�*���AH(��Ă
*�H) �E#�H("b,`�"���"�
B��QdR,�$��REX�FF"�+E���H�dQ
A`1����R
E��UT$D��Q
*���$$(@��SL� �)$
�M*��E�X("�$�$��R
AH)%F�
A��$��R
AH) � ���R
AH) � ���R
AH) � ���R
AH) � �2�%%$��R
A
AH) ��aI � ���R
AH) � ���R
AH,�(
�$D��R
AH)�M$���(��R
AH)%2�
AH"AH) ���PH)H) �P�%%$��R
AR�R)%$,*�H(�AH)H) ���R
AH)H) ���R
AH)H) ��RAH) ��$��XP�H) ��I � ��) ���R
AH"AH) ���R
AH"AH,
�$@�HF\�Qj-E��K��"� �R)PY��R
AH)H) ���R����D��R
AH)%2�
AH"AH) ���R
AH"AH) �����$�����XʋQj-E��b�S%$�$��R

AH) � ���R
AH- S)%	 ���R
AH) � �RJH) ���D��R
AH�T���AH)D��2A�
�-�B�-ImR�"�EH)
HUJE"�%1H*���+�T��dH,�RRI+DR
�X�"��%(,dX���b(�X)TY ,"�-H�dZ�Qj*��Z��R
AH) � �@���%E� ��$��R
AH) ��$��R
AH(*� � ���R
AH) � �@2����YQ
H) ���D��R
AH) ���D��IM
H) ������"SH�R
Aj$���R�R
AH,R) ���D��R
AH) ���D��R
AH) �*��K *���b�L��R
AH)H) ����BQ��R
AH) � ���R
AH) �*"(*�!L)�"�AH) ��$��R
AH) ��$��T)������YI) ��$��R
AH) ��$��R
AH) ��$��R
B�(��"�AU$�$(H)������R
AH)H) ���R�R
B��RJiR
AH) ��$(HRAH,R���$QaH��i�)�����) �
HRAHRAHUQ
H,��R
B��R�R
AH) ���R�R
2�iHRAHUb-FTeFTZ�Q���eQX"���R
AH)!UD��R
AH)��Ȣ���
AH) ���R
B��) ���R
AH+���H) ���RTAH) ���R
AHUQ ���QdF�R
B��RAH) ���R
A
AH) ���0��) ��� H�T"BRL�KS �IDUDJdP�1-�jKIl�%�"FR�b������ �)�H"(
E���F@b �&HK`�D2̣
2�j)����I�CQX
Ab�T¢�)�T@�
ȋ���)lZS,1S.��(i�� Q�0�%�@E$P�RQKT�Q���)�%b��S"ؖȑ�e�%$FB��2J��P
H5P) �1X#E�RU�IMDR�CUJ42�� �*�VM	��)Jh!
�`(���J�II ))
HRAHS"%2
JA�l���b�L̒�X\�KIb1B�%(
����0���J�TZ���) �AH(RĦ�2#"FAUF���̆TZ1��dL�s$�,�YLS,������E�)��Pj�d���RS) �R*4�����%2R5U�JDJJ)
d�����R�R
B��)
U)+��4G��v��e�������m��SM��j�-Ԕ���  c �v��n���ة���V�)�r��p��]�
��Vݫ�(��{� ����6�@      �       �oˀm�eP7�'*� cm�����͕ݾ��{]��@ 8@
�    U
�;�[=T     �  7     m�y��-�M�( �;���8F3�� ��X�< ���p�OY�������` < �P�1�p�� ی�@v�w�l��	��8@x x8  ' c ����<��{  ���s�5U�۴w-���7��ʣ]]�y����v�U�ݞs�Κ�m+�ת�lwn[ ���綶��j�T�y�pκjp0j���x==�����	��8@x x8  ' c ��@�1�p�� �p0*�T�8�;o7 c ����a��� y��(cN ��  Nc�c ����`!�  ��   ����� �����q���򝰇��p0  N �����6x�=�����+�<��0 9�pV��]�/9�0_���+���\[.0����Ve��1� *��	��8@x ��	���ϐ  N ���y�k��8@x x8 �8  ' c ��� '�<� c��8@x��	��8@x�`? '
�y����	��}A�;���[):�A���' c �6�O]��y�p���^��N�=݌����]�z`< < �-��˼Nw ø����^���P �m�    �ZJ� Z*���  7x� �M�� ����ld Wslm���qwU��P =m���` <�	�U���ys.Z޿f�1B�"�A�����m
���  @ ����   � s�Tu�Y�1�aW�� ol�c*�   �  
̢��P �@ ')�o�             � ���mݴ���Mܷn�  .c�m� *��U ����+�Qٞ���1�r�m�| � Ǫ�W��W�)�����*��]��z�Cl��wR�ea�ݶu< �T1��PT�<�IǗ3:��Op�7c�@��<u��B�@    ��T�hw6��   J�`   �     *�      U    Mրn�� ��6�i��7<�@     l��   YATp w]�  T  �l@T `    U 	Ͱ      
��  ;��d�  �T*�-���  P=���ڷ5  �Al�     *�` �P ��� m� T*�   �  � �    l��o`� �   VP  >>��     
�����*����W���mޓ���Μ�ͺ�ܼ;ͧ+ب *�  VP  <�U�P .�Wv�J����'��{��璽	�Ǌ +���yq]��f2U UU�7�{��oo�Y���8x� 2@ 
��  	�wT��Z���g���RͰ    :�z�����<���*�o���?=7w�s���Lةn�qܞ�v�́۵J��[{y�w��9�_�jlq��Wu�x�Zz�C��  l  ��w �1��e`8:������j�9{{��l��m�p0�q����   �z�    l �   `��  <    6r�  T�@*� ݀  ��>6��v@                               �;���ʩĪ*�         >�    �                                                     6� 
�           ��s                          *��m        ;�   U       T             *�      ��  ��  U   �  �  �                                T       �  �   T      �                        T                      l P U �
�                            U          |             P �   �*�*�    ` �U        
�                �T         �      
�             w            6�J�   
��m�00   UAT
��������                  U  m؀                       x                   w   p                ��   �    6��    �         �                            T����J�      ���     p                      k�@VP                     �-����       ���                           wp      
�� �                   -�             �k� �   T@         @                 ��    ��                ��                   U �                        �                            �U                          *����}�                *�    ��*� l  �   R�@              f� *�  U *�  T U U�    ��                 �S���� T  U    6�6(*��            *�          >����� ��uP              PP     5H@T���p����N�r� � ���U�ҍ�  �            
�       Q� � lomm�����\P�U8@  ��� � -��N ����	��;�T��p � �     �6�` < < ����P�TNՠ ��"p6���p [;�������$u��HBA���˟��	�O'�O�ӚI���ϷK��ݚ�k��뙮�Gk<m�ٽݣ�y�  ����m�� �   h�h�v7��z�۰���OT��v�;�ԙ��m��,y��0���	��8Gpsp⨜��'��P co ' S��f��z=��ۧD�'<U�1�p�� ��n	��'g'��m����t�I�ߝ�Y�ն*�U�厀��Z����l� .-�����s ��  �^�+2��kb�����s��c�Ye&��͐AT   �*��K@/TSlU6� �m *����l��  @U  �B�*��:���S����y9�w#Ӟ;��v�9�:�ov�=��=�^u�=z�F� *�*�k�l�����w�S��x���      W0 *�T�         T  �         *�   T �      *�*���          ��     
� �  SlT     � �   �   Tm�=�   �    �   �   �  
�       VP��    �    �� U     
� �   
� lT*�    ��  �        P          �  PEPP  �  @U   d 
�    
�*�   
�h��k�
� 
�Jcw 1�� <6�ڲ�T��T�U�{������?�7����U�t.�Se��U�P� �
�r��꠵ҩ�6�qk�n���ݛlV�ZTm���n\�r�<�J�ql��m�մ�D���\�.�v���� �[  UU  [h � � GuPP��*���mP �6  UmT��� @ *�TU`�[ ysz�� /~���NA�m��A�I)�D��	4+m��WuUm�Vڪ�UUm���i&	`���I���2as��C�o�{�0�8~�Bit��nHF�t���m��g��|V�/��,$�$ۊ�r�E>;�_�8)4��.�)��),8f�i�#nG�%�|<m���m�a(�W��Λ�-�5�}���B���H{e���pz3-�Km� e���P����r�4�6ƽ�"���H�>Yo�"�i���i'$mƒQ��YL�����G)dS�%�#���O���B�mT����4�H��|�i�m9.n[.*��W{�l�r m�lUZ�e�ATz�-Kw5,�9��}ߩ��ޏ)���h�t��8E�A�
G�}VF8E>?a$Z��6�m�����>3R��j�����<v��ڇ���o�|�R<iϐ���)�J��$l&�"�i�`��)�B���~��,�|wD�@�R<i����)��O� �P��m�Aa��Ƒ�ۑ�P�)��_�R��!�y�E8i�>��鸅#�>��˄��G$�$@���奘)��>5�lRͨ|F���S�H��c�
�<E>7*?�A�c� �2#jI��gS��^� ��PxU*���
�U�g-xLl�B[l�Če#Ɵ���FE0��7�YO�
G�M�#��)�%����O�V[��#I��HIp!L6��%�4�H��F��0�~;��G��i��h�b�Np�>���*'$���m��S�B��nD0�|nZY��>3�^F�,ڇ�l�ye>4�6?2ZIF�rI��c�+P����g�e#Ɵ�����L4���o�S�T���dr�E>;g�.��rH�m�܁��x���]S���%�4�H��m�ͫ�~;��G��i��-o�v��{�om�5vml٪Ԁ�� �e*�� �P ����H�JH�L6�"�4��鸩���L"���`�CO��ב�K6����
�l&$�ĉQ���)�x�1�j��O�߆|�R<i��-�dS>#p[���|sQB�r	#d�#l&�r�E>7D�@�R<i����)���@����G�nFi�>*� � j9$&6�m��Hf����8t�eM4�0}r i�i�ܢ�Hf������q�$m���AK:|G�}VS�H��c�
�#N��+H��-�0��i��Q^R'$��ym�ܛe<v����b��@
�l*��*��-N���*�I�,�Ƒ��}��{��e�:DqM4�>:�&mƒP�܌�i��߽R��hx�p��(��i`��@���sr�!aƠnI#n(�C4��J�PRΟ��U���<v���Ӈ����R<i��Ĉ8�q(ڑF�ç�|0m��|i7�������~�)4�]S�#�M��m%�RI$��g)�|D�f�F�����!�|F�����"��馑��W��2I�HY.���|8m���g�С8����x�'
�  m����Wv��'b�mk���nǭ���� + ���Y;�s��۴�w��G��ݼ�vV@@   P    ʠ r�*��gp*���T*��6� U w �U b� �  ���R�m��U-���*��*�ӹ��]�^��m�ӽ�c������3����x�dڨe*��m��#I6�DE>2��)��>J�PRΟ��U���<i�z	N����A��ҒI#	�G�?n()�O��`����>:o�9����tK�H�x�1�)D䐖�0��>"i��i������z<�3|���f��{XM�r8�Q�-l����4�4��Z\�i�"�)äx������I1�TNIM�p� �ap��X�G�?nFE0��|��H����F�}�o�����m���{f�κlλ�@6ø�����@v��#LE#q)$�I�A���N!Ѕ0څ#���i�چO�}~�yHf��T�&����$�n7 m�E8i�4_�T)9�Y4���ZC����+�Uo����SR6Kq"��)�H��c�j"���_���_v4Gx���ƹ��7��AƢa'$�&ۍ�u\�D�G�>"�b�mB���)��G�AnFmC��6����J%$�����!�~�Ο���|^�P�x��d`ӄS�o�
D4��O�Eb�5$���[]l6ɫZ{u 6��*��Fڲ��*���'UwSnH�mAK6����YO�#�i��-�x�|f՟1��s��2)���xj%,m$�M���u|^P�4���R�E>;�_�8)4��� �0څ#X��i0��Y�%m�$�H�r3�"�������?|���)�є=7�x��d`ӄS��Uy�n4���8)��q�)gj�����<v��ڇ�����H�N|�n~u��F�6p�L4���|���)7�W}��G����,��eG�Ze��1�12�q%��ش/�� C����lY]¨+)k��A"!�6�m���~�|D�f�0�~;����C4��'��S��#E�zeB���W�J��P����p�|m�X&
D4�w.5,ڇ�k�ye>4��y��O���Lo�Q9$%�̎�R<i�,�ёL4����|r�y
G�M�#��)����H���n���ԍ�$���j��)��G�AnFmC�㾿z<�3O�!�y�E8i��A��*'$���m��S<�#�6��p�|m�:f
D4�w.5,�C�6_���G�����ޫ�p���U��l�s���]�����P�*
�v82��ۊF�6ܑ�j"�����a�{WݍŞ8F�`�7���Ƕ۔�)�׊��*'$�&ۍ���|i0�0څ#�SM4���܌چO�}~�yHf��V_�j$�2F�RI$P6�"�4��'�T)9�Y4���Q|�
F~;���mC�,�B��	�N7%"c�)�x�<�ڇ���mY�O�g���aӤ}���S�!H����܎A#l��&�sK?����
G�>#M�/�Qs�M 1l�i��}��� d.GgwB�S	�v�� ��C�;��f�p�����]��lW0��I��<.��۷b��*��V��^��w�N�����۶�����߶x� �@     � 
� x     
��� 8B����� � 
�l  U�*��|�  �� ���<v��v8����N𭫰U_Z���ۨ�ª��*��ePU�m��.���l��M���C�;�8;B��#FW�T)9�Y4����j�)i��6��-�Ĥ���j~Gu������׌O�#O��g�e?��V�di�N���鑖\M�[m�$G2��)7�ig��E�C���O��a�;�i\�4�O�	JaH��q��7�C���貟���h��"�:p�^�P�x��d`Ӈ��Zd-���$���qL�4�w.5?#�������|i�k�'���Z��2���(.Zl$�GQ�QKh�wt���PT;��^�dmYAYKu��FD�D�m��jBd$i�O��ݗ�e#O�m��Q�����F�����a�;�if� �J%$�I����@b��C��z<��?|�������.�o�Ͽ�J��4�b8$b�}�ln_�X���|��\�Tc�}���~L�ّ�ҒI$��#�ݕ��nU������[捾��c�"��rHKm��=��1m�Ų=כ��}�[�]=���∤�)�a�U�ݲ�]˝�e5'n�@6ø�����U*wn'%�[*&2r]R��S1���ݨM�~�cGw}���r�����*'$�&ۍ��_{}o���^n��n���*�~�~��Mp#LPF�n�I�Dm���av���u�}�	$ |$�$ՙ��\&e�(�����*�1	1��(�7u��d�D�N7A0~�O�߼ԏ߸�{jI�YD��I�I߱�h�LI8��a;�{(ݒ{(���N������#�~�߯�����<[@[l��z�o[�2La8�bg�z7	���>�O$�!/2��.�=��n�%�<�y	��g.��BfT'XL������8�~���UI��f�`�ª�UATm�P["�[g�OotR��n$�L�#�?S�~g����tf}�n2�>a�'�ᖛ��a=�$��7�I�C�=�2���ޡ����S���?����IIq�$m�Z���N]g���5d�d�d%����$�k�Oz�8�;��拒l'��e�N��8�<�L�i��۽mֵ�ֵ�o{ӭj�E��h��7����<�	���n��L��:�>a=��Yy���'{~��:�-���{{ֵ�k[�����I�\�Oz�:���7��ߴN���CH�:�e����}ꃯ#�¯�6[��䑶�	ɛ�y#Mv� �%���Pio����Fn�B~���y6Zm�!����r4�l3)���y��T;���ŕ����9�Y�Q
2LQ�m�$�A3�"�gG?������ȧ�щ�]�G�/,׀R�^���B�j7$���r`�a�hbK��ewP��cW�>�����O`�_��VuzNT����I$�	<dq���-S�R4���� �1]��H�^8�/��x����$�Q��pH�q�^S6��)�s�ω��]2[#� w����m#MfIU��rHKm�����z��
FG�]�++����{� Y�1ѹ(|E?����H�⍠ۉH�,��r�A��Z{�u�����ø3�ꪓ�1��S�yu{w������-���Ǌ��g��@�P6-�� �m]�^�׮{�w�5�n�O\���;� 
�  T l   �  w   VW��
��
� cl@ � U ` �@� P�>�k�*��rܹ���kKW��֭u延�t������� ���Ϟ �fe�R���q׭TMvي����{��_��ތ��ŽZ���i��o�Nb�O�	���N|�J#�Gm���ﻴg��ַ��{�ntb�f�L��}�XJ����m��e����[�w)�U7�:uʴ�V[w�o��ވ+Q9$I6�nFd��޿`�[����{P����y�Mm{�&�$��7�I"�����껻�Z��Xv�����۝���� ���!N&�y��s(-wm�� 6øUW��*�� U^��-{�K�m��n����F����4ɢ����]zvGc��H�v`��Z������G ��K�4)&��ϼ$�F䡤q��%��=��vz2)��oG�T��5��\&�rHLm�$�GNb�O�	���H�!�պ���Fy��6�yLڇ��Na�I��q�$m�~&���eﱑO�{�W|�#�ݣ5���z��
FA�.^�\i�nI9���jGN�G���twz#��|E:f	i��ugT�8��5Ѧ�I}޼��;�����J��q� C����lT6¨*�f��.��㈳m��nG�T��<>���)�Wi�A0R<iD4��P���1������)	m@ܒFۅ��mC�S���韉�}�y��Dq�zZz���4ɢ����Z�x��D�[q(ڒ6��H�Hzu�ⲻ�x�籫��xI���CH㧼;�ͫ�N�(6�jI#������oG�T��=�o��)���}�LG�"���V�"��,�k�I#m��pH�Rv�6��)�}�����V�y��Dq�zZz���4ܞ�T��p媧V�,�U8��l������Ve�
���h�u���iI$���`�[��0R0��.���C�G=�_,��LtnJG1^(]_t�l��*�j�G��j�FE<@�-��j�B���ݾX9��>�&
G�!�}�&�Q��R(܄S��d�x��!d��N��0�>=�1�"���W9�G"ȏ�Z@Ӥ�uT�M&�B�V�F��/�X�)�[��0qx���
g��i;}qG�s�<K5�I$�������L%�B2VJ�3#��y����O(B<xl�U�#�g�M����ΉN��fζUMws��pw
�����6�Tw[eך�7�$�m��{2pS����*�	.G���f���%6��=_��Fb���m"��߯��__m�15��q�/�[��~9k ���9$I6�9�t;�+}���K6�๋�1�c���|<.$dqF�m�a7#;3_�l��w]���3�-�$?no�_&|#,�Sl��i2�|}׾]�^���C}������{ۖYwc�$n'!D�#Q�l������[D�G����}��U}{2 m��ٻ��ٌ��[]j��؞�K��<�z�UKd�ew6�{�,��ohm�ʜ�^���@*�      �   �  ;�� <GlGp
� m�� @� � *� 
� *�J� /��� � �ʡ�wR�m~�N���zz�e@=z�^�@�w|���|�n�ڲ���w6˽.뺅6
�u5yo������F�o�
�{}pY���\,�m�$�H�r=�/��}���")�+�����x�'1L�j��IW�\"��V�)��I*m��S6�N����q�/j��傟�]�16�r�>9yf���ط��3��Q�$�$���a�=ذS<��#�o��D#ps���:lHm���Wi'*��I��H���p�#��ܔ�7�1U�#�ew��a�##��)��_�;�0QM�ɎF�
�����ڲ�{� �w osT 娩P[xn!
D�Jm3�g�x�b�)�W��M���8�o-�\��`��a�~�P�5���t�l��$6�!�-����a�6�X)�V�#��5p�F��:7Ҵ�:]�QF鰩��R7$P3�f��^�Pi�<G�[����\F���G�Nyh�}�g���Ȩ���HKm��x8�+W�v�x��!WA2��V�ǲn;�Q���go�>#��/��E�#rI�&о��P�6:_�Xdqˮ��\"�#��ł�b�i�}qG�Ә�	.�uj���e���X�ެM�p����
�l 6����.��vh6�I��M�WҴ�:z`6�zT�`���#�}�^^��i���x畛���n%$�F�@�S8�#���u�\ꘅ�!yʘ���:}�}3�G�x�L���r3J6�n+8E��1�P�0�J�Bő���f�$���^:E��b�>m$JM��$ڸD#��:7㇬��#�Zlu�1���5�H��L�<i�d�	��nI"�G���[�}�f%���֎���Ŀz��/�cy��4�~*��F[���#hI��oU*��T��x�`�*�z-�������;���y4�HӤ�i&�PI7p�2VnU�"�����ao�^�b��˩;%������.&�-��!X4���i�cW�a��*�G��z�!�W��G�|8�Ţԑ��H"��/(G��}��"4���0b[��.�uˮ����x��}�^;e"T�M��I��7�,�>��FJ����Dx�G��uB!zh�c�غ�$�?&�J6���0q�9�.�oۼl��RدL�z`/���fÑ�Zi�a��I%��a@�W	P�� �ffP� �PU;���	� �1�$�Oͺ��x���������Ϲ�YI��]�͖bq��Z:˯�U�&(6�m$�H��.��Tį�Y:}�q�"���������0�����q3�%&�iH�m�hX�<r�	�,B�s]X�˯�W�Ep�F��b��x��*N�
���d��!2�̕��v�aF����Ȅx��ƬQ7��	��`�2�6��H�F�!+�}��S�����>:}�q�"�����r��x���$�$�s�kY�h��[7���VY?s <   <��U�l��v�� �� Um�����x���v�m�� �3qQ�����y�۶�6�{�^��{�����O[.؃����[��p�������'k�u < ��v��0^ݯZ�נ	�S8x8 s���< �6���x8i�x����67���kP�Ͼ���U��U*�w=�@�L`{����U�;� �.:PYA�   60�Ck�z��;�P���:��z��i���t�    6�	��*� �� *� U���'6λ *�+( �
�<���� �懸��w Y3k;u�Z9��n�ek�'#�nۿm�;�[��d3�����Þ"�UŰ��۹,g�w�S� �`'�      ��@  *�          @       ��       d  w                   | ��             m�          � T�(U ;�   w    �        U �
�       z�  �    `    *       ;�@      
�eP �>         U   �    *�    
�    �      
�  � �    T
�  *� �@   QY����     �uy@��0-�` V�	���_o�~�vkg0����R�1���i�W�Hw;aU������ooo�G�/WwmJ��LR;�UvѱSJ�a�s ;�����ޮ��l\�w�ׯl�߹�t �   �  � �P <�  �   �� ���S�@ � m�ت @ U   P� �E����~����*;�7�߷-_+�Tƶ@�w
����6�Tw[fS�����I4�I�´���3��z��#�.����&�Ol̺��.��%w���LN>4z�x��Ĥ�I!�G Y�x�>0Zm��V��4�F����Ȅx�wޏ#Nyu�L̨��$�n7 ��b�8]!�.�P�2J�B��2Y�N��a|{&�E���p�Q�l��m��E>#��ĵw�q>}�/�,��ˮ繣,ķ^s.��-�i	���K�9$I�)8�a�crP�8��[�Y����h�F��F�JyB�P��RM*P�g[���v��v��ר U⪯E��[j�
�����oj�p�P�I�b��]�9v!a�8�^�FIY�\"���A�u#��P��l��I"RI6�M��Q�����m�8�Gt���Єi����#�ʞ���0�.�_䍸�m�n,�.�!v�W�a�c�rP�8��FJ�X&cDx�0���-��t�M�$���;��F��o�����Vm9�Vb[��]h�z����|�x��vQ+8E#n4���$s)F���v;�Q��x)�h�"����%��"���,Y^V��kD��UI �j��n��� N���� a�/fR�w T�*��k��t��U�{�;΄/.�x�׈�'m�p�F��to��<p�[�#%C�~��I��I*D$��a
����"��7�Dx�W{�F�B0�'t�+�aA<Q.�P����g�x�e#���s9x��VUu�����Ĵ�L��^"��i/�D䐖؎H�#L��|��iAn,g����ܳ����3��4���6�
2�jF�Bc����ƈ�N�7���i웍X9��㑻�<Gt5�D�J��	t������n��e ��U^���6�Tz�U���L�6�,_���gU��qy�R0�?����j�藽��> [���I&�I��M�Ch_�aF2��Z�|�DkH���O������s�@÷���D�J7 rDr��4���~F�O̌��z<�x�F��}��>�ټ9�����I$�Hd����1oG�eu-/=W�/�ƻ���Y:|.L���V�nR!D�%I�ZIF�M�di�tv1>��i6�g�`^-��A�C�}��K��>!a�}F�����˽{Kz-�9�� *�qUW��6ՔE���]n���UqI��$ھ Y������xᐗ�ک�ّ����oG��Hҳ9�&4YqI!1��(�x�yY��x9-�fZ<�+�ļ�^h�B��k/��4�nx�X�m�ے6�nL�M���e�<p��	h=��<F��X+�� �!�k�����Km�$�4�x���Nۊ��g�L*��#��F���W%�Di�.j�6�M��e�Z�E#Ow�X��f��`�[��.�y�WS�y��/�Fx\֫�9��Wt
� ��=��p�<
��c��¨8mة��S�_Wvz��yMV� ;���e���PQ@{\ m��uq�H���x��׋���*�P    
��   �P p    ATm����6�T@� U ` �   T ���>��w ����[�ٛy��x<��kdEV�-��@�w Wu+2����PU�1�	��Lj�6�I��#��s���?j��w���> n��'�x�#����NE�/����m��j0b�H��`��}���|��!�w��#�i���r~��K�t!�mI$��24�������R4��}�i�Wi�I���H���r�<E��NB6�i$�D���5�ҥ�����-��og=�����7}�YGɡC�4����a�=O��{^���_������K+�=��kM�)&�hR)$�	�x��W;^VP��U@
�l ȫtNHc�F�G���R@c��,�����u�z�u��x�nvu��I2�n)n2盾ι�vT~��ٿnwd��.���r�x�����$�nH鄐���rS�=O�]{^���_�����G�%�#q)$�Ha8^����Q�xY9�Ǎ��n��}�d�90]d(��$�q�!�N��8J�w3�����S��}}-�Rmq�J���^���Mݽ��s�x��P�*��[+e����m��z��o*��U�!��w�և�m�}��|��=F�l��-�^[�t�Gl�"�H�J$R��K��靝�S1�K���P�mIrzŎ��L6�M$�IRM��nߡ�nL�\�v^���Py��}�\h���e$�IS�4�R���M�]����r�m�1r�Q�[-z�`jHۍF�a�-����˲�/�^���T5�`n���>��R)VX��
�v��2U]ղT;�+��J�� AU��#�]t�@r�_�/�:�޻N}%˖�C]ܞ�P���TJO$���jH�jY��m�����W.Z1����T����f������m��*����I�c���I�#ps]�q�$5t�g.4x�^)8ۍ��!&0S�O�N2cW%a�x�ɹW�v�C�n�a� �qr���"x����T�m��t.0�2�\W��O��5p�zW����X)��Z'��W�#�_V��,N������u�*�W�3;��U�*�ʠ@ʹ��u��A��fF$c)����A�!���[傗��H�n+�Ft���|p�8\��m>fD�MHܒ0dy�Cܴ�s�a�8dƮJ��웍\(�;�:�3�����7���B[m&�C/+�~�.0�2�\W��O��5p�zW���X㇎��Z�.�I��M�Ch\������/��6������lweX���l�
0�2<AX
��"I��r$G8��|{�,.̕�wLx��Hpɍ\����&�\8Gڿ\�ѠSn�mKm�O�U��[ݺ�R��գ��ǎ��m�<�#q[�w{��'U{u��h��z���UB���� ;��m��������oU[&��]��`      ;�   �  �  xOTGp
� m��   �   P T P -��x Ų��UV�l��/��,��n��=۽�w�@P�U�-���VS����]�M�퐢RI$��$��#����y)�ʟ�\��F�g���dq���\!+�7�pQ9$I$�ys
|i��D�j�x��Ϙ�|E9�t�i���`�yS���q����-��m6�a{�sJ�p�8z	V\!�*�ǌ<t����Xa1dH�Kh �m�ZI4���\8Gڜ&y�p�0�(!�ʒ�����.0�0_Z�҆���$�KI4�m%I6������.m�هH� ��6�#OM�."��E�a�΄�Z�4PH�^8ln�67U����� U�
�R�wT�
�0��9j�U�:�ʒ��Se8Q�Y�5Ѿ�4�t�2��C2V��s#�0��j�6�ML��j䧔!<6{*��!ݩ�<ѱ�2�\��4����pلi��l��T�M��J�*w҆�\�j��[�'�m�t����ShB4��~B��!��t�TI+i��I&�Ubf>�&U�^WJ!M��Fg��F�P�!�0J���[)�`���TZ��m�R�D8a�1���P�x��쫇�v�L�
�#8d�qr���g��� ����Uu\�U��V�/T� 6øUW�l�� Psm;y�{/ UI"[n��f�κ�%"ɸ���������t����Єi��MI��8b����8���X�ķ{fg*�w�̣���+x�ķ�%�u}(i���i�i�m�RJ� 雄3ҷՐ�6Ga�1���U���$�1:��{�x�:��g��٫G��^e���ƓR(ډ}�%#:^P�l�4��}(a���Ʈ�����.m�هH��iN�m�RI6�0�ҷhB4�J�!p���u�,B,��I�b�%��p��о�I$Rl"�)��m$SUJ���oF��m��]�l���eKm�<^��6)�;�9�����]���0J���[+!�l�0ä>2cWҞP�x��쫇�6�^�D�:m�UUT�m�±�L!2�JFzU�F����"��������AĕT���)4�����:D���ShB4�O,B��!ͮq1�/��V!˩(x���"�m6�uT�R��E������"3�.̕�����:C�&5})�G�`�SE�m$�M����\8D9�:g�V!a�;(!�]ICH�J�B�����}(a�"!��J$	i�U��e�,��:�T;�7�U*�p U++�m�ک�nU�}��]%o�p�����0�����ЄiΞX�ÄC�]��+�0�ZI��j�I!A'V!˩(x�6S�E��\�W҆���U�fJ�Y�dq�!�\!�QN�I��m�Zm_JyB��'��"ڝ+=J�#8ge8˩(i�*�\8a}���ĒM$�6ꚾ�0�|x\ܫ�a���8\�DCfD���ShB4�J�!p��U���a)�i6�I*������L��Ԕ<B�)"���W҆��4,3��ܾ��}�Ѡ���ҍF�IEc������c�cl��L;����1�q{{���wlm�p��wQe�du&�l� ;��j��.��t�ճk~�� �@     *��   x  �  T�6��m�T�   �� `PU T   C� <׭U�@��V�u��uGpN�U���;��%@�w
��PF�*��������򩲨�R�D8a�1��O(B<{'���mN���Fp��q�RP�<��!�cID��I$R1�|x������=sq��#%o�p�����0�����Єi嚁F�$�l��%�m��r�;6!a��ɕb2P����gx��_JD8n��I�%:�M��M��n�ڱ.2Ga�1�⮇��{�Q�/XV8�|u�t1�ӊI$JF�m!���rE���.<F��>�,�a�sr����6����l���ZH�T��2L��6Z�V���;�� U�Uk��UaT-��m�R�m�(s��e#�E�."=g�+�<t��V!�%�J|Q�,��s�&۪��i&Sl_JD8lt\/�I�V%�H�:C�&5})�G�M�7p�!ͯ`�PU4�I�6�T�RAX�Y�젇u҆�����Æ����P�!��n5p�d��G{ҧI�M��Ȉㇻ�ZE���C�����c)���SF�"|w�X8�rG�$�E%�H���<F��W҆���F˄Y��Vq�8���ɍ_JyB��%Z
��H���Խ[Ҋ�n۳� *�pz�J�� E��[n��އ8�ܩ4�I�p�!ͩ��S�0�ل!������x�Æ����P�!��	$��M$�S��WFJ�P�s�a��uM�ӝ*��ÄC�W�ˎ#������iFQm(�"D��7u%��p��<�*�P�!�}(�p�2V���2Ga�<M%�r8�i%-���C��}���#�mN���Fp�aq�RP�3ү�p�4����H����m��)��C�Ǯn5p�d��1�ن8<A�T��=</�\8D;�}}Tؤ��vT�5�{�j��3{d[h� �eT� �ʥ��fT��7L$ՈE�t��2�C�RP�
l�
0�3��b��"6:.�J�O:-��UE�m���ҲD8a�1��O(B<{g����I3�;�0�(!�]ICHY�n�Dm��I$Kt�F���C�̘���^�1�ن8<A�T��6�^�A�TJ-��A0��_ȬB,ç�I�b����Se8Q�Y����P�!��!�*�:M�JIA�7fJ�Vq�8���ɍ\��#Ƕ{�Q���aX�a���:�K��=Eh��h�U/^�OZ� U����*��l*���wZ����[o&ʛ��MP������*��#O��R0�i���Y�3ܴ�'dDS��EW�Y��uT�M�L$��ZD#M�_#��\�bf=bL����
��K4�:��1D�n#nC�Dr��)���p�F���	x���Lj�S3�sm��̑� W%I�m�����m�$�r])ݗ�S�3jC�}ޓm�Rez�i*����)4��+�]}�hwI3���u�[���\ރ�<��;վI"%ۉGm�(x���{��N ؠ*�pn/ '����[�I��W�s�U�P6���׺彐Q*+�� ecݹ�oWm�;�o�O�y��~ m��     �  S�  <   *�P �Y@p�   �   �  @     n#�T���}�.܀�w�W��פ^���oqg@:�6��ﾠ�w�ԪU� �-���^�w�'�.m�l�������z	�޾��a�o�oi�~^=-���*[h�m��I����]]�ޗ�I��S�/z�!.d��}�Rje�Sf��I$�E6ԩ2pR�u�t
��I1���u��=u$���6�Q��8��~W�Uf���4��
0�FW�)̐�4��{�HlQ�I$�m��-6�JdB<{&�W��v��y��0قe!��qE�T��ǈ�Σ�I"Bm$��&8d�?v�۽�n�q�j�Tl;��e p m�$%%!�($%F�q���%2��S����\!+Hॺ#��<G@�!o�_��p�oj�pF�4�m���L؄Y�K�*�/*J!M��Fg��F�P�!��A��d���H#*WښN���!%h�pä>2cW%<���ƮD;�:g�V!a�'�b�˹��i�J%$�I"��#L�Q���C\�j��[��DCfD��!k3�*��IF�) ��p����eCbf>�&U�^T�<F9�F�s]�CH�L���TRO�n�I��2S]�TJ�7 P�UwEQl���E���)6�m&�1$ԍ�ps��ܾ��3#�0�����O(B<{g����N���Fp��PT�6�%$���!yRP�3�^!p�i��>�0�a뛍\!+}C���l��-�J�M&�i6�6�����=4_t^<Lo�{�������39Vc�Ve!M��FfG���i�m��I&�a6��JD:zh6\"̕��Lƈ�:C�&5rS����j�DC�K�"\P��I$�3$���<x��ߘ�J������Æ���P�!��n7p�d��`�PD�RE"u6���)o��}_P�Yz��� C�{eR����UWs�Z�z]���_�����o������}�~��O�g��E�������Xىn?=�3�f;�fQ��ʹ7�f�H�-��I�����;�^C����%l�1��<p��Lj䧔!�e�A����9!1��E9Rȧ�I�aX��l�(!�wP�3үÆ��K�x��nx6�+�m�ܑ�r<��_jN�G�4�.��M��C���p�oj�2�����U*�UE�E��m��L�!��8��CӯZu}(Y����,�[+���#�n>���e��(Hd�2JA#�Z�Wz�m�
���
� �V[hݶ1� \�7IB�r<�������ȯ�#��t���~��r�*Wu#=*�\8ae�\"�	�a&�m�)�}(a�O�dj��[��G�x����ShC�L�\8Gڝx��;M$�IStҦlC�:|ęV8���!M�0�zp�l�J~���ap�2V�y�'Β��6�m���~���dƮJyB�&�W��v�L�
�?CfK����j���K��I#m��2)q�i�>�0��ϲ5p�d��c��4�.��M��C���?/��-�$�G{�˝�{w{@Z� x cwl�m�ٽ'U8   ���U�q9���] ���m��1�p77��q�m�7���� �d�@��1�p��ܫm '{8@y� 0֘�1��g����W��6sh�  �p1U��8 N ��a{��������-�\ݶ���*�zn��� �-ݕP*��^ܭ�
������f��@�*��  ]u��T��J���^ٴ��-v��-"欺m���P   Uթ�� *�*��    -�+*��m��UQYU@ U� @ �Vo�n��T��r�wgZ�ݿwm��mݭ���p��m��sml�%兹���e���T��@�Ƿ[�G��{�h:rw�8V�      aR�  J�            �    l U    T� 
��T                    
��             T    T  �  �  @m�@���   @    �   pU     U�T *�    �  m�   @   @      w @   @ �           T        P          �     T*�  n  VUP    +( 
�    ��   UlU��^̀   �9����`��]� ����g[s7w��3l/f��`�÷j��Px���n�Ų*f@xlF⵻mm^��M�i���^� ���W��m���mU ;��ݎ��X�ݴ�wu��Z��w���        w T <*� w  �l�PU�T� �6� � 6�� @ P B�@U�x 
�����=W3d�ᕠٴUU:���n�P�UwEQTm�PT�׭���]k.�:�[M��a�.#��_�T6!�>bL�^Wu��C=��7Ҵ����!�*�:M�JI�,�"̕��p?��N2cW%<�~�m_Gڽ��q���c�Y)�MH�mƅ�.뺴��W�����}+�|�#y�3ܾ�(��?CM"����5�ET�M�L$���ڇ��p�ok�1Cp��1&U�/+��F94a`C؍F���i2�I��I�7Ҵ�t���C2V��wa�H|dƮJyP�=�s&�(�HѤ(V&�T�����u;Վ�@*Wt�W�T��T[.��ѯt�06�e�������s�1r���r���#��|���*����)4��+���Z�{�|'�\��w6_}���~��0�Ƌb'$��15U���Dv������s6�=6�{�=km�ݑ���7 rEr��n}�7H�n�����:�o�lt�n6�-��(�z�۳���6a�H ��m}���O+��,�ˎ~��w�\Z%��%�"k�ݶ�{Y빰5{��ڠa�^� � �
�Z��'m3c*��o�ʒ����x�>��to�}���Y���3�:C�HlQ�I$�m��-6���P}۱���N<��0ӆ����U1��Ƒ�"ƛq���(&^@q�g{��!���P��?��#мA�T��T��_������m��B�V<p�eX��I@Z��(�}���JD:f	V\.M���v�B�I4�I|��5q�ڑ\���[r�d�7�92d�uI$����M�m��%6��M"lT�z� 
��*�� �6¨*UWu���'q%�I$�F;;϶.�2{�m�*L���u.OB�u�6�3�S��I��I�m�������B,ç�$ʱʒ��Se8Q�Y�5��(i���E(ꚪT�M�àY�E�+}X%�Dq�!��)�G�l�5p�!ͩ�g�V!a�� �CA6��HKH�F>�����c8��4��䡄C�ד\!+ޡ��:"0�=���T[M��m&�й+v�#OO��_ȬB,�+��X8�rC�@�"Ñ���������-���w�c��@*�qT�R�T;��J���礜�sA�m��bH&^C�8�yg���^=�|C�o�ͪy
F���L����\�s��$n%$�G!FH&
G��iiuZ�#�Vy�i=����<G.v5��m[�������i��M�Uh+�DB!�=�����4��~W�_ȬB,�+Ot��Ԕ<B�g�H�%�e6p#H���:	���!0\"�uoVu�Dqp��ݍ^�<�#O?��{(5$�Ĕ��$�(�9�����H�n����R=��,Y�0�>��P�!�)�D ��n�-�yEG��MU��N���yV�S���wb�m���6��p�5ݷB��Բ�[ku�
�۳���qb��2������.� �   �
���   �  �   @U ����`� w � m� 
� *�T U����%]Z����m��w]Q����m�nn�nZ�h ��
�P w � ��H0䍸ے6�r/x�m[�p���11��;��k>�����}��x�ok��Ebda��(�$JI*�F��]IC�c��G���_F*�P�!Ħ\!��ެ�ƈ�8���a%�n4����Y�}�)o}����^9����4�4څ#>�<�?��j�4a&�H���0�F�\�8�|wh@�:"#лA�̡�0�h��">��[�V&�i$��a&�B,�:���1�GR���z��W�/�G�����t�V���i|�F�F$�b�m�75,z�PTت�� U��E�nG�?�1���G��#��t�Ư�]��=��!�:���Y�!.�P�?h'�I$���l��`�H�e�<Gs;"�C6��9���C����6��3��.�S�"�m������gdv!F��U�^T�<F8���������B%;J@t�l��*��nώ|�r�E"�����i�w�qDC�t7�;#��Έ�T�j�StҒ"0qg���{<�t���P�8�]������c�!�#��]l��Ƚk��ܺ��m��׫� C��W�T��@*��m���j���D�JDL�f�yo��M}�9�_j�K���nN�6ѥP�uM��m$�!6��lޚ1���t���m�������^x�u��H�IF�H'__ZEVۃ�B˿n!6��S�ٝ���G��N�qR��4�%&�VM]�q�;���f]K~��^<LMx��Vy-��{9VbfQ�f��(�6S9$H��0f�:G�����|G=4.d_��F��:C�&5b�#��y�ɔ�~e��i�$�~H���l��WU a�^� �
��l�z���*T*�_:�;�������H������j�\�NG���&�0�~5Ԋ_|m��-���#�!;�<$�DCfG�x��C�÷��Y��q�-��#?D]�%�ꛦ�J�IՈY���n��x9���"3�.�꾸�a�H��#,��nI$�c���R>;�1����ް�qx��"�{�R3�s�e>4���.���i�IBԡ}(Y��Ɏ��G��	1�ن�g��{�R<v�9�8��8m�A&�����EvoR�J��׮ 
��*��F�UU��j�ߵ�l��&�&�iX�,���*�,�CH���<�W҆������:��d�ꉤ�I��D8a�1��]#O��5p�!�:��#=HB�mB���ƒiI$�C$C)�|e��چO�}�貐�?|��1�ن8<A�̡�a��Lii��j��0[���˒e#c���L�&U�Y���n��x9���#��3��|"����I�(s���m_\h�0ä>L��.�����Q��*���g� ��m�B�N'��R����ݍ�� ؠ*�pg��m��n)ƻ�Sw�w�N�@պ߮��ܷ��*TVٳ��6�U����o;����ݚ�W��*�    6  @x  p   ��@le ��
�� m�*T m� 
�   �<V�nwhf�Tcwn]o^S�sM��.{� M�n��^׬����l�U*�
�U��t�;��L��-��=�x����e>4����P�8��gc���C�LtD6a�{����$��7$��"1���R<v���x�1�y���g��?9fg*�v�Q�2pzx�<y��]ED�$�q������C�ӄ3�:��4Ga�&U×C����\(�t�|�L�LȓJI$���`�x��h!
Y�
F|ny�Ƒ��jE?����C4��l���D�J6���:D���2������˒e#c���L�&U�Y���reI%���z�7vի��wke�����Uj�+�J�;�*�@�mw^�6�櫺�@�|l�g5����C��2Ӆ�u�M\d��>��"^a
�l��q�S����z��ւ*�����/�؅چO�o��$~��rF���_��c�!�#мA�̣�Ǿ�����cn�׆�<�����c���t�%$�m�:�2P�-��a�0�.k��CH�M�t�x�U���a�H~�,�&�I�i�Rm\*����\(�t�k|F8{�)f�Hύ�!���>7����q9 u�T���a{d1��� ClUU� *���
���u�Zw�/��t�_J�!�ٓ_���2ab0�=����0���!p�ٝ�D�KI4�T�$�F��<t�eX��+H��ð����i��4]8F}Sͽ��pƤ�7�F�q����1��]q}�1�� t�%�u|G�>6���U!��A8��"J6�0��|in!6�"�����e!�;�<$��6a�N~3+��m�ZfB�P�䑇�g���8��,I�bd�"��#�W��J�!�,J:*�H�'B��l��m�4���q���u@�w��UWR �����#I%�9$��f@�Y�a��,%1�t��Lj�W\F�gLj�DC�Q;�
G�>3���i7#I�nH��9�|��/�^<|�;�����Zy����W�#�v����l���T�aF�$�m�Sc)���x���q�![�X���:eX�ICHn�����%��i% ���2F�,����4�p�.�"ȿS��8���ɍX�C�a���Q����I��m��%�#�O��-��}s�Y�wbm����b�s�f�|�l2SnCu^�n�J�v�ko[�w�@�w W��@w [�Gv��ݻ���k��_��v�\��Z�ݞ��������>����g2�NIM�	.]�?tٷj.�c�E�j�%�)�m�GCm��uI��i*I�*d�*c����H��p}s�Y|��>ۗ�͐W�I$�I$�N�u�ٝ�&.OB�K��t�%�%�Gd��
#���I&��T�N��%�=:���L�f�]�W���Ύ�A�IQ�ЈGH�:�S���`������{d�6�nr׭�ڷ/!������Kd=��P���U��J�
�X��ʽ�������o]�֦U����i��   �  Wp   ^�  ;�@  �ATwT �� ��  Ul  U  �T� m�� 
����TwM�l̰�f�m��M�]l��lb���Tm�PU^���Cu�U 8c������+��_��5o��*_Z����I(Z�W���슫�i��.[hx����hϘ�c����j6����2B7�~�ث�gp޹�zvuͼ"�x�y��Q��M�ݝ�-��͝-���"q*a��,���HCH�4�:H��K�I$�d�_>#K�|C#�߻*��#�::"�4�6�� �|D?n�hM��`�+j���JU7�ش��@P�*�©T6�T[;����������|p�!H�c�C�X�c��0� Za�g�sn�qf\��	FI�'"�I"
<�B<^ތ�<i���Lj�#�a���QG�S�g���{��A���i&H�K4�"i��e>4�����F��o�R<i��=�ᦑ�9�I(m�$nC�����o}�����<ۼ�ݝL|��2�qg���x��a��\��I��M��9"�#�S�xv9�CM2Έ�x�1����4��cW
#���������ݻ��T��]7���Tl;�U{)YC��@Uݶ�ז�(d�Ĥ�I?(��H��i!
Y�4��P�|in!)�>?f�,�x��
�2NIi8���DE8x������w�/P�8G2�Y�������Y�o���x%ц�U�i):�X�6x�3����G>�.�"�/�h�x�1����4��h4�T�d��m��j�Dq��/��H�O��B��i�r����>2�BR!|~��T�k�7�F�)Ô�|t�숊p�H�g��p�#ڳ�3��̙t���!�t�IR�2�)N��������j]@��U@e�ATw[S׵;��ƫ��WE'V8��a@�a�0�j���񳾣�a��t�D�Ӻԑ�IB�n,�������,�?�^�H�O�E��,�����P�|ir�&B���ܒF�a5��p�׼���H�{�DiçH��M?��n՞c4��8m��H�6�m��pG���Nǻ��a�t��_���F� y[)Hä��Y��Y�F�aG��>:~!��\?q|�cW���L��~�1L?����\���1�$�D�EĥIl�)O/T UUz-���l��l��)"LQ�6�m�h{��#�=���>m��U�8�:��{�m������������4�29$a�#���n��c׎a�ʳ��Vx�?'xK�X> �p����M6�)"Yr�ψQG�#^>�O��g���Q:fӝ�3���"�����QH�r�,�w�F������9��׏���_S�H�{����#^s��H(ܒ$�I*A$/����A1_�֤g'�A%�/T�����B�!�#0��d��F߂��W��ueU1��^p���n ���F��7��K��7
����v�p=P� �Z�U�k�λ��S�w�n6�nV޻���  T� w    �  �  A�U �� *�`U  ;�� m� 
� *�T U��m8U�@x�[z��"�lݫ`�[\�V�[ �wJ�R��QR��7Oշ�Dl��]�ml�Uo�~t����緣���.��rH�m��a9��|�����{�u�w��=�:]nt�KTK�$�)4�����5��xv!�&�p���(T96�I$H��(}/싾�h�֫g��yt�w��#1Iq�$m��~���^��:~:�5?#�H�}%�������zQi�u�S�7U�yUH��`l;�U]�PUj�
���ڎֽ�.�Wt�M��V���%��Ο�i��Hg�����i�ٝ�\e��M��m��s?#��C���g�#�mX��vB<i��{�r��\i8�m�]Sn���0���0֎��g�O�EO�?io��p����a%�I&���I4/�F�2tʰ<F����Q��Zz~��p�B�@G{�&�-��nF܁�G��2��g�C����ۑ\�.��>���M�C�$�3�ݥƕM{���W� *�qUW�� �VPVR�I��&�b8ۍ�ۉH���-5��|G��}i�n��)�������������%$�H!�!�|@[א��p��*��L�v�ӇO�
�����S�cd�ܒ4�b8$c4��f���c׎��r�>KOf��9�g7Y�x�>7.�o�E$ԍ�$&(�3�h�0���Ɵ�#�i��� a_�pR0�����1�TNI	m��{�\���ξ������h�&ӯ�_�� Ӈ�z�����O�E"�m��A"�m�ʪ�n�J�ޭm l;�+�J�;��,�S�p%�j�l�(,����"�t�_��4�|p�{����0��ǈݕ�?�D�I6�E6��G��]0<|g8�a��q�?G��/�5}����S.�i4��D�����Q�Α�v���S�N�_�di��&X6|�A���UUSIYMݢ4�a���#H��p��p�:fVϓ���]�~KOc�zр$�%'UTѿ���\#Ӈ�`�׹��ӎ!]s5���O���F�[a�D�/yƺ�yV��n�[| m�p����
�mYAR�����g��-��hRIr?~�����#Ƒ{�s�?'ɘ������}M��Ϭ�T��I��i!I;�Γ:e�4�xK[���-�|_�.�q�gɏQ����e��%��m�����F�C���������)M��Y-&�I���QMu��/���!�g?t�*���P���J��a&�i"�hl{��<�2��<C:e�6�%���E���ֶ�(mݻ��t�㄰�  ����S�u� i� @m�ݰ��f�Z�< =T����������3��������X��
q���T[��c �����sp8@xN��N� � "wD���r���[+(U  ' c ��uO8 � 
����{�c��8�7����J��l����'u`.�y� ���Sdj��]�� �� �  �w]�E�B���pUU��V�d��.�����x�mU@     6�e���  ����@*�
�kb��Px]�
�*T  PN��UPk�e�����y����W����Q�q���� �y������ݹ6����m�λ�����v;��x6�w���'p'�`��     ��   T             *�      U@       �                P                 �  P         x  � � Gp   d    6�   �
�    
�        �X  @   q    �       �P      ���       �                        ��    *� n   U *�
�   �@      -�    �^��n�    T5Z�*T7�*��  c �*��"��n������y��j��wvZ^����w]#x��{aNݝ���Վ��^q܂��?Vܓ�]�;�s*+lٶ
��)�uM��׸y����u/U�  �     l   � 8T  x` �Y@l�P � 
��  *�  *� e]� ��U+��k��ͻm_�דl��[u�*z�5��TP�6�E���TYuY�!$�:I&�J���8<F#����:F���z���x���S��S���-Sm��)[#N�(dO�"��ܽ��#�v��"F�Q���������K��IQ�ɆH�R)��e辦���י��<���s����ZgGy�8F����M�RL�䑇�,�i�x�gS&l̺����|���h]n���4���T:M�JIw�t�q�0�0���q}}ޏ?�߸�8)�:k�M��4�u�UV��n�m���������dM��umE����V�\��q<g�(�'�^̽��|�˓/��p��3-��$�R����MȒm��a����;xg�`����q�H�H�;�/��i��O��i��#I��I��çt�p�Ǐ(�aB�>0�#O��5b��w�R1�M&�I6�m��8)iyF'�~#�(뜆R)��v1�D#���4�Ӈ������q)#haY������.��p�%�t�j�f��[:��3fe��?%�����6�v��y�%;�f��ʪN��y`�ª�UATm��*��\���)���$JH�r�O��E�G�Ӈ�����Q"0�4�Ǣ|aF�v��m��I6�T�j�����U�N>Ofѹ�����e��y���ћ�at��~?�2F�%�ܒD�S�u�dݴG�dw���fP�0���!��wGspii!İqF�m�,�~gueH���ȳ��i��哏�eVsd|x�!��0��.&�m��e���YC����X����
�H�^����CH�ݞC)���ͫ����&�wr���zEm�k��z�J���U^�b��VPUܬ��;�UFJ�����O{�4��1|M�}��x������Q���a}�e�N}��S\�R7$��#�<�GA݋?3������i�~�Yu����N?��-�'�D�M$�N��#�����O������e�3ٔ��������{�iBE��Ȓ�I$�	$C)�W���0�:{�ɧ����6��24��"щ�eCH�Yt�&�$�4�b8$e��?w2�l�c�͙�V�OkƾO�����>#O��{��0D��H�WKu��ζ++{k[H�m�;�+ٙ@w T�*��u�ֵ�v��	�s��~�_���u5���̪:�~�g7�)ïr84� ��Lk�Q9$%��Ou��&����+ٗ��h���9�@������0���i�q7M&�!U��x�;�.!b��(&<G#��� �C�WC����k��TNIM�$�(�]C�4��{'3Wr�4�<B�1*��ó�5b���F�P9#q)$�@����<t����:�f�_S��f^���ӯ\�/}C{��������ކ���/o6�' �85]�C���M�m��ʽ��e{��\û�]�VP��x�oa^��b�*������{����\����wP       �   �  ;�   �UQ�P cl@ ���| U 6� P 
�@ C�U
��� /T��a�-S�w6]�U6�]��� m�p����
�l AW���t�4j�OG�I�i�]h�Q�[ϼ7�٧�ن�t�4���~gu_ q�xI%�E!��hVr��>#O��8����s�4�G��Ҟ���T��͑NHLII$Q���or=}t^h=����V��1�ݛ��9$�Hۍ�#l%-��$ݵ���W{����~GvH�G� ��	TM�[m��ş��P�P�?�ʳ��i��哏�eRoN#L#�m¯G I�!���QS<�^���q� C����lY[j�
ɼ�IFI	�O��iȒ���q���|w׽a���
G�#E���G��H��V��$�N�I!��_ݢӯ\�^�ηt|{�}zN�KOx�Zz�x�;����Y��DHIM$�I�n3�����wb����,��x-�g�����{'�����L�6�H6���da�D�ԡ�i�tư#�����a�m����CHN����$�(�d��)�W�ϵ#N��d��L�>��24��"���7�<~��; �9p�P�$P�fׯ)��T�m�p�����Am��ޒJ,H�,�䑆 ���)���3�����wb�L6��(zF����U�P��~*e�o�Q9$%��E�C<sjߣ�B���EO��8�>Θ�E>?��`�x�6��m3jE�#8�jF�YH�|]���?~�n{&��Ny���2)�G	���BdrHKm��He>�);G׃���
FC�݋0ڇ�;��"����#�8d��$�mC�S��3���U�zqa!�ԧ�����������b ��������j��V19=X m�p����
�l AWu�{7�oeکPM�pR<i�����=�q/ye8x�/��.JD>=�r��<wk�+�UD�a��RF��3|x������,�)�l�q�n���x�m0Rͨx�<q��	����q���6x�>�rP�!���C�3Ƕ��8D,ä?j��q}�		ci$���$��G�Y~:{��H��o,b�̣�g9E����fsE�Qi�\|W��l���H��H�P��m�!� ��W(B4ߥ_��p�ok��bf4�$ت_�M
eo���ڨ�u@�{�W�^�[7Kl*���m��w����m�
��M�{���~��_�u��oƳ�M�Q�c�e]�%OV_c�B�:E?r��E� �m��E�W%mЄx��cW
"��se�0��*�bu%F�2�0�3����R�I�i��A\�0�|{2��0�^�{mp�P^�B��_�ÄC{W��a)�a&۪��0�B,ç�$ʱʒ����#�2Q�(i�
�C�3%OW�?�Q�M��o0�f��{���8��6ھ(�;��(؇�l΂����Z�!��C-�䑘�*$aD$"aT���=Ȩ�8Iø;�Ӏ�PN �p�v�����Sն��i�pUq�Y�Z�^��Ԩ �k��<["�s��VΣ���M��D֯��T    P �   �  �  
�wlGp
� *�`U  ;�����  *� �@� *��@p�@N6���y�={���U����;�M��꫻�w( m�p{32�pM�m��S���f�������~�^eg�n�/�ew�x�w�g�p�G ���8�9�KK�9$�4�$Kt����� V!�>bL�^WuSWa�"7%?aO�I|�b���M��LȸC2V���?#��e�}�.�=�m��́L�d��W��*'$���Iġ�m��{<�w��h/t��%ɛ89�}~�dB�$]6���۠�t����K�r�2w��v*�ۯ���ח�$�I$���nsqz��wv׫ ��U�
�l�UU]��Z��]��P=�I���(G$�~�d�1��vMmuvg��TmU0�i:��m�M1RdΒ�9$���s�h.��3�&�I��u��D�m��&c�w��!��6�)�	q�_�:����.��'��(��I�i�z*\��6Ď�RM��9��5]���P�?o�d �6�uT�E6ԩ��L��ɝ%4"rI����)
�I<C�6�6��){:�?NgUT��q�z�P�*��[7KmYAY6w[eһ����B��Ϥ͜�ڙ2p��ro���%ǒgcr\��p4QN�D��m�A�Q\����,�r�2m�����o�$s|+�j�6�ML�S2^I���jT�л2�199�/F�wu�F'g9E�l#K�p�Ҫt�I��m��
�(i��̹p�2W�C���DC�"A���P�i��~B��!���D��;I$�ISM�m;�0���2�B��*i\a�YЦJ7%",t�!�+ep���h��i���%�$Ɠ0������Tl;�+ԩ��*
�wu��p��T�m�)��!f!�u!{g����x>�*�#8gAh1�y!_�'!�F�m�D�!�l�4�e�O�B�˗�%o�ps�h�pÄNA{�eF��0�E�UT�i��.�B��!��6kv!a��eX��IC�)�q�gE�	��4�:T�:$�D䐖�$9�"徬����t���/��Єx��cW
"�����0���j$�$*�St�H�б������2��f��-
}�!��e�p�d�z�=���>"�+�"��E5�(���z���otUV�;�UUPU�Tz���d�HKm��H{���C���|/�\8D7�&�n�"�:}bL���(x�4�0�,���4�m&[i&�ʓ�}(i龕t"̕���"a�,���B��=�\(�wk��#j7$�&ۍ���`�<x���A�wY�bp�_(�m���9z+}�����p�d��G<(�I���)4��wt�ۍ�q���9F'�s�����c{Rl��B,ç�$ʱ��C�E���p��m�ꉦ��7�E���f䡤C�����d����p�Y�H~Y���#O����N8JQ&K�E��u!6�c�<�ly�ֺ����
�cN���o׳h-ݵ@�Էw.՝��P kb�lU���-N�תʷz����o;�       �   ¨ p   +�6������
� p �>�  *�    ����J�x+��k�;�Pn���η��;���l�Jn�ewUz.ke����-�S]���Z��?:O��W����6bqǏ�*�l�w^�18{/�^6�|�����Lz�j<�m$�I$�n�'p�d��{m8�;�(�}Y�1>{�����6kv!a�.�B�$�I6�B�N��|��:�ϝy�ߋ�b�e&=w�Z̕���"a�+��Z
(�I�m$�-��)�G�l�5p�!߫�o�6b[�ϳ*�l�wY�bp�ʸl�4�i)��I5UT�)�W҆��^Z�FJ�P�����9A{�eF�M�."���5��:��^�r���۹Z�`P�\5@6ø�J�P� �PU;����,�cdٱ��$��Cn�P�4�0�,�2w��O��D�Cj���I#�ɶ�I�m�L4�D�q�j�R>>��j��8�׃��Fl��h1��R7��!cID��I�!�p��)��G>�j\!+H��8��Hr��T"�����cm��H&�.#��vvGbf,IqX��|B�/M4�?}Q�G��ǳ���o�Q�ԍ��(Fq�/�K����:C�=e�V�i�v�W��v��0q<p�m�W[rj(ڒOڥ+��ob��a�*��F� *�g��C�z���m2���s����Y�g(�m���9z+}LO?=�^���ZG7-�!��*�:E$�7M&�eP���B0��z�Äq�����B,ç�$ʸ��a�s+=����JIM�$�(�;}}�Ev�?��_��a�-�}~�����]/Ú��4��H��8�8orX`�1R)6̡pلip�B�uD>=�j\!+}R�i�4�6�U$�J�Mݢ!��r��U��>�/�\8D7������X�*�/*J"�zbT��Pk��k�[u�J��zͽ T�wUz.\ͫ(*[j�U+{�����)���vE�2Q��4�t��d8C2V���p�Y�H|���%G�Y)��"���%�Sm�M:�p�wk���V!a��UYbu%F��.0�.hSڇ�N^_[@�F�m��3�fJ��ps�h�pÄz���2�#O����L�؄Y�Mx�0F�-�H��M&�l؅]ICHSJ�"΋r}(i��J�fJ�Y}�#�:n���j��3rVmG��ʱdq̭�
���)��.뺅#û<�qG�D7��D��b&��|��[��ت�׻�eUa�^�R��� �
�;���k4� 9��Δ4�|fe��Q������YN ��|�#���"��Ԑ��>��I)nC���������w���|ʎmC�)���q{�ҳ���[I��A�vD,�!x��VJ���j��2�?H*�##�Q�8�V�H~�N%�Iq��d�$C8�#���0��E:n{�#j��h�~�E>#�q���)�bfB�P����`�)�W��F ��/�|C�H�C��TsjOǻ�_���	I3$E��I4�m��R��5��;��* !�x��޻���W�swVP��x��]���{ ����@ �Ө��7vH�=�b�sW^�z��      U `   <  �   �
��;���Tm�T  � P��>  � lT T<  �T�m� vk7{�:���K�=�n�f�?j�l;�U{(
�l �6�֞+m���3s�[��}���7�1�q5��;���F'_}=�X�8�V��X�a�!]Q��t�jF�D�88�V��xwg��#�����af�>"�7=�R�{�4K�c"��t������HKm��He���B4�J�!b�����B,���b���4�~.�<Fݖ~l�䑸di4I�7҆��,�fJ�Y}����t���/��T?x��cW
"ڏ�s�
��"I��l&�Y���ܱ!wRP�`�yB���WҰ��^Z�
�|�s�I"�P��h�J�+wGE*���w{�J�ت��-���VPY��-�i0�I�	��[��!ff>�g���rm�S���v7"�:}bL���(x��ДF��۪%���ޗ�ſe`=Jz߲���[�[+/��!f!�2�!=�A���$�uM*hRM���x>�*�#x�2�F�wu�F'e���O�����?C�5������JI&���p�d����"0��(/uL��~�~B��!��6jf�"�:z�},Ӥ�i�$��X��IC�)�q�go��W҆�����d���j0���q�nBÎF���7�>��! C��J�P� 
���[gFP.�I��M��E�ٹ+v�#Ƕ{�Q�׃�(؄a�IV��7�%F	v�f�~^�y��I���QJ@�j?�;1YHf���.���>#��!oү�\8D7�~�De��m���I�bf>�!bu%&��X�o��1o�_3�쫣x��[+��Ii$�U*n��ȅ�p��Y}Ւ�#Ƕ{�Q�י킬B,������܇\'���I(��F�l7W�F��¾�0�|z�ԸB2V��=���8G���S(B4߿��_�w�y�x�z�U�ߵ�QU����Ŕl;�U{&ʩ� U y�����4�m�UI"Cmиl�ojM�����X��
������0�:�F����?�{���NF�JI$���Y��՝j0��Ys�%G�l�5p�!ݯ�X�a���mWʓ��d��U'M��(x�/(\6a\2c
�P�!���R��[���">"X;�M�m�"��D-���1>l�_h�m1��3��[lķ�٘X�]ICHSJ�E�re�*��ۉ&ۉ�'/!�8����F��/u�D,Ä?eά�!=����v�㸒	(�(6ST(&�UT�6���oh *���U�ʹm�)Y-��Uy��&��I8#Ǐ��X���(B0t��p������=׍IRf�yH�Rt�UT�M(�n�L��n��\�c���q�\�s|ĆS�6���Q��:i��.�q�r�tٯ�:�6��b��rO0}�RI��$���R�f��I�:JhD�I��e�(g[�2{��@$���Sm�M9Rf�{mL��n��\�c���q�\�s[��(�):��I&׺X�nۏwF2  l��U*�c`b��vӹ,�ͷ7�e��vn ����V�k�l�R�Ů�:��u�Q��l8?��` =T�w�	�x� � c ���T���극�� ��	��8@x x8>��Մ���g��rp�Q���{ﱾq����.�n�0 V�[b�l��yl��˪Q��=h�+�`0��� R�   x5�
�
���P<���޼��Ӻ�w���6U@  
�A��/Sg�� @��� �Ee d6N�  .`  � ^�)J�@G4�w0 'U<����%�ۓy�w��7��ݼ�P3�Ry:�pn]�{{j����
�l�q<��P�>�� � �wݹ      Ve   �         P          �       Tp         � P �>                   
�� �           �  UY6EP�  U�    �   x@    �        ̀ T    w*�   
�       *�     �| VP*��    x       *�          U     x    +*��  �P      -� U@    ��l  
���mi����     ��
����öw x86�����o�X6]�go1z���g���ujp��7����6���۷~�u�]��ܩS���[��^�J��f���߷��j�M��oo�͑��gU��� �     ��   �T  �u�U�+( �`U  ;�U6���� � R�PmW���T�;�V����l�����z���̷d�w\5@*�pz�J�� AUw�k��5]�$�l�N�~%��G���E�
d���|�����&����=y���x����I��h�e��[���ƮD;����W���!wRT#AyW�F�8�!�&i��m��j�b��Y���R��[��ՈpÄz���eB4���P�l�w*�H�C[I4�T�m���,ç�HX��IZG��pلYл%�ZD:o�]�%l���DYe��m�çba�e��%B<{'����x>�*�a��%�9��q��� ��R$��x���;����m�p��d��6�l �m�.�s7��U]�￝�B4�2c
�V�^Z�FJ�P�綬C�#���c�fH�j��m6�`��\6D7�&�L�"�:}bB�*�J�<狆�"΅2Q���C�+�S��m�RH��"��[�θ�,Ä?eά����cw
"��}�U�0Å���M��R��m��!wRW�����f��&0��a���p�d��{j�8a�)�@Z_�qI$%��L�2��ˈ�ཚ�q�!��6j�a��!W]+H�.<F�6�)t���(�OPvv��� �b��E��6Ք���m���a"j�I&�i6~)4o�i���p�d���q�Y�~2˝Y*��=�\(�wk��
��M4�U$�I
IѸFp��h1���:fP�l�4�d���"��.�����^�J1$l��m�&,|x�����2�lN�!p������E�t�^.���(T<�LE$�"Tm���fg�L�nJ�!��U�p�2V�θ�,Ä?eά���:�'�$�Sm��$ڸQ�׃�n�=�l��+������x�sf�2�����wm��L��/R�eRͬ���q� W�T��� *�����߈�9$m�[m��Q���[�Q;~�1�3�k�������}�����s�|�f=dt	�I&�m�����Uԕ�r�.0�:�F�"/�]�%ORΌB�6C�X��
)�A$�m��f�ڄx��cW
"��}�M�qǏ�*�l�wY����s�xۉ�������ۊ$�A����8��>�B2W�C��ڱp�2��Tʄi����q�8��78��Y.5rI�H�E�t�ą�U�J�<����"΅2Q�+H�K�WA�,�[+��ԕ
a+�Z��U
��wq���w W���w ��P��m��U*J���ba�e�VJ�x��cW
"��}�U�0Ç��A�]�J�sdύ�Uz���_$���#L�f0�J�!�ٖ������\�ՈpÄI�՜�������rII�Ē!�l�ok�t��!�p�ą�Uԕ�yO�E�
d�rV��r�J���F�T�m���,�^�g\ba��eΩ���ƮD;����7�}ǄK�N)$��N(�3�x^�pلi�.��U����.���P�綬C�"�M�F�M�(�Sa��f{�� mƀ��s�4�*���
v�{N��5~�K�J.R����ٻnw [X� ��Pاz�W����Oe�{�z��V���;�*��     .`   <  � PU m�q� 6��UPuP� � ��U   *�m��  ql �����S��WQ��E.�J�wX(Y{n�J�J�����6Ք�3���/j�)E"��C���������C8�s�g�s��a�L�[W��Q���	��$�nFĎ#��l7}��΂�e�=Sk����p��T�<Q%�7�I$����#�a�R�.�B0t̡a�#�La\��B9�}��m_j��&�TNIM��wV!����U��4���U�dC{\�xC�D#�Z`��|C߁��I"RuUM��]%���GK��Y��d��"!i�\�M�#��U�m���^�qz��]�tm���Һl��U*���
��w]	���F�NIM�rgG��N���G����(1�IP�eXg��!�WܼG{�!��X�n6���Hf��T%�mX�CdN�}S+��c��W��G�>wdY��R����%$�l!����__i�D>�/��H�t��8E���VK�B!�<=0����I�i$QL��ݮ#Ƕ{�DC�^l�|Fg��bu%B0t̡a�#�p�Ҧi��m��e�¹+�u�R��{�ޡ�ڱ%��o��ccڲ�)u�$�D�M$[rm�Ih۹W����Tl;�+�@� `�ed��B6ۍ�ԍ�?K3��Ӫ}�ϼXg�g�GF�"�S��{�z�_�k�t�M��aӱ�\e�u{�#M���8�8���gl)#ڹ�8�W��A8�1$m��l?�HE�x�21�}+�u�R��{�}B	����q�:��Yʑ����R�"�m��m��dC{]�>Nȳ��񂗊���!�C�	z#���8�Y�k�Q9$%�ɑD3��j�^�b���Xz����O��;���r���1W��H�m�S}?6��r6I-AKn�/. 
��*���VPU��l�uU59��P�����o���}���#:G��{�<��qH�4�wV�'o�8�0��
7����i6��꽯���=W��vt�?��'�X��Z�j�!�!���KI(�nI#rr#���z��a�[���S�,=e��m}����DC�R^�*#N��$�n7 rDs�۫��������g�#��{�<ڿR,�ψG��-�C�9Q��RF��L�O�E��,���[�"��{���M�/���7m&�e���M��mD�<mlN���� *�pR�T;��;ܻ���	��H�*6�gߩ�	���R/A�a�[����!a�e�_����^�H$�Ĥ��r`$S�[�/Ds��n�b
f-��w��G����yj�H��Fq��m�$�&�HGެ�=�<~D{]yW����l�ok�����g!ȕQ$�I6�B�H؅]I_uM,3���&�WЅҝ	�a�[���S�?}���M���m�[7ޭ��O��;���r���1W��۫����j����=@<8?���b��m��	��^R��C���P1�p�؍�+u�����cu�� w7����ٹ��=T  l�*�uW�ٞ��N�ݯ������^���jT  @   �  U <  ��  �ATGp� *��   � ت`P�*�� *�U*�
��C{m����<w3n���Tw��n�ܶ�]�ޚ�7�@�w
��P w U��m�����mƒQ��?w���G9�i�AH�w~�e_�`����qϖnS��Q��D�j~Y����L�V�گ�t�~�^�����w�BR0����BI#�m��mH���Cd/e�jm}����DC�]�瘫��C��� �b�~��G�H��I$�X0�;E�@����W#���_m�GGz�,��ٺ�F�M��i&�"IN���N
7�}��k4n؍��ڭc�F\�E���Sh�U#����T6�U]�TUj�
���Ek�z�sml �f������������o���{�;te�#���}z��8���d99��~��E�n�H¹+�G6Կ����cG�UXM�\n)nCC=�<�x���g�g����~dC���)X����t��v��"6
��"I��r	$g;��q�:�}��T��C�x�\ڛ^#�l�;��w*>�4����m��n�N���m\��1w.#æ!�z�z����,��?#����ra��a��z�9��;>��R��)�� *�pz�J���z{*�tv�i��S3����D�����˹�ݡs4�v���|I��%��Q���wGttnJ�!,:�}��ԗ�C�|z�.�ik�&��a'$�&ۍ��?���h�����m\��1P!�F��fq�+�XD#��I"[�i'#l%���|�	��G�]����4��~���^ӝ�2,���:�I�I��M؆���#��a����Ѿ��B:`t��՞�.1�q���&�-�Q�S�H�1&���7m��z�@U�� VP w��@�H�2rF�n7i8s�{�i��p��w��_�Y�uD�.�J�`��1�gx�h���a&�m�Yi�}+�s���GM���"�:�]ilt�W���#�I#��M$�7I�o�DY�L��8x��K�����p�#���gN�%�)S(��m��t�qp�:���0�M�|h�6e��4��w�14�;��>�H�J6�&�a�<o�G����e!�?��v
E8E����a��W���+@��Um��z޷@�m������6¨*[k��+�9���%�IH��"���ߧ����V!��H��Xg�3�F.#�*p�c`����fF"�a��X4�8B�ݕ~,��>�q�#����u~#��r��G)(�nI!�F0q�O�1��b����l�#�5/�G�H��"�!=��6qI �$��/�ޥ�뗕~x�~w���M%������{�^�Ν���(�n7!�㹿h��>�����b�Z�}��zSe������#ݎ�Y��vnk�=UD⫏F�<{��{b��ٞ�m����wV��U�m��az�x� 75*��n+���g���V��We��� `   T p   U  ;�@ <��`�;�ؠ�� T� ��*����T �l  �`<*�����׫�^�ȽoG+�@;�ѩ�̠+�U+ԪU�AUݹ-wM٠�U(�n����2�h�6�<�<o+f=N9�g7��g�#�5/�G�v�戩4�%��)4������ ������*��1���&��m�<��2�ǎeL���9$I$�m6pC�C�'t܇�q�D'�N��o�"�O��|�L�#O��1��I'T�i/�&�"{�y�龳�n{՚6cnec,�w[1�z1��X~�J��0]$�m�ZI6۪I����IB!�:��\����e�^6�����[��=��X�]Q��k���c��e]�{[l�a�^� � �Usl�{Wu٪e$���n,|mZW�A���'tܾ?��9	�aӿ,��?8E�r��L�a�ےH�qf����&R����G4������6�`�2:G�ߞ�z9n4��4㙵x�'>�B>;� y%�8�;���\���\6G.>"2�MS	6�I:��~kO�j�(�W�ܦ�ψG<\�\����b!8�:w�{�J\��6�m��Q���6F�&U���=&۾4G\⦺>�;���m�ϸ����9'��r6�n6����Vz��
��UU� *���
��֪3DID��7�&��ݑ���$S�ٚ y%�8�;���\�6���$�F�m�$�g"������a^�U�p�W�ܦ�ψG��\���H�e�R|J%$�F�0���|����f����&R��S;�i�!��惊I!-��qF0S�է� �x�=ޏ6��d��HgNmI,��ȅ%T�N���e���7u�6w7�x�y�߽�[���G��;V��w�C�3�r57�ځ"��h���5Tuf���P
��U+ԪUWvP
����(�+ݚ�ۍ�\�e�����N#�j�_9�i�>��,�<����d�Q�w���H�JI$�r�{Op��6�~����=���V���_��mmϓ�*'$�&ۍ��g�L#�y뼮����U�i��}�%o[\�V>6�?��)#��@��-�Lx!��#Ҵ�=�%�㞯gb#h��4�- UJ�d��m$�rF\�)DS�xN��{Op��;U?�p̃���x�z<ڼ�aD�Ii�ӄZ�6ۮ�g��]�{�� m�p{( ;�*�@���ڭܪ�	��s)�����wg�L#i��Ť�9W�K�>���l�NN�I �m�!��>6�?�Hg��:��=���w�n+���m%��ۍF�h7����Sf�}��;Op�m�8fv��8�.%�I$��{��N)�����K[�(o=ߞ�>V,�=�H�4�I%M����>����k���۝Jy�y�/=_0��eo޽���������m���ӽ�̞�V�r��ӻ+�Hw<;�[`p����W��wN�1��7f�t��:ٻ��زT���P�Wu���Y=�ww�ݻ��{f����T      �      �    �6���� gp*����� �  @� � ��C� �P�����N�=�Mː~�QYV�r�V��o\��m����Q�ATwZ���*�^տ�~w���3�_]�s>�ا]�a�f龤ι�
p�?�PN%�zF�Q��'���=������~"����^wX��5�|@�=���$���#���^?fd��#��eY���+9��S�3����Ll�B[l�YH��v�v1�#���W��|6vG`����9����o�n4���$�
a�@A�I��a�N�G��~������4g�~$}�#��m���e�̑7[����g�� C��
�P� 
���g,r��Lꭵ�{����~����U��x������s*�x��Y�ψG�R���16ܒF�"��Ǻ�|E�;�~��̋��u_���l��F�weL�eD�$�q��#��wǨ�N|���'���;ޏ7P���>!��~W$I�#q)#o nO��j��{mOs{�3������@U�X�E�N��m����B: r;�C�s�#��,��?B=F�Y��/��T�E���k�m�ի��sf�{�T m�p{)Tp[hͲ�ۺ#I�����H�g�>�U��81�����a���0�6�<��
�>ȋq�!1��$�RӞC��v̏i�-=t4�������� E�~䪪2�n5m�[��������}?i�Ör����7�r��:}�}}!�!w].[��ܒI$�Gi�!���}�#���fʳ�0�a������0���-߄�	Q$�%B�r<���>{\�ӄpW�c�Fh>��� ,>~�F�;�����o�`�^:̦ۊ�@��ٴ�PClUW�Tm�PUY�ճ�9�R%�a&۪�Mp����*�8t��������Ȯ?�LW��g�j$$G�m��jEX?B;���L:@��^�S�nw����:�<���=�*�UU�M��!J��z1��g�ܞ����M�ȏ|u��g�4���m�UI�n�Yp������X�:~�5��}�r1zp�9z@�5M9M)$�0����<t�ܹ!�Z-��0�{��4�4���>��!פ��6R�@�	Bdf��8��1ֽ�u@P�*��ت�� �-���N�������f ��N�O��A��a�dƮua�y8����Ё����gs	��Q��Q��k)�CO�7����㧮@��f��F�B�uVw�!�W{�&6TNIM�p������1�a�ܯgb#xwe^�b��}�)DS�_x"��"����I$0���!�=�
pک�����=���X~N)|B>9�
����$�n7��L�!�w�z{?�}Vs��S�����8g��G��z+}y{�w�s�! Ͻ�����k��"H���$��[$D�ل��7*DI4���6����[��I]�"'��������|�6������������|�N��;?o?H>|�Z?�� BA�� BAo����/�^��w?�˗��	w�?�붪���?]�/z�:�U$I��"H�B%HT"ܤD�<-��[�@���������o�H;����q�Y��rk����9�H�h�훞=�=ΊA	$H;]��H! �}��bH6i�v���j�����5t�kz1�j�@�������|?�ݒ$�1��׫ەݽ�H�{�{$H;�[�:�6��U��������ƻ�7���Ӈ-�$o��j�Z�g��<8���qt� ����~i�~�$~���Ǘf�/�b��L��U�,�k/� � ���y�߾�����                        �^                 ��                        �         =U14ST1�P��a� `diU��1hU�5L 5CT�|��^ZUyk��
\ �Ю[�� � S��aA�Ҁ�� 1 �9���          xK���U*��P��UK�UT�کYi*��J�� �����J�f�J���U��T� �T�mJ�X�u�\l�����U` n�W-Ҵ�;t�U�j�VZ�U`          UJ�l
�w
�R�cj�S  ,�������j�XڥUb�J�  f�Ucj�V3U*�ҪLMU0 �XکUc5U,mUR� 2�U1�UV6���`        � �U���Xڪ����Ū�� j��-P�T��f��b몕� j�������e�T�*�X �iT�j�U��UX�t�\Z�S  #D�-R�cj�SU*�Z�V  t@      ��WM\l��ciU,m�UW  F����@b��X �!��Te��Xڪ �X�S��6������ -USb�ceSR�� } j��M�U$ i�  � T�4�x�US��@   �!	��S0��iCA�OSA��<�T����jR��a  � 
���SeUT�� ��24JH2�@�     �N��u�we�ݻv���v�g��(jp�u(s��*�,�"�e(d?_�����TEc��<�"����	J���4��O�ɤ
O�'$�����[��'�'Rs���
M!�r�@<��<�]u<�B�@�%��N@rJU�k "�Ty:PF�DM(rN@�)B ԉ�@�*���B�' 4*(h4��PG@�� �*'P��P%:�� )�Ҋ�4 �u�H�AP(!�@��9 �l���s �r@�aP:��4"$��P�Q9"���(�R(u�WB�+��?�����{��m�kb66�ƍ�EmY�U�)���f���jI5�+b�1E���dhJ�
X���E	BD᭤�4U44%	BR$D���1Q��ji��i��])�J��)��J��)�JR�J��R�)��J��(J��J (JR�(J�*�iJ�)ӡ�*���b�b�ZV`��)�B�(�( �(J��) (JJi��)��(�(J��� �JD�H���R�
�J(��J�i)��B�:�� �]�#B�LF���N�
D�� �t4�R�R��f�ESm�bi��&&�4RQTDUMIL�TD1RP�IBU,�UE�R��h"���E�������������f����Q5�Ԗ��TE-%!4��R�ET�EEDkkkl�)�m1�b��V��0SSDV���QELT�m�(��B5X%�1��h"*�b�"�


a�1D�URARC�b�&�jh���LUE�b(61�c1��I����h�f$��qSh�"��'E[E���D�TMDST�M5D�S1A[cF�3�,�h��f�ljƚ
����b ��lL�l�6h����V�F��Z�mF����Ӡq(&��D��D�Z�N�H��� �B�0c)PFPJ J��J��(J��(J!(M	BhM	�(JBb��(JBhJ��"��(J��(J��J��(J��(J!(J��(J��(H��(J��(J��"��(JBhJBhH���hJ��(J��6�P�%	�4%	BP�$BP�%	BP��4��$N�4&�Д%!�UC��i���%���!�(t[bJ�b	X�B[	�C�1�bt%�&ٳ�(J��"��(J��(J��J��(JBhJ��	BP�%	Hm��(J!(J���%	���Б&�BQ�Д%	BP�:t$BP�%	BP�%	BP�	BP��)V�BbhT�R���R�B��X�4:��a֝.����C���(JBb�ք�(JBP�&��BhM	�4%	�4&��	BP�BhJBhJ!4&�4&�К��K��Д&�КBP���0hJSBR&��(M	Bi����&�-	H����&�J�К���QT��D��)КA�КJ	lD��BP�BP�4Л`�КBP�h�"��$����h��T%	H�iJ)IVqF���k�Em����q���u�u�]�F6�)j�Kd4�5��h�MTM%QVōEFةE�՘��,i�I*�Y)�Z&��ͣQ�[i�ͨ+h�Q�5��)6�Ѫ,�U�,Z��5i�ƍV�Y�i)�1h�4R#��-	JБAB�R�M4�E3҅ 9hJ��J��(J��(J!(J��CBP�$BP�%	BP�%	�4$BhM	BP�A[XJl&�КD�4%	BhH�Д%�N�К
u�4%	BhM	l%!�(4%	BP�&��1	BRE�&CBP�%!�uI��V��3�&�-m%bД�RD%	BP� 4%"D&�КD�4%"P�	�4%	BhM	BP��H��D�JD�(I�Д&��)	�Д%	BP�%	BD%	BP�%	BP�%	�t%	BP�%	BP�$BP�%	BP�%	BP�	BhM("CH�%	BD%	I�Д%	BP�%	h4%]	BP�%]�b��Q�:4li����֜�M�ZH�4Um�
)b�Z��X���4��M��K�(Ka(J	�biBhM	�6��PiA�)�4&��4$BP�%	BiJ(u��4%�a4%	I�ѥЖԴ&�I@V!(J&��4%	�B��K�l�E-	BP�&��(H�К�F؍	BhLBP���(M	BP���R�4&��4%	BD%	N�BhM	C��Кl%	BhMPH�&�A��Д&��4%	H[X
��4&��4%)�(J�Д%	�4%��LI�4%44%	BP�a(J��4&��4%	�&�Д%	B[!A�EmA�DBP� ��eWH�H����H+mh4
�SE Z6ؠ�e�P�hhF+D`Ӡ��J���)%��t��)-A4LZ�D�ӭ���# ��6E�ZQ�4ꄢ�mX-KE1ih�@U.���u�]�U�Ah�kF�1��lh� �YƇ6ڭ��E�b5X���� R��h��J�Z������"���t�Z� ����H��dt)PM
s;�AS�̘���l�l�ZH��4�J�&�҉�"J"t&�V�Q���bV�i+N�e�i"����F�4&������5����u���֭BQU��*�10Ri(��Embֈ�ZMѶΘ�$:)�)��(����f*�j�P[cf���:����mUb�ͳEl��
j����b�.����D[f��Qkl���1N�E�::t:ƦvuULU�HhMQ�N64�&����M��ڂ���#l�&�6�$EU
a���TQ���c5:0Q2D�QT�QTT���Q$�TD@[��:�Zr�&���T�*�������L��PI]]��9�������ܣ+훟`"���{�����O�B����ζ���^]����e����x�����%_���77 �ּ�9^������   S����T���     �z�{N��k��� �	�     �  �0    <  �1�p� 8@N ��    ` < x �  p�  	�    =�0�    �  N �   �'     �T�8@ � aTU ��� ���VĆU8@�*z�'
�` <U< ����� 0 ��p   x x     8  �G>�< < �    0	�    <    �<@N      ����   ���	��   '   <  �    ��	��     ���    �
�*��p�^ U	�V���UU@	�j`    N ���� �� �TN
�� 
�S�	®R� D�j� � �  ƪ [ �U���m�]�뽻�����i�U6l�Tn%PU[:�e���ѹ���n�T=β�@N��@8@�(U*�۽�֠y�����o=�3�*A�9;�W��y�aswcf�l趁�y�3lk���+5�1�kj����mmɴ���u;^��nomT��[
�ӗ{����qs\��Ky�QoG/w�ۛj���Y����;YS;��nUջ�6�Y��[�+,��e/R�0۱��   �� �\�Im�QW�T6���< < �@ m�6��
��n�p.�T�� �p0�9�+y@�8WR�@x8w<�8EP�+\��<  �����P3� ���=�E6�P淳�ܶ��h�����C�n�z�Q[��6���k�����²�9��^���t�S��6�p��4����>+]���nZ�t�ַ={^��ֻ��yjW��VvQ�  �N �G>�< < ������`A�Pp��m�t��
�<� 8A{gs�8*� �U< y����1�N^�Y5m�G��J��ŵ�p���\-*���gͷX����a��;ú���y�e����f�V�����	Znկ.�y��W;leo���w;r���R�v��{��os[Y=��Wz�����v�w����7u�[eeof�T�{����6�ݻ�Z�u�ol�Y��fѱ9Tཌྷ���n�kg�����Ä�Uz���Cl-V�ج�U�c   	�ms�V�[/E9�v�mK�������a��]=�SV�������B���
��� �wVy��  ��VҀ V�Y��eTR�M��;�)[[�V� [-�k��T����Q[����Q^����
����c�t�;۷Y���4�Kkg�[������w m�r�0��v��YCkksn�J�n� n*ʝ�岅�S�ު�������lb�������u�v�o^��Ԧmns+k���+)[fmJ��v���i�@[!��;յ�­�wm��QŲ�B�fr�U,���U��l[Y[i���.kd�3��l�ی�M�v*�wq����������j�
�\�ͩ�UY�vv�mn��
�ٵw6mom��wr���slVm�[v��(��nNZ�f����]ʪ߮�}Wu[%P�U����V��n��m�-�v��ۜ����U�V㽶���ܝ���C<ɼ��MVn�[F�m��w��]�k]�ѽ����:�{�t�iUZsVɻ۝��Z�q��۪�g�=�:�k��٢��r�����'�U�R����l�Ų��e]Hv�̴�m�]fWs�]��^�i�S�ڶ��m����m{�m]�x*4�\��t�xrIRHҴ5Q��bGUy�ؠ���wOv�������m�7��o]:wow�|��gW�fU�{Y��^���������x+u������w����N=�Uwv��T��T��]qn�ٍ^e{�^��m�x�r�+�q������-\�o~�����V�U�y��q{e�ړݹ��n�2J�_�F�S�����V��Um��J�:�����Un�;U(kJ{k�m���e6��{;���-�wZ�u��z��w�{x���n�+f��uǭ����,ں�S�s�g��oX�9�ooo]޽���Ool��u�j�㒭,l�	�T<����]��;Ni��  �����_1�zٻ��9�jg���Yݦ��!Ν���v����nֆ0                                                  C�                                                                             ���                   U                               UT
��@     *�[ B�[%QR�  V�M��m��  @��  0                                      *�   �>�  *��   `
� � 
�      T                  *� P   � j�    ���u *�         �                                      p� C�    �              ���   �       
�  U U   �  �        @ �[ ��*�T�  T�EP m��        P *�    ��j�
� 
� P 
� �z̴�n����l�P 
� �
� �R�k>�����ʽ��eN��{MN|@                   �                                x           �   
�         R�     �}     �     �m@�r
��
�เ �      < �         <    �             z�[  p�   �  �Wߠ     �                       `                           eU  �       �Wߠ        
� �     P�m������h��2�*�*��}���     p���     Pd ��               /YB� �    
�� � T �  P    �� �@T      �@    U*�                 `m�          P    @        U   c  T           x          x               �   *�                         ��Y@              �6�   �   @          n=                �@ T      UR� �+�U*� �>�                    6�J��e d *��T  �   [%P  T�ݮ�     �V   *�  P�} � �@V[�B��     ���P[!:������;�+ң��Kgc�x�l� P*� |��PP�U׭<8S�s��6�V�
���SsR� @l  @    1�b�UT`)S���|��ձK�Y�����g���8)P�  �ll;�VN�+@v�2�]�{J���w@�^{�vپ����N�۵���M2�M2�<}=J��R(t�2�6xH��;�������O_?4�����?����o������ ؠ<v��	�   �`U �ǀ@PAT�� � �TN �  x x  c ��o   Pm�yPN W-A�� ��jU6��8�yN��m��U/So5�ֶ��-t�6i�7{���m-��� �P
����� <U�1����l�UV�)jn���k	��̻�v۵�^�UD�Vے�yT�ʂ���Ik� �v�R����u˻G��[�מ�0w>
���6�˻�h;ݽ���uͶ��J��@��]yle��Ÿt��q�m�W��y��Qm��J���\�1�ڻ;��*���w"uU͵fI�{���b�k�j��-��v�UU��Wu���d���f�x�E�R�벷��5��ӭ�����wͲ9�w��mn�*��׺���Wq��;��Y��ϛ��aj���x��          �               �            J�m�`]�       T U  *�    *���(          U   �   8 ��T*� @b� �P w��wns@        ;�   �    U� �l  �     
� 
�@          � *�   ���hU ��   x�       ��      
��              �  �   �@  w  ��P   AT 
�x *�P�P F����-�UWn��+m@ ��ml�q9���獲!��_�ٯy$����)!$��7��qT 8@ g�Rݺ��{9��]�e�=6�m��
�p�uv�6�wk�˻k+U���V��i�|PN���ݻ�x�0��vզm2 
�  �  \�`Y@�� GpUP��UQ�eT 
l  �5ٙ@ \� P 
� UF�<���m�׾{�ᶫ]|�uV���kzݺ���u���UWu]�[�j���UUVڪ���o�z�����H���i�/;�S0u�}�́����n��٧�T�țrI`t�_��*���k׆�1�K�0�s}�X�دC=���m� F�
i8M��s(��>�a牞t�{YA�=L5n�����Sr $ @)�o�~�3�����OԎ��>���s���u�S��� pa!�i�S�[��>�є��^�m�����m�;y�=?d͒I$�E����٥KֶM��w�lb�׺ U��*�W���n�v�uUl	(�3ۋ~�l>�����yk6ެ���V��^k�^L�Q� ��oy�ܿ;���v�������;��E�y���t�d  ���w콻�i����g�<��ҽ��Qf��py>��� �c�������z>���.�ם.�r������I�\�$����ܒI#D![=�{���ߪo����?}�~[{v���ݟI*I$��7�{�Sa�W��7Z��� *�qT�� @����s��]C� p��罬݌ə�͸k������{�[��F'zG	#llr�E ��\��c{t����/�u�M>�l���׶km/�JI$�6��Z�mn'X]{��+��o�?b�^�׫���w�mh��S*F�$�2J�ykoMu�׻��3>��{�e=������$���H� �R)�V��[��n�{z����׻�z�ſ\6���I$��n�v�z�W�u�׎��_3�� 6ø�� mdf��[sx�ʛ
��
�=���e�x{�O=�M�ݷ�m��w��o�)4�I`i��；u���o����n���|��/�cN����H0�/��k4�f��֘�9�X������n�}ԵVI"�G�	%��een^Zٺ�M�3O:��/�ֽy���=
v @Hl~�����{�f��ȏ�c��ǻ��~�ݒI��6�P��U{{;�ڴ��^���ª�T�
��-�mʍ�޵�ƯUR�E�o�|����{�z�{a��1�\�\�O��l= @$Hzg���Ǹ%f��+֯ukؾ�k����=Ν!� 	)�y�ʽ���?|���߱��m�?L�&l��xϳB�v� ��=�Lۆ<�۾�c�<���+/"�{_ly�5�o�!��$�"�^_��}L���\6��ܼ��ukɖ�=}�������0  	��8UC�٩��GlNm����N7����6Ք���kh�B�j-E�(�
�8#
�����s�λ�շwn����kv�ds��       *��   <*� wA8�l�m��*��U@V6�  �   *��T P}�� �[��V�_*Ӯ���� n�����6�w�7o<U�ה C��/UT �AYM���:q4��d�� �B�^������L�o��yz���f����ץz6P6��H�HV\ǻ���Lۆ<�۾�c���{�����}(7*I#cq�r����nnOm����ž�l7GX%{���v�қ���"߅����[g�u<ٻ��\>�߾��=�߾�k����$��	 �
~9�o����n���/�]4߸S�]��x��O��I��$H���TS��͞�k@l;�+�@�R���l�u)AnI$t�)ｾYok6���Sk7g�׻!�3ۋ~�l5�����	$m�I҅L���ukݵ3LA߻΋\�7�1y�����-0���N���t�W����4��^���Y3��C_��͍:T���	$m�] UZ��i\�=x[ڠ��*�)f��/w���t�nP$ ��t��'(>����xo�b��tZ�7vUd�P
D�I�)��H�;�ܧ�t�`�V� U;��*������@��	$QH?�~��{^���z����~�h<ƚn�Ww[g�*��� M�{�e�yg�OJ��ڛ���;͸��v�>��	�T�Ѩ���$<�g��p�kה����/-���k/Ku��}3]6��( 
Is�{��^��]��֞=��?Xھ�y�
۽h�o���� I!��f�5�����0�>X'����o]�+�������� �_7n|�6ymof����� *�qUS�T� U�n��� � 41����^��3ۋ~�l55����]�Zo
�� �%��A#�������7L[��+��{{�=�~ח>�e��P �T �
�z�vLϪf�5�������yZzV���4C$Hlr�B����i�\��oV���/�t�����K�L܃o�$$�$ �+m��E�~�:.�n�����}]�<{�+���5ק��*�y���r�;2� ;��*^� �
� N7v�̽n���d�i����36�z�vL�ʽ�����?�ٳɖ�$D�% !Q�IY���k��޻y�=�{�~���[��CZ1�F7 $J�_gav�i�7α~�:.띷\]���f��%DRI$����N!m��,�h;e�u^�{���v���)�P��� P�Cטk=+v��ޅ|F��Sk7fMۅ���5�<m�@  ��  �� 1�8��+en�����v�v{Y;�ޭ��Qά��7�P�;�/m,5�v��VzS��x���e��ӵW����[yۼ�       *�   z� � U��6��� 
�p @^ٝ*��6� G � C�PU ���sd^��{נ w�ui{�d�۝w�}�����w
���U1���YJ���[�Z��DI"P�$:r紡]���wun�L��l��k4͏v��֒�c�D��9�^�=,�߰�n�x���}>�L��_�:R$�$�@�W������b��x��t��ߛk7u�n��p $.{v��ͥ��}kf��Y�����k�xRPI$m�6��b��z�}����Ttn�jnlu���!@I$�!�~��u�{���{|fP U⫽�P� *�qU�{���n�PVk+����~6�ǻ�����*=����km�_5>����@޷$�H�ǿ{l��
��}ɭ�'L�̬�d3��O�Q�7�+O�HۀPԄt�E_/'���20���yJǍF���3��♷DU��V���57�lnI$�!$��^Z���
�_Z���m�Y��}p��_/,Ȟ�*�Uyj�O7�S�I"@JL
u򉪵Y�mLZ�U��ۑZ���_-ڿ��V�4�j.TU����}��?`z�����s���n����;�+�@�R���n���D#�����M~�)�[��yef��vTŶ9_!5V��ٮ�yj��-�L`I�JJ:-U��Z{��U�YD7uDx�����2�dx�{�S�*�ym�(a?@r9$�F��*��wz�{�p�����;�볯�p�?�Z����*
@�߯�ݿ���9��J�:iw��W��Zibk���v}�Z��se��T�UJ�%IMP�r��	k�'sv�Պh�>vJ�!G<��aʽ��"E�2��5Y�j�[Λ�$F���X���/��B�Ȩ���t6d�d�U|p�p�뜻�
��I��T��� ����v��ڵ�� ���^��*�� ["�2�~h��H�D�Ǘ��>��<<~�HOec��N�HdB9Z����]{�<�b߹4��  �N�K�QW&���R�b�*��}�\B"D4��
ՖG���������?0$ I�%���^���D3�!�*ȑ�'=.�Y��[yD��Z�y�⍐ 7I�.�5[߮e|��ߝs�	�OP>s��оy��#܁w��]#�WԎ����q��������_�
��h��萜p	$l��k�<��C)�pj+F���Z��QS��)�ʭ}�k}$�I K�k�����x�nݮ��r *�qUk�ȫЪ
�2U�����UYz��40�E0e߈�K�2�g�?	�H�!�>y��+�G{�ߝ^�}J�'�UB�߾�z�b�T��.�~����{���^y�J�#�{��Wμ��zG��W܏���羏H{��0�%{�����~���r<���#߿<
�80 C,_�~���y~�_����|���X_��${���zQ�r:�};�tsпe}���n���|�н���+�盖#��|ۮs���s�p􏒏�_r;ÿ9п{����G�^���Α�!�<��/2?z�瞹+܏�Gܯ�^��z���/�_r>���ͪ`I"@	$u�W�_�~���5_���s�~J�#�Q�u�~���r:��e|�Ϟ��~�?e}����羏B�ο~�~��W���_�-�R���	"�I$p    T ���]��r_�V�V�wYP�mmOn����x��@����{o�󪀭��)֫ٻ����wn<��{��z�:��csr�ڀ      U�   �  ;� �/@UQ��� �U  �P  l*�
�   J��}د ���U[����&0	�;u���W���;�ݼ��M�>����@ ;�*T몺�yU�]s�uչ�9��}H�_^������+܏�Q�W���ι�p����+�G�Ͼ��J�#�{�}�Ύ��W��_�UUn����1�P �N[�k$�A��zW�cv���{6�䧻��\��ԁ$�#���=�۝
-n����7dջ�Ӿ�3/�%t��I �I)�+w��+�����|oL7z�~ϻ�e�Ի^ÑI7$�D��]��xJm�ެ�+S�h��t���"��ݰ �I�8I*$��Tu����o5�ͮ� �ª�UATm��]�Aӓ�c$��$'�w(����4��R�!�[yUc���<-���1xxC�+�m*�	*��d���(S���߫�f�X���݌��ub�7[�;�TuB�6��S������^H�EUUI#ÅJn��1b��ɵ�w�q@{��LX��:$�d�ø�yO�g3gz`�D���;.��H�jIL	R�yH�K�w6���7KyU�4C�Z�϶�.�꘱L��P|'W��ΰ�^'*II%/$�Wf,S<&��Ԯ�@�<v��>�]�!𘶱�$��ub�w[�:{oͻ���ߞ�~�[s;�T�]鵴�˅� �;�m^�d�����H���\�$�$���Uڝ�.i����S,}��������]�)�$�u@��w;�a����IUURI�i�0C�b�{�۪��"�,O��ۢ�_���-�WT�	k6�o��☱w5N��I)jF�ԇC�u|�{�ݺ�1b�!�5߮�w���w;���vh���來�$���0OW��������A�j��uB�6��S�������ŋ�M�Q��P�w�,S���'-�2T�$�H-T��q@�.Q�;�:&.%�λ�WKR,R����p���7KyU�׈xK]��ͪ�'P��\���K֞����U ;�*T]����ueb�UUQ%J���b�3;!A�;$�@��.��X�xMw�]򁍯����^����5��᩽��B*FUT*�I8����,Oo]�t�~�|��ͨv��	��p�|݁Jbŏ��\���-|���=��h�(��)�5H�]���X���������0B����WOOl�-)��nb��}��1Ѣ2UU+$�U����)b%��i��r��gd(<'W�{;��f-)�p���R���C�;�6SRF�ܒI#Dd��.M/&��6d�4{$-iLo[�:bꅷ�@�ͨw�:!�|����`v�1i����	����j���smlv��ֽY a�*��TS��+ڻE\�9$���%TUz��~]7���Uo�/���/ٯ�Ӭ%b�X�LZ\u��
�����9��F�8Gy����芵V+P_f�W�,^U�W�/��O����U�ݞ(�)��I �"HL_�y?�i�WZ���=
�X�m�1j��Ff�b��#��c{�J�@!$r)w����Y�l���_�͘�V*��|B��حn턬Uk*�4�y�H� $�R$U��*��ֳ����q
�p��;C4�<|k.��_/�Z^��-�RI$�I$�   	��8J�:���z�붻���cw��}m}�v��Sf0�u���k�^�魳e�ݣ�=:�qU9kf��ٺ-D�	]k����%N�9U6�       �   W�  ¨ ӠUQ�U
�� m�  ʀ  @ P @ �U�yUU�s�*��u����� ����ݗ�;�l��-�d U�Ҿ�v�\�y�*��L1׍���6Ҫ�Ty��U��_޸^�ھO5>���U���zj�Uj��]��W�#�Y�m�' �I$*����o;��{�!��9��\��)k������0KRwvu��P1O����%I%I$i�j]�'T������)�OV}�ً�jn���1KY��9��/6����-�CE	$�	R5N�(�m�f/�`�Sx���⁊Z�f���قZ����$���'}�׃$���H��ً��fmC��D�>_n��`E1mc�ɵ�:b���;��L]S߭������pk{Y^�*<��˽�^����@T�.[w]Jq��"�R��*���P1O�7�s�0N�����gLR��Og~�vb��Z�����4LR׾�g>8�$�J��	$�׼��ַ�kv�E����]�[vb��	�7��l�(���k>�]�%��k;�mR9*A��E
�k[Q�m|�����X��|�Y�P�qN��|���n��1mc�ɵ�:b���noӓ�������I8�vj����Y����P<�˛͹ޘ'T���r;s�)k�|'�>����@��.�F��*��J�E<��,LR�{>ڜ����L��Q�:�P>�۾�)�y�Ͼ�%�i-m|�����0	*I*3��ݺ�9�v{�>/7��h�ª��D�l�����s��J��UϾ4KS�k6k%��1Lo[{�˪�����}��|�䗛Zߛ;�c�I7$�D�EW(�G��&��zb����μ;�)��7m�N)���Gn��)�>���Pʪ�d����ݞ_�S0��X��ug޹��`[��/�����.(w6۳���+Es^I*�	Q���L�(�?-V�>��8S�Վ�%S��8ҳ�����{v��S��|��	8�#KUU�IQU.��ymc�&��LS��͖���[�q-M��N�u@�>\ݶw��y|��~ ��o��v�m��o;.��wUn��`<Aբ�R��n�f�I%I$�$���k�p=�^����@�3yU�p<�V}��r�S�򛝜�����u����ʪ�$�T���ݞ_��	�r������g�˳�tO/W*o�1H��zV�:|�l�yN��\j�Ti�U2UC�� �>_n��K�"�[X�I����:��9����T�{�:���˹�����UI�*HE�]��y~\�Vt�-qN�2��g����-�V)�<5ߩ���N]�jy~\ͩd��J��g����$s%g {��*g�p��>����<V��ЭB�U���$��n�n������1U^wn�8 6ø�⬠;�EM�m=[m�˕�R����~'���ڇqN�|����`E<����k�uq@wl�X�6�%i���*R� �@ )H�~���ۓ�8D��s�����{�/ny~P-L�^Ub�Ibk��5�H���!&ܒI@H��T����d������-�1~S����^���b��7y>�]��yz���HT�EI$Z�$^5:b�r�8���t�u@�C��ֻ�p��7~�������M����9oW�1֔�p�Q���F�^/*��$�]��q�bC��2��������~�����o�U�k�H�(w�����}���[���\@�����  x 	��8@   �  �� �ªx x     �   �  x �>�8@�e�V�U�⨜��p��UQ�ۺ�n'um�-��e��^׻�:�w��s������^�6�,��y֭�Uw�]@�����VUT�n�\��˛�s��绮��f�k ��'TT� 8Gn���m8*��2*k�ws=�ž/M�)�74��n��NQv㻫sv�ͽ����8*��l�Y�m��lU�ۇnn���y���w.�̫m[{* ��R6�{<��íٗ5U�ݻ*������J��;�n8��޽���ov�׵ޟ��O=ަ���mw2깚��=e-��\f��K��wM��۳=�����T�˻v�������Ͷ�̥�q�k[�z��Wo��������O��Ƿ:�yU����{�Aޚ���                                   U
�  
�P �         @ �     @>���@          �     �  T  -�  �*�-�-�J]/�.��   *�   �   �    ��SeT      Y@      T     �    U���T
�@     *�S�}}  ���    �                  �  l�  
�  � �@    �� ]���TllR�x�G�@j�[m6�* 6μޞɥ� z���7�C�7����}���ߠ ꡌ  � � �*��m�VڝK��Ԫ�c�'z�R���������}#׭mJ6m-�J��y����M��;qƜ�e�63��{����j�]븹�ՠ         PW�  < J�]��
� �R� �  �T  6� P @ �*�� �+ԩe�zAV9��ܞ�ۻ��vë�uvu ;�l*�uTF� *����76�$m�I����I-M[gx�+�Iy���7�������[vy~S�|&l߇��b�Y[�k�<�I$������Ur��'�����)K�8ҳ�����
��C��]!��w~�������6%��RUU+$�UC+���uq@wl�Od���$���ú�b�.o6�z`�D���WOLR.)����kUU$�%I'��>1~P-M��Ub��0KY��l���/�g3�'W�כ����޺iZk��i��I$��I*H�L�(���3gӗx��ŵ���R�&޷�t���7z
��i��������$�F�)��p���sg�u��nq�]��;��{+eT��KdoV�7eHb������ŵ���k��`���9���.��$��ׇu@�-wM����:&./\ۋYEII%N<GLR��Or��Y�_�St��[�C���MyvT��L�u���:�P+<���\�$����%7f/ˏ����⁊Z�s�r���ŵ���R��6��C���I|��[�c���� �I a ��	�������ŵ���Ts��Z���ޘ��/�&�ӳ�u@��k^��}	$�$��q�w�˖Vt�-q~Sܬ�nb��'R2E�0Ť24���0�t����� m��ݶ�mW�NK���\ c�
�+(�
�S��[�yE����!R;�U�ɽn��*�Wt��d20�ĭ���":�pJ�E�wy
 �i2Ҭ^U�]7z����'�`�G)�wxY��+W,Uj��iW
�����%�24��["��ǰ�7����b�Uۯ�MV�Z�f�KΆ�IP�b����mm�Z�,U�ͷu�O�I�X���p�m�G*����JP7C�$��UkwX�yj���wY�x�=�X)�5.�24���~}�x�����ouw6˻�����ª��D�l E�wv+��T$�H� R�]r��QS��s� ic��E�Ǎ�2n}���
�2�㦫z7˥
R�@�L*�EX�ӍD,<c�"�/�o0q��<D���⪋���`2T�Im�82J�#�9_�x�,�#�%7.��_�]���uX���u�r�$ܒI�K���U,�[���_�o�|��ugt�QV.׾Jw���^_gr��S�$��Kb���n��_�Ui��P�8�<V8�>#��`㧈���>���V�k�����r�o� C�����UGp�
����]����r	 ��UT_f�=*�W�b����x�ܲG� Jn]g#���<�tj�rI`
a�j��m%�!��.��<E���Qd a���Y�[ϗ�ʬj���n9(H%�����s(�:@���l�#
x���q���b�|���b���`$ F��8��<l�/Vq��T��ip�$'�b��pU��T�Դ(:@ H�B�Z�U������D�5%�*��I�6���bz�!�Il�wwj�  =�   1�*��p��ov A�����6�w�'�����s��lw{w.��Mڭ�N��]˸�6�8GI��У�j���Sm%+�      6�W0     �� *���d*���T c m�� {(  �� *�T  ��j������V�7  q]Fݚ��׆v�_-r�.����Ve};���PTw^i�����P 6�ڪ*���K�����//���> Sk([8G�­�40:_8�ڥ%I7�8��UE��w]�/,U�$�՜@�9�[c8�#��5Q�ǌT��qEP$�(ZU�ʫ�ޅ��8�$�����:�X8�<Aw�yb��t�"_��  NH��U�襳�wv&_f��%v�j�w�e�i:�
��J ���k#ܟ|n̼ϻ��<�v��<gז�{�$r9$�9}�ݻU���������l� 6��J��S� AZ����cm�حf�d�\�H��]}ނOb�/�Ի��;�'�?���G1��2�o�+�W���2e.�y_Q��g�݃])5$��q�t̵��B����~�|n̼ϻ��<9���rnI$���$��0��5r�"n]u�zI���r��S� ۀ@P�I;}���v�7��}�>{׻���������I"�I�Z���Y�^��K:�k� ��U��eT�UQl�]����ͻ�W��^e=z[YA�v�SA���%���;{�͞)��?d�6�lRG׶�*V��"��m\����˧m�cAS�pnnI a!��?9������ ��x�騦=�J9��.�����@ �A^�r��Y��,�n�fZ��j���ul}�t�n��
�d U�������z[OS�e��5��_nz����I$�IR�ldI�Aֱ׻�ͷg �w�ԪU� �
��T�
�R�@	$�3�V���ح���=m}����w�^i�n ٞ�%�oo=�#}�omf�u��>1�^֯�t|��T�*l"
�B,�����g�t�Ռ�և�lE\�"*H��"�,�4�J�UUD �ʺ���]}ޅ굪�Y]�y�:C>�fW+�F�t�4�����m�e&���$� �_/-U�폧,!�{	sVB4����ذ3��!6��j���|~�͒HE$�T�"Cu%�sed�����l;�U|����P
���J�cA$� ��z�u���օ�,�g��X�ψ�=���W8ϥ^�U���
:EJCc�$�񑅛3�c�,���m�3����{оB�^O�������w͛�F��HJ� W\�=^T�~8���ʾ]N��d2�`sn��E�Ł�,�[zWRD� I$��W�֪��}R�3�3� ��e�{Ձ�,����5Z�V�;�PrH$��8�G���R	J�Yfa�,q��2M��Z�_,��j�ڹ\�I$� U�  x8��r��u��ͫ��@��a�n��u^�����v��N��O�Y^��m�ۋ���v�8������m˷�O�>�|�U�I�ו��       N�   <  � U��z�
��;�
� N6�  �� �*�UT � ��x 6�yT^�e���k�|{�oWO:���׻��� d6�U��eT�U>����|m��*7$�D�D�ܫ˗���:���j�Om�c!���Ըp�Y�%�Y�Ϗ8�I��A$��(��֯-^T�^жp�U�s#��b��=�m�0��opW��*HUA�øtda\�U���R	J�Yfa�,r��]}ޅ굪�]��MӒI$m�@H^�|��#�R�W�j�{څ�a�!c��d8Y0;��D1K�K�� �I� ��W��|�+~�DC�!tZ���F���!����[�UkV�����I$��Iw��͎�ص�lV� *�px+Ԫ w PUl���75]�Sj�Z!�"C��l�da^�*�c�i�RR�Fu��%�1C�/�2�M0���rB��U|�����Y�|Tr����Ε&�a�dCHNz��E媾]�lt�PI@�It�{έx�{V24��C��L�!ӱx��S˼�Uy;�9��\�S7�=%  ��*��嗽�u�˹�*��g#
�W�8���J�ʍ�0��tԗb�T�8D�J�yr�V�w��� ���'j΋�T^*��X����;ʥf�G:�?{�$�J�I	��\�lw��������U�F� *�\�jW{��hm�]�od:Y�K؆6��Ռ��Ϭ�:��DC��[P�5�24�Ei,���!$������o<GWXJ�V�g��X^5��g#uW�*ug���\��g|EK�7  �!_*�LהӒ���y&جf�_��>�>�q������C�ug"E�����Uyj�s4(Ɛ68���/�i�C!���.�/bD0�&{VB/S5�3�9��p��9�P[R��F��(1�|�:�^O7㊾^!�Ƥ�F�#,�9��ƢC��5Z�^��o�I$�I$cd�(&�ܽ�n�r���s �m����sU¨*[j�kٽ^v�qM��˴��߲!�Y��jji�d�a��<�l��Z��ݞw˾u��l�?8�drI`!%K�U���yԬ��>u�,r��#<�佈i�l�Y���1�Un��$��� �L�����>!F���kPdiY΢����,��欲���T�M�J�D� ��V�j��'.1��:��iY%!l���54�C0�w�����uʾ[�mR��J@�� �G|����T������)�B�5D4��}
�[�j�����^U˓��I$�I%6�5ݼ��wNu�ո� P���T � 
��]ժ�u���R�)p�<�+6�,��w�r�Vs��C�8�Ԙ�؄ae�ګ�E� 80��y��u��w�����U��膑��W�L־�V�\�U�]b�>R���I#`IE�-֪�ewg���Թ���}(�dm&t�<��jhi�C!���,�m�_@IȔ��:�X����;�/S5��ۖ��0�ڇ!�A��^oGW��o<[#�J��Gm�8Á�����/�q��Y�p�7Uy��^z!�!Ҳ�2���T��1~v��} �  N ���pIƫڪ�s�AU�i���{�0WU�Uo�6�l��ܶs�\c�xy/n�J���;��[�n���n�=ڤ        �   *�  � T��*�p
� M�     U� �T P   n-Ī"ۭTu��l�|@xv�xݪ��ٶ����m��@l;�[|�S� 6�֨~?H�#p��%\��|�o�ҋ�b����!�^*\�P��,�Nk�Y��μ���T� �F␒E$"FyG��!�C=���Z-�DC�Bqj�!�A��:ܻ$�`I* F#��j�� �B�ʢ�p����ƢC��l�dn�}u��u�\�����*�7 I)�z��3�SNK$3>#�M�X�b�v��Hqx�r�B�24��9����I"@M������^T�z�;�kU_ˮK؆�,d���^�kˁ�)���o���� ҡ����]�nΟ=��u� [!�+k�EQ�*���婬iB�ӀI$	��+�y֪�w�UC�8�Ԙ�X�ae��5`�j!ʶw�j�����v6��M�H� �P�U��D4�t��El���L�SNK$3>>/d���k�x�;n�!��7��(�"�IB�֪����yT�j�i�C:-4FyG��!�C�yު�z��obFB7$� ���->��v\+da^~�C��M�k�#,�?j���X�C�$�@)��V�W����"���UꭐѸFb�MM9,��0���m��E��_+����$�I%H��n�]ܾ<kN� P� <� w PP�ӱWw�ͧ�T�h��u�qx���+#:T�E�j�iA򵪽���V��)z��*� ԟ�Gz�y�>u�7�U���r�����5�24��Q�qq�1Q���5���(����$ZZ���5����Tح�,��O��臈�J�W�����%Z�r�T�o��)�	80���[�Z�oL�/��y��u�:�Z��t�4��5�܂�C���S\����M($�6�/�uj�b���2�5�8[���0��j�$W�!��oa⯗�o<E_+�I$��8�C�s�T�Cf�׹m�h ��
�J�;�lr�n���Vk5�}�F|{Ձ��Q"��l�`��^jaW�:V*���Ü���5��
t��x�I�-*����[}ޔ^��j��I�u��/&W���,�R69�Nu�W��ʧ�8 &��U򵪳�<��"^Om�22�5�8[�����q�ni�%�Özj��Rr*ũ$�!W�ʷ�#�إr�Z�e�y�qx�C�w<m�,�_Y�����z!�"����PJ�	(W��ޣ�6-�!�a���OX��X�#Ǥ��iV��>�>u.�W��.{��I$�I��|��Fm�wy���t/p U�UTUO�*��u�%r�/m��γk�^5�I[Ad8Y�K�,�Y�'�c"�3G��-�Y�������$m� ��+�*�V�o�*�i�y\j�"�0��Vkƈ�OL�k{̽�[*9�I$h�*�F���M�//ˢ8�ψ�sҋ�B߳�놼�ak�D6@�F�uF���G��G�'��B[��I��w}o�օ��I� W"�=��qeCxbp����wR[}nb�?������߯���� U� ' c �ersٞ������T����Nu��ӻ��^q{��q�V�r�k��/=�M����ڛظ�z�5��       �      p*�/R��B�+�m��� l   �PU  �  @ *�U6�
��������U_ <�{����7�v�����\� ���@�PU=8n�[�ڨ%_�.����{mm�I�b3VV��7�Q�w�t��J��G#`Hk��}�؏tO#���1�ι�ۘ�*R<��$��NN��ͧ;�n����7΢��uAR=.�I�����Ԍ#��߰�,�v��~+��Z�;a5l��Ƌ�NɅ�a�1��H

�j��I0$��
�W�;��/P�5x�r�c#K8T�E�r���&9Z�r����7���Sۤ�$JT�C]l�m{;k[@pw W��� 6�A�( ��7=���_-��ұ����8S��g,�J-P�5�2,}ni��g3_��^sx�R*��uX!Y��sV9Wde�g#uW�����x�sUA�Ul���Mg4�O�d�T�IgC�Y��3��\��u����!�^*��X��,�Ri�_#�yS7��(��RQ$�HGYFyu�{�!����d#-3^\�H�p�]�r���;�$�n�I9!
�^U����+�Zի1�X^5��g#uW��C=���~��ߟ�¨��������֣˻]� �b��E��=s���X��)
�H�RUQR�ww��l�C0��d�3V�#O	;VC�8�L�>�.�W��.��:<��I"@A*#�ƢB�+P�p�3�<��"^Om�22�5��ۖ��0�X�QD� I$	q_#εW��{�p�����=�j�9x�Cl��kU{���U�J`I#l�]�C�C�M*+�e�i��m���y&جf�G�	;VC�8�VD%Q�p"�I ��u���y>�*��CQ!c��d8Y��%�CH�2}�|�y�>w[{�T�I$���1@ǯ:�<�{=�� C�{eP��z���;_7����+���w�;��(��9j�+��P�t��eU�FY�sV�D8�z
@�V�ۦL굪��f�^������ѶFbf��rY?BΑ�M�X�b�O�M�EI$�@ i��U��N��X���w(X�(i���
܇��<�������bѦ�q �	��Z�E�f��r���,�梇!�A���C�sK�s��5�ERQ&�$��Gu��F��G{�����^r��z!��6*6��L�SNK'�-^U�����I$t�"P�H�~�i�o;����^� ��
� �U`�ލĀ�  80���[�_���3Ds^*��X���&cܡ����z�_+Z�|���6ҩ�� I�ha�Ƹ��X��Lא�nZ?Ye���P�5�3�u�p�k�HQZ(꺠�@r�.�~��ɽ�u��F��[;��F��u��C��3 �������t�)�5�m�%K��^U���E�A��I�XΑ�x���b�3�8T�D���5ו^�w�	$  M�J�8Y�K؆�O	������m���j����|�:��*�*���:��z}��m���ì��S-��    �x��1�     c ���<��p0    '    N p0 �   c <m� P
�U�J�TZ�om��]ԷM�ۻ+(*�mu���n��m)����q�ݵM���z���� �aWD*���P ��w �[��*��v���:����|�6kk�p0W�]C�A8 :�ⷔ< s᛫�N�{:��a����� 
������J�;���7{ȩ\�U��f�YZɕs�
����8�گG{�U���wR���j�Mݱ�����ީ����w-�����ol*�jb֭uݬm����x��v�y�z�&@m��{�2wwn��9Zê��o�y��w�lv���X���m���w�x����Sa�ݹ�;M=���ݾ6�o�融Νֶ�f��޽ލ�                                   m� T�Te;�          �     P    �       �     < @   *�  
�  �  n�6@� ��ص�   
�    w   �@     *l�    �  a�       
�           
�*�  P  �  
� �   �   d P          T�     =�    �  �  �  �    J� U x   ��
���kKm�q���� m݂��+(-3B� 6��Υ:�U�S����ׯ�8   < < � �v�lL�֛[T^��^�[��Sb�Ur��㸼�<�n���)i[�un��u�Umۻ�u�W�rr��]V�      Y]�   x  p  <c�UQ� U F�   x @
� T P
�UP-�ʥS�zm�<𮯛� ��W�����f���]@JTUU *�*��m�V=��n����rI$D�u��ʳ^#�P�r��VM�;μi��;��p�7y��3���N�D�D�I$���]�Gϧ�agH�=�+!�L��Ob�t�k�T��E����1�t������(
�s^4֐��Ր�dg�y/b�D3|�w�����M�?E�U}��0��I#lICq�|�=_��9��Y��eU��,�5`�i�!��p�7U_6��Rq"@��$�6B��*���b�p��������0��I�+�MW�+�<�����\�$���:"������l�ݷ�= ��
�UwJ��
�W��x��Ub=<���4پb�;���������t�y��6G 	�k�|�]���깖�}���ߞ�bə�ͷ��<���)	$���IL�cߊ��U��b�1�����ɻr�r�|ڥO5� F�
a�o��=(�E���c�S:�������ͱ�4� IE"E՞�0p�,C�B�mC�֯��~�U|��z�Wy��X�[���$�ILCAQ`+)�B��U$B���l;��� ��W�t�������Ƣ���|p���S�g��*�MUv����r��/�f�X�+�D0B�	(��[����~�|��y���gҥ�Z�i��+�z�uJf��z�ͪ�����u $�ि��r�m.���/U�!�ܿ����[P�5�=���_/*�x��}�����6�dtp<t�9��Ƣ��|p���S
��⒮^N���*�׷��G�@����1w���p�7~��s[�YC�)��|��f���u��I$�ICr�lV���M=�w^�w`
�b���Tw
����l�������N�c��s�=��5���jd���;��ɽ?J�I��*�yV��PL��~��=�j����x�8uW����*��_*��e룢����A�@�/y�1ߕ�J�r�����g-G�I�u����������.����*�A$� 7��y��u���5�!���(�^�0�a�5M8��Mo��&��tj�V�r�-�]*)I��B	����u���o�|��9�;�ѱ:C=�y`qx�C���XG��T�7��x���+��۽w��[:�o��W0 *�qSn��ʠ*��m�t�H$��$B��u�T�p�j��ƹM8��gH�olVq�C�(9޾^U����ui��@��$�1�$��ar}C�����
Ղ�8������Te-���S����~�?9�H� ��ˍW*����G�b�'��+!�K�A2��#����GX����T��	 `;��U�>�҆z!�!�Q\#-q�SN;$2�2��x�u��[�x�!$�@�U]�(��L)��anC�����
Ղ�z�m޴4�G��Q���5W�� k�1�p��� �۝��-�.�nm�V�]N����ڴ4�h�֢�w���o7�l,��n�fx�ko��wO+��ާgi���w[��m��=z�l��0      PN T
��  �  �Twx@�*T �   ^�*�@�  � �   *�� 6��[nbwm�}����Hu�]Q�X��[�;v��{r 6ø�� ��S��{yڒ�_7�������uy�!�E�f�#J�ꕟr����	\��b��c��Q@��%������b���g��*���2*6��\k�ӎ��t�|����n�Cںx�U��ݞ�ZC�J�%z�`�7��.*<�5�+�t������ERl�����V�bƩ�4��Ƽ��!�E��y�/$�w��ʷ�+�tߚ� $����Uj��-�]o?�αU΢��������3"�p��ƹ^�����n�v_6�<uwx�������{�W�*d�.���z�' %%\���t�����|������ҩ�^�X8��4ɄP桨�5{��@I$�@ܔGu*�{���^ҼC"��Y�/W�[���C�k�N�-�Y����VR��r/��o<Gu�J�V���Gu��5�*i���^�%g�"n�ݓIJI IB�Uv����ؕj�t����`V�����܇Hq�Sl+��yU���qJ(D�������>u�7���S��[&:�X��WYj�W����]��U˕7��$�IP��ڛg�]������UJ�M1VP�T�HWy;mڨWVs��}%J0:��;����'���eۚ���$�#rI 62����=JU��c���re�5ݾ�e�Nt,`B9$�6�rJE2J}��.�٫[W�V�}tW���ƅ���g<�ן^*ނr2 �E�j�\||B輡��F:TC!�AA.�ƪ��^����ξU�<�<��F����^X�����_���\���|;�^ �L2Y!�a�$��ZF��~~~�������n�v�ۀl;��_2�����[wa�lnI ��/*�t���]b��g�[��4A����X�#<�yXеZ�K����a HR�Gx�jW��Z"0�kj�0�Σ��j��>��+Ug��{ʗ�(�7 �>u�:��,U~g���!�!Ҧ�F��.S�Hf|G1,T��� I )�B��X�����Y���Sl,F�:TP�h2�<��Z�W��گu(ۂ���!�cD��d^��xD�DC�B���]:�X���9o:��\�I$�l|��m����-���֜�@+(m���@�
��ֳٳ{�]�j�%Jp.�U�_.��;��O�|�u��ǈ�U�Vz!�!Ҝ�p��+�uG1 ` 2�\��|�j����4�9�Y. S�b�24��8h��O]j�bk7�)��H��ul��3ɼU�!�x`~Ռ�����D8a�.�T8!�a�n�B�Y�H�`�U���N���Uk.���8��x��k�#5T�:���5��6�$��/�]�~}jK$3>!�b�+C�����d4C���}�N�yb��J&�\|$�I     � �[Y.x�m]j%u *���*�WO���]������ZwN[U��<��f�6纖�W��:����z��9        ` *�  ;����܍�P �R� �  +(P�l  U   �P 
�z��T���<�A�[��uM��'��.�u C��Pw
�pU
����^�2���ګ� ����
��p�3ɼU�!�x`~Ռ����D8a�:�*X��99	8Et��*���8��8�K����ǌ�5`q�0�˖*���{J@���*���<D:VHh�#1�a����y&�N:�^_Woy�/*�t�>(\�@��$�4�)�b�,^O9QY��҅N6kV����*Ɔ�5�C�,d^�~n�|�A$��	%�rF���^!F����#
�J�2!��]U�Uk.��;��O�|��U���I#��q��U��;���t�� m�p{(S�5Ҡ	�k��g���*�����5:����7�=0����w\�����g��N���% ��
�S��aN��c��M���js'�#ڽuj�j���z� ?1Uk�-C�9h�p�]�p,C�§:�d8C�!���<x�&*(n�h�$ F��ռ��h�C�n��S�=��Sb�p��2�T����\�U3Rn�� @���]+\F�欇Hq�)�qx�]+5�ת��G�굊������I o-ui���m�Η��nPY[b��P�N�
���sa�w��i����E�C��	�XȽAj�b0�kj�{�J���H��@I ��8�z��/�^������D�^0���)מ��C�A����.]��dPrI$�&U�/._*������q|#��() �4n�H��r��,^O��Y���U3|Q���  M�Dw��*����ڭZ����XȽAj�b�B�mC�b�0��bk��1��$�)!_+U���
J��x�� ��0׌<F�ϲ_��U�˯��%I$��6R�"N��;۲�����dl����U@ PQ��*Q��� Rq��Uۥ�dPXf|C&�`�\~���Ր��I�>��u���yqt���H~#c��P�u��_*&�w��*����Ր�=�Cӌ�����D8a�u9�`6�G$`�q];u��\���Ca�A)*"<d٧�(��:��劽���Ų�PܒI%1+��D<D:Tب�#1�a����y&ج
��z��s�Y^�Xa#�@p�B�I�wX����U����m{2{k#����u�[�՟vt�H5��U9�[k���n�k�>-������P��� \�V^Y꩜��q�y����JfZ�8⳼�W4�gft޷���6Z�?ʤd�6��F�����+ծzi�);���p�<�L�#3����XE$7Hs7�p*m)���!̶շ[A�^��|���'JG I"N�[v�>�ގd���	��>�R��*�K(Ν���� $�)�{˻���~���wyw|E�w-��W��$�$�H c �  <U 2��m[��f�յr��v�Wp\�^�hyTm�D�uU{�C�Pۻx<n�nά�	gzZm���J�˫ն�/R��m�k����`        m� *�^�  ;�  ;�p�TGp  ���  mP ��*� @ *�U*��T<�r�fԾU�o��@'�̫�W��׮巷m��� �ح��T
����w�r��%A �@�=�oz��e>���g�o���f֞6d��T��� ����	��f��*d����a�J�"�/��:T9 �A�]�7��>��w}:�ݛ�u���[Ϟ�|�&�� @ �;��T������*�t�����Z�?'����Z�U9����JCcrI$P�B�Z�W���5P�V���|CO��R"0�5�G���%[��w��6{k�ݧ{��T;��� � *�S6�;��MF�#Q��!W�ʻ�:�QX��,3ՂD6 ����a�7UNS�!DV��t�T���$�H+�Wn���Q!�
�D��X,�#O��u��:[����*�,^]���(6�$��UR_b.!�
�����&�S"�e�v���i�DC�D�QR� �����8��V*��4�W�Б%C����j�"�Wx�ʯ�齉ҔȂI`�2K��C�t��x�,ID�a�2M�X,�U��oz�U��:���rI#Щ��ԯU��j(f��4 6ø�)Tp[hT��v��m�7{�hdigJl��d2s��|��okCe�z=��i�օJDUٻ�F�nS-Oܭr�S�~9]Z�Ui���Y�"CHP�!��M�pH�#UH�ҷ�$�@M��k{��}��D8T���C36�$�F�0�&I�E�U���ɠS�PI$��$�ʻ����l)�������̆B6���Qb�y��f���}��MS�A� �DW��μ�����r�˕<kT80�#
�J�2"D�(q������p;���Vl�Fݻ�ׯr���ku�U]�F�UPW���i���G�	 �r����{��U�GY���5l����#�-j�ܿp? 8S	��^_Woy�:Ch2�`�4��Q�A��j��*���y����� �(��NA&�d^�<#��g,��mC�q�����z��u��M;�  ���#R��!�<E�5����ܷ�j�mU}�K�|O�\��U߆�P`GL��W���m�zQuX������M��.���,�D,6��;sn�]�N6�PD��S���iQ��x G�U��� w6�VSm�\�ЪU&�c����W�����b���;�T������V�j���r��-��&�ʘ�BI#�!W������r�b���u�����yW��׹.����Qn�(��( ���D�P����-U��f��~��|��t��.���Y񢹵I.�B�1��)'��_��8�._*���x��V�����O?�.�����Uu���$RI$7%8����㊺�n��=��v���z+�]�b[�h =$�I��W�	��8B��]6�U�[`���8w�6˷a8mͻZ^u_ 5��w���nۇ���f�w\����n�����{�w)����Y     
� U� P <  p *�w
qP �M� `  P  l  U T   C�y�*'u�ۦc��]vT��6���-�� pw W̠ � �P�͵^���T�$�n�$�����ٽr������v��0$�H� �8�:x]����b�u�y�&6����
S����J�ꪡ�y}}���=S�*Pq���{����Ur�䐈�������`��6���}�%}��y:]a*I7$�0��b���iu��*��Z��y�V��V��w��賷��U��M� 붕�n^���69����_�ª׺�cU;��*����ww���#R����Uz�;�U�������,�ҥg� �hx�||o�DD�r %�*�T�kW�Y����V(�f����*�����[%�($ �I a%]Wʼ��{��~ū��wc�i�pX�サc8~�^�R%� �#��b���;�/�K���8���qb����J�1�������ȣ�@ 
�y|�[}޺�Uj�r�����}�Y��%I$�H�C�+�&����[���̠ ��U���p V��Uwq^�]U*�^���}�����H���8��6���4��L�.�Ub�1ӭ�4�|ܒI#RQ�������A&���:K�#�?>���Eݭ�V��I��#���0J"��&��qE8kL?as�}/�yV�X_qR
$�c�$�p���,7D�,�������g�Z����ʼ�^Zo})�%DA$� PIZ��dx������dY��]�w�U���V�-_����$�B��{woc�m��)x l;�+�( ;��* ym[ܽ��zTº�R�x0��H�!���.C�C������*�^To#˗�^��'I�I$��S���*�i����嵺%_-X�d�T�U�.��B�o��:��l�I*l������yV��O�Q�x��ݼLUb�׫�����h���I#m�$�t\�b���g]Z��Zo�J�5CHqx�{&��B4���V�U ���S���v�t���9*�Dx��4���#K\� �l���'����[ծ��v�b 6øUUUT�ܬ��-�����^��H� �IN��T�������yb�F��q
H+Vq�*9W�Yx���q@z@  ��%�j��Wgu���?7�`�8�*s�C �2(iyWٱ���`$ @K��X��\�i�Z{O��\�|��u��.�� �62B��_v��7�[��{�����}�G�=�w ~H.PI@ �!�N��&�hS��!� Nk*`��	q�]V*���Eu�5���Jߏ��RV<`us��  < �   <   �     1i������1�     �p ' c  < < w06� ��U����w�.��][�=Vel��O�Sk����8^�1�{����vݦ�r;�zZ�!^���WvݷԀ�T��^�^���N,Y&�e�����f��Z��   '*�`��uQW����.O8�(󶶃mwt�g�. �s76��u�X�@��*�� ��������.���wcb�
��ot')�޵ݶ�Fm����j��{��)��z뺲����d�u�kp꼮�M���w]���T;��s�j-]�l�`���Y�����zb�׮�z�f�mOWJ��j�X�u��ov�M�ػ������n��sܣ�u��qn���r�r[�f�ݱ����^�ym���Wo.��u�                            �       �B��*��       � @       P:�                 �T � AT P\�
��U*���ԻoX   V�   � c  wP U  8@ƪ�@  N   P   �                ۲�  
� �  P �U    p            	�    *�     <       �   w@
��     �
�|��  ;� ��7k�֠ {�UR�*��  ����� ����`<[�g~o��{;�p0  ��	���p�e��z�on���5���W����iJ�W8���q.c�n�m��*(R��M*'�J8R�Jj�e�Ѳ��l       ��   ܀ � x Ë`� `*�� 6� <   � ` � 0� PwT�o6�J��μ�����;�M��^m�����z�w2 �C�������UQf+wz�l�qfU�w�����̏��̢��4��k�x�+Z{X��8�y�NUj���$:��I�;J�aGr�B8�>�X0�"p.b��yb�����U��Wt�H���� M�Dw��D�wY1TU�]wz�P���ǳ(�:F�m)��4�Ω��I1�$�F��;��,�E|�Wʶf۰��4��k�x��4�Y�4�8y���2I 2ʢ�.��*�r�H��B�#���Ճ�'�,F�#����� �mv��J�i�˧|�ogm��wm�P wyTk�AK�P���T�c���8*��X��O��:�C���ʾ"���`�q4G�{2�:�U�U��)��H	$m�I)���0�t�Cu���<C>?;����Y�c���"P��Jhr�U�
J�E�	(��
<GT�,B8�/����V*������6�!N��X8�<Ar
68�#�RAZ���,��&*��b뭹��R��o��#r@.Qr�U�ʭWv�uj�U��q���q�<C>!�<XF�@ArX'��i���o��{:� �ª�U]YQ۰ UT�[lw�{4���&��Ui�>�z�ʱZ}�HE��C(���:ܡb�iq�
��l���0���$�����u�����X����V��8�,I����Ŋw[������ m�^*���̢8�D�L��0�t5#ʖV�Wʵ|��m'�Ӹ `���+���0�i�f�<G*OT�B����J�\�}��7�B��Fې��n�W����wV�vR޶�qx�Q�C�<��RAZ���,Է� �d�ܛ�w����%�w�� ��U���*�*����m�����lA'���V�.�\�QR��[��a�0�ژ1!�a^�R�#�y4�MJr(� F�֪���o[��Ki�׈�V���Z#����A�}��ܩ � B���W�|�gx�"C���Ճ��s��i�IUR�R�X���U��S�I"�Dw��j��Y3έV,]~�������ث�Z�����b�]��Kʝ0$�m�(Buj�UV�+�Z�V��w_*��ʞj>U�O�/o���X�����I$�Nnwj��*�^y�n�Z�����J�pJ��wuձ�Kmk�I�����W��U��U����J��i��j��x����`�4�I�|��$�� uu����Q��y�*�u�I�oP�ff��A�4>הG#g[mw�� G#� �R�GX���J�0aA�Q�������rCM5*�U���=����$m�B�d��<G*M��Q�B<aG��:�^_Woy�Z�U�θ�ZPܒI" �Z88�<A�D,x�Hq$�E�&U���q�7r�� ڐ=�BQ '        '^����ݛ�*�v�8�N+���5[�]�N�Sl�Z=��n�m�x�m;��m�Of�u%��^��Ǿ�ns�i��m�v�8�ݨ       �`   <  ��
� �[ �
��  Tm�  +�� *�TPATP *��T<d�[e^���� NU9�۵{z���۹v;C7k ��U�
�l A^��b��I$��|S%ث��Z���/���0��TX,��2�x�x�m���n���.t��H	�0W�,Ui�y2y�Jsj�G%J�q�8�_qR�:�^�&��)I)$�@	!J����.XS�����]�&���#����.��n�$����^�����F��`�8���Ff��T��F�6wX�c�+W�Ց�0�=�5��8�Rz�DrPt9V(�}oI%I$�H�(����kr�;�{{�� ��uol���l
Ɇ44/�  p�B�[�U��v��#����#OzJ�c�rC��%w��T]���~	� ��C��f��A���הG#��J:�V���uj�Wf�nq F�8Ԃ��V�WM�wX��*y��Wʭ?,����ʱy>�'*��3�y�TT�@�$T;��E^U�7�\�b�/���80,F�4WIT,q��dۍ82I$� 5%�*�Qwu�<����n��E�����0��4��T�m{��}������ 1{h"�/^�wy��ooP ��
�e�R��m�'P�lnI$��A�U��ᢱ�a�����Hx��׈������]|�W���T�A�AI wʳZ��P�l�G[���4�G5`�Y��R޶��W�*F���@��d
���h���;�X�|���ֆ�Qy�|Eb���(�t�#ݾ(�P��F�l)�EuX��}D0a�&�U�#�w�4C�h�Wʮ�K{FA�HۊHm2���(����J�Cd2:ܠ��u������_k�u�t$�I$�I��.���i��I�uk�� m�p��UPU`T�����06�J�ƪ���i�H��!c�Ш�!c��n������؆/7&2/PZ�4�TrPܐ�.�\��yS���~�X��tR��: ��F��֏��m��ï5$��	�|�b��\Թ�4�aS
��h.Pt��6b�[}e9O�b�.�n�3�q����uk!�@�f�88�<t�r����(�![��g<R<��W�"m�_&~Q�  ܗ���|���c�D:|p��L8�b�+9��!�<Gu��UkV���I$�I$ ��;�/f�J�v���@P���������TE����ٽ��*��7�ߟ����u������j�y�.����_*����
����1�gf�ҍ4�N���de2IRI d)ޣεW�+�<o?��]������+��,tZe��r�g5;�U�}@pJ �_��ʹb���B/S>�8[��"0�
MP�9h25<����yVsŽv�D�R6�����agǱ�X^5�*i�0�7Ux�A������(\#-3Mg4�@� �@P�_��ʳ��sε~���,gH�T{B����]%c����y���~U�` �6� �  p���=z���3��U*芺g6��
m׻#mۊ�ql�ww;�nwp��S�ck���Ev��O�V/s�m��*a�.�S       
��  T  �  �6�mjPU�*�� l P6����� � T P *TP�*���T�/U��o0 ��;v�{u�����]�n ��wz��p�ȩ�b��oq���T�������>�����^_�d���S�W��Tߺ��֫T�y�E���f�*I%t�� ��V�5�:p�r��VM�;���5�"��Y�����x��cH���I �¯U\z��V���j��(+�QG9�k���
7�̥UV���$� ~ͷ������=ݷU�6G�rV5�fߦV<�XH�b�r8
��ݩ�G>��>8]۸o[���ý��:���"�I$�$ےTE���M���v��ª�UATm�UUY�ww�޾�j�t{�����&ʡ.�r�H��.�r��u����\R����RI$�R�k�վ]�*əRE�
�.fl�j�f�l�.��O��NHܒHS%���,�\����1QKs�;���s����ыR�&� ͻs�W���+�l�����ӗl�)��߳O��G*H$��UUv��ژ枅n�^�RZ��|x��ﻭ���v�+� �I���kok��u÷Wxڽ�7������U=fATUn5�v�eP�Ug^ؗ�o���6i�1[{��T�1�(�;�t���**B@ �G��Ӫi��Űl��r(��i��$�+�p%N�#p
{f��]�o�;���}�wZ�ߪM�'���3�u+]j�{�yޫZ��}��6�d���I$��]��CH���w&2/S5�����"0�
=P�9h24�l�Y�q���H  jA]r�Z�Y{�w[��Q"���#uK�NC�C�9���Rޭ��'�|E$�I*7$��nR��WvN� �w W�T��*
�40*�H(9$�GP���/�hɔ���<$�Y��x���������J�~]r���J���$�� Ԅuz�j���{����*��g[#-3^\M�L�!����C״��/�W�b���n7$�I�:�V�y�6J6!Yg��X^*�"��#u.���������w���Pd�� C!i���B!�!��
��A���NՐ�/��а24��_ ��U@��@�(A���s�T�x�Յ��Pl�o�B!����E�gָ�u��yr�[]�$�I$�D�k��u�}�&%.V��pw
��UQ� 
����a���m���Y߯ﯨB4�r�2!�Ƥ�V!Yg��YY����*����U{ϧ�zSAؤ�Ӓ��u�^N��S�]�[V�B!�#�ey���:$�Y���޿��#d�6�!N�#WZ��W��D,tVe��r�fj�o,ٴ���*������O=G̴�y$I7wuK)Vf"!���3��#J�u�p��q�1U�Fx�9�E�Q5�>��	$�@dr!��媽�g��=��*���e�i�T"0���s�U�[M��rI!�I�8@p  P�8G{���'L��S1�;��=Q8����N<��ݕfu�޹�Um��3�]�n���u��vlJ���V-�[���0      QV� @ �  �T��lt�m�lUP � @ol�����  �  
�  *��
՞�0���"�v  �[{R��ib��m��]� �+����[*���*�e�ݖ��G6�L#����'Կ��;�U���p�hB+ ���kK#yM�ҽhB!�6��y�IU I$��R�p�C��؈�L8B�f�F���(g/*�x��	\�֭S���>�H �UV�8�j!�T�\adn��=��SeP�Fbeځ�B!�!�r����Q P @)�w��U�������qx�������)Ȩ���Q~w�y�굪��y���Jdm����x�x�Ҳd#u3^\M�L�!���i�!�A��s�J����f���n��;m��n7��{^��K�� ��
�+(�[j���[�]�3��H\�֯�޾.��G:�Gy�dn��3��#H�
�*��37�A����`B�v�TZ�U��S�4G���n��#��L�Y�$�T��hU���������I����,��^��!�VT�F�f�OfQ�gHNj�!�o���@�T���NHB���f�Gu��TZ�e�j��x���<5�����[�4�t�x)�M�crI$���U��.��!�,�8c�Wƈ�4��m�3Ds^)��WZ��S�����)!%I#���]U:����w{�.��@�w
���� J���V���ʭ�{{�eDx��
Ռ�dg�4ޑgL`�Ld^�h�4�eΖt��HJ-��$#@��B�Ui�ӝ_+U��ӹW�Yg��X:yW���ٚߨ*^�H$�� I+��5뭆=��n��n�r�����5Ⰶ�AT��ܒI#T�*�Uyh��+9�&B�+P�p�3�l�V��"/IܙO=G�7���t29$����ت0���r��۪���Y�9q�}D��֭Y{�wY������o�BHUUz���{�]瞫uv���q ���UZ�UO+(*�e�;�owʻ��Ug��U�z����iT�(\#-3MA2�ن�L�|e����~���S
��6�n���yVs�=��y��,�Q�"�E�Z���+P�p�3�^�k>y�4������$���5/!i��-�e�t��r�W?T���.5&*�A8Yf㚨�4�H�$	�wY��s�Tw���#vU�A�����V�����r�<���[�U3[���m� pd)ޯGZG�;k�����didr�c�~F��N��:�U���7���I$����]����nk�c�[�� *�p�ʥW�@ASλ�j����=UD��?v��W,W��MU��g�b�:F�t�CYTUs��#�� ��� 5%\�֪ɽn��O��!=5�q���c!�ҮJW]�[��:T0p$�IB�W(�ʼ-�WƢg�v�G5�p.hX�R�ܪVs�c�����C��	�(��V��>����*Ջm/\�E�;hx_y���#�i�!�L��FQ��F����$�DwV�5���)Z��*�fۺ�#^/���]�׆��]|�����~~���[��` m�` �
�Nm�e���.���xwVU��*�Uw{���׷n��\lM����tӶs�4�*6mݒ�z����׺��7[����Zٳ       U�   �  p�sۀ �;�[ x
�l   <*�T���*��  *��T�P+�UQ��p��_��x��^۳�ױ����q� a�U�@
�p *�^Z������U�_�����|����~�j���9�����ݞwV��C��[�S���-T�z.�$m�J	 ₫���X���<�Uj����}>^?3�;�Ȭ\kP��Y�:F�����$�  �Q_"�j�'y�:���_�ɢ���b��m������?�y��֪��O7�gⓄ�� �r�z/�Ҧʡp��˵ʄCfGd�
��A���NՐ�/3ƴ�UiI$���)�d�u���y>�J�v���c��c8Y���Գ�x�z��r�M|g%�$�I	%&`�cD��)�ֶ�f\�
��U[�5S�T-������8nHZ��g��Yֹr�kk��P��ꠇ�,���/�/��.C��7$��
B�V�W������GJsԅ�/4�*\�V�YNb9֪�w��]�%I�@H_!V��=��z�֪�������D!�C���)�z�=������"@)��E�G�#o�(�tä.�a�k���m��t���w[�V���T�m�~H �UkE�Q"���#uW��9�2U�f&i��ن�lۻ��ݫ�Z������ۖ��˺ 
��
�R�T;��*s2�n���z@���^��W�;�оB���L�#m3�Ԋ����B�,���S���-�*6�
a�;UZo��|Fb�Z����Q�=�Nx��E��^O7㊾^U��^�����P�l$b��V�|������s�~;��ő���z�C�C�9�B���k:J� IƤ�ܢ�򬾱�G:�<xIڲ!��3ڎF�g�w	����/���p���crI$RJ#�p�3�l���E��x�ӕ2�����ߢϡԡ����r�?iC�����q�w=��k��uwz�ܮ���wP�;�U|��� 
��]ڡ绻�heR$#��j��-���+�Zի/yA�i���SMC#uW��Y9���O�mA�7$�@aWʮ=_G�d"0�;&R�5dx���Y��N�}段W��.7���R2IP H`��C�X�X�FyM��Y膑gr�B2�>�����"0�X�K�6�$F�H9WȷZ����u�Hqq�1Q���=�-5�y�j�y�;�S?l�F���K臈�J�(��f&i��ن�sGZ����_!Vs�h�^�  ;���;����m����u� *���U�����J�-���7��SbI$���N�r��/��pT��h�\�サc#zl�u���gn��kW�z��9$��	$���g{��m��7|�}R��<��FLo���)=X#5%wTR�iZJ[�^3`ײisԄ�iι%�l�<}��h�4����I`B�v�4�30(��R$�$X�N��_o���>�z�>�@$��8N���~�Sf�0�����(Ls�;T{�MR��d�]�ڔ%�PI	� 7mt          �   8@  �{mTp��=��  �	���� �0  �k�  ��;v�1�p��G���USdr��f�m���g�ڹ��3r+w��[Y�Q��<�[�n���L����
�
�e�`��S�� �
�*�YE�;��;�N�xN�ٞ��NɌ�+� ��O�o���pu`=�j�|��'�#��\��J9\h��,-ݻ�u������š8{�������kaTR��@�U�J�m���ll�VNm���.� *��]��mM�c2�wwjM�t��V���66KgFu��d�u\(����^����ݺ���m���M�n�6b;5�WW{w=�k�S��	F�1����N��oo��v�;���;�.�Pۺݦֲ�R��;[{�n�][���y�QS/rw�յH�j���z�                                      *��� Uw          
�P ��    m��              *�       N-�@  UT U� �U��[��`   @   �   p  @  <-�T       
���P         � @� �kj
� [F *^���� Y@*�� EP  w          
� � �        ]�    
� @  [  m���    
��T  *�@++l 6ʟ~��|}� m�)ݵR�m� PO-�����nf���{�ݽ�	c �  < �  od��,�\[1��'���g����zeon���i:N�u���u\�K[�m���yǵou�z��Y�d��S��j{����       *��   x  ��� ���
��;�VS `  P  o�~�Ee@ U*�U C�UN 6�{9ˑ' <ƹ����Q�{��ԭK �w W�T � UGuv�~���@�����/�|�+,��^3�g�")�R�L�Q�C�Q�4�{�]��%-H�#�%�sǄ��!�C��0g�digJnU���ʝ�uz�j�����1~_�� J�?*�j��|����yS~�!����CX�Vs��C�8���t���� 8�ʭj�e�)]�k�uO�#uW��Y�D:T�ENUv��x&@ �8K�Qq�&R�2�#Ǆ��!�:/�^�8�yj�}ϝJ�q�V����I"�!�I��u��EK��͛�ր��U�(
��l�r�f�j�k�U�g#<��<��a��;�1����!�ߢ��t��L9bdiQ����i6��I������x��b���2�y�c��Qx���p�dn��'/R�^S{��$�I$ N_*�zk�<�!�!��W�Zdx�d:Gk�����Y��{�U5)X�������Xj.!c��c8Y��哖�3�Si���m�,�H�� �B�#�H��
+�sϕ|��u��t��I���0��c�ËME�Y;�9Z�^�>ߺI$�I"JIf�ܻd�;��ݞ� U�Uk�lU<AR�z���K��ڧNS������C�d���34�y,CfCɔ��U|�����yV��i<5߈�I`J)S�U�˻��J�v�'ʝ�
Ռ�dg��=u��H����S!i����J�� #r@
�\�u�˗�<�a�k#J��2>��f���p�-b��R�����U��N�� �I$m���Tr,��\���E�!ұ�"���eKr�4a�<�J��L����D��G �;��[����}�w����R(������Z��,��d�Ϲڮ_+��zJ�I$��r0@�7���Ǫ��2�� ����2�� Ae�uU�����d���}o�W��o�`�L:B�a�e�F���!�ڬ��D�V�j���|� �UGE�Z���Å����z��D:U�D\#12�G��6a�[p�R��M� �;�yꯖwg�|�[�`�hX��Ε�,8��P��
�z�j���s�������v�����Si��-�,�HS6��P������Z����b�!�r�	r1
�TZ�Y{�V�����Y;������^"*j�.��I�>�~w���;u�婃{kv��8+����{( ;�1�`,�R�� 	$���._*���s�_,�;VC�8�S{B�F�t��a�f�ӌ�9����-UUT	9)�0�|�������L�e�h�4�,���Omj��x�S�ФבI��5 �z�Vk�w[&���V^����z��g���y���£�����DlnI$���W��=B�+TZ�Vc�WƏ���j�t�k�0g�c#K8���t���J�  ����h_*�V�3���R��sƈggr�B2֡bF��֯-^U}����HE$��b � ��w
����9g����NTw��{c�nv����xUJgZ��i��R��
�w�v��۷���]^��u��ݳ��       ]�     �  T:kCl `*�� 6�  @ �� ���U  �  U�<Sr�ͰU�6�K�^�c*[e��q]w�m�%w6n�j *�ت��TUռ��r��M��{�޽�6!�L_!b�O{��W�ʳ]�]�r��W�yJ�����}%�p	�@a � �E%z�xVC�kvl�T�#��+��4�7��}�9��y��p�I$�5J�yT[�éY��Dpz��a�/TO,�����\x��{�d�6���[��L�	�f���U��X��q�1U�1V/�r���!yS��K4n �F�8,x��^.A�:C �uB��Ƌv�j�Z�&���_*򕛾�I$�Tn%թU�m޵]��O� �w /UY@� *�ηH���P��+�e�iL��i����"�E��"c��`��^�$�Y�d2%������lp�F	�^*��R7��V�T�o��_�5���w\#��k�}D�`$����~B�7�~��Wl��ڿ��j�n����!n͕��j��~\	��@0���,]��=�Α�iL��id�!c��-U��*��*�}�|&�A�	$�
a!+U��UïU\f8����u����Qc�#�k��}o%{���I)�Km*�jj�kw:ֹ�z� ���� ;�l mmf���UfiF����o���<�E�}�Ε/*�H�MUv�B�u�U�$�H�.������Ə���߷�9�*�S�/yT[�éY�еTͰT� F��!WV�T������ʵW]+�z�O}1E���V�T�-S�Ui�h5�R�6��$��U��x��g*��z�r���!yW�yJ��Wl��8��yV���?ͪc�P `A�򫷈]ЬU�}2�<��׳=��5Y���O�o}���w��??  �[�V����rZ�wu�n 
��*�tUF�l��ͮQ�r%S�i�9I ��9��+�g�^��Y��"3wS<FZ��7�u���t� ��(�$�� &͜f��_d���#��R_Q�����_��|�Ԩ����9�F��F@�H`�*�_�Rz���W��!X�*�e�y��Vg��yVk�޿����F��')�*�Z�ok�R���l�-��_*�{��B�_�5ڈO�A�	�u�j��� Z.]�/®صLB�}�4��_c�����V��W���_�T ��q�ݛz��w��nӽ췺 +�
��U]�T
����Uw�y�($��_�H�ǼU��b��E1U��d+�x�<���O�n�kn@�� $�J��i�O�U���[��{]�r����/�*<뻻�_��*�@��ԒH� ���?��"�W��r,S�/����{����5�;�?
�]�&�k 8~`�����c�R��{l��~�I抦*�~B̅b�X���o[j��P� �w��_k�x�#�ҝ�=c>�(��!c�a��qԭ_*�}��ɸRI$�I%I$T1�p�  	�<Smuog;�ګ��Q�rr��m�Aƫo{���=�֯f�J�{1^���-���ڛy�۽2k�W{;y�w��[nm�3�m@       � 
��  �  
���UQ�UA  S` P<*���
� �>�   *��ؽUl�s�­���ۺ��w=���z�m�x�jǶ a�_2�� 6�*m��J�&���u)?�O?��"�V*�<���_�k�V�u��1?�E8�� n"��E���+�~B���R��{t��~�I��S\~B�n�n�  5.�V�*ɶ9�/ֽ�헩�,��f���P�3hR��h_��:�6��F�:����n��Uڤ:�U���_J�X��kT�*��d�S*�*<�NW��p[�g�^[��+���e{<���$����W��7�5���ת�W�� *V�UU�ʨ���sn��wwZ�{[�ml���0�����6����=���j��o'�����$Ht�+��h_�u8�r�[������Uv���~B���V*��_��N�( �GS��{R��������Ӂ�c�n�(�Wo<�����^��Z�T�{���^U���*��~B̙+b��s�^[ȭ������9�WO�H�lnI$��9%_ʼ�,����v��˽���r�[�z�Z��\:�A�����I$�IS���z�+�7-���뛞��ws�U ;��:�U]�[A������֪��h�J�֌�Z߷�ڞd��m�E%_f��%$m�.��H�1�J���j���S���&J�X�|d��W�n�
�nI#l2K�,���did���E��"�}C��B3�,V��tn]g�Ȗ�<
����'	��B���Z~.�7Ǝ��_:k���.%L�#�f�m7^��4 �)!%�s��a�R��#Ͼy������#_~��.���V����BI$�!�"�� �����rv;=� l;�+�P�F��s���H NH_�_*�wwޗ��kJvT��kC
rUX��dL�b���o{𪂒B% ��_��dG��g�K�YTɁ����f����'3O������7�?�  q�*�����q�+�#��س��{�Α��Z�f��~����j��	$�Eux��!ۛu�����M�gHmw�<2��LI�HX�Pd_I�/⬰#p����j������*��bܩ������02�Yf��qj���� �ϖ�Uz�r��/i�2 *�ت�Z U¨*[oU�n�nt�*CcrI$A^�*�~�;�ʅL��`qg����Ş#1W��3X,�U�oJ�5Q��@	Wʮ��*Xd2�v��dh28��w�]�W��%�*���zRi�����#DTpt[�x�5z��Y��=b�Y��ïUz=�\���U��q��	�R2I 6���Z������yV��9܎T*�ꛜ����>5��
)8HI��I��4U�f-y����÷76���߽O<ݠ�R$�I$�H���    Ԁ��vw{����j����媯r�{C�n�h�l��1�w�V�q�:����6���6�*�nBB3�Ep�T��U
м9�M��4      P�   >  ]�  �9۱
��;�V�  �     -��T *���*�@  n  ��͗i^�n�ͻ�ݗn�i�Ξ�b� G�Qz��� *��m��r���� B�L��?���u��~�ū���+��z���+<p�Ȍ���t�&Օ����@�� -��ʹZ��k�温��<�����
�CGE��-g?|����6:mHI$m�@+��U�>�G���j��ESUKy�#6����j��ޅ���~�w��V�' F�
a/W�f���V�
�_��.��T��uYg�b!d^�$���?29�����I��%꫏u��ɟ2����j�?iV�ynäs^jv&r�Z�L�$�ILBT�$JT��TǺ���� m�pwe�;�l{�6m��[V_57�~�7�ދ���TX��=�<�_���n���Uq�8��s�b�[��biQI�I$�����UV�z����k�gZd������!c�n�<~{+�/T�"*� F�80���Z�]�qש��u��W�`��N����TY�\vF�_��UPI$n"���V�3�_s�_/�w�E���t��y~�3ESU__�W���	$��i�=��9�f��q���r�#ܵK*z�z���y�������￀c�ʟ6�+om�ov�v��� *�qUWt �x*��U��.WJcn7%I$Pc�_ww������7YE�_��<�|�P�U�
�I&2H�aH���Z���;�9~�^�;����B�~Ξ�ʶ�e?j/�����&�.���$�A�*�Uv�\F����b��{о�{����O�Z�j�ǟ3�>�W��;{ҙBt�M�Rp:�՜���[V4�/S�z�`����νU#�q_5��X���n��:Q�#����渵U-�����}���T?tS�z,���T��<FZo9� /w�����ۜ�w�j��L��Pl�PxVP 
��a�]tI`J@W���Zf����y��s�<G��u��,��n^qD{�y��ҪA���$�F�rz�P�5�c�f�<~{+�/S�z�g���|u꫏u�� �^�2H� ���gÍ���sVY �����弭��_�W���u�;�����:�R8@���U�f=������������c�ͷ?V(a_n�B��Z����*~�m���&K��_cϙ֟d����g ���?=��Y��=b���_׿?��u���)�6=��oh�^��ƶ �wP�(�V�]�n�T�	P��@��'�U����4�}�!t�欲w+V@t�r�W!U�����)�J@�0���w����TX��>�<�_�ʫL�Vɘ<���ok��� �4'$;�wo�s�ڠ�=C�Nj;����ȳ�e$OO�N'  �J=;qN:���Oretp�Λ �����,� ���0 1�|���w�u�~��������|�F�����׮j��1��|ߐ�   U  Y@c�:�f���w��R�W{4�vU��6wVz������n��޴�5]��)wn��'ɶ���vo��h�\��k��[�v�      �� *� <  �UTQ��� n!Tx  �   k�@��  � �@ TAm��� ۼ�<�0|�2����͕�۔ U�Uk�Q�*��+���AS�`��_�VwB�\Z�E�ݼ�����T�1��mAcZ�*�����R^� � 41��T[������۫�.��Mo�D�q�8���1?8*M��$�)!�U��l�g�~�����x�)���t�Zn�|���7�J�Pd�� �A^��!l�c�����?G��7�
�T�3���i���n9H�r���Ъ�u9?yS���}�W��i>U�'�;���~?����=�w]���J��g@TxUw�P�@U,�TP�H�$�F�nSb���q�s�����Z�ߧ��u�{l_x�U�~�X�#���I��$	$�!H����<�LV���q�?P�U���_k��d��t�{���N�B��$�6� "'$����ԫ��8��ѵ?|���g}(��~�F��P|�w�J+ВH� �d*��>���V��^�e;��kY�d��o�#nI#m�#��ت���+�W�y������ݹ_�U���_c��h��� U�򪪻v^�/s���׹� �d�Ī�]m��V�7��#rH���{���֟t����Ԭ庬�~{���X����#�-(n�p�% !M�U��}M��~D�9�Y�]�Ճ�,�ʠ��^�t��p 80����[��U�}?b�:>�<�_ʼ��͢j����3n�|���bi~]?(B�	#�j�e�M�F�{U[	��F���|��M{���*�{�������@pa%�*��f�A�:���M_�*ﻟ-ﶞ�l���Jw��I$�&�m��7�s���a�� 6��*��N�
�6暌�okOQ�S��~~�n.����7�����Z��ܖ��6�	$���s���:�W�z����on��m��o���d�crI$PT��${u-����Gm�OH���7�*RT��$aH�����6�n�}���6z���+�p��J��h�M��$�9(��{�8�37z�ۻ�w&,�y�O�����zJ�I$���I��z�����v��YC��P� *����Vݷ�^�U�=��}�{����չح��ܩ�-��-n�_��Jc�r8$qf��o}>��8�E>������%;�nPU�]�U$��	%&�I��������Y��\;Mݾ���ϼ�_��H�$�v�wb:��<�+�����lV̘��s�Sg�5DA$��	'Jus3;H�r���c��Ks=\zSz1�.ߦ����?^���$P��T�~�q��zg�IX�q�%I�n74���1�\��1��jLD(ш�ZbB���$(݉
��d���Ql�)儔+�n[�ͮ�i��a%P�*(K����?N�yc���_���_����_<1��g��v��DP��<���BT���a��(c�����p�a��d�ͧ.s���"������4>��k��[v��������)ALB
�B�*�b�a)��,w3�d���UDP��^��_���w�b��v�Ç>��(d�:3�?������ׄ���˰���ݖ����"�μX8������7�Q"�eQ4��GvT�NL�F6���F����Z�h���O��~�8sc#a�Q1���Ϫ�������hi��)�Շ���βۊ�(c�N�.O�(d���r��ޮ6�a�c��Li�2��~��w��l���M���N[�����1��8pÊ��:�lm�ד���z%Hz�_f�-6�섩���S������e5����p	�}��/���}����S�           �Uϸ �K��CE��t4\��t�@���X�E��(�� �K����uUk�uZʸ�U*�jUX �-ԪU�2�YeR���U)s��T��B�5���R��ҥW�P��T� u��K���EV�ԥS�*w,�    `Ld0 �  ����@���M12d��a *���T��       "���I2�*       ��U&���      �D��!2a��5OMO)��@�"~��<��?m���� ����$�	��@$������� N7��1&�(�6 �%a�@�$��,�@�k���w���?E� � }�?�L��{>3��8�O���K����$h�+PP`,�$DDb�"E$PV,*D�F��X�X##X�Tb1QIUQmB��
��QE��1D����E`ȱETH���UQR*��*#JFжŀZ��)lDQ�c�X���)$P%�XE�Y1PH,J��`" ��Yj�d���cU�1��R�FVB���R�Qdb�(�AQb��U�FE )��`�Ȣ���Z�E����ER"��Ȱ �
ѐRB���Kc�PTPjV
�PbŊ��6U��K���"�U��"�E�EIQ$+Bڴ)#AdR,�ȬTYUJ�QAU�PY"²E�TV1E��R@Y��P��AE U $Rd*V$��+P*�)*(H�T�UB�
�
HE!X� �B�@�
�jIX�@�+	PZ1IR�I
�
ʑB,[hڂʒaR���++Z�R�bԬ
�P��+-�R��XT�Z$�Y-�@P*E��J"�(�%(�m
��F��)ڕ*ڤ�hT��-�*�dH�YR(�H�m$Y*�E-�RhJȢ"�D�� ŭ@PAQDdPY""�R���� *��T�)F�"�
�dE��~�[a��2POb !��i����������;?P�lP��d
�T 6�;m��  ���#�`mu��5�m��sT V��km�Keխ��I�+/��*�eͫqe�[�JdXd���S���ضwUEJ� @
�  �  6(T.aݺ�-���wM�  w*��ͪO��������d�����
� *��ةYB�ʭ�ye;��dc U
�    U � �  ;զ۹��v�[q���s�Y@�[�@ءT����n�QVٲ�YEP�
�P��n�l�UU 
�P �
� ��e�T    U
�-�+( V�    e �   �J�T  P
��J�����m�
�� *��   �
�� ��  �   
�     �
�    U*� *�   �ATUR� *        
��UsU�@ ��EPN`n*���  T��Yn��{cmP*��c-�VR�J��b��*��T)� 
l�TUn�5��\ʠ �� UU  �  VP �@ s
�� �[l��P `P�(���x� ��c`��@
�K��@6��@ ��}�T AM��      ��� �i�ק��m�ew:�%J�ywUܩ�Z� cJa]vc�5����Ln��Qӕ�kT�����Ͳ�6�9��ݨU�����Lj�if1�\&WW����-v�ę6��ʋ�u�mЮ[�V��K(,ʲ����R���5�5�A�]�i�����Qn�d0�75f�ҷj�v��J�[.�I���A�"�T-�6V��Fl�@T�M��͵4��m6ہ������]k͎܀  	R��@��l�U lP
�V�6�m���� �Vڨ��{�  �ՠ   ^n� ����������in5���+�-xM@��F�6��-�t��̫M���������I>v�	I>�<��! $������ �O�ܙ������@�-@ �Kh 0��������  ���T \���*�)^�*Y^�l��e[7zm�[g T �T T �� P@     @� �[��l�Ud��%EP�PX� =���.�TU  6)ܾlk���wQ�Zgm��u��]k��l����d�%��L��V�L\Uw]ú���U�m�5Yn��/�|=Iϟ�^��0h�nͰ��Sl�m`  [ ��UT9�v�Ҷ1u"��nNQf�����]�~1����Nm���g�|�unI��G9Ս�BL� \�W���X�ol����rŘ�so���5��9��o5������{U]�vۻ�6�e3T�Ι^2y�j�o<�[��9��@��SXw�bs��P:�ΐ+=哴�c=��n�aǤ�1���{ܘ�����3��55���8�g�m�)<�d%���&r)Ǵ�jNe'~��
t�gV�q��J�ɜ�.]1wCS�����
��s8�άS n�P*[��e�;MLf�u�1*w�3-��˴�`�-��ל����G�59�MMLg�9��מ���,S@ݦ�׺���yՓSXn�c�;�yӳ�vɜ�'�������0�Aw)=i�x�!ݷ�P������ܼn�Go�a�Xc������8��w	�P�箷��	�jA|�L���5y���R
v��cT���kĘ�g����=�!>U�Ƃ E���U@�VP+mJ�6�]������gkaI���5Wl��d�@ͦd��VsY��)3ׇ��t��H)Ğ��f\N0�v�Lf=w���ΨbjML`���fd;�52�R��G3��Vb�j���u�yg�=^T�խ�Y�S���o���P�N�C��vg[
����ʘ�&���V��]d�MLf�u��9��*W�K����ju�9߯}��U8x�wg�
�n��)�79�:bM�'i���a�\�=n�Lt��%�p�;�O9��\�t�L@����z��'��39˜��|$g�,UV�m�ݮ�k�q��1+���b//��N���jbz۬9�^cseN=�n�P*s);�eS��:��bW���y�˦!�T59�N&�!<�t���jd-f�ޯ'��Luv��R�73.��jc6�c�0Y�\����'�w�C����Rq51�\�f�^���yeL`fS���ZN����66k�95n�����Sd+!��� U  �@mm;���몀�7p�ZJ� 9v�m�X��ιՅ�yγ�d�E9�'�W��'+���{��0;�Wy�@�̤�Ͷ���s�q+�OY�T:�OW�}�fp��+�7���[5}�i{�퐄�I��s(�N�*y�N�S��36��1+�%�p�<睭����551^Ѽ��ט�&�B����lk:N3�a���f%zd�>s32۞�31qB�FC�r�|���f3,�7�fq�;��03)�;�U�1�3��rؿ! �!��#��a�
��T-*AH)� �c*C��~���R
AH)�}��Y5� ��î�1 �'���N�������wBa>Н�	��%I1���I�`MI�=|/ð�{UUX��n,w\����O~�$9Ր�kr�cI�9��y�&�%a<I$��I�$�����I���7x�v�@�'[Bj@�����1��$�so��v�BBnX��	�	�@3{�������S����UU�ܥFۗ9��g�Rެ	XO|���t�N��'l�
����$��	�	狀�t�8�t�ā��'�$���@�y�� t���d�q	�	��
�w�&�	羯y�,	��T�Nr��d V�( u�����[l�JH* �Ȋ��*  �@@�Wo&,
[��Grڲ�v�eʪ��Zh�e�N{��v��� La5	�,	�	XN���g���`z(Y{��Cw�W��<PYP��泵*}V�A��   UVF����;�r�Us�rx36g�Oc�����\a�ή㳤��Nf�P���哜_y��q��XovT��'y���8q�2��jc6�bz��c�3���ڮr�B����Յ�Փ��
�|���}o���;N& W��a��SkΗN��L��ͤ��Lc�fl5�bW�'Y�T<��칓՝�N66k$/h�O@v���V.�V�p����)$,�z���̝'հ�\`��2w�yq�ҡ�T59�N&� T�3-�weLN2n�S��Rjy��v���N���+u䷚���>�\���R�M�R���]�P�(js��MLg�^y����l9�N2jbu�rO\���i1�;�[�M���̢�{I�I��-�T�^H�^O<95�^p����
1UP�&��un��*� 
����*�w���Yܷ�˴{e�ݴ� ��*��r!�{��';O7�� �d�(�ͤ��_2擤+�\aά18�z���q!��
�8�]'T����9��;z��l�$IU�p�uI�V2��y{����=�55!ݤ�ߵ��Y�I�H/<���3E��ݤ�+��usXy�'W�l�r�������L�^�
�)1Ă�����<�m&�&�Y��O]\a�Y�MN�8�����I�LB��Lq����a�l���O�N)9��u�����4���(q��q��V�d��G$6�x³-&z���u ���QC�I����f�	���\a�v���p��N$=[�z��ν��.6P(�0��=5 �2u�P��1�u�&!X��<˛N2bbC���<���kRc��'Y��.h��T����`{'$����I��<�⪪��*Tع��U�5Yz���j�U �ۿ߿y���ѻomQ��n*  
�T�7Sc'�Sl -�U  Ql��*�P    U  VP �M�*�Z�e[j����b��U���V^��ȩ̪*���m�mB;s���ύ^w�Kf0�Qĸ�1Uٵ]�@Ƥ�uM���.��ݳ.ý�Uw��U<�dQTj�cd��3?��sy�hU��������
�  UTVPU�*���\$n��5�t����	�;l���4�Fm���#��ί&&$>O����<B�-&5 ��73;�7i7i5
μ^z�u���a������rܓ�)5�fZLk��w�ݕUUX�(�r[��:ĶOi8��z�zY:���ד�Mcy� y���OHVe��{�����e:n~u�,%s�2��Δ�/]��i�<=�H��-�I�����z���o7��n��ȉ�r��%�`
���_�j�f�,��x��������_$k�� �t�S�zL��m���R��_p),�j����Oi��w���
����^'�<�gס�H�B�X�,X�P�P 
�QT+(��Ys��U�ƽ��������Cm�*M����{J�5U���������z���N�Sְ�I2uPq����h^��j%�m�}��v�.hGS0��nٟv���([K2��1��z>�n��15��|�?c{��e6��|�崏Ԝ쎖�UW+$��OJ��ָ����9��+�E3���͹��[|�Ē
�k�ʛ���=�|��i�Y�~���v��l~��p�~��>����h$Nl�W��@UU UU��x *��֛V�ZGj:� ���l�r+s&��6�=<��u���6������ ��f���:č�@0V�e���O�mq�����#���{T�
�U��ȓ�.�p �p�1nRX�$�<�]�Oz-*y�{��Wc�$���/�w�ߟ��0� ~�%��U@dc/��1�𘁤��Q	�ַ�2P!>�n{)�� kԈu@Mkv��O��,����M���x���T�������z�V�܆ݞ����8D�dXb�nw6�PU ATWve*��e=\��޶x�<v/����Ww��G�ؖ�sK�){�2�`�Y�'�u�ܛ�.}/��*�ŗ	���&���	�䀖V�K�����6�
b2�]LO���m��UU�d���:����Z�7<��J� ��6>D�Bf��ݞ�ow�}L���$2���խ��m&�����*�����*�oD���bq�HD���q��O ���:�����c�+����ʠ�B�>UV�khڍ��P  @ .j��{l
��_7^�:۷���6�m�)o�f�6�����V&{��!��mX�D�����M��q�� ���q* ]��<������9/�SCUM,�斺"Ro=
�q
�w��*�����k�%�ɿ@�s��2�%��4N�U�� ey�,�T��w,ԭ�$�I$���N�#I��kB���=�k�=�h�!���@;VI[%Ҁr~��pcj�a��0��rG���ޓ���VV�<�R����9���N���n��t���*�"���uޑ�嶷����TAUT��=W�l���V[m�͔
��l@ -�TVUPd U 
�Um�m@@   U @  B��*�1�l�S��@  EP�UU�ml��M�dJs8mm]��V��ӛK�Skt+m ,lp��]�UWV�6[������*�`�m���;v�8G��xO^��n���5����wPmc�Twm�  T 
��� Vą"ݭ��"kAG �`
����\�R^=�%�ٹ�Ľ)J�u(����=<�
bt+%��`Y'	�Y�UU�m`��]�I����ʠT3���˲��&��������t�os���*��`������ v\~{�RҜ%��t���5!ҥ�Zs�-,ݲ}�����AP�� �\�pt�b
�q
�9*KǨ��Z*e�A����g1
`�Pl~�'�+� �2�,�w�l�9�d�tm�v�d��dO;����^f���R5UX��mn���@  
�e*���VN�X	���o���J�ݹ�J~w �
|W����������mcu\���U���tz�jN�~�	ᱴ�ߺ�ة��7a��̋�������Go�&k�
��&�⭵�,o�mY ��&���3��ʹ��HI��N̑�.�>�3��dEUTm�\��+�$�\R������j����%8�N��a�� V� �����9+��b�ik�����&Uc�2s^~2�'���� �*�Ш�b� (U 
�p��` \u�muV�v빳��j��-mEUW� �N^�2_5&p*�� ey����5K���H<����J
bY�P�H`61��Ilg��r��h7�JtZš� ;PL�ˤO8���ID������}�`����jɐkyo���piҥ�s��cr5~��?��"��|x��;�%����N�{m��ڊH�C@3yɳ��@۾$�u�%�H^��?.�������ܴU�Tl��}��K
q�T�m����٨���N�Ìu�	��ۚD�a��;Eq��kmQ���U    ���m��Sq+o�@�[Ku&5��]*���5�C���#<S���ݺ�V���;V�x��Q�U�,Ԗ�6���� _
��9?	F@ߡ3nן����֙O,�����
b$|�Ұ,�Y���U@-��\ȍE]l�@~��۹,)���k�=�h�D��VΙP|�x�oUUY���yb�a���Q`��G2�V��KA�n��V����}m��Y�*ܔ���<�^�e��A�o��y�/9��O��t�3�Y�N��:wv�ݰ�@  @)��*�A�%�+�(��a���U.���UT0����X�s+���	�! ;�ZvfU@�J�����ݶ������~Kh
���W�����l�� }+��R��2�k|2��a[sR�Z�1=�-�QY�k������Y;�OY:���ؐUda��y"�4�x����P��׵m U[L+�e ��)� ��@ҳ7l�@~5�˺�C�_]��2gH �!r�l6}�[o���YEl�J��lQ�j�����տr����>����-��k�lj�ΥT  ���rm��:�AT��  *�۱ua®��e^��*��� `   QT   *�� AUT �U )����&�R���؀ T� �T��*�` P U/e�J��[m�;��Uaq�8b�%�q�[��mn���B�\��M�6�:�T x<�w��q]�-������g����tw]� 
�  ,�eU�T)Z�e��٠Yvع �ʖ ���ăc��O=���.3��[�b6�|*�`w���K��'W	�Z�ƹ������DA������9�ǭD�������L	���}�, t8
�[]
�=��L ��l7�C�I�M��x)tt�B����d؛#<^!�;g���03-�j��a]s��Z���ԩ��M,V=���*���ęU��zG�3ȒAOFH��#M,oսO�U�^�lM��7� &*o�ڔu�[VΊG��]/k�n�t�    �� ���;�D��Ճ�U�J6�`�k������)D=��ۺ{'���˖�;��O
��dP=�oɽ^lC�V_�{�E q��ȱ��R5���\cE.��v�r���?E��%ˇ�S\�]�p2��$� @rb� ��&�w��� �m��*�H7�<0�� Yȇ��� I}�z�����@�?޴��f�Uٙ������� X֌�
t_��9�C��+����[���ĕ3� ����g�p����]�m���p��m�*��p�t�8Z�!�lVA[k�mP�  �F�l 
���nV�虨�n�!���ţ&R���f��2� V9�?���öS�ϴ�0�4	s�� 5V2�F��23�V��[ܕ9��$��6�bSJ�"bԕb��I�6���V�&,��#m!��ok���@���o7^j���nY��0n�����N�;:%;v� uU�d\l����7�9g����'��$��X1OX	U�5�\Hϳ�ܪ���ū�%�.���N��9? %��B@w3�ٙ,4sjO��e�{����H���v��  *�*����fջ�s�˞g�u'W�uiij٥c�I.;}����@�|���'�s+d-(�e���eS�/��
UU� ��
�O�r.cEP�*������<ʬpvKa�������ʶ�1ˁ�Zr󢅷ޒ��#�O�������$��n��(
�N%�UUU���2��e�n�Ej�I"Z�vc�/�J��t�m�ILb(Ͷ��l�$��Cjx~�n�����'ꔴO�1��p�*k���v�K�KPuV�/T��n��۹����  *�UUJ�PcR�cj[y0�l�;~
� ��˅jBn|���.��@s�9��JF��� KDzG∡s�� ���ڒh�̬
�Tݖ��oc��L�j�t���z�'��lm�GT�L���$g�pY�e7o@�
ۚ�������:�,V=z�[�@�e��>UT0-r\���X��J���.�,e:�@m�����H��_�. I>�����ad�pdC}�h�sϰ�8sC@%��ȟ�J��āz�����Ns�mUdUV%�����u���_~��  �k���w+���ڶ�  {u�;��dmm �PfP� 
� �-��[h  U  *Y@ ڪ�T s�m�T�بU�T+*� �¨ l�U l��.���2���@���m��Uݝ�R�Q��:��`�aIm[	�)�e-�U*z����Z���s�ݹt��6�%��YX�uղ�w;� @��@U*�R��{-���Ǟm��{�|jT�E��b×���dg�4ɻ��v� ��J�
N/br	t�D�z̕UV�-+K.VG�x���]�����9�$y{�Bm��B�֤�?6*���ŵ&�\@��k��TT�sEٙ,(�n{.�O��il|���M�z��J�q���5tt�Bp����m��(�e�]m�T�p7�~����>�{� dUUF.E��y�N�'����[�}��2�2H<�zs^~R�7���V���>�Z��hl�,X��P  
�j�HH �A�I�� &1�)#E U@ �$�$l ��IUR��@����J�:�!�Ӆ�q�IU$!�Z�3*�
�{�\���@p,��ӓ�]h�@����N�R�e[�'W�T#������bW�o�;�+�󬀪�,HV��Å�����ޜDu+hj����.�T�T�W}�3v|�n��O[�UUU�d�
��^}0��� o�.��r�MQ�� W�»�v���*�����$���*ն��޻�T}���o��)��t��%WT�պu$���7m"��<0`c����@)P�Y Tu�U �P���Hcn2IC
e&.K�wv_:�[w��R����X�[|���\v7�>�ex9�W�]�oL"<ֺQ�@���ʐy#�O|����Z�L�f���ޏn��h��IU$��~�խ����{y
ao��߭���H�H��t�wT�&��feW���u+����T�P%�F@��]�w�|�o/�����2)apr\�����-N�=����r�@�$��O��d��*[�v�J>�&��~��Ɩ��Qyy?!�w3$��&�`��HF�Α����)�����|�����M��sj����(5j[P2�j��A6�`��P UU S��UP�3ܳ�zշw���շV¨V�^t ldD���WZ��s$�������	�S[G\""$;m��N {��vOY����VF�1"_�*�wou�ɻjx`�}=���{	�<���F�.y�%^��k��]��UT0nG�`]�c,;�aM��q'*��7ωN]��ܾ��D�˺�w����T[J*���Tm���Gܣ0��V9RUI�5{�2RR��)�գ�ЙU KKl�[XS��sd�����;u$��S�|�pyu�dW�n���I����T��W��=��s!h��j�.���[j��m� @��M�]�*n�[��yx��	�U\56����c|<��V��[�[lG{}�W`ӣ�ZLSnH��rZ�է����(ȭ�r��doE���m����q���ddD���9�]Y�*J�S�ms�㻁5F;�d����_�J���F
{ܴ�m�j�˻Y�ӎ�_�j=�'6�/�0{'�M͵�v3~��6]���*���w��ۦ�	�q��}����uם{��'}�{@�6�;�u�]:�z���㏶N���׿K������'Iǎ�#��s8��n9�x��Y��I�3N7?9��Z_�UJ�02�.�8zq힭����5��I���%�<C�t8��N':��^��˽0�݋���'9u�8���N{�n:�[yˬk�7|��d�Ƕ#Ψq��MMu��}lW�b��$ ����O����}���������!7��А��� CH@O��2 $�#>\�f0B�G��d�
��� OL���\��^���%>s�~�<�?iϤ�>��뉇��t6|�@螥�M� I?���y�O�H|a��>�I�H��$ ���H���������{��O��>s�}a��! $������IN�'��Gð@���C��a�Ϙ�}�����~�	�9�'����ù$�P���@XI!#	O�!$!�}�N���>:p���y����Os�����G�������`�|���OxO�Y���?��c�@2I����Oğ?�����}3N�`P����?a��u!����?�=�����|� �|'���ȈS�??�;�8��~��� �$�C�B I?�?�0����B�G�%�GPHO���@$�3�����~`xu  I,�z9�h��d5��!�����rB I=����O� �|O�>��O�� �������H}�������|֏�)��� ���'�t?(I���	��ПL$�~p��?_�:>���C�PTd�/$�TI@����C���ó��'����;����O��s�C��y����>Y��!�y�NI(~�l�'� I?��O�d� a��|�?� ��'�B�_�I��OAd��v����!ߩ9��w$S�	�`